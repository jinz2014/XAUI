// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jw2ugRC1rTAP7IG2Vob12E5twc30vPb6r6RYnE6SRJRgM0GAON3zgleFY5Z04B0D
9LWJ0ushedQBQ+rgNaiWkxnKNc4B20MuNioiVkLaiAneRHZraK3kaDwDRgOYTuP+
yiwVvUkgEhU4xObKv9d3Rui45cL+zA0OHxbA38d/AT8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8192)
P++GybaCHGmrIMB2mylqs2doVeGlyppSgU2CPRQucmLcpLKPQygACg0OC0WSnLmj
XSA/KSQfxk7Umz5DmE2TL1c2morAykwV8brBXow3Pk2dI42V0+cAw3hp735gl2sB
SRcBWpYBHjsoIC+uC0YPbSgpnTpNSGGjiihoLAldw1yPk+CfHr21r4y5EusmAA8t
N+um3qcWUVwZol+wovAhbMBgZ4/4G4ANIOrQkpKijH9OBwcXhlprxP3dhOMQli0Q
FC6imgNvYWf2J2FIk/+GMxcy/xcii2o3Aduw4u/jP/XHzX8H8DmvVFnbwPjwbDv3
GjJv+LAx51KmGEv7ibFAiMt5P3WNiPQnEZy9xtuqWdLN3U42/lOsEXDdxggnM1GC
NWTczvEKBiCQ1CWIuYTBZl31hfqjIMtH0ZWKzYPdvg8o+Aw87LmTJVGR3iFm3efB
ac+oRFRP77ZOP2RUQIgqyhOBkLo4UkIhZTUvDy+e3ajMEX6MUPfNd/8GFHnugLse
Rt1O+t0+Qzz6QnfH9NhOOoDpJeFnTNg1tAg9GcjodS0GgzMs1CdjJMVsN0lpqlZd
5brqjxmpo4fty4IR1qG3ksxA9lq2gvFaBmxs7yPCaL4QABq/53csRTz3KvqpiAgP
7cEmxxd088/veDTrS2RbHrWSd4XaqmdqJ/Tt9cn+Cw1V5Lnv4PjWL/fZ5/JH+qMn
ultyjVS+4iP0+TjPytN6RuVvLQrNgYrj03XUgh9Prhnl9TaoQC9IfPJJLys4XbpP
PwPJDiWlc4CK6EBMFScJhOuNiaJegv08LYVGKFjAaGhUyXaJ3NQUIEHhEIM+gyVn
LqT8Mv//naVmhJEkXip6aEjEPI9W/hw/iPXjiIqW9vgVl2MnRfGEBzuR3+i9C2TG
bPDDu95zFOuTzHcPZNgcMSXWHYBZzguolK792jqauNCKYjn1tZRR6z/zqblGZDo8
r0s8QiVNs+ZUW+Lhk9f/DT5AwUUysIW+Z+SVFcB5MV50Ciff5xJccOVGXHdayIXv
FnZioO5NLl+SJinAGynW/9ng6fOWEICT/HAYNZR+UpVHuWhfbHqVJnQ6KI/tuw5y
y7PH3GaCMGjVQl4ZsifqCcmKscGMK37sPNamB+BzI52F36ZZuyTAH8D/xS673QNd
dGlkQu2uq1Z8Ly7tK+75H4qswuzRY9ITqfnAuSMDS2rIiDzBlmIouiztIZ+vYA9U
LfvfHDMYulZYile6mqeYI2U6ZHD219xTXqnZWpIwhPMttoSmjuf68LYut1zClQ0d
rPm8WN098dFovEtZl9rnf9h1kwW7BB/QSxmdDWfO4WuVphMGTpBEnidAgQQoRHJc
s2IaCJuEUmJO2Qxl6PfCLzwkzV5nn7JpNBrCJB4vQ6WItUWGG3fgbNWwsucoF/Ca
zP7d3Qymb+QmfieZaISa/t4pyBr0Dc1aFhATlO2uwD4EkGPuFjG0Jc1KewrnTgs1
+96MWuo1aBtMXPdz2r6Ne6MCRZhLnNwsrGkNFmvf2W4GWQgAdcD1Em0qNP6T+AJy
jo0D+u4NIjvm6AVsIh5xKydYhCWlOqWgkXhIj/V0l7XxGYZRyY0gu+Z6Tc4AUhW/
dW9Kzt4tHmbGa7paS76NvMjXMdyfe2sw4hRlavKmCfYpvhDJ05bU8gExaD1ys18K
Yl2w9m9h3TfCNNLLY8lujfeqwox8FdycqEP1nJIAJg19NHERloboyGvLuptgziKL
hjC2B41p0wSGV1DBsv3KGSXa61G00nL+xfCm+gPf9TNJg/6peAZ8sdKw00DODFq6
539cJn0CGBmZebzB3OkZex/wsCLUfjQh0gk0XUmQL2eZuOnZahltEDUIEJos+QYW
eLIWFLy1bvcPX9M49bwwuppW2BIYs90C22DMxGhLuNjNusYYQt3oe+A2thNhuc/N
becFmm5vuWoHrZFa16rNHeRo/EkJbqFPvyNaTil+ES1W564T2R3Uko054bGFbSPE
QIMKShQscYPYNTqTmbCGH/wp+IdV2dkJ6AAkQXYiN9QAHBVqeVxRDywiay0IQoD0
tP7eGzbm/ME4k2GIiSXeWAUnkTPOFbXw1tbgdyZ2EAr1ZQS+w4/C0C6GtHLDUJR8
uMh+bOq/yzpv4ec+MSGtZPS/6fWp1ylGKzfPL0APhCzfMZGHaeq9ORzkX/HhSEDu
3fcsfXrlQKkq7RcuJrkABlozWwytLvHjn/jNRpckAOC1SBA6rhr1tRJ0u8/Ts0R5
ptImv3ES1tzlZ50KU2b/HGjvXKCfDdHJ7PTOwa64m4s+Y2M9TUqeedMd2/UUkTN7
RJGcWraVSjfIoChDd9Xzo6AMPFTHkEmNolV6y3TBYDhOHHWBhv8goyETU7INZXCa
5Pm2xFkC3LxcSrQ8pqalVOILUAP7OJ5Wd4n9NLfwOXZoauB3XPZuCPFN2RJC3AXF
cxwtsCFMyGBL94Px305pbP5nGOby7cNjGCBwH6KUGcPFE4xKwBGiYj22d4OwwOUI
VpApD5XIkazZF0GUGy/uuA+PayRPvw8Q6BuY3z14/gJ/8U1o+KWTlJoRghImyR37
JyjdK5Hrj+gFq5mRdNYxTHb6SGYPNpZKNknzuFi9FOVtT2xryZbwufCZQgv9hLkH
5z7cuH9UvDmTZ3dhyAS6ouRoxYwcKoNJy4MIgcPkfIzSDH1K2+aWbx+BFtYLhpsA
SXfjBo9cwd0kHJzzjUGjo2CFA6nCduVS6jHUkCQok3wU8tG/40hwXlbRIJm3iHaj
TmYrOHzKxT4DliEL2rEv6+Tf/60AH5McvJ3aBW7Or+xT183PcjmL+aN+Mx0TnQMN
okTWeJIf8Ib3gbeown57Iek7T3IYFxVmMXKypkgsTlVZmnbWp5UH2cqP0E9T10jM
yszyngVawnauI5RRyvUBUgKKepu7+ftXegUFef3uYox7U2vZbHQbqA2q94RR4zJA
sxQOltb67Y25e8mrQgFenScraOc20slIzkC4yIkyAGXF395snl+EFWM3V3uw89PD
VS1jJofope66ieSN8R6Jrn0UoaaiMH8PgvEPvEjDKYIdwn2Jthwho8QDEEwtXuMW
0GMnsT6IXJKou3xqMUIwlhKP0+ajdITJi4fL28HyqvBw49pT4rlZ0UKTkCRfshpv
HPgB6bjF373Z0Ales6iz3ipWyac6yO02/8Cpp2vKTCSgv381V2fdwqcgkLnqXgsH
PZW73KKJLj8S4vnkJtIISfXPZpkercLv+lN+1zZKOv3cPiszGVaklYy/CG6UlQjh
aKLaObowJLIQkRRvDfep7vJlzboPRZ7ttK9BAOhNsAzdPlmiETXCZ7E+S+gs6veE
w5foqgNKjQDWkGrD1Rw+YcMaDywec3ySS5UPSS6Lg+JUZ4RC3pOy5gxro9VNUoIN
wAKi9jlVK//wa7yLTXNypU6UIkEQAcS5ldqX3AEBDAg2lkTzPYHqqROvJiJRf2hY
CTb1/Ezd34gnsN1gOkTfNnds7ZzVDbs5HZV9973EHYj1u7Ph1K8ePAYPzy+uXpXs
biM4fMGAgKATomEVvgUkZTsvj5i2KAiJ4B+cQjqQK+iZ1VDmDnuQ7CROe6Eur8V2
0wy29Cj6bSKsEyywivMU7NPU9ol8i6ENH7yCj3f1Ll52IPUxuo+rSoA/5EHetSZZ
dsHT2FY8lKVLTVkbZSCtOkZeEetb4nFIlicSwoqJwl7kkBio5lSROde3QyaRhO12
mqwQLo4AqfaW5rIBNVnLD72aLZqzDVI6hgeI9ch/RLYIeiu+mhFnlJWUz9NhzKmq
GekX0wDWJx11iXKX7GaSUVqtD58x22vvGx4RFZuwwbPVQmGUjn7F8LbT1O+BT9Jv
49qZrQcDMxq4bivmGAul7rnJ+kxc4aiHIZUNNGW78BIRbu8PQVqUYHGYt/SL7Gje
K/QE6UKoRPzstUmqZKsmzkQmmB3G5Bs+W7dzgw7K8nZkqTaxehvhL9VMoR949GEk
dGsh6AeekR2qjikwgfwgq7t5EnBMn1z52NVqNuda0+82n9BYwOzJieM5yPGgRRw0
qfu3hMorBSjSvC0Bsa1Ij8FEQvqLA5kMNi5BejP3J/dsOhVRNIY6NRk6ngpjJDzX
4yoso/3St/TdCi8BhjOwuE68LIJkcTBfEqXLFY+v7gCgR3+hsXPC62a59E9OEp0t
QZQd31NGWaFIffN3bIPjBA+qM8/Se8qbGGDx7dXSxIz3VxPu7mu9Sxx1ZeYOLNxK
kpEDiRvD7wUwokLKjJP8qFyG0TFYBxFyII4i4aQU2uML9cagAsR7anDRt7NvAhc9
h4UkKZ7AACt/49y4nq4wdbxa6Wyeccm6XfAWABxTDL9+9oJKdB24kyRQ1a9JSeFN
pwxijgIfrNDaTyafx+BF2ajphukILchBk51QRvu8ApNbI+63nUkEjMLgi6kQZuov
npfHL3iuuUVyeCzde1AI59B5K4/gC8whLqy+60iPh2MIUHHHc5pY722GHEoEC6xF
IN6DYTt0+l9roSqE5lvv8S4VZHuxyizE8oOxIeN7WahQLnx7D+9eq95/aGi7TOYW
qvR/PIYpDgrWQmUJo2mTaBVp2s3lh5gxePj0BXThhn7uteDwEoeIP84bLB45zZ0r
tp3ZiUue/2xY7TfdOY+4gM5bzns+STWB/jezWB7t882Puflxuu6KyMfaS0/TiPgQ
wgQlWME8C7KcENwkC08kcPd5LakrXwbLivddIjepi/8Yqha0wNpauqmWAr1tWBpN
M/T1le5H/DhHP87vHs4d3mU8d7ohz1/l3/NbplzaeIZkltdXHrra0YJoCtdmk4te
kV4SBJUNyxQN0bicj7fS375dSq33RlTTIGKYgHK75fpN+uQPNC+qLgbBd6ixKdgZ
ktDc/THfIyseUW16Mo9GXJISg5Ggx/nCBfVC9q+2+NB4mIuSLs82VbWwbHnJkXnd
ow0Mr2UMQ9Wm1zJoFwjrWWKdg6nm6AXJB9aJ1YLGrQALI9i7bILy88tDROQRqDcY
PTCg2usrY1TWDkQvRFDt3/osWhh4WUEwKSg/TxKg00rinao4nXBKQyPDCjdNKpKT
Zt10+/emWRWA9OeCW6ZB8yCkPjL84RdL+J3PsER6YvzWqFYmZIksMiu8Ms7m5l/e
WSN/8BHMxvFOKSq8bgPQW/fKco+cNeE3tZIKAYHrFljpIEbEAvi0h5lTnWzZRscG
Z60To/eHod2ahncHEc/Q43BMleiF1cEpMcNfuM/AM6IhM1aF59Zfm4iMjhc50mAB
MJzVA5nwEDRn8Af2lJaXpt5ajH9YW0trALDBq4sNPSLiy9InteBcNoFEnyFJR/nd
AdXEjKtp1L9eb8cEGSgfYc9UMNJCc5TONOS3RO+h+EG+5VTmP3zSzI6N/iE6yOLK
UgBr7Uy77uMi+fVlMUluiOCalym3+h9E5xopdgTUW1SQrSLBxuOa1pDhZkr7aQh2
8Nug6sDyScQ2BOt+EbUeb6mB7Ln5qxK5+cMqKUAKOj7iGnIQx8GTaCf5lXkuIhHQ
7C0yx7UynNZyuweL+TDC0+4VvEbchzJ48if6GezCYb+kfRyWyR+GgQ58fWWQRkgM
9N+Nx+y8Y9Izp73XpJrmamYsj3SVlWW7rWBpKfBVkcPivtCxhhotlsj4gNJMKx1A
85gtOWqMtI4UMFuoN3OPPc9J5WxGiEh/Mjon/+3SPtknQ2ZkmBpMHMEV/K18g1qU
+9PAat7wTQMPpdJK3sCBBb5/9aLSClQ0QjYJQxrnNSFASi5VfSPLm2cIei3j2tzG
5tuGGiIn+bkvOLU23sMn2fM6JTfn6JNqMtUQ3N5AfpNdk4KuuH5Z7fAPULTcBl/d
MLHjnhElx7QvFLWsn+wJ1d8F6WU8ChP/rH9pEkJxKMIzkT9y1l0a+VgR+oAVL+YO
ZuG9CrT30Us0SoqBpFX1z2/kGspHBmFi12BORq9UpSOP13MBZApdyj2Mdsaah1WP
GeSbfpRBNBS7UFWzCK3nd3rXWlzuNajgBrBZetIeipx4Ju66vH1rEw/sTFpJ1O/a
Qg33lOOoDxGghSFUqn4jUcmcivIDAP+Lr6UJrtSL1wIPKv77f5bYza08U/yyUfL3
tCTvalVXoMW9DjpdxnRwUN3xSbLp9RiHWkrFRtGWWzkBb3GM6VTmol2b1LfpOZsq
BKoeGjDIuPWM9j25pp6QrSXLnkRLfbuDw/M0pk/wgqSx2lUm+d6P9daomGnceloy
i2VaL20ZucSDut4eBdZtoe+iXVBtpOTzFERx4ZkNfWwiPQBcLxR0/0BSg/kZ4V0d
dtWnRy9HOsZIZQst0Cl0tLIwzZ9xguC8l89P5m2H83lKy6JeRThNoFmMAgfqpHin
vPfhkAjVL5dAdmuqXeIH6dwz3HG1Nogx8cnijgQ5nEJPXCarZ+AtkMG+Z+EymRQ/
7wBBHfeoSDtKpiW68i2H2I1c/Jk9yb9OECWyAfL6uCAgQKIwdU+I4Abj/WlSG3Rz
GO+aZnJUonHLovKgR5tO9bBIvpqSW/NjuTUiJyH6Ami2n1ngNvv0pTxgLpRCGJYF
hkY4a0mDBP+3qgSpF2haDt6mZZmnLhIcnRTkudSplXY1In164+DK5h7hJ5VMFuof
vyYSh0GEOCx4ihGB/tsF+ERmuopF5PdJWagjGFWz0nuKcG0Wk7cf4EVhRP7VBuae
cgvEYxmAwhOK+TfVzijt/OmqcPVVrpq653ljiCwbCLQ3QjSEzOKWUNik6cFtaWJX
cVYCsqk/j2oJtK3ahPXHxW8dPMLbLWw9FmwnL6h/uts94Il/m/8uO8312y1akTUB
L+ayJwBcggra5eiDhCuwBpY/5wKAP4CYXMZ0rasg+PztQuSedRQU3SGGqYX2oYK6
fX7DdkEpd2Kz3KP7FQTPjFfbR/xPS813UEtklnxrsz4JAgmnskn8MgcmZ6UmS6K/
KUKWlWdRgNsKPs7P/fDnZObyWQJ18o0bxcidtdQHwbMjx2hJIEXZq4RzLtsKhf9r
edMiepdZL4I9ifaxxaimeFGUTK66rhflAWGJMQ9utlItGqGvs2vlXALzNINAhSqF
IWyej74ZIsN7lmfolTeoNQeHYn4TdLBFN3NaqTVh4umW4BIUrbjbWz4WI84fkVxG
IM5gsYZYiR65qjEDOlXgjjSkry/aVRkxj9ZJ/d9lMaeqwlk4HkZ2xC3Wf7BAAKNz
y81uaJAbZF4iIRDF3AeqtrNWrJc5pOUODx1taR0NdCLs1nc6O9ToMI7RbOiD1/6L
4icRK2rGuwGA119RqT+FONTs2VahJc3p2P+hEUawj14gA6FGLsNewsiR6+CEREk0
HDeqDP/ARp5AxXXOuG3GD5y8aIIIickIX0CZbBThtZHjM44U3xCiSrZ11Pscg/tS
IhZBR7RbPETa8IRWjXPMgKylmTlD9sUwvG+XEtaVdywz5lUrxhIE/WtQ6QL0QIlP
uymX5c9Wf9XtR8B6IuYDEdNcJyvAE7kWanvD8rGhwcatsEdnwYLKf1KtrS2czHI6
869R2dXP4dW/WgJ6TC8sF0QEKqEE1QLYtGI7ioxRlbRJ2n9SFsH99H6fVAp3DpDg
Rn5QqIhFPdRdT9k8SiDQTwJp4H1S0WQz12SkRu9X2Dmdfz3iXEB8jlqWjXFhpBFN
3l/eK24OnZk1tqYVLp6kHFXwy3b6r6Oc2oMQKkB2WHOegHEr8VLf5+0u2MegLZZ3
sUtePAB7bdGYJZK4ejA6D1cQGP9sR6boDLVO/wVVWolxNLSo7RG3kJzdWx5f0ur3
M23udachmuJn6C80CMBLaeDYSnYiUp0x8KDUErJACSktLmopjZx+ophQG5h9n7En
BvLZQxeKtRn0q+E+WRX40TOWdlioNCRkMVNRn1MhP1kUu6DsWno9FtCCbloLJeQ3
fxfm+yFJ5t14gIrfL6ygmsMpOv3oBC/Y39KKV8K4uXbKwavlFc7ykzTR4CVssghd
9EyU6zbWH2E+v+NjBXM0X5GuVNKDMtjtyGh8XJOz6Uz3hhJWrz+XfrmsQbAucn5x
e1D5hi0qBUGKBh9wV87WIkY850aNtJPuuUgwFImjFhiG728I9Zk8g1seUo0ZPprW
LYIRIIG3YT8L8FVhSZHNMB+KB0H688JJHSg8nF/iom5tHIyfd06oT0NpXYB2DO6P
+5UgIlcGrIwCFdzKt6bfayoGTbaIXvrYTEJ0sK58OYzGGLAtKBPAdyLT0z3uaKDT
OoLUQRHdAhxpRgJo7Z5gcilg5njuezAxCMV8nomCiCzzfVTESitH1oojUWSfLP/F
v5wtryjHLRcuh6zQ5dbBYXecvLpz58M3lyWDE7Gr9ek43h2E4RgtIFhWPqxMrkw5
EJ/GLsKytY7tYumUUak1OqtJBCTZv8LlMnhH52YjjVpXVCIXQkGddFggTGPu05Gm
xl/uoOsMyRUnW+gEJ3fS6O6/LbXW7/BRZPObKulg0rKMb4kxQPA6OkOobI/bTMSs
4y3GA0DLLMcCqwsoBhYilJs+ubyUNT57biu+h/4LQttZ5xAaVDYT8Ksoj8GVliT3
sGg3dWKk+Y1UX9B6tPyt3Gi56jNVFMivBa89rslR8tVt7cK6LraNIdDPdiBRU8+8
oIBTGjel1/+ZT+fM//7Fed3uR6Pk0er4ElUGxWwfohZ3drFYWP46ujWsM/trVHi3
gyvsGtbjOtkBs20L0BU2kNwnMrymhDWNQ/5d53diue8oruBrWsCx1kUmKsg3Xyz8
/5dELxzS0pqWeMRhcdw41N6SjnqvUo+RqAkhdfJyKA08f9BcvLUplrh6hPG0z4qP
uAHnHfNpdLZ9xHhNmKz+d9IiBMKYIZJy3fTMgcsqUn39TfbwFxZcH+x1Y42pbZGc
t7PVwwD+0MHMKoC6Hzb4JKiQqrDKcjGOJbbeOKkciRvTrZ6QgYc40JSjUwY/40e6
9gbx4mHUI8kVVFRLYHxwt1AZGzCkQsemrMmwmJMevoB7a1tt4J4/EIAWNz0bbEY2
1rD6QRwdsyKV2DULMpGIK6pIFfZBjiczMSRrZNhASUbjgN+Yf3WfAMVYFeLz76w/
3pVNAvPYIjVTgV2WXj0FbDE6nO+a5KkD+8TNsAIxeYKMBM+xjTVKLk/1sin92n5c
7pqfwXRyTiHvtBZEd6tCinNVSHU/H3qwYji++V27zdyd9hQhFTZQChx1eQeBTg96
tDPSSHRUsR7ierrgiR8hC6WS7uKd74CoAFvbw4KwbGGGaCKmxWwmpHxrsbve81Ns
iznt8MihXFimAj4HLEPGikwlbEAaFFqx+6ku8/UkkmTpgS//flRLfkHY2zOl5BBl
y3Zpqw7iB6s6pm07l5fIKKwWjpvMpXpQuSKX8+Sm6pNbFjEtb1MWSI9nhwsuydys
STsBjjapzWW8IcA9rNJqfS58796lKNotKyqt+O8Q26KjQc/etyw4bIMDsWZnxcMp
pkdKGKwQAwddS1Lb4VOyIxpDWQza1lEg0Rn9K5ZgeKRb+JEKSes6IpgwtGQPV2Cf
OXdigu7gnb8mWROeWZCLFN3Rqz1+66CgBYtekTAwn/+1iLBDfzvaJPQUP8lKxyjs
0eEtgNL/IKFlhsHhEA66HzVmmXffP+hi1+OYpRoX7wm6C+7leekSsZj5r7LyBfkQ
Pm1tqJc/tgy86FOwr/uzR+Xs8WTBb/wwes3xFLvdwcIvlaEXdiPFy4YqectZT/Ok
A2DhUWDauBry/dPXDw2nL2U9ISjDj74K7XlPau70Esnc29CP0GDJLgm33ggkWpsa
bthmSBOWYmxytkT8K2SvqGek4S2qRcRd0fIK/878wdjhJ1e1WHrgSArwkcHttiaJ
lMrPJ8cVGH55tWCNC3Ed485wWi/dMJ/72XG1uul2HRW9btNsNbMzZY3Qy8gkWwcG
8FlBQ/tKLtX9WJ3cy82MPt7ZfShbUfrhpOQplf12ZAMglvWpENmlvsnZGHZDBc8B
umZry5gz2JlCRV7FjW6LocycmNylCptbMlzyaH/vPmwY4Nbrk9Ns7OYUs1I+lhrs
TdSUW0fph5ckEy0b+ON0mvIR30lJsyfwaVyvyfshM9oY13HXOIU6ABX65mhuOimb
N733Bgodx1arM5QttQw/CDbtz4cvWu1vh0j/OcYaLJ68lfELsa4Zy/97ffYgN03U
H9qO3O+q3XwGnne+a0JVLP59ib3xsVLu/lr2gYWv4Z/8Yjy6VfsS8RvADstFaB4Y
LjDnrZoYH4IXokEKIrOxif1S/QL0kuuxdbFFo/bXlIaJ2U6We+8KjRDcA+6K7Oha
J8sUlezI7/IOpBbTT/5qpIBHB3ol9P0mVokguNe3lXCW1puJ2IAecu62TYcOayEK
/rtW2FgSLV5xNeGzhR/O+2y2qr37tDjfSNGiKLTZrVsMTfWD+Rt+K39WhKMyHAEn
/J2xR6aBeybshuqWSPIFW5PY3oW3oCyfdUgB93nQgENxlS8q8HzIjRHSnilbbvOB
K31l/NsKP7qMH01fzCQzAXOLMvmUFcqiyNkzeMiNg+Wa1NYkR94TDDJk0onUm0Kx
D4IN1XQVG88A0waOeLzsj6NExwyPteqCNp6eVDC2O5nSvmX6pTGBI0lOUj+IIP49
lundbVuBgoUlfwoGy8ImgzlFOOsPlXpbDZOazodWfsmn+Offshc9OQYIvwXb8VJH
Z3Kg3lyKKm/6haKwILzm4ja2sl+VJZ9++03ScATEMIaRQ9nYKKJ+CtS7u6vsrcTA
wXIydKZxNTZlvO3IMwcP+nRcXwYN7hQEDah7UZN8CFybyGuAtY1rQebWu3x6qVOk
rPoG6Nao10sGPKhpoXOzPksz4VB7PbqPXS0kEy5zDdT5mf99fpNtW8V8Il0UAcUM
CESsKC86L7qUFm/pcNxH3kgJotYDMybs3Xss6vCjTJPuVBUTHv3cT+svKKpBG+dQ
DkiAPd7QN6xugXPl5OXrTraEVP9ehkHcRHh7eGjXD3U=
`pragma protect end_protected
