// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:31 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k8yXjAApLaMXEC/jtuQo0kh49iUa69HoHrDSoLupM7H8vWN5LjdosdiU84EZqlsq
1u4bstwFf6ByXJqfSkfPXbbCkdDNC4rYM+NrR+jpnrp3pCDgJ5aBC5Gb3JCo+8iS
az7wCdxQttRTCHzR04ryzqCayZMni3YcIaVx1pc8HfU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5952)
pW/KZEHGUFm9IcMgmKjWevkrVbtGodlF9I8gDfPAxke6Vtn2Q5oL1TGrZcFfBe+B
246WfZILcfrxr2Kr4zAjU9+51SlU3mpEI/R0BUy4KMnCH679M4a6MD39cBneELY7
rk31rr20DtIflYG8HTJlXAuY7movzrSrkCZl6QGUw1SDDpPjrc1UOfWrAJ0sY0Wi
/sxHHvKFL1TugZuB3qjBN9shyk7XQyQYKKj2UQfnTAoE5f6INF82174mLZ0KbPcI
gnpXM4Iqn/w0xjUx33eIa6YRjJfY11nDkSQ/4JOrTbO1iyCh16Pffjh66KHuZfy3
h03JEorIA5MaXbjC+7yZOibEW8lB4sWWWNzOX6Fh++wQfaf/+DLgy4dH0rlOtN5u
1fKKZSOQsij57SNjv9atoVHRxoysR5oPnr5MdwIm5SnAQNm1Oi3lChLtk9BUYcgv
w9wkoFzz3taJEsOjgT3zjfR/FruvZv01fIj9km2BRWX6Gs3YCXvBcsBJO8O2QvPv
MAHFNot4cG1Ela6qdcLLMDt2rIN/VzIzB5UoLomEvKaBPEPTwjlUM9wdHbiitKvF
R/amtV7Nk6Pp6RIMjuOwNA47ycVbUsNxNVm5USJ2RrXBgNW4ZiD3XEgMVx/NnqsA
SM02czQT3D4I1cf+mPOZjkVLPQYZTVo09z01CPujd1SSfp2zVm/G2QVva6VGC2Bj
wL8V2L7Li4iR9i9vHmcrvgEBqeK9bb4iIH2c/4vKOYBAaGGg7gcA5YBwTGsbeRqZ
uJPKa0t0rmz0uCkmPMZ7Ho8KCQi8Dex0nej77+iimDC0UXiAXkiHPkZeV/M++FfC
sVsdd38ESGfCTp+B9dtTV4hrP+orQfJGSMlMJkEjR40fCgG60edBgWB+PgJuegDX
pOmNb+dYDNTfHjLN4NNHwNF5VXZyH5I0L+dcj9CA31yScsadSnzpOM+TaZWW2uVP
SLF+9+Yyj3eDzNQi75df4pUx+bukgl8chtJnwjK7W+m2L8m2CqtuCge4tnuxz/tO
m+KxR+I9+A8vMIHjFk0UXRBk62DGKWeFDIhPvWk6N2zUaNteC1QPBfVT84AVVbk2
oCwDgyloVpMujxu5Of/I02X5PIH1r24wEWXDH+4CHhCJrqAwVM2qNkYG/rzyTkJc
Vr5LX4K8lieGgLEx9UQYmV36GhDmVVQhTiDnrIkkKvI8HK06HUUb7ucbJZNbe2A0
m7rFBwalndc0siUu1ps+l6MZteVQ0gUcWUXzRjbsHAyhnMqTyOfoejfxh78mOVMX
zPC5bNkOjXddjr82ct0OXPBfzgAEjfTos+ZQMLNQGs21AqjuNJa5XLe5d2ALLrz3
IM1xDQsml64ynKkgUMCrtGH7VA2MfvR/JFBkCFCz0uDC0RVj4EzkKbMXnbRrlqzB
4ucAE5VYKw8xIQtG0c+IWqkRyF57OXpdFvD3vrxbkFt/BvLbO5PN5lBhMMUEEKVp
vqeGRXjwujBArFuyoSMC4gWabt2snpgGJclLEHlCRR0WeVjksOtq09NNfUxnEj8s
lqoAvpZ6BXW3QMOSx1KL6Gu8D77dXdGx74oH7LAaaEAAEQtCLdNqvbOyDyzPOwhK
zSC6AbUccDyL+d5Wgnko27Rkhu+w7B85kPtZScD0f7QK41e3X0dewFbE3hKJ5c3q
XNFE7cy3YfrvVeoFRD7dDs6Q/ZRr+ZhEh0dpR3+xEHhbcvgywktleKKmgDWTp9WU
nvoPxjS30FgFXkb8g94DqLNnRQEHeWraezXpjrXTDarzAr6djzIS2GaNN/cTzqCB
dQOr41nSNqsLpWBm/7ag3evVbkXltJ0gxEUz+GzNSV6Ln6ozRfik5lQIHC5jKJDL
tc5LiiV5CmfVThHywTvzLVWVqgZDFEHwqSBN0WNgjw8XuS+20KyhzrTrTJWoPhaf
uoVeMMo8JnFGgFzpnZ9F8fBs/ZUnxGIZGHHRDSBW1v7EgnbgvLBllMbxCTDuaCSi
2uHgTTQR7L160C6Fzhr6ufr16GmX+H6fEeGXbbr+M6fvgUOLok1HhTYdn9O0NkH2
mVNsbWMW4dYQmwhJJ4CTocY3+GGPQ2/ioKhvYe91Pbtoh6uxN/B++jpS/OdVOPrY
oDon9NVhaWLpYH2lfupylIqDGZdBcntsfJm8jqH0Qd4IsJ+Y4OzybX83LteEMkMD
RxCRifxaUUB3/zDOhbU28l7IAzxTExLiEjijPoWIC+yaNnln/clNYeOiMdWQUADc
824nLWG9Bi72aAIA1685p+U5kewA+inFLVlNlDsAAP+Wsyieqm8xgz0RPFWP0vYT
jbhaqePHfWDT3AQDiFvTxex3B91tndUr0SOicQq5IQL7p0dwrr9v3b38qjmZo8Tl
/wY9ZoevuG7ux3r53TlBfg9NegZhZBea+Hbc8CQlSOHT58w56V4MbmLMFlN/zLuL
RN3KXVCCAs8igQX9OiTeiJ3mPvN57X1BPZsZnMepzQr8fCl2EIiOUw8mQQCFQfx3
k2XqC0unqHge25EFMdFZxCT92unWA0geHD+3kO11G6+gUlmSpth90U7VozB2XsCq
WxOuuzuojFcgW4MYoCKoDIh4Qnhb68tUL7Fum2aMriaKvOfoKntcrEeBswDl8LaM
3ItQ9LM2NYVsEeywLvw17lhZdFoXF1QeWW5UCzlaEbsDWF7TKIhzalTID0S9W9Zz
crLZpBBTG7YeMr9NCvSdGKQTiS/nufinBgZPeTlJ7XrCBmlmTu+FBsI0FL377hLE
BLP6H40AndtC/CN99cM855kIWdosRqBShTcTsQ0NzXgKhZ6vQTqOPIjulDiPFA0l
KBFzayevsa6uwjBlBHro+rbiZDnPgsTv6qtCfZeJIT/dCgjh+wzJ/dRCZE/yXC6g
e1AOVaDeo4wRRrnHzNVFjtlMUVnR+aF+3X/9cZO0Y4gzLbSbNeyHgOyRD1msy6qi
LB2Wpl/3Zgr9HjZoeh178fwecbe4cehCyjFI4zRJBC91syuvCK3j3ICSDsRth9/c
6arBHq80kWfs1A28/RvJM8MiUszabn34SmkGjdicfx8QvfSG7XA4EwocJ29gUM9v
CppJHKCTKtq0vpTySCh/JN6nNLGtZ1rp3insJsQUTn6s/yWD6SH+OM2yXWhL0HrZ
scOJuyjvJGleMBu7/fimdhiuCspz8j7pTn3sEoYXhQqJeclKGp/wWd9xjAoXnBVm
Dcc8GuUtl1Co+0OhfVV1WOeXL+rwVpl/vmYhP/CsNeaFc821mQv66er5UXkMCPpI
Kq2W/x8U2CeIn1WTou7d1s1jahY2rrEbIBYcktGN7Y9hfl5XsFhGzbuFWId9LnOb
qVvwtJK5n2PPfD01WMHvSBet7UH4fKnENmJAapi+gQykJo16Fr6cg/9n1EVGwRkK
9JmqkM2GCkyTWP5EYvTlPV8Be0dr584bQoKJ52tvCaqYYG5FnAvx4EzjlXlAkZBu
iGU7k4Vt7OWTBFZCSq32b1j2N+Yu6AdUbwYLmVaVqmTazfXAF0vkYTef0YVdj2th
mU+9le5SA6VWw3TBxOPgCMA3D3gGbgF/dCEfqKvVI1SH9G6JoOHDRW+og3dBqXCN
I5/QMyeAbED7kTeRtW3SqqSbPp+imDxgQWqqpZY1+hIFBEXp62aVsUVPNCCfxh0v
xRFXvdWcDjXIhEnLhaL1B2IPOhFFmk9PpvASTe6w5bGRRijcMvUrc9d/xufbtQak
wzcCvwyNTKILiQKxvkrW04KIJN8d5DJUTl/MjVlB1roWh+uCrG//ksqf9/Ra0jYV
dwD7T1/IK59U89KKGlcpUtanAV8qngWJyfIjjxCFB/FcaotXtNG04oNmFchmxEfb
2m6e7mY2oG88On1C85L/tRjLMgmH+2xyAeU9LUvGnWarsc4zHHvPsBOSl8ZSKU1i
Be7Y3LZfA6I85cdDxhO+NyxC96tdy02yuGY2fqlLYv9ghVMbPTVP+2pPR8yErgPH
+N0HRCmb4L5Z2+FFqsH2uPh6LNriGMIYPHuEDpZR2Xj5sbcHaf//8OrBw2Vr797m
J/+fMwRxRscYtvFhXan304Ar2ewl9PWlpV2u5lc1YG4v5MJNSsGcaf38xUqWNxnf
daeo+QOX5mTxsr+cH4NmMRzQN0cb1INdVnY57KwZIpqbeN2CR4xw7jszDytzqBhd
I7wMCDH6WVmHnOzGAqms4/4oubKJVg5+vBsYyTePX2oKqib/a74Ka0tgPXfa+UiT
BcMOl7DbZIBDxEg0isolZjmJVKklBjewHv6XfMcrXzq2g8uNYeAy0RwCOMfIk3P4
n5mPcjYRKNdCoOFeV9NRU9mciOmWzBCidHlLxHAPdw8JPvWTuc99ZZ1/95JEAPD+
ilsugW2a81BRM2ncRnPCT7zOwe3rXzgPENR2GkojRgynJ7HMu2RXAUmT/ID9oEol
ATIIlw+Y3CqKFI6Dff+lNJLybo4vlBXwtLcWKlAHqZOTxeOfJh3/6MVRgDyAz+EO
/vFnVl3WoVRKqfgPQQAXl90ZlAUnEhyuKPs8z+BpNjAiw6kCjytTtbyrtEkQ4C3F
N+pe/0ifMUo9AvUx+yry0CyqqGXXRGorhdGsFBRBu8pIOcAp91MjRmkojN+Z2htu
u7WDN3WkCQXDhRGw+yL2B7QyH/noSv004IDKx0tSTCTLovDi52h+Br5nElPxZQyO
xv5Oi30plYwdGCi7L5As5EZnD8+Tvk9xBYWZ1ouv4xSRSZBOfFSrCPlPERBIB3TX
PpvRavhwecAsFsRIcZoo7TK4/ZnJiKpUuqNAiKhjIGhV/hxFvhZpHLRUATSj8J8h
UV30dfFQJ1q75/++wIbzgyTdi6YS85LJHWRUJ9uszJEPP22otSEDl5+JxVsrcDUo
Lzj0jCkWD5YgKXguZWMdr1ZEh59iAII6e6XVNTwTYovr8MG+8gXt6sCaT+MNL+Gz
SgNKx0+bMm32Mc3yoUIrmgMmOqqLkkmkKUdloHx6r6dnPDxuEDf/TarJWhnXhhO1
JfVeJehVs2T7DaDXoUkI0YFNtbl20hnxPjkGW6FZ0tgDZqlzr+0uchzTTIFxsap7
32yvRgaop6r58uPnzC7NkapdR73stz2G8oFXeBTtv9qBjfcXW5uFReAVU3Z0hvlk
eGt9VPiBa4o3AkLHrCZoVSxVHJyuxozHJMSuJLcQmAL6slGe2n3f0XJRn1WOYqEP
ovhJHWuqGG02Lhm4spnT1kEmMn0/sUx5KjOkc0QA9Z+PI+Oa/FOjL+E/+rYRTQpK
qE+T1yP2JAiZKRYqe2EhV9YL458urKwLP2+MnpCbXv7nX5HBbrJCZiG7+bA03tu2
qpwy3rUP1NyHYOcHq1ZDeDOkxHFr9r/CrFQ93TSNqF7pU68l9Le4WI7dTKq0AX/0
JluBsBs/scxQoXIOKSoGm2AIvcX8EJP33munYBRMfeIJt0V9nLgMkaPcD9PzR36I
rXho5Y9dUZVhJOcT54/bi4xKXm4htKP3WLlb0v0OwIgw5N+lgLqpq51sI8Y5v+jx
avKM5doHqbMTloJ6sshlkNdgXKCx4jcYVr9eIjZhZDRcX8JTZCrMwAlk+zvb7dvb
mYjeu9zdLOwAMUfuqS/ir52V9GKkVdWcGnsztm9zgfVzt8W0f4zhcGjUnbh/lhlR
5OHN5YB3Vg85y5pywVwgOr/HEHH+QTRGUWwRCjc3x7qNTeT7SSG70ikEaXudT7OY
9wYgYQ3Byb2nT2DLHqQvqYch7faunIO6I/mz1cD/UAd7jB1+glQcl2FsGj3xX3FV
GtOHPg1W45LnnUCfcWhFv/q+VO0kWvbP7wqd+d4mNdPVMHbnpifJ1lx7f4FSv0/T
2GBRMWaiYdb9wRpN01XWysRfIJXQjbBG6Kaj0oYZyhZOkfLKrk2Ig6K9Kt34gwLD
bYi1a3MLhJl2OlnKj0UlTSA0YoX4sJaH8bumRypvpD2f1C+GBZRFybVVCIdoPGJ8
qHkTIlCgdRjLQWsIM/fnhKXbRKGcpFWwNXA2q4CTf+xOkj7xxLsMHFfJaA58u/ZQ
ovSK4xzpydpZQ3AT3PIP4knwvlvI4bSu0GW/3P9rBy3VX7lwu6ICUFwJyAK3scMT
O4xzL45x5ZyVWksiTkIwaKdEIKqVJlFpl20HFDFMJIzTtA/ZvTfoU0Wz4TTArJmt
OYj6qTxMyXXRn51fH30zZ6b5dfAsymwPKdNCbJx79duSvG+r8M7b669/JXV4/BDn
gtXSbiTLpQegp+Y/xFkUTpyeus0HRo1A3jdKsagJurYRS+qa98umGnC20Duz1/w8
leazBgbvAa88Cjy5kxB6zljMqO307UVgKQlZHWwob4UFR8g0ehzZPybr5FDvPgrB
1v/HNZNrx0HlCeiKp4LKSzJYI5NTqys/PJn4ZKUCWBdvaxqw6yonSwbjZKKEUD3C
YpJwiMycGMfjxYUJcurWTprw8a9YQyQqbPH7fM1pZ0EYFrqim1e6WBbvdGxouSrD
f4EPuSt3HeT5Pe6oYFyiAsERW2DMw2++d/MWaSIoZBluJLQF4gHAVmPaBwAnAyvx
N2IAtrNGcwbc5K+GEda/XvR02b2BDxSt/XpqC1cEseB4YjoEVOw7J04oAhE30Edi
+J94FaIzhl8G+RqxkF9ctOrMlvrkHi/2s9nPZvl2TfzCq5TruaSoPxUc8D1/o5Na
QYhfqMSqg+yQupnyJlHVsGjlCApChkPg+t4MAVXyc8MhvLm07WhEahb1hIOl0+uF
ykmwTknt4STPca67Ii2rwO+yO/f0FMB02R+gynrorZcm7YIrg9g1hS8kmslZL0G4
uNTK9Jq8aEkKs3PUL8dmLLj7lkNgA6AoWOVOjdz3X5gPq1puxmUauc1DRvZYDced
EMBe44KZAmqh9GgGs7j1PArnFRjovBEUDlAqGoJQd1Zr+Ny7OeVs6zIl5GxEn6zo
KBHuNDBy4yQYa+Xkiw/+HoFSDtTaAWz64Vf6nTu/uFeg46fDs/rizK5muPqM5LO3
du+35zC4kn2GPVMW1CJjtokmAWyShByCsNZaeCvfUHx0jGG3WmqDxafIvKYKf52v
04vukJ6IVWGvz6sGSTOaYAahajTyJKAM6hQ1S2OehNIMsUhrwXPOCgKeFj1P4Oc3
jaFjHbzbk8uaTTOrxm7T1XPmem90cmhD1n+6qrCRkrZmqyTwHC6eOY+jZpQ8xitb
tqsKfvU170ReFaBgx5EbuVYn1hZ5XsfXbMKq/JUguZHZ4pUZGwwTTGT3Nx2KvZkN
NwlPZs2aPJOx1hwwfofCnzzBQ6Vv9rw01+Quu/wMr84VdDqFDx8EZhvZlwgb7spm
uR/aLj7W57OqMFadDNXTZyRUxrE0XmCsSV9EY/WXql1Fk279+AowA35lJDE4jinb
15bKJ9OV66qQG+GdlAt/NDBaAdgfmO+Ux5UqU8dfN5H9QC9y3L29iOdtx+2DNtqq
uXx1qk9MIZ69W6F4mN/2UlP/k1LvhVnoYUa8OOktjfiSzLuX9j4K4bebdRxHEacv
kdZ5xfeUt/nQOltDjMyfH8FLMs8mZ1X0K0+xdjXxU8MC2lTMctR1/L5NTS8Zdt9h
+3DsAvX3hDcqdetDSH3zN2mWowWMPqcwcd2oM6lV8ZnyOxPTzKRWqgzUfw09syYY
L66ckcwyWzgf4O2/viBK9wFN/+XCemSwuSc/2auAcLk41DhnfGX9gS95RrkMr9tp
LWfA3w45L8+Qj1mWZcnG0Ebu3q8WmrRX/p/mt99gbWbQfrO5xO8UsFFMxaLEpsZw
UNsJ9su/Hx1EbQuVO0bJxaAb2ZGaDnnWJrO3Dc5QzeHglMzgNQUYvZX7MjGRmR1p
M488PMAqtbVkBVpL/rYmnfa7oKNhf02NOaWsIHEeQth1WtiEKpZ9thDdlRVpZRwc
MIzG5+OwO/1+pbEjo2yPDHVXDiXIX/T+AQjzpXuJUlV9wEzDp8AVmjQMaHfEaR1H
`pragma protect end_protected
