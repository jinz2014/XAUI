// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LsSL0Ztq9d7+15kXrR+T0S8e/zUFDuhRDCAkTrmkQsqGhrrF+UAlWDIIIB1UPeHN
447i1J6gQHd+vSxpCZP+InqVkdSenc0DfWa7QzuAwwkjs9rXooZoisRyfNYrEm/r
kFpuG86rcdavm+45LWJmRBBE/5tmvBmWSeqOMhUyTJo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
uX2XR1abHevz09UTpaZxfzKMq43W6AML713XOq7jKduuZcAFGtmFdnjqOXnPCvjF
0hlkV3cxp3dp1LDULZR+C7e5WFabKYZvxOCyQKP7CKyrtgDXJh7EoEVFK4M1QMeS
8YFjfaC7xGS0fz95mceCBIxpAhw/Ova2jlCmPuLYcP0tEOVtGAw1/nIoqGjSr7eS
KX/DMcXAkOBRQ5s9rwRINpzsaiMp2WUiqCkdKiCipzYPuhcuL0ZGUsAhjnu58Ps8
XfZ42IHur71m6pWG5S0t+Lf3R2fUuJF9KH1lADpLpJsP4saCUrsFt6yQrw1pA+EV
nb5VcWTsTwPUEX4/WEHI9X4xtZAqCWnHHcrT5dTeyuo0Qu/Qof3GjRPxrZ1MyVvV
ruGsOJl8HSAx+COpgZm0YsqUaCggyEQaBVcY1OTOFEzlRJ9kbjh1NThZd0KUFFwz
Uu8OACBMffTETxSolNIQCeHaaHhEPE30ld4nWYmbpuST+v3bqFFNEbGtslYaCdBd
un1cM1pqjZI1THeDEXJO0kQ6t5WrDxMELArtlqB50nPWHy4cxV8xxU76FySUlUH0
o5rdN9pBNhY+e/SL16fD7PHQ4+gbd4DH5bVMcBPdbFD08IfW0LMl3vwHQu/kWZ+f
wxsMo277HfI28UxComiAlLy9JNb2FMjlXrpUhPnVZ0vuxhyfnRv+drGkPxuMsUwS
cKpbwS3s1wZSf3F0HjtBuIrN4ZnfkAaNHjIe8xDYr/0+hg97RXW/4AflxecrdVuI
mJnwgME1cGsEVXeK73QbhCb9EivIX0yX08AyuaAhB+cPqw7KTTEtH4U8wsWgCwWL
xim1nzoJnnuSvFoVE2RLKSYpNyuCur1RRLConkLUBoSJmBNw4KGd1vo4Ph1sgB8+
f/jy65ix4dnyhKYVk/pOVQeA1oFzRNpcRLaVTuoHxF/tgoVFvNUcvouqUODTW5pm
ih+3xD+fJUzlxX8xCkHT1n4lfwQo2ZnH1mN4lGk+TKnOlzZJCEjxiFlAUKYgDn6P
NWWme7nOqhekS7def+em2YobxBXZQmLERhz6xYNF/eioa2RPOqVO1o7FUannH/Nk
wzQA/YzUm4vmTzZ+6NhFnrfPtjk2zO5sJvnv0taPNwECk18yKFOaDWqlRQX+MBFp
w/fPOhAZ6CimGQ5Zj7s6x1iD8oNNN2tB4Pyd+TmiSybyRMoDp0dW8OLS7IgN/yjX
hJ/asIjuZrIPrrrn6ENfF4KsnfNuRlzod2+OAsQaIoaXREjzS0kC/4/1O5YyMtd2
FqRl+yEaL77yuE3apvYTFmjAaj4pBDEAdnwW9tvMe+RTnQh40uffLBCvXTBJJRET
pRLmXoO/jS5QXWzUeZCAB4iNBwc51FDObInbkKN6dc6n1mz9a7MgWmip6Djikarr
AGbGBwsQ8xxFL3zYmA7YRfvx8l1cE6/am8ah72A8ZiuIdqwC4X19B2gUk5lO6B4C
SXd7bYQBcMfJfZevn7lwwcgZd73D/f4MO8c/LXepE8IVvykgEunvoch2dko0ShCN
LlHqnscEjzkQHbOfd4KTthq0R4nUb3hm+XC7f99f2yxPeJv+HqaCsie9tCUunEVW
NdL6flhVqy3iiZlTftgtf/zFoIfU2BfEfVYTpwLW65X6pJAEMjw9Bn+wjqsclPx0
JL58DbXrOrT6EITMO7GcO1IbtqI97xCpssttVmprkVvvKCdgeKWStMgWzl4H7Mhk
xreXWNCRK76IOp/MBbcrIo7GYd2MAu0txBhbieEjR0osvLaFrUe/koOkdAeVSlMl
txkrdZ/e7EMUhB1E/vtCvAfWVR5NG8A1lT6Y4wDYVNr8wp2jP6/8AHA+o9CKw3zx
jLp3WQ46hm42lYCcrdSSa2YbxB+4G/uchz/kQWg5dMFdR+nEEC4J+HSe6noqzaUk
2d5OCOImFErRpP3GO9M/tnuUT9VREovtP7nd1uQlUhuyiSpRoPcNwY2iS5tkwDcD
VMXOYtC4G84spHmKYqTePlcxVdovEMhGpx8pPtBulZwcjetSwcfTuRqdp9UivzOw
yv2jg/A8jrNrXK24aCWjG0If/xoUgf+Yy59A+OQBuE+YJiB4gfivM952gwYx1pke
VUCvAQs72th5bzWmvh+yZstVVj/hTVIfLDuAHOW7ERq21riP/rtVGXmopDw1ONW2
rxqP+9FyDrqzfc/8Miio62S++RGs4vTYBJVufuJnLsNUrzhZe7ex8+RIxseJ8d7O
TdzFcJgq0X+EurwLOHwhItbBN3WX4R3HmHB8TvY6fofZwzNE8CBIjdzxHt9K01uo
RM58tKPmUcPr+epuzor/1NvWoeDIYyBUtO1EsRLotCdEFf10PbX5BV111EfYeB2k
VR8A7YZYvpkDPKRU+f9Ve46y10yKIqxBQYKQZ9FcLbD6qjIw9RxMEjNgXIyH2+/d
XN9P2qPdILq6LzOTYAPFmxlRXjSpI5jM4KwMqKr2d44NnqRFmaJ4YexGgcR4RKLa
LKQJCakt9CrToW+WxvGJFV/u9YYy3yXexkmqEZX5X/voYygjvcNgv2OQ37835qUm
+tTfw6avaynEC68scdO+DpiTBZ5+U+hyPToPtegqd3yG+Zelxwv0mckAelzpkcI6
i79pxEcCgm37pBIgUVMWb6OFE63yd4hbh7NWRWt3W0lMNmObPsH2GkGZ7idUr4V4
cAxBXQkpFd47KT3X7XiNB9MhgCbWsyIEQO6EWaB6RNCesNrqOIryb3DXuKgjBgGv
6YYjNZLjWEK6O1soloAPV9lvpPlEHu9BvmrLrfF59cNX148MfupSM//f6KInTojs
dbB1a8p4dFwi1umAJclut4Gd+a6CES4b/g0zFqSQ515sXj5Bf8qI7tfcqV3ro4T/
a6lXQATO7aemmZc9lb81VoHlEmdQIppWpLsRBJKKtOhGvpYRvy0y/dYMXJoVAJX0
6iyy9gIBcwjDnPCVyqGraZKuRH9aMcN0Myf015swvQ6RCLXNkVfBrx4HeabKehDE
S8IvJxtDgwyRPFXNzO8EweYcMWTKFwwOswZbDJ0r+QrL3chwWinsbiOxhDuOv2/m
HJSGyo2KllF72DxlTj59FiMzp82ot5ttD4leCc1vebcTSIFoqIUwpuqJElouO6cv
LUWFoWwv4abpgXpCzJbONOBcND7sHPDOawQ72r2xT3U/zq6hTdG6r2G3DLPL0Jo9
IY5jmIZkB93OlqdY2uA93513qXbb0QyMP2i/VSxZjO8cakkqqW7o63i/51BjK02R
Go2pyOtxtJ0W0AURLkkAi7hGDj2lYBbkonvqlDrnyYuRejYX9H7gOXvnesw6wrQT
t5M/Q/LLhb2lNcojYqYqihl10jGqJhBDpw/Tqtd0Wklmnzi3yu1Umt0L7gCWIhmE
Dvj6b7HefIhJBWs8oax0UmlZdc+4meEh9Dmpc3tt5/oAUKzUgveaVDpFnZs7RHmA
QOrR18PuTG1lZnZnxuvvAMCmSM3FmPv5tiQykq1F1utk7ScWzphFtnlsXh7bMpCD
zfv8BFpFWago8PRRY8XWqR0TMr0phHlmiR72qy4BekT575EUSBvefvF8nhChLWBz
fai5fF8EyhWWvMoQXv2BYet1sRYJuIMfAi3L+dB8FF3cSdpRdqb+ur4dFCHS7YTy
6g9dkTlt8NdizdebiWFDyCaMAuISCeDcy5nah+KxlclZPsTKN/G8lITFgVFDlldq
TnO5poIe8duK309kK7/p8AO1cvjnME83ESBXDqc/m2DfqAyZLsSzEN9IAsDaodBO
4/J4LTF9IUet1orxNJQXHaEWyiUFAlMRa9jQ9rxlhlis07nc3Y6lz7oZGQbgDH2j
XWApdb6O58PzEmO+cltLKBNeGPb13FJATbaQYG58CmZUVr/dAwG2Hn1CF78g52xo
EuctVegyH12OZKmMK4YpYSZN/FcPNBWpxo0h9jWdwMpzDed/QZZOlo6SM3jqYN0D
aJ4W7PJQ9Hr0EMVsbqMZxG0px/4Hlh5o8vt0tZx503kU0x6Ejqi9mAYAh46Ac5rx
Biap23lzZHjHpZkWxob/hxhM51PFtMbJvVgjNP4tubE/ckrJNGOasyxKICoUNlqP
bPDC/D7vMPK3wreikk94cNVpE6Ia9RVyqXzR+t6Mf5Fr8TTXUYnweBy6es9/t57j
DtLD3nDD4NKRM8w9GdAicEf8teQhIq5Ko2FyzMFd8Z+lkYDt9DXfP+qN0eUoI1mi
bWBMOdlqnaM7cXCV6VKfGEH3chr6ESH6SA6Zm+Ft+PaVVMvCeEuMENedS6rgRWzO
Rvb6T9abJYDzsEAxgtpA0gK+yL55dHxrcJ3byv04LhhLHaA8zMHj+LdgQlLIp+ZJ
LYWmF477/NhJ5ZrxYKTJhcBAdS6t3XmXsPcDHo/dfhMSqakPkADapveqcTqUdkZ1
45N4xHwFidjbEX39q3CAJcRbD849pSlIBDqtOyXSZjJt0Lu6rtLs8Hp+n10tNq/L
fhRybVvd2EeWAvuNwsdSevJt3GU7PlX2oiHxdYVeZETIBIHXO1zCNivDM4EC/UPe
9IVldmw1bDXXuctZTx9IlfroUbqfU69oq6QDbPS61gK2M6mW6tuI8tUWHxJ1VHGw
TDRE754xIAN0mw2y0V8f2BYgUvUMqZTU0l+pbrtoMpSJa9lei82ezw9mers8Etqx
0P60z5RxeOtjrlFgM4wolCcNxMuw/2vqghgZmDcwGvnAgS05C3dtnldVoC+EES0o
tibku0wZrPh3OF4q294z5G4I+w/rOpMi8cYEKyZNN/pztggDvazwG1w/DM0obpRD
FDGPBAffCuw3gwxpEEut/6fyzvpI7iaEllkFdUdxyUR4I2DZauc2roMCysQWpzeU
EXGuwO7CPFFC43Yu6QWsCn8Y0d4gpr3+r+vb8PAwsktwh3bBAxOzluDDWQio3QDF
QKaEh0T8VXTfKZdRmm+Xo7B/10VRoV4H+bDIVnIxhB2UD8Xh7zTJSyiiumPdPvZ5
mPLzYqik8TxqPgeXz52iYGrgZGvpkJXZKXxDuSX73iuP/e0Sr+vbGoXIlhOYTleJ
oXo8nq9BLWEXBHN9/498S0oRXLPc/m52FyP7F63LDp/AkH3DVvhnxBIfkTIvIkfj
QlQi+jLExjXJ7Fr1mMI1KgfUY8j5Y5erKmw4X5zehSg+8ScAc5NyQL5RKa588D67
XW6ZpDO9A+CX0nmVl06zij2tFSku79BrznUlWqi0WHYvzf/o+INwk63F9am3jXws
9I1PHLSbGKYo0AgDGOvaGLNc69+0rDYM5pvNgwHtjh0om46y+YObsVOlabjJVxuy
q5pe8QWVw5bs8m90Gj7Ovd1STT9F6sErOlIeX+/EgvH5SN+BNzQO+XVlwEmKrbTb
E0kEkg+54ivm3rM/gKMYjC4jaJjYHAgJ6fDtBItNYU6f3AYfv9CWS5bV7wXSpYtj
cR0BeDoEegxH02f/aL4TQVoDDHac6Qa8J9IdU3X7b7lRnrJGDnRVqi7W/ASPkBXI
u9PwWcTStr8MGWsoaCdR8gnhqqOH5H0YhTWKFTEqaLa3zM/48yJVnINK2afqPo29
u9nPG/fXf5oet0cLBBLSb78Qe84USnWyREZpfKYWXJTqeNGwmOVv60JMHtq9fqIc
SGrTHh238EUYiiKodIYFRxKgEJSwjHn5hB5lJjk5DRmDkalAgYHtdICrOgq7KMcc
zdIfULogK86+za1qEa3hh1NGlpxlOx7wXbmH6Z/AdlJ75zbfiMncnb+dVJD/MLs9
sLiXh/oxzEfqF02A+70w3JKFuGoIbQQywFMLUWmCb5no5Z0JteQkwvhQOHhnU6eV
+92wEMC3bpY42q76+34TJx+2uI/iVd56rsWKHg4wUoyVzj9wagfEL5lIb3SZjcWD
URfUYKzOavQK7IYQcREobvLUUcxBXHbCh3yKHAsjAC/gwf/8qgs2SXpeJUDNBrdZ
Xjl5E19tyiddcpEUyPhQnzpZscvnRkmrjxaKS6J0bU7vTtdaWQHtDzl8kTPvBvTS
8MGsMf+pEYzqN7H/O3pBr1t8T3Df8IOUA2516QTG9ctMePrDVCEl/6w40RvFuNoS
7ZluzWfySyDZZ3vC9UgV43rQKjB2XEUj8GM7G0XblWaJg/LchAJxI67M5Ko2JmYI
ryy0iLtFp46RlvpxEhnPetfjlGIaKDQmxmJPYdOZWFzS0XBl2jfyaF4boqwAUjGn
TeluRhJWt0aDayg1nxtkbAUfigeYj49mBj9sjC+CXm4SrapIsnMFYu4JzOvxxUCG
QVw+7EOsW3H/RSg/VygjIFWxAGdFbeKCTSVfnZ5ayT5k+R/AwsrvSBahgxTjBsU5
IKZ26tqLcQ2dP4dSDLQshcWyLuBrMIUc8tM3/1e+JmYFrswCFpu7bURmp04kntkp
52yGtb4e6TTEgLOJVJWkzGJx/uv3RlLkXno1j1pLyjq3sXfqz3/FkdyloI+Wqtc7
3+SfCT8Xb+RTkPHeqmtIysG9IaykaCR/ErsUiVc96hbeL4Gnz2XHc2ZFw5Z4O22L
XwugzifO4t/MAvSwSOotcUGdz4DN0s5ev1rvm+HI28HL1rYgzSTVgP0QA5yvrLVC
9AaWw2v4+xbdRHpqMRIdasKIrE8VcHCPUapy6CtMuKFaXqIsJnZq/8PTy/TFUIkt
hpDCIrlPzAUrI1ZSTCgf7tV0Vv2mrjh+LJrzxRvZT/UA4DUIjoQdyz/T/yBDfaUZ
nonzw2nk8EfFKz5e/Iqmeiv0qKhEjBGKfrylPDqUHtNo6PUVQVVynnlkzbcL4rHK
Zf1v9BVt2Aqwhtz+qm26IRXs5sIWwSoyRrL0oGw33F1lL8Vo1YZf93hFxraroBwH
j1Lx8z1b1BwButlsCk+VCbXKVlmpopGQ/CZWGet62TZRNAHZ/qulowYaaIKKfsEh
Mviv2c8ZqWHDU9D5CbWI6B9cmpc8/mio5CfnMbt6jwVdAQvFurc264ws0rQXHe5X
Lw/3kAAxTrN9tXsJsEyOLtxOfJMha3sMKj4xO5mWROMguxg/qz09SVVk0t7EHv9l
QbBVRI7iGW6ijQ+3sK5GrXrVs4KqEPwAUz/mOf8S5qZYo2NAqQodN06ZnJGCpS0X
MUW/M/L0v7TBQJlbqzO6TEnjr1Yf5N8ozr0fUgT6Y1iCD+aTgcH4bApuAQz1PsEr
xnw8k1hvbQqofsHoYQxRAERGLU1tIKchFNN920LjIlDUOYSi7iUKb0F7dKefWkd3
K6RCo6DydHskWJLxIG7+2oENrz/Vh+ltWCH3UZEBLDMLJ4j2hnDcaIjJV1ZHJLal
8JtL2J1iEtgZx/Nw0GuOPyRAW5QHxZtehHlrqEKHqX52Yt36yvc8GR+9F156tUeg
vvNtHA27+AkV7UVTC8aDca/j2JAlt5Ccmlwkcs/tQpvrunOFFdwO/Tw0SPrDhAqH
D9WUfHBLm6UTaxjfHJksLMTDwCfyIdrmsjmhxuazLk8=
`pragma protect end_protected
