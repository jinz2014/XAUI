// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c4ttvVa5xR9SPA0t8gnw5tRjriE9INieadpuSNRyM3jU3KK9/n8q+FUrVdWgeLVJ
IkBkcwW5fNx6caI7Z75VjKYG65HI4d2DaLFADGtHJtUaHAy0zQAVSg7Am7/H9Ved
e2lmlAu02YobuQQliE9X/Ymr49NwolqI+u83BDjA0Po=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2432)
ek60Gcyz2JXPUsqozQDeqlkCYJiFREvd4q/m31Ds9up95jljDiJh6Kd16F4ZT9zt
vcGEQewyAHXl00EUHBtf6HB2T0q1bI8oWdWfvlMbHc2Eqp++U+eUs5/3Ejk6O+Ow
c4CgtdbgUC6uEBjE4xEKcFoVxeudjLHVwAmeuIQQopk/fZIWmt3QJjHupTZVvNZh
KiCf6Xn7b+xw5JZ5/APOvYRTbAq2MfEOsr4eiNfPO2CnpSMUZcoL1v0HZyZdMp2O
XnTNWoWoi57GJE3Ij41qQ9tPJyHUuWhozloVKrl572SWM9wvOMA048Qi6NF9T4W5
/CLqeiXywKs5uZgRQeDvfWeq4dPifYfFT0NiXKkK5bk3p4bDVYAFx1VfFQbgyaYJ
HXLjI1QRWgPmJW+hDz1M+fpdfJ4xXeDpbTbVTtUazLij1HRtufLZxknICaf6w7lL
CFS2Ubgm0KSGTgIkb6lNLw6WzZhYCin7W3l83zf73Z6J5dB7iP0SFIOg9gptRh9x
OCRylFG+MPqz4AFg3Fo4PxC159iOi4nbPN4NB12IZiIhpV+2EA2JEv2QOmbDC8fj
kxQhTgdDvApFmzqCbVoBCKIyO1CU55FdEeoqBx8RilTAamh6m1w6GeGosFLNr6/3
SkbfHEcrXix7VnwPQ69JsFZuxoQ5aGnJ0wCoVDnMxahznKMmI/KyOeVu6Lf6dB4R
0sc+DasT/gTsUFh3AyfGqjxtaNTv6XOYY9nwDDx8ByP8A0C6HpoqpKpDv1NYPQnk
ayxAkJ06xpbg50kvOkHDJBFF0fI7lf+vbSF6cFHFfhyvPuMZAsq6duvhEXo1DPPG
elJkG++wSPMPhWSiN3Zyuc5J1RhULpmSROeepes2SlICLOugHnFzH9426IkKTkrI
VGcmyT9AtngNb4s+WteRRyfj/ssrXzZAIgIf1JhH+Gn/Vrgr42qiX6CgYtdUiuhe
N83/Zyf200s0ISdwbJ5o9oLLxwz44FdGeitd2vYW7pY+mE1co2ivyGzji6JT2OqA
a52DlKSUpF3G+TCkjpuW3ZAZTNqM/o5NH9L1PZbiDEsr/GcnGBJzTfbcHfy3xDhe
odte++u3iAI9zjv23d+VGgRdhU/YVE4anY3cIwsAS/2yE/3K19DEFjskT+8yL5uJ
NZE+veffm1dTDi76Ca/c0rDINcsc1pLD2pgnuvBhRllNQ1hR0COpGj7t8yZmuzRE
ZL+hYx2Qfc/Gjg4vTdVy+KRDz/px9q/itQXGKafcu9e6eubXUPkW7cVKxdgBYTEk
ejFSnMHnVfJz39i1GeJTgjcn+msut9CT3QrN3JWZiwUPVTusQB4nja/7bt+cQlKP
52uT5Pi6LwxfW7htPG90ZTtYM2/WbywvH3aIMkgLwsuQRWGXEQwx3B1v8O+YGx81
6ovE5nZHrCZXbw8oRADDTWaVd/euIta8mVzuwcm7oPiz6ld3+AT5P5rbCOPjXlex
6mrg5P5gWIjaBBgN4BdrejOzaAIYwG2n5Qe6rQuRppCKl1MAE9FAwoDP1KSwWOCB
cwi1Ry9lDoH80InXOOP6IiZ0colj47ThYxVXBAu7KXK2tvmpMltDya8pZTaUA0DX
PRXkeVqEGnQLh22dXs0ouBc1ykY9Te0ej6Jl61WGzGo1dhdMuzUgEjSwffKeIGhw
uPxVEUB4K2EUXQa5VsFxqL909Viap8E96FSXnC4h3FDdEZpb84C0sgjGfCPM+Skk
mpPZNr9dMezEXvdEbHzXYZTFSE/Xo7gISMu1l7545ALYnOcwpoLO6yUeHPgez9Sk
bHKUoNKVX1NVhBfWPBuVnQ2QTDoSmpzUL+b7ZlPBLdq3H1hAZgZjeYfXhE9IvtP+
DQrqzNb8cX9yzfw9GZb56TeEm/jGmRYIlfK+/Y7CDmd/ep4LbJ8HJg70NXW9yCLA
PpG9TS9hZh57iDG1cHtVu7BN5DKJAFmIQtSCZGbb7A7Ltxl8LKbB9Oh7jR3wZLFt
dJ7ZHqfx4SRHpj1Bkv3UdtsdUBwB5UN/Wv8S4NWkT2mmEQu+GXJeGxfPlq5sT0hV
lWbd9AkGWMiQBK+V4/dAeAqnGntNOEJxm5rCS6c35hW/eNqqCzJTx8sAvkKKQbUh
frsbmSUI4zpJ1dgnTTZBaiU7GSalReikGHBY0gialLsmp+Zb95a+zItQbolK9uT2
x8VaY3GPLESiyNB7ARoBKX+lyneWGBXN761GetCumcPvBPsl/fsXqAx5aWsQYEJO
54SAtobxm+7+isOtqxDOZCmeWiP4TfUTnVW92QUBLUDRJIMPjC9XhLkdCUmYr4d1
kbjGhpf56resaumyKsQkg3bIh945XbMEqaasz9ga2mlFwYEHEvPRRbrBKJGKOTVZ
r/obRdG0n5mmiLCblijATxyVRLM5LdrgfZVi41CcRjGLUwca4qGYxl+2DFET5crf
cFDPavpNPN5Q9wk5pE0XzLry3G3cJYqjmba2tHy0NeufFs/7PxbIKOvx6M8yjVTA
UO/Lo3Qs/9rfbiNCdHRWMun4nwxcNXyUnwboqwQuElJVUhNm1doC0kHUP3HpbLFF
ML0ALZm2Prwt9N8aR/YZKKbAy+tVevwSsoZyB+9z7fkNvVkY6w7sY+ARoSK24baq
M24IRYj4EosBYZUdx10UJWh3I+tHZWsL8e6JUf5HYR8Gnfw31uOTOCeQpPUb6M2/
HMQZOvDIJxGL6DKwcDKgwAEaSQwWq2DUn18cdRXhssG8roMe8xI7PHHNodsNosKD
+SloPNtMFO6juutqa1jemQAd1xDfnYv4q7AIco3Mi7I0UtWNWs0fIl9nFq1OD6HS
wAGt76hYA4Oc6z1Vv+/gFVpnwugvY/CylVbNpeq3zQ79VZZpcD/dwzV3FTst5yYb
HzgWMZ04HND3LM5KG+xDNAUn/KA0EJ4Ue6zZUBfOlo+/4RIEE4Nw5dM6p3YjuNRH
nSidfQebTJV5z23bIrmHBuX6X1F80NSD5IYCJRKNVNiKfBS7wz0efElFHXWyB0xv
6EJhHP0R9HoqIhS0QTvrSmGecJSH7YjcLw6U0Hz2/4lB2Q6CoMhGe9zgTGccpQ2J
+4r5OhDMZY5IftjeeSZa8q1uSZeuO9OJlR8Z7qwN38XVf9aaE0PuRjwurcB/b7R6
dNWV/lv2lljJyhvwJ4/hZmywTbDqwcweTktcEXRnwzQpcFHqbBVvhaP5SpCN6UW6
tIqaXLAfdn0y81LAF/AKZLXMNsWnvOZuTNKsmANfGHk=
`pragma protect end_protected
