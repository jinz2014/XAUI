// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L6ht0mNHsVpbrq3ynjHqrUn4vPn5CJQyBqyuE7FIZv+X9OYxHw1KloSUDzlcVsnq
0IfMgiSvEvGIWgpcPReCqwToe6mYcsYEo97pM8+QzEq8KEJxbMyGvqI53iw7Mumd
XBxJhf3+37MM/opVNJTCJDcNxtnAWF4iFHfJWJRaQM0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30048)
ORe1GkWevd1KNrQjglU5euca6udrMHSSB8DjUtgi6xKIviOBC9WZEuRe4sdQbLQp
ReoypDse+z4T4dimSuJS3Szhz0MSwc082w1mqoEBmU2xD8AHH8BfDbxWU+D4U25f
yD+nqtgLSgENDauo1uMVZGrql3k2pi7agDpSXd7yenVjZHFPbIY+JL8ghi2oakFV
aGALa038ki0DhunDLrhHeEsSsxK1kJqSMGiVuZwBqd+hiCHRNLTgvtOrz4ISQxWB
A9aqOklesR7ZYV89sKuvnrKXB32lmatp3HrqbfrgyN+tBBxwsUa6TGiU5zj0YfkE
PxRKiUOlVqQ4aA7Ffit6IaRaQ6gZ4rkSnf6BI9a2uMx+QIyrL9/y87aAhpD7JtpY
mysc2A7hkfBOuio9iVu7zYyGMIb5Bgf0Xgwl1UPGnSQves/JQZbYmn5Ne/k8Ng/T
s1wnrBz4xDRCIYEACkbkkDP2U8//iBv0aBiBSKXi+Bb3dNyWyNtiwLVmqRPX8fqv
b3xUJoYPDtcD5VTcX2ZGMjLkWiZjk7zLytRnBjqLWnVFE2fnPZrRsqSFoPkcPFZj
hyGZ6YGYhnGjcwoAnpM8mwMWbVkVEBuNdNCuq2bp6hjkrnzSX7hkspyWgP+K1FUh
RldpLON2xeo35XGl12mziZ3awY7OpzweNZ6z3PcmzkWN7mX/tOJqodOSHSDRsZT5
x056c+Lhsr3HBiYjZ9ffAdV1LHZeHRQSmGqYEnUPO368vdSIgXCNSh+Ll+TwU0+P
luftJgylbt+QJn6MtLfYkJQ9yxo4PjivvceFg+BtrZFslS4gQwkF9UHVw3tMJp0e
mpL0GhzALzPi0ZptzQL1+OocQ1WaJoY5ok/lbuSsV4kkcq16PRbHcjGMkcbr2E3n
DWrA66uAUCH6uoXo6mCUEjDzYUb1b/1Ez67viWNS5aozKNxd1eZ6GiV4sIyYOdNV
EllSX14Zisbjv6s7cFEDMBM0eyce1ApXp4/xyutBQoZszuF3FzvCCygomrUTlcoP
4ROtlv5nN5/ves0tNDhG90PBzKSra7V5qAEpL3qWUKH694xe2iGapLJIgrHdWJwA
OEn4fl5OUO4ex3GMf6BzxG5no/M1/yfCSWQFVJkR1LVRBzAgJDcNqJz8PoLouPuU
A2H+CPQ4t9VTcmNhZ90ia5xHwWidKZ+jFDSG2tjDDBlISu+c8KSDlG68dNeyV7xD
7oy+8aHIU3eDTJMytjxCEzQhbHud50vra8fplRqNu2f2jhS1s/7c1jGU2DmFo27h
j2Nq6pOoPyUMzOzDhAZmgXcke0DQi/4b3In2Bbz8TXVciaf+DIAd4R4nrORHSnz+
lSZZFj4EAGAHV2PueDdh0+ltZW54WyBN4lLs7DCHYjlc8Vt8zfgrxuv6ZVDXA9Xq
OUUBbVpPBCW46Z8OUXuzNuFDsjD1S4sdsDRzSN3Bthqh0cvAQHcajFWxBFx8R9JW
VtJFNzjzzgpFsbpJrxO+tWlp3K1m7D2Fxgoiiw/vHlWldcXxHldB8kYx+/lb46KV
RLLVR9KYe63A8vT1qP1KqvhxHvId5sQl3Dleuya4ee2NUTrqnoESshmPjugH/9vh
v64TDCFzEpe2oOrampkoqE6j2TkZ/UJTCQvFVT0mhJntzMs+T/xYyvzv2uJq+zV9
v8crSoCtkZ3bttvC8xZkJgKNVQjayLL8OBU8TQreH0a3Tj9Cbbr/ldg1pD2UlCb4
ar8ldmfE3AL8gawPsdsrIA8xXbzFkvj3+QeLU/jTM15lsUgB5UFAPpHcARDYML0c
XWGxfjSMRn5B1xYqs0ATu0a9Q70pSMSnceufLbOQZ8/ppVdSm1NX96wtvMAuqnLb
rzDP40ieYNsXOrTjW+5u3P0iP5QAuqNZYtaVm2XxhCNe0Z+TckK9UCxZji0MUO6j
GAMkbKTMEb8Wl3SJvqmsu0uZ+6ICOL/08fphhRCmen2FmCaKailmGP6ed7k/IHBq
TNRJMqWnNuMTPZG4+tZCl9hdrd0teE4rOEXES+dr3IdOJmNT/24CfLxHXFxeNH4Q
MVk7Sd/i19VzfGyGIzcxxCnLsZDpWu4x8QRW+UUGJv2ffVe1Z4iFAcHhtzMiIvdT
PZxICL0KBeUKlhqplb2Mr8gQKDG5A2TyFVzVHElvqSg9Kkp8zeXz7Hn3MKr8U8Qy
f0LIZgo9eDZOvGBOT1LoZEn6m9T9lIOWNfp51yom1Ha9MDheRl9HMYmsrmnikunH
vKtsNH8Ehwg2yIQhCQYcCGZOIoR4zpLRKj6yFFYJ9GYHYgDcAJuyyWiukA88PHgH
Vu+ZxOPZtZAJ2UZbjhze13yzKxWrkkzWqJ4m5a2KEL3+giSls5Cf1yeDK0c08xgK
uoF5WDz6/f8VxIEdDw0WqNqQdjxzT59H8XB0pnlnMe/hASm1QsxQNE3wRmwrOZ/4
3VqLPnlPIu/1J8fbwj703i8LdV1EKCdS8Bvdz5sOkswMlc2svI9JK8Fv6ZJjF/vT
wETWFJX6Tdzqcl00ZLSi7tylourxLLBm+68DIDHpeR1AXDmURFWusvT30amuo5yI
xuKpBgPyLPJsloppCqPIo9QvrYzSNQ4jF2d0zDstkqV8x5C3zZWH5zYs/N5XFaVa
LpZOrQCoZEyrmLtt5WTt8wTRYk4OBNBfmpAs3YCn0pRAbZk56U1RiiHgJc2CxSEu
S2GMn4q7EOKEln54KSbmbYQ+dyBzRPRqpb6qtbN6QF93Hn/TIKEgUsX6PM0p/D4N
1VsBdxMIqVcp0ALRnjEfgyZXCz8MOEEfBwyTVnB7Ej+HUteh16d5KsIKqdbHbh9b
bxawNN/a4AWQBc+M8fHjr1hwa/yc6ukCACG9Y0OXngWpp7gvLDG/qLKb5jEjhNZ2
xn7LJjDGvyN6sGVImlbAQzIbTu3iGNvW89SbW9d2XAyy2RHHLSXIcgDG+OJYRP89
9UZ4Uj90d/GOv4VUQkuF3vr3xS71QVSSomQbkIdlo+CQ624rQF1xqniShTK56EQI
r137lmeDCeNFQz8uoh28uuBM6R7+8hAzSRcOaBjSXs4wVstmKMzckMI6Kb/THzqW
Ory7kw68yN+2ZDPIhXAHXWmtAAHwBYVyi6gf9Gv7h74wPFupMkOGBgRCkCwKcWvQ
wmHHcxUpsIA5RZaZwRTitw2YodIgx0FHfnlgVDk/ZPVDoCb9zJb6cHxRG5pvaToH
oZ6Cug8SFDM1aXyylV07TESczz+mXI9ltCMWvnpliQXdjdalUXMpGOXkH2IFuXVH
12KlCV9B0jhaAli5wnCSYsiS1QelfogipF9Kcpa27+bnyr961XFKBieiCjvYGJzJ
JptgM8N69ytwkJ7/Lcww7OWfYe/NmT5O1kVDQ8lkyc/torOIrXjzaw4z19OFjYv+
hFOzABMMTu95OSzrUa5U4QlV/oK/qDDN/lza14Z6UYM7Z3d3gsOr9lA3QKI0mQpE
mwl1qIekYyEbtQggcFqp2UFN3YQc3XmOE77/Id0hZcQ6glr89DaLGDUG4CuHANlz
g+Yld+CgONMgftTlZ0vx4NWf1/jk8wbC7jDJa/xNfzN/cz3Lel1a8kAsSd8Ei5gv
Q1w5Fyo6lT+AaQpumTH9X9OgNFkJXYKmk0UJWWPXbifis843lcor/WkLIfN4CNUV
/5VcqLWhtY8kVjVBC3dUO+8sFfd0Cfou+TRMwljUamiKaFBJggk5OBmZwbaaTeIF
WextaBkzPFY1f3jWf5lKGwNFiUgJIgG7NGJcExUQoP2zY5VTe0VOuZTfsdfMn0HY
N5lRw/TysZ+KRPXDZKOcnjSCc/NpHeyvu2uHwxdwNzkgAQwPFBXiMgb/vsvPwCEO
WZskVEODdI8MrAY5O3aUzmqwdfVIGiZzG9kqKO7QeR+735gcGV2Exe2dHktmZXJ6
YUS+x9GKq6dHM0FTSruszBNYdHqcUMA5ZY8rUSrLcdQbdWtlprI+sY6gJheTiAQB
uO47d5jhjNT82WeKYFcPlgqFpReKWn+02986nLODhNp5mV5ZZQcOmPEN/TIcicpg
3FMqHfobh8cPwFP8Jine5UoknNpyc1y63L9zDKlkMB9KMI9Q9L4JIs1igOQKlN42
m6l2daLdxyvmS5mU9t1KsyDe3dSb3TErJkq50kSFiOrUjMXvMhJ8PPsDioxcEEUf
fTNzIoOOmWbr3ZYH8wRW61iKCLcsG6GeZHqzr8Glq7ezcKjrXohe/IoakyyifiXd
RNX1DO3cBXRvxWMgEelQGKdXGKtLm1g6REa4R8XLyyuNZmNVOjV4u5TEPd6mNPIv
t9iwMMp/1ibWhEe05+KtYOM9ajmbw1a8BzooFkOKKhwNnTXLfFGFfKUoLBDOQk3i
TeFiq6J26fbYlGduLUpjEeIkasIBRVbEusQLu2/zkXRmaNf9/V+pOnElarkhhqbF
oZ06+V/7B27yp1lMaCLYpgalFmBmyGNowI7eIGuTNabqesQcbAPD6JcMZy67hKdN
EEa/tEZtIhcvELIGYAzOuU0xoXGd/C/WsuunIaLeXZS4ybEJlPlwlBuLlPbI3bvd
/qqmkYcZb0+xXx2lxuKyC1YGwlCHkSaK+D1sQeo/gySvBWEdfzolvezltUyFTl81
lzNcjNE5BRbyfYHebl99iLt84xOHVEcaOVGcnxxS7IlRu+ikXIALWs2FsnNtKmZj
2O23tWlq1m/x7RX6skHUN2xgexKEEFswfOEqL91rCD0I7kmfcU6uyBcc5d2Teq6k
GVcK9fpwp2kAHAwmXw+/9kaKSVCzQTjJPQmDlXpBfkHCLyjKfj6Ra94Ss9f6QQcL
bpWCeHYzATcHwbi0IS0IrkMGnflmcrZsJtVXOOjvD9Ae6DskVmLonRPfmqjoXzzR
rQw6hHQLPMtkKfnkuj6KMRZwyU++wWzoPoBytCIkOvxwBs7fdVoDrAz7Fqkf0UNJ
ZMLM7F2ZeHEImTRvrxulbTAQMXsOSZaC9Wcuuay9HyQ5UrwEEvZJKPK+mjBuRxJx
q9sJUQIT6KM/1wdb9iv/6vPPpkrMeqiin7jeTCUi7oOfKfhSAh4f4572ovmIb9bf
w1IsLoFSW/9+ZI/rPZU1WWYYQa98v59sMuGGHs30vQfuH3AMOmjZgfcGzmnUWSXn
Axs/onOyZsktFcK5seKmA/hNylpw/L4daW4MIdgnD9SsVj07uQ9uwr08r62E13tI
URA3LTwxbQJW8szD1fOrpwSW00uxypGIr6Sy7N9OhJzU5HabBV34Rvd76P7mQFx4
J3eHWRgYArzTQMJCCwG9qAdgmDmx1Vl9Vzq7uUKLu0zhMpaJDIfO+/WrAXJN7YJ5
Bpi4bYo0wCp1C0nqLAQMRzlVH4l9qXCjaWEkYky9GxlnSn5Of8/yoYXbXYXuxo/x
GV/4MEMXTSHwADkN6tVhL1EUggXvm3Vr5KF2aytQ74c7TXMYWpCNehLeKVA+vl+9
2ZiCWHdBVkDyVF3KgGFRwHMtypBA3TsIRv4Rbr66FA9QSSFW9mFGN641aiPuB8yG
XPGYnAR8J5S1EW1P1wtEeK9lN/Tu8T8dH9vWwmSPdWp4CWLyR7INbepjzl1CtCPZ
n0xuCD+vD8hlDaoMv+ROqUk4SOMibgBcZbxT9CR09lnT3CVA9jdya+xKkIIopGE6
wDWNsqAKBp+T9Zg0FwyIPxrP9NU1Ub/kCjI4r53jTSj1y7jBfCZ2eqR4oyJ9dxmY
4yM+3txMaWiZl1YCXH1xRtAcXpplAIBbiUQNSAczzp3ogP/I+8B+GlEF4xCVYM4a
xPd4ecmAebQYS4RXNWgQ+Fn1rhaqCiNy10+LpgUQdHL0qbsTbDy1xa03o6nj0tAC
Naf3hrXfjJJxSEs17SvyqvtmgCMcHqA1rWwrL5WHF/1yvLvOgbKI258mbSbMmxe9
iFAwSx/pJMHyRMTzK0qJK0aZjVCqAs0hnGcznA7jEd/SVBAJVwQkZxaiZU313Kp9
WHwtjk61QfbkCATBMS2xphziUkf85CsvkmdW2bQ9xdut+Z/lfrptm4X+dGfCRTvC
h0CR9qjuKx1vxX9kCn9HEB5ltGQ4lbHhXzMqV50tInCsGQj0iUL8ElbBZDCW9psZ
T9QZ5SC+bm2dwomXT31mwBO8p4aWsCwU9w9Nn7WaAHJsidCHGZoRWQrFzooCcSyl
E1KwY8MtN4irfihAn+3wwFjCwSGZbTjKnXQVD054ZGaWNylAm+F/+HKxmGR6fLmY
/ERT6wmyf66kbIGOGrMM27ssrYb9ygCMmncT8df+LJq+DO7fn+R1XtIm58RSVALD
+v9KrpIB3DjpvVisvXlIvw+D+D25s7D3phNe9S+AcQv4htVUqP+Qt5233SpDg9r8
QhQAEv+xt3GLj1vFv2/EN9s95H1f8xf1zgVw3n7gMemlS2jac6MTZvbBlK02vnTB
qeREn65tcABxzkkjupoRJHLJ4Mijj99g2BfL/A1LAB9h3UUK1W5/i904ZYbvv00f
cVWjz5QspzjQtmSdrB9NWjhUKMm+ngFkrbKuDPflFDjQ8o/skbQ73YW+Wj8dxjC1
mo0Djh0Kd+cMB9XA0C5VyAkD1JW/fza1XVajEF/xHksdSd7jfpHsfsPZS/fxIRdw
RcLPvLWnlNWXYe4cYDQyPcuTaduOWkvG0NxYZ1rUvr4tLgs4ib14FdRt/IW42knZ
9ZVD5kKyQs7PXoJbS5JJCpI+i+EU19yBbNApl+VfIt3nMemSJPZrpCzxJlpVQ3ji
lSwMYhvsL+Ji64Bg5WpNggFjC4jxnlvEHHa4+U79garWuTTd8cAFppSaZrphXP00
Hl3I642ML95A+R9nzLlxzlQyhj+qyN+5j3653OPUPY7z/nL8MU4n6oE6ALZs+fFJ
6yFNsQAQDH8FGv9TYe7yKKB1wVM45kCDW0P+nzvU3+XZQrQ7poT1HeWwfUT7uo54
6lE5COoZpTfR2qZHafLW4xOmrlOAW4br5xJaSavl+7yMGIbv3DNmlTE6DhjeTQBM
GVZ4meKoNc03cMXSYTaOrqPZRZb2YJJFhEk96VuNjTea+POSRNPbJDDY8Vcu5VHZ
pt1SnWdhAkyLav6fldt9u1JGR5A4ED5f9JWdUSWnYFkgL7X0ysWCnluWFVOkY0ss
QRDRSqaSp8CeD+DrIT6rMTVH6atZ5P3rX3b5W/Io00rTmCO73LMWiedFXZGFTX5K
JdEzhB3EpIa2v1CF2JNcL2HLC4LIPxdVAnQcYmWHqdGwK5tQrAB7ZWtT0fsdogxR
VY4FkZ53w6jiEB4XIcqN3b+BRt8i1H61ArhjdYWQgpHJ1bwLzS7shFs4ntix+F3r
oH+MoaY/cHW8gN5fmAznNxNP4m/yFlp9A2/yV/Zh6i6dwzftacPJnB0oLXlXfNEa
vb8UEtKXfkjMyclprinSzon1M/CUopzD5+gGedCEWSVFa9xwMLXlFIRKZRi+351z
G98rXQglb60CDQ2YFmBFXH3G00dBWvlS/fHYh8jTxHnNpKwo7RVcBhACm9ogfG6A
golTajS+DYqvG62xdfZaq4hZUNdZtdwMNX0eBN5ZX1cyElX5OElH7Ge29TCCvDb7
W8TWbp5np0w8VdNmLF8XAY5winBpZ/irrDy2pVW9Sbe2Bt8x+Anr6MXxYxu/mEiD
e3+vLpRWmXE8JRDhsIS5V8LWA1UzAAdzw5SYw1GnpsjVHXhKKrJPRwqgwEcCuTna
QdrVulfvw0oIod7TZC+rZ1ELaTXy7umPVIq2Qu35FC0iHpA9hmRvYCrLe5HOYdaD
w5blhVpO0tEKvBUEeD+fVIgtXXDvTj/HS7WDYs+0jfv+DGssEGaIrE6u4Ccih0mZ
XDWaYvXmNR5AA5q8IIZN/nyYcNzPZjXaLvAPEi03MmJc8dA3scbHoyOSwlkSXfKa
Mu6fEevqdU/11SfalHp/YAmHxdDJnteCGxwCZ+s5X7w54Fx18aqNDwM9Amz2J8/m
GntH0F9Nxz0iyJr4eFTjcv+77Xb6FTOXg23xBaFQlsWnPrU2idZx/o3GvrjpxZtn
kLmnZKW+nRltv5kcPOGxVRjizKe3CyIXk0rY1dQjUNLtC9zOF9gDsa1rdvmNXduq
r3bfk9Y+P7FFL8gM6avsVrbnHXT9obo8vrcK8vpoIaKhfIw0rYSzqa2K2P6p9s/l
hzwjpMX8sxanHzmcX/ozBZF/+2pcQBn5cV4+apkKY7tGwHbzrYVEPughohX1g2FN
Blov7+XsjjbroI/lyhqE4ZzInR+P11RpoykyTT2lL47w4pi7gV65X+g897qt5tCY
Y/NY0IdjaKd/5h/xfTc0qQdY9V4vmWxo2HUuijNOQUxYIDK3lpOLfnhXRdqsofTx
vuErDQSiSRXMp7G+XJX1gS3GB971gz7ikZgHZRZa4MnODicJq814Zj3bmx8EkEFj
guPnyYjfS3ApHXDSt1BA201qnlpB6xO+tWXUl7MsBIKmD29PSe1qUfdg3v7ywLNn
ICoME8ymKyesHWOOoDDOLSVtRKU9QUKhpOvujQM5t6FxXpUk5fsN73FoX0xXvx9Q
Lz6xN8XSw8vkpuTb/6J586GcHxsYrs5icfGBkKu9gTA9LO+d3kpPH5D8dSNqHJiz
r0t/AenpTo/MQEjPhA6SlAamLBQww6KvvrygiEOZsJyoM9Iy6/pej68FN98VdQZR
i1jRsyhPWvBKae3q6cg8wElqpZm6/MBB+8dAxOcVRn8SusedMB4Et5MzXF5vt9xx
C8/1AsVrbOhOsirS3jwcnNAsB4UAquNiIMrlEXVRFx73uW77FPN3zxSP5zW2HJTw
e4dej30m7RK9VjoTAxM6fNWF6HsKRZCBzryKmLgZBDUSrriviFJ/0kvj1uxJ8Eeo
cP/SJhCdYJsVMutS1+jDn6DHx/wYoJZu1hMuJUIm0mcxj9IeEKTg9J1mybjMVNPq
gbPG4kGbK5y8yqZ0KlHOnspjkqiJhJwVXVoIXcxTn3suR9rKCXQQzK8L8ODrtIxa
Jd/Hb3fD2lALUfGe7enVvaoJjDr7NQOQBNSP3A1W0wBWPPZy2Isz7wJVW5RqZLKR
4Brjub9CR0v9ion0y1dY46qchTOTdGmeaho+OnT1x3F1F7EqT58cou9Jdc1pMNPS
q9zEXRFooO5tO+4v7HPfluKX/veejSx9MqR+uaGfWhSbJbojGyQpiL7XscOrjzoV
ZlQbbZXdE6nRfQIHDIVIUdf8XbkI0dFQdQNTYYkCxO9eV8erbZUFEdJK3geRiUix
X5EQ0WFJKOYPYkyLqDiep2oKbLRW/hFD0jXUwlZCV93VleBkB6vZiqtJ77cpFyC5
DL0Bc4t46m5Lo1cVoZIDf8AH1JnfpO/Rk30aemmTxm0NKc2bYHduBXGQQWrp4FEt
bQnZ54lqCCCIMDnSTCVMt+Ht2OIqAM8EH1hsP1qT2GqQR1JtLkbr+51U1FUYCmU6
CihiXXwZ2UNSGgHF4ImDnzsOzmLkBf/GL7IfjhPtHBu8jppLZVcU1xEil8Rbs2/h
xVhwcQJB9sUcoIQNJXIugWYOGnAN9Sf+3Agkhfr/xG4gIpTy4/GWAfh0GcjhEvdp
k2Z/gP9jOMuuP2FXTc3fQwNmAsi18AHgRIM8nnaeZKsalVxOEi53ZtgCdvKaxwzw
AB/WGC++RCM6aReQIwz7tBgo40lWsCMM0IH6yzI0611fRmf0REGe1jx/j7CiHAl4
Lxd0lzH1R8YK0tOXo4PRp4Mb0Rxo5PDY6qGbFtJIy+rK/1YIQaXNb2Fp/YV9Gnuv
oA0qW1e1NVB4vRQPkOgrIV9usMZgvoldoLaXpeaddfVrxQoW+purrHaW1nRyj8d9
Pvu73/YMwTlApYfYnXyV+x5QcSzZ6PknnhiIfYGeoEU+K75Ivwu9PFkK5ztjKvrK
bjuLvf+q7ylqkYh84yHXdfeVofDvskVBww+1h0NBW3M4Ey2w1BK5F59I1SH006E2
BA2qogzQUVeNIlCG5fmP9zh1Jz+R27z9RGg79tohD9G25ObIu8o6iOGVZLsr2yoo
Hl3yr10Dzw3xP+lagCNFabaeLS3lgKVMaYHh+3hcJdNHSb92NcoKVNNDZgvFEH4/
CctqaGTyTjtIgSwFzOHLrTZDI/D/nzJ52N1hs4uWV8M8QrY6jdr92BKKzU0c7Gyy
Fve29UN2WcFrwK5iP2k0aYHeqfPYUzvv/mm0FLHCCYEEmskhl8CVVOaHlIA/HP8+
owbOQno/rnk1OcEQ8qGbE2ccmlNt6BslUEdpH7XwpF3iLVFjPHyK4UGmaGiyvBu6
KGnjrhXSF2//fW6JDSAfCVRGFy9ey19V9CCFTcRCdMwzbG4rAV+dY7xxd7fjcF0y
norwb/ikGDdc4Ao4J6Gh90HS8vNvOvKRW+IecypjRm4RNQFZLGA85nfdkEme8BT5
2MTsZkZ/iSNdFW2OeeqtKtTH7cCMvqselyidFS9TCqSbtQ7klVXqkKAdIbAWq+E8
Odn9zd5UtxkAQQoj2LPWAVanFzf3FyhWp06qX9Q7txyZglwtLHYnv4TIEtyVsGIf
C1pBNNC6lb3auobs6x+7aIkvPSieCAmsEF43T9Z53/b2wp+ZH8dxz4Q5FZxJi2wc
9/MC7n2XUiMm48BLrfjj/A/Rmjx6wrfmNzJ3knydN6+T1pGD0yLnyfp6mwexeboO
WXuF6mTCDZshBD+K5cfbwdYiVvTiWKsZ7aeJ622tebtBKyNiq79lb8qMCVYfFO5N
nWSrDH4x5x5cQR1vPc3Rsox6mpaMcoIh/nNcOVJc8yrDfnA98XDwXNwRcTeJbXBX
xkb6f5SGgqVU1MMbVira5nReoC3qxs8yd82yZV3JMEJXRYHOxbtNN8zHUsgB+Tol
hq3YetLWcORkVX/SSbrBwgXuhjluoj6INj1LDejvxIPZufIjvBMDeQ5fca7g++HC
4nXN738duhAssBBwP/WmtXu40CPP60NcbN/cvLTwrEUOSDyCoLwj0Yx3I/v/dC5X
79yvctchEurjvCSbbKl2om23DqR9eb111vKLxS0EDob5BnkeKQSHuuDL86ttDEwB
kNwwgATjrKi/NLbIl3vpO6jlhDK1fS0LjhbfKxP/NF2GjBSLmVllzhZNRoqGy1Ii
zynMjTEstFggxuR7vthIa/8NJo6SSZLqjy49x5WMwwm4B3q0KmFVxg9aPT48Fuvx
hurEJDspQDp/OyUbaa2x5erKkRf0avbae/u/2GSDKQcTnUI2oqXenEza9SbWYUEH
WNHETh/6opeeLkj1coWna4Zi+hQAMRojRdLmX98EKZoLDrH9sMG3rZxA3EvenguF
bVypqlg35pevjkVkXRzJp6E5uFfgvThaP3JDdjlz0HgY9/wLU1k5DGn82PpVxEyt
sOi9Ip/NZBOkCtU3akxVKtcUagx1ePTh49gz61Yam0ThwGECPbUdcU/iD9VgVB2+
kzvISP1fzTorQkqogq+5TdwBTa73pdkG5f1nUF6F5rvOFm3xg3YFb6eq/ZYNafI8
by0U7toM8AM6kFGvvY1Vij90Q1cgNswncKMVw7Nyu/qpniPQFcDhmqhqR1IHx5pg
e2BM/mBZqRKrvwB2EB53Y4MFLXY1AUdjpj/bbDyY7KhSUzVpIvgP55qVZlpy8Jdj
b/Bew8cv7OjhXJJVKGM6ImZsRIQuSE+v4gAw+Ik9jsFgQR3fnEtGcibA257Yr+zz
Y1bRJD8slM7aW1rO+ZeAzqOZJPaeZlarTBLxYcDILo94k955/Cxx3j1f5Hga5fC1
8u7TAtd/64Kcx0dolbzlLhWaZJRp5e1DSf5z6xGtFdycSAgvhHFwT6Kp6N6nbi07
d/H+vcqvmMFO/thhcshbeWABtDVlWk1Qzy6bUmcQEhNhMmCT9B4O15HU0LJ09c4Z
B04kGukRY+ei7CQeke11+KgBqJ8UzH7iPT8ewkKcQgmyPtRq0zXIfYDxii8xHcFi
0RJhFo/e8yy/C3xODam3S9EWPuF7WYLlPHdVrFVoDecu8Mog3KArN3MX9qYweTQf
isn5tcSVRu99G/RQrYb94/o7d+v7o9P35HxaBJY4KW0VgVqF62i6uniXXs9gZApX
T8qWZWTjwm+1nE//QUILYkbPVD3otS7QFIXxUZoeDyjANvKh+E6iq6EEQizJtDbB
bp88pDSWnjAziXH+eTTdP7FVdU84aBskIgcAXCNKHywB5YWcIibYlQwqJdV/7Ko4
CRUcD4heI8AEZYuECt+O5UF/XvR7ov4hSuNFAgBjPxMt09atBQHyBUA7UzOQZJyi
ZH1vZ1+hHAk4yD9uGTjWTr2OpgzCp96dmbG4nUAkNzBeHkSRJK0xoVbpCCg22cfv
ed7zjgNOZ0HBYb/nz56ypHJn2OpcypnIb521W9/K4ogWNcialB1tIMVHBWM8szB1
Pn59so4Hvm0iGoYRfph6HaJMHH4dNolYZTK9FfNDTw1IXdaP1/VdsjOxDppZxUYM
XNc77fE6pialH0Kqd+eGelkdFogESwkWOaRJlodrtlWMq/Y9ZQDfdw5mlrpQmiGh
idJGFLJcDbqxIRYaInO6OHd+eAJNJsfotKm9htOasf9cnUcJ0brgqqbRdWqCrkGk
Qe32ywKhiO7+kmrHWHKwOrAD8yMAOcScwTMNHCzQycSMgWBDiTVLtBpPoYxhO04b
EhRcNq7yq2LFSc1hcKpqnYI9mTsQacJ9ZnWOdxUOUnWAMWYK3au91+Dr/ghID8q7
xULEBYgyDiK/wjNZl4Td9HFX/xHYL+R8KayA9HL6SroQnEc8ayjebIwJcAwcTRKN
DBzQJ0poUVRKlzADx6gHoIKkU1gb+t4kGuscfLy9zsxqJGxzu8nugpPIrikhoAnu
t1p9KRban4wN4GnU6ZQWocE8zG3h7NOoVcn3w5r2ytRKWtzrP+uoN+RqX+B5EmJi
m4PyHanimXLD6mSA5Yyep/cieM3hF0Rpf8A/J9FSRoHkOB2ibbhY5YZKBY+HlhXi
2euI7ncgoM4yOGbfEduQ70VeWsVPEGKgaQYx/3yUUAszIAB+nQZDR04VmLtD8OMe
+iIGMJUIaVTLSGnQ5pr8e0UbfbZzmfw0F0DmPhm1PDwTkQYdV02HtwTTKzhH3MWb
3Th5/JhOoNaU29/KPkKlIZUb1jqpsihtQ1tUHTuVCvKXkNt6DZJJF28tKvxYj45d
jAFRnMk4P2TLo9dCuiodL/k2k83AKeoOIJDyB81iEaFMCmlBdDZiAFTL2SgCPO8U
hjUFzpVECH0FqMVXDD53rUnOqYwL370CNBt/m70xqopb6qSQPWF1UuPgWzvKudny
JGQEwUshZMxkvS8z1dPPI8BIlTnmffRuXbTYLLdQzMsSVrPxzgUxwawI7NxYW6E/
DIp1YsM5HBv0dF2mY8XauSAHSunr5WT5wJ8YQo6XklEpqGlSba5VL6Hyt8C50CR3
vnRuVwWGAdC3Cyjt23Vf4AF2eHhJNnWaDtL+S2474bkI0bzZY5Q8v2rx+JpsAN4X
Rm+jf5QDn0Z8pT2ZeVNJ95vGgi4rg4sLqgpIq78h1h/hSC0WADpP+R9rgAuOjsHC
cX30TthPv2dV0bI3n14OD1wHlteZlztSHpl+ocT7S1hKLmYoWZmZjypImj21b/1d
K2boZ35AQqN+JdhgCiYm25y6CGGoOyXr9izYplhQFMtL9pTXB/0HaCOOqFKQ23Cj
U1/fj5zf+2V6A/kvQBYv1aI8hbrOyyuYlyUF54p+WiNsj12n/zZb2MlzwxT1PQRa
k4+atCea/vBHQd8bewSF2Qxz8lmFlYQK0xpJRC9f4zr44/HjcoTk4+LHfqErC+J0
oZzlorxWduGkZ1YPXb7GxI3AwS3Cp7XlfLHG4kFz5E7dfADRd5fT6IAcqUJpgkJ1
rAAwQEw3cX4ezv/JAtGiLwyAIL7DhJ43qL5L4cVerIsKRj2LsZcg5RpMqZt3PNbd
VAP4sGMoFb/3JYYQzDq85eH6F3w4f5I92GzaetDVEuH1qmYLqiJ73mPGItaHn7/R
fTrlYH/7J6NvHM0Fa94J+CSpyp5BRuX0KSZVKTq2Ym8Y9ScNsFKUfzlJvFYOJEtj
ZNh+YeEbegiQwbKh5H7zyJxH/qeWaLJsDFzLL/9HGFACzkWgKqSjoq1UIvzScRwO
LRga2Vi6T5Sy9Jf7j6BBUM/omIg1Ogswplg0WjGWIen218tCZVhRvBnEOwLldx7S
IsKU54vGk+xKVFFrOloXZOXn86lut+QWTisvHPAQVNIlBw7lmVuW/kSf7XruIPAa
F+rx+mrJ80U02lXEzzMylOD4bvWM/27z9vNjVbnMbFk9VYP0hFjEL58+nFRebZHU
jUqNEfbantiH5t5OurZTPMaHhbYXMLwYBBI63T9SxAf8Q9wbGe4xF1cs9Dzox11E
JYVz29M0pqTnRXxBGstH7qIGBJvzhUAgawdz1eg9JQmgt9gL3nXYNhjwoX2uaTRw
tLdGZ7Nl+iwxjnJnTadvEvbC0LcOC2bM437o1l8aEhV898ZyD+oqV+v9NDAW72tJ
7m8zmVyDmCwDjBz9O2yRiywcm+9gXWpGoiSckWTZ+WyV4+fOhoumF6fvzEL2mH8y
yp0QGfvodF0dwY9apSETCoFk7mPWCoD3b4/pk9w+W1Xy+n9hc7JXuPGWJfi6FwBp
5NJ5j4/5hkIacZ4n+lNDkhavrXmF3yHwq6WKvPGCYW1od6LxRr1EDyqOgATEsr2/
QN/1P5gR+zOFi4seWmCo7El/2CnlpfatGxZOlcds1cMtxfhW3yMom8lsxMJDAIyQ
s9o4Uw2Y9KzCscPZ49eHBm6DQwPvd8dy0201agYsZ6ghDcR9qLfBI+ZNEDRJvcae
5jMGrujPuKllR4YFGvjAWonBrmEXloRt0P4TEnumHfupK3Fm7xDXeiduwXcwX46M
sVDFX4P5M+rIYQ6wlX11TL5aNGHocrE/daE6bgLTmQrc1lvIFZLomvRaNKquMcjG
tNfz4But6z89L9pagqB0NptlzD3lw1siG0PiE5BmBUN9hohpvPHETyooAkn5LDnm
bjpkT1tMzqLfcpn4PPwkj24/G6uESSYFWgXjqOrdBagNJJCzgWGa61pEplckFYgD
whcThNMdEyy46CDG+tnG248q3ww5w31PX0fbzo4vQmLkFCOVbDf8mezI/Trv2qJN
PhMgYnsDhsjWjdTITzbJZeEjbTMt+KI1syO8Uxw5430rjZr2FZXRShMe14Vne0hN
tDnnrqeAh4DXc6HnzLe8JC1ouopaPF0tdq+DdR6Jq0EmrHpCFX87RJaHrmKkgvXd
w9Rb9E/2n0M6n+ZwYEqIx8/pW/t2rarHbUiZZzBUoishByFabnbD3TLs1Z3Ypy0D
BwUqXCQFHMmL+ppq4FjvA7foIbBHiIrNpTwjzkSvjTraMnS85sqeL4uAx2VC2moR
aoablOJU1LGIui4rf1QVR3HIW94o7hFzvMgfUoziSmsgIAqX7gmDnpOtvH5n1iri
HVsiygHjTN5DjS6Q0JxqFueAtxnznjoDPWy2T9F1bGd3E3FLdi8mpIoh40Hv9yhq
z8kbAIV6+ChEwmZ/TUtd1Uywd63hzPAYAM5Rc7P64WlRz8Ohqg4c52k5549I0RB9
01lUmO6RGqSahwVD1wpG9JxmMWUX1wDbMkQgkfP7D5TYLlrGjm7q3ULN33+Ws/or
Ke9M/oh/LkrVcBUoCH5iWRjbXZUAZ8lZ0EVGRCslP6lN0st8ut8v6c32rmt6EO1f
MAEFRFGBYKeOhrp1kEGXpjeqfhp0sCKlL09S6Psnk8CBUOvVUpMzmZetKTTqL/Ro
bIbySJb2UN4OdnYt6rLX69dd+x008FWhOWBbEl4V13mo1pxaQhUTwPYVWlAc5PSQ
p2XSlVRgU/bcPxyh4Xu+88WzUxL99hVCQ+BOC/GOjC68ZCtrVoapRAYB2j/OyePB
PHArybwcuE7E040qw1SQFVQx+TgFwbRXvivpXiJuP3rerkemFPmbAl4S9aAbjabo
00tJHGzwsc2dhJWM2K+OGDv6OoP88HdqzRX6kMyYjy18zGbB5DGVdq+gBmiRfP+X
cClNa1W1lGKM1o7A5PVqI2MeHce//h15C5nFdd+ZOxtcfZIy+5XVgvqfZeQcIr3Y
M+PFAG7Gwzn8ZxvBA8oKkYFVN5LHr1fjGGvsHslGCuIcyd5iublN3nrzpZbIGioJ
lz+BbnvgGbNgJGkS1jsG/LwY8M9HUq474MJqAKKdwHnknP2qvWM+V+pmzz0+qHxX
DZOl4pgj1wEvgXfiT8kRnjBlLfre1we8Ty0OO0lVxGs9PLg0OudRRMsbFY7cFWeM
fWS8uqGylq7F9hQkUOcS+hBhm4qrhvqEc1yectfwJ5Hhu4675VcCRTf21c4c9o98
I07Fsn3QycqHGmx4qLg/lGyT35yPl99mrGs+C2D2CgcRgZ2+NLshg3H/ih0L0eKx
LEes38aSYq0Wcl+rICp+qn77Od9fcTebnB0FuUlu+8my8lKwW9RRYOkvEndApSIF
Th96VdDDDnqqbpCe4DdziW+xytK2soMSZK+gFOW2uqgHGcRvWRwJw/+xOqHKHKGp
H3jM+RvFzVhrEG3GFCzWKV5VnzdIFQM5XoWPNn47fZwPnIoizPEt4nAM2CZKlje7
T6GcRB8cpXrGW9f0+wgWu+AZANDzR4f9oN6EyNZj81BsysHQITc+Mk57QjaLfLuI
ATMTzzY+01H59bmFsnBtnYFrYiNHpyAfExLDUqqbxy6514WGz1NGStK6RTxcTxSl
IZ6m5goEeawCG3BhXigtXtzdnvKibvRjUlm5pWWUaqcKrnjxuJI+A+KPMm+cNz6m
kazrTL4l1Iy+f2iBoBp4ondWeOOpglRYC1cxBCwBGGX5+O7JSWGX4pOnN9kn7z8w
cf0bXVdO0uxjiGRPpV3Rc5SgC/OFOD8OS+Cy/KRo892gJ2EAsyQunI6l2mbahzik
l/PDHVMf8ZobjoZzFqnmlprMC4hgGkfyBvi9Jpgr6cLZUkFPAxU5/D1mlSR8G+Ki
AkALTzVS87ncQ8NwgjsAzAE+ZbdnqWX3tkxI0pO3EhJWrLqHsobi2VaIaOt6V8kJ
XbAvjhvX7y9iWl9Bl07Lyia8g3Vn3Jx1DCMtay3RyWnAAR98fseQuMURytmcrpwy
bi2NgbFy4+u7/F+QWwIAxHyl8E+bUWQ4A0jr8kd1FGzbJbWXgWxK0j67C7PhksLj
VHG9wLsLKG46eSneXbFhCKh6KsHLs+94NHFQI2CIkCqngsmxYoRak+vhsLeJFQc1
+N+f5gae97g5ZkbcflshXhSsN3d+LN3dEu/Kr4XstyAVaSQXeEPiAvgPRiT9z212
iI/03GlftD9eOqbOuE5t3qYF+EXxXmuExDTbBspGlVljaAG+b9zYfWvi3qDzMYNs
ALY+586tGi2U610XDZh8SpQTQ0hzU8Q27guqV2pluVZM0fhql9kJzCXVN3t2meHG
DKofPn5JJW2FC9c+mQhcexNbuPTzoIjmv+0wLUe0IY87fXESGcMEXx7g2iIpneTY
o0Au8nuSt5IV0xbAjsbjVzjUNDbE5IPdO/Z9vPEXGVQ24bs2Ygh5ZxWj8Lqd71Vv
BDho3JAwz6Sb4Dlm2ypDEYDAWEutQ/CyiDGYyXpzXYEIteXD0FKHXFug67c9KPa1
gu7DBVObwLCd9eOV6pQIBO9FCtrW7zY3hQFzA0zJQUtWhMv5VN6wHMnM2Baur7ru
lRFGN7tlZw38AmpHAseSp6ADwPmg0x9TtBEesfpgUcGCchURZ/2p8X+bId1tCUyP
jI4F4STo6rRwV2cBFaXNzuIz0un43E0g9lIR2UtTLvW0b+HJ27ZCOfd90k52nf4n
p19d8VYtihHj176ijYy+w96u5MWV/18i9to01V42Mus8bf5CErHNUMiEj3kMbIoO
ECDeTqFAhlRsV7Pg+HFGbbcEP++ElsHUDl4jFdTUJVa+JDm5/C2eWZ/SGkFe/Rnr
DJ1fprQucbSb8WyYVORw0hXSEx4WiVh64z7B7vLLmrFoB612ujoItkNcmJeVHRux
ZODrCt30v/WZlAdgL89VuIRhQ3oOmBPT08QRsFYzhN8qQyJab2QCx7zBOaU6Tp7h
LwZlhdyKprzVoalLWSH4AFKTMR+hV8p0+nIVVKTv1xo/NtUyswvFFyey8sIeiY4u
7zepJdyLvFdP9q3XH4lBTewrA4g1pDSHZ/9Mh61Ip5bwk4htnmHxC7T7zpJmrvqo
1NQNAEbgrcCjdiwmGAWgsH8OdtxTAzqKVNkbvdo9LBF9Iu6skz1/3rgxOaKRdG6H
KRSk89DqKQcfVk0wteRakuhCpHLsE66LnsGkKHg/biLBLzTqhWKteDEqy/qyocTx
h7idS1f6PnKg1PtMwSmetJA9gUSrzRbCQWmwy8lv5SXT3jkddTKMr8FiIUX6sgZV
bEnzQCLXrWUIGTO6caYMymq6K07NS0bGiFN89/TjYMJCcxGfCUFkKH3vcCzLEYqe
FWGQy6ya6hT9CTyu7vbuFGk3aJnbXAsrrYy3BnkTVYTlDcD37+gPLrzuarphHXi/
RwrpP2kaWmIKV0Vpkf4QuDh9+j5Di+EELo1ahAJbsRvuvfH4CfOzwtJUuBufn5b6
nd8wXf/gkYux3hEdj4UF3zdDsV5b3VeyyT6W6HikbCO33Qva0ZRCWWDJaaRzhy6B
6+73wFajbgDi+UT4eKyuZexSbKmINHMyvUAHNXGc0qoOzDwPzfZxJhXw9pcz0E9G
UKdFvYPlTzE29Ejn5xtvPDD7nykFyaH1syls6/BIdt/CJ5QshdnzVeBk6qX047H/
wid5YF1ZdQ+cXcTIAB9iVMzDOZyx3lHIgEU7CLMgoGisNyWwN9xiwDyVNMBHX+za
mwiMorx24KiLP3ZIUMPcmnkr+/YQ23RG59aAVswhpwXlW1kThr1HRF/1zPdvKGwq
LFyHobbApg2Tk/cdNUyLiY4KyTkLMHozSSRFVOYJwqzXSYSMBwyKYf9NP1Z1LZc4
hAfS31+U6wyGZqMao9TPdpNEYjTU2QxcFDAatfHNxjtZtY0ytmhH0RVUJTckV7CL
mgox9A6SP1ASD7WjuRVVOptWEWdVlSKcNS1Jsrb1ObR0FA4434lb1ehkdWglCxLN
0SWp8u05M0UO2K7z1CYnJr+SaJglXOoqpCrXJMj+8SgL4JIkwInIdYah5GwqNNvi
nzy53GqIZxA3sldLx7rXeS5OEAThMw5fSjxo/CPfn+J+s8aWPkgXWi3Wm/CfQLxC
c2Ouc5bggOfthMybvsd8asqUIQGiWcYD0q3p31yDqNAsMlX6GiTEjHM+ehD4K8oB
2QDyDd89tXUlwJkhRWS0P97NrzV1mXb8TgchjpAIu59ZMWBHKk21H7FeDASmplAk
2UgciDDcNF8YjXYzrcNhgRxKYW6NYzntTZE3mbhcYibvrILj/PQsoKLpqE7jMU6c
OFSwJummLDHkApWskQ4SrKUGWBINU5YieokaUZ6b5FG8fJx28mh+sTTXJdlK9PIk
U0RTgO1Kosimy2gnyzP1CLTO1kzAtUnFzD4LtEhRSgtBoSvSktAqsHforCCmLTZV
fVC5JhYQjJDY4NBknQqm7lI6y6QUNaNaPcVGl4BcQ/kNYhKdaeOG5TA2s2zIXyFS
GVFw+SkGnIrcBiNKjAfRyDNCmhjutWWWobuipvinABdksXD0dAtYYgwmQeuBArwX
zIb4OcAtrYbKyMJUnTOzcLqiX8EoO8dXfWYx3PIrX77fTSM3cbcaEItDINqyM1qA
axRPTNGi01xwVz5JNTZVu/wM2fQjDxxKBlmqsr8cEuYrZPzSFNcF9AgPyhAtuYQZ
ZTpEJ8NSOCzT94gWMR9Pr216Q6SwyNHk+Jl4icAuaWiDeBvROO0gmGr5VN56yYUr
vrCnIkjFur0jLRRi20/IM9F4t+ZbJt6Po6c/WH9vLZxKi78fxQGCTxBzE9gKaNGy
02Ekixi43YNlDpzUmGm/om2Z4YSYg58sBzHefuMH9b0Gc62iMB06j9dkDHVx1BzD
k2/KOE79T0ribSWqBsXTJpssAw/h3uLKwNpuh6FMqnlKyWPQlMQKm7Cl/Dw9M4Bx
Wo0hMky+fC1u9PblVyIEquIVvdzINRHAFBRMfAv3D/MD2wehplt3yaDe0QIhj0t+
N923m1UYFC4mPaLvghV0LfwaWl3VtOM9PA405gEghn96qKN2xDHsIJCWvzGF7Gs4
JhhFPRoollYpMCNrHTKMUyOF88rc8hJNyoCiRQkkkScS1Rlcn9deJZwiHRN/jLTk
UThxcJM9HGTMC99Es4D3kadIKc8PFd0hvP9/0kzIkTienCKc1KtcarBl+cp6Hjge
WlMef1PURDbSdpN0MNAxJNyVdCbsgLa2BTmWJacjW9VLLp5dYhBcDPzDnYZFqm1m
WGfmbR8se63juInHjJz93dbOdsT4jU9Ntx2dM6pacA7MrykdpI/iQkNT/fxNOK5z
XQfbcFkrpv78/PUI3wCE+OS0xoYRWQhMfbxTCXFw71garDO0mgvIv6owxEww9CCl
1A09OI4/dSU2+iuLSjowqomBQpBj0GKj8aIi6brj9hLfCNt7FtMV259H3y5gE0j6
ObsQ2mrZL5/gqniJyHhfYnqsI/PL/TcYDTiDBGaVUedGkjpPDXr/BtGbjeW+O6dd
Rq68h2SRUiPaKlJPxnYGThk0WHPWXVeZKoH/urJ4OsJ5aul3PiqzKfciyyWk9s/H
PdF7NpgCN/i78o2qnmFrJdxTBiiM9Rtkus+5HN55+iLZ+dxNWRlNygbkU/IWhCrN
kP4vjN4MP847Eq64AiN+z2BB12lZ3pQ7axhoBO0kpN56R6npU1jSg2WlLGnOVkN5
/B313tlgdkJf7xpojhSKdAUO3seHKa+MV4RehwRxWl8b2bgmS6fPANtk28YnZAwt
kPqAuIpWrk3TyWyA8ykuwtdw5dCaRgQh6r35FHf2oX47IxYtWcSA4jGBa8Lv5k61
TwBob0KihjaVq+0Q48DyfAW3T5xXxHRNBhiNcH+UXikM/qi2MwNTl5uXRCTf7XXB
c8IqT09kX11bYanYCmrlONq3dZpHsG5oBI2DiY9CYnd2K5scvQ2CxhsPOX2uEhfK
OClRgRoO22xydSrl+jbqw9sKLP3dnlZboS2vpD72P+Ppi94PdtgdqJ7bqyYrboxq
VXulLjcFL9v7jYp1fEvuGr4SnzqmXxbq0AOJ/yLvCsoq7/32SuNk4ZaNHoq0f9+C
s1FKLNjpLWuDv0VNyZ18UKEWTxdTUqRurDAH2UUkXe4NrUqZetaQdVpW2PIP+Vqz
ikC6nBKsDBFXhlxzBUvYiPx9lP2lxXUHKQ09y+gXK1o9VyuvWu6KWCDVBXgCNZoE
CzSxLSe4Wr4nXUXdWHxgxxy0M24qHHRfTMGbvosiAZ/G/NBzggB4ALJur2b8uoVx
jpu6+Ft6LxTC/8o1F1NroBdQ2h7qm6ogwM0D02svz4QMKQq1ztlzii460geAz45r
TIusdM0bBCgZb15O1nAzMpFMRNKbPTrkY4u7k4f+IY1gJ/N4rs1X0FSoEki/rbRD
MeUfT3LiJdKeaPqgQoz9XNklpAgUhJF1aYReqrm1+3sKmpT62DvHD2C/OTbCwmk3
KkctFI3+c0fdE9CSPZ05wFWzkieYSLrhtslKo3KxDBX8st9CTDPTf+CLSHIUFPx1
bwoUXP8oZ1xWaI4lp2Kqh6gCCBBOzx83bAcQATwfUAihuxqUoK4SQjgZj1gVEJMZ
iLGfDQPFYU9r+Eow0Jb2umEXlh6BGC+BZWHtdcXLntWbqTg10wafHmX8emO7IgyB
8ZinWfEM9KVvufVqPONv7tviNUC5FrWzxhEC9WeNmlshJbE3thSBN/HimqIvAa1F
ur31peS9AcHyjYaQ+N3dcj4lfksMY0qydrl0k+t4ju4VtT6MqO8pK5COSi9G3cSu
D8CF+lGXLv56URhTuPb+pofVlxvbr41jEFeNTHMTaXfStLoqNpEOoGKbCT4YiaXm
aillq1UpYSU7sHmYXD58bNcpDJ8p0JOvi4O4Lk1IQISlXpgqYPkLiUTHWWKl17iZ
vVFZCJdLi3JHyTY+FS7KfUJEm8YmqfKY9c6vDjJcaBRheHLyMPdFTfi7cR4yk+1Q
KuN0RxwffGNJLHHnW7B4uAh0st6imthQqw8AHIZXDfKfOb+GaZZGugdhBJojHNuE
WNG0lbEOxg8looIFVqVnSqD6e58rza5uHjaHhGJnfCleAHHNccSf/7ouF3ckMAcX
k4F1YjBmnlBRcPR2q96tnybcMHJDZ0nchhIDHr3O6tr2AGHgH5YvdCCbUSFkZs80
r4kp6PJ5CV/0/dIF5kyiCmwB4rsZKSQp9Woq0vkFO9hrJPUjcvfE2m1CJaMivlhn
WIoE3pnwulRcMQyx7CwTWSVY/JDt7RYcI1USwlV2GkcYtSGLLd9k5vuT6nH0BfwQ
T4c99TzJYnFaS8DPVTMbpeMV8gVkUW8aGJta+ZO/EsZXQsj9lRUsh716Yvcftsav
AxFO2+SLkMhSZRmvLsuZ9iCfWQ2fNVxCPNU7sTvw3KR/viYUE/upmd5nu+HD/sgR
JVfJ08ioeQeubEoKo0P8BB8Vr/qV9295gUq8A//YA8CHScXxHCQQO7JKEp57qb9y
jcdiZoFQghHPKZhfsBM3TEDFt6QwipExnxwogYIrnVrl75jojWW5FFiOh+mPrqgH
aAThQauCNcIaxhR2yWSezvz/rbH1+W7ZKPP7nlWJ6Baao2UoOjYXLlOIW8OUx/lK
zljuc+d3Q/pWnHXvBTJl2S267TzCWbO/ekI1PBOx8Tq4jKi+6mUOZ85sEpWm8zqd
ISYbOsutWs1hmS/cijILUVsx2orXJb8HPQ9xNCc57B5qqOJG3QBzDrqORitanEXv
ZGX5RkbzPL2ba3J0xibW2YrqFLWKwM5RZn8+yN0PfokV9omKcXpTTeaUPsUeeaJz
jhRS0VpaP5JcYBs7ih0EFpbcsLkvcF6A2+dFyvV1uvlOdiAzCtFYn0oHAKgKlX8N
avKK5X9ozVc+ZcJ+jqJXh5z+bFvtdP9cIj/SCXrr+7+bErUpvEalfAKAOC0zWFKD
9Uf02t79RRqE714Yvp//UxIhTpOiJVFL0drSX1jk7faKKcYVq0F/EpUoU3HOLVh8
ODX0EsfDfuuFoGoVPNkjWSv/DAxlmi4nt95RCWmczVE+Ume3Mbd/KwN/eGow2RhO
9UP7/KDqt4j9C/cS7qm+D4p+97g25I7bSFHPjt6OrikwWXXjdqf1CI2fOBbwJSWm
J+OLFHO49uYM0RjWfpSLwTM/RQ6YxaYYKrqSbJvbFaBTHATQdPQfJ2UQEeuVxEa4
amN4v26sJv7UHVtBXFWcEGunRnBZV58bYTxRsSDzYVAzp45k0KP85A+n2hobL2ta
rX1Dr1/25Y4BY6eK5pbYyp15dR/KOaXlPjHVLe8NPmJwnv2f/0/j3aQ/Oo9NpXWw
0rgi1EhRuo8g0E2KeU/UCqVWLD9P8ZKcOF9yA6E287iX7fHFB3dJ4UF0/FbFy6t2
nGS/AQaR23wMDjjiFd9kFJNGqicW8A7j5WiUP5MHqlDBGq5cTRayDzLVV/itfKRO
3BP6He6Es3TOIgXQMdvJmptlPRJiC9nP2CJ1UxHycGe3F7vxs1GgU+n5zTWTebqF
1oBoToWvcd/vzR+HYIznLjPKrtUsgu+8KEmfa2uNEAFqzLLNLDNCOaZuDAafvrGE
sHwkyzA0x4ViKDXNBh7kK+efVsOHmSc/W9JIbmS2qdbb/dIJZM7wYwzK+rYgYJXz
QOZGvyKH3TFqF4AIbOVA8efhb+bGC7L/JUq6DeDYSy1vTE2rG3o7YRyzaUppQP86
Z4H047lPkGrW43iKmPpQpu1YQzW6lqymPVO8lM8U4AkmPjgpOFjqOzr8tyR6y5VY
wv8F/iRV2B6NezK9SUiI8ohgeplNss+b6xJSCyi67GqxJ4NCrEPWsNLjCqGlgsRd
2XJhyrFH4apnSuZltNjYl1dp0r2WOS2lv2UPKvAIHbIkfOSP4odKPlqWTdantHMD
9jYCeaR1iPf23PfqUSETwDvywfbBekC+CjOEPGN9/y9Hy1ORLSnGISv0FuGLUSvV
01HYsQ6DqmjYkrrGOcRSlZyKGJCItq2a8C0uSIFWbe4zioINT+9OObwn/REZd4HL
qzroFBhRbkTEkw2CwqehdHPiuTrjzftOgnW/wKWnJwTVPLn33Ev7x2RHprPLtgjl
euWRS79+0SwFvx0MCu+7nirnaJUeg5fbf3dm51OhnyroW4w8ADoyQvNnfmWfFUxs
31aPcH5TWxtYdYkVvxzhX+ZH5sq7Qbp6tQjyhGCmB8G7/ZU5QEQ79rQA+NFX/mVm
qdN3Khsh2fWxe83ZiwTNrspWcU/9PLTtZqB6jJuMlDtQkchhBjUg4lTkOzaG37SR
afJRNcLbYgXbQ8QEotGAGXArj1gGiem9wnkbRhsBUYkeQg7i33BNPmR3W1M0DrdL
fc1BGZ85JEP0sHlZWlCNpQ+Rg08yg3aCWFuTT6SnHtZhLnbdaVvIR0nufiwjaRF0
8fcpfjQH+ULJgb1UVG/Mp7NiM7mZDi1Vu9qUZBCS9tRJDK/IGcbtfxT52HH6UQIp
98ZFcS9NKtMvdWoJKDbYjzlrkvJellHX/nsbpUl2a16OgJpXPkDJRZoRmvmPahnr
i3bWQ2Os+3JI5cFNngiKmvg4xQW+mvniwfHaxAroSLheADHFpEPpm8GFNiYrirOU
740UuAwv9CgDbIgRAhZV07lqMpX1ehH1tssVnmEXC3QzoSs0lEAHd4qSeYj7m3lQ
2L1XWx/oMCAHvsLDS9vrky3RMjzFQdKOH6p75PDO2e9tZzVtGJwFIlaTSCZHy8Cr
85NsbUDqhxGBqlrhvBSEiqu4LLdgWEiRQYytCwgAoX9kl0xdvLk3FwHBYJjVYqnC
EZzjzZgE5cVMt/KYi8RPdnSiFD3nFiCoyL3b2y14e0NZDKcOUrLQ2Zun1SjrrKRU
VHZ/Eu/UQrjP48bi+4UOaBLxuk4PhXsIkOAr3VsE/w9saxrEd60f9ia/QFvniJ2h
TaMNuQ96x1Ti1HqWoqKiMY7VlK12g2Vdp5PZ7Dq7tfw34NJxEyi7a/Q7ht/UQr7p
grGlGbN5BbbzQ2JaGjl9iH4ZLnFn/eH7uA3fL5OwtF0ojkDfJZ6EUMiuLKOAIA3t
bEDvNQxxBYIKgJ0dLCsvBILzmOGfDh/q7aaMIehFEBKk72qpVX+OqgQt6HytXN7W
q6TFYXt7haXCg7a0Cz5ZBwxQlBU3s1Cfa/UXmcs77pet66XkFm3ZAY/gizjiJBrM
8nmS1axiv4rgBagl+j1K9BC8gMdo+TjhRMNJzpG8pOUfP7eSGLwMPxDCK7zxHvG8
Cpyo9MjjiEqULFvq90xXGefGt4OqURzGEwn169j9qnkCWKjIu0WtwleE997LB4M6
qej2EkCkBesoFJJYsYrGiMCfSzWPzU1D209khkl3KObOt8Fr87SzgTcG1FVL9t4M
4lZfbozTIwRtkLEcxbpj1NWEd82sXM0glV33Bv7vGwXDwdFa7mS15k2qNjGvmo2r
vrtFmSYtGFRYsFRsHd4v2jz7rLWXoTXqKM6YkG5azgbusKHaK7tL5q5SVfBxWFc3
z32c9mveqZRxGL+4yK2QLNsyagcTV1HXmZCVqr4Q22LozMbkWa9DSWdePOogvzOB
jQP9X/ACMzTuhYsy7pGTXkH040zYz0V9pLBlBiFr4tpW0onW6tBWjXxLwLE4gH0G
IzHqz156tYGb8Ria+ITfsgTBz+sBQ++i0qcU/elEzQJb+VMfUFBNtuzQ3QBfrrLx
VylRtI9iE3ZH6XZUopAiwLXi5YspO5Gp71cx72AYz7ZdHQYODee26sXHhn4kvUl6
q+1KWY1vM+wnZ88g9imxfpY+T/xG3ErCHl9kAIlOZOl47NqB8b8Mr/mYuAmUTTRa
G0TvoUC7Lv7mbIy81XTYeGUaH5OUoHM94BgMoTS2d3hC9rVHw+OJeCnYZTMuuyJo
eTS5OLJq16jcjfdDYkkUKgWloLXo7dIoGwfiaRqrIKn0KHyGUPsI3ckNCGhu0V/0
qL3iByiX0T/scYx1rEYA6xsbg2DzNAA8AHfAjT+uaNxnWPqVDoZKLYFJBnVTI2x8
a3kqIluvXjl5fbjV6PBWdxMpAJXnlruuUgsmBuxhVwf15Pmb6ZJeiEzA+CM8c1nv
H1LWsSBxEkaYrykiLBK/UktBjekbQ+7p6IljWW8DLSY1KSm/yYXCqEkHSRdnrU4o
BfLYcxI30+aL4vmyVPSlzMpK2dOWjBuOANj8mrT7vSuYu5RH7Yry7Ndc31DZA3TE
gh9S1N3xHzbV9ODxZJYxBxir1I8Ud5Co4DvPxumKrfYf9NItOb/N3oJ64OSzkX7W
F8CXH+UkWADEuiR+ci1vmmPuQ0P3F8AZVEtsDYP8HAg9qwyLa/ilAnsdBDi4dJBw
QWCXqtp8Q9sBXPU4ikEHB7yQwWgFLRuo0cttzP9MB0BwnCHwwgjvaQMAVGuovPSP
fvHABQMBoWG5eYRxhrLQMt5sa5QlCT/43C+bLnTou91wr7sdOPrVVRIsX7SAjCAz
tHH+Q/OLT63sharXqHabx0OWg/StPH8QRiL3E+p9pn4sE8fnXUBOZEJQ8jri5OBY
fzSNKkopkCisJy62Mn8SPN6CK1vWOCz+Yib9SwliqmQupC/GEkQMjr/74iK4wENR
Z7DBZieuHkwzytV7iWsiz2VzsRIMKTxfkf1LTgq3GjzEVr5HY7WfEdaKg1GzRHtc
KyvvwliiHIdy1WyzrR9LhvsBYvfEUDA+31If/H4a11NUilJow2KwExDHxJOQeARa
6WaOD7VkhoXzuh1BYLFUZa526rX7Mx6kvNDtU8fVrZpgggMhh/7+sN3MK1EQQvOu
f3yNSQpU+QpnrA6mQbIuGUFGp7J/zwiT4XTF22i3j4NYh74BUDQstDmvGCViasfw
Cq8lERcnu6MQYv8hNOcfYLob5ReY+9bb88MKBdJEZJIEF1swtyjSdBOhLSyqjwqe
0LMw6ATfTnNgYvrb3IEHr0ARwBDdqwprHVUmzvz7JYWfCPTxcjXruOHptBAjC6S7
g2DyppCFty6TMNqbmfT/FDNp2b6Jx8wT10TF7BeB9A8l0o4s1P2OviqhJenq4yxu
cLmIYHhh8uMrhUJhB0BVV3cAnlyou52Sw6QIRFh82qeMZV5aPf7uTojjdENF3Z57
SFBN5Q3XyFBzgh1tFJYrz3SPA6EnWulekfGSvcQVC2B3+bLKmhHK/XvcpsrLHtGe
H+55B+t+aO5i7qcAyRClfpMQ+GXtKG4dYEOYzoTOSAAnWIuaH67YqgxgEwZquAmF
QlcUzIhOGMnEPtqcBeVsM2jEDjJdVMfRL5pttS6eDp8xqQXx2vPA84k5xsRbI+sL
R9aFxGYd51E36bn6eIykrBin+C1pGybxmNIbma5lum8nq/lg+ZoZWAXjLjyhSMV0
/JKy8RTA+aZjPAcmKvOO1Yl+tikbiFduCYUmsPQgh8vj61XlLvxL9uritXm41jDE
JS9/4U9y9kZZLIcdkXaGMZ6Y3X68iHRv/YB9ioe1ZQMFtmH8uuZ4oUYx+ZImkv7m
6xflvccOxIp8ElH7a7LJTIvvHab6wDWVJh16zolakruYmnb6Djkro4SL2Xeq3xup
hrVnE1E2fv4Ow843wwGpMWIMuJxAbZTSahSLx7RU+5d9C8HPoled9sVyaL7yxKTW
1zsRHjpp0EfICVG0ZyOg0LGgVEEropAaHa1/jHj1ai9hC3EEMtEwzL3kpYG21Ik+
FNA16D0w5AEjFnZDv0DC04lu6lnaqPyquKvHEmTXWR+yO8XqKECRjFXYNVPEjbeb
UrTvw6UB/mULVmkgh181W1hEaxAYKoee8UVl+CfLhcQfkZlogXylba6py5POW9o2
ClOsq+AKVXIKoLyqj46zxLJVfc9Ypo6IV/rE3If5fLLioke5Mljfcsfum6PCJ2ws
zM2B24egOhBwcLjOB9vLaGcK3UVYml3NfCzkrlM84zl2GgXrMG1yQE8DnwHGS7jp
k7mV+3d5Ri2BwWM4WC+ZgrNlbIxgNemBo1tRMqI3OgWq2AF3GnnFev6zQS1w1WDP
UdzxhoXTWz4I4XvKm1tO8ApikJSf+IarHSCibnKu9qgZAUJ4S2SerwyS9K3cx2u6
X1+Beu1pbQIkqyYMl37bl2sUs2yBCkofPeUlTvG98BlNC9U0AGFviJ+wdIRGkOZ0
d15aBnXBl1G3fizl3+p/t8WwQ+fNzqfHWMGLTcIIBDWg0eEloK/nqDC0zQl+v366
AtHXHmOeDi2nGkY8yaiWYMKws5U7PppwjwRvUobXrIjeC9r/iDCnfuk34ZHrVep8
4uQQwsTlp64S/3m5q0j4ED58ZYXJk/CdVwYhKVJcz/ZyCuqx9k7vbNpryF7LtpAc
7Hl67CpfLIdemAob0tAmYumFiQBiJzH6STSEDLcXDjBNVrGdMOrK4RrYpZzU7at6
Jm1bQ1+9rRMsX3vHSXJ2VJkvG9O+CCN/kNX+3kfDIsi3bShM/Krn0wmnGBgTxyYP
R+sdwroFdmX0gdDKeGatx0ia1483N5n0u3bFFZ+d9yHA0ziU4kSn5RlrUU9flfqu
xf8dHur9E3Htx9/RCsSbiC+yLn/1sBrnLi/w3GXlq+E5yMZKtKH65k8uRVKJmVbh
RUq1oKx2gpXFBrPqJJZduqgJT55pD2lmXKqRS/JTr4Xn1yUbaKu5l5RXTR95yzEG
XPO4M5gpaHBEemC3QWLuO9xGyF43jWkYXU09HpjGaFz7C7cZxKFblzabziu5Gwq/
p9qJMHPr9uIbiNktR/vYJV9sN7nGtYwtIZEjTtERcsmyj2KZqjWTK6QpPGhqyDT3
dA3v3r9HLdlzO/Qk/9/I4wGXkxj/cMvKTBNY5Tv7Ul8hbfpVECp0HMqOorB2hLwl
BA/IaZI+3hPnut0HdfKcBTLGr7X6GquzITjyaFjva6+MFTimGca7EfHp0Lo8g3Vp
bYsOeVjvtZY5hsejptrQwUGqJPLISlEnJIo4KzTjSxJcvclGaC+whYCQc1YOncLY
lic3V7gEMPP3H92IpR6ByJ9nGiI8XaaDeOaBwbDtNW320cj1AWA86kR/KbQflUmi
/J7w/h6jT5r2CmVCH2BmCxn7Qkqpak2DJR5AO4+mm/jQzSc2murjTW2b+EDPCkL9
31ab3xv+3E522jf4Cq6tVlaCsnnNA2nEOMsp/+662f43AkC7a2BE+UHZTMGusuZ4
FGl+aT0ikrX7bsOFbYhuS79ctjPN2xyW/hlBQyZe2fV+rYl5N+qeu3Yc6FJXyJYN
2grytjgMF/MEYRwY8rgetYNTzKP+a6Uj3cjAhqmXm4TjRdbYbJoSpeFIIkm2qiaV
Aov3W6B7Mac9B5MdqwiOW9EBv2a4cuvQKm7Po7BVP5PvOamugFLNkO6dyW0LAMCI
rNDCHfADM1dZJ+3QHmKOY8BD7mbvJJnY2KjOCH63QsOEWR28/xU0gF/d1aiiv5mF
wKpFIhUk1K4wJCrFZysvjYVKEYKpvDUu8wc67bsZjFh/K1h6EJKTI9fdoX8FsO9b
XX2Ekf+r+9wNl0Q/wH1ufDA1meYhCFkVkOxQXirsu5Vcpv0GuRHh6iPpzS1lSA35
/MDwdUFFWi+FiEda1/oeik6ZDS19Suv0y5+9lGB5vycF152JhH/fW8BXjhrwjvJ5
S50pDtF2rd4Lcgq1tCrdnXvC2f33Z5wlpixaaMsXRCA2ZOG4sww/gVD0PNmjYpd4
EfGNuHl6nsgQ85dMqH0cCYg1/5XRaPnNv4aU/JNmSM6YsPVrNeaW+7RsaVe6Ka7m
hwmzEYuC90PZpGx7QXEM25GSywvCObXgM1XGuEAbpOBtFol1yu1ll0ota6M2TiVl
Cw7eNaEwC8L+e05STogrz8XbE7JOuNRLn3xWyYvCJTuM/2LI8K/qoetk9hRe30VV
vpYm/2C8u5o25+ne4mNMVyDiQHc/wj3NMO9FDFaEqX4P90BqGwLeakCmR7ihIOx7
S9dJmF74bxrbqtQyXPZ+OctBgqAyYxZ4r4H3VpAjBgvafuuWEFibRZ5wMoDL8AR1
Bkw9RL8nUTiTH8we3MdjYTY0cMmsErxoNBO8012z2u67s6eiNhT2jvlAZaqdR8nO
VqoRRd6+3/Ya7wDB4ojJA+0DyyCRLPNgcewyfiDUj0g9gz9JdAm2iRluzL1YgjLz
P+XY0gs8ULcU+ggy9FoBmSW7tebKPoyr895af8TiwDG7SjTsc739ZTIebqYlgVpQ
rE5PWxnfo8R6d5D5aIRMO2xgUc7J8PLdC1j+k9hfl1roaAWuRBRyHH8Yfv3+psJa
WlJLJaZFw/hKAqn2w+/jbARyHFJDlrNt9IheK17F+kwA64H+bxszWkzrA1yRpcZi
RtqffBcD58kDC3IZugY6T1atEyhi1PjqNYPGWaps82bnZ2VZbX/aew3oJ9VAxQUR
5N4BI4oOWMy2YG3hicheB7qxx+/i2kKMKL+VJrT80l9i28aLRD+oB3hCOzFeLOyd
Rq0F0tSmHrowlyoaasv6U+YW3QSArTP0pN9/T5WlcOYJC/0ResXTVETCaLJU2P+4
R+lRi0fXmtUfWvRFdzbb1mTH4bgjmqTSn69+po6C27nyRknDfO0Ob5TrYbBdCIeI
i6wUVUptyUM/oTchBpZfVkKApu/8EtBBddm7Zlyi3rDwLV9xLK4DbtFjcb/GfatH
2p2GnUDHKQBw801rqWbqSC6diM1eGqzdyX3t5Sy1nzR3EYkA9zFRsT37Iw6nqvMd
FvFQBHcY+HwmbfhreOJEJTJ5+O3Y2yciiwd66JcF0z+Y+WIDs6JEUF0yMWUyw3Yi
nZ9YiCEp91pL6IcioN8JAfwqrrYtk4Kwi+23Gy4yZPLuBG3MnGfhi8osEESf3Sf+
e8FkVVjboNlRhZKjHlyo1fF9d8pYCbVnP990cfrk2vz+2ZGkzAqOxkB9a3lh3KR/
bq+a38a0lp/ViJaQUcdLmqskaJp2f0Agj1q/N9MYf8Nphj7wY+Ey9NPqJSLiN0DQ
VPSdkjKxLmGRqRipD/xi53m78rSX8YnsXv1VFfhinHHoRSRN4vg0QETop+TMdqgd
I2Kr3hmnOGvRwfJ7woh6rEInNFU99XxNiQxA9K5O7pW5NXAfJrRXBwAFb/tD5E4x
rgoFByB9f/sQ3BAq1y2FlTrD1b1sQb40qXyPLhS+ohfSmxThlqyaIQBfWeezwCbx
4TB3ZbNrcgwmid0QN6gLHpF/5lxJoZ3mX8J7v6tiOYjA+NlhlJ/H+pTKRIfBC1X2
Sm/n/pYmtqpA0YuyikPjwgTJYFKo0EVn4jnU72pQ6mUOu7pe4sDL9E3LessrHQuX
hHpWgqMtog8QRvRg+sgm7qXUcn4HQU8CD+9h+6nT+laGum0xpKiPjmIkDAj49h2G
VdOh8ZoJZi+OeKcY+0v5AZNaOB6ijQzzzFF2SAWsbYbcyJpFdkUwJNtnI9eWei2K
+aTFGrFMd1kzhUZbisCMWofPcuPhavGb7/sILV7WfdgwGKBiZQ0aPGfn3zNAUHPq
j/tcofxF5xPMheXIDZZcH6GAHhkB0fYc6l7GWDu4M9pXX7dODCh/6fBMkjyRow+M
WdQsQgFZ/V7OwxtEJpz+wultVh88LHP8ag3yLh2VSGsuLgYloS9EedIq6fGKLdcR
R3vcTHy7utuqnOuOZbP4kiK2og/ZemWCIHdXVXTjlAD98903lwP35mAmppfk27D0
ZSUaK2X+0uD+mZzotsIDErATjlsV6sS5TIm/+YWwyiSPVXaaB2e8oINN4w3woVQd
/fqO12sysJ943BYR9w1kXAQBdYPNUTYn/MzmnfFasFhXurI9AaiiGW6xWa35dD3Z
8TDrqvZEPRt6wummAVEZaorfax54KCsy//fd+6K3pOnb+qdvaU4Rdr4ZEbeOsdca
EzPDOC31V6tamf5AhEid5yGObr98gIajHKsczROSB8cgtVNMqHcTpG+iIQUQlcnn
Yz0iNUXJmD60CaLOOSz3iUoajQvlHicq5CefeU0JONezSv/nMu/RoZleUQS1Lk/n
XVEX/8G9O+k+H1bBluRWXsxSgStFRsy7PslY5w5VR18M5g0Ou6zm5gFp/fEu7v7i
UhTmZ+NRpY1jSnSQCdCCkA0rwkx4eyLtc5/PQ7O0CDUZdNPsDWEu7NnWMeMLhOkr
shpQ+WPYrtjHmOuMBJl3efUjbAgIoLI9EGNTHIkr1tzVruoLpH6ZkNj8Vl0dmYtW
oTt+tKqmx6tmcXmYgBA7PKmtAUPazoj5IvocZjzuqHT9YULEK2VlsGKzLpqYMuVG
R42nA8RxhTHehRE9Cn/O7Grq7SVWXu/DCch4g/kRJ2Rm862kWPtCDyjQeCYhIKO7
qiaLE27pZ7WxrcZWpncw1cpiXIO0Y1ve2m/0iFHqoe5Gn6Gnf6fbkVibtGQ6iHlt
JOiiTDX3fIkJEOj4ewjjrF1Ag5YjnWxvpy/ARkJInn3Rppl2bMEIDBdnn46E6rVt
8DVexFKY3XcDrGFJFBARS+DC2kpWGMtWEHeF726c1ct3ZrZz7DWtZsmpVq7tlFHD
cUPZAMrugH9BiTZqTwiTyO29fqerZl3GB83Y7p3fyQhVzdjcgzRZB8+Dc768iClG
MbiSHLmf5+VLgo23cTbDRLlPOXW2DN9NVphqt/7zwVJ4FdMn4My+0VfbqK5z//pq
jYaaf/zSL6cW4ANwD18W/7IYgGSjhISUCpvW7X53VBU0homkvI6lrIpZjoReLQSW
yX8AN+N32YGW5yQsxUqZXl2ZC+PoVPqDfR4JHK81mb0RrG/g3/R2BMpwlzY5WTr6
yg/HyNbzM8pfpGJhWbDMng+qJTM/ryaN61/CNNIZOt5wRwz3IkBgwAkOV3h+7nFk
BP7drjqqL40maCTXdxL6KwUfgstgjBFZx+ra5E7bSLjG/QJ1cuT2eKsZXaJ6RNuO
5fovRtP6qan3mQl5TLRv0Kv+BY1JSlYJ2EISlnhp7WYRDh9u4ZGP9z01cPwkHF1g
T9c4xgind/+H3mTJWZ1Z8JC0YHWET//MfCzWuoYMKGi57z/mjf9PAIyAuFoo5+IL
fKP+83T3yYbbGbnaHuthwSfrRZbLcJH/rM7NWI2itohpuDJcJDEWIcEzk4x2cvp/
1LvYvRkHGbhz9BtJKiHM3KuNaFA1RnX/ldcp+iDqf1d43vlFPvBQtxafJWJIjP9L
ZWBA2Cbw357iW1lybexiYpgwvzZ7GQJYJ5ZB7dAeFw4BLVXoGWw3LdTbxk7B6gCU
KtTCCdZDX/v53GklCjbr/NRI4iunGedAYhpArn1GGVdRllKsKLwBcySDhyErBlxu
FRaYDbpre3A9b+7jQvQifeaoou8iKzvTnWK1CF/+LxHgOFnTXZ1tbncoptEusFKR
/p6DKl5I0moCHEufKHq9r0jp6gKEiHsrEmRMtGeXcgonNEHbW8BvNf1Z0Sw5U1Bi
A+FIpwDoGvU4OWfRsq7JhuACHPwa0mmddfiKl2vd3Wvl2N/NCV+yydNtVm7pz9Iz
oWZvIe1h/14WSKB9oFDeP2lWo5/ZeoSR9TIdz6jlJ/8yMhOt7C3cXYD2oAxHhAN5
0HCKmbrzjevVmy7g5Y3LPBCcOxxTk77KW017d9gKt4bTiPCzeYIiMP+70G1gxrAY
ufLB6DXHp8pFsPT6Hh2xARkcpqiZbUn0sqQgOJz/eOeOuHl08OI7DnjEDVb2tl0d
9Ovauy43o7S6zHLQgFmHqmvJe7cEbDcbe77SuPjxJegNeUp+3ksRAppHDF2EqEDF
e4TkC9yYQZHdepWrBem4Z6U5eGPvDJEu73JplO5G/uROH5A2aaYdEZ4uPdB786iZ
tCos7A/bTG42bab6m4Tu3R9JeUwAlV9kLQd7hYGFSdaKaDR0sxli4PdTB4PAXOlb
hwb3yE6c7oKZZmcvVtaFrym0hwYotvFr9ZdE9q/EGAC0qY9sWk0OyaXPvN4yevrr
mxx1jYHAQCqpkrtolzoIYDMp2L5yJOwoMuzNN6b1MCVsxFMIKsSxqKnvwQwrcdi+
8CbEFZcYkbHlDVAQBCxdEcoNGflEShKxx3SHv7C2TgOHzjjBJWAEhcGk5boGR6++
Z66j0NLOmwwDrIILgUOAqQ12arT2oapL3KQYxzx05ruZpuJPXUkqyQVLOrxzjc9M
3x06/8RqGBySVvXeuy6/3cW0tLItIdVoBHfSViBU3Mu1HfSquuPRJnF0XQRBR6tg
XxgVYEoaSNUuuomo6k25TgDOydEEXlP6qwPUrcDwESk8fflxQ93WNhQBxYJ98KF3
X5ZSRseUg4G0bynEf5WAp4ehyhHBdP/hymjSbnYCe75e2l2cQPtdmZfXJ7L1Duap
2QWl3pfg2ZTiK2Dyw7+0Kk46vElE+foy7aOz7bG6RomcfqT1p6adQmN5CfjZ5wNN
Wb47VoWowduolJIME2U1dM3hC+XK2isynHCli6tNI81twbPedZCxsA1iPfO8ObAG
I0SRyx4to6aK/TKY7cNnRwoU+CCnjfanhKradqGj+aR82DbNzHiUk34+CyVNh+kD
SnnyfvguPgeYqtAvggzBT33DzDxftwOwIGn+8kCXAPs54HJ0bCRRuGl+YoRppsAc
jgu0vxGP1U1uizVLL4FOaai/dO5aBKYpT6svJ7grxUVDGeof98IgbKxUiqtaZleX
Xyj32NLs0AyVh63f+f5MOZqSWfIWKaN2MQgWKIiGFtROxmFk+EyEUSWlhDE+y3ID
Dpxe0sgnbbOeV2iSvmFiGOQvKPmMVTPcR9l3IeGOVG2nK6//GhEFIviKdCrYuYLb
oG2kjGhQZ4NGDCf4r7Du5Wvk6D4xrshVVT+t0/KAJ2gMVmVh8SRJlGkab+iNX/I8
TfzffKFUONHbitUkVhRok/ikD3XZjox2f7i+akloIxCebyYe3gSK7l/NLMKwf0ch
kmH+DwrytgpW3QsmRf1V82MqQF3NlNQhTDbmHGqeakn3aTgxosZ+iCgWj8Uv0OJt
01geowMq6DIMw7CFAGsPaVvwB9lDdteh3TApk/aNlVVpdQpoCuZhFyiAdMDzHxh0
b9kW1L6zRA4IWHy9m2SC/S6r+p6JLydI8aLYGn4ZCKPG4g/Gr8HmEKVYRDhDYkLG
YTFah+jbW2Hsrpy0+Qfel/W5YhiSrVfefFQ8FT3PCTxyjYoaY8Pt7SbaGBrK1W5U
14vit7VxAZd6sa5BNx2owvHaf22wLvDlMDpxhdJ2k6Ig820R7/7dtIerc+C5/Piu
A14XIralkGShS1NnhbTBI2LuG0LWfc/TbIqDgQJB5dhLuLv9+Jn/Nl3Vjdn9gbwq
Yd3QUrVX8pbUa8M42vdukDdVf8MukzbqOOJ0vI+gsSS2mqxB/r5uHNm1nDEhnmsL
1ekYKWusbFDUlkFvUL7UY78lz0oaqsiPD4hUqiIgHQbDaxyLTjEnLjg156bHIpX2
cYaSALwnxL2QY+1v7+gmz48els7byfTFWYAy7tXK76okdG3I0zTPF6xMhqMR5+FY
iNC5xdzQU27F6Wxq1BBua9vyWa/Xy4E6NAapw2yGxEr8EBO5y5ifmYyTQZontOLP
iEki/UIOPxczDDNaMkul41c3E/m5E6Jt53Gx4/IhbHEPLn9uGAoEm+NETab0RTSQ
v3rW9XBi/JaC5m7pnjrDaXDqkWebWJGfr4csujahUlfGXni9pnm+PW55WtwWh6Ju
YfdcCYMUl+T9mlCax4qXxunX7pKOiqWLO2zEFsG/UiuwbXge7mES7qVqD4W3GpWX
3Z01WjI6bM5Hza0DK/03Eoiz9hNc3Q87zLs2h/tg/NrFUIJg2Vs5kKX+CZn+tTIC
73dEmEhvfRo34jbkUqVG/eRGq9AyrJ1yHmO4mmY9vbyqLuSts8vimsCv2pGX30wr
oJafBx8PmfWNQCPAOtzmYdEKfSwGlwVp8aLDH4gMZaaNez47UtObpLPdZp76P8IN
3G2BXAZik5uA8G3VMQ0oAzYH6+uNNKR96AM3lslKZEeL0cd2UETMfe2YW5VNf2pW
zjSuvKaoYrv4oE7no1z9LYEMkIxRbUgTrNLYkf1MccORJhHI8vQ7f5/ugur6guSC
Fc07PYgyyKMOuhXIiDI5/03BEhX2XOS6jMkWNweMZEq3bprWSi4Y2URTlh956hCb
WBoh3TJBr0Kha2NHWrr2T9geAhlGi18Yu6bwcR1DLLazVAdyIRSTRFxrbQj4OuXq
7DXt75nDJ/LvTK9g35SCTzOt5B+BygZe6ChinbE0igautCLDRZn3/TTqwLD38WrD
KNjhrYdq1H21cc9FnUJ5wQcKmSeKjOB2sEP2TL5ZXgSyCL8655KQuu8WBQc8sxIY
DaxlnO5ED5wNDcTy9pAUbAYUvMc08Y40LV2uBgp/vWrAXIcj5LmasHY0gTBmbEV9
6DRCjBkqw8Eb/GfC7vTPyz6HUvLbleY8jx84Ixc2mjNeXeQ8CKyldHa8h/tAGLIi
Or39AthIX5Ll4KCqq9cgtRMVrU4Cyc5ARceloFI4V1VRcXEsK/iT42uKYU/5MrHQ
ngGNqVAKPr+T5AQgLTL6DQBux1QslBj8eGixr0p5t7QWK9bgxABuf9ofigUZDdIY
VTb0qyK9EX6ZZEJfpXcCULjRHkxrh9Yjjq+detrVabsLi72eBvQypr4SYMVhQ9YX
V6WdAglE8A0Eo6s4jkZcSkKwIE7MWW9CCKvBy24oQKXZ5KHGPxQqpKLc5DDGR/0d
77rEIYlif9XHxjxzr9nWA4PazPwljVUOZL2+nTMhnvjzbqWn3zToNJ0ZvlZHus4y
kN6j0wRrHJm+m/0gaMK7sGaMFsH+GamjFNosaDXrYq9pug0AAS+qHISQk0N0Y4FJ
5x9Xe87zJQvMf67xM00YTAEUS6jzS0JyXmLIlmdQbZcdA8DlW6gYguHsJzUf4bVX
6htKyciI5IZKi3uLO6caV5fi24NkS84jxwaWyUjk1pFc39Ya/Tp86IAUd1WsgR4Q
0GVZnT9fnq45EvMjR54sWb7i/YLC44t5jGVPLAsog7LNccSWZSh3OTmVJSrpPdTA
Y0Qf5MH+BhHbtU/x+RGs9a99rSDZVXeaizhB0KaAK0TJ3YclHrqmT+OCRFpbDK2f
i4dphNZah4VR54CtxpBqzW7V2o3VyrzfhaFMpMPevH1dycg6xo+QpcM9q6hQ+KTb
jzueQgMUvq2Dtyizt90IU7wVpNKboYHzl8dHENsYGk4Vu683jdSMKPmNNS/Out0+
KcdXH9eI8AMH+d2u59cHjigM55Uk+gCp2cuP13k0rn9jRbId2+lrflYzJUX/qf4l
OjkHPYf7597KVkEG4Pe0owJMdh4D4jNUFR7ZLVYNwpCrJ+nek9FhaHfY3obZwz0b
6APdSQZjTMR89a+4CpMXCEutxPrWw2x7Pi0Mqz0lVddmvqiWvro6k8x0Hi/bvbAo
pxIE0ubRMSJiWIgrtQhrFoReVVXfjTPLubAPKY0nJSiu09SP8kaLsCAbMhFAwyQo
iqfr3b2CNfvYFAfDUYgFZuOdAMf4sfqnNUSQM8UG33c8uRKeNjgaATyiUXuO7PpF
jykQvEsKhdeXfaaFqOGG/KKhMg5p12Cr0b9W2c3z9Q/hUvdP0eUEy2UQ7v9qyL3v
7gKvzAqOLUMjg5nx+bjUgt+667wM6Asx575JT3D6kNc49NBb9q7aGlWieSChcFHL
iOgemzoTmmWaxTEe+36FR4DlmmP4bw9dQnmBLBVWOnEjamRMqlW49DvatnDKW9nb
juw3axSzkqQMPfJ+GT74H1O0lhNHnuuYEa8aA9z0NgWSciArDJw4XhKDDzGnXMrZ
4jqYhMB18pXyABaPXnv/dA8ZBZFh8nXhMDryB5asu7SL5k+y+meS5sZcq2H09tf/
WB2mhFZjw4JIhriMlBKbiPNN2B4MwpxmPZIyu6aRJd84nceCGvrxX7wcdIove4QT
w2s+UCwp8sPKxey47Lfd9r1y6WCeBWnfdQLNi/KGwIPBAjSOO+kqkOmZ+a5s+9iJ
VY1hWbT7+UpgBprGLGdnxJkfnMkH6gpezSyXUjllfPHS/Lc9zeDlVm9L2NZ8xfRe
PMnLEP66qsdDwUMqkEqp01vzFW7anv8oaEiXGWJXfCkTwab90OqGCosgiqmSIyoy
T1oO9LfZ5MRFK5/V0aI2nELu0IH6+ggqCmFv9cuCYE9XJiCchQSDucMmK7ifQcbD
+CDW95aB8gZurT0CWHJg+qgYGV01svb7LG/Mav3ySKnhagC0BmlZl566RtNcIO6u
wTSsAzTdBvvv+w9andozjsHFB7/XeQQKIJcEaagBfd7koJxajfTUQBHD6EkXWihL
8LXrSs3liM9VB0ZzOaY+4nGxQXef8aWDhpJedc7rTUBgTaQggOp5xxA5nRF6gesZ
m9ftHLvqdQvRaOzhVedXypseu40XiY0YK5XOjeiGtNRHGfq11cBTPI/v2J9lhDy4
heTRD/fvjS4ldsJPxFNx5iEfOy3euCPcac0yrc2iMPykv3W5WlHyM82AH9a9rFqp
OKJNWlsOieoKXn83/17LgGlzqC0+4C/kzhJAVaadW7p6oL7gV6T+NkliY52S4dzp
8gESCXbby32eeTp4vs8N8Ls22bgn1P1oXVgJJfLTfqFevwX/5A9J8bLp3Z1ZFZMz
AkxfiVvsRkst37QhrLDmjhytCIRuVB5okhwbgKd6JLCzOeh+rUD0lHk504v4ZnFk
i8XaBO9nkARHZzhDBJ+5CRsUegPG4sr0gsRm4HQACNt9DztCJYupeHA8tk7lX8c2
dtl1v7cCN2/7G3PWbco3qKPbykbRITcozgwrY3dID5oYck2/dz0XUoSJVlZSLBF0
AvlM9+T9fGsMCysvVkDqgqQS3TQ/MYFR9ogKM8OVl7zDQKmikQV40EkxPVwr8bgq
80pYyWuo5OY3+so+oYL8OlPAiEp9xJwCGhRYlokg1gHHE19ugHQlZbvESskFktn4
1IPNfHiBoftDGT0i1Vq4+RwWyD5wFYXnBjn80uJAsNC2xZMhCkIJYHIEZDdPNKva
1K4bIlmPM7WIFVY10x38tkwCoe9YIlITnjQkDAcbID7OJDAnex9/Cp2D24Glb3r/
PQ731z+MGh+ohMDcxz8F6xhebsyfo34WEUY+W6I/Oqu/idlDoQkDgJGnAjeTnU/s
fIZ5E/iCwJi3KfhMEWn/itazvKHYOTwSJ+8/bDBq0jmAdNRme7kiGeKwf/Z4b/1d
Q21HTVbHcGQ88vbAJmazU020HWhxuUH4em8lNYLqEqknRkH5gtQ+FZ70nCJwc0ql
HJFBljo1QKSyxsD8dKnsrsd5U5StisOwOCxqqgiT8Ffq2Gd40CFYthK0uwT0QOvO
WxgJJiRdQZaLFU+ZSJMKz6AOWzKRKWdnVzaKte5hAa4HdK2Ac+W8g9wmgASHJGvN
3r25Ar5bp4HkWwtrkfa998vmSTMfM/4sUVyqOZvUOuxEZzBQ0s9vKUjmgNRO7ZRw
jy+3l4x9bS8W+m2whAMbczHnyzaaEPMhPzfZxK11kJBOk3LJs4I4xjXBPt2LlS+y
wXsYvoj5MSXm4g7I24SuaRIfgnxv2Li5g3RFHtzVcvNUx5p4wzQI4NBOQGObYUHz
ElcRI+PZ3om3SUA6GzCKQLmsTBpYlxPIMspCzPnSqjyiClAJdrkUguNwz87ka+eX
zvyBw0rT14wVgSeCEk2Xo2UzQVThMGgzGIt3K5dHBNZpvjlPX0CsInm1+n1dL89V
WaGfMpf/gb8nwbQ4sJw98ZbElwiqjrLisIGP8AlhJ1V0COj12OqFrBD+enzz3gep
zXUsuWfbwysmh2eLixa4CEJWGQvRSH6N2+M184q9CXzqJH8DI5ugCBZN8+1Xx1qC
8xmonmjNCjSjAx+bU20ki3NpVkmPLnZTNqcHlxpASR5/eGSQz3K7gQTrhEW6m/3w
k3ve1Rb7cywFsZvk08CfL5yH3+9iimmYNEeTQVt5U21bOyn3D3LPXKe5WctzGKt6
/2atI3yNmX2RxSO7UJ8C5aXhMUeiuvF1/UcjnE8JZ9MTnJCXM4jhyldDiDiWEI90
`pragma protect end_protected
