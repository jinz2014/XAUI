// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WF9S3WFmiicELv3I9K0oi3UexdMSBdWGedofK2Ep2p7hTD44DKrNg23NMgN4adNK
eCGQ6qOPnfMyxfheJ46uI50nguGxB+q923pTS61Hq7vCbZwVJDmCf9SvJv0XOjaM
NlXwlg1EYZkZ2xqpgmPtKpttUi8cDQO4NZiffarzmiY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3808)
W8ORDEQHDoeEHNi8aDu00c36OgRlm73x84Ym3c5OqrWwOTwOlGVEVaZVpdwbz7Lb
xPdn7IllIVMaS1I1qbkoJKz7NFDkQ86Qim48GgSCpfG9wRVTDsmBRl6S3hfpU9Q3
oRIiGMsOZAttKNOJWmOHbK81iNFZIQ//v8LUnO+pSyhsWwSJ9iJ6Fhz/WPSU3bPh
k5AA4gvRcup/MhC86b+e32Er4gyCYnC1LMR5bwcoVAWwQvHdtvCu3vRkQnXwjsS3
bDTfeuAYQv/xDD8nLYS/iXakJknRp8GINMeDVCQ+6tlzRDkJ4GTyXt4KbbMzfjFn
UFUMnIAdLeIpG7B1YDbH6WC8KU8ZMy9wD2f6qj+8jHDbAC8vluFrdw3MC9dhQibI
qXTGc7wALO3E1H11a52Qj4AXRrj3T2VdFePpuo8tuwIDC1eCbE8I9wXBJ6RfTg8v
+mRHE3m0ZuXZ1pK4uCTnyoH3QmNmzWrbx5bx4NddL1leKzf1AHvxVCielLZjQcmD
gYgjDv7hG19wdYtht+Z6SKZ0x3GEzB8e1BICcmbhfIgUnJ8mLu7EZ4A4lI71ZuGh
5FcEs2upi0WcispDJ1Uw0nn7vSkUAMLBqy3xuupaZxng5kKCda8iM1XI4yEjfNli
KimQXIzr2hSDuo0ve0S+3ibUcGliVORAKHx+c2TOKp0S8PCZ1Mu7kg2nLHUST5+i
cs8GC1AwwD2bRf2b+2A/XcFQa8pULiX/OBTNhr80mXsYoURNqzjTkJtrxc5Fxv8o
5EmxmQp6j1rRoqDJXmy9GKRnbZUF2sd2Vc/A78x0AI8Nq7zl71O6bkcB1w0FfMxM
4NOGvpNYvBeZbNUl6w5ppanFrcSKfKF8RUlRDmQOjyumylN86oBJWYIv3i7lt4Vp
ifLYadT2Y5nUoTldNpsob3NPXVMng/ptto+2bBuHefwRhS503DL5VsogtfQZgGIi
4wCjfvTntYxasxqL6SV6xvWviRdNW31tVqQ3JI2lsSqMq9qu1sDm0AbRwFvSKELT
nv51AbMgg8GHJImQs6PR0BWBDzpFWLw6pZUvUacukcoHtyiLvvIgFGWcoS/OrPG0
etYH50kJ3Y4R2gidgsj3g5zPVCPkq+asCAO0fCJr0MVXo+qx5yitZc1mBFitPtPc
1XFc4yAkYCVz2A82sYNG/fAU8evjeLTQsVDpBxI0h1giEm1q6n39o1rR0N2I4VYK
JH+qU5p5GSEOt0MVQPzGyRZVPrWFemCvpCkXyYWlrAaimrXn5iyYH3yWFbKEqVkU
kzzRnNzlKP3J83l7+5EuiZpP+nIGJICNp0BgXxEO4zs/8kV3ayB5EcDcxxKFBF7H
z/DDwpWPGrtuPx5tsEWivPgbmcKqgvW1fjrR8xhed3fF0WiEAlmwWJOHzhuCDBF3
jH+eYGEXJsYxXLCYSsM3etGJjkVtNBQVPWMPdB/Mk039Xs0l5CP7eUatj07aP8JR
71WWvHsu+Z6qXFKEVqkxYuvxljoOTqpWfi0R7ikSKzz/Qc6VTUKGS/CBMB4/xxUr
RD5iDXiPPp6sgP/WttK38J3kFxeOQ7JghKIvjxlmrJ76oE39VihaO12Mn2gs3PTp
pj0COjCKA2lgKlCveKfx+P/0OjI5EYWsdeudcxquiU3eSm6jm63533/nSVQUkYNU
iuGvGWZtj1EzzLy+R3X1gkE+PMw/FhLTKP1PE8Tz4+YvfQhhnrz4OlAYhw6U6ppw
mIZb+8Ju7qdGKxK16JBUif5EivNp3b+xvjjEmbmySyAnqKikuWEEUBom9j2M94NW
09+RFsskhdZB+KeQAdIwsC1iAyzAKM8agkPo3ZZjoRBAlZYNCxa3BY8h9bn9QmAB
wUh9VNv9WVBlzAsioBcsrO3EIO4Me6kuaGFvokGqQAO69ZVUvVMmN6pjAfmUZSC/
JSJ2oh0xxnoadc5MnHQLv9yvtsXbxLgHWTvqxUnv8dt8c2FRQ+Hp98MwCicEjSFD
X+OIcPcrhzPLgrJpTL+wjjuCGwyuTp5mS1hhU97Wg/zH+YXa5P61aRPtK+4gQ5Cr
bg7ikJiK4UjBuDl+itdeylOGQrbAPEmeTnw8nr425wzqEMJXYHZDj2bHBtQUwPU+
TackZIaBCPYEHrhDfXGf4D36BZHvKi45rcWF6rDj01CzmZcGi9o2Mj+clcABbTKS
BfweBkaEEo3HcbZCjA2wxDvfQzIRjnHM9xR/Bd2DPTgneffognNOwEHryGKjh9qF
4MGlp5sT/zFxC9vi1dRHrVOzH9i0nntisM0BAbbHV/Zqmy/rqxfg7iS5nv0sYRgt
j42B7j11T7yAeSdn1yuX+0t5IShJqS8uFdU6l9TyIYeVp3sng/oc7vOX2dALJiE2
AAWGAg19Hg739aG5d6HOdbduwiBDnDuILFxnRoiTWtfX/ot7Zo3jrhE2tXTFT4XP
Yy2B3OjODdIjS/ckEFI8A5q3iPoKnwlICxkYbKDWtkMuDKvTiBuKOBpQcSzT1i8c
D28XOLbXeswxAqOIEmI8keofNVnAB512hVx/JrKyokkT6jGjpz0fjx08GKb7jvIf
iV5PspVLPbQHbKMox+lURrEoNbv5vfc+zSIN2u2VVYejCzJAkMqS4qyeTMP01oCv
JAQbmPgOpVkxzB0CBbbh50FkhcSo6bLF/VzrN+XmgdShTAoa+zM6a4cT3RRJo4Oe
PiEmNHjjGi9Gn2Sy5tM7YiB+KKPrGeST85V7b45iowkMIFWqH0n+rIYvD59cGmHn
ocH0rh3zf57PBNP9FqVCisjmFJH8l4ewCSs1FRb30Oc27QxUrQMCd1dT84+a9tvv
XizTPJsrGXct+Ke3VXtdxT/mQTqK7/U091XjrM42cYU/KrXUuhrrBZBIb9UqXyot
fOmMxvKnNjJVxupjs9jjCxfgKJhM7ou1aFytqRkMSWXTwAj+CCQaghM3PzpDdjuv
mXVTVjYxT/wuuTU5lMr2rJq2nFpS6uIFSO+uPWQBXDM3CavayvKyXedi2GuaPuF2
8GRMxakDkHNG9iSZETksjvDYJuEHCaXoJN2W7drQT41s6wAEhw/VoF+ULvwq1tbP
G+1dkrelWjcqQysaSiJ5Scc0L6feR+Noz1hz/rGT2b9JfUske7pEQeSOLgi5vh5y
z5my6/JGhm01EdRNG0z5eJZakLQaWaLpV0UM3Li47/In6E2zbGVOvsrCJtP7+vRW
HP+PUZLIDDMGJQhjSVVAVRKVowceAQU6ws+0gTHH/+E8v9BL9TkrqcOFDfGJdNyz
tajpWC+MyW+hDwSA6HJ99vHvdJ0kucLgcIu7TMmf6JE9pD5RaAx6fdntLuwGVZuK
iEoChZY4P2vetILk+8XaTEEabxkEDoC0zaTrA3m9H/1fi/mZrwvHCB3fDbRAct+T
jVoVtqByubEJ2XRaXVXixfkRdOuUy2yHgnv5ZSgMJR/dwm5Tmwjph+Qio7Y6ZmEL
QM0buWXDZClH0XHddaqC0FWR22bM5OZk59Z7IF4sk87GVrqQ248OPduj5VUab6Io
AqXtUP6xZcuiN7XttQ18ngfwxCvs8USccNHE9IzjPHsjsXztpFS1HsjjoMpkVgIK
lTQxn0+sJHDK8FRqd+e2f16t4uiox8Npozs0xjgTr+oGor2ePIAsBlPnV6dYJEIr
2mNR21DWZ6joSLiCudMGaDGiSCgL7+LLO3KvKLe3RbABtipO5Gvd+HUMRmopynpc
gMi08a5dQW6KJ3W13ivPOM61Atf0sjgeFEcD2pJ6OFBiWXtSHhhIIcRCd11C2f5A
RDRzpZtYOmKHTVWys0DdcEJ9qZgaqCXo0/ph6Ns5jKGm9SehoogLWQnbwULz+0E5
Bl+yN0dESAETDi7IIC/3FzgN+48k/OYZAuqUcttyD5Vd6UCUmcRLfONoNvAGhGLF
OpjMlhqY1NJlisO6stZu3T4ZknkO7hgY7n2v/HGDmmTfTcqlgjvnzDTDepML+A9W
nUZHEoqsoUuyaORQv67TfdE00HAHJVlG/hq49cPZpS6k7kV2ixAnkYroXMpixqsh
xEr0HAtf2t7Gx4aXFdNHBun9qhQyE3dnpDNzUa4McMcDCUxIQT0Wc/eRifP3yWmi
F4ulvgBOosJ2zvjSrDAIIJCLLunJlo8N4XUp4kCazYx7bWAiOud7UzFli2w6dbQI
BSeOaC28IlEMXd+Kz5hlqwKLHRUkx9zd5Q5+Tc14zz40oCwLNvo/IrCgh8Lm/tlZ
pEXcdp8qhBlD4pjvn/h/mgjRSobF0XwSEVp7JDgtDpnezkeqHV51auoPqnp8IKhb
ulyy3sg5d1gcu7+f+SRk+IQB0hsVYXAZWPIUOLtqyzVw7Bqf914W24cIg/s797qa
UNhYCH8h+4gtfbh7YVlbiLRIyNJVI3PrbPayBQfi+ZwRt6Pzswhbpbo9TlJy8j8s
yXiHLrowqHGu3c/HiJPrXdUsFImVeh7GlUwQf+a0YZuccEVri0CYT9VXnePq4t8H
F5Uw3udGXnDfIByhoStb80o67Q9BYQrWujdJKx1R5Ilmas6e6eKuVjJtv/6sI6eT
+moWAhGd10anl5MSAcFZJje9BmxuJK2jkq5455GTUhSfD/VyM/LxNdAv3Zq3IQKF
Ni+l7jVP4QUjodp+4oN5G/97fQMf9BbTI+t4VrI2NqYbBkF7YZNwQTZKnzKW+f51
8Yk1t99g8DvBELqBh+SYSmlohZ1FXys7q4lbt81v8rPa8L/+KIpVJSGCEwkzeW7S
8AKSPivc47JE+IJkbdKCYrHfDj35Pjtq55RAlTdQmi6W2WIuaVjvL9FSyzyifqKu
oXly0f/4yYfpv7eLvDCOL46YXGiehbBG/6hSFXwl/vxS44fkxFfm7C0TIcyjAxFD
vrHWfcWIfEKx4GDS06e/AT+nmsUNGqjHFa/ytWBtckjNggXbzCF2kZ/YBJEjSYFs
XBcKpHi3CHDTs0UobVo/Tr3ABQlROVgUXjdWBfSTKhDQEdfy8s1xim/RSObtzl6C
Ii4uqoBa0CvX/578t3IOiYatjhRILG0JzCeZ9vOM0hnDgFLPSLK8YqGaodPoIriu
b/4+P4vMe9HCWvs14dJ1BA==
`pragma protect end_protected
