// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OJ4Ey9ipSMlkhknOtPwIGjZxbGXbVxpEU04LSMcrCTVfqbTy9VyBYOrVK9hwofVO
+tTMuiem5B5Zzn6gOafz8TYACRaRPmEh8g8FEQT3XpzdqaLGPDMQ4tUBYd0EihlP
YWOTUdBlMluTLk9KHjbhgoelmevubdmrX4VClDp3kd8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8112)
RbHieayf3Ym3GXwplirYEx0WytEhYvE0MoQIm5dROlm6BKOcikJVruAbysfiHOtG
TOuJW7T55C/HTQnXS/gT6zQvAjLRrS/CY9i6/hUHksWs2fR4ndml2fR59yfezNlP
CwR4YPJCEDHvmXlxed00DKcHEBWEn7L7DLaEPKk4+VTMTjbtcYgC17g0wp6/ubns
mjWoY8/iVJvY306gaA+BFhEB9FvtFjyhHR3kQBifrCL/R5RCek1HC/xY3YCzCrYe
zBN3DeAKOD/zqzntqcXgjaB0+eTUWmdZ5TeOOiM2DRYShLLXSd9fhacpdsupHSWt
yy2Mtd6in9ly51wv10XD4tfCDkBTqEjCwzjW7+NRLX3IInJn7mW0QaQBSZPBwptN
dHnQZq2LJiM9sR/0Svo1yAElYpG69W3c98atneTBsTaq/KN2l4VGa168SxFa7NhK
qIcACU4Owl25/p02HG/fxg1ZISJE+mDrghBiVTlQYBNmPSr3AQIocImiG/dAGX0w
67+pzgl+J0lJSvMoz6rvo8msg7XrFcXQlrOPzOWepwko2EmUtX7Y1JWOUTnfHMdV
3Sx/vq42wg6IGigRxJ7s2anSPlvg8BgvLiiUpRB3BFKyH2hyzQBG+4x36NRITD60
cdjQf4kUFwbF/F551PfWX5DC5KpJXySBQdcaSWKAPnLQIqIk2fKn3P71adt1ZOZa
dU8dc/BHGTEE+8u+VcHqU7JFDAliqJoq2ZCdppMOZzCBlxIBM7s3UH7VEmTp3XJx
whk3zMbPVCSHReqvWvH2FD4Pufgfyo9bRfOw6yFvaMI9U9ZJDqCONB/nA+GdS3cb
DkXYQ3FAzHIzINrgRRJB/WY3qR8DgdESps43pjGnRsrXLR8LnbJfO1+sqfg9Tlf8
FaSlqfic+rOcNfYqmajB0lMHi5pywmHKV5TqlUlvxjgnCcdyQkpfbYTeUd6QJleZ
4/DyW4ZXYFV8osMuT8czBNrHeL+Cjj78gacnIHIQAG8Ni+rcAih5Zgn1GhjwqnMh
WH7cR7b80+H+imk0NKdB/RICvlXF3oC1HY8z1ILuxVABN2cm9TaX40IwiVkxKxTo
8F2WhPtOQcUmbTxn4mgZP00THF75WkeIRwrrg03q71Rm8Ihr6k6twPVik7EeY6Pr
Pap2mrEZtd+1hsGtDwnblUTymK+aUweoFjmrFce7xBMl92rOlrMz6qr/VBSsdZsj
/pYIAPMQEYU9UNnprwqi0EPvp8VOgubG4kyDJ/58bpEEkKJ52fgWg7xNY6RP+Mmc
DMMhfqyYfZCEWTq0oMa8FfkzQlHFTYajMO/sgZbtWpNxSFB/HbGmmaeDR8DDy75E
xLDVqmjsF9TR98+M19ii40vIfhActGx2YLD0nhHuwWW4iUZCx3JHpcmpY6rcvyzk
g/2r3UvavqG3/XgSmyLeHw66uVfEKTZw+2PqgVo2BjpHHh7YbMjw+BwmCUD1P9Op
ShLhZKNzyF1b2TMfEs2/ibQDRWMNw1pS44huJmV8amV/wEKD9sCDJ+sFrVC1zoLN
U8fD9IbntDC9uYCJjHT8l9gh1WXfuqW6CuM2WnpQfxJhmtL8ZToraVAyvdyxzje7
+UKdDrZ037BkgpA596M0QVTKt0jfhsJFQp/Z8W7b+zlWtpxHArI0M4DSLE+7SfyH
3O6Pb2U5alC4trATFwt3GUKIyTWR0axBzWwb/BD3TCc/18vlgOKvlSqYUUpNRuoG
SPhttoN+L4ZQfwHKWRDuUdfCcVSXUq2leqL31IcC5O3xmXf5V49ZXmfWf0ssqhEQ
Y9TbwPVC3/j0a9rnm3mYQTVgsQ4J9vfH3a1927pvSiC/qa0sk1SvuMo0xhh5Nh2m
KxvPJM1LikRT4qInmrf6xQEY/WvBs9BwJXRVcovydTLP1ijuMkSNKVcxF5Yyq8Ua
joJqAxSm7Ye98uHF9VG7KvhfoXjzYwne9VY1LmuThGyor9VLf2E77YDo+RhX6lfW
rqKLva+Gh4jrcNqyxy9PrYsJ0LiLwasUvctuFmIFSHwxYSepd3yvUsZpr0dpobaM
9ZcKy8A1C8LOG/vPRXmqMqOaBgwe2zJpmQHQCShOCupXzdI7tnPx/E0FfqeSwVS1
j9caBSDyCX0I5+sV7ARg/XX5g8yb216xMvhoKj14z3o6RrCFaD1xaQZ1cV3jwH9o
cwkpIhXDH+jSL5Gfj2kXyioemcQsnAJ6E98g4krwSShx0dxTHMP5dYXOBCcBVG0P
h8Sarp8BsPUxzr5QRk5EOiFF1Ue8ow/IzTtgUxEhpyEXLN/VB35z/W+t7/MokZmn
cJJo4dS/x19mOIhp+bQWlkkWekLfCTDdFd+SGfVvhVU++rCyufXCRMinNnY7i2Ie
ETREJvxGyY59MMUtH+RKR6C4eY0lAXctSRvZsM9OImbICebRw+4MzDcXZoghAlze
feaVTJ3nu05oIC8yUrqPFgy2TOfdT52ismB+VudjNuaozZejOUpqos8jsO2pxEov
bP/HtRZDsnfZPL71l6YZHlMcfilD4xya3wm4SfosMaXwkvkpiybUZDBdI7tzRc0E
JbWxG92HKBEmhLPeMZ6IGXyTuo8n993C9BQbs+Q71ImkRQEm5XfRfAE/VzInUrIK
PaAcdX2TQ1ZopQB+G1TyWDr2mN0G4D9qpYSjuD5i0tfnQ6yn7g7h1AMFzC5oWTpE
uMfb6JvcYAWSTGQ+pW6RBTR4hgkdC9suQbwIc4JkC3Xxnx9hwaxoj6dM+mUXe3KU
yoe+5n3eCTuqBJWQirPw036jkB/myt4/stBXtxwmhhmFnmcKOseubNnGMcQoOUhg
y12Lz5ur416dA6rLxJRv044MWwvPXf21WUtYOxdbOA6aV0aaEqYr5kZr1dHO8SXm
LC4iKYVPcY+fqDPBI0/i+A2uW9jtLNsTsHb/kRMGx0/RYqUo8JvIft0Ph4qOS1Tr
oboXv52qvb7DG/uzRHVe5mVFAtD2z1LvN/Z5t7NnECsAwpDhAW0ndugUW7YzdP8f
9+Xc6KVjzzpbXdqmdybzG9NxGtTJNDag7TepNdKwwQ4Qd7a/6GuqoSi2T3JMArEk
8l4DV07tgtcjr5VOCSSnfGLHmUEA8Z2GkYuReg6WHstGN5PO6tZf4wNNt7/t6fsL
8A+1QsZYaeaw4KvJQnNh6LBybNCSSrDPhMRaEBZlodsMqj2mkdXI6KZFxPP1RZcb
QN8XhChOP0ERu5ImZ2JSP1inbHAgK60xtV6jy8ORh+dYnV1XaPui6Ifs6aX168+i
FFvu+9djiuBOaMD3p3Z2gbj0b57QfyRHhrtoKE+ltbXkS9dC1U1Fw/0l8a+T26DZ
rlDpTf2EOiY3g7HSrSEITwcyDO5vU2lkKSi7brYENqjbYtdadxheEZYbtrpbAC2z
LDor70tzJ5L61rWKKoqv63/nG+jpCJdnZp/n7mscxyZGZBukltXHb/6u5z0C1/tZ
3+AxDia4aIh3b4CzYPjhrDrILZaShXh7XOg8p5ndC/mrNqj6J9ABId4REvs/zGVi
p0Jsj8Jbj1IBIl+2Sg+VGE8oII8s+WjdJ3werpM2OUigOi+uhWohuvTULdF7PKHp
NGa1cyAFrRLaIpop7tmKJPSDTtVhoKmzHYndAdMbPNPD/truFFP5mOq1W2/GWHLc
MzsBzxAs8f2T+CHhFZ3Hk8AVr4ujnSW5WkqDM12ej+uMO0umTu7Nf364Tl0W+ckY
ojdU9ng+ueFFkLVGYs+igE5GobBVrl5S2TgfJxd2QOZRFY0hJacxuN+VXCX6Re8U
aSA84O5A/IFRIodW+XVD7cGpnZoZgKATUPbHvQTEez4c502dn+psWcgdnDiaaq16
1lO4QF/xkShD2Ot9qioKFSv+FBLZ4uwuyIU28KFe2lLa2Ie7HmrQOAB0pMc/kKmp
WXwJYt3eaCB9knvgYecto2AlQohi9+RN2+yeXSIKDZzjSJDxDPgrul87/yBCO3rE
luz02/dUOweaYgPt0M7f9LvvAoFdIX01U7+0Qj48xuQLLvTLaDJhU3Q84mIVG4cL
VollA3wMbdgxOdHSsLQensKsOf6ZujNyGSttVJVTTTaYwvWMhh6QhcDnFREyVLJg
weN+MonueIe7mzg8cQpL8BAyQ2YF+ZjnDWLFelWse1sp7ElXjv+3xK9Vf7cJ5Nhq
qnBDm3OwrymvE3o5GJ5Ft8fcDWLdOWqICsAdYTCkWg52Fr1WmCs4pUS7rQZkH7bl
NKtxxktCB+WnkNhYeLuetLu2yxPcTdPJ2esk+1/F59jGCtfel1/Np5S2MNoed1UV
d3C44XdnBDFPWgmTL5iipeEQK5pV9hFvi06YM5o1bhxIuDCAk9XZ+KPkFimMb48k
cSeh0XCGyp9udAqNr6ueHhVzKNRr9oNj2/l+WiRwUNl9TLxq2tBAB/uZIsEQ/af1
2l1H8Bn6I5Ji5ws0eHg5ajA5Boy9/fX0tZwHnAQ+yLwcl+PL2jUvyKlrlmKCHVi8
zNllSgdBoqC+L1Q2qvApx2PSeE/gl7yUBxqvf62CVMvsq9UoOEshNXad5F7zOs2y
eB/e9pyogft5cp4ms1GJr6cHQBWrDuHo2vUf2kbZfxZnR0SRptUX4KwnsicZsebm
29Q4+PEUJsx7r8kQQF07SbNmpm5wZxpV1pnKRiqjd67wHBJMfLyXmNYWw9BE5LPi
EgFf2hkr/hjLJrLQA00jviLAzEApq9xlcMfz4cfwlFOdKeSVLPuhdtUyABpmCcCJ
beQ0PTnkk9RYPgb6UW7z+/CQrbiomJJLEToyQiARkMdWigpuTEZZeyrhGOoTorYF
KYv4qeSdD2z3R27gZcP3GSpXt+jplnP5sA4ZzzFqQgrKd9I+lsTqrmq/pcWEWXjF
/0c+LjksCFmIcm1uA02TJeIGi5m+3Fcv/DskZ9CRSiQZ85QluGiES/oJ4l73Z6eG
MAooKue8OsRWiNjDu7kGqPi/o4MvommQdu+zPstNoduWxNTEVn+U05pJ673yD66n
qeBpquF1YdLABk7BQvOU2ynPLxSfXTGWrofV/fJsUcf6YHy27NzR4BPp0BvLjaUb
gjFMw1S2UKuvwjNop8UKJKWQILbmSI3VMGxMuVK0dBc0GoJAnmEPsue5zgxMVMwN
K7MPOCj6MXZKziXL1yo7MAw5L3SW95hT8igYuIEocQOKEr2zQMPFoTduC2OPlNYH
l7Yqk9hi3PUUf0RoAgvAvncd6A0mlmFWD7pHTbsNfMidIlx+Fm5B67cR2nkcsV1V
CIvRTMpp57jsJ6yy8RIvOcIZOxNse75r6SKOwbosxWpX2kptSaBUpfASA+1NdYzy
pzhCe2CHrOF66PvFEAzKFoRiMjL5Gl2LvfJWU4rKSmkwF70uXgBgihkYeor3gTSK
EjoHohxy6sOVtrUWLcjpoxvN2nCLtjC8QJkfh2JHSnuCCszXPliEDGSALE1yusif
ENetUZqD0g+pRfcQH4T3CVxJ1nC1whkZDFkIj8eQbkJSSbv/YrmjzYv2R9HMVHk4
4rW2aFmzWrwWGomv8MuiAHXsK2SSZBYfe7wpY9kOoWrHzvguQ6s2s+BLZ/uH2TF3
p3xZcyqtzn9q8q9qNhJoJODdtZ8aAEXv8ED1LOlvauYG0cpiL0tLXYHD8idNn92e
wdGw73GnFRQ1Nx48IVMw5elScTFzepfJT4fl3oXQIz/+pR+CGr9eLdqi3qDRNvq1
5nN2hkWxvTyKYE40sDxinMKm4BTIfWt7/6nk5QJNGMJMXJ0tJMJK4dOGIVdPHgKv
sNSAam23rRYLbdRZG0ZymtCz8A1ErUyFFDl15iOpbmhZK7aw++Xy8D2iY2344XPg
UKQ0GD1ROVvKa+TqNJ2cHDjsnBggnXY02ZgdAMdBtNtnMtbkW4JFSGAnON17AWOW
BHgjdppZppCFy3Sy8EPQ7tKMCtNCmCaT1WtgF3uRA49EpocfEMWRTBV2t1VpRgYs
KaqYe/8+WUuwJWdLVqAjUWrGFPGH+y2qKz8pUVEwCfIKT7EU+x5UnTs7hcXYupen
EhZo7OgxO7sWd04n4n8egsvQ11vGLOr3HoZt0EW7ugqsye8/UxaREKsTQQg1Obdm
AD5Xv6+f1Y13UYytM0Ubja4UwTk4TZIWmjDrhjPv8NysM6yWL80RXqowjtnSaGiI
gdnj1IgH6z5Om6+N6wblXdcRdMLThqQDxXbbAxJ+2UYR2SMfLoZhxqL3zl1F35jB
WY+zq+Hpl4+svLVhWjbNESxHouopgnzvBerT0tkrVhRiiYlQLStWhxuku/ah1Nsj
i+22XVErL9ib2b795d2yTau8+vQZ+mfVJY42nax7IpGjA7d4CT5GfjcSFxgGWQ0w
gcQA2obUh3DuV4pk608hRZ5z9OClCIRw04lXZMiXJREj51wd1gwBnF2m+WBoSNw6
QuWCGuHpRFp+BEXWW3BcWpuGv2y+HjVJDR/yjA6vTf9Q9yqxdMgrlmHieO7TTj++
DPBtkohvEC39JVmbdi/sWEkMBuGvHXDthUXcMxvLLHEmzA7z3DChsZJgEUBUEPX1
VIO4qTgNOty19xk2pAuEV75WX3xBlxNvrEDnpi1VpB6ic4471ur2bwiDbj6UgOzC
Pzg1TrgSbwCwzp4z8YPOafexHzkMBGgY7xs/M38nLbC94fH9dGz4NRVKr985Gv4U
WffKSWlnHVtR3VUfH8E5NODnXMjlyCQi3NyoBVGBMSq6q6OZOZ1E5Xesi0CdEK4i
Zll2ybA/3lV5zgkndFLa/bn00z6x+6m+ojkNIrxxpqMlheVeAVWX0Hozitna6ds3
LiFm8XoD0bMLZ5E4kjKGRPtU6yYtCozsEmoU095HdJ9xc8hGr5gpq2+QuLhtmNYt
j7vOfvbE5ogIST16AdsWUH+xb1YKcOn/L5LtHLBWG/2B4btYkaecznjYrhPI37wu
EvKDwYwyBTRgqVTllOQZpEppHXUSbjCO/vnvhdCdb/BRnW/MuoB9YU/zgLUsDutM
1TFsMTwzbpSQLqGuiwVuMoLf7JZreeHPZQbV3/e9puVtdEi3tV9FLcp/eK8JjVFj
txkelXIR+NrSBl2YKQEWPcTibQo8adTFTDF1g5zD5L4USIMSEsuYEDerg34tZSPz
/CC39M2TlU552ooaBvung3ptaveGVc0iDQR8s4dwOzeeWVOaR+IVBtD37VCALIL4
WsYklS0gH0ITCBkpOTjRJkHYBcf+Ft2W0aCwUrO51ZDN6FAeNtBQ9Cke5syB1fM0
OdSaxMz1WvLwfo8ZSZ+GbTv/FAlomJTY8TfRVSeKdb/IGXsOErW9aBIPn4FOKqXA
ktS+BkaZzlA3MWh/g0lOtuK2/5xK4lr4zT672cEZ6TEGjTzsct7xqi97RATPDIso
oHXmbjD9eWvKodtz0kwB4t4ppEt9811oAGxu7BOa0B7e0wIzv/nudaT1ixS15+87
6z7j0fcmnRPh0jc2H7oT5GK/KLcWV9hI/2vYyUVJfob9kSHN2BTFMlSOiL+j1+bk
7z270C/dtLJEQvwYsS3wzGbbGdornZnjDmK3uayLHhS6EYDQ8DtgzfgjcMB6s51K
Y3Lgb5FOBy027c7NBayDhoPx6vUSe2brHeegOL1/FdaRBD4p0at8DwmYVduoSBQe
oR0GgoUMK0RQa4SXqnWRJZ20vPGT/egfxvVx8d+fokvj8E1oOkFUAYFAD8xhrX4j
5b3mTPN93xKdXbl9GNrQwUQIcFzUP1fuzCOvH3Bm1TcSq9NJHzE+D8zLOhxj36ZG
KKtWNgTcUyZn5Sx3Oa++0hK9UAmfXynIVuLIsp4EpZ3/m63WhSPnzCny7cJPOF3p
9jDsip0Ia7KWJ5SuOWkYfmUeOPu9vnyMeRk0a5Ey9+feuGldk12mTcThxbInm55M
KVu4Bk5C954/Y+PR2zMfNub6cXqNiSTalOL2DFH9pdDWvPb67kDD42sNY+yDEnKQ
1IARJATIQX27wKsl3kQ7z45Hl+0kULIEn2SBUDkDwrDKXLmtwWc84VLHWCRsLvZI
Re8UbXBCBk7n6mff3HY7otINO2ElAF1Zm8RU6x5sf5XxFlMqor2uA/qnUOAzOKz8
fOH1d69tVuviLZoD6UOXiNL1DhAKdZ/kR2dcx5CtmhSRgJ816w5yLX9+pJUf4Gzx
3XPAOV1PQkVRNNEvw9HMHtfhqROV4lOaj47Uk+DWzbig9PqgFiNwI4mrqWgZ6Gf3
+cNSO0hYuMXMD4K5kTKqWFnW0N1+OmFRlQStKTZj6vp9iLRPyrzoOYF8MeYZlF9h
snao3IcVzxz+LPGq/J1JRoKrZFo/Q6HIFf9DHS4vDnBGo77IkOmmr9J9QrCrRsyy
I1z0+7dpAkBQqbhwNY//cJQBXlL3rVcpWwpoGnbcyFJHJmYSoCBn77oFqVZrMXnr
pHLdbM9yy6XOJ9dH4BN6eVRSxvEHDRTctMHsEHf7KUjmlIKIArIc56c1iDBAV8ck
x9TS63hzbBck1cuvgU/vNxMp1wOKWbpbyUSahtsmPTIHoR+TaxAGdVT5ZzqXIeBY
Ow2A8ljL5oJREWf8FaJFm1Ah4N4IdMXGuMtK1v+ktXqjgzVuo9B+xRaDBOng4vcY
TAV8Pciprpujy6XONdS5HmGIn9gQsyMDCJZbwrINgU0SvgM4qtjBBRv/hO2bo96Y
Bh5o4m3GEd8/6oTtVD3ewDsT3xKu5mg1yLIFVBpmg0supk6EdpDC6SxozmAlmRqu
yBYrMG4cDBgCZd7PP1BqkyxlVxCqSiESoj1GcpF7L+iNvwOY/HlGiL8rsY3/B60y
96ZSeSqxgtziGJGH7BJTFoM8O0q/NdA++gDd3S1yWge1tehoTAqYufxWP1jwUQyt
Zx4ngFD7aYQZJKo50lxP7x+RBMpCo+mykqbV6ZR0gzDeWxG6X8Ik773kUrBKR3VZ
2qJyElRV2BIZ6UVY6SrXTlb1MBqyf5DdX8WLha2nzOg+Vj2GGDGD9pCk/MOjtvGc
6s2GfYkOaCdbEoiCQg4eKKquycmUupDcLgkN9/nroq7bwjo7hFhDP1v8yPWK/wQZ
C6Nw7ZeLGEqsXAafNsnyNxG2aFEpTEC2lkc/Yh0FTRu8wIlgh7UCtrRSK4N5Nju2
TEKeNZ0QXt3C5+ITqWREB4KDHaSHFCaU6vzQ5HaZubyfaYITErh8VSWo8Mov3dP4
VGoWWLjzHNwaQOtXXriMROyxnowkMCVnxmqwFqaIbCBdFTjZclJqsS2JhX7qpe/S
jxq25c9EqKivDbHdwQZSDGjMwtXXAjufJ++zSylWApwXPzuev2xgEDEBXrvKfj/K
e09jC1wSKhb3BnpDzbv2LsI3K8H/B7jfAsILkjd9Mjbce2CIG2ydEa7rAeZZsDF0
IHwLzeLhRZvCyG7pZfbg2Ojw2ABQT1/HuaDT1HdUFbdg+Vg6Ovj62VHFaES5bNti
aVI2SRbT9+T0fSHyO2zaWOskj4RzV5mgeDwh46VT7b1JBB+pYxSK5q81hWr10AY1
bEiFgFkE+nrjtFrFrij4mK67kEtLTTDdoC7djUIiwjybcJ79PNHCMe7I6mQXQXdg
7tXeAj5rpIBnsJ7V8/h6cIVlK6xyV2H3RumzeIw15Cr9pzRLaaN8DSIluVM9KVs5
ZTqKouBOH9/+cpGjBHBwhpzMgVtzluO+VkAzzfHg/9vPSvRz5k/JtbMsgLUg34zk
wHawkZsk0atqLN+ColnQoc2nIxwa9LGIt/clH57NS+oOnIEo4cDW7j9BsA8keaDG
VBJKeKgs6w3YMwypRepSwAoq2q41cCmdBJSQwh/NceiGLVjBTp7vqK8zgZNhssAi
9rwlsmU9X/916EVzOEFEjouuk+nu9FWMS08M1d3GW+rEckuDc/fVrWJR2t7hr1i+
nWAk+tPyOx6xNrWpaiLnMZNHPRuROpL/wwhBlcLNe1310YGeN75cog7aHyA7Afx/
rCnAn8G/Nksse6l3/HgToAA8EhVoSgaPk3UVOP194HfJ2m1iHqnZqkZaY0aoQVtE
+X+YpWdGAKFcMOrKh/5VVqsJ3mHMjFwhese1JaGVx2FQv37u7g6KNvOsTR3Wm5OS
mGOj989NhfEtVSbULkNbBF8fOLJ01mQwMOERdzu5VX7KM1OnAklLhBmTePbgsTA+
vUEGPNHiOoxZ75cwtJ8zF1Y0Yd/ZUWlMNAxDZ3mTGnihZnwVSFsrCw2MApdKEbAV
avScDAaRlwFp1d6O2R2SEaOsNvytWqfl6ZSZpi8/eeSr+S0n6p0nsRxdJgxWXPDN
B8lLJTzgzgmM88HQb2ej0Bvm67byFV3vsVrsRGjs3lstoSTG2hucFfpKpbm2WnRI
TQ+n5ss75PmGtrIHq95ymE0/wMNl0AAtkmTQYJDFSbAZtvdyLYKEDacNIT4zV4cg
GDN0fEr6eMyXdjQPshXNvMpcosvxM/7fCy4IaGeIbWHgMLQUwugJ8JqvYPEZoHpN
+TQEsBj1FG/R230dNLrHNXLvlCktfDx582tp9VXaE9/Rg0/3QEIGRz2GCU92Wez6
YporFv4Crc2ZJYh6l9H+jU0I/4ogD4AJ6FYlA2+Ii587mpgqGXAWTOEftjUdHPwd
yVCRA8CgSy2/Pai55Pt1Xg2hsbdC3dJGKeFZmBmCFv3VAp6PByKr/Uyr2mCV3Oo5
hSdzK0rYqCgKfoJearpjXBLljIBKQDr7IEYVaoQTAQ9I8FcuTtzjVFIyXzHWyhRd
oum6+3W9Mg+Z3Z91vG7LmavC0Nq6BCxKVg1rbEkZxqZj7P1azFGZ+v/qQCBNnBci
/EBbw7UAnhdndI/HWR5Jj+KRtRVVQ1wt0b0kkN0PATFSzy9O0jHcOwLoY+fVNkUP
`pragma protect end_protected
