// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BQKBHz53SDJjBj0gXz1DWx8pMaX5IqmEsl5GjcB84VKJeLbnKwQlafjknXtTCDSv
5SRtjzJcyT95WiAzeYtGEUgoyfBhI3Y4dVvJB8o9IsclhiQRs49zuvm2SWq8oQrH
9p2jDGt/V8NFP8qvvFMYFbJ3wbLTFvLQ7R5BKI6Jano=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18976)
pAAdHcP4mskVxUl0GRZeCV6ckM982zUcyldcQGBMyMiLJw9MCGY0LLwXR6MHOyiM
WGXm9J0qa+yusg5Mmm1M4Z5APEmpwjtvRhHB7FcbGq3l+RSvwMxUTy6M9PXmp4z9
da/Vqsj1UNFISEzTVK/RWkmC4IPYewO4ZThG+NYSFEGjpcZ+1RqXDb9FsWku3oin
j4C4A8n1ecneKE4RLFIK2XXj+6n/ZlIXwcADqttdb+9GrH1Z0a5Ofa9gsn5ojbuY
tpjIsNE9b5/e25HFE3xof8jTU0OmLVvh+bJbyFt/ycwkA0YSu6T2WmK3D7X2vZqo
Vo7i7rYV0N5DZUA5JF58spmNeJgQkBl+kivJFqP2gba7dFO7qnxwo4kGunBTsHdp
w1toyeKq1Ci0TJjI00oss5W3ow7IHBgd7PCp4G77DNOeAO8EaULawa9GaX7E3uGM
QXqTMnLOAYSf02TvfnUHBL5+HsaUXaB16mc1hD/EDphuTFSKeoR94M5B6V/Xt1kv
WKIooc1DhIpCI4RpHYRG5wRN6fheTF2qGMaHm8NGnxlg5DKQNLhACGg4NY9TZAxF
aia6fjaiSBugue6ap5xTNpa2FehmF5Y6G4PYJQ4ZzA+/fLSnOsNheoNFr2VXlUr2
fGf/pRgKrDFzfd/XcmFZElAyG6kJDQ7t+/L1QkxWWmJZdG/sWebWjDS/k1Di6dNz
3k9yd5y+jHHUM7/JmCinlKKAql36Dws56aRo3fQi3JckwD6/DHroxaKzGJhEwtWc
huVnuGVf288BRlP6MsUSwJzmDV3oSjcxX+q1EYLYD7eKceM3PB64nDmSAlndHvdp
Bfy9hetDuicX/qRMvHjQxeJlTXdd985Thn6I+Pu6tawvt64g4bqFxav+uvzSIOpc
jU8kjAaatC5c95+3yHTDCTsywtjLoGP4sYzm4lPFS0cxj9/IH2K58Cwu4kCUVOIK
a48cp36O+8j0CxwsTkOMvwvt4lb9WAAtNIH0pF0554XhFXcapTAwOkEsStW2ohqj
DgNSPLDg1TmL2vIWM8hdHcft5kMqu/Tv1Y8vAG4vEsPZi0Owo3xBGna0QC7XS0nZ
rE9Lsc1mqzzsSv87x09+fc9mGAm/L/PHt+4O+7UkYZpqlHhNPD81pojezQtUEUyn
mnS5rZOrR3snnvLIAcX3gTQyCnYFc6chv5+64IRzrkJzZLVV8xuHl1rWR7RMNjHC
80kNhBjpLmlaiTkJIVSATZexGeN3/S3wgAoCP2NrNzBJcuRUIHuULxJuELZ+lHFM
jDt00T2NeaEmXtcy/f+HgB/nClE5Afw0DxtbJy4FDg8OQOajC/tOfsBEJ4RZrN8q
OY3iPenk0y7FsbBJhkB5B6v3YjOt5Gq6BgI3k3mrplXdwm9MK6Cm5g1JGbmmAFGh
KuFWOIr7PZkURS5INBUis1lgzPs9kPFOjEtj9Ltjcf75jt9+fOaszuwczgy/9GrJ
UAahxcqX0dMpTLtvrxcDImqEx5UOEqAiUkox7O4Q4maB7v2QDkqbWLE4WmzdVszt
q0+AivbLJ+DoTm8jZAW/0JVi8v5/vmo1AIHwmPN2CTK3oBn/BY/L83JfusIdOyl0
VsnvOMWesyXvfdi7ODgJe6Kf8NMBDDJS0cN+ZdN8I7o0kvjr1P2sx8RTilNmoAQ0
0wFdnOB2LItLJ/uuuknIz1v0aiAIYf1gRjXszADEEuEJK9Hh0JMrmxwYelF0mOem
YseAanTrOH/Gz62VGAlW9LKe7Z9cgO8kSjFlo2/uX5oZTejtaVVldVSHEVfgVcMk
fxINli1+b/MrEbU9+irlZeFxzp714zU0JmEi8baMX4qHh7kuemprhCA5LQ5c4eDM
pCthVbd84TrFnGksii5X+sHLeIVHvHmb4F3rZwPNV7Z+H5YJek8pbuPjPnE2+GWo
wfze8n7U5YQJ1QPLTzKoBcSW+S2YWSC2YT1JwquMuyg1U61W/qtjYusHZ3g6fyGj
36SJ+7fRlFRv1dgs+5KuFwzd3pFWd5ZqH/v2b6YNhwoZmkzBG+CgjMSmmkGHUtnd
B19WtVilbHGX9C2GSB7G8hYMvo0obWCSNoK94Zn+YK4cTnwAS8oS98e91iwk6opb
7KoujdHReV4DnaszrWWSPdAAzqINQLFJKhIM41/zybox1QayjA3ICRb6DeIhR7jW
CbLZd0wReVH94vP9zT32pWTDr1hfq+eYEvmqCcP5jjuUX5IVjymAXddPt6Yzm5J9
vLaS6kym+iBeZjFVNCDIN7PQc1xtKHL6jz820giiJBSvkavf0pU2VaoKsyXPl4/c
/EV90nd5IlfzN0m7idwZAP/uNDY/ksfInKn7HEeNNqtSKLdTUGXSkcU7/o6Zfscm
/4JD/H31C2+Snqeg+zYJb6F1e+JoV5CvpKa54P8TqtnmgT0ciZFuZ4AOgz7nM17n
8vS7pVz/aWxRYcsdhMkQqXCgDk7bP5TcYUpJZ+0Zn5pLKC8Zcykr8Et8hqTlBSni
mjnfk7V9EoTkhrf4UUvYBI8yIy/Hc/YnHQnzie6N9LrXSC5cfKh+Z02jokSxR1Lv
6tmXu4TIF1ViBMbOsGhDKUYPVeTb75DibUR2oJVzjeAoiks57yBiEmugl4fJvA7i
njndEHSGv6P1D3KcfyfCXTFqCdmZ1AuACjURpbLFOTh/u8hi/GVQb23mQzW9+Ppa
qQ09hwx1oRTXLMS5hg+oOkaLMu316L5rHK6SbL4fCMvTHUvxNq5k4p7BClSo34yI
n2rqsw+koOCQxtDlmgMx0G8bXj40GLZN6UAeJBWS88h1cQDEH0LtPRCQiAfNs1rJ
MP2VyRg3PnCerJQ4m1LQsZdnhbmyk/9oxzRiDrRcQw66qi8qX6XZ49BE/xi1+xK6
w7fi7ZY6gi9nPxcJN8zkwuHNRHYGP+SJn44WiJ/TAZUQNAhgMeabAAuz5TBj/iEH
kfs1zXRJIa/uds4aK0gWW4ayIQ3uPRpFfomrmv0JvX3UeU52SW2qBITHOvLmFOWP
UAopexkidHImUFZeBURtDKbK8vm9KVtcEUFiEwtOcIonvcjhBzffnqEfQk7EDKR2
IQjeyVFoXWldfsBZ62GbNFGhquY90K4umk6YVjn8b27lTMM26v44a+lN4Dm2/Qpv
jvSYAqwNMHd7Zl5ad9Ujcw0+trwDYAVZiZjQDnhKzd4T1mpj1+cxeuCWVUtFbxSP
wp+7SXMQeykRR46MDhxPvwXzm33erUJuOmbHumqMEEYiS/HQ8V+F7fmbkMythL7w
uWvPIau/Ay13N8h3Sz9WUuddE1JGCZVDYHXeMe1BaLvOjIYlPzT3JfM9Nj8L5KQF
u3ttvyzipk4UGt9HX7XR5qkU+isSu6M0uDfVHYqmJhihYn9ammnlf+oHswVmMied
v8Sh3ob0wtRWAL+v30Q83QS1mU+3WkBPqes5M0q3OoYdR4Bu4diyec87ZLyq8o/6
JkJOykTq7TwvLClpZQ0H4Bm/8cHFIWodm6PgvRskI6oRA9BHW4AYPFKZxTcqiFFw
4zQYF/UibU2TGKTp5kdnK7JXslNWRAlBWgjr0vqz33wcow2zFEQJJv6/2g/TSxxi
dQKgK8X0zYRJJ+Kx2u5QLvNRck83XM3vSyFyNVDeEGAWnx+YbD+FMrMeXI4bD69t
69FJb7z0KEqmH3CHT11zO0uIsoqnbIFn5UdyncQ2M15hNzs6IiRplQ9aZTIKCpyQ
wOnAekIFzW6KloU4VaBfcjlDqgx/OTehXK5OPcVa9HYQSt6rVXhdAFBktWXorvkF
KufO0uLfC7fgCZm2sNglmASe1aBvf6tYnKMAdh12unHrAnDvStNU5KLepwyFQj5Z
LUplLwRxuiYf+RnSVVt5OwyLDDsqUbEIThj/6hP7Bkyd6utJq8Knpdh30tYDIBRt
itC7pkig+mte6/n087yMDgVR9xF+jj6+vdfcmOJjLiG/fg8wsrOxCO+Yrg5I4ty4
IGH2665HYq0m9RETLGiH3Kc3TLo3DB1c6E2fl3HSqnmiRD1JnehvQvNhgm8KAOSu
oeQ4G+WEHIvhCk77bv27PIqQrKT7JzudH5IetWYtacdOlNA8HJK+0zjlCmzWVhuB
+9Y4NryFi8Eu6cR69v+hgymN67yoYrUywM4S7aZqZatjFsdbWQGxytEggGKU/xAO
peZ9MHHeh0owubqpl+MSU97TGbRYhOlL22ptz8Hip4L194SnDmjrWQiIycj73Ab+
Q2AmM4wnn6wzA6B4ZsfvM9v89624+Ux12Yp1MoL9Axif6o1P8YQYU5n0Th1uh6BW
SMWvDbcJxG8OsAh4+cxZEAT12EUB8ynwPaZRXQlT+AX7k2C/NSuBEwgBIVjVAEWg
M4zDq3R/pSYmkdrE05N/Db17tgiGZNqJDnB5Ay8cE2LLUAezzWTLXW6kmnUcqCkl
Do3pf9+e1jitN7M042AkqP5GUB4dg8mIxIYRKHOv44Wp4irxe55qI16z8ZjrXXnF
ngENZyrpNOJ48IjRByr2DUXA6rhy29nChdeehiN8FXmDknDrHtHcAFRTjXJnd38b
0XCC8KRlMzmix0zrDOKGayo6ZlxAEObBW39S1PGg0YBks2cNNWxW9eNiak2nzeCS
dSBvd23nJxJ3+oPCwD93IL4M+rfSAmCKRGQ4OWM6WiMajAPoWOCE0yxSq5BvDfPp
4a1yVdouoM8YsmDyrTrOjvsGBe7SGJCTOx3JwqBjd+sJGSmObETRgjknNpHy+TeX
1uGvA2VzM5UsJIzwysv7MkSVF7egXNxRVfzDbgtnZfseiYMeBsqkK6yFpALARoYc
ysAwIfeUuZJz/7XCIeey4cbtmrQUYRLh4ufIIyMex1FwrMp1WEbH+vzDcb3SRlbS
U27A1EntbxEML/JaCxEsP1r1oU+SpgPJGSGhfWApQUK4rxz0Rv4AruKJE3bfm/8r
P4vqxUKCUmPrubxIYvBIjKlN9Nz0DaPZ+zJggTyAu2BB6U8YNHAcd95otDVtiH8H
L8gj0BW6p9zx3QYV3sX5/Xb7aUmPq9GySP1K7Yh0KgtE/SJLb84TFOlJ2dwEbs+0
gHsFFyPEMTAGiq3ABziMO4d7KOHpGZ9sxWksxsDL1g5TL9ue1spYE7V+nyXQKEJN
lEtEkGEguAEJnh+9KeHXyeCkKdxBX3xTpGByXuxeu9io5KnMUzqMZWcJfCCY+RJK
TusEUf8Tqnu5agEp6JohL2qEeGv0vOO/CVbi5qSoCCafjXLh21GUrZv18uVtISLS
WVOSvYkDi4grulE8qaAXUbxxst3IjhPwE84b/It6Gvmrdi9f97dkHVs+RhiI3kC/
hvPMEbj61SvsqLNCxOl8fpJ/RY7Gu/LX9ugG3XOhhWgW8Q6qgZK+6bWr8HNprev3
zMo8VkGdvruCH2owF0uciIARLKZV09A7ObyF6w7wzUYrUhT36VS4xtVbv3MmKWll
NDWz1x6B9mLLb2DFYDlRSFIXAVdpVbOd8i8bR8dhPBcyMoWQ6SO4MTAbnmH0ruP2
m6JhCG/jWl6cSROveUphPd+JcUeJzMqLvfKttwYFHq3Mo6wCsnugcSpH2pkPPQ9u
TTywHIkyVEk25Z0L533IR1c8bvLW91ervbwBwyoJqd9tgpUBZwjGAbx04CjhA5cD
KoO6X8JLPDk6QIfclklb7OUC4KkPylvNZ4k0PH+hOuAjyJK1NofCiFsALSbhmKFI
scj0LrT5S0ddCVzX+xn0Iw5AAjGmhT2gCSa3jrO0j7TEEVG50Z7VeiplCJKBNkbo
uoQ7BfREl4dVHgPzLMi4zsNJJ9gSQPBBMgBJ4+n93czKasc4XFO2POZ4DG4LdqY8
vqGz1mOV8n396JoF6L0UI6XljN5PapE5i627yp/aHszhOCuvuXIlFkCSmvYYqiNa
WlfMK7mTYT/AJiCSZ+gRYOPdRCNuULoA3dYvdx1PMRGZaUShrQ6zeqaT2hlDMevd
U5bbozEJSscutmc/dyMyC3eCHP+xFyAo8N1uCGG/4oUnHadVE5UfHyGcsW49qvTs
nfUWhCNlNn9NTx6WTsSbzo7T/bMIAGDFSnTsdoWRrjXLEsM+iRCrMWSLVLiwtXpE
ljY36lZL0suDBW9IggLuPOln1EvJjKIfa7TxdgKHUSGxaKVz7bFuDvk2Vpf9gveg
kdd9hpy8BFbbMKjfoN0lu9byDbLdXPAcIK5CxetwDG5NO0Uw5cgJ4XrdwZcY/uT7
iJHe2bRkdOu95yVX2QiUXMn4NEMnrKG6TZTntBYuM3YpkdCy3PTZVcCFKi9xpKrk
MjoSRHbWABtMEEvhx4xr8mCIBB4mGG56pXrf4elFr5KlMRPeocxNRK2UF89NlEQ6
EInCYNq8lBXXiKVc745Hrj+PW2F63JTlRoeZ2l1zYLyfEmvIHw1Uoqjrbv5zwtDe
1m/6eMrXWwvONsfTygjZ2kxGMiIL9v3W8nDHMN2j3/FARQ4zr4QYq+E/yjJsOQ26
4UUxbpDlmA90rG3dxfJ19/+fKHVYDc0fRBHub+MmdUE64PZJLGSXqhScRiLmp6IW
yni7GqFxvNUo0hiHYLVeITC1ceYe+tIHcwBCiUV5xV2czMwpa452NRe/2DvEu1TV
ODpaCGqsbHo6DftEWoa1QhLpnpk3o1YoR/XWpf9S7N1BieALDOCWSkNnLpL16dn7
QnquugJ0tinV/SoWXib/pcmQjvnAmgtQkvfQUkFJ/uoIb0XVyMloDiKQQzHloSk7
RKDNtj8ZI+sPv1bSdDdX/NxtgXUL0pG2+jfhK0dM8j+rgRLbz3bc2+SnWb/lw4YS
/rql2qU7JLvZv4aY0oSSkKF+iRtlbyuw0kspbunt6S+LVED7LpnINeqvuYSlJLvu
fZwItM6KW1CsQDXKEX7uHHMLe9IjWsZhR+SPGTRbRfGUaR2lQyojHtV1osBCr3uF
YdUYQ5wTbXSEzcA+mlTv+8pS1HmMTS8hbUQ50uVVUNKJ1qbW7akN+WA3zID9TiwK
APJzqhJgPGehl6zaj1OrO1N7EKpfTuxItoGlH0ukxox4RuoQSwO2t2nitazD7AJ/
xzWEdtoE/1LhoPcoloorpbaRPgKSuT6rXBFUmXBVNIB0SrTs0h3SZ6B7rfTxvl8H
mUWLzUzv3aDIqYc2ztPyvXIz6EgZOOLc+oadsAgxS+Or6vBrFKeyX78+1CNzwe/W
UNIa2mocCI27hMQvZcx90XcScy0iTWj+CqXDohnSA/V+NiTHb76FY/Foq/7PJ11l
KPsY+13Dpj9GlTBpdN8JtGttKZSYfrkoeqeXW9wA26OcdxY5SkzLoIHgnB7fLI+7
8Id/L6IAS3Bk+lg8SwcohdgGxUxywQRIG+jOaCBL9fY6LTYeaRqJzUSwwu+KXqlf
7W89x9WPfRmPFxBDd2kYCJN9DZOzeD9aAKrw7O/uhUbzs/NPQuzMK6ZoS8ay+m0U
hDVad1kAHUzTQOP9hrmV1b0/bn09lO/QV9bePv+D3mqDyFL7Gb8XxszwCOSM2uQT
KSZFBw4qvGuxsbNES983O6aafY113Q54TWVIhQEPYTj8pGFzcmi1RoJlXG/sm29D
1KN184TUKQdZGVL7avfyisCGPKkWLNankvbbM0caSWiT2Ak0jZT0SeP32TnVcI/Z
GWLlFTLLAYZBQX5Uwo2/40JQj3XF6lwGMccx1gevHZ/A0B32xo+vOkRGxmWszOvq
HNQbLtCHhYNqvz7EGmdZkuYUuU88Q6vj0P4Dkqjc9NRmRQ523uQU24zDNvAVrpTx
oyOVx04ZgGYn4Wg0S69SElEbREJdSn8nRpoIlmmbEI8GCxwgfBHR9xEHZs65zGLp
BHj/pCBSjbtxn9gxLml2wAEjUevOBEKev7QkDXejaute+dwK0yhGpdwt/LcVo2xl
bMRlpLIGKSCK1CQq79cLs0uebRXlsRuEv2minvSpuR1pAeB5tW8Uqu5vpHyZBUNS
Hrjy5ygeVRmW719B8BVoFEK8KbkSdoNIVVQ1uw+bpun9PuvczPSjBdmImKRAViYj
1EOD+2yeMVezjJlxaPK2sjKP1/tYPJqjcU9sRN6RvLeJvC3qJI/GZJjOx8MNrApu
JeeQNmHHMKbLKgEefKMFBUozlumlWv+QYbeIXYFqWgzBfr81rDzDwVWniktp2hji
xC72nzcmWq28ziCh/4ksBxZgD/LJk4P0yghfJ3qmQy2rmP4DXKpnu37i4MP6b/kr
52jsPCmFPhwSAG90PcyEGePLS+ToAhakwH5g1f1H8wCSuKae5doHLE/yZJjmZELk
sCSr5+EHej1X28uCdV3X6/c0onJB5qU7iIwfBICo0xUoICZ/1xVBAIZ1DmW1dhGi
KzSS3mu8Pyyy1SSrUZNfhv7grOlMnP6F/aFDutOOq+/gLhmbnhHAwptdLMllqU+L
j5mFKklKTloWhFf3SURCla6NHokWSQOmMiA9gOR11A2jQDUD8qn5GGFB9qgOzd/z
50oiMrXq6u+rNTUIa9OtTPOhIFA1456ZyrpGEnSUI7XsEb05CO5G1Cdy680onn3k
q7ZTRwcykw8uLrwM0A4BvB0fhYqn06QURHoskVVSKRCCMszbNKS4cQbEj293TN+p
sRycJWRC6FY0Iu2U3AmCrs8wXBCQkfcE6RgX/+5GDuIf3x/SNq/I5+sI1jqLQy6z
sQ0UNfNli004+5CGvqz5l3+0rqAkQD+71R3DDJNFK6Bw5UDQGSorakUX4FcdJ+nI
X5pxd+q2/mcn0qTLsctsb+qEvQzP4SC5PHZU644Ttgn98dMkCmGCyi/fpJPQYF+x
GYRuDOt3vADsFFZAT7jpRkEE6vs74q8+Rb3WqptC4QBnvMe0Y+Bx+O4HdKT7x8Im
Aw3U18UiqNrAISXeyjWG8asnPDYQ19Rz3Kts/yp62CYVywZleDNU5FOD0q6RNhOj
JD1rHP0KtHSU02QfiKdGflyuYW+LjtBBLbzeONp5AVPbGvox27tk96aCIk3b4ycO
Ooc1Qghm/iXbOsAcUU7h4lGIG0ytR8tiM7aHUjsPcRr+sY+UH8PtHwe6AlWIl82C
sFD1kBMNNiLYhMDxlRWAPqOKmABKndlRoU97Ay2zRbyiHPPFyIBv02J0Z52HuXVh
u59oMUcvxRA/hxUeVRRaQAesGXV/yvHET3fMcGL2uF5YxZ3ALXPV6N+W/EW0MTEN
fZzBESE0hVZSEP1UpiO1742mWUCIpyzoQYF43H+efYzW5BYU3VIsoMELjwRYM1Pc
3GOAIuhUJNmC/W0mygmwSFIHFmBDLTB/OzCeXVZjUisqJpldfWWzJWLTwWrCHvHQ
MK/QxffMBrufS/XFXqR7+LXeVhA74aQSCB3rzJCFK+8YIL84f4Gs6I9jlh1ogr2S
+vaKzmJGitcTpSC53ZSsHMJ7Rap7GVN8BaORnmkDb7m/XV5I6mst/GZnzzAwm07A
F4q1xSRkYV32e/OLpfcmoXieJIyjprv7iG6QLOUXGeV80kwZffsHoERF2L2Nt0bp
DJweOWOcHp0+JLIdGwbVAuyxoyLgBFrldnlVl9NxaQlE76PH/FjVNWz3hF0H3mrY
DkOpOc0WnZnju7+Y7QLSi2VCXzvvuGZ74IvXfMWKNd7uNYnkkTMizLUtCadmZaV2
8fN/u6dRfmuhtcPn5mSIViEEvRFj7nWhNiJrxtg0MYMCATG/UaeSQQZpfXuB/vcS
Pm8EiJISe/mvXH8ipPl7QCRF/+49WFF/ONJrtOPk3XEr9Zl5vEU7+AtL01B1csao
RrW6BcqUwaO/Nxzi6P53G1rWv/bqs+RnwYVvRKmbdWlbsYNcFRgjC4rm+bVrigVL
Q2kRhAbVjEcu22qe1qdfKOzqN+qDsV4TCXCZSdTa+cV9oP9EDphcZpPb/DvIfmbH
TmQMoI099zAfyHhfU28hxFdxo3YpktVhbKtxpB4S6MUojZxOhpIvuWZx9vZV4cLs
Z+eCSOVFgVF3Z86Dt+vFb6eC1qh6hEE8QdWviAsx+bcAyeI9ZqgQF+6fsFoX3zWh
Ps+UW9wlil+qXnDTWgaBFYZr4Kv/rgJx3WgyA79s7jK+tq64I/PdoHPv6EcEGizl
oQJeWcE4WIXcrIm0x5r3wh5Ty5Uc2HGRTVaUFgW47Lu1a/ATRBhorUKHE7A9Tt2o
O2yZ7c74edCK/fps+lBwtdrM4r0Pa3WBS7cVWG5YlFdNM0D8IphhgCV5v96qR0Ux
3Ec7kUYaooc4cVFpovg3zcxjYisZA07tk1JMJNNJ6Md8qrVLR+y5Nlgmn4gDTsmT
jPVG5NxridQAWoEulu3aLPDUUQ0h7dMTGLyAElTB1vINJ9ctzeeaHQTIDlIuvjh4
sZ2zjr3j9/aB4JDe3MQ6g2CHuExo7bTG1l4Opz45X1p08UN2n9OrVKIX9JfqFp7J
/JnTkmZ5ZS5DZxWxoYM8moO9RL6vZAg/hN4Av8AmIhV90C4hzHa7N+AcJbZXeFJv
R1KM61HumeQXgZgbJRmIrJtFPJWZBvsc12dg3vysYRbkXhBER1pbKJ8qed+QKACL
v2XrlaiCO/KPSs5GxDJm91SMMnWnHfBQsncwjMOKhiEQpxK2x4k8/DW33e1le+uD
nol++4VrWBn03HQZ6m5KsRS18fYSRx+ofcJfgsvbl1iXr5dEfhMD3YOMdUR//gKX
GGE7YvvUDxUAy1awEAggp3CG2ObmPruk7fChl4y086ZIyYjo5c2QUnUIqs+R6k0D
3076BHForqSBDaI9S17GW0rilueJ2s0aw4NWWCvRchnyamO8ddIvGRroOPhweHhY
GtouQhKlarYG/6sOl2axhp+9b88sqegoS6WPgcTg9IhdkPmM1TSgM82burRi6Nqg
zrwJ1OVOKel/o/qY1CfueO9l0Q21qVRwtCOUyOFQs5+q470CoBa9lq6zhW5GWFtY
dhHzTEjzvQtJA5aTQXfHHh+wV0U86XFwq0xYUskcDw5ZQg7fvr8B5HO5ooCTmU5k
Poax7vvee7jULv182GAO4L8k5TDAsIT8fAZnp1MPek72p4IghRJ/AR6M8/NwJNS/
2ceIItYXjexGudxcnVkRAoPLo6J86OHIYve0WrKrjqEYHfy91Vjq2R7XI8URRy8o
4shLODQ+ty7TCReWwNxe3RDKZQFi3bUZwlJrXSX/BFh5YJF7nU7If1SqkoJF5VPc
JB5mpxfvKgzJ/ruH4lUcDKaT1QXozSrtKy5kkquDpdZB18QpnlO3EpE6mrCHYNE3
mEnYnoEy0b7hkr7s9DZ3bkvB99Zm7UrGD0Yf4hjwhnR/LisGuEZfPJHU3cUUiq+K
sNUUEEVSG1p/KSebbe0dhoF6ckuPj8lK/K3QLVtTA/ikhphri3XgLTNccKQX4dpP
I+7SOmJmb90skaLY8MZv212UuIvgYs3WeBNLQ9YWyGuQa49dnjmqfnHxNwWigU7y
KFK0t5x7VyWLdmCmbYYPGQwIYnnD/ejqcWxaNHCqCBle70GgXWrygTGv4HjqUF8I
FhJ5jd4aSyfaaByA+MkmqW8p6wv84qg+/BBTty/4t7/EOAVGgZZ52CPCFEyDrCls
EjbfimbEC3Z7iUpMK9AzIuKk4utQ909l2d92IbLaQYCCMDBjz5UIZhJjaN9KQG4F
CnGOZlChivVTs6iFF6xy5ElRD69YQFHmFWQQn2KCo0xg1J2lFd8R5EI7D4EP6c+D
6St2+oqxH60w2mMxu5llIJZz87xlaKHCXtxWtpuFi8CKQX8WMKgq5xaHYNPhyEkR
6sp6jFr34yVdy644ICn9Wqn87wc18VS44iynIFcviEdQJrLs1uJic15abf9IVtOL
MazjQesnSkNicvq1kUB61LkSkB3oxhFda1LBNL8jwjR8U3hYTV0FL2ZtprgU5jHx
ZdKO4fqWSpwbe4FpicoK9PD8/Du29fngrEOrXLkTLaMPX2dZXlcmBNszVt6UDKfJ
CjQgR5DXtVbvixjF7ws3cRh+e2O/kVqEhyuidvEAGNVwYsVSvFstYlibcsPvDEJV
QRq+s+G61yWBJ6wuST6TP3m1CfAnvKljWhG6YVz4OoudJnffP293p94c10NvUYd7
vZXCt+HVYegCR/BBmlnB46o1+NspBNMa+lHMsfmCDNSQ3zcURjpuAs1i11VPh1o5
ZS7R355431txcMBIwSwPmxRO20zYvzMekXmhTkfEaKtaS5eSDshdTlp8Dg+qwLB2
Knc8DwpOaiK00j7ZoT8FmMuzeYBSzNDR0Ji98NRbuQTpizd/DcwHK3Aynv+WKw63
uzFzuSXv7FkTGmQsV9DoC9BQJLeVo9LqevNFaF2I/YW/Fr3jBeNufRzRH27qkL81
K0dOTiEqex7V38P21OROhw7ZjcnI1il049X8UL+WfLNF1uFcrjYiW/kgeYBYSZXx
bzQxEvQU21zx7sGaMtFOngO4ulnI4X3WnzlArBgvzM9OoAPVovFM5eq9vMBH+KAg
7KfQIsXm2ezham1q2grfNmqvU00g14ujxfQRY3dBw0WChrcARzBRY4tGVgBsF5Gg
vmBKprlAaLeaoguc75B5IbDKtLn/9tfswPyjncNbxbr4gCwdiUd4d1hC7lEosat4
/wM4joxg+StsRdMKvaNQ8DEHWVHMfHaFHpQJGAPEEaXlGUig/GTaUbjxpbtZXUy1
+DI6tgZyzqNdiyUbFrCkcyVCJktjOh+4SrFD5MtFplzZSrgNzgwc8OBSHRJ5u1Zm
3pMaOaAAr7o9YbhdkWAYzQ+mweyT1tpRFWWBASQojn4Sw9aq7Lx2YFNwsfJno/xj
mjqw99bYuwTiCVzoggfQuQ9iatXcqpJKDUDBQ0Ia5V3xJgq3jXwA+A56N2vGrBwU
iRb6pDWvo7h8UkNta1wO1iO5gJ8i1EF4toHx2lBhX+RL8mFqtA1g4cfF8pP/OcGe
iAE4Sr4cmEjjZEfJlz9a7c1JcSHZLjfUsL8NwrKAIiRncj+S0gXTXCkFgxfLw978
UTWP9z9ooskJxuV3BgW5L1+yx6jVirs3BNAKJnquTD9fEItqFEdUUIQUOJhMUfWG
0bdyiDItc9PdH/ymjyjlvUj2fLgPpBs0OH0QF8Wl7ThqFQSbaQFZmAIfBJhI/SmB
bquk7tZ26eht2QLX9WUhItLSr7ov9qupPwXko8r3N+5CBob66UE3mnz4ziUMRYut
6uZ4/OvOtP1GTNGRn0qh32rBzN/RyL0exTub++1k2y8QHtMFstalpTFF7AApbFtx
44CdBSIsOvtUGSd7eKSMXH7Nkh8T+qDfp8be0u2YQSBXX+/qZmb/ZuFKtMzU4ZTu
bywZ0NITlDjpVvKXleaJIxWgFMtCABehs+zNpXqzMbitQryhvi9URBbG9zuhyM3u
ElGRzD5DUQRu1FEJ3ARpsdfw0B3Mo0I86orDqWf0aCCD9jI2E9WEjQx6GlDjiQaQ
xHtszWpZYAgx5sgg0/HClyVQC8b/cCpl37JAg5Zf8ktrVbeHE0nHuXf2+ac+TOYC
90bMwIDpc4bRl/G81YywQcp7X87ODqUJTStLHjAQLMTre1n3P5eByJs+7CUG7RrB
mxaLo88oNRoJyAXUWU2FOyiq8FxGy8yYlgTaSPvsAI9FSS/uetrmNhgUEOR4UiGT
GKIjo6wbFfljUhJZxY1gEemSeUX/IOuB9pKW5KWzCuH99wjMTWWmGlSHlCrkPDgP
nGvfo0uf4O6ickBuV08NXOEk53AmXh1Nf2IHo05kIPw309QKrsgf0KMEt0RfkxAK
ZJqd/AAe9aW86HQ9TrPn/W54pioNYUOCcT/OS+7ag8tL3yEVwUNcLvFVCDXOS+qb
ELE0gpnSOC2MehMGgjH0l50Hd6VR3qnAll0DnUXLj7Fbi+B1wQVyLR1fx/04dPQs
+2XU1ZBL92thDPbxPKwo42d7v2I4GJzIhBi7eMejfC+UdFu7SQeNebxWCzs1ZSle
n/HC7saDzOr5eTR1OrhBe7346kGzdquRj+NVaRR6iV6MN52rpA3oLjk/WBbLr19u
XRx7lg0YGh65cz5pfvzbGXoDh7jZZ3rltNowtKwXJwCuUTN8NDOvWCIticxyaBtt
8OCKMtXy8p0PqXi4fYO0bPLNDM7KOxZI1ttuDw4Y91L6IjLuGl9FOpSLoLaAgNvL
9WV3xy4JqpAAa0O9YGIhwR9kkIyfCWYQmAg0lDbqW0WR0g3kl0dpO7EqL9xeZH7j
F24mQCEWOXhoVrFGq+fqFPtbCe5kFxJmCDFkkmrF4oGTWL70k3GAfxG/Xibdc/OK
ynNi4W6DnWcljp+SCWaVBaZKvCVMwNSme43Wy/a04CLcJg9hlyMoCyCO253CYvXc
fam8flNQK3i1EL1qz71H9Hm1qLc+hLWDsgTyjluYY1wai30ao8U82n7bL55mIKmW
OM6PZLCgBRSzNy18FiUzCPQ6XVeAyDhSM1hLwvEf5PtQklmBHCDVUDkqegN9T+3Z
gL79NqCMsErB1TaQGd3Z+LhiIC/5SaxnYVkkUxvORq7Zcie566IqucO7KTFB3go0
vdRZu+GsrJbJ6YUuo4SobqhofPPrTKrR7yYvdj2oiKWRF/r/919o/dR9VSRDtBMg
bGbV+vuyQK5Fczf24oCnsrtDwRT6W8GYYurceA1q6zORb8FQUQNR9xunUEpYU51B
Pm0TTGlmP5bJ1bKYakt1rCSz+OMloqegK2Qybbp5nQDZKUpvpn8PiT2re+yB55hP
ak+f6LwIBvgBH+kZQjVs90+G30iUvTN/7kbPbJVWn6WNJeeL+geQeqf5VXzuDq+R
MRdmbIvBPahrPnQZhKaoke29AIwoHc6k9fgW8it+Ly5g+uKrVPwZKgrhSVH4EH3P
S02UaO8u9egVySbP2J9ejhO0PkSc2Kq7yu8rkYDI6CCj//JrMsHusDy/2l9UQj2A
b7nl4PQjrYWU0/iYiSGyXm8VQRIKUf9KuLnlvnKey9wlD8hy6YuExPk0t+PnHDxz
5YioZV3JZymsTwhx4BiJdL74B8R0y6J9MxzBue84AgJdJCUE0rCmZebHGXTehC0l
llQSjfTJDzqA4l9KFHIy+pYsBxN4ZVl92kxIZ9rutog9ykxlwnqq86L1E7nsppCl
KKzFDMFQ2g0YCH7vLnl26TGs/HCgFbtKYAlbTwN15A02ZZtbgioWRz7Q2P2vc0T0
qT6LqHLI4Zeg1kVesr5J5rDvYPo5ShkJKF7uMlbym28/7ZHL/gvpDjGxx2+BdNe1
/O0c4/hU6vTDEHULPgj50ZbYStk8coo4W+XI32k4HgJ64sHw56xFtQatRvL/a64q
jw6NI5wipAYsl1UrJBVu4sb4yLxF4pXNUyN1Q+CSdx39Rnt5oZGDauO1+h41rETh
3JH/SIJGxpLg4ndbZ5fnZ1yT3xrc5gZF42rSq6tuqdWCthQv++PTrGEtnHei8XSH
J/U0GpaaZuu1aY7DuKskGXMuHioWuXcNpXoW+rZPvwlpnvJmEdD/pdXic8DWeiVU
iQBVEnWei+3LHH0wdWumiyABb52J6SwLhD7itbWkAkS7QsCX0aujEPRQ6o4cJZTX
pvmWX+UxwFxMW3Jn0vSxH5Rt75AEDmUk9t2W3WpJaHu5iBPBLW00g4UXqCFTBTML
BDwwrfTmsnHCnMdxHa0TjgmO4bIhLP+deqEvYFF9ASS5siXrrs4Y7d0Z2AkCIEOD
fVZvoZOML2bOl7VCNQ9YIBXjyWdEBxXkyjverK3ZjqJxhIuKNsYEuxnmcKblQX3o
44ZM3/FSnBYxCvwucR5FPjc5FWmGfO0M2RsJ7z0mWkWSXSx/bBe+aofyk4TvM/eS
QqMDb6dXpB+aKOZsyvG7N79MYg9rjQXnQEGR8oLH4kPVFWgiQMz1R5CVociih+Fc
UsWFxbducRdMGJkVgBlM51OGx55yLY+YDi/UyGGkgmQyN3plh8UkWBF/mJgxgrmB
U4ppAePVLcUXTKaZ0lKathI4aXbpm+0JFUyUmh50Je/a6PRKnVGgfPSBo49fJhd1
citN4tRsesCKlojIltX55fad5x0YlsproM5Jab+rqsawy3qPDeWb6S7/BkQYEQZm
NRQo6O/MnHbpOlYbcUq89oAIY3fLMHjmgWuvXKzgJxi50DbBkI2x5PY2oC3FnlAm
AP516xsVft+uqwvOWt2R7hs+cJFf80FgFJgh5bqqcsWSrQM+bmQLxqsTPQxN5Jfa
51tHvSyKP2soClufwXvW8Ahbp5FCct86iwgAQDe5ErgeIdbbzml4GKlIv20iuQ2t
28yO2ulGSreVGtMe7JFlwZjmS9PTiv4ELfEcRVQsdCmo/RPgv/ehx/uk7f8ig5sv
SNtTZofophRTTG1D2HOND9z2Li6ccMkZwiAuU4uDHW4HafiNgxAOuW2K/KR3zBz0
KnlY8oxxMRkynURh04Ts2cnxDzLcxfxy9Xl4XNYmayFjbtxXGFd8KMUD1FynB+9l
qm+hEKrb3h8Vrxtw4edoZp2Y+3QRDu2lHzcuf5/6l/5ZXcRgw2hi1xVUDI4/XBtR
vED8F8fPSFDlohmIVZZTQ/I4HiKfiXZhInGdnpAiVENc+/XLshJTfnL4/b8xISs0
U2XH/APQhg3vC7/3KfD30RVmE1yJQUTAug8SOGuQAc9NKmU3NZ6loCSCL2/duKlN
9pK/2LjYs3p1xuqmBRgTQemTSdKrqxD/GZ4jvFPzqInGf7d8thhrHFPGht91CmaC
sCAycBR/g2E++6Z4c1kU6ve4BPC/+/tdyDR0g/oBnJJ0Chdy/mSSxUMNxVVqPqMG
QElUApdDNszf704muRsSKGxdneZpIbs3qW/RDNCtWEFndNJYrVk/MX28oYHyvnZ8
X0UGzRjKGgu/niqWaHM4ZzTeCxFSBHaHka1P+qhmWYXA2avyZFtHQgDr1M9bcvlm
RBmkWA065bvgTdYJp8RZfx5R/EWBh/3rP6pTbQQe9qFHM4RFjams/KTSiEQieOPF
6laq4GGM9zEZfRBmHx4LgE2e8Sm8TES782aeO05LT5a10GO+o1NgOEEKAyj+zJjU
8TvJZpctp2gNANm9v1tgTZnlLOlxvbp88OcVRyM3iJ8SWcqxDH9Y9Sv123902iSU
G4DgskrLuhsGjE0uvmgZhJMY+ov/lASWmZ9xTkYjvLhGTeX8rtWG2OTvZi0AVmnX
b4YiZnawHP0EwDwAKGVEnDVARZX62G1ROnqHYK82wuiASkAKpXaT4qPzMJ4uw2s2
kFtJ1ez85mkbUW+h17EvpeZ2wP53rsDpkBcXtAqklP/AkiIrXIrIS1PC/lmK4DJ9
Y6WwpXzo126M/mEekm4FVZDivcdenG+wYr6bRREKuPBgSKxts6ChIR8CDASs7pf+
4rHMkDbHUTbNPVG/o8ULbBHFh77lG61giDN5owkPNMLSwgjOK11iNgznnkPyttQl
nXyF/mgTdeHN9RUN2Srj5wsafIFITIfsrfX/M2rJc53dEapgTo4dyR07GcmY+GBc
QWzbZezYq0KTmjGiVVW5TV7AtZcSRcR2JJOLs+Ntm58JKd7S8fr6+rN5lfyZTao3
5Pk+bQDB6gCtKwddw+W7GdHbMpPGJ9b4zpOfUTXXXLZxA7IemAZmeIiUXskcA3TC
iQXtYAzeLmCcHDEp+r0zr0c1JZZbj39Ghgy0maadPFFZdk+N7Mk9Fdn0+brx9jr7
0+veASIDDCDLB1jU1eT1dKmJOdr1sKRL4BHxmqraA3CSBv/Htnl3nNx6f86t/mAG
F4vs1mbAsT1Xm1RmrIn4Q0Fn8LlqXqaALdnwZhZAmlTEdcmypj9YcCz5N3deBcX/
H/r6P3jnUQMba4oFOUOWJe4GZ/9qi6m8Mm32/E5PK8QHgWpw5JZ98j0v/cZFSW1T
sPJ/vlyeEtI2xCJFXgFbwe8d+6f/LUItuE6hKt4aOxZDuLS9hUHGlTuuLfDYD1SE
uk4+29ws1SFFsYbfA01XsDfwRed4g+r8ATxUQVQVBYUtGPQsaBBU88ved2vEXOfF
i8rbSuwwRubOJEvtvBrKXztp0weR8Kk0y6nnJqYukuOQJihk5DDTzQawuOKA5X4D
NQNMY2nkO2i2sKyPbmZ+OxJrndePaMU7hbVOeiP10/nss8vk8DZ0wWIdXvn+VGyE
6Ql6BcPgNeBt3en1jHESkR9Wh22pp6RHrmgWQQK7wUMhq9Bh5i/sYzEL4Pk9xq16
yfUUOQOTG3TpL+5B6PqE6k9ZKmg1iZ7hVHieQUz5lZRt2efB4XjFIYPwMDTDYV3x
z4vMfimQeDiYqCKckXNvN7zJclExYSbkLEdz3wg7PO04Tu4vTWyLDmVu0IvXFoGJ
L9lYIoCf9+VSSjlZU2S7K4tVJaDQYe/A+ZULvBh/TcuLUg9rpCbAURA94yd3I2i6
gizPBpdUiSjHChTJiJVOEMmLE2uVj71gkOJipAQCPoqZ1IpIXSQg/0yG8hRwiK7j
5k5ILU8hdyqI7O4DVGIWn4BoOeTner/x6igKuW0axEo1OORtxZY5/aC9nBwKpqua
e0S9zo932fKZhNZJ7a4J5Mbv/tyL8MHyih7ST4gdxTW0uVWbagiVUdXf1OYIRaPc
5ZVH4wvvHCFFh9QRjwOJsDbX3MUdCr509Pa7yY6VQwPNV7Uai/gIRsynf9mMhfrv
z6RGP3wN+uyLAxaE2ryshUHde/WnoWOCjDDA4/JCfcCwbetNohXT7acOyjZ9jAZZ
Yiz2Sx5xxNPqDb4qcN6PwgFXJmVSi+3RZ/YeZkYbN17Ets4lilhPD/YI+OLvR/Hm
hbyfnYYC/Nyp2r0MpU1uVbumRJVzz9AqQVzzRdg8kuIxE5/D16/z56JwIBGMv+bT
4IF0IZcUNXWAtIVTsJENRu8RlDQBeHKThaxSlDa62ynYqG0q4gBvsN7yPaWIsZS9
7X7LQpzyV0BG3PXAYuNdgq5QsOYAGaKmrPFIBnqOQhIrhFEIC5irSWK8AnOHHD/Z
aqpJpr/XqaGSaV2ZEHjUe3pe6JLqLNKi5kZ5TGiXrmX5g4gHQ8YsxpqiIg6OLrvr
z/fMmSxPV2DnFjT1aYj43bunXHUoDVW8CNNqv3M3XF2tO2W4bstCwzDherAOm4Jn
CY5WAF4+1UBfiQ7Y6kciqgxQHej4swrLnju94QdgFwt6nm6AfyAlIpFjff8WfkfW
/4BxcCsJukBDVtB3jbywXiffTtMfgURKxlQ76JCaXCi1aA6/TKevGpyFmoahnwUD
xUy8sy4ZaazSXFxAW1TWAfKGDXk14fjcnQI0E5Q5abMAMSk/oiMiGzyitDpe8FRp
FfrAXiyM/ZnOrn6ZbLTaw2OFz7LSSJtnJBSPv/NvQTi0MSeJ/xC//vwgJeJC9LZw
mBt7dWGQaavFbXDkBbraprA9FCrsSVSI5TEpXxuYk77785CXD3S7zP9DRCEPXzM3
yR9POjg1rcilNRAlJYNfQ/aXON2FD26k+2ASy4jsaFa5/IV/J2HhyDUtLFuxg5LL
DJ0KAVz2Z9IXhy4PvzXczoUsG6g/9Pis/vZAV01R2RrBIULrMAumLQtS0XAwOqmv
KeAUpM9Fn3gcSVlbfAHN5UZExBirFBar8vmjkfDW0pp1+NUJgHfnlPYJJZd3vHB/
sk91KAOVY50EOr17I+gUOYI9j/mbvMvVpJEK3c/24bZW/llQvOWtLRwQHHuTp2CQ
+qbMvK1/mOMf/jyXVMeSRwBA+24v6Ni7EhBr6YW4iqfWqPIjhW0rz/8xFXL6XtRn
nrgTzx2lVwe7Qvb3o+6lHS0RADwKz6fvAcgglsvwXu1DjBfiwXZ9Glzjs6iEhf0p
/7hmNdR3852VQSf6nK/7Kddqt0w27EGv85SUhujLt7oLLTqLOclP7F6Sukahv6TW
//fX6Mtm9Kv0ECbsH9As+xCF8al5jb5AlxY0WgpF7Hg6AyyYAg0EppYjUm0Im6Fa
3oaIcAyORHoGJHJnnzBcOVzigh10YUohVKcLlExKoxVwra0IxEDabEqVPlaHj7Sl
i2nGWhUkb6qV7oQOlHGucYFxz2Xv9SFCAQLOLtDwowzWF8x+TcTJX8zdLzY+CZub
cJ0TzSLSlFUHpA4GGDcSH1F62RMrequRVCXbg28xCELH1WOalC3oLsE3zKKl4K6h
h6uyr3PrdjrgFGZOI+I127mqfVRqwHM9cr4VJee3wtipDWl/Oi2mqnthvQXCa2a7
FycipB+OCUXNRIHfqm10j8V1DRYP6oUbgmLUNcqjR9faDspifjGoXOVGJeT4cmh1
cMZQ33DjOMgeT4Uk2FuYi9icMkT6vp6v6MaTBRsAROp1wRpa/mO1wxRWbSQGUb9Y
tnfAaqBN5wbqfDvlmEpx1lORqJI/b7Y3hOjVL6eP3jl0c+tsdvRDVwKUVylSSZ/K
JTPWS1PgFcrqyOdhlmIVF+juVEun4epSKhPmFfVtGNJllZkbUpRR/pOHONN34FtL
WAbXEtz9eYR1umVLpDORAsAUEgzGR9dr75n0GE6ARzDESiSjBgHDXt/p5CdJlIvH
psbxGsXLsi4xOPJiSGW1lRNK+uQocyiX00+7k+jT7SomqpeAxp1yFrp6CyJ1j/Pq
COspQnB7rl9KWWQwUBWlStIrqXeCRqdQcjBQg+wgO0CIjLS4Gf7p9m6tDiF1m8GN
fVWYDcIOrv6ycJDPeDP5SL9YSwKBO9SESd9shuurHit3YydyxnSbMqomqtcKu1WB
fLzXfM2fH/ruupVF6Y+JpaCd9IaT6BZfPhlQXT+M3vrKvAB/stUTrZkDcpC99q5Q
X9KZP28UMOD5mCGtSOpu0J3OPdXJSSJtHu/cs2UQVx8K3YAlOLoKRX85Ia2qqzi8
s7SkmSRhLpSXU8av+qY5fhWxHEsVbW8AMlvjAEDtoKUMh60SGjaDLefrIaVHwgP3
ozWWcc5wwrg5mSKRLbzcHKltoSLC8xWkq16AP6s/CLPLK/8R9T57kA9t1pYmCBX8
rIK2ODxTdmUjb79K89xbASe4QttYtQQCNpiKa7sxbzTPC56cw/dctAAlZtzmzVqT
BMUMPdobMb81qcOH7IjDqyp8oTtMm3DTT5IQ+ghIUhJohSvuwCRxeNwdVXHinkJD
yCqVzkvVfepDfaEMaG/uUu3cd2N3LID0HplbSObu66bDnWUk7+bqNMKkQN+Jhx3w
z4TvAUeN8xyTUruV0gBwVmqivPnMAi534Z05dtcdjuC+ccV4pkObqpi3IweB+c1A
lthz+r32MWuXHcc5SnUEp70ZEnaCXIQcfs4oUZLew8OkzwC04oK00ERjx52X/EXv
uFihD5k0y6c7Z5ygqvN4zR2rvKKSKMF9S6L9NigfUT/ptcgVR4jEmK+EJ0+Eg7zS
0doG/pjlFRkg5rwkiIi+oF+kDTTv5G0/tzadbOwThfBqbI807v4JGd/irKgjFI/n
a2hAZnwkyOLOrikOTWYRTC0ff57oRMEeE0bCWT0OdyekQ98hSjbvBxlBJQwTGQkk
Dui09M/yWxoePdduM+ZAg2lm5opH2kC+bZdbsRJ6xPHtp8lDxdgKwfyHmr2wc0dS
piT7+J5XICFHUukvqwjFbAhANASoRljqSsOTUP+AttXpcv+exwNNzV8KeM5pZulK
iRRRqUD9r8WTuHMr3SzySYKe6EXOMA1HK92JwCOCNBF7UWTxBQlT5nDy/8qg7iY3
WnZYTM728Z+hy2Tq5VN+1lnqaF4wrVpRRPbwG6e9gL5MvBKmG1esBtOAJ/ur6v8M
md7C17SvQRBgYxGXMwUmevZbKAHt1HRmtpS1+CX91zixWD2WgQxiExLLRiosVtqb
VZp2+7HvQSMu/+fLTh3My2cR0morwQqOfJnMtiP1RydYItMxH2PHjNRPtBhcXcN4
liWvW++XcLb/KqPn8e0S1/ZUODW+it38O5LxrrTCQgM+wU4CNoAXTKmvphCX59Fm
PeIinKCEduJJH38xaY1YCIMyFbel9MaVd2vFg8r3GMiIXWOVVY/t9uQXoMIes5fC
znDJQ6JlKMUAKddAJ8tpVk5jIsYGHzmsu5/AtXfJvVWZNytzxTa8yU+4qfqy7guu
SloU8TW2kGZZlT0kspuVvpnonxu2KDHRLC5TT4oW4pJMKIOLk0ypVceg3lbOLNFu
d3Phbn5Ayahrd5DxZfPdnqqCJjbNFEnTDLF9jcxZV2cdv3067N9U+50/MLUOnhh1
XXMKqcnJfLnwFFAVqY82sT9aQOyMoSozpE/wovnjE8IRaHrl6Wgu0EXMx1v7Xlyn
+MX1cHME/g8GkU6coOaUbspED62Qe38pydYMjSz5V7pfWia2ErPQ7rsIHLJo2/J5
yElUV8ShqpZhHGOBzq483XUATR7n6Zz1g9BA6Aq/1/ogec7Zc3aU3Nq2vinO+Z9N
iF/2C9bQjTP3IjpojTXXibDRqnAvDZ77XY70Bz9dRrHv5YhNA9gxCUP6m5c1ZOfc
mqH4pjNbY9sC6BBlH47o4A9mXflj52qMmGh9+sRxCDpWWcwa+JeSsIrtoC3ZnVA3
xaPR9qbwGBRz9KOPr4BjGYQh+p92FBZOsPftgZcLPRsC4/UpbnzLTaXcqqSz+hwT
ulWDy93upIyr9osvNfNSYff628WjYxSgq2T5orP1J49jgQDSoNI2/uzMUJaHVKBs
C+PEQal7w+hLQYVNeez+YxiDjQ3SWh+Yky0FPgYde0YQWXKyj2dyEFLDXpQr5aKx
9+ErQ7C9IfAM8+OJSxTP0I8YmriaA/MDgt0t+ELK4gpKMZXZFWUcXf+rhX8Yso+w
cqTNUl2GYSJQoxvdXHIDC1rnUsBTDfUm4tkIz1bCGS5e5ujKMdA573hXp7M6Y3rE
EaCMvyRCz1wgijRurO08aOBUKV9h5/V5fGP+K/ZoBN/EstuaDaZj57GOkiw0Pil7
v1ucT80w/W6zi5nh822uyQqS9iI7VlKYOWhURNKJ8BO3CVNl73bhJwFkmzIF2NB2
3Se1UP/3R3l1upuTSkbsGrRajGLMb1YOsdd9sCq571uJhnPdW8gQM5tO2sLT8ORJ
tEW6ru6d460sB0sOKGAJkpyJM4wLf9dWhM8TbMSGPtcyRU5lhFUsVHM7bvz1v6Iz
LtPMgSChd3QzIoxk6YOjMR0vCK1NEACawljCi7ISHUH4kSlByAKdLpYrYpn/ZJ3v
6jHHkME2c5C+pV7g2bvepBW/0G147cYTGDITyTjJRxcBiIMgvBhwkVH92H+zmlAd
Ld4OpH1cOQK8oVcA/tXf+1SK39WGXPFp0OBBXJ31pDAjXO2RLz2wkkvuiqWVghhN
gGPjm+s6x+3PX+9ZrMZznIwXoqLTlDMXuwlRsENLG0RW+JekLJSmT2ZHKXJ4n/Q5
wR8A9mtnuTJsOUZ3yocG7SorI02/zDwvTd86V+CQgP3MigAIlBFeUthNtd5GZp8B
cOTJvZlXaUDOoAgH3ps9PDI7rc3OuE86RNt2GI89avU9f1DrBWQpJ/OXrhaAyXeD
TvN4xzMelgQX0JW1yWrY8orXbBcNjDqTXzZ5P/JGJp85pZk6ZMI+u2RwQKLDeg79
PGI9Rq+aTsq2VLc9cbFgAwFOr0Z+MXaOenLJ0IWQCdSZOj0mYURzf4UdWSDZ8DZK
zKIWMxPOLwVt6dZt8hassrD9ktzuSBn7OeApe1Z5Sx08rmq8oH4OfhmphcQp6fq5
ZtzFc4p3NhUM6b3aexA9hi0zonK0ef/axXrWhRo2GmfGyIOY8eIyJS/nbSTSf+Ah
Xt/4+BUZelf3ksc2wOsFpWRpo98pSEPn1JP47i2RNJYkpSpKtVf1cQvha4kP0zlp
IcU/gMyOGuHDMCMK+mA4J1bXh9VTfWMGhnTyUCn7/5DFservwLFrlsjWI0RrIxOB
1QvacNMiym9901ishlr/3eYBQ5ePdx0HkdOufebC0SO70bkV6zL8T78AW5pUMBlQ
t0FuCqYRX0iOI3/qlSvsTcf9z5L7V1RNc6/91s2lOIm6da0X5p+wkydiKV9YTvGh
HKCzY1Z3x57SnFv49R3A527oOXwb07EGxOd4/5ibTvOs7oE5l2R2ObGoE9EcHaNz
F80qg/RIUfLocPAvVrYhobM7pzig+GUE2IDlOsV4sv2akKDkg3Uw3rE/0hwxhRVj
e55IyQWGxEPHC+j5CEDkljOQiWkAiB2NfaoT07L2MA+4A+bJEasFP9+CVt5/VWfY
mwFYW3OdvI2R43P9nKwehAdsK0DbUSXVVQo8cGE4Y8j7bp2Jj4OdyuxBwPSbzmO/
JdlzE1WMu1beOHap70a7CXC4jeWCkYV/SmbCH2Ug5uaaLl4pIG10NfbYH+sBEhHo
Om3SfENLZe2p5aCj8V2tN1Xitb646NulSq3+nufoIb8AlrnTNu1xsRjYpyhF6RN8
l7YfUb4fvpD1NOpUN3pAFGIJRtBUeSaVylf7mP9Te6rQC7xynuXUP5d70wdr665i
e+Nv+fN80thw4GNomfDfbwf2yNmG0uQsVKWlDGkCPCEZkB1vgLrXiYcCbFcNYOKT
qaf5GvIUcqisWRPZTqPc3+4BmxQdG07S0HWBRQERa2P9ShP6R5Dypo9HG5B3ISDL
cINrCUnQpymS19r1AriLJu6MFp5jUc0Xkcnanv5teJaFk/AFL5EVWGSiVz8ZlCxk
hVzFSfrEUtWnot9ozh2PX5YcV1Y78R3JKGFZd9GTKTa8PMyujyPVT1WlTe3Px1X1
NDR6hTqZEJdYqeJnd2FL4kEaHjr/CUUubdm7ZuwDUD7HSMNtn2L0l+2xHpa/PIef
k5aVT1sRMIgBvhgRBBOKkFho06GrUbL45O0F+Cm1XsjTpWk6kLxdYwPLflygYdp+
+5K6ZpjF7+9TC6aCZuJ8wKGqypwY0/UnA1sR+AQLR6rctUadcza1vuF6gQ5/sOC5
xbxV9s85M4usR3TWQXWBBnEAILzAgXwUY2BYatmXrRF3h3TWDDwiHixwIV+fxBuu
JOB6XYs5XbhlG5U/GB+S+Zy4F41HAI+YOu4hcI4K7EClqhshj819ITJ4GO5Qqelx
Fs6lH0XnmnfBr45H3y5WIjoGg+XYIANsiBNgpECPac01V08HyLHQ5tT6txP29qN6
NvNmemn0ttjOjgQydijqyoSJsgRYdyG+z0o/Ew5aT4P8UQ1hlORJZp+LpyZdLFY5
Wy2VvQXqT9oelx9cb0/dCbyO1D1X5SWzAFTnB85rWqH7qum0u/omNFcwPL0xIXDv
cPV7YFt3/gUBBjDDG5tY5t1+rmoXzGigyz+TvMPwYKylx9P11F9K15Ay8zTo+4nS
RYBc47NRXLC/7b4nZVmtAsbHW5otKpTX5oHlhk1i6UsaG5jK6OW1GLmQW4vPJ9y1
akazbokdT1xok5JPPFDCqyZ8jKcIi1/Ahvi59p/QsnPKB/7TIOZkTBE9+hTVdDlo
7baebj5Sl+WCQ9W2zhTDcQ==
`pragma protect end_protected
