// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qQUNJQvx26Mko5/ivBIh1t0PpwTZTmLtMP9iECvAMmnNwJ8QUWOf77Mk/0fH1oIO
+HHq+HkG57j6GktUTgBCCtRaomzHqsv4sCt+Ec8qIFJqmK0EG4fEO3RgcUM3/XCx
kSa1/bDC4jx9HotSxlTVLala6n88wF4ShRenYa2R/aw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34896)
hQ8gGNzpnkYvuIlgsA7fGAiXC34KCU+tTcNGCRAGkVZWwJzaOM/jcpV8MbvI03yJ
o7fj6BmqPGaDZLHC5ePO5jOy9OzHRs2mS8eT+be5DQ8Y9jXoz0E9Y8TZzBNXk3S6
2TIliKvSf9TQRR8JXNuTpnwVY3+UjEk0smvsApjLohjeYeAKs2R8eRkj3UZjUARH
fJnh5ypB1otbFUjgyt1QAbGULpY3ptsAMg+K6b9oisLojNOJUZHqh4Brx9XippBD
WCDtK5u8GwwMUybbDfyPa0aI8apUvjsCK8PrnPe6CB3VVPbJqWGEj2AVHzN7YiXC
fKwKtcrL4GcjIdgQRN7e3ZvIc3lsSmUOQUEAI9m61nEcOCCeCMFf2xIt3oCp9THq
6xQGruGU35X2BBGHykmLvBCDWdFvPy39HGyWEwvq2MOzTcM8IdAXgyk9HQOz93de
yyBFXQDkyS6dxQ+5cFoCq+vdDLC5RmNo2kBlOro3PlAYUh28L0VRIPydmPMn1Wgp
4zsGj7g+xOllN2EpjR/XPYTru99p4VTWWtiPofxOONOMG/D17PwviOQqJK/ghbZI
P8LEo1q9hObJ2G4Lm5ORVH67Rl3mR1siuP3qwXT0YJN3QZOu9UfVNzT4Nko3c1kp
OlPb4ifeizPpGdt16yTGF1o2LxCxHkShIy1SlhIH/8alHyMw4y5S6PkVJ0jWRR7p
+OVu53t/m3J+6TT0zPz8iiWioAkbAxC41io5sgnAcWV03DNcmtJ0Zc/aFD/AUC8l
HPY4jhscpotd90kL9T43sCcUQgLB3JuQ9UR+LZ9H4rjEabqu34PYE8ACXAr9jwnm
ozMA5A4HZp+kIv0YE6RaIbmXilvgidEQmQce5l0rpHLHn0J/Jg4sKHE5Mju8QLEL
wnzYFT4DXoGvLv0Sv3DHFXuRRxshpeqHpXwwxsOGdSJ06LTE7/0l5Xz0OPVkumn7
cqkSNGG6R0t4mc9NdjDs+G/Nmn6i8SIG+IVYshnWiAEXvmtwGKaOfyHZqUKHZ8Gh
uGy5fICpoDJmjdWs5Et1j0m1LknQu9GpoJndW+TPdk9WFJReHy9A1YDhPIrRWxIQ
4VfDwKGlvKWg9iHzXVdawIWZOHLzrPulhECw54VIQI3kq0/3jNAF6qq234hcz2JK
1Vo7h0C4gdA3W2ItNfYaLnL+dM3XlkLfX0cnrAMN26UZF+4PmXVh6eMfsa2xkxDF
x06YasS9mA5KmXBcM+ST9saksrBeYcnb/jyb5K5pBKrTFfy2OyFksEyp24ForZ/5
ICc7WHfiSpjhObqr0Dt8XseNf4V13GgS2N6WzonWQovuOebF/36sNh8vf3t/oBb0
hobqRfVk5YLblFjtIaacn2atZMC5Qvv3WLsvgKs2L0G9sc3bkUqzR79HNwwUt8RA
1P5YWzwiKzF7PmINW9I5xBXGiIc3iuEHijKvf5CSuIVCnIIZADoZunElLWFrJhDL
uhAN3AdQM1WOq3EXnnVdfoL5g3vDHwjcUMpXeeNkFCOL62wKGBle0/WewdzvBeTy
w0ZzEb9q9YkBycVzM/kBxdeJuqMChJCe3astwMNQNMBbUkU0/LL68NLjWlDmqGBR
lhlt4btGPGVb6rmq0Hdrba5vonbKpkSt6aEDnDwN6Q2DuCoNieKAfJp4xvaF1hO8
vFfmMlwxKQ8zqDX+WrFLVeWc6kAxxRzsNiZGPJaUkb9KIMKKpvNq82nowHtbgGVX
lvhGUTtsDvot+v1JfPS2+BhZjLfsmsNaMbdnexYGjq1+65ioqkHnnIkt4jLPwm0B
I0hHybIT3fZ4RAT6g9I63IJFKFoA0nWpFz1ADCIyRjNiXds7MGTz5j8gqEpOEFgM
sYLzn+aYyJ0l/4S0p7kunRUsquX0lglah+p8v2RHyyTZWi7uXJGsETsd6vKEVmxz
oy7lOKuPp09SmCDj6TwWKq+OEIUlArC9fumvUtcctvk26+gjU5MVAkEwEFrkzrLp
6JECAtAE6FK8wKkb1jrHNBTnVJC/uKMDaYaXBse7p/HXpDisBiDOXC269USRXC4z
ZrjWTqvfHnEJj1hppw257nzW6NPurFpQi2DZMLfhp9hy7fnGs+nJZcIwccewABu6
6IVX1qB+KbyBihnFThSioZJ4uGHrxQLbiI5Dfa+wEdrrycEedJh0jDWv2UWNACzi
4fz5WeOovfwjr4xD3/sR7CHjXeQAGsE99Lo8tHqCbAuKTDkzko+uC1G6usEK7K0o
Ko3HBg8PbC2WM6ZtUslQGbTiUKC2yaxhaV8OILmKRk2b1EtGZtcNsszx+86xf6VX
uSiUgsCktai9+8p4T7otWC5EOQiiQzNLw/HePZp0wqyt67FM8CKnKZFnfZVRmcU0
2u/1Iz7384rJhHl1xZrmlkvKzP8k9AHh+ahFTK0QOEbM+mMdZEKeis3d8C7SxZ61
AWeDNS0bpCSJgwEJl70qlbnbrGQdbTUMYOlUvFWdg4cyiVYYq2MgBGsP2VL8JFeN
ao5FlmrhQ5EHcKu3oVpeR+NbQQX1aLYxgWK8LPsO9O6Z9fhG9nNerNN4zBNzvxd5
d+UmCx0KVTUr+biaF+Nud6yGvW5nR6fWZHkmURcvo6fnwMg4Xf7I1u3W7/UAOI5d
8KsmECG8CtaL0UaqIIcoc/LRLmnA2hJUk90YGRtEc9kD/fRvabooAdgmiCcmWELL
YI8+21Q7WiEudqAD2zBcvq8YV316gI4IPvu6E9DvSmNWbyeQYjuYMnjZ/EKhtVEF
h5qfgWnaZqL4DT+5RBvijVszXbNfnHbGv6qEa4mVzKkQoQ4cyhP07aQ8xRPXNrgm
szKA0O7S6ODQouMyij07K54yauXqchFAyB7Pq5LCwqE6Ys9t5HS233FMElbRlRZ9
ibUu16qbCSQ2pMAa/WYdO1NWca8r3NSGYEOa2Fxphl8/nw2YP5EX6qFg9S0TdVPG
VEIQH4rJWDnEvaQkWgctTW2+XpsapIBMmAoM5wa3/EFsB8x/AC//Lvt4dHuTz4y/
K15vwpXJ8no6C7eIb0jyLCSeiI6/jx+0vQcQ1l25QfD+Bpi4QKKgXKur5xEExS/o
Rdz/0zrQIuMMWJhv5JW9xUbxyWSh6IyNiI8fzAp/mydgZYQxTSngTVIQ21SXt001
0WR6SSHSt/R9LFOg3+TXozbLbLHfIsQnWxk2lZFfhhyj0SH/Jm67Y+i8+dwAdmNb
/hi6msng2VbNTNErXfiDcrb1YtGlL8FatgZdcgq7nHsvCAWtxIhOmgb2HB4sUUjy
CKiKObc/xp1+4EYvagwCbuovfi7deH1qErpZsm2FgfNk0b2jeEAokwqWNh7wjUsG
l/r7bX7DEeGun/jCczG9Wqk0/2XogpKAVXWpggEKeRnbu19ZSevMZ/kVi5C+9b5k
rYhcD892NdxLywYimPVxVL0grCNui07+ongDWfJc7upqnfN0Quy5sdgdNVHLZqc9
FiP7ye2z0Vgfm3biMh4DOVkMk6GlI9FItF/+62/xLgZUrbS0wEZEJFAfD8fDl+I7
KldgXqA/+bEJT/ffeiq1WQz+Bd8Y/d8OxV637/bh/LFldt6q2Eahhr/F75CVRgP4
nQkUJyrsF2veBCCTgbWny2fHhDHnU5kdLhWs3U42Vt17y08HkIkHDv3yXyyEdPVF
RZqPRYZ+U0KNJQVn9IhobG5CwoPhVeb8gvvjxcdGmDkgnbsP8M6m/EMdx/pQoEdC
ht8690M3szMsrYp+eSH+oUTpb1rXBsiF2RrMuzBqfm3HQhYE/QBsLHdnRxvf6ZZV
2P/xZqLTkqdxxqDumBE9wgOXAZWxuISNgmbnCEMWecuJ/swsqyZpHcdUXFrE7uz+
jAH0Pu1KbeFU2y6iM9wXy2g95uHFbAUyyBZ+ldfJ5cURkbnXaQtElCqH0V3mrZSC
oVZCkrXRlXYNCeqsJgZraXiFYJx1dxOndrSObcM3CEx9g6z3+0CJOf23SD46SKyX
886ifxJTKX3z/aiyVKkOQA07xijRfM5ew2IKcZT4JeOq62OZEYzn0ryn9QA2imp+
avVLUDzE40CcqkKpoteU3tP2NDQ3iC3/aD8NWJIjkOzVaRY4yXYw1BW1T8wX0JNL
NboBy2Rl1Kh2etcEelvaplPolsxr6OD8vkghrygZq6wdW3LbbbvmtAxNvVtSNm7s
uUH1mrm2+KBDrlihBSPPbJHfVpCM7FIFxelsFlER1LqVfj+CxMhbBqKdzCXgNHIr
Pa4sXRxLfxoftD9NhU2nEF3I6IjyZP8yFm185W3pPNybeCHOR9ctMlFpjcbJWr8R
hskCD/8QAa6RuWxB5nxxpz5te28mtViOFk/FlPt8j48pYr9Qo5nT7Bip89MNYJIO
62HcLl8FdIZ6zOWDluE5t9SyCTEqnxS1o7XCIPmOLV9a5S+ro+kCsrGg7XFCXpPU
nq3peyzLCXBzRNNoGoS+kUDXjz7X7Sy5d8O95KAd+aSbJkVV22UKdGCE9KXTsbhN
St6UspM/WZKJFzXiETZpzU9xxfe7+sjTbEQdu4cFV438mS9FRYA8xXT0JTStLO/5
l/yciIM1pK7V/reLpPNtor14AU8QYDPl4eZObLODZk+Pzv1tKu+gR59ZoZsC+fdc
Lw7LgGbEk9JKLH/kR//r7Biw0K6zduoeoK+vo8lk3mNVcYrCsA39Dv6KyyPaaWmq
LKHy7zl+RQ4SjUzrXtomoeMrUL2clZDKS5jocwc5cogQJldJ85AtY1S1t/9X4uf8
Oym9Q5kQ9XVk9FPg+ikgauXN6BR0i8z/bNV0iv3Itw6eoG0oyx08yGE2Dbgi8uAd
vSay/6cigNxfZaDitm/z/SOTw6bM1Z3JDF9mkLruTXCYBVlIdbE2znZR5ZIYP0/G
mEm9ytmP5TO8yowI9SiSLmX1Uv/3UQkX0I3UEiuQhSGiWicWWMXPGKpBVWFKCu8V
WsKW8M85hqpDZTRr/Idkq4ucWBXdktNqmtCcQDtPOiLBiF3yzn+tuZZwhtvUrTYD
CmW7HDJ8E7N5B9tXr33IUUHweBPaRCGOXIaiBPeK0p5qsXxUaQKb0wj30kuuuiGZ
7/iWEIPtgo+lHYAnygG9juJRzMlp/b7VWUdii6udzv2kXwBxqye2ArrH+MzwgSG6
EaatfW77jHncKxZa2ID0B5vt6t4asBm45JW0xQ+jx7STL/sl2GM8K9P34BjqXTFD
XAdQZRcCrKePDfaQLdKolbeWopMVgb0B/z3UmGOOohiN7FX9n5DsviT2PSHojifV
3tcmOTpgZExcWIJJBg0HNPTo17qd0Eg3Xqkh0KDNr46REic3H16QDZayqCzrYmiY
eNv6mjqyC6tlGyrGiHIWcwLrFH9R+9nADgOe0bRRoGgurNmgMnQFfG2JHktSlLnc
8aFHF9qkZHZOixXOeq/E/84d+Jdf46GLW38qUai3XoxHZiwEc9a//ep7bVHZre8n
CLmimiQ3iPKD5W5QkK4JbPcHahl++Vs4iIs/1cjKC3TjJClMZ5bYOs9V6IzHI8eV
l5hykhX2Fw61QKiZLoP62KL7NIdC+HN6Te3PjdgvfoilLL3oqQSH/+on1oSwLDJG
DKl0XuTl8ZqxmgNQBZAMDjtVCmFUKFEzmBzCUlb7SxFrZao1LG6QlRRLKh8y4Mfe
zdHsavr0f87m+mG0GHeE/5s1e7OsEDlSoINXTURnCLaGBhkKDSGwIx4yc/3P7Nd+
GT1N4mQS3e8sZWCgJ7QS3NyE8QpYFhcafO00V9uzV/kqQ8IBBAd5ZRI+f33VvoxL
31VVNT+1tmRE0kClsi906c+Buqb9gVDd313xKi/1McHBpcnJxOQznPpd4Ru4qZj2
yhXNG1iSAXMoppMPa/ONAP3sR53/8/A+/C/7wXEYUz5RkLu1vGUzPOHdCbC6+3w6
jSALqMlv1rk3y7WPzxWKg2RuM+bHPvk2eYlzeyM+kJP1+mhBzTa1m2IWemd0PJr+
tsUNHNhQjnOqB2wypd0Ll3zEpFnT3C0uIZdCIsoZhe1vOB1467g3HzWNtbdGVRxo
WBCEH3nnRbdxK/UvVQE1XRjoSutw9SNRpJ8WvTG6OU+v23aZ3g4YuH3ZDvPm9Qj+
HSHFpILJ6aG2vKiBktTavnU6owsyj779rO2K340vyDHtFuhPvfLvFvXMBby60HqJ
9wfaKwEp5oCqunEbiXOim0EdjCEj6MElXPGR5B8RTOwoVB373n/GWCuIOugvzJ/q
sTOeNLIJuC9XBFrAE55mmOoZGSqFYkwh6Pw4zMJRW/lsrm+JtaVzyI4/FQzLNkLD
Lba65hqoLwM0nck2npvNP/tlN49MiESxK0JDMLVfeQMmxj6H1W5d6mIEqX2ZpYxu
DnYZS7hDVMrlHdxzxnhCCg2YkkDHsBmTCwpas3tK/6b8A1hVK3NuPc3YHB2EivAG
5jPvvozGCJO+GP3zLLZbarVlhsS42LYih5XT4yzP7IFxIyALEZVkhMfZIBeAzn0c
9796aCcLbVmbuootj/rSDC6K/VHmZ6yP9d4NSu2v4BewINPdeWuI4rv2ri5CGVw4
Ve02RcPnpx6PApVO8UlLpVwDqO5ojsuNp49J76DIcEmuYjpPJfS79fNOGwZ3HeFv
EOlvoHwJGQ1xcQyDnuE3fyK6ey091ijqBE0/i/Al/GJXy4pcUeqgfLzgIydvzfSz
Hr+vcbS64uB8ut9Ibs4m/07bqdgI/kswym0bMRn6pQ+sxZ3SC+9+wyj4K5dipKc9
xSx9DRtn9dAe0KsD0uxZvzG7f4sTPa5GqcfHMVWt9X4AOpcOLBqnTTyrlS3e5zLT
NHF1YcQC72mLtPY290AyKzlRfHVtMSvv+Hvo52Yd6RlFZ2+lrw22G+EqAvUzfIzR
gJu4CFVq3Dlyx87QQuiEbFSWp9iLlK3YzQBTw4sZ76iqb3l12qtGc/tDzAfFUife
K7nK1dyQy11JP6nFtrOgoPU8UqAyNurcXVOKPB9XyZoKjMAP0vJFcAYDmcOBpXjY
6pbYTEkQsZ6HOv1EPjE2JwXRmY0+LviwjXay3IUkqHPCeuR6fCj8PrGXmCF/+Lci
IZxcyjjWZmlXDMTh43JPaZJeT3cnfzZfxzncgZeLXhGIxsM5gbNMDsWzYA3bpczO
lkiHlQyIT/BCxruBAwj/m/y0H5LkEdqIlwdlT0tpXDkiVfrzvA9AZfpe/fepTpgi
0UBJJGC/CH1JabL1f/EHUXRDOvLSHofUVqRkAyBGAi22MqlGWfcgPOOoWxx1kPps
K5h7wtbONKfgKTYE86y+XTIXG4mkLXFDIY9k21uWE4lgU0BzUEM9XPUNCKRWkidH
w2b+ynl5DhZ/NbUhs8gJvAg1+9FupXl/Z0AESVZPGYz41VGoFVTMzsnHCY82CaJc
LfB6yg53z26OOAzVna1eUFXMK3BPbHUE9Hxx+9YbegqEIG5zGAawSvoBT+e9tSkF
Fnwga0VKB4+T5gh0+tNxIFZ3xZ2F6QL5/SLRirrY7oQOny2zKu2c69lmu3161O9c
KQbw6evVgko0oeV6J7uX19UGctiiateQnetN8rKCCO/3whSSiM3n0jCU3nZztYem
LpiOPDxq73KGzEnaUmisjlWxrqGW9+IA5XGp2SbNbOwcr63CPNeU5bQZ725c7Gui
cdM5zNVrwF4C2RnObu7QRwBYP5LQcYAs3ir5+or4Zc7Tdzd1FcQUrllrKzaR3s4Z
l3JwRVMtKWZi9aiOHaCWFfPtmwnVDq/B58HAqSBOJhuxjFPklyoHE9wiNOjoFMfo
K4Wfrc1QyPCiL8lnHTS9iftkrN/P/rEyIC0Fd1HiApTPHCDxmajd6JYvQv3FSqn0
PFAJxeXvEl0dF7o3BwIbSbtqWHuSkIF3Wrq6i9c/23lubyMGiPfsBPb/wxp7hIlC
g5psJ049ni8KeX92PplSv4NqTKR/W/muw+Rvm4TA0u2uTfvAwuN//GQLmBY77zzm
fwrMBszCNORjmu2OycMnUQ2g6eRjc8tdvzJcLhe6GRFnFgwDqjB8IIZQTYy3xr0y
ZinyIgcrDCme70JAK0xieZNBRrxztpPM6ETnvp6qr0LrbAe9a+sz0xXmUNqHjgVN
/0JlLEAw+aZvZa8FH/VmIrp5ZZkynVyUqqwRupmVj9XTg+0IAdFFjDU+FeuP5BDb
1AUOtcDdQiUIe+sIE3Q5vbH16SAQTNAZESuHf343iE6MPLx6HlMclv6LkkZs0nV3
PlA3QQY72s4+U5/5Oq0Ud2AQXc6qwXThmpBmt6FG4BycfuKjgmX6Xj0tom+51WX9
pGe+VQDU/cqGkRqmn42UBByJeySd3yUu6VfNLkxKBnbbbelyqSfU5ymkSbNVxHz0
0aordswlRDWx5qvpCbNL/Quz/cTh6gQu4DSXaU4LBQOmLJ8Lf+EwYI5Bxu6eqqaH
d2/ygh4cpxswlZ0542IxRBWFhx09xfzoG2oUq6zVxpVpQ4QKJgqxPVjLIm0X/FJj
4D49s7I7QmcNnVwY7jE8eoRs0EcLKYLCjg504TkWJOziMFHIZyNGWHJbcecSwFif
NWZP3Y2LLBsrXSaT5PZgBOAb4DgF7D7bKg0t+gqRJwtqFd4FRkjDEbiREKKul+il
3U1oOLA84224c30wUuhRq5LLPgFbcz4goPuPosAUWiXctN0jGmin63LRd1NZ8jUu
8QgoLlP8fe/p81mPeubLh8p7KrCmf49+HsrsTkdWs3IWOImTkjJOeMYEPuSxtpWv
B5TqmYnVlsteXUcuGogh2F5O4ICZR9/oGa+I0zJCEGLx7OZPsXQxF/u/yp+FrMgY
lK1oTOrI++WXn+p2kpi27XYP+0JeDk2XBYFSpk6Mdwg0fjnIoqcrBCkRYCu+gO7V
1HiJYkRqN2sHdzR9FhYibPgiwlz+/lQP6kAtBknYA/mfIA64E4ucT+WAKp4P9ivJ
aMw8XvQDi6ePOaln0il7xqZfwkndQYz+aBlAMBy6ZrBj0IeI3X3AIJxYBjeCDKwR
jkGi1Yztro3ZsT4GClDKkEQyituFkviIFM6+l7Zzb0XdJaZo7O18nN/WH+EhvTG4
QaZAHRrfhEG8PW6ZFEon1h6zhJhOEiTrQ9/QU9HYWYG2ZhDaRxsaZfP+qRM/F/4O
McDesCiZEWPY/LcHRp6ioIBeYUXCzKcMFIZaSkpT+kjzWyEfbggdw0pEm09qrHMO
Hv+Mr2qO6G0Zr6jJrOOjaT1LfdGXEFEiyYOt1//91kAj8OGKLHz+cvzaww0yIn+I
1kHqSjRpXD4sohhynlA+p+Eljr3GHyl0Ve72s7t64X8uQIVzH76aWUARs5TOlPmm
vmvzLrtZMqjybZL2aTm97zdr+oZ9pOTIg8mHBCcDRB0aYiyHFLm7ZtfoZX7z28hb
r/0i/+6ptvJS3G6Y6pQhwyNnIDZ9GGxKkRWePqR4Lm4Sc8ERCKfSpmXAHtOoRRMK
c1qG62R2+MUS4j2lo5zLuBIN2aPGsnJuTUhJR5le+83rZ0fZeI9OxXZw9i09ENtt
cUSiMdA0WgACp0X+9flgfIiuNkC01mPDXOzZbEs+nqzPuvGv/gG+57MOA+906oRY
3Dx1zW5IYP41fyRiw99Lq/o6f+Uxvc62vQsf8FAnERVr1bmUkKKuQMBejKoCoNDB
NaTk4pTVvh0K/vLfLoMMj0fZamVxyfB77fIwm9lwAlp9fGgcaHko4mZHlNDZ3f2z
Nzsm0rqQMrGsl5guk9HVL6vUeodbKwCYzUnBs6My6sdV9UaCqxJLa0N20s2uzMqi
py6MWuhjYwVt+TMe+5GoY8nW/RXhuQQzCFpyt62yetFY6QZ6k2DRRYiaFwtSEg6P
aIOdvDU8qhRtlS2gMzwgg8xQzjZalomJQnp0LXW996wO4lTneZqct7aPw5KpaARe
Jh0Lo6pKb8smokz9al008U6oHO35Nri8nAqIrNUeljjWqtAsd1isZjG+aGIoPRe8
mFp364ICIlNpjVk6kwRoxc2moN1YKQQwH+7lEFhyEncnCXrBRX5Jm5uEuOJYsW46
QlvwDaf38dcJDqJHvseZ3UKfJOl7yV47uuVp4yZV/KwRCQxf1g39kU3yxX+Z8qpA
/tWO9JirIyCu1O1ZskEsGUKgwOiEAlsnIwWRoFxDRFYlil8f6e5EjcBxN1CrAXP3
srw6ndSJOdLHfmJXKtJKznaDaVA51HzVKntXZaVXEvkIikhbj6+bwn89C0rt704e
d7wFx082udyiRel6H0RgNsBQAIls9D8RDnImnEF9Eenlw+tYEn+8YRPGtsaD7AKd
n11tkxgSTmHrIKcZhpkpTtf2xBUhOIRVkvf7dmVNB/rwZUq0GyNlHg+Ho0VYUCfA
y2WlvIAHPWNex30vrjDSdSdR/ZOptvVXmBySRMi36388BIduyJj2TP5GiBFqbY6Q
PxIVbXZJdqM1YD62ROaNdgWeCW9qmwZCCByBKQc5qkPkX+NkXPhSjy1vhMzpSUq4
fCsz6ahWnEFeF3hcl8n9xNMajbQd/8f4f7Jyw5A5JsGsTj5iO3TOTiS9knd4nC09
Z+aD3MEebvAJGYa4wfy45DZupIss4le1XkF1rEWQjj4zS+5bpfvcrr/Kim3E2vnE
JFsz5EV+Am9bu/Xoc4AYhJTVEij/nPXnhG8GX3IOIjbnuzLybVFFUHGIGaLklDzD
AxNeG4h7/3zwAuTT6ALjHng3dR4GSZVn5wSIGfLfXuN8a40ntlCaBxoq4BsBpdNU
dj7be/rTCuSMPhTzR8eZbZG6VeYaGholWHB4rNvMxGw7051T1QlOpYJmqLNjKCI9
opMbEbsNJPv/DxniMCcBfZnGQX49WFohLGNeRBLp36lHAQYHgL8ySzTNE+gTbKDj
zuxN3R3YYjTS7hE2/kMn+PmMPvNLzJfGY8eEZn4dAY6Cn+Q2FrtM6ApPsEvNGhL1
7zBLGVlR0VHcaTlvqpD6nb5JmQVFy7LSLqCBLdVy6rdCFecB2inICQsJAEDFMfQR
o3fvmu+Bg7iPTn8Phmk15F7tTppeyKozMjJggOZKN7XWrZ6EaJAn+3DIIDi3XfEt
zs+0+NeXBffwC8QvVBY4qepOaFQyKjx4RfooTTzU46zpccL0TGLhD3fyYH/OT/Fl
GUtx1Uh2omYvOdFpaQAOrs3fstD7zZwD1srbvw7G2TpTUy1eki9C4TtouGAPNhEa
OmK8SFRWEsQUBi/vRCb4QyeUx+DdMK2lByNzRZQBmn5kbSAaHf81DEQUWNnC8cMs
AzmSzc8WBMS4Xe0U+PoTLfY5sh/mGWOYya5K6cJ7eLBhpWEZrjpAYTnFE62s2QVF
/JScLOgAb8PtCBYHFd5f6Ss7MVRJHYDxwfl/VEq8f0qNWNE7N5QoTWhBvEkH8GjP
vXH+52PRJKK5mlSp4h+h9y/GmgdIhhNqmXbzGctT89BSrCKiBYQ5n6b3MfEUN41B
yWayr5NKwj4GuTf+FnnIYMo/H5wFwZ6HSOMdOPHAC1ikkBcaHZ9AeKXnd6sCfOPB
rIrGY4geeF8c7q6w2QytJSvUG4c3dEDw4eYxU3v5q/pcXaK5VY9wrVJESBU1TUfo
f3KGsaOH8FLzNStz1y3wnD2ujTDbtrtnzMQ0zpjoVCmcYkofUXNa4Y8lWcBmabPj
VXIDqDGCEW3ZxbywLWQb5wyLpz5y32BTkE/MQzrk+tllyLH0JVPZ/dzQw7jWMKzg
UPIu7sogy3HzvotmOOI2tOFIzcGbyXgr6An8jozljGOXNlrxGfodhdmsYr25lJ5n
FmeqBtcxIhCiEQP6hD6gVdWDyD25ykspWDOLDzRKYGX+uFqET6Pxa/IlFnUORDZ9
vvs5oaQoBoiajbHtguA5iAZHOLurmb1vvDdj+HI8F3e0A+i9K58XokjZNcnfWjq7
oJ88ww1oRGb0YUcuyqs+W1BCuQRVhteVRHq17ULk3nAhC2v/IY+S1xhWTJiv0U/l
tBVkb+lwhu/NDQf7jT/LGNvg1AzEwYX3VWRJshaPh8Xv8tovWMf+G1a0+XllY1OI
PifVUoaVG9fFnS0Dit8Lk6s/UnVeKIybgXXD4dTUsG98pBBrb7uPl31dbziZP0lw
BTIu07fDba1Ho8V8sLhhwt5a4leiaQHYqaaTzmHNArBqx4tyT6g+jE8ye/6yIZSh
UYSd8DxtZS365uxbLDJsVZDkEKZS+iBdNIubpYm5IkME3bDPGtS/EU1gVUvSfiMp
Xt1qND7OS05G/YSWcmoGDxyvkjD0e7oxY8mcu7dcc1MJ83RVi1LiAqB9n7BLkrAi
ebicIzuL7RZB9sC7KivvKdlHMGyQ4Rx1vGeBpBpF1BF68aGi8jGixR073d5O/ZRE
01EMu3YU2bA0ts1ojvNA5jKT51jRVjjGhcVDF22PPQhtvxrrF6IFnkFQZ4/1EYc9
LWInEqwNRoHsHwUrvj+wuQGDH1S2eezxKkDqdqTftxYfw0Z95/+qw0X2UCEFRvIr
pArMRz5QwWxTOHIzgzZc++EVvGJGO6vjJoGAi13ycuPwpYdR/DyaBkzF8jUJCFa3
WE79HDUUhG45ueCo+3UGfbeUHaKft+a4dWmx/MXYyldD1b6Xi2ZfD2ZUdbz0ZXjx
D8sLpmQBL4XSe4PKKFEE6BVXvnnXDQzMkJNgLYkUYN5qjMu6H2rCSHZ8hE2HY6+x
2g4pTGoJjTjSTkeSu3+PE0I6wx//htGmpV3wUoIIEsQMZAJklLats2M3/KW8Laia
Nua24rwYVfFyOHDtu9pr4hTlYD2S/4bKav7rzZ7wJuDMvtx7IUSbVb1iFsZwDhIg
yYkP5tva+m1B1Kx+EnY2bONOub7QYcx65MbpVcvaGaXjxK/ZV6iMSGI/lv9eMePk
Ahrm26Jf5senykHeW3/Gc7uUFh9xEJxlUr65EceiWtsMbRjaO5xVZCMu7WzJvBb3
80y93V+9TZqxQk/skSWV+9wTnzXyIvS2hQjQJIBjoV0cNHrxDb4Ilet6sN1MC6ct
Ov1hbvTL1wDPuIE0spR3Ij41f6DZeCNqPSWq2b+WlHkFnDx+qNyxdA/PhYa4HnHV
TIOdQJpa4YETMgHb28L1TGInN5Lb03nxIETd81o8wnWJG3eH1MOFkU7WZuK7CNUw
UCF6wGmWquGInL9poJhNFzMIHfGhCfWtHTzkawwhwMjp6qFfFIh+p4d6jx802lb7
9XafPGiyoWzUyyr3V+dGfNi9mlqE20rlfTZfCESSv2l33cczmHpiUNmiIaCrml8+
OkPg6Gi3asjki3LQoYHYMiDzFG1bzg/xc0i2DbkEXn8OpUP2+qa79yaRnA3gXO27
/cY1z+2F2PJQW0R5TiSbR5gkBAia1iW571peSAR8eZFgQJIy2wec9MqfnUwWhvlj
a5mQJSmbNaz9YwKZlsj+YwXtj3pigFZT0WxK4dsIByFIEQQ6Rif5VYvQT/H425VI
3F/sAz949mO6QWZWh3ahCeqWqdfBdqzhnsZnWSgqnmmrj3a8an06F39oYXuoyIXB
tN1Jb394rPtQffSi8+7rbgZXrsjAp/6kmS9aP4AZaWs89/HUnXFplIJuqqLu5KQp
RaAJkSzED1Z3rQTQeZSv1F8agm7Ot7AZfqcA1CpjTvy21cpX1KiiTHNwVF/r5seD
PfR3AsTYHOskdWJAOB034JQ0lfGrrZlTF9AV53J5T0kwr6joaMi5rs8DYWSoOgBW
UmsA4YPmm7yD7JrS1ZoBcQjz72co2VmZwPSYmyOACxbQg3QyJ44jRrBOvX9lh+x+
7Y3rVygyajwm9Vk/sScqQNi87/KrGx9n6mo/UU9fVsU+sbtvi6x4aNnaaTXB0KMs
khhEwBtPbTt0rAtB9KIT9s5MSyjUIhULJ5sB3nU5Pm+ascxRQoex+lO8jhfr1l6a
glbRAGbqtFqbW37PxmOcObN7fnyKz9AjVYEASpV798O282WbCVd+B8yU4D+9PGRH
iVqiZEgxwl9tB7RYe25WcxYmhJg9IQfTBvk62wT7RY2Vz9niBUVjpg4S6SWWFGGl
PmjjNoMsxHELCHg9HjQt8aTktUrzcD4nDOBE0U7D0mx41QH7NuDt+4BxMtbg0DFP
Ll+VAG8hF9YKvGSiD18tIeRtisDAUqQp0HjbvbI8xb2XSZ7XKdZEpaEwpdQUmoqg
tW/Tg+fj/8dO+BTnqaXNqEyEplytqlYdfOWOoxVL+OQVyMSjDEXbuhxHczCWbbgT
pnpw4xZZccDYgu1kpSoYAT5rUsunfdqkciKnaxrX3nC0LqQ6vMfW+80ZTwllFY/g
i2/xOqn74AAm6OBzcFqTbQfFE9HpmmA5UWMy+iG0R0PCusqkguxLDtxwB1P96yXk
nzrBWXYc9CbEyHJmMTR+EG8cAEaI59bvkr48AJTzbAQECoUbuc96R/qF7+QimfYG
fClLr2Rz/rrVe2emcXhkSky6I+qvbMxtFPnuffcUsuJoL8kw2nhnfyk+ECQ7uN1w
iLJ7PuO2mpekaQDmuQhHDZ8afMmkUF4g/BSkXfE7n7Bo4k/4hxqyCjcD0BUQEhmL
cXgDZ+MK579vS6dJe3Tyq59lb5QwE0kt/C1/gAn0iVyqkFWL+lioXBC/mOD/MmKc
0Vz0JFFwYEYkRBm3MRYwz+376+37ZVSIuJp4SlsYvQtAi8oA3GgoggRLBu2ztcFu
/rpAGGHRYDaPiL5Fv31TF/DRylxRoJEbA5qxvanHVvXlYbAzjvrPAcKBTkrWyoU9
o7Qrrq4ebaW7b+L9zIQkFmHI28bJW7NaDd1VuQsNj0YqNdgyc6tvS8PwzQ/v5Iuu
a4CktSIP8EXtnW0PIwc/JGcKlRG5Vgr9pZQCwBMdogW8BO3VEY7WxybIRi7fqmcm
CnEbFzpH7nPcZNNIEnSbS2IcjkpQlQr1H6AX/bwnE3Yb50lrReHFv/FybBoCIlq7
ky+B0alkpvtDb/YBZodcAUGHmMlpFx3nZu0zB3hzhbBdikc/6chqhdnRCzOL2KzX
NY4WDW8B80amZUxsTP/n3MwsQ9sEhD8YsqaJ0QUahtYKRz+Wtf/lKY9ndLgihK26
O6lEcDuC9IYlUGlIWddKgQUmcj8H/8mNoJlsgtMlL3fVFrAbUCf6vXvrQ2nKkXwl
zkHJxzeHheTIAnfQP2esDDeXgq8TC7hJYkfW+lSuvlDUgvDuT0B8zXnSeIavKBAX
zNVXcHuWRnKIBakS4fNfoTXuZNbAKGzOtZoenOyvh6RRrXqMxUWlku4r3IcVgsAs
vSrYPGGlinxSFwo1Sje/XdaHT+vv6p71TdQFTJHEyImCWUp3qgJZWuoZzD9EwffH
GX2msWxbjjNcL3sYRxuDpT79VJVAgeAgmUJyY6Mg9jC8nsuXNQZ54S0NLcCS7ak3
Pvt4VbK7Z/Kd1JHFibi/itxJ0UbW4dTIZ+jVcShNORL45CaT1WMqjeJzebf1nkSy
qGJVpmkakEt5r5QlEBoJLyjHzWi7HAe/mrLY4L8e9LmFy/029dOKmYW+6WBZ0cZD
8OzNSv95GekaBY6LIw+r7pgNF/3VY91esun5JitChbnbBKnMoABhOWtKfYGn+rO1
Z2He0ymVl2/mtGhiTb6munMcSIbDR3nT9HOBojj51dzBZuuVmDWETWo4phsklWlY
OAOk+1uZikTfR4n8aRRpO2c1TaupruFoL5mxP473bXi+cwRbp5ByiTBbkIx5Pv34
xQdkJTTRD1wk4iaNXKkKuVpiWJQSFeCgxsN5fqe5AwmfUkzVSstoE3f8niCFy3zY
rgi1A0bN+9BUDf46gkcHz7hS5OnAzaxd4T18ggz1iUANSiUe1Zbqmk7TITWq70kG
xUVVchjcdJnHQTu2ll6jYjhEX7O2ZP+3YvUZKkZ4NPQGXosxUDC9YnqLTfeBj+tW
BlLQ+z07MD7QHW4EmSeEZTOOWx0s+mtIxObzQRjcAP83GLe2Tp1b76ziv2ZQjltZ
CeUa8pRHPf7JGv81Kggv9PNgpXSWWQbTxfXM8ErwIAUwMk3saAlyVEPpqwnTeiO/
WNcNPq1WYR+fQAeX1aiFtiQJwr1o/aJq4wUpQKOnMuG9N9UROE0lY56LBf6kzt7s
hEUNC7fkCllBc7amAcJW3uB0oeQEUzkUfhTbWO5dQ9/gEoHub7NeIh6eg7AcGa7O
hY+tbHcgWIYu4yTYJ5kdMqcEeXBlRR9n3N2zpiciKHPEo4fnphLlbcqw9x6dDAot
cmjPIxKKUnMR8SyRFSM8JHjeT6j50peptIbcMaU/XRkRbCjw5eNd1f5oAx3l6CM6
l1lKDsimRurpx2NHXZ2qfQ6qMm37DXRkgLV78AiQoqeqdumyZfzjH+sDS3U05h7x
x/QnbC3e0nxW7nw93KoIundV/e0OBVVsVRGbeofipdh7eEcLA7ouk9XJNCPmBecG
DQchF0GXDUc8oMJWPszpYSE5zwG9L7CN2IIZSQBtoYIuDGPQaji7BTnBfkpnDOQQ
/ovLYwCjOew2lg7H5u9Ak9Sqcx4zN+r2igl7NIAsAoaRyU5EZeAD+bD7yxjG8LHj
Bz32H5Ctk3nLdXi8ttETBA2kFX5uX0JC33GgjInZfAS08TeUUPf4xVOkpbJlmpYC
Uae99WUofm7WtpcIt1XZ8dqsPnQS3U8fClGlVOIXT+AhV5qtjm/0MACRikqI72Yf
f5aQdN4jCFXwjEOQd9rxXIBxPOkSb726/uIQDzgKsSduIjcC3c/SyGhxk3k+FGZX
xlDaSOYE7v5exOb7FJejr7hNgNXN6aj/NhDH2y6dmH6SL6Ad2OXnn3M30ildc1hD
/Ex3skEjiyTyrkauxBaun7hhC6+kvFEHrAP6nW336PgECSe628TCVK4ZZM9YEg3X
anbBZfyy6ChsQhDtgoaou3f4c8+6icXQbEYxaJ5VMmUWyXdYnFrJYO9MeiBIOU75
U95v2jUU2Gu35iNs2tzqev0FAN22hJ7KEV+f0HxY1SsnoNLYc1o2BjLCMjsGN+Jt
31jimZ2SEK95t/uwZTlNqHVR5EJvk2o4adiek4WZlOQrgHF8py6EytRAAPTKlaKm
/TnhwkObQ7jfKqpdNNPHKZHNvq1q85UG6UZov2PxbAIYIuaZEHzLNGj7Iy7R2caK
8H7XVjeN5+FlJWNcuTx8e0UH/Kt/YnWSSYdm3ZJmKkqFJgHQH8X+DghABSEiqFie
Ggr6m+D+/WDPCFSxsQKiHvn8Xi2kE4GmH+4K+WvGFMCPKJqlf1/4C3kP3vLaOy22
GOfC7Uil0b0Q7L+dg2hkBt72isufDLySO/+kgqdrZxKwGteC7vbChJ4MwJWYtJeD
ktHSn2VwToylGkHHLFUIMtIBUQaR3RSp5Dvg+GKfk5wnNARhfwyy26ADZSxkPsbc
7iWJa+VI9/lPuOyqipR+Wsc7j7f5dYKS2LWKaayWGvcuXws1nYmugLp3UkXQo3bw
3E5kA9wpf+JnCv7rPrxfZ2PcjqCgHAmckZkKnt4mCiIUM9awmBmnRy7JF7QyDK3R
FAQWJwjgxAfUJF97Td2ugo4EAoFfkkFdgp1SNAY47SrS3YOUa7dkbZ8WY3MdEfO5
czTwTltjsdWX7Cvi7vmG+tDcrOzkVV05yxmmeWwoMv0UVGWNQArFuWF26tiLCX77
PGGSE026h5Wq2KP5IIuJfMqc1DXO8Gf4Q45RRYXur4rzFSXZHUcrtsz2WqHzcABX
zdChd+iBoKRDDY5x8efajCBpSHWLw7/VlXlG3TNUvtV1Ik6kY0oJRr+mX5UUs0+J
WdnVePCIqoKqQ36kkjbLexsmtkXpN6f//DFLOLwub1YaVtU+Xd9vYkIvvaKn+20K
g3OqUuZu/mDxzuVDcri9zNe/owXaeC+l612ijjhk548YNx9KkCfHyNLIa4G5rj+f
18lPP33SOZ4Truuk3KbrNXhLgo5cSHijA6rEC2+mvxotT4YPF8DDTkVqClw8ev6g
yDx7PnvThNGsPOKS2wudQhmZGkBItobgRbOmYIKRXe+s6SJceJhIYL+JzzlLuEF/
9Xzm70cs0LdYfaZyv3uhtdbgLIJLVl+xD4IKABHMHXEqKOaSuxWJbe28IcyPzqB8
dH8U/rJA6Hk4Jq+HAOj/TWiU7X9SNIayHUeSC9XSGDtrggEZlwSz95XzTN8cgN1l
IB4FtB0g3fycJNLcFkJNcVwKSJI2sry6PEoW6tXYKoU+rHcaRDqdmH6GAFD3c0W0
YFoHv2sEZPN9qXLugzAZaH6V/VHg8odJSgAgbdYlGiK1//jSD0wFlD64e5iVIlf4
wA0dG02n206+AGPPqgK+Or5d3esCsZiniQKJnYDSojsGVF2QYQ2SsVujjiSXZYsQ
aVFhy2WFsiz/0Ybb1U7BvlZoxP684WQTxsjECwBxPZTTVwV+GBiemt/LcveNg9GU
/arMp1EhZSnGsaCfKZnMTBfaXPdrdSB00oMlh65a4iXQ45xk4JRvdMzNnJWh5Les
28rbL1L1IDeEXo3U1poxTQVLy8VVUP5MiihOdwrmsZ3UfNq0E1p9BJ3JDWTTx384
zXmpv2PW/34gkZuCVIQccx67F9hNcTFirpbqOc/U9aHHv/mDiSCudW5uvF4TG376
8Q6W6NWfiF3H0KTWb8v1Bj8YJR1qLLlMv50ziqdVK5hfXJQbUS8yO5xVHxmEdsHd
1G3eWsN52kxwT5Gx+qnuXJ/gwY1Gt3gFhKnw0dDFYgFde3als9zqdmJisab7MpLz
owrGMj4dGCZRIgVSh1gNFxIltgQxZKLuW6QGCrKSazjucnj0MeRcdB9XaN+9HDZ2
8d+BhMvjWqkaLK5KlLf90XMqavqtgRzqcwL4mIihiXBHQhsEIIg4qmfiEtI7ogpH
84aKMMJTQGqbPir/TL/rruurzSH060MBXODPd52Ote8ysEDzJos76SQsUuUa0Gt1
bm7s720weOw8W+MIHJoyoQeSeapnJAXw8MbsC9a5OeLzniKLfl6Q/f5bnbvaSdRq
QyH1cMQjKXkGinVolb8b9T4SzOwJy6Xe5awuUixzS106jeUgoiqt704SqJ7eninV
byRQ2H1Ul/yWJ5C0NipXVksKLWGesC6n4GtGCxWAWBdNvvjBlm09DMwPrTUB7dkQ
InFZhR7LdfZ9OZk9QFNQwpTUzICwBPI6tdGDAQtmpP0cBAMxDGnX+3sC5BbB5ppm
4khw352koQju4zGywlIuDeUFqFy7ZhlC3AinHVdQE0yr44jHgrMxkIGJacw6v/YN
nyhWgxsEQz6DQbyitGy1qgApRNRsuYOXD1yjn5l3veTPCEM9eihZI/yqFOtkntZU
/ADNQG8FmZ1V2JEnOnmjDi2ZsdOrAGURWQvDsDHG6HFkX9pcYO4fTDGrCbQ4VktO
D870AhF3pYCcAsuMFHq+upU+fhRipDQIhlN5mc60z7dh4+5ZojeDmcOnznj+Z9pg
8s8Y7gzBuetTakWgDKqNzHrQXqH0teZFv/uTmRpXDidPqgRUqhFq8ALok7ivuQt7
EKUVokebdeVzkR3hQfK3GeGkjjx6cnsOc52/DWZgm40vKqXwhAxqDBiiI4nYtIJu
5tVadU//sK2Px5NG5FK+vJ/TtIOzUsKwnPHHl9f2gMPJOwvaMXWs6th1aE2u7vXD
0TiIdDMwFzwpD4vXOpSjl9r2QdzkcovmezzvlUB7OMQq2NnSO5Y5AbQReWsEstqT
vXiG3/+1ZkNm9rBWu41ntjkYhTo1pt7jlD4R1/BznnbiLrCM0/kr7TL+Ue95YR0c
6qwWSHmwva/fPlQ2+DncODzThKcRd8m1HZ7HCofXgcCOtOsYLkdMD0OFm25XVhzf
aHDHvONWPaBuE7snKpqmPz5bGWg9wfEPXAaBC/xWxck3jgowTSm4vmsJ77A6K07o
mgMYZvGJRC7HnkSLudbCoBvlx4ihsptJTQkrYGZz8/tkCUyUs+uFgLcvxTTDs3eA
zEYcFOO/O9AFbHy6mk03JbtBuJMxVkGkdLCezxZLBg7q5S5EMiG+Vybl8/QiqUmV
nXKxh9YXoVP+Xxv8h3q39iKZRWzfdPFe61TuKdpxb3Hyy65eJNHVq50q55l8Ie28
Isob1v7a8PZtNyUnJMLyh7dEcgkc16f6yHmcYJAuEdhRGorGUCkRNat142tJyCPe
XM3wC9QLsYixGla3NZQG3uW8B8P4pmksqvEVsFdp2N/cjjzmbiAiAfS4J3wVC0LG
nQ2+J1lHpXeNCLU/ePFVPo/j+Gc7Ka7g4nb20apW4uOe5yZ6OZ6zU51rqwUphrFu
LhQV2e6hHz4C0YryYAi6QsLhASmHBVEoq2uY9zkk9IVS8V0Vf+WemhrxcFndISFV
D0URplyHqy4kLngbAEBHjebcPSCElE/GaH3xuZBFRT9naClS4vJf5sLd/tXIjL6G
qye1XKjXIeZbkA/XguQW0HSiYQ3o9WJiGIqEdyP/mRMraFaGdg5F0c5OV0J+L+UD
FrK8/4IgiBuX8oj7wB3WxKHioUE0iujBqUcQYqn8FNhUfR+v9iod96bbbJhzL8Yt
WGmQdpZjQ9gKSSFQJBc1aRSVw9GdKgOOMZwWpHHENw7TSctoQTl+sShV00pUPahq
KoI0nSge+LX8JZkBWu8rRX450/j7yXOd+bQoSuH+NkHTCnZ6BTsL5JtH9STQIK6O
7t08exDoWq431Ksf65tTqKekWfSGtr3OLFUdNNXE985sqEyeeDh1oB2Y8JBnhp3p
SZY1ii1Tx/5jGeJee+pojBI/0qL87fhgDnFSQjxaJ+dd/vyUgtBRdH1skxIJ2H8C
qbvX+Vf0O3ez8WoMikMtl/rCK8D2lT/jDRK2tiYLEwJO3JKcTGf1Yyva9Vev03nk
yXBfSK7raF9DjSVYeKVvL239lgDXFt36HIccC1PSewpjrD8y+i1Mq/3gdqCYjDXG
0SZlhmtKgC1X0Ec1dZAhx8o64Rn0HTb8/Oy0yLDL+Ixsjeo+LMbnyaxvWO0w0ML6
mMKhY8G8LcpvYseZnCrAItU6/px6cbgipd3+GCPRkXB7nN36Hvk+M9MnNd30VDNh
Ici6JnFlyrIQPAC3B9BABwi32Cn6DnfuvcGFSwyeLdEq0gdlVAvoy1TCgu0unkVW
KM43S9u7AQW24o3WXUJbzM5n+LWZC+W+T3zVeH5VBupvpGgNMl3TOvDaCoIPT1d9
QNmjJMrF/BbOKPW6LcN3LVBTKzb3olz8OcCW1DNEhrVhfNQZsQvxB5e7FbAUiLXZ
xfforE0LvzECvAAqgGwPUH4jycl/zabiQq+8JnvDojEszyF0fTF+F85Khf96Rlm6
Rj4C30noRhExMTmL7ivI7n/yUxI8xQ9+bIbmu4t5/QWh5ymCNjSVfcaCANiFUHWL
4WtPeZFHdacNzA5STdlP7UsO17GqpE18vltZBGitq+V0ie52U/WFvstT2ttv4/aR
cRJr7KhWVHUS8YPPmivZwt1SegO7e0wpm0qrUa+8x+YxEayA0EH9tG9LVfheOegh
2J7QHTY2vfzz3b1Jq4N582xAk8e4irb3RRqOLdcZpffsPNI1QEQKGHK3f1pz6hYb
S7SjcYSm9E/q12xgT2kHy2643Wa4dKGdgSOYdazdzxjH5Hqdykfb7qwiWwXSPSAK
CFQYEY1H7kAyxxujYrmwV5IBcA0BMZAqLufNmGDoROJieJJU6BaZndUn0rIGHH3m
tN/ViHQqxceO78Fu03qzQAvqAEwh8SjTiCis0SaYHkfMT99c3wUWwGE6Sd3zjWID
sp8ZE2q2I9s6k5kyY8B3JUXVXa75SVefmN0u4lpqTcwHXxeVw+pS1oWtsqEPYlhn
klOcP0RlT/ge2igL+3xrTv+jQ4XSJErpjWEkRqxonMm94/DthD4u9AliHtDaKQ05
PgkRWjOZpwQ7Kf9iR+c5c4zaNLWWzVzk4HYIHrcUsVVAacko7nv79ZL1Bd0vhb53
b3pYf8fKl0bmuoskw2bonKT+cQVKyxYcKlvRo4NGW/L4Gt9ZyH1VsPlgypedW3dE
vspWILZINmi8oINAfNsI1Cq3PBPcre1K/yWReyb3mwBixb2yQI7BwOLBtoi56dUa
dblMTkc8X4B3dK6deAx56D4az7R9ItoEp1q3prgUh3itM71eZbMDS4zLjLc/RzyK
O0CHV0zhYoKzazUBZm4YmOx4DZcKTgyplgWTSvD9xyskvJWIZhFYC64tRosCJetE
41UDVFNh0H19c0iSRdnvGJbuMdFZetu6y53wOnrCQMy8YZqO+RuNt39H/vXxlAEv
vZ8kX5jeMzkcSkoqf/4dX/dvjz9MIqzqOUTzcgdMbVHiaqg+0VK00CH6q8pkifuU
voxuf832Q7iVk1lLpR5QQl78th3lK+cgffihOegWeE4Q9tcZubcPuBeI9eCXE2hc
mfHIqZdcq4OPRU1d1QglZCiLnZwdGmKUjV1iEso20fP0XrPgjP7QyOawfLpTNHdd
MTgqL4qyi1fR6xs5cOO9LLkIhh1O0UJhmJQ2/te7WbgJwUB3F/IVaAYl/YLFfjXE
9Wsmnf2p+d1pN1E8B8ERicWIdf14wrwreTTSvf96z1y0MPvFmuauGsMlhaUFUYn3
sg7P+AabeLET+zofQzSRTuPTjehxeHns8OMFdnNb9/dBQilgDugOzcmWlmP6VQLC
3WsA79vVhJ75FHxgvJ4ogBCzds39e5XAOLZDi3JvBltk4vGE29FQYj9UubtdsCOY
BiS+8O/lGRXCBVzwae2g9s9da5kqCIVxtgGUV176l+NAEg/+TARlYWe9O80LMAWh
a5nuF2EBF+0Foz5etEy8A4aTaYP49QwKoDlryd0OtfsWdmA5V1/BghIFVkMt0ii1
1hvws5xbQImTPDb86+mRi5b8h104d72iFuxEsrv7fF4WWb99ArbAHj6ruPsEPgG5
HcM+QNvbwArvSbghiwDrsYtyq7DgmviDxOP/i6rDclzwnfF4zGdMr598xXNfqqKu
YCXXC0XbrCi7000Cc2KT10A5PFy6qbekRdX3KmUoRIVOw2ZLOaWGg4/VjLMPoYKR
O1wyaOUO+ttl1wUsZviqwzmKHZVWI9OAM4cOIBqwDqbiLrnHs+XWALK4ixSGJagD
s+e9NF+E7s3tmhyVmuiWC4iMJz4q4UOq7jJQdhGqMChYUGngp8iG1CEqhmIRnUFE
LY8XyMU9yQjp79dXVXqtxSSw+6h1oHZIgS7Ks+r4vGwn+rrp8SH6SFG2DARGed4w
2K5DEsuw2DVx3al/9sUbv+xKjDAw++zcxb5vt2RSWFPMGVlGqnf9Osjs4uYJoHCC
6FGV9WkI5Jgq0zUlufv1/r55RbxR6k/cr+RbdMGvVWu2h+VgGhc4euRCgCx5MrfI
7XZq4yihXGaLFYtlyVvdgt9sobw88XqSojhIFxb37YhtDQJIgEp4DIQ3b7lCiWir
0tW8x6qkwtiu4tRbIAv1tzIM5IMGQYAVl2DuA1i2Cns+U4Wi9f4yCZEQyhwGeXXo
1j+31Ghtz3MdUu1NWkTnn5ag1E4yrgJkWkIrRp0/3VkIeVGRxqZBix6QO+ZZM3Fa
lxqSyzXwmneYMiypQLtelUTLnBmOdoVG2LvIR00D7woeHqweFKuV3nVvJGZ9GJhv
rxco95kBigKfq8cfQUdLjgLIfRXRrLKHCkXM+x5YaVN0ADMzWPwAETtB6wvVA1fc
0K4hNJO2cZ8XxGaNIBqUIT1yQ06VKcpWcHfl5IG7eMA76Ayi48qF768PrjyKOt7Y
HtMmhRb2rf0Zr5NlFfdyfXuNL9NqKxX3y5oeanutfCMgGHds0reoMD5ztb7p9ep7
KI8jl71rfuF+RqaKXo9P+hgxbkdLO23ZagCpttPp3COGlOwzLMZd4qBTiLpb86dG
A3oqygO255+Lgtl3I5MgNmVhxkVzHhnO9fPtgvYD040udhMN3THO9oEW/jZZ9TWS
fAtIaUenz8ff9l9G0ter+voO14dwbt7/YT5gOoltE7hpW6DuYJwZjSsWBR66VFZl
viMd3NzJ2e/pzErE0CsMnS3lLwG3M1KtVU7LzRMWZPPzh2us5NXMyqX8q5DyGkSV
5PzfPygzMzpGom0oEFOqe7g5RoUjEP0epxiGvGGa7i1MgRzV3VBAr2Nap1q+Xz+J
k+9L+it6mMXnsX57ueQGYlVxzIlmPXPWkd4UFXPdOATsWH/TiIn9uygU42YEC2kR
V8ayZ3V6hs/pwqt6KdLRtCLwpvBV47Lm+XmDsbZOxzimxSy814wHw+IAIHnsr7ID
C6p3kqPy3eTmvLknVC31u7MfgZMXamqTgEvUhB83AbDqrb0kI0wK4qPBJn5JPtUk
B8MDectlk1TZZkZekALmjmVdsYBESUZ0RQrSBqQUtRLKJorcCPERZvlz0nkOxiAi
9R0RCW1FRoYbKlIREb9YtJgPg78n5Fz9HguLEmAAWY4aQgH72srJ7455iZ9JfFhs
9oH1o4nHPJ6xTOzojGJ4TNaP8C2ggsujUsSfgKPB1vkvqGBSWmLo98uBy9pF+tOB
nAkoCBqKNjUFAuEwOlUnrgfrnvCe7O+gDmyu4Jxam/NSDz8y4g7NBczex8ymv433
jRVaVBGbSEiJc0FDA8hXOy5U0FbCwhhkll0LcWcFbfce+ct9tA6uaZFUEpMBxC3n
Gn7EcwxOqSCdK/DOPDuszu1su0eYxBI4vQBlE6canc0Ef9ntelEWVNNzApUiiPUA
hpQuOTfBBEMnMHl43+H5tX0FtZDmC4qiZi8BGVMzmSqwfMw4fUYz10xPOhblK/2G
q/nnUODIjYbTcz9y2t1m7V/CI0pwFE9X/Uu4Koyi95OlygdLoDz5YFceAh41c6R2
H2OPyaXvd5ZJt6ap5+hp37YUYLJy3DZcXVT04xNjckWeJE+QLk3PSSFk47VKMIzK
BNkK1UMlmw256lTlakdWbmb+huRpy6PMtSiRL5uLYoGqpMC9D4PsianIbYHTShfq
26a8c2h/AkBBe+IXKkSvNBQ17j+ZM5wQAy61d6mOwHFwnKds6F1St60uxaXM5ajG
AyAAcmM2UEELRR/Q6ky7Y+oP6OVpm02Tfe4lhhxtnhW4LBCGokQ41mNh+GLehSQA
/fUu8owu74p4G4eFpEBGNTFcKtDGJgBqjykzINYArrg1wV+pTZm9466CQQPvT1sz
v2/QNWTg8HjTw7fQoPvFb/G+in/h4x9oa565CkogENbaCPHqOkOZmuKNBMPJDm9Y
xaIWNOnCUcRug4jNjbqRmwkiAUY1160fw1eZa36lcihTHEfFauVQ1GDUHqnJBlLl
V8G/xk///G+KCPL+sufArX34PG6DzwugmmJ/3iud9aKMZVXw9rsuJVMNdwQa8JGS
gpdf4nagJfXDW7AH3gY39LGEo2qO7XaJ3Z26d+7/OaxBi7jy9uUWnhW0d6wqwaM3
bAX+2Na1/z66CAh9UekHBi4icmlqOcqs2NEmLBaCVlk8gRFvilaz4KNeZKMpWG/7
Rxq88qtWU8eLL2KBbjAUQYLyDA1auu2/+ZlaMR74kECUi53yw6EhyQcMtNH/hkNh
gwCnbVgcqcQDs+s/qh0V4aV1W7Uh4cvE4B/QoS4JV+nMnbBNVWbSJ043Dw7Mjkhs
PpUqnf1pWEIbr/C8Un46j4waa062we0JBdhwika0co/Auy8fNIa7FZrJ0Wo7aCrI
5h0dtsCPnULZhdUFfrpiSjYLarVScSEI72axmciyZ1y/IwSAW97x4h2sZSD+yEs0
3VUjyipfYfGJb2xtpjdOzeIFSy82errjf2xmRy0hi48rJzkMwbNR+AE5UKhoo2r1
YH+qM8lMlDkmpx+omQue+95iGx9Nzwo5LgDLa7NTyrwTYMs/auzlNhi2HBnyXEXg
UI6cB7COL+DInM4K0+KL3aJVq/r2QBfr1sLese+ecseHHK/FsCiZ/Hzl+QyPNn6H
cc2zQ9O5yChXcM1lXhNARuernD0+sAhXqG/SHDKo3nJhWaxoFU8X11VRV+pHxv+g
mIu97FvooL5tSn029wx11BuVun5VBpvvV70wCyTnvkmSqw4o+xFkQ9pZxAzG62Zm
D+XkgHf88mn0wFlXHa+vDitpipw22d9ILJsrPzK6LcFU3Uj6rHkLhNm8dwyP8+lj
4rcP2wp07naxgYjMKz5uPc3EmD5iQvRQhDYS0QyYruIUZBQdgRDu+fxzaP+SHGGS
mxaxnJUfLk4/6Oy7ycKIGl2bAB7u/vWHMUYNG5+vuqatr0nG9GRK+tl56g8OWZqK
bG3Lryj6YVvP1bteJd3hnE2NFhOI0cRU1YhqbdbtvpBEtYa3lg+TMccyj2pjBUBu
95cth80Xfs/4LIGGwAG9emGCpzMRocGDM6peNJNkidt4/ri2QO6zClGBnp6H/pOu
LX0kVE3HbEQBeNTpYwTEWW/VpC9uyin+4Ialh2gkYUb+sE7t11sy0nDJwKeAjz0j
GyVZK/sL/WzkuM/HWlMngl+CN+UwfyBPr+ihGqYkRRJ1/C228NptlHnqv96+kLoP
J5tRtpiER9wvTZKRRJ6ijNEF4atsGogagop7I4L2y1R9EW08s87iihnnNVgnkLrk
8dnDSffo6mOOFQc/dpWok3sj0VxW8vjMLQfQc/sIuNqc8+UBoQu6RG4LX9wxT2NR
hBFNe4wzGYv6vOEQPJK6k/YAnOQLpifgRnRp1PILPyz95OKS8WYAc/HgqQdf4QEQ
PMudt/u4RDc5i1CGwSWmvPMDFQRbz3wF+76KXXCtKQWbBCiSMDr1q7N9V+Cli33u
KS/KMkfCssIYDDc3e2cC2znO6Ubd+gF3U3WxCDWvePGZhybdsJYpfZXM2/R+qEbm
f1BqkmjOtLnfXM9mLhew6UxzjVI6cvEjfF8T77whVyveHSwKLjogLiiNXqXP4fRb
rkr1bVKH8sawzLCBZYOCMKnF9dgRyjlBqVqlRtZO27nOARJbmopUHZ6ovIHCya1t
ykagUX0oMImrbSLQmYdotWhYVtp5ygtd5bSXWjNhcJQp9Xn7LlgVs6TcU80TaszK
XMzPcCjf4jXA0dUmEVwQtGN0EBZ7ltIhjff1T7edzLWHVWKW6vwBC883Oy9mXV/O
BulpaSOUVQIx5j5rijYoxgiJpc5o8DE6bCc84jyjbuhmIWoES1ql4S9CpMQ9NQKF
imNTeD47G+vvzgJJNiPQsIZeaFKCLNKedzScPn8pLIU7w867YEBec4yP5J/d6krc
/fDbEEZ856jGdEkuIaesT0eiSYNiqwBQczQngc8FMiuLBAeeRWCc1lPQ6r3FOwLu
SlQN6xuAcupDVO1uGrwdXh0uafY1tqTl6ACcxbyj5jTWPxMVDTVEE1vnVZrtZM08
lME3X5IIUjLeWCH5CU7gxXhBlAXMG8cB1nG/ZjwNpgvwFLAU+zZXyyAVFV3F4UDM
rAjxBjcCKGDBOPsPByY8OfzKxmEAVL8qdeTD5xjd9E5+brvbvG2Oyb8qTRD/SOQr
YVeWzgJk9KV0PVkHyLwXzRqGN82Vvfy0ae25eTq26MhH0eAWqMa50DY9WtV2fas6
sVBxJv1oqXmOxazS01CsYP7eIQQvdxxuJYSRYn0YDB/EGm/0X9yEb8FMxPygXU9d
Qucv99jlgNnekL8Qtdf2mf2AvgGkC5YUih0QuaWsFFiUNWcbU9pDaeVtpXtrM7zL
0vMCv8hiBpdGMgfZMlVfOFNkcJthh9cYx0Wrgojze65yNlHTKfh0pnf7vaaPuIdW
xu5yHdW+t6Ct46KMuL5Yn8Y9rmrx7oaXwYEzpXqDOJ8/yr1xCM1K8KW4l86O9BpB
vm6S23UDH5I8vScFdYsyIqUlyTePgGT7z6X+TuqqePz3wxmpTZSjGax92V/IAPwd
Ii82ZDA4VArzhON+yyjjEotz6zmNug+xXRXl/xD5IHzdRr52g4nxTGvHcH0lVSWC
/LTGzPb+OUd7Zf+5OJ3lFD/ATssQ6g3Q74DfO7JIjPL8gM/BowH7l+ufbboD5tEm
+hV/jLmJmAGrSkCBF4uGpbEJiyAbhcENoePLtuhrWDLrqexALbIc686fmTs0xyjU
Gdr+w7W4fbn88th/iKZ1pMHYjJ4Ui+9behpyPHo7yYYJwC1KMANXd50Tf7JP76JD
6eo2xu+Jk4gTucnTDK8lopdyZ+zYbwjOTaiWmhm/9Zq/RjXIfPplcMe1Ra/t+45S
DaGi44oy04F7bp3OBolQ+a4lWKb5n1QtOdRgn09AdRtvmdvWuopinGfhhrep/mfB
cnGWO/4nUyxziorC0+nXHpPB6Q4ffbNx6KGJVTp8ezwc5RdGv4U/V7ROFIAMLusJ
FEMhuFehANf7nWsLFXR7a3nORHxymZONrdM62S5tt5RmTMdqMwUZFS1SauMdt73t
odX9oMsdMpJTUbdZbcpI6GvPow3CmDYNkamC6Hfu37bGPkX1M2T44fMe8vnsHwul
MCwmm02hUVeV57sOW4Gt5+CrG4hMGwBY7cg0Vomw/633NqRkgSXPX9ON1MNxzbbc
3/sWrPn5t0ARnAWa8BjAYvXcxCLGzW5ag3oHFGUHVOMyc7is9WXW/mBfsK/2OM8n
CfQCLfrBTaUdGhdZgF/0CHEwv7Zd6NBIKVLDWow+KtpgXQpHRjkb4gmcwFHlsSDT
v+XbF+6PRmf7FgS+dPjXiCOMXlFUJcgmp9iKkjLhGj93bqS1lub0D4w34kRrzuWT
TPFJmcYvry9SSRnCiPD3JXrtAJcHwpmHE6ovIyu70egQ68QDZC4ewQm8TSf29cBN
gPxXj05y80jooOHKYNXcj6Pb9/fLGcfPOQPb6oLMJUyQPT6CT6pXjHhua8mgDZ5p
EJf2RtxbjBtQm9YzPX/8ICEIWIrvI7N5h31ue55iMQsM7y7EaOxeMJs7fGdA6ahS
jN9YW2AIRx0oXen5T3f0ZUpOK8eTlQEtJ0gjsxMxINbbPMn9WWQy2kt1Lezhx41x
J7w7dZ71Sf3BQtysdjPql9EDdIO8S6Is4qa4SAXojMDRY8s/g3csRmhN/mghl3Ju
GSdVv9z9pJgv+U4x/BdqXOUMF3h7S/FDK+Oj5owMWhnwBAR74HnuUqcpxyqoUXT8
aFtiXOwktwC7nhA5Vz5v5Vdc1fojYc9uArDcDglTNCzXbBeTtmuewTobRkyKpLRf
tkWsmcWtyDzrYf86qRcuCUnMybeYLknmznNDuryIFxMYwbrgLLUT4uzC8zqETbdF
kmGWNSqc1UteweHixBERs3s286zvlwDeKL4MloxDJMNvLfHOKjJprQaNsuPUrPNm
bhDInfUqkBCISEKlZNXfEj7C7+VSa903eFksTdoxXbRUs100CgXxZTiXnyWTv8sk
Mb1ElMTh3zY5v8UEee0MWRbLxB/xwvy1pVykWK7IT4GmIWagFBjXxjVkufkBHk0k
ZRwSP3/eygHJZyAHzXQgpx2hdVidBDznDVTaqrZYtD6xDMLbK8augA2CIEU9cV4e
NzZ9PbQitRn4FfypauwUSiuCynegHRGpAhEx3xePcu2YCmHfkSlK3wRTUb7az3pD
WUJpup8UuoVG2lmiAY1tMK9+dlKugacw7GsgeFCwaRYTw5nj2f4fZBfSM7BP5tl1
ZQv67G6ZAxT449YpFrLXRzYuP0Rr195IRnvXk4FMVfRBFUVnUYJ45ACnqChYHr2X
MqKRciNi949j8ytXCTcqyxPN2lC6dx7DFlTNaabXqFEToeps8oW/1RDUvLxZaZUS
wFRt3Eg0+Rwj1+m0OnubiVz2dMejrOYoi3rTFvTvw6gN6AYxpCVG+zgVh8cJKKvu
Nhw6oxwD78icr48ix9fCOjo6gPVYmq5P646Iz7ZHC7ozuJXnvIGyKJJsexCgAyNN
pEaWHz7MEe8VQGOZ45s28YGLEoUkbUsGY4hul84boQvc1SS3YKcIdEjlSszLNj0M
D1CzpFmeTClFeKE8dlgSKLdAyB8mCPfg7/RQFtbokruJKj4na/8YQrC//hUAPyFi
4ROipon6guQVeS78dWjozmp3LQUIZ75455xsBFkbubXhl7D9AIMCSh3UNe8wMG2/
mOSLMvqKK1Q+SH4Oz4WCs5f1LQnuQV4+iMVsCPFN2v7J09mohQ18YzXQCUgNoAb1
lB12bgoHKF3BA/2cz9kS/1ksNmDYk1Wf2sGavfoPxh6r9Je09SvV4PDypPAWIewQ
zamQxL1eDFfnTUnKwspKG5ZQqJOwVUglaonMYdOw22MJWdj+aFZ0sPs9bDhqaEfK
KJATrwGZ428P9ElA07tzm8/xeYR2MaSTtvaY1Bu3GNSdsEofcC0Rk2qQOeGx1mWR
xBe88aGdzGPbkip+vSkgo1pXv0l/1/N0Pfi+VQWuJgfj68BcXyRMELdxutPSV1fw
6pIBFm5JAsEjyeH191kdUL/nggRgQRi3k9tVISPdCB+zbCpb55b7glz4KpzXSz1F
tHGPHkTPF0VnB4YHdk7KHyd4bj49+nuzNOG3dIoggUmX7xTDCCWQrsVSpjb9gLKx
9/oF2K84l7cE4CdJ3TCy/TMtogp9BwEkUPtQ4hFrY97M4xzLIU4I0RBMcwdDpm3p
45r+2QZKqvcyg5696yiMkULwQm8lU5MKAnqScjk9sHvk+TE8bWknGF/ZyX9zhLnB
rA2MWkg2sp0cSdowiu3mOqMEcigrDaDqcUKKppc9Q+D0Fn/r2gRjQq0/NdtqZMnd
NQmNuhtd+tz9ScL8/QrmT79CPZV/XIpM+CYpUlneu34bp98RuF1YXUujxxt6ewDS
edXveUsrwTA25XU0GSKxFS9X0h8D9urPr+ELbjx0/JI28+/u59gmttZXrT+Iacso
DZD+9eTToojqlJgC0Glrp0tsWt2WRP1LZq1I86hOWwZac9pbpRO9M2cMBmrZCPly
9pgcZ5kzUmAuvmw4gIFbH9owJEaty4ktt7dIBR0DD3mqPIgeN2AilEWwmHDz5i7r
6N31YmtsDHzIPI2VOPtEn8pA4FD2l5rzpxEAzGmisOePZtQEc3buxnjPPRdlvb9Z
ayq+A5+gI/x0TBrPL9Fm0wr9+UHry4WQSg2GpYlRjp8cKVR6ECeRbELTmVkyBM/s
+TMsNK8ndZRFIzhEaC82ePRUtIbia5sKP/D3uN6QyCYZNuFVr4iUKIr06eALWhK8
+u+dxyiroY4upQdG9W0Ba2Cr+XQk9E6EmwUYfTfxXHiHzIdeCHRnxn2tsack/xgj
Kh3np0oPvXYao6BuCyVp55ooec7wPzTaL2lDu8QZsBznf2zI6Ha6qpFvlAoHKoIZ
NaZyrdiC8UoGa5W33k8XsaAEvmIdwyfBhRVu2UlZPDOenJHBZYFw8kJlMBrbELE1
CZwbFoGYw68m12Keee4g651OJpAgnR9bUsSV5z/M7i/+dB9T8g7wY/pkpeUz0cxn
j/jgBIp1fQ2aaSa7w0VjBT9P8nOsx2s3Y0UpGdT+TlWREkJLw+5qx1OdvplWcizJ
TpVHoGa/jcnwFjYVm68doUtyz+MP7f2+TVijAuSoYSrpPY1ZxVeauUS6LY1wwXMc
0xeBcF/fPlrl0Wizw+rlUbSFG0mglUW+MBmIDPses+REPhU6PEsXhbuKuJcJ4q+3
kEh7T/cxSjE9A5efBBSk2tZqjTPa34zhdcpoW1oo56vVOiniYu3Rqcxnpx2kLsd5
cHOpitWvRYHCJbFh84Sz7VSBOaYJESmRpwzhz20LfhwOsTOJdCSwpUPLA4FsMzAA
qqUHIn5Fq3laSe07oWX9eHkxkxVj7K2a79Z8WxeSlvAEr1UMjGEdONCwdGDJCJ67
+V2c172eolwCNcBjoR4Dtz+IQ4mMTIESmCNZfyzWQnOShyfnxJBahRChkfqxC/Ii
XxgXKzFNKtCrSrFwShOe63n3XUdV3eLx6TAjy0GzDC7nwe4gXQRzrqPDS3gt7/aq
3Wh9R8qxLkUhCWV4VF6tHr8DzsJHniJZqQT70SL44brfR7kJX65ync8iiZ2itQoX
ASszAtS1/t4JjEPoWx+eh2jpCF+ZGifUq3oj1iHkEnTlQ9FvZTVy1mmNrA4EiieB
rYtnMCR1x597OfAySF/OV61fk+WzkLtVx+zmgtFTBOhQKmjmNVFPLHMmbULHSFSR
a5iWdsFsvA7qDKu1tqHR6NlljZvDrKgkBmyWbb5kmt1N41XrkZEQxSr+rWwfKtLM
cZhnZH3qrl8KbqvboOttXfrBI766uWfDAQnJcoqf/kirFK+ffUJhruC5GDiIgSQE
bBv5prn4RSId+O3KZYm3c8MqWe2YsmYKXeXspF07qNvZTcg2o/rAva2okY4Dvnpc
XG31DwrLtN/qF5H+eCnz7Dcaq93KKznPYM7o5Nk1LEBLgJAF+5VzY4MjYu94lsv2
jo4SrCN2sk26RQTAhoVooGievLJc/LuNGeeD02Xfo3d/1g9vB6DHRh0NNwrvYiow
LcHiJPUFhO2fiBK82Bjty9sJmgTjId9CYQB/q3GSi2s8ZafuDaLTLvJDIIl92n8F
dyyhw3EcWhXr9xts50MasuQrF7SXTHdeVOnILQ2sG+CPGN2XncCwKwh4pq6mTuyu
gEzrVbR5/NAay29fPyUDIbeMJRAfVpVmauUR7doPKqywaQXZw8+l2SZamecEuYip
cL+dP2ri7+7almwYDF+ORruwiWrDNEfn5P7tmvVohZSl5g8PZRE56X87nN0W1u8W
k9qxl1qTzHH7Tf7CWAZuynHTaxIQHxEANuLCnge12Zj0SzwL5PeZhtvIwW3voO1L
j/xHsz9dQtfM2OPmAZyW5PfsHxzSBteO8ueVQkPOsWtfhkUGIhNs9fVjZJbAkaNf
HKt2Rs8/VYD8+qv7D7i7BrO4Tx1vOPQiRH8Vl82Eq4hpO6S2sa8Z27hQsqwF48nd
oSokNC/kcJjj09PAY3APqX8s8UOeoFpdJPQGgvx2BnL4Tl1jnA9X/dgbGnaDadyq
79IiwCngd1mKcNPaDfZsBh2/XvViH0su17hz1gRmYG4F7P+TjDri1mNcOKH19ch3
xXa/eUxgnOJIdJseiIlthAkvTH1J94qJWUnL+uovsQeUSuHxqUcY4NltKLNvAYKo
iUibUJwmlI1KAtP/wFNwV4Odo7+1yGSIB7OqdFr95Phik21DXRaCofIkuedUR+yy
215mcFmYpyFa8FShy15CGWZCIUyuPrmwDE0uz50vWTmKbZS4cnpXnXmcQ/q2kIt+
j/vfQLBPryAZW3ifbz6zLBflGwHbA7gKW4JEsmMYa6aJZLk9ku/ZBKflT4YupBoc
h3s3xOKoenwoKkIeQgpnBixcdthiEjIe6luEDtz6B+4+cveYO7jhvQ1LJFchTpzT
G2+ROKJRG40LnlcqC+vPiZhh2F+eX1ZG07KIy5EGs14tqpeEDq6pVWvy+WOTY+1U
5mFl304bcKKBWFqMzBUlZXLONWxtphb0wykJyRHlZkQ6c8YUkQEgnRIt+SS6OGG1
yoKJHDteNlmOeuMOtGc8+kLWLCbV6uZJ9O68Y3CS7lekk0kXyGC0/dq65R5upBux
x3GULm99gDVYnWLJ5OTnqaQTdQzAMmBZooidtn2cDZBIMygPNbC47ZH2Lukcnhg2
unvXWh+Tdb/Y3t6xQK5m1TSZtvJ8Riw+USU/AG7AWXcfSAaLL+trheCLTGgKX9cV
ABb0iccfse19eIsYPlIB/r2873nOfOvkjJ/c5wL9KhmxUprbThqKl3rg8CoOir2D
fhHxVwhRnOPmMJGSi8/uQoSbijknS6/S3Az8hal7ZkXfavgE6s7Srs2Q8Hx/q6GV
forsRrDapiRRUIREAVq2TLgcgXiNFVuMQA3RMGFCcPjvhFd6xIKfgfYs64e/8H6i
ctqRWPe7gjRGjX4N1HQHC6dkgQ5CumQ0VbDJEnSUDMf/XhyW4Sq8wH7SNrX2g0fe
9DesCQ01XfG+J5tXz0YZNOlfIOCauJwcCcSjzZD6dY/0zm0xoFPG77KPM0ShlFbM
RBUK87HhQd3QLyZjY6sCRZlr+uLr4TfgXdF7X2xeG67gxhki7YFC3h43ZBTiAJl1
Gzx76a0ZOV5hLxz2CC/cquzrHWFOFsJ3aA8W0qPUqGmRF3HrciW+fiXgMuZNy+hU
UKCKYd4oAurRyYxEdrkrd2tpXkeaHRlXyJzR2061qUuZ+qdcDV/IEiqmE4cJdxur
vNPZEeTqTeOGtXCJpL6SxLYGpFzDzMjpTv0aEs3DC9eVuFJ8gesiwo+gbbPaulc1
XBl1Bx1NndyYR2t8upOsK48ORqIU5bpQLRJNQBgMY+Sc5AkzUsw/+5d6pKc44tTe
ZrgTMeca8AxWGMZtPGiuKckc+sOA7+2oNpsr9xOiHiLfIxHWr3gfMJ5KkbzsZVgd
o9qy4iDblPuXziPBNQMKKuMuyCyd8evSAQxX6k+fIFJS0bwGBWM2Lec8M8h/bsG0
qi8MW9F8OaYzgFzhGodWbfnmwslBKZWs9e5YRPIuDQ+hd6VADH1oc1gRzhOXDXmw
B0neA2Upe9XpvsP42LS4FRuWkOa7Xcl5znuJXCzXqTAYD//tkt7Hlij98ZGH9Fqk
y36DNlwczVqHSjdonAmUJTT12LA8d4k2rpW5lTauHQfrW5wz9g2MSNa98cJ7i5c8
MMsBR5zarMQfXftnIvGBi4KAAwKYgNJd5jYWoijWkqdkBqwwiwYr2xBoQ/8rCk/N
8/zypjh/iKtgC2dmUkdkYjU54FdTIeasR0Xk1Dto4ojpi5RhndpSb1yu+SWjFzCk
CRvfhAXgatsJ2X5dMpKLALyuRNEdBJhXjm4n9WZuQzPifOANw8oe0+gLDFOwDt1G
WjG3xYs5h+fYEtMcrXyqC7m8IyeZttQTHUZKWQ0Fo8Q3iXAcPZBXJGYaf2yDIZmb
aDDgXH1czsXNirdDOVSTE6Cet6AakK6UstJU3s1bFAwql6PB2yWYB1JV2qs4p+QV
1krpezjstOj0x1z6/K9sc4igpRJ+GdevgW4tGpTccnXWh5cZtfaSd6SAgPYBC1S8
yvPhg8mQ0iDyrtg5aNcqHyXj7kVWRpOJp22O3EGZpfWKCvGsoLxU8W4OXeS97Tbv
c/ClDxZgjHKG4sYo7XtF97BczBKcq2cFM5pgWr/551JcZ8Z1noSHopUnYSeabJD2
lOBZ6gG0zxNWRO0fQXR35rrylZNq5/iC8d59nhjII2HoZ+tRJ1oYhQlseUbl3WNO
ltLSBRvjeKUSMV33TBZxRNuCH8SGtpr0Lr7b8+QoDVt4PE3mjWtIWqcUyoBiB3LX
z/7+JcACLer628uGy44SFF5sA/qjJ45Fl7NLtBWSQXW5K4EOgCtOJmra4IhN+mPe
9Ja2481/BZO0voUupFQOIeIEp3oIjiQHeaXn1O4hrdBnbAQ2RuQA3OSmpNrLdw3x
gy/XjiYxnd3l81mCStS1KaTWctlJhf1NNU616cUJw3rmGSjOAkP2Q5AmisivzFiC
Zr+bsdqYw40KTKRohTcXLmAOnWmjWP3rX6e1+x+Y0/UZ3PY4IfBgZbp/DG5bbaAA
jLXKFscx+XwwR8YU8grdrqGwrA3M6d7lnev1fPTK0o2ANac3prEudMN+H0FpLyVl
CiFQvoEhIgkcKGQJdzNoI6Voz9Nxq5H1uRIFejExnPEaV3bemklub/S2cBy/XJEL
VhnyC2UqmblMapCkvt/mObhKN4sDRQNvp2X2V97D9yfm0MjOH3hht/JXweYz/leQ
ip7xKuQ2YaDBFYwviZQ/jMmaDajf1fRXvFOl/OCM0Lb2mL1TrCIWACqbb/82DN9S
9ZvsGkiKBECIKdSjRj45Jvp3qjuXBbl/6qWpT2I/HfuwJ1uVIiGv59MkBd1sus90
stgidIFkgA5qh+XVQiH9WOZU4T/0IduRERY4CtWv0+2++388HYjp6ruladCF+uMu
3GZ6jnYjKnQUByRWBdxyO8Z6y2yV/6zV0VVhlwy51k56O2jVs3ZUc9LBHnp++3u5
T2jFmur1IvELMExizcqYbdXAj+oGVN5XSlOe1psbYxXW0GOnbrnI8iqHhZXZPt3N
4cruQ/gQrDgci/jHIawwyZ9yyRmnx3tpZJ+qsYoSuY9Vv1Iwsn5ALccIBmu6HyYs
dFULDN1gJj96SKSyuCMTTLYSwD/8Pgzypp9Age9MqEAjpa6eGTCxd4kJ/i9YQvZ8
zOW6cBFEV0MFB/Kh1mbMZrHTkgVMyEijG9yWYGil5GrI4+3rXoYMBNaI2872BDjl
jxZ0zJ98TQSiL9XOj0GOM8oVA5nbToVnK5edQTND8hrOO9MZ4MpRIBbUkQ63EJgl
X0ViIim9Ny95LFtkJFo+R+EaYpo6Pztz5VfyjC5hCC3XZ3CUcTWMMCRFFtNGGeFn
3zF24MDf7Ggu1SUh6iwL+eN9HM0RzfJBqhOgA2Uc+he5iVoNwA1sdBBnZBISVPap
dXrKkFdmOeavaE1VlJ+z9Vcs5W4v15xuO0/md26iRc6L/7ja8vrMGm2leAVLyYmS
zHGQHwwIC9FB8uiB+5ogOAObUQLwfRVhQQRFQ7dXm2xE82Qk2YRg3/+hOSB/wJqq
ZcnOot2nhSupCF0XC6ziYsxSTFWUsddBdyVAidX6vxVS2QrfGTWrMU1PqSJrQWyb
O3vWlyMRvMS46OGj5ZBJWFp72sXE4ZXzeJkQ+LfgjoBtD99Mams9kZXFI18w8Zci
5qq5MbIoAllw/zb0olG+/iYFigSM1g/7fI6G5xVWsQMc9/eOfAWFKihpNRql1uVE
NXeF1eg/293oMb+Pe2BxUXqNKdURXD7PD2e3ANt2AYfWTfEJVbL8lX9RL/pM+CFT
8V4m/KUXAz9iW3roVcWyYIpuf4omkWTXuFSvQTkwqpQjz9K6EIQuommaDwVlBjD5
jE24cZAZNgocAbEZz2rSjk01M5jzO18NyGWDZByNMKd3sG/RFMFCinIivmBfZZcI
1k7RCkT0CW5NY9AD4iExF6VhuObw7gp5J9eJqUYG3wRCw/hqZmP4+IGkCHK9Lns4
WXFnPLqB602VE2/Idw3+lxVYZLxopzKn/EPYAFfRTS2f2FzOQIu1I20T67ER8TLb
L7fsm3+QjbQ72Yg1szh3zz4XRh8DhzFbroSwB2i1KcIXNDnpHNBr4Pj0zR6JwKCd
COm3rqnMcX+KccHnp7HAbtAc593jOEc9DPxvzUsyQBSki2oG/p2eXKsrY9txQ9xb
juxJ1ur4X1getEYBICYfsk2v/07HcW9PRRe8Lgs42HOrOBwfeBxmOjWZtQoY5BkP
11BDsdyC9PDjV8xIBx1hjy4DTdCimHo9PYy87yFSQk1cZgVyJucJ1ENcwo+97CpE
VGL/85kdnnOr6A3auogb64sQvqdWY3CEzJAAhmIiU1wDiwRSgAepcTLTzsfNApfi
pM7tGdtozhlvO6DVqcPOB7ZDG4mNunc9ZTCiAPvU84+LCnKrIpyjwospDZ5rGpy/
P+1SUxpl1b7WZLZVWfHKDn58NgCnDdDX0s6Zo+txWvTosx6T8q/bZlBesWULZ88a
i5Oz4ovB3hVtYoEQo999RTk3zxm+mAm17DAlZKPk8WB74aH7OFhWNFgKUQWhwyAg
AJkKQVUqCgMaZTdSEFdawoCtie/NmJr+8kH/a4eeJY7oKLIqXVeyxlh1R4yhrKEL
CkTmp3AQA+aKCzuObsEb/CJE3SC6G3idRYC24pFaGD7HDkAMvPWar/6fr+v+IYZd
1wRVTUBTDu/uray0EKBXHhX1jI7qVilvAgjF/QzzZihfh/MoMCpnDA0tIRKRPSnA
8Y983POz2LkpclJn0hOuNM+8AY1j/ujl06iWLdHJluACJPGRd8UUwE+T6j0te0mx
JLRj1+ulPuFUWwx9SAM6cWDNIms5lxFE5PUkb2adxomWQIWzmDG8mTDis4uivaM3
pBZUHCDcef5UqmOAMDNE9iviM1qbzFrrsELNWjNMR9Wxr6sav7pBC6Y7CivW7hQC
G+kYH6/ACZOkQEGvPCGQyNVtXt7BZvwB5lVvSBXLX7FbDXKJaH7VP4WC/wnE7VjP
kAJoiq5OC/CSf2cW43VzFIy4A3rmBdCCXcwEMfrnxsDUimV0eymxDr51e3yVSV9b
onANKVjUtlUmju+bRVat2SvPVxU+BFWzWMg12tuD7aPcQuyuuBsk4nrrm7ZZtNrM
oHf6kfuEDSc6GnW1INzcwQHFKll2l8liGPZfgc8TfrZ+egb+hM1xgqw662sHz+Ha
vXwEk6IVrvMQVHHLHMo8ocO69X/7ZQFbfDD9FybCPpcWOugoQjZ8722CS1Ij2ZUc
f+dcfNCRXEDjrBes0lWLZnkbitQ/mQqVGmRmKaFzfBU7gh9UJ8gnSiNmx87gTtl9
XIkB8fYLhXVbGQ7a2ALSDvwN/SSVi9gjJt5h7YHzmmpHWxH7du6VNtYtAQd+yn8w
w+Q9oCb5aTBBXp7Xmw30wrhASfUWUnS4Z7IRV/I0DMwou4+i4mVkvf9rBdAXS3QH
CNJA9GyTZkFgGrQ7rXivLSewTRmcWjbZe5FYDSSoF1ZD/DMZKsdZ2pAkd+0BPYEs
Ta571y3Gj9FLZCWXKU2XLxMutORrvh2SMrIYbywAPVgXbYnh48QQrnZ3OZcvs6Gq
KaHow/tf3Fj1e44RH2Xn4PVZUWfEwmcWvPF9jb9r2A+XD3gv5myE2S15kWekN+wh
j+RlDZ2GxFjkKbrobaq3N3gxmw/56faIDdcaSuVDVT+s//Ag3qEjaVfGTAawGN2q
dt9ZyvQjLN+IeVbQDqJRJwssyJBN11ReQxs+QAABSBecpqJAD4QBBsh/GGfFBsk0
TMVZax4gqJ0KncM5a4BAb3cX3ymSd/0s1bOEda6Uqk/FCAySAfLkHvHI0bBe+MQd
mafyd9V8PFF4eUMWG6xVKb/PXgwJlYeCwzVJrGAl6tPRTvBidvCyuvWbG6AOM+9y
YADQiog48f6LHRDJEolJJvmjwa52yA8PzSONr7aGx4oVokOHl3yQH2yMPNYtzCYj
GBA/HCm7YalRl72CSOzrG4Wvwqt2A4aSeTLNF2AA9WnSX4xnHaPjA1CRKzJZozOJ
apAJDnmC8Pwz2iqfKG3DPEj5kHZliEKHLY461lbu2pVm7vkEohwTM37+zFjy4zPH
Uge7n2bW3hrQAcasKswHuOMCiOJ0q7bzL94z46pg3kTOn6q5NG63z3plpkeSCE89
/qFhotEWxMB7Evzd1+h5ki2CvpNVxlvwnt1z1Te+gG5/XdjP7somb/5mRv+IQDQI
AkEJnTMeuKgrQM3sx/BrJLVZW+PdG6Yj62P6KSV2x0xooZPiFHzolpc2PgePtGom
YdaAew2FdY3yHgJ7Xd4+eYGdc8AapfH8v4ZmlSKUXpvlzerdhTn/syOuYTTVVkVE
sHtMi/7LpZzGEgQ4QNTN1J+QUx9EUuExV59Siiuguo9FHXRBHb+hmngAGXHyV6YV
t3ePOYN8qRIrc9brAqX/PbQjT+u5QoJIc+hATZWuYYPNoJGwt57bUDmQYEs2Oo9E
nmt/QvFU+t/g5G1aei61CtcU9r2gPj2pVQznafhJxFCWDysClKm8BX5Jn/e9fRfH
22auxKdgJhINI5XF8Qhg72c2p9guL8MEF6bkBmqt/g0lYk3fJ44u4xKttJ3VnL7c
eaQTUoep15wL0Yq/qg0ySf/lSe3FUreFOyn8uBhY7Kep4gH/sVNrFdf3knr55jR+
Tnv8IeqsYftL90KzsJ48qqL+G0d3fJ1ghQL41DB0vnRDyWmlRrdjwkvONHBcxTIE
i8pR8Sab1sSljv7YldUHWKIYxA0KqzZShaSODpNqFWWIAb/PoWa4PbT/dqNz4hge
fZZqzVWPgKFKlhV/ez53riToGHlZNpk+DKd9l0EUWCgp4YU4HH0z+z/MMFQKUFtD
13G7PB3GOiFdXwaOri5/SdaEqF5OxByenQlyVClELzZIRM4Bd2VP6jNnaouTQpUP
oM30NVn5D0KURNBSDzTRSjlkxh6tIR4+uspHQpUb41Ny0mrba+oB5CMgG8YYqf+F
KIBRwM9h2qWSHavtT5xPrtdxnNhuQkYIc8bWO/eJESfR2XaPgtu82Lis/+mbxcLv
ziukKTq7Qz1i1YZSrKsXee5zZf5Jp5VzGFa1qucZKEeXnqqX9skEd3soWNZygeU8
rQJu5+L7ZPn+jp9fA28lE7MhPj1+9dvhbmGVItfxXzTHmvx8T4qdMOjRJTT+42Ka
y8RDN0LT6CGPgp0ygNAuq18HPxRxXNBqJO5t1Ch2hu0bsoKrJ1/WHdRHNEX6jMVP
npPUEFFV5x7k9gWjwXH6JCzUSWqBdDbqIuNy4DaUfiIiKpx8M/HsmvdHBokfpHav
NBzMUBkYH5CBeISvkDi7ANjSY1RUGKlFfI1lFguDVAq3ztzbSbV99BuExTd71UJt
dR1hMh/od/B/T/iyUQBo+pMptxwO8Sd7B1rAuM9oebhF2JJMwv1qJxxwlzHzimM3
tEKAtxIZoaBTtSsP/hsF8K5JaOnMK3Ou4A03CJ4nNCzjXrkwLRWeWWilAOcHu+fN
KKgmP/Vv9TDrsPHIqDuJSHcSt7szYXCqaxP9txcIfKwJaz4Br5r5X12UCDzioCmg
+Rc0lQxYJZugm/6z7IIcCGA3RH3h1UoAtb+IYziGkaD4WIf47A/BkgXT0GaJ0qGK
wtYiz8gExgmr37Y1fB/VUfXyjLmzt8IwLUxg7wEdflVm1SIGsiHIIBUIurk4Et5D
Kew5B5nP7sK3Q69tuQ5xZIjjYa2oFhHyROyPo3f0NHTO34QdKN0ab4DHDHsFtXgs
UL8VJtuZntOXVzOXij/qdc+wA8s8WqZ19TsXZtiv1CTnocgCIbp8YI3pZhTYi1Gp
7Jmg0YwnpZzkDHgAhpZDri196Wl/89i1ea+xxvSKrfyxmE7n1IqXTtqe2ezt0Rsa
hvCff3y2vjkfeJ4ZZoeci33Tni7TYEbwSmHIWk7e8txESBDSi2XsuVGwpnsnj4DH
sb1kGbhoeGnarYQ1F9FVFYw2QTtW/kHhc3tP7E/U1y/34kvOX8wNYzQxqoSLKwWh
CK6EheeabY6O6UldsfAl1AFYgn/lvJ6Iul20ZsFhvCVyjjIAJCjz1bg/4WvLMzrZ
dEimeoCMuumO8/QB4C5C+WMJNXHszRAsw4sISy3UkjmVpOr/YcwVBhyV/dcd1z2X
cM4ij2/LJVGtJuIkjnY7akIR7s/qme60Tdy5Z8csohaW1ravNyerbijdCceEFJGc
jrIxd0F7gmExv+LhqK4WnGEOIAjY3RUJHHd6DfHGGKnz9+EiqsHiez9umO5mucCX
jbdy6wGpTJnGPK1IehuR0mBdJWrBzYHk/WkcrFuyr849aVw4YaH86GOMtKpyBrbu
WraZSS4uGK7L2ICuOM3IqRXpUSywrFWQRMIkgF3obM2SdhDTY8idgkj2ubyPEP6b
F6D3Js3/rcHQB3UD4pqqUOst9y8VLd9+w+SWIYcJq9CQMveQX6bfayCdkD90RPxs
oDsvGTnSvfcOtxy1Ms4Gef6jnh972ev0PvZHjxvt4CrWk1WTBd7J+bPLJ2wjzcnU
srWnJJ2P7L6eSuM25KK/NjQnpxLpP2Th+XZfL5AeROEMswT271E68eNve59HB2go
azJHzclnvfNEABz22xPeUwl9ag/zT8/AkvAZfEfHjFcrUEj422W2wR6mRI3aRqrd
pPsLhPiNsvkDol609QTGYCOz85FooLwLBo64qbaKC1/ywYNAf9/YD1gZ3SGsJRSs
HS21J2ws3i3sAqpvGtBvkjhXqJG4TFgQ/sRASKIYPE86dJX/mLJC6YuP5Vj68gAP
XpLSx/x4qGytZb/T/n8LBEnccd18Aurn913eeaD6AV5Bdor04QkJyZYd7xBtvd4X
T5SbgfeF4cH0g3YlSH6LRRGh7Vg7RZhi5KTQVjWJkV0AqouXOxjLv1h8yIu5z9RM
Xag14Nv163TSejJcL7jDuGacjWW3t9fbN6TEG/50QsqMByNaiCgWAJhf6b7grDJg
FRqdjLXoAM5uxm7CoR2tE7hRtK+Utk4Q7Te0+mam3P9gaSH0U8SUC8W/7QqyER9+
7hiS8HKafr8qrvDt4JxjlAWsXC6ZAzpUs5AlcqI3e8aml8hIPwYl6r9iCWXg9JKB
Ysnlc9h8gjPIplpHZXeBoBuid9neXZvJhkWiRITCam4O3B6AubnXrB0OVypTqq8x
YuueIDg9C2sTrAWx4zZeBx1oWb+sGa641vRYuVSbTe5rQd07n+FZk8IuRcyLNrgI
LhQr2dwW0Awy2sC5kj+WA1YTeuMZ1J60KTqbzAoE6jpoj2TWW2fjJB2wQuTXBW3D
WgiqAwTW/F/hh6F0AG2pv4WLbbol1o58zFT/neNCcEQdXZ6vh+a0zwsW2Nepeh/2
Fb1WYrm6EX0cBS5TTUQ9DQa5HCszEZDPeWUSpCXJKtmKW6RCsrL+XiprSXEbPeVA
/KrhZ1VStfeU4wwoAf0Ffa2g/wY7qy/Lkyt2SRqn07RKWTQ0HNmJNDXG7gbouWSz
uHTJkhR2LzTyG127SrIJmwkJdfpBORWskG5PY9uSlCbbsVVFRfYW/iIAt7jt+/ZQ
L0XacfYxkqr3fnR9dl5+U4bEwwkmXmb6/wi4XiAvpSZ9ID4lyCsYfUXbjic7fIzE
RscLZcXloFY6rtUXguW+Njf2qgZeG69zfrXBT239sIGeI3N2VMfyNTjpYan3YEef
rdxiy+7wKu1ZCLrNtXoZBRFB8/kPTfQW7CNJDl1H0AyH/SCfkuh8Cj85iXnmwSIm
z8ZM7C5ocMmPyaw1ij7DdUrxXPGEmSgWvUoWIHdSmUzgbHH1nxqonkkATPIsM/BR
2Ds+/25JAIplqpXX8Mo0Vkcstw5GqBLp66UDUsYHPzK26YdI8GYDqBk0InHq591n
3GvLU3QZaJRTGrcSKLjsuk6ur/d44y6QgGW5XHiqC6/QW2yRz0eYpnDHwWGLOPad
yZJFBRSipjWusBHbhL2u9sSyMtK2VSIjGekNhhKblCNQzo1Yre9Hnfr1F+zqjf0k
4FiYbzNrrJTtrEvmRM0v6uNmr1JTXb5D5Htr5haGfi9N0WL+d7kXLOLhzsi7ThXX
f+C91tTT5u0ssKNTg928mZ8RaupquWmXEB1oZDrBsZgpmkAJqBTq4i5PT8Yv0RVu
hwd3EXGZeOlpm1N/5XnGB2dJWyEOTTIzt4n2zvN+vFgKxHWFdB69m1x2p0PrPUks
NWSrFtBnxlZ5acYHT1Fd9Hv6mlrO9GjhxkxLoPk54tZencfnnrQkMgKt3QwjNDRe
JYR1SlUAvD3LpUfyfAbI/byxbYljqBwUsOi6aJczNqV0bng1xHAkFXO+grZQEXNs
lng28RoNnfY+3zjHdgZetM9RKxRf69TLF0SwRkVYNNX/8y0d5x0gmH46uFjhApa3
kFekFXJvFwPP1BTrGK5f3uYA7cWznn8MpKpVL6kw40VXNmZ0UsqV/8Wd6UiRlybQ
OubBeAOHMt6CSj3TtD9nb5Fye6FkHO19DNu/sw5waq4/kTxdjJ+VxmCKSXpBYF9h
VtUWG0v251BULSbwMNvjiZInovh0IV1BpFaWFAQL5ql/M5SgeyfoMNR6KQGRJJIX
6tV7tdW7swCN2YJxFXjxBg6DjMqJ4JypXYr0C2wWuiqEqKa/1PaGZGO15QvvH5IH
OzO/AlR635KwDkRsHP5rYIkwY7+t+rRjt07Qa42OcL867xTCIsTVLhGpDghpaSSV
lD3GtfRUNBddMzlfMtmH8k8St43+xZ2APoviT3TWFDLqzTOt5VQbtqBqF3iiZbUv
kDqBEbVYPNP6hc3ra4N84pYcD8p5tUK6eS9yfnqVS1m1+0yKFOLoBHP/HJYeXO/f
Qus/8ICKtKl3SbEkkTY3FASK6GQ79Z+m/2RPTAj3SvbB0bnijdbgFchD4ATi7fVe
khRWCncANAgb4NYrUHkpcEB3KPyA80nQtf8LgL6pyaL7XExImxasiD3cxuTWHPnz
i5ejepAkg4bWahzA2QAREdnDYIN12jdipPmbTFIrBrNx0pKnvtnjV9ioeUoyJH1j
FbnyVNWtfM1gcw2sW+YyRdX9gaqJFrmmrOyDksHYGDxVOnno1Te9w0XBgeECEQBJ
ZJKM4jeamPPeIA5s5whtS0FPSW+CVdWkV/bELI/nZmGlZB3z6j3uZEQHMiLoTBDF
ZF7JMrBqgWSbCF/l0d/RWKjMUCtAcLFksjmz6aaULYClPONg8IRpKqLzRlSRvJOk
beIJ73WSXlnUMXphKbFa6UkVPRWdnSMOeS2xGGclC7CXoOlYmZaecHRSCWIvIdUt
mhWzdR50lzW7OykvpVCwsCuiH/7fPv8VJHKpFktU1eaXC9WOdHO4cR1SUwfDU/KO
WSNsHl7rtjzDyWIXviGSuV2L/FT3LEFU5emfcwD8VCAU0P8z4CEvm9G+LAB4d+1Y
XUq3+y8XjxQoQ5hG35vlvDpAAY6kR/4BeY0LsuLOL55Sp5T9p9Npi9UCvoikTREJ
oJa0cA66yakx8UQumN2n1lrp/i4aQ05wjOWvoE+pkn82c0cTrGGaBBvzZvMd3nkf
czcybICMsENVv46o3xXcxWF+oTkA1PdQrdhp66Ypqf8PMQ9UmPpAoHLA7gAbv50m
MuzIxGQa4jmGbmTCUlAmvOH8F8vd0Nkp7flg18vLZt6o0TCoS4an5tkcB5BMHiwU
DqhEzLxCmxpgI82IWGXxsjcLbDGh/WCJEf4t0z407TAuyFmnUtf6T0a8pBQ5wcrx
bqor2Nc6a0D32FhRjS7/kRH9aygeMZBI79FGDPj0XwHqNdi9MA4gAGLJahC/jIEG
Az2AL3ARvcsQ7QMGhFf5f5dfyqPUdzabXJEWx+gbaviBV7Qmx2ufU5wNE+YpFSot
bEEl4ujxOMxDZ/Mpok8YOrc2b0Rdz0xo3HqQ/4p+MKSDTNNRYln8ymL6bodq9iNP
kZLYXH/teJpK9aDoq3Ae6fe2QvWnDhCFGwdAREZOBQfHld6LbfVngqfR4R/WE8Km
lKOvRTZlZ426zzYv+tW5IcWj9XWsCNqaR5XOY/MEiH6rB3/uIv+fmnV52RN63o2F
dAu2QGUew6G/jvR5jfifb2yDam540T3vOGY1asBw7KqCB4CVU2t/UP7U/XsTfUNV
8jUJkCh1mBHCi/VZULodas80NyupWdYVzh2L4UxfxPO0E0kKUdhPu2YUFaI1QdQC
daDtVU885JLwsj8CqjcB6hoVUTWC5bUqGNF364Wz/UyjT9clPN3sewtP6Iafuvm7
xb1o3I7gnMQwHm7Dflrvph+nOySZDNMIsdVAxY1zot9bt8/lrPLXWprN8k2xCv9O
9lHpCqtTYLNtkf7KYQI9M1aXXQoXm9/RsKBDFf/GS3JiYz7rzvp4QuckeyQRHNf6
CNG8j4nOK1kNUXJiam65w2pYbTVv5uPLcWAe2zG/3urEPf9TlWPpauCaLNoQnWFn
QLBt9KdYtz4DQvJ8/KTmspK3ltShiUAlI4QdhTypaZz08FsYad/zqvAITrTZCJxf
bMRtstresAWYBzR29A55umTqX4fr5OBoxS6AdiTbBSHYDKDMXuJfy4iBWMt9IalV
lg91tPAYHb2YjVmoABvpliUH84OUoFnl+GVHTSLNTzS0eA/PcYKzlIaZtFIk8Xrz
jm4jvio2tQPanJd+tluMBmU0h8EM6F7z6syIFV8OztIL0T+5LSZnq9DRfx/4MURj
49Ez54hDj6st9lE9MecvZGycCJ7XAOYidby0inno4khR/+NMePwyVFeREIv9ixSD
zFFIVDPnYMpH7dRHe9NPtXS9otDA0rAnKWHyHg7R4ewSeULnWMAxvYkuS2b6XwV0
gH81ma6rhUhXWlHKYPG8iCxbaPSmVFzXBZyltAd8v3Pc7SErJC1HtQ9bE0I1KZ71
/Tw0rTccF9UpwlaaaAN9lxEHJZ1xW/mUYVA9fShSUXTgZ2PJcGRg39AsvoGCDxKr
BEKPe5stz+gBpZtGvFifxMS60WVVv+pkO4g2JK4k/uuHNi4VWtOJIUQ0ufgV1/XT
BtMDdPORlKhjPZ16xBUHPU/PC3O4BFFxLPLx4Yt76Qt0AHMN5SUYAd6BOXi5fek2
I3TLgYZX2pQ3CNpF1AJpUEO1TxsS9JbhlhDMg7bCswz+gA8l43TXcWH7vlV3rd9S
DFbKMySM9PN2dOaiPmVNJfTkGcwcMRpqlDaE6V7t/ZGuqWXIGmrn0MAqkIdyP4OM
XZfDaJ+9lcIRG70g6u2EseEG3wcTrAkfyUnizCltEufEf/LmK7mrpp6wB0AVu5eZ
0IsYnv0NXQUwpBsr1HMTRu8zt0sVQP0ucl2eUf1C9+ud2oUUuR7mJTtijmxSQq5y
NtQeYkGbixsNGBGPwu08eThWM4QdPnYZW4nkMrnSNP9+S2Qh9n8IK8d2lAzbMsQP
IgwunkDblioHUe2ov5fZZw83fL1IvTWdGVOwtFl9gD2+8Ont7mxtFIQI2fFaDBmr
FBc8Axin+KfzNvMF79KKnqsXS8+YczwSSloNPTF8yTzoWbLugvtafUjKWJ7Jj/qt
i6kYdr+o8PaOlPo8evAPV2TtdvvQFTBMhR/Z3IOdwT9l78n82VguIHBvVXeNIpfU
1BinblPk5vAiliy8+PUk5MecVAcCE7ESg4aXGq4Qy0/OjNP4rXtKhpXvhBFD7XJN
LtpjEmJoCh2btw9D5/mfn3fnRCfEo++wM5kQ/n9qFICvG6j22DepWUv6Kc/C2eNE
`pragma protect end_protected
