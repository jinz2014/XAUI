// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bhbpn1/468Ggi7YS3IoOVwqIPo7VMRdsuneFtYP5KAUUbcEqbqYzkN0bGLveTuQU
kravaOZtw6k9At2KmUydFPyQ7R/vkvdoDC3OvL+z8Kmy8mC9a5bAXfTpLin35qbW
0ngsDLUrqa/3Q7bQn3bz92XYOSQgDZlGshTQ9eieqS4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8416)
nuZ0xpqPUEVPJoea4ThFlwTBTRxirMBIZNV5YBjQdIFBXDTq/Z3/q04ZjVUMDP2T
wkbY/VvaLd6hgCmIBuNtmwq5kXEl9/YwMrC68TwY0iIX1lo34Y0FFBspuyYrqQRp
CeY+j/nZoJOwogX/jbz+613+8K122YPSaDxKvdhNEdggO+tE4TLzPUAhwCawRJ04
SM0n/7uhrDxQjNy+isFyq0WXTdQAKGZEKi7zrF7WGAEejf5OK2CsqY4ohCTtF4RS
LdLZK5A9AI4VX/6u/kD4F+6XRXKjXtrF4bwFbgALBDyrpUzCG82fqg5h30+Opoxv
iCyJzP6yjY3xR8/zIeQwt4gVKrVM4Bp8xvhRyVMGlRyhvjvDVZ/XqTEwydCZ17YO
DcobwNhrJnEq16OzlsjtK4zvz6QYWTKlpKGGNx6Bp1Wso52GSZCChhynax4eDyKd
XE6S2qt2nGUf6gupH1sY7psGa9gj6uKoVDMvqDjlpSTRBwfznkbasCe1WlTXDCMT
DYiWoU03mgXyEmEH60G+If5twjwV77BbaNqFBRlDMoxG1HUU2yDOnojWRPvrUcC1
StHweHEMv4K2hNFrYVEzuDe88zrFGpQRcAH1k7JLzu8yQkSdce82fHCaFQ4kQs3D
Kmlpjg0wmCd8+0XdEYYZwrR7azMlaHO+uXllsGhCIMouC6qP6psQdbVVQQygcaWS
oIuRI9i88acGKWxVdoRevJO8ccntFF/RzrNUwnQl9OoddkDwVmL+slQlpq4eMUYs
Z71ta6bJ6DLVqrG/Z5kMQGALfgkdLjOQzQL1LQWJsuk9FgEVPqtrPiDUmqo1cXzb
s9HhykTyssFy3tsnw56J720+Orc3+uTpDfPz0KQ6XgNBnM3RRO1wcZ+VD60yY5kW
xEJmQIgZx45eLh2V4za5p1s2Q2ylI2Vk1u12hHtFzxR5ECf7l3o6BxdXrMeZDqdi
S22ifhAGm8pnMjDzFeCJyUiRnv/l5u2pNz+kCsYSXpSWyxWdr9PnsORHHTX4zyC1
sBy5USXIovKs80uhnye3onubFJf+vv25fr6qHMB4G4LbNBmUf6AmqeigQYknaGTB
h8diNmPnL1lsAFQFKXz/QG0bbl4sSlAepzKfzJ/fQXZsLiuKPaX7VLogHcJ8iXYQ
RKERFW6VIAySoyH/cSLVw9jYMrwtmDS5Ef/lnIVhh6srwwf0hdFHEDSWquAyBVrW
FOfkNHDf6eBi+OZuKMAqTRikPDcQRmDQQuKequW5JMoaUp76ljqx4aQFg9VwN6Tm
gm3OUNmNBxM5CD8CqwbJ2AP+mnTeZ/+FlJXJN3pGfLz5TbKx+lIYA0HPxXi010OR
7FgTueXluyAfffA96w8erRf+U6tCTbd9+u2h+koSVY0xozKsNLMGLQYIAvDQ5u1M
iIwLvyfDg3R5UKdqxWlPHy2f8dtNthiON00SGpRb3bvuiF+wsKLBwaoPm3tksIn5
0bggq1ton5d3AwamhEINg3LxdNqkuUQRgNbzEtvGDpvWS1dQ7OkhT5UyGLSuP5O1
N5c7u5UX4jFiUbQePEq0tlsJ4jeQAUzQkwwqpa4FjN5v9e5XQqbSt5/UiLZEOJi+
anwi+OGBX5BPFLDJUmbnOvHcs9SfZSA7VEXmUklINVT2CA2PxZxAk+y4MvuOyXsX
g48ebqMxu9IN7Tcj3kBBarejrNwo36KFBHVyEEneeS/9txFVI2FqPnMBELcDgtsL
JMFV3nIc0Japqr9QWVn89FqotRBBcg2CeZ+0LSzUx3m8D5IXjqI7N7ScLv05w5dz
vBrjo18q0j20TtDkanCydGDGNMHVyjCPWdU6CcKfmeBQjmiyEXGmdwnyAs7vkq7N
pmpY2XR0cKdaL/outfySLZ/3wQdOfVOcV/Q1bO3oxBTOdz0/o3td2Bs+eREFPJ84
fcbrGZUlHELtLxPmg6gUI6KIalQuq5ekJ/NP9gA/8kkHxe1gNmWPZP/2yGSyqlhr
j4kZlGXt0YsVaVEHMJVkodudMT9MJy/hwChuFJvy8V+H/2HlTJbAhzF0czygwAmj
BEW4iPRw1OAZAgadopndHv+6yhBFL81D454DM9dQtdnggJIyX/qDP5XcqXOrpm0y
ZVpWKUdxM+E690jvr3tcSvxOpzCLOWi13ae4EbmVbwZ49aurI1YNSXBkwpyjXMfT
bEv/7Tgg+a6z5t+M98PiEIoyfLphh/DLq8Ew4EMS14O/8auFcVSr3lyz0PhFe3+U
vJC358y1lZPXzlEnbodWTWem5xRIK+ZqaHpPDrLPXsangpOBJkEDmHgxXb7GljxW
a+adb5E1fCS0HYRLtYrtUjddDN7Grz6+APQhDRJo4YBuDrpqZuTy8BtlhuO0NzJ7
0oKixk58a1H+a0OJtWkVPGqWUqBD1nJE8rQHAMsjdQeAa/cOu79dEALN7zNWdko9
R4FxLpqxKs8IIV/QvpWk+sqS+CFEeZuyVh9S2CjRikhXPlAosObgui9iOAcsK2Bi
HTqfD6/tonVCyMGteo5uf49onJHU0amyxB0sO0a2UceudGi7SP12eRLHil3pTUXb
jXybY4jPLzNEbCIY90VRWLR+qJmGalGc7r6Ar/mYJuSHkZttLJtx3HDAe1u0aZY0
x4VgLYdOaYi0L6z9I7XZowQdwieZii2Z54VP9Nt340sCDqNed31Xjx9WaoKlchJ/
M9YVyV9v9G5ih+SEHE3EsX6Wf6gIFeIbW8Kq+fYW9BW38PrkaTsNip3MZZA4DReV
Jd/siZet4ivCiAFFKupUFSRygixMUyuURKlshts26vIgL0/RD6VVKxZKN1RFSNYG
2tU054bKO8z6sYbi+a1237axay438xuYdKMidcYmE0wUCcJjzVJswt/YvpVnVrvq
+OsfZ2vxXNzGKM8frLSmQucbICXI0trj9/OwaxLThVwUpF2/6qK2ynzh9Vb08Vqw
2SM8NbF8RWIJJgDRjfQ55F+JT5/favKkCXnFFmwXOmUg7C6QjIUj//ziQHkYNEmy
hT7zwb2XMiS+webDSCUgbYejDti6LG2kFUwIpNjpPSmNWJEzK6ZJYMduRvT//H19
xfbA2goQqeyVBachpinugu7+PO5m76Fa31okY3/lR4cWmv3rIsxACW91/WJWR2Ev
OH6SM213y3msk3T/wfJam66aX/6/rMp4Idyz+DclkXy4coXysL4MX1i5TXY67gzm
u7I4lY5pZ9c9fMCxq1NKb+s/BwuFWJ8/LQRiFAapN/++UoAjf8WCzDXupgUYWaxu
Acf58BuC2yoO6aBQhQpMO3qzJ6ABdvjXGTPVmRHQBv1mp2T2rLno77Cy5YdsrBCU
PydjCFQ4+RmfNxVgKulTPVtId3wr/NvaYCSi66PChhybhOoNbueGiGqEKZpRqwGw
15xl2BWriSiqAmJRGl9qrvB7Kq/TXOoW5nzOy9aVeksiOP0qXZFes0uU/3YXp/oL
dGgAXpZQBYwF0LfhKnvsh3FeCpa9RuVd1J0a8XWKz0CfaLU4vtyvYPP8+Vu8s4uH
QG/gHECSNnrI2Jw3TMs95C5qlSVWsLR8FqrioLfE/d3jCc4dtMd3W/IzV3LSSNW+
LXVZgHtZKTdZ+1Rre3NO+Iinfb1m5mwbV31nv2BeIsrgeF78nZ989Xh82XP1QyJQ
JUSyIgu0TfDIclBKS64wd2nUdEoK6b0EzC86IK0VF2Pfo2FMG6x8JpcIzxdXicyV
yL4CEvo42qfrZEfp5Mba6Vk8OIO/MGaB+LFaho7tOCX5nKyMEphnsVskJEju9vgK
TVYl75LOyaKwIbRM3ZV+J4mafI4vV/JlPfxYKg569PIovB3cleNYwvpQkUpxU3bF
2c71nQabFJe0x9TXvebYjZC0azIudRgDU7NVl+S83QMvt6/7sasE/vhDuYhGQBwn
nK62tvtBzTGfBmexkeyi4MbFI9RFIxfCAjijCBelf9/G+krSAk6XqRPfyw/76WF7
xO29OOevod7WBqP4q1bUOxVOwvLXxRvvTggyZh3Uk4FFGTh9gDF7t2iwHMVLzeWN
tO5TQCsDRK9Z1H49xEFSNuZlJdzPYQsaspPwan5TQ20ncqUViOEtcVVeLgLrByqx
0P85mtAbmKyORUmHnAR0eNWNbF1g8P/7K9Z2FtBXD1MaIA8d1devke5X7Fv8uHLU
9GUfUvuTngDkURmdMDqisyV09my9qUYqDPBBVZBpk1+usVgQuffebisPS+KFNnkB
kR+6S/PJ+55702HfLAyb7mbViYnMl4i/XQvfHvNU0xMi084R4dixkEmvyqIzr9if
lYxDWntytn9JfyJ+4R3PUP1Ud+xgmU6REQaZ7ZRAMKjQ3CT4vP5M75qblhHEELNo
oNsGjdpTbUfKW+cpqDWQoKXWRkqsdEsvwFvq5rY98QCtWuD5i7Cje5aenmhwdmVm
9D2k6AXgegXchuDx1NInYh+lOAbbTrN512pXYnncQGM1u2vly3KbdkabMDizf0ad
rkOOzwh+NeArlExWeQt93FmBLvXXH+h40xs7EUHwlLji1IW4CDpIWy+Z/nt7HVrF
7j5vA6KHsFDAlQw060z5lwawehNCuk0EsV/w8HIaI7uAT9Bpl7E/hIL+Na3vnH9h
edlz2cYgTjzF3Ezrmuy6YGtzq9oSHYfjS0KC1JDAopSdlfMlWfXsCW4Pc7i1OgpC
j7+5z++Y0qyGpkUeGq+U9dIHfGYpDjXFrGdEmghi5QyupsRlfk21bkHCafIHn5li
/8MFmRUrbCq01sl/s5aUnE3Si0RiCAhk9APrHDRcr23LNQS7iNmD+C5914jAOXtd
QwtBwY9tEQb5cKe/gotYfOyoN0BWtCEtqHJkdwAsxoYlD/TiBxsxx5xsmDlL9Ti0
brIvhRG/vO8fIs5kzhHASiu8ZVbaLzj/kCm6Hg1kTfWjxX5qRx8+6l8XL1Tr7e/V
AHNv494sU40RWaGT79yyI04ObR77+gOP9d7w4LN1VcS/HzbZHu+tEx17gybIDRyg
mOLjRwTQDZ5Rlk7fC0kvfThO+KF0Fr0x7ANCRryL534ykThSNU5KwAj2oglcUghS
vEToNwmv539cS/ttLFA2VlJgnrX5fAMvTP0gjUpU/o33strzxgaQM+D6pfw4v3bt
oqLmAPoiX7a1mXkmtLxHHCF99WOI5kW1gEY4gNRtntpBCGWoX9uYZmpRokzzX3zG
j5CwMuOqfai0gfv5GgwfKItJBARMj2q5WbJy2nUf6w24MaNvXhw0l4n7YQ5/vtM1
2WXIRZr7dPJQqUApwzei7nqdIS5SYm0EnRLsbQ+TpB18mY3VKIZB7VRa3xZj8o4f
b6s4p0lTtxanT6O3bzXmuB7w8KHQMapI4jNZx0PcF/bmJewSS7HCHvXMMYsxiJEe
JI8l4eQLoc2SzmXeMi2hgeRuvsTylzeDcQwy3beUc6e9M7Z9BS6wUUYj4iukE52I
KS58rcD0ej6rWgxdRHCja5LoqCxO5/amvRvyqOWaT2BQKXs2j9vRuW8tfggaUMau
veunGfF6k4/zxO8ThlWl193sSRTFq3jj3XfhhsuRsEFskrIiLf6K++BXtXO14Sj+
ISu3KLsRW/QtbxAwvpMVBiKe+LEfWJf7hDuJirU21dZOQuCJIpXOOD0EIJ3ZPl1d
AqAHZW/6ps6z9tHfF0xiKjkjxCHhhk7Y/iK80w7tGymTj7e5Bc3zGHghO6D/8g1Z
SNOl/9gBel3o1wPjkrHfmYdeSUdcsIIODXuq7kKbcZtO9aCOa9CXo5HrKB6wqDs8
dFWZm0Df9D+fKNaUPbxbr7zqfZINAxhqznNnkBW0Euq+d2eyXd15UU+++IRtA9Ah
/4uvoz8iu8L7xtHqOpznA7HFsVYxbcVUYAfJsLBUdTYzjteLW1lQ4/SJyqqj8qlw
FjlOyKDs9EbFGs7Vhhsyr0laudQK293XPTyR+eoAIqcg9xvDJac97jaZRM6TvNNi
7ZRJ/MMz9ISyiO/23/xkxtenGAIBHyCC4RJb2EVMxvtoi+Mzj7xU80iQFPfszFHh
Mcmdf+uZawozC8ear6WwXeH+762RViMA6+nzqsOjHYqXF1izB8yQP5/FYAQhuoDr
T3MavAxXusBKxp5PFbg5b6/LEvTGXcjeXX8U5nH9uj79qLb+pVKZz3uJcRr3jTLd
wb8FYUM32bqqYaxBmA7UZHsuEesAvRxkmi0/MVhZCFUYEbqKze9LbkCKSGjCGubR
u35MH+d2OW6OYwWn+0MgT2oS5u6rj6Y5VMCbhx3otoT/jtg2jJHBDgQDQNyoaM+s
INHs9mQtsnxrfHCOtof6guJTvXoDdYGG8bPUtkFoOffzMk/H4ThLomrta0bNzznG
peXU/Ydr0XAywud688pip/ci64YTD9+dHniaqUVTBA68vE6rM5MztBHvLJuCQiZ4
QwEB93mxFRbHFNBbDpTaom60zaMIhVWrrbw3+1hehwUlZFoQX+t+Ie3DWHjheiCQ
HoXP0Ii7hi1ctAom9bfNV17mSqCKEVqy6my7W0/uOalg43FxWtYpq9C7T6gJDKUu
yFXR3JJppBDrdJaAI5u7xHdPrN7fyHNKjg1rN8n3Lkd/LfGSSFY4DF+pJOFQ2K9l
/i6KxYRQEGfIu7SAxus1EHVeGRCm97ABSq+GVAaYv3BEMq58QBb/2Sg8DlVRUvlb
RyUec7bR6voarF1lSPc1wsB3hHj/Y9EtC/PfPCRo2EKrW/jw3aBDLpI7jRvrRKz+
RYYG+Wd6dk3/o7v4ESC/6R9XptC2+AvsnbOeuMBMM/ETqTi2t+MQe/W+cqxX+tuI
jerwYVE9jfhKaGwsG1jOfUXs4qLrk8onD1bEuU+AhGBtS50DNhyYnkHG3s2oojuz
pDV5OZXrZDQfCGaJY6676ZvTBUgZZ0jtq7gK/BdOHPFOebRIqFvFJ3Pgt0dNj3oK
Tu27ehv9P8fdXnY0LjX8Rt7mDUfPqTWXB3IR6sR2IeksL4tM6B3NBOM7pWZ96VdD
rxlPKuqoR1G+omzAs6RUs8N+E5iNxh1NGisPz2fRCJz7IWm+d3Mx9Lo7I2iEf94/
eJA5qh1eZyLqqGNFhD0K4yMProlo1HiVdaDNSjGj4GWQ8lK+YFsU4vpPnQXHCg2f
Xr2PcSqxOuGdQB1cq2LAbNCpsaeG+mdwLNk0KyZjBAVDERxql2TMiGdsbSPD8a6D
HDafIKIl9/gdAc+XI2/t7/j+7JainOTnnS36r5oa32m8fizaKv+3rMpRALmbIliy
SQh+AsNLwJtZMG9Hnhzr65vVESnzJamd1h388kR4Qv3Jh10Q7hJoCSfgonqpj7lM
hIXm9mrJ7GxBdJ7FE0amK9XgRG4snT7CfsHTglAOyH/0wv22F/y/pgC4Vjk2uvcR
nGDFXLXGRqpxdTiINELNzrRRCnbzRrhVGG8b61XC+pO7cgUMmTSyDTjRBsFnOpkQ
z5KDguj0AqFSe0KVnWmaZVxZ6QMPAIohYYoCaj83FfLSRwKkSM5pf8Wm4HF8YmDW
cpsQWTEBECFCJ7QCAOS+2FKFDhnVI/S+d10h8k0ss3rN5r0AMvZR+P2Qb0ncFmwy
jWzt07UvXTHujFg+x3vTMxLBRz7vdFCQbizKUHq+Fmeuj7WH+V4mv7AaHONsRbiV
6NEJVBilGBpj1sjXGi3djJ4fXXQGkKh11fYanFuOcHezg3ln5CQLMLn4UGidWHLN
QtrsghEheoXn+HKbpXR2/davBVsvriIgCoTDScBU8HJ+49r1O86mga7KtjgClVvA
uqlL/oFV4gwIjJ1vIU3hW7dFvtk+5AG7PQlUZu8fYFfSCpF6ch5hL6lJh4zsavIn
B9ck95HfPZS0q/x/zlJua3ctaixExEC1Tqi6J7Zi8Ex4BIDc07YwOgdkPK1xHmea
vfqtsNBOY0vSPJEAfh66su26jxzJNQbc40spL2wL76sTaTWz5wwu8oRQ3pHlPR6l
yI/qBB9msIrHtWxeotFj/h14OgJd2wRSq2c75y8WgryZWStkxZuS9SrREmDuE6w2
pwKnj/Yh1kTo14IFVNz1SLc/+wYTvry+pI2DcEQTaHWhzg46hEWbOFB0Qfa2xlmv
dYe/tP2phkBPXcRWPx6uPEMDFcndl/cyDYj3XKegP1ocqRLLx2yI6Pcw7eRKimbn
1TMI9QbN/4zs3VCWQ7ddjh9MSWKcuVyBBgkk020i8c5ghN9ELPvUuSYFboD42hMy
uOib1W7JNn4zUGAFy3FsdGT0qHdfBqYNABN3vEbGFQlcEjRqE02zmTvvxJ2BD2Sw
rh7lWVO5xz0EO6glgdq6E0rqQ8Op1rJlxT8FuUmi+w9KlV4b3lFIkIKWwKvU/N+f
4Baw2jomobNVC2koVwCsRSuUUv1v8BjC/FTLy4QzV9RWE09Jbq48KyyyxA/86BEG
825E3PfXqZaCkmKdrEWmdBYScabn7F7z2vSeqgZrrgvQytQmmYh8qegw8QI7wab0
Wnw6iBcMhDxY4+mzmMRJoZclCPOUHaOKbjORH2A7N4FLyiwS8EQEQRWFQlundTIi
Vo+qDCBpc4yQlEZFzk2YsODG7HL6N3svqq/3iL2oqmySyfq2+XJ/aWAr7VHb/Tow
o0i9IiyrokSbZHxlRk3ebiBSP+nGx6lHG5eDSmLHjP/+u8cySkkHCprHAZ8SdmB6
J66Y6nvmctPPSC61lYbVfaakyLpZ0UzNAueCjqyFo1KPFzNhNE8AVKrey1mtignv
ApjNgtipyY5Gy+ycHI9pyT2KgtkGT+Enxa2uT4nnlbk1hHtdXplcIA0hE+HytVio
9oYntgmA1Q9+tGRIZQFoNVcepDbclrs4FhIPYdtKAo3SG/m3Nbp0YVJjzoASTZGB
OpOX5CazrXXp+RhGIhjfeNme9mKkPg0X3z7G4ROx5FLmYNs0zukMM5/RZefk0/sb
Y+4EOdYIjsx7wOdiCTcwZWIPxwYL6dOFm0+IIe0zc++s5bxyo733CnLq/x/9Lp35
LsGZ82qqRRr2NtjS5mbQ7azrcbG3rTixiSBhMvdmRM9w2q0RKNrsC3XjTmD70c+h
AubpXg90UsCuQWgpmjBfdJ9yPiJ8HzoaGyQhZRiZz0mTtetxIFddJ5r7YjCZc94/
TyxlzX9MAnP4J2fmJwoidMkyy3Nzy/6wFJZB9qKngJLVDPTbK2N9/QjkCaBigQv7
Fdu+TZG0RtQviX1m6Xt0oGeMbZv7vs8R8/qzk/uBfcxJTG3eaWKTIt9pzuASb3ci
9eOdwlbuAX09GkDN2oxqf8xxuhixkug71VvRUxMiP+jA2OerR0wY3MBc3wPsE6vW
wMtfCAUG3DF1vN/5H0XYM08owpGs9sgqbMg5uZyzqaWu2USQOYLaY229GKkX5wGk
qAWa+3tMOfn8k48SDLh0KLXIA3zTkxYMiECGLhKPqURPdAi6Nq/lLkUaDkIX+X2X
Fua+quXViKmSSGGkUjpZZvPVRFwa60eHSLFBryo74n9Rw/xVNCPrRxDJY5vWqymk
2MJdlXM9hBnL5C6wZ7ocv2yRiOWe4N6vGnqdvqM4o1DMsSEjzKqRWi8VNG3cMwT0
RtaawGhGC0cdW2M/O1KjeJRJbvBthTihWarikho59IdeOkOdH1UPqsWZ8yN1jVFY
YtkHrbLK0LP/4ilNgA2t8KYn+bz7r74EVdr+3Q/rlFvHtzfklfLLrLm0BYU96DZs
kAnkv7oe/kTwGiJ0fNeFHYSzhrLY2erRfRMUc+wio0hfP5HayHx14ViDDiVQMmsX
k96G5U4bB58/EaP14iOq0kiRvUK+Fg/fNN8KBcehjbCz10sO1dqganjbr17PFXxn
Ve6HX0a5N9JMkKj3zd5LCacQVNisABngykw2OZZMBnaS6vcIQBnn2Neg/s/Bec8o
xpVqpOxWNPHaXCB/pR8EcqQcfxsc8I2sRG4q04j3mqfoLBpqhPajCJwNZ74MsVfs
LRkcw96Izxy5ksN3de8yd+RmxDXykh8Ln8QisJshBlRQyq+ijqbZkfx9nBUMIRC0
s9bamJzzYsOycxn2jLkP/toQT0pJLzWNwEGofibSJBmx+vM/+jJdB6EFxg3wp5pc
ETePbhHIUa1sSleQllfPKih6FnFR6OJzTvFKak61mAySp85UFNMcf/0LWMhGQcyu
9zT82mZUHgBl3D5G6xlfYbEsFo5O5UQB38RfZAwFpKdF44C/dJoxdcuJiEWTmYDX
zleGjDIU8y78ACVbL5lutYXUMAA28J4qsu+nRPbDdYl49xbyasRK5evCUUyDwL35
RBAne742MXngTN4yZmX8T8L92QfYtRi4ip+OUAa+o8Baq7uYFOKXgsqNv8jozUdP
OAhhyP5jf8CvPQbgK+vGSSXmKN6FsJU6uXm/eRVoud6RmxzMnmmUaaJ9tcdM8ovs
isFbLeCv3MHeSN+r2dZcPXGVCnhGxrN/oHx+rxanGt8F6FWdzTOxaJ30CPfLDX2L
12tlk+/XPzzHyXmBV+1UUQJ4JaWWYZtW2xqGK/8fnSnUWQgQ043H3JIUNZH6qzTe
/5X2Y1Hn/G4bNojHpFL1Tuq3LohrVJ+4zGt063hPmeweglMaEbD1+EGzYDVF47BQ
WE/xo7P7/+w3kYyNmwgkFRnoj6jCZ+heyKOxvndLLbDpj7mXn673/qDqsqzcAIaR
7mB3vzutV1htwUb6Vn1e1K25+PaC3+sn1U/RGkWMcQlLoMA2jhERgWda08NqTkqW
76Ji6xyt3a39mTLTDZSoFIeRs5hFdYe0/ar/WUVcYvkZ2yomNIgJbsl+mG0qjS5g
5HsocrR8drap2GcYlCnXBEOyi5twRDjFrQtI4S1to2GQETecGScT4Vu2FsHrQitC
E0ZConWCmCJ7keQov3obtTBLGAWGOFlMP+pODD4NzrqpxPOjOpPA0i8yDgy9Fz0v
RZzgjvEwP/WFtbl/ek49qJS1nRHKsBVjtDBmk7dE4hZX2tdFs1JcukTHY1mP1HXq
yFiu9raP2rNifz50yRTSIrV4asX8SGNI24vj6AmnuIHQyo6DOd3QH1bt77mYoQzJ
mxRPV3fcpimlbMgt68eNJppjgUkAk/LTceEwxxSQa3cKcH9oK8IFXCul5ht7gajj
m4sctlU8wWUZ/sNjeqba5GSBl6y/0Hv5KcjpukpSEqcNhjWwa/nb1HXBaj3fkR9Z
r9txN49/5veuAuIt5LgDk1Exg0W+rljEzVDDwBA+voBi4qkBLgF55vfXxkkHl6iU
7VaF22kRPZRfZq+rOaMf9Q==
`pragma protect end_protected
