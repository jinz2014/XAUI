// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pbkm/C5swxPcVVhaUqvW8EpJR3B+EHg77EXY0GmLfMIwAeKt/Ixue7zi5ALWPsI7
LdRGG3bE7Hw7TatS8rzBVUCNsR3o3b5YJOVQIm3J57kvnMGs4oL7taD5fUkfoU5c
IrkIiIngbTOa5AxLpWMV1H/F46uuJLrg23Rx9Itzda8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18144)
jyDLfH3aa3oyR5OkCPu7zkdYankdVOKBjYE+yCLqy6vrCqv0uuHgNTm0ZWESOENA
VxQG/mwSE/yymGS+ovv7FTD1vo4wcVc2hwoE5qWZ8K08fbnfcN66P/SGVRHs9kgM
lm12woYGGFjBQRlW4kyPfGRluPn1maQ/nabiAERJsQwyzW8epitAxMcbzEO3dgKp
okRFeRfZqaGC+rcMtGOgtzDJWY2cLST3O6TDkThtPWmTg4dVJLNnxULDVkHooCui
MneRkXJZY9FLOi/7rIMZ2QiFV8QwpAKpctzn5ejU0CJvHDq5lGztHDg9gVVjBdff
3kzB24Ny4wAVSPkGFNnZrpdHcbz6+ieB9oRkWJaYVK8orPWgpVr1HDxWsVgivKlf
gqlQ//Gv7nSZnw3NoXs4ftEdS2QCs60UZtkBuKtnmEcAiJ0bIp13OXlKCqPzVjVH
sAxMCJ2Oci6Uvq7dfpMpDRZNpB7CPhZQHIbRttARyB4ingUnaov1eaqZGx/IUu6I
xxI43+4gwAsLHVDRJn+8beUbme3LZoMlbQY+LWXFDGaIMoIYIp3qj53TPlEGI8U1
pqpHhgY47uSgFFyphFdpzzvUjcDiitmA2lCAUcKCCljFADtw3MFzqAK2XW/uC2Ls
GrTNIYrlepoCbNdI4PmsGesV805NOVuCFpwDloy7/ZmFK6eOhTr73NggQCjjwPLm
tvWQV1bHwlQ9R9jHPpZpUNUk0RYZIzkpAHAqNRQUdDTRLj4s4bIQiDXkclzSb8GM
B8G1mCP1FKANhEl9O+RzT8FjzuePQEYk7e41UQTqbA/prN1AOWYSrcWTcsQCrwhA
Ksk3sjT1BbMJ9tMMAYazed5Vb5I4/3qAHA8Dgx/DRe09UjPCMRsOQMrITfkv4Kyb
U3/6rtzHlCtobqeRxFuTaLY2I1emtlKft0beRZy93api62CT6E4wN9pcCUI07aQQ
LAB71m0woPzOyC8AKYRfPWgGPI7tdi00SnRcxlBsScst7Gxm0WbggZ0yzrgYelZH
W/UrUUiI2GfzyMXPPtXx/D2UAOCJcuMTuacba7uueMnXirIazG9yIuuc/McAvYKa
R3jU9xNUEEk93cvWEZg//A9JntbrfzeTgSwRbwBD4CYvw+oJIZpwPiReeHC764L/
dFu9zsOzw661ByDttdYHGofSbYQAML53ID4kO8ZyhVaH0Nkdz2UWsx0Paury+eKY
C/nlmz84hJnxpOTHziRLkKk5RF43DJuPPgh9i/4dWnxfFNDgyBag+gT3qJ3Pz/mJ
LmS+/iZupTDF7RpmxwJou2+dwukjxn6+azQfo9iRVMAm8mVrUIRh5p7QtX0qyc7v
BTLMw4Iw/4/cJSsz5ro8iCrurzSXBBc3It9hsnUmmJpYEmBGdvM8SJwuR4ZtqaTJ
fbzyMw7jOtkzVfkv7nXKJVmmQRChbn5yGPbV97AFsPeBQZa+g4nZSN2JF5fD98y1
u3SdYeb8w/Mm/RbS5Bn8FB5kZMZSnP7elS4b0pYmGGAciNYGSILlru2IFZHY8cW3
Qx3akIMrrokCDDRoov1ONGIMTYl/pBI1t4Ctyhdwno/zWznaM9KxWNDWtWs9lk9j
JsfJbzIqPJBeHEVrS9M6HUxGopbWPHbUcDCSrxECIjCcLMSuwusm8J7iE+xe7mst
DK4kZru+WcTzhY4RSS7bGUt0vDiymeHxe89HM2K4EM3yLlHW3TbTBFrZ0eE2drT2
/9JclXmHvm6YVBgkhczPAMIVd+bukAxF8KH0G062Yf67wlphZtA9HSSsBk7rYOga
0aCKL6Y0iKXTe8GvVmvyqmaesp0LT5rlJrGEYrC6ZgNv6AIbNA6FDP5U1nsrf/XZ
wQAlaqTUuOvMy4sLmlIoFyG3c8Um5rleSD3QIgHhIPAeD3OBerMJtZiRMYUvvZ6J
Il5SQI/NHyio+VNmt7pw1Jpoz7bjbA+SMjnhR3yXWNRNKsuwjtAmUOWlU7Fs8THN
ts2IHkJTK9UO+8SQHXttFrtUr2WcJpbxTKNotaaMysftxS1FmbDTvcpEkdleK/Pe
O+voSUcSraJc3xtfQ9g4I4eAjTLU3i9BwqEHbB6VjWuSEodqrBw3ZhMIdXUzF80L
qFpvAx7TxqDemuBn/FOTeqK31bYRWhYFQ7vDzEy2xMBz7kEYfv0qb70H1EqghwDd
sIhdcpRCZhcDR+CtomSUK0HJ19HkeIv+ZiC2yQZXvjKIpJmBSUihMsNnhfJXYIEk
V1DEZPZ41dSAcWZ+LEdssYLrZ0kVkzY97yE+dSXR90RIhtvJtarLlEYXELco1a9C
KflwVzdPH8QRKAluRzI/su2RBVnp2Ry04OISST2VsMxlw5w+jc4D5ZrectK9oCYY
OzHFDvRdev0tt7saGej29s3vD+UGBPDrAImE6jnlqMs1JzPyLNX/VBUEFJh2WEOu
79YPs/4vtgGxIReepzwMG6/SKwoiaUYo69c0t8ufpAv5r+pgxYPRKIMzHgZFhivg
YMfyiRUjf+137Ft/h+jomD9jUEZrjaKrQZIGxJwEGGg/6m3tRsUdyS14Zrxz3WMm
2NojgHSDlCEvP8zUr1/eknquEizvXNTG9mEV3Em8BiKsoMzAt9ZSG8WKJ2z5ytFk
TE7xSm3V5yUXX6z1BDjfl9GzYqOtgmyx+mpZPENJDOxbKt7fj5PjXMXYy6R+whQC
+EIxX2W7vYEa+VUg7RU4EJ83wclHCWUmo7Paxgp1PU1yMLOdfHQnTtWSXUzREg+4
r3RmTWo64A9esVabtvXEQQ0lJv1SeikCDO5e7wYmzD2kR4pfqvepJ7tzQZoGK8uV
6hb5iGegE8jlEIkwUsrOJwFfSXTyRoy2xcohmsPF9Sf9Hl99mCc+yzVZCvWslEwL
hVmsEFgbpd4Paf9M1ia6m3Gy6BtvK7wivqs2k3S/IL64BYg4XbR5l2TsfdSLk03g
Ty+bBsNsOpCmUG72roSdBNVMmpN48w/PBArY/I52pHf35Yt925IxXRbAwLiuw0eh
OpZbSXmxs/XBRQYj/p9wylG1NuMxgGL30h0PC6tt1H+GcH09x+/5xfsB/ThAR1YZ
Ndc/L/7VZ5oGHEgR3oxnef7CUYzdjWgwUkMRywJAhXDLVVQ08bGYLh9GW88eTZ0x
JlQFg7P1wZkzvHhdSrLPetzvwszEVCOl0mPpAI1uitZ1LDbQ37QFnZfcblsw9j0O
eIeMVo5ORp18vvaFpNjOtsfc2V5PuXQgegwZuQqjLjRsiN5OlqDOEyBAIendmIsJ
Mh6PExziwPBwrNmKl7SCp5WiLtsYPlbBuAF+XsAU5c4mK4UcRsLXsgGS1GqnTzkV
K0PxD7mQ9l7XHr2W/6B76b/jaOFUnEW23yig8iaNGTT7UdoHnz4RKzFhbI4At6Kq
vib92/miTKUTLbLKzlD+EbWx1pn3hlJEeI9aYDQaStTsR+V2X41/4K3oLyG1BsCc
LpNwKf7h0DBB7GRXiyG9kJ9/UrmP2qRDTnA7FqvYB7zpgUXfyn82rIIeCK7qXtSE
g3lkUo3RT8w4FcMZEh5vudQyk8q6hagYeobiiifH/cCQOmkvH48sCrMBqm0FGXIl
oN0ig0jmSkpmDRqRHupYisZaHT1yDAsRnSKhqOIcDgubxb6X7AP14oZIeh5EVYH9
kW68ryXArpIegzg0IR25IxzlHUDeidMn81ucf94O9zktO1c5okt1wvJ/VKkimOCg
CDJhhSGYwV7jqpI1gKe98uXCL446aA//oA8W610mgxPaJrKc1j3aWJrLirSp4Ba1
3veuQ3Bai9FBFYPuFnlqY08buUSylVWabrVeTQp3bMhYWC+9GazI5krX7rCNVSU9
E3N3g1UNhw5hzV2rNGm+5xZPdSG0gw7CGURXlL/71pVNodBZ9FEOc4mlOfS96Np0
tgB6wY6n2SlrByB5pZxlqeTTjMz4Zzhux3YHNUlQLvBALbCsuOvnMcKnYVPoykU2
IqaHb08luEUnslN21ey6AmE9zI54nRhej+AA+fxt71850dWinbmXo3Wkm6YL/DiW
0pYC4LZZM1BQ+GBwqx4LyJtvfNq+DrlVJUw+pSM/2RnnUXmdvollmXqncHyveokr
R3B8u3s4xNdVZVMGIE6KOXFnVpTrEqKtSjnjPlU59lXy0SyzFoM5PzPjwalOSGEj
8C8db4ZJWt5WLScJ+mftYc/EtvNx6/Fiz7WhBK0RecLwKXRnKO0toqIdbTvPl3jH
SHDjZqPEV/Y0WfpWG8btVLz6M+3aZnHFcap1XyXzg+vy/wTqqDBgRftOYFUOJCL3
5RwL92iku1UE3Xz3rnY46ef5+Gg6cqboTBflC8M5zyhoAtrzFaNX6aVNojE2HEHz
Dmw+nsZfWAmvPkSjXKEddsdkbpJOm+6k0h8aYvlxJJOAivavuPJOBzmakNExJepY
hN+l0tGz4rHT6gSFrS5WADVWbjxlHT1D8mvTLjCihuGBYsPbRjNnEiHf+QMhNr38
VwUR3WcbutDgC9bGgHVjtx9NEedRXn4BMx4ZzIAS3ZxgYWOdHZovCNV0+buIJuNZ
vds/yNGrTXzur/lULUn3eXYAb9SlMAWt/TXxXMB94ZzQA57QqdkM0485QZmeogGm
UW3g8ineJJ3MOT6jhGo2hqqhs4p4X0Pwger9+ASrRRLDErrU8dTEPk8kcBORs0Va
C+VFC+nzV//zEyOyYl5+O23zMuiUwCw6Xk/taI860LGq/xrQt2/BTkiplXL+lrL1
6DSfE555FMmGrvERJ6yu+5G0KfHns1iHc0oUiRECKa00nCB257QR7epR8qqoSm2A
IhsNsc6BvyMgPfYL+kUtdh/9cQ+6SlSDjeja0u57x1CiXbtG5D5lOKqdARWT1zTi
uRYcLsywcUEEsLeT+cUQbBsImLAk7UydKhOXSV45ATT5II/VPH+FYSEyOc9hIvii
Kf2RRz+b71MjHwvuaySoEfJ4zgLp4WeWf6eP7butMPYuVWvJDDrFThtMMMlWjatz
NzFSDKLTNIgBfBKTDn6qDvSUV7fssH5FnfmgDi5O7/Cv8SS7vk+HtmPbdRZRj61+
6Iupi4SGLLEN4sXKwXJiAKM0pKT7vrsocxQAkXSSVAUHNH3jM94ZSTJVlomJx9FZ
86ZTGNc8b3KmwK2OWaa1cWze0GbnfdpsCpFKM6GKJ+HoyJCrUjPVHqcffvsqdbuD
C7+htYMuA2K2lktKdBU2OStoVbtlbPGC9+A39jD6xENW4SEAnVyOENBqatNVdNBw
hUxBs8e6RAd6C0Obd892rIMrn7UqexhkUxFuTtaBS+nwdVzf5nOlmP9Kuv4D+u98
hh2C+iRQ+3S3rf3okZ62OAzJVx/AAZX0PaSGjPyxpF4CleM6aUN6jUxiVRNlVrtm
MVoB3f5M6454EtiP4BC+DZEC5ICX+MbugTWruDUtvJveJodXoRxVH7mAMTNhVlVj
UCnMwYG6ANxVsyH0hTG6JrwKvswHCmoLGEZ8JdQvJ0ukYZAcFe5J6Jlq99aDQj5G
myP2/PPMPGjESn0eAasCddqjocZfJ5G2498W7urEz54XQTHcqO5dgTGHPD+AhRas
xgEh9XEbwvqJsm6rGSTPk6uM7ISfRKAZzbbfmu1ZxqRJ5pJT8uqZ7MGb7dVhn10r
FhNJ4DHgtxPUYDbp5qQhypoMe2Ja5bATLNjqAb319UAmA41vRyrwLp2Sazely5KY
P//rlUCgOgf701r9J/uDLfzQb0YVlI2RqgbM8e72DyuoxCTex6BguX6O6WCrWo/P
PjKbsQS4Cnb46LsSJVxLhuqqx54cA/iupQbR0uctbimP8qxxAgvsSmjZ8gVVFd4q
WT/eFWQEFsiI5VGuDFsI34Dmw3UkjBlTx8sveL2GwsA5tuZvfMFrEJScKX0m7qom
e5sW0sgvum1yieM2L2gVuknNIHuLEadXUeLvOqo2U0OTkay+j3fqMPkMkFZdIHfl
yGEs4qdIRgtaBZ9lSYkBxQknO6mTwZ1N53Tb8VwBtaSN3OsPPgUJvt0eA/mDxB7G
tcj14dc4B9HDttvKWFcztpJorqlN9j3dcZSNJct/EfXKfckyr6EIT6tjczSpJYej
iuFj62tbuSOBsOysXn0HC4Rvs+MrK+dOLloMmyh9cDeveq+S98uifxIGlq4ow2gh
e5FuKzmrkku4P/116U508dtl+2JcTcguqlNBzBNrsiOuTdU9MJ9rEc2OfFcc23Rp
aYySxTus2WJiEUA5Nw8Dv/UliTyQBZ5uZE/F87jmDE6FvcMZSumfFTUf9pTeErSy
LnFHa9j7MXTPUms1If+b9nG3E9/XYXNkJtoPvugLbwivyGB2tOtfjunPi3DLefGi
S7zMuyfBCniBBjqN2Ku65sYkJHkSPi9XGREFyJ2ZRoUSPY0HswFcCAMcQhgY7BLp
qLg2WevSWoUR7nLI1KAbBrqbOkzQwak0NqD36J9ud0PVQWjerUbQ+sgUyrSSYDWU
qoUfA46wUBfiDAcAKmFtT/Rnse81XKzs2s7/hsRXpzxQYhexnWZZ5ywPoAAyoBhG
3VyNiXBqLAeBJYJjR8TnIiyoXe/X2mpXoUa1bEyLUX2hub0SImYsLC5jqoyBi8Wp
pnQOxDbUIehWNj/SDLX1ybUpJ+hNMPppNYzW6kRylcgERNx7ogEp8pJPIIZ2uSuB
fjBzv0s4vxpreHOGXAaquWijeCijFvg/8otLvZH2UyeOpuj9Jd9nIN9o4C9LfMT1
uqknr9PgnvpmshKEGcRP7Gr8fsBGOQsgLvv/MFOHtEAKShUOHFxzQVQOA+eFyYiu
QuSSbo/rKmeXGVsCZDDSrEgnW/psqH3nsRq6Shvo2dF07nJeUqMANaKg4RbrxPPY
8DVAFC//iMLY7UpCRDkdjGFwsca600ZBS5t7C/gLUisaQymMrGDQTq0lc3GakX0I
FQMvrWcwbQzLHraw7ClI2fUkERa1aQ6+5hrcbBziaMuDlDK8gvpR7iouQ1C0B+Z0
YF3TfbZbfVSUfSRFDcPPfzVcNrQKU84wLhKClXAUDAIZBC/Gaw1AvtQDhr1VU3Tw
7c2YfFDMDv2E2j0Po26VhX/sA7ofGCUvJJ31rcZUWAP0jjG46uVRFFQTz+UJ9/JW
aZhiQqUynJImd/5V3nCNXldaCdWkqmIQ2/hUge3Mpmd07TPgLj7aCd6Atom7+0B5
Qo4AY1EtSWDfsswC/1kzbWkiBCebHxjhmtXH8kx1i1WEm8WBLzL6VfrpwYRGSfYN
bwvw5WSEuLlDBkHDuyW8o9v9jSB+L181Ebc3LkA2nV4/cIF5DtxkMZ2w9+hvRtQ6
Ud4NNV5yZsu3rlGPcD1M24J5RnjDqXczzBgGxAvnrXe4PgSsPVzdXq831ivC5xue
W0a9mq7oT9FO/dctP0LYw3lMBn6J6Q2IdWvRJ1AXNO6WOufi4/HYz7q0TH+qNf6N
SmrBFBZKm6AuoTXqHbpLq95TwC6sWLqhn1FwogoHLDRLgbyrU/AwaALJOBFesUg3
qEsUqd1jjXscn5U5GHL7j6/B2IIriETAm1/znKOy6KGgrnxi8oLlzHxg/N9DxI64
BmDPvxyufcxGMzjjTzoPINv6TXA9XDqu05sObkm93ay+pvpwN7YZ8t++UNfL6aJj
I8WpV/AX7vllZV6F7VkWM+yQwWE6d24jQubTYwWnho96Y9UBNS0juN9/GNYTbuSe
jEHFElJaG/+HM8+N11U52NXRSJKLAdn7uLuL9+UeqAMRMAMZet2OdKMZl5MzVDEB
JAhtR11u+QNuV/9g2ArL9Q02h1qegmWj3alxpOgc+V4Qlhh3CO7bBKX77QvWqMyx
B99Ao+bUTAM8ZWOjEqP609jz9ql7LhFmAxV3uK0RcAXPOyajS61M/d5fQrRutlpA
ObobNYabVhUH2u2Wi4pgjW17REHXeKSQTsOiDIks7hBh9QGMvjvKZMcwRK4Ki1sc
JZJxyrinT5cOLvwghPlLQ36mHlAF6pTTzWul5xnZg+lLRw/HsOCISJuuu3ZeyylO
e7ppu7xgJQk7tts4HDM0cKFs/qIBy0NqXxOoQejI5VfvWMFbx0/WMNQw9ipUPCW2
42QBJLZ4BiHog3Guh45+fe3o0VzY+DMRfTg5hWfh/eRy3diLUMfcc4S80l+B3CUJ
yKeuXY9MyolTLd9YbF+G8JpymBJ+e4PGyP3gShoWYOKGSZ9T8osqOQps6wcHgGuj
LQwGlguOVEFtTIda8I20dFAkww6iAPOH96+pnesFpPHU+YzwhRQe6P57E66f1XOm
oNNrppSHiIP7wny5Y9VbG+/ehKMHe+kGYoyNFB6LMoPdNP8Ux5L2vQCQkgU4Pc6J
wgxuwrjDwLHFEazEvD2uBT+oEY7ZSW075P7JXYabTNBbMRQsM3sCz5vkXJLF1VGq
BlVxQti98WLiHl7u8DldMOZgbUvUhWsKQ8XFytAv95WN+uehyER2nTfjI1cogLrP
c0wB88Wfaebgw7vjAWRcuAWWI0skjCNX0hca6f+viEDtdBqMkfYxo4/SpWt6CTg6
3leQVa8X/IUTV4cxEIDXA760jSDcg70aVzEjx1Leyh8wZaWmKlaQH6MPxHyA5/a8
6t/72frRCgw5eu6aClS9YyRuQKyiFvqpP4cbgqIzNlKGqgJJas/AQFXpk6hFRd1W
VSfNXKze/2MgajOeQJgsph1R6E88f/VOfuWS5nwF5A6ynry5UvRsBZD+tfNvtEsz
gmgXMznnqDORjzAdcAiVb7bwRxSRbOYWNmKZs5RhGy+xzD6p55Mbk6izByZff6Mu
bsWrsxdeQzT3oGs0VK61vn/QidS3n6D4bBQ4Z+OKmvyHkFpCGi76mqGaUNQUBm6p
UqW84b7fIZaYbuUzYpnC6Kwft3GJbqYviz6JSiS2o4rpsURFXd1ZIpi5zgZzoiHf
RSGBJWF5ueKtW0ePstHueWCgnLPn22SIzhilyDl6q6ld6cRezXiLDjbIwqcuyAi6
Eft9uPJ8uDuFIAhebpv1T2XFxq4XiPRLAEXhXxWnFiJ/lJLWL+yjR/MbeIZKSZhg
sETNWyzdppdHiUZzARrzs16O4pmRnO/DL0742LgAwJ8QvV9smJSDkbj1yzNqMGHm
L0aYbEQg26ZIus0Z1BjRlNUlzOOuZgjFv8sn8uoVKYRxQ6SeVH9h19JJWreCj5WL
+OgMb6CeVYXlaudRVU/oHdBkfWargsscRrnlHb6T2raMWBJbdTc9WyYJo7wx6H/K
WJDpvbHAERjF1fhbiT3nqfcXceDnI70XJdVyy20bwoo9Glrl11i4qwkW+2zZYS6W
9ZSj/6dUfhzove6W+N8k9fWDfmpLCGAv5Ze1bUo0vFkvKZgKwmA0lDJ49xqOkoiy
aTBs+EtfOS1LXF/Bjg+bbCx1OP6XxZxirpg0FJ1YcZ/ZqYDG2E8kU2wGs4bzVUYV
NM2YU8wXfWl3hzbs1hiH3tY+kAkl2CA+JwBJzPE8iC2bbYQltma4izk5LP0OCr+X
OLS//Iej3URu66To5eEXYPM4UC1uUy6AhQ69lv7QxVbfnzNqJ55pZAwW61VUFuMF
QLQ8+eYWsu0iJBFYvbViv+dTg/rWVbQqSOong9hT5vPyeMrM6NrUbvsfiyilQz/A
mAWKbo35QWTk/CQuJ2Cooup9BgLZTDFx7v5ADZ2LIJXpY8XgIbZcnGA2giUQ9/zL
hM2J1tQRaB5XQdU6A0kSEtLKZqDfSQJoG29o0AKr9zqjGwo9b3RpWLGDG68wsnLx
uyriDNdnkSu1qqCIsE9GMnRaf2OOtl8SEic+N+HexiDpuKAsNqKmBduPGtNh9VeO
IC8lK+6YGU9niEMTr5e5Tb2TlDLbPYk82/EIa27DkfBcxjZQRGepbSXDvgBvtYdq
qVfoTmPr6X6CcC/k4LIQyy/WbDVZpOWRmK1CO9UKXuODrVkkEmufy0mIF8wtzRiz
NrybnEEmDGFnT8yANgwFU3IGLGWnlqNutV5Jbeuk6lkdBmXeKwb8q6FV6rnqFfai
DSob9JwbzmrmoVPZ8PhZkbkuuZSSlcTok2/l6cHul+ZwUEstI/NgTFQJ0XowEuQd
T6hDuaDNg88Kj627pbGvhGwteQWv/ujQfWNtoZbZWEO1HxJ90RH57IRraK6pfitD
cZd5NBwZeYQKjfwO2kc2stUvKRG76abL0rVvZZ7oyj9Zci4toXBNOi2tB3B2ldhB
0QEJulzMxwIaCQsu+AvqvUO7GRG42thZ+PpUOLiMrWqCrt0j9T/w4JW0lG/S1n1Q
ZEr4DZeY0gGQarp0cvnikDSDVnHlA/pbPG77dLPtKhczzXJ4uFHgJJFQlfsSQpQu
8+FJUzDSwsBC9ABIzLy7pPvnnYqtdGAnhk2F1NGIqqw+jB1Hb3Fm4BCgMpcHSJbN
ChnNNjs39JPjjXmlIJW3Yd05AuSR4yK16+2gub/MJ4Dfk7s6My3V6t/wJjvPSrQk
R9BtCHeg3N76LAhNfrKaNRYHiRMJALJ+RWui6Mx/7qUe92MO1ni6ZfVfsWKpERK7
2LHcaq95RJgbgN1cFxuy5+fLt6pKK1hxG/CY0zcdF5daIA15sRA92LZCnRAVNdml
gk/A4ocmbYJmSudL199sU0MtScT2j3OsDYUEXZG9ld+UPbEoBbj5Fff5L3uHFPSM
nI7+X8607bGOdYRIkVJhZmYGWvCMLC2T7y40pha9m1ufLkp9uno7z82v2dTsYJ00
GS4rjS7MCQlUld7R6UoVtSLLuktp8jW4/APuhKn/bmwifM3JqqJbUBXjDXMzGVbv
gQPktE65SQckx24I4eHQb87gP+P7VHein5VOSUNzncV/nbSAJsYDD2F87u8POoRU
7+3ckjGYV7oU48Ujhpr8U/6PXlzkNuV8o8a+hCEAVSDyfXOQZ5D0kuZmtcUyySRK
GjD7HKomBU53a7F/GET60KU21zDsDJQk9VlThWU/3YV2jz4gI+oXQbAq6gJ2YJfm
A3G6Psds8KNTEBJbIhNpf4PMfMy0WkRlucg7gXL6vUNyjldfD23P/DvgbHoyBvsz
kJwvwlixq0miK+leBS2ETnic3xeFFulItuZjExeeKUuvNLgiWbwCnF+/3hvf+J/W
OeVII8/NRB74kez9HoEE5s4N/dqxZpx7qtXTjV1lOc7P7Z3WwDW3bEwaYZ2bo3Zv
ZTj0U07MiDXRxnsfw56jivd7m6L1zdgzhufLGREvE/hy2N4LLgA6rb76C9XuZnTv
yCDl3vOJa8YX++gjbashWOCbCnQN/FxTsGxYMesSTle9CG/NGG4ohpY2UvO2/5v5
SNtlGERpEQARy2k+dXopxgpP6XEdv+sesWzGVDWkvbTsFz5lnXMl6bjWG4to81Vo
JXzzISEKZwEwBct70L/0h6XO4Ig2YdwupIRwU8b4wOTlAR+h+vxKbEoeEjwVbzeF
Y2JGfaZuflBlRBC2w6Yfki2AFjoQw39/qo9mb+nDheB3i0tHTAYy3vH1iXFSPSpW
OrsCE7oUu/MRL7MHAejY/cdjSxuGYL1pkABMRgCnDs/lb7P0ljjGJhlsKg/kkQhu
gEQYIIqfPuWMeH/42X+FoWiqD4+zVKUexOnB94Nj6YwEKUHJ+dtxExRHl5F1YF5l
EBjaS0DwR9ry9H6/FnplCSD1loP7uWGPCTeo3C9x1E/1cYPYCasWu21exVbqVgbT
ASB+MharkOdOVo76Jp++z7med9yNrGu20Gi0zdwuTndNS8Fv7AdfaV1w0UXZt+Qs
bSPwT2RctQ72HiWBDStM+3H0oRtN2m6Qkr9WSq8umINWgfO6qV5yRCTiA0RjpRIF
67MWAcSWQPNdiDMsYX/3PUYcsda7ZgxAqW2dtXINpMn1ja9R8oGBaH1W1JEO/HP/
W9e/uBN9CyNycrHW9nbdU+7gZf5i2OeSloB+Tm1TN8+G/Y5J0HyO1/AcI1ZjsE/1
+Q4Oxc+sS5rboG0A1xVQ3wr+hakrjauwYu5xbRPC4Fks24aTQ9gYAW6iCsflR+pX
OHGYqGus5zGRHdvaLciz5ICLWQKdZn8HIBkPAXfv6NxbvlnsYaZbwETi/ADaBgMV
RTag2BmOQ5xm4rNBs9Y0pwz1ZiMxH8s/429b0YfL1kXhqqxCaso4hvXbojd5vdms
YnFX0Dj6C/Iejd3bboMed6z+/nBwV5oDUnl0PyZCaQyBHmlqtim1LQqGRvUjYvYB
kRTNB2Rct5+s/L6gPZETnLBuRO9apFHZbQHzrfla7F3h9PDmpt6rjR1oJA2Ibo1X
LMR8WIoHJCyhMPP2x1tN1ycGEgT9DZO08qik9sBnWXnfDLuyCXPJwYrfvsBpfhfh
4om0EyvrB2Jfk4X84Zjxg1mJdNhHYflzBPcbC0VNITEP5aSFgiTY75DHb4LfoF01
8kaQw4eAzU3wn3oLnVlMCmtUUFMugF/53BwozpQYnXdyXyIRxnUMmAOjcbKCh5Uj
SBm/Feli2fBaj7kSX/IwGEriGT9o6HOA3FoALyCpHE4RaAX7KAVj7xRc1EAp7yhu
W3aHZAJI5QuB0spYLyW0O4a7PnNv933Gfsu6FjdgJ9umki0iUj+ZuRefI1pwJqgH
GVrKqpILSikMqrIM4/z/0oozT2ZasECXxoZ72ljpLvwuShFk8diVMurudKnXMKFd
3mS9nKM2B4Ul78Q4+QBBGxc1m684bM8Q4XapS/BVGf5MR7P7FIG8ihWTqg5f1vml
KnGkMDEyjc04V8ZhoW96Bg76TJuvUjC8dU51jx3OJ++PNgZI84M8yNmJrCS+246w
Vr0VCbqMwmhoX7jj5uMDB1sgKFij11aqihzzKZjaTn6osa1329+e+bYDcx9WHNAo
RB4HQWBUsG9aAj1bTWiZs+IYcsNt4hQdmUcuJBEF9jEMeR/BbrGr+u8WWQ4I04/e
8WZ4iNOiHF6d3xVHcIiIOVP11HxU0R4TtWwR7w28XG6AnlRXiWhzscdyE6h3e/M8
u9h+zHF+wILTOMkW6Jx1sF4sEFctUw0ldIN2EXFRIGThVtnHcvOjhQSrEMEyEfhi
StDg2GB850dsoUfUA/9PG01clLRMuX03NLaD3d0EPYq+1qVbD5exWQF1ntU1XGin
7Pb1HIhZVQmbmubxNdmn4o0ttHtGTI3Cj86g6Zf8ox0BxOkFFjMFMExZXfeSaqEV
lhBEMXlOXafVCLkaF4OxbjBz2lNxBAJetxVD2nbJw4pyTQ+HcWUjJGPY1ENTU9FI
ZYZkpkpGJyhWnYP4WZdRjnYrG4NJ4Qz3SjNnYeBYxD7IOW4vxJrKNcSD9l6gih6f
1k7f2fIX2JXdnFi5po3v2DTDfUAAZuP+Ro6SA0UX7lJt0dW7XvBlCJOLsaeUcFVr
o0wuTmqUjY/3dsZrMxhMEA3E/Qd+ZI+K+DIZsjDHIN+prDgLIxStqz1un/NGICRQ
lB+Tnm9XZV83KEGTARuFN/zVEsQ0rbmrhCBB04GwCtp1xn7n/q1CF3LZzWDR1/uh
/avEn8p4PTTB+WUfOfC+cmXCGEKcv63cf0gBPqOc1qJT3J1Ofnajh6jvFSvQk85d
PrHdygWethiCmZ7J74gP86U9WKptqGH5ZIU3+Jy9g/7zBpJzoYgG9zslQkPgeOsO
0mS6JQMk2fBTn6cH3mwKzgqWbW4Oqwmz4YUyMyYjTeyQo4y5EGRqD8/yMXfEJ/Bf
ZQg4TwAnoIyAe6+Osc741HOOr4XMO9I1oyErVWqhU0z02Zxg6Y6bUxjiQ91GL1sd
f11V2JLcp//Dss9xHVVOy4sae71brJM0rx6KBuH/LnY1g9rlWmv1A0t0tJmsVvLC
vjU4LYyM3AMBU3zTjK2GnmA7nYQ3+LYMGL+A/fE7ylE9j/wQlZs+FMTfX9eBEET1
bfuwxQeVmZYlgrs9wBctsJ2jVHQI4CAR66TInCVpDBDABl5v0f6CX/oWD4GylCpB
ouPYy9pbG56+o7S1wXOS3eBmlaXCZCLHseuQcvGxVf5t4Jnmk29Ni6RkvjaOL8AT
Gw6mXUxUIWhcvaljODOmioawSVJJMZdO4BDz5CTgMTBvPph9AU0gzQuvqsPY0g/u
K83AB5waE9bj3m587ZI+NlW0cAc+ABvMn46hLjwwpBZ7TmDj8hDbKGNWDfZ9F75O
U0yVsH10cRvNAOzVWQQK5CQBLxs9+OeVHALRLN6WAspVeOgq7KOJmXXrNq2n3bt+
uO1FQtkwReyvXimDQlrZQE4iINPonS1nORa5XnkI7JV5vPs5Zgsv68Qj2HDWu3IA
YAiIsyIoKWo24IM8eLfnN4nFLPWHbWyL6zVcpaloDgpD66LBSP8bTivLRw1T5BfS
+yGCebujfJTZ1qMmd8H9Pt7yZ1Ytt8gNqXojZDWwpoaz/OWv+YHGNUVWnNm1WH4Z
ew4QE1sYY1qLVRymEAI8+bTBX4pPHV7EpG/8hj+KXYcJmpaJchV8OJ3y/HfoCGdg
kT/tvi1myIaoDcCkWARgBp0qvuGM5lN5NG4EoZf+qGN6yScVq09OKYIhOoiEwF3C
IZ1k7ZOL9zWZywt+1fb0lSy1x/78YyStlrVrHW1P/gnSYV8iTWjw61HZzmHkKRh/
TmDEm5kRprt2U+08XZKXqo1Qf2xCJCfK1UHWTcTvFdDmU9Oxr7Imv7dl/hbgz70n
nCYNSniJ2xDSIKfEyQV5+cn8oB0/WQBa8KykW98r6dbq6lYLVEu1AlSiapkWLCQm
DLCDrOO7+G0MvtJPZJ2oOj6Kg3L9WLBCthgJiWhrnD+EXkC7fCLTW20rzxHx2jc5
/6ubn4PtjtMKVynnBm+hpMjk3eiHpbTbmEJaNE4kTIu96Ar4DW0srJK3t4/gGSzC
kDgiBF6gYaIa8LkXUZ0r3/rV1tamVyG1F7pZKIDh1H8avCW1wIRnnXIaVZiYMfUQ
Vi27CWrb1QuCY0awAnM/dHOcFMJ/8bWHzGUxOUktfNhcrcRzUa42o6kz+kdpU+KE
iUKJkJAKaJUM5C+iN0y0IZynJ+n5rsAbqM2r5TaVMjJSU2kvBgAjM2rWtsgvD2Dw
0xLYJOMa5i4dlRkKKC/QZthWuh/zFs20khVWzJOq6qnZV4WcBSXDt82UrLWIdA0k
/TmqOWy/rhg1AlF3DTtCM7PGtKmO30MiWHZNvcFD+pZfwPbCkm7LjKvJDtyh9GL7
XBySUusuboIYkPQzu/3tbAJp9PcAY44KgdTkb1P92FDsYzeCBiVmQNMZKLV5zXsR
M2Z0XMfkCjdjTw8ByciNmIwIEJpkXYYAiaYsyI9xBmPRYbp+K8/LBCoV0sAVCPAd
EQKFbiv3s3kRgHQTM16eAtnE/YpFTj+Kh5vXBVG8iZ8Vg7jJ40kQwF/hqt/T0i+m
M4gFyyOgohW65Bitud5Vv4bBKA0OknGMCFmucGJsCAfucfo3tq9ppOv+rdKLZ37s
Tny9KxDQEHnV7NG/cuAn5Ik9OQVaRGt0WIP+sWe0NeJOxWfm7udFdowTTIhlGSTl
dT0FO49OuqjSw2aGF/CuWtlqlTURkKd4yniofDaFP6p030i8zigtvH2cY6mwKmKr
D9PM9foihyYk/qI53okx5mKxinEUeh0tIwSoTbvCYCyvJojFelqf0IaSTy7k3R2q
FQe2p5oWwsxLalPr2pW7m+4q+Pr2D8Cs7kQziZFJQhTPrAsC0LBEBWb5G0CXzn0R
OUKLRr4jn3G8Ao2mEtgsKR2HchRnQmQFfCNv48zZ4JJeRKL7deizuqPgaPuf8gIR
k/wxsUrFmHygSaKnxSIol0hQYcJWniUmfnVlnmxhbyNbREV+1WFzHMmWQ50MgALv
uc7DAfBXJwaeG+6z8VRr9oldgM6KKkOfpkCeKVEkfRlOqAIeN2CwtoYTXCPNPrAH
NQK/y1S0l2vs8GFgYiXBaedArTbMjN/yM7oiL3OzSfFBjmAatDBwWSXQLBy0QJqi
fud4HWcgkA4s+CheK32Z5fD7jY3MACh4A/md4zL30WnLC7hYiE3jQ+9VsIZGRcPY
YpXiXTNxwk01K1Efrzi2lSID7WRZ6EjJFVupE9Pzw52h3NkzkgIDi18iDGze0SbK
i76dqBlTBXaSgKutlCAl8buJBAwpTFOLEJaZc2iDIN4i20KVgicgxryF3rgTIyRq
aDN/1ItwhbUvydzNjbOrfB0n6T9sMFiMGOUo3WeTNgMYjhZ4fXk8AfrswHxWX8tT
o22f+A5P+laZwBGBw6C1OzMl9T6R4EStSgmlgubEn9kXlucLpX2RN6DjJf3Z7PYH
88rXXyOTf+nHQP7S86JYHesbU4DdNfu5IGcrA7GpMkKitQjphYcYYUUa8kTsoz+G
zW5XGkCh33t2tS9z5MgGNVkoAssBmvMUBI36rXkkhFHrpbrNR5opvZv3rbN8ChEL
YaY1eDUPZ2u5fevTxIkHvMNlqTte1hYOvEqdgblbji2LziG96bf7gWmAfgA9C5Q8
W38CZg5SJAXFr+6Ip8vA/+bU2zmGdrRjayZBtfVMeO7dRSMDq8eRcLRiwLDocXoF
wqlOTh3kMI1AxDfvN2gLPzfmtkzEE99cpkrHddf8wMZibKRTQ9rdAwCujVjBErEN
O+/oBd+kM8AfOAtoRjMXTb7vuSLZfLicrGsZB+jKR+gPHEdpkLxybkk58BrPT3Da
8ye9xwCpMF1Lam1MrmScX+KFFwCsifPqfSFMCo2xtSEwUFCzbkF/n7I3cPT0Hn3a
LPU8abUWSoY70aDnERDjuOWBIhKWK3rQWoAS42LdCtRz5KC5ak6Ysu/YUpbLdnUo
pKI53iyJqsMa1fmMGlQyR37CNqWevO54P+L9LhJ6UHHsUwe07luMqXZREryvQKEz
cPxZ/n3VlZrweRnnl22Utp+q6Ozten9H1SGFRrwy7/DtHTuS9bzvZ9T5QpGekR4/
IuI3AH73MrJ2jHWLVsJMVUb9gMc1BE39YYvWgmL4uBWL2pz5041mhp55N34OFkRj
+WmRxKljye7mDd121y2gQzuFbOxY6CHQISk7zjO8UhAXyu5ZPM39sFa7gOKq7N1B
adsbM3BTwyOq/rdfyBtfTS4pQmP0ueh7wrnpM7Mbo3bh0ChoPtJpOoYKME6aMaxe
2iPSVKPvF7dr8dwU8jEewdR5pOPDIu6WzntQRq5Gt6N46r4biRRwef1CQM0ankS5
p0e3uaH8VkkIJbB6buerzJeyfhgber75yo3OXIOputzPgQPY512dHnv0zBWUNwJr
spOpoGj4Yf2SZ9fHp/VkAg63WkXT7VjmIgFClPKGtUHlRrH5vPtJTF6QKVC4kdSM
WNGZ1aF1NcFbSxPSttgVIvZdBumb4IsNxAJjcBrXzJb+gOPn2dzDyn4J5nWZjSRq
7xAfqtLblDVzHaIVg/0DRZf7JRox0Cx9gNAbaD6H/4QJ6hgA6cXY10XjV9ZFwQGa
+eTs6wMimFIZoIs6WsFUAOh78/o0/bmZjP7Bx68sYXnctxCFhefU6UU4eHkHKw5d
Y6qeezthVWhRZN0Mw6euHAiIk9oSLnH8Z+GF61OmqH3wN/yiardIx1hTJ0SmWRjf
0wtXX/n5nL5siPDUe+Lu2qIHqDP0R/C3V1KaeaFIzFl1fMQj8hGBIArkwWraCYou
qncn70YsGZM/8IPRwL9lGE3lJCBcgCcUB2ZYafo/MIccxMJpB4a7v1JhKAvejSWc
2niM1jZxPQwwq8VtgfJDnPhJqUtjIoajST/sfFP/zXZvMK1PUqdB/jNEM9Axl+7f
2LC7Mcl5MDyzyCkP8IUOn0bbKdM1PKJTw/mkY5McuB6VVdLzHXiCAK7gW8OlifyI
sG0ywJDUY3F5urAsGSNiwjD6GZ1LPBw7tByrinPXVEd7YG7cAeXDUqOpvURWCZ5M
fsSQBRsEPBYusecdFExaE4ZGsTdf9BY9NhmHWHZCEt/4phJaOe+DiU49OYHwR6Ta
0/kD+3Os6VAiT5Rk97TmtzeyZdlLBrBu6lGM9xbhu8l29IgT4ufGr/IJRxfkHO3a
Uv0y4mHycOtkC5a1ZasVsnz7U9I1IS9HpiivycJl01hSnBVBBcZbPA0xiuRlGiQA
/WzIH9nYi5SsdKW+lTJO+gEwxNfSIbkJV0DW24fr755vRw4nZqIxS8gKJg0kJVl3
jVg0cL4f+qyA+g3qjS+vdcn/Npmu1LVi0ViUsbDzFhucqLofVbDyt9QIqKXy46no
QUne1WQoz92/LsUXAlJzaGWqlg+6byE6MjVXLRaXTbVgLD/JXFtIlAclmTTQC5NM
pPPO1I8FgqWlmSdNGEIe+L1qAf9+og3yBsmyKShY3xUbnlReUtgJIeXmlr/gF0Zi
Ap9q8ljWWCR8ENSXRqcsbfNkum75olCVlQs6M0MF/W5SuvbuhNp7dYgsq/xH0PzB
ZqVBd4IHCfVreMZ5bRk+nhdiLPRnJl1LVxDBgonzAb3Yy+bI5lW03BS+54OBdgyN
JrdkLAn1oUP6/AXOIa7Ui0kCzvuVw0KMLvdP8KrtXgnfPA7UFRInWmpQcGYz5BBy
BQrUwS7aNdRw+x/olnpsFORSm2O+97bwSAReA2jI90HYpWVJaz038pgeeHBvPkT/
W9DfxofkrPFV4HM5LRi2x1g69to5SVWVJY8D+KId384EoiTLgntBjAVXeVJ4rIoC
q0Lk6KzHiULrB6voQFEb2ahRP8VHKgqJwUCJVYnkv53YKMYUR8H0sNt9uLDsgbvJ
2uOITxHJDjwJVhPQQI9PO7qlhI/ZOiXZQn/kapPcLJWU6toJ+Qlh13MKuaRhVk/0
vBAqsYWISfV/o6gXLj7R4A+eGXhQ4TKi2P3inHuGrQSzhXOdc95qOBFlDwcoSURi
kGrCNcm+0bTv+70Sw8vnSgnmducR2X/KCLJX1DR950IdDOfiZBW01r9HJDAYr7Cj
SiUKS0caqUoj+S07QXqaaxx0uJ1x49hJvX0scVmTZm+21gNq3xiQowEz59xzysyF
KucRX61X9UvwK10I11kFKKQLmgQqzd7K2eWuIWgtgDAGxmRvzQenpf47gNn5OA35
c6awNdtG3DhQvKMtXTLPp/Xxy3slxXhEMiPog8vpt5Vlrqrfn2j5454WBY5NsXbm
W0vjIq675uTLlzUz0YR1xxdklNGV7XG8niyJETJt/prStj9E2YnJI4lut71N66V1
sWusJpT3CdVO7XaRwMw7BrPzG2i0QKtYiX4n7Sww0aTn8LiShvod2otlj22y8ddM
Lah2S+pWwMXqJiD+WJnO0tUurSWQUc8+rxiLJDnXCDyfz0yduqVM7emSahMI9KAd
zfwkxFoFtn16FSlBYDe6HtkEWTuJ51sIrCt6vkc3RIgh2tcHbHQEZMskzeECIVCY
rs88IOi+mn76T2ylRA+k+TnybEVbJG5QoOPDcMimWF5RAJp49XlTg2b6J+lFReUa
MTAdMzSxTzpw7lcV6nozybn8FMIloIgfhrTjshaJclwTts+jFyYGyzYQTXAPlCde
z2Hgl5vokIkBHjpnd1bOgFKP/33B5D3wFJrZuoslb6jWxux4+hfhrNjS+jsYiJQ9
+ssyb9L6Rvvbk/cRWG4h0d+KWOPAwj9WcuHV8R1Oomj6zfzOIBMf/kyPvGTGeRLX
Bd1ZbJi0WdShXzwg5CDjB/dDC7CRvn5Fh9uZGa8Yr4U150Y8zMfQWDwuFxTjacmn
kT7h/fvvA0gYkRxERtcnw0G/GRanqRlmQ9ZWwuTgz7dpavFSw1ouXvwBY/ltNlaP
MfjrFz15AxYhjgkBi7wP2bqcMZQm0sYbUeA9TQpaHZ43Lxm3thPH8jx6AOjj0P/T
h1c2NsOsX0pBR/3zd/OLw5jxkqIER7EewR7vwSRvuFbAef56S/qbMTpTB46rJ+I+
5OeUzrklmqxofLrOaXdCwlqyLwukuKR+tAZE53TF/RhUIql5L/ZQLlc4FqUWlIAu
difC5KkkoL0m8Soy33xi28tS7Z2ZAvMQLy2dGXYgn+SGvPw73EV2aKwF1rQ/zOh8
xtbOBFoDiAk3Cymrg1ki/NHrTliztzyabjWQ654o45UgkbLGEx6lAxREcQ7DSgMF
xLhYUsyb63f6YVa93HE3lgOPQLdE7RY9igrxXaJOlQ9A2t1e2D/r3t4oWbj0f4/p
2m66lUsmKQ8Y3m+2wfDuL65GElCtR01X7w3PPSqaansn+H1CW2IO5v+j8SMWAtpP
bsyv8frf1iaDCIf7YZ23U5gAvTn0LSMTAWnUqR/n0SGHf6WerKaJhtdEMyZCpZRZ
vm0+AEjPF0hEoiIfizT6/Rnylm3kv9YhdW7JDwmrh9NHMgzI7giOjGIj/xYK0glB
qOlpf2JwGUYQI+fWZ6p3Aq+jZJXb+O+oXSMMZgV3aO+xjYlhXQi3+cmIczDr6Qw7
BJqBjyEO+l3nTFGzHv2H48ZIS628YmA3mD7Yr5JZZvGw9oElTc9vwNPnt7lMLw+N
TPW471Xh9dFs4y3IkLePo50ufpxuNA4m/qoe6kuZETVz2CVcrG6XwSXVVSvoZPX8
Q+/glI9gOa6q7zG0kvLR+3sNgcePN6XS6ml3ZaiiBWgK2s4hGkNv4RZUqVhIQflU
CN9oe7PJiq002SaLc5tHRQYYt273+Jcz8WpnjGvA1tljR5Pu3OjDPhONvFE0GVwW
DqzJEcp0OV56EhMOu9+DLkADJMxZlheBWJMesRMpDsE7Qe4wUp9gYZpGbjm9lrRR
gTyk0LLeRPjGfjqXky1Jixkpj9VvAdoykNfaQIpeqYFJEhxMpuTG/Xo1QMJpoqbT
K/f/YmNK5+yM0gc0i0iQIkEmOBUxMy52NYHqY9uN1X27tQJhB9GwVLKoOI8wiQjq
9oaeHUzejWoUepYbep5zLwQZk6nTzcXlLR22k85Bo1vviCEWl962w+VFCwxczHnI
nV9uAj9tXbRiH/9fSpQkEkh1/w6LjC/FEa1sI70u9i7kZNeJAbHlJML86rjoFZ5/
JYt8oyzF1TK4ibPMuMSkXwg7o+dJsswD/ZN1GV7nvho/dg0QzjYa6fJLK7970HJ4
RJf2uetlVB9ElP/IKpQTvO600+1vytKegdGswd7OCPyIxy/0nxLp3ZEc2/3mlQMM
4ImQsjYe9srZLYMzOAzGG1fp9IE7IUpsC7JbBsTImJP31ogdZs40A7LHgHrb9zwj
dvmcswBt6YyJRk5pQC5944K2EDeFSMrsOhNlkDPtYJr9OHYf9VI9QWoX4kyrlcO7
HOuHWjJaHn9piV7UW+JA/xGBHUw1YaPFnC46zNezR+98Q6vfifalNY+DnJgP/h3C
8zXXjCqci2/64arLZ26y3k5C6pLRoD6uotg9+i8APpGGLnWq/uEH1xLZpsMLbAKs
7RmoORcaykydEmHuHZO1+KD3CCOzacjnnHkPFxB+mxLEfMyEDjiZ2P+f3SWqZdTU
6c6QOtW/EgjYLOKvhivqdhWrHEd/o7t4Xyl7p+3lnL40Goaj8fXr5VHuGMhZpgrp
J0hNjtEAbUYNN7nembNLaKBCdEXhEjAzTv6Y7la5PWlWXMq4Em2viDlvcH6AP/rL
ffD3TS98xf6g+qKFYos7SwnkB014Tlu5eOZD913z3JiDNz4meczeh973twoUm0xl
9XAYkWUhhUNbkZuxQe9d1RM2Z/27GpwF7UG4SJFRTtB+KT7uiWC8HnPDGwL3jwhR
myJufRKqywwL0bOqKOE3f+NUxhk/+vUkUClaZWSI9HKn8npRQGc3LxaIg0JubPIK
8nLog3kc3jXtB7/DrKRUBbZshU76Ux5XyRZt20RTb2cSfxTFVPp9AJn7DsYILP0P
Iy/RdYsaJnK6Q6Ru7WFvwzBPgyK+XU6WmHN7dl+GrUm2o/VPFOHhVk4gkYgmoOqB
a3Sy5OGZumppELN6Jk6JtQQ1RcqJ7vLObBiH5b6NHqxp180EhUbDAUFHc1GLRBM+
uWJgt9DRfSW2DLWbFoHghGxaslHPV9cH+H1xxWMq/gYb7JfpKiPQU07WAPE3fEUK
v9t4FYdiAwiYMoeTB28vNqD569wo46igGKyVmgde1inp06sTDPcmM84VSkTVzNw8
SoXCkmzoWaal7ndDlmLw3OuRf7lLnUiAm5nLlTGq392PNXCP7XsChWRUsXmQrF8t
CVfoe+YAi8LrhfRxp87rWcyGYR+q8hU4me1Cqj6Of239wPhufCk8b47BKCJE/DK+
7bvoFFQt/kM1hp4IFquB9I7HQvUjI+JhxgO5paK5f/t5AeLsztiiU2LzhiQ8n5B9
nqOYWkOH4qvibZ9dWVLGDhQEPSIGkCGrr8my8JYGZVWKTRMOy3Kkwg55hNEWvRIL
rXZtR2ot5QSgJKmEPyBGXf/4WAJ9sqeVit0xW0qgX38WplGrYUD0V+PgLjs8QKNn
Bypu/LlI9t6lgG7krNVMx2TGlcGrrGCX7yOR8oypkdWpIuLD3Ss6C6zCkX9Yw0Xg
TxZh3sTMtYZ5G2o3RWrSkQvCYj117LKdOz8XU0NxNfCTkBRweswq3QHWyS9N+LbN
mB6qeCxnZ2BW54wyPU1CZqmjK7xUHpuBezPdWO0ZZLrd2IaS5Ypuw7FxsA9dnTCv
dTubJIXRguowWFihYHnKxK2fbEoCEUruFRVnrRTn3iWRMditgI+6krRJkQpTwWpj
bxOddtXUKiNPFEMGXPFziHROOw+wQxIAh8pL1vHInGw46yGe5wtSThrZXSDUtzah
coLZswP94arbeCELZYz+ys6FHwRXp9VGd+vlfSQUi2stjLBHo8+AhHyNZbafepwP
t7OoB7KLEeJbUx1hlY/AhbIWOH/jX2cpJUH1AJREjQIWK8tsWQKdtxysNmR+bnah
MyhGUiebsCgYZHZYF5/7O546nWWJdViLKUHBC0Qv64tP0ShCwJvdV8x2ODCPMh3h
Hz68B7PZLK0xSgG05OGyg1xCnIqz1mrouzrsppKnUKbCNuc9iokii7RxZ5U5LSk7
vnzxhsuSNtiVU6n8bWJNsfHei9dyzEvfM/5Qyw9IwF7uiUbnTwEf2VJJMsmFTCAu
8Qp4hsS8T4GILcDX07Pcw6iTFxC5nbzXBE4hwl7aQs2mj2RxAvxijjmzHGnoksxO
msFSctPxFuNEyedDJdn4R17VxDz4nOOWXwkLIiyuB5DD/TMW4M3gr5+LPw+PDFKh
V6SguaEz4tkg36QOZvdisRkEvbAC9glMPd2kzqax8nsZBtjiSaA3GOyk+xVWVG6p
WlSRywWNB1RB6kcjJ4VmCglvHemRpm+/iYzx05D+J4web4jf+/NNdMBq93UmjM12
ynch2jadvpCIxb+z7ShNpPfyMs7VRJAjvpDygBDggZNzNnuylNcCWvVYM6d4Ho3/
k2XXYUDxyADAaKB3G3zmny8vXRz0zBNnkgMj3bG4Tx7sw4LIePa06CMoPQwkpbIX
Xn6SjYbZ9ZL1tBBXk2d17oLoVzDVkIn++9XMXMT7bdWv4BG4Kc3mqBi47jnHx2x8
jO4LLC+29b6cNWB6/QlHLZmZb27npOBuPfeSKvYPBw19HKgQ3vkaf76K0FoaylOa
k5RC54RbvZ8UWwwHOlaKQXTO1NCiWmIEjapI79x6ZusApnrTbB/YgKtj712LNpxb
DCy7Dux2sgVE2WXWWbwuPq2oXsWxnzK56bngd7Klso84ru5H4Lx9b08HnnO6CDPT
Kpfpn4a1Oeo6qnhnP4WQc9jLviA9xSoe50gyqoHId8Ep1cQJdX3AYh/yjO0WoJnz
XbhMZ1ndHLHky/nEsN4+tpCi4Z52gCF4BAVYPQBNAwf73BDeAf6i0InznNcuKbck
TnwsvVR91Nf9iTE/PHQDkiPa0fBCibFsKAFZrCg1sj99um8FvKl50IXsokSHIgNj
ZcIerTmAd7wx76maiGvq+pKQANdLIVDn95ezkjO9zQolW/ptuTjxv3uBEkydb79t
0c9sihByur3RMyDzh0eFb5j+7KW8aBLH2gwJ1MtwKorAHUndm5n82VKMdFRvTqkB
ZVsMjLvnrLhCFjbM9XKTdWcN2QbcFUib7eDY5lG2EUiUAFEig1zU+bbeHP4fERru
HvIbFBUCzb3Fbdh5qkXxSAhnUULPXGJx9HQU9LGOkrSTcPnr6aVsSwGqYCiG3aQK
jECWe0HeotQltKVbHHPdOmUAdm9QysG2pYvQ7md49ElIQf5CbrCFlFNOZJBzBjFj
XCra2Wm3tepaqkkuT5uljB89A5Q/Q0oqu7lh43vqhSbQ+KDFWGIqw6mU8CoHOSQB
Org2nZb3+w1Qxm5Gk7DpIOnBA4sT7u4y4WZ843P73Ccy+t+gGPc7OlCL0Gmd5qnw
`pragma protect end_protected
