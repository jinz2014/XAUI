// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qnfi0RpSpMwdnyRAfRbv+4+mSMnJp6xFHYSTfBq8MINFi9KWgG1j5/AXY5eh+kI7
DgfaYjnSpqgUIMvQRbzSEH5eZdVW32zVA4PH53dDY1ApHpVfAp+eRoZsNOHYZPe1
+KxeQz03JVhmW+YqDHq75GOkxnICfqC9aCoRTOAZnYo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2885024)
awwZvfeIyTjREquPc+egDDZ6P7juftXozyov7dqYFkMfgSDDzM/qrtgubmJfv/Wc
GgzrNa/Ml2yrHD98XGpc8sjmH6bxvaPJbMA/Lgo1Lnc7c/9Ij4qdtNrDGLZyIF9f
naqI14xB5j4B2SUCMWiPxrAKFaNfMPOkrXmPzIgz5FxuJPFGe9Xo6GCuzMyLky+p
oNgsquvA7Tbt0cGD8lZGM09HUzXd5EzVXQ7F5fAS0e+TJVezDbYMhH05hpJbYkXs
drtNWCcnqOn8ah6qIA7e0g0MmJsXBpniYbYoq2+4pAPcTETsEbb5h/fTIu8hFVcW
Uo7ZqKIf1w6oO6VFcEC0issZJcdGjg2V/fj6khut/rrCBD8tRlppuL2/uEVtd6Tn
V2nEWjEYzsMblnq5IT/uaIYVFv6jwlTRmFW1V0qVHAU0yCnM+gvPFWCJN1OMzTQp
hxrp5SHulUWrvFI+cpz1jhE6YEcpgFjdhb34G9MK/Nco4nb7VVtoZRT3hYJavsMG
QDiwyiNM0ySVl9jHqR+4pgYepN5eSxuYPeWn847YkICKaQYrBRDozteucv89dKlQ
GWe/y61opapY2BYCMGwfhdPkDcPi2KSkXeNBEzRqcp1vRUEymtjf/yTxHnZLqrxk
VMQ55kUUb8s5kUK2BE26VXpX1S6K35L5fo+ASOjfI4/RBGSCYs1rklrJ2SaaAi7a
EEiCsKa7Zv2dajUTxXfvWo0cPnbWyPI+2MAI0kZ7MJpUJtEK3rhUzDRSggEAjP5q
9wNXUeJ8E97e/G7iZrImfu6sIoERgOr0mYq+ptf19vN/Xwicrs2vFejGeYOBVYoC
IYSWOjFvk/011yxQ4M+AsB0Zdm1cnazmS4/MxYn1oKuteq+I1r4iCV4TGoBERDtZ
GSEEGN1Bg++nF5zYa3WJVpTdmVnYzh6kZ8WXwvBwbyLZJ54wNYzW87UoQ4cUWlSA
mQT/gEhW4PrtuFqrxFwupvh9jCqb03FnHLMMUTPo6wEm5tvACUmBmIh5Hlen5C5A
aGmTIDeFs37ElTbDMDbvVP+hdhSfG1wDu0xe6AFOM4kNSJgoRR/Czb/zHilC6Qnq
//UbZCaYMoZTQ6Xjgoaacgyna/hfcaruic8Z7+KH5sYx2/7KWBNUx3E3dXAN9SZm
iYC5SubRiYiIsbJSAk+47Z/V7JGIO0S0NNFSEWAB1oRrDzGGFkQGGYMGvXWu8ewY
wBsXy353u8KLkI1ZeArhL5mJqPZLpCwSqz12GCiAqCe+Mj3nL0P3Jf6yaYT/sCR9
sI5eLlPvgw4HbqFiAKLe8i1QaN7SvSvC8ETQFshQ8/GxV2X9aAsOGyuAmpEE4PzX
vxJwRL/UO+rt+VrBCblTbjcbM9ZxEaJ4Aijl4Hgytrm5qBWBj3OYo+JCdfFxnvBV
jiPC22i62NG8rYbGJBMo8k3xqg0QQ9odvcqxT7zkHe+nE8rWhoAmN+efu74EuxPn
q/qQB+FtrmfkvvNVzZN0+vkOd9uo72KhaN5OE3TMCDrIXweseNGNYuxFrEW91Ys/
RYq+nJVY54OgckIQstr0AQKG+VqjhZWONf4mi40FtNBTenudf7Xqht49sRE7xdLE
41pTsHKnptHXP8qawgBYOz48ZG/X2RxbtFfvVSOjGtmthost4FGp/iYPVjKUOlPC
E9GgaJQWloizfmYc6+GxSkZ5VJtmLdL2hj/MEFqw/jNEpMJNdBvS0Jl2HYVLqasM
1Eia8E4Ex3c/OTQl8pD8QX6ifIcO9NpdT5dk29UYYO/79cqfqjitreSBfZDxFchk
O9p0ETG+K2baRB4u9NKuOlEWpTkl3hw65d+NNwn6xqjbSuJvR07knXlsqfXrI6M6
qx05AhLI5J/PsEyaGyHA7Q0X4gGEKiOb8ubK8eaQDhViAjoaTvwM/MqgTAx+EMKR
VeaO1bUcD7+yU8Y6M4gnSst/PrJuZaV4+BXTRsXGrQusZnOjX6+kIVycIDKrHDmM
iuor1Igas2SZ1Z//nXvsxsgxbWxzFQe8aKAPPlvvVwvYizDL0jyxFDd0ht6P3PuB
qRy9n95dwJzNmWPm/tmow8DtR5GOr/dYCI+tcGzV4+s0I5A6BqvicNvhnuFWc964
ZRFzTnzsnyXwNKkL7Svv1HC9358zOVNBJQNm23IQJj5mVaflknKj80L7aL1YKoi+
9A/XM3dK2JnJM+X4U8urv46hFk5weQiy1a274WFoYCwFfGJypi3RyAf2DT4tFEyt
Shhm7igtN0xwmhWsyha54npUZsEc60W1iQ+kd+ggWz6MRt2Bpr4ohPH9Qk+wRv2u
rv2HoZrPkIkBqya/rGwcI2OIGkbeACdJS/b1DFzFVejTb538r5XeuT20NHq7JNt7
02G5L6URgznuIqe3A6mKw/wdv2RBOHJSpfqSJ0DEEfm1G/dfkJog/wXMXQ9jCxPq
eNRiaXKZcsiAYYlrv2mOd3wog+HOpw7dHVJ3O7vwp2yPrC63zNJe+bJCg/og3nXq
bctxklEiZqfGzhvwpxLIJfEAjYIZDQAd5Pollebr0mTbXJ3zAD6zuUljDlsk07cd
xI32al+OsFm7kqdjNoWgtPOLF8a4aS5wcCyj4eCrDcE4tEZEzZZnlqlzURuzeHEM
hmiGSjuWxMiObnH52Bdl2BCUve0y9QHxCUkL7CeiJOYTVtiFgvYDQo+J75v5adti
6TG4G33JSoSngH8mNTy5M1LigwgRkUFk6tkehJDQT8ImN76K6q1mgcYPOq+LXmYg
I4+ZfNdiCyADD5aBa085WXIygHVKSlh8h8FfwIv9jz5Qp4dO/Ya/BEZzHXQVnqxh
KNZPzEqmKlFM1e2xt34IKMfyHnR/nY9pb+h5OiwNv/LNGq5NfF5rpIKJ9SgNOClS
CPsXsHxhaLvcdcz/h8XddSzpj7cA47Zt4ZomDng+3AyjEJ3XggNeHft0NOqpSGVN
Fweq2fuy1XNgIwWhCQiLIQZJ1wL3GvdXR7yDzc6rp/5uIQNEagb7+Xe+wtM+JU8j
vZUDHqDgDJBaEiFObMgtkwvOB6bTuhzR2KZGwzbkNEKvezP/jwI3Odi4GoliLjIW
hfNoEKn/tgMN02yLZS8N6qkncGwK/JhWme53Px6A3NZjibBE8g2WRA672IDabSEC
RI9egHZrVUMsY1V4gcdpe98tKEq/QCubqDhmGoOrL7APUb4Y/x+zlFgcz776eh+v
H4BCR9tP1HSRyjxVAqeqFx0VN1tBVDXGggUoe3eJVWgdLskhwZqMGfPsv5DVtH/f
h+uISGqRujyPiFCRAtnkeHFNHo+dDugE0jPjuOn3AQtk0cNVGtalzYFGtn9q15Kf
VmKcNvfkxRuFICwW+Wj5wBvA8P69G1srXc996SiAOVtIeHaONVaAOvqb8In1X79f
cw4pPjDVaHKkctCXJs7YYRhVzmOzYcZG0vxIu5uEqGkJPrVR1HeYyum2Ydnn7hDi
Gq63N3UIPmJbnP0KeafYpBBxODpxdGY1IWcbwoSPHYNOcrT0Tj4pr8bqOVXa8Wvp
lKpTSbQ5kQFyX3XbMW8gHLnMif7oXxlMLfFiZiM6ngiTzARVw45giDB+eWgIURjI
hsk7CuVSfZR6T5ouI3jhbyDXsGuywIhbUh3ek32Xedg9NahNIGqqQ0ZB+96BbxeZ
3V2aaXtaHmLMqE9Xqs3PhcNhUTxP1GFSh1GW3GigmCoNXGw9BpZLftAEQiW8C69a
k0xb3T+oBHcC9a8Rc0kVnEKjTZAMVHVIYXAwHYT90T/e+zq0qox/Eede0p8vz0cg
1i+rzP2UzqydhmY72tj28BWj2nI1Vxty2f9HwtoQxcp7Bp6qbGHju96LY6cDLCT9
2PXSwZIyvFpbK8NiOKk1cM0LlAPA8P9m0jf2nmaDT3iTbN/X/sRYfjdrNbPIPPYE
GCgjcfxAweHxUBmGmAwWARrpqrxXsm/oc5l7OGBYfGZY+0wka+MV35hgYtQsYep7
cX7FoHihNGRAbZlr8r3D7nw/fzz9Ho3jzuLsE/VqhMH5rEOCjHjCT79ccxVi7qkF
0aBVj4Ifim1A0n9bKsNa8MnDV/eouOpVGaWOx9p23s+KMqnNK+7SnP75YWVvlYi6
QT1xQpDAeMKFNBzhI8TZplRnqmloAVDsu13LFIYnAggAZY/7IouzPRlcjj+jYA1D
T/WcoAURFuWA6c3FSlvPd9l3VMJKgGIFEzd1AtrB1ZfQrGQu+eHWoE9j3qP80Vd3
0ckprowLRn9b4pjwlE1QOm1Tf0y0hvS9mbcTj5770iwBRP7wh9OMDjW+gy5CLiFE
To/HIRVC6rGJymaFKVBDbHTNqtAn9mmdP8M94dFHZiJ6uE05+AYPlu4dE8ipHOtr
R/fWBi3rxoofOyWnNbVSi2B9M1onXvhSaWFK1LAb6Tto0lgduQa16Sa3nR4I24HZ
a07YmsJxYnIMbv7Vq77TO6/agrMrXPgQgan1qGjExKVixqY379cYmstx61K3wPko
CTWB0rHM91S8N7UQofrpeYGdrrZIlCpqGo07pFNZVtkVYKfDqaSnc6vwwA7dY8KS
L6uJyXaZBJmHa/SNIq6TIt01rS1ctr5aydFUvrE5pVCXpbxWsQA/4d3s9OGOz/yt
LbsXz/Wz/K5ocYrZmh4tjhDWWjQcsHuli5EGrlxdC+tg1MNaYN/Mt6SIUyg+CTMB
DaqFNSxtznEkTbKLxLUYOdxXJEqqQyC+UWto+7hxRXBDYHkVqbLYZseJkSLMQkO/
EWCED5YbztDsnyvpdoja/zvmsRkkb9+u5kZjTF/jgqcmlaf+XuWpDaroJFniQI6Q
vRt1MR4UoBj4hVJkJ7xyVPkAr96cnsECZlRhWVT3uHfznKwE8Od0iVTNxY2UUQD1
cVUNcaK41n3ulxMNwcbKNnTPvjE6nWNe5eAy8PTYFljVVCZwPHX2jr/SWA74WYDW
kIl+CmuLq255g+TB2ypOs+digTATUuLSihbYaUohZEBG9KyjKcdxvFk5AuWRnDI7
p9pQoQCu+7FYvVRxn7roiL0xxo+sOfKQJfrs/gL2nz4doMgIxRILKKfzyO7jofUB
F96DojdALrJcO3IQiHwbbq+fZlALTsdog+wkdHSNF90JYpLj7FpJW38UYFC7pyTO
0oiujV0trHnza9+WlWvUWPGj0LzYiQH3rOZm6q0XeSutuG7IhHUFQ02s/+PJ9FOk
TwaLglBMuX94rUGnBpjo5YQP059SaYEliMifR9KM6KSl/I0Gege8OqDLFTgKIPgp
7XAinV1PaOMQiZC1zWzSmLEI7YsOGmUW0ZzfL3wkAVaUvadPmJuLnoqBc40lw3xs
mCueS+6MA22jwTT8HPfvkrdxrJNbAfogOlVDE37S0Bys4bxI5TSkobE8rNchOC1M
8oMRlqcHK+hgwGqX8uc7AYaSkGC8e36lqoeTbW4YeTYNy3ORgMdGwdH5lVvp0CUB
pRQlxBTSsOvi9ypglY5H4QIOoLxdBIbtsWsxgs5M3PGi97QRjeEjjbYeR31Eadfc
xc388XgWGnxaqc6DSz5C3zLzaLY0hsQWsNy0qacdy8FVwpudkuUcDPZcX20m182Y
+DKlgT/OyWwwJZI97KKkGD7ZrDjap683ACTEQDNhB9hzgeGWcJsy0altIhkq+L/r
ln/TpmIxIR+Dx8RwwCjEN1SQXJU30xU/a8Jn2zgVVzfiZXMRiIqX37yhrmkAEn86
ywQwFC4gQprVvnOgLt3hMiPOb8dU+42N27gpGZZXTaX8XehG9UNZyhOEm4A2+5I6
7tX8JXUGyYWGxK/EvFOXP4ngJPCs1hITe3juf+qm9fG1bTiyyOkP4ljqP4vyGlhB
rFqACRnmDU0dup5N43YHGozCr1RwY0yEr5tkhCjKOyRy1Se5IcQzTi2RdFW3zcLJ
jBaNEzWT7HWVoUNj+gojcwRcpxk31Yj/i6JBTmvDrkPIFGud9+2RZ2OSeGlp04Df
IwSgT4hWugFTGxL4QUvaX4btbj5hgWQLCNZFNTuYUNzrWPGKCxFjugSlq1CvpFqN
/jDyiitdAuLVFC5OrvPy+6hnXMV5JX6OLu0c8HbsK3KKt6lA0ida7h76connW2eg
BomEjRonZsL9PzeIX5Kggwnlzel6gFZIIfOiUJ5zNf74vbdDourDxeVcxuB2KuQj
fcAExPXxQO9aOfPXN4E7QZmjgbHYYSblaHmnuhVGI1opX8myWpKPvDuMX9Myy0SM
xaPo//JYCgsBnDTWvSPyTfMVWtoVUGzcYl61uZSaGvVOppUEK4eg+61ato+EAZrM
6ragQdXj5i/ziZ9a3QOUAScVVn/bJo7jQ652R/hjW0UG2e+esB13DMnUlu47VinO
se4LEyi6+vdhB+H0clpxeY8Kt3mhGiz9lQLldPFWRuYQoW0GIDk5zXbIykDObbkM
kC1IpH0HKfqcAzv36bBVRHywfU8ofa2YhQTRfzZZNUnoWiO402irc/TUqzN9n2pM
A/iO8CR7GH3PtXGTZboF7yH+wRFFG3GvYajxf4r9J/EfV9itPhCZFzkYVB06EzLH
ctYssp/iRKsnuYY3243+pxlB0PvGmBcXrdr9rCX/1f9tVl1MoxJ7HIyhoIwP5wjU
MBieaYgfuyHFDDHcxHXsCJtyzVcWTUN2PonngOaei19yKqtl5R8lSz4O6HTzagkd
Ku/BMgmDwTl01R28jo3dzWVUYRXVu5TjQIUFKDmIS3Okhhh4sugugFcFuwFtHyAf
4cu9Z3dfHdDGPsEMKHsTlmQ5jM3QqnCY+CboueEc6hbHkf+ducEqEkIF8PQ2SDhd
myWgDbOjNT6pL6T8SLCTCE533dLQpYNXm174CSoJgBsx4TCtp/msRIiyPWTKatx+
41pwe6T+uJj7W0zgd8HtkQeBlDO+wUTBjZbt4JDPlLhy9fN9bEAwI2kPdTQG+Zc5
nYIn0d293SLQn5/YaKwosvtC10+0vz1Ei8I+Sj6XOGbHee6lqZEzdhClINMWbZ+9
QY9zVKDmdhQs8b8MIY+87W8PBc6HJb3DO+9ZgfDuRrnomR1Vic9ahW1jld+K3joZ
GQUHigvzc7XGeul2lS1LBhTLMskBzph8b/YTCobmjYpkI02N+Egz6DcXcF3MkHtm
p2xiYHkMiJQBPHXvCt5VCinMf+fl0Mfwfaom6HAsgazgOHP5Z/zDnfa5u5ypFGIt
qlBbfoI4w7qmURYdEyQ6tufFd9O3e6bRFERSKNHxxhtETyT7gnyew1ZaC3eRAxze
u3qe0a6S+1IKRPpRq5DZx34pg4bdqyGcOC2XYbcruWCs7XK9yGOSeGRvfvJrCW6D
HfnCwkPNNwyxaTdzDZXTXwgz2CO4zB+xCW3NG+8V9FLLrGlZlBCm53cz1zfDYGgW
MvKcRcsOEp/iBDz8V3tKQo5fOoscX0xYwJSCOvqd/8HhfWvinZvojxxxdRHC8Fvz
De4m6ww0LSnT0UWjtWlCExr7ERA4T/LoSCafUwcNjBczy9jhe21pLjUcsxbIyutX
Ouuc0ldjh6so9c7eZsi2/oeD/rQOizfUnRw7UbKuxEw+NsLsTitsjnsXpomYcqbW
KWpylV4op9z4cJDbVoD8GKWY2wMOccgKxRvRXKuevrbuYAhmHd6aL6EGaL3ICbFl
ZV6eDbthze5ho0+S55GVVxT4ZlM5OrYHfsaeVG+THdGJn7aZiTqgserGIQhUKQ0d
tCNBvSXW/JvvMB+JgVYdXFGs/cpsDpIe10NLYXEpGJ52UUGhgjC1jY+EN34/T3RU
SPG7ZwMnXitx0jLPyWecx2qZiD73KP5JFCu+RGyH4IQ408BE8PPEYq3OqAgJGp4q
f+clvuxJ02WNIKtUIDy5tHBdGduoKtYx5DagkMnpwwIbIzEqxnhkc7vkOPVGxVru
pdmFbfkFEymoO9toHU8Chz90gD2A7/QoUmHZwc5xg2ldA5E51o7AjkNeabeE/8wE
25cckihhNJYm4415gJUAcfsbURwac8lUsyW4F4hBia0mH9gltQqgzWnin4Qbb4qp
/Ex2WUfZknwCOg4GAOM7zoJZiOXfjFyaO1LM9FxTXVt3rjLP2dLRczSddHOOsiQY
BqNA2are2PTjpJ65rOnz+hIn3DuqAbimHiohfmYCmjt3g27BqIqnv/UwPp9efsF8
xaA7WlUbSXuDJ9S6ARDPzY3Yb2u4mVKYqikf/hWhdswkSis6/dXpk9M4uL/mEIrz
1dzh5WhL85cCq3vRxKob7dXeL5TNl90NH0C8UBJAHbnUD8Sly9jQEzKdls9a61eo
X60mSVdGfvBy2OzyVSTxAGJafZB/HV2JiPzpwNZFdAA9DpFg+lqpwvayvXUF7oht
RD0mDblAhEFim17TDzTTjJott42XzCDOgofjnQu0COcMIXO4QbnnZQaYilkEMzYb
4eIEnfT9oCQW8rOZT57TDkB3VdHfHKH1ptt0j5rjmJ01/WLDC6ZHH4rcnrkNBco3
r3nV/BjFZNi18ltsKksAmZlVjj2EOSTg8wxC6noU/6+k5/cdDFOC52jp+/K1mNh7
IwJtxMRTsA09UKKD/0sRm72krDI4hIxET9rfhOLvICKv5Ql3HbvwGnWlyew+Nn9x
85tUkxeXJOyYYrPVZ0GYrkT7bK4isu4yAXDnO0KTvDfy1T8liPI55GKeBYkGDwUA
S1nE/ybN9ZnbhA23lsH+RtXys+v9DK8wCGb+PpMKYgv0jBvd9g/9Ig/M8SW711sZ
6TX+5kZrShqNb5OZGHuGNNkutROVg/fE2ik8de2MkW1rgtOSdEffMfFS3gQAnebT
wvbcguu3TdvdPue45yrXM1VjbQk2S0y0mmIoUQnKHckhrDQFnSiHzF6M8UpjW50j
OuKFi09YRL5B9hK0MiDxEhXORL4ITqBNeoiF8U8GMXjhYX5ZdidmyzJvq3XCGQyv
jdZJVgf40at05k+ks6NGhpAGuPtjcdCjTVFq6ajoE7rxjjUfJ+ax6r3jDAOnSW4Z
qSTH5U4mV5fMK0ktPWy4ySTjt8g8DEkD2/qv14eakV+f/PjfihbbQ1W9YxDGKxqi
NI0qx1StANTR3VhashHdAHAZSWUlfT+lxhe6/wgSDefsmpg0qZo1P1+hxBec/kdQ
a3Okr++bR1OuYRIYnJf5Rj5nntBlHTpdNub+BZ2X9/BRBIF0IWYjNXD8EeskV8my
gZMaSl6gq3fC9X3GkhtTHYJR5EUEA8JiGHtq1FzcfSaWUs6drHEWy4rYJT3yT8Ot
iFzoKCaj2Pypa49eWbDP685KVo7hswhxArHwiAUA6Z2SQ3bLufI+eNKgROzz2+i+
OGbPliOXQWqXfgdmHQjpg4AX4GEXyfAZIjsYGTFzkbamxN0BKtkJXYhdXNW6JkNJ
ao1h8iJfQRwTg4rrUUOko6UKlwzA2ofK2c1QpopZJmhFn4l3ZXU3gGcUG6tL9c65
N42FDDsc6fmFxyNF/OR7+zN65yGeQjncjh01OaeBKpZ4lLytrau8V8yoYvUJBnoS
XODEphf5lz2xdpaPhoQ7iwuVuOn68+2p9veydrvOPjJTnk8BmZU0SFl9+Tiw/0s5
ZvRsNsHbe/TxoBbAUMicOkA6Bo7ZS2fkbB+akvQqcC7WTA3xzdyH4gnIRlCVle3H
TITL35WXV+KYOg2Hs24oDNU0c64IhZuzx7hB/MJL0TbR9AU4CNJV+D8ZG/upygWF
tmyTq4BtAl323zc29bblvPSHcXkeryrqpEPW8vXTgDdmrhLcB2G1+GfrltKLrIeQ
B7tjLVAqq7fYeeZ651iFNNll+HfJFFeZeKQ0kVMBT628hjeI6tobJPy+iS2tGw1Z
4Z4LoLrL38QM5G+olJuXCaY3f3hEQ0uFhrtCviI8AjfuTqw99IC1LVaAXpKdfbUu
gfWKi9uQXAbA+peqpCFC4X/o2FxMH/Ks0Hl85JK3Eg4DvLFdGEh45qWJ2H35kuC/
WiMwRyZGAASqMiQj2wU4k272FzvMwfcEJ0sZcSssz5iVUtdG2Yumalg91SPbJcEu
W2PbXSch/jaULMJ50vZE6u373/3ncUzKrWqxfd4FI6ARmJpXinma2bYudVDguPRD
mXT6eDhaxrSV2eG4c2JZTJhy8K3lm06vvoMZPyd2JL7S4QJU1eFxcmPmQy3izMTs
xqWEtBPj40TP2cbAT4fhU2DJzX20yMGVJLn34qli4gJ/kgi6vKLlGjDtr0rpm870
R2ZaK1Zv3zTog/aqZafpFEoomB11FwXMyR/KH3oxNXOH2KvIsrcgAVQ6OKBbo4eh
H5fdOYE5Xl8kA7VjZy02d41rpdRPIVFj/x6v3UK/LgzDDE0OcUYaAczrIiAjFIs4
IanIaMHFrMo6BsIPaytlaB4wbtfbY5LiU4Os3M7ZlbmjFzvMzMdk/p0GU8qLxHCd
osJz0ybZik2ixq/YUWW9cp+ePgVEUFl1Y1FiGAtAitCi1NNG5ATEnde0fEPEHO1d
KeVX1Bwkd10WlPccAbfg6AUJZJb9+B1P+xiqPx8Ps4/QZglWPxJomBxx2JWyqbl7
1d/zcf5rrKWjflgJMBwMAOKYpuETCPD1jQNs2JHa71sVqINIrcVQbEw5ZhFtgvw/
umF23M5wKjnXSktCtO0loNt7OAaLZ743VqYHodtU5kdhiPrkB5VTh8ewR7P27xzC
wAiRmMwbQ2BH+a78vNa7hzyObhOP9hOyVSfm75t12cHCg8uLG045ZFHMkOLN1GFa
JoNX3FPwfeua3kAvHSwsFPaQEK7tMpdwrdfuozTPapjthVjXgDyEVmdCzUH1IB01
JCpzS8zcnYb5CIdpoyKSSRO+pUAYj27EOLqnHuMWCSsc6rLbmUv60xnG0RGKpR0J
vJJ/3K3obm5DVDdNW5lyFWTG7DXgLZp3/ONzk8qv+V1+iKVxK8zyi92iKVC/73Ty
ANiPQprds8BOEagvVrZgXJiaDQgIM5GdC7BB5TGEC3H6FVuJCXysJtpKtWape7fx
9fXryprCjAOd6bP8/AsAm+3ALzUpY11qTuuG92TG2q53lybsR6V8xmwYgQL4iQj3
CqrpmWIO5J6rYdQD15lTLF3fBW0cqYnsIsMlkqczvJh0HZiRVYXAQ4C3nExcVUIW
+mwb/AZHkIcK/PWSGUB4XjiwyEwcNImWyyfloONtlWVspJ3zKWeuJXQPApOfnIVS
Qzb3y3hoqOjeR7jj/GZ9oEuZ8VLrjgF+zazm7cG+WlW1iZKML6e3bQh2pB13bErx
JlTxc5NZg17Sm28Qhiaw2NZjbkOMU1U9tIlDPewpHcpW1+C6EaxxNmEajINNCrbK
TeYgBDNeNsIY5h5DRTwZI4U1cDJ6EQpPj/A3mY7ZCQHn8EnJCVpFIVKTGC61EOGi
lb8phNHUyYGuz3xelUfE0oxwGqLUzGAeYkiD/NvWhAplzFlBhi3j51vtHLy9di/h
5JS2YhjcH/nbpbHhjtQSb27p9ziMbjgWoQX6oPavaawP4OiUJ5vUMTW+6ByD6a8s
1iH2/BP4y3LTmhhXG0jv46qkefgu64NIJEDv0+Nmq7O5EOW1BooPR311qQpXMUf9
6GdLQUnuGVB8UV+ydfQFCqLP5KCPnCjyi5Ivzf/HF1nGrrHE5PLfQoRNZ3zBJAkR
mhocoazBm7e7TnM2X80u2AuKWfMEl2A3wkwU2XtAHuYGy5ouEablO2wykRMwbpvE
u90HqLA7GrIH7prUAxQYmrr8tkZEr3XZodtx0DqHzS3h9XFzc9MBmeIkxV7pevy1
v3Ix1ZVqUwVnNM1jJUx+ValVjs6MpSIcX9pE0skVA80YRCihOFF6mCQuGuhmyttt
deURvN7JF2AsEiq5Sjvt79W5BX9dLkd0YPcfv5OJeeWaNkMe5P1dfDo3KBjDTEar
ue0MWbnNx3zclujmKlkC00xQ3T9e/ja5nFKSY5V3ZTzRQG2q7RCrAoD8fokgzzOB
Tk5Piyrlfif5Fzey0AV8L65w5m3bxJonct1cALqg3ifLK9UCz2/08JF1dotUbfRt
pfVomcBAZmmNHKfbVAhLlfCL38j7ekopVXfdg4UPvBQBYR+3aubUHeMjUXFwGAWZ
RmYyQrCZc3miaqBqzE9jinM5fmV1yqbEjWszgHYGrqdXdogNS6Ny/jLpFKM6067T
LVnQj/R5OxC2PmIwBzs8pXbtOhij+G6yBCXK7aW7RV4r6LtidPCb3vSd5sBqwAmz
X+6bQKtMtK063U+yeCGwMKcm1RDLf1DUWJDJGRIHOyeOGpJQIeAqXmCiNC2P7f4F
h2qh39cVFulIO3lLOxO8RD1sJfpEB/JXmZ4K+evqTM7n9rDF2qYyoFH6GvxEg7yB
mM3mObVZE5h5gRSS6qtGj2Tmva1A7iUGyvg2+IY415NuaYMq+yn80XJ9gXW7kSvV
Pr5ethsOFqSm+F5mhTZXOHsTnMfIphle0XNZBd3cSsA3u9BPeyulnd1YNps3X8/S
SvWtJu/4Cl0+OcvcQ4C3oPW4yeky3df6BNYWXf/fuju8x12Adl4E27mUb4U+7ZCp
+vHkjyI6e9Dfmq1NHZYHeptmeFN7fe5zCGd9YFCY7w68wxjJYaK4pDHHiSK6XVZF
f4sVZL80ymjTB0npVbDM/slGoKc8wkJDhDUog3yCkvVwcnb+FzEvqWA4yRacx/w2
vVCNyN0hvjIGKX+9QzcXe2+dOSHhn3UVn1cUX9If7/9UeE0+tWQ3ws31mAJqh9Mh
ApmhuiGM+P4A033ssdcr4PwLyHiVwOH3L+MiK/JvkZ/uRo8D5n5QiqiYkx31dO0x
3BnSZtmXHlM+NJdcjdSxef+dhSndLE+UB0JZxdlf6wj6LmSveTZPiwjm60xaZ2Jy
MbNiD1nCqcjyHrP0tI69H+w0AXfqTKBuFGP/OYrgcy2sUMZFsJI/k4OnznE4K9JC
mUEXtkrHWuLfaBWQVMCQsDlq5CGClvGfOK0Gyi0Rzzbos9f0yj0O2hjbmIZGY+8v
MEsHR+p+55dvG0/MbKphWr71IW+QItXKTGCQtQe8k+D0SSR7iqcXj3Q02YqDO1fP
fWjiJYI6wwxNTcpD+ZWuPMO93/t53bT//9fJye4gxQt1hqoZLrSAzQmMobeyHhOx
iTSkQs37cC7dMk+4KPj10mat7rXO6QzFJSBuLPU+ggjJGCNB4Z2XZI/gsN7nyWLZ
QKU/lfYiIhJZVUfqEuwYvmmQL05BnFNM6hjxe8KQnuvfd6nv0Ib9dyJ6R/a2m1SD
5fy6qvd+74AwPvzojeop3EzrBfcXUrxzLihrarAA7CDi1gOV8qOTOOmMrQLXWIDG
LhAW9ir4Bb9T7M9AS6hsAis11z3nTbA/TDLomSRXWZ/t7L3INsmGBU3l+TtIH0Rx
QeGDYaicJtMtwxxRwNF1lkkE1g3rxX145PbyadT0YVOLWoStUEfnSBa1dgQvX+6Z
EA+awn2QwxWiw3lK5yyVyDn1nXJ0NjEJaq4iGJaEbVz+mD4gicxn/oGzkG6mC+kT
0bGidO9sltb05bo9kYr6my+e2EvGelu1Xa9Fd2cEdy+yWuI0x+8Zq0IgiBOLY411
xOF2AsuakYBmj15UZm6etWT9hnJ38sMGYCGzLIZCSYBXjtIeUCWZgtCpH6FPib7y
Z5f4q8mYY1Y74+9uGSv7vYo9tGQNUF8nDMBoIBIT2xZQzO93CBpo/N25mMn/zuh/
ps7NMls5u4iz/g8H0SNYpdJ4ghiPTrI+ZQAXWBpDdmEdcSXGqvrou+W6nBhaOofi
QvGvasP+QsmHsJJoijr8/4lahvcH0QfEf5Frc3VrrT0bXHi7pLulgwF03sC18Jr8
PDEeddEz+dxq+Ue34l7mp5S4XnhiWuMIVoYOqUkyKvaxTWNJ7bSNN3530JfOglYW
nytXlUdmQJguyKtHY0voqqL8pgnqNo+qAAZjPW54DZ+9sMMpYIp5kMOqRm+WObBu
UCkzCMPr3NCfPU5BaFOLxvhpTPAkIZzihwcXIxun4quYBVehPXNDT35p1imfooG0
oq77EjUpM1midoDGPtvTd9u1X/Q80iRDHjlalH5zAJshfT0/qKp9q4cIRDCu2cc/
91W83jyQJmoRpTC7ezz913CKPmhHV863AR9te56dlgFsmqLKdQhjVbCmkrUEWIj+
jHT1KsgDvd+/cYsgiSA08Iz0Ln5AW+ZjBVmcPUVrTQI/fkkeirPrd+zNi0MKZuYr
wePeNx1wdiCQFW7knCacRD/7eCDbL6A7gT6OoXVz7uJPdjWFphEPgQjkbF5O6udX
z0kgE0r97L03Ucc+T84tv1dGDP4zXQaxqsuvYJXY1Wg3THAGjiB89HKlGyDe/RX+
BxdyQJZujE1i+37NLIOrwqyzfGDRDayCRHLWUlkXv/wQ/BpYyyK9c2LutasY1Wv+
sT8McKmh332RxAE9lLtbIdUHpsPzyyU30jsmX+P150IccQo+liNDy7Ie86RL3OIH
/oygUI4HOhhQQHEZGPRUPVncsVdeS0eUpLT7WuYoWjpYyMn7q2in2leu8YtvPrN+
CsuCPX9z1bqr1pN8GpUysL6TgbDtORltaJiQk+nAdo5xCH/zaxwsP+dhNIr+6mpb
sWqXQBUJ8LydV30qVBFHUB3AqszD5mfMj/Fv8MncNei2FFsqaMHSmMLhXnmRapcP
mrQfWd/HkzsPx9kwczyFxsprqiUJNK8mp3h/kXXoyuS38obrEaKI4hnOK5xE/X7t
dc1//qDDTDZUM+aIFSLhH/3Pnuctz2L58pdDt2vztLpc3NnJSVZotVMZD1W7aQP1
nu5ZHzm51kG9dtNMl7t09uY/kvqWCvBfC//3R7ca1qMV6TM0+S8qj3F0gIAAbG59
TZKnOMwjpYpHGxRZtuEEZyAolD3Fx3x+zH6B/yq94GxMkuVh52omS3Nc/+p2gu3e
MhWKGoMszHv9tD5WsV2FpqYYgAnwDwQJJUAPTCO14GFCeTMpFHVA1Yaud9IDyA2L
zfOl8p8o7MBsrkcCGUwnnw66lYCiOtzSYJCwSyUOjT9BW3oqJnRobCD3CLoFbfEK
/wGbDs8JOBx99LWTwY6s2rtxJODCSCjJBWo5KnMOfQ83TGSxq0/5FrZTpTuFw3LM
q+dMkT4Sl3KH9z+cfAc84rE9Fy5cbY+YAiJqRC79P4bENBgA5+mY39fy86wUM+RT
voIwCjRelEvXvGjeN4MrCUTM6rtMlY6aMwDSGc6bACVpfIs5+Q9gg9cNc0V9+Hss
ANxnwfXZGAc4exNf+vZ8wQEEyfC+MbRD9OrRanrctRomkKMnC3UFHiHPH9lueO3Z
A3jYYVNOYGCMfy2zhNpk1iRbpxIJZoq8SfBvwLoQsNmFby2X1Jo25+ndJLgEm93u
vnVYmj2q3QbdttSTTKEBqk4AJblZt8Jt7/V44CSRGaZUHI1QPjoCKtFiNsc//467
yJ+pQ0klx1P/Uk8Y1ZrzN1cpXJhoP56JZ3IpkFjDrayZtBoeDoSOFgtWgtcuDFr1
hW4Aj4GFrc9Aw4UegHJnltC2RdR9I6NRg786kvhZuA/8HXmpndN4Thrptt9GcLWv
KgFFdXVE70Eqtq+l4je6+7+/iW92zfdSfw+0F4WBHpa02hCyeI8IeGSNEse590xF
Xe5cb7Eoe50V5YejY738d3PIEhqKkQkC4wLaFN6fgGN9cKGRWydUhq8iAxYydYKl
JISvfGhW5TLPLSUbVaH3gyNE9KNu7SPdElWmLsaV75qH2Mv6YuE9DSxmf1GvetI4
fU6z0QtoBIJPdVgQIjGGMS4Dxm2onhXtpzbWJvyRtExLiq3aWkaGrp+TzooTZ40i
X0ElMv+xxZVA1FknmQRW5x0sLksX8wl8Norzd9vrH5H/9cpQjJ+A1N2ZUf1y9MDB
AQIB6A6bBUPJSzJmB48pOFjAet61uUVzH4fNErsYCuot7VDV9EPOWivDrM1aCvzi
a1Nzst/sgmmlK/lrtTIV59qlhkp+HEonnDhgmW7MIB04djFUKEvGwTJyRnFsI98w
Xhcr+khq9JyY1WNVUUgEQXR9lxSNVJgyMBSin3p/k7vli8W+QtzPXB2sDEMcfdBM
9tS8ygUtHJGQMRtHxiZG34AEdjpH6r9HDeaBqkaSlks6N5cTwDWfHnwBtILkKjwA
3kxEobvliB5yr70MrBjWl9XL+HetPF/EeaoZgkKlkJUbgEls+z2PK+UGcWnii0Zq
TSJ6X8rqZ12Qcu9i4i/z6fsl8Nzbh89dw0Q6zgK1RyjlesCr/nPhWx65bA09p5nj
hupEkWU36SjjLbMWt8+m5PhIzbQvfQ6SayvwK1MYgJa93fa3FRadx0VJpeHzeNZO
WqhuGuUHnZESrN3EgtgTtVEZgeYvXis4oTdBkvUsUS3KaH0muGR6Xxu9eti5WS4R
N8WqaPmemmcEINK1y/bPY9tl3NIupRtfSeb8PY1tisq1zYLrUvApveKjHlRGCVb0
UOTr658NgpJJlPgjN79QqW4jGSY1Whr2VmQ+3q5bi5QdkNZNJ3NsFYwwJb8N5lDV
F1vEwR9WnQBkGiWFl/5+/qC3vhvPWY3p4YVgeG+Lh5MTWkbwdn5KuKgqp5q47nE4
FnOcD31C1o9NbGD6Mro8ZU0YvKx0wh5S987KtsO0ubZkzoGw4mMs1bp/i2ce9C+9
QB5AJL+j9Q8jEvF7DNxu+5G0qj5SJw7p9LZR6oBF0LCfr0WjVWkyHyjXMz3xc4gx
u9ze1XSZF9QUEnhlyp5eTqrnEf1cDWV01XpV28Yn1TNcMU8VCbE3UcW/1vu/9AY/
vPeoDSxClPQTGkXKK8XHFc8j21ll/1s6aGsWNFBuNr8/VrTRN6bFKydOV3YD71xm
Tydi7vNb3GgFppeH63THU0bqfRptYWJ0A/Wlp4gbtR6WQGvW4AENMzy515XFNki/
GrtoCbsl1v8eFu2bkqK5GXR7sqDvZTOeLz8E/LD2InyUPuRQamSJTI+fbPtz6xV9
+cjl7L97w6VoHZf7a9EBWtvjjOyHTi4uM9uBTutGBlkh8VZlzAD0bF44de08qxZQ
+qYHYAH27jZNbjsD/BWcwlTEvkmhEBgT09lRbMxHIjIp8NNM2vDD2yXCLVbTl2FW
T0Kxby2MXPU7AKS8cLdjq7ZN3j1h6gHKpfVK9Fw8UE+qxHH8gjCjnpqs6lNXpxPs
7q4bxqbewjpvhZleVAShbg+20FVy0nDZtvc6g1KqAHtTMOrJdyXCk45yPLvtNxYo
MXhyb6fDwfiHjHS+JqeGsvvnAyXTVV3z0jULnctPK9S7YF8qI9mOXGggxyo6PKZL
gvQv0Ft+RmUxQ/2zo2AFVIdOJlRKHuyiOvsg+9wlVxvP0aUvVIZpQu+WmDnL1wGL
eguIf4/m57BxWjhtYEGcP75ZuoFRMu+FyyOSOJUQsKNGX6dHLmwP1gLe8M/peQAR
Rm5FQJ8m0qNKP/xTLIWjMhXJF3+rTK/Mff63EfrIKw7AF5sogNEJfe/xoruFUbGQ
i9QkiZulDG7N7CFbtxg5GEjlWfbmx73u6VkXN2AkDySKnkFY2UwROsQyPIxKah86
bR2mutrzADtgYcswV6a4LzV2A4DvOIsiv1mtASvF0e/AVhVjroudjRduWOAxjQ7M
6v66cG5/3XxOuOedDXLCSnSCvwGai64p+rM/sD7c4JoXCNBZ8+bGcGPXDw6VEZPa
xORsLIbcs/edxb6KCv3IJm8T3ZXbMftrq7u8j2C/hVxMgBdugQ0KQmmd6Ovf2Myr
cf7Rgqtew/MJOes4MN71muoLvmxI6DyuMNUBIP3gA7ndD8NvQwGVhMbMVA6qcm53
cnYIUsX3NoV551mKbefiDGJ66Ux1TjGntFkl0IvL5V6tyrOp5NgV/Sb9x/ws5rMA
f+LHppGgopNlEjJNXzE0WR45rLhPvlJj7us0rM5DHkrBHjq7Lrxohg38tPeERh9e
/A5jpJZhPbGNnRjPOeUHt5sqXpfF1MVKCCct9qZeTcdFhPL6GmImC1Q9HrC7db4P
UWq0FsQ5niz0HX5+Kc6v4VfgwPoOfwLIhMf92QJuhM3f/Na+o/yBw3SaGsp7nU1B
uG2Zv3SnEfABBPZZVOIUM8T23oKU/QvVwGPYmZtjPBpBIKJokTJ3wpm6JkOeRv1q
8VvZgY5wHSm8rlDvZiRUqPiZNw1cJROZaPnnBQdv7I+U4Wcoebd8ye1mt4R2XpsW
v15yhQKLLzo7frvovzNjtRPl9HGfi9ainI6dIQbjVg3Hh0SVhDVoO575cT9A9dlW
Wu4sOK7NcRtzx6nGdzjcaPaZr5iAoPQjJCfU3sNxJ8G3jHQe1R5iiepU8LxRNghn
mHMuUYQqkJ31IdgMe8VqDHbg2FUVv4p1Iozf4xn39OK1iCBOZNoZWoh2I88WVuVv
YPk3ZGIYdLkcPw+7C1J3UE5IfejDGcpZUul4695fsZcTnEpu5VsFAZtFcs+7ys/3
m8UZzVuphKOMXsNOYo5xzzbZNXz/ceo6gZAsZb9Eta4AGAwr2C2gCmsQr8YNbVdJ
9hokXohjyzxSBQJ3LOpO5QoN2QB+02LXI2V58bE7QJPd+cBTSPJfsXDULRohEx9n
aC5SvSeboZ8Hwae0davwNcE0bzVZoUwqm6TzeIUBgIMfVIfJoTa1cO+Q+n8RbNDu
SdHCjytGjHZAL9xxd+naUydlI347jLTYUoxmoXV0HaMZ9TyIrGKjuuTGcFwHL1mI
W7y7Fe3jWY81vYsxNBjiG8Hc1awzoG1P2BBQe68NUodFazLuB6d6lmhMR1gjWyz+
xo/SRbV0K0R39zftank6yH0A2TmZCld/StN/C7cXL9pDKw2uMWGfW3Ed6YZQeRAe
oLiIaehuRUBHmsx6YZlpv853pM9CCceSDRr6l0yG0+AvgdRz6OTygH/jCzGFXUMb
xFDAh6Ap2vrPWHfVwouapHqhs9Cn7hpw6XHgFvgEobq3IpE5IwNkiw0yBRQHZVN7
DnaaEwSa5AzLMjHHVPo6guDe4oMJ6HlYhSY/wQnR71thjdD7lgdJibPIuvPBpmCT
fno83fx8tKH/CmP/1ApylZL7X3SIieSkc93oIWc3Ryt7ZW96Cs3UH7rGkA/D3eb6
0ZmM4ePYNoP8GGJwyTZ0DnwCgq558fuLmS0abwYHvRwOP86i4Nz1ihJY/QhF3p70
8BSPrncBEuiM0hMGtAJGJjAqu4OxsozBSVhRqj5gRTk5xFiDhOjsQUeSwaS0h9vh
1BvgjhdKJNgf7AKg/Ih535iLn7anoANBaRgcMU9bAe8OCSt2jSr0DY5pAUT76aba
dBsOzRxdkvvN39dzyM28B5b/4Xw7Zx0zhdLtJng0Jggh/FvSHekVNhlcKZIgeANH
55Qpe2R6YMcyqSWNnvsZAwEwVdkG7FWOmyV8GXTGCFP193KmFmnq8Xdh3XihuzoR
9KY6oGstC4BQvPPGeqq3hH6sOEhqo83S9RC0crfQ675RTy9FXyWS0cXPglupNnri
cMWmO/MGrAzDP62woMqQLOybohcLuw0dSZ/ouaYM+8xFJ9ziNxHYkp14iriD0jqJ
ZR1c33UX3rd5xWl2ZVP1y4slj4CQlFVevxlb/datPftD644a+2FuP7ALRrHKd9G6
zsAkaglUFa+prKKDXrBwTjT7In3dsUfPdrFZGUl+YT7MR9tys0PgL1CuoKMq/UjI
V5N/bPWxSuZ1U3Y5PX5hl5QY/S2csixRHWb4npIV0aQh2HOdQe8SUdMHW6k+KObn
AzlXqNMd5IlGyLrjjiuLk2FEw47cKAKklEuwKAAk7DzoxMCb55Z99pPbb7M9wWRC
EMl3D+APls0ztS9q184OZm5mUy21uzTZDgFWatcJX6YTBFo+7sJxT7YWbpUTfPkN
N9cb2+/o3ZzcxgohVdw8UwVWZFenOoq+yrwyXfNxy5t1ZYVEypUqwxdqMRx7y0Ek
nzp6GsMyOfs4tHB6gZaWjHP++JMDoipuWXI/6i7kEWxRgBmeF88ZsU8Eundp0FYV
bhehNXdf+vxNfnN7Cate88zrsv4AHVptHm8EAneRCIkZf3s2NZuU1S89CoQw6ZLI
V2DiXGWr7xZ1OadRGwqNczJ805cTopUKoVkMljlPXE9sKmfTJHaXy9LFXKqdzL6E
Nj37W29H2jlexht3fiR2q3L2o9t4UaUbeySaSdIfRILsJlXJPPP+W/UBmT+SppzF
ymq9lnphbPuK3yppeYNqDx9N/QPgnPqj9oh48Nqj51Wrh0YefXzGu5+dcU7o+E9X
qE3Rq/qtvDvbG/+AWvUSPlkxEGx+SLB3sbOXu7GL+2vq8yb48oadeOecsVBJY7cx
jy4OtE0KT/cvbPLwKWyFfCmVVlOft5P8QLhs5jD1K9zYHCzA5+tef8GM2XYrr1yS
XWv3YK5x4zG17+qxE6ck2dIQorrmhbXpJ3bYmKwVbrTN4Go1Lwmd8QJnAM0RTTxb
uTyTxL/cmkhFIbFB4cw2+R4ZBZ+LN8G/tBjDWA9XlFf1FMNDXlP4Z0GFfSPOyXrF
3WTMNxZb2yDxDSm7wzFCpGiwo0b0A7rq9n+BY9mzAG+RpV2Hf7O9jGvjgCHbWRRL
G0f4d2Wrm2PdlJWsyxFrsAEPrzktM/qOVXeUK+jRN0pVQdBTpMSbBpdpQiBR2guQ
JlKqM64bC85WTdDs/0ZEVBzepq1ubyJe+PmDos+GpsmeFwwsWp/R8n3mih5fj5hI
s9/2ta0gXyaa/xdjw6V8O4YGP0vYNws69Sba30ZubnNHgruL2HcAsxCgdjmRUTbc
QVe2ZbfGG0GGdXc+DsSjDOWdLYPsMZr6YxloxSYzl2WV6AgK8ivpyGGSVpeCHW69
9P3O7ny2r6tmjDYlerFM4Exp8pb7N30b4Iu+kc5Tjqg1n8jygZEuz+O52giaCc/I
++y83vc3MyLBRx6ilC8WR1HP5O4lAl+r/xIBvckGOK1oHbDhAMxpGoFd8usm9clW
TAbIUvFt6H/W8yWvzwwZo0Btuccctl0RHEoQMwRrrJ5JLyQxTsuISajxUT7VlZmh
Wa7d7s2rPamQdMGGQlx6uG3KAFg4CJfMWo8dOz8zeiBQB0vfisStxDEYnK7XWNyK
qLPkodjAVVwZrn3XLW/j5xVM5vuRuKd6RgyaPi0s6VXzzx7WX2AiWB4PqAFJKvoS
RyRvyHoXp7mItd6KRZoaMtdK4mps0CTlBgnbcQf5yTf1patbUt5G+WMw22kqJcaY
TTJ6BPVEq3NsfCwHRxPQwJvFvW1XtPp8HZ5EUAN4dt4LZNLe4PqqUlcSsRkYgrtt
oMGD5sTLcvvW04+52ht2SwefegkPZHtFz0A4h23TEgC6U/odrA/Dhdkcp7pVgsmV
ZNILYejE1QpX3vWCf10JAsAn8Kxw6mSqORmwes7bEAGIYrwAlRcm38OSZ/GJYrwf
z0kwMH40ZTzP5erZuWVnvCm3HFIf/AkDcDmeKSRK5GwOpSglnLNX5RGacMjRHVMw
QuaGgg5znEr51im9WHEl7VPRfHvlegEUHqDR+3dnNPnZNwKoaDoMuBlppMRTxLwa
emveYS7GAYClvjrbgQz4hQVkYPPvVq5FbApxaukmiupe41AmzK4i5QzwiKfPbdKV
T0kC8X7DXM5S8me2K9Fli46vzPzENX2I6HItY9wWAZXzAoQqGUT15PL09DVMO7+Z
rj3NFPq9H3NJqLSHTV0AHinYdL2uokzD9llk+76SOHtTshhZlB6FsXfndDT+E86m
SL/HWd+dFoEN6g8RnDOEvGsoq9XXk60Zp373cMlWFeFDQHbdmH96JDV1fXXYlLcU
7kR7Tg4DaavJaLhc+eSQpumpXcmglqsidaWcYgpq4ohYX2nAxcjC4TqjaOwu3S19
SuOIFpOljybpiqS+r9Wvosnd/0ijZ6axX0eHspzoZo3Db8v9B8YiBYOUO5ziHewT
RjOVGqFpcdrSVGgBbYn+ONCcAB1gLBashPfZZq2R+we8mMQ9JFhG+Z4lT94HLsVM
gTfeeV7C5vpeouSZH9W3rTr5/5MdLnYiBf1I+NL3hjyCX7tSnib7KVFkfZRupAOg
nYZg3WviaHJMob168swLlCPi9xWG38aUbyfnmY8YXTjJ+tbZ/KxUZZP56czjz7PI
K0SDQyYYUysd22sTaEfRvslgjP8PopxYpCpyxNYiy+EJNhFN4p9cirq5E0nUUii0
ElZWt9HBIz/I8UTewiMhR3Z4mAO5u1s2UlZZB75BkSAM1x30nYo6qM+7T2TQAWP3
iAHUxg34PBzUEG8xpAZvAA2wsny/EgRW6b05Iv9ONwPmAhtSZI3Yd4G1NvBaN3ox
QH3SSN2mj2dX5D4Zex4bEKGQPdteHM+0hmygLKJYs6RUEQVrRNGV5TVIQiwe/74Q
qcvFuRWZQQ3CtzKBlh3t6USBhYyLOR7i2M+LB9B23yAl2iO+a6QENL+0+hgCH/5t
MREsibYNepFJ2fxgvrQpDCHVSTDQL6y0+kCXzfEiB5nNQwM8r5l/qt9+8cWmI8YR
Jy0Rx3mOW7/XDm4SrLo4paoL+A/i4E09goDVyOPn4wQ9UCaeCos/BChdMyK9sBQB
IPjDtE3by4XnmvSZslW8cLsiQV6R10VTB0AodWTA33ARmmt5VqBhgknkldHpR41S
uv2LaRPDIMPMKTSyJD2VcdIy3Wip4kGXyf3F7ahQswBrUHKyMwLPs/iV6J/n6EzV
ECeqHblJuJ752PC5ACsFy+z4fwhZhzg1cWfcDXGLKTDLxI9H933N811U1X8wr1ie
q2ti8Gq3CeI8h+RkBlkf/9OxJZnD9+sn4mHncYlvKPx9Xe/GjddyVd6+ex++lv8n
G6iKB4Lf5IcbWP/gXUHwWUwhoPKdasfchDrqWa+Y2IGF7xGeK6G0bBWKe0q93w3T
FO9cGNbs/jQ2w1875b+Puo+2ogX19YbzXih1MOoxFPsU38FYKGS9p3MZJ+9Y31Qo
gQkUN7Cee9UVgwUhJX/79yGkjb9NDVvf4uvVfjZCrKQEZEjEEfRZJJvFMSoV7iW4
PDcqhGB0WiYsmlM1tKi4XuhnxtHiJurkoYy+9fEYNHDG/O/mxV4DYilGuiDtMfvB
6Vc8FI43F4KvLrI3gxrW3XIsTpgSPz8P7URRxDC+3ae4hJh/UspewpI2Y+68dADx
9W+lTymZwUEzliGezltHuWElK+DvZ3j4u5d72CYlQaO8/HUy+q3K9c9h/D5AN57h
mCSJVXT1q+a/6LfHtSWowg5yIN2igxTrknzvfRGaFJGq3imnzKz3fyrPb80Xhh9I
YRS5zJ101Wqv5qdwtsKPxd46YfZs9+qUKMOrJM6XtqoIZwKbtrODjiiRA727e4hI
zUWKlL0/CFkYv6o/W0BZqk52mZNcePgisaE0pnPTmclyfgS28w7aet9OhaWo656i
BE2z5obdTB7oSb8MSVnLZWu5/KINKE8NxtVPWFVY6U8MRKmEZmjgbgvC9xXMpXfS
e5oyEQJJEwVBwBos5m4n+BCHJd1skk+ooTl2OMWm1S9B70gw3a/V1uarcKnt++gm
f6rowS7NkCUD9F4ubl1GeL5ftBaedPHBOiRPIbrh83cRp0Jp/NobBedFBiZngeXK
EutTShpotUTx0Jl54sOU56NJY/D5JpWQfBL3N/l1rhulzscBpRO0nVQmQLazsETD
pzAZWJZd6/6/MTIwbQ/BIcj5obQN6iSEv1lnNScGxjMVrdshgvbifhaF7DNxZjGn
Wj/vNQMV3nOO775Pp2WncWCpE1O97LbsI/bVHY4tYAXtdKYDhuo3Ga6E57tEc19o
1JlKTVPRUgOhg6OVLSJWtWh+VuTvCWJFopD1SDTI7HYS6rXThZdmjABeor7Xh+sz
pXYcuz7UEAYKyWjohPBoFVsb4HjxsMy/KNKg5JP3dMejuDq5S4nv59Szvoqr/ZJf
DwLqykGSI7o9NebOo8RGeW4ip8SShSh16okv9c5BYnyNn3vID/FUmPuvS3kqamzZ
AB6m2+Vynl+Cnl1mcWxwryuvByIrQf/yD/ybtY4InoqYVprnN87Gz2sAGZ7WnJVg
SLmnSRHOr5KzzH/QpUpgG/8W3o1dOmDmYcf6ZW99DXwCrF4URTgSewX2c8pbLf9g
Jtl2UatJtBoXvBgA37VscbKcJOPEOxYyggqto712aaIN4mcmFCXcQ9ziAZOLomYD
JzBBb0sEHKmOA/gL2rZzK0xw7jth1R+hUCV3Yqe6sk2Ip4AsOw8q+L5Tj3Ppz6A+
fAFfv7tY6SwWl5IwPel1x9EbOUioA3HMsVHaFlvZNwKcA60rBwEDYMuSupL4q9T+
yCJpvJCH0xoJL+J+3McCudeg4dlw/QZvVptubrrro92OB5Yhx55gQ3qPsNNWB7Gd
4zv/CdkONW2aBtJ1fWKvQt0JcUh6P+ATofLz3NnvrzL6jVW/V7G9J7LJjtyphkL5
tMme9wcYvcCllT/TNPFNyVPMO4bDv3WZB0nRm1YrasAKVYQhD6qrzhw5sgywMHS2
kNpSVKk3IvhWh4oUswv0EHP7CSPYzgNuEdXSfbdEMxnaUGyZUJN+Qg8R4Pd/joAa
xnPzS4YYqLEVROk1rDxCag+V00/0E3k+e4wJLHgM2UNxpeIe+U28SSo7WL9q6EZ9
Ue6BxKZTep+B4mUWQeazO3waU7xiebsDg+D9x1KvXWJV3DIZLS8TmskxoKu4IVW6
eGjn0OK26DrisrQpdtnDrU2QgRH0gmvlH8dixNybD9Cnt6X+E1Kf+5Nu+JbpZuFk
zPVx9e3lxcDFozNQ8xdbHnCjjWPF0KAdwAtb1Cvlzij3ZyppgprlmKAreN3TbEgF
7RT/e4gTZPUTB5wpxZsOkL+5AIhVHMuFaOSZOUQ2/SY8udYwHeSMQ2xlwZgOZ63t
NJIHcLHHNqvUfm11pClQq7JqrfO2GpE96NI+YAVehNqgLYnLffwI3KfEuVBZA9/x
/UWeQZJ+slZvC9k5JWI7NSfoE6rC59FoRm9gJtPjuber4v3vV3DWfu3QHujMwMLj
ROqgR4/FOJxdgJJ8hyKpYZvpEe6VUtlERQS+Rb2JhcNmHftHJ/6oHSDKJUIJ/zeF
80zDh82F5Avmg2GZBpKBWWK2DrFO5fUBQEcX0hw/4QAbRB6zZAVjvMbHvsyf/BSW
QKtahbTbTb2Dhkl+miUaAlchWJsS+LQXuoBE9UCiJ5+87htxKv3/oOhC8R8nL9GS
xAsR80OXGVmCUj30Vw1gkz9y8mB8bx9ARCGcQjYuZI1X0gev96rvlbsgBGGEFCvB
pKxM76etseA7sr/P15LDo+VDdsg8A1xnUt/akzU1zM4s8nNoC0jM5jdTGU4w0dz4
4lCZgHJntoVxi6rkNmUOobbCEQuW9+ExfruIOjxWcBmzy8D4k35Sene4O+1d/C7L
HJlQEV/9diensQ1DHp56OG0NaIq1rsouAJSwcy9KPGgNGd+XTIeP9O+xgvelYpsr
PeQ5qG3LDyx5oYtrGjBK8VSLl6Eg+5R3wOz0cyw2JAr0NllvXxfqn566Ui6YTHrD
w7glQKd06qHz1+4OlhLEPilsC7TU8kKxUgTCB8M0ZiLP/j+xDOziuiqTnXx4+Twr
W6c7MHJQ/sf9VWefW2YRIeTsbxvcOvMKM/y8HGhfCrsZLS5KM04uOCZ3odXtob6N
/0hAxtIegiJuaVm4vuix8xb2bXPPtO2PEPueB9xq5fAtB6+MFYR1HKRrWDtJ6W9f
K8ZhjBj2b81/a/xV0JofjQU/FRfr6nR3+lkMdM0Pys8YO7XwzbISjBrA+NF9Ad60
VrqPAf9lhJ9TxVonMBGn6oada9o+wstSX/83kPSDyH0WHXXzgXrrikMumEPaYu6x
Qh1ejanUQBnhbTYpCGeeg453XTNV/RiSWvWsA/0vfcBeKQXYOsY/B7idnvRNWjdg
iI735q4jnfn7XjWf//35AZHLOFqyW0T9WvZgoxhFtqEv6cP9rW5bZx0ukCFQBPWx
Cb+sWzk7CnpLpz5GrZulr6g/VUSsFmriy6kRJnDXKC1BFbmzLXrOxe2iCyhJMbl5
8Luf33MR+3fhohQEdGc6d/Ul5CN93RIXtB+REjIPqlEQWCGZU35dkOhgjFaxcSKo
/O/DJ7K4VAesgtFb8h0I880nviUVEr5HChw2wi/uFIMIf1uzXLE4caZlX/toV1b3
7g8ZKKluT2M7ESTv9pKwbnlOmi59LgOVYjczJrA9ulaFPwZFGspUA2cgdKnXB7Dn
FxdFXyocgVXYmXhBl+PZbhavk0HPwrrJvR63aHfkb1secxkwEH6Ky8WCOAg1XjRB
F1KdF8OUlSvTRSQXS9A5TkjRlmup+cElyZQd+phmnk1BIdrqF/LDZiRMSvsD/f0C
izM6pXoJjlfAH47QhvfE2mQWiEzWJJbc0p3FThrH58EkHw5DDcKuSJJz3scMFNBa
eLz8thNbgSozlsiTcsXbvyQ0or7UoyGbaepCAOy6i9+5dYCS77hWGYKyIhQivNp2
PgP4E7RiNpYtkdiUZ9U8mGUMtJNznWX4/huTVGlj6GFrUdTEOaf6pg1kmHYB5BiS
Ic1064itvqMCGXvfDX05xicnVg06F8pNSikYWbXDVpwmHKX+rdSbnsaWbceYjVSg
Y7iVXTNKR8NSjGvbE0A77CShsfy7xeKc5cYJk35Wcs/9VthYGUamyR2lDZcRQQvA
kzygBoerNLgtnP1x+EYhwL0HiFuNArFiYR3mQjrVVvX0qWGOvo530QgBYGtC/DW7
TUrskchlVeAzVAutauLTitBPz0GK6fK3Y4euNK+CqM/Py28MUe9Au/OXyHHs0PRK
HLMe7qppNUn2ZKY1RaLCviGlAloFvkYVg+/RvqiQZujTeXyKqhxKpHlEOBsUKDAY
T+GwfiT0t3rwnZ86fg7cNz4m+gDdcmfJLcD0B/aMoY1Ybo23lHS2QXuhPx0dkMSM
35GsY53bG5IHD/6LvBwuhN0hE6IF5GqyvrlrZ+2Ud5WzAJgcv0c1fryAZIFvuqzp
SABSjs/O+9jeyuWPo+ik3ri3GX3R2Ifs9iaVha5XZB5WjGtgyMwspJS5VNqUWqGC
7XHDqaOi/fK5ISPX5vcYXdHiTgbGzbhrCAemKrHL0TTMJlZ4koKrweKX1n0AIzRK
4RNsT91wabqaX2ch5g1b4zTG0hPLkLWqlXK2lxbfO4HU3ApaF5gklXM4Z4aUT+2i
Vzzn9egKmb1RWs8ZEzbISVnm5TJqjmAO+3Ev1i2v6mguc0+36HMo8J0atWSArbA7
iiMfpEXnhqE9SKzdfyIYz8iGknM0rdlIqgdHKnWmqzRAcEQ8ov7X9q7DNNgafMW1
g/PV3HaxqjL8aSRXvtMaoAQBV7Qehegf7MmeoBpoqGDue5sR6npTcoE/VHV3vh8Y
rNS+QyIaHrITLw70WiEg6bNNdGKNV/A3oVA4ithPEkMnvJJ36MejcYLB1mYp+yGH
OOQiCPzNzXix/P5P8nTPbDwiVxCIGe9fViA+ouqRvZrwwDbhcZNyw8h0pV1/h70g
i0hL9yq0YJ5b0JFITrIdppdbDmGlXETGjls9b+ARJe2Y0zltri8bXMJJe6a/H6Dm
DB2YzL95Xh8BLT8asoSYynyM6kj6MpDj/soi8/1dE6sRrkpkAeXdD0tWlg5Aojc/
i1AqH9J8ZHTuK8+q5K4MIh8l66tfiXnqxWqsuLOQFrqX3o7oqcQM/fQUwDp4Kv3r
YOwp2+1zp8pjDM3Tnqhvf5tcfS8P0o36dQOAX5FGCX6B9k08uBHJfRxNBRuCwjsX
cKGrseWYhDzPq2Ndt3I+ykfon20av7xXZWRwDybtn+1kGFX1RZWsaUVfwA+41BQ2
O3AlBhMx5pw4q2RNdeynlfsUgELNLLbH1Ad/HrbC9y+ATPodjATgOCAxMACMuIAa
/LOqsY5/gmDypreYbKWJA8MZAd+SXBJUmrBN8g8avTAJcW6oBxEvnpL0eNkQjOHm
rUACNv5RW458E0LFAKnmoX/hmUV+/FtKLYRB/++YMexfxVGXnrc/nwqUJtP1oUmb
tffaOz/dXLI7BqphmSHGo7oIi85P4hm/RbHE1PnJU0QMgRcM4Mu35lPvzx0ivjS6
r2QdO0iPPXaVYZFQNM9s25/VBvMse7AvUIvsAzJc22bjHE/SCEW+w7h00OOvy1lP
aUJtvQs3EaqaNqUuM1AVNxJDmTFJGidajicFhx8Jq+5OI9YKKVYlGfcfUt1ayupZ
sauXyTdS0XEikub8Tiej90aCbYZ7/EVQo+7dXNkXERPjikR1PmcLcBilkOab8RRw
F7Wz/x5lGB+UX9FAP+OQpqDqNwRoj/M8DCPsqrL2ZMXezjr62Yn+UJwMSvnyugte
gNqcUvX4K+AnczMgo74Q/iqi3zyDlxG+N5bBqVvyl2cgYlJn0k+fW9W6QB1blrX+
fBG3PcsSK/zr5PWOFKzyP57UtARVD/BGPS9gHEXY60fR+2GpH5fzKIFsyR0/Kbw/
EIU6I7uGDiI+clFRTjDO7FtlFa6xKFl0d8xODGvOgIqzxsu9hoOY3nsboNDnGs/Z
F3IpCiHTwYNHrM0a+cE1JKnBxktFUrAFPxRhGMpKeLZKkl9/91cT5RE1jgeXDE7Q
hIzbyKcLmGI7rJRx4mRFazif+aMZ1a36eA4mCkFxHR/WmRPcrbyeqL8M+ZBSmy9+
/UZ5t2RLXeJb1OIlpaU2oSsIRUChe/aNCmYvpoXOd87myO6AuaMotOqQZXcM/C/s
49p2gKMpBTyQSqal9fJU7LjY0eDtosYJNYT1SQwPekAZq1JULTSAUbmd+0i6tjya
LQpmXrVQ9HlXQM7ju85/RA7RqCiSP0ZFQnjupi/FytJy8Cu4VVd7mFmnoXPbKFLD
rm/2jzOVZGWn2CabEiBePBgVY60Gl9uKwQo9cKkTFBG3NRPpZ5KrTq9tAdyPuM25
UjN7+VhyAavK6294SZfCFAXOp2NH5PqC05Kb/d45QZXqgFdfjmcFfV50k0ApAsyS
mnMlMLm+LJSy/sDmye0ERfO4cCMHPwaE4JUq+jRw4nXw/lYrS15Gz2YL8i4YyBn2
v8sStaX5y6lanDRC7qqp/WicgEoRGG52Ketevvn/dBA5fszHb1nN6siHZqMNbH33
LjN0HEMxJJpz3oO0DEV9+2HjzEEWvRXapUjPmrcCWxfmO6DCqVu6u3IiJ4s6Eh86
T3eRpUMt1cXe53lTNG4j0x//MuMhAEXX7r9vYljH3mpMvbbmB4PmAHg8XI+T02Lz
8zBa0w+IlI41vKilXZEzie8D3r9WkGVENry8WJZvwV0TNoK85APi2oAdZxL/tzYY
O+zBhien3Nec4nVywSRjxP+TRJajH3TSModqVxDSrZiO7QcGRK9yUm8hCv8pXDc7
/xv+4BJPAFTAbiB2vod08/X92CVueKBjFD7MxIdorti9d3EmuAnLTc38nXINaL9T
Y24ENeFvB53qUrc3XIVF3FIgmO5j0NO/k/X97uGVboLvKQ6baRKzalvZOkOo2mXT
ABhCZUwW8FLz8k0yHofXABCpshsnZyRGbsHjUT2GOslhH0hB88gYudSxxFMQL3lv
5VQnhksUTu65tFjb4XeYPowxiP3aPHzmTEbKhhc5bU8bdZpK+7ucOtJkY0nK3cNq
4/PeraKS0LWhJiBFDYuQHwkSVTgD2tACh2NuAhHGmgtlvI8IB2saBlNwW+bCGqY/
LVYztgwkXhzi2WjJ1KCmH29xhj8XVubgoNHXC+G9Oa38VWI/Os43xsUNksUKlj3u
c+imcTuUMQhfoDdOLA1ZWgYk6Xs91dZXznw+EhfdNRMbCvutTDiphbKgO5rILvKd
yTIFB18pRNTNhhesB2BH88iV5yxWaSOW7kG/qJ7qZg4ZNeHwlBP4KGp48//VWu6g
4MQK9HJp4k+J/dsLj+Gv4K89CBSdbyui33B8HLxPHOYEBsID02ETibW+CoBLTdYZ
GcdHtYDiSAq++bd4Eowx4UYDWNskKCHazachpctncpEJ/cMb1QApkvC7Dlkl1Nqy
gGgaLBsWT8LxtCi+8PteJIjjyKSBXzi0XNB60AYaw8eDSisjAabXmgJWsbKyvm4j
8yJkXp4EjTH0UrOhMFPQKR1jBNyP2RIVZfe2qLeZdPaUB2FIr2Wmr8jeALbljrpW
zBl199Gp6TWICzepRpHhIF+whfeGw9RAqS0MQJJ2AKTkWFFBZFtqVENX/hQIaGhx
xDI9oF16Ke4el2uxfK3DoOEe4wTlCZYYPH9/gG+p7mskqMo9zfox4KTTiCjbLoaE
MtbAdXRRLeWVVrQYKu3X2Mx5rL85lNvhQxYjtHdKWXZqLydfWxgLInkBvot9lr0t
jYnTldjOKVU3Zm+WVlnL2tYGIS0xgLlwzD67Gh+smYpZaAu7GdKmXlnIvecGVRbS
8jgAizqZ7xS3oce05GRdVPmrh0skSSDQtUO33OI7qM5nmNnRyaqIEXAaT+ww2Wgk
ly7EXu/ttjIxDwqyiAa4fRyBlWRfnE5ZxOVdlH3ituC71JAyn53Dqe5TUywpA7zX
7zRkuWhof15U9J6YTCxrUEIT/3/g5FmRr0nUz9Ayv7tspTwERhgMxiXhW8ioSGO1
ENTzbMjA7sNNKXnhnGI0A4A0etwHTG0/vBQsW2Fy4OR7GV8cAd6BOcIttBdMdfXk
Tk/89lhfJEQ8VLVDHymfs8dcvV/tjQPtreWxa99Um6rf4T1Tq0RHRGl95bdRYQio
EoClQOd0cbUAuR/dLqGThSCeHXDZ5l3yE2NLo/W8fJJwq+6obqtd5WVSda6NK/6u
+LgvbaP6nDNplrew5BMyvS42XmxySCtI/iheI+7BYJVZWZlGXQdpVozeZy+rj7jg
LmPxH07dqCAmQp6VQjDh6NJ6uL5snzt3QHznuQDOnB75Vu2pAtscR81qPSNqlFdU
fnFURylbTFrSjjeRQpg929O+yFBmrmbeQGO6fhtOAA7ZEhBT5T6DVJU7Vpemzctj
skxvJakHWKohl228pKJOQ2lH4k4hye2dVrlrLTatizbaqaomdugObzJbB0kDtAXM
/obgLUXbHTamUqs7w9XJI8hL0DGjaPurpCuViJtw0ejvAy2AD9Nt29uHWu2jG23t
qAs8+/DlRrnBGwjkRBj5KxxqHZa+qLZaB28zZ8hP+7fxlAGb2oUdEDizPodJPssB
A9nlz73E+tm3dSdRePLFwCgDetOZvITxEzMoJCC2MqqPoWPh6a/gOeYPEhsLshYt
xN+kO3MPFnbBwi440ATBJCA389wphleshN8Vl3Mj6Kv7R2aPdKvEZ0YlaZQCqiKd
qm3Vw36NnmkT1TfSZe+kZGjeUylAEIuGyL2Z3Qk1gu3GKWjdvOBDQjbrbwXNTnzZ
2z+W/eWWaiextmYImFI9A56usTfpCVUo9t8iXEcc7u4R4YnGtbvgNhoLCLPUsc99
zibfRTiqXAxuPETbz5dtsq7nPhrUISM1hvbhX07bG1UJ0M0ft6NCi+7znxC2ctxY
+bykxmjdkPFLHn/dADb66dWlFK4rVIllaDsTfeMYC7Fu7+tkzkhXxO7nMGAR4iZM
znukyccH50u3s5IJlSOLZfEqMI+THvsLfiVSk7nBiJtFh2TCIsJBzBe/Gw8XgFRp
/cijBi2hwpiG0hngGQucZ3MzMG54VjGQTwxjoETbEFiqDRidHCIPzNQa4FNzFv5c
69GM57RVQay89U4l7FfE+AnGYDL7q58y0GchOAnWn/lXhgjY2005ZtfLcJN779Be
3sSY2a3Klx9j6CLu9pDkgCo4nXxMZZxwtdHPab3Veg8RmXQnIrb+ozrYDR1B5XYX
uxGSMe1vnceVmz5e9qESSfKAn7WPFavmYsxkeW9N1ivAWgygo14yXxJr+MDapWUZ
mv0ZufOlxzDHX5ZHmCFztD3mfGelNqRQIr0o1AGh9t0Oq2ME4g5IrZodNHgEzFrV
B5MsXafhj+lsiWytTB6SNEtbOkYrrzBdcF9KQFQbIgP5AJuhgZcEZ5ULe78/LRXD
eOciOjp+WBipv/HDnwhcY1ThbnOOASc+Kjp9bWPc1jEKduHRXOlDvrxmv/kFFf8B
keokim+gxmx8zUbRCzGtvCTCvVS0DJnLlSbMzLLkkLrAQcGfULLV/sUr1n4tPVad
oQ158baqNK4yGCGtR4negj40Jsju80CZj9kLo3OcmEiD6IaoHq+AAaF5lpS7hRQe
o/zNZtcBHsXZS9uiKwPkUMHQABKkqwfZxNtfi7W9lbqYfamt+NAkdw1t8qziHkWF
ppa1cSmmnI8PounZx9uBvURMEf1sdjTd6RECoRTx4OyCb+EH0RyaF13Swg0gIz78
4IWrNaRAC5BO4zbnmtmm0o2pnsC6fdb1AKbzUGBZVLPDnDU74S85Eld5XIBs/ey+
iFDNVQuPHw+Bh6yOEQ0C0xzStM0gndgwClDqLOyY/mjfhP2D5Q5NJr86Zu7Jxubr
97kvQJgEefbKq6CYdx3g+jzSBxmHUOj+L6KRcnntvlyCJWVD/MzbdSufTmlgGzQx
GZFtZAOzCmyKJGGR+jnRGhI6Vs/cSVYaX52+UwH4yIBg9OxfLjQ6VD76BBpVO0fD
B215SPjotjs0dn8eYCQSVFVLO73cDEVgEnD1UzjBi9gkk09Rbs39j1qds43lyCVl
nM4u4MXiEZ/dcnbUsGdi8AIApZ3eQH5+ThYhyc90ERnNaP3tzbAKyz3MpcJOlucr
XCk7O4NQgtsR8ltslRFv5hmn2ZkfWPEhePzj4lB7X/We45URX+gkv+ESWPU+JWRf
Fcb8/Do1StrVyjqHeWshEatBmCYUYrj5ibK+8eA10d5Tz7rWJus4I3I8hbP4cCxe
QD8eHe4iN2abC9fooe1nWCc4I4SWkq7kS0XX5LBFGnGk+GBlwndxk92MccYFOlm8
GWw35nt3rk+LtCSB0Yve1/uFT8iUVHQrS/iKBu5giBd1732vs3pQggRT82gQawxG
f6Cb69hgmesyBs7BB8xlokOoeXKSVAAUWiRiZMsMtNB6W0eO81G5gwgk4x8g4S2V
t/ZMc8ZLaR4/STMMpos7oZ4bMiDtAVrw48iKDMzutVkevHV8mjU2H2Q3+Q/KW2vO
nSLCWJP41q0dRPaTJp1DJjLitiI0sVGUV8TJw7zNIP+j3IENYJ07xUiml99Ugt9+
08bjH8FBfDckD0+H5oU6DFRzcvNmN3Ty7Y++qw6MlkwuG2JLi0gcXnH90t3J6B1Z
mJV/rNupYV/fR4ORAkA5JzN3MFRTjErWhd+v57GNXHR0bqvNIAtAGz05k52br4bZ
GhstDBRHr6rDVJrP29EF+d3k7fUMdslB0x6ajO6v6CuRfTywO3MlUBVwM3lzwDp5
EhtYwnZCm/FL1CcK3tkct4UbPu8sRSVIgSj85t5Zn31PYJ1ao+idTxXw/OROy7P0
QWIpXyoVaSLxfGD4yH+gec3AGcSvI8Kd5n9ZonRVHkkDF3vDe8JBrE+EKi/D2vSh
KI+Y+Ts1PglqNQ2lWQJWeOgFmvFzalaDMafPJhYP0cXBPVs7JeBmjZg7ZQLRO6I0
eJuKaIJ7a/ffr0KbD2rolzE9Hxy/wvHYHHCRbWl9e6FkaFDbFD5AmiQ0F93mA7GV
2LR2QkR1NCeoEw+5QHDvQY7YRMD39MLCXBZWel8Ojoa9tFRATv7eVg3DwQbBfbd1
siMOj4r68JMF2y6Piv8IORqa8dA117lEexwpCeCkLDFcCMnc3P+JowXZHBhcgZ1j
3NQPZqfMTE+IGgtLBrTzdOjM/zjMqhhgCJHsloX5KnYW55n3+eicWUYO8nHW15mN
qRa5R6YRuEpYBNO+7jjPW/HlnA3qM09Stx+5kmhh/W9Bf1+MS9x3n17tQfnsUfPS
0Wp4P67nBRryEnN5K3SUTchCVWNE9jxcaL6YafHRBglYnbg1UytG7uYH6dxOu6fm
KRPR7nwwt7J5p7/PnmqTtazUM8yL+PnQajOmY4zxIf9H0WEMicLyS4OerY1qFntV
niwYOu+U4NB1WaiNqWwyY1E75Fh4KOQNs1O6n6uytdx2HdBHBv6gxkGg/7YSDH1R
xPSzv5YoD7LLStBH1WSossQip/zvuoHnDlA21dlAgHMthgvstpPy9Bli1lhZf5AK
rvKMvdbAfD0IlShsHPqasukCRBPPoDLcfKofrPJDxNExO1TAShUYVVxrBjMlWz/O
6L5tR1cpp+JW9hqofyx7bxOPyaNwomBBha+pynQ3ESaVbJeZ17+BFalM3LpRTLow
Wy2ceB9xMMMZbQLD5sByO1dyH4iAbLJaVavA/+XnGnMge1hzxb7+P9hyB1WguGlj
alImd5SJq69EqzV3BxdC8e0OH7BqMj3Sm8DnxLNH7h+ufeigmq2g4HpAeJHmOHOU
W3hwp/3rHP1cyB8aaR45Wrldixc8lwnaR/Z2s/l6pKztKx2/qVwEHpy5QrVnOhia
ypZxDOPnKru7j+EuLy6RqNfJtdoYqbt9XOu+PtDti7tD5VM9bN6aapaJZpqGRbOX
vz0UbMrcOFp6/pMFT/gVDt5JpSCcETeMksa/+qF6w9ubk4BO4qFSDDX7wa+36rmo
PE7H4ozckZUJOMCXkg+vNjE5gBk3FGmGTWeH5lW4VT0CJ2i10LmQNvt5lXFPpuhA
n/BWvyOY+CqlpMIFGexzHNj0r8Z+t3PiuTcZmIOM8lN/FqYS/Hrf0BTzEg+9dCqf
JjnGoHWaQm8jtXxNZzEqCyWAlWUJa5zc2nwtvz9vj57e0EAXw8ERFXkUpHG5Tdeh
Ex9JXNDRAgL/S/v0FoCKiZEmK1EI/rga1e2kYNLtKImPkmsRhaNhSHaN14LrQpDK
TMaFmaorF/uftmc6dBxXnyWUewH3/IvI7JYe1rhh362i7Z+eJwivF6RuThZlL4RZ
cxSi8xa5APA/IJnXc0EnoglBjUNmSYEpSeHwyUXjXzzt+X2V/YHAZYhtKzdANmQv
dQpo0KzcMlVQGt5kyTfnKnRIxlFKwySbzQMvhEEsXv84WQtWHkALVzLou3kzF2U2
VeEtoAbf5fxfMcpoeCig1ZbKGtzdkifPyK5op9cs/vt0D1NBLOTI4nYp1DvNG6kv
eXzve4mMO7eLiBWY+de/7e8X4HunoAixIhyq/XFkJqDAMg26od7oPpQXuFFPz6OS
Cm5PK0ijzuLflN5rMEJPYXnCCmZxZjtrv8AGCCGhGW5YT/kMK/rC5hGXhy0MC9RN
vw3MlWZOHrBeVQfKcuEYS5qZv2dFpuNHaBuc/ljs5Z8sz0HuDkANxbPfL1CIHGmc
m/mA3CqXw1pePSW+8Nz/UoO7hv1ort7XKj8rQDUvq5WbO5k8vZYgmIJW6vqpMkdl
Z0Rqzxq4JV6MnMtclGwiWW6t+/GHy/Vj7qYsmtGOADHK/rutJbYWZm09SqMWqxWN
dEqQjUYSSJUT723A4PmSNwwK5cIOtXvJWgOkYzdR3/+ffzvoPFUvlFqsJFUkxfH5
uNsiCVWpIP7SkrBSuIDFPcJBUiOWnKoyfnLXBuJsHDU7vWqVqlqI7NqHNkmZu8k7
XdKgLXPy2Gvcq1yejjwBe7qgoWml050YTuw0ZWqG4R2mQvYtEwcRwQKI8TPo+sPN
gQ3/goLXuZkTRbg36Udk6p4YR6TK/H7CS+3t9tqdFbO3M0Ljhmk7xNAgOhIWK9LG
VGqiLxTCV1TkHg0+YeKqiZTjEVmSWTjcLtl1zrz0w6YSeD9lsdLAafwgMKiTqVyf
EuEbUy8wOI1fPOmeclDl5InJJRn9Wwg0e9DNmqUCe1t8xDP+WefervVxK5kETBz6
0BxFNFZyg8eoG4B1jc8CMVx437s+9Cf+6YZ71bGCxJ49AC8ax3CxF6oLEI/hXRFy
aZzYPgvqZoNTIp/8H5erjinLo431xzrBcmt52l8zp/KswyqeMNnNQS3vtQ0Vkak9
yeeDCGqJNICpzw62knswMDeFdmnCqzcTRl3lLL/SqXkQs6l3qbYoGXL2XGyQI4HC
hqFENfhKOVJVm77tonlyncwjftUKe0juKlyb5ql1fPLMEoBFKpHltBZC5nkkm5be
x6clb1QRpwnQm+OplaT/FjJcoa2liprowCvXgyPMTwtNUMIBH2VQdiMstVGTmA/X
6CmVQWHfLk6QqTXwNlRYd4Shw1nZDeErXSfw3dZTIqWT5jfOyAKO9E4PxjVoxXlQ
Niv1NfJYtYwtU0IF/6ZOPFefRwHMEylkwgoI6tBsoLt2wI3IIk/y6URQKe+q+3Lb
M7dNp7YB+4DaLW9aCyZInqtkPHIEORVb+ydHtZXwhbk2UUJlmlHZjkwwwoEsu6rX
clLHjSyxN5CD695afvztWkxpNAJyw2kp61n3BOb9dRmCriE45G/lcuUSkKOhq0o0
oNrE0XbSrbmcf0WefAITmnGrfS/+7CA/F6BUH6A9gKSvU06pW+559QAf7ue8hBf/
5E5tnkiLdAns5hVX0QJD82jofRNKuwNSn+nSXL01lTWTV3mja/IU2stZ3mPgWt/v
L+Rs8D+biABn701O5ZhDCtWxrGm708AyIafVBl955IoSld9YJlNgP9ZAG0pvHzEc
xxCsmW2CSWxBFitov1swL0JdyP+6k+ucGZHergl5kJjTn2IMBzQjU5TdnoyDnmYt
jJb+AzWV6GXtlChfe9qPm15NJnn5JNb2MJ9lM3oVPYRT4nvYchj9jcVnpeBlHeIY
CRTY2keh7DucmQoxH2m9FQvcJRfBIAoKXxoWFcCJLNbGLY3ByHP48EH1Ba7FR/d3
yUHDt/jfapS7Otd/O9uijV0JjWvDruUoJUdmIlJ1tZK0zQ15RTvfyXs/Y6DeMy++
3whPFf0UhPYYAGicg+CYDrQT6MTRnngIU3U9jtMi2fy/I3g0v+kdem0QUJy6cnQI
SA0UWo1f9kLKJP9oTTtOazM8Jpz3sdSVoNXKgVE9W6X3+h83nJnsFlfTavhnECTy
vztDcP66bwYvorU8834vcWi3v6+bxWK4bg0qfdVF1CbEjvD3OlBL+rF/WMzZOFXg
h3zNlwuZzZ7DMIb5404Vn8/gv1Zqdrghht4aVUvqr0huIvGJxFEbxVNnD/j177Rd
vt3IPhZobzioa6rRUV+597Bvv4sOO7s2QfcSVhhUA7h+AV86JB1ia7G22uh14At+
7P1eZ+mpvlMhSG7cLzwZfXIq8XQiWhYD2icg5+2mrrPxZHo+AYwsH9wKCDGFu3Ck
CIiUV8T+Yj89cLUVXf+R3mjhojlf9Az6hgzb00eat70I+O9gUkTnAOaZl7zW3gRr
4AvcvDxbqflGwl3h/O6PkzWiGwU9c2zSabP7WWHlIGtDtlMW76S0UZ2qBztQ7M5i
ehQe75tAHXcW8I903TkPevBhzXp0TqX1kVuvhvT8A+8tsENrmAZpL3olDkXl2rA6
xDcDL18Z7i4Qt2iccO879QJ/AwnYTgD+ZgpUBUnVZXKVRbHjguShCP7JevA6z6tm
8wRQODt+PWThHSUpcYZskqwEJnNyxfIqr3XbyYB62x32rvM4fFplisxPz+/Afw14
qbMDEMSvw4LPsKYrhiV270E8rFRPJcozZgJYtsmVnM7XWNsZlhek85kXYuCFfrq5
+TRnoh4bvrYBEhqrAAsCKSPyHuXtFx1D4VnuY9W+NwL0yrgpLFGLs2/kYpNu9Qyh
gjudcWLIY5p3XLLLbFN4H5dgvX9LM8BoBF6QoqWOHCt0FcYZT71I3o+qVC2J3iRz
xncczLlBkwbaw8LNtSBbAf0RwPxjRJOy3zglLfv4eFuFHoBrXyEHSi5QuDcOA6Uh
OwlPG2u9VYk7nb8wnoABaFL1JvLnABV/ogceT/5P8ffZwpPKoWaZFLTxtfxi+L/k
aBTAbcyDkLJIs8ARiUN9cQPv7FS7vaJvwVhr/OXmUk3EbWPO16demU3n75P3kM4+
Krtp96H8XMqvzIwp7hF+0ocdcK/P4Mj0deUOj0csorDkT7DwWh+d0k9XA3TdjHq3
o+JSBc9IrQSZJY5TG1qyjVFpsAqlrY9/szuE4BMgki/oeebbOVXNXAHuRm3JxOnl
ooEVdg9DoWHtXWsP1ZsCs/nGBP8vKlICv6ExqpFYgfLYpZXnUZNsDvxfYZ37/KfK
Y3kSi39sKWzFx4YpQGqQ/3SHIlxz0/tPRpAUATXGqa4lVUr0R7hY4C2UTeCIAzgA
3j7a/ax8gspA3YSst1zRsCPU2+2m+SNkFl34sD0CSIyad1raIbtwBggwR0xemw+l
1y+oBB8IDHoH8+99na+pq7MZuaFH1qrP+S7KdKK+h+2S6qDx5HWETYeBgNrJMjDq
XIF5lHusPI8wmx9Q3PeZ9Tx0CG0WWfWFkp7OPH+Uawn2+rbHobYVXX85gYCzXOkz
KojSllNWCG2CKnotnWz3U0VKqD3Khmai3XXUHXNen6t8YKvDg/Tb8u6Ere8TtbXw
z1RNTIMpSLZgwdyDoJWbiJtgRhM73KhC+tRr5AAm3adxuOZLZCmQrR2ki1yZiZec
pGXRWNkWbNh0XvLo4eRZPBDWPif2lI99TXfQore+4eiJNoBKx7U/6YvS6Q9OmVfe
6hzkkr0nWk2/qhaGfrJ7bPNRvuJHuSzNq9ZjpHOZK08fxioq+mhvNGuCCn5OCmob
UlEMNbHVDqeu6rtAdzPijlxwZygHaEKoX/B78tgujdEL7xnrYOVkaIS8zW3OQfNs
dHCJTJCBPVWQps6+3tSl0d0BGnmgiD1i03vfDb+r/HvYLZdf0rDn2XzZx4R7ta8x
/9v39LmD4hu4I/Y915M/h9Dpa4acOWmwlAgyLjQBfJokMvRFAUZkITgUWQb04z1v
RI1SfSBk9w9mCNIe/R0QhgUtYs88KsG2YKkAoSEa0WwoGowePD+bus5Oef4jODUQ
+McQRH9Ocb5RVkjtBWERjzm6X89iXTyDIBzvBTztaf+FXJFdXeTD7Cs62IOXDErv
uy/bQSGgbnByTqM81sQ8yJWU/SBtfOg0EaP8/M4tk3czqCiUAp9V+vjk/3d+KfLR
SW/F774pKFLRqSqjeYgwVnnzSS2VVbKNTR8SDEyv2ac3fLU5reGSdHDQZQqb1iNJ
JIbj7d3PE9Jd1seGeYBBQ5DeC/1HksvdVeMxQWU4PWkyTn2Zo0YqHqGZZ8B5wE63
f2IwIUs9netFeUFU8q5pYcKzNSppqHvauGrFLyvFZNpDjNt/ug0B6ocHJqt73owP
kUQ/N+u+2yqOsYqgK/7YDyvGH88CAu70aIwPErC2BlGyEPa38e+QbKW4GR9ZFvin
WLGK/AyYh+bnxD4wfhafSXMOyhQZXmiZbgI5yrCfozp6K4Z9bhi+WP3QoKwpY1s6
xwba1aH8m7yb5AaaVhcqINP9Fx4klvGXH3W9IQA7SxfpBKxQE+QGxSrO1kGNQK41
QnmPws6uVaR2cy3vnPDllQzZKrnOufDrwmwYmdNjOh7eyLyZFVoGNfDRgrv6KUBT
QeolOVEPRcPdTSSAQ/Q6PfKyQqWDiU58Dgf4WIyqtCmGFzxJxbNMZV3zg77SBQe9
FHDIp3fGwUBjvF80rVrjGEk6Zrtw86ZBknIxqBztQLcdqaXPH9CJB6MLYvgvmlMR
5H1UD2dmrHPkmVwDxgmI8SkDCV7sTp2dL0lEcqgozeN7txnZJzjCwnfIrGYb+Qmn
AmGGOZgGBkEpkHeDUJvPZGbVxGvDlje5q2AFGACGdyh9j84DmrkW77nVeT/HIWCT
iFMYAmz41rJPr4rEGvHk0+orNnlsLYF7BJST8EhvInNWeYMxqMoFQkt71gki9vu/
y/6DFocOZ4UGIJ6jjjcPx1+w3Z87QqBIIP6kVKviJNpwPwTKL/Dl/pdwprMRsaRC
N8jwfcHEkdBWGSpagOZ5L2MWDcMmMZ4mKCpTKWYWBx8Kf9S2rnS56YtcpNVdl6w/
x+R406Nrx+Yu/1mnRFDt+cGD+Id3Rtt65GPDg/OIxuWa3QVq9H7bcBOABuWDG93l
7X1WUTkbig1O7pqMcG+RPH38rrEpWpTzNjRBLjlliN+3lKqcgmKAHMCHebaItQ2/
HxuOi2UTZwlC8uEpu+g0s+u/SZsSwkDyR67lYhu15LTQYdzwAqFjN0MMHdON+qNy
wELLnsa6n7NTq6ypp1qsKYG8ugPgvZXTs5yGOsdBjVO/kdC24KePXoB+Y5+V9VEI
nkY8pvojwWUxPmAO7UJZjmAqdC0reOn9ZMahN10XrL+SAILVpRZBv3JxbLFV54yK
swqROZIs363fLPdYBWWo6Jw783qj3Pkc4x4Mz03Jof0mDL2wIAiOq/Ke+8eiv5w0
Ki74awG4Cw/1P8nDwfzv3bAW6w5iKVu7TJ6CCzu3jow18nzz50vl5jbJ9W10AFdE
jB7Xae3yCa/sqpmV8fqHxn/4yIFH20Mh+KTjW/OviL8QTMSoSH8a+eCK4o6T4q14
JKQobEds3i2yavoXFpl2WCec5mzkzYZNjsoiK0Dl8Jcuvwz8F8ghQ1QbiyFU91LJ
bNxPGPx38iN3sLQpfmQ17xdl4nmAxkUnT6kMdqQd+URniksQOqGlUaDK5vPv4h8m
bRxS1LE/Zspc1ozx5ovAPE91Vmzue1lzuM+Iba9dL9rrL3eWOl87Bq5b2F0HmRu8
NuxbLowA/Zr+I9PmtDW7J6DABVPUJv0fsvCRChnq9+uwy8311yNj7Jjq3KsHmxN9
wLBtOV8gFHj58aOTd2PtO010sLolZsNwZC5xb+7LfR5RNQSMW/DLJYEntduY3gJR
C6u3NitdOXaQ2qlhEU0nFEGhwMeU0zoOsZf+vnzHrpVPi0Fqka4ipFl6//NuneIH
fUOh09NGzNZqw7X3D7sGOq3HXmJYbrhcwRK+sIJ1hC9qgvwJWkA32lYkdCbRp1oi
QS4IczM7K4hS9Ypt03yhiPtHZ1C1zUEn6WaqjjzHYFoeCd3/KydhW/4cWKsIl1+t
7hxaZQh991GfkgVcAc14DFeVc31ctEZDZtniVhyZVUnwAX8cEi4jSV1sFBoOLdx6
HnK0tQpI61PI6sY+6au51SaFTISrm6zxdCy6hHymA/QaTHXI8psfPzmP1i4lBcrV
zp9i1UIq/XctrPIfZqo+RxFKvbhOAuORugfXpMAeNhntQQ0mTbSqCySbhUb+b9g2
6z6qB/v2uK0fRwaea6lV5YAcRUP+823Hz0/GByi3J9ovJDqDSuUBh+z2OweWquRj
EA8ym1cKrb2RKdOQ7jOXWqFweGPeizrxf6AcDWkQmpVt8aJIUvwaxQguoBnlCWMX
6DeqRlp9gdh29KiK8M3+Poc0If3klSuzEZBBZJYGvE0ezHHW7tFok1yyRexySXrt
nVZyFmGhJwt9VGho4W5FF4Co/xfQNImxRkKHccQolBD2xVUk4fWbUHJRQJRLtz94
1xJWO/Mj6qjcECnUOXRympCtS28YA2a+ZJYXqYLwxaAU255f/PPb45fO+TS/vBHN
Xm8WOkxq/2w9sVWQbudBQF3EtaZF3ZG6znK4L/D9oozSJdKgoglDxJSjR2kP1/KS
dLv0VNBIOHSnmGevLIMdP4DGCblzJ72i+FqnIcw37YD+HdW0PI48vV/apWmbYo3K
h2kZrna6osqF4tx7/R/zajLgXGTiD+soIUS7Xq1RCWYcTERFlX7ag54cR021iwZw
o93JTY9+xf3wp8NU3jlefxqgAR9igmd+LgupyaQg5RLM4LP1LuId1XI8NNO46fT4
jI7znNSTqll+0L5QK5EgUnsNQkz71YEffGP6k+ryO/i4Y8dx/amtKhG6CSXk6VGh
SbMadQR+76nb7TXg3GhJonlBWGd4JWjlRcmVYcZl0GbZY8cy9wWbe+r/pDzsar9E
laPApOiBm2MUk/haKCfHuyalYmyDOuOZIDuisIQuWEpCzQ/IqTA2ieAvhuIgwB+r
uX9X0ZnOuFCDqhHptEUzhcgDlwxBTGUhJd4zhRqlBUVFUyJig1ZpPQl4rRFmm+sj
wbiR1SAkkDG13t/aGLcIO86woyBIwYUmlJpAu5Syo36IfTVV0OsTG13GqRWeTP1Z
QmX5qvGHt8od7+ffFGzh4AXm+04Vy21UQhYm+/jKarI/sc0MC195iSE43Rc89hGi
Pu7zWIYC+jZmZFAu5I3qt3hDBLQU0407q6J9WaaSfQTW3GJ9GxKLSZPNI8ElR+bf
LRn8n+0EWgexH2SXRDQ6nif3m18e16NVigtA50ilTCRQSMADV2aLGmeOGt8Xmbx2
l9Wa9koXt9l0IP3nsAHXIUDRbkeImcAj7Tg+JHFV343pIZsvj9kwd44LhJE9/NQo
24GPsYobCAhUlEwOTFMxUKH+gJLHn/XrcnfDuLcllSFchHgI3/BG/XCSZ/7YNr0F
kGRlp4jLrXH5tKWnziJJ9uoOs/vqecKnyNpYlbD6kmrGs5vO4xD5wptat0JleFr+
S7xSDs2Cvo2mF2BBj/x+U5sDW1x/dEgE0cs/JPu5BQ0f+dM9HiH4eEXSrUvfAiHV
wS6rMAcKqDPQX7KTLQ8Ys63WfO+zaCEgETMjM7vxUIFPWh5EpsWhZ/p3xs8LeFvw
G/KU6ej1TFTGXBfyO/UOs3a6srj8IhdqIcTnPMYhjnn39Vg4NZeecsrAR8OIjz9R
QUbKz6pMxhYv0jsccGX3AgU9o2cXpS4+GOrdK7lyEeixEec9c8xAK2/3O5GjEMMD
08ebpdCgABnr7iN5rIjIp4tMsUJZJ8Bsz7Fra387H2/w37bOl0mZ45dtLb5lt8q2
nzEKpUOt/gwg/KO2u3dihY9gl6ip2tPfg7rpt9eFsnAV/vxDP6Yskm3JYQoKvBa9
dWfZLzmrR9YKkuartFQuTLSDhc344cUTxdWdpmYBWxfhjJGJe1AmvQK4o35byClL
Toc3Rbb/vopOhW/izNb8KFaZ9/QLjT08kixdkfjsG7QvL6QQ3FbWEMCQ2SIcaPNd
9ZOUXZsocK5t0xJFbte5myBWIRXNntlZKrdxGw7ideJd6p+tvM6CL3AHsgrJyJGc
00s/kPv31mvbwrFpmrsv/jINiEDtar3NVguyqBWTW3SsKhBDGV9kiX36BByn61Lg
CALDU/ck+tkIQOOdCzEGuWnckcmUZlT+91m5GBZkiA7PDR0X5lAxYqrTE+qJmGDr
PraBZliEwcmXWd57tNWAJhEuWc/s2kFjQXnEYnAy35jUhqlbDdv/48hB2YlwM/y9
dDDd9x2bbuQ3/Bxs4IXWYkIz6RQUfxP47TiQ/LxrJND/Ct2PKPOdj8WFqAj1AJ2+
T7eeSFwswrhifeltDmZwMN5aK8nRGVDqxZTIBpBRWm1/az1SzND7oIrg9QkZChTw
dacTOV7CrX1Ik01weHR2w8Gb9bersXFDqBhbCaaRFvFOGApQHr71Gx3K8hRNfLGB
UT6//9350rMlxRs7tiP3VEMCJNpWCbvJDR7O3u7TCmc1gv8vkg0JWtCritQX1+LT
bfs3dlqCADXv9iTiwG2F8Sg1Twvn1ebczSJx8boIMwdUZ0bV004tUJxozFnmvsPo
sXcIhOBm4rG41tbpLkUE9AVc7oT66ZxNToMoXB3FoOTteD20O0JPrEOlw2mZybux
pmEzvN1kuY7R+IVs+bjvhZg/sL5iu4rWk+YIlaQYaZuSQLBWiJBWDihABJ47SvhZ
uln8IkP1nJY3r9/Y3Q4IVQOtoCguZ1F/fmqdrfLbqNiZNZtAw05LNb1rrwOBYkJ5
HnJHCRK3ebylRBEIyvwI/yhhXdNedFfadO/nf3VYDNx7ESDBQCznukfqwGg7RQNv
ZbFm+e4y8XUwy9LAdWvmys2OU2vB3WE83awrhghp3Sadv3/6rTt2HIpAIs1isyWg
TRg+LPIzCmuvYLDYbFJ/7aHvNyHarHBYTo2+IOxNZRitdlsCV3o9T/vdki8rrH8P
2Y4QJNzhZpFsHXkgtH8wOHlSv2LnifEp81Z6Xclzf7Sx2ftq40Iw6CnMvvbUwcKU
tAfUmDH16MvxC3T8Esid+uW9pidqREO9wTHb9UK0XBeZRR3ewt6lAsBIEHvbfKph
+rsJUeEH9SJysnSTG8fNRcCL/uVRO6mRV2sR4i8eYGd/eHyzIrtL8zcLipssw9XF
VaPohA4pvBlLDAnaaMdNWA3/ZnPGjt7GzZilPATr+e1TLIaDu9c7s5M5ABOzll1X
FEed9WklejPfRpJNxR+6dlQhNWQyewDKp86W06aHpIlhQeMPUV0uVXSE/goT4FAc
HLyEku5vIDjWbZwAlMUjyC0/Aws0wP0Qto0M8TGy3ZtJJEzycAC9+L1GJIGgyXlH
KNMPw616MXNxxMtuJYnePktRoxryxaNok+1F7Kdcw7rmUi13+6jhspppuSlwQPyM
KwowyLAgkdGU3uT64N7n2FdI9paE+2tHi7mpd0ix+kZpYbOyF+dm0rt6/WvHB/+w
Py+oqliHzsyBHXScvL8BWpL/cAoY+Vd9YSZbmySTfmOAfEKGSiOZCaNTNbVuV4QK
rWP3IBppXPgEJZxb0EQlpurEVlw7cjoPCLaZnu2A/aUi/GPNb1ZE9SKzNkS+eZSU
D2UWWgZ6xkDJls/ZHUPa1R2ITCGHUsqhMQggfIbQQn+YOKkTyeSskrHiZ7yQ7jYs
ExpnDzMcmASkpzE3kthqn+nhMNsaEUfV46BhW0fWkzorG5yazcCLW5+2t9ATH5or
ZsPZ8Z7X2WlhnBqGMLpaYo8VgKNJ2TCKS5W2kVOIBT6O0nB1zW/vXEMdxSBYdq+5
kvnQ+iAMdnGBZbhO0v05mQq9KYH0xYgTdQkuvis9BiST3i6pEPXFOrL1JT6jIuz5
oZ4eOgrgRwbN14tTpqXPVabybwgVPVeVxeYBl61rOAhHsewqImp769+G1KAqWqZA
TrifVayKrbortgyFqT1LewPWz8CFxbzM18OfmRFI9+cajFt/w/SNRL+cB57VZyXD
4bzAGtY8S8WA6gzl5ysrb/zX2JQazPkzT7riox3YrTJnjUHncMQ0W2jU81xzTV+W
4AGFjW6H9FRtHTt3fXiraTlPSV/TB61FVZV+WQtyVKgCKYi3BoTET0nuRlaN+lIG
Wvxyak5gcTGq9X6hdwnTk9A0xLJG/LEmSKPwvMIQdiBbc2w1qRo+B8t67iNljG4n
rpNxe9RG4fZXoa2RetV8hOoI1kzhB+twBzonmwxtLyHFgzvNcMvVSOAfr9pOBnZC
/C+xa7aIsM5K0gznBDlRSGFbkv8GeY4w02ePDnoG1a85ZEMI2hexj2QWtkKwwwZ7
5BROdOqDsuTDx0sOg+UbaT++pbqaRti1OrdMMk5q6ysq4UiKAEryP3okstVMJ++b
jg265vtDPEfuraIqi1SkoPHP5/K4UQbWc7GuO4+mNLUkofQ1uDa6UsGYmt641k+c
+lB9k8A9fpqK8+qHz1qLuSQpCzl/Rr9M+Ix0p23pLsx7GOvN84QAJHihsKjiXhhb
9xs6pp+HW8U3xO/QEY7SX+iiEgyFkt1+zCGePnUftGmUQU/CLP0gc6peWMaLVT5h
AJwOA7lsHqkLO+9yl7RdctCgFUU0VWB39AZVTpd3z94+MCYS7IHE0D5hE1DFVAWu
idXCLGp+rIlg6ypI8aYIi8cNvbmq2ffZao9BNtNHLINP2UyjO66pNlqDynS2usov
IZQZ8a0W7xMHyyS94tY9GtEv5+7Umt8BWyhKBuoO9o30JmZ0ik39VDdAuPnMJTHM
k6V+eWWUa98vuRUkjVIzbvuvR5EFA8n0pr1x4Dm9WNWTUkQQjTmohr9m62GZVfeL
8TTSQhHuB+1AhaiwO3Ox4nP1UyjnmgbGH3qf0Iu/0x8rrGUdkcVG0BuJDMqUnInV
fyMg1xhB8yCRL91ot2PjHDx64nowdnTzMghN+qWPd4LdwOCmmPzBS3c8MXJFAqNm
3d5Vpfl92RBEg5qu/jkqV2bvTFwT0soo5uByD6dfyWaM7TR9n3eVK0tTZ8iqVUMF
N7uigJ6S7eZoQaQ3j8h47EZfulcn8KGyIv/dv5KBGU3KQHxreIvIvPMjRs7258/x
TTlOLD/WBveKJNIm+0obQKQC2bCHBJLibL8nde3DD/oUrDTxOy/wsFKIcdfr4N69
ry1tx8ze+zMhk5/rXldLSb1uF1L6VqTYrAna8zYuJIMa7TtLz0ofzWb4Mxyss1mN
EYgV8oe5e2JGgNvNJUIldgSLtpTyZQJzVZIhm1EpbhPJRsEJOhfgc6T4O5T7AL7h
xN6ibmujcwFIXJ5un2GBB6gO9xXTnsoJOlrDeQ+UhDK59vi+u43EYZllH0e1MBrY
LHdw3lXH+qrRtVpzF0Ll/WPCfSRVJCabbIFWQuHPg33SbVmWTjUmhQD/XHnttYAY
3gaRgWPgMw21abRigaCc8AgQQjFZ3UTc1+XRFYWYcyL5xY1JH+lXfgc5b1PkuILO
0DRcl1FpspOa98dc8LaChCdbZXwNCqEvEPGXoXU5KPuLiiYpgHYeifncaKJvDbCR
ovUX2u98khowMAalCabn9mlsCk0//CRWqJ99zAnssFzvf4jgjFj4PR7TDD8X9DU2
I5ABxKb3f7vDyZVQ4Np8ikjsK682+j5AHqc69vOmXikv0WbYEyT8zmgVkQ/zPbpa
pfjeqAFm2q/RlUqUE++2FgPXe/Q+xbcMzj8LtIffcn/+xvfrRW8C07lDPXx8RLLi
Uo7zw+dGP71QM8+jAbGOSEVI70dlkKXDAnTsblrPirz3Kbv7Tas3ukLnR/zaSY1R
bktPQocWK+dnFRScHjSvVD6UKc1AhTh65mY+vH/t9aleE89SrR9qfeVVQEK5y2ws
K/SJL34kwHb2C+/ibmWdAwkZ667JUbl36UExv/u4hEBuXsfPhvOX3zfnr7Yp8m64
CGDTSOPk1tGlGdXc7cnwTX5b3qLqFJziAy9hZN391GJZgA7A/o5REAI/fc2tHV3O
jtc7D/9UlW9aqCg/XI8Chiblq/LtE6OnW4vG76VfOovPjPbQp9Clu2Oyi4xyGScJ
hrvj+35Ghh9fNtmH5dZF8DksCLDjVGTbaLf4RWwr6YscYUqd0+9rO8biSPMIF6te
3EjHJK42NbjKcJigdi7EkzKQii5K7GeXIkkOm79rbpgLV1fjrTcrdj8O5qI9Arrt
oKkiUxYTTHZmQqPRwr/mw9AGn0uCUBAK4O0VZb6Hot4eT6zrTs/wds57nqNH/D7u
St5vvLHIKJlWwcl01x42sbw4oTaUhA8JsQTORhdW3AAmwMgXRbGXPv0SuLYRqWlU
gcv19OJbyTY+mtI4oy/v5Rpqms8//0i8T+6sC0z1tY9aRzec5z55ZpKKebv295C6
U+Z0boGXMz7U4WtLoJeBAqEs0g4g77tQ5GMtq1iumJX7c49wuX0O1UFnKmqOfeoa
9yv1TacfllMLR0S/WKBaTGawWqYaekJZCg6xZ88a4CW3/s9gbrIQJ44MiugKMTH7
nPaITs5T9nzB5ZyuzTpWLSS4EWDbzixbErC9tAJw8yxmLQKbn4XhVKtiF/eG5qw8
Fj3IBYxkjmH+26pmtJRX0f0q6p5uenDU34OlTUfZmuzXV25h4DAJ00sq0MNfOAVR
ukJAINW0Gb+5efwgGBFdlH1coVzDZE47PgSbX/kswdBkjw184WHVhB+M9/h54UnJ
fE2vL1aKXSVxKiVFc/SxsX5cPJZXSziEXOLD7CBgw8gzlvyeqbbpbtyp8ZyZJ7AB
ObInkqpAcv02hVt0RgvvM7lkQvpvXwVx06bJzcfEoeA6zDdeep7hfsftJt+kKEUg
r0Lrca/83ww6T+XIZhdhvVhJnzxazbIy+jPd9Uzkwa/YxaqzJKpD3WZlShRRKGBD
hb7+0AZ/R1yWo4H9uwmgDRR/68GX/wFhqg1RyxCOwwy4nufqlcsEmfTeBcNMadUB
PJNRNIdV1xRvQZ6AjMQe+4mzAokATkoQjYfx6sD2NaK+CfLodDvou9V344Y3uPOe
A4hDorqxT17pjpNr/HacUuoge63awuTWE4j28dz+3LKMJzFnVHxPk35ji1dq1kOn
p+PkgGjCm1Cs0YTs+DSAslObI4RXT03kYQFGhE1dbgi0UszHbRcWUCUsv/+5KcFY
XG+18whbmqJv+Ly/vFZuArB4csLjvUKsSfl79jP9t8tHJPBM2U6ym06s8JccLESH
MwFfe0Q9UlOjKCe+ko0oxB1BohFxAJZVxOtp5PDXi9jWpb1j47aec0KKy85x+01h
5WVkF/oB2zWIITecdRCMXIBU10jowu+IuvNDZY5m8cwTv/c5GA4FohpZCjFX1Rtu
4TccKx1K2Np66INcIcUf77785RsdVYJorNbE/JtQNovVNwabII7A7zx/7IeV5UiB
quMUlasogHyWztt/pp7AyHRNEcw1yUpjdAh2uFtigB5ZQjQ9JiTztzCp1V2ntW+I
IoaPGSH64v86adB/X8rmiYBBsJicgV/zl8H0eCPLB65OaN2IIbUo79dzPXcns6m6
HSeKtf11CGppz140VC6uhJcYw1i4oOhV1Q7NL/UI7dIupDmgaj8YdW8nQKEaT7Hy
xiSC5cTBK4ZjfdnP0ZGCRqLYg0VwbhHe3eCbHdRXJxkHyUaKzvZQ6UlxcypYAGFV
wc+PsZRC7NYzcHXGSfBfMCMtKfYpKcqlYGuxZAqEpoNb5iRpJDBSPORrRRcMO/30
Gys5MamRu0xI4idZBYWDGuD14KJDcl53qRaSxnj4JcSifEJ2c8TIvY7/0B8MNPeG
W0Q8zb2tkdS+eNSR8odDeazpV48+nKZO2pYJiqy5Acoy36uox8s7iRiCjl0YX6Fb
poGQY/5LPIB8ghdB0/GJUbKhYL/oyt44WtJUBQNxmKftUtsyDCxz22Z7Rc7mLmD3
DVSK58anxWO7quQt2JSB/2PWcDioAj2RZgD14d+q6S0RRbsfmteEpPAiqUda8nkN
6KGyDq/22313QEWrA0VgHdpqShKoDdFph2hQOG0UTJmWnn9coRxXurPhwtbaoaZJ
hHyId4/jDUpwPuJdHvfwzm+w25IF5uLEZy6qvo6TZr13kl0O2O7GQ9Fmzixzdsf2
JLC7sluuo/7y7hd7pnESdrag9u1oBEYN6/aAqZe0h7TEvKpl5+U+8/BItmez7bVb
bYu8Hj0hD3SK4Gq8C2HA0zgl5E/coKWvBLRqhbw8SGqrCSwdYm7ReDpzERwc/uOd
CXqOe6Q2gGgC2YRHzvrhrZ2eyrtIKLRm1v4ijNbak/cE+wxQ4RBMcqIUYADVrWQP
C5mtW0Kv7MTqFMKbj6kKcD2dN8ydr2mowhhvvjddfmyMgtdHNkiEgWY/Ic8tY1ZD
16a3EMZ/ZAhgJVtIAbQQsuAuNZ21YU2mbR4ztCtWmbfe1UeGyh/8lrWLanc5H0fV
uk9GOElBv5sjEYNasnxe88Pctpk2fZJfbxiwjL6vOU1uBVlBALm2ELKTj/snzyku
9cD6lm0S8hJI6UIUVyw44SzC8nb/VvUZE6Ki4sXuG8FVrzQ1QHk8oohIHuW4Ty0u
AP8hQUFkJu3scfc6AhKy7CH8ew44JS+0PhPcNcyYbYSsN1Db0RHGlH2CtqHAFYGs
oiDCRQsxAtpPnSnTcHfdom211JyYrP2Oc9aTAEy5LkGk33JbVDL+PgNvyHJe23U1
+VKlGCdZ4CPqx/Qg/JI49nHFeaTjKh3SWnAM6PupoydE4Qt+Sq9O4evED/QpslAN
z42z1hic1zzDb6p1NENIXMIp0TZa9Ola3v/h4XM4vbxOEj3BfcpVSOdkEFWIRuLA
FGPeA56c4g3I8S5nPBSRKFoZBc/TtUn3IHEn+aedFC/oeIAtLzHghhGvWwA1i/jh
GjShjCl/a5/mp63rK/e6JrRkNSVj5s9auou2xR+XKfqwmKTqMBh6WRe73juoEGw1
m3Uf88/n8DQ64C7NxJ/JRxNoJPHTzbNCU9LFBc2xfKsV9wRrOuS+1Y9r7g1JvW9V
+gCyGe0WXg9z6mqs+cZAYtevB72Bf38M6J1JXdF8TJ5QvARSr5jUEAFaFGvtEEY2
9A4utCxftGhhgUQQKp28tUMtkluWghzKoPFcLs6wYNaZXNhPD7NVoDICL8axhmby
JuFp18Sp/Me+0ghp83wem/IoTub4+Rg58u7oi2gT7WwpYo4Hyu4c/RlWY+tUhfqL
S0rNqNjXECSJezlqPRpyxlgQWa0ruansaqKt8oGZZitH4Wutkf3C1b9AOqKqHs4C
eKC2V1c5Ar2pWUPxzMLvYHyZox7qp3n2nZDFpIEyx4wLbB3fKdMkGFLM6oPKplLf
gxxjYOa4mNq8LlqfAaxImtToezCIDDyz2fWf6goWdh39H/bd8E81b1bdvGb6OhVc
WKGP6+crlwjZV1/DV3lFmyjQNtBbrsiab2ql9tF7StNSB/Y9fzSSCgG54zbhYku+
Fd9qs+ad7FuO6cN/G3hLEYBgrLNv4kdChhine4sfcbgMONCUhaG00SQYtUSsUl/7
hSSrUPDJU71b73CuexetrceQAlPZwBGYJPUxbyrh1peSq2g0sUvh25JP3ZsUQDjO
ogrw89L3hOvtEslTQFoPTglX0+N1i2DX9mWiRCz3cckOYkesClGzuSmFGcDDPNS3
tD4JzS/wvYv1Vwc2MmmSO0p8dr2Ed3bJBdoCmNyl6wyk0//nZD35ghxf3rHf2XCd
JttWLBZUI64CXpKibV0ymBzlC3g1KD3+RosSRpGxP9y3+vogxAe+Z4QuUAp4G1qO
tUDtSCDpGD1KuLKKj7I/l+81mQ1Xnzh+nmRwKgXt8aDWw2QzpC+MQQY/YtArgVPB
43vKe0UdXFvY0Ri2nrkn+GFvCTVF512qbfaCSfafTJgInkbWvgvf2paoKsEpYjdZ
6jYdFlQhqdci9CT0oTBs0FV+b6bY9HJQnA5vvmEkXySDTqmTan2aGSfSlAA9jwSI
9Qt/wwPAOwFIcrNcL4ZpOVSzeps5rsSztkSxZE21F7JhpkRSI7/uOHZuqC5rQfqA
ex6TxyYaf2ckhResOzNMNqP+V/RJOu/MGi7CEUw9okZetgLYPUxHgxphuNtGdDbx
s/rG3ik/9a7kA/kdiR2TTyTf/kvqaxhYYmgqp12pmoN+bLp243tLLVD3/sbIRceq
hZ1GC1vEA0fU28dkFhE1p3gHAh+WIKzYsRQteU2anULVqyTaZZjjHK6ID8dYPVIw
cdswVp8wh8adr0qyf7kTXqOwQSNE1NuP4jKwHvLVlPvry/0EPsC431UYNm5T9uVI
ZUE+b05MtjMmb17fFuY7RdzUfboD58rWlEKUA8nipNnCNXCTgsKU+cJCBUJzOgiv
NOlT8XhUUE1qIVPagic0Ld7A/32HJUOibWVI0g9bgbcIcTCHvEX7yFU/HaqtYWUp
CtIpsSU/Le9ED0OgYKYJjoVOIbfpizAjOmV12QFpMDgGibMi7LDVdi2FDm3s7qNO
W0Q1wswBG2cfIAQP5loxMjwniBHTcDKiofcCxRuvFoGVHBWkrU07lXEOtuEhV0gi
0/NBqAqXXSfAG+SsmS4t0GgWqREtEYAetVeHz/3hAA/LyaQGmgk7w665zefAeQRy
jTxzIxMtuEcl1BbGefXzDmyVLCgtodaviTeucwL9UPLFTquWWqreVp0sJGMJraGW
BszLklLQloICyA0/20dxk0gMX3mUQy3PtTDoAHo/pZe5u6Uo3+dpjKlATp6Nkq/G
OE7p2tTpNqqG3TS11xg0qLY9c5ZFaAYXUzF0GvaerhZ7ttYd2Z15nD9NcOKwTwJ1
ZQjTqRyyTB6Y5EXu8m9OJrJRlzhPKWUy4BAN81Eshx0MjqaEKUV4P7diCPOdCWRO
pM2Q7KOOC4sM/38EhbwzUy6YZ+nJFKJysE0NHzbOtGI+IiEAo+fhBQHcADSUJ4tZ
lUYIm6d/2zmCPxICheEURh+yla1YeipVgJ2w48ofJbTpqqQv+7R2Y+LpIXhq8pfX
v8BOYiPpximS+zMOo7WeztovCGCFOWFbk2jiQLbbYmTyjqsKS4DYxlHtPGB+cg9e
PdFtaw5rmLRsqF6KfKglSvU7b4IhXjqnzm1tluMJyJowywWt6tqFaMH4lJoxWx/e
wg6nUWm5oa2VNmrKQUIr8IXtB58AxM68FM/tjKNMY9ORdhqywZzQeFI9y1hvEmV3
XAB7a+IUZNwrugHv1iChlZe2xsr5BKM1S2NqxLjkV09d6dBeiDMSmdyqIGcN03tr
eeC9BC9AUqg2fCLWE+u4QhPO6IBt95hmaBmm6YcM3VJj1mJtksEvvWnRg/TqBy1x
11A3VQv3mDGDXkQjaIlRIjOriuFqZGVlYjr1CJX5XYpCRbHxWPgpJnrB4WYiFv0F
Q25rwKCtkHqDZxGxwC38FV3+pWQEjZDUFLlNSp4V0KYsswRxgA1yarvaKdZ1+51Y
lLMQGcWPMUVCQNdt+wD2CZQ6LgX3PkC57CQW5xYgPfBxjKhhE395XcLaNnFbMRB/
71DlS6o4Us+8BYE4Q2z6acALyNRwj2AS1iiVUoRTA4gOqmgy5cdyQctS6H0EUpBs
LoWN5i4rbuh5W9ctu0Tj5zlEX+FDh4BBfFWmOA8iUEcOjE84JEnggxR7NQVbehFF
c7LR5yoaXDAbrC7EBrICf9uW8RSPa5cuDChO/eqYSt6585UGcDq7tqKhcNNCvtCx
5knCQNqb4nOMyTWkcidnclcQqKP0yTIhvWkmMgBUx8QszFf+YDg9iIRAT/E6dIV9
xwgFAprjvePJ8vrjuVCtkrAgI2QUqTFKCqGD+rNjgp81xP/lgdBFsiuZowfb8PEZ
YC81Vor4u2ThGZoVCUHSlUxNIitQtbqkg9Kt+CJ/O8BXIDovk/RtstntMrlXuDYp
QkAhFlL2qFd5UgHDuYA/j5kTeEwWHsncG7/xKmLitjRYEOfIZ5nfrb8kyzfdpavU
pcFL3IO4nieoM6n1kHrR2MWPHkmjMgFm8k729UBj1/HFgXLQpxEwJVEWTyMtBFa1
7Tv5ya2xyvOSjEKu8BO6eewl8p8w34I18heOzFwZqLIDiTzlyFkkJbQJvUIHKX+T
3Vj6DQKkKIU+WqFN5CmUN/aA+d7r2zukmYicjdOy7jTR6RVkf/qjOuItctKtNreL
cd1GQGRLyaoWGpQeEkc27cZmpZIlhW0mPsDx8PSe1fSVWqdzArNxoxQeTBucfHyY
hOi65N6RO3ZYilOI/SXfoSTiwT8M8/79/lxiMObGamM5lbmsBxS67z1ma+1SP+uB
WGxNRiuOYwbXyDTQM6LhP0vNFV5srklrSv3FFT+qNl9KHMdIvPzhiOmLPu3U8c5h
V0Bs91dvTeJZ8wi2tE81rATZJKD20Wbmw8taTsxErYGlrZXm42TzqSeZs8/ltfSt
7YXNnFp5CqYtkoyiobt+Og17ACJ6w4yBrMTW49b05m8cfexLNKWB/7AagFsh+g5U
vzN2OT5vuoaJ9QDUHPjUPbOnOPGxojOhgbAB55GWnDxVyYgv4FaQ2zpY09dU8htG
osDz6aKuTS9Reskg7d/ouZvSKwuaym7UHXnZ729JmmdP3JMMMdwiEJv/+xZ6yJTJ
OUfPHQkSpsADOzB5aPklaAp6IYh+MjAmg/oNp7iUttZaFa46/iZm2fcsuYNMWt99
Zy1JaShemWCyw7X6QgAv9rRHsgyPvEn6wQQbfRAm4NMbmnFhHax//msZQY7avNSP
9TQGABNOkTObn8SCUEKyPErUuW9JsGygJ4QX2GJe7hhXYmb9/vgid6Nh+eVeYT7z
XhbH+5s6qHIp5lNOz2ttvuNwusjneSPNIsGeJqhlms7+Y6TDniwZgBNkYVR7VzCE
2vUUBOQTslLD5xLnHws+frNcF/w/fsxcBsU+EOD9v1ldXln5j0xU5eDkbBAHIVAZ
IJL/bRIw8HhMn/PX1NLInJe9Pq9rCJtwNHNyrn+L538zUSZ/u6/eWYsXPNFNETME
6brkfydPQG75jNomewFoSL9IhpFNwJf7El3tnbyDwA6oGrqPROBwjonJ0+dmlF6O
IbnlWLr2ZGOj5sodvUDRw8u/OzZIYgSluAisDN/uAdX9mAKljgz4OBWGeXDhvTai
da6jr8iwzF7BtpVfzwI6nb2Fi1EnTF1/iyxBtF/fG1bZ5K68XH5RAx69RIARAGIa
WyRNa34cYky141/jgia5nA+Nb1RAweitqWcHxV5+6DESte39o9u+N6Gjncv+Heg8
JCylaHfPdJETEDytXqMJACnhgUS2WeQIHdH1I9jSYeGz3chGVx5cl5QkQIzLvnKI
5X+dT97dTLEXzUEC0VcKgEpGBQ+QePzuw49SKIJIxM6uebylZCMeKbCMlYIqhzWI
Xez5+rT14QnKP42TsShUBvAoF/oRPymmqTIpNOfsTZ+CHR4ZvbdlFgBYHP7xSVoH
KyBq7+0ghd/+2cfxKl9VpbcmGXKWi1mgQpUmlFYANQHftloKJzbLPE2mnNRo5JxP
hHd5dyFMzY/+tvwVBIeGO8K4hjd2sJoQkFzz02DWQ2aZXWiAUYo0ptjP3glfAfFl
030pf4TWou8+jdZIxyvyBjTMsVdMpl9MGjyrfnzDTtQTBo4spY9G5cYEjTyySweJ
4NcrlroD4/45dn9+UjRg/WAvq8+TaczDOKJFbIwUVxvu2jdjpYl7RmjZQ/recCF+
YbiCSKkEVq4Zuc8b2QONrRuD1Zc5FoEImC/u59GTc4NtvmMo9m6xeRl/FFLnUwrd
GsnMYAngVXeptKiv0wAh9ybtHAorQLUZFzP6m1eF+md0w4tju55Ye2LamBl3keI1
A5XDRLvUuVRlRhrFdXahpWomPJZzCiHTfSOEs15D5qMAkmCf3k7GRW3kPeWzSEkS
udXGeHCi8MkRAhDlmTFr7QYvJP8g/TUceDc3fJmExQiPoTM8O7FE2nq4ApUrUe4V
ZenShltEHU4f6anwgjAWBZ8sV8S53JZMfpGeTrkmS7cQbg4AFTvx+yPbzw2t51rr
Yoj8cybN2qfL6/sSa6AFOdaO0bvxqOWhlTjXfgYTRHyx3DpcmQmlBrvqHQM5UyMm
doy1PHneeqirpJT7J9F8uYo5oVp78YLJFMhv0BAM7Z8Q88cX8VD1ToK2cE4WyCfH
Dwtz8KpqjqmcggeJ1IrD0pJlOadYAIW7OlNws/+XouM9bP10ALsXFg7c9jpbkLiN
8kvpVeuLf2N32IyInw1BH7zo8jSKAnv5Z0TATjjwzEc8qsxm2QpGG6j/tb5pjxp5
PdnnU0u1nFiUmO3Q+Kbd4VWMSIKvf6yuYQjh6tozvFns4gjYjXKFTRcyUyaTXDq4
JlP4eOsMZSDMvNHta6aGT7xM//3cA9a+bbrZau7k2cN5l9ULkhjWx7TxtQczT6/5
SzRka3CX7QvpoE0PnP9XM2WvkYJkU6nsiTTaAMvtmFfkhc3g1JnAQv2FDAAOf8H8
ULpPm53x8Loth9PzFjHH5IGvBI2d8FnZtv7JvVilCeispAUqfJl9KolXyv7iekuH
wKD384dhVNI4oijmPzbY+IdacWO4bvcvCi8H5C5D4J+3nsfLeqUgMSR1BCXBjtPI
RuEsmzvkj/1Mee+ATWEuGp68Zb3rh0HXdfDYUdnodeEUyvMPc3HEKiiP/btlNL9n
0EP6is6CbIlKIT2dGA5I9g9wUvzxVM8TLe9q3MeRz+Uyy0dkibvujyBx3Q0TpYt1
Pi2nv2PPo08xoTr0bPqGD+bLv9R7UP6KbhLmoJQlk0x+wDzlCp7FHwwmbyEjdaWm
Ej8bTwnggdp2U6yOgMEUUXugpNpxSHCSs5aGO+xO4knEKEDhO8dC2Q0RDudKJXD8
fGP+cCmSNSIay+XiAmVjfoY4hBZdd6RTJH1l14m1vvO0VNH5b6e/nJhDUqFdkA6W
RF0H9TFGdoPA5qVgCEHv65O4nknmU6v4MhZjiwahNhLm0fbGaE3XlRQcYEzsyUL0
p62WHwCOXhzqo5V/algL20SsgNIUD5c5SSnjqP61b9VwoJ2HT8xEvOj5NkeMeWgR
O2MO9N1Er4AbUBjYp4JaIsXUQmW0Js3czWDC6zR/5pWejb484sqQxdUz3QXN+KaC
HY4YhNxdrIeZryONTR7sOFZAVj9hpMt2Bq817hWicysXIHEfF3Gtq+aep2lKq0Vs
unYCKj0FBhkwTTHBRpp+yQGoh6ZMqzLR9Rjy8ynXyU+8vHvFjWFZ8qj+ymJxC+7O
pJ6SmhEZoO0Gn2QsHkmzYtKuSSJfb+Jp+4bMsf3FHWPZ/en9C27HAOQlwOetsv8u
Lhyc5pdWnP1uCODviVj2f1YeBgAIHME9pkRr3skXP92cNMv3T1LDjFHxx9bAfrEA
hQ4VrxSLIXR2t5fqDjg2YVOiC1rvQqPBxXsdnF24+WtQ5EbH+jNvRY+2g4EDi+uZ
TTwi0N+Dts2hf86NrGiZRUb0IsB2rZh3u3saDN6MCNVJFpp3PMq76TbdzDENJ9MG
CeNYMLPjWS/YuUfnW+19Q1t8s7/bg6Np8snErU3rkCL1tlU0impKWSzSaIakhA0u
+ajeITWwGffXugCZa9oOcjQ3aDvYcheg8k6f5cyGyFDgfMU4zy/lq36AAT19VMjb
zVB0h9aUyzrFLg2aRZkRroXF7UbjzPgEPEeVEnUeCe9/M4iNn61WOPqLWQjU/T8j
2acWDIOldOUSfEznZTK/A0kd3mporkp7pCrJCIb9/VNztYCj6rGBy5kXFcfuGzfw
U0m7AEpDmz3lInFWpH2tO7Tz0JMDPNT5zuvXZewnvOSHn7ylIVT9RN5wjLKYJt1L
tSod9SFQxtdIgcl9VGhKXNGb3pZuUnW8BHtbH2+Zqoi+aA1hj/hvHX5cPdvL0lCo
dEbOm86VRI8pGRPVmPrdhe/xp6zSwXF5Hge1OEpeLSKg85thSw+uir69IWECADpR
FdDaS3YNt8VGXEcBQ5CNjeaD6y679MIEFIPYU5gVxpMHk9AyRTC38dm+Rb0Mqqsm
CyuQt3iX6kYJGtgA32LXy92MGo1yPQXcgfO75Ddd7Eb9ozThm17F+OiLcc1I3MTz
z9zCMPNYkF3YLUenB75CZJXadscOYPYW4U3BlHFU2B+0N6XtiswCYjhYbXdijOUH
gDM8bDHvwZHRi9Fy5rIiebYrahmsLfCbCFeva1NGjR1R9LtvR4ZaSenSeajPoZXP
ETzRH2kCh5xKN6tm7bsNyz1K1pJM8kfYJJPeQX/QXuYpV25PFtA5WcRiM6Kt3+vK
njVaek7xuDlfDMvNwftU4k5p3+2i8org7qABTkvMPQK2I40Cn1q2+Sv0u2izwM/a
dNbVaM1KMM5JGtXQp6kQBYdjUK7iU62zGvRQhFmqokl+b/fRR62VtVTDmUPnD5A8
E5B9YLaAIAKzcsLPpRgjqAY77UoSbJCNyWYgTRopMxuqhnhi4kL63UrySQwfbnMS
qpfqhRMCmWUEJ2yyJMsPJF2Op6BtqsRFaESqxaiIgFbzrNbkpz/vTMemovAR/eZU
n87R6x10Rg5sns2R75DT5EHXW/7XYdT1lbT99mXNlqmJ0Uvom+4Jvdb7eh0uUsHR
TdlC6KW2Agw/utbJ9ibaKcQFm5qRqdFWs/ycWlsWPLwBi6Lcaki3mDEsOCn7qJxO
g0LZm3rlhWvsugRyecw+BqmiY/HcT6wp5pQedKeEgW1uaSma1ZjfUgPA2o0UeV7o
8F5XCLKds78mkpaCfYDHUHqv9ZhPEa91D1aMA3K811sqit6V50/mj6/1+d5D43Ls
UausWEEOgo0bYynl0Z+OrNq0aIMxgN8qAGqD8R2OfpAvx9jO8KMn/ZNwi1BZSXLA
2vRObaWxQaCsx9rFRe8Xkj1AZeetZPG3j8qJ/PprQfNWlzCCg7g11omv/0QRRSdl
p2QHhE2Zve3EdQVoT/yxcXuM+JZy32ziTHEBz3po77fvcfLMiG8Z70RMLUDFXFxZ
2L5EoQug9CFRdYZRPDwXNo2xrKXpVcvv+PNANcsF/1WAlKvZcW3eISVZBiB+BFv4
VNUwE7oE8taZUCDo845pFksEra6X/fCuvIqtLg+wnMQ+xfy3+mZupObsj2FcjwCD
+finsrNLnaikI9zMIncqkNu5FWMP27+PhtxmPro1/kP5B5qaxYSgqRg9zcjGkTgm
t6FtxyQa4TfeU1eZiny3ZBzRu9h6+ZkiYu++BnWvnJHwIFggafGzqTgrG3jVud4W
Gp21xMJyobNubnUc/0aXzATWiv9VtGlVPzFxNb4wxCt8e1DS1PyRKnv4jxzH2MHj
h+SsvmNO7O+SdBL0ZHk4ZvVd9zc6PmRNYrP+jF1/VlfzgQNANjwBRPODFj8l+Oo3
5nWMfSr2gWSS7qbw29JDaHppjqUYju4/alfTHyO09tchQQPyhfQJHyb7KfzmCoRi
8DdqC0xbB7tl16zONtzl3l6Mt2s58bJbeySObTrfbLpi9WnA8G4jyPEmx9loxhIc
bDrHRlvWUCWPNKA+90obgE9Gdra8SnqKSv08HXJT9xI3W3gbavXiWeMutm/SC1fR
agjaQ8mODIHNI6z+Bfv8KIqsvFMUlzZgwq0rl3g78DMGLxrXwHVdR+EjwM7kuvUs
NX3AB5xkhVpIbrpHqMGx/uInnlNOzEKCEvBEzK6H2oruqVrbYBzqHwe42IL+LJ64
3M6cnTUsmV6C3EIXf5HJU2gvNMbRfyZZ4EAZ8v+F5S8/s9hz+jN8JEFOIZdpc6zY
kB759g13MQOE2k6mTmyXx5EdmnXapuaTVK5SZNIRVDy1oMPa0/SPGSTvw7x0HuPr
k/m6uMcvTD7ZkG7zT8QYmwGRd1/H+Ztodvbxbem0bYtnQDVLvz+2NwNFNbWodGck
9LGEylAYKUuz+JjQP1JZzb3ndAqD9mVVKZizVX+ZmcWqA/C6Vzy2s9LoO/927HCJ
34NXMqH6XApq9RDFz46DYtCB1ro8psfRcVPkfS6FOBp4sOQaOnLKMovqv0MN2s7M
ecYLUQERhknMt6AWn4L+pCn3Ez1CLu52o3sGcheMMPExqjYSHuXYlLPw28rdARaR
ObXkzgEB3VTAgNW3ztIPDlC1MXVmlU5XTA1+onuZCGBg2UXPBQmQdXs/Gci1fva4
/uva9gAJEwpadUbntquq2nuctHxSEL/LOdALvF9fuNhRg0VKY7cl7LsrPe0IpC7s
VH7dfKSf758mMCANHuNeebouWrp33jlnQmvEXfEV+BC4Pnyo8rxaaxjxeTNqZ3Ws
Z3HMR1FxvCUgHZEk0TIETuegnRnb5Teka8PaPfYSjSDEdJsfVOAoSgCpZF7ghjeU
IT2sCLeEnFsP7r3JynmUjxUnDfsXMN/nTGf0J6Gb0ICP+c34uv+g86ZedVoJXdJn
8cd2xI3fjVqgAYNshBAoUU81EAp0aOHno2V4hWOuzlFj24DoZmgMbtcSa7IAOY90
iu228fSnytxCFa81IrpE9pL62APd9NWRbUhVqCVjgDnAyUo+/bivvr3Z2afSoWrc
kgumh6yWjjt0d7mLk8nqis0r9yOgoSyrc+FUWOZAisGp1jFFnzZPuRtl3YZFGBLx
GWuxmKuLAteWe8sWoo7evJiTIOJbZNopWNVoYCdAfvVsZXrgJY9FN1BCbsuKcS1d
DS2udqxCFOX+HR8tj5YW/UOdpNxhUZsHaPQZgEq2nJjKmYZBYeXqv7IV0vZuhJP0
uDUvse72Mpuel9VnkRsZmW0atxAN0RZoNu35w2kbHp3ZzbcnH0Z/luJM9ITNWrMc
LFK7wElU2BbVaVad3vKdooq6kqjohjfJ5YrYulGCNu8VLM/cMdrxutVtgRmCiiQ9
ZhaFtdT+3XLkULO1jPYS86Jp9bvwoy8pqI2cKRavmPu5EOK5HYSkUj3bdr+KayEZ
k0E+87vIU/Cc4otTcAtOKGdcbVHHw0TsPnlDfIvVf04OkZoiHUT1SCp52tIultJ4
7/G9j4/9oKD5rjt3/tZrttacJ+1yRWNoX1ydWEH1p8Xfx7rXVdTvzG4mNovABwJo
9A9By5wcxwxU8gietut0HjOugchJPH0A0+QgeVLPqf+N2eN1aFYlxHXsmxNO2TzY
Ar7j+TvgFhQNieoUtkzt17NB62a3YWHpYCBYYZCUdxpAPM8bPKDMznm+swIlTIDk
Q92+87zGAV6dJpQUV4cYje+TtFjZy55c7hb8i1Ss6iBZ7IEPiHYNLJq5J1zchQsY
XOiGAhBmQYeVsDAIPIcWE9bOkMgNCVNlIOxzwfkO3Q89SKLIqTmZ88YGeNba5t2U
DHQv9Htu+UNGDu7XXvQ7JUaKsnXTK5hVB07m4ncBO90XcucPQ2Q8UsoZgq9rnwin
OZWghDmGJdQqdlFgU6xi3fqa1NQCDM54rDRgg+wXkOe5wQW/QmlQtgbraGy7vawN
5umY2Y5e95QotuuS2Znm3QEjhVN9lTdxBPfAbFOpUQ1NPcwuGmw1YNhrW9l6729P
G65j0OKooT462eTHyOlwupAtBAXHTMh4bfbOzjFMvksekc3lEp2QmGPo2Jz3J+OW
pf2SI2stpM8ui6ocywDigDd+Q2sO9AqKvCcYKAYVKXYANyiazlJxFxgj73hmTR0T
dnjVKdYtc8VIdXzCukr1uOmavel9LSy0ZKL+DsKNgsNBc8xtR8+0El1DRriuN6wG
N2BdIChxy4NMHOamexrgbPss7xO+c+Za7pJcmDfZzWY3CFrAUUiZlswV9Ojm7cI0
30jJQ3txPP2PQ0hKmaDqWHks+ZgUrKASVqvFh1Qp9CJU46u4FbhH/R2rTs1RiIpx
ltvUyx8YlRJhgBA9UhgICtCBcVs7RJJKIqmrNzHpSIx7IydcomX4dGc+n++2gz7C
MtHIziKc57gBsT+7WlRuqSIsNPAd24EyoQTOyCR7oe9tKRvnn22ZqLj1OguY4Sxz
wgD73EEKrwWaVsNevw1ILXjeE4zM9VHVTG6hC1QdxWxxAuTWbBXDmvTrUD0PeOD3
aNW9ls8jW+vPBOIAuNnx15OE4C6JFe8hJeZIxRl3qWT2pf3f8SpvVeLiqnwQvy2e
fAKMJ9fto87dh1L9BbKCsSVEPcOdpZ1DqU1wldlcSbv2ed5scWLJ4XiDwekQmfyK
s1gJsPCNEbNvDa6OS2QbIdqHdsD8E1PrEHuDaCaNmg1EDqKSD3vTn7CbZN76qerE
uad58nhgRwHhYaXL/XOa5hy2EKorQY3Z2zpuqkEqeXY0JbvkfSyz0gbXj5BYQWqH
N33QtD1qnULITEynax57g+/pfgXTEgy8qMmOc1DcJdLEaXMyBbrf65v8fjcKd8el
/J65QvPH346eNuhaMyPhrfUZFYuIyfDYGyhHXEAOnnH0FoeMvRyut+vObXBNuKla
UAgmwW0ZAfA4u/eS05EFQrJq2OTrra6tYHSUHnOSznZxjV+TkBzgSmA+Su+BCCBY
WiNWRGBI5DoAzz8GLWG05LG9NLgtU6R2WXdr4lB9Djhz06jyvFijCw/gvn25uNLL
Tg1jbBO66YYxIQCI098B/ehkNtz6KZrkQGnjpUT3MdZiCSdX2j7QOgolekrREXdT
McP9BVQYSaKUteZOXiv3USgvvF3Dcemyz8k8YQz9EQlkYCSuOmuFE22aGZGL5SWq
s6+Kq6wQDmV4ifi+9apbP69wZ7YalfmdE9ikcZzdAfDx+jZhD6dvewNPpmX32BMp
vNI+EPM71xq5OiKyiJTkdrSlSCE4Dg2v1MZQtM+ghthyd1UoiQbt4cwKT42vz/10
LmQ6b/OK1J0VusKEfODsUAtaXY6dIQJPKnc2cpHivdSK4apDqCZueLpqZ7aMmi7V
zHj3Q38c8u0760oOFiR5Fn/i70SKvO6dUoG1eDTjFWvKM6mF73eOyUPuf4zIcXJb
sjNqnmUCks8JglaOo2DgZyyaj6kXNFH6LdyV+gwEv8pmBJNqspTrDtmvViSD1c4Q
xzx9ekg0epCM4YVyRxgHOxFBMJMoosxvv9Vpw3awFwhoLk8LccPldl+P1lYbuQKf
cf/HQ/58M2eV42uZjNiThWW6H4Wrc8d/j+/vcFo8/lOjYkSEdQ7MbN7dV2Yo7GUp
7J3dSoNNy6KqBeXGN51uOAS80cUGq8D2TYp3gDxj2vg60CsWJHOBJdpCqoXr9sCg
S8RZ2AHIdQcfAquyARIlN/uA0CiqM3IuVj6qaPB36+ck4AhT1d6Go1Be2rgD7GdJ
VNgNI6tPaPeIJVozkOp2vHpjdQGKnHUoQ4ETjrb0w3Szallt1w5CAtgiVUGhpY49
XgwWuj+6+JZnm5okJb1LeFE928S9DhKpPhKwO/9qXRrhq0BAzLVjFwrciewnkIOX
jwGgcfEHkYOrsQuEIpekxEI+lyOAwAlUrf2MtK3KCD0GFH+jUUoVveyUREOOAlo5
yfsD3D+OgfCZzVQNwv+LZj9LqJGA005fgyB+QRDsfi3xTSyXOxtHIwnc69t3Ieoz
nuBdj2UjnrEk5DX3/XKLypK7XFylA8+mmFjsovgzAlZi4lK7BWMIL2UQZQrgRfX1
jqEpfcaZlSXAJ8IPs7L9JZ7plk636waccwpt+9QYlaAyl9wBGHn0eRetcuKzWEC2
6q/cCj2tK9+paz8nebU+w4sE79E8ibKauSoDE4Oocjd2Y1bjZP5UlnyrbVHiwE2S
QDkO8ybKvLC7K+sVPX+keBW5LvWsA+XNnPbWOHLhukaNKNZBoB4zZzg8+WMfDoti
6Mis1yVeJQ8Mh1kUoJQbaiXLf67TKDQMeBaNP7tQt9SM2JpJYC53DPs8NrWnQF22
fHBwkl/MkyMvAyWECAzxKaPbRWXL+tIEuHViPjQ/RkTAFDzc3u66iGh5oe8tYXxP
jqHGOZs5IaGzJEcX2mrLKOyJEOwhU3ZSt4nAB7eCsABEieiYJTOt100VRRtEuPUV
HAtof8b3ndyXaWzaVtVlz3XYzxo/68Dwqwa6dNyrJJOqUhIsr/JuQGssP9QNlC0i
tYjem1RYPK808rUxof4ipR/kCl/rnU5TeI6oS4GujkYr9UusQ8I0NMLYpFKEdh4O
yMu08tu+jgYxTEtlt46chV/OYN+gTZjU76xQFmpgWUiYKK8MR3/kYoNffe6ZCtIV
2fcL7vwcotb58UpfY5k/OID3hwpSjRiZfmkjscOOFJWeHXnOld/sCdu+tRDh5CUC
PqMADJ5eefWShehbungFjQ9WfVBat8L5jApmcu9vh/CFSlEf66WmVvq+KGALJX6r
XT6WQpHZAdvQs1L18ANBMBKosmLDGa+bbHiDGB3OKqUKPmtVqtb5PMbU83AuV2+x
7yCs9W7dP0cYrSboJBqOS7MGRhADLdIyWNDaFEOkVPJ+K5HwKNHYCLwE4ywpCgQI
ywRFpTWX862bJA+BbbTuDSWF5yI1KVU5mBUYI9hahnun3VvcV3Yldwv2/YuAwn09
6VwH93lbJZGSFBtp2Pugdumy7SFfhC6XuO7i9RIek0mgmJIFfbHYClwh+I+KuaOe
RzdmUno0eytv5YrlY7+x+l71pREb7oMKDHkauc/yC2C9Agb2eqhR33WkjFKfxcRx
eEzC/G0cHGkf6quxInCgH2HH+3SXuo8W4daj8rtrlUkldeimsfXYxafRcH4w1Hn0
8ONtRp8pyaJhvBJYcEuWEI75gFCjBmFFEqee0rxKeLLUNKOGoi7X+AkInvuah4t2
92B5wLqOSNCo1zV1Ula1BmM3tRbMIp8UK8BtFFWX3ko9Ox8ObmvVgf77kSpHfzGj
gwqK1l2I3ZiB62HNYTSHZTfUBaSkgVy1TQXGbd9HMWd4TKkkVDfx0LdNBE+Qsda0
/0cB8logWpjkcoC0V0yaeJX7cIwJwTHZ3kIJ1GYHGKYfdB0526RuYt3OVBiDe1j/
L/wybKPMeCMFWP9EOtC6cl4mMW0x8d2ECGjz6KfA300F2yDmoDBPKk5/sYxdIB//
S5UD+5vUUavCqK6X3T+ki5haUz2JelIt5P3zTG46xT3j/OSC1DQQoqP+7K8Pu+fZ
0cD+d4081J7qA45wyn2JoPHym9eF8jYpT7BzSM/fkh4Q9oC61BAlX1WQ3pZKF6vj
dCzXhob/oqH8IUBMGjIVta/v6WSKGrCDsGwZ/+N3vOHvqHPiJXFbMwEio7qfyBrd
PkXHgVRdPUVIPAzTkVXzxQj2hes5qH0otgmacHv+H7MpwdTPnhWD2HAMa7pV9FKO
cC1ZVm0PTRg6bCmMQEtCSWbU/eBVrmswOfnbApI0MnRGX828o4tgzvPGDBlSalpz
k75sTa1fzB8jZMDzPkP+R/eggcHTFt0ANoNqTw0QP196+CfS5gVRvxugXKpCmtqP
WNMGgwtyigN86owrh3mw2HL+JZhlfMRSUztXbXNbDsp7ZcR9gQ5gw6kumKqiCCen
eM6mhZB0Lnk0w94Nq/sipmUwFmoyw8Mq4FQcn9i+roH1s8we4ct7W0HPudS//dKB
ZjbfcsyvCJvPb5FZfSygeLp69AcA3Y6t8I/b1mgIVGnMhgDLUIHzNA/QsY318WSW
eFD9lsMvTDIac/CQJDWbSht1VlyyKTGq9X8PaNGzqt2VjwQB7APGHleC3LL7MfP0
rhXOcqJ+bnpJJTgZ94cIx0DVkntR8kj95Wl3ur+JEGS3NjGWopfU5b21NtGsAb88
CxPjK6rMds1ju+4tW29hG6S6ckYH/JqXqyDUv0jfHVQPyaYYl72fWP/d6bRS0qOq
0lUv6T9YAFX+NNEkaOL38CANRsWwcHGX3iGs9d2cr8gH34ruAAlHtWw9ec2v6ZrW
X8xWEI0PcSpWijhm1ZZQ8NMbz79Xd0zBTgZBfAdi8co+bbGt0NtqcLU9rr2caQmr
ta1GtCPKhNMaQdH42VU05qnQp0CLCuuacVXOZ6STQMt69dmK8RvRYIkA0S7rbcKI
zJ+ecfMht5Imeln4R+ZU8Ni1w5NHZPColCRBdBUMnpPXEsj95WDkMzi/P4ppBzdn
aBoIpqRTkJBZnO+NvUhlMlYbt+rRcekN5w/Kpqp5cdjPJUcSk78bjIAG0xFKWKlf
sjqf4ka96mKcnbEwClieLOXb1irGi0um4tcZyV4Kw83N1sjJt2X5vssf41cY/tHs
vBWIHzCyKM+imjRR2oEWjJB4DHJowA4c84lSH9O8eJbHfxkyOAlYaPSmYFyZ7HF3
8XY2j7umYk2uPdUDm6gJMurKO0TM60nTSRA7TI5BLG63wUNOeOfhFTBqdtt536kd
2s24jFDqN5qn/wEmUIpRSphaH3d8IV9yoYG2euIQSMY8XAcgk/nhmUaR1N0/1U0T
gNrb9hmLA5i0M6lMv2sGki2+F6IwUSlRIC3o1PvyFAktJnilAT4AhpnmuGpbrthc
HCmaSkdXpD+8oaVdqV2ZYvZhe+OMsJUVDXKZj6brYig9+jvPPKiiE1RpxhlwemhC
KK1mPneoDqA/QSAt41BUJgreqzH+53fU4CMcePSw0vJ5O4JTfJsaWeQ7TIUkD/+3
EGkrALQqpx7w6mOqB3SQWHzhDwhZA+Neuua9OZqnRH2aN6jLFNp2kFpa+hUTmZz7
e4ggCJF048p50rG1i1KQC78qGYnIX408n4Zpn+uF2VGdngY/5aCZ0C7AHSVWVVBn
3Sg2hbndQmvBog2W90YlJGFoao6GOS2AyFlotRtJ6rvWKbpuZZdi/fPF5Ex2hsHn
hxNDmwWSXVoZgVlSBbjDDEIphPWwtafMeyvXvNmmDkTRJLa9NPjzuJw3rzlhXOrm
2EPjsJeIe09VIWGHu0QmN97Xpp4uu5dpINGvtZynVTflKCmI2H+hYRFaw4Ryeaci
BmrdKG3GgrSQLyYIwm4dtVQ6Bd33GgrQ3oEH+ucwiHYB1W7/ae7kwpbNpkGdI1Jv
qRh7QRO4rCctr0zrRkzoX6QSADX9Il31Kv5adK7xSIv0WtWBLwskhLVDiYhxaLgN
h5mkUQv5Q3fB0g6Br9o5QTC8yiFl73KzhrIUl7ahwjDzFbvEt7RWiyx8JeXORuvP
DyZ6sdvuQ8nSbQZx08YjLaEo1Kd5c8Pi76lRK3WCQaL4IFrWMroAGOXkZhzZaMd4
tyEKOu79wwNtWqk4cflqcEypJFto764pqHjPsFwrIK3CET/kiG/m+NrZK8bHma0I
n7DQn892gKmor6k62UOxtCn2IPXYAP7qjKYBzTLECcVav+SssIht3Eejh26TyQdO
/JJCfBDhOWuymcWuQT7fFrl0B71mSa7e9UQkwWlN6PlbSJx07IjpYnGRuAHUykzk
Ztwstq6XH+/SURisqn5WL2A1EXaYRd8ZJITC8+4rza5hEGyVwrynNBPyHWTGLzI1
x/UO1rpcnTEZ7MTB1irwVMiCEduGkkdJtyrEIK7/fjgxpxk6AJsJ/Rx/+UPa8nHI
q4ValBHboW+8/YRL4Cv7zTqSVMnjFIKU7+KBU8MQBfISmrcBEu8m07l3TqWGifkb
26yQbJfxOCqygpa3Ks5cdcZjwztJ2JmsKocPXOfplVlEPqM7Cyi/d3ylmyY4Ra/5
snrsk6YseuxhwezK4sE/Pz2k1hX7B+SxZwa1x9WS5wg2Shb2Nu7lcPc7Abt+16LQ
Ddnhnzi5F24BU8ohd6Y1pxBRjvSweWFPQqY+r957Ru2fzmO759hESZsqO+F45jfE
AJ0EZodx6rj3XU2zHI4h0MFVA9EVjuhqz6zppspF8vDaYA2kIW5fzAs3fMbD82Bn
/onJq4CKGCL2sapSVa0usysMQoalmKjZrIQjyfAWYwbbn6CGoArA2iIZRYw0lhkn
D+4lWBb/nK5ezkSZVz8UPtgc4qiWQFmL2czp1/u84kZnXVb0lEpADLDyHnaQwIp8
Tl+YhHlLeUxH7I72zTifllxmlJIyR5GZFXvLkuBV03L6bG+Yn3LSKd+3PaQcS7Xw
fv/GRDzUGs0lDqk6RSCmXqU9o6hps4acdRmzY9iNApLI2yNNUU0QX8MvV9KwMhmn
fnlLwpuGMkDldmHDMIUQCT8mO+b16SUySgGIeJ4CN2FfDAfOuWT4CijACJLTtG0j
TWN8iIhzwJXNx6UxnRgES4LhCBXV3OGfXCyu1hSXe0broK0dzxhFZcx2nWcEkrzl
lgbb9ZCiD+jzZhGTLIfNVmC6x1SKR+h9Dg0JTHQTwATDjT/g3OQPcHRbjQXDTygp
Z+BtGfvCToLulAH027SZeVXyO++iFzZ+KhXylkCcuAe6JATds8saW8ajs7JQzRGL
TPrC/DxEi4CKqtYzuIBs5z0Mb/X0EHHbSsk1DrUv2vRWLPw2qAgM+DZIO9Ymzdfa
fSooH3aTWRwIyaFLMlzKanaa4atUw4zjc5OskT6GigOKhRmF/0RB8KqyJJqbYyfs
QjthlzFiKP6+2IqJZhaKAAcAEgNtSuOXpzE/xdRI5dEDBOgWeqiPzNFdgT59b/W4
/nZvX7jDm0+rjNRhNuS0wET+VQQVkwdXxEp01MiGqBfrJJv8f3KVz7w3dLY5vLph
gCPDFX4AAD76i0XYnars9pQuoGxMpui7LjJBeBB6keRoEKbN8Ea8oY5fJr8lKXdj
NfLTQIkvuVTgelBeEsvWRBZ59sRDGN5jroW1V8s4M7alxfWEMWJWwEX8XvdLSFBR
WrkPCL1UHP38Co0+Xzd7Hp48OLHaNd/bVzh2t7TDcU7YN5mSXTtiAmMlrmfCee8h
52/y3IA5MNbC+n6HCr6Vi1bF1YlYxr0HPiiADzfs1jO8zbqsoXzfkY1cCt1AvoqI
qqkb/umDT5qP57By4g+76mkGYqvm+wRrVXqnco+rBnkTderq0ImUCAU1qIizxak6
+bQ1HUyTxtm3lkNQmmZRMnJFxnMD8gCFttoB5tP8POb3KbI7GG/skT1nKS4TSv/X
idSBqa5a8cdp3tnEIQbyXgbESeCDIV5XBLkTrv32qZ/kizx2IRQqZSD5L/rw0AZk
keoulqC/YDz5E1o3bBqkz0ljY6TDhWvyUha/ksdglg7bpen6mNLzBmSl/ulwq7iW
Br8vY9NcfoK4OjiXy/QbIOtRzGDTWqZwb/pejYYiYNvyEi4cqjvqq9WTVp7IH6Cj
M0Gro/OpzzBB5Z0h9nzbXyI02oyelxwrgT5S6m0okNquGoLupct30VHmw+VPPOaI
MpnN48yU9mE2xdhfMTce3XzwHFIw5r2Jkd+N0aVRJaMeppSn3KgNZApF7umbgiyj
jj35W+d0w8aH1CE2MR/9Pna6mpuHTjzGUx+mobMHnsYcUei3uJlTRqJXdRODGZSn
RTjPXcbMzDgGmNjincFfaXFOFR9mHGVlhNjKZGw4kc7322IHbEMPyIb7fllgr6HP
h8IXl4dzuzSvrHIIRg17POQh3gBbfo67HW62NgT6iTZ/OQFbavbSk45CkCvtniGI
rSrQEM7JSwEA0U4uimkrVmPqzCtMVznvYI1dMehlZ2o/RRK+OPCk9TftQ8A/I2Pl
FNHFaYvPMU5H3avbDjtUA4hMaO+b2ONgga9WncRwmoTfhcK/fHBeI8xEBXYY1swG
NsaR39LXKN4Pdf/zDnQUrQkSRMfw2uKaVFGeYKnnuVbZ62UEA+642+1xzCp/kdmy
rmzjuFcAd3adY25obdR6vWIzSQJznonlY/YTuhW2MqaRUSeV1E81XlumeAbDfoCW
Mji2pzHDkBnSbijw/b/74qk4AAPghfDp8Bc6f9FZhYYWDWMbza5OacaH8N43OwRy
DLQ0lZ5bSW0C9thrBqgRkQhUhtqDt/KVIyQhlYWmjwq8RJy7j/SJQSRsb983sYJV
TQC+iyK3TOjW0RshxK4uP8MFo8VH9HZ3mEIQV8kUrgfuUC9nhx9sA2cWMhcEJW6j
PdveXq/2Vzf3SWlxmBtqqUHL9c034P36Ed7RVxFBmXI5yRemEaC/AieySArJZ/Wt
89+HUc7I76ipTr8FDrGa5niLzDFAGwc65v9usAj+4NMUh8K3Kq1wyomMsNi19Q/p
ohM859L/Gd9aTql+yisYD/DApR9PLMSrJI23ab1qwXnfBCNFFzvoAjhx3RUbdnbS
ynIckspky+kMeNwW11oUQK8st/H1pbvfvYdPN2R8dzAs43rAJeWoMINzzZgQFim7
aqxkaV42PX3CwuJ6yRbcM5NEgEzDhXMfKj74RyE7xMC61KmeRdtFDSeCw2B1rsKu
dohNL0JVX3u/S7Caa2k4B720re0KmqG9BXyVQ1oV+EvXcJbyJtaCqA3XSLKIOzKd
9vHTfBVMLaTC96DRUeATKbGjHiBzJ95eKR04INIECUCqTXsEKps0Ig5mOSDHz/PV
yMQZJY8TUyssemivi7FLfmUa15NV6G295/aqUmn8Sf6+saiIy7TQ9kuktr+5JRPS
XKhWVV3ACOD6B0C5gSSbVVpFQPQ0yu/AxhoRieLL7Hb54vZ1qjU34bHn3JsrElQ/
MgaKKeNig3zOOs5vo4iy8NuKwKVMkpE6YzoZ7Ch40ETdBJvIiF6exuIXxCjea730
JYi5dF9xMlFN1O3TrgaUnbmxCUV/+D46saXLjsKNNIDXR583vWCauTCKQyc6vKgd
NjZzGugnr9huKXipz8I99RmlTSRZViTW/4dp9q00BTS4UUopwLEI5rzsOE2GpV+L
cDm+Hc38gvW+pK+60oMEsZkiboYDlLivRtf51nYkomdur+f31T+156NsfbzrQrVn
wmXmZK6YBkkr8NeodX+QuG+oGFm3TZ/Bc54BgcMSWNwYCpJFV+l4m/bDCmZp6sx+
j0fDoxZXUQA4G8Vg2UKadY88e8Lpa7noKZin3Jy665uBDtis4AedKH9i3YWtLtQu
JDelwfkvjl4cVF+bHg+N08zvNCZ7t8tDhu/8+2+gU6LVWIU6EaQQXY+EDvdXkTaL
HkTl5hwg7jhF5kM2kXnGzTp0RtM1oOL0ZKuMxmpCtptMID++zKEMf67PjAdy8LUX
zIaMYxbKYS0as5V8vAdgTFpAx1GrmRODfmoIkmJm/VkU1dletzzSXF17DY2RJbt4
l3QovT7D+WV4Kva/ERuhR02UU36BLJ/qKR5/YPiPvZzmy6qqi3lpbru8oLx79L61
xy8LlSo/QUJmoY0Nqq+ekhDugAOFxD/TvGgHFcFzJ6uGr61ay2QxRJz+YBR9SLeZ
SIzx2gtk7A/OEnzVu+aCQyIdaLC6vy/1j8vO45zbwQr0x60I2bZKHlLaTJMZbZsP
LivkQAlTJYWtVSwOZLZL4qtgqZ+en0CxxwX16TZ5TA2LWL3Yx/OvnL41OEqU2BTD
6JkdA73MYpaMITffWp90t6/moa1GzjSgrT0oYLr59M47hBEb64BkujLFuLvYaSYv
IiZl+GFcaTxaGDOfAKV1dcU/Bg/zuuH1r43XzsibcsI2J3MgxYwddxn0koNh+XYV
NKX20AtOz7HiaC+mkB07wVMZ0kkSlxLG0wS/SlqCwsbQJuQsf60hMuYbFsdX0/jw
O2Mno0XMUsS4TD3PUy4KwC72Fv30vIwnED8AF6wPOqY9N1WdfIx3aMc7VQeu3yuT
5AJM/1YROD+o34flyQ12J1dSg2XpPqFeEZUAP5oDxzvf1CxAyOBTB09qejaPTh99
hwoZa3M5m4Nf2Nn4yINpvVTzR5UmLutepIIUu6Ih5/pbwYLqyABwrz1eXe8UIxW+
yP+v6nfK3zR3tFafSiQl+qyiauFElIid87vVieUqxxAXHZyKP6cq5CSjHvmI/EPX
iFeWZ61JZ+0wR5G1oLdOXF3/abcUBebUVrgkK8JaNXsrBtJVy1ouIJPgw1JsYxJu
BOm3/5fONFfWUzG+o57g0qUKNJMoyXjsTHAJSH+H71fEM1rZr8iG3QU9govswzaG
hQPqNknSHC6VYQYiXPkAZC6R7x/aDfzybbMQSww6FRZ/ZK9ehbgexYkrZAy5JCW8
/f9RVBjttetyxp+bF7zGfsWP3v9fDz7SoHs4slQWZndkMlGsCXyVF3zTObGEIaUM
RQIph612CEqqM/DVhAoNT0EfpLhcbJjCJGQ1OrIYck+aWD7AlGtl36r0KSQeeDed
pq+UozaQLK+AvkTKW9Qdp59NJeN673mkemrT+45uU9vvhTbd1YAHKXTwe9BVzYFI
rQiq79PPyb36jqSTa6SEosUbRRnI6/VyPahIrhVOpdoC2Dg9W3SMUQbmptMG+0Xi
IeBJ0cZnGTgfs1rgcY8zuCr9GptWn4zx3h8DVm1AOukRB19BFJGsC5uVN53pZNA6
zkYse2pmMmFdiOCf493RBV6sSPEg2Z9KrywQSX/O+Op+0Y80nK6XD83PLKLmz6tE
pGkqhS3e23P8EFlFA8fnhS4SCWxHkG34/Zs5E+eYpp1fLYf9P07TNoNpMcEemSpE
b5n2OxTUZCpLXFqJglFz5nh4GNn2wWaTneCfSfh2lMEdW90JZ+Nr6VtHr1G8LvY1
Ae8hxNB9kA+0NS7+NWdz+iQBNGRVwIU2nt0KBhIkgJCHquIJHoHqUWE2AIX6ad0s
cOlbwxBJtpli6WLz7iOYPxjHtGxls/pA1dK8ECxgxNdCrCoMeKwjxgQQtG1xIrKU
hqCpiTA6e8/V96x3gRdUid9/wAqvIRaSvkOsSw0dzZ2KAPbltughHy3IrM3NWqle
UDBpjMUq7OYaFTSVFZQeGxRLqYPE1wanGtOn9E6U4L4w5JJ6BNOEv6MoH+jHVvF8
LzLLbxrrk9KQ4HCPlvU6QJYFpy2XZi2g1mZJxRe2P478CTBpAjkU+ALKQPwXeL9k
dEMpppRPOfSvHtuPuf7g2zldywVvdsuKKi48Ziv0+i5Z6sREHrRGPhAY8f+eSP89
Vjhm33TMbrI6ZTksx1tishuhQG9Oua5FwIis7l7pWxtW4Mmdj1FT36j4D027Ekwt
n6uR35ncRI2kFnDiz0udFLzRSrBSxlavoEFBM02TgcSNcFM8VNZn2XeXHQ1hLLCF
WwzHXt16e9p6Fw3ZKBzC/rglh4r9LkpKxTX9qBizQbeJ3fmAcc/ZpUxN+fVkfELR
UkaR2ePaNXxo4o51Mp1F0kGaiak1VSmhlwX4YKMTOWe39D5F8Z3r92TBRWAGyTdQ
f38v+RE2dbX/t1adbODxMuGNDuYdEfVyi5gxzDjXr/7buHe7dbQ2PabrTMXjh3/6
5bkDr6U6zsUOHO5QF3gBP+6zAI0BRsvWROYzYR/IKdcAFMyCs3QdBbV8FZrrIO4a
8cjMHA8/cI4ICTsuMaW3c9c9ygLidCXptHGMPDNXs5JUXLiSbpJXjX4LUFoeYqHz
MHGopiWaaD34lvMcvQLZ1vCqxU7l+gSqav+Nq1b7Cy3+RCAhBOZ5y8quhsoRM59d
PbStASQrz4mnxlZJYarsSN21er33ChIpaYgLyIUIZtGLwkvkO6s2qu2PLpCtntOO
P9uZUNpXKP2tuq+zyxFx7RM/yX3upEpeCkMwE+qcTNFIFgp+vYAFEiPXWNyVywz3
zd8MdxMTOa9/t78oqcRaTkplB8+CGKsdvY819IhbI8bCtaXlb0O/4T61EOtj1Piu
YOO3VdtNizaYQVbNC0ggPhY5DvSoZMYObMmGWeVJabUtCiP9jgpYB4Lb0R+AbzfN
XZFJLlms0/M/IcKF399gBUWgYR9UPHs6d2vVTZWqdu4NXiQiHgWT4catvlXCsQNu
OzRruZxKtJ5YtW06mwgIJ7VRyIGpmyz14nkWOq1zTfEl2tlPpgeBPiyPVVQWSLgm
0DxKWXhnw/5jVDYpDHCS13Puzwn2iMOKepuUMueFQJo/gMKu4hPThg8iaR1VFhFU
qlSZT3NBhHjSpDRN+KdBHIAt3CKwBlK3gpIjCAUypX33SlS5kogDN73S7/bfRLIa
VJ4NlYqRSW3RDdJiYt9tqaiHkaQuBYJnMrW87vkIF+RYopLNjbrTvRXBVwuYQq37
UJ8DDCpUfeu5v8QCNxWybJJQ5HQzledolZuYFpELVYUxAs1en6prg0eLTovZXKbu
mpNEy6Fzh1d2t377CICrQ71aUMVr3mMzRDO3Sk2pRaVHpY479Wujaheiv2WVO04W
NnVLstYOe1X9mKr5+fv9LkXHGHXm/69CGCCDMi6vjzNi/U3cnyS/64GzVcGe3jSz
vRAmLu/vvUCsUYuccr3x1dDfDnAhWlTbOjDm1L0Ys2F3VBakMzf8UIDorUkpIgNA
sNtWxUI2Drjr3nJH3z+Reks9LM4n8TioDu0CaF2XC3WcKEPio0uUziIvf7zlobvh
/YICnLbN2zZ5QDatUcLklMPOcMAShwUHGnOahPks/LCkuc88l5OQeNv9L/nFgrnr
4Y1RTFb+7HsHM97p5YbcYZpbxRVBugrNJqprIviAAOKYLyXQ2kdlO7wZPeP60DHd
VG18pBiYIZQOoXT27QkgI+8y4cM9i0ZdVU3YNOTAEuBpYciMlrRhZan2LJUtWbU3
fMEeu0HhJiJLzz30/uQ8BenO/cxK73JLwwZOjloNRbRsHl7M+0kwPbWKjgzzhq6/
dnS/YrmRV3cXwy5ZVPPr8m4QWScme8g5royLgzwp9BeR16koZcJZtn+5UfzStqlF
jmdK1JZBlrojZD/JffI5MVj2G1tBXgG1738LYUoEXhiIeb/6Y63iG/sSWOvOx9au
/3NbzJTYKj/5GfBLcGjAbaVn70GzMxVUatSj0wzQb7v0Gm89vYwmSPlGoiix8Wau
XkQDqZzzz2gkoKylqNulUDcrOVDRAAbvZX60PiGGaVjOpKt38iCedOr7UFB0mOhD
sKfaIFPxIB2nAF5PoI1j4xpeaS4Ey64wHktcaEPQhVV+Dsx/QhiIdl1EkKv6TjjC
2zwfaBSTvsljjBSBzE9IWgdgPFVOdS/dYqFQBA92F+HX2YaxVG/PB6mIi2RfVy8a
mSK/m71p168ZMghfn8IKA0gyRWIGVjCY1e2269IAb9zbAP4hIoNvoL06thhZ3PuJ
SEG8aKpzpNphmYJw5CBOcplAdbVFQH26/JOsMml4yyixSCKlLc0Q7oyc7XLq4S4c
nyUFPJlNRlOfjU0CRDRFos52mupfvNPK5n3CuVEUy68SXBAe+bRmjrJg3R6xaIU7
p+FIrFUTUmgK8Tn77u12/3NmIPpMkmQExy3Dm9Y9rN0qdc5F91FoHUz7apXS5YnR
tkYJ22BY9/2hvjXLs9s4OJLgNMGNmb8RvMGr56BABX375a+pQpk+RWhqMeZUkot5
tIfyd8Uy5gSK9ik4N5rs/6kXTtRKTEvPtiTGmwlLdoygtth9SaneZAatsKp8d5+A
hEDeHMsQVxyeEYZYoj1pJr0PPaqUDwF+XoUuE4aQhiD+usu2KhrChNTJxvXL1rmo
LnNr04v8sqPIhDpbYkr0yWydmQzusDlyyLTtHHZaWnZfQZfRDxizZDEq78Ui3A4O
E4RGIS59fC5b0tIYKE3W3TElg+kfUQyV9alsOtjiWH9oL0SrVnkpb8wGJ3wGuqWx
s/peZm/q9dlM7SG3zsE4Otv9U6ALp/p8DNG+ar7f4IDftqNOeI53h/iGRBqaBxJU
H3RMgANm202WYYwZ/lX23o6Pkf27iOSpiLrs0AE4gaU9jCPJPEcyWad+z1Oq2iXR
WrOHFsAWGldY4D011Oc2XmlThsTwgSh+Ae2KbJ0GkLH2vH8OnBHypf8fR+Cvkp8M
OLW4r0LQaNd4BwhFCZ6Aiup5DxI5c6qjUzEke950KCNMv2eNbtBJgMqUuowp9imV
5ce+5PJO2NIDwtYIdsuxuADI/7JB4SlCDSV46g4vdbxgVqVE/TMsT0iX+BqgRNWg
2NOmD6Ns8P9RDA7d362C8ZRftW7chlI8jSKTNi+H4SA66hJZVB59m38B7uG8CAHn
kOpZRsMg6Oz5/1FVdVepFx17S/bVB2kNNTkn2jrQj/Tp3rtscDj/h0YXAlyvbczD
pmbbDp4mUv6TZZ5nJyt+G3PB7NmyxpHVIP3iG0UmLu8uVoXzpE1qN0aWKLrV2BEP
SDJQHp509f9/68uJR6ZhycizLfBRgmatHqWLXbSO1+oudnrGHCQBBTiblby8cQ9G
nbzHLwYCnS76RAWlKRH2k3cDQ/pHNETOkCLQqPHhwtbYYJ42jtrl16dqS2+MA5UX
H7nDs0J119BlxeL8I3HOHQ2dGlldGa8ei0IvJv2q775dDaUeanFAB6JYZPp5TR5n
xxYS2cuS83PibWQAqNaYQ8HuQj0ULVHPgAONAv7d9Epega+mj0oOJvxyHX53fDzp
wApT2Fr5vtBAkjPFWfZsmK2ibIdn4oSJG0YIcFk9HMebhE9edlhWOUvbswK2GyQh
Uil+EWg0SauMXUMYcJ51ohYY14FsC9zeLRxeBd69h3y/ATAPkZyB8G4SAw81qtJ9
g3+tGrW+5Zs6fM6eNugS6iUoKysUapjeTYq1HlNIKXYiUFKwN2QFLlLE9uKMvNde
3R6t8pJfQjpi0V6M4m2j0LzwSxGssgtExN8y3ru//fenIQkXJSYeaB/6LsF6KJ24
bphbZMuyUSBRkHomd1F9VVHiIeQvwNbkemkAPkSuAa1Y9h7YbceqPKTL5V35J9zQ
rtdcYG4jxuLLZBn/cOWkf/e4GNOHPmGI1LxltTCOSUKtgSY4uWTYIxbDyCCDKLeX
3sz2qWsY/yUa9GJwbj/be24F9SzamTXlsXnzW+nu8vNWOxEysFZwnCOC/r4lNBvj
pDpAIUA2NKQ/acINzRwhwSGOxwEQl0ex39nzGrAgE1KcCwE/QN3pC0N9TYS7oNkq
jg+x2nJKMZWr2oznS6LkqJkmzDtVkt71toRVQVOhka0ncyWqzqNSeddxmwjz5J44
BO4p9/8a2FGEmHdfPg6KNRA7xTHyxo0PNCYNTssJayLdGGtbqqFk+K8oy/GCpl+e
GWwIrXc3oU+v0JQk8Ye+Hn3hlpx8PS2krFTzRDvAr0TgXfuYcOLQK7Lf1CI51LWk
ycT8+x2lnCxihIfvFYUeaqhQiEl70a/DBPQPJ6BD+oZb5Ufdh5YgV9LDqtFD4jW6
9qtch/0zjjdx+okU+ENayF5KK5Nu7MmyCLRYZHYIIXgzVhYHVnLoNzrjQyRjoCOo
p2Zm9m6kLwncl9FwHPrybDZPu6FV1cbRGrO0e7pIZYjgzbnPfyTltov78Sb/hzU8
N6TEb5ceRQtnb5s1ueKa2NuUfjdt60joAfkF+Swmw32GOiVnkxjzrh1rZsZEGs1m
qt6T8wiirk8P6fzlCMVL21m2sVx9VEXzAD9ejFqy8d3e3dVsuMbN2mxqNlk/9LAq
D0HcrSAa+pdTaMUhMEf+aQb3wBgCAOMcKHLPdPsVRzCyZtIfIv609c+MqKAWpzgL
8kuXfq1q/ogjHlop60vz/W2Xf9eDOgTgkU5IPQdfc8vqAI3N+HPRF4kHhsxViJG1
FgqcdOJugoUWOHdTa0wYKy3sNZC5wy2x7otjD7jMuriiAtVaEiV1ZQAN+HwJYSgN
d6QfNfrMiQlZB2vEZVUlHsqBWRymSDE1PWUmVbmNKEOFnQl4wF1tv//Gy5hwqen9
TOTqZH/3e3/X2l/MA34sbP5nol0+W/qv5T+zmdYauxLV4kpsOoMMo9db6NMHAirJ
TLzwi+1UUoefzooA1olwTfODwVLGpFhurmU4zywb3DTHOCZpSaXM0R61NPneG8FE
sAuJWdJx+uVWHCV67mVmrX8L02oEwVp/RgKZmxXs6Bei67WyRQKNY+SgeL2h+BmC
xq3OUaNKGxPVX3I9fcJevjGxPKvoCcv/HTKqnNJ5JTP3GL7uR+bF59RHxrOwZKjN
Lvq/3Sklh5XNiv466lqlfrxdUGq9pRTMNhGLZ2hf9rnbvv1S9Ypgvj8M8DCdjUFT
uL7HSJBayMqdX9yRZT5pW/8sQ7JAAS36nwB4MItZ1Ncmb4+Qm2bwt7LW7/R6Nx74
JQdyaox+wGwVJ+wkdrU2DxpSYCTgvEkoFVumqnE2GhJRBEORQUFC5o1LOA6lqRY5
Tg6X1ojU9WM3diamp+D1ggrJGYJcx9OuJ6w+FTMQvEYoymIUzyOLRecs8XrVmC4c
yTitJklY6nitKYUaoaFEjnt5WNSCojyZ84s3p2GmRqGsLK8LsH7dTbBWjNFuwBEQ
yMKGAu0cDw7W3raQ/ZGPqCAH8wFtd9ogu7D7d+ni2hjs9SCB2Ti96JprCyztmVYx
mSP8C940fldntftoQ3Rd4O01ODVFuWGnCTDt5e18LaGdWY55Ck8aaJnBDsVeu6/U
Anjz9g9eXb94foxKyywBIkToOTq/q7jZDsMbY6YetvjRdqJ2s4XnDkvGVdJpuRWf
NRXLzozcd/64KU/pt9zzpTKF/XcibBwzKmjZZYYWsjgHXk4BNRxxYF7prOxoLQSa
hVviAeYOpcpD6kIAIE2ciC22XqA5UNmoliDgn/uRlzOHu03RUqy+7LwmRNOBNHIQ
dt+o7UsGW+lGijaHqs8ew3Bbv2fK8eYoPrn3WeL/uBITszxgoNwG/wEZuh/f6yiU
RtsetPz+OH42jhWgxCAHKmSCEov7HHkEtnyZTNqhORuo7pziRAEXvyxqGtJGApvB
69dl4VE7WQOGGlBJ464Q9zmpMuCwCXXJxK49WXWwMK7HCxPG9hX3D+dKDxxofKi5
5t0qDYmdGzopiN/YgQv0/IONQRxOC2iTS1HoE30Zz5XTEmub0nVWZOPzChMfwVeS
06grOGQ+PPNW43uAEXxVgW90QtmACN+YVYf/lSLdti2RH1T/5iI3yLybyIKt9JbA
s9324GUa1X0/mtQok7DSk1LGq6uOWnI0gQA0PdYHsa+pfYM8rtl87x4HIOBRGOpH
diupy7N1OacX57+6vT1LfvTBzNCRPBb2M9XKB7xBBWFxYweolzHA/nNpeRuuWz8N
Cve9v+y+Iatiq5qs04hZ0cVRG/a+q5w2/4UacMRdiHWL8WjZW0dxVh0Ib1CAspJ6
56BnwKuaM6svzill9EnieZvfalUboL+IOa0HOGTvrUhHDFfSrY18iUPtiMpBzhVl
xOa02hkapkXI0t5ZsccDUllXCd8H/GPxsTM18olG9m/CIoCRpQvToy/Gk0FtQCA1
+SF+soWkO/JSJRREiK7diAXDTz5TCdnojJ3BkrYFK8oZCrZWJY9AAI9DrJXAgJUp
bV5J8bqAKp9Wmea7mdpZPTp80eACtIDOR0wSycYHUfXVjR1R39s9SXoK78GLA7oJ
4L6vBOC397UycqKGbP4+03d0OzeIVNPoRtbU/nrqEva577l+wuS+WTPBr4Dk9iDb
Zi3JY1RJ/Pum/259DSXJxmW93i0L/aTMdxxS5OQ79TUTrapqIICdLwtVnoCISNYy
KJkLpUQEnFoCiVmKyFNgDdfiYxEzRsW92F0bdrkCRZnIHtJuyu8sCrPspDkIlE+x
r57/jFqHW7nw4P2j5tYcHIYKga+R8wQ8Wv2vonenGzOgv3yXuTmn79mICpkIZTZd
JDmRIzNJiKk1vHhR7Qawh9xA2XrxmZ1Z1UgYfk2DATUyZz8A+mkQjCcuvyMslqZt
UnkFTbCFm6I15/krH0tTcxwect3c2lGNBfyXVjzgEX/nsI3arNg4X6scaUC4B5fk
VuhZ3gEKlIP2TAtg9718tReCYFkNlRFehutbN5/wGuVSQcQK9fU20B6ZGwt1gsgo
nzl7qXZQlSIJvc2LdE296Nkmtxr6nUuMfhkExbu68xgiQYm3oZzi0y0GDaZWlyWd
E2nkNZF2ehuxfP2/aHsqgyuQa/9c/kH4Pn4+K+TlKgmGdiYL8Ek47bWM8/8ki4sS
NoXZwXfIcLSr/qv+5uI6GcU0gpZ65siMNLjyeensi2McoJNgEdRkmvcD32e0RhUG
gtmlEINyffUXm2lMmT2c/ZJrx3vSjS3+bJ1o4Jcz6LlEn115qn8ZkBd5KfR3DcA0
P7W4GlEXKAFSTyhg7NFCl8JszqtTFf1EiM7wsonEo6O7qUr+r36ktEYLkpdZLs78
6FAuj9dcpRN297Ik7TEjh4j3oALy6TaMpbRWChKBrOgt4ZtZMbi/T1KEzsjoeBUg
ZCz5U33ne8vs8Zu0+7fO9BBZsCgpHWTLXzr3SGxxvhyWw60WyMvGSg8GjdhgBvPj
KKXq995Ke+H0NGwr0JxCRtU95yqDzxQCR4Om9TIq7QXjn72aq385KgbfBwPfrEXh
xVNvtAiQy0oW5ufIQOJ1IWMik9GBLo43qJE6u6s/JhVAa0AStw17GjGpgqI/1zek
X67rwB5suIfMpcJyYSZxZDvRgBEHrfa+RDLFZ9cXKDw2Q2YhlRPS7FrRQ7RaQ3bp
TWY7oNL9u6fB2VbJSYmW4yq/ZyxBzFgTPjs720aAKLO+jlS3Kkw4aJvgoUMGsg53
OcHRsxhJJLwaB3gVZoqPuKqwK+4+BzizSNzadP5ekP7zansmcfliprU/yIuYU3cs
xw+C1WSWwoB2eb4BIUnQhiTqRc4mS+2LtJiTvUquGksfj3mXbeUj5/P3F4ooMZ3r
NaKWELODCzO4IKOWr7furVwZka12Q55NoSgEsgHHAxWpMcXWgDOi3iuZGD2RXa+G
9hKSL7/DDzPz+/5ljau5D6461sl4sV1lofAd+E1Kotp+4MuBcfZWXlIOhqs9xf5G
z4/j/094Dn/HW9PTGCCykN5eWCDWOvE6tFgAipyyi4dKP8a6P9f3HjPr3FgTBB+/
MZw1t4ZLiOjebN17U8TShsRDjTnQtVmi5y7IxDOTfPwUwCG1IMXMZ11Jzacq3e/+
p9hQngoIWeb3f6EOYwTNddJUPC0ayev1ZhU5s3XJ0m7ld2bFvLnXjhoV0M0YpQdk
fCQm+dU8CHPprPuuzUgBSfPQxwap1ZdcNAKTt+VrGlZCHu4habf5DwUC3CiQC4N1
2+7rRYRTO7GVwRfCTJOuPK6zKoL9jW1UEVOfUV3lVHsdGzBdL5Q7VdPavJtbz/B4
C5V26IY9moL+tXwurPKDKhRhuwDiH0evLDkxCwHL4n0BEBni4Ce6ZVv+Fh/fV1nY
qr7wCNaT425lfzmHtKzVl6Nw24kjs+xX82Sip6For5wlqPPxyaFtj3MQYyDq5Cxx
PxFY/YAOTRs7QtHBpNxHJ3toRDoDDZi2T1o6cBzSCq3dcLRvT92Q+XZ9qw9gSgJJ
J9d9aALV1+rpdmw0THdIzQ8Cd9xEtdgmQWe7rJw4qo0xDof8OH9i7aIu3XR2G3d0
6ljAKc5/rrD03noDAMy8klVvgkugOOuPugir+Xkqob8sLq6dfXljZg9GJTx+5awD
LLGz9UoESo/7cGtbG2LwmIhtVV5a4Y5UGRLj1QwK475HtLO0jrKrD7LeEAATx5Bn
6R5zR/uf24aUoQBLKnFTA4xb310xD3SRxr7mxSOt/hOYmrfCbFaJJeh14L3paiTa
ehOsnmDaO/5+g8Tpmq7vKcVf/CYCBiLRJ4eXOfBVW//lP6aWW3HozAfa2auztYwm
m8O3B4sNtRmu0Y7uE+aGRjiojOTK3nLlaO7WlmrjZHAJdn/zFpVK77llqAsKvdfd
4WlJ0N3PGU+kSnM0f17GB5AdXKcMGjPJQi6eQLO7JQsDX+3K+A8kwdonz0rkpoXJ
WtLEJbS/HfHFvkOeu654uverVXUFnCNOXSc+ZpWmkZP6DUUsKt5qyGAs0/QGCrDt
J0629pTpxbuF+J2CeNyv3SapDLVIfR2eFDL0tAuiAMRa6qitWIpyF7XMtZguW4vb
pqN83Buv/bFnONVCaAUsHpoiFyxeBcZdjkEVx7upRAG/WkqCCj7D3DJAKFNGMBM6
7wz/vh38iuKPYY8R4Gssl1l/PonVtLXeM3IC4OvBxBRpQBg1bDrgIawy57FmPigj
FECCtbI28j5SWy9KCHrkUfooYn6lpSHqEdwnsp5Ej9uHdQw9IaOdwC4nFu1qHHie
qR47bnsHgMCZBxIV8KEdYc6BhB87ixUJdziwJWysvyp3o6hKU1gGoxqw/aa4AmPo
WNdD9G3V8eYeGI1EkueqYW0yJ2PhGeAMtuJUu009aO8hLem8yd36VcUQgmLJMnPP
3Qty2jqpodHCYUY++DSqEKk6z4x6so9ti/QyombpjZu8r9LCZaaQy8YFVs0FLJUA
W/7XcmJSaLT1h4lAV0zCxGJY2NTrOni6Kca9zCwhrEoabfIfmJFzILeylhck8I1F
N1JKCCNG29F3T5Ci31MkrnQLO1kDmB/G3kzzCJYXtudHsXGkRIz3wr9Wg9ARFBUN
FtBkBY4xQGuC8tJzO4YFkVU/rXu769REJUJkNoleHHhY8a6vaxWYQ7rEnF03rMUB
6pVbQ3IkMFgNaL9ATAXztP/HN+I9M/g2Hf15b0acjJIwEyFjv4goNYtTIo2Nbccf
vOkFC46QTkS7FOmGB8/lmpGOsgJ6LRVRv2/oAPPR1KTKUNoma/FrqO84YRqkvpsH
sW592bGlaC88BbNdCitdi2v4YAWnP0RPo4tQ19LR4w1GhXXlAhu8vR1chVZ6wzjx
7UrEE9rKuHAXizUfPdbjlb1ATaYmZaFJX5CllUaVFe2L/DL0PL49YmeZwZL/pKHw
WavjRJkzWhBRZCBy7RfkPj4RC6vFYFRus1VpuAz2eJCIqxK8cPTE3adUczLoGKKD
4yjP5J+SGhklPHTBv4uEvwvcZJ7/mFfiFLrunj/FVNXnuRMOj4zHEp9OgoXgFUAh
xz8yddVNbC8lMuG7EOXxF/wzFiQfSECAhdxb9hQTO8UcVjHFyOffdj9tjBBhL8Mp
CDgNsa/OYxK+YhZYKSufsT9xPWxj9woifrag6J6L8l9ussg0KKeaqIwmgRysK2Gx
C+ucoCGcZ5v/G5vx5Cqv1g6zkM5hAWuI8IuvsVW/gQ37cl/y5XOQuCLDIPzqEl+A
+hPtvIWQGfOZSfV1LIbzO9etgReuVk+IDhU/FzcT8uEuVvrwWTgwC0GTmdbZ4ABa
EmUIgOJ/feu0TQ072DBbulcwaLQLXz7YTepNFGq8TN3iZy1oF0EJO9QWd3fQ9iB0
SUBKeUa3eRWGeszFO0ujm/y+1kDBryhdfLAqHFGU/t2DraVKEIN4wEHDyZ9qtjBP
USCSwXzV5qDsfAHHJ+PDLWZ2W6weG8OeZXljOOO0iom9icJwTYhXC5duuV68c/tA
CHpqfJGoywIX3TtXoPqhgVzMvE4awQGwoBpUAevEqrfk9VZ8JkPhfGezeg084/vo
P6iI4ReRup6G2WqAMQi4ksVWyHKn6KlxKjaeVr0mrfU1ldqyL4nwDIh7Cbt3tJ0M
HDXoAksa3M8ee1+JzYZ6Xt8AXYFgl/a+deR9aQ1tZVrU4d6zrlAykcg9EoJngETe
kzQg30YVoRgu+V0d+d8JOitzuf6+BZmHhA0D/MF8zAmf3fMuIAODpG56NvPjfRzH
JHUs69zMmOIK11lVYe8uWQSxwGiC6zJMddBSIfmfvixwZGFMKYlXhPPmNQg2Puia
msxQ+SCA6GSMiP/udCs+ZdffgQoZhTD4MNts03xO0X37nQSWQgPvDAH6WZejLIXg
rBev+rg4g0ngWQwcCRBqhi5+XYhbETbv6bNzX8D97HKujbKNbVedxDXqCPupa9kA
29JHHN1Nk7agrvoIVPJeiyH0Kpm6qn7sUm9P80lw5FB7eGaWAs2CIaSmJLW63pRM
sccA23pOkeeXVi1PZqaK0JaNA3dhH+D8IRt8qZmI7rc52LN33Ov5wSdx9MauwHfR
8UROcA+T40GtJjK2+ruWbG5+PgpuJFeDXQkxWjsU7OfrHsk2+ywAtIifLiB64Kxb
b+Gf5EaK85AAI+Y+LHDN6FlqxOZOEaK8X5xM7CVi7vsrHHYUquej4LYxyB5wgXC1
mqI+ftYXTz1KBIGEF3a5LiHjBuVz+VK8+23Sw9sB7U7CS8W/+qVBv44y4wFqj6Oc
pyv/LnQ46FwSQAXyETJq67JnWAfYjGeNmA6rODVwFKxTX+5y8ykYDErFkPTrMZ63
R8UGO4QFTa8SmowHK4lBBpTnXkBj3xP7ud5BIdE/Vuo6LkgZncKRfF1lzZI912W1
KId3qpE70I/QV4ty4ry+hVpFO+PnhL8EfTZdov1FD9GJkYMneqGumBb75bRa4u2D
mPI0vT4xojuI1/rDzpNWA+SToV+wmpXYl2q86HYtKB+/kOP4eF8HkYDCoA/qZMQa
2nU6QckX6GzlZUSCbm2XF53orDM+CDtWCqpI44iT+k2FN9LD+uCI0zxnv/yjp+Zy
BVigGggPJXhLKOon/Wpfd9jpu7ITzdB8cvRrfbmTnfHLTn4aces1u31dlY/tYL4Z
rnwsrUNxjcXNCT/U5tsBD1iuj+AsKT+HB0f0Dds2EH+uu+TwVJ3mkX6BuL3E4LJi
U7uQ4heul7EKwFXJM+aqoaEF9z2DpKIfm8HOiSUcGNgDTIBKspLF9yaVVR/6k5wl
fqAgRnWBK+0Ruz8ekG0Jd61TurZ4w17+4hdxavsDlLR+8RmFfrt6nNkGALBILt8w
jHLKmL0ET4Wlgps/orcD4N1nGjDMOZZBwKCeHCkJZ6Ba0LuEFJFYLjupEJQLX3OF
Pmw1LFaO/R75V1qafUfcTzpWsCljyr5QQW1khESgg/f4k4xq8TmHUi0tclVdRZjn
n4XZ98LN28atzmUo+vn0Hj5/Cf62BWg/74dcr5omG/N62IJOhoD0t61UGE4qPFnl
TFOySbK+jFqf1NVTpyaU+c05ZmTs004LmCp8WEpkgazam9/oeA3eu9Vfoe5oLstu
4e8d/DnlUZU5H2Y8HEOkdWmIP4LVg5Ss2PWwHUsR/+iY3SbxJY8/2PF4IWXZC7UW
gOWTjG9fAcTGIFYNg/gsKpof2hz/c7YVq6XfJqonnTO8ioCKl4Gi8GgvuM32QXOb
LA4iGnTXJw/tXGwmh0CGjoXet3mT3pYsWWHsyFG0KDfPhr/A/zO1qaYc+2JnAEkM
T25s18FOwJUhj1raRbjUp+HuYsaXOlCMQ3hp4ffCBd2T2XPGWi9naF5VSAtJv6he
B/OH0gpkGO29AqS8ltC99C442MymKJUVNkBsTVZvE3zQoUrfq5k5yAGRk40INShq
WS8yQ6AKiAfDvA45SG27j0aBby/hFgv7hiqk6etunrKO9mhs1HdMBJh25xZBqWmS
tUi8nUk+Bja3nEtvAsZeUZyljMOc/nFXSeibivoLispjw/plTlgb5xK6mvE51yXu
O3BpX4U5pEr2gr+AqQs/MDfkWYSb8XvVvtzP6Y8JKKEO3U0vkzaKVbp5B2IiE5Oo
Hzmty1NWkDU5UdXNbDBrxLsZfvbdDduQxBb6MRXD1/Z9kur2i9NqqP+bDWDvJnSv
dLEW6xohXSAvN4ejbBxdmr3M9vFaJZwW9ssrS67LbwbWXS4SSf/lJCHC1A7sBDj4
8fu01Wq53vDzzEsxzoUeWqY5YKAPV5ZeTKZEJhyIFgFwHMKsYxCMKVVXYmtNVw+s
JRXthMdASA7WZAIgodJdWSUa0EXZciROKu22OvdW4hPljLe0D7/ogtJ8kmb3XdlQ
hncGXGRV6NnojfCVI5L5ogmLJ6DcEy4GossG19HoJfp6QsMzsyuo1uf2qHffOPWu
DyKmI+DjXnpU4Jvf2T2Yyz9jCEt+qG2eoHyTSnF5N6u56U/yeLA5NRbv7V9W/m2C
FjqzzrH2GMB9tGCsAPrKQ5PfUTNhPidcbX4DOg3kVqNUcdwbUYk6YHEveJIIDN/9
7FtaxjPzuOif/H5WwtnWHP3gSvpFcTwvTNtehfmAXNknHkEDEgOPxxsuQzCOmD6X
wnfNeoIyYZEcjFwNxNXSTxynLrxKmouU5iLmbnEz2i6NzmuIHZ9n9/4BT6MeXOj1
WHA6mUQbQooj6CkdD86kpof6TVhPBXJdr2cyiNPsYfSAgUbKYO+/yzsTFvQVweBl
36+pittPODZDkkp9C45zOPMp+dlNfdyZHmPOX05gwtTtQ2s5QgEeh+1T3UFYmB9e
qJs0bw/aLq7AV6mR0QBi9t7wV5IS7swQUUWu9ichJAWzFTY9+6ayY9zmK8V9CzHO
Y/Pkyabc70l9/c2vH/6UTSjFGIGqpIXrrxMTepcIQuHN+hYe50/JAMuwbCyED9Ao
rYN21DoFdy9o29WsZ0P1Mmfw1jRDcikq0AkPA+vG9iWjqum7Np2PIZZuF9oIWf8E
XZfwTOhEUgwqULcvS1zMcAFdZwDjwlIf5efNZzKe2xG0ZBbqz+EYqFQRAK8AZYTX
O2V/EDw6/sRTd0KFXSXloqUN0h1nQINVS1aYtQ8f081RlKD5j7+hjmJKVnvKen8d
gJmCksJvQ7J1SDSZ5+Qy9TvoyP1zQZFj5Kpt4u5KdUXYVr/NOBKjqDiaQT+cV6Mq
QaRua+bh/yM4yKSt9YAta5S10znbqC9jmyj+PrAwEdI62wqbBf/Vg/HuRlNKDaLS
h77z6PdRyLTiuYdGAij69dd/iKw//dXbFrmL8U+IqV0Eb6BlKISJCMn6onxbRmqN
DCs2x5BnmVgnBRPCncxxPobLXOPNXVbtW6g2i4LQcSOW7N97JWMQZlEM6cbrYsTN
ukNnrJYCSywYhorRmFy8hIsthUqj1wnJ+IuoreLKQv4tkUDCQILP+tIRuf0MGuSm
OPcxhe7+/79EnTJS8IqJuqJe28YeS87xoBBSwj6Y3LYkKhLQ9l9Gv3CCNkcMZ8OY
lhuHtRGPtQaE+yX/5P8fzA/VHOpYzL/8h0P29A8nSb8WJMx0ezAgf6qGC+tD/bBM
TYTk099G5vkQTa88ZxM+i0M4U7Aecmg+EFzLdHkRi0CvMvLHvxCJYlG1spT1IsOp
M7TZtCpHPo1u4mL2YWiyqq5w0ATERwGUid6Z2U7PQ6URF5ZHhqhHcvFk/2v7Gkg3
TUbeX15XTQuHN2sVvBJk7Cm8HNNS8vGusPqlYuK4Xvi0kDWWg6BWCPBSlT54DvrA
58+McME3zPJvtAWhp3wEtDVkLD3JtxChbNVBOJnHLn7PY15YN48LZ2xseIDMfq3J
pTzDTl+F11swlZXwgdKi74Thp9yvDlKg2kKJ+23e1Ac8Rj9t4aVuCyBn+vli6Gim
QvJoAvArrMD8qOloj2E8zKtWg6L44GA+fwK+S6gGCvPkbrfDC+2nGC4zb5b9CtQR
7BUs+D5iMkyjFmE15NTRRQyIaImQoaqOvKhSDL0VF5bBDsk451K/VwZZrAGp2X2p
tUeBdOFEkiPx3GSzUF+URCi16WRlMzhsEwn8B/WD7gyud0t3Eimup1ngl5JhFcKf
HVVIlbV8o8eTwRdSB3Yzi5SPnsn0nFq1kxunomInWg+Yl6LCZYp+Bipaesbs9EaN
GchFq7OJWacz4cyUHdJ5xHDxKJZFimEgdDjVA73iEutRXq6TfjZxiCm43bFUxr/y
reFU1ZjqtATBkywivrCrtgei/vHVuhwtCt1wBo0/sOCC1PM00qoY5miJ90NZXNhe
uh63BEEdIup/rptqyyDOaJybU15ksx7cYYo6sipeKScmU4RJFMs+ieJmzOwULMoH
680E0eCJeFElCXfEqMn9dJERHijidp3i49qJN5LRtXJKsxMOJET3BUa0MqO7hUjL
ggh1tukbeRBsIs1RQ/kuznO1MntWB0ysRqAjDQQeE7S38NAJf5V73duIgkhLiYDt
1ljHk8pE8vXf/i5uFjAXCJfWBYBdK+6mtxawu1NxoMU6aPlF2pLetgqj4HF+nTog
1vz3jx705/353Zi4PtCP7w1SBBDF7D2aFGTxGECZ6rPJTOauCwZSeK0yBEeavZL7
dXdNJMNVT6oeaB4yRXSjiAQpSzLroNCZRJerzI34u8GUjAwNWbCe2XBvQu/O1auA
EJxYZRiyMpSkqjNfA+CdLoQ7RCKH7fF3qi2vG+mVgbVgIH3RWDqjZS637hJNlmbF
nx2NUQDCv2tfoj4Sf3rTC7OpLbVa8ckELBquOYcwu6VQS772QFelop7a0nCKJCzc
zgqIlk/LFfJWizpeNZq8gWIW/l1c/q+EncYqNT+q9KitPSJ1ZX0lcpxvW4g7Yedg
EGdTKvrVT+xMvLOrQd7RDwLYFRTyQpvvDibmLHV0weHcRrKuBmMETz4CJ8SRDayL
JKUq+hthbDCl3d94wBax0OMsORNBF9JFUvrIJkI4FQ954zh64usmuIcLqiODYom7
dWvO/ygkH2choK5Ee3I31owyJIFgZaEvhZa5WfjK2BZICD5zGZfwS7NUse++0W0c
ahTg+cFEWWVZ4SsSyjajoyALqXT6qtlbgdCh4+i03uzcn6aqQme8mzcAFTT6UvhH
+Z3DuFiwGiii8z/CUBVQcn7EqVHUHiosTAPc6Olqux3oHtW+GJ/eX0VWCO6A7axh
9+Y7JGLIbDjCZPxPKJTzqRtHXbeF92PB/LuRmGz6KXPf8isOr0eK3wS/SokRA7Ac
GDJCGtYTJoBamSQlk/+0+JQhSrVNrARjshchAgegHSQlSQXB77/YREhlbeSV0j7/
WPVnV1NiJ794C25+1EzDgwL4/nK+gXPiZzQVxHMtei3CLIrAv/gMTYL/YE1A/NKV
R/jkzcO8dY5FNRzahidE3/lu+8a7C8QkTVohBfeVVOQ7OCSqWWRM0mkqMn7YLJgD
vaFCP4+AADXFK248RQqtvKl9wsnLGUUwHIaaIbLNJ5U20RPxKUGxQ8RKyZ7ajSlQ
NcWOfIJrENl7v5qN+RZptYMrSThczqU+0SF/mtjuUgKGt4i53qz8ocxI5HX1S6A1
5QO+QvI5KbPUBH0SgCDIOj0fAByrJz423ZQ+KY3tZRr4LRJXmpSoRIzaE84avFTt
IQCXzK1C9d9x06+kRWiUm2v4Wq5CKMhLxl0w/8p+tjS380MD3l6+8AirH7GhinFc
TsHEBCyWn/xiKtToJTB8JX1OFPd1X/S6T187mtGn5YlDbVwS44dwwc6q2Jg1Imfu
snxJ3SvlKCCwLWWCkVudK6x1KkLgGA8r85UJdm1MsPNWEk4G1YtEuV2D9nbsI7Co
syP7gkQxl2A6BI+YJyk9hP5jL9eMakK4bfp4d2FY1FhDQdIEjjLwprZ7PnFrqrWa
T2nDJCqEZ+epUGO72eSDiRgd2EOrbPmqYy+Mha+F5W26KvAoRixcNLnjTU5a+7/B
tDGqSqW7zYgtbhuJUv/mikRtD+rdyi+C/B+eo4qiuXPnTraLg4sZ38jepVlZOR/z
wntzuABNvNF7L8cStrOzFE3RtBMm+CMjIoPtplXGs9a7mztBcxSPN4BEbxW/96xQ
2nqQVt3+VRxLvEhp2b6dtEOw/9F1az/80dj375OxSbXvAm6+xby0pW8XkjXOnBVk
LcLx4GVsiYoz2kb2uCegNM37O1jklvlC1PIkVFrHa/TYdqUNmLUY7Vw2fh4Fjyrx
a2M8Y5yEzZRdDYcFX7POw6rK8+CQ78HQK0ueoFouUYi+e24rEGMbTp/HsH+WPqcP
ELljL+XhLvbDZyUP6af2b3x4Lo/oSj/5dpvmkZnkJkdvACYn51CM5qyUXYMDxzFu
2h5mqW4kbu6SOERC+ss4dFxzX6ranu7UfxB7LnxftSVtrtycFx5r/nLtM/ST1TjL
PXzRFWrHKIbWADIGdrgGN6dOuKJeuxeL9MfAMWDnUcCIZ09NF3HfgWStQZ4DfMwg
Fl8ayabtqiBSdrI1yp1CT679w8syL1KDwj3jdK9Gp+YaFqkGPkQEKP7vaDJ6BspU
r4VJP8BOTd5Mnssk75Ip/LrfERi6j3/zRH+fWyltLQzTbthtMxcWtATSt64vYvt3
hp6N+CbJGd0nP2DqF3xllihSOcDXtuGWeirssbp5fcN0q7Ex++yRfSowvxim3C5t
daKE+7XlCo2qgDsiHcO9xB6eq5KkNYbtyltleSwr7SVcxWtS4XkOfy69OriZjYaD
eN2zmaZzqMyWGbjGv8JDe42ezoE4XaERo4gfVPv23oa7QZ6yCNZKFqoNGCbocXS/
C2+uj1cX8dPUciv+N4JYTqCl6pcKLPFgRi1MIhH4hnIfpsO4dH5OI4SMlxVcmJah
joRxllU430C4rZUTLLUGBRkHEEG4yXit/S3an1vmDrNmy1sjeBagn96aYuUR2Id0
qIS9742besFNcVXpC/VvRCPxGwnjVBGUVi4ArPviKrmxVBOsGf3gH2VFV0twke7x
pAl2JueV/laXSAsB5yyh2MCFiYbx6CwEJ4nrqayfjiY1SJhyQaWqHxdibFaPBL2t
GUj9YrMtcjFuQjZNFCZYlLipc6hBk1SNZkCqTkc149vmkhmZ0xrVQIoQG0OV1COX
w4mUVieDUUcAVpCko9HtBMqHDFymcCfpDDsRJeBBSMdXdkZLOCb8wOU9n3v7zhB5
FeMKHIit2aaoVZe5Zgouw3un2d738tXlBbtqZVzkyVrPsnpvKxz6fnk5wbl2XCSu
KIP4NENS2g3CiaPpaaZlTKXhl/gwZU775wKpMauB1KbaX6NlkgsYAEDCVkwaDLaR
Lzgr6E7Je+Gquo6FdRImH2WnuyuEN7bIC0eTMDAPt3Z0NCmvpRLAzHfG5WmJVHd+
MVbOfaHuFYKJOXqDrAg29FviFtOLb/avyLyoDIMOHznGoCegrlaLkLtvUehnp7yl
Tf18BW1sTauw/y/mNDhV3fkwwYFPGZ9p+xFSQl2iKO8MPCLusC2jOUtGjzmqDDEq
Y6rQOzL2AI03Dh/qfOaxeqVh5s10KR8FbA+xYz172tzI1soKUyLTMoDw7LEYtjGc
zYnDAHl6d481XvrTaBfJHFixQ2i3GhoxZdAdOfJ4IUIoMx0f6HSpD71AJKHCnJuB
+jadhSa9n7Rf02WSjVaGhGV/8UTbELJFuYtSnLaxr1Cb0gCHJrW/A7req0jUkeCe
F1eFTCoEcWLosL/6x8XrcyOQ/2Lwut7FmOScHrUkxgAdWVfu1u9+QEPbmTk2TS+Y
2qwr/+d2OWoC6AM+u7qsiGGu2tGTvGfFRxk7qw48ezmheeRy6x13UlnHjdpWHcLc
sNG2JVnshfNltpXMlMqdVpXKKk8N69rnRWO5Cha8FYgXpk/LlQSJS3qp/9+E6JQm
AasduZTI7ntATubJFhM+54nhk5yFSpHMLrgHdWQvNww4FKMbG1KVIOXupF0ZBIgA
M3vjHbRshn/te7i0i1s5g4FA21nMNJK9YaNJG8+wBLhxJJncedyiuDX7tOzuXLk+
xp+HrfBQTvCEqv6Zd4KOtYjJ4PgaK7Q+usp9o651TrN5lN5jlVjdcIZpiaCffk6m
xObTufI32q/Tvca0fYYndu9cZ0EYMOqz26rx7lsMmS2wxO1DsYwZ5PlnxgoVCdL6
Sfh5gG0cNEy9xnzMi0J04rQFdr7GWxzwecLM5Z88Dl/eKqJx67huDF90GOsRf4eC
xq57wj4+6aDh7Woea1MzRRNXoXmnFl9kNuizN7+mMs8rkWQVfUd98pYMqYi+nxgH
5F2JU+8Vi/DJgTv6PMIry7DJ33BaoUW+wtBvByxqv5H/BwPbfx/h2IIpqD+2l7wA
2qxFHgU8MiHuqZ37WOaqWZR7B2KYq5MJXBTTTLoQ1LFHux6jshMmCvSqlTXNcLhg
kMVSaG/xfaOv6oSt8+9j0zzMGd9tSy9ejbNrLu9SOzldtJaikan/ZKRqAhNHTTFp
gLPyBCqoIaMPLGCutSJp7Mj2wYmjT2iTYLsTRFU+DfGy30VNF8s+iBFxnyvJutXF
kdOqlwFnpegbzlNXqFvAUZYWhFUhtaTXzIvVUXOsdtq9ZD5iopUtAD2UY5bdWEau
O7AtI5TF9U08dqVYmVl8WIY5jZ2DLTnhIyXz9e8Snll3IGzRY3aqQ1YpgIsSB2c7
5cl/t7cr9780XYkUz3XpbTV+/uMOmGLtkmmQgiNUTMs7G7mFqh8dX9O//i1wbcz8
Ea1ALeollzlHLWbLAtRhnHNJyac9NkRX2QHhRJQBQcCLpiTLHCL3Of++bqYAXXKR
mL8dwQmdZZNp4RTXfGlFG5uJATMmbESBH9vV3wMsLJPlkDC/fuQK+sKhpBm2zDBk
KxEFItxHtuhGttiRSzC6GrGOHv9vwqavIeaaAc8b3sEPqCBbKwNxGRU7eoD1qjZ1
LSCC3Y8U2dw4NH/V5Rd1PA89idFWmREZt3JPcF8/dG79vb6M/C/dp2EjFGySaTaZ
jzpO4P8OGbXg+vlbv0oEHPJ347WRO0pNhEv+fx7zYKkMnax1aBoJgrdIRmIgAtaw
sujpXXx61umbFSWuk5YSE2NLE2cdiJ/gDhDda47qUbAXlKSzJxYaLyjtyjwag+N5
LpUMh9Bp6lkFi2QXTeYLFu+aPReXWtU6vWS1x6uI+B/mv6ywz04Z4/kd+AJUPt36
5jwItOSdRWdCwN/yZ0bTj4xNxZ0M92rK2NkERg0ir4L1a5lgiznSTxIEbxCsqrv5
pPT5JhzqN5HC3W8blzMt/IgNlU/Moc2uIaEl4omAHclojuZ1rQOT6TEcqC5Ef7r6
LqEXKTn7+OyNw3nOHofbYdXnAE+71FMWkCa7750iI+gw/XCFwbRsy0z45zpEgkZ7
2X6gaIkKxmWpINeMiSF3JHysocF67VbzST/qhg05SDSXJ1iBh/2QKnMM8mwBDkN5
VErJbu7ioHpAEQ0bJ+4FqpN7NOfFx9u1w4SWjFz3O9FhwnEi0piSNhVBggJlLTYP
U/lIypRoZVZ5oVcw9bSrwbSw7aXrnBA2BP8BxsSA9SqzaNG4xRhnfK/TgOcloPjN
D1FGn2ugdiMz+dwnfg7c364HoSten6rg42vUkNc+Q/dXWpZTM1YuIr+YFjOwuLFq
+s+lTHpl2gpL1uU/9xQpT2T9iNrh3oRy8NbYZaxXZ8g8Q/kUc8izrststiF7sgSk
UxQMYmIMTLj2tt/gO3xPLo17kTLkI5K0psKVNQ6E6GA/IW3X0uWo5pEehBcEfDcE
ARLqXF+xfKRr+z80smBWMXVBkzYOeEkleBh+Ledq/+FpMws+PJ57/jVpswiimQPx
Rm+ctQVLTLFNoJxCaWovqbP8cDTn22Y4S+sD0bWre/BmhdKRcXmmdDucy/tNxyNP
kvSu9FXukXZIQCpuF/fQqWd9uXDmqu4gXDQpCfp7fRk4+/ENpOO6W2ilHdh6EdH9
UrIs/oYyFjtnNg4eQwy5r/3sgZeARxgzXhrcgyM3rfE9zRaJxGzNsd7MWU+eS/5i
cJrG+qjfYlJVemOXCDapKcGIL0Rac2w6INDjul53CXLGuG42lEU+VF7XiutcNqbf
BaLe6h5vypE3FRHldWe8DuXLSjTbqbJMhSYizpLZCrQMFI9/7TIqUjX/ldhRWV+U
jua6A6hq79uTpCH2T5xWnrNyehI7wH75Ik0t5ObBTqFxLVpiQaDweknXyJBuIbXq
fRtm9ZVGZC2lhxCXHK2KZrbMyu/V0azOqBvNVWBOxDN72oCaCa9YrrZ/qn6qebzE
Sx/71Tb1YCiuBZwMtSJhFQfks5N5M7PddnZEnQIsvcim/HkfVg4S/DK8wRoYEn8r
g+dZsWec75489vd8yQsxynRQj+8RjRqEopJG8mrAg6FZJyRaEridrxo6acRcmQ4+
b8ySsQj4XrdBiL+PdSuNYfx6qiGi4VZ9nBGuBXW6QpbfA3iGaGqnjkNngXoTKbOH
67noHuV6A6AQ6nM4UU5QRRLbLGuPmXKttv1KCMT5zh9oHBjNBJtdQ5nr8quOcqPF
e/Bk5z8yHDwi47SFsjR3b+YYtWob0lU61FsB+qnPvElxy5gWsCTXNvBDytFnVsDH
jNYhyaqvXbOzEmOVoSMzgLLQXW0AFV+TrfKT8i2Qu5muOV7OymG0sf2L7zy/IUrH
KlIyyMkcin3MNJ7JP4x/pFpu3L4ZKVZHAyqq3NoemE30ozc7GXd89Lt9MeBFvzPl
7j803cVbYzArqB3qF98TMpPSaHLc52lU1mGE1kzmMIemVLioJI4zDfES2hNZzwEr
lVHqpwg59GoygGXO1QFraIWZ7ix/Iszw8lov3+FiERJ6/EkUr/ma21xiDPO7qNzJ
8CWQuCt8F6BcRL3wm1GYmIHXMyA1OtFf+j6a/tchOsWZ30a6hGCSilIy3hRkhkSw
sa6ptKPmGLFVR2b6IdqHDbtBqCekua6ZQzLLg9b9xWoCyiW2rJD19jxD7coq4wAw
hij2FkrEtQWSF2qoa/jAdc8R85t9fGSh+gUze/6vPMyUwO7jn8eSFSZU0MZ9joGg
YPz7hp7ov4nG1eJQi0i4NIti+KTdQwO3tCohVEnCXr6cROOs6hGRO4KoYynR9bNe
auC3wzdhxTq9EO/JWeV82q2Nl25YGlaH43iC3mziJZEO8zM8Goci/XqPD7+75yhc
W7w5GsDD8hJy+Zz6aYLQX7QWItVJmdlS5ZxvXFb+b1qkC/yyYFxMluRnBdxLKXtO
+pYJvqsuijSwO7wE34OqMOZSiFQpGLbRrhIGE6rfVo4dkoiSIr8sX0uOnbHJp/A7
Iie5sOG9zR1r3fWBp20vL/D6/G052jl7vQjl8jlbiORQQp3Mb4xNYLO+mescBz4B
Z0rjy7TZV504dRb3zYEOainFeFKSfMC3/qpruqEej7JQfg7sBxZFSl8Eg2cHGJp5
X760larMs6dzDfGqWA85HckA3UaABq3lfRFFoqIxo6EdxHhD3W/F+I7O1v+IRmkJ
CaI+tiBhl9rHvzOIM/nmhyqCXM1v1a0aU0uHPkF4nw0OkcWGwAsoluF7HRtjfgSn
6bj4fdaLEkLtDVUVIwWDIFlG6isu/j5mR2pvdIvnFD14eTT9TYfZWQmc+M12ETcM
wmXZGdv6gS1fWjegs60/mjqL5UASMLtWEWYqGTtL8GwtTnMP6ISbX1nsDMLGC5BH
/j1a87C/DOu/0DVz1uzPiSS1iNHKUwNIJ1RpDW+pUkn8FEhPC0CG1B7kimlCcOf6
BtbNuQAOkX+4Wzc53AuBYBR+qZskdJ+2vz/mUqOYWp05iJpeXDuPihirT1rcIL3P
pL+qvSeMWV42ENUy8JctGCMUtBTva7V2i0gxGQtn9f9H+GxYm1XKmZs6WRsTUF/4
2p9fhwbHDui4Kw7u3KvWbOhI+C7AmarC5FRgqULXZwsJ3IHxLk2sQ6ycgzEp53RY
xBB/TnNglMZtilSJgBdbenip0IRHZZQjXIHI+2t/kiIX7rgTjErTgbpyYb2nR3Wj
67rPZfwfnPA5+zAyZ2N901q7YqpCi4JqDWLDV0CiRGduOLmJIXZgiATfIV1wEO+W
KfkJqHWpgJE9RYSQFEYy5TrAwQ5kGDdl5ULDdAyy+zVx5n2itUVL0ycgxedhU2Wq
XNnvkbro4qijFoFpYrd1PUO6PSSD7UuXmZm8K3tMv9QvHLQ8nWvI9i6bSZrr4iiD
s8iA9p8ExUN82WCm01vaov6DPniDx92CXmGn9+cYlgKCnqPWiXrwaSw3wfvB5NI1
yTqItDt7AfitW8RSbdyUkWR3w5rMrxxzC07PmdLEus7+vRqlCUkGPRFbrszd9wV8
9rVljOBND2AZrnYSdxGZsGwoPKxJZzJl8Tr0Ec7kKKGakBLA778QQqQJvi9Qfqp6
eww3su/8VC3LENWWT38181Fb7IyTUsRWWkPSyiXNUlwsFJ4DM7Ws0XK1UrQyZNRW
mFHi0P0zO7e+lj74ijYuyTQ1MkzYttlUeyHKAfhqhjnrhvDSSgByHenEfK5UU+x9
ySsGuSu/ssrIXGdIluYS+dJfLAl8B+h1lRq8merztwmWQ3KmPpCMDrbZ/uXX1nxN
/axbexGRW1HTOVonuiRFW9EmlBkF80CP4efE7JDMhux0iwuT5l69Crpyt+SWaWRV
evJEI+cG+HuTV9/d04DjRQRps1CSao/X/p+/Q/tPDt8Gte4lKkEec/SSBiBY/3NS
GSBpVnxUomd6e7P8quxitZrI67fxUa1Ao5EyAxjTRCZLkfTX7EU7X3RSbdennKRD
FZPEiW3tGnKHVSWC6A+qCEIqwu+4MiJlrS9RLHERK/RkyVCGv7YVHj0h1Txv97d/
rGXiJqTO4KMPCUTQ9M5TyTSfPbw2m75TvQuQ7XFuNaYQRTVdHVr17HdgLkYafFDw
XOPA1qcFWuhUmVGGTit+j76rhYN8q2sC2j5ppH0srujAqlulre2a6ZGVPpEbtSqD
ucNd0PB8WWxuJd8sXuFaVO7Zj+aUCy8AIz9jH6AEy0rnz3fRtCUwoph+D6oQtBW+
ULf2jHufl4AO+lMSyFJ66Vxt8F01ov6VTR/4yUz3qiCG+RoC6NU+CqbN6OQ+5SUN
TqlNLVNmXve1hOxJDIOZFWKLTFSSDhqYuM7gjpwVdBZAtPyE7ellcAJ7iuTdpjQv
KlCRPs8SwSAz7RZ03eE/58WqXy8L7IMEDYF15/M2jkV0bxEb7eDtcPj1/NP7aHW+
J8Gv0OOc91MZbaM5dZEAc0Eq3IHzNaWqbNAgrVF0JSaUTNNjpveUOxISUpQGyX08
dmII7YahBBjAYGJw/iJO97rHZHbGq+pktlCSIPsrZSfWSSmQGoYPdXN4NQgtkZx6
5a490WlbkNStzYIpHX7tFwT1SWwUVCSRfcrLkQEwi9mryLhWUZBFK0iAe7x6dQxa
jfetCwo/ixqMlr2dOXo2c/Hj4ys8Uko3wH0MZUtu9TrEjwwFQR3GqbVqZDsab64f
qGsVBbLUKpIJf3urQ7dTbXL8MoZtosvshMjBJGMA907+eecuY6hgdckfYTLBWJ6w
9HzlpK/fy6fMunNplo4aTycgulfKxRV465J0lcKGRNcWl7NMX7YTN5tYlbFzTZNr
+veEqfeXMuJaP1PJPtz3qZGS5d9DCLGULumcggNaPzvBP0UD88L4devLjtLtt5B/
StCMJ0KimJ9mIZCjyRCW5/JrxorVoQTWw4/Qb1y5lRVwwJR2CoYjxFviZruDKKnO
kZ8TFAnsNWK5adgju1V2hiQfqWiOTunkbNFeoPdBBQCjfZlP1Q/DmiWRnjpje2W/
Rt6MicQE2R+q9Wi1j9fmeaHQthbxGQJcJ1uffLAWVi6DsK5RGz+THjuUvo+FdHTN
jYqQYfbGDMewl3qmXv92+MVV71/vfn29V+t8va00AC7rmhehyjVvtRTuhlRWdJLY
CzZPqrvQdUY1VualyYZNUT4lRHfB5elgmi4jWMHLDfUPIZtrhnpOPakufI3nJ+tf
0s/2q3+nPZo50prB89tbgDb3VPPIDlKkGBriCLOsxVm7/5kqVJ9WHeAdK6l4aVpA
2ZXkojfaCVRIqYIYNW81DZ7RPDqABERfv1CXrhVFFClCRRvecCkfAl3A9x1WRueG
OFgerNJPSfh1lnVtJzPWYyyIwDvVP8xLfjZTqVMqAgj2t62UKez4gexF6k0je3cA
kM3jP/Adwbe/sxqsAsC+i7fhNsZdiVKzhujRVpmnne3Ws+3lCtCzyjM5CA6KMvQf
pqdf9zzI5h2rpmQsnssoN/8yLIE+3No42r0pXv5gsFbQJjrH3c36bIp9DNzObU7N
Thxh6IrWr/RjLT9PAmjO64SuWXc1gP2E65i/Z28+kos4ZlEveDvtzKIfJ9NoQYiF
VA840CjAlm1oS77oT3NsvjNQRrKYgfZ5G6YCuQRmHt1Jh1Tf4MvjVzhoJtNsrvPb
tUzG/vK6PEHDfkwZs6uJMz+7xtak9vCtezXKpc02dxEMsG4A3/HXG5eY82SDFoEQ
aY4NSu7SvRAVQM0QZryHIv27ZNgE/oGzsP8rJmdZNUqtMKHEDRUt2qeI+30H+b9P
tfGPi6TVdHD8VVlEsQ6YNyELdnUlbQHrNDEZOhhYLvXJCIxBAlJHJmtHqKj12/1M
4D7Hfr5CkFsp/hDRZBQPQMGtgRj74/bCLMIIVMWwi5MmJC+64ypKLeVAv8TOy0p+
9TypFZgEX2TtejLb9yHfsA6eC6lOZ8cTezqfFtg7PV99VnESulk1hTgg1cE9J0ci
aizCRevOC6uTRq7BXS429qtR0SIYUgiTBkbWiKwMkRZ0DNVOIsk2eV5hKbeL925R
hefOKggvs8wz5LfixB9YF7dKEP55oX4GNbT5PEaSOaZ5KFl0V4AeiE/IBediuXXj
NCDX1MQPpo/89I6HafhpM5D5+dkveqcr6zCNJDPwsFr5pujoCdKOW+m6TLntlVlY
M5nQztYS/nv++OddluXmQvyB9AeNZtVmjr2VVQkEz/fR/V6+Vk+GKH+S5KXs8Nrd
MUyy/ubEa2WDZKfe7DMGAr8dYpWvJWyEEmr9pEbLDYg+TX8djJgaXXbtvZ53nncd
AltkJY+GGzuWtv0eG60sTCO0VDFSTesYOMFw7wHlaO4scEBA+GLilZiW9mQG187s
Px/SZaY3RXzpAEFhkRESX5ak1Sg3ua7gXqYMBHxZYgVRdd4KW0FVUwvpmBSAl0s6
IkEKPmS1FcOtjzNl0tfvOwcj+2Ftnj7jt20ySFPTRnnqGQhQuf5oOBdAKgJ9D8Qe
T8NOQggs1qQF91/oI2YAFCTuENfZTw9DsCQpuppC1F48R3faTXO5hqObE7C4166W
hwz+TX1uUS2SEfXnzx0Qdu3OVeOj1tUE7vqVlx3mMxAC2UUEiTwHPmtycgB/gOq6
vL0l6I2qNEC3/ENHz/Qs3NYHSwTr/z7mF+n+yCSGrRk53zvMG0NNVSfufslmg57l
FfJszJHrNMoEH0l/nMUxOzUH4wS2fYbwBnysxd+6CMEBi837l7KoLNEbjevdkTA+
J7/YBR5A0mQIUSWRE59C18YSpx6UciAHZu/wzwTfNOBHEYLfcu4EBD14eE83trVv
x47k+DtyollUtuBgQiPUYGjT96MmIZc699GjPVVryNOZcsXl8XOaWpY4jWSdnpaj
t7f22+uytS/oY6i0AvoZnphlQtmgXtyodQukvYS8nd1BUlCnv4a796AOaQRnvCMr
4w7PBYug8GFfqzsTUDQYzq/GtYUmRVtwNVh7QtgUGHbO6Q9ODH/LS7Cm+s5rI11L
fWkK1JPOlkW7v9QEDNBgZ/p9d6Lsu5MgjKQI3IeaNxCfvIufH+SDqB90P4KkZRVP
4KAPhMF+6SLP/yML4jmKPYjZC6Y4FXmFd30uowTLL0cZUs/Gwhm13elWgGc+JOJl
ifwh2zMtMZvtdLDs4mejjmw7YO5yUhbcZu9LA4rRssJon8iPMjUNRGRlvY9+0Bzu
V9W+a3KusPDEtAeq/mZ5frG+JZkPtqoshMc0cxJ1jw0EIQRbsQ1eOfjoLeOhNOkV
laWXoDwLycRbJubSLC3gSji72na89PhP8KLgQOdYPb/WZPxKsljMxG/MeAhTeGle
pa6zNZkRdaj8iI+4mqDmNqEy2RT8neBV64Z/xdoxdnQVaFeiifnPE8E5kBopFtdO
DJNaU2B5lb5GB7lgrqjPkUmR+SrPHD12tF+nuCftxedHu5uU0onjm+5KhzW0RzLm
NBv12sXnYrTkAO5uh0QdodsKzmrB+P7ZamZIPbL3J7fK2jYueq5/TETtpK/MF4Ic
ZpMXWnOmHA097nn2hjlyvolFMW3bVWpiznJJP7/2NCqllQOgwjLq1ih9OC4YgZO8
vSDX9Heo3JaT2NHPp/Dw/ec1l0sUY3ZNwDpWe7Ca0lit2azPscxvM6J1h9vk8Sq8
f/a+OwMx5WjFN462IAV+9dCe2ZgdmQQUmlD0FIgi7HQcIrYZvGNK7gV3uuPMDnHk
TYLrzjjvlLz1qTZIrJ9vDwceU4zNNExci0tQBnBtZno2qkwUIsI/k7tc+CQjDhBB
p3EZHIUk8YGeCUKZBNXUeEz6rKQStohRpGMG4P/GhNx9n2PAOhZN3m8nlLPaAKfO
H7d39o4IS6e+2fXn8iaYrCBt0Z6WRGEFJoKuqK5xXgHceRCpvcxx46HVHhCaFK0O
+t0or0XuqL18MI+louIzuVHJL1yTXOc5nkxoXgF1HoRVaIdSIV1Y7ieH1YfibMn3
Hqw+yCpm2Z/LK9lMcgTT/ygWZAY7DTQEpKRnDBC+rz9TOwwYUVziuBGR47Wd0piY
wJbtDoyJhaVh8CWzZxaKvVcTspLMTJSpWbVZck5qxVmcRQq412znrqCUn8PE4wn6
NrHG04U+NQDJi8PfjBOmm68ttnJktFlozJpJJxmQnPNZ7F25lMPx2imLP/qoS6AJ
IIiWlEQQrzOrQwCUayB5KVmGLQZ/r3cHRQkcMAVhF4RCFNjiQ5h9nneJAcy6e082
eKEs65lqCqVaOjFmtLWoFD7zAsMf8zrAEZggWwy7nhSyhANCZRAELvkuSNrFeTp/
OWbJ3J7/S+ZT3U3CjTJ80zneygn9JtaIuwDhDH+k9g8zPC+OrMhGHGmx1k2w85MV
gRSDZ0mgAIU5dYkn2zQs4YSBT2rtal3S3MiQr1HlAAmEDiUmk+acRJiQY6r74+xC
jp+NXwa1pEkJ/n6XsgmqOIF2Q+p33v359UXKGBCc0vnykglj5lI6RGgy/4PMkQhk
MpdltLxeeew8G09ybSDAyo4DXikpAJpMR9lxzpGjmf7qQ8TFZRwfpt8No19KMXjO
QiWr6r78hvqLGqV+KucgSn1IcrGRWaah+Bctp1Ic/L0UCJiTQHFWndKYVbcqGb+f
mU3slpuI/+4tyGnURWBcGxlXrx69s3rIjzaS59sjrly6jSQPWgqSCILWyEgFi6O0
Sg165P+XvGUfeiESu4+B58By6UG06p6tIzcXGS96k+vao8IB8+1L9hgEJUR2YRNX
h/DdrBmgXGT8lBsDXLDGpckjnEW2oHUiQu3xDKynT2MpLzzmXKfRVxcIbAUjy/a/
3b9fZ23/UTs+GEynQHHCfGm79W8f3ZfpM4vcaJH4rEgzde6ngmJAAZsLl+0GNttp
8wG3KNDUBksaaqdlDQybVQTzYFMjS3AuF5FTQdnh1SoNIJOXN9PgHqZPIOPm0r8e
EEmFkwCY7mXdCQYgMsAefFGUouQe6dQ9B6ShVCqPtE4oJ4hMCx078Ga8ORhQjLAA
My8BO/eildXzSSNPhlr6qyhZsrqheHW6kPTpQd128GIsGFegYBQzrH+afi4fs/U5
HXlX71gpebh1MmCLc3VbHZEf7doLI8OSxvmT/kg4NCLFzaAkFrKuK/+gIWotky8W
FEansQ1RHxodnAN2zQVZTKEDyf6pMIqe81gwyDj96ZH0TVnAGK+DS6QmhUSerywB
xeexAZDCm6UVoSqkKqJy+fvSC3xq4f4rsMhfCEe/heaO6rskZVmmp4s/pZwO5H2x
NEZ8YRh2ZXv0h1Ff1D1Eb6nYyLpOpv0wzD8wwl3gTv8N/zN5aA6GZW40++2J0Gyn
sZ93qjFETZ6kXRD9Xdih8KjL9RCAwfpZnZVEY9crWwFUGma8Wu9sa3F7OvP9BH26
JABGQ3XPNjS9uB7XEu2/AVFFSgkB5q/vl/fZCBOpnL7L2pavOwJ6KmXuhDpkz/Fe
H4Vk7LeRY94LND5pzM2njHRZanU7bf+4XycKAfmwtPyW+yp80ddfPa5k26jpv/MG
yQDwlSHm1LY0ynNAiHn2o+cSfHbHpnmv266QJ8VfLxNncTN6cs7LzQDTl1KDGnWT
INSOazF/iuhWCyjhKR6dQfjKh+FTLSt1Ncs6sjCKW32AaG4TzUUNfPExBsOlNab5
BMFo261bNc524nbrEugefvJsAVLPUgmjSZMfMP2JsKqIdGXrsNX3aA3BET8/JK+m
SzcyCGI1CQojPy0Hlz7SyqZ9Q6bT0wPml7AXlJPv/6iKTW1Touc2lcwRV6bEAGia
fcLfnhrhO3YMmP6vvuJBR+pkSwUrE5q6nHxBC/S3xS1yie98+EA+O0CoqX02UzL4
eexxHrB5M2bb8o7s/VtnkHsegyEnI8gKxk6JJkuxaMuoTHPpVkjE+cMDq9RGdA/b
XhL4IzecshkMMwf+TH/CeuuGQxAdDh3v9UxEQEXQGvE3jbXH9T8u0WI44LWnTtvR
UOR0InSWFvDnThOiHxGj89pOB6eiJsdWpGyB924izbRa4pn0mrYcVnzz8hssNK4K
63JlmgjHCqcevf9hWlXGs/bXxrq4BYukAXMqmjE4n08AvJ+3BdhWttCd8wcRTXFq
gZd0goLyrhiB9k928YM/wyFQcEs0EHyLZq2OSPE9YbDeNnzI0Oa3lZthgDL5YG8S
yYB5Wi2cpWHzUircEkQPJeQS/k27Oa4WNMFNADN0gdD+kDD0LoW9DIaW+EqXYsZA
7g09g84i2GjS+z1zJTlcoXrm81aUNxWOU2TlRagAaQ3x0CXofeDGg/l1GHkCdT7M
RxKIBj+fl1auklvxDDQZORCkkME65WDwgFWkQW18YoSN0okrEDoYADjQuWAOeU2q
0IPU7JJqTPJR30VmhBCWYEZ489IZaL0lsTwRwuhql3OLpaBXk8EFB+oW3HcR80A8
+N5AzDWEkN2vSs0Y8p7MRrnd3saycVJqA/sns4uqcjPr7Z2BtjlsZjiHzcyYluQW
Z1yqGomSmNRf90j0sJgg5b0FQ4eAXbe4Msc3JiCedseRg02dyKfrINnlD9at7ADa
tRYlVTuTXZwwVAI4ukBAPjKwI1ScOMWvwrzImt2bCm8k/xS7fVIOuS+SkgTRgvmW
jgLZ42fnge7YLHfwUvfGuaIqfk0ugR7pVR9YBtBR2bP0rbli/lz+B+GaXfEMcMJF
YnidMaJWSASy+M1KKuoWaPjfRrgpxO5f0VYVxjfLl6C0vT7ZkNWEDQRRn2f3nAjN
hnDuOrkBs1Y+DH9kbPPbYkGHSMrWrDAXqcj6x6cqtOIxpsdwFrCIX5XL9bQSeMpt
FMKHic6kHaw3OW/SN7Jwq1GHZMZPGMvEAJLNVEeWsmGo+MJviKVaGZBX7guxeGR3
SAn3P3fevyv3K/adwLPy7QNM2J+e66cUJ4NGN+rPTG/Jl+krcI8ynZNG9x7Onp6C
+Mjr03tvrB0eZqgo3BElSGP8Vl4yyjZ5puKmdyvAhPFJYjo3TgJAGtA0DlLcwO2R
FwsZGNdyQucfqAr0Hx74aNyaLimwTUY7s3P5+7+CoK48cdPYIvoYdXRHiveXByN0
EBynBgqGek056Qj9OPHR/hDvEzGtmIfjvBgcShYFVLCCHKBQS5JyWqTpKe7R5JPi
eTyIvTu8dHN71OPEvxkHWoBaDvgAnJXAJ8/GjAhE3noa7NW/5P46+lbO3ko1a9eh
g1BAOEEK/a5hlX/3jrm10rOkUUKDi/QcUJofwCRiDeG/17JHjVQftdKsd6O0oHml
4xUH3cTcKkZq7WRXesE9Brl0eLY52hBmF/KohrNFkLy6kAVaFEShuLPhAv8zoIfs
8icYX9cwlNq3Fej2K7LDyGXmjKQTRamzQ5vKgyFjBScwP3uoTWc6NG+EbhlmqagV
PcFIFHmG5YbE+ehzhE+tmh7HejwQknlr1x1lBSwZKqksq6CPWksXiKloXf0itm5v
ybMxnJsWkHQMgMDET46ClQFWJ3ZX+dpqo25UpPgLLUbb42iCFt4gvOhtdRF6zi4u
wspn8zw5GMn7luW8HT/TVutth3ThONyfoGsGT5Wae+wh5hLw9frMwKvw2eFYmS6w
qyyn8RkdFiIHRVw3Xl0OYqMOrnpnxk1X+uS/k/L/ke74qYfDMLBvgM2Kvr54KmaK
8Dw6a0pSG1x+FOAV5z3h9PbHl5AA3D7EWeB5v3w+TX9QAV+fX1RVkQ4+aOn8Eb0H
7GL57CpW+tcKi9Pudlwxxr5MShcCnMCwg3QfDElrq+P0KQklDiA1cNXakmau7MCn
duYc5Ok3BC4vB3cbyLdlF2MagLfJJL96/LhlBzx5U9HDHMR4jW7+pp7z9sYIxymH
QkflcRFLV9YeF2gLdzSk4LScUePBgVaFYxMUMSBBOxaYOV+YAQAhpvTPogxIProA
lo8z1urBR6VHkWesPBng/WI4QQGy+JmiBSgYW5GF6J40Nb5Ega0d0m9HnPiXslWh
NZ/ZZjzaqeXeYNJwX8SVk3FUp8eKvkW5OSu/49rbJACVSwp5/Pq2Sm3X7z7BI0V5
TD1zBm0g3dUwBzAw/hN+vnzfwhAVBu7AwgqMXxntrwSVY/a5qjO/MuXdOL3/AHb3
fDYP1fyGW4QUWByh9arPXI+1KFcFGkC8SPUQqlyDQPR+YYez+8AXAFCqurkyVo2g
8hZjH4zN6ti8uIvVEpKAuGs1Oj4eD1wFLnuG6uWSqV5AWzyva3IkYlBQ2lDi0TlO
0y6Q8HkxKi9EuKd6HbiyXs9IzeZF24jtHbGSqbeM/Jh3rmcEoaqdESA/zmnsCxdz
xjq8TXyhVIIWOtEvc9dbWFd50SvAGHiS742IDCXX7Gk6zaX8p7f5BpMjKCLcDCgE
eG1mPtd25InCKpRIsmhE7fycDLav1PvTJqRGMEsYcfGwEl8bsWtT3AAHL95i+TNL
7PAtL5XoZNhbYdMxY9LbTU511r9sNKQd5sATz0Krh7cTCHPEXUI4Nvc3nycJP8e3
EnGgFJY3P2cjcPntgotZJ2h8nX1ZCn32+uqAgtGfGy0pjc+XqAQZbVnmKlb0QY9+
iK3MdVnu3lCxzrDJAMZlBrOWHu4PitXNzqInM1kE+IQtcNOV2c1jCVxpFV/8VGcp
czAO4hg4ESwWkEUSlmwticENVH5IZrIR2JxdixrU4KEDr3Xt+wqcBlb0rsvh11jH
TKXbbHOKt0DBZ3F8OOQiSwQ1swEhUEx9/SisYKKqQCcaXBJouq3y0KIclbVvHh4N
EY7CIpnzagK7RrgUDIoylOsmOvtmn8w8cFnaHfPX1aK5XMVVZR9WZ+WzqxQXliQd
gu9JF1LFcisq3C7vhLJObyvkLDmPqjiiBjewGcqa3FU0tv8/iePuIihh1v/JxdRB
1e/Tve6FqaTdmJM4VFoQdgiCUBdXmNXmmxZQl8xh1t2kd5OdUeDLt8sc91sCLZEh
zcCzVManrPD8Z3zi04+jNEgRrVGBe+lSpL7WhbyKKnELAl3HR6QCdd18lZpJ+XWw
azxE/mAsh4a/lBggEHI/w7iWeWq/pLgEKdWTg7onySNSrloyxtRBLqIc+MtX5S7l
RiMj7y3peVKmsafBQ1IWnpUQAgG690Kj7u03zL8hl0RbBAMNJC/BztEHEVCxk9Vs
pFuhg0HSbymX5tH7+E2bc39xFIYxW+nV2rKuL21HhJVFDw3LYUEeMiUaodnvsBO5
OnFpXj6FROxiV5ru63bv9t04hdHx8N2T/4yfVXP3W5c6qnzAEocTINmnMbEFzru5
u2HyCzxEOShgEmp7xEDkjLZGEVYrEgwjCjur8anJRPAGEprSbgnPO/FupyoJhqTL
A1Frp/7paP1tn5PHsCbR7lz/zgY61ZQ3aHl68UIq58Q8veSpE/mwcYqBobGfLgv8
gZZkjLucqqaN8skTaB5uaNaBxXGuTpQutgoLJozyaXBoAlg0CGGFW/J74lgPx9mD
lsdkkwT6RmOO/B6087SR10enNDvHSlXY7j8A7d4UfJCphjb9KvnhhUdapBJ85Pk1
c0SBRJjKV1mnX3PWIrfbsQijLHEvvyjdwFkkM6aidsxHCw+TmXK8OMLZbGh1wX1Z
vRTfHlomVgeOJqEJmZlifGFoNCQtKnYuSQzmHCQkpLDRLECpZj/ZULBF92V+pnWx
EglQF/6SSa6L5Po0dAvK+PR7kEqWp9wbfjgUtjzCFwmuv6T7+ibb2kbnQDY7HHZf
+eCDQVWzkTpOnFWkuUkmdAWOl4X/rx9cELy544slht8MHgMylMlzaCQoWidMRKW7
e2oIHHirrwkFy+8NjO4MU9jQDBlDRuhaeFS4cIbxQ0V2AEslv/164JB26AtvLRI4
bB3hXaSrZHF+g08z9D3WnitvSS1dcrCC6J7eP1mCxdN0Zb7Z1/JBT9beLKxTbEnm
uinW6r5pXt0tGqQN/5nYD/3O3tYcEXh3mka+sTe5ZShkuwBy4TKvfaxsmZrL0gIW
e1PbaC1VCmPtiDsJw9N6+RtKedArEQJvomLZUk7vnTxr04zSRMqaIcFktbZ8B8HG
P6v//iv3+uITVCCD0AXcbT+1xi78xa3S2vUtrRVrWkh2xO3qUDV43yrUslGH0Sm1
4YDzBKTQ9Yclt301XcEHd39m7X8nyHlcdZhQ/BzWhHtK1HPRkD/XaSlJ9NnUXX16
QCslxwNTjwBXVR/Oz3AGS7kLR9cg2nOloOrIyPao6o5yPTtckQOFlYeTNysuRVvg
0EfB5+5laiCYaDCPK5onmUbmwrQH+gQ/8St4R6i1aGQxNOGh4ZYBSq3CagGt52Mi
x1kH3qaHfZOO0+f30/gLbK8Pu+gKyhIuIgLB7NhWDwhAWp54FvrgxQBDaI3i5sIB
v+PMMRrI0j4pk7LXhLEK1v4INP3H4bZt1skO6qpuWDjwZJcIHANu5B1KcY3mQkfj
SWXVnG8gqjdIhFVMCyL5Z3IeQIq4GkiBSmGljcbCzwae9leT9fAEDvneg2nQiPF3
7tMZ+OSHY28o6fd3F4SJ8rRJODHzYeCAWjg3PjD3uUjgbxzw9pFXDvDz3YlI1u89
n0qFADl9o9iQLoTGv3zTCGV8FvGueUfg8rL4qXIicwz8G8sB61/LmByiYIrXfgC+
/OU+yoGFTSueUhbleUxzmaeT++wdOdQ9qk4jweJfFQxgjeLfTWzBNY0FRsTizpDr
RY2MYuwBuksI9NcZr01bhx8Sv2wH6h3xK7/vsR3V1kk4+tQEDp6ZlsfE8JWABmxz
Zm+opeRkSKuP03oPBZD82oYlOMttxN3c1IgB41srpHn5UCLsM3M5tCSEiF9QViFe
D7y3UwBxQVn/MXn7E4OCNiQV+iGvioXicmbNZDgiYD11YUJCPJFFfBIiMWqWQiFW
t/2lvmnjBE06X3rJwYPOKcDAvbKMTm8ez4ULb0jFNQxWoZhoVWBm36pzP1EaZqxM
oxFh5q/rztY/5pLtnhlvEUqVxn6NWasegp8kAoI0YfJ12yFu3wTjm0D2dCPnjO+K
K1tsTMaF6o62quNw3Shxe5AB4Ru6oGq7/s2SS4s3JvLSWKgPM3HESzhGXk4Cu9BK
63meXCpJd9+NYdE228ftQz0ZDSlicoVxstMQSWjl9cXzIaXJ9aWg8wxUjN5w9Y4y
W1Rnl6HsrYdBJrSlwHRYj/yCqR4HMniN1yaR/XwX2vrXduhKNFG1dEhSXviG+fIM
uy77NpAslrb3udPrDyoxbEDw6DNFIbqQpQTyYcyGJydK1beUG8LGWN6GNI728jzo
9wJiV+6gvTios102F+D4CP3EErkEt7VTq90bJMNmnfkFg5sbXnvBi3WnY8WcG54Q
H8OF1BpPD/a2IvRjzVxIfy+JOByK4reJdNFHzgzOoVZ1jX1ROt+dTLS70tFP725x
Tj/xiX7WiOD2mxKKDtDTsslzdPSSCwwHz+5dFNC+rf5SmZYosFa3IM0eF4JlhbaD
YPRGEKLKOMxb9c1FZFgV/bKneJi2D7olAvtdlr1bGyvvrHGpQ1AaPxo5IAtnuEP5
+iHm/8iYK26O1sPs8GncZLccuYucz7bQK4xbsVxfSWYl9q8/Qg0McDWvp4kEACfq
4sp3QCRvWF4lkizugqWjHxfSZH2ZTlN9nRmOtSdiiYDQn2jzxPxQCbSuyXaeDOWH
k/XdMvRDLw1eT1CltQdx3U0YYLvp1EH9EVFzB/FidtrqgSyQWKwMmpYAN0FXOeRE
Jl8gBIjA1z2tWhfqI3PpO0Hk+peoJPvp8ulm1m35F81jqfSceHsv8G9bIO9vkhIP
GL2ps6TLUFdFDqXKI97Xbl/L83magrfZnxLsqGlYkrYOd+oSrNHtSHmiwpJGf1hi
oDCD/5AHiPVQj/JFWqAKFUuasMkR4onZGdvPOHfAeDSZfy4RmTxP6P6hZ0slHLDV
CRBeMLEzYi+G06rL5fS/NH9I6S5JF6HCMGEarcu0eejCW6Maj5/t8Uy/xnoLZyg+
jrtBkjGjv2dW7qEFYIGSJKWX1RJQfWii0Dux9dDp5SGtL8bFrMMIdsUaCF3/GdW9
6GfADcEG4jEi2FqJC5OdCiDEW+WRTheioX5DfoBuBU8M772jxR2YZS4Qa/WMQykK
eN/TnuefQWg5P/c8EITZxUB01MSO/4lOqmh7Ar3CaLZ/LXthrmUkVLekhy0rxoMS
0uqv6Xh7YrnVa4MXbxFHCinCfKt6qutkn4fhciZ+g6HiThxNcib5uVxxd3BD8yEZ
W4kBMZ/x/Itm9J95bTdIVrGOGsSMzbsdqX2aLXK7lZO9DzA8hcHgWe9zB3J73YIB
19x1Tgq3QR2WLK77Kb4RuZ8DAt19oYNZDSNUInzTI9h+E5KAGozZOiGXUSVtT93g
r/KiJMB5UUbS9GLyiiL5HFwhvaBieiiTU/jPVMtuqr70bG6bbOALPfWGZ38K20DF
pXSFdPiidN1pKVqwTQbE4i8rWS4qudOlw6LUrbWyqtU/5BdxroovnKpKX3b4HjP9
MUpwQ+EVE4KiaqEVpziQc0GI3P/l9wS5oPkvdYwhUfcLxhTFqyKBzi4ovuCQiyUg
Y5fu938JIW6ErwaIJfDG4Pd01EohUtCegI9x/n/IM9X5D/7+bE6aI5mYgw7AuX7k
8m9+AiyPYyxrdDR5Ob2KJ7itSSz+Vhry2Mf4kpYxk0mGtZ6B7zqo1Zdx6T5Kw72I
PSZCut5jVuGAHuuT3f5FCIlhQ/NS5cGDxkfYx3fMkCfJOaaTWz7bvKH2UFPIo+QO
RRREjULamHQkdGmuQka3NjgLkZlDCckmUg4pWk+7aSbhKRKfMUPt5vLzbabOZ1t0
qZEM6DsA2M6o37rn1neQmuoloRRZwyzb/oB7HBBtyukzfVPFi1WxqmRd/xLk0QtI
m0+k6VI2r0UEuG/mSZ6FILbPO4EHWOQscvQuFvUWWQg+WZCo6jrPnhxLWbxNo2d6
/icbQC4JelP353gdg4QG5QRzVPLL2IG2mHvUcjJjI1eQUTBgOsTeC8So8OP8AneW
xghkvG2fyH+Na5eI4RSMupfMk9gyd70TJxQoRkaY38xQ/JcT6Fdks9ER56Okw/vl
aq5uQfpcv3JxjCZhpzUSLIIvu1vpCljEMSUQfydqQmyNa5A3BAK16o9iRq+BzcPN
A+MaJqi+QP1RtejYc+UEIJEZVVw8H7SRfUJesKpP3dXsoZwq6WkjltO6YVcakc3D
bYlrZgmQU/bDcE/sdRKbq84XGm+xtGsji0lhWr6hqxgILEbPtyXLc1ISdd4ygEqx
BU0Pt9ijhBFpL2S7CrIIit6Z4eJAlS2hOQpeV8UCqNE78YwqkB94iC3In97WB5uc
ybGrD6hWcWBdysv1RnXfS3tSvLIRRpP6hfbhSHdfnSWrliO8dfJ8ZH+jkqqdB0I7
REdZVhH4XEIwqndNQyaPineS8Jklz1nP+Gpqc8b6WuLLEKVqVFeV8wmqOlN7kUFe
Ij83u5RuZKPDsxwJmX+hUCdop1tgppN0pTs9iP+ZSeCLKgrqzzzv3ou9zkMm315q
xnjqvGDBTLNPF0uKeyYFJkpqTPSAnfLzNItnlY7S0rAjR9BsMw2JC7Xs2nfQQcUq
wnf2+ZfWLs4I0Pd8p1hD++eNrr3cKRB/W8iKU1MzD0+1hguVzJRigrlvRfTPc/VP
vZFKyy1bwqi64fVyHC64xqBbaWhaZqI24//SarY6D448hBIG3096y1XUbULSd4qw
aSmdwJTj0AchM4RNzLcyjTUH2QvX5oFLv7MgT2sV3rGKkjh3jnjzJxnAZKhX2sjM
V7TkEGtv9auA4trr+miQIXfO7/agi0f/XDh2qfPJgJe//585NpkqAq8AFipzrlCv
2tANRmyePTObGzGqMJ/6Criz1fao7UiaGGDXjsu+w6GIYXN/UjEvXOIgwMYBNv3J
No3n5U1FhcLGG08YoMA4UeHwPL1KBQ5ULs1BPwcflbhZzrR/V6cWepKwwMHCmlpp
15RthoUs6HBnj+Uo6lYWrrH13j7X8vMBjwYxs47SnyLr1FI6u8u4KKf2oXDvWvmy
UPHMLtvJ3x7o9zf6dhr9sNT+N7mUEuuBaMG9KvnpzD9/MbR4N+wNXyUi0TlQvG6X
YOxtNZZOBQdvb5eZvr3wp9aayWFdcJZKKUfhcH6UxGN8wyFFFnVkcy2h5lCcRkpQ
tvWyLYy1ml94DJq/OTk5/peqUzN5o77ZXt9AzhRbkmVA8/3VQ5y9aCKeQ9u7jmFX
kERsaR/98/wrq0vNP1EvMtgKx0YvHg9CwQxkzm1rF8mY+oIr3aqQZKAGuvnjsowR
yy+pPbmefV+HVyP5lVHTw6wUWWSNb2lOax4mMO9SmJZfTAKJq2g6vjOTSpyr3tlj
FebVXWi22FBZolYV+oKKBu290+mu6/TdEIbZ0Prq/w6yNDVNLnLWuTl9EKMoSpyU
X0qUkp62Oo30aaFX0lO8UqFF4niPyKiuw/bBGcCZFjUd/cfV3agg+lqPxPRzbvUK
R9a0nQIs0hL7ZID6iOiw8sHzI9yT3zd3syKc8n/lnYuEcub+jw76P6tCPKV82sv4
fnlI3CnOzsOaMtNwaBQ/wg/QbYU/0VtX8/hwo8OBny+d+GeO/UyTjv357nmgb1X5
K6khC/D5nLcYDccOF9io+3hv3BQSO7Gx21LR6A7CetwIXmVTHq0XaBfI0xdbSGs/
4z/A2/hS6CcYH52R3Sa+Uo8vNTXTv8F+Br2MfeOoJLc3NMgSE5kfd/dNxuL+l2iU
7jTxdy8pR9v7ebRoB9sazhrdh4tHtJlGR/+/JCiRFdWDqOOgB0KnRnwHyPejfF6s
5lf5G1Sl+M5WmLzGG6G3x0HsZHk3/G3vb8PnawTf8UMyPFYARiB5srlwfh9RCiCH
o/QDHiyEGFtvwv5LyM99Zh+2hxv+8ua/UxWCIq5QwIHP8SfC33QtdQLSMTbo8y7C
ygGnboNEG6g3lUKoUiZ5w5ns9yNniGhqo9S8rOn2vpj5OcbWqsvZI29LaNcaE4aD
oKk71z+OdOeAuz5oE0otr5hb1lkqsHHJt4crCLx2Cog3VE2Jcp6QYfNJQ8ZaeUZg
24kjT8bwDQcwO6/DzJpkYjwaXe//c28k/1/B93eZDvdMShx0mEj+aKhxqHprNCpj
g+iMDqQSw9o+CRTij2qkaXkNH5BbDpVBPrcqemQW/ekz3LCb/vTx03NXmwFywDvV
RjK6BdQliJgqUJsp/FGE3J6SdobnkNdTZQXmM1lCHwsKMZAgGPWbDLK3g06YgY4e
yFi1VmRSuVeOY7mWXtm1vnq/U+dFeIp5p9AV01i5dwCsQh4Axz4pNzU8gUH1ScMH
9pcF33mKxfEhic2NdTFaGBKeC/gsDY6uFr+9wQvCjWbdk1gbYiC+MpX7dpLg2Q8f
A4jBn6wn9C8IX2hNyDPKrsiG7T8tqkFG5bOWauRL7Vc4ei+Gdfe55TDBxnswak9j
/Tx0ojspXJ9ECECHh1SMHR7KXB/alqepLm2mSRtLeTK8YEfmJlw5yocHU9qRwzNl
rHclRQF1PZc75vzJh5HDalJBg0WdEHxPq0GGKtshs1p4WISpVWlkv2GVPg4gdVnP
8Vu0ly2ZG1OhueFQ5wk+1gdAxfNxX4heWB8wkYwOD/xCpssgZ5v91Eqy7CfFMEcd
jtRmhR1MVVFOCjFQQG3SNjxqfbDvZ1N0xkGN/oEt8HmzPz6q12NPUXBZ/02nlgds
vg1bzVLAKuwunxbYhy2IBIl6Iit8HllbiwVCYxEcv3qbSkNO+GGy6q/8jlwBNkB2
fsTrQuMveG/165MEjzjOQV2+ASTws6vDmMxJhcNqYTKWsI7wqzRyv9QSkR2iwE72
dXOHa1CMd5lGpEXHouLZf1iGBniA8JI2fGhAdHUKGG5fdM3RJkrU4u8uKn8MnSXv
Bh6S4iC/hb82CX6NbD4hzF5m7opKNIT1IJdSdO8qOLi1HjSm3RIXYvbWmpA3tChF
ALwDLJJUP8j8MbLM7UdOJYZdNT2KdMrVNst7kLv66Jq2JZRJGcoZYaGeEfsBDCcg
M/1nT+zxaUSjryJ/KZGS6+tmBZc9woB5vUhoDESMlX/VSd0wMfGzsAAOKgR+gaBc
f8Ji+4z1bf3o+S2pIxAYb2CfyNi3akYScYN/FR9Cup5bBmli+h3OESdHxIWskYBX
t3Lqb5TVxfUzLabbSEzhyW8BjSe+BhHIEhHnyDpJjqWEEDAJm/j97mV59LEaDDuU
CM45IjKSPmpcRzMPVyFwDmqObEZc3+TQ3poJ3REQpciDJbfPlS5iyBcCvkl8AyXw
3r7EpD59aebJyRbb2ZiBxI1uC5EoNf/aAd8ibffQ9yD9ziOOSgITbR3rfPpPEA/Z
moB8W82VdYS+WKesotk1a/oHh2LxISpfXRV/x5auQj5ji25Lj2ybL2XoeIxaZeXi
zBPuBx9VC86fOzZGcecTXZkMiqEOcEamyezAR+H23h6WYBh9S5gWJfhzraVdNzSe
LBCFW8nWCtRPDRYSRiXgSu1SY1eRVacSCj/uhBB6KzArkCoQtv9gPX1emd3hoGNR
xMHG6iP0VcbD2nZL44ywuA/aEgIIujHgk6RQq2HWgK4GN6g/fSoo3YUyYpB80rgp
AehA45Ve2iq4s+DCpRPkeacv71ezcnv6ElzV62wsLEs0KrCNmBRzUHNt68e/uAx9
zsa+W9ml9D2Hv/opvppQc+s3nTiVH/SCrMOoJQl8uKceWWNkiMDmXpgLPxIrLEJu
vuxJneknV90kGag4UUmsV6QrsBsdP3deLPMrFS2a+EGj6UfXGF6LH9HrJ6c1ZZrO
6JYcw+LFURkW0NWBsF8SbqedPB+xDqWvXK06mFShT8fVV4kSePZj+IYCegS6zrFI
3z6jCL2Er2eNnWmOhdAu6szhxgd8cek5qigNa1RoD+NLdajiBuQWL8U7vQ5W8QyE
IGI9FC/MzmpNjr00t9At9i+X06ySFyBorogzfumfHGe3lRnqldzOpji15mynl2vg
81Cpk1VU+m6fXgs6aBxtEw54o8LzsmV+hQmbqoZg2dqKmoDhC5QqNK4RH2LrSmMi
tVHfLBJtGBKihJNqYnNgz6XUL0rXA524/AuIpoZyPP8FAbOc6paxQZlBe/uv4wyi
0EuWVYJOvTpqxcDJlq/7A6kkEu1rADhN9ELT6Vk4wyfgYTRTVVBEU5oa07apjnSU
Fcdk6f0R4x78TYoYMus7KkHFG24OM8MNiGunAeDPzNzJRVAPnB6ych/VG4p+SCqg
Tro8hiJ666AYgC851PgOfspHoA4Q5L23u/r15VHY2ifPcbh4Qald3V15rzdvBdig
raKhFRoMiT6sl17VN0pBpRnJAO04JWaUACZbzUl68eLAyx+PgHGtO7w9IzFfuZNa
jiZ+Guc7G86aWgeU4gEQATaBSyyaPpeFCtYCA2U3bC/3etqt4zgFumLJ4UCEfBAN
gcFfXQANpVe9jUS1FJ99V9O/A7sOV4/39Wa4w4AfSHWooz41ej7ZbuJWbEGKpR5D
0lTsDS28HK9IztFwuP+ht3E1o2U0JxfE2gnAQs+tGCr2vteQS7/hMYgiuDPfHTXm
TKmafsLaTtT98r6yvyNoT7PvG8X2bgMmJTjHQd5xEpLeOaXD0W364xKRwREotb3o
Md4cpIoEP96LFCxSHQxSatsa4tMhScp+yEqnrb8OY1BjbJm7XMwFiNEKuFZID5zO
UunU4QY394vF2k2MOzpkcWNRSgljv/jxDqeHRMM0qNtb9fFc1ysJfne2ujUX1BxH
EKRbWs1PTLeWam4tzhEbbd0CCH0W/sb7E5wbiHr4XCvdLBtGdiWqpcP5l2EwRChh
Z/HUrJv0V7ECxbp1l8TWkK6UpC2lR70TPePmEFDppmN2gugoN33klxvFj5sI9yr7
T3lNARXbRjc9cRx2OgqpZkoa5BHIEeLxLCt3dUkBFmBByR/PmQHF0CHc/bwcwHoi
F5jLLolthJ3FbACKX7rWtV/PMvhkZglhqOkjWigNZGkS723OJtawUsdnW6h7g9Ls
ftN0uU++Cfqc1H41yV/3iOr4NbqPQAkgC/Xe6axqp7nNYTwJ2lNSE/TTqLjiMC4Y
8bkykTFV6zF+vh/E/+m1bA7xGMV5BbVDKIq93lX7zH/CWDh6ZR/I2UMGXQjQgHgq
1UNil3pTmAqN9xgDAniJkqADJ2QsGt1vy0Tk4rtsqcFUpkzSjs6jOe/HQk0oGybp
Hkht2Tt5G/9xi22vYfpwwQvEQHN/FFwwzb5lmGtd4j2T1IhgrOJLe6UVJQI6RwYn
UWf79oX/owu8jKgQ6bNpN3B4VZq4QNawU4pO52vlmPRw8rrNSDat3tihw+904S72
lPtx1YpBhzFHqIvpIc7CIaYWnG7p0qiJaC/+by6MguFb7fBbonXdAeE0v0z+Sasm
3GB40tNH+2pd64+fszKdnfeDh2/Y13IYSoXYyha79KBdHPeWANZX7iPQG+7sxPcH
37P+hz8JtY8e1rrz1oLhSbTKqRIgOiyYlybNRoj/MWxe28g1hbfkJ/B6yYMjE6Rb
L91rlWR71+Y0rLzsBqD7GbNv609CLmfK/EhJs9Fdq5flRa86xFf4hsIelHn2eKU7
CgOKhQHfOYaRJWpdglTy8dVdWplEWdhFuo7/0NEem1YJDq6257I4OKbNqxQmNmta
UJPeTJQ7mklqiKkqMdThXYkAB438dd1szUAXlX6KmyWYrpzOU2Dyb9j/wOeFKxZV
mk54hqLgFTshZpo8PUDZA8/gzaLoO1/BMxPVmevmFaGiqk5LuUFHbcCFnCcsT2xi
RN9/BtmU493rmNGpJ+GTbA9QkCuOq4gh0eff5kEbjXdZhcXthg9WNQqqlwO+kV5l
7SRMSiDghJy1AGUKPpvlXTVvgjjcTGmRFfm59A+V96cBeCLDYuGL/67xCeKEIjmo
HPHM1V4eE3HusrrjT1Vx+54gitILEhaWAC2Kd0pJXuEkSOLHfX6mOckRdrFzjXG8
BC/jHpmQ/TJ49CabFC/Jzo9Sx45MsjE57qE/MNm0xI3nE+KCKI1hvzmL8/zqvIWn
lYYL0GzWZTTlQNEpu6/JmGcvqd9mmlqQT5Z0474DrNMC3YKSJWf3lh7If8Tkv9nv
CCCiRxdg6jQoWSwhsyv9jjUrxMgDypnzSQF1Xjh5AB8+rVFP+F2qTgq43k7alHSp
hTg5LlCh9DqYWmICt79eOAaoQA6GkVX0ih1wIvzHiPDchblO8PnC+TefL4S8rJj0
4C4BP6zQty8vqPRiQ6hiOgXFI6lbu2yxGK6M3uYyJRhGYg9Z4FeJvEbtnOFZeZ3q
edMNIwdkkqv7Dsg+gqKhDQCz8Fm/rCIN05PxGEqREQXMJRiDbfHjVivLv093wBJ4
ELRiH7HHBiYJyDpue1yZbFmEhQYnE7x+MQMd0gtYP8bZ7t4c2MQhnbn2fBR3nOqq
d4DcM7VaDNb31HZHnbbpewjiYLH11/AEtTiE2bANgCiq00pd1LN9bLAcZpvTFr5w
NSh8CSsCtzKc8FVQUBCGeJ4OvuYcyFDVB3BKiMw669pOtrySWMxNZJIHN4YOnQ/J
CD767D6wtbj12+xMecByc7KOJkcdha5ruK0iOIaAl/ZcWVbEhHD2EuuyxjCP4mAB
bhIkRp2jzeZQS/6+EoHSJ6Ea/ABcclD/IMKhZvK+SFNR+9FGyem4kTuyLyOasPLb
i0eWYsQ14B8ICLR8kqtUCd+Xd3VC0Gy/ETZO6vk6IvcvT79OeUJyz7kVxQQVQ594
+IwNx5kzdMzEykmcUjrGPXj5yP6T9CWcU0OZ3B/TojUc5mJ0dSiAgB7vs86s743A
9+4u9tMX4CXbNzpKcV/nY0ZPDbWT2tXuqBKOTLOpYKiKBsaBHWuhReQ+wfFg6Kse
ME8Q+b+1e/zy4SM/gTgmM0ZArut8nQDdwR6IV+muTGRkWeWFFty1QWW1rkVhIyhv
IxLd0cMM4xZr2Uk0R+mf25DslHenKtom+shuaS1eK/m1X6lY3lRXYTvyFvg0Yep7
bhRChQ7vB1VU749mvBArrzrH4XFu6El/O/bNSC01ng/gD2pxznkS1FHzxxlt4xER
QT5NCmHwNI+eeojrKtmOXsZCtD5fFLAa3wIkoAaMo3u/E/7W7BgDdnkFSzpMj2bw
Uw3uf91d7QwoYm5yeVAgFdEC7wWVaI2IU7B8daor8MLj3BKCRbix8m516z8vfh66
pfAsR80ZYCm8y8WFCfWCQXTWUBMsOIBbi28Pwrd1xAkRTuW529/NiwdkplqJn1BV
xxMx1mGSg9u/Nh9tvxq1uMrK4tC7QnHwkzTJ18UdmbTIAu0NzoDEy4vXxJvbPoD8
X5BNy4Wln5hUfFhjdRVoJikHwZIAIiDw0y1xJ95w6+1Jwhs2absGHTKgMtzXti0R
UGtDM3IS9+Rb9WMcPtAklTocdhfZwCF35ss+sR45nNdwCLaM3ioRiIAQWLHeBfcs
od2K0sYv5V3C3FUT8wlbVnvldnTH1Fs2ABarU3ME136e5UFzwWUtCjd/Alp9N+9V
gMATU7yhLlogsbABNr346FPPmCf42W0VyMxJS8hEsZawvvdl8AETMLd3erVaAHEq
40R7YJ2AxBTR7pWREiGPDxVkmOIbGoWiaLsnjnavmNZpZ6DbxFWA9jCY24k0O1BV
JPxq6HaOuAqBc//HLhcA2mjAdSC2hPC6jFMy5c3nD893WBM7M17NM8U+rlOsMJ93
jXhpyYCzaICTsGWTRtidj4JGs9IrBqqaPZhW+GBxbOQNXc2LvqhOf/9VFIO8VGHv
b7gJIhZ+LC8DQwiIWcFhV4UgtQc9jT3GtroWAkIz5Cn4qWIb4dj+8BQ0Jc5tWIxz
LkF1IDuptUHnJ40FUOfj1Ow6+sVE2m3KlavQCp3W1bS82bqEympLvI3xeKT8TrJA
CR7BF7wZzA8q2UnYO78qaf1Q5+vA65ouZEWOB8SPW/tVVlwG7Ge8EHLBRE2avvGz
lujUGUZaL30IMGgmm/Vks+AQiLJncuhqHiWGP9/mi5TdHxDIl2dO6f0st02mhMTF
la+NzrEOgAFf01zvgbwbrjZkvXNJSEVFE5QLWHnIHp2h5MOmAsJcGpGA8yJm6Osx
6r/aw8nXb5JPgcIGjTsVSJPBYw3Ou7mtuz4WmDvw1kB1HtAvc5PA7zhXuLjkSigI
DTaGZ+XR7grEYnXUPh+fTz0iFFOtOm1CNp0YEtQLHyO13eDc7klueFLEs+pkCb7H
2cu+EwbwxMYTgAf67spFtYqMtxNtuoDT06YMQ1xcOsccyEjVVfJbDdGYbHH5UbI4
3k0UFe7pCbqIenhkNia39TF+clkmP/AR5y5k7iPPWTBDEl1qm/JbYHS2IcFvr5i2
uniLTQH2eQ1fYv3vhe88uQc/GRNappZTHtZvXGZFRR6lk1gH4hFd6DEFNtURqeI3
eFyGvJcyqmud4rdm5fuv3mCoo9ASiLP2PVHd1XnWOWgynpKN5KHcSsmDdSt5aEx9
4395IllZMOFn5xP+MrRvCM3Oi1kHNf8rBD3G5FRVhubdIhLz6DMk867Dh3RS+Y4G
ranJHJAwWldar1+CsdH9K4jWSR6tKQscR8itkD9u8XxAH0MNC6FAIAWb66tK76uv
O7E8g4QFBbWgzYo2am2d36AISyLId48IoXFN3crMn71NqB7M5MGmWu3dgaJuTm1j
Tp/fSyiwnyzzQ2CdVWOA6Ozy4EjvDLzNu3NKEZ3ngoBZXw/tBwsqzGH0hRlYVylV
9QL08E7a68jMWpl9Qr/jsn5Q5T/LbMnP6xtHqnnGD0ad24mnFVttFJ7tDfCFO2eR
b75J4r75gEBGws0uMXH//eSDzN9djgBohAXLiGnKo+dIwgqViygnTNbG1uTD9AcI
aWEGa0p6AVH3AZoOIGSfj63iKfVj62YMbN1amcQ1z8XBEVq1r4ukpnoN4sa0ANm2
WaieELrf7JM9Gj/322vZK66CoWa9DJRV9XwijPjMPTds/TuwOPKWr+0c4dOqoiHX
2NcodUezQkLllLl8Lh+IbNKYkq9XlgdXEtY66a4QtV16pI81CeSYYE8llmzDq8BJ
gOV2wiQtRqStazqSeeNmrK4THjaMQNKayUu3KgP6foGCcnOM+uq3qNCrbeGp5SU+
VWzHKzeDzXbIrRMXHE4sTucusqXC1QOuEPvMFsxePaNvmpITjEE7QypUtUJSebEN
wQZc45Yf3mQMZ0Tll9ZZWIzMxZdEtAHs6ngDYkNegS0K1VtL5v0C8vC0TC1UOvuA
PrM1zbxNZjTKps42MCdLK/YByVsNmZLwHG4+jD03kKIbBEQqibZSX5KkQWyvcgus
5dGQyXm2Eo788F4gb5LAcsoI8UGt1P8Nv+hS/AAHfjYsMj4dVsOQQYKcJvWN0ma1
GEGltsgx/OH9UIM7VcmbzZd8TUSy5HpKU8qGWlzGPIyOzm0NSPdCvcPtdLm8n02Z
RWEIME4r90Xgtq22dHVcypuidNuCSkTRS2/zAwysFPHxm04kNHgMHv39N+FLx0MZ
+zC41W6xZvMeD018chwSFY81wOgY28gfp9JpECxddYUuZOhDsFiDeCl+Yo+7zc/x
nxjQ7bulSE3P3FKTFHk40Sww0MzGNIvYjKG8NnMDVZTV7p0yuNLO2lL0rlrJVYsO
rzHEMHbBW720UI1zhqWJ6bdBw0toOg/O0L3WuMkEmbp3cPBiuroMjRHRcb7fsiTa
PgWWCi9gXVcTsvBKTPYQz+54oSpj5xfP3/iHOz569K2jvu7VzZ0rNIUKl37kjn0U
7fJuhNDIq9w+Qw/uZoXHiZFFqzY5hmWVOrGZ1Nn0KcasGd3qquH5m1Xmukfz44HA
WOOodQTpiRCCvrYd9xi5tsDjHmDqNaG1cWa7NEz27cZNcs7CGCxOj7+dJcf3Pwsj
rHpK/UYXTjm9ZqZPZ4RlK9YuM0Qg4q+uep+LTKNdXCJwoabxx6Jpc4ZxIOd7nZgC
9IZWEix/CH6MIXJLGpns+NWgnInWJ/YW6DOJ8hZQRUPxgJKa74v6kjJAifnVEZ4o
FQkGyAxvQzr/gIhF44Ea8mooxtd6V9h8dPq/FX6STHGZbgVImwgyPM6byOP8RciA
HCQuc9gIkHBE2r2xnfIQPp4NxkGn9P5ezo7F44qfOQkVsKuI7AHHq/3Yi97T/VfH
1gqv3Tk+Ss6BRV6Dup7jmxA1JhhfcMLPuR2qpbMSHjmmlRSElM4D0YuROXfthVQA
uWa1B6oxJv+L7eQT4i2GYSRTMFVMX32t9c5kqTmM2wXCyVdbsRTRIc8Qkn+ulTHz
hRM6PZWdrooR4J0oJ1ZKVoPl4Nd0oqxHi5oKQhqIjhZ6oF9Q/WJqO+dpH4DnYWaP
7HPcOMgIvdlt5sJcfL+G1Lw6uof7R9DqeRHE9FxeNaEm80x5FcX9je5iFCI2dyHQ
PWWdGKpwuL/TFyeqxffvBMEqTMx+snCp5N0/qHLNmCCuIroY1zpsbaPr0N3bJLPC
5Up6E6jvOJhFq1dDrV2b68SLMUgjOdO81PNFSsPSI6ZRp+oPxFPyut5UPVh/K7GJ
s/XgDub4Qi4iPs5M5P44RLOnLE6M/XGik+fd1arsa/QrZ+tx1FXO8RGnaQ3F8Spe
hgmDBfjWEeSYkf08MlD31cy+ngVJjHGtHg8p2RnW5nUzDANwKxeG6EsVSP/ULMjz
eqoMmN+UmQlCMLBZQ/2ML/RsZRvJvTA8dJZxpdtIAghZ6G73NSEbDzgra7fVj7xh
LLD1n/RTJRR+aaKUQlPAjP4qGQi/aY/FCUQCKrpzWzJ/FvNQmnHdlCCW1oWIpl7c
8Rc75MOR3fzktUS10MB52wF0S82m9aEuYW9culImewnF1IJttuBjYUyJIQIUeTD6
lRNlo27jEe9hf4eXyp2Eb554NGgPOgNjndEmehDU3HwWiVit1NiOb42v0GULmV86
E+daQbDrE5Rrz8u51KaXZVRVSz93xntZ5orG7Mzi3cmwXWUH2cZebycE2gNGvivj
Pqz7Ho0/VNjZoKUuEs+pB+8UzaajQJJKDODs9lwXAjDxKiAGBiRQ0OyB20hXdG7a
12I26w5WQr3Bl6dhcM4VjLUlX2yorvOyq7plmUsuawlCGGbLoLdxn+XYWu/fvl5/
k9kCmnHunuloSs9nzKBSDN3iftdshoWLioOxd5Hu4YxrDomq+9SUVE/+Du051Tkm
wa+MCTixGlYV6LtlOcMDmMun7+AefxUQKurDBecdAdVd590yQ8j3CsZkq/PTu/l3
zOWx8dSY5uXJ5Gt+QTlKXC26IaOdWMPbx7d4KCI0dUlZmzr6CQaq9tIuPD6sHTW/
osK8lBvXWCyMaGXMHL539qJnhCMCdPA4w8IQT9kqVlt7RUKNepr2NHpf2VUa+dSq
Q1eXjzYQRKp17huoGfETP7FWvSC0OJzSp4OM5/WeZVQ5JxQzzihSh7dkpz/54r2I
2wS/VuaG2GfRjhKw/Gisok+bTFcE+Bbbs7DMuuQq4JOzw1K9Dqcx09CH4XuzVH1o
XQJJm/i9irWQhDnQy1TG2fndDAQ+awuYWqDOHPeh9QfX/Ordj8wWcSjo7IIhJKvJ
7SRU1+LVtIGNDhyju6jCmIVVA+9Dx2N8NTyW11KOIpNqZV9I4ywsO6LtrsA2DNF9
rMchNEIxZ9ZVeUtUu6AIcJ0NedzjQntI/3tQo1djD5qEJcR6P8Tsu7xsTJMIXcwF
D/TzxEyM1c1D+9WQI0kAneOACA2qI/CvDTcSAvatTUzhCtJoMmehv2STAMdUg3R1
cwOZ/DsMEgmzj3Gy1ZqFruKP59Hj+uloPk8o7IRcbTiIQc3vhXlbiGrzJkLXXORT
+QoYhhtdbQLJOouaSRfL5MkQ+qguia184qcPGP9dPn1P8VNuBKZgtSW70O7CDiJ/
lg2i2kuN0Sb+NrtdWhgMfPXXGO1VyVA1ZwdQ8t+DYwQCIrbKbDx9dnhHIxy3OS3L
p/nRh+y4358KFplZu9bxai4PYjt2AILZmm8WdLaGGhzFc8MIh4swN2Rchk99WoSc
zWIEd+032Lb5C2rCvsng88CYmvavA0dqumNSvNzmWcNSlPZaOwoZxJsenSVF4Zln
NTKfur/zRqWFL+m2Oe0Gc36CY32pkjvvIPT0RiHLT8kklUAiPYLArfCMnG43BMz2
CwWt4/xK2rArvCKu7OCKWbXUIEsWYe+LeYjlW5TLRtd1r9I5W72HyvlWFecOlOmG
u/Z8Y+tyMnhoINq1oxNiuXO00ifGIgNK89tw2MUC0gkO4L/6rH+RxZNnvHqgIe0z
ay8k3V2WSHSo22nr9VHtB8vzRBGJxEplp92B/IzDksVoVQNRkPbzAFfnR4BxnyH2
q0hSxmqt3lzXQ9bn6o607YHbzmnx7WuENUKvr0zwy9hWqXEG1AFDzJf/gsjopi1N
r3yMFrQEL41AYjFBAEc/mdRNjPWed2w+KTXH7HbR/T5zQChAaLT/KSn6dLur2Rwl
14JILRbno8WG7anhWxy/tF8urZ/B4N7m/CaTOj6ob8/jUH/6lH/c6mHVK6wtSxYM
Wd9LEu2nCDkWsrwQwx/4U3UD3HB4Gy5LzBuaYDrItrXGrJ/DMd/5jdnJGqG2cCId
VAxNv54PSvfmh7tk6HUwh+/uzgfWnCPar6fm5AvWG6rbjogdUOnHuR6/2eChzGI0
AKH+GaFtVb+0khLFCGCXVk5XYKG4NsMVTBAetaIn6x/w82DJJn5IW/mK/kUi9wZd
VBqHiC150TvhXaKHb1cw4njxGMjKSu/Z//fbjScXvK8cx0mBU04f+3BjH1V5gkb8
BCKnhQgB7KA6+HSHKmX+/GWTnCDNKHBE5WyqfWSdIrQFMJxHHhMJNHUyaqU2GQ4L
31DiW316EUSzdUW1mPZBzFkPTwc0oZSCvjtjBlh0KjtkPGLKIYxHDfGvrYuazbH5
ojUVf/QgXvaY221dcDQA05Fw19SzJfhsH9RhQMrMDwwzAScB5xTxQYI1FK069r9G
sv1GqJWWvJ61iYyDLHblgYQlTVo1I6gCIByDO4GlfqOGX6gEuiSiYDUawPIFLkv4
R06rRvLv3Fqf/N1uIk2lWPb4AI+hyrOP62uDL5PwgWNwRPpvfDC4h4Kz2lWA9xnG
fUIDnB2H1jAcWa5Nq7N4cF9z8OM9OLtdLRz3GvgY1L3U7hKT8Ri2wthoBDrLVzu2
rLDsUf6Usnx7KwQu1wdeabXm7BvB8duFaZroGebm0+LLkpa1o5GEx+7/UXr6t/vt
HDTqQA1I9QsEccvKtM5iP0k1L4qPXA0Ru91HESKOJV6OB+3yIone2KgZhni7ZnsZ
kLrV86SNBDIqIAeF/ej0JtvrhcBWrqMfNkUBnaScCSKEKYqxMO97XcQ3EI4ZUJdM
Qfn1c7+AJ0/xgKmHobrAkz3XFXm42B6kiakQNKY6a3aOoMVBSIj3QjZtiGa7eAnK
KZxR/eRM+uvoNKB/re0h1ZcmCwGv1DBp/cUFTyrmB8oC9scu4PzjVfzP0oK/vumb
bIT3JqMveJZevpv7YQRtjDTh0fe4BYZbZlyLf8BU7e0CPCXSY8dNGX2mTajSc9ei
8NdfDPfnT61wTwUVqQgdvFwtC5Qg+l0NBFzwCXxa0eETFcA/sqQEuXaPAnrUUIqP
PSRfWsImicGQ93wI7N8KZQ3engzipLOeJZz9V2UUl/FDnr4jcsP/6d7ov8Xmtrju
3DECTCZ5KGYBK+3Ic10Vtjs3HeT51dMGxLBqPlWZzB08YwgrbJuqBp3Is3rWFkzN
Qbzs56BleoT+Al9J2KhYthEc16OYg9EqbIY35Sufo24huKnaNL6gz0DO+5SO4y1N
PGy+VeYBDhC5Dcq+PzSVLSDSmanuIw8BwC1GucdHBAzXPoyafIrcvMAvnDPz5JLR
46LzXdoUI0YRw4UmxrbHrgpU3Jdb02TfX1+K+kSvtRycEsglPuV4xFVA2jKwlwoM
ZnhocXBPBy2j+5Bm7Q71eHjhJ0TBwEkd48gFSptjSdjRX1RVTM+mgvMICGigtT1w
pN9guloJdKqU6KGxhP83/ehZgM1de5iD0kGod72i1fE1UNx68LwSJ5BodIQGhPTg
mLXJDSBYxa5dcyPvhxxW19kXjo0VMTyuqYTbRBTXRjDQh11yQgF1veYfmn11RHTL
x7oCvuiyRO3e5/kPz10GSvQvSzJhaYhJpC5+0t3kW4SfKOIs8XNHmFUgXJkcgilm
z9++4THAF5HkLM4plsRmsv9XwRlCMYO/py4Jq0zBtG2S3PclKt4s7xe6/npJCytm
8otFAon/MXEyK4MfMwOkfO+qRAYsGUTOy9qON8Ow8r0nA+44h5jb1dmssY/XAO9A
+fdC4BG/2OmCZqT/qr0d/6yyyNREeK8G9sC6B3GHXQnTGFXTSPr1ZLdNDJX8+EMW
3YeBqX6CD143ksy4qEebDhNoy8JLYLFgOCfgnQrCm5CjC0t/J2HqDjfOPtMyYy1I
wU1IqtVo1Oq3TKiG8ARhiQ6LQkgNVSGbcwbOeCs19gWxraf1SNJ9+lSH7VGDVx/Q
hVFeWFGgcGlPU7UNaJISKbp2qTzqFcUAm95WwZ7mPVSiNKUpMlGxLexDscsbhqli
i1fvIcXjG3nwehj4NS3DfOYDz+ersqgAAjhlT12TN2qdwK7vzRTB1dLdhNR9AxtN
zT1jVO0jRsGxf4eeJ0ZTPbU0s8E8jVerxH4EIQMGUOKCRUqpWmtxAOJGjslMvPAv
kYT9DeAXVgGnUNIbOIUTg+Dq+9ou/TgPObN25bbARfwsz6qNTEm734NxLony16MN
TiSQwotLBn+UB9Nt8tvR6W/rpvY004ISh0THZFiXukUrYRCCfIwcP4YmViL7zkOd
SXIX1vqoK6B/wm5suLKr+ujLXcphJPfdOQ89M6sHGtk4AQi8w1yHpyBQM0IY6fRj
QhFAhQdFMBd3Rw//M74lueXeXBGTZGF+FefGxbSf/cxqEXV0n9i/jCQqDojySeFp
WJEL/kv+wSywQQI0q4+H1BYbFsEZ+zSU3TRmJ9jO2RtbzMkqqS90b0YNQwArYySy
kQKDy5HMTVeCIK9OQPjzE27GPzlLO7eE6lI3j0CnSzk6nFTK1hWwZOTJ+e7mR9FR
QrqgZuHNoPOwy1hai4gdhjhAzwFtH0ZQBu0ryOMkmTcH6pyxVrUCbdT6UlkZ5YmP
lQfEjUqW6zkZN4r6qZr2HwYh+NTwv+4m7X9/ee4LINNgoFQN/kvAFF6ppoxW57Hd
BDsxaZtZAB+z3hcG7ozAecoDlLug0jkjjWOrPrXCeY9dL50MqtnXyFZyqWQELALU
AqHDvxRHqz24xHQsL78lGmKlDD1+k5QLs75kcAYp71+YRobXoqdI58Ifl5xcGrmi
U6X71KsUlM4kbHgnt7FokxzMB13qZOoZFk4Tm63qPdaBVjg2wE6Fa2qIpzYAqas1
ksSXrfsKcELt2QIcUKkyeRNN4xReVvqrZMMdaGNJuYl+3HXtJ1yiL1f06JKTBYBU
tAqarR1285RyoGT45DnFfTgRHJ/EGxvSA1XMkoS5dguBqC4r72iu8Grqnyl+c2q7
n2Fv+D2RVh/w+eSje8cQ262wg7Qa7HxVmHpqSAeU3t8yv0bnA4TdYD7pwqQRiAjl
GHctGMRbdJE8IHhsDFgL34TVN+xc/H65SCfi3KmOBppYYExkecCw/Kon7b2H5n12
AKsozPipKVicVmNmlkxWvjKZI3HSfnGWB8cuKbsKNtPXbvAmbwqJ1UUsV63ExB1C
zWLHrzcLYGwmmDfuBJbNnvuRXj2fPLLMeWqZoNTABnbghpY3i825UE12lPNJWEXA
llH39ACmEDsuHFkNPMBkdZD6HWLNygXOoW/SZ7F/CSm04EFS7ouVvyPzYBeOhOJL
PAR7Eox/Az0W6aE4Yu9lF6rbQCiETgGjBWR1fkrB81jPVavJg/blJjjxkEyhVC9I
4j8z8+QTVpaWDkFSo0EO06zDPgIzLmoF246f+Qr+1xkI0rP052yrJr3smiORRbHx
CrB4bXHzYE7Nvt8Rv4Gd+8g3W6ObszF0NDkOMCl3yTbpd7DKRlzL0YrN/L9e6Z/X
yFil10z0OzLZ2n7VvrpsMn+8NocdPrano/oekCbhiSI+gEkDXSQMIXk218oRnBCN
U0TmsRBkoQR36zyjuw3f3jQeRQXEPg0NF2Js9CouQkd3qjhaz6ZWv5G/UyOj1gjO
VNK3ka5RdVoHeM4P5ilm939zLOjr2ElFCSMlIJkFNsDi5Os4NLbIQofov/x3pWQO
KBOFlp3x/iRU+tqeyLltuhQfMXoaSSzx91DWvPq+vV4MeuAvd5dv5dYJuEXpflka
E5TwKF8K2g4CnM3VP2VfhKMs4ifhWPRy9gWyN2kPvSqG/N1bDQ2OkaIQ/n2GF8UG
xG5k96cYF3iV3aW5Au1cMyCCN+hMwiX4OuNpujaTOsT5MK7B4hYizwIfpgsbWLV1
bWB/88RZZGQUYeG/Y3WqXwR1CzqfNzf8GVhT4CZZu/3XmTMKbRzTTGNUgO9IaQjt
TUSlMx+p5FJLhWrG9D4J3T0C7IkpPBLfZRjTZs65GsDQVu3ERD/eBmhP7+AcWUYu
9BmyNpCjbX4s0X80Tr8mfzRjlvUpLm/HpDXUGlRTpROSGRBs4i0qwYLyRxrIz2rf
ww7m+Q2HF3GRIwDQ4JdHXjI9SMuPSx2fPUPZ/TdnXw/B8KFROyqByCBEwN6j8f52
rs/O32yvVN25QrE7vLuvzYuhFlc/gvuqW64znFsfabAcyCTIkF4qvG7WMHTkRCFo
MntNCVXZuK6w+CZVaIEM7252Mbf9GkkCGC4wUK/iPOxaExoHr4hKnDFTixydq8XK
KCJRCneyhusEhdTyUvns+/aJGMHiZfPekXbyoNmJtaelzpiZJzcEVe1sRvwAHZng
j2RZYDHB6dD0+pg0/EhaVZavpb3qBYZPo1PAAsxhDAIDroFKpgZRGcsPguUyU5p9
zap5pgZ4p91LisAQ0JSjrC9+E1TIO85b1qRWjQnAx/UWcd47oggAoIWiAn4w8y1m
yMflygfSs1QVUfkJU/KOBx0vriBQllNYR9gCyeM8P1/vR1dWJEaiSU3zmdLkvk0P
557cY7UztoHUmxYj6u9JEqWWqFucCJFpS7D/w9MWjdJcdUEGg4G1CuU/A8tZXbJK
Fm6yMEUi6Hflf12dkUC/Hwrk3Z+AhCCmXmt5t0CgzI7kGjrcqyaN1pNCCrzNAMli
BYcEnvCLdcZfVP3rSQ2mSRZ7ILE15sWQU4LFgpLTSzTJCNP7OITRN6L2mg0EjKJX
7zikS+Arfaop1JvLi8RmCn40ELgWbFoVvw1i7JF/szeXuMxW0iFAKGgifoEZbl14
9dYj1lHGqrO+qOTcb71dheIeAeG6UyDcsthdBIkEhi8ta6ZjrA/uscwu0uEene7O
RlVK5U7xkRxycLBxOJQa2JlekqqavdlbfxWoRCdkNzGikw8gvDLrxATik/bTx2ol
2flh3VBSn39cgiJKBL4WdxISwx3yOeyXxhHSlcCxT7vMrOuzAIuIp+ew3lDLVImY
vcaXL8mFUculWRjxd7dTIk2wqGpRco6w/Mgo0vGsA6YC8ccAOhAfzY3Re2rWoiqB
ETcPin6FetkWCqOE0Yj9WbeY2//5Xh0FPLegRA4TWKuvGclvsAL6cTdfNCnKUxTU
AYTSvwwAw5Vbow9xXD2CbNqT1Ov7F40elUusEOKOJgWxkB0uCAPXmjF5R0+AX25N
bT+yFtgKbjnO4gEU5ykYU6y8yHINRMrnU4uESkmmaDz+O2uPdeujdsm/BqFHJfDW
bIKLLhbKFgez1ObsyLvt5b6ROs2vyaGJqLa4Vcr82oZHD95/RxTy1QZEUKW98Y/6
0DARh60iRriPbSNycj/8JLT0/kxWGmtY369vnoM/qR3SUyBxPAJd6VZHACiufbks
FljqUHWacJZtRzYioSssAtZV95fHjeabWx04Skk4y1an7cDbi6r6kPQb/5rakZK9
2/pm9aubgZ3fGmdDcaKVbNf8spOYdLkgTTfoGIdBzD7jH0XGmuEvAOfhouC5DMHO
AmFZiNI8E90FwfpLDRHRbi1FNe1HpaGHc6h2ZHHVk81AKw9yYLf9JzbZoYo47ZXp
3r8he+OeD63CiIg9pHKXDtV9k5MBYqIUNHgCGpZyS0wpODHrqviGFEjtDU4Vs+K5
yP6GCaKIsT3FoCq6wioJQhWCVnLlChJbnN21hIRlkjZAlpz6s91w3dccOIS8mgDa
3yplEFwsYcFxno5vWBt1mId9SPObBLjR3t+gZYx5iKMTMFETznfVKHedbNbUqTpz
K39C1GeHI2aaZ71hCQqV4Fb/PTrZERpJOHM5NkwOANQ2Cw9wAakOhX25nA6OPliD
uVeOP7HwZ//FGGzQzIwJLF2svmaY3edywSQphBI9KdeN9yH+/hfxMV/sl+Y1zBR4
64LuWBsTkwjzqULw/q8fU+CKTJtZyCyTZxzUymcdfdSsXC5Iyu1ct38mq8WFxvQE
IJoHLGVh6jKppQGCj+XN4NgyHpU+jZzrC5YcyWgFEcIDa2XnN/sq4YR96tjmgEdM
wj2mWTHl7QgoYEwhhlP03WYDo9NrGOtrlRz0njqBdwWPAYkqsgv/cnCniTxv+vFt
xIS89FGVjmDwvRULRdgG66XfYdBluIrhxUFSXZoGDSPK1lcmrGoDHpf4xpcw2wgt
MmxZ71Bl+V4V+hGniKv7VxoM91uIX3MyNlEHa5DwKhiw70osoR9Wh+DKqTBrxhTq
OSe2O5YXxZ5h1lp+MajhhJBpIlENgzSFVNykmHy4HkoRK5cKubhginPkl89mZVBj
wRLfM5qPNArfV+MSaK3QKISVHc06OL+2zghNGtPTuN1tTpMGfScB5GsQyS29Fovn
duKBDTYVMd3uDh01oS0iDpyhZCbsnogykxtILV/rbDzE5TZbbJ2YxlO3XBt3jncj
j8wbMKpdJAe2m5l9hWGhEWGc2BbdRaethyQox/b9mc3aF6GjrCEqkR4TKYtkAq7p
5qVsxesAQzNQ7imIrdrXOrENv9u1jxx8q5leN8OKArWDEY2qiIeQn9i7DeC2ivlt
82w5HVwbPuwau/CMoJfnrQqGWp5ktKAaBFQ5Fh29aHslwqPPD1HGayWp5opElyLU
GzzoiTsSqYWdstJ8+AzBB8J+Itn9huRlG68hmxJv2fdYLArO9XWTzA/mIvKAd2zk
59pTxwdu8rNt1p84bCgJCkCcpiPhQotXA2QVduAdVngR7dnFqKgM6mT9l6dm3Ncv
Q1EkQAVMnSfj+Y8IlK5WcdB66wms77BRHETTTSiM5LCAww6y4u0tKtfc5qyjDWsL
tNIYxAp7gGtFvapFZOfU3G9JfIF3dqTBlmvZPEVrvk2bktFfsx+xCubZqdnuVLV+
jaHmqLyCWmvaR8UJwQRB0BMdkrypfEDzsLySUvABLGsQL5HuVB5rvADE+BrDadC5
ZcrnyJ25QnlJ49Jo9VfDRQvJ7r4U/527/3u4+wC5logRZlhUKwQugsJXsRVTy0fo
RE9zOARA6CGpK66AEaea9sIwDaxNWtthggFr4KSsXVNzZI5KaOCbRE/kxsCZX3hh
4MmHKFT6ea2CdS8H5QOXdFq2ifEWshUkDYu7jdiIMCwoZfzgeR7fGSGJ2Dx5+SCM
SZAyQnYW5+ciWmfwGu2H8/4oxlsa8SHQ1RdJRDNm43qUg5cXPvc80ktKUcBx5ops
+X6xfVQq6vjmyd4fxEXkOno65jXDeu4EKsgU225zeitL0hTLdp+kpPq+dE40DV0p
3v5oSFBIJy+mZQj8f3i4/FfNfDQ1aHTH+6ATvrti4b5VvrqWLEK7G18Oi3mfF8Lv
pLZS6YYfZIMICSKRo/9s7YbaMIbz4TLz1WbZMJO9B06lwXIfjCjwkMKynIdmW/JE
0tdrIZI16c72+KTHbFXJw4mEUn49KiBR2OD20jt62ov2Ll+LjurcblkA6JOLpS32
4HrirlVB7Mslzwj4bSyiLHPH9w1/8twv6iyYn+8GYmrdxnjq68ADbmOjES7AYwx0
lwhu4Xc4o6bytj3qla0X1nik2qgkydd7xtdfvN45Slfh8EzE4ro1ZviQvOQgv0To
1hthgpt2iMXoMdjhQltstiz32dzmq7NscnN9AeE3DrosoDUr7bAUEV/P6PyXmZGX
FfYkV3OBWYh0vSPYE8yTjzXODWcb/n3F0qsVMUiD+ef5aEVZT7lK2G3vu29CozvZ
M/KeDwcpmqVO3bB9vLCzk3OvwjtELqYlXMI3+fiT63rFD8i46ZrbdzoSrdBMKtG4
flIqQFuYl3ESwRKQ3J21zns4gM64cT0q4vTzXkB+45OcsfMzh20W2NHH2E+GQFOv
SZiiLaQTkEJjRBHQwwBu+xM3CccuFsMcaoaErtDTERhsB+14xlE91z1ks8ox4hRM
Gy9AfDCanRp4UGKLEgOZSdY5noHfwjyCuMpKO5riGaskPWG3l3gOd7prQx7/IjhJ
X1uapD7DZrLOkTs+IIY4XoFczedcDUN/JBEm3spLIYN+UTlaMeqoXpD4/2ddNjil
pvf+jeAf2QVLZsqHj1dXsSgx2o8s+sy5KVQbO09PsN13f7obIjALGmJScBZ/CTc+
GSKFhTign0OVxKFL+aDPIWYwu+Op+I+avOGEimxNvCkw0V1CnxYXS3czDResc5ki
qKlCZsaj8IHziu8AqhEexcjMgQcfckum3lj/rsYdZUzFOkHDxVeBuAIcrxHLtnB8
ub8YXQpwXMsHjVtj+0io6lM8Z8+zglzrLXerIyny8jwBmIzqrdS/daNsDalfBNJ7
b6crZ8Z61wU36jSNC/GpJhgYdamlErOUcrntNA7XS9Iv8w21ed/a0gJi1tRszy73
DIu9EfjsQ0rpa2w0qIahKoA9Ktn3MC9jBGOZoSKPwTyVQ89UZc52gwH4qBPJcrfP
9j/AKL48aJ/2FkV4i+oR+34zijrF63zU3UW5kufT2FjMj8R21v6SWTYA78OiVbIc
y49il6Sw19omodhih72ZyAqEHq/hRbh2WVs5CI3Pq0nnRcYTquX1pUOf2JpwMvJJ
TQuf++XpkT5GgMRcjXVpBlVIuGWgxohmn8TxJaZsUG7ikvfo4Qez0TpQcxh40yYW
hVE7XRQoAYB13VT/jQ1xCtqy2XoTxkfoHg08B5xRul3k8jfnOpAINwRdUKYWfWWS
S3vREXasQA2UaBNnvypJOnSC3fA24DUC8IvjG9gxFInxsa+pZ4rVFdvl9ti4sEff
AavPMxAqM994YILe44u564OHzZ7msarG+mpD9hM437oU+V1CO6vuaglGWU+4CuxS
BikQmBp0p+6YpUT6D9ih2FOfOwvR95NzcEWRJQ1SgLemsaI0xa8+i06RmvYIG7wx
eL3QQGdoW9S4hrqO3Iqdk1kJoVsqE0RspQ46CfQOG82JeXXW911rX21T+C2yNNsD
HEUZ07DH8jE5eec2XM/ZAyMuvedex+T5EScFUWTP8RiK0RTs6SQPtSu0E4NQ5lu7
wpe6I5sR4AMECktYslZttveMUDMGpTGH9uSVIsDkqIGFXgVUu6Tq0y1Fv1pnVvQm
vc/PAaY7Fj2gbfhIZ6oBNdyf0hzmmGhzXTOmdbkxlapWbH3oS0O86NdLegAvKI2T
xVw/gJEouEB8Db0yOZDAUP3S/IqN5Z3BVOjnRQeai903ZccisHu2mQ1qXdLaqt7g
mwtwY8LlfNVVCHeUEMMSfMAosFIoDvSlDhKcxaMVUshW5af4Ip8lQHrlRtViqeKs
otvlXQLXGclbpMwcFd52IFAAnsIYI9H+41npVugy6i8jh32+XCIA0q3ljZZBPJ9x
xMd/CFaGUqmPBaxlGCW0hgLem7bBn3X6tMSDxSu2jIbisu1RPJhnT3EMzsSq4DNO
nKy61B3G+BoWYfwUtHwHzYOcqO37Kbhl+A5ulyEtiZ5oV+CGZmJRJ6aENw/XKQae
7gO8vB7qQI9f2X9PFrM3ageqVi1+ZYwshstuBlRcv3vTayQuXJ2iSN1DQt3QD/iL
AZYuC/aLCZW8N0MmgjMSO4eCWBsThB4O8DCpHLjVmBZBJrd7I0AMnRzQcII+3z3p
bdnTBspXfyM17yUsHZcF9YWHlr5Y9U8vJ2ONK4ubpRyRJF6Jo+W64q1U1pZNBAWl
N/J+6jCML7Qmm4nulUkZryh6bg5gMoSlbivGioYCvaNR67CkPusBwdbGduu5RLNG
yw2ui1inPX3W8XhO4b0kx/fIoe7PxVqwqepcr7Md3jc3P1c1SUwI8KYoSUCqWFqd
ZoLqgLnR1K3vPV6kmDVCWk7qZ+8eGwGHInSwtxQ80IEp8WGFdvsR8vGjqE4TsQXY
KCOwpOe+wtuRj8WnxnCNaQK1E3SSHI7sSifkANvfyvSYpl8SQTZmZ4ofC5/YB/Y7
dah4xfotPSigicaMvK1zsUZmaXzF6feiWbUPFY7OIMG4Bm7qOMNG9d+c7Z3y6mzd
/0QZPXWHjbys3EOcBDIkuq7hD2Jz58LViDJpCzUSi6SFK5Yik7Y2GBx9uvxAGFkW
nzV1OJcxoP2PHVJY91c+4ZQRg4lLe7zJLXbDT/CmDvdMv7MTT1IP6nmuAB12lmVk
oymxuHdZlBWQfxALfTK2d8b0aGMFTXVp0FNOZy5mcCVJCP6hPjw6fRKpPzhBBC21
m1xDMJd6x2WLst2WenxJMLTQQ5tKjq3T5jfC9s7ciSYq8S0l933U7p664IBxZTUp
G+S1dYaS7wSJOXWNFLHmSw8tLhtAzr5R0b3DxFa0FKdroP0ElJioTFhNFb7+FAQU
+yWuRXmDMOOvY01rFFKfUpqY8I4mj9nBhEUqieNVlcWid7Z8pH8o6lxz+/qlJ9Q2
qstd3z2V2Sg+16kK1cLDWPiJZWf+BZwHrs1UWE6kW5Bwtd5WjJCy+qYn9m4sGIHt
Q7EXDckxjmQDttKNw0zMoXrVa2pvJvzQj6Z3qIKZGX0Mj6ojjjCBZtEPrdLcjsF3
PlNJllK4WvWhidIGeZ4UwhX4Vami9uYOxDLTncoq3kNNLmQHZ5UR4McHaUDP04oV
rP0IcSi/R9E/xrjV44wIxY8OK8DCT7B/UFHA5l7OBe90D30Aw1pAmaM+t6mW4ICd
NeY1WZLkcVQy41CY/VjFpeWBYQFSw3tEEA/Kw6Vb/eXDdRNWHG5fEHJV3+OdKisy
MPtVYQkfbkMm6O/aKezK2vYrftLcjnvxs+ykRdjVpHDwRJu7gI0oCNkR8xK1zBB/
eI8Kb+PXUUeigTqom1jmNkB1HYu3KuJYt/63jJqGkJDHHwAt2JgrEEvwA8+YmYaF
LVdhFORls2OzfClCGtY9ooXKiq2DKkmLnHUA/3+dMJfU0YbGIs4LhFc4vK9cxF80
Kekx372R66iPtS3g427Rg9tXePY2dK5+zYRSaMGUxcXFkOMDQM9VbbvBfK8lKgOR
oBDGLKJQN5QkSBXtdLG3hQqQxonNPLn46V5qGiKYV3gKO5NdBOdRdXozLzZ/gXUQ
DCm6/Uh2ZEHce/yST+wpN+NKazBmzj6lNK+5zCt6C6Z/vb0PddcuUoIL7P/HwY3Y
ujX6GXepxyaEsOIjILWFs2sE4vES/SyHSwxZhbZfHlE8FPfy+ok+x3D58XfYKZFT
jAYHITaiw3EbyPNE4nokdfZRcSzKvdD8bbZhXtn0UdU9likEfdeoZKrUuCA4Ennr
LhFiGsrxC/gHFsq0ex11ujrWqIAV7lqjJZv9UPmmNReEehm9MKDwtv5lGtgHrlLZ
CTQqR+rNtW11eGfc7XwNyLISh9Tv5E/83JgTFARQt+Inh1uBILMAvrFvtQQ3H6ft
Nr6BrRoSRVJ0BRVVu42YZlzNRv0vjNoOyoGkc4ot37ai/PKhWARb9ZgZ5JpT9NAm
4A83gu7bZZlzK4gGVjMsH8SVYUU6Dh0mzKbx5/EZhpTrFuIItqzJ4dn5Ysvk1O3e
yOPBH1oYyXa7yRpShpBH2m+R+qrDuBBqRXKDUh8PIxUqbWqPytC6PEETvHeVVbcb
DMwaTfsDGgVrhZhqmRhRmM75zi/JrfV7yJMeVMqnSI8oYymr1xzctRFSjljRCOpI
5Iok3d5Y56Y11N+DIfT2xMkJsdGeNpQ9iRcoq7cSBQizqFk+dG0TwsYqMn/X4XKl
U69KbnQ4A2GWsqJwEufPJxkBgBJ2XciqOgZKNWsBv0HUOSoHuHzkFK5wj02woyUZ
hJ+D71ARNyIxFCiUp/2Sv604uQHf3YX5rLAmSNVEdeEtGYBmIanwySFBwnxCLQpg
dtD68y/myJfFdr7mUqx9Yay4wocrB0+CxjbqjSIm46w4F3Y0vRMH4U1nIj4OMq9+
g/T7XO85+/nDOd2MO4ZP4zvX5VHwMKXXsRtCAXJZLAjxZ5facRo0xgNVTJ0/pM9Y
3CNSwWWdt2V0/0kjw0Mztuf6fwGKAR/zkBvLu3gkK+TVCuIA/gT4NjrIv8TDbONG
T/keqpPNVlq1BVgtIgmMfVcqu/deUyGhbUHDqzaNqjE/knWvSnbV4c5RHW62peDB
D1815SA9i6m/iWKQZV55qRNOjcIWJESwhSxh/jvniYJ67EXwFPmFOAg5fRfmIXwE
UBBKCgDy3jU0QtSDnam4D5aVnfgMvwclM8Zc/USc2I94NE1v9f3JtztrfbtmMrBI
sp7uB07+m3VHdNdRzRZoldckLGHeryIJFdLPAqJE0WGe5eGybsX6JOqRaMXV+C/J
u+4e1kcZ8YrrPe89t1+RjHxlu5VSRFCSBnr2j9qu/+SrkM5MClf4kLaX79omVpew
RjEZSUBRFt12+uP81ICbKNNTyCHofjZ24w/UJJ8Psz4M3aJfv3xdc3RPNef5vmft
5ZMoRmfgZSnSj5pDpy8HsGNJiBvsQxbobKA/izR/CcAJYths2lllnhfKf22oHlK7
PG2fyjdstYVsSCabMpxRm+4Z8e+PaniYUxpMUlDhzAmjTxJSNFtdf29Grdpu4BzF
4QuDDMCatgZpp2uoWMfaT0ZPt0yZRQkGZheUlSDbxkKWzVgA47dleh2EbbRcMKD2
15bGLMo3iznEuJou5I5/Vu9tztjwxvZ6jMJ/HRZIEibM2rxVTzRL9NbaGU/WMXIg
yF+SSMGiewa8+mZtLVZhkuYxFzUsNGhB3T9fw7OLwI+rb1DE6Bh0VWyN0ZNUBnO4
HKeDI2Y2+47sxGHvwIXS2hO2tcV/JLfOm3T9eXBHUaAlLdzCFA5TXNO7CsFp9Xze
z9Xc8YFk6dDProJsS1zB98nbvxLlRO87mKsDLDmzmmsTZ8G8046ss7YOA6w/Je7G
o9hrWEBEAKbPh9KFQIyNqrBEDqUchBaiIKJH0Fx8G0ja3Q/IsWgBbIYAvLrx6lJr
SLKv29rNnCwmSjwiTKTX99LDF+FfXGlM10JyvCC34VlNxaiLd3mTvxHdyq8lL1Ro
zJTa2BJHa0SPzbGHi5V6CUD5gAPZoaR2jtgtoTqnGmuuZWQijy2DX3FCsetecoW0
agHBUYE4vlGD37NwNEorSnMsX6FNMpkO39C03ddboPHTUd+tYNMwzhAmg40uILXv
I8/7lvMaewc/EvHgN9sSpzJhlsIAazC1vnMyCsD7gjlEegNpFr/9s5yT4mrlr66T
/xEFMtABm3n5hz7C2PA8vy5vdo8BlfiiMMNsG6lAuUDmrLSEkq6NABUr3JvwVMKG
PPc592gRrEEjY70H40EMadkTVPhrWNeh10F20C787jalRP+UHJwnAyX6Jv1frnH6
zibKBG27xvdqxmtWuhyVbSXasi3Kvw569AgjTnjF01S0FeCN2vaXFhWOdgmO+9Pk
WoBhzr7bRlZrs6AKu2FK5UGExNkOk89w5sl3xpa70QoG11EyA41LaQN36ywo8Pyg
e9Mhzvsc32Kf8cNxKRhSj0/q7x+0okB11wcf0S3Jjw6DaySF0NXeJ9xQKei2odVg
loRoMt7vX5IiGDWuK/ReoSDvVUAQaGskymwTxGa9fGfGAKPXcjGG/sqygtUH0kV2
H/0gGusCYq/+UfRylXzXs/ZfS9XnPpUpP2fu0AwflK+XPKlSDJW1wjsS+OZ0scN4
T7aCQwopaDs2qd+Cg1jTZqk0JL532X3MFWLoHvTR4dHODl2fWiUDFtsVnIF/DCSc
qFtwlty8GsB5siVOl6bgxfkshybkqhkYK6UD3HhjOPPSYIob8tctyXj94tWMB2ah
K2hbYFBfaX9BzV15Xo31deMRYzkD+e9qNiGHC5xqvBafvNg+zmjqfAIMr2tjQdnN
6gcv07wCArra+80VFcq24s1U5qeOEC3YYuoYm+u8A/hQZornS2Ia0WOxXzerTxYG
vOe2XQ3e+Q3iL2YIoTT79HCKY/eNg1s5zbniW+/FJziq0KZ9XevJz5SvVfQU78f/
r/gubSeYV2rFLLJ+q24S/hIActkFEqC7haWcAnmBvOtomPXgWcQM8HNczAwrbNYG
nieoACyP7FYOBlX91LyM9g3Q6JgCSjZkKUBHHA9V6b/URGF4nE9PB/j3HPhhXV4f
Zi11yJzeWwMCQhdmHAUfYZhKBU+VHuIrh0gZbPe+iACdN67E8O4+SmUqRNevt2Ms
KTgCHYVwgs57My0QToRDNIrKH0fjOqQO8AEL6Ju2P206++WMIBZak+m/aDSZgV1N
nrH1+1XTC61+MGfeTKiVegdV31FgvgfzKPTUNkwgKuMrfa9kkadn9SpYrq9A/vZJ
4FJuI+NZrAL+/TKZ/FRruINflslUkWCOLc7BU9Ndues89yb3jLWhKLlTAuYdrCsp
4ufezwXXaOPP8ZxzcbCP36+lwmU6erhWU7XGcsHL05MAoGnI7vO4zOscC2k4r6CN
Q/pFEsqM8A53cHvvC1yfFIkU1o9Y8cm35CsYACpr1mZcXfp2060Jp46hSOqDF4/T
j0NpYK8i7GOLlElMxL3tiqxtLIwAZi+9gaTC5/b5zD1+PK6oAtv0e1hCbcQ1QhQo
0UZeG2+K3FGcMu7cZa6A4+x76f1wZkVw/6uyi0DGtwjT+CyeGTcDyV0r3tvkIlsw
xuQPgpSwnQumwuj1IZxad3Ugugi+PtVivdUQaW2Gux/YSwzgt5hoGam6Vyje0qeP
fgz3eMFa+QsCfjgYT5OP+h2a6fvYa3j37QFkj1iK+UTLdlwTHcYUGhEKonld+MqV
W9ZWBCAzrKd1QXW2nW6p/ZRD5n/GelIT8D/DbBKxs6W6UV7BNxGGv0zCV+nOsUUu
Qev/mjPVVyrOMmyoOcffm2cKFuBhFuQQCRkp5aBAfhJCkrzyqPTUCBEJuRaiUtnD
UiHEYwOcSbLnf6NFZdlaqDv29R0wvGOWaQ0lyuX5mkcxNZPF6VyLqbSVHcm74U9E
txPP3xSPFuBCqMei+LGDA5CIDoKPWzZCyVWjvQZQk8fd0OzQH2ZvCCxNIBZtzUVF
lVmNar78EnSKbZOtxLCHSoUNi1P4hGHUxSwYwNtoksuC1FAOpNrHdLRgO0FjaLUD
Bu4ugjaV3gIZUBhxtJlpMBHjexRbY59mGGmX+AECqkEn7Zgn0Cej2uhpDD0I2uB6
EAbCTavCzNfLnKIUDoOw7lCdOiWkZoBiZzqfhkJE616kWit2t60AKg93C8STP5uX
LV+w/LEsGQPg4EPfBQidje2jMIxHheQQRE4keROf8RAMGjYbnbbaiD/HKcRd+B9J
mroPSMHVVckFOxA2yNsJ6y9GzoFRiNB+MQLJdgx0xDgSHZ0Bfs0NH0S/8eTgSRyo
2wlnZDLyQuXx3BksNFD4Ois2ZextRdDED5iP3qOYmlFKkWW8mORQD54dM/Yb9Xxi
fNPYh8Gh93ocZ1mk4M1u9NEPwKiinRUs7pdYrtWba3vWeDtxLZQsVOmidVmn0vD5
ZkCyoh5hNxgXrvJ7u08BrJek2QNRDoSO2Jr03Yd39NtFAMv/haM3KKRHKmzg2uSq
OWQcHnbF9Rp3kU6+xUeaHptQwEcCOk1yaBtsFgttAKsh1yzwqLextohFTJF3gUbg
BDSwwt0xPFNYGbNlnSESapGC+WWW7Jj9i0l6sIMIEwyF42IF+cSMxfq22MS9IAVi
kIUpq24Gi86bjkDP/P2FfHOV8yaa3TzJWxMQU6UBVvOY2Jpf+yCLvXqVMzIb66B4
9YJfm5nQnLLwgf291rAocmZyKgpbzPKTbvW3bcI0Qojvi9s7tznwYiIf2u3cuk7i
u4/W0OQqxIYpGEXaNw4FNx3QC2+LU1F/xyrcOSKnXRMsYXLF53oddFAa/8QCpCzI
4qDj9TIsPteCHtaTZM4n1nWIlq2lic0PRN5HLU21UcfSCMzd/Wq6PVpRSPAT/jHC
+hc9r0Cve61KqkX4zwWsl+6/7MmPMJlHPcyEH9kTbHkku0OybI/fiQvPB8+b/HkG
yKzktr9BlXkiTLh6YO09/4XOZqR37hNf9yVb71sG1gR3Kd9039PaGR1z87lnyoTS
oUO3F2aJOWhhRPDg+esF4om2Drc670aPGlYBk5A5mciiSIxX6aeYvi2PwCEc6POR
f9VZs7dtqK+zHX0+Q689hEfUawvWHsvxPAFiIpk5NXIium7ieBn+ADNGnNnS2PD7
ktLOfuKQceu5w1Z5cByesB9ueohXrnJ+UZLPQERmG7MHgB1XEjbkjSQGVPBBuaeM
XX86oSxZsIxfwoYLwWh0jTF9rGtBXhP2NKL1/h1XGjRosNAkCTKgWHoXVQLbUGkY
jfCzhrmAGS3wwG1O3z/nyBoI5xFLt7ltXoB59FxeVOM5U7j3kU4R9SGgYcPJAavF
EjydpKTuCyA7GvDSzW2qMH8YwcbyMWufDVd1m7DMuM0AOxWkp8mwg1QUJksimVJH
Aqm4Wr2uKtLvucZAqIpcw4Fuj+wGOPRDjuaAmqEobYp5+oAcs8eIR4LqTRL2Hosd
eJUlq4G/cAaG/OdsPSabcDwbqaRBSY/wCQ91Yi26RjdgN8gYHRAYj9xhjYfE2tY7
zNUCrBrUW/cmbTWJdg0M7FgKFRQz/NdCkW+xRYxSgiPgPktF7K6tSmO1w4Dxy9KA
GDr6tLBZENM3Joce+5JPA9TSGCAHOaceOof8pPP3yJdSMDp5fGdbV6tx35BJbClO
sEUj3pWnVSxs5XMcqRSrUjTr70qWyonqED9bKCHKhoiX8k0PHT1Op6Cc7LJrEG4z
0XfyE9/hncRM+LQM3hMVMI6A9cmQs9Siaz4QtPEpsjvXFjxU4G60cvi0F89KxiHp
AZs2OCz5dtzx/CRMsP0WO7Do0q1r0ceegkg/8Fpzl7+aaiHA328JmQdQNY6aOvoq
VGZeLV2dC+HiPs2/vLGPKwO+wVfpw8r7bOlBZAu/5R3NPmkXcc0TPn2nXrWQZXRy
XWAm6EL1/W+ZEyAT6KOIwatXxrjnefGyZmBQw50uSp3w7L4nEGDyAi3VcFdHMbMg
kDa9XfQadZH49jBPcdXImNL3WseeO17PXSPLFl5108/Sb6sGW87v14akPAj4qAFl
5PlgyMRi1SzyQkFegsoQ10HlUwul6P5g4uFL1VXDBZW1GYId7GDblFhkPjKhUVvx
NWKYCg7hPqyM4cTWHDvhFpC6TVOc/s6PKA0j+PZrivSeYX9ZClO9Tj1C71jc9dbS
aRUNVinXnke/RD+kQIFrq1NJScVVhrkMcjYiknmeSO8rUMEFh/ACi/vo6wEgG8oG
ioMr0qF0NKsgbsWL8F/tMA17JSkCi317hsgNvFGgys4p+pPSMkYcUur4jCPfTqq3
AwAsNDE/F3zEtK8CF8YawBec4oozmASTXalS5v5yNttXCoNVnUXf6mRsSeqZsd8y
7SCD9EBT9GUsJxcway/tJUwTm6aDGRbp1kJ/CSbN3fzhvVq9ygEiWZQwQemgz162
O/RFDBvfaKEZDCpAbDjVRtCw6OiMao5TCosAj+iI8z0YptZXdRHZPodEBp5q7fSZ
WT/eOUTw8S0//ZGPEz1DRShsFMPNJc/MWeta7q0dWzlw0y7T58ThfMjsNJ6jg/Tm
WChG3M2O47mSD6WBCWJYEm2bynWxp07sC/ftvvu93GKdCyqiJZWA41VEOP3S+Zg5
9oDjICCd0DuYZ+wjWpvCLWOJC9RiSz88Lnf6EkCqAL0kJmTpQyoxApRTnYWMZqfH
L6b4OfK28pyuVLB/8sbhmBlTXdEJ47MBb9ertUutqj/z9ElRM4vQyNUVWkqMAm2j
z596kSFCNoIOOdKy04xp1aQN84mazeIC1tirzqSD14Q0gXeJiTeWvvnhbOW9FHtA
VHFS1UCZir2TTtR5D2OLyT4YpicIWBhPpx8HhnzomW/0EpbUbBeUIJ2qS1sgWjCM
RVR6XbQ6Z9RfVhIn2ZylAHyKBrVhpIrCBs/Qb5PBa13W9LynDd2Ri+D/OdOZTZAM
6Pmrh43V0rp0KTDp7hH0NKqIvtX5UCSX7eVh7OJ/EowLwQuoAw7stxg7kRl9nPi4
Xa1LrZGfbKL78E3NP0q2Ft++O7/VtRBmbgc/76us94v+FZrs+D1oKFG4LdqPg6D2
l8v/qglDgaUVSCdybjYoW1f1qXLJdk/L29O3NF0xGfrmE1GQxkeaoms+VXRVONUX
Ca8MOqbkDzncfyfJpk6nUwgDlQ3PUOwUFncxZbFgwTJQ6lmK3Zz62vcEp+HfZUmk
57Adfo71QnSFQoGPXh8gqgC5OnH3dscz83q+ge8DE7eQx0X7QiEKkt1M60WhaGaC
OuQ92cpFJJ58vXIHrSKi1QjNeuPgfWDLcNAKOu/L3yWYKvrrvQe4IzOs1YnVsDlB
g7iKQmkWj3PhqGt39QW7N3El8whdWMipz9FQ8ISbwo5FWqvh3T5XLgq7LHkpvG8h
+LOiS4XEEGuXr/5YAiKeB7AYbSBle6Tima5Y2LanRM/6eBXhcKIrCHsIV499xzbB
8EDhQm7XpB+yjLBcZfOHTnA9wq4bH5G9KFeMYSgCZkYahKi1uD837D/FphaibmcQ
OjKLxor4XzUdcXDKpaVEa5mLxv18bhDIjrSAZWHBF8Z1yfL9PW/cBzTi0oYwlJ5J
rtC2zQHTx92khjvX7cXvupFg6w7So6pAYhUeR7ZxoxbHn/VPdKsOTJFiEnV+P7mc
KS1ZDza+yPyGFKEhy1ivZ4tI+siNL4lHoUkYScVUcsBKrN2vOh1UQI2rEtk9hbZV
hy1IHLneR2fYgd3vt15gS0UKlYOksUUCwnioiG72+8cM2v1k2r60w2QiMrNNFdTd
Y4DG15bE5B+wZrRbHWmvcAAAr0i5ZxYjeRAtEHKReeA2xJhnKrL+ZxwFSl3zfeeN
Ow2Cy0zbKpa0eZomWxQfOpYKcQ/KKxSxSTlf15mJ91oSOciX4A6J9xMsIvs34exh
B653MyYlS94hxkKrG4JB0giV2dXjeoRB8r+lKuoeLht9HB1aUCjJfWPnQUQUHJLP
mSzVbc0GGn6LE1HowRfomYXTR4zj9pleRaW2MyDt0B06dh9gNRr+xB1L3e+R4/7K
QbiwVFL1IRvGSy5nnx7q1amX1LEWsu80Dq43HXZETB+RZe/gLjhiylRMczR4cWeW
nuvDWeDVnbI/bxpFZmHB/HZ9b+Lg7lKxZdzLTm6XsYXTWpfdmQw0CIekG/ivAPW8
V8ynfVzArpKNDkSRnM/R0L0K3T0fqPMUgtIPWL74QC4HPyPsfpMfDH2cIsmTHFdY
T4N9XJ1ZlQ6hUs354sZC65aTkKvTjjoajv9clf35Zd7+sGINzNvWyxRUpedGEGqr
QaF5cJjXzSbCJh52g7SG2zXVTe8SAUuPzRCd1ujkm9Hqle1vlhN3KvWIvDv9wcpR
YLTVO2wUYZSd5vw1Jm2mXFSXtwfv6SnoRZ/iUkX5M/q7PNLTfT9I7lCEYuFthAu2
oCm1ZS2w7oGEZmAmMA73Lc34EqpD5d2BRKkKZiosYhwK1dEvXOfgSGq1nDSfsNa8
siLFtYdG9pWKUhgmSnVZOn1oOArdWNS0xHvk8D3GcPEfDzZzIZr0epYF19jZrLq4
XpY17sig3qUNySwh0CuFCTDIDMfydJ6oEplnTFHUq5BRqs5s5tgj/rkrWXGxT6y7
oqZVlV6te8aN90fLFhwbrNPOb2EwMq1BT/cmfJuFEhi+VZUkTFiXuaTVhqVXxW3f
Uig2il5yB1FXM5SCq28IqP1vcCPXzEr77ShwpCNt3+QdLUnLXOhc54y2sssDbIxw
x262mTu7yE5TZsAcKtGePmvLLLlKvVPA2yYdccE7tik/UVxBExAN0BDM+MTANrML
6uRHQDkyy8BsyoO4wCe1DJiu06L2mow40FEbj05c+P1Ier7hrHu72w66zMEdKSW/
h1O+7v45aX8UXvcDpvJT/yjYLes+cumW3uz1bQaD8aH5KDLpd/+gY6jgkwXgg9b1
nnSIf5Ig14EgMEF7YvmmkncTkV8TSRo2cvCMCxWOkMApI1a6+JEa82+r4oEJFE3a
CaRub8/p6BEwPRho3eunZQNqii//4TyaquMW3lsaY5SNABsPBVkTZ2oXABAjnX+Z
GXhPjUlB6LGzLc4CQcz7PVxf55B38Td+Ba3x9yWncFCz8X6SjbA/TfUaqOCYDI77
15HQnYqQzNOlnlnDBSSCUmtPr/Jxwu+I2iLssYurQTaJ1vw14kBLxD7S5z6S54VH
1E4a4aZLBHgJt2GRhuoyBj9dJ7GowE/H4STgRHsAC/TP2c/CaUiQpnS70maTABaU
k+yqIGj5oE93DgwegEkWfywtHLk9p5vnszg12aJJfxLEmpgx1xevsKdZp5W7W4CC
p8N5LfWgu46hGzDw+gyhoQ3ipktvGgB2Acak1CC5zoWtB/+M24jGfNXRBf755qG7
INVwpgQFCDZ80d7MMZXoNRh985exgAgYLGYKJ+t7x/1rSvMDoyr2VSNDTg4jmxR5
Jul8cLgTkYkohvcJMQ8vxedmM48hETuEUQUJqhg3KJKkArzbhVO+V9L+sRcFS/DN
zJQSU1kat7TtMby4MfE6M/91xRx8Hm5w5BYFJkVXWImJybcHCNB10xCqdL9rpbni
QoUsvCAWSfgtFohj9PH+CR0yrC9BoBJ2miZOJkAHC3jEZjjHmWXBrNWeNt5oYY2Q
6eQOKxytUlK9sKsxZOSQv0zpOW76/q/e2izERFx//W8KrOU8xODszu11cwqcJoJm
goB5KOeIwiDKh6zHX0BWLDI442OWrZeAG5Oeeo08EmC4VAXeVfXc+aeUzby3wCgO
hCCso5XiAQiIThgjDkBf23U047tcE9zrYfT4d5jlppw8d4nQg0gRfKTPcrL6zk23
xlVRJDbSro02YYNafoKLAH9IFORETiAh2Opq82IfYwtBwhc10EgtdVHKzHdIGTxJ
rauZm0R2XU2PliOFKLA1yGZ5qPm26k7APGfXXgq5JVxS4JW3eN+olW3BSWQM9lE6
Srz2P3dqeBUcHnbIbQK+9bGBJkh+MxOEA4atWk9pBJuNWxa67nc4Lx+GUlfVtZKx
eGHqIpo8fEva1EXz4oVxuylUtcX76So24OAr3D1Yyqg8CvMuNo+dNNXLvPpLRCsB
vuL7Se0CjuVJxilNlxCfRGjFn4+XsR1h+NbWfBN7Y6YzcHERm6yDPVZ9dCtQQz4m
tD4qKttgkbDrUfLuR9FcO37LLy4BhASWX/7uNh1VVArVJHH8dXtf2N37TAQRWHlS
mUyYe6u9sZQlGvhXe/Df/7YVc3MqBFQNcNJCOy9F5o/veiYgi1WI0TmMeWvqXGfh
Hddosmod0jfHagAz8FsbfWOEX4K8dh+Tt4D794b2trQAKiIaxz9cV2+Z+x3j7grJ
kHWcyLtKBBSuB5veZdWL+zLkQ5jnKXTrV7ZdnDJQW0wbW1vqwW/I3IH0Rjf77g1G
TAY/k4AUPbm2XTLrnD3BrbPp/WB/mI5inqlnYXr9EqeVglqWxVr7eLw55g9/rGQa
9o2nHSHZO98Gxq8pIx5/FFMlNtMiYuhJa3kjrE1MLnJsI6U+3DetvLm28QWGIqtP
8SxoXesBpHOZJ+IChsmxg/v3jRwdHMhR1rwjNdjv52LjE44C5/HzrGv7fZmGbqmZ
zZWbjzO7Mp1oXShv4zLZ6OSeXE5GI/loA8rP669T7GTsrwyCW5i3BDu6ytUDj2dy
W3toq5rx4meoQGrUT8a9OCqxly2AxdVU314ow3cyNTIZ8WhlEP4qNDZavUV9O58b
plcpbfpG4Xam67h1Sb6t49uV2sqRinGzElpQNX1mqbwekOxu+3K4pRFCnKe12RdC
Hh5tPNKbI8zi2/L6L9N7E4+awuGDozT3MBY+iSkx2z0P+AsEAiPm1X6+HzTpvm9I
M1s/9OYQF/GO5Ja0WkG8vqsOa+VlgRgt0ax2jTWWdA4v5Hs8+dOApt3dgIuDb17A
CVz23OHMyZIH1WQL3C67hjyrSjBiV3qlD7KpcVXHPCLMHO1OKyAaOvD9xHCWZWCe
ImpTR9e1L+R6er02Mn3cHcs5k43zM8GR4rf1hMBMRxRn+PHaSBOE+2U9UHpcFVRA
SmNLD7H8BNEFJlqbHao81RDfpCrRLNSVz0DLbv/pv9Q67YCxYoNCjTAJHHIJFwbq
0AYmffw9etEwHV0jiOC8eW0c4EXEcQcHiFZTeQkO1xlR0IgjffcizhDQuHrDZMKM
SUXFkcie8wTowRz5H5TyWgn3J6qFJrf/EEuMb8Ot5OjpEvzKumGVmRsVn74etZNF
KBKdPiuUWUG0bn2vmjoBxSp3C0/LprScToWkSBUN+eHcFs5Z5LVvWsXDhJLx7c8o
Wb7dxOMlEtCRW+dl+be6PhhPMhpJKetX57P2DG239rfL5PjP2lX/g1b7G2zGV9Vx
SpsO5H+VpuXoYF5eh2EtLKn6E536OhTQhldQD7iJOEs08JtJ9fC0+ZjmawziwYL/
w+q8EkLRWUIzAPeopOtCCQ2x8x197zH0TLxuJS29k4mBmr4T62wdya/QllPVNBhg
dmbdDOizmrsvA/Ni1cMVarweUL2514In9DFCWB5DS3dlQ9tv5LTk0+sPT+16L6Db
yCHbagL8pJSObHDmg7vPGoe6FotqrH4Gy5qFm6yeOvH9fPQ6A6rV4B/dcEW+ObkR
htckIVQaWOQ+PZ8qLiMw+i20VoAamqnzSAO7yjCQfTo15d/l/Keaq7fzKnIlPu2Z
kWhuImfTq8xz/My2XJB7n+91qRgpFINdNT0wGLMJbVH0PhNQbkCvHwmI1YaFcYq6
kCXIHV72oke8HstYtnwyY6tKcDWVzUchrW3j09GIpxbfsuYKPE4fFdCMKnqOoCLf
zi7v0MbaBT5YNWjEgR/gqTFuFfeIVa5LoiM9Xs4uRoIA1Or2sIfovSgoScfb2sa4
LPwH5HAkgIj/iK5hfpOnqt3QLYhh/E/BWM+GLPVjB7ABOh5C/ZCAS9FYsn6oSJWG
6/V6Msr5ho1az4ezLgK568aXPD3D5kyFAHWsbGXRmS6d9zK1E03Dh0YMVTIkn6rB
IxRnEht6jdZQV5bChj0zCqFc9QBoyrYP1GoVOkhS57Ejx/hfB9ky3GJcyhhLbbwn
XqyeQhArUYMxsNc8/mRtA5QTuH7OdV7A/tz3Chw4fEGnjsxgW6+4YcfK6mQOKhUT
wsEy9FvNP3GWSaes/Si4jwMxohwcqlmuvke4294xremRAMAvOmaX0B+nk08+V3DP
6F85dgfh/JqxM2XEyqO3QtCE/OAVhY006UCGcxuHGCOKl1KaTg/mRnvTXmpezEk5
iPBG+DJltretSfAYBF+o8XbsdFoRHoPl0T1xVhCkEQHXMTefhu98IruK+TL6YKA2
dWM9snnAPDHdeuY2OjZS9/EJpRt9v/yEHG/D92gHZeFTZIAsRikbYAWIi7NNOXO6
qUzYTil0H7lpvVPJfFGOwAbTVpqgRdHYBrfXC0PzQdIplM8oX7keJ8inCrG67hAs
DAgYZzkBhn73LtaIffyecyz6qIW0xv9+KcoqttpdNsMg5acgJnQBxRB0YGy+0GvO
SI9GtOkMXe+33SmnjBIvDo098ibcfytxFmzuxEmxdeebHAtTNBhMTJ+xY6Lh3sk3
T8oF5gHKlN+gBLFnC9KmerJm9a16q3F2x7FDwmXUJpmbx3HY15cWX9L0tnvu4YYH
bR2VH+/R/cucyZrovG4VvwqcKojbmWf/sAhv/XRZDqmLzv5U3ybZk/v+UrRBFiGO
0laU8tI/79hNovsG+LunpX9W8O/8kPRfBnkxDxb40eyGPlwalFTDC0SUkPSM5ZRD
XYrqTWulnOUcVX8EJrUFDJ80k65V0qCv42sUoQXWuzTREr/Q5qHhMTxqOkxOu+Ds
EHNPDAA5FxY6bFL4VD01/1oeoleBCBnzyVwZC/pDFGT5oguMLQoQ2RyAStQpF792
/ARWCBNxOh4kjkZlm7MMXwSol21mwwWCOHTN1roPvJMY0KtpubXP+BiDgDxIJNv/
aHXBhHqKkrYgxnYVrYSIcB7FpawG17rFs/KYpRNu4SD9hOB1AEMl/E1b24QWpsW1
8QYbqM55k6An5eC3UyOkfRbnA9fD/xBBVM/nG3mxIlqv1akn5vMuwM7fICCL6PYK
izqzfqmntSiKpXgBaIfV108HU7B7zs1wmIoqpQJnSi/krVPmJB7ITVS1mZQ3care
koWjWnUwn5gdwcGLNYcQeuLxEhr9yfalO1sdZMMRzLywCGomq9Mbdag1L8ezZbqK
goxPc4f5PBYWNskgzp1iuYmyGEpAxiNmFvTvww+f8DLyUZlvTTskP433/+bPvz57
0wqHW29fGmU+aOK/jIhmBiYGcDWelNP4wT9aOBMJu9OM12nyThp+5+nDctO6Jmgq
y8hf7yao5Tn9eS5t9W+Tu+xHlsSlIugSb7maDcFIj2naeQQgaD3Mya3i/idt9yTH
r5DQ5VyRq8HY5yS1fcPajlvz6A3PxwATdDAZzxKpMjTyRH5zKd358sfCcfTiRqYI
nZXfPJATq8D+JLuJNR2WS4RDkdy4Q/ej4BOD/387FrwWnb6tP9B6uM63r3eBHAqQ
0acUTnpjPqULtQWez1mAijF6/NjiwJpr7LApoIUd05ThXuWkidY1gk7cf80nvhgp
bGGYWsJX+zqXKO97bn1Vrh8BfspjBIMnvtr09qpuOwwwc1vBaQU0wYAOs/sfGYIO
5q1vx0V48APHukEznslLsfcPwwAFJjeGvTsdOPOm4yObi/OoY/mAXvhxfqWwXN+2
67HXCoMPZEFcgzel66F2R72qXpV7eBbab9y5WuebNCy7pVSlMDg0/FG9Bl/2x3ye
SH0OErqbFZohaxfBzxXkZAbbq1ITuJVzRJ+nGZMOdEB5zwSwbLCboaij2DfqCxeq
PTjdiNfW86hzpPmYaHLx0B6fJ0AZtyjIVTCiStsQ6OzWSD1NPQ9RQEgKsUE1ri98
6rFn0IlOLlIsX4fA+NNTbnRCvtDt4byGP95tgwQgMudZWnU1Nm6R+V8vl2V6xULq
RkMwRF9faxI1HFg7H2npgurBdFAscy6/4FGYBaa7MJys47jituTUuhnS7sULUfJy
YuKHFmIJudEwjNU+n/YLMVPsWkip/79HaFJp3LCLvmnefbiV3+QXV3nX6oMKJ7mO
YLrn10YnazJV+OjIi6Eaup7F6VFPzH34G0Cb0UtNAnEXwp10J5vZuy4vju5/7bxS
4mhqWJO59iHhYAfdHIbqc5CUE6/JPRuXWXfgO2An2TrBCbqHa3xkCPNfdYIkJb2e
R13Q7p/Ssk3LWuDu9q2Ro7UkbfBLwtRMTsxMTvL171ox8su5KbmGToCz6Og0rUtU
3mEspJ/tzKk2QqUx1vlDfjMkURqhmJ3WY/d2wob5XYKbF38fY5EzYSHB474tS2Q0
onMX+ZjMcvXAM/Govoji6VBViQ3fgco+kZ3SsNRN5IwuFKQmELcqtm+sumj/wkaT
juaNwDEIY9UrI2+YQmODz+7VdtxLGYz+wz6mU0KiBsmVjLgAZObjwwMl57bagWOC
to+wLNI9so+V04LuXxtt0Kf1m55m6tUNc9bNfAFmxaweAE9vKjWguFG9XkAIKBU4
WPyPg+U58+CmpNQHf4DpP305xxSE6wYELrU/KsEFWArW80AfoMxWlmcqyyf8+Whr
QcdPbunxv79l1Tihcp0pqp4G+dTQJWvfWIOc7bTJ9bminOKhEn1bpVykXiHyhlqs
lRGDnudvkikdpB/8yAKHrsLs3X9mmsVsTTmBwcVLnHbjC34Oui20AjHUovw28NZ1
NDUZYsrrxMg4YPCTeqHgJ6URv3ItT8Cmb8PCwi2JTRaYkXa6LSPzFnvjxPQg5+CS
rG+9PoGrayyFLkdBtFJCir9XvTVA5YBRcOFgkm9MdQzLNbIUb21+kaVhPr267xDn
IOzPXtt31Ih3hRwGX0CSC9jLedwHxtw6TKUjxw23Se6xSTJL4/x0aPfPGqAYj3iU
mHkNnj50GekpGj4JaTbGPmiclsmRi6u17W1CZGayNapO81/Nq2cdTOIkbZ0PiQ2n
AVa807RNMU9sm5WdfA6Q4+vjJND0YEtvRd7NTOr+A+6E42ZkWIDrlhFl4wbwdGdx
REkQaAeaXo+CCSykT4lqV5aK8c90u2Gkh4TW/dNJO8XyNZXW2nRxHz+MMNiTX6n9
2njlajPl6YEtMkXZgrq5UEFM7xkfXyRI+/A1X5CX9ypwXsXI4fB1EBQ3M/CKVmnT
RYC4onvBDMu9B3PYEPxxwOhD94CFkoLaUDjmoMMutbloQXNgND+zj3IdY4D1wpyf
QK2ykQganqnEAnEEhqYhBbrjdzeYXK682PIoUMxOjhtpL0RGIo/FnfOlUk0V+JkL
s/ZxwGEF4SRtHQZDz45FODwX+L1d3Wz+fRVU0Zw5WzRI+LnhCL1RflpUJ7PuNwtl
nf8OLlLZjkreN/6Kg0qUiio6qcCeX89kXXACECT+NUwtboJ0d9tekOdUH/Tp7ihx
TIBWHcT/clJy3/05z1qJ5b7e1oV7qK0nkuMERDbxDEar+voA1nzMb5IfSKvHLjzM
0rh2Doax79SPhLCfjejJNAwUbg/OrzHimu9ixy5sgAl46pWRhkpUDRRvFx0XUQ3O
QKrDEsrukcKjFtqk5XZsa+kbfUjatt6+Pg8U16huBeWS7HZiGEibt8ogZL9r4sl0
i1Tv+2pw9GvYI3J3bIhTfu5JbbfcPeED9CVTgI6LGypiXE+3tjm3tzY4Mu2/UIbq
3EDVmcsGiMP9wt/ZADfyiR687IPsC0ZIPhC33rDtWXaByEvMIOsOlLUUN4gGAzT4
IN2rDqkAqEPgerV/flEv5A9aN/BdXi3J2eGVviOR/Pmrix7A9ZjAzbg1jnZrYFNA
nNVDvltmor9lPOMcP8FxUTMFaYbTJCvf2+coPxazpO2iladJ58Ib/jRPCRoOl2ML
t8CVy54gbHwV5MytQgDkSdmmpSDrO9jY+Vv7/QrknFYq4zQt7HaFXi3LjpxT0wGj
xhBRnjL2CXHF8KwSrmd+CbIiicuMPyORA9LNaqK3XvbqRhotuWVsZe2VafHhWRw3
J3vsFK7ZB7Jno84aGIe33XRW4VD35VaZw9HvGnwf2m/4A9XjispwvVJ2feO3LLOE
P9tlBemzevJieLYBAXZwXLftAuxkp1XusejWO15D5HO3y7vYozXDSR7u8Ke8FLok
vbWqV4x+SaQEXaNfQhLpDMlPCYJtF2ZzUclQAnUhiD2KEZRWj0Hv51jdi21OifN8
XgNThjIL/3Ot7Y2X4Hu1mOiTEWkU1vM7HZLas96wMaU3x0UsxNEOoHj2c6iw8K/Y
x+xRQUxi6ZJDoZDurXlm37WtK/tNSRp4Uqj3wepYgYXYoFQ2vpNlyleklIojOsrS
wu/rrfDEkpdJVU8d3e6q+dR6Arcfn8sWZvpt17lRnK87Z+D1Fwzf4VLsYFH0FNHR
ZyfezjKIDFUlfrTKhS9eYqT+Yr1Ftq36e8GHj4197Jhl8LxoeGDZo1Se0OrlHg9G
h6vydyh+fVX360KDtwboEQ3f48JA6VcIiGXyUlnqP1giqg01fmBphc8MNxzx7i5g
9LL3fz0O/iXf7tkCAJkD5p3zNBGnI1/xzoKn+k5bpGoCNDR7aG3vB+XATnr6SvR+
XdZy274yajorlfwDqeADkfWsFKYzOGlhSqGp68QCco1x+kqY2RFCRxj8dD8iNqfa
hMDfhQSFRUbbImzwLOUpompbhvh7DGl95/1o9uuFz5/LLH6rSKyUzoq+2ZhsuDw7
C24a36hC6d28vxZoMSrttn8CJ6/KlIl6RKh5JmpSW32srdnAMcfE5Ygy0SFfHcWW
LhvoJ7ydhXqh4sYXd119UYHEzDCPbeYpHdY9PtRYVXtdxFznxYOFv3TVA14YFLWH
imPXXSvjSNcoDJhpXeABQptDeX1AakI7pfVorYeO/MvnfeJrIv+TJkd6vACyqTeU
8rXoYY8PlNWvaZ2qfhjj83/yDjIAVSv3j1SxSNV0ZGFaFdj77dGAn/pTqUTGwkdo
uqwVOPSZwCbZA94t1ewrhEYv12JB2FCgI1yqtgcq59aLoY6L4EtQVaKuTkruSW7u
+9GMOzGCXlEfI+E7Ao0A390GqsJk0ibc5AXldM26x5QeY0D+a15m/RGLE92+p6ni
oIWxkYwZlLF509nbRb5Up5MRwD0gLLclLUghRsZNaucBOaUaJkiDI/7G+Ufhbwma
mdffF22NjD++j8fsD1Ih4xpBPuvk7UOPFBR8+PLZYw8BBRJv72NVBr7yC3BR4q3g
ASUbbjhkLtOIIGgER39kU6z6SA6rPRPY1h6PkgssXudJ5MytLpMm1uGOlgeaJj8F
0ZBrbOhT0yW6B76EV7nZ17pktHQ60l7/ULznHdYEa5aFJZSd//izDCTia5+o/BEd
p5uNTVivTMIHvq/h2Dz5XUeqo/lAxjpa+n6cWnVeS8OcF6SrciGQBtc/M1d9n8Jj
3+HU2xjioiyYWZtRH6fucXcPbmaTMfaFLFrQO/VixYcR3P8HDRiTX5zbn0md64Qk
JeTx7xh2x1oHO0rrHJOKSFkgWeBokpby8XJ49UVUpKngbKFn8pwKtqndbPXsSPhS
jZQSPNoZ6onZAYtE1dokISRCnizt7ecvPNM0t236MpU9YErkTfIPt2a7Ta51v+vD
MwE7hZ0sxmRz3zA8Rv1ZoQ15fMv0Ktf21QCyLUTUHc7bxobKAMEFpaL5MHqCIlcJ
lM4BApaGZOW/mThopFZhLvndifYg51PVp/BM6aN6ZMY+mn1eV5MQAlNky5e6TBaX
/lAVKHvW6GNBePKSm4Hdmz7M7S0XftjATIH5EoOHnYJP9lK4vQN+RafUSdtWFSBr
KJntWbKav/2G3ozIJxswlub1XrG4ppQFejJJi5F4plFfhiq+Kjd1UtPnNIir7S5k
LO9kbDCTZROccKjsIThyLJDwZ6eqnEmm4d3+O/EVKUtgC93iTqyqhvbZ6vf52JFu
IX1VsXJ0IzxFks3z2rdP4g1xhOrBR3TxbBE9L5LJ83BdzCXn+58v6QR+l0zzXiV0
72kRpcbzqpBAPVrLKt646blmWNfZ2NqQ+mrmkPMcbhJjETazr4ar0q9ep2nyAM9t
mxNSJEsJxQviizveZgZngpphNhoFjVGG94cUomA5bvSnIbgAIOGsULzrAcOOdfrt
XOH9c6gyDCERlSGr8uj1I8qXJPggBUtBEH8mt16lzRCdvA9g8mxUhkSe5xWFDRMM
VPt/MpZbCUKyCV4AGlBNphWsAG/p3S/ZqyncZLB/RPW9bTZAeXfBTFox6QaN11Lc
dgojuAAvS5A8zYHFd+TWrI9uldztJbZdj5TUD3sdEbjnciEQ8ZFdiFNg0v8YTzuy
YnUeCwPKKzdM7nGbVUKeeh4WogbGefMznqH9X2gtaJZ5svIp+4xngORQJV3MWEXL
/1L8/xup/KOgmwZaSVLTRhLrX4xscbeBVoxmIcezTSzQCYLWEhdXWEhNijLAaJwJ
FbQtlMmOkv/Cqg2LSHRtZgnU3B/IJxC5/hrqHthyk/8PzFSs0w/QYvzx4N58sHmX
5EedquAKonacKBZHEuGPkO/ziJxv/lfBPP9foQ15fhp8XF4gBXQ7CeGE1a99g7XI
WrdGh6fnB38A53xihotaPQpdG87KXkdVkI9BkgFEXwvc614Q8cmHLpwzwAQcShf7
BWy4CZ5QSghcJgFWEW7vk6c5a0DvlyFKdlBj5SVBVQ1Y7I78O9S3Hc0ok9wo4apU
XSb2U9r9b/KlMymzfsjNmCZi/pxYeHR7rHy/XgC2h/kViQldqaMWLPAtusFQGnAT
NMv/T8iPg6p3/bkW4E5sULM9yCEn0TfxYV1iUXR8cqVpBJwOVQZBKamhErdCf8sR
9jPo+8h3v1LAYFH1yPrASAPQRZyHCKxtjPm/my+WZ+UWCkCnxGQGTsS3Egul2S5H
/cn6854GnJyGHFF5jsUZjG2L23ZPcLNKnF9CgBJgZRwdosSQMd/njKzlZsTKrsFv
9i8qyXx5sBqvL3u91WzJd4V3FRVorFhvw3JQSb3m4LO/T0HVrkYELgDsatXGMIec
8Ei+uDjjKM5MbJbYaTzSDsxOx3qlWN60FY3tk3U1W7C5e3Pevu7Icfxb8DHNsNdX
pBS5E2ynmUNwMyABhirX2+oPYzwapOmFYyvhZxLBMz3dV8eE4Hp5W8PupmUpmByV
wzpE+thoChANTJXKqxwVzqZS1BvNVQBCl2M9pFzaF4Y6+kvOq+KBos48PY0b9MDP
3Y43AImPI51TsYlr868ScChws2RMMpLsXZGKaJXl0zOB3qTu6UnyEd3MUE+gRI8f
qhIBBEojn4oi+nh0Eb+YZQAfsZDRgCOA+LrKma4sw0aMqhXJH2e38O40ggCdgT3m
s/0QMVK9tdkoSHddh9d1oazMzI9xvdkrJqzCVA/3Frf+hPIQL6St4nT9Af66Elwg
9qL5ZQlKCqad46CYsJ40aWS0sW9NXEPOCtX4Sf4tuDFzSJNhnLcXda+gJkW9hW9g
6mJRK+zR3NtDxbv96nqOEDo85pcgawkvfN9TC6L62zagCYJ4lv/UkwaiZCTeo3dX
b7cufBMY7N91CsQH9kLEOAy0HNAwePiIO+SUqDhVsskNbGjRMgK3mNl5hoNUn2Ed
w64U1e89MZPTl3n7dEefKK5NSE1+WuJYlhb6fdrgSBDARV8EyiMkZ0gA6cGJVxth
iVCuSCajSmmSHLKmTvd5r024QnKGVjxx9MMx0HlHMcCo0jf9hPp1olI5v+uIF/YO
753Jq8UrKl/schJoHbUd6JiqXsUOe3ph6cA4tke/u6z/smQzn+9nrlOeq6n4vg0X
H/Huq7FH4iju8jiGxIUXmLCJ69nkT+sYDxyMO8/50xBVBzB+wg6IbwAO0Bsn0azD
4YDl68HQ6iqg27TKthd1o1cuFKkxdCl1QorcKnie+jI7BnoVsdVAOqkabbqAq+5R
hlEM5EsadD7Zl+rj/czTKkYF4J7gyZlj4/WtZhJwAb7w8i06q5VjfBfb73lY+Cvy
xqMeO4+csytdSK0Ok2K5JXaI7H4pgpzYHsr89uqF5/ygyuMIJchqhLCB72XHFCFf
gqfvQu+tLdDZClbsH5kXV/pQ0h6EAiC/py707JbGfQ0sTz+rL/jUBpR4GSWUm0RF
HhmtcrA+UaZ0bOpjJEC/dPlOK/DH9QkWhoABwn9etLha03TBVr/LNxGvXZ+TQOZ6
Tw94om7AncZGGGnBjxZd3SU3NurftyCHAFVVFaPADLsj2hCfJ+JZqMioVWy5vk5I
On70u9XJNYWspejYTQ+iYHz51q8+4rqNHyHHfFoSMhGG0LVbWm1GjlrRS4mhzGF/
Y5DGNTyXh9j7ejzHj3rIolKNpYLi2eycRU5PSx9wrryHnvlrzAn+EAHtbjzg2lwU
lgi1w3QRJoO/cwWFCVu1K13+g4eLMzXNggBZGsolLt7LI6qEAnIAP2iLgSvgugy5
IZIi2rog5/3PMKTog7jT9oJlYWeeN35Z0N4otObMyYtlZ98lXydu6jZ3dZaqGJdS
nrPfSLrLtuc2znXKBqI1UrImLqXrRY3VCdM+1LbC23Oi5UykmM0w1gYZvOcIJ+bJ
RrNGrCXCWl2PoqNfhIA9Msxk2tSNow81+lpnlnIzsMHrhc+QhPf2e4Ic7dhvXomg
x3w02Dq04VYReWjTTvV2mHjbxYFbsfV6SX6ywPsTNtm+6OB1/kDQMHhc0Zgrtfh3
NvzXa1zS0d9Sp426pIHVW2ZkA8rt2Qhfs6c/dOsko0XJFOTJWOSA3qo7xCgynSWF
mBUhneQ0vS6yxEJluDKSVmlrAoKlsne3ijfuflHTMtcLfqTn60wMIYi7C50i6fW9
WYg1QzzqbMXw6Q6BNf5wYuoAVY1nRHbN3JwgnV94x4RF00rYdpdqdWnknwhQIoK6
T0cBEGncg8mya8BGbQ+s7VZTV0rn8Ojdpd71JHm1TNduzJUTzdlt7GelTy40t29h
E8h152duxEhsep59zDMZKQPHquVPFHV6sCoRnXmTNWRz62L7nkZnU6HwczwCgtRV
HAjmKcIBYJEroRkNJmZ4vfJYBXY8gsbwhIFqvtDM+XU2AY2HDfMOePPdxDC9Gzer
/CAjnxb4/Fy4CSDaEkXuuLsMp9YQU3ESrwg7saTLiTMXHlVF/6SIzn5yyE3wMaBE
gBj9nFMYXj6wnLbg4JF9Lv4+6iL5yYknlewsG7E8KqXhKeYFC8rri3zSBl0CvS/1
1FloBA9sEjuWam0uYgmOHMPWQW5mtkAAW14AKBjJmEE9oXgwMe6RQq2ScHzanquh
AZQSG+BdtA3ycMH0FVaUor89VHQtNPaYZh4dhZCsCM6lAir162iQ6Cdo7edJyrkJ
GjenoGibFG5sRJUlC2nbwJ68wUIVcNfyUdFM7HSKO4NNwt1apwUJ2YqIns/wUU1B
RLqk1cZxmL2RmQ8GUsF2XYurYjhTLT9zItPXAUUG8Mhq3GW7C9V3GUfRHLxTOa27
3PWovBuV1fBKMsmvRMysVbSuwKFCIiTNDDQ6kyYxpUTFrUPulml015Onf/f2eSqu
d7QtxDqDy7dkVZB3NuuCnT56jPENPpVkfZbMsH4NZlcNqP6RyAHkk9uDBxDO9whN
nzrdwoNO9/FrKVZmjU5PIpaP0oN07g1L+Jq80n9LxQLZcKMdeIkvskfWgW7hmEAD
Uu1xd4SSVPeAmu/vX7YD1+bMAFTivxt9GkVZvq8tYDyDUdZDfuKApYdbPbl89xhj
kSnRF0V36WKCtlmvoTAzZs6CBSSpEKTx6XhtkF7Uk9LaoCvzrDgn1aiHNPbsmDt7
tyxKlhO4MY0LQC0Aj/9vU1D/Dd7+B8PDg9DrHpN1k9hNPfUW8WIvra6GzztTAFUE
WGBfWyDGlTnsKWETQOPmDn+4YdGcFb5D8MYM1xGqn8FOtUBSI4A3X6L0ryz1R9Ni
MIAtlYrqlLtldKUQEMOJGOC0AL43KLISc2Gd7m5/+sF4r5KW6U0YESFZOLKa5Tv2
n+eZmXlUIv5RkVUxyzUZCjF474V0QtZKFMylyyNhwolSncYoRbWJrxzTxp6pGPlh
sYe1buZYQCcO7Ol8b8cM0cNkvNOKGUBQ2sFQ4HGXW/zNX15JNBRqR2tUnQQmQqgl
gRA1OJsf0rPgbmEkwcpor9Hl6k6V+nSe+he/oSEi0JiE7DI2G2SJV/AKtRUmShcO
+vSsWcHnJy8zruOiCQhp1O/sUYIx0WR9RJ/s7J4O1zIVKebUor1agnjOJ2qm5qb5
nuhWAdZLvCbZ+cGI/NiiPK74BZhQw5bK49NmoZzRZz1DfoPZeYiDEbm+cVVUBWJX
NLjWyCjkW0Qhzxpo9ndhLDzxOpKB3TFJTzoswnL3MJrQVHY2Fo1X6mn3tMD7vTSB
AFE2ned21cGlmQaSRtfE/JLb8goA/+2lfXt4rauuHNISeJPJQYcWUrFc6dgjiRZ4
M7G6OxkYTqhh7kzKN1OmXCZTgCwq6UxHU3Ban1VvhXbQ9UJaJ7UjCwpOEf0+SwYv
qPU1ndcgsrp/IOZYOvBiqYohQFVhhE3GLcSE2EbacYzwYrk+IGy7Zq5c1fixSWGz
bHKrq+sY2rmNMXZiX7yjU7NLxTJfz9NDvqVExZORU5O/rd+ZFIHpvo48yvgZEzz/
5hiE33Tc83jzgLoZoSuxgKOOwcMQFZ27q4KAOCmn8YH7sZG9cVerHCbkMwqJm7mf
YNgr+YAmCDgRs69ENP5hGZqwHeJ2xFWl6/XnnlYs35LrJ9A2PrVAwcuDxXgI+cG/
E3BedFe7qSjAl8a36q4hg7ZlMvCIWnamT3igALigPpqdlpWE/2vRdxjZRFFhhMFc
VDw/dh3vG6Yhlp1/X8mleLvURHYIfE/w01jGXBSwjXR03TYjB2h4nFgt88Mqkvgy
eAQX6cCySmPp/ahv/atvN8ieJodroLl4ERY6KPGxv1qLSI0CxdnGU+946m48n/uL
/ffZKGqZaCUSlo6+HyTMqSxqv52kqxFjEP5GJj3SOeOYxVhZ8lbkYJFVKBxJo4vD
F1V2SeosLgrcLWc5BJpKlrRp3QKGWHt2JHMfkqIIARK6U+YDVXgcG4BCfvCKfEwx
xfMmvttB41GZ2zznC7r3prOhMNZDkupAp6rCpvbHI2glRDbDSMBRkRBx2O29XKb5
dUV5AO2jod4HhNsu/z1jeOrxK8S5FTjfd7xNebhmil1GY/wz94ofNnXAYAFbWVf2
uCcC2zNPProug3sSPNafNiMfY5N1+NIcvrsDwmQADYjtTONdd4AS7Nx+LD1Wki4s
Wa4i95SpiyN131vYHoOTFazAyWGDV+aSK8eS+zhHFbf6/ktSo45+78I2yQMzhETg
NP6BgV/VAdqtrN8j9ENk6tmy1Z+JWWsHbudG9UAEwV8Kjb1wNbxylYLBC86JyBdg
aMLoMbssG3IWEbHTLPMECSOEgRWJjMJ1K84N4g+Kk/mXSxKTn5V+fCU6xe9lFGaB
md+bK1J5BOqwPuK1BgPB2jgLjFbCN+5LXGuRrWVxEqu1w+r0CuLZXIheiPdfSqkE
zC1UwrIXqnMzmr1Qsnl2q2JwzEReO7N+izV7+JYeyjI2/gid7ySsVfES7JqnBPJK
bgdxFZ2LEeYYBegWjOAUYxTwklb9V4bvKS4XgHBWkBle/+KrN9F4JIamc+hcvhFP
1aOs+QPexgHgKiW1jPqgUvzHf0vySaSfj4LXmWu/mTM5mxxsSnDvu5zF1HUkF5FO
xtam1wJ49vadVwQ+TnfO8oQEXyUKeFLhcod50b3DlzmxZh7xp1DToHBBK+AZcR8K
nTH9PH2xQG1IrJMS7YIdyOtC8S423QWvLYKFwMjhgcFDVnf9zHCsFoloe2uUMhEy
IFtLNt0t0JTV2kMuwxyx7GUbjUO/8BL+x+ZyDkpmGbFfrASXyOC7o7fYvwAXKkFi
TeIWtEgNqeTF1zk2isil4SyumRdjZI1VYUnJgyCq7a+f1NUQgKSbBYbj/9yEpZbn
aabQx/RMzaXM9t19npuQTWhauFMlorjR50laskiSUzysXaJpB3D6b9TvcxvNwMpY
GD50JVEimnW6TYlwXv3EcNYgZCvX97Ks6W3lJHa0YWlKZ//DlIyKnchOgBpM2uHF
ak9BmFGzQHUxXr1R3DTtygXYrN7y1M4B3JkIDKdMf8KWIKRJSeFEK0qWqWJStxtw
QDWYWEw1QRH6efrPQQsggQPcVxjkLCp9by6tmzDzau4ODLNQcNR5pdYyiowplQpi
wmblYEMHZWZBbxDPid54V3TL6kChb04iurLa2K7M7mRDrHazVtxn/f8G6xfuIX76
dc6k8RegqyIZnzvk9syesuzInyNkhEItAeDbhP0lRCR3470wctyR7lZuwS+Kvx+I
kMQ9O4+VXiaBtW6WiAcQD/ynym5/MUH7oxuDLybvIniungrSUeLCfFj3yMCB6RIo
qYt3RUDNTRy8nk7lZLjVe0/LRM0L2EKPlti8Pz+1Fn+Ohf1UMUBB3tbMK+Q+e1FP
w2PxlDsKmx/uKuRJpZ35OjASQ+S4HLiBUUWo32VZvjubuXoeNuz+XoubpcMr62zF
bEFatz1z3HuZFd1gsD2XAsUUGj2Yud4tKkD+WwRJTY+B3HL6m3Q9y5mOU06Oosig
w6qx17zQSN7Ziy0t5PPqv6uKOZReqCiuh8BiOA3wFEYgrO7aiU5wy+eVLroS0FGC
MSy/ZiA7omUN26akcWgnlUDnOfmwiXCJnawVtDc6Im15Dic5UkDShlYVq2mlUzRK
ZceznS6OJx5/+4nolEjPQHBAJRbfpieLKQrsHkuVkKuQ11rpyx4xGLhX1cltz5bi
C60OndU7d59Jjre2IKjJycJjj31raR2x5/C2i2NYTY9HAfOhIsNsU3+qMKbCdLnI
3gNHnqtOib9d7E1/h+tVdP0C0Q3ZPNhjwFvDlBpFvYjv6Kzstx06czgeSvyYlvRb
VBrBe0uFAIZxbFeSaU6KTqZwpft4ZcVHGBeZwDUuiD0Fr3wqSZi+aQMWRmKxWN0y
hNzWxbBrdhU46ck+6aD2oDbYsWMQCfZCR48bE+iTZbEYpkqEqg8TfkLGC6Vi/eCc
BJH61xqdk8yfgwZR5b1WFaVBb7CiV16b/SS1s5woXTNRrH38N6HZeaG5xdiFUTD3
6crdv2se/ns2NFSM3toVsYZIWCIzpzZWnyIlGco5OI5P0HV+y8mDi7xJ0LqOgVzl
PVRbPkdy/a+5BnOIgGlkhzQZxvIBREQXwh9JwlPndxOnXOyVF8yMx66swnzRFc0p
CSw0RZpxBmOOmozwyrdCbo0CXdyX01iqCxmpTXdHP/Lyjwzg/HqxfqW4cmgS+tqY
rPNiRFBVxAADZr9EWc7faX+s0d3RYt40eYGQtVYHmUbY2eTQFeMtrMatPpVchjDC
Y40gN+NLcXaxcQzG8y0GabJSzRAjoxIX84J0PUuBIFryzQNq0azo5uS7FY+0udg/
yQ/Lg9RNFz3/g9sXGF+tBxN4DpidClG3IkguCjC61kAUvXZLA/9UxHX3FvTpqFqj
yGAdl9XMRKhtXtx7UvUnaeqMtzQ2uLuCHHY/h/Cuc9Dtp2ZiAf23WzgyCKRW0msw
6iJg4CXeyfj+gMjkD+uINEii+enz+Hmf5bDqmmZOZMOhkofIM0GY0iXUNAWfD0nj
J3JC9f/B7LzC6b62rnNw6C+qR2mgu3ubCmJHgrncs0zphYxNWPwe89MRIt12U7aC
iN1c43OYEee6a9nCHcsPh0lhNTyKgsB0QBAoUH4otGm3+jI+ZHB8X7USdvw/989e
0Isy9JIPVxYEf6J8w2j0Cu87U8tklhrl7AJ+CuJY34p+66wpZ4crpSWUCZnQuT3+
E3UmQMfS3IfJFp6/KZVXVyE5QyNiDLa5Um8yCBffKBsvXtvvm96g1hDzozQONvXX
2lh/gjKcbtjL2LTsGlMHlCorG6KU8cPikZiMndcMWFrLf+UOsq0cWMkG1jXHLEEj
RFBxGRs8Ipr8uM9jfHWahb066YumVSIqXGQzI3VjpvRpLOA9G52XVNa7bIoWZpN3
kkwTQ7KlFP/KwjuoH8/HC8Ro4fGQKrTw6qk8OFIH3H74/z0/TOccOUNsnLWGVIE1
BEJ4jDPa7O7UWxtsHzwt1QGtgnqBd//vGI2onWSg4dDqhdAO27D9rs/ZU6fhfDZa
DxVl/+PZMylAKNEvjulIoalWotnjnvDPs5f1lOG7AXb8/8bPHCKPYe/B1s0vC3uq
Af324IarDdPHs2KrsZuAZuJzGQYDOu4+oGy92AcwgSIHsqqouquSUIw+wUvt6JRj
YQpO/FNhAwgsZiycRNp/e835+MjnQd48fBiutSuAQ2IKTCDGtzj+V8WsUpZ4O0eg
a9pYg/uh+h5Zbyby+oy30I49JFtGVNPRuQGlIidGtp3seC0SADf+cJJlOPx0oSfa
WgmndidW62hMNdYiZlb+y2xVT3izUTPwj6BIpPjQGKLCMPcacdAACJuB/ffB5Ty2
9SO44pdhclGKldv5C8ZRIXBCbbTPnYwckYd9jjkoSMJBmZ1+e28X6gpCq5XCE3xJ
DGI3JYcbga0w5oH5b8X4L7g/ObAWjYpX+Ze9OmdoHwooQBJG0EvdXw86VSd472kS
WbhZfvryOF1K590a4I5pitO4sq4/u6wyOdyNTteH+7PDAnwaRorM3JtpRMfcMoO1
hbhpAGLvTyvNJ+YLmYgbCjDjwQVjMH514wzgQBW4Q4qFVk1B0FWiZjUu7UbQ8A3L
a1dE5x0fdvGGh/361KVEo5lBFGFXddqTV17V47Mac/AhOCGmEH6dO3/Po+t3s2rY
dgl76KQ/zWZyHbLpLCBL59PLBHFQF3csbAI6+sOHSm5htb3bwdCc0yvLQPDtO3uT
0KKtrRljTZHXNjnUxBjfNP2cHimv85IDAAVVOqDyDwrmx4P0Jg0whrYdIhndaKcW
uQqWBeyMvSKvtbOM4iKcZLx0GTmnTlJmycPlHLaAqlwj88+/UrYXCIzFi5h4RRaU
2Q7na+hCjtKkUZpL0hA0t6zeGQoWQdVTkFCYWULV33CFTXL7pvYOOaFHdnkQzBWH
LDM/ud/nCVinHgPAwcd71myc/to8iZ8eOL5W9LXXP5d5iX1J5/m39R8RMf3M+LIB
R6YfCvFyGR/f1Zpzx2aj+mOx6yFjk9b0ewhxlSdhkI4sxr9q1bPcW6wXqzghsRHo
Xb0yOgLjhF2VzOEewpSRlgGvGqfL/vr6inGKFNg8QhbDZIoQM7MMqsjLtVyrWfv1
XSihOuGO4KjibS6p7RvyhbFEVDx7//MRENWBYAKI+G6MV7jJFpLu799SCfSblGBK
zwMzxs6W8mukkTURk+n7gr9OkxRPbEkinRFQVaXKIsoYwQfLim0WAMhCx49nZO7X
JzWgISNLy6GC4dk3Mqnn2SXpU5f50hUTz0sUxiv7t61kkkenykxAUHsTAm11XMpE
xCtthWo0LplA8H8IWjyI9Y15lunl4WM1mU/iPebbQ7i3isTBdCvf6GG5WGivuycl
ZqwUtEs8PQir7qVc4SxpsCXERV22qp4Qgy0weqL2zY2W28Xtl2fmn2aBXpHdT2G5
OnwQsbOxTgVvEkTyYIs1huxqkGRT5ghK0UDhehsPAFKkUQ2RwWHranAg6H5nOeir
X43KYc/fIFqk+mMfZKigeN8tkWlP3B1mQf5PqhTj8U+YgNbTTD9GKs6O5Q2o4rKw
nYac9P7lCLnOSkHdL9kVy6hkIV7EzG5+ou57JrLwizLReeQtYxmEiE+4KXkbeU5J
Al8sd3rFt7yWtHP/mOFDJyeWOpx4Ub5OfuukMII+jb0JZuDXdchlnndro9eUtwWS
2D0DjZqis8GGlrIk9FFzsxS2mfpux08mLinp41dO2heVj6+3c3BQAAzx4jub3gc1
XzGflLaEHqsQP5XtLvbJunf3myFMR2H9GvhUvMb6PFaUZZLcodjLepO51X0g6pbK
EJ4chEa4aTHtl3U/PWS7CA8Nl8OIsjd+w4D4Hart2g+JKGuYUCK5aze7VHy3YCd3
dnfuJNR6FxusyjsEIXckI7QUKJyPnXVcUckZcS9P6mAELknmclQDyLABcGOi4QQL
uzHo9gmEBDxy7WTVECYSbUVBpWcMt1Ygvn53IBDWh7Ven7gIY3/2fu3CK0Fq9XA/
AjY+RW9cWbmXIOQ1/U/zHY9W/kz1KJH8U0qwgfXcf/ZYGrQ73Eqe511IYKrO3N77
OkLPBfuyMZ7lenPtW5hHszIm2h+i+ajXnN5mT2DBGlDg1iyHwXyHxCet5FtSzvz0
JlYjf3D2Xq4W0JG68AIQh6tXC+lXPZOZF4G37DraRJ9GyjopgzRAaGyNQHWnWuir
ClLrsw/wlVuAxSFBnk1+tmCZiGLRUuCt1Y4HcAWbHL5U33CU4+WAxN5Wl7wtqkh4
Ly3q3QT/kfXPpUzylYIgoDu3FOpYeB3iTTh0hhFYFfF/bc6JVQKwSTCuZgIvAsW3
DbOZflozOahGGNd+d3aEiY1gqqFNwTu4iStdF4vhFCm7saq1LYYPtX0rvgheEFWi
rg7qIf0KcDNhhdu7D6KWR3ssTzgKfHS5+VSwzD5y2O6jcPVJql6ZVF7/s41dYb23
7s9GKJtCVC4/NPr9XbiDaQVpUY5Y+Vbgy6zBtzZKUMLIvkHgQzhWyzXDJZApqgHr
JGWHpp5h4dnQTl6vJzeKGGt5cQZoDxhdCdxbuaAR1TIGJRqFkOUAwH020eg4j65C
AdKLZY20NKq0P0fPD8B75OML6Q7iImJgkjaJ5WZOt8eDSp0qXWdeLyfco+LPZHK0
Ip7j0ianIqCiC+MZ57gZ/+XSig8NDd2ib+xP1XwB/JDRVe8FTtUkHK377xKIfiIU
TzMNxbcJd9Kz9CW8VhpnxDQ/qTIcHy6tHJ0AlcM96hdNRF0TjbzsJy5BLbCr0KF9
lrJp7PSyyjchTPu4BZep7+z8DYrXvAKHvbFhCPifi1+tcNhXWBDngWHHWFzQgBTy
3nHtdflspSpeI3gRJ27wAKufuj5i8bTLBID4XaxAM6pZXwYa8dCWWpwckDYRl/aw
F63bOVCHfTU4dNPDFGkKlnu5QZhvuA18sS8v2IYp2nlatklh0mU9Sfjn+cBhHkhM
9gSlax97xPScHNBDTaqZDu3L88TJbvqRR05Sf6Be2XrqXxpYJjRBNHVPgSXgYaFH
5DnArrOcTJbiwULpYdYUNcmx0ZPuRT5eEHvu0tmmXvohE4fDyecm1xiKWllq+NEu
cx+kXEUkphXjiE7ffpriMcjCsqRJsaMoWHpF77vZ5rQOBRZBLUbdk6uCjclwIsNb
dp12r21IwBT74CkJF6UyJPAqWNgx6O/spKCSwxcrKS5mCRoS9rfEOMowOKf1hihI
STw5JqdENqhOjHy1MADA8ZyeYIS5pVzd7IDgkH2txZy9OVzlXyzLj534350r3HU6
hbRTj29CvTv9okvk29i0XfnZbwYAYFHqMLWMnqQ/HlZFezdtSlVnAbjsUheyoIt2
cMs3Kul54m6fPQyMKl0MnFvnRgM6GWV6tQFRE2nXoNnaqiTmhUzxVIQpnsytW9J9
wTfoF9bSkTecbVA+kdg5UbEN/NrIyM0FY/zqEK273OhqYpq4U1qtR2YWnBVkbKhk
AySn6qrVxjxra2pj0OG28iTu/6CvYP6IV1TOMJb5U27vXKB2LjLjsiQUHPJUvmqo
hvHrm2ymD3FhzJF9lM+yugYq4tJqTlRqx4cK4Z5FSl87/F3NJRLivagZBY6WPLjv
27N+Hhu8oOSBIPfrTF1cAJd23AJ0HkBjBqTqMKykm/7BPYW9Aq/eBHnYZVOeIJ2g
VsoGv2dwfM5FM2o7TD/JJ6hAAzTQSQi2tRjabTXXtXWBMJJX2YSgcI/+pz7jsO3N
GJihIns0qnM/+mletd9W2rfTa5k6ubASD3cMMZjxuhn44H+GnLTP1iZbXOnn79gT
9qXATwqZGa3b7lM5JANZTtTcfPeja8KYv/VMkfsfZzCFK2aVPUAyp/CYM75UYa0q
43lo/dCXr+4U1vrDoDz5fdVmO2wYyMEJb5nu/qJjnqrglnvHMR9gdLRbAhb2HyBw
lXMqV5dfHUGYfqcJZx1iAkIRKLUKTnoP3nJAIjZqOWsl6Lq/OoyL9OBc8jU8U+0A
ZsSNrwBDyasOuvWRJcJzgLlsBE2HldXY6QglXo6UI7dLE06oyxGhINPJq+KGt6PR
GEzN9Ef4YG8maA8KRo/SSyvlPnd5o/pDCDLcJdDcfvX+1FSjCVQqJ9+Fa7lsoSok
h4SjMIptNro0RSTD2RuKoyzbTsY9aK0q5sdfT3YmTc9k+oj4DUiM85KE77JiKM6E
Zvlm3rLccut4av4X77iJIt5G6T17YjsgThrSHZm28qzIWW7r6XiMoSgFKMrHDHwl
loDI5Nq/oslwc6kCaYHbUne3SSLzW+AvE2Xrp1dX/1VnluJQezX99IBieabVjdk1
/csauT1k/4nqBpJ1PzATLkN8qBFwXTNdAInWtwPOqUbAfC8PFsExX3Wp3gvx+RbU
O68+OStxjiGVcjVjJDaqftl5lSJb+aeMsVrsqOsMJV0Aje9r1h+d2Bac3PhsB7BY
zpAb10k6N3e3xP93+3q6ZyJ/lImSruNHEQt/0UQYrI+SmTKGMUyIWWCFIKiI+ALT
admgJulCE42oF+n14UJXeBfawUETzTqc94xlAze/6O64rmG81bPG3EAmXE1EiYEr
k8Az5UzSQT0wPOOR+vDHmkG4naycnU7pYxLn+HzJ2IAo9kpSiaFP8qBVqq8X6ILs
Wp5/IHxqpKhJVZECcgVXjVnfGLGGHf/evQSB0+vuXRxfsO46Zs5jRyP3Gl+BKa2/
ubtpnGg7ud278R5ZnKD11b1xS8/ikcXBYY3K/W4l9fUoNclK2o8DrSQqNjA5OvFG
F1F21PGCUgCAcF21hb6lC0YytG1BNcFt/OXmj58amGf10rT1JchUlsCW39YJ7EGn
r6aSPfV9CYOmpwWEU50WEK8aZFHISfArh9PCZtZvnyAI1PO8SVb1uqRR5rdmQGSK
Is1ja0dq/nj8B6uU4agBXaVOVIYrL2vMJnp2LjQmuukMKhjTr9TyW3HVn7uR0bev
dJts2V76RV6gAYsnDvMUfbpgAyZRmqgivKfd/tC3hCGqLcj98Mh5vebi7yHsfbCv
bjoWDJ01Q4ozBA8ql2PaG3DahIf1/i7A8f+9T4w/V326YgO31D1sAvfzw0TUp6/p
xrjNyMDbew8Jt0fqaDoCe6x0qJ8B+/oNOU5aRrSWfCsz12kc0pk7RsbJI7X1kfXM
g8qzHyaJeaqEpau0TAvinqUHO//+9+iZG91WggFRzXopmdvoyeiftnz8q5OiSrdB
oNfcxVcbPef3k3AUZxJkuFASukqHdhCZvgJfY0hgFZGBrikyYB8e+FNb/rF/ivPX
LFXuXY37NPMaGyAWZ0M8Eixj7icymw1gJK8FGPu1Lk41hFtLfwqK3OWIjOXKrfMF
pZeICjcEU3h8SC1Jd1QczIl5LoXGLHfwhcFljcwHWghxYAUl6sHhbgmEjtYRHpQa
nKYqYnmXyW9yrUj4C679hURb4qK7GuC1jVUM0GdZjDjHJifLsNz7B7njyTOcplSJ
39b6l40lXfV8+T2OcbW9gWdTXyTydDtTpfQaFO2zLmiqVrDfj97tbRPuMNeTUHMA
BleC6O1RsX0rU2dnCsMwULxtc+WKONA5uc1e9raIHgZgYjxhg8Srk0vnznQrx8w4
YA3vRF+UHE2vjqjGFgFzaaPh7pcn71PZ2OcBORwtpB02qFnMTeJ4iwsR542ymuaT
HsR4krRcikHnoWb79JgHW9QCi30tKIXfMmiPHVvjehBZyjda4j4hp+FuYPQ/IU3Y
3MXfqZxUGXxlONKAKJs29UaZBEhK4HnZ1BzRQweSdCJIMixtE0OA8l/o0A+dSSgX
sLK7KK1N1o29huIQVbQi40XRkuJE39uFoN9hbVS23Ia3v3K7uZlZ+FVSYydI4uU2
GrXCWqhNkZuig8HSVthR9R7BUgL0G+KmRbeGxn0v4Ulg0BkRAU7x5Gv2Vp2jSGUW
Dbpw8kVBEZ3PRhfb8IM2KLoFR+9MNEcsJ9SUPyYc3ZiBhBYjPDlDdfRtKuTuweZx
KdPTJrsQ0MADL0K46bbb8d+3ruZLfEXGTtQNKjpwxX3cHZA/qaadpFm/A3wmW1yT
05pLk/FDtiy0/DFC08PV4FGTVXVsbgdW6xoE+hgef/p5LSN8Xzts/C6XZ12i7TVI
TIonv6O6DNY970bSiuFqGDqR7JjgE5a7E/WYCR2zJselX+SyU2jG67Ag8affazhP
ILpvDLRzqdU1fbYmDkmzNq8PhPfHC06IUKUATPekL8dTkbcmCThclZQGt3S5DxIo
Bb+HBQuiKjsnbesvV89cuipVdl0FI7QJo6uwIvLEn46SUx0pjoaN8QXKX2Qz2A7X
HJR/7qGlkknZYdZ/ZmZ3Z8EXNof4lxoyavbhQj4kDiLFReVaeuGrAupvPG42BFPo
q84GE7duO6Fzim/Bpw9HrJ+D5IkPz+9IAx8k0dA+1qiR2/VRm7OZ15XNc9vkreyA
t2H13qDUAHnSSxi8cTKqkSqtBJgo7hvIhZEN0o+LUhcwIrpEeuGDzYiz715Z8jR6
M42lmx8cwhqjR4ZVCarVDSXd3+dO7Het5hVtUEnFdMHyqV+d8eOw6fNbnYebIU2l
9wVlefXxkL8aZl6Fe7Gekd8YEn+DkDTTubfSpn6EF1e7wec5nnYW6zvXLoN+LQzk
yE3iDpsZoPhVrd7hU/0/znK+Q9LhnuCxxN89oePYk6SrauXVAqmmx3ELLvM51CeS
r0C8f1iz+w97hQJT1dQxunC/aQMaN/xjQH9487I3Rx2d3kURCufUwE7WXrKhsf6J
IPszxLQcQ/b8EF9ZUCDhUnuws4KFM8ikRvlLsDHzXVxzGhrgzlEELsdPv5rZbZuf
JpId9BJ20sG0kOg3oKgfk9woAguQqkZlD6lAInl3ygfQt44OCBC4XIynDe6EZ4ZH
DqQjm99zAMrKIxOZLlvMkS5BuwrAj56BqLmpGiQXLxyf2V04eShp+Vrm3WmEIdMl
4xVLodZU2wPIBNUfIk+Zv5B9opmSgTic/WIAF2klh/yD4PYE0Uh/rFh+Uj0+zMua
5tsb/IQA0AZCo1qzdkFrWytzhpQJ5cT0E/fiNTfIHIdBRyhKeMtEosJVQ2cJhZUX
O34jctMsT1adrcdoFlhc36dORwu8MhdDBaY62ln5aLgUEuGmtrwhXWX0EL3oHqiB
Oiw4xuIUcHe3CKl6i3PwR6l2Xt2BROakTNKGljSviIjpuSKsgNSPCnpCHknXlmKB
IQRm7xdg0QdNexYtVKEqb8O9Qo0hIQ5tx4yVJDeQdnsm9BrBRfMAi0bX5fHqQjJ3
6K4noRSddNbj3gcf0k7KfmyNhW8MYq5r78oGA4o/mnapEfjtlxquCKp4IYJcIdhc
FGgycbcpjZM1djwy55xzDNkclcO4OOY26m0Pk9vu8M9pk11iCntTf7J5ucMihNyS
TxTigOjabUHw4wA1Py8im+0Hxj7tWDH2jxpxcdyF+yOJAJ5SNziaZ/Ag7ErsMybQ
KxdI3sf+sMjqRHXG8XCg41c0QqgZO1SFjwdL0l1QniveNcKihomfgmHarQNowi1a
KSleoz8QQ0K7ALnm3x9tEoLTW7veqKbpEkHmVH7OzDzR/MrcQVy1iiJOeR9M5F3J
tU5C6FY9t9AQjM353bOBob44mIMMfoA7JksUQQ4ZjzI9CgMIqVE7I6K92YHblcDw
PqKwZiLqw1Iapu47wVU07OUk5Psl9+VDQLKyCZA/qHlEWXIuoAV5A5R+6WeS8Bku
zSLMg5wsYMLr8f6voQ/yf2NEqVOW0OlH6szeyKC/nUTJKg8+Wjppq415gk1+mOk7
IauzuDHESDYl3wOk8q1IA7b8iWG4j1jVy2mg0zPhNKzWGwd4o7XwjGmsQzUJzBid
IIhkh0EoIeKkzTKK5uSaBJRzl2WCp0m23TmBjSOGInKBEJhk7FZWEnfxuDe74z9q
9HWpP/mMQGeDKjJ27o3u7E5eKnNcmr+UN+M/OKZ5vrWAvwz1oB/8XsF9Zm/FCCCZ
txf4Ik+P7xBtUleF8jX6LH0uAnDuVo7fn2LoCE0Yp3hhrFzf0CAT+FtZj6j9Bzsw
UyIsPvxnkeU5PQCNTyPZmhXgzQxVa6gVH9O/qLch82BhM5dhvlph0u13wzVGOpq+
XW4iWUWrbyLfACst+yR9uwigveLS3TfMXEXLHePUu8w0YIOiHCsBZQB4c0ik++L5
k0AQIcHv5tCrCdG4rMMOll0FqPFM0aZ9UkYM7845hrXRi5vJo46dEWY+d5OiI/Ka
HzlaDVQke8prs8gI9dt6CIAptdRFcy1dEGqu1B1x6n7N8Uq9WYg9rbUlA8GBP71I
14riJYOmSqru4BWxX4xsQu6yL8872nyj8z14ybu5i1D3izfaiAdhQ6A2ua+KaV8b
fK9cH5ivE7/mvFQAGhak3BDVBMki0rajEkfA20WOGU1GanobSkg13ZT0ZvrQNrRP
eap0YGT+WyVNCGznh5we82/OXaLVDu5kPPAKxzoORHV4GjuIdaqe9FCzDbDRrpQp
C8Qd9+qVPlxVSvq/3sVRdYzj3QeD/620Cth1YTKkj2c4mgrbULMfWnvX39mxTkfP
Qw+XnmkownxukrIqWoBgBSazvSnFPdyZZEOmXCHqpvTyBdVehMINmXfeZrS/W3rj
oxLQQdLo49g8coyTNdzyl6Zbgjd9jZi5GEYvs0GmEbtojmVlHS0EFNEWPWgkXMQE
I3qTP87ReY5rpK1gdEawy71u4IbFwotkAjIRmlAjiBXias+uNobCXMp537Gc7eRu
11mkGxUbNFO0n6jGwvc8yilSoGktIYDaAoNqUt87JoX4q1oRBwCr8ocgWO1DcNVB
oRtO+/Pr2qQIDaMHFGG95dg6NyoXctT+4N33vQcQ9HoqGxGFNArhCADNWPmTNfYi
o8mM12uToGoDjMgpxJW3oQsb+4+AcZLqxU8oGK/zJJgLpWEXuVq8gYDcAf+iNWtn
G/IFZo4oGomJ0BIO835lcTXddwLMjKey/tyd274CD/Gg8T7fzCWVPrVC9VlsdyZ/
KnBuIXAiS89AXIRFgRueaFE4q+wNvUTTjocGyZX9V9ZF8swixRdQKC6cBJkauhdM
AFTyjLmI4cuYCJg0J+TFjG58Zl2vZLEG24qQ+lvr2xu+LRCQBRYWYwxU7zsfr1rr
fy9x6W6gFZy+YYOjb+BvuOp16xm3Yr2jv3c/RZi0FBMPVcD4b4lkcyHpnTzJCQlY
vVXTL0bU5mWzbjUQraILeWI1hf7CKK560yob9EM+NaxuHdSSoLPNKpo3JAc0sKyX
ENaDb71ESyZozw/uTxn5HQ7GQZWEJ0mSlUha8L7Y6O/MjGggFRAecBVhxTSkvKN0
1qqfA+8PvrhhNH1DZVdZVwfZ4zzOXlQqIO753ITTM17irZ5ud7H1qAcX2n9LLbR+
ObLYiR0sfNqpPcz8JANT8S747q/y1cz1ThEgSEjvmaMzvhT6DIy7b+2VnginOeRU
PSuMAupdL+iB/wZ1fFkFJraOGRseyjdi4/JsbQq4uHmxw+05/nLZ77QRx8KmLp64
AesIn6FAbsYmkewhtj56bFxytGk3A+IZpyEbPkLkVlgYB2VkrCewyqwCRZTpsX8G
xS4UbABtbNs+utRN0oJoZGjsjq3zUGFFZBxYASt8NWoi0gba7ga8A70hbm7cvrRb
fKQvXus2TlwA7dPVBHEvL9lG+Ta52kydXJyBkRfGaPlPjGXjdQe07heVgmqMtM2C
3OoEohzJ0N4w27+zTtS5MxHsKYFbYEO4E30QaueOgtf24nWq2N0pfkrYMyeCO3KY
sJu72WmnYoxpS/XH0L74DWuB/ygOsXY7gCRGB4FQz8BNMpK/VGqPHgZ6kAuBk/Mi
+GEPG3XqPlBO+Bs+ZetUKtJQcmUko0Mh5X614OYMZzHY3zEijt6b4XmW7C5uYDpa
Al5w2cbxwy7s82Qj+2l3IQPiGOjPYwdKR9+6o/QvMEHEkF6iGuEfYXU1AtK2ycci
DR1cZkDSFLrHi+chUOgzjsuT4bhlcoYUOniWgilzqk0frWvzYP2vZwYUNi9iloxR
BBIQDrgwYUbg0h8q35bgYUkL0OE+4DQntSVZ11btR6kdpyp92KYNnMXT9ItSG7H4
CGcDmvG/qlS2IStZiLLDtEWUgUt7n3VZFOxx7Ug4icqk/0GL04kX9oqRlXVhPHTq
DZ06OrUiF3IvKaDAXyDcXHvK3wnlYMux1MbLkMB3d8jQCVGjCxyORrsFICE+PY4V
wAcMB8+R7c+03tCnLr3ci7duhqHO3sInkEV34X5h1PV/wcI/ymXRY3fRNMan1VPN
ForRAGepiKjrJkdY1uxaIxuQqQ1BMFcKYhUPAy66yTim7E5bUy+7Rw6W0BSvoqpr
/QuKhCLpGxv+rH5g1wntjHno1NtIJkUszxVRR8lWNkAKtPHUEAKDQ1giULLJayEl
+SdSqJtaCOaRcw6y9VXbRDbWgxKeb3UiwQYe8QAoPd2rzJfOpxI7rxw2WQ0UDn4/
+9b88LpRtWZTuO5SiZHKAMRZj9jzItKNlloO7G+2EphoMnCzBavndMx0POgGnV3C
81orZGV7D9Oi7hdeviGKdyJu6mBZjKjVczSErNUiP7yx8hTlE3/lNKnJ23XhJAgH
4RGrwMos/DCCFvp7ydZEwk3V7i7B2DHOFZkTfJWFnr4BEn3Xabl8pP9fGhM1cGcw
aTC0v3wiobbUeDndKkYl/5QqQFVMNFZ5uNm7+4tWfJC1yxl44nUh9V693gfbtq0Q
luhoAo5Xh3xGecZ3qxe9UlxAIN8bW4Sqpl4boNZjVUiVO+a0adb9f4pSqvdJxGaj
HueRo+i6nLQ/1G950a40o93cY5ok1qauQNmrN4DzXylqwoaAZ5AywadPyKef7ted
yhbprTyZn5w/lxaW0Thd9nZAy7UWGhmd414/CWoAV3al2GYZLCa08zm11uxsi8Z+
vBhLhcsREHk1OwXw4ZZjOZkB5lPZCGGH0JyRvohBQNBS6fm//D626k4DYLiYd+X8
xzfYTHmzfywlfH1YtHCyZNsKYq1EuBxZVCCE4qllmhbJ3diKYOReR+LMkhudSIo4
ppLsaaQ6jkrcimJfj0RWPQ8fZHOCzc0C6AZHmGuboFm0mKo0HNCbnMxIfhVY/tEU
0d5/YQ+oJRaIu7FJjRxCCa6ZYfZyG5+cDkUVB/cYaG3I+TzrJgNErjHlUyywn6Fq
ux++LuWt1e8mkLlM9oUusTx+gU+WVFZclnfw+z27qbF/Bclu9TN3C5P2qEzI5xwK
2yBC9pPR8WzzbQAfJOhC3UDF7hXCR5l1kHa4v9asIxI1L7Yrw60UFgPbNyEcbWZn
9rZpkyN8WEMO5hX1zi44erj9wNx9ypDldt8M5KlDJNJmZiJzWX21PpT5RSoeFDtP
ZZbK49KPj4ackpPTTQgS4ZnSXyGjk6LDxXj7IjAJ00qAP5WX+QxMHfETQLeNqY8k
R2aX8nFkQlVGI/jg0Sekhn+RD323Faa2wif1JFB6i+BhcwlnKJvOm3dOv1z5ha61
J5bi/lX4zZApQIYW+QxlbVVM22pJm0ZGboEX3VvnoyCw9DkItDAURXK1RNy+eVfl
7KFvO8VoTnwl+1Xszz6rzJX85l7whSVjrHH/rGl6Bil+ST/Lr5CCEpacK8hr41aA
Ku2TvZ0AoWMl6PFl1LErXKDy1gnlMz/Ec/PHaIKbrbsmbIyJGrYEavob6vBbHvOQ
eJ3RJPFapibiuDTy8VNIq0+N9ux8/XBCEs4HhUztpn6P/ZiKe2uIp94hgU1mXHkH
CIXKaJaHBSv++LFc7fHJuN4T3O9xxovJNYj+jJz35YWMjTHw9+26p+DpzP+CVXGT
5RpZp9J3/XMnC5eT0ZtVcQGuz6RXesCcLO9L8eUlH0RHNfKNbeMqlmWJ3/ChT+Jn
n5M0DahJVkaB+MM7mEaiSfY9WX6f70g2oOF0FUdF1UlRPFfD2ZC2i7n3QLdO+4v0
6F4XKXdnlKMQGMxQcUTwR3ksrzwOPMG66FXnFqKDOKpe0Xc5v9/Kd4e4EFBKZ/12
qlBFu8YoDfzkvLqRPAXXDV4k5eyBeTPcD7BaOyQDvS9P/ZVfrmHBIff0Uc9cZb4a
YrySA+5fPwurceJn1xI9xdyx0c9g6pO28J/ZRglVkrdjyp/lr+ugFWDNv7jgFpaF
u0y9qa1el6ZZE9Sh8mZeEof/FegrpaCfn9Q69YsH7NkHSdJ5hibf3Z2gjSyAggQD
+K1epwKY6HkUwBBmicSsaLIJNSYSDelPe+GdfVus5Gg6FQcAkHjU72fJZDwA+yeP
6UFO0WACnlwqLHGzqTSqcoiGb8lEBvZ2IT6Ur5U3hKK5yM5rmwwayFR/GUDusHwK
WIIp91WUTOztdbeXKPyjpYL4yJ+QnOjY6+2o1pG0lxV3Xsh6MvkQIAt8NYpknjdg
vlnyYpUAts5fHwqbu4Hc5caOqLFarXHQTIiZdzERrTQGeuu4iq0lcJ93x2Vzkwuu
rEvfGT+PxKL+9drIagfELWzNTtauT18GPrNel2KsupgkFn6e9Xbw0wltWNWjcJSl
ytMGGLylMrrVZ8wuhstH7Ehk+vWN75KCsgJiSOsCDD+H50AbhJNQksLy7w8qaSJJ
sjSbH2fdvMmAtRfuxP53JCX1E2KWu3L0YVacQ9Gec9S+NjKghCGP58IG1RXCnfUB
BzQs9GyK0UMWOW2Ox/m9ZlWSxtenE+6UbYNSWPX9QRlZHvwl3ki2W3eZPKDQjNQH
5zyXDjemP7Xc5rEI9Ct3/dvtN2qVcVEMrVh4//hFfiaq2A1+XUQ/Ym31NW9kWlZk
z7jhw9w1pUcEUA+JGLA3QmuhIkVQHer0jJfk9d3UQbpWhQvwQIWW7iEsfklHjrIj
PcDQY+iUGXzbn5K/FDPdvj5QM6IrDAdzNvF+uLJpzP31DieV6iIH2iGnUJ8Wc9J8
kM9q4QWXHEZymyNrdDUsuKt3P/fNeFtu1u9CZc0zMYoT/WND4rCkO6gtppl181u9
A4HNC29R3kpR3KbmzjMQKAH+TsF8KGIpx8JavtdDrYZlPpD0+LzZQJC1Eyxl0rnM
d/ncPz/X2EdTU/HNaxy95obYplomoA+O4NB9Gak/l4/POvVe38z4yFwvatDkZhih
aHfMVV9qsjg/Auz7ant3/Z3HaTXW4bq/axEcSivrdvMsJiO20GrLvT+9ra+UABOE
EZUe2JpHGWtrfsbe6kLTqOoVuWWif2Jz/5InwAL1GnJaKXxRYthez8Vj12nBFYEw
VjCU/miWKQZL0Axttn1EP2ZT6/dhRRAtvb3pogTiFQ+Uks47Fue9ongfXM8P6Fqr
JAwt9mmN5yYOnXe4ODNNF93NOt1fyyoTw/TuK51cYGjO5zRD1FcDtkmWaH4cg3xe
tb6pYpCVHe8+cXDLoBD0eqL+MtsAa4jpAV1o8BYTTYzBZddik5F5AibfkGrT3E3e
ODOllHSB2d09SEm7t+ih6QFiN9jnF2bNamZSzjUjCCEiAZfMN2NqSHCuhGWKxxYN
wYH5+OvTr4Y8PbEn8PHV/TKAe9gtb2oHSNgTtLUqaBk6kzWf5Du9glTVntVuu+1R
Si1RfkbLaSijWI4VKLu6HGrLu2BA/2z90I53UM+fTa2bmu81MTy2fz56Bp4bVh6z
faMfFr2ZQrN9f8zee7M11QxWKTLRYaxQOnwBd6goj3fw6rXrwye+G/TbOdGKpupj
dKNF4Ny+C0Xak+XIG81cWHvWb1rsp3zAu9edT/SRQ6ZAKicixexXoDhM5DNElhbe
r2Y/lGZeIVl5BAS3Pqbley/lBjYHCjSK/rwqto2C8lxNeKbvX4DVe3xyhpFcxyL+
MdVohx5P5rF7/wjTHjQmfUpR/AbKlRP1TSt2PQYCIrU/xYPQqfVJv4ZyKtLGU192
ijMdBbfxYgtBHqq627zZXNgtBsxci/yR6syc980TGmC+E8slGmGSu95UFdAlUIUS
fIsQOCiIbdgRH1ZeV3OGqgs577Q3/W40GmVPAOK4FdO7ZEy8gVpXHqJAprsiwmwF
0icq67DqVzbe7KI5G7wCvHfrQSFAUmDIol5PS8W8qP0k5Q55VfL79nH94tlE7vCH
ZXQklLSyNWK7kXhWgyOhLN2iiymx13AzLRsCVZDI8O0hMpo+FlOaB/m9DR6PX7s8
099OzTZO08bsCx8XarHWds6I3hplEB/Cic2iMV9qw78yL/4P2Ku9+92RN9ZRL40N
KIfjwz/3TGTrxW0bNE1KkVAlgor1v15ugorR/GbfouxKPod4VytwceUsKfSt8rmd
xiXHRroWTeEvwlE6T/A5nh9Nri5WueXSD1RxsDaZTK+kTYw4xPAZ86832iphSuLy
EO7Yj5WiSgviLWKQE9CofbUugYbo8DtemICavT4SQP3nNyuf2ZIcyr5t1u9TKPe3
P9j3SzijoQlRpJZHmSL7Xr2qPhSUI1Ojmt1EGPMfrTWE3Gv5LVXpqdhp3TF51UDi
5cfTbQJFUPj/lWzxJwbBeQ38/RvV1H5Jf627QAF4v/PF7VKwpSvkZQZEorbaEQIB
dUCE6wI9hnU3Cv6x+tIAUzqA1DSnNGIYqp9W1w3vI4In5Dwh6XSE78BHtESbB2PZ
QfkrvjCOmUlA/EzDZVEhR8zKMizVmRa5O3a0vBJIzwmin+8x6kkrF+dU4lHfNH2L
fNCOsev3f76FghR7RYAqzsZiY90m0gdIdHX9oaEkLK+mRYIQ0IMgXOJjH2W1WGbZ
BoGsXy/gOGrlzDbpyeKZJVnlgrQye470/OYEImhMlizTC0tR+18A2OyHiGIxX1im
AuHyU6ZybF2NuhaqS8o8Z72KJa3MEaxZFIgyywNR4dTzs0SY/g/35rr+PbQ6miaL
tVeES4DuTMEl2w2RBQm8dSubl1xJyQ5AXO1XlyVKl/WTx0hgMAhOO/hiD7AJpJvb
rRSQ9Qz5lzUKNkA7jk88BLkYOumDBlEFZWkTUWQech4TjwNSorvxzctfWt9xeLXU
CbjNclX6YQKGwGdMr+jzpYgwwl1DmLOdfuKVhuw0mAntTPKuO06t7l2YsSy1fn2a
eAAmuFcp+YGkolZsaZn9gSHn6mfvHXLaE+EPNjd86nM2n5C7R5Q7c9QERWZ5XMGM
MF9DQwOfCFq1ngvjB1l+y/wN9VaF6sHgN5wlTuOzttGAhlCTXhAbm0scNtLKY3EN
INcR+m8s47QJ6lYNOeKuC2Z51+F+MhgKzkYZ+3AcP26uzm9wh2KdISBo06Ab1+IN
vGCfZYtvTnlXk68P5xdJSJXEFlFNW0NY3vwzNfsVey6vfRcBVsM31q5eEIeiH78r
KY467A0jGOI8PMBikkR2BuYg5Wk8XxogQF5IUIDFaODiLwRnzY6TpST9hHb99DQr
p6yuzU+SkaTRXSRaMgZO801ui/MKI23ChmxcLVsINVHoA/nchcQLCwnzz5kvAC+Y
jK/j6r8CapqxMMlFbV8DfIhq5CFmy9kty0eUWrA3R133kH7Grp4PSDIApfT1Jdyx
zTh3kFeO7NRWoWgRjWIBMyxi4MW7o/tB2SEpcAY48CA4t5oYuMLSbXwBNaIzBUSG
eiQKINbkZe87CTgvS7kfgkIvp9hLs76v7Pg75+nc8XuRY3cnoNhrRey3kyfybk5L
3rw0HSoiR7utv8giqtcyMrwUE9mJZMffAuMvW96CMkGRJYtwFsna8/ATASznhnza
m368d8SwrDFRSCsOaf0nPtLDindJGs5/6lD01HHXOQsLfoZ41hoJ/j313bkJqyap
IDjmcX1/clX4me7waSrHGFC721w2mlXu5WEEbfy5786BIOFDxvWX8P5+CMTJ8Tc0
oHMOpfUPL4DoWjXOMwAR282T9KXFDPO22KZFyqpSI5tkmalsXiXxeGZ226Na5fe9
U73CE18uecg8TFXG5iR0ZjeqYfJHpsEyNLJa4+OthaGWMBajSxT1bKjUj3/Ic9KR
SrVEkbnBQrAA/bw2eY5OgaPWWXav/SvCNZZiQl1MsaP9BkhvKhU9Est1gDJZfCzf
kiu8pjXse0Q2aTICq0kmd9fTfdHXE98K4hIjfN3m34mmfuRkpmivS8V3joBMhDX1
MKewlhQcWKDVi1ilh19qIGSffOp1dYKUf7hGxErqqpbJSX2uAU2NglDnyp6UJ0hR
pflGXxSfXPBxzECG0XgiEhix9+BJ/PqlJBMz3RFvrJg/bYuTcDY13Yc2iVbEVqnq
CCY0ZhvpJrh48e6n+TZrld5ba8OVXcTPINnvq8AqvCq0jJ1CRkgCZeNnerGmdBiz
YYjdd2aVyL+MGZ1YBHdQK19+NhWm51G/gxLL1HtLhL2rBsxrp1Ed9R88XYUJ1d1g
4wYFSqIPU4lE0mNFpt9SPpacBKScrWF+AosN0yD4CCh+Zd/TUUFyQV/9AoF4uMo2
WWlmxBCY0nuRUP3XCoNhgjZ19uTryr3t/7AOBJsmAPz1PSk4mu0O+pyzcQFio+Pt
nFCQF4zXtI0NUzg/nQv3OQxYL9i4WfeRnRN0hwQzh8AQU+LKSPVu0CNhb1oGV0LS
2zpaVBH5NmWuHF1cJ/STCl+0frbi+YkiDd2rzHEQz1in0ZG0lQ2mo4Wm1/kasv8J
H5HzN1UJjmk1WwpnNUkF2K9i5Z0rg6JFUiMW2sQKa+lrKayTq1z8Xm+WnY0E0nPN
0PZ/L79EnpZP7zhkEH9THv2GUwem8bZC84E3tzQAOyJzANfPJEUOl4afb3EIdU3X
dL1pGs4hxjuDWZugOxWJ7opD0TaimbGVS5zsBeO8/kUXMGs64yEody8ylOGg80gp
16EO3qYGbDnvlrQ0ZIM6UNOO42R8vAsM1yh1pYwIVLIBUfKCV/kTqop7K5z1q5Ft
swUl19qbJMgFlseSYYWqXqFIdDhyMnc8rGx+B0TRLMwqFaHrX2Flr1r8KDZ3tADE
cs9ZEyklQxJuUyuECJXaGwxfXB9MHhANk08eZtHyYcHIo2IwdNLdppHE8b3rDjuj
v7vj+f+HW03QJIP+gRIX2br0SwVTgkyEYkieI9FViypl+fiCkOd01lmEG5aRUt4T
hEqUKysSsLeuyFS9fyTe0AheQ2O11ZsJaPoIANiZLx0fQ/j4qe9uCUsRDCmP8sYI
KiXbNDAXJxSrZv5V/8YQ69wNSO6RqBI+33iScjqGMWn75CzEVMnKPMTnj8yQ26Wx
CrdcFlvDck27k08tBrDvjUwrYbND/Qiba0wLL8JXJD0xQ/i8dFIwIim7QL9uhj51
Lw9qFyfV+B7H0vEk1+mKiPm97HHupHYhdfO9bf8aaK3HnUh/EQNV6GVz1Se6hR9H
uK+p8KvS4+P4nYV0ZKs8e+VW7TQ1uz4L1ARchGRE55X+RREM8FV2LitTe1fA7QQT
oBC/P1Kw2rB89Jgkz4rmmmu+lDVCu/0SQWL1JcQIwMjh8BNtTNUiH6/KV08U7h3G
vDWl4Xo28qFj2cu/FqNKzXxLQ1HRULKBhdwiQF9BO1HxCgLYJWysclp078p5qzmX
zcf/LwJKXpF61Ly/xgv4iHEVlX0wcs4X5rrB56zzLTA6GDhEzizeO+5z6Nbzi995
5D5BiB2bycmiADpiiukZrOHiBxh4vy9DiVv3rJ4NCCG0O/SPOCV+usWjdibHpL3P
aZTlU7BcEwmI86Etfv/BMiwwTlAtMF6Yf8zmv8uvVSxdwF0avKDN/oc4QDMrxoHk
6eVAvyU2RtMzmw9UXr+QvkGxpTe5Heg+m0uLCbA38kIEvr0zoCxF80JzX0I2zlNk
vy1NxkBfmjTck1zN1lhVLTEqn1OvtXey8ZXAM4zJ4XgrgjKeGbs49zwWpRpFtzEc
RcaXTJSf0Qhh4/qIJ+WYDzgLWoevhG/cQET5ysSuFuLzYJCk3odZxdKKAdxrp/ba
Zvq/mAlvBgakCdFOKpGB8Ld62d/zaYLBx2AKuqMyQzTQYBXMu97ez3XpzaNcLVEa
YseZXsqwcMmG93agyEVV3LSZjFMDf+iEf9b1nAHrbaGsBqRGBmo8eLYeKuFZ/fUU
d3HvEAkwFX3+tKxpCRJj7UByB/Zp424ZXyv0CELpD+XldziNflSez4TiFLzouIjM
+enFsvMgIJh+I+FkHrfJpWU/cMz07q7t8KXsK2oYCoUWlILXHXLRemxk5axCzh2K
pfdUNNqm3uch0fZ/ExgBbnf1ZTDNIIGvw+5h2C00PRQHuwsAvRpia67ddmNRx1md
ZVE6YNJfgLzjX+aDZo/GgEB/wQVOvXG09s85qMjBxPq5seHgtlGMWOHdxr/jvw+J
O2/tRIcMu0Bd0v+mvvC2VXUV7a9uQymfORAE/OeFZEBSlbX9ze4PgkDv49CQOvIA
P38eOK5dNvj4oimeV4jZKlrfzfJB+9kVdiY5E+9JRcO48xICafoJLL3dleBaSeVU
/tH6zB93j0RmLMoT4Gh9ApaOyHg77enidBK2pMePu9iBYHJRA0RrLDnBfgN/+3Ky
BYbYoRXZByqiEg2Z05JowR4N1kuKD5wtdLwm2LxB3Oj617pxbNwAC2QVvzMrxfV7
KyA5eAMG46f2t9ismGVzfkASbq9ETPuhyXyp3HQg5inJIl983Pdb/9kkiAWDQsJu
sgk7ykE519s3iGbQuTNL0SXn4CsCCLIYeH1vyfWld7R/ijyAZvofGZuYuR+WmC97
RjynGmdA0Q3qUWAfKwov7u+5FzaioDCziWAbRUv+qKPEfCrmGE8Ei0/bJ5C7X0tJ
vbfW/y01UZPlfW5Ye4+yQip2E03fPUFCYekoto6K3gWF72uqUiGE8Pn7wAu/+0ar
4IWFEimoCz57oPRo92G21esyrpPtgbR5xX32X1b6U2XbRSiUjN5OJeC3LGmx5i+s
UFlMKCMEQL88JsLbeeOuXFYO3wEmrONBamQk+OgdkWRdIuXzmF+Xo5O/2sziLR3A
L1DO0MutVkvv0/tAaz6T/xwq88ZHDo/Fy1nnfRpWkqDxP14YJtxIJ4J0cwGaQWXm
eG+Irj+RBECMqKFoMhjoMThrT5kbZZuFHRhV5zX3HuNQjB7hTeiUZ3Ze6vlyDndx
A74dWwXGhAZgdq6lFeOfJSJJCzJZhyVHxK4MuKvabkiWWSkhnpnU+Twre/SLm2fF
lCG0xU2YSk3B7g1UqeWg5DiwPiQEZ7FL+uV7Zri/sibATR6f4jh0+RM7DCHg+rWT
Izb9dT+3qrnbfH4CtPSQwXhd52BjzgT0xAUlZdlq/I4qjH0TkHVVSipYpLx3FtD6
B9Y1G0GFaxNR2vL5yTqGduaaShEhU109a69EwLYVBo0mAZ53xNZm7A2qgPTN94CI
VjBYof07WLM4wPlYaElWoFWRw7uoAFeOJ4Z6edRRxCx5nXmKL4IGKeGU3HDRfvhW
sZlMFxwSHVZiKGG61ysmQJIcAeb7rUFfVm+cn5V5DsNsQOoGyOmUHC8PpsdwNDie
YHXo7JryD7nTkOEB8ZOwO0B04gcMzK6CgTj1ycUrY8AZ2nl3JPuviOgBVwhJhrdH
TLskjxMtLZyVu96eooF7qtGx+9lXVviGiBVLwoK/0V+HJyhJvFL8woI3VqbrXmDK
IdzZoTlu/aDY2s2CVJ1FzE13jPtn+kBz+311esiZcMWY9rUicij2oELqtFa4ZUXL
tNieFSLkaKUO12T6zZ/5BPzUcefyX5M9EB+jYTwBh/DM0kL2M2ejv+pbGv2YFwG0
NKD8xmt35Xc1rabOnohgaK9spGqT6j5z/1Ov/kQ2/xlxSQDWHddRoS00SAHiDNQT
pXJ1NXBkikpfLTUDC9jwd2vcF03eCvbtzQ1KdFu/xNqiUQV96NlhLyINip7WHblw
C9Uzfao5z5SQFiQppHJFwEsGwMmZ6ODeijSQgx5tY8RAyEtDTer68wEp4f134onK
OdG/nw0w5GY8VanmkxpMTdizGuFvfUYNwP39TexM4SyQ/dNhJZi1WIsWikzHH/Ro
lnSf8R09kWGb/YMbNVun24/WHq8AqJF977GT9yNOpKe9b6bQ1ASz+Koc4157xIMx
p4yq124Cuhj4dlIyUv5ZRNCZVnniozSPn5tra/uxkMO1nGd94Eu5r/c9iebZi0LS
PdtAkav8JftZ+UMLnecgJJm8FQoTkv78mi7K56t7GaD2IuIuUo13I9lc6FhG05id
n/9+hkY6rSBTioBxliw8YMIF4Ax80m6/xnkrKKNUzUWbjJm/ZJ9GGa/k7NUOGTYQ
4XdZTr1NtAkiaRSJ5sfOH60YYu+qqEy128o8u4V9qhAeyyla3wdnEMlKO0L9VSLE
/zf+m/mhZatbKx9uOqlWYK/46yYiKUhZngeUPJ71fYglPGu5hSSNDGWcUvRc2Jcc
PMOEUQjjnIlrxjTjcEKpPwwL28nbsW1Hp+rlGsAmGk3QV3AWoa5zMCTDoefX1W6r
ccUT4L0QCkb9IqbmJVn5ROaEAW7YK/vzeUpvWECzY1JwVs4VorNn3+CmwRJb64iz
m5DEfjrizhpdNT7spKMRzxKr5/1upV8uyOSAnB2cb+o0+uhHw6hRNKyPDp3JhvQA
+9byA8NGiHWA9KXS6vxLTpLGmqvPoJiGJkhn86RXatmO+4PcRa5ZO7NO3X/yZB3B
uXU3TRi4NdJVbEqkwTr1pSmVf70Bk/Bu84xzeLbW+UnEqdIT7cxJ1nofw0thZQAH
i795hbd5oYe4pAXjAq+hwq356OM0k9OpzAdVsoP53hke10e8THHllGqivRIcAsfB
wcPD5S0gec1qm8LhYvkkG0fIqHCmpzrem+Nwp7mUD5LYgtF1CF2oK2pS/Ug41TGG
ST5qGYeJ3AWkpgJnECcvj3EdMVV9yiwkeV6XZYPWqWOUySIbPv1PeqDg6u6/8Hgy
72qpD9rqvJCH0PnJs9KqArHGbPoa0CFSBxsuNVjPFX0poMZIvXWy6cTu9mBLevZx
e5H0uNOyhvb2CkTVBAGXoKXsbR3EbZWUn9rqLwX6A7Od6npLhySjfR/2POn4g/zx
6bN8Y0P6xReZihG8GT2zI6P4iELdL/L84qji0PdKGoV69RZS5RaDrtL/wQmd3g6B
kOa2V46xAirhnn+fRn7naNKTvVqrRVZsloxFD2iMek4Wa4uITdGz3r0iSPB6agu8
RNsXl4IEgC2R+0mbv1Paxuc1WjZZfYjmvyQsONmxRvfEba8EGIBsqgi+yokJot5u
PAt8cXpGjgld/l0dG1zMLSJ5li29N5xwNmJWvD6ZSuAYIE4ynrLzA8kAHPXB3adh
ZUm3RKGMtY0J6ikQqFUPiGzTcsj9bKx1xP+oH9wYDhGroHCFxwXqAmEzMtZhY26C
Zfwlx2EPjMnbtsl+6kK0uiNtvWgsHoruJIXJ7mLfQKYKsGpExOrIquk6+yjmuWiZ
W9ZQmFWma18IExCefE1tJczE60x4fAq92AElyekce2iQt+ZVmd76YHYR+yTUVpP7
dOdvh8dx/1zWyvNa3mLHjSGQm6zIB6wKzx4G9YTIurXorbGkfgGfDzBYh1XpMTFZ
fn9LFRVYvplzepfVM6Up8Epme6wji2utSH9hVKn6VIZDxeLFLzZc3tj9YYZgUO/p
Sd0U1gt2YzOqOEjrNdV4m2+2ClrmgRUkYYHv917BdYq+zB5bGNjm4f58d3MZqoWA
CzZqdrQYJUCCgos1wDnWgczhtfZ+BoDYZfzxAzthPc6VdRa8SzgrWp/I9m9hBL8q
qKtnsgPyxaD2y0/8C1zqhiHCnUSn4qccjCXpQLtJJ+LlrM8GnlpZIMAbyBHTw5qw
Et49k59AGFMNQSRZhg3S6jAmdEQ926GHs/jYtnRxMU9/8xCEDGbSWLwkoIHPfq5s
VW5MsN5Qr10A12Dw8lZNJVdrNWTLJB0QF9rUa36jzU8GUNrfYxKo97if6LXDKLoL
o8Sx2YtcQieSPAR+C7Srl+xP73RtV6Tu34rwRGsxh+5dAhFoq7idccKjpaV9FOvy
8k2/oBmMTRHN+5qM/Fi7tATsLN0sjK85I3qkVu7SSJinLTUm4vmoKRYUMKq4RvL1
yX3xViBcTUgFOpHXb7OtROPpLJ37qHvjkDp+/xBcrQ9IFQAx/2t6gsuBbp7Wz4CX
gdeyVI19pjta7wYTLYT/6xWprvjtQYtmFK7wZDEOnEf2ZuzWOMXeMa2g8K7F1b4w
nFcHvci4JkmbyhYOro+g7BDavLlN/DVgrFkDvxCdFAar1jJBWQHG50cOJIppD4+0
vTYwP0sPNzcrppxeNIAvvW4n9EMV29LYqO2rNUJbRALA8L848itMd8oKAxd5X5hH
l/icMtqdrrdDCmCeOQN4/y1n1tsBHrlJ3FInaHqMTrVGyQYJD9gHjfXg9nlkC64P
G1rrNqLLBLqZv2OF8JCdlDWh5wJrikn0hdG2bu8UKS+pLca0CP/I8+Ey0x0JXxOV
l2VsKCEU6p5EM1iGZUzy2pmwi8ph75lFfi9DgQPUZC3MUkIxpbeyhLIKcUzgz9nO
VUg+05jv+voDkJL9mewkaKn1o//n56MUbNhFfDn/XHB+2wKkLRKQ/YCZIm0RSDUb
ut7WGg+0nghftmuWhimcic3bLNSDlECf3INW1pNKrwi7kamBERc2He1I4g2C0ViW
6XhXNZ7sUhRcsKGTHaWxupJ0nougPpn9B9PNBiVu4eH7nQAWmcJKrxKqRwzHOlj1
TcFB0jicxLcJcXiDHiTLV6Jwzu8p5lJMVMniMv7dheFhzgrSJ3evBLKKE06wMuXs
ZX5l027wfieRyTKkRLwPOmkYMuP5covtRnen1I3lSSjtzS0ASMtuTiPMXPDpvsqt
4Gk5nkQ5+WG6Swjdms2pEezds4SVGn6kNZDviqRBTqC7+Pq9wJvxht/6gzNvRZ16
98IVMrNIMuA0HIble2gkFidQph4ePHLC5jSiTaDMV3tzUOkq5emr3KgendNj8KTM
QkLqkfutQk/7oG9VPORAgVzVfrmczxT5DB5Q19eRYnU9bt4WOUlL/zlqmESJmCvc
GcEnEetA9Vg/hiCwOcDweeUleg21pHh86uTUqn/IYYE+9R461FIVXbio2Inzjzoc
ukdyjXrFBM/fijOWJSCvW8TWGSbPOobeyVpllypW9PweK5oRCkKQL9VeR4GciQV4
QOT+2yAVTn+5EwB7H//hGQ8RQ0KV/ARtWdGue/WzR9JQbeuToBrOwIZqOqh3NUCM
lI+BE0j7SNFFRGAHiN3iP5+nhZc+v2UYJ7xbXBgQSsRNWU3LedI/U7NW3aq0M7tK
DtJOavw8zl+LDHXMgDbgqMY6gUusjgI5/0t8fy2K3Xxl++u3EUuDtQNpAn7/lEHg
a/pFV7iMQtnHkTHXur8BdfYD817csq4AdcnDvyIwf5osIQ8kyd1n4ZEi7Srd91p0
hJng+u+HJATidUoGcIfIZupqI5WLBdfIJqfof9FlLjwvfQhP6VR9zN6tA3n6s5Le
V0GE5RHTw525NAw8cF1X3moPBulavTu3CQ8nFOvK4ohs9+ms5YFuXLa2LUc8/lz4
InYttwSPpVKJjKiTm65j7HfuOa5o8uPy95KeWWtrnJkrF0wNLf9wB+BS5n0lkBcE
I9g71I6Y6lpmtWwHHb/mjx1dGWFyXaEwgdzHJR+xAjYKAtfFKeQvubpQW0dIsARe
e33iYfC3z9bObqv5EJhZmktYXvXDJ3LwpLGXG9NTkouz79kzIe1G78ukyqo9eEG8
zSVw6vMz0nhe1URdd1/tgbKolQgwR7xfDb0Rd8YeTRv8OkZt4w5vuo+p6C7QGhLH
ThBJb5p5IvJPxFgVE10SGkwHqD7QGNAduWTEsUYYPAVkYWdwvQzAcR9ktCoJpagU
JozMQYsUXx9enn/dQSjlRlJ1TLCb+ylkEKulJhx7vXUhMMH7Cw5XiHVcIi3OdOhA
ZzMvCYIg5sQ42C4mCEtc2s5LtmvA6FEhQ+6bIyvoovpRx0Z3bbJj+TCZ3Ro36NYm
OEo4riGN/JU7fL24O4XDYwDhctK3kftl+NyoTCD3QQgkWJhgTWVu4ZQe8EDPunHj
H+/81R59YQP0+L2zX6owrpJR0q34BlN3rIDhIK8WV1Arsxib6oRWBuVclCLAgz4m
tfSr1aCySBplY/4QrE98n7X4tWUtUqDOiUnuFkjfhVsRLGxSMaweyHm5L4Ho2SKi
jOJUv5Tmak/n0zfjuDBuoHXPgma1QMYOq1glOpJ6Ta8/o2ADGRd5rzwnQbC8Vxi2
8NtiKjcnoOUaRHX8bqEoJpEZI4xwz/IkwRzBye7zyMd23d9CPZnJnRMJheZC90UD
aUx37y5LEIBzcSDfwric5KExdaszbe6LNCNvKy8Rd3SCC3DzKyKb1UsLhVppSyNJ
5wYYVISfykh/YbiGB4KESokSyxPR8mTDdl8dpZF2d6uYf3aD3itfHFvHt7E3Zj92
DZ6Bd6ANBZc83nKBIEA/cv2fbCWjghYEBNF6PNrR98IhXRToQsjyRq6DFtn+249W
LkreslSLbAXbAoX8kpGirezR34Q77eDOZdSqQ1IGdsiUCmK7EXY09jWbGm870Iy8
Wy4Oe0fneR8XhhL2jAw57iiZehSPzO6wc5PkN9J8LDRWDK8ZUDETSy5oRcVVFVQt
EmuEVDHXp8BrniUGjOBIb4puMpzU/N8t48TDyBxAv471IDo7n2RZEacakzxTxwIn
dEDfXR7jzVGhZgnTeoJLjGapuh0Uh/ul41Rkq9Hn4j4IustUrhth9urg1IrVqdCj
HReKl7fblCYP3Ymxd8IYYWG2TcDHmpq6g4I9vTLhWexwVwAJIdgHFhCE5v/pv+sM
5navlsB6y+Fuw2oXPDPZitzlGTCLYaQFXdECBqoj/+4XUOW8ymSIMB7TUPwzzvwy
FlTl8GYHGzqp0le3d0XQm6R/3EjDuE6a57vNEEX/LMNe5XqZPK6yUiYK2aXr9YNH
W8fzhh8sdRZ7fFiEhYl/x9KRjOcKjD2Z8ZdSa1budtbmnm78ckdp1TEJ0Wv7qeoX
AYGXVP2HyWZ7vnyQNfMPm7MY2mp+e5DtqTk9kWSyyUzJ3Y+GmCBnmaO345KrkZ8E
hTF1ebGv3TMBLzKUE1CcxWhK0Cp6LIvR7YvQ3X1HO3jMM44hq1mokpNjFaiwR6pp
2OPXe64p5Gf+u2LhUDk8yRVNZFa4/np47iLwiwP8sWUwMzp/9JKuvBEOLvHGt/c+
0ZWZJRqk+qYC9ngHObfgLsRzjsGLTiXUaXAG/GWsR1Pg9rQLFVgJnZd4F9YWnmjS
WpV/7mdJhgb+EDgb473PGp5BMuWkA7XCp4HkEcCDM+At99kAu05DaOSk7NeYWgAR
Z2AtQaSJLd3Zx0iqCywDmPtS3Huoc5r9xoENVySHi1oMiMr7a8hX+eKu2kjLZy0t
CVhNiZfvMAkR3HxQLD6BZ3yklfI1B0I13yJNtT7LQCMIGzrS5vCcSLwtPVdhamYt
IYvCqt/mmCne9eN0WiAm6KodLjiNSalfs/b0lYS6bOA2aflVu0sHY88pGaRdfWp6
4ky0veRlG0WeXi5XygLFXGPBucxYPlpNRs5p+9P6aVIsEjvrd4Yuw2CeAEa7f+mp
gHskNGRUt7PkzjyRXE9iFlrXtQ2dmaridjLynRAeC7XA0R/M1EMt+/ABqmqrH8cZ
ymcpJAj8AruiHGDgGeeFt8NGTAfJpWoRNXsh+VZMvCwKdsB0mhAgIMCroJ8EVyfS
LEVgWDVhcgNjXPRg+CqQiSzgxu6MBOzWz9JT6/wBtthiIPrw6Go3TxB3237OQOqt
SBhd3UGmDu8O97NMCe2lFWFF5oY7fE7jVLH0dXG8s6WkrZG8EvKmiYEkZc5veHn2
MF8BL+IAbzCcSci4K24dB4JfPtgkZgafDT1kA7HwJ3PfJug9jv1DdcHjjNICq6ll
cy90bmBI/HEkgRG19LKJ1aHPLtRJGXpYcICGUEGaGEJ5CzrQkCIv3NQWHFegON1R
ALyqXgw3Bqw71rzzHjIYhcmP2YE+tyOeijG9a3NoiT5xvHM7NeCkOtCgKJZRH3DK
D7Qmze+pNcu7jwyMZyiyp0zjHztjj2aOW5qgvSKODwesImcXg5M/qVJ6eAm0oazT
JOoPNtMOAgnl448VWKkHAObRXvQ3HRdW3OYXOK2h7vC1LrKJboQjvZs5IcHzpCkS
N8Ixn2kI6nSKUDzZ9FyN4eYdsvriddNhmEPzLBzPMNnp/CCO+fS2CTBLYWNTnwZ6
64v0Cr/s2kcVCY3+uga/Zbr1wiZVWI4GYD+CHfE58Zy+YuBdggPuXwfvFlK4KXqE
1jVgErvmoabbbxfqDra4l3eDhQ6p5yTrDYigU4/dALchs7eA1u4zYzcGNVl8FKSL
FN9jmrLoJdRRwZ2kNFid5SEoaH+dvnz5zqJIv0VeEZy5gnsRf20H5znW1KLcRtvD
dsFqgpN1bZQaVNdP5ySijBuIxepFBcRt4ihl1bmiAtmYOW5k8Q5RYCy5iCsyCwFr
1ZuYFizlwWgnyVSeC+1kpA+l6Kg1TYNGZqyClW8BFz5WUhwwGHrND69NfxYd5WaS
sAQ5pyyvshP+SjFmTOKXThCHBLNoxXQpTOBzkJFaGzMT+G5tRCFXAqusix9SJsGt
rdvhit81IUkId8B/vk2uiOAsq9CX9r/53hAx1R4JznZZqjraCTIP2QRTnAdu3UJm
pycix8/As2uylB31BOQ7SsYeIsHLSPAF8zP7n0eTlVSqJDwtYblJ28m+/V+6Tpod
VTOrZ0h8en+G7HVI9McVCNAdWCEuXdO4lI4CgUfKYxrDsLpYuo2Q9AoxxwnVRTIK
fKFRVJVRh+AHm8VcjHawG+mCOpDjQU3cW5fyZco5j843bPwv9Xiu4BijyDCHNvFT
7G8236F2Uv5NTo2BRLMgRxtqt9yOuMU5QdcC6ZRPk0cX8JvHc7YOJEIx/p+VLYmu
eHJAtl1GA+woigHOvn42s8fTD5GRfQTvtwJ7MPVG8DYtxIbaEbDCQ84G/zrU93Wj
GFYay4AFhdVQE3YKQNcNqMH+3MIsAkFmLJ9F+zUBTvEk+DNjl3rpYBxdjzjnY8/9
VOZipzitE//fwbdfOMoqgOiqZ+pFkHZdiclH/OrhhfxILOtj6YxOon7PPyzX/YT4
HaC1i41l5QhfOaYOONnwFwQ6PmRB2dZ4Zk+BLhzZq/YqRNd9aCdVMbVrUfzmDOeA
J/F7yaXtCcZIMTznn/Mz5IRJuv4t6JaYbyHXtkbg+NesVzQS+m2l3dfq6C5BvQ7G
+C1etnizL2GUlOxOj2YjgXOmCFid0i666NqyxfSS8n+52sNMa3++TAB8a1iYxfIh
vaegDRlGUws+qwVVzxmzcANxZB00DUJe7HVDC6riieeGeZvZSMzv5EQNm0tKNy+l
AejujySBDR4JGSOfFBwENjn7AASHJh6+eggT9ZK3NwLZIrNdVwxiTt41tey3coeg
Vg1a9x0j5yWNWRPJd7vXCsFlA/15jUeR2DmCi4ZSPRqa9kx/d+sHvkziOn9G+NLI
pPUENjIHR8KY6G/+owYr8M4E115MNJEy70CANpFPp+GZcKJlJ/qCDbvmId1i7Brb
ZTKgB38quBsbWyYNLUl/Ez8BZEf47miUa4fStMjSaneiYxi7nFYu84HlwSa2+Wi1
+enZ43PSfqC8He5qSzJMg4+4A+dACQfGLewSrP/CH74tiqhlR1PqBzqzzPWuiABC
/Wt1dMlSLSed4wT0sSkO1nfUQodgOZ2y5D++Gtf5waEIGxHkM+bGcQZv11iTInyT
SztehC4L6oYnkmG9CB42Vy3cKp+eYSOJn3dCkrxoPOdmT6hBJcU/N/0+FGnNZHC1
EHesM1c7zQm29VuCeNVvbLTfp4w2mUTNmNdTM2Kj75py+JcBE8mF7m85+KujccHc
TC+n6cINQV1xGW4wziGGHhbn0i+Ijq5VDMUbZeRtFQ2UBtdssKPP/FcNtaAPtpAe
XVG9+FhFONpK+pygnvDe4ioO3ZGpMNAAMrgt/UyxQ5rFtRWcxLjWMbW3sbxSNHmu
VHeFJmPnqr8DA3XfNYoUDhnKj44aXLZ4gvZg5/lY9vIOIxayaZbdyxFjNKJniyDE
u33oIHzwQFdWuct4miyje/pU4E4THd6NEleHvWFqxIPdSMlUvTPR9gYzIsz6KiKH
O9TEdXou2twZ5EQ5UhIv4d8JGSrYgvDXbrJzo9MMRbYqKcyxqkHrBwR7SB+C8S7/
RV2gNwtWb9BXVGT7lyw9YwfCoSNfPNW0aN9KP6QikJTAOcQyhcTSOj8fF5k9u3Nk
a0RtIthnBU7f8l7Akk4QsNycVc4ykJXv6xd1vCS1M07PLoqj/MqF8ymVL53UP4wW
V4y37/fIIiSz1kux+mkMmf22n1JhBoZFz4liyt8Kbxn1TJmEozM72bTf2A57FVP4
smGuzqWvWiuD7YXsEQLzmJ866i8mmhJGdmHbmizSpqnYPnnrDGooTHYBEYEHqcsm
htZqqIVjUJmAoSEljl4Sncyu0nbph5lUaC3VOha6c95F8pwYmfWWbOXPAzdW8r+Q
W+QjCoog67bKYjb0hRFHAPnfKVLJQmO0i7Dri5s49JARoCmofpMyxDT5Ps5dXPQ+
Hv9l5OBuEU2n+g/55xcl7s+bU765GUvtjbAuqOA8HJthhHo9grZYy9NrD4RrbRp6
CkNg1tmkmY2FuknXMf50mzzpy+SWYfbprgaIPEr38iUD1QvulpRbRMwhuaeaF+AC
LkuACHn0a2oAxrlkxb6UOAuafsu+5vZyZiqsbhWrY+crsmTKWkpKLFtBKmPKjlYY
o5124/+SzL+IZnTkRpIhoVgrCVi+6s92FYSSfBVyLuJl5c5HSB5KOgYtf8YG88cC
VpQcDK3DqNv/Sy7Ngf/psm5eu3FbRqDOjcxyFdlpuEaOzk9eVPpoB2yrq3ItHDld
AsX9MbewOwOBtbC7Lqn/CIG5/5TtjqkVU+8j1myH3u5atCrQGQa2CColbKHZIuI1
IiABgxBVGrijlhcBmh4y4nr068et/c0LLk5H3p/CcxyaFq6w6V35yPvu/7x6N5AT
gbwZbRhWiekg5GYn4Y2Y4nO69lM4SdNrHLy6RLTpCn5SaC72ITbBTN4P3eX0dhjO
IXDmH7+EAiMa76dK4bzun8sMfa5NE3pF178dTBbURNgxhAb2m9N+OFTbUt46vioi
vmrZSQKq1cwsgM9SCvT1HJ6G4Ij01eJn0Z9ma79wGK0d8m+mV8dvlO5Hhx1FUnt2
E9UISxOM/cE7Lk/LktFAMeaAouH+f9RXZCF8IGUEqUEVJwGRMtbQ8XsSBLSDSc0S
ZOXTdceAR42LGR5+15fTw35edEzLACG134C4nZAI/oTsP3RYaDPM+TrdT3sYMUOD
ZOv45Nng7B/fQFjs85t5TtB9bbMgN9sq1cQ3zMs3bRithjmFV2k86vaL2uM+yYHq
8oBmu0wrjpNsPn7xZsfHYUAnGX63yCVyMt0knA5zOd55Un5w7zpbSXeu0+fvac0j
dmEWqJij2vS+kzvJCmA15+VG9QfyiEcOmaTveLY7M/yKpgEz43vi9dDQMFNxT6RN
MxXrdLWa8ZIyFBnTJDiyQnb8fpj6drEwBD95TVUjiHrgd3pHuAkcC1F7NW0u8thd
xvaLMfIPZP2OKydks8iTCRZB0BLZnQ+BVH6eKefaQL4aDIZki8Ix5aeRIBDgmH3t
IgUDJAUzlowZHfII2loiFGREVNOElapfHTxdJsQU4+IdmZQTUNodgSdCscMzwpv7
uSAAcGlawFxALa+Rz8Dro8sxrKYvEL9YQwh1W47ElTAKs8d9R5uTLAEOMwM5fvh7
U7Jk5xiPESDuhdLXjD0lCjgf4BxTTHD/M2CfyxVMTbOvgGHK+MwkCfxFO2lcmaam
sokOcpKckPDQBkyuwibYcDp1Ugi1o+QCQkiVYqUbKvjNEERTGbKIexKWfBdMTrWl
H8IHY6wRHn0zNwiuJoiynNACWyUi77y8vQcmZFI/+Iu4pVKrEbLEuJC8BpXFKEa9
W4lWvekWBZqUBnHN5bDLoPyMByz+c+/nCkzIKiR5pypFoUacDW/O5Ijh+8jUjl0c
06lPxrO5SerHrQrqJSIFkOXh+1xfUSCB9iwPUuwXsqQ6crnPFZz31Tp8AMGWOhO8
FUy7x4mUKasmsd452dMNopBMgW/UAoMqpRpaBuCdXBrMf1OnrwzIPlHUF38UGol2
OityQue/f5ILUrnP6K48VJylYgUbUJTvJpd+HfGxmm8XUkP9mC4Td8Bm893axFvS
Zit9bSaj9mA+cTIo6szcno1HQq+UC0tqA1p9hPpMqVmcrbNnJ0nUZ5dm7cVc1bOK
z7beUn3gyY50iYl3yHsMeieLRdaC833GheuLcGPKsWnfZY9a8Wmzu2T39O9YjlYn
4Q/P/ylC+jqxvIQjvkk5rLGGlz44k9aPuOfwjqfaIT2nRN/8PGkb2/0DyCzp4/H2
TvKmtvyX6fAmDP+1s1rTNZU3oUnzYOXHpft/Gbldf/xm1MN+QYhLxaVZD14TB8mu
keyWcbAFf4GmUncrBWR3xIxPm7oXTzoVHfCC+3/Y30S3jP2DACQyJ5nfcjKwJqpC
EE4ZmvOoUd1x4c5ko0N31cKsqY7gtu8f+QkEd3NMnfRpFeehzRVceSuo0MHG8W5z
n6Y0f1mAr15XW8vBVZA7VIod9Wp8VScVGLrsdltZ66sWLoViNX2NUMunJyZ7GDPB
dO3Xq+QWJpafUnQJGoedOWGw6Y/a/7JpiuYqVlGaEvJLBZynwjDc9Y3NliA1Fztr
ONHMmDbIck6XtmYBNWC8gkc9ha7dupHgBs+eEVv1zDQ5wP7D/EJnaq4INIitmMtY
uv/MsqxS1pMBdHOm3SvhPF6FYQH+rfwqNAGl99AQMh/McM+fcPEmLXVksZWPPMbH
LBsufiLpxf0aO4P1g53sjAv5ssOaRQWXVeMVhqfinuqfkWcSWnih3SwycUt9Ly1z
MsijXXZ4Dwa+JZVVPRYZjh3UFMYz2j1CyQbLprhsQcYhQlWbGkBvk9Wct+2RzeSf
PX8v7kKKi9nHm9rRL1AMWyWKkLzg6PqefCW4JybK482ALrKyteNjkt51gUdUnUcn
9B1pzvYTpkfY5yFrzina9GzGmYHWLXbbWvPZ6kgDOACDKvxSneNeUAQe0RlyHCBi
4W1BVEbqPHhjyDGghazTpOLkWZdl48l+8rTrAz5LfwettJ9AF60aw5PwPgiEHpMj
1akmFqHcGZFURpg2ebG7MHJGHABkoprgfZ7RsUwoRvxkxZj32wVbjzdeFfgngcFr
HsnZHGvMEsy8dx26ffGNBa6svTIHQhkLatG1Lu8mtXT0LUHDadRuWe09l2IH6SfK
n3xYSBO5EACc5UnH+3WMw/c5D1lnd557v5KKWzIQmHOzbO2inPnP0WbFNS+1mQwP
NWu5c6vwU9nC6fHYKTJtYXAGTPRyanIllG6hOTlUg//u5SpYp/Ue74ngWwzcmZkB
q5sdDVmvTEMqhgctSRe70f7TqEKKRVnQtVfQ3FiveAiNgyLnzDleGQKD+2PqnsFw
o5Fnq6myBnF+D9XA0JKoYp2p0nVg81oQHL5Srr6m98aC+DFuSIF/yznYcydQv+qX
IMEVFyMfWIKPmZgw8aOLRrYmxswJ+aIpnumPHqnK3UaTvMXXDz0raTdCJGiq0yoF
Y5+CeEwJWnJ2ZGeopNbSg2UXuCxcTFbFfy9HqiYu+7mrPEF8W+4wwtssO/3mtQ4Q
Q3pQqxWMFfxof4roUuNbhL1s4GGOfNzoFwPRt2KMk7X6VCYx5PSEdJuf9YFSGfTL
44L/nr5lKLc2kiI5OM+llsAM69TBVbIh1MJyFRxc8CqfTbBI5o1h37cvZsThwc2R
WN48hupdZbEd9rcYG6IfGAWAqv1EUnF+PblUBgtQeZzrs0lv2d6Q/sgmFZSGa4Rd
f+pHTOvzPysKLZfrNqvZi8Lv6go4Kz9WYSlnCZIuBvCu0gpaO3nIbxO7247nu9S5
oMTObAvP+HljGJ0EKR/fm3G03EtchVOQPmzLypTK+aXrNhaLHZUgzTrwFZwZR7UT
+Dm/jCM/usrsuHoqVshJgiq9uBMbgRqHgkU2NVOCsEFgV0FQlgshvZvsjx7X0DFb
Dalc7dlqaeaNLJR0KfB/37hwHUl+aYapppGHij0HryVOPxbPO3+EiwRY5uVbDRJA
gAVHrD86/+Z5gxm/AzenklJM4SH2jMDHSPaCa0ZyiKZYAycMFkoT8sZAnMwMbIn+
lnTxMndmuN25L7ukJAqZsPOc8wvYQ/oCRHdxopaAI6Z6b+QyEsVxkTd1hJrVJk6s
j6LY/ypqOuVfj6qtM6C91VrnfxViE5qMqAud+I+HfQpyEPu/9l1CbpuanfbExKjE
7dbzCqYvlenPKctajs1bjSUJT7q3bTKrw1BAGdE2Tkj3dsd9thYoG19Y2S4AQT5z
sO4EYJU2NsBLcsaH8Boi6/nXJGGCsw6l1dcyVrD72NvPZAxNqZm0cnLZRUJpQH44
DfErtuw1VvICFSP+zAiiDBfXzKtZCs0RCXG0IjU1YrZ5oE9InsLB/BqUwPmrrmNU
oe97DyP5lkXC3Po61Zh9C9aDnnaZUDD+RDS8ucRxTg7CmFApaNrk1newYd4g5+EW
5SIQWbYP4QtnRvBzoYRcyxBjS9IL+p8LpmmCCdVSivEttG8d0+/oYScwmugp3LNv
vEda9XWerV3vycHm/rluy0vt5rwP1yed+4D4jIUwfVGbIiBlSgTPS4edoyK6//f0
cOo8OvVYx5tz0XHXCkJ3PDKxB8BZlulSSKxpLW9jKFPjJaoJRCtMIP0Iixwbwnfi
5yBSg4kqLdUGTuS6CZB6yZEcFlU3nP36cVzuyFLLuvfmc4g9ivwuCEj/mM7oiwQ9
7dEI0e7vltxqTi5YNKiSWRWnfQTKJxzA8S+MVO73bGKrL4v0Qpd3uyF6AUsBE0gK
vXvU//xUOlsEMbOmTWpyUPuVkbuN/UTB1q3gKp2hRjK6WyJUOinGsYKOJPN6kxKO
1SQGVeiBriWY5ls6gb367ubld4lfBcrLkbKylqRRbcqZoSDLJTLOyrVNmIFOslpb
MWY5TCMeAhkUmQtM3cdSS1aQDszCufdS0KJsn2IXcvWymV0VbmBagOiCq7TIZvUc
uJnQPqQ3SeRZ7w81VHz+QqMjAqpitfomOzcSs/irL+XM49kVxB19TyDh6tIpQMFJ
tS6jyxtHv3Hf9zw8pPg3ewNtsZo7BRfn6jeTYzLWI2ueYzwR/NQ5cOJlge2dqlgu
EDAhC7+Ivzr2LR9AchWn6V3FnvlRA3blTwyRM30ul4EFPd/sjpeHwIjj3WC5os34
4PqPnrlTzyz/3jxuMxybcaYCOlgas43cm8KUADrfRLci1Erx7P04Z1xdBFLcgFx5
/QT2J4Z6ck18NV6SeVkditj6IELTW0fd+07rn/QzcIH3I0ryAOjCOxvhb3CJ/T0a
+Oz2as/RyF7DWQzOTmq05LzPdUF+RflLzdDq4y01HIORKQ10+uJJ6B4XRVNKRYAf
s3GqdBDWtKDHKl7GRa6bSKDB0TPRgojiYvzkkq9Q+DVAarFkpLtPtcXU1YG+VeH2
aTuyq8O9kJVoLIYK+hqOuNR8fv6YG7BP3MFx3uwIJjQQkWagsfKLW0j1btThgggC
bLSYmKuYt+ypcRx1vJtKPzYbmwiFI3kvegIp7NIavddCq+wcFWww5r6oyHiC44rF
l9lnSORAG3D09+v/3GL9YAd2mP1xCbkm1FOCKjHsqOMu0dbZUhXfMIPN2vD1HDgD
sNHXyd7LcOugxHgOHz4hU7v7sIZjeeKmHsbZsSOPqWkaoBUN9wZuw/4uS7ETfsog
XKwbhCkf1YbGbwxJVD+vvwf8zEVRLz1Bvuf9NVgacuCBGzM3UmhiAV5kk7nfzB19
/ruSm9l/I+5ylkPuQlw6HhzcILqlxJnNBYBEauPVMX7J3Cuib+O8LVLjTiyd/V1R
O6VU36RmZv9jBYoDNxEDlhJHhy67iC7Ep4aC9L6TXZ8nQ5NPMzmLmApTPJEjv9zO
iOfCoFY5nvwuCAKt16ACkU8p9RwBi+ddwslFe5VYO4cpfRSnLLBjwP0yEhSxZfon
HA27ksCaYTwV4ybphFPLHk6nfnZjJd1VSmnE+gBIx4v31u472kuZ+w2gYteTY7a5
LUp6IPlkULpAR5DGzhk2cL61w6YU8aw02aEsT2JH07+ONoKxfKcOpF58iUXJ448g
FcfSh8YND67UxVBC/Q/uaU6TdM2f0g6YnVFthp7QPnh4UsnTMGz4Kpjv/ck5uxFQ
o9kB29c+SpW2m9p0xgvfDrCkJS4FoCAZ8eCc32c0U//UUSc+F5dieuIc3Id4N4Ji
KWldLjKTvcQG4+wjzfiBupoFxey8pyTmKpgDSGFXyTBZJLrGLHEjQfGGJFvgG6+y
81wxyepE8iXNjYc92BrMBryxhP32DDVhmSF6xGGvtA/sqfD5bXgvNtLyZ/rf5Plz
UImZhfOfcSDuvTmM9WpHbF0cYxBZwTmFV5cCRy5gnknZ90fmopB7Lyqp0fWea9h4
lyXg/5XRH+S8hRlfJmcFqSG15YUW6arSVcwAj8PeW7ziUoFJOOIP54rFj66/7h0s
76gVFM/NDuw8YsUT8W7Nr//a5xNxwD1Tv9xmMlz6idSsW6zmJMjQzMLw5faGs0Ha
/EbTE0mn3SAj7kovxpVeKCK04z3eGQ80PzaZFb4cENDARYmnpfA/KTlKGdBoxquR
qtYg/fjddXwPbbt7/D2K/I5iW3ThOpus8L0i6F31FlK+w29zTeQySSnYST9qu/xP
oeI9WesbIGRiHrTHVpUOmyDpIWJrV/3DCHELfmmMYATM02SCE5utolrJhWUMHNfk
bAp2XFxHoC0RJ7jQBkFEJMunvrb0jJ9qebKpTJiXaNIhiZNSF/xS/6RtnPqkcDM6
YYuJjmQtSWVOvVWu9RFiTRESuLWq4orh0zUmYdRsI6+3eDSrUw83LfS+nKJeNu2T
Dq4G4Ljto8z6LiafSbq+odlYi7r4jkiifykd74MOvpckbUGfQBBW1/JgtRLtXyQb
sQSNzpV2XYBjiXu8l9WAKM68EiGk6x3YC2NomtZ15VpncjpO++39t6Vr/De47TZu
zT01WoZ0NUcLnwuq10DPmwrxZ9zPMwSItV+TUQNe+SZfVNHkzNJ+Mar8ZIZlkpYL
e7a3W2F5xpqiIRMc+0nQO7rSvUqSHSnRS3bDtzRpUTYuWyqislK0EIZDWua6HdY/
H4vY8G/qRuILUb5tJQYr3D6jf1kElNa/08U/Jo0It9kx65W95618ce7Ois2UvLlg
K8yiJaJa5CRzWC5TSEyUG31oYuH8cfC0QM6Xpu263vPc9SnBlil9wrgYl5L88zJf
AGqvnRIyV5l8xpskGqu+Dv3dVIoia3mS9SONNRiXoROcsSaPr6pAIw6hCf8tkk0p
0D1YzyHgSwvxUQ9BvYHvYsSbcHSjFC1BzsaR25TTETm0h0Aj/Oc8OIIBb7Eqm+IF
Qk0PP72gifO4o0DwGkFfGkiiwIrs9sDklJm3VkqPoYMkjMAPFT9IVvKKqWyBwJ1q
sm7/zMkgBnoFgobn+EIcPxjP66KMkKYehCzbiPUaPt3EDYcu/cRfXsbx30LHnwiL
uH1AtYViyLCBTjQ7UqLTjaLuDAo5Hd8jSODK0ydAyPM9oevGIA6fDFuhgfsSMtHh
sD/iUQIhf6/etgl9LyTxBdm6n1DXKMA21H/u+qmuCKxyCaIkggQHxPid0c+Hojjn
7OHJqZaJKWt9qoHnxziwOq8+pgl0wa//FerU5GWiRkhCSNPMcSXiVHXUg0b8DDIS
6rfyl3AbuHN7pzhn2zeLPRorn+AW79tpaAEbDgsTpnRluzJGKUpRsKw9rTfXlKnj
GRazUv+NOPJI4sTMFYIT+FQPwEak690nxS27j7LFGRBU94GBOivWw9PYSxfQUy+D
sNA9C71cBPgS76l5USEUsiwAhA2DYW7oTbphLafhhdw0Dtk8C3yLRRx5UHTrzFGl
rPPzWG//ASWDvWnnNnKxIi2AedgFvbG9KxnJ/5s/W8A9QcfQe7RnmWEpk1zZyAwS
0GA50vVtbmZ/g5+SuKCmKuczX6Vej4n8/nqkV+CCHl0tpU1WANiM9EyVT9FzugtZ
Ot/TO0KmwDGeZvQM5iOZo7B/HyEOBvRpJ6/yccWyXLfl9IOpX0Y/KqyfnDd+WiK3
Vtsp82/6rkW01ovqE1DzZQsNyt4b3jDFYgfz29h1fvASBAL6EH+SUTs/JGKDqx0x
t8p0Fdc1mDMVhcT4juTylUVsEH9dAKP/dwbnu4GONzG6OK1YTi/QrqBRowDV6gR1
9e5SsippxmYhg6G7ZN8Gu8yZ5UWDN+kglKJBhtrAGySVvOphcJhk+nWuUg4bnSfL
yX2M2f+ezhTw1xQV3OoQHM5Vl3CY75BvyH3JrBDeSVTFN2IW0sxyI0roq2BBYaUv
dG1zMRA9s4w6c3QP4CMczxKxC+2yaVloCJXhrC7LKYlM7yKzLJc7V6S0+UQWkEig
Akx5pNWsK1fQJBs8NEmcKns2zXdqtb/XElHjrGgo+tQPSJnj46WOYGGIU8BcPsoh
jHV0osfzQ9xAaHdCHklgX7/3KdRWA3pzum7pJqaQ7qAy06tftTMQADeAKDcYvXVc
fz7LH+J2ZRQrqNni6N0ID1JcbOOKpmfqD4yhUZbN4qc7aXdNoSgfRSzExPhrdG4f
58n4ov2lrSYntlhYYLcySGB0YKt5KWZQK8n64CC55rjIG089heWaVkkx6ViJTm8o
3L28KHaLa4wTgYesLE5Bp324N/MIpnTb2HINYpfoupL5lBLegPy9vVBHPnpMt6Al
JRIPQlYqBA4YkiNJX7Ijw9PxA/tPmBv7if7ErMRnXkP6RYjtdvum0c5bkvGITYqY
etgCk8OfEC2XiVpigIEWQyzWx09jyq8M6Nv1ETbUIc/OsRfJQOnI+S7CP+bvCq7W
GtgOzEq7cpE55Ci49TtMCgybGtzRpY0mdEyFdFI3QoQi2UTJh3IiB3hvWLfpJHDR
zc2rhZI+HfkakmufWen0G5zwtuWqpRztS2OwNiS2vaDWWcYqFJbk/7KmnRVizK7O
Osephblb7BqRLmbMX1TDBQUn6A1SjpBgDA7omT5mfsur3psb/IzNXGhf4n3n7vtL
iLGDU2kcDtZsHnS1PvvMWm2ZHHuS8v9G6SnpaAPsG0gMgsdJ6pJZi8fsMqBgCZDc
tIOhuWT4zXjsin3Zn8/tgbIfBovyWqnckTQVLUcXxUKxo/Ka8wKl9lvbOvma1Y/b
pDyuExNcnj56b/5R016dbY4q4QItaw3nyu5WJEj+s+ULNBCnUEWJ0yWOd+8D+tfb
R13zsEiBN8IF8h4ObgNAhHhyKBPmLlbgXakecmtYe3Y6IWKmXSCfCeN9rkcdA8Mw
9TlhGRe+0E+qdY1Uq1AmY+rsDgXTQsfBF4kkyY3IE5KxtU+1KHe45FP/EEZ4weaX
qej3WNp3zDeNpo4E/lK2MBWhJ9ezK1elMv3aXqnF1ME2camHNnbZMbxuNLBrxmO9
+arIRCXxDhVxZZlTjR8qtj3op6+OvNIRMldbkKYUTTouvIaAAZVOXTNuuyPHlNnW
MeelSFFIMamaw3NCcesIxIUOIffQCtpkuB4RA6L4AU1Ly30FS1XLV0hrI03cFe4O
kpAi46w068DOYnmfpb54KCT2u/RVBwklXHozNovlXQAsGwtZrZE2ORC/ZmO8XAP+
YQOb4LewVBrZDugseb868gKlkLrA9WbPsbp9L3dUqiVbRLFzQEB/FHLVsUbpiBVY
UhYpZK0gqVkuQ/6CbxAzTQd2tXCqFr7bf0sSBnln37Ehp+ugErSJk5ZXMqMJKrIc
yG5J6ChWJqUTcbYP4mN45SWkbgefvanmEzoo3p/uBSztF45vE163u2hDf+UrcqJ3
1AL4mXimglq/TsHpMv7kP4RufhDwHZ+HWn9/v2N4YcCN9fSwgkn7lxK3Ov1c2Hjg
CocryES4jkMjvWQANCOxRgz32r90qHfs+QRuEsL2PNKzqBVQXE12mAEgrQH4OMZp
hzNI8A9WeJS1KU+DWjyPaMAlT3zuF3dGcw9b2HBbSv4T61q/qpLlt9LUsRoM1umD
Gz3Whzqyhig96fkI8fBmmSH7TpALuaS/o66bqZ66usviL/ekx/6XZKgQdt8EPTyO
PjP2aPeROiWp3S8EEzvh6NFrFOFp7ZRRo/ipzh8WPbn0x08QaAvgTdlULbXkiuUu
vPLDI/xO1rKAvavwgLD9L8mEXndN2rhORPbcOPsVYFM3pSP2U2tE7PbICxOBmdL1
pfEqPNLT8pXnJclbbbj5JcNifULMxWOFw3HIEoL5ek4XRvnlRs8Md5BWejMNSPU/
ioT7hW59VnqjB1gPTyFpHn7iRoG0n1tFGAOXdG1QcsskYxTtSUGYWgX7Fd6N9E4c
583YgIhZVKPu0i7hp3Fe0TzNnF20arnt6iLBX5wP478K9LzIhpK1rg/qdRjHxPzz
36mqIon/KLVB5O6A3iKifXuXeuUxqw1PGQF8tgAg4KWMK2r5d1ABNEFiLyeky0Bt
Xk0fDw8CeUiKdDTwRDbEBjhzt4r+LnbRtt7Mi/Ls5B1ZpBo721S3gulihq9i5wGc
DphmG6SgxutxDN/NzdZe1rRBWy7p/JSSZx9WfBJ/EgMr56JBawIaI+FXcC+u0EJr
926jwMSr6wgac8uZyoVJF6bZfW9zVodjV3/O2ojnXD7i5AR+nCixoZk99Qqzl1C7
/ZafBmbWAgyQx6K0NnHzAFOgmmsKKviFxH9cmyYIZ5wiYsA6O5N+HW0Q+SWcJIqT
UxQtL1n+nXW8zV/OSOIsIMRcQ3/cXEBcHI29hgX90Bh11FzxlMDeroe6yyqlMKhU
Lzabk0pHuX7wfTlEJewB42Iqdz6RcTmwrI/n8m7ZNhxjqPAu2teWvTtCPK3UzaTI
o9x/9FQHv61J/ZUJpVp7curM2m9hh2VLfwLwS/BNjgAh3p6UTLT9xH/OP7Blb5A7
kgxcVkGfXPPmvqHmLV25lXiwwy9FMCVUaLrzw7/3SzHtktTmDw/am78EC3kOC9/M
Y2jtix5zuHCFot00CaIEoImDe9mpcAaq1GLdBTmUwcadcQmD7eTUzLZzfLtqmU35
nxmf5vnezxtoOK24mAwSMnTSPHPPcEhQyL7ca/aQPU5nRUW8PFjOPM9r2RxkhCGV
1F+/kDyg3Py7QFWLTjXi0/xHSG4pid9u89RRzoTPJVyx9X6J7z5XC0uz2nCd/OjG
o3Cvlci24zZYScw42h8aTjxd+YIWaCHduy9e96rUedwAARqOBVDpyjYd7BHai07M
IUnZVb27qQA4klT24ots9z1maC4rEV/dXHZZxnAQ6AnXPTC6fN5fA/mXQ8duj+gl
zvAIIJdHGJkGYUXKpeHzPVeXpL4Hrs0KiOfQWoz0pP8F057IkJuFAhi+GbaEAnAJ
ZCEsw7B9oeWPmh4F5U8g0C8GL9gMoEueY25tEiZJctRHG+xu+HabfeBVjGMSxHeQ
qYWvL8brPkKBvovLFcKN1nGyBT1S/K+kXkqFacG5VhsIR7xKvfa2Pp6Yj5A1lp9b
l8ObRjnjdPNmiG/zdXLTuPVRhtosDccZr0u1WwwwxMpRE0feBvaLuvnewj+emqIP
p6XT+YgDWQkokd1fp+R4UqzUjjg3+CpkFhP6w+lckOcNUrrqP/5KEdfUsbOTBgdA
91xDnBSeiERc/xU4ZfKKSb2Km/Szfz55ZDUu9jQ+byUoCoxijvvOovIw6uR+5B/E
aO5W84EiK6z6xtUJQs0RH9K7KoVVM6bT4Y+x5bY+BPT0EJzeO4+ZM3KtNPs967zs
rav0JHbuYcjKdDFzRXzSBKKcq8DM/Nyoo5i2uM0h3hSsxOr7bcVJlpf1gOac0H1v
EvM6vROHDAJuLwn5vuIID92hcpEegU+cQpyTcNcpMj9xdP/L0hv7RugjCFQEiUcF
Wt1jZ/HwH1NZXgtOnsytIOiz+991GnFp3EuRQmgtNsUJd4N6iXcfd/hZoP1e+X7j
xC0p1X5QI0vpfJdmFVb58Kel8pIxG9mYJOv1ZFPLWN//kq42fvHTpW+jZCKxxPs7
NUbFdcwCdWXxYTE85AwXVyWWSRuJJpWbB3iHKVJv8RF7sAbGo5FyE+tsq9kvnEtq
8gFVf5IfjadCFAJ/0lcmug64mcUQsmrDlUp2NLKIsLkaZffnbSAkKAlqICFTi39+
03lR69aJYOHwpjlq7wtWo/3RaBFKlLZlhPIhkVIrNLHVrGa0nRVvhSe6Pyf1M14K
cp+vWvON6M/o3BxSWP/tpZJxhJYx4oNmZ8woYD/J/Zhv8x1hmHG7kdbOnfkfIbqp
SHoqVU3sz3/ZRIi7i2mxD/YgeJiHUIBv2U6n4nh2u6jRM/qiK6khz+y7YzLM7zhL
kbg4vmOWaijsbglMYRCW5TyMADOhR9Eg2V8VBBvEgE1h6XBWdx+S1162QpBmvjjk
xuvLbIOkuFqsf1gTswiOVcRw4rE45D28enHD7m4kNOWFW5siQL4MVDX+1R991+xO
Y+DrdHYzyWY9RZJjfFk1NW410edmpFEWvyE0osNzO+rj093eEYe6SzShYDVD6PRz
8F7ny7hq7Q8CqzjPKS7/ofg+pkcQADEFHUXnxj2bObMy9fu4e/B7tc5QSPdzZ/Zr
v04DWd3DYDAt0kRUDwKUoWjKgaqGDMpOZ8+nlW0lUNVZ0kTWQddRnnVUIwoljRLx
58RfuGxVZN/MQ9gXgMmAx1sr81YOTtbuXL68l/aNaWln+pVUARRCUw4kU3HSkf2d
9UAgIsso/SQyYzhAktWxlbsZDD+omuCnM0AzItAhysn/7S/mHOzI7FlHnPxo5eGX
wTAsvm1FbmXnojzWTDLKVvRmLh8DfkkcYsNEZi3VQpEvRI9FkmPKmUAqB8dOlF3R
+Kqg4ubJj6HHHq9rAOMIi2FAwfCnyDD8BSWh6fD8Wopsz7ZCjtnJWu/GHnfaxE/G
fET5naNrJeoV3w870jqcbglDShVhPwSMIVphBqOBmXfwShj4OhH+dCwqfbdHbc9x
XF26iDb5n+aqB20bHpW1c/e915gUWcA+PiB3MF/kcXmYrzeBH+Nbegn5FXavhYS/
LsmCTwP68WMjx7aF/XagPlGvrSZNtHxhQsca+oybRKF59MKLDmxnbKqbF9FsOo86
0cHgp0J8I2CzG9FxH8Vc5+bTMwwaQQpiwIPUpXORLF70AZu/jx6a46nw3NRF3Ara
gnE1U61EdK+vkrkXsEQc7gR5UCEfbKGff5TGHUIU9GIodNoFh30Mwhl0EW8/7Qds
U2+pe7/GIAW2W20ll+kzwUbfOjsgf4ZcXOf6B2qeUJy1WgcU5Afc5fz6mD63FFY0
b5BcgcQA11+rvVtYtYAmAupOc87G5R4/v4ctIaSZfqWLnQw4ihC5zc3VdUQdZ5c8
4pumUtvZHnzTVfNCtySRaq6GfcymL/scJwScI/i6KnUoKP/ZomcOKXMN8VH/z2AG
ydwSa5N9EdF87kiSdq3L4sutk/HTff9C7IJusX+dyGbt1uxpRBZYxK8oW5xL6/1k
rF/RxSeYVIZJiH1UXPEU6PJqRO2DZd7BmCB88MbPoWfYLTknDG1mVm0yrK0RBf7+
8RdE7QHkh/vH9wEE8SK3vOzqICai+730OrA98PzH1BpgT+9UF7KptUrn1yIx8po2
SWaT1box5pokj1+r2JQCbguX+tZ3TdKEAFFC5PCItRID0WNtbDHI54rPuoS14TXy
pun//mDfmO6JIKpyljHaRZDB3mrHi90Hy0xtSt8Sj3w1f1BJ7Zkvb0uWM4Z7Qckx
S3X5Um8Knhlf81e0pXLBFAYEeeswS3O8rxp22xhciUJqQdV66jaF6M/Skx0+M0Va
QNjj+ES59zgZYdRyCHoJO1FwSEQo3BE4yvB6nKh3FVl7gYzDSvlL3HuP9TOvcWPy
aBphI/GGH37hacx/xW7iTlGtL/EvdDRhoFfUw+M1Hlf9cwQNgC1MuPFvyF0R0J8U
YLdcyAhBziJQtcT873GJe0Hg7nG9LnFraSdHUKOXfXzdKPMa//xq0nrB2Ch3qpFe
vAKjmAXEREsbkd5SAbi24W/YHu8S/tDjgHZbPAcMWQY2GqjjAueCWykHJspP7XCe
4ZQHn1rtJwZbC4I5ylrYqSQV20t/7mmkky/SVlwLhUFYN4Z4TVzzsiea9QpEa0GS
uYxRWWgJ/Royz7r4TgPvLo0Z2FOb5gfHN8/ez78f6dvprTALF8xtOS3lVFSOiNfo
3i4GwjVS5kflHy17yxki3CXCFVR94uqGInED5lLykHPjgVaZcwf0C2g9p8H7Q4t8
Q6PBiT36bM5VZLkxjHdIeTdeNe5xfAb5n1nkFjKgmC/eY+Zp7Tl6NVq+dnUnTR+L
iXRrPpmj35p+PElb5FODI3CMibJgZ4kjO7H2tlX8eSQ4sExsLQkHyBk1/+BTp2L2
gyp6kRLFlPBTUVgNZWhNFL5+4EW4sHajHYpUvdnn6rJ7eVbTYU15PHMT1/BqnvCX
3r96JwzR9CTBVAnVSfiW8fWPQxKV8i+WGW2VThJ0GFdOpIuESii0nVFUcIlFNk1O
u4+QqoUFLQq10WdJaSzfJqT+YZG7eqhO3093wEtBdJgNTqcOsgJN8WRY88qmZI/0
T3kXd7DtXHXAmAyq516zF/yR5rtxZycgeO8MEW7aqTi6F/0ghAnhyjhASOhuCUim
FpfsfBdwvZfDiDs8kIfSipseDRgZ+t3g6ETjjOCNWLai3r0QjksNBNDbrvW3sbxa
g9diM6guRF7JKAXhnMNybYIcv8m2oLZ5SVCPKpTLOAfXrYe1rnEhrXFi+Fn0Oxlq
nbsXVahKm8S49yYix7P+wOUpvA0EJAI2X2tMH/sDWTYzrJeMdCMxXY4+MS5uPKpr
FV2h2VbvMpesx9eh+D9NM1vhvskRdangzoP6FEmUQuOwMKiYOJRJlVdcV6zeqMeN
JQEV6x0RaTvBa3Ia+myLWSS3ZcEpAvxQUBI9nL24Ur4337BO7TVrmOR37XMu0UF2
Vlcbt3p19D9GuB18EJUEw5qpMMEJdPyyZmmkmPk7eSxBGLwToO+Ib9NJrdBqOjLG
LPacSvi1pssUZTJHaVFI7kmOo8fVBAj1aBRpolqW9hbQ4B9qYTdFuf1Fx1PAKB8h
VxAFlKobqKheFuHR1/CBFUMxc6dyfJBtuEbJ+XrV8KgNiSh0NROFfliiSpqp1+Ys
sT0yR+Sslm5AHYNvfLnAM60wUAnL3eRsMOOUuF/kZ2puFCdjt5EOyhQDjH1QfjYp
6psz5633F1TwDQCwPw/UCSweELqApBEsIuCfD2RIWfdxAGuh4YI6yh+wcEV+gR5I
KVGlgDQ7nUdxxk8CaBwu1RStn/12ULnWsXxGSYov2CPDJRJdTGlJRJOkmhUTOdNE
s5MBXwRpiF9FY5iMxDLbytvhmabAm+CQ2C60dqFhJEuy3xKWAKNDxrCKYV7Uh4JA
omuSL+jEd2DCrHPqPHZKjnu+oAj1AktQLhnwbDK/45yj4eyy/tjJ6PvL8sVcmViH
ZqBMm8Qci6EwZR2uPVKW6zixBJDmS70l8oZae1mjcGwmgV5cGg9lc2tpfWDetr07
ow6tbOZpkWVF0gvNbLqjGxhCjbT4XHdbi8Bu0TiaYYnardMCxSSUqMVf4mS3DGtK
b5BNUJDh56grRqOLmk/3CluxJKiiIEPqKl04FeLtkATvGzCFCfYnkFI0C2V/jUqZ
SeJdUEy4BfpgHlN1Kndc/SJE6jOdFXfVjhYxYld/vyQlYvTla+vzoT2mlQ4hoDTI
CLlW0QjWAOa48a1YTl7hNjaBuDTrhXGv74eJJq+M4zq41QXN1hyjEQwrS/BuKN55
2ZxSxQvZNZiDS5SIjvEP68aIpNRY204YFJngENL80m7409JcdLvC5D/XxcOaZqGJ
vv8rHN6WnOaO4kTMvZ/3BRa5ovmzXxmsO+MIacjxipU9dX3CWNX7Qyk3Nz5RwKNV
jGjIBdv7OL3TF673E37Ylkf5mzbiEHJyELlEia0us7gwn1D9uGL86SSz2/2GY9ei
o6ovYzwS1edBZaqw6o/xVx7h+WDpcEjv3F8AJzNn8eWI7imAxdzspSgvF0zI/Gju
8aHeK2oLTh3ImDUh8DIat3PoC1VWsvxAglowhfNy+bevZvutiEBY4z2F7BTCDM78
BI6aQJvbeZ9JZ/hTdQE0e/NB8AnHerPsyq8zLV+SV48SUHgS9HYmm6YC0vGMqJ22
vemNePZBGV9er/wKSdLmMqQoAaiRNAB0H5NkPAHAkSY1c/ixPo4AlBhyp0b2JZXY
3YQcC4zxbh7kOMg4PPsJ08WOw7oIhgIXueYdFWoBORCQ6e4B7BmtoWO6WCZxRlFc
TwWDqDh/rXo9zs56IW/kqspdZV8i9EsI2PDC5Xol5eRMfZesrRbEV1RI9cFefUZ0
KLooKdAfSJNnDQ66joKr2yjm8hfUidwIJxdcim5eh33hCShkEGiO5XZzVaKOb+DP
37a6Aulli1qnIQxHcNArSM+XnTG1V9GbknMnUk+NKZM4MPBlGZ628D7iQvqMuOhq
k5I/Hm/LhbAX74v8LducK/if40gBjHTFgkAAFUhREMZtC66v9GWVt28FD1/PwB71
A5ngAo5wQSB535QCuQsUPNb1tXz9bW/LYKQTYlldxwQX3ndqfgC6NXEUEireXavS
EIh2D2jNauTLHVDgcj/XXDaTGk8bWSatBsFnJoBAH1M/MAXPLW/qNf5XQ/ljYFRK
y3g+IlzrluH5UXOqX4249YltNWkp+RmxTAyRh/UlLbfcAgRSX+Yp3wUqRcT9ik6i
iKb4t8dy79KI7ustUmJUmrouqpHa1Y/ZHkpyBUv2tmYEdcm818xMaLn94H72W2iv
YM1fJRvc8psxNzVBpHu11ZpANohGxYUaIDxc7yvnlExdA40DXTfJ9r9bZQfT1Qwb
ari9Ql/oaG0NMJy0YUUiSXKi1adO32YgqirUgHHmrIbJHvabOGEuwjhoXvftoTKd
RFp1dsneeRP5/+hMGz36GWDUcM/QESCXZe6m8LLTImeNSYcxxEETLktMiWJzpBbO
CV0XjsjvU7R/6Yl1wB2l/hEIBy0Y3stwjzL9kDx8QTYl3IcrtoH3ZaBAn4qNKWOJ
hJgz0YsT2ICny5yePW3nqhRGlOudep+Z2ZJDAcw07cAV4zBZQQlZHnb10QMj/WRC
mUP5A+FmaCWoQQgHX0VSCAL+0Vhc0uVNTx7XQt1n14Cc98mi24DCquOnLuAWyLVv
aR08jZzSgk1RnhzCefmYR4yBANWq6ZKIsMvasMbmJ+YwlxxLTcW3UYmqpijMpork
prQau5zzn0Y9Gn8B38GXw8JcriD6ZigU/eN/a0MfYIvgT03CPlDLAkn5Owy5xfP7
31mi6b4rzwh5u/N2YTCkgIEElUrTeJnkqn+ZCM0pGePTk7VNgrJZuHGyT/1pDw0P
NIy03lJIrN07HEURHo5mDNH8hasqOCP9HxiEB71/fqpbw4NNDtpxtL1/ORURmn3w
wlJUVhvtJoGNSLyK0oUyOmkdP/YvSl1+Ucogw03lgzUT1GDT0u0NP7URhngWTbFo
MFp05Dk62BiUwXaDNuRnY3I+K4GbtwBq2oRWt68OPMcGDf5xJ0Ivudf4hbJbKvnI
59o1dye3FJy/20qiwOtZdla/HRlkoNoCQfIprOY4ieTbtj9baPi2gVLCyA/fBtlC
Hl8rO48KuOqwdv1hEjm1KnRJMcTrLHUCqv2vbZYujZOllq4bO9Lp/rTwnNUln5Zw
L1ozKmboydnYuCVtiEzG8TqBr36yKGprc6vLOBIdMl/aglMe3dCRjRIABCKgzTZ8
LlP7snbpJSI9nTOTi4+RiZvu95Jw3ZsD/dkwiotPoVm7TDN+Im8OCEhnYcFIE5pd
6/jMAjZkqqku7hVXhRvyx1THzQx1YZDBp7l7pGUb7m1qGyPkQZl/ZdXVRma1pXzg
j69LPkCuiAxa6gIeamy2AY8ezThqae+RwRc4DUgZ0/JhKz2+QxsmUXuq4OunmhEz
FYBv2JQS49DyZGdKqWXEXIj54WnnE81fdWyrZZNZ+mg1w7tJ5THnE/0JWo7pbAV/
rMDzmJuK9OOX90tkAWYL8EJ61ooLkTu+5qbTE5QcovrdBe7pz1vPwGwvAj536Fts
zU1FZJfZMeU84rbuOMcGQOjfCLQq8yjX9wgMh1WVHT2fW4gaCiWnxw3+n6x5TO92
bZj/iejLLTz/lXPg/ItLflpCopwmTzTpfT1L5H1C9cqTDqqMCekE9Ffk1lZxUEOC
HGAr345NjnWqWSreAMR8YPCye6hQx1iN+JsP+r9uEQ8oyD2DUddfz1Q7E+h9voQk
jM/lF+bW5PdHN8rwOtwQqse9ijiukmUbQDBxJkcw1bIn7ltSNo1dLnyMf8x+rA6G
YcUNSysITmXlhCobvJOmvF2T+0/wNwXlWUFvNOL4ryF7BzuqDy8TqYkhA7W4Q5wF
wjjC787Ktov/HXiZcK4Bb/u7WYCzDPpt4rQlo04qyyjGJiZYa1eFwLfbsHSt1v8p
o/baSRAwV1fBk6HXAGQPevID6uYSHVZFctoOZZ4IjdDv7XoTdOPrN3vMTnMHrtAM
I3G0DS4w5yWLDz380krVDsYwyuNSZyJt7bw4hjGKQTUzVcsvxO4dhK3gNcEyS8N6
2xbEX7Ef1UOmRMRZdSLc/qdhrVq7ZEKbFY2ijc5YsJ9k6dlc0+hlisU1kRczatxg
XgRevogOfd8FsOqj0p/AMpeP1WsxVHfpWM/EHcV6JVbYuzxaGRtAfPAmdbYypImp
9wC4bQ7A44AcxYT9YKDFJVjHbVEDjFHwUyz6+6HSpAmCAFU4uLQsUFlrtohRRS3t
+TNqku1GYTaXtlCmtUFyRa+e0cUCrqdyKQxK8XsStaeWJK3NVnKMCf8ggd5LIvU7
2q9/eijT4v2fWh+vrF16WKvAzdMNNmh4jgQTwyulwLofngQ5GI0rIx/QDmkI+qAd
jPk9BDN8ixXvhuqzChZ5l6Cc2lPpkI+TLkFmIIZoagk3JEOZj5utRNNQAbzDg4f/
0uHSB3DNKLXZ9IgIp4fCQxwS0ko+Xxq2rxYDfglHGj8ikfE3HaGZRM3+gZQanbX9
Iv+3+jTSnFwl+GH7QaBwJ+UnxcYg0SEIIKoa+NEGn9Cqm3rdu+CH9ydn0AEuQPVL
Z6tLUXBTy2BVraXOzyS9QxQrRXlBmFNeWCbJxv2EYaoPZbHnVG7wSqOQk+FkI+ne
I31rM4pS7utY6dUGDGJm3l2i4TcL0aeaoSBzXUbL6uBwZyUnKjfKQaflDjMqotWl
IkP+b+JYRnDvKx2yFK9npSlc8x2Bnqxo9d6J6alOFDNa1mqhMlFjzhP4iLyhRx1B
tkHdEwoDYY9xexkI4vrD6heTBuggnoYE4CSfsVV5wC0Gm6GrpLAHHsycy29QONNj
+BDJb41OI67R5EmlKme1lx+bovmySAj6BcKDtXzqVM2+m1GFNXhTGrTAKRiRrohv
l2NcLjATFivgyk0X00QKYHsIIUMrva0cga/MHsMftyzbNC+/z2LvKPrfoZRBqWFr
Xr+brcVV3Os4i73ffCUIP27bS2JePqOwikakHM0q51W5SO6f6vqpjMPGk3v3nQLh
tOLsZRvyT9eAgPM7P2NHKUm3SjMvYunshJziT+tb3Iwg8EtDJeOz2Hw2m+bpFPgM
/rnTXx/H3ok0pzDmKDlw/206JmaJq165s+sDn+vZYlgKCA2Q9v6ZSKtLDNf4TPry
Ppf4JnmwHiTGS+p+2b41hMVoKWJt2u7sQW9wvxkeS8YU36epZ2kutd9xZUiFDfar
5NOrvlPZsX/sVho3el1d0i7kv4rKXr96agNOMr7Avm3jj8i+WwntEXNGtuPqnsdE
1hcspunz9Zwqns39pMtKrTtSeoL5n0i6/zLldv0MGShersULGHgDZR28j3ZVVfSj
L1SAe0VMUXMd0vw2DUCgIplThj+yv9rluPnyXprCb4Xn3mWL1kQ7o1+CpK2HaBop
8ci9Lw9z9BI5T0fEzFIUqJT9fXx6zDWFtYgqqAPOjRohQU7U0s902gYgxxRIfkLV
x0Dm4/ruEFyAV3UuBtc7P/z4sa1FukHYawym4U2lOTFEgnBzERHYnhhJPNEWb9Gs
E9Xwgz7RM4NdBiuefIxYLvK2yJ8XPrJh80a0Ffzln41papkJjywwOpBaeHtIYID+
HzGdo/aO/mWNZTTS97ySzqAnnuuUFfIXMxIgVDKIkXiTGPqprtspRbYBQRvNSVjj
XPULUarwyMrtuHW9CoIiBYvc/KFNLxCoI7zTDTkKFfAInyKLfk+e3cUOmHLbozsp
fAJSUTClWbpDmBRJtPK2zywgPZb/cm5w+yevmPNiuEV3hZPF87LwXP+TXITGYaoR
D12UTcH06TCrqh+IkyAIj78oHD0Qd/rPm34q29F8513i6xJvl+lx6iZ7MqdFDWSh
IStSFRSWipIIa4j/r2rbC3zT2OauGfIh3XC3vahz3HVbwhC+2zpxW3jKC6La/r+F
Oh9pYl3wY+39xJlpaG/Ew8sbtWwIUnfLYH7JQEiJic2ISd+HJpP8zJKwPms1JMmh
TjmvD/GvQ8xX8YO7Gry3TslrDPV2SzjX2bG4MGbeqIp7QBJX+Nyk0b0GSQ5XGujl
m+Z8KmxPpVTr6O655QG9lMv0Jx9kEQbKoNVYxkE+KqUP84b8kMtbZ/bScbxNpEP8
p8C0iYC4qaW7wx4fhZ6of/hODbTBlNSaQ6AoTI8qC0lqNF53D8bhEJMakYSWVm0V
8PsGYAhjv9UBx3mD/uEtoTaQ+tbUuyMhgDHgxaggwOESpvzbXx3zPG1HoHq/wGAY
IKBMniO+7YvN4Nspadvf0QVP0ZiS1PU4Hf7onSaoIE4VGJ4V6ZWqrqjUkxYP707l
v+zAB/7Abg/QTSZNeCTDLYQK2KNJxj9ZlnOXKr3N4iTRneMla4Bt18sKYv3JoShm
E9cfIAsxfAHt6JaFxVPeydeMJ8UfBt4CzneMQWrle+KsbgZWPU48duswGWvs43s9
NPU/mqucCgaa6fdorEU9hydp+8VFVt/n7Th8NLfVJOPexAPGIKh+4rR3YrTmyYlV
mWYejHQtijRsOqSdNu4Lh5Ydp0DtWyZ2XEQsWK1Pv2ZmcVgUuUY+IhYpFgX2oDqf
wXXe0Sq+L27Y4YxjLoujq6dVWEZAvHHtMHCRrM/3CcEoYFjz7iiAGFsN0TjoxIen
zAe8lRtlbGx2oGJhkAks3gJo+YN8sN/PimyxJ6fw6OHdiVNi0Ct+Oe8moLn3xaeJ
v9kCnGTW7+GxwT4QstnX1I0nVtEOWhfRL7XswoQO5TQ0Huuw0XsDRyUzNpKzSsEP
ovRSY3AK5EmQtRT/hIr5L6Df+H0wrjDWxCWpH2nWUu0CwL4edpfmBgZTOfNbmMd7
wjiKgiNgJtXBIaM6vu0u7koHSN7o9cVMniwGotGNlCMmAV15QNuIg6IfCFr6V5wt
5/mREgdKKRpevU1pxGMAi6mqZo/z98RWSRe+x1d4MnInFkYBq2vYxw5hz+jjKnDd
bVRmvIZ5Eorh2gLu5F8kDeX56PltUxhBEMxXDd8mpcj3rdwIf+NGZ+tC+kE7tk7r
4zsak41AfrLYAr5K5vLrkfh591xG2Eil7k/joiQVkZz6n8L9s8p41VsjguoQvEiG
mw5QkRULF26CAchs/uzi1Es6QkR3aUNd1FKm8aWICyOhPgFXCGz6LlL2zSNpC8N3
bEbnLSIHPFiP8UUDV2w8glZSyo0kRge+bYMTi0/fX6sNqHudkdoyEyuLx4cU/Tyf
8CGFZoAUWsCO2J/arI193sgC7y2tk2jj5sHtik6v9jPCvG/PTOSBTaXpcpEmPbal
r3FFUiLHYLQkhn8mDYDXxMZf4UhKP26aADr43OfLEAmuhdt35Mq62H/Ix4A8RLbr
hn2LyOHUTeqi51C2aoPcG2cMl7IPSL/KbHxv/yJCq8W94BNZomh+VBcHtY8jmd+g
OFCYgxx0b9CVTMIpbV/fCdeyZ53us8BZm1/E9VSH1qPeBOCeRD/gacMB51jc4t95
PA892w+e731b/lV6/+lc15n/C/6DtbraghXoU4Mriq43WsCzNRfnFkVrx7OWTiM5
J7sAxGhgseDlqnKNFfaSSCQ/PvJIAkgYKGO492Bb5b7BD3WGxUCGdtDPB1qmMWxt
CJMCFv/ASQLxyMpJO6WIaIwSf73Qrc9mD6Y3/sTBb8poZXKuC/yikQn/fo2bIM2u
hQHv0Y5sJD0NcHVlW0AtYkTyPeOL0S81W1e3rzmjJmSwtkKNFnlodVV8Jc9P8gQ2
bp9tmy8/+W/9arPZ5i+V8Tn0c7Y5B9xDA8WLvmlC62bHyHhogI8kfpJKkyoRdow5
I9Pu0jhWpyGoad74cQS5FeY8pT/ZNbYhwV7hkY/XbBiht/oKiiP2DeeYmrwINzA3
Sqg+xwABUMuZLuTAydOyS6dCDOrFINH8FyjPgDsqRs3KCIukulmlfiG8D84zO2y8
68Rwj155AgE9INGuOKG8FCPol3/2StPd9Qy5Bdsyf31a6pyiCv9lba+tjPWWYd4k
fdOviNQo2rp1OA7d4nqM3Q6GoYQJRWK+cY04QwOSw9SGaol7uNhiI250PVgOY0pX
KJBiTWgmGrAzarsQ/O7xs0ZHjj44+i6TdjaoI3d4MrDaf5VqkoHlMINH1RGqsNjK
F5JUTGzLRRSp86h1vr8lE+sf5bgXLT8L1AEvBtlL5Qxft0wvJQs3dWBe5QGrG86v
AkA74sWzTjenVw4klPjKXrW4Ts960oVe2Dg9wwY6w8fKMr3Fgqn5ZLpSwKQAaDqC
UDejRLdUezEK7K7vIXr+UpIuSx2LfWH9B8lngyIrVB0tAd68HsbCbT5voBQojJIj
tXlTxBJ4Zf5epwI9/BytY8BA5AOxZ4YM6ISeOWOG90o6biDGEzylZmmKpJQvi2XG
jhVXiKFg74VnIe5sS+CPn05424E7du7OROEOHk3hJStGdfbUDfZrLavurmgY9f9g
QqQi6ijbGGU14a1gOk6kZnMI0hibIhgWv0ZO069V2xfjaimL9GuBHuUumtpKOj6Z
3bp/KKZbppsmCNDLhB+fHjkMP9fFEqq5bxGN4BoyjbB62hRk7/erI/PuIOcjeurq
F+ZH6SBKhRGD+AgMi76o7E2UFkKnmyLlxUaJAw/YjkiuFTgdn8BLWBwvs+cApbhO
EFFnjl7cKB6k1YZtlBWjL7gkypOIuJ59bTZlPfSDPSZp7lxr7AamqvsiubT4NLZn
u9NddYwkuOoeYR9VsGII4c7Itlb2cKhiZOc9kDMNnE1SYOYFg+lH0gQWSuS6wXjC
7M45phbr59nonLLtoVFTeUHqvJ8JBd4pOKDlzr5Pko6sjp8eDOs57VjSi7+VnIVf
O2Ostr2UlIMlffdWglc4TaMuf03GUWCRku7zhUwNE+GvTY0BfatYgWg/7/jxIc4B
tr7bggya1b1wYgdrsUQrulg1Dmqn+WeXW/PyvQRGqaBf6VQD22Eu9Tlg94uzj4Ay
mANM/K0h2NmQU16rkCA4+9oTWomr0GgEeGVJOmThqQgBQl0rZwrQCUe7wm4dN+Nm
OGP+XFOCasxUFozLYORm2ddMzl85vsEt2X+m/DfHvEgJgoJY1fGYgK5FELishpej
toHLrDMiXYWP21GDfsenkIcY0rKwzM67p5W37g6cnSQZnV7fWdL5Y6yMtG7sk7Wt
D1idGraq4Czghzj9d93tbaVmJQPYbpEZ+JyDv/1aZLh3t6Sb9nrT8w0yK9sBODKA
HztysFlasa8ChOT7K8EqCQ0/oJXCtwOUpyslvZXDRIVUxP0CfXL1b9Z17EMGZVJW
0RqmbhPJCrdIWBbtH6aJ8maumYkK8SzFXwEPs6v9uNvjVQ/MPZVWamm+tXqEEeP9
Uikm/Lh7z5fF9WF228106hECywQdY+uwjXHxFR9qpfrlNbKgm22B5lHsTe83jad9
uNt1BHJGse62uvMIt+8qNx2xPze83U0L9hDq6hTHeyR7bHb3HT19Od8chv+wZGYy
4qEONLPhtLwBQz4nhOGflcoP7Xd1WEI94DdHvn/EuVFoAna2Jl9VMQar2Xt5wD5n
t5pkLwf9Qsd3lV12YgCfwMW8TAurh4FQCG7TZVYdsIA+kpQue3KKxZfAbRpwr2e4
r7icg6W3hOwCagUPjwKch8MD9FO92KgeXz9vBaq43Lwpwi2wZWEIEmr+TIMnOyZF
Y+SzTbiICRYLB5L4Um1XXlhNPX8mFI3VFUp6aCJjdukOQ2C8Ec2x8xIZW9tNLvWS
edNNj9is747vzFBoqCNaV37S8GyyQTBgImdxmoQ4/Bmk/LL5HPuvkAiwNa/Qqolo
zKyUm2FrEos206+6dhhd0FqlobqNLDVb1vG3WNd8Gu/INaSbosRAQ6F/bsyYnFBi
fqb2MRb7ZYGnlcsxAC11kHhFoH6VMleWQqykbslV+nz8K+aFZwoYlqdxEoK5Y2lN
S2sCw5STPTTX1qwwAd1cPnMP5e5RJhzoF0t9Ar1/0KB+8m6iT4SbELJZ6WObJclj
eu0Cg+485C6GwJA3FJ1M+hoGdd8ZoaKpL97sv330zmpv3VLO/fnZwzi5XnHNQkeJ
7M3zxtO5/BJYxzCe8wxkwZyO6QUqq6DaO1sN8T5gOsiusESrwHCQyrmuwXOG8E2q
Vmb2ODnglzRRxlaY+359S8xQD7ZwlclF88ime5vYNk4/kLxNt2osMGsRSEc1c4+G
Ey+Hef7iw5ytNENzphjTOrzZzDyvQwDS2mXVJPWsfo/uosV5iaUoAahiMIpGfe69
YNZc0Hi+OSdWIbBzK1kv6J3H4wDfoaBVBAPW2+fPIRAknTkUEYpCanoZbZzmYosd
p6Frbrm8yp1I13tAwfMVj/1Mx8UAT9MTsAqff7pL1eLTmfAziySFYmJzLnErfOLP
s17fwRYlctJXUawseUDCrSC76y9hDPLza5aLl+WvQrpH5PB7kwDi5+4M2pmocV7N
ulDxHTLtu8E8sUdzwQdtnTVUhz9OOLqqtGxyg82PSsDGe7hky1y63KNHaaGjrUzO
HDQyPhEyA3/AboOyTQCuT1Wu9vWM7Jj+ITW1xFnbvhDkjYWbaHGsXOP+C0lVMMw/
WGtOXtYapw7XkcFTF7rcguWkzNec73LljQrKtrZo5+YuCwlw6kZTsZsf5EEB2zfC
d0gS/S24KHOLeEF2+4ZnItzks159hFdoQRGrGMRDRw1JsdxdaYVVoxlipp8K/fjd
6aeFd5v0PCJtMah03HRSdQEKRlQk4OUS0PL0PMoAXy78Kd2KUFzY+hGe4LlZvg4M
KMb/sqnfVM3oOytYVLeGzcG36WrAmCQcWJk47gsIM6qASreSK02mNB1G2v5RzKJE
taFSMBuNMqbaxAIYUDZWwhV76aPn3Faa9AnJnhW0wqYUOpryZEWBL6aCraOrdBIV
oFBC9m+hDvELaGGdp5kCyVnfOLp3xRQoal+JXaUD6KEM6a6NmijDm0a9gCJskK3P
GMV5n74EjJPxa0HdsulIjHsre7tAQEXDiC5L3mgRaxPQkuA9D+UH6f7bqn2NP1eP
Meb6en6/cKwr6MfKUiyiGQ4nap1kYrRjK002sYHcBtw0ifml2CijGXKWxbFoDQsP
lm6tlok46I0lysBS5W0Nj1yxtVgxs4XMR2ixl2blo+V0zDP1DIUjHXSLfvVn6Nj+
b9MZCDx6kEL8hv5YYUn8TkLWFBM0bY4sbpEjNbDPuDZuk0A2TaKrf2E/BjIhH/MP
ETICKqImP+l6o/7bF3km8MF9qh/TV9hvCRhFQc+sK9ppggECa8hrXEgMMMWS4Xec
qWUpSZIJBH1J1iHuTY8oLHPc3zuAFwTb+VYib3STZ+wc4wlcfF8RYW4NQbgxFmIL
zPu6NH6VBem+DdtdhyGIumFsG/xr0kB78Xh9F/KD0BPln8rsfcGRevhgVHSpodmQ
PrHIQYOIe6wKFSNtbHuVg+H6NNnUXtqJAdIX4APp7ANKOfoJtNryYCwxNeBxkFX/
ybR8VUFD2R6lMY3sx/4e3Y0jcywwgWpu0P4TNDobMhvqF4bqlDMmLBewPxy1UPGw
JJWLm5ZCRYAOz7aeKhUR0TC3MzIALJ7Ae1y0LWrY2OAsKo9cK53fcywekWcDbKlW
pygrKMG/jFbrWaW2WsQK8juVZ2e95rXa1dZynJEWIEiBqeX+5PMfbwFlMIHpMd/N
UYDydZ1hc8h8yvs2OnasZjx6YYf9l7DKJNxhUzkPQObwC5d8Q4jNz0LWp4O116R5
qI2/Rs+3+LXxJspRvx6H+P8HFhtjpSV7hVzRXnFOE8dc4v1m3SHtLNfkPoVwafQK
LvaLCrhfKjXzmCL8oXARjGaGF+wWWAfmPkrRbRTN3kxIwPVKGezeHgbrQUsVjNs1
WX5WXVrXVvahIvVEtq71nVHgq9bIRhLQDSE1l/hTqIqTeo8u4oroRGY5DopKd9zV
ewGF0eN//HgRv1syI5sgHZyMMG2dzmtWCpHHUUjOBYJphRU1EW+G1mkLzoIiwK9L
uPmNXFbYx+LCKN733o2ro1UVxNJIggmD+6dFOpWzIijMfKg1J1BPK6+Gec8nAwrE
y/7540A9XrkPkgHMY7QIwqHiNbQBRCJwhmu0+9wY7rsew5SHY5Hl10jfkkDRi74k
rZ0CcUgDOMm/ngWhX7yaXjIkpTzRNTfsYgXynKsGDwGLHY/y8P5gWPqOQircPZNb
8+b55Pd/vd5vtuC9CysepDF1x/CCjo3Bdg0a2Pqo1w0wPCLBkCfD5vDtTKxVfyk8
qJkm0ouiq45KbPzeaDGwI2h/JA+WnfobRIhv2TWSVvQEKwNEdVI2SymrkiLXqvUl
KVHL6lEO3Q9wKYSbQRRtUTrRbjolgK5QEfNc9IG0QaCsPltzRR/CY7XD9tusUETp
hxnx/BsSiY26pQyxdkBhLTwIeyHNyPpzzsdPu/ZWeYk8mzoDN1TQmUfcpFWdda/C
6hmadFN/pBy+dzui3FM/4vCdZZF+/Kr7na2tOxNXU4iqfRfuaFBl2kL8qcjw4axg
KyWktr8wOPSb5W9jfVw6rGcr6wot2/Zg0TxFbc7MFzzDHHjhqz071PvxPah6TGWy
UBeWXQkHM7yqU7/1/dllCDbBTukIy+mNgNRS0B6IsM04oc6UMPzdbJwSzTVDGGQa
5NtCQeQuplkjbLJAUrNSpBUE8DeWcr64D+870CS7XP2wR8FMWgBAfiYedf2cS+ZQ
TzsK8IXunrMXAZhi8LsqGzPoJYkpsY8CfSWzWsorpcsEKQAoM7ggt2BfhpE5rEuZ
yelwekM/9adGrCcmelnikKcX6U0xIB2f02WkYQ2g6J26PYHibJSesxKzkxU6A8OT
IFqzPnEGDWEdkod4nMQqMBKSIqnW9ywT6YfZsNRX3UNDhU9+lSjpXM6OZ9l5s/2J
EirXynBWX3d40u57tXYW/DfVbgmVlbyuqIIGL+bH+9KSd1f2fWSsSjPm0LOmkX55
FAMR7tbSToqyxbXv0MwvNqMOPUGwdREWShzZmtItd78zazGxis8av6l/ZkkrCc4N
Jf07t796ffhEQWe+yDVPf/rbcr6G04DvF77OXX18TEKws0I9E97y+hwH4zHA/zb1
MorrXhelGv4MagHdPLc0Ttr1NVWx0MYoq8Ow54bRF56L/ZRxsrQqBbIKU27N/UL0
zyrNjW5hLy09pPh/Upq/r9O2zZIi1yZ2l2mtKsMNWHI9qeBtORNCC4Y5xpN9V/Yh
4Jt4CSJALa/3WNpp6qyqSk8EiaxFkMYdSUE7pDgPv0MeY0YSJF6/3tan8bYqZPPZ
ZVlDXqY6EdRFO1WGknrNRXI4bTzDWRVWgmHj56YcpGDTkT8LSSVQokzDfcC2Z/6p
DYr6yEv0lfCPYd98aifwsV9H2rXJ8esV2vbYZyou6uWemWGw2gtbwkN/lrXukUuS
nRmKdY7KoGMB7mc2MiVlEJd/yMjxtNR0b5eymZhi3f5scKWDArjs7pnlZ+MTpvE/
hhtZptBzpycNL6d5pr4kxEbc41VyxQ3J877i3JusHGfT9HTzTQ/8P30+PsY5QBFK
qJyROPEBG0sSJXj+YDHZAV5LZ42TlKwFnq8HGVhaiwv3RcfmPyQB+oA2qrTf1bVY
zugEN4Fjv7vh/TRQkujLID1Ob0V9E3YS4GqVreaLAGiF1qoLeJ6Zfkp2sAU677Ju
pn/wJcCz+1RduQHmIA/WyFQOLSs4BqoEwuDFMFknyrVFG5sR5EYjT9kb7hSqLe1B
8WelA2fUR72iSWFagDyABHEJceeGMkR9XwoFwl6N4aCnJ1eSweE5k0iOgpIlUIoC
u937TP7LfJ55gYiZB+fEHqjFiJjfKTiuJym4YflegE5eIEoxFkh0i1OP6Lrw2+JU
FA94Iw2tbDRpWOPPxCi+qzzg8tChCEyvcMiCUaQ1pIKYCBesCBm1e0qVrVjvilwB
pBmePk9Tr5XblTHFCshw/+C5Y78RcCMBixeHiN1tGwNOumaU9z81wrVbxqILFEtf
YJYYMzTF68O4bV4wVO6ZoqU0BJsoSl2dTzmFNUCCHBgqL/FmpSExfgdRVDukBlk3
HUscxsq/0OeeMFlJOIzNV/4LY83xIiu8V74LI8P/J8rKTnNo7kGKmigujuy40LkD
LfRZWqFlkOBSZK5iNO0TE4peUYy6u8A41WFnf94isjQtrEHjQAc/jEm2IoLREN6q
cTGTilRf3adryaDYL7LM7rG0CUQMMvetI9IxHBzsQHKvd2NYh0W5WWNNmTZGmj6W
9AN2bv2qDCbfEQWGIhdKxok6+L1+VeL2vfIhX3xFrEZ9v/bRcJhgQaPNVuequF3s
xRmdUs5RPlZ7mYkvuEwtTOBLgftPIAEVkfUZ2TMoc1lJ/y2UZnfHXFVzwq0t2AI1
FuqWCLr0xa18OMZ8ew0kjPpJGGks8ZxrsS0Czm+ibnUNst/s2tj2+34wUL+DxpMh
HEa1zIyZlR+Xrc6PMunJCCO3wN9W6pDzwmykkWHkzZ/R/Nia3KwMA+TmLcwdDSVu
2aQEbzar+q9Ui2xg1fbVLhyn7ckdMTAPVo11lLnOtPGzv6xtH+gnYKoTuY8zbb0h
z7MTf+KFjvOcLMY7LQmAdiBYOi6lqNSnGYu0qZ4voiYBmdZkWObRtMULABSn9nZT
CtjfVkJBTvsrNqb83Jvgflx6GKQd3QiYo5wjWLXwnWywn8iV3ap818VBrR2WXpbk
8dy3q+QirRL9nn9GIv7jC/blUkg4MG1J2HkB/qYvj7YC004O5jpa47U9z8KcXrpa
G+orxw0UnZWxpuYCKABiwCFX4DpvzAGQOGhq95y76Z25TbOZmF0Lyq/iLCm5PdfK
78uX6thpmBjK2/Lv61dyJGzGoYoNVvKQk4l9m8foAv3enncMxrYL+9bw2bor1hOp
m8qCu6yueUyRZxFwhRYVe0hMR/atllVAQdolzYxseKf8cVXpUUVmpjXb9aNCOcmg
wLhXZhm30g9UxIt6GrMGVbSZA460d3OIfvyy7ReNScL+J8Nj1pKCWfQR1fuaTJbr
EPlZHuW6b0txjiY3McN+STSKsU3w2C2Oxqs1prLw48PBWiDQyJ0IiRxtMd3z9Nm5
E4ajcGrSS9sJERo4S7Tx+ZY6RaI8G9dFA5uBHt66MvP+pQIuQ3i3ZLJ37I7FGI8K
cGIBBM4i/FOtgNj7mt2OIeM5MqGf/MW3gsG1cGuY3Z+nAcxK1kX5u5GXL2ybDhtt
e/2xfOl8ts6WZSkmhZEp9Kgx9Urt0M997vUS9BThSBX1fDVctdHQfzgCWYr+b16s
IducAm/W+JVrc/JXBt9Mjj2LTJIluNzMmNVh3mAcSdR3eFjr0qeFWGXspIKh6Rja
MJ+Tq+z1uWwEhjNb1loo16GPM9a3639CpfPIjMfKseYo9AidXXYsZp7UhK45+kPq
3X9uIVTf549B+7xYRkATp63U4zLYpzqazoGskshuqbRZVE8a6G0yWkIrSDVZmyzL
9FiqmvWFX2pSRSdqPj6y4W+5T9evHsO1kXDz494WGvPYg2JfupozGZL5Mzjw77XC
NH/YK0rrmslU1DHuCyQSLs1DNM8mLessTsi7ukkXI6j/XP5tqzJ8QJ2aLPH9sT1n
iVUrVreivq6Pu0/VBcI4vBCe+gSciBgS7Ve5qJZR921qeAr/G0NV6JHHXwBfIwn3
HtGukuWWv5OT9PPiJGH432agPjEzSWqKNr+Zl7lSIrrXYM0Ky1SWGjItPrHe2jzz
HGpScna+jUpx/rHWHlApg7NOP8WPRebjFsckRR6WERMd5RdOYYITpsZBAjry9fsl
IL2OCf3vsN4GNvcggxV+GF7S2pQc5JosNc/rrNo4e9+bIBkagfdG3mFnTvcWiMdz
Z9ZLUgQosHCi07jE6GAKNAOBvI65lXJ5QfCeT/ypt+1D9rWH4EpECWLZGYIyL/CY
q+0JaCSXUMriTlTOEs7skBnIGaF9B9lBb61v/XVnaHlaZeK1igbdkJB/46MKVtli
Hp3Z23nZRy6O7MDQZWZd1KqerIRlg7IHfR8poU3sHagYI/jk5+kYh5afQNPOMA8q
ZA3t8+7+xJ12bXHPS3behLxc44PDNEfey/+663EydT1N6pTqcamYTX98qkKkhHFE
dk6vdH0zNs28qKrWNgytzKVbvGUrarlsUwjWYYKudiEWkspdZZ9Slo7gpmFqXM+K
6QSV6kxOtG4l451Il1Zam5prhl+g6a66kdLIG7jrLmFZnPuNCce/DDtUuJWARccw
aLezC2eFVam2IQi1ILEMpzzPHekKIPIggVzgSuxsqTLVF7wzX1qRLBMrQvS6P7jL
Fov+nnVjLJXaXzd5jThkLNz1hOQlrvkX0v8OJMsd8J6N/w2ra/b6blLJ6aBsfCt7
eaLN1zM4KUU6i91yQuSYTMsG+QJrfcXTJsg2mDQkrqAgYihQvVWyC4ciiBbRCVmR
pj7IJvN63erDoS926AU1Osq0H0u7PCKRPGQpYrwGZQ1qqQM/YIHteQeFgISrSJgC
kMN1bULLKhHwlyKoWwvbWlpesrg+yJYDKU+tcQTweUCzyJLcWfem65Ic+Yy2CR3v
gXT4ECtxM24LewKkzpYixCdLC5JZtiEJCXr84UYh7kIKyCyEQDy0YwJw/yuEt1mV
J8XSkv7/ag6Q9J65ZIAZeMRGzeuhsSPPtn8Etuxv5+4qszSdoUSnCnwrT9SjgzMR
qw9HKlQNJCPR2RIYxI98TgggZi2BPIguOnaciSr3XIMqEK2JrxxGOud++RPYLVoV
QHDH5yprxGbhZ2oc4pZl0FIKO8jms1fwhLRvonBl95/bPw2FHeEvPySPu+izNJMI
GXiUGQ+L7d+c7UQIWHCTr89uQu0wT1BINNHTDwZ/1JITC9JXwaRI7qDDr4v/e9EK
aYuI9VhRwk/Zk7zy/tUOh6Gsv7Ad74Og+bXAvkreu4YztCET7/35CsNIFhNDT0ts
X63n3LHijPVQ33YoJuVMT8+1Kv3B4ORTM+gHGRySwTriz+uHvGGlORPGgyysttlE
1IfGNHpCLOyVag40T7sm5HI3yd+exoEJaJ0obrEBom7RRIUoDMMJLavYLCiQ0AQJ
HXOW77Rnwyz7xW+RpfflwtVwd82m+d3ZqeqyNiXSqNU4lqO5/Usm6kf4JCrLPLUD
CXkE7AJ9BMpTrACF6vE3RMBBNTuRlquXlHhCxdPYJhQ1k+Vb93xdyyv9RbBrgjOe
zwxZlifCezQmgRZQ3tlBYuIvj5g03JoDO9qa3MhL37TChoI6eN3ya+Ty4Zf7ehq7
F4rQ4WhS6sNl5NC7xLLOKFlZD96Horm9OAVmrin0y8jvnKSSa5Dp1BzOGuEYdOFL
uyyh2dNFpfyIYLqD/fl6BuwxRUF3R/FMCeLxHAdrXGhE7BRfopxnquFn2zr/ElzD
T6cJUuFG/EL+iusfLxj5wkOvyO6Jf5mUv7gkj7AplTg4f9ovTwRg8A7sTlSVXc25
GUNB+zsBOVlidYB3cUgTksjJGpd7Ws2iEiLHjqn5KnM5wtfvZD/kw1pvdjHDtwva
WyIPkbbLptkXnkDDjacMJA3MSRPUhRGvlyjl8iB2t+4AH6y32mOA5K67ZfzFEE3C
Lcrlniuu+zwZBMUcYL/+xEugaMbUvwNNunhRjQU/AK+hAK9M7Q3iJYYJaAYGEvVC
wy7UkKkp2zc6YS2aVci7APMfdXdnHT1YARllPjFQwOzJmxqnuytNCDKn478YMmZ2
c3GUZZGTvYErQ9dBaaDUoXCU31tkkckHXqkf/q687qK9Zf7UsieRdKglRExfIK4x
U8RGD6e49s6b2h3kUdNz6Pb95vtlBox2GusRDk7FrfFlhl0EsgfIlPZY7xTz02Qz
sznSRCL+FX9L7/h3KHHOofTsR8K/JUKtI79bS2xRfv+J1AvfLH7VPq7A+ZZhGxO+
gtKqockhFMO7Qt75zMaUNXDvsQwMUVQ++mJ46kvOfjPIrbx1Vrmd6f3ZhswwJyFD
LlEJtm8FtqHODqQlBwUbsOMAE8ATJNdUHF45uW7eIqR7ftPN/37FuEgzj/Umm8F3
Z0Ksdj1anAzNLh/6zPv5gtyc7Fi/ghoSkjF4KHmoWjHufQyrWzt9aPerqUb5hg7J
jsj5zixWqNqAb9iGl/Z11TNtemlr9DOZSfRXsRkdBhia9YcepA32FKMHTannJJYQ
aRpNvTrrz7a27/ZHUL9K1HcY6q5DkW5ZWHHeCUaaE78lEDc00NXIpRIeLq9GrTuU
pZXj+Lq8VoQt1h15ZGutRkQyOA64z/59RmASqw0Mf04flAv7ExG4hD6dIv8NTKQi
8HhbF7ZpZota2YM2JQzgG1TZwtgBLxxjcJHdq6Z3wQwQFGVHbjjON7g2o7ijrp/q
DkJwVdTHY7tDXvWTOyXjYP/WdbtvitMpcfbg9bCeVY9qBGrdgo9/Z8PIR22+AIsh
/srugiPsvg7CVZtS2KaV1+rwvWZxWImkM1Vb+CVZPKxMWF5GKA6n2hPDnS+RSk5x
/YoGrHTHVCcgkWXhr8HCHewpp2ZNb8rONIsvicjLQ29pBwoFvS2OB/E3m3leu8SV
5air4JgXkcEqL8j+7EAJJB7JoKtRhs1blM7tJA2FPOyCNBpopTVcr0xuxsoXqyyH
2InK2OPN3togoH1SN9WSw/2s/KZwF/5qItapoS0gLYRt0W25mtqxuaw7vf9GjFko
7kzqXQKYbWRRVdm44oJJpIz9+HJSTngurvyRpWUUY5Zvu1QDxn5AuZ6Cdz+LFKx+
DASx1e0sixWcc13cwoEJFlueBdnK93NK5reU+KwqCKY1Ezheka+kSiVXRUxTFcT1
AVnwy8TSOYAN9WxSCpJFANgDC7qa5Ui6VVyJEe2+fr+1CUF0v+k3va+s+9AexCIg
3quN3Ij3gsi2D0iaAvFCgDGi208/RtZGPbWAlPgrTQcdezOj2o3BnL0ZM4kD3idx
pq3pcmU+EzDytaovvvLSZe1UtOo/e+6A5FaXPQ5nArDobeGP1l1fukcrTJJxqeOS
udpFWt1iObhyAbnvS+mYddFGqLCiIDr/7gYnsTfy17ag+0Bm33A+LgDwkaSoZcWa
tdSfDEIP4oCVhnrzu7u/xU8AA8wLzOFB5o22P9qyQVvlEGTARSKTaPY1S3ZKTeJj
4WeI2axaNj1znCUhy5kOktsGiGsJIYzCcftj4YCqW0KRURUPmRSvQ81dSb6XEw/g
BDaUQiD2Wo4NebPCqO+NDhR4GtaAaVNNg+36kQz5xhC6KtyjJ4mm1FSxs+5JOh1y
d1M91CGzRZt0wahDjfzJrNFifKnp7dk0iw1HLD3wq+W/O40Xg3ywdSgeS+9ox0MV
f8saw5CPI1NbrV4Q9gBWlw1UJM8LlG2yo0LTg8GKXA1rsZ5VGqovWTnhJgDTX7BD
sO6RMC3K54Gp0owpoO5j+cUdudL3fZXLyNyHaVHnjQZo5dqz6U3OCUb5sVUjE+qn
755foHDBb2zI2Xg5ZKOEv40DDkuRWG3UvNtEBUXKBRiCEevkV5l+9nm2zZCSKDID
AUF00UStX6Pysr4CaQhwMRENQN9MPFUPDtSnxfDwFHRghdKZoTlO6av9rt2xt0Hl
fcSC0EhMxqIbjqgbJ8UE2gD3l332jYGRucA2Pivt4gBLoHWF/7DLvFMYdsY8JP+z
1+hGkOr+mao6Ctmn9NmQKT5x2I89JBXMOOd2/LQYBAh/7HhEQsHhNGG1dIcer/lQ
nnLVtLvZkw/6C7uvXKTiEnwlpoF3yzvGDx0hJRq8MTt/DknesrxPZ6edSQZ8KkOA
qc465cCTUJjl14LfF6gWwhIdh34H5gWlT8lqAGr2B7wHnmOb3eYmre5mirmA/kFr
HNpNTzuMGsLiEUsT4kq1EKdDazk9ZCFCfx6dKij0y90bR+LTxHBVRpOl2qd4KETC
g2BPgSMFgav2lHvVRXtqbWlM0q9EkrvcC2LHoFVyNDDSLnBpSBssr40tW3i0vWPj
/Dic7UVApAJTIDH7aP71jP/sZ/76SdPdfPjREjsV6os7/1W/B/Nqqf1hIHF7C82x
+XtVGp9J1tSq+Rqnpi6Wpu2/oewfQ8Konw0QHWe16ojycq4I8FCvBgQI1Zxw2pky
irtAcSTSYXGbSa0jN4DK2J9ayybL6jihdIzrQ3lm58/fCUSJEU1yUBsRB72Yv5ym
bVDiYFet0IYP0NsWAqDVZGRFionVJE9QXAy23vjOFulR07WUUIoxBR7lm/E5yui0
JaIpcQ14aQH8Ov4dL+e6gWRPU+EmJUr6ngW9oK22FzKuiUq71oYcED5YJmKfZ3ox
lNH/rwMrPqxlRucCRQB2gvRLdYk2yaR2LkgyKvDqHeFY/cFvtCEH7LItLmIakhAy
sHV8PYUA+NTdBmstElPMkSKGS92Oe2kGaQwj2Y7hGI5F2RAHjrQFzPsGVXyeWF0C
K8kA5kIZ70ptMEurgK61XL6/ztQW1LHZ9fG7bRF7ksr77h8gvOkFyFugbBgkR0Xv
Sy1IGfGKCRg8qwizHLCTcTn1HipIBI5TQtfrXzTLtrIp+jfEdFjNjxqw3+/MkLEG
DMDO5W0cy4XTCuGc+yujs12tt86ns57n6ZtMpTjEocgQThuqO3JAyQU2cveFu5jX
/vl8gXaYFqGJsEclFxm3SNwD5SFgYJuIsdDac9XqTG0njFO2PQ8iTTmesEiMrZtV
0bCLa2seWjGzTjTJNpXQAn0KKP5S99WaGlvRQcCrbLvNFDeMlHR1AhrsCYr0+LTE
htvfxzWsDYB4WufzkmjLcr0dY/2JalIvUiFitprcOoWRNKOMSlfMUsiT4s4MVw6V
p6gw76MJ0iyy4AxpTZFz1z7/NAmX3RkLhfR/q4Hudek2poLjWXFNFmg8HygH6HZx
McEpOhDy+7ihqRluzvJ1SzuPKun4FvtYZQMsJerm1lgoE0rFMTQL7DZysGSUX3ZP
Jghpl1+9i66AWFqW+jGphM7L4dhXToz41J2AG663Ivqs/vqMqAjL56VWXZzw6AlS
Htg6v5stMl7u/mKMiwjvOhbvLzVFszVMR+3iFKynZyLDaMur/J563vslQ/Feq+gV
j6aY9xtbjTzW9b27SsfWSVPCjULTUFkpDslXHf7jk1s+SiSyJCu1FULfI8Yn8Wj3
1gFTq7Xc+B7wdT1j/i9MNdUrzqOh4OcgRjteph2DSzWrptLxIeC7Z7UqjTohGrYk
ZJeB/cPA6RqJ0iOPJiCgfdJdG93PUNsM1T9su4rY+B7dcA5+BPwwWo5W93qTwBrc
pkj7ikqH9BjQ9+oboGfAUhMT3Z54GtlKwKCqnf7DwW933d/0rEAEVYSzP75UkzuN
HOVme6k2pcF4Q94p+UK9/vpbDWhhFRFaeCekD+oWbuEY4l/0MX6pQzeWnEB4i0Kc
Dew+wYIbNPzv0ClaHt+bz3dcrJdE5i/ShYbJ8H1NC8OjrHMpnuCsJgUeFOOtj3/u
R5Nof/VMw1rH5nDWRhboDhV86dpQo78uZFckF2xHe5dJwHRtPmiXlUWfU22Gvjq9
L/ZkEgygDegIGTw7KJw+oIYd8QAS2db8hBSfnbU9cCFhuDtvLsQCXBPECu/zyn85
ex6GY9h+v5eHM+7BKlU63irmowo69v9lPI4MpQqp7MpjYDN9XnfpPmgNVQQOCJX4
6Psu2Kdtd0vlLXuwBfgHbPp+Xsf+iRnZ/mx80TTiq18CYjzzn4clOZm4t38U099H
BBSk4NBPnrohbMlj4+sWPjqjIzgX9VpPYDQE1dLv83bopTun8CyRx1MgLxuB0HgI
74/QZTI3Zbztk8zoSDuEgWYAAYTpOzm88tLaWTHVpgHLmIwicRUsQRIURpE9RmTy
l8d0rG+61UmgW5zeUVAxSvIIV0UGyw5Ywp7jhsvLjEBGMIqTX3aK7SXLkuazHiFF
XWrS3S/hOsp+qQHGEjt0JVr34XcZN6evvz8Y7RlojJgxHGUCAQSbGkfHWnwOCqxw
yzTe7u7m9uL/SKcUmkeM6hjbfjdqxGidCmO977TwQUZCxPuK4cwKkDccJUkOokS1
MMZs4iu9qifmBXEUYfU8qtzr1dgoV2LL/6A5evKC2VCo48PASrTuSIgQDnnj1olL
xHDyLhsm0e9Ej+QTSd17ynkggT6Ub6HYRIQBSFFgnK+uUB8ZnNw55/m/tz0ye43n
++tR77gzZoCUC1DsPum3OxefmfkUrbTdV0QY7T/n9nVwcqDC4yXt9AZ3NsdAo8+5
v1T9DYwB0kKIzvqt/h/VHSUoBpRiFf9gMWvL1oJ+ep8oE42PlhK89pWTfZFoXSaX
LdBzC8Q/c2IO33qDEPb9zIYzWT2OQaos9PcVcRoLN4le1inUutBWql7xfPQq3tTI
+u3NX7BARC8w3uvwB5L3YC7NAyXgRJC25aeV/BS7NSYPbfF41oRPRpRisja0NS4T
XQcHi9VRjhdSw1eV/q8pEmD7L4r4/mwtBgO3mSYpRGexjjIrQImpxM2CWvVxtJNj
IqlQSFiCRRez229BO0gULyH4O4yn/J0qNyYorhi2Iv/2bkgFHhrUnEVjhAGXsceg
5r14Z3wikzlEA5YZUyEuSp9Zt067oJzPklrBTOQU4u6bGESKJI6ubZ9YDdPY9aE7
GOuSjIeDkEkzcbHQACUAqKzf8mUFlno74EaHgM64l1sp/kmW4rBShB3XukhRx1Ui
Isam9WP/oLL0G29HvRnoIlrgYACT37ymY0hblx5Ze3g+r8CNAeJu47fOb9fR6vbA
QwIGNVfDP+hn/JpPT2au8C60Jdj6Cp4XbS8DMOpNRWRcXqOZ3v3GkWlHo6+Q9z5e
jQkJsrcOvHEeBQG0zdhPNrjhwcMvM18Exf9jsR3zYGe5KaA7axCwGetjXbGulW+k
ykMtnei1Vjl3+zAOBZttTs5E5LuvvNxGwd8Jxfl0OjDMOhOj8Ck8TpZ8c1ejLsPo
nQEBNKr98OZ4hczThPzxfIhvcD2FtFOIQrckt3tngtNQ9UeCnOcGpqhMReXEX0fT
e+ZpSMY6JKHibEo9iY4445Gi9AeuSE0ZTT4ol9Y0b7M9Hr1eeIy1EvXLxs7OC7TF
mha4ANN/UbUDEpl9np7ZJT/+olck/2ALrH+a7/zVwI674eFP0Ay7Xzhx9smjiEWc
5rHfgYnmO9eZbTH8iT7xFUdIrzEVyci0pYSNdzzApur+Mn68he6lZoCUEPB7vh1h
lNZP1QnnY6q96uIdkPTH7r24ssTSmPQeizdWNZsLHAgeUfxn82ZTmLWc49cIUXCF
Nx2ZUuZZ18qT4bW0NZAHROwToItpH6IVE3ftfpEYqrYDb/muMOUE/a+CdlVmrzaK
2gPwuYSmvE7thoOQwLSz0arloqYf+KfKImfYkgR6HhBRK5rdUEITn5rWgb2u2kDB
SZ4u+mhyNpQGpEGypfozuhurNNfRQUnN4RUHlN94N4nQKdG2w5OKZY6lMiKTAqJA
ndqlmE8qj46zgTVE0Fd/nlwat6uC0Ll5TF3ezDSwWD52gxzGmgPHGfiIDmwAdm36
WAS9BlzPl8f0TsDF4vOdpD5kSLLdSkLlpq2MGFnj9iWzcgfn8QE+LBbpaKwAPmDp
MV7Lb4IdtbimgmnCT6uITczitFIIXrV24qPVeR/iWYqAZRHQNwbtgrGhfdhoKKba
5SoNvbh0ZPIlTju/uYOOfT65x4PhNtTx+m/1P4oBIH1qjdA3UDA90HED1AfJmxwT
wyZ474rMmYoVtzx+JIaqQn072Rg9lh7OZC9WyGVLO5NIo1ElaDX7OGF6I5vKwgv6
txAHFIGNLK5F3BNRuQKPcjgTHHJa8ywWwUTCu0yDlLneKpM/kgQ/7T1PtA3VVUh6
e58IJPtfC2iS/LQfyt5q/Q24LSLsr0fkURFVOTxm6DtCtTWN4pA3BdOq3llQLtDO
uuAkzWp/eUKL68eQVzo4p/t0BmrjWgBXpdwqxd18CQBIyeDH7wqwzYPo6zRYMYgA
/XtBS5BAqbRDtfg2+5ZJyULCHVTqjvfC7IUVyniGyUUfnH1YTz4ELaumDW51Cbhq
7C9ToHkTA8mBnrOzml+KbwEeBK4/uFas7Ks54VUl3+486v8f+TzwsGftpC5N91IZ
yLui7pre+593nNeaMuNy088pqITxNrk6KmPanJeVOwg80NEnuhw5DzJkCQnk50tQ
oumKUn3RI2QPvtmOhGR81X9uo2o7dY+c0ftwz0wQczcMA0w8F4SVP9SOjuyF4iEG
ihwKdCCJwOncFL/Td1htrkg1lsn04EyCcggGHclYwoLE4N8Srer7wsJHuhvjfQaw
X8UZEqlvhG3XMyzRVF5SnMdx5xJrSrRguGCshEAG3lhlA+o8kehjWQZlNDEA1t/2
SofwtOHa/LKVHjdPD3+4PT+Xctveu1mI+Fjk2It81Sq+/4Q2scbp8O270Ic/9C5z
Rw6LVPRS3iGxPZ44JcUXXe2pYjAvPIh5m0Odo/uXpGHAYiTTF438wx+WYERmOIO/
job76FMNj0EvmCbn8KeET4VFe1b86a3AgH3zq7r6pmYriAUTPhF6TQxOusaGpFc2
W2z9HAwkQdIoIKvbtiNsQFMGEz0PKiD5QbAhq8NTKrSB+6GVoEXFUY8eHkBpPYiP
eQQwSN4WEdXY3VQoke75mTJHS2npL1V2I6Kbmpe3UA36dj+8sFo18btWB5p8lqtQ
7YtfpGD6ZfO0TAYAA71BRP0T3/bejLqVPkOp5GrNHicLTHY/bVacQvjOOrroMe+Z
/pNbJgjAYhticnY8r3mRGsrFncC7AiCuRzbyJxoQHQ6PLoF3kk/qtR4+8peO0Xse
ZZc6M0p+1FYsj1CdH5CigNWAHXVFoDbU/4a+nBtiGSehjBsXJik2xzg+lVbUWCsB
aPkUAOprNEBJ1KrLOuXUYAw093fSuGWuH/oYhZKm6d4/ZsFi7lc6k0XO3MFKw2QQ
QYis1kNbu99eMziyfbXNe3YX9uCWk9hBsPG9vzI59AbvpgW6etp748qTxP1Uysgo
fKx7aPF4CGTWFPE4aLLj3gm7dxmYwDAUJhM7wsHGoI1O7VJXBR0L7E/1bu0wosge
PT1R9dyjhC3WqvF7SeH7ngqfBUjW22xc1pBu8lk8+hXu4jaOe5lLXe3knh493Moq
SAWZJtLSwoNPRUf9xsa/QnkS5p/cmzZKdJ7medaVCBwNlNtu0ol4CcIrw+539PXq
PqS3rEiJ8h7NUnRby+bwKlVyzHFFhr5b+JLa5Xqn7Bk5shqqOMjBEX5QL/pmfq6T
lP7w8SqCUab7qF4qIQ1uaj6m4ZRQYwSja1XqNEI88L/qWhvc6uHj+MyHl0mOyEko
VKqapmo3dldfDK6erHVBoyuXUdQekYhLyrx2Cac5mOtma6+Jbn/R95SQVHQ1XN1u
XY8FBgmrvTYhjWLQssYgaWjgmPPdXo8ULF2eQ8k+pxdZvAg+AgeyuJ59qzkR8P2F
WHY1ErBiWUA/sAH1aRjN98b/SXrDTwqhy7SudE0XPcpDXVCe0wu6VPR0aWhhlIqW
j+5+x/JFu4gQ3N2v71qH37ditqH9tvtP/m/zzzyGx2WK4CVhlD0WmC9qFbkGb0m4
Gr93IxPXnv68fiHJlIdCk+j6s6X3pkawd+VCFXClRzTis9e0Z7RvzMqo8iA99rUk
iJTwaxnnt9xFBH10ab6AOXXBWQNfihTFoU5mNr7OBsD6wEhCJh8+wp5zEnORwTC5
M0jS0BTn64k1fqrJidx+8fBqRJvV504Da/SLnu+m5pjec+JU09ksJSo5QH++Evog
Ae3Ypdgus3Mmz6Sgcy+Xnd8/B03nFeALzPvDHsknT+Auprp0kMrmd2d0ZMNZogrL
j5Tk2IF/rxxa7zJf3HtfdtcTl6IBc06/7TLnahnU/tl4thcbFfyV3JxZCZiIWVuS
XksH19LTlAa0SAvbJtdcx1h6U/DIVjVx3nzBDfSVxvgmeMCbWSSnPG0ds6kXJOsh
EdkCOAlxoQHnX1Ofrt018VzdWEY/WYgMdWz273tGmSz3FearJYCQZmufU83S4cEl
50kp5tB8owwnyUZ9hhnEiYE70sJnEKMNqtTfr6JCdp+HzjVE/GKjs0M7veT1s7kw
CDnc7yzoxuOMvjAJ0H/lQ5A66uYIxzv1XAatoFPEyXzs5uP49eLh8azkIo+NEeOL
6JpXyniTARNRoDGxo7NivX2+ZPcpQxL2j/Z5nG8KWIGUAfJN/iib9Fb+NEO9tT12
429Aq/QbbLq2twaPAJfDUkyh7lcokuOB+Vzrc7WFnlkaXk2/6N+oP9rQi0sysLl9
z2Ek2HPLaE+Cm5b1U/bHtB/GnltaByhoyyyO6KpO/xz5ZEEk0EZQ7huqEAtdpnTQ
yjkM2hsYhORUaixtxaIyqT2HiVf8R8ffIgenjlfKGlLgxO7R3nwil34Y2LcIwXuN
gzWEhG+LIRqFVN9IHA0Qd46mLoM/cSkHYvdt32RulA99OWDSsQffMHoSPmzZDYbC
vlYQYkHx8VgMu5DzynHGzi+y1IxPBWG2uGK3mMfVjdh98S29j/MZP/6JfEY+2fNn
dPtOsuLFhiIZksUg9rDUUCTvmZq7fG9gmuMp2NlMIwTQMEvqdAp6BWbS9wMCmLVj
HBJy4JdsjHeOURivXr+TsNIOXOydT+d9++ZdbAticaLNl10sDaHkreUU56V1tZWU
DjIo6tX7tB1HImxiMTWIQw+ONCg2AT+Uj9ewD+LXxwjYOvEdV6cOt3mSjS8ZlHVl
rpMPLIZa5Y3G97XMtm8mGZy8a8ucmoZYRfNB8ezE6ruoNV2xiDV2hrkFECdUkvEt
VsV+9Qc9soMQc04pmyF/ddjsqHVSByNRb2Rbu/je/nWej5wcmapZqcPA6UUUTzar
V3wwarlGN2cXxpF4LnSEmPwN72mogb6JpmsYfjYEaZBKVXKetUWmcz+dS9GTxLcb
71rIMuJXSwPr0napBp4z+SsdnaEXc1FM2Rw1RZy9zwfh23xy8Odz5VHMVGhjsHlA
mWjMfMHo1VnQfUZay72LejwOq71eIjKUyhbbNrbKALQPcfz/DtKAjcueBF4iYb81
15OoF60Ekc67Owmu1T9l92eKLYbAcaM2dS1tdKbt8bhVXz/iiP8H13kZT3s7mHmf
A6S2V76+NOetoCCTEsPsjkMYVtud9oJyVo7+B+c5xiPhjBIQEUWXNkTfgVCOkpqF
pTVCjNC6N7a3ar5rON+vsc3nXpFTVSL1UOiKp5MRgG5QpWuCe+E+7uHxOhM8UfIh
J7H2KL9B7MClXLkY4n0DBm9QHI4GXUUXoJ+GczTyJqjVn2fUP9ZcsbSEYOrQnpDS
TDtpdWvVTG7awW7y57vzLfClAfnD4K9QEyUrTRPW/nXog2y80ZPHQAePIG/f1HSL
PeXgsWuT52KXJ4Ep8Tb3Tld1uwbxrzSomxT1TpKnEZXHuWc+lYYiqettX5tPYxlo
iJVPoVRP+8fbgRtImy9cefHcOmVoIwpDf0cfVAKHXse2lc009mzBfMGAtcdVvwyg
6A+A5i82k7z3JQAeTNIZEpW//cYPrXjqGQDn2Vi/dOwEybvXrFBP5H0R9UEwt1gU
fC5wgU6D5IjAWlODMsdqQTJvtMxSH4P+4KJ8iiX5+HTAxsxyz7P22tveB8U4yIbw
x51Z6R/53nuPuXGcUdZI8mxPGut07t/3JijIG8QaSalpQ60FhH+u9UDl/eLVpQ1x
RomQV1f3x24NrWV9cK3uD9+RBZnJfWqA78CdlpUkrdgcC51yWML2aqV3PI4MjfsL
FDcYuFrsO36Bi/7JJMPaL+uDVZsnh7StHsnpPxjotbhVwG89WjxPhgk7ZNc1pEO8
FflMG/ASDMD5G4Tifj6BmPJI7d4l+WLAc+i1vAQMCtZATjwPatb2KhmHoLl85UZW
Nu4t2N/FEuekMv69yHGhLqEFvFkR4Luo4mTQ+PlBFTUyn0FejFv8vmHwAydZy61y
QOyQ4PpI9FFNRORCkEjFa4DIgkQIWR8uK+xr3LT1QHj2WwcpOaYecXCy5n/tmzko
Hojomb3vXt9MVR/855/nz+f160KEbv96YQwqemzvW46Ddzfc8U9plYvWLE/Ws3+X
JzPEHqvNiITkqEEFWj/xkNh9ilnyKQO9Mw4qYToPlC03sy5HkU+MzHwpwFcXtkQJ
HPTeSOm0+K2wlqdo2tfLDkrfWhYMIS3xPJNwT+Cge2BMvZ2VLIPKSrqM11ImQv1T
QqCI0hJShXdg34xxq5dLdscrcFzB1jTEPeirdhLslPvZbDgT1gS0phaRRbSa+aq4
bbP3f+yZoMfKolwu9ovr5Ve8jbhI92KXaPbssemm/T8F/p92rSFdZM605OJMFpXu
MsIr8o0zcwY1TxPEdWet34UD1iOIJYC0hnCAtNb5X1aDqounE1UpjgGZnHVz9YMI
IAR+QkkYn65FXI2LmmPWXcyMEmLIYc4OIroraF+6TJklCs3nM+ZFWGgwZ6n72GAk
dH42po/Ts7efylSkulSwNKHrBraKODSCxqqvxth0fv6NTgb0eGkn5NH5FW5G3wEA
dylGwbhSa1v7XtYI1nOreJbblR5vMBsL7pKzYJudOwIbCeIuF+06rVaRCpSvPZA6
Yrifmxh0y0s9wqwdv9K4xDiRMqkBOGjOS3kFn+hA1ExJRzjJvv+8sL4T6XYadWrM
jz3lb9ElbgB1hRgSyBvok0AV2KMv+yGNDoe1DLRxUN1ZDM2iSDmO1N72TumNP9l/
IEAjMLnlLyTBEn5dE1K4JQ4FyN0aELX74nl+0+p9sNBhNUXr89WSKOoIAKW6KJ9a
GxzIrQ0tVJ2UzAbqwqLIdQSTuO1XwktnNgWtqgXn8Zbm+qs1ac87hR0UojB3TuPT
Xx495kT0lbgv4+IaLXFM9JPmVC0ZM1yjfUf2Cg29mEW3qSjWRqbgnDbTwSuZIQJT
/P9YpBmMpgM83OeT4dVW4tJ2k6SSTK5lrso5Zf7CLOzgS9aH5YACzEKzNX1DbEnx
QTeYUas5Bxx0PdjkWzjnET2tBHqE+pPEuQ+bJiEtYmMvFrk++Iq2Y61dcUw8HQzk
QQo0TsP9BSRVpnuQwQ61vR5Ei+eMHvvde9ZeV7lm23Z4hRkx3PpEp8F46rekh+zg
yfMdDECiCty6W5SS5Jk0zaZD5fzBCwk6mTTCpqiVKR74OZAYXWwORI/2JIw70rts
3qaGzkT47/70u74FmIb9eWznWq30oBjqr1EWyQY3jb4iBELju1m4ekz+qKTBuzv+
SJOrUlD4i6aHQnZjjllrcUTJBIq7SfmxRmAZik6G/rPO59k7KOkHKF1RdawUWNSy
4lKuV2xOfMEdAjz85qjb4f9t/dISzQGulo9NK2SpgZPdd7S7KxrzXqaLHchO1NDx
KbJ7GKk9Nq9KbQRBu4hzLmo0bQjUUQBbJFRe/6OFVhFiK5H4MR2FJDbw+zfreU/i
jyD3HQzXLBhrre8yL+PABs3k+pX/J3EfR7t3qQD+C+AmFiyqzWyLYgnf2YkTh32u
b52hoJKBjYOpWuwMdE3RMfXemskCX2lESxJq6xml+xM8s5mvpTFv2KvOdka9yRYT
D85OjUQV4fkWbj2B7pHv8wWjqjTkB0FAr56AOLq1fAn7v+8yxvlWN5w//wSdRD0p
RoBzStb+FMu+wNmks/FLbsgogTXWvLm4q98Opnt+mCQd70lZXc4Z14lIbiwuWngs
5bY49e9eNojoKc/tpoOd90xBMlxykWbykG1KkmCCPY9bFjML6YxVRQctA+HKugUt
DOtJTFjN8INvgp3TzkUczb/ec/hZCC38z7oqx/Q6Er39m1eTLudZB62AUeiSdtEq
oxbbpKnxghWa0z5ppwEK7/df2gO1pC+UH/x6eAJuIwDYES9DV4CcrQ8P62qJjAfn
kB9YtQRajaKL8i82dRqa5oiMGjtyJEdtcsv3VwzAq9mvA8iD4dujzm6MY9mPl9Vz
wUZQuLqUWY2wB9tPDVJrEAtTdxlWyzUbSz5P4f3RXvdHZNlG8hctfN7Pmhhxjxp8
6xWuRn15f5TL8fA3mf7m+yF5cWIcMl4Ms9niEsgJmLOEmqy84YqUYIT3EHJjmr8P
HqBP83vQ1gHCQPO32Suj4RDjbr7da+PJ+vae6q8qPYsr3O3OxXQ6hhl4NYkpLsla
4j63iSBkxGS5Wns2cg9okGDC963HcEAiOl0aGRzMaVHWlQl37/wEtOWoPlJFXIUc
8HE4LVURs220o7+/1djhlFF4EX5C/m1NJOKpczIaak6FP6qumNjcZi33ueouhNCh
y0VTTyoY4cev+AO+SFw3PWnEN6yn4U1QcmYyzXDh/yIZW46ts1MTtcA7mtm6royN
nLAOFDFoUCqRvfkd0TrWyCgQ6kg4LIX+w+3vlhRrL66deZOPw0yjr4g/Fc3pjHV6
Zky64bE8Ttp+FXjZguvNKqe4DnlJ+AVpVNuGHuFZEo8tcVwOpr9/b1J6VKn+/eSL
kCjdUvs69ncg9Xwvo/dBu9AzRFDW3cn/xDkuvZp2eMNsaFuVMyRH0aVOkoUqaegz
LWnUVuGRVD2KWN8s5uk8SOFJLXpPh8vFTVFzLjcNWOJfFXcPMgU8iunCDNyR51ff
qzjvzY7oFIZ7UhETJcYoWchMA3FWjpIUyIq7Y/AEv3/hhGirSce5eM9mcRu8qUFM
flfQgF3jj0o1cYWz9xLkffnwFySprhUDuu75YQGErZ/EsBIElNi+5ztuan/sh7LF
r3JAyUb876NPOwOhjXsRPOi0CYfySqz+tRYvkZm1RJqFsO7WRSbYgJg/m+95K4Y3
xOobDFZRhm+H7hoCrYVEMeeq9JzNkDxHFIDGqCPJc/7jk+PqUnKioG8cVGdH1FX2
0qa1T1L0QrlA6m6vwuClES75+C2ENCKwELNYfEBOqbgMLOIORECG5H55CvsDLfRf
7kefFwcU9KSesozyjTMlzcVNmfJ1j1rPTduYYqTylCgF4bXJUyefee1K+A4peRgs
pkRYKvEgZoAV3qW8HIzRnVONSguSjfjVuPfvDdJK+olZb8yCecHlGH/UqUtizUVO
4GB4OmEUDj9TFjX5AzLSBtjcMTtklVu3Yn9tOQr4HU3SYCHwJVT4Yl6eYXrykeFS
D93zlWMc6wXujKF+pIodpgTw98IJG+YA09fY6YySnsRZL3N09sb02LIllIiAmWuY
NOuc5cv8+67qvek7G937vp1dXD9WblTH7YyZdXeWEt/HxCDgkSg80eDzuxXoI8Hc
yiaKTT6M/71IuzEqJu+4vnsaxTYp9dyrAt2gveQX8qkR9uayzz2iDSJysaO3stfr
Ndq5aoIGMTq+MriFZswy0Mklm4TcWvvc+LpcBW3bhrUegjXMH5XcbX4+absT1BQU
GoodjmT36N/zeOyCw2jqUqW3uTcW8V+gcN1DFJjltl+CgRl/NRezuWrrHWgSQjOn
7Du/8/TmdPwvN0qbckn/4Y0s5K/SLKhTll1EgNzYeLr4h5P9fCmb5xbLfkN5OMmi
qgnzciz2wc211xOvH/M15VQdY3brcvHLnMD+lQ5QU+NncLx3PjrmRuczYrt69Mv3
rsa3T3nZNmRO885vsmjfyHY4AYPRgvI6ouHtk9WeDEt+3imanwzLMrvU1m4oDzDM
h1aKSYEeNpAi4jjpwXc1d+/a0QI5Omu8ZhuKfzf4tm7bpMhVmxxVpVIb7JfCEn1q
CDChbZmF3Rjv7Xy9i0oPAQ7ZhF540qOdU6eW70QerIplYqTh1tyfL35O0VCcM7Uz
tFm+Iggb1+l1wKsli5Y9vMThUy8TYxbPgMv3C8RAkUA+UOFfc8JF4C4RgicIwSeD
9tKYBmdHO0Ylljo98CRZqzybCDCo/ZUOXaRPxALsiVltfCvjNNBZAm8DKsqm4lHQ
Y1XUVcZpp7f1JBn5w79EJzhndh25jT0YMOJ+AuvZN/PU4MI0UhyjB3s16jPyonte
tgKsCcxudfzhddEqA6+HDCnFN0lZPGZXa0ngsoq/RTuDhN7Pg+ForZ3uAkZDdxLL
Fd7Pwix0RaL3yCvcHlRw4Akt65VekOLcoRW1If1YuNo/AfOYZYovr9kb5JhBXMN4
Pyr+DBmE+H1Qjta4yL992vFF5aXzjgykuh+87QwbWiZuRrVXdOtEQdVGmpEkJ+MW
As+LUGy1EaiBOokk8HnKgI1LEV+vEudgYB6aplTS/hXq2o69eBp8nNQfwVaVMcsH
QU1M+hGGNNpwbsUqvrIV0wP1aZnYU+grovmB8vI+mlnCUp80P1sxDoaAeTUQY73w
2vqkJBH+U8BEUqz4t2KumVD6GncNeh385TkN6JrdfgGfoGOhcY9H1pyEd9ssf9+D
WwKNCKGuOgyRu4Bx7WDGKgyOWSn2S+7KOTVpOcooqA2qCmYpQuQGu8rbkmEstbKr
djP9y7HvYTHC+QkOOMC3ikAAknAgacttkb7YQKBNJzKSf7mAx4+t66hpJ7QNIwPw
wfGNHzJdQF1sZFoQTQSQbCP3/ir5diBPqjVzZlzfoA1/tuGY4HP1Ggxbx0eg9XNw
XlIZNyTrAfUZv2mJAvOAH7aAtY3ddPFFt6SgIFuvHDB09A5SZS75in/BbgaYIHzL
0G5mYKEgb+X/ISuokUc4OF3knjiLuf4txhf+UaZtf4k2gKkMgyOf5icuXasiRqoU
iBYveW6BYU+kQUNUctg8Im29DRP7LWfED64qkVy6oJv6+aKHarVkcFrSMueTF1Ng
Bc4JdbtPXk/5qO2+4k9VeIj3GQxKKMX8yyiwFk5OexexiV0W//lP+O3HcE62LAF6
kogwvqGUDQDy0fxHhaANAucXdF4E9ZKtl4BgD7HQ9tk22MVd5atmR/80y90r46lT
qvEHxMRqt2owtISr+snAvwHO4pHGM1vujisrrtb+dCRiXqwmkaFoJA4Q0GdH6oJ9
92MjYalpy0U+89wd1nDbr3nvC6f7LfC3WxwoxwBitRQaY6+FQJr/hVJVSRhIiNc/
byKrVKc0DG8h3EfQV00okgY7/iQfwRYTSH5eGBrz3FHiOo6wreAu0sn35K6XdbJh
MqtSAv8WpsPdVMEVQjWdd4vbi/UpgkISqChvzaAGQuF0gD5q/x7U3nQhulOf5QTg
qlT1AT1kX2Vu2qvFRrkefuW35dPww0CJ3YzX/4Wm7ienQE/lg2u3EnlorbvIDZZK
aBUkYgz+eE3tZsKSbBgUympwvrMXkaoFUIxsJ5vq9HmdoDxxXCYg/YUYSq/S+vtZ
pixlGJe3CwdHIMG5YKItiFvzQcPJAz40RaKPZ3+kob5m0Ifsdl/GOmIf9UyzBOvn
1Gpb5dDq4gA3J9u3ImryXU3EfVyplrNR1Pux6rpD6dEkYTDlLw6WOJYsVeFM5tKj
NKqwp166f3qO9by/74HhZQuHfl4NTKw0ppoHMw1HnhnXkR9eA0ln9ckgQgtAL+AN
znziry8llViCmOp5joj1tU7O+biBeQXtrwi6LUpssC7XmWKEBLOxaHeiZuMpMtUX
+UkLVk+uF6rd3SFvX0YX5dH3RfmXfXswgaUCSbPPfCYmSyr3kvnEZl19bI+iZqgx
0yOpfL83WpUmW8J4qDhdmhcTW8rZ7pmdfXt1YGS+OofomLB8+FmR2tJZUxFXQl1S
GUHOqf3mmHCVYtQaV1bxxsflU2dx97eRQE5ExZ2RPqX8YYYixZqf+VQtacXC2fyL
WX8lwKc+7qKAFV2bWRMz2a/vGryjHuweMecmjxXhEvT0qRa2RHfSLnYvyQ8xlhj6
oAhoQzgNK2WuolV3Ev6QftwlT0YXdk9aaAcS7ufKVI5MWDeYns7lkR6DFgfieubD
FH+Wp9d8jZ7J/aJm5vjDiRltxKpBWEQZ5CqO0EHF0KbjFTdrMLE/wUMwmEIRgusu
VmJ0PbACBjStIDoaFY7JLbE76FKYLBrZSAwjHs1JEN2Jmp/EVpGzuIc8ReNyNU46
AHv8zrNjXXElpS/TTirXtdvS160609LSvQGfVctdXaBV0E30C3of1EWJclzmKMWT
OOEB+i5hbssdC5LiWUtGn19x+ogMKJwpw8aOJgZ4A2Y1gLyHxXK2IrSmSdtZ9/Pw
U0zjpmZ/eG2AnWHZZhhr49ZacRNK3ykfZLC/oCo0zc6JcXBHSdbjpVZBKq7C9lM6
/iSkcJtj11Q9xHhVnwjrs3Oa+pRthnFTh9oyrQ2ereq559cI5L5lFFx7IAMseS+i
AdpGRC/Fj6vrNshk12JGjc3n5MvKYBrZN7RkQVwd6OiWCJIukp3Hfp9pmKqS7DJF
ubD4jhFFTQOl7FD4bnxjo9itj//580StppOd/m453e2EJnM8RLmCDG0wCbwZqqgv
gGHNzkfsF8Ao4zo2PGLu45JKxn36jXlHVpxYdw81pygKrZJv2ddvag4ED4jAV7ZW
RIf3wuiwmZvdBNfRU7Cum7qJPEb6MH5E8Mgds6i6guil7JfkAt8wewPiWa96xp2S
wQqydw9CckRauCb9q9u9Z7QZrRDFLt4Ixg02uQ77OUaxm5MXEKl503yGboq1l5VF
HDAGcRlbp8Wo5uYXkGAiKlYtNK1dtWUItTfnyBUxh8+MEueea3dHQqvbdLg90SYB
3s17eCNH+QUzPbdLBDC5oph47ltOAJYv2KJstPDEAEnumjCguJ7vXdVscSl1K/AM
fTKTRDFBwQReL73fz7lPdXtvQBUTo0Fa21PDu6lnjInwE+p54hQj2nRtJjXznCXF
qEDfpFXXzyvA/2InHdxfhJ4l8RyEYYyhOp430gMDaXvHf0n0Nq/Vll/ognD8kOj7
aDLxs4wn7hbvXTxz8YJanmmbpQIu2Hhhdxpy27U6dvGSQfisSVjIZygnbxABhkk9
hisQCuab0KySg9IcrmC0ZpScDyA3JLZnqzyPIyVq9Iavb9HZrEdR1h44l+L/Alb2
XPb2DJZ/gixbib+DvlRlpRF5/nJT4EvMnlS6wvrWivLfRhk0/W7Gohu9w9q129sI
jRhATqs8QCXM06aYQew7WhmJgKvisUvBzY+z3yoASfupIH3iA5Mz/uTKsc8TFQBU
gpA3W3mfAnbIAzofhTWNjd1wdRsKlp27V0ZAUKeMI2Js0+ugYsVqkkSfwonQ1Ow9
DiJU8fyLyLSIVfuYr8kNblt+X5szdGcY7zq2yuL5x6R1sUiUd61QR0/YtR7rsF88
tgjm4Y2KHwXJw6FM0pZDs7/Dnp9GnoTKzigWtXgAC1oLtkngynhpLSBpVeUEv3y3
kJr+rJb6Zl1JIqvEX02gKlQa5GR4E7t3ts2w6gh90D6/vCZPC1wf07T+ueYy/zzF
cFWlUv8jcnBk/UjZgDhN5CIYMEFPs5rd5m3yrsAYstMxkcj1aAIyxlHqj7dCyCkO
qJsvX4UscFqfFzdpEcIaJ/m+L2OSsqZzFg6Oq5rEQtb8R1d8r4gnJO8TfE/6zt0A
wkV2vQpMpviJV7uijLs757Ausye7Nvi/We/OyUoFWNytnX5M4YzjHGxWAxjiN6zC
mavLh/YoO1C1K1uvBQ8tT22tzil+NAUVc89x++Eio1qmMJ7udm36YTOWiPKOYgHb
ciV3IecVBdljS0v5pltGRe0uA1HUibm9PLIL7votaBAFmOD72JIchLcDA1ILQMKD
4z+QOqEeStYG7/pMxflh1fj+LzI6GZdp6qn0u4ZW5P+Gd4hxASBeXMdohYU5TByo
0mGvVlgjtEgR5Z9XXbtCbYShpf1CKfP+cFEA7QqxKuq3xl9qbXCA+4H2uKfq1xFv
rut0gfaFc0VHJOprfW6aSMocyOHOMQlvZSZX71UE0v0CD8dPHYaR+wpWmEH+Yygq
mYq0sUj0Oe2D8D2x5sir8cGz1IdCezFkAV2BolDYtGE1u/rAdNtYSqNb1pqvRMPb
aoD3AU37RxT2FYEXyzPmBdVebLefiJv9vmwvhYpnZYFkt/5Xryim7VfACG7rZ/KU
O4p0vmGVQGdsOAvcyLiIQ6iEcwdzoVHDXGwdtVTI4/0morlWOgtcg/oqpK1zLRJL
ZKMMhOdwGfDdeZPOU05Cb85CwqCnlWtMj3aRWdWuH4RTFO1l0NaUQhTU0p6gY+iO
gcWIst+zwQMbSQz9FV4iPK6k9UYkZwVzUM4h0S3+9UpbUCkz7W281+f4e+lZ0Gl2
J3MTcRb29Wfc99rQH7LziVTEJ9GVcWm95GY1DUNeq0kQGg0MALGl98RB0rSzQm5E
sHD+KsJEMHbs5lo2xTXlUEkZhgrcXxop02KqdKEE69owiWLmzjiwzzR2ETLeN1Hr
LWn0kbfGiJQtKM5tRvFClS/uRH7Y5725zYut0/EKti2tSmFyiHxQELfYI2KLV8Jt
gaRwqP/FTzcH5oK6W+WrDPiMgZZq9yjWVP7v0nIZeM7ZrhOLIG7JjUy781131qsp
DOp5TZC4nswsKu29CxnDzdFfrxNHkNmMc8U3tSf35gTiOJVtVMpj48gesjLVnAYa
EXx3Qg17f2b2a9GgsbJHPVoqZbKo2NCSJYTyYsVANB+Xsj+fZQv3BmhAY01wWBSN
Yg9RFv58kckg0ek6T0Q8OAFirtWyiZQpTWGv0qigqVRLbl1PaJUJZtuTydGUZ2Jg
3DiYoRhUnK9R2y8WgK7999nzYmxK8rjGlOQbgkoF3QRivsX43BHrSwiEuMOBckZ7
o4XBqHuHPOhZGGiF0tyPfT1boW5gi2WNsiemTLLDmlDf7g3VLRgQlULU68CKVboF
i2R99o+TPeKbBiRBcs2rfYNhDR6zW6KfH2HmRp9Mr5JSzEND4iO3dcr6ktjB5W5X
RPkmvGwbQE60GNpmg23CcbMllf/mEJaYhJJ9esIcAh1hQgSogaTsRd5SoxoHzy92
MIsGiLy/xF1jQFTXYh28XsrX+ra6nyyb4dm/zKWJUnHZA/OJaYUid13Zdl3hQ6jh
Of2Dlbb+pOYFHF1ldxniPl1y/but8BvcmvU0X1UBe2K8mcvp+J7UYqb2YpMa5bnP
Hf3hgrorht6tIaM8SWhKYWZ7g8mUfd/WxaB0NmgRC7ejGGt2OrZqNfG5mLFRksOW
sdXvcbyHAfAfiONJFe5Ainth+6CoACEdVfmhrjM12peZ8TpFY9Owmr1qDNzh4oCf
NENl5qfMKphVtgi50MdkefEzHl3bwe5xCFJxm8rzBVc8cRsatNMHFqRtO6ydvT+a
FUVyZGkjmTxyu4SJV4IzcX3UdSGGMHbk8y6PeTCmkD4QrVSStSSubhCo2UHYOoFh
pl798rrLs3/S1ifVIVkbL1Vd+Cwd1oWYiUyk6eUeGej9OJDWH+yMZv2m9dEF6wdF
89kODsaV5f/xLc2J4AW2re30HllKp7Yk2YIIEYgqgA4IK3CPLz6jT1f1XL4Jbu0w
YfrfOCRhm5q3SpUbG38+cng8BTDLsi5QH94YbH+cz2hBtxKyVCOdD9yH3bYDumai
Noy7cp0MBLABeRu114ywSQGcPS6ixhJwDx43RDFSp1uc9g1E2/tAlfVn+A9/AiwI
5+hIwdrJTnzXiBGvmGg0uJTM+iPVgldWLeMs4fiOyuLWAd77qLpZyjNU1iDi6y6/
1qkvBDDJQkLI/Zj113ukISwgwEJMNk+hNWw4QdEqug+zXzA5U1hOa5cX72yAuk2A
R7YIaoJ42GKuhYp8OriRcAzIJAE8JOtNMETla6NhafD8EW3+pJfaPmqDYZkDcPaU
vvNC9t111HaPOswmepQlS3QjITNiPj/eLKmJjDGZU00uVipUxshn+coYufTwrMmY
fQYehluCP7ALr2Ajr5bdq2um+vqQM+FW9zoBPdnkoMLgQl/fknnWTw2kz9I9Ub44
2W883pa3zo4dJnem1tyD6w4s3LQYigDVLzPcg1T0Eupt7DsOP4eYf7k2LXWNNAmQ
52u5g+T5ikNOMh+z277e2FcAxpF4WntruIWB+ByjlaH9cDVMWIhowz6RFL46hGhq
G7jF5ShOFbcxCp+C/PdWy3/RYdXGofhn6KGfr9E/BOpM24gOrnt/OAXz0n7FUjzW
NYNzdCms2DYySSZ//Kpgy5W0X8I2hWqJJEUCdgK0rycKTrMjV78jg/7aFb5Ut5fu
PXBPuLOhMvcjq0aAMkEYpVpoTNV3SbEHNfUgS99rw9DJlqQax9aggr4oRYOLLvjl
UQPNvuof/estpiT5ed2v08g03lO5ILIj2elswzoHAWxZ+ycYCYM+RL7BOGsnDfPk
MCi+eiBJqleQARVhq/z2WeeCOQ5RpYwEhiX2YxS+W5+8tKnWeShtxWhqjiukNeT3
U5l5Iwc4D2fM6OgqIr/DOK+mJNFDVTdRLCJ3qrtqAlRSn2xgz4IG94xjkohPD3m7
tDphpnMjM9jC8Da+MNPx2mLs1oTcsf7Wck3f3esmnHgmjj8TBnGTd7FN56Gw5Xb7
K9wUsllx/7NQ+7ZWy59KeZPOB3M0x8iFK739H1ygK83fUrSiyBA/s5dGG0eRB8mv
5pqH4eBk30xj7CqfHhJ8vz73qdwD7ARZrSFBO8hJp48cRHBQaGH5IHvOkcBIf3/y
4D6cuwdtR02V+D6zwPOZhrLvFeQ4B3ldINUG7emktUUSAR+C6tT6Vc23iv6qJvLK
qK3irty+SQzdrTY2BQz1yKkbjQa1YWfsPZolMOkifz7EhxRN9r77mIYTzjKm6azO
6/MqTqnY5ZcihZCTKk7DNpUeJcjIcb5m0PsDeYhNsBiOVYM/SGkk7sQMnt/dIm9+
AVlnxYM+f4XWcxh4w9iL+3GdlYW8hZ/TICeoddL48DTDXYlpb2+Xa7Sjk++Kw6sY
XLYq+9v6OjW03ilbwXqb/qsbHfUBb3m89PXDWLO0CNVhbPr/sX64euNR5Kgp1qG4
r1qUgCLWYjiCFy6LvgV9UFnC7VtFvFang2gzXPx90nVA3yAy3pAGR5pOIP1oTEW1
8Q4yTuwz76PQzuznAzvteNsoL6RNqmAoTSmXocHqfiGsWQIstp4jrdZiT7nLolay
JMUCvTE9c9UtK0vkMECsJ2tsE6yKq/MLSLQVR4bcXE3tFPOtksHAd1QcteBVGJU1
JHtum1KR9F0fqHUNV5o3gzQ2nNYLwEOHV2817P+PYA8we0Gcjk5oIBL5qO0Ev2gY
hlGytJm5Sv+mOkgTDQNBcsWwdzhvF5uFRkjCD5IYoqgnC2/SZQ4Vh2/A7hUATUkg
j7bzOV1j9EHrdeQXFKP8G1F/s/qgR8kLKFfxwy+LcTAshqo88kUnngrPrahR0ZWP
H3JvO/7dKvNFA6i3tXA/namfb6+j3QgWpDFsmUqtPcgoKZbgo2424b5yUW+RE/cU
KTvoD5k5aGCj5ennvLoEEdYL9iaWlDfx0RbTlK8rmUOM4Q9YMLWp9/USXnr58Big
7vgBY5Uv61Zny7/+CE6BFynbqyGzgg/H0lXIQsqhmcGCyBVc/OLbCbsHTCuAwuub
M2qWxpONbrI9P1v8VFWvyDEquCwDCeVOjHsAAkpD5NIPeNYEPYIALRx6itX6UcMm
R2eLu6NuxRWJdKgBZQRqoixYy5C5vSiEGk7WnPBn07QZFRQ++BC1BMPAXasMCt5f
IK7vSR4k0mApV5thHJ+twfmU7o0F9l6Ws0f4GIzsUO9o7GsTAK0Eb0wQVCoOfsb3
8cnkS7PTnhjm71U+edkAmrAT/wQamQ7BBa3RTpVqA5bKhF2cycU8rs/1k8lqbvuQ
7a8ScUav7U/VH3uCMJVaWq6zzfX1Ha146VDQp1iCjsYQ8x4UWfM9Wns//NCR4DpM
ocb9E3gw7i5BZ1DWmErEdSWL9nLVVH7HHNZlQpIrMs3exhbrWf7frvLweUEh5JPr
oVJG3xeylLKlXB2pREFL7AzADUF9aM+JYqax8vE++2nUr/pym/8+2lIWtbQ0ccDZ
HIyb1Hmei/ChSeGqNYVgT8KdoVYuX43+y3p8c2D2IzPo0XHsReuDWJnsG2KJOMmU
Di/iJHQj2m5WletwJRPK35BWoa0NXKLOY+L1AMJDk+HCyxczOqBhahayJ8FI6wJH
2ksQT4Y8IwxTFMvo3lFOhP7qJMBzVoIvXakYKNbwkvwykKeeKdxShQARAfv2vpjR
Al/C0yZerTiBhH5zgKwFeII4fyGH7Rht1Zd/ex/gKqYyu9q2lgc9wfLl/SHuziWH
wbFJA/LGpQJqiZahmd6g/mVZDAMwi/dgIh1a+FQ2gOh3+jU+wn4QhmTC+vpG7bEq
b2345LLybxdMMQteUsJQQ1YrS6HUJtQZSgXEI55eAWOrhXwSxZgwXTZ1QAl6glyM
Ym8ONt7oT5hQOL3Y+XiWbyPi+s2MDnED70j+obITqs6jtggM7a7rSVG5NxhSBYYD
dUW+wPwtLsuiNk7VtJDO7BnAYj7yOMsgM6sUoRRC9Hc5cTjuyUumPfUXRmEMBUdZ
kKvJ6xbOR2slZC8RkwgiRuetAQW5NWNneKoD0PVKRPtLhMRp57d1CuSPuE05Nat8
9uGAd2pTSJ8cM6iwQeU5rdyu/RcDF+xUcZ9mrTCEDCatu7bYe7qJgHVMuL0khQo1
zKUwIUft13BpcgB6XY6ldL/MnV8pTlbhdLTr0l8fVj3uB6kz52QWxjEmoXmgM7oR
geiiGMvBYAMsD5hW1LxKsah6m0RqXENX7sKcnOu078PEeHS54aXyXTfqMtA/9ct3
0rpk5GlW6wZdL1lw+QJVm7PISVOJpDNK9nB6vrdSbAg7LFPncZrrFa1qxz+yoC8T
wrLQjBCegrW84YLcLe0f4jIiRb78lginNakCJ29BfCavgSRZU5zt/G/yGRNe1gBO
yNbbLZMdPXlGqOrQIrnkakZEUuJIIIbY+h+eHhRZoMqCTJId3sInTCZFXHMXg5/1
XVxNXQA8yV9upJUB+mNNtVVDJ7YOsr/sxpVar4L4vMgyUM6SBsNLjaTuY5oJ8SRx
8BD40obQ7gTaHxgUxcgOMDRnp/xfHYyAX7DgYBhYBXV84vmN08j3X6yMXQuH7LdQ
OR7jg7e4vdhN3lxSwre9y0keOgxb05nZxhv5jRuEHKqXWYafEQl/sMcK5/uHkDh2
BMF7dsQ5xFy+32NLM7fGAA42F1r7zHwZt8KJOz4TCyl80Ly9gFbYe3y2hsfHuAX7
8dQpeHlkqSHXNQqKYmknfvxAkIpjvUE3tSMYnsECJ5v7n5M9xiVrmJOUy49b0Rs5
ti6lClspgXOJlsPCCmab4FJ3xcU1/HyS+89KPAkdlgXwdeq6Av9F/fZydN9TwjFB
+crCWcNO+MZ8voqtmY6lBKXEKMqR+QVS+N+VT5/4FncCfjn/rYBfXw7l/nPB5o5+
mIEXqavra4oKooB/sPgCburZDKzikiC7PopAetxdUYmA8NbxVzuJsgTV5WhUs3VU
JYtOWWzahTDWwdl+o4pxjptS+BBOgP1joYYkcLAm9TUfrlzCO/W1kw6mIHVRzaFT
9GPs1PImk7QSlXKNIXBET0e+bSKamP3Bz1jq/jR9eEAIqdzyq0sizJnfiKQnek3m
SIzBVbC6rnosw+l0RMBaxKyQhXm28q8qF6tFSDJzW+4iDA01YmJ6oKbDk+aEiRpP
yOv8Px5KNkAfkRDiBUw7nuw00gL15RQaPKfI/oTo1aySQdG1VeK9Kw8+429+jTpD
ctkBemIfFRizIO6bWgYdjETzCRkbBiipoSf3jXeFC0CgT4BhRSOds4kXHbQ7bNwP
NYNTa1o+Tz0BWJ0RSVcS78wNCoJFCsemNWpau34hggs/v6CIMrJY/wL1DZ30T/W6
Tgcj+7V+11jZBrc51Ktx1VSCxPUsqUzPdepfru5ocS/EYiJqc0V7GNd1VGYy3AIt
VOXpV5vRUGU6dRSr/FyPZKzMq/ITL+Rn/aNUW3FR06FOaeV96RuOeuzUQtRM1vhc
CZN0T90lGdUzc/ggJcroFSOIo5/mDoMzimm4u0U7fkGYxrEwG2FP4mAh4/1CxIi3
cpNCt/kd3GFZ/2jREGvOplm1zMAR0SR/JEBFxfWHHrsz8r1bF1EMWZvanIWLaCVb
GiXHA3KXVwcL1MgKMUWLqV01J0RZ9TY/rB14oH8yla/CvMiu4aWz47IvKJsffB76
VRdpGbutlYFiUFrwI+qikFFv3/tsTvr/R1OzWF7LilvdCcYq3tfFEwB6bScj9qrk
AW6G576YKVjU/j7x9mU5sXNs16OPW1SVZQbP3hsuiBqjiaADMqQRuowRCWuSdmMZ
GpcCH/pslldmDBYZKSMmzGTl54+5pwlY0ggZIqr1a40yUWys9neR68ap3V8+eC5I
+dQgn+C3Xq0NTn30WvEXyTI6FLtNeYz/ZzXazVE2FVfBhc5xJ88GLRRijH4N8ZjI
l1X6O1+3TBy6w4tugi4siT5JgBgbn+vc19UDZv3MIOHfpFBm5dM6G7NeWoQeQZLZ
1lEdlBGpQSLYmrJG3uLNaboG35lZNHiVviwWEtG74yS1Tj22odeQsYX+/hsppM77
9n8a45HdtT6oeQXglc1XRylXfHOq2/cmYa96cLlASqSS1DLBcBn68hhYrwh4Tpj9
zPJoFv/A7foGEF/cdM5PeUFRp+ifeZaSaLobRa3dMUlg75mnSFuoxrDDuoZ6GXwp
eywxg/W7Ls7di71poon1mufQEpnIYQkUSWA2xsG2Wp6gDDgN+b341+09o1z8YQSJ
Og06bRgZJdfORZCBiqlW55MMtunZ5vylvg4DHpklmU7GxAWjhOabcJ1NiHrNvZqR
d7qLhdUfO772rmShBypAXH6nTADk58xAMTMVTBHDfsj/dSKmB+s8R5OZlP8Ifx7d
LOnCKOF5JU7rU3AerB1RdF4q4/usdE2hZqsvgG4S16NZEcopELKSLZ9SnRwTL2fx
qXbwSJfOsGX6ihpLWMdUORQ5M0zS6EZl/Hr3lDEuGLbgCPT/AdE5zGS6W7K0ZWcH
kqcrYYUtNG6++uHo9byMOLjqefyukmPZZGOzRlgFB1Fr6PpnvPpqq41H6prBrRQJ
bmzCWesSNfR2VCQyd/KGCauop8aIqUtGbolr+vDEXrtElE9KQ/HbJNu6Wi7AMbVu
hAuNIyNRmOGIC9KTcrbL7IXCxqxoQTo44DlqUruZsIruR5fNCK+yaRlKIKcxHljP
R1E1TgwQyHrh8XPWrsHrK2/c5X5PPAvr11RnKjtuSinDNGK+6+9IX7J1ZGjtGUNH
SxF7zCZslNTv6TTf1fYrkna5KX6y3UGwP3L19lBClPHaaXwrgPJJp693SAwSJUdK
Lmkr26TGRwc7nV8le5INrNmWbKJ+DfzwLVgbw1BVoVdAzKTMUSDjf3xKitsVSD9g
GfM9mWw8+iL5HGziJYowYFaiVxSKAETWiRuVCEfiWq0LzlX3fAwv6LpYyei6ZDrK
6poyepHjsE0YtlIDR63B5KPMjm6MU3lwaEzCCKI0Ji5k8B9SHLEs8lFc1vdn94ko
K9MUhYxrOw79CP1vkt7ltZRg24+OArsxU8iYoXQ0UmWQlduL6Rn3S3kxSjFfXJZk
gNGMs87IaxG80E1mmw9TBMbQPUdSXiEDXuQ/Bnau8fQ0mCYQFhle7XybFP4fWjUW
hLv91j9PhJJ5KgY4IqCxgAtbhhrfwVRJvgQnFbSXaejnPn2ssBlWgac9sXNMj17v
UuJ2vpItJBl92MowzPB7Z9c4SE7O+Nn78DpAOVBG+LbaUUeybsEzoGlqk2hQ8wa5
MRj7fZG254SfvK8sBrC7Fhqv3YgFKo8n0hhG01B40xRy722wTkPZOIiXz8rGwter
I82oiQNLDbJW9dGC3Cr1+8P8Z0yzAXY0L0aS3KP8nx+Iop9xBrGyhR3u7/KTvotF
EDmh9ZXfmWAMvKbLtsZyRkS7kaOqKX9Fm7BB0/gxetGTMed6uaBoferlFQmFtNwU
xfnjGXBXW8hJy3s63jSTldp1pw+ObVLWbrOUAK0aiSTTHnk5qIzXz//eTDiMZTMn
81bA4a5WQ3r5Fa/s3895r6WxR7wZTWbQFdNd8x+8GvodYU7UgmnfPSACQJW4OD3S
fNkjmJ1hh9nkBSDKSuVy7IiJXqmvpaLIdT7c9Tb2sEDjH/rpdw2GjeHf9hZOSDpa
OIbGrE7ekX9snVOmVUb9i264CeGt1METDgelidx04O9DuMiiOCb8pLgGUR7k4In0
UCT8opDOecU9UeJvR8ySrkIp8oEnQJJNmFUHHpTRdP5sJgMG+qSiS68pMMHEo9li
LYmXwx5KskokvN41lS41MZZ/R1mzPe3H1cGzTKRJ1Hgh+ibYC/SC01otG/KNF0fJ
3OWgLdfo2JbUjWfNOh/eOT6nS8kGhX/cmftjfaM7M3koKibNSvnJ/0BodtRb+Zva
17db42pv3jIeErkxhDg5N5k97Ia+mtDleSMKQFqP11D4U0qMt746KnemM+n8Tg3e
q+VlZ3qL1pUl/cmScx+7dxD08PSAYM6xVwaSfFVkgYe0VgchTtJ93JGzpEl98IFL
XGkHeSwDYtqRy7vtdOZSX46cfYIVxg6TjxDNa/gE7gtqmxqaGSxHNLszLVerOyLf
gPatydFpvOPI0R+qQyasnkc6G3w33qOBEFTqeEP0IJHrG49ut0LgMF+T5ADxI7Vf
nNXH0401unubkTSvI1EKUaOSz6xKkUkdmEmLHG/w0bKuq76cpw7H77WxMNvW9Xoh
xFPc9BzdB79oco+q16eAYpTYzglJQvT73Hf4VKhiUu68oROJaoPb0XHH0zJKLy3B
R8brR8KkX1Ztbm5hkteymaMKnzohvHSRtSAZRYMdMADuourF4/uzRGgN/JsLkvVE
7LTe2ZPaF7aHgiTrDJRuIBr/1d9+64z2HXJAOtdlWxhg8kW1dDDUVgjBKkD3d7aM
wDRAzB41EviESYfwGvWc6gtJ9CGangtcITvw8Igr+XcFC605qWY3ZMjP4M8vlEuj
Y9Lv4OY/5aRuEM8wosx9fSxAuofbc8yXtS2k4Zs8UQvkzSIYcbwdiOqslSbpW8p5
xTp/qqw5Kzksbm14AluD4x+LHRgZcf7FmbeCQm7f/uctvZ5cEnVUE30hfFxQsRlA
Xa+ds9LFBiTlLEX8cAo5LALnAbJPVwN/bON17gz2e77cG59yIrJRwkD6ZvsUuPwC
KeHMSOxY4Gf50mnwbYM4TmUAJ5JhIrXrXrCSq8rdwKZcPlf/A8ZP3E8482LXwfws
0TYJZ6pGlP1ki894N7VQdZ3LdlytzdkoQIt27HjcDnMeQI9Xpl0M9q2rifhCul18
Z+fgpAtCOH7HQ+Y4p9qtWXDccj6eCnpIfGygtmIZ7WkT6PXoPiGkrYI2O6d+uRTg
YfEdSu3RB27ERPz6fHtWbDNMPg2ZAbR0aXHhLTV1Dz94jcGk2jbkHw3JAMG0rYwi
eKTppSX+Sd+Et2zUY8Nh48u1pItI2YPZOMBFAdDpVWP+I8lP8mMHE203diVS8ies
/TOTgMq0+P7iAY5CHY8ekEfLeMUhyuUjxRb2MRlt8LdS4gCls4iIQHSZTc2j5Zvt
kZ4w7V9yMN3IP5FCrXtStJWEMTEMUNtxX0msN3PulbfJmgT1VhXywrDmL1vhsFTf
/n+mMDlDNZMRGbZHFTGOhXmPL8nkyyCI9FrUhF6UKcKASjrSSBSjdTO1DqSw/II9
n5LmaVy9FCjIom8L8+PEJLPyMplbwkLj82RiyqBQ7/IXvRnGsEu6zqZnzbYGJgM8
AgCcCtth6NH5wJsMw0LmBSbI1o5HE9fpfbf17Pz+hNPXAGfzQl6tVZMGvJfcNVMR
WXytInFJ8pVkJ/frYhzICNmAZXrYfIOzyY6WtTPhK7KWbc06ZOzjxClp9iFwH5dT
A4tB4JNjOidpCb2B/XjzVt3qOUFMaCz4fPe/OMpeDnDiNOJFHrv3mtaNLG4vfUgC
crIQAvncW3UTtuVp9oPGiLUuWw0JDuW8Kwf6TttnEwORfsxfR2ycSOLRgc4mUuWx
do1cZzqM7RqLLNT3I8Wgi5jVgHKj7RKtZ1ne1m8vQMdA8fZrEtE8jFdw5S77TmCd
0N11URYUvhAonwyJ59HuwVtXOZ5KF29LD7x8D5xXNd1hgx/9n7Q8+eBorcmnEj+s
CV1RNty+PgOxGllv2+Q40OaSdOjP6lBFMC8+hoZEfHmZpFwEFX03K6t4eCL/EyLH
5k944e8iyWs5Z2KVZF5iMRM899KYqTw94ezZKYWA8RnDoEnztvIqfydOll35WiJ4
gQUkMKdPGbK/ZkabP9LSgie7N+CvPQQCGcm+Cnp6NpLzIzV8IagLMc0E+fY2EzL4
Ff6Jty0AQhX2YiR1ddFttEHUPW/Cq0kx8pAQPR4vW4QbbIOqnP2LZavK3vQSy4MZ
SUjOONjv9+ZLn7/HnjgTfSIrKR2ReaZwZyCnHJ/VIdcxSaTQoznU52qvUPOhhKek
USiKBOftLG9VaJ9ZGPM6XpORUA2d0OGA4QWx3ycpyuXkzNCYYV46xOwqulfJcQRg
ZIccr+vgVsKBwYGES6egmEpjQgF2MViulVi77lSgVxElJelrD1ECs1ux5dAQNBOK
fBUnJMi9C89xogFuoZ+++8IxbwUMY+GLcAE0QDKcV++BEMmT2ENgA9cFmKsK3fLp
X0EKSjOnXc6NBjz4j/t7BR/40AvPYQ+JzpvT4dDHHXoMWIBDIuT4TRvICI1qWarH
7LXwUrV+sLW2vnlqn4i7obJ/ThocgDKC3lYizxMiiv4GsKcIM/xAxgpzECYxLIYw
mM90DJbmzRYBlmthf0ZIDgZIQMHTwiaITDET5WDwreKxUt2UjW7JhhKlEK2O4YDl
wE27/kawoUtPPSkc4yixmp/bfC8syb3iKy1xE7R+zMdFV9fSXyh1aLG6gmM6ADrw
5/yDyiVV/TyJHGP7S9GwDQYXSPLe3wjbz0KJX2hk2K8sSwp7Qpv/IcF8L0A0MAKq
WTxUuFqbD2CZnL33A55p6tWQl2302mhtf+0RXJKupxVeFdrw76nLQ7XMEF2DPSlx
X+f/VIhCOXYcBip99zosW914mHQQ7yges8+OnniLCMcOugqKB3dkY6F1zIvGonDW
rHBIj0hfWinWu/MmsjJsjUDT/RhdYetk0DL7dW44dVYTK1plsve4EtpN27bS9oP7
aLv6uPueHTxGXCDJCK9RWaBN1UO5Dd6DAg/x7EFj0V8HDBBLnRImoVLo8nEw0SGI
Uh0e981ofCik1lQOo6rQbXdZ62TPedqTmznnffQufnAiNAL5YpzJwhBWXrIm4ceF
MjgOccGviMYGq8XCbu5a+jEBXPJvGEfpsR1G8Ok60Xj9f+rrs9uipI4x1TfyW4B/
NDpFsuHfrt5jZ4l/6Gz+Ixrihv1fnQzGMDm7qgWlZ5czmIb1iTMMLOXxaYG2+/Xn
Sp5e+0llIZhehVxU9rfp9OApUpyu4UchwT3dnQJLhA84aJR15dfp8RCHrxIeymSj
q9Cv9zWIfTzTwwE6bK4vuy0jjhF8B1ZFDRMyGETrdGdwMjWEXHMCjcg0NgJkZ/uF
GajadUfemfcJC382HsqpJiTMZ6+ENZRRimnmpDNUhPy3nmrkG7WUJFrQNruQrylV
ymPealc/XbNWwCA5ZW+mP9JXt9HyPmH75sddtPl61ogEeSQmif3RWJt15H3+0pNT
Sqofdh/0De6CLGDPisvzGUWGy9U0xsnf1MM2mwfV6j3C18H6w1bq0wq7MUEwiery
0Kqhr46Yc2JcAYx9BicYm02V+iqKAQ+wnUxwkt/xjZ/wS/kQiDS7k2uSZsSCATcj
+c3xbpRRfkSVj+wmGQ8NpOTHdV3E2j6oU7K6iF36iW0jddzleFNIAh79Pj3umt3u
uZprBiOGZHxduKzHum3+zjvBmhj3Ph3Dxsz5k28dQLoErMgqHumKPwwINZ3DS/Yx
7l4BzOSdrAXxnCNqyNsvsrljaFElZHJm81JR5pp5Aqm3RR/ZqMvo3kfWd367uyoT
t2v3PuX8e0l6WFnw3Oshi4OfrbmjAkPpvj30JZEq9Av259hsqsFTZeQOsMsfIbaE
MwxvG8iCF+JpemK136Awe2vAV1roq5xfQw/LxRd8Hk1hQP595HdV7q7zbOL9cqOd
vtgYkTRgfH9sG0OLfHnRmuYmIJzanfjNwqzD8BAveY405fk4scqbQsKX+x9Jj9aI
iTHltLuMKaD3ryp3joULWdUoH2PzSLiFMCcmf/bgRAuaR1pLgstF/7XpxyFFKsyj
JWxRJqqVkvD3R/7KWvLlqsHroPguT5/NLnK1D1mUlmi1/uOLv1bDDI3oqKDdJvmH
jSetpmuXEUbVzw9Vtq6ut48ByG+Isgou8tgAnhIRE8kkxihvBWBve1Ib3SoTfeEx
wJJSlYoeqovkKQkG6Zpcypth2iT8s1YtgClBFc5IlYS1Fr+/OaD++oJgEAorxll2
76rwpuk0QkEOYmb+7M79KEcl7xOgmcE9z7qp5ruRAJwMpBHlUnZNpScCQLYfL5QT
pLBUsclMt6rLZzDXlMJdmYNWIzJfgj0PmWMt/SmBPeUK/hWdtd4xKT5uOFJ8K0wO
V2Js7GBGcKRW4yoHci/ymkZpBRAJVVRAt6rpCTP6JYrebjQg+2iGmjUpvKUrMqAy
UF+Zk/8NgnM51oZbJshyTv+SIGxTa1KMX1G2Wkf8t4Xws66i6fpZ9yYUOVdgXweL
c342UfXkd7+/YZnwBeCBegylzGK3r5IZjeYwjg/SnVGkBjRtcWrnsT89r8UtxLRP
vTuLLOQEc95Fl0BsCh6RpiMCHsmUTEAHZK4GAJC4eXJrrMiZgZc78l/Aq0+vEpi8
zKy6gsLb/WSHLZmYPKEyPQHqUzoKydriBtouiEWOctAQgZpAxmlm1wKadj7Yt51C
UyseSR07BUBXSBuTkG8KKn154eSlvrooPVEHYYw0k5E48tYEUZZlG8uNU55WaN2T
MLBCO0TZEprsMjU+I0+kjL3rGEWk5SzZhv8KLnudrN797DcAQe6pEldeCmllF4XZ
2UES5qPdgTgN0V7oI7sQBYCQzKR/mcpkJUggx0T8hRBbj3XTrOXISi/VZeETTAj0
BeI7wf2VZPA4Y8wJjwYHYckflfHBDhlomMGocOftNQD8WXzNo2fuGQFEI2Wg9Z3r
Y0bQYPTKBgAxY19A2D9nfSlS3OMV4nO5ciS5R4DtNlKhCbUY8tZ5JzfzyxipcENI
jOTg5Egk01p689uY0riVoK+3vFyiI6plPG6hnr0tL448TdW7VM4mFhKA7mW0/kaR
wUR8Tkj1mAslJ1LK0XR9WMi/t/jj7HfVcccDUnAIqYk3Bg3zIlXNAc0cIB33s7Uc
SoUTqGpls6+sF7npue9xZbgNYoNc+Bhi5AcdJEKlHGFgeXspHpr0XEGHS2KGzTSY
wtxLwCGRw6WymcOG3Rc9uiK/MoaFV/lHtv7/hPn4N4kHdS8zHaVYZtlsutpR9XRM
Jkd97MKPYoCX5BFu+jLMFaQqHSlV445YzEcN5wyuGkEXh0bCaaYOIXm+b0B9xY9z
er8OkaJoq2awFwAhkAj/0A37mQOohxvOitBkO8phmPTjkZ6qHtEUNt+oxHdB6s7V
+n8Xjg+U53B6f4R2CmGpGAL8+XSQTCXF1kHz5z4j+4glG55d5JR/CIUk9e7RybIj
FSpL5An1fU0v2Y/Aqv1muZ55dHR0yUeWkqWHUcXOMHHd95APA2amRWiUNiyzeUut
/iBw/iAZcs7o8MU7HHLrYvX60iP+dSr5ZPGoBuftRt9FnbrmthOxHi5lhNkdgrY/
UBL5+MYe9edLNyoiID87ezTWxuU1wFJB3kkZ52tnuDUjwUyqybRwUDjtQw2xjuZa
2TROlyfBcP3r+rMazFGzjJ8ytlFDQlF2y2Y5l8ixHbNUiAhStsD393yXJ/Gm6NKS
Cg79/Z8D/a0PvOZ5f7Ps1g2ZZFxO/8RHBD7CawRZxcX4k7EkCZWstQ1T+H88Sxyk
LcNdiqJDkXFmwphDJbx14RbRfP8WZXt/JDGP8UXZ42CuNS9DxvNH3eupTsyKnyny
QElM9+wKk1ngwK+dDx0N3A2xZs6k7SvAtnc0V6WTniGdfXoscFU7g1Y/KEz2kN1V
joceDlBoNjuKj+cUpQU8UB20g1liQ18NJko/ep0TLh+xHJAAjD+rv3q+3PN2v6z1
oSYObZqKvjwMIQLpv2tic9lAgXnSPelQmP7aimmUrWOSf0Vu/jHIlXepKdfpw3d0
ksc3gNNe6QWBKHOvDzQAZUEP6HZTnKrfr4lG8zWAyROmoLfdkXuuGVD73Uq5Lhhs
V48B+L+yLAgeC1H63g6TKGlvjA8h8Ml2RBHJwVJXA5FIRraq1nbeqfW5mLd1/cJC
Oj1SE6LJGoUB5gForOS6sURPZWH2YX4Uec3Vs/HYBzPaujqjMf3BqwxcfJlroUNu
hhxl/MUOYmUUsuOn46nh25yEBS48GdpiwPFuAh3xQfTnRcW/rRJboLA3Ziw2iBT9
4QI+4Z2684cJRFSW4OTgnmvrZFRasRlOy4SYdq1mh6E83bvyRPa8Vtsp9LD0Adth
RU5A/GWpW1GkOdJL+51k0Cnnr2ICXKO3R0eTxzAOck3tJlJcuiRgfGlTJLqpA3GO
kpwxnKdD7jTWewSlTvFg1TG+NiIW4TvALNqFH0ZJvDJBWSPLxsWzUZkenqumOaNH
UMY2iykMgoywUQtgNcaAvL/WfO2nVBtl3iAoEGskuHXKCyowc+xRynCQ/P4/BYwo
KNTM+uNdBS6PORUd5SuccfhOj0bGPPiGvb5THsAo6ryYDB6eRWk2/tOmuXdY5KaJ
Etd2o+ty1a/7cCFZ7qFFaOodSwXM6HYoKgFJxCPivsvxWeLT3z2xWlHTUKNSsuva
0UvcZaz3Ey42w1zsze/dYm3Qd9yuislZYOryNCD7pOyG5bdfuraaPzWq89yQD2Mv
770W+SSw4ic8yBV0J31tobJSNYBTYJ63d4bzkmbsY3Xzs/axSnM0wGqZ1xO7Y034
nL1Sp1oRLd7pjiw1aq1UaQBzXsHaskJFxLRWCZFP2cERCiM5carIjyPlGSj159JE
6z8waLn77Sjj2KAHRcfmt/DnwZnF5USRD1onkvTYQwNtliBYiy6oCEXIaasBBHcz
Vu98j5TKsig7OvdDQX5rL9xcgLenhwHH2cDJtB2qE2UU2fKth+KAUI9NVg3gTmWk
3NtKZ13GQs9Sz2Bi+RPXufp/XW8O3q6FWUVoBcIefDS5mzJ97/n8D5EcsGkEaFdi
BalfB/KURzfocMBMKFvrWd+yEe0NGQJAB/aA4reQELiaccQXlGYX38WvlwOQXCX1
i8nFPOa9lVDs3zLVuXFGvoDWfX5BRWtLCS6KA7zoKMPFvF338rQfy8aSU529vQqG
vmMLfu/ETs3oBQ6pFfjpT0JYnkBg0z6bqXsfZTZmVJNN0r2Id62V67DwffMsWL89
OPBDPnZyyOHa2jfxW6j1DXgq9yV15a9okMYnE29e8yJTanF3CJuCLXJI5nrO1glt
udnWU5ox/aTJHQwpTMXjbWLCqD2Wj+WLjXRtZh7w37ZAA1pvuJbnSacnGiCQWLcE
EgbJRh0eIl9DuaJ3NIUa6r+P/vgVm7Q1KI8LJSZrYecKiwm0V/hKQLNJjh/tj1gl
ZCnxLrzlirYrINlNQTtTvYGzL6ITankrQapvQipJO/ATsSeG4BXmxsh24miQAlVu
0Q4Vfv66vONIfb+6WRg4SQ73klS/FDX6lXTJCLEORcglFHFWN1j38apKXkUe7FxP
ubTpNelj4ADGzyekNHBJquZfuNXEqA6X+AzY8sWvUEf6zuyXYAHe4kuPVxZITyNX
+ZtxI1dvu6IuHGgffIlDhZjIOHhpHIIvn98CEw/gkgDfyQzNLyEfcZzF0+ghEWi8
/FoDyAfYdO/GcSGK61PtO4flbnfyv8nWrRMaw0pWVN9tW3Xl9ufjqfCnroiutH0W
2PqkEPCuTEqx5+L9r9KbH3mAwLOgxJJYy+EQsXwBghIjpGVXSUfRDQK/UwT7J6bu
zx5GZe+FlJ2y67QCzVt59N83rLvN9zOp5TCtajXsZPBvI18lCHPrA+G+D/2PoMvK
/EOg196j6jLKTxT7oLzqoVXKgIbaNnD1RIqLuFgIRpqhLLSS06h80GfXjZ8sDI1r
jd9ENZGxWnsDr04sb4nzL82JtC7iSDoZ6Tpo/tnbELoQbUxVGc3NuztXmLV5zt+Q
RdEriAg/hSCOzI0hB0Dypjgc20MMhE40k0EnNSYQEHBSthaXMK0dcIxjbeK3cGlP
Kl14h0cFD05yHosG/vJ6YDWAqYxZvQql0akp9ZezMVrjUB4Z2bBV7+JYdBgSJNv8
bAKsxF1F79Fp/30tjksrcwTgFxZ15yfie7yZPvRjzEEP131DxqfaJTU0x78CkFHk
WEfYg2sjzlMhGMfFjwENubpOUITPcr3eOkbIzWfJP5A6FTDQuPzdzYCfLiGtC3C5
e3RCkwTujGiFWf8oud9cQs63pUlPfH/UGosmsAqdr+k+PbLF+OmRTOkOa3ttLYeI
ryHWWbNfHp3/njHCK6vLt5dAchm3Z2ybhhnKGW0bO6rPmfhrqtYoYPU8Va4OmCrH
blbrmWj7DoQOKqL6drYugWQr9YRcQIhzOo6H1Tq2f73/oY4gv0I64yIeiO1i4G72
PYuCT5Z6tziCtjwHgkLQEvIN9Y6n18XH9WhmY3dU34HtPOKDuxf6DJbAZd1Lx0hf
Ugh/oHDCKLSUrrUDJTOAGNZB/Z/FD7iXxuGSRa+wMlqeIaHOrh49NFLK06f2M6VE
/MryT4Rj8uJzVSIBrb0ZpnJnCBVv6z2j0aRLQlisjq5VGz1iP4t9XBbET6gyFw+j
R6TS1y2lFiB4TqU01IuvrDIMeAjPgFtm19J7fCDUVhmSwqZ98l/IpwlMxFfzgHL8
yQJt0ctCoRRP+ZRafZEf3i0buwalv2e0CBItHjxIkBifmGGWgUns4hJYBRd/v1J/
j3MS/Li/moDSUNHW/V4lLvmrRTsXpA4VxfcNH+Ivu6jG51t8zEfqgtBssyX1q9ci
JF05cZmwnPIjXSeDWBww5uqLlL3FlXruiEm50Mgr3FFu9gK3F+bazFsuTh+i7a4L
/VrZsNVa5ErC6U3Ny82IPIwnFmllut1uFZUve5kVyRLTr8EI3URDj1XpwzQi5b2N
Fbtg9ktR1LOkaNVB0j/6Ie/xSlgy2G4PPo3xNOkA4fPJyFXGmpeF8WeMj9Nu1vET
Ee9591wXtItTp5QVka37EJa1R2Avyp6i+Br82SB0/AZIXfxzq5zA3/CnnXD1FzEe
uebrk8MLoQ+50eLNZWlnePujJoZucNDbOiuUhPWkQVfT2l3DMg5khXOS0v5KoucN
mScayLAn5U3Yn2bFrtr40XzEWt4izy19huZWPFXeSRdB98zRJ0r3odssnIhabbKg
Yj6JAUs8nOVNWoSFgvkUvvPOloPAceJ5VjnSu2FM4f3u0VMOoDAUpq/HRta/p+LM
b2wGkYAzWDwbnBCnuyFOLpq/yagF8L3KKL3qe+kSruY1ttR+O3kAhNdXiQQa14SB
kLDeF7os3KB0b2VxoIupc9Jpd0uZfZmYNdy4+1L/txmqedX0nwEQjyALjb+6YZYR
ZXTRIJ3qXJaEph6JIXfv2+R/rop9HFERt3acIK1I+SkgYI7fHKaOnZYsrpI35QPB
gOec/Nl98LmeSGcB+cG9EwcHpzl/vildL6GqpxKPSJVSgkAe/iVjtxKalaVWr4tx
8Y+9GNNzdOHDf7LVBulfE8wDf1hVtBeP2ENwhdWIgvTW+bCTmpJmnvqhfb+g7sZq
e7pE0WAFsYQy6WCXLsoClTfhc22bs+bzBmglXFheRWOqxKv/dEYVcbtOn1N163bF
bFkVkPYKpVQRI5PbgYETsc9VFIXwNYIASqpNrn1zNB8qE8azLT4wL55dK1zZPTmk
/rnhR2cP//5E00KC1lejcY3Y4t6K3RP/ZRwR/b7h14x/qg52IwyeHrLbJ6nhCZfO
7cFR9PPJPY1z2Xf5B0Dg2kckNO2nR9z1PWpMXocXnDo72VUmK53wYYPQf3IyfCYd
V3BOEA6PX9kXrjBgWUfoq5w8jmBuJZghT1sWtxXuFWLi4IDTJ1KhRxR6xdKM+SR/
h6gdPqIPCe9pr6PhkBKi8aba+0cQkvV8Mz9xg85kADp0+4KmFh8TUdxZALF3x9jU
yedF83OZ/Vt79CU4p54Xk1/ch4GXuql8WskK5OeNyCni7mqEtbtplLsm0H/eahiu
Z8nyXX6luxaoDCaU0/sti7Yjz0Dp7pYxNLRfwJVwcwTyzA8sI7t0yc9qBJwbhNB2
/k1vjkMj78HHemQ6IJiQ5d5HaQhnOq7H0S33V9xHpdRpoMtVu/dNz2MDlG8lYn5B
+jRktuhzCg5PoRKrq3vpTsADLWyEKWFxsm5UmFppsyBkGfuvhr3zwHOf2cqOCi20
LmDbuS+K/pHYLtmdQNr8xVqtGPacQp47BG5t6iPuIw1MDfHJAP9nkkuH/dyZc5vJ
nSG4FsfzruIi4PhvSQFAEcamC6IsIXTvGzdDYfpLPrjd+br5tWO8xfglgJYGz3xy
tZ5EltzzSCZwb56EEfihR6FBVglZUvlx4nbc3pNatQ1+VEJettOWdPpwxoPmmT5m
YWpDSPDJw5yDbsnhW+geGB+CfrvL0NDSYkFhUojnKpxNGOrR1f8MrazXzTD54Ta7
gRn1ObqKdaMH6/N3x9+OteDdN6mYaetUSLha5VuPAwZg1FVqIHB6mxlUvy1yCQiJ
xtoRoYTs65IDGG/JOs74nkFfZKaUTZ1KoOYwDD+Awf240BExQb+n38IfBgtOSggr
y59e5+0SoYoiYNHl44mefjRQTFUmV27vmJhfjjU3VtDEfwIgNB99UUkPpgLT3vzf
6qqHPfc+pH3I2tOaS8O6yLSS176cn74SPFAve5tHpIOYiZD1crNZnpeslXUR9QJz
lvNcmj+Nd4j746Gp79l3Lty/PvbY05AhbWWVU3YcpBBe6FVQY8lkeQwOxUezgiyf
YtDgb/auvGLG6768zChUcq5S+Yeng7cRyhC0+S5AHQy9CjyRfP2O+GXBUFgMwOQS
/7JImQXFsNVIZD8SJBKAw3Dyds4JyATrB3tgC84zlHGE6Zkhop0bRnvC8VGDjqEV
8TKWTs8sFOenPYXYXvahhd3pns/t3UNF2Q1ZP/pDvMceQZKAeIMMUNFMCs2ebgwj
melGnc93mUlD2Zwy4CB/4RzIg7wW9gi3Zx4XgJBJyDS57fsM0yKusrCKfl1LJAGT
9/50tXZRH9I0wr9IHTZsiaIAmtoz6+9rsIh97uCPagW+PNdGDJcnad8/6A1AAkNu
vSyua5fhf0VkDCq6jrYJ9tE32JfGtRVvINkm6eL1O46Lp639T0wgPnp27RkfsVw4
B2/lBgOm+q/Qn6e4hqOAXSLpOZ1a/rIOqm1eypt7/7corH8kagRmSc0Yr9ftFOdq
69Fvnp/qH4Qu38wrW6tzQiyddiD64E/UTtaEG3cqU9MzM9lAXSKIbxGlWT2dZLNT
y3/GsOCcFH8J+H2YQ5AEHt+i4tcZhGwItFsToKM4fPLodXOdkco3QLdYU32fIlyo
o/S2cHb3FkiFqiQcKtYqIP61GCrIZPF9nkPLsaRqgV74GaXw4VyZgR+WD5lSHiHn
F2Z8AQbaOLFzTcK7w3Gxg9heea8vArgfnX7e1ZuTvChpBDQxLzrLPKq/1Spwbtkw
Mb2J0hw2sAMmipaQXzD+NZfTUEepstdHEdd8Xfd0KJi+0U4/Od/zBvHNOcPI1ynw
Uyv/NocIeIeznWxqvipiLFesSM4hleW4yjET+pEAZZFXoWeHwfow7hNdPUja6cU9
RG+3Kd9/89+x+nL/sItY00Ap5vvpKgG6dlC9knETZJdyMLA4rwh49+E20hsd8cw1
20n8ij+Y2439T1auq/01LBQ9vPxDAy475YK58BhT8+eKRX2Z30DHQkCX8mGHd940
K9uAhAzx4enL7TKTMu8ShrrocmBJmYsnUIOSYJH5fwv62cNo1neVpy5FvGzd5O8l
eEO+mNYnRQSj2CR9FbMaRucP1bZlQyoWthGR4mayPxTpdCMnAW0fK+7S0w6LosdR
RryLhyJ9G0Va6lMsXiWESIxKLy+IrlWtUAT6RNQ+fiY6bYS/h4AS1+kERzykgn/c
1IOrIzhkbe8Np6ictqd/s6wW2lBhMCbOa8+fxrC3WSu821rF62+j9tOE7pVmuTrL
hybM2cGIb/HDqI559CjTJEcONCm98s0NsCNwXMTq562PYrRpaU2C4UiRfNhU6QQv
Vat87Oa3WD9t606PyiGyN1W55tuEanH5VFO1FEJVVh5MTitjX4fmR6CtaX+0q679
qcu6kpFa5iI2WV9tISIO8vzZjKqk6FEoHfMOxTMlAuZKmMQqk5OUrvtbKgs3xIeG
Q8ItA2eWv5NjTYfAOG808sDJhMaS4WN1AkNt5TLdqgPCPLlRmE865uoQADBnZyiQ
OK58NZniF/plgH7qzzAbVlBzqTAFJp3zbKvwkKYoIkJoxQ3VEIM3atAgDyBfo4vd
zRAWfHqs8yDw++/V5e8O06DKTwz+wfopMhjaYbki4lZB+bzdwlhIbMPyLXZA3s5q
Dt0XrQ0RIm2J39FjKbvQU3Zykmqkbyd32uE7SxkdMxRgz16Trk4KovAjjqFjIQ5E
POHo0l5jnhqgE2FfeCNWUZGhIHyVLGe7qMC3qRVPBaTd2WlyO+QyJK4ctK80nW8t
hO6medcud5Lg0pT1xRvU+ufSNpy0BxpNODdQST3fhAnjm9SvS1X8zV5bOFr9/mKR
5a6KbIVZwst17qvVBNILtEx8wfUot8gsShtHwidBXDkf9Gvfjqp3P+KPJpdOj8Wf
+cWBGBfWoP+L+v081mrVwO+v4ICDB2uFwOMYobZIhqaz6tgwP3gn0zcGr/qLl4wH
7AQteqLM3rY7UhbeeC4AV412U0CvN+EbZeGbQaLuTthqfQMdLxtf4duFjNB7Pk1o
odpSwVlai9XmPmudH8B5U6aSGe8pQyz1fLVdDfTCGmlVZraXWdXysfAZypZIkm8a
fDDL7mcEeou6k4SiaWJf8jnAloiz8reV5kwyqR+s5LPEJIEkRmfzu2JX9GMjpSeY
AnhRLeS4jFdKWLNnKuRjrTEhlJIwsrz9NqX6TmDDoNVzgJ/GTfC5FtIFcmGh9Fmp
6dETq++9gVY03qu2EE1kbMY6zxsUujCKv/znp/5D0sX8VUtMd/Dcc9tg+PiQpWxk
HPfTbaHYqcsvhaP12dobplx+wM4Nb9THCoGZUclIRKRIMeYXanCw5q53OJZW0cHI
nY6A0VRY7DfsMn7vXBtIP30i0t4ideSFN/smeOU3KgTpZK9a3tywgJPXDF5USKNA
DN/RL6PIOF1GVe5Kqn8oR7qHn/CCbfM9pwZC/HyciKKvwuTNG8Rb9euISulOPVCo
79MpCfmCFpQ7tRaVoI8S3a9NcR3Fozq1kgoD7+h7oz9Un+TTMV5EMZDpXCW3Irwo
D6qWc/K8ke+wHqojtH7HISg1hSBQsBfFzXluJq2vozFuOIdL72fS1XqNhhLzdMCv
HZ+TLAcYn5umXbFUBacZAS8tT6nGvytfTeZxFlVxo3MXQvQRAhOL3OrktS11bs2r
Ka5+3NZALxIP/D/l8wdlwTGOkNL6e7O0p89lR5m0Pavwq66iPRbzp4G02eGf5SpU
j8SEmCFxn3Z4gcFL3UsYpd5ilXf9EnWuqdDr0SGpenkfxGtPNW9Fl+px3/DplG+X
rnz9RckR/9croZ5nM1GgrE0AdAr2Bfy4yJqIIYFCBueAgvK3G9FWUT2pyAY+0evQ
56Vmf72qIeEd3RqHcOTungNbk+mAVsNiuQkC24J3c6m8evxPDSE3/IzCxQH7JlQh
8sCrqMpoqomMB90MagANy8omGYFjcdJ3/TB+ahdd/dBy6zStfuyYyoAddYmc2MMt
OiiVRr8as2lYJRdAYuToyTDqA4/6OwHPjlJehQrcBbHLfdbYHMyraiobN7N/DSOQ
v7hoJSP83pJFtbNrw4BGaccQaESrIMIX9V12xOedURG6wKl53fKT4DDB4+SMqK1F
6d3wB/mJmXPIxbAYxAnK5tFFxC/I/nQPo0Fw7IlSGq3PhD9jxWJLJ4E5h1QiD8/t
bdobazrIDJPGAvcZjE1w/wMdR6EY3VDMPjcUTWSLJzAO2dvxTlpXapQeb1Rpdsg7
Tte7MMvh9zum9tkmQcnNs1YyTKJSzDc8mbsrJp6eJOupDCRdh+RveEAdbo8hoWVA
cwel9s5j+Kmg1di+qCFGEgeRExd9WFDWBzAlQb5oLBezAzC1yi0Ms8Ab4BqjeT+Y
XRDQWMiWqiSLVRdVYdbTgZSxXLLlPUOnTq3E8Ngb27xIIVD3CMRiN3Ono1M6IyPg
UKlewTAycvTqb/1iWjjWXtjjVggYnnMxo7SjLXZXIQuL1ua2xisoF6O+8fvVLfco
RmpsAwdtqWN3WaJHnxLhD2clvmPATGmnf038Aa5HD84UN1P3MrUoUc4YgqK/ylBH
wU988LS6rCciT0S67NJgAGrubjLrZR43od/TCE32bKN5OoPcuBQ2zDeZQ7l7Ryx9
nv2cVfhri86BbhYoz1UPuyPSScnHuz8mc0pTcSf6QxJGNeobFtQ+tBH2Or3F8FvA
jAMRYVIyGosfRuGmHc2Dsl3oKSPbr8HmpfevrSjsKv0yS5HbUhGQ6KlUToUMWed9
v2BtZT2rsEqD5Li51O2QI52igF0XpOr0SRmDA2BApHDV8heB3NExOZlhknKpjB9F
aVcsRg/UZx8kaLdi7fEMGd9X8bng/RsQp1xoym2lTdwcIQJ5u5v6oA97Y+dfEvk8
G3gmAvlAmtmj8ARxmbwN0iNnaO6l4dCSuxIT70F/5Wd92nVGjs4Vt5p/1HrxxC3C
qicY5mFf44BLmwQo/pJ8llyh/BLUM3fXtK+mKlFgGqCHAKRY4DslydEjwa43XBYZ
IzoIFZ5QmlR8b0GcVYdlRxbW4bx5k6nGwPnxSZc+Ru961ywqmr4TL0u02jk6QnWS
0tHxM9Mb91XTNRLVUWXEUtsxvMfCdVmsrTAOTck9HzY9xFBZrZfYfA5ysjdIs+Ad
7wRfigd5RhJyJeqjzCts3suLTdD3m15OSeYY4E1EmqxsEo1NWqWBg/4KhdAaXAuy
I0iEqK7ksidOeBGmE9T2n49kwj6Rps/fOEwcNGrZgpg7cVDvpK6AiRrWauVVcKGn
RnT4eJeNiA1raj4WGL5i3MNq5uWge4X0pt6P4/LkQ1nRu53Vt7zgb0akAqT9XfHF
EDXo3lfKiPWOWg3LSRGIg6a/Lq1Ybp4kvVRtaRWIbUH5X5A01LfWFLTz/SUb6XUq
69xkGtlvOrJmn3zio/oUY4+QE4WZiBGSzGrZiySLbzO0LVJ18hK7WmaDtcOnJDxh
7cNt+crWQw3f2qjRN01A9UsEclisW6WjKVQOXWCKJSwSERSvGRrWv61X9je2uXqw
fBsHMFb+3V2WOvXBXz4G+WbWo3hBNzfySAsAZdvYmaDUJVJgYS3w2y8Ippolt/Z4
VML4oqQwlHWKs48OOP65y+GyqJhsc6gG/uQt6lt95uQXcn0YnWrNZDTZAFcvpxvI
YIKQpCPfgiQg1YC7tll7PsqZFQjUdj8Ib1ekDzoN3cjxRuLazYLDiI9DsNN1DKKe
D20wqpcIwWqqw9/805pIZ+CKB9LxePbrN1MWYWQSDiSiKuIiqAKruQVTeNMxtD0V
1zDpjynPGtog0AjgCL7aAVHGa0P+8duIjwI8204NqO5Cn/Ze/in0xNr6pBtGdWcq
AkYUbAHOGb2asplJub16kXe+eXDVrYAZXnrq6INm5sxeZPe+lUuBxl8i6kcLFlxq
NITxyTUptO+xLbJDUW6EdE0AER+NkilBfCZgR3HW/z10SgKig3vWtDVvcNTTo8w4
M+OxVwBVWJ+uEGZ4YqUV1X6h3CToR142BRp5dZ5azkKLAkELM9t4X5YvWNa12Auq
NNLklHc8sm2qJOBbKNQNdXX1NFdffA07b1GLlB1vQZy2+mU90DAbbJyyiqvEArxS
kkhQFjb8OnwB0xOLfLK0qhGkR7/bB7+YsuCy1XGc/kYGPBfGzxSIWOZ1GJ5dNZ38
EscmpmCTe5EuyCuIuqNKAm0dDBBF0r7dL0PVWxLvy/OX60YOQSgBJofMYnrEP9IE
KC9qBYYy6NvwnjAg+EkqB7exbbXq96lMLZJf8RDqhNoJg3K6sSBdTRMu/5quVroH
tUyRUktibbC6gV6orn1ayk/8XAi1XWwoxP80v5pSQsmGoKDWmvpewQtEBLceiu1a
AfdrAqpOk+WnqVQ3IXIwWIuNIQ7piK0l3rt4PiV2IEto8AXqJHcoOznEIkx17Sum
UkUGksIWImx0Uq7amUnEyh5ujkQYsScBRuTZ6E7vVDPnGrJsUFaK5WlsnZ0IEYQt
aFElvlEwXOcMezRaS36iUfvyWvQ791Tlv6DGIbLBOsWgkSYcT1tp3ez8gLKlFa/6
zQLapBx8vWNzZKq192lI3Au+6IUqulPytDKX7jWMJhjcZkb1m7u6ZL1uHwnLCnkc
/5ZJJYTUoTO3cGhiOCOHFdrqBzlmqcGZIblxpv/U6/XEGfsInSzzfKoWDsWyZZfo
eisKnAkNr41e1EqIfYKZr2P+Vf+RzC7JY9WBKELF936NGh7tMFA3dg5U9j+MGku4
DEWSrxwLeY50/7l4bP/pCjEEnCdd70V9pfQfvih2E1oDwlCeis+/Lp/MyZ4OAuI7
I+cBOgiRBRI5pILqI36Dzr4DH0Miws6V8nOAYWYw8k0+iC+QJBcB57el+fvhVDXa
FNVkpQbVI3NM/+ORBmAXdszVHZ5rQblCiJiARs1domggPtXHaVFWgNzno/mZ5vDz
ElYFr0xcA0js7KvpU2KYKPoCsiMtFl4agHIbeXEfC6o2md8zmWaxjbUbIutGul5l
lVeZo6iwTpqq9zJXcLSrrb3xbZ9F7U120fc4ZZuCVPdqBrWvqA4NxdgqYA06k2bb
MteOoGp4w4kh656vsjm92bqtuwJ0Lqwt7e0u7e6xTuMVuiQZEHxByEi9rvGGeP+O
cQTXnbGvIpTn3h/pYCYCAbRAxCP8hxufhv4qYF2dmcdgvP4ICTZWHJCTeunj+CB5
fUeoZrg3H40L59ec8F+64U9S1QLOSfSNU0M1WXec3p4cjQzfCx7OLMY+TYyUDhR3
lnxQecdupP7JXmynZzRfOWNC1lKeA58I43eD2vPWmfVhb8RiplgyG/kSLUR4pgFw
b7GRCIMZa24RLIshBxUovIhf0JFgcwl+oREK6shbgRDStPMGwnCdy/CGbMk0dH0m
9/5uzXDuGsYejxhNCCd6AeQAvzlQhrNfyXmWoEf+SNFpoIG8+svP0HAcUdL9528G
8kkq+oiup0v+j06FgwXLVL2hjyxR5cwlusWReGYa9InLKFeAWPwpBcFXEEJHDr20
rxx2U7zpMl+oncCcLtK12SXqjQJKxXR+0g2OBdyAIyhiO32z6XdihKbsaMY93/UT
sTmGEPDDSVBTtzzZSqZr8wCJbns8tXtG9+Zbkn7CBy30NbezbYMBTmgJ9JxcJVR1
POv6oOpLRhd2KR+pzTI0GnLm7wmJIdNoL1TedtMKvF+UP83CK/QOoKWYI4U83Eb/
NopbqIu+qW/yCTKt3cVtOOl1pzq/YYyDaqsjaJf4j4hGwAZzCOZCqoNIjQlkrHCO
qNL6Z1ByJWZgNUmKt0g4FK34lOPgkGx0wa6vuQkYdegYVYBOaY0+MdlO6FCORxkj
jeobE89GwTNXE4ekDOShNzTzE7EGSXGUsKkI9+JrX0/d+MbpB5v4dNnsSkTEG9MA
W5vP8pOrFjU7Awq8+u0+1M7up5LVNZoX1iZWjcnXI4Dx/l8vFaBrW3cDvsZyqqz7
su37EhcsZqJinJuOIgeni78pKL9DXRUnpKXnbCzZe5HyR+OEy9cvkMkhp0f4Yyla
m+c61Zkwa5MVmo8rTQ0kWs3BlDnEtD/gKDTGkSHBhf9QUB9vlFmgc1p/nT/QoJ6/
N5m7GIUrHUK0oS3BixKZZifOC45DviBLyB5DpXEJ3OU7VwHkzM7IFyQhi4LFfkkc
7yqwrs1n1odmaiMbLlQuzDBFBbErYlXjtRpLj6weQLy6zwoyDisrawCsD9B7KBOg
SFppchArX0Yo1T6M4XIST670yreq7YvJE7OnBKHBkSs+Xl5LYIUIdS7roeutrgkf
O5pjJyvMXZ1B3n2XyubQ6Qz2m3RpC+CCwj8UiWOWVFSOC11kw4WPN9NUo7cbZNTI
Wfqjt6EtNTvl/iPTBfDIae91bkjWxDKaYqPvtihSwnnebgRlULmsrf+0Fu5XOl2l
odkACUkZp0DL7ULRx9fRPYvkadRPeeK//pitLVHGhoJip3B2HgrvVNGKJG3FonHb
r9smlgxGbSXCuTcniXzSfdZZ6shzljGhO4nbgPM4kq77Lp+qgXauJ4AFhBq10Dc3
Hz8JhhSjfsF41dFPkpsHbPfP1IeHqTZOs0osWWezR4IBlVrVQb1U3N6H989yHNzv
a4sRbMEi7yIR8n6SEAvGLDN1/6RWAaG3rgHF87xd56zlAlSazZr7Q3kmuKcvoD2M
S3k/apN69V6oetFNC2340bLRbb4ojQpHkk7Phca/a1UETmUtDyICEE5EItHSXHb9
bz2e+ItREeMapr+em/2mltkl/nvi3VHb1LxWjZQIWLCQhcxRYd8pwBZW63en9Or0
T7pvdPvH5ajzESkgKIJzs6HXl9wiL67rFnletN0fBKszzOElyUQTzbayYNRcpvb8
9nliqXvoJCHsQ1IkjaxMty8/SjBr7wXOiK0u12y3thKj3LJ2wGJSbK0lbnVPPyr6
snUMSnYPZWt7QM9E9Z6b28hCFB5dxWWvEMf4YMDnQu40mgW5cVCat9RdBEWixRK2
Rg1UevnzcOx4bDAn/Hvd0aWE0yC/wVf3Opb4y6Eccq2DvKRLeeCx57sRajszbJfK
G3/LBeE6yK0cbNIyEArbBeSeGtGBr1MnsOM6reJiTOUEuc/l6YIhixDcf02QEHwV
AxqbZn74VhRJbahRWyIX5QdOAiIVRucqlS+rItu3heLISMgr2zFfUgNAuVdC/frx
77ldwVgF1H/Pi2vaKNyh5dFafSdVV9PNsKJByzE873G73o5O0FHFYD+DZxZIQrQD
pZNeuETls2YxtyeLeZ9/gJpXUvhmJdDOJDh5099F4JURM1lIRqe4wj5V/an6w3dM
TObiVlGq2Mcv8wWC00+zxNV7CslGftAgAm38B1M9JtAjEKGRPvoRw1scL19gqmbT
MY/3hGpngbH9e9qkhbWiTFVMi19+i64w8/Cv1ycnRhhZh6LeFdLY7jlHbCZ6J6R4
yXrfNEeQSXB7QgOt8DCN4fmm/91HO/w3FIS4ALEi8PNrJw64PI/bu9Gt3R9xY+3Z
+u1Vtdoga6CtafZL9qkE4UEh6ACv1NBFU6pfi3OFXprT40QjOdB6QKJyJ2+wtbxu
9aGxEzkOJIje46nIP0CuzEneewGd+yzM94PexaPlzRhQVnnGocjSiW49JreZIdVf
AMShdUSZKN3Pz5+z7gD2TLluysGSNs71GKoxWy0cz3IbNqrePuq/XWyhmN+QvzWS
X3vXRPA8dt9ZumksqsFMrjnoQHapSajoDy8wa76xHYUfhbcjldpwJ7EMMT7vP66R
8cFVDBac7cfWxb4XjhPUfL6oGetEuYCsMy78KTIB2J7iXGbCbjkpMoxeTHLdR49t
dpC9xLvfNncS70NNTSYTIFTZqA6umym0HjVUSD52Dfwm5LVk6SlRzBi/QHFkHJoh
I13qWKKMEuDjYTrT0umkR2kEP65dPkDHrFeUt+HEqlPtXprmuF5OFFNTFTxhlh1z
+yx8F2LIbARlZ66ijC7y6G7ZDg3eS/TMG4FEwcOGsfRSa2DKDmmU5rjd8Pbflu9n
NwlLnrsa8v0jRHcQ5kEF5+bfBwN2dxFbNictFBvtwpPgcBxpMKZj7MQcmVRvI+6t
FpgOIQdz3Ir5EhhLJ775crU2W3tMaaZe8FImKdg553RzvDjGSWRPkNN1urDRTn23
80hfxLQ8sc3suwk6LV8CLGSihiAGlMonTy5te0QdJMohGqOkrRQP6teA0qa/pfre
BU2IrJGAkPXHAqxnNjA9QIaz1/v9DfLpFWJsr0OArihWysvt0cEhi7vq9EY/IBB7
d2DMZFGMEVe6RTepzDngTtqaMYH8yK1SVyJWGnKvbcNwPKBeUVzMDCa+7zTsTwiN
iNMUA5nTkjm+16PqT64qcD8FUd4ToL/GX1mHdGk3sx1gEOPO9od1UTYM2fLUHPzW
kisN4KC73+siSSIsi2VqKgiBg3QqDxW08tP0BsJ/ztz6+WdQINT5/+aIXyxd+oXG
aopfV8vjlz4Ri1OgSLCthQhD+3l3nBnCks2m8gc7Ajp7RS9jKNNMKmuVNdzfpc6p
VEYE6jeY1YuIUBXCMabS1e2Y6VGTOMqxikx0IPoo56b3u+UhEtVUHnFC/TQgdRAr
hBKO5SQUbr/0yrWdv78ExLQJeQrjy14m6/I5m3QIl1sIE8TXwVzkMjoSaxHInH2e
ZAnicIq6RJw8Cdi9jDz/0i1QpA4qiBkO+s6jZXJoIgDDT+IS9J3JKjUlqyAKC5ij
3UX5f4izdLHL3hQg039tRsEEcpnA1LlgGdbjiXyepkHx0b+l83NGa5rbxifvcRup
Ue9vSurL2PVclCTOAAfUfW3/LBeaI9DrTpP6btCJqErnPZN6Ibn5tYCtGrpCp4Mj
Euszk8Q7nLRHTyNP5ywU4oSOGU+5LrhCaox/OA7g1t29+wzZiOZPOlmAuuTU5e7e
Z7XG/u13ZLHZxm44hH8JhcEUoCzlX/IvxLYcDweU+/SA+15B6cYS/65984GZyz54
bdCspGPhnIJqFk7cIJACB0rWEviObhlC6OOFKc+dT9Bh6SdBTbFvllE2uSOLqWTb
3WcHEaIZfTFBP5/YS7JncUDkYsNgIgXoKyd26JHsKFeWhXBXTvEVAxRsLEJ4iVGe
W1P+eupENqf3G3457TgfdgHbOpl/LC/VBX9yAfR6vU4ZuIs4lHjDFp/pEUhojvmu
F+kt2C6odeJ6w68ygCY06e5tJMWB4gNUPdys7Fa4jDuP7aLA8RQphOH4FKeHYjEI
iJDu8Cvc8oww3W8BAzKlcmZJDOi4kWhpumyVg09eEx+3xZE0SMsYKTNJd45+0q+F
8Yka/CUDKfEjafzqrM1Qq3Z7nqozGu/jlQ4FQqFz8Sv5kk7hlw4lZK8J/3zqTfvu
jHFIi/mf9B9oexP+M/1Pxz1uc8zvtqW9rnU4GXTtZ3lH2T4lft65+gBzjegI+l/9
MA3a/duXbfa+IaBHIJr7WHEXT3HRLi1mqUpmHkuZzT2ngD/Re+DB9/kXYjW0sq0M
GHKEeD7owGebCIHet6libISNgiKDYGUpSMEJbfpBJsVvbqKPuVYa0S32yXup9Jmc
ysAzFAoNJByOij1cAMPelSkIvBWLLTIh2fcUJiELP72rqAqILZQ6GcXicL7laqAu
jNnL/5si8JbeeX2BKvFrQ03rf8BC0KP69l5K5S89Tkl8Sx9J2dXgstz87gibIgI9
6+nLqf9Iub827zVCzuIGyYxbBZSSdZ5RwUCnp0UPTxUF3uI8DR/LJ2SoZcMlrKoe
i3A2hIi5xe/rmviHSeljHcDFWNRaUxwk3FyHQSPhRE6v0qWa78zCCYe+hzDWgZiA
rU1HA0+/PSsl5b3hK8IcaRS2dqiOCs0Jlrbs4Q64F3yqAVWWeFaBQTJdH/vdu/y+
WqK0ANCSrBi8btAjv1DVeGgOfyCEZAI91iaB3zfKPWj5i9knU+ev3OCRxqwZOGby
jiVkYAQx9LSGaTZjvX7ucNjjleW4+SirfY3MeO8XdCbAXqMXjJ9c2xtUwIEnCe2T
fkfRSiJpFmaNzoqOnptqYbG8b8a6/03+s+UmHkEZa3gskEfwV4Erl3aWmWlIJsar
YBVME8UMr/i9e2zmPWoWimuwrErPHdWSWaZeBE6dV+DVgxk0gMoqW56f0Ka22X/e
78SpXZ6Ou9D2PJbSFsWZM1qfSPN67IydLw9mByzmO0z5OlQ6I6ZNG3IOq6yJL6qm
xmuPtP0piediVkCmPS6KwduiCBw7Pr42avg5kTJhizzoeCMA4KWi4Pzk/p1uM0Tj
Hz6+4ETd7emkKqIu+LA3QWJaQ6qjagRLEwL7SOjlJsupzrYIHgvIyd72CuWVpYPb
Hc8y03b3qs+Dul7j/OxmhmJnkr0sshHEUR82NJOoi+mD1I5JpAcGgiMlGbiBiF3S
KcR5CNcu2DT/6T8AmvRV7vexeotMe2WkImdrQHUY54c12UnrpGFW7mQ1ediLJV8d
AC0Xf6NyBwPsrL3goZdcl3B/47LSgN7CF/AE88fZmTWipTH35IXROO0SgLlQqgYg
c9YSfvfiKmFItaKJF707W8VOv27B+ctHHlqWOf15ZteZWN2i8xXof2irbxzzfj07
eSV3a36hcB0HLSfoe6jSWWYkwUxZryeoRc+5iWSrvoYDBRhiIwVdpluhsxi+4koB
2r77fYKEhoNRDB3LaYbaTZzmjFy04whT/LrAyPuZyIRmDfHHP/WFsnN01MVun2X/
ujIz2xhv15Pl09fb0A/mL/YD3YLm//NIBJ/vK8T+wo7Yy3AnRKxQr4rXI/QzovAM
Rw2kvvKq4v1wl8hzQtPdCNZ5TjbJMEboFEr9O1LS/LT6ei183D7tGd7Nr2fu36C9
oVkz7yfdAIWGJI8ul/vNl1deur76gooSqLl8FgFpRMSWns7TKVcQ4H1s7/5dmQc+
LbOOuM29YViNKIFSjuPid5KCEX0sS92KMeG2mJNB0usBNhNj4D2ri8YPGP7IP3Nd
lB6S39KrifN3y4x0z093EthbYnFhNuRY0k+ZiYcEIQAPwK4U7slNADRu8WtACmox
FvkP0n5ueET1YabgcEt/gdUXH60JGIC3sYhwqJTzjEulYermXnFvTJqJtsxWLxm+
tusXaGwzNxZfXtZxlqxW2dSKMu+MRrvjh4sFa5Ek1f8hwZbw4wGlHYRsZ51sI+oN
Pm8i53QW5R0ICyNlIE/46reQS4v/NdcaR8mmaNB+gEiAhEe2bMbqWvO0ccfdlWCe
Ri+6s/pFfEuMtW82xUjIZd2wuA/35ig7dfInTkE2+Nxb2LkUqbryu9NtV80Rxh+W
+76cXSwl68wLbN3iJz3mCURZfu69nOoLNqIWkn23++jo6PQlwKeWGWLjGAMZa0bw
lfscuccg5HlUSaKjRaMToO6JMj8RUddoAhqEvkygcCoS4mUpQH/xNPup9yfhxTqJ
07DOLyv6LzfytF8ESChCJzkCvZoxoGA/hamLLGlcjuauTBrc3goZDORvMh6jRlZz
5ysVM5VxqhDOiTh2GXiiM69f5cT/CpvnUx9v35sRHaITcE6ABN2c8ZuRi7jpJu+0
2VTCbrAxI6TXDGDe98Zj8xV+cdLkRGyDlDNH0YmB8KHrwMCmXui41Ko1UQqoth8N
cbxNI9Bg2cS/1uLe5gO+510Y/a9AA98aiTbn/PAPh9ZFKX1gwyki9tzDzt1ZSv9U
Ttuu2cB5EDjPregwkUPxLhL9k0UWEz9X0ZvjDVNqVTrMtpx1Q0EbICmo6fLUSRBK
FlKknBH2+l+MWVMu9VL+jRGO8ly5TOyrXyZ8Ei346AbsPXB1Yb1IXWPHQTdcDb2a
r3YFYrz7oEaqvB4FQL/mkawDPLEzzMMt0s9QypL5ZJmRPAybxZeeKA7+LEjre+py
Lr74BEcAqQgzJa7dumOU1Fa+gLMOw/qIojfvRTAbJBeXOGH0g+VnPdgC2dTT4om3
Kj+OZ69RhqwmQaoh7evkmSIm+a2mJKd7cjKcQrQu8C4mvk7ewx33P26kcPSzZhuu
W9ixm2TLvV2kxuFZ7h2E/z0n8tnsFl4x7JrRzvw36ceBknoIUEOsVJ3TFKqkUSDv
A9T1Vtmo6O+s14j14BEAyn5iPUNHvjG/GTtzxkO1noccZUvau0Vdq1K4f4Cua6x3
+kNPCZMPlZDFZtvUpfiNPi3q2hNXz819qdJ1zb/8qKqRR1sgUqRsRYZ5BqzfI6Ji
TOwnN3fIbcKM9bMJh8NUop70F8IJlwiAtu8W+qV5ai1Ov3BU7giTSl8HrMwK+bIF
yK3rgH1bMIYpCu803ZSUay40SUOdnFDIo9gQeD/6RNXRBJ/4SZNFAZHxPYXqCvMx
4fajb7SFmf8l24uCG+sFrK36RT94kRelLFU/g2LoymzbIr3iUFHf+PV1gzYoKwG5
61I21ta9zwBperEUCTUH94B7ES2Po13z7YM6mg+B9pbL4/CBQvjq3yx5dM3+/VLZ
VZaE2tcq/FjSkTDqrgLt9dvJnA5J+uc4gdRXar5sSn+VLQZC93YBX3+6850bM6Co
S+wLtVBPvTHccciFFgBIM85jX7kUifCnFt6X1KnQwQXhTHumOsgu96dNdO+foyNo
yex97zrjrIxdQl/YstyihZpzmCqM7AHT9ORteuZqnNyoGMm1x7Dvsh994CLquj9h
jSjrproTa/9hj3bc7GTLs5qFUJBNeRbrtC4vIw2i25VKZulZuoluKqQdaUF/dPah
AdC3efygb8+uAkDV49dUx3/PcjYDLWe/idNnruaAoKx79YvqcHDObGVQbOs+taVG
25cZzb17/Gt5pwTe+eIbDrcJjDYiWBqLqX2tHrAA+trzOsM7ybaZrEsGm0PoKIY8
sDgJOkYyX8c4RjdcAQYdVK/F8fv8yB0vAZqJ/VccNfaTkAN9ioHVpZhTnTBRK1X2
Y/auqOcoCWlebKDzXmhlGBTC8lyAVtZIhkbxKZ2BHFwQDiC4oYx0Ekq8E8taVcKZ
FWlAZ6d7VorJnObzIJXpeUGtP2yCNfIKeyfViTD9fIS9Dw2kpyVE6HWRpFb6rpPR
WOKo2r1Mnj6WxwGE3XzzDY3PKDg/41pJFlJAaW5K+L3AiN1+WYgIFlChL3RQI6Zq
prWoe9IP+BVQWwFMpxxYuwOaXkGL0j3sDQVilrfSiaPTLzGUVzPUhxOEwfdMtxak
xHUAALxu/UCrK1pmpVAEDafgaSPGSaIPruUuYxLUkzZcYWqx2UTqKBLgkYgTElpV
2d9lKm1t3VCnzW3pIrcB8XYzD2WglZ5x1SouXcNe+QgacDqy4fsMnK9UdU54rgVP
vOHj+eTiyhMbFoX+7iygPgieTW1sW6dm6VKMp6X1Jdaz92voa9/loN03rfIRyCb9
pMh8RlyThuoq/GgQfyyfvbYp9rcg3XaWAwsLtH4zV3tVL9IABq0AmSE7TgKqk5vv
mPYVtRGmvXPzbs6gNVxo4bEBrjfhTDI6IcSrhqQ/IYBIwX9Zjqj++6izx/TrIev/
WLfHu/QZvh93vqo77Ozrv8GRKiROLJyOkZ2XtqKH6/9WT8MQdnvJVmVxcTnPsr6r
+XMOXJObnxpplb9J6UNi1M2Qzs2DiFrEPMpDFxNEhyPlQRjcsoT5dPUUKDyTH2KT
DsrOHLYawbAdg/tupO1uH3H1mJJp2B71R2PrzijHh0NkCFQ0TES/YUk2bnQ3RSTD
4HTHAAttruaExGAyn3ApCdlceuTn9h+dO5v+9CI9Mu9qBFwB/YYjZYLHSqcwhGYZ
AbHkNmX7WicMmChqeoKxhLIykvCL5f1hLUc9KR460/sP9+3RNcausWSOX1RVvBE5
tCLwFisFwMDChrdS3VrQX2bBN5fUdJe8d1q0Lghfby8QmlWDY+6BXSRr4XTsCT6/
DaUE3GYa/2dq5+YBMV5ll2qZBoKPlqjansvXMcX29IDXvDnszW/GakUENQq4mG4a
khnEZyFqkXnJnAdwWRRroyrAfprXKmYaXvVQRU0GhTCqm/aIz/gBimjq25qRX4dw
XMBRinOSjeSXrZP1vh7tW4tXwBiqaF81mvRBdR72FRTZKJBojISDeM73r5/Vedxg
lJyCevVoFI4NW2Cb0aTC8s8NUg4BN7ClHYnVwxAttA9aqg3H8n76cPphbrApUrOP
pGuRFO+HEsUj5mYhYahweNMbuTuzNKtsu2JLHALl7fdcvb6jSzbcV0/GNM+YDysx
DAfXO+BxarC9l8Mqd/N8jWSliNjfkmpCZYXpt/FaTv3xP3f59nFSSFhAF3QUM+DZ
Q1lkz6JLYTBYpLQAHVETKf43Rn+d8k/ySFfWhqjWLBIYT9x1jSUn8Q78zKkzruTa
YAKMENlfBnVHU00aZ8zDlfzIvMrZbB1GUELNIkQSsDqxt93Z+xbvMsNo63VVhskY
c9IB30jNPU02mn885zpAsr/4u01F/PfKKLOH3inz7cKLFvrFuU88oNEBQ3r/MKmr
QR5E8M1dQQBxXK3wv2LlfxFiUCt5g2VuG97JYBgTPWwrNl3DIULTUFY/BOBoUCrb
cL2y8UeuLGeEhC5A6ctATu3QZbgykTo3fagLFejxmN7Fj3oWVUaL7AGbnMk9n9j9
OV74aSD0SW62i919euSW/3YuHzuiVwVSQoyulDdwsfeFNZgaDLXuBkXMmC0yrPvh
CEWohb5pQGB7LNeeWW3aVuGLaVmSGNL+a/t0g5LzmKY+wrCRxfv3beRRWCfC2No3
SPI8MWmfchEHQTT5yUVNtN7mzSEhEwLvCr7Ykj9z8oD/r5cOFhoXyh0ZSo7N6WZc
TWWeWIZblrqWcKKw/7WPugdUzMoYmXwlxGhBxb7QwDunkSjtYbGT04Ffay5UBz4C
7DJFK5ax1stHfrOjB5cHm4zlqvFAxwRM3hCgYuiq25yxLuqniuI8r//GnaPo0O+d
Yr29HU2vyIVG6R+xXnUhnAfpmk+lUlX86NdMeEdwvbR5xY17zCJOlT0h1u4uyWZj
QML8x6vnhjFk5imOEKp+Wj5fOaVrAK+pg6/S7Ax9BGV6V0RC8WkUrmvdbL1Xm9ew
BUwNPmEr1/6bCNrVdY2+K9jIjE6XBAB0Gcrc9sNNr71JxFP+CFhLbAFk1auJ7NO3
bGiARVVW4nWsRXwhADj0il3oMbbDgeJHxohMr033fvHnIok4D+L1cT5NNib03igJ
v2S89GOAXi2v2UBBCQo8GuwN7WFP2d5vKr/Kdho+UVC5OScLAVnv65ZtVAA9bzpN
MkfTBvszd2B10+9dZ8S838PwuRzCFp4pGjL5rBW+ZghB7Z4zk3D4qOuukBISwT2y
8gbLmQivQq6CpWmQI2jQDf4Y9gD+rKP27xBMkh40bOiGjnzfsQ8fQ9aBUgMRZA6V
4rlibgUfjjM3PxXKPzQoJmBMIrx4LdHAhpm4fUPtKKCOZY0meLleGCdlY+57NtTx
4TZHRaWRyeUkrv5IDjbx21qbSL5DWBV17nbMHyUGDy2OPxIphqmTKjSPy+K25ae9
04T5IFDPku0B++XMGwYqN3j64CUZazXrcxPlDjpJAw4fx6iX/JurrCblItJhHXxa
qa326ZspXtoQQpV4BcJC34UCidxGtgsBFnBXYbmC+GaqG+VExM81XabAmevj00oc
T4LWt8NnbMaK0bCV+/atWc1hZh04UFHSRGWPtFmGlDXEGKlmEqMjrvDFX2CT1glO
bJJyqHaBSZ1lPZlQAXaHOsdxlgeZ9a+40wqyAriUd0ZJUk1cqr8PLBeVBT1suTg3
+l2My49HeW5ycrE4Muj/pQwY9UyLOJMM0/lY0z+tdAvC2Pt/jRorYYQrL402gTUK
MS2AWMhUoI1t8rzbupGjb+wrKjjlZDbOXnACbcSxQQ2YtdaMCGo8OHk88zJh5bAB
7AzqsWT15XI1jFMYqM6YjmMFdfvB7skuMurbjbGnAGPTwsm44W+ga612quqVuA5a
S8N8zQQAkGYg4ixANqiMzsCsFWLc15LNDvlVhAM4B0yQ2cOUXe7BmGOplmqKNk9S
H7Fr+eGKxZyBUle7vfUY/l4X+TJze4LZdKxKePzbVDMGoA61toOx75wVTr7CJ5R6
/6rpu/xWw5Vf63AM28au0IdUlbGwWYFvpvdAcGiTuPrqp9uUu2SNFqfLRxHOaqhz
zCvgxEarXdjwbAzM5TrTuoomRDGGt3DI+yCrJpv7khmL+3kRqyd/7QbosI08MaDW
UJLcXq0zTVWIQGyAfETro/iPqmY09XNLb61Pcvuh6zVKbMpQZt+Id61SDI5zP6Kr
/9nun6c5lYG6JeHNoVYK9Ad9lk+81EgPOUhbNwjXE4xuHMUnr5yVgMkFkA7YV8l7
sgrm8r0BalOq+II2VqHZpoiuOQ+jWUHFv0Oa2VIw9sG2IMfyO9aKxTjmVGSREBRH
WPuMZpV1mmbTggwJUYTAkIxd8cAA002XogE2Yoleg+g5SrFR8e/JXYxlo4ygMQgK
Zc+OHHmszIwgK8g1R1LMhsIQbn4Z4aKF2MAgjzpiGlkGgLFlXzrmIr1ez1JGe2Ky
v+HOLuxMbPpCezCjQUVrJ0GXZvHIHNBEhdCQlbkFp1D6CBn7FiBWinlk/aPyM4pS
NoRGHfgr/gROVDOfIhB2ACJ+6RPBSCZneKKJf7neCobeXPESeF5lItTj1e4WwF8c
dSXdsRKq3oryTUHaJjCx4KhxG5X0GKYzQx0ZWAId8dolzC5XYdpSXqie/pG8knEg
3K8xuX+9jQTg54jt+fiCWvu9MNQxbDYkBtCDdbeLTMQ72U8FuSz1PlKiikijO/A3
C9sibxri1tg0ZPl5YSHgIPP1sQv7exfbxa7tK1ssVzpgTH/O0ezL8Km1L/OJeV6T
mUjug5q1j2/yRPJl9kcz/ohbnGKCQR6YUZ2507MS1Fuu5JNXxlLrOUbz7Hmo6vzM
Sf86Dk30ERw+1DBW4uZh2AcIruvaOauCzklOD7gZCivkCoD6gayPOzr7BWIomql6
yAZHSz46hXRJJqn/4oI21NXxM2H1dd6TFwZ/Dohu/Ac9gAMaMIFVFZwl+lV9nK+Y
lIynLmJzIKUivMJCVp7cfkjmdi12Ynlqv3r5FqSmYCIaCqszcGxvYDu9PqjCtdKB
z54YqHX9Op60TAS10BBj2wqONkzBpUyR5Q1RYgCLYTv0VDwV5lAcwxW7yhnxPT9n
+3l1JNfmlp7DupOKBcYCT+L4KVlxZ8Ba0sL4b4/L43TziFcPJ50XgdG+6v2pF23L
OjS6hzqVsTxl3eI0/yLnDmazRCnppJBVJRvMeHOpyb7rfuQZj/JvdZm82F/RvzqA
WPYkoAXy0SshQzcT88HsF2MzLC3sYQ0QKa7/eG4flrSTockKkVCjfdVSf+QRx9CT
Fe86OniiYkzpNMgczNFd0tXN9yyrrzXvjmRbZ2C5f9VpXlOOneIWUaGFnwK3CzxH
5ymoe/Y1xHH+Ey+MZ43JFnHexAsbG7K5JufCPtRhjsuwgmHlHjyKh5sXtwDN79o1
NwdZBZGhwLRm9Ub+2KSD7a2nCbRT/i+HgRaoV03w0OmbFEHbc70zcymVZPFj2DG8
xOMy25a3F1zFYI+WbOTdgYMmh+6i3nWKld1wIXL/J/y1F/kmiQBGuqO1VO2NvgN/
rFBcbrVQnwBs8WHwk9W6ieJV5A7K9BMEphhsyj2FC2FhLdVAjh9JnmAqEO4FQ24C
6N04mefaNWSWAxuc2PZKK2EKHyCRM/NBJq8I29fkBXRYQasAVhyB5WWGJwFGs2iG
/p9XqHlwc5GETOJtpvIcQnVVF8HAh8rBF9T6hhFEgbs7K3i07cYZR3IHp+gTYVNj
RCb8yF2C8GJxdUkhhmupZzRCsIbRctpRunLz2mzwtzrm+AE2lv9CJITlYiZ9pUlr
4XlCE4Wjl3WrQFzINVPws5CNKsvQQUsGjjz5yk1H6iyQU7bEekVTi5IJ3C+0c+qJ
N0brM8AbZgDwhwk4o21ZtUjMGjBeqN36hCLneMnDkzzJT/8ZWw7eP2bhbgSppFYA
tZWzIAAxv0Dk1Hr8JMry+TIxCkeMCI3kbo97B8zAL9QHxmg9RzOvg70VfSIuZ0ff
ARq5TaZEPrYmgSDm3L1vsv6wGFj2Q0USfnPign8enw/84Gm8TmHMkX8+rZ70BIPT
J1QawrkfVPOFvkAItYtfEwoHbnegRXs2JhLJ8aJDNHk2bzSVs0ed8jCVD6+myuHv
hoZvXZX/NCmC+kVmf02RBrpsaEWaASsz4k12swDn1l1D5bexQFJAfIGtxOYOKcfl
yFb2JSXH3iVS1cpGkQV+3omCo3B/oY8oQXQA5xeLnHrNwe4kx1+eo1B+E47jDnyh
/AD03e2rEmIN2Z4dGQ1bW0GpNCp/QqO4yCJzKLPfpaOWzowlsZJ5WyYMWukfO+mc
ovguwGJaJyKsE3fWfaD/Vpsc4G4G4sfNMsGXJZhVJx3eZwj3aUR9YjZWmTfOJ/4I
mquMkuTRUN8/6/ImiRTuF0ldYvx4K2+EkmhK++iLXinClSDw70btSxVbZExur1n2
wmIHJLWSxTVYnN+3s+F6mDvJ5X8HO23WxHLU/ECgKJsmk70i+MaKq6j6MGVnRUvE
bWX9pnzT4fEae59NCyR2TePDTmIj9xWD61jI3OlrPhheMC2R4jNong0SIn7F3xEy
8xcTNFs/qHG6iI18J9oikmqGiXSnwl3N55lw4eErgGacW7nvvi3120KTycuKC4w9
dLluNyMvgJTsxjp551To0tDgTHWP9cTeYcrUessmCKzEZ0a79J8Hfo8oqGxBV/CZ
JM0Edx5IzfJBa72Z5vysuNhEpoYyhNiIt+qLzgdIVTFtkrNIzXsvpmrD8+9qJrle
DdAIjmshNQhdjJ8KxGarizw/V2YdBEIhM2sQT6WPGhv+IwBS/XisQdrrXfoGUoM6
BtgIL1P8XKPSZL876IeEEFI+Ti7cYoyE9HSFKYhRdEcxNug60aArplEC6BXieeOX
9xSn/nVWtXit9qLHPqx8kZVwh9N/0Bagy1+pZAJRO/JnxZTqKpE63MuZm42Rnhg6
KgZ9WyfnJKAwbt/D+rUBrjAyNPSOt3piHstR2BaskMfX1MPHO/wlkPlP9Di+n+8A
UCmFSnLvxFocHyXdDRK0RXVR2G1jJCSUcG6vbsF2kCQvhB2c4YaZpCR6MQhcyzfI
220nTJ7fNYyDhVxaACgDoRUb66SwJxYAB/lDYb4uentHkjlPNzvRimQpoQ2OGKO2
Zm52b7hlfQ5mTdSbYOU9wOVSOBt+6pgbGX4yjw1x5NgII6HI6Ptrfecp52WofwNS
aVcvTDURzhq7+2gBQfTmLCMvC2DKH+zm1te48K+bKKg81bfR2FPNpQEXOGv3Z9rI
4G0PvOa+ltZTBdgF8Uy0ft5fqCr6xYTuKNe7z6ehlWAwWYnon7XgL5r/68rEIQ2E
2Wk11WKwzNHGh44K7ZnHDcp56C6dlgXZt53mkhrijxEefK7NqdR4ok0gFBgaBbxw
hODdt7LZb6Y8oG8BV/oG/w+Fwr93+uZ+BZ9WlK+XK+PemY6Fi1DHPUhnEp3ZCd/H
PWIUnNiSlPM43arkKp1/pr9bl5LT+SyPA4UZDOSZzYfeBhewSR1MNVJn/N4tNKMg
VG947P1uGIGPNOxD5mY2Ly+TOwn4AD40OfcFoeSm5lVtxY5t45Z178q4UF7jNqaY
84kbZVJsX77X/a7/Hp3FbDFBYpgO31SWlN+DDq64LZGjbv5XOLXQ+/AO4w30HTjB
uTf8sZw274Ax6deVyzwzlW0Sx2t+yUIbFSCn0M4NGGXT0JJJ2MbhVGigX6ZXCYzr
A9uXLk/lp3JCKri5ncdTnxvAJIsMDvF508ufJpeDv3HKI9Xc/GnJmD1nI7wEWkaM
hX0ifAhshSJnrPHntSonCBmV2tHA2U/+Xm00fbkK8PBWLQWb3ZHhG+1zS8rCA+WK
Cf7lm4DQw6DNqdOgb+KJrYVfuPCTEWE7FmVjl3FbqYIOBSsOjGFJ1GqqIDfFmndR
3iqoJTvEacoI3hSUL5KJu0AhPlkTqhsSTkwVZrTtWq/zVGtDJtWq0jOmYoLpe5v6
ZPynp4Ep1EiwRgRjpjc131nHOrKgWYuYkFE14paDXWggKeTJoAVIfa51yUQQHwJB
7fABX2NBUlJKkhZOxihJjUlmLYFzTmfwGu0T+ukyD7iFwoV7JgW4xHUAi8B688BV
70M/FA58Re2MhNupuVHpTPm1jorEND62scOs0n6zKvd5hbPpbPGFgy40xg4knA8R
H90aPI0TAfZSQ28tjcNLoiiPBEFXSc+JBpedkjyFOtx+mjgvBgxIMDtoaIcD4eMv
chhOfBEDfY+wOwIfSyRqI8aFzS9vbiT1qwLWS1Jnc9JuKSFwI9LBjwKUzhDIaqsT
1jn4gJxLeOasjnbpuF4xG/AnL+TPrmE5OB3Q/34WGcaSG4CU94AlxuPJ52g7YGzD
v2OHmWykVT2HM4kHyY/Qd1QzECOV9ADD2sANMXyVXxlOISYrVlHQV3G+DJEaHWH3
bGHw9LanygBTDI8e6Gfgu1D0OCNi9m6nfmxQkDA5+twXLlIavmpyQAUqDufFMIbS
TbwGlWiLDTvYVyz5oist7V6d+fxnSq++56RdDVuvqbjXrT6zaVXkY2Elqz/21WxZ
bpzMdRAffLpwt+lpFlRM7YGfAiI8sjzBmPZ08FewfxfAQ8Xp41naB+xWOOx8qfor
GfFehlv8d+FOrXlt7qAl16pKqnmkR0OHkTLXrw5Px0Q35dRT7OEdDg/xa1aUp0AO
Q7gYxpYc2Q0NhQ3UXvXvK70YLWJFOG4sCA9sE7wQg5E7qZ9JnNxG690a2RP9qIao
GXyPNsj54zB+4Nrzn4XZzWdlClDz8dk/5y66Ewn+8NYbS9nbHJmdWjHaidKk33Y0
WyTJBw2Q4L9dq8QPAYODlerHNo+VhvBDbKeZ6oiPF80+wjT1DYnXJUGas9O9F2I+
CLqJPifTZIw/uh7FjsqP0hRT1Gq0Z54giMfZUuwzV+ixgy+NBHyzuqxT6B7D5jYg
kwsm6Q6gORAYucmZeNxbv/HFY/ef7uCjunybX+/2IMUeID9KNtUDotatsVEyEQhX
iVx9TwbtJnBym41oSK7RR/66bRNSNbCbuFxk3BNUpMXMda0IGxKfO+5zslx2BfJW
9iZdu4TPNJuruJLT57RXivXFJjUMoBMQeBVSvUANoBg3SJwAE7RGQCHgNYIY4uFf
JIw1xGroHeevpnHTSCS5sLTn07h/cUazmvayGKoyifa4HWWP6thLj6pBdgHNZGD9
CeiE59BJ/HqiWg/6+zojqVeGEUveFAkWFc+azoOrqJm4scDMaVahGXhH8n8JB2uA
qv/GXNKscOnPMqwVqIzqkvTvZmNd9YnPgFGREWClg1Q3Lg2TCipzatI4ueVQDp5Z
ZLU5/2TJRP4EuLxqxPmX66So5zDCAdCSkgsPp0SkPjSER729VBkD26qRF/ZjkPFv
euqmylzMn8ImjDLq5Ql279NnhSKbxQ8fzJYZ94PH9NcZ3T1S41RvbN5SmUjkw17g
bcr5HBkZXM1A2dP83NjlnlsSCuRDR7uNv8b3OR6mE9+YEOUwNzrUDKcldHyZHDK5
0B/J+QYbuJ+RAmz19Ec6o+P5ww8fnL8QpQuhQ5QmH9WZrnS2jN9IQp30voBLfA2D
dHt5GQktvLuJnKjIkOtSBpR1GScrZqBRLcKKyhXVkXwBzY2O94HDQSuRqRr/iCMU
wfilXomDm9+1XQToKIXC2Y0XpdjBYUM6X4Od/jfonoo9ZxMSp2vKl0UP9lMNz+TN
VcvIwv+3e8oDq4NfTSoj1xZ1PNCOK6q0vrVJn0MKdM0EvtEB6Jip9QkfjaP47lef
v7DtSkMy8t9SWBj2/P5gXgBEmXe6jxgEhfAHkEY1FU6FrR9TRrKm4QwUl31Bo3Jg
71WgUOS7OXkxepFhLVLcAVdb/m21Lu6ULGze0Y3YfyK9u140bhVllAxURZoTyQFx
3GAR4DUXasQ3BblvOLthtU1SzOPAosd2T7R/Bo21OqESegxuKO3Hdgu0l23FMmcQ
j+Zc5mbkXPC2GedeJU4jlvwJZzHi0uoXkeuW69GGl/A7iD5sFHcQ+CnHqCU5rmal
pjKKtZxCfl1IlSjk9YajOkSeL2U3WkwGZ2qEQyNIVn87sV8Ic4yL61PPrRVP2G3U
wBCbNd7vH9Xus+FHMIcjaogthnGpUca71YQqsf+hz/bw1C1DcGOT2v9fv3uUGKl1
s+5ijtqqXY3c1NpdTe9mEXAiVVl+LrM2yXmVzAZZ2Yjh86AFHfaE/mgTq4y+/Hez
8HuWWOqO/75837Po+3ewxYNVwnskKoniTlpKM92rzOn0MLl3HO1Ku+djoxTKkFcQ
GhOztVQCZxsA4+LaUhETN5TzU5TuKkukveYHrCLRfK6vLOpFYEldZkn97GnUQCrA
FxF2T5MkbTGZooeNProRMcurzqzrMHmoYtEf2qJJh/yXanlIiKWfhMbwOwzuDbFw
L7KqpUx060G2Td5TJ5WW7jczgBFxFbxqbKRL/6bi8k1lm36TnA+L94YAlD/fCEAa
sF1Sx69B93HvKi3JnsruYrzPceHPo74ozIfquUVDWYlYB9XaB/RQbW1qBgy2Ajpk
/eC1bypXElNUp1NU+D/AYWIYSN3Qt9LlGL+WMZpsLbb/Dax2vBFLGf3Qx/XP2ErW
8deZVHK1AkqdW6l/hGYlgisgh4lnwmtrLy/fnpFqchsAR5XtyZIzTabhuqTUWCOS
++MkSpG5bHaJ/P388Nhkx8DmsFJxylXHcTgtvGKFTrOHTRKMbhAG+8CmcSp1UnNb
pw9HverL6is63Lp9tysL7NmL1e1U9QEA64F3W2wagGbx2iwyiNQ3HH91jQfIVPg4
hXeB9wJfEKl/vXqSuuuf3zLT6j2XBBGTtUF/CZD4DPnR0cLsZ+oyzFo56gd5esa/
0xueJxZn5/X70BUPbdpPxjhuW7MWnDOsBPQMm2sUot1sKLb10Gd7jt7+/8/2R5aS
gX45nUpi6x6M7BonUnJLtNgNJYvmMVSz4FpMOQ8AJl4Jh2SNwCRMI/adzcLSlYIg
259O+MQ97244cB5fzX4ixRAo+8DtCLdeDSP8R/WyGJzhCEwdLX9uBLkBp/LNIyJS
eKA0pxseehx+AUYsjAsir19oH1e9bplqTxnrq4XXr5ttLnFib+imZelfFfUgKBZs
bqFoh7yEtHFFr6cw6uIoyWvKiVBvaT1/fx8H4kUsyXlf6Ajh46ol34tgSDlpXeSh
Xm6i7GeusjQBRYjTDtzBUyjWzwhLcJBM5dgd9py7csUmHEdzanpVbZD9Xc/HBhBc
p3Lxe0+OsmYo08hfdwz8nfRcmm+3evzItl/Z0enrl9SSTZhZ8pFzgCuLowQloAu0
pm0W/h8rIF6ZhryGS5iokSEU9L6xCqfRkpSpOu+sRfT7JQLp/oU6R5nIv4zPybST
Ex2yDa76W7M7LgeOXpPuFCKk+oNMqdfO2w60Jq6lG8ACV+p66KJmmHFiTcD3g3Ub
DHp9rb4hYywPTwvq3jo2ss8v0ao+X1J/NV7G1nF/cwvWL6a348D4k13iU6SMGZtM
tyzWuYnkiG0qahkQMD0wYzpEuP0YQhQvcsqiovD3pssHDqDHxnH+1WRyfVW6hoUH
fAQ6gLH2hgC1PzhbkjJxsUEWex/hPf4Tflajx0ZyJvqmdtXanKNTNH2FBG8ytHa5
fSQZ8/8t3Zx05uXvUAB4rMzMewlYcrg9HLZnhGPso/5zIgiQgIHgxoNA/x38qd//
5kOf+Kkpu2eZ0FaXCVm7Tq3j1ou0VYJaup4azBmWd7E5sstTwt1MbA6lbmG2gdc0
fBElAMIjgY9ez1Rim8dpbf9V6F5CG+zIq4nZV0CgUdQIgnjTThk5o7L6c17L6nFS
jViW6A0kO7lJtgCRQbuoUypEj7m3IBg80FgazPNVgBXMsQ4X0g6ums3hlEti2ZBF
Ccx4mjUQeQqzAWhnkM62qCbZ/kXlN2oXOGelqATzHY5hL0/Zg27ZeC8xDPkhj30A
RqXl/sPMxw5QdPASOBOYyP1mVn6OMId99HPG2T6AEuqhLObkm1ZuRBQ7VZ3f5OfZ
5Je+YmbBzIiUdyl/m3yDczLTXmVt0KWf1N1BZvcRZiLXGAwf6f/6e2W9wnzRWSxP
aXipsx+sedWSHKL4nzaum2MVuUlM1J1AR0M3F8U370QB9Qdf0pWB6s2FHm2sIwPR
cneQoIi++URTfeWGglFdo/24ACYHcIs+iylu+SJEjP/o6i4y+Xvv6NG+JU12b1R5
rOTa0aNDPZWfUu46/CxcUXQpzf+oSTMjFrYTlColQUMoSRxWhig/v12pzdTjWyrp
BVzRtvInLl42ERHMQ64GWqTcJxFU6SzqyOywMZjRfDOFBHD/mbZg21IowfnaX8RR
RuaDZ1fJmrqbpU/1c025XU2GkCGS5rVVwQEycPBe3JlfxcTVsVLU8AbGFsNB1vrR
gkPAPXhUYaK7QFRX7mfNzCorpB5T1jGyuGGrj/crj83N2afYZcszeMh4mxBTsVYi
IwHpcDY7Gak91rKwPnHczBqtOmjnpgfFnYZzsLWiYXUZFLmrN4PWIYtzrmuyMRP3
GrI+xSWFecT9+B9LQC15dZkp3/1jdVOS7oq7zUQC9P2FuuXtJbKZIMY0XJGroaIx
rZseZKO//4tkAWXOZqhaBPewQkieJoXJ1qryhlG+6Na86v4/jmdVIJiRES7F3GaX
y/Bf+m4cslTZFZrwGC6EQ9DSFgODOp9J7NVEdhJVUcGhirKgELwA8fPeBuuGc4Eh
+KFktPESYUWgWrj7yA5nD+KCDYDtiUEryQrBQuKOSOiSfhfdrT+utBpkVwejSeIT
1oeIrVfys7fCOZ7qtpCe6hMgBHlAddSHxOSqQp71vkBwYqg/1RjMc6cXOlHmETnn
HOrVAxL5yl5MghEu5iEq6t0TiQDu5a/+WSVVvdn90IU/Hn0XOERsjt9fP/l57ZYn
mmx6JAp750UWP5tBOiVRlrWeG/JuzPM9/PxKQlmH4Jnf8p3ue1KeCn1dtarSV9RF
Jeu0MV+BCq0fUqEY7cVCDYAEB5j4gyDyuHnZtteBTESNJ26Muy/L2l9mO6tzReRl
+JaJnDGE0teUqig1b31WQX101bEoc+u6fcjTZ2TK1b8TvkDB4ayyNnvl1/EHmb+n
wmMCxUyxNG7qYIIlgg2pYlL8hGqzfIlDeygXQeDTtHoIg3EzHWl/2afcdAzRgd4E
kWPR5q+uihX3XMMNvJe06ksKAG7LWHiH4q6WRN8ZSalSnQCub5+elxnAbqmJHUzP
vZUOZRtgNUmI2njltJ+3AfK3kLbrqkAr4YCbErWDn7iPXIczrMi3JF9EpWE+Zouc
BS4jnBIZvm2KLPYG63OV2OFYCGyBIG6KAO+rx1CjVy50lCqImERG9nPq83ZXjr4k
hfc9gsJuujQhAGadzFAY4xcNM6jEiuDfwOiVSwyVfeYlAW5SNSLYIvcMb40BkSZ1
Yy2ZKqnjfbHl2v5WSHtaz/veiM/yKRvi5/xjYEyslwcp0bhE5yIlCNXPV4QLNd+F
3+l2XdAZFWeCqo58CKY/HlHM9cha5bb595KFjXFkFYzVi+6/AbJu7zNi15wn7ne8
Po/KD1TE1DImk1VgtLJWMcB/gdO8OTJTHK/qzc5ELqvuwKm/gspE/zBacYDxHjgX
yvBwIjc/yY+rTOWpPAEq4tEZpNAcu0bCROKFPpAhUFRV0rTu4D8xpRvuSAxscnm6
pY8HAGXlHIT0ELc27WvQHMZJeGfIjKqc0xPfd75ndLPWe4iHC8JDNvdQ4CBrMo23
/VbyjtbBUn1mh2DcUNrGQAbFINDl8PXNMLrAdfWNVwnaPMqouKnttYYXqGgtiaeJ
wUdvkurgtcec0wUKyzEJY1C0GYpYVtlejfBoIcF9u9MxJEaZTk9/PGHofMfQd6Sc
2CL2GObSu37IypnT3VZA9ZLaq45mDQGdx9YROs/UYiIVSttfOy+6ZaGT5WdiQ3+b
IXwU/yg+bZevbOMMuJTntBgEFPK1/9jUuIq6ihB3CW2FiHKZF9orcjnjQFeEcy5H
oL+s21CiFr0qxtR05V7JLRyN3MAfqwke2Hr08olyv01TwbA5jLl2UnDd5oEsR/mK
o61NY48a4QbQmeoGVJ0ven/tjUt4I4FCvDntW/BU5ey9Ai1MXkQgxfTJRyVHUcnG
iVI45BIqMnyGJ+batUwv8L8N0ToxhICoEhulqbfyIUuzM/pBAxdg16TDFoDibecG
NI5fSYbTFmE8G92k6vgwQbCDe5uvpDCfF5OHWWSvxMlB5essAfUGkFjlFHpWUohZ
l0oUWZKPjMORhOLt0iL0dweIkBHREK+OdhLjeHMNuRzCso3Ep+yjnYsit5pTJR7n
ZMVPS9r+OfodlEiCdv5ZL2QtqaWpQmq6pVK64q51LTxi/aGlriaGB+2bzqQulq70
jCgxDlpqi3tLt0za06e48PIQqrxTKVhiQPUz3IXNRuM8iDXbGIQeSFHZ0MaWxLwd
WvZ8/24BbnsdNHzcKuh0QnjQG8J5LQP/gGK4VspbMu40QqONuuZhnLalfH3bhLxF
HKmOBu35GOvUb48bVJ2zT6ThTAkcth5oi/8aoWy51QTlaLTVFUIl/znKqG9JtE8g
ZHWG1C+S3f5SjzKbE1koha9sSQSbI8EgnczFyrZDZQf9yDcnUMfHUriAjowIp8ZO
6d29JFGCy96DYmRpNgBMApOWIg+yA2hjTzGRqu3WMB+mJRkEUUoZwzzR3SL2GjCo
Y4Trv5E1f6A5c+5Dfgpp+yVPXW19FzUf6VvfX8Yd16wtt8HDbQO2aAVfeb8r6NWs
ypuiTxd6NRPsZATHVyLVOGgwMUn+lWw0xOvTP33/dKVT79/GwK8ELFRuUL+Zf6DN
w80d3C5m0TISH6iVth4VswCiMrIvzh8jbIUUr6Sct/zRuqJCgWw2zzPkYc8sUUiE
X3R/T3iI1w1yJ1kLNZlcfR0izb6fNp5srewPfQ4x6jmv6Mq3G/VFQ/i+moW59Cy+
nHjaZz/1JuxK4qsOgQVt687upj3i3jxqP7D5IQh49B/SY5VNV01r1EcEEzTYMa/F
y7d4z30vDUHoVWLGr93VnhVTLlSckU+mrwO7D+9Gi412urfQkFL68xcASGwr6k0V
XMEHKFU9r+Y1w6o4YJ8ljIeIW7Epg4BqD0FOydhhYKx/agZsdvCHFxZDyAptJ6Lq
oUz5OLPo5KrCtHIjU+btVVjmUfBh/aWFeMKFygtScOhnNMuEc0HF4reMxgA4QnK6
mJq+I/amTYKVdlrXVkGnjyvBL8PcJdKrWzvbHUv0yiyvCiSkq+z9iPLqFGFt2fA+
Rzva5RZEfRN6ngL7KWiFnS8H7Au7xxNPd+aVpQSLGl6fsTuGdajhaXxd0FWC1ms6
RlZ4AbZyDZkSwulr1iKmSYeWfpKfPT3TdGXXERbEJ60jSCn9oCkkPPNDsNnvFLTi
IUMKw8tZodqmmwTgWmSfuH66JpF9zytW/8WIFTKzsfeUtevWdO2opyOa/9w1HAbe
IHUiyjGLFsVQB7oea/P1wujsqSSQ86yIqyirQTm7ER31MTFwZUtliAizSJ0CP3Wh
nXsug4CfSu+WbgW9531LgOxmqXNubC+vM2b/9aOfA3AA8CyCrXEGbUzc5M9yOfnk
5j5+Szt22jInBw6v0fOOozzYLBLK2In+fw7mz7PW32HHgbONbBTQ+2oQnO0ySlGt
hs8oGLUGL4QItYErHM9Dwrgrg5hF3z2u9XlI1tEJdKs5PFEZAM8UMVKYBaCfljLH
FGrKX6C46nJcu741bFkrfKB4YucG+Iiy+Ud2+m/p9AGn7A49+2X8k4mWjCE1hwO3
ArNSwW9Fx9atiutK+s+f416na6Xiumwo0rX1Z0xuMyK8WdL3AmR88MyPmY5sYXQX
ZKKC84UmAy+AF74WRwLHYkccRfmSJIJ52Ahj73yacT5XOJkD/HOGhDMI2E164iNI
dWN5tGqIUAICwHeQvC6KogumdNtCJdNT++tdDaVtIM4VdvTs6MCV2NIWOXXmhsT6
hcNRzJMuQEpPcY/QhQw6jYxzAj1Rux47Ajyip5jFQvnCmHLLZw3qYVKTkWT3xqLm
gEvwEz1fUg7p9JqdPfKSgmkKw7An4LMfSbmD5rXvDGlh9juRdNAlPm8cq1hxoWSP
HjeRj7+5TKNXGjnoToZ/91TPyWxyQTR9+ab3g447j4SIADA1+xkAoWDE2XUzTqXy
qzYkexN2jDzndtMD3mfyxClFQ3V4AxW9aaHnXkp+36xz28YmnW9nkKYjx77b311q
F4e63LBJhuujK/hBmPormvdubRO58+DkFiIeF2t3/hoR4bkP8RbZxE3OkIw320iK
L/bGTa5Urs6HViZCGZjbiH0qEfRZQJG/zxnrUN+a0OXW2w+YELoU5i2QXMrCmIOC
RNFeFngKQ355Ku36DuacNWGBOkpgaEMbsEJavAwLtIn1lnU3iyGnosRiHFwa1FpM
BxuBUun69YjaijscPJNzZuT5RG8KFrmAeAxmvEHssg5RyzidZcVQIxQZpbIRVRSu
PF2C7oCxbazhUDBxaRt//Rm5O7p1Uj0SJNQ0tnC7QcJQq5chMCu1KGMb7fNNtubT
nqB1mhTodi3s/6S4DzXtEJvdHJMZ7IDvw4tGq66Xq14XXmKRDPCXr8k3rLV9ZOkO
RYF7m5E3nyFU97HDlE97kVxkNfQ9oj/vY0pWIaUPI/96pSw2k9ieJ4Y43ko8xEZm
xHmomW1UdMESwmSMYqixoQK1eMtj/2P7DjP+3hn+ZMjhWZw96hFbNPlFqsjrAB8C
v3TllaUZ9CQWQZxSVBdpJBQV0rwyCcNdDZ+JO7NKMDLs6IQ/AV2fEMaCIORIhgPw
a91vSwNABefHTW5UAQAQBXQ0ZT/8aGB5iQUcNo0pTm3FHzuprxh1zKszOUdMw35T
1VHOSNBBvHpSFvbvz2/d2/fazoOdNnWfi9Dd80x8XxpxD/w1EO7FvXdX+GrZYFjg
KuwqiEgmlMYL2SjReoXsZ6GoprficsLMkogJNXtFWrve7gwomYYx/h4eQPulh8d9
f5KE67YXPApHyFSB1+CuNO7f0Dme5QwfIheluaixd3bgFSzK5RzoBIN3qTtaFbBB
6OyFS0t4YMFrrTiHv3ogFFWnspP727SsghYtmyWZ1LNo3hS7ELwFbz5Nl/aMaRMV
MQfCKy/JtnOi3xKAnpbUYlq/pCc6A3aGoI7UMO9KRngXTaWnKvKqy/teVMW5EzNG
83dndkotJgl2s1vtmaYztrEPq8ES3e3e8xQq4rrByyahC5ZN5YfyXp8F48o9MZKw
T2f4asS+xF+x7EPUHUZ+fwIDx5/dgopgbTICtLPtOtE7eWpnc+PhNpKGSrptFFdG
40qed29Sedg5WnJ5NV4FKVJGZ0FzWHp1jXRo/Gh2Sgs9hvOnjUE9eicouP0jq/H+
TmkehEo5qV+Ut9wamo2yLOS/usOLou/C39nT9cSOQtSG95H7TzfCrJxPd6VfYZ+S
pD0/Mf/015tO2Ej9Dy7xowz1Tdv7effFeNTB1nsdcwAEKDAjCFlYcejR3TU07Fv8
gqWoPXoamkwaAQxqWhWYc+WBW/9mMkmsqC12T3hygpovWWDyhR9W7tM+IIKM24Iq
Ir+Nv3gq/8b0LtCfBHzmzaBUi7oiNgSBwNTjTkdOsVsOtCz5EwgGWPMD4TiNW9Nw
8g95X6W3Ssok3q8CGlW0vl9LcIPyM5T+96xnInCwIdHfWO53LWcrAgOoCKP2g2jc
J6Ez4e8EMpEO0JKqpdBxxjuZ2Q9GgpdwTDjuFPgtdeK/YLZo+AMD33vL7uTJ1M/x
ZUonjvaFvSLBSfDfRYXgxSaad3rV7IliaxWAYHQA1quJ7/1aC3Rr6Cm1O0TrNC3S
uy+oWGeYIpWYErPTf9POQaggchwoCFrZAH3sSbbFLN5PKgliJr/fKNNdMBYljcOS
6ONaLWaHXtrbt6Q31qPgcJ3vCW4IP0Tqt6O0fQvlSnQ/on+J9DxjeiKZpCC3kgEI
kxdYmD0KhQseVWm4BjS1wo8nUjsFGPvNXrVqwcmG0G7LHr70qRjm4ks0NS8VQyYP
CddAFbt9Nj9w4AvxzsUCTHrNZqw8DSVsHyNT29EQFK/oS356FHQfmhOdlxGHDbX1
oTCFgO/aaKLeFrBUbUf+8OEVtGV7k9xZszsxqhxg7iUrnvhmRFkmxBCBd1+1/qAa
/KvSzlJ6WQ40T5Wa5X0b3yz/5n2mr0uxfCj7SBMAiv54aXlnYFcs20sI4NVveuvB
Cmcqv3nlJcnOUjIpV0ZcXw3uLaf4Qb02+EyvopfUwWwY+cyniY6gKZJfI06AwGcr
YDk8CL0TWLNdxzh9g47QXoMzu+3nDlflulQ0pt7tfIbW/7Se3qSKlcxEbuKKYw/a
rzach1em9rWQCLQ4jJofDZCu6Ld/zc3EiEDxjbNpOWu3b1F9NtP55wWnn8kBWmdP
09IqMk4kp9onZSMcmgquIfMR69NZuNxe8CkLrIIQI3yGC2jRBvwruDEh1rFSGrh2
kSZrpANklRdgaSkqp2SqkGIv5EZc2WFroRhdWIUJ2tlwfTlbknmmmUQtz3JWRDXc
5lx/tePzIjR6zVW1j5G0lFlp3cjOkOL0BR0IfoPEkYt69shrmPIqZLwrXXd1mLLT
eS/PgcMOTUevfvM0wHnmT56nG3fAn7HnpQhZLY/2cfO92gHac1ob2DF+BE46eaSf
M1IgVi98mdadb9ccTQ/Jpzp7aUruf2lLzvwRd0RCZvF2+VNMhYbQz4ZiTzEHk9hX
AhlUPAhSolXZMw1gI0tQCT7KbjORbNVJNDjpbbJ17BFWwpbhH9ZH4568VFE/X4Oq
4EVrqvRb7oLcuGQHTvklJUGWQwiRZautKrKE6fDyww+92VCXpYDYTi7pYd2wZZuh
9xD3Gdz0afcbm7VhIV3+ifZCvAeA2y/47pLuGwFbSmHuTYC6DHer+irKwkR/h1UX
CPBC2bGbUxtvKYn+DR+mW1opnagj4V8w4IZKgbYv10ZSnbKj6SzQSSl7tu/acxOA
Xv2zK9j9bWfhpk3Mc7Aof6cyfKLyYmdSAi7OYNM9mLEeIshxc2XOSCoaEKtBGxal
teyDkZiGhh15RaOpfXYYB6egeFWFjc+ZHI4Ys53LO3m6bO1JsPClSFY1GgzOOe7N
m1ADP0q6XR2pVmjob6K2KHgTaBW037DhHTLMJBgxzBdPTTyG6lGhvUYg9uI7oMPb
v9XHBJL6ayUZQHXWZ2N+FFq7q46wDBxW5HDmy/4dFgr4Qy0yk9W6305VAxWNPCxg
NCudCtBY+L5kKHPrnmd9nFpHG2BKrP7STHEIKQr1BvAmPLNIy2bwLJqwMb0J9KG+
+A6UOGJ+h3Dm8J1IgpRWXm4Vbz9DUmzau93aYeLKzuEiK0ODnv/VTreISgMeXZMq
jVcvj0+Fn+PZEXI8KE4EU7EKVifsYl0iHFieJtQAqgbAX7NMsla5NOs7KJProp2b
fIc2++xRVzeWDxyB6+tzK61IMCXy2ez/mb97S2mpGMcA4qVNQ/euLqw2xY52i+YA
j0gM0tttDVcIWA09Qht4GXJKV4xol1eFermAKkaTgjJbZRrKlp8vv+gbUwI4kNqB
5j1VkjtLnsbOjEn1bPe33jFW2QzlY/S5CHaLw5SFMezUonFOWU8pkMVkfimKvE15
XIIw/zDRja2StWZJPL5OYRRo0hm3nHUQpZnacfpglr3mE6GHU+n6uk5fZAkpom0z
bw4R/4Ol5Cxu19P6i6iIXU+LoqI61b+7+P1zsGjPYICc7WdSaZCZsWdCKXplPrys
F5amF+QL7jk45pO7EjwUhTYgPbPdGJjRC2CWGGfsDgPPsZE7ITBwNvloK/MbywoD
UmPwuLuOg4TtTirC7aD8ldoQRczPne3oyrkyjoD2alFgEdA0qIrbEsoYMcb8uFq6
6nPqVLsd9mgXvQ6Rdy7v+UQp23VfEFP6BxSw4vgdV2ZyF+bIxFTy23G776TnFPx3
YgeCCzLLzsKnEJhGGlIw8A4l9XI4aR6RsijiYXat/l7QukGwYIwb172iV4Z44ZZ8
xmkdWfgEPE9gWkRxg7+1Bc60BZmBpxUa0CeIHFpimnwocfQ20mUQLe/Qn0GRMGat
1PRDcNdFKHs/xozLU1VDMv5zvncYeBkgNGkLoazITH+XxCco7IpE1tqW0TVkC/fj
QxFmkvV1GpBUBiWjkGH5VwE5aSiNLxgwD0G++ExJ+1obpKU8KIwwAX7Qzvezani7
QbrKT02HkUhmaSlR4ikjS3QnyXJj7p5QEuEWoGhV7h+zzGDqszz5Xe07WsXPJbra
iT4RnysFPH5qqhmylw/0wP+jbr/dEFmYytcIUru0pCMUN9hLnbXeDcRB9INCVA90
l35EaQ4N9wfQZlJFvo/a2PFbtYMmkRN+94M7vk14Dfeg07ELZWQP/5CC4Z01Qj/N
/9nNMJeiDAUvVRl4UG9yManARtpT6wiMb0ANsVK+iFOiDtc2BWKvU8h+tAqNToN1
3FSOC1wKgapeIN0npZeY3UGBm0ldtevP7xIuBdxYTHvSaqZFhEG6XD4TusTsNiJY
rKL/8YH1Y8ow3/2QgCnn7rSngBmMUZhLPfD8V7MjEl1ap3UYDyXxfoAn4h1QfiFp
GsdGwCz9l+H3VLYPM+ClitKSC2Df/s6DPUztSdI/nYXk+2K6YVXBLxkTjWmwM6GX
LQGBV1GGNpsJwSzmXIU8quwpPmU6iyX7qGIxkfBObQPxd0FguqYyfMIlGBZhQeKS
ecVIUGvDYEGN/wHquX7EqZ58QYSeWocV5F//z8TW3OPw7m3FizzbSZW+V768P3u4
ZSqs4p0sfBFcmhSBxw2QuJSVxZ6RSF6N/xi/EKnr+dkujS2BpaAXwugwsbYb18Rd
/ldEmac5Ix2GqaK4gs5DVnyggqI4vpaTRWgnhSaaWLf69F3zIsvqBlxNOOMbatsf
2QduGiBXhfbw5t55R8JgjkDTb++HZBZLbnyii+TVaRoAlVcU4YXDPVoGk6vO3meB
jUV3XuvJWCLphIaZgsqbcGjqsEBHbU6Baxqf6Y1czHlPeAfTueKaZX0k0JGpOIu5
v1hh93BHce68d1XYk0mcViqKwBDYElnbSQutczJJrYyfFPAttFGNLJrKMuR2bQhr
4MzQpEtbsILWyB0PToEPgEE55X6Yp1r2EeDC1LwclKxPLxzy2TjtKKiP1Q32eXGJ
HIpW3uLbHUZfmPTZUJ2Ztfqmf45QiRDZsoXgHcggVpD454T6ugEHgEjTe9i33Uk7
sY3Sel6VYyWXDWVxVxL9w7rqXzdnK1066wWTxjHwBRV6tVFti1mGAWvyhaMTumF4
2XW8++7YfyMn+l2gtrpvRYDKzM4rUlJ/sVioSxGc8/KZtJGOO3entjT1u7NKNF2+
icuuE6+kRysAglukYSxUd5VkZAfbRhXUoiCh0588S2IIKqxbzvoLWF1kavXm8vkG
ChQqMLsA7cU/+Z844EAyMc86POJ9MbwnmBH02HXC77/xocDkFXqnE808iRN52Mig
+1tDSvH7AtnOM7a93cytqC801VADxoyncTSdLYsd8xUMW1jwG3jRgwJN2y5vNtlh
7yq9oJyB84LV1aFs3imBpKMC75M2aojbRQtUdhyinVlIzHG3VopWuK0DPi49/uqz
xgF//IHYyUBRWcVs3/398gZfCyWGliKBcBETQ8WA7hpB7cNFNzxnI1F3HPuHdzYb
5kY4Gf9B4qNiGrZsdJZqqrYiSXMqZPY6WyNrhZrpqr/v3rhGIC1rKNSOQLmv1fWu
m2fH/CmPGKkFC6tq4XXJ6fe4vB/tzdY/cqZHcEIXqOni9+JzS5hvCFHRNNyDl8F3
y8S0ua50jjwcoGIxKZdjX/zcYgbgwzKW1Y8KeUF8jts+NTIgezfM+aCypPRs6U9W
N+YTSQ7iPYYxh9orBZCx6Iv1/JwM9jmKDY8cMd8fHSKg1gIlKoKP+lt6QGcefpUN
9amxG09HdGSZ0R7iteOwiEC88nc6rWKgKYJCA4ucIzVcGwmHXAnkZZTJdBEwXuBn
yPBG7MC1rCEitMcKpW6FfFJLBdFVRsFMjQGxBKpV//psKD21porIbAx4kzOWpyVo
1PWNgAtLMGgwol3QIS3X18LUtVosfLQf3r+8yrTG+Po7hdNjzqm5uFyt80kqwgN3
dvJRdSKp/MIXrNn9JRyE0Gpr/OtFjktd9/aq9aDXQhlOK4IvTuX/uOO3uce6P8pR
GKxvBJdx72wTvk/HLoyYTAL+eY3aCKYQzwVOoHLxl97CpSAX4EpeV4DdaAN39ylc
VdtzJnk28oTrEY5V57B9MTckijnXmpcMR03qwaG6TDtcEGEpCQ+um8eei6PKr9WS
7UpOx2uJJX5mhwxnXuilJuiLtSo7swdn2f/32p9p5ku7XaT8Q5vree/8nvVuWnlr
HsIfg+dhi7nwvFPULjvgY7fYjmnAyCrjgps3odbyYD7s++lMOhmZSPQXYeFrM4Xh
ggyOJEVAYqhojOm2JqlGksgE63jHZqpTNdv/Njk8SfSoohgosq8zRtpbAwiM2D23
p+mB4l3htrKm7zl5FGnhql05fM8ECLDYD0KCRs4ZytwnhO8NO2ZxIYKGbjbGZtBB
WzGljeGW9mxB8B+ZPkG3JY8dolaD5y/fk2glBZigPof/O75xmi6//rhxvADzZnBn
WuGtqgSMpl1VLKlNhPlrYlqqb3WnuHM5nT9w2/a4/5e7u5KAlEBAaD2gX++FpGUQ
vqEsnlJ8jdE3g/8nHeTx75j98ARokTIPe5L131DGZK3EPszetfGpLE8oZjVtparb
ix1u9tfADWLBKW34GFJPE1WdiRPMMz/ZcNi6tR2V9v1KH23wNU27KI2CI+8Ec6yj
y7engGC2qZPCcLFxKj9D/L0rlrM4EoiIebHXUXyYMzX6DOY+OdtlGtKfq2/sGm1+
AqCRQW0rSmZ1ZNy/sK86mgTrDUgN8PH83jwSdk0vzmmae2eCRYZoEz4p6GGP37m1
LSQo4+j4n0qL3eH0dbRD6AA3t0te5oMzZVxVVdqmO7mnDd39+w77wt/KnbKEC3uK
Cg/05AMmi+jTdAYFTuoLBrZyVRkLQFT94LuKuzdwCiLOw5EBf3oe/ZP2DL6sKZfm
fTgf31N+BEc/uHRzb2BlHtyVuhdHQQa+WDuO89nd6Z+iHV2ANvPcXNLAgecuNx4a
PV7W0tuhRI+gwsm3jBNgzs9gEYgOqW5e/4Rgw9B2iCzc6h5z3SCPyLmh/JwGF7Z9
cv+Kc5XGFIMIxQLkeQH3PEXBi1bo92s0q2rakZi84V1UT4689pc8T2Slo1a8MUQp
8IB8+DAB5hljRVv9N3/MX3SFan4pGOcBqMyRReAiyztWcHQIt2RrnIihszoYirfF
1Rnc4IW+/VuDm1yRYa2L0yg/skWKlIB+dYRKd3PW2z9EINDrylKOFwe+Pq0U8OFg
E/ggr1vzjqfL2bURiMakVSW0zFsxVUi/YYF1bEwJzh2HkjTnVEv1xepYk0W7pcRf
4Ehb3TnX/tzcyJsZwvcVwwlrBsXYuuF9eOHy5suqfTHbbDhQaxV/FhC0chhJYW/M
pKgDWzqbWo26z0gG/Tv4Fdi04jaS18UAC/8n/vkIUgeyhjOIBOqFSBPFo0KEDdO7
DbFQu1hBpKbUvBmrqPP4RiV05bEyQMgU6wQO2h4tBAylsKH07hF9dnuAT3MACzmw
lOZXXDUR8wgZgByAX1Z9oV6G32Dhavzv/qcqyD5HVNnvlooXaUko75xD/GD//xc5
0ZFOZHIcXUCIkUVax4jnwApb3zvx3ntplM3t8iAES+dcMrV2bhCJy5/UI9ajMgKi
0Iwft/+LRryXfZfWZSX6NWMEyYD6FDfspDYeM0X6ppXEWgCNaI9p5HmTKnPMcnJm
D8lBcxxeCJFJWjiM0NdI3Bd4zi1IQCo/YzuQWGGEllv24dTGfTPQcNHJ21itRjAB
Cxren068jj/OeN8cJ1IF4aXljLBufmTHC2bvFIoTkfLaMHmQ9S6m13l7gSMmTjNI
bHzQcpF5VhcK5xIAeHxjiynEy6fccFCbQ1HsT8zuh8SEmPyRmTdAAvGw3YCF3VBV
8+RVfc2saiMdNBrqfQw9hzq0scO0XA3fuB67C4T9+FNzsM1T9GUqtdPAjmBDPCXu
unMf/uxFl+XymSlX5fWV+YGkj/N4pREggMCiNrXSs/9p7HiN1nPmrF5vrkMRBqdf
q7IafxDyrFUcXikk+En3h3HQgDS2R7eQFqQTI4vOg9uBUSyZGrkPBd2hdptlZTlW
0avtKhiBczHm8GyNQtRX6qTg1MTRrTbSs1uzcwDYyMMESwcPjPIETg0nDUmpN6OT
mlgtecQSVrZRMx4vtEHGsUmhPv6Jau9gijG6WoZgFj/xxARFP3wkAMdO06XLyUiT
SsvGCbq+iVPe6acU0eTagGIGL4XhCMa7Rbk4Vz2YXIEhpoF4c2F3hcJo1xRQFwaw
ekjru4aqBFE0QVJl/Z2eZE2HyWwklkKgNicUS4a7Td2K4bpE+lS2PsVNdANbRlXC
EbniiUNPlScNeEGXQDI40cLN7TyxCDQZQC07GLnuUUtuqvWvHdH8RQL77qeTmqQi
KuGeua5CLDacb5P8AF4CWDqV5/e8S0iaH+PgnrECJunTdKOJF3LzYG3G2SkM+h+d
npi+NilzDjM/8neN3MVLNQEtFK7NPb+7u7iK14Iz8hcNNba8p+5B70wiRQY9/2qE
0Ui9AtxbX8a0HSxVEXX3+vdLAwiG5RWYiFxHNqteJIGUijar+K29rTpy7DJQz1ls
Py9J3wu3eCFkaQhymfu+GZF1Gzo4mvLrwvUpNZhvxk2uqHO9NlBc2hbzqE9mH68B
dh5Ht6mpwnnPsNqnXwLbEoGlXG3hpIi6PxAlR7vfxMK4mD5izNWPKL/ubeUK6VXM
jhtcw85rstIjhZKFkJ+Z5hUAiF42dXXpTx23BbdrIafSpyXcsPrRcHqWF2pukVZS
8XBezsiDG7l5pQ2u9cnohC7z7a5O3Y+uH4yicSRffa5bHOZ1xzrcx+s3ck5KapwY
cklJM3LmAWId5eHGirDPm57/PxLODlj9aoACCqGbC96tdDdSO8u48h4AYrL90C4W
C9OC+kWUMwgnQJiyxmxW34bRjE61MaxhIt7Y+qgySd0RoXFS/WbPjP0zlmHXISpD
qmQ3+HRbBMfIXGsdOAfiq/hPgEE/VrPBTUpKIl94/DrlejqdTxij3V53sXQAD/fy
tVN4N4it7fSIeRirLAcy3DJd71gjwRitFUNaIoqKbNeps42xd4yxPcVOwu1xkhoC
AlnnctjVRiQQCCBOlakTt0ZDpjzFxCbh03V87Z80qvYo/0oBAuPtQQqGzQVLOF1U
DzfiANs47ahcf22QiBRZPpBcPLLw+bX8jJaMsX8TBh5HgS2bwichiwlxf6+8qvTj
0PFy8yO0IMzZ5gyQ9C/EQMFFnWXrksvrQgTes4PNQqUND8R6daxVCFpRk6CJI/fV
itFKQKhK7crFqlRJfmPE90oCByzOP6MGONdVU4T4wcY7I6YQdhdqsPfBljd+Wlvn
AdG7+G4lA9w2I7a4oNE3RoTKP8OWUxGICwt5rHb7aZhx6CkFO4tyPIi25XPdC9mB
6jKD/sG+94ztVCiwGoOp4M2wTSALiPY0C2U7CPT2TZjKTgIPGkvbU5cY7VoYm2sH
/XAyR/Rfv/j6rTGH+XHSPR0TcCAPNQ4VDS9U869sWdv4uoRdsK94lFFtjehngtj9
J5d9GB7YZtczixcgDUD+XcJaZCyAc5LvkQYGRqWLpJubNX5MQ5XrMjUi3FtpMvxS
t1dFG1lmgauu1Cfy790Y51T/WCW9XE46dTtL07vrWt/vpSi/0KSrG3srMhcxuxO9
cA3Cid23Xl71ME7TUHUCCUXG8dvT5911AokOarxK6gKV62zDvlCbLAB9hi/Uk4DY
5aSZNdlx6uZ8VSAxCyzmmGz3BFuw8M+IuVvTvpPBLod6woTwBkKlsRgq9YKyqwsB
9An3vbaaSBsUS0eEPHlR0PiCF8P/jQ8GaF4w5/P5f3ilaCNsxM3ECVkoqh45PyGk
zAmlHy70M8RrQMD85cYT4tqdpcCCp1b7F2QBR25xb7+y2qhAjTtFzkWm0bjIHOAK
gawevrU22D14V2xzAgOvWC1P8OCjLVVVpXMsBLbivmxWJmfAm+6hfe1BGdVw9EeK
bx0eVWvN3FdAAr3F3F84ZiGJKokBDaFwLoZ3EP2o6DMArtXZvz0BByca6a1jIWGB
fdPwJoKOzxuf37jReknP9i+y8pYbu8qgGdSFFtMipUKMiatctBidAqVkundPnUrj
blCtqqxO3SPc8DLpnhn3S7NIJ74GT9EMUi+OwgxP9RvZCU2uVScmzmCqIs+tj+ZR
QY0v5lNlaWT4n0ykmCzjnS6d3MekCd1YuUV+XsHIGoOhlp6pt3AHfhyI8eww5iWd
vC22UtfP4z7aeCawm0vWfVzpfOyEtf1pKFgXfKdd4RRHn4AW6Pp4K+xgnmqlbsUf
/t72d5ZCVXDG5l/mCodWuk6S+mhyqHilTRlk0a3m1I81A9bkr+cIE9xfM4A3zrw+
zLKxoe4vOG0IqjZULnU/xOH7XXKPxj8MagSzyZbwk7sVKPpHe56JHPuaN5TJoC8K
R2O3Fj0Rb4Z5KR4nf0mHHPf2G0C+oIJVVQXzTdfDu2hNv9YIZ4pJPWXgTR7xK6eB
0E9LHXHDaBmyuJT34Sz+KOMIl6igXobwPnxdsjm6KI8/NswMjiHMQD+l/u0ELND1
CAvaTHSdGT4oTl2H+fW+VNg0RxosxYlHzU0NbfELg5ZlVZ2l9E7Hp1ppXeRJIgye
dEHvchuSvrLbtOHx8CmYGArrw7RWwqj3G1yF/CekIJ/akSTZ5rDCSZX1zMdrK4Tr
/tl50FrXHg4Oy1zOEzLQUVWKWSShWzCRUsW5cWBZvud0WXE9kNo/GggpA5dueRGJ
8l20uYPTXvYtb4Ue/y94M9KQ4YjT2kydN7iqijbs0cZngbuGrhFpXedf0ubX3d9T
l6s2k8FPGoMM+PnRyAVJj3MryNXzTjzrxaijmAvwQSGI72MquCof1VUp58CTKRM1
R0NX0KMBLau6ka+0D6V6f9rCuYb6fHRtNuh1r1dwE+yI74ad9WY21azB+c43kfT5
fM6aMc+5jR0ut4MHjU2h2nyVxUCZUkCw0DJcZwu0vyMPMHXbY0/CKf8nYeaXYSxD
rOWtfP70Gl3yWuO/m01SRftXF4vBw9jvBV0eFWJbk7yDkfVOGrtoz8IabHEXkWhR
GA21czJqkZi9trdnFYicsb9D/btb6tC11Xc/GlXIyqtsniM0kY9zAUAcUHVb1UEs
kAPD8QC9oGCx5Q87VgVkbdahCM4W1gr3v5AnY/gSCVdsebeDB28E81qg88XIbbcq
f0cB5//N7x+82np1fZt4utYTmqKv4ywJWM0sf26Fzm+Hw1DG12Xo2p5FoQFiaB8D
4WDgq37AtzX7+sSNNiaFLKRL44SlPPqZEQpCQKBipwvnSwuSPmAUKdg/Gvx9jit8
axBBk+nth0CymQPDmjJd/tGjFrYt1COUTe7roqv/kZeMf48M+Gg2HuGNcaphD6ri
+qghGnT85UbRbVVSCAQ7gtKRHkA+ce2fWBol8Ms0Kgxrh5BA6ZwRAny8q71TBO/v
Yh0HfSh4pKCNm44v/8RRRmZNsMw2mRy6FhcisE7rXUrHsVyZcI2ot3nWZzqVcsot
3n/LnckB5FlirlVnctWUu0cGf1ccBOi0F1beLs0fFx+jp2V9IFwlRWasuQFPDS2z
NWt/8VU8yJoJ3BAJ3EypvbZx6u7HlQZsLm/mb0kaA9elTLuCHC1+y3alce+vC8zs
/DyJwQUbZ8zrbcoy38Bp7YFSbjstWHJJnq7rA4DDAv2iR6snH8bfZIaURaGTjsSQ
3hSRoVxy/ULRGDfj0+r/NvbpSjshUIrzgG04xY+E5M7WjGvFHLMimhmoUHrUCr/e
DA2RhU/TojSkeJaDZ6qcSC/AP7o4HqHxByuSbRRxrAn3Vvd9E4U+BHJRIMXGJS99
lLhSvJU2ulO4vxRAmyBBVvVdpKvuV9ys0fX/qftnQPg6Rgde/g1rgbMsjuqtIZ9S
sOpB6twM96hwOUxZy0SLQNNFhzowyJ6IeSqgCfjpmb8QrVUrmr+Ed070J2VwrqxL
vKSIErAwR/P69iRM4FbEGSdKRkHczZuUcd1Xo/FTtIQLKBgWff6aEBouEe1KBNIh
0puQpPlzan14ypYfIjewaBrqqrRjIFJ8r3AmC/DvmdMlobZ9Gnx20U4icO93Zmw/
SmbRmF0hid+JOc8m2IloIv4q7kRiY8Dha3JCyncOSPcwZqP99L+2ilMBmf5Smf9d
01qy2LlQ6edX0DLB6ZmvUydG7qts5xOCd32Dam4LdwmS92ZIuZTTFfK3Zh2gaXsF
NCcWKTuqIml+j6PapNty3xbU6ZIClK4XhDSRvfsijzf0LfA9rugsE01avUnVVstV
Li5Hj6dfvalncrxWI/qF170FpCYUL/K5ufbiBz/IDNQBHMI0c/niSZrkbphLW1ss
Q8O/3yWMTYWrFnChgCkdsdmkiD8MCgy5IuXtOCzRz+MS4XZDiOp1ZCQv0jS0ToDL
/e6OnFHpmkHFyGWIjU8KkszadUZYaMxXeprL9lW97zUxa5A5w1QkWnLyXDmT4Nv8
vG8D2w35iL2Rc3bj96pkWQD2vWKNWMIIBNrGoc6/Pz8NMLlbn0MUZU5+l6ChRLEG
ZyoFM/GKlpGeGSAOXrogjxwkpI9AYl+3/pqclPetYn5f7IGzx1VSMf8erZFQ4Pqs
ALTAjLEMJh5N8DFnpal4HbnNsc/+Bj6XaYq1uTjGltTdAscBwCwyRuKYRSTmyJkT
OHuzFqkxzfSqspbCctZLSP49OhFnxnjxr0aRfqFy8CqKHUlJvyYV5Vh3uCAtezdJ
1l8xBIzKYC6rteChTPoyOzXHYE6Ef9reKFZ8V7GMl1QWOS/92BdOnsSQRHfpW+8Q
Bo14ddEkcQSw1VcW3D0KCRA6r/XN7tATqPWqV7U1tEnP2hb7ASKvXHMus9aC0Ha/
zNxRvTxUAINpBn9SBctVYaRlRnP0HHZnPTCU/tWCc0OjfppZ+yINIso+/r8apCwY
Lkml6R3uIxmPyOOcCxb7o1mo/2MB3uQwS6M31i32RnBM6P9K9unjbOA6dL3j9TtU
BD/D2I1QaOeEmYQT/DzQvsJa5cXG5ABfK1g3o8S32n6BAKOKQPvpDLNlK+FU2cJT
ynRrPEEUnWRDdU/2WEIhKeL8OEw3sLJoflC27o+ffA1pEUezCIZkppCWe67xLreX
Rsg8kamMHcG187qyDUHMl5lOCQohYXOC5oxJVwYI/7kx5EZf0sOic7VIIEo2o8mI
VP621hh7HxMrAR6FIufX6KYHqtjjshEY61JJb6J6bqpMZ70tJZrXdOjnT4/0wquL
vqQ3zoK2iWS1yLc6r5Ay1+Nadi8vU7pAlE5rEjAraJopo9P+nvZPKkAkDl4vt5hK
OsUPTzQWiV6IyScFLcawWy8q46qb/bQSfMgH+2w6QrRmkYz7mTd9nAOO4hI+Ph/s
UytjPXy520rLtRENfqlqK7XQoDfDBRYP0eFtSvdpWQlPRXGLF9ctsBN4nCkTZbid
S+A4/IVu5ct2xdK5DKrLFUPr1BNuNO5z/XObMc5tk+Tyy/DatWw1pQGQts8Iz6FW
WtlQ2GohOtd+PshHfwbpaOwo9bxZx66CxD6uMxHZIlDslXd5yxsntK8Wpnoqote9
mzn2E9yLlhfBLJF1SH1v87QkgMHPf71kwIGY8eVapEB6DatXjReE7ZaEt9fTl04f
Bvd6csJdPK4VMChErBU4HGMpN0mMB5725HaR8YWnbi3hsudRZgPFTEM4yZjgKJE8
9lpK8vVNAaWFY77mfVeIjFwZgrngLpqrPlqrip/HNz7zIihjjsUZsMma3x5GIg7x
sBu2cX1GbFs2azgK/8ab0mnz3gAg8gApsX9nk2CiLcEmET5eOvzIbeeMr7tafM6u
ijVxYPHLmjTjYlph9dlkDyoypm15bp8ddMwgqLJ19nEn0k7i6B8F+rymujrg6MVE
m06dN1h8YKqpSgBXbdT+6a4ri1VtL4kg5XvYfDa2RmBfBRXUk06UGdH7zNAbokk6
N6EbDMmOwwX1jC8m8i6b5Wx5a62pM4it9Aa2Ppm2hjgTJNKfdLLwwViFqppayrZq
CtrlPauFFdOcLapMp8/zs9iEUt6oyuv99ZwCavd6pDepEyfp17Pcq6yK7J+3s3iO
5r/8gAlJvkVM1ilapL0s3Vytparml1c2mWZEj0Ls0PIEbIt7UhRipHcQPghpbMfF
7lJm003l5yztTbDBI2jdJgNJ6Rwx6yFjLWRlPXmaWLPPkjJ18hBeB8uzdkMwqYeN
vzjxKXsJEt2NpEqsAkrHvOGumAj75Nt6670uFOTkN9f0jKMcsQnhp9gd6ULV9xb+
4HfBZkXB4nBtosa+Mo62KyOc6yrlrIURbPI8vOvNwOa5Rqm8mwJfpsdBLWsyEbo+
VhjrI5y3uUd/bk79p3HYn9Bok7l4aqar39hE8mxKzwqH2rl5jac3r3kU8QNHnOnZ
X6p/LsKp4in+NjI6Z7LwiXAfn3l+OAXaFueS+zHwU4vR9bTK7lt3GHR0xlBmyrm6
l0Ee/v7Z623uiUgjuzZkyKn/r/5vtXhA9Xcn6LVvPUMCwvU/bcXpPpTf6POsJbHz
p6mvmlD6SJg2XOB+NXD2SG1Wk+W9GyMQ5lrmsuvpUM5RBW3vT2kdeeET0JYRFy3S
hEUK5zT2o+VdGRwVZq1nU33ZD9bJhthftyo/XLE7lTM/6EYH5xVzBc0+EPrPqWYu
8ED4w0aoraI3PIkzhR+6IyiNkPTDb3mXAGScDwj+zM6Lnl8zqm3j0Ml69k5a5Le3
T61QQgipoRQG2h3L7gT1xS93D6VrrbsNejxtF5XYmrchTC7iHxEubtN1DXRM1Ttc
lABWrF2qHhYc8XDIL6unurkIOg3lx2k420b2ZDb2DvoNoxKDfMqRbxDDnhQ3QKSq
lz9GAwfGzo4miB8H/CjNp0o+5v+U7OVwTI5k0gYtenagrXMgt5W4wv6dfpNEzDHG
YkOipdRT+tzBZE3HOcusLSH2rI6POpww9h8t/M70mS0wIcHzz2bzA7WXr8GgxDo9
4Prk3cvyYfcYNG6As9WLKTAE4PmU2mJNToMh92ym8cGmZH3kDLzm7QuPaLVz3c2K
tYAmpTN5xP7/C76XtD0k87MgptKy/4SYHUtpfDFGe0QwLt/8ilHWScLXWi3giiIF
KMkoIHgNP3AXORx9A9wCRGDXpBT8JZkwB5amq+k3E69bS6UDNQ6fvH5sj5DDoGR0
hDK2Fl1H8md3JC3Wrl1jtfIm0hxgnBszIpdYOxwQpFY4AEtC403mxczWe2Ry0Oxs
5OcdRIgG7tOecITQRuevCc68hBbfbedAsVuz+L1+13FWwkc7hWmN93VAdc+xpJpm
hRpOLUIXPqXwIm+CWPtaZ39l/1GhaW/3eH9erUDV8Ni96jBkDPjdWulpr/jm2iXd
rgSqPqqQmcokWznAj6wxVhxjVVP9tzWTvtt0PNDL5E4Fn53tqeQNzYILDJ8MrYpr
ScpWk9GtdmWDX5PQ4QhFLs4lWPMUUC+AFq9PC9naLOovEjt2XEcy83Onvofhpdlw
wMz28wMkKJkqkbclvFIzcZOEOyHUso9iD7M23K5h+yx4cvBQwlIfzU1Q5L8viMel
FRVTkP+NZzxz7eAEXyTogy8CmepDlS9CgkAG6Mts4K9DnsvhSALHcQn+NaGXPtlU
XsNeePOzYpbE5YiPQeCYYDqvpWqa6ZMgrSKxg4x68a1ZCZrELdJ4IbinGmzCMFnK
bzFyd/k01uCSNIgmiiPW7uRZCpu+Z1b7NsT5kkwn8PzgO3A83kfce2LCkehADr8h
W5oErjCLtwOs3W32zzqOOTETR6VOX1c1hL1KrNDMgnKeNqeOhAT7IMtHqAaVi/3F
YQ5GarbALZBStGrPxR5blfgHKfe48HuP1FcvFqbi8x5h2gZZzMinF4cOyVpLgvcz
EBr7vw2lIQquybnccSATNlmc811rA90WXWbOj9ZrCeFPzImeV6JdiynCQlmH+GR0
w2RVeOrvl/FKfBDro7nuY6qLkjseXKzgXJv7eJQ0RgfMK/RbtRnNpKy777PBO+vw
V+sjkQDGPd+BmUYTC1GOXObsseJp4lJMG5+W+w8z7chO32IK8c5ILSBiqMXGdeFD
FYsZBobICJ/LKpyfw2cz+cAkZ9T0nDC5kK3uYHMocSZa0R8oGHkjntGJaCE2brU8
UWLtL+vKH0+RnzJHR7sG9uM2RbzfpLE38fsAB0mqWHBziAMSsYCrLuEvgb55GR6B
3kfYxZucJDwuRmuFxjwrYNqrxRiU6u+6xqiS4APYt5EJ+wBjyObMzz+yo5DNuomK
xveQ+pL8DcTsc2GXgREU6FnBur6h6Oy63fmv4SB/kINApj9zUW+jvW5SR0GyUOHG
WG3cOuMflysZQsZDN+lxxj2Q1dc6wMBm1LYwW2NgoBAKULeyp+X/+j+qm2aKtfKG
2cqd9AwgnyWl6yAiKoF+vzKbEjMTBW1ZHoPa139v8Vh03BAUZmqEN8FwGlcT+rwB
i+OME52OcmcVUKiqVa4duQosl3xjNBKF5IoW3g1rBPl2KUtyX2s/omL8zyimrCjz
p801dT24DEV2R0slb+fkrduF9qNTjEtZhpd5D6ld4FNayFB6VJIGcCoB3pCkM2kv
r9bcHehdlb2iJKFpu4tFkFFUhZNRGe2eE5GUS6SLCI5xjDavLE2YKLd4GsJGgTd8
X2Fpc5XfXF6OTxOBavPj4kvq4Q8cuIcD9ut35EQk6XEUhISHhAG3/rWCxRqsLr6M
bb58Yyk7+FZRynZr+vbf6sweO+xD4Z6U84oZtWkFl8EbhET/a5EVVfp2gJ3LlIl+
iDD23I+PVzkV57Lvk8W3NDQ8eqGIj8nGYlggUBZ3VnCx0QPJxCER2VJDcdAjYwpK
vuB1DOGT3Jxfq7pEjL52GwEkU4h8pHs9vrdnKQJ3pkZQTLmBKOlj654443Ry/NJZ
xvfCg32Jv7PZhZNqY0I78CHFjG/zRLHa3ah7Zr/Fqt+4AA/yvlkSWTXVNARgZrAD
JA4mtimxovhje6L/uzv0T3YAzC5ng9SEsZzCE/kvAWYuAFEh4VB9IFdVW3tzj+Xa
hePhbok1kntQqRQbpamYgVWkC0A91mTRbEEpKSinjoL5RyjY2qPWeCA4QRWX5cdJ
fOx2qWa904Qc/LoxI7ebKvvR2Lf1Lxao1UsDLQEumP8iZhDxGdT1BvxvzMLCllki
Xo9dVpkogSuIOwpblZvHVEulb7crgXjYcZEcGZF2srhrtQdF2aT1vXvDbCrrk6WV
5aXOV6IIF82rWrrmtbBuRehbVaVzg7UGh72WBgjthamXMWE5ArQBprvYPDw14/w/
VYzdMpNkyiE+ta5ZzpRkPjpMCyZkWSlCZQhhgTGlbgwvtEti+HKfj0xDgfXh75Kh
N01G3+rfmwuXucDOT+VZoZy/loS/exP2pgjg/xvAza6WwbRz29Ea5gdtBM8DIa0n
Az6mKTOFH805HGLEImi8ZVp4hBqODP78XI2WHupSC5o/GDba63S3YbNG39wHZN89
2pUzM1fXPocA/qM1jH2KfqxlFmLkuJeER3sK2VMtW8i6Lli4XVhFnjpYat2O3Of5
8m1yWR5efYsX1cW49FuXhfVS+K+klxpoRENr6X3qk/XGzzUdeRYO3x/ZYKLFiaon
tlrEGMoN4IxZUyffrjQ1N0gkAP97JQ7DvbShwVSWFStpQIbzh1qpeFp4JpY96CGi
VqlcnFWrGYMxReV3mvgbXL31fBut2BkgjwzbIhPvNiPNNCpS9z9zwjmdOvxH+wkq
/PobqnZwviV3nQOYvLZTXFhmwxCR2chmfbvDBGbl402d76e4udA7PcdE/SU7jOyf
TzxZGCMdcqOIIfaymLGdjumqqOm7W0ObuWPopJ9gbHhbh9UxXpAqBtE10QZ3EQGJ
jJjAA8AZD52xjAsqXdW35VdXzqTFmC5AgyTakKzYr6caH9eRWx1RxQbMn7PXKdw4
wwW2V6EcqhRV2SQgCzN/rDeVleGk94jetEYobPD1xZ4sGxdrrA8y98swE97rtcy/
4VACHDcnm3Zy6y0Nxvc8M/4lZ5g0NNkHYKFz7uSRcEBy1amssQ/bY6FoWCjXzYCw
VCHBBuVgiVUK36uFe+UQyO1WzXu7v89dfh8knmqmPA6SHgxJQpSGEjIs4p7vKGSv
GdtudttWHaRde9HodzAtrCtzeZqtfLY/Pmnk0UbnWHxXkXZCy4eaCK/ssoQpdAXI
ut92lnhSjL4d7wLhCnnfqXj7mkSNc0lKAJ4xfba2hmC+W4Blw0oean2coWScIp70
YWhVABSrbtuMFr0vAOY4Xbd5HQkxc7rFDlFQUwypPbA0996OK00J5OpEZ0mbk9B+
i48u5VQT/zoYGrJxd54NKMEQo0fB/nrNqCuHXbSKFHU7pdaJzREeuL4eDRPLFpJ8
pBH5vtwOoFl9pHBEy5yfD/AeI0+aDuNkRWVRrSm/pdcLlEOa1UBQ3X9wMtlod/wm
zj93GfPMSooSt7DH8EZSRPlwTnlIq5aBEKe6M3b3B/3+7Rix673/g9l7+cxEjNpE
CDwrz8YBzp98w2NaNbwcg7N2hi8eQ4EaZMzLFRUR4BzQgUblfqbtwHMMVMnjwxUc
jAPTMk3v5UOhdhBG+W3xFce1usTSUFpo4/fxUrp1F05etumz9vtmFAWZRnfx7+V1
4iK2fxxXJ6vl75FBYThe1lScJxsU9gLXWKmY0v094SN4OF6Lj7vif2qxV7xlA3d4
8GBWvbPq2rlWuG0zAKpSJnhfLyusvyFpelVIweozKk1yYEmlBJ09SLIHx+zKr8Ya
IhzgMBjFLoOBXbAdMZ2ucG7aU4NoLDE3KWGMuqn40eJpcDRjJRKKen6h3ishaPIh
swysRHIWlTLPif9KcGRZ5c0dGrTzF5ojXkGczR7bnGO/s4vY2sN5e9moxIpXY/+w
gjU47J6ID2HBcVPjAkNF22X7F+08TVAX/9MLKrKzWF94XFC+miWB5+ej/JzdP0Te
60XG2phdlt5M114QQihGsBmtgPmUUw4H8Oj7C71zT5fjBV8J2s+hBI6r4a23KhvQ
XplTnBa93iUirEh0hfAdAGf+qhs4TsbYSd8D8f6Pf0GdYx57XjwsLxW141LoCE+r
z0jOIA0X7C6wfgHvUxjSFRXNNVEbRAQtPBKNi6bGCqmYwJJG/eEZyB3/z8pdu2ZH
nOhlNY52sEaTOR1Vvx0Cg3ZXXL0/Ncecpi5XSHc4t+cYuWDytnWDuFwZLYyXjTXg
DrmTyhptt05xsTvKyhhI9+HMzVbBfHp6bXTLRZvugI64GIrruZL/gfQR7ZIzWlia
F3K7xRMPLkdZ1dJDrYd0pZ68x2knA2hMPiuCjZfCwbcwrgJnmamPyScVx8ZrVNPK
QjDUGHlxKedMLZelCoZZbT5bqw+Kzs0JFuUep+bjfhTqBDqI1LrlNGbcuCegtpD3
w/j7RyzSz18UD95p8GL06BaoyctSuEmwKHiy5XIKiWiTahvr0rgldhKQgKLI7D2i
3VBZDD5JQGw04OMJLY7uTmukwDBwZGuAOeszydESt6sO6wr8xV3O8vgemzxuY8UJ
45sdqI+7Y8eWkVdcFwEFsh1er8I5tyIv39w3ruh/CctUGsvyF+pRhFCCsoMU9QlF
Qo5ZO2a5qCPSqhvUh65g7RPbMz3QgWLNXOHjp17I1i03vdTeGAEa7dwigjxuQwSy
hgVSzDrSBWAc5Ohwdqsz0onNcp4wjVlN/TabqGsPMwX/ROLf2yK47+iPxv9TojBb
7LOupJVzQmMYnaUzA2dNNdDNdBCz3qbi8ZCjZ0uOuqbcPAEqkhHDtW5nCdfvvk8V
UCR7zZ4Qbzd1V9U2ZDEQLeGU3+3WRPFQORFgmq/B/SOGqmnvhmJxtc+oOAORlvFj
mq+f/ldJKawJG3HcZHJW0fWghoLSejWr2NioA5pPJC6s6nq0hAfWovYeEVzt2SVD
ewhEkw1GXKUpP2dHy720ymz4MU7gWljtlpEcdux9TOgBdX7CNajmHIPicDM/xxOM
qydbayZha92wdPpesN/8khxmb0pt6WdVmoON+nLVUy3U9EJO8MBfE/ieReDOniPw
P2t60IxDizjnOYZzRQB+hREmMb9S10Zs1zZsXb/+VfBF4oINBQVUMQDIok4RgfMd
eNVfLWElTz8Jb7v90WJaXbnQSZJ9jC2V8gGyKX0sDBz1G9T5T6eRVbiD8E/C2509
zJbNArOKlPV8ZQ9aWezXNfJZjhlMECBVnqPyyaYV9H3n70SKaf+AutSlT/+g2PL6
OyuvvfjR2Te0YgrmuJVij99ALNu3xbP39iXNsDd6mOjmsd/kidaZOQShdgpxjtAD
1xo0p5r7D2tTvEjFfti7MzPlaw/x8r22yxrZxquowbv8bE8DEnMqOmqAkvVkZ4gM
3eJ8MQ5PciDTrC/0GbNHMiNazlwR5SXCeyfYGzGftR8pZyBIXXbh2JykYYAdazb8
GjHf4ccdaODr6A77Cn/DnPeMml7c326LMx3x8EIPlUPaYDhqjGquhZh14Q0vE72E
kwmF62cjplJOWTfCtLlNUnX3CY6JsxoVf5KigVncHpTQWgSrnSo2K+XV1rG3ZsOa
4yQKXmgZV5CGWurLEMoBwKKQpfuzt7q5PbK2JHPxIgfToU3+qm8oX9SUGhN8qsly
KSStbUYd9vHIP2ex7UZrB1JAPolqA2A8LeloloLeB0ubk8uy5QWO0h4CxxsoOf73
IrbAS8yuGC45kMpK+2Sg/ktUV/Pa4uFYkuv99lrwQe5bzOpXfdzsQ+85IK9kojD7
BLghDODl+w5DqE+sfljaEog3nKHX0w3R/4xyxKoHT8Cy3eFGRwFjDd1YaycyiVU1
7Sjnk0ItlvrVhnA9VbAjIp2owJ3LrqkQgO/ndWmzcR1iLsduB3wt/Xs6YqI4IUDt
EVCn1xHiywp6ITFFivXJ3+H97ApFOj3UQTBQdC8RKqELCpoysJo4biML17sNsL7g
S/W58hWrm20U8ypBbJWlM/IqkZDbQekj7FzKeARmeZjFzEN8eoK6/nm/vahdvm2K
+86ZhyhQHu7lJgRzrMN9/Oc3O7XXAzoI/2foj3n9TexcxbVAXwiW/o0vTzxK4qlt
rEVSbgpw4FU8TLodMpqO+VHO3Ppl7w0HTrKrHtUdUUdh3oc66KfBYtXfY9F99aLM
LCC35+ZwaELKcSX3K13Jh7825+rJYkbsPKv3RfmrnxEnHhX5byagxyfO7uxpmZUp
SLFHFdgEDs8imcmnokzZHkQdro8tvOCq7Limm7BERv7FWTBZ2MbgCHynhUbqkkpO
SPUV+Yc5xpDOZqDLiZ8PgSeGzf3oPkfBA93myjKcx5zXHeqej8A1K3rhbaUWE5ao
2ecuwo2NyrN/m5O7/GE5jjeYA/QhjdsGU5bfBKQUdF5f93jHKekZcJiYtlKZMMQW
e/RxLWDhtBLoT+J7TzKYDpBpkvX3+YC4WVhJr6XQc3A/jCd3ceNGtuYlX0QW8QmR
sm63ZFKxz+WPiWamVDmXzGajIF2aqCXfA3cgFFIHWCwM1HbeiFKGcGM7WxqrItdL
1CWiGmVkn+E3RBDVmDCwwihSYOAfsIP/YjpWW6c0L3cMWDtlwPij2i/zIFs3WXOO
D3Pq47oPkYK4opg9dKW3UWRWuLY0TJjB24ni9m+xKCsyQfZuOM02cYLkfjwCeJGF
6xY+ngXm0nRl5DnW9XAAIGdntkU3OH9QTdHM+UnJ/EJw4JhIgMWkN5weq8nYHkFe
bjeV/wIok+JiMnr2fY4U61TVvNFnTUt8YNDmja19NKADwPPkK52VTlRs6IcAzzRH
WZ11RIXs0EDjchO0QTs0R35bpHZTm9ZCJX9M9kwrTWBLFS8cMIjjzyb38H91X7Lu
vcRZZZwHbC6/kf1XCh5r2ABeUklCUxFHZs5sXFy8e5cgEtkrcU3SCFVZ+iaSRb5w
hTA03XnUY3Y2S63Of7D0GizIh/m4w1or/snS/iCzsOrwbNk+RNp3XT7ou6ZwqV4z
DqPV7tfsmgTTDh6xSkgTI2d8o8djz6u1ix49XLzMnMgEB29lEdfb/x5UaIM4YnQv
lHPOYlZ0faOqtmir1SuXlN8P3T/iTYNKv2Aq1xHHRh+7QmvRI6wXc44okU+M3Fzg
QV6RNLDFrJ5Gkpf3Nf9542fLqpLhLiCuudDf3xFdYJ4+X8UmLHol416xpYKRb+K6
0qQx6jhASRGfdAMPRQh7U4/o9h1mHW7LFHIT0TvfKakB3SoknfpxlEjuTmco6fLW
5wHp9GPj9VssOHHORcJZoMjR+OpEodvSz3L+wePnwxinFbIg7h0mFKsUj5mTqUNF
kuFmk+lbJPjkFJHSEsjTeBaqUo/4qA9LJTzsBC8l03UV5g4aRjNXpVH5C/HgxtVC
d6UCqdZSKYNqvFzWKHjOdfHrPln/uuQSR2dqdovzLMuLB6LQo894S+7LpnVw9YSW
49/Xfly272Byg32qCpOj7/N0foAt1GHEywv2cL5UxQ2uZ5OITM5kZbaK2aIfDH9O
+LyGK+38k0x3z7EO93BJsBiCIwi7TXsVG2kJJgynNXXPZaihxh4Z5BF2zq1KV9oK
mu1X1byS9LP5LMT1waoZ2Diu3ox04ezL9Ewp6UHUYW8NLGbvPf1G42fClut46cJl
B4MrXm/qagYHrmEJ5VG57tQDKSIJU2DgktLpN3WeelB0KZEOfG85k46C0oIr2cY2
B8jh6CSNerToCPH50s+I1xoMyxkNl0CZhcxJoaLyDCp1oc9wk2Mx2kgr3pApJWyW
9dnbD0HD7IkDrcO3gMyZK3KgObMf3ItmcjU7n4v4DDWL5Fn+/Z5HgAFpxDXBLplz
vW0pQCCBdTyEAOG6s2GkhskqlwRDjM+WJSkMm6OBXRMb4+RcetD/jzKBcjsL8eM+
7Q1N68KF1ab+4Rxfi4RJbElYNFYjw0j3W5vuSFRySRIh26Yttp77YTS3UqSFCls5
RiPQ/36ESXCJwmmbVKreFYpMc56NA5bhnkv1wW3o6XYWBVWl9F5qsEJGPixnrFfp
cyxiIZmyVflL3nAECNtoTYpRlqteJ/0PQChXrM6begjrwP1B7+Y7s8+Y+DEbkCPs
FVhTZMEFZCE9nDRWYdZl7u83pdDeWIHQpssJRNCvZf9LK8/kC8wrjmQIr0RsuIl9
BcnfncyNa7fwoyzc+4Sp/D0+PW1K/wLmaTuDNgMBdun9q18HpkV2TEoXljx1YKg6
+bbVte8y2PtDetK5wQfqijm8F05jYPPFjJGIRfGrVeufsFKWgYraFFUlrtmov4BE
0rFRV4a5u+0KFiBq8j719zX/InTpMVldpRkHtK7zKQh4TUHFWn8J2TwQC+xMkMYl
G8UxaonIxrO+La88ykbX/DdD309ivSqfqE5f9BIxCrrfllbPowY0kzfUyUAiT1O1
f8+Dlutp15rcZjyygKyLnqECZrij7EkQ8lc1FwXg6xILtJbQCYdgzmkRfATTnP9S
OzjezlhvagyIzky6xnWkxGNgrV6gSjBKQvNK1BXUKlmhRhImmTCkMuJ6wxFmtpmL
h3Mbe83MVVvOliPX8dTkyPDlhHs6T0yeX6nexXC8mT4QcgU6gezv6PwLvRIh0yv4
xOY1mlh4DhJRVwYOqP9oaBW+JKlyA58pNI3/eIIU35Q2yvikctk10zH8dIMYB6qP
Mud+wAmy2rziwDCAyox8HlRsKRVV2Y7zzbVN6T4qUDXNq5AKroUhS3dJr3l8POEg
GNGxQf6S55MQQ6tXD/Zn/4g3ILoKkxtwrILa+7KH+k9AGzGa4AXe+gQBKI/iPfQ/
6a+RCtJNSjLiUIFvg7lztO3IUeAa2dh5cKBAyF6LX6Y7a3hwhQeD0Z4WyeQEte7/
Q1SGjXsFxHhP6gsVAk6VYxKtGIWfSVKQMlhF3muRxDs+gsNPyzFCrxl6cPOBh/fh
wXGj0Hy0HqcobzXu6Hofg+khqYtiCRWR1OlhIYMXJyNQ1hLoPbYk6jMQK8yZ80HM
icSm+H/NtLVGm3Zl0Kf6CROSDM+myP71VWjwTt/Z2RuwBdMqc2tsV57ovIbwPZx+
dLtmOa4NUddhDWdKjEBiPARJE69wKX2qxdS9RDRMnpFFFcQJAUNcHWY3ew0pI8rP
Ew+RtoEUDBkxOYGgzZEHeBrRGWZz9WPaklmDoYiwbaoaaPPQLutMucQ1ksT+hYFx
L2QVejLWsywl59AUkZoULV2/ZsGl3OCrias9yoFrPtv1Fd7zcblGH0G4seObud/D
Ame9v9WhGFwfjNsC2DpqelUMlAwN8idNA4/p80YX7Pv8tqjfM0W95pXv3/Pm+RBg
+jZixQXRBSW3jCG8UBCExI8num1ItBuvl5F9AIOaMnvGWXDWyp1RbtAg12bQmMKe
+hniYtj/s/4uV6HYyE0IRMd70piDV2Ihq8YPWssxFl0zBzDurz7p/Ig1Xz/27ups
UO4YPjdbh5BIsnxmZ5dDEPwuuvFo+GzwrMxFDZEjpYhG0Qweb/pH7Ceq9UJColch
fTWn86syiZCNwuzQk1XCaDm5ITDegXkMdP6H1GxBznKsw5us8qxYX3a5XeEbIAS5
kFsLZSaInpNYtq/oknUXS8Us0VOssoGoACNz5yo1YQMZKgKHPvhcevQ7682o1snp
cmlqZ+SWO2SC3Z0cZdz+sgvKjl06PWA2mL5so+LlB3YRWNmwnr5/1QANk+ddb0xF
hVSpxfIpCxL8cAfy+AnXdPL0QUwhEzh0zCEQay1u5uSj1GGKID8TOGtIPTEVkLZo
XO3zX3rDGhAqwoNqa8aVXnFf3hmvw2WP4cE8OlK+S/OELN/QNw7cMk/uORWvZNzH
eaMf1C1B7q0Xstl5IOkJPbzOXWCI6fknM3BvLvGUgRpP4JytWNfNTJ5LJ1RfGEiO
kjIEBgieQ/W54fGazdZiPHkqE9EFMLB0grp+ycCCyVmYD9onX3luAzHHSa1xjGCQ
vu4tP5apALaz0S6K05g+jE19K0mhzKFNqZ+4PoguvFlrx2EwkJm9sb0tUxsF54Px
5IpdCg/MRGDHICdfLD+tacvu/lPwER15PcOCthof89qFnS+/0VlcrxuqGHB5LwD9
GVcz8CcpGsANthcz/MGHFRRD0sIoo+BKYaB5XKqOMPxZo5EY3MoMM+w8TVcghdRJ
0tn0CbGAeEh3rIsVPYvwfA+mh6fMdaplNv5rUq10+7mB/gg0ZM3EKsMJECXn8jNc
LFrCpGQBC/BRVVDxAe7JtUZ1wAknHErVR1A0ddkl4tT+EwY+IdQ+95i2lqcvx081
MYMD8ehcei9+Ssz1jvyl5BtODg1ZJCh7aFoiA/5eg1DMSJysDHthBEhZp7i0rCrV
I2SQX3JWyYQFzakeXtTY2wQMIEMXj2qSSpzwgzFcaQLmEuzreHeHG79fC7Uc7qRs
FspZTeNO4pdowi296yFxWlhAOfuHp+SWjYb+dQmHzA4MiBVGZipcylZmTZ3nf6+L
p4v900cWqk12Q+N3Y+wiCdfteq7fcAIr/ywvTrrgiKhWXNJndVPF+3tUKSySmQzR
NzLtRgDdHPr9yBB5FyQrVZtpsp0ecNPkKStAfWJP7HyLi0PdmUuX7++aMa4QbBDg
NnMtgsh8bAJjS69hlynCBnJVfeSqNctgIb9LHO9jUjWFulDiJ6g5PyvloKW9b7i6
/D0g1aTFehgl/j0XHW2S9veoghtN6IpkiAVokr+skCjVFwWmtn/s8TEXOE0y8lDt
QC39KCtiVSONcuiVWjstDKGK/0ewLqXulsunk+isVEpR7yjYWZMtl6rZxvk3ftnZ
PmqhmFmQGHHVAfsNCBGqu7OsHz2CQKqT7ivNxM85B+kVz1gAAhM3vHis0McspkTZ
/WxseMK9s6Hj3exLI73KnSFQori8RiIBmFub1tiQPCN/EFR7Mj57QqrYPMTEXnmw
z6soSf53jkkb5fNDC9p5d1AEKxx1f03jBExGDdA2oVa9be9qzvylx7pK1BNJrcJA
x/y/RnFrZ+z8V1DZnecAAdXNbpsZ7fStWfR0Uv3Mtj+ApVAC9VWkxNOB3+aw8RNq
QD/fKdZF08yfbpIYk4KV0eahpfM2MFYT+lue9m4xjObJJ72pwdhG3+hEk9/fYDS2
hJYDOXupfCBDGt8aJ302e/IPXtimUxR3TtdiwVIup+T1TJ3tgeNtZTRN852XkAS8
AEYlUNO51WkxsT4KMn3kIs7CYqC+RGrXk/44Ll3VQm7ziv6edrpNK00OG+yHPCgv
AIT1UekNtfQpBoI/n513dsu/84+zcHP/XaaQPFInHwEJ++fjdFUGcBw14Uz2iuFj
NXwWQV7dPx4FbYpP3GSsMw2wPiP8pF8IsCcce7aVPWSK0EreYfKER3rj44/R1CJE
oN4PUnJ8gnNBYO9ZZkYasnLJ0IRriEiBfbKg2iXcWElE2sE4rC4kZu5YPkS29HQm
BKiAre05LdRwUNUl6K9KwoqB75bpGCMvmnrXU9hL+ZmQZuVrOMI1kEDCI516WNd1
zLHl7zZmdyiC32XeNHdGSVjaSuqhesd/Xyluk7HhvvyNw0ZCabrH1NavVXq+Gx0o
2QEZJ0wN4RkOKDp9cra0VTo7mRKG4fFglxuacJ4vkeXgokIBhmrPPGfB5xfaktBM
D3Xx8KDQo5Mm4ic7dsW7hKxbRdNKKFm2T5U34PmAu0VYKAQFhPqjyUyV6fzBZEUO
+hWxArRI2fJjDp5VelBXCcZ9UgIwSMu5hGqHAgzhOpqRxyP1S4oBriX+xOUmlbUw
AyolAz5PoXa4vN/WOA0fG8jrsdxoFkZc1DARwBGaZFFaC+yjpyltPtL68Z/A3gH5
P9xsY4U3FSQmU/lcXpUjjdBRWO6eoycFzRswxhxss4Rjp92YRz8OC0phwwWusdsr
XAfAh1w869pCifCcbupO9PZxOTJ3TISwTG9+SR868YWM5KgcxPSwpYsrm/QlXxWm
RfqkxnYYe4sHUWigOuWUcQguq3FcYNYQO/0xy8IRiZUr45elP/Q2PBAiJhQfzgCh
JKjERqmZD3MZx2Drryx4SVs371JUeU5FkJm87fKa6ZfvcEwU6GIePeXcgQlv1dku
JEr5rMeRPaaes7E9zyXh6W6pqmjU8Dpg68EaCEaAglAmphWv+K8kp17kqFc+pMbq
gT5Q2GJskXXOCaPSVFBSIu+O4hjoThC/o6GAFAMehYxBB7s/fks6KWDUuwJJs8mQ
Xc1zZrwz8xr0Ce+7LE4eV5GaPKx4c50YbPmIwywGRyTLYEgNUUv+CsKxOSvZC9wX
ugqKutyeYvvNa3jDNRmriYWhhObI3oXHaxwTzKNXO84INRkj2gquGDQ6ItF+FIiV
DTedJ09715vrEyeHco4DKZfdaXgJWor5FASaP0ATl2P5K7a7iLpxymq4VOZyATr1
owQc0kS0qbuCtK8a14bkRdQRcw65YfKyKKL0oIy0TlG9+Latw0JdOqe0ZC37xqPP
fsmUiWEA9xRnLi3OQNhdOefSCpMjtgNv6y4eH/HvADNr/H3Y5z+6J9iYK7w7Mb3Y
K53pHYc0dF5OwQ5mhSpq6PPI3wNkt6c3N+1HAAzEIDBR1Exxd3XTkoXnzPf8jwJi
ey8cxNSmWhKZYwzjFUZIAcdDdJVoaVM5SwmEKtX+BxWrP3nVdY/ypuYKJw29zML0
SrbfjMKCDFz7GQ9t6P/OZwmES46WYJ/Y6uTbRaY3JuGpt0MQ+/wPzkj7OBEHnucT
pMWj6/xTVtaLoduaGWoYFE08SL5s0R4++vIeq6xPF85Tdciz49r7B+DDwCufA/TI
RnyUZBcMz6Tc8PXNJB1Kl0UwAiGjvY9aZrim4mGDP1PhRTmq8CvnuEYwD5ggkwu9
VeEJu+HCBxcEd4+xRGTCz+ibEhqfU8KfVVyERBNk4/YfLA47CfWpUySANvp3Bqx4
VeZzjDhPt8UdCmuL3jq2RT5K/iIvLD5DjEilvBqK/Aii8A2aVmJKOr8ufFiCjKRS
fNh7KbSo7zop5Tb1M96w73yI/5Zve6WIilTt9wNYfSBRJil5Hdu7Oq7KP/C5sKlr
ei9lGmitLKcF79B0xJ51HNVbX3GLWpR1Jme/IPQzhz5in7/IhMFNGn0L7jhEAW2C
PXjG7lDaU+R4Cv6a+F+h+FR8IO7l+NirwpjXGp1f8DB0OKjj3uoWc2P+Z/lDpdCj
i2sMKt6rugRkPenZNJ5HAZAYC08YAblgcTVDvAjqbx3aOZRwgCWGOPbz5R0lCD2Z
y+0N181vXv1E+XfxdeYWkjH/bhYEtTxpNSwH1f/b3dynEYQSfn7FvJPLkeVWlF+0
UPBLYrDubepRLNj7F7gqp+DTt8/j3YKWUaJ1TXbNLvOSn0YCdwtfgvc0k0w/JJtE
yFNPT+5a1T3r20o38pgE3lrY01h6FP4Qxh3PbmtNIljM6CfyPCjFHAmlC5Fjgl6T
cwR4s/4vVkN4/vumD8SDmYGmp4WcS9TS82rOmgRvHZigsec+mZ7Owk9bBmwNZaME
Bc6Ra6wyKoPJGygJuWvaZss8cBFPL/vAMmhjuS83nBL/7i7Ln34vEVNoc0QPsbxF
RSrnDqhFRD2sqz0jtzur6c/oDYnsl3+XTnhL2TzNB2oyObPl1koANhkTWOTbbuxS
HNzOSx3LseS1czp2dfIhbvxYyNJEfkVztz+LcEUx/p6U2zBMaBLLz/FtBmLKMd2f
XUeEIHaMFMglvRCIQiAZIMhIDyXSB4EohvyyDIu9WUmgw6YBL3SeBp8XGJIzGV+Q
8mUvgZKEwvezTW1kzQxJgDuoGSYr/ibpjxNrcha7b3DhhyO1T0bP1kFr+5awN85M
62DbNLj4sdm2BfA5jWvDDMGv4NFMek1dNeaBPdYKZw9AmfrL56aoKH1Z/uiLGsta
JdOGIDdswYBHz1TKzqYXsOHtdOx8bh7eEt5KTNd4uSeO34YcVj6IBYEyswj1Uxhw
WTHpw4Dv1MUaHcUjrsyMwJHmOZkB6jVXDevmGKsKn+dxyEAleH5LMWL0XHBTvayx
zKW3MldUdkH3c3CrpQzkTaTadiIgqpAmaDXfm1RzK44JC9FLGWzUYlgpRxN38Qkw
kzGMfpPBRrmyC5i4lWn7Q45+Y9oic2xnZWHoNsouWNJoqo8FkJB3+hJHW8og5zNx
I2uUB+LPoMrEIGgBAKIAL2VnAoXqJOFaz2ESyWH5dLU1/Vd8+y5r2FlecNLYE6jM
oTrmDxA1RXpkXlN3j99i8SgTX9iQOZ7BYWCbUpSwMGdDlJfpfg1m/j7kwp+RiGcj
M0qN0i8ZBdB+JxNc8A8zQC8OgsqYUCLgnwUUbfpzEf3EdiY9D/TOBBcXEMpGeSxs
+UNfjErgVCRgycrMwovo2uNVHc0on81QEibWcVMgGc5vREb9d8XI+EgB0UzX+2nt
TlmGkLPAx8S1mbNAbymfXhI0y/L9d7Di2jjn3LlMWPOBzCWmubZ7+tVa6GoFQDXX
7bLYSBy8hJnxSQkvuglAj2Uf6WNfxQCb/0OfPJZOTPU7kTPHM9TNI8rXtezu0FCy
hNDCQvfB3LNJwCJ1sadU2O47glkDTytKzKb7QeZF2/AWB/fRLdf2RRb5n6NLRR4X
qvXQ42jyibr/qb+O/t9K1zA5JI0QiiLSBnF/Ch99laNoyC4gJcAxhQ86ZLVXtMYo
FLvDbOdAh0sCgICy3cLQ/vp0L4eeQBJZlBKq3fIYREd4HhaS5jehzNCGQQ7IC3wx
f5Z5jCU+9+hDsyUuDJp/vKUd5JAobxGDjL68VsT3C2ETllK4Xs3akIHw60JqMoHS
iOFy3KJoGFN+SfwrOZm5JQB88qLWplQDYxrCrdAjlbKw3kNdlFov7s4foYjHHnQJ
48NL0jS8A+pDyYG+K3jPEApj4HpO3+SrSEhzBc+E2kSmVzmBF7305QAeQdgInJeP
B3yq4wKi6J1s1IWgZ7tvwE+ZIoc4L3DH7r97w6c1KjQr9vhTpevFa802+ZuY8+ZN
KxwfrtX28Z5jTmvh5POuhG+ow9f3U4yQGlfXgspGaliWVYjxu7fxgIpO59l9lOXP
tWIemUoPwHs7ab7qEetSbgRoJvHco3BzZ7/3BaoRxLJy0ersczBJsDR6c5h2h3X7
mVJcCaajnQAmG0axSgxx7cY74mMtfRKJouL8n7wj7g1VYduqH/fFdR0EIcrObGpK
smpwZtkmTFNrowmh4gtG2IM9mVL3k3ZuBxQ1cS2zxD0QmdRsvpeblgzQ0ZyFTm51
asc06+dwtt1odlI+ixKj9p6genCb7ljfUpLw/Qlaa8Z83xrn23v2DL2SocXMxTKT
cWL4zMFoeh1Yw/XvQFPFRUPbP9Kd6/GH8mvWBBNPKQ6890DDl/fdVeim+5ktXEFg
9S0WoUaQGh+FTaV8Dmo4tTrTkvC7PSquE/ahpdXMTZkmPTq8OHGcZbkixyKIS52/
gz4L/x8xDRTmrcL5u50RJXfPjIM5Em3pAWNLkLGFtpfLcG8VqwwuxGOQHQ2VAwfG
1fSXyLZ6jMUGooeB+zxkWUZqM+ODjx7fc6ppyYChSy4b+QDQbN0MUQ9t0nZAWRhP
OtucK7mJzF+DQkFTuUH6kTcmRPz8zqad4cA3w1ylJFUHjVpGU12o3lxlZQHXrdKM
+SfDspito+p3eeYMLh9X18z8YCfrETQc7TU6u+BsFfK1kevbv/SGiOZKGoiw2qpt
KDASz521ohfcbUGmrXwN2b2d7Q1or4olLiIMMua2sv5J2fqWnzQIcEYKRtGNPcxu
keiMZACIoJyvE19IuzYPA1egHYzyTZB5VquAbnAh3vidBDy0BJsp66S6TairXMJW
aPglpoKY4HLsO4XkdTMooJ7eeODXi3Nsrnz7Fz32VS4QrQNC9es7s0TcB9SacuMa
/J5oed7EXXK6pFquc8HmoFiYXV8W3/aAIOVt9BZwmcpTbWN9/XBbvRn78P7LlQZI
c6ZVEirZBHUClWSM6C2bzCWm1IZkwE5qJVdyfALrt9RP445jO+hvUOnPIfJMxVr5
zy7ULkb4D6Fo7JRXqzsBiq9+F4UO48C6k4ofNMAaAOw6uxwIJ5ND1Jleb5JTJyZE
mVNpFDDjhw6+C6TL2THSI8U3SeezVUQgi5SPxRmPrG1ojxwnZ3VYrgjgwmncgvxT
A3gpRBIZ47rwwfQLBGrRYtoAS125jVNkD+Nvp+ufO7BmZIDyifDWYH8a82enMSS4
3DhJ8M1idU3TGo5TOHdSkfVgk/A5WOIaaEvBHwWW0Y+ajoJoPphuIQI44t/TIjfI
BxsBesrAsLH5Y55yF4ysejrSIfA7N9h+sZlfetf/84nASesnxQuaWQT5sepRz9K1
iJ0OrXFOAyd9Yq6eiSXxSkCxUurPwXVNEVrKJZR72kH1A7v5j21Hfjf2GBnRcvn9
tOfiVj8nKMTGq06XN+cKLbYWDqcjCzM0urSrv5hAi9Ss4u86q1Onbt7MwQQhRA2M
l20uP+75EK32MwER3gY4w1PS6YlNAqLpsXmYmcEtaLDkYTuJGGyRVypsuOZVkDn/
EMRW0K7q+6khXwXohTpuXlAHOKMRpHGHFRDsloEQc9k4Ionjk1c3w7Iv1FrRC2aZ
OOWuK5fYYbcwrz9m7AxeX6tDA+9FwSBvUGXaas1VlwxRqMS/emOuJtH8oDPJjNY0
oDyMYITWAuXV7GjWN0/KxQB+YQr1+pIbUbNfAeXw9W64YhprDNNtFA1bHFL+9VZp
8ZqG5szZA1V1oMy0LH88EetYLzRJLwJuSP23OsoK8clB1lOKjc1Crw8IjU0vhCP6
HJ89CBj1WeGpoUBdiDjg4UqW0fhb1Yqw8faURo0UEii+h4rbjKGbQ28c2bESfvEu
uhhY/LovpxBnf+DLhzhcKQhh+rz7lE2Xsw7u3btBk+v3m19R4ujfUAD6bFFb/4Z8
7zQgR7udZmCdpgw64BuKzcvRvBYKUH/plSFbk9tWRXmmU1q7i9Cr6vDY+p8pfIq/
WilsyMtD042+CzZsd/Bd1tKz+9E8AKHeeZ6o1UFyQe+936Gy/JCTfHjn4YoM4H7r
xypok9+gHBbmx/jOAxnP48i+qrnZAJg5xPRe53rqAg41ydQ0y+C+VWuhAWt0pBBv
uczUlMIyikXVGrXgCbHJIRq69UtUavAL/kSzTq0lfGYrRDbBk6huOEE/i+1f/yYC
AsP12Dv5SMWDw92w1n9cLGqlGhb+/gYeFikToTLYMEvpcZUOj1GDeU5Oa87nwUzi
Ng4iUt1USeue//PHSgN4LHrkt2jbowL84RTgwUG6+K2Zukj+BAxlT0Uvpyuhwxqb
hCkbDG9QzM/NBJ28L92w+ajDLsnn9Iw47DXvhDksWAWLlKI9ULQ0eGfZRQXmJ5gE
7hHfubC9q6f3DL4IiY52g26r7zze5/gEwJnWCSVrteMrrsd7FoBQMOhB95R5i4Of
qS/0wI1vOiaOX2MOvk3erWoAkGrulQLdX6me9VsVT2nQZthHE/VjjFtrEAhtDzDq
lDU21J8rPaPAYT36qiQfhXvHMzE1kSB7QtBktbPsbgN7RyqdCv9vhSnqU4zi23Js
008YWAv7Fgfg9WlW3lRSlqnm/ZUDAStQo2wZTZjxOhKU2VLFyCSLCDR170tgkiVA
/cSTBlxWmqeh8TduT9v2s/+Y+iByZM4WViyuXAI2/eT8hvXM6wLvyGVreaTMYVpY
jmWO6nlGPfn/KJwvUlB9kjJOXHUPXu2UlXnFoBfPPtrecpvZXE81PBqg5Sn/tZ9z
eu53h6GUVnXnr3ARWNTNlDY9GXZNSbvR3/AU7FcZFmuuMrDPDvfxUVfkTr1+y58U
CU2Il9yHhdaW9xeDeNyzMAnAhhObDOFH95Q5vfmPyvSOKbnPHgeejhgMvba9DJVb
88U68q1PB0a2aLvVjYoS8jihVThq1xZUNgSsAq2DmIZy2lB3HSK6MH0f9XUWco1X
8Y6AAkc6UCVWN+t3almEi5Jer3Kj/JAW//bOOUitTCvPkrEK4+NzZsK+QZ7IqQmA
JYGUe3RFINn9bVMJhr4uWeofTR4oK+yf1EeVjS2BTy85EoH0hPzKuAcqMeWp88Ho
3NG3F1rnhctEJB3N0WUexO3+Xa4uohno3xjkI8jbTlm4+XxgWAAE6t52ePr9n0FI
hrlOPaW8ZcyeeiEaL2fh0b85BdVPgV0RhsIVkKm6NqE3+h0QntCoBmXsm3FxSLp/
8AQs0c6Ej3fnKa2hAEvICQC8SCzEt/sET1KHDeZjwmUChptIenr4v0mB/nOEsy+D
zj2vAwH0pPskHZ3FR/WpCzKPAvtFXTMA9PzK5B/eLBSwozrxB4SN661HtmpueMtj
co4KCDcUd0vlMPebN+OpmPWmR7putFzXhCgEAzJs+ml4toUiipW/TXCcAHfY3cIC
DceG2tqlClLFimSW5wmy7TSlbqefxCMvD/01XYmTfomFvt6pX/pQgjKU20yrjpzl
dFcwEYV1qMgVg/BnrSHCtIT0uVwTcNRjKlX2SqjvzR7BBG6qysq95FlGHJ9W5ex1
BzZnBXrMvv8lDygaLiMfKrnhQyvLLoYxPerib0M8jNmFFA48PLNAd8xSLTlWrOeT
yhht3LoZcNBO1M7VSBWfMUIWU+HNV4pxHySPYhkh40tn1WsQLGZgzIxRH4J1D6v7
ANukVBzgV9JQRokmImGqytepb4lvAP7wlxY/QqvPH+hN42SNFT43w9BT8zIE7Go7
aHqaRfENfSHvVx2f4Sgp17uF9KMB+AWINzZOm9cE0JlVp6IDJqs/Il4xIZdYPwi0
N0zJYufkj2jJ/GnFSw/TLwDaQMgauGgnqwdmOo/ti1AzpXWmT5Vt4+Yi1MZyfBF/
Zsw7+LUMtCQ3Xru3TgORdzq8XEkrpkoONRulAT6kcqQCkXjB6/qVGxivQI6Z4LUO
635OhkJyLNoGAUEmo1lSa2uxCHbPN54zXorQSEfdjt3NsFSlGBTYyr/mmFsXK175
J5K8wjn0bxbp3kLBTSLZdvSRup/IsJzDbh5O8+y+JWQl3kn7w3a6qwQYrJe5q0EA
2vyhGz1NuXtirsA18Cw3hcTf0tho3RUrvXpClLjaURAMyZUKuH2XyNHiHyqdfp90
X2Y9FxK1AuUXLjLM3MdSujZLfzFpIkAyVLWyMDYWvqkreV4tHnMmxDm/7/YU0G+j
Q2pk236Gmh8fapu7BFQmJrZdHeaz1IA537NGAbaOC+JEZk4BQxA3MeNJ3MqQ/jrE
0hPAGgdzjxT4MzEAGjnM2ID/8w6snm7oHwQJUvZQ+8cwJBp5lW8/1iYjS5a4T/e4
SZHlFwtQGg+Qa7TqvunyUsAZdEuLFj24OAIU1zcLh4wrdbQr+kbLT2wn6kbny4mP
6bRTToy05EVymMbE/lqqZtW+aUdlCEgQcrni531VFgickGyDRm2M8iP2MVCBi4LU
QhO+K3E/tB5wRifrF09XeOgNasXSbXQSmfHACjWatWhO4ABfrJZVlGMyg5VKYCzz
G60ZKAH3a/S28bIUOvrC4F+H9kvbxzSTUcgroNTUFdwkxym17WBLdb3FZ/1oadCc
YbYSJAiZU0ieXjKHPg4QYgolYnD/jLaGuMcpuv8f5Moiyu2H+nw+WHSwig8nyqvV
uv07tQk5gxyEiC7QlKMT4v8Z2m+DBYu7lV0hV8yHTQ2pvQ6SdTTg3KkhUn4ZJKN/
5bFH4Zw3Vx9RRWyHvIVz0EnXT9VROkK+juR6TaPbRbp+oynCHI/F76FRIvcBGyxH
DblfHPrgLIS7WR8L3/tdOpkEBI9XlblY+3CLOY+YQR1pKyKDdgQhC1sC1ShEMErV
OSZFyDLeowdyCaHTjJgje5PdVtIt1rR4ejsJN/2KH/mzlaSUssAtsEjZpUpHEXXc
efn8Un9TPf2t9Agvl1oZ5D40eaTo2s1NhfrFFezsFaZmSzLN658OIu5QsDmwxH72
x9n8VCT+yLqCI59fbbAVoerJdsqk3WqkbHLxy5dN7SciAb7gV2U/xXc16Fu7zhQ/
F/YUX88K3fxHSdAJ3r7QJ60BqM6EQp2wgEJ+dyzFIgdEUbn7nAaRUhKF8EQ179QR
/1N2Y3QJwdw7IZMrNwO3Oq4/KhJCqJsKpTPrIWRRcoSL2/QPvULT5XzLgQ8VEyZF
nWHYdspF3wAqS7bogWpOI26vibBcdrYWLZcya66g7eug1BwPhh14uRhWbzxq/SgO
Fd6VsrROYivhsMW7IihsPzHznuKWE2Lq9kU02fEo0RszwgDKK4x5hZAOSRgEyTFp
vqWd7ZM+7O08uSryJdpd8YEP+/AvNOgqQ6c2TAaZOKY7SdOlfaB+XsT19ufRqaYy
qVqHf661vVXjkVB2vsWg417+q0jUnSvxUHLxF6RQtprDIXKHqqMT7wQn9aIH7N7y
E9eMgWWI6BloQUEzkHro9fl6U+L2j5dCJMMoY+y72u6lH4mQxid9++txpNw8hW1T
X2EhnimFQLAcQNiBetjNIA4xRxdS0xAdsw3cpI3OSqWR7Ir8v+0HsnFMvnDyiDXD
ycws5kiFrsZuS63+DB94iWGrWQUaFFpUM4984A1hBw9xnZDx6QumflpUDP8k8kdM
e9Yj9erZNod4aIF8vO+mz6EqT1/Suv02I9OswvkycENKPHcv6wYxPcYHn6lI0lD/
vPWX5++mRsUQxN8o4vVS0R7KsFLNWiqM3i9QyrTsX7NdRmCMM2JjMxOHNlYSmcMO
OyIG+BMU2RjV3uHtcva3UXEik0bjoLoNE8GP83EOvzIHPI7lAuufOP/AAe2B9Ld8
88R7q8mKqD9YSkuvAgNIrd7fF8jfkTKtnFmyx/GIV7VrK0OfT02KYOl/C0LfKclf
nZTvRdHA3EzYvVzB+gJthoGdcFXPMdsKXBGZmEpeEmqJcE616SGH0JFuzIbocjj5
tNu0LSUwtyi7bbezouUW7qAYy8qLDlR7eOkuHr3jcylTwGqMCxiNh9Qny3hdt7SG
ElW9Pt3SrBLA71byT5WGmd+BUfA8KBBRMTVoxAKTA3BaWXj6Cqz9fVF9s7tsI8lD
Bnw3PVnVQwmb1eF3EM0s/8Pw0VoCtP2+kZoVD3kvijbkhySgJu0PaBWLsic4NbjZ
3cIsiGV1WDazBCQXSsCCRabvjLJJHjs66/lR0s3bfLl7DMSy8+PMcxNZIGjmyjDo
NauUMTlhXon8wDM9SV/BIf4V4tGkVEVWGIjScIaT4qBdqZ7Or2YYJKRHZFuBlnDl
5jsGwUH0XcEBbGp9vgPRm5VwjRb/fYA1Sjx7agJWxa44VEuQ6Yj0+kH2CTP3G+GE
vteKkjT7WCZv9VFL/+J0kSMknULPHNz2ffhE/pufBLZ5AqnWM5HyehBdfaHazDM9
zX0j+fEcaXgLaQD6HfJ2cSm2q6TAB5Yrqwwv9dQx8VHcrCEH8Fqdpso0zzV3eBrx
uaafBeQw+xvYocUNcsts2GuBDEKngLJtrKBTJmklWhPZ+zFz0Pt6cviyMRpRL/1Y
a12Bv95qCr5tYxJXxovhMwi7lDZh/RXljZ2TJSAhTzz4O1u5cv7gluEVCSGqEVSD
TtHXzsarsgulNq4Li9PXd9j/FIdALEEJa5ctNmTOuRjqCmDou+VoQvyQZdS9P2Ih
eJw7etsadL3VfJIBvLKvo9KQCKFpmL/iZghznzzN9y2ch6/TCqi6VSFe9IRqcveb
xO/1XZKk1cpQYia8KJmBVDHIbdDnss+LGun99TyHpr39ZMdTxASgjwef6V3PPpm7
CNjslw7dSMRsDKXEEErlcVIfv3l5EbevRe3cKScYwwHZCrOXQO+kpI9OZoL3w4eD
mmyKsePja/mOzpoB8id39mZyJQgBLhJbbpllEJ4HOJWbQHs5N60I2HnN1nGE3ujE
JlX8fQH5s37pLTTWm6E1G1g9INM9mi6HW8R6VDrqzir3INFEs2Cn2HAVu6n4whFL
HQ4XVlgqKjadXLn9sNUyMm5RWf32QKEtNms6JI7Bv5U/Wq1NNqAG51HZqvwwUZHa
TW3uRdSfvooOAHHWLC66eNxJV+oizzqANbskcylXo4f422kOTWmqwQBN8oi+P9oG
JZA85klK0MIfXN62Ubcn6Pp4ir46n7hg37v40OMgvWuF17/hS6GwoLNoOnLsyyRg
UcVnwbjZEPYMfc0CWjSYZpW24YVXL8LxAq4q1ZrL6fR2JnIK3I0dBWkWNGj5Zkhp
p6sHpvKEhYUKUTA+Mk1+AV7FBPM3Nb7/VbsECSdZsIW0L4ZVI8W9pOteC4ktbCZc
BzZohel9F17MdSjgawXqdd9F1CPpSXNTBHp199wjbLVaTUk3iIrmVkhnpZdrFhoB
ZuKkIZEsjaKffGV4f68+H8hr4a8mZ7TC2oHuWXaCV81qlTkT/kcdg/tCxmTFGD42
v/Bj6HG+NZROhAP7zCE8wK6GmEaQnzVCJYt0P0V4iK92pPDoCaH5o+mFdz3OdTgu
iCnx1H082mb3ubo6cTvGwea4FsfrScWWBVFUjfeJkrRC+lJ4AqtW8k3LZOR7d064
2s1JGZ4bAJ27DhpWqAFhvCQJ7d/i7S/rKWW2eW5pnZIcS+CTGkYmsJrWF96JqLBU
OryH8MnZ8zBzLn2j1cjjMMrbZFnKX+Hxke+NVVRyAKwUcyF2qLqCbKNFA1pHaCBX
TguBUnOgobFSwbdJxKD8HX+I/JQetiPybVbS5NuwMW+zWu6rjITypSTY/UEQL7NQ
PjjFkMGSBmWjm+oXC6TQ7iKQJ8HSaiN+BhrjsaKcyboVLqixZAaymcvFHmpwpV63
kuWdENxkZ7cpOqjhko4LI42pH6giDux/+pxAnrSBKjhyq12PQ5p4k5W7WBls4n+T
rgK5rfjwJ7vj4TQW/0rpwicPqYp8JWl9dih6ScjNBKfOVGI1SSsyPU1clOGQ5hGE
ws+U5pPIGfDBAeDHHfxpNq3aeN7V37ZLYWXqCV4VUHOoiPjzXRN8fWqAMuDsElUg
7azRrJuthbwf6tKJHn4IPWp3EJpfiUQbcFHFsWpXZXtDvgrzmiEnji+0sZ/NBajV
jcI1V3gEwnH/80iYysSgkJ6N/kOOJUvdL9Z1EoqmekEOVGMdCtnoYzYFVNfY98mf
LNDCPRl7uCv7l4YrAbmDGkdBAAlguPJBi9p+KcLlExTXifdaw+7nsuJb5OsKdII+
w3B4o5VB5gB0Xv6Wc68ZiWJoWQ3JgTRjg5+7nJEGJ8ceBX43g7DGdxS5peL0Y08N
GZZYTYjwVUD8B6LApAz7SUML0/ZnzG6wCVfWPGOwrGqqPiPRnPgE+B62l5Z0K9Vo
JYw+qMojr3Ak+K4m1ZOYP5Yc0qdXfST8+I5zmqiddnqMsO+H6/vc1tkbG+Bjluz1
cFhlsnLzkjPPhgHQC2tG0CaKbLhCXvTsSrG/3xGXVoibTLStTrrJzL3K/Q1EtfPu
wqqQzJWq301NNPSFwquundqBmM7Zsk9BTDN32EEdNpKOSyzmDtCDxKF1FiIC31aI
cL2jt7ZYqaSjCm/KLRNIO5BiXEieZf+856GPEcxtPcWUwiKFRyicCaRmKVQ65R52
aKnnxPnEOa+9NafxnRDEiDWUKOryM40BGw2LWO78GhMKGFroogDqrfCSTSrIumfK
esrR7c8OKIriUhC4ey1PaTAefTZm8ZQ+w3SrWqtVtBGxUrBjxlUGTmx05P+fgrnO
63MSExSyUQGIGzdywyD9HvMsK9jFmvxmV8fVMKpaTMglJpsaswoo5YwUSPyZO0sn
A0uY/8iiwhdyNcgqmYw82kHV6UsDrYlipiXm9EQttnXC9MV3tfLCTQxEJstgQz5x
sVyx3f+SBkRTO3wlRzhNIsEJeCAAK81nR0mNQkV7a3v7zO7+7aT4zX7ijIqY4N2X
JitMTqqE7urfd9SQmG3zpjlO6I1COeKJagS1CgCqwAg5fy7BS8styWA5UlsUSqz0
ZKYbu6Y1Bov+UfYLEQGrZgJIJV39OibcX1SSkpPRCINh/VvIc5X8oYs9PS0Zw7fY
QEjvhBr0Fgw62XLXIlHyzAYoH8obKj/asEGqRcYBHm3AObac3Cvh6POA8r1R3NDo
STqoIC3B0hLjdG5MW5A+fRFWXDyWzSUZFkDjxk5wv73HUGX51KQgPneJGVXLGUqE
uOqYKOGlxZ89UtrRBp65NMajUCTOjlbMhMjvNO0RmO2FycSin6UDTixXBPZi+QQx
jUPjkhJjS1ATY3QPxOni7lyqTdDCppZ6VVxE1UgvwlWXFXCVYK9W9WR+hhUCVUli
3nJJq6IfeLJmiOsDBkEjNYKIiLkZEwiegYEfMk11eEHXvyjFTM+d2CeWagsBDhGo
cdfCxhRm5886Xtfh3nhYcdNO82b6aYv56c2/a/210QorwJSA40KCiAvx99g/Pa8e
7nDCSFoF028ctrcXG/kcNR67JADyoL8HKEiwgxrjzNoBBEvxjw5Vferk7AD7RCaY
vpdF5F+Imd3pUF3EPCbonM4IF55bVIMsX3fn/9i/JxoketQWpp41+1R5JrfCmQc9
bNku0qdyrfvZTuUAbGvXU0h6Cwb4y0qaY06jEDibyMGjHfYDSpzlV4MSnOAmAzhi
LZJOaC2fKoI9mBy6RLrzdRghQwkPLLJXeiqZHDUecFHferv+qzwjjHc2opE3LvX1
klYAQqXQylS06+dVjWe6NgK9I0O63XlNeWg7Cpdav56jUxJUjidYWvZIfvzDmXYo
m1akGA31abKwi6tcOnLtHyFWSbUcNSeDiSwDhwD/ALVAxHyKIitd9GEdVt79QQuv
9NnvZtH1B0FnggnY4X149XOCEJvNnA1MLJHet/bc3DcycYHV8dgE8VeijNbwKBGV
AZUUHOOOxcH9tJTV3wKN1hzoIIlavJQtAkBMUWcQmszNHY0cupHlTgCFxBkYFlim
3P+f2pHWU4ajr6Ogci33ZmL2MwVBW9gSVrQ2JKnByk6TdscqPxOQzaCViixcLAZu
G0KbIE9CfvKGqe0RaMSTZZcT/5J3oPICsGUNAZud5J7/35/iN7w+lW4Ygfwi5zLa
EpobFkM4ZvH2rDSQJwf23yxjLjjddM2L0NCd1oR6Eq8JJHLnOHnqQDD/Ks2qFeBq
zAOvDyvWAC25xlSs32m0Ob7ZESWFHHYMllwKsp0Sweiakj0cyb23MgwaOPru3swU
nYQ1aRba+fRp0dCaDEqzq5FJU4k9XWLjacYz1szjg/LeG14LWPHBsKGfLs+clwT5
VV9OmG5qEDT+nEFbBlnlu4v2a903qBPUcKSUfMoM2T92hexsJW02rb0aL56nO1+t
lMuGK2eLZO2IGpNjbng3Xz4fMny+Zz+xttjA4ZZUVP7mQRnnaBbMm58WL9Nd3YgP
tUI0Js0Lgnw+RvKtEud5H16QZb0IIP076EROmOH2aE2AREqxQeO0fleWPG9aYOEz
R44pzHBHx7uWDyUQ/IcILJGqhyntFpdu4xFOpeeknh4440W4gM9CkF3dEvlT396v
P4i2dqezZp+0ge5quztSC1JExzaiZ8nM7CHdSdwYdQnFneVhet3CEGAdGBmGednu
o0+lt6Lhx1h4dnWFxyLZvWWwIjhn1IGgs/073Mu4BRHcZvopQoO7EUMHZrV5wFHV
0s5KuOBGzQ6b9Nxp2MGN7rbxrJCM1SR/Wym1H7+5e5RifNxo0/onR4hkB9J3T3yg
qfvETL5DQsYPiiuctpmnrujMb4jXBcMqQu1XXKeRPivEk7Ax8j37bwRXrbkNGsh8
w35zN+bAm6yoUOXIChKhQPOiD6vBjcV1NfVR2ZckolveMb2Fvh4R0Dy39uDXqKiY
LZgXKDMN2M7oyb0U6xD3FPqznmwU5lDqjM39vlYpISaZZokLPsGPwsPoGbyrFrMF
YkbGNcnt/HL0brVmR18T+VFM6E5fiJQY0n426tvUlGrmuZkygf4C8BLaI9rrUi5d
Y/6G0+fOniNGCmmNNXXHrWOR6a9wElDKh/DeV8mUVFdoVE8ltWLMksg6MhOFzeb3
zJ8jcYSiHJb9hjamyPDJpmpjaXEGF2Es9FfCk4pCoMpk+o78XfRayGiyxttmd9D0
TDBHwQrxd7U1ZQFO+2Xl8b9C7ke771gKJlS/csqqfI0ZQDzUCnt9qyKXoMp2NfV/
4RfcW8psU/ZhkjBB6Xca5AyLYVP1tz00aUUerV7VH0v4NINTVoeVIXjSSU/uW6RL
b+P4/P3A9IFcocK17vZpfVYIns5E421Z6d8VFDnycJK5UeRknUdN7zOJXVNdeEH1
kgGzzdnocZjC708j1ceBfVS88JP79knvsnh6fa3yG+BXn5zSwNbrBnjWb9XinPQz
iNpyLZJvLGKPkFHmOeaIYXZshDZwUNZNvmrKdQlIrG7xOD2VhHBmXGQHPoWLi5BE
R6O9tDHusZF5Oh45LxdOsYnSbTnJqa5YG62RvPXrGlAWs292dIbPtHFEGElAt95Y
62Bfgk5hPCfh54FL0E9Q0sVsyo3saO4EQQ0ud5Zi7oN+R/sdeXymu4eEeb2uwQlv
yt/8qOhiWUuZjdLur5yFy01gDFYkkV/vp0ZoVIK8HdnuSrazERbbZqQ1wgrqYyMY
nRxeyUHRSlhIfLFOxvFKhZwboxMpGZnjC8kJI9IkAKrBkMo8V7uc27T9gDzwzbbO
1Y/NTA5g62I6cRxpyw7wU0GOaCvGahwlIZdUj8Ng4SZQmlf2N6Hk3Hawbj9/nyku
PwqXFSeA5r6t3EnPCDbBqMsqavCO8rMQN789wsZmbjwP6dhGQ+KildGbeHCsQV6j
LP+NjO9fizIpIRmsiLc5knJQXUylwUIiFaP0r8gOAqKjhJca25u9WCwSU3qKzDf/
J2m56EU9fQZpeDY4twnHvomI5GOVlc5WFIfIywx/CL9sfmSga8/GEmmDHb0JJhcv
1/gura1lpNqQDPHQWl+RQLLYSPK01zjdeGP2dCJxzGHqZ+xsoWPdEyXdwy/d4crR
VqivfP4LnI086Y+YlaW0kWIBVHf7pyfN6Vk5RUCPDF7Gm50zvGXbaqrvi0d67M8C
TEt11MszkBq7dHnrVm5IjiQvnti+0JJ2SQKqFveBSQvb/fuunHJy0eAeiQ2569/8
kSxaKX5u+T0+YCwgZnMPmjoM21JxXONUGQxcVUS/Cqyz38ixj9OXfKrLzawbWaAZ
Gd5zJQOCIu3OMj5s0ovZfCIMYWD9k5i/NuuMMhsQHQ9NUoxoU2kSGYh40nJWZSkN
dhVUZQZFmk4yHBCFMlxaQSHieaMSbt8ffWutG/zjkp8eErCZWXloZwl4wQjUPlZx
PHXVwo9A28dSyyWS290/lQTpMaj3n5NWRRot4u3qdv5aiIYIiBYiJMfdnAqtBweZ
myVfXgU6ZnoiVNvoNDvRcG1K3JPupszypHBSxz6kwozy7DC9xUnf4tnvt6H+uY7m
HuZdnboNP3u3KZHYYU+K/1dC2dstyf7c6MNr5D/ldVTAxwo17ltn3jFii60lTcj0
z9c6qCMk/+cycN5sfunKfoMg4+Hq49fJNaeP7YtoL4KD4Fj+4KvXmOa41FZmcxv7
EQ4b+ZrBfTDZkxKgaaYEcnEGICrqLYi23QCEmP2bYvh+U1XwI+dhQC2z2JY1L5mF
SaR1mW+HxypD3KkpA0uCQuh92hq74Z95zL1f4iXsr8wsKz66rC6JRgAZYDhMB3wa
mS5KtEsqiaauy1oQbuvtv/jYYTrziORPqs1MXBvnSq1LNF79pD7yvnBH2uxAauFd
uUI6sMaHTVVOdzMpHzRisW4GPh7K3DQt4RzsIH98mmzrwQmZ8G5V+AQIzgdVeVfM
7d5G6aAXsA0ne+vzJaG83fYQkkEon3brTDVUBBQBlrt463AmiFwkgIrLEVP72TGl
eIYWasp5nY51cnjKto763tIyKpGAa7iKffwLw5XmQ7/Up2TtaNJf6yseRv6Ls4Mh
EjUDRrZKx3TCGNUBqe5VK7fMSpgnrGvQf6w1M0DOI6tGMjPE4vcADVnovNhKA8VZ
9JVihLjWdq64h+gdGHua8zT/r0RFTA524FrHhItCVlkFW8l2EaKzMMmhGVbOIoV8
f03CyYwPSVUaa6Pkoh3GRdTiqNx+zzkZ2X/HbcXlUTZGbLnksxifr0xw9nrUxkA6
RTkuOGlr3HyXhAFf4kUCykOgfY3YISCXy0v5IFhypf0/g3FNXG5jYjOFhDKxw15H
85Tkzg4llVdmPEV3sW2LBg3B6VE+QENFaVhvN9/MzReX7l9VAtvlHYayM0Cz4Yuh
44otgvNbFJri/SgDltBPVhZUXiWa1dLOH6RZUdnMgYDQB9ZtEgK6pN2wcN3ihKGO
/p3Dt6tptRIKOIxIs93xUT6OaCn7rjiG7aipY9NcqEcjEwcC/t4eVACljHq2A7ss
YbA7MCpFRTKLVXiqlM3WNCf8ExNXuhKUKGlBs8+FK0nJKK8pktaIFJNe/LtWc5fF
foB3Coxq1KuT1wvupSGCvmGE/95Fw2xoskVfH+OarzRfEjdSbTFyUwtcxg31rNTh
wl6kxALy997dAKcgmejVkIrIET09E1nUrYZA4mWz3M2fJcJYgcZXGEIxfURFOz4E
BU0U8BzgrMEKf36jrKQlHAyfNRGCP7MbsDwRfHDSS2F9jeH+ZRaoYQfHhurqZlul
YcjjfaaGqxr6KyL0L9Et/JW6wrMEFl7/hioYsFroo7XjgAyi5eQg0m/1cOmDWWW0
6mhVdeh7V/r9T/yzak8PHXWJx1g4Btqs+TpUFeBqe4PwKgqEWrV9uSOeFaVGwqpJ
XumrufPpUxDPUmav7f3Pbn60LzngEmDrr1YyQRM2935sbtMrLZ+fDQO5/hKhnsPP
CP3qi+dXj+hUmc4sxQKN4W8W9cAwwC17zUIPYICiIrAH2VJRFLrzCyG5HgOCsrof
Q4pVySi7Lwrttf+CklF334WyO1tCVvdZKcjw26CWxUUjSJgoAoYnKU0G21NgSCd9
NciE/2/xVQqMg45AjbglcO2EPMXGXeTg2jLck1NHKnA7HNNkU8nrWo3VIpt4FzZY
p8jVna63LfARFxGGyu9cqMCpqU8CAUNk6ClPJzV7qEwSvIcyfyKVTGE5W9vO8wgP
WdNcCf0L5lwkLEBMwOoIgmov+IBVwbs7cgwmqSmr29YGdX5akXSHpwgxw4fTANPV
KLFTQYYcig7dCyOURaf7nushd4G4XOQqebx/Y1bwzNe1PUOGUuAKNw+fZhq1sHKi
59ywB0QsFnxvzpArGT6tF4l54h9isbGLHtUiSo4NdR0pTm63Fgxp0A8IGH4cAs5J
7WNDxyzsiW41V/j3Y4gNOQbpSqx2aCloqhSpzjsRyqAhD1NjeasIiBlxt7LlD8mv
4iX1NUyO13am3sc6NLLfEHsoflX39FDV8Xmt3kadIJp5ff+x800AdgyXHgAvT8Pv
2fVWBIOgVC2faGs5z59Jyj2O9KWerufjXeKgRs6TDf92OcKNLXAiezucmpaZrypB
s6rSrgM5BE9ihYzSBxRrFng+KFg+3z8n+PN2tautBiY7J2y+sUSkKTd5ccU62Vp/
9CGduzlQycDd0sbRFdJQzPoCH2Al0nr5212nOKuyjTxN6OwikXCZrJZdTURjxwJP
WuTRmrkHbOTNXjeG6BC0s2HA9NPcK0MpJUqcL7diiAimvkiWzcMk8YZat3gydZTa
WiwfOhGKZoFpfw7VzrJRfEangFWgNMVXuaET1BFyLpsF1zpJEPcJfUvjA2+MSzJy
mRJaKMLTREFcTXfViradOrCHwgX+W05xfSF8R0rTK2xaLfOZMY+42FSRTsMGEOAr
z9G736c5JtQLJvHoMSY/OrUvWwdQKAylsVgXGwbqYHZvV+ac6hNqQSToe+Lihtyi
Ok4Kjto7BHLUpf2FZmK2YIFURG2TpnkF/Wzgxg0fQaV6al53RQppcaZdXHyjiR46
Vir1l29HWoaYGOgAGqpO3lo0gHKCerZUOt8P2VW4Sb2QzA3lM85xanD6N8eYo8LQ
0pB3iovR+s8pf0NJtlNdLgSG4QhNGgZdqEId3rr4cf2HQH1lKpwVEMHJri9IQ51w
t6xsUN9jEuq2RCIX6yZWnc+TW3Zx8SLFw2pgYY0ckRbd4HZ/VVXi8TiN6hJ4kgZe
g1ULE1a9GuS9PpDR15xcrM/mbZ0M16lKk5emqq1zPwoJGP+z7EgnjSNsGV7nD4SO
o4InYYv4oIewwaQqhdp+zDYW0LG3TtY4Es/ABDe57Y/4bSNlt+6yQm9+Cwed4AnP
/b6yuc0+EDGwl1hAUlTJWT4+3L8Q9qqcBa99ILPa6pvU7JnYw8FPPcr5z+417blQ
3G7yMlRDzw5MBmuKlw2EsE/8xIcOaesCkgAjTNCT2Tq0zImg2kMspbZX26c8Nv0V
BijankN/1LmbffSsDNrgc5dtkeHkJoCr54WasYApDGrxfi/MHLOmLoAEoAknzRdN
dYgvOGHnOmzdmXK0wa0hGGJOcyuqgPLQwmzdW7uvJWPt9JkzDw0g0k17Zhqk5uj5
ca2CGFH3jcXNdYE6JjY1p+Xb7XAAAjfOveHVGKk6TtxEzUlGA7HWvTJbzHQPmn0Q
dwLObFxfTEadfZMqO7Mn0+uo+vKmEfv2SmO0EfayUTw6/zxGhRYY9uzWyI/DTyak
WiHaNdF68LJwLJHAkOAA/wwdvdNyTjCrgSxska1EelLPF5fBMiRC0rirXIcW4wNd
YY+wlje/wZ71r2SS1vnmWBvQPtylxkjo7wBsUKKEFlIBKoKE0n6V4AqAYzIGKW13
FneavYUB3S71KFsljZEV0TOUFVoL1PrLxsqakEvgUq7wnQYoVG26jPmhdAaBtWRx
2ZvUTbzRhp0qbHxd+LUZu2vYQL8evuOWrzgriCe10+DEpa3igaCT/TmKkdh9aEm2
pO5ZMnTcV0NeKnaoQTR06gborZ0F9rE/TeN1Sdncsg35UH+Gt3KYAo2YLbRlSCgR
iKAzi5pIz/ny0D5JTeYAW2lgw4dxZp8j8fuzDYjgu+AvFWCglzhukQV/Ks/cjSBF
BWFhI1rcse9LcVfTqUzVOwHD9/m7q+lLIsjSbqj9ZurANpcyqsJEanItDejskW1W
w05gT7qrfAZTRBAgh7HZhWq+m9qbdjCkJh1rMVC7HcA6en9lKoXCcSfYvyse9irM
ZFmohZ7QK791XKOV9FxiWz1MkESq7hpAbOgRRAfjtCsr/dtd5Firb9VVMBDXKKwg
Cp5Nl4D/OpnmwPJM0VLfqlT++RHlkoFVTiJmKPkPGmy5cL3vM6Wax5/W6q+wKZpc
m6HpfVqqRioHEFItFZrJBZHeIPZRxPFyUwRU36Xx+wgZ5NXm2vEtFnPz381Tb8wc
zxNFRAvLLJy5IT8iVHDKyHZf/3hRhtc5vniI6AktlgAuo7SrgDgiT0yz4nlRfmOt
Cq2k4CGiFNHg1uDm5Dwpr97K0+jrl4aVnL2OALdQVm8xpK3ZEMmIquqQnmy23XiT
qr83//VU9/eMLS3Pjc+Ul6ClTAswJC0P2+cgcGobFHHJu38Rwmn1XzXeyuasmYzh
+QpVPBYyejekjDUKHRElKRVx6A/kZWD9KwR3F+iZUiXfnKfJ6HeFE8Pq1BiKiTr9
FFqa8GBbQjk6DyAXSSULnN7Qidcq38ZgOf/r2oDBqT/nTjgdsEArAZ8e3BB65Qjf
iAKZZ1YUTefMveXn3CczH3ty00gYhFgpiIY+86/6WCJLQ/fnq3A+ueEAc6VyTYsb
nT/LXAVHzgRWgHgCLYevm2goH0eDGa64bZncs9MBAOEhn3xvyDFtTsY0q2z7rEuN
EYBe4sQcEHGJ7ktd37WkOM8QgTVQ+C/ImKXOxc3MW0Lqc9CKueh9MhbahOeRJ8DL
wHzHUVhyuVV/2LrA/Vu10HSukLKaGQ40ukaObWCxmu+UejkrWLEtrGeas/97ZJda
PlqOVMPHS+nH2bus3M3hpflXCytCzIMcOA45ZV1M5juBvhRXWbN+5XenfbHAa7/5
Aa43OVO4OMB0mQdgTNIO7uTIuYXZTTr3fSGaMCcC/NNaq8HjBH/J5NpR2YSqZuFd
Fu61x39hNuZHTbPgmlYs6dOfHMQTz2Fw6VgECAUcuMNtvLipwtEoUdiP+cflModF
dg8QlwXwsEyFuevArWdxnHQvqawk5jrmmkLYHZHLH8OFcftw7gAlBpxVxg1gyNp+
wxGKC/Z8ihpsrljgZ+hKOMXcfRm1KeC+jWW5CSaeCCYLaIZw94J97idLhg3WNAd+
OfG9UuT4m0VwcdJzo0wXTo6xnfCsUsLkVq0LeE+ZEXwiFFDrd+0d6DOF5K4bhhNB
dRRLMXa7Xe1emNzJu6vu34bO0DRAbMKjPnR9yUF4c8OuoN4XLfZ8bnI6u1WJjQ6w
I1EawUqJ9cHRRmaWF6JVP7jP4nBIrw+k8YGTy6COszSUGh9nOiJ79m2yS42WKN2J
PVlzgorHu91z745Bakc6x4AJYl/kymP9sieb0PKRRhkBGpjrV6XpLbIq0Ve0bC6z
Mo4LN9m/IV4d3azRiPS5OvIIbLeN7DQcb4dH0/B9iCCWy65ebcljS1uy2QW68eks
hS5yRJZxVQ/o4aBnlsDCCKkTnFYIwjot+/9lvyNZb6ey74m3sgLEGDcBkW1qz7kI
uIoXB/Gc5vLaCDhTaMYw0Y2HhoJzERRZ+MkJwD1PSRRRcBFoXWLh5tfOb/Z4zdkP
uF7mkIi+SDQne7Lbuo/i9BVbvYz9281cecYdjDdw7DH204IWIqP3j2EhNE3dUUrB
e1GpYENyuA5OKelLVKh0ZCA5lphrZ/2BB+0aj/VPx3na57WSd+SZe1N3pN6Uvn2D
83dLZW3FB928tIgF/x0VoZYraDsvlCArmcXXLpawk+lfOEbEQHOnu8shxlXXN8fu
8oLH8gAjdYTrpSyqCzUURWAkeOxs/Qypr1c2kz0KvBD3eHTkAnyldAf+EkI5YyMl
58rktnSKUvP5SFQ6PFz/LXGSqlX0r5XBwuVpe4jw7fe0rkSMri8cp4kPyC6O2pFP
Vb96LTv2Dy93ewVgtx2/CILv+Ir11DuI/fh5fcQfh+JfwdBTJ1N9RmJvKZZfRSCN
sMHmbx8ET4cz2kmJkunD5dhtEd36+7NuzWKkLRFF2sTuCAKPjMxie/pPSKXgoysx
jwN+Sc8ML6/QTEkgUBxx8Ie3YvEL1R7R8DW4mErq+8gbY0SiUCF7oG42KNB112rg
ut8lyCDvqw3R729ydo8tIuYcoXPmvRn1AbuFZNfcEIwKTzozNOrsP1NcvjzVaJEf
jfgbbYBNQngViZzx2keihuG4Y6ewDNADEHmIEoDeVUH4HzGxh4l+6D1r0rt2IejL
PHQflKTKDdfOTHR8DkX6Waziae01BRY3RKGUrKHsiQk6rxkU6Cax3aoZB17l7Yw8
QgG68uJzbYEk5Z0dd2mVBS4CyaWSlrk320iamGCLi7C8Hj+jBQpuZtnC47LEttbf
Uza/muCo6xm7bkMkxP4MLEBbS4e6nwJUZOI+EbZ4D2tk4pZMP4UJgawFYlHizatT
sov9S1NKCKZgPtcUtK2/7cjlHsGjYKx/HjGg9j2jgo3fic4xNf1rlmn47c6u6BO2
YCVaT0CMunw/cfYtCJxmKPV4rnNpL/HRsq4icE+YoaV9YlSP3o9HMPBhrq1r1xwG
Eq3LVtrdSuFxdi1DLWw0QSHaJKdLxsrsxV92PaCVjAS5nj+zRQITG7502mVxM0TS
bR7z4ggZ3kuKc6oyWr+ufbeGA3F7SrEdy7c3RpwdPGlC+NOFofwRSCreROfBmmcS
5jngwS85mNuQgKbsca7pr4kymy9G5BNOppVqatKC9pOqCYgY+JZkoPAJcm+oDZHB
3aCa4Tak1KYXYQECgbCdAPNKs15z4k98zTNTO1yNTnOUnlUsBFMxAs4HXCjgugMg
tKTpzamNgn/YsocVQMMbLVgkOU5ttsDo82TJgGsfnEUkT05Hq1VEYRNIhxJC/R08
BYMTqbrDD1utts/vyvOoKUBpX/HvB4aJhKodEUFyQyYmHKx8ofwyadQOWp5UGbqP
FieXB09nNaLBBsSOJQXUUPgFBxQMWdKUZq082xzpr0KP6u12CFrt00cwRMdputrD
0ZdasLozYO6i0UZAtV9tqrZRfycUJZw4No+QZw4Jn0XmevXd+5wfJYEeGX00xkZl
t8ZC9mfLmbbObA2lGHOj1D/qouiqtur28J7gCr2ZiytmLkC/XjaALhg+qGnM/tE2
v7Wb7SRqOkgp+zjAjYQBRvy9IBNdy2r1VUa8/uzgWouso468NRE4B2/tMnNf+rlR
72nZwb6mf1s86rXPmLK2ZgQxcckz5z1TAO3KS5DAIDCK5vUgPh794ui/UGfMy50H
1FyhjTt1tLa2b6l/wbS9YrkWpMy3oaRAgZg0xRGxFAyRgGn0XIpj5KEvyCKTM61r
JPQ7ALud6rXfzxWzoZFJ/sNoETvENJw7RFAAeXTJCQ20a/fBLdxRjXhl3+cEMn9y
LqOKXdIUhoLzPyQ3liTJi1S0+YHKIdDvJzWfleLD0EEDol8oy5HHKEJHPSYGMZDU
oA23COJ1LMEzME0id4jR64dJxyvSSrcNt0LqtFzhjn71gWNPBWkBaUJij2eJD7SB
W4a/mOoFMhxMbDh00M+sNR7z9o2ux0pc0n1vkM4Z6vcj36MnM6UfxNUTJRJGBWU7
uAkNIqDi5LgZOBruwP9iExtizZyt8ZuiCNk+v2OAgtWqP6OhVuPjwK1HF9fDQgsx
+IDqChOuYIcZ9N8kgMzrGy67Dqfbs3ZyY5ujvAAJTRbhYmPbHXNqa/hhPQruyz/r
K6zxwh7JDOzdcoq6rucMd+FXf468vm4Z+sCNLRNax3tQRfNlYTVZNxjTnzoaGFXx
HRl9/+Dob3bgLUCbDfwm3Zhu9nvqtPlURbKw0xaIPfuRKPbUC6xKImWRkC4pfmFo
NdPnxHGv5dDGM5Sb5qOBMmxeFnGi5LiMLA90siwrd2jkrDTYWT66dxd2CzRDyCxD
uYX/wQrrEryBM2T6QJOgnriVsRD73+t2pgv5yJNJrUvvvW3T9F1SHlyyAtJZsPec
9gHQHBO5VXx5mdjzhcwpkThETxkS9xc+A1zrmvkJCONJ9Mu77juC/YIIUrAneTkd
jgdtT45giHTfM5uMQ5lRL9zH53qr1e1HHkb3BL6sBuYj+xWW//DncB3YctJbmMR/
N08HeIreiJn2PWmy5B9EeOZkkLweEFA2hUlwsHeoG1obbxqsDBNfzjx3bpC+qmmn
VcfGU0/K5Kn0UzzC2U48J5L1uBQZTf/7VqnyluwfQpBZ/HS585gtvwvo6QaNxPPg
WNoOd7QiHQ5YLG0Gfiu9xMBsfHJG1Zg1VaL070ceFa48ICFmC1xTX3/HaUc6olzh
XHAQB1Jq2Kunx5xe05UpDiWe91qIL9W3peQztJiO+sbz670fYfFkwgRPkoa1xexM
3BSLOOwepEs0xKgmHBlproXjFd67OFSLB1giRYVgIJ1OQ+CWsUhAtu3HZEUkULWS
UccD1u3mq9hgvwNnIGQncZuvT17WvTGgBt3otlzdbw9xhy08z0y/HbK4zx1uHMTk
tHWznirZsA8nBsKXCC2hHtkzafG/071E+ub6/mEi2KIhvaMhpWvPMBQX9NJi8n2G
Quxa0enEu/bfiC6ZZAsTLTqYafhP5EsYFFQmwuN5iwhgp8Vq1yx1mBklV737z6XC
M2hAqIlgIDIVuxF64I25iAuOPjmcghL1ltDlLRi0eBhnVeQW8hxzyHHO4UYlz8uX
ukTX2mgJB9G9LdaPp2u3cSKUQPjyz0YbuxPkr5YyRwrqzeIv1nVegEPOGCcDyCFI
bgJuVMUZmHwRQOzuv5QySQDpHL7O3IDFIUuO/d51wCUJAyWDQjMg8c+eqjFb+Mti
Xrac/B65ehLSQBzgwj4I2U6D9H6bkCVNdch376Vbdx7Mxo08RtLs8wq9c3NCPMDH
pqzv1V82SYrM1hu3KO9yVwH7LmIyFxk8hkVyuEWg6ol+r6x7/nIcgthrdhTUnoQN
E29lCyiGLKGWHPWAgxgjg03v5smVu7o0bYLz0F+WxFdXzzxuttKv5OTRFftSXWPX
9qr/2+048BqsZNAovKkscviByZiwRg4pr5PlxP4OLmmyDe0TRIQb7xovXzxwBCHL
/Yd4TRtrEnHiRzp6DJeRItJyXTY1cUauuQXR4riRYPnOAKPdW4XGqvsKAyHTLF0w
Ldrfn8QhhADv7Whdd82eTorwwfvmBJoi017ISmipxZ3TO/eE8SVMuPQhgjq7vfYp
3PBMfGY5mhrVOsTSQisV03gSWk9iHqRyGtIbz5CRqHG/2I5Tx3aH/70+OfJ7OEkD
H1QRRxEFbqJ3iA1mV0JavMjjkxald3dWp839/LTs735eMzFwzjIWAWHUtSSTXvky
lbix6YEaV0cCLCXm85xpufX7JDO76/GB3Qm12DMjqErdbQOjv4DhFuZrdyAgzI0Z
Cyb2toXF5SEZqCtIA0tm+/axhs1R5YM0Zp8jtdeBeSiYbmyd0DhaRsMsewC2fzTy
OSM/tRVXb7ZG76WObzR2WZ6HYbPWCa3jt77t2SJ7DClaJBsd/RdrcjbdZahEz5V3
mj7dL6BO29ayIFIMEGEhNAjeOLLsB3WXj3WByC2Hc6yuA+2qTS/6hJbvDcXE4aR8
XZc39Opvy15vtTImN1bjup132UDtUdQnkhtzksz7MLti/iSL9d0gviAwnWlq25o9
/pNlUt1xZ7jysz6ixra1i8WGM2PSeF+ZTlzIol1kzY3JUZYwT6X6daa1ya26uS6o
1yaxRo6Oj/8TCuUYwt+fGyyZm2IpmsADj6DEEdwokEyuxA9HcebnUlaznh+4XMi7
nrHAtoN9ectPg9Jp1U63y5lH4sluoGjYAcfBpKKc7e97LWXqfy/v6hF9DaGPOvzm
EMSPncavKl4cyYNX+pq4S4ICTUklPDndBU4gCdtrToOzTNmnA/0FpEsOpFyEjP/d
E/GM6CdgJ+XMCoSO4ZECJhT/r+Ub6rofQEy/1ul87PaCQdJECBzmM9ZIQiuMVOux
/1bf8nd/Lm6rsrLLAf6+6LdNQIRD65nab/KI5bWhWzyUWu8T1XFa9KPkkynjuqN3
IoBbKBzxwagy5n6sWtpNLgWAC2eYnc0hKv1LAs49HFUYRryTJarJohuV0zVSIWBc
kUQvPz1N5ZhnTwAe/MNjkytJEw64AtJ2x6A0F6qxGW0wwMsTANtKIjrGYq54uenV
/VfWHGaXgwNzgJjh558x5zukjZuGA90YVQ0xDzG87k4+otEBH3gG+YGhqiibBatJ
b/zHlFyo62NIcjmOeTQ2msiKybUn6ZSItqd19gsX7lFHhGF2I+aYXbQi7LRvY03c
MylZ8OA+VRF2QJZDRWI2KTuCXeaglTBSl45uutnzgEJp+tkDfdbhRElF0HFpMPxF
MWPO1SfwfRaKsyIaO6z/teIW/525PQ+GY3dj7A74sYd10QxvmlC+Ap8QnqMwvLMX
EjHYsltzjBH1rExZn74sl/BzaSOSemNU2a0uOXeOWB4E03tGcyWpKQ1t4nN9LG8B
RZqz6G90CecCvnnxv0pntWlIdOontgu37XuhCOHXLkResxODOMhbiD1goBwHR71F
K5FoXY5cP+Q9oNrFXOexVMhvUD8NLGXlsmQWeFwyFm/2gUghEDkfLkXv0gCrdQ9X
pADaPELsZoENtnylS5jleP19SWwJWHiw2TqaS4xcnDm4IMbYB9nX3EcTwcj7jAtm
plKcKVXtPLiC8q/Ukqoj7qAoNKrRYdTkVI8vxPtVCyhoErpavKLLNGJkwd2IouZ6
1qAduSi0+fscVx2c8OtrMkEd1ZL0L9poYWF0wTXMgNUZJT90fCHRFzxS5WcANNFX
icl7fo4ow9gsHauWN7dfSCltNCdct33IDgWsasLx7QqZO3VmO0CAKEJg0jEjpiVa
uuifQwBUNgUNb7nzvXi1+ddk6cVrgVIK+J4bH/0zdIC5gobdgIa20ML2fCeRMVG7
R8RoyD8Znm+0ZjJQQIqg66MrgrpBAXzaROcHjIZzv16C8iYsOljcaQ07bNmaMoL4
6fxuwzLvN527IS8OGPIoBm5+Ox+VoU2m/dBOTUIEIrzKgwyl1H80+bXOgy3nwRnR
3buPyLGqXGfD/00p4jWhA4dRz4UCkRGJR+93lhYGnGFRBC2n7EtKUDV1bZIGPpj3
2W4knCQFynphbxgNjDWQcMrOhAg2uPqxy6c8CUe8UYSuEZCANnCB5mudTnAHvRCh
6KsENDMwosxCdE9PVR/Yi659hhOiEmK1reE3R3+LqKZdbHPAUpYxgc0BCPuvq1Tf
glcyfluSzkS0l6VZ8hU0u7folMQGDId/6TYVDTVX1cB9WGsS2T38TAlm4UbOxr6b
hz+Gf8lLugGOoVvGuWhB9Z5bgW/ZLSVj/Mhw+rwJn/ffWB1CAKOUVpCnoHuhhvQm
yIJDQOxRFEFo26zZCMkNMOSfmGgDWDf/qSia/0LTSG6CF5OaPTpFPoiNoBd0C1Rr
AwGov5AMrOuUu+Kc4Gl3sFYvUTLN0Fk0qZfzuRfMDqGO4Ks1Xve/DbXNEfXufNQW
WVj8EvGpfJHEQCP6fGXGF5lzUQ8KihSjHXeVgkPGFY5z1m+cq5BADxyJ//f//Otx
ksD2SC7cOC0jTPV9M0JXe9ygNZyzTqTdXrUPliREGkt5OlVw0adfOk3GPL34D0yb
plxmQ42ddYlhr1x48dMH/yaC+SdEvyUFUBXT8Tti9lWoZhlX6JtJ6Fr/KyT7r0bz
FzscRdnEryGVYaq/8Atd9lMNk4DD8q5rRpfUduagfA348A9GSmuTsYCqyO+Ge7/r
qUNlk3Xnd6RkUlRqBPYo4OfXv/Wnr9CI819iGndyk2TK5XnK56/lwrTxJs8QgWWV
QrZJDBCZ0IQCesSH3+UcaYGy9P7bCl+9M1VGX5M8BE0zm6rdcXSoWG56AIoG6HDZ
QDB51wG2eZOptVOw0hdNYnyq1XDkTx2ZufOeOnxT0F0+d77zn1/OTfpj5Rkgl437
QU5KNEv2fBb1EgQgoETiMID2EPWoEH0arJnevn8P/o5zAVBU/EoNvtFlyA3Krwrt
rqPHJvUWLlk9bNUc2Hok+JWUFhNjR7rklkDF8ezTTnUk0SIj6tVbgz/IpEVbb+gP
rELe4DwoJD+0H+zw7P5q/cWp1my1lyCh7zBIt2cuX4Rh64iPaTHDV2VYDdBcjkvU
1jcujjOqUfc2OGxD5y8utjRdig1DvICpoqTFz/khADoo9VT/yXCX/qZeBSJT/oKW
rZ7EH4YX3ZjqOELP9Egn+SphTAqzFCPqaQVn58OXwV67CFhR2qI5FxJ5xI1aO7N2
OKwZUvaL1bS7P9WZR6rr++IxO6Fa8rcbI1SCSExQZAVvORCILxYPEmN0Chl/QSlp
pViJjDX6LxveXYFO1viduDgqDyCQxQWIBJUd2ZpG3a3ztdw4zGlFZGJC0B2Zt7JG
UNn/qCHoGqFvuNQJidAiZSP11rKdqO+uVR91xqpXiaxfvOMfWQc4nGxfVpnUz72w
eWH2f80hv992RRWJN5u+0pAdpjIMPU3SFdbZu6AjVhjpaVMm3mj9gm/2gQn/p+Im
lpJGDPtgZhWOYg6a634Oh2pojmxAXU1HIW0VPNhhRNHFcbrJSUjzAQHWW6DesKc2
oHdi3W9xx+wTxZsQO0I7jeERzKCOTwlisW59swJrj7Mt9w17uMreGqRf1yHT7P6w
dtppbACeJVXZyzlkfrL6ayu/T0MlrkLBRrOIFfGoqSItnRRdnOex1A2Aod1TfAVM
wlbvpaT/vh5GGWiM99FhMBZgkE3sIuwxo/HEWJqfD3rNjt0OXM2KD1SBbK/fe44A
P2Fg2pXzTx2ldlOhvI5G3jDIC4uPuON/nsMWqHtw/d88fUkCTebhP88Dd7JbBv1a
38aiSZ/OWkrBKpZXOBcRtD/sw4RUL3a7QgSx0mKDY7H81UC/qgT9ZI3NbATQf8Re
LKm85eRSaDMLvKwmdWBVmfqEDpugnH1Kg1JU0GhmIKhHY27E/GwH54/YJq1usVfF
XzqQBqf2m074qoQ2E098MK//9coWfE3x8YY1MNcu20cG2VLWChyfLb//UmVFmHfm
YkRJkZkU8UroQ+v/M0SdUWBJT+ajdL68ui2jEo7kfABxg08EAlnscb1GYju4C84B
45HmwJyoqaN001R2bQyBvDLeSXmeHQ5i+wvoy3+P02f38W3hliCzDsbxDuIH33KA
jydQgSLHUg1hg5/kn/hwVdvxcmZNtBi8rH7B3x1SXf/eLK404oIjlmAaC8ATFWMj
PuE0L3uXEyrA+0L013n0fcLeutUtP/iLSei0y3TOshj4zmeBiXhrdA+SIEJilrUz
mYguEJVJokqQpCNF1mEMgXPzKl99o/G+KTI0gwRcNSL6OWQYKFMqasOS1QRnLx3H
W+I7PVcFLSnzW/xPn9N+RWKIOYggD3AmwbAQlFuoBGCk1TD4dU6wvs9NGySPdFSK
7r+qkylUd/R8M8Lsi/qCzARVxmqI0VjwTNl6W85+P5a8gATWw0WlPtSxH+eRQ9gx
32UwLTCijdZkD8ck2tj2BKsm7i776rfjFyjz+Z/4sN8VSyge9zM493qXqemA8Cs4
e4QnK4Ikp8DHzhLPDambiVdig1aU8d1mkaBOZDcYKgLvvZfpL8wVyESlsn42Il2Z
LimiI4zvlqVcxAg/atMUKYzDEQRHUYBvelcHVnoTGKqE8lD6H28la76YhLRVL0gN
3U2jY7DMZ6IzD2QyoIfnq2dtR07y07hvx9/IenUF4YJtJtbK+eATql+MQnRsQzeB
eG8oaEu31CLVF3NaejEeRGJm9RV00yLncVd6aYjquC36wtHS0AW5ShIXIQabdR5w
OzFVKXHUddY3fOP9LF8MisITny40nZfo0Dr1b9X94vyVUSx0JZ4/FGCmhkWYFlbY
P50ql8kOXiYjgyB/oztJIh20Q4yXkMVaj0lqf+rhlDaCNyieA+BwZhqwaKSpgtQF
aCfYUW/98QfXiZMZ8fHZxFNM52GBIY7h1RQDo6+XUKGYupdOzuKFUkcHNuanZMBy
DDU+K+OytUKJqfj262GphNiYYFwR+v7k+VpT79/lql8TKQIiEGUWCl9VokAiaaR+
ResvS8b6rdPg0LoNoTOBNEitEBVeZ4UbITo5SBvwMHk8xgQGtyN9AMswzr8sVRbx
8FzrI3MVjrRLMKVsHCMc9JLsYcmMvYZh+pmK6djXSTsdjlgHA+52dyYhLMMs3w7n
8UtjAH0OgQ3DdVwAP/PD8IqAgwdVlChj5G2DDoH2drsOe5sSr1v026xiG45HSZrV
7n2pj0/7CgjIwD/KJlO33LfOlXpX8sl2UDEgL4/ZHheOO6cGcwScvgpxAj2apgtJ
H+K2NMyJO/f99xOGUt5t+Ayi1ortGmLrg3XWwJvgquThzwajb2Btj+9teGpoQP2m
TwsNRJhVrjTC7b+LoKSE13rBgXEk7nzYgXxusH6yGQuXC657sN0uz3Z2B+8SgUs5
xEIXj0PtFY17EfMI5KibF+K/gIwI66SNGmN8jrZaUY6ZjMMQMhwm0tjpJU86lUOC
vTx86LYRSRWmXL1/w9X7EEpvI31jcaI36kIz1H8Ez5SaFODxM/4i7h4z+YuMbdO8
tis3TNvS1M2CD9x5HO+ST+YBj1/XLmN8H/MeFWzGr2BJVouWqtUghnSxXippqtUz
IY5b7lk1rUFcefvkW+eIOTVPUNUDNS4GL4FhxLkzEGqcDfg2crAyfYeKn2317o1/
8dSYKhv6yiZXnF53BLO9nmf8eLe9uEU9e9Kuh5y4ssibJohheo7C7akVhlpwV2rs
H8+BuTjP3BClkaqhuaFzKK1Jo4HI53mT1qRoDhM22al5Cz3Q84XDjiVhtWb0BEp6
RDbuZewFuNp0rykgbPzDodCHlSOqvn9cftj+6nFCjpD/XVArUHxG69fH8zaU1ex/
uuJABpDoE8bG0u4XN6+pPYdTMQ3d4Pf2dvfLn9LdRbFTx0pCXnBYpe+zZ4gdcLXs
1q16blrP27yHAMn0+sOR4hRPgqztJvpV55lJLRXOqKpf48E0LHxc6C9TWTZ8T0/u
o+YokVy5zFQQBF445bPEH/rZ8AwxaADxH/Zg2eNJG+SuDJ+6sAD2GimpBAlyBk1t
QkaCaMj3yCH/KFmbP3j5oN8nbNd4ub2lIBGkR6vIREXeVT6Zp6glmztAWn+/7aOZ
4UnL9+x8ZJgqyD0c3aq6hojLT4FkVH64p8j1B4VuU3Gwp8by2ccFIeGR1+dNuneK
VGZnpWmH+exwo5le4Vt6U3BjiffShVqFnqPYpTXbHycu1/PqnlXKRkjY9L2NzlWJ
fuHeTYADtK8WRDq89SJcF7csuH+/vi3UPwT3cDdtmuJITF662k31c9gAamk7DZW7
57sVHfE4Wdm2Y9cEUr6/Q+ijkNXknnBKR5qj2xHbMxRXhIWKfwrqVSEU+UUEMwBU
rYFa6+X3uT9ZYFa/W/SB8t3RvMaRuXSaC2O57SWYC4Iv7HO1yKX/AFKTSRCYZlyT
KwFiFf5lmsl8erC7lu+GluH2iHHxWgb5vqhtNI+OozMEIPoDf97Q6vM96KH6nx0H
YWpsWxmT2hq7TPSkXst0ZTPwsvjvyfYjAfcuajzuMlbx6uIPoYxFxxVacrJYXo23
f2PkxvO0K8AtlFiO6/Fhz7y7fSkVeuDD6PrIq3MCC054nW4rtdXLYbSOaKbeUEnv
XGlqf3jubOTZvV/E6YW4m6a/+LEaGpeWgHPbxQ+6pAezxAGgSMW1CPgeLQInTwNo
Tdr9iPjRAvDdOomQsdOi8nfzPZpGwvZJfO03/ncr7f8StrPWrjgkY642lqnUSPBQ
QoFLzcqUxERbpSUWcSGqkr4RTjuuYW/Y9vWi0JX68oFDkwvKkx+pUYK3AwAZCYpv
hhs3LvSbnZ+E6ylhmnlRllE6me4ZX25CCpwFw7ug7+6m0qd/Lp1jQQMuPNyMI4S5
Tv7ZMTl7gMeID1voMrZJ4GFPbNnRSq+Y4flzQuKL3OMOu64feruQQEhe68UktXPY
w/rMX08oZYtwhi+BhL7YUhft3Xtb2fI6KZ+3qsKEV9dpEHr+NDQx6A1XZNig2yi9
71yc3laL6bBIb/DcA+kmsbREc+sSuk5hGNzWM7UhLjX4h2WWBVlHn1fPuVjSfTlG
I+8Axm5t7zd1B/D5CNizmew7v2JgOCp2bQnpsEZEGk5JxQ8/1A7zeoJlhHlmqltR
syPOk4PzaYprcFKvWbPi+LVlWUic6dOTQcBRl70QyEaswigfUA5cFej0SCtRDnyq
ncqmzQhj2ivEHKoPrT/N4AUwCPsbMsGAMGxRMYfWDsxPj97IWZrGZWxuv9IAEKk3
mAMGiG1jfrJgLs8NfHV1oDXe1RBmSlJF1XJLEn7BFkcn3SOVBZH7RwWvUP8laIMS
Aq4WWt6MgJOngi1ZthWL64ZN/vGnQSZKSch9gwytFMz0KwyzSYMbLqx5lv54c6x+
9sO7wIUtiJU0bNJ/zX3lDs3mu134gBL6Pd6c+pC/Pp96Y0Vg4f6lPIQGpI8+fjF4
1JpmM3bkHUsAWaQQfBrZOOElHaE9fRNGCRvwnxk/TxzIdEJAOoSCXA2omXpMJc2j
ZYoOpwpAor5msqUgHE8L6v1yJJNeEKGoSJGDwOrSNzc6AY5N+mWZ8ADMOt+BkpEW
2/COeQkL141USB9OcS14DVtDzferHDKtKclwjMViS3G4LeNH+5p/xAdWfPAJvg7g
8LZib6uMH1q1MSWn9N9qdn2kz0l1yUrZgNcNukR3lKxgzd2N4T2ueigpG5Pcb2sf
ZQ30DsCKNXufAnB4k7sWiZ2FEbmIXZuGKHJSmejuCUznVfkMSPxsNrsu4F8oU43I
+9wMDcQXly8xFeIPcUslyJkuzpXxWm93jVOFsA7X9kEpMxxwFcHVpG9+mMZZd5sK
XoEw56VKQYmdTDJnCW4eG/eA85ey3O71tCsLQ8LmYzDTSKppjYZtLXG1+Z4lreLV
T9dwi5RWQn6DOz1UDW/Zet1DP/mcZMWn+Oe6B/gXS5hka8fujDznifQ6+i3MdvKL
oxbR7dEP+oAUHo4p59jKo3LQGOhjIQ3uMveWKD3WXYeKvwklXHescdG0krQk9+nw
Q6PLY8j/J/RLYJhnVEY775LuPn18aAYkFf8CMisNvqvwk1TRIE4YuLIrw6nzVJ3+
+BjJHcxZktrCVpZoip0sJ07AZZY8Chr7Se1SxHP9KTeOfvCaJFsZVZRGoc8oq+/R
vtsM4v51p/6yAYtJ3eRWr42D/YAqJZFX1+vZawXHGZ8VX+ZUzQk9aJTDZ3i98OeG
PD2Ax7IjXs/RahLOGOB4Paj+I8dQnU2HbMrBK7m3zsvyMeJq5jiIgYro+7LlS3Ep
ns5pzUxEDN2e+1SGNcKpITgHsWNlYc0+a1cZa8c4XGgd4cx/OVlg3LYGV1HXPMyf
l7B9Xah6yJecRASkImnkX1zUy1x5Dzw7XleB/+k1NS03WOlJ/Mvq9XmhI+LwEUta
yB6v0LBl2F69mEWFkCies3tZZdFZ0kHGmiRMoEX0HGLOv38gqoBm23jD6gQ4IAJg
Qg2PkgxqMimbQZ5pA9wqGu3KkkyRhngVlMzK4Om1KUo/YxIVTtDbnvm+/4d44cOp
pRrbeC6m25ZOG/iaX+8V6UWo7gxU7HYVSWmQoOWaU6a8t4VBHqpRIWu+wp5ZyWcT
RZF9cgQ1yOv8nvXgXhc2yejMMBlXq29HSSpPg1W9ehaFhkYO0v3wVE7AgQjYrsbV
VuklLbxr0B3fAjKr+lDNVOq/377CSgzmGNFa74ELFudxkbZdhf3vzQ6QKX+MuK9H
lZbwq/kafm67dBYEuwNCVKCmCnBYei8TsKWEFJabCAV6UT2XnN3YarIOJ4boh5MB
Xp/PDdNfVMTfaF8h4fr/0zJKVy76gyz1t9VDGvaq32QXKISKOmt6RMTNW1J8WW55
1TUeZurqe8xN6k/k5yfYIqtCAi1TP4/TY/Jpr6TiQHG74+pNUtUskd6qdKQwM6qq
mPidraqkp1XRPr9L7tMYf36A10ADq4Gy35+cwCLp/B20uQVkX2qIKzfI9oXkRT1H
LvPqgGaA8Z/XuUGx4+jiYIyMs+zyC1Zyw3BVQx44XqHjNNJd3qn9RCZQ6Y9XcJDc
Oa1NysHkVXbgI3p9rOjn2t2yCighMBzteb+j/xDd7odBiR0wPQJQaSbfL4mRLODi
hQU9ywoTPa7rrJ0KrWOEgGWM6b18YqEeSHFM7M2CwgIRe2wj0XXhlbWBc2YGyBi7
EF5H+deTP9T1D803QgZF8ikBZgFu85BDUjlA6k+jwZHjHKQW9QIU9G8G1aRHH/C7
+UpX1zC5q5TwF6pljFoBBb5+XRTu1ALHvETa8A/vQtN5IH13xDf5HOvOlEqUpVep
Qfox/ySGJEJlMHm1orfG7DSQzVB2MBQdGHNnXqmNgPdTAB40xIsRojv79Bkn4lWU
1LkhAz9aaL8CAVsHjr1t0ymEyiHswk4/jtEL46R6jrrq8STFNU8Ggy9LAbL5weRi
oxx1mEWcyzLrodT1bnmfYrL1r5VJ/jN4B7geDmE6Ca/Us0/kzJLYCg3Wl1XgAdGn
pO8garZd4wqTLjH+0kh7AovN/3n5lTKqQOpjEbVZwOJjtrIHj02dhA7NKWqtpACp
l8h7avgEVvBRzB/zZv8E/KAtqGEYfchcFYxylTlK4T341rcHZlPTPBreEmHwzora
5r7WQ1bVxvOzU9wRYO2VoyFFDOUOVNoFOPrWqjAnVTmrmSsygnYY5VOXsaypGIuq
akdQj5K9Ie35rt1+VwEQNHybidNbfbi++5gQ5O14edvrW475cxfzGCg8a4S3wuMs
L7n8RhbUtiIFewV/ldvoTQxFSu6NvAPgOrCjMoZzpcnQwIms4T5Idf1+Au7/YTqO
Xqvw1F+xHgjQxBcZNnjUHD+bcE3wrXIM76kE2qHy5kQNw0BP8NSxQT4zCky7/ESe
hRK87e9VU5rVhHzI1xOWpuH7u23sdgeYocPF6z0il0GULv2aQwvui4dJ7xqk2q1Y
yakIMcUzGN1fAz+MoT7/Jz1EX2iMnxLjS+rJQUsdBAvoAI6zyatMmfH+ckGkf39a
clO+6WoQkZdi+gTW8BXs4t0HrSD1T4+cLRUT7TZZNnr/VZB8JaaKlvZVsWOIIqWo
oZoM+58+Csm7EvnJQjeoGTKjMgjwSwaHbe4pAfl27bxfxDhn+nKHvRbzGyOa+o57
s+39HAo5BMKEvqgseIPbjVDFPD/NhTAPAszzTHFzH7iiYWBbX5eDMcEuAf66WboW
OrVg+mn5LHw65htI24NbANFfcJx3DfOpZ1qCsBtCVdGDTymhEyGJbvCCXbPuCcwI
dNJckl8e8xvGVp3SL+fv3ExAkNaUr6RPRUMby708/xx8JAX3/IahgyH1jmRyIlua
vfgMl3PMHrGSbujfsAP3sVI27MbjpBlqFofICz2qi7z0pLbVlZv3kU9z+kajAdFs
NjtwTRCv2cUgvIagY6Ew7AvpX7vbfZp8ItaixgtMbZGWAtkuG1ZLgHLKkTf2jm1B
ZG0j3uQPLOa+bO1BIu0uzjsXI3XkI/NpDCz38UOuxidalrbLDIYiXsrdh+9PUEv4
J4h5nSpfwhv/N4FP/jKHV/knpnZhFKjIQGxV0Ib6EEnSTFU4Sqq72uRJTezKqPbj
HIwE9q4+d91SulQ2s9MZnSNI9XA9m7FPVIOurtPq/60k6co3VRfW2lShCN6poREQ
sl+0lgEKL3UcI9KGJqfhHowq0120YU07Y2CBz3RUa6wtXN3QJuMDYEzrHEiDtzLf
el3qSBReODdbx02fsMrXN/rukAyvz/npdjICy79a44BCrplscNBdB7ANev1WFWGI
EdQCzVkB7DI7tpqXHs9w5pS+hPWffd7NwEHyLmkP3I85/VeupHxLHooMl4GzXoRe
3ivZsyuxAtm608n4PqXdgLbOtdlWNj8eGp3TDgkbcTRGbzhqW1cHhDhMJyJX2Urr
RiLTHSF6LWEgy5phW3HU377700mccndTZcOLpQYIdQnHcK1KdTSg29jHdTMCz9rJ
xuf6KcXyhH24aNXTg/ZeXFo/2zRdC5UYiFto4RasktZyyiQS9aoZvw36YpAbMHxc
6yqh5pHYlNaYoH1CPO0gBt+uAw4OFocCfmgiX9omgDv81aPSxiOz68wbRHhhUmBl
lrsqMNDVpv25q1y9Ql843XpEb8nhW403f3N2qVxoJvZangEpCZKyWQA8XLS9xTOt
ZCO0qcoq1hWoFvBhiBfhaqVPwoTi8yd2EABhFwmts5cV17t4HcpwlpJ8y8VOHLlz
iodQD5ysCDQ5jEtlYZkPzwmrJeS8U85fIZ9WZZK4lr4hqfo2cve6QsCYCgjqsfIN
qP7vvNFWJ+DloPiq602P6pknM5pjGXqa4IlBm9sDwUar9IOp7bDcVm28R/SGZsV7
Iw3Wk7aXmwowrueaaU7l5KNJrKNvwdCbS9z+jKww8wAZSSJ2KbDSksjbQ8oqYi/H
x2AGP3rhzwM4kqZ2VJBO2oIO7VX8+HEedPu1XpKm9ZI8fCyJqShoZJescOmUORR1
Se/Y26p+/k5zNhqAo0Dce4CeGWOTFzpibmcRgu2msDMbcCD24/faFMAE+q0ZBm7R
cb7X2n9Ko1IOCRVF35jVRLbtPlOMilicKgwFYQQr57OOp2DNZL46G7wYh5ItLHNO
ZfrHMrNNs9MctWjh9NkjnBg8qOXr75GILA6HaU7gNFI9YR1CHhRIdbuA0CvT6mR3
nq7bSgv/E85yqa0lIPi0+vOtup9UEQRHhTF86QmN3ntf0JrXyTfhTBkTdO86DCp7
TuGAKQ3LGsEghc0ZkCd5OLFH12dI5ACGZoZpwY8nljIGNRA5ZtRVA/DXC1J3QxeE
tkZF0z6/T+XM/n8yh23TRQZ7X4ydKHD7cOpiC76sa22RfSCUN/A5rZn0+nNE5A/1
KjpfuP4PKpzPAYQesXGhr3Dliw2xyR10PfzKdAmvfTCIKrTf7BE/YnWcje12hrtF
1d3Hcsia1H3oa9qDNgeCk7BlG82gtUTwduBwS1fYkvMZNyerGwkHDRWAMekT+QLP
jntEzilkxfxuF1fGm3dkwYePebZO3M3ICTpCUiO3UHemErje2RBzD7zUxBYTcROv
v7WLZBqujX1FVzk2OsA/XnEexsm4QkvSVUN5X+or3Hat4NwWTQfNAHedsypDDla1
4AeUwcrNKRwBZpib9t0nEDD52ipTwlGfVK314F6r9SV9TigfME0kdZXi/YIv3OM3
I/t0Y164KyLz8aXGHfQfOaNAnYHNP9jUhsVhgVequylnVeRarZHQIXkxZUbAkJu/
RjOnymUaWjV58lxeH9KqQ+v5Jy66/e3JD60D+0pRMcFURvLYYjikDGmrTN4ib06x
yNtrGKUi6271pGGRpE7Bcj5Y/Z11NgdwbJKPBk/jLqf8aFWj4YAL8PT0+Lf1HFuH
4MomJRLaWqT1DBGHt1rsPUdTE4Um3vz1rHXl1bSci3dmFvo8u4PWASZIWISPS/q4
j+U1hTDoDdyYJslqk9QZNKOZa/H2MMCBPb4dqU1CPzWkl3iXZjfukgMsV5knJbdv
IRAFOD9jCAu+/PD7dhAMarFdwZpeVs4RHnSakq990abU6sD9USLVyR3iq0oXITwt
TblHw3VTsN6E5VPHK9MHTf60C43MFL2Iy375KxoHlLjuCf741RAGmS48bRG6v+e2
pydxqT8lSHfktY+27r+MynfXldvrvIsaTX2HapfELQ9AZE3w9QxZ6ZT6YDACaDe2
yMOo7/Q/ggz9Lb6TpU4tom2mg/2BeesbvvCmBupcmZwWly4XB6xAPltihQEmJtXv
On7EyQIRY8EzfwJQlO2o9t3cCbIpagiLIOy9neIece3uDSQkphLeBPYs7ck8Ookb
GDpSSCbxi7Avl2sjTMLwPFSDuW/fKsBLYWSHgPLDOcX4mDelJzftnwIthFE7PVy7
HGxaeMys5tjT+RAuXS24vxWG1r/eOQ9ucgQY4Bc4lzO4T0+t1vgR4jRpJxMeClEi
mXHl5eNKzBVF3TPYBnDJCbm8EfJV1z4nzAGE4ULtcj2k8IVbh6lSf4fCKZbL+bcq
VePpjQUlZsweOcaAbO5h6y9uaU8hfjdqATtecF8uMRKt6sgcs0mhKaTzYt9C50I5
MAnadaDtcMr9vRk4L0zDul2yVuuzUvM0Y+3vjJ3KpfPNBElsTrBow8yAlYWzQEh5
dXvP124sKHz3GSua5/DNJ6VgGut67Q0tCW0apKojE1NNT+4Y2aLnMSaR7FcSteQM
5h+tdzCdc/5qhKrgEY/k/SQdjpFSp8saaaRejTjBpB7+FMCtyGmHRHS67OPGZPtc
MZsqCDlm+yEamlhDxtqZQX8Rgl2mfY0zqhdaRlRuwbERQAP9iAQjPZqbHUip5VUw
Hq1sVvca61HjuzGCL8z+WIwnq3WWoJrH3r8GyJy4k5W5+NRitEmrXlnPbCz3d6dV
kfLJ5qKOgaooHGHGLgzBIqZ8EckFufF5OkOWNssmYEZP14VFLNuofC43CId6eM4y
ncfdRGj8QWtSjjGAXPb10WAHsgLf+hsF+ZGUxyzMd66Pw4kmOIN+CC18qf9tbe7u
yNa6wvkf5wmmn9t+bvzjoM9uqplamRppqlJAyRDSsfE3EZdp7xhRbGGNZprjN+jv
FYOKyk+73147rlt9wyFhS9nZxIwszT6/NP3KvKnzcX/7guqmHzo6g263H3uZyJPD
yFZkCPZexy4B7S+bS1IRZ2k5zqw/HCEhesVEzBRyJdjw/wt40zbZkEa07A31KFJa
lqGZxk52Tt5RFuwusIbCmhldRuYygzn1BPP+9+JdtyLfG8EBvpCiC7z2c32ia2Wi
vPfFEA+kIcMNmnqOKT/A7qskXIrN3dnkRa9ubhJZLMfBwla4VWryRrF2uPc9teUb
yBAKXJM7E8ZSspeZNrYjxM19i/ueZTW8kSjbzaTdqkvjzD/uGuT6LPCl8flHR2O/
TAdjZGMvp+8F+2CWUWGW1uJy1boTW4Lxxfm8T8dMmuWj7QOxfRyOl94yAi9s2Gsm
QV/cbohEjCPRXD8yGPyg4Q5wE43E4qYaTlz4duSHG5x+28iPAP4ByrYTgXp20GOV
YcY4xbQh2mk088lTfObuK6Ikn2E2HunAGjhU4rIv+wnB+3E/dA/to8D591as/iRn
xDzAmFilmEvKIJC+9CqdIQ2eJmLeFZZjq+FqfYxByPDfobIH4Q2nzEXrLcguY0G4
p+waKLl7LHDOjgRZMVEdHIdGN0meTD0fSCqNnjJwG2J8k/Z4+nAJ1NrZicr81ufM
bEntDaWqRmbPFwarAHFWPThP35vLwZfbFOji2+6AZvJcJSrMMboilVvtw236CaNa
c1XY8jYcYjHN5Pd1odD5hPHScd33zVns+xickGS/MJBJVXHdz9jaXmK4nVzXvgG2
/8q6xVVWG6zlGhp+gcMdxQl25p4ui6Luq6pdIIvQpmmo5fr9grYTMYg/rW8pvE6e
MOvNEs/vZ6w4pO5l9DvCVPeD3lm2Rp7j3ckTdujg4lLmRlWOy2gjr8adv6o7ImkM
IvGK1Axph7YRh1gIqL+4F+66mgsK24+RnBYXoRlOZgIClLJc5oUDudzFvAFf5guM
NGiBjGzruJkPSeGZ+Y8CwDien+9BeuP+Tum6CX+b/z3HumoWenPkLQ1w2BSImOtU
V/yiRqiTtWVNKQWW7G35QPzJL2TB46hMSvsvpjWCFMnjaTZYAQIljWklce6VYqJL
BxNCHAuJuEMOlWdX54hljkqjeTLrRYvFrDhNmljBxFQQPbkq6OaVwlfzAQAWVU/9
uG1O0PUk+kSW3Au74pYNJ1V0Dd4F6MeD6xUSwwuZl+GssYjCKwhIFZNqXIw71B4O
MLFkXF1GQntoSS8PAUlc+SGs+u8tbhHA/HZtPycCU2FEm3Wn6HnaemN0W4zcSjXV
ntYDGv52XdmHmAN6OYniRzelfwW8rOSJnEwFWfRnA19zPqASpkpmg2KV4mvrfoK6
zkSEShPtiT7rYUv7c8s3u5W0BLp6lYgzWnpS4h+8BFx+JdKqHHdrqF9klMBTEp4T
vPJtcefBH2ScOfPlqNvQoTf+vOA2IDpeFkmNoelb3gsI4B50pHZlYgV9saedpCum
qe6UNWT5a5uU/csZ+Qn0qTdabI37MkVI1lKVTWMqQxtsAnF2LXNZOYqMKasRxpDv
Njz+qkYaw3eOVeRNLERl7qjr+t3J6ize6oSq8HASk0twNKjxTyibzwPwz9nJSBJe
PXT4OyeqwKiztocxOa+Z8P/I5wRtbspLKPHwtSIyKx0pU9lt0MxGFjtid8eBi2/E
3NkL1Ymq/8q88HGQDH4iO+H7TXSJWBL7dYQ5DO2ZbdVNP5j5o3Evnii62xQ9MkR6
6Bkz10vPUtUsUwGslp1dEer4ArGkyWBZy/C3WEKNLQU5bfDo2FJrHKJTPNigMV0/
8OdF9gu4W9Li1VD6NfueFL+hK3vQ1G/TUf9mY4N13qr50KiSJTYYFeT9TzITB3UV
X1xudmD33eUBneoF+Rz4FjuwIIIPZioVWRlgXxs039FJgMD1AC0UKba/dbUyxT17
2x2+tM6LId84twPdtuZR2czPtYZK8balChj810ktOA3QQA1waEpfcq0S5mTtzlWu
iXM/qxtuIvZydQa+jKEDCpEv0x/MC5kIld69gi5xrzVYe3/dCYPvGVKmZtRjU0zH
TQBbigtvhfExq/ZZDfCtWhbL+VRHbGyLaX8Nytx5nugasl58PhIy6MNxPi5cN8Zt
8XeaYnxpTt5i2jiV5YItkdvhRlaFWeagYvexplEXfiwVHAZdtJMqU69xJHfzUaXV
PjYdUvLB/T87L+UO/8LFVLOr/KPEWD5a0DhAgFh/2js3TEd7cD587Bm/eGyI93gU
UXnkrGJSU+ga7u8J3H0mKTiMZxCfG4tLcQAfzlV/XCY1r9u0/hO9GnUO5B4N/q0x
hHEw089OfcEOUWZHShGS7i2ap1AXEO9tJY0lRCTMTrP67dEq6IkLJr3+0J5rHPpP
Q7GGRuDtDcRTFd7XcDoioZxy1ImhFNQlLDFEgcKQudZYzbD9do+oq4Gjp8vyZ/rR
4uc5VSq8Z+GaAlcnf14MKWQmv3iNPOEp5ULuYbKXCTGTJeH0WI+QC4JlaxHzirMq
AezcTfSpxlGFab3Dq3Uw0r1/FV25LS2HSTXawNkb5GA9BD2HZU+Z1PrWPJecgmrA
QEqAHkTDzxaCif8UviWLPHAaaeBxLgEI7GKftFgsV228o2sEKs5GUT+46PUYHqFT
zR+fa7HAZdJrecMdj5GZkPUpPumABqmh7PY5uuxT7wq5S7PBxshj7wwaSRXkBGWN
uwsXt6JT9a4taktBdOcuVcrJ4acUDNhjqjjy6oCGuKfZ2ZQq3snoO7C9UcgJgnN0
v/oA0NIO0a+AaE9W8DL3A+BI4MhbDnhGWuTTNY2hFcL8qpX/WVugmEjzb2HcIoCV
40EzabZnnhShRAy87UNjOG33cyOy5dPvaFmzRPeQRWLvZVW/qsc5BOGhk61bD9xv
UQGPp8+KTNwUvgf2Mn2xBpleKyKdkzx5w8QiUe2Pz4TNXSavWW7F3jBgfH9zv4k2
MfEmPHXnZFBJLP6mNLchscpVPOsPLmeOgi3nw73hknSkRvXu7VN5T5qgOCfRiogv
rOifUHgR8DiLZtHz16pHzZiiDQ/NwfZStRqghiyoaaUq1VHSsQ43IjfW8IpeM3yX
TzGINkOSN/g0T7VXCAtSwOJ3p156/l36+5En5OZtgr7kWDkeW1ZvA+WLSPXTXtm9
COUhD0pEWGaSipD1UcjGk0LIJxwhA4SWceokYKRbHI/pL20gD8A9F7bvCnwBfQ+8
a1F7xd2lw3ql+DavLnyWRvpgM/WW6F1C5EO6++Qj5F2HvVErBmruraxBwD2vq0Zs
i8Xv8aK0yUkmmwL9CpgQEdKYSzb6s6WR5bHlrwyfChlHTtUArvMP1x3jeoYnyG3n
IUeZ+MPhH7XXSzDJlNzjtMW7JKIgYdQpnlNbxFWN3SM50tQXZyrq7RqoQI1FE6Zw
+9dTb7RUrpXC8w1OJldNFKFCGsCruazUug9bodhhYCKX6QyzFq9LtnUf5D4WSo+b
TSexhv6OTfN9LjNS6LjNnNNqQB97Wkk9hwnYKkOCs7F8lTgXqYwf5sdyl0uV5CnZ
usSgX1WTiODqN85CJgnPds8If9Dn/iSpQ4t8IhJipNDJW3vAlnNjhDWkxc3Ui1Ix
MZZV6PmNqw2i8ano6IKeBWY2xjU6JL0C/Q3MCvntayPtzAonK6rmWEfld34/rJrw
oCFsW6CiSevx8IC4Z3b/aZ2ZFAgm4/L6K0lZdiNmHtq52O0kWUNvOI28t5uGqTUc
Okd017A057Lzvpi4v6JH7W0zexXXaaFvjNDg+f8ysjvAN/+Th5nz7RCmoCBEpzrf
Bl79u93XyIKXKKoW1n4+0MU1PDYEEM7QVzn6/ZgsUiAdFWm/Wa5kEddXbjBluLpX
fT0rt7I7EINaUU8tzBgnjxfJVAis+Q7dE2vXiZKYrbpabizSTkzXGtEyenA/uhYI
d2VViuzuOS7ZiiGw9eiXkfbyo/ETZz7vm+e4Ys7gLnaL/tMlHvmWgYXzi6YU73ST
IjftPcjflwhbFRnZGteDKp4vvA2mVbC8x8q282jgPJ/Nqb3U4J4FigCxRnAukC4N
Nqlk5jyx6NI/32SVA3iObgpC8y7ceEgZaF4gCeEqNc3nI/W0h1h9ZmeiRPQygIOn
UHcQbuwkyDUvnotmKtWyskSR9VfRTozWj1AClbW8IxaF2BtUWA38KVapTZrywVgv
acNG5l0LBOpew1kmZF8XX+of3TpRgXmnFRIU1G1+Ct/0v9aIJXiMKILj+iPL03sE
qABrmXb+8KWMQfDWr123qpcLmyx1bpF2ws9Ki5sDvgnBKzApPjRusWAkyzlGINXu
XGwjIIAf6fl8RBlNPH+ln/uP9rRKhF6Lhaz1HL9FOl4awDGrga54JUBMl9GTCBm0
OSFArxRHVaW4UO4dvmjh7jgJdOGGsyNq3tqbSzQvud4fIHG+InRp7Od2Fah3CtAB
O5WET5X7w9A6YqxsTO81FemXr3qm3YCWGR6UR7sPyAgkRItBXywuabMt/R/UueDE
NgEcELu3KjtyAgn0h2sm1mjtdB9ccEarbEFFn7KrS6/E2aCqFtSEIPbfYSii5Icg
rIt+4KdhKdF/goFpSlihmBWEm3gzndvXJiCgc71RtLIHVWx4znm5f8ldX565Fh0Y
fXi+9kdrPMnnJ3hkoha2S8ms0boqenoUhLiEp9MenEez+8XtHiryUalf4fQBBKfp
LVU8V6B7iKYUd2JtuJjIP3vhZB3Ouj/DepAC8ONusAfU8YGlwRESuL6s8AqR6hCZ
fQZ/WjLocxGrEwt5AOfza27OhIM/XP/l1TBM9GkiPbZd8rX29fZRfonaucTiqlvf
z76PzYj+kUc/eWd7Xs+jdQ/k6NE7zEPZNzFnFFD3SybqJ6MVvvH8wajakJ75DFHD
w1k2z+fpkhOLh81qM7elR4OommOdUis/yer9GOH4FlJ+BJPF48B8L3QOd3f7ueJZ
dAGinD7FRlz5IGUdjbYY4wgMTC1ePqlhQjowNRN+HNkKSr+J8e4/ydv/y74DT7LL
nVcBHe3Gu4MEN2FyPajAu2TzAGVYLA5CQk2dIyvYU683F0me159M/v7YDOZRy8b8
sUp68tXEIRaGWZJ8ZfDKxPsDvyUQQQpK3/HFvs1qaGKmGdBDfByu+qzc+yO5KzDl
s/COXld0V25ApBpvew2euFtPEBdnwi/SXGaH8zT52wlTyS3MElfK6w53B56lixsz
2LVJWZvyfjekjEc8AI/1l1PEXvBd1lme/h2en7lHvfvB8dU/eX5e3WzpfwK9y0Gb
3IKHYi4ncd34F8GoKh7HZpisGQtw2O9EHP5x4fObpwGaoxRvvr6Jw4oHJmYloJlJ
PyximL2UNumx5Kvl8heRvioaO5/koj3HE+DG+EjUPcac7Ga2OPfl+07my7Hzl1Gn
nUJgUauj5NznpCt4I5l3Ma63KJZIebM4VOJo+dpDqrg4sToXruwfyaQMQTH9pVBK
cSLKlxN/Y6+YgZ77c3/1PRnBPV6cttOqW9NPmaHG/rNC4RZHyicB8PvxCU01r7eR
thpUDUCR4Q0vNdxS1UHQvdXzTfSUhQ3tyM4khEFI1mTw8/cagwsK7lgzFLpQhClD
eM0ixT74mbYhNUmDe41urWlj9FJqmVjYGN57RsuJ3wLkUa81ldSgRiijy2Kse4H9
kQCY6Qj0C3OZorMCLmcH1e7gsOx0gUrttwc0jv3Pr19/YDByAwfIpP3bzIdfVvIe
OMF/bFWUkuJJ0y3td4iCHXdQU5YCEmYfiDin2jEzu+3BC3dXKcbTGBi6Jw2oMkmP
2AlEiP2XY2y6TFyqYhr5kz2i2GZ8V23imAUdzT1wFe4eDEuVuHkhLYEWMa4kaU0X
xXj2hcbRMn9boTC08pbizbNIMdefxjyImiJRsK40GpaCn2gnO7YJVAIkauJLOK05
+jFBcR3nsnsDmdlIGGERR7Vudr0IlMt2AaszoquZbPQ8WNGMtmHj8X/YkTaNp6G5
hB+tN640Yi2nsHLppVP907brDhzQ+1gdO8jqlpiO4rz4vCIyeeEw70kFIPHz53qV
xhOixjC/T2JxYq4FCI6qL0zBuIgcwRM1qqiWgDSYR3jtcsWBwN92Enj3xsKnQcCi
pKMuJDwiguih8Suta1OoLBe9GegmWTKJj6hxUmeeY2ZibZb6DvpkU6dJdRv+rmvL
tgTWxtgYkV7BryPVqO0cLex0aUOHKgyAo/cKc70wu3/BFqgJi2c0Jt8O5ZRSoVqJ
2zbJO4OpmWamqA6dGu0QUEe6X70FDnu8/iSyC+aMLE9rmRarCy/XdWMdso7gjNBx
xWOsh+8WNYIa38MbFWiMEKmXcroOAv3oJeFrUk0OULKtz4HW1IGjhuXTcZr1QvZ/
b06Dy4Cs/ZfGXLM+ACBNPz0dHzRgwx65RTbGU5ymfYFW8DqGeAcJUaurzYF52c7u
riRggNmwcIlMzYjmFhZnCvSLf1RpEs6LB0HVWMQ1Un1sELOxVKXuQ3d4pn6EhryI
IS0ZkS70HylR3dldgZ4bnihEoq++ysuu380qkOvN7XfqNnpZ7FRB5GC8IUoKP2iI
NESwgKD0BAL/toRfOJajzhPjRyRBqLfljq+aVl9/jolBgSoo/Nmv5x0cFX6DYSR4
DZ5xiboxCXmDs4kW78/+8gdsAOXi53TwsSCm0Zf3IxbeEY8PdG3rhjOoPYVg9zJH
0pXWA26U/ewcuKki/KuJTOpcuzLCZJGJXMkHoQeLoybr25gxuIStIbKw/OZOTWUm
IUj1tAAnqcXE+5oh9m1VTElp7aOb3853+dAewCh61bm+tZEWoe6EVmh/zu8ez0Oe
ykjKgdIf9W4bkZaTZ1QVfXQzPqpLzVSl+0BzgkINBMu+WRnfUztvxAVbpNxqotpL
RJny2CZwDl6tiMdZZA5KCy/sWbrV3EjiMfjZYk2v9BlU3eftg4DgnAQdli5r4FqF
7iHsREAjTjmfXUY/tPR0+n5X9HGTKN828IwggqrQn9LizuNQHW3U+NBDnqn1+o6Q
XwWwB/rMxtY6ERaC7Mm/Bxq9cEwjIvLIBwhXXF4Vp2XND7MeMCpDpybqm8Y4uYZl
602Tqhl5saV10dhiU3OFOqtohx+YQfdgRSOaS4vl1QEevj4l8pqmej++v90el+1e
YbnW4U/pJ/mq/16BZ+vo9KZcUwnhKh3rtjNGYZoFSAeyabMcTj6J6X/b/Mo7+3zi
iGHNAm5RPlcQ1PpZo45O4zIE0EYKcnIXyYDjpY16kb3KzWcivmbzOJ5sA440oURq
Prf+8BACnNySZ6j4vcfroRVmD1xnaEmcfssJ3HJeTvU0FkAv14sufh2Jpjt+Y1+N
qnktfstek8S7yzOCdODCnDpxAN6lCeMDcxUuVm4esePY4oNn9qxP496XcJtkcTck
CAYNv+rf69/587kZ2uX0rqJ4xOxscRIKAtC95fDlgL7i7XG4kJ/M6+WfycNaHtyu
c3k2ZuC8CcSTRHKOJ8ZGwKGP6lIeg89yevMR+n/KkMAsuYqpetXdK35Ye85AHOb1
5IC67C1Q9DS8ZkDLbXB38EsvA7WwxDEbReS+HeuR7UQZ0RJmD5XvGIwtO79xcgtG
2yJeoQjAsgVfpJTdvAnKyTxqI3tspv26NGaj5HS8qZrjijoUAsGssl1imRqE4Mhr
IqLR4s8UGOfRoicIj23T9s1ga0lv74ppAyw/548NLY4t9AvRZhl7cHLEWQyn/SVC
MbFeMkyNcyAfkEXcpPspHY3H+k5MFJvNb4YecZDnf+ml3FLFQAbd+kA9hWmfwsuY
SEglDB1xexzpxAPP9IRUkasHFacT5EYQAabmbeVH1UAZEXkMeo/2VO4U+HfxDkm2
9ZrtcbFn/nd4DoEyM86kbNLd4rWx8dZjhUccBcYKLp4Nafj8W6WIbOx6yKtEewrh
6iTTQ8LpstEl/vMol2sUjIK9tllPlQFj47+LGcTDPS+uM3n0QqNk7bkNzHFPLVQR
EnOVDja39mivXnAtEBoYmmM/SLM9k8xgp1Ct5Cqv/IA/ymalmbgw2ytiUQadWwfF
cvTYZyoC5uQJf/VHLWkf2pYhqcTlEqh3dO6qlp/w1o0ekp1HOqUd4HOUmO/3x9qT
ORv9AqAZTa02EEmTX4GqCZS+zo0ixy2vWdxJzVaPB1Cl7+SsIApUCxL85VvcTdop
/EHYG5hg2zKRgHhKIYL7Hjcx4XErctF8NP73N27K1LImoPeNDCzUPYrgYozKc+UE
NcCntve47Aoc1BChAL0aniPTI7Ll9eHkHRJJfQddlxywlZZ1S7/UshhPgw+yDHHh
5LUylRwb6WPFRalErYBgqZVg1TrMTVqXcNZYqC0BxhM6embO8HlkAnYmydt4Gqv6
hxmgM7yDgIm422QYVEdi51uwjOQRCczDpPMQ/uzIgmlSI8l8X6aPYU2xxPlQq3oL
5jXXe+HM+do2iuWiMKZuyDVJXUG8R1otm1p6rVc7rbXmUFTRRMOam9SBkKnHF+3H
Cy03P0861TJ0jCZ/J5uyD9gRk3duiNy4Q0R0hlHUMakzmg79JtYu+FbNAQaBaJzf
7FBxZORaZe0B1IpygnHiu3/jR2kjWo42aad1dTZgt9Gdqn4a4E97AJ5ykI+nLbUC
KkUl7BSkFTY01sX8yC3/6dPPh8HziYhUraxqQLVJ8MJYCqlDACnHprxN/c2OzBZ/
PsXmrQwGlnzq4ZhkvdkUnW8Zu7AcrmvgWCuO+KpZfN86+/F3f+L2o/2hhQZJI+Ve
0ilgvLfWGxzIFB7A5HXYBOW4qHHtgsPcU1EnI07v3i+lAAKYSykNXflApqzmLesP
8ZK/wEXmf2a083b0MDVBCYUxt2w5oT0vpsYhiBtvi3ZrwC+NogJbnXhE1Cc7A7GD
g7V/Nnjiknr41MOQ2S8vrAvgoc6FABXW12BbJY1rR6kZNdDbWD6lZDsCobnWmkT/
i051JGQFlfhZhV5k1WRmHkFdZc86h3klJK8J6NjtBpo0P/ZnrwqkqnF2nvv+5kT6
JSm7eGuZeR9mu5uuKoR+8m4P3hG/T0pfR6C19dzTLP0BaIU+MhbiTecAomnPXXiL
Up9RUQpCcvp2WX9LDvSk6Tkf+IloyrSymUzSTrj2JfApGzD7VyDjzumLnJAzHBp9
pykZv7zb2kgbFRWULpi9w8O8kT8VFNLMf2V/U3KHRyqs4Z9zcS7Z2np3BMCOC9cG
YxrqS9btwe/pEjgodCCdLjQ3gAQaLBKvpiwrg2ht4ISpJtfAxw5aVl4oew2f7DAf
LWD48whooVukfQVQ8RBTT1eaNdKZemh+6WLZ2/R8bdcMwwH1U1uVaLCVpcVrlL8Y
Ftlifkc/G0SuwBQFS4mgqT9UPeLxIuWmmiey5+9dcRkLJtSZugpM9XfdJga7u3mS
2Jpu8IuY5lr6yDNbotni0dLuaaj83AYMxoRK74q1VWZSZkrtT440iR0Fm0BIBFIW
j/sEYd/u1YmwRx8HYRhmtyKDV7J9V4yPSSG9Csyu4HDmmdIyRSpGfMuwjAhEfyAq
bMvbGvC2NHqnlc0CHrS7c2tjApvruXnI+3TFTzWW5pM+2LarCFzsCnCVi1thyF3X
Ol8qlcawZFVzP0UArsflIY1hCjqSqsGT3JKVcENVWX4cOtZ2p1AtPdyV4v/U8sg+
fqOzvCmxl+mARxBSRgtNEOVLxdZec5lucpHqiMLs4hSh/pMlw29W3w8ozzGeeXMq
mIy0GVtDR3j25oww1+Lomn41o+JUlxSw7w0+s7nr3fBFVk5abunu09b0NSdkONMl
m00pFUUHTWbXTKTMeINy0dhDN/WSiQBSPev5Hyn2/Jv3JgHL1uKK8NxN1O18i4fB
6uDVqqFMQqmOKGm0yNxUe0+S1QsmWnCrMXqWCG5YnZ5xbhDw1xlHgAvZxbH+4lyj
eune0H+WWX+atycH4zUpjFksKUb2vNCHz+W84nkO/7HpENsomwDAPW10fZI6dcYj
xo5F7bhYZVVs2+LyWxMZDY6B+B9KiweRWuBLXKMKmBpDyXLJ2xCMLpvMrqBC40zJ
EZeni9b3kohVK7xdDDQXIi7g72PV4Vnc9uXb9LefM0qccLQgcEdJiIEmXvpEnhcy
d+fRrCq83Ia8PdqMscHPoNxNLe5E4F6RFganVwPPtI/28uYhVvfa6sGx1gbgofvO
rZwMGphHrmwfvFAZWggcChifH8ovBrBcTs01xmGB01i2pKXDJ/Fq0eyHA/E+py5P
hr9IeynLIRmF0glww/lrBflGcT1kZhxOBXR2QNQvRj50pldCbsJnkLe3wcahk0Mf
iXfcONcZREsuTBFeLRydA2a3DJ+LXDBpxS2nJ9vhmN52+4S7476qjMITHrJpsR3S
4cGuiEu0rKGMZsM2sLjDE5mPqzsfFHtbl6ztI/6kJAMjB/BGf7ge9svLC65CTber
Bvi0y/USdKCU40iXrh67+/PJOhjYAS43LvtytFLFuxZr3xIrbf/aJdCTh8x5PbT5
ZfptZajM2X3KsMKx6zDAaLHvzl6W0i/bcfF/nsvORrfLrIv3S5Ad8xIclVCua0Qt
WSaTLtZBJOFT2yKN+X6zoYAOppKp1Crk512y9zEk1y5yIpYxlY/FPF+mLf1AQJEp
8hXKDpEKmfvHZ4I9IvohcGsbx8OtSp7ecAmAFD5CteID6fv4JNqPHP68IqDfiwWU
F6/VC0Qs3jI/tetX2cEwQVIh+j0F+Bgrwtd/UWD4V2yYukta93l+sTCKau6n3e3+
cXirh0WHf7AGlMeGiIf2j0ji12nka0uX7th8e0FCBihA8kgy1wtjjQOCsRA+OSIw
8pRTJQSe0xXHfHLS3ft7I5/6a+Fhh2oWJAXfyHgUB4I/r3sHNNWBaKkqkfLENDez
Daqna1ynFhfyjk3WPfPGeNJYCRgRdMj+qWPHBtTB4fPc8oc1GomUJH7Pyjcpllk1
m6w1QjlmnQ7kKVqdxhHDyXPqP8rg0CTuP2A8mC9jYDn1zZivo8MfCuH19DvuWar3
EFtMV84bPyMe0KjGijkw6jl7CPeYAF3nQVAGzcWNGnOnZnALnNRO50BAT0cZgWaZ
rzK9mSvchzDmA7H48Vz3KaF7qR3AwhHq9Ju/1l3GArquUrYNn4og1xCZguPCwr38
k86FehBSvQ+axrKW/ZDaw9wersF8V3GPtZ5L/FvQU6Xzw/df43g+X3hw6l+wPUWX
KSvNE87T5+GIb/3zlvsKJ6EaTT7PR+MU/8nVX+hAGZAsj7G00JyBnUhBfGNdPbxP
5mHPTdgHHogzRDLsHJUwejSPOCJomcyKNZuNPHYrFFnHLcIiB1R/XNSB1z2+cmlJ
z9IHzDy3Mk4IeYSAoltE0r/SxMKPLeskepNH1CC9MGnI+PlGIyz38G4VTuS7ghTc
R0Q3W44oTcqiSqAcv0fiE1WtBhnffl3WPuxnrCf0C+jTgCOLoCazMJQxgO3gw6a1
JfRNelCtjMLxiY2k9nnb3iGN5qfY7F7jwonaopNhn2ix4f6zTRznwuwz2bK65gme
KSlBAh88JILC9c/E0cetV/yK2UtlZSqEFK18s0wp2mquosLAZj+gkYdpOCPImJrW
dKakLbASqQMt4xAYLniBf+rxHsYnEKImRWglMkL2Db8pkMPf53Uvtyf7Sfhqk06M
LLbGRHktgqVwn6uvKZREB7FgSVnAb/+DQAGza8n1pcbptCGpgsGk7AkVywdCwvnG
CppYOJgJWs8KJ8FRnhEF0xca0Sj/2+ScdFymD08Oy5zZUjDlVqlVI9oSUMUZpPl0
JisarH19ds/MVn/9xvmXbxnQRheRcgvbw27ophnVP/jaPQHaJKlrOVXYY/6Ijzam
O8sZ5DsfL9H9o4LB/YkdOKkxFGV/KqRZyU393HTs74eQDhq5lJU/pwYGO+634M8Z
kCFYCbhS+j8aMm8ngAGgiQBNaJ0xkN3jdQ4hON5xdtgyLA5b4EGTb90laWaTb/4Z
opBarKIQuOrADl31ZSkuoybwR9owRwZCvXebZCgi8FxiptYUXK/oZ3rEhnjh6wNv
RPfWpp6NHi14Pd+IZpGj8A3k1t1EYnOgLXvByWLSbj8wzy2ZLpDcSrTIDB7Z+a6E
cGUJdkwT1jbxvMTK3J/pWLI7sUfBi6Te6jYsXbSY04qmg84l9+6NcjEKDgUmiOCt
YwGkebUqbWyOm6JpZFhGgrh3txwLHxY/vk//9KZvd/Kkicd5iY87YDe1QyeF34U7
SRoDzVx0wyl42AK7D5kmaHfMQmDbGibyAdlxwZsDoqEDlJ8veYPJsy25TWk48oUv
Rbx2hc1eK81rZWRMuuw8MqpeFMGGS406YEr0NgxJV6xOjRJjDEmDZ4V/B5GXh0ft
pfvT1rAT5Z9K2ArUK8ih7KYeFDbgSSzL/1djVUEvzUclOXywvk/eHtE2THixgvKH
lqEtxKYQbgUmMHPAWelhC2qbPHZrtjgaJ1vLZiy02uFi73gvbrwN48yYsmN95CPt
LP6VRjdnEO8R34xuYroux2XFk07gl5vfjc5zqzpJC2K3kXfBoUvGdcUSYq7l1rXy
kYmsb3sVTuwQ8Nm/brCf11jX8y9ACr+IhLLj7NLKdqAyAYHmsZkWRqKG02nj46hT
fW8+ZHkXQXVLJVN6zmgTCA4KGotQOJACL1OKnYa+bow0ciQ1oxRAqBgvSKKsKd/E
ZJyeAQ+A0FmUpZ8GdZomQDMVrc34qcJMQse2CXYHdjhhrkvtbBSapmWgiKITYs4F
dactkYpFun1vB+UjgrJHQWcPVzWZr6OIt775LCg0cQGnfSFTO58ev2+lZgrlOd7V
j2pGwmQq2mK2ImoBRImVaQYpl2ptfg97ktFThgJpfjIupqvxDvLftW7A+Ev9YHaT
2GEzg4Ob1fkT++kKBjLtMuRdvGwoyH26M8wPV4nRstNe7HSPUeE87ytPqyz4IelQ
w9YYaDR3i+cwvBstvt6ZAJPB0UlybjHxXT3TYdNF8hA9Jxl3tU2SOvXKElf3Mgaz
au6adxGIyr6duC0kzM3KzRGP/sL5nlos4xJZ6vtwk/yhdbu1Xm0/1M8dX7rHNRnm
dzYat0zKSCmpA6FTs+3/qd2tt6PUopvFzWZqtVpgOTdmPNtFGozu0vS0KQsYGjJZ
GA2mowyX89r2A1/VXb5KEfKSu16lEILYiGwD2DXYh80khgjvrTWLkrrR+IxTKrVy
FrHN7+QKBQ9g3JPwltWRLUvY0gUilmHvYMRYQUIJaEkIzionZhgHKUTbHjsqF+kA
axvTmovTh48ikPnMVMA/QHK9B9iviFdpn4CFxrQlCK25R2/Kmz3WUrZd1nhG3Fk0
GuZpJrWeX9jkk9VG0BwrJH9Ny2dN86EvLlF94pBwO8IeW1QhVoxJKYXJo2H3BqmL
+JrImeOFiUjzM6+7Yvk7GQiu1g1obPhPvXViJdqoC+16cVEKeqwRX+9ASvCO2GCq
HKR/amDZc0Zm2bnD5ComNmeyaSvojYiiyMuAdEaNjdUa7gKoDJWkZxyJb9TrTcD5
L2utRiS91iBP6dV3pe3TW+kPbLTRdaiCXiaMdTC3qG5yEzjKrarc52pEBau+JBXT
57z9UfRYXM8BuAj6QyJ+9MDl4GGYVVqxFLpF3D3UWjLWF34FVDekug3ilfNWsulp
92wlMS+Ki/rCAJRw8VAqWXQixNPM1vhfsLWAso8EcojWO/ApPuTYymvO52u8dSUa
Ji8ODpoZM3mN8Tmfp0TMFDl1HYxPTXTuIkALxXn4NADFiBUfhaPBWKnaya1LPLz/
NkFa3BcTZhHCKNAlJXV99su6ISA7Hhk5zT0f5YwVEQumcvNZ3hJO1QLziSA+089w
9e83sG1ynO6/KOsW8zs41iuLd8nDHo1uHzPBuC1FvqaLo8OCflPHUXOd1qzA4CaF
RIkIYsilBax24RsZsSl7msZD4+QV+vqsimI6/EkCWhjMwXOWjOVH/LbPqrXms8FG
r27P0KPSwam80/8VvNx4Jzeww9opoK4WjnRmf+qPRwNGcHXBzPEZxe6V2lSBLJ4W
2w2rqdPNl1KpOO37UQjbkSEtVPu+x+CljEi9/bskyf3Ume8DrGWtLetsM95whIn/
HxscFM1L2dvtgWoFUbqjQC6cLp66kM7pKxiuFTZ/KahJ5taUfBSO5+9a+wKdOgNp
esssBB9SQSVCuT713X6W1Lj4jQCTLHNpQopnOcsDe5v7mbRv6AzkTFMeIyn751HF
LjNRoIvf04Cob7EGXDEt5BVVefjJXERwoDqLljUth0wFARHl+Mt2fllHg34kNCKV
NQh+Rv0ADdDi4tLnczuucGiYFm75OPHRBTyhoElduXM2iXkKdrDogjaMF/31MQDp
pA7TunIDoyjDHWF1E3mAD4fAYxFkQ0BfzZjL4eumCPTHrG0DKLLDe9/G0pE7dFMQ
wnx2JZsJtQVJLVhS4IwkyTOrdNy8jwClRqu86eI13BZyRBHFqfF6VTvLzmoI/sjW
df2xHj2MZx5gFbBC4+aRRqyA9ykewB3LCTN2aKrEZiyO0/KLeWK5XH8z60TYrBMj
wG4K326Jqm6xsGctcwm+PtN1Nd0m/jZED2puLM+SPHy4VGBXl/hv8uRCPm8JI7n8
ReHl981TUkaKkBI6v20NWNKneBzExNTQJ6ZdmOrgsZtVieKYbNiDuHwEV+hdsvqT
gpZEuPCo1myqByLncOiywMbaQNojKWTPWyL29DBhOITRv5BQjR+zBqK1XzbrYCGR
ipcRyZiziy59oSoZlVJR/DPjLny7ZT+wCO7PY7tkj/APmlYzMT5nFRXSekjZZQql
x9MFQ22eQDnKKf5nNVvBj1o4kSv6oOKNACj8cyfW1b/Lq+PcmHkNMdCf60rYrKB6
IMaUE0o/AndzWQs6NQb5cnyOjp0jwIi0COkGww0PVRrXXX4RE0RkScO1kZqCU1rA
9OZYYJC+9B7qXeBbuAB/bczDH1LFg11QfWR6MmyvdT07e2wwtbDtg+BEh6R2pAl9
RllRafou+EDBD3qZ7z8cmW0kVzNckUgEEGdJtgQ20hZ4LLScd8mzIxZO0LzuPUZI
BDoh4SxfJoTcbcRvaAkEdIqspwK19nI0GcDdBH/0m1+j/FiWfTYuG32axLmnWYyb
VGz+1vFq0QMltb5pcQTCqPIJOFEcRa7XbjF3smPZi3za4CFNR0k0WDaZSJJTpSjX
314EXgCqalp2OCmBqvcO4jW3ioQvsryRb2N9rWhQCEMGakaB6Ocfh9Yqn0s8Mbmg
ANh8Hnpz7MUyEcuqx8dOY/SDqtyo9lYpG2bRXGORpyXMIbj9fQnqsyqv1DoN5Qz6
xtlzze0BT6yd3xVAGTMhBj2uL8357Po9FQaF75TnzIS+EhceOjDIAU8KCYhaKmzk
Queo2ZECVYLjiSKRnS3gpnlt1Bbpuzout/dd0bQYwtQ53w9HoIk9Ocb7QBSRAo3W
RwFQJXGAlYb3Fo3By2GjhgGHi4y3sklOzqzfS8+3eOj0zJ3FD7jlrwLY9yC2Pp6e
TXCwqj17//tk49BJKCU/Nm/sjnhJKlTFWGRpzM5NZzRs5GScpRQhRbxiSizO4EPd
0PnJWHAzPp56+SDnhtHn3zd7maSXt0Ueb4ALRXpdb8nnSUpn4aMJcSL903kgvqM6
oF74SaP8xDSlfgI9yHoDMSDaqAeAP3Zbs0uQ3JPvonh8ltLdq2wN/cp4eNfV7grC
0rHn1jtSogYMkUBMZ26ggZkZeeXg6bqNCvBNxTEMscGlvaQ5JszU+qe/ZdX3WIN+
C5qrBzqunRjr6YLNtmFL97+tRZq6JL80443h831YUdO5ZO2otJ+fZ20eD9ENndZ/
HITshAwBW5Hc75JFzJPW06EOjXbfzTLzRxsKwaxY9sV40t93OGCQY7qJu3DrqH2f
YaGrNhjkyRTtdp/2KTc43nkEBa9Yz4rRfSu6fXLicKg/zb9KylJNcKnru32RBfmy
nk4FVEy8H5NUV60KU1iDPnxZzo+T8Q/VKL+QK1KcRLaryZvqiwciGmpAtFjlngtG
KSZXIS0GwmiVwlvy1kNxROITMB7gFk49Ms+6vI2YnZrW2n8l5X/ZhuK+KinpgDKD
ApmId/BRCxeLPahzAeq5AwLyls0J/ef5z/uw2w09eQYQm7bbM6UvCL4csNf24waB
g7wAjx/V/Gd4l9IVynmdaf/DOe5bguOemUhDz4QqoQkbB0iiQO2Ktuickw7++euX
erVBFXN3ONvkfNHkYpoQtODnfeW9DXxvlPDWuyhTpWoX2rEe1ACu5YeiHRdLxCVK
uiBK+ij8uZOlYXi8iNLdobZP99QCfLTzaGFfCD2VgM8/Arr3tve6J1ap0bk+P8U7
Qblw1zIoG3K6uvO7F7MY7jH8VPNSCO00WFbvV/H3AmHQDniqi2MIV6oX4XWnKp5T
Q/lHkfn4+YAqXk2QaFrmHyKYAIoTmX8R0Y2SB2jzCc69GtT51is+lOgWc7paETZr
/33A5j1e9Y03GM2Uevbgxp+sznTKQuV/ypBFywQfX/vlttL8agBU9CVpZN/yfoid
DgqV6LhOfhxr8+mNi0KaYUJbi5TStzXzB64wfIo1D9pGeoWTRRkd52iFSqTjyupm
WRv6UErYdWlTzmdzNSvlRr1FQmsEW9pAaN7vkw4cWSVrMHTr2BVQ6MXq4Ymhs2sb
sq6G4OhX5aKEbK4uwJ8bmqBcgT5Q+54VEV2xKsfS0BlBqnKms/k8LyRZOzKWnQcu
VoZExuIeuuFdnTR6kXfYIHtg1aCAolpxiPQrp931wLLyj2a1i8Rxd8sJT1s7Tspt
1eUkMwlwFtrAFGBXg9QiiX3rVrZYgjkb5kjbcHJW3V3R8ISlwzyG5MO1P57aDWuf
JV9jF1Hy3DTMEn1Vk9JjykH3g/5Pm/x0MWm+ERdVMo5RUjPUXxb0VRsY68NiWB5v
WNZzRuJIWCosmOJ9Go1sh5qThPLJpuXntFryL4MLAyb9DXqi0jCiOxdLdP0eYQLW
TPxSZBFiGHzR0xQC/BPjwtA85v9chSPLGuktpglyAQW7Z//8QRMuIszh7y7SwENh
qVlxABlvBIgMehYt+p1DUaAwm/gGviHtli3MmU89pYDTFyjp6Ri1ukEC45l+OqLf
sfG7igKRL+JsVRlGh5PtDiLUOAueIls1fQM3yxla6y5+yEF94P2oEWfwfW0FsV5J
eUlr1q561e70MWxQaip1NG+/adwsg9FCySivPNCPfYjF/sEIMxw5KdBNWlC80O31
Xc4k9C1Zm9uapndX7obOPMtJhbiI5hES7wiFAloNVjnSLxeQUCEZ07wxwoPybvIq
8Qfxl2/XQPHNg4CwSxSuHcimGwhcGD4kucwwodLF2x/AIuYAuDLy3zSHk6Kk+yqf
t4+ZP9YN0cEGN9edM/xcgXu6VUpACUpDvCxwtf6w1nF5Ms33HKH93SWm4SsmJnBZ
jpQGA128P9/5gsfIEoolm9eRJSJGMatMOHhUEtlz20615kINs3KFRDrsoTJpsg24
JhPAeD3X7OsrVV81ZPvMiamS6bLl3laWu88xUcSDVINawQUrlIQoA3un0GOJ+AiJ
el+/yjLnDSTXD+Jni2WbqZQ+T4KSvgnHEsrYOuYJ6e0uDrXGMyLUcMQYNNKPFsjf
3rgoYZT/FamWsIUhaHTYlHmIPS+803vj87a4DZYUi/RZeR2RBm1lXWFkUY36mGQf
J9SWexSh1cpEYR2fbgCM5VCNnVhBO0CoZ1BfYz/W2w/z21bIjUTZE6JzKbBXV+Jy
AS6sQKkccAGLXilPQm8GMsSehR6F0C0IYyfmzahIsBnbvHsdLT/TKYdfyumvNgsE
MKM32avhh7e7XualL7fi1+C6/oLjruKuyTHhA+TahbDH7tFD59jEFH9CvMSrDPDM
em/LnlYQ1k/ZcHqwtWoF4BuF3rmbfr3zCJMcala+AQn/+Vv5UoKNwRdARzttAeMi
EUlWGRQiDq8S0RUlOsbTJYU1zcn4ADtCPL5Y0PjQEJRgDfECZM4KGY3jhMBX1cyB
f16T5UMGFotHiwQwG7PNQxeCev9018mW7O7gHknvKp+smVHMmbdBhPh4n0zD4ARD
I6FornPbYMoAoHQllVHsor/lv3nTHJfCnLmwy2l82f5hY5J8zsGKl27VS/uq/+tT
FbsrU0+xJzLx4p5EnjpvlA8g58sd0bl3DoVSHTL9thvPjiflV+EkUl9FJvxqJ99P
HxLb9Lx9PLcD7a4tZb/Tr+Op0NtgLqRBy/0eC0A1kfr5lA0rlGKUl9Yd3xMOJG5J
Pd9RMJT9miPUqknESKQyS3Svzhnw7AojZ7rP5zRWqtgoNip4WzUoY3wEhBIuyF3u
bU/JKg+xjxJhkRNWArUMWkBpf1XtMKhvsfdu+D9qd54BpNaN+AnuzljlvjmRjTWk
9e9iey7Z1neCV/9iUaxp0djKAY7kH4kuj0HIQ7V5DNVetsNAo0jXQ+tnbZXv9vo4
6uWeYn9uUMzV+k1VqyNA1FT75CDf1fJD6Z49fyxGG3+0zkA02xORhWUjYHX3TRIS
DE26qHY67aTVLwYyX/7HJorZH2Y8XQFbDL7l0fwe1tUYjt188gO91O8eds55xFdW
Ul9TgpKMc1eRU4BNpUNg4cPGkT5CSGXqz3NkGVjXrn/Mn+r0mvH6eMEC4KzgWL9i
V+SqmtqtCdVMi4SJbOtT9/r8nedv/2kln2WL7nbNikcr7+y9+jN0jyT+TT6RcZMP
hXm5VdZ3Vk7TEoi1aA3Ms3rdy90jSvyWqi1xpBtU5NvcATDZ+6VPRpa41Al+LnZ9
ijuMrFpuQKKb8O5xx5w2esKGv6siZTtkSVqwjVCmZ8Gv4Ns1h4zlD1pinvbsmghZ
FyR44DPpJoKisJKe2LOzoN2irNO2bwBLCS6C5RNUbfRJ02Uz+CygLsYnDHZeCmcQ
axT7YKFD87780/MOFI9agiKfT3vHY23MxdHYgb/oXOALAxXMY6jNTG2LrOlz/AMi
QGhFzzjS9QWWGoXFeLUtDVy+r7sjhaqNJMVy5zvZTl1+M4/e5ASc/5DvQ8yuROJJ
bGkd0cVg3vFUSQy3akNO0rW/dinq/xTJfIBqkfCgwopkGDSUbzZdxbEG7zgrG8E+
/MiCBsvJ84WplmwTLibFI7ojHZlFP6ZoW7XOpaWpbnfqTLqVelEw68eMZzaxXCPl
DHfPcOjOf0rBLT8JHQ7/1+yTzBvT7pyZ3gBv23hG4/rTncliLlMzjClMC1gvQ2hZ
9liFyWhsi/bkA3QCaTRSfCRPMfidUHtIbymYuUKOOGdjGbuK/rAAxgrydP6h7X+Z
sCwHG880gsRKSABtUrS2yHDWp5zaFtSZuLRzyxwgE76AKSZ3sKQlEBrUulftIemH
L69fGKsJt1HM8fa7G5D3nQDSMj20liYh1aiyG0L8hRsc9I7hXlMQ2Npki8ptoo/0
RkAO7mZ16SxGiTBnn02/lfxP7aSgR82ESLolFWw4E6E4LZ1cvMhUJNP2XdCC1x1H
NTCX8LA0hE6huIwGD2csfkpiXLYg7Tx+jXSoZuANtlPH+2m3bXlypqQCLEfM8a1Z
K0JlpCGCqkxOCLjpEVJY8lEzXGCfPW3Own0ztAU3DR2wNQNqfkFUOTt3kmcC/OPK
LBx/AR30jU+N9K/D8+fDKkmAAH9reTWrer+VMfbS5kC32vqMYnSU4Du66gHArGiM
voQBfMWp8o2i90hJMGBwacWywSi+789x4PaaZnc9BA7d2qzPgXq+xrJEfmEDTBmF
QrZJWmzqyND8T0JtPALc+DF5HwCiqlmv9CabvhZXhgpbbHLKAFQzWXp5eb9gAWM9
gFjP0xrn5A5x0+dpbl3ggFNfDHDM2xkXFX+X221fhXSCmYgGOVRiavWBhANIk6bg
A14q6i4rgrPc2isVgSNXZvJtn1bQ4oV9PcI/mMfj7bGtUob6hJ4hQnfocFfu9nT1
EbX1nsuytaczxtcJRXFcFIx9BCn/U7NrswzOyhTI8EiQfgQB1Wq+WKXzhztqjhjg
U7n0iWHrS+Zb2DALy0NQbeNeL9NE01gq6LdGtVRdXEfgfD1H/OYzzewq0m0BWPbx
O2LZm8PRmoMOzAwNCOimcfzdwaAPkOX79X6oIXbmIoseJzf8TCO44eqoMVBodzjI
1YdT6TJC7aHAI9XY6ys3J3hcvATmyCMLtWWZFjRWj8mWM0JcG3KmTgK6o5AaW6UX
MYkKuRX70usfwU51Ml5n/VkvOKEwhoVnwBxDuS7BuE/mNN/k2t9pHwWfBdOUgN5v
XasUFUIzW0YY0Z4HA/RLYvrQIXRdv1oVlEe3Pdx1X/cwtA9w6nAyzKwSblDe0J1g
4BJ1968Qnu3h5jldlPbpg/8eWOlaDrE/jEdELq1wfNVPaXGng6Ez6vpGPo9z/KdL
4t8L7PhgEdIVNcePdQwiXK6kynEBB0aoAJCBOagUA7Cs19XdG03vjHMiHQ9cDJ+h
jr/dNHaN6O91ZfTdIT1ZAmOQHQfrPaMqTn7w0yPniPJspVS/oANFGlwxEZYLL+hT
GLJlFvrKEXDvLaLgBnB0m9yW/UwAkcEQopsl9JSTJcyz39+mz2yMNrk7UTxN474s
/wauYGMS9+qTEF45gB5CXvEfeUxnABHZfFXODyKCo8na9WPuP6EqERxlMtBl5Rjy
9iokorXcJqJgy1xNjpIPTmBl3d7ntq61By+qn3SHUO5r0SS1RHnr0SFXMK4TDMa7
mliaSieb1vo+Iu+zqjLYVq+iQEgY8yOvEDyBiX/OMwRQGHM+uFAfkALJIaRE/z5c
J69c1iGHIs9xGd4jJFTYQx/WnCYXZuRmQQdH18VaQVySXJbyMZf0zJQU4IIhezk1
Qb+mUHlZk7qBXTVczQlz4LiORTFbuvYC7+IUnypCq8SWbcsJio+YtdlkZOee7ajJ
Xd25T+uyapi4rZX+ZncUWBU/0r5hwGnm8mGzncZW83HNREQCva2BWoplLrxlnt5G
+TQ06gpwDcctT3nGGIfiW+nByFkQCOSdoI09/+DPah5HV/dW3OtxXpSnDkLT/fvc
132UIlB1/MpWbNGwl4wjWNyzKXPepmL3wvChI35ftkBBAhIZg4Lye/jSOUCIhP7D
yfong1HGTqit6J2zg42hA6XUS71qjkN2Mpl0++joby6icPiWjOXlTD9inH9hgWeT
s4r4vfrNhxpmVKl+DlgGmSP21I9XLsT3/Gi722WKRnf/XSxs/1ZvMZx8wyifhvH+
fIdu5aP/v5ObxtdetubC1mj4vIara0uuvrdHs2YaI/gpMYAFGq1zMCvZXXmH2gqX
pNHPA2cia8qEwA/eHxPUx+I0qTAD2DrQJh6yB80vyWEMxZagp/zw2LT3f9++QXNr
JtCCFkH/iYtiyr+kLb6e8R8Xn3PuPK6U192tDyQ2BD5KSyNXtqovkGG6sG+vcc3r
5T3IL4S+8VMiiq2DXW2X190bKl2O1Tfw5MgCRhVDURELDRVRfKVpyopAfZvpstzo
6v/sMYswjUxsA0p3ujhhV+6JXKH2224bK48E5821GNc4pwFeoN1KcRGtoHua4gDB
/08inr/Ra0EkX92C+GQEL39X3jfVVvkdQ6TteZbrVgSCHZ3mUjepeT9li5n+2FVT
mSKWjGG+DMIH9fgYqD9pR7XxzkwieOGQ29T/XSmXaXv86c6NCy8ThWaFbALhSi2J
XKXDiIPkxaefbxxzTMs9AGSSgbe1fNHEkttqMmJUPBoKY2I8FOK5Jynle1mygipA
ZymK+wjdBCJVDTkXW7Y8su3aGmYLkq4AV/gup2EexxGYU43vO510BwIGs9Rsnojz
2PbwPDghlaWqE4Gw4EHZI+GRN+DU4xI+oWpFag5gDh48Z5ulWsB97vKD7z0F9BhN
ywSItHUN/oK18QnaWPvWVWgdg6rdC4DPIjARrpkcnqIkBsbWYYAQTUafks353XiI
x3z75u2dSOC9dL+XYT2qM+mRLDhgBx5D6vSL4HTRpPv4Cl1hfJ4MbxWQL5sxE88+
/dsXoJqtfdeIQvE/G+zjXnzzfv7CUIYf8SNsUsVbVCu+k69qHurXpt3MYiUTyKvi
uLLgH57m+6MVX9xSFH8HqHLdTAc3HU/GBkmTIL0LZmitRUpEEs6NDLH+H5GlnqiW
yxjH9fJHts2lyoaHRo7jCdoJeUe3aJVZoeFDIBL2GsEJ4GFZ7Y8nEYQYB81ipK7m
tWoir3vJ5ZN4Eaj3wyVftgUVyHdRenpxnARZVblIw+yx2e6gBwY4kago9yEq1t6c
iNHOgjyKruJXoqV+KrnRTZ1CwitbwBKtCBWkx9DK4yL6kU4eIwIYSQ/YOCHIhq5r
AvpTcSyxZ3tVti94KnPpYds99OLTsfC82+RUXOr9tIYAJLJAlydLR8zmCJiVTTCr
P867U23g9UMLRALpRA9YdohUQ1KAeSEMy+rim+nShvbY9fDwZHqkI3Ittsy99bSs
ydzSny4pl+cVFcr88ipOv0vPBVb/cF8VMt4GymqN8CWM0Yk6pKX2bcAcYy8irpbY
m1Uv9SDvsQnv8oRK6Z2NV6tdQLFSD6qMW/0J/nfBwfSOacveOENp9CyMpw4NDoUQ
EKgxAWX9AAWRujJQh0DtSUwNHbZcN+RbHnyhdicTB/HaWZjSivThngCJE6T22Qzq
gQ1HWwpFiEGf31iYH7EiIDzKerRwoKCQnrcDH8L36eN+jU020/NRPe7NwWq61hCF
wcHpuPC3R62AjMRBB66vRki0Sc8si7awguGeiXYw1Ou8FYvGAmclQpSnvRVY1gtH
4NQpXMg0bOqVUEliZ/nSDwUEkZOhrsYbCPGBpGAjvSVVONaAf8rkJqPrmPRtVsXB
U+wJ2KBZDo/r9hnoKUGIafogaij1QkwyRKY7ytT+PK5FuvMxtRQFvgFdo4uvUbB3
OUXb/OKbZjyit9Z/LsS8UN0/ePhifg7C0qsO/7kzqcx+YwOx5ePkqdX7B3/3qsbs
qVbj3arV9aV47HHNYUzSKHGlZAeYi8kzJ8qZC3MYgsII2L9QDHMAKMexOyK2Myq5
Nv8fRU8GJmy3CjhzENmGO8MisqSYIcrP90J/J0MX/x6Kh9SBmPx68yXdD2aPUsNy
WYUxXYcWPpCgv3Jj/4CyrGNsj19u8VfFvzvADqC5gLcL2qXM6jNa4ZJBH+yvvmEg
641KNI+w9kJFHX0fMbtPMOYJmrUuMgup0uI9x0LyUlBzeS9YDOrbENjXNGwtcDtN
8T+Qx3hKl52KwG3eDMt4/e4OE0YU352IY+XSUNxgKBUpEeLSulGjZwZopkW5U8cG
3bnMTS3UGKUtoArvwf+dzEAIVdpbCqQJJGSTKIOVUL2Ux/wryAT1t2u5SLmAA+kv
XHgCMHBaE+oeDdjNUGs8iIYYaML99gysa6ddwmAqPCRVOcHS8Tiw1OL1+cxNBGfu
d5Pw4JFDCufELp+t6IaIU+ZxYKzrcPCNZQypG8rM3FccSI9TPG8js3pS3vXmjpOB
A3GXF5Da2IgVsiD/Xkwz/CuvjWqrszTW83NBcsmuPD/tmIfJL4TlYVtR9uvd5B5q
QoWnBC1s/gpQ+SlTCPj2iJ3F/9jAFwyFUKoFOhU65wSgZREMjFdlkQwbyfTPgOVF
1XgCcH2g0vhKYXtnJR4+ZvWpL2iLtCYOROGhcXoZFoCOhHI4P13z9+mlFOtXtORm
/9lVHmLEbOa0qIll/v5KrcX6DY7OhMm7qIZSvon53u6oYr12enkdunItz3DT4NqQ
b2m0MhM8hfQOLRkHfZ0130GTXmklJpM4Nn20qrbcpBnzEtqk1xehoMwXPeUUaB2I
IUu3ivMF19Yr9K+RBSd82s4OOO8iWQR/SJd1I19BMT798thkCPsWYRrutDHAIu7L
JqidcDYWe4qmTWTdmucTTc1c68XF9GOpobkCcVfjNoUtM2Pk+k4nkc5EikenPVLh
Gs92pjlJ0BSx+LJ23vNwHuk8FCIG2M8aHNm6UltjwR7LVqfPB5XzCb8kibqKCsp7
4WvbnsSIUVSh9JDk5JKO/yeBpGETPq5nEn099jZPivovVa+NaKycl8mwTxnjx9hD
81TELXOKP9xUXrYnqSMN6lIIn9WF7Q9KD+U4J9OYFleAer2HLgARs1tfiIfWB4Ua
nWgR51GgMHh+nqANKChUytr4oswANJPY6FMF7uCCVgd4VYZv/TA3T69inyf2WmEd
Jz12DMVm/CC3zmB3RnO3Cqglpx2xDzfDbIC4CwqJYib31EV8ktQXDIsjiqwwPvX+
Mq2vIRIYFrSHx1Db7mbylnZhFQOB47kqdbPQlEq7ZQqU+24WXauVCMPd1rgaMG2F
dSSxCQa8zKBSO2fmPxR/cjFlgTcbPEMHiUN8mYio/ozvZngF2lREONGve/Yysd1O
R246ugEoXKh5JW0ZD+5EFX+xU3WtyJjSuCavQwkl+rbnkR5VBvTdYqhoengD2+Pe
Wx6PlU6puDYhF+/ZJ5TlLFHc9/oYldN79ogbrQHtHE1zKWhJw3rKrCtuXtuJJExa
FgsjLximEmcIdrqogpd2SLpJaoZs5rksDe126Q/UmVV27xVVwmLwu+NpggcT543z
9hDsZ5qtVbqGfNnVxSEuRoBzQMzOsTkXYiiIBH2xVKHJVXgch65Pub4n4KwrPG05
dFYMYgtE4e8SHnHjjbr/cDEuGYCx5qXuoVXNE1K95YFkZgLRfU5Oc0Y4I5MuyMJH
iouhQ3W364/pwXMJuw2oFVeTK5U88ZMZumfL8beUJvgwF0ffoxoGdaGpZZNMIdQH
gvHSxYFUfzEK4bvlAF36ng6coJ/cUVTICeqeGRjQ6KsW3nnuqxIPDYAsLBbljOYq
2rOeHLmFrJFDYggdiPD/dWvWXh/RUtSeb8dNv7MTjLKfVolrcTTTK81ARfKdaUDl
fJm9MDHubcfLKb0UpTFoQYyQVQauKcSNJm8FBx9tevSnGqcxeBbkFXlmkZ3px8mN
rRXIJ+2n4/Zs+cVfFG4v7uTbHIGNKznVr/TVtLWRBFBzb7eQV3dqZUKHUDq7z7rI
Mfg2ghEvBXMbS+hILjDZndupTPwgoDwCc7Vadzxf1QGlDL92TqtS2jlRnfuL7dxj
kgkjjuu43YzohNrEobzxPiJDa7ilMtEnYjQLI5H0yGrhL7+nTf8GR3GKXnYO130r
qSdnYHWl9p39T5pzTSwKAE5ikHf0hTrjVWOlaP8nNIuRAbh01ucTDcPDj04VIUAU
dCwa5yeoq7Hluv3A4T/eB1oarEZ9tqr3DZO2vzF8SMlapt8knTPIKwhOfA0hVq84
7tHWJ0wclf+j6xxq90zFy2wWGPlZartfkARO4Clb3iak1b5sq/XTrvkBT2pUagBT
RbNkPP/glLF4QnTxxPIyNIUdQt2ToK6GGdO2TiQZfrrzVlia/0ECJ/4wD+EgNEc3
qVzYcun+YgUl7GUDd0tMwpFB3rylkVsxe1aSBzAkxOAPdJKZ0bbVSEcM1ZvGTMM2
ZRjxZrCch6Umu2BdiGZ38ApbMblxA/CgH0NyxtWnDTRgQJh3Wf18riFVBvqp8ysN
JeTSet+zGZMvRi5LDCjywXGvkvSdKPL5ijjWozeEoOMpXYBHPDT48CLvQk5+QbVP
/WX6p6buNCXsM2hDI7VhJ8aRqKZS16XNoGoFdWJt4YDBcXSIzObvTaNZb8PtD+NR
F1Hy99QTlLFRP7rBBCJa6nBVXGZxPLh7LJgE14Qj1fdbGVS7AOfvXxyaQjhydboy
mOtNtwUhIvsEHh8jxEdvejBuK4hi5R4/rbSyFBxjaO7GNPSbhjGPe+wV4wna76Go
+c2Ukx7KY5Dyq4IAv25duFVdr5ff6lnveDlM5cwUPfefmg0Ev63JF3WdqR130N0v
hyFy3RoRO5dgYJ6lTZTqhixzE8CFOe6ZvuFXAceVGGO7GDV+OrIMYuNO6ouiRvVo
1HQ2KOHjSxYs30t70uwAXPs06vrboPUrtcy7/UJuHqLIDD/5OSyazVI4rP5lLtBV
KYUBdvQlPV3kaFFjTA9Q6noAJsEqOXXetul8nvHdcg5DJZ9vKUaA3ldyTCeSgeQJ
SQD/HCODCUI5LwqHUJzGib33HW9Sc2OpjhDD7j3pgrih91hGSD4EnewxtUqB0Eu7
PBwFq7PNh0cYQP8/x4ddtKk0TBsy6qK0AanDxdWdk2xYX9FKHmprUSXZi2Q3zECm
n6zEU8ddqBAMMOuGQkNwF/TZdA98yOeOuTBbaCmMTp5tJRLWMzDg0FeNPKIH6yg8
FiRO6KKSXxTDfmH3PenoWpMr5tJhuS/IrDWsQCk0sPKqaUbSL0+BzEgAJVILoCoW
wD1+6u4eQS4XszTmGQjYmU/rHjrPQcm8Trd2G7iXKKWfP47/hQVkwOK1NiwOi+Ml
wuIRNlISubSbWjRzmz0/NZ+tRNeV2zRwp1XzRUM6EOqxQJRGYGCT7/3ThumdsPJN
McGXDpO1wnavEVmUY3pZJ+ub6/AktQaXdSSLdF+KaPgQhu1cjkipOoOjxRPe+zv0
gauLuCvc3rDOoGN5tnhagjCiIaWhkYyF9wO229lPC9zFhD0mlBJJOB9+Ev5EpkgC
049Z4ZFekJi5lL5Y+urkVmta70RqTnUdAUHUhH9xiMZo/Ha2GcYYX352HJeJLzu6
oz4UHaQjhdkrh/aHc0YI1r1mVabnJFIY+O0LY1BEHzM9B6Mh1XnL4efJJsH0Ldeq
xnZxgU0NvUSkoIucxWLRjHPI5uJRVv/apvremt9gA4beoBpabEk3ixhADoWR6/Vs
g1HuQy1jrw8olQR2uheb/zevisQAb6rUxi7kSRDBgoYcAo3X2RwTClLgvAPJivvD
h/SjSfs52ygk0c5cBx2wfQOS+MxeTtJBgRGR6g7lPXRUhbwz4VuXThX7auTyWlhh
YHXyqAar83EQsFtv3wpbyMuM0nB0+5FhT6fZ4M5ni5Kl5jMDLyq34KXeak1CDrL9
iSooBcZnYReTcrZXKBI80/SLDnOTIXNHvDmy5yzR8i/5TnHOKDjzLTrRVKckvnkE
m9LPeR5A+h06NfGMPdVZOHSc8Qlo4bpx1zcizab6yeEq78EQu5rEe0GVTeInbmo4
8SXRtnvYoRDsSaQVtx/lm2NItLmb0Rr7TE8rwh5Qd99+Dp+wYXk3jCVtZANfpvo/
eC717xxcOFbOTvigpdDM8iiqv3Cz80+BRZSOcmHlM7xWMZH7f0l7nX3qxljbvroG
+s+7NOYCglmtOxgdMu1eYB6QJuK9rJtQm9pPdyLd/dlcjmrS6ZEUzy4r320bCcDL
F0SPIjnYIPi3CYHnRERJok1BurQ1aQICmsVkF2Dk4p2WxL0EGOt9NElEK8N6FiPp
gSkg1lEEryNa/SFURYuEwmtncKt/zyiYBF8t5Bei7t0ObrwkZxPYmVnooOHGcBbD
4dMEShKsMMFtcRKzOJA/7rbCcHagwQyEHEsvX6OyIugswwGl9YSJTKTNhJjB3JIc
ZYOk0HNN6gfErgqXlZitNrvhenhaRB6bBZizAe1g1sp3vgyEomgxrxy/nPb2/8TX
AE8Bw4tK+cgz9bGS88P7nOv58uW1jd+MsujBY13aO1dcvYtppXasxaRmVhXG1Z6U
jWbu68PMCHGVV0j5WtPTFVSzmwYHaoEtqhwqDZkotbUzFlqw07meZnWYeF40gIFR
u9Fw5B6NmbNviBzh5h+9inb//AZ6MMUBe/5PNRLaPsSHP5xW5zam9xtfFZlCy5Wt
21lXazphRi2fu9KgGyx2bz4bEhx484U7QSBYQw/tiX7qW1gcdDaAimBXX/Ri2SvB
OakIbkWzofN36woOljmLXVCJ6nQOdbl/nnJYJPufKbOkU8fA8Xp17IRoJaKzkHXU
uWYlsFL/OhvpyAUFbVqfIT57brxm7Omj05QnWzmSQy9d6zf5/hBvLXVQ0JQ/FDse
Cu0FZWwoaxVx9yqRMYGteQx5F6VDtMR+JOSrLJV4C+cF1kfiiXxbvliL5oswO7dR
em3xkvnJSLatNOrGdEA4rmwTb8Ur1EKGhq3+WxFeHmO/NMK2FHl4hs7ncD5Fb3EE
epa3oQe3DbcQXmMo1R9dIOoV+8vlrvcbOTUTPUy1jS7isZNVUOfGGgGgPxxW+U5c
jRcqT7Ijfz7tSL8TAt3ORNjbX/5RaB+zFtVAIVUgL+npzi8NXpXkYl74s3eF4qDc
LNsDr87KCZ/VdFo5gym+rFydxDsCWgc7BZjfzkpWd0SoodxhuI0b+jMMbKwWk6tB
Hu7td/K5a8PaUE7BwMDy1gJZA41DKtgVg+4UCmw9gWPORfUg7GBbGowRAlb4d9Ir
YXJ+xX5mQZ6Ls2X2Fk+V323m9jjYwgIjxNUQ0r+khTk08D5A2RicBDArKpHplqo4
tBCk6tvu+ZJr5eH4fsfcrkh+FWJZEPmkkCytTTVxJMxOdFegpYkqZoLUNqKfiMsa
Uji0HQMnRGOOkejBX/jPiahMgP4s1lSjvkgNqrQ2cppyUXBu3V2u8YinxtRqlmV/
UkW8svuMENbCMVZozAcsUbry7T1xJ17G3mdrljuZ0hoPYviZGP48KUk1MMw4B8+2
M50FCfiI8VTeL1B05MVzCSyXGkDWRzi6RGSeSUk+KTFI+RN96A+tjThjoPPHwWhl
Go31GnIJNu+UrvWRoqog/fuqKpCXDup6PTnofTPH25Tmr6SOOvQDs1rQkk/zFC+Y
QcqJMMQzapiYv/R4wblJ7Gpe/MQm4cAKfs51BTyT1GhYmDJ3iNPBSINmue0cEshw
aHCw8Pu0MH85lJqyjgPDFCFAyeHe/Diwj8pM79Q7/61JyS7tu7A0BvrxyMGYT+wH
eBkicW7KVN4ruJL8uZ/B0LqFNz6mCP7OThd4S8Jcpcp4hZtL/RjHRB9Qf/WNQgzY
iodcWgWjXtcpy3Vt1HCViY+xFW0LN1RXTiz8T2FEtwS8xYzEQS2YjOn/n4gA+OTI
tXzKk2fbZgrK7lKXt3mjUgMqXKGa3qgeSYjDGt7zQgK1yyiTorRvFDzpd995cQaW
EzOLD4oxLIEuU9+3ghqROYJKV2EnC250VZ7iJd0llpVnOprhPTA52k6AhEYvtBfW
k2sfnPLeXrTiSt6EC86DDs5UdA5hBdNww1KAnjeMNoOPcT4nLZVQyqrrrXLPOTwE
0XBkvmOu0FoouDwzzgMAsrScAkEgL6mgjxkdBueNtEImav91buxuyEf/l+5aksmb
TW4ddhzPmEo/ukmGjHCCPX/u6wTssDb6ixFvE/SfgBh384HlmVWiJGyukictW6+S
TdbdbG1ZfywMW3VdKuhoUHTx/yYMe3QUIJryHVrSXbNXgEHKgGWQa91kP1pk8G4p
Bu84392B43yVQtGvf6uHKzN6oS439EVmM0Zf75cXsctIkKcTQxPHVPxwLV+7fM8r
pAUwWFp2yVgcPcdZ1DX9ydWDD4FGMZkOqFI4KyelmcCFCBZYXsPYwgyXMFeKSIEh
gD6mM18ls9b7oxKYTPmmf75r+F5neBvH4lakrf/54+Zr+Rc4RfuFQ3mtRIR70Vfw
Ehm+jPnJp1ilcoq3KPGJfWP+CFbgzlv5su73PGRWrYCKqzh/RK4JsAV49w3/ukes
6DKS1qLwEuL5djvJR9OqUSSB04dEvPebyqYLW5tOhw/HFgiD5eZJuey9obS6kotv
g8Kc8iaaJMqI12pB68T3rcWD91Is3tNxBhCWOhHEd3KP80FqjWA/Plcf3bbRY8Iu
3IIsFfXa2wk+fKAElrA/tHYVxGzoabAwwnbkxpo7CEr9Tj+vakHYynpOvPF85qSW
Teu8vu9t5GwYD75aCZbr/SgBhDUqxmuuHYjPwt41t8jQQQBUghgtO77Us0MBA2Q6
L9uNQqp40WBu9poP4b8GBHoD+urCUg/oRTru0C58sccWQ3ShVublLjpXDmeKWKR7
1R4x86jJt0uqqr45o/h+/KsDy38IR3REy+i9Up7CzU6Hkb6em9KbzIACWQ5w7IdO
2A2xfF0F0cKhd47qH9xtNp8hykoaTiTpnUPjjNDbQOqUMAn2Bih8BA7OJjvoJqEZ
gcuGS8LbXPiQcF70z2dwm0DMlP5bqzATvBuFj+yGI4Ew52+wz83BpKA6S9vtEdEX
ptQnZnuDmKFarzpyTeckJTHW/Aj5e8eJd/fOr6utFnX8Z1/Sj7F6I0cXYam908f8
dQG1xoV/x+1mz86YmW9mHT/LsH8akv4oFIfZfmSgnGtdvfZemA6YoF2lsNrEQ3j2
ZeggsfM4Wo6PBqO/8uOTtPyzdr1iHI93Nphj70CrsUOlJd4ap6wOqsSuZbhRAtLy
Kh8h8YcW2xKL8Nn7/KCNACykYc4Te1GRbNVuywdfhm9VLUa9HbhLeILOBuxPys+w
0bQLXRuSOjs2pCZhCiFZgu4iFRf6rZyB0kvMmfvJ+LpJfk3eq/ua7PmNPBGXJqGi
cmHFA3JxhJxWDicjzVNSuh54eT0vZn1cb51Ix/40UsLthera1VjWZf2ysfRdF1AH
JP+YbumB+HIxj4NC+57iO/Mm7QuMVx7kWfcsKa25vr/qHM6PUCTxp6vzl0lRic1t
rfiw81bPEKIuWbm7TDa72INSpXEAsy4AIZOljknMoqJD0EiKk5MwWlNmbX0oyK6/
hQU9qR5Jdy+jI0ts+SId7dHNSMwr60rbUu1mhRiM1UechjSDj5DGi3A2n/KnRaCl
bvrfPN/CPWZq5FmWtghyMa6BXoHDS97GlEkMhAUgeoXA5dvupIfILDbjSwlvCHQ+
d+IvtWekhCFUAnDSxgjdceMANk2lEoGUqjWhk5EmJUO8zAZqMojxNs+LdGAsoNlF
/CGJIqipQSlkxDAa09ZzbhHxtwB2gGq5dtDb6a9YAypXkG8IPp76HTGtbJjMGuhH
hY8EJPP7llNs3TlMvdxUuvz+BT+hNlsVG/hJygRiLylBFKP1AjDoiwTuqdsoM8b+
Gk2XtznGbgIxWsK0lCOrSH+CKdt+dU0/RNEa+gP53S1XXEdP2nM/gPz+EHnq+Diy
BLIgJDtDZGFCoPc2lqdUOeItP2ijsp/aU/X2up76yvgi0uhzbc3a1Q3PuBxInCZO
6UAqzoxP8534oX4ljI8tNsvot69bpXi1W4aFT0odUpPECbdfEvhDEf9X+/4umngn
uLCfF0zlJbufU6SxcuNKdwUeE9A7aJvWnHpuKF0C/DG4UUMbAM2c8kIYDoC2VNAS
Yu717rK4UAmxIwh1qqMeBMysjq15tmdudkn2RTkJJC7szhdkXtZQR6IVFiSAjMVr
DR1j2aT1h4mcuq7zFSMyNtuDN7J+E8dwqIrBZGYLglDjCCmNHFJLeJiMreFs4CwG
XD5OayLSFnQQI9/k6+/tnp52EdCFUwwH+vjGfuaG978b8RwljQx2Jk/DllKT+Hkw
1A52aA0OYfm5RQU8E6fO92isvjULSewmH2PP60cWhqF/KwU5p/yVF+lRjL5N2z7D
XK9dTc3f1NYvN6C3j1mag1rFM2msbqVkdR7ET2s1BhDRl9S8YmRAlA0Zw/iXppeK
3dgBsjPKu8plobFwpjL35vphr1xNi036EHumrVjOkav9rH5ePXWzX84na+mINpT7
sP0Z2pqlnbZYoU5gzH3CW/42lFbiEtctmIu9vehhn2fQinV2oDFCDIoDkw2wwWfV
PzpTP0L/6jTbK9Nz34R1iVAvZCSy2sp7r30IfErB3/GcmVBWb7gT4Xk1XT9QjmJv
prKmkWVY6hmVPSQdmA1lbRBBg4K3kh4IBfWZiZ0Q7dcDdTnM06FHTycVOtk1VCzf
FUcqMQDlrraULjdN52rase/5DuwL+GxoWarH0pfD8KArvdILCRaPAh8lb+0tmXSQ
HHTod7lYbJoIajHU0QKtzAT6CUpOgcgk5JHJN6vjEg/v4GYWB3SOGOeJ0IRP6I4x
omB4W8dPzOxSQOo1GTWSUryFVHaDRWFvtniRXzgHdttySCxyn7ecn0avk/bTp+lv
8tx/4Mf8r76WP5VUgAxSctPG5GU8OCQDdS7DZ0kV7I8eO6LAdQdk+WD49TqT8eiq
8wR4LRiIntAQ/bUxK0LbjXLX58Y3mIiLzspP9SB8NUvZUxBjCA58qDemPUL5f8/a
mXfmXxckZg492Xo22LBx/usViMRe+oQzeC4MsbcAot+8fRC9YN63mzef9EKeC4x3
85flp+h511sqbo76qwYiwEqvrVv3cekqPAjbLC0C5a7hMqKcUGrJOAAzh16dxmyb
5EckULWgYi+AJmmM9G83j0nAoUZLjXufZQDyfThysN081KJE5BDxaT217eLCITFz
IajZyPIsaYMuD69wPRRvhTCApsaqClPHDUV/q1OYfKuXD/fHG4dK536nXZNIm8Ga
uIjfZFQ+viTTR0/Mnp+x5T6fGmiSZPXtIa6q9fgXolYwwI3EmVGkgm5HDJo1Lhmg
wGjU1zyQhZdU8xDCdQLazxKp+wknqOl/7cFoVIpQYyyu0keCXHYCvq1gF3Dt5Z9w
zaESvRJ11iZT+7o1NPzLvCca0hetqk5IGVaLVZILWiU6znjCcIGMFX0qD5QdEGSo
nHodJOkV0jcoQK3cBBAg5TZUEpm96+TYD8F6c+PdAenquHAnG369/I6b9CvVSxo6
49yxSRI87maY4FRWBt6fUyNX548DJr5XH0pGUlGKDDI3/Q+VKLtmh0VeSvjAEMfV
CyVMtSQdOsPpXW9N9oxTRyKVrRtPVFb/GlXsLNA2kM48gfb/5OVnd5dtFbr1YN5F
1O1+aV0ZDUBrlaoKXgMTmTNJb+w5Q6h1CokYyd4SlAVhG+JgcouwXVYG450TF1jS
tLEA3Qubxl8pff9Cn5cr9oj0jvce+sY/SgZ/31O9gOMXclpWtQZ4l9ricpGzSB0N
9ovq4Ob83dtbjpoLGAbhR2tm+LfJeMOAI2mOlfSFDqlqHvAeR0K6aKiOYIXObBCf
5TNmT45z9I2sYCRuD3zCv5BMMl33QG7n/7A1UEz94Zm9LnMV0Ya4+fPuTD7wyU+J
NaEVcN90vr52AKajJyqCL8UuqorFrWwBYixIjLtRVDFJEq8+lG15Ahc2dWWXRhem
KOrQ+GZaekFFJwd8xwwI4pY1tPQPRx9Suq2WDTHyHKsdjIafGHKxdIGin7GUG9s0
fWpfQ+xyjf7NUWdb7G4JALBIOCfk1M66MOUDSznr/PQ9eluxR5nffRurdkM3fNuG
47V22890s5LwzYDMTnuRkex5aKwnhdYyAbdUkLvZ0LbfycBrPymcHg1dFamFH94g
kdUqg3r3kEaY/bWGN/Rb/MlQkT1iQGD+6dGO1gajh11S1sZNJx94SMXA9fhAnuqk
2wQid+TiO9vKZiATIj9bjVg1kC8eNXzhLzUMnDpaz+VUc0mm5d76zzeDEY7HuAJj
0paDoXTP/Ygn/tWHQIWViRH2BXQ4BOzmDOpX6lS27MLUJu/oURLUerx2tkQs8Jtc
Yxkc/QTEo0s0aTJVp36ZsxhhkxJGLWKhlc32wM/TG1UR0ZhVgfmdfY0GR00F7wSp
tqiwh9eDjZHZNQauOStcMuD+lyE0sbXFo05+KVRDaqj6an/4qoMqiYXqy3D+wnQ5
DBp1Htv2VT2h+x4NaRKq/HxPnmm1KXJg2obOl8iGjmQpRMmU7sJNj2vMK5tri6Xr
X6xX2Jphzuts0ff58bDjT9AlHgXb67a6VJdaVnCzZjeP38i7FqcsIPjO+8pKWeJt
WVeX3SxrTUzvw6o4NcHAXofU6/j9iqKDytWTx6VUra+1csQu7THux0l/QLG5Gbyi
ZIF9buxnKls42RhjhCUhnw0cjmOogJY3bod7T2HfxD+KgBzOyVTiDuw7lZoXUMiz
bY2m9mV7MGEm9JG1dR6Cz32WTwdCCNmSWYdtn5PCyuzWrgx9mrxmk0411J3qc4R+
2stGuDArVvjfcooxvZKRULNqturN5lyfQsEfsWkeC7Y/p5RDkYPIZ3/PBJKorLgv
YwXnRzv4zY9NBKat8jWU+TPj7Hs5b9QPAKhsWu2tKqYsmrxXh1yXKIYRVV9oTcJK
gX0b7GUB19FPB+lnAbHkPAUcheUVN+XHDes/APjLl9udMH+vgCQKohDLERySIt7W
uxnXTubEnhBPzLDVCVm0gJFeMnM6nIGDkttSUjSlUC86wOJSz1C7rfK0Q9dZp3by
67QnM3hI4p4KgrzJCVYE3PKioSlFEjFHDDVuVdlyTNaYY3CIWUhVW5ZoJu7vYGya
b8AkP9ts482phdwqKd4I7Se/iltud8wYC9ITR90TsyKjT8AiCZrXsSHN/ZmiVs4U
jL53nP0eoYjGq2HbitIQr0TXbXUhWWWH1QNUKmUV/vPT69A11TWr3GHaKasik5O4
4aMBZDMHDWZ7whgSqXcGCziJkFYNzFSkYT9dleaDMwb32hkwjuKmhRsv/ZcQlJnx
n0lxJxHWDo+UjYBe4q/oJnhGoTeUZOj+JVQxQeWk8UZcCXOWyj1r+uyYv7ORkpeL
fVAtUygAeLkZtN1EaOQKc0uHG54xi9NeLlLAC1f1QCJ2fkQulm01wEUXnxWmqOaS
EYlmLISo1qpMbdj63yWPNEAESDk+XA0nQkTfSfWjotLWExstiiQJwDmJhQOK/EbS
AnZycXFz2vBEzrBappFKUEbM/tW0APQUODQCZ+NAqmgiH3XHn/bvaIJeJA3e33mo
YacG5xD9zjP6Cjh9mwdwJYjEKvHBDMLmWpsmcfApstn2KepNd6p5CDJwKvJ+aDhZ
22Pr1ach8yOwpxmr6oH5jrKXb8coeFXEyCTDIdUTM79Y3oZZK0+8OxyVcIfEekC6
mdNPLpvZoX4BaFkriIeRCN/Lh4HdQ2n5TZCn1yiuwaF4oQG/X6fnr1Bhhbt14JFh
UX/A2OrPcYtVn2xeJHedAtVCkHFs7IKI4iB8w9ZAjnQLn7HdAPEDBunFwUJge7wD
G3lSJUEqM21ffiV47rUethGbkAzgu/gKLeB7Ym2kM4aAr68aEmtrh94s16yBdPtQ
EY/8Y9VL/e4AI0R7V4oCuyFT7jAAGGCchZm2s0GT6Jd+yO+xr5OI6qXYjCjmhipM
mU85yq3CVi4AE5PU0qxb93Ld5/Z91r/KLT28YT3DxbSYiUzb3G0om5v7rQbwMH2g
Olzbqu4ISOO6ccv1o7bn1r5kCGRNuiDdsd2Cst9H6uPKKyxxUQ5kHnmpxC6/SGj4
ed0FUILA3nxuTzuBQSrjOQkArJ0QkDBiA1EakBCAv0RXbM+CILKHM4lyFdaHpk2/
I9SOrPS2XFyeTwGRGyy1SxJlp9SMI+ZWuAy0Ejp7WQHWb9GLLG0ygOAc/UEFnvH0
liFRsreRByodZhfxuRdzuic9NVhUt8HF6/cCGKefDiSoEqVSAODCMeVHLyTWAxa+
RYCPvKsBJl7XjJTXYkXnvHIlgwBptbvsV9g9XS8sRN4MJ2i412Ais6BiagqhoWQy
RcaP+xDculh+axh7PXqba0+nUtRAS635yvU/GcHo4+IoW+L98DBghn1TjcCA4P8A
banfDDdPlk9UiY5AJ8mSoaZR53CJlkaOt+pgvsmCaZADyNZ69u8bMldECdq1sRgv
un7cxQHVq5GfrViCjse4iU/xnMUH5P+kFW7AaKNkQ8AhY/vTCxzUcGMakjlKitMN
Zm+IRuTp2/XPAgFwmEShdocttVGG0fs8MWq/Lney47H2JKmdNH1qeRsD66bxJzsE
6h74oXNgzvTXuNofUsGHCMvLGGRN6kyAISbTT5Uey7aNvi7XCGGMjCR6e8d4vw03
ZxgtfEbYE2k3jkJXNRqnjbbAfdVGqmdTyRF0yUvfGaBZQDGbmMjzydBKj8F/N6qI
N039rsw/4StPgQPQXD+/s+w/hVnb7vgzrrEvqj74hFerxO/c5b1XtQfLqv//Vl8p
AC5QaJeX+SN5B6QUQ4yQbshGzBERtl+jUv1cd+V2ncNbpTNpC5qQfR+D/OtAJu7G
jpM0GZje7zH3OtkVPV47zRCAoqnxYb5Ydz/gY8RV+eW5e2DMssJSy10GiUo7TLAV
q2hZ7qSr89Bep7WibRzVNlXw7Lf/YeDm5TIfdrjA0e7meF4xMbBPy7pThjHHqi9X
pplSHk9jxsmPg1l36kJbBRpCvNgOQ3oY6xk1TadLE5J4ITB5e6G7vS2ArSDbrK1D
lY8TpmS0Fpqa47NqE4k/p90teg9lywNK189THmmgFHD70Z9MaXT3ONI9pSVirDUm
Wkjlju09R7MCaH2Ezmh6YjIAzjJr3cBA2/NZKoWmXnLo7EceS6bK1P+fAdDyn09c
DRYC0DmK8INs2NI39mT01nhF3g6X4+y+nfNncQu7i9msImbsPXBEQrhAvktLSKRk
DTHM3g9uwFfQJoxt0Zy9K517U7c7BsuuvXz6Fdzv4rFExKeCqlKTWjw9aN4rLAw0
8qEgBn8pp8DwKIOnhqFcynl5PzvKnBQcxlP/s+mLQreEwQN2ZI8rwd+AA935nxM4
9Yw9dvnxLh3W1l/hFnVsCsa60eX19bTBw/SLUTTpYVyljRqyppk3lUQEnpqi8PPT
AIbr3CjO25C/dHNAPo6Cw2ZmO/Mwd4ZoFs7C2PbSn1QexVoDoEPKA1pp/50ETTXC
JAq4rvtjfvmRBZFzHObIahYDWakVItxT+yBUEvBGtUhbnMPXzji+HE/OjgG024yO
ARx4mD7Gfl8/JAuWu/SqrMx8JDWJouJHy3q08ceSLnWVNq0w6wlAlYCsyqoEUviu
yPplr4THpBczVCLis6xEBAQlEcZaYmFUNvlDKqK+dAtJr2PVnvuJtLxJQv5RLbw3
DzCd8R6lZ+fglFqiCKs+SEoB5auyyHIukbgs0mKq5+R6Uzc/7PVX90z+3e6e4fbx
R6F+fzDDFP4/Aeo1aXH22JZIVQq45tqt79xH+8sdCtJdxQJrR1o5qV2EmCL4o8M5
31fVcacWoHF6VvW2fVcQk/I99TB98++RFXfBUOgjapPSBBscbXw2fybLVQFG8AI+
wexgflQMPXrDqsM/Rns3P1KIAkU+pQjgaYzwZxuGGbFH4aSomVlGqelNPWTYaw9v
fMAeQSnASxhjE4mfZVhOzIqNYmcf89++GAqeh6u8vMZpMDXgJGu+Pxp3Ci8Af7iy
kLSC0iuc2UR5p71aBv9cvwMYVsvQClFzrpad2rDZAdM0njNrcyaV/PEIlI0X4nVJ
KoPltMY5iLPLVPfA8ynZMGT6GdF/0JHVkZgJLTyCnpQzfjRuG/a4hzITsOFHVMMp
rhxMJOsyXi4ISHW8gAFoASn2KMZOum22210Jy8DHTyUdex2pvdB0ZbCmvlt4hlyI
PJcN5Uu31VYQGHLFD2dYJSgtdYo5VNg64C3SF9RdWQKTp+3+zRBHPuRwfeKoCzci
9wj4WVQ8hdPZd50ZJGCkknVCNyg8AaeJ73xovxSqkh8MTfUcPCokbY4vSKRsO1af
OD0khlWOiKM3JXtN9OAeS/+ArEACQzt/Hjuq3aAb24zFEFy6cWbYs84dL8jzxfdf
O/hmbXsjJiVVQ4FcFHPfy3TGp4+5na/H2h1uEnI/kqNRrWVSB1eUw7jk/SP2Cj/f
+wq6M4wcWsYOEe8JDZxcTyUltfmNoXQih+Dcu9QyCRX5Hqme/gw1fnbB18/Il31r
wl+rdcNzHDJbV+Ha7Q6OtN6E8hoLIBYmLoS8eazc5T8nWc57m5+6kN56QT8VzwNq
bdlo1Nokfb4JtyX9JpiZwSd7zoAmMQLq1/z9XmFib3u5PWdbNG+45XBAV/RKCLNi
Kr+udV8l9VtZs/Viz+8u2+xBD2ooY4VHbK7oVvsqKpDTz5hj2WtI884BefGq9aho
qWwQpnw5b5GcJV9I6oardEewBYxpqWC+dkQKuL+elYt9nQpgdwh8m04f6XQn5HBA
RKDR+/T/HNQ1vPnD1Es4LRSBTluFH3L+gc+QpSf8PnSKQdH1CvNa4P/sjWlA5XIb
Oz5cUbif2ZYqAowG7xl3YUa5oAIPiXxueIPQWZgwD1wBlz2RiCa9+SDebke8O4tJ
rR4O4eG4jc/FwqSOI7MZKtiyCOChbMpdaM7VYC+X3ArkuLZxa+QtBlZkIdImjE4q
pHbKWR3E3QHTGCPbT63bFbhPQRaM5TtldSGN11UH19o/8emC9G9mSntQr8UbRChY
6AVe+HGLP/sgoVeXYbrwY1wyvTpB8OU45Co1+raUZk65IKPjTgWS+HeHUfdZfSSs
7JvTX1s2+1dcof/FB2zMqgmLMMzxTZb1cWxl1Vou7tBNJsSSrEoSwzNWirBiI2r3
RZhwryJVTm1DNBPqzGkosP/Of6ayzHoUZX07V8D8HPrpdtUao+GfLrNELdaKLOW8
f/nMcq1JvFzsu/CFwqumMzri4sdE+ygmJgF1jjYpjdqlLvnVDmXAu28TSv+bGHOd
6nXmBciSH4dCj5idYvjvg8JnESByxSvRFx7s4rFjGtZ2HWS2LPoSG1ZA1GQd1jtJ
oQz8ya+XPpB5dtsRtWTtKp9/rdwzKH2tUEPx/R+obrtPV0vKtSF6gzpYkDWE79Kz
KwZ1lbDCcZRphgzulTtpTgFj2jgwVUSxD5g8+sTcH5fGHx9NqF+hvxIUD7af2gJS
NqP8cHKxc5wIfcajJILI1fofF4XO5b/iF6Amgvbx4N590hAqzHJXscjvBYUnlvck
CtZafwm4cb1LuvlaU3Q5u0PRJlItQoHDspNy87GUzU65Q8HGoGD06lTxGS8I34k/
f2tjByIKhmG5vDZMpLr/s6ipG0ZbU9t1IP/54W3M2qU8p2ImJPT6fhX6UhFi4xKF
Wb0EAc1L9O1JqMD/M0atQX/nUGmApZvi6akOFq9pIPZ5BmIwX/YmQZJKoO9d/w+p
WYOIpAQx8BLmz/sbzJeYdbB3wi5wSwYpXKDA3vRVP46+6LNGNJl5p0nclioySKtv
otGbUvkGhuO9fEqrFNmw9ip2CJ0eeZX9aVLmjopD9xUTVKreZ8c2fj6zbYU1cdsl
L8NLSiI5rUB67htDVBG9VQFgTwMy+lt3WYv0ypaw10ON27Hxt4FZFMv9Z+IX3uQm
gxDpNRIM/VuT2tIJMs9odQYCzNCbCWgDRaIEZgnmqSdqY/GZ+Dp0YZ0TdP2k6VZ4
oDhf0K8wmQEMvO88UdUxNeIIZw1RoCiPLV0Oh/nOaPuNbOVeV1vr8bYSaWXi4snf
RvwuKkobql0KxmtO2vY7tNaowaCW6ZhrAPa7YYGE/ZIIJsMvXmnWrExuRXBWMxLU
dukqMoz9LwwKrsrxAjjxXCaB/zuGPjignFljpjtloD+fTEbI8dgSASyDvxISv3vJ
3pkJwSQowxLA/wiw+3H0JJ0Efs45IEFMxYSuTnkFSiYIS4oKEPpE3b9JHzWzIJIt
Y4qmJXCpmkKykby5zWc5s/JoVOdxX1nJAGJBY5wXwvA+LFLEfLuuUt4ziNVNPXaF
2vSvmHcZM7d4id2WXcGnQZkFcYcHgrxVi1W6CGizMqINuRJ+zBMr+kPs9AO2/gyL
ARnU/Q+q4ZX84mrBgBlq4Uck7xTgE+JPVzgmpZq5mhkuWEiz7uQvQEbYYCXSnJOB
4aFbduOhE1Do/wfNWv1gQVD02CORKfw/dOnQL5F2SHl9elbyoCQqwuMYfMeMenFp
MCcSrkDPW0AldJIV7dNWaVDYDdmIbzdJp9NnLtNcCb9Mu51k/lyUb6QJo0Y26/w0
WIJYHP90WVJvIVAwlNAE8+zuKFK7IgsfW+1W0ab7wZe+xd083wXlrvTxwFy9kt7Y
WFMknVFR33Df4RH2YrzrAsmtR20RldYlu8LWBjbS7ydkhJCo/+w8I3eXdfhktebe
Ekx0FKlR2zRAzz4jOGU2MADyU4/3jjTL0+2FcQnIUxKFFH+4zcOVwYGyCXPp9VIT
zS7JM7Z8iQR9OLXDRjpJiStgdt5gIJfmoyEqiSvyLiZFaKseUMzfvBqlq5aDIAmL
mJ3IJ7Hws51yyHPulb2et6/OSXB+o1VD+j+dQVGcC1OU+FoNRrkNSzlroOZdaBI1
Z8KnuXmZ9+6vNrkmj05MYtS0VFja19phMAoCj8EYL6mSlya4ZW8XbK9m01+XrAiR
0E3x0qRsipGr2nnjR2LkA5SHYnb6Q3qj4EMBZRBHA0wYfOMUBFIvcB16S9SeDF5Z
bCPs9KOgSz49KHZBrV3+rxCn+fPZHcLoKFXYcOGcQUAfpTj/OWhyTm91x4bfsVRV
af/pKk5jUWA9loUzJ2TfFdsoFSO3cbnBhG2a5vek6Msu0P4SIxWw/+Z0Yz6XCU/m
sYVZ94J7xNpMMw77EuiLpaiHalSqpyLwfFtAaakeumNJeDWTlO49sVLL+rEO4An8
j+abLVE8PrqA598GkguutzXO50EyiKCYvPyiixUproUb0bpSchWZ2Iq/PsUzJ1H0
QTCiYmpyjkOqiIt1ssb0Y7azRAdAaItVho8rm5Hk2QzCkBNh7r0xDULBraihdcPp
kCdkfZs3pW2dpjy0ncxmQcHNgNsDUsktkYSITNAaOp0SVh250rUPXm+Xdskq7dK8
LbWoA6SqUmDoeV6xBKRNFqO5ANemIedshd73ffuLJMORI6CF/1R1vBIA9zIguYJO
rB2DNRK3bLy/JSl/mlNziu57WE5BkblDiTuHUZAaKyPkk5VQuQWDj7IrQGBWfrjf
9vDiIq3UsdvXLwZdMx9EjQWMww406TkcjB7R7b8jK76vjgd7cVRNCsUaZ65fGYPT
Bj+We7kUzG9HmxpvtqzhzgrFt5ImqLnKjVr0YBNaLk16utr6DjFwqUkFSbvfXSkl
jTu6yy0B3wYJZurAdRS9Wfg2tHrH3EiimgwSvgtg5Ygrd/ZRyJqux6rxy7aM3QWd
xDaa7Qu+G/PrblGKV4Uhgq9IPi1w7khq2v4sw6sgfNLhnoErrA9h1Z/3sZ5HiIYp
HWlKLJI0B/Af923K5IcigvyrvG9Jhtd622tV23R0NSTc4SsxwQ+FEtNSsd29ZDoa
bbncUax+J//R3q5uTXz/9ZkzGDy2FbTMq7QXkolVbypcw+56z9TaYYkrSkh1Fguj
UNlO3gAuulcXKLRBJ8tnzob2exGTVJGRmK+53ldyx+6ctLtHtxyrYxq+8XYWwVFP
WZJFD49WCr4pZJV+GHW6/mLorcIJ5M6cM0JOL3QT6Riy2keiA6xqHJemmUS+I4hG
boF9Za945RLWsgtad9FQknQFQ2rudhXfto0DI92OH0tO/pAZhJuTBUbvG+/bqPeH
0qjjnLwwjgwF9I9F0fWHo/K+n5ZjJp6glx2CDi2IvN6DUQNiNorgforkI0gFJse2
pkgN6Ye3oLFMmqE9if4oxwRBwP6Af5UrFlbxreRp8s3Fm64I4V1ns6e1HIS6oC01
Gg/2PzAWZZ3qYyHyxPheJl7nqV0GudDCs1NyEA6cq/Vu46PhyaEjVGKrBNbxZ7Y/
H4VaH/loc3NHwUm0dJ8VLgpduFxZcbNnyUl2yE4yh5hjrvEHt0SpBnJ3wmYL7Z/p
o5dQ5jKAhMtJt3ItOC30ZTA7Car+HR58s98pqNyrFCsBM5Ue1aBMQtwKTvbu3dX7
jBC8X+z+GO+zlTqj4f7Npl+hcVssEbuADVQDbfwRwmW1/NPz6EhTfU6lakzulfht
a54phRBqD6+V094jxxhpiIS6hcD75CA4QeQ5Y0vcVAH8ivWXISbjjOppIGDekvMV
E8h9U2A0Aoz4mG2DyyigxquyHl4VhIEMpurJl7nd+V9ae0hQaxLjPdOvrZCFdjGF
gzQ+pikXBJIOLDjvs8swZSonw12adaW2Rn5beS4Xh+9Db2Xahuhpx5+kWmL8y55E
mzi/8HGoBObRSsmV5f+SCGtQqyF3unHDMJ3eLIImuJANCsuM6IgpJARkdjr3amTB
mOnFyNGX+MOjgl1HJHw8m6YHROZl/mB6C3R2cltUlh42Sf7BxgN695+tOXYR3m13
625vvZ3EdWK1z2qLKXArzfeM/+KD03z7wvtE1xY9Mm5N8iv4G2POGFFi8hl9A14t
/GBWepXlzswT/DsolC1++srVRJXjF8+R77suC5i68aCSxbgNvnCusO1i11bEESEN
pogD3Tzoy/RpXFc2Ey8vW4aiCKNb1V8oKr+VRRjb/8QNC0P+4gbA78fCQ1zmqpS2
ElyzrLWkUbHOC4mEOFojd9sa47QEOGe/ubIL6WWhotlqruC09/DlOYLwt8X0zZNA
4k0m9bEKyB2Xn2dfe4CJA0wX/PddOiLO76FTee+Z5hM4pkA4ydBmxdbjdhTwzsR7
c2NJCXZr0vAWuwOjbZYravKOc1gOGlzMhLCUYX2kZJ8PVS9FzNQxdnwlWIePDhCa
DXaO4qjrvHWTSXSnRPfmJlDwgJHKWfH0zz0++iUqnjujUrKSZazJ5pjXj82dVgEG
RzKo6s0yVqixm3+FjfKDfPYSqOPG+PANGsTG1jM9A/kBdtiAwsuMOnr4iFJhyvjw
goN8LyT7zUpgOXX7N/gBIf3f0XqWgoTefJ1hWzjDDNXEcE5g+6frwHvDhAC4ZRwG
oyPJqLM4kIAUkOBEwN2+gMEtw7H/tubo5g8V4p9gizODQuSjO7CbYKU4qu79CpJX
zyam3C5LIT++eFKUrttUMKwnN9OERIOmvmOv4GqNYYpk0lS3owYDz6LXQOWs8By5
SBTR/WB18zfaZz+W9It6FUBSjsUkrE6tvGOXpIi9IppOtqVSfLXL9HZs2f9W6caZ
t7wDKL3tWpMYibMAmA/zaYwdq/v9G1lFXZFwN9UU0FpNpdkPR5r16AnGR1itKOcb
JxE7RhCthAvgrfF+oRWuJ2oqNAFMxd5wFUVj9a/Cu1fJBaHl9nJNh1QRwRRiz3yc
DYRafv7JJUBP1+DUN7if/sgplT8ttqPygJg277z/tK9mJvoxN6j8ZpBjwJdprUZ0
XhTeVlrFGGrWqero3eDA4Vs0/AN3FzApz9umzDWVRFEK5Dn3axvWHz0bEY2a0x94
GCj0r2f1fq1UxWTTT27h+jkkbFqg6hYT5vuua2tN0Y0OionoN5gjJ/9x5Byt/plP
6EKcGsKU8B7VHeCapz7+ey51nzBfe+1cOUBHKOkDxo18O0bduvDr4iywxzFHzGi7
nLs5R7sUVp39KRvALqT2PnBsDAS1VkcOoF08MHdq6bTJyVzMXvWPP7Fjj9PVLuGx
Ja9ZPPQJbhPJ2vaoh8jN38XhyHdaIp8dlPw7bK+f0AmBOwKdpAJp203MMu0eEy41
FEpeieKjpNiOTNI59AE7ExnmaIL4rzOitJBwbJ9K0CUWRz5FYBHVbN9xQec1VCJV
n3twuTLX65IjOgO84Db4v9MrkkNpF7RhbnXToaJ9FTBObviNAcmfqMh1xY59fUuR
G2HcXeH7qam+RjjgIK9Niv0MrzcZmWR/pYeGvhj+gRHdtS6TPNiLQEUIihHeQbSM
oXacpBOnMFTG+Q3/GiSUaEnTgvKedsJVYOA9/+csWemQE4+hVvCsEVA5CWO9c40g
a++U3r+GhQuYP9ewf9ILH5Mf+tq2BAOKuGtjCv7E5wS4J6+JbJZ2QSyXRdkSPPsX
eDP88JIAe/TpA3SWkUuDfpaReCixgy0YV/9dcHZLVQ4VtgY1xEsnh/j8bv3jz+mS
zerf/y+q0duVQMRZkVuMS0wCEVTobUBWZc40FSMntpEBWQHI6kVmCuSVY/sdm+/x
IaprmL0AStclNnKL6W4qaNYV6A6hI5PbG/NYvfk3nt6JDYNl1+DiSZz2cRqVJ5vr
2BIIQjgdC73+MesMTKhJIXbinwKUxcwlX9eQAY26V75UvzPwln8xGyALfY7VL+Km
IfBS+vh+XhwKVadOOE8A/X08TQIySPmbv1fgn4J0LhSdQnbYFGpyR0yU8iTNeXeF
BbkRp4cytA1r3Meut8YKxexmNMcv+nCC7e22NqzV5RlxekPIMSTO6qqsp6Hyjjde
v9IVOXIJVDS8PKUpl9TK1JPccRLwVL3SPRo13B4EwaGk/XOVpst91qk+bWcASqnH
3PAhiqOirhAy5ne4zerL8GRXn9rBEI/lhmEGNFrznv+aWbEAdCjZv72Bwh2JZmBE
vMIbpTHgYwgjZv99gJ2fONSaXLZ1V0vtMQDeExk046vn4oVfZ/h9Mc3wukL4YAS0
inQ6a5akz+imDXL9dLdsQ1GNRGGBQl11u4hKm6LOmX2A6ZULS8nNUYqiDAif/SbT
Spasth72BBpD42ihZjDBHGF9xpyxo2Rnlsz19/Os1ULzwhKpuv9EyyqLTo39Ul9d
DEtH9MDIZqXnBmGb+FWiFyrDKxsawU+EAABASsnpXFU+PvqrUjvC0eDAxz8R4Xq+
JRs/59aikPYnb+Ypl4wz3l/hrntgY/GWqckEQgUnCBADmPhN3wi3do5Y/bq0Tos1
rUuT+iJapzg+lxG7088qKHepyDmTDeQCWRL7usAL9YeAvuYLf/lByZ9iRQPaezpl
Y/5B5tQqZ+o7lGOVM67BULLbMfFsLGveVOu+PJ+1RokY+vGyjwN4R6oiG9DyErkt
VdVEh/p0nhUULWPtbFNal5spSlv7CweunqQ4YTOf8lq/hEGJnN3kppq2ybU71rLH
Y7/lgi9qx+Xhbyr78aTMSwIJCasOaUlc+SxSVskxEnanqiJMnb70uijQ+JTj2g7U
6CosbF+x+XP6GSlYzqQJWkU9gF2qUsHSxs9wWvXSnn2eT9zh4IQpYk0k8hh8bFr8
hQUjPAsw9WXeHdDD7aUmVZJYQc4ArXMvYs9PJbfC46xy0VQICgg/d8ARLHiHK2E2
rErt0r23ZR/PD3hsfe7Wkivl6ZkevOgIz+X62TSTutO+d4jIY9IC8FDEKtTwr8Vv
JrO0LHmemQe7P2hqnuwPiiv6X1nw2uywPoHTV8R08IZJ4ZJDxg8FoSjV2nN0yvIx
RkYpsbfYdrtp0hmVpe9nQqQZ4Z0y7QjUpN/AFtc28jDbAURyxsdrIKfDqHs8ml9R
Dt10LHmd1Nch2hjAXnfljTEZNgbw6Pib8iHgl01q71k+DVUAAQIsMwRcgn0wFyHY
7VdVbJxWpDHRMyu+hQtVijIvu7R+2IagvLnk9VzXTVvL0S1EPwEMEEdzK3cG04IC
ySEns7L65NRpsV5/3H+uiVETdR0eKs+XVL8u8F9vDYmRP7FvHLEGqmqUrs5Mrgj2
17gzmSM9oZyKw9xQ7LqGxQzhBR8SrVNsVjqf+ZeacbPS9PVbLKiVAtMzhZxfsNDK
OGXWpC2b2Wg8DD501QMShidpi/9HjxGLmZi4EcfNPxiOfJDKlERaAlZC+smOJdzM
8RFc/IYWCMQEaL6QhPthyFttE2AgwwcIjdplJFqb6tC2JNNQacfTg7GS0gv/pBv8
xbSsapxUSyiuQ8St73Ff0yCak4fjYaeR73qYGtWYIrsRPwZj4ocsxp80ILNyHH4T
yk5F0SOc4kVpL4gxy5kP109zsdr7zpTuS5uevpSXJfaUAGn9LEv8vMGCW6CAj9Hc
qp3rF5q75rlr5v3gQ4VjxRvxr/a0GM32a5t+VO1P9n9YaGUC2dE/O3BkGPe3c8PP
I+29lNYB9uGdvjs3m8ULA9gZqSub0TfJipY66qhzSKU8fTZZi2aK3im8Ekm2KhcL
wXzLQxXgvqfKcqlqwirCKewn0Abj6HjBYG10+ZLGJ2ow7Uk/wTY3GXelkR2FpNd7
NqbXT0z4EuGy3g1A9ojstlMQj9GjcPi6HG1WGAILJ9zDVVIAN+etuO+KFLBvEc9r
/knrHj+9UauQSTPpVKBohbaFTqXI3x7EznPQct4NhTfMRohwlvdRHxOmPprmVP3W
pwA3uUoOnTWcFsuRLiZutM/JnOAdRmyPEZioI/j0a2lbxVyfQ4EYg51hTZ17rhNB
avtD4Ou0X7c6Wq42FDJUySMFwfnuunXCVRV2uPdLUfQtkw+ml4J31R6sx+W7rwrN
u7s/AYw1qDwE/4Nx+i/yzBS/0zBMvy5Hd/gojT6WKbAQvbLJv5DvQafqf46hIy8T
SPNXD7AtO2R/EYSv9pt1iE1nJIWHh3Y2Y7TsSIWNoixp82dhrAi6p86wjY2jDZ6Z
o5jWX5jGn7CC13ECly9wrpLuKIhAoXOwlgDuotvDg+EIuyzxM70TLL/6XjnfMcuj
Cxg4HnU5P79sJ5qiKeiokDI/b9ceTWhrgEQYKdPl/fzblbPIl+wuuVRd8LxtGE1q
ZzsuXTC+aqDAoj2fuBM1y9P7TKu8vLGn1stp4lumsqU475/N+GJ4UDrcjQX5Zv87
r/uNgihJU3gezrQP5nGYFYUXiPpI4NimldFDDsUbWJVEbEAd6Nek4Okv5WJJfFEL
dgSkGZbotX0j7a6o3woZZcUh98dOMmcwG4fk9wJ1tnHzyx88qc5zy1DHs/MMDZud
h/WxQ5Rgk74F1cYmfPUICabfQm7bk1sEGOoKsoG9+Qj0u9ZERqukiyfi31xzw9E2
0kDVGuuWnl3xYKEo6aD3D6//1XLrvnPwNgfw6jpRtlupU3PkIrmzXK7J6udgU+pD
GypGa71RzdKN1GFxToWCBvIIxhEOWx1BuI3RKLsr5YqIKH+zptQf3orSIU0plUXf
RT3yJcHa2auj7X0FVXMq58wGcnaxI6xWV9QrW9jiFW4roDr6gE6FHGI2kLlZ9mDI
VjIGw+Q8CFnd9+2L0olBB2JTrTr57DcbsJXNBbMvyMoFezq+fGtVOqRuOZ+0Cj1D
ek1mwhdAsFTk/vRt8srDC41P7tQ9JvXO0DSABsZMiLMmW6faKxGPcebU/J1WbKqb
VS6KfIk+6XqCxkDinnIhhtIsZuvsLSJhDik7/lCM5KDZtssL+tyXrF4d/QndWGM7
NcKe2x+F+4Va9nUBpz/BP4MmFXFPeMZ1RiIRhu5Vzfi2wAnDHMoaWgvJYMKqON9h
6dkSkqLGVsrHoN9xx9LBvajIL4s8taXa/CvCS6j7AZxwuJg/1gZP+Ohs9Dj0/HXa
D8RTPDunq1krQ7kcMKZY+3lV9xBzyC/8o1mUUU65TWsIqpA/s8JLO1WHV+nqqyMA
WAWLirUl98n0yh9sDRnsPiOoyAbH12XDVjSkYSGEpTa0s5E6eCO9D9w2kHZnwKjj
CzEJRi83VLtTIwJwyJ3I9U6KHhyXyMfWKyiYqyTEZimfcZuXP10dNDRb2QLmuI6E
qNsH3n6IpEbbFw8pIXbN8ov9l/ovVyeP+Z+UNcwQ6czMbyZQrOBBWE9B+iBnUoQ/
q9fV8l+dlLLqd/hrYpTMPtZyU/e88Olfa1taDDdiY17i78ssK+0aefEhBl/nHzBn
idaS3ekcprmdq/rND5AxDDTniaNuAqcDaZvj5hZnyJp7J2tajYhCBq33X2J15RLO
n8ErAAMliSTb491oo3FSYqIUO178hTKizji5pXA3TOIFXQmPfKnnoyLst/tLNYjo
duMcFzI1sNC/BMu8xa7B+qwfEHDfIs+iG+qnZMAZ6LeO6bjmsgOScl/poFIYBmuK
g+xUl7qAHXFTs/Yg70YZDXActlm4OXf6skEInNRLlLeZ1UxdjvjOj25l4+2hzRlB
UUb5hKXSLtEquul6KGfp+9kleDQUrXARC0xByM2cjC3DmxP5nC4Yf7jDLnxvUOHo
o/ayKkfoRDeQ2uEidQncBfJ4dg8+Ru1V7yABeeYudzxuqa6KZ6d6QUvXyt6Yg/CM
wrHs0wqJFHvP05CmC5TstYRkjB2sDFiT3vGXoqxMEIkZwLIWu2hFe0Lm/ZyrOzPv
LUNREWjSMyEkbmmOy/V/eCxqjQFJ/Qsy3ucHUMMIll5OYKQDdv4ZQqfWm9t444p0
WyTZC1ovlidRry2/Frh6pNnD9dwjjyn5RnqDbgdjFboV2MyyQ87UH2yOZNLQEDPC
BUYVKv0vTqrHo4t2Vnw88AFP1IJk1O8ZReucpk+Kf7wW/ASInldHQCYSkruYJ+X4
oq0rlPzKIL1btnlnx8wBFCQYA7y+fOHlcK/rIF+l2PKzIeTvtipWi2P5THQyMwIl
1Rwg0Cb7T8vYJL88BwaAy1oKWNGRkxLV+SfzgZevNX6YcFWPZZe9EnLJPkJDe/bU
7ouCCIT3efORu1Wf7qVajEYoFyumEkd4qAAzG0mo6Xi4hOsqLvkVLgPOfiZQjRQd
SBhGqKm/jN5zm46UBqlPXMaqQ3v9MiKD2UkDgLsFZT34j3ZpEsd2G6QmPoUhg8vq
tp8mIo/lW6foqS86ussRqWJMDLmc8FNQESwDKV9suNh70vWO1a8/wq9JCOHl+orC
6NQ8TdkinXvh0Yh2OSisdz3HldMURHq2dm+VAWdqb7F4l9iUh4PGCYykMOorowwt
GeFQj0TFQcA5KJQrAh/dR/2N4nSPsuNC1beLNUXDlnDu6CLNQSrp3aFmocBohRBT
oJRzf/Xb0haKUScO8VxoNdKeYqfqE0JFeJCJ2NN7DuRLuIjz3rGMyAR50GHLUnJj
wDcn8qBfR8MKwEBkZI2lQxX0vtUGLYonrlUaltvb6U3Pa8OpmvB4rTBlS7E9Uxiw
m1Guh0hlGUP01G9U1Ndrh5Lxt4jQz29riE2Ox5GZYEI0Hfv2OaH92QGO/8YHos6T
7ueI1htW+UFsGpd/qD16xD6AKLs8QvOmzGAe8q0lt/QpZpIfp+bSvTO+hFLlmU+f
WuvE5+S/c672XrKvvSuQFCv3IYGMoGkgovg9T6LYq4xvSK4PPBeeu4+E/FaiHslB
IH3f9jZST7D9T2no20Xx4tGFm2IueF4tfKUZk0MdAezCZIOoQsXNP6oK21OAIrdi
rgSJfEQlyKmxgi/CwUoTFkblgxAuRWp/XftTaeYJFX4Glx60YlKhY2xDfzueMK0h
iIPPq4xBD7/ubVMtFoyHq1PMEaAhQJCttP9uIXtdXrFv3m0nC5Qt08gIUMwRYTn/
wzPedHPP5da4GWby/ZvB02CL0z0kbUA2Tc20jPOsPA2jpqyMNlk5mdZ9e3nsqIgw
urDyYEV7hxLN0jJ+tKcEYXnqzMpWrqTmbNehz9SlyBwq/9zoDBaOBQpF1DCR4AHc
Z5YGwLMHGdu9B1yK2Na+KU07XJLvI+x2prsslu44cDJyRHHnZ3JbU2R8POmLSvr7
JvTZugPw4EZf3dVEnPjkGKogS3zo7rUDz975nYt6zAokHo5kZTU3RjhM2IuOvlIJ
rnAaz+Ym0/VO28tROzossdhOJyJR7YQ1ng1Pn8D3zyguhzKtzwxs31/oFkUx6ixk
WHAcD88kauwVlx5J1pPoEkDfQ8f8bcPJo9akGDLGi1B/9umCLpgdWINYIIGqxoOG
ywZa6qgsacKTuFGbGP4OvsRPD+peJw5bH8tY77BAekuW7tS5doO3ShuOm5L2E5q3
LGwqAtwtRacunA7yCIAF+D1StaA79AldF9lUYFqc3+gsADsqLLIcq0Wv14g8dPiA
1wqYSSeljiprLRg+ie0JIspXCn4ZdmiiKqK4Bgc7Qkau69Gb0Dxr8su31Dph1rdY
cyIMZDuoedkeGX/aVDTCDy2MCQla0QNU7OflW0c0RwEELW2HgKVQVDUjBe8EfiVz
0tmyOUKMu1qWyFqtAR4QI8qsd+0NwtUlcCaZLjlWbk8Z6ECcc9sksZwZc2yXKY14
V2qv19B0y/oOgMEePam7zmEUatcl+tSK5XDh21pf7M6LsEvcIJFMafcHw4Xf3p3o
EIsmADVs7SaBPgdxZxLBUO2eI+GZfDzi0hwHh2+Wauk6vf8T9Or4YFsMUrFfNabf
SpRdvJcBCS+hLqhDp9Nk2lGLYh4GT1flvZo+br7LxoAqmGhWNv0l+KsZ3V8Hl6L4
6FUy0ynXUQ1gLOJ6EOFSbaLh+qG1BKO+8PpD+dq/82/FgjLgXKMYDnscdtlbz/BG
TNCicIw4ZYS78BN+o+h25qP6S8Mv6kNbaUkNcmp97AJiG77RAERINvkR5S+cNstR
Z0OvXiEisHQnDzK3OcAActbDMfX0iei1RAu7af7oI5mZcgc9z8HgrXLVGpOyIzCP
6QeC5EOOPPrOUIaLaftF5Z8Bxt9Z0SPCmlYvUEa/PIPjrGqR5a7BLMVgSX2I4x9O
7PMT1m9lVe8o0Ii7eZnNhJz0r7d0dq8tWQ+AOgs41xDpklydAgu1PoPjmRlQz5uM
6a8WcgIn9KvvzkgNJqFQEsbRSLtlmqKCdYuvlEO7WvHIidpJSIRTyN+GtzfIbyNC
LiDDNi9GwoGUJi2h3N46Zr/VMTk5EIpjce0laug2kn+2xZxlSHK/N987OLlzXFAO
38txNW6jKVWKyf+WjC0PR92IwKAjuX1niRo9tqDHbr4/wlWlwo3yF4JLUQb2oqhM
tgpotcK+l+Vuc41n3lm25Rd0JSH0+p6OyWZNAZeOFJ8aCYaNgReHdTKZOSRZqcb7
Tb2spyajjet5+n6TnqaffeoKfD5vXOHahtFNUlgN35bnHsT51dAbWGi5Q6WkBjNH
nohidwrsAa+jSVDx28rgI2XpYoCGToS4HEuA3obTce9gyceSpZtjfvmGRHK0ZCsj
UhmoJiwtOzMdVMMOvOlur+p1CMSkZPiOfmC2aZPFWYtShNQWyNITBeK6Lk11pker
bkP9s6a4PWerJ0AlJ2AM5fmaRZxqlOyXj8E4vwRnFxdWe8pQte/kFuoRQq5wov1w
6UD0IMF40OHG+wuxGbnvvkQ1Zzb8kWbQYGuTm++yO2ZllLiCuyILLB7vxZQEIsO/
WkkQXL5N1/gWwYvNIM8X2A/9JQ5o6Jeq9ePfrho02Ond3I3vAO8SPD4jqCGlZESL
2t5p8FX16NmsyHfcwjTHkaCesNjpI+iOMge5d2TdSuFTOCrOsurimqRXujFtPT/F
FnrQ0/dG4TKBTf+EJNvhT9e3UYMf+AMBhPWKxdGtwtDTm+00902cSVAzfkpBbZUD
+OIDpJthJPlXpQ7CDoyWXP5vh8vRsXAefvqH3HFgvppUW2f8j4fzSAYo6p4KgH7V
kM1Ivrf0Uw94fDLBbZgNRrW//3/jwn2l3hJBiTXiSipi97dXaEeGglCTCJkkmaJt
IjR10sTX4Js8kyLlKYX7S8eDxDs+vd1tSKbZ7FDeb04Cw56iLudiE5K2mfknN9yw
0CLfJJWeMstK6/zFIKqqTNcS/U/suw+8k1Sae7YoYavX5eCi9A3mq3Z7SFY1Xnzo
4mUFMmrX6GyjseHSUnj2VXASHUf0avfU9QCmaeTFK5vkwcO7uIquDSBN6CoNPmKC
PMtvoj3SA8P1AZhFq0dBxk+qHWvfH9hH9lr4HZtjWAhwXtJP27CPOvlbgD6JWRL2
Le4S4DFeHSxa01asjMRAro+ZEYBthnBSk637HzrDOuyMppeGsyRkZaxzyYH4XlJr
+nZUdm9lfWTyKes3BFkFvTGApb3eH+Fa9c+y4q/Z6JMLy/oh8p6zO3jdlRkRYqR5
im8FXPJTczuoq9oF7h4EMTCs+U1PALBnZxuwdBA5ta6898DR9e6SSdlvn+Qac3xL
847o21SgW9KGhfNGwyHgCMagxnCxBPdHM7Esj5qNstfUSDMQJoro+JR5SASM8coR
NimXKLqYnSWQaGSS2rBJN+XcaUYtdNOORPg/IpdxuzY8T2GD0O6yLVr9Y7CNCN7I
ccL5q01hmgMc2rUoR0Pa2i4QikHiE+Ydi9wGkneyIaQ1ksupgZlWtnTeRswF/Y+T
LHrr0Dzpj5PjT/o24jslFfog8sG2aBBLKApAHzw+EvqIpCz4EyJ3GgHxxSfGHjb2
FEGTTbp+2G/fGmIxzVDcI/TxVg/sbcVctD8Y+qTPOVb3Kkp+6bFzTSCWZUloCQhK
u0wKbmTosUQRLQxp5M+1Q4wV/1YTcfqAzWq32Nc1UpYwJpqzLHfcDVKTmZxwHeqE
P9EHeldfSWxE+pDyetsjwfF+7kbQ4fN7+34TneigRhZw5lGBuOW46Iur5w1b5otl
3JDbbI6ePokLH3B39fEwNGDmfIJT6PRs4NNpf2Ag+LmIdbroWISlSMXhdMA2LDls
piZrd2DyIgGcA7QOyu4ipQ7ssUVunrPmu8C0hxHKdJJNVZheGiaCVbc0HtJT/zIs
CAHiTrSCYA41a5mmRhtg2dBiPsuFZztjZLaXEb8EpuLNmXco0zBQdrVy74QJWnPD
XYO+5/CTXV8JiMK+G5+juhkT640jGfzhBWEQtpnaMy8+idY9Oj4yVjVf1g+yp9Fa
t95Gue0cYpjXTwv2Mu5w+QQfKFSDWQv5JycRh9jfyWmkXUJJy/F5XBZlXe/C+BoO
i1gz4x/nRCYpwYGX6h7Q3ed/YmkTUkdM0m1H4oGADqsabFfm9ZulBamE9LBaWOEO
JsZU5Lq9qFQWYaTlH54GFD/Q7xBasIxYLb9XBizDhowjleMm7LknSTsl/GblskPc
Hsc25j8nJZIBtu/7cWyBjaoeIh7uswdkbFg5yWkbZ6iCkenLCK1aF3wOXjpjkZ6H
kNcKYWN6yM1ZRB/C0+FguEvCt0ZwJDmzmim2rKTuwgsGJRrPLw0ThPZbbpejAXgB
BRAqSgqeEioKQbVJHjcrkr5igYs/iAKFaweL+5e2QB5h7rc/N4ASp3RQaQ7R0RE5
RjrswGG7vGtWcFuR+/025clZ7PJKhWD2h14Z97MHeKrx4gkTCNv7s+lVra2WqOKU
gEDijRvx4KqalLCkh51XPsXVWvEcOlxYRUL+DrUIFKg8T5zYKpqbgtjGb3rSe6CN
60WoZBvXBBlCwOeWhyw1ae85N5gf0Xz6FSOpwGFkekizb/4qzY7AP7cd0PDngDm4
uiEzGzpp7RoieJ6gMiG+pZmWLQJlhvf1PjuDdGndgqibqbGm0pE1FaI1v5oybWWe
pAbMURBYl/zZepGn5nJfsOYePZtJFW0lkqQzoVXjenJbhoBzU3RGBV1V9YeKc9Wv
OeQXrMGjggFt1EZb5euMiyRn3qk1P1BLrj5uffXUApd6Ix902UL8ktVMe9rYIj6Y
hZc0Sj6ya7WTOgS+hRimzpKKVX/H4p3QouxClOdhy/mBD5IuLT+7t498rkg0kHdh
J73GXm4aGXlYRWC1F0R7s06oCUcZyJzQqc/uo6SNcBxYrZ9ijYvog2kTcMPrDinl
EN63S+FVaMIxyRzWICTtABNA2Qds8SCtSVrCoOhfypVOMlAjnTzFTOqfXUy+RGi9
Gr/NyeHgGsCD3GMMvlxyiKXMfDCq6LJIRZ9kHykvk2f/pgeg/8V1CUEKhlr6leLp
z5GDns4nhiAGs7VRl14Jjdi7ayaS/YMafZoLFN08AKq6AJwGLvsr2x2wc+nE8MR1
pzBPp8Sy/wOFLyNRCjIBfsYLnGheRi3UTjD3OB+WhTReKLiNTElfwaQQBRwGtnnW
xMKpYPBEsw08wlOShqVSCiiFYcy5a8fKcACx7dEUZzZZIwxrcl0Tp5CnCgXTJW2N
8IoqIJQH3MsaSYuaekY/Ej/tTSfHTUiD22mpfphRIgmINJ1jHo0qMhxKZBUk/l12
aJ70PGC4281/o3Xx6kl/zEQdbueca3B+bXxbjCNLrBQZc5zp/1eTwdY60IwfhRy4
3/Qsx/lvqH0XAgo05yqlp77mLpmmgzsP8NvEMRnlcYq1izhhTWaLbJ4GZ19bKWUc
mYgXkHrd23Qd6Qbw+06bnPvtv3JPpAZ09petUFN79NjeHfhVMIcyjB3ni4E4liHj
MtwvlzG0JFky/SZxA28fTjvcRcxpVlC+QYKmun2TokFh+UUel/mBLuYQEBmII1v1
Skr2Nt7xDt0NcBRv6+ZLngs4gK82vK9rIkNGqQdwp/GTzARlvF8kk1pVHwodRrs5
UsMQvXXYhsoC6Pqwj1o2+uXJLXmj5mLMNYMz9mdZK9PCraWZXIUkWaa6qVjFGDzt
5AMjl2dCjZmqnrx3Rgubf0VEsfiEXF6deI6ZEJ8kfaNWDzjO2//cqQOj/6G0v8bS
ku/XV7ZEycnBzUESvJd4Chdn32TwNXsIDUqBnHbE8/JO+2UnHw6Q+JSAWjs2s112
Z+s9hzHv+tSf2iDSXFQwRdjX2GJ6OLYeykHqrveNdJsgek4H1gszbXYnI0tyhIJb
Gv1lqwBI0o+G6vc62KdlDpwMlkAT2yne2OB3bcENYHMvFyyLsodwhCu6sOjy9D2h
Q4MvbyZ2G6eN69cV2rv+oT8OlsWCtJwxLYwaKM8MDALwGQs5OU+t0qVKobcftmYY
lbTsFRs9XwdzkBYkkP4Bs40o1CtQaa9gOgjldmChNCpltOta3jnweAWCT57wjMuk
2Iy/9MkbnVNmxhiM8ybxtg1HRgT2P8PpWlycMC01m2cjxprvhBYvHBfHt9uWRJcI
FNGCi9IWswihTiqtlvafy8Xo3OP8zS9tEmgAqtHWDC5g2eihsQkGghWzqZNEBvaU
Q/2ZiXG0TCts3d9/PgWRzNsy1hxrtstCJ94D0KcDtmxF1LkS3hWl4U9bSmKsRInf
aLxCUMxDRSLBM3CZOLz8xxJ/lFahcf092fTbnr2QjvltUBUlhvyWT52ZAfwoLJKF
eYduf+XW79C7Mul4eUKu/uZjj3pq14ihfR9v67sWx2zv4EgBSQVvsWuyQnEwypZD
0Km0zuu/gCUHOQ70SLNXM8ei9ll2fbjj9LK3Wj0bwjTJCIRZ2NYxcfO19q84cNEE
fHJe3sXmUAiQ0eRjq1JvuUPypKVf2bqmXGRHedWqWnyL/JNlym2wB2wCieUAbeJO
savL9V9BzQxsGLdNbiuDJfQaft+4EmdHN+sOc0DlcIX9KjQYZEAVgGIup/HQ8T/t
VjLdPqaVj8at8S7y8sKYuKLzvsJdhET3JrMAzcwH2Ets/HvysM3nUTWi3ozFwnu+
GU2VBI4pkG4E+Cw0+V6zWiHbsPWafE3U9iaLmZ515YzNRUsUvjDJZTG7PtsCqvgD
eODZtUOsqbUT/5G4O6+fVRRiAW7+Xdo8oowvgoXPlJB6sQb8cwfZ1MJzaos5qUC/
YMRjK2S6FUVflNngf+6RRqj5c2nywxFtczgjlVtrGz0lPQgcZnj3VqJXNfAdlBSI
1TpPA4bKlWjgL7RvSenCr7XVE0NiXe2kKhm/rpQz6/qmm4HEaA39g5uywemmBl6u
Z+RCZdZ93yo4ZSY9ajP4rkpom/cV7PcyYvSH1sExv8vrs7tD6TAyTgzZwVBJpodM
K/pSNN9156+I/uNzynH2FES+kBmRrsOCXqKJinpJCosHn0WMLgXomIVo8sM83jQs
UACKKw3pfbWOiPjkc6/mINdZHUybYBXLMy2HY1aUxXDO4wZE/mlMZw0j+XSKDFxt
iSCiPsrkXGewRaHL+nioJYUqbDxoaDXshI4wOkhIaibNHgjNtxJc/ieM8B4wgGlD
jzHS/oL+Pi1tukTvU2P5AG5HKUW3Tl6ui0yHJ3rpaeBZmQg9nGkV/0z02MEeqPVw
4j/Zb0afnGZH9xJ4Qawj2bBIAEWfct21ob0JRp/YFGFLN8jIT8stFbc8ZC1mupNN
6TwAxi4shLTidWN7ZWExwgzFVdZAL1CCbyP20EkAUFwYnQJ5WEyfBepSH7nPtwJr
PNZsEe0yJ5usevMzSXJJGsyGU082rdxkkY3J++giFhBRzQ8U50vyxUWoNelvZzuJ
sPiN882VSFzYooApVQECfRQ1ircY1wtJ3chCvUwTyqfELur7NYb3x9rIuKnQtW6k
lf1o+sH7zX/DqMT6Nm2ZBS2DjEFq3GoWzJ3AnqgXmmTPuwzlR1dz3nwIJ8BxyV/s
Od67haga1BD7wRwP/KlsqCoy6cdhYfcs/SyC6+JT5TDwS0cIdepZZKeylJxuVEDz
bh06/cZSiZHR99rD5kEKmzsBFV/COGl4yknZaHMyWHACzo+VljdbN9drjG3b/nQO
bVoDeDE08mI4O89vfTj1yVJSfOPTAXi+w3FdGUb80IDMse/BeJMS1SexkeKlDbPY
sr0tQOL5tnGrwCLvq0fe3zhcjMb26fhIiTiGdVYwFCPq+RxNYW5XzJlH+NSafOrT
Zc2SgQsYr+ohjTjSz/gfv0ZwslC5aBDdY7sg9j/fjCInJhnB64h1renLfnWwl3G6
8g1M5IMrc1WdvbBjtnCOXn3M38Gz33fw3vUkipzSn9A76sFDwiWZON8MTxTODY7S
ND65HdwtEqNfmeqwAar83SOPkM0iEfW3M3CgQbAa3uTx10mGufmDHVl/2HHc1PkX
LbuH3BZ8JrL0MU5vHWZtvaDK4kr5LfWjU0wG3AJSfcfMLhmdSw5dzdRPpZidEFdV
JaEjHQ52Cyy+bma4yeD9JklIjkrUITiZK+4esvphcFgOd6crgWN072E8T4tMBNaQ
pxHiQiMg+GEDXd29gawavH2BulWts91wItbXmUW6KgwwH36vSdZPfa7vVh2HC7lE
cIQ5UJrKy08IIN1yQLq/gQXb3wGBYL1BGt+HFMMzM0sTA732sFaWjF75pqdTwWSg
KQ2Yrg5DqyX4vHGGDRy8JVVIc9b3hAfoCeq29WRZ/MZ5ZlmGb22PYAKkboJoyHRs
fYU6i4hAOvb+8crCeBUrjGPaXVdhbnmMuJTGNVDcDD8f7tzolIK0OVXaP9vBMCdu
Vh49JUAkxPM8kG2ckQR+I+f2KSsxcqLR3KhFdBultnxQtEaGZVSs1y2/JpT9Tz4P
B0f6d7L8mrdT7HN9/81cUVe9hJFeb0EybviSbs0me7RC6lLjXvD7rpR8MYZBwbyd
IEKhM0JxFHEKea8c/iObxlBIVk6BOPLeeXOOOq0NI4ZfbQWFrP+OHtsPAqc9wp1i
MrrvPv1se2rsYtt3dYrKcGS7b/2NVF/IWPmOyual3jhxuxDeWrWjVxbEv1pQ4MiI
3QdMRWPtDCyVcWEUuUHW0vIsTIgCyYUdvilP7osu0RHNzG/NRxU2WZSi+f1qT6nX
2qCNmULdIgEcd3cBp304HtaPYMqgETBWox1J9cCJvnZBwjip1mYDLYik5SZ4DXWx
lI6nxurg1tu0l42FsL0pkkD3ps6J791il6TbVoaIRAbuDobOua3FRI5pTtMB3aX6
R+s/lP5dAhKCDzn0U2SIFs6QyGtzsudug/TbLNrXNZrHGUBGufVoV9wWc7jPeP4a
e2Px4oOHcz6avuyYvyQZDIT76jwGvDHsX8N/xaQXVN1Tvv7koQ7l4ZyI7RSC5wCB
STAOlChaqeY/y3HgbqjGxReJPwv9+5VOZZt6oOXxowy4DnNXQbA72WpJrXqqvgaX
F2QV7SqaFByN0Tzq0aFI0KlXNFdFOuTHXe8ycMnmQgGXzsVJoDk37I1/aotODKna
D3j8RbzxcZsprGO+5GUV/5ppCpUi08pBc2foEfeDlRfUawVO/vkDt1yormd+k6Fv
kx6oX7VMLFxuQ1qmcfVtH3Q8wTv7pKYPvOX4D0ujNVezKMN9aLTNfqthXF7BL9aR
Y0F3acRU81SHAd/cwTEz1P2qk9w3Gh5/xpEiP673VJIYVvId2sYWXWMrjpyXC2Dj
G3nSMeqSbnKOW5UgiW7dCIT79Zp4DyT+xb4dBVDl3gNgg3VOdmQK5dWWlxe3M+qr
GyeO19oecETycj3g5a0SDIxXnlhhyLgWRADnyfCTAd42302ehIiobGsKLIvgffLS
GDDcnReXXTJEMuG87K/ea50w6KoTUTIDcuKRFMUIaCDoOu2fpd9UtRPh2uxJXpVp
2XSHHvYnDnB3zWG0j74MYTXwiyJpbP8ekXJeYr+OU390vecZ+zeGp3RcpQpjzkLJ
Dc4EOQfH3pJMmjmFOhMvUoDTnUv7sKIyk6ZFcbXUQ/JgicPxrQx1TZRefWGrVKpX
/y4nSnghWTGOdn9UcC1NZCRGGeBl5Fa6KADqD58BuLvQxguYGuC0kb8cHjaDNBTC
ncUjcOfIFWjNOIYY/Zdu2kKGG3QxScVAm7CwoBvAedz17ZGAe/F78n41Sqg+5w27
tPpBy82UZXyFpF5Ef5MgIjTmtclp2FsMqE/yPoc5oHkJxSWx6CcdmeIZcquVTLGU
iWlDh6N15aBHrO8IumWHHeINlWmZYCzolsBdY520c/QuHssdJILQTVzkHCg4ei3v
EfMSz3jv9q5GCHH2SKQKsX4QA8WRIhPIAOzlhixP59cB1XGak+vR4VFKA+cISXWL
0OyxFGl7vj6/eUGe6S8ZWKNnb4CCAn12z/MjTcq7Petf6t2cEMbSqvRdz70xP8pq
Li/lRbk/wfQWdx+J08XgCS2vJ0uL/pzO1pG1M6Un2d+2Odsa1JKneFlMpaZRsdvi
eoaYpMiQJwH7ddtetsmaDm19/K1tjvCv/psbkBZ/21QSVfj8q4QoRrty2mAP+q1q
Ze9oSYmwh6q5GLVVuPq/d3WxH+PLxeaabIRmAgAs75TwcjYqX4fgsehB2EZj/S+i
yDw0rmtODjTacVKR9OInEdiKg2FrpIL47gGvHaL/AzlkkWHLXycRIMNq2/tAP/e7
NgjnSlaDwt2azV0zMvkNDfSsayHg6eR5egV4GAk9ZHxFZHI2Af8UsfzBpu9tRMo7
HFhTv55XebcihbwZnPIY4Pvo9gmeTMB79S/KjaWUiLa4zMkMbVZ/GefuRmdjq+Gm
gFWyyGDTAJCfYe46XHi4zpwvyvqSC9dK/qqbzbLBV4oF2u796F+KW9SbhPB6BXae
YrmzkCNPaLUiZo+eZWTrmvDLRGCxq+5XxLAYhRvkh+xS9354AHWVPCvGBoUurDEi
5A6ISxUF3fbJEGtzczWGTjHi5B6NTMGeDdzkmLXOsiZ2GqdLFU9RXQ8G8R1DC45s
YsMiKYkLgurfTLiqi8Lz+1MQentXZDko/GTUzw8AY/88U1W5vF0CSuY5cPRo4tBz
T6fmiFhmAoObx09k3r8af59lalTR2GcWPnimCtgOIVhcMQIbZ/ZC2+c/ejWZ8xsX
b/He8yieCakrhAvBiKBPdj8Xern5sQQFKr1RxBp5cpbphrtlgdbg70cr2WlemkKt
KrL9cxiLNk1aOrMQPmjg4LYG+AeOGDhMBoDg19GcNyYMadcxq4sW3redyOspv0gc
vVNTT123A0Hczn4+U3TIsDgNfYy42NrEs8gCixTFsZAR4XwTa7/J6GyJeo0qU1jf
tAM3tXd2qYnupYR3/dBAge/rP4Twq52q8BMNar/tbw8E9DZMz749fmVk4kgpWudR
3hCDYEUHNzNoX1UwMexvFdAatC6GaxwZ1CP3idMToORb7N8CGO1Ew2iV0t/Hf4J9
gFkcHtMjsZzs4C6r88oEqO8I/nZFOsOTGoLpQxCEVAIs7tPXzDQECxW/iT2O2Jmn
54s0jMRVf8OyQMINo6VOTrNV72I0N746aPuO3g03ZURddbT3AmIb9NuKDPmJKxIG
u0CfnwFXLv58dcv7bud5/8BlFF4NuBHdQ8koqODMQJBoyXYMSek3UZiLDK0NWG5Z
XFcsyhlmcc4LUa1Ug5ZcvinPE4XN/TrOaemb7fjQz6hv+j8BYTjEgb13BkLKVJV0
fQC1HvPwg6H3NGF5MtkkICCOAH0aLgvCBqiXNsW9sN/SLZNfaqwipMQ0UZAMFCTq
6vEEttMI0wPAlgvYwMhdpX8oi67Fg/qA9qH5MLQeLiNVMfOgY47P1JuXCcga+x/e
9bATY43btypsSSr3bK04MxQHmhIqP1JKm5dVhrRBg61cS7+IU6y4FKnOcqw4Nz4p
Sgapbm68pnI9TvfIWgfFgz15ZbExs94n+7cUKvOSS0rmAb4uG2I2sBgAvFrkRrs7
cu/VcaC3pJsE6PzA44UalYlyf8tzqvWMzx90DrmGxjw5cwKqNU5i82Ar09lKgcKe
l4XuIBgKk7nYzH57xo7BpuWaEROmai9lCgCLyFE0dYkSY6tYn7Et+MpxBfHmv7p5
kI146CHuh8C1w1Le6WMaimZFNQR1qP1vj4p8oUefxVByMU/RAEGfrKjBYOqa7Bc4
wdFDeGrUAqXfOhimjkXCFgnSizEnCn8HYgF5iGJDfEz2J1JLT2nfImG5zxbaUGZg
CLHEQ7Ec5YbBZyTRcSyLylEtTPKW5/MJ3yoMJqCcNaQZp8n0HvvHxIhsl2Q7xYj9
qJ4wu85S0mb8rtF0PeiVvJc5ikrUuKQkczjIbyJdYgI/BEyRtM4Mx8a5ty8xUOJc
/FWAfkDla8fQVWqxHypkG6PrrIZy/oXAZKfeXLsh3v7gFs+bAbGPGY7EiVAUyIPv
FE+l4H3edq/w43hDQ6pdtLK8tJVAOE05UAZzSX8yXGnuZNsYpAPoGj7UMcM1JQkZ
/oZmCkBejgyPkKsWX6pRj9mIVt7zY+eU8DMxtJTWQ8Y8sURYpSAMSXvSOwyDwXxT
KfKUd/lUgW9rzbzwhHUfQ9vBSgTdpytZDa28wkX0VmqDsTe02VVSFPSJeVEfbvhW
xFrf1djAKHocOeiBURbMBJCfPON67b8MArr2HdIuaD3sWono4YsgKJyK/7gykBH2
StVZuM240s+5EWc372GqA5CXzt6hWxY8iuEkmowXWjYVBFy3AmZMwdhzScmprx+j
GnVq6yAMJQMv//iziRBj6Bof5FL6rcS4ea7SYNjvdaeTSNU0qcU0A1UD6lPpET7J
9QvFgEiukS6qJRQ3AtIMftj2B4Joyga+1Ig7Xyj1GVLzKK2EePW6O3S2peTPG3FX
hJC0f5anI433yz9Sx30XdlT7dHVUAYr6D/qZCM9iBSG7NGX+LioilW7WitHbaIsO
UVhQH9BTMN9GJC14ltwpHf+rXAicJemVzOPtUJx2ymf36oyqb+Gt+t0Qj3A1Ezdn
yO9cw6wkuifpXOXIq12CXIz0b1Du1CeidKFomUk7yKSRHpya7yiiGn2f3dLU2ryQ
Fr/cReJRUN27PRkZ0SiHrsklAFUelHn2+oYMdt1ErEsBDQy9SeJ7hO8OdDzcbNAS
cuwAvss9Qmbd/slky1KQLDTRpqsLgfS0bMrQf1U5jO2ENMiXg4TZ32EqzUZ1D6we
PsvGMIgoDCy127CP5EnaZRVWvdv9TNRABDzuTQibwnEVY5E+MMIb9kD+yom0xVG/
iWaGARsFRrK0jbYfY8pBglRRfWpmAk1Ys3RIZcOp/ulsCbrDyMUT55Tn3SR92H4R
7Z3BZxNiCQnrD0uHAv6kcAt9HmKGr+2Z8qnMjWK5ZCJW95x13hmpe5RhpWJuYwEx
eG+btCUpm71s4Ly6/CoJQeFOopHww+sNEoGFQa5UCyqqt40obzSQ1yEmOmQlKQ7t
Lf8ku+oa9KpB3GC1UacYDdkyPkLoik6yOqyNphsKVWvtkaJ55sRam0CdmsP8G/B+
PxiKKG5JKsYGHN3nPVWH4GYCmIcFIJjoSLnA83aj2CPrBn1kQkK+6mgKr83jptw1
5luMgEWtXSQyneXDz6Te+g/OZlN0wZFE7/yjeJFmlb0DaImGw+ikZoeKgMAc3IC4
mvM4L471hw0vF+4wxRkxqJONDHRuYYIRej4gVb+/luqBk1kFJbIXE2fTfGTyvMQb
lsffDQ/euNr9tsVOCmaL0O6glOtWKuVp5aQvKGL7qQhzBBaOJLIb4QM6rODSNZq1
BV+XHqEC3HcaIE2xNnYnVzU5+6Me2NMHV170BsQrzT9TG3TZSztrg/fuNjet+8BM
cVSTnRu6WDx7JP+G/s4jyXZ+eA7k3FI4jyb75I5dEv9syJKTYa01BLOAwC33i3ZW
k8Phgvt6m+ngbKPvkxbxJpMkF9sEAzcwLjbRxWFR/mJdbgff5rn+hkeeMegOXxY5
umhUWE3J5O5vOVUeIIFyxJdVUaGGUQAbXKhOOECex828rZ9fRT+/R4EJ7McR8P/8
Fv/pv8Yt+5MUKbjhnN1mSDsG1Qhpjo268lcTK3JvyQFHEQe3utZ4JLUH8tKeTW+A
vFCr0q2iZgrTLx5LONPwr6rwsKQSSIzNk7bzp6JMVaCmRoTzOxLhPgzGTT2vGagz
3bKINypGfZz9/9ZlDSBx7ELdDsBf19VbU7mDJqj/DAllL9uXaHHDfRpWqolCiaot
KD1nxo1OYAxIYdVL418YsUekSb+caX4ySZkT2rLEv/99WKgxo76T0n7HYhVP1skV
hW+3bt6pjymkmY/i3ZFdEetUW/VUAE+S6+LnVPQoxfeVy6biuI0hA/JHTRadpPsZ
TV2at1P+4Lfabui6BJ4IqIDHihBdP5X6KTcOY6n5sicCM+lv7+loOx0FV/kPLdX/
wbEkmXFj6bIJY1IUqoXkNdh3DyA5YVjL16re0HUrCBs7d6S1W8xTOXYK4rOfpds0
PaR308OC8JDeZdudBSqiMO4V0UAKdkykHQXJesg19a5gDQwNG98UWja+zqrHvwWo
SrS5QT0LFQaA4Pm6MHvOXyAuXnkDqsrvaLubuxAwO4qUR+bVasxCcnp4qL7c/8EX
Y4ji7FbVxdMjdvy4bJGMAAJSP369ilrx2crKbXm5FpPOxQpjCL3Mc+m3q3kjGAdi
9tu9NaDAm8TA/vBM2q47poJfJp8FlRADBzfG04P3vFmv1zve5kMoiTJuENBa/Tr0
aCN6pfUurDZS9Fl1JU44MP8DDdyuXF7x7xdKZfEk1Q5GOw4To97KtFla0vehO9QR
N+cvuZuoDp2FsEOSjRB6kSf4FEN6AyAOmnR4nTw0+VzFjzVlazaYOdCermrA+09u
LAfYg7WiU7VLka11mSi207k6Ywwsf0x+SIRr25rm8E46CpyiK4fmhez18OVtun1s
m01xMupquQF3UqFoo/xH7SpzE1BvRrAjjfv8TRLOiX7aqf36ry/gOt4SL6tbChB1
XYJt+xBS8nz9q4dfIYNUZmermRkjIJ+6IMec87b7V1AXIp5HhL+sBcjo3FWh4N8J
g7ZegETWL4UV2J+cuLUoQPqPk9ni+UmrXX1FzP0UaKCxBGAbQzqmaWVNxCzeokGx
njYY3eoU8A0OZdaGExx9iPaIKSjkAO7jqXrno4IAj1c26NFqdm1wlzlmB2STFYBY
Y8lHJypwebLv5sroCsQL7nqqNyy+TRsIdkLu2CzbEhC0v+RFN19nmdgfhQld2igk
8aLujM4SaRO4FPnDFdegS/QixHq7uJQayqW2WQw24wcGOXuLWWT0PbYvAOYhybhZ
Gf+jJD61Y4kvvYw5DP3T1dfObhfWqejBDXyrY4JCszZWj9Z/waBDCIpWIYRkfXCN
W/DJFt2FoD4afD4VowhfvOpQJS7TX4P9J8tuo6SRE8j7bl4oSWzuvH5fnJe+8ixd
K3oEH9qzaCwoXnG/X0AUiP+dSPqeTpban43QYAkx98gz3nWZjmfrksrexrDVi5I8
H836TW3xITbMrK7Qrh7GRRz5S4nRNj9CX4CYWFUhYVdSjGKg80cmTcphClesLYxk
fG5IMclsAtat0BefTHc0RNOfeuHgdzg2tv/QgjS5dqqk+U+zgPzFk0VSD8qjw4vR
iiGR+e6qD5MT8PvtZIRixVYx6aCPXrlgV+HafUcwmHa/w7JLJpv7/03fuBTEkCRj
3of32GRNUF9lo7JTJL9btDqyYB7h0eXODIPVTcPPeyh/Qg+nHhcbe4KdG2wASlHV
fAXrR01SNbpphm3b406dYap8Abgq31Bl6MHueTlo2Fcq0CRDubkeTL+mb+R9bTfK
bfUUJDAf3grWClCFQ2aI9fvYaNWT2F5XP7hJdMBkRneI1ekOM9pCXHBNvx1XfupQ
3a6uWhJPc5tAfEi2HPcE2ZP0rz5GXKDXBTAJPLLumld2RbJSnhX5oSK3wU+6JPtl
lwSyrW7OEKs02eX++ORvS1hnIK5Bik3eX+RZzrNzmgwXSF//ABBvsMefwK6LiK9+
JbqXKf4S+cM7Xp4ZxDDeWZICv2a0OE9cV0iZnRzg+EhpnOiwjK815r8sTkslqhJ2
sfXg8+Le/zgH2x+TvWc0J8wGKDR187sR+9MorWgFjwi4UwcRpQ3aaSR4Gd1mxBiB
K8oJzI2Q6k38kZgk7typid5ZAYVZ86rq+PObtAVhZXO/TdIHJDn6kh01JrvzdoB1
v/yYS+OtqcuOjJWc4FuSUI7Cpe6KFwg6Ke5pR4skP39geNOjl950Q1ae0TuA6XkW
ciWQQo0WAh2F5H5XfhC/UG7+EAt3JGJwTZN0cbdtD55gxWqqD8oq7bUyavagmb7m
NuQwH7mO5ahZfpaPk06ZajX9Y5/aJ7inD4MBWNE14x/1WSKTrj+z+gqoWDFhOg0J
KNoOqQEtbIWTaPLBA6eZkEcPa/bPC8qIYvYyVGZDM6o4sKC9HVT92Z5B1jA2kGLW
f0wc0QdLbbWNLQJUg2rfH0OT7X+kexwrNrGVq2DdlYBoiRT0yHwmuz0F/v55dUj9
Ayrl6YdavJwOhSaZ/InJboSs8PJA+upr6W2BL+0HsjRhu9qD20fP58x6GrXlRHwl
aGiLUo2kx5evzBh31c2xNwjl8dfkZHq+op3un6IhVKPdlG+9fM8kV6CqtGnm11G+
Oj1Qq03eDoYSntTL0M5Z/9xNTITvrIWrejiED7COmYQndDgWxM1G4v01tc1RfTlC
4ZZuOnXIqNpgOVwRvsAgdHY12Ha2lWTAQHeCFtvKDVVFY7XO5Qaoy+7x8rZww4xr
PWIAloWnX/h7PItzPFG2AbKf7KsCBVoi4jC1ByRFL3BmWIOKvJ5sP8c41MzIWvA1
XBI+yXIxTrGqttUbg64HiwqORdzq1fSbLZU3fOSCvTTU1goUMiE77ySfRFLD/R3/
z5AiL2piNaHUxHUjQTzy3JK6QdG3FEHL5mdncrFbrdoFSRZvAlY89OanUZNXG124
FoOZfhF7/VMZbaha4fvZwcGZ/RIuK+gWCsVVuj5yzEK1mJ+mKkbfvu0F33nJQUTj
CsahyO9c4ldx9mSKsh8izkoN4wdNRKaOzMdo0KSsKE6bF8AIZ3bqxhZWFVrLui85
CRCgrAbgu+fBhhF0TZxElMelWwUWJvQa9lS9ngMErtojz8qkHKf3NOMFhBKY3EJw
Bzva+IhehqCc7w5n+5arGlXkTM6iVVMR1ki+hva+sFy0exPZJ+195dbG+I8vCvz4
+xs7xX7UlcyLEXMLELood7O/kVeMgxaf+vai0gtmKn9kM4n6bXMRyTEDbLQKk62U
5PM0X0AcnpUfYcegbV6RjnCEHgMYnuQqy/YZFGDmJq5Q7g1pHuMLenBDx1ILhppx
HSfmYmePcVmrL2n0+HpQ4IL3+FkwFl8Ptz6FuH40D4Cs4vAd1Kd2W4XRC28bqxwt
K5tcPfaSZxwwzZuQFjIWJgYlZoTloUUreSWRxDTRqDb+kxDiVoulZtHMr9NqjSBH
cSUkYUkGtB80VZ5ubE1VPA4qrEoMwy+6T3SrZ/2NNPpAs/BtFoiS1DDb3sy6VyDs
rrHIAK9DSBmmHehi+Xx1piMNQ/kGa2CJsSVS9Eb3ykkyfnljG8MpiZn1AvuqEchJ
cYaL77hoetT3RapxP7434w9G4IuOfphoseeS6e3boFiUZVFv4OWI5NNqN0SzL7rA
CNIuKwtPdFltjHWcL4UqciKSZTs+WkyG/L8sVaoY6EhZFf6P+r3eqzeELQKCg6nH
X9jmBvZV+fda2Tspon6q2hN6bkEtjgFqI6nRWYR5dK3X6MwVjS+C83ZYaHHo5oe0
i6EnZNqppma3inH7kD6sXse9LMnw+Lq2+6rQq+q/G3st8G3ab9nBbajVxtB41WeX
0bn2n7JIHwky93AcOHrXs/GjQC1VhyyeX3uVtD2HjcVfrGRDfNgmbtICspc7Sx+R
7QWkHq/a/zpzFQp9bqMwM5RMIGsGvkheAERLz3FsFnzQVsxOpSJ4Q5H+V+4QKd5c
qomP8VZkRHPf7DP12TAgnsvVm9F4IMhdXdr/rPJBsNDtiZ9VCgBLygeivnLaCwAO
ygftqWLGJ3CiHGFQC/oBzGudHqSXyPWmM4nobMz9Q09k2pYLfSwHFium4qsp/RZv
8tJEtk1/8Dt15wiC3YaHrVkcGFG/mRTAG+kUN73i7AkSg/5RMpRfHNbWWklk62yK
v++/U/QSza49dQ+oeYURavzXeejNRpBADAjA/5GcHwCWKoKUZSnhSwT9wHZ0mEAt
YdaasJdFW1OyRybVq6FSz1kdsr8XQwGUkQ04NwSrYLn3KQBjJNppw0RMg6wYeqQ6
uV22eegjnv2v9MGjF6jSAj7Bz5ay8A7EaL5Ge52iy9cT0BaE+2FdTnRJHuo1tsoB
PTNATMedHz4LLMpWkTvf3u3vsGaXUFPAqJuNRn52+pmElb5sPw0yqtVz++36mNw0
9kAIo7/xtfau4Z70mLK9E1cOXMaLwZ9olQUBzHJbjdi0zA4W/gsL2od6cyXdOjIH
990bqJ901GmUjTmwe+yxNbTgYZHj/9oyS57ead91xRbQgie9Of4xtk1ndOB9S7xC
rnZs9tebac7qmyyXCxkkyLk039iPOA7TNxhrHeFi3OMX8BMdgQzoPDFA6w9PovCQ
LC9CNx6W80xLie/jrkaVXXrUUXq4E/ncQerd4ngS4se1w62McukiSjMpFdU3GTMI
hoxLwvv1wg13n4V/yBl270RoGj5wQBKwg0hd0A/71Pk9PiMM6rkL/fH3V68Pd40y
+V1jfoY2orF9kF/6IeM5JKKWDzN/9vFY3qH22LBWHCImrMYMP9XG7lzo9BKlNAs+
qpQK1Iy8FAkhAwSHiPhANk+h/j7EtnoGfWVwGjFcchVj9aiq1RPrNST2obhdUkdI
PjN13Dbefg7TH3mz5za9pV0fXjIjo8j/YjX8csjJFD5NRlcyZNn+fXUfLK4HX+T4
Kl2ZghgHlYtjXDYM35yKDuUV1ay/S1NiZYZervN7I5xr+XVzRcpVNL+MzwtMv4yM
5ryTgd+dpDA96d1lrH/nQuoQKKNEgUpkoOAw+uIU8Nwfur5X0zUTvYdfiJ3y9Cs5
hrstF6eYOcspR2gSPB0HCwA9iqCuv2HUyAlTW7WbsPI+DDY1DxAys1LXp9TJXAXM
HGB4NqS2jkf6F4aDmVXcVp0CTh3NF1VRVE5cSfyF5/BNumPTk1Sp5pMBZZns87/S
ppq7tiYvqW8cXMC2iZOuA1GVO52oCJqJ68Sy8hGCXtfL6lHU7GRnWnn79kvb/KgA
2E16N7Bzh/K8A3oyIshXl4+REXt4yVBGcXwGgPmTL13gdynIxln9tXebiYttt0Ly
JMxdnYNZsuc9IKWwuVy2+bOOmLgGY+KALrTsJzSGxlj5/dya4odGog8ZQ/NTDs0U
D6U62EADAsxJsAU8K8M1Dd4ZDxeXx5BwNmd1beXHT1jRhECFKTxyHBHE+RM855RE
JmaTX0Tw2WaZQbqpoUz6JpAeQqLIgZYaxljAMeknNid7Xg/zQC9T3TCf+yUhjD94
3NlEW4F0O3quDk+XENO116Yn+crElsuBDFPEc+OL87tFxpsPWj0FddKIitTbmIb8
SwH8c9Wsr1ONBlYXlL/SwHneI5r4RCdHXiQzoqcqzTrixUgEvYtRU0PfiMKE2xxu
jF/9XoEP4+EcRngBvN/RZk0CoXJawZSY8iZQ55SmC7CJ/epK4cx06TsF/Tph641E
eo0AeTrCD2eT0cZSJlFzeftgjt+ttzBKYxl84Gkco4GE4KP+r7BU298UJxdN7UU1
9pEWUIacTt1sdBibT8VA5V0fOAs/rDxPLtaS/SoFPhd9CQWp+qEzg1IPEeByDq1/
eTnMQCrjJPcYPtwRgNNO4jc9tUCNC5mYTvKiAmrXJJjmn7UE9atfkK10bIGtEiun
NuHaBcLIAIQ+5F0CF5j7gqj2VoGMOalvOJbTHz215WmQB5lgzFkoSWPOW0ukrz5w
RYTy/zJb7LJoZ8zwtg21224xWYKhj23QrdnH7hgCPueM6G7sjisS3T71+uL+4WQ/
6DcbTm2MEWRVGKVLWzZIuj8ewxj3/usWvCNkplcS8wlEbqudezLxj3Fk4WjvCM34
8q47eE9/SuSV0wNKWlM6i1jDfyLb7YYJ4+B2dNUB4UfCAYIPXGeZjGAIeSm5Rte9
+xqbXGyxJ0WnIe06o8WG7fm9rI8WCuE8lR+peDstgZ0/8it8HK6xnDfMaqiWUBtE
4eeQ+6cLK/130f54dYAI+ak+Rv13lRxSFQIh9eOsMvcH6IO50FC8othk38YJMHy1
5M5QQ/oG4e+HKloMsmryNspyxE8vr7696+OhLVdEauKU/FvTXhQ6AinrJ5NIlARp
2y/dLyq6Z+HF+Hp/mzljWCT5oME62Qzgg29sXx9IobwkJvK+CNKau1FJ5rHp9wPt
yrJm4wjqQVBfS2g45bmyn3JGABd8H3aZDQJSKpsefj5tz9cYEsfxIAuUP9sCUa3I
mhtyd3YvxricCNGLxdT4wHEshk1SFP/cyT5tA1RqBZUmcMtIJNBOsO3FT/MygsXe
EdL65aCq5RTh5RDY0y4di4HMGgaRohLho3sYGqn8w5oMfS6eBlmDMludidTAYUAO
Xuq5XAWqVSt3vAdeqD0VHmdzZKxpUV1gJCrurIyRcY9qhLLEI9CwR8ZUbDc0s3E/
gNzXQhuawpTdCqeDpcWy4hGKx+5D7k76BXg+bhGDG0Si+kydxo0iS3flArZubIKL
837DiaVe4oH/TJTU7jJdsBBOQ3uJbkljivkdNuOudNL9CZaprnwpj4x+QqyVq84U
i5EDzIrONTiHhHX8dTsy+bIDZ7IVUcsAKM2056iZfXCej8fy8WI7JSl+EKziN1tH
V1FpeOrBzuGQwc2BzTfQiWt5E9UP2Zcu/an8o9p5DGZBeBkR4bjD5uSWJLeCyMFK
ksvAzJZrRO8ZcxNsDRgSs5EbASFSmSlcz+fqEVShpF6pZxCEy+qxDAfnLImCDGzZ
40PBSG9VjAGBQRFbLZRBmMv1u1uajvUptQVaYNylB+tcJMV3KVfcdf6m196lfAP1
D/ikkKeTLxcGqCpymjNiYNdBVCm/Z1TvipuUfkCAVUq+4ck/Y8iqiY1x7rLECNEZ
3i7lxZ667OWrp17u6WEKOapl4ZLe3aATNoZ/1H2fH4hH0dNTQO0ZXJXrBfMUh7YS
HlU47PYdEkVmmI+WGBHJ0rYQox3yay64tW6o1Trk46N7KxgzLWtg6txHpGYgMxPV
NMtL1frAzL3uwRYID5wIsrctrsX/CbF1SCxl6dPGNUeFhrVNoROchhew9/2t0cbi
xS+jhW4K+Fy7XoWU7qLKxZ+wlHEgPbMtRkwtFXS72eG1z6CVXmGX77OTEImda9he
bhxJZUX1n/Dq/3GbaNYAAUw8C6V4DVOpKsJE5v2eFiNQM18ZZ0ffdWGgSmNISXSn
23K4dgkY0OJ/si8P7gXo/VekVSdxD9yhA2doXHUcOeM8RA9xNm6Vi/W904/XHK8F
TgUQ3ly03DiIupXC0bTi/f7YV5oqn5kCtB1+LTlAexgBR/u6i7ZqYo3R6VFcXd2x
xqC5MM82VPmxg0hBOOWxqYggmk3xjNuOQsBOMwyd3OaKjMkDgXaoRXTh1FUdWw3/
B/37eIzrc3G7QwflBdfuGL6/se/cTOucTmkUlcL8hqGPS3m7qnaELsTfCXiUR3RU
z+3Ok0h31+AA+2MEWmYpxXUQTNnIbXhbEattfzkTjs/2fBOKzGSbMSqgjGlTNI/w
y2Nc9rcQmLBdLkl/3fjYRWCSLfSKdVDMRQXqT6F0AgCBtgll244Bau67H3YUSgZq
9H+rN1DL+JWA0ql4OyftgNXJGfPAoqkwZOKWGc9k+lk+hnkO0xXIok3fo020hOvN
fwj2+1PuJINchgi2Lvl1Fbo2aSYQmEei4zDM15vMcKtYCN2smsl6TeUhbdiXttnA
pUlLpj7BbG+huGNCLaRZ5t85jwwtsam4IcG0Ln2RPtvavEcvShXQ8kn4ONxAxtif
ANBXZlyYFbaTzVb3tErLK9Bs7pbCZerkrOKny/IQZmrghp+21obpmsVCACbsXqxK
sWYTIyZEhyXqb96TpHE9xN5+J2y8bR9O1JODUNIVC6bnnLTNLWLUz05QVnhHbaGu
QwMF4+3UUTmeCI/npmLFi0N0oVHJKvUaHXE897xUg6p/SIrRd0TZWbAb6SlAP+zr
5awv8aHmUgRfAXByJWt7aTZBBPwP+Ics67xn+rv3/dSVASkZ9uD9DDOwuH7NqGDg
lq5yr8JfmpAjNEaySP9e6H6XEp+KOOMLZkMzDPUhuipD58xv541ZBNenDbrye2fh
oXkpoTfXwQ8P79sGaCQhbz66kYwcKqNYhjrbyi6WWQi60Sst0tAv99B79hO6J92v
pvJ6Igk69fWldFeA9B3aYWnMf3N2juBnUyzHGAONH6PtKKlvFUsEyMg8hiwhkhK5
d6pPBE7taHQSAlK0ei55VdyFOQtbgq4dS3nuSfXlB5TCD7ZowUbpKCHosK1upS2d
0ftLssxA6alc1xRpE+G3yZ1zx1k69X1idfNZfxP6m2oqAiJZQtzZk6rBeMCEqMwZ
+7Y+HHYoRwWGCvPIzkIxLeQMjN9JlRzzH/D5dPLDAX4tcRqFah0GDZRMJnOYZZJf
Ipc5DX99Aanh7p5e+I8ZkDbZNNmL+ZmtQiHTeockH87IEg26D0JjXvxr5uGQky+v
sfmJoFNN9LiFmvCzRBo0TyAEMlURFP7hXsaog3QVl9cvFvhCRpaiEdhor+BWug7X
ImprusauI9AYv0sZtu2W5kgjWSXoCjfGx3Y2ITdACA54yWZqE/MV1sJXtVvdca/g
kTsMEzOqPOlBrjWRQmUlqwuwNzYwdQtuS63CN7KIJFaCS1jn9iaC6Y7H8aOoY5Xz
bdo6lkPWrWNnXYREhr/gieWTk+8d9Ol3l7T/nBccBipt6VhHH9p+NkbNZBUy8tfy
+1jFbtKTi5VaYRPyPHld7K/R6KqU5IvsMGEVNEPLzQRP7K2GEOjMmv6/tqDvalbF
UUA2qn7ev6GWbzzDMvYqYX5vc7BwkRq82NGbmDvEBzS9bhvDdhiWRjwrnMQ28+a7
YcOssDQS/2PcHjgqNSApD4Es0LT7xELNqmI8AhMebqOprppe7rSzf0x2/mksJESr
uQ2BWGRYXEolgkHi2L0lkpmGMl6RKOkyXN+sJf2k5QvBXQhb9gtLrXpa2mdZWA64
YZNk5kLdjIlHAZrnqmw85FNz8hxzK46UfOGZpiYMF1iNJgpnZqqCxNAd+fKdHQZe
uPlPg2VxEKbPo3wMqQVWQB0wXzgFBhf8K9RBwQMJ9od3OMxUWoFJU1B0DugxMbF7
BgBsyvtSRN790I9OcALOj4x1+PZIoi1VmsT+FcJVS1x8WwwNXyufj7fbhtGrmIQ5
fQhLDO8O1KjIDwW6mAfH3yW+I6gemFOUZYMW2HmgF86slKA1sOt63d7BK0L5BZzn
g4Ol0KZeWi9u4Ucp9MDvM+rtvE9sqMOUwNpOq8AFpYu04VJIgWLNtolNYOTckv4A
8ILRilam2E2m5T/LAJ8lAr10jnHbAZY+sctAqQxUyTOKh2LszP2x6/pzksOaPKLr
L4UhD3fdk350TJJFkOD1DwMz/5Ijvprc1dQGiDs1UreSb1rEVf1vSK7ZZkmjpz0f
yRlsS0unUxudY1wrE3FyVIeHdJNlgwywgERDmOE5frsDPkK+z5E36R+GfAmKPrFX
I72kwwAl7X1/YkYwSPgbkURVeESktujkc71fDlf7AMZYb5zQhqj8OBn9J11KVUYw
/POUu4WtxDZNobc7IaDbPf24wp8TFa1c7hl7l0Nn9hd+l99Ra3VDJqXAtRVIH02C
gWYBxB74KiRTW5hmn035JEBavbzezolfrkm303bgRxVo5InDguJ3sA+xFDLhZstD
66GJwlpTBxkbSYG/LuIRYRXdnZ3bYqglsWeSBUol1HKD7YHmHkuLlFV9MhQG315h
EFtxEABj3V8XqVQis684j2o2S2RIQweBu4D/ZRqWFZJMTGOIxZiKHy+J4z/55e2t
E6zJw7OkYKeRnUahWAzm+x2IzcahUOPntGRcQYQynEicjISejt9FZ9emHRK0ndDW
4+XMbnCFaZRui/ernvWwil/i+DMnv/WVc6SuyIGLm2MNtr0UD+bI3NGpOVfEvWTo
XIFG8NtzzRkDp793gvTe6p3CwnsBQSejILUjnYVHprk7vPw0vT35IiAQRIiKsptJ
F7XLjxRAEyT28Sy+tacL1683XDepfMifghVzmiPWHk11q3alSRHdrx9paxd0CUJR
dtAkSuwojBBpyyjFpchHsOpJdFxENbuRgDiotSBRZ1U8H3Y8pkCVP5jYlkjdmTO0
tx60hol2n+qdizSZWLsDIl6D411/8d0t2iGKdjWM4tTDWg/f2Z0xVM849JAw8RQZ
YCRgLXsQW+gCa74qjJLp5o2n4SNvV0lp6VQmhypFDy+Za7ilhnbTIftuCpF8xMRC
OW4CNBf62kA2S8JVqcrSDDhaHE9XZiQLXKw3M1vtDAU0wcZJoUMkcZfjz16bJbUC
QKo0DKHsHWdeLCJCfGrtuUkEqVV4HL3zh7QwXYxQuxfBYABks32DEO4eEC2lLjkf
ZixiFhN3xt/iDyGXBOzTmi/52zzWuZBhMphk6hH8YN8WSD9VdD2WQsIRqyzedKRy
0nTR3uRXdFtlprZWBtlhswcAzffhNLov7QBJ4kDalzSDEDQgqwON5BLRjMERmPXJ
Ofax7o+FyaL0GACOq6srMo+77EcLs31ZbsWfw60+VeXzcA7taAaImDrD9k5oSOJp
8aaQO/6y9PwblDP6YqxL8xKpscEohixnNUzUy6H5azyqg+8/FAhQuGcneD/D6y+2
aNL5Rqk39buGgLc5DbgyRpo8Z5SsdTwxp5IIYcg71PgLfdJ9HtPF5tfj/wKnive5
VsI+38CQh/uh1Ujn+DYPeSAH+va/9w3hxVh9yT7pIP9xewp0mBqnvABtaiMjs+ae
wxMgFoHkbirIfQ+S1+uT4AMoDbki/BhYD5bnl4vxnN89wW/oTmaAtuxsa8wxEJg4
1SZRuOdKFGTwykB3eANWp9vLeMTT4grTitHWi0Cgnozarjz2gXP8cBlj7AThO3tt
xoQzJfBoggUyzF+GkmBEPopCqICLylv8Jc2BVEYZH0yZNNiKGckpNfW+hQK5xVqZ
ZnPkTIxZLj0ej3j1sFuDlYjkWRXXRMiIBjb4Z0BlcVsJRQIWQKazcnYtha00IHWu
cNndjZ7Dikmn1Ulf0jbV4fLa+qcxAAYndE8pcS9Aa4Cf+eOoFxxAzNaCOrMda53a
6aLk2sN2D53EXsm8NU4iWb7UuK5/ek6+P23DkCvDfVCgCxSTguHqbPbeVPyCPRI9
7k4Ww3GfXKg7332cwtt63JBeWNlSTiFkZnVflgpw1aFn5B1yeWPYtESOtLYUUYqP
e1VBUkBVWW2tsL8/eTkW8OZO5m0rey9jUhL2jP871NsLiGNW7dgTR/mieKo6+ADW
ShSgr601uCB/E4RofjV1Jkg4rVX01ZY5VR5kSQmhj3k8QPgKN+4k+D2HkxQQE5Vi
H1xee9f4Tw7wNQVDXuWxZOgPQrbyqVIbF9xuqgkl220pUUET39tLVwuOjh0OLt6m
WdFmUSFfqAGireceZvjpC0xzRXahCOBLHdOxWUbvOWFIXTeOkrGnSHqQktj3UjOA
zHV0wvzGVL/6YzBbk9uEoEFul7AVHgNTasATaPG8zz9WZ7R/Y2c6Ycq/mbozVZKL
0m7D0n+ymcSg9EHkmg4fknOeAVTQgCKg5j28uzC9m0Nuk7tYJpRmTWkMR/yBnCdz
wW8umiMjmdN0fw0TOAa27XMhs78qQfAhHHbYSDlv4KZIZ2XoAl97E6LgWQU+8d55
U9HcQyQB3A8JSVk20YEFWRpvhEriQENX/lrsm/sv5QJ9cDp031huQ20n6pQEGtLy
2k6F29a+oBfH1RGW3N7BlK0ebVB0C2sOlG8H0Li0OEEdS6X84Y+/SHw//ghlyMAU
R0sMUN6aFTYG05jmfkeTqc46tC6IsSv38TGhuGn7GzmOYWTU5GZ0LcQBrrMhXEmJ
Y1qNxiOmxj/0DrmCgyQaiAATtMkfJ+tJhymtdW+WoU+McFACghrzY2nCaXi4TBF3
E7J+Lz+oy9doPB6F33UEzkRv3Z5IdszncOFNLaiJ+n0YtJIx4mWPK2KEvZGtpymd
93Y8QdpRn2lVqHHBc8o/s2k0YqhscCwZL7lgqRSQ8KB6Kv4w2MjFIxkaogAIBB79
+nb0zn0XhBcYc/EPi2L3hqp+vxBoDWpMbFqIVTnqnmkqph9V0A30qPwNpnqvN733
Uh0jgAMaYNDvs/YjAkmeRGDMARksXBdS08S2J4npB6PmZREDGk1Vt4sThPjb57yy
ONo6Yjd/c5Zt8b4xO22Q1TK4fWf3oFolcuMXh6xyRgsFhEpvpsugN8JHTfcTpepY
FEEuciJ1MytP5SLyjWxR9lCCsITmtUFGSwqvpelFHT5M03soV85T6vXrK1+Y1fJO
C73oePw8CdtsjG6jsQH4k0l2OI+xbFFl85EXXUI6scfi42bDygA2xyeYzYtkRuqm
17Och7ae4pBW3rbbbxsPlc3p0Lcvdrokgh9d0fUoP8/YH4TVhgC1J6LPKF4EjjRM
P0Qbjm3KQvNF7pKcg38FaXDU8M7OiNCf8xktmHdZxc1Own80vAevs7uwM/C2ktQ2
SVWqGrZubTLJe7puwzq3Bx5+ci2IrWmEs9lrgpVNc5xrE0thJnimtZDQxOHK/bbA
MzgpN1OOQIejPwgcX2zilacpDhHFAgzLau8uKitSkLCQxQhEfP13n20mGkT7YpCB
/wfVdX+OBA5cPIuTFokuD3G6eNHzw3NBFUpa+3EOYloRDencWqmp1jW9FJ9nF0dc
oMVxU2Ikebck9W76vSPKf8xV7vEe03rC/ydeveQ/XVfpNCGBq5qIqYNnAGx7QrzR
HocG23hqFSuW7Hee7w+R/z88OYoQQnDPG2fsUuYh+PMrXwWu/sho4DUpw+3EVM0J
jo3KyqXTLSn5lioJP5OqCNcApHIJmocbknvHGp34TIJa9YdrUckQO00fsJ7HbVC4
oaFaMESavKUOUz5UbDvWRDeGQzYxImRUR647qwI5c7VmDkbF1uL4cWIWRRkQEBrN
wcttTCwKHqzSASzkyVw5f0sZZKt0vxsArAVC1mLdxonkUgZBDALeCc0MIqeXjUHX
lWMLdtaJvL+yqh4aCAa8dKfR8PYDb1fh2CcEMHI/KLjnfAcikLOME2FFrus6YnSn
0LOahnHkyMzUv7T0w6BRrB+5rlQLZ2mHUSten6zXfuRg5rs7rer6AsLO0NuU+c4M
xUYKjUk9zysYd9ePEIqXC3Xp+yBI8yplC9XIsljYtUgpmIr2Bw3YTcxPR5Y7prM7
Krzy+0igBmfXkYCG4UvYSkm6TQAlKVOKqzgHt8c4gGpTjK5JAF3imcxloIMngdan
P18DIbfow2hv0ncPtUcgqg+OSOITXYxgLZUNefdhquZZYNdHco44XQye3xUh+XIp
h6BvTAdIRGpsFbcSsdT1GBC8oMs2ln4/PV3CZjEN0bT1PiWOaaWrNaJZN+y06OlV
DWsQsD71jhsOPkkwjgEKAEf9DmN3BMhlLetFhIeRq9JP4S0rgUceGjOnyytZodl7
oZsRYwi8m/TF8uLDc8CJAmHPhF+zv6QnH2970/6lSoU9fI+1txyoanPnZTWvIPC3
95aSeTLs/6Evt/bs/H3Bcp4Mw9h61G8PyfMB5YDXqGcsHrTT2iCNEsSRIdc36rYx
sNMaWz/SqQPY7xQS6IoNwaUMOUAR1I03ValPEr7KkOzhnZZa4Nptj4db6xph7aOo
Sm5Vo+kbbzLt6POjNPFtxUk2oyIN5X8O2Yt4ye9PZm/h0Dj00ORDQRiHOg9eHHob
gOQQh3SANbRNAA0fWISPASfOkwkrsJKBJ+KHhPF3vHau0rHS+3dZce3pO73uYK68
L8tfpB6d4OxYo8rwT/wpkA6cHuyyMo8dHeKeI5jHDPhw7zTu5dc0O8E/dT0FKJMG
ki1cDFXSJfMWnzfzkWAx/INGd1q2MFT7lG/PRNMnPMzU94Of0zwhzDX9Qyt77EY7
C2ctcESeamRxUY/DyGFPNU4FLOgUfu59x9rb9UcYUYJKprKSLFzgSNMe7KL3a3U6
nyVPUSzviRzxVOcRZPaM1QUNUl52ABFPi2ll0OMe628L6OeuW59xLS+iVE2vOALy
enqfsENU1BWmzupnqiCCxdABLw8Oo8OVSSTrZ87+cB5bUzXA82HxiO7+WEfPbujG
1S7zLmIfXqCJ9+FIdZ/+WiREcYiGPQ2ZaIfGwHR2BdnJyQDp2AQY+K4XhUH5mYzk
qKxpliZkSm7Qiw0GU/DqoWpndI6+i3PgJuGc4N7HUDDQoFHCfqcmNNtlGsKpzzVV
JoRbeXeZqwzclg1qTjheU2iExA9DMIjhQylgmT0SEcDnbXh12jmQw878b5dYX0mD
xxLDP2VnyumpA+yM2Y2YVw1HUpJkACfWh3Nhs2P84MOUrmPNbAVaaZSZ7jQ7gNmB
enkVw6pVjRO3qSRYzWBzvX/s3jDDQqNVAHssWkzn4i0fFFPNFOoFkdmzjybO5hGG
7FsdLYceLAM7q1D0irPZdNSFJeHi5QRdku4jbLJ5AQ4cGSqfYm1eU/DnZj+mUagc
733WMxihI3KLjitcK9mW12gcsy2kgzIiChOU+EbOjBTfXYaYVDrJMeZSf16qkZTC
h3Ict+tUd0K7zun6g1B2bm+x5CYMYKe2WOW3+Qslh59m3Mdn8AR+5D27KOmm61/D
yamH7aLg2qvHOlw/xwutR1XFSP1wIE6mkR5j3n/eIxRap2rYopL/Ta6+6z4YpXkb
KAwPcYyarNN+Qvwplyz1g6RD6E8JwvM1ig9jd05mQRlrAOgjG2AXVLMxvNQjNAiU
6aBO1hmpqPGXw8nyFhx4v+tOw5uESFDJclqM/S2TF2rkq034DeOXREvtePIkdNmR
oRUKCim4UC0/GV7G648Jmyuq6VJUKE5aW5QqfjAds2M02gXTPT3DqwykQY4Jfd0S
cJg0slnY29YczpmXiXhe6D9gRxw811gaziV+yFSMfxa6vm12Q5LiI+n8hcijW0/d
PT5or+Ut8kmdq3P22Ewl/dVZ9VqATNDVnmbO5bX18ztu2KAQycHTc3Gy9NLpSN7c
pAdULeTOpj3JT4VCBXJjE+RpanBwE8FqFL+UCedfOpa15GWaHKov+OkQdTfs7FuG
Btv3rstRla3mzQs/DMCZz472ZlHc+aE2l/jv4jeJ0V3uEciYojEB9NmZ3Q7iBqy3
wcD5ekIZ4/3t74kJMSaeNOhWrpLlUdD3REK27yJJybtR+CAxXwIAdq7ypD/u5b+e
vcAIFkrO3tot1JyLjHhnj8MiVBn7NB9mmQkefvR/j8yMfSdEB62DrUgD8caqEYrb
mD8X3fTFXJvBY32NUo/V3wqucZILt/C99UbdbuvviUDHIrVSMFUzZCSP9amOLH2V
7CCCiX3qNzbai+robTQg+DZLM+O0vGvrh+U4LD4aa80HzQa1FtsVMiISljWID/CL
v0VJU75gh2fAEQb/rZepdSWBBf4A5NsuMU9u8/7zjnaXWtoPAEcpQC5HokCchiyT
seX5szJp5a63b2qnKFcwse1O7SvaoLDYayTT518KeGAILqdllqP6/8qAjXA38Rdr
BKwI3HbFbFTJpXPQKv462hU5+y93i8lXr3Hgyx6+jNM9hLu5RX6ZD12at19wWrrX
CK25rKju+EYTdmzlUVN3Qgs1EJwd5UOMTc/3jcHuh1K5XvUjsow8szl+EkQ+siEp
CIUY8LhC3umfZQM01Mudz2oWcowS4Jr5FUtLXov5ioB8wCay+3svFZeXVt3nzyRV
+IEobsfrQrq2FVObNuMnjFN0/lVhAtwRPhVnxMVmQ2X7RxlohSfapZO+B13LO9bK
n+V+tThOMdFgC8Yrn2J1rv2rxNoDArsaQs+fES21TuHTIXFGO6RrkkwHjk3OKof/
ulyQHeOC4OIcIj1pb/dEfvKCMCMmut8CoffUTX4/I9ke3gCu6q+ln3ceNL9bJ3or
5UzN1mHQd4N2LRoDRirzHIJ4g/WU8Dhwqw2kdDUjlNceylmMew84d/lHoE9ZS6c4
7KPp0kQHdHNS44gOnYIuVDVZDvD1ATSnbJ1YvX5zh418fA2hjqjVGg9hP8lyq0b1
DjTFVEs9RistAelz+7M2tNYb0+dvXC3BuJqyShgSaPF9BUyeiWFI9ESfeaaj6xZF
kRDU3WECPmiRZKiLnmrXF15lta4905JyqNBiRndOmM62IxRyLP7mg1xpO0DFcQpO
t+gf6Oy+nxfXNOHSI71DFFC0HZYyLN2LXuuy2mdlE5F3lTq5CrhHyvYcp5t6XnjT
Jz3DVHZoJr9ZXSpeD7mEcKmxcY5RcLkBkqdyYIgk2FBTPHBSFywtt7/dJBShAYTA
V8KqXZwiB1PVDmcb3pmZWIaibK8WZLZrMz0YzR6f5B5P8sLpsssIjl+KedPxihL4
eCKiY3c5k8U3Pv4ubigJctHGN7rYFIy6qBbWAj0tm1Y5uONY1Xn+ZlXVk0zE5CPt
aG0gD9wCbQJdsLp/f+EbTAd37qjj1qI+4OXiJ9dzswB/vIl2mC1JaR12F/PQvZsW
Noe00lniElzBhPFpaLKwh80/M087oJ1F0ULIW6JmkaXOGomtPEkvvggAC7MvT4tu
eptJJx1arzFqCqbX2eaYsIlvtC8EAjnbpuD/8dnDINn3nPpdnYqSDOzz01J6sPb5
q2i3ZIj9io7g6O41CpL4wJFQY835AcNBc2S3MGP3ifgipFi0kjRth5o7npl47bGr
bGZEPHpOW8YOX8Qfy43zTckRZKSLCEu/6obbA7+jKXjR85d8KbFTipjlnRPfXGbR
z1bOI/dST86AQuREbk8iFXUfRwLNK612xHBzXLIOmHAEaelsPqBuaAEQjyEljVH3
3ICEhU4bcsmcvgMYgN8bGDdwf6jUDToCkQLC04QJbggnTTMQoE4DQxF6z7PRYVwp
BIoLLSjqjQ0STBs1SV43wt8Ie/pvufjHGKi9uxdIrLkHND3gX0ksQRLdYUzsvM2c
KvHm30vHRC22chtBB9hcbxx9bdyueTW+dqn3FwmkdvYDpTEqcDmQSGDnmC0K5/Zz
HPn2TSdTYAQJrSVj/FZ653NZfhMbFP1Uns4j9pQshg72JR8bjblTIUA2pujnjdYd
WIMmiv8UVfrgyo7pW7lRv1h7MB/BlU3Au/oF6enp7UtFrY1GCkVqvu2cfpieTJV7
r/mt0SI2/m/NCsd35P/6I88wOgyh/jj2zQJtNaS6zfO/pRQYTgrHiQMCHRn3ZNSi
ZvD0fyMZCM7wGhoTrT7M72kz7YlFjEQyK7a0zFDzHGKnZguoj3Ly1rzpR04eJ9aA
jiupaw9Hnia2JhzHHE0gLuaKgS7yZ7I6HHuTnsRjnzDv4p6o5Bk93V7BQRTJ17s0
FQH/J++sb4HKz8s3tjJE40RVtC7MJn3ZxVvBPVdqX45V30kN4JMrXSsR95I0Rwl3
BULppYcqWU0uC/3H80l1m73af8WK0tVBAxw923hrI8GRYasP9wn/5GMymbZ8WyNt
Kjm14kJbkiHBp/iH5OCBUpzzFKkqEJTwWlBRctiWAH7w4QsGExeNowdap/XPfuXU
7uL5QrAQUk86WkVrP7ORjYYf18Du+/M9ZySJ4J29D1x6W3iUrhABlRl6vxcvCinV
ej+NL7qTgjx+SfZ5W0Pm1FqUYw9YPa32NBvM9pRlkX9LTV8HRx+yzZugTT38oYxz
9roe/Qa8oGdBPknTt1fI8/GeYweVxhSJlb09JkRFlrF2/mAk5L1bTCe01FHy54bL
AdtMiOsfz/k6AW7v6/jRI8mnrtnZ+OpDOfGa7JNwNbZ4DDcLgH8vU2tLToM1ITQ1
tKwmCUiS3+7fmvcHZn9+ZnadwuZs74dJBi8D9ilFUoA9++n+b46ePchV/j6i3Xty
Vv7oXDavdsO1SOVXf4bG9+baoK6KJvtS7+B9VnOeNQN23c4ieg49YanF0lLgolXQ
SWNYT0okp5lD3ZMSWM65sYzM8GuOWAr6qXdQbeDGeWmcGg3DywftR9c3norrSw2J
Shk98Q2rXZpaHcU/HYxgKDXHe86yJsfSHTuZpMc/RFna8B/RZ42IFVMCNgcr68iC
ys0cok8XIPSkxF35a63bBtIgth2yOQjG46o1X6nVuofuuto7wwJh1Axm6zu1J6rV
MCS6VcSE9Vj8eB5BZ0wPDn+etWI69FncdyT9FXtDr9QVipTchHrXiinOL13KELID
DT/bOrn6c0rzqCDsGyHvIDxTvfRwRx7+zY38HQdfx8aD/MC42IdZNhI3IBbPKFac
+Q5+qefn1h+mjPhLYMVln5f4sVC5eyDBvQRKhAIFryG7AbKBilAhkzIQHPtoVGi9
FDC/Yr8iFWrPBanFCnBm+rcsGCiEDNv7S0kz6bSmjcUJ6yebY1LEbpr6hhE0Wf9y
cAZ2jRNXlGRylWYXSZTx/XnbaQUWmTXFPXA8Od+RKKYUtlqWV70i09oBsPMIXKz8
d2DgCOAUqBl7tcsMaVBo0I/u26cXxGFE2nlSN2A2GaURz55xcv8s+lfeCah9gbOo
JI7ocL4FDz4aOYCCx1PytxCMI137H9bsAWSZW8yy8GxUx8VUEdQpER5uHbNDz1RL
/AuZFlgD767eijSJVyaMX3dWk42YgLa54Z04RMn8wT68DLsySHjgUA2ZUycDY5xW
tF6WqqMXgr23oEzRVf2npSaDIE6JMmopfXxi868EvGF/ILmUBtjL1u2Acy9P28MK
zQZh+FzyKbDprpj6isYQT8WeiSGqxXW2X4R9N0P2Vjt5fy8By0dZWZplDRj99NLo
OnIPzTSICL9j5O9U1HxDxpw+CcOauh6Go1A//LSZPen3kY+B5n0Cb9aB3WDEG9Gz
nBqGc+K6YqK0JDmmWiImD7wDrygEwFdNwO/TeKF/pWutZ+wACyk76IWvvpHOw1uM
oqyOtBqk2z8pXGrrVsfvQLlvpGqhRU27tN79T6W2lkf+ImrQ5ACCIIxs5zaU2b8F
UEsi9f1jHWnPd44QSza/Rjio4ZYWXV0hCyNMtoLmz6PBCxdfhyEsonzLhaHmw1i8
4yb2tbQs/IEyIshYo5NgDp6sfeOleIg5hXa0daWGwds2egvE7P8D2d/l/gWo0Wb0
33GUYWVkuj3SL60IIchbw4TINeEP1V+TZiqwQaFU+mQ7lFPWjvMkdRzhFuGc8SY9
5ZVuht+Cf5+TJvaD9D5vHvIPXnkLtqheKD9PeTp8ZxcuC04vPzygY8R/bxPETa8S
OIjLmfshVcuh76UcirLw6p1jM3MEaToZ3bjjG0H0U8zanM7meh6ASpebHMggNWJ9
OsJv+YsXSjNXskuARvbgtFfpbHS76ehROTm9QoN0RnwzpaFuCDfH/gGgZWXw3xLi
hGYgoZUp1ph2TFyzIx3jtEW8J4SkmBY8mAcjAWyIqXvxcuVjaIdmCmJPKsxZlUJB
dEexFFs9OaTOg3ZxGya2BmCpaGqzumUBhVx7PGz5vSZf76tzhJPDuTAaYz7Gs9TZ
uG5dmlkMpZqC/BcudlUw9eWhQwO12qC85wA4oGAGX2JthVXy0NSpmK/uUm3baTYd
8RuWzl2WddYR5/vugS1lovWoT/4KfYkrR5CaqjKPFZSArvvqkhoW7ZWJraJDk+kf
LorAkjbkVVSI/JfyshHx3Cy0v36oIttkOvsR2Ph619AymEzPo2kXbB8JGlWJrQJi
3BDVwxCPYJYmzNFleSiJzTOP2QSkx7vT0Gs74c7K0UIJIztAkASHz45czSVS4Gn+
KHF4NQa5KwtJgbGGXmVBz6h0O//g5cm6s5WXMKwdbcNwykk9OGdg74f3B1Irjt9Y
O11gWOQIv4y4SWBm6jRQdukXRBd3JOJ8dm+o6iJ54rMkiry3x9DNchIu7tx87L9Q
CFSEKtWHSqW89zSRajk5hqcV2UuOaBIJjtJQPwg/O9AVAmw9QOWO7fekjzauz9L3
V8fQ64LfG2fzYpbZaRt6dBSkFxDMye9V13ZxVJpsADuIREr2fQxmvrsG9OctjBtg
V8Km83TU9BQXRZOOAxBPTDN+bXWGlTzjeIdbdxKekHT+gj7N21GmmMEJvXOx1lxQ
dLP1SUaT0LaFEe7lbdLBwAnEKizjMKdn0wQgL9ZNg0xHCjF61DeyYqvT63vuVZQc
7I4bmpbJFY7bK86yp3LN60OBtDSN3CYXtM/Lc6nX0b4HzCMRYXtyumg2XYhyNGtE
GLZ5+6AdCBHoIHw+vODTyihFDpe5Ug51/AA660RJJUJane7lfinhm2a9SvHs3us3
rX3ee1ezVEnMKAYai3OmI0q/XDRg09UaPyV0ntgJNwOu51NNl34GvKgxv+5akrOO
wtVF39oANafi8Iz6mY8XYSj3ONoLXQ06vL3zd3OuAC+baNEpeY+ptGY/6boZUGRq
Y/gKQxG50NrUHOtln0Q+gpq9F4sk/tm3/HMEa2KY/zHbSra8cmx8K6XgfWlGloGk
XveKM4AWo9KfX4b2aaROvNouUmJUVFWYvjfKlMySllIqsx+XlQDCzrrtjs8OJ0Hj
fxLFxOj1jjKh6EFdY4ZjACCLeN/wR+XgvyLd24J9S6vpvf/+l3ZLeMktpODkAZS+
e4IpZ9HgJqHuebSQcz5xr5IgZNsnOrg0skjHHBd9B5zPe+1e8DyXX8PEVSuhO5ef
FtTk8mmVeVbPVbGrb8dVE5IbGGKxzlxr541ll6l9cfsubHOjrl1GM+UNSIbsO5ol
FBT6y/zANqzGsZrx3ZjXzjc5bVnZS1jKqzU11tl/BJ3HxS1GoSJozw3yvD7rnv6x
JtKjgYJ5jgomTNXmK5wRYhOUBV8sRM08Kl97QJpTd7TBQS3NEHlSwkVD6KC4ZSw3
mzg1C62a0k2sy/+SyVpmJ+Guyhf3UrIOjuP9k+Qx+INwEfRcWXdztIAiozqHZAfq
cnV4mvKgPQQbT98vvZ+syQTPVlsnKxqRsa2Q6mxcNlGUbh6jS266ykBrr59vWk6F
zjIDaIFx2LY1IYy+cFlprfRwaFMJHor6jxrTdiHlRlUhmbC7mO2IT+R6r1g5Lhfq
/rE4wHYvVsFRcbF0xhbnOowaQRA7UrHWLpNZph0dt9xH5uYDUIf/IBoylnVFGWL9
a31dereVZst7DUwGXkcIT1ncTRPAQOQyG+/iYdXsc5Lp4X7C9hp1chvcNIArXGWi
RHVdvSvAHL/t5aNkIUIuPUlzVtUH6P3H2XpAAuYA4R/vqSNPhSLzQP0ZcdfpAiMe
ONQe6mdn9dJi1ArDlKL7W+ORZcd0F5aNzd6s6yD1GZ6UdsNAdKyLnA7kvhEoDRWa
Ydr3hscn6FwgDEJS8p44yoV0vkmySYvCYiqaqglBME1rKX9676mnOj674hR4LLH1
T9LGalBgUUPAmuWGl71W4yefTjCqCQGg27z2uvLddRwoFdaGS2Fg6g//92utxeGy
0vdnoLmCrlqnuFQ1YtD++Vc2RY1MiZvL8RLtuu3t/qAeMXjUCL4FiSuTDJxhwMzG
/bvuY5HX0zZHBlJ17M7k8kZe+HgMK+gnW7y3gNK2bNC12zLiSbfTzgHrNifZT+tO
lsYDTSwKj3i8/CQH7z4ZNh0ifb4/Ial/i/bchClJRhN+y/bMwQQ4QTDlFwtRsP3g
zI6vYaxP6Y5W8n6cV3PeNSQmBNrXSS4VQn4VEkgdgZVC07oW70iP914Qro0HTzjY
hCKnuvJFCelusftjmYjwmxFpETk9GNWDAN5XII3aXEN2Exxem2MFeix7FIXEyEUZ
K36XNm0X+KRyc1bx9X9eVJjB3sdwRMkvMV1VONxuSr6DXTpOJJg0N1GEKYvnRcTQ
RfRJ+UHE+6IBfBCQTSMUcwqhB6+A1djOhNj9w8KCjzieclLGgDqccvWmKGH8WuJB
pHAzS/nVygiFKHKaElCOoDRjeXsGm3bEDtGr0WILlJ/8ijghvo8UHm8RV+slApIx
WuVw1BPHhCToot5UL4jnpa4/p8zMqIOVIzouVV+a/XJYyip8O6yabTDHyg2Lw0j6
I/50BbKjIik+9jA0auk/KU045bgYQzOjN1tgPQkT/HJdgVKV/XjowcSi+3NAdFLh
M1pPybM24lpZqX8RgJENBIQyLxUU8eHbkgcizFfcTNtMCIc8/0gBQ5TVaqvQTBvg
jEW5ocdDyonnBLd7QPapcu1WwT7VD7oS1Oa86iU0wpD+hnyJqX/ERZDZHtqwfiVm
b4ATOnskbHdU4MHL6p1vUwWOol5ZfI3M3/M3N0rYJf6vQFAixta4K2iHGN56kMzo
YRaSLeEdBQJjYnQeE48ZYeV2xHEBJORPcY8F1ihz81SDozb7aLKVpD7+vGklc16t
TPvdF/zjgCWAL3+cC6oZt7SIF3VQh1I/K9tL/ie0YzowYCiWpqCicxuaub7raO2D
Vnd1ml3ETNYTprQVf3On83BO0wHL0sZMomrvSaGy+dM53fFDmnWBavpN1h1gA9NK
YAxKzxC1+2G4xSnGAXMeAt1svzBrEdepD11We1f9hPQmas98ckuyXV1/lcjl+e90
OsRqiKNdhXuyaTVnHw+YwH68l1p5Il3jGvMHEX2JeNkJobiOUfLiLz+HxHzcTUR2
0OTbYs6o+lXeqk/fjQ768YeNGKxFTlyvjRykzA4zTOaaSQLddXrHZ6X3QRAxLOXv
5tuaiEejxM8CZO3Yw6VAAQcVjtTZHHV8UL8ha+/HUXp7CfgR+vo/7ewelFfg3EmH
tnojB77tzHVkIIW2c4NKdJReZerHIa7iErCYJ/MEsFgfkOrukNchkONu/16q0l60
JLuecCOj6swuVVa3WBc94Zoxr8DaJkLzz5bs3c0Gw8YfKrm+GZRtIgzZfSCnorZ5
I9z6SssZvP9vD1YV7DNRHfcILAw4Ge5vs+hFtKYZt+ryoDitzcMUiZ1yG1v+zDcQ
g2Fzj+eWVwkN1NjaQbJ9KnT9X4bnDdqkphDI7r7hoV1u1DUPEnU+DETiOLBdG2pY
yZvH/021EqcLSdD0AAMeF2LOhraT6VN4j1eZ4sEKhO5P1f9PbpVkZgeebSAf7alt
O12Ko46iAQedMd5PRnHn7AZ1YuJF0IEiMIP4u31tB8bqw+PbK+GZtpEZFd1kWaUm
Ns1ktiUVvJtoOJXnerfZK28j0WM6bN25+aSkjTB0Y8gyP8R6xgOFyAv0KGM5MSeZ
CZ7V4K2Bq1MIXlK3/Bv4q0FvIqXbY9ZdFThA4y8mr/Mc1CqHbgyRC85TGIb3DYiE
joKlTeQH8LLeDDM5jZF61pKOFsDeg+CbkJp49qsq0sWaDveLu36YO2YSMK0pPYwC
/M3OXRnHXPz1rNYaUuLxXa7D/TuGMg71TbnbZX+BujNE1jhgvptgiGAbHdSCoBs5
s8AH0rk3NyA3HVrRJeLcUaJdm996GON0BbTGZN58xBDubf1nbkCy+F9EUg04dpe2
d0bKzVueBQvNahRmzzboh4TTGNE0hsPo6bHViJxE9lU6Irmy0gJXN4LnUPnZw3oP
qkufdzXbtAI6PoYbYT0R/iuUYTDuVhpdvqJ83RBKtwnZFFdWHPjVd29/ObQgsPw4
NDPK+KscQgIvZUaDWIFCrc9uFRpIVGH+BpQ5au0IyrRM9Vw1qJfsT6yBf/k+nc7X
FdDQlccR7m7KzL9Y/ItwGDYCdt7q0dsORxaNJnFwxeT5NomITnBqgyK1OSIi5x/n
Zu7UwGCRhdbYrXT1Np4ZtZ6lMqh3fbtow69Pgb5awU/sxbjfz1W97So5Sm/bNOzX
1I62D20VnWQfFLn0R3y/l0cj2St4XD5LmW2mC6u6VRm2EsbWbKPJSNCmfirXG4sK
pGc9NQUE9YZ7rD2v6cs9KHt3xsCn6+hVYpAsDM+BCEM0KAgjMsmGYuYIxNwI+VAI
Z+RxYGpFMd/5Qlyf6qQpAI1YW74X6erhki1Dvei0Mt5x1xKF90FVKLqEr1MYZB2r
ACencn4YWyAaKvUdtagIUAMSm8yI93eAhdSydRCzcyHW+mh2RjdYd1lZrcuTRyNP
0f37enDuAK90zyvqsQ1m01tv9yWBQo/BDzUqvSdW7tnXq4rMYNLKQ628vz6eUjY+
YikTj1q3jDzW/CQ3HtjdYAqtTlMU0PKMNwd3ndiZ8wAuTNDTU1geTLJMrb75xKty
huUfuwh1ZymY1hYh8YqhBhUZhT7Sq1fsTWKGiBN8/TfGO9ettTXZpc0L2ZjkdwW9
kKVlDxx7ypdpM7K+KuI3okiZQgDvNh5++OkTvtTDeMgPYu630o0MuyK14+fyFNQn
Kium3I+tkGht7M1c95phW+Rwyg5A3sFn0v6PIj0D2nmW4WfNWcs3uxC69f80AlgB
vLcZrtojTiBoR4amXpzner29TnVnk1yz3+EU1MPZurW0P7fo/0XkQd1w9BMESTqh
HLN1rvyUIChcLYHRlUnjFqcoN0h2KkPv/1H2XwhfF1DpEziQoV0GChAoTgxIDmcE
BC7IBJ5PS6xG4ZEPqO4HZOcWLbfyMlbm0hb6V4onNX5r2g5Pi2f5BVMLvcXN3c6+
pRDvuGDdE28E7dWzAOQChwevR5igyUf+y83cVmY4jOFqfPUf+AMMTZsVU26+inEM
fuU71HtFVyx6N4cITR3bXcJ+SV5dlHTAknzibK9l71X3Nb0nMqOUPyxSBeLhVfC1
wvd6KS67LMwoyOHhmiiNLVJMQf8+7fknQgBaKGgCOrhwSX6g62BBuCB94PSBqm6k
Cq5dHpLlJ8Ehovx0+W7SCVfLAfv4v5BBVbhdF+FlSvuTBh3kc+aaZa+14dGxq/zk
yAzyxYYLVutrmcUmnIGeBr4X2DKj6Lf3kMHVMryu6xv321FzbRWgVvWbbYyW4yO4
ZCQWX+6Enw52p2JHxUq7okAywmaJRGqw7hfZNQkyclz3/SxMVfDF+Qw/oJapb3/+
cT58hj9xcSHv3gp++xuAMVr0fK1Gh44epGF3lAHKriXc1xpVBbo/2SMmNyRAdTXv
d062YRTWSeuLcz3prsked8WGwalW1Z+GRmWvRMJH/dBMEp9jPtb/dSrFHCiYUbAY
D+rkquxZH/yhOUpggCW+K0Iwm/9xt+Ozrjkv8SCTwSoVePziS/twSVeV19Ssglry
Qbf+oHbgUYoIlqYW4l8+FVt5RQ2BHvj4q9yA/9ECFXai9sLjFrcAa6dyzLd++90N
HJS25xq3DL6gcOrwvoz/qWbE+tsEuh/xZsrAx40Q9duzImItL/woxbTSL4DMFX9+
tArmMT4DiIU4nI2nDi9PhIp/YHWL0DiVW/d8D8EviqiIIyIPBNpSVA8SPf5LT4G7
Y4UVqovhGYDH3Vs2PIWzI1gvc9nc4AtvjqgFQDyM8OgkSeXm3okLv/g0oOqNV9Pp
CC73bSv1FjZXzBTU56ZiWRT5kmoqY7EdIa8IrFkB7qZgplVVuhLEuDtsCkzGVqR8
LzsDxQoPceYYBOdrPirXMVO7qzU0kRqL8l7Ud49dNOZhdernm8MBz/7LwMyk2ND0
aUJMj8aJ8uOBzs+qJPoQqvW8f5GDgZv30ipA7D/0Na34g7u7CZt2Ic8sJEjcJU6Y
FfoOJEPo5DszIE7QPlsNAt7FSwIy69kV7CFhsR5IpgFSD9CsRV/0enkC/ygtbIwx
ERA+qCn5bjIN5gsuHMibkD8JaGMg1ixJa92hJyiC5sSt+p32hShZvssi/SpMRMUm
ywPp55sD0IKkhN55QPP0nXJMCboO6PJOE+a+Mt9YKW2xSZoIOwoKuCwZ70CWZZXE
kF7IWjoKYrdhdMFQHFJZrGsmdQlB/U/ltkSSzBnGYBEnxX2YNOsAZBQapulGsZme
Quf8el+YBnu1otEYFDxVoQuYa/JLohOLB+hlTwea769nV+4ZycoT0TCDR6mtN6hJ
0llyKNKh35z6w6fCS13G07COkR6Xs3NNNFPopYuLd2YZ21u9a0d7bj94uc563koB
o6Z/NK7oMKWgrAOLT4n5S2oObfhScFae5Mzcefd9gy1PSqxNPnImxSByF+lBbJ2g
gNfsZkOrVYDo9LbWjo28kO77PD6h/WACFB5yiJjHzGiQXOAytnlWoyUtXXaPv1kZ
9HxPwa0b4tABY6hR+9Vb+bcq7YmLcPAOTp3Uj2EruK2U+ag8vO1a1kbwpbaXcHDQ
yZSBe1las+81rgRDgUFoyDKDQWR9ttXWRXN6G8iC8REVLrkDIHQgU1QVu7Oqqelr
k4tUEdaUmNfQUWdgkzTozgTwpOPIY+KErF/wVwS5Q6x9KzkXWIvR/GpPkGqr3C7c
PAVaRSKlWnzLH/YxiUv8unI1tANJxOHEjIflNHXHV8K1fIhCyuzaN3zo4YThJVGI
nAbtSB8lXUyH+R9MOFOCq2GqmDH5PdTSjhOKIROhESERktWxWyxR6ERcI8K1FSWP
WFpPxoUO+4bXhT7qrAJ/h2Ji4iwP30KGUBXwBxaT6XBmQZnoB3VYgezUi/aGj1LD
MZolaX3rEJabLXnpSTFRZKAeY43MfUpN9xrLpz/Z5OyNhsJjcCXqPAmv+lv2Hudd
T5y/z/mAUoi2SzBZT2pGAPG9qrT6O0M5IU0SZnfLPKyQSWAz1F4B50b1nT7e0E82
UZyvxeknIbkm/Bl5H8OzhPQTmZ9v5irbz0erx/KnbY+apGtNP6C3g7RwME8WZEDf
PZtpZyJ1pvc2B13ACBMe1PGp2wOn8NXOeFclY6c4eJY5OnLTB6UcxCu7nDKBnkDu
IDACffFql7NtIkiPDv4wTukupqT9zseqvL3Cj0Zn3NgDIMY9agN4H7vtRY94ZpDR
gCvQDahx3Zvv2B2TRgHQv0cNSy5D3tdavnmP23/52x/QWxSKH8KJczSHkTkPBrxX
437EeiDZx77iVIHlyDx2SpXi05VU0hLCGEZN0/R5DV+zK9hRme9XpJGFkAcnHgoD
I4I81os+82laZ1hg6gNC6s3IP+38gRbv13vQfxrKLnIla14LYMd/FEldTlSsBp+D
ah1eC0OTi8i9afgxtBx3dDt77HyGWfQokiNgOnXPzhKUyva6kqC5ekk8ZAoc9F0i
2GR+iEcrl62RXe1cyKkuMzlrVeAkmivX4rZaeObFfEMZEYyGR6yJ7bIoUsuBJF90
SQw4hD4QcBMV67x0CvQ72fX1DH2Vx2FQYsgx+Wt5HoLCMFHleIWbXpzO1IgO51oP
kixabc0qTojvkS6oq6YNcvO8CUnKoF7dLlDA5Nsz9tJbBZWF7rHHC7j5Scp8Tr0W
2b/mgLwOJMKa5Zrs6EyJBtE7hXrkJkucYAECk3dDrMsrsNK9Cm/oMmchUEplG3RO
7+Lek2Om+6v1onK3L2B4BDySqUFUIFaRuER9KewgqTI+y8u1lrebD+echHFO5CA1
8Hfn7YGll21ifMefCo7mWvL5w8aMAOsK3Wrmt8h5LPMbQwA554iIYAgz5wWlceAV
65hMNIW76a2qlsU+SM9JBtbspIolJJxPT4OR7Gz9z0S2uprPLyhQaebTS0g9jVR7
/AA5Bpe0jqwmo5YKxE65ifq9g2zP4nNrgYAz1OQSbCgWpMoQfoonxFCf7L6jJ09l
V9rSD3J4iVr0wUAdJYNk3s5AdFDPl90HEVnxWbx/ZJKU7rUtbz0ei9+pCHEFeENV
+u2NcQbFEmOQ5/OIEpIhLfm2Os44LCdieFmRFnFbLfmXEruwK+Gro1RwkomnS7wU
OBjj+TCRX3WhgkU2dP21IKV1Cm/bWIVQvaQXkbtVI7nlOBmMRppSokzfUz+2672S
oToy84TCfOZvUp2NcM29r4kUW9fzliTOjCIlFOrqG2oKFy2W5BoIbTW/vIj01K7z
4l+/D6+O0jo6O/Z5FAUEIrThjqvfWYJWjddYsB9nTOyBRo1GKuqcMHJBU0GXnDMO
WFuVa5F8UDp7CAxiDHKOtF7VE3ZniCGjX6pM1EaPmq9i5Q2Mnz4TCxdG5R9DPYpw
MwluNvHCmtamLZ4cOaE3yIK2LLRFvQjQ7RXQaENPUl+MoDCFeCpO8xPloAbKz6tn
ctUb7nq2wLQ85b8pv5bN1e9F1Rebi7Wceie2iVQmI0otvW6MkcPZmMJk8eq7m1/9
3wc4Zla190g2Boa8qep4doClC3ri6u+R+IWQ6/cR92QUGlSY2EPKrHUdP9ZlBVsh
kD0Oz8QkoKIRHOqmcqA9bzDWtIZwUhHNx0GUgY1oNKbhZ3XtVEYorfV2M6G0aEfA
cLz3AM7UaVSa5sv+/jI2NdpPxaPwYMC1cSD085y8smVFxFVPuW790lgZmG8tAEGq
GzAxfbx/3ey2jyVr0q4uy5XISh55EEyXCUL+DlJH6RHEi8y1iglqibdnmRHnSj+w
2r5j0y3snd02F7AGg5hiFKcaiMx823fNLSnQ26/pGzMGXX0K2gPABolC/ADerTcm
oKOm1fnjNS660w5WdaI9FDz2hKl8u5CHrBvALkrwPK8Y1KyXpPmZjJNb7C/tFLjm
PShdDLFWbE+mJJH1i6ADXxjT73UPM84Y0GgaCAkkSKP1jbseJ3CnZNLzdUIjIvp8
Kr5HpJh8TrXdjq2V+prH3umvEAQQcXvTjnMKf4u4o3ZAr8cqKXCkPXhfxQa5qKRx
LWtvGgv+UcGZ/eEoWbZun7joiZzSpM/rKleDf3bvjFt7BM5rArCWsF/pjUWg2LRX
AKzeDchvEGmTWbNXvF/ba9RRCzKe+/mr4vKuFHUam3hQ27CPB8A+NMBfGUbB65BQ
E6Pl1xfwDdUO6egA7AB6eaKsxj0uHozIgh0PMpf6t9TA+DBzeUHL1GgyVEU5cHoc
3UDPeaY6SkzOb9whRCKyGxKj4cLVfn56dPgChsL/v91JbysAxb4YIOmf28H35hI3
2iOn6phIBwmijxS1vd+QIk8G0f+i3kmr160JLSXn6VPA106VJBtvw5t058H/gelI
Lmxi65DVLr8k2aRlZNV4QyCtKdQWamzSBXAwXc0Kl5rlZEF1l1qVQ4SRWM62pFZ0
Z395AD6g0lJC+ze+ZmLMzPeIlYJouv7PItxYaEzMaSbE6rGj1/WIyMG5LBj/cJlq
P+KWpjpPVfNPPYIvghEemLaBg/TqF8W88LnQVPR5RdYebe8dUJ2+/aVVScPt9ix3
K2nrXycJMQ7IV52Dz5+BmZXtQlRWWcEQ3+3ingRJpM2ptrxSOt0WM9UliFfUgxmM
nKlQNK5OTKkyXTB8xDc8Sr+QRkuBGkqBDSUVl/EPPS6ys17UuNsHrZb0z+yaKPa7
7WJfoBbs08tjTjYuMwC2WdHwlQCW8OPsmJzd5ERf6iQ3AhExPDyVpSSD4f9AuzG8
WJpBUMqZkiOJCYvlzoYdgCzc24kyakIdpOsK/G3WtFqpB7awXLJDiWqP3h4ZUQq1
C6sNqLRbtzxI4HmpjpkMtt24Lo5ougMgjBkLrqu7IqoXAJA55UKE2fDM44AWpZgy
eGQfuuO0TlEfJfvFiBh/1IcdxY5nLTvdQ/cJrgdwz4SDH1GCjTZX6Gdy5/COcc3M
JjtsiVV7qck3fc6npxSnhtYa3mq/UXlNcYP0e2jzu4aKOcRgk1zJ6DYaz22hJEPK
Nnp7x2t5AUgJjxb9pOzBrcd16tT9biIGsF2tM8zO08Ou4n1bsoD8kOqRzFYAUdox
89UJQw1NJ95cnwG8u8UCt1WyyWsz04Hw+v4Uq37hSzaaF55qCqoGArogolZ2FqD+
Tz9d7etu2TIhjTFplK2Bop2oWSCwpxy61L7jJfQMifo4i1NqiG3zZBvbML7fAW4i
nnXECAhvIZt4xguaT39nIkTd/gitzZjt0J/LECkp5PVDx2V51O44D1f8MGsARrdV
7YHxs0LBP6oU14DA56HzmbLmPe0VaONwarDBQGdidBM7loaif8aKLhZ49WSLWz+o
wxq1J4s7pzOazzDTvSVtXd8AX91SzA/SnTxviLUEWQFaRKMUoX//dB/tmVFrREaj
fLcn1wVYXHh6vw8a0M3/mipCqfCIJpFO2RaNNVg7pfRC12WzijIUOPdW+VNYPP1x
ekRaTZpYIr8mZn4vayyc+EmuI285XBZhrDj1CbaBRKGd/aT9d+lX/fGbMvU+dgxB
9En4rLttVeCzdnTcQi3aeXfHAGlP+uT8s4+ViQyD/vMNEaa4bazavVPp8ixeWKYF
0q/1o2Wlcla/JSLMoMwt3o8hIHeaJnxDU9zmBGXPf48gejgurqQ5jKY9PSXtuy6x
NQcv120/hpfmp5WItqdn4S+vUAUYM5l89ue+NgidoBkXoq18AbYvf9etHc81Dsr8
CmQnOM8QDUeyCNuFa1KGgHs009Yh6kSGHpmvVDrx9EAkqwT364/f1E8PgZnblAIV
KHG3/Owwxgc7suXepvdrMn/buI+krzb1fQNLDNq8/lwS65mAhyRJBtHyswtOoPgB
AoEcpqgm5P0gmHOakftzHWZiOOtru3XyhIRjmnYthkaDaJhRCo579pxT8pmX+Ti6
pvYRP/gZcSvxxPoMYTdzGJpja0I/oczVHwXzXrTcclla7YsAz8WpyRbx7r48K2Gw
bJ3sDPSbRPjK1nBEsmIwNWunRIA2lty8T9lbdHntItF/ADPKMonoBCqS6WIG8l2G
36IOa2iml7p+n6P9Zq9yAJIKT6XzH55CUbc+hZJ8R0U1SqQWWQ2nqq3b/aQmaX+n
4+bjT+C7FC5yaMROXDFrfHcDwF63OX++F9iC3H+KsTlxIr69haCy9+fdc2obFiUK
sihr0TM/FN8xYan8nm9cjQQKCj4LVyIq56aqJ8dJ7E/daGrYBStWxio5Zh5Lz9X9
gTwwKE97btujiuKeQsuQT9f/gMmvnoRwctNJ7ZPOUZm5Vd2xss8dZRaLu5rI8OS2
voW0W00os0VIjgZLDzkw0iYD50Vq+eLaaZsZm7gXvb6itax3qhfzNrRaj3D8FsTc
rflH8qwrDJTwO2BVDMAT5aezeHPNdsKXuzwZAQ/muM2wn1ynZgHyvnJyaWGXpVrm
XyL4EQPfr8HfU2Cv8V0VDbIIjpl3EWEerhnXUXIyppF1cXedpEmjqA5lDfej2/E7
52xOp5QW7lvmvUS04y7K125PIOkyDxDGxBfxxafot/G+AFVwH6E0M5ilCnLwDRPd
6QYs2sebGWASDMwL5VBOER1HEAzxX1yPG4AOt2PDPjI0dFazV5LyqPW0b8W/Dcv6
OzE7aEX6CfbMngGB7gfHVe9jbhmO6/tw77smFjiN0wU/xP8gC9kNd/mYhdrFkn/m
UxcSgBUZE75bUqTIpXlD3BAFBxT2dO7euu7cGu7O47IS0Gffm5dZYQYSsXiqquhk
3B0N5d5IfNm962yQuOgg8EJqXEG4xaGHh6xWvGA/EmG8AjmLEOV5EV/i+nUvsSnJ
3oA76mq8c/qCODaIgNj1zrPFXY2Hp2+Fio12jkv0Uw4UaIFsPZotn5Gm/pw0cQsG
89Bew3rOAXLAJL7Sl9P8lSQLGGz8RY6bIdsrV4SE5O3av2iEKaRXJ3qqhM6jlb0V
Q+SBXvZp/HkcDsVYSWnJ3z1+b64cU53QYIT8otnGVjS9qjnDzn0/dPtPLgShBK2N
gWx0nZz6DpQ0uYR8xH1jjw9Muw9BMdd//Ik3ObikoJV8zGMIh5muh5ZxnemlPqB2
Mo6nPoaca70UeMhhx15/aVmh2U+we0BU2jvBYVwNOs4qj2AI69UpIKDNLLcUGBEA
pEsnjg38t7pudqjYxsoWUayDdhSOZzYJKimqiR7UtKSU1jfDWi7lVej+6N53tH9t
0Nx18p9+YzOzoWyYpHNGTZNCcRyLtFTVgF2bka2jr9cJBp+KybIUU/g10fZN3iGq
Zc0EWDfOiIs/odH9MjRGldrGWSbYgfFic2SgDu+rKibiYDHqRGJMstCNRAjB0imo
RV++6JnR+NL4OBgOFR8KMwO8LaPOjCw74js7IOlx96WPCylM8bwZwmz5d6H8IbMZ
Cj3GPxIWmqn7Vh6jluCCtopwCC48Qg8KRZSxVMAmDiaTj7rK0FZVWvpZlmhOO3v4
w8Ys4xTCks4QR3Wik02+LHF3MpQ0YQ+owRK33LCz9W81cvl5ybRGUCvvcNA4n1Yv
8Pz/bnSdmKKW97ieo8jJfnxs7bwqb2NAj+qRPnblUCZH0jMaLaJX9BRDFLU8N4oM
70NluGS7H6J20BxYDPDRy9gSninEukhoxKIl9OkR60l353kiBsj0hAzdQWE4Ukzr
IqsI5ri0sIG84JQkgt/xVKRsd9HZIQ0mmSMyiLh7/uM+iho5mEc2pMza0CqWj3p7
bD8ml2Q//qATtz5/FIStPhLxah/L5IlszZ0jxoqi+XN/pbFZpmWLdMe6nvoBlxYa
T1l5DaGdLSicfhjY10tp22dXKerOU0X2lFXuaAUiu4bzw82Th47awhG0ah1ImdoR
Bu7KXXn/J0RzPIzU6sVXdNAu463RZIAHURiH+RhZQBTSQi2iri7CgOQQMlgdF5p2
wbvH9Y9vm68JEPifDv3efRlj0sud/XGDpqN2A6PXy5lKZflsU0DStvHYGOMJAJYQ
GXO4iyZrd+5Pt28Z17DmuJKwd2rDkvUOFAu7BRMBSL1u2tR5t6Pr+W+vV4HsMTlo
SVJxLrY00WSeZboNzGULhqmH0s3f+sXnbIjvOhTZz7awWa5eYiMGBI6c9VmS8sH1
D31AQnG75nvG/ImYDIcivEY/9RkRsqq7ZpKMvWRLXaVNKELz6hxmoWXACwzy5ZMk
7aNl7842wGlE+FuqPdW6DEYa0WJHVnog8I6oXPvZs2O7RyiYMGsbXB+Sdhh8jqzQ
ZvVCfEZilnWYC/Z9JigSjQhm20rqB/P9HtsqKe2iWmacaY+A+f1QUFfMtPnTYoka
ZWcvKLN4qPKqNBVOnJIukvU/AOVX0HIr6wSWoWAMqJYWMQ+tCB5fVlk7v9f/+QsP
A4ebXcjd0Zt5/lvdkupWy8qXkTU3yAwGZMv6gtItvXo9+w787GX5jBk5HrcHtF9N
2qXOzpO5X7rX0yjtStOQbuciZEyOD1rJxRX+kxMXP04NRyzfQ5DB2koMseigMi2o
RR0RgSM6aq+za2tJ3AYfWA1XxEFSROl5FGTqmnOxVeJ8GuB1mZY6kYaO6QsYXb1i
6++rxwMogZ0kdvDZ8i0XrDzRRTBCJMaNsCadFOfiOP+wNkjdhNWFOzPX5z5B0n4V
2etROy20th9zuMPO/0/3vRp4q+rZWyoGMnDNfwvM9mL/MdiFRoJLv6OetFxNdKtL
h/DI9GfomrRiYiiQVh6iWOnXPpfTHhIZPh2r06ORMpDjj+luxVLjRUSRRzcK0Kww
6yWXsIuEw/M/ICbUP+uFkeXXxtCVA+nWxDgxDkuemxet8DWNM0Fy3bjGvI8jRSDj
1eF8+yh95hTqIkZ+fQ3dGIx+AqbvHq2nyE+vkD4sZntpICkQ9CYj5Fbw7SZL+7De
2otJnSej28H66ST+xPzhGuR/uGatY7ZDbXe7clx4LYr2MkheuBlxciEqQf+IWkg9
Cya9JHsChr72CLjPXnWeoBZFzPKsEuZcEcKv0UgNrr6NIGi1v86/647Fb2901zks
y6MSkpESkcYn6/PPHKBIMSFH0O5rHidrNpVco52NMBxMniHBkH7JYDR0neypRvPi
oyllX7aJD6DMXKHwKgSFsfhoM6C/GLe9IOZ+UXeSCivCArDrrEr8z88uZWukIOCp
l9Zz6EWXAW2AZTS9WwmH1//Vp9PUX2TnOc6+VD3cCtlo3dwtplsqY0G/HdbqolLE
UcKAppnYtIoMmLFzLpCsdK6sZn7cPuLcJPonZ5YPiG35h3goQVOF2z8Fv3GLV5ny
nBVTRS9t7GXA7zISiPmNqGA7Re318qd0R7ErhClGPfyIPsQZNtYI7BGSKtRqXGEb
VDIegALtt7m2hf9CvOtIBqZzKtsgTcMiE9tpvY3BGc1fTxnxEeynU/1RyNExq2fz
Dz+gDaLOnO6NKT4CjjTHl6upx3rgxQkIApGgBOaWxYLEiqGuhlS/4GOXUS5uFv2V
ZMRArTgmne1a882BxzIdE9itJAOEazmlSI05OU4Sa9TwGP+jEPcQx05rgE0aOyxH
Bpaw8OIAtfzPew2UcJ8iG5jZGFR1r6/c9UYWCjbG94dNdQ9v+iVt64xtKjzTVwYB
knt0PZdixz4fFmoiTMCb0Q2CTGxYfHNnjqHwUL9cn5mP/4geJP1s23XbgHLOkK2P
UEbsGJcctJmT8ceY1QVOLy2EQADjI8eER4S9p24fYs1ExymYpm0hNgwcNsDIlPTW
VSA4fw9t5Z138NJmRgRkMv+0JK81QFeMsEy2RRKEEdh2mvv70Kf51bKZBMB3zcfg
A1x8895e/jCXseSkzEtw8sGiKYYrSaQUU2Dffd7X/iJPVUAus7Q5/AmcZKk06PrT
Xj9XFtil+GJrxULIXrmcy7QrJhh/y4DeWncFyj7ztdGJ7UGiJfEEAOzQBJ5Ue8uj
zO6EJNth0OjLv4BCDYcvfgz2ccLFPhZvDk+oyuWxDAZY03Clb626H0dVPajjDRVD
WAZ74XNyJSqwhNDDoPwuh8pMKlp6UPBGzDt5YcHwMVTZjvLCoN9Bstp0Md3VSrIQ
DQ/3kF4wG9QahaqP7t7xkPa9ep20juYJBoRA0c7IvaXyf9zAdBh6YnIxJ2AhCDsu
CmYUVpumgV1KD4ujz+L0bS3jxm15Cq5M1jiDXzYRq7zCx095RylXe2Uo9+6nJFVc
vsPkPQRaiW7l/MP33smNKDJ1RidM08jKZii/pz56t/yKHdDQuqrQ+8wJiEOs8Csk
eRkpNq2o3EauSFPFW1azRMmEAnuQbBi+opVmlsvc1TpPdIp3rM7uwS/GPpy01GmB
iy+BAAyasE961R/iXk+36tkNJ0jI96lfb0NNacJwf/PGOcjMo2xFTCyTe1Ck7YS1
t9yqG8OP/ArrSbXG7WTlV24dlQxqB3mksQgugPrYwwhsSwMRWi0Gd+CkgeTC4WGn
lcY9DkcK3lz0YkBSu720qGbMK/i2LqWS2EKKGKAqjqEqfRIpCnqegKvckrP5Ldur
sg+OXI6m26lFLk+ERRpbzrhGxeXc075Bu7FTo1aVVAzigGp80ses2RoLvRcAhI9c
5zYdiUYk2Psl62nRl6bGeUvhmBu+fovm0LATtv1cDVyPaiufvIZi3/WOBwoG4DD+
vpU2eIo7y7MtDOCSOAfOn5GOuSXpRpgKyYT4mCgo0I3GYfxqmhFT6GQOnXx2F7dt
v7+bkf89lXtratpI/kzM3TDN8ew7SikCIH6SFgwt+DC2xUUkWKcaJeof/uKJW4pb
ekVL/LyIl6nfb9KlVC7KO+LhmKe9NbNO+GmFhMYCy3sP/Es8Zj2UqK/3h9gH09iL
MARc8QJaMeU6ji2RVp+ikqbB7NxGuS1skwwOci8aQ2UM7pw7JDR1N4+r2BZNZDjQ
UvOwUsNf3vIy6G2oflMRBHGExpiiJhaKygqITC12DxloBTboJJiUG8DVEGLHSH89
69F4IJ8vD46CNAoigA9YZFaUzmT15Mn5cW9NytWmTSFkuoqsthu89s78H1ykND0y
Lr5yPFWWnDSbYJWF36rhf1KwoOpqW1qjmPIH77uwJ22AHX6fWFQ145lVsWD/EjGl
iz5lrCvP6yWCYbmbHsM/sgx94TVOlofiMWHhcCfOV5RogQbaeQ8MRRFPTfllBP3c
u2U/MnheMe+xR4fj/5X+wd4dFs8ZcYzhBunUstpe+7BxwBg8Cx+hp0gpdbYrlU2m
9i6lUginow/JPhNfX9CY1JaLpvUw/JiLMx7A5dBmeKGRY/8dAAnFH6K0e9PIIFXF
bHlCuNV5DH7bTb3yyra5vCfHZq3BnwnQKxbGvrxzkC5l1Dejk07Bx+lPXLtXTz5P
yPNr/wjQmPTnzU7D8h2fnDhRChCgE4+j4pcmYo0z69IlQBFNA/ZHwFy5LExbvfzR
NyCx1pYu8mnBlciAbgcvEQEz0hSEZWxyMmUwWp9oQXSR87UnzipyJPfowosA8g7e
bo7YivUgGLTbV0H7cqYXT/RF6IQUWOr6gMP93AMpy0XKRY6u/umIrcZjrs+3qa4N
xQH9ilsGxsTBdOzTgkCLaPW2gmjiV2ySY8GSAZGxHJy2BOtOhwwIOcC2nONUDUfl
RzsSbn0ZKIdPvUPx9Y5IiW1A/vUb96kcz7fv4q//tavMGqND9LpFB3WzOu3y8Ybn
Q/bKPw6X4QQbAXyJK+4LQKuwqhtGrVc4Pjd++Njv8Tdnve4INyFFvrs0yVuVMS0M
N0pMJRf8Xe+3TTs/yDnpGoC5tsaCzwcQU2anv+sorIxoRm3A/EpIPM7GBHsqQWxO
pvLefN0vKZJEPZW9lBAh1QRGtS4vWZU9wQ/o/CZ/uvbHonZjW2OpDgh00ZajgwGQ
uTRrXYjy4Im2Ry7t47jjVNSi92k4CfTvH6flJ3tO9UdeJ+GwK4Sh6wD4VP1ZHLZG
xF1MT/feMdu7+dOeLWPsnoD+HC7HTYuj6rt4K6w4/klSxJZGnTh/e9VsBLYnyEZw
yXMl6iExjEcOG2sZw3uNIk1CuSmtCH5NNtN1b4qgfPxeFTOVL2vt5/5H35Ac0ks5
kmDc5w9pG1BDzgskpw7rwcirfulNAU97gB+zJeCSSULe0Pw4IJMqUVbZTYY72GLQ
DX4ctcolJ2eB+2StJb/TAtlNZcjvUErjUv8alwpbHZEcIohAvUh8KoBMrCdFsFB5
Nh3njRL/d56ytEdoHAeHC04aZdcMAHDqt20N00WXicCtDfPJlV7iQuUDgT6ZFetY
hpgRCpnO1C8D+8xjcd7zCZhdoFayGRIVmM0VGq+kL823f1pOdr5jZ9mwI+CnqmlX
SK1q2TigsxFjZGv/pdgj8We8E1nugmo+yMI3tDMA7m3jB8/Z3RGcLmCZSU7CwHBn
C3MnjPsBAxc971aAlMX/KEDqkFYHY1J1QsnQ4XFFKXkIE68cflHKZPSlJT/xVsxJ
cL4dOqruQlb0U1yES2B3x+RWsGy4Tty62it442QavhxR5VAQYzTSt0v0FIRh66qH
OHP/6X2MwcO2klHCDsRUyXzvRfCHqkVkF/WlYp1QVU8Kk5cJ+ZX7qb9nmEBmkUZn
CbsVplLev5c/Ab+73KXCmr8Gtx50aMYF831UQxxGOeT+qf4YAm/4JsWW0irW2CGD
sVB9FvtsN9wgdea72oITlO3oLm5E1WXjiIpsAkEK8PNNSNfIqLQ16Fir2uTmdOy/
NpzuiFeSSPNP3OVhEZZvbm9PAll9WERcHZqlfWc8hj3C6orRXUgxSPhsQqm0x5qJ
UZCCY7a1eBK67yDU2wROu6brin2LdNgeufdMzBgaI3EaKoZxjyRCRFltYYtWqxmD
ghEhoPCj4+Hlf0DBmxv0RadCmRuBethPX/1OLg8SbeqSyUS+86DrR+081DEURiZ1
fUc0idqOwc4Wp/NyzdSGvY9SPSK107Xfgh/aCW7DoLykGaj/ZuhENjqCdas7KenO
Q4Z4iBpR2KtQdGk9ghVOg9P2wWlTSz9ETFluiaWwDD4mtrZ15ifl/7EnwswcSohk
6iZ6gejVzQbnDOmxbhwrFoVXqtXx2hfjbJSZPW+6jh1GigxYlXwvliS/g2P8m1+u
/lOX5JAz3ZXyRkeSiCpqpXAP8aiztHj8FK/qFSyA72M5f//KRFMltuAxbgARrPLO
B9QQn0ZT/j9xChjka6SvDXTkoKq4JbbSXg2DnnU13aDLRfbekWSBgLS7QoX6tPh/
EPwYRadjkZ+7tMd8LX+HqB10SW45Ce/kD3DcdE4vWTUKB8w1lD/hlMh3/LpW/3df
fdd3jzuUfkX/viGrntNA7b+UzYAsaDu1Gw5q2YVqEBfonxzXFIcxQLHPQW9/zhZK
gLZQ12PX4xRewU5VdoBgcHLskZjt5OjSUgtPamsMnG2bP8XVwaatf+tFISOWyDxO
JASTP1BlaBpiBnzLkP2Kbx6PUXikvNK4xSyjGbPuoBHfvVndVi02HbfHNkctKaOP
Ghj63Lk5O1OX886VgscdqZ6tpKlTz8bv8TDr6Eh8C9gpAAxYXBpbSp5vng3lZ2sS
OmIMJ6VAio591Ij3IWNxvmpiwvVZ4oMmDDLxrVxso9Zp0o9jltY5SXEK4Ujy4te1
ggX/YVKG9zyV0km6SX9xsA9NyQ+3KWL32kD/cBydrTmnLQ2F4a1wQ11ZJid9DCnH
a5w58jpA5LWupL5ZISgfWlFH1Bz40Hg6pJejC1cfFNVUN364xDuHS/MnhRE4OYX8
n8d6JwkRJtoR7t4wxPwEV+d/fDX7Wub1o9gkiCPTuiG1g8PXTUwXlhIXiEyUoIF9
j/kaRVfmddnukq4Aaf+1tbdX6cQlvfpoeNYxuR4eE1JTx178tD57nNMxgXQ0iIkY
zZsgVvLeUbcOuZCJFyddr8xEUv1cLMyJMp9aLqcZlpDYi8dvyJ2lLFMZrVSVpMDG
j10ioNBRpmcYr2xv4xHHbIuBcHEX3Pl3wVhaW3G7/79VP2ilxdLOYqO3ukhIuYdE
ZGk1g8bI1G94mOmPuQsui5kCrcF6pFVYF3WsAsQIMggIrcchqXsC8v7XzKz+DWtV
OIshXWMcZeD8JPUHyzQA+sed+jiTQxwjPUo7vEXvOCeb7HyaoXaBg/dHa5bb3bHT
nF11NYr6D2JQVzcKZg61XFzb8cjz6u9NL77bmSyAxlGXMZKUJ3ZcxpIFFn9tCmpN
1m88Mw2RMtu/xi+9j1AXQQg05JSwihVjUsCFlbBp3P78Z8dhwEZAHKPnRX6IOgge
mzM6ozW2rA7qH7YNTayDcZTUc/OH+15ekJG0D5uA8XqxD8BwzMtWlSkmRleZVYJO
1notCV+XLt4ku4goDAYjDgjcACYy1UTBHiaFPNuEMNEkCYj6TVIqz3ZU05qVEnEB
7CN9j6F5oyhJ0YCTz05TtDXPm6KNPmdIGf+nmNScW30hn+pvG17jAt57WFqZ35ge
jWg8KXlPb16bhi9mxo4udtOj7vKAu1n0yWHHI3gak+65dNBE04ne5mkvNvzuS3a+
rawFMVb83gQDS8MN6uGDnJYJrdzJ3Jkz5vqziZ23/ANnFwyfUhRk8vOX5ONnwI5+
CnTrMZlFjJ3MEV4cykgRBnSHDp8WZ8B4qgQEraDApApu3815j60pk11QjaYIk28O
z5jqyEEVTlYe/HlB2ad/OY2vIGWkvM8t+h0IRn+LW4W5t9K51GQ/TcQPiQnXwyJO
uixxhfbzxdrc/rV7yX6HOjnzUfvDlUOv6vW5GChuQS72coKyOVNuWd/WNgzn/cVm
R0p8lOab9YboTnBJFEchlPmLkQoUqt/Unq3jJmeMS9iMx2FHWC4QsfhE2Iv0+NCW
aYhRaDU2uxKleM9nDlkgbMjNa773t5Tk6T740PaSCif4rSHjYwJuWBfGc+nCvYSH
yxRTEwN4YcRRdNis5NvgTFU/100UUwQIuJrd9Sw/guP1tl3i4sQ8uiws8kAiZas4
6XTz79vna+b44dw5OeS2xYLi9HPZzxt7SvmvyRBhLo+YAKSoT4a89jcReZtIpnQE
6qZewuz1DeR2x1bwaQv6EwNX9jYLLpM5SmX7w4IPfvnCPjTObSCCakq+3Y8XSLHX
65xAXnP/W3hKszql9f47V39WvdN/15PLr6i+I+UHPOzhCf6UT2BH/mfU/kbJPr65
ZNMKkwZHFueztKY6SMaLWV9hMISlQBdISOW0LgfkK4kbBXaRI0AiBkKN6J6LATSE
zh66GxyYzkPUkIcrWY/TP60IKsxNnNXrM8bTU2Ow3hx9x2XOoNLeHa2eomLhLeB8
f3xr95FXGIYXsvfHotVGIb+G1/hDCgx2vNaG+56VWfnIntVf4i71SqbgYqlZ1d5b
ZAfWUGsPiGnJkojbHtg2aasovXDXtM+dCnb2z07mE9Ccdc58Ot4gpVxptgwwXxtB
F6zfu8JIhEZvCwWWe/pMMJsXafyofRzKbXLQtoObh7pU+Lf9rWCVAQJmaIxFY6tc
qK8UssM3wtNIIbEO2QrS7/x36j8/4xNsyWrICAt/BLxfgGgw6jmAQK9XDDuA8bSr
In03Ob5kIewCqrklfMdrT7S0jDealTaJrhB+qavcZd8WAKO35bMF74Oj/M6vTQGk
E3svwMwsG7Jua9gACB6yhMC08ztiC9HJH1TAoryqbs9S6FDirlF6k9DOMvgpu6im
6dvcfR1n+jItYYGOdcDZr503aiYPV/d2BjgMphwLtZHNG32ICvWB1pfJSKbyTY5s
UVhgmU6uaj6GIAWY5DaKxYRyRbQ+iEtvOqgLraKEQiTGtbLmvFjbNA0Xn9NKsjXs
9jJmwJySzN/zf1YmaBhODqZy5GJFv76Bc6omRpzhPDHFrciVSIaLmd+5ud6Oeez+
s0p+U0BWy/fLTbut83mxocle11xZEAWvM7vLTXwIkqB1stpl0cODnt0OzuRn8wyS
iHJuL8LquMcKNG9epIziLs7GXOlEFrUHEigU0fbeYAO4WZbIdE5HavVyjWwmsgrO
Jl25pvj6All2O9EE9xEoIdVhDqoXZi3ghy1P7l/Djg6nnXxIP+wtFL+v+Rrgad82
W6f8ou+YbKLj8bhdNUMidzP4E5/ES3Guyz6Pq47nIOo+Cibyf5Yn2582E8mUZAdU
XSHzZYk3B3+Y+8od4HBN50hSZBMTmYLZDKUsI4B7zIeI6l9MsuOupbXWE4PP7XyC
DXRKEH1w8TgvBt0S3vCLHOAUCrS8IunUuypW/4GNDHHPH1sEkjPdaz4qeFquK0LU
9VUYkoH+fp7l5AnwQJokJCzUtX87WCoBR7UkTuIYmKAOjfx0rKZLSHLtX6eo3O0F
3R0lLLh5qumuT6+22H/02oxjGoqTuqo4NDQktuh9oxHpmZHdv2cNxLN5SWy11WtK
3m36ddwsN14iOpbsGeP49NA0QxpHEg1AN+xTQ6DkUAdZW6ad3RYxaTCnmvYso+oT
KK0kzmxOA92jR7tq0ko94a6bExob0cuJQJSnxGh+LCyGq1prWVWqXxo807QvAMs6
qj3cJ4bTRDT9CYQ5Qp76CGDxGh4fI8pKEeMoXpRibdepwkIjhdfNevoHrB9O6kkZ
d5qYUyr86aiLqzMGMzCSsehtBbTMu4jBJbwDCAV/3Rk69k2B+I2c169e8lFuUeH8
C8W+WcYry5L3T5nhBlR/N4CRbnSutcY7ef1UgWjV0Rg2I7v9HW90YE4AhqIYjHDV
9gm1Uq6qTq8r4TDZ3SIIaxlbwArQtt2my1idHdvotKbq4LzT0+nqg6EC4ttB5Rpd
bUFN6vh6zTO0/q8U5uhP4U2vrcZGdk80mCgsnc1OvMTR8MBSAXQk8jj86bnx9aDq
zPhFFuOV63ozelb8opzTEEWLAtjH57sloBRGdgbeBCu0ClFaoboM7P3jt81OwSTK
JAE4rg7OyxjOHyrKIpnm5/5QWckzPBHqG/aA2OV6NGrp3gtnBEuk3DZLYvSWQqoX
zvo9Zohmc0vnHXGQ8RlkYCeeK9XHHP4QEV576CyGbTt7TlfLcRCs+H+5fRjeXGWK
2rMYN7txLjCWQedsEWN3sT2w1OcWTc3i7rdEx14w0pO5L7ZfUIouqtgwdqVI7wFL
h7bl9TkRYws86rA2m50vdye7h+lMZu/F9nTdP5uneE3pZopt07/QaAJS5lBWnSBp
ppUEr/7UnokGjErNFg4mV8T3StPM3EfPFopHrOE5FV1BGHPzHdViraascytCk/XH
9S38QPRXzpUHZOuQOApvr5aVjf+nz6Zr1iU32pFnpeVo+0wbp2/erpUhVQ3T9/2E
m8s7ITJxc2RlUsqPTwxBQqy1tywUx2xXdLM1x4P+vdc8LKFjgHhqOKMbVDQuXaUa
kU8mWUtyt3GQRSZRcgnsOd3jzz6ewaNSm0YW+I7WooqhcpppNMHkfvfo5KzmKoyJ
tW0yQemkBOqJL5x3MC0ruz3BH6Q6kA4iTfDRfOKDDPKZmJrOS9SPyPexFeemYfdr
+BnvOuYOY947nBm1EwWv2TnSWTixgBa/IYQTeGxycrh1WYCBTzJtjJEvZPiO0SBV
EFUUA/++D5dRxwVCDvsHD80YZBBv2Tk6OjtfTtNHN9da1yYgxFS3pZmqOhWx0dw5
CSPs+b2riUTyL0WPl1bTxJ8afbEW2OeMw9D7Y7Ju1cMvJyh6PSeqzWTCtliMxXqB
ieZQQhtFLEdDRQpantYK/Az4EAp05GcYLRC7RA3f2SKpNk4iap2s6yHvMMqMjuE7
obU3n8jEr7evlQh8WpfVjECohRg7nP8zqPPZGhz4QHTaAcKHLeBHbsSyAVgvGBX0
0D6HV0u5Fj8c+GB5+BruRU7z8HR5BqppscOdd36Yl9GkapMHIKtxmSTGvJ8Felnp
2C1wTeiNNsJyfMIDx0qYR47WXK988klt/Vfy9pLmRwH9D2X0oR3O9HUyR+Uo2ajO
CzFWSYa2qHh5+I6O83m4xKpveoX/gDnGaFp0xVwJSRJJMrbeI6bjyv5GHyjSwRAY
74pzlPcCy7Hmr6f3ZuJfb1BU4DnrLQOUkcbdDKG3jOEwgvyceKEmGLLhIiqQVHXw
kCPv7+LccADWxSALbmKRyPZWSBdgGnIyNst8j5kDko5UWdUHX5188W87NawenHaq
MnriVw9b/jFotmVALhG8eG337x9ne64pI2OfvXQfDZg7+uOg2YSpP5i4MA5AURcH
BQEZjBiHg7DjZehEINuQ2JasmclLaqMNlzeWQSAZ6xtJ2Fv6Ymw8JUKKKbQQt8Xs
oOvIFVNnKo1ZAzk1oNv/z4MdFqnuAsp2KK6pORhdFsfCVz6U6nkN8jOsZNZjAPZf
lpim/AzhDXdqrK7H0WcgjwO6zxV5c2onGZySvLy9s0m6CzCkT484AkB0L6PjtkNg
H7tr978wyw8DEouZant59mJDMwC87fp8X000W/tu8re0UEnK8NvaAbELhdIZ+Irs
X3eJi3cG082ZC0sF/h8UIQkEYNuEKJfHzA8ja5wsCJJ9Vlf9X/p1fX1o5kOKZM1c
hrQW2+Aj9tCM3rF6BlR9MBjksgi+NUxOdnn9VxI3PWZuIyzfTnDRpBw1iarlyFDl
1hDpntQZTq01BKTTtKA2T+KkgSO5h9uP43X/x7Zqnp4Ci/iHdbGlySLgk2ICGD3K
haZigRl61B5EeMxlIy4TPfIpPCp8+ycmBhPn1k/czwAjw3k6X8zsMT0LiffM0oti
8iPkVsqvQKVpI/OOnHo6yvEKp+it+u3bTKcfVIBODcg8l4hKHEwcjnLj2H3KNuD2
m8lJBVQNTHUJbAYWaGGl4ZPjbAeh+n4ufaF/8t+FyqwJiYAW3Uc9U6er+gyFuK3O
MFNzX7z5wYGIsojPCHDXyw4XWR8fwvNuI2cW5DVvhY5Kr57BJHAhmNhJgZqyLeuU
hR2W1sOSnGh4uJ2gepPXtDg2qv2pGt0gICantxqjjhOKzOwZqh584/aTz/HwYjzH
q8W8vJapOBpDl+lGdVqGWuzTFvcxTR1aWjGfZAahg0kPEGozo1wwKrkEDlAibx2g
IPD6JWJFAFIUP0twhlZxJsIUX5+F2lzivgg1ThSkL0ubbBu5Yswuo7d916uc5y0p
8uMtVGhZYMaDozucOEpAyHETm34zIZnf9sxrzqSVH6Kkf/J+Muqfu1212A5BPt2U
xTf4jT7KG/90xludnuLi3/gEw5YUTHRs+B/cewepUK+M2Ol/XzyfM/QHgvHRTG4E
jEy1Nfd4lBZ+HVV88xBeZDyYk60YHEWfb3i2ASe1wmeo+Du/p0GWTzhwcMANpb12
w5Fm5pV+TLeqRC+09tFz5XK3HrEUZKMaMhFvLBZuNENlRCi+wYqUKG4z3c0ywEzT
/bj2a6YjJ0iSHP/tI8bF6qm6AEQxUKZ9jim9fzxFDsunE3ZzS9C6PtqufMOVMAvw
1dyJdwdJmBAoXe3yhaAdUXACidc4ujfdi5peqEbU7jaRudZdpZj1Wu/eIFIF/q7P
aqFZVvA21c0isEPBUreKlNX1SpcX6ge3xGpXNYiPP2fR6xzZD1emgN8EBrGSZUQy
wAP1SX2i3DmepWa4rhuj1hVad0jHCbHQ2U8acSVJneegwAR20e09d3Z5Nyse//K1
anD30PMqIFywVrTk8ShVBds/NY/6UDB7Jll3meyVWBHZc9KTKiiDS0pTTAA22LKz
YYQGikEOeK4lhc2kYogs2miza45dhE02Ls9Ot0cetEqhLL/vswX5XIeEwQxCVNrI
8mVsCIbYzd9grp9Cc/eZ4FDICs8dTkNe/sc2t94xjS9ItG7/uTgyloWAQWlmkGvZ
4FJpzjDsEkBAm8f1LryjemTjkmVR1HojO1sTZumQGUAGK+NQcQ9dCGoXu1jXmlVj
WrmxA5OkKwPJqaB4/GLuZtPiZANRUR1Yj3mOaZMQdCiNqhH/mihaE6FWZhNkShZA
avTo2s3aej6pgJ/4sWu7X2lgSAKdGH2ahi+cbAJuVOjGuVn+6Vtpn+w0Q5gmPMk/
37j/SJHY5EnXvgEwiPYDOnHf0nKKwD6vrzZ9QnxysYKpKuFEJOs0VBx71w/WfjNE
0Yfd7Pr9tFHHil0a8MJFieyt96Om1dGOPIosbzvXjGN51jSueekdVLZ74qtjKXFL
LR9ED9cHPR5eb4nBDusX4QaFdjsjInQBXScPOn16oKRx0DT5KVjJfwKdi8KOAs+k
Hush8eNOTDGGKqqZFfcOGMS7CKeM2+hBxhgtc2rHqBOPJqN1JYAkPPXNNRuj4dy8
rqdZJ0XhpPH/rsS5RxW/aUPq48pV4rIyEbdgZhA9dubOfRBvNJxFNXEbZ/fdc0C1
8Hwk7BqYgoGPDQSOt7SkSiV9VpqrRDy7wPSXQ5aTiB3HdC0TAG4fsgw5LiGuH6/Q
5kRECAUMaUV4ACFcTXxbmgcQHtWMg2H2lbWGOXEllrQVKWPDlcwZAU3fle3YRC33
HkziVgcS/YasTToodQEg3PZfeY+3Er+Gl6QuKeUhYhOO7wF8D/GM85LZ9a8YmoFF
dZ2/nq+2eugpbp0zkfndyUBXoVqheWoeaTEEKlBMtEgPy169hRDfDIIg1LBLmk7+
YzPsAItE5jQtBD33tYrVXpD5wb4paMTMYeiwzAGIv6L8JnMFPTACQs3Mvp+6PJl0
JD4M7BWmPUpgUUKQySg0t0wvKbbb43Q/0FMa+eBvAUGGXk39Hj+zgtnIQtd/RPO6
0lw851W2qae6zgHLmWTY4Wzu6TEn/7zFjBA++8nnx6nwfKUpkMCuXmnz7yu/Z1bT
WeyEhWL7rWrOCzbb+OlJJ1yZ3hgMbA2lw8WF/xhqiIErCE448+4IdY6GvonKyksy
lsK1IqX2B7SR3jIOjgXbyHbYRClaPlDmgegcp8a4CDOLi9QR5JNOSZLGge1B103I
s+HfW4YWaXbv4mjeqSAVqcCo2VIuzSLX9sSCzL6n24YcCBbbS+Lkayu/OUgS29SJ
0XYaYQ9G74MhJkt6+kTJQ6bV0VPcANNCU+zg4ZarvF/fb13S7aPHyziEQt2url6J
nGdFmjjMON25soJPhQLoNX3CyuIuoETXNPAUFPbFlJuFbSa8OomkBwCQYBehH73i
5Svx92C+0HtA5GdBxUdh0Pk9qe95JvqdN9UizSCbBPAQBt2n5jx9htwf/mnuPaKP
QSc3EENngRgBVaU0Q3T76TxU9SwEFK12pLspSdUmbmNwGYyTb+YNH+2Mg+DJUFvu
C4Zz++T47/yyKloBWw1bSJeki8uy2tzzx0AmDeV+gu3UGCFIUH0q8KbSv5Br/T5o
CAwMaC6dJyQvObWdjV+ubkpRPkMOpb00snPqTEUb2iBhWFvXg99cTiwqN+m4/Zzq
hnxWs0FikDk7nh5EciXnNs2GfMuBS7VajVaYJyMovaXx9R4t4PSqiJNjUoUBOzh+
EpDRv1ngG7Dl02thKZdwSgtQaaRqh+PTH6+Ea6ApHgNCO7vPQdaQBmD8FJZ2UYLW
VRUKleq8hjQXdnFupeNvWjCA4GJ7g6lgPpi7cLISjK76dd7O0FgxiBSUwRIVbWsb
0ckUr/G+4UKHlMQ3R5hrf/HhXJcUkeYF3Q3qZIl2YQ+Afu6R+h1PLbKZeHJs3b1d
V9ZzPfcUNQy6OzzQKbHAgTgHdh9ZDaelvf3pl/r+I1e6oABHWOk2K6SiGw0YpLgT
mgbevhBiDfVQl72JjOCNyKxGJZKD36MhCNSqs0Tjl0EHAajzp/Vq9xvSvS9HzaBz
i+geXDN8LojNZAXDbdtyFmxvJpYaRXvnT3M3hMtyqyMcH6rPxJD8XCLxcp9EXrHX
ahqYfUtqPQRHCocvEQuz6qMnGs2Od63Yc6BzUdrepYCHFqGGB/RCsqHZIOkjYWOF
qSGvenGNU279TpDx4eHy3zRPr7o9oam+6xA+QnWBUSN8G4xCHNaK40t+jJG7Yhgr
cxauwTzmYW+b/YaKfvFqnC1rVs4HZlD97A0l7VIbm2ELvg9F+uHCoSheUh7WhFp2
GuMp4nAnM1hsXCChlORvPsGOkfwBIncy25PqFJbQadkx6kWZPjM1JZPS7YESHIZB
AG807BGFlqO2CPoeClAaOgMxP2m0TKN9GPI8/DDoS0soupa+FSk+7wH+qFKXqiwV
wl11MbDaazx1GQQNCB54SnkG4wJglirRJLeamm8c3vyxxS/18PR7Ps5jfnOt9pcW
8PhbY/atrFWZbwKHOF6f4J/z2rei46gO2lJ0cGrSo5wsMdO44hM+uoj26wcVo2/p
AMeRcH0zdc5+6pG0aotTj0k+xpRZYh+TGNfINlqbsm6YJtVElyEeMPrMkf64IEWT
8MhK8e9YNd7KkSWa9RiY0GvMZXjgmXHzI70meOyibt8C/zp8xXaF/rBb27f1JiJn
D6+2L0JVBD/YkDk1q8NVbQ4PHMpVLJvoLtU9hReJP+hXtY2xOfqMualxxhCrh0l8
aqzBVPDkV131qPHo7HuX8IF5x8TcdcNfmsjO2WoSgTUMmLEI6kWiFr67Kbyf4hW4
WEgHEzvnXVaVKkKXb2nQ6f1lVGDIK6Ze1WIoNB4gweOLGbxNR4y5QykCCKvutTug
pnYbyteFMywXhQPC54E6NUYeaLQAFRluR1Ge5E0WR2gBIH5kRZ3drseM6+ZdGKrq
Ft2TZySzyFpqDsHCGKPWqPgebuASlpdXf7TTogoliRPkKsPxgAjOY2uPO9U60DBE
+iBFlPeZDckzzNih0l1W7HMxcO7XwO5yVciXBDTE817rKCvhgu5FGAf/ZnM8vmW7
6Nv1JLM12VDdbZRJTiNBZkVGdNQDVkL1eohTJ++BjDZB0ieMdVveAzImyPpH0hLY
kD9RweNaf9F74kNLPiu0ld4J0qCnFevmP1trahdB9FlXdfJKJ3CH3acbUNxNC2ry
yxwXBIhi9b51lvXGQLCPkoPIz9INQIG6K4WlH/gHkRNB/GJl9YTgYE50Htz6ma3+
oCi7Ku0cqwpffCwq6/dy+XsDxEwqyu5BfZMfDIyutOJgDMC60ctDXBa1jwSIczlN
iwfY/F8WlaTNEAkjuAum+5tz9X++Kj4AKx42c/u+bAb27WIq4DAHTvMmVlrQWPqu
79LrN/SEK0I3je961CYyCwOxmk6PJg4IG26Ygi1KXkMeBwdWWHyHpMrxocTnztpg
2U3JnLsmmEQrL1MS6Wk08PInxv5GeHdzyln5U7FC4t27r5HC62ZCh/Wfx4BO92W7
v6Oub7Lv+0psJKWVbcY0zS+H4Gbqs5bxRVDBQCjz8EncdBoIE/Vwo2ZKg2HWuFrI
LjOeTQZVKVu+utp/HDtznx36HeDY5bjkHSa3PMJyA/DfsHDr5nhedvWUS8wCpH11
NpIaN19kyftdBv3j1lTPdiPGWChvX9GSteUF6yFRiwej55pDZF8JTCBs/XMCXxL7
ucbcfoRscjjIe8jdnVbf19AT2n8+haSPyUmpYYygBD+1qpQdtzn7/1T+iWW58mkh
XLCF3ySDF1J5sO/AXtPo+p0IJ0lcnk4OO8Dff5RwGH4SFH3rGMTUX2lqp0Jehv3E
C54GaSJAALkjzUjZjsJrL+SofKb3zid+hrPTlBE0C4EotvvczVlGG+uPtQFsZqdQ
iTX+CPjIdtMwLVlWze80NJRL56S3rZc6IRdGB8HsDHTU+toinvfPz2SOhm0TxR+b
5LEFgkm988V9NlaanI1CZOypTZI3PVAdo5sdhcKbNTuYhmZhwToJ17F9sKGRwFp0
8P9ja4W02YvqNsV0KTpOF/KH4ZVKZZme/olgS11yA6QOjhkXtQP2004/cfuxJVPX
bw6JgW63ww6mV8rlqCJJkZsMSBhhzqhKYHlqPN/8xTY1ggegYz1/H4MdWmiUxdmE
k4umH26GrcQI37cRGDbVjyJUXDV7f/4egr2f+BO2el0t3COKVOLn5uL7LE899A64
FrnhbBVd5mdVgARh/1WpiK1FeTDPa9RMmC4ymqMXHpWdh/Qc/hU3/faABEOKPMgE
PYyjyat2+Skhb1DSZ57kTNeqSAbZEvMYoEoOkKNgKHjQpwE1zgMLlNE4OYl2WmQ4
wcWoBDhV2BGfYb021kwofoUv20HmQwX9jBEdPFq2/dg07+7qNIqp00ond2kaEkO4
uz4pXsBbOic6Zk/EgU0YBAkLhFAHjPCcBEq/q07/TdIEzGRuvogjCDv7wHMEf46A
2l2Q4vczaCiyqOu7hOUn+TAEInnHr8bEGPCo7uZj0OmJfsWctscuU+436/1psjua
DD8FxQdOCzXykh78ci9hOiR+htDN6HTHwwn318g+6owycIHT632gWO8S3vPo/ksD
B1jwRAZH5OnFUoEZfWhdLNoplueNelQ5j+kYhSGlI0uIev0bEHogyO/+LdNK3SLG
QqTsbb6DX5k1QugmrT8GXe3MLvDjcebnNoBi/uAQf7BPyGRJcnOrqTA1PV9Id762
Isuh3FnkXk8KyHbN10he68VASdv0BxDzL8LZEIv4lsJNYw46/qWFuyD3VUZAWNyX
ANi3joZzJhRkbs916xebp+Ay/Mb0xBhR2jX5nvVTw++Dga2BfWHWSSzdgL1PObPC
w+/JGK5c9y/IPKWF6bwF8FGhE78uBuKKQe4enlfl0/5ZxZfxkXpPfUsPf6tasDDZ
hcktqujqlJKW9dQYfbITSBB2NnP2NrOH1SOjt0bQQdqGc3ZLIZcz98uCl4Fmymdx
+xCn9pFcnNm4MRGJ3G/mIiaY7BQ4DWuMmS+VP6n5l50j7RHXL8bVI5EgoXW+2p+A
KrvEaOFL9ELPJxkXTOYqZ5Z0f8Ny6VbzSistNe3W5EUDl43c8mn4xmEcME1tAh7k
TErXMuhAD/wPE869i34REY8msRrB65elbTPK/MP4UsCtGEYWNSHQVbx1JnDGfQvO
PfyuVWzOovELwIDYkCshYratW27NGHcvBb4aSQNBbuGMGuJAoErlIRVijve3NQis
WoRzLE4V94Dx4JenB7XJhr84nOKRDUqhutUugk4ogQ1T93+ZMiAmH+DSeOxcdl84
cGBukOyPP6p03TUXPpTPT/UMn57vnjPEpmimYVxn6S/bLtWm0BJ1klFQ3+OP6Xxb
6jYlVOGRBNPEv6bxN0BJ3KGNyICjBQUXRJbqMTVU8gUSa4oRzLmr6su2giUBYG48
gfgWZEA7VAteY9LXCJpJ5YbWLoWuFqUYzhOLSjjr4QdObmaz1evTOf1HVo0YQ/ST
ktGW1E5ud626FMF4nfFCHER1bSUEGY1hzYr5naaUATERMGTO4pXVWKn7eTIIPjT/
jJWCdKK9rd2THFqAhrVBKpRt/ZOBbpjmrSWZQLRuq4+jA2dxukrLhJ0yI49dyD8F
WQdzlGOB80rFFl7CrfGCdHPmc58LscFHax/56TcMksPCOGM7lp00yS1gc2jLir7/
cLv1CgbNdFr1O6OJganYnP0kMBwJGZAI84M3SOJ6dlNmUIwON41OcX1XCNEPbLyk
y+fmUHSzDIlRa/pbtZpHX6dWOJdp+DB+CvnDBQCNNAjGoOkwTlOg/soI6W3S261J
W2BQrxnKaljLROhGNX+ZElyIgRq0gYB/Go9PN/CN+vu7+S1ddW6EfvTFTBUHHvLq
LXqDzbgvcdsGGFW6KhTQxXeAxSwqasU/gjkUdYu7EtBhb9ls1y6cl+XXallAvEeK
qHD0nNsAF2hJpG8cwW8KpMQHc5BWoW0KVoPOjNpyeHJAS4ScU9xqxwKBPcCcYcCM
ax3NyAbtMSP+JRRFOfV4evGYeeKSHGWsKdRNPLpGnk7NtFEZm9+MQeOZstUGW/4w
HAtY9TPwE5R9i7OKWsmubWFNXGsukkZgQ5cT+nr2Ao9JieispHfd8rtUDeuCb+IL
Myrnn0eU5huj4JAdYR1BAHVoiydtZBnvTBo8azFC4otITdL4GTnVZeM2pXwAORma
1JQ+q/ySmqzz3GyYEST8Xy2GUkrk9fIHE44TgOTY8VYreAwRhgXrcuwzy7n4UrwF
FgDRHvWIv8yNM+ZXoWuo6rO7nv5dF5Xmu37NDV1TqOhKOrltISymJaXVTsHg1rsk
CsBl9JceaCcXyyDL8vtcupBuaExtNcAZAHxpdsDX8IhB+MpQK2Ex8LHWENm+u7J7
ZL24nev368e6+d3dThJIYse5QleBr4QHWVj48iH+dx9Eo4865KQH7WN95pSneiQT
n5QIdqNeL1PgRjo4dDZiNXMXCKessNBYOV7b0o2RApCdZJcZVm/U126vhinb/9/h
na5PW75khbqqbTTuck3mAOiNmi0BdcrL5TIpmduH9SyyzqzWz6ybjoUbn+N4kHee
WhJEOo9o1l6XpZzMWZkjIEdBPZGvw+uG0bqYHoAeZTVPj7waxGly4kqiJlLcTrdk
oQRTuS6JmxZxLtkr8956n0Y6thpvqNI1yVUnFUn4QQlH6G5RnBYe43/A4FRgBk6n
QFLQ4h+YSnwJGvZ2VDksEgqO8ZWg/MuWmCBpEUt7dhK02UfmIOWJ+5ahDltOrRA4
nA5G3kCLiCK7pnWqDIVhHxdWF52GadVZBc9nFVSCf4LEUNzYFtOyfXrR2GAKQHcP
kZyDfDQw4XnJwkYNOfcSDw1ZuUq8GsV4vyqRt33lT+0nR90Rd+vl9d1yKh+j3Stw
W5NIJ+1rIEbZ6KdeqeR36gvsTpf5LjMee6vqVE6bmZpfBcUvBgGOH66koHcJ2BVy
wuNI6q6Slu6UYCxVDmbFQzNMHeoSijEWVqoz2ZuN4SVzFimjdeLXjLz0X6LVbxQV
k8y0f9fhcQY+sL78ee/emsysiyhFpgr/496bI1Vo3p2ArWdG6l5ZbYI+TY1wBTa2
uoIaPC3TkhP6ElX9HbVovAVDyM3U8UXTSyI5T62hl7DbSpTUhypFg6eS74S0IJxE
25fvLpHXLov/3E7HT/O0zw/jjliwSlKs/02GC6hU8l8kOowjgrPTEpSXjnhdtLVH
9mo4cM+hU+mtsWM+rH7Ohm6/ha/dG2YMD/i4KdRC1B0wOJS8nzopUQjqPpEJx99v
mS2cUq+vAutWeytOg//nL6MaaD0CBfnd5GgGlA/fPrcUEn4tuOv4PHNCxLtqBoiQ
lo/D6ZNZaxjTDiUtZWfGPazcD5Z2hChi72CM8tUQToGic19fPFBhWvJQj3ptcuW4
ykx14lrfw7ahZjOfcm2j/kx5m5o7GM2N8TDb6gDhD7ud+arJdXfGEOp16rGXI4LD
s+WpBucnqPDu9Yx+xF6oM3gz03OgdQBwtsgXZXCsCvPiY5Lp0plT096SXAfBTYsD
IBJGsMVZo48H1SfBfY+nAtKaOgQ1a2/rpfQ4fwglufTU9UGm0c7YPaH6X3vCxgEm
bSgH117QcXJTI3YFetvHyONhdib9V11kcrdnumhPpAO/wBZS5Rvc2ST8oTsmkHR7
VwR4/P/X8AgbsHZRSzst0DOakV51JFVPXjkA9QAHY5CFAgwDB3IXaqtzYHavzjXz
sbMQebLRDgqfU7gw+ffKUDSSYQqsb+7xv7N5nBCfg9ofZ4U+1sK6oHPhygaVugUT
fblR3+5xTNe4B5tkoXhWdTsh3ar7rD5HfV131luNurGQlXkDx5yvHSqwgOpN2OgG
hNx0uwcpEmrOs7g/LHHj0fWqgKaHDkdfGzuL9h3l3UprCGak1SfkHZv6ov3kF1pX
hqZFxHXHKOIc7x4ie/UJ3N389cQoBfZKsELiq1SE2eeE7uWxrg+OaNfL2aO+2GJO
AG6z5Aclpnb85Zw1sxm/Z5E4Q0qHSdcGw0CF12bW4jIpEtROdYs07izWTbOfsXh7
+b6Ssho97OUXOLH4VMw+R+qhz6sZEjOIL1gtHQyXDaCy3/1H5FVL1iMfLsFiMy/O
ologzjvEWPD/28bn+1D0k5YSFCc51FykE3rHSRly8xXlnhTJ9D3V8MMEB7fIjyxM
uShhLWEhKpZRMvLqIvVTf7MIWDJAwuuggW4hYMiHQxcK1cTnDxX5o/8oq8MgQhPW
uAsDPKfty+njGXo26UF/OviCQhqct2q8Jf1mjgIKTrftOexzVZsaYIAlOE5OCNwS
IH2MGwyjyCknDx5hGN8+pvIvfb5regvnxkMkdKdoOQbh3V8QVqZo0uXn1zrGESok
mrxWXt3E6bU3LUn9FJ0ZXxCpUX6AImKdFLdLGSffO6FtTYVxXZAK0fUDT2CfEj9e
kSlv2LIpoDNHINoCATSI6umar+CjtkyKSXUBPS+8U5ZPcDHB3abgluXX6bDxIkCv
yjU/g56f1/GNVqFQi+2nVYQ1s+xK44AbOcD96+0HHyUgyacarsvFwOTND2jKaQq4
+IepDHBgyANwbSd0GPJj9vqpBZ5J+DUDwkjs4sC3GgAE+D5yvEp1yA5InMeMQU/3
6tGWmW26qGvW7+LRSHUN1OjLtH0zT/7MjmIps442d+sssiCp2wrnD2E7P0PJd37G
G2EPphU+kvTmuVNHOWd5vcoGHnaB0vbt9wFEKt5xS56RNVwiYrSA7UD95O14bi85
A7K+4zN/0sSlyXwPOnHIdTw32TbAiBxCUg0xREMlhwFna8kI9e4uAmXgt0D8LW5E
Ki+Ld7aUlrXAbSWyGBmPYDeKl7mLeTEyPCc8k/rkHTxSYTa7OGoesv9V6Qig/dR2
RnDIofQRW3vSs4W6rnwShnOwjVOg1U9cSXq1ACznMqK9TCKZUchbXr4ltCkd6xkI
SEEBVUoqjFzRQRzwpPvyjCHmeClFQyV09r36/Sd0N8eZNi42ZoyHh9jNxJ4IPT+3
QEiK25LIhG/9DJYEVNsIxrWb7jOHvmmarDVgfFCw9k3injgiBP061kGW/vX7B70a
aGy6IL13G0+R5IekMUg7gYfgOF9LGTjZ8V91eeMoEq6Ww9pUwS/7HoUMItz8rMf4
BQ15s0TRgK94SfP604fejoi8v5dyiuqjCIRiLgV33t+1p5qbXvhZtps/7aiJYndH
DXGNqbqEP6TeP/XeS7N7n3va15vC5XRzD7rRZqUZnuGUNR2BVkyjoU/OgsdgheqH
e6rAeOQJFqOiXy6m/D90nsTB6oH7t0JoD/49DrquB+59+T5B1gnXZjTxhlV/ddwU
IJ7K98AThv+7aYObUFPM0BEyJi+/oZ7ZbG76c3TJDq1nf/UCtGXYrkk2CaJxDDor
x+R8rQ7OfbnnG7taqpczLYGG43orpJD9HERPrPq5TwfHeAZkKJuBCu4fSf3hC+xn
LT7baUCNwopQQsct0C4fAy+JEiia840L2488BBIwzEgX3srjMWg7WqTNg/dElMbC
H+2Ct7iWnY61srPniRt7iloLy7ewkFQ9sphnqb2MZxUcQBWJJWtFeG0CUsSimq7D
WdEFxv/Px4JZN55l7yZ2LjlNRCbhiaS7WDKR0e888VSKg79CgApZBxurXhn9acQl
a8hSav2RhyXq1eu5FfClge+BUPxrWwe6xDjZ85y9F8mOQ6lGtgkHFqNzlcTJ1RLD
FgeWRr6N0Ks38WPRo6DzJ4r/KsO7LZQWPGELolzCLChLQJqgnb9r/r4vdYW+bgBg
QBhmLH8tSh+xtWB3JGRJKUnPpYx4L2kGw0oERsJPdmogAMYcqVlyfA4jUTW7p0qM
EmXuQI0IP3EDGd9L1t8SPgjkgTMsL6gskj480B7C6l9D3crxqvYFkXUBM9sxOT2E
4WBS9YBk7v3MQ5BG9S65auKJWQWGVywN9WMpHO74JXjF89GR/I+ubg1xVFzpMTPu
mDYlZeNUW5D5QHqLxMhDbh487P80e7TQ0y8AukeZLYkebHVelUJb7sge8LxvXfea
9uuac3quhVPXcznqqgmiedoYCu4UG4FuUURePjMDhZ8lXkRSw/JfgduaapI/ybO8
s//MvbzdIjChQc5rdiEwiw5z4HNS2H/YUcQvk8jgRp/eYkiFmHQe/17UkYI0+3ah
9LbOaQcDf3ZXP3Y6jH3jmC0p8cnFYoOOCv7glXHBYR8hBUMt8MSKrzh+YumpeQOZ
AuEJWYvKkraOj6CLabIY/7RZBTItigLBd1jejaGvfdIBol33w9/mZ+ZMNuJ8YuMp
6Qhtajel5oKvYOHTZI226i4vhmqmXpiP1bFFxi/Vn7xNoRkkVNI6zNppOAug+Uf/
IFjmrC4Wu5oQeRb1+EgbS7EtkKeQfXc3klBmG8AD2DSyvOz9Tawoq5gpLpeN+ur9
+cs+JQ7cjvnl320k971lIww/dLmS18BCUSjNBWdAKLSRUUusZydbwwhxas2e5m32
1GlKmR66rwhNqc30dxJ6FqWyziGoZC11MgZGs5U/b/AYh2Qn+YBTy4iT6jjTwUUt
989i4DonfeziibwIj514bud483JbXWt3QKR4kpmB0X2DP6E9GCKARGnGMpoEjLCW
O0H6oHpElTcl+AGpO0Vxd6bLR5cFVSj5SrjRBS8JRFUw+H+OCRxQAC7KkZ+JKQ8G
34Jiep0P9lYJGYH6ODEn5mmaO1+KeDfCv+1bGs4rRfU/At0MqnJkwy/by/BvYb/L
/J9SqNxjlcHGyERdSz/94KWAZ6C6SnWc+pvdd/s+DDW34W/jRa0jRbDPo5076nzb
Bw0FaViXGIOB0nC85hQvSrEkRE5hfQjFCF+TJ/yuZgOmnmMSB1DD9nRfXEUEHNc9
R6Gcd9Sn3Nox2ljcyEvgzy3Ck5MYVpUmwiwLdCFfRuR1SSKeaDmbWWtqbuYoDVFd
Q/0BYwBXEk28cC6rFBGv1WiHS5SGSfnhWYiroXX5Yp/XkLBMbiATOnKKWCwFy2Ks
Dw6C/G86ZVWd813Hha2Mi7Gf3x7t7V8cm3FHhegMLkjisTrSiC/ktN37hvV89etW
DbLrvSVHwbFOUA/7QVnsVcTYAZq/xP0fVJaCbeZO/dqObu0ApIuULjLiqmowdHyk
+6ewUxkTJtoj6Vbj7UBo+09YBZ014hVeBmy1ndEAdLXhc/835z9tRb4HfZO4lokM
j0Qppb+RwsTriBzG7a3o+Nd45GNTDGebso60nqRKp8MBeCH72vPqDTkMeHHTdJfF
iRWFkxTAmth0MkyE67T3g4wrLlt906/iQIbev1HPM228VWlV+Zxf462QXHaVG455
iaewCqsZQLFcXUv5kx2RUgG2kAjKfLn0Kt6N8L76GXQvyGgNEakNSoE0+WrCEtZu
s2RmwaOj6ZxQ48zb+1QPkdWV6bEctqk453WxhMklqXjgFwAZs5eXHIitwn3Nr1up
AX8tQsvF9boyU2r46BrRsgiEzq8ze57TIi/vJBOCPozJ3T1vpgng6EBQFBSm2GAZ
+AaUtJjaNZd4qAFTJmGU8/3T/Eyh7PRvBbzwKiwDhvelVodA8UuLC0iBRKtrfeJ4
EpVTrbKzs2d315pmjuTTae9+giMVZAmyS6BE2p6UFprqp0OeqCJhdl159Tt4alBw
1NF0JHBLh4icw1q3putWvq27dAk5cXVVxX+UGKXsSNoGXfYGIbseg5qZ+gjzggDd
7jIAAzJyLmSk/J+17XlqV50JdeSgUFpU6q2voYKdEIsaZqW/c9ZdRaToKlMygcut
THVq9SzVmxm3kR9ExYxJxsTGAhCZ6IhTx9sx58k5Yo0flGdGAYQhkhLAL4a/dnZk
Kmif+H1P6GuJ/TRizji7thgzbLxONHjdQm3cGrNUOCHCd4PQyPmIoZesRuIiLEtb
G56Na+YqOpCyoCg8HVbJS938YQhabAHlC77U/0OKc6pXOpE91HbPJEAiePKkTvyJ
dlTF12GM8jZawZ0YDe1JFepsh8DnzwZgScT8gx+QejX4wv0ZnvbZNFp6E2FlmwXS
tABdakhf4E+ssI/AcImrct61//BgmBLPE8mnOWWhRN2DiDWxueSFakhLds2PWZkb
xX994LlrYqYUh57r9H0oHgnXK0QW/Ae9OdSUwOfZWTdU3vI+8C75m6cdIv1t7WVX
qNoPXYaU/oehzJOPYUyJySilcymqhBl8TPguhd42r449CsXSj93uJO8ddq9V6B1U
Cb4GRdeZYVDTgmwmycB/UJ8UCiNP9RHpw71+d49ryUZazruMAAHd/E2a7N+fnVwc
BlqHvyWKOBNfL0Oksv4SpZx1NscCG7jYQ8GTQgMuPJRZVloip67Dgn6cE8kq5xRF
IcKivYTWL5drhT8ruSE87hCxDJrqjusm82hLLUr/hkWuJ1H0M6TFNiVTiS8/zfNt
e9g8gacoOqLbSu5hBBQKN7Mu/FYAoNW33ytSOQw5fWBovsqRnvv3GbAXEgXecz/L
j/S7motCmCC8uWvMVaxBi9St2WU0dD9d3bIHW32emoqY+GdehpdybC2hbLtQPZy8
X6sTdJEcN3e4NiO4PeQvq1DaHob85viFAuO4NjoZib/PoCRYzOsr0LeLeH+iV9Tf
992duW/fpLt2vtHKCAYbLfgepoI/a7NCGZ2lHW02Xwn/pEgTarpoDGoT46VTfufY
Y7MWtRXJBFCieOadZIm1CUdNRSwrNM/EcqPbNj41KeGsUsBGQd++ji8gVHMRU9Jq
JX1F2K1HjEOFRj5X18FybYmYCvHSlQPGTXSxQLCXoR68Z3tiJORRCTnVBK+wb/52
n0SpG4prrrFveIT5Kr20cMSw4RE4+dRHO3KWkNSb3BzxTxRDQ7EHcTNY53iDr3Ge
x/vzUsu1V9nP8WjWiIq0+e6PE1eSFycfQbwkkTrHi4puwKv/CtxammUFbBfxfDmU
Qa8R6QYmfx12c3lGiTqkmUHCP4G0rZ+QJ5CRzIifLJ/RH7fGez/Ku7xu8GEEM5MI
Q2hd2UNO4CEt1oMCRJZ70ymD4ciUqGTx76J6XN6xkFPhKuCsYUYFHaEiZ2u2KXAW
ZZQ6HFq3nOaHg7DLrZTomaTRqMcH2u5H2jAyyryXIQ+KcaqGhMA/u8vT3s8PM6Qb
14OGpyt5lEtDWhca0F6QfKjNkzzxSfvDBskAZ49RNXMM3TgWEvrnm27gxeWqcPlE
khN4Tsgv4ArxHiTD1InuWv/+CxaUYfjY42wc8KogykYeigpoZn2nwsGQyX9JSQaJ
rvnkxXVPfdFN0r80iDUAqYriDFu4UmtwBZac3BDR0MHp0LzSyte1Q+Z0e3y8ODNF
N7K4Cvk70aJ6oJUk2kmorTPIAmokAjEHJsLrl+FEHsbgI1oeWeQOvtYM/yGr83Wm
P0sOFndFhbJM2xCrJk9QBDEw/+j2u5MGY4odYIhawvAp9t+KukLpUS6e+8gHcb/E
cH5YwiicQ8NxNmYn+PAekPC+Bv/PsyaCz/2TUeVtzOQEyScXMYhZUw88rh87ntfD
oejKn4wMM5CSjJg2PfUmSio0GOvPsjJ40iOHBWj/U0WqQ3XEoutbQxSL4uCqKHz7
pXdHi5zIz7/iioHErgjFtRgmJPFp6KciXGKBSwEhlo8h40wmo4dsEimbSNxJtF62
ozTn/vwArUpqY3k119bwXPd0ki2X2q2anDfVBmrd0eSZBHPlD3n6H4p54hyLLpOX
6IFME2tl9sZ2hHDfaQ7hA3CTrJSMPjnFF/GjvYAaDO3wpmjGNLEuqEPJz8zBNZm5
d4Y9SqLP+36cAgE8uEdesIDN9ZzYC91d3zLnnL7FwM2/wIPauNNwOMOd5/aqJh1u
Hnt8S7yZ1/84uICAsPKQ3e0kglF0ogv1t32iAEgRIeNbQdPV3OgzwNHQMvZmF316
G5c0g5M+ykhbDXZVuq0wB4tZt0wf+Nlc+Q9OjGS87uMI4v1wjGt09sfnGcSpkIlP
ITmGwdWGrTnSxUgrGNRjxpaBavIpgokGzkyoqfNwl6yXjzfax1b0xfN5VmfIN/Yq
qV9rNQXERyGREKDp/3z/1OOgjowXbs0eNF77L4hHAtUU7RZIsqzimyAaOrqH7g0X
HebSjZ6tivnY/Zv5ypaXsbpWydsT5LPhiDsi51pGoleyszHJiDmpoDPH9m6odEYH
JE8FSxF9WV5yrrOUNLq6RyjuxHh2sOvJPPM6J8cDD2TDiZPmB9WFMqQW88k+bw3P
5PMhSCfTgYTg+NPZimkqHTopHK6DHjRjimWvr1+taKxqex2PcXqA+vjuHDNgREYh
XGfu0p3jAJYSK58/iZzbytYOZpddHjGqpe/B9kKk9YdO02/x50Vgwc28tsSgUBDD
eBtcql8FNiHHHawXkJnAcveGj3WnD19jXZCENLZSyP0qwIHsUHuXUF1hnIa9TXbb
fVTfZwoy5lrODmf/1AUtH3jh+a9xTAV3vBwoKczxT19iCWq9mmiO+n6ED1DLhtBD
vF47tTiEpJFQmOg048whONTmlnIVJ+ZdGMqanQzm8Sj6pX4ELwqonNlTpq+HnKJ/
aC8YwmAOpNTLXqzgzx4HNH80Qhv5MscxdZOH561xmuh+2nY94+WaPg3TsKt0OH0U
OUcp77FitSN1/W7CLfk156Efva2o1JXTl+rl4iFMwsLCV2sxn2p6KVW4HcsXgTS7
ddP9gJZHKRqWidCkcXsAKKTU22FV4J/4C85rPSf+JjiWi8IZ5ns/gC9495RSqpQe
0OvUeSjCQfJVeXqKbsf1Nehmy8tvzUS9LN5Vf90S04PcXdvuz7RtKQmlB44TAqSb
NWMgoFdUAvxV7ekTAKRRfqgV+TlJoiP8SOUTuFIb5q4XIZA594P2CQ+Y9Wz+M57h
OeepfY7zuO65QA+Yl/jrjn1wudzQevuF6PdsKqgn9mvd2xc9/a9/X2Nn5Nl/W3h0
DES/KDzCtHK8SgRaH85xLnqb64/KeJzGbfe7UTF4Q91Om2MDQOdT5snB6FvMuGds
j012YNl0EMK8A1gsqoVWZq69BTbSQR5YDhvkwWke37T6dQ1z+aQz40u6WZQx3I1o
k9Bro5JFolcRiqR9YRdaDlRkT9xCMYOueJRkRn3iQvCaaWV5ScEX22uquJmmXv1U
abc+tR2w33bt3gZrN+uZOmyFJyZRDfRW2rfFomqIo9Shw+yhJHiP25O+JOUm7hUv
X6SnnXA4UPPrqPE3lbJgRA8cfDsHyVFPOlUE7xoknaH4OBl9bGvsiQHLuAlpfbxr
jbI8RT85ttKyaLfANJkc1YTz9igtz6YREA2qdwlbfk3GfheTgZspw5fc3zYxb2ri
5U/Nv1oY/IrmI4i7+cwqg8o+uIOt8SluQtosAi7Yhm2xeeYCmTsMCfSJmc465LuX
r3Q5+BtjAGBGflVjmPGO1YW1NsC9Yy23X6BvBFMbqtxQ6PL8EYDBbL+z5g49mMYi
VQL0DIbmQZX0+EjdfcSxwxVyH3qSQM2oW59Q27Yhm8kkBD1os+TliY7iTsaYjhkv
ucyObALoExt8zixjWwuo4hookx1LelZKx7xTuf0K3/zOkxgUbRWGCw3XXznEcwjJ
U1zUmxfq49WObA3L76fB73oaTtCZd+lnPRtmIZbro7YW3BVqfT3j1ES/2dj/JXw6
iSuXkhrVNUWOtwA9gkuxw3DQeWey85rDG2xYyvkYSY77ccBp+QH04b125957+TfY
cSc3ZtnNQo9XU2ncKw3WabDfZT5p+Whm8sFWxi8MsYCgee+iyOakbaPOR1X6NOAc
UPL8E6ukp9apa2Ynf22DdnGC+0mw/BH2fC8936rUlhM+5ChTY2Gc4K8TI6BtkZlt
+RiIq10hBjKbCT55VpgX7X+cxq86EMFhbz5hf8SStjpL2S67LO8w7xezfd2/oKma
/A0wTO5LmdMumr7nCVBkYrGzlB4j8ZIYkZ4jTRchmXnipJNW5IN0eyOviNq3TYTo
gEvBeTBlU7HAaYF36BxtkSQiDLrhoMN0HDh6qnBvqNT5QeWcQOd80466sG22jodA
vyDkdp3ZEkR1q8AEUq2dsKfDRpFlFJVkDRQlylBUEoiihejuaUWyN+ghYBuK6d25
38FRVcmPwSq2XrnywdRlj+mtiBMmrvqyjDH7FyZtXerAet5Vd7pyoIh6YKVWQpWp
7xqNECr91Bm/lLdXzh8XYk0wD+f9RAHanjgXWdIiGY9vAoeYgpCIkdn/ruB9i1yH
8wlEl/DVL4deFT/xQUnxdt+H4SGt8VQAjZKfWuP2SauTvEu3cwjElnAIFg9V5pk0
kliZKvWehJoo6fIB6L5f6Dhyhp7wHpK3Jfw0TqogC6kVGG+a4BfDvyfWknW6fOs/
1zaGwP6J0DK7yLf02ZrB/598r5MvJ7vWzRqvoB0KrICs1E371u+2jiuIxV70Iv/Z
5oZ3aXb59xSnCfkgrMAk+incBl58guBp22mzcB4jf+jgNLbxF65KmQv7O74z0r3x
oSZNxZTTYTaTrpQ71Np7mKiH4Lsyyj+HVJVS3Cb2TdysWqMxqZAg2K+SE/6OQkbM
8e5cgAOVyO3l429G23VfR17+tPcy9aLULBq/JRy7izLGQJDbi/Kut8LalQFtspYN
Az00n4pX6Twcjt0BiJ5fmc+3tufASsTILQOJ0xExXZqxOG6ljBa7sJn1cOiw6Kul
iv7UpQPgvDUaNy94e8VdlGkbkh9mBkMMLwFD97LkQQG5GzCA3PJgL2E5D4gYWxCZ
qIe8uV23KWhwhm04XCfpjgqWjudbJ9o+TJVwg0qovsfQoPc0Ip2AwlMKjHfSyGCn
yt1RRjwc13ThvIZ1PYmI9lE+TbXzFHqhm03Y/XmqWpUuuUnwYEkgDR3Sk9zomjz5
saIlr/cvAK7tYKx2S/yrvB0N2TbhWG5TEhcocyPrHeqPSFMOP4mySQ1XK+aimXUt
fqmgdFcOpAxzAKeHFlpsl6btNfwFlT6jsUtshDd43yCwFhHfKzbG2PCbeq4UaRld
HxnMgj/+phyt0Xaq6M7PJBpQ4DIg1/bRsMFtg0dJkoncC9XWymVmofFSLi2gPDOB
8OiemqbRVokeiI9Ny0oQ+c4HcyREm5JOSGWgeNdRyvoIDpQ0Dn5FlprJ946zc1Lh
Ju7VXEZYQYEY+fsmvhDMP1yG3R0xkSTPjl3bFlwB6Ol3m5mztw67Rdu6wT2CuLjl
Xtxi0pHsgy5NI5hkvxCczmMxOzadMSCrngp0ozUQ3IioGIhhqn6XyN05nWbH6Clm
l9qqBErDYAKUW1ylJazUXrak8Mia/RSIB+zSuzKxVohQYLcjcuz21nD9RmoF8DFg
UaIuQB34pEZVF1a9qulsB6YvoJPovwzBKAnwrqhfVjGB00r1u7kUZAMwZ6gJIFkh
8kC19syP7cIL/iz8fMLKY75innJh8zYSgV+RxOekdJmz2OwlCsP32osbPnd/62RU
OoRqxCTX08CdEBGrnDUeA7DaonTZzgTm9v96Or3DMLxz8xwtiAFb4K7t4tzz5qgT
nFN9xB0psvSI3Mfgjo5NV1nJbbtgMxusyIDZ4VmpZt7BLKT8+9lo2RQDY09TkHMe
RvZkGNkhvncaLxEyZHDqevBcbe70xDOFimQHAaJOQg6kX6Ze5RjggP5Zg246AfpJ
bZnK7bI2MN5tqG6TirlLJ9bmRZCLUg6XmDdI3EHmRcaTuBgEc/3OW3LrQfdRcZjD
PijIrKcNfiA4xpRHcvnUA1Y3YbFKvR+3Mc1p8Hm7m75Ot0crGSYJ74KeTG4YLLG+
lyZXbC8qHllJh4foZqJCdyL93YYr9FjX7d+CWekTA2pXcDNRTxKekhVtwTFzRMDW
N70I5Hv4eW4m/dItjygzV2cCpSlVNN3yf6I80YXEKazGqkwVg1UFD3/QCoJSTwqW
G20q2WqLzQESjlSlvFf+tYKF9bFjyW0aaN8CCjXIka3oEdauUvz77Y+XjFSY2jlu
RiCmBvI0iSkrLHvqhN8btQAM+Mrm23FXtbhq/gWJUT2yi5b5hyQ2lcr663CjJgGR
lgDlnvIwDygn3YVvY29UH5i66V/yo+JoPyVIprDqryXuKdYydyz2WM6qYl34jpWL
B7aWA6tUrHjryzdN2WP9yzw0Dx2FzVTnBSNl58Wk9Za8NLgZRRPVNIS2dQHrjnIC
cknF62Mtukz3J1tDHTkzlv96s9qzAc5hwnILuvNTf2LFZjY7oKolHzv111xxIwA7
nrMqR8uaL1Fx7CTjova8IupgumId2Fb1AGwyvOy9P8TRd1/uxSkSdvL1IgKRJPHe
bSn2o8WcG+h5MpS04AzdImnNtNAoD6ctkkTeRttcedZR2nn346zZx8FlCOzAaPxL
TsUFL7cLlu0R94Lf+zFnCFgAyfRusjkndcLLwvJOs8ukusqhzxg/VSgNxSl9Q7oP
O8C0TrBYDPaVTqoBk4YoDOHeURB8NG0UQqfYXU8Qwg6d4bCusRNHAwS/NdxdB9jO
dpTdrZfqVnENYgTwfI0K6iIcm6UsWE+DrOyVntu2TyK852I/wXGgaK9s6wLOr3WP
S6kK/jJXXYq5FzoAXvdtuyq/XSaMRuxwvCiTBsJ6I4cOc4f7vdrOpt5IovoJar/r
21hmWBNZpp9rkJIiqYNypJwyedgFKwwEP0NtB8agFUo8eYDY5zlyRwA3l/XIJF4a
q3/b3Jz4TvTRJjTI+T2dAwE6JDieuvfjy8ynj5K+QDW/poIbEYgWHI0p13eW3MJ/
AmWWu5FKXBgrc0t2mSdIQIiMlmms9BfpPmYyk2R34xT6iRdrv9hLyefsmEwoqhf5
O9Z0ERFyRlIx8Zr75SuVsomQo2F2QjSvUnAVsprs5hnbte/D3AUJ9f7Uzbb4GaZP
IENrRo9jMI7EqCdnk0gDf577JYwKXFtmV/hL2cs7Lwf3j6rjTXukf0KPMddfaTIp
ZNClATisbd827bQHeNEFqRnErlQiHwShj7CR4u2zcTwxoIJQZIZNOwhLtkC4wyso
eDje7ZZBblhrprixJYd+4EuMy7u+TcYU3FREDNgNRvUFHDf5VS1j7l17mFZa8z0s
FDUml/e6AIGdE+Gai+Gh3EQGw9Lg2sxXuVTQ3hC0mQ9hRNh67wBzv2rRuIGzc5TX
1ZGZBONw1iFXAyZqCbF6DRVLWuiIQqYq3RLdQdZ6Sqmfo/Nns/7w7R2fbUSVZXqc
SOjyShY8d3JTOLoTg0fIsBoZXrsXMReebEwpUAyOw/N6lEQlybuWxAwRKh0LUVkd
Livi5whdAMWombbdiNkTsM0Unjiogz29AD6U+Ms8So7FT5V2WFDlda23t0DPmKnd
tW174OgHQmEUwRRGYr0e8Nux2G+t7Ns53OEIcLIJivIJ2wWXeBC7nGcB/OtpgtRW
dhw8d8hIQf06GSTMOQV4GMwXSESaPWyaZScP6ixzANYuWPjICYTpderl53kt6ouS
l6RYi9EtdZ2vuf5sN5kOBEUpvkjfywR5dbTQhMr8KLCv/txzWBSWdnNQgb4I88pM
CPpJUIoK7a4bUcNp8PblQ5/6bUMGei24kYDZCTiKP4NmS7XAGzIIIAzgd7mRa0ub
jM6XJH3FWoRfmgbvC6xU3k8CElIIpHupv88GFdDjf82TFHO1LAOYdBvQJT5sAbHh
ujmm9o+NQkvFx9E9Pnwgp74N4Fzc6QAO9aA9EoMy1IE+sXhYXEXLJ2kftdDk7a//
FFoqfUWY+iaLm5TFdOUcxt0wk6/YWMF7/PzNmsqtiUgbXkC9u3VNQProwHkBALck
Mh37EQLu7NuyXOqG5WXGtJ1omWD+1qPgWeGXGi58GFgWYNwIm3dnE7igdC61TzZn
rKZw25xEn7UMLDUdlCBTeCnNUN2+RW3ZMKSUREQfxws0YILcd1WPhIxJogRoHmPl
JosgEOmvcfxluempd2+hdj6FXhgeJ0N5es87L9XXsw48Vp//HcYBesmasFh+gzBx
TkbZOTPLjssp+U0xnvC9NHzAuF4ys1DY+DeHrany+Q4kS5DwQeDVvA1Mqw3CEcNs
XIjb0pw03PQYNfh/2uXHlCWXpQMpQQWEejv8uEdzhcF9LwPXlyU135EKEniyFov2
HCI6CbKsSxnmXthPJyUK1DXg0Te5RSLwhkL+v330cmetfZfw68uNWcguVSYb0HLU
XhwwEmsf41BbBR7JSLH9/b4+P5lFPhf2B53XQTD+TMlOVjQhO9L8e8E7iHx+ZqRO
RnwYTcNGxFuBhNJr5oNiZuXKY5DUCoaUbDvoj/CHcqV8joAyQLpvgF2Nk9qJd2Pj
ZBOAndL31cT96zYDbz5Hp0J2Kq6l0Knx85fBak7j2SAz0UvKNtBX+fBZrPtBayu5
Zp5a2n7tu7DW/UTRntjdwlqcOoRk+JdVJBUQWiLv31CVWbo/RNg5OrEy07oAd87z
UL9GvGZ3IPwLO1VVDL75aeB/lHnAKRvRBqNtWoFQdNbNkCWlgw9Xm5US2TUW7xED
zsOEmb8PADiujeutwpcMRC/4p8EnDF62CWW8nHc+nBcIf7kDCr8TgZhSYmPkUeju
NRW7w/5du7HJjkMp63F2KTq51Ml3N7ntKIZjVl6kBD84hwhNYgoj/tW/VfWcCo4M
AWxJH6zu+ECFp7GRHZDgliVFRC9C5gub+v/H8nH4vytq6Nih4zBOcEPuHCkFXM3z
ppPj0oC9GxJSm2Pv8aAIzWhADX8CR0Ts4B7aU9Zpd6WS3sSochzUrFd/nOB6UUkz
wChhUHkPofu+jyKwQu8184Kawbl5XMVpdbiCqdLGgtPkp7h+WZxfYTkQMsXxrlIH
jlnZAng2lQJJNYoqRdi0CwrxL78FH0Im+gwCYiY474OI5X/3DKm+nK71SwmCShD5
dEnlN/X3juUeOJt92oxRf39qPRwTLbE2f7NGPsudiU9TzvIAkrC0xdosQMqnOWRM
W/Kz6EvoGoUoKFJb6Qm+TaDAFkM+Pbc4MGMYe2nYzKeEDNi1CKsYzlPdSnSfoL12
DwznGGClf5IS7mqWZvihHqn3ybXP+wmQ2/Qlaga8RdKKIYSoSx8RD5O2ijx3DfQa
wnNFWYedOwbm62X4VGNfOAfXcth6D414zZgAq9oq6abETfK1QRcYsSdRkEfKrimv
vwafvfdAxjfsll9pD+sV3xki3IJXkgpgppmAaPz5+tPaxdUqxPRSm6A82ln0xEqX
iWA2VwENYSpuEaEhwu2GyjD87atFg48CvMCd31PElZLnNGmrwoPvbttSWX0CZxMo
MWlymPiEAAmTvOFPG4YZCKtN+1bvx9AGHOFxAWC7v6TATkMUz7ikEOQAIN0NpGhp
DfvkJXppG7VnjckFniZ+xN3jBjKngxxstbY2RWfjQORJLy7gHvGLMCO3Y4aNPkd0
GC0G2cGzq/1QZ9ELrOaBYqu/evqHW7c3qkNLCR16VAaePlYpL1toIijb9oXL/JHE
OtdXyRq0sYV4uc2wM71dRaOH/t5F9Y00/IvngN4VWxzRjJP0Ez4ZrJCcGibGMnhr
iGQagBOTBs3YapVWJ00+h/scxGKxHHrYTb70nLXbNb2XQp1cHZ0VtsbZoknKDDr4
UPcy0D4z03m5MILWcg46OFe1qGmJFzKip4iyTwwaXz6dRLe4q2/97s8JY+iDoYcm
UNOFCSc+y/z3F+OBsVdGbjmQPKlFIhdx54oNHhVoT4ZdG8tIVcf3jGU1dCGlfuxI
WTG2cCTrco8KV/XgEu03kIzGFb7GJ7Cqxbix8aAYsO9ycP5/a8Vf0SdbIf8Y0wlA
Q/m6N/aDre3CEjPs6vlYVpHShF/H9hskdtUmsDzKgJbWROdOjoT5UWIsEv2jXewI
XN3U8ngFQc0TT3WOq7U0iGe1NS+G6lwetn6DBvMxgA14CGlsH7BrWgfiLKmv/YL7
ayrtlT0WMLhm8ATxm+PHsOOboZ910zMAz3KZbpPXweYcUzgF1NsuIw3oeKodb4nm
KheahGE4+pqm4wR8pasHXz4x3LVZHb8RptXHZIg+HqUFmSKqXWm9g+t5kw7Sqsv5
X1tXabfUMB+U7cpYs1jt8Yca0HCsZXvlcvfEo5M2Plm/KJRBG52FBOFCd5sJ2sr7
hMolCFN+GLDPrnA4IRs0LFcxPnD38LUp+zr0FUCd/NbY4KE4SkuXFEJQ3OBFOvmP
rchR5glQx55cduA7BZWzJwizOndwdIj8iLNhtavgeZqS+zgJEwhquj4jz87y2NUV
lxA3Ed3YZ8agSFCEXeLCf+KbGPIXxwJ7sP2VzdNC9Gppjjr3yD/1xPngstEycKWO
LuFhfmlFK7Ib1hICHuDdoGmd+G4JWGEljtv19MhavOWVA+LxDevwmjTkoUpPJqGl
cy5u3tac+J6YaE+Gm4hWMROvjf5cb+bE5bvS7eV4QZqPsjG7LQcisZjwVFIhHX2W
f8n2ksL0FAZSRM3x1NKy7pvbaELLJTAUlKdWtdMOk5Imag+CXAciegF6meINoXhK
ZZPQLownZ2LVIEbfcCVIUgHcFEEPlhtjqyfnY9q86wB9CZGW3raKMPnMJry5LOwi
ILxuYcKpK4e5I5FE3W3FbCKaRIPc9Azapu3aQJ7Czp14TXbcLkdk+MCmBpFNN5Ao
/GzP9MhW6u8rSkqvsmgms9iyBYYpgvwnF1GxEBHVspUaSDte7dcnDfor2GKvcaS5
NeckrRTYs25F1AD5PHHMS/tLcYHgorWy84lI2l5swq5PCDTpnaRJsgwORdCIJ1wa
QySN+F35mMYUesUrQ/6pO7GYHAo7gCk5S6erueTsdkYsm/MNV0pU+X8no8kLV4ul
ewhazWB9clhc8kHTbDGZRMZwRQqojQU+OzgKmQsUguMcGMiq31T9FCMCf3h0tVfO
8iqbMbhbSLtGZ5++2YYITC3bztH1Q2ms3GoctHhxxHxzmu+NaAFPePvDXjIXy4mm
7ZLjf9uSSo05p3vywli6BWSvfFucMD5XHmHmgIjBKLcJEQ3eWLgzQLCDENVAptDo
c9Ov4hq4FAMIhpC31vpCbYiWjQ9mMClM3j8o+l0VZd70bnt8xNd99fP/HSrx4nGi
hQ7fsgdkXZ0zF2yKKc2KeoJ387DYdNnPvvk+N21ZWWzk396bZpr/diJYQTD2+kF9
Vy4G9wC9FFR9PzJ3RPt/r7OITK8aKgXgdQlahcZHRBIddfVKQ7tgVCcOWzu0neYr
MlOkgg9O23raKSXPa7ZEQNYvU8+pHGA6FA7eEWvVkENZuT2j/krSKUyyQelWYMI3
2CB+gqFvc0Gq0CdRQGTEqK/A6tJK9vU1nA96c81x9hNG/CVRiVfIGuohBYuHsCL/
UErmgZpjugMNwLNndeiErRIT8MQzGuw/4M33xXnG2MQZliP4H+P7V51wy9nWxCJ1
sguo6mkGYFVce5MWBGyLqVlQVqxvgkwWvMyKMTGebTwnVCcWnRt2T0mIZ7MoMSDb
LYOt9qWo6gwuzsAsUwczV8GtRq6vqN+h71jsUAKGnbL7gwcfEOURU8r04M4hzqx1
lfkJLaiExCpb2ZpxnwUqjHGx7rrewL92CFcdnv+1UiybK1aPvDHb9FZyG6y4HKva
C2kfI25BBxStavSZDW+zFYGPIFYU8nt6/wolcEzdGicykCnI32+dyHw47TEhOeBt
SKScIr9lHMmD8eW3bQ+2CN0DjpAFvmDehALI3QWQe/OTq4YxDPRW+BiDlaVscQZA
UMRZgNJHdWsi5jYdXM7+bNRIct3pgPmCNHa44uGod1ayGNoqXVjRATxbRT3kitBX
t79UXT1ESAmLDEQTpJPzChzuye5usdSrLKI5XDdbG0JuaXuXvkkLlvdnM7T+TXKz
RcnbKZQFZrA90nnRpOsYPwzENcAiEe8Xd0g2lPDuK2sBPgH8MTWI5F0LKesivhuz
nCBbd2jNmiK0kDDhiVeH8JUhMYFGK93QC0eWat+lw6SkyAXqKOhQISm49tFiujIw
4Oxyeur3hM0f16q4VJ+rwkq02AIb9CMJMPx32Ry5ZrkGol52sDEeGn00vYU6Ndju
79wck9QL1Z4xR1s9XmgNB88XeBQu+2pNhbqHMjPRfpyb3YtAiwrGohWVFV3iTeP1
od6nMzffcIXbX18pd2MrXxTG535SmqKtZjMX/D/TiUUOGbNBrJhvSXZlDoF8BQkV
Blij/H4DyRIkald+FOxpA0iwoBzMfF4y8ysU6nsKLZt5fuxF7TqhbhGsXRm/P9su
p+536nBh9ecb5CSXhgp9ecKMNsbNwW9jcWTtVhxt94Gn7X+dekLZJvORYu1T/6g/
ZXkUCSS2i/38j8VDfREC/fuiwn429SO/QnPH0MYQC4MJtZ6PyRfkp3jYMzMOSWsQ
l65neQFJ2H+xSKBbu+tJVoPLX99gJR5/QcZVKijDvbtcYzYmJ4IWZii4nIsMiXIv
kZqxCxNgQ/NPmiHCizYDILvrPadtqZbgWHtBkgSx6xfTQF87W5IIHZDDYsMnJp/F
eVqlhJi8493fhwy6uyM31XspE+v2dNp4qFI2fAPwm6BWJvvM9Wx3BIl0gFFjx/+v
sEC3IBMI61VmDaC0YrAfpv47MEtIKhg8cltKslRquGIjW7q/ZIeQJjL5638H+7O2
qW8RKzcKrFy3RFz7P8+JOaSSaSxfrTmP8VtcGx+S+jyV4XiK+URcCdesZvVudR9i
aP2ZoeiplNZNhfjJOWt0Tn+xHBf2x5QdxeRRHSCTeydDjVTq1AxZEBNcOH0YxkmX
A7fOmfr92PaJdwREOAAuhGd6Zomji/83CoS5oKoVO6W9isgIeMBOC01w5bdgZZZK
CwXZEmeTASOqXKsXnT7mcKxlP55vqagkWPVslBWAbondBdmZsvNXoYeQBJ7hNy1W
Q5G7KmuJUXfFliDEEEke6ec1Y13sUHEDxepF+bEBmRqL8HWShukNDBtcgRqfzNIG
UMXd5bpjiMrVGoQEyzscYhJxNtM+ZLysoQ9yvdrRBB3oZIjujSUN3E28CIYce+3R
98+LVWX/m5hu3mJhaCSi1XBSyRsvWZexaKqcdhurGVYt1hI55HtJLmf6hyYXGnQb
aRAZsT51U4bi5wCAE7tNaSkVPT4vKaaCCf1RDqKV/CAZLN2sgGnjB8mmpt0lN4Oe
UV/OrJbpIcGTfYmDEhTKgVRi/kbPheUl1ta8Buu1cnVs3XWdh+68rqKUFVW+kGp6
p64IlCo7iNHg4KzjKlF7kat6KtHSoDAA5l0nPui5KcWQ21ml6kMbqlLk1yrJjYgx
OPI4riqc2sewDm8IsqKd87p6T9B3UsrBw+Fueub0g4UZJNxfIfvKkK4V+kvY0Xdn
u+yUtRDOyxWebS4C22iibysr4Xob2CBOuRiZJch4wcd+kdlZX+J307XdaXVDbe83
Z7mfAb97/yGR3HiOVhbvHLutitnAtt7Fc/HZZoLXkuNYm8KKOLsJTs7m+6+Iodu7
xrKoD50tgT0P3rLaf6JLERv6xEDn9pK9B1QZoAISTe7kDc0NlewkbKX+MJwUQUU+
hirbuswIZJLGsJxfVWj6EtnomCL/XjLfhD6Yu5Qfb5/LqRxV8hH9XaxHx/RZNBbH
jpBwHkENdOrN56PH+8XXOauL0feaQcEpSPK6YmglfTO1b/XTSAja+qBk+C4D2fGf
Q91HpHelBXkgS5qI26CwHAFkIAnHp8gvYJ0mlnu8TMPZyg9eqCuLvZQ3jYhgH/BG
2XOyDibuktzYC4J6nQHJTOhgmJ+jk+2yaLj3/3wPIjmnr1mBYGo2W+6bor17xgSP
vqDiUhkyIxL2vJaW8U5GPZSdJvG3aL2/2xOGbDfm2N7JwdE8kqaPzxJpoWBaXd+P
6qh+hiaZQA20Ff0b8VRck2Eo13VUiE+m8ofhuuLQjLuKvXru3YaGE4d49jgZxgSc
WtEZduOg0sQAUt27qSILLppaiu/CFaPaYMKB7whcpnIHMIgyCTfdNWQkF827p6Ul
NNmj9McErjdsFYH0+LvV4uFIpVMYXkQw6tbRUE5pFvKoQ3JwEg45irs/U3nICoSV
cNZzADnbmpijSCB8IJF8xeVwfKymvAhXNJSCPyFGHKZwdC1DXKg+1wjunNQXAeG5
PlQEPdXHWLwQu4J2UMk+L/r+wCNGcaVGhLvwYnXv/r6vyFh+dM9zsvo4ezCyCK9g
MjydzqSunTlatZvhUU0foUXFbfPeLnndaVvkBH6UuaSNyIaGMfhH08ZLmggFyv/a
oWTBnaayPsl/G4WEe/UhhkTDeXp6R8Sx47I8ffNqkCbOUj7DYP15Nq5s1lInnV+0
MjfbHHntOlrF2oJO6r6DphgC6GVmSmWRk9OHfYznbnROGnytE9dsHOejYNbzGXbp
d6nyPIXPcI7wAWpwFPaIKJuzYN3KhbcwP/akI5knT/QXvWvIpL7N/mZSF4w6ZWb7
hzet+dkubq/t6q/G4U7TKkpvcXP2VBvditCtUf8eczDBVT4RLNcZJrTjeg4Hv1Pb
h0zhmZWV8qZdV85rvfcrCeHqN+wwoTfNaGwfn26rz1ZAQtHnnC4hgADXlJye92Xs
nQUssTanYd9AC7Z9mrW8BRBNHAdnGBQFBvCJTuocWml/h2rLcuRjkfzWWJJ3h4ny
QCKFQXRAstTwnsmjtcnt+Vh1ATYxE81XwVZ0tJRqdNkSEZsLn7u3hvGi07Yw+3te
+PNHyQttIXRuwHlKbAB3VeCkGOFmGuXX4TF9iK03BacOm1DKO/d2bKYSboVETQ4B
JA4r4nhZ9H3+8bCPmmtDP+5S2g02dqaCKan8LJKJP2eyF1ZObdUCCtuhLzzd109L
TKEDPIu+2qW8eYhjkFKKILTvkK0O1d7/HG7h07y45c50m5bUr696jM0OxKKNEd1o
eKh0u+kAliO3BPRZP7TwjqVfmuyTJs29vAOBlajDuQzVyYp4iTFeHU3nbwcLsZIc
v+N49j2DzP7ZIDJx28UcP0wypplnkWMrJHnhOfYw4EhMJXrdf7UVyII+6aM42Dgu
lyrooc7kHyaN9ecBXls6iFILjenID1ITl1DmH0Vf5dNfM4KwY6TxV2oT+PXHirRo
cpEx/BNxQptoHLltj9lw9svmVg3KeBTDw4llAO+n9KBvR4CA3vRiOF/0lYRdd2fJ
MSTLZ9ENl0g1+VczUKQ18lsdDZjOd5O1Z/5hYkSUUGL7wGCTyEvlZSrjCIU/KTjJ
/7593M29GQhQcKzTeAeLMHRuXqIQpCluaH1mKcnpreKUAdT7r+7LGIgz4pWxgisp
HhAi1SebK49NLfhegivieom2El1fF0mVrJRMLZ4AdRpvVTNKmWEbwv86YlCAs+uE
ScmtxsbB3WCBPOzw71HGOQigQbdRntrXykyq9MqePsSBQdVeAH5qjVLzLZqBxa12
zQRuyqzM58x6SaDLdt4VAXVQ0miTWUGK/rov8doFxwieZ2/a2DgDkzuIyNHFZlA5
6Q8u9JkeOJ/Gu1qiWclc1G9YFfI9LCibTrLC4PfCSVT8jrndqcnexTbTY53R9dlg
pV/2K467rJ9CheVv7INBa5KtHnEwKPfKtPX/t33N2IL8WTMxzOR7eKgInlnyXEbX
s4NxGUNUttbTIiDss8f1Y6BIKZ2I8tifyWAEL4EBSXharSFldLOJZtf/aWvVRrsy
eXJQ4ApTObfShhDi2j/7s2X0gPnZvHxNP465aBzj9NdFM/YRGCGLDHBFzbfondAF
5vZ1K0QqbvUwYKTGVxqHDMQVSJEQXUpB5G8oq+E0NQo0FYcxY1D/oYCWbgHNRsfC
JAUN3vDbIyc0QSvVpnyndLZ3+OP75S0hg6hHREq4HEpY8fhwU2W042hByd7w6Xif
/LkAj7OxaUqAei/uEwxxMDCQqxaeXyjakjxsgB2Q7Z57ExWNYHBVhqtPyU40KPQi
kkuXOj1ZpZ2pX/kMrTCAqABKSiOVqSL8EEjgMDMSSBcibl4XOKSciaL5tm3nK5h5
r8B6jFML6AOxF2vJJD2uk1xBraLhUuRGUZU+y07OKBu1E9G4c6hVfQdbQaJauUK1
7VrT/LdBpl3pVDyzFdIoHfWS0nfb4++EU2Z5z6w9PQI+D2KIxxtgWMjVOt+wmIZ8
1IHA+YTOFxHO1tx730UKQqPFUerb58jHVEZXms2KAHwFXHPYJ04b3R5hkBRqeF7Z
oZWZSCLOaXlc+Mo5moMSNba++iSTDAoSUmuKPJgtuO/+u+nXJ3mMquhZsy2RMCng
qDBkSXEEqnY+dgtIrx+7HP86t5N29rK3p/AvmkhNMWFuGvbRZ5f/RpApgEKriTPr
8Nk5i7iDtEAjMWZ/hg8jeLnq3zRPx4zn5zjRML9SYX5zTa7fhzD8sYChZ4Lc5JcF
bj3eljv+s0taBfrp1HRb0l/5KPrP9qeeXkxpWGPdKMHOcH6ZUPgFA0lcTQOoS8QL
xXRqE4hP9TQ0v9EO5H7h2viHE3pusBjtAakJ5tF3wSNdTX3ngc5cEEtJ0ltz8m7L
RQnkAkc7Ef6Xgzjs7qjg9fxo6jkgVutOqG3WYREI+ENIfhT/DqbhiveWS0E3ove8
+wrcg8tNkLuYW1iOgd+XV0BiSgZtD8ruvKBXDvTHpiiUEQbP3B0lM7Zd6JJVyl9G
07tHFZ0HryAHEc59XX/3CXItJl/9NkkSXRAwpdnFXS7Bu08S5aR2kzs3divU6kT9
WW2GYqGAG20Ku3h7Oa7Tfr0oDt6RR/nLLR63x/OA2MdidycrGbL+BbHP3GN7qkCl
AWjx9gTwMnqygKp1etxgW6ZKpfWg/5XeMEdVFWkAZ6XT/CuSPaCJ6FwimxV4B1hJ
334+OVvlOIwS3e278hVCvvrlv4ZKfpsDABgj0Uf/4g/SRMnHPCq4KwvqeI7pukHl
tbenm5d7z+NJUvb/pbOiIdOJortDHjS1kqRQJPgA+GuAf5se7LmskK5yJDfSYP1g
pCN0tX81YyQXrMtmdAAIEmUBoKicALDkAcviFgiYczm9djn7Ugfit9LJA2O1z6i3
mNv/C8bINbve1slx7diXVrzJwn+92Tndb1dbZE17SrBRG9j7CnEZeNDGMdH92Ejk
63SL+w9yj89dxKcWqxSMjKKvbe0z7cWzAfxh5E3AoWJyUXleYjTfk/mpl1Bwfo+S
FKgI3ndcBYy3t6uQTv92JuANfMi6V8/G7F6QRQamaR/PfiGIm8j8wFttQBSAJKI/
bXGSamkVI1CdX4Z8Qwu8zlHD+XObwnhvLT6iCww4H/Y6nzvW3PszTg6cAsYZcnK5
ZYTkTQrhGKa+XUyzd2NBl0Hry82gT2iVFSRCNd3zglub4VbSL+PABNBMRhDYLG5n
fXW7hXbaX2sSX30RP/ErDWqHPmV3YiTYam4x1jt6CQwDMlutQ5zT173SS+2SlEJF
2WyAhtmB9Lhgr+4GihsVfY2VoaLH8M5IlS3H5rh4i+Fxp1PpsU79asSIJo+qBC1G
WGkERID4ilZxDOFWNYhScySQ17AqpfaLh+L9/jCpKYpHwqboq31DdEEDHfulbo06
BjpC1Ni10lgClWfRKXZMpvICWfWIMUgK70quh87YAbwJSUu6kc968T9ioV9Dsd4+
SbNFzdmX9ADqm5kRQ7ifITtgmSVjmqCmh/qVaFiaxYPimJQt+Qoz0qF7LKs4Ekke
dKIoojtzST18xV3tKVDlXs2huWJgo2VRf/c+qf5gLd9LHKnxEAJiF0GOYW37HmP3
29n01DfiP/Wu10Z2jUyf7fEG1TmCAFExY/niYOv183n98drm2r1ylg7gBaJoJpkI
G6pFqd0kH85zWOC8UnfFpO4KZlk/EZm41CYkA8MlVC1CFGh9FNzh/L4PQPzDU3ol
S0Dk7xkCPOY/W+iljX0U7Ppioo5I8yVMndJLKTyr5x9k0uCQc75wOdi6wLZweHv2
w0drTt6uPfyU4wD5oTNwg0os7sMI1lx31dkAZnuWJJIIuYZJPNq1sFQaIOhrUiuG
eDzjOj09eMjxqA2PBa4KzSX4Tm8+kuJ8LR24lXEAniIF95JfMC/Frfxgto78p5vS
BspPsC0yMjJOsiU80tRE6QJZJoQeeIJ5naekWsS9fP0BwbQAOal02LmsbRfpxUFI
WsFUw8YatUigiZZ8O1opPDzi1NoQLZBBPlcbyV/WrX0J849bXzrLNZBnYJbvKAyk
SzZGMgAJQAgso2Kwze4CdlDPSX1jvyYvlYGtqnGSaiStzjf+x9TCC/sYNd47Ll/3
m7A5dp5sTM/0NN2kGPtDqd4Vzqvyl87DKxxQA8RBYd5bRrNDsvQHZQYKCYXLwDNZ
RWM8DSNWBomUvhlQN3/ItsqokAAAS/c7dlv9q7shtyfSB2HTW6FIzczLWzhrIHle
zMyOMHiu2LRb4/D2sAORE9aclRC1xC6vWUEkTWnwVZPV56TR1OV3EhThygVvwPLn
Qe1kF8rJnms55H1ZcLWpnD0EdhO6w8AiDUI30X2EqeK4OL2gjMDXQM9QfS6mS2Ac
vG5HGE3Vk6zLpWnmLCtxN11QAOkx90VWNmfjpGk7icaTOrgvmhC/CABTG9Lf/DA0
FwOVi2ymICtM7DIXExK8aJahGPj0SXegzQl9tVYO80YeTdKU0xICM5Jx89D4YdSg
wJhcZNtgP5SAWt4GI5WgvVw4GdvhLBIZ2LZSgyLyL92EDy9bRdaVPguhr7A9whaj
KfoQDNZNVqF/kQ9go2Vdv69AuN5u604WExhFt3YcP4UZC2UTBwhZoJyzltqjhjTy
ErA0ZPqF4iO+JlQOEmy9JkY/FNeFd7acdkdWr9+Fe95K0MwH2GdY8fKYo972sWVo
Fmnjg2arhVjAzXZCINVtHK9B9zAxtomsI8IpEJxjVEg0HMAqkChPjk2WRvvwCrKA
UF5HxemOoWKie833VMdDkg4dvXJPWb7zDl99A1Y18oYHyBPY+NYzZCL3R0LHjdm/
yBsN3C8a1fXLkHnrjc1CsVaySqih5lqbLcTZW0CNu1ODA5hLZUp+sSu1nlPorxh7
SfDQKUT6FfwZ/pHlaAmkno7hoOYLn3LDNJcvV5ugpQrsz0wrBsnJt9fB3czELj7O
eEpYGgyB3MMIw5DrGix3c17INSWck4Xeu4WXnAYQcA7wiZznVj1vBasGoWePdkgQ
/3UfZgoRj4Olliy8pECxpmaKgoOgWfiGS7pv/ndJnGrFYvgzFlezOmuBVQqntV+L
iOcVtNQX5Coeb+29/a/CDokcEAFYwktnZOvNLPXA2xlOTPLPEkjYiETQaD9gW2xV
gRf5x4+8geS5ZJOP7XueJGIZU1P/NrNcCPz1m4iAuy+9viJMYSVyc6WD6YE6EVUR
jQX0edAjRoXnbQXz61Fwie2BhD5n08seLYgRC2d7GT4fXKh/8zh/SqjBb2hWHmUd
iEtOrk+dBHtub6u1OskYs2y6LyVG8p24a4WuuvHiFUyG0qUyUukwowKBgPgaV82O
8wTJBjJZDKegTv2J0jvhJMFYUGEHcTkMEM+StyFUfDIgKsDiayRF/yYs2jOgd4Jr
QUQomFLArEj969Xr3+eb+c7qntabPaM9JpkkuxrNSvYLf62kGBefVFq+MgbDtw0M
ztTi8LFO9dDAcv3b/Xgrb5PdbyvC6RHbjJOhouiRS5xkxWLcCyWDrikErFDwnLCW
bicHQWJ8YRicbCd8ZYGGBUBNfqYXxMJTDD8WIAd7qjrxiN0ULykQL16g4qmrZCkL
X+JL2LwfTiHnprCKP7/Qfo/1ffRa1iD6vAllLM4bxEfLRiEmZjycLfGX+OIm8Aqi
lRqdcDrOojeqH0vS4M0NYxEVKxmmacBR09lbQLoyW803kUDoJYIwbnjb1tYctZZe
FIBkFgh7JuzuWlrqXY+mS3XSGU5ZdoScLSkgdZX6OOc/actul5s+uWJYeryzskQ5
NPnMQd70B1bdQbwFkUmB9IBGHAeIYzicFBax3ml3yi4f6Vy/lcWTErgaCTg5sQqq
bSjto3/SpPRUdIory1oU0e5yLnhtG1f48bnnnWThAHXQcAB3W+mdvmreqA6jyTho
L7OdphLAr+dPVqgeDu5dqE/1hf01ENRgbxBjuT6LtkZWSbpsXdLE1G4nR34a2pdX
rfZbwyhB4bfA+oRPEHAdsqbR7JySUsDo7R37FbMRh/BFgNmAjgzqxnQihYaOVBOw
yPvxQ+Mf4+JUSPHp46iA0Lahzq5kPEMCArYlWSdnpKXn0cxM0FcAr4Rgy+tWUCah
8jny16y2AyKU88ipStWcnM3ayKiKJao6gFalE1S+Xzt+PoGf08Qr+A9d8QDxbhIN
+6rBHeSVZS+QjsW0/P6ve9HPap21u4QaFMK/cMmUEJi17HdPl9soaq+4Vn2z3Tdg
nw8pqLUrnoiVKtE1lUYUj/mdIeop+/IEj09jmqWAl/LU6xu2VybiyM0pUA0vvp0H
NHj6U4wf1P/Dbq8tipz2VMVL6BsMMxaAJKNl4XC87g4mjPjVTh3Lx+gDGxW/Gw/D
qis9IpqMwJhqfht16v3uffW8o5xmMpZfEnfKBzKFuomi/UJpCZvNYWqcQ6oV9reJ
HGxYW5NoNv4qqSikzsbkQKlIYqDwBb/av9wNEqg3rJMbTSrwYMIBQNQLQDw8fbgR
6ftn5iAn6+Gx6buTVCWH5ifoJSFKi4/FxVf8dJGgpwm1dx+XIigUURQ/jF5c42G7
+EJdfAeQnnr7SK9CRRf4hJqv5jKzBuJFUrcB9ssYWKVRwEyy7krknKZoQFdklDQh
ogo7Si95xeEagO7VPkNVJ1vYd3NzDT4AQioHZZLBt1EF8mqj7Nfi6m3lqqd2P4ah
/byJeJCANJFH30t/bOw42SwZsDPhbGSerVhgm3ygSM5xPQXXAatmj6pR5c7MdMgo
s+BfPR3A6QdpyJXrAvMtMqpPxe6VXL4/mlNbZbHK9hC8tWCaHT6ogOCN8wBEJRS/
fupdhno9GBXlFV10MBHl5nmMtm73LPGEmkDU9VLU2H4XwPu/O3xXYFxru8zuu9OC
ARnmg1zy34EZHHM4k8w3BO/5T6ZfcqvkJmpEyQQbPOEwUBzM39FxVrQOJfBB+7c8
piSRKe1nw/jmZUPFTN4G11vet5lmmpNlna/h5QAjHl4nKYepQNjfFRTq7d+sK+t+
sJlN/3WSShIRfd8lvl+4/VeOQnFRMJWrP47I8GdwZu4zYtX9BFPEnabydXfPXmAF
OAxqbIz4ZbHvC7bQ5b6DExFghqLChUsrHBaNO0T/mmbYHveaOxiBMJSwNRLJYUB3
+YyOtPh+JE5979/bTtZdITGZ9SkS2TrSLby+aDKSmNcbqTynm5AT9ewdq9o3EOcR
zdaaoQO1dbnE5E5dx9iTEKE05yJEai0spdHhatFhy1CTUonVlnuKnT7L4msOWWqU
7r85axdYELGQ163cra1Wa4l7zcwqVs78C2Swd1BFOhmGJOW/CKICiOTWesTbkzH2
2Op7zsY9PibFP7KnoUF3Ahuv8+p5l8UUcsHR8i9/oGrDDXfJktJnfFXdlbeeBGNc
DkEQ/PkaZGTJraotcpqYxvDPBxfPPSlIBAjz93RVzZ6jcjSvKuyd8uXsQ4XfYZMl
C4I6k3N6Uc4M3Ozb1TH83YOISk6dYbrzXvvakMIpseSBuRjBH+BBTWW197vCHDOX
1iPb8GdcEpUeA6cTr89BFraU8OFLxPPK3qAl4Fk4FVBTGeW7UgtuhzdZRvDbSdLw
4Zsww+xkSBcSZieIqZ6vWx+kJls8QPh+aeviSjNeANLMRLJZ9KAkRuo7VN7eM6v1
1jGeJBmdaTDXoFKwk0Av5WkgxFHtczN9QXMylk73y7F+OCxhjoyAmWC7rPelEkut
2SPSyXT3o2Ax+8cydSXMoNpxBxfGNnIblcPsW4CX/5zde9owsLkSMnpmKbUca/bs
AOHJN0BiDUG08jFDGjISHYFrxez83Dg076m13V2PvYb6oCYwtY1Ky/qLmkm+QSme
tRbJFXuX94mr0VSBK1uSdFZgSZDfyvEJaILSgKNSn4gMO2JRErVbtaPZxhAjYNeW
gJGe9bBpMTmssRtaGKOiKYaJT95Ivv/2vN5udtNi0E9YYJVWiyDFeMJjpP+mSlsU
TX1GE6W4QCpyjEXi2du3ZRkPM9qage97AykfT+fZ07xyXauUNaJQ5SCXVM65BElb
rA8rxAUVJLMstOYK3ON0uCnGY09Isk9QhWhYyVFdg8O40hfFiFYJy83DG1Y5DMIo
l86Yucys/agbD2BCJJZCpz+rDlVz+2ZPwhES6yBathbgKGZSNyXsHHB2VYfWIZ5E
HI2zIkrCW/cvGACTEVbqxWtsykoqw385Erv5o5GRcZ5CcQLvtTedOweeLu0i91Tr
YTp/LwkMI5WX39Sb8/kz5Cr+5zwa+hJYc2fJOcvDJakDKgcapb5+DkSP1JedH4gF
6Qj2j4Dlhlj1tHFE65nnIdxvMMvsl6qtF3S+o1/uIHlCKrpSPX8l+GiwUA3FHNs3
6ThhdMaDAudgsnO5D6qZkpD919lHhGSVBxXaIHcJqhpE5kbh2TOY4ImNleantM2W
75Q/XWBAq7xWZ0wPJ/eltkaxNRG3AN7XuCntfIDK0+jOBvcha4P4lL2CdgSu2gVf
c+oDZRCXS236NRdLUbioPSP3tBnClIBaV63UyJC9U/OSdvgWRfs5z/bjT4k/HXAu
lFuNcJNDsXAmQRF1p5CeqIkowIU6wLJKB//tWWMsdFICY56PJ+mjLTO0V4uSV6xF
RU1zjOtsOAO4EGjKcMm/YU7PC972tOSe+PE5NTCvt2JU5mAPoqShKw/wSe190Sh8
VcoIMAvkFg3ySdMQ601g9YIogImWIjtH3Sa40f/TrqQdeQm0whVw1TATajvCLk9q
dy70iGZcgLZSwoFmANHXtrevJm9wPhV4OVo7djul+okdstGnu/dL3amruCMJNQt4
YFZJJnV/2/PLfDTfSd852b45JbERfdz+Zwa4RKf+XbEzlkh8Ixs+5yAluIWxDCRw
4OLqmYwk8El2fTPGeMT+OdVw8noleIxmvnuE3UKQnE+tPQ34Kam1ztuT/NNS+rof
i4zl2eKO4tmiUkqDGcjnX0bD+HdwZ915SrXYOnbkfYNvsjwpxEMdF0nKbePNo5Ic
nwi7OidNW1X7jwsX8iXOeGtKMR0KqZFgV5WrCj04GOb0eVZVH2YMc/D6AJwiUsI5
XHpMWC6o3jfUog+hRFdDcbh4VA5u+3DI2TdWywvs9nOQzShN4bVB9DV2YxvWvL3k
SnDLDehIc2nB97/0gnivpba1dhbwTZOjbbIOzpc7qeJK4EPlI3VW6wsr9VPedunB
hLSR3X1ZVg5BRSN5uWEEyHANNKcOJmSHbqz1aP/thL8LoY7IdHuO2g4vmmt4R0/w
7Dw2+9f4f/41/2vfJRDn6doxeOSXarcz8iK0fbMz/53bLHYS1LImhvw2vE65gif+
dP7mbri6L41se6HuOnnL9apjdnPpsQuGtrK8DZdB49brpP2dyrB9Pz44j35Tjq8L
UufxKoqPiUX2L5IYW+/C/QY8EF2s23gWCHqnnM0MyMhbQAzOGA/hpqDZ469oY+YL
NDsEC6r0Svl/7GhhE1OGOS/aCbCT7CRnRM7ZALyxd83bd/LsZOJ0dhokW3kO9cBi
IoTSbtA8jTMvEkH5FgbEQ5tevTaCJXO9Ot9+afoyIwsCE2UR92obfN/As36OnxSh
OU0SUbiB83Rzh4RT0W5x5FDzp01bIOoxonOcvMYZWpLR1s5L7UkkitEWNqBbiPJm
HyNWsYWay+kNRUK5h2KCgFkrnu2rPATdcbjYwY3pxQyGqm+wP8PzGLOdMZcDDAWZ
zcGaj8A4h0d0+lMFLjfx0gSCO3X7JYVX1N8C6XjnR1g2bwT2NixqyDlFcIo2Z2Pl
INWLCBFNfaxAQbGlzawkoS0ZeVe416heKQZBpz1kltKZbRT3xBkpmwkzCJjm2f1c
wzp33cG8IChplFIjmCPeAIU/TBpgEkqIHaUGsnd6LankmNtFVLp0y6pgamw0uiuB
XfHgCfZSH5Ky0b76CdNtkZ2at5wTe0njjfkw8ZPzwYGDguOwXM1en3WzA5kwBIq1
FKpZInWeTYm1c9G0zxxHRcCNX2IyiOuaRVZAGtUOqcs2nBubqOB5zW0sTSodx7Ev
OEHQeMeX4ee3BI849MKZhaXxy1KSQrR3LnzD9/kiCDxVsAl2yXgLQH+Bp4zKkpg8
4ktk1ZngN73eXJZBJvjjcOqSPzU+sUlm873PcV9FKHK5N5q+7bXUVpfwtD6IccwB
lKzD93PHSIgYRNwZLzccZS3QtJdXpMoFTDv0Y9/TxwaV7p8uKz2K6HrCqDknbB1S
tHmuKq6hYXV9eFofSefUepeUqc5C4jnjjZ03YaFwarNTt7VcnDx1cfssnH8DXo8E
7EvgtG/Y5+GrOED4VDwYV1LPOh+WFP1w1PYu2F9lHBm2WpQD7bkiRiitrJkm3/WY
b36EUVCRTjKXacnA1FhZGrjpFTH8/miMZzENlVhvd58mv55Wq7Yb9U8srr3Wwf8v
skTTTPY6P7RRYUdy8FpOQFlqO95Psmlz098aND83L7rvVpMMvw4r+EEwy6v89Ea1
vE+EPFlZZj76/ZBhbx8c05fh1nDcPG4T1BqJEYnem+jWSQyL95jXw3u1zJuKhPin
qEf1D9r2ih/pLm/DVmV2h8Snt6e25oBfHcqQs07bWYGC4ni5FktuaaN6of7R5Bsh
J5jQdPXdLzdEQndT8v2KbUd/H4KmilzZIVaE4zvpLZxlLpvCeJuWvxTF38ehOrJA
Jceo9OyrCbVVW1L9gdv2laWMGUByE9hFoHP4Qn9d65OhYDqjpAIkLzIdjTsP/6qo
UMV3Ce/uegZGnnEfmj9WLNe9DZIhKVAaF2tf9iVodo/1SR5ffZ0GuwpoUrSkkLBx
JFKCtm5pxFSgZ2bWzq9h1M9neIsxYmZdlaGYhMZjKa1WJNgrL1prFR3xnKMcKMzp
i4pjnGgHbQspWVFWseXIQeSZ2yFTXOcE6QXFfFZsBBr/IN8mj2xSuqwkm+9QSYVM
kBiuPpcSQACAKc1dVotCak8/Xu51XQt7S7QSkr8BcEptaF9GOz95Fdm3Lu2zguqu
pNBGpMKliIL3NnOY3okrTomCkut6+A7zZEwyoNE8zjIY9XqhUjyjBDPWKnLsaF68
okVIyemLVFsPG1okbOKd7iiC/wROr/wmIOaw8JkffQ2gMig5BT9s9F5eLCKAbbva
MEfu3UyZMKAvi2l+CxtPHDgJ+oasWq8137byzPN/+uuevSuXRRuTCSeLiOaSxj9X
nzG+7axNgkTCF5mNcvTG4gUpMK6ihCB29U4Uf97/6L5dav43xpbIrhacP7QQbY8L
B6JNrLV0Twx/d0YwPWbu5gDW4nC6rAuveKQTCm9va1mMtVlBLUqW/OwShWp4nDBX
mnf/9s4rO5cb0fiJU6sbSUE047x0durkMihiLBGZQVukoonUpB7WdQsY3k3YaUW5
NATwQpY/SmyvHnhnuExnczn/GRC8d01SUDh+tC90h2B6I5uV3IR4fCHznvjwin5d
L9k04l3EuQLdcOXLGZBF8GjYm0be/whxzcGz6ByHjJhMIve3ULTcuFzB4pkpYOBZ
D/6zwZEVx9fqxd5BF6HSxm8IgIHCeH9jjde4aeOayOA5487n23M7FqPPrfhX6LTs
crPDV7zIP2+KhGILBFcOOc+nRoAWTBY6rmX+nz4H5lNswdSe29B2j0tgFerEMIqg
W2HHwbWtsFVZBBCa3R8H+iR1Lf61Lj+FAPK7va7wuHJ3i3XvJ8ERUgKbom8zwlVI
cZ2EmH7AdthNeQbiGCxtaLeUsQ9qBcexdQ2I+4GGs6aEfrrMl5dxgjSIjnd7SQpb
eO2XJP2DuZ/jISg4ARQLWCVSoRynVR02P7ZVvyDzqS/i2t4yC3mvdSW+1bUY3URt
sQ2e5UvAOg3JUp706LgPza28YnIwUAolfslmzA10nykIojG3LUqjrSZhIxOcCV8l
/OhJ9Ax5MZ6isFwqLzcHuFypkD3BTfkhQ2qTptGz61/JJpNEw/2N6EGeTkUQxV94
u3ptm4MaYpLDJSF/A2HmlSHjLvsl0Yb2kmMd0eBte0m8nxU5eNMUlxYOmcvy50Gp
/6EwFW9hE3wOXxcodQ6s2uUh/RE56GUpOMATmKopIwIfnYNR4xX8u2vJCvNXJKqB
Pkw/6UnpuLi0ZS2gAWsXVo0bVh4hQJ/3zR8XjkfOgEZKHrDOAiy8vFu9rnVoEXBc
LVi0wBO7H1vSJQ7H7LnaAxh+dkanPi5knU2S+c2U+RzpNGd6s5QwUQyyea0y01pr
DQEFUiOStZtAhXJcZciGdKcmJ63mwby3Qzq0JrJkMdpjJ6fHmzqkMd0Cyfq7+Znu
hR5hgJjYE/pdMUArPPRQbTTDNaaDM4EShT83xBzzGIYtm4Vua3o7wxhk8dLnERUK
cgyVDWTcfosOgZYC7fsaY29VFQVAca97RCVE7UBm9O20yEnpHnQr5D5k96pgRrdr
oBnJx/+cV/hYAHZPakL8NV/vP3HlA8KpG4WFW2wsn10hU0z4BKT275I8UZH1bWqS
Ez7M71XXrWi7TyPekX7pafN5v9OBH0tUGpk/A+rAVWDgA4E/udHNGqhEzGGS8myS
14XoydeHdMk2kpajwifINRzOZosrmo5SlnYgM2WKsnUzhITZUZeD+Wyx9acyOb2O
ix4WaXMv8B71Fw2dSM+owodtDIIa7fadWHc5rBzk/ZeCaZT0DJSB5HyEUS5kFKec
n82vJw29xvK5F7n6ST8X2riw+2vCAClAKmvpa4JavvcFuLFcq7h5Bv4xUV4ZfNgS
TGalsRtmykRNlVN9XkZUhl0jVJvCHWOHuzUGvIIXjcNqEMoVDg8NxcnuVea8FSpX
BfEKoR8eDXtiyH0NZfzc0Jyc0ijE1jDlphp5lvAKu2dyv+deIaXiEX54+Ne3hF8A
q6vXCWHP6pzRnuGQBU8Bpkl1RN2ZqwEbKeXJ4gjR5k3wG27iFJ/d60cU5HFXuNlb
qiFiqlPQWrbCl5u/5oSBrcHyvzvJqwErPUJLwN/WcL42B/n19C6GVT8HaukMB13A
wkEZzAnfTDblS0uqY17ApCGQelzTDIF/VNSEniAAwZECZsHBC20HLGuilGlrFOOv
WodFfR+4s0Cczolf5ac3bRTToJ7V6NcWxX9sdVWVjNB3ZvwItkQDpnL6zLreCUwi
HZxSkZUvoCMq/eulelupfLeZLk+1dkWK50Ob+h+rzCbnLTwbFX6MmnYfvGFcZBmK
PyWjFkrV4ZUf8ARH/f1z7MLQ4+3dGTxMAI/bEZZWtYcvLuugxzUl46WVEw9o3noB
RT3dyRSBpHyH8zxh1Op7sQ1B2H43jZPp4BwypvwDk53709+LDQXiJ+o4wIsM4LSX
PG44LWQq+/1UZK/XCgeKByGlvRbs2RJAzOpki0rzmfpjHecIREXE5WW6xin5QJcl
JKsXOxRpIsjViMy/CwBJhCVh1xjFo6mXhaa9InwJVtl8l05ro2cXMTYnZzd7Tf8Y
wgfhLF92yx+AaQJ6l629ie03NmkmoYVxeLQHQ/ePjbaf8IqbeB8lCiS3k2/7YpOw
0vhejrS2wOrZX5sCgFt8qG/mzTbLvqDEQHsTCA0pSLzp4oEr03rKiKK09dEOueHQ
zTN3D5PIf8WqMziKqRVg84xBgD9OtIpvJjAzEENx+REsfCsVTmEy2fnJxmTlsaG2
3lPsh1f4441A7SMmXwBnxYBNy+4GCoH7KImDDUGvPCsq6ALWpUFfC8KfFWweK/v3
oW0V0DMaDSYkCmfHq7DMMz0krI1irZfbUQAkJgRn786Hy+LiBVCdxh/SB1W3KH0E
bbYpjyf3uWBp/fa5lRIS+Aq9dq790O0+5UfZiggkzSpOxFk4mp80t8udfGdIwCfj
J2datQC6E9fcpvyuiK3mxmKdGdh3MpDrq2j1D+/fu7fVNtuhPHryJO32YQ6LVih7
TDWL9KvWDs/kXROn1v+Vz8S+aDPNCB1sle+vO4WZLSb1hSHacYr8yiwTQDy+K4zC
54C1fUgnQ9U2moH0uxxUKgJyb2/whsZkae5zaKwSaSExsZTVxP7ZfkAP/7dE40Gb
mfGf8miMjzlGZHI+9DmnazlmIZ030RX2KUmlTAR+3PP8kDE33Zj48uhZX9z0Il4i
Op35/zne6ZLXQObJUXsJ2mK2js3LEgRjyvqaBf3kpxX8lH6z1Q2sW2WWMyu0TTZW
i268uYlIbkIEmmF5zImQhd0s5g/YamJyIhQCeXLCYScMkvjSpEk4KR8xRCgEFjcp
mUxFv33XCy2zMtWJIMtHJ3xx71Gy/egjovBSpPwMPn8rUf9aE6svULsgMZqvmDHG
Bj8yp1HE4slz1bIN2lN5y8oz42zW4HZ5jlX8YfU2AumrT9hCzyjZ34kZosliC5Dp
bLu155py5fk3NOQzPbbguFuFjOxf0qypyJApCPtEFicfvIqm9LxtsQ2kdAl09Nae
SUPgDid0y9wnVMeXbK3XWbEXkDwbMQIKm7LiEfW4j0mr3njgEZPfE7YJqHxUChQB
q+ATvu4h0jOV7PZO8OIm2R+8lOkWxj0LuxoyKohkTcuFJC7Skb1yz1qTIZZRgz3A
h1oFMxzkFXZnhX8EklX/OM37bvPYLMZDVa//5paco3aB7UwudDL+oTre0aofVYsy
zOfgYeaIl2oLlqCGx+Q02LvW7gWqslStIsbvu2iQJFsmkxPit1VxtTgSwGNozn6B
IyktxLxkmWE/wC/dm6vGVHP12QjDizNT4YgWijOBffpEijb5xJWphajtGuj9XlxZ
jFfRL1RYDViwJo3SJXG8N2XFWNVA6d9scphDoZEjDDoKfLiqp2G8PWW03JWAMIMv
mPQhHPF2J5oyUOCzD4HUDoEVxiOcs2Oy3afDfz0aU5ncekj/jKtqTX4dwZ+olFUS
yzAx7okTdlQHnTaAsq/8y8EaBfPyqoc6VQ6ugNk0Ax4j9Zti+fl7BNJ0MiqN/DKp
O+SXxA9JVFVeS9+gylKV6HwI+ehOUBUfybld0u5jiXgggOV3YiwPSBEGR/LWfA1o
bA8MJx45my5x/Nih2fMddjYJShIKppDy9t/MaLo6QrbDWGsC/a0JcnzUWvJ5Q1Ez
k/DTD4SS68s+kxEWdPPtzRODVYuBAAxVLmjHscThhSIVC4hDQe6zHfB9ExtqQIWx
EGBw4u2RSO68oGhgh0I2HArjHQtagtrEVsjyW4ELxdrQ2gpkSUvmvUQi6zESiebf
C1jJoS52ACFCjVUJ6h/u3wOGU7a1cIk9qpQcSY7s9poPVeh404NtUL+wG2eDXqRl
0j1iR2vIZDTcFNPbRuJpwzaXaneRiJfawVUsA1rEs+jesIkH2vjtPzGlGuJWY35P
PgF3rwTUK0pNUF3ONqbN5UBKm9GTlGoEdBc5Vtli5fkNQx/ARvcWI+XaTXuttv6B
41shZCYcb72W14W+4l27xXniJsOnOxOqi4X4bpzqaD2oV0uB7MXQqfqC6Cr4I9wq
OXS++OoDTfsNkLqjby/6V1pZK5LAa3Y8DHRZQEslMSxQGbNlAqBCKVLSoroeh+JO
9xUygLsRG/2HU7GIgZ1rWtY0YvIcOEcnH1K2vca8MiU4x43om6MQuFmRMmotAr1C
zW4bLxT2eS/iAVZS4N3v3BaXSGYyX6EHDREvWCKNZqVDNnr+3gMpRzrfElRTlJVr
BSfBeRU4+Zw/LPXPVK53eRP6VdoJLkfTMDtxFQOvrM0N4yQjCep44TsY5MQMQlZd
89kLuvo3ubNMfOx3kM6d5BaoCZjtFsktyKosQ/VlCn3/kffeBBTCGNFk2pXXacZe
tGDVhjiE7jhmk0KXEnE8hqBCwP/HRicSSNH7XC+HfiWCIyEh6Cpe8fyykUJ4CFU5
yVjD5+d/SNmw9BFU0t/X5Y9Ur1aQxDuPj0uX9Qc43qBCZlAp5OQ+wBt2HwnDInmJ
tHvAq8QCq0EOJqRV4rDqbf8gRmEePfsPgmKQZMFqyoPTIxy3J28T7w1emiyApKit
FiIVTxNivoig11w0dx7mg3telkjaS/WD4u1u3yPfzYWY9Oi9qEP1wcIxU67xjS0u
KbeiuMJCWdoekrxXJHrgagL1k+3f/Kk60rHHTDj4i/xfEfUlDDutGZ7/uggpdsOD
IO+iZyWHgm1Olv79nZ6CaZWDyvx/4NXJAKAbj+hdoBL5djLGmesJMBQgzqSRjBKh
XK7RPdc+hXr/uRE42GqaKVbPF6v+YBmrX5K6j8ivXwNCPaZJX9AFTvtddeVOaHqc
nhAChuRK/zCwGpaU34H+oY8/t1UdLU9GfZTGX/JnqNPxbzTmOFIw/5NY+8DGxkuo
A2oP7AHlqK95OsHiVxaXD8w6G68s2Y7lD1eRogQMvO4StvahGo3KbKIPPqDzQ7om
phxm+WVT0OHdmBys3PPPE9k3f+fY+47SONH3Rm8jxZVVX3ApCnpA1ce+FNTifyR2
LRVpCNDhMkV4WYjgX2r4zFCjl5XKtTpxrJxLk1uKrQRt3sQ4Oh+H4gd3ZOOXrjhI
JsFCEvGMdNSss4lNp+evVe16yQLofZMbNVf2mv/ar+RfLk+pfxec1jzVAYzOxLKX
Dcy28USNUYJm2KL8iY4+yzB4+8NqIipzeP74SEQkQs7GsXB7iTYCIfHWYYg/1aqh
sVwXamxH7ZawH+UssJUr3RWJqoqQTSuK3X8vVZHBW2/zJYajsBFqf9ZARp+YwalI
c5dhXJU2e5KtfVqSh3Ut8NgAcAL15zp29RB9GB9U4rYgHkYCF2UhNxKVSHpmVP0a
COUtj3w+FM+eNTdNLVOjX+5V8qzpKCbi9JgrbXQKKuONmFvGn1DeBwSyPrBJnarq
SgiQ+/wb7GGrkTVzzHy2QmwhUFaymdmhLlIWuH7+ozXp2fsTs3LWtsf6mz/0JT8g
w7pV5sQb0+9plzz95p5qb/vpMgPn3uGlovIes8WjeNxlN8qnpTbIIAD4bj811Skr
hD3ly9VLc9sR+VK1py3I8Bc1fEBhrn9fL8mliDBiYZ95yi9uWvCziwTriCAx7eA+
OoCPgbCorayAgMPQzQeyedFzhYMuj6rbvsRUsmIg64DSDKat8Yi028oATFvCzSMS
EHqsqKqsU4NUpPjJhhmO5EAD8vUYTcnaMPTCpP4x/HaKsyQAh03RHOhIaPadD/sx
ZoM7mQN53n0q0e//46GvJicmenfeGL9I0yu+NbCAYVYzcJVfH68N0TPyqWqoprM7
w9Ml3rACjpXVDwemazwO0AVtVg3S2apQUg/Qvu+rb+vfHK3/VpqBAvo9UMJk4zoL
b35zT3OMyI6UUJ+varsUKBP9yEm5CiwZsMGLZHoxGwBMlLy+H3r388hVr03Woj4D
/0rz40c1CFl4zf0PgLvZI1KMzBNMM4fwklhV7+aOgQ3afq1lrv4bH4+/BDB7r9S9
JcRz3jfI7Ubf0ivd6RzVgvOMcIKczhwSNhh+X90K6zossRN/CaKwnwn+nl00ztWZ
qbWkb0rXswDWyXfiyQ0k9FdJY+SOiR6ggCbql8dQ1DFJhRKJ08L/O8kUigCp5nlF
DUSTuMuD5e+ALX2A4HN4jB7kO0FQzC5yXyXDDNS62He2aaTErlsd4DwzZAY5MNTM
IphFoOT5sKBqrLuNSaP5sfHgvh0X615obyHxtpIK3iCXin4YsnU07sf2Dk6j1Aes
phQ5MG1uxoL4+x20VBquAlqYnhFloG9rpBTblOhD4ZbioeYygED8CTGt7sqI/UUh
LWyDvLp3uJDjj3e/KQo7DSCTDQ8RK7CVvQIOw1tX+kKDatYCsPRNtt6Ht2yvwMFI
SlpKcfauwsWpffwmFxpt/3iLhU/30bqbyETqSkZZhQConfP6yup53S4QinFv2lOR
EVqyS0O/A5Q4RlHJLz0RMSLeSseI3uBAC7iNmXU8nQwCmhw2tJVVYPtMw+RCEBtM
05oNKnxcZxg71zbAPejQu+pmwx9weoaZ1TOHVW0wYqiIdrvMq62yjrtV9UJhIs5t
Vtx0ivwXOoK6bJVW8voFw4SYiVxxUrAL/m5c0vOyPw6ue4AiG0h/k2mWvfywOqo6
iExV4xCR5NFFeKLT6G/U2wXC+1yI4cGGxzwOEgfe4KtuQG8XOndaDfZxZlCW7rSH
18imU88zmwXPUH9yyL/TMhzQ3NUqvGlgVG4TN7a7lw7XgbI4oXpEEUk3SA9vX2/w
y6RBu9qis9TueBRupAcSvdpJYw3WbgUDz5LcT5PaS8zXblp2NC3pwW0DnZFjR8pG
mKoXto2zsoFQphCNN839STWfjFlKb/JjMAq236jfgVxTDuFjJ2iW5CugFUsIZ1Dp
fpGVl+6Pnm1YHYeFL9Pz7W/hAhTvcEPZ6nErBDkj4hpigGnxzGq9VsP1qItCiT/8
FfOtGl018EfX6orKl93oC8B7XG0HLCkj0NTAzjMRmQcZpCAtHnw1sdcv6SRVjyut
Xf2mAvCnIV04NNx7hOsLfkJ+RRNJg3jxZUce7Ra3uoF9W7pz7UEqXOmHwh0nK4I3
Vfhgd2FzCSnBQcJzgNJGdLOB+vG8X0Aw987I3yGvcIg2J3/6M0JUIu6K180YRsOu
HtOz52yPs6gcQiYNMOsTO7LbqzPCVvPPi77cJLaVoiyYMHKXxKxyRnQTtApDzYts
PcW5S4Kj2kC5NqEBb/xd7Xx88wrT5S/c3HDDvqYe/ymNs0nspBDfAlfAnz8Ya6VL
pyE49w42jfD8hArMKyyZeZOVL5jlEbkrhcNwnf2Ns49akl2utf7OBgUWPbGiZYjp
R4Cbkn4bRDW3bDN7PqYRcaIKjvbZD0w+lA7a+418VvtoSqGX6sWR18KlmAn3mkb9
JV3EymyrmLfKMgZP9OIiQ34UET2WW1oJ8sr/lM0mk7WUNs7XvfuGj0/NhK/Id5VI
x/MWsM/XG7vDgciPBhZUOA7+g1iZDlVTWk1gUvgcUkWazobADxKYTzPXaAiwSq4C
X1Bbh6AVWPzauz3aIB8GIa8YgcMqfKWTKKQWzSIblZCMBX2d3YBnrLK2P3Hqhmne
ItuEnGXIIQ3unc0HLCpRZC2V7Ub9piyDNNQ9n2CqQAtgfjOleVnfsMaePAyUb7K+
bzFCJY7xHM7zGKOE3BHlofy3uet6b+KGWLFWMakrj2RAGeDmEeX4YKbDLfDTc6HW
XowVsC/870Pph5wI1SdQIIwcfRjKZcfoBF6UotW40BHwQVPx1hlm10ITrCnYB8Jg
YrXoFAS8YLG/LhU3Uk1+Sp+fx9v5umE6FWFJYFS8Wn27dcGB6ZFKrF8v9KHWLETx
gaK5w0rylNobpJnDv+JFlCdweQqxaX8saiHAFYVTS/1jw8cGSJzcLpF+MKFmwsRN
SKFSpkTgN55YJShuCJm7Sth2hod1f2MVwm7tPXzSS1oQP/BNClY4+z/h4/w2qrc+
YEtuphQMlSlDhF25GWARL2sF4d1OoZ4m7OZULt8w7nggMcynvTF3cqPX7ziitxSl
zRViBCS+RUu8BX/Ag5TmjCSogPtZzXi+dGQS1HwJcHUjfBJgRgXLI3U+IZNYgvXp
sybHgO6Zd+ZYt0XlpKxlcMLDDL7Ja18IQ1kR5omnhR+Wvr4AHzG02fsbzqUnlm7s
5Yl+4CSY5jZDOpMGCsKBXEvB5gKeDXG0h1Iq3rTmGdNgL1OlNfGwSotbGYHdFhJD
sG+PLVWHCv28fsUmE9yYLasKGBg7foyKOMHt50NsWx70Jc58f6TyfE1qNZ2wP48i
e6bCCXlgFUaZO6RbHDd0sIkZ0kC0guVuOBvYso2vWuIzBVKOipyiX/dFC5it2EtD
NRcLXy8y1SG0QniD6BGf4K4FQB51sAt8ludNU011yXm98PFPaXkodbs6a+O15p4U
tmaxPnZ8HcfwRlbbKp/8QtXsCY1h731xRLK/7G40/Y7FcT3IrL2Ba6xgG7lL/1Pt
NLhX+nDHuXtXWdjhOtUaG9zOXeJ3EThs+lh7KxM1RStJXxEuB6VMGeEtsqMvonuQ
DmBJ5/wZfgQM91dcBbEdzX/zp808Z4k/Voyl2yX+yllapraC/gJ8OLTL7v3cHGkJ
fPyOUDjwdh/dHDUAaHfmwfViwA/y1Qd9j4zUdrUZ/hA0f0f0GNwO8cHdIyWKXiBC
0QRyJa7uaVLeGGmcuPgsPMd6+LafF7hQkUA6R+pGN4Nf67U6DFKBnDSlba9ufMT8
4fijhZQnfhh9ix3S2bovT3tqSitk59qH2rtRLUCv9XOD4nzsv7IIwmdH7GofdwOx
FFgK2TUHP1ZMgxySFNtxP8ODffbCJQKaeoFG/n93dtGzo0RqWdyflqBdd6sST1Y/
9AN0+fXHBnO16GN4ZVT1m7MhGlISn6ySQkG0NDYzzJxt41KSOKqUoIyXz1Ga2G/b
/6fEoG9PLsBQstKo4s9lCeIKYRohuLjUo/GOlXnI/S3l4ofqCZr0+YXj4pJbzwr5
JfE2e6nAs27mBWwzWrA1wRlxqdRZ0O2jp5jSx48typ67EiSWJ7fTH38Y20M64vdz
W6LHuyVM7comGJL841naiqNh/w60t6JCdE40RM0NbNZSljRxijUlehiagFmT1Tev
ihe64LWkYLsy37AR1lMgyoNna+ExEz5AdTT784Cc+EmHMND7gaj11ItRvXAUiccI
mz7xHJ8dS7pHoOQkfRhfslFYA5bMUAiF5z85V1nBHmTZTMEXb5KidPf5ANm6VUep
HHAj7VyTT7Gu8600kf4NHO586wzqn9Ho4hbkcTrF8auL565iq35CllabqtsqFP+a
clJyDMvRyPIh01OoUBG9/2PA7cdeur6OYZExmVqYcLNDpuNSFASAt42NK2qRBIQh
ZhXuBW+3Zhu32Li+2LFL9trseLt2HP5q5uH3P+CvYp8RATFPq+ULE7+Yq0VWZ739
1CfSMntJ8XF0XCDvtVGtDBdKPRutelmJltyR69JvibZ5xJ/Aigdmi9VmIJ7UONiK
OvyaV58eKGwE1wn7LKNcecekKRjJSlfk/RPgfiASoOdEHWVMvmLQTjFLtOHIE4Ce
51wrYGP6xgCcZLPdifPvQw4TGLgIviAdojvXW2dOu7dkIE6+++tSARGZ36E85mQ2
N7SG8mk+84B5206FK6dcr1lu/kEtferqTs0u0ztCb7C4E2JYGNVRcW+HMKQz5cnS
qdnrv6sK0UnkTqkkRcNsS9POHwdnHwQEMxhLUnA2sFCkoDtUZpjt49pjFAmQypt7
/gRKIoA8qVqSuOcIfWlcyW2lMJ+b2QtPQALi1631NbVOQWUapLsSOEHKAvOP5Vl+
DSMHZ4Ylb7we9eDQqaBiIK7LtUQWuzOw0Qw5ImjyrwbqUF3eoE6viIWquIWuT4a+
XFVaSPiT6KeLAZlTvMhNSjh9iS8BIBPzcCn2cH3zbzNwCnMAFKh2gS/yaKlUlUhu
haBORXRf+5KKiGArl/QlPhxoLzeYvZoy26+/DY5pMzjvIGHPq9rASm5gxkL/nKst
2d3AQkKU+JR2kbpGLt8rjhBMtw7LweNj+vSajStpxwnKdtCyN00Q8sTqX8pXJWcd
Z1630icdtqLiJTXgK1BWvOF/kC92ivAYZEMJXc566YGlysZRlCSKpI36/wCY+8vM
gdvGh/AUDGWzCDHb4vswp45+vzHGyl0OE3/LIbWCvfZFFQXmmN0iXbcmL1OCYFuN
+cdBrGNQD643dlqoDYjJz0of5R0+r3CP8h5pkyGV2iJoSy41bj+r5WG6cBnHRW6m
PeCp2U//UM80+5PyLBU3cxekSzBLggnweNRpAN7YB5pUyXtYxU9q0f4lGaIsKRx4
djJIxI7vkRcsGuabQA1ay9EsHvo3w1FCmuhxcJ9eJN+qlvmuasJ79K2ekzTuDeaf
Z9pHnzbh0w+EiZqPSaMn5NLCAEGhqsWj0IWIgX5N7IZGezxs652u8dXHXw8/fq52
QNhrf0Og3CMmubg7FWLottqUHymYpCnUOHiVbC9111Soy+bjdzn6Kd2t1Wa+dXK6
QauNunP5JOfbKNXSr//bzixpxEpZZKQ0NmlCaawo7Og40iNe3/8V2hl/KQulsFnU
R+EVulJ5n4vVfMqkYBfbwzHpey0Y0ha2tUl5co2c/bsVBB41ZZVnjnT9o6ktrvsK
ZH1gUuCOntmR/J7I7TAjOiW0gjDuB9HQ7yr3zXfRWcmooa0UjCG60YPrQ0/q0Klq
Drz5AhD6OsNf6UmE9WC+v0ELagZF6jVRM/8L9Rb8XOU/rK8THdfnidcbV3PJGG4o
3hEoUXxAvEbIMWoNB/idiSGs5jXRG/PGWthgXUfb8i7QAPu3rNG9NE8csFtTsJO7
Qp/Q/FWCJWspsro+xu5NIwc7MaI3A2aZ0ZxRrlXl6/tJc7k/PFinqi3Tj0M7vi2t
1U5pgz9DLnRjiWJFvZCpdIJLs6YQe46LEqVFoLHI1JvTo6XV1MPWts/LW4US0BJb
eTr9KA1IzoHK12Go6Ma51vwdSpgLbCqXlp1hVYOPt2FxFt9vqQ0J2IvvZ4qT46Xc
ld6yCnRV+EpXWfp//N8J2jWKCUr6bXkxJVlMXHjzqjwPX6/NjpeOYkIR54bdbw7j
4eeGFLy1m+oIkMOel/aopicpR5VMWHTiuZUYf59RCp4fKtzlphBC9yTw7LfjH/3B
M1yJu+pyldtzhl0xfZNPYDN8ETZLfMT62erkyxzErSZudshTP6IeehdrhzymfxNY
wIZt9QLY2LDMHL9OhZuXwWArin/MUFVIr8JN4KhfbcrgAwVHXa7SNOIOcxu+XvnB
yjATZO3A/4LV4thauMUm//eBsdOFWQgIbcQt4dFrBm7khnzKtVd+tSbOP8bUw459
CsxNWFgECUO9xu1Antn+mT+TwHPZG3VpXH5/YjG4Xe720gtXizaFw5dX5YhAQ6cb
2575ni31hg4sCV7HXR+9GFPg+giKiJaEbWMLkAxKO12QVM34rzdkDUWpDQJUZ2Ee
FqaspsYEcv0k2oY/cwLSCpCjrHkStYyBL26mgyBtv60l7Sb6zS5ro28g//BupZ61
XT8cwnE6TN56YTfkSzOvaOakF3yBEmXwWCgzEJU9GJdQmfQWfDwlX4yng3vdDJue
hOXSnVK6CWQl7Qp3ZJhKokGl8aTMhgT5nO0qtSwjyOpSqw/ydtwjWHNGyu/U5EU9
eF+9lP/7EgagVApVYyI2dauaXjURnUIbe3Pqs0GlksZJ4FiaCx7fnZZu9qDlk68K
bkydTu2NjroP+ZgXenX18w0kFi2GrEObr3NQqEXb8AvkWYCfOHu79aGFB4DkzK97
QGTQ+sBp3Asx+jWZZ1h4Fb9DdLozsjmNcIa0sx/K9AFyBLCacsZWUNXqLpJSc3e7
5SY4ssj4zFi+Hv5XjSsxg5CLLRRexOlGsgjIMsjAOXn4LliyLC6quO20wB/RmxP2
QjYxYSf9DUzWrvZWzxKMvqlcZu2ioKUAz/5XO6BtebtYv8hdum+8hQ3a1GV58N8s
o43jxISDjsJpxFutRvS5NIjuLVuCxxXHac46qcJgblGqJeiuDduzonm+uL358TxM
5ribWFFXuFkqLsTGTkvg4ckLsA1T+dcvonYms46KxYg2toKlFmUFl1RkuXEyGVVA
HVXEloySWzkR2Im02HinZeQ/o4RmQyYljFHsu9NIug7ybHnRVbiHvVtTN5TO3ujp
ToBfPti2jUQ3LE4IvGtj0+zFfxZR6HgWFSLc/nwFUXCGIMz1mVzgA1+m4YiRVvwf
JeLaflEW5ozRBAAo0uD00A6tF6Sk32zIIVIxWcByEp+pM3ouq9GWlXxRb3yMHOiK
Z1OOseEyU6I2ck9GVQjGKpDzFrMHG04OvGgpV1nZw+9EsVCv0n9Dl60uvSelFbVV
JcoJ9qaIwepJM0QSBqVawohdaK4b7uwjKN0NB23ZWkl535lrd/jKiTVVwPfGxiUY
6q1MOk/TV+u0j6tHbDZ0bTCT0qYupOUyofkFQrowgWvw9KdWt8LLVZQqnTUr71dg
52pdcnIf0NNU7G9CMgF1DEqyxxXcbiIWbIxthZmmNEWX9+gwFuS1KP/jgxSX9jmC
iHjPPNFZ33xCkFCDJAI7BaesV3zTm+GoL0s3jwb+mUGtcMTroIbIZYNZcDPIt6uj
CVacJq8LMZMWRzwiQ7Aeq5Cer9nMhG/K23Y3q96ZlfbIK6gmD1E+TqISHRbk0E35
67vIOSAn/fCH1XVQXklUmxhl1jmhga8xx7XG4oKsscE2jp9Lv0MgAPmGtWeN0vDr
zYLG0/1VOh2zpC7bhANVTPkIQPnBrpgZr8jmIaIQsTzx21TyjbOttNNyKSt5Q477
57z5sj+eL5OrKF2FXDdEdCjWChwK+Gt5t1FrtFar4KzlAE2b6dHz07h1LtB2Z11c
wAUH0J3ne/qBm9xuSlSEqxyPunu2kzsDvZoiUHy2GCTeCS9//lcVodBqoYJehod7
FZHhpNuMYU8Z/BP2b+fx9V5zKbQVjxjZLE9seWD9G1N1dCFSWcZa+8c5ffqA2jHd
tbR5oaQeJi4UhfVSdUjnF6lW1PlHk5pMVXCIYuna5OJ0txC7GXQeKZ1HBkjr+6tK
7RMkxIfJ9sew5GVMjWpdk3uVOy0QyxdJfC7+9DvV4BTI+jx/MU5ZNqET9gdQSjAV
/Y29y9YZ7kkjVsWNeeT1qO0XE+h0DbQItupmPnYDoLEbTqIc+slz6kRV2OM1h8IP
JY1HyBdfJ0A7x0TK114+xZa86STbwdRjWWkEQLE0S4jFvdiPrLnb2GntSapFzXGN
hlDNh5wK2ADPwwV5HgZS8PqK2B2UPuM2ZwbHPKHQkF3NGoiPDr/VRThrSR8/OquQ
I2eXESTuCSfI3eKW/W9vEzR5R+jkxuw6JOJSNOKFRjNzug/HmBkf+xiyTa9faNei
pLT1h6bJ6nag3VZa2YGVQj4MgwgPTBcjsVHDIVR/BpWHeeFyGFZSx6R+aT7Pno3/
ntwPDWUniGYcjjOGTeB3tcVbuPtYeHnSDqSTAR3EgXfOo+sJfgG7WI5J9kDhahfn
1PVh22WRhcM25xfJ9kpw+zAKdATsMxYZFd0atRM5YAnOLVVTR76EiSjT5m/uI5wp
IIwDTAAV3wvW3VoSll2vKu4qjjIOmXLo1OFVUXs86nFPC4+qUuSHYLagKFZvMier
Ol8/8jUpPBwQziVApTreSmMR7mfbKnwi9lqRmOdvqbgNHUza8/3HAp4Dy42eYpUO
Ybi8IBvgAn+9HXwJD+ciQppXTKknuZeKVsRvUPC/o6kMIlX6u3UDJ46r/TY6qsGH
7FUxDbwVNATFDVsD4VAa83vxm1smzNp0dKIi/yI4akBAL7n+61fY3MYwAs2Nn/7x
zCJvTSoGNcmKdsLF1HGRt3nlf1/7remSoqaqedT9xVNFj7vJ9zCb5gWP6sjaeufD
VLU3gJv8pZZ4HqshkOP4muLzhTVmOeGYzsNh5kBF0tUVR7zPHpSNwn3OtnFYi3k5
I+G33jweHF8xsOrAmanxbvhe7MtLhm54UoiEr8zGKqpqGVFCCPhGfoMPD/loWS9/
8fYwvIro1Utwgz/T6Gnopx9mhu7A2aMOD+f8Hb+07fQhb0VUkIrzO6eSqWcPNy7i
9ZahLsW/uoQ+wX1PSA4aD+UtoirpwyDCVTnNJYLRumSd2JBmWo+VLkY0GBzDB7T+
xNmjG8SLZ3NI7qhVZYOIgKEY9nEKYbi0QZXlr0VpxU6NxnItObNeFRSBbAY6n4zw
sez4zm6wMOO45s5FeaTbaUdS5h2rlS3mn/s+O3om5AQnD6JVsmmx1EXr44aYLOfT
WUI7bFxWJkET4UihqrxqCyI4YikJWl7PVKnFQhRlTZHN4ORIxXO2oZyBBAvyzcxj
GWxHRGxqq43RC3tzI16y8bKAv8RbzWvTl0ni1SyGGfBO2eHOlQUZMBII5KwULyQ/
e4fK5rIL6T+IbaPenEot2Ywh6SKyYqEwqka905DYehfsmfVqHUPnJZkIT0e/BjHx
qCZ8pR+WAyOhfYE4ye8e+4V0ZIW8toms0qcEBufdHW+roIKZTmDsaCsFk0G5hs6Y
JBVBRzUJfaExmQxZbKkyxuNsqn/mLHkiaBAiCgZiUQ4a5HYZrE8IvJZkdb2gsKLj
VnM9C/ob0aSK5aYOT7GubsYOCiM/pifndyy07TUw2e0Kowj9tYWG0QoT1C0SfhKM
aw5D1FxMwhPfJDLAokiJd6df0drdjCRKL7tpLN5qKJqtsFlwfXrJ2xuFlgu2gX++
94DqDwFcL7iJ+5m8pB8rM09P7NG7TXnuDr3AN2HcGrfim21WfxaZLe2qVHKcF0M2
hTKkxMUZ4HLNYzhjeciK40Y8fLmcVlhJqSmycbteUPgs6rNFOr15bSnd8um+MtV7
q2wxo1iZAEPlj2zYpf7BCaCB9Why/9dGcQrzwu9Kq4HvhwELsjJDBBA9kZvJIy4S
T232fHKKUXRAEHc6bvap4N1X97z7/1KprDZDSNNhzBW+DWainZdy7hOwsQEJaETh
7Tru85fEBxrDE6bTfrzo830751tY7Ibn5SqbitFz+SP6Pej0Zk5Wkm3KNcJOOKZr
YFeUl+tmwqdnGv7Wg3eLSx7woF4Dotz55tJ2NBaI+l8611WFuYeeI1akjMtfSPNh
BCg6jGfVtGY3mXXQfSo1XIg04rdAV20taGEVVVu421ky/v3vnwpLuCmmwVdZZuWz
xeeJ1n47PekOMM4iHYZNit1XPTRkos4KCRYjJAknJSrspNcrjYWXIoQYsrVGbtCg
R5bsNOAdsTQlsFD6DJULLbLXuxFy0U3TDPxtKw5sEVmX65gG6/mO4irhvAdpdVle
giUrEEaYOOSfNyTjJdOQd8X6qYZYrFsUCbeNGvt715aU5SPLlIJ4tnZBoS2bRhiF
Rup12hnINx80SHRv0gY01g37vOtipOTwuntGktwz1b+K5fQZ/UQSDd7OYZQFZOBX
SC0dyX6UYSkogQV+1lYf0DagyN1oiO7QUFeDXRJfoLzwQRNBEcibe7bDr0hJGpcE
LE57uHNyHpkynHr7rdqErOBAYTiEA8qGqtMHJIHf/gbs7/P35/urut6ndgR9vs9x
Uk+V+1bbb+CtYy0p78IJ3At1hF6iiFlvcd7B1WCQKXt/ZfsjHJobBBimfMRapsi9
Sgs4wZ+BmEfg13L87f4U1+7GG/y3GmNtBsd1ganAkGhdUTCDxKQaatXmHJxIq4mo
SqJEHHA9NPoDSh3oXOKOfNndnHA935rArIlWXyRr+cqWQrcjSOvqSi/oLUWHM/8c
zRUXdsJRNWkIvIr4ofc6Stpav6FvDHG1JBYPqd8Z0eVT5W2BWdUz8qTgBZQIPLOE
P72jIz7jFrYHTkWOVM0FFAm2upcCtadIUb70niiKDw/Ydpi0RV7U2EzdG0bcTCfS
HG7Q5M+3D6IDZin9M2e9E59JyhgrWFC/h8PuNqxOzeDU3z0Zzg7uOGEd92UeU+kA
4SDHe8iDKH93UfW//bNKwD08qdiH9f0UBNRfW1tlnU7ckzVtGNsUEyM39sVBQGtp
qSQubZlT1W9c5EvcAGLj3g+pwwkxJivFb5LXIeiqvOBX5QxE76g0m7jXxEFxPa/S
dKU3qKEVn4zB4JJvgnAa9pUEJ9XTS/H2OGc0cHUD0EUXnRctmt0I9aaK4DY1VpeC
V+HAEDABxSVtYAbEsn39/Hylorc0WXJ8hGbHzb0doReU02O2jHSLDv7/besoxtgt
sH8yUZ+IZNKQCxCpOG8IIzEXCEZ6kRvG4b6sWc611jw59FAwwY/mdT2QFw9/JSCB
YcWhmXJw9qfucDcj7OQbjBBcowxAg4QkRb/mKD/x7IAKqDAP2UnEW4gTaJPa25Ww
pR7iwJcCASLw2n4XAM54mMuWNuqQ6Vknta/W8BFK7RkxjCljD9UQg6I0EFmhWrD8
Upf59MS0By8iXkJrgw+cnzDrNnxzlLV1NP6aIEjUAOI/DnZ32LRAaMpcoMz+44ua
eFXMuvd6P5sUL4vFx4D28y8GiHugW2dvJiezQ1F1FfbA6GhDKar3Q3/qQblrc8Ad
U7HWT8eCleszx05gqhXces6bGcKg5smwHTzSHqTStS1erZKiQN7PLkf5tHv6LbUp
ytYOhzKa41yily7lfAEHSAmZLmWmxQRWeYB0a/eRqjAj+iIDSbSly0CxHfOUS7Qc
KNpLEv8ntqK68Ng5kdxjBwzMQn1VfhdREvSIa1y7U64i5jpgPppkS0LPbUSWa0FC
yXCOML8jpqbN+MJnLvgNebSK23PghYQ0H76KL1B+nwIdP6nBx1m3gmHikAlPr56H
j3TA4coAsXO3X/Av8C0e/Kb5BV3a1FDwAVaXLVdThN8zwpvFGgSeAf7wGPw148DW
AuPlfyK9cBxj/wdEp/RJg+5PI2LfZ+NYfLIKVMwY6OA5zYSZgMtGiGdI7n5yCiVA
ZhVkaJ4hdmW5fTuX/jwaVEHazQFortwdU/4ipe895NSeTAXJjRupLeAZjCN2UoF3
VQVqEaAIxsJpE0g/8qkIDQ9ArusHDmtFdsyuP5DD0hIwtCcGJGMgSTYfhxNg5rA1
D4OmCD8muoojE3QSouSbCpGET6MU7UjGc0ZjqJn7WZ9m0t+sM7lAFZSPa2p0Fh1f
nl8Wpj6b/FtdJQKGYTMQgAPt61+ZfOGTjfYfKSmrMfOAsZ0ffPUOvv1JowMzr4Bf
XRe8JR3aLiwCJe03vu7wVqzhdJ6s3CzPs+Lwc/M4QmNanNc2vVuX+8LbnxtafnqD
IZrUbI6K+Wcc/tusUeVzAdFiKGLLJIE5dosFFOqxS7VGLlCQQfpIZ5f/nv2gwjns
YYMpm3eDO4lPr4fgUknjRPv/5wmlRVvAP0ckZlCuWZVmdog4foCOKDKg/oN4aC0l
+heAK/nC/m9pu0XdvKnEbNoFUv6kV3x0luaPZ/hHATEf6UWl6FX9wfL3tlYq65Ix
SkeXciuPLL7t4vcArrLKiUdwFJkftiAzvRHt+U5KlolRnEQRy+s1koVVbUIKEdVA
gXRQBpi1r9aXsRtGd03kfgAOgICEAOYzI5JfltR9+i3kXxS6bq6BlnXn8mtGQPeM
VzqNZdFsoSqbax2ZRxukycGDQer/kztL0IonkuT0I1LiR+ht6Vsg1G3Z7++eMav6
mSageXrrb03X+mz72zN+eX9G51/09UTMjG2dcbc0tcZR6X+2zzWzEByGIqzWlR2S
J6woWV7MkGUSPXty7tMlYUmXFN45Mn4OfcWkMRKuty2S7Kbz7S01IzFUQp/xrJon
2r4arBdzSz+7iU+UbEanJ2Cdsn+/8fdUY6jYwMtLZxnMu7v+OkjiUXu8bURjCBIa
jZ+oDHblULooyGI9AXZt6cQklXOA6DxGfJKF8a1WRURvmEWUn9EbQIny00KpE7Q/
Y9leQy1Dk9gUa1HrV8q6TMuAWEhWSHMaGdFADpqHTewTvWqfhwcXreoO3/EJIBED
zCzBnh1W1WJk5Soz0fMBJlPFE/4ERaxL4LlFFZSpQPrLTiXYlDpz4jeWQ7h3CiCi
dBGOVyZTSNIb2Rc0QAk3F8erqR0Ubpnb8aGlQBUXSfVxmhocRrg3gpyG6IYDr8/Y
iJ2dExErwiXZGzh3GtzYhidAToywpDieSyZJTF4bJx4dWqkSsz/oqtEeZEG7QeaE
4bCNG8UKBVfeXLipIcnV0TPKh/qY4781T9QwynbF1ria/ETJXKsL1aj12f6HXNDq
nrSFrvnpqrDU6ZCK6UWVK9ELiSG3spZPL3G3Zs2D2954sh8cG5UyjyyDuPVyPr1Q
B2CAljP3s4geQAMbMI1/NUIPMBtkGfxUGd5xwBApiH8Ku/Y5SxklvpzjHeci0MyP
o1bE22xq8e3knExNBtp1d9iRH+lEP0ecPsfBOC5VihNpidNgk5v+weeG86dWSjjq
bADcj8vC489H+ckC1gVOHXh4L2BpharMEJIWdxkdCUhSWQsSi8EUEEecddyV1zBs
eufcVLLtF21ECW76/hySOjkIKv6QUGLuNVsx1AmT4hbjA5VN7cHeTmknn1kWj4Nq
k81siooihic4i1rI/W65N4ibnfSttkhvtoAfWzyIEx0NIZp7dajYuE7PBBWBmUUf
uR+UL8BG9u+FZz00EuoRC9D5WzSy5QoXrH+zIfLyqOckfDx+8skf0MQeFbAI8QJU
bqDoA1At9o/aIFlaVToElTgOCwuVC6Z6Tri74LW87rBGt/tGinDRG49OgUGGFPSd
9rMpbY4UOxmpoI3R2iT3aeqj2ZG3Lh8wqEHETd07jNAa+gDrvaz53U4fHt+28peV
wj1FO1uOpjC0BRPCpoJH8dPNFP3BXBZMEcIRyFA/D87ftEw80QG1zfzM8DdRBBw1
yjc5sA18qa7PmsqeLonfKFnhmj3AG5arJGCOAm+KIn6MWkFe+S4+sKDL4nQvBeS3
8oA3Y2AGLWrIOjfXzAbIqrJK395mzxCrUR4VjY1IzbKAe0gEMYfGgpHh00CnB8n0
8tK2Vh7l8S+rfT/Fke2Dtsk/wbftsjIgVPMbinbWrB3lY+Vdeq5N0peQK6IEfdIL
wVG696NrMhuojEhx/LcWbXRW/r/AT7Yk/tZDU+8K9KE5mzvWWY87IUM0PYfr9Z7D
ZfuRqZZUUJaJ18+Q4eOKksi2o1hIXmr0RHLZBs6/cCtnAnJPpBxBED7PK+C5J9Cr
3Gi15M5vombyFsx7OITPC5jaCLwwHZ8YnP0ZUrgBvXgCPNaKJKF4vfY15mmaWlGQ
Z18RQaEJfWPZS/66xDhFa9UKrnHXfExvvwrCQz2JE5r74vZ3xMWFMAUEnKkMc/bH
AIqQlYI0jCFGdWcZE1V4v85ZewYwO0HdT/Q12k5SFW6ZlYmCMouVHnOOFM+/N1v5
UIuIxLxTa/9FABaq99ZSEuB6TJ8oq+/qapGR5YP8825brFwkNccUFQVvuStArlXu
LMRigqsdq6ebxMew7RDZomb3Cfsh2Jg/B3XxwxMushe4mhbPI8rBLJCeSTIIUs48
8UKvMZR2yZ36GEuFWQE/JgzuMPbi0yTsJSKlBonG2a/2iazxfCqd90LH7NnMEUi4
5S1h73vMqzCUXgZBpnFrxRKvA1LG4tOATuc52p/ZpjDIuO1keyTzXVAL9xbqRB2E
GM4mGrcWYq7wC5Wlbz0qT8i6zgdWjBkpnhoObOha/5xuKkd+TU2Tfdp0KcuAbWIc
Uj+VHhcttVDnvfh/7MO4q2yq/iEb+txEm6bx9S0E4PrSxOkBveXKtn/ZQhC3xQeQ
Le1iJyHCB0q0WR+dPUsAEgRPBmhTkFE56/KNtaZFSo+HOT0Do61gtQAF1sJbKOtZ
vNouORAGs3o0+DME++wUK/R6ISJEarebQ9dblbs6bvXc7catxOk6KfUDs4OFbGpK
d/xtUV0OTsS/lFXnq6iTtYENbKkp+ScBI6Tnk3/BtOr/ugxo+OCot6D0uQweiED/
eX6XF7tp+3GDUpeSsmACzqE2CEm2CYPPnEMOTgXi37Vjc3jv56MOOa1kE4ptz+MA
tcLFP3KMRq7EKDCeaW3U2FlmOm5OP48aD3NDJA0fD1fLHHKGfCrF01dMb5N5lAU5
/MBZZOtlPy5LAPTW3WuZV+qoYehAOOf0Of6OmfegTmxyGgPoi+Udzffp6UHWOgrZ
MpoJmHpR5poYnjyJ7GVCynw5KrpRiWzJ1D9FxR27d4M9INMYXPOw9Eaa0BYwlWvB
e9z2IqU0/pbtI7zyDjbVDWSRH9YlCA85hNcfsf5VDvTeTll8ShVxwZ6A5H3BxfI9
m/5q+YtZaXq4+b5qf8lnXOqK5YhE/MnC2Ws5UqnBOHwWO52Q9eruk++n7zZ2iHBx
3MYp/EEJjuIrrnsk8YQ/66g3BeuiUmXcMRZBhifhaEN5j8kifNdq3edzU/K4vcUk
CapzT2maZnUhFSSSngRnorVMxvLJi71EQ9i/9HITIUcvGVGkB+AVOKafds76c7oj
zq+2f0QADAKmUgtnYEtkt3OdofzGHROvjsDVzYl8Felyvo9w7qsW3ifzFj/mLz+B
NUcgZZQ5P/7w3zP9ttdDhz6up2EgOfIpYB4RP3b3WB1VWpbuNeozr+U4bGngjMi2
4xVCujEWM7BM4OUVhehQtgNJJ3mQn8t6YY5ZtZTFrUZeEP1TNjYaG2bM4Bdo5/Xk
ROQSUIzT4aevK2fO/Jd/8bdOZ9FhhMoRclAvBnuhYgdQWfdbNkywiCknEX8S70Zi
II8iTUmNMYwjL0qOQ1V2p1xFyZi5HtLEAQ5oSQLVfEGjGCqykuuRJKZw2tS0SlKI
6Gu84mWCTqJkindlwc+VbQuIhgmGjOEccW+/KCkZqd8Q9Wxjxn3iEJbdceMs6FkO
kihag5ag4BCEuZhgN6Yg/TbgrYr/Zw7RKp0zMAC2+Xrqbh3wk68DTIVK4jM1Z2pG
8cTKvPrQ9bY1ZVKekfW1Q0uudhwFXB77Ng7P63pF2XWw1TCV/OvXb7+iMYauAMzI
co2w6pRn2Uu5d9lR+5ZqWUkCKFVJtFKivZt9nwEEdwSSX/XD38dko60dNke9I92J
nPWOAqCawkyw9vHnX5hLINj7fH5E67wkpbpBHJK67yNaCXmK0ujaPUt1UJKtRXr0
GPzjj5NuW0df2i35JIS/xrz2gcAQSSHMBvwNFwqBhNIHDFxFt/106YembUrz6pqp
BcOAhLBYvNUW9pROMR79Je7R4EnvtrsHxHq1w6M3a1+ChEvgZyHhNBMp7TQKkuFH
o5vZcL2gRsJMBR/eFxRbIZu3NYxBb+wC9xKtqidK0gTwnmPhK1hw30bGn1ex2yLO
gvwrMJDyero4Rgye2q/KVF2XVX/zrLoAF9lXgmJwKhAJl/wgi5h6pxAUM8KtL61M
MUICAshfo37C7nOoPup/FoZ64n6H7DpXJ3tWeYa1O8EDqixqc7wEPB2W9hYRg+7h
4eDsVSljKIBg4jEiqwhwT43bg8dO/OeH/cy7VuSSx8IVP5c5J/uSr1554vYCBtC0
ElV65zqfQaQLX+AbabJgXzHQONKAHTbZOel9Rvo+/lKoDcuqXWkMOa77m/kSmMLZ
xu+lDgqDaVnQgEnmIYq9XEho4NBZSfH/3zarhE4Ro+MXn+kWQ7JBeUh+y9QNScWJ
MdQ02jfk6og5qfJssung3UZjrznsdKFlTJeE7A/9jiDQGy7RKoPJ3PzpTXP4VNYd
o9x71o6j57ypVk3RgMk3AT1EhNdlSAE4EORcAWQVRsUA5BMyKmWgTMNpBB8dsePL
LCYtOt1rS0lURodbpqGtHtoRCRTUtXHtXsm6D2qCAQbOfGElUZam73GkR1PFWIDb
h1JAZ7sZiTzfeKVUShnuVe8gT6/W8OsMkwFR3gPXqtgdP2Mya1SN/eN3NR95NwdN
i3AIUYjyfWiPSBJw1J/FB1iZUpks9cG+5+/9Cu+mV9+nb2mHWOtAKPVWWjciovbQ
XI2n1DQqo5Vqe+Dr60oekNeTTjpE3M8OOjEBrqrpcf8XevVQ7QeipWGjrOHfsFO5
tIm4hdNijzDaVybtu5RSYTFANpAjdtu6z1NJeC2CZsLiLgWLp6HF7rdMqhVQdptg
da7oyXdLm0vQWVzI4he5d/crnM8ojhP7mjuoaIoHG4QFDmD54SqZjpv1gixKQnKm
61zqcOD3joYd/m3ftkHjGzdcGcT/juNQCpEARSqipCVMNMYjViHylJosRz3WIlhK
hMtkWkaIMCpUSsrMbzI/LnQLlMPL9QkMYYxfnLD3QcFYypEAPgzdANv+3zgzgSL1
+pBrrp1yG57EerzMoIBbCmscaiauTaxk2/WNbOqNb403z3XZNG5LPSixYW7zaf0C
ZslaPjP7B5Mzy2feirAQnoMXcGJo4r3cai/12ok+T61/4ETa4dP9Wb0gmKTe2kU8
6oV8GDyac6u3ylLYII5giY/NmAVS8I8XqYeoIdTlUu1yn7ERteo7NpyJozHo5iD8
s3Ty/GydUUPWeut5xTDCIFkC6IeDGxWm2FBD8lTc41dWW9qBYdpXl3RMp/qJjScL
7cg+aOtuLGiW2GYpgly7nkWjcm5OEeOf/YMVbrO8ndnM4b22mDl+b2IM3deQWSIz
zjQNuFWLpvLNnMbb7IuLsrzydJAgjYTC0+XxO4kC71LqvVgBjueALbptipb4cHeM
IKqFs0Lqa4ct9rPnY7NDzWSH7WaNABeAkM61Djv2lZWpsNj3h4sf/CmV6dvcd2wF
DbrMA/JVphTJCXtjD8n0h00fln/lopd9Y10z9xwy0q1CDzAozTLJiTarBHsuxZyT
F1pYz7xYgPz25iZLhjme4VlReVUJ19n/SRqMuZRApkQ8n5TAQFev69wKPheOFZ/S
gXRl7WVwdoJnfp5/hA2QTDTa5CDnfki0ffh2qJRo5wHJuUYI5KG3jtXlQxzWVIMv
koJt+EQi3hnM5laUPVmuEtUkd8toqTvDdj47TG3yTvHgnxVnNMflsqn+a4cVd0qZ
xZOqWGncqsR6y5Ksh+j3RZ5Ohuwi1Lv8pWdeMpPcXT+WrTa1M90c14dF1IThDzJA
RRtA2mef+8T9OgISCEKEhXW5XabGeDxxvJcjPshLrS5u/P11BWpzxWigqVV9bRRs
CcMOEeTY5DJ+gFviYDfcP8BZBWCty88/YqgqRjsV2fpshPkkVvc2tNRCRvEhYWAt
hyMmu8t3jl1JaspL15pgC39Bu5y1b+bEACj80WdCvJawLzQNDTJgQeJdXX0ermdE
kmGaT0BUq/IzPon6Vney5bV62YQXhZUk/Iymok8v4RNxwchwdkSlP9WvWCL2rIpu
Zsn/Y4B8ClyMTeY45ID12bCneQMahLmYwoRVzymfHI5jUitss5QwVKiPxj2Mb4M3
4TyFCdbdyj1X2oJf3FSEfToDEzGZbC4ybOzj+h6eRJVPfcVj9VAjgNNg/U8Vv8Zo
pshPFzAMe3kciP2U9hdJ1Wm0RRlz8wsirRN8ZJphUMJZr4u5uF5OpZP7bhCwyHd3
GKvrhyVD4wZ860i98f/K9dAVw8/xtSCxE8uHgJd3gvXXTovFNQyKnuaUSJewnzgU
bdCLXr4sANjXF1CkD6aFALlknK5fFb6nmfAryZQhzcQjC8jbcnO02m8i5NEwM7md
oYQvi/bfrwHMK66kzo5AW3KHo4gLNB6oVWu75XYV/NRxp+XOA4q7oW3LsDavAry+
8uGsKH5+bMwpX08VPeQm7HmDC6b4r834yXZukGYuzBO3VeVAwyYE43guczgjRYMI
mh2huiP7JNovuadaefrwLZrKvzwexJbRr1YDv3ij2+iwZErfOJAW1tdmYcpeyZHJ
M0AGzDXuDm8gs/bha8Vz6KRkNqzVdXK1n8hDD8BnD9D96AO0bGwK4XdeIbbZEURO
kjxKiRbSihc8lzRXyLDM5qDPS8ofTCZ5nMlvZ3ZU8e0/300CBHlSk3GYykvSP4rL
frOSV0+cbNZpfvP2t7cgalXQwjuz0OBPAxxyULdlSX6aevTAQABEXM0BCKwGN1Z3
0h4soWuLXQmF6BOOomx3AFHKNOgnTUXWbonewNlRhGgKvgE9NXD/MLsbEtHuAXoU
KOGJ0FwET4SMMNr05o7+psP5yWEyh5MupqbrzkJHcY60vlpVQqSYQWWrxSj+xrIu
FB/wg3kh9dea90+deZFiKRBWVQVq27ep8LXhsKcU+v7WsYf5I+WAHj0jh+pDfW38
qalKKXCb0QI9ZeS6BwNrN1aj6syz/Q5MILL+THXe0Ap4l66+txVlK+OxthmfQJFz
DJFxeW9/ikCWNkQgFa17TvNXnb8fu/1/Rv4/PF4YWVfKzaBy4uwPLpYrithj0pG2
599tfOv+rX3fRuOsFs3yxMj7/8e4tGVpeKnSRHo82Qgxpx3T/IMP6xd51rZp3yRn
Ow2A5aJlCoCT6RQ3AXwEHtqB5LftTyf2IKZmnBvjSuBtydw0YVVahv/5jbeRchLp
JZZPZqlNj/KwfIrp1yT8agaDFLqMSIwC7dilvDXFTD82WTdEeUOwwYINdRj5PWsa
hMX4FR7eEYfwEBwtiGIsqlean5Iw49MrhC/jRdovKS77JHec5EDelPWyOHc162x8
BeRaieRwTHQErdGpIBAxv/I/tw1dkLJpvfbAppS7U7RUkYMPTF5NvIXEPxOuHdx4
LkC9LUHyqGHsyQEYci3x+Djz6EUhHtZOnw4vW4iMaUGKUIvzM8W4QQlhmylC4LAj
bKTHpnZsLCgwPRqKvmWkUlB9Kmw0Erwptwaxi+F3WbN62O4axW7UmojlYFwvRQYC
KwIZmpc70lP0VEiLS+YSz/PPg8AmfHkWPZyC8m+0N0cDHYhEY3N0rOxzRZ+xacML
dfagvFs40UHAZ6ICJMySWaFgqBtB6EE+j0u3nxm9V4i2di+Do/FO+YztdGI3SDgw
9xJs6HzbzXrcezvQlbT+Uyi/bNHoSS2LGxJnZNI0mFf6yMUomzZiHW2RmI9Ub4Ti
oP4l12/8q1NSwmgeF+qdLuR4iMStg1PCNACS/xre/E4Za9eNeMtH2DpyoF2Lk81Y
CUQNPAGO673MUfkI/rPRL9VPB1LE5y5BZMoDXPqsYqfWZ+ehv7OXbwR4kvHGW1Kj
y+2i6TACyUvGh1LXMU0rgQ+QPGU+CfBE+Bo/Epn6fsiiXD3cHq48hTr2Npnli6aS
Har0o89pn9GiXl9ndItf0AFxtbQfL2QcxYM4/45oNx7wHjVDVSBkWUJ5iWE+lt4O
k5G+23MQPaDnDP/Wh/uxZOxwJryDc+NXx/gO0tN9K6gsqBGzRTU56S9h5mMJyC2o
dyjgRyszvCnXd4wynea0SvQne6DEG4uEe7kfr8mbM4ysBo+OIyGOZVbHJdFNDr/y
3sx0Y2YsOIYGC668mTYTQVk0OUcmfoSfyLroj6kGQzZJXmEYNCdkhui2wYI7kKQT
mSWen+oPkjurVlTCjCfNK9aWC+WKh+NhEGJH4yYgoRutTbhpVOc8/t4jCYw08C75
Q1DyoHMArrDkgMnJOdLCb93xGxOStrP/xHCVJuBtyFiZFZarA4eT4kpRIcZvvYOl
tjlMSJPVgx3iA9J/HMy6M/Ni6uJ7PioH1RQQYx7taT5jvnq/PV1bs3IQ7Ywkh3aG
eMgCAxGdMvUkym6LCli+RTTo3kma5993/ddk/DEAizVx2BPWHz1hFKuvukbF2Ywh
2/2BAXIb0c8riaz2PXXt4kQKaO+z6sZ75wlO0oFJIxGiqa3u9Hi9vMCY3AAVvjwb
sK+kFTj0PFmIuN097LvWaL7KJWWHvSBY7nKMbBWvde/9TTaLowlCJpXdNltftAEy
wDNRl2doBqOQryQ8lRXOGQiISy0ha3F+QfsVCTqp7Iu2bpf+tN5vla0BVmK/88q6
39Lk7aTUHKxaPmi06vTbgg1GBNHCE6BzyeJ+8ZC9o5zkTxqpxu+Z7vqPIBcI5VwB
eqvq+2xzRNwmCd0KXFyUEOZhoF7f+GlUEy0lfoLrCKSKVLHEBR8n9Dmq6F34Xyzh
ZJoBuJc495ajNaihAj5DSASxkmUVNSCYYTR7KEEH4cINsYEIitZYxG9jayb0Df8u
E2d5wbz6aJvETXPpkxfI9dJu17x/xN+4nhzBA+bSzWg6oqubWzuO0Qh+BJTFXdaT
5AOTKUW3lTIt7lWCtREi+F+FAB3Wn4kP6caE3nOKCbO49YTG/fIAxH4GRxbwkWWB
R32OS52FZihORw24KTtbx5wUIKTm0oqxLvD0vT2hiL20OIKffGF3NG8Zfj7Ul8ut
+frRO55E01FnUowjnarbgQHJp5x4yNgun2aMglZVWKUMvDXNnobNJyvoP3O/DFe6
qR0FLFq9P5QTQPdpZswcrUJnldt38tboS0JKLw2leDWhAoThvJsDxI/Z4OFDrF+X
0osDIbJPcPjgFPNOUNFW80tnsZ1wG4lhkB7p4P26Egd06eGr9vOaHnk2mRihcVCV
ASoKl8KE2sXspZDrh5qPkbAFMMP5x5uiowuntCkS9BvKfl6sPcxIERBqaSRVhXxi
QB/Xkfq7D3Q3e1dIQbIOODauNhbI8LkSqoZhKovRtRW+BqpJdEn6n6fcBu9TU+RF
W+J7GHD8Rv7qPJTtMK9HXfUyrMVwZGqaqSw2tK+ui6Xs49hVXILXtpl7XCvd6Bk3
QBStT2X/ObmNwTdGGLN3Ecv/kR6ewGA0DAe3geYaKowFMEVohNjT37ZtG74cdhbo
H4f9iNPvAPwPBmEa1pnnfQB9GeINiPIr8s3RW4tIce/hf6w61459a20+uN9/wh4x
cnSAo0QWJNnNSWjk7LgMT/VdEJKxGopTD7jVGgVJfDNlmu3V/y2B2yC2mrVPUeu5
9EOHbWRMpb2F1+E8SQrqlOp4T4oOIjKOZjMD5ViM/iB4Plffpyz0h8CXHWTmCFZ4
teqm/LljkBHVJmfYUEDjBEQix1JxLIPpuATywzl7VZXNuQhCD+HFJP7LXZQoV0yw
v6zQvOYIWz32T4pR2MU/Vntx57IcFbVWaLsyBOVhzqZGXIq3cBTmFTNRgHU1BntP
bV0021dmvKrdq90SLZgcuqfGnX4/qepWiNodlQ5Pth9+i0Par/5PmtPEDKoT9XA6
YVrjOuECOR/xHuINwCNX1NoEiQ8l/GuHoLS23Upgok5sHRhV9d0vK30Lm222cz7h
uit0gjKlYI29EiExBHkO25v6BQZH5C92T/PwxBUHrjFDsvqiwTadXGFR21/IpEca
02qA4rySGl0OJZ1QZWtt4REdRHVrp/oQ9+MTOhiRolLwV5WpxsMaRkMCLOvaeA9G
17/UCNExnWzEXQmM/3P9fghqXPdtD1Qzo/YEMNC133j5+m376tIKZRqu8me0RMGb
yRTzToHEp0is+kcxIPN7Cq86j5jzks35aQVDgiqiFx3BFY7w3QyT8m4TAwQ873NO
JTgJfr1jd//agAKcvyTp7hu+rUYKhAzINvfR4KvnxjqZFZ+rwewdVMlRsCHLt7Vr
RSiuUMi7MIUQlqgFZR1tPcOHg26FoX3gNgGtqu1GfNjhzzyBV6gQyfsyTdrowvM2
U3oLu6WPvfICj6rswlj17PpgmlQrREzT5fDzrm0sIQZ4I+n2W4MO+swiPDzvllBP
yIj7C/O1lB3ReeUAty47JVmoFwsgszuMKN0ZbtVjf2e621o6iizMK/4zIu3t9OQf
RjvX1iRM4Sr1SQO5nOxCyOpcBwM6qh0atB317s1ziVj5LNdd8VsCo2D1HDYJznDO
4SndvfrzSmBoWlLtPFB1+iO8as/K4yaR+/6breCcSGT4FAdcXAfXY5rs1SDIuw1c
r6tmKVFtNyxikRCltiv3xbw+/70CdDjv9wbC0a91upb1WkvhNlo5pJjx8V3pbqiI
9CfYDvOT0pPPOOEcWx6tXnC2N82pv79a/G1v+8cyIq8aYqssUCC7yryTZtBxqXox
QORVUt90dvsuqEPZfdT5d/hJVSOTW5KFu71rKAIrEYy6epcaKnAcCTgTdIeXgSCI
fPU6bxjnOX0bG/dI9ZDO6JZLnTwyFZKuHPac6Ujo5EI0P/mHGcng18hj32b5c/EO
+FVtDLNEdX0kvA0bac/WU8+K9B3jpnD9m362uJ8oce26qrJSm7tw4rRwWQd4wk4D
a8v493M+T5S5SqW/6DXDAGj/G9FBjms5iZezgvjENYK1BzGe/nAtLPSeaMWKuMxJ
fV51qLy9fwrxPY82Ad4Z6a3xBKoJkW0Xs6gFf8s58WiY4HW5fVlGrOy0YQgOXFV8
qtCHD+YOIGXI3Js3n8MimlBivijRb+gnav74Q2I6eHel/r8k9FGGnXxu9xxq/gYr
niwNUVxogU4ANbo4TXuRoubDicOWLA5SaNXerO8YE2LyMTicu+p4KIpewmjUxygl
z/BvBq72Sa6LCl+Q5h3HN8LAM83yTkDpbHkB6nj5UJ7T8jHj8WDflUdQsbXhqsNK
gsnZw2AO30cDXBXNtpv1mxkcYzGHlAiWkHlnxU590mEZYRBp3RtSnMX/1D5/e1yp
VnArOK5hnf2Pt/Gmgk2IRmF4+QwHmQetxJTW+GP9x9+jQGZZI+jzJFNvax40g9QF
N6ga7N4tU9auH+WaBNSNGdRxtvJtQNxWfJxhTnQ8R0qqSsEn/vY0MnWvHjh1AAFS
YbJ3oaA4yXdzNztVD9NNdyP5zBQnz/OuDK7p4a3G+tZFUy0r81b5N/Ndj4fdIlWG
LXMq1Njf5kUpxLLGzjtTjIdUpXrAxCixJZAYzXStglnz5Q7BYV13s9wpeYbuxKar
Qko3IqAgvzKaEYj9oZWd9JQMffQo1MHHJyluo6Wd+fXiu8e8Ehobb2PNUVmV4Es4
Wn80osOFXCuHLFY6pu5UhSMVO1kBL1PTr1IA1APIAaMAcFJ8ncxrTR3OEmaYP3Qx
+GPpeJPEeJLUUQE7mCNV2IkYNM5n2JgHZZeJ+Lwxsta+3fKsYhxs35xPJUyhtqKz
wU7m3b+qt0fvNdgf6TCLfYemoqpSIgoxsbyCWz/erF8ovYxPUU6QUJbiYE3x6Nkw
4XaZXmbHJyZfuB588/5Ix64gF9dzLjU8F6EXRHOV/5b9BUOUxWEyR0XpJBqkfNpP
fODbp5kDLqA2jGiYVeT2RtvLfzylvzj60ll5IQiRcFuS4gvhjk1VvOD3cOhsoDuG
un8wTW7l+WDH9foDNWkBIxQ0u895IT+PxQCwnem6JxsMHWMXXaAkgU0Z/nAhaKT5
pXXDHzdgH2OoQ34moQs29Ef260CMyXnnECThPMBOzP3dtdSpR07Y6+7sw+nfuCwL
0dBwfCO0DA9Pw7Tt2gf1bfCWnSG1vs91qQEyAg9eGeVyz7LYxTuEWN1BcZp/VJ4W
y3TB08El+quKqy0uu330YHxTyUCA1aqjWL5kTqgU9xKnkl7VhVdO1X+DB1JFBAZB
PciYdB5NC+48lVQK8zDmtrVkDvWFx+N+6WBwjy08WGv1jtJv9Vk6rqne7C1PpFq+
l70G2ctKxhiSTgD4kyrefuQAO67Ksm8onfcq4d4+l/lSJzs32kVVPNRr/17heMnx
Gjncz2PB85UgC1kTeymFsVNlnwVi1AqoC9K4fOLIxYE9v62NJwxTdfX8r0VgDEYD
Rxe+x0ungyPBsjaPc94FWxIYj9rUwNeREBDwwY0W8voS8H5AbhdOA3ycEUXcZmWt
D48Ng/6JupSD5qOrLLS0f5LL2al1lU+b+MhimB+zwrzz8f9c71mItdhRIOhxZgfv
MBioTn/rW5n4gl1TrtybOZWraO7piOOQinZnvykbXmwJ5xhW0BZ0aCFkb4io/3g3
x8LIjZxtyzDBz3GqHr6g1LAr0GUJW4nzQ77U47VA2sneYneU8jyPRcqGpwLbFpSF
fWCHnwH3mLh4SdpLTgKrtCDg046AbvCPO/loR6ygRhOCpx36a4GPWJiE9xO6h57J
CnCeimU+TL5DSPaOOlj8tWgVALOrdKv+1YqBn1FuWg0Whax4CAQPtmS/dPyscgAn
JyQTfjZQpblJS+UhYgcUCyO/m7vrBQayHQWZrgV/BbtCJh/b2rpRoueDywMpxQLq
QQzr0uWyZWNARV9kpX3sWBG75mD3lyTTZdUntVV4MNTiPoh4A7aXBmb9jRCAroXc
r1UjyVWezT/Mpkr2ls11xlLt3lX3aDZiJI544gMSsudwiY1/qoiuJdeNkqUZh2Gl
SOfR2RlqeliMBiDYpulSAe0RbBod3Cf0+FzZoJM35NYZNLKAXXpplSzC/VPpTGj/
SFp+gyziudLymaeovwygOGdl780qhc1jTKvsoYkgS6w7qIbIdZAlszOwz22apaKm
bMXKJSRwf8B53Q8dM7HAccy5NHo98s/4E5UMlFMoYG/5TLBWTp7AboGnQ755LR6I
Adx+r0zwluOwVjzf3Jxhe+ZElN5le3mWETRn9N8gcFYY/rvRlhhQpW1nKQhYo8ep
zpLg+hiAddhQZTe0zWAnSfgdGZAhpufVEKapTfqKwd3Iu506YPtKbtUq/NCBbult
AnwpaI1lRnFqg3PdzPaDq+lv5R4DsQ6BAL9puDelombfG3pzEDR2/WK2Mkckr/0e
4g9jCmr9V2IKwn4Pk1HYblMbaSSLPcbVzLCrVPEhuHnIclgHAowFYVzraSOb0ZcG
J88wLXYaNFx7Kkf8GO4Rqojo4tPrtTIvID/o+wp3vn0WL3gKZNLPHRhYvF5XLsi4
9Nfk6FVUJabycKupHYOzFMlsGH7hcVHJgmfcUZE92g+kurryVLRLrQrEci68g1x/
dpVAHe+df/bIuqKY0RuKmhULubHj4S1srUqUouxPbu1wz2itI74PlDgDXrtgRoyc
Jz/Jkn8u/Ai5kOeLQd/2PniKXGxHXFwo6CDQYZvv8Pg55sLcZebNshNIVi6tdq0H
Kfb83sLBol6DG+ZCjK0l+3MLeOeLBxekTR4tz+M7aLwK+ay4Wm2YE/1+2Sot/OyG
nA3EB0yTjfYLA53+l7+lH6NX5wbqd5oXPDqW/Kcc+af3+AuF/10+XUhcdVCDeK6M
j6prG9roA9EeIWBejxNJJYul4V/ct6gghcrXX00iIx5U1COlROPMpsdGqaZ+xXdh
X+lPw3+hQiApyr5zvxThjKGN596HQ3QjIn6a4P5Z/fPQ7jroIGMG9Jij48hFLKld
yCXSzE6QVpGFus5M19vBPXyYsOdzlhRSImjTfL+06EeIqyjAR+1wb9RhBGDLYeiv
ApFQrzfM26YV3EBz9dEZzfWxstdJ37lsU4ipuY/1bWxNHCvZ1k8ktjY+wb+Ojnxt
hT2NCKvEeEBlUIMai+Aetpeg8nxCnFAROmZ1J16O9WxujHSVpSg1OJ5kYtJNftRU
shgEuqkvpYy+1ExL/9RXzZ4+XAvmBElyZPC77gfVe8sbXxgwa24asn7/MTNjIlhB
3gDsLKzMLZFbqDhARXIRV8OG0Zs14D/xWIzUxkO6/wJAZOSbZcGBfVInneGOGLOJ
Ui5W5MHAffFFx3b13qtVgQM8S+Ea8rcE/ZJYCd3vxCh/OMWIOLNtnQYK/ZpNvOyf
cBUDV7rBasPCgbU0dKSqjn/GfoH5kQNvRcxZ0nrd5jdXQBpQctNaz4x84YJqwgH/
WpUyxAv44f5n52nfkhIUwfl4hYb0U/ithQGbBLwc+KLEYxY863uqT3rwkYEp1ZkT
LmC5Au/EkA7MYKPY6S2/Dmzb/0PG3khLzm4gkfXtTVNTIyw3zBJUFUBc5PSybFgq
l4nQy6NcaEGZRIGLIJEYbmDk8x8IvNzB1h7/kygOZw/SDzjAzft7YjqzYxIG6xY1
4UreKUda+JWljljGVxQXpaL9veaij6JB1XJlGRO0+VwGIiZ1EhBDCjX0Xwa4kFUV
n82DjnS5FuhXMzLZ3Embq5K8D/03PLzLCj3BI8KGIR6DmGUDRflqk9WBy/8BGLUb
6oKSGR/jLZjnaffyPK0jLnO/w2O4yuLVOeWt1S0jC8h6sRXj602XbxyXxOnqPttk
9scSrJfFJMvdDpadUzhW2avnz9jg23KX91fzQAK4IMGwsn2OI37V8JJDRcmVimV2
bKe3gJoqeTvz9SEyXLvpjV6py/AVilIzxqXYQ4TgBCUGzr6WEFahHNpqbr91+dZA
JH64qOVzZEccd+Fsjb9kUR7qqio46g9Qqqif3PhoBvv6h4u2O8TyvzTJ8qf4d1X4
Db66fccsIqMttHUka+YcsCRZkjJQJ25YTU23B9IgEVuTJcFOhQyOxu4IULetDPq5
NDRTbokCygW/SA2vDI/ek4j6Uy4m4zEeCfjN90u0UIwFTqBgW1qx4lx9K50bFWlE
un/qQYxrc7ZbVUqiAl8NNtVEO/xIeI0uYWcYkBxHmwGHgnECVpOeQgGaIKkc2ZbN
iju/BIzp8UW4xgu2FJBvt4W2TA5J8LhgXRzb+DccxkzQY+SSM5iDLq9rfXcUjpbR
uq7jpFv0JiKz013WtKETb2VU1F6klLHzPhsKEbAsdNcknSsTB9B2vPsGAp9hVu0N
G5Zai/5Pbt5mjjdPcjsxi2+15Rjl0QnqdvGX4/AdjquQLSpMBBJ+hkTzRlVfM2qD
LGJGcugZQACQTT7F6IyAv8TFglZP9p1F4alZy5/jnGj47uXbfA4obdkF2SAGTb67
bITP3IKVYKTOGm0X4DY0Ohp5kUJWwNcp/a/F44V9szajBzgCVCiaVKXIhRWHKzSM
AgJgkBYlLvyPyau2IXY/R+yolUlFcS3eXKBgfN5q5+ZVAIESfN/XyTKC4PM1SzFV
h9AFjXO+SEZEoO2S95f7QHiebXxgRGe7370iXvcosRmkbk//1+dLDSHQHd/C/ba5
/i/W4vVtbE1J/pzKwhScpw4OpAbmF/cFulg0w3M7D8frVoHw6FjfaiD+Atc/7kUT
fzpxBTnQDFiyZ50XE9iLP9kjdK3s8lGosV8+Wn1OJEd7c5KUT27uxjDVY+bpMeA/
5Oc3mMLHp3trgufjxv6+hp3HP4brmrVz/sLG5lWaVOEk76wi3Yigb7nFvv/1T045
v5txyFyYssL8ThyNj1vpYQhDnyQv614HnUYNJgjvT27NOQkJuMxUAjTQR/1mu1M1
UVzx2NOQi/ThnhJl3c8rf/v3TBFJXcyDFVjohORX9Nc0ii2RLWNKYSHFWwqSLxq8
OKHmwgIwChtPYh+PdqmY6TMMkfCTjwaifzrKQxvCrFzv19w3EUpkiiG5ogfPXmPd
PzVXPzOnVPLk88ZcQ6+JXVUqiTb2FYhakiFO4ZtLX/YHqQ1xZDxzBAQJjMgHi6Jw
ez8s69F5FRBW+g+yeijz64sHDTZUfYnc/dLbjXsxoQXwnaODgiHNRJfdy19LewGh
M+9qVjZxPxL3V5Pd36haBA9QQWfhLCIpSi0V/DP6y8WI+EPX5CuIfTvpVKhSAiSy
n+dp6SHVOGUxbScAiid4SDwzoV/EOm+pjC1nzsHIWjrGDnLPNmWefJMRG1I13+7d
jBr/0sRjObfNMoZGLE02oTfJL8fyik9O0cS0QsZoB49XKtlvikX429/du3VmhIpT
dPi4lfTznlBwaqBBooZMZAwq2klOKr9QalnyokXc6UD4wBahUbX3TkYBCL+EVk5G
R4MlzxRxEOC4TBSTbqVWfNDn9G3NMkNin9nWFILdcQaMOMisPGYn+jhb0NKi+T/M
Q560xxggIVFXrdXPHWDBLRtzCeYGOQF1PKoyr5PKQOjR1go0hBe6uFCy1a6SumCk
lcdhf1dKA3WEyXcwnWozl/MsxOspf5MersHqN0VyjUuhf7f4tT10diTwp70Q/Dfl
EGXuu9E+a/2CPo4bsK1bQcxAKkIA3EmYUxY3dIof9ehM28n9QsmlwjFR3JHH/W/E
M83ktHP972NYi8nsG2Wf2iXTf+/hwtt6QtBYQpaFz4xN8lDWAfkvpfb30lbnDCLq
8BPW6g7py3l2vi+xkI6nQR9nNLvlWjaz8eeXPK9u9uVO/ZKQTgxmj8mXr0zV2mkO
BAJiogYRyTYRGmqxU0tHvYMxTyI3yUkTFcwLKlKkjORKD7/E/1gKiWOGiULwO2cG
DoJuMHkpj9McYRhyC40KEqUu9JcASzEPXKglKx3Xiln2FRZSJBtQXOycIEF1fFNB
WLmBH/l2fvRbkVL1Rha2lZdy8409/Wc2H1kMrShISh+qf4FS7dqya1iy/KReCx2T
fauWDBExIB4yZF+8lv9p3dV0IlNnFUlmERPf38USja4Ce1uxXwCoGBYR3oz1Xqqn
mpSpcMXUPZiHfqHjkp7bweZHzGQ78cbjVQf3MfLOQOjWz4geCcupsIRQSnzD0jK7
QQwZ/lHvVOjqLza2nF3x2Km0p9qE5aHb3P7KCwjcMtU09n2IjKLM9BR80lMX97sV
wZH4alDDyzgouoEx71JQar2fWb7bMtpnO64DaYQtzicOcC+VEMUVXccywwKzs2Xf
bpacZ02vcx8BdXZ0gr7lqWbpQdjVPT41OXOFyq92XhxVMJn7QxymC6TqbPvWhFLT
LVTYUrJzr8Z9MTFfUGNI6w4mVLxD9Bvv3GOwumlEf1gPiTtCjAdIhVS43lgYP8SR
kDvjzUKX+N++PMLNTJFn72bg7KIlTByd2s6arL7NLqfWB2HZf4QrhaMp+lVkOisa
2oTeALoFO86O6ZESRN6iXYB+nOyAZ4Sq+5D85XcJvcda5OFCO0rg17zbgfHMq4sL
pSUO0Q8j5wlIRWOaBuLvdwyItElhtI4tg5SnCxJuRY2pHiiGB0UxKXF8qnTh2QvZ
z/KePgYOU6bkXUwag4aFrSvKP6U2EkAzMJye9h0h878ODXUIU7r5Nm7lL56ajl4f
fna579vH0xDyr9GxPxWQtA3+o4CPuop9XLVf0Lj5pZdUC+y8oOMQtJCSA6TIfKDg
Oj3xMA57c3O8Ev7ahbN0tVs5a/khfEwSIPzFOM8Kwk26j639gKeYjdCst5dRymVp
nusQJP62D5HcZFX/bIzlUaR9yabT1xboh3qNfRGCTWQSXX9gw1oY+Z0pYkjPpqp7
1wEBTqWy6v8GuPyBzfoVHLMpv09ribtm6SPlmbRTgxTF68AFHQl8gyU8m3VaDdF1
mdzSTydl9dEglFoGP6sYmKL4Imu5Rk0hSjkzYA3RVbblgBJUwB7XYMhgz8VeQuy+
J3vIhOM4LyOT0UNiYNUS3XeY8zrRoNha8B5bUoW/UFEH/Z1J/eFC5boh4MRSZD1E
5N6hqxdQO5Uv4VDUhsn2mhzetFgdThwINYnaGV61+cAYiugFjdnBooC9I0ssZt+/
V+RqbsfzcrKcswdX72w8SU/p4AIteq2WZ5AMjelx6a14XCuPGcOULrRpBW7vw+r/
LkONOiD4BmB0R8PScGiQp2fONhCeMGBiq7RHwmdQFV/8BT2H/oTdzkQAvX8h3FAA
NrOAIODW3GNRu92lYejjOZ7Ayq6vzqH1q7mmORH87AK81P2EfjAtF5o+Lg2MmwrL
XzbIyWtbtNCHyeEQaBYAgGK+/mSuuODnrJOO+eO2i9KjsWQPPgrtnHFU7iBY1Wxz
BPQ0GB9pW/v4oqYDOS4UEubXlqkXtGc465GLWdFpD6xYNH2q9AGo5rt1Fcg4uk2T
kXW5uCriIRzI3cjjC5sYMnUmaOk+2eSd4hPGHE89mpxglVZSeqdvppQQt++Q67Rl
IMwHyK1UdP1P9UUsAVHFqQh2recazURDlzXXSIcX2aLC3k/+aptbuTVBtblLGKNN
ox3a4oFBks5BZoYiSHKo0LnvmMOmwK0CIuOh/flTNjaDHtTGGY3dT6A7Ce39V7og
F1jAuYKXLVWbiiKB2RzpPOdLEwMOvMXTY/ijQVexfJJbw4K2vXTsGYI2q2L9x4kJ
+roYY+FWPLOs05MQjPnjmE2ItlJXELXvwAfEgo4U6Vx50RkEC/CXS9++KmtDRwQz
SomLFZDkFkckK36jNHkSfuc8OmJ4HjXwJP0U2fDhLoVqVD2vhVqAGadYCQf7mGwS
h2757/pkbQw9MimiOWD+x4Bfyj9z+dlcIWjAURlp0vJ/jHmHUBcE+twP8N8+7F+3
l0FNXj/x5yQXAIcmzYETOHkSA6jaQ5amWzN2m0CGLKJZj8pJ8A3WpO899NolQ8ek
1FhgKv2uWtmhoNMGyJn3dtE7q/c9fnsEWxMrelm5MaY5ppX4lxGPcIrz5H66WHVq
QamwCJTFYAN6vck5Zns+K2CZv7pw7hWuXpQBPEbBOhCSIfm6bULV03mtFLAUtiDS
egPU1Mwup+pfF2beQ4cFpjYAtjqL6/Ih0jTXgk3gSU9yGrLa7Fys7r3k4MgL5upe
iyxjEgeCycUVRKtS7i9i2HlIzsA1E7/9u53g+st7YBBgoD2okAKUWcpqSkuI5s92
UqUSmVCeIdEhpKtTAkuudJ8CKABAGK0KmpVL3b7s2y+r3ZCV0GLq6cjpk/HRVFi7
URNqEsFRphiOzxyHBUF9dPgI9SD5QM6Ham+EdhGVAuqrqB/5W/+mz5ELE+2O2XXV
DaiyQT9JsekoNb4/eICL7Zia3kXoHfGmqxojwEq+tZAs/KDJ3w+7OFRdrLL3kYCT
OpSKGkK916HvFam3j8rP7Tan3YJOJsGx1HKttkqhMkZYzRVs63xhHx2q38QfTgI8
EinUssaxdF3sGnvqTrCjdyN2yiMk6VqO4y0RdKN+8KMXT6caNYlQ3hxtnnpWqgX8
e7mj2nx7zKr9sAvLqGszDOmgaq5jePRriP0emndzBmE8oi6oQc2wIma4fz5/SlyG
wY3yPrfBk0pG+fVGQheT+mtBzmOPYAh3I7xL5cNaJzszeuxwpDy34V9cFieIBMdG
GqHRemqlhYs9uZdACJbBib6nCjGuFBbqJvfAyJvATHhOcrevJPnfZZGSbpGz9gvk
b6LZSWtqXhB6f4B1kOgLZeZx74M6D7GBnb1NvKjveJE3jPHETbrJsuu6KEWjUyHI
dGVuaLIN0rK8nMFJggeTMvDiO/cJrxeHqu02Kp/6hZzHzui3uvdz2Gc44ufFEa0b
rKWCU0d5EehhgeEIZMm9CRRoTa4CidCwqyoLAwyvOEIJ5ezcvQ5Znk/17F4NG4oL
9jB71xqfUF74T8wc/ixp7rewBJc+qNV2XB+SlV9UkE3yGY1Jf9k6wol+mECYC4YV
N5y3pSOc+b3F9t5HqatAAG1i424wBzF81AXEp8Q5XCgw6m7bAwfbuqXRPOssnryX
NhXZnde3BwJcMeFfotWU2acidwcZtSxbDv8bX5vUDakRbYQaRjNNWxsqTcpsWVYx
+hGrHtk4ex+l180DI4fKDHHcn7vejaSGe4XDfW9cenFIsWz56pP/q6R4r+JyGzIR
Iteng6xoRdNUPjNS7ETpb/KvK7omqe9yycGOnGpQevUBXGCSIFKv8UmEypQ9J0SR
ztRvBAibDRNCS4owk1jsyoNO3AKNeXCgdKjD7Z9Bef62ByTgnTOheMEeolpdni1w
BwBRu5UkoNI0lrRadMjYWdcyErlWKLrsvl/EhHrasMwrLITMiQXfUizNXCbvehbe
cliNad6x+L57S3C9X7S4A5D0j3vuRBJsQUu5NLLl7fHgnXTuR62mjE8e5uaMbqp/
DdTPE7fGonSXEW3LOOphLwbkqXjoq/6vYENcYC4H1AkMwm1FjSLxk53m3jBJznd1
baMDX/Cv21AiQ+g4OPKvHXGE6gWV6vnfYzDRT3r8viBVEBVOveIWJktQeR0JeNJT
m2+hjN54XjenyihqBD/i3ireTTUWz6d2IwsDl41y0gnFTg46AwGrPre8hlvhBnJJ
hveuEBydf/tx9gI1Dmzw0DPoovvX5fT+3YK6V59OeGSS157ATOQU+H9X4YJdAw+9
c0WHYrwOJifGX//lSh7rdWwSF7YYQ1TCsDw1RYoAY6caadx7UaWImKbDEB/MS1b1
avurvg0Ru46Ri/WCh7bQZKv3+MM65suZbR/X/J7TRT6NCeKnGV+JUWNUnTayQXXP
HE9yVChKRT4uwKCeFtI2BrNQiALrle0oSnhtsH5eNwVT7JeacTfWroEe1DJ0+DBc
Ae+25hMpr+HAIq9q/yLIq2ni5FNrSubDZTQZFcRDRU014UsZDnn9w3fIPacT7FPr
BsB4yMAWMv4Jr0LWzYUCS3AhVhajPx8zdST11LgeRF8fiR03nTv0aMq9dSIdzuGG
xbqRU5pGNcZPzxDfr5DYCNCSipEytP/bmvBsLBTtK/hUK99gbcsy7zl6Wy7dWOdI
WlMWYqFWBxahYBM3BGUSbsPZvtKBZ/UnmgML5w9ix8miO5x66/2xDYgioyHQIdgz
2QBGIxn0By+UqokMjoyP0eAe9+JunNjz+E8OSqdOqJKNWGZG4sCRZ96kC07L36IA
Sf88yqVRtzwauNS6XOQtAPgLzUw5zk/ExvNkILezrn//dsIFbQ3l7bWytjDF4VzZ
3jt2xqp4A5HzIp7hN3KsimwpEWBByGIde/fIIv8hGQSINGJNgHevmsLwAfX8aka2
Y4rEx/tkeIXG36eMp1Bpe9KjN8lKNza/w/MswWImZwsF68XtTby3yxR8mA0jcIIA
dElm3A6p2yBcmOvWVorQV+QdViTqeEqXEGpZfK3aLiXWv8zNzeG+syCaVMYJbL89
zpgYv6zOlYnGg2ZnRaq7A9i3PzMtGBdnwRMOoXsNoy5O71utCCNRSWSNs+27EGeo
5xEdmUK46hsN0X3A7dimqDaadUdhucDD+riFPCNHTTfjeJewzKicW9Gi8ATwyPQS
Wq/Rrb0YxQ029Ua/DefquVyTFVTgXnKSnna7cgNJZpENku63fo8WGdpWGYCAKBNW
kszd6hiCBP9Cu1fF9wCMlu9tVaarEN8vXku0jEdhioAZ2mzC4VZnC/SJHh27fwFQ
h09M36JUigYz5QOKj/X5Lhitxe6Ti36+dmmuXVk1n49p0m6J5pbfk8FoY889rnl/
r7YqOv3Aa6RTvS2z0yxq2X2JQXNHd8xDzybMj35XTBptnoCnBXwhm+7CiTU65oz3
SeV9aTbShIMEAsOgBP5GRHTulJn1cBNTD1nnnSc9X38rFrfP5p313DN+zYQyTzbC
o6m5fPdVJ7bOhGK8DFEBcHve3QsFvrf6hPkrb0f5ddfa2zd623jEm/wqmEQnsj5k
RE2BXZ0Ca+TK7r/CpcVtcugdtq3q0hZERrBJEcXkur/S3gKgvoeFg8JwnMbvwp1B
ZLSJmsFu+5u1HpvmWbjEYBNehg7lWXO2s2oVR318y95J1gvnu2PF9GH9/r14be/Z
jZY9v9VW8uzCQkMdC+2TsCevkHXqUDwqW6EbQF9QKxyK3gYVjgudqQVlNftKG6RB
9j53D66vMs/vJZYWm+oyWs9litT7Xsh7nA+LUZJa3+AWT/VHgX7DZ7f9+5BjHFxG
q526Hd8TtI6bwM2pETQ0ogPZ1cXfgnzaGcQV+runYGfRd2fRZOTjQTvkN7rSl/mT
mo2eJTb80r4d0PZtPkGMfI1PgsUZYsraa8jtGEszzSuKEPFRe/BN6zONbGeGuEV5
XiDGvdezBZ1/QDmK8Bo4/6YwmYigrZ0q3v5Psq0afrZiVpOzWuK3XbtaqskX0Vcx
gaSmgbqwAmMCbavzkicGwpZQxUJ6IYGJKcOHK8xUhya1CXFse3KX+8oBa0gsDSN/
FWqvY9AOApPw/54tjjTDPg62l7k5GnKpw+gI8xd/74iutJhElkD/7/nuUjRC0Kpa
A+BIf/I3PCxft5NI7c2AZ04te6XNMQJAH4Ofc6BBnopJD5zZ7zruQ/q3rA1IlicX
O07fBt+fZfCpxZdw4FGA0jXnUKxBLrjWncHToNmb2uGlETuI1NToeD6FhIIaFuRI
Ee7AEJHRThKlgcUNt9qBHf10bDq03QU+auyeopKB6ZVxsrjHeajWrEMMGcNiHp8I
vdlD0LqIRi9cOGigQ9CeUUVIhwlqJ62neajqYXcJa0P7tc9TDJZb2RAw1sfonqoI
rylzd1nma5p96zZrpOGiDQQ1j/wny8PBBi472EgkGQFjevgXxdJ6C81tZVECbb9j
7NYmP0PVWAN+JHT7YaWzQlDGSG6e+qa7GsiaXmRZPNGJXK4Zbb2DwYGwJGPTFRES
ty9fmA8TFefJc7xkYJFlUoIpXS41DsnzCFLxzHz1Mvm7S6vVYoQCk47365C9hiN0
6f28m8zd3gGDaOGv3W+XiRi0uhfLKisdFIce8xl1MghWzbYb8+zfdDV2pZVph2ou
FvGqxoNR6Vj9bASagdFddDlx7Be8Nh5zpPAQ/UZHsymec1skpu8I9ojC9wffsy27
sSFPnztBYt9xClULIwkwBaRdZDDeVVTdTvcT6I5kpgtOckw6X3rHH0QkntGPL74T
XU26PsgnMivnG41xEu7C9es2n/Cih4R733/06/U57UUyrbkMqFnamm/18xsxjRUx
Fhwxtft7Rw9fmNwrMrsSgHC/s5oFOEK7OKcFpwtLK2YM7OosqZ9SsUnEjTc6oMBZ
Rn4vj1QiZoPSA6zIn/qo4Ko653CLVWIU5faIwtglfMBLinp+6OLOWYkdAxmjPUrB
0rkahJlBNHqwuHXZyGE8E2ZQtjEnq+YU8rrDTIxTUiKa3G8VwldK6DjyxiPxKKxd
bAyZka1jC5nyCRPipQJdEghYdgqI2BZ+9m69L4unGbXY5f7qS60/ltaN9Iyr4yfa
sQstD0hky8DkLvjxqbj3jVSW0cvmkrVFI/yq41VJBcgqQhUGXCnUG5uxzGBg68Jh
vTTZkjUH51cp9amqzbUQdn5asUCwBUnaKqkv+0qtTYk2ZmIRpVsJE3Tpr1obCyLC
a9QoGNXlYkTjwK5kGoMxMiW5ChOLKk6kleB/J+Qpswe3HbXKz9ysEkFE0Emn7HBl
3umcNAws6vupt13W4uDEYt/bQlmNNaqFaAkxZUo35le0CpnlZoQUZgqakH2LfjEi
sG/WBYSh1vL73DJZIK8no7Yr8NIylOxU6/Z1Nvh/6ucNAd24l4zb3IXzKT/NklhG
mmfI10H7rnl2U9qrCR4PlCLf6qML9rmAsgMxu/w60/p5Dyyv4dQRO3Y56t9pIUJi
XwmwZQe7rNZAZHQ28FVxPejwTZCj6GukQy62eCrVRo5/njKwsN4A0yScJDNU7tM2
1dPATqphcB396PZ6ODcEeJTkdpj3cMvFecd8FPxSrqDp7FOZke5z+OVEVLonrgyV
ycPgetCRIMSFGmZOCsmkBaPOw5MM173LjURXxl5kC9NJ36Q2Dk8h9/OyDrBVE6+t
FlFI77g4ykAmKdN+vJJi3dSGl8k2eLRdJFRGMt74tw7Vr/SBvROVW4JjjqzqwrQ5
1gC38AgQpICo9bQtpCBodkdgsJBUDyoTjgvFZHbG5wKwYGOQmeqxo46jePqJYdcV
GUeYbPEMWKQubGR+37ACxDrMA58wURkfyb03iTQvyE5s0UNsbe5fL7Q7X7R5fy7+
HAVOcojOsz6F+4d2DiZrrI31akZQ+s7TV9lXAgTDRDwOOK/Hx9ocEyY7bJmTAHtY
3cVP9L7UTEEjGPwobnd65Z1qvjZZOSP1mQySvU9RXnIMSkT/bjffxcv6/R0GQNVL
7AxXaciWsgQcsYYuY9U0VxVOKyw7F4jXFHrmNHPeNAvW2sScQNtFpfBNA3m1DT5t
uDgjG06doOqVK2MZFxrvvHUQyimkB22aUu3QB4XpKipcIttPNM2lKSSv5rYgebO8
39/gnYH89NrjV8B+XhtmHlJofFVweocFgPlk65sFN0SliTiQRJJGMRk5Ym6RxoFm
BeSYtrdPw3nkTSNDnbj7xge9mi1jV0DYZmkw1YOAV6ERU5RzLZqNnyBYCIBzi1r0
oVb3co64pt1J8+LRhHDHeeXsChG41wewMagtEX4E0L8ODN1cfqMMzKqtSB96Qisz
lYSF15Ji6W8FEAFYrIOJ3u21uIBaOpRnSZlxPGXe2KWSvwdn+UWkKur8xJVi+8BN
mCEGcGpdZq4/LVn4WPlrec5P9DLH4X5N7cZl8ufe/Bv+Z99dFdZ/O1OOkNP5enin
+rXNFCdWRgj/Z4kM6H7oVB0CO4/DkCYMfBxfUCDSTf1tRJ3v27TUHZmoTlIPqQKD
CpLfYaw79lxhGi2zxIwmlQDJI1gV1f5PiBdTJHk62WUc7ik3KuUGGuRHvdMzBkXk
l/7azmbczLCt81yuxB1Ghd2ictBWlF/NaEdsV6GaJdMEpiXUpxR+MiCs6vPmmKdH
8x1gBwLD25b3Um0UZq2nLqzc9zAnylI+9Hc63mv2zKDEk7bGKqHIeHVBOgzYnDbQ
0pQtJ5qShYin2cKDD+i+OPWhDwEOj6U1yVF6WnRlatwZ+IwxGOCPYEn4F4/ymGd+
sX6GjK53zDrZaJp7ViUk3m+ggQUxcEJhtYuphjV5NFvOkqfr3lpC9K5XA27TVmEG
RebVDjc12rrEQ002G8ktsB7Dy6Zes+lLbajFLRSGg17xE/n8KEINFjd8obUiPDX7
gAFH4SoawkCvUX2wwwZyJ4ed8VoJ4NR58q2NtTHlztanxGt6PG44KQD4MK13uUVP
ft9WZyzKjCtbnjkd7vU3m6P7axOEJ9lVjsPqnmjTY2CbM8/VCcSuJsT1kOuEHMyX
28fjqN0B0EY3XA50V5oSjHilB519F9q8jvTRgocZBgQ0JpuMYhnWtL1e2j8tGZyF
Y2By7Q6bIdZDzJMEOM4f/SxlpmD3B0L9gnvOJrLFHJSjUZYFmkZFvHQXBOzjM8O8
03UXWFaxEKGRobST/IIumNtJOvesVkizFzBTiG6ChRA7lM2ldTyqvj5yXnqeTt51
2o7+mEvNp6XCj2TJM+KeiW33O5DGMpDXUXyCvjoLgvUPnjT0O5TZbOq0U8py48Sk
W2OAaO/QiIuyYhy51nisdvlZiwIPxVag8rAUTc/czS69cCOI2v5a60QTTWmdZ6Ym
AYfbyLOiacDRO/AVTY9EGRhRcmOk+WT7eglRRxnyJ5ZQlIQeUaX/LK2/qi47Wq9f
2di6zKq68pGXXFIyQiqOqwsmdjwGDi7Vgjxo8JvphVpwHNgX1dqSX0dOGYouwlBA
/7oacUm6MisaZBLER8Ed9E4jHGHmFeWn6dllZWab33YJP6D6Vuj7SlrLulv4TbuB
ncJfN7aO640TwRcMVM2F63SZq4Z807sJRKb7YNBQSNV3D551iNdOAcFd2QDsK/Cu
wTbALKn33+eOSlRU8iWXSwIpc6+XZqapPELIThgBWk+LVnR2KUClIYUsbEUWAbxg
GouKA57dr+z5WiOwpURW7axS9OQjOp7hdCQKOQKDevLPjzOJOAFnYRN00yFxvwzg
6zin/CRTd1cAvf+j0zwRqPFkVkcNbOIURLO1hKJkfyrN5rTRhP74Q7KI/obF9gbF
FvbI3FX2Sn6rJhrAf4kv7Js8RqznbxZD5OFOu7oAmiSzKQtZh3hUAOmsH8uJ7Ep0
lyeTR1sbCuy7viO0LOsno2UMOUFUT11GymgMvX/173gluEerDfHkTmYhCXaHB1Lg
TeLpCK/NB3YT9f1+uQ87QJueU0lIrL3PazM+OCWGjwhtrig4W668BnVzQ+Befkkq
FpNbiZ1OPWfSDn8wLoJIM6Y2nufgmYu562aUvEcp0P9xDx3nrc1rkQi+WC9Vtdgt
NPhwUKvam1jJy92qHklpImcJqutMdZgsek8FDvdzb8x/l3yOBqrbSnWKLeBPtca6
XZl9VbaXnojobZAE6NvKkaj3UV28hAn4zpNL6Aw51cD7ZKkdDzsUHfbaLp5kYAvX
yNhH/KZXr98epb7Y7Y1OcunenbQj+wUewfy09KprvCdn8bbuSu3kk4lVj0/z4EYo
7/c/9hBsyh7Os+vh4l9mHMw5tzfL5BFnPUFMMNPPdPVMH2xVs8hVs0PQL4DzuhnR
Oe+LfdpMbmKSoAKd5w8PS8ONMBRuaRsZaB1qOEWjhPMMXWhA9cwMXJfC5uhXT+Lw
txN61tHOdqdOz8g0ZykiLbJZMuPAxYM41KkP9F43ZN0BIw6kH3AoEYDv5utLHCBQ
XFwCM7q+9OBHK1x8cxCQU8+/FnjD+xOgexqEWtMZQpeiTNm0JPCytWysFjCJFimq
e7VyiFX+9526fPttVqNlnHsXmwbeMu7MERWdZsPlo31+RkiybSa2EOrtuISNJnSe
2pKNAPQxaVlwectccrU14HmnQymdCi6k0mtIOOuAu9/i+9f3UCFyu+DVjAEcg2Ql
NYeiDZeupn7zl9c5Es+QZjy63u1O4L3bT8OKtrmDVx5oS/Ikrsgs6wpvXLghauLN
lOyUcX2FARO6x/VluVWuMVIMAsjfRy2UNRKJMPb7X2V1c0FR3B66ffkjTtsoSap3
tQP6ztV3I+cBma9fq+VqKufHVk39Srn2a/wzKbH6P1moyIt0h4nzroj7vPCrApw+
uhYWsZB53kdsO5qfA9UT8xgAAQnQ7PIk0ZAylh1BZm/Xk9rYPEIqdQ4RY8RJL9O+
4YabUf7KzsNSl6fpK0t9y5VUn62QBxyYShXTL8aEKekjpmrqqs68TR5HOEPS1/dz
RI1ZEWfFH0CoWoWlG/SlqGwjvphD9ofVXAoTJv16n7Tla7taS0jJc4VEiIf7O27c
k35bbKHR42ZH3P+CpCHAemoRtvYo+cWCX2bhsG+JIofcKvTwKmgvCiP12h8orpg2
kAw6UriHd7L7JPmPi4cu6v+BXOn4ud2jpg2gpDJQxpN9hRnyMKICTpzHUv3FrC3x
qvIDuRcNDVFyQozUa8vWAEJzCo/4hgkmbN5nRsZo+zSjRV9pdVyyrvz9tgFTwIDP
z7vcZkya0La4VR3/sJemI3l+zCyvuR/NRa9ghGSDoRnI8YFx9PmLlj9vC1ucXiTg
O91u9U72LAklobo46iaDVDNohaUjSmr0f2D4q6IU7InrpFzWiO2SNiUXiqk/0ccZ
bWzAvJPp74r4cgdFF1MQuPVr77Pr9ST5PAEf7lMwHH3gSPyfRvLQtSvUvLmyXCBT
Q64NSqycKgCE9G1XUICQH+DTB1ADeY7DXVYkNj9kpoZgbbRCGcFvZS6z8rM7Lz8g
1B9ZLMe/e2i1hnwUwElZwORrP6kIsSecTiEm1M0tcNPI5NJmkFUy7PnpN1AQy/x4
UsL+YdWtpb86yR86YNtEoZr7m5AsRF+ECdZbFS65wNDXEWvyoIVnPG0UUCYpnoZu
bxl+1y8YDDVOsi9RrGS9dfLmhLZP7vcwZVgAfAP8lDvSS8+78RAAdYuilyPtQwlu
m5ElkDlruZu9OwcDhveIbWGK8AAJDp634X+PaWiXI7zw5jvUoI3YbepTU8QrWMbc
S3cZkwx7+tjtnvg1INm71bQZjajhr+TGJzGsa39uSnHFw7gtUB/6ZTybs7KUvSGu
OoWOqfVoUUY2sIHUmHMzp/tDyJC5yiClRTVO6MvuU0MEjuOxYaIQas43IwwkpP+1
/LLzQoKDg7C16qFnrLGqsHDNI2EZTQG6Uum8LU1FbSNHZxmb05Nfj1c8wucsmrcV
E2Es7Zv6VfbouxCdL8FiAwzDMla0ZfnbrMCvMzvlZ1mOj54/3IrUuszmi9WqhHqx
9S5WHM4tZ5kqCpuVam2Kq5h7JNqEZg+1jlD/bfeaF+PJanlLbkJrDMNXlik+99QR
lHdwyOdJTG1Q0em11FgA5T4S/CUa04eNijsWRUN9ZkJPHhZ4fzeyVUa8ffrD7d55
4n2oqS9IPB97DIcxFdxpTJjBLdsRdt1/fgac+JsnWAUUiuQqQ8SVYpstYv/1dafs
T3edhUMUIGdyVcD4j2LQhYoGEkJZuf66CIEbA7UemEjLmjD8E8i/mTno1GuiEJ+i
ojY7gZplqKLGddhSTUsyTXwMuxPviD7xQb4LLKSbPFCZxr34dGybrjAyrW4wzf+I
0hKh+6eu2dBca0KxHDwm4TlLqcDCHkA2HQJ6ThtPnq5+vFCw2R5l/zdQ5Rr9MR15
AnDxXD+RiStjqR69wlF0RZOopfEYkRSdYLXO/gtyJRI/S6XMQIy9DZX+FdPhV2Wv
jKIFW7opfZeiFK8l72H0asP03cO+C3GDLVLMtrBfOmacMH1EXdyHre8Ao5UdKURn
uPvLaKlUGP4UI/02gNpz1GhcpOXbhA9c8KFYCVsTQ99HNhn6LWLzFvFIGAKyhl5T
x9kwCMc14xPsQEbRFEQVkA9PmIR1CUU54+8AkqpzTeiiasS7kbZ6mQal2ZcdDdAe
bD8w26MW4tK3znhx0K84vx27P4R3fLyOu2q+6ZN6a5AHUT/qUSBf2YUDcWGba7HI
kBqoH5nhbkxzYg0b2Wh3Xy2O5dJDXFFvnoKlmSG+YP850QsKj4ZJNV0z+xTrA9C8
u9ocksX0CYraoB01ZN/CYiJB3fCAYhL1aecJNoSZswprmIUSDC4CyYcq65RP2Dvb
XSniz+2ysK4RanIJBmYrsEemR2F+pHC9XdYoRS6MLumgHzD34U8gAk0/SGJTAWvA
NjEn5zkbB5fH4Jb4Aq4zZfNU2XolX4VJFelRX2lO0cvYXzT/UB8r450CqFc4UhJk
4uMPAXo8GzWJyyyGH1g9DHTWQdUd2EfUcrAlY1KebY/h5kXYO8lVVVgrPuoxC3Ce
h1oRMbNabhsQl26mF+ReKL4j30RFf1L6yEEIbsxtQ9i7K1vaT7jOW/3++0cLPyMJ
zJl23hgxr5PziWaJvykddAZvmniNTnMe5Vhgj5kmRhJ35oqvbYlr32YW0IhOj6vP
N4T2H4OnF97LjwaXQ6eKZWkdn4MtVhfVp8hMflba0DJtSQXPBAgig0HlzFlQcRp/
WhFlDHnOChoK0d9nLbkp+H48cr0gtC8t8P5Q7ndaHeWXBJNBj2YYv+rTAPGo6ZZh
H9vTIhhf0gpZWqBshRLmFRo2K8Cyo+pnkHLVC13uamSqgmYJRABenIFaWwAODRBO
n3igWtpWOPVezmrlm8Cq6tB2Wg2UPzwLuiNWvoq9Jh5hPV8yVmp1SvecRGC4x/Sr
FA+uzWk9WaA5Oe557HE5dlB9qXV8uvCQjHRlKv2cfGshmVfWxFTvIXRykG8NyGsw
AQlDh3/XX66vO7Ip0fPUhBMEM04KhmEdvr1sTAWzCPSRu7K4mZvGUJzEZg8a8cIl
skNFl1JEmdQnha+9DuHfSkXkgdwC57Go/aHlxpISS0e438jKskoJ0ba0GcUqNioB
l2Hz26R5DNSI0KSb+ljOhUSY2c+keZzCf9hqN2NAIis7rqpjs2DkjDkADQqhUuJg
IOFlYTqJejeeUaaZosR4NTdoKPuQs9bA5HQi+Wk2ZNqO4iN5AVtaY4eU0igJ/hPV
GDt51JiRmbvKpzZHl2zCaWuc1rYpLOluEwXcUfP4f+9ciy4ENz69XYvmfyk+JAnO
d3G3GGbIM7CgF+F8nFg4hSqU091U6hBq6aERjR3kwvRKvrRAqqed8LDbAuMT6TId
bFt6W6wkbtVeO+OInbDMzFxdVk1DsKZDbTuCEwudqZuOmRllYm/4RPCdUohEZlET
A6v0GrFH5beET7Rj+hroAO+8StkOkplLrNzCjFTlVymQRi1leQGjAi/BD9tvfmWm
tGyIU8rbWiBerT1TJq6r4SUPXFC8qVpxcDBfD6ZdEXn9h7ksO+3v+f4kgrHUzsTx
UXeWGnZwFibtbaRcFn7EOkYz+eouVxHfyU6QFP3XyF+EvHbtR1AzdUq9ZXj0etk+
+tEhHqlWMMNcicg0mkCLyhpAFrpHtRyBdUj3pc41CbvNd0qLo2+aFcyy2PWkODqb
wOgyoJ491pzh0R4ImKnWnw1eM3dmYRa9pSRJnCMI2AkN9282ANGuqikER/N3qevL
jMLJ8HUJ3Cb2K9jQSgDGfY9/1V//qDVqpD6lyrHtXwcqOQRQVb6SfazrdOgkFV7z
/WMQkEL1S9n3fy/CVxQYxvsl4nn5y9kQ0jvt4mOi+wCcz9EDl7LF3Nz88B+V9Xpe
/mfHxRwE2Vg5qsTqIrM1RKxTPx2Xy/QfYxnGMsvA4zz6KizUuykpSC6UFplKDEwT
h3l33ZoK+JD0vC4T6eRgADaGfgwm9boag7zMc7HuT/BsL2dYVd8L4GWkup4kXW08
wszLZ/kGkZnug7l2iVEks/Vg7Af33dElVNyPR2uAGgtDln1vDjvT9YdWde4VPCvc
z3IH37av32hz2Qw7z5ASSye2W/SXB2MAw+bZw4tzWPpdGEx5LQ640lqhiAj3MUpo
3yP+J15K1fvDnKKprgzQnb6aDghKof8+MdobgqVIIYLM1tnsPXDeJoOF7wgWBm3o
HCL6DqnfNeBCCMl5UwqPd7A7bkkBXVbJ+B1kS2PHcehMkG7udhUF9gkXqeGupVKV
gXw74xt8PG1Z1CXTX5MlZFxefyRx0PnHXBFUIyroMdFSMY4g1vJTfiyWzJQ8NXYh
TzcOltBF9tHwuXk1wCS59N6M8VkWYBnvkBQ63Q9nPy4n4XrY7zjL+14v0dZI0M8L
iDF4cUPYvKCc7wpJ1PHaRChbgk37bZ518ACal6Yn08qcO3IU83WlxMGhlvh2E288
GKslKgfrD55Qch0Tgn6FkIrFWP40soOL70uv4djs9MFAsm2xXlE0XO7NhLwRVBbY
LQYAzM86SON+CMhtyvVMJTbh5YUGf72Bf68buHr8rJvZDhy1XclPxKPftwddyXd0
9Uu2isFlivyRO3RKLIYFRR1dUMWvJBxggZSyeghU6a4f1eRDejhQztLGLKkyeAS3
hBvE6qGUNLYSIBLRdlZjYNKbyz1/Eonn48m82OTcKZyJ1C+T8twr42TvOdlN4FLg
b7oza4+YpKcLBCZN4HtKo1weBBRs9CGV4B2RN5sm6y5Kx0WL0fsgBbLtUdQVYAtK
DgEEQ6FwtDQk0QwrkGxMKX1FvX6gcXNxFsEHMdWQgPHZc2Hwg/c4Tec+lW/1Xviy
XRHbB2pVA0tLyV3ssHTH7/EuffvOStkq5iUAgV9HuxjjyOpFekGiCtYZoiJvwRAh
cFub581GaJQlyn/uWwarxqBEuI8EUGKRXlcn9ui5pI5zfvnovqHUHspeotZ0e+su
EO++yp91NpBYfMqZhwxa1QlGI56nqsyS7WS0TH+7I2WudLMv65HvHiaVv4qJiGQy
q6dLF+v7tjysPxQZN3960GstEANHX4RFTCFjQUcr2hi7j3Pv50/eDwNIsls9QV3J
7LynXzUK3nN49ZLE3i8xlPMaAxp7nm2f9Zj9oqBiahBz3MEXfnUurbQptZTsl/yQ
3IOCtLaJfuk0f+hUqnvseZ/gF1f0ntVgf2LxNMoARKcgqa6AjKEiwkNh6HneLKzl
gnjISLLRTlj69OS2hL8BK1UVdZMMm2x5lDyCQ60307lEy0obLY2/DzHQnba/gaFW
7bIdjwbJH5TMXENMeOeXDtdB9K0Ra7GifSW0YALG9qCZFrpT8JuATVy2sYlum0Or
0XfzHvFIFJa8qLkwxKwzRdF7RZexJgVLvdsbUZP24A5g+7S2IU5p3z/PvOFDU0X6
+oAGlpYXvxmNWvbG5gPWiTF3h6bPH42WrWSPQttOWFtLnGBaLoemAdZmNl75s3gQ
klNs7inU8XuyrvGpx+4e52Ggu7FvAteF7H1JkZ6YMCkk2AKtnvkyI5PfMQAR/Wmh
lF61q0KIJ1O/m1ryJcMpKBxjzKEaMYvbtTFPEaZ4wPqniROFbFBfR/SmydCIxzj/
b9yJABVTQzizGN5/S4gZ9W1c5UabbN8QAHoFbw1vj5zUhYH5UYoN0uiSe0kGoHh8
NGM7MJvYV55t7wjjp1mp2Z1yYZw0zyVSjBcMkPPFjU1SYkomxXmd9rxPo8fJpHPi
XukpeKHE5COTfbDQXztND+TkXhIan+pHSI9V/9veYtMTl2DHgy96agiXj4tZwvxa
HyvHBOiLUb/BBFMHpLfKw+6MndXrthjEap5oz1pkzE6+bfwejI1hJkckJFyvKZcw
UBEqK37zVk0GIs/jxiQdmQvPPYbyONqewHFaujoENkG6GifyfK34BK7rHO36XW1B
3wUWhhDHRBpdsr82iCk/60uLzgT0Cwum90oydE6BfMUmMxt4B6L+hX8X0gFRb6Fb
wM/+d7d0H8+t1x4bU2W3h3DQQsfVnvdrvLnKS7emnfbCDi9LtGC5uNYdftN9NXHT
Dfr1B3yHF3J8m5jgBRItpoLULPq6QY/2mrNinEd1yfEpshcvuNn9zRV943SFzhlY
FqPVHkXGFfYrlE69xijthM+62OoDwFcF0tD9/AQOGOGiWAoRZSY+/HmFlHk7Dy0g
+uEAAEAjm8M5NVX62cYC4oqLudLT0t8tiei/OF9X5r0AJYcOCAjs30OrRPMyKeEL
p8RevIPsBcMUsqaTtfdXYUsUI2eoILCJf/lC/nNnqTuzOgeRwzHg0sJBKL4pwnTZ
/KEXQN6W7bYF34GwV0Hv6MZKrgjtwiVmU1QZsWPVHrJazIzHQlHH6y5yYWnfhMM9
aKrDGxFZe1XOcMbHfzuCE9zu3ryQavsbJF89UFUU1T0Uz96aR/SX6tHswL9BPqEQ
UlDZZoABtWYL9lL1GogrUWvC4xC+cII6ly21MpXp2A8HWkkvNwjIoo3xIo6TGc0L
PyrNt2KOOYPSZBueB8ITZB1ikR6WaJlBznc5PCGFb1fJyO2uCkkZm4Jqub3lQeDl
54bU8trccRHS7CWgYJgCjvAyToadqr6hqh8jP9fvCHdVTdFcFpv/6N3IsnyrH+U9
HrzSUvA6QpsMBVBZq2aTOA8HxpnXKOqZGf4NuEwe6Wt7okFlhAvGfJnaaWIqGm6Z
RfcDP5Vz4Xyxb+2U6qE/JKkQ0i5oG6CSY0zpeS1kZxLilRZ0irn8Nm58K5AVlbuu
PYVzAXv4urs0QWxpEOKwErESoPt4zlJSj5AhdnWzszQNy3dvOcJQ4Ze02/gPWpMC
XPqeYMcIEHsnqCPvRZzLW1EbDmpJIWF3VSHPrDuxp7ytRiy6zojoP4hnNysJHESK
6PoM4kSVZmVc5oRFTG5sYvxkPOn5IHW9xWpqMiYFTIlMg4kmN+QBxg2/jYOjVSyQ
gnoPmmPP+VOCcbhzyzKCHwzY0rPqTHB22ENXOzo+Ioa4NjEpHplfmNRsvm6WKPGm
bKr8WEnMfLIIDxkEeVQx6GHXdPFPiHcCSvWYMUCNrjAEFvpFNMd52hEmdOYi3p8Z
qGZJGod2cBZFeBqUdhhPnXxO9vaeaPV7vugE0VHiYFo9vXoQ36Svz/CcnuvCmF2u
57W5mIwdXspmFwrpFm5qYfULXN7fkZpOg8zJWf8tcN2iOoxC9ey/LQ0lPgcpxWyh
ytykKHzhlJrr7ifm6XICkutJV4im0L+uqCo4aVBlJO3hgS3cEUFtisz2pECYFA++
QnkGCGNCicy7NxNe8FimZiu4tlD6XPAeyAnaNlg0COHamAnGoa3OKVLYzTMG+pYc
qduTUhz8IAOEqXbBvtbdwQDC+sy3VISsbi0U1tMFckC9mkewOGgKTTTstSlUH462
1UUgwX9ICpKx/jDmhGi+U2DMQRgzLk+77CvpwZ0IfysxwGWWKoSnXqjnODzQO5S7
cUDqMccX63xtmniVZWF8m3hANfv1MN8svK/gHkCXPl7aSpoxgwyLA3q1djkXreRf
Ll17WpRs8dyxo0v3kmJ0elzBytPXMoT5BLnXcqjcglrUYvGZlaAjECf5HX2n1U20
5Pgoz1NmOQ0AU3CLBs3GUogEhwnI0mYyvs4MyZzWOFKMpWNzXVyKP6hikDBBaMq+
ycIgj03gJSupBpKT5kGw/6LxUnVksAEMORfVea6lpTFE0mma9YUxQR+TcVCi0w/+
AaHtBXX1uIe0eRvAGjHNjk/eMhxYxVF4ufSF3J/6eYs/PwIPKbO7bSvkTSDTZvYb
8MQ/E3dIZtAisF+ZoTbNvOYwAO1VK36VdjA94I64zP5UeLhW/QsnJLdBexjDHSJp
4hKKbqBAhyll+QUd2LVyw/jjP3MLqB02uJbsXQwb1iea00uq8AiUt7qK2c7pP4eq
TTbNLoT8N3hNf1nGWN5chWj4fyzH0uu8j+UzflRTVYdPC/Xiwe6UOgJFSwACxiQM
EGV/Kgae003vu8tCwAYVdKPCfHiCoVVMUP8LWebg3n2Enz6mgOh8fOFR4kIlQsgo
+keaFRRhVIQOY2g1g2PJ9+FlzYdl3YRDwwC0zzB4nZVarv5YbcWBG3ufz6mjFmrZ
qp+S5+euni955GuY5h+TrIKwXHsdGhqs5DCX6bID6SeAfyXC7pqApVX/C22khlIG
RWVfp161i3InuvQEmulFAmzaGjHJgtA0OXa0Gc/go4clPPKy3NuyzMAo3vMd/64Q
OcLBCfPnJaNNhCdtMUcfyrsRfTqrY61NpXrUXyhHC3FnTr5pkkhcvCIWj7DHnqlL
+HCKAZ2JtaVkX1ZwzIhIETXTqYt+LSK0uRTYKyGdkrCneOe+1LT8oGZqLWa0609A
gO+cnayd+WaMDi5+oU543ajh+uUoQg1JTvhVWes++dd41+N6bFDRFFt15sAVOA60
iCr6V58tM/ZLSquNqFUn1TjlQ7XlgrpMkG7co3FcgQjK7VI6HSbCLS6kdXHNs7Pl
8ztp21ORHfb3RFL5qXEMdbfvuQ4QZCr5s2DnED95bo4SK423aaN7TZWQiIDKb/7Z
1DEwR+fbIRPbnZaY18FbihOX7efwHqUNIWhBDujiQwabM0LMPKmM80BloVCejFr/
sndCM5sUpRNJq/cWGqe57HBJloiBstggDEDl0EiGgQrdCviPadQC8Pe7lZrhyrUp
/Fkqyq6zpEbAJ9/IRPRgr5F1UZHa+qzXn4SOvc1a+seJ5Bklg5kGhHHQpwaGWi5X
sR4PgdEHplEeeuqgcAC2rXABkwUxDFibiSeprTFkp+qHM6WyghktTJSFtkziVvdT
EdSty58+ZMad+n06pXnqOCN2FPmMY2czxUfn5kCfGnkkHLCR1DcZST0d0wXXEPei
SLvk08bHImmC+H1i91uHa0go35SBIsupl5mTwNgJdlQQXFum9t5MZApZ6T4Cj+Fe
hKeMiEEKGOqWzrazrd7bhqJNN8clRIfwFA+mZna4wBHiyG0Y0D0GEouBSDrcUQwZ
TP3tl2CiNjr3sXW0w4c90OBxLSmjPEKEOcoJwyZW7pa8p3ucQEEtvhca2wawgZdV
oiD1X86iAYq9woUZjo+3YqInu2XuwEfZUA/TM/LkRnRy73d0MZLsHUSsn4LWOzNL
Vk2uDIPFS5v0Zm7vlMFMv0Mb43EPDAw+W5hY9wwem17JnsvtIrixHXihEsk89isQ
BQBmH549bCA4l4u1Pb7RGGyE7hWyRmZJh6Zhnnhhm+UpaEIMaYXXQh2NBkPasAzp
ym5gv4u6kjRysWrch4TSwRthYQhzq5m8P4A/E/Ry3YC/RZsEBiGRF5ugxini9+Dq
xpezYI/J7jH4E0EWO8hHMpRbBXTYjJrZu0wD3Ac0rDXZuSC/MfLFLk+w0mHzpiQt
FFplDi0H3n6PWuaON0PEtdoCfyC1d0jqJACZBwwZ+GrBcpzE92i7agzdA43zxU7l
ntZx1dRgZCvFouMPK6UfRjlCtAedwVSwd4EA4gr0XC9fToiUh3Q3dis56HWrC510
U7/DCHl+UVtRn39HCGqgyZ4LJ+tieNEn75kXKPSHQp89uk4uNPdGXU2OCMKRL53D
7Mb1xHtV4M+aRT23JNnebwdqkc0brR88EeMrEzHlZquZ+7GhHXU8Gb/gj25gerS/
U6U9jXl4Hms0lZBC7Nh2UD6Z2AK/FBFAPOFoZwOUT9MZL5XbDICDtujh42m/4FsA
5fCVA5/3+vN54OMAtUnxgitpsYOW7WELVgGbB/g2l6aVXDLsF73/oAah7lU0ERgT
qKkmuJ8hqCdGOXP6ybTOQcLoYVxvEnLJhvjAWBOil7U9ihmHU7+7lkcztAySyR6d
sg5GK7We6A1x/eCQ1H4neAMrR9t4tXjPqEZpwWdFcml6dA1vUftWKt+AKMWTi2Vq
DFvHvJqf+6dSmPPdQ23v4Cup5arYvC+F7SlHAjZE0lYknbQby7NOPJH52lZ9jPY6
eYqyEJR2+c/LIDib8APjeKhY8YMCgPF4BM20APJOZZnwW3lxs9v0fcKKrPK1/Qs3
qBZ1L6Y30Cq+fCeCydEl3q/I0q8lQTNbIJGJTAI/OL/AgX7BXhSAoLouytUvz/qo
s3ag2TX//sgpGj9dEzpfjSViOb/plPT0WW5O3outZiHQVdRD8SvX4c5UUm6vMc0v
xk0o5qp36+gXSeVHpaFZY36U9qXHXYpd7H4Imw3/+fsd1Hniz+8QUOuwGPmYp/d4
j9GSs4TdjuHuXw4o/bI4+ZYYSAwoEzpYUSDAxi5ZTWxEASeAmy5BppPZkEnKZHAB
6NZFEEuGU/JDJFiwcAE2DAs+ZBMEZk7Bvh6CCiMB5+xDvjSecr7B5VH/cnUNvCPz
yD2X6yWGxEvwe5hAFUpFIeXi1CzBFaWroQ5o+dBmfPoK6TJTI2BpzG5OWods0r8L
FDPAUp3kRoybvBiTEJCr+YQ1mJ2uflgScG/jCHMgIm0kLecp+Z+wrzzxsv6OaeFD
4iOadx+Y5gfpnavNw/MfHVxG9/fQUDifFHw6c44JEYSTx3+ww9IC5ou5dD7AxjA3
CnlCNDIpoYEjU0zVFKoQqWX7vk5rOOuIvXdxdLquAZ77MD0IJgio5jQMd1xZTFyu
lPNuzZcb8aFQ19z8UszD8k73Ix/RQmvDyG/EfHdG2r7Xphqkr9FJUdO+eT8vYv9q
JmP6pTEdkkXV5NMH8TNqT8tgNas4DB7N2YjOJai0+pFg5iB6bGzlDqnApKCVioeJ
sgUE/fTh0yIOJDE0/3qY4IggUTix/O/POHYPUcGJCrsm5qboy0UTIGHukhqaGnex
mqSrNOYMyweAQBogvwPN2jwfzuZkdc1zOnZ0Anxwr1KBfduXqQ8sD+/6ZSZPd/96
OeMvSQFWOZpgIyF8or3yKPVBTEkb2EebD/nhCe75YMtlfiHzl1kN+IlP5AN5z9HR
LhTB7FIZgAAqbByqXvkcLwf4yH5fsmqLiG5rFHPM0Edg8rWVJYS9dILhmzLTYzRf
lKFAFxnFNeIme9uo7D+pmpUgklXCEJu2Z5HW+x6iYT6K31tp62SWCbq23ueTCP/M
jREZGnFmiPsoISbCX5rz/wYnzvJdL77d3M/PHflQew+nelVhoUgDaNupQ2H6v/ai
fWl/Uy+eL/4zwqU+T9Tc3Gj/+6FpMgY1cPK1ENo4fJz6vAsr83LDNsKuDu05c6qs
Hv83RLqCr55LXP72l4MziEdyLjanx/RZ6Trb7aKGIFwYqTeEDcWVzN6b1fUCp3U/
RFb9MvRROdqvcd53OIV61D0gzGgi4xYLRkC5n6GnfMk7fV9dcs1q1zZ/B1SHpD2v
t0T8EqzMHqDXcv5nf+Tgn7QtxGfD5LIv5UaDH8edr0byyiI2mOed5/aQNNeaTe2o
S3yDPIB2YZALKKioB+8prgm00MdUxg+QqnhuKDMeyh1tn07dd2+rbHDXpr/BQRpT
DnWF9J6W7cWAzQJoQ1f2MxEh6wtQJfYA3qwrpZU7NimM0dPQuc5my8cNUeT8fBfF
CmqPGqPKOoaNn1Qrdp3PYwZAmWlihygseW5QrCeH1Yh/h/PcPgtKBQ+wyqM0KijO
EuuQ0UFjU7c6G0PDCkp1uqzaWnZLbnF9wennVJQYVY0M1oIUPHJvVvngzCvaOgMZ
lspQSEKB6Lp8ftRjoLDsWBvkApcmoLOAlsgZOAJpTNIXcGKo0sUSWAsttz6uQp49
VAHixdvSgj/lkTtPMiGy9/evphcB+VGK0rPpmuPVYCr4mgfv/NpjT6Ie5OtZvzAO
YNHG6afdxW9m+T/F1Dy16FS3bu65LA8vsYKjTD3iunjnhfiVnBL1Pu1PTZF2Rnu3
8PYL9djzTynXttYz0xk5yU19aDRNJmCiuh2IRT0sMcsDcslZhvCYvEjR1rm1iQJx
HBDGoZaCjALCrmVsP1nX3XcQYPmhp3WrstQBGo8LkqcVbDpV1Ekwm7x/oaKsEmCM
duSqAaCXMOlITXkkpLxPi8LTDwKnYm8vym/I7cXBARbSCmYb4AgofiZxIq1m6t1B
SU+093krLlRd/6Wh3o3pfG41eDSAVPwj4pLCgMovD4rhS47d16AR/W+3M6eGZphf
IZ0dfNQ7hOdbgHIBAvWqaPjlFbMGXd7Lk/qQfLDEvWJCWyS17ddo42VwEohix/IM
GNFkgio1/xOmtOxoVMODk+EqMHuT2zVEpn0VdYjbUaZ/N5CALazEZlqqmnkE9cvp
lAWBasgzB0u7gQoFrQ4IM9xkhFrNBK9BbDTW/ZVw0OEcm+P/Tq9VAWuxAx0WXIFR
TNkXH5Oes6n2SKoPNqmqFcuDhVzC94B2iN8I8LbYuFHax+Pvm/Ou3o+SkA6U+Fiv
cc5c2QR6LOdpd5Z5w188agnHBJbn2xheDew5Ox7uLMyFW6SRhSDEOdOEapHFKGTU
7u/gQ3uMKOR/IGDl76/fE66wsqWZg0kt27TTrOZ3kyH8+GzcHYh7z3mPPjxkodHq
LHqYvc0WYB2JVuXUcdL+NR3oYl5gByE7tnxUurn0n6waAFq8lNBMIglJKn/wxy2k
pfMtyadO3X1PU01mvw13v7Z+VdlsbYyXdlvWhlsZm1V7JcPT7cvoc0YZNS/jlLHA
79kamuWmpoxA58O1cTxZKJWwV3NLnYZrM5QTWEtgz6u0sb1I8ztypS4WNW5hTlqQ
IM/LVQA392FkyF2+YiyM/Qs4mOVgJA/sYMZkxiU+kZs+MKzV/xyPaM56C6cm8w1L
D2lziPaOsRvFSnqNni7s1alzKbFeMCIr6O8kneqJEyZTE38tRfDfvcpE3LpKJ7hC
6Mm1D2QMR3kPwBFUZ0RTMNsAQLK8qhPKb2oKGN2hZuAWSvkjMedU0wmY946AKpxV
dmLn29Mt7xrNPh22XkKBohAXAWK1tcfA/SfIH+EK3iMjdFHE4o/EVG8fTpV67CBU
L3wXbcvx5n37fX90VqGvRGri0ksYRP3rGFpygvCzW/dNUxpXjbUwUuJEByhw5CEt
tEFcbxUD6elHl0QqtR94vMnwqbzSP8cR3LEW1bV60CyzKecURkQqdo2VFLs13z6i
C0TcuDtsYfmPuh2Ofej8nTttYSBGZ1TSOU/Jk0WLzo5kn5hkV2qoWPKcGtAd/gp9
a2HtK8QyHlzqG3rzGcUfp4+w0T62ULc2yvwSAEgzOsdQM9GFpV5qO1WzfoxJi0Dv
dZYSGWZg7BSMfRt0Vkj74MJ6hlyFsHXV7zzoE5DwEvJQ++shKiFPoGNLqiORGH91
iHYGk7bMQc8nCvG8HbzhFbJIRMz2qORMlSKGLw/6K57TglOZKXeH9Ng56NIxak6H
U7bNc1GqB/unmLiaCoPdVTJPFHO3AG717FCsVSUllIJpHFpaEjsPlpw9JEb3DIiR
4ZSPbGkmp4Gu0pxfI476JZMtZBNuInoxvtk0QITN9u3WNs565YqA31LWjyCI5/wt
bXXrL2fEPVR0NnbMfj//R7BkweC2T3ifF6NK6aP5B6qfQ/fNJ+mUAkV1r2/zbb21
FYPNw8YSRu/vIeQUCXtJWrPkjelH0MY06LrSTm0rzWtprLiu/xLZcDNcuAkTu0Xf
RN6YHKm7l0MP+b5qbSoCgF3iKc/4qLFKItqTJuvcgTCDLw43ouVJXCPXXw9Izjta
nV25aWhFPjptilYr5CothJK7BGxjk3nkFXoC68dTQzasqYdNKnFgUpLj0uaHddg0
TIcKlFEju/uBpQ70XK6ph0B2b0Wcsftc1jSwObTNmtFApN6LWUzkF07EyAj71F2S
YAq5D4RlRRUDd6NYWX/6Tc7WhxzSbHvycnxOZDcbkyBfPvbWZnWoLTiT+QU5/0WK
gl3KSz5wUrWH8QnfylHZcW6Hd+yMb1/f3JnVcs0qQUNZ70ZJbYLqcUpJAw1MX5mk
M+Pvw/JYMBunSMeXb0H7d2+1e7b5CFvTy50aJ3okg8mLn296Zr0QBcmW9uVyVNKz
rfS1quizO007+2iXrkou/zdmuYz4fwWZmsMHLkb36lkey9ZuA+U049wWvfUafMbf
HOUR5Bk/+MsxTOfSttuOUCksFS7HzHvoIvXuUTB92zyw9ZAFpZThmXKlDT3OECO7
SqTDigEecNt4tn1e5r24CUGn71aIwPhmLVjAe8fS+I/u2dncMRyiSb7lIFGUb2E5
1vJdxoE6mph0Z27Mjn46qU/OrrV14hTNSpZUmCuNuhr7vcJjTum79t3Y3nti11t4
pNAjPhOIWwKnlPxAuN4jqgVjZ9tPLpaHEEv2ORBU8C8gQqoZt5BWzcGs0+KcL3pp
moNkfRyeI3tajA9djjlNTgCnwOLAHKq07UvtXQ2T6qn5PH9TcoE01fmvTdhNzixR
Jfyu6C+qU6CbAd0DaclXDnGIGffDvMGp0NTp2mu7R6LAqK9ODFe0vCzzB8oKTxFk
ljETs0jj2hhFmYpmwV8nlTgN23oQ2kBKtY/VnIdboYbkKXFJOieUGDllS6qeHkiz
jfSjtvYiBqqvyl+cTL7SWIs+KNYo+tEVIv0qp8dh8nPv+ArJfxdcORm7d0bXZRH9
lsug1dTqcffHJGWmBVvv4d92vzvFijIAIEii9jHngtgCWl+Z2XL1PDhcWKJp0DGh
DlcZfcinbwi5XKGmRZjaoGj0Zyf41F4eniuAOQomojpxVrDSWueH+fW0JIG226ne
BUuNcpxwy6YDO8ZBYnwaTbSjIrDtovqgSMq4Fbzm9WanuRwhLOFk2qjpv4J9IKxD
rutbSmrxxh9Sb7/G99/3Do52ncS5UJZ9VkHGxBZDWl5/R5cgg3qRODujIa9foTye
aDXvYK7Ltr/ovrG7r8kQAccCPHX5Hl9ph9+cScFcWf4j+XewhkzCqSpeCS7NYqmE
Xx/X7G1dECWJGYiQtrvpJMJhE7fnkzgCUGt1n+rzHUE5rcSCkVimedczNJA4LU88
ubAgbX/rjyBFA0tenSOFALGGS1/oh3NTYpINYoX/ZliyHI/G4j22JhQ/5vWOzgAh
TDUNLRrAF+qnS1okfc998u4LrKOD8qEWO660N4AV+n6OIQFqWotxHkUtlvFb0hw/
4CxSY1pb5Ts4mlY3dpi+glTzimBaR2ky0Tr9fzEI0PjXJO1T6E2ALffnxmAEdsbO
EmlE/5GD66CuVNNlItCQGLrkrnbw6j7iV/mzEYQ339rbgjHDFirR620N3eN+PfyO
zgmgyYILstNgVT1zroWXa66Mkh+OfSABucUtFl8MwaNbKq3rYxoQe0/D9l92tJQ8
y44uhLooF3Hh1VlOGBbN7XOilwbE/tBRnonT9tenhz3Omjj/0ls9DHP20gZRmE/y
JTUcwE/giz0BbxoXkgrulSRVWJMJuqxUdAjINN0cA8+FEof4Aq17tdwfQEiUbzA1
uH6xD3JFV5g1p3lhcxYLcLjHpo0bgpaMvZ0jlz2KF3+LjKv7YL41u9WDLvw3Cl8V
SEZpcsfQ9lEmO8dBX1BNh4RILgV8trxDAN9ShBjNGkdti/nmT8BqyB46e6rPOk9R
ClCs7WhoRhaUr3IeuVNFRK7DmAW7QaXvWQk/EClJIc80vKy4mwtrxDMQYP8xT8hG
vR7EvTR/hL65dfDoJieZOXY/vNlEHMb2xh7SQA4SMvhwg4ZULFH7lgpW4JyUACdr
Gp2nwMScLvc3mxQGxlX3mhxdHqcdtQptePCO2tOckOKnYlX5bcxUjykZfAwDCmK1
qVhSexwgMSycTtcjcl1dA0J44nAthuH8MPm2vgKOBfaFzkd8HSDa85tSpadv/GUA
05Je+61dLu4pgwzjNj9P3LyE9udHSUb1o8Yq1A/vkBPV1I0pw6+LZEy+KezsifKg
LpsvY0nUmevU+G0kxItRLolRQcnugeOGdQYfTeKtmv4SEmP78qEFITztIJpqBovx
G/3FIEbNGiEUWzal6r1NJxkjaAY/E3MAtJ/UXoPae50aJIbYVZ7MU51Abvi5fmfn
9KUjGJ4elU8xKHlO0jtRzQmRa7UsYtnSNlliII9KkZHN3oGKEGUQad3MWgmISwDW
Nbq6Gq/LVm2yma6DBgNk4fCfDb0wYa9FapHdhUaENzmWzobZm3xKCw29MUPw9HHy
Sld6P5sEJgkwV6bwGjse63jrjK9gpfVwDub6xc0MvvJlxvAE4yUEyzYmyJZ+YY3w
b0HOt5E/E7S6x7hCflDiWwUivcE5xfeuhAMF5lbJHsByt7zXfGyf5T548Xw2HGbE
zUOR6LKrKvLA98Wud2BinXQPaxTOuKMEBuHh7hTheqeCgtrVsj00DnnQ4wvZuBok
S0AkFFp/6KdtfAKdXMqVSsA73aC+V2dAV7nAp4hiIpbH0/mcTr1rpqyUizoNKpzf
UcaA8HEk5MkoLnPsYW9XmMgMnE9cWbAwQ4VqP3SBZEHcrPgLwL+krkDvPXdbvVc9
aFypfr6ABUtbMvhOgNgbChdkU50GK8/n+j0+wvatEmTVX+GNw28HhqfEf6mwo1Dc
JJm32yW/qzuA348iGWRFKHYiXX0m7bE83COCDVMSdOwQtTKH0SHm7+EI5WV2HDbp
ejIB+NDpOA0cZoF2/VJbtH+gqlymRrHHd8mE1VToabHslDwXIk2IIq9OgoIuzxCC
P9xPkr3GMtTMmkfNFq0l2LLndnr8yy4YBgORlfKWGOndC0cp0tWNlchw81gMKHwu
AyB5Xf0ZAzJizEWZtOBw7Ld+pxqz6XKwWFe4N7fZrEu9FQdWDDpzwvZoGRFc5TV2
NePGgc/FKF0ZQ8UbXsaB7eDqgOV4WVbdIVZMxWZA3iKwvj/72q7lG2vM/BIZ5z+E
4fDlfe5nZKNrlOD9teC8O+j0kHatwvaEnD9Wm3NpRKjUnya/iOC6wYQxPQDJn1LK
wIH5ViDvKZ9ZD99Usrbb91dubRnDL24D0+3zE8UWPoyZ+d0CfKKwjMGqEupa3Rge
tkzskeYdxFq6szGZT3c3FBsmOjhhw7B/yYTlIqHWoOAKSY+yvetb8CwU3b3M33MC
wrB2OcaXxMNf/2Iy4mBtIUkqTbS6/bXlBsC4zo/2QNMyDx+QDBXt10EtE/S7XL6X
AZZ0uYKyFhRimQkjOV4ezX+BNibrSfKPRMutQkclkxVHAck2uygJziO47MoDBMCE
FInf7ouPcJMi6a3SfFGdbueJ2+r8MNCXqbCl9JQJR8OrmXO9NLMK+FSUWeV/kRaC
BdSotMJUf4CKa0bKp3M/kE1CI57zBvqaLk/e7V/aoX0Z7wk5MM0kgUMtsdm0h7YA
RpSuAD2MMFdKCtvwjYFhXETYHszjo6jGzNz4G74mXfT7u50MEpzgo7/SlAP3N/AT
DaRYqo9s3u2IuNNwFIhwTQgoRiihw12LVlxuqodHKbs10HhBvnvp0S4ocDpRxmHe
sdo7jCybGbQTuYOUB5UJu8pVFJdmF0YsSIdZUU6Z4I/iwY8Mw+cHZC43MrL3J/9C
jPeWlZO/iV7VtFTVHjR4ClGmCLEvJibzbtXjixJuxK0qxOzWLeid0NB2Bhq9Nfjz
JQ/NcNuBFA3UDdxCl8v4OpEsIPW7LpCPGjby7BVhDBnv0wuVBulThMqrQObHxGWF
EpZyYSdGOf+UKbMc3LFUo+6TJw2xmMXK01papd4xdlJq14Sh2Aew3vr9maQ89Z20
xOds3bfSTFtW0D5U7xMOc7nRFdZT49Ylg08HTiGczAN8bsOSEGS7Eq0L7JS5wjDv
AnMUG2+19VKgcGAIBuuv97OUhLkoe4BUIpcvSPmbEgkBsJvsPB5ZMSboEvlbwiFk
ojW4AHoI9F9U9xdYmjHvaH+46i68hvSenrqRIjwerytI//ALzHL0okXEqK0Y/+nM
kNH9hs1Vog8Qb9GRTR3AIZrquSLHp/2nwMy7BRfvKeCiJB0aBtpv3vgLRZVWUIBQ
vnqICxzyvdL/3T3d/tCYP1kpNXmTygOdrVXOvzMT101izwfGBavTigUsiNvKWbKc
Zh8ydoSNz+gHR5iDtOirXY+CpM3LY17xzSHwZUKTrRe+pGWZxzfEQGv8FLfhBuBn
RErym7trxLTidDr2npJaOtSKknei+YL2wVk3t8hR07jNdye99bZiYm7kS9B09ed3
Mz3/xiMuy2k+UBurvgquSXd4xPxk2zQVbzaOM8Ith692k/NQ5/CFK0foN1tPPHcl
CopBsFEV1lmp5tLM05Mcb3SCXS6BBXdxJE3FHNuzCRxtwrjL+hwF5OHr6yhVv+Ma
0pNcAVysG67NR97oTaYSktKXs838WmcKrvQnI03pY2J7XWwTNOrKlrEyRJxv1vPs
HGRPJRRMk0ioIH3SVhL4Wg6/XdXXslv4SFKdCZVsrxguF6r6fM4fix28zdtgjcvz
hdoDjxZE4h9/8zwBW2MmGeJQjc0of8Yplg1TfNKCFJviD2XzJlg7rXkP3RCVu1fE
PPcYilNd+C8y9kZnCRnoGjtJOtKUXtWkOLDRbAzMfxhFpmXulJDBcoD7AGscwlI0
qqjK6VCnA1txdEwu6dn31FqvC9d++BmQ1iZJ65H+pOCfHTyWfXB2EW7QLHOBuCum
kkkpGmR8o3pwjwgP2hwgg1LW9S6frS38qP0KFlUY/AQip2FVFapk7iQPg7w2zkR+
Ph10N68DT0KWQfCFZ1H5jT5823HtULJCAjo/NnSEv5w5tfpS+RiJvJImnTPiu7li
YQDLqh8EhQA+FOSiKzbA/tuUekIHxN/HvocrMW3OzDH2TBnb6hYuWLOyoXUttd61
aQAPsvMlzAeOf512Z7yWsTaKNnyr+4B3J2vI3W7iFYoQ/mK67IKqZ76Dc5vwov0K
XeCKxyIRsjOPt3ceLyW+8OJZnbt55XAg2a7BdB7XonNTzU/lufa4bLBXrEJ/G2oU
uY66M0yXmkgwBBxxzVP6M57xt0cGpFNFRDWWpEtuVP2Fc2M5hiKjbF6i9JSpU0Yk
EfKaiP4+lF623JasxbjuoaDQ9fwTMF78ea+9tX0T0UMgQ8vCKJ+ee8XyxI//EPIJ
WszOeY/ks+a3OKDQ+VgLgacLFOHkZPrt6pILXlXRSPP7hX15oBu+mFh5nKmT9cNc
dfZMdWEa8bQ2wqORZjUF3ppXeWXXo6rpDo0VHqeqGTXERBLS0gcZjZPgY9hR5i/n
Y2lGYfLDrwgtPe5qdB6ChA944+X5dWllNH8OOtqMqdokFN3MHW1EduYGMVWZIqwn
6CAWbmN0SRY/ruNmHj/0aSZwGvdZoYsPibP4GeFdCX57ZL82cWGZCBdrm+umQc6+
sg7v2UBMS8v79JdvUdXc7FUOrvOUtLFh14aVZnef4uw43UorzHcwYkfbZ6DXcfqk
/ns2pcFiYngO94JWfSRk63Kq0RJVzDe1SiQvsoKuvBYgaHsEcvz8540EtEwFDuo2
BH6S43fWZjjD3WgH+8+xl91QmW0W+xljq4xn5jibwULBz4gz3KzLVedNE46/asQE
CByI7FN2b8jCI3ZDhay8lJBqOGi9IS+faUP61SxFdMCt+Uwq6ZOs3p+jHQsnnWw9
O7CgUC9YN5FXi2qXLOqUpDvd4aQTtUjCzFCulO4v3WWRxV98NPsI4CkbrnDWSh+K
+4FMj4n6EcpTQEjR3cijIOLRF7pkItkLiMasyWjDhALRrVKYatde2ZPpwKj03goo
Z7pg49j8ese/D8gmeAsw28H+AwgBdONA3aSG+dCHM0yoWzfYwZn0OvAsvgvn4QnO
0jljukAqYTKWTTOkUXRq+0jxdj/zvacHIAF+FZ31n9r0AovfauAOu3bm4yeLyv5g
rmeDoEPTIIF8fCKTRGbKNVZHq5jWh53S2s75RSc6GiJjTH6zvlQaepV9Jmbgl73D
9lX0vVpZ8taB/PZl+GXVDoB8OHfK9VyAfdAZTPE1NGl9jMYOwTUSdrDHG+ZQaT7G
eWbjR/RmLnlBvL6NbFnmFZbnceIdC/9i5z8+1WTHxsv0kkrPLMqt4z0LUw0p25fy
oeGZss1z+5Zj+DeVfOAYte+07hU0u9njNHbHyCZvOzNEhwV+UOc5oXhtB6g8Z0VP
2PI90OQsoNjluAL7H4ODBqMu/zq/ci5mD125TGYUAYRsFkWDuPJ7oHQ6S+5I7oHr
o3My9T9ErZ7StLhZPE2TglXzMXU4F2uC0gAI0kBACdhkPfV1mc8Gs1ul8+TAVhG8
zXiEwZa8mhm2nbITf0inIL+oDsCIfykKkndVjzGW+eOAdvjfNNhCUxubKrk6rs3y
iObwqf8lsM1ddgJ2I/kWMN/noF2dRp8OJCousvzdHed+xVWlq5iL8ZN7ibbbIr79
kqvj72owMQ+nkTeYkFLbeg/jeWqoyvfxkCYsIvJX1ia0FNI2xMtsb8fH0fKEzm+G
3G0nmeb49zutv6VfNQStFB6vSnl3p8WjXJtxyC390k4/r14TFo6Yi74x57eg4Ahd
MroFY+scsEQHx7wMacEHhDZDwFFQY6GLeUzghBCWyVEzEehPesvvPEThbhwyVQiq
yeKf8n4Trr0sESEgJ9pQaz1HrkxD67uFPyU/Z+LEl7vZBgQgDbO1M6hg1HnT1ZQC
t4anEZ4OvQDzcWsLl2DNJmS7z6/0yvkkHrA6ufYegK5DC9Ng47qECMtRD/M5dDB6
vwmi0Oz/rQrwEkYTMvYSAJkhmJQZscv4rGflwMyVS8eYcFottmeIsvX/NidkJ4fg
ZB7KUl0OLavEKMGdzmlehHuM7TdK8PLBByjXGpddlNWeznN2QLk2os/ItJ3whPd1
qp1Ak93GDMR2B4H/ZjTnGFAc6yIZBLIpETHpsE3GfKh2E/EAyjEiavA6ptrtb4Nd
YQcLZA/wClKbBl6ICFoKgyiElhjyDf11FdNbpVrpN/P9LB7BBhsXwus0NF6bgcTD
9Av4qWKmwov0sjaEkX3Mg7B7MhGJfi7e5mbffLh6TgPs726lBwKioJkHr1g8D3gn
wdbhABhhKHWXQTZXyWCAWnbvmNU9lFYCyfNHZ7mHWsiLpVUAOVysMzoGFmqbvmda
sZi1M21gAebo23lbxffSfaJ0KfrNUurmK0JBmoBEF7JjJ3CGQASp49hvqdNrzDXd
LK5fhrt1jhtKRRVkKgw0m6jPXW47zeUEkJ+5wRbXrxSYwebiblTfnSQ4AZLfBjB9
M6Sewfoogt0jERlVok3eI624spcvilh3GAIB52fwN0Ap7acwcWVFCXnpoQ8J4Y4S
TplC7MqQQxqsSoUGoX/CGzCx9ECp+QgGVkGW25cTMTlT8iIsrcjR05jQL+9SjCtm
WkueV+K47EkF0cW9nEL1ONyYVm/Ce4hOJtoG+xF1rJ4WAy7mjs2M+m4/a+2z0tQB
QFL4fpH1GXXmiSnsnB7If5Eqg9GcAbp6UvWVHPlZEwVE9lLyv0XTrigMAasT90K5
ObTHGTyWlXGEEbZzAspjZDLYMc8wDPHpNeK5Zsj1kUnMqk/REsMbYSV4LaM47Vxg
UuB9gfzY2N+CfqspEMfLj1py3TKzSFcpQSNJXcLNw0SFKQy4oSmTWo4lEusA8NPc
liqXoKO4vDAA3DWO6T50QLrqIINJeCLRYA3LCmDm0VwWbB6ZIOrvivxbIFULG6s4
/wUxzn50WrIAkdHL9AVz2N4uCnuRC9rjaVj2lBq8lNIREPKhxAacvGUyqV4Hul9b
/XCj/oCgADKq0WhvkeTCJK127lkJUeve/ZBW5k+FhI3Ev4pAZ2DFaXg6hGB4Sozu
yNA2x9BjV8LtlUkqSBzR4eDhHL0PTxFUi5hrPLFuSUQq1rQHNWMmbtWtRInMigX5
Fmf9ijfpR+x596pLKjYa7QeDqJUZCTR8E/bDUHNTW5rMuT6kDBUQlYJk6tS8uxFM
nIyfY6y7RPV3CNuhSZ60D1AylwoBGE1sDsSPZsCpwe1vF8y6KDbNp7cXUzjJVoQm
ej+YJQRpfl0GyzGiBmnJ7leiKMEos23XcdZy0BFpcHHB7GP0+gDayacoqpVa+KAH
wKuH0DnWwjqNZDkz5ujdgcQy0tH+qqRs57CToUbss9Mpp3LerFa8Rn7LOvtIsoXr
b11rHQ/onzBUnWwrni2DjdiEnyG72vHa9r2Idb7mAJAiYxts6CpbH9hlSL6BUfvY
nhJLq8HQSR8Srj0/qRGWztOBMY6cZJRhx42lhZKuM5wqsrqY58hpWPD4phwiZFjM
OyJZL0QmR9VOsYDkzeWbJW96LLu6KFalgLjzC3NuoHukZREFlBnNhFibdBqC18O2
+2NxunMODH/3YgAXKiW0h8F9kXfOAVC1J2KmgsJnW3yDdVCmzooF95T4CnDJi5K8
t59diw99GBpZnXWoYHj3RBPk60PHO28vjyitNISvzUPM18dZ6vEJHEpyRvRX5nJe
sv6EiaRgzBOpIh9BqWpBH6A+CeAN3fZN4QVL20Vscw9V3GC8DsJcqTuyBWaDW223
U/yKam5dBo9+8PhPE4+2Owf8ZE083A1V9vTOwigCBh+6kCo+HYttAyx5w8PjP3lZ
svS8xg1WCOiheQULOnP+sAhVGj5JwO5mQtLW/Br1jlTQsrmDJ2Ss6azs91hUtC8R
L/f5BDSaa57Avi4GTq02+o7iX0bD8OiKE145gXTEH8gWqaBlRR53RuY4dXw6vuU8
RuCmcVgpCOLOexSSr0+EqY+aqIhlz6guXs+2X1d1PCd4hgiGKGgU7CuwWnTAQ0Bf
H6J6vwBAkLDKDQYrc41dBvrVdW7I2rx3NDquzvlHpiA+P3K+uylFppSv5XiMqhvX
a0JVzh3s3kwHab329gf7dgTQz6J+LbQKp78GdUDYbwh/GzEEBMGPttsV869+rsF9
MXjspAir5H12dFdllxhXPk2vFSyr6FZfBJrr8eNea+/WBxItx9ZIZo+M8OhAATCw
lpl06ejVoTyH11FKpQiJ6iIQzrdEzGZ/cd0h8T9YT9+MjpPOsSKPPtXDs+K2pwcI
CGrsCMpHSki0y3tfdYkRrZKkzyEfg1f+JVylQVg4qfHYX1t+LX/56JSXMQot9fC5
zqdJyHpjP+vQM6ANZLr+RhZr+Ey/rznvIvZfjOVLctaM0gXKlOdvPqaLvczY08ph
ZMwtCgjACJnEKBY5FwQf5rsK0+Ht8fpG0IqGEPA5ue/zPdn8VKQ9pls/5KijagJb
qhvHr2iKHqoQwcIIMZ9hIgwbonlWft8BkiFv+H+PerRRXVW8KFecyfoxDaY48NSO
cVlIoCh9ltFeb4oB709DWsUsFHCeJnAf5yzmT32cUs1vicXer79BPUzrHDNz4foo
1ajb4gGLShwi1bEzyrR0wdziuDewVHBg8x6+7iLGGcrjg3VQaBE0BHbqDfyutx8B
cPS2Deyh9y+HlzqN1hf/liq94MPCu4Ond185bW8SqOAO8spqYphFKEHFE97kBShF
qSI6W+ybHdoklCxhkzPvZRpuaT3ODSzDKaUew0+YjLzlfRGTj0cbUyoHa//GVRRP
5yxoMJlsC5sqtARrUIKKRsuIwxuKJtF5MfmIh8Dtb6eexTrwjlnsgjMHxpK+F4Mv
o6PssyxA4AUZajpw0np+jSsjzfWqm7qMhlcdyHmbsVONHzMjfFGBqKApNL7IYDnd
5xscBImHG+5ipQ8C71I4PdzajaHEXbTH5+EwIxD6JVVvjk4AQiezL7bsVxoVpNEF
lnPq/q3zE0Vm1T8V/FcR9MK/MlxSE3U/keoIodc87Ub7aQv07hzBb46H6vw7FW1M
fokOYZ8kJQjJPrE6SXvObC2d290FwqEO9jEe1gnZDAiLSdbloGVINEa1duqnL0bH
vZ0a0AdCl5sTLAVpDOQ1kKbDGoYuqvpmsjca2UJ6v2P7iNUv7OVCwQou+r3/Zdo+
vg8avZ78PNQEfRdg2Kdxmy12LC5XT2EjCKEI2vGrPxGuJWPZ8FHRVE7YDDnR3vkE
p6uFwvztZRq+m7QJ79n9/uJ0mKIW3kCzb1Y0JAmCCNXuNhIqtiIVSa6SKarqntS7
nBc4AP+/364Dz1h22FLE86WAd5GU0Kpi9POHT/5RwzKxApZHDfeVYujwxM+5mR3M
g0DHZvUGcl8PkqVxkvBQLDcm762hDpUc8Vn27JzMFfRFvVtk1N31u63EsskHfUqR
DEZs9AtcmUpEaRTq5bfaHWlVFtTgrdBGhtHudXJClUK3R6naCR3Sm8tq83ypZUjS
5Ls3rGwnYwJHfmszhJeUIloQBD9dwP8E9TmiTpG/SwW/iAJhUkBzXc1onXQsl3kF
J1ckUMxG2Ly3OjjCxzbXfNkN3YN8YpKQe292g7rqs/2CtwBFKznF9u8VihJ7eQDq
uVD/7/83h7b3yVwL5zN0bHy+JeSGRzIzNCoCk5qOmeseoboiZtvK+afxGfCJ2mWR
tDeogs0z/yqWPP8HAfWN7B5TZ3cXyky2e47+3GR2QHxuCEcQLa4oVEBBLh8R3mHc
3zAJq1YmOoG4CkUaBGyy3PYNIv/GJxRtdweOJ15L8ZXKZ5TyvpPi6nJsCMLtYrq/
WvaPlA3neoKYw+MepxTCE6H1UzRkvodFznkbHL2J+61tnGLfdfgPzPOt0/oH/B9Y
N5XMaRp1YTcmfA80rfa6eYLBXbXGFvaaoQmQyDtaZL87tEw0wgnjqH2tRwJFdY5c
jKPwA98b8KZmp51e44djkc4R2HtrgUBfdsUHJ+MKRxa4EJ82YG18KS5fX7dVzl6t
/Dpy+KBJ9KsalyprTBvKmHH0F9L434CeRzLgn1BHOuHgGhfSS8e76aGlh0x68E3i
aGBpAnEtsdmAoLw+OhRfTEdDA1/8zj7kOy5+e394ZbMchu0CU0Rw2gAc9frxvgnj
k97pNnSzcqoRcv34KuvcmnXRZAcJOsDUiIyWfKB5VI0R7M4ygC4H01dK+4+GZqAt
cOLId50PkSJu4u+KiIS3tuiFEC6oUt7eV+jc0x4VTF+wRUTHFJi1fSBqaRVPQaoS
HRJN1QGIDkuyGny7fIbqPr9ZjwrL1yJJUNWeomw1R5C1g16Ds4M8wb4Qo+wF13I6
0ktjiB8lAz6RxbRsw0tdk+ImLYFf+xQb/rGUk+YWTLCMEA4qk4aJoE+jeUsESGNC
7Hb4pUNeWVcxu3TZqhEIDAskOw+IR0F4GUQFYS+JyscexK3WG9Sv8Wl1fP9EnKdV
uJU8mCgkgC0R9nXMYnJsw03BayZ8KRw/dk+4UaA2B9JLqtUZIJPex5gVTEiwRG9G
Lgz4tE9/8a9Dvd3dUY6a+KLFyg5oW/eIDIIqCM2jRSEC8G1wcdILNPIRl6VVqZI+
aClc180Rwb5Z5YyIjWN3jr43INT/dAiaOFBF8r9PDpC8AK1tad/3rfrEYM2aYDSr
53k7Tx4km+nDYv22hWgxYe1mJbidDCOjU8vPAzV9MOzFeQMzj35SRXD6AN62M/FB
ryREoLI0WlVyHHM1qhVfiuHgC/aIEEFn5Y+2sdqHwHYQ7eSM9Q8nLHqOEmhu+xYA
HWFaF2oA6ZyVGpqy58Fw2bVOa7e4OoybuC7rZNhrBoLm3lLwU4oqjffN/R+Om0Ca
FiUIGytMnA+iPieEXNCwm7fSlLYeIF9ycWFMDWHvU5oHlumv5KmYGBzbzWS+7n7F
cphWh9/klVvfaNK9zJxiiauMzLkPck6vW9kyqPgKeo0WDNIgDbAcY7rT9vGGEN6S
dAwaEVZ1BDkgdiUlvW5d5rYYKwplzeuGzZ32Fe/fsEwwhBcVFCB8m+fgbCRBsCvm
WPP7r1Llx2FPpPIU8pC8h0fEMHryyn/Xxguf2I1ybLhMU/9OaWJFSrxiSQV7hl6a
DywifvaZFnNFytfKUA3wJwp8cU/ZuGZgzp/tnGxvG8uwTQbu2HOYw4F4Q0UbOy0w
QvUaYgqnSw43UKIi0GYPT+/Bo3rURtxVY13zwQrAHxoO69yx3vYKn/MPzsx7m0wh
Mk5jGAdiGQ/FMpDLPeUzM0YJrJFDRRXVxVPTNiqu08A+LcvOMBsexncmyEcgxeZm
klTIwWgfrHy5fwZQTprpBN6cernokaDLSVlQ9p5q5Ar9yZx4sHrJri/Ft/9qFgZ6
lP7BK1e1ZmLABmrcGYo0gupDAW7/rLZ4W+tpxscO7yPbzU5zFBVidczFxNj0YHpt
OXFex3Z2hiIF0XeJ6iXYEO3/r5TaBZhJNq1aU+kNrvvzgxcWpW1QhiK1DWJ7CoJl
9zAaCrzmdUx6SVVKNCIGHdBdv6Dz6lova8fYtvzu7MYSNTflkugirxTixPSWBAXJ
9AS3mf839fCyNE9b/qFJbJFWwIj18Urd6vZCFnaev0xpzWWYDvFPxxraLvmazXH1
FewWz7p3qTJwG4MT5uqEdstE03WuhhjOilPwO29icEMc4bh3BvP0wrYr0/X9pg7Z
QdJPCvhlRCkAW8PjeJhfx5fclmvGkLDWqEoxmZ9pmXNO0WJYpy5VmtNnzZBH7/5R
34D1q4sITTiuxhlZA2bLYFs5qUh9HaNzcjoebUFh1QciR5trDUeIK6E3zSnMWhYo
ip2ZmT0+0hxmhiswyGjZrPU85mWGIfbvuSO27AO5m9U2HGKqX2jWnCxTbyqwslR2
jxx7Fx71vDp9KIc3UlY/J+uWMFpRogKjJl71p9yvUOBlVMiZ7kMW+bhToCBJ7DDS
4HgvWNXDC4qHwDKhUIhpJu/TCoN2IqG7ImEIKUV2w/JtH9scBisms/Modd6Viq39
QIPC1vK2ubR/4lTb2AEUtryJ7rgPJxD3pz7to33SWmKaKGrW53StGif8ycCjRyqm
ApDbYUWubVDOmxW/IbD8wZvoPiG+Vzj8aQy2b4ObBQ0UoUm+ybipU6R+xNFdffqP
cxoD+gUkU75uA9hjL3CFtcZkfzyo6giWUidTFwFIV7zzLZxRdbdBRtLQ7YmJAPQB
YsG5M03P9CQ4OFC8dZTqL2K7k4ROakLyqmCJVbY28S5AOjslQ9fxCfUXVU/8mBqK
1J92hAFIkvUN/zk1q3wW2SSPsIsPuoK2eUyJojyVe8mqCvMhuExy4eoa8zEQ31x2
wFYVRyeVK/0YCQCJbipzyXMtWzT9H200yozXdJ0OxegD/3xZPGkNqqbEk2lAvczP
5KU5RinOx88cSk65+LTjD5Fh1dgNAaVpAqSCaUle3yNvx9Qz6fSmdfoJEezUHcRO
LMkGfdWSX3WUBSpGBE95EL0ZC05ycYkpEh6QJwheRnhQr+IaaCxg5WXGwuRJhrNZ
fr8CNhmCu4sm6OITf+iKYA8Kn/lR8quUX6XyDGEK54EFHbvCwE4fXkArZ/fMZLs3
w3qtqZRj2bJmjcIkCbyPXAsjcPlYkBHnPmIw4vcqrmdSss/QD4UbBGnOw7HmZnpl
vxZ7zZbLRyLnRqzk538FVW4Tx+FsLpUr0WLUA5+O6BOeC5eqcvlVq9eiCdnoTozt
hN6zDCH5Omm0jWofLoPsOAF0gyoJWQna9XYRcYFBpxU2Wi5Cbq5f4IXzID7l93hg
vafIchxvwi1pQ+yU4X9djaLxsK0K+34nFznIHPQ4Xe3Z4Ei7n1Lz8bnGqzvB2X5C
PR5tk0EXbr/NhJ33BVwvySl8fzxfm22iXb9SwLXovm/Ivje3s5KK+Iu1lh+IuPaV
DrnAWTF1Zfee/zGwKpEVCq/ikkQYE1JnBbhNKfLFJn7M32w14dv1eRg6QfOw8ILL
3VQ3XY2bUBxfi2uA+U+2dLkc8IkZVgY5npOrGJ1oBYzt83MbFdJXkTLsAe5M6qy9
CMZgRjIIQ6OZJSOGS+OTTYVZF51M4rm6o7xGvUMcjT0Q8meDw6U3hk9+DlacPv73
42ZXJVR7+iO8itXCMP3fKUREWYEthOZKNPjeNkvy9hGmKNCcp6Hw69sK5f8WUDwV
opiy9DxYxXj4ipOZhCd3UuIJcBdVHmB5J4IjFgeKSDrds88oe1eSJSTz0qelxsUN
tCcdUjlyX/FNeP6AV9fwdY2te0Pjixr4RHdCIbZN7/Hvd3ZAaluiLmUwoeq3HjlI
oT4ce/ikzBA7x6+VIqT524HpytUr1aQRqcT4Qmrz0KuxO751NPAoLNHYyHlFUzOe
Q0AdPe60y19WE+UZew0RJl7STd0B6R7Zjkws2OZqZcc9NayXVVb9THK9FQzAMx+o
ht9FdyxQM93lu96HYD1euTPKExIvc8PVf03pwg3bPb4yeyl0Hg9JpMmBegpajBx/
yEpcq93iKzHT9xqiinh6sb8dea3w8DnJXxzk59Fqdz+IX70H3uIRpz8ZkWtyQzY8
SRrh2wqOrzKgE9B8uxjePKEbg2n517bdGAM50PKonZFj7Z33lUXSJw0fo/L86Z+p
yQxRDZtGDsPwNCJ4+BULUnGxgcyuNQYxbDAa57ZQYdBIIOva36eeA58Pd/KBr6lH
STxsTeH1qVYr3wbnt6rDak3PMWTQN5a4rPkpGSWHgt2rNuaYQh/PhkcfSzOBtUgj
LqrP+O06zS/t5QH3H6tjolj5tnEMLL6TxCWIDnsO3klKCaGjpUYAr709chiZMtX8
QoahFbMWjuPQTwDoy9+Lsih25VoLGscnStYvObpmYlqfzQnN3QBXx+XuBgucQz+P
6SE2ZgZSnfLnivTjeT7ULCL839NKdIoAwqq4G7Hk4l/IvcnQbJV2LJluevQIBQOa
IJfSJN2FTo1K5tSuMX8Z5W3r/822bbU9wNMX3HrSAV2pO5gmEKlYig5PTkZ/aZYV
nZhPCIR3O1wvLcijusYK+RqX4biFVhacq078v1ASM9e8tDSPR8fvZETwxDpGgxzq
fg9/g1zjc/tHGHnLlSup7EmYzukFhkbkhI0wXV3g2dK0GjmlNbu0HcXhTzj0dGVJ
N3Crxo1ZBnlTDdGeQzp4MFmJLxUasdHcvb6/5V3FsfxsvLK7wf0W948jZ2O7ppTG
wwXzlr3Xrge+VFul4wO4/uL77V3ATeNUbhSPtouq2kUFX8vcVyCdB9e5jXeiCbYc
RaPJActLKpae0E2tRzhNcnFxsk0HbMl9A6ptxlXsyrAS/3Izn9c7qGjkmHx3domK
Z2IAM9w7FcoXOexsscbzOgPuA/Glc1tP094qtGwlm7kfVnJoboe8lXYPaQTuE54b
DrHxiEQNYl9mkMtUgOb6JaTfR+sC8xHAEPURjWQzThpFlDNr6DFeLgy2eKhchngP
uraZR4hXCGXvuitt3JiqCllAsh8DPcnp8ZjxqH5IIxDUdSE4/yzatrqJlmLAzskK
rO320HU6oX3c8Q/HmgjSvpRJcivn2QEvoBTS7fc/+LQ4rxquelHfeENikNo6e5Yi
rJ9FLniiRwFxafL8Jvs3r1anb+Fa7PSH1zKzTgS9P6iFYTOm7UZRs6Px75T2e8wb
B3QJ7fsFfkBFm2LIS3FQ1vF/ASCzQr3qulmpsXn9PVScBomensFyso9QC3n1gveU
Gyj+uVfmcT8S9E7GDp+a7OlSNvrLRQEAM4ZyY6uoT/pGRebCENzzQWRD/hf0Ju0U
XNzkLqKcKX8gnJ9KKzyiSlVW0JfkWG69g4yz0tMT1pHlXqCK3ahKhZnFCaExt9pP
wDl4xQa4N58lLf29EG7ZoVOQRLEj/zkh/RN6HhhKmI5Wk271uIjBOawDADGFApgH
+VG1pMmjwmE5dLTd4A523XkgNt7YHsJZqbFw+j7c1DK+MDBKGklfVmsMxnrCTk9v
piJYsiw2psddkbYAFGBDbBe0JgEUdtPIhEVZhM96t1RaJd/htJhtFgxPYmRwKxYw
9WOjuJA+eK4TZiMqeZrN47yHNUOxQ6r4c+gIm+e6DuySRl9FWWQ4mnkFfrZVQ841
xqj6QXzCe3CpAXHn4iDtznLzK7Tuhk7aHP5N+MY2M2lph20S1DAI27yDN/mZRbWU
SiScWAzVrtyki2RU23uKimHhfLmWR7QmdLsfYLTk+ofGjBPQXTacbaH51/PpfX/7
TleVauAkEj5G23kuY17+geR9EWWOzR//ctirx4fR+VqoygxmicHdVA+h7ajSvor4
SKhIbtYLGzbb2uQ9gVMBFlAlK2DKNEPm+B0hh7Awj1FP8MiUHMrgsyEftESCNJAM
Ysf/sM35Jci0k/1M1Qe7MNyNUzZpnCsmcy+jtOmImXp22SBAJvV8DToKHuXP1o9v
xOBX2Qi+mTd3iNCpXlKuVYZ/gbx+4lnqIuA9KQKkpMyg/7LfdClWU+0HW08xpsA0
oj8cjZtpFhjcREphR4sfudLVXHjTxeYqVM0olcZkCaoEbiEDRJH9fqe8pbb4v3kb
yPi+CN20Wdpu6nLI/n6wW56yDjizyDRv4/HqKGKGEWWeu0Sg3YyEPwEzhcx2srsg
8rdqK+L0xPyWLAFUpAWlvwc1RTxqSO061inCplOQcHbyQMEEVu2YqdIpjlbncWUa
D6GPKk1UuZ5W3sHdLC77PDjdEFoKZCjwZ9NP0f/4PyoJwNESk2FctGDw8TDWUYNR
g9p9rTjsSBC71pyKnTktkpTqWSDulkbup+MdcSR9Ah9k4v6N//h38tr4LLavNuDW
ESNtTz9c94bSl30/fzgrdoyIezLbj9nvF4tXg07UYReWQqtRNC3RbpDQr8brX0fV
K6zfx52k8DDq+B1fXJFzodkAqAzWtwc6jibRzWN9reDLGYXFlDueKzZhe6xjr3E7
iLv1eEpJJAoORna5qjoOKy7RsViHHwBOQytPKMxh2pe77iwMNFKlERgrK/O+hkom
z3oX3PWyb5sEPNUelB6OwgUW5yNPeEO09RsaFn9WZ+yn1dpfQPhO4XYlMvv2eaiC
QAyRg9j6U3yGMoo5wjxd7lCTPdnEImJxIgBEZbDF9eAmQl6BDXkcjtL7RmaEe1pQ
C9jJPsLvJIX6ENjurQy8NvvgTdpDxlDhFrptJQNIjqTn4r5XiZJsO7nv58nfhVgK
mZkCw3GwY2VahwuXbM/rAwHgpAnS95orV51P4p2lEW45OMdnH+AfVgm0RGTQuzt0
3EjISTn0Ug30Y0Rk/SRbUb5IXvPWQwBB9k1BJinBWGB7xtOd+V1QrbLI1YiZb0wN
XvEItuVUBmTDUIFtTQWUb2HNOWad2rpvxDTHyJgdYgiNN6n2NFYre0uMetDbrHAS
Tga3MMDbfCUlSdvSZ4e4tQg/hZe99tvgVJQNiXHviySSjhujpM4S1/VB+UFsnasb
eMi2+IOgjZhLEOR94kDf9hLsQOUrW2dr+PldEUHKx3vDCsDJjIcmu3d5b6SDve26
OkMgEgrWeTbDf9sX3e8VHo2I9ZPf4zU36XsLfS1PfbaCSqG0glCC82IC6aY9vQGQ
wfNE8NG+H5Wct47GutCtIWAy/r8y5/EVt8EDd2yLxCykNcs1KILfda5ObvZW6pHI
sbm8dN9rk97+NcBqWsYIxGQ7dvL07J4MWjCvV/MEMk2kIxEV07hJdvwcoKIw0kRl
d1ja9yyLKmf6F+MeLnxXnSvuqHS6c2uT4VU3WN1FwMq3c6rCY6O241sCQYmvHtpv
eR2OaAf/L19lzn+GUZ/f4sjAIpn34IzY+zfe80QFUzVBWt1MTEyYXTOqCFVVqBYe
+5W76sMotIOJ7oCNd5i+loUZ+dqeyLPVVnw2inSMEslIJNT5Sx4P9iDTflwOorPd
zBRjJ/PUosPj8kisFOnZOArCn9J0h/8Mb8EywYinLb/vaJLIarcM6TmFf3KjX4pF
4VTjCCRah3rCKFyZVbkDFfsAMBCORHkz1QBINGh1oCdjCNKGkcTjhEe0nrrrDKws
sGfbaUHwQw+eJ87E7Ij9ZIpI3Rbz+8ady40MsjfUZYvl6XbGWGPRWTnbz1vfd9x+
ipLx6bSTq2Y4AT/oe+COER1BbIWsfjuae8lLATDLGN8VjMolnG90Jr67krOr7Hte
30w9X2RhiPFN4GThhhvISXNGOhMH3+f4RQWONXQG2ryrFeA98Sg70DEsmyQjnTO7
XCGJioxaqRwC+DkNMUx53+IB12BeEeWhdIBCG+iUqziEeop0/nOquC6VG1Ip3dmD
UvuLU7g9zvomkeuIqaOcNtvbW62650+5x/BDRoNzpq3jIkzx5+r4ChW/cNRdP8wn
2CNFOvusvZX7sw1TPA/dEBGylGV/z1Yf2d1REFJzA5WQlo0gn+IWlq2GN+Kgw37g
bHBqCtUv5J2SE3Jsds0TPTlmQODku+GeGe+owKIxe5LVMEp3my+uCKiwtulV2Oxp
xiWaEvzBu07/O+GIZAfv9pnNQ5cp7t4eH62v2dDEfCIEdpm9Au3+LfN9RXqg66wX
Pg9/6yo1t19iPAjkdPk6NxXpgOrMz/ZcAQHEGs2AGDBbJbt0k/+TjvtBrz5donv+
ENrZOFu4+zdbGq3dY5yPqOIyMmltfPB7ehxKECwi3RmI7G8lwzGU/q42jnZ7pGfF
cfk00qk4dXqbEOFu4oxtWtKyz82oDTARsah8S/HxyHK1yR4bUq+X2peJhbRpgyr7
Lz6OnrNoR6jSHr0TMhcHMNGqe89UQJe3CCkFwMlMh1zevfV6QEiy+sOj8Jeo+JJ+
C7+niTksQvk7HJHHL7cMaXo64vqlgdua6qcHSyRoztqBupJuOwHMDeX6uKCswCSb
+f+yf0h7tU/N0zf5BwRC5l9WRFBxE010FzjeXMfW67qaGbD4zlvqBAUuf1xTAN+C
XKxHg5bQ1Nk1JSLrMyAmPM+TejydmdWzzV+dYqNR2cAiutpDn9ZVHdhrwZwuOPHn
HvPnMm5XLDAglFcKVY7SMW7wJLHuu77ETRnRvFucFPfCMFN2u1towelj8gyQZRQR
RRqFNHqw0pZMSmEdDgmgrFKBZuCNouH0hizRDF8EfKWU8oe12zxtlUFrZIoqBMwP
gTpdrPV+ZrpAOLb5YfkX9DhaT7ZUvUBTZ8ZHZihnQlFQX5yAMuY4ecI4dFGIQZ5e
0cyH6UE8GRmoWkKmCNF4gLetjexYNoBXUUUoHSph2opj9yRDjs/rOSpOEOol825E
uAiig1zAkmFWK8heSteTOL3wjWOnZgGgw3ylokKRAitF7ljGGnlVxuJTTC3p0QXu
jvRiyxAv9I6SaERxZntdWCB9n2qWi3NMOfv/5A29S3g4hW6OnqbdI5Qn7xKEdD22
htRHWvI4nuJMY6PnLH0vlwkF1dGQ5vAVap4HJRlZ9mAKXlm4i5kb20Thet1Ya68t
m9DzlhY1WAhC5xemsUNczNT1cRLN2Er1+DPPs5OpsPK0nI/3aWZ+x85doKUdw0Hv
d/tz6CcQMBnyq0eAhgaFSIsnFZk+iZH8teiJ+YdYzp8+dcKGs8bjRM/ZZBlNKqry
1uWM46yQUVWrqtfq4r31V2/Eboi+VRz5+2rSOeuwPekguz2jlzivj4iI6D3iQXNQ
FtdT9M5qZQIJBm3mGDwGma9SOhPa8lnxLW09HKoNjNYdMzVT82ilnauRrOT1jl/u
3OFe9yJ+yHLkV5VWWfp7JQSiinoi2m5QmfFe5FLDW65QRFrsRgyVUuxt5gf0pnIc
7/WWHsj6okLyP9lKCQEcuiW8CAYNNWFJoNoKY1Emsb7cNZPdcPUckd3Ug1H/MTCF
0K7sl8gFjHflEuX8yNLGpwC4mPAfYEdnzgQIn/jlaljKk2WzmxSmuO+HEurGBCx9
gWSC0bzUxJb5VAFuLQFcw3ETiyN+av+ctkGyHbC45MGd7BzOQuRj4asfT124sAYQ
waWq/M/WbyfO6P7rj0MHApgJsDedI8GzLHswoxVw3ZH1KSauT12Lenm9f28qF44N
jJNW+ycaeGQB+BcyJBlRNqmoClMO4gutQ7eGX4lPJoG496t72IZF2DXvsvAelxFP
lNzR4aMGO1KcsX1Wpu/rwHnh7bVJNWExBvHQGjbaNilSluF7MYkn54SlY+fB/xEk
0o2U6pXzO4JVsJzS/6LE94lTmX2tvWtHot+pYBVOMHCGR7sJWCkc4DEZf48vXLL+
09oFhToWbsrd6OlrYKgzxWjhKCHCOHbFAxDvenl50XLsH1U01OlqtHCxGHn6CNK+
pndltQsyeWyVCUupSUPcJ2X/HLAf5lNOTFE8ZoBwX94G+ZglMx4VvjFZV6WVQDpy
ZEQnGW2mpmvcreeCcIOz11DVYdtbyYPpVjW+pA/7D0cnzpTpdjOjAktIcVeO3UHZ
QVt3X3qN4huwzbbhmed7DxZ3flXiz3pJQQ42He1tY4tj8+UdjPseL+kjc1mQgA9k
rvjovgvjsKYzNty92MNYICOknEAWmMLIIq/Rfmns4slU7RAn7K9R3ezo8I13aODd
CCBhtn1JQ5dKfhT0NTQ6K2wolGJjXY4Q5vAoDALsBnqF0uUag2nqWgyk6KX9Ol3k
Woea3p3kCwBmeQXf6v9Gq277Nek4+cNu/5NTvzNeRFHYhrb01qTzNykpIlI5eARI
+weMtgLjixqUlXCASn6aDaghgaBlzw98bildZYuO8vyVuCq2qWFmtQJif3pLZSCG
QEJVItConQUmsLbJv96R0+kXitvKC18zVqw7UUh1LIkSHgHtwJqFk2AA9t0FiuJb
0gYzEQNzIw1GC+LB7EvkmP3j4RMu/ZqO9uPKFyS64RHsKF40u2GC3KFX1FegBGLT
cECKjjQFZGQs7OUjoszSSqabIDL2dyjs7OydthU+HAYVTPsqGz6SWBBy11Yjewon
Qs4QyPEvewHKBCZyRdaZdr6JH6Ej4WfUJbDmFdJQwWaEDWskXEeA31b3YY3K8ICo
ZEH1VyGxAi3t4LYqn9j/mIAMEhCQ/EKFsa+57KE5sh9z3Wv9gKHiudnCJJfi79oS
pki//kVdM2QgWLMlUouEwymWaToToR8e1PorEOefVTwumccU8NSNUYApW5/8iLZq
Az4TOr6D6JOybwgQ2XocFv+7yXSOX2mB50T3h/RaBjM0LjwNx2kIQpsPIYEU0OFn
PHuCGDTOS8qf9hyVfVqA3dpMACLhVxkUd0Mka7bbKLbb7+REhvokqBVcuzqeBysv
ngJOD9NF7/IFkxAdzivk2vHR78gTmqD7COeoMbqWkuRlbtEI44d77JFafrM1t2T0
YyfsVTiIK20P5tyFJPNO8PxpvFLS+fXewhMtXLJ5B9WwINfDJvkJ+G7rhoLU/IAz
rbeTiNQpVoAxY8ofJB1OM8y4L+3plMof6WDwKdW+Pfb2MA1oprDrg+MhNjLs5GQf
VPityLHfa3TWO7RPvMi0DFBgz34TLLYoJ7aOXHPcCNnmnY1toR33gpay0Uq5zr9n
4pm0xUiGKsSFYEWS5cDmAAaOZMqx16KvDXPYNHJRwKSKlDRIb6SmDWIjYM4da5jx
CjnzrwFpCMuR166n0Za0/JrSnuNqCnXUvw+Q6Evfmex9oXhkiXnTSsHw6bR27scl
najsCXe19hn6nUlmXqHK2X2Dsy8kuNndGv9IJB6sjsxMnx/Yzz3mqHiuTAklmlc5
fDFpF/AFLgQrVJCKJ9xc9wzvqYLxrtBlRtkiJJmT+gXe64+l2vbKNn5msGzTuaQu
j2F4FSGM9DjSIPHKQur0fTgCQ4cpKSc1mkRQFn3O0Es+dZ3bCgk9dnaoKGyLJjWL
OiZ0CWQoMlUA94XIbkD4uvSehsxbp+jx9+eH4DyFatUuJpaZqXoFV9IdaHrvqu0A
lR7TwNklMPjvoMnUwcIN6qVZm5/JPLOXXJANE13LQmFObUH+v5dBHdjAvc1X5LI/
UQTaAdIA2v7glGkV7SpN6rFump3nDKgR1yiLJHQ6aSDvtAIcGnIWyi1YgOuU/7P4
YuUm30AviJkclXHVfgq1UHY75263K64ODNqvxLOIk55xCHRn8uHTXtD4esRVLsgM
POjpcPeUYxXlAYbiYgSujxCRWb6LxcAwMTE49+UYzDJB/PDhlcN/Vhdbe6HVlJeD
i0ZGTU999BMrey8iTe1KwkQa3gxWslDXU6X+9jBZZkUd3XgkgaqvzaV0n64/w96Z
I/AvQbcHFX0hykw5wOIBl3YJUmN3Txwo4Cy1+KNmrhYGi47PmOw31TDiqyeuhFCc
THqLBBBW6X9iijU8ZMlLP/ukhbhL4X515QZ0rBSd0bP8eVWu8pS2YOlxhTAEzVKD
H3s1Kb8mEUBgXdKMixSqw4DjqN+4uNSdE0r8/G/Uqq8lm7zXBTJBo+UAgI4dzwkU
/pJwp/lWk+j1ZusNHwb8A3xQboBqJjsb71mKRFee1O6zPvC60GTvoQwgGr5BwGuq
Ldbn9TCYt9w2HaWIgoacc3/4YAnGR3KlIm6QotX55P3fyMZt/Eq+Ndkw+FzqkIw/
Vvr5ygOpiFO/gyvrhYhPNyqe+9xfKzcGlyD2APXD41AMbqAhsuD1EymeZSwwkoEz
g/OY+wF75c3b5Hu7qHPAf0Flx2ey7yx7Cu3nxVCMY7AVxDJ5RpiM1lPJDAXuW+18
Xw008hwpbd6L90bRSGnmm/dtr2pRWinlQ+11yzp7+JaS88VetUaWybVIR4Uoyjei
ERVZF50DPCu3wnLZF63bPXNf2OkzNmaJcHoFMaOa5UfBSiIveWyYKHkDG5onuA+7
j1/BpQsALuUUVa3+c5lU05f+oOn/VZqNE9uBDU3vCPUwc71q677hhV8wzaMXDPuE
WIkH7NYsu2dnqxFi3U/Un53nJuY3maxBKnjiEACnA/LyBaqP2LfdtaDCYY0uDcIn
wZrMX3uZwYGrxLO3qPW5yr7oOgWob/p62jMc3XATgUEpR2pc5FEYi51L0XbbaVHT
xWLsoj+YJt142bFcZQStrK9XS0XukohBvKWiiLBccYE2MGeSE2EgcsucVD/K43nz
PfPUCk35AqFf0eJkgp0ezibVXdHoacH2JJ+hYVCUzLDwtA/YkaxquGaPYMGTqJy8
BxaspNLrXGzTp8W/UtbvpF+ugKE+Y+pb8HXm5cGfJeiQtfe19I9NPj7ODogg20dG
d+pi9An99PAftCg1Je1Vehu4vZdOFouxD3lnNo+oOE+52g6g/CNPQWizb/89IBZ3
gHsfJP+a+VxIPvGd8OqMjJz1JDpzw6QLTZaPMTdiGGbeuhfhOy3LvW9mc89NVWhF
jqErlnwsL2NUspMxhCfDEeBlZsO/dJrW0fbEnsnBh2Ref7WA270F/7NoBlBouapV
HwIX2ruHW8XAeJdzhcLxFV+xYFGCVdhPDQubF2qHYpMhLU5C9bnUWI8SM5maQi7I
hHPXlCG+OGZKwccou8YKpjGzK/VmeEJv1E+mDMSh4XYzKxsgf7aUBLeah+1utJa5
4la0Jc7iYKVXe5L6ZnQWJ+7xuAKjjx5aG/tuQ8Qm8GWVKul01HYxgXYgwm4LUEld
oCTnaW9hTnlQaEkncURLfADWzq0eIP5eTAIrJ2bKFtRiDZTLzmOUV/CTF16/69iy
Pg69dSfvYbCtcZul0GIdP2RX9yqVIBxSId+uaReoPH8zBg7eWDABj99gn2lj+Bdm
EbFMzr4QenPIPe2zcfDkz0gq+Qe1CaUjVY8FpGqkXtJmmNfgIn3KOGJxiuoEu7Bi
DTtm8mcZSWyZSR0TL9upeEqh5f9hz3U/RvJh8LEYd4XQVGGVYrsaoZnmEFaptFbN
XfSJxGMiR/XMtmoQqoiceXRJhhhW5AcCxrwXYhbJ31quP6t/7C34i+2UhGyMC2tB
6XiB+iAAfYczqvMuvvWNjOc7mPtNZiRzCAW5u9litxWrf2Sd0kk9Ldxz6p5Z+PaQ
fPSJfG/01tK/plzh5jUwBv/TAsB+N6rKTy8lfjgiqWlBsA7D5gr+W0ztmVEiGXdj
E2Pf5T5x11nBY2+aYVXFo0pQg64QeAY2zzLmVxbLAywmft5jZK+q9VJMz/dqqNVZ
U52ns3sbzDueIRJ7ILLMaJ+x75orSWJY8clLmAiwVNrIuwOiRcScfmr1X4ciLkaO
BWe0pdPLXlaL1d6rApxgkpYeqILfc5st4sVQeVDzVqBKKNglfukbKgrUteBrVSwE
7MgTDKm7s4xTzYX/9Mk2w8Ds1o4U9FyjIzILq0j7cMV6MRsLMfS86qtVHaLVQIvb
guPWruquK3MAv+SBZzxSEgYLmUyW0+LBEvlgExqtqVddW1ytAhFv84qTFbzzUifG
+NdV71rudWaMXg9gF5jUxJhFn7BgcB4Eow0bW05+6e+g7Z7EYFIRR/bmCur1LXiJ
iSPTCAXE0/bChd4Sabilx1autZprF0iq7HbWs+AW7xCJf3nyBbakYGm0WvW8h3fZ
eR5bM3s6eOPAYsMZQS8ls2bJJ+mHg5ouAQFuS3mPfjAsdfIOVNCeuNfqLIhLdM1S
WTYUcZgmv7tThkl74Hv023ilwJKYK+nVSOwJ3/Brmk8YpLgONEuiX63K3H0o2Z2p
eAW0TdaLVeBShdNhbWo9+/hv7B/l29T2fW8w3+Sszxz+zM90SKtjIXN60hdf8StB
CxlqyOgNQsFnIuSn1xJWPNRi0/4OTbj3BpNmmUcOCkTkjxjXoiZJvNTTeVl99ZGM
UprWSlZI+ZyaWYhzcv3KeGOIv632140aeZm/FRv1pPe8ZQQaNMRI0LEE/0qKfcBv
ci/KT1GlRyTR970E1iWmJ8SsZj62+tXB/FxT8C5CRRUShxdY4MZG3hDAhlX+hDmE
1DqTwuubtVl7dDAj9ssdPdZieOe35TXvXoOA/eWen5Z9fBJbAjMP6/lIBv652kHf
0zj/nEfm4tRz1y2o1gE+TeXvyIfxs2+jw8iwy7vB/9D28apMRQ12hU+K6FndP31D
6egNDNNlVoH9ZzdFvtNuJRQFJRDMroRMdKIYr4kUtkgrUHUfKDTYwpBHAlcXegCv
FpcpPI63ZcUBq7swHEzXJ1SA9kLqYy0hfoYy8Bhs5bOmuxRbPCSMWn+XkxGB7V/J
JzZQwTdSRO/6nP64PK4t6AFYTRn1rxhIu7xEIKEL1Fvzjq2afYgVeVjPtCZIUbub
CoLuaoKRdGVbyzqCNfqG6SWK27IBs5CVX+aRJNJVnZxJDT73365NFuGUnZwp4Ygc
Xxznre1thYScQ6Mj9tRmQYCUNv/J9coYDlZAu1KpdAeqld/2VTIUE3efJEKjG0cf
nLRPBrIiAK7yG/PjRNQ0Adr0v/LSPYtCF96VobZHjZucUrAdJjS2q5MqOwVN1Vkr
navcqvYQ7B+v2QPnjY2lDI9mTipr7TCtzY4x2f4mzotsP4L5kgbY8J189PQpMAdZ
Tz/zQrIZS9q6SkqKD2s5urmBpO+TCaHwopkhevi5eYv6ER9YM6Ezn4lGZlnnTwy5
Od1MNfsJZPhkSXWTgIi4W+5ppiJ326hvuqiknUbiyJHfPI2ScD90WL7wfwkTWGB3
HJsDvXBtNfhv9E6i08zqzPK/JIBgJQC9FSws/IQTt25sYymHEcHAGP88/F5Ht+M2
ia+eUadGpKeXOVjED4M6EqCsmoNUR/F+N0fw4mv390UQRiyTK0hr+FhNANTFImH2
rB8d/b5BjO4Aa7aRZWZLnQvyScNnUDkcQdW25p5YQp4iGJVetOJi/9/XE3bfCJQI
iEScMKl1x5mfD2/QodJUhs8jp3MxmmkUuIMAF2aNu12PSU7W+WiD/tGQTj9oPNng
GMfjVrm3Jrs4fzKoUyOTZENoQAuPZX+eAcGj8YAFXPw3b1a5wYl+VmWJJwcbLkS4
Y7Y2rVxeH/1VmJeTlzaJh00LuhFLOgnUbygNXA5s4IMtgY8SsWymzI6GyIHfBTEU
ewDN8ueD0go5+Xb8KxHOVHfGqtqI1pXb5VlTp6dIZcbXqIzjh3zqDZFl8c9ajzgy
HoZG6jZpLQnpL+VdPgvxU+wTsu+GjX+qeHQksDwGZPPvdUfQDcx4MYjzfTccCHdp
PZyWVs9dTq/7GEuUmupZFBOk99mB2Y71Qs5P0Xq0iPqNTUTEquUXnSFlSRX+KOkO
UGXwhIegtZ7QJXdilbU87Dy4UvARRYkt2H/Jh6pFmKN+pmT4UOhyL8CZb54Zf/YW
HoSi8uQNGBww1TMWUNdZZYTVcyBJ2RRb4Q0Ikm2v+JTcd8VbZT4qBoXnqtpvMfNU
TWM5LCLhfsB1cacAqmM8M81sxg7XEffT0Df9ngAsEi4QlNYj8YyRdla8Nw7tWKSo
j1NLbQcT5J1vUKTgIJCMmK2yUtvkKxRXGiS+mkpg3bsKGMBkl4WuNB4lLva4aKY4
UpKsuHP3iXcSwhXqn9CnBoGBxxazE/UWMyPBAHZHZtJppExYywf+crkCCP7JYF+c
BCsTqrheHI8I/Aw+N3A0pYvcQmPCEzQQwVdHo6uxhaI8ClXorHmN6V8QrhuF7RLn
m5EOiHDasJwV3Vy4+6YUzoJtDdOgonXR7BRC1PLqvf8tOp03TQKfkWcWKvMwXr6Y
8A90YmpZMdlUlj9r6bDLLimL6F+Gl/lDLfVXHiGsniZr1xNwdXqKLVwpSHu1sy88
BVHKM6NAlmNKAyB4rWmIbAhdK6YfPDrK4Hp5yTFR5nFHGDEcQrtVudwwuvbnjTML
ui+7jV53g08Fowc5IKRfHSZjn535Cqeo/5oyUy+a7WeMjcXb/NawGHnLtDCmtYQd
SfWjZ2NX22dehke1Qve861t/qXN0TFGMoNRjOXFsk1SG11hX/EEuGD/c2wKJMjNg
ZbEI/LjHCg0e3GW0eoMuTA08UXNmCk0rHJgOTxIPOV0kblybDDYS5X+coXOtQu8N
pH/gZ9Xj+l4UuxN/uJ+RmJ+eBaPanLXc+TNmvR+a5ixT4iUMtGGRgMJvfonhhiPf
1AdGzPmbn7CXSdWnyne6XXbSwfWS0WMZqnfed5SGphC4JJapXyfHP7RF1iAJJqNO
kzMU45eYEZjxGiRdMTKAE3iZ2mFiteUDK6YJowYtgayz5V802vNTKgS1GRZz6+Y3
D4I3kSVBOOEGV3xRTAdeh7RziKU0QWFkePDskO0JYzYXyL1Rd2pRYb7ZwelV6kwC
YFna9gaRTcR/Li7C4YSlrJnjY0sU4HztnldqqBvs3Ze+TPMY/LzSOVnCanrYMCzo
ZU221baGoLpHAp17jHdXWn/Il5Zv3GgBnwaKhkjV7GOJMX2gocfYuJ5ruRogcdAD
Hl2qwYNbCUvmsxIPPN2ezb3LWErnHA0b18RHhVsULbvtM7ewe9J9e3mObIR7v1Db
V3VO0ZVoKOCcHhhCjKBoZgB/zj/GDLxY+sFx1xJpPUhWU+CJT0WR8p7A4TvDzTrK
xOuqD7LJWgSEO48pFzyahAakIOyrg4pQhsEq1q6jvLK1KDS0TOhbDwvW1Hd+OWc3
xlCREKE1R4wfYSYsgjOJAdvH2KhAShEG4IT0x45kUK+VjLoA0yozTa+H0SQFAUq3
Lbz9j2LMQ84u1q+vrrUcOsx8a2zD5FVQo1vWSoTerAEmapcQ0LeE8zX798KYgnk2
kDIFn0eIt2iVJubrssxCLZjuNBgiJdSyR026ZeG3HyvFRNuFJC/lQvKfQ4O1vGEp
vAAUjHV/IEJ1PsZWOvzJNQbnBZtwMoiHk1e+vsZIMycXb/hZqEt8YRrZQqWxQ3+O
fjlmj76ZdWkTuKE3CybBb3l9ZX0bbgr9h9t95Nzc3Qi7sYczLSEPs1lqwGLqW5TQ
tt4ESXdI5AW2Ghq1KUKP1vrynJou2VBSDNB2Lzd5q2GteVZmLeJMnr+FepazFFCC
EX5V+puOdXNcR+D10Ulwqor9zA83y0TBRbfHIMT50Me6XYyMfumOAlL2V2z14gJf
BYQR+Fn17kOneFY2pLmDbHhdlut+kH6fHsngxFVrErs1w4p43WZdkRVDkihDIhNJ
pPQZVksTXMBdLL10Rz05qHLKeq1CMsIRKfAdbNyX0fNozzREmtt1WqJxPOdBwcY2
sRMEXnnFWI3BwAG33q3aHXDEAquI3/mhXCWQ4qd5L7bb2U+niEkZfmALNVxQQyCO
Cp9HqBPUPnsphlTrgL5PNpoY9hf65kyy7AZDnb4mULtWBTWFotd4E35d/LjE7FXQ
wveu9LQT5pSndBNLueRjgeZUddw6cF2INQTulcYGKMdxjEXVjtrRqoJVUq8I3Byn
JObR0KM6NX+4Tgp+lbOxBHyBSiR+5p96F5mT9OAmU1md+ZKdpSSakap6YbajVWNM
3+XpnE9oUV/EaKFFpd+t6OwsrxzQPnBiEbRYY7BDswgfQbXgxddxIosiiWZGKjcv
uW3ATwGZyxfvMrb0oSRxbugfKGd9mILOrloIqrsyOxPtwgR9cnSOsF0xunSVrq4S
yblxZeAAh34zzSLHUgmilcmtcyxN5ahQ6zMiaHtIEru0OpD7/AeBB8noEU82+f4T
BMkOJXJyvAcyGOCvunKKOh3Y1GyLjnO+Fehf66hgx6faLQAX12yDBNHFdjttIvBx
DpqwJWpj3dz8JeTUkY0KVQk0rvBiNmp1ZFDaXhg7lxxIfxUuISVlBpvQX1z4kYe7
KzDxDaGXPbmJF/acCU/QjEIk7v0aUEYJlpwkUQmijWA2rxIZd393c7+ZO3QtXoFs
IWTZEIsV87xwknc/vK6yHAhX3CfQis0UTWF/nZxVkMY223r6Y7Z47B+gYVVpg+Z9
t4At29LvVKpa7HflcsvJwMELYPPo8x/vv/DZhsne2463fNtvQBeikqHcMmfAGe8l
ZQf5Zp6gdFTvKvGnF5EvcEykGkMNBS5UF1Ts28FuEsThrQDaV6FxVrfBaa7vTtmg
NP3aLuCP4wzXjDzmRxHAqFR+DcT16buH8Euao485wAdapqhvmp470jpapIDAsC/s
Re9WMwrMs+mhAIAoRNoXmtoK76uU7Vjq2gwpExcQeE4MqYs8TrdwI3+07VAhDYd6
nDUcDV7xJ2DK1IaNFEXLZOP1nxfBdFDrO4F21iWqSgPDETGtPGEg812fFRT5W52s
abaiRT0hm8Nhz2KhyyL3qa9ikMqSYfnEMNR/5anFirPBOjhMVDZxymJjUcedMNtV
qEoHGSIWJ69XglKdZRmolEFGfi4Ev4YySZ2snj1eeb8BupVDB2aDdAAGV22m7M5a
o7Iwsyz3g9M6DljZd8fXv5t/cgnuwTYldHtnJSVKkOhRU6fsu+RXCpdtDHTSMiaH
5Hbei6X+aJr6scQYSTkZBJoH2q2A2gPPEGY/JOg5gQk0NdR2+gC0w7dUn1ePMsga
e8xPJtHjJyGy9mHAuzSzGfWNQPDFPViISyBiw6i6wxaCHg06r4tyNsqtOC9e+WI0
JoKd9+2K4vBxfupMtbD+Csgto0tnfEZHiW7ZvQQwMtDACYOel5TfIMb8HVN8JDyQ
Ugz7B6/fQcnJUmtoalBAVAdhM4h69Iw1GflXWkE4D506KfS8j9eE+u+Vhx8Q14fA
XZvyhk6juVs2xnyDepKP5AJG82UpZJTCeqYI8jmBz8qFcSaP3aIoSNINNs6M+DqC
fcr4O4dck9TMOS04MZM1RRCbn6MnU0tTd2HADfG+6ewoeQ95XRFfyaKxImy2lN39
o9ASBggyRq5FZ48/A9ll8QhQ3tSmdpapHhvC5DBuqWLriMRawleXMwy6SIJPRX9t
1UXHeJlV65ZxGMmNNnshYeMxFVTQLaIZWrB7VH9O5ybIoxYCzNhrNeZK4Jua3KCe
Q1zryg5K1B3tzqc7hJEs+kodiDMuucvS3P3yz90bS0AtJYdZzBRLqOKlbtxik8H7
N2FkX0SmQFPz4LgoOT4DR5dgP7vJ/wyhOA98s4ueT/Hb9FQACweocxsPQhevFATv
1V64Fc7YMnboiDGbY1nF5PneLd8GWe74v8vG64UBq/rwBUhdmPY6Rtfxy1Q+uAI4
veTH58C2npMRrQ6zWUn08K9YiP57CF6vQpe7YyhaP+mHg2p5DBwTLrmEwXa/M5FW
fE2H+gtyXXQnghG5TsLNDhd7KqjqeGoJDM+NdL88EHyvyg0UNmzgWydnE0b+19EJ
nU6qYCmOhycoYpSa3UH8c0baOZvLVPNAs9UsPEFh7nf7U1oxZpbQRKZ7Ej48OcyP
4Hdqo2X9rdLqAUPuVZScqXCEQ3ovC27qJex2pRLMcUN61mOukM34W0u0a0vF0HTz
Yg+GQtqowXRz90QAqbYsL+uW0eg+pnaZzcNaG7CfoWzFcB+5n6g+WIlxC/JOQPng
mgVEN7JCxJppizmkUUXbTnaeCUvj5Ko/V4cET2XVzP68Ow/cwejoBgafep9yaCSj
n5zHTxDhrJVBy2nlFenXUCSwjQJNZqbO4ixvYsB7g+M1+hfQhJgeVJKQG4EeZhNq
VcFRRqtfUVCPJiW/d2+9MoK1YyiG4EDAlOgvV9hxSl7+s1EggjQGmbrMaX92y3xm
awIV94LN1Pa46PfmQSvywJ2BxbmYXiDnLrpyxRoM73hOmf6VtxGM1on2PtTd26hX
8+qvByCZBVc25GTkGngqcJP59880328cFriQHgj7QgXK4Sn4C/qNWbWWWPWq0YFA
ACp1O8gCKc59oeuDOkT3NIIP7KsBB0wX3+TdvuDkm3vyfyrTa/uSIqoJc2gidJL6
IiHxuAqiPFLnxxYIK8KHRekWsqNqMnmTwNvLKp5RszUm3r8PKT79so/BmMTdEco0
5X5eQV9TotKwDd9BpowWBKpCL0W5V2Zup8S7Jbmv7ZKOayjOUjWiWBwJT8vOoxiK
CfT1Co/eVkKIWz7/SGubX+9zTqJd9rkSzAReCsDjXjiasBW7hYgkmjIHohpVAh61
y7cv7jzsSPClXuahH1iQlzyhJ6a5S2PwMd8d0edt+4Pu8j9Q274dv6lk7ZvGnjeB
o15kX75cfFqM8eLMmLv5uRvIFR+gv+glpk8lXG6ZRUvyOF29tilP+LZRlFgsCc/Y
0lLLYXhNMnNDqLDYQbI6BfjIvWhoUGS5BklG1QEUpSjk8J4z0F0zliKmqJLhdCtX
oyig/B/g0vjq1JPnfecnw3kKPTrpafLmjRK55UZ1uC21rVPgX7YSgC/lcjxIRhrs
O/Dp10P03VbB3rebTRx0Mn1X+8ogilV6gI7Rfn2Bagw0lAhAuNpt/CbHYNfWjgsn
gmRjNzt0m5e/eiS/acYU6qLCu9Ng5y5oxrKGd3MlhRT+5g6uv1QUj8ssYcuYLVND
nbMrP/ufdGT4mnWFppmaWpMZVRmbyX64Vmlis6szJMjZUwt9/cFrQeVMDPchYj0A
SJGv+AHoA0fwgSI3jv/xMN8TT986cDElA6k6s5bRHArd9D7wv24GDrwioiVBcaE4
8z78GGbGmLJbP/w1T4McV68CCnBQD4VHhO+pS14yYN1w3f20YncP8y6BmFQV0wfa
fhvX4hSEWF20TaoU63oykY3YusA3HWSLEuzA30JZRNZdAJOT1BDuky9yLFRCCMN+
/lSQYKzQbBa75lRrKYw+xZmcdzIb4XuSs6/5ZD9gJ5svCPvPacOe7AffYXxYDvhT
sl46PXJA3f7T+pHYSF66uOzHjscyEDs0rYTu+7EkrU2jnvMgjqAuPR/aVP9C3i2L
k6T8qhNmr0LEPQsxIzc0lMtu2ColqVN+wc/AewrQeyyGoEKx6b8lzBH+ORhAdMtW
i4KjmFowNseN71nDnjFVpOJTvYd1Pm13QjfhX4kZokdGjYOjuPifXyTwtbBB6VvD
sviiuIWMoljWrEibS06JsXq9a0RJt+CkRFu/UbEh0DnZLMrWjm6d7EOLZ3b5e0Mq
T6tuIJKypxqXxtJV07XLde8yOCabrzHz4ws9Kq9wS9phZq4xHQQDnodfAU8t1Hui
ePgbUF5hqjkWe4HmiUxmy1os7+YWytp1PL4u2KAo8eNJkiw/lFTmEvRiusTe3Nyl
R34sLxOKoskEboxfjSk7vVmzEacCGw3WVPvV+50cItgM/waNqVXgluRVDt7sfN6D
MmA1NtTCOL3WjEgCtw8lZumNzVFq7E3XoXSMnwdAIQB7tYipHYu9DfJTy9GHoHwd
Op5wMdwZjAI0HUj4qq5Neze0qmfGARLgZQSb27mEp9LZh6zbvFqU74ed5/h7Clih
U6zQhllpd/6zZ9ctTuP5T0NEcM/KSSwrteLVEbof1Liumk/NFWRFQ1Qfl+CYMwd9
trbjq+vNlZe3t4tFilyPFxES0y2M32K+np4ZIUZaNQEiFzlk06hsAtoLZG01H3Ro
q8/EqFO5Y8Mhn48dljS5W7LiPhzJb/rWgFKv52eeEooHQOIBARiDw3PNB/VD9duL
Qc3sU17nl2fzUsWEFLOdZaiFGFDXPlif9tdu4iBS0yK+vjXKmWGafPl562KgJ58r
sVSpYGcGYl9qoBa8uZkTxFX9GI4Jm79JWzsKV9zsa2BkD4NWoCMbJsZ2PnripGUC
yuZdEw4rcM9ni1zbL8EnHTk8cOayk7d9LVx5K9DESdA00adXcy9NrN8TUDyrxmEC
IJDPxo7NKIb+slK9I+bmPadi3LXhRFuS4zaak7yGSPyYgfeN3Qm7bIYBEl3w2MCT
5Dwo5j6jG2dtiSKZuwGnFkhOvS+a2dS+Wzf3oQ+0U77GhiZp37Xhvh0b6Ld6d02f
T4YI2CzQgstL4G7tJONrdU361yqmfIpfiFLFH4sq9L6yKanFbB+1xmU8sRW3XEDE
R4bAnFcy2nMX0r38gmqis3LWiHYqnpi4rkdbuHloNymbf6C60itgAIbTbr8f0oqW
AmgBvVX5Y901f3RYxlyRG8gIuOmKRDRlNTE10n30EH0HL96yhmVRxlV7UtqyTvWU
GjadVJrvpYl9ERlZLJ9EuxSvk12cXnrLPlJFFeQvixYgky0ra3ez0vwX+XJ3k/8s
xlijgTiDtunejj2LYPBS4GGM03v5XC+rlEv9TmLnLrX4x8uYyrrQ/AI/BAANSXSA
R0PeZhUMKpYa1+ccW2K02iktAJZjAxC4k84BOLu4EuapDIUdDj4kcMv5wfansexz
F9Le0KRfASQOBkULHjy4pVwFW5Z+Ad22LiqOjU0bpVj7Gyx/X1WfpZ82rp62dGJZ
Pg+xWdgsPPZBwCQEUWjs8+jCxuz19lKPqryQtN653loCsD6mpHj9yZXPYP+Pv0Ft
WJDBqwG/sjPn8vnQpY+4PNqCsJurJeZyHNiyhDWycOfMn0rCd75uvtGdrxR3EP8i
lyKxTJGCWnYB15eU9eY9Qz3rNxBbYf/aSrm5YQV1vNRGoBMNYDISlN968cy6PMjL
fkdp4aDrrb2NdzXFGqQlubHWj/+NKGurs2UHVXAakg20OnvPnqAphthDvrGxxKaY
7FQkwHkKcfMJy+CGjJXEGwdOrljnH0baMsYuZol1KqhXqK7ry4nzh1GlBkzLuO5P
hjhDLgIzFgsVDX+U0/aQxTPAOtJ60XLyqbm5mxah/ZyibpfMnYYNsjvISOi7HL9c
jvyRML4QXVsprayojlu1hVYFfOd2KismeewXzdrVMw7K4ZE3s9mtvQLkNFsF0P6F
2OXyW1qBeC3YOlxmXQ8D1GnHzTHshgkLa2Eg7pd1rvROMwlRdezk4BrsfZ8xKMOk
1ZCdhNTqRiioslwHJV3hTYKlGmPCanK6l0CGuNWg1P9jP1Z75pKYuR8Ieu8AvDL8
rqufXAyxpHlSY9T0tOHxi7W9D62PLXMRSq2Njd+BhtT+JbApXDYzsHjPxNWrPUXo
j/8UJxXZF+7kYPX2jF42Ae6jq/uQ6l3lDC0iJr3w9QvanC6RVwOtkEBXk40DhsDZ
3KtZegUxS8wlqStEVr3qB6huF0Yh92N1IaXKTo1wn8jrn471hSNSQhD4j0DtHwmQ
zuzJALAnlXHdPWzE7r0BPTKkgiywDeodAnOTGkU4MYV/LjCs+Obz3OVr2YNe1xnw
/46mMeviErPUI/RdrjUb4AkbCcD+EGAxB9gMsfy4QPKcJ23nfDyAtw06Tz4tSl3G
iG9yG+nXdjwnMqqQygInoX6vW81jcvXFH3XEzOTdS8GjdMsdS5tQ78QEv3HIzERR
cKQwB/pjVWB0gDFUUDnNbOvWHBvnRskulwdkCiLVz9IWfNwboN9xbXn/JsFtVnue
PILxF+ZMKqYvVvMuWqyMngDANztVN72PL2OzeLxOZ0or8mWCdi/4eL2ZkkrRIWoD
tld1fTY3MzyvEb63knJRlrntFF+0UdjWqcC8OgM0nT8mXYoxKRmWIRQkpxhI3nRH
6D2XebwyM9s19azCdzHRro6TIBqVaunieTLpD3EP1yMjja504/cvSE7Pt8lAPbAc
X1BWGYzSffP6gCGR+63rB08RH7pnPA8dyFiD69JIZFJSzBRt8v+1vW0SxUjRBrJW
UTNO7KgzimqDp7J4Hdqrg1CEq5NGfrIhy46/xUYREecU8eyjFn0+H3g6u5dMSBfO
zZUgPyG0MTJy8T52dqbJNVgbka3UAVVQGpraeGGE7fSSADmDwytjgaauxoAt5WKu
FFwbXSZJ2FMjmBM0V7hk1mZwgXshEFQD043GejoFPDTzY/yDOlVysgvULaynrpc0
AeOMqnr5nuvEodSbGs7auA7WODn3IKUQq4x1BQPbr0FCv98GPw4okt7N6X/ZtA5R
9cKEuNArikioOYw3oz15Rp4mGybTuQMd00IwGj+ujeKxn3SKhM21FFxZg7/7VkHq
whmvDzEJMNyY1y99Vwx3WBcyMTX8cHKjHBkwuElFGQDvmyaYW7w1jklKSgT8ZIo2
3yxpr0iOwyWPSSS1DlvCRHYRGzBXPoLypQy9xV76OT5sjMhN6SyQ8TwyHTli72Ya
c5vTggUOqRkENl3VsCM8aBX6jPsb8q96IHiT7/10Ohe1daqjoK764elTqNTY4Lop
uNR52xWbNrFAIij1ivi4/3zk2OtCbcJ5lFzqBRarTVR7Ge9q6ezHHLLApbPlaBYi
YujbbSf9fCtEIvL59/ArP/EnC648yHnMo7gEnb1HUf2vlv2sYGPPjmSqTH72Ahl3
sXQDWjyYJc9PErrKBSwEXy6CVuOm1nE2NOBtD3NF64OhTRO3nQJZ3bsbOQfXT342
ORfqZ3KUdn0C7J83kO05acoUpW7ILx40sc9Hre3XlphHXvZqCFT0ZxA+FIX5rCNB
VT5YLydoMrO3gX3Iyda4LYHNXaZYzcQdiiQkevMneU+/6V77Mp3WDX9rGAi7qm9P
aSa/7/G6eg1lE5EhDC3RorUC3MPJOwv8L4Fp2rhX7ZJfGDxi/ZP9KBiX126fQj1T
uYZPgBO7d5ty2ROpvLac8SiBONNhsNde3lBiwP1yOnBkZbVGIU4x0EKcCJbK5pxG
JutbK4f4Bc5laNcXGAgtxsRG/LPfVStCbGb81/Q/DqQV2c7bovkNhpfXbZFf13eL
Q0/M/PGaQ0XuomM85d8f8durjwU6B74PTQwo/7pePYfppLonKzJZzyvbAGNj6T8u
SpI0NekmFzoDIWGfZjnsx88WVF34cNb1Xq66V8BjULIf4f6FqmDRo43SY0k22Aq9
IGHXYRqdTh5EIc+QBWnJyMkWT5tAOdU+PAVeZGXhEIMSAw6Q50lXeEQUnYSGMVWo
BWzSC4BO2WJKdFVHhKSbjVSZtmm1RRZG1vj6BzPrELx5EB6n/2mSuROzObjdF2CM
7dIDuDP1vUJ9TDRRJviZa032NMhrgzQSnP23FdgJbtBrrG+oquOfngseclhCRcS+
iS8hCdrJI9qT/O9wwEynz/Do3+lYefGYvW+DFPiHM2JYafS1NJnXwQlE1N0UXrYM
I53etlZ9Wcrdr114tpp/uxvyThLuKFysdIDfA0LYdNyvNQYQXxY1sZz3zQQYmkFs
t+cfte2GfDRLhoOOJbdvM69VboSZ1Wv0BV1w9vnRr6fHfLWm6Yht+CBNOZZ3VZPu
RkIsZiBKpXGTzqvUMxCHnEGfmD6vlA0swk15Dut6ljuA3MUIOZ0befSuxoJsen9l
RiOgvHUj1OOhvOMC58n3glbUiql+zrJXiHGAFLvlNqypWpNsVHf9S5T4006pLhjT
8mAPT6G81Yg7HKoFTaoDcRrZfp0m/w6lmS+zwWAx1RzXh196xtC7LGRHNRDOx9Ia
672yyhN7UKnxdSzpbKJoIEenmf/bAD70dEBEXKvxpR+z6K/lDq4+dvrt4daRksms
RaZum/09G+py81EA2YEpJxjCrvy4zMr6XxviHLppEEVFLWFnqa2tZStXvE9riq7Q
FkQSm9vLMKGYerE7TKCRjYefResl0MnZRD/M7YI8WSe+70ZBHQ6aJPIQtN2F9img
prhQGw56La+ll0dx5jzh1R5ThC7TwoeL1QrZRDbE4FAslSeJuQounUjFCY0qhTHA
WLuEy4gH1tROW0ZwGVT9Nbv6QMD0BRsL4/+dBoCEwjDJSYq7p92D0gD5W2z7G5H1
H1Uukb5+gvcOaHf8nFPWY+RBb0VKcsNC4FwZYLmoFrDdI4dhU73kCz1AUlQAsD7R
vRzOPhDjtD17nWmMCh81wAaXS6u8EkOQDTVAy7Q4z0+PyD+Ff95CmrfaQDQm0axP
h2JgXXFDIOuSUSKwaL0lMLHCW4WZGuQdi56VGo3WyYjY9K9ddf/95pDBn9bJaE++
WUaX37oO2iKBJHZTatvri9kdjHfPn+vzxruKkZOSEMwxloW2YUwQKVZu6E9bUJL/
qaSGdUXh9hj5FFVqySc56ApL70xUcIVjrdqNxPbTf6GRkQ+bogGG827DVu4OgDBc
yCcMinYAaJ2Rk3TNSECWumt+qYBCjj0jLNVmALzuq6MTsxm1WQ5z/zwlij5Xylzv
TCKPvgcwCA3QPamLcwnOpVgJAg/NT2MRQWZA/87v9yRKP5nbbKhu+fy1FItFr5Bz
ojlXdTZc213jobFFSldIaQ+K6wG3+ZbwrMxJygecRkYeoxfv1HoF8MwecJSMtORU
wyZQ6nCqXHuVi1PrNobRuOs8Zw1N1bnixmTeOHO6D0ri1KQthoVe31ILs92qAwoj
CO20ZZEsgsB6gZJtn1te7WYQSwTkrB2rO3rDFO8i6xNoL7xeXunnXNuEDHtnAim9
l5yNCF5NVR+7APVRnWwffqR/Zso6zDYqnfwdpR0ZpZ68/BsvS3dD3QhkOJJ6TM0+
7/fqEzu1KcouuNAQ8RRgEfYxFVF3ZB0zgwUNLpchskt5SpZVCO4RUM+cWDhqJXXp
MuKlZV8Zc/yNoP7+CwL4DwG0pYkh1P1LI+2V8dZhfMohNZhoZWfdUJeJ2U4S7KaM
bIxj3d5HEZ0biRI0gfDTE/QueQBD58yr2egtw7uEa7SZW6NazD8iT9DkyfgiAkXY
zrIFXRM2YRScDbbRtmtXmv66jjgYVVsMghRsydcibeRDMSqATeFrDc7+5OEZztva
piCNhsqSGWm4C+JoNeNVrDYOPSwwkp14sjYGklfw4tCnSxbSx+Dgb2wOnkC8z1oY
Ie97L6PX/mqW5HU8GLtlQSEvJFsuOP9rvV8eEvZJriDt1iWvLH7iJbaDYS21DoRF
ISLK7295r6MSKNABsHtTE8UzofUslmH+Bg2jPHdrI0FHuM1SPLEGO5jGXCvd0iGd
raoA0U300Jp7lKfmYncCzX1PNWiGR/GMvcH1TyDjaM+tdnlNd3XBacq3XR0u+v+q
4iE/OXckeKD19g4GbDiyH7lxx1W7KpZI58RF+JuRuAmHJZRkaJAtaLn3Rjz0C1K2
1hX+Z4+IZnm6v0Yl8jPd5Qt3lVft4MdNmhAQ0jZafn2rqh7k3iYftf/+p32oIWXo
5PKb97Z4XFqibc+FzHRYmgskfBLkm/B/xxlOzQZoowtjUTfwqcJeEF91XSkSbyu7
JL+/Mft4Jd1hOMrzDrIIFMUbFYhNd3veIe5wzdoTiqQJhIcPu//J0fADy5UCgfsQ
PjyFT1POPwCZwpQ5B0iSiH75+JNMpi+UNZv4OKjyMRD5++VywMFRc+CZm3Wjhkd9
RKHVMLEOpGe5CnCJWdoeIo8UZYInVIeroahwqtRnef09scTyvNDe/iZUfzyAkXLa
aLr8LFiYeKMK0jHEQOjzV13YJ+5uFtF2yyvIFl/No7DNeMfHpWAhocmhF5ulpmRc
c24C+X62MV9594v6zwBpHvHfCCptPR5uY7pqAhsXj0k0HK/L3BmUgVzwLWBDJyFe
zbRmNLHMJnCCG+6Lbn1BtFFXCIAxoKGn+9BEAgJKDZk+McxuiIImf89ruquj0p7/
oiJkNPvRdnJaN7h+QLKa6/BxEAQ2gFxp0TLB05Oi0lFmtfk5hptGuE1mPwodS+n3
qlUsw1L/LX71Ml6WjWaiMpar7suILbWXJzHuA7Qj2xJXK3SbVQ9+0Ct2i45bs+bH
YBE+s2/c2y/7pIu+2WsOczCgfGg+v+Ip6EAZce1Fy54GLsmZdbQ70KsedzlGuDTG
lp0s2T/exMgHhkOvr14juFfJVRliFgKZz5iyDwsmo9MaL8BHy5giw75I/cpzFBsi
yoyLtdfm7PwoEBu0Qt9CPGaWTufY8q8qtCoGcdolvKD0HIHZ3jco89lU6Z5CdNpn
YZ3SM/KC2u+dsQE7K4plem8PBkD4QAEBD4SzDbga/gZ1YJ2ZNZ+S8RXPWVQt8kTo
QfK/2VU1GyqLUk/nm7Go39ryFNEd4X3myXqCxDnLvLqPondp8vwtKQ+PFn3GgVNw
qHpzmbdvLcv+E+0ht1d0qLu5qIvFI6DF4lmWzP419H60/Hp4RtZZbUmRrade0bS8
7tXPPIZOqE9NRwhTxxBx5Creuq6WTuRTlcvq55piAmQLA0YTKOcBHWhZDima+vFR
DyIKnJpWeGJSaDnzor78r/CN2pyNv1CLRQoW0OlHrSXLXr+exw+Ms76Ocd91W+ED
aSfXMeKbnUl3ztdecBExr/8djPy4OyC1YXgShi79WxnNmaC/KLPtJIysDdNhBh92
9tcK+d+7rUaAnsttaZ6ZdJaCy6up7x21idBaCmtyH4aYVMT2bRjbExnKavranqkS
izH2r1hQ84obtdQlhUSY9B+R894OC232e3FcXwYp1mXtop8Q9I6TNpVNAadL6RzD
/eU9c1GYmTv7s57zk603iczyaxewIo2TdVDjdi0kTIQ/HXe1OJ1dMTBYuj26BRaP
y7wilZIySStZoXZj1XprAsd5vWiUDpkePYlEwWLrrD9FAQl8TES+22FRcRu9Fhnn
oiUuPR49s87PYvzvx3uBS9fZhS3+kzH1T5k76CN1hIbooh0kS+p0gBnzKfrvXu4D
eRbRVcjReaipDKrTZuiKZU9wP+3Qx/2DDdLTvNPxuWz7tEw9BIWWdztp8nYc7emd
qAPQ13nZ/4g84AKHEBrCqbHANh5962VUXt6jB8vy1tNtzlNYinpr6EpDqS+G1OSC
JIJqZB/pcA4Vv9nzcI0ZPJw8F+xSovU3tcDfoXf3BDGWrRzV/6a2y1FnApfE3H8M
L5dbCFjVshZulRBjkQgZ7Q0BFblZw3wDqgnZ1reXQIVoZWvfVHoEYAbpM40wXmIY
nxjYwqlbB0N5P31YAiZv2RA72G9s/mhistU/iSqDBUTt7EAvhJwaU1uUtWo/sq8f
9E+Lye5kl3nZ/mm7niO7Oii18eTyr4pZha9ue1t0Sv/hiE+mrmjogeApSRRlDnHG
zeaRuwClRWR3cqEtVGsbM9hFQQSBh/dhUej2l8eeG/pjJyBDr14GQPNiJDgu10DS
4lBnlCKDyUtCF3mqo1GrVtv6ckYjY5DoGYsJerQO4+GJl0Bagssvn+eP0PqhPJtR
vwp4RI3MMJKyJT2TxjSqljtrf2Q9O45v6gXHTc0qTK3xerUwz9nMrnbsshIv4GVG
jCOO23IRZLQO2Z6VPQoQPkOerw7pdZaeJU3BKquf3yX48Iwosep1DAE2MksyEG40
kGaXJ3HlUkZZUUIVgMqyaE3KnXmDaEeN7PP8WuVSNzo9X1BLxqQT6qN91nE+1gqE
8Zr+dvGWkl/U0qfY1apbr1RlTz1Df9KrigrI3ayZxxjulTIkdyxfC7HfW5slB4yj
ZwbJAYtQfVsesuv+qwvQSYb3kU24ZTuQEfR2ATf5DPx73sTel8A4QLv/q9kasUEg
k5gtPyUT1NnJm6YSWJ6fe0U7Byg7BjwmxCOcydcKWENCUXubH0vkc1m6J6UmODVH
oSCZYkoI7f/Hd96z05y1qeiF3CSCsRiVpQfAO2mZIIxWRDau1XXi+Gff29WjWdFL
qixhn/gy0X5MRFnNw58pFISlUR9s/bvt4eq+DBjvvTcuVx91nev4o6GHK3+9To89
fCqYQChNX35scrW00ZTLsWdGBuN/Z0bbPnTqdn8fw/8chn3ZcH5gmsyCpmFDlPCj
WPyih6xGIbqfJ5J4Ai4TFBxb5/0qCCi/m+YDRSuS1KlFp7tN43UlGDZRbZwHBNRw
+OmVDGrjNB2PlOtKuof4t96YMGdvyMB+Klw0VB4ubwX1cwRjFB+uBmR2F/+LyOXl
nKbkJlZgrkhhRKredoPXHq7pSVW2YGum5I4kXZYJ4/nU5lLRt/OmMF7DlO9N4dgr
DAjWkBDR8mBCYK13CVFwgrEfbvNUBtK3I/jhc22XAWviDfG+vL5Re21APSPI9cgF
97kOMfOyXoxWvnrJPBbbvQoPTssv6YUnve7iqNE0Q3Dv28yVnOot8ueYOsoPW42R
ZHS/bnoJc/fZ05CVWwJBDeQiamgYiGgBBD1KD2h2sIDCsu6n/4QhmGlBe+R8La59
ACcsHSvSoo9Z9qrxvo3NdFtQMYnwAVvf0fnzc3cXVR8uTck6XH/5KvyyyDpzCjXU
E8qHD0XBIq69qGT2505yNoaVj8PE2Us2eOBfO3zPTT+DIk6qiNCjMgDnsq2XyFNJ
JIPpwklBX0o6aMeT2Y1VuLzAp7G+c96bVxGANlNvxSX5QxkOq+NuwJQdt1+hAdEe
aZi2BnilExjBj8rzfmQo8a83XAx8zR0kv1ana3SErQu2GZ5nmsJkGdly2MsT2JxH
qzxK7NQtdVPks5mKuHvF7I59CGUD2rC8UyJ+xNh78kurWp3Fnf1CHpzr/OhzANVn
0M+cBm69LnOubQhPmEQPJGPG0F+NAYOKgg67oY3oxUbgKq+8o6xguYjop1X0tf0w
qWpm1vbDq0p8/Y5BtaVYMGIYeTYr6W2qBzbg3nNH9GiD9fN6iuEl9fNLD3ElDsNz
irQsT4NTIOZb+LERXUULUdQ6Ya4ERtV9tUMj+ART7q6rFyFBdiDSWEUEAI0y7uFF
Dx9QCRfs2a8OiT0+ZA8rn16l+Gn7XKvpu8xC8/y7mDws3gvGghbV86U4IZTAVM1l
8s+8zXejbMsp0Nr26cKy8H5Gq34LoBtBiDvLzKoIHA00nez3KM86yULgZ1NY/Aya
sqpcN+9s11g68RDr08uh9tYw7treRx+18gaTDl12AetYQxvhRrd2ocLHiBXmMWcg
U8cb/IpvbprTFJtyy59sXLnjynmAqNv1VN+YRrOQcJ0PQW8gob658xxJKamsoDWI
VJQXlbaGO0VLs5k7gkBvhGV668C8XcLo+8WuY/TsxteH40BdJt+Jq5MYfEMMRC+Q
Nz1Rd7viZkMxAwCpV2o2rTk7M1ofMPu1DoO/oMUbB4+uDn/7MJiQ2hKLShc+NfQk
phnQLK6EWrP9+ZOF/STJikLPlu75r01g10DDe9pwQU+hvP7PRybekLEASfgeDWuY
wYkqkvwB+AN6xxH+cm3BN4lS0T4+cISIaSaF4mmzf8EJStPUj+xddgL8dvdPZ6AS
c0zvBnQC7tOhbDWhs4z7EQ/jEQVv6l7+ymhKrhvVEncU1jCuQoAj6b90P+HKZk8t
yJUFX6XPbtSZ8xLy9sgEUK52zz/kCIa8dVL5PS8O7P3sIGrGhECG/5e5qW6AInjn
mrFPBqDf8y/Ybnvd17FojUvEE6u2xBXHVJNRBSiEaooUlFViktqdqotQDSwaWd8p
tpoWg4hPH9pVL1+viU9w9sdQZqfAmhyMkm9S1uyDuAeQQX0lA7oGQdxyFEYvC3v7
n1VsxMFXdpFp24TSkz3QJrhR5qAT7CnvhBp9kHQu9QTPPu5YxgqmZvinHmt/YBSB
Z8vsixB01TKvO8p1HIDE6w//BnNvUJECvUZXpGJQish2YOc9ITprfe0oa6b3DIRn
AVbhz8qLfzscPkl6+waFIfR4a4mycrNMrfZXeCw844vA6XI1fyt5hgl3QDnqr7J/
jNDhjsSvUjc3XWeczq5IgfH6pYrmUK6KnrUtb44J7QZvMCYp38h3addc/qQ1AiGD
P+X+CQhbjmuRZK4TFk0Y1syGgA0vUlCsBrtpaOXnSWOxVvH05eLkaAdxfmKm3S/5
xD+/TkqdVXT/D17CinSRlNd/OX/j7vRWSa75lMIATevTYag1KOSSuyG0ga3oBNcD
VY3HC0h/mXWm/2zWtjfro6CpRj1gtaHDIuqAR/KxFx0mRQzMP+oGi2MX0bJu66bq
7Jpnw+zn6NXOKGjhJO4IQYm6SgQX5KmNYYnlCRUWBC+hbEwZa+uNFC3IK8L6+ICR
6A0Mod7Uk2AAu2NTJrrtFr3BHinDdyyvV3iFhTw9Q9U4fz5ZCbnmiyV2j3I1Eilg
XLx4QvZttQXUqKyVM4mBu3UQ84ITPAABu6PVm3LnGOW2dBxE1FfGa6QNWRkXlFgp
KktP/U0HmmhvMbL2aibRuCXFWkF+0GCov5mgiKGxn585eSHLw/ow8AbxPGZHgopW
4d/CPy74hpDJ7XMT/LpOOUQWf8tPDfjLmFZMYwtB1nZLKTODVZkfAvfcD6FmJD4F
zTNKkm40XLzfkgMZ+JsII0p121XTiM7HDNPLHwJrPZ+sw5jKcsHNdqEUx8UiIlnd
T7AfqBLGJbMxzw/oNhopekAVcRaAlPOaZ8Msia9JlmffU5SNA9jPmYX0p+L9wmDx
YQKccSsOfRvCuYVzNoTL9wOT8rOH65a/39MzShr2aQoEihHm7ZZMCX1wxToZSycL
8unosWJj03dAOIATHUqBFuZZjIwFTRLB02/TCLyexIh18C5yH1ZhCDPkw7T9O5JK
zIAbLb/FdHUVJAgxHF2D6rl+M6qjHPmKLZ8ESovxXkqDRBa8zdHL7HYWsL9CxnHd
xl2XscisHdyudWNH0SVgKsxIph3F10hc/HxjxjKyeeSR6UfGLk0uOz+20wMhPriG
rtTEZ8ODpV8zAxiuX1a9vy2jVzHoRMlYwINkJL8RC2mRS4ZbZ+/yh8hFOPXQP4RK
NwzNr3dzYFQDlVlNKY5B3KTBxBNVyuER156cnNKgawZo0/XkDPz3orK4KwACiq6Z
FSZcvpGXbPL7xzpiOVjJTw51uEFWQkF+oLJ9l+mnzeameqrfWuQ9jr7IFmwML0S7
jedYUQwwJoI5BCPZJ/DT8PX0YeQeSQVTQOJVfoOUcffvo/LRKLTXEVz8gUZYoYQT
lPik6P62mgoP/L8P6HtjvleGrLECdTXCEIYmqNUiuqxthj4bD/MR6hcHsxfC18ga
v+YmpbOMmreNf8krUVYi1OYFkvZQTXWS4eeKtQF0rS7hsd7Zes2FekA0BlDlQyc5
vwR/45lPcKPy6fJ5Y9EA9rrE6KsAfT6ieVVoTkUDCHU5Uk58F1XCY6aCKh7Ysxu9
8+XfKtjirFZXyAPb5LZ4ZVDO7ezmD0QX3p3UgtMoXpPcF0E3nHHOAwXYMBQzXCQ9
RxPkq9ejlCIYHJ/V+NWFZtOD0eHFJu0FvAbsF0zY9Z46ie/9tewqzhBgneuut30X
B+Yrxw/88BRi6wJcvNuS24wkJKK+LS+JbdAd6YHpVJ5g3bSDj5C/gv5xkC3WRLFY
CAKuhObwcaiHk3+v9cfsvauP4HXjQbd5iLdiXzZ8DwDVR52HpCJ75EQO3J0B7iJ4
LXax7aPIjqGU6gIS+oWbsbcbFrBn2zHjV80+ZWHjPULhs0UcqyNe8muZqsWXQlt8
BCUCmEbpSf/HxiVkNUmiZOAgxoUwLV1Expd6k6tI2x5kS0RDaMAMSSaYObOvhQ7s
KHI9C9AvDgHG8pXv4QN0r3rGdtGW3dIZWSiSSTRN/fsbpnz39pNSTHE1qftr01Tn
Aj+FyrPm7hs4Zs+OtLFPavRkIwexl6H6nmIz9irDogG1oQMXUyJid76JzQ+5USDL
TdKTJxc1gZlHVrqx6P9KvJO4dFse7vVcLdk0HXTg+aOfXd4lopQA3GapRPThfuHC
LjPegvDRTM78g+kJ8fC3lIZK5kOu5osYU+kXAHbJsdJl4jDwnHWgEqJav75OKR6r
SCNx74V1aQOxNs7chcFZdB3PCXIrF2wMUEADxUwJHeEZ6P2zazXe1LoX3cAjBx/V
UwcAaoHVw1HUCMroUR01h5WfvM6tOnpEHhyvREAavxVO00XUijkLoYMc9Dyo9mPv
t/OEvzzwSYunKoqorex8bX021vyJj541gcq4IjIQUopX4yYJlExbv9e2bV37CEDs
/vfo3VZ6APFJ29WvF2uQ45Dnucx4b5D1a9BRJJOzbehVcTe/p8Eigt+FRthuQUSv
Sj9X/yzTPHuRYDLNPFMq31BXgZqrsLNToNvbR7lWxSyGB5RUYbbw1isRG6oIS+Ay
JodN3W1N4bgkOcuWJ9HE11OPT/gpiJVZvItzOoROpJM9/vZv9AkbU0Cq2A0HRV2l
WVROSRq+hrmb/yt2rGjTip1k4lRO+PUaDUEUcmITy6qHzwX6gNzPmQhjhUzx84IB
psuBLm6yfgrw2NCtjXdbsyVQWVS7nP2BkCEr/BEKI0i5VJJJnv/tjmxX/wr+fLPd
9ga6H0JCWPknp/qdhpHP5T8rolEynBLnb3ckSVFm1EYvn6C572q6xIlwHbQqKbij
DPmTYscUSPCbFdlN3ssNYp2f5a94r9EIeCfMbR64OXVzI4nvGq7bK4vOvJo6dgS7
w42bQsbjUqmbOimz6v+yd7z87Du5hM42uWWDq0Ib6E4lLYvC1Ze4ha+R8UhQzetu
NHtlnFqCZrX5IrDTmLDORfY+WOpuGlvXVW7EHZ0BxOdteBJhME/7uV8OM83Yyn3X
7+lxXrgUFNpK2Xv5Nnqj879N19dbvLEwMLamqPNVeU3l8zs6Td80UwU1ZXVXx1DB
Cr/39Aga8LdCz63wyKQimjHTJ7CqMGIzy29GPZcgTqxSlb3A5N/WtbFvIPnDnnpE
hTVPooun8w87sobMgEpd+pLn7xjFXkG3Rv4LfzxhuqBAhYGGHB4Ed4rszzPFN9eh
a2TP39xNk8yjwBGDgbvkC1CZ+GG/hKPTAPsjPlOHbcXiPWMgt3UhZouWLlIqHoEd
AFNYvy8A2WK6hYxFyMZC8n1KTE6LZjuj5oUEg1mGMt46s9tZdcQspjilW977muu3
6dz3/fq77oLXIjKC9vFGR1Hr6CN2zjSxv8hbxp1BcymJW49TULU8FOVP8iIYaUoF
3YCMCBpXlFukec3p8lH2ngfdP5uW/RfdObGhObY6IyTMUMgXcSgguqNW+sT798+Y
3se1MJIpiSiIhQY2XqQep/UaJuQBOlAN5T0nqTzGkZ5eRy2ldER/595epLN1WJfk
x9bHieDqOrRsUgpTmL1TZzdpgF+rTG5Zrgy4ky8otrAQ5dk0ZO7QFN956BxqtPEH
Wth6QZy3H0rjgOA53vFtqt08Ish4h0+BspijJtG+p+zdkR/5+v8ciOEsLb8fhyMW
sOMNRRc9CZef01geuymxhvt3HQmlL55Nyk3qsx5baJ5IVNljBSb91cSlj+UISYdD
dydZDEG2lm1ghrznffMjKGA6Rop7HaMuIuYCFr8hH2d3cf5fRhsoQKTmRzzeOr10
fDfcEvCiPVgwPD6OK6EazRNyto/yokrX0Nb1x3TN0OiHP382HdYfh/VqvUvmt/Dp
Aqxmae4KK78uBl78/bkl1Y8Zl3SNqJsQ9TOnp+w+09TneqaEr0oNHLvevR21IMqu
FQCg8gUXW8AGTbATnK4t1Did/i7envuV3sB6A2sELBlTBdPh6EFKY3GmvaM0Vjs3
vjxJ2Ow1PsgiSwmIh2C6fV5llL5R+PTzpS0QN8BB6ztBzOxy1LZo0WnknwxhxiH2
7IJtMxzszoBD1fhVg2lv8m2oj/0Gc/tupOKDGNZ70VrpybFwXg0SRn6hIuARC7OV
o/JYIw87XLt1xuInBT3sXZScaK4JgJEm563r0TKIU76Yxy7kf1P8YPU/m29a+L/y
GvtQmXz+1aKhE1s9G+WXnU22VaRXhFm8YwFJf3DU/HFzT4J0ajxeY3XP0+REM9zD
6rtq874UXB7SKMaTjMLU+EyDQdLpDyTGk27n9KShWW3c5qD/sQGmJ2j6cB7z8WKv
wdOvpU1SealwukrRBnHrp4GSDI0ijQfE6xmnkFZLFoqwo/u7ftH6AAZOVLKtnBtj
BngPnOPkGv4/IorO0deFGmAY1N4Q7uc4F2TP1q26HL4Glsa0HNsadxrR1gu20kQI
bRfFNGXkqu3WthmWCo/BPQYgzQay6MQm23hQkK+4RU8vvU631/kPFDnR5uTtV/5e
A9hpdJo1PbU5bmnZ5/IKfUFwKaWCjQcfZqnP3yB71O1qtl6QSbXwCnH83ugQ2V1s
V9OxkXpA5P76bbhe9++/qBidg9jI8rpbPbKMUoDv+SEYrlGk19kMlPAP8tkXMOP+
yyk7ek5QfWUCLHN1rixF9UdkMIgf1bsbaBu3dtAUIs2C4mgAw9JBpWkvtZ6lY60q
lYcZYKu/FV6pCszf/yJpGO86b5i20WHRjsEnC5v4skdBqgv/dQ2LCuPgg/ir3LLf
IofYvEKCKpQEw/20eV63+iijZmg9a6Y4NpIv82m7hcHUGv3BmBSkHYw2hKqtl02K
n2GPuOH+JUnBqnmJD8KsQ3nyu9oqObWf9RWE3Wb96qGimTy68OuufEfemmdB3hDm
6knp++/2tEimd7zd14to+zheQkZBpWpZ98rVjX7eP49CrZ69XswDbPoYfJ5ZMa0d
kM7yDSGaOhPhBQAA1o/bPshJA3tMB47N4bEKj0rImdDmB/a3DAz8z78Ag5WAGWqI
nl0x4W1KbPqL36udTMUT3BzDItWBGcUYPgYiFVxL83l1Elhbe2uW1pUC2a+BlEHT
QX7VOoxpGlgYItoPWtvjcBljlaSqp+OpUUGIPrPjbcMoXkMdCFxX6BnhRAQVZO30
SBmSUw+/eOHtNQnC9FvbmbEY3fqbB2ziPNrb+DE9WwnlJ8cY99UeHO2ioFEFdCBm
BK81XRKOPylZ5xGbfzwOwn17JV/0dHMWeTa+jcjtcOnW09Qs72ETguXdI6y5tagU
qeFsTN2YfsVz3kGzMSU9RHExLbJQghOkaURme4nwcnlBLho4COUs7217d8GPPHPQ
yGCGttJ6/N7I1Vkso/nL5J/s1/NKJIesBuPXhX2pT8aohWJgd7qJuVZadPXQRkIa
yGN2x3anQFNTx+iqBosLr7ww0qnpxDQN0M2cceUmS33p1IAZkCnTSMBFzQ9b4GHy
0eoO1V9j3QJCHxBFF5FTn+e499pRUnTRWaSyZIxUq1beYZZxlX+fyYzlTz/beVIW
BfHRfVQxCDpaQzzHT28AQVSPOtfpYAZnXewONPnO23KJvUBX2ssZxlLiUieSZAVX
OHjzmG0a6zCikPyXnV30lSYghaOGMjkgAbcwBf73bJ4iGFNe/64AYVpVaAqT3dqn
0Bg7WC5IFFYnLMVCoFr0LNq6LifpjTE91g5B4dP1GRNK61XvupySFF+sRewbwAsP
rnrT91XSm8yuT9Q5kPKv4RpX6uFBzx4hupjUIm30o2ajBhZZk3RRnDRqw9NOqpbc
tXaCXLChDezzbXgg3xvjcCrYpfZ7ZFL1sBSA9JaA6sRHQJUm067j+UTTAJSqLE/u
mBHhKLblXpzh1aHvo1/S3r6MoU4alS7FsdPb3yyErkuj+4Ik3VMX8HH5x7e2qCsc
w33zUeZZYUQtVg5leizF3WMefUDROdyreilD8TFvsFq0QU5JIaJk13HmYO+wg8Xc
socCTMgy7hl7TQjlB1fapIxHvnrcfDPQG1RESZ/KV+ispeYS9wuflKeioPk63ZI2
UwnuR/ga3Slx91YyjXtnWiytGlxCneW7HF0R9BvU70qr0Sx6FxpEBgJJbZJhme7a
CuzQwD+mCZB16V2OZ2PqLHj45J9rGU2g2d0r2j4XviX7+RxQEQ/rCVVxEOyfpCNV
DEmIkhGxujsJfEQeXc5VYgL9QbgnfO4x3JUow2ZJtnAitpZF1Bzv5gerDPv9HxYB
lXLe4v1QY6BtvxOSzzuIng0mtA0zbPDpmuVrMXsx0TL0YGk+zXSmeH3H6dux7BKo
A1zG3pgFjPOXHjbISYRRSUXe+jKjVCX8ajGU+SAPcVCW6UaNNjyU2eQFJVtG6dDw
uqch5ny9gVqUnZxYx8pg6drX0PYwt8RUWLQJFtmozbG1iOXWGJiznI6H9s2nW4mn
qIMCkT01G1TgHdfKv3RP1+oPkQkHyBdJTmea68PTOH65RTiCop8Bjz6o1nbela15
5ghXRz+9TvIhmjqAkSY3uOyDkJxwGFvYtGCykm1jmFTN839vVY5Gv1udDK6CNMzX
bq9Ydud3ZTSiLjdm2PbkO78TQ051Cwlh9pCzzG5p+U5Zq8ROinDOVNK2aqh57Dnk
PsVqfiRi1zR28MJG0wQ5t5WKRdVeUJBmKgpkxJniddZB3sti3rgkHstbNaMD4Nzr
qhSnrgGCpBAGb0uWB54fZ4PvXd0XgUtKRcbPK2SXLgauy3oCkYjRlFScoxWo2cGx
yxadcf74ADGsi1MebHOBy/RpIw2B3JhaNk5SoekMbwJl9ajnmNivx3T0xC3YaK6N
N0Px1MgPdBJZ+k0XiIPNBVeWgJ48shGQLepUK63Kh8ZKs7yKMcwtz1wJ+stKXtAZ
IvF1fvBRBuL9o4aPObbQRWadg6UbwilOsbgJQFPhm1T1W3FDM+cz6eZPBB1/8DcT
y3WOE2HRurOp/bprXXDNerlWDERs0QnSA7TyR/OCA0J5MfPsSWfF/yMi0KFPEPMo
GxVYd80skAtyTa0A3GtkSzu4KT3mzj7I04lkO0UP2dbEDuqA1C/bJMQEmFeIRreb
HPygpeJPxC+OxUNLlzLt7bqvg4XrHZUuG19BeZe7FrvyhjDnxpN1bYdQEO14BiYO
l4cXBUpjxZ2M+56zRdUm4/RtDy4fztb4HySKQYJYnC+jaMUN/Y7cAIngExoJnJ7w
xoCxN82+oa++rfAd9CPS6DqnOxLYHS36a74NFr+qw2XH1Yz1JUOjymDUdJrAYp7d
w0uc3cdvZYUYPlKyrHRZvLlR6mzyFrJobGmessIE1xtl/oxeDcl94kxl8hvuf6kC
cJKoKQVzH4W5USaIiefIFVsZaMEyVPUfDr7zH9jPFJbFJKgKA3aV0FJOQELSFXhs
GzvrjRJUzcU6D1j8yTFfkAeCgxZlrE50s2p1Y/04T5xsuAQ2KLO+wDhAkEto1nRV
3jHawgWwXo4d7kxDCka1RRM/WSgSAUfiKUPozCpdJToEhG0g+eGVQ2ZgN3auONoM
uKyMUbd4QUJw6ZjfyOJwhHDaUcnn4j3ChCCEcp/mDaPbQiQwQZ57FNw9ylujiXc6
43iGhGLcN6z7FOUBujwd2Vri6vjMk9XeF3LorW3PwAQ8MY4sZkIQJKzivCVGtMxh
QRyxotWtarkHbQOhs+B6vvPYs2PiYuDIjjpRK8qgFA7mN54OrPptUtB3jKWc9gmr
jjmpPsbDWgg/iQkwGUCikp9ekA9PRLi/BsZANTxVkEiW1bbm2KhupC1rwZ1vNRuq
AZ5l8kaJjDfjTdqKCAYEiyRc0czcjJYE0OtWlKk8TAO+R+juGYtORpi1LTR2PAtv
uGCoc3A4VcP3USyZzYnv8Zm/xQcs4oQ1fkm29bu/uXmgxIJhK85ya2X6888mlKSh
sWM495Awu0rP10br171+oBr7QEcg9mblSfs7Nwk6jCwoBSAPnHwQgqI6ddbumrNy
9wQm4Yaet0ZpdXvS5j2BkJCOL+Xx/1VkMAaY1wvKlpXdAbT9o95JwkXH9EDqkrpO
zsoN2BfGKq231Ut+axDQFGmyxqKFY4Q9+H1geBmDjdUztKXbakql4jHRyniia5o5
r7CbKWkSgZ69KoqHj/CQw6LS368wVoZL77kNrM1Uvw4nxOeQxD0kqofIW3zHv8eZ
AjyUvXJvhemY4J83xaoL2U2ANuOmV+CmXNxUb4ruQXUVfVo1M+z3TBFsPk3Re61+
1Ng33NCFzdRJn2NuXhz39tcRmd8VOpBc0hbe6uLoQ+qTlj3Xo+ul6tMiGO5+dWzo
vpcppPIk9DJR524Vnl0dsJrn1Kc51ogA1X0zlhNq+f2dXZ5qNS0mNZQ5Pg+YJshd
4k2dAUZVQjzg5mm7H4BsLuTa9JE3ePsEG6MEEE3tghGIjRDBNNvNz4LYKBgiugM8
Kcwifm8wNT1yHEDKBvZPHjqCE7XNZoTfclgXpNG0pjwSrteEyxl8aAxbW0DcTP0q
V+sn+BRFdPx6dUfaekxvsyRMHv99z4Raorojr8C93VxJe2bubMOsSNcyhKT6zJHR
cZFO4zpTdyFePUrQ5jLwqBVSzV8yvRAV7hBqpCyOCOUABb3UfPUhfy/7WZKOA7/S
bqMK3o4mjXnHXOiBb3Ls9xIMfHdphkq3Yyb2DM05celp7UJD7QoxTp1gfpbFKoAW
MIWqWdvqvSYOWaBMzV0lF2yPeBJEP9BwAfNvekgRVZCiiR6K32QTMJHjn9peiBwd
a6QDaGxeSBHht0D4uyZ4YZLXHFoGDI9OXXcQTsrK3l3EfinlkB2Dzsg2zyeViJxM
cuzvtJUrXUCnVJo2168J6rL+WCo3KIfCQf8MhokN1ni+pVuo3A4StnE6iWWNbyTK
nICO28+lq1RPsru2SbGLhtcgjUgoVgoqHP05iIB+lRbpQzi2lBx3POjXJv9lhloH
L2VSn6ACVb7du+iAjrl0f7+SnHmwYD7RQVBcjEfe10w7NDBf4SCBQ/eynUZZ1H4v
q0sEOLrhTs2uRx5LoitfPudRobHEY3PF/rmGRIdGXG+5zGPtQ5hbHquCditqQ0Bj
P0llDhWwl3FnnNlGrIlckILFU/YWOC/PZ/hpZd70F1mRLXaLiRnN+ivsZm0LA2Oh
Uz5ZKNH5+KrBcnv00z7aK6KkYRSjKWWn4R4CtZEQ5uGWVVVIxyXaXPX65DMhZ7a9
0JH2lW3wJxP6ENdNkw6H6h7uCricni05fXk/tGr0QDqOnIF+HkjmfpXnR/3T/TkQ
e3ZAzuqpRhtQX0l75HguqMeCTaPXlPyMaM/u6UxC3sMJGcVC9il09PYcMdzuYAcR
k1NcCWmSkAcUmczn3Hyw+KycJ3416dUXcKTmdes1xKiXf79XjwLzDnUKSxr47uLo
YWu/ivEZHohpQfbBm3lo9oBVr6JLrtgiKZJ3F9+NBd9XBtV9ydoro+kwbAxnWB50
AlrLjVLSo/5RZ9hiKMksCGDksuEsqI6vN4xmpjUat1zm1zUSkd9xeIkYa2VzKBdf
Y90cLLbWk/hmS9nFxqkeL5wWDwNjeJw75EgoxzqFh7NkVOj8DhT4RN+XwyPlNj0f
isoTXER5KoWdjsUQC+dv5Jw52hLOx70+cenQe30HILO8xD+s+W+naEKB5rdlILSv
n3Dac6rseLVDjtFb25v7gLEso5dG2kjTAjtyKIg689WoWWbsIiWWw8WgKwuLY4L/
RNIBMWv4hFk8sThYxCVcv27ZrIPb6u3MVWuj/6T39Yijq3TFt+uqvtbMfnXghnsg
VgZ6ZKeHflI86PeblDcXrFmk9RKiCWfAl0IyOM5lxaerzNfcM0njwmQloCunyFIj
xvvrJbwx9y60VX7HnZq1kDjI3hXtso/2OInADgGqcxRa6cRrb0n6sioKV6+EdhWw
co7IreDV8+6Aln8HL3MVG9RePduuYzL7cYsnbRS0ZnPelZhEN9zZ3PEKVvNajiRk
l1vpPQYeVPy/0av+FwQPB0l9gMLmyb+5Vzc0J3vg3YbhWT/jS/Y5ivVcC/ibtDqO
2ajzaUDjs7hGhjfEPaWaVyJDFs9TjUzHvw+EVizk5jjLAlxSALrpByPICFBcRtFX
zmt1hBO+Uo2UVjksamhIT0pEz9aWey3wH5r1tZz3xPYaQL1rlvgwk01P8LuefBu0
OKPtvCxtcjCSP2CKnTkgjSmpfmvMo1U/iD52s+EEO/uoBMOtFhWDMdAkPR5ZOw0a
Okz78O/BYAwzb2SivNtNr67Rmix/Xg6vm2/TtIgT9OwdRejbx6oPSK9xjxpktrgA
O5lZMA8r8X1/Bp7ryLH6OZ3EQy5x70QilBEEwxj1vqBJxhmYbbE0WmSNLLLpUKAk
nfwX0eq9auIHtmWQ0HUnxiTUXZi7khghtGoejpBqZG9HjyYsnX2rvz1mFJ6AUJsA
Y10em0+8ZBpXHlSk2LRu6/1rR7ifYt76hSyq7E6LXZDRbzW/fxlA/Rmr2ScID9NG
fOrVxtewaDJWBVw/P93YnZXQPvtL8MZZA8xoVFEEWO7/jaQvo7eZz6aV7pDWNiBB
4kRTxDmsXqJjkhWAumndWoaLK7xpH5djUI10624fmb227b0yRRr62IF3eRP5EDnU
PbWmYy8iqJSGxj7PgrkduYvXYHe71zDuGRJBv44DeuJHZMhxg4N/McucfKOHoYTF
PCSl3aQReY2h0GqqF2UsO3FKGHG3LfizvacJNZhSh9f+mTFC0gZMKdhcEshQqAtt
s6mx86pFGFE/90XV0fx0z/iuPv97qjucn60dPimjXFgsgZ3ZrVc51xNJRUaTa1Mt
d4Ihez5wsZYz9kLrEVQuOseyVa8HNs0KWz+tWNPP81LibIWJGmZeILFnECz2Z8mB
8ag2yaOEA7yiu2OaSejpGwtG4ZS/OqnX+Yj/Z1Rny0QT7Bf8vDLJrU0eH/U1nOr8
0+q3gtuqQKFCwM1x8DY5wE4TpGQPUEihr6hW+ZxPQNhBwxWKz4zIAJMUl+/iYXAs
DVh7VGCGUnsA/0dZzU+ksdoRT5HSbYd6d9RCsSZ88XiCKZE1Fs1tFkwd+NSPTACU
8jOJjn9/GAEaqmt2cg5m5dyg/UL55q4WR8gfZnvR0YJ5TFrHIIROYYihYiMbvl8F
YmKjeg1Dq96i/3Yx0U81phggiLADWXPm17v7JDwSTFCTWGyjyqe1gLLjOs2QGl2U
wlOKEVrp76MTbtD7LIxlDDi89PDgHtJjMyCnlOD0GZn38alSH3X3RXPdVaaz/jjc
IRhk4HwuIF571L/NPmrko1qTbcl8LjSr/VAcrl5fT4MJsQhXaXbWNAIGAw/uIaUa
YhZaOSUxQ7n1IoFH8Ke+dnahgOLhd72CEW5qw06eNMCO7RB24ka4cL2TD3HDUVcX
roc7bbnbR6LaJFJY6V3WAV9IYEswuXzvEjnUAMcCmG7a6p5zO7j9WVUHqOE3Sq4j
GVt+YKR36i2sv2IReqO8PrlA7fcTuh8XZqwb2Ybn87qNe2cE/WMfHnT0wZ31QzDR
Jw4wyz1NXvh5XuqePCsnKcO8G8Er/5mdAOplTSjyaQNrBhNdXp9kU2WYSGlmZ5On
Il80fsNuAHNyQ6QwzLb3v8mxu5PN2SYPrGip9FKtO2xPiUBTte+FLrVmlPTeHH4Q
5G9z84W0gzyG7DzLhT6Nx+UjjJwMzTTdXIZ1fd/OOuHVtWjIsV1qUPtO7LR6BSAR
1qCOpJs9jKdMZy1YINEHiUZnJmYCtVhzet5cgg8WEIbTUIgSeOJkVWIHNUGo2LR1
M7MuVtXM7s70TD9bJQdR95cFZmFwLmvXcYP4chJvayNRYdJUcYpoq1LxaPr0IzCF
RE/WjZZ8FeMvBypQEybqDHPkIW4Wok4Mg/ayFEITtq8dZWXQ5A2R15sjJmbbEneB
IbuVBZmf/jyPqMeAsSUM22lun3/mRjYRXN2bjvRO+5w8WhnkV6l9YDgBhFSWuvRy
u/QMDLXCLLAr98yQRiAkKtYQu/U7QpVZAsQ77/feSHI5+YCIWAhTpzf3F6nT1IUu
9QfWrPMI3479GZqtPXWuwwzgvgkj3OpPAJYmCSHvMTm5VGKwP6ZOFavNSdNQwoNK
lUqO4GoHeX15WXlF5ebLVhVRxy+qyH+6ZNabc0iqvpBrBva95l2FJ0gPaW9cI3j4
Z4hAZNrgHr3GMQDH41ye8RgwRZD47L+xMeOYZgu5kHs2fpK1Q2K5k0xaoEg63d9P
CNuQwIq9VcY61XHc6pT7cC9bPYwn206jB3hDnVmtpwc4WZ07Ms3dE6y/xYpH2Ssc
pd8fQ4FY/lb7ApYAa91WB/a52u5p2on+R4ZbvkiLDxKGnMzDrFe/GDnC7ouoqS+9
X+WoUcpOx+gTOeC82mPeqmYnlfrN9mslPe5Ujp7nxdOPoVUSJ5nmhneh3gVCIQSC
IK/PAtr/O/RT/0SOoY8HaWYHMvIHYbSHoiPYGOPkdgjN9l7ZUZTjg3sJKxbogcMe
SD/sYe8AO7fBU5csTLIDnsvB3MRpjXpI5NpRyWnBOk28CP5eI9HgTLTzn4tS7c1n
uISdkoPYbBJblqLb3R9YrNsksIAWPXiOYt5XJgcmco2EkeDCccowpU+leV4vmZ7Z
t56Hoq5RBNHlYlz+RllihGUHONtt3gqcULSVU1xTSyRdjfS+JesL5ebbT9TX44by
FOUWe0Yg3dZq5rfqp/Yb6oT9+3iPfGYwTjRNK3NTvM5SUf+LP7jYRpEQIJzin/nh
zvXBCkWERG3CbFGT0XKDHZBUXfzfBr/NuApoPbylpZDUEZldQPP7akQ0XWBexPbD
GehpFI8BB8sFJ5OiMpRfvlhKhoBiBGOygEvRMR1t2Fz2VGrf0ErrCxcyhV5DB+ZD
BoWC2emEW7t28Gg+gS+cSTcnUh3blT/NwqIRa+IQACuKdsONG5nJNiN0A90kEgAm
EMAIpcJroAnKcjm6T1J1ozvRiZ0S46gJK8viFI1CPW5EY4HHfkzO105irVuioFJH
9Z0y1ACo2YuJ/Q6glCksBenk3+wMKlnSo7RhSMCaUo9jdPRZmDxbmov5s44uayRJ
H6olrljEM3tlQSCOHncGZzA4hlYJ5Nejix2NtipjqQdrApvy0a3ShdpzcQIkE/aH
3MtaFyDYDlXnAyexjOD9kK+Ijwlqn98LyMq8POcRB1L8EkzsFCccMyEGi2r6w6hm
Vq1zpRDabpMTcErH0I8qri6Xxx6p/KkhGQoB1gm8XFhakPY9pAbyc4Ub3lSA5sa8
A1YoTZuvFh17/4mISzM/RXnDG4jIBYNAk513S7TZIDhSYtJZIg0TrcT7cdx4u4LX
/HWepKipRHhYD37dAho2IiFg9HeRnZrGzwNOhnn54B0SLJhTzj2bb4D8ba3xIksV
usmB0jvNzEbvF74A58hOLZG6j3dzX6hpwPIz8Uhr1iEB4Y7r0IDq/wJPl3SXnqaQ
7l8mytIkgKimAWMFDb49swWyovSzAbAVVl8IiafkvbzkwPw1QAdWY6M/3Fa8wKhg
C9GtKXAbLIonHut2gtlZvblsvaSv/tn6T5u5ejDMQNvgeps3tpbai9FeYXif2lv9
A1G4+Oo1qAi2d3pHbhmwqJLP0i9taclbGnVkkc8hJAnziMO3fNuF9j6t2VIgjbSz
CNv87Z/If0kSJ8mDmdPfm0FEitjbZYOVQC4zcH9bQtkC67khaZb93CI5yHhY5UL5
cu9MCT7+T+X9KCUbXCOWkq6MLn+z1n1duYnke5ZTNLhyMhTVpkPDcWS8TLnbK8b1
w+0ycBiYlxfV0WXXkIQ/iquZ+/ul86doZSwZE08O6Z35FUsRsAWvDHmV97NIsoDp
dDwXZUWfN5u4ZwG6OT559cOG4jiU58nWs3DW2/2iJUAtXqX+dQ/EK6ZHzrLVOj0Z
Vr5FOjD30xcxw4rIUN1agQJv4jdkCsEwfR4hkqcJImDW+lKwJBzEkN0OKiwbQPu3
PhRwh0VdOqKEobXAPMdBHUW15Zftfw0D2xDDJ9s/7VYD+cfQqJm8Qf+cwQ0Df9TQ
Fg9R3gKfurczuhLtr5c9AmH4XKf2P57m/Gzz2swJIkOdM0N8WhrxiWLKXJDhaA68
vUcvW6L0yLGrpr5ikSQIQJuTHhBOKggVdHdU0UehmxZEY0bgV7RWWFX83lbZQtqn
//EngmaNnD5YOFpEj5Hoi/Wlflj3TJXv0ObFkfeWD5/5CLdUmWdatFD+vMV59D+A
Eefr44pIyftyUjTPq8LdpnHoFHulwyHSmALZGflxIDNga2TtU31W/zAAjaGZ//AV
SBsHVi6mS4MP0v6DJLXDIr/a895UiWf3EBPJCZL2PB1IrDQzGQyOLVwAr5w9oq8e
31RYtNk4Is7ZJFeuhhWMeLOLDJyBmcpU8chESWlBjYPtbitoG04+CQq9nGkLEYs5
GtZdsORLjptuLI3SzL4yaiUxHTcmNHLmYuxwme/exhuAA5IGEHVyTKmvmOqvhLTA
gkZj/4/1vO5t3K9aiYENLrnrPWO2/hH4Xg0v01gZi5gwsfmt+iqooWx5HdYrlhp0
Kt9WLbXyh+26AxK5lPpiTtf3vwsQwgaWjR9dQrZ5L3aJ6CfiM+/mvRtWKBOlz1tA
STcHbjpFfnwiU+f9rUK1chqGa0THQsKMqXYeOYCB3z3Zw4C+HGIOHjpeWaSGCTzm
OO8V0v2FsRFKkz8aHgp+cnoOV+YyWn2PsPqjmCiuOcOI79a8lRAve8kZiqaJStwi
fLc9rudUpeDqs52Tg2aXDGM/jZvN33L0H0tgV+x8yonJvZVIc2UL+RTLf3So1xTv
KVeesKSN+KmfkKZLjIy+rVMXouz2hxWTbvb+2V20+ejBwEruEQ7b8EBI3PoBgQ34
LHHAmH0Uar5HeSYUWoyxONra+AOQY8ervrt3lQCwp4O9JXVsVTOb4ySkgIJCWJYT
2UclYPT6VHbbUkvPxrko1tIp0n2eP6Kd3iKDZv+BHH8pTQ/rxKTH4TllZBJLH9Gb
B7lzvwfbnZLI5MwWVSOOXSSyuaRWfMPXBzA0JXAE6slnslNh5zweS1kDuVlk4SUh
dOhs0ldR/Xxvw/Wa37rIAy4F0fRSOCJ/29XXBw0AjLHwPJk5hO6TkzXcBoPy0sag
xb8uqQXRsfkXgCj3mI7Qf4n58Rn+bl7oaD5QBaiPh/1skrQOCvFLZCeY2gLSmk6X
gMVv6pnOqjqb9i1X17/1zFVm/ebpUvO2+ZpLNdlAIY0MOTSezWYB04EsHkI9/NJm
/tkeD4xEjoFj1873TJYOdLhAK1KYSLN7IdxNYUojvxqIUsuvHrSmcmJes/hvilf8
EgOyYcgJOKjMClV3mRWbu+ifGmBdUvPo59XBv0g6Y0Cd4WbhvMKeupmx1I8w3jkJ
3jWG+IjKz7OR1BxQjCjqblTMUuWWkmpgnpGaI77+sRiCteREsCl3AoU2tFYaHtTv
mZDftF1838sOdLl+7BmcEdk3Adsklq4+qOi6k9CyOVmgyjvLlgA+alBKId+wIbTI
8mXIwZTPcP4Wes9DpqW7M0yU2utw9UrDlITIvplWMoXtjX5eTdNz1s5LfnUohPh6
EarHUusoTtMdTcZg+gztOXJCxx4+0+71v8P2QVTenBFIZcz0SDOXuXw3MctYt4mq
9x6DsQ5YkuTLCnMiEmFyRad56rfX4Pu560DqjEmR6nd65AbCn4AhZJw5H4Pilb/8
zL5EeJ27G9+JjFl3oWc1mtOD1VMZXRRhsNl1bXqdhVP3SGlNLix+qZIEhy8srq54
gT8PfG3qBoFXgRPnp+cmS2sZZ650u+GgArzpV2dQBwD9uJ9iTdb6r5HmWkuvkGjk
u+tZtzeDdgM3WR+KDwgM1QZRhidNIF3nCfd2zSCC68KdPnPLIrhs7nHD8+7gldTd
qH4/3m7LzUhDYn6EaDk82CcdOwB+mRPhXiBmMjbUJiDc3LQThwiVBJsGWg/yuXAd
46o9A0ERTtvXKe0Hfv88RbtYQ+XNlGaxORj6L5Ob+claa1lzlGBsb45ERFphaEmc
SG1FXbSvt5KKItKGBvcZ/Q2S/1BBAZCNzey0WQohh1Np/+FMtj4wG8FIbsKCChhx
Ulc4Hr9XctF/Q2GnE+gQj3RBPGe0/t4crKdt4zVqzGJPfaISQsMBMiLQdIn+ddsP
H1dgLjgBtTR8LCA3pBlKkHfeTkev2C5PgQDIpYP5g0cEbM7F27Y3++eZgHDsaW5H
3y27AMWUMfYOixsUBHuj29FpLAGYk4VTs9nHVwoYuNhl6o8PYpbpxmOBDeaojPX1
RxLBBpB+wPIVA3UXRzjf6p/t/AmMQZlVXGw5amZEYg3wGXaQngVfLYBwiIki4TSd
MLOfCM21j6lcOW4UIHdq5+M2ywJizzsZoAvPfhi/r6kqGDF7rPrCUvti8DN6uYT/
3v/lTjniNgWsbeBktHDXmSmulNWLXJ584HexnMK8FsoZK5V8hOchUjqksVUD7lT4
BIzm0d3uZUBup4+X3fjPtjX+eoLgOBRrc0cE+QMygSl+nCodkAz/0gtMb9piSUFV
30ueB/dfYmJGYsjS7RtArE6ZAw6/ryAmcWpCM/dLGnKnH8k5sp+70oU/pY0CbAoH
wbwP3qKzQC3TcUyWknzKE70JBgVGJJdy1vNZOZiYxgbIGVQ10wSGOlfWA77iIUpe
1lQG5Y0CQQoXZluhSk5Ic/ChH8buUceNXDNHnL0g/ogg8LtNMwDgQB5TXFJr1y4L
TWGh29jKXL8Gp6hZDXd0O4NIoSp214J9w46IWj0+5RkVSyTT1C/xyURuJ0LEuhd5
F18j9gar1fGdfX4zFsd2vgE2g0m9PHjJvxgqRyj/meN8lFY4aajwj/+EH5xN4zyF
lhp93Lk3F2e10IKytmHtbP68TthraRdhnrAhF0tu3n7MX+lEPxex2vWZLItVqE/k
JVGpINSSvAQZxkSEMxI12usBbh/LqNfqo3xyrO+ORXiWyTqiHEwDhmn0+o7u4/mJ
BnDUWSWXV3Be4CXik6ov4fqwnIDRLunRPSnNmvB19jXuQts4B6yOL8XjINNKVVlV
zIhouUTGRdos1LC+x8H1xO2cqlmNaHDvh7bcOgJNOciBKCqiK3uB+UHHJKKp2pX0
jdf00Rb9QbhEjBQPs+99GtFlgOsSowP3Yvd0g/AzWNpV+yon7ALNYnsUup2wRhoA
DzvZIOpJo6bIei6zv36Y5Q7EI9ZSQYSElHcH2HtpiSpV30Ctlj9Gc6CrBu65sfZs
H7YVfdy123GUtB8i4VssH69ZT98SYTKTEkY7ZbiTKjybQBX4GcX1venFGWtQ01bf
4EiI64aWd5ecjhYDqt+QUoMvQAeLoZDU3vJX7sxVA0C3wrWvlAnsB71pXQKa/L7D
KKvfdP6SoSDQsmAS8lV/uKAFVOxNNCVNBwE4qfOEsg8p0lkO8YprdANxQ4uczsLa
5ZKjVuPSmC1tlqv9HS4k6kVmhM7sXA3ZI8pVVXDxuCpmlHByIfQUqIRRAq2dhC1U
AQ5JpTKlxe5ouY0e/5xVDAiZk5G+zedHvRAAzLwyDvXO+dgk9XUBIAJdXVfyDED2
Bj8Mwh3oz6REk983jRwLKXKVVMe1+ohs2ZOoVh/9KiGTvsaT2GCIeBgSbs4XLtc9
l+8/bPWTb3Xx8WnW2qf+G7P/wOwsc+qmLtdxnbAN8+J24z+0snktbRIo3jr09yY8
6Ma7WcTpmKeIxpzOnSFDaDGi6g0/0Jv4nVPIMg/yF9RreJ8v9dwJ0TLpJjF1F5kZ
9+Gm2yMs7nRJ0fHSMxL33rNyVtVCM1/bc+WJsJrZauhFifY+RY7/VWpjU5YzJbZo
HrFCiO030kMxqin0VCA0Wt4IeYfz3ZmPMQo++D/sEzCBbGYaBMZ/3UUESFDpQiOD
RDqmjNu+JnfgysnDJeR3U1tUu3pYrz783qvO5xP857uZFBF1ch9i0/YEzXcSyEMC
dUHBHR294A3NGHuTx6MoZMwwd66nG1VvRS/R3ph59tAhPxM4zh/A3YErPsweDIO7
fjij5Qp/wpW4JsFXUgHDEpIjFvie3xguqR7gr4J6ioYGve4RC8Ex8WQmBUtQgV0A
kkpXX7ShlHKLn2Fqn2ISHmIaRtzuJKmg70Pm5wJfznYKp2RPNyYq0Ibk3boPQyMt
IM7fjO1VFL5GyQCtnHMVl+vs0HAoRWjyOZQYxUtSBFRLNih6Kxt5cq5a/WRZHWCz
CA764ZO0E+gA0CUxxgL6aDlwUZNKa4NyywjHXQnFPuF20mQRpwRL0uHhHVcsx2TB
poI6yvCLIz2B6UNXvKxejQE/WIM+Qm85AM4jySWen9KhXK0u3Q35Ij5UWv63T8p9
MbjMAmxpRlVTwForh+LxFdxv++dCxB20SGRL4flRxi3LciFDPChJ6kqEz+33qOMP
tYvKGwnpnuZzg1KnIFUUHe0xXOm4BK1Ggk3pi5VDUOp9y6MUGfgAgD8cBD2PhtWi
Zti3RuhpME+24FedcTBKFVavrJiIqxykOn36LHlBNHA2xl1pfNKGSmPhVHOoYvkX
kb/mieqM9IM+QDPMejDUeb6Zt/DN+CyEjAZxRqEuL0i8bHy22i8/7/M3lXU5j0Wz
5KmiS0WWg6ImQZQMOPhl9Slb1mvLbxnoiSJEJmjdTVnXU/QKfFGlizMkr9dkbe5d
t4RxXQvV75asXxm39x8sSGwOJH0MAYfZXZB4UPISHGGn1kOrqsXVF+mxTVlCBtGI
s6aZ+qWIaOBorhljvqzfGU02HTY3AOdFaPAFUgMgUDBooedi9eSpa9mTElvCiNcU
abfFu4Cw//Kcxj9t8+JXJQwW/4MHHlKFcrHyeVaHjPAFflXzlIjFLm5MHEzcWDuv
/9bKM3gFpky3AeUmLdsAJcGFfDcGryCINPlaTd16bwWmRw6vhe9qLLN8Zj70KKJD
seZxkZ1+73xgy395dkAylPqiEg3CaBq7wX/JALsyWzUqqNBXss8b9J92p6610pRx
ZvC3cf8DqtNGfvnArad5Z0V4WmIftX9L1WUI89gMufaQLc0CieWRXSlQvE3KtDmG
VhudNN0mOgFDcSP1VW1bZuGF/xi4RA2HMyUh1hpGtjoB1P4vYBtLOqMPHShYfN9I
XLLKuoyP/Mp2DXDsLxxVJHkkHte0bEzSJKaxJ1OtFJAw0T0Xgt96uykzg1XuLTge
Mz7ClvejGNf4lsH8esLu9BGSq3r7VGCL/mheXrMnsCP/QgV8xUpbdn1D0saGbJYa
6qdrZcRG7X++3dYE2fWB88gwNJP3GoWWS0UdhjnvRPxCWGmor3K0K3e4vbhSsmKo
9jDIz6PDkSj5GxQ0PQlI3LsatBPaGkOFgN8GIKf6P1Z3Y6Fb6PHR1xMJXqagPIGI
vntQrcmZUoaS+dilKQ75kYXVqORRh/APfv/qvJ6dr9pnpb+GuEehA1XIvnpQbEIR
st1pP/xCdGZjutizq6tvqgid2AICEWxl9W+5XrxaGzGrFybyTm2kYKX5i0mOslSD
vdMMJD/CAagcobSx36FNeOKg12U/BunpSeauPSQhqepWu4bANyxd9NYhU2Af9BZ0
4ARi57nvvj8jqeO+i2mzUxUu/t/qmU+Gv+uPIi+XOV7GpHkLvzlSY+teF/9tmZyY
6wA9fc4u6bCIHE2KfWuxA8OXqsh5/Z5RABrXkBt0T2GTCiUC03l1orqrXZdtW6/w
B8llHW1YVIyQrvTnyEDET/0ByRyKTJl/b1Wd7eREqRoH9o6C2xIxNMkeEuov7F1c
yTUqGNcouH3iQjrfi6WI4xfhDfy91IMACk3dVPMzbTTaI6jZvs55hnwVSmKx29dN
/pZ/AjKw4SttKcUbe32cAAecQOaPnDWbPqjoBv1vj12t/x4QUXTPKVlxTEZztd14
0UxorPKeWrrH4VWTmmOYVzR78NIVldriDXEdnjS3CyKU++0ZKEh2y28wZ4b5g1Zq
ktFMR953Cf0qNovJIrkv+QxelPz7Xl+FMvUUZbGBraDcJCmk39V47y7s4X1Q9SFc
vIVMJgc28jNmwDXPZ9Q47Srl06m9fPzy7zsotMlLpScXAZ0yOJ82U5ruIqaRxnhO
fen/tm7SqTf2P5uhKpJbYfS+OKnLwMYQAMQbGGfa5GFbnSBfvhrW0ZkdGgt4PQTL
uqUE4DoIhV5w4JmKAgca6xu9zDA0y2xbPKD3Ov0C3iIoR92f3MKOxzKV8hfbvdLI
c/Eyt7kpZoXRs6i7kQi66hNLap1E+j4YqDEFsyExbtWC7G9lKcPxhmjUOUPHuqXt
QYwqElhTkaesqykfOx9/eFNRwnJ0CNjCak0RagcllZWoC6mF+kFPF1M+iMRIr5vR
7VZc/8N8zKjg366p6NhxODcqQPrGGdRAamqsiNQd20Kqme4e/wJNGbOp+++MkdAM
j5Ti5624EA7ehwttJmyVKoV+r8+Efw8BGDZnZF1/yhtGGRLJP6L/2xpFhFvaQkBj
Y4a+W8W+MMOzp5tEAuas7jXlZIcUwxqzFTM1zD3ozOQxRIe+9eO6bl32PkSfZG52
anjqR9YjNoDfufN1vSMpxZGwvLFJHGrj+xK+l0bcqxahGyC9ydLiztNGWu0sY0k4
GFQH1t7AYxCTG/Y4r1WhiZXfxWjASexFUGq0sonS8bNp/P2CWBUk5HobO4mRTAKU
85FAkrNKZSzDMzOOf45+lJGlV5hLH+GBNZvCaHvLMarDTvbKrFlsRvOcqX71CB+C
sz0UXcrxpi2yX8BXRWo2omLz1IT0G08IQJb8zcR3euHch2Tla/REC1epnP5krG28
qyv+SrTG43sIia0K3rpmHCawGHnhP8pu5UUxQXCClRXnbT++6gfAWZqKNUSgj1Uc
JMFdXB9Z6tsGkodtFOBU14q0Wg8I/qLIIQY5rOSe7a7XYUOt3GGgwrsJ+RGLHJmy
XvEd6iVb/C5scRNjuACfrFlfmYZ7vqpcGpPbA4WL6eTZSAplggZSFMnkap6hJNSJ
WBOII934PvCSMW4feeMk+gz87wVAnVc8djcyoeMZun92W+kCor/pOlFToN6fO1Y/
QyES0gn0RRuodi91n24aVR0O55SgPcERJNZppep2l7c48qFQYu5u4zH003X7Cu8k
7XmF7dm1h8kQCXU0Se4rmQJnfdBgKqfGFOtGRlXSefwtI/jGtCh58HheW4/s/gvR
J36yi9qzREVNDNhFX00aOb/dQ5ouPJD3/LyP+6iNGD1P2BQfcMKdVvWbBEYyJlyK
k/b3JXPAmLB5vRhVALGn35ZoeJrVOTTWAULrLBA5EwKJWVIhgGJXtWxhroo73Fay
6P4MuEPR1aPG31MeChnMKBGVHivKpLuiuXuCiProm+aN5qi28FOtD9c7VqF1XePd
aeuHe1Aic0lt/u8iy8m3T0sMAl6CJA4zzK8AKacTPS2nyphYDEexLC6xIvX5OYEJ
ogTE7gkpOpqFFH8yKJfNLu8Ti1vBZ8NMoWFHTFFkp2qqVLKJMYjVGIfgcj1sFR4F
em1E8rwWmt7laLePvxG0JFR4Mq/6Akn9Y1exYoxlUBBZbxhtgKaufju8O6KShqyr
O1fL2At3KQ3PKxdCWIK7fZUVqX+3UYAZOLSVG3CMBng++zpSpOsUW3oulBNFHP4D
kVj8AE5T8A3RxH0PQpMLPqQstryTxc+CGZ+WBnhy8PXwAuqU9q4n2xhKRolc6J+O
wnYjHAGbRAe65U/iMJLZ8xtKoijO27J6H+xq9AvrBqeXaA/Ybo3AXRn7QdYRhCjT
QPRq5dtNGYKEaO1i1bXMnwmlgE86FUkPbcS0frXLYSDaaLXhwBC+gZhV+fobEQK2
IgGfKH9A8CwNJdKoa455/lw0MT7GUj9pswbOvMooFX6I3zZLZRUihryUkGJSRrxf
p8sUnYF3vgXaIgL+cOqp/0eGIGdWTwkMli801BGm/w9zs0XvFAq5BDZ4IyQPUk4a
2ezXZXXPEu/g5t+4x7qHTZzPsnzk0b6kFtBJD0ELKDyDFQmlS+G/S+0FHmbHpxvf
5blbafjHGbk844HnVUe5EGKrO1TtvcKogHcYtd7Ade9QyNLolHtJ3RdaBn8RkGhA
K76KKhOHJdf62j9J9yoLfCDtyG1bPiwTUR0RnHo1cVEGY7HtGOeUcXWvHLWFojo6
d9gVVMPsngekx74gghaxvUBMB1YvcgVOOcPnVeLrzP2PdgHCpg5wGjuY+5UQA8lx
kfuifxx9pt6hgOArVyYGrE2G15mnkphLpiROsJZ6S19LNJgz0GjElEMlglLAsqPo
KLmCY8sYJJCnoYV9V9stRHTTtOZ+XXMZHEJuNmKGTkc1jWcIqZdGr4Ry1c6huG9L
Dxwh1t17WLDjf3V0Rj2hJ/vVxWIvjslcasBLZwrh9OkdJiWIHr0XEKWFOVma2QFu
cTCR4DENiSCwwpTp6fPbQFBD3p5pO9Ke7h9K8t4MYaa4qRXD350UELoOaOoiJar6
Fp5Z/CMF/Rx8akehGQphgbe7vcUMkPizHZngo/Qbzx6goyY4geTnY0Jc21y/muF/
8IWecXQ2/BwR3d58u1pa/Ux0ruwOKVGnAoDjIGyye+USQk7l58n+Jl0pH3UY44rl
eqoydBvmepgAAXLx1pHuvhrwHMoSJkkxIeX/+5zgZP/IIJk+QI2O2tsjzCcxFiyO
pOz9TQqF9p5j58XQpaXvZUGcR0SBmjumbsanuXaRZnAgp5eG+4fkiofX/Hp+k0k9
uTZYzDe16ylhdnROZYKLHRNZNoSSgrw2aLufkwGwvYwQ7ZDwIBQp1X0834AcbiCk
8nM85bsUYsTxiTeKUTqoYloDAc/rz2jQHz/pQNsREzAhh9rCI60ZfjHqVZ62FHU2
bweAkaDL0s+CJaED2FgoD4BoYsEYDerLAyhYPXQgnt0EkiIgLXTnDOzTR58AnAqC
/aokd3g0AmYUKj3sEUffDEMCYxdIo1VTMM6YdGbjDVcHCEucOcOrJj1f9ltqzoDE
m+o4fn7VoFQHIMks0fgNF9xfPy9swyTjNEbpcENkPBUAIPM7ZNQ/1N/X2/SFW1vG
Wnu43l4SWVxGfG/7d0eTIED+aOvPiRbQq/DgPO1jQDzL8Buo1hPUTdWePwUSOx3y
eOfu3xHrEksAZFsWx8TojNLz+30Lkybe+TesCISMFjHhO87L2r/9Ybsf8DU+O2DU
F2Mu9qyzB1OX5FAJZeEx5ARIk1l4zdsTY2kEnjU+of/D72OTXKaomU7dPoLJjUHy
0cWnCz8g5Rv6ZGc0456jfqZRsAVXfUjtZpkF4Y48dgBXwnu00sUeypsahlRSn9Ap
5CtWxfLPqHTeHNx+cRJmkBWzVqevPXF7/g4B3WIJkmeil04gU0Gip6xW7zQhSQOj
4MlR/aOPLsamdfuP+p0TkYBoYJ2R4qnRWFCA4JArpuGpJWHdu9wR7pX/65HUZHah
0RNU01zfiy/HLe2xH3QG3nnbrRcYGbLxOMgkTR9wK9T6U0CVvUe0iqI2Aq4ZKJKh
bK21uW4gmXY7mpXllCQbcpULRqmgeB4gT7q+4B2P9lLKT1zMfOGhOMxSeSE4pPw9
g/KdF7qrJJPz/80wVZtRnZ5Jhgw8Ygn3OQLOjDCNr2H7ejrxBpC49kPD4CkdJQDA
9JQNkJOf+EJsU610J+IuHEijoO41SvIpZ+WLe/GZWayfCyHa8OMf9GAzQYS7Bhou
6CNLms8RnqEvglXJ7+tOH6yiMigOc7W7nG+FYnRyvv3VRg1Xm37NwwH/7S/vLw0B
bv2i2dtPEVME3ctJRVEHLf50JmmSZqOLVNf7UoEJyr/I9tpt8Lfz+XaDu0xL/QHD
FMB+8CaxjLckSTpCOE/PYo8WM+5TbCJ2IP+8jU+nKDHUKKv10c+f4QOu/bh6Fm3/
vMjJXcIkBlEIVsOp0JARhYy6lnhVLHczHeH38GAUM8GZP2RwW9URsiqB7NW8CIrb
yAsX9YRMp/t2CkRAftGw8FU31OxlHLyAT7DKaJTEsL7yoPk1wIHEX14b6opabKEo
SNJMaU5C+t/hLkc6sRLYDkO52I3CVc98T1mneHih4x/m7Ns1/nYS69b9CcYIMgFe
wE727ORF3jRk34ALYTpYwDNvHCZSyq9lytRAC28VT26yJtlq0cPh26Mhro0/dIA5
WlOx15R9IkmzEBxn1AclDiiGB0GNNBLt8OMeotgJPaT8N1acvrghL3SJoYNllcQD
/QPkU1ySXMn5r/bNUkPukMvMWCI3tzLzxeploeoVanXbi/ZRVq/wAVyMGlSxnUNk
5yyGpCNrNIu7JGRiQVMq1MMUEaFTnvfoRx0dX9ugROmeOaTXyf/04+c07RUvLo6Q
KI/cLYhJf4doaf9tefGv2kPZBUkrFBfb1hYvFJA1SEjvA9TbGY+xDQ7BNvnmM2Al
sc5IHYQ92ySbOn/aRdd9Jgj0yf2GN3BXERSgz4tdRFUOIsXT73fddwVbCJEb8Jm2
NowZ8yKfo0xA2FYK1jrxvXCEDG7oJUCtKlru6lemYciFHbC2/31YU8FVlJ8HHZUB
tTKxYEi3tIOKclluHl9WkC/eCelMUFk9xOFIWoz4QfdZAwqBpqZzy7L+F1kANrzO
XAdZpuwXZkOuBYwpOX9h/l8qAenXY1DfRGlpk2GphuZao7UzGmZUFPECdyMkzeB4
xif5Jy9lQqqx5Iz8ANkqtKRZ2e0VkY/ugfJAuuCNXK0wi9u6d80mPdm3kZgYXVL7
e7PHxNmG+WAUI4NhhVKua41akuq8HwltB2PIPgPOsTjRTVULsInx/zlz3E64eyAC
5qKTsenzbr+FQg/FeeQlQzNjwlrpsQSWLS5O2cZhV9ScHEZYu3NOfQ5fI+ifwAfo
qNqJyBKnCFETP4Ulv2cHLJCM0UdNtTdqWxK+dJxPaoanrAM6gV5Rr+QfW/q2TXd7
7Muats/VueCh6ItY4gfqzsN9269Ma6uReBd54czPy4r6RfCF8owvoAMZZhuT95fc
wv0Ndjol1xscd3QUXXW/OG1UV/f9AjuAuYr9WVj7eh2dWobXBam+NOowLhJlNsOV
ChkjnxZx1OU4K1zVXGNF7rQfWX334SkJ2qDKlBkdL4k+t3v0L/GagaupNaeJJTu6
jDT4cmCJIIUaLbdvFLsZ0FC8jMh129gTvcnjfPALE8p9iXIuKCGFvw083JvtwElJ
7LV+sx0SFvrjuBP5OWanAgLiguCSDzmFv+aIi8kpq4LMWTS/Y2dx7CYkEkxVNg/e
auJmc0WgovKH8nLZFMXZsXjmEcY7+rBbMGnrRbwtbrjyFdZsaFKMg1aR4VLseeNc
3qqo1LcpuTfFIsxWuncRQwKPvmXokiRMegC2bB1e6bCQ1cGr2OYVfQdeXGlVQ1gE
11x658Bp3egoXH0XR+BFj5fTpZmCVyfbhFwMhJl+3XI8IpEkWCABBd8q6OcOTDLR
DQf8Fr3mhvjYyh8vPU6pMcqxaexJgGir0ZukRmiFnx6TjvlQ8eATHryrnyIhe1nc
XO1EKDCvn5Bv3sdUSfWtEG/OZWomEISQ2a1HqOdMfJKhLSPf+jBW64dbAlo+noVJ
LNAgwTZsly4NoMef/ILNt+FIq7ZGa9czNCsG5/bp2cRKpXFQ6dJKQdWC9efSDSAP
2BcFx0xjCM7u8eQG1tlgNijYPiXJQjYEv408IMVS22GKFemLJWkAzxFLOldiP1Af
UH2r2bCeazWhzC6FvQ3LdbOllIu/CgqRBQJ38BXvhYeXkSsxBGYWwV1NWyu3nT9g
IcNsm+1eSsKuVW4bFwyJFlZzd9cNsgmCr9SIjW7knsrqw0OnLP4FaYM9dLhXIU9v
bdyRVmMEdbTFhVVAqSt/h3gvZf3u0yKzwd2VtudCYfTmejJT61PxTpSpQgnlGYQy
xKAxQziNn6UjSel1lK9av8kk1nfbLIlZ8HgP3Z8gGQj/UaKqDUEXbE0X9FTX+MhJ
TVXqIdjHqXWHqY6h2fOKVG4y/VG+raASscGJrdTILLdmvcHKurikHFSDB+GWJ79/
iqAOfcatVQnICLReAz17g2icZDv20ZXg9sB9tvRmot0TnUUzpy5FAJOcMGQfNMbW
LVSnE79vQg3wPTCCNUuECvvn1Co6565aaagHWmGajvXSZDPBQcNVolS+UzY3fi6X
z9OftTniSbxj4qKzwPz4e605YjcQoObyyubQcRJytJ2B+jE5f5yCv+M0AfAonDzx
qb8uFM6z02YtEJihAbLWSAO4xaYStZcAm2AIYH6qjlxqFjL6Qld1kgkVJs2xIBwO
i7Y0D23LVFsU4aujApSSTMxMKhh3snNdxglZ3gOP5qMPiQkTlmH1K/kOaigcseOL
6Sx//7cZ/RqfZqm4MCH7x9cutXjUHaHNlpwIdlDnjJ77DvtuzoHF4ET6P53BDikV
dCF4Of1ocoEp0gYUZH46rIAWbl+lUfDknp9uVZ8K6YzEQe84cymxAq1iBDsf9rSH
b5qOgV/pJoQ8CP2gqq8ifNEOftokjcd2Df6NqD+2uiDp62dbQXdWqQKwGwn39Xj6
EN4LEZooQT3YEHsYbUPuJQ/hitJcN3B1Zc0PKB7VjARej9pG9uUryGHfX+bb4tWl
IY2+LFwwzf0MfKHH1+j1EDZ+QfyvUApZND+AyJwPC2nyRJ0EbOsihzCOuYPhAjlR
JVietRqSs3EpdLIrBVV8ikGuc2JhJnNOlaaXeMDN/xipdrXZ8sOhWlzzUlMNUqSO
Sf583XIKLz38+vNE8OpuEKoT3G1BK7/VC36dDDP/+NU4IkavW4wQyveYY+W7xoIZ
MdQQ2guc5HVdtEu1nB9Y4z3yFu2q4DUxSmtXmPVRxaIQoNipEQ+FXaWY5VrNfGYx
Rl4YdbEXqaPyCGL3BgQ9OvG29igB9Upt5o0AdvTUw66UoYbpMtYcARIK1DCw1pGJ
FFk/jIUNhG0QFVIb5jvgr5aB3ll+4+0CcPNnG137Dcew11jllJYCY4Dm2Os0H/X8
6uAwmNXV7QZP9ECNzxEeL1hVX9kBLG+qHyghkwxY/GuUnIFuQgvbfBjZyxa77Byu
CtnYoQnwsoNwtd7KnsXOsvPM/6GPXTpEtpF/zkIO0PS6AvNGwPUwwTTU2Xmff7sb
NhoJ6k5ak+zBSOJVXamZPcTE3eRJR0zQ/gHJSX9xwv88hMJtjlszSkmyOsYFk7BO
T1hasKTvlLmJnuk7IDu38LOyF9HsKVfp1D+1d0yrspKRXYgBEZDW+kbTOUW3bG6J
Jt2ej1qXZrnboflDx01lp1fFZJlnh+uwlXE8Nkzi1H+cMLk44iwSrVgqYlsR1R8v
15NkuiCcU4RgvL25DixmcyBDiMst+awk/UmgeFRDyV11xUjk0XSCMpuQTBxYIe7l
j+wPClWaG/Pr1nIRKxH3Y/74MKp0ohkwQQDHzuaFfxasNMe0QqR2n7spSRNJLgmt
eBn/9zOzWf+cUwySDQTGU1dpCMeY8jJiGOzO5j0aWpFwn10arCD3Prh8ZxyuBCXw
StE0O0plZER2Gup8M4ZpNRMXos6qMiPxnxXBaRBY0KoBPDBMWe9InUNuW0KFYXbp
kn43hTZPw5A14AfqROFZ7H99LRNVusUDJi1HPBNH29UeesvTXZd00zvo0Nm7ItOa
hs85QR3DlJ6csD9EdceP/wIvw+1923qrH698nRLpCez40+mEJ2uFIqinTAhRFNp8
8O1FIkvwAK9MQ7yOI012ANAz7mS/3CBAxvxzIWAeMaqySfV6CdXlt+7SC4QQa5Z2
U1jH8AyH4b56/WLQo3y8y1jx2VFGAWpZvtEABDQ0cu0F2JCNAGI3EvXOZ+Him6+b
CpK+O9osnNyQy5HKYPhry4djixvlNhD8IYe78oIxr+Q8OXeJyxcY1L+YUJCmIhVT
4u7O1nIGtwcosdx6ybGC+4Q/bq8DzSLZmrB5O3YY2kMbW3yhyrsZ2M0aApqvLYll
uDCKpT2rCGObdrwmyqHJsvsZbhS8SHee6Os4YcEWXIW+zE+iAKGoR2Ts0l/3dz4t
48jf4dOEEiGY8Fo4v+Bg98Ad7wWmbgI1hZmOs66BBraFqIkiHjEndhZ5nBu6bgnb
cCCmljQvasWLWj3CtNCRWYf1PpWxeJGNFtfDMVpNhRyd7TSybUzFrqKRJLTMjIwb
58fpbPmc4uQoBwpwmtbtjbkGKoe9h4cf6kp/w2i0rzs/xjckGkCVyEl8DNdwmYgj
8oluvFSErcrZa+8VhBqCAcPQRJ+/CnPbdxVVcXi7RAKBcxo7bYfPgpJsTB6PO/00
esyH0hCjRd8BBsLlsABTTrD5xPTpRv51+BqRL8kemWiRHDenu4HIXdCPXfYPfk84
mpfVRzBoIooIxmZqEDWgpeZK1x2WP3ePi/lqgVw8md7dgu2ywVXOX7MXsB2WtvpH
Ya0/VcMyWaFj88FZz6/iCXlN1cmYoBgerC4ttQAPhMLv/V6DYH9i8elS5w8UiD79
21jDbIBH+gt4W0kI936sCrDxReH3SYvuae/eLWi0hLRuz7dIGvcgjSTqOz79+yUm
iSRU5kpG0TIyuwInpLiwzUhICzW5slCgyzDngXniDdmTDl/z8baiDvROgAHMcnPJ
8xnlENZRgKxUzhRbfpYHUHd5Z+x6U7MJ1v0q0xwFzO5ri/OKfkLkooSGOuuvB578
D8MijjmrM54NAB/oxGuGssLcJmdJlmqFuQaoCIoNw+hQW8V5Ky8TpkYr7c+IgDge
ES/pYjXZRChJm6htWhw4HceaJRZV5Odaywk6/fwa2tOf5q3mUSAz92dC+DADkIpF
0ZlaHe+rqkIV89NxFdcK5+K49/rtHrLz7ORbOKs2ZS6H+9FzRCK86mdMutb6dXze
le58XOw0l72kujPinecttGMyXEsQue5A9HrbB/LuBmUN0Y22OHrFR895/PZCbpn7
6P0vvyNM3ZjYAmjATeNJ75GV7qnhCf8WgfdPjCQintTUjFfX4uLbxpgSLPdESiTw
KSU59llno2Jx9nlokmmWa9ibFetKFcGXQ7ZjALnQvvUf3OZfr5hfhDsxyZVd0l7G
55tF1RO16ngHweD/cOEhl3M6AfFkjbbJmvsoF3qrMOPQ5Dxj/4b/F95q6LE2Z6sj
P5Ne1syo2jHEvqAG/VX1JVNaJAGTdbekqYiXYNbO1RyDyU5Uz9iX88IbAOvUw4nO
HTpezMibz6YLcw5uunpNiC2Qp2x26HTmfG6ZT1CZ0nZio35XxeQ40xsvcAJnkecq
woxcaGePQBfnT1OvTzX2ubMbFTV5BEumlrT+M6aPvLfrMbLmCxQ6SDv+P2J6PcMu
Jjy3Bdyq+jlwKFXjbMuz9Og+cc47iFlwbRm/P0m9saHX7Y3VdK/PzOA52nbPuQLD
wfwzvmK2E9Yqz+6n6yr6u621YANIXyz8o0KF09r7O3qL01FYCzyiEui5+vTSRKUc
OsmZnilK6R6GQAxdtmQwKT+WFhZNqxoA1YvqyYFXSC52MvToQ2GR1JCUPJl6vH6P
Ood4+7THZEWXdfV5eYpvnO8nTpPEOJqL/N6lTpp/ynOwaqdQ598o65DRx9YBWRhW
l2+OxbIQPF6AMcjLOaIVaiZTYtts0Mv4HHqn92566izdKRwlwrCbxFg1VZ3vYkeK
PdiokFObxwE30Y5bBrz7gntOX8DJqwFgAmHFk4uOdL8gKuE2hNEbBVV2HCRWqJM8
JIjuaXNx+BIMkoYRp9BLaDhIrr0cek52xHZy5qZ9QHt0uIigX0zncRSm0EP6cV1r
sb/VlgkRVWf+uGkCbfJzJqpvrX0aRTCbKOuU/t6y55lC8AVkEi9fXRHrmIw3b/lj
I0twD4oa59oGoLcxrGam4gBvfHQAtg5W1dUjWXanNweACKgF4hetXD5BDaHuTwC2
qI3sQt2toHmYToFbgo5ENtFwasmN64uNRCtvQ5khiPLOUwvBda466ZHuc3NgTIwh
7eh3y++tmf6JHQkhUo3Pem5HWSWkKPT2J5Alp4YXMcJiT5TGAA7Jzcg4/Abfu6n/
ccUtTFOLFWawLZdc6mBN21YxFlVamDoBN9X8iP6Uhew+efS1udLoA4A1fnoNeL5m
LJJhpWczgeV2/I/ZMXd5lOVg3ahASGPmBRtxMYR0F0/LwVdO3Tqdec13C94E5oIO
IUL2nc8pc4O82qOI4IB8uScy+spqZyO3fEM006Uc87rvtoX3SdvukmIVFkzzB7Y6
kD23B3QlgRky9Nj1b4hi3Jiw/0Mi1oz/QT1vjnVYxTZJb/a+kHM7CKQavy2L/kTS
kJUbYh/8WA1CayyTcriXmXfzK2LfiAuKh0GjOBfhvOBe97PJIGI0AzWx7E79qkvC
XDqgpuU96VWkXGp2LA3ZVKGUODnMvxUrcOSVezVY/h8omFd21HPSZ2cLbFB4BNhC
FyqBuuhoct+juet2pKhd2ZGlmBxKr/15HdHtWDjA2EvpNBPUqmUyE/nwE2CYhG/M
JtzbewfJOAHCVYYgVIkuiShSkWspl6ysDCVeHhnoUswa8sQq0bSeqQcaMcQb6m2u
Q6nue2yNSkkEFC54fRAJI4sIxdeWSdM3ka5uWVr5txxPDTIDaODFIHLQMOaOnC96
y9WvJ/Cgd0Qd1HO/oJg9yNMhLSmjPdDcV3tZU5wf9HQIqK1QLOVBy7AtAH6hX18s
KNmvwOoDcI/FjuJynaAguJWBMilmaxm3A6FrjUaxtPgY3Fx4X+GPBfODAp71+Ii3
Is5G6acBV4AeAv1pGb8E4Ni086XAj7++nFQSbA1VxYBxk/9HDkhMkyHibswme5cQ
LrE3eNtU4NI4p4SN0uDyj02Vh/07mj05Ru38uGv4zs1KN1r7cwU7vIzCdkpoZsTy
AaWcu/1IzjiL1vk+a6g4AHlAOXcw9UWm5c3zikj6IbMjE3wmrC4GSrcRx7aRkObq
2EgbgCUYsAU7lnjLT7eOw65lqCTV7rUiNsDjwqcr4VL6utGglR7ymMDX5Q9JyXTn
4DfHX1mKJjNp1n/6P6mTFSrnAeS+vcqn9Wr9CUpGT24SKvjIDME2GRKp8hZytyeD
19HgdoBjdFrrAUbIlweX8XC9Hd4+aXrOKgNdC7lTRBokWmY+EBWHJ6dJo/YRGYNB
BvKCoKypdpf0WWkVhrJpTg44vUJuZKdU7zOuwW0nBpAosKAS8XUFce8NxEESUDs8
3WxqjqaKm3xBAQkeGu9mPi/YcKn5YRGVB16hSmcf2Cf+9rU2XicFwg501Wg6D17h
TUiqLqyGbwDffQw98WvPZ2ZaY1e8lqFGUWg4fvPMu6DL1FiU7xyIZAMI4IFcYM9r
XkoKcd0/bQajucSZ0/ZNOGG9bYmkRbO3MekszrQXbqsLKi7wQyk4DkhzYpjCwW4I
dAcEsIwSMv42EZlgp9SEzjU6uu2sH6M3ALCILgIpBvcsaOAoyVBiFyYlJzXlWSL3
IdSwstTotwdMajEkAfaRrf/T0EBYmrVqDBYiUxBAk/gT/mUeyEIsjoT/+Ip3bh3l
XwMQDRts0zR+Vxbb+Xl8vLRdPTEcJeCFZTHLkzcLic59TK+1y2uV7sKHxOAT+WbE
C6OO4kN3FrfGU/Z1eVOiDnQGvk+lxRPlfOqBlifWvhBLy3NLEvRCEWc0wVyBdtUO
D4PU+gyzioooGI6JERAAhrRngt8lOFncy90DyHW0AvxIjVC5NJXeH3wnrUyKR441
FN1EwYnGVkTYKp3RWN9jkNFpmgxB1HG1t1IgNhNCLtRYjLcQxa2OgFJ+THn8D8FU
rdSLaTbVRUtKRBo5at2oDBJJ92+FO8TEzZNgoOMDL2tGh73kJX/SpKxW5OQb1TBh
Srs+KOdkYIZxN+IL0hwZajqcYv9Gw7jHeQpiqXdwAZrYcFVWMU44qYTW2B/HsKgA
lIr/nQugKM5NXKhnUZ68Mt0Ykiw4lpoSXRsXUMh5d1ST34t1IhXwgLByipoiGi0b
sUYKumMn65RTtM050AHw3QtxLd1McH8n5tsFGhC7gjMnfurZRFGwWwnDU29PKxIA
JYgFtl5jp88tpaNvXVFXGjlXWYRsvq3qCNHh0pryzS/E7jn4cxz/xq2RfICh5XWQ
VtfnFYyO28MLIjJiHJ6NFk4qp2LF6cON6gR0KnzYIjg4GvEU9HOYrtonefC4JAjD
UealbVZYZWVfbnADnCsoZkvkOTZ1IQ4utdtsNWvjpwTP34POiWEbocGIaKzLArzM
nqXIBf3qCD/6K32IlXFR1i8B+jwI4H70vmFoNT16LOMoXt5jgfi6o8fVkzQ9a/fL
zqxbP4ey3uU1gjGjzP12xwIakNWXVuHYWLP0aj3+fLSlKzAHX99ektSoBkKqFbr+
u5e9LYelpAqmCi7p6Jnj9FtPKNqAqOkESaRDyF26vcXpyvF3JPu8CXfHCg5irTIP
U+GFwjv7IxqKqt41jROlrJHZ3V5TiabMxl7h/tfVY+Ha7oCs68WUDfXu/+sjdpBA
Ak5IwogT6ItByi3dU355iOjNAs8NRHVeqJ/Q5au9XLsz3TOm29I/LXgdg8NKNEuI
jOhiFNapNNn2xoVHx98jPN/EB1nmEMP/08Rn6XzJZBvbPBfTg+zSGeuCdvHROahs
kZS2/Gnh4mwIvqwng3cAXDRiL1AWKZMpGPDfBiKls6XctcYpnG9Bnmfjqs/HA/ME
vgK/CrycIrbBeFZXZhmMb6FchPkNteL9ZbkfGXJ+Wgd39gLIYbBlEriyYdTl3qRB
f2s3gXb75lXz9qpbgYHx8VNqpFYUpvNAP38YSwOT7PSuAg385Io5oZd79VhkR4f1
4icHNFfZ6jiZn9oeOvKglvwjq/Lbt2pYkEcjpR8idMUVhQTH1uobPhzbOOJIm2wa
L4Wb2SgVoqXgj0zSzSe6Gv0QuO4TiwgE5sIuVkYfr5p09yTtO7SgMQsKXtVWwXC8
jwBL+AZ+esWiyBLShnzrbYC5BfpuxZf0IAyiFjaVxetYobqcGRZrQTG/uciU60zq
g6Uh70ZIuzqsbLOF8kaw76iiX4qL2asNTwjUKZwUFci8AJir2Wozh1s/4MZJcBaW
HWxUID+hT3IZGZcenzM98fnaGooV3DAgb33k12HPaYQfSNPtYXoHAV8Ler8FtmVx
j2lif5fQT5SsFL0FT76+ohZnMUKSwb7KLW8Fq5ERhmsklCFmVEO8O97uX59Z7+Sv
et2lTMEictTWHo9LDaVDwstgCdAjneawhcAsd7TtNevzaQgiTdFRLy3MUHi1ouMF
BMjcQ2vYJzMYlV4teZ4XjMduSU7NzFHBnsQfoYV+tsLVUJskWbqCyXZf+Hdx66J6
9JsM0HKF0RFSB9MoCSXjW6vGNpNosP0Pu0L/wkeDWuQkXS4zOSYoz+OGmF+ERnOA
8R8EZr1BdP4oeSCwCj4UNzrYpR83riIOFNLrvlqtOJFOJezrYd+eIW23FqHApeMr
z58qjn4uVdNVaX8IDN9cJ0XWsetRL9DDCW0XZYaoRNo2eqV1FNP2tCO/aA73YYDY
bdpOxbwrnMwXZE08jEEVONjXVbUUtaRshsS1NiWnR8Fiem0bwWw0c7YMYep8njxL
VVOsVcOeKcVYSA/AT4k5w/UyPBYDp9RPRlxKoMhP28/JQxf94lLdQV54zwPVzfY9
TKiy9uxIo/E/BtMC0l26K0oXq4XGhQMRZoqW4gst55Gtu0fGVir6iD9fXtLGNscV
4tLR43OYOAJ6j9qu+5SE6hsGWtH7st8JuNdUfsN5bIzhiB18xRR3jkY1eBElliub
LPiXBje3xO5fpOJgLbDBa4PL1amjVpSMcLA3GUAM/6aqEISSd1itwN8dDEfjxENf
NNQAb56iYODHZOF31LPgItIWPzAe+mTyJ5SRhxq3klVXjC7ZmMHpyVm6VZvLwts/
0ctAOY/O5xKt8vNS3B5cTGuyUdyNjrqJI6jLosMRV4hVHT9vEHcmKI/rG5ZK4yib
LI312hjOXSEwHLRkPzgXBVyqEX6R2gRG24mbtAQSXi9dmHV/PiRwXvP/ynBGDLrj
e74DwLVaH17zAOCqcnzkmSaW/JnTcf9z5FfvbGlr/TgRIjG6O4sMwavpalrMlnSG
+K04Fm8AblzvNRA5Piy/zoh9O0TEdQnOocSUBZt1dXm3fsCwMhYEl969w1q6DN0H
LJcTxxMkM6y9iauVSX33vWsUybp+fJjos2WTThMHbDq8uyXBc10qEJ6igAVu13gq
IZt5CcMfMEYFz9i1tddVK85Ia55A+odW+Ra+waECqHSZi5Hk/E1nBy2r0rT6n44N
hTydrl3KiLnVZ/FNrvP/zXsjpgTpBpt7fMa3Vt53SkCc+bOzDkyFZUWpo4YgpWDE
I5f1QJGfxsbG13l4daxLJMPRTARhwy1hIiHTSfZ4vaVw8/6m+qSIRys7A4FDFbj1
tmRpzqi0Rs1a/JDLmdO4NQf9b88daUAaHzVd7qzH7ZlCfu9OvA+woAvLxBsv/ECl
HqL+GNIaTiFGbP6GHsWEZRwvNngJDj8+Q2iuQDuYEFvKyS1Z6ri/n3+ZRb+7ufh2
y+U1lvqEbYTRrRSwOfPsiQq9IXzHjAxs3Z2qWwl6Mn2hTvrLAscqvJ28VoJTn6jW
LAGTk0bpQDZRn4nzQLbu529oKdR+CtgOrZ26hpVn33cgAOjhqZPcDvdTrPS49JDW
w/tu0fBns4bPzIgg4AQeQhBNcBfCIXjbrNmKQX/E2rLvJfwngUfQD80ub/zPOOWB
cZQ43IlDQ/buwDQ4BjZkFycqKTQPWMuEiJuk/3K+GYtwM5W/UAF92wLaH3GNR10T
sipdt98epkWCSmj6lTaAF+W6WNZLS0CMgYKtcVJjNltM93OrQM/aGbM1CjZiKwlS
DgN27CdjuSygUUfUDRVW9ZVBoENfhY5nrb2zJ6YuPvW6MZW+gw2KqzcbK70lYgn0
kcKFNzI4vh5zCCPXgNd/UB7URvN+KCvmTwgklL8VAel7wzU8c38385jT2dpGetAt
FFk146/tn3c1jk62Cgl56QtVZD6zUss+VPBsLbiUEJ2sFL3ag5ltCLgHP3yfia5j
eKcTBRz7BpwioVeyaNsWyqTMGFMW92vgaMqjwIcZzdI7OtnGUVLgcmlhUINwqwmx
m4FTdW2wB5pX56pDtLhXUw+IMFG5EYDh39CnsXmc7VvmdKt9Efeq7iImWOEVsgzO
o30qbH8zpPU7iDqD5jBUiwdX+6RPT8qOr6QgB8ePXSGseHWsVPzVZTU49ysuYf/6
NwDmqonVWCRERsVbkHi+E9vbZgCA/lJpCVX0yXOkg5CQv/xiYnrXWgxi15PwZg0o
fMbEbwkqGddrw1FSdof+X35UgR2fSZzdqVbXy6A9ZGT/Bf5GjIl3CKsUrsIi07Bx
EmJcNvE65ejxUGhhPzSeexhGs4rsSiLX7v6ehQwxo3YUY68GANXjhUn0Endz9kzT
YCxcskXDVr9SBxhgSuSniz8SheeHIQbvtzgtQngzDQHfVkEhm6uFweIpRCD8M1rk
SjNvIO2IMXWLBOjHJicqp6FnkZTjIJ0u2OQ0V5aeVcUaEVGO/NlwGeH7LvECvW8W
T7JhN+xZTOp4jAJlxWava3t+1Yo6M4j0BzNsrPw1xAGF9qH79HJ95Z4jSdJjgoaG
uHKZwDGZs2MvpIfM8Leo8xgI3UOO/HyQVCifPhGfOEUpsmyTzihooPoXkWcoyDVe
HLRy6wexo/Ge13XidPNXfssQ556YAdBUl9lRcjhFAA9ShSdNI+5TWmQJsVaTarV3
OIfvYdqD0Es1iEKFRm/yjNhZNr1/IyPKvZd+G4qaE2+R+4xxXfP+xC1+HU6DpvfC
EKpEpDhYFyCm+RgMsfcZ12xo+I9WjrK+hyVBOUSPEjyRhCSGb/+RxJ16Cma4usBe
8TECq2QZRnWe5yBbdfmjT5q+dRbz9ad6tiBlBD1k+1bZGFSdUOPq+GlQ/ZOa1061
v9ZCK8xxircORWcCArRb/cmk9L/YzvyInc6PZe+VJBSY3Yxh1ofuZHs9efqYtNxq
Sax24fYC9GWjDAXU+dv/d7AYAMkYXsReqUYc7JkIafLVZR9lMY8AmUz9gk1d5zjO
N8NOLJzVh+FfXYoAZ1fR59Gez/KswC9nte+7cDHhOLgjon3LHRg/E+YlDPysabRM
kseMwUPyYOknpcnGVlM60GjOBnENF2st7apW+azFYhJ2bMZyzMXMqVTbbG1eneYD
ULR9LjzcTWPNMSJ5ICv/GZNNEgbMqcYDoESvBldb9GvW9YNTsiRPlmIV4DpdeXew
B1PzGvx9QQXrus+xUVoa+YeOCSTcsLjNzYS0LmF+X+Ma5muTc142eCLQO3gJL3Vz
vxFBvanFcHaTsmL5KB6GvQrOrm3RpUhwiMiWr1Tinwq2XrC/C/mGPb3irZjmA36H
7CsdvyAbLHGA+qAgqiuadHbs291C7Na6XH+k3oH5pQeHCObQ5nYnU42QsgF3J7X3
PtL5ma2W8au+TCqPi9O6LSsWZIdeJvxvVub9N+vAGdMmseKEjdYPb1+7SHYcpVtm
L6NmNLPWNLFSu9bRMNP1Mh1Ce34wm9rJwkIsmLpB3Lo5tWUqsxNSRTV7xfr7neQs
mElDQmVf75uFAnp/2zj82YoYCATZb7ezO0wmyd9y2DDq3b7l4i8RYtrWwmgpUvJB
1i1baGlqfIL+pUeOTrIKKO6GUKkaYxropoWB+YkQt172i7XoONC3S5EZdwO33Txp
0tZbn9KGEH4yeoDdGN75vbru8mpxgwzjUw6vcxa6PkBqPrZNA9u5TIjLaOSYNTVv
9pu6iDi8gOJfQqfYobP4iZgN0B2KasNpywsvAfHcNbMK5a/Q+wmYiix2Wffyt6mz
3D1rw+tI+JVP4wyRRGMI4f5NIiTrs36IrEln+JQekRxkGLXq+uZyiTN28I1IjXCK
g7lMkzIF8YMpXzRMpXl7nOA4H1WTCwg4tkckC4fnX7aBAIFYcB/hORwcKtEs/boW
pwxd1nnjPdHXsVUVfUsCd/dEavkN7z9YHQNBP0sM6dyz4Dj/wVWmDw+r8lk2+MpQ
XNvYEFZb/Iu+KOu/Srs4/E+ROUYKKqWmsdxc3qD+QZ6HVBoJyxUP712Ro+c7QNGO
v6M6nQZcyhLWPzQAYIKi2DDuIr6PTiiCxz23LATKT41yigqFYM9JsPNgJYou50TU
vqAdyG7bNRwe5o+zmGBg1WFHYGSa9mDC1NJcUJybL4xZg2kHaZE6uHmmLVXTWEWD
nviRr1F6/+JODe6dDe0l2irMAiD0dCIQRjy/cRGtWh4k9JIQ4ROdnsApQLkUFfnl
utceD2YkxkhKeIDLLdnFz1NE5Z6RccuRlkASDyRTX2905gFL7TiUiC0zOqyFyeMe
rBmRUO8JxEUXCS4hU5tUQNNhd8M3+0Av9mc8+H05Rwjr9TCXg33VC/P7aboNfPxm
SyC82ws8ToZI1R7Lgzx9oZbZ42cqKQQVVIIWCkXIArmrbikb2S3Ko0ZURuQdP23f
W+oQVYRPygHbXOecf3PUy9bQ/fNPYQu3xa3WHoc4WiS7nslrlVAfThfR8KYm+oQ1
7RBZWzJg+1GuqNFPUCX6MHN+pEUleMpCXE1vsaaf6X+AVibp2JD1tG5/mvEkqdN7
upK/VEHAuaMnIhlYxamcJCMwA99WwgBVldPxPALsiDHAADC9iC934iQ9IqNNkrBQ
30AR4LmdRBp1S4oP1IPnI7k5WkWdZ5M9ixMgyz1FK7nCI3PiaKncnA+kfvXrz4Xf
q06H8haR+I2DJ8o1t7gnx0gUhCTvx2o8DqHyZBZYwdt2yY2zNYMExHDPH2vhsLUP
LEn1ox6HTyi7+nlrqM5S9AonU3ToqibC6SdZc0WKYNEFukp61nP8FvHDTt1GfeEX
pVxVSDcQFObuN5mRMWOGCaDN5h/aiacOwFHhskWtmuP9OZsdgqDvPSf4wLe5KhjG
yl2C7h/lCKdmp0K5/ILXi9Tg41sa44mQh5jAG6jQTc6a2MIwg8/VF8hNt1DaSn9U
mBHlcZ2v4JtN+QuriOW/9YJco4f5k/D/q7DyBRkMSQvuwCbkA/WKy17jQisBwnSd
IM+Qz/NWCnkMDp71dQ2T7HvJI25uzEyT/JAHdC3AClc6b/KD1cMOws+0xtdZASDh
T3gwFmLsyGpJ1cnH5jrOCKDUtX1J2JIoXdZxRuJkDkQ2hJP2n3bjQndJuXC7rX+9
bx3+aaXSA3jm014r2Jmhdz4VDQuVHzA6w1Sb7497bWXnl4u5J68DiiEtBWa6sDkQ
+wdcdCxbo0K6JxX8xmLBrqle0RY930ahNBEBQGvGf0nhHFgSWAYzJMlA5B9C57Fs
QIytzO7xTbO34sphBsoRHkCfGs5nOzVs050pa6aTbGQ38lGxTSaPnQdDhzxfWfLD
U+AVfaBUHNJO/m3l6HUhowXeNiG2WRMN7p3KqdTQvUaCLOe/0IJp218rJr60HRzN
3CzlMYZlihZ/8WZebVkhTSk3O909dfFq8Pyc+MLrcjzzSd/BBGSQYbRzMZNF2h6a
tDwEO+EbZAb/sxrL7iP0+/FhFDUGC3YMcXaCxSgpw7d/BwRg5NbeDrw8F0knBYD9
Jfpuw+hCm5lIJj5zEfU+geomV7LmT6QezK6AdLzgtQhvXAL8q6woalQvIpYSpc9i
o2ietwQjgDvbHkXCoQIiwkyYBHjevvR2GJjv2sxDxDqhksCDNb5PAKy/4DLj7pFe
XTJzYYDEf5kbLqWoH5Y10DkwufBcHa7U+4Z5mC84YvPeASyLQXCuzT+N3Dea6+qK
Jk3ww+9L7vwedg6PNwk/DlzpyOVHF5CpZ5PlkmFR8fTu0dFZdOP1c4SWih0/nNfR
Ngs4pq+LzLkmfil6bVAVhVKlbdqN0OIYuN9IieZxdCL90FeXd/KST24ncY/U3VQD
kVeaKFoKIUSPBWLFb/04L1+v/7DbATaaS2AS45M9lqIeG/bU+h4qvNmemybgQ3NR
rLgQhhoUJTzjDdhrCYWas+0KfOOP7MOYDecMbzTYHyCFUqme8ZqhbPsEVCzABgeb
apDnEQYD2I7HCClL/vLADt6V4yd3Q4fjLzFZhIhJ/KX40kvTgPBVox6eeV56j00A
Wl/AjKk9JTfD2sr2SLXSHXNBdO2VQ0jBTyjiXENVBekFyj4rhTCeKSzOjlzGUibq
y9gtoBPGZW6mUrr+DfCbJPDQ1GpTTtk7iWQG/uauBrrWz8jJ9nHKnNPMz+UwFvd6
aaBXlWqYqIARa4YZqtpBmGjBht1RuhlVHlqhTqovlrHnlFZdbn01akDZ6PAg2YZs
Yo6buYWcaA6th+bhPi6036TkOSlIaCBn8mYwBjEWJ1F7HidDNPfbED+1RYdLqfai
7/5ZOolt1TFo9bkRSxMXGkjOoCllhaxNHuAsw3lXI9ZGB6plfpvVhP4iTpej0R2g
csFAR4Zq6ptTn3FXppLGT2HOmBTTuwNZtvUv1T2iLxDbA48tnExclkhdY9N9dF0V
k8Elod0+9BWbGJ+7L/xNxTRQr9NIxqHH3Iw3tpljK1nw2oHrsVGLIUVtGLAPurJ2
+6t56ykSVCFa+YvPzq34eGvpmv7Jk/GhXPDDF0xpN3xwzByzuOsTYYAxOBOy0/ml
P5o3FmsEemq99hGWqj37HEDqSI/7cOdtxTWDRALdcGRwumFGg43ZWI1Putx4MkHY
5QA3IbTErApMXyHimneJRPDoMu0zX3rBRfpqTzLoTlCI1E8U9AW6QtRbZnS342FD
9rwlAmgYx2UX1+5iVbWjTbi0i2gJSHfCsxeTHGwJhhUtLyDdSUdG2CB2UWjjzne0
z75ZoTgByeRRt1+bh3VcbRImFJaaVin3PRqfDNfm212O0Hjgttsn5CqgjIaaOWXK
YPdpapX4cy59Zl/yQUHua68fN+5B+HISp5JRwVCfu8ZRc13yDORcintieDbmgMd/
UJ+1ia9hZqPkNi5gIHWBYe7kL1Ig9+6eGEPAF/mGH9oTp7OGOh1P3WRA+4zJCrvZ
AnFIoY+5zq+FMZphQfYnm6rp5FYPaZRWa8LE1djEJt3E3ZZEfgmMQK4Yi4ElyIwg
DBZIh/H6Kk7mgrnFFHh0xYG8SHsYiNyA6giMfdYvm93tRTzVw/sQ5rLL0bhmAgac
2G/bwXDrC0d89HITBPPyxeUR10jheDi3ptAFPSURPVty9kOgauTlR8cZm8hhfrnM
5zwnt1d/gu/c15hfxUL1n/IUgANgc1vuAu7GXnlsyiD9HGCKgqy/Sy7txUvuxBCc
wCtU2kEq34VbN4kS1VKFoo2HRRRXPW6bVxLvwffoNvckUScv0/iycjZZHNvXWukj
H5QFur7Cwrf+c1YsSCRLyMWPRt5TtgPWSoeI+c4MKQfkI9NVHTkhLSOvXCVkNbGz
V8hBoWiUSeFaHfv8qCAhbvsuqnJNT678pUiIrrNKwlhSq70z7U4uDvnIiIq4PXXM
B+uwB2gWo+Oyw88EWS3BWybtrCiUxv4PNICsMe366WYDwr8z/ZuY2T612XZAsdDo
61fEuJuFdi+Se+MsNSNH8P5vvxABGYb+C10Utz4p6VfBasXx3gpuN7XE0kjrNmAR
nirst376NosIvQkjLCJFt5qe9k0lJKijmoDmnaOAfEjyrVbTZwrH/ZhxgO753KeD
7tnpAUIW2/DaBH+MgdCYDSU5TrRh1hUEOIoafSFvbFZl5QRI3qDo5MYW20Wurf92
FQBt5ZL1XTqZ6Oiu0ykOZGyIpP+XeQ0bzjcxS+Pj3YDwf8koRWwJKuqhou3JY6cr
ZNwPTqaUmoJ4Zy10rnPFltV6vnTERJq7Yc14GGvviAYNR7Vb6iv+iZW2dFA5v9cj
5ECg8LDeClnRAvG7pv9KI39edJsuDpz1NuGf/uw1Hg7TRoS/XrErTqWf2RmaCAD/
6PyCFa/xPu++VJ+/t/auQ0lDg5jtLb+bsjESNbZNfWpJCih2hYHoO9LI2mft/6En
9svxm3xxlisZHn9P9DzEXQTm9l7NwuMPRnXjBpfwKqyL8AIbTyjjhPP/GRyckgv0
yYUWUiNIJGXHKWWgw9zLASP+Y5mhYFmYUclld0dph0/UN+yFboTK8tXcfGM+hd7N
nEIHEthGmOz0E8BnVPx7WkA5+YrvdvtzXeF2udv1qWrcx4Jb+ePB5kZyJ+xMN60w
Wn2Z/V5tM9Ak9Wzepp8RGJe85JvAZbnxplhWt4YG/SjqVvsiWH9SVWzbMJ3jnj7d
d5Xr52RTDxGzlQDcnOYxWFbc0WYhSj4hjqAMnIEM6D9ixOF9hennPmPUVlQOW4nG
Col4U92PWu7cYjJexQzbHZM30k9MHiANvid3dQdWfSmUKfbybkZ1P1R7iuUOJqh9
3wAoIxWl5FxsT9zgvI1Hh5EU8fCGwIoiOT4oRQKzqiYmxHFCKtBQYBUcf47m5MD6
m/LWScxXkNxKd0wwEnT4ST/poJHDywTZOX+Gcn7fORFy2RVjQpKwrg0SOOa9GWqs
/uQeSU0YgiXwIeR9a1KyFDqNPQzLlSfXM21zdnHAVByYpViITCfOTa/N4TNoosNt
7AAdeepy5/nuVBd4tb+oOuuZtkr7HmmTgToiEOZ8QqA2y0M3pJ3ZFWCsC5CzFc9e
Csoxucg76sXSkyLBtmxwomERvePJtEsXCxLFaxHBpKDsXWJ2fLXA/T410uRYt32g
cgWplGyyzofgm7CYdbN6Nvsv8WEQ/ivcgWgmFWEkWgMpIDa9LsTV8x6/npQ1A1Ud
W1PuX3n7YTL8RbI4b0mYh/QM/OE90nC2JmP+czXe0Mc4oBXza4p+26s5l0QvWEt2
WbdaOPVGG1BF4j5owSQ+evMhRWJYD9RnIU5Nn9ZjG/CP9AW5UUHwd80fEtkO9+jt
lsYYpFh5DdPhtjNE22rmn0aR/BHH+ACWUNbtLtqmv/b/IvAm6UU8AfQtUONxreaT
CTQ5mHIqj385bPPXh9Ma7DwH5t7q7phVOg6fYJFJgaLPpOIz9Awlwz09kJnekORs
HYzn2zbzbE486THmstGuyJu7UaYtxptPOJEYp7hy3SRNNI2alFrN66Ule/cBUdVM
qm0hU+S4khbhpgBDTiJl5R3FqUz4/N3suwYSEJl6ckgHAN0BL4tLY9+mpjlAZhM2
xO2SIbNjnhxlKNEq9XFCP6C+ioCC0aDJs9Blem64gHoWMEvwoSBwU36x+aGTn1yF
gvFva9ARt0qrrFcRtstSeOtpZseBskxUO2mVca3Bn6UcVnx4GzAtrNo7GQ6gBwbA
uirEJCgm+4pLazAiNTvdTTydAfp6xiFMsg2oS/ybR86K9RNt8TlHeF4x8IGKsTgd
KYl0vpWubBb+3GYinPmp/phS/nN9kq/sBWhNTSKcDX5jczOEjHFOGhAVaA70qpGA
l+Bt2+WdeL8BpbchzZHAQLliaJ/CIh64Z2ynmkVFn5tzPxijr1eZhDpAWDcexvE1
6/vG7fuENlbkxVx+OKWvBXQgAujX/pCfDYFwY9KHJtB3RX926O1diWkQ3zDVHDfM
eGjgvx3qIpIhMXJA4/m/fkOCevDuB7cV7RSS2Uc2QcrDunnsMXGKPvEWIVkIfdJq
A3sbTCr52CgLJvMbZRcyQ3H/BWyGFoyTKPVJ6Gq4mHcG7aS7CY1aOc71+IWk6Fyl
K4c1zvgBVIleekxGNu3hzqx2LzB7SCcRu08J+gx7dsj77bC5K1lClFFIjTaR1FdI
y6iZ/YJVCfbn40C575ZJip/D4tDkf5cswbfsmhUrBKMtmZVtPLzECiuzSJOD6LqF
7sd2EbUuoJqrZPqq9iMaXfsXyk2bHM+7YznzgJ4+luHUJ3uQFjabS+kCTprCuxIT
OcBsxCpdUqfwa9UgNG/JfpRwKgh/ZZ4ky3TMPph0CAgpv3wlSxWqI9sLh08AqzF+
XLgE79f4yA2hUvSbrBxOf7De4pMGAmHma5z4ikRnfp/zWXEjL+ruvvlxxHlTI9ij
I+J+xjHClTIVbLTQfDMuulPM0WbZ41ehQV6frU/dX7dxGMh53ntvUTqtIwzL/RvV
WKQq2NU/dlTwtOfOBMndrGTvlc2oG+I49lDkNp+tOnbV0dtxa1pJmSQq1xpFvNRm
SQXEdWON8kDE16b+WlaIeSpae+qatCPMQ1kR9ktnIL3ZEr3a+HhnqrO+SPXmkqWF
0PgbGPUSBJt5LGz+zcpL0DmuW1nEtXfqfyZWGDxwa4MNryeHRXEZ5wnvzuH7LR16
1BOl2d5NFqBD+haV/ZNHuHXbNv/pcrMY/1AMOqD9CpVyWd4xDuB4ry5/AJzoDHW7
PKn7PP53VeiWPn/wbm/Nqncm1JCDGr37wCUPdw4x+LbkPe6JohYiIfpYRNI6SVpS
N+3cdWgR6AWqrzaLEcVz+gwEVvZNU+CQ6G7BwovyizlH3O6eU1PtWfDIx3a+k6pZ
2ayAptYZPB8A0loe7j7YcFJLvFiZqk1kyoZFIhKpXywiVjqYq04fMRsWkb+GwdJ6
RstsU4oTWXeZjFsKAczpjgQ53M/Cw24EBd9QjREp4RKOSEQ+ch7qe20avRDs71i0
Vm8/di49eNusa4Bqlb4/MWKmjlytYRLLrU20svH4SfjUqZC+Fqmimrfu7mW7uHLA
TqOO3R321wltLoLgDTIATvg502kmReYiGCO7qc9MEXZu1Vrq2sFmTLyuEkZk1Hrt
MWGGrA+gtbgC/UZG5uPqYNK9YW34PBS4r5P2SWSWj+dzp+ppgvN0UqJk8J6vRk+c
E1cQzkmtzekB1Wh0c1xyUM6aZzVBOoCjA+ypwKKUrq6RuodsFz+Jp9IrIGRYXwoT
80JyxvK6XVw9JKCYOgOCyyF2a9siQkZWKZ5mBOYGz3kb8nCgiG0wGD6kZTHSwCAR
Un27GM/mAFD5MLFxb9nLjk5c3f8bEz0IGEdz/rPp1GTcaR9gkuEiz7lqjgzfW2IJ
6h5VS4sK0RO4WI+zG2NxjnqBAPFvMQKEuF5ErxrCa9RZu4cInEH8NOota7ek+A4M
/BxdAOw78Hq88OFQ545sQnwDmI1OuhtCb5R+YJpmRf0u0ynadssrs1ueypYC9nzP
eI6zKUKZPx6EQYumWcR05WQ8X8C8v34EwOmSk3ct7rioPITB830hBa8Mxz7RxFEZ
O3p+9ggSCl/VIfYy8Y8VZ7xKyC9TcAO4p1RUpexl9EzYFxFwOTydnBSnk/Z8TTii
qVQ/kx/O9ZD6zgnHbCDgeiR/USuoCI2NFg5nDEWmaRNNpaUNcQ8eo3li88LnTYLO
lPVxzxH3eJxxrQsP+QIzYLJxEf0J6mmQ2/dcSsW4RUWONi8ltiuqY6goivK4056k
+wgkdGIPqq9+YUGcYxOa2kOuQCEa7a7aYa7ZyfrEuT9uCZMjoF73QZtrUp3soKNY
gxMlwMozHlw4VXr+KLsdZ/SVauzcJZ+eRjXm26jchcXmvbxhj/51jCkPaHFPnsf3
u2/lX0T5oac9cL2N0kkiCV4W3wA2t5j57yUTyCGVv4ulLvVBeGAm/UvDJ3FiBUY8
x/pdu7KGVpc35wRjfzqq1HoRzB74VtL07PqJsVpUMvcjP+1JfdrTawNtGcE7EIq2
utxPhL3ZgI/vWksND9ACb1AK/km8wuFA61NIpR2ktEYRCbE82eLXVT9hUm2fRanN
tIJexM55XJWOy/Rnk6Cp8amjPt/tTFABNpMHibAprLASCHp6qWDX07+aiXl+wrfv
OCeHu4QukOCRPCiIISU/YZt5OrrZZ2/6YQxDV0Qt9FVW1qMdnkIG2xERdivS/lVN
h7Ib6e8jRbKDAxt13HUitgFSlOHEq6LjRCqX2J2ya3dqWkGsF5Kt0Vz7xsu8z/4C
s1uV9rxF5Q4/s6GXGFsVNxzOrmCCCqnTNkrE4SL1CGYFxPBHqnq1O4GkU2R/QcmS
HeWXYyiieNi875t4uJIrUTBmON51jK70kehyeaUVOKxVnFgHRdB9YN5NHkfP4I6o
H2Q3cumlLmwK4+DuC0+aOjWqIT6ySXDZPkog9Vryaq0K209ViqtUJm6PC/ioyQTZ
bYcajcbI117lQpw6lp86eEgzQ2fbpQs/MRi4E0IWcbUTXUv02nOgDVCC8GujoZvY
i8XlsQmUEsQHv3RLSagmpBFQknuU/ZnBQ/VR7Qx0apI39fFR8njS/LBI+Cnp9Jj4
yBlJhVTOm2KJDzgO+O6E8SEupS41osvdkL5gYcZv8N/CGkzvIdu0lHIvFudUnoE9
3mL7qdHMJ8UiF+PCTp57+3oJVDD3Iph7KQIE1AkoN4g7YOG1L56Lb74Y0KCulBWI
l/04Uxp4uGvOcr4BaxlQSFOtDUeEsb99x6oneM86qe2vCjxnaOkLFLljn6fkf3Te
RKUWht/q2p701ExHF7akxQegBye42oPkhh6cJFq6P19YEEsfnY+2Ar40mtc/5z0X
hXf1YnkdP2DckT3XGVRycYx5HBZ+Q1XaIESWQ6MDDT3iRI+fJKvjCFu47NtRP7tr
lH4XcDQxju0v1JaBhouf6F9zL9zZyLt0UoDcyP5DyVuvlsAPIq1papRVL39aKx9B
KmLT0GnwGmkW4WS+89nNjDga/8OuYC8u7jIXbPOrn3Va6/rbwrXB+Tbei1r935qq
UXEBIBddEstF46xhJa9TlhdcFBnFhq+eQLRi3jOl4v6te74GVzS63nzZB7mcIv7I
7ElaXHIfCHcEblNCMyfqBIAxsmHKvYerKSAbNSYR5VpwLKaWfbeM+pgUZU7HVaev
aNiOds9UjclSVwvJet4gNUHGHugxNa/h+tCtFKRh7VZV9dbKFaco3tRfuKV06X7a
+cs/JzsCC6Z6agcSN/HKUIUTPo8HzzLt7Gk3To1XzpjJZJUxINyAX3eAA/UCbEId
0gZ5st1UzqqlOp/Kvd3Bnlh+5rbvD87VGyTqJxvCnte/pcNU2dHuQHjJEjqfo1qw
lsq04p6gxSgDTjaMYoecbQl+EPCwKCN6lS/1fdHP8nISRDHZtkCrx9WgOIhvHwkP
23DYyWzWH8G6TsXqQopB9zuj6wqIB+63RLKjifX8pFB2omeAT2zv2KoMlgwblC5n
3Ow93OteYGtMS5enBxZ1q5Gj03G+LdUKjY1wtK9no5II/4RwyIH/dOCWFKuBQflT
DR5Y74uPfXMbFvFv/NhDIGX5GFErGVEtQHgm0PpE8IuJhnb4wT53/iOJ/F7d1LT/
zGIiojjmFYS3fRLoGOJ2EZzi75k48mgPipJTydbzrrIVN7nJi2wb7mC4wfZYRaXh
YV/QFfcroaME6xiyXcWObh5DzQ7AmCd+DM0gjDl+fV86ed+lEoo17IBQ6G0BwibV
9ZjDgM247wsrWUpchHbzZPxa/aB/JflILQUQZGdyleev+ZMmeq/lYRfEy82kLlck
GdETcMYiKZmYYjgukuR0Pum7e8kvDgmxAmkuXFhtl0Dm8Fk4MNlyD3OAOYesLAK1
c/tUYxtgc684tdcRQ2C/5H8b/6YBQZiPyiLA7Cu1lO5O3nu4d4BTslo4px0sG1Tl
r3WVlzgo+UOJufRlSF7jrmVKwaL/wk6miba3dg9MWwa0Kuct+padlv0InmFvsONe
7moErzk7RM0f5VXuylFE9TZgjL2loq+uBmmx8Bjy1VdK6CrnC6pVrhdJIM0ZhsD7
uVxXAJjUoFg8xolib5r8eUdhMQgDX3Klbh/Cn6Op1T91lYC6gAICP/Co7G7ODDMl
tCk/eDe8KazIUWqHcnNpVZ78Xa1g/r7LMgeiQ4EWwOd8ydPdc22nDBDDITmNFpxc
mMvWWbRqQZd1izh6DvBE1f83YaV74ybfufVQp9nunm3Vr9sYUe9bkhM/i1S6xOxr
CHZA/GJfiMadUjSSKIp4RqOJcsLGpWP6unc7HE5WfHxogWGAkVGZjrwOZWxnt2OJ
asZV89gCfRTZSfHcGsBq11M9lC8vS0nenMj2P70AUdE389mF3UqED67aOesnRk71
uCqefFinLpTt5tMxVsTOWbelktyhJY3YEZ/mOtqmcFxPjueTTVg9flW6eSHk0DcN
YchrhoBinj4tQFVBCnI6+wIC+WPL276CuOCH8+exIOZaBiTXqdmO080MPqOZxohK
zbCB5MsUgQAovpZwnaTmJ7ZrqsN9QKKvPNln+0ACS1fx5sn+etTfe9q3+9abGRjH
uQnGcISoOKWBqp4KHjOrWb/JSJoLq7Ak6HPukF4XHICjIgdW5OTGXVul1yLPylXZ
FsyM+F9OAGv5g9uPgJNFZDfuDCK4nHS+cXqbyyoSi5VpelwNdCj5nlFNXWl5B1fZ
49gip62QJhBRXsbykkX/ju5M+S/Jbvh7nGm3ncVNk3/L39TkvFN8205OrdpRh7Ka
8DdoDp3IdHRbbD0iKxpQfb5dDFpTdD0suy5lPK4lVfeUccqpF4ZmXDvUofG6zjHR
GBA2LTS8loga/awRrD0tk7XogeWesMdeYUIbS5YC4MEme0El3r7pqwE1RurntXGs
gR+cFYgdCZ3H/aAJWfpmy79g0L0KPlapysjksWQmDhuiqmJv9Cg/fJcn6jvVIqcq
eehOADV4YRhmDEAESXu7Bq4X5xQq1FR42ya+Rk2E18k5P8rxms2inY6hINaaiOSI
AMps0xkoExF3sqfTM+73vlx026CVYjFAbNarDO31407f6FFNMcuqSqN25C5OAC8a
3XOV1cYaYILW/yUdHC0VlOEQv0mkrd0IInra1hnoKTazbJa6TEimzNZu8FAhBZyy
k2TBKEjRJgsph1IPWhQTPb7hzKUYSA2q4ZW39Phn8D4xes4h4VYfCbbySCLr6FbX
1xY8zRWOy4eOprq0R+78KMcr7kUGNd4dBDVeMGPFDU/G5A8ExZbGc0cbLwYw/7Wx
ZAam4ZEZ2ZxQmH67q0TMHei5EEpitXndsIWlelSu8gMufuj34wffAE6DtV5rBnJ7
EQQo0Tc//vqSscbnHh8nmHeZ2s8MmVpN8LvQ7vT0qnTK2Dmt9TWYqFLCi8koI1jo
VIJ+p8aedD0XJLAlJtjUgTsaMnsPsyD6awBr3DD3WZ5Zd7p1jKzGex5QrZT4tCFB
N4Z2QpjLR4Jw/omWZqGrmWnCKUsm5BvkmWX7m4iG6kmuv4OB75HHwfpcmIEaN63u
P2KDmF8ERVAA0ri94f6GtSEYx1j6F1VSXXjURGmOa8xTHhqf0pTHiFxF4FZPq15Z
YlSmvuLT2igkqPNi74Quqx+0BSNWzOk6Oltq97XstEUdl831ipynnlc2T4Bz98LF
81Tx7qJv9Do9Lg5MyNGhNIxNeHlQ6Bygi73gzWm7hEK14YfRRj8VJKmHJqd40E/b
QlmQRbWY/J6moLdDZn9S4oxsrFNbdA7hDPuhLJfS0vWIr9bnyxtQNlrL5Ar2NvGs
oPNmQsT3SlwvNmDz7YC3owMcu/reYn3N/m78QURYd4jN4tw1O0VshUpuCn/ZoYcK
yUZdgmsZRxDBVA+ykpci7pthitlee5BPRV18i00VOvvbna/lqIeLbcNEWyVvNE12
3toI8bnoT23jI9qOXND6a2oS9xA96WsomQhfX537vsLBIofVthvlKIfG6or3KSNf
VPuYhY1o1d8qXbmwfU7cS6cDZ+gKAui875AGplkWjPY/89E6CalSA2j88LY15/2Q
Fd600CloEiNQ7XNFdcdKoLK5Eb7qMthTH5KBTyW4+LYAh8Fwp0mz49tIeV5KyqNi
JunlTsN6ZfH9r2tkErfz3frZnYbHsHEAIIqToF2BmfXnGdml/gAAFfE8orcX74Fb
/vlhB3rpSLuVfSYvLv/nuVeikfvzMZ7dB8h59eMjYqi110qCXoo2tOc5Tvi0gA6v
dtCVcEOloZqTn3f4FS/h6Ade3ZXRLBE2ZgNbCj83McxhOeLUsHeeMdacVL7G/UIh
IJoXRTrJ1FyYfBT4CUm+zJuZRPfG+Cb8jKaTOjvwlDpqWXySTie/nbIqSCZB/rpd
BaVFSooQi7LtP7ZL6smR8WRyrxYCjA96sy0ks7WlNJ9SB1cARKp9bZkpvXz4i8T3
9houOHpRnVLk5o+nsJU8briigOUZTqa7CG5SAkjnV4w12kVhlZgemfQR+i/iA17q
3rqmVbnOw2PWEQdCtwjrpYxzeu41d2xNcjzYSY7KvLe0u+xOtQGx66b+CAih7fSX
KwPBtiCGM1afMg694uiavnY8qoihal0s7CTX9gManUIxeuv7Y8O/stxQFQdHcgVO
uRSD93N5lomIcHsB4FkKObHbxWYrG92vrp4HL5yx7LZwgykTY2dsyD9CarZCuyGP
FNh31l2eqUJeHUj1fqlpKU7/B6TNx+cl8ZnST1KK/K+4CVzY7IwN5Vige9dHvLoB
/+WBANLqG7mDg0RadSUsZsa/5fxq9FjiwYzxGFbo+NkMKoPZ1Gvlbuq+tuH4SU0w
XaikXxS797gKHBW+hpvBKz7EYBhxNvCPXrtPLGVvcj+CyFHUUtfa9hz5OjEwgsMB
LdgZJJ477sGGIlIJ4B3mRdCZn+9YJ5fzqwqj+r4ImZ+kdIs/46g5CIcPsg3eSeCm
CVd5H8rEKbRIfROyVHWfqncAGOcQdnyGmaiWBp7fHk4fEEewqry5iEFMhzPAeNaA
rtn5NXG/NCNWPl09/Zj1VWkD7nhTjVSGgHla/Hyh0llrYr399zqowEEXNWgaHQNX
yXqMOuCIy7/ew0yCzOyDhWYf4vJlhaY+/DikRr+2LNRITbDTh7kI/WE6DpERmo4v
3IgnrFvgTPOi4fi32DFLyXLITWyCPM5uIRQSF41husnbQpf1rZ/GrENll+hfPXSc
W7XadwpLumV9sgNRVekzKGc7aoWLXWs5xTDmRvmKFdpGExQgx+QxnZiudjCgXJAD
S+9prGgFHOUx0t6tMGtaUYfNg5DaxTwReS5il83YUa+xMBRiX/X9RcfDpRewLoKB
w7wystUWF/iQi77C0leLEQfuwlPipc4CLy+53YbKMqGlQ1GPPVMvSedARw9VGngZ
GAoDiGCGh+nS1/tg/fmZ9zI3y3cjtmpYAdSGgAo8gZoIBV4sfJXriecSX5rOUtYy
TW9naaO1H8e19cOWyCAeg8ws/Vz07wzma0ObhfnkcawDSRQoiX09Ypx0STxgCO0f
iGGs2HmiBbbKA0tKV3L46YVLMJJMpgPU3BaO3vB8V6gFl0R5pIXeeWQPMTN8T4+G
zRD3psSIZX8wAk26eXwViu9kzO1QyZG3VU+WEzUtysQ3Fjf5LP9FHr48svl3AcUn
b18/9alJxmXSBSs8fcEofUxdTzZuANJz/m2VAskh69At3jILY3MPeTey5H6bZOfd
K4IpKbpwNQThHfRDZugYQEWYRd+zFTpf9HJ7NzqW289TX6HPfmk43k7s1RHrRZIi
tggPKKUJAScm/AUq6fmiqXbe/Hx0aBcNCr8LdJGpmarng9514bK5aCESfHHrTK6x
CqDy6JWq/KMZxd2qleLbvN+z2N/OXowipMjEqLIz9BzXxmk6pTs4wzYILzmG50bC
y9ZbJwEeZ8EWD1ok0sIvSLvzaZhRyO+MflsOzY5NwxDf5jtoOs3riwI7ElnUQNDc
cj8KbY7XcY/NQMv7tiVo7Ym4GveC9T8iqlXKNvjwDYE78SWSiOcmbzsOq72ECqnJ
wAPfLvcdGlBBi0Us4/BAnhZWe1z1rs+YvHT0sCOl0h8/Mn/sR63F2K+OV4Cb3rS5
6r8GyEUp0vasjJ4G4hlZiLRbu7G8uiNgjDPjHWdB50ZjaRXMMJDsjuIvgW8tjCQx
e/JKetvhlEdYeCW8IQLZ9J3FYp5Rozsr/6Az1awcX6H1LeDiP4IiLLC0tbcOigOW
jqSjo5eSOV04XQp5rVgOEDhR7xf/pH99yvHcTBRWgPvIe4W/WcgZ2mm5thT1A7CF
hVSrP3674iTmWW5LrNXoKeiF6g80L4PkITV/ku4XSOVfAiiOddMjAJ5TVrvzCM7k
4jaHWxcRowidgsL/u11HjqfVtYlZJO2krQSaOB02N79dkORW2lL+7fcGHNMR2dzc
2bRNR06k6ncwtb5nQWIEfT59VwXSiSRbHgKB5Df/BX/WgGPK414n019e24UXYaSk
77CWE6l81UYPYMk9tZl9u9ALEk4nZitUmK1+RaEcjBfnQTgGetEoJ2HMeWnBwaAv
/UrtZaApA9fzQAbU24D5n29lTPjFt4J5eDo4CvJH2uj1/Qv9cFSWa80BIwxmyNWD
/duACblZQ1izLGzmm93al4Dh27hJ8dmUA48ss3rhP5vzbzaTCvOjI9DN5HfWzOuU
gRDHhGbD+cTvw2dEVtThlDdmruLFRHFv08PR3ncGeITRJJ2yvSGpZktUF5pSEn6n
Cb7ufy6+ptcLDg5cO9qU7UCso7eh8XzYK9z+tRXM0XdpvheyjUmNNgbWGXLJFxS/
Ando73VwKcYluZhDQOnd1eiaeA8N+ycEAGYA1le+3TfST6wMoqjzU6/mv1q+iNMf
BMERFALTBDLrXKv6MUvLbDjCC6gKn4aL76M1Nn9p/ozGDTggNdJieuCdwIeH8Lsm
bMa0QQqmNoYFxd+abQRx7jG1kJF9077pAaQ+0E0ydgIS3NAZBlcU3m7iFPPBmf+k
QMwn7MWhCpswfREN4/cAkiKAIpUIj0YkgyovOEy6wlKLcKRPZgeVqXWO7LRflKtz
7GLsUVK7S7KvpHVVm/E+z4Bd9R/1UTm7HCA70WBh8wJs7S4KlC4IGNgY9CQQmMLo
/SwHTUwIqHooCncf7Xl2UOGwAhnHwuy543U8z2a7lJzRNanPzN2R8JLPzZK7LZkp
uisG9hJIa4eNUWdAwssEn0iMGTSunDbgLjrZGeZJzACrrWIzicTYJJJHt3MHRCpP
X5oelug+6WnYUF436kL0OTvTptKisSmnFViCnwx2phkW1MkyWi8Shh5D4aAuvhya
aYTZHun+v/IzMx3QJe03vmL6WAV8r8Ks3NYHP+c1Fy2RwvdmmMc5EdmB/btYTnI3
WP5NwsPoLdCYYctakYqDZZCt2/yQLWRaBGLfKS8fR0wP3kFxPIhISH9LiadL5Mmi
FO96+Z2ggmVtYxbTlpGaC25Zti3ncytsBGwDL6h/B5Te8yoBhrud1aCeNdno1WlB
BNenfN5dpbJlMbWlHHtCK7rlBSUUu526FnXBMVsx/eD791gz5zmZln8ioiH05+F/
d7LlMbteDJE5sCO04PLO5SPtLamYLpVJdvY9UgZmdZGruFNzQxKUoSGsvpWRuKcC
BeJEo3aUBm4bAjzzruC/Ryx2cB3dO98gpxule+bgf9NztEx4xpVpnBSTqKjD/xQB
Es0AQ5xJnH+EUPIot05HNVCbdLICSb6EMMiuxeYwcNjWTjDbraF/G/l2TeC+pmfq
NO2eRIHVh2Q5B6NEt9x955u3DWmoIM+8AZQn6ffdQUMcRc8d4efKVAFDBknh9bSp
V6ZFkoMged7wojla8iTL0Mt048fRtY+M80TZim2rt3Z1lh3soU3svJwlVdQ+ZuS1
PByYZY9k+DKVvV9v4cT8wqiZMq5pUqYP32qGQvUOiAzqpKrxru7J4vw9Dk2vDS6f
S6/+LdYz6y/2mER0VPPRZ7Qn3JkjQKCJyDKY1jTduySh/tm4vh+4ehuTVHtdMJIG
DCQwhgDN5C8kKP8lUW5+tmFxUW+JBUnBRpaVUuZb59u4jidtXBBgQSQc3zmtd3Pt
7InNlocqrblTdgcQVzE9RJQIUkjz1uNHGeF9jtQBGVQyJuWhbqpNZRUtohf1oeXn
Y//p0Za4dHoak754HeRknKurDT60FKDD26Zulzh4upceCnjI8WEcZtGwYms4GnMx
tgZOShXRk+rMe02xyUgK8ym1Ev8eecyWO2bXDaZTIcBWpCVqPaLhsJE4E/aTgBmE
GIbTHkQ8zmkKvZRCqkRmsuMNY/F9uTbpVF/RZDYrae+0kc2ugxb9YFes3QafExgu
wJ4qTxLkxeIKr40KQNhKTYeDI1lbAGFxfX18HBuesgOOzV93J2YP1s/oDIpmmKDe
8OuOJU3KOCwMmkxx67qY3YwQImjqQXMBzN3LDSRitZW0QKuDdambtKXJSbl/3AbU
NkP6iJaZl6pjhIN2l4NQSrDneM+ct9LsG8MAr88+YXTrvgjgkjXlgIOtIMoKIruX
Ue4MQ07yog6xXKpsM1d/JM/CL8bgyelZmAqviqv2x59667gTNTfv7P872FSOmqcK
uTzBXxBrbKqD31h3l1sOUUjbTL6wdK6GnBCnA/PYkhRGpsFpXG9wLo1hstsvLkPW
y5m98nni0XSqr99uXRMZ9j710TrrdOTSxGK5raQNjt9tdH9NQuknSdI+MmIl2+cP
qWUhq9bZgWm+ZLIGvOEn+nkKRCZ27yFH/rYkgEfWN4U9xvIWGh6upnp6R8tshuhO
ScIMt7HgQfAzeOT7UcC8BDmQg7MDWWBl+YUlKM3nPiCPXZpYYVVvMxLwQz0TLGCO
8DNc/136pM3RAcC+tg+nEn3R3nkzMcgsfRY/8NkkcN1Fhtm02s6pgPG79owfJ7o3
dbhjVAohIS7yApXtFiH5UWzFcOUWCHf8nasMYsTpRwt65WTVyKNHGen+60+o+Xiw
yUBqFL7tVAenwtPZqXWDed3xqP6j4BrI25EcuXiLPOq37gQD4lfsizy/tpbPQt87
Zofujoi7C3HoAomeCyEw+uVCFlUiHKXwPRWfNXJXzwK6bCDdYi7Ljq4bURrUAd56
x5oC9za7a8v/HwBgW5kz50UalfurAeCiltP+It+qloURCDEU9ZYiW52kUP93QsS8
cH8v74wllI+j0bwv0/pNuiIIwLEXM6HNUzQwUCuiFWpTVy9Y7mERUvBYyPcqTxhd
1nCnCcuTIAMi5m4UaNNtfJo8SdnKBDTG0ze5vxYFXHtwaXkchJ3B/TgihfX3zdzu
AuEEvtm1/RfxayAF2+vzhM2O6G7br+M9TH8AAcE8yXxq1j+iTYirg8aRFN02GyBB
yHYzX5b6nBjAT7OG3WlZXW2sEwgS7m+7dtLEED5ZmYuCfDqeHv7Ob9eb+vtoQ/IU
xQ1AksZ/aDpsDW+Ppl3yzq6tVZezsLW/eV1BX/nDSJUweXjBLBTwz0iYUKxgz03O
bcAXPoIeLQCeuGWDJAEwCGL8kj2pH6n26gygCvqJZY4tBmHF3fK6dyLTj8gC6TkA
6+YYbl06InC32EyNLhDyT0Q8mOPhfA0xHGUGOBlW9yc9+zjBOjfvRxUtMesJ+XXi
/g90VRWRLpReNk9Tnn2elUdQB22CV8MfktO01K18tXxD4GKpGXru8gggp/OzQyDP
KVh++Y+kdpEsYAM1epqIufH9unMSsumJGqLK1tqQoXTZIrrH6dkAWjyK20Ex1UwU
q1hcN2KUzTytyhSpHV3duZPMun/pr8kmnCSx+SyzB/F1+RJ+N3MZVwK+iZANaiuA
k4rEIEWPeUR2NXGpgK1iIP8GX/CY8eOPnDHL3PWW0KsnCt0Ks5C8XLX3EYsHuywr
IKH8Wu5xF8RqWxKDEuEAlhw60kZrfS5gx0jK2GtFGLDIHoNuPabp4IOt3clM5mPh
2GNf1ioGCJN3IHpC4kgaJQgcoOXE9ld3h8D3Qf+bdcvTycJMQvhTbvp+1TMlJiX7
dO6NxwjIQ6xZUrMl/DySAFWdZ34BUqA87igTkguw7MHt2G+E7Vipn4pFK+ux8YCu
nPh6owZafn2tOIM4XeIfP4ic7Xg1WdV2Q8FnClp3VJ1NdEnsJLgkF7b38biNZfcw
4wT7tkvr3zg4Oxz5t0R34lWoeLeAQHFG2OmptGXT2/7c0Ryl9P8uaCLc74xUsdHi
D/o0EZQy561WN5ghYZ6TkVwsuJDVM4hj7Mqph4fxsV4Kq2S9u1MlVQ9u4IKAY91I
oq5K4v0lZr+mg0u++Laf5R0wcPt+/dX838UpMrM/kwvDGHAmlmQ5KlgMgSoYEPCP
mIykGS4ycmqEAxuA4zY7losU4JFFtlVkdjnkMEJxkPkE+gjaL660l8k8kAXvgTKq
m7kp0Ia/bo+BeIEgqesClF44rvhUShQ6GXbYKzE6cnAEij85kPArbZBv88j9HqXy
IgSIMmuCEMDDvXaXQqkAYHhmguIq01HCb5hhm35PN/7HY2512bQ6LX0uBPKV0mep
HHpjZynCIJCpXbryH2RGYeKUNNU4Ptj0biBF11Imt08fAZw2v27Bcob4BKZjrpXy
NhMRXWVzm30c7N+rOz82lN6mTL/rVmxxFmC22MKmMYR0FG6gH4oSTj7/ht5woQmg
hYll8g3G43E4xMgcNidH7DkDA/ETL/W+3CAx1bPParDMaNvD6hPG2wnTm0atAJbm
qfivfougjPzAWHSsoK8TvTALz+v/SFaLEgK/Y3c1CJ+gN4fzBd9Sh59ohDkSQKj5
iieG02j664v96LvRD4DzeB9ypmGhH768dOvxq+2CJfUPGtIfUJpEAW/2RfkONxHN
DmGzY1EmvRmr/xwiHURb44rctLa6WlugBw7BJGgywZ9I+1Geh74sg5DQsmF8p8ka
irBfttdva5SS7vMTUaZjSyXeO0Kw9HpeYE9g3AHXVrd2UKlgcTNWgugdSQt2laNl
/Kz1DYDK33vm/FnvpC/0QBlAwMnJBTh5aZuvH3W+2a8T+35A629Y0+jusU8wg7qQ
gPYiVyhtPDWAi7pSFgdh980bb5kuzzv6NYKWzm77xotkhBreDOT23XwLDCs83RYJ
rlrupFuz35nVi+tErdhp8wnJEuFXukEr+M83UwDEnkvcmmly/ERp4Bd4csMm43zA
5rv5OlCBNMLfejLvzU1GWSSiyr5txtgoc67VdHX1cKYcykDPACT6lXaUPXHhSiqq
WfIPRGxidfxjjzxZApR/9khBIqxgUJBXVkPJ8DnfslNmhDQIEMnVoSd42AkDsZB0
t+19oDnwTTO45rPWo1ZcMM2BEl7jQUpwkNk3M1FC2utDuBRojhtsYrnXpX9LzQQZ
Op+YHJiuGGVBspWwTlX04SMRsopNIMJfLbZ75V0hpnGM6cxgRtOYhVcQJsPsgDr/
Ep03J4Bx2QD9FtAoARAsOo9gTDO1Fqc2MCy/+R2ctgmrONG6JEFTQzT4bMJmLHmL
6ktJzZMtL5ZCQu+f/vIrkpz7hdocQO9Dqs7XVo+/vIOv6XYpFY7G18XAn64fCg6l
tl6f2WYY3aHCCgXEgH+kWeiCBKr4hymwu28PHhv0TZ5hh5w9PsgTmA3wAAd35A+l
fm/PSu1kmuFi2LsFKPr6EwV+yCQYZS6i0cQKHSUt9eKLZYDpCDIXDP+z/QkmFWjd
ZqgtrojSm65k7BpXjkYiY7AJOecXF4vRlohgUhbI0QDeV5Fr7KbrpkgYQ8NlK8MP
UxSynS4XAnZOJWsvDNjTPs5FPjIpwRl4zwTzNIGmp7JJH/fxxriML+ZhWqyO5e9r
i1Uf2rsXwkCpTEt51rXPeXKR/mdM5lfffGt6hc56d4Y3P8PZrCKy5D5hIp6rk8C9
Ps3zT7mL8h/jzFu/ST8Lg4lLcNoThnYl0rc12LEzC+RkYuUnWj+h/yJ5+3c9qyij
GajypXmy0J2L6AQ7Drp07/ab42WjJ7wV/CZ+5MgDuxVXe39nJ2siU8DtPu95hpxY
vHBmQXVmHuYD/1oAF/o3hVk4VASdDNHVzkin2e4Qp+sul9Iq5NtvhYOjvyexs6kX
cwmexqwDqraGGbtYRk4nilQSntA4k2eNehCO4W7HtX2iENaEB27vtBa5H8qlJtPI
8YcAXVfprPMJabDdeeKrW1VgVakX4s/W4mdOmUPwCjzwoLnUxdBiaNf9f4OpLOSl
nQirSbxiv0WAv8ibw5VGCCeH1JZGDkRR6sYtHrrs5u8Co1ou7y9sQcOC9c8UN9Ea
TSdz3ux8S1DbCshcOwMEm0YLJJYp3vsKng+LMJDyFjNXlFN56qVvvB9VsVsEg8jJ
WGshCnZsbKW4Fv4h1myR2mHAv8+9ODZccR6kbxv5sjxQ+dbYDY5AafCllSTCyWJI
E6Rxootd80Kx+1RWUGcQNwQ2sHZUvsfs05tCvhNefe/G6mOAIamr7MuPtnix4DBH
RVLqCDjHW3ekhq3o7iT2uAxtM6wSsIU5nlbVC/T2riUbUOgTaZV7Tc0V/nwbZLDl
8bDJggQ3nei9SXZNjfBw9kSQNeHkraKB70SgSm0wQhep2TmOwOinYDiaIdT9j+zs
KY2t2O1RaQdWikf4Cy0Lu3TFX5suUyIztFNielmGj+z5jG7qPyMMyp3+tYpucxON
gv0sjUu6oQ48G6EVxam63sDRWRH5llHy3+i2Nw4DyFfJo0PUP/H8lNhp4ziNKG50
mbF3Hk+5DKvGajjGWSY/QGG6BWx9zOcH8qKjIh3rQDVMEVfh1nEv6HI0mPlgwYYu
uEbggnxIpboityGrHAFyRpl+TWnSdxeXyBdg+jwWKBLqTkrtIpFVOjySmG3mgBYr
H51D0cqVArJKgM7DaKHpYKYrxB6DC72zLDR2Lm9MOYCbOnDnZcVMNZFzvWnWFXEY
ILkDYWWqMOlb7CbmlRqCMMVUilPTj5D3ztCux4Z+RZP5f79VPnWAOhwQSp8B1Kz/
LgsggPYdUeetdhgWBlDrFWVDFran3kdwQZOP7VmoECcJ7t3/sIZzdzsoZbwLqOAc
0XhucTORdgdKqeq2FBsqF7GyTXHXhOc7qFot12rkIMeHgZeXbtUFIgB0lRuRXE4e
FMEHRBn8vQgrDZctEkGR3+R6IqUgydlbnm/i2/I4wKAfbSOgWIQ2Gaaa42DyEI9W
Fzjcqi9NUwdJptlNC6NxxjX8PGHMUNmpBpWidltjxCwmDcVr4GFrudOjgLjn8jRs
rr/lPTySO/T+j8/N8WXRmjTjixtrYwgTIDcmpKsr7VcCRFg57bIbZfRRCr4GVkrc
aTRK58HxJKkaE1ax9jPeusR/rm8MSEeUI5Nmq2Dla+ruMigIcRZw+s3CQNmNEOBc
Xa7zosflfQUX+hlk6Q48OwY8Wukl+AJP48mx0lGCMP1LwnHnpggyBeyXep8+3myY
kRpJgD1CO3k9f7lb3A2JG+DbnzCRxTaXRaabgTkdVq+1U+TGkE8AWFkWfddbbcHh
eynP+c5gKUZ+fyEmXlNiMIyqVae1pDoKr7zSjKSETlfiX/OVZUDnPtMvf+tVHiXr
pNklnCzv4EUy+Lxh5BXK78z+dhd8JiYWqT7r2AWLCHBds1KFi8iftOGuHQUFRNIv
HXLzfAKHPMRVJw+u/h4dGkMiT9kJ7rt5YyZg9Y2YWiheT7Xbf2iO6KkaERLBaJp2
gv7cxzDwF2btEauza/qCV99gCTa8ydux6wL1hZJWJ0UCh/8PbJKk6BHPf02coWmM
3hl+HGsbeiC3HMRHRbsL7r1h2Ehrw8xbL1ZtwPoiCQNWeosizWbEjYCf1cwHUo6k
liW2Nv+1eOuUNZ6NS0BW6eRWYxp3YX8bfaRZaklvmUGBO92Wdnc/UV+BdH0SX4ny
zfFp2QoJV82g+LKUe4XnO/uDSL+y07eFg6q9DhSe+8+TskrxAgkjpUQpMg7h4KsI
xJ4vV0Q1n953F52pWx7v+QZuu+mGpgvqz4FJNwncVJdu2tx2XewJ2TMiOtUDxHwX
CzIV2p+ooE1q7hfGdZqv9kFpWTJoTCpUyrLiblRqTjhLTRNNfHP1lgmdAhxx6rtd
jufxqiPhxtRDV3s0Fsje7G7fJc1cCpc0v/JKjE6MyCXjYgV2xOSmdirflVDFWNHW
dLRAGVxmEShRN7mXeIrFmnHMhwEToVTZROAQpIcendRBIueoW4ZYtjmKFVBbbj30
yog8AmM3I64LQ6YvHlCPdzD2IJf0sxshgxNMQmupQAc4sqKIrK9AndOMjzoxwpYf
+CF0HKusZZdTul3SN/qqSwc2cTngPA/1B7CoFUT3gIIMQFBVaHjinY7fAuQUZ2Hb
hWe12Me9jDkXtuv0nL8CsApdxtSBXfKmSE0RAzw80HPsLtHgK0ykX9RYyW/Gh2G+
TvW39B6krm+lwgzJUbKN4QtEXWbI5Cr+wpPuuSbOJIoGVas1uFXkuHlPFn11jj5I
Dk+LU6TfC9XOAJHjxBo6cX+sn3pKsr+gcivP31DT6njXINrILEVcLpoPxeAkrbSZ
jSfxZv6DpAgjMiqytysVe1lNBiQWlA69EWcB1lf0xAwA8wJOQPjDAGONIjtvPaQb
Z29qC9/sYcFm900J314KrcmQCq4VBt199F51cbyKQGmbavV1A5SpmdPZ4KtLrqQN
yFfsL8ycWeR1IO7tr4cL+L1ezmDSOnMCgGtct9fCcqKrhkfoYxEgdsDK9tNKI5+Z
vxsP0A19HonvZfnJWpyj0QJctWL2IXWZ+xEVW8yUMgN6UkmiuPNusddwQPIaP9TA
nz6rgL1kU5k4TfceC3b7yIYv7xR+ifFzXFKWq6VtVvHedvQhusblIWlVDKAvh8rs
jmjMsO96oi5/LCS4IpzY1gvec2zUdEK1cILyN0stxMNLR35Y82isKHVgz0wI2Bnv
lM3OnK5ivQsjFZB2lR/Eqdv92L7i1KK5lAxhnEAwc7kf4zSZEfXbDhWdoat4xe70
taCMSWz/pK4y95LHtsY9KLGxn5gwVXTz/vZacv60H4awvJPesCrl+tkJCO6pLWX2
Hjk6zMuqUX7ngTuvzDFm6jlRcbAhTvsoVIFag/C8Mq1Q3w/QUXRwY405dBEtqFTU
RaoLF/k1Bj4GKgLYOoHGtVH+CFTn3bZ9C63/w6bMoHBnMAno+HXsUFgdidlaEXaB
zh9c9loskeEvg7OEcBy7WBQPLcYZsZGMr1rbcziXUHixLOMYpVRXX5VuTQPnkwF9
a+6zcAHEmpbXqp4W8sdi5shUzMr0VCKD5JJpJV5nstN/On57iWBWwSlS3J95+oLX
sfU3ox4Ntq4++DwdHtV1Krg94/BPdA1KXjrcemAwI53NkLyga/ANZf0heB/bml/d
ycXvVPeJgHe6MATL8bzJ9PcTxutTd4MN9Wb+ytXHxSH0n6VkP07eFYdff23SW6Lh
n/izUQ/6vqMEe2UzvyFbX8pMEpbpIWfzP6b/ypzK/KJe6IeHpRko7RAr4YZNCN/m
mKEHoQjCZBsHqYD9WFTlv9mlf57hdVpp0n3Wwtuy5SiO+sRn1sHtwnL9eoPwmxvD
44972GfR5e7VzdzB9SApugyoKXnLhm9Nj7NA6PVeIJIgRDTx23Eq8byeeLbZhWaU
igimSPBFN4sZ0jTLcRdmW4cJoJPum7ZNGtBFuCC0+sOVJl2YdTrAZpCkTrq80/Zr
HhU+OBYvqBL58wkWJ727tk+U0nAHdiIDy945GIsBAu23WCcYBwhzlU6K2c5OaVFA
WWX530nBVnudumNlIPRZRKtHgMgLEVkZY/30hGVQVT1ertkCtkT8fEbedyLhMjXT
9T8gpL72RZewleJZGvHeJVULM0VY0aznKtiNVATAd6Yl2M/YTth9A2IcPucInqNI
hp8TytULFraOryCnES9enhC4Ks/2R+cw69tHIknVrHuLb14WiUSehH3i5wRzwNCC
SqJyEFXsnyHqFMWM/z40icAplJrBFsGnPfIuzlXMVU51c/tbgkwE7pE+1jjidjg0
Jc4EFeON0h0ZII7mwB48Oug8cqv0m7nwtdS9Bk0JyH7cLTWADdKxZYpJ3a/wqoOW
UxVcqbBlhtmQw9tmmxK6Rk0Y7FcBaVkdF3E2XrybemPH1SqkQZdsi0XMoC5bPnRA
c8HhEgSJl+HrHl4zkT85uHunj7UJIAGe/84NMSoXUUz11IFbwdF0JFCpuhmshSUm
8+cx2pZ1e/l8wzf7vfVnD1XGIY1ISSgOQ1sU60W4y9yNUdwh/YRrN3SlrOgfHS5E
YVW9aQLceQoU+u9bOXzSCB85NMTXEtsNn66aVB64Z+3AWB7S8l8EXsqoaF2ct1kA
Jef0osHZodp8lQkXbD/r2LT1fZQ3TvScYd2Og5rfS9ZJ2fvqYdffDYlS6FgaLiV+
COiedgSlBMytnWM2Pqpm6w8ZkELAyZxwiwkNS+c0cRGNoTc7HCPdyzdZW404VGpR
ulyrhJB8uUaGxSHADfOR160kG32vf9rTkQWAtM0esOC8rDGEwUqqC+70h+BOkYPx
gWcEofN+Lk9gwn3tlBrt1/BEn6L4Gpxiv/HzDzQE1z2p73LbLa1loC7R1TG+kcVN
6DFfnURFU0Yljy57qeZKf063ddZklMCLFKmCHXD7emjRkxwb4MiA40Hwk+7pAbB2
YXqTgBneezyubJ6Du5edZgC5YO4M4DPEmQvOMJSYAPBBPYN9t/OhGovYzPdIZzJP
YRjxwb6BCwPRffl8rOd/j4nyIj+CIlpYggvJCTUe0g8js+WbAmCXOMDXDItra1M7
Gljv60mZRSCAowmCUiKRW930bxFVgU42tkUpDX37yU0101vrkNpuxKcbH4FuLEVD
2dGYTzEqLBJJ3iQy6lfZzdg9gi4dadZJH4GoPBU07G6TURExpj/t9absWP4La5Pf
zYqG9iEt9tC7+Un3JbWR5/VmeUhILheDNP5BOa4hMaYj2isOJrk1EvjVLqxNTNhy
hMbW6RtrDfXwEN6UUnvxugDhXegY6MlvDEcGItVQ/p56yVZYblleRPB2Fm0lX6Wy
MyI9ir1R19zv84/JZl+Wi679LDmOz5TTYnADzlRaNrnpS2ERUYGhQHiyuVguP+33
JTIc+BuCXV5GQaKnPJYZTFpsR/zXLjnF4wwDZhd166f9/FlXp7rQDJffXqjHc4lO
TXoIx/I4jsLQCof71e6lOy9d2J0XgK8B2C5Hjv43d6k6nKNmWLdukb9LcZx/Ez9Z
jrv6Dh6pQhVSfyzyMKAwP6bmgM530R+X3N1ULpibMe356D2sfTRMQRr5GqAkrikW
tHOm22gMdG1pnRFRnHfY3koUM3JUn2iv2U5Qs8vbrTx8L75yv/NfeK9MDl4ZlcN5
ghtNtCLM0sGJ4qCup34rcTvQ78cKpaTSv9arbbO4HuUEesBsFmn9lHkY+TsKFS3e
UgRWd9lV46Mqh/tQFVjxhTSLLg+Vthc0XQlTeDsCVzQ8l9aXcfCEdkei0BejeTRz
GiQw38i2dkC4SU//23bxE4YLv3cPSuDhoShvsVI+gqGloUJnEBSxAbQXazdhMu90
ORBtSHMVyfndisxFVeMsZ8rd+Je22Rxnvejf45MfXo8OnDmy0+nWdD5k6GaICUC7
YPML+ztOwuSGY5ZVSdCkEP4BHP0Ba2/19/7NlBVo5D2G/Me/dcYLpGUPNAJoZUK/
5AuxglcgfkN48q7MMlpYlSzn+Ut7cboEqc81jPvzFjlAhZmisxas9KFWAz6rDxi4
DZcLFXajM/qKVB0mn5G9GM0UcN9j2tDw41CBgfLY2jFQ477eWMdSWayStFqMMZx0
l2UCq2oXxHbG+t2gKt8QC9AHSgCPU5fT+B4flmDv7cdzPMIvq7dkfNz1ogLBZf3c
u2oBgmihMbu6+aFzVwl0kgTaXNiHD1XySBQ9IihF5V+cWOAkxS9jsdK/J52alyIu
pQ3u9JP/au204U0Zr76k0TxE0Pt0dnAKL6pAvghA385EdF8mvw32Tuz3wTF5cSJi
8RFAPWnHTpTlXQLc7mFQqZ0PcuENE7Cr3fBps1RhlPPL/FnsqBJUne5BWo1dW2BV
YAGGPl7dOS3EICKlrhaxiRQ0dCv6omMLY/ZYTbpRubqcfxvNyraf7cRUfjEAesCK
vAuLaSOwskyAYu3sE9pnnOw6QQ2Zbo4itIXEDcp3Kav753d64F9NBiFQu0NfIdqd
FEMtKUZ3y53lt2FpvG+mzjQA53uHxPU3Ks58xGndf7fdn9el0k3hhCVHSnKelIem
yhdUTzOqlw0X0kx8CqvTQV30yduTd/0zTAiU5uY4+YUrNlOzSUp9DSySbWAcTc4u
tTRB0+BJ1UvhDZgD0eQL+RffsH3w78b/EJ6XqVL9Y68O7K1LDO2KwnCT1+JwpOM7
ETpOdswOwLvS0yp9oKMaEbapKhVa9pM8jJBX360DEPhzWxMSFKnz46o9R9XD0tTb
4XnalVfnT49j56ychZJLLXSqUHVFb7h8mTb22k5hyAF73bN573nv2To5oDw4liCL
85WiuqPjtJqVqZZBMsR0gD4VhnQ5KRl27z2VOsHP6iUfYTBObQUsKNHU0mxsk96U
MoyQmrBq79/aK+r+Q03hBJPTz/7Usgv4pz+tXiqH/GMaASEaBtbmXSQtmgzAcqmz
+DDN7D6ClCCkC2ob999d4CCz+w+YDHR8yB717VJA7L/kBTVK5HKM6aMPzHL7I8Ei
wOna0Zj8bl1YyUqyRBs4ND2/H2+Qf+Fp2J29zw3MoGaO7N8fszhzvjjrTbj92V0t
1cCV/gsMvEow5XTBg0/7n74Za8PIyp6Raj9KDa2RV96dbH4GaQxH+wxo9txEzggw
0RwWaGJdPkm7wDh3+jKjjo0UgODxNOU3AjFxC/+/H3O6FoaIAnARBW3LLxxeKdom
WP6yBdAWUReOwJVoJdWhSn4EIqzT3xtT7A44+UkeaKtnDECmNW2jZUH7d1oRgrzH
KTi4sj4TVCDPf6m+RkkFdNXjBvYbodedH3y9WJfBTDNuK4rzLsWF0O0W7aq4C7Lp
b3xN/U8IOeL0Yr3EpRplFxHXRljLiCoBti2Q51WE5FjUk/pHOtkR22TnXUd6eIZG
mD2Dvw6u55Fu2Z8EJ9xo0+j2CtSlUU3Gp1yD2OMr+DahyQiWO11Zz8k4frKFJp2/
SovqolJQq0gsdZObbiImV5sC4IxFGsGuA9hJAmFtSYRr7VBK0I6ILlAhVgwoCUJV
qCfOZWbkCZ47ARnBOkib3Szp+k67lZBrPTPeQdGmjBRyXsZA1FhEXgMPNN7W6TTO
9DYykX2pOzLf/tAgjTxYb0GAtbedF0FbEHeJWcMfal77L9dCvLf6/flKHeTmc3pE
0lrhr3yhz1/+vEid75A6tlB2d1bBYi4lJFTGbVVMkGz4604VSey8yYneq6T3VRaO
GWHpVhxFcX0xARM3XTR5CMuzjd8xuBLgxxra59aw1CtTE173dX9ckU6gKywbIoAc
Wvbs7uBqt2MK57JxUiqHQMZ5ieY+jXyd2ELgTvGhgQQtjWoMxz6DNImhY6KaT+/O
zNDRZqTpHbuTkfeZbn2onB3Iucz2zwJiFH3wWMDHtwRQzD26xtIsUAz8KF4ItfCM
g5Lc9U5tRCNE8xx2MHTdeRQSp/20Me5FkI+29VcmLglMta4snTAHGqnh1Y/+7AW1
E7iES5CDr0I7D90pFUe9BWNcZ0qTydYQBAR+ChWLcyzaV1GAxIFxcZ9ZvSVXo+uC
M3UOTxrgEitRzeGMIprZKP1ZaqESTlcFTY3wlEdgjemzlY3bq8HI4+mZOL4rVh7w
CtqfgEIE4qqcXoPK7oI2Aaur6lKEgVIhJ9cNJveqkeZMq57mq0Q4UZcou+at4TAt
Dh6Vsua7Ofnq04qWxi/sI3TAHD39c4vgybpqgxTS/bP7rbUn7Eq4QGP39wjyXfbQ
iRSKmpiofcvQ6Vz+RIiYReXtosTr50YQctHsVE4sAZgecrD37Y3eJfH8FCiScBlo
+MbUQGv+X0axXbDfng3YuaQzWC+QT8pjVl0yqGeYjIBcEb3DCshyW2aNO5QhSMEs
D1jHi8DLE3HkPY5NqmglEiSxK75NKQ9IuA5Lho3ru775KMPohpz70lpPRC5707LK
5lL5bvOtwIqLUe5XoO/DHsL2wHomakYsfYk+XaEqkKg78/9cvpokEqaJuR6fI/eI
vUZxfZnlUEqT14njm+Cbnu1UWVLyS1xSVRFOt+NcbQGROVJAnfv43W2y7FWMosh8
JMjywEgN2yQMtho1w1Crdpm5YOznN91WGGJjt0I75NBoZ/3D8+3s52/TYDRnqe+l
woLpdFXj3p9wlveGN6xsC9gE2vBinGhHhNNX2ZdUsyaRAmbU/wUF5Po3Pu0Ofwf0
RTzIoh2OxxhiOSXuPLYrszGuP9Pdk0MtvHplvt1EqQtbgdASwwV6ndGq9QBETa1i
cIvN6D1LFTnLxuaPYHbIMSa3E/datVNw7u0Vw8U70YIvogmQNnqveU0KGLKeqjoD
4XPZephnNY5L/prL/xBV4+y90SwuETMIeVDxCd7wtj88FQ6RO87NTxgmIbcBWwLq
Zx40Q5V74vwzEtTkuOHBAy68abrqc4xwehYOV6jzaNYZudvqs3Ss0NSt94IlKs/y
cmWpU7LK1P0546nSGhKvhhEgIxFmF7AiZl/WR69tiuoMKgkh61I5FuTy6jgiYq5y
eYKrhEWX8s50a5tWuNBiIl+6kdAL7AHjHLVkeulno325XZhc18KSF5tsNd8qYmC8
EM642/kq4nN1kkCEDT4sjBGBV+gp+qpNkho/DN76lWIWSSyv6MrEGS5g1Yj9YB/A
pOCstrCheVaCzak6xyJj+g/SNkMbLznIXqQyN1FhTrF58UeYOZ1YlOY7hlzR6Q0w
Ryvab8xgcek51nO/Enu6FgyPMq7HVYqUHRUrYmZqQ4lenn58yYvlQCkqRZaRftOK
tjX/o/s995rSLZhqHWgvxKjkpu4JQZYjgLbzAuw8xflVMeHQ4BCc841egTrEQdLa
iBX1Ez0xfO6vFmpmxu90fQwgOc5xJc5iLRkAv91Ac8p9FXN7hdAYUN/GZGq2y0gm
VsrWyJbaU0cSvzLgqxBu7jptAxWG3HnWHdyaN3meJD9W0Otv+uVA8haXdjggiKTB
ziClUQ4p1UQtKK0WL5POqHwgJOo1vrCYIP+fd+6GaCmqIES49cyhZkfDHLPofvo+
gl+Is5qMEZrM4WzbB/18g+9gbwFwSlBLMr9Jp2k4F7YhRJiHhDzFLj6G5d16MWo7
+on/p1c0tLQruyMYo+dh9ZrSsiJqWTtTybqfFTqmf8iINbk5YWBwSWcbcV6+y90e
5jqiIzwZPTzQO/eQS7OC+bqwHutaaLw3s93S9C5eJ/ggF+kQpaaTXDdjbmn4BBYe
h/bnZd72+ShvX2AJSUwQFaswHjRT+d45vQnJ9TSi284EysWlqmycv6Nr0x6iw6Gi
6uRxAaylvjvunTDW6Lr+afxeVqCjHx0RPjWt4I8DgnffZVJzXMXnT0iyZDii4rjn
jutbYbkyMrakWu2nEm/a+TBl0tTb6wZqBBnJwCMvUmnx/+TKPWHx4mTbEWXfqaV8
DksFd/00DBFKOFjgi7h2JlyRZ2L6NQbTx69dOBGuJ4y2nrV5I3OQjCeMEJwOrBbi
Bj4YpiDi+GD6klrWg5gN8j/PMHI6TUz4muF3+rT2om3HQeMRiTtmpyCvA1jLfC7I
f1+xNUNic6zTbhdwhyeHKysH5QXiAxzQKAPtYYxMg0F59DDOAS3TbgpjUAuFY71R
ZAJPLcfGAnibEuY4u6VQBWKRomgST86Lhd2Suo1hUWcH9NTYKeZOk96Qnl+Bkh4Y
kpKimEs+uG3sfpLAaXLePJPPLva3BZhD8xgwM9q9pRy7J07pL8s11HqJIfmjCanZ
NGsf3UAehFvhc23wP5haVmO5W11n2J4vex8B9lnGjV6I0Kh5LxURaWRFbHXnuuCV
mwjgHV3Ay5mc8Ft3qRmrjvoFzob8cfzX6YGBAKJD3AdVKlPb31kjJJJflWImYP/f
L4D5FiXEnYfjkG39cIVZQ3MEN8pDvCxZJnEYetupZWUxJ4SdW81cgNMkkynQPn9H
cZlRPa+qEH8fsaHhlT3H2YO8vb0+S5mxRi3YxmqBysDo1jf1MSZD9BkQQHmNaHHm
4DQ/EtxnUoHosJMB6qZ+kJdD0n5mGI+ht49xac2f5zbR8YwLuNR3wNMN/3fRWwDM
ZAI4gly1KWvX6iD3+6EeOb/5iVzOGMB7qIq2k/5W1e84BLvhonRWfXGh3PK6kUO0
tvsGCQmLFVowWruhV8HA+W/oA3dHBjRr8/W7so7VMb+N8n/IH71vYGq7JSOoAFdZ
CuXWE16rBm9McrspHEE6CIxZWkqxofUmUVk01q/acauJ6ixk1TJVHUdgBOUFQ5R0
+xCwl6N91CW1Z9nmvlD5FqsE9tB1mJs2o7qvorshiMrAFpSeg2CRuT1tjXuLFsU5
PjUlU7gA5SJFdjFLxjfpgVAgOnvkMiRJeutspqkwuc12iJYH2LZNv8npt02cLAQc
RSxIeOYG5qVPH4mQJSjMDtuyNiJYjuuMWNhyS2dwswoBTjMBjZ2tUVsYV10Xvkio
9RwycwFbSSf9eWGmtIn+kWDBWdg79nJ2kSUSwHj3vwLsFEYBQ8xjSw4qwpu6LG2I
hkVc9igAE9T7kK2oeZPWOuNP6FTHo0aNledHmSAEHhDRdUWZfUhKBKo9F/3FKHVZ
yuPfX2LIhlOSi87ZjKx1L6KYS7WtixNdL7tT/POZaE/M0omOMArj8BB3b1S2yoYn
KGaPzHWHgeRpHCbPk1Vb9z29FJ6ALZFWZ6ULoI/qiKylCSXzWi9jqUBPezh45zlg
LV5hOzCbRemd3buJguImFvnImI43ywRMdg07hSntFPqoKa8oxGhjhR2ruksPulGY
GCwFAATvZwttvA11cCx7F2nAoCy/L5RfKyM8rESjF8xhYE84+y16RkHaSn5p89lz
0U8UA0jT6riVUn0F6p+AgW9sNraGNipCC8aZU5ANgrKUdpvsj42YIGvHyu+rMJYk
85W4ylaeg1GOPwefwryqM4ri8r3ApF39uAZOhOM5Gm1jpt6+ys9BAYvaFegpzKt0
sUwxH68kDmbiz8lvIVj/rGqeorudhs0oSJLabFm3jhC9wsnFCLQqFU/FH/4qxPfy
uUXV6Ri3tsk6XFm+Ew7xkT5AZUCsSfm6D/aVOU4fhqMwEF4mAA+xPwxHyAiz+AK2
7RxMf0WhGsM3hFWzCv04Xq2UUIbkLxREGWfXswEtB/RR4DtEl1jqckla91cBObDM
nb+tGF/Up7dnCP92ExBz1jpylFFC79qhSzpkC0J1loOwqaOu+GRAkadHx5e8fvN+
n9rKg2b0fnoX82nigEz+ZW1i6JQDrK5LOZ4hAPBFXMJzZyz6Aml+GwJL8d+6eQrz
O0vG7qDUpq6h7m3xAZRuwiw2QkINu2Sf0ksFDGg2gxOukwvS+oZeRiscvcTzpPHC
p32FS1Cj/iyYcp+kPepqy+wB0fBcXNt1l4+w7ZEo/FQlnh0Jlr7Dxv9Ek9uJYjPH
Eiitalf2bFrjvtXvJCveNGBU52pE5gmxqPrPTXvlyiN2BCjWIxwsCLL3pxjzzKQ0
yKZOYbnASyki82zs1R5aSMv36f6Q1NTWrGxRMZfhtGXdTXBIsHFAiXRMPGDpI9R9
dte37aSDpLpC8v5e6t0nXoo+i+qsdQPO5Sb0MKWPb2ndnkOyYETxlDce3ywiviuK
KzLjFS3bbgc6EIjcg/v4d42AWlQ5UV58E//PPmgxs0YdGbR5vMPbtJRazOwK05Kl
+jzIOjyJS2+v5Fls+AcVp+Ul4p7WJn72HqTGRttmdeMeHuTwidFONh8rtekh1Oua
ijOhtbC36NGE4KUrp4hMiD3pS4LMxDvxG3yI6eChO1nQdikYKwFTGMDgV+1V4HUd
TT9P3nGWO48t01So1DhNSP8lTrkF+mhjB0+09Kv348TpyF38kHz72u7ZMfPV3jYI
wXD+gBmTH+VcCgeoKtX6J2jcHIo8scROVNnjUGJdB4GApvOrtwjq4Q7Pyo4MYgp9
+P8+JtWhoEAoK/cuP6TU+XqzldNgpaF8N3V1Afingw4QcoKqjl34AlRcKqAzcLbl
MCJ0/4OO0FStOMVheM0g21jaMYCN6poQVsnNBMdigiGt+v7l2QojqXEYsc7O7KVr
hNaML+jtKsCS6v2pW0RpV6yM2ievx1Hr3xKM/oQrbtGXQ2TC7R9sRavL334zhYyV
n7kwvuzpL1otGpaoNI+zhfca3x8u3xYRqXwKgYIqy7Ud3vNLp/xHR7EZKbsGKZpK
o9uOOxElYplnAyBPILsyAqeiJGdo17mzR3xWh1Beoc1D2u/OInuOrkovYVyEZodb
pYEoc+Su2rXTF+ynXIFeJT5v7GlC6p2atllfUn8ZKCUbrF6oMZYvxLRGmJZfKejA
KavPw29JwUHhEITbi0B5Tmra03y1VI/vOgn8UsM0W72iAOO8XP7z/YWiKaAu1L9k
6B2E7QaoFYoK1yy+v0qHAi4X8cCQYxktp+Egd3Bc02FJ1sz4A99EQQ69jTwNGzCq
6RUEfD05yaP3KelY6E8hSTOfb1/kSMja4mfpPhwi5M+SSOEeWK95ltCO/Z1yui4h
4vRXCvRhkKR5+MWMs7qbBvTbwsheUHfjRuErmBSCY3W+aL9N0dtf63XR9qk+hn40
iVI82faH2Y8etjAf0OEkHf929WDWZMaGEUDuMPX5AqvlpBgehOPZk1KwE0KhXbMM
P6KBBZjqyRspjK9vIe9QU6MMJxyO1WUn4Eaijwocx7+a0wIrKnHf0ZZNbM+KB/yr
8R7gAc1epkrno01y2WLjZwcDHDMTOY0XusXE0whwJ30ODmVuhz4kYAVUEmH9zSWh
Fof/x0SFpiYVVCVUkJVn7qK7l7wt9o96sRnu4VTPNGvKtKJ8TRz+Opn58qqDXXjY
onlz/h97jzTHoKIdqyNM7IltsCAoOcOvdsmJRy68ww24PKluJRXo43PAZ/d5lppZ
B5q6ygH3zvLFXU2AGm3qFeJ2AyuR8TuGdMN23zcRBZQABJ+waXRtl/W3NcDdB2wX
vWFkwC/kz2VkgANVnoHah5++3cIsew+FVnyjeazfJKhXzFOrqeL1mwn1gHtl0pZx
Qff2ee5U5BDebtgRNhTm15O7ylPFIBJzlISYY9HcscS875Yo5GehShl5vv0ZzFUB
AadB8cFLRG4PweWan0D+I8bhNXSUUyptHGaFHb3tWgaHdqOoYdG0vJAe+JVTQSF2
7owwokJUIbOzNNaa/ceApqCLD6i+Px230yde+zsR2OX+9Lky+C2SdtEXwWeZOn8l
q1Jja0IdLae58FPuxgyzubR12o+QvRVmSczj37h1HZnZPVUkkM7w2GbIHyefXVQn
azWzRpm6qvOcxAeCeNFfwDSMS6dvQkMsNlAbqU0FW8O441F3vpCtyR8sIzZwr7go
iidY70g3I17ZD01jTEGNqrTjxMkacRmq3Nun6ATyFDrczg6/lsDYdYrC7VsG0Ue4
IYpyAAzE4ff+cynuxYSDT4E/G7nC99PKlUb5em2fJ58qNuHI8hQVYFquo03zOqp/
NK5Ow6aktDHob7rWZi0O1C02BEzGxWHo6dpZzqqcrdYT9DLYNeQMPJvA9sHYykmv
ks+gloLdTindMfCjwPIdU5xnvqfTTs3fI3vhpk742btj2A5Ntk0qPE7O56PabFQ/
J/SZ4u5rydlE5YUwz7ClZQRy14H0rdmMcBJU4u2QDtmCDrWp0ZofOWgfEW+NpvVU
zJ6Zq1+JOmAtbrt3esouxgt3ezhNJHaC5bPCbDTeqc+S7YLGTE4mXceRjxsYsTj/
cLbjQtdWD+xlZb4CqKvUP0lcsJOIN2DM1UrdFhwm5QKOzGANQ/1/jkQwE7KF89sy
3cfDgqg8XTyPVtP0SrrB/dL76vp4k2M0oAQO7tZt9aMA5e9vQsjVmPvYtnNoAWGh
6s9lS0ZZsjymkfAXgK/0f/I+m4srOG3DGdBNBox3cxg7EBJSagZyLLEJt986X2je
oOg0sqBGoFkO2xN1kFzveB4A/nD5lrnHm9dGRo9Rx3RaZI2XihyLSPibEi0OBgEX
lb0feoIYuwJYMYMM2sgLH35nLyj6wsEEt7dGS6PecShwnndwxXfjVBSBvhe3qHm/
IpB+IKyjaCYsBp2qotJCNSh5XY4hisNRhZZohG/MEbjKl+tA4shvdTRBu6TitqLr
kIR4qylcOhA3c4WqyyVautIPwrhIN2/5b+hNsCSgQkBGlmMysglq687M9733pRSh
e6Jd2qMACQIgqYz5hiCCq1iZSgFrt0IGaD/GO78nG8dWvGgieXq5sRufRrtLmHlk
rmPZ/EmkhKcUqTO2ERXzEq9Gw27cpcBbZDSo16YWjmZTGpudA1G58QGhhL/Xke8P
aRg22x2iuRkW9XCWDEwVMJ8DD4RL3VhSO2CPZLsb6QjVTl/g1713+y+/ov3Moms+
k+Z//s9BJVDlNxlB90C5UYH/r8/F/4zH7dpiL4LWDHb4fbxJExi5NVcP6ke496+k
s6zTDsfgNr4BKMi8jqJpWkh8vNVY6wN1B0aGsVr64htnG3v8pLM94vPheusqQP3s
5zMvCAO1ohou0q1MsQP9DJjLosThCwCTpAFP0QfUfA8tncz5+6QZJljEjjC8HCJD
i3zYBY87LYKRkhIfBZVXHVIAiUDBLzf0E9FRSpLXGs8PTU1VCerhIpvg7p2n2fAI
tMtSPkAwQYLNKdL79+Jm4ldT1kqcgp6g5IVDXaRk3GG7A14OqOGoYidbG6sXLkJQ
1DFy/K6WZsh3mmYEYeOuVfRdGMQfYnbLgeH/uZh+k7+mqLgpXnhI/Cu679+T43+1
2F8dZGl+YnTrONAZpU6+EH6DdXHZbJepHf1tb2JBzeSSA4lyd8mcmD0Ri7pBva9S
vXLtQhh2ogsLuJV6LPYQm0sVKa6denbL8B/fHJpPeMkX7CJrNj+Y60ymRQlh80uF
ql3EM9otAO8mzER1g5zX+K3IeMzrGvfqh29+7wCM/HQyKBmS3oUHWIYrYS05zeOR
R6c7QcqdyT6joYBrAq+ygubkXJCriHs++ijTUc07SMOirbC3SnSzS14gRgykvbbS
QJJcjv0EkG9KacwXne+SfZif/RRsMr2UrMocIpNajKFYjhtmP8hdw569z+Xx+eE4
mjg9I5dfRxWmX5RusVLQJr5apSFVhbQU7J6HK+TpgmVzFQ6IXsaJ2LWcnzh1llFx
nk7vQ6FMw9ToBrEQHjNFNrdbb0QLoYHcH0Vq6Ig9jIGGDTfn824hASwctcryT84H
oJfxJqCm72A3MMhpZvihpeo6YDb7M9fFr0mg8vjA/ycqGEwLOiSRQOtSwQ8wN7aL
S886sUfkCCaExM5OZFjh0zMlrld8Q5rnQroA9VYEpK5XDAf3riuYCATpwY24zCZF
XrXK4lSwCcuRDEfNcktrS+I2Yy5pnjg+L7uQ3/S416OIfeO9OpkXuOji7EgRTuUs
djHktatJmvEI5zoldQdAtxRat4FH/T2Gl0Me0aGNnYVUcabkxneKkeFH4uH4ZAYf
KEPqLwA4sEx6v9ub0GRpYP3CNjw4dTfw0YWTdy/fB6OS+8UtLh2XKrzwgdy6gGg3
UZCIszSQKhhoL63R+heWXktpqCzY6i4HS8bsHJePM3FZEe7uFudncbJwbi13coB9
bwOh5v/ICr7TGSLu1PsIWbZP2GHJloraNjxbFAdA7vcpl1lV0lPW3JAxxXqwEhBF
NdAVBnbZjABKV5Hmm8CbspruzrXVkcpwKlp5taskxcgpeVyKkailrLVZmt9e2gDF
Yq9UprQvf4L0mzSRtJcG25M4zCq5NmXlpbiLHd/j/S0QoFNenz5abI5icAYoXBMj
V91UwHpSU0V24W1rhxA5G1xpuKUSn1F5e6LWvl91Eq20Nl6ug8qSUSq8Hfd0+hc0
FiXf5pSsZungZN4QPd/MwDlR1kWRtFLAHrkziaz78iC8jqwLqtHXYc4zpApR5GyO
dhbbYgJeCWDc4fsD4PdVFh0EErwSq9WDb1PFAykiFSU4lBVO4afua6isVj9e08Wy
1+3NdwQbXZmoQjcVPGiDi4xlf2u3QMG5TXAWkcqlVwXQ0LDssdIX3x+F2IQXSR5r
Kw6bAKVaWTHcXMi2ZSzkOueixRf8Nr0E4wqYajTK43xjTc+2pxZlsIC83+F7VPLi
jq6DCol/9ZqkjcHN1gR6QWbzq9AcThbTZSHk3TyLitRhlvS8zRDgT02nki4k16lo
cqeFzrTVg3U4dEQjw/fb2G2CCO5fHZ0057ASUU2/Sa9vNk2mgpw2XXdI3QmpP8oM
uK0Rr1L4BD8QbcfDtIaLgZP1Y9tzwIEYCMRlsLvhKQ04+yksJ9tVBBMn+RpBh6KP
OgFZrfPkdfkAR49sThtCKEi/XfSafQ8enqa0pTfUxwMa/IMDNvk/i17kOKsGLh+G
ViO7nd6dTC+5480MYLHXVZguLrDQOlrTHeN7VJ8JHef9nuDl+3T9HHlRDeYls33s
CS/CWu4iokr0k/uN3mkAVpSIWL3eNOxLR9h/GynbQz5dHv5irJdhtNEqT40E7vRb
6dgPJkSJ7bWeFv28SO7KL/YHh0xWYVqrkIJPW5ihPUo8DWCmKGdoNAbtf54lTIjZ
c1MLyREbwfeuby+f0tiztgovRFIoJA6eGsb3sFKe95D9t50+fVrUxPnY8kWlUeCe
6mmoNKs4Y8OQrnZnR9q+99Y2S5ifRel/WK1P0aAXgf+rUq/vf6Vs72EynOlq3QOP
5XPVDD8DKueSu9U+jZFnn5DPj9mM9h5+NIVOzGW7I3vUp00g7WS4+4MrDb7RgRev
/BEj++SBwExN/ydl4NLe2DmBowWIET/qm2AwOwg5Gb0hG3epumZMW95arbnryIq1
0kMHqKLPQF/Jto/wQD113wxDLaYjXKlfWTXABCHZug7jXb24Ssn+mZVm8r/7tW2O
BAAYtJcUnfS4NvU2l9mnbsNqROiVB811GzZSTV7Q6Gqm1L5v/VX4uvIU36HGkRga
9AwXylIXqG2AdtQKUs5qjfAHUWs4UprXt1eUithflvAm3HPZR8j0GpLQFKKbXOmY
83JpvH79T/bY6U2siEbeqq/VqnIATE/ShNn/WAYMAZwdNjFa8Ai5Hz8Efp+8hf5/
xWYv3VajG8NGeqGUvcZ0mBCImCTIQzBQhMEKMV7nfF0EnJXqcyBLpOrrKl1X+4Od
2Zkf4qZOttX/ztdp2PxHOHRH+zNKx4Ie5BUbvq0+2Mq8mncYxEO5VD18d4Gpdlcd
tVTDtG5TeyDBrbsP1bW6VT4fkQEoEiTtuMQUfXc+9p0GIBfN0G8kdyU68AjmhGUB
THsmqPPAmqtL3aOPkHyu6yekMiLQ9inSaHKhiV2ilLii5+pOaiLHyLPjoSSDQNDw
SxHXjdVoi1IiF1ZeHUHaWooURitEWa89XUwwATJDlWtwqQNUGjgaeWedG4O0+Yh2
vn/gwXsgfi69xLUbkpWeiilMXt27v3TtrVq66J81pvySMLTOS5JualhwPxJmUKtR
Kl20/CmVTeQOwIN9WrzSASoO7h77vwnblg4iQMz2f2mWio5Xr0Hr/XjaM3NUQ74w
WfZfNkuUUe/KkBxK+Z+PB2Pay8GmUWuWY8HI2/kh39MgPXyVwe4eAbExoDu6Q4OV
V8gpXaOOiBBnoaiVaivJukOsd9jEHs3/rG4zq7WBVI5jKnMfVecTJG+uv9vKd1A9
lJ8+FR1w6ouVoVzmz08KtNYuwmNEefo7Gt3cSJ5002z4bdA5YNw95q+qZ0zfp5PC
7cqk44o3KUIAGCEy6SMPvngl/3wU3+UaLK47N0BZ2Pdf0RMiG5gDUb9j9npNKU6D
LudVHttVyJDcMs5b3gF+5MIzrWW/tSHYV19WItqiF0dF5yjSqx87LwV5JPs5QHeb
s9eVJbo6zwJZ/JyS0MhHItMca4lbgDh4jjWqvvvrH+ERbj9HhdMWeBzEnZI6K9Ss
9bcP0vuyep971PgpXUzLbmyNx+yYiTEHcrOWFWzvsbh11Wc8bz/MaMyHd/tMaw9p
CkYAcYpCsMC87wDm5au/CPZ4ouDPG6UeWhXSJrjEABdMBokiMveNMrUBiwfuID03
OHjc8QADM2HziSspKKzEwSOLhPcijjSsZuYTlWSgOEjsf8vh1qx73WIVnIQ22aae
MFDKs4wo7OAgqkMUimJfe375w67kkQzoGHdgcKdek/B2NiQDZETA/tyLdli50Ekb
acUfOcAJ6+jr1Cmvq20H4aHQ84iR7HkPnOw7QfDrJOyd21AvFl/DEGwUrDuOUkeU
fxw5taH1n6c0wEquuz0NmLM3nVfBRDeNHDf8FGYfabuFkouo3vlDBVsViujryHlv
FHPiFMg8fYpBAUDpkOpamZh2wzNI5C2621WABTrXkjs1w9w2kKGAiEjHg4SVC6n6
ITFZS+qJSM8qozWG+KzVzdmpmW0Xn6CQN8fsJWUptuHcLSZh1EDa8hO9VpkCP3wp
3Qp2Ie9ZFDLwxVmPntuEoBQe8Dov8Fd8TxBy5y2EZCW+I3Ya3bszkfCjUPXeIGZr
dzKNC19GBzE/MC7Uu/7lgYGcN4Bzoj8TpJ32ZD7C5O8GiHv+ZjRKeBSoU7W9bLdP
E1jb8W34LmMGbeSKAhgn2Mu5DZPGnYETrQr4zp2z6pbgBTgXN+i4MW8tAnQPcI6m
zIwAX72UwttMOFHSOrfpUZtnZ2AK2Wrr+swq7pKXSN00P4pwyBgutv/heal5zct7
b07/5jt1fbxTwFHY1yzYaBcWdESplntUW6/8qYMzNS1NCZ5GatccTaP3QgpoK/np
MFnSVs1xha4dFOXzHdbvIR1tuG+pFIYOAHDmxkVSxM4OepK9QeWxI0TjiO7UbaJP
2UxHNa2eBiqfwKufTZBrmaVxNY6QXm2FMN5Zy0CGelcr7lNg8g1099LItq90J8S7
0TeXpQ3AM0GZkqqKEvWldhu8TY7I4Dj9zCj20PFQXs8uQNBy6dS1IWoaTiVdk+zL
1sRFQuRyCFRS5UY7cXf/dvEbjRJ5A8wU3pl5f0e/TjmLHpq7jMmjvp7INgGupwZf
TgvOsMDaXatmQen02BFIT0eDZ5682mFg6jC8+tN2Z2En1CCSB/gAmpFWtQqHka4h
rAsZE3wv/mkhtOuPIpi4ira48kB0gClBlMS1uY54/7D//xwebL7eXFsppVJk7DIz
iM52pdFp5pUnioa3NbU0guBMdDYOICWxZaQJbPI4OToXLdSRDm2TyHTPo/w3g7Ki
jcXB0PY7jRFJiLV6lWBUsSJab6RFsgVgdxcK6d92STETSaRenjFqbobFzKFukAI3
VV7ZPOzjG9802sGIdfpESChEpmF7svjr+8H9xxI74Sh+dUoU6HBKemVdL+mb3ps6
4BhQB3AQPF2DtwEtkAkHZSjG7pwUWRSTJSXUnw0I+PF5bvu/XUQvjY7u7QhrrsOn
SHf3W+3uUnNlejV3jHxlgXxU9fpkULVKhDzvr7t1yDIKo5fUFK0RM6lY+IgkxkOq
bdv5g3RdvuravsW1HxyAuvtE0GFySc1L4KgYoaeJiPeVPUM7cASzT2He39Jx/OZk
tzFon4MLQFujtMXeUwwWzIWM1Xacof+P8n0Y3IJLz3Kxhm+994WvtJiYOKBy1+Op
qZJFkaUjfaVN9WzaeAZPGgYX6kgsjFrGrwZdfy9LbkuDTjrlzK7svTjCAfzuDoqk
WsGTI51Znt7I1FCkNaYf/N2IDqTtokx1ePd4URYYAfY7oRl58Ii3lNFoqRw2sWLA
OQhIm3ifyIt/wGn0NjZJsnb9YvZh292BM7NdzFz0izp5Le3s8Fp4WevGwlr7O5Kt
ZABcwaGnhkDyInbXJp0QjKq51oEKHVm+DkPOjTJ4A7JrUF9r6j/+n8XVqvaTogj6
NEPVwnHdDfKtGQpwlxkgH+prYsLdf58Kq+q7CKf09a5ep8Jd84/Y3NsgExMDykBU
k/G6HBjyRThayrMhi6t6HqztN1MmaHuwqT/3jaAGYWOBcvgOLakzYcuJ5DaxDPnu
IqFxV9aObjsBAvmOM5diTp8LdtR5jKUtiFz0C8IOrw3D7+kh/ZNH7OT47PqX+WQV
iliyRbGtvkQpJlAlYWFqGOT2cYgM94b6wTVOqSaxpKSrnnT8VfacnMuFesvgB5KS
9AiTCPe3/P8XNvMArEH0nT0RD/NcLLiGRjpLdasRbldzhNliCO034YtsbldZC/Un
T4OYxAF4GPR59knVcvfhOTxKbKdx4G6caHjcGSxrrz+x+8mGmGrVOgt8epOgDBGM
igN6Z4LKUxNJdaO7zfhy1+d6/PFieuNhfzNcfF9I15811rk9m51j/LCvN9hWKlwU
0SNzPDDuGkW7Cl0mw5nief7+BEvRFNUFOwHbbmI/fjmnnAMnsWwq4PCEeq1xvjXq
7g2+x+dT2BGraI1ENtK1My1QcOksPpn77AVpHmWMbccn41Fly7nX4EYo2zYgNmBj
JyDssKeNcOqX3CDFBPbNpIXkFCC5Pakpi6dTX5gfmCChFEWffZUHz6NvthStwuKv
MiHW13EWrRo3vk0rSOeA8WZ60O6EBrRngf9CC80AuEydkXrlWSCIpOlXs9eQ238q
AYZPbU+xt6FN9KM0VoAg6MOQtzcc/Iy3UtC1XaMMVecEXAfh+TUtJHDav/UMmumz
cO2I2QAyYlCLASWxdyXwe7iHFF+FsfEN/T1STFKhZVKHSmfhc7V6Vqh+Qket13Hg
i+qHdrcy2PPMtgc5dXdNjxX1VvVQwHdvV1PNVmyS/Fro9gU5WWJhVCgIdwgBEACK
AQEJV2AnBvs2+tZtShA3xsfkEGg0mDIKKmOXugz1Dv3yof/7LV/yI63h3rfDZgKL
AE4+FweElM9V0HIna9hlryrzREhSiOK0cD+caL10U/TKfD08RP2rBhnlExOumb6e
5zKSRe6MeZrN68sLAkpzpbOC6Byf5ua6EQUPA40pIyI7U/AyMXNw8hx7lOxzSytX
GRM94eVd4ii+iqN3oOwatyPXWLwrzgN65/5kYmpTjd2c/pHy1/pG8UsMrndHBg0W
pBH/fGlj1F2YM4M2iIsyRUmi7vNkUD26jks86BdH30EoiQR8y0jS8NEX6nGA4S7P
Uw6qHfpZPPyGXJv/gWajIk4aoRHwDtrgFq2c6b4I3awJOYuXd3t3Lf9e+fT/AfAY
m6sKWRCfk5SQpVHDUHDcLwwovrfCQHEmshoDmnBu9pOljnVHmi7WIH5mkvdXhvjq
MQlMy5Cv5Ccbz/DtXQSwV480cSu13hWRByD3oGZQArRfCVkdopgz3iBzOj1MYqU7
Xa5jyN+gHQURJ2nYNdjBi9dFeXtWvpuffN3zYTGuZcrGhHDJ01Y7tEK2qYLmf3eO
ebplYCOk4FSITp3INyishNLRNzxR18eSnFEgu4YIaoxA3yI5zrpYvzapOCM+x+3C
AK6AYz7zpN9nrznMVuYMuaSlpQZ4cMfUyibmK3xG2JpvuFUVsXICKX+7ixpNzqAs
Z8+96hQyZaMV6CsyWX+gkBfRr3Lm9/z/ChT6Oa8GnL+ebOXBX4uYfk8Tqnch18By
uDJRgb3ZDGiBhRblx0cHVSqi5fNtZ2g1oNvczqo3mlHzxUb+ZDd/OpHZFlHSd1GZ
nb5CW5HTj9CgA//QT4yqJzw7ebMFjz6LllPaIN/n6f2OvT79aoUFrqcKz28X9yj3
EJHtNQ5OiGvZjI77ON4a55K2goqxBS/IxlsCSuQIvo/ymjnoAt6aETMrbHLapqjX
aOlifUE0qZzehzc8aEtgviQXR6sBZ0r+lINkekowN+JJe8VyxFUDul5vszxvZ44k
JwZh+7vaQKOHqBQWEXPQ+CVtIaKwY0WhZbBMShfXCzIwDKsLG4H1SABeorCBqVcK
BG4Oqc3z8pryFrjmA9WYg+OdU0NhRDHuIADsTH4CuYD2zz/YitKfH5gt02nrVHBb
hUVvlaOaVGcT4oSVnydAGU4w9BAZvYCNa4EU4VXwZsc/pa0yhO7tFZRoESPx9W3w
Jyw7AWeJ0GBVr8Vd+mpcBCkczKTQNhk4zkbuMZEsSxhHXwrQbhWPBpjx1rt1zg4B
PBhyxnNY8QG8lbVkTW8IpTwbHSVfaKoQtmt+jwRJLanrMIOEqMCAzjAoPV2axU4o
qYwMFwlHZUV7B5Y18CpaxuimjUHyfIhzk9vLbEnXVAenmByoLSfuWV2ILhnMlTn/
KhfMDz8i9E1UN4WoOHHdhQNaYVWfzvCXRuAGgL1r+uGY7HA9Hlf5QM+XGFZEaTVs
+DN5AqOmln3RWHU6nyv6xMg92UKOkZ+ohqvXIq2/0kMuJCkOIICdFen9hZUF18ZP
nB58dpf8jforuLed7vA2rjKKWem0enyKhgk2edsuVSMUu6LDof85L0rLVR+srBuD
KeyZsCgnV6ls6m3mBzfjN2j2RLrPWehjWOW63wsdHeyASEylJlOmf9rTRWwMMNWb
iMUKf4SNIxdlkl/OEvLchUCZBVVhDF7regAV8kYWQCuBt3llwtBmUZ1X7n4owgvI
xA84Y2fQTTgv3cLhresvO4sv6blN39xgxX2rSe/4lRvowz73QsWNMYcN18O4ai1X
wg0WnxxM2L6Lk9p+KhQOHeATnbwk7AY3/ozu6pKngU8stGR7UMNpWBC8iDqjSd9z
BqWcjdpmjgc4xc61hwAankC3IUg1eSOik5UDNRdewJ6HcI1VI4yLZU15Mkk5f789
xosugPAOWeBy8B0k4yMLcIYoTQI0YZEFvC/8uTo2r7ZJWa5iQ/MIfaAgwJ/vRePQ
IR5NH6HDRsOUEt9QhnmgnI/j43GcqXohJh0EC5bfrEjJoZpk01SZVVfYV1Shjd9/
tKCAtBQnhst9bYVQsDvXQv9Gr0QMjCiXciUuMw8SbX3kTxv04oRqz5HTakpigJO7
4Ng5f6Zt1bi87OVGh73DqZTFBcwGiI4vrSAEgPJT0xxSwIncoERXJ3Y6XCJGt7Hn
7Kd4xIQLqemZ6AhIt15oNTPnO9QKWB1cTukbL18ccMCmTCF45Al41dottW4VLSUk
idYw35g0hpfXxAMVT3+pIyuWmOma6xnvpHriVgrKHxNTUsT2x6oVBGOrhvXNosYT
/I0gbX/xY8Jx89gAL0tslC6pEyHQZyJIipqcaHa/G73PeS3GfBpOTAxwuR5qpKCs
WuLX5bPtiYWn4e6ksCKeu4bN/2sNGPMPB5E6hxsxKhcnDVxEzhVKNwC/P0vBOcGc
zm4RBgARAB/erGCN4S+ODD593G91K9DuPR7prVnPV5q+KXuRgigkMzn74XEWzJkC
HT7d8jPfUKcP0k3neFunjhnpRZVyFGCBWUMqztIrh+aLNUMj6JQCdehU1n2RbyDI
M35CYG+agaIW07bURqOgHa/VXEcBOajf2HJd2X9u7X/AISJuj6g01N8eEydE5Q7q
IO0tkWx84lY1QZJZKhj/oo+m3TTJBC8ip2FWevyu7vNDYIY84cXMnV+o4KcXiymw
TY5OGXh3CfsgmyXymx/dlHhZM7x9hssV1yWVmE4PTH3EY0zfLcnsMcAFjGY9Lh4E
do1yKs3TfhK+7ZsJ1LEj/TCXC9nEk4WoqCpXvgWFIa5+yMGN/7WuBVhrVy69cL/X
QBAXosUGmA0bmCLi8BQs+nbRF7KBL7rufZW3nLsiPDRtutMG9TY6uvvhx3QHMb6j
AJK8e/IEOxumPPDraagezEtqfOu7Nhx19qA5az/EVzBSJMevevTqKMTPIo0Fl3yX
mHVUJh0ezesyR+LE1l+boCROYwAg77s0DsO2ME+tBuRM5s9H/up64ouOoCyKaGnH
CWR1sX2pXzEg4KA7i5N+ZPtjvO2ylP40M5ltlp4wqzfkJzogJupNQsC79ENYRIiW
pev+UJ7mVIUtUEgLBCMQp7kH8SdlTYEO5scI9973PCLEK2090CVO/9qZ+7fxqa+4
cm2KesVFQ8fJvL5Dl8txIJSQPJYl65l7ajUWhle6OqpP3UrR52YRv7xQLqFE51ge
prTSiaxpIGRUxM75zNLm1DWCEPGvlXIl6r24OQMLd3aPuPhjXPa9Mvyw28iIwZuQ
94zwzWl8jScZGJAdsjiE22kb6y5UA28eOT0H05Vx/DSFG4FRtEbPba+MMFB9I3XT
HNZu5h1SfDy3MucyB2PrE2LvwrGZTwShZIXwQ4bFVzswhg9WjuOuvWY5G8yxXYEy
aRmrE0pxwdpzMdVr+VTeVJo0xVVF+GQhqQRsQl4cGLxZNtB1hQoMI9kXEfNx5a8w
L8+hwRlBraVTjoDwyjRKFpl9CBWDKXyfQ3vX4UbgsGpMv/vUN6fsrezNJbhb1vWr
eeyz+3me4xPirpFQe8gG/5bZ60DtR5XhiQDEP+vHRrQVisKE93TtTKMfa4W6Fxpx
D3pYByI9jMHVoLLgs6zWM4t9zzDToI/GZrnRUPutKZ8RxTei858otTUzfqMVA9EA
m3yLP94dUgDxUvvvATUnY/v4TPU5ml/OCbpOqpgn2k0S0Zsv2OUBsEBrbg6viANS
8RM8uAhHP9nNze/ukqjjXh8lVqrKkG4Ab9Md8P2MTZBLw2t/yAGjaJpIcL3cqNgL
wTGv27Kr/G/8d0ZUvtVePasBg4Rb7WTNlmD2nxIps4p8f+8dPmVioxsKo6tyV0yM
JE8nULTmipRNvMQY6tHaua128fLNdadHfFDZJYlnbxRsX4dQefEYslJbs2tUPMtS
l7F+UszF+4cWHEmhQQ40X5pUKt2l/MEiGsMpeRiNUepHB/yQAzgfvKnOZf/tXjuf
29nM6KnH0bEJo7f+tyblYv/3O/5LH6BmILambzRjBMjc3U95xyVK2qH89zlxHVLc
KjArvngPTrrT7TV++/Bx2BURo+2VVXc2NPeoct0W8n/MnpQdlHY1mv/teHxUGXqY
1JQBGBLHqDc22/QRArtEc1upJYHVbWJx0zxmMz7B355TQAtxAVQ8LDX231cUr7uy
PR9rMI5+945bQYJesIEIlac3ryVpUYzgSDcb5sk4A4+No/PBMQP5dP0nSZe0eewp
Rfu1BWStBTmuTjVBjy3JMe0FArVmeC4nyU5mr6t6cZd+9uBGLkhgiS+xPuYhAVJg
mM0Z8qPZUJGZ0Kud+drdfB01YqFgWhbjQSsCE/7taAK3zX8Ixf/HFtfdDHVQgFHG
LwxzMAhZrkksBrFlXRV8E7JF5OTiJDEjp5V9uiF3XDbHT3O0v9KskpHG9LtiRbtY
fi70nIIfOHL/MtwfHCjNR9cZVN/JvO4c+VaQg/RiZM8lCrY7k8wWk/Aa8SIEZmVf
KaL1eC5E1pgbIO8/FT7oGpHgjqxcc5Ezwi9UOpvUVfKYbTnzOiafPK1uD7GTBaSl
RaHVjTk+ITea4DLV/594TP4Dugl3DAoIl3zR2jbdwUZKrstsfkVS2kMid6jWqx30
V37Chk0u9FdTlQUm05u9/SvafKWeDNn/b9C5X+cPNnpr3Vts5zLUL3vtRjpTD6wj
vicwxH9v8WjuhEjICO2ZEAyvLPFSi4pI4IgbmWWSVYj6xfcau+lL86w8IQYrLhi3
WFkRsdep4xwp3co+3jzmbbB3Opxda6QASdIuNqCjNwUDTBjL6HK2JhUZGzPeTbO4
A5A09ezjzkR0YVPLYoUMEXXhzBhNaivYyUkGsJDzrMn96vfxIj1rGRvp9cW8w/NA
nkAYhj0ehcW9WBfnvCOzNyxGwQteE+yqs5SMAUhsr0mTluJvKqEIDANYINmqrl+T
znjBRS+C14dhlffLCmr26kdk3l3nu84ehES+SzsamebVvtG/k1e/ClCwJ6qBG0Li
PbrqFDn0Xw002HvOh+9vIqswe4aft7LHywh+d7EN6MQkZgjiXVnJCHyZ/NI0ALDX
vs8C88sL4yYb+g/RaENwt75XRI6iLFCsfpxvts7mZjoIkOuOFlIds0l7pnKYAt6e
yl6Cqi/3eXXlC9eAMmaaYIL/CBk4kIGLggGd+iKpp7E0+WrB0RsyMpjqKmnXnl3W
sNeBBnVyne6itQGgZ/g+eSPJqn19eH4YHw3326JkCxOeKw+PVxJZBcoSlhudIqmE
+TVlEd5Vr1pUzOG1293wtr6/yM2khX/e3rvkXKAq1LMEudR6CliQpqkz6aIvSqFU
G475QgvN7JYihLzjOTGjCxofVKw4yM9Bw7vnwVmrYti6xEK436l8dX74yeUmH/y8
mxjYbUcjc3q7wf1kQwbE+yYmQTNZlP6ns97bM5cAGIfrOEMZuae3pkOtxUaGsD/q
sxHk4u/OggW08bOMBz1Ihx6cslDWMDYEpknmoUVqQjdqVV0FgnYKCj38QSyzjbaC
RcNS7jteNU8OkCRhyK6nM2KuAyTQAe1+S1jbk6sCMRvoSUOITdqCGwOXRDDzNaIK
d7hn4g0pAHIuqTsZjM/AnwjYAGXCYz4huAtMVLpAxX0DvsoUp2ghQGcXuk5h4VVd
UrAO9vHcct8Fl2UehivGrUr/RovCZU4ZQQbzD/2azrLiLlSE5rB1lHAqqEUQubKM
RyHmZfMxR7KxIzWamUXXvvNgBWxecFf9rt6LGoY1giD467pyM+IAyJUX6lhK5hbP
Z0BiPThfk4r+OTE+PLYqEthfHS7JJGfy29Koybj/hi5SYYwTQCMyqSkaaibMdlnL
frxzb2AOTr8Liz2KVYEPcFQxr9carE8ox1+oB2BJoCUulZxUc5yOjuHFGeDnkQ+n
F8AMsZCEj7J+eRrD4AslhJGgGSJBREo3yIWUdLybnNcmh7KVhtwDnSXiBealtx4E
Z5AIAmquyGZ0jOlu9tRsDthnN1mW9DfV0gX+TQB5ozbIseELx8APUvXazyBs49RZ
0gO6SflZyrJCNOiVUk5bTBhOCmQeY5DR9k9YnZKWmuDJST1cI0A0tz44x+vyCBuE
xFTzYFp3OLch4ZhdP0eoU5QJzkI/D6ayU1tkVfy/xDzxwVcoaPHi/YdEaAxq3ZQe
hQHFWrrriIJuDFzFPkDNGfLpgY1ZiACrQF/D9PBlxVCbv9xW14Yan9phuXf8EwpU
bkwxL2632PDbcgtg6Im8CuLBxB6mFBA85Eu30cS/Uc5vyMBe2dDxaAOFnUOANqft
Cm+0U/g6rklsQyCMet1k3cN0Cdf36Xji9MBKrv5eXsWGk0btHpVo0fzLyykwp6Ag
Vox5FfCr8boyWmp7msST+mBGVwGnQnQ5Mm1Uitc9oe1Y7eL3JxDk0ChlADHYIliU
QFsTivTDLDLZrbewIEPocN7zumu4Vnus6LNAr9mv4NK8bevyAB27bPGez2AND3ej
ooSetpRkuEp5TTdOkMM9Xy0Y3U8bgq13F2wjCq+hRfvDRIUpLwBZXP94ORWG8XTO
/KrLcs8Ht83/DzVqPXQPYrRteNJSGVrTW3sh6BVixGE74HsnWI05oeZRb7B1C1uD
74bTnZk4zA/WLbQG5mz8neY/C9vI8zrUHz98T9xzSnGuirxZ57iXKPsnRrEOAmi4
ZbhxwSxhZu252wLBeZUCnHJY6Cbow3EjVGXLmB/jbuavv/+j1Id0voi2HlSzBfJu
gPcv6FNgXALfqiKPU1GCWmu+LoM9GgC91zhttmN6O3imMYSt7aee1C00ybg4vZr/
1lBUjaarpnKdDXqn/n+sLnNxUqUHliqf/4nz34RMYWR9SBjcuzVPKPMj5qww7yLa
opc970awR3LEHWDSp3cpifP5ge9e6/7u8I6yqe7iDwWGlUUUwJW6diPbSEx4zkfD
fCo+c8OTMbBHXfYmJJpqtHfOiluHg6+2ThBgG38qrxsUk5cFpMNNSlkjKTY/zNil
nIYueqK7D2YjbxuJaDVPr2DCIkDmyTLLVq1ePHVCC8wFxJE4UJvZArePrNBKzXZ+
cwOZP3HyxO7IQIe39/3FuLJa2Ter8Kv30jWfOkQk/i1uWy+LyRHtLxTNENIQ8iCE
eU3iHd+qehm9H9C30uEkIzykkxGc9u+rXxjKfTzDbgRJbvrP48CbTsB6FNIIRc5Q
ILOWjrGRBHLzXpm9R+2xZtn+wsG8L5lVU0teU0NzZJWgbgxAMZfeJgf5LwJYUq/t
YjqTkrKiY8QF/rudyWSJLTB6hzgoSBsk1qvo1QCzpzHyzFumVwXxCp7x3zsa16DT
83pnEOghEo+UnhSq0povnkAmUJHS/eGTsveJ8Hm5350xNZKg36jVUpl/BMe3LaO+
gRFcCYK80yvcwx3+43GHAOFEQaUb7QUHtm0MJylHfO9MATJUXvicrcGgy1PgTyXC
l2EtuX0YBJStbjo+gm5KTnbxo9YQ2Q6YQYWXRTCbGlJnRLuQI4bE4MFEbkrh8+l4
1KHfQYl2DmIgYBmd5HxMfybeeWP+P/Ca6N740yK7YQb5PblZLGheFy4YD0Uqrqb0
Sv1l00aZI8cHVZLD2bI2jGLbDFmy4kQHBA30r5MndFjh+QwBJc0g3QdgDHuHy0Dt
wsXrtd3sF3BfEtG554tV2x2OirlcxFYyu1S4v9oMwvyQMpBD+2diYHnawjz2Do5G
KE7qaV0xE2UdQJhXiO8BFPpxxfbXjwah9XJBEA9ufy0y9wedxo5g9oRWCxVpgIWq
ICoWpVXpalYO8mHMtJ5ZRp90EtRBpPKWGBvibjPhEZlVP+bYI2pE39SxlImnTbjj
BV8oVx9AZyqxmS80H0D35K9sY6c+VYqfmzAJ/OCxl9DnsLEF3aarkM7DAO0OPr5/
VV8nl8RK9REPPyTwEX59YhEoOUutmFbNk6wnuzgLJCTQ2OVL5P3DQxTTBppwbgw8
c/LSlSe7k7cypbdIRLBORKGrEmi2TWP00NFYJHK16BYuQQTnHGE+bhd7nANgiBXf
f5EGGZZAN6w7j7n8WbYUqtUga94x2x69/bVxBuc7rGkb3TuGtNXlMaQJf+qsSrMo
IKRCYhbDghvZ5qm7qNrUyJ04Lpt8eVtM1v6RYSt3KlsUYuJ8E9IWoGRra+YUwexK
vFOHasfyxssCBSAVekEdlv/R9R8hJJ8MRDrkcF2Z4E/BJ7WNlVRQEidt9ubt2cXS
dnnPWXhXKsl4/iv20SHQAAwGjr4QM6VCB0T7yAXJojCQzpeR0WJkKh2xvaaMITtB
f+f1jQ6MacgYd7pjvEK362fPQ9wKovnnyStAlOqJRRu4uMCQ/xYFAbwWSiKP3LaC
JzF0ann1nuNqzt7jGPyGfReWSA5jqyG5ZB2Z1/wvWYQqUThSvfd6xHVerE1hjbny
KhLKj91s6AZojH9MAod7KsJnNUm/cF4DIJG5wkS6G9djHJRKZPqaLCh3AsCmm0xI
DT8S49iqV1qkunCFNKKDSq6igix0LObW2hp/YJqcvxzJvjJtrNSPMYydQPqiP6hf
0Eg5TpSC537F49PKsg9bVRe6BJ1IrCqt/6lZCKzfAvlNd7hgS9OmQsYcenKR+pHJ
9Nv6uREyNI6v9fbdLar8rVmLEQbZr9ftWq/gO5pCJMRfEFSWik/zPfrgAxfuT8Wx
kSaUFN3jMDuLyv086noPle9cJdHFE+nEI0yYmgBOkOEWZYpcqCLOyH+5C3VqKJ3D
6wMnt2RjeAlHsqvWTIcPeqZAQcznZc2I2Ftr1+kUUvHQtMiIAuDWARgLT6YNLBNl
ON/JzqGgYkAEFeo95w4OSjQmD9cbqF0hyIY+viZjoARFlUesV37hipLssno+Kqe4
hjei7uArBfhG7C27+whVNdkpuy7BzjuXyJeLsRff9iXKFp5Cnj4SIE1dCInTHkoJ
ZTdPZLdE0W4uibNP/qZZLoOkQXoDN8RjDbW+cujGs2qnmd8Hhr1+ifnEap8ITYJL
+8hs3OAL6GOGvfvVr4EBH/xRY0XnF5WN5KNOvz2CZKYjDGr9jmqG9De0a6QGH1rW
XBsusfqLhgx2qr8v+LQgVPFQEfAtELJC3HbJtO9+QN6ShDtHCrbCKHIh/PM0ox/f
SJ7Br7Lf+FvhGBptwehTIhak1WGCM5Ze1TnO3B2KbrTbVSGsk3jtN3xiaKiPKqOQ
VTV8jhlKZQhqo6NjYJpRzxMH7YflTqrANpwi1hkDTykrAzstkxvZc28ZinkR69/V
z0ZiNWFmirAvYuluxuYeO0PN3zmicFjKDCRsmJ/aHFgddrOsbZ/bdNpYZmNLBKGu
tm616QaJ8LtOhKcsUQTrbXlpmZsLIEZTvVi/VKh+gZu6SxbICSN9ZX22yzc+X195
Jbz0LBbQbXifL6geJ7IV7MOmNx9+yJQZaSczkrjj+vIQ40hRMOA9gDIDr5X0npiy
e/SrVFu5sHKeum3YtgVOyQTasLSoe25zrmEj8pYU6cTcieM7i3AzBZDe/pm4G+s4
1FbtTeo0xcabyPeGQfzp+I84cCxo9B9H5NRCGu+eltjSXrpQ9+BRDnl8OSMaGyIB
FiZOfIUbIpoemU/7jM6nhjUqgsQStheLJdp+ElMRvwtkNLq954KqtpSDatADqvM5
OiEo4WN3WRZ2r6FHNSH/QBb583ZD3HDJLTUf/zAuWKuSKMiA6RnOF7GxJLpiPy9p
TXGAGNDDkzJGnIuzh1rzeSBsDAc8a5f3h3X2kD+P/bbZt8hBLMm7bvtCGIwENuMs
PvuaRKLIFPRo15TmbU9dH55ttG8dHLRUxbOdBV+UyhsjwfHEJcXimo7bTwBG82SR
a8XEqngnWs3TEXXXWKaWnNkKBOMcqdZJpHluKgBIiBhMP6Mjugfi0BfZ8r6j4TdO
EmbNM9aMGQWsXH/gtAHLd1QPRv0LVP7jNapTa39VvsuwRrXUv/qLogAwAR9+VYAn
X/9FaCtcZr/n37hd8fFkB7vz5lZM9H2W2yUZoETLNHqvfDYuOc3YISzsnNpeERyo
9j1q2/Ugu7N6JiHqN+H7qcj+TmLk2l00sxA0LMzJR0G3Oaij9T03qEqci1gzJspZ
GLviwdJGW6Ncn1yj7hg9OEGwRx9/W+MQvDaYpUCfrzjOcQkAo25J4JIb2uNqEtdK
TVVfmaA03/tNCWrLSqGOjL2FuU4XolHJ3sObU3+Ud5dTO9e9+bDsKfNpPJUKmnrZ
kN9ONxxrZQsq4+9uQZ0cJWhJ2y9N079Oyhq50YRXBM6eLhPK8AOao+fACrSQ2GMY
VZTOnP/MlGorSMOFhfTAj1R9snWzEsBJA2qlVOf4wG3S0bnUZFDMwJgHUEKaPBMt
6m/bhfWBVbnXIpcHT/WVgrbPnOZYLSVPPRxT58lVRR7iuvWtNt8/3VmN7UUvF156
OoRS1sps7cpPLbeRjGoP9QCFPz5CYs0x6qOpPvgGw5iH6K7jZvv6gc5rIDyyKdVK
9MZRIvOK0jfw4R5OLJ1P5Grh60e2jGE8EABL2j/a7eeMm1d91lbAK5Ei5SfKdFD+
YiP8MsMDwBUmeJgvWTYzwFZULsJHso4NB5lR8F1GkJORBkatO52oEcy0k+aUHA4W
shoSm4q2+3z3fZyIXP5bo8a4YQluNHYH01JogBXLQr02ojg2B/5b/KjrW28/U+yR
pUHCFv3FXmxLBV3jQnELrd5DmyUriQZTfKdRDxRKSrjPBHxb44H+1HeyzL3T3pBx
pBXpjlz/FuvHQO7AQbgcG1Bz1T06S8sQC0SLXRmBGMhjAskjG3wDxoP7Ic7ZG06C
r+Hk6CKHKo/MFbmdFCNaA7Iod72MP5lQf9J9wnOWNtl1P5wiAdGBGwB823cUkZ90
Y89VbkwzJbuklPvTmxf1LLT9M2fopDGULxpZeqKd14IE64IpzSbGnv9jmk2csYIN
WGSW2OLRlIFoQcVZJPzb4dzXpq+SPz0L8j/qjuaBJpXLbPYmxD5Asx5QVcXlKzfi
jY9eWfmeifI7Q/V2T2k47lVCyM3g5DZxAjgX8uI4BW3yq+ZTGV3kj53QKKgvGGCJ
pNKE723HbaL+DTXm/C49VCIaoX4mg94SSBnl4oiijg1PfrLovlwAwPvf21H9G6+e
Ar9hPu/2ES8O1BxBri4GRCAYf0hW7xn97SmzDGMQIl1Z19rJF3UDFPQEqEko5YsF
Sy1B1Si1EQBM8KSk358w51ygcDB28/IsX/dPROdcKqjIe/ZVVEgF1YN1pj8FRQMA
it3iM+nlQFkezRIYn8nfhoMfnIFbGon5qtPfbH1+VmcNH+vqETL1IQeMUdc4jjKe
Ec/2gg/RAuMChCy6eKEjQsIZbpc3CDptxM86FAfXAT2GO3ZaG7iKoCIAIoyI7Ura
KDlZ33q2z2nNDsQX4VZ3PfUt/zvhwc4tlu77ZNr85xcficjXH01sQEwlVDFM1jG/
QLqD5QnSHwMoNfUKTqB6653KT+eLehhnrD3mW7I3CyZvkRQiXB3eFGTvOKfwd1jq
N10WpAsbM86DGU+jqJWRZZzNU2YXVOGkSMmXR8O9z3z8HBLmZDx0P3zEeaaNuOxB
IOiZBk73SmWW/5zSyvCN1DcpdjgMVYm1DmRUG1g9xl4VFvAYwBfbsuuUbGiGiE4t
XdpB2qyCpcecLkgFrtu6PIslfjn7stH9NjEgpke4uH42WHQF1XZCIWhcgp0vbmjD
l4t76Uf4jDPzoeamQzq4n1LW7jk6ud0RGVX4ZKc61iUb9kf+G+AOlFkwlOMmkxsX
d5T00j75kD515IETdOtjl5mBiJipjVFgudqBK+mFhvRFL1mFocOXNEnyGR/0rQEQ
09hyBEOp3IajaCRhTDU7TpX8dV6U7hFnZ/N8onmFiCeEooOzyvaRtnJp7Po6Lhh+
Fbc3OBB74p6aDaYV7smBPGVBQM8fY1/z6GcinJGsTume8E5H0s5jOro9hbFEWuBX
1tYjXkm9QM1W0ocIaWiObldJVRFTjS2ZLr0nRbU7vzlm/1Y4UiHLMxI71Z9gQ8nV
t8gm5nu27uMcrufdOh1qUr5Wg226glWH1S5n9wBaFBUWdFWwo6L/us4XgESnBPI8
Z20Eiq535vfpz/IVLnkrONv0REfABP40UURBGK2bMm+o9VQPR/l+HTAt9zkjO/Vd
oTDdTWMbm8QmTC/7WlXye/WGyJfrz4PBtjjO+4kcwZo+wfWMHP54dzk73g5jvLXJ
yx88iADLhZfvjuHK0R6PUkz5cCIDjfiJswc6hyOiU5PreGBm53A02jZyet/X8hzG
EuQEVXPMXjwE10LKdhmnoz+ufbml1tu5zB6537m0/bf8Qf/JXOkcFYvAQDwLiqgK
qjzBLvKPbkMbE7cmMR6fP1HOaknb6t6+DMZ6LjsXmAXOt1pAVZ47Mfx6j7HcgVK8
u38vQvXzwJmZerjR7GuZTxvyXliWHotzTolpLsuTpW+rbA1nH0iVjw8bnTzhztEv
7KG/Rh7Cr8gNY/51sxpdMINhJraLArqIni2JGXBd98IKIi2Z61dwQpmCqfe5kL4+
3h+tlAQCn/dLF9ubjckK9eXkmpyS07CqDR7tcn4br5+roBII2txPoQpF8ZGKAjNR
6W4RY9PtSQcoheJucRktRNOrl9ka7c8bvYTyUPbw1ZOOMWDSXa3viN+Xn1fRPFkP
cC31aM7ETtjzdonmhG9qvv5Ep3XvG/cpcARJ1Jlm0Ou2dwEcsE7SKMWkVKyP4/77
1jVtCHTNlKiO20L8vOtk7pAXJ522BhumiD7rnRvwscSjBnEZb9YQxtBBvetony5w
24dvGp8XleeOi5pDtlaRhj4ir4vN9vNum7t7VS4WYOUdbU36dBTC/B9hSVWtqvCF
/vK/SvO+uQb/Txsn9jqx9pJ2abpVUfMWcuyk+Shb3hvE9GYvAd8+A4i8am/M6OpE
FPknsliHi9fR/LGRCsa00uNApeId5IvrB5ty4VZDTKnb6pI2xPs0PPxo8AZRB5g2
PydcrG0NvQUJzdjc9iukgt/OqMjeoraFd+z+6O6h2/5R7K51lINBNy+m3H7ds0YG
HtXlas4vY5uxXMptcDaP+DhG0VN35y8pxIg0rewZTYjiS0h+fPllZYkXJAGF7AX8
MEMorIFn/b2WMQQNmP9SrJAO+uKJ7X75o1nLw6BkJnAmMltX4QzqIg7I27RgPsnZ
5qdu3h9eGEih7vZe7uq4w1698Ogct5uozs9vmkIwYjvhCUawMMtz6r13GM7kGpqb
8GIi4HFPTNB3ZbKcBvwyT/dOcYHsBtNK3DPbvpBfmVvVcEWLPew7VEe6zYlZxsbx
ogGAOrL7LNv0D1/HHC10lUrgt1xOVTBO7SAxrGzX0Xa3eXU609ZEbUleme9OaKoF
8hYtiIyUqrOxvkrUvPaug+uE+8V83s60Rar0AYDX+6T1vJ0F8YPfSTDUglcLISv7
WyHyuJhexZGGfqlI1LpfU9sq7ZohL8JBMrP5CUu2XFvNlbutYMux+Lqa3/qca5lA
Cc9hoE88BkCg3XG+0ev5iH3o1aJjg0IYPZyEpkGKtV6wRffAnKUfqfPz6gGNIbar
dO+gzv9XO5HcxYlBsWHbGWqxdQLqji/hDEH9U4etu4Ibn0POLud7Rq8yYblFlMry
C09qrT4Cp9YWfhJgMaHleiH7MJW+QLYU3eae0RvSLlAVgmtDfmX71ONL3CZa9WbS
LuWxtHW8ljndFTnQXASN8loxpGFdLvVnwIiVKWZ9xAo1w823jMlcMMugqwmqYphn
t2GqwpNWkg6t50y8dbzx2550BbqqDtVLMfJX3U303W5NVq+fNYVPJgxAeoW0t3n1
xI3MZscAq2Mk0ne37ACWqQnwer+37YrbsyeB8h0ntNyS9Cw391F64SLUKOrEIn4B
Ga7SsF+gCe4BbrZusfwCvIY3VMKFu1dnP5Nvi/HrtOjaJdasJnf/oVNHMW+YP8Q2
Wofe7LuS8HZ1MaErVkRypwo8jf2Swbx/O0CIAS4kL41nZG7swQuMA+yYfDGQC1CE
kDwWDQ2uc+WvV59pficj2WipERScOdVk+7FEEIDJ1U2DMxnV+pN0t7Oj7Lq1jZdt
YAcRnfzn6YUb0ZHfH+xVMAFnvSWd4lUoDKsZ8ICWcAyJlOhmJUl5Xe5Avz7cSXS7
CIV8ZYfIEjHeKFuHns63K5Eqa3e883iHAG6w8OXkYVg1QFdmC7WBdeCMrCk65wKg
4LKAVIfOoVHwo0au3EuMSu66WRjP/K3EEezmHwrl+3iLcquN3s6W1C5qMZ9HjqUL
fjP2zxvqxD95WwTOT2q08Rf+fqqPTx0lwNChFdKOczA0eqTLCHOArX5Lu34fdZ9P
vYAydu0Gqp10TfjM5F+wddsaDQW2rEZGdBFVEq2y+5rA4lR2kDCLxSwon5h4u7Vn
KVsm2iqNsUJ4lpjDbkcAxKPObRNklzVaoZzDxuO0X0j6UmmflnVCo67RYFft/h6D
ZJE1egcgHh+NRHOuZElVN6tpRLFbFsrSV84jpvp90OwjJAUjxF60UFc5EgZee/jq
sGex7SQQSBK0sCHgGpPgQIFIEywEv0t0Ra59E26s7pUte379ho+Ok8XbBD9dZjK8
Rjae753i4BYe1ZBFYqps3m1R6CAeatUSNo2RGM5X1VTofb1b3I8pUXGnRXU/5rkS
Mr09C8Gk/vLhfChu5GspYASpZkfkrMXMruViHh4gB/kGYzbmZ7YgtWCi3g0Cc6wE
/9KpEZsq7S8AciPPicnTGOVSGtIVszwFErLByqBb8qe3RHEDXbkzqtlcvJeIRicO
cBlP42cPXOWDqTrNw7qftYiucmgJD/BZ5oojyCqSd/2RDY7ZfQHuWrUx3rbiswZl
KPAZbwL32vPkqevIuIA3OjdbWG9nRdJS/QeQA8KNwoOnoaAop+xGdtj+Y70tYa/3
q8jP1B2vWt7T1W7qlNEHe17rvKAwM35MqP5fwHW3RtDXULGah1TfRJTm7uOnlMeT
qt3fE/468N5pDr2l0IPdX9Jh7OGys5mKHltwLWT8PbkqwJ88tqYO5gXA5PFZ0Hh6
pqDbd5zHLoKAGQ65VEd6VchA2VTIfKzLPkhWsnfIZelbX622RaNfQ9dYO55/MZU7
9KNxNMKTsEOZHb6/NtuCjsn996pUtvzKKe/vaTGR1ejQGsj3GKykVolSQWJopyHv
cVIm92DVUI+n9ujiHnDLMd9a2blttSs8CZIhExNE1dIG6szZ90OMzzL3nSa9TA6y
6g9S//iPdOlvDyYu4kWhmbKdhBDKfUCfPuOMXar9J5nwjVcRj8xLYaBPi++LUO1v
vwUMB8YkZpixcsX4NYDa0JDpw0J5xHh+RkXSoVIL8/3ALNlNEFGOJgekt+K5dPs+
bHbLPGtXIIOZWObKzAHyvoJBNdznuWtuF27wtWLgV4Z6irO3BZc6Kr71N91/XYVS
qqZvkCQCyVFUJFhiGlZcSneqkbDKAhY3a42FZSBCagBxTbObGECREzT2gV30+SV5
hA4du6ledLFLHTso4aYymGlnW1N/rCOkbgd7moqzqHjo4T1XqNg5TUySZG7UT0t7
UZ00EQJ9NOUqfBBJKN6S0vlymOroUSme4hRy/3ut4X3Lw4rq+4K+Rid7xZlfrQA+
/iUOlBk075zL4RuOgkZxG/M+rdz5elAJ+cACg7QPUaXm52sa/bLwdQX8KxqLr1N0
W2C2bgnlccwcUk2ATixspqdNSGH5M7b9agJwlUtc1tx5VfjxQZtmYvq5YGmxqaL1
qh85atyUt0DH5R4ORRq+g4sfi8BQ6yOTziGxTHl8Q0yw779+Y8acfHks2x6GeEKC
GNW0OA4cxYdQKlYd+fYlMl9BIeV3frYbfOsoK9pOc0zr+oZO6qeDEzZkK3UUJKa/
I2KMkTv0cs0gud5o2sfnMW0CEcbtr+qEUWoV3qf9DGVmFkjzL6Y9M9El3LJJmpQC
neY/zQPodqvze+t5rXybT2lNoSRf96V0FKze38KI/+ybvacl8vT/PLRs98X8ASMH
pV0qIyiV89mxxqyAGoitkXKwYBSwc/6GHa2afzRDNpYrGFC9Ezaw0ua07bljrrVt
ik2ED5g7oeOEfoOTOZcG72QxFqo/zl9NZLUnzCw6Q/Qx2OTgVbHrrsvqOEdn/+K9
LnO/3Q4OfTbE52oWFihTwXO7/Xl7XR/vf6KkMJ5Ypl0eDpfzykzfLa66wT/MT4bw
QPk9mcd/YmjqbJyFDvgHsHYO6EvsC9Bemq48SdnXNJJHPfKhrQvAto3VN2r1n1FG
FeQ7DzWFL/Y8bWmHNmARCg/J6+30LRxU/qJjCREGJKpKyWn619LBSYZQOsD3a1k+
8IsHTFOb9SdzjmWo9ZA3JowUD2pME2aaz+Brx9ynDYAw1yS+KNb0VSCKE7YfKFis
W1rwlXHrsONGIQhGQ4NWFBfbZD1+am+m3xxZH0zLxvMOHF7Y/O2kdMojCIynBGY3
1rroHnVlXWjJdJPbEMSfz7Yb41hsZC0BXHfe0vPpR4a1UW8pA/IqVTU2n4hb1S3L
S8xbpsSwk2cJ27dby1eXydxy1v3TH1LTHPabHeN9yiwdD3kIOapdMFziO2V9I1nt
kJt59/o5EyTgoURlOdUMor7IhSjNtbeOfrmsJMb8ruuXmTCPojVzyeJuP3pAMPmf
tbSFptQPivqMIJG3VdYJ7h9d24cjl69oxZnc++SHwtrh7kq1KfrKSKzpats4EsHy
smY8+Cp/5cQ4DrOtXZmw8bORMnhIaOISkyHJjCYzqAZ74thsCa1GveQqa9lKrdS4
SSQvGobUu4wOl76zhOmKOn8/9r6cr9fyJFxUpfjg6LkbWmcOWeiJV28dYJ2bDQbW
HWiGzDVoc723uYH2ZuoP/vrF0NHMUlU8W0bORNUFwbiEqJKyjKqiZYsg+3YXzn7q
TW1oTbITrw2B9RMYsYbwRJNKn9+del9kDp5AuHXUkZOTc75nkcQoK0ijh2ch1kNh
ujqsvNtQtrGIEzbm4CJaw1gh2ZO+aD3SO5tIIZix69wB376qZo3uTrh00hUS5OeT
Nlx5oB/HSYVixfva+5OHO56ybH9xY4kNiH481RtCrZYWMcARAZLjMTV1wmHmTHGh
0Jlr31K3yESU7nqmoypkXFyekAPtIYIVkv/gPVLZt2yeWxXqEpzCm6SFfUcXAxAV
fp2XkldUs1gbiyIhsc8/1tkytBfjJG9gvi5LOmxbUs55u2nM3reChUuXD13OXwpt
dItAKjSdN2WgEvaMfdduKmcTyG8F4kiIBfiQssbZU4q1ISbfv3XlkofOCR8wg8jD
/hXNaczS5ODLNBPkqhmro59vgXrJwaqD5uF7czPZ7/ne5rVp+9ze48eakREc5SDh
QdoBiC4zDBvi0ef2lAANiUbrsdf9qXZE9q/feF7uyd8NFzbiV8nvVHEYxxg/JDzS
AtmiCaZ716j89JQbEkAJOog5MGW+/sbXjlEMt2XRNqG6Sa/IKRVDu1QgNn63isGd
QQ1PCY38upCsTXt+DJOEO9Dw8gXEO9i9J0au7QMbrOWedOQwpGnUseKbqAnZIxdq
CWGZ9byVUtdbArmyRI8yT+HB0ma2M21a9Y2xTV1tA8eOP6NeO9f2W7x7XpH7U5hM
myFUesokVjJjEN6kv11RHovN5i0GoHCSfeYAiHfgQr8xyR3S/UTgcJNCwVa+jxYR
Ae4bKl8Qjs7r6/7X7/nL1tr5xKqKmxfkjshOkt6UqqaaFbb3Jene5gxr+15z0B9N
cKj95UBkNU8QVEjMkRNAN07pnHVspj6LcuEc6uGMV7C2xRgaMqIuYETUKefvc+Zx
yrdrhoEEgsCn1wbksN68WPpKHMA1lF46bGoEWp3s+W70MbS664Dn8YkuF101HMsW
+STLTLwodhjPqFFjODaQ/GO4Zv0Ysr/lYOLAubWwie2abJHLTvvpSfkauvMpfY8N
YYWJzuJ7de9+nqhsVYUGvdz8vHCLmlBTCDXFmQS7tD4S9vYYGjmBAWvQ0pDeaTeZ
VFaIl82btQpyxWV1lu0EkUVqE3A+NOI1/posfRjTR2nC7Ojr1vjAZHmks6dmRPdM
Vi5kDC4HrHIVEAi3nLQLqrKebHJuv4seEJBmzGtUXuZgb5yayMG408GQEi9DqjjR
oDNc5mw7jH7NCMpjY2I1yzbkbUuQzH3AU87HdHTKX903CyjqpEeFWXCBu2L1I7/z
s5r9X0vh6KwafHHLbMQZeWzTlhwHarytZr2O2iC/gekrhyVq1uSWIauuWXQ2jLfv
xA9/v1CYxOACGnxSvqODDdRaKzEYDf0ouOwJLbHa/z3pKqTuigixEHgr9YNHb/g8
KWnmo++Zut7R0Y5t53nGMgQZwoglHZ4CTXukXlMx5KZkPYqeme/fhZTiHZHLh9i+
WWQJF1BSKSzNaR6SrlJMrkeRMYKXbfCGbkLAK0qoZG3coe07by4KmpF8NsSVor7/
g/2B1SX8fKUvu0uoqf463jrSsnKnU959HqlPJjvML+EOJBeEPEOkLp5qI9Ck2dWT
90EjtJP59jic0NgGxSK0ahpzusKsGQYSvF0nUtbTMbOcrSXw7NADRxTv2gqbAC2B
sKzX0eKtJ+7y3pgTSUou7p/vccKexDL8PTXT2n5SdADShf7F3KiffW21hchzjReO
AUSs8ovUoJXyUq3QgRuKUArfn6DKUYKV9J/j6wjoo1wTLC2sk0gTP81wPAcUnNaA
NtmCrfAVgf8utOS+AVLvK0bScXeOO9rJP1/8tm5LhB8/xoiI1D06c+yEL5POmWfa
l+NNh0dyF9cW3Pi6zlqVUiZifCJJntUeHpwS2FVkAeLLzuw7p7An6Db76/wOQL1T
MAe0uz3FGNLMHU+c5b2JDfkSKTrj2C2viE4ToDXW1iwj//I/zMHrwdgBITb5h8jh
c2zzlhl5n8TM91WghX1JN+e6+aRPcQIZBXIJB+nQrQ+kUYc9BBx2qumCskfSnUUV
PxhXRqwruwNIcwzDycBUja8b/+/N/vHYl4H7vJCZGrhMSLgSovKtpgpePahKASJT
jqrTD0EN3+udSzinapBKrPSO+SaBaMOuZbd/mQKvDSWo/XQ2qfbYCk7crIaICGGD
jEr16IS0E/ZT7dQO+jl1NJaWrka524AeavOgYNKB+GBv3c8hWohunqMdclOHmLoN
/BiPeYyQjti8/E8NGl3/O1qhiFNn++mOI5tip8k7FtAp/MjGygVCosn4l8ncq9K3
GpXl5TosKGVkqw9/rcUiaCNZ9NG0IsqqtxyO0cdLI3F0bw2vjkRyGSp6QGUlUPfD
UACjh2zFd/eitJbNVA5eJ8pBep3q1W0B8jzRU7375F/f81r2XS/slE5nIzCahUsM
NbcXzFKmD3N4Ck03gEGc9axLC6Gc3vmIse1RsSdIJ7JNui1Wkj2JkZOWSC/2AILD
5iJ7zqzzxpedacF4Ealj3ap7A9aAC12OE3S2ewyM+c57jg/25jfqCgNq+IzXJwp6
SqNcXB8CSM4u8Ewk/0G8pwUBeYkZvldikbLEom0NKLFO5WSHa/TRbmc2G5gMzKtZ
XGoFnduj48jL6DuXmHytwlTjMyHjfN5ldB/XrxaGsBu4tY2vy5j6b8LE24V93P0W
/dHRG9TzTeQH5otHIOX9p3qGg+HW4DeutX2nFk6MSN36E5LmSXbLbbadzeeTx/2P
XCfyfrUQQOlHBwjBE6143CPmldCr4RGyhQG/Zi6CfbyP+1pc9b/DYpzq8GQD+6gw
uroeUiHi5PQSCs8dM1JQDTPfClPWkUYxe7j+VghbROnHKQPd+FRCAUeum7MypMnI
4JqWhE4M/DougRmeVVcd76s2lQss1gsmpfKGG7RKDBCA+4Jab8WacJA2NjJQ16FY
jN768HPwaiqf5WODx1LycsjR70bfzIhY2vpg94wkt83yyqc/Qk1nwUAXidS8EoJR
tp9CQmvgOUO58dPq04Mv6igauQZZE0WApTcNzvlloGeCA+uKNZr+sWLgFWY2yYjq
7UniIoT5Gs6k9KHTCIw9OrRNJhRyhsLlpR6mL5IMN8n/jpv5Jy1vrrOQ3TMCnVC+
mv3wNeNGM4fjY80hbixRibsmc+CBrcstDe/FQ51KswhYLKQPzP9yS+nMmiIFeLwq
NRkjpEwtE5oKsKnSRzh7f2EqUU1+1T1z1ekLgVsajuehyoxHif/LsaHIrkmTGZ9w
6+wbx1l5E8IrEqioA6vGAMgvbUqShib4iNObqwft6t2xgdMFJOUvegege/BK+bwB
OKg5eanE53PoIyWV0emkPpnKejKP/AzZi4IYwFGa3+ihm756cLkLzUpaXSSKRFdg
or4KOZDM1T7BMJUrlRsJJJz8aAPCVqoUR7KpyyxgOyL2ywSBhFG8gss4TNb8SyxJ
0MAffHU3PrMZUII1vhok6EzxwpfcwlIhGxOoxSRPpqofLhqFu2b/u4tzyOgdvsLp
wFmqyXuZhfMQZxiqXQ+1+t7TsXZSCiDibPtbUg1bEF6JUO92CEnSBs1Shq6WdO/E
BS8o4Bkf/UVTptFE78fijUPfPPpyC16QtspFWMwWE5Rskm6JuiSymYIDKefOUuqt
1KwYJh5HB7iXXTLFzj56ueypFNf+fXHK9jjXaQ1UDNX+ctsJGsYNctaZKkMfN/SN
OZsURxLPa4FlxAfby6vd7xHCa/TV7GL4pNFDYddqpgJmr1+Fcd+1RCXvkyd2HyMw
dMI+978Tyq2exjZUBTQO+jWQtzaYCSMr5H4VYir3ccuZ3z26IHYdjqahBj6l23wD
9O5nOMAXlDlYy2voZkM3QiF/die62CExB6jwtFGzGFNFHQtpymRJnFYNjulxvo0S
n69A2Ya06rsZDEWr3s23YpwKpivRUExpsYD7vNBBIDVNq7y09pEwbadoaeLzhiYG
n1QcqCG8vvrABrWgtgZUx0xADdvNYr39ZLVc82Ai1yY7LdENad2GOkSOXRaNWMBS
tWzsBcTQk0l4sqAjj6xbsDPuXvS+SQWmH37T75OPs52CTT7bhE3gy/t0Xu9ezFNd
jJdUptPmHPsWrtZM1utWSLhKTahS9C/HDI1eOJLfPaRTPLAoOQqt49zKBJFkHxRx
nO+68VdluQG2fO2K1LnK/MIY5b07zbQdN+JCiNyKJZAIFQWr55zKOtTxBGilaJLR
Y5vwrF8EC+mYqzTwBPxoOy8SzaEMfhBYbaoeA2bYF7YsZDOm9zuMNyYIcJ7qoS1U
OJaIlRnufazKgPc8zTW3Dg2IwxlDC9F1sC7lFKYX4POuy9SG6z6Op4stw45Qm61q
TaVQO71+YSFHh9JoiO7cEBRKf19r30c/NPcwP4lTtR5TIR2/65kw8uuSxdbGJvxA
S+lmDSoP0z4KnMyOBxg0xwVemoxEcEiRQ9hcKKfQ1m3K3FDfeFMuWe5isveiCFz7
9EfmrlGG43//vxQQmomDDecMQnNnS3EhmxSwzoSd1S+waXPPo5DUf3jfxD8Ijcal
9Hdgk+O+Ns7JxGGoctu6e+LQfg55T4XsJUG83Oee44aJ0c8FMqi40DbfcQwZ/6n8
BTC+275aYi/n2YUip9EAhLxzursHs2bVilcIbPpWSHJ/COfM1ivHhGkDeYh2prwf
VClbFSDBB7eKrx2twDw1wqunPEGs6TjWj911rDM9G0lLhL1JPcI7hGR2NgAYMVNM
d7JPpyuEzCJ+A+TvU/xP8R3UAkQZ+9+kR0b702DtUKENt2j23el12mF67LqLQU7h
6TC47np9hT0RpvMhB1rAcxKz3uolTZVzmn+aRZA6JGs32qPpRk0EWSvQ2FdljRdp
bRVM+xdCcP3vcS3iN93eQlWo1jbgvb/BQRKP14DV8g6O9SP3ZsjcDM1+hmb3uZjf
J8Aw0pYUd8S5nSarqHkb6KdyevAz862VGRwmjcs09FMXhIkeppkfGwiPA+gFAx5I
KQehjtxxEWHV2o6lk5ZUXNODd2gCzfMJ8qmuqjMe/sv19Xqix58jKzecEqUzy1I5
eUAgSidGq0PGO0OGfQibReq+Ow27qx1txsmmx09trhm0Bdc8uT3YIqxaS4NhUlic
xl3PGT8lvJqeAfaOX99JltFf/G/har0TKflPT59AP+zj5NRcKYrXdEtoISfASPMq
O5TuUCbL5GLv4kfapP/kuWA0gdKoXIQgl4+iyC/x4aNNCmO03z0HL3iqi2fx+Fuo
1g/18wGnhkp5OkhY2++RqTbjUWuYE3nengsghafRbL79LOqUPibFftQne8mti7GP
MS/TBVDGvJYI0dWFIP0ydw9OcY4f9fueAzkx9AXz8uamMy1oWRPOZIOMWQx8wNO8
15W4KEWGi2WNx5WVu2AUgMIXESN3sQqqsqS9JhkbCrbkcjFgcJXAL7Hm73fZ9dqL
h1goZFeW5nHkPAosRYjn1h+RflIkE0JJz+es2iBVO8dLcoSMWVB0KnmgKItPEqNn
4HePJoGzLzi7f8uX/mkEpn0g9vMmpubkT9+SfLVkAV1BThgR/Zi0Meu4q//xQ7i/
vLu5iJl9gKVdEmXooqNMOh3Tbu6Lib0P0wmhi8WPPoh0rm0GqtGmIlmHh569xxln
I83tBWH1K5c6HWY90uXCuNk7EYDpMFhT9tPTByaKQg9iWXU1I07kEchkNsGKsaLO
t6rVq/D7vaixecO27ihZz4rFRqd3u9KiLcTM3jNnsCIbdTaiGQd2ikM5OXqovf5j
BQtN553mx/FNEl3WN1tEXDUUFB4slaQKO2JAGytHXGo70I0CGfDmvycZyTtKYkVJ
Njvmr2uDUXu6AqFI2yJaGhLHwqoXhVycwLSq6FuJzqdPRvw+nRKyfh1CjWiWYO8Y
N618T3IoozHYsBys4s8rhNjPgN8N7wvPyDKncofdaE6vU8Zh+PslrLYc5SiiS6Fe
1DvR2gIayOPDLghn6o65f4HcO9+/ILToMI59s+EFVKfiDed+24WXMQJZmKzprOmg
kDeYbawJbnRZYDH6gWGSBn+hJOqt95oirrGbTXxVBQyhdqI/refdc4x+ihQhmsSn
Tjb4q72k+3sPtgTd9mf4dNefTxaeyq8SZvWa2CaQfXsex1iI8HddvhNsRmQkxmQb
WcCAH1GIsgdPIr5JonIYfr2GLEQJPAZnNy6Xxb45J4NAXHnlwwFPJy5PjGtzXe4E
3b9b8Grf9bQsCD63l5qmBPf3XcT+LTCVNbAVJq48QjCRulG5H1ICeKyZc0jVfp6h
uVVSgqH5fmgBUoZua47nP5aQGLtxYHwEjHA7XmTfjo7zIvlnxnguHfioEUR0N0Be
sV2vnDETHHselJKqesdmfpX2+nmS9dc1FajGApKykzjGUBsUio8X1Bz3TCGGq26h
vK8qZixi0PAoH/yg3sLq67FtkIZK4VSMDsYchhkX/DZtwtNEEye8x9/O1oeiUeeX
PtmjpDG1Rs++RQjlVxkcIiX0uMD8Sn3zIT2x5MZ5Fsz0L7z0y9VEGKO1AWoCeLQR
9y8tkbuELlf5SbPbOdoWtBy13VYS77rslpCu/2xXKrcZqIQuPfhwocIR1CVHKkNu
Bj65X7vr2hpkPIA8DcRuCwIzAcY0XVwSBuPaha2dDxoz018M5FgdIipbXkx1WDwq
EqY9OTvdoC1G+YnXEMaIgLld2zavdd8cDvObribDAYbgd2G5FSis4rtKVCTBCNO4
0GwDFERGhlV5vLuGWkKQeM+z8xWuZte11Ho6ej1VGbNNxl/Ug8Kfeb63OQl8D+Ky
vBvlfXoKTumEa0lqe1fACdRJc7LfH0VabzgctKdDD4EFNdFEr9Qn0zvFygMVSZPl
QbE0oWtrmRLHjo+NYbvwluQf7KDg+GNTA88l6/sdOf4sUMWsEsE2xaiyf0mWUHb8
0tNea3vmVPz6a6MOA3Q3uljJOl9xbRpDK3DplVqAx9EHJIaOe/xKF7DEFIwP1fwt
KAH8P0firVExLp6cCGXh67K3CtogGpOJDFxnOsHVMS+GZAo/6y7C5xmVwF2GZlkN
xP9TaEQNZW38NMsl4INM82YBCqeziYtmu/PZdlmXjJAdGxaF4UzFsqNzzvCwG0Xy
D2x/MSseKWvaV+XBIaj0bIqsfQ3sPVFfefOYaRQu4NjQi13y5d/o7Ox5JQpwxbKP
SeIfLZaqrKHuA9mMLZgC1bfTVUvGli0fsgOSrWFj9FRSVjZIBrvfJnqsur1quCcV
9JJqFtG15pVkjcuAkVlM2fGz6yskttxtvXnqa1TBR629VNPCEEK47zNjiiOHqQAf
eSp/s8eSFr0KrfkSGaAnYFTkLcOb9QuE/+bxbDI0kSlLSRArR4bPFT6aCNKovhrw
9a1ZxDyN20NghBtAm17VhgW8OPQz2nGFha1zGcx4fap9tbbGu5I+r85fqx/bcRBM
d9DUEL48mrrCG6z1vzlQWfz9RgKhHGyTh15UQ2YV73UcApMGfSnc0DPA98xApKpg
dzx9U89aywxZSdl/SFaO7UfX6YxQI05HbQ6D5W7nJzcDg9kEianI1h37sQK90l9M
Hi9XLhDth4RfP+UAPQezAs7LN5z+JizUJD8DlrGCwIvIHK/znVlcMmQiJqyODB9I
FO9rcgEbTZ1fesxxcAK0ZCubn+YWrzhs0hF5eXQEpVArk4eFjMek00xzFUu6vL1y
PPR/S1CrgZWHUHvVPtSoI/gjSxWo2IDlI7JL8c3BcavMhwd1ZgtsGPLeO2soz+5p
ZkiNnS+Miwv9/7iNgNdFNZng5Jo+P+EHpHqvZ8WOn7UV373RFqmEZuM/g7wY9yMa
XHqljnzOK+gL7RsnE9qawKp4zphnZLU65QPeMyfDdcm8qHGsPBosTDzja27JNdMg
KjCCHCE5MW+dXUgKagt2yR8HbDl7cI95jf5myAIGsYauV7XSgM+MXdhzO25EBwuU
8iFhsbUhgbt9korXGhVWTTmDDelYI+yEp1Wts4jrHrLu/nBsonWLmS/roFJxBl3H
dzsgPloTnX15xcPt7Pme6cVd0r2FK35wb05r+Rox+V1vKYJrITGLZ4MN/3dYbg87
jasXhW6siL+Qrnn9NyGoR1vXM4qkTo+VYO8K9REuxK8GY+ONK3B9fbCBvbPSbmSK
HJD3RajgNESGTpFjiS98TGiaGvRg4f+vUMWypU0mguO/YDc6Ng1GgTYdtdFPt8fV
yzt2t4ylj3DoKTWf101smIszyEEPx91uzWMU0o5XeS0CWkDXBbQRURaFbgQddlH6
TL5KnOVuGQFt/I2WUO4uINeVKk/uSjeoTaOXobwGxzZANOA6srOD3cpW8QNvw4Pn
w+KPI57tqZ+c9xR93XEe8gcM4/kw+vhk5aFcsxFsiIjKl7JQKHsjcdWF8ouN9r8A
FgSo+KLfPWkiutOyrn8b1T9UKCzm7W2o/7NwgvJVxjDisal85jgyj6VmUGlzBEvr
O9oUaaB53cUZpyRYn7Hmn4PrCp9hABG0Fo7M6bOdNUXfefUOZzNPPBiJQdzEHAQU
IEw7/+9AiIzxZKtVHFoGpAyQBC+PjBx8uXDyGIjWIbJj0FTE/ITCnYHrULs0Cvek
9rKOLo4KcBQOMFKTpejlzZmhVWTG7DNiAgAwuZByQHoCFMxxiOSBKCmIoyPz71AO
4203ZwNlHH91ShzVLVUZ3SUN9bctmrGwefa1nFa7HLWScIF9qjUMRZ3aiacgrygV
X7juQpZGEI6u1x57QXbSGfRTMKM3ng66oRSiaurMZYfvOYUj+Z3VmSn0LRa70rtg
vd9/mNGAu+MincBgvqFhJs9X1JDLghfTZI1D28sMAz/norxv3R7MSbEiuSJHna4a
I4DUxEDLxJ0yoEM51fXgYbtED8fyrPEq6r5uDWX4xiOZbk/mM/VorPmfjC5mun3W
TAeJOk/Gfn3tez4aPz6Dindciekk3pkBjlqivSOd77I1G/R1dvcGX7k6qpwDKRyR
i8ViApsw3LscM4SO6ITudrWu0EeJRcvDUuky56smclXsKPhCfVVOl/1VH5ugDgZN
OXHvjuqgksv3cJxZa+ghBzsuSSewK71VHY6H/6AZP15jzPw6lmo1iL0xIvaqSyFi
e66P0u5nZ9KehDwaDe19JiW5LAbBz/N51HXzroCeZtr1x1Kz9G3YuCOXQJjMnzsz
9qBdqO6M3BL8wKusZgWnihJfNoULGIxG8gmiRCkbP/RDducrujE1IKjZ7G/RF5C9
n/om1tT8GQxHtqJ0L3z06/Zu0qkzsYC9Gz0LHSuXdn3cSzhktRposgFe6FjUzDdd
9paxYXxdpIWbzcC3va3Hx3fI0JgNoPl5uhZV/kpCSqgyjGbrrlLwhH38+aXw/HIT
IDP+yzwtNep1D8beVtWx7Ilcwlch89ddj6wZkNBWRamocOwJchBDGPgI2IKF/uxB
MjA8gIeJpdeaWnRPKgkCqnf8AtPSH2j3NZIKwH2k823PM2PVAsKBFlUkPqQWBQ/y
75K3xPITJb4JPAYMxZ0URN5hZujVY0ASX8JHmVWvmfv8/K8pwppGWBtROzgBua3B
mwIYcflPtxkeQNjRUhIxGuc62rSPnRu3OY5Zb6ZI7DiJvTjKpYD4VbsWpMFwV9Bi
yiwzWsg2RNAtQz+/a+crzKi7GVFawl4J/vbDIgYWDJgYSyrlsh0Tv9i1rPtNa6ks
Q2RY0prrNwi/jmD9wbgEXOBhgFt2nYgOXwBRU4tdfquQnUZ6cND2qa+7iaVY+Wnz
zfHMWp8waa6qw4M2aYTqjTn72s4pvPm+uC/zf6pMdoFQkYEEAiZbIws0pIzTXnr7
Q3wJXpEy2Tvkgsr3CWDXHwyJtdXCJnDh6Cfsn7ydEyq0CSeLpiwURxEExypmoX+x
fKFTUszs6w4YmS8rYtSIYTE9w8/D2fqq065kj09qBLRJmVfn1xI6AEhFsehlg7zO
LB+OVfGHdMBSxJJhDoaHPJz5o5RakKUI1lD7ZbfndAk94ZCJx/3gfwdP6RD3hNyb
MDZva7ltShmfIRm8mCwicVyrdd0oUHl/bE8uwm9XJYbrfj+yQeCAyDuwWHCGDFtN
rzJvGRo/dcMtxJSdK4JH90B6YYdYK5PudCtZPy/ffy3/mX9aeflrvDvoWGN30Y5p
mGMZrU4X7Fw2D/QSCBt5nY8OWs498mb5qps8rAqGKa9/VkS7WiqHk4hS0CeYgZT8
ep0bPUZrunODeYeSXC0Jxv2CGcmrutEQtcITRz+Q+3Y+qq/B/IaTmpacdS1llzQJ
MTXeMxHZDUqgp4BPrfJKbFp/RyuUT7SoAqiVKlISBjuaxvm90rKzYNYanJHwQlmu
vfD1H6K1VLWYgZpMSpVzXtmqTFUbpReMrABJp8XZ2//Q7hDA+aE/ykyuHUciHy3E
GwHQOgspeBQrezkRqc5W9uDJJObQHXzjQWX0nG+Gr9TbX85XczQPdYVM1qpn9bI+
sf9fzmmAUZTqhOMnqGxyi5EzW/MvnIN+q+1PtcIoAYyF5Cy11J04IqrndOvoL6bF
q3Xc8S76TTLvllW6zNDfldsJ2vND0rI7GJPoJDi/b8G19PaskX2Eck95ySYWmcbq
lKxLyrRQlr9rVNUEZmeSjigcRdNB5TSj7KG0h1PVF5EB62mLpla9vez6bSgOV0K/
z3h2fZtXIkykacPKLAWAQqGJcr17fb9KUPA9yeLD//eqNu7h41c+l1kED+4a6Y3A
uJqjIDEmPe8VO85KEe+5CgkNBlE4xH8X4cLXhYkDQhY9THWUR7J0z2zgpuSze7af
49g6HUJhfRcTVpgOB1BBHbViT/n6ggPotKZbXAosvNZ0cqi+VN0MXB/L7DX5t+2d
NoPgJtqXlbhLy7AxzkO7+h4TVCSOqaWAU/ds22PKEbVb7F1JMel8L6IbNvdxFRec
sSn0bDwiClQjrO/JbmMDDJF/QP0xTyriOD3D905Io4r1rN6d5rcNcS+an9PCCP19
AVtmXUdv/uNxVd5zREbkzfBpAVVfz02vh4e4efpTdkKtGP7kMDi86VOSEPmtekoK
dcoOzeMnN0CVEbUqY3+c0u77BgJUvDUfCtwshAM1G5oBKQuHh4q0yuE3jisIne3k
YXIG35AAxJ1My1KOreeU/WalZ+j3DrTczLoEFMFPpejb7C/MQG+/ZMcTcAiHnM29
vlDeDr0AwMzVOSXA6NX3U/TSc+2eSlNucWBVEtyk2yLyE7AqU7CdKcjb8+B8kBNg
vCiXMkSvTk5BU2yxRbg6JswsgQXHgkfQgG+4dTrybPOBhb6YhsImIiPwbrCX1s4E
9H+Gta2U9pYeTlOLqGjsOqMcOykKo+qfkxk762QMf2QqVElrlsLTKtLB4CJG1VFa
Jfx4VFC/bwni/qs8Z0oJIK1vYOw00a/ibDtKGHR1omHcZClGuF9r5T6BDPIeSqx4
jT/hvlz72W10ZtMn7x9RSgeOqyfqrf17yLzrrkHIM0uSaJO3yFQYkLJjMQqrjDhg
jgNPLp/x6L1TTFzES+0g5iTYsb2Tat3MoxqJEAl6CNJTtg0EA8c7YXVjTduY1DXa
Kt9KzamTu6SK8R2nsRQdBdd9qQrBzLRajEPRieMoEJEPzhTTNw82t8wgZYt1e56G
JzDa7PBqKWL/MoPCb+kDq4aC1Q5DaBbl/vHudRQ402RES9gmShO/HtpIKOodwCQJ
L/6hWGbewtw45JdB0HxWxGt8tHlMuF2Kzgm3Y2Rk8psbSLB9XBbKp1RO1+FuHaQ9
rwseANAl4PpReDE2k1KbdbfISoc+PuRyr0YTlc7y+TW86Ye+h3P+lLoro/H1It98
BMCTk9+b+vNEL1CYEgOZ6NAw73AOvBwlukslt7yJOljQSGT2IIwxb5souMporMnJ
aQPpr8PgKcXMGAvlZ3arf/9DaRLqp/+wgetzqV06L565zoMYxxcO2xQmTv6r8d9U
RtgXCVZPGjzzgMZwUeUd6/ooL9+e2d4+TSTIvHKu+HpJy9K8mzupOsGs2wW6sYuD
UeLEVztLdgWEmSMa8a6rMs5rVW97z1GZeqyVK9ndh9YPcZTMjUpsHpMCHMOtMu7C
S1jEVoGCIlIL87ZehO02kHf7xOtzYhlN214oPXRWq2a2Nu7yi4+nTLrsIZ34Xsrv
YXpKxX3nqrKukUC0S/Zhtj/M4Wvku9hodkFKJut7pnwK8BudjcadgElX77Bc6aHn
n9BLxav2MFB8LgaNewsLNTc3Knb/7jNkCCxBm85W8mz+iR6qPOxsl13TqWKfhUqS
2WfwRQTcxlTHEb+yidaiAXR/P9qpPg6NJWzIkuKUwOTosK1oBmyLF8nTBTI2NOW0
+z/dszvskF3ViYNgX8ZQNkxVsRoEJCMSWTQwRydAkDBZ2EpZn2cszWK9w60MFLSb
QtBKQNt0UrxELjkvdPXT3id0+qQNtJDvydzSJkl1UvtVkf8DYLHPcHjfh5sknrYI
SH7kcmCUg2qWSUI+B+BJDiLAw59Ki7eKJuUXb7n6eZrY5t7YVnWChwJSSKYYCOP+
7yossDdJ/Y80yYeQYGXHgpbK723vfR7ecvIy1Pp47FsFTiOvyX+MKtV/D2DnMxP/
R9q3CY7SFgs/BjpmXGkeKjGI22rMBjY5BuapsibS4g7o7GZeyY/QKP3Qoh6O24H4
zra7GP9W6fM8M1jURjzFspeHl8D4XH0X9TPixY5jpSLNc1+ym7Gu6W+2tzoC23tn
VoV0ZReW2CiKh8kYUKocBC7etKLdGIdnnvoXf4/IDen3TtJmD8pQtCRuA08CIWyB
LSijzYKvOlT1fyZ6mXdA2JmIB+N+3cGry8cjp3jGX+h5cK3X59lzsbtV20uxql9l
/m6eMG9PY5p+BnvIJBu8u2kuCkgWI+uWhPpmkdASmT/nojxxc8X3IC106tZC7JO1
9+/uNHVl2wCltz37ihEFUdAwS11D2DA1FDGBLaJozfnNlK2DUEE7e2EjPy7OjE4e
Ebnikp/yFJDqR3t0+jqogbE0XEtSJ+Isf8GJosFUqx2jLvYiAkwd5ix6k/Q/DLr2
pOwzK0nyFfj1aoSno8mLYLgiJFygvRmuH6rru/2W34rPsYoiBNSYNEqliVD0eHV3
WAxsSsfQaScKPiKeZe3Au5Nmor+Ep2nlnHXUQiEaPn3na0ZaTWrXL5YiM9qRn2nc
BIAZG/dVHjgPxHcf9Q8eGtlR442izwjM9D/PpoPzUU3iU676cjncuC8JEYLnmnng
Ze0MktebcrZ4OVBVzRgXTGNDtIohVcTghlDchGmVRb6NB26JTC4PKkFVeGY747Hq
pM1J0YBB6EGKHKJJmTGIcOj04KOfn8SEmblxePZvtCPDsyiXgKbRy0GCw0JNcKF1
AYfnPtDPuAAU/Pm8tQLCYe21QKA94PZKu1vBs17C6mYUZkzdHFFXETGOHQIBSA5/
u/DwJBxNOvyfn1oQFtAx7F4qV6HKBYCpbpdD4JY2wwbH83C38SdCyRO3XDQkVVZf
oR6j/E5hAqdWPE4fxQDytPi/vvheucRmG5KqrD9DSVJHTl5OQBI8YMkx/R2L1L3Z
psS9A9X1/nTMtpoHjse+Vn1FlEEeCSmbUXOR8VKQkWSz+cM3HXT1At+7PSXeRHhw
RuXWy++0ZNCT++6/Ducwa296vpGII4JvWUoV8ytDgM251mVADEXTiI9FRdNlDuaT
jRgcLk+dF3/Gi4POYcRdasyL6JNcZJ1yOZXOTRVzCK/y/W9gQ2dpL/eIWyAksW/C
gkFx/+CRX8yr14v0w84ww/34tEKGm14Y8DZi4YcY3qV1f9SJFQ1s1gzA35wrm71t
re4wM3o0cbMLndZ9dFrNC+5ilt6Ls09taIgnl95yIX0W0lheEN1cGsfmJOV+Y+Mp
QL6JoDPwrkv8yew+t/tX7ZHRUQa7ETPdZZrXymScr4ve00PUOKaT/2mma1AbMSUD
saHNws2hc8aEBPecZz3p3ELziG6YnoD7RNFGHIumiBNhupCHaYBeohdfVZVBcjhv
vuYXQ1g4Dj38yA1Rwh3RqxbcsLXlhAUcTP6qbTRl0kF5OU97pLPTrPqiP8YTD3A5
D0Cx/KWelXYpMnPWlteWIaJAgrzDBbmOVW/IaOh5iGx3cqW4UitliVKYW/wpTHxE
kPhv2D3My2RPrmp2AKMtgOKxAetGPIh1JqT2JzHvFhBvyIYVKNE8BJb4sA8QAzoB
fg7ZX98Vt2ChEfKeeKbxKG24A7B4sbas2ekLMN8VruC/nCAGHMTLpoT/CH66SSKn
Mz2kkfU3dqY12YIzkJjlIGx+fO8sLM7ks4QPv/Axh1D7v/AEJhnNazHnrI8Gncfz
aGnOXZdx8LdgySkj+bZXBha9jZOppHHYIB5KZt5PZHmYvfqdEiTvzL3yr87GLKsP
pHbqcUvHUuFjgvJll1gZPGgr42u2Cc6o4+tpu/C0uVjDnS4lTAlWofY2xaDPVYpW
Sh5zmYEuCrPjhkWIVgjHc6Agiabn+3st4NEQSQnkJLRNwYTJv+dem0x3gXvDjaCg
nujL27nUjHGRWvCH7Fe6bYrs4mXjj0nc/zd8ao0pIjGfBNf7PMwGvi0yuggEsgFZ
7H7xyftYIWxn9O1hrChS58ZLwDolg2XTUds1pP5r6pO8dufa/GUFkdOoSgNlszKz
97/y5jdg/0j4bybMEsfsrqtz0D0THlEmmcuRA+ASEs4mVPgCbxH56z1IYJeXHPuL
4uq+MCdLEhmsXZtI6PuvZWcIkXS5nwwy/AStgFBQ2UQEKEe52NYGinK9bplEpDq6
+tYHfhGX/5IuTUiKseZ3Dfkq13c/Ubj7jiDPtT5XrNuA5LRWkZZ/dJE+X0lsXlqQ
scLO9BWucBgY/9RzQme0gBb2oyN+Soxt3HSAerAIxdVPBOk/Pmi78hDYwxiq5P1c
8qJmih4Wys/NjsPAtrTWgzBIEcR6hz+2zlum9vxy1S6RZmOTwZtK5itledL+NMZn
ozmmfeG92ye7GrEEBPmGBJKS37+BkC2oW2ZIA94Ba7whjOVVStwLSxEpHfoFm5T3
pUUeFRMecPhaRZ4k8KCAfQzckCLO3/fiDnNdcLvGYDLP6lXi8Yl0ct3DBTvg4k82
LFbzmiQ/O2FO3qjPiZVCg9PJq7sAHtFwGN/AO3XQblE72ITuEdpAD07BDZyzfQxL
+UynfzazroBwiJ3h7jOkY+50chtOaSC5/G7dO9UYzRviZeJqVNypnFppF9IE/Pgx
zG9h4U43F3BpaPt3wMHf09XnwGzB8co9FqJRie6HyYVweBL4SZMswWnWelMnVjcQ
R9QgEBqWu1Vp0ck8/vZ0WueEAH8Fz+01aheSgx2+ha6ZpCCmw+7ILBo5D7a5lKle
cRRNgMFS6/intphB5XVwDVMABnYDiXvr0sNF0/em5MEOFfzX/6TvtW8SapLNoMIk
U3JPBg1haWphBPJ0W5YdAsrl/4dUKy5vNqA4HBa8f3RFdzJZoMaFI19v43tsftnc
eJDkVbN6OOJDNskyhUKJA1HCyrj8E7fdm4Ng/gVegZ4hAVvh8Zr8uSnH8T6NUXvg
gAe/j/UvvKxWsTT798UwCpDp0UlToqIoNavzP7bTW4Ne6B/Iq4VPtaLuquV+u0OL
jODh277UrzqvwiLkZfWOekAg6gDbUIcLSIo81VjUFSkOC65gMH4TIGGnQBxehY9U
6TlYmyVBrVKIRq3fFHJ9jaYtfqTw6ONFroKbLgeCmKe96Y9t2al4ftxJZ48m7Dm7
dlpK1zkyLx5vte/zKS2DodGwe6Ex1tQe/Ex2OyBH6AaQpui2l5f/6912iAyOgQC+
j2dZ2L+oPn8sUbgkwAez7BvV85q0z0Ns66W/u24UK33WDOJ/q8EFdCzcrlE+mhdw
X9oKMU3LTcAfvi2YZPegjmwVzxPnqZjYLybLw7dqv7qgjooLhHmYRMVl+6pWAjXV
0/xSnRS0VBfHizPklJmH0ZtcfmHJDIUDWJPiiVzdwLcG//UM1YTzNA8RM6HBwzvi
Iv/Nz4Q6q8E398l/E4bUNXWDh/H+17x3VbjqnmkyVooUH03uKs8yezuqkTbnqV4G
nHoeqQp+k0UURSbCUpqWddvPX8n66KeS85w+1BmWXxbDNTiU731ZRiCdXhydoy4h
dpPP5JNREbWAd26pK6SJwybVt/fO85E4QTHtpKDvsU+5ywTgOK8gAprR/1PzcaiT
4yTgcMwfSHcVRJ7d8/ivsACYeyhWEZjG383hJsKgQ2Mp90N439PuMPpBkzNiW+nU
gwTNMlB39qXxRcKcIw5SCDRC4yPAW2Fc7PEMrs026CDf7AhMCnmYH1je7eAeF1CW
vt4fHrmZ5L4SLKl4YO4s4UQFqyjG5PUbYJ0G/yGZbmmMZD/6pcapbAuO+zLaKAsF
3u/mLlks1SbQoGewRimMTnvT0nJIXpya9l+aSLzuGuDI9dyOj7RC7eKQpj1jNQfz
PCHbNUK1s+qFDmqQncQp7S4zoZL0/c3Iu/AMmQpvZUQzZ3l4At7V6DHUzz7DKrBJ
szZP+NbUs9wjlxf/5MDkLaV3vCP/rvMdffsDLnUGUSNkD8OHLooTsX2PQ3jg3jGo
BQ8KhP2jPOWcI2D5eX9wOtlxg8MvrGzwLpHeSi+fLamLDAoimz/UGJRs945dDw8l
sSDbVy/kto5FxGtPUlGfS+ZezW3HsxIjIMLTwFPH/tgjK9S17XDpOSlMtvZRQQ+v
hM12M7ioahx96FWRh6jn2MV90zsVJNPQuYXDtQ2fMxoafVtd1HnQpVxRQiCmc6In
2tS7uf++ETo8uZ2lO7vdnk5eHIjqRii69phAPbjBkN8A/geyF5w85HTH5BXUDIA2
MGO3NSOd8FbT2SqW93e7zUEN2W/BpPjqbJzF8b4mpOCn4wJ1P/LAVFuuPEELtY3N
7Dr5K580WTE/1EBT3R20ODSXEar9AEoG4jD9cF5JtlGAHgBJQuX5/MTxC1llQNhS
+O5LiMVHxLqlytCKV5r4ghv3kBS4snNYwLx5LP9P5phwRCQKjcb8Ib6Rl0/IPwTc
tHn8bUIMzFXS7QTzVkFXvLO4+HeVZvy9WuFLmxKb3dc58iukMeXdFpk5nsWNIuvt
JN9SK1Y6ciQfMB/9wWq0qyskKisnV4Wd74fN6MVowK1ciF3MdjWyGL/Ivc/Jtm8I
4CQVSw8CUTys2db97P1Lar3ed1bJIW+HpqmIAPkwLJ+xykSaC877/LKGWMhZfova
53p+/IE71S8Rzo1LMRLagqtytC19HPeVPah8q0G6rRAMvIuoYmS5FqIuKr5Me4zj
zll4Xa4lg8i8GbEWtefrtszwR2wG6TXlUmPNrFYoPpor28MnWtY5kEN0dWmef/S6
VphS+2hzQvwruXfdpsoNk4apjC6rR2SFnx1RQaOwhq92AyvEEEs1Ge4P7LqU+imi
Vy8hmZm29tvA8OYyUjqc0SV+ljqM4dfMKitk2eBDufphPFkavEcgb/ZKslhWBVWL
6RrcGU5I/NIxYhosearx8yptpgq/ehKCHiOLu/sAzvg5bH5dCYdDa/WWCYAn0/Ry
6bYZWha2y5Pnr/xsueMArB2aRdicIcHzgwawa2614KJm3WGrRVsaizY04ILEBSXi
vesVHCnzJGPq6V9xhMdZsrGcpkZ0xhUjASvNIZjHQVfdKPIAKlKIOrxAP3Eisd+g
/DCsIS4zEC2yE83WjqntHNeHbaeHd3qA+vt2ybDyP92yp9Ay1RUhYdmKAVkeegU+
f29PsMbgLzj4n7/DBKTGzaV5GMGRlvSYn9ilP/K9ORd1R8uV3eDZJt1X5SJkdfJm
FtBtVpw6l7byFjaJYxDC8qp6T/5YdFSl6UsLya97p7XMoG61+EexurnbMOCnKheM
Cs4CVJe5LuJOgaXHIltVmhwoobbenQ8j+UTwWO7/f57U+TIhuk4dq0Op+IJ/VYQd
t4NU92A2ZKFE3vQgt5456+t3ARRxs25bkyqM7j6FA76aiOMLIZh9wYhoyVXBVMgK
GI3Pmq3hODtLPruXSypbx2g5EaeZ4Hc0nnMqsfae/HxevKL8R7n8ywuKfzefsfpk
/+pv6tqROdeGnZuwT3e6o7iuNjq3OXd5VmiimWj/p30zuUcwyeT09CHGzvbqTzu1
O8IBtYDZ+GtX5uToFj/v3UcjlyKmXQylO9SZXi/PU4JlJ4k1L5DhArfaTmnJUN3f
/OouJk+7YsPenvV69iDydbmkD1+9dXcAQriwGJW461KutUOVqVwL8/Sx9kRynqg0
S8Hd8LE+nUAWa3BIO7Yd6GqoAXgbiBQUXPizCn9I6nCHcKxY+IA/5qkxXhIOYPH9
dQocc8ZyLfB8jgsXX6iOSlR/EL/iyhNnwyCMd7k1yAJ0os9WrWXvJQHzLTnGanw8
CbUIb2dA4M25BU+TWZ17AAUgovedaCG9Xpfmzvdy4W4mYARYle4iiIPXNfp3jO1d
PXgrc3gNOnNAWEvqEyIblfLbl1iIZgmMrXE1LPG8dkG4KU7CKgQ+ErZb/DtB6D8W
0sFifVVcAC6XcK4yvb4ZNHby1F+SWpEHjc0or8CbKm3ARzgq1JIQeF85065G57s+
pCjxDE29B+7AyxZRUjRm2xM0vGtwm/Q3fptioqkEYFUDGg7y8eoYlPMBjoUPn/23
46SyBsy+FdCQCwF85FJwKzOh7qotEn/PdCFLSldlwGYBa5GWU8xwPaUQjk+7SjEw
4u8wF++La/qeUK3M7+xez317ehRP9gRyjqSnuJ8yVHGLBPXASfpqALx+Q1OZLJu+
igzC7jwQrEkWuncCcCdRdkUnuivf1HIBdOCOsOPXLhYQP+SlXOkMjJ/gAuecYF1Q
C5EfjPfVaZBTiwExd/LM0PBMRVoalv/FNrTv7akmpz332kR47PjnVp/60SVxXO85
mb2Ueg91JH1hXRG1PFgtapDoYdP7DecXtCiBplVM5PRY/2fcu+6BjEuG0dnEghx5
TsmV4X/9PQ/SZUr5yHzjnUdONN3GTRWMxRSwD2+7KQztGSSmoaCzi9hnLri9jGlu
/OjOJVcTGBEI2lKKFt0RiVVLGWokmkvIDhGKeqROl1cuKvyhsvR9ocxZ85bFeXSQ
ZCDnCzfnPAEfAndwZqSqCpbtSyIxIuXViI8QO0tH+P250G3x42cR8ykfq2mdNw7i
uMSCinfzcA1p8FJsGE6xAun00z0eauXDZL5VpQl3o45wp+33PNg2e8KqNbUDkmdl
M4GetUYUI5nYQWHpppikxvmikKwM1sIHTRp6cIa2zOCTSL2DqKGsNEldhvZe2H3j
qu0ocF3KqzcxesX5dyoEg43B9DpnZfoO2tHmHGO4LVJkyIGZVlNCMksqtwekgWgg
ufYj+FSL1F8ScQ9gJzzBpbdsMV0kT0Eb36q4qJiWx72fs74Rm3/Ij63bSW2geDVi
1BFs010EIvB2zJmVykLp7eWkXrSXx2CGeyVTeae2giGqdGxMWM9PWlgaHcEMNnDT
tuXdR/0rwLGLMuP3ah7hY/Mc6CklccGhYyAuVtsg9A7XaDH1vyyIxRDlh5ZrY1pg
ejz6FuJZcSJ8UhjZZM1GrW1Az23WS8P64o2qL8UIrqIGPNEqVmz7et3bcOZi7wPr
aAZNa+qBjpy/4TAYv7s9ev2kO8z8eE3LbZ0htSTDrTt2LL0pL/hzI8hQR090sCrP
xYKyrT32PFahNga3qDP8tGv7S1VDKJghzv4r6oExtjm4qssp0NBYbmafz+lGSzLK
frlc92ROWnlVfEIDXkrxI7wTwo8qxLw3cPwzwnU9OegeYfFlRrFiR5F7JmiHIWh+
x4vUNOy1tQMgWzt7FFz1Co1j1Og3IVt7K3ysOFxKGL+oqmy0/e6Jg+ZXZKxK9Xmt
WWlv6nCODPjWzni1gbsE7Z72QcOOEnqoERYXXR5KvxWeMe0FTzVIRLDcMtIGnSIU
gQzKntgFSC7TfwERb3ZQoAgmuIFUjM7N17XKVU661hr/y8x6Y9VSvvBgyv2HQZgf
9iLYA5DfYgGY1F08zFpa/xnwEkvsZrBRG2e7kZ9+DvTOiDMmwuhIRwPHMxys6Lmv
OqdnotebBLQ8+tCsWVf8Nk3Az2TPKdO2bjmGG3IdOH7NAcA7scHUhNtDEUVoeEbr
OPQ5cYVtHvj+s/yzEM5p5LR1TSlTmNwsGBH6ouo0vvbjRBkcRYbjkIGIOKbn5LIE
X6wTrVodQs3C5E+HzRfkQw+/HvBqlqqJ91jZgmT9OzzASkKHDHVKuWWjW13GdrkI
4O/xzXcSi5dJfsc1zmWJOW7eY3K8kuAvoHkQJT+3Kg8juqT831/w/e7RDPJXcVb9
cbqRBe/4Z4l7VWqvGa1/B6akzvknnwfW/O8m9S9GqSqhsH8D1bwcd3wmgptXR+fI
/l1MSRr2Ml52L0Zm+6AfLJKxYEMLk9GjHw2eGST0F+bJx/fNyDmzHgzP7jV35ZsF
rQstuVQ8acVYrQlajbxcSZJka1eFqm9qI///aDSdMTGzwUxAgarjEmYXEge8k8v4
Pv7InmiUwp9yPBC6J7LTl83Q8qtN0fPBcmeyFm68RXIVZGJ2dvq+HhVcaQ06AAHc
WPLm7a2d1D1L69xK+Gs1gcIHdygJAIZgJDy8Dxu/6m6JNIF4wYj3rX1JfXJ+Zptp
yns0V7UoPjydrX0KLXbM0rzNq0jLhOhoviA5dOp+DIbJO+PWpjMITvLoeZt8JEle
Xm+LF0TQkz4oVqPG13LSUp4u+lLF7JpCsXd/CJe+sALRsH8pFDTWh24uiv/Al5Eh
rftSLE0NjctnbwqT94tlUTyAWWm1NfMKTFyxDT9QHpINNX0pagGnXGljpXwl+8Tf
Ja7cbHlhzjwqc7uRqvlP4ihSfnYRMjSsLvA3tp3LZ78h2EKpUzxkW9QMlKYu/+VI
5IjpAwlXSwzX4VKt7eWET0fvLYkxAyP/7jJ88J8MCB8ZcU6oy2l+3qGWtR6JND4W
q7+LoGF+gyhaiBS5RoNNlzutdEcP0ptj5+CYD6PtJIGn6955YaTxSfs4FFCK+shf
hj+2+bpBgLjfX9eP4YC3u8hM56zFOt3WIHIYXwNXdDogDfj96qjfQ7atJD0eKGjH
OrpbeSlBoemQ86Gsq8bXh5jiogLBKNMZEYEF3OrxeROg1EcvgdEaPSMrsCOpmps2
ZmZEnGUUI43jLzMqiGkasLn4ILSHERHRw6SH6OW+mI0JPsy3J0cNzFHIuRWWT/+1
tM4t3OhBsUauuuaaFEvfyrQUt2VMPWl+20eTEjXcR32FB6Bipz+QWUWHmSSv7ops
j4DnKTZ9De+rIaDHilvDBq9LLIYAEZGgNGm+iEY6CDmMZKd39JKnvPvcruaLeIJg
Rua75hjHMJRJ7b9nmBs4deoldugdqcM9UIfHUM1f05duvkOKr7VvlY1RqvSgy6aI
q9FEWrWJMQ9jwRzQHu+qI4cObgeQIdIKjf/JnhRw9mmG8ldRGUipQuTmvFBQnoHL
TpFg3r4WtT0TONnRwv61LG2j9IAhO7nT64gm8CpROBHNIKB0diQw1p9w+hotG4lW
yGhdc6xQp64dqREV7tii3j8OUn6/7UZMAmn3rkvhzgPIUqkJDzuZCeORiVYL6aPL
j32ZxJ5Uspg5vgioDQ08VoSfb+A5SCsQ/I1POVz0GaMxdu20SjGz2I/gSluffuKy
M7QMGzHcgA+tc+loKW1wVCFcFwWX8BFJGZH3LF5vUWCWwol7L9a5It8E57++IWZm
AXKx7UeywL1VZFqXqHuO/dy5kid4xqL7MQsvq1qeukjzLZfM8IN7Vo0tWtLdOw0X
lbgfHV1yvav6d4rXB26VQx8SMzknLM3mNerNhkiqqlgIFb6P+/reifAoDcGzbFOh
mcXs2e+1+tIMAfvnu41yk6yoayxGVZ7E5slzg2f07biE+HfA2swFeHPuHYoByHy3
6iwljT6lqlHxja4naGYdvSvR+joxldeED97lvpy8NA/Ii0hT486jNRAsCeWdb0lZ
tK60kUZ61spPWAGmVjFrJdPwZVULMLpQA/O7sG8JP3XdCglx4qnDcdb8Y2hy0VSS
IZSzNZa3icZ3/CeO+QK4LJwrcJxHE8JfacG0KLwfRqrBQiMIvW7NH2laW5rywxyD
U8I2e5CZHHeboM+fQTvVDE3noomWmsUUcuvN2SemlkeAj6MCHvLatQjDZsi+Vgzt
wgVsrawUwOi2XuXgRz6gkRlqCawxfpyT8EnTvMz/arQv3PtBApLOadsHyqOlk3FR
g9HyF09OEwblvJj8rNd0eHEFVtFeucsp8eYUiLdaQxSPM6espgf4aZ0ItSU4YXEo
4HirS/YkS+6m8Z4V/yXcR8+el7jzsDXbFyOZFyTPmNDbdnkSqDQ2V9gwzvasUtha
04X5zD3DVZtQvu8G3d8IEA1fNWQjuKE7zGuXo5B47lxrVS42PChRVZ/omNfJK1Wt
tgLYdQ4aejRa2pByp4FuiDNVsHThZWIIhmp+Tiwb4ztqnBmduyWDZ/FMRT9K4vmf
Dbw7A7+qQBpKK/rzo0vCMZP4zEj2LXuhU/NFD+yuJwIXiFAYL8QNHgVBWzoF3aA+
pjXzVgbl9DoieXB5X1jbOOMChSaJxsdt/lhuWHDNceEaSV9cKXmDSIPprOjX1b7P
0HzgZP9LeM1G2jC1RpT7OhK+U5sV5TeEYSZE7Bl+NY4L0gGtRd9/dFMC9aZb6am4
PR+yLfPTaSKuGs3G9twWHIe+O7VmlJc83/RRKwp7JN3y2Q6Nj0+w1cRav872pES4
/0sHBah7gpF/i99VgxusnV6MliFqh+xNok7jZYtlJFBI5ctS7ISqowLgjrIePyzR
xwQ+4nFERK6K5opA1bsZ1SLCgOUh9rIWmBT+w7dVG0Gg02AhOQdE3iNkWapLzrLe
8J6xKRxNSL2gDIpyTO7Ol/5CsK6mVXhfBpW3C28LQhmkbSrvqAhl/vYFzcUZYcJl
3f51QH/O1mFiyk2cnTNz/43T/iE4U22DB/IbDKcioIWgKRfD4CGOE1LxXDgOyT/B
7Ok402JiwH7mLFa0bGcPQVoW4GO/jn4VDWmKw+u7TprvK42qBrqcwibWoR+0MDV1
0zvJX+d1gckFRDxG6ndnscQedAdKwqxCniufRNbG1rcl7EM4G/QKiNttDLmGYWvp
LSmJ6+YWbEjIPxt9OxI6tMXqX5CazXg3jITq4v2npn8qe2S7M43u8SC+1Hs3RPOs
CKN73qJIuTGCXyrcGFbP7U6iXZaqm8uRELFhphjkOdg3EPTcXIm3V/NCwngEaNzj
GI1lt+IiAzyUgUHx+3/nEW8ThEiImPTj8NF4f1+nUWt48i0D+xcWFdoXBpKLa5WW
ngoyPAfFkNCA7j5JguLUf8T/FkpeKztxZNkE0TaCFS0TbmuGkhd0fFx7tjTlwTxU
PvaWz3saXoWgiaC10Ta+S+lrRZg3I6YPSHRgnn7WabJXlbYKKGBGAQcVjsGuEd53
BF7MBRdIBuWxj7tyhYifhuSapkqMp3d/CtfCAJONspgXwEyDZKS6rH9y3ZubbxVz
MdVvRw8NWMETTBNlvzORrjB0DUExiYsmBnCn/Y4Gxtm+OWxW2IaNJZRCZMvDAnP6
3M5ra4ReejhklLHuGTNqyApRSCy/cebv7sws5y9B1sJr18cuhPlndp04pGZpapJj
RnM8bPHKTHDPa1dZyn4LcFPhj/s5dh9wrn0HXnVLpSZQViCkqKNzIK9M2sYeQqNE
tpZAmH6BKtdVzRaFQhl1YNbwtuUsbTegN+A/1ELyMmqRDJsg3eUXWA/vDl8LFQyV
pgkifSBkvr+7WM73b0tK8NgQMqa7mCM6SVDs+emWNW1ackdw4SFQu64ooVulyZkU
4UpASPd85swkJD5b9qjTUiea/c6rmd0BLxyOIlwe2BZ9h7Y/Y+14J5CcNXpmp8FU
DLO6U157q5fcnN8H2LoDGCre9JGSFznnN1Lzy19tw8FJah7aWlF3TXydqNdKASeE
+GpBPn0sfpX/ZpQGwULKT1vX4hSj86ybL0IEqAizZxvlpHDgu3wcv6IvTave68Jo
tJ8ber8/AFMaI9D2bV3Et3jO+OHj7j8Z1n/c0U3Bx3ZOZAisavBNbQDMVW8EkPu3
wXn9PqViIDNw7QYmP5snRtW+h56T+kugtZ9AgFgZrkDqqZyK60wm9hECohT2Dtzk
ChYRnF3Y55eMgrO4zmI0k/pRKSAVdE6ooD1JHi0SV9Dogjr8u5yAFLG9cT3YMYyr
/Wm66HVpqP9jiwGfL8I9eRKayoHH92hu9lI109fBky/EfZgGSxKNVf/P4lb4XDsT
da7wszMcCRBzTj9HuSFpiM/xyl4vynkmLD4AfqOmaul6Z7mC3aGi/EwXcMkdtZSi
zsqSpzmvMxZDQ/4wnMSqe9GyhHyBjIGnoj7lv8m2aYRdb5GH8o7IWffIJd78CDLh
rN3jPxS2Tv8gdX4i9JaYb2hkQswL6O0V0rSQ6dmfDrJl9xSxI0vBy+yInmufbI2H
tOjxF26Yz6SVMFlT2u1sAU1XYNQc5GulPGwZLa4b2XlaRez3412rhRH/dCZG9C68
UB8nHUhSBHwtW6gr9LMiRbXQjhYtn7j8OTcQINwApvqF8PayAmKEVc9oAtts//E/
+pUVZHYL3uTPgIh5/NvrNyaq/NtTmCJE0Tfh8FnCSd1h4C068mpGNDi1Mm8Zrc9o
wgzsEolf8q9hn2vbqr7HRlqf8CPz3FmUFr6kjpTTo2YUvMCyegIp9EYyD0g6/P3B
5KMymO6GfaFdgMqWXGqyBGvS2g5nDgaR6yT9J8rKN8KfRhuy+t3CdyLb5zI680Hv
GRixTWnzsATTaF3UrwAUDHWnky611ibHjsOB0pLL3MBjesoqlqgMbyD0ZK5hecUC
3zKDrXUSmnz5L9eTPHHLGAjo0J2IvEuEC1fuspvaBjGmUkjfcWmkBgM5oH3lrHNL
nTW0lOmvPl1Q+MSl9vuP3PbW1Pz7/yDrzk5S/QSCmr7NU+NysVO74O7r2u3KtM0A
cjJaY1bQ43Kqk37qElYed+SCYCbcCrpEoaSSYdMcIlDu8AIk5SswnWYslQiM4Ec3
QuN2oBtJly89QyGmFGX3IHPOIAT97YlstmE+KOHIAOXPb5CNqfDUwA3AD4IsFxsk
KcS9q1Irqe7Hij3dOBfiv41kK2P8JJw/U+apYq2xoClWZZfV2iJF74hMqmCbkzgB
2x9OpQUY6aSEq9FsLtTptl8uxf+8kZSGWiOFgXglaxmCbhgETYAyZtAN2coB6Oxn
PyoYL63xvhT9tQjfUFLnyhWamlpFt+JQG1ozsU/zZuVMEmA7Qtm6sAzKTmcwbYu2
yLrutNJ5ZfLMBTRX5lLicVC5rT1pqUqT7E1a1qAbxQ1fnI6Va3F0gIQkBEGkYuEB
ffvX0voUVbwJVsgccFvLYcsnjVXo33MJEGby43e7MAzmGD5MGFFYdN8aL7IIP4+A
K9j0spBtudEgmKtm8+opzbLCF3+lJtvscBrmlGGPI0mrPQMPFZx4wyyeeh5PKmqZ
imPIY7QXc1WDNf8Z7y7Y5yxLXVaUe5k6n8eHvqY5Ar8C7YTeYOo+HjjY+somRh4U
X7pxaparnCPWVD2wQ6z4Z0qJr9VxUZTozILL8UaccOoi+EfdV31zBfYo8f7tNbLU
ASSZ6l2NsAxB8B9w0c2mgqCU/3wHwbI5N9kcp3L5oV56KWyAUaLthT7Aq5voGqMa
BO0AgPBhOzYD+Ur59TL5ui2l3bTNhc3zPMb+to+CUoA+t0Uu/hrDAYK06HjWTUX/
lPIAGjK5miZcoBeud3s3X6QF6AVN82ELcCrPNbNq8xqNJ8fqjnCeELskdaCfrAj5
v9g9E7hdv35NgBFxBpw0QR9vS2mT7VbSM+010hkZWQM+A5Yf8RalymN0qHfaGJ1p
pIIV5MsG2qF+El4F1/33ISAxBrej7Dpfd1bMamQLTS/hqydqu0JT2dJrCmkWyqws
WluYKWl/vJHvGg2UaymzznvfmvT5w55xrRQjd3N+7VU1SPN+Oux5gnqb/j1Ue4Yz
mYRZtVeF7mQwcO3Mpt2pivhsU6hlFpkXE95uVj8HUDbIhkHVKJ36F6EskUNsrtdt
qKmNgruMPjOD9yZyRHtSTjKyOcjDvfM92LTRUGVCj87IChFSuFaNcZcu6pnZGuKI
6jsxtUriI4mUFJS5yltwMDaKvABnsWXl975ubIJpo6GWwT79Ab9c915+C960+2Bd
VRYZ/S77618IhxSFvQDRTmCYES9wt4tJ6RW+mih9p7pGHgcqkNQa6/D8RPNwQdGW
BRE24v0UHlJRcAeNg6C8jMmLRrSyqHGwSlXeZG/gCtY4N5pqOuiMT5FGdH9khD/3
ab+1F9OXldHpquRKnrRRduOVF8964A2Of381iqvTMA5Y6t4AGW2jdzm7cez4iLRZ
fzg3csxEVWcP8qrxKyw5K/+MEAvLAqhaqztDjWqfzbqS1E/pvvhNbdVFabTQ7Gug
LR5qmGeMOfv1zin4mckPEEbKq4MgUnxPOsygEf7YxsFbmEVNij3T3VEeqzOlLPF3
ZJJ6MacIN1fWASKwQ11K+glUmvNnYILoxW1qPX0WWuHc8tWPDdSyB905bE8oFd8S
saKnj6GwaGmgpTgp6NfpH5F2IR0bg6k9TFs8h34cNoSl5nunlrCPk/88AM0CVGBr
EPN7poiXOEMZdkFWLqfnXvjxzorqtFyHpNo0XgL0yP7O3E/0zAuou53wu9ljBzKa
dkGIQEbKFN2ef9W+isNaB+juBICx0TP74MHEmjFuLJWM/J+cxUyPSODKyW/EKUZR
VsnkMI5EsnjE96wmo6TPdSDHYfajqC7fmx4spnJhjodT2OediXKUSSfwsqtYdeFK
RWeAmBLyn5KKebr+poQyKV/vc0ET/iMfjXcEcUiNgYS2cEq2U/yL4RE/sGd8LW/w
X2zXesB8oUz3hUtuBJ9vX/RQtVk2qG3CihaVEVKi1bAtnV5na/Gd/cEJc28eZfRt
ScKeXOnHH3WNenwWxBgW5Qco/n+rHYVSOoSFhyvhIa7uEFCSDE4lNSNeRmY9wo5b
6skRXnfByrPURaiooLdWdbUDk0AoHPfGWtEMBC5t31BPyc+kbG5cWAuHUgiOMLDY
S3KbPWZyGYc2l1qbC3nJD4d5WJE7c9nygvawoU0KrgwztLe7LiuDtY8T1SuIN8rF
szBeWPRpst9wvos/9ZiK40t3WZacD7vVGoq2NTLfRRqtA4Ua+sRhWWIwAyoSVcYV
u8j/46bCrTOEm48nm53+UmKOJ61FnW3rT9s7eGgP+XNmGmAgYiyQFcj2tZfXdzL1
xOMxXw/VDQ5uFiWxBpjYt1cklOk739m4wFPcZJJw1GMqiwepp8Z/5gUsFLE9+iIL
vxiZ64QIjQATURYOgxYUANveQTdiy7fFJ55XNvOBj+uNeTdoy2T39quPgq4M6xAr
PaqB7BLPyyOojY17XiU2XRwmcy02/PLOdR3778fW4QpIKWJalpx4rb0tjVrsN8Kw
YbwSwW3Mxtg1OsfIiXRPyLN8lB7qY9PT3+6CXY43GfmrwF8U4NV9+p72IaiHM491
xBWGEwoEqSwSwk88HESJg1MuzsThYQGI5HNJ3a960iJGIMIP7BMPOvkrmg4uDQQ2
8vSvw4B7pfWXRMBatl8Dazj+IrIBMJKHdcYOM7mvRoclonfSUu35OmP/rkAZAoSv
T57h8t4tdBjm5IRnApjRZOTAODrSysL2WlWsf5UAAy6HQM4j4xcl5cEU8mofUid1
+Il3bYgrFtFtKN9o3qKuTrSQjKbsnxsAvAAy7dekTrZw3eJvhGbFDsDA7pPlVdLP
9CVNqcuu2N52/NVV7ppPeG4Zg3tZzNwErWPAexnv4Ss2e8cvjquliaBhoBcT5z9x
TR3ov+iQNxBDDFPXpfiFuPGAv9DkWUdq+NQXdYpA2lgiM3I7Bk19mciVhtoZe13K
7NzQO1bJetcapKl5gigVi3Rdgey8LHV/om6kE+i5HK23gTqk4/X9qr5UzXMGYyDZ
6UNabZUPi7uep8Xqwe8kC0IYwz0uI/FCFdDG6QRMsuoz0XQc/4dwBiLGDF+xn4yc
RSObCF/UwLFKl8ZNKWtiXR/s+WyKyrx41pwhoNx+uBlYHKGaV+rVOISQ6bpzhbCR
58Nn7r49o4NQC3LFI/WhnsRP0wKiC6MiaQX4L8bei3tyhto/VqnK+90YJKXU7dfJ
82rRFzkGK5V0yvuAZ4c1Reqxi0RLmupJv8TJAb/6qfxPK3jWFzxEczCLS4WSn4Ha
JFJzG89qZSvJWiyGiIY+IFj2k2M5tj/ykW5OBClbnFuFqSl4v8wU5VR7HM1dBi1p
3cW/b15OkQ07Hb08AtmP0NBjmo296S7s6qUoZXE+t6GAfAP086dNj0+wATnrL1ZT
EnOhlLuEKXltotqF0nd9KRKGLShPH0hp1QeHYZ5+ndDRpufp+qybc64e2f4xSYhH
7MURZF+iPRYHOSPSJigqidEI7v41lsOl3o3w8uvlX1BYfUh5BAnJSQ4iCA00OcAF
nV2313TO8I7ws7fVhMphcXZ57N14Nz0eX2+wom/iDnUSbUXg6dhz/7i+M+NdSYCA
dcV00PswUroMn5hadmcyzt9bl/bkmUpNNXjcfqj2+FVPuxV5tQ2xIXuR/QxsDOli
GMDm1i63TccsPwbFUDFlwcnYbBuvEF1uFHpS/qiVAt0ZnAbP+wtKOgof0F3lpBDh
uYmYeE/p884KuMIFdPmlcLwXQ7N7ku2nFBQMhG0eZF5ThcOSJ6HtvhUS2XlfuV6w
f4f1ZAP35qGBIeEdaHebFt4BVcz/XiiOHDVTvY1onpIqYhVoV/SVemTxqsXfykje
nSQBkl83xLyShtLYtW/KDEpS9d+Es0sjE6bo6QlGFwYbiO+E6WEcDETmPRiAWpFF
s7akSXElEvY8IPS+q9LiY824WGmdbx2MH95H8a3fJBtIjvP+MIIWcM8LCB1K3UiI
VW6il6B86VWh4b2F4xtyToOdafah4HdYFrsMOYm4LqjfQxn6aldAvTgWC2+LS7ZL
SQIfWv5yHFf/EcxaUMgHkZ0PrSE0phNKQUGm9uASL4a3YHgEZhzCMlwEcFFYnOn2
M7pqDYdkCDQB2u6SUxoykn6UguLCzQkSj8sIWrHJPQID758G9dVEK45JOl1am5Jq
PXELyyTGk/IupNGWI1M5IQKIYaeaj274c4U0KE6UOFCB+tbWogrmRhpP6P6+e0li
u/QqrOuJ6neIjGlpLTnUMKZJsBi2nzQYOxNqoi5BLDi9XR2mmwBpYND7U3SvVI2m
Etp/3CHrk+gyL48e2fDDo0zI0g4GUd49DYZNJkLiFam2cEi6Yi9stVGgD38PZ78x
CKWih0kClkAygL1NJzNdZZc7xz0WIlxpBR0tuWA4NNiKqC3mFsWPedKyfBQpu9Sk
E9jfsFAL4DfelG4lOYxXbTFCP5wIynni0HRT9F6Zxx0nN0TsFAlQdhFB+Kow4fIt
07P+74uJSGq7eq5GAGjWeUiEPTiEM4bbhqzA2MgJcyUZYzMXRFz3rlrc+fHvqqnl
yu86SX9gPtt2+rUeI1eaXDhpHkBMfIIS3mn5QXnUzKKcfuLG/gOTe+9Of1q5lCrR
J7YJlKiEYLScG9mOgEUwQqTniYPAMlo43ReD2GR0V0S/xQf4zc/MHmaopiZU9AKT
anJk21lsqxxH+BOQF9WCehX6sxoG6NP9fTAk4hnF4a07VJPhMAyH1EdA78dEElZI
O+PkY5lp/fTQZzUewkLr0Pc9ch+cyrYRI7lGVgG91K8Gl55/drx5I+cHb5MzISJA
vsGdY9H1K94/pUJmnpkVMZiZSmZpuFURIOmmSQZ+1AV7ASVRA58tN7HnRIwe8CMM
zNnGuge2oM23Zj96bJWscKxrUuEwszty5UmhX+vVnHb2Mpz5BT5MLmLe4JD/0Qj9
jyMhm8Z1TiYLAHCwpQefNSDMBtis8hJ3qXFCPB5ecIGWP02CxEyisYebqD7daBLS
cK2fqV4cB9cdhSaNKGmMEqnT+VwZXWWylXa1MtQtANsb8rPzxV39CoWrH+fw3J8e
q3aBPHDGVKZG88yKDHwa8FIZ2A3VGMVg0Nw1APdffBtuY85XZO9QZlM+fEmgQlKU
8guIb9DIjKtCTmnmE3KM34turJ6fL4KxIfeA8N/HRIPo/j/kYwqQ6feQL59Y5Y2E
u7PakD/h8vxyC4nYL/TaFT/KLzjO+UyoCPyVz7ebjgillkV0KlNUZTSw6M6o+r4x
sat6mj/qw69p8jpg6PY92APKv2X93IyzwCwNi7wvKqwtBtcUc6xrdweoaZPxHkcC
3uN3AAsAhfnp1FQBxLAX35/zGC4Q8WSWLWqNDzTCEcFonrJv65dXlx+WEVUL65TI
SAhjYW9yX8deAH+sIBuByvd0xzh35FrZDOWv10564cNFi43GX3z3yxOo4f7xXwfJ
YJ9eWj84i3KWMRGPL2Hq20YbDZwAGBW/L72FF7kdKnbtnIP1O9GTYN0xXEHafapU
qVXwiG6lvUgLU9Zv58di2Z4O7CdEQm3z7ZM72VnV2gY9RokAPWJv8PGY4WmVdSpB
7EFsRteLnYLYcUZ5mzaJ5GaFjwioxqz9HG7CKO1NU3dUkI9nLnTDm2t1ecgQevVH
Ay8IXVSvOQURxocqKhKUTQFhqlWhXhcd5xbAs2wa0c5KMjzSntxhkXgp+PaUOYaJ
Ne6s4cjenqns09a1dttTSlThHv/eKWeW7Si4Uu7DE8ZUXSMAQ88/8jtXcQNdfdnA
tQNhEkf/pWkMyMyesAnY+SjX0rZQwJknYEVJM0b1ig4SqHw6zFD9vMENFNSO+r/C
Asgfyq03Ys3iF2nedu3pauaRqmPZ4N/psDCuwckWR3jHFKat2ePc7JAZWqejktMb
3zFsGJo0hpDm/+cA58J2Uc7COgPBzpfRvSphp17Yhu0LA1geLsQPFl9QB4HX53h4
YWXKI1xxbsRJwVxZvyNs8t6CNlCma5la6UO+eKB3qLN5Q+yKsdZ0brk9cM5xLQZR
MoYGI7Li/n6vcHUrGFEg1k265jjhq33NDqcv1NyzquqX6p+kVSbcX6lT0JPhrTab
lHxvwjHLiBarrITbvlZmBkWVHxDlQtk0c7v/Fbi9LlNZTNxalVMGzQHlI7A2YV8a
tAObVIdQbC5PLWGXHwaMZ6Zif3bp3fqG9QdVDabQG/K3N+78JUB9Yl6erRqLnioQ
zX9bNUxb8oS5wCnpKq3Th+SylpcBVjgoTeoolsL91smMBA8L9hF1J4+uQRVia47z
syW6Og3Sg75YaRohbxvvP5amJ+l+3gfrAEBY84ChKhyVDOkhHbF6dx+W2aexPoYC
+d7n8iBGc8kt5KpGaqBjQNC1tjoxadoU07ZJfzd5TLss9W4zRUmcPu7J4G3LcsRA
upPc8cjwJtVonZ1rFLiep941lRQ/Tz9pGCF4zo2dOCRW07uAuibJWWXLN1g7ZlS9
TmVp+JaubqcN+35EORw1ksq+tQfzZiXD5q9Z65yT/iG11YZOZYQdLnlScB72hSSS
xENB6Xk3Dh3i1jOXgKnsKET+t/TMl4Cz29xyFfjbj5kEvTKBRigEmGuw3HuiJVQD
ZHC+s/yOPzAWmGxIrIOdLrwaiWDJU2gmIJEDnOcd/Fwlxn5NHEMpo8jxVGd62bCb
AOBFEBPR6xE6xcbAsLUSSwroZ1Y7NpfNhbjGw9zh5JckoqK+QO1R3QWDWEwJJcwm
iaKqCNsl6zQMsIyQzs4ATeDCZ2mpbGfmUsVr/CjsSiB8U88TlEf0pzkpaCjYb7jN
YZnkUVV0ETsS2QptyjulnxlipOkqJ2gOeG15RWboeBKsYF2kEN5irR4nmuZgJBoL
hIokI0Zo1q7l1WwuqpyzEu7ZqLTJ4aYsZNkhmiU9OoIlJq8XQ2edVeuyo09dxJgd
7x7Y0I0VjXxktDiqhuib8yftOBGXNLWkb4sV3DLWjqQjbwpfLpJC1kMRQ3/fO3zo
FZxXDG5MQmxL2QKicNY/K+cSRm/jajF2Nxn6G/bOZ00z//1nKHvHhVck5fDzpb6c
f0/oPt8wxTvaru+bD91q3SBvEjIKh6t8XQryNIuTzcy3Lpdq/CrZ9DFqfeQdP79M
zSNDzhu52gJMkd4eovp4ER6cMws8MOPDJI9YVX0Uit8nFS9Qu91hibIEKHk+2pyP
drGhjMDXABfAfVZ7j603IgvU7DTyKOefWaKaThae56WI10wgg2ubXXcWwBzktwZZ
FcXCBloMmKTzG9uocU44ei/H9fcNspCeY1Wykq3x+l4MFmX96bWCcyGfg4g6pNbV
J2VkhEQfiDDyfQCghoVhwLhos7IQXTIFCH1Rk4yIy2TXbVIsdR7OcxXrPcU7xWhN
Hhraqs4SzGvjyACc34w0JtLCh/wp5QokA08Gf+D+fAMEGPIkIx4v5D8kMT4A9e/1
5PGMO97DwiYAqEvW80sjuhG83wu+b0RR/F7/HFWMG2YX7wXIuiy4es9Z5T47HFah
X0FGQK7izRcsYdOnoz4LNigNd5ku9z2N4Cmg2vmgCTJM9fC4FSj3CryQIsiSxBuo
hj72oGo0PQKvqR1WYvl6pwkbhkP5RmvDzrzxt4kTrL2Yqch7MYdut2eiaH/nrAT/
Pts+Banxasgur1AeNVwD3T8PXjV1W2el5/pnoCUa69WPBiTVg9g8VSoVn0gQVEkR
tjq9bp/M9XDsyrBsCFM3P/tyrMJ7Afwjxfh+8K1erROafpnaSVZf7Yh5dnNy8Q9r
H8DXUcG93uTmHhswn90vaRsxHhbyxMCxs/qqVETBaPdDrrNSkfrAIii7wJJx/HS1
9sWN5lelkKeu8SA2zGkPgYG5aZzvbFCWvkD5AbD6ykJK/theJMd/TswUHirvRBH4
pDJpE3WH24O5GTEfTol5eUaxGvDlk/+zyXbQVxiaJ39aoJ2uXcPEfh80ODEROrgK
BGt0w77TrDmY0jJPyWr8r2pEYEJdQ+Uj8G4cFBNu1wLZFOsc3ckGiZAaFxTnGWHZ
YJ+QNTZrceatjLFi0CLq43DNam+YX/l1ftLyChWg/dZMiXuCKYE3znE9ZDNkpSH/
ze7irk0fUEVl7DqLHKV0t5bU8OvDDU40d/20i9rEoKNc6ZP7HF4jsD+5gvIcj5DE
cexykNhrAbFO7WTDyHRAsns2ssocWb1a+oWY2J1AZD8tMiQXrUyZYcaXeeXGu5Ma
MHDGNYHy2W/rVmgS02BIh/s5lLOHjL/NfP7alNovxkY3JC1JWpLin1H+GZvx6n65
TkdcAUnixHWBYHaAzhwtHT9kRbEvf/U/1FWChZjnso/V45DxkGe9tWhqRU6vA7xk
ngqKR+N/bLfkPoHPIRWsAim39SSGV591OjCZg1GWi+6hsVf42BUWJxZxwM2svuCN
GW0FcaoOJyDPDeM+obon4sSYg4P3dPb7nRbHkGGKMZ9dAIuN+RFeUY53EexHnAmc
LQFPHzWTvwATlYmotkfvL/s9rQHFocWVAdmdTdR//umxPbxXtxZMz34dltIvQA41
EkHfUne4jMBSPsU1V1N8TC/LeJkqB6ypn82PnkLAjs9i7z9RYEy9uHhBPR6EbRqb
LYh2EBUuuwWIWvi7sbobRXPhND0p9G7XAFNvBYkDoB+4Qo2v966yBRdyHG01LvsL
Ei7dz2WevKpktcHm28qYYCJ87egO3tR+G9aMAb5NRiKHNH30YTKRLLDA0osvl2oj
4P2UEzrUvTkSrBvCrIsr8Me9JnqxgJa4yBq6eeeYf0XmCAPotKYnpqAaKoxINsCe
ytLNW1A0On1FjZw1j08Rpu/s8f3oHfO3OkP27uXHTTKVv8n6dWR9HsfZjzkk6hbQ
CgXv9SJNRz3WpY9fRpqAuEPnQJZm+oS+wfBj6G8mT7VkpK4/byo45KNp1tP9DBms
+UJL645f12vC+BgyZUZf/J90/zo9L/Hrbx4jB9Uh5mOQMGzPkO+SWKY+OHU7HXUd
INCV0T+HVz+J0gjz3u5KTbtrqlD46rJ35TmWT/vrk2BBk/Pe9rzFagGrL7BR3Acj
/9os09Gfxqb/c7poBaTr+AmrsbTXYhjNdwzExngpasc3fzkJQ4ba+KzEB2qTMHUl
ommuw24FitIm3LmrYp+bhE52i7/UASkhX8e9h4q9LhBSaeIHh8X6xIMAzKCkWMz7
IXw1EjnL4J9GaPia+LioF3S8uLVxcR/K3PF6/eOGfY2rAcJUULvoJX6HeUDG7Wek
ZV/HkhPDR45NllZFYde8SbpcyRbIPpsNi0vx3BTKzCvp/tjnIzAIRdrXPZ4SjgfJ
IQ0lU3JIoimyCTIfYTXwUK8n1S/09VRQ0WeSC2g+y+jaQS43qoUgHriNHvVpQJxM
jPHwFpmrVwNyto579TPvk7Lda6evJNDDcSrqROMlj/6H34psDOE5V9t62fq2GPcM
gKI2tqUCqaZQNaWZtB2vWG7iHyrsRYUZqE9VLlfOtO7KqLGV7RNw9+jF5BgvjKoR
qq7ZbMO16Q9K3oTKUFK6pIwNhTrh/H+axpvsAdwYCTvib84GSB2db4XYJQEsneNr
7wqf94CxRWC/fubSshdp3KyNN3G+CXyRSEef1wIwI39Qf0Cuf5pvVfdRyG9sxaWZ
zc0CimLw9KVGSTKxCsRB2AcKKTWl/F68RO7/Wdnt8fSKCD7S/qVW0g3iUdG6veP8
H5KEnb+owpejB6nIj6QWIzKXt+pE4cqJTXuvQ0R3ldwuen30hsYrEdu8c3p/YUjB
PS4T+j3qJ3iYvzy/HHLyuMWvCk0syfYT8gJ5rMVJ32TS9RUWoXnDxLnFUQQCHyfh
tAW9360Q0gDU1b5YJ2hRlmpSLA7f2WfioQg04rxRdjUDv9rHubpponkq/Hlil5pZ
giOiYRbsBw5eINlCHBsnhTtHjWXpMLi8iaSw0ua/hL4KGb98Zq6/1i70i6a9jmtB
RwMjLmJ+l/TOE4tOt/mMOe9b2LokK/p7TYbNYOpUmql19n4XWQBoB5uxnpxfmY+e
YSHClBx+F0TiYZsVkqLZzajByqrkys3T335S9gxladtcqot5deIV8nVpfM14zHkt
VRX+QOntOpuC5bggh31NjaTvQdqmQAgNsF0Vvx5QyzR3yCjLVltMdM14nS5+aKJ8
hIc1OoMf0MmskVx/Nv204qeHdWwgnnhtbWqMk7RLIdDc+057QCipXhz369FS0iKh
9iskszjtu1qxKDpwPR9TAzjhDsGOxhE8Kg7WeA7SE6/Q0v01Z7b7Y4rsGavQWSI2
DXPrQ+LPObNmTpvPSdHtYXtGHAQ8cuFZbAVZp3mO0ZJ0bEq3S70wSiBVfhxtrWb5
PsrxaxemtTgx+V4OL5TrSXOOudfDjYmmbnWFbpn4i67TG567R58iIwiSVjuhjnTg
CC/cYs8Db2ofi/ByAdCTeRr7R1CFZ0SJgrVVXwIW9Vi3xn1OcCX/6tyOS8la/Pau
zCoJfkbh244HBmbZXyTRfn2OpWAU4E38QtLoSEm+DbfytvFuSvV1xts/iTTgpr31
yJ/4U+ICC/ypPjzXnZCAaYUqgh82p/2wFAJ4NBnmAku9uV+3jkljbEbn0Tf3VpV9
C/NsnUhr1AW8uaYa0lo1fnrRchMIdx8+XKr3pCqJjhhoKqWi+PHdIjwVLb9HGWg8
zCS5cP0d2rLr9dCG5WkAWIeqqHcbHt7sxXcrNqKkAVS/VLt1lIqKunQ8oqayaTPL
9sYvbu+k8gmVbm7HARADnpRF9fAPpyP5sKBNo5WJFdw20dvMR61mYlV6oe1pbE4Y
ZmNTw85P4PyfcurXd4ARFHcqDagGS95hg6woqluh++QozsydxClUIHeksIEFz99f
ra1XcGWGLQpuNBhsPi0c4qr2LvMqgxeBJUsvm6SizFHp4BgATbTO0aYjLJimrOyi
20bKUHVvIVErIIFZ7EFdf7Fn+9OjAOeLSiRIELOm7xRDc4M/8tlrGA/gQcjwxEqE
uSNg82OxDGSS8P5P8pAPSt+QeXxY6Mlftqg5HRJchdo6BbrlT1tGaHU80o3pspZr
5Za5D1mFCYnKJSJxQEsegShlDpcSYsY5h6M4MnnKue55DTPDDUJZe+9SHELX6thU
UisrFMpo2lAYBFmhMmbjR/XLFzYm0AT9onzvaNl8jz/wwwxMhh4MTDhrfu9LHf58
A/5ivU0vbeMYVppWxINBGTYWfcb3FNxF9crAuQvlzBRDu1/3VlOlQvPJVdJm7AaI
JEJv3m1rK/uihWpakoIgCM+iPI9vqCwYnJ/eJ4yy2lfu/Peo22bObtO7iwsAcnbb
uDDgY4R7OmYytC0SplEr8EOzTYQJynsS6C+ivLNfFkGBnojAVQFNvfam2Qwt+otV
Kr3rUMV6A4hApNQZfZU4OoD6h8OleGSRLRcp9Wg4V4TBQX4Gz9JSh4GgqgbhKntF
7B0wyv0WOaRH533M5uRoiv5qkDlk5W1G43rJ9HknfuMrucKSj51BRfxycBB/dXgi
Pl/DaWRlpSVRNxXfrNK3xFd+ev5XHaRKM1Jo9rykBYZKM/Hqe8HNkUDEPQ6RkaUE
my3jv+fxRbc+Fqi9GyEJQaYkJAtl3vDvTHtZy5ywe7MY/0wYQ6qbCcPO2FK43hGU
Rqs/vnEzpZA8GcwIkWDFnlH0wbgH01+KZEN1a+wAbQoJuENsAg1A0ZZw3LzPBX+u
zOuQ6rxP7nvrJ0N7e0IAtnpBtV4PsqY3T0Y9mZVPckuCmkn4Zi2BqNNpvs1usnLy
JhCMX1kynPePYT8JvBXf+AqaN5JDnJrDNNkMqgs0WQTL2dur9HuW/RmpJLU1Zn47
4wrglZO2E8pJIRJd+k/nvM4KSqn9t0XItYotVhW7H06piWYZaTyxNoYNBKHvBX7Y
q1ku8eaPUNNi6oe7kCHpSQ/eF5XB5M1RWnh3mRiIki2p6no+VN7o/h8WoOYGP6A8
28AARojqwf9Kc1ulpGm306Y6OFzimPutwCV9QQSapoOMxZkTTpI62RUN4QE/d1+H
h46IT2TG615eZdOtv8YtvlkEekoez2xhTPC5rV3UiPZinINm2hQU0t172nlW4zrF
smXNUqbqV4bnGPGptYxXtKEDogMKQ85G3MssuTV8arML3Y+s6XnSN3bKAQn4OK84
BzP2l+Wp7+aIwURUp75b/ldL9HWfmx6SeGzFhSR8EHUk6BMfUbqAttlMwI5SBAbp
LAEn3wDkVEydxNn69Kl3DXX1zWZowAKbQraoSuh+qSOztKsnnBGbcDUE1Pe0KKN+
mGrkFM6YpjcMlVAvhdqt9pFYDyj5yfOw+g7wD8QSVidAqsZB/bPuoTZpBgga1MWA
zeDV1l/coLw1qHOhC+1IL8UCH4G1XQ4shGjBTTfSz9W1rlRZKjtPHvhE/hQ3ICCX
9FNHQhmYIwDd9PHu+BZVyqaFvCTQj5X/BZed5Yoq+m/SMmtWFzoyHGWbNTFDbmro
Df8YPYCTfadRS+j8vSNA/6+ceqezY7YawHqJe+DMzixan6Ru1gohzvd+m+2WCG5q
AvXRtIyh/wmQPtyxp45vbW9San8R6YmC/Z9c+y/jDOMlSWdCnciIYI+p4OrX0Ycu
7WCbuTxe4LHPBW5ZylnR2ZiKOGmqDnHqJmq4ZrUgmri/sKilAAjcHuZE7uyXwUi/
1n6NuY0cIIV8KFVRdfoRa52SMLwHolJK+28OidttHEutZZ68EMk77f5uyqXuxtv9
r56R86duWKi+esdr2Ktu24nazj9tOtKopB1KqEHb0rtzEfi9RFBHb8olhoiJ0j5x
nzsu0zKpyoIeG8EaZcVeLCw3butmFjkD1qitukrV/D3jHJaIoqDV9dZ92UH43mVW
8LVUYXK2iHX5QqaRcOier1gdpPUwuDH4dhCQE+TdluJPf8oAIL2ENAXgEpAdr8+O
hYRnpDjMCtYtUUFghvz/cgLtWYdIMCCLKEGwzF8oZ/K6OGf7KjVJaXCu0aiY2gEJ
AWNEwuTICcynF2LXA0FgTsfwE/oA6IDS0zEPDHPqrUkxe5vvH/tFCl4J9KjbYQ9C
Rd+FmPp5TZsXU7AAZm1YPPBZf8ZojnhUBMF5soavfyespl17qmmdesMfboIWqtK/
MAPV+h64DRPuWvbTekufEdS5zOPFhlYntCmNs1rQVvkr9Xw02mwDQWcyMH9Jsabb
aetJfSxLt7f9w8FjXCRXtC0LDMaU6iDSf2SH6+OMNlkDPXc3UOAuNNL3kXrSfxDR
pVG1tJnK4rh9pr2v0bU467eNoQFo5JV+Y3w+CO2tul/yO45KpTgr2IkaiAbGDHzs
el03M1GAZtJHJdcUZ0fGWcfdOFEg5Wmepa8VHRtXNumA8mH1hh2bQuSS4Ge+fAYI
uLJECsGH0N0OQROv82V2gITlK0CnJEh190u54ivJ0t6DOiEtkvHCa3ZLWQ7Hb8OE
IpENE76BTRK+6i9wmt7tJcaP5O741/JpTynnBL+beEJ3we7o4YsFubCDRNv7J2z7
OM14i0BhLnz+2pKrE2l6lFtrf1SKFw78ENv/T5fxdSpKaeS4XxW7qmpRFo6pKCwT
K40+SX0EXxUfCRSBAGPDGPXNYMnvaO4TmVlEtGfKfi8Wyat6PGWrsyIyckMRJ5AI
0uMd9iDVFtzOs4oPSfKP0ikGnQrLAzURbBjWc8sBykNzfeSkfsS5wGg5c0ogjc+f
cHO76tmFdfJLeMAPyqAXVhEZ2S67p7cRNVLxq/rD7ZEW+eJZ4n9xG2XCgxueK8Js
wvkhRe6xkUJRWT3v8pd5SprW2NC+JnHuYSkm0GG4vvrGth6ZPPrWnJKZyBgRtKjQ
CsK+xCS2ExXIFnQoWSpUoBSjtuf7tv5bgRgo1E7olJrUJWzNpOwf3DZ+qIRn7O9L
wlj/tm9ibDNruCF/Wy4m9Coau9JNSzE1Z+4YnLf05puxY/NR9H0p5S4oewk6R9+f
89U83BKRCo9ZhGqiBVLh29qOAQfGopeZZDu9VOD/ud9nzlYybBbIYkCtvpYi3AIx
of7wOGz9ctVNCNVvu9V/Cy8vMKoUgNe5lN2mqmiTusM+xrwPnZOIf3xBHG44cWjP
HdhK1oFKwi27/DLX0jIb+mhDyWCvFCa6KH1EHENSHa9/+ubWzIMUyBu2JQeLItMs
kWrfu3WCqDzs0RNVIyOmCT0Qk6evRUGhgzQog7A4o4dEC4TpP2V8CnZK70a6O7UX
BsNyjm8iNxoWMZ8hvomPoSG9GK+Xu+6fetZtsb5zK7W/e6t3EqPR0e1uPw1pVlEu
vZDdfhmT5ZgpVpEs2loPiDH2ntT1VZXz4N9Yg7BapTn57ikX9UiKO+0MK2BmeuTS
rK/VuaZaEPkVIAXAL1XoTHhd+p7tNwJLRvusFQB0qbkVRRi82TIbnXDqra+wRMIj
K4XR+QYuJ4hQv/fDNbnK/ymPoUGPkeXPYFHK63FzgOU98zc7AFXzmI56bIPxgDjn
KaLep+CJMAtz1qzPQBtW0mGDRWmiHiJnclp8ipQjxt5tRwcsP7i0et0sru5xEebR
mDiOqAYBXjJ9LzHWMuk9xPLuTu4wSh/r2OHqKPS0aqF0WfhoUzSRmBXV54KZnZ+x
T22DlGzcCwzl7IQPxOCIYZR8YR3gk2bF54y7uU+oBYZlFPm+ZAayIk8TU353QEdQ
O2be6vDNtj25TD4097+XeIEhhmsXTR3uJkbU6uiDokJgRlNt4eHPWTZ43Owd7naB
aNIO4HD6+HggFcAtU89nufuZG5tnu9sIYWYQmP7/cBxKl0lUgtqfe61mPoAo4mMq
7i1Z5gUAwYZ/eOq2TGTTJMa1P4DZgEy7xnOnczzsDLKZ04OBa+4vba9oHvE9w425
Yd0nRumV6JG37whzFnWVvsVSK+6qCl+LtXkiH7EtyAwM8Vm0rWpGjNH6E4wMWh/P
wpumOsbuBqFA558WGDJKYZL0jiLXUvA5MIRAwQqVjfdwxNqxw8mePuHmMQ3ewhKp
WhNO25PpiazK1UsFgaXVzk2Z/rKs771VcFeOf39BiIdzuvJmZan6zxUZzLixxgjc
ab4Dbcobg3HCQhgBPgBIUg2nwBLV+t9I18k6XTkcDF0zjR87Wl2vnDC9VcuPv7zh
UcYRlvGOIbC3Kc+m/ok9hCEDAFdbZn8E+Zwgzt+dFU5Cat0a5kqZuos3bgi2z32x
rR4gacXwgDlQdFPk9o2TMIWxpTTG2VjmI3yneXoshHuE3y4gyAllJmGsaaFrtnTJ
ONnyspbf5Ut7tA+vAu3fKXMj3xYf3/F61UWp5BgeYHdEll+5CEltkHzekVSSiQem
mV1Jo5ki6btEwpGTvwoVjqOUfQ2UgWN7wHQ/04ZFhY3PbaEDQNvFGYeALbjJPqZo
8kd1gXzYZXOU+evCr8G/NM9viyeGQcw1OgujBDiKz04ouqOM4p/tHqSiEUKG+wvE
vwaiR7oYsnIJbcwB9lZJR3O784wnlD2OqlBbyPfB62/g7IGSLpTC6OS+kVqHw2mu
+6MgRFLysRoyjD9hF3JxZ8dGpIwnAHtjgwQTZIQyJHL2hpm1BgUlGqJduDvxXTxD
1n14gpcJy728LYZW0xv8QwPCbgNROU4Byo2jYfHQl21VpBxIzYRMe7upGJodVp1A
wtvYQbNjsV0P0XNZ+l7X5BKd+1wa/zlfuYlqyiqMTWa2bCQxZw7nvPuunIOcLLWm
pvps47v0j5CYnAUaC8OI5pquo43qrSyL2vpCNH/mSHqvgt//mGElAbBmcAEuvEUI
Bfb/o6QNUzkOELxlf29ZnGzXg32uw0jKBz44i12jqokNbpuYCU8tXa7TgRqspMIK
D9SAbkFjKz4lKxS35E3moEkCXZS40U2y+/35a2D+98V1JTe2vPH2CfxGRrZ2sRLi
j2RbUYclrQY156b3yylK+yrSz8VpyPO4JXXGxECIXgUNfdwT/oU7cVLrCbOet2g8
1ZQEdFAwFptPCw/WxxFy72yAVvmLVNpqXfsk35qAJE9GzL1wGG8ov9qGtX4UjKxl
4w7gFzauXlGPQLYESqgz3vMxYiryuLW3HGY/pVgWgqCn79BIUWMkD/hcEotQ3xl/
aRn9rpksWRpF9cpy2f4spIUeJCgUbPssL8dqpS5oZoX4TG319bV1hzckwzq3m5sV
iUBGejzozuO9LRb5JUdGDOul9GaZWvrEtC3Hu81+1DoFwb3LJrLC4G/lsGrTFD00
4ReIY+QMZ1PlPVqPmqRU0WIzA810Sw4M8WHxMQLAxCt1HM+QzUqTQB+YOZ4YL8Bt
Ri525qk4RzDbZZCam+xgU6p36W8XXicP1OFmsI4XdkMYEMhZj6Yk+mtoo/RGtSw9
PtjrNmRQNjonro3BiUrH8rU9/EbXo+qzAKC8U49uPtD99Zj50dA73jObj1O2hqjq
utOLhFpJ2zJPnKVgOhJ4OdtUXhzoCNq3E+a9iA01xneqZe1TlLmbP7cx5Z1ldIXL
yBY8gMDYRYWxjhdHR6e/TToaFNO8d5R6RmlZ/1GjGmEDw43ujdlPKMPXJi60IiNA
hugnpRmVOBlydEsvLtckzZiC05GC/2HJ5XYCWBrGTfsMfKJJsTdiMoGgPUb/ohLe
GyUKGbjHFmE9U39K/fsCwbYa8g/7OdskyZ+2rreM8rU0JFYFegHjuAvbZ5hj4RqB
dyqvlLVTl8V8ziOnYZxhyIk+G/6I/LxYUOmsPKOSV0OmyUD0EoJ2ZDXUWCuggFAE
l4wT2Nng85UZHGcWhiPDV6xX6YTmiYZ4r+LhJb+xzvBB8ZUnQi7QkScOjo24x9M1
DAR6vmKYzJTYSof8ZgVrgTxVkwiakxufLAx9M1BZb0usWyyd8TBJ3u9J8gnAsW3P
VfJat2miKhw5M2F0JTjqRcQGtVblTL4WLcpPwT8uUO5+YPmkfj4GWMTYfHiZ+7LG
D16mOSVFVaKgP4Pv15f0lvAJEU+WenG8Z2i2NO77mdvDXjOjvn5zf8huYQV+uJr0
pd8rjtVeCuCIqb61K3cRjA0RKsFjPoVq2wZSupRacHYhQbfM/g+4VO5eFa2zYIzL
lZ+wcGRwUS+/Uzz2p0816w4xvvi9b+rXbf4w8r1/IsIeCYw4uIQd7ZZyPDR0aa/x
frrlQd3ukm0tLysppNbxFkrOq2Lb8C6pT66LUnhCHviJd0Rg1+ZdoitlXPjtFUe/
nvcOW9GeBlb8SMAmLol6m4T21Za5a5TY+02z+nmWD+Au2EG1IG6N7/tmGOe7CLlu
XzPHs1EBQm1fgZPrMP7AHXrFA7lyElNaHmE8UvcHiklQPEPHMEuBrTPahFh6rZsu
7XVfL/gll932lwoBP/lJNsuWkx2L/5y1mLBDiipdXvMYHplZtKNrVgdPBTPHihVI
kh1HNnCTlinUquCNqi8AZSWSzft9ltHo0/WwjIVLWhO2+TVuL/RX9c7msH9TyJuy
mnPhQ7noD5kBywIvzuS30r3Zy3ZevgxhTfKwA3UHJxNcBdun7OEeeklnmlvF5cWE
slZHGR9rU0JsBsLnn4pwbT2KUNs2sLnsXlU5UWRN/oPocPRRuIy9r/qEVF82C1t7
/5OG7B85Ig/sE/jG0fTr6fPx+6q6eCRgWmElRwIzKGzvs3iZvVnsAL8Klsg0oxyE
SEI92QhBv8kWkEu6hXeLzTKXUxIVbRUgrvjs8EPvhbrOW/p1y60ATEYh5zgjr7Cl
vTbKlljBoMDnaDWeXF4fSAcN5KYVbugDoRd76zfCqYWVMBDtHZt1almzGKZqcLit
kWOmeMbEH6t19J8D5Jx191lPBSeFKg+wxdZESta5+uPqzH6Cavw7NAgqrv6AElgd
YUhNpCzNZcv+Ts+ftWGZgT5SSha++BTbR1r+jK/ueQa1QZlgKrqIIhBvMxu0tBcO
hjLg32+EGy13BYPeHsUsahcM5drp+stuyFGUS2AVm1IN0XQ22u1zxKYLkUyG/VRA
lUR6JT97Pzzc9rFzATQ6F6AghqvQ5pEGr82JMPXiatQHi3CqkOhgIKg/WvI75NBn
y17X8yhaRqEM4lR7YLeuIGh2Ml+Sf+ZsA/NF11xqcXqv9G9MIGT3cfAHnC+3I3vV
PK6o0cciwfteMF5U5fVSKRUs9lwVghrwlsuac7NLVj1m6w2166EqYvTD/aGdADJZ
WWFNg1vBbkkiXxaPbIULaQlC9dtIn440c3K9Cnl+vbEVsWUMGQrK0o+UQkCseSvI
8N+8IfJxWLzhSbbPBjwmyfr1TOKIOX16IorFshTLI9qInPMARpclJdUYrD4KVLtS
/r1c6GxlGia3NRO7jo6jOKT8Bvy+n/o9askHF+cBqqREWLE0EmAmH6qdiUsi36gE
uVB3dK6N5wPMHK25gY46bi4KnaK4szM4OidIGB7EHkyCUZj5KNnt1Cevl0P5vh0P
1EOWI819Bo1jBt2/LIQBlrs+VG5V61rH7KQhXrMtr1sRA1GBP6ZeV2qIaD8JiWjL
VP6Anh+K3e9KisceuF8/gBUOSp+3cqsX/0SRYtMvNn/MKcUejyzMAG12fBnJZHHY
pIVE7yBJFnBjDCgqI2OvjbBPDNUGVeq4WVlWm7Jj+MBmpBz5ZoMJaqYcxL11Uz3X
sQn1s1Tn9X742QLV68fWTAP18RQtunv3AJGzxiCqcBoCto2cNPS0Hi8u1kVGFsBL
wUwh0uKcPXQOAvkIVJoAFVTI3CBIP5Gay3yy51tNRvfG6uoNrFSLwy2T+ZRYrSlA
1tA6ruvXqN4xErEvzcK9b8ciyCPstHOvgEpkKs8iAB18q/B1A7Wv3Nm+vERfRzFg
Ue1784cl3GKu8okDsGmL6+b2wthrO1NuZZN/FQoMxBNj3UGAdKXlRQN8XhISu7gu
rmuNdGPt0ZSjxN1LeqRmer3/bdLTp4SyeYff4wWz3PPpZ8pMHI4/EVqRMnnL8G8c
ccO8E+beYwJTQriwwDLPU8HOGc/3XzUuwuh5FpSfFICegOUI+EYsnvBLlPLDfM8U
aKH7xjcGyxPfHXXMG3Y/BMwbVao+kpqJqZaQ7SYMofRrB8MD2GnVdUYN9VZx46fh
vbD6vIpdTRtep+djq9Wp73BPz576LLuVTJ/PmYUUZX4eVoad6DIe+yXxCQLlQcZx
g7LMucwRJK2fafYebgxgfOZv/+8l26HOhhydg0RJPCvXu6gtcCMViiYmkkBd+uC4
/39xSzn77fC2LakYiIVIODQ81SoU3Nrkc9b5F01pYfpGp2vOdrcvVv/228UfvzfM
TN38Xe9xIx5O95RHSw2sk2iEKldSkvxI9boh49GltZXd1y5GW6sDu5SYK395MsNO
NQJaA9IswmKEuhhfMDkMM+ujws6eHsgnLIaEVVB1WVJrXRkVMP5Ute/m5g9rs1Xv
onUcotXhk2WpnFLeflz57f0AgTXh113JYRzvQ2AnfLiAPxXf21/qcuHgmPL7bTPL
ZT3UMC1jZOxGXszL+ujQCY4jFJvxCo5dX13UdPL/ySIaZGclIktDoE+db5P0BAnX
fUJtLozraHpHh3xlsgg4ARkD/BRLVdSEEDPdaKTCKQXVXkquNTJOOZ+98DXqdLZ3
ZxMSKFTHEDv+9VbaewWwiZ15ww1w0zPS+A2aAZNRGG1jLSOAb2ib5zTSK2Zjm/Or
qe19x6bgQbygce/B/2n1RyJ8BLcUv37TOZxGZe4O900/BAPbWvK+Dq3zXC7wdsKh
NLq2pKtB2Dm2bXElWwA/XzR2eq95eLs4WrskROgkg4ykOMjc/lZJueVkHiktTbgX
TcnYkQl6UWIyknTp0K/ZRD9knJ6MpSLV/vFtdAC+ivHz1VF2qZY7jtSsdzYUMytG
HD2SwS+gL9GZtiuJDSyfogvJg/NH9c8/XijP6ylu2TYJTYAuIy3uPLc2ABlQg8ti
SjQI4HXifY44s2IHRoNZBYIMjQc0rKxYa/aNAcg3TeHML7+o33E8QNaE+UIQXNO2
3JcnWRfhSN/yMDNqKu4JBL+6lXa+AOUpaPOhzdhZstWzIIQJER3/1UVuvVyfVWmD
FFaZOonu89T5hyb+89SbAHQ7GVomcJO/X0J1MDpXFNQxtNECe7qrTk7IrfrfPfBZ
tr7uGL7hHGUBNY1LVuZDv2NjNSABMd/vkIOHVpP6cq7R8EG4Oao+agsHBbP7feLd
Q/8EqbLe3KZoS6e0Rinfyk4YQMzMZ6CoPplndPdkcwh/MVOnvPSpypGyXdc7Mxvp
yZHc4aHsjX6jx5jBa47rswJo7ae5/jJyi99+ydmhcwCS09Fz9tiz6SwMYtF8hujz
1vlety88Pj5kGYAFSfYYw0Ah2euPaAYqx4MeZW+7hhoSdHIydlPcUaKUZE6nwB4F
e5T1Q6YrdAlQ/fqWzVAGMHmquqCw/W5cNyGa6J3ouoQHO+x1uhjWlqlE4zeka3L0
AVGDDkZ+bgEX1f9eVGNl6PfjfaV4xnK5tugTPcs+94iDkkLFYFQm85Uj7ZkyKg6+
uJPQHqw/PUpEYDCXdxZaF59UWpYypab1aY7yy7MUdF4WiPiGcgdJqJId33wV3SK4
SfRb5jSL/btID1y2mYPQV1aliHEKha6S6ErghJe5VRqSls5Fg6rNONLQsqFIf8pC
raQDNf7WUyv9Ltmx+nBIyJIIBWyeuJYfDFjyjZ82NIeIikSAPa/kIY9QZrkWwPjn
f33PHXh0cOK6dlIEo6ZmjeBa5hez4mQJcIgjcHS3yVb3hkelWBqxz79rtIzDV4U6
ECRMo9ItCTyJ/SFJ4u3IycHM/H6cm+pupqwfqOaSSwRG6BJcemQtLH/0QV+y4EIq
xd4FsHS7iLcFwcOGmXXIKZAFFo4VFKvqOHoFCA5M18WoL5HApulOqyPwowpzb2zD
5PmckVblsdNDfMevkoiYKDOy7o5uPfCgSmWgQnQ0icKWNFbm9Zk37F0mbVjfOeF/
jZvsw2XoyyQRDrS3VMDrAQMAJeftoMgCeZJ6RN0COcHlBFcPUc47S8B0ye6JjMZt
D+Fa1nf8AtdzxwF095broyZcCwfESGSVbsFIvXqAOnwwcq6JUkZ+nS08l2H3OZvW
cMGTRilJIS5emNkTeG2DvhYbpfAvXmSR9kjYtz0TevHdG1x2XVrWmgnms8TbyYh/
dQHNazoIxhITLfMd2LlnVap8xZES27Ip/5ykIcZirXj6gZzhcCgIAZj7LzHa48w6
kR/tCjJBprIWDC1tuKg9dZyWYvSVea6Vtl7e2/0nxt+C6AB5B3Yns9aLjVUs43+l
r1XEon14dkFt7CPpyuKo724vXQORsw6+Gh0BwrTdISaML8z+qZx3n0Ff8k/pMbPo
2BrJeUU+2g4pHaAnDErAO4OIu6CUQguY7hdI8fEIRCMJal+9uHWC3E/nq8+fs9TV
SuwhUwkKlRniLn+fNL7G0753bEbJwIlOyGK1v0R0BIszTLrHurG6lY+FgM5xs/LD
DzASkop/hrZGEHV+SofMcBx1Li43nb9ZkTWjJnJ2YKpw5xtFL6pjc7CQxBor+83B
b6aOgayKvE2vBzmyUW6IziXdYP3lsMDc2exLrqG+1M39xRrBr255KvKf1Z76KaNO
PdRglU0fJy719slO8lr4JmAEU2u1toVPAhnr59j//yleVb/7Lvwaxbl0etW94xIK
KzIus0/6tOWJ7QqewIh4J/jeXYYvPA80zT5Cp/sDGyeRnQZN/buexPqbOjngsLxJ
w/vVAeY7b7djnbfVGA1q8NP0mTO4yU7IyGi2Sw/2Q2I2JkadFUg++2KNV1Uc2M+b
w5ARc5ivhTBlnfZ9oJLQ36kVDoRsIyv0p1PvKY6DjumN43HaKiIEfj8YXG4f4B2s
zLUMrbXznVmJiHgC8wKhXlkOMrkH+tMZfdNal/OVfXfAEZ8D8yoyv7Ib2Y8ObrwZ
GRhZauEeSAKcvwILx+qxJQ5XvJnWW5n6OMBDMolShm7wER6Wi7OpzoKVUivPjJCZ
UWdW7t2TqniKptANkh2eoVUfL574fQP3Jfcb7o+wFguKpfnlbFLG3OiddVN2RRjX
Us5Xue1c6xb3ySZp20+F6TwdKGo5iNPLQt7KyhMhjWTIEje2aaNzI4xJbivbOgPs
XY+Tlp08UGxWKyXt3owxochyZUhcP5vd2fUuGgLiUwSFmFGgTt5V8sO2saBlLpoo
FFF8EtuJDhsTyK/yDZ9+sS7xpdE1dLxfJUF+L3ymQk2TXZdoqiY/kG2AeeF4vWaI
O4Awq0z9Txfx0w33sotr73er6CdJhSuXdaoVz5ntVgsSSQyzjv1LEdIzxHWIgzjy
7KC21vVW28qOJOrNQhXJczPlIrLJzPSW5Sm87+xEZu3+SgrIUKaFvyi8eg+FUbdL
4ah202swyajI1m6RVZvy27dfomfWCJVb/MB45yRRLbY2juVTLYgCUGrkAlaOpCTO
/06O3RBhx5htSf8q+eflA3+nMqv0mw/cQKb6nYuQLE8MFbQENQZawdbF7nqk69l6
dCUJH5IHg5vlDIzoYPeqEzpiYJOcv8vFzMMwp3ArdJa6IfXfdbwmaG8Jx70L3AMm
1CazAN7lFAs23StIMruAZ+SfC1LHt6aEfwPK32Wu7ikHEMRq6EdrbkhRc7YXbWX8
30ln5b7Btc9yoJzAwkUOPWvR9yV7Qo6dA2lv25etNlJ5cu4+ZYaOWgJK/iMnPXhW
Wa1IvCZb7G/gVb9r3BfVvbC8vSIaRPi1uGI4JOOvfkayyv7zvfIR9aIgLBev67XL
0PkgeUe0oe33P+Qco8pg0jRCLJgWaA97Janwa9Ru4lG/bhEeTSGtKGMI5jZ9UERN
F+O8yc6HWyNoX9uc6lqnHmjHqUgyHV1WCsgMbKzkT6j3N+MJPFKl3fCvuI8Z9f3M
Ich2GXHyLsPMes0+/xPVnV/fz8JDD/NqXWYKA08l99/lHGa+sJ7fumktGjNzRG5S
LcinTI9bafC+ma3RGtTSAmiZ7pLbD/WLUClVwB+1DqoFDBmCeGGJW1NIjt3oKmxH
gr2OYEgr6QF+AAf98hlE85Ng7e8kzJTvcu2c73LFpj84DdqEHCmqU0/GMfXIolbO
kf3J6FT9nPtIiD+9Ov+Ha+vfo7F0HgPdIva7Tqao6Edci1vdKQ8PJlEQydZttYAo
pmoI3snfwI7piqhH10A0f0V257jflN7mmLwc6+V9g8m8MlMvY4NyBppmmXvJSQ8Y
bpsWgob0K/hjkwK6Nxw7f+F7jVU99cT/jRqKrmIDqCBJi3R+h/9ngOG26ss4ThwF
nedGwYl+jJqsGNzqIjcbUrr5iVtvmWULkfsftmKL6moNKx9HRaYW9mSjlJkJ6D88
n+S+XlPtqw8GDRRwdiOtDlNvm1m5yxfZRalG3M1+br869kyRhunV41+S/l0wgj8c
1bl40eW1V1PSs7Jco8ty1wAnArltjEJrc9dYvtzErc6KUkJCadnF2AIqPZ2ESFp5
qqFK+VXOpwUXsclt2rep/TpLL5HCMH2B2Wi8s6caiSSCNmn8kZrPNbvm+SO0TE0C
bGmsXE45KCQe+ivLtYHIabN5cVt89b7Qsh/SJR6jJhURhOKCIaRQR2cyBiS3AUbu
QOJ+Vn4SXQl6LOaE8irAlw4+yEXhV4IekWN+bGRxafkvi4unDRzzV5uu2ngfTkT8
V6LQlpFp3SzMvZedqVjnPYacjSAwkQSAXSJ9CEZEFfiQpaTEB27PCpqDChccmF+v
JUSpLZCz3j4h/p/fGrHBgzRj/QPw3IP7oThS3tT4O83IFyVTbWkH5K1x3trxL4G7
+ex5UUqn2Dxl7KQX/m34fCGBZJ0vh+ab71U0rhTyO1CyeGsYwkGm9XL6X0b5N39t
qFdnonn9Za97i+05Upyqm8c9OTpyhe8H7islGzdDYFAZNFYVb/fBS1V+ZWWATEIS
e1eAcHpwKrsWa48OFUupPl7Re+Vx4klHRK6wSqn6IPERIFd4PIdqtjFl0BoXatir
qrBqzukYiYUPjrTywuTAgQb9p8XLYAXoAKL24KrWIe+hNQfr4JLmmysZPhkOSynX
0ngRqL83liKUFaWnOgzNOCtZy3K+KX1A1Dxt/gwmzrRBEKL2DGGOAqfEYhcEUnpm
euwnrRIpePjxFVrL4TPzAILJ82uGVshU8W+/hpyR0qq3gay4UEO0k0u+HY+VSclm
9aUwrHsPhn7+2YrUlx0gXeHgJN9HLZPIWZWmLAoL4golrqAm0wTEtCEfcSoHlMwp
0hoH2qoz+OD6eLhpODnZZA4ZAdyHkDgFKq859TFtwpx1GAvgGFZmUWysNZgXeuDc
SYIysT9or+t2x4gImjRZb4bzvIBbHodWmoKaU94wGSE3kTX/7znlrE+i4MvBBpCQ
LjFQnv2bLTR1dPl83kZuuw7TAE9BwuEV6e/Ln7d7O2LmU5aoIKH4BALNABH79WG8
ZdWY4Ucw8hQ8j53JF95zX2YP2DR+J4nSb4+CmT4R6BhHVIb3QtIUievXjImD1twe
u2oxte7vqq4W8GNyYIc/ZvPc2IIR464zpTedotyo/xXHcu/vREJNMw8AFuOc8R35
P+1O/tCMA/zXja7PXskXnVzcLk53xVfEKFHJhirZ2+Kl+Tr2z+M+ctkC2Kj7gUTc
tPcrMH52Ijo/3cIvqdMweQrIjcg1sjygPrZW8i/Y7gbw3fG/ngYI+mlzMzVEOpzm
liO3DiuuEhHWsfb7vMHv0tINF5R/FodvDXyJqfQb8t6L0ldl3ZI/C5PIjopeivyy
jAf4S7NY2Q6ya1lgsZXeo1l1Pjbmm8yEskOM/wP1Viha4MmucXrms1gCb3nhnNKD
vicL5CqsUa35O9NPKMENbUE2Y9lT4KSm/haP1Pzrwwu4cLptBrU+WpMSNL3a3NKB
/APChALR9nI+JHgCtRrM2Ta4x6kxJwqYWaQFPhFkd4STsrtj5C0B9I/kSaeagzqc
QgyXOqpN1R1L6Pz6DAPRnD8D06TjtRvbiKYx2XtTC+l6mtf3+hywgt26EjzXfx7U
EF8scSc5cNyvH8lP57z3L7upJWj6dlxtN+FBJDnPehwLWnYm3HIRy85WfPMkHbkV
WHAVQbA0c6Ok5YUBiv7Tgd44ZM+f+WswKNlC9d5lApZz5qVwUIpl5owUFoeMxXnO
KdSz3j0uAO8ZVep0sRW0suzMwZtC69iB/jK3LK3BrXFyHyIwp6B3pLaM6lyMkHHo
5VB/ngqhPUbGgfxVHrdmkp0jU0zamEUAs1qrZwSlPStdCN+CmwN5eUGdH7PTplzW
SPde7Q6auSyLGlhbzxy+9OwUKqTdyIJB9rii/y28/2j32M+0wGFA9/RMkUo2gUSo
AwdMA12nScKdIc566vumLJ1Up73iaAXBM3oW328rBSD/x0KyMsD9SlR96dloN2bI
aRUWV6hZStq63pQS2svzoRcyG9x7tGCqoI6P1EsC3aayNUBQgrLApW4A2PZH2qNn
1vPh5FHXbTv9TJwKcLo3qmep+KfstSzcJqK8gDbfT8323IP0mNErSdg1nxkNG7q/
SjUSceQjTQO0L90VPEzI+a2GYA0BThj80YyWDyZasrlTRQJeGfqr8OBfWkfx5Ztm
3paVlxWWrpcU42gC7VttZqYfDHEwFmKBvpd9kc6AKRorF6Lg6ljhNDIDUzBLZ/5y
H5TPCIro9lsiMpvSh7JikZiTP1GpsEwX0M4u5d8K2G8E0hi5LAt6dApU2CGx4Z1j
k5OtgOx9JbUik+TUXdZHSoUwckBeXXHlH3hopok4yo2dHYz9zg0PBUjG2bCDZbOn
39GokRQdRK1pfhFvi49aCVOGkmqm1DqZNZPhduT3i1vqD+kJkvHokcSclJ4DuCm2
xIY39WOqZDuqqj8sAP4rDgFfJ86E1CVMIzoA1gMUQc6BGUjNShdgnuftJ8jNfxq2
7+gefoEXPd4H2KahC1G5WQcwHsxbGCK5MGWlkNQjmiDRMc+u5a7ZAeUXopnSLx/T
zgVLhd7kWNa1um8QGfzkdtwD6MJgH+Th3me1MoIeCZz5ijzZroX2SGTozddsH/bG
OvV803zkOOsQ50AcGqy0zv8VZF/vsZAoXpydxz+pQf/cpu5c0iVoOipgi50NeHbg
I5hunfhSfaeVtcKZ2ieEDf3qAvu9rumy+HoR7XvifRpm7CMHrL1CYEFHUB+tio4D
CCeeCq3Uipskc4dBCpUWDzfswuDvDcpD7wp+Um4L1V1zM1uMsKNydqPjeDmmvLXL
C7mtrXCH5XXLpUERco5YPDRL+wextUQEmcgs1EdVM3AXAcyTHOjtV1i58J5zqxem
nNJr2GkFY7fG1+bH10fyoVBGjuJ4lrtzYAwPJr2G1e1IZ9PujM7lX1AjLC4P9Bh4
RR3HX36Nzi8ksHAE3Pikyfr4Onx9sUDGkqeKWuG5jnH37DAhuMGGR1QXWzEj3gCY
4TIK77qMPF6gsFiJBjSYtRhwqsKQOEVZcf1xEyji3xV8zWDdsm+W9UHJa32HRTXQ
x8MK0Bf5goGsV5E61PCRa7qgDeYZRvXphdbM9/eJ+cuQ8nfbWrH8UfXseWaDccKv
xBcX6To+i7cYpJsfPJsqfxFqlaWA1HVfAJd4OGmHSPq4gi//gKuaKm1tJKAMDeWo
Po+69vceuHqX0mEsIU8YGwl84I7bKK6/eKh5ToHmXIXNwddF9huGeazegWtnsQeJ
kZHw2Iddpq5Ub818u9Ec9VYHFMVNynUgFymf3OqTIvtaFTansQpMVVyfqqM337t6
D6dBznFg3+d+SLoGqrZmhQazCp0+2IJfjw5ufuQKHC0XCw0XDK1YyYbXD/2zNifA
ZLZ3AVGnYYp6igsjzmr1oDb6EP3XwSiBgOMGyA5SGx9qQVJXFxO7wtD7pQIhCD58
AS6RCLs4Bi66jVGXKS6oUPedt/5otslfIgjsYsXaUcfkyvCdKNYu2GHswa0ixJKU
1hZTNL6RsNQGV734BC+RPs4z6Of9nYywwI9K7TlmVH/tU9fRW9CJdZ1S3wgGKETK
Akrrpbl8iE4GFmvUD/JDu2OunRkgA0ODl5Ue0WCk0qTBnCUq/WI0OlvsY4jijFse
olH15QucMOHq5FC349PnAxUPl/LUFdj9RPkAyCOQQEMHHQYFTOG8QIuZUUVxRm9P
N1A4Nhfg1H6V6A3JmC7D3AB1Gxoe5gSUEcCPbhzo+J+Rw0vpw1Abf6vIw2TZaSSK
OELT8+2S0V7oHT+BFnpRvMK6KDdkpgeYWwD7QH2I2uQWY9YxbMM3iyqgNHmcr4S0
YPbhBRUKpkoCjimbJnDv6Ks8siDSi9pSYJKVktAS31xfhk6dwFCPnhXLOYiWyydF
oue//A7YQzvyUC+8jlOxpc44sNcl0OokUOVXtnZVqi7ZEcp4CpzuqYtwOBqKK2nR
PiwGLIl0zBFoDB0lK0RgLQmrhLHB5s0XybBaHf2q0+K4Y2OuiNa0+E3jOAdrkbqL
XKd/enxhqU9fb875iI62acfREQEfuTyyVupR2Tg59VE0zeZad5ZHccgQs7axFUVR
gsOrJ1Yc42nZrjRIb1kITWWm2+I+4bnW3gE1Iasxx/1LExDZvh7lzXh2usZhZEgB
afO9JdRTTEny0/x83Bj090QGBqvVO7lS6ue2CyqVVakVk4tOYZKEE1yYHiaJ9z8t
c8IcBZkEWezH9vFtuwIh/nZAbzfWJAmNNWi2c88+vUo+XbPkwMc0bT4jW1C0tAmY
oHzStnvoHk/6JueodfRtJx/dZRWiJdg3adiujI6iE0BWHjPHrzgybVXQvmnmZ9Te
Lp1bIzMWjczm6rljCrOYJIN1v8aWEMRngRaJM856T34/YBL4U0eFtNM7xw7mG/3I
/GxY4qXR3+quT/nfO4y50jpxZusMeN+xwSGLdUyqXD3F5UHTZf7XJHOGXMRkjftW
ZQRtrrB9vx4bdRm+rWCkVHGBuDp/zGn/K5ayC0/N40fIB2ifnC7UQfDyX2KeJYNS
RHs/TvIXDdvmH3oWl+cLR3Y0EfxdiSVrM8A634z9dbLUNzoQcboyeTwk6mzk8/Gt
yj7SiVRv2g2XM9Fqbo14jGJZUesaiJTF4u/p24EmzlOu971PZUFpcK/l9aFmKFdH
+rwDKEGsLk/+YRwIb8x7MIjPjvqrbdt3tUzhB4JDgG0qmSIK5IoqygvaffSTBSma
2wXj/W3cD2V484s5oC+rG66io6YKkEvIy7D1x4/bjAMRfa4VD2wAulzC1TnjDzL+
zcGTDQ3QyIabKYpmocKBSO6I9s3i4mSkYwWJiJtBdLtcabWWPC+xhHXLlSOXVe1J
vg7nuS3DCcFqxVluv+vwTsUgwuOLLEUaNK6e6TA8xBKng2Tp1/9BA//63bsIZ2sn
HXu0iXsfJqXZn8hFRjFXlixtQiddFOnHJoP+6b8UHAxhwBNHjzOi1SdYw0lKOPWz
94o29sLG89r2mKodcbX2cTUiGwsTICUb2HYuLS95wPBcG3m3F6E/2ZdFe9SFCBTo
9ZCsg9Uob40BVsDicCXxEdg0FQA6tRr0bD7GvrSWrnpxYY3Zlf0IQrgs+rFuE8FJ
GGuVzaYrURgc+QX8re6J375VXp4GmE3ALz49OohF9Cj2TTS8g9izxVs5MrdPLL48
eJ870rx/Qs8OaiIMY1bpowYAbisDhgdbelpJBfB1CRwLNP3tcHF2c7I0MDfofySK
zma3Oo7YnFY2ChVA4e23g/wRyS6F0d58BXadCQ+dhKCNBi4T+4NUTjERxBrlfNJS
xdvfl8AxsBWHeSWBcJak4D36SmqlZidpzuxqjMCNBY1KrrQm/+Gh9A3NSuhjo3Su
gMH1ICGGxsK7KdIjij6ylTHBCfm4Zr4iCR6hZM0SSYQin0ac2EhsSlkQ1B0Wpq+3
OlMVrboVL1PLh3DSdo/F5w+pIhlJW4AfTaRe8ZX5MjV3yN+7gixsFwbTayJWBTaE
0wJH2lMYEfJV7poR6Nu1+4wQqIBNBIV65kf3fjifDQar58f0KbP2mjOQos3oLrwk
eUMbzZJv9oZC//XSSlsQIGwHTPhCpU1drTS1AijK+D0BT0zpPqZaGSWDUzrGjHs7
frYpaNp96vw9v1Wik6ek07Whdbg/ZUIYLpIn6Yntdtxjmn4YA53yxEN/LTHA+ECz
CCQeiWLSM5LUWH+aiTaunSKiSm1CC/mE92xtu5DZudORzH/cm7++koe8gifI0sI3
V8kX53lvngq+gPSmI89e5XKWhx1sjNwJvcdRwrfWaoz7JuhqqvZl3B1OoB4+d1pt
7f6eVzBf7KG+LehZNkSKf/FXET/rEZES8FnlZRUDavia2GI6hE9B4m4ys5/VIBZZ
YcNYcVWym1J9uVt5Nzivp2bQwVprKgAATahWzJD5pVz1BfudOPYsESjNfqszkAWz
rJzX7piFpyeLWhkcXoCyu57DkwfS+/CRQQo5LHaDbwZ6/SGC/XD9xGrKBTB1Gal5
6Rqe6FhYhtbtuuv8BprVSttPedfa4VytlGVcJ/jqg9BCxnw11xWvb+8fdEoGZiA5
xJzWwhewSsIUsQVbtOgSf2ctfKrBh7wB9R55eyXXlpud0LY82djXlq6jgadSJQxp
Hs7CaSfNmwpcRxkIxO1dTvVDTOgcDjVXTKdXwJKmWQD0pDPI6iogiY+7N7vTgALd
94DCtbkJ3ZVjJChDiNU1xlrRPIo+W8XZNKfPLU3nl8+9VIL54MPQblE5DgDJyfV4
wscscbiTaUx4o3d+A1A83cA+rTOKBaJFJo2GTkmPdzFGpIrRKU8pyvIYVasL7WvX
udUSFU0JD5A5BPuKFrIEq8YtHdMLMix1AAlsHBCylzEP6d0ZaNNpVpE7AalZEX7a
GEXSLrtMFnC3o3Va7y2PELb3IP4jdW5ZLHma/LOJKAwKYdgbFC5DXnXMUmPLRv2+
hdAVsF6ozpBBjG7GArLGcS7GI+QHzax1yDLLw69GEpfYVDdefDR3xud2iKNMX3pZ
snFJ7P2r3PbSJrH+dp0mcckb0Vcf29B+Wv42Tqbz8zGEYzmxL/jVdQJMJ3+XG7+t
3PrY6S6tkIZihzdvwhN9PklR7V33zKULcUNCaL/BcN3bZg3omo7aRwizc8vWd0Rl
+qSmKaCWlOaeOcSYalNwf7G7581peJoqFPmD9bBkdUCd2yQSavc4SFDC7LMzxSTR
6JHtkRPxSnc1GBsc7aMhadN1SPZAKrwyPghV0S5p0kK0ZCcpdqmhqSDzHzOI7Dnw
wQI/u60mCYBmCMQfjEtA0ZV637k6kr5jxW9mDjR+eJOjDrRUvlD9G+E3DiOadYHK
+GCAqWHmkhQrNmtBB0hPIbjal+4XDl7mymTlFSX3zbQk0tIGnxBFxK2B3fhtgODs
FxBK14PD4l+tAsXMgp/ZiTwg8yls4SfQprqJS2pXZWADIx1T9iEr+59uGVPlZb5n
w1Hs/ehpawA1aBESN+iLNMi8bRTdA4E9Es33d8D0zmHLmnwj0/PqQAIpcxRhYOMH
PZqWxxRiXqL7439gHK+lM8E0HvQLxy/DYQzzNk36maV5x8ZxPRnmE8kl/qWQ7XbL
ks+EFy3ygOmeyf4kdVEoDqsGCWfvrBP0lcN4F1leq3T9mBp0r8H7WTl476Dba9yR
GgxxLqsJKMzOMCjFZ2AgRDAjUgR7jvgvXXj+26TCwgam6wO35x+045oYplJrCtpL
0geg8FWzNGhWTVdmEpJCToZDelJOSPOTYqQa8hdiZ4jd2OnaEgIDGBPWsAMi+XfW
XBbiHSaDSERXeR0WcmBIR3msgR85x5RVeOt9t7n2weY2Ym5abaM35vKfLiEBHYX+
eG8fUKF8p4F9X1luN5y7vpiTX/V2sKI+ndd7+fdA9ye/4ioDkKmrVf4XMbNValS4
2k5IJYJWxsjo1M3fVecudWXdZukW+sMPXQCS/tyoJsxM0q/h1j/mIgaefE7K8CnA
HhApDf24r9JaufrbfJwkMxEHpAAfJY15C7nI/WFTSMfZh6LYSxpUs7ExQV6oiB3Y
OA4grwnpjlTpl4thkKnM44P5TbfUUtzp+XgH7LctWCIBSa5EDDpGafWZ76BLU9T7
FtDkHxBenn2hDjFqEjqk3WDDYzZcnGN9QSo2m0qV65URQufD7NMvc27ZWHjWz9qV
KF0qNr2CgVoQGW8y2gPlCnPGB7m2H2kh9P6IANkzPSizKLkZ1Lya6D1qgLItTLpD
waykxJCaYsqDeNQcNFbOKt3l/UJXmF68JPkMaxHuyboDH8r0fzHIJa3Moe4uvBex
Cnc9btt+mK6gs3FePnATL002QwLyDMuQorTdWL4rAYc9aGi2sGsL0BYKcNWvnQ/R
bn/NbyBp3ml1zQC3R54yEmTUnjLTJ3DCctUAOWb6bgXH5pu3PtP6czMy98apNyVi
7aTXHVdbyeQNvIYvqyNFmw8JOFtl+FiAdsdy17V+gYordgcN7uppWyifg4+YM6/0
poQ0P86XoCIaiyEcEkt078O7qM37XBiVoq6vDHkjTxZM5suGJVVYJv/+ytUMl6xF
YR1uRRWrOmh+DuU3rp2Uj2DHYVxu/bqh2uTYOVq1bl52KZ5eynUTnuyOnGixc7Y6
5zDAmoFynno89lxNsKeFjZQrEaef+PzI3U3K0rc1/GLCXkaqideOpgjJtgWhCGNd
h3O4YyXOOVsuP60U2rbDwpA+J8iULLWK3IO60bJR6qSKTUzmgXOnjOpv/Q0L9kDt
MaqgTsd0HyJouqR6a8klpWsrEKoxwbYeQRc532WkLPnnbMX2QI3ZRDuXTU37zzju
iRCx6V+cN0Tmt5M8X43Xmi5w5uAOEmIGkUzUbqmBL1dm/z6HSYm1wSM7cjEC+2BB
TmE7ZDMUxZyaLPeVwTEPHuydQ+/xyHZuilUEaHTrTYklGsGxVPvj5iLdYS5DAIkX
tUn42OOgfx2+3oN+gakF/CNe9YhzgJ3XhcjsPQkhElPuWm1eg9rhpYCEqzEVr/yI
3ENagA5Wz/a/2Zi2cQEFd8MAmZyM5+/mJcZp/xjRQxCxIjduS+JflL4JvyWapGnh
K7sgKY2dzDa5uy+QlJ7PDw2R8Fsl6Zt46WjrT27CwXcn3FTcgcpy0QP8eE91kAjM
GLbA6yRMZaGeqEpvxNTEZqceOXvg3M8ohb2RHTMsX1fTgu1sDltdBNfVRCfwJqAr
jIaV/UNfmb6zPMrKvilu3/1Ydehr0opWUhlU5bFFx8zqnhDc89fVM20oVXxfbdXy
rjRE+nBD6i4hS5YB6XNisKGcPnbCnCSGPitUb0hwjlWiVIFwuy0Ax4IN5LrHzjuY
iMDp1nd3CE0TFWC6w0nNTa02UPfyq6ESkIcg+HDDY4Bzzj5cwmcV03A6ZmWzTfZb
VBRCUqSdPy8CViU/ItNFaxH8FTJGNnYAAz8wOqTBfqJB9qW7L/VfFCQDWB8tzYv9
QRyvBdzfCLoxSNWf1ixfXFbtkXKVOzOr7bGfETT/Ijok4WBtTRA6N958BadCMPKP
RwU2imkCveEDXlUGLif5E8IGlYTQ1feosdgUUW2JW2tRZ6f3VGCB8BsqstfJJjqn
fBd8fKE6WnFgZEcdIk37ZeFiU7mJegTApOwNczzo8dWwyN4RO70/HncntBQD5GpJ
5Nrr6E8d2IrF1d7CGurKNSraZ5fmGWoCovhggKwCSdawZI0j2BWlqlzucj+VRAUa
NVm/jqFLjGKslhsVOVMCeQt++LF2/+H6EEe94/iTCb52HCMOJE3IQg/c1oBuGQIT
CjFBSvfzbADpbxNF+2HwP/PP4BfLOpVLZg8zbk7lb310uWdCLDy5aZfTpitW8LZ+
BvH47VOpHeIVIDd6q5T3IA+j+uaqtE/fXJ2FujjOE7L9KC9uBgZJndNbyJ/RA0Ih
SXWuPeo7s+vJjxfPohOngLFQ8x8Xk6Wr+G/BBajWQkwHnQehydBqnry1DJhCg4/G
F5d0KKnyVckiypJde9g8RBqUWPZulhyihA6V/lxAv/DDJ8s2uSLylilcB/+X86m9
USwfuXI1DHffGDf9ZKjdrV8idSsp4kvKnPYmcENRyT97eaUEqSPveyx8ewHOl/7Q
6g//ph7XDVmr33i41xbdGK4QNj9xezwcwzi9rSgH4DqEObJqkR/w1UZpNjLOU+UP
pLyPfJy9wzoHhqMYKEVjzDr9/37kyrIahZfB7ekuTWke9FoWh7fiADFU9kWPjBEh
0rXpNUXjnhXOo+xi94hPj2QyB/8ZF/XRNyI3Fkw5rWLXi8PsJYNiJiALDpEPvB09
lOjmFwu+sKWljH/EEk6zFM3Q9QF60rYCTFYTDPdvaademwSl0IbIogv1AhtRlNLC
rOFDmWa8K3Uu0bT0Wl4lVJ65Kbh1RcbARghGl4Mu0jNhwXBUOkkZP56HzKT5A2aK
ZnJzsMftVufEtl+CQL2I1kdhJyaeStLjbz500tdNMEtjkgxLPK3N2w9OreSJAlZh
kDNrzeY9xC2dGqRYUA6Q9buKUSyF00zHU4jXnzLjwk9MCEas24D0RZ2uTeyAkISW
kMPxm2dU0xcV6ppP+etXqSAUxLnVd4xAysoBRfBHls/tHmignHl8946bWdxAH1XX
Urhvznme+4UaiszSoU/2MitAFh4+88pWEMkSGILq155KJrurJ2eGdvL3WIqS+QL7
A/ImeHNThccyzjWXv/eCuJLWZEb9fWUuWjPuqEr4etsONuyq0Rzeg0QhFyCrjB+g
8W4on6heKwHX00bP1fQZTkbGfst9eERWk2jbwU1ruYaRKg5zNp+IiIgQ287D9wei
fWzaYArZEB49X7Iv3A9vyLJyPWNNxYzsIc4C5+BKJj5kYa6ucSpsPF0c7YGkC76J
AXIL/A6w/GfJbGmwSWDfhMc5LTGcsEL+5y9aIFDL7Ll77+UEwGNuLMt53Nzaq6Nu
2BeTYibvvmhIULbFlhijS3Oewcj33yBQxtKK3h2I8kyb5YEVM7q5tYkFh4nusM/D
qnpwXqaqozV5CpKj0Xq0lwV+rt6yvq62XkzxWXkUp9240tH6XFXiIGT3SxOFZK21
KB02L7QgpVCcVVonAOWmViT2w1PuswCVsFabknQekyn/WeTyWjOb+y+3ukMHPJsm
FNSIkubVn7NKZWDd/0/DrIbkqJiilMLhjRU539NnAWueqZsbmeV143/4/IOxAobN
9NDXgopyrX42+4lXWGX+DF/E5UXkH15eWvwtXijssbL329UC6VjF3aUw2FTzH7fH
EbWIFLSWhZ87JC7cP243fSULwSdwrfnruI0fIiZJdEdoNtxX2NMakMFB3eTSEI+T
xKgPGv9c1uYzY/IR1MusZk+erb26q+D8hNiuxRrK68E34Jrs2rTOf2mBI6x4UrML
C5DHefEcpiRUdcj+H6mUdsFjvXuXRTDibGNJ8f57VHrcbjK/E8fw6t6KgCkqfu8X
0jaGIjD/flxwoVIW55J9++ISxgLPQC9PMa0ZMvrhkAteEKpiSQcvOFHU15upw1xV
lKGTwkE+aZDkf25qfVmt/OBJAxcT44oTvXihIrr/qJndtmpHIThS4z+awEHLbUP7
2cpKkYcB+YoQ6xwBuIAV7vD6bEDS+VwbBgFaND3WvTt3LvMF96dI9qZ1HnD4wLEL
dfssOxCKyMrU6L78uURpfXUbOyoDhYEyp5nxdwynpXlAOKzwyxmpyEyTAw0LkM0O
2lzdgM5A+Z4zF34PGHn8SuEdGIt4ZHAOyc+R7pvr7LYaFOjhZAT6v/kGd0QCAM11
MbxBbxjnW8H73+DujNp4RuspuUC3jARk0z4v2BoTY6xbHRZ+DlvIN9GHUYUJ+PG3
JyerFsCm/xO8320MCKYvrYYFMpJ6/fJUuL11JxUV13zDwS8b3J/bgUC4cM5AZAj+
pT4yKgzhZNQtWZzaDGseISVXToeCyvTC6s/R35ks/TGFPRlDEEJaXJex+p+X0o3z
9/5EdSIyPOqo9Wx5Cudzb9yNNWbvey64WJ34wpm0O4irwdMlNDQ09i8bTvvtC3eN
C6GrHacLBvQ1Wm8gKTESFnrfXxSXkUMqaKyoB8hP1R1qy5ddB5LrOTBayk7BsFwD
WMaCW/QG9VGCDtQHUFR3v/2EAZXSjECEqenlFsSNzz8bcHs1Ug990sIEjzKSySwS
KSZxI0zSbofszQiLgXpdCem/l/Za1Ppt8E73j1E+QrH8P2rQguUskM0GxN7fmors
u2Gy0EqpKVgY3w3XF08xBvPdVO/MCYkZTyLkwlKUoidlXu+UiZKgfLroQzIJb2dX
mZYQ2trYzWQCVdz5IPUEOqH9RZKJ73xsWx0QEnv0d2QWgkEqmVOyttRCmHVJaWwF
J5MYKOel7pYTi0JO0FWEAa8OSNYb5w4XAztFVrAfDVymv1zmdpRphvCWnkr1H5nw
rEzrTaFzpzEkuxm9djcAnu4ZmHKyex8S3fHVdNuaM8EbZ6Iskx+sX2+OK5OO8u5M
+d0oDEG4FZxp5xRn4Gw6g1YxNmp6UkVBO7lWmCqQaOW13mKWtyjTC39qOq67WZg5
pebZa1U30JopD963q0djtj+BdXNh9gqbrLqgjZE5DrIg5U976CXD7OAah/zBMPiK
F47k4HLCh5rhScD7WhR/axAj3aiRosFc/LM9uMqZQ4G29QdkyR04+OH6u0PJxr2s
u4wGBLbzeVcLCGXs6Elewva1kjbzxmDex4V/olPFmKEqv6lzH5XC0k3yabbZznP0
xeVvv9y4u8LX0fdHLUEB6AHbh75jROj0cWu7Qnm20pol29HMsXeToR1ABXeJI7Mt
ydiyYFd6ojmYJqOh3pkI+PDFX/f60UdD1XBRTcJJqhaskEcrepCMFlK0Plw29L0y
nkVKe6Wwljbc/DVgA4PrHwaEqAFk0pUpn/dl/IED+Yd1EixqpQH812iJVxAystWx
Yn7134qTdgHjGiEipt0+ZT2KdRIgl2D5m+w8yeqGPggOs6peUPVXp9V0wfQwC/ec
aq68ex9V6TakjfiHxIdAJeaQ4u4LlEsqlUQJGouQ6RCmx21y+xnt6a18JiXKtXDQ
sRIdzJcp/VS9DhRuhwac7GPJHJ4q60/X4+jNFqnKpWpNRskGd1y5typFhjvvcn9U
lxw90KcQSz7o3g87k8FZAs29Qd35H7HojtrnLRSZCQgwwUA9H2f5jushiYwkgVJo
9gcEVXB35LtB1HkXqmaYKZG0eSj2Rj7OFkR0jr8J9LB3TVBMhQifyhXtvGkMNJBY
Eowxhrc7zaPFDPpDOV600J8w+YjjLIwLzaEPftqU7MMcj3MClL10pgk1PU3StXGy
7uKq54Zk85NEV4wkgGX5qIKtum1olp4v9c6u6cSfaveo0FFhY+8A/WL97uItg+pa
/mYGTkmmAJMQ5CkBnZs3Uk/IiAM0k54jKR+WlSXYnrF4Ax1JJi9a7Q8yg+bjcAV0
lUvJCs6Vrx4oo7KfrRjQw5vuCAzVAIVBe5WC0VeKy5Wbu8l0GBioFcSGte5p2AFc
MT//mPIK6ZQUVH6++7HndI/a9fCito1voibJ0ZRCOnLoaUaB5SNArriN91aLRiFa
+3SE7xSdGwOOpaQSEyeWldpNBoRHAR1bKnxtSTV1MYObGzDDnhmz6/bMBDX9Cq2f
SEiF6QgWNS19j6K81cI75XLoUST3YxuYnj/VxDbocktDPrBKS8ED6wFXjxXDisJp
E9WwtvevAWW5IkVtwKaPG/3tR8/Oy2j1jKuZ5Ay0gtr4z6g2qgEq5/uUStMgv6M2
KQ9BLryE5hCPbPEPw91druRw5N1k4vI8QGWVcaMQyhMyWQU/ZxgjGCarplE/u0+h
xsexHQDhgz/95zwH2vHYP4OiRIdmK8bVMfTbVJwePhlbx2K8a3xo3QdFh7XwxYs6
GKO43f/3997HLy7BPgfCVomDlGEnTgi8XoTO8+qfw2vS78Nf4pBgvP8P4bEELYCE
87W260tf3OJoth6hacleSyZ1My1HlItFiIFPmYiZhl4ol4Dlg1cicczqUuiV5Pw8
rWLZk6ld8ymoTwDFw4R7YNwLI36jYcyaCYyREpMmxLHOt7JM7yyvSiz7maIxviEV
hYGhV5ubH1nJoGpPSVYBP/452/hmAacIGjhrTC346dj7BoSIKqPn6Rb4t+ZsFbTt
WP/9T9XLI5qfyKazuUy6cPdh1Zsc9JZkJoGDI6Mjapfy7wRWkFeA+86RzpMfokGW
+dVQSLP1IiVmsoro3xgU1/EOyMy0RS4a83iNyawzEDZFdAxTD2AaFQkMK7pBWNdT
rzHbPQQKximFWibYYakbIWO9RQOnR2v+Got/C+z0ueunPEQZ4I2MCiCGqwOwZvEp
aAiwIQgy2MzHy7FSjhk/mo1HpEKtZSYGZqEot1dAktMOM+vbfUzJbpHHd4ndHX0z
FLNCq5/4sDZ1HsUGObYxTIwW14WsRKGznUYT2fDzBOI4h2PpEgIigBsf0zJnpmi3
5HKZD5j/A2HdeWrJeJyDzexiufXAsMWZA7E/PXeohJlObguoq6YCjGifN6Ebc5r3
7RcU78jWd5BmqDQNnOffk0HIiuhVWtS+ubZ/773YEElbn4od6zu8zf8Axgyyg/YJ
W+PRXBOTnihjK7x9rnNMW+K15DyrF0pEtllUkXwEd6Afig6vPmgUpX2FLRlP2yZL
xqWi75vby6ULfm0efYo83qqlb1dLQxunD+D+LM+EBuAK7HDfqvXREUT4qJcD8Mnb
6SHonoe2LJWuhOBc1plOynlG3p0hSsASq2U8XjjDcyXw7GDa+EyxSIzneCO+KuK7
j4wLO1rW6KIS0n7KE4ymRlGg9GWsMhJ1M9nxW7L2+K4YFNBfzBCa63ISlX23PzJ3
bsVZL0qmkcN5c1sdv9EXfxzSV9A7t80vQQO6AEqkuhLO+KVAMyk6NmF5IrnbU511
ChFOF830WNB1HxSt+KMr3YYkQdKn5m7Qm3xEjNZXFYsgWn0UDVdgrj+MbSLjhMwC
lpf6FjMApeyFSl+V2L+QPFidQERdCA6Spm78dFWPe8dq7BsARrSBv0OfZK62vBcy
CIlT0SZO+sYS7MeasxQUIW5Pz9/UAerRfNaSwlBmISW4eBpM5iWI9n9kMonT6KFy
T0YLd6lU/R2Kbe5PbGKUyJ3pAl6gf89XHsbm2IKW8t7r/F2TOlIZFt8HhmD/XK9r
LPIffh7kh5W8rR0hSYL8n620z9s1iPW6YDsV2Myurw/GSq2zrj1myx9G37Ie7YT/
hJiTErM0huv0iqAVx/b2WdNHeL46qRqRBelFETeUZ6gjKYciM00OgpjPDGqrmEra
pq2AMjtZoPcWos7H1IjhbHCGBYzhX/cdkHC+zzWkAyb6YCIxIBu9b0SKBZsUwiXc
FaHovFMa+bC5LDmdKHFhFQJSsJmsjEKcXUhPT/tiFTypGvlzoVBlHzHe9I6rLVs/
p2PnjpapeLzTmF+w6jzPahaWho6M1laxJwLqjckq9OX0S5L5s/fa+PiHNRshEhWC
TkdMGiTJMbuTSW4JtrT0PI0ojza6Q9V7ieDyPNjXVywUZmgyy3a1M3Pb0HXuDGGi
oh6TpnmxRyKU8mOGMdg3HEkj5bhemZk2ycW2E3tQaeNK9095MWwmM8oOTDA6jPc3
8stcwEzkmvmZjkhT1I4UMkGM1m6/PeIUduO0l4CMp0gRQ343N34GKJ8BrHV7pQE8
W81WWH0vN8B2jVjRjC0gCiU7Hrh/T8r6p+BmcZee8MhKqubdE2HaRXysGsOOhm5j
B0WZd2+nEEdpe8ii2zTbXoYKMZbr7RRbgZHyImvo01okAaRM2vZBdjZTbTQS9Ack
WzP6E2QQvVicVUVfOzBfzQwBb4fpLsievYppOrSp6qHa9yM1yuQ9uOBCHcSymOln
S4nxP3Uz6pgY4hvf8Rd0f3eSxmAX3cVy4TOjQ3Ux01Kc/pTWo2y9U50lo88oYLjL
62LcZQdS6+tdg8clsk2aMmv40+y7UX57/Zw0kQAUvLdsmO7E48f4oOuQDKipSpjv
lnPcK+3lUEVu8njMyEk+2X6OG58dUYbc6dtUF0ANIn5U0QbXEhKhqRGOX+TZTczm
K1KiN5z69eH41nd+vglAWUXAkkiQeRy9pbthEjY0+dpea5NS0CWYCHcSpZiiqJe5
N8uHvYq+pNLTidWDHpKkSws7qj0/4ZLkq79qccOW1oJ1Ygd6a9mQEdRTmMpYbUXT
1wO6ZAgSyp2XEPZktgqdqiiFqtjEL1pCO1tZLku1idt+okfahILvfc9UTEM0YHKQ
G3tzsTfsRMoUn3cCAaNdDZykC482NHdvNvhUO4QdKN3hI5n9PsH8f4hdDpGqK3eK
pfuCNpKVF+93+6fcI+tWFbEkoVXma0ljZVj0udTFzjoHfSb5MSJKJOXvde0XD1ZC
yXIGqSNa6rGI6m9BgUzNYKUzDMZUYD+fdYFSLBebSjeVCEDTrQNCWVQ/kNE2KODW
mUnNgX5NTzkG3wkHt92a5g15oW/g8a921xVLEIv+cBLuLcqWB5ocyyZV2Q4K3U4r
IlD96t1gsa0tSjqtA23cnuzBI9jo3uscwDMqamUO2s4omvYfYe6ozL4hyMbwieXg
yxU5jH4jAV/2z/DH1owmD1zHmsCuX3KGKhpmdSzFZYfFd2x5kKH8PiJhyEdaqDTD
kvx9V3UJDkscoow7MnTkdpF7U8fWrfh4Wp9L0n/qrUnUtzelptVDRGTOQmUyOaoR
DmdJMF4vXGO6YheoCg/EdxVoA7RHF3WGfiRA0bTGhDdzuvnnqZmRXGTgQz+Zgv7L
ebETQcWe3HLE39m8qRYD6WWdsENrUmKIMwp9LTAaedPcIknAbwGqVCxqTJaFaAcj
fz024e75phmHm0v0SeftqjMVVQQULbZNdf9SKzm43YdvG0jhSN/JHzPjZ93EvzDg
+Z/ReTT+mN1gmUE4YQ2AlMK6GgpCbhqzLI+itKXzCMJXbUBWEvnrSpgv9aCmmGzj
YxTBHiGZcMfHDLcaeF5XFi4E4kWWM3Y7SlYbPHkNRMl3TacH8C521u79BKcvwumV
V++5RdPbnL+dsg9ZKkppUDnnZq5hQOW1Yrh6TVqpAqDP3ibmLlIivwylw+G6w31M
ZSWsiJ+J+aLhk/5/4hzxBvU2bDkKsEnJUcFlLUT/IUIg1j23S/Tq76SqFD25/erd
e8k9nrpljCq3S2aL4JR9jwh3D5YlDT7RD7pXypWewvlUI/9XCHpWUgSBb/p1j6Gr
RQo3pNTXps/BRvgjx/cLLWzrx+VK3ghnBDAbkIvpuhgL8ZEzShZ0KK6ClsNTejoN
Pwd9RRR1sBMBsdtH8LegUaBJwIxuM+Q/kuYLvvlmvcirrXG7qH9sNdS1iyhZIfjM
/eYDBxO/lJ9728qrul3vMZgJfsJihYHafTizM4qyZoNr0m+3oMtu1Nosv/LEx0C+
ynbZdpd8X1VGRXlMVWpB/+/g9MjNro/JwO4ZyjX4WJamM3UFgX6w7KJRCJ3jKdcc
VXieVhJnyrr6CklJGIrt03+fPKSubDrIuwrxvsxOlZCq/DRzRvWDtzwjhp24XN1k
ZrxjQeW/wOPyCDppgjfaWCFshGRjznximSd/E+mqAiSOlcrsKpYhscAvnGr3f+ml
egAxDECVSnui3gL9NqMeeyZPPshzKJKwngcqBp9arQoN6P8w/pGRJOq5if2g/V4F
DxVZMdz6PIpiES6Pr9BOkQOvXY9EGkjeCO9K0xSr9lrxH4BDdxe/O1IG2G/ahyUP
MWQRrNullX5QX2yHkpJRZYYAqgugRJS73ZAYDHcXbSRI5bKib4NNwDJHsJqXmRz5
MfQIlx2G6nI7PYO7dbvU//AuNR52sa1ATkVymp7mMvkd8AdMVOoRbYXmm5u19woE
KyYZqbfaMFH6ChVq5t6x3QCUM/CSXEW3CflYFGQ1Y3A7oJEY2mZSv5ChOh2D/J/9
LVKgbsZRJvGRlF6q9AMViHpuGJ47R3GET7cpiKmQ5B7yY8FeWbeD9fBdm5WFVdjK
yeqy9uTFcKx5IFHFBmE8Ro3gCvUj0L3lWyRFMjmROsgngTvairRrwRSKrziybaRG
jZTTbxindnrd+3knmot9b19I3UDa4Eljl0Qb0EL7c0LGICC8BYvNRCaw1r140tDU
tsAgwllFW3SAV/TE7FDSCUbH7plvjJP6lrQwqA0YW342mKsgTDD4iyTER1cwLX+s
9O7ruRYXLQco50dtrdluTyMfImQEgix0euVapSb8tATk19ji6g0tSR54vF8zSaHA
rpMrRDvX5PXtM37LquUuL+2bOOjanPuDEc1gG+szwcy17Xzj8yUEAFJeFCRc+4Xn
MUx+gnsXgzruqMElENm91w2P0AxtQXk1YS+TwtaZvhppDr2RcSwO17H4UmZTUXgW
VKRcJIE7XL2whFKnzXQKtx0iqG8ZXwC2UFHqQgV6XIYpqjxSyDkgPTQujjrASATs
luXb/2rvLZuG1+pGOOZ/c3CONJnlShOMxTsa+yU1tU8liF7kNLEJx8tZ+RzAeoP/
WWOtQBJmU/ftH8rPouceXFFTdu8zlykiZWdZbcbZVlAdB2RHXY3dZ10FFzPXgc2E
rmCE4cKpZuhRHVGdBtesrVrHXJjGYMnsTI+2vM7s6x77XsIDEoN0TNu7aYQrFM9l
VfCHajgPrJcaUJEB1AwIS1MTIcqM9N5Tx6peAXK/ksMMlNqZTe4g3FLK1MPPEwAU
GkLfnG+uih2VI8VNg2RR0amseI2TQSg7ghvdTfLiHVo4iEIftvRXOhnNk5ZvnSY9
MK1QfupSn4Cf3UavYnwQ7YuHNbN0sRJsh/ST8jSJWWaBzV7y3UCsggpNWFhLA+dD
W/UvuQap+tebRrPf+L5EdIWgrUA/ylB3odotWovcdWknHjdBXwuYaGgmRpx5JBu4
+07tzKmeKXt5Y7i8a0iE/Cgu4jdA4ZT+OpBMkAxaVTeMMPj8TI5qXwQGMcVKvhDC
ouAyEgGBE1QX/JxrswmyU2Ex6cHsDbciDPNRB6OghxfBrzrrP4gVRKron/8az9Yz
RqKVzl8nopE+0Dklggap+aQPHFZY2jU2/BlDQTnANM6MnO2PobM/iM7OeLghxCGj
S0ZgR/xITY8rwte939hCTaiS7FrZhJ0wAY5pykdZSDR5VU33suCLFVM2TrXEaWzF
WjVIhZ0Ur43C4316A6IcBzRUrZY+jEGkIF+8vGtI08UQwRhuFNPJDcf8R1ZpNFUl
iKCGUl1YGrLf97a82vsWXO2Ww9s1tEhjngsYD655f2v2+i+n+DfyrjD5RJOQjSC2
2ZFPgemOizTLZhxdFB82RBt11x36wH8RJEfq7od/ipWG/VAhMWkB5sCqaHNBeCAx
JN50V1N8YGXGghpW/x7dH7YItVhXRLFZz+n+w/i3vN5Bwq0b4sf7ThyLJ6qE+2j0
94HZIKXuB/DRDZM7dmj8/6EX127+0Kle4GjuiEkWpTtnjdOe8OQBT8cI4lLJavjt
koRbqQ1WkjqCQYAFRLL2BwLa315O5UFt/AngKyNLTJkIo+dTTA29QFpR4OsFWHGU
XTnZfUz83GSr5Z/kldAsvrB1EhqTro1ONzqqco3447V0bW5d/jtYnIEa1pjxC64e
HvjWqAnFJgz6yqg2fwMY7zP6t0u8iKzeQbaTxWhhkT63IygUvlTinourMF9DTMjb
dhmyE6OluVGS+BA8jUbCmpfH4d7IPhRsK7q/ldXRK0+ouRU0EDIr75rSwUzu5s31
qjpOmPi5SaypP3iMzqaSfZ+EmU3N7l2ALL0snFDwa630nu2nwHzXmTmZTEgwb10u
O4hzklF42mJ6iBreTC58Ml9K6598pDFQkqRugRVfhQ74kAupodhQu+xfo2oJB5R2
yqfCOY3GIWoUlvH/h3xOElexC0Ej4ieRcPzohzwCEiBYbHjN8cHYCJNp5EG6TVOY
NGNNszhDlStLnDid9DPc4T+fkNcWB0xCo29KP13m2DWG1FZwcUkkhvwHCSALMBoP
Kn8zgnabJJDgH15amkTYyoXxKsXiRDpXjuLbDz5qg6O8sA2UpYK7L+YgHucfW22X
YVzVN90Ep0UMa/jGLqu5Kc9ajKgLSRV0Zh1Z9qnKh/iYCU0KKQ4jgpDnMYriKYHi
rMuLaJR9or4goKGh7ozPM4mnI6+WQkGIvLmuAMkD14lZFPgEniqf8LD9oStwRpSm
JT2EV3xVCKT0tyAf2DZC0vXLR6iSlyHVT7DXIudCofbqJGp0S2abTCimPAg7Ag8J
atDFzGfDhfLtEK931vcTUEHGrvhakML/tY1b/GQwMHtOnZvVIMobRQpec6RM+Dp2
sRVIAM7OJfhIvbFt2uQHobclq/36ikW/bTIDQV2ioUPy1w3GwfgtWVgJUEX9p7Oy
MJKD2CbMmrUmT3AFYChOoeKUQlPN2TseqrWpnIcWHcB3dYM2Kqdtq3lSRC5JfjJp
3alYZ3h2sEc5LfvKi4d3XzXHEIX5LXt05ex4LazYkZVCYpd5FGqecVYIx8P5H8Pf
D0bhgtFDP2WLou6yify5Rpt7sFzoqF0To4s5/yVyfQ1V2cMYO2PObEZM4RgGsOtC
rsQkgDX2Rm1kOe/+grbGO4z6ocxhqTFYI92daPTWUKzOL09OgRYP5Dqwz+ADR9LZ
PoCOggA/NdDpY3vnPWHgqF1bVJVWjbOGCFrEGssQtpwMKIBmcmZl/sFRNpqgkeUA
/1TFQRHeL0cbbDPmb3HqbIPx/PcIqv+FzNQjDlvq9yIca0L/iiu0V5A0ve6ShieX
lSaGwBiMZUnmzJVqLbcuBt9CNR5nqQi6VirUPhDsrQIZT8XFAXeTD+5vGoCPexnG
Dett0iVjbDhw1zUmDtrrZyRlIg1SSmORxqBvay4SSYQ/nqKVxcEq/llj/7u4U6gw
0DaEppoNSE11dtX3TAqFgH5bwPmV4FHAkygZX/JGxZUKAGu/wBqcGl38VC6DXGFC
Uhhvw6/S43hHxHdsDZDTW8jOhR0z0gxdGcl8ESS0IlXViT6M1KC1CNmps3HKN1Ip
fEt9d6AWP33gpDVssOP/2GWQTfQXLptfxL3J812tvKVY/1PRZn7+QA8fxt6WG6Vh
HQO08UvdhjdWl0RjHgPIFR0mFks4CFrhCLv6KIYx8+CurqL3mGtyKD00bXqghp0n
uU2o9e4fLjVxa18WkP5q+p6HiYFlgv9gCDOWlbrFepGsiP9CMcjRGgDdPAVOHdoi
UdBOS9Z/XA6Fc8lm2No4U4bLNoJ0LoO32nR07io0mv5+vHqyYxAWW+jWTyQkRDKl
Vhk1Kb8Kidw3PuSddVkywhrrB8fP8YPaqu3UsHa2AP+KILm9Fz3cT058vnuv4cXH
YS5EV60xONmrNTf82ep4bL85TuWPuTZNT83ur1XmzAHjxF+GFpQjaO+BOunOucbi
HqxRWCyoxSgldrR4JK6krWELerNwOu3uicxEHOuXFlDmI0DOmm/RcvRsO17/RRBP
JLVCBK0jBmDIpVmf0RVhAAJxkOuwny7HPxtVPmHhYW6F9iS2Mt0pOK+A/AsVtdix
d58C6WX4T2vjtgq1HcyPY+/US4kztOU0U+I9uDPk023bX7EzvQmhRmHfPCZMa0D7
Lt83GEvvifrZcCiNa26M2CQGybzAVibI14Gqw5Ff4Inw0XkJORphhiTlOs/JVSgh
J4Ue6whggBy8ME1goafAoDJla3qLQSCvuqyPnYr2FRSDj//imZgcXtFHwXOs4Bse
XjTWAIYx9e9cbwpcyM8Nf8eaL1guz1kTFAbp+dFApz0O0Jzs1FLRxmPU46TIE9dU
oPLI9LSiE/6QYRObdeUYwLEIKq4xvjFxD5cEPIFrs3pJOFHnXLqH4FAdikK1Nxp4
faWw5ilbpJgqQhRRJGoIbcWPylAH1aURcyEkFdyv8H4sy+OzkqVTyQUnx+UVra18
VBxkJiAGdClg/qRe+X97j1z0wLJmKDJx+UTz+yJ4atFelON63V4z42qTJ1hLegLc
bFBm53ThSuWgdskCb0tr5OmcXub7tTcwimxGhKNRvJSxxmjxhT9MKTDWrNfxrzSh
lK2jllrOlw99tdAvbcWjC3Ibcm92MND6qC6CUWkWP30NjkWRPVWKcthoT9jRx+hF
j20nVB8+T3BEk3EiCjD7ifH0enQLnCMF720C/6Ta6Ypebi9YCHlVGOobgLu74LSp
Ho/npZmYfhthAkbHeiYxnObrIGEm+a4euzABjjTmB0jLrBekXj8k4Vt76NhJpwbU
FvrkTk+ViuOOQaryqNlk7zidvWIoLLOeyjGO4L7vU3xO/lor2f2fX8m8lpodP6pN
A+tBAySkmQHmTanbXTFLZKS+hfzU3KyeKUA/sMyEk1z+zhFjlVClgFf183JRry+U
7xtYHyV5GY8ZW7pY3pcDXC7Kk18BKDp7s84hjU5nZwJqSSpGi94zW7nj7W+S5FoG
TYzdf3Z9WhkATlAbxbD30fWLRF68AoKqnpX5mqRfeCh6QoXwIqrrU/r53sw3pYHe
5HtT1QKGmGmTdz2HHnLsYVcJd4n6cBJFC91cnmvY3w//yfnoIF59J9eFW1Bzws2S
ldpyFQ3qTieZBJG7raznzCtJFmNePemaflpVFSF3V7lZV228SDabQ/BxNpqOgiIo
BmpROQvn2YffciDBBNh7Qjfe/gz9CM7W+tZtSAF46STDNpH3rSwzYiLNcyoSMTjS
gKY47E2qCOwkg8/5H8JF4Lt75uCTot32B83j7bmK+roNeB0koulR50mgNpUoCjte
xdz/SyhYI7dlW8U/L0O+760SqpwfHJW3wwKJPrUzVAhtvOUaK1xulvGxVMr6cO7P
bGHzE+p7Bh+yVlXbDoRh5ryYQQ9EcKmIdlCjN9jenG1xbvRBs69Rbft7jYpS8KVh
g95NbllV3xi+ub1xaXxBAAqdGWViYb8vYPTFgFP3Nn7cErZbRoBvKEfAwKF6sbK3
r8q4HjPrp8UduVQZVbbN/yJPCwOxNQWHml1Uvy1rMg+uAPVWIZPx/pQaqW+J7Sfi
l/yBNsr1c22fV5huPgNFg9Lf9QSFrCENnSOr0/ZpUrRnjd/edUlhCW03NlbcZxi1
7fpiuwkvs0OSl9w99/smnR5CxA69qe84NlvU8dfyPcfucJKuFAU008jORK4Ou/xE
ZYakp2WHS9mXNmyE/mwpZnbAn2TVK2qIOTcsb/fpik7Z5o3jxKWw8yd3vqHAeu/8
4K0Zow+iYv+KxFWCUEWvQpVSRpAmw3/bXzAPeFjEOohxPEQPdxsVA4yEffGp45fq
xGBlFLSonC0F4bQc0asEdt4SaMIqf+qFrt7oYB9QdOcAAru3F4HX9Sd0rEUKwUp0
E5LVvbm/mQDUuRTS8NmwLOHBzUyPvn7zSDrAkIQh00fh4lmmmsCMlVgTVNsgX6ak
6K+3H0VD8t3RqIX1p0Orw11E0H6kN0WCgerA23s3U+26RPAKZ0DhUiZ9UfCJeVk2
wbs3V6X3dQzqjl1EbbFnjI83s/1KXl8s19mmrTejLBEp2ZieBsz1foKufU0re/cT
+Gnu2HxLNo+cvYlTyuAMM6lLX+himl2xNYg06e0fpKeJzxdo4Eki2LFkxakyCvxW
J26dnSOQ74AtPW/3gmsnBnmb2Fzf2RPLzuFK+/EymoiO1COlavuqTrZvX3CncCqR
Ke/Z95+DJmdfBgK4edcH3NWGXGoTSM6Ghtpu06i4sGBLwkhZ0CFpnCve6gVGryaf
w7XuOCnX5iUEEFoaF8DEyQk6Kwkcrs47Rv4+xw/AdGfvjsBHXmwONCjvmyPwbUvI
4oCWDVzha6oI8/w7KMvqnC+9nceuCt0V7cSq4iio0ZSwFGu8xndW20UUiYgj4Z40
29e97ttCsOQNKWrEmzAQ+1gyXkKsyUoMF1ZoDjCM5h5VLjh4dHsmMWQ972lZ6yju
KmjwBlWqP1p0GnQ44P93Dd06d94AWQ7iPS7GADsOkUqrt1g1+q6QZHp1g34HMch7
nZtrDfsdaFQpQM/iT9QaxyhFDIdxq3oJhsmzR0SnkbW7jgaOS2ScaGEvf3X8q6pm
dBLiYi/ZVC/HJ1cxKjNemF+Q0HT+7+bnBSjox2ELPEnWjROFahEUri0PtcHChzXR
HKmlpmAv4YhSVj87/n3ocquPecY7fyiQvR4rWKR8Hy904n6lhHthWTuoic8GRkgi
/wecGvuZkjoPRQoSJR2z5SGoS1k7uv1kLmWD94xClCA3Zg0b7LII74me+M9oZzHU
1R3zO8nXR7JNwOiUvbOrWTFDTlHODKZDIUuAFwUf/Xj5NnMvm2HzqFq/CYm16rqT
rKGsPrU9Ya813pZ0hkUAGjUUvzXaBlUEhQdJyF/dMF3bsbx0CNi72GVn7wyAytVs
FKj3ULjMJSWCHaCy4FbXgIw527qpJfDBdMrZ/z6M7ugtgRbEQlp4GjFCkEZQidZo
1TczX2HaYaro8pWiZjfJx2jQkjGAf40zMu0+rcCuhg/7nOYGikBkBcnd4Wnt5GtI
F3BJoeSZib7NytJZIhvjJXSya60uj9I9PH/FsvOXmoUTQb+d5LoHNxLk3CKWDyxM
kfl1g7dchQVdICyjFRTIVkH1LrFFpEec8eSMYUQGbx96X9//g1m7BZwaPQpAWxRU
Hr6GSV9Rzzh9UtDvpMFPYHl07H3fTeiGPiz9jOXvMICutbBPfDlZkHUUYLzKhJRf
6+jkOiJqypvsmGW4Ovr5IeMc2kgKBnrThLgyIn7O/u3w8G8r0Sc/XH/M0dWxvHyl
Z0A01yctA1BWoMg4eo43Dwazf7/9WgrEt+Z1W3BZytBDVnRxxzaj8tjlnjmE/j1B
dTIIMcEM+vFkvKwD3H5oNNLuIEfnWRrKRwdKGWsZkfGOKImPUg7PY6CzkSd7FS+d
e5fhq1QckNfAVUIuOigmtw36hSgzDt0Vhu7mursX5OrsrjX0FGBmgXGCuHWAu5L8
RM9wNd+Z4Imw6pirW9K4BuiKEqPgS0jdRhpcCfAHcbDe80bede41RRn4laD6CF+R
w0/ZQUEG1tG8o5oTvw4zphLXauap+f49zoQgScL13fdtvuR9e3fPKBCI4U04VFtf
39aOrROwI8vyyG0BA0phJuTR3XyHLwaOBR7i2FpflsEDgevPwzbgSsJ8er1K23Iu
krNGsqyAaHWqmq5cElNFvv+4hK9t6CEzgbA7eTC/yNDOY9wbdzONSmYwb5NmQrNL
tC0LHimjktIE7qSo2iYauO/uco0X411JbxLf9F5iA/31SCzshugBi1cus7J66YDo
eHjrCAIXtgbOKm84Q9PaZc12TViCzY9HTidTNgdoSkQhcXXGOigagxUZtOYI2Lud
A+98jMS2aTiFsqqn76v9DNOQRESctS4lRbrpNXFSSX9lJszKKbLnc+RmAcv/CpUi
jY2AFtykPFAuBHfxPkWOjNegPQzz8X0ngxYb7LsysH97MqSmGtQF8kUx8SVLOHur
nIEEaFYEHWGu/LZua8Npy+OmgVt7Eo7fQsP9M6RH5P8W0PN1B7s6NDNcWrIOmbBG
NV9puRiM0eHZPVZaphL1mVyqopLYahh6WaZOe8txCOzGM6Cl1z09z69Vqwk3MumP
fYcILEacUzeSlTohdLWjxaY1m+Rs9aeKCib9wac1dcQTz9lifqm9mqoiUKk5UnkC
6N7lubG2YoXr6MTXMXi4D+YsUpgGQ83G7cbulaQsxJMBjshc8nr4I9u2q4Y0uMhK
BdM7Ig3klS5uquIBj3yKsfUZaiBZ8KyyHc0LwvsQ4ncjIJkSwG3MW6FIi4iR2qlp
fXC+J/fkgW/bcqq4H5JmhZ94OAueYgKMEdDUHYJdBAuMWz3K2IUbfCw5Hvtvp6ED
KKViJKIqNdedlNWOEhBirnJdL4PgGYqiG5aADMz94ZuPSnZXgPdt6smZYTWlpDdM
EtqIvqbvyefBJJFuVqkgYCXIfJU6xeCeSiH7jGPkW/EQVc6rSD2gCzLIoz/IRXos
ljBP2kbb5aHJWRfDooG1HjRzFxjvcCVKFiDdt3iWh4tafi2dcwIxa9JH3XVQdJju
3iKPxGFBZuRgf9fqq+RO36OKNQKa0h9kYlpGQlSAnVw6PRyGfMGa/nzForoxtCB9
xNTu7Xusk3PEFINWkJ0gtdIbqGSrYJemOyVDFX6u43swDZseqK0BdrDiOQyuyLWD
Gg+Tq7bGg9SrgCOxU8xv18PbECBd11Rs5ea4WXhPN95wTLqxAyzOceSWjZtgXaIB
DCHi7EyFvJzcTJxnt5AF8ZCAkrodR+ZX09vv93QLX/WEP/CSSWkJP7E/2CUIan6Y
wIB91tbiVVUAlSKuqI6hSN1zklkuRQZx5nu2HD8j/qaROZlT2QW/1iVKp80LyzaS
GRnE5JjKQJU/JVmjewogp0gWeZXE4wVnLdP5oYMWdc3q5Q9gIK3e111Qx+IMhcm+
1LfOMYx6S26LGNn3MOCHIBowsnAR1k/C1/w167TH/wtlCdX6s7J4YuAQTK3NR5BB
lbMENDaCw0P0ZrTw17dxigM6z/FYUYYKavuEBbR85CvJGkeNVjlKdDY6AMn+LFv3
yLejIPKnVaAsi51pr26dOwJ1cuHFRQ/JmPb41CaWU7Ncv6Gk1k4UbHrAZtRjkvmV
DIbagh9+H7j/8j0vgIJme8HuL09FmWjTnQgGc6//+2fC9unLVUG7rnBHVo+WglGu
hlK5tcdLy73k/AN4jAfmWnIqRiE66XvdJaUWU8WNYgdvq0XR78xLh2eT66OsB8kr
q2g614obXIFVaw348mJI6HXUoPz1HSHOD9KbvmuWugHOhgV5gVkh/uANEme9P9s6
clAM58rvtxNuK9EoR3VNeg0FrCNOWjLLz8Bv29YE0RaSOz4MZIRwk047+WqZajdM
4LBesc4fMRVp9VdN1GslHD2sA7J4zkIP40NrkmMJjHJbTCFH+N4fNLC1eMA8nDMW
DOZkXaOJikaAS/7cDChfeW2+/rJbozfh5AObU+kXpHfoYMGL4Onuc+7wLGWfu3hr
06ArLCcniu7PiLezd8IF/tyvVHeU+Sx6sRF5t4KDqQ5lj2AWbOpJtT98OQXzwC9W
z/yiW993qqy/ZrqBRc6QkgP66bTdsIxlP1WWlM31D9z4eStXx2or3H5Vg9MXd5zg
KEL3FXuopMmDTBnkT058QlKjA5Hk6JIuuRCw4uln6NuuaymAvqzUvHInHdpkr1Gx
VhhWq4WWbw5O29TYwIq+vNLPwqy9osD8NhGo7UWViHHy+xWU7URExYQFntQlyL8s
aOoNtOPNcleUAGxknVPdsEGJtGCl43jFT+bjXCaPeTYbXSFcQWpyJlC7s/Z/Tezd
kAdhWzr4MyV0BQc10wW/sWUd3C2Xl4eMBQmbKh5xrWMchEe6LlV63MT01sCPz56e
e55os3e3PN0Onn+YF3ND2ZdBmsRbRCBVtoecrcDkDuF0a3tswJJXLTDh16ba1Omo
jFyB8P59755eJkdWZMmHIBUZCpzxEWHOT+Vt6Cs28rpYmgOtfVePeHIG2aXRCppC
ORrWN2YNmWNlcvqiSE1FPpMQJt+kaeqWKMrdpdiBz30gmIDmk+s4Ii6Zp1ZXRm7V
Oc4pzId3uXkcb4lGT9TC4/TTBRVsdGkj87Lztf710fpxoPwIUjgpg9hZ3s6MuSqU
f4Nm2vcWgQkeg5MvtxuqXYeOvP/EtsolQqz+utFOn02vAcJUOFUjPTQhf2/VeqpN
b4vr2peJHrsu+IrQ92tp/jh9fkegpqwIyszlN6wpbBV1jVlMhW67/Rv/NWd6NL/f
FYfmXUAYcla+YgequWXGGfeNsS/g6DZiqdPiw3NzToNMf3HDdmdtSClnToUnQpj7
A5orfvrnw1JRFm5oiqqfP1b52un0SP5LaJS2LCPSvQFS1jsyo+3IiHJ2oXSEH1WK
JZ+50FzppPYOIRXrdBPaxb/yFrORK9IfY5xRNaBO3bOPW7tnhLEYLkLJ8bGVjvlZ
+jjNhLWogCv0yLn7SS5lBIy/DulVEE545+XurCQbi58WbtkAXLn+/32VIq9nNaVl
xSVLBPln424Nj99RhjPAGaJwzqMEOyisgCSCN4uVF+7wA+Fd3BppUTPo1/q6yX9s
qhbwgKUYQvbp8khXrs7QC583aotd2zivJQLyENYfCyghnPtamGsvAtFvfkR1Ldan
rOW1pv2l4UfLwv87rPeDvX7385QclCVSIxA3/GA6LzEuUw4eYGOJJPsUM1Cv+F4a
pJUzYkvUcWZMmkJ/6n1r8PbZsbNepJRYAhHOgCPlffqiTltiUBOaiXclfSRQVI+2
FFPX2pjNmxc+Ov0zXBN+aG9S8pooPuW821o6kj2yOF/cAOyQEcuDy7V1fFyU1FEL
gLRh83m9zsLJXVdaSou0RHVL/zkyj9fsnWtqs9odLvTOPtFf4aO0mefa3yzNinhq
ODDlF+ByZ1jrrU9CmIzKIhumhcJBJqHTAzenMJlqK9t74mRIQgUy2D14jJfYFg2N
59B2U4kXkQFSw8x0X8C98tjCHh+wI3LpSwNP/TGeGGJHp3OJp+t3AcZycv/+8xEY
thgwsHc+uzz6hQvQaEnTGOl39ygX1gM85Em4BFM0k2AuPLj/oBQzpA5aDkuRKizb
6p2nLD/31PZHnjJQU2rG914iSCWMu5TfSlgFmpbSqZg2gnp5vg1HYM6MF+eDOZ0z
sDQiZxzhl9fWjjKxc/pjvHqi5RYHrRlGhhN/4msNSl9fma+t+hz3dLCW/kBVTfva
jj8U3Cdhotakw6a+nsiGL+L42F1RjPPzn0dm03tUL4ioFKJifEI2exgQNCtqxx0F
A+Q9G1tvpnl9PG8mqChG2cte/QE5lEjjXDqmvUX+7BrAW7AZgQ4n6jNHaGfvwBjg
wAltnQTouoWU5aY/OTSVfmIYX96XV8wEcu7Mh8U60MmPiZU3yStXy40/dL/kmjHO
gfDgbU1NjozbATgm7taWBo6JlXF0NVaB5OD9eVxGKJp4msv2UQ3YA6sdTsQR29X6
OoOtOujRy0lFLWzZI992zh2/xDc9vJWwavJDfZOG0FJZ2i7VpPEQddoWtXBq6Kb8
ZlONEAjVcz0+qqTSDMjZELEyCkN2qDqRtqM+M7NqN71p1h88FxlI6eBR9VuoES11
gMGQ6DN8iKS+UJY6QGtL7Uv7evaNRaCgqyhNUerkdXFDeK7StxjxBCS3aA17Ir3E
7LGg2K/JoaDVbdQAttzOLScC3tsCiksGjjXiDpzaFgQMQrQE5/c4opdtSdKluqvE
9QxLfQ7/isQWUtHgyDKBlpwqBnm80tbMJyWe6ZlzCfWm6YGyYaph1KrgjvE0u0h4
8y2NZJt/fnBrM9m0HsHSxLUK6QsXWNE8Xkwbdg6sQIEsa6j/ccQK6Rj6+Uz2j85F
kJbxbkOJZcckPB82WA0OGCbDVwH/mj4GbWl1ijiZpeEp9awdf5Hx8do3OtXaQQkO
qY0BLuEXDSAN8WkSa+LCfFNeYAppmiKs8aFTvI5TnMPh4ru55HhdyA98fB83k1bh
0ZxNxio4REDaR/WOFEc3J+lfy+rPpuG808X8Q24S2n2P7Lh0D8oauDtBRzSL7Tnt
FkI3PKrbBRleC2hHEwMOAAcJMeEneIC1Rxx/RRcJOMLjVjO5mC/46zKbuXnOVkwU
IsW4RuzriKmVcF7mGEbFnMSWtcvzQg8pDX/bc/XrfF5clAwt3JzEyFW7pQILzlKY
sUv9DqE630fg2eFmrGHDiqFw2g3AaYxp2MHj3/Vqzskdj4jPftZ77xo/r6QhB3ES
OC/QYQC+iP01igigcgon70Yfa+e7oMjvPzw0cXrcGNxpbxYYQvj2JyC6DZul7var
bwfY4Ux+v4v4S84/sUCtmGbpv0Hug6vQzoc566ydI8z6e3yzws1tpWGW6sx2Gr3k
5ZI6+2U+KfHE3Obhhs2VslM7npvbLCaVzIbnP5YqBPBefBzWnmGZ/a55GqG2CMU4
1XY6/9pudCAM3RVHTJh00zhGoUm9fgUiBgiFH0GNN0Vu7EJnqdFsMrvjFvOsojon
Wcmoyd5yeJIMmVoyU3J5W24+Es2c6qsLu7ESeeuWnuCSg4FHW+WBCHxqxIMQ/EGh
q9JmGW+j68d4eGIEaIjIBvlZo+vZYkceySl5XfEcdrzb67jPxegbqncbkrDlTiRT
LElNcuE8r61w6fcE/sgknNIqJcP0vkbKp2eSBszSPkQqypSNrMcOdth2MB3Hr/sC
gn9zcisIfjVribYy2AjOjbvyTUThQEHRC1iad6Qxb4AAjHYQLojebWjur41Zse0X
0SmjivGX3racIOMbdMvjyFY06Fce+fu86mpvReI6qbh9Fu3R8gewQDhRQlPxIgOO
QpIxkFzqgUGzGdSjXk62CG8Ysxzr4avfMUHNOycku1aVi9nsf9XtOkdHbKTZV+Nw
olCd3lnoEp5WZ5yZcciNlDpVVEdx3F+yFPuFxY3RfLGEQGSrvMjp5qTYMvl/FL76
FZzGj2xzru7YS3oFhGBB/BeVlEEaTsyJj1OXNq64kSxFa/ZLN/6odYruf6/ZkRx5
TsDgvNymcU179y2ZKJuTfCz09OEEH51sAciYmU9QtXVRo6BGRy1m4iIEGowuII76
LkBVI1MriLG6zkPrX1VrvZnKaWTNTeODngQiXJhFiM5+oHnhS6CCrPOfecMd23kb
JjRsAwSJjv3qhdiBCf/f1tRD+atoYVAW52G81oRu+0EwV+Gl0EBVZMAe6NBmaBwq
82PmDgVRsP1ENfqq0Hm+iEXlJIjS1bX5DlrI98Zz1RYtYQ8hCFGePI3YhD9Dx8YE
bwofeMSNGjWphauuXO790Y95ruGIMmtY/7Dk+lkpDOi9jzEQg40PqgbaDs6H3BCr
VMW/8ufbTfrL1ydEIDaF4aItz2P8DCEgFUrN0mUCEMyOYzr5B3dNLnksYF18LF3l
ZbqcT3hpZFPCuYoEQFsqy594mm3HrYUAxYzVuHi5IyTsQS9QJlZf/u7jQ/poqYW2
csZcJiziPxoELQnyfP1NqnW4OwtOCE9iSGwCVyQi0K++Qr0gXU3ESpgxfiReG7Ay
tEwIjskRTT6OCx7J0hcLoPgeMsWpdPMzKrtSW5l3H78YmxH+KDwlMb8dUtQGQSrQ
DmxZNJZRcAmxfeWsZDcuzlmtUWJn6aF+WIMvKmJ5tzdXAG3tapg2vFQf8d8IkOZQ
N14y6R1bLJBXTGqll0U23eKkOQqfl1e+n94AQ8au7GR108SOjOirTdBN1Nu9mZ3S
kGSRRcZofIm4olJKzXY/QVWlPyjDIpCSZ44omDxiD3L3t6lVtiGgXlbSHc/zWA7c
dHDlDhrkMc1JLaiSR/Wc6uNpLQIRBp1vV2fp19NRLLhv9J818RrCFP+B78Ph6WId
Mm1iFhv1VStcgLcUYRCLsY6iatzAHuRjgBR3Q+Avv0LgwmBqiqKOXe/Ivp03g9Us
XXMYCXjJ2baf9oeYzwhhVaQ4MbtqfpWiQBzkhFGhaBw+FPi3aU0I0lUEmL5hrdJf
cc63Ns6RSjjJoQO8HBARb8N8yHTLpr6O83dM7IU+BpM9T49axozmoJYVRZXGCGER
Ai0ZSmWtDUT08n+8B7XuVtBOZJceOM0EZXpLi+n4pIZJCvUwGJzKL3K5KPr2viaN
IhyKdyOwlZbuySq9H9KB6uGeW3h9AwY6xFBXqHSprW8KuP1MdKtTfmx4PwMwDszg
Trcb01f8nL+92nDabf64AreEUeztXVzDqZqOGV2ns0+OzilsVP/0AIhBNslxdHde
8x5ovIpICKIS+2PaIWCHCRLtR8T2VfeRla8mWbqIbKSK8uBFGtesessFUIKRo5jr
UyhksDsQ8+KriPgKNlrJIe4MhqycHM+8QovHnEzNT3JSiN/4ZGya6h+YXdDzeZ4B
RCWgF/d1BfbYJBWxuKM++ced1fKCdC5Ix7UhLAY9qRoyoh+2kRRAJ/OuHtI5lHmq
gw3v07xIH6h6KTvHRFoqKZatqlpBCk6/ZwesoQr8coyRiip/LXZEIU3yMbZTfNdl
Q9Uv683/+zw5ubPZQUj0vh9oHolyYwk0gA91M6gfEVf2iD8BJVjvXP6ppZcg9ToD
6DMTS1WD7pLZxyXOPhqjh0/0LrbZpJRGtuPJX5TfgoflSNhn9nfhMY3D6b8wEi2x
O6thww4wVFmEfaUu8zUI8y1EMJcJ8hfipB9BrnTUV0UZSn9GqrryXwnlZmixz23k
f+fMMi4m5GArK/OEOKB2VBl+uEYkey1xYLP2RGq0ygVNttg/QOxrMWsiqRBs7F5X
oLOhB36TREnYrJHZGN/ep5TmOrE2xV3u+I5ZjA2b5aXDcBKA+Rrmx1NUL2gOfhDc
Ehv1pebtiXs1/wjMlgYZkMj3bORYUf/FL018yCVebdUWwniUoW/O6zl3hTa0quRj
sFEJv/AXSkdjiityZrml3PXxPptHpUlsO+95SD6pbVC72LLdLdmMSJgkAa6lpwBW
zFa6+/GUYDaSu62iNrDh0Zug2gwVn41rqun1of1b9gSbwB84POFi4IelmYyquVJK
G7DXTlEApWB1W11mN8/znwqfHdm5KbUInTpGa8RpYeZsfhHopFnZ03FnG0UkuAEN
pbvvkB57L/c8eCS9pAwx5LtdJE3XpshAWdHVwxqTRm2LlAtJLiZmBGqe2z2l9pcZ
j/ocuL+HZVK7CTiBOPGUBFeybBw+5Ik+6AwsWO//LGwVjGetjhqj7W753ejCwsAm
GXItzNLW5t2ayEnB6YI0z4S9Q1p/M7/1nzX+hWdncroOWYhiBQcsPT8P7XZZk2Df
fz2Wxc94L/eyGFmkLhUza2gmeXQ+9RKNXtXXRGrWYqSgYLWgDRuPBIEBJL/gfEzs
Eq6t0wMjnaFAcw9QhNe6T1eG86QCtOxzvME1h5Zm1ct7zdL9xmRQBJtsDA2wnrs5
Zbm8vifl68VV8Nd2AcDtfv11kX4YfF3pvbchxCXQXrGZiXUngXTURG59CKQWRgY7
cvswn5yRF27JGIc2JKkDaqTDxpLsIKd92kOGppSWQKgMvkYFcXpIm1edFxkFk4Lo
LVXD6OFTKDJLcqJzpZltkeoLeexsG2lhuUY1cT0HFWUGg6fXEQCb+pbtV1w65gOX
YPSdr7Z+7U9UfrGZVn6D7vumkXzOJhTMEwJ2EagY9UMNHEKQZSVdDTV7xjyRlt3m
03YHv3vg3XvrmWnDYzLwAdu/pEEAISUKa1FoVIl3e5feMko4DtBGAetKeAd+DFUT
rVlk6ZVkxZ458A8TAPH2tbhFJIWTgo9bnwHzhM7nVC+5QWmR5DWCdQ9xYtHO4Sgv
weupyd+VAijUVqVA3NRf1XtwdK7GqG8Tn8o/0sDJ5g2vxqrX1KwCamXSk/FKvCKO
nD/yRLJb1TrPnWkXoviQuxrD0GJTUDHllrCsLD4FCvNVZjDOmYQeEDIRr2uAfGAa
DCf6VmOWrUiNQ37SBaVv+boPeeb94uXUUVRsBekYzZlHxdBBH3px5FQQsPlTtxKQ
bwx7JGFkEGISyIaDYCVc3huw2fg0ARPK5OGYB6IM4/okwTG7lhad1bNttovI+vUa
IalExxclkHaLiLisSUfzx5hVCjanhnG3PpAYpXdVkFcDn3Axj5xW7k2RTJbXEpPd
ECqfW7GrreODvNaCiu4Ocm1TsP7nu3Jg4Y7SGWSp2+LpzRwk72DG1B437VVZJPR7
DVbB4ttykbXIJ0J6dvVWB15RGFPSU1GAn8agPIlqMAcU4xStrYNbRQTygqRXwY9T
865ya+HC2ub4ccPxSZcNVhDa/onHu9vtxCJNaFCXg0cs0D3nQKGKnqtYHNk2mPoc
NjhqDRdbdhrfkVIY6Woq8SN2vlcr70anralyZzJT7usi+Kxrq9sEt3LHMQtQovGi
LeFh2aexCTjySy5b/n7bBPi4TOZ2blIaDB+GLomnTrlaxjKHiqTlWD4vjijvm3Zm
LPnbUt6l+NXXPaNFsxqjL6rjyp37KC0VJBIhEK+JBHRxDiKphcuKG9dGsQcAnRVc
eLyrRIVY7G7SyVueRBUWppsDAdZxYZ/PdnyG2hvPEI0gItw1eunBc8KiGqqluTRU
SHbcwSpE1vP+l/NWdneYjNvOHs8t3FshcdnDEBWH+cOTJJ66y884d7E7/uPTcDJx
op+VOnT4mW46QZIoPStjUWXFwH3cecRQNBNc9iZP1dL7SX4e1Uvh8tarUccWL0Ej
v7Eom2V+zJeRZuHzh90LA3IcV1Dw65ytJbpiFAxeXCtdfGkSLYuS5BcwIVCrv4w1
AtwprONigT2AZmXQgKpWERoIhRw+1+TwYK/uxqjohDgaN9uLXjQQztSFQZdc3hi6
klxtoZ6yszqjs7UWHw2d9jvVLq5WKcoBpW5/bilTQYrd2wkJ3lU8H38N1oMusXBD
8xkKmahzXHV2pZLj7914p3H9cmZkR8ofT14SLl7NmAQYU4GDHASS9RLlA7SLKMrC
oveXuwjPQk6W1ciWy4o7FxBs5YNYtkWL/x3RP4lZMJxdxTVU3YjPswbjodyvdX6D
cjuuIzwWzgpGtOOnVupPfkyUNzctvmy8atpslplf7exVOXRIIh7b/ZIsmphgFvLZ
0iqh1OC5Z40qwsQsU9qZrAkzQ2ZZdD5/MGhrrh9/enncRqJmXJEsknkBqtVnN4fu
zLVfwISgVjQBw10gsglCG7BZDEBb+snWN3dXs3wPyvrJF5L9EV9Xq8MrBzyhCI3b
JWHpH4DUpRetMBJZoDw+F2CX4j3GEDEWJkZhCsEXjG7rqntDWCFDNALTmWq0cxvH
cA5cP7TMfz54O/AQly89trjOxDD51GqsUbWjH8ZhtNFx/rkfc0mVffzieIngfzkZ
VLqHVe2DiJGDaF8W6T4v68W9Edww1sEnwwCkEMaaiSj9ehTXpiNH3IWJOCkSncNm
VzEKnFxNJi9kURw2i8dEyvzYL9CUK6qrf24Un7Jas/OoynDYgIv7gqBq+IX6kVKn
nr0lBXb+f8uH41gqKy72gJ9mDRd9frNi1b6lx5MOxpIjdNVN+fzmYAgmV7q3mg+A
QttJpi6fqxRzboTfR669tZfG2KjcXKprUUcWIFHYtOt4OZQhyJF6GugcvZZ+L6MA
cTjHskUbbPtRzA6NNfgNf05Z8SQiab4WZqsutHqTx7JixeqwoLB0kO6c/rd6mZcz
HzOGu04glCq4H8CKXmybIKZBIDze9mYKQwYUeAHUMzEKbhO1DDx0EtsMGUrf7oWa
qCIXwHqe7SF1yhSWO3kAKhX2Nmnob13YPHg+SpGk1j1Z0Mgoz7LRuczb/0/A/2MM
S8IepCyh7iYRA0L+gKfx9yMNCrrLjXTPgt91MYAmQe+n74865GasZ3vI3zjgQ+rN
Qi1KxCeXd1CY1zsKYSrJBIDSqq8CPO0xpNJJS51hYPfyhS8cxH9i1cqPJNcPzyF4
wAMkZbSAUyPy9PTfZJ9UKdhc9cM3ROaIdrg56TQS8qF9617Kh1CDnlcVSJgB7uoC
VydTfO1XjBAxQ7GDQlFIMOwOMTyYpa52ZBCQ85UGQ6DcbrWobbs4wSK2IW99TkSs
PoEjVtc2pyNv0OdUCI44ghZC6WEyQrkHWK5ww+OQimhfKUANSVfa0IK0PYg4waNk
UsalxMftWcThxv39j0ylNZ6KGrVnz/6c+AyOVlvzMMUKrS2FsieTyNV4ag7eCsPs
aznwkjH9VDhrMgy9nMVRlQdYwgM+vF0N0FbnWT6gjxr2nRplRQG2FhUhpAvtGhR2
KmtQyc6LZxKszrSZTfIYlO1tl0kwBmqttgRUXvVhrazHQ5Qr3KyKb6zBpVBxsDke
79WnAPFNUBwuCG4oiWKq7leQnFyceOgFKM3qUFBWSdK1uoC84QMUc2SbSPcXrHOm
R148bB7/SLs7hwqpJTP3uBkeTrYhPx1ghhFKGc7273DizJCDBladPE4Vl7fNrpTr
mlgqGRnlROVSpTSwmGmdcOu91ZYz/dbdM3F0wq7CxeZZb9bpqYcfy9W74NgoafxO
yVZUqz0RQ7zxzfPvwTclbAwt+bIp16PJooXNO4uwt4z0Wqvjr6cujQga+ACe6vUZ
hP4zW7Ae9DAIXjOAYVWKXl1k8gQF/TJftYtFvojsFYig6tPZ4Y34zm0DMYtoQ+3H
dgOjqZmVnNfUvxqljAV/0vS7CcATaR4sh2culiTbo6j3rPG4leICJE4ak+D4iFlV
2RgfuYcufsqgSTh22Bf5a1o8i6stoxVjn3Fq5ltnDOHjJPnYZyRauSVLscXOD0HI
i2CzXxK2pRmJAbSkQv6GIsA4ieCTza518Iuz49geDIfE+7CebH8af6SIhgDoGyri
BS1TvJgUtZzuoY2YQS+zPE5xY2jhdlD5i1oJ0n64jk4Ens83VTekq+n/zB5evwLq
bjF2UIJm8SEvEUYnZm/VUNL3Uyz7wXIJjVWSYctuQJG53IKDVQpDfUwTL+1PiTU5
Oo7mqqZdSfHxuAEHhyyH5boG529csHYQNH3xKErnJ8fgt8EBdfUqnErShybsxqYU
lcbocNnxOXRj0Kieh3cafkq9+SLXQpMPKsMy5GNrGMKM9QSOO1c/aJRxzoJBSwFJ
J88aHKYNR4Y5L7iSK5vEj5uoMpQ0n/axw96n7sTW++i6ZsZ17zKYD7uY4tl5A657
p7TwC80lo0HR1HsUtB7k6REYwdXj4ccD/iIp4D6UhJJlAZMWVyEFm+nYmaBnkwSY
BDsn9LRgGp1w3+B1nx9DUHA2pwFuuN/AffE6kWLaVIa4lXrKnII6Ewf2AfkJQQIx
bnAvBFtbNMrjMuNgZYxl3R9v6RDblrS27dd1/nzTmYKN5MiC2g7Vk5mHS2itGMcB
Yqlunk89PB/+naAKVyuiAps5EZhQNPHbjaSM7tMWvqT1V9oPY6l7iIbEM1E+dq1r
UpezMPIFgnfGX2bCdgJx/+pVJ+4c/M4kgc3q9YR716RZYzHVBoPV+mNiTExqllKu
sOwh9bwEA0WS3oPBsMe1ozJ+QRcOsfxQ7re2AF/PISgBgsog/Cfb8J1fkCwD/XRC
mBsTQsnT8Lm6zTv7Q11k3PcXjsxuggvNQ3j2AJHOkFaSTe2xFEmV45EUt3WTI5Qg
fy1DMJpyZDY/gNu8Pt7e6Lzq5fGskjeW5qIhfypcv8c01fNZVCPzSJumPVGK0X77
BYkf4dOqA96kquxyaJKphbBi/HTgRZVr/AMPdi7D4JP9rGR8P8LsYBVG5E7Hxy0C
6cjHlSgnFKwv9kauzqGTskzgb0AZm2qwP2/jXNcB2RGpA3p7FXA5EFatC5s1VpH1
+DT2Iwl66aPaUnB8g/EsGrAtcZnXRZkchLdSQt0b/+u8k3K0TDDT1rKoseLB3/hh
VblWY9/ygjuX7U0r4Eu4qC7DtzhS45DGpUESeZEEJnJ5HFnIf4/oarjg5U6fF4Vq
5DciMyj3bQ5Vb5+TJ55gS1otolChjnIgMygH+TRVoleB3Pbe2UOMHTsNM4bWUP5P
r1hRIutRN5Tp7ks7My7z9ahIINVuXNwMAgyxFz+jThcN9At4QZfRTgCyARZ6Dpzo
aH7Fek+kb4Ei6I2h20eXlpU5B+7QZvNcppLXSvJNzpsyByHFdKItj179y2vMK3Rh
aN/PCd+PpjYkSAWgisNlHqfMHBr/4cOUFtR0kvtAB4jV4joA62RWUKcEppHfLYns
ifpbSWdAWb//KXaHYu5JFsz3sm8+5chQ3OjaykZwFVc9wJTltfv5tDQrLvm0TUtu
+AHnKGzS3SbHA6MPKc4NrG++Ej59pPO8/KyycdiGoherRXxF09UW8Oi8uZDkDWwY
yRa1vGCQm5ER0D+t/JdfXWJoIIrnQSDQN+lpj1LCb8xGB17I+RnWIKLqk4ckmZsS
+WgtTXKgUnYsE2I942HA1ZiA1ZGjxmZNtRuCaDOP//sNQ/CeYAh7mdHp6twegv6C
Fs4CSmm7GlcFEbVHBGJ4GyPx01vuExmCX9xwZsgKYQTVMefvXBdRbdtzjn8/JkGH
984xmFlvNFUgHCo20eAge+okbR7pO+J81pot8vPk3ZaBb1qFkNc+3aJHUcRN3oVo
l51auhlx+bI4k0cVpF+WlqFkqJFwZ46cpCV0bclByi08H0Xn1EQ6h+bbKsEF5JU5
SO9IRiBX8jgjVuy5wPs1buv+37QW7NV7nGOEk6lkWQuruj3DGV96HqIAckqhdA6Q
SXDim4b6lRyK/zxS1TX41AmMa9ocNEl67NhgxnD2oN/d/s//A9tAfxt3lbBQA6Qn
c2DVg5F/2fYkfBZH71vkwttf1Eym/NeunJNVxbaSJHiRMcmPuLa5oB8CctbnzRqe
4EUiMch9iQV7VVfMBNTrlGv+m9AclnX5ExnSQlZNuazy4g7OsUJDFhK2SXiZNrWG
WXksWQd+nVOhoFglUOEjmRALjj6SPl2SmkHsmxw+L35iZyPyUrqerUjMFaw6l8kM
gr0Y6fwKkQQ0AOuNHmpE6aFEU8IULpShfaV33cqSVnyCMf2zuz+MRjAfJP9otfPJ
zQaqwTMe4KkeKaAuTPXILPp9GfeBnVBxPEbFtEnnNJkdrT0NcHgdbyML/NjEUyzK
BhZ5E19Q/xR3EjxsGlTshn/BfLNARkQ854kKCl8OqLtsL/pzDpvP8LlLLknIvFkU
/n7bPW+xiP6uMoXlbD6s/V5C2ojDQLvmJLqh/QufL5CxNF69kwo/eIzdUH3t9XFh
jP74iuLwrofaW38uG7J/avOOSYl2BjV/z/RvBIvGJ20vt9EG4EZ1NpsPh4P8fcDl
yAtJN6xMsglsQcsG2bhfgMtsg3sGApov7X7VZUzOmy2moLD3D5ALlGdNK0m4OxLB
+RkhYs7NKklkIX/xe6Lu0XaOOroF0VU/DYso31uFI1hWixWEB1yOhdsoZJwUNM15
G4CBwwBGkrVtxbudzEb0O1P+NGGEm/qAI0GokOd40XVHvDWdRcLWltVtaetJ4nw9
fhXTJXUKvq+8UH59IbzJ89qq9FA+Z6fNvlPmtOg4DWLaLLSDkMnBcy58LmB9m/zI
UmSR2s6XMhsc9hxfrry+e/FeJoCSVD38pxX+q7famR+qo3ZgKHEj4o0tykXO48eM
3CC+0gZ5HcRsyMycE9mPv4GIhWhFob6/SMHc77QXMYupnmkUu1eHN2xdnGdR2uei
qLTP+bUxqnJh/ZqcI1QKhHTlKTDiXdDITDiaU2CNxqq9MCD3zvqyZU9/mvSlemGn
ejT93DBh/KbdWut2mDzUulJbAoiwPEtlsqNGScyVde75EPUgNt8goCRVuasul4c9
Sr5ws5Mdc0yyH16x8Lz0eHgvHxpgdshyZ49KYQTflrgqXTXo6nYgm4F+FKWJc9hL
8o/BL5i4IdMJGXR6D6JOrHZ2+sbVCpfwTqw4HVsLJKxxzH1PSDUDiX8zDHxF/poT
UYGBzXYF0hsQzv/Wj9CtZjY5q4f3YMqRanQ2i1ZjyH7afhkD2vOFqy6b1Do4APxb
5cZz1Xpjp3cXU8yS5ecX0v5vs5K+4tPQ0EnOTQXD3DrdZsqkxorBqd5wGDfJea3z
x4DNC98WAHuMauBdlpK2Hw3ncX/Hi/jCjIieRJnaANZrnaam961K+2Y5iOM8KQ8a
6cgkMDKMpYDzQMCPh2CQ0dPYoJF+u5bvECfxTUxFQyYLjrD2NGiDtq9BKbJ5Z8fl
zeFqiIzkUW1Mc5+cqeQTrA8suIMU7trYQlLiom25P4opzRCXJz5+y/2VDHlKbALl
uvZBJ2nU45kgLAd4SMeIGsQp83tPZYpV8/C8kMYFUfW369LC93wzJj9oS0p7mEif
qJ2o9KfALme9rsOppURpL0RX7gd5hOoM7R3PNsJ26wWsRu+7J0iYbWG/74ibZ3ca
NFhmSz9rhnXNRzSiBVbcdVgKgxCcgxE2B/wMkL9fveZm/YZepk2lt2t7kksIQql2
HkPCSItFEiIqMoe9doTN/EkKycjyRCC2zbdN/oE76+yP2PNgtnoGDxr20HJeK/Bp
rL7/nuJtnK3RdycNxlqyopIn0cCfN/PgNM9GOPV+7+7Ibaq4dcmIb2HhvdUoVe+J
PvJelwdPyqB4RJqW0vqxFz6+BqPuePTputJ6Lao1sN+9TAlE5PApHh16jnMHeWtO
oEoiAsY9vr28FiuArfhE/1Wq4JMvuXNedCM50sdKdM0HBUfejBK+h3ENVH/FS2IF
nfBovPIC5FWO0Aw7mLgDvEWrH/yIjj3RJBJz7c1sQJCsnyIprcaWLWjCmzxMYvQJ
rU60/N5ESzE0VTiYwBwhw5sWxI/EUm8fMd73giuCTo9I1M0gUGEq23pFDqaQDDpo
orYxPkCmzWPpTj1+sjd9QN5sh/++YPMs0unU9SVG5FuElIPXRxKgAMxu+Uek9kbS
em7GpSLp8FmmZ+KBCMvVLjFCSuj1yhH9v7mFf2MH/dlcgMFaUZqyl61QwpmWff7V
S3IIars9Lh8nLdGg0X1VJO3KsvEoPNY3nvUVmglupEshpxNijpfmyFS2GbcbC96i
l++g1DaL2RjoEBjN7eQQZrWBM0wkvIMjsOWXtl1ktWX0TGMR2sIcahKc5OeNNqlS
nAzakGdls8QI3Y5MGATx1xMSKLR+1Tm0w4+Ac+SN49udFFnN95tLjk3mUlQrrlyj
ehWlwAQ0iWWXg2MXEAJ5+Z0dz/fUAchZxs3nQY79uiNnmGdKR+++yrwAksHfIBZn
Z/0AEsUByntvSBQQpIJdxxz4Hiv3fK0RXa36yNJMVNY8dSgqDK9SI8IFKxAKLIpR
0hsXkQkTxT4/UIOUJnPlXdYg9u6WvMV44mqLiZJN3jaHAd/1mnWfXRd1zaYPaD78
Ys017BeYicDVdHk7uNIYs1DjU6sUGaCyzLlNJ9xu/LcWKijCkOlpwx8QgAGOZV3q
tnOxt+ccQ/lkxSE956DC9Ad1FF20jk+rM/RHVLQ8GeAJ3gB5f+nyO4hlPRIeWXMQ
XHEfVGJsiEalHaZI/9qQAsuR9s/O8mEdPCgo4ax8q6Q3XmxFNIYvaCPbMAtv/Gg1
yoW3pPqYP9GgkAzCefSeXDtt+BmOOJ6wVRN1yxLQn6hN2yGieptBMKuSHRorJR4+
TQc/sF3BY/4mWdVxYoKjzKDd4+4/uXR5LvYyX5RpBxCyipZp2vEiCmQEz+zj+nDq
acVSaAcwsln0mcAKhyUBg5WwvJSOe+T6CsxleRHe/pZh/py2Dktm64IJKKP8Zy/6
OqwEz+BUhG3oxaUW081fTpzGkzCiiLQpkK6C0Mp5sNoSV+0BhtHQX7VJw+zZKGlx
MO3IpKXSCc9T5VCBEptGm4U1BEn0I57J83qk6p4z8J6Er8P3qTzACrQOBiWYuO79
MbV240Jgj5foZfur3IX11lP8oX5nD9xEzRkULEwQ+9DX1n7Lx/mXeD3uq4EvA43E
TDBCc3aNiB2Dy9307t1fnBOz11VbPTZ30OpLg93vU+0byayLJ4C9Uv80c+4r4UP4
71ANohcm4sCE5fDeUJfIfHfYJA7bQhI7nCsI9TfHvbOQg1nfxzOS9wJMBG37vI8s
/LdoqQhMP60QyD7ltO7NO3blpj4zfE+Q/OsQ/hq5vwc5fSVwjjCIgpxlaSPNoEj3
rFsax09NZTjrOQAQ+gzs6CdZJLqGwFO0eNr2IPdusjF07tWpBeB7ejF/GUptlpgR
CWpUkwz0H4sGP+rFTWdqhLdYmz7+Yta1Cbitl6ra2djzZE5A2YbiLU0gJqwav0Oc
jxVCHiEFlMn5JFRmaRqWpyrCqXxGpvlJhD5AT8Ib/RNyohL1aPKSqHWo/jLfRvOQ
q6o9EULFL16mDG0WngtQyrItJWMogFqIMpmHgTJjdVZgVIaKDFSn1ov/3CafPaMO
33wuEAPeJc2+fDZv9r+8tY5eGG2GcP/y6gMUeBYLHG6qwu4ZzkHcVtBVRbNdK0uE
KBiXXy5bHNKRI1tmtlmXM5Yt6wxxMrolGa+XFBVR3ft2coA4ekEIOTp/N9CJxUK7
oYcg56u+fpae9HgClC/S+9RNKF8nv05rcMo1GJbURQGiQSyDa/HYypXZHjtfmkIZ
UyvmqWLBQEBNivfd0bfZE6iYGKFbTskFbX108+CTxPsKEOd3382TfcAnCx7YIyjI
eHIhg/UzJHfQREsIDy+Lw4IMBzyHi7mhckZ1bFAK0Ls0ASliQBFom84//CXR07sK
BPw/H7yKiDrLpkAcycYA1+LOb3PPsXyg2lcOnUg8T3EF8C+6eJr3iGwjsBppLogO
ZLFraLGVPE1EFMfGHuV/nAPzbp2Q9bw7dln13XK9kto+k5PIKQohYsDSp7IQEPAu
cegamlu5P3zsNAsVW36DqL2pl3r70n46jRaMmL1utOyI28AcEGsOCQFFQg3lQ/ux
WXT5Ttxf0uW8yYatqYMdQCiO2OxioXe4pRW7fltdzvUQi4rsMyr8juS8dYAP7G/8
6W6XsRVSP7q24Ch6Z+bXTNTRRgRVIw1EYvAeLcAvUGe1tJxpR6a8frZlRtzhV1xz
nwFcXuMquvmdCwxpiEuAcnUYsF7S6rndv4AmnhiJDRXxOUrMmN/5AmovBsiVxrjS
Bx+6gtN7FTjxUZ/NrHa9JWX2KNigiCtTqgxI0Zymp9lxu8UwbNGc0bptkEXBR/nu
c2PPS3HpjJzXaTUAil3JZkZtMVA2/BkYjBFx3Ci17ylnkcXjic/WxHmchhSAfyfQ
dZT20r/RE9j7qhq29kXZMpQCvTTM0NjLBkAMwPorllqGE9oaUNzOURJIddX7XajR
pCjzP/vf46FZjPtqidmr62NhsAWatFc04f4hXn0t/YXVIIOSl8xVQ8jMitnaYu7+
/XftqxT+nlE8wHhxew6dqi5idqgGmLxtCUF2evrXyECDWFg/wv0oq5sdcbaW59c9
sr6C2eODeC0iYi8pJbjM+OAcYYIOlnz/87GQnUL+Au9IkHdRFdNAuFXUpm3OUZSc
USp/44XbSppDiq7HqvyOyXUrkzEJ5BmEFNi6rawfzAUBbeDOhPpYiVEXbANfUCAn
sMgCNbc55aH5obXh8ndgg4uYBuaK67ZacHFPKGJ4J6A8kRKltO+aabpwzOlr4yR4
eoV1gcq/4WLx3hoNBQeqfan96TXWrf5PDxMI+/Y4qBlEABa9AgCxX8DVzsIhvQ8l
YdW9wlHmm0hd5l+dnTIknVFqXhQOeyHqBpKT5kGsJ39NKwVCcpD1/xxf86sdgWGd
ghjgMywgSoFZdubrr0hLmx133Y9rNk/G1EqiQ+KinNSQL2bItUMWm3dItozmjXMw
iqXxxkWreEYBJJmQLNl1ON1AL4nqHuotNIb/xBtaSZPuUow97ToBjCcTEofcP8Jx
tIU/8mMaJE3HaAuNL0wBS0BggV37IslXhjG2/TnmCoYqlHLlydjvey8Sc5gau3Oc
91NEBSH0l0AmU6UjbvVb+vw3Z+ieob8EYIMIhVUnv3d6WjLpwetYMg0VldoRw9bw
R0aUUUWnCbr+aBjR2fsCiWvJGoKG6NN8fJxTezHyiYvGMadvOQ19sTULGdADD/Mj
/r18RgTdTPval2ma+YKHPsUUCboHoesFOFL/b/J9NaM2tL0ZK3V4wAbur39sMcgZ
vIfUU1r0MhAOHadIbEe9j5KmtPpKzw0xMk5HO2HSfWGWO2UMvpTsmHFUx+lRgVmv
to44ZXN6EoCiidJbi6eudtLcgxtf+OjjZhDApZ/P3DHhgcXC9qmIyEgveYSBuxDQ
456TSoBbnrOSvumCFhWbQnfROFq3Tq4eyHug0MaIYH0NaMnvWKx4E/4Bz+iYn0ym
A8Vo7KxnuhJOSjEWfcLL2FvfdmzdX+NzzsB0/E8tKLXvrzvuyKYdclYse7ATTKbf
VzVmW3d1HyJX6990dpvP4MA/jr+4+dNMfENom699LDOfKcRxn3kEWKAzvkE5XHdu
z/T7IANdAZ0T17ORgfbg3d2CzO6bxXH1aMmFckmOrcRHw2ZmEMDrjFwf6abLpN1k
xIOEw9cz5o2jIoyWLAYPsnIr039Lj3Gh8EOk2CeVTF0m762+18z7q6cQPrJ8SoKA
8moUIQBSLVgTI/X6wag61dINfckbLu3UbqJXAE/DtKZaNYooOhXTBbt3Fei1RZbx
c6qa8jy2oSUSEKlgR72rNsv/YcsQv/HLgP0WuEGyxUNFi4alYA4gKGSfsj6Pomlj
ysHZegQk/UY4yfQy7JuIK0UKMbRwY1q/sBKjlIwReQRMAg9B7Fgkzwn09T5L5ebA
mtMmx95rrGCuZ2uBkvgBXckxhJZNktzimcqfUULWtJMztfxTIZSh2+hnhPMI+mzd
UWnsFYDerP063ZphjWOWNjUBKibfFFmR+fe5CuKBqUGsnqyHdhZWJ3KeK0z47oOi
pE3lwW8q5gLoQIp2T4XgAoOSd/tQZeVKI1N5t91KFMtNyg8KT1VA1juV2+56H+I7
+9MS/3rBQ4jcS98jKFgsktDun49LMo5BOI9McpF4qKZ9jaGy0gL883qoayOR2Z2G
exUuISLExkDxcBJhEpPj4kA1ymTKKr0Vp63oT9PLP/fFfCIrsnhfUXdLaeUfSmJI
K0oK/UqL3QdeQVy9LsawLzqfJAgJKNnlVgwqqMJT/hvPaZqPQ2qfPM1fiYi0wBEb
zRbTyWfOn/9CgMTCQd2Ff4fLrZqxUZljiSqeeiNIvaqkvXPKgk1lH4EKj4jwzgl5
t+/KP0SEWF+BXVntsSlnURlizJWDua5Ege4HdlYgttcffEQgtG38x/2FwM/z+OKi
Cbath11KQ7kQXgpgP5NWMb9Zazl5p78uIQ3cXxi9jcIzf/c+zCIBAc/S+Zh1UcRN
5IG1mI2D+oVX/A96nFqf3K4JfIXaFjLnpuLV5QBknXD+FfpDfkyO5fKG435k7A5P
k7cXNNVdppuZC6tli+X2lRU6DOxsrP0cFrwaiWwTeWVIXpRiViSBVjoSDKu9rkM+
azrlq8N8RpNK4gpqwnUy4+NuenTYJtPQn4qKd1fQDPPdQnWHdP71TMm4QPskuPGI
w3D9qDX9P/LaXXCEJnGEEiFHGlfN85v4Cq0NeBa/bpakp4QFmNOYyI/g89KnGp8w
vEF8PdcNZmIMn5eibvdsIUvluxRZaJP+e0OqwrhggDPgF7NhgXPb12fqV8DgunW6
vHxvLSnf++9POCOeDWiqS+cKPF3yWfH9pQVeB07LLZnFkxu3J8dx2gzqZvByxxqT
1W/ExfqCcGTk5n2W6E3KG3jyDYYqT5xtLBwTdF3TwIw23CKTnlPt79NragyeKZ+X
ysDJbPP+sY1lqCua1Y7b58A3VIgoIx5D2axDUNNrgS6PN97bQ/qb1/LaL5Xzm5O6
XRcJmIbI7IVJyAJ2UctsS9x7SH/BfxQ47S1V12qjngQJgBvmDBd+5SAAvjxXNiTD
0cSrjl/IA/D7XQ14+MebpFze7BH0XfRjZ3uhx/2jPzp4HRIaATKsrV+jT6zc/Sgu
ISdPYm7Rz14FooGpuDAHq8Yjahe77v2AmX6Tk8aIcR7JatyRrhacm/uJsh6ClUgi
/sAUnszuxe0M5Xt++odXwCdvQeb+TzpNmEgAdrjrvk05HndoAPjegFUGuIu+WM5n
RRU+bqV/zX1LvRhMdrc8vcPQCs7djnWJk1GeOYWuVY/WW8SqCgoGDpSgsgxsUaco
COG00ZhPhzCZlpnrDyaxBZApOLaN//CV0zcg/0LAnlYtVIECy2d5nR3lAZT3oeIv
2LhW2TNxM207iWZt/RfiPowRRJmfVdr3Y/Z9kvqxk7o45lwvjBSmbQLtr2e0sDW7
HRoyI/7dlNS06edXCWWs+o24F7UvICOpZMYjJt23kJbvgMrG5JVmsAQLWecIcL8A
B2DQnyb9cFga+LntfmlKFoCaj2Oxqcq19V/4PMvOiQvyFbkE5XBXT/ii5XjRHvde
6RLPYP3C1Ajv2VBAUG2Qe/P7QMMimHDU4gWc5Jsrv7Z7ZNdQ8sxkSZxOc2keafds
p6M3Vb/0hdU8T1bOHc2DnG4VX+N+aoCgohTWi9mi/+q84JA9NRnISy7LikPj8fnp
5kP4CrShj75KsHbtR+lbHW+gpAUR3iVfZf+7xihVYnAApbrTVCsNxFNjK5aoDdlX
JE9N6KKJW68BayO3lnKE+t+u3tE7NvliD+3Tn90rjDtouPoECpifH8EsIrTC0KM9
k/Wc7ukBnXoR1Z7w1p1IQ+eDHyXNPWILHmKL0WZBdFPbX+bgwvSMjMoP00nUxI9L
pks0Daczoe+Ehj050vhS4dKsDrqiX0gqDW96hFmIuHwHsS4n2qPXFTTQl5KwqFaI
iFHQqhzJhrXy+S8zARoX+VIOruCaDhyqoc0vaIOilacLBIwAmX+FpNI/RlB2PMRI
jBhlSbxQmKy3/dfFGwEKPfFmjCVistcAt5qlDjX00+bSvO3Y3uevEHx0IhXflQGS
PdN5W1VviiZBO8JLA7halA91TPPbePI9q8KHdKgTFZAUvdwE6u6IttsSv7QDSgAM
fbwBanJeA0vVfiaLsGCl/y6Iygw4q83+sBHDa7+DxctaIthK9YN7Apbj6CDE6P3r
m2YC2AQn6TyGuxA0mi+GosY1bB0AtuUFeud7X5Av4C+QIfvqX76MA0nNc494QEqh
DFhsw6eItnAzhseiiO4OsmvRb9AB335XwRqDp0QW/z+g9HdvhYCJsfIN09mW/qi4
Hs4u+nxmM1wIhICQGYXJvtRLGZez0LhyuNkaxZAjfAtOFUM7HQ+bUivk3lwa3mNx
O2+USfoVeOopg/JhtDHRp/Ci6QYAIzyNCIY81pngQUYIUd8eHYk/azRCW4gvgzYz
bQo/y/wr+OBKk9MTA+IDVNnkaiZTYTMFbA403W/4nTFKqjbbb9txJnAO2F76vGMS
tkFSGCgPyrpRovQInpJrNrJ+5GnMcOgkHXcMskcu7uAtEp3r2EtSXhm/7Kt1LYz/
hBMgfXw/EXyGTzxk4E4CvoUH0jtQaTFLMW0Fy4VkdEtcVTYjG1reT3dl68bojyDX
dUw1U5BNunjmZ76dHtjxMwJUF+XpOSOdWV/c4Xq3ETfHuZa13tdg6O1J309lYzAg
yMBSm/gffryUffP0QDsdXv7zvb6Lfo8JZ5rfghPpM+5EaYLY4NyZFdmUepN42yS/
/Kh1hiDS3J0NqltbuvwFboqkj9ljxREAESYLjhCxyhfQ+FR1p7Kaxjn7pMvChN04
x/KS5oN2BAnJQkhAyoKMhpLanZkn1f/q9rKDx78053WSZQ6tQPEYvn9K5MY1YCPb
QeGXSqahvkI2ZopcArFyjgea4cY7crk0IuGxpAjlOqyDjzHmoh0q4m9j8aEUWE7q
8zXrpbfEzKxF/nA+7sptrJT37L/XQWP3yeKMIVUC8dV1tMpNJiv4ExZ7uwTala2X
ZwRyzcThuTflJdWI4PMQype/ysq9D98IJjpguaw2jRrW7fWd/G62rbVIKrI3yNzt
GzDvjfYrkmZEuWMGQqrdDvS4SZtcnNutA1DYO+uuuj0QxdV9OI7v5Y/FRcgYt7Wv
7J7wvi8TnTD1yAxQOBfdbYJgguqn6Q0zPjaZr3JStSSmM/+ddIuUTj7GAjXEBV3I
K1qpY22pct9WzQ8M4a1ZuoY0ncKxq2XaByEU9cmSXWYIhuB9YJetwtbeWwzVXf20
JvNGd1EMZV5Nve+occUxtJh4Xh8bms8LkELQjQ5sTF5nDx8S5uy4yQIZlADEujU+
CacKPsLecksZb0rwE6wNWOO6hsPif9x8CeoXWckrOqcMX7cx8JDOaBv1wnnaaR8D
cEZl6zDXF+cdgqQb2yEgYR9pzvrvgNUkajfOLVjD4RMrvscBH9ZNizIUeoCzH9f3
qHem2zWGKm7yFlopOEQFmsZsKeaYUPAIIdcHuNCos30Iar4SjEjQdo2iRTRAl33q
vUe35cHReS0/+rybaQ6UFGqbabbAe95eq5XcEmyq6zsuRqvTpty2jVTKog9m2BwN
R9oCBa+6bfym1iXkeWA3CGqaIf9Snk5hFYb/cJ6Q1JCEAhUNYR6Ia/qognIAKp40
6QBPB/Z6ekF5delS5Ds7SXKqAKPooP5M8+eXCH5ZoUuVFRHxZwItut2VPknz+nza
WG2ZPD8QxO4YTUyI+Z7eG0FcthI36cs3GKlvsRzXOpy4TRVhr/BCk4GgQxReUa8H
UoP+hsmHJRdbxff9jP67oiNZSiofA39aEDarGsbD+LKJzriCm+WkZcze+ZltE+8M
/gwh6z59XZMGrKvXIkZvzsS+qypDbJEvUXkmmzNUoFf7Nh+ysbSOyCR3a0ooV/NK
BvVbJloyQIjnX9EfhPQsonLZx3hBKIKEuIy3BylE5ryeRBnH5Qwz6+mcAzqTNYvb
moasNJWS1lrQyRlDlK9wDlbOn93wXlaMPzDMEtM4P1DNA6PEmeTp6r4cgoDzaP6r
gogrjqPLHgAb2UhyWFSP5aaABAaKvNS0YZzhLV6e4q09wVSv8vinVEFwA0/45Lx1
n7mrSP4gUbn+QtH+f/GEeiND79ON3dI6wvYhd43yKYiKM0TPOZeZO7AnBWaqvuLg
VbvY52fNBiSjjOVCHl5owOpN0oXbhb27aaoKzesIb+HlH4GcHSvIieHbjDq1PINH
rHIvIbHqLO3WOI2NChXBi6HECUXx+BlDDpjAvrRU4DcDdzVjL/P3UIU72BapHO2H
nHofsNy1hhMuoyn73sYEzwxMJNxS7QDAQ0vdBaDJa+B3ymH6Llk+OXEeSpSCRWBx
cC/BYpBopEyUKuxI6UoCxbMYCIIDlkpq97sfHXmhMuOG+OB9uPa2HeYCDi6QRVWt
mcBeTDYkmwtz8SDy6Ntc/4LNDnghXHvjLe58/wk9xWky/1CqiBB8pU+zaZxG9qSa
viIKZQmWF6Bmfx5UtEJ5eINEQBFjcvK9E3BDXjapZv8h2WcLQWiylju+QTGgdIoR
QTscMLv7m1PtSxDq8Ysoz8g/RDO5H7aPMxiSGPKJwxJlIO7gDtJTJJT+ys6gEWcD
FsymA/7esPTZHJ3GPDmF9sDKVNiyw5KGy3cZ6thZaGPejE/A8HWKB+sn1qKhvkqa
tr6TRxdqFA5l9EmvLohjxXhhHMuO5RJ1uro/NE5Cf4LunBeppqx4yAW4x1HkWRa+
IZ1RSUjUOvP0fowQQNeLu+wuKpIPGqqL+OF/QSppDA/SOFYZPYGCnILe7prIpDww
qZUtoKUA9HOGve0BwaczMnzlvVvDeiQG81ZXvN6XqNPy2OwLNmiNF2OcP+dmOXIk
SDhYrwFK7buPnS+ord4q5tMja7n7jczup+UzFljPb+ma7rYJY8qfyyM6CkAZ2OHv
8yKj82cjWpzzRi55I3u8TPQEeiroQW6GfH9NSsk90QKfY1hy2QNHC5UXLEiE0G0G
7rQgUce4ajLEdXd8nVxzCvEWdzf0rLVTlKmze77w0YxJ4eifK9vv3PeAqt7RJYeq
9KRAWqMat1P+ZbsXr+TyftQdLwWF3aawOXq6vVzNOgbaJiFgeRQZBhLgC8GzKpyO
mOQrFPQgOmk7FwkKa15/35qPymBEhramBj18H5Xe/r9K/0Mq0gtT5AbqH4l+91Ja
T8+GjjTK3PDZRHt7DpiAC9Xvd9PBWQgMbr+ox+t+YldUpwBKSd5SWCDhK5vzKMtt
C+lzdvg7ewd6EmAhbjfZy8qB4y2l6iC5G5nc2U6uyiAfRdlu31KRSTwdaRzeFdNO
aXqo8NQHRmmugMHaEuj2lad+K8fh4Jmd+BjcqEOckSyRvtTxDVdOCHr5PGKsE4Xz
Mf2pZU3FZJgfdtUUluhXzccN7gPUvmr8CcwDCgnG97Msb1Gitf+Ko5Aj/obWc+L5
gKgKNT3q4d5A0JAtosXntDyNvIQGqqnAQiph1HCfwv7QQIRduKe3zVlg3ZekpTlS
uOaWuc9Tlleo7aKOz7Hc3FvOLylDVT/Zr15C0BL2I/47wPwcnxtQPn72hst5tE5W
icBt71ng9gSp4qWFmnbQLcM70s28GOjHmhGpAvXwpeRB5ITkXhgT6wLX6UjgDeOS
txlX2PGUJV0nNkkYq98X5MSTE4euC2HuQVhqx+iLIa2z/JOJOFvHih8ocdaNQhpD
FxLeWEXOYzlBAEyrSGWOgyYogKsuR+bVbqsNX3oXfJno9AIH6/jQhy1vjW2bjVH5
YwkH2/JvfwubcjRJ1dyMpa7mBPkkM3NLkvVtfwL5YwOYmk8oPm7Djx0jGwV0v6sG
c0I/nuAyskcYlfcMbMeIf7cCp8nCxrC7fIO7J1MYWRaPxGNK/JLZAHRbq286+XhK
d25Z2w3zhStn6zAhm5XzkA8qLB1vxyBn5T3lbqHPI/GEJsx7PhZs2TYrGqYDjJN5
Zco8Y0sK76NitmdXFgj0iLpGCythDq3rv46JTF7OumSBfj5RctMsnP5W+wjRWNdn
VRugs4MkXXR5gHz+iF8MYRA52DmBGvyn48VsNdf3AEqFi8aQx7MYi4k+HIJ84v63
kScfTqAn7tpS5ZOKHZfIoT/BFlHRWtmNj5DSjd+eyLLG1Qwrq9Pejv939dOc9uH6
aY4UaoWkFFIqwWRSCHelOflLsTFxLLL4oQjg3FTdY3/VGNpCOHv+yqTCSflLfUHa
UYlzslkQpTS/V8Funiu5B5ErobinDFWLQMKRrIxCLuiddgh1W72h6tQVPapDFFgB
And17LaiOnaBeV7EzHUpzyb8zLTvUdD4+MgDXrOXgPXMD0KtFd45hz/EN2nauM5p
6/5rylSNGWHzNFj9NRNnldCnXJ5CmmRYa0WB99zyAJFrDd7NeqpqxJyUVhkPEPK8
lsCaKDx7eWonu0tAUNWpgGdwF7kVCmvc+BC+VO8XZL7dXqALkUgHueqFiuVK1X9H
F0aPsD1iI8j6UCOlJx+QejFRyS5qCse+LO2066j1AvQVtDC1EZK4byD8mtG3K8qb
aLncBVzC3aTg4RVkiltATdytlV0+H8v/vbXdZVxoGz2kYEzXOUbkyk7izRI84O5t
8NDSGZCyoyjERZSWWSTCLk00MRrUKYji+mp7CQLYIEYNOCYHhMywojryJuOxD7LV
MsoqwhbOdk0guCzVcQR3m1c9ddHJGLg2IJvQHz/FA05fSHuoEulAiGPBN+QrfcZ0
FuOSdY8Vzk1V6aagyfGMt/qNOI6OcckqbcotTpclmH20/mejVHQRGb0Bhs4ndrGv
+LEBP9sGkM2wiI58G2ZzLHg3UPjfpNmUup2qUBMrgD+U48hJoqIec1TYuMzN6JRE
BF206r3zVdQxSXAoeGmWbbXHvYeF0CKTm9vNUZTDieFGAVrIUzz7OWGBidbi47OY
FNcZxD0ob8f5LJ1oHN6zLkyvWv5KOM968MSOKeeB+4y0UNT3IARslmtZ4cH304gU
mAd3GmhEIkzG7BxvZO/Hemfs8PosPA2Uu6Rd0MuId1AOaGX9HbWBG+Ns1s4EoUE8
5aPHgcR49HEO5RDRdy97fVP3WcbqxGXYeKoKJJCcNTYs3V1gKBQydTChTNusbYo0
vMzL3AKQq9wNpXfJI21zkmIyStbXuINbbWmfXtyd60j/Lgp+6UtgHps5B87XOotv
jQXDlLxgnYxSQu0AvfpFUT0/o94eW0wiMA7JDZ0A2ADKl3qWrf+J1HKD9bg4L7iW
vbRKJAZ5Q9YG0JW+RZePsfOwbVJnSKFpau8IH5Wu4o+G2T5D2pY/zPC8eWkRimR4
n/u8IrEEJt6XUN+7yZsJ70n0bgWYTCqxK5gM8Utlr9YYhnDFbl3IGrtm7ssblfZj
/kV4QHIMPdKHRHWCP0QxD2K3dl6PF/Eupcz9fZdCXSGDeNLfUyB39gdslUixREI1
DgmMy976fTy6ZQTCWT+FpSYABGxWUHJPs6KHd9uNajWPqhSsuFpMm0V3oGC76zeL
y0jQL6x916d4F3RxfxSk54dPoKNekDTMB/atkZ7/iLNV6BXLXFWRZHnc9VOsEr55
jme0QJ0JtCGXYIR/Bmc9/uO3MD4VHVqSNh62VqHjm6PWeGytdwIAmhvsZS7iNFLG
esi1pRg0CAdUuXAMGB4ulc/IHM02ydSJajbOPZp9rJECm8dZBIXElTgWsjX4IVxM
dp9sAaem3ws4eaLbnDVjkWTIJumtTBacAHV/Iq1XVk/Vxp+IbXNKhM9qrstZzi0n
9LIeX9G+c8HcqISVK4sfGlC7RrD8dguemRWFUFjX6ZrZcJNvVWg0mWA8GoUyA9zy
v42u+aizQ5RDabUcuGGKL6Msz3lnORSWneSBVG71ycw43zRfJvJ8NKFTq7yXfkrC
BvDs2RMTs7shKIVUhlm1l3WPs7KLL9zZ/Go0uAxOwYPRfMArOQKkFR2isMONbmL7
wOs8ofkR4CclBDjWW3upUdjbAU85Qdx0xd5W7riwiUF4e/d5f6WcX5kOMeku8R3b
2dy5uceR6EIAuWuEUvRxPnOPj6Rm/O73hAWL2Y/JrE7jsZG8DN+eEovJzfi/zXek
N2vRml1tPvR8LK1xui3DItvEp14M+6Tk2YZqIg079B73lHInw/IPlx/YLHH5tusO
eHjlgT8Fb7QrXRyhY5CdoYu4i62Rpn4KcpAj4uDI7q773yrQJQw6EytjiHYDsybJ
+soLwAUnY4ArV+4e0FuP9O+peaBFcXnmUjHQ1agvEIR+u9EDoQJwqQM4k9uiI2+F
YLFbmNUKcjhCOKz06QRt/6KjXIja8dSFNmh+AmzTRZT+IiGOhpCXi5p8tw5xTUuy
rmOS/xATKsZtPqhL3YyyhMAESefMREbGh8n/cxn8FyOsi6JvDHkrmP0IwwfDADxb
Uo9/yJSYRDIihG6dyLl7n8iBLh2xsa/MtdphLf+myiVKHgxGr51Eu3agGjS4X3X4
VqItuJ76Vk4+qHjwFL2LqFUuWYMiodNhpeleCwoDCcGIC3ZLcbN9roF8wUCqkfbl
p9eXdFvy0RrH7Vpetv2ZYkI+rdSz1UYSILW5jHgCwcv+yPrB1YDHP919pv0ud1Fn
u3tCW3Q2d3oxYOG6JsEBKBAg5dupE9r/cVUMSkf/r2HuYi7QFKoEMWXQ4DAoyryH
DS6pf3JKdgyP+6WSaRVnh3PaLAdGwOlR4/m1oCTQCAeEZ9pr9z9If2luhMzax0yn
sURl6MGW4mq3kIZ9f4R7ZOdNFdYqANaNXKyQnYbSTdmEZDgbsYstY4/PYC27wVTZ
VGA0VpFnxwp3meMsefdPkKCJr8sDenPvqLwuNaaqibh64qxbHPhUoZYw1Xtc8Rfo
Z7x6Kft7ViYNjkUuPOqHMHOArC3pgGUQgyD+3t3A98HXE+9r1Fj+OMtm5S4SKb6+
WGUwrP7ZXagilwmOciDUa0urFzOMe5fp+9uCSZ/1t1jzmUlXKQtnr89Wm1x9V3hC
WLofIweQwpoxrgqo5lFWTB/rljClMxddOLJQgrLi93bnsam2L050toOTrTgiszHc
O7GjVD1G7S2VXCouiB3gEBwQ1xAM9jVjtcQp8vKR4AeZFjPwzF58nNwTHtc6PZZ7
alts5F+wc5XAAXxh4f7awqkpNW8V0tmjhRu4yOm9bio2yrliKAwfZ8lOLvCtvcfx
LxYNWeHFiP5U6QDPIDo/gUFWFaiXkQTKDGw4GLaNSJMAm5q9Suzap2mpuJZvtHip
IyKt2hPYmTEisQ0ubEJJZK7rBXCEwuRT/PD4RlKPW/l7idsVOcBK7ds17KBOjuuF
xfFCbAcNFqSlIm3RZfAFhv38rco2T80huwkevtIy4XfhY8W8RYtWMxlNQE0vsHmX
ZYfysSWis5y2sVh+mMRcrtS/kp9HtgCE5moZx2iheLPgXNCmWGkc0cvOtbnIc8WH
HjHW3ejnthOoTQ+kXJw3HsnMyXHZEBFkFd7R/8uWlp7ezLE27j9YzGUlM5EMAQK+
mV12U5nMbzS/WW4KxDH9dW8FA3KlT4Iwiw+lVoAyJkfxvPoBXmiiKWDZ2TKYh8uA
C3/TZMGzwbqZA9i8t6YQiv9nmQOaCvaWMElPw9WPJuq6Qyp2DCELzup8aKY7+0Ol
8pPZ4Gzzu2fZsGWTvYdR5rjlElOZdop63Q/cprVQou721AYitV6LrUUhxwbjq7Ib
WZqwUbHToQbW9n2DQxCHDMJK1OjjPfSQ+THbkLQepVKp40ko1tw0BifBb+JzrNcd
HiaSP9jyhlXT0DQD7arNg9G6/3suxsirpmEQ6CQ9OUjbAhVc+HVmk9gYYxSRsd2P
hXb/SPaYTbKSmaLWDepvBiyrmm1Be9+32pjizQMzQZWWAa9EoynDXicZgNhkv5P/
hzQidG7JQMKFzwinyVZPG4n8GdulGn1Ihd+PPZccwMD23f9CDG3wj0VISdm0RRUo
pYJbHyyKRvaQ70XQzUe9OKdNZoTQrWuVj5lVa4xT7nhiif5Oux3J207XNTMEguRe
R6rw6PVwB1HlLuwMtrWHi/svslZuiYO4UsYTcqQlZUTiNPZrcFEJ5lRjrPu+Ojfm
lbJGCf2QHR0KlX58NSxQT3NgPGqRt8fswMJvMsT7O86w61CvVkovYbxY3WkLuTAp
WPDZyGCEUqBJcZayheSjGYjo2IrI1rWxJvtj1pI41VG+eNzeter9DyYHgtcjIZtQ
2UE/s04k7fWb2u7M8tNeWBWBjFsuN9f+BBVxduPazw+2iWwoF5z5cJTfM6TfVcUi
3DQOjSrW35bp8BaPQkVgKPKD0h0OAiHdgneF4CGDoxuqaFwYPzr8+bWozEVrZhpa
kaukjt5GJiFHIrcTZ+GiB/CPjex2Rf9QNqp5YiX7ukBQNpccVsHzup1XpMKA8Mpl
bCOUNUNsmCw8sEbpc5Zs3xghrMRMHqdl3nScg9uh9FcKKgYPbRKGq/fglmq6Orp0
t+TEEODsGSkQZruaTUefwLY78/Jogw6f8vlT5HbnrPgEuEy9Pt0oZ6Afx4XKTSzD
j9DhKoUJzN9suWZNULKCjfz1VNyNnPm/qDNLek7qzTksjnxBwTpiZbn2bQ5WV+04
Ds87S6SR3Al/bnFRTkIxETEMZl439sBqhF6nxfQJBrejCXUBZcR7A9rSCq8EAFoF
O2vUtc2gYK9q7ytTYPxVoXdkLWD4L0fhs/vZlOXkdtgMiX6o0A5e6+mBD/ZcVPJ3
56APERqy3f/YY06uEulmbCNVUK7kLiCJIiJSDtRLtAW0GlCJSNYNxlZGwAyr5ybh
y9w3oFkaLnIsH7c0ryVOvglmAwj6HpSX4jkY56CY00MgfezNqvNLrAQ2592Q6jVo
WmaQfYlPYwzacwC20xgi8nWsFrGiKiAn++otdmCCa6THATYoesbG5/wdMz5xig0S
H5miwaSSxzBruLFWmi14e1o03ZtB16HvBAj0dK0p3skJF7+LkabwS+l/8eLWlUym
T0BejjRXC57MhBXChn73SUmSasQgeR/FJEbc8N1G0IyUfdge85HUKJXZ5SB6w6qv
ZihfhBXIYl1IgQPrVKYsoL8irwFdYERl7ZlwN9KRKvpfcnHuqJdtJBRSeOwpMxJe
bJp/qdOP4sIAFWPXKRApDMI2Bf3tZYtdPkAXNvNSV93H8A8DFqJOgONn638AEHxg
UMjc+uZ+m0wt75KTDt3Hhr6L0ru03pqQgNqEOyfOWEmC38L3Gqn2gmuZ1rXkJlTJ
L+nzqgUCDLvWIJdb2Q59rADed3+ywTNmv4vpLtdGuN5OmO8ki9nqBHqNROVZXlOT
mxytsyb1MA6DxoGvvHVOwQ/waWGt3XW8fnxsOtEH9vD5ldLBpUXkWwd7+/X01rtB
pikVDXJcs8dByWXRZ3uiVyyD/yYiPVFq1RJav7SdKV/oTFBRu6x6Fp49+saPkMHq
pQCAL8uW/eA7p8fg4AMMaHOHiGMCX/mcT9HP8ku/JHvARZq7Mjiv3cRkev2I4O2I
iFYMFNPWFa4Cn3vqOyWDTc+TGrC2zO9kQy/qTkh8y4BDxqnwSZJ+1696uiLSXpsQ
EPqjjgTHNWtVHE8K+/ZlUaay4fGHPehtr8oUit2m2IlC8UEYp9rS1Ybsg9ZLgpM2
ifWovcjlxG+54IMkl/R8NMZ22cRFww2lXsG7oUspFpqkcJObVcoQp6JWMO6WFYfQ
MA2eRBCMYz/0usExsMrpoIW4yqzlP+nMnLIlFWqUndhmR1yn+cEqEYbZ/NM7bxQt
zJe67cBoD+pWqRGxUMVyYofXkEdJuf3OnNc06NvlqLx4N4TRK7hJFDiJTzbE774F
WqsF2/42cSA1rnLGQNVERhPiPk7gItvQyVf4s4FanucU25mH0NT5f5QhpfHpF/MN
K5gaq+eAoqoV5ImweFKSLhZVyqjCjZG5aGB2E0UBQ/90MRTVf5bSt0sobxL7WfxI
j7TEVZgFKDELkPjnnTC+nDjEnm3L7H8SEvm0Lf9FKrVt2Wqt6E5A1JWS3Io9y2NR
AHFf9OCmMGQm5AvpNFIIpDBCfQdRFdJLBkqPjIynlcAOXL0ASVMEJTlfUiFQuYDc
2aP0qA0PTtxCeecr5wKjwM5w7rFspiQ9qALPsRBlg2MQYmBW4nv32J3k8hVZ7puA
fBV2xC82kfq4yWg9ed04I1T0h+R+Yy7jna5gU6JHVhuq8hjgTwSm8e9paCE8hdOs
OlEhSQNUJoFbNm/8LiElDVvClaQzyOKLIc1zDiT5TAlvKsTtsPYnLVKz/U6UnBd7
CjQWz8oaJaoJ1szlBI4Plv9xSUB9BkkBBpDmZDdFBZc0/DKAOq+6ruUbeUCAjyKD
WK6uZGYGT9VcIxJ2YKmk/uU4lFLiE25fPOdD851iXOL6up2m6yfkvx2nPa0jEDO5
EppCi6Y/Jk54zIT5R4JqxvWOaILp9VqFPhgynrb2BRCVHuVjFldH0A3t1FxaqPkT
y0uOWvKF3jQQ4HfmErnC/LnFnwV6yMCPpa/VuMXBfWHSls3cr72DnlUhbkbTcV34
nuqADhfhRYDbFRjBpdVXRhyZ2QJL95sgcECD73hfnyVkhQc8FyaqTXtTz0mP9OU/
1sZEQ1vBtZBQkamXCDGSZcpA83XjiuJ7TtMUlayJywUbs7hjnhPKX4QdnKIFIV9d
CfJCgCMTNbcBxYHLMtk04LJVfsFrzDjPywTCK65TdU89XqcfVnPuszgO0YLJD0d+
YZDeCYfpWrqzsp9tsKQqI6aRCV3lCFMXtbnVp1VG10PJpPVekXbyENgdv/IfoWhd
LUQW1y0JHuwhWTzHSZ2CM/0SM9BGLFW0sbJp/7YG6KjCc6oNXXYHnGMZ1RSIRDP0
PRoohcOWi1kiE8PJdkFEecRF0kE448fKDtvoS211pcgmjy1axgqfYXgPlaO0Zs1P
wYnBsL+CIbIQiI7Je3nIvU6uh9F9OHI+4gklfVygv+8WWJqxzzr4biGoJEvpRSza
HF2gnZn/sSu9fWbLCghq2h+X20VDl2jUJYjlI1QMy6IHdGx77df+28tosXnvFO4t
W6ysplLPQod25oZcKT9kdr8D+ghYVHFqqLUbM115mcDoj6KQpnGtbAsUBRmGNZiG
VEpZU47jU1XIX7pCD2cveUNJ3urK/YU0NYNWk/NLD1cqoYP3JIlvVxe3eN1Fu1J+
hMNF7GJTqrWm6NRfeX7ezlEH+XNSCafPWsx/OMtaYTiKSqprkdo7f35tgs0m7KqW
t9f+ql2iAvT+YapYX/wa0JpNGRrxfznak5lx0jLd17OGZrF8Tb3KFx6WdpFsDwMb
5Rep8+qWGxt8IFKJ64/V8QUXtQdsLtr0NxpaKWIeBHXKrqZ6z5Us1BcfNmXbFTH/
fhVBQHdiKiPspdgdRaa/DIR0SBm1oUbYRreXJ2XIHzRTbxb9PhShbv8hGXe0jHs5
ihjtQhlG7nBASu3UShv91kcvuHPIig2aItpVnqQ5boj4BMQfLKO2tyvrB7fYgDTi
cWVyCg0nxPn77kD74WG4uv+m+QIMRjU7YXusv606KZv58bO7nD02EV88OOcENBtn
rAy3bu/rtvbhuALj5a+8L+Q98kv6hsRq+2hPRhbmYEiX49WRWSBxoGH0hNZjd6f3
VaJbi/mKmyTgu0ZuhuNNHlwpJitb4Nojimkql9oCXMIIlYqyHsbYMlTc854elpzd
2TrOM4rkRlbiEpNRH6ZAiAUzig2iwnm9n/rrPt8J119gaybOycYw08XZy1CeBxzD
8UERSCMU+qfgGabkEKzhpngDgb+PbuLm4A8VHKD4nqeuJiFoHW7ydKmFGBP5uor7
37sTr07TWjb+pm5A8CYrdhluUHysdcyvg5DwM56tFroZw8qCIEPAE4XhmVkjUNmx
TleUSR94WjtyiV0u0ipha8rR4Xt+JmNp8O37T7tJxXXBThvoQEOYGy0NmdnraMqe
wa9PgfPAE0rOt7vWggRQPdekXruc0KGOeZ3QFxfaKSv6+1DIyPZtCA09vSLspe3i
GixYmFpudRKNcy6ootmH57ocVvfHewE+jkhh1qGpsjL8S1QdbW0DK20onY8UflkL
5DsM3lqBoueNIv5MD0NqFkM0p5y5f872pusXvi1cEKzEGaDAoY6aDj0RswRjcr9C
icnOTAERqcjB6c21Jkq5Kqr4amlWecG96IRh/NM0J+1W6jGuUjfnqdTbREb5+m6T
soEqSKUCurT4r1E3dbhy2YF8ksH63OYRcslJL8K5pyGXNf4a895aeoVGB4m6dsdj
NXH35NpzB6U02fUdOpSGlJe3BqMtqWa6aLx/OFLgPYD/ZiRRrd3YV0KaB1vyvURm
7PEQ5tZ5sJBgotcbEcVlF35EXuh8aMYFXdrvm58SJWmR2svLbrEpir1O1IOq9TYx
toWOJkivg5uG8TfIjig9+EUYmixzzrSHQOUkTl9ajsUCJsbZzuwtcRGUc2+djyCz
d6+jtHO8fiQmQL1WqZK57vZgoNARlGMWGclrgBOWs3hFnqGhTqEYjUH+kiT3UZUL
e1HQiOLfBTePdNe+VyTHT1KrMZo1fG+D8ZzAs2weQmE2QvuhpMXcV3wDKj/qqqcz
8DBXxqlWvzyVYdACK7GksdzRuuczjNNbJ+ZC0eSpEyQ1tE3f/coMugY0nDkCDyyN
N7o4DBoL6D3gHRwxapemF6HNwk/X7aaJMwab0dT1zSC7IeVHHC1uSWuhzmxRGLC4
kcNz7FwEWyPMR18cliUxniBNP0XbOtVdqnq7HhJDk5k7sYouF/ibOUQ+iwH1Q+Yz
VndV9sesJcLYh4XUYSQ4IVmIwXh51RTIEE4VAW+Nj3kqe30qYJsXgA73z8cEmnhE
erkknh7yuTSE9Gzzg8LNRrtyA/f6v2Yi8QLJ0a16mJ+/Eij04ExTSc8HOQiD9FX/
S/tnKp3STze4FzopmxuDvGf1yXN8IELYqG9Btr2q5DjzK/d8mjSIcKgiQ7J4DqyI
RCu7Cui2ykf7sdeJDembNfLkXNviIE2T/uBU3lDNfPnnJRnjFdACmg8Z7MkCcw4U
QIWm5KlctHcGEnaC7LFx68YfGvtVBzHRCeXSyXdCV1kULevV9IEGg9Nz8wxuHiaq
aCOQ87RVVmlIwga4pnQvG686NdcCgTNM0DeNZl7vN+7ugUtVUY7KFkGFBRKThvUD
EAT5DSMxdVejBDP0iRoDKPcOHGhJtZkxpbwTE+d2GRyuCyHyDTlnlhM3kkxE41L9
i0QRhLw/CWmBmYAhwkP7dMfJuzrgGIGXKx7C7qUmH/8tlaO1k0OwXM3hxUdmt5Oo
pQWtqID3ymnrZRij7lwhe5H57MdSgBpRuMkXM1XIpivEl7C/cCEwuaY3lGY2fXYP
HUox9KPqeryjvuBna0LBvCGa4w3hbtW90THxYp2GflcTJQJzoMOPJBErBW+ijCfg
vBvkXLrV2IXK1ytkSR7DNz14QVg1r4p92HOKBUvVu+g8nDCXTVCpKVG53xNKR34t
ZxHruaO/T5Bn0WqzvfSH2tuDRRTbXy3BKV8fDtxIJa8WMXmOHRilSU2LW7Za+XY2
dYoTqczU+yODPb3WiS+BUnXbEaA9IGZXYWv/UVOUBIfd8vG4ERsTH3Qn0xCyTT4Q
7lUwzS3bAY+bvkkmP5YvsxE9uKDM8M9B6n73KsMOM0ULSf7fvhxfFzAAm+8y3B7L
T8UtCMM7b4x5v8Pap3P8JS7jD+Z6AKk73WYeoA7HLDPeURH3GJoiMpZAssSLouW1
hO8Jqyi/vkcrNuI4FRE4mitnyR1HxXvk2aAieDXA5UFp4WDCdyehki0Bk0BXDrRz
fC44uMRiv0WzYY2wrnUBCXIZ17iHcXZOJf1A9+WZPqMNL2a5JepXfmQCGu+uFRH2
x38qhSZNHu3QzCCVz4B7WtCS3g9M2WNQZLUVM2Atal/bHNXbtrR82agpahD+gP7r
SxLRFnUwdR+LJMSP0tWmocP44lmaOISn19STBKcLcpLCqFi9NcKgxbEQGinBLKDy
IXxPWaPBg7jKMjf+CNhLRFVvvdZUCYy6Q8FO7ky9ZxWUNOTX6G2qVFf56icSjsob
w3vPn3F6+DlIKIWxa9s6+ZK8TFnj3h38z5vAiCllL8Ocn0BChqP+nWBOI1/RN0xA
YU3yAdr2GBLdrJ8vbxHatgqOvj4BlTz7GS+vhtJAuFizJVmtcxqAxIj1s5auzmli
coWb/NnTxH6NRgtmRpIQdinGeflC1wT8v1bXep2a6UMuyd/cJTEGEUryiwuJ4RRo
aCMFyg7WaVB/FftM/qhM17C1mhYeYsBG4IOReTNmGBetxRwY9gmXj2hhspFciRUi
03ns8HPx5DoqZo8pqIs8iV9J0exa1rapAloK1JAQjC5KSQu1pbOzaOY7/hhbxZ+f
T7kzvUKJnAfnFTFbDfU8ulleonaQ/JHuuRSnq5C3IM9yWt5A11Zglhrz/OOlIao6
moJmtzW4JFlM9NZPnwXaip1L87dH5kIRI3qD40vYl5e3A6h/7Yo7Y23u/f+CJ/mI
1etwZE/AO+TedPvThJ+UGoHdAvibtlDgs4+EpnrutVWjhUprzUU6yTGGzsS5Fn5M
mH6x4bzjtK5wwyvncRvVz8tXt8QtW4lfb82TiPgVIrg90+kUJ1pYKqeVcvlS1VNy
m7e+c7uQEXC33tY9PoNzXADT5SL1Ew14mfkSrkHlgfiJDmRvqYAVqxkOWNdIzXQe
TYSkoMjF/FKqse9GbE3eTuxaXjMiA4bTnOgyK1FyRhMy+9TEpNq+LD89hosYnxAq
ObD+wlfrr3qsO9wVCTQM5bo4bp5+lyk/82MzkgcGbzneGjw5R09C7um1FZMGBQzB
FF5KJLqWcYd30iKquNprksK+u/uVb7CWDHFUNRcyFD9VqbbmPzq6d84zeHRkrzNJ
43+ev1kK+BzCe95sm/78k1tFBRGyp4jw/gKk+hqG1dEFyOj4DHrHltnNE6Fwy/Ir
eorn4VsdStIW/xg/vlmKzlH2QXHngCJHgzqxIBydtOPKLbl0MZsTfy4n179dp+VN
fGhwImJV9DKTU54Mewsce5uGRmPIGF13TVfCTb57xZkmgpwYDDyv/N6tvT1ePEKI
x7SkW3u6cUEcF9QZUWEe+vavvnX9VaJWhr1+lzXb21lEPMH07r6rchV6KH6khuEn
1nIkKW7At8EE6ADNaL7Ag7C2XW8eM1XBAgjDA+95Njntc4UH2Dib94nlaBKZWTad
84YEbp0DPNmcK+vKcpgRPiPNemTLOCb6Od23XoMflWGFSCydev/RDa89nPmREJay
8aiQQq2aKZYlKqLGdOT8grZSmu2+5eMdyRVRZ/hz57dBvamfkyhCOWgumFAwY5SO
ZLPnyragXpGeh4vELFnDm08lGwKLFgVX5C1O28AYLXIyhTgXdVhMX2RhF2Tb7uxj
j6x/JlRnGSORcnWEiOMpmlbdRwbhuU54SrEB8Y4Bg5vy7A79xr0vcr8I8IchgXXC
XYG/ft5RGBuOpun7dO8MrYmyJnsLYl6XPXXZ9MqEYa5AEIyOrLy/wecK4VqfhRy0
fLf1i0nD5UeTTxEhTOj06U5dS0TW7ck3+WkRcesPk5ZFlcVKHgRfT0xc4+Q6H2R+
et5UabPRbaAS3fxnCgmOMms4PxeVQXO2z+qh4WnoIVqsOgQPh210rhcezJ8IJroW
5rC2Vdyry2J4bFt0QK50MV4OnnkoOcc7OKWwwedeZfPFbXYlHMASTXPHDEMh63KZ
DPvP/xukgX7o3oxJ4PViJChdTSX8vtRPQcuwpLaQR7lXZJDbDU04FwnwCBXXgqW9
tu2Dh4Bn9eN7XQUbS7cbwWH/P3M6dn0NuF90cNCwAhKwXdzhEaUKg8EA+hOBulAL
/54Pl25yn4dznquJi6ztw55DUMk2Ct85i6OXr+sUXGCMSchgdnrSuBNnJ6GKO8ZZ
w7rEDAo5vUoTgKj4M4tdWDMQll4sHwqL4GCms+xgEoDw7UzP6CWdH5jr/oky/gDK
d8NCMz6i39ozWvSGYwMLvr3LSKNz5ddfoIOIych//DIibKxMm4/gYZKvza90oS2F
vYN0Bpk46+TDZfcyfWpnFVBa68KJG0XTsZFtG55yj/LJEqKVYMunwawHnFaiE7MO
fFPPe4stsRHYLnD3Sl7K4iLMmZ6LDwm+aNIIyTPKobIJDSubPRQJa+O0PL9NS95h
YbloEfB18XBIhNVn99uBMBs9VH6U2ECZKexcxMFcu6TgF7xLcTu5C2gqQkrIvnWn
lPxaofCKhr8ObqJTkUUiepSm5A8cQYBF+0O0JKJjeU1pWvBFfWN2LwVZONqhuhiG
euk44hnthMri/74RdgfUH2VHoK+bAIZrXkroWneyUzW5aXPyk+FifWpTkWq/JnNP
55UDYfUPoH/1EwFraPB9JgHVigvgyMo14UToJQThHwNs4fKwH95j+dsh4rQg8j99
BTnxY76XI4GxPWUf9QMLkxC2Zc6G5z5yfp+X3Chu8EPTAzeFO7sjmNvQHIvLdQDI
fJl8JC1mgfDHo+9X9qpboTD/CegUmnvtfKqGwSYIFrAhMEb4JdC0btEYVGh0qfEw
gtgazFuoAP4Hk+Me+xHWQDNj/hmPc/qOO60Bm29GOl+FdjYItna/0/ToBuGMgYPf
mAe50zZVvGo4RlCsCY+wiDSaZQDN7To7ySby0B/Nf1AOo3/58RP+6RZUo86dVB8X
5+NKq//XTxuuGQtguiyNiRCz5+t/mu7vok92UPfZc046kk7Xd0xmdNPfotk/2FDz
xr7ivCuLBFwO2HDZr6uGwbHFIFDkvtg5vJxIhKv/ViFUy4PbiIJKgM0GPM7g9oDe
Hb/ByqFuKfEf75lz1yw2DZIcrAmL2PJPt9v6RVhct+YRo8pKepBWygTMANhqkaPl
F6twlQ3HR4hofOTO1b+HprLUXNtMVg9IZia98DQbt4/j4GlV3Dao30YklFbKv6oZ
WCci6TNCKSlQwpvY/ERmjMrHChGLcBOP+jUrewmuilDjqBfoYBKaC8hbVncHCnKh
qTPZtXLQimivdyk2rpjoVNIUmf7B5JcRp7nCA5yRDjMCcXShPX/B3QR4NVM8epXt
lVeTZRizYeWPEz4nR0CTeyFp3VYSvSyAwblWXikbDzmbX5fot/RUmspXuNFf6C1l
QiBu8+F8kkcwy/gmI5XxJ2ylLlFdIAE74AaLK/j51q5VsQhVYPfDb7T8hOWicFv7
Rn81i3mxAsTgSbAVAsaIC5QhqB5+gGAhGmXR4ZQWW7toWbKzB2DlgVmZiAkWWvHc
2hg9mM3kq7oxCKeuoXNMif61ozi/TFgWvDQfUaxnwkDXfpzfLJRVItdck17g4o3h
MkKh+CYidx4HrL0rc4vP7MdACaFydo5mmTLwx8ErltGCLD0C/UwbVGRsREOT9NA4
cfY8osu94QqF/Xf6cjbU9IsEFnT+TeIOe6ndIJomOj6b+2CXnAIIgf5+8zeM30L1
4j96p2q/CPd5sqwSBux5BBfoCtuQocBt9J+Yq1mhrGIe26lJZ+pvZQVXOwSgSWqD
EYuXr2LMEL3Hv8cXSQmBMVqe+s9whjHHhpIYbhMnw/H7W4YHcJN8U0zO1TyzePcU
iaKgW7TCRXcSwmXFkqfl1zuT8L/VeZDl5w8xDLynIqKsnJSisfc2pLS1LqWrpVEX
cAqx9LvyepuF0oEgMLZ3EYYu2sYkvFB+USVnib5NzBn6wLQcrhL/Mk2RHbgYzC0A
+XdueVBIuUh+Q+unwzkQvcKdVgIQcAPEDKsDFNYBhrhdTN75B5xnC3KOOJqM8juO
c9OYkqQdPn5gvkrVLoip+Il59IGebOR082mH4HmyLRdDFYtg40Mlh5JR4uejCcJ1
5VE+RbBnUNbp0VIxqZzA4fswBOCAZ9iJ8XipZAu0urAHYJt72nFXHsRybAq5M5G6
GqruOiDT7NtimeC/cZDBFzEa3L1/aGlSqgDH5Qzln3mAtizmf1zeeh95mw18bH8O
v2dpgTAMzRoMcbqBA+RmiewPjJxkuD7NExHvux5/xih6O4iOUhL9An/LftE/zc8N
PpDY4cRPeeXTJwdm2DsCaomik5dI35V5YRJtqzsCY01VwRHmXSm3+NTC8qoFssB/
HO7MN3XOsVlvUixKGHkaOsOCptTQGnWtLWcmm6FA6JgQqSKpI6pgkTgz1rmoDKii
aQGakcsWCrk2e793oTt13VO315TQeau3in8umMGbRWdyj1iAkskFLO12/HfflVdM
2OkKkD3tmTEqXbbdUCi/nMFRJpSWTvNAPnJ+hoPjIXrvgof96Evj4GM3+pydKAmT
EoMz0fHsPVA627w2J/ahuVOrr7J0ff1fTL22Axm3ooCNQS6+iDGHBswaLbI/YZGl
traP5KmqHlzbBLQVNw7gtadxM8vwUCw1L6LYj8Y3YLdbvmu6uzfgBmxD6qrfEcYe
siqqjzEIqW4mNZm7ZTam1hICPo10nyUDaA2lIV3agbxvSdJ+CdysA/e16VJ6+72C
j0EHiVhtifoAsbgCgNu60HX3vabTXAJenb65ht0Z/1Kb1Kt3rbZED4qgioWK2DBj
qWCkUQO0Mm9Em93yRFZdyCqQe4pvJxCrxISNYaYCtEEv8JQkWdK3Z6Pp8y7r5x8n
92sv8eV9Jwjpbs2nQfUgYRAvmtBJaABc8NIjiIQaWqIi1mbpJCGLgmJxrzK2CIj3
FOycDY9vul1TwcSnHFOSAPYI8usdkfyOPauPyAHkfjXRJBAuTlUGMF5aCeWJ/ZHA
L79oMZqbi9oqAmo6rk94oIObTJeOGQYIXNlwMzQuIWzlt4ib0JBBD9O49iaUkPs2
MZ5tc9kIXs8IdHhGLDLJltOzCCmQfeYa7wpW8Q+R8/OpMo3PZs8LbKGYmEfmAvUu
RjE87mGSdLKVvlxPuM2wldV0ECgP07bjgbRUeazRFIcADDmzL7WtKIuqQcJfLz0i
kP1tGhT0GvuNAQsyxKMUNGCQng89GUUZqGU21fy5clfn10uouHGaSs8xzSmwtW5B
6jQghsqnGSpFGTYDBbm1I+BbU4XhDCwfcPiCzE/VFSCjhAY88Fr//BSy6obnPM9X
GAYWcw7sZN1klDuGnMiHN2EQ30ThC4Cp56emj2WLaNxjUKTwVx55l/D1639MjvwO
E+XoiXsihAJsvGcMSvtFMcpZLL2HX3dslIDjsdPd2LaQpGhf2kY6+fuhRtc/Ntgd
s3VtkdnLp6c9ShuvMFP9P56MWyw2i+5w46kLWRVVFNrg0SqNWSNFbKz5iNnUPHEb
YTwpZKN6d0YDyf/u2uoDefR6e4xAOptRPx/+JUxM/ZGVRi7su9/OYlhgrCKIJfbC
BgQ+8SA5xFc8uG0yGZEhmk46YM1Jl12BEQUH2VfvbuZF0XIRFDUrxsOVNX5ft1vp
h+PDuWCkwLomNuKc+Zu7VtLcOUylmok9q0H2mtOxMcv7UzubTkp+kuVLPN90cDAW
K/B5kbZS+nm0UMJ3np8z72ZjUBewLrPnTFkmudPoL7uMg76F1izuPzJuTLYpf3G7
pWqz5zZfmHMY8P1paKqtn337GBfkb5u1K5BnMg4k44GLfC+f7cd/UfFJviwNOiZd
60FSEkuDPkbNJ9jAgsj/dRfrtvIcQAZr2T5KvSB2uiHpFIX+icSlnvU0ydeZ4rtk
H/QTFpOnZnap4xCTxIx7efwaRHS9AIrXded4hyW9qO/RD6E0HkqGcKOfIb80l6J+
jLN0nYrnCyPuYI+KdzYi1cANj9gERYlPZJd/kgHBki7YU2PiMmxwP04roaIu0frP
hz2MjWYYgznDT2zLaMtXubdh/z/S32yoBO7QZC1IRViy3RbP4lvAWUyMl88U64zi
rzSmQLS4mpI6LLZ7YKr4yG05NQPVkrUcrZYvdBcMoov8hHJZXKihVM1+AbWUe0Aa
SCdhEFU5Hw2gStcXBU1iuvYQHIlZUnkjKzz13fEfr05tjppXsGUJCYrcm6yIpuBh
sTaOBEHhhvQKNEkIwDwvbXiogXFIj3aomFAD5HOXNQyoQDOCod5mG+PXF9MLB/E5
zJWKSTkiFh8neI1Z+sNpG/BaLx+DmgecgMcE0TQF06FI8UtlQwsn7Wipy1yqIy5t
00nCwKuz2pGAGFgSgI5feTRlgRHERlRM4ULxMET4202/kPwubQJ3zN5fLmdSk2ed
YkFTDAgLCiq13JHbgl4XpURIDT8kEiTT5keV8EctWE03MSkC5Yi51a35cV3dHwDh
Vd6rMF2iA2tiLRmRVt5ywmSrzMwiSQdQ1eZdIDbky4APW/51lAxZRGxbe/NP8qay
E3Wsgy/wJEgRw39pDIyq0tWrhVk4hXxk0iENY+id/yiCpUkuIEkjOQrVEtu6n2TP
KO86RrD49lafVTITAsdXBNWbyaP+8p1Gpq9Sj3ewz53irVSYnPhe1e9fYEm6QPEc
g0KfqD3TAM01jM0fO8Tao1go9KjbilSdxxWvGYvxjMXyLUEIq4Eix/Vobhph68ag
mtbxO6uhoG0vNPmkVNyizoKjyBWslvPYvvUauu+SXCR7/d/p+NwpN6oVfGtqqdkh
7H8y+6IS8d/Aq6YQ5aI6KDfBko1M3sy2QadIjjEFS4Ry+aR7G+uf4t4hGAVvjohW
n6tezhdoZcpmm8HYtIIfzxfVQH5E0jQCNeBM+zy8fyp1M8Lh4nMTL/iBrG7PF4PD
02dMxYxwZwbzD+ndMtY8ElAOd9BvyOgc9DCJVIdajT6lm3ZwL1dNEqLHgJT+RB9t
6xCHsieYBZMaYGUtfu8M0GL1tsIm21yjTSNRSg6OWxdKj4ynwgcWZUDzTnozcTH9
bCTr5TEY9HflYrTCcqJXp5Gp3R8emULP4t5wErnplrh4+Ra/Bkzh3Npb2s6DuqrO
XUuAgfRwA/K9+qCjc87vI9Kb0kb3jbGZad/whZ4YOyyNrKMJdiMnTWPy5rNMl8Sv
9o70Dj8cDMYhsdlOnx5T4/14mpcMIxVjKqTnw+VRPcFGlC484WR22NpzAf/S3g7U
Ejrc166IwVRqHWT7WpUHqT0PXeEIjMwHZ771C9xT9K41vA8u7hlQiJJq1xLeijF+
bGTGyvuLz6zM5l9RtCXw8JZqLP+mYGpMa63yv8PL14AKI0dllEbS5WaVly0jG7Xr
07xXGzjWXrRnFDY+ijRi3HeyFpPwAwYklnPoPLWsHRxnfX8UQdPN4f3nobES/ivz
Nlay4Pb/B6toBUe0mOKNywSx5qenJLPY7l/s5wCaeQJfh4lpHrePH40A41EY+Q9F
e6mBvh+mbA9qKrSOv0XDezIwFLA/GQGZj8ZKKoByw1VKmt9NuQ/8Pu4SuuSGcAb3
4dIeePpZA8Q2L/xW8znqSvpeAFk9ohCDEaZ/44OQqBEhH1F50WevH6Kw1jAJkC0I
5rBE7xtZmZtv/wp81c0rnZXGp1EqHG+ig70cOJmXQW+rDKiPJ2MgO7nM0Bk1TnFC
9JpNeEcfHEK8eyNbLLZO50wlp7SpKoZYG06EDLf5c7KZIy0/uIqY8WajMXzHjTRG
nZbN9RAKaFn+ag+ZA+X3ZbH5dUTm0TP/zgl1h+fXPNQyA2zXk8b+9VYlA6ZOFC62
CSvv06CbfTKuPytp0pwFegMCWFksJKdVx8BiFwtzI055Fzn0+nz/0Qwl7G/9KOjD
SwKalsN4Tm436Ox6e0bta1C8/H85bnwBMCCjhBnGYkN2DGRDtzbQt1q3dC7H6Vw6
vRjM7BMtpU6cqqLbRGu39uFstaTMOAqGXNF/BMWDtwmGlrCVO6Vn7QxilZALHpJb
yksGXcJkEawAxwvcSrEYxoknNFP/cUq3FhTQgKPdt7AwvEMdj5zcJs2hMF2p+dKh
BygT8/L4EHkYPWCyt++4FC703kiKYNVo61brLmL9HiWDz4jJFEoxv4Y8Kj3Ri49H
OpMBPNLpxL0wg8HBQtVJxkUSMW3+Hc+XEVzy6zXGiAYUsHGSsbYMtNxEipE58YgU
VNQ73TuTJYty7ts6zMG1YxOH60StxOjfuLUwCX341LQsUM2ELdqfxRgD+gasIS0m
o41COHtpgCzcMLmZcht1YeerkkjdkiCRSXzlHTIMCd6I+ihAZ37Oo8FZ+HR/YXry
YtEDtE/IS5X7XhX8PU+aky7MKRitkf8x6hYDDlRfQov3NFXQV2TBozNNRbDfr+S3
6NPfQT5kSUaVFmjcwIYeKkr9j97AJM1ik2FGl3/faKMlH3Vp9DQSdN0VhYibxWCS
279lUraDZESlFPihg/DdLn5GC5htFrcD7xU5eh/oM3k0giv5Ogz2cRt2r0/8+dnK
hfi5yIEoqWRUmU05V4pvmquRbUQxlGRYv7QPNNUWP57xJPiqfrVqYQJkxwzZaBFv
3L4CZRUmHu3zS4YKq1Hw6laKzuU4KIDZLVJlHSKFOUWPnEEZlK0mDOIdJLPLuKXM
8uqIJSkO1NEOnKYAG7pI/MVuObjCOrBcDu7v9B/e4KlGS1ZRsnwGHhsnqiS5aDS0
moqN8X+31frfa0iw2D8lTPjFUxdyiLbu4JkYcAUBOGOPlRH1J3JnHA4zoRd+w1kM
3x/uvdSoxenaI+9ru0/97wD3x5Rl+uRiq/OOYs9lZumE4LXrNSjewiFuh6wspDjL
3No4Anlu49uGWhSUalw6X9udjZKFlFqjW2iOOEysV3+oEZV6Vm0931IFMOlLiVSX
QT4iMy2LMNI8XWS3A7/xq6OMPAIxe6JHuBjrAZdAnyxA7lvMvmxXTmpNpBRaHRXw
nXCuCabtCXZmQUPeZ/UZmKcX0twqwoUjyfa/4JEYJZ5LUmqybxfOJRLII0bH9Iji
nlFF4hCL6l+2SYEYzmfhvr+tH9o3CWb8ZJRjQDQwWMl17mCFsfW48X6/t3qdtA0M
G019pn5qGv/cq87ncVaSE7J9Kzdj2rJpk4XelYujtJRHCSGQ1xRRTpNZxybWiKtl
iRv2Ve7MzFkX6PTD9APH4g1G8XUVTldwRdvRFjMa99JZC4Kx0Zx/udHc6wt1muFZ
2W52A28Wt2ZH0inI6IVdaA/Ns2Gz0hyeXMiNI0736KGQRXVU2gDvgYtt5svg2UCw
lDjRO7pyp/Wkj5IdHjOn+8G/v85kq5xVD1O6offAXST8GI6V2EYFn229LcwR/93R
ozBEvrWFuTR35f4ShGIVoF//wDAmy6KHK0XrM/Qh+yIB8AM2smBi2OhxR83q5eAo
fym8Nlum+DYbyo0lDkf5fi2XFyOXGd5DZ7Ahr+dxDwVRPPgDVbMBc9nVJepTlg4l
smxAI2zM87+R+TKj0JdWohQaPCLZ77xR3/VNhj5lOJSc3JR20PQTCGO9KcLI9FbD
rOqrpjZcSNIG8GwBsgcCN2iwpyTXX7gx/E2DzQnOSZ+KSgihbDgcEr1y4VPr371N
yOTv3tklPcthNfYKxqUYFQHnx07eN2AqHxUxK7lG6HGWDSVHa88UpKQzk1H+duHP
2HWMQqPVpTDPdKLnb527k6pp6OkgDpSlwbf3Uo6kLCTigHO2LSZoZ+7zCE2nvffS
x7QeAOxK0TXBFm2Ygx2MsqQKtYsTtek4cKbsAxWSTIUDqudr8XdtDzwyHRprEQGr
szwZNp7Y4HbCq8QPn9Cx2smMPMqf8vhfXTk+LbUecIDDU4UQoVS6fdAD51+yAgnr
Dpl/AAASA2ITB9ljv6TN9humZtndbBUFwFZ/ukLcbM4Wl0/NMXou3V2jqoKN0odG
y0W2VYk9zXiUszsjnljoFUWxL7/VBwasHxP+Aq38Lenv1NdDV903esof7gNyTxrU
WXr3bTK8cDsA1wb/xLUwaPC2Uuxgl37Sc/+/Em9ETbv6fkOzBBb3QGvlgMtc8CKv
g/z2IitgJzjiP3rGUXTpIBj3Ts/0xI2jwyF8Wr1ngJuqH8TEFXk5RtAl7iFCH1cg
ai9XbQfkPJRJXzZpAGfnqjGNcBnBP/1xLDU+KzHULX0OGo0hyiA6R9qAXrhMdTFE
5QwR4ejdIcAXDdCUY8eQcs8BbBnWJLgom0MWQcUx9XtiPlNYpWeVgOTeeKY7uJva
OCqftmOvcFNL3krM75TGFRTGkJaSHmG4NfauBzL79LbI/VoxlBdPfqxUMIo4aXjE
wXXhCa6vF9DRH0cZHMgvXXhi4S6HeeQMeYA8Tydi5Q+QOu5szSGUIOXCVZn8IGCI
G0zDSTsNSeMgeGmUR+pt8T+KgolAABR5qXL7IeYv5LUOJwXjT9nJOK5SXEHqbDYA
C2aLFh3f3HQaCer6pva/C+Z/Fb5DfP9gcoR7JCKnEgXBHFgirALdOiw/mdTZO0Wh
l2NuSpNjUxktqmsvZdk1ZZzro4mQNbnr18dkTXsyQwha9PmAC+vtg9h5pIILer4E
ovch6rJ61RUNXBVezGiZG9hbYRLqNIo+xF09eEjgxy65h/7Q1s4tJoPINVTPl5A+
n0Mky1Q1Tt8+F5/a6fXgH8a+Jk62YDdTUGEy73kqrCVV4dEVCL7cKIhmGGvneFMu
39S3NQJnlYE931cp+K5yEk3GG326fwjQKvEgzlYgEb81/zqWup+BLUwgKOpuAdkh
M76oQEikWFbo2Oh2BLcOvzY7TL1Dhtb1MexYzNSdnQ6/fTK5pU/tgezWUEqpTzRK
k8zoIIASnz+4MZSjLnSNNtaMvDnWj329+htwzFASRjBWd+u7paw9W+aCveEdKZhk
TP1+T18+bDXQfaYrR7YHl1RF9ouxYfypr/nAO2ylOTcIzFixGyzVS/I90rRKzP0S
7jz7M8C2bBJz5WJw6ziIGwh9ZqxUGc+C88pjQg6FbvqIgaZQGds5VrFzp/arGOfe
GDl+AInkDTlZ1YAI5TXwGpGhNIX/wsTVN1pLa/Ks6pAs79+gIm6bYOj7TQCWoRcU
TZPcDi/s/XYb0AUNRWH1oBb81HT8pVlbNoztC/a871jMYFrIRcE47FXSzL/X8WKu
GqWMzLewCra/3VmWj+3xEXgEOOvYImOYblA1GJzKT4n7jam1SeXaAnN4L0+G0Hf1
GeIGhLmnDmfUAgS4gsCqHdcTeHPZBQ9sBJO4geH7A8eVaesAcwXTWSxi4m2QdVwa
G/GiqPDoyL4Xv6ClXXdhPDY03Qe+mR3QPza+wsA1iO2ymKX+ioxaCsA8CQuQGN7X
aJVe7oYAo+Xar8p3yjta0NZCnb1Vx2vhWLQEvTud18kyhE9iC3cZpWdLGXFZwq0P
/Jr+bOCL8pgYLavZxS5cAo4uFSra7VYf7IV/RnALcRnWdgkUkiIdsj4A8geLC6tv
jwtnWGeqMAF+m51+NlLy9ivs+xinEYZpMbrVQiEt85+a4ZT31YpDEbRBu4OHg74C
teuMJ14sbVOcgdFrj+mG1tJWsDm+0mf7zfyxHHZr3qQ5OIxhvXjN/Apw8ZJnH252
EvBc6+T47n3FBXxECs6Xt6Cmyj/pApdy+1bTVeLYIlNWKd/Zwd67IFQoy4IoeFhd
zpVcFPxlNlkkDgVNX5fUWf1SyqGFm6yBp5jYNW859rrE7NQkRYetYK94RYpj7ORY
vqDKxFzh51SaJQPnER/a9R37su8/4EMgZ4UTZWG63GqK1tcaxrJ5oYX+x2SZcgKD
qq4B2tDYFAV+9XzE7rYsSmV9/7ghq6MxJDzXdfl0Hcf1KOqnQDrNZHbVgoILFmvO
lsieHZO5+VGwRP4ps3dI8BLvu72eCDY788yL1jhjg+WNI6mPTdiWtAz6t5j6jC4o
wI3XnOeH0I1kNIo9Q9KM84s2t/c0pBa4KUeZqGyzrG24OpgnV/+ePyvvLxyZ50xz
xbMUGal11dsvtwy2qKpRd7O7vvTbFlHyT//kcMZ8wkG1ns+mUPpvwUjpRbZmSFbN
vksb5lbaPzhT3xA191qUEFv41msDacQZEY08dwQwlFnJPQCxuywcIHCickRnnmh4
8dVB30mOOAHjKt4KCNC8jjYphUA/Ld4+EOggmwmsWTLHLYd7AG7SAM2capntIItA
a1BnnoLL2S9DfS7C+FI5NhFpgEt6zwIouu977S7MbOlnyrh4b6uDeY5FGJZwH8gE
TupicS7zBnZt+591hd92yQcFGGYvFi2J5a1/U1BO5WizI+urLdSDfTGDwOFDlber
1Vwv+kmtLr6s/pHQC/BJ/YbN/FAcsuZ0/n/O329sMEkVCZ9F1RERieXIvfnDOtA1
kD1dConqDnJiMANEIN84QO8KjiVukXF13HPpLSKpvJcyQrWcP1EjtQ6l/Hmu3icO
fWwDEebIT1eJmlVeqCf9HwtIgnJ8lUcCYn8Nduxj26u3uLo3dH2oN8sHtQwVRQV9
5+cq/CIjikNMhQnNlXRUpg6gCtvI4Xd80zDsqW9cgeDuTYLWvI9+nYYdZHl/lCbC
LAsmHUinbi0wMHKXb6+QUPn7YQJLJh3EXSBBbuTjOBPj1kCCBtGuraBJPURz3fEV
HODSJGVeNvSml8o8WhWpcyI4/5TR887pxxx209uAezeSV1YQmF4x+j4o+t1Gg5U5
kR+2DxsypuO/iPAQYnSL3o3D2Bf+GIaUqjykJv7aEH3x9iwqCwGTZpcC1btusH8W
zFHgpdVePRqo9cAq6vYkj5Xh4cNtJbEHRb1f1rkpyCPFZlSHHZnJzaGfSEgcMpeu
rwZlS016NQMmS8NcW4naR4z0qg+Hgv4kNxiIq45jKBYAabtwRlEjh8n1Nbu3erSC
Hajb2sG6tG9TfVcY5ZmpOnFkVijb6WIHp2GBylhTtpdxe14DYJLZOM0EoZREJEKo
D4gkDkHsWqAagHHmyFEkq492QJrq0FgPSWGiPHPZf/zEBTjoKfcCPOPCBd+oQwNa
plVp9DBlCzM/gPt66NfE4OKYz7SoKnzfZ+oLZa4AKPxmeqngdzR2ot4+lgTkldij
jqfwLSIExdlFjVxF+uhIkTzQFCrUsJ3Hh84uD2Mlljp4I+1AT9V90sRdqwpuc0Ba
YfUT8JuH8CZLnFS25kTKAsnWB9ZYVXNINIZVSRNfHCzM+Dy5ZLUIhjI4Qj429bnh
Ym2Wmrg1fTUlVBqw74DutEdKlkrxpLBP8km4Bq+ItPQ3kP91w4es9ylQBN8xyIqe
k4g6cvwLVtbnmNVbEFPvW/+rLsnLeqsYaStBuCCUqW3A5L+YdS01K0Nre9XqRKVG
b0wB5TkmbewAzqI3gys4cgO7G/7iKE2nMxam4rkAKrG2N4Li17D3nA0vQxdvLx35
dQ5w7oIufkynxNzPrZD2js9MalpbJZLrm6NQ/RGmbdiNsl7zPLuY2rRCYY4788sS
Ii+rIE6x33ANENflQNXWpQgfvBLexZsFzeL9XyAOcfiSmjsgUC84tXJJPZ0+vh0K
lBTT6IkD+qBfMarDyAE18q6TwySb1eH2sl3r1kSkgPeAXNOqL2WmREIdGvrWwoxA
XSsgPXlTQt3wzR8XwUZVr89RKbyHeUIYLH9BOmyZ1VCmxAKUzDgpylFjbV9oVWw+
pCjJyI4Gz+SVq1/bSKxoO4ufsxDiz8TRK9Z6NwTYBLMRqdfi4Gu/HViTkosBB46D
ciIkNjJkekJcowkBZlH6zzoEZiRW1KKA9IPQPhrYymxuamJdbMhLzWx+ucM+y0JV
yRwujbfLDnYMGdjNmY5qcVWzbKZjliHYr4qHMZcghJJlqerbfbczxCNJB2aAcN0I
nMTgSK5Nj6G5mdfUiX2VIAFQiSDUN9awksBDSjLdr3oKk2/+tst9j9T1tIsoU8Q8
Aap9GI0i7toWmpoKUQ4QwzK/ldtG9UU35/3n80kd4aIZVXwtTrT6aLpH1yh8CcAB
cMC+td9sPgPBuQL+sBJOuelYxFEsRbesnjtbvrx1PgaUJtjFYJCKv09mq6m/Aw5J
8NOtSVRs+0fiCvz2Cap/aR6l30fJFpa0txNg687D3c81maxIhRVG4WUijx4wpsiM
9ls7g0Q99Gi5qDHccL+viTcDvegTPim9/JNG93XkqWwYm4ZWPv/sC+r4shvg2tZx
VRbhp368fTwY+N2H07PUb+Jl6UX6vlQ3kYXbeaM3pj1htonhAIHk1bcrDDjDPSar
vto1qY4JQ0iKzw0T1UjGgkHZ5T5hkHFUIfKN+FcRnH5SPk0BKOK/cEFZImzepL2w
+YnSzylHeDegFLu5fSqy53tlKm9v47+/0MuyQVxhfnzwvSJ10iW5i/ZVlQUqCy8/
a+f9N2XZVscEmt0qYJFsKZvEb/ooe1s799VawfsFqkanXU+XM+ywAer8C3mZ8DZN
9HxvL7u+1DZUNh9w/lwi9XUlMl2gfRzIWIAJUEPRRXDqqXNJh4ooga6S0PeRYjfP
l8jK4W5NxD0VHTfHY7QdVzc6eLgcWXRG5p6tviXeIBG8l1HPKmURATRhyh8pOjis
H75ZA/OFE8W2cFxciGFOotla5dV1uf2sPJwjB6aYhykjW/f/5jUluceS+/7ZxNoY
USdfClC0s9sMZp2fkZVKV2EjiuyiLxIiAkLK3VojplWDvEaOAkDnDDz/aiDNwZme
qYzJ7UTwkyV9iPKpFI5Evrl3ehVjn2HHUZwq66o4y1p3vYMd15dlG3l90y14sylE
GG1xVpJMeO91Iq+Lp1ArMIi+pPk4NCpR65luUuAH6vjxNWOcZNB+w5gEG5LIjoPY
0CSXTMErTfA8xSblNKnM4Xcz84xBMeyhd0INMXe4ngx7QosQtav8f6yQhvGWYuAE
BJPw14Y1lAQoDYHlRBtG25NQgJ3x5cqL2+ahkcF+JoqQ+0TUhGCPzCQEB0ZyNZxq
XUe/m6+G70nMHlVx1ItkhAF+Y1udtgJInEB+hIyVIS5nVGl3nuad4IDUOd13kw0P
XG9y1ufobNv0IBZ1fyDGKkxWJatUyO5WVrjunA9rWZRLAI9Csb1UhMTBrjqeLGcU
q8aPI/yyQiV3BZfWZrXQN+Rixqy9Gjm08aWocSWsWupGUA6/iSxi90oxuQrKp6hN
joHF4eRTBcWIYJnCq/cCrnY2hKavER6chklMcMLAcS3yzKG9OMMW477ifek/6bbY
MBfR4y0UwseU+NC7ThSQH2oMAvbXmz7LQD9qNSA4t/lTu469qsIWO/Idg5EYZKd8
gpmEzB0GHO01H+bdoTeBUGAkQLh1aaZ4LIFb7YtuqdJexapsCBC78+GMBTmK0UtT
bMmAAUQ6137s15c7uUbT4GYLmmP5EbFSCdWpqeEfz0blD65g0gtIl6hCR1UBEZ/K
gB+Rq+lOXXjSjWtqStlTA2Pc2I/Ms1fCOyOHiZBhOrfaqp6iYil5EnbT0tIb2rOy
Rki8qv2PtoI0AprNx4qa1czb5Didy18HuTpiICd7BpHhvAgtnqE5dH0kdHNmTcqO
qZAysZWGCcs73OnCHnM2lqLuodNldLDUv+yUJAwBZc81qgFe11oygwjwh5TuZIMS
5TYYywpk5T0tVci8PLQGAwG1zSq8ZtFyAfNyoPimj6huhPFW5x5+94HcrvfndYSe
q1QPzrQgQ3BJ0hoyQze1ctvVVzElEjmiy9j+w1QWKXnepcFlgzJZUFZGncez+6Y+
NzZSLcVi5juIlhNymBXzxiYO1Uiro7HpCjQi0hE59vUuXJ9JSpmK9duc9xBkeL0k
6nKILJ4KzedydpwBgq+kUvMaua4HlWpsO8/OUcM2no4nxIsOt7vkGHRnCb68oKlS
Y0d1+bkA1Q8hY6zoVloTPFtoZiegfkcgrbFSolrjt896rKiHIgdhvjIkfQHftPk5
SgFz6sgE0/U+a319ronJqfYeMdnjSKtliE3KGSl+p41AnO1sIiZp//lOY29nSdMb
5ssCUl5G2dvt5OB5jMZ7qIy4dpeevdSYfuzoQY/zPpG13gwl9TXr2VZBTQI8L5rf
zKgIORJ9W2bg1fRnt/5OJx0/u9ZOb1Tq4XNQFwfqJaMaiuwXX7lfSiwFveMQSk9S
bAQd1P9OxTQqtX/xs/7Vu5GHhwCeFlgvSe6qvfC33Y0oPhbl6qKWpg8PQ7m80prZ
I6HyCMgcjUKK42TiHwA6V+HaVZCiQoHhQJPCDsSa/n3iQiutfkVYAMakcW73JGm8
Rd8C4ji2o01xg0I7zZWYieqz3zz8iTxpaG8YvH/dvhaPE1/iAv/qOdGuuhM+aXMM
Y7+M43j6xgZ47frJP+lAPjGMnNj/TF5jgL/TVyUPVeNq4sbz6egrCD6TVq4JpbJk
4wjp4KvKl737FcJKufbdwxyJK/fqtOYjPWK10qoKZwGiqgdzfLCJ49i5Ct+4zA/l
6vlp3eUtkP5V7x8xOd5vtg+R6o0bqdlLEWd2I9b3+1gpDbnaYY6J02TCEVlNMAqe
rqIGV3q3WmWVescutg08La+wkoC9lOgbM8ljLL3PYN8dsVleTmASfIwhtcYE+Ipn
qjToyTW+wV9F7C/wRyizb6RV0ponHnZtDYog/03/KlxYf8KpW3aQy2t5Qig0nKhe
W2RRLMsX6VqzlLAct+msQ6ppmzBKuq8w9S/45ZKMBHo4krposVUPhaMLSrp/76EP
vzRXUM/bsxl/fBkd6fsu2Ka6LsTYKrdObuvM+xavTGWUPdS30v0Rf3ocTBvHwWg6
fKF2RL07mEO6Lv9HyWuzVrDOSjurgeYavk3VMdBChBTTE84hOJIwrRHHm27Ky/VK
v/6kTgy87pcr9BlvvbN+6TnMSNWS/nEy75C+FL4WdPUac6/BMyupYFJtBZWoWOv0
Ug0yZHxYl0tj8BxDN4r9oOIvrTPYBwz6sDshOJHaP6rLIT9hL8aBxe1GHm1sRR0O
DBJgweMnIYEvCBfgY7X5aKa29P20SpeYzljKEvXXBFOFHTIeQORIMTHd5fxek9tl
LM/jJfFxZjLhFvze2SC3SkQHQFmA5FCm9SllBiqV+t/vuR8/++VdUUQJ0L6rvhKv
3AhCniqHGRsNON5nS+BwoBjX0ik9fVydzD5wMuiRs6RHbs8EP7e/ovkW9KO4uqrG
a7AoM9piMH7srNPiLVtMq7EBi6kK+ncdBuPT6M+8m4pAGgOysbOFhEt0GVf+G93P
R+x8M/WOAYf5bQFfA4+PW1Vf2/DQOa+VTGXWwkRhkjL0t5ziAutxrRPIkjrEujTD
yZ2/CN01DkDZ97vfZ/eRpTpDZmRDrQ+gCh62UbyDZIUuZxwFGFXr7cuTbYLoI74A
wd4Y9GGQKUwGAvi6DZQExuWo/UdAnsyE1nLPvzAk7lRHIaqgiJKaYHVupupthg6s
4gkrgpNLJMRFT7hpztCixuW5EKwxGoSY+ZoY2hT7d8QxpqFEDsmlqPh/DwbWbs0U
qAVKaDwkZNJBBFtHvK/NrOQRAPTFZz3eVjBJ2V10LgaFLqoqBenmWU0XmFrSwPAv
zf1RFzrXkKhG7urlkuPoLKZl6+73Ep0C0mumNuhVlGX4ulStaG86yQce4gj+AQSK
T7u87OakPrW///QhkFfZo6tNezBUFm6nZbB4yeGmP9rEqaYcQM/6ciXOxJ4SPc7E
kjIZnjiWGNfyptSdNw6OwXZGxw4kcEF9yCXFI6n96rhouQLiZOEaojxuOlB0qKpT
pgZyr1Lf/aBKoPJT9wb1eF7APHTLRrAMuyS9zgjshvW2LxappMokxeF4tYcf8Ueu
hWBrBi2J+raHBNH9QAGJplmtHxgQjSRDOcXxJ+Z1B94SPMRVHsMY0BmGj/A595b/
zZXJAOWZRawLykXUvg4KgqkTphz2XU6neGCZQiGuM/dTZyHvXS+7+4QaF3wUYDCu
MQuuIx8nlsbXiQUMn73XwHUvYdWEUrz2Kf0eHqnXnFzkkNzVTSrnzT4XI8I3O7Fp
bj+igJSihlwI3rxdwzm6shO9hSDdKJZ0bDwPN0nn4mlypYdZBOryP0ytqYFm3/Rm
ANYAZo1e7FZJ/4dzede4SOWLh8xO2b8VtOO14vNQEUeEsyUxhIJoAwKpaGQ/YjX1
X3752zBWuWtZqfZhBJ6iELm3WIo9/3c2yt2Qn1l9FU4ynkrdQ2xxyuI7SEs+JAUW
M4Jep6WF6XF+2C953PQfRzZJU01mfrMpvkkfpZpXDaNmJU6kUkWEkywC9ZW/fer6
dAcqsM7ZMbEHAnUKwFDnLTPoD4OFRt72dprwbLjBQUYcHuF3f5zT15zP5haZLdjj
/055bRsTBYFjt+W/12zAxjIGVYX4dYUO8ZYh0/S6f4dOyL6kKF04Cv0f6eK6odBr
82DaKxkBuffs9P3IlTy4EoVMhL75smRj9GVk30ph2/QpISVBpf79+nFyD4z3Fdda
d0Rw7tz/uBuJtcazaX4uivFV1u9H1qnhNIRtdJmBM2FDClEBla9CiOrAoAYtEfhm
BiuW8K6XSoCSWBraI5xKfKc0XcW4HYTteBVt5BleMzU+ckruOCiKoyUAD+mel9n7
+Os0K23+nQeBUlcqTfkLKibrTu9aqXZ+Hq0+Wdbus1m2RBjESCt2T1VYHi87TbFd
9sH5FNrPriCFi43qWZWEiBpsi6XflXoi4IZQ+GsC5TYBPskKOXAKyi5eke+uyVDt
VMcl7XA5l5SlXru+ekb3QHxozPLyvSRsS/hEoZizKiiHLZ354atLPewxrWWbFHMu
kgnbfwz2MctMALNxa7nCorCaJS7jXCcmaS+7dcmd26cYyxUS3nZZPzdvHGf/nYwj
NlPcPs3s3X4IvfeQ/kfPHjHPC2KIzvdarPSqCMl7r3BJcDS+aC/XEjbqBo7t4NA8
jzQLEZb5kotqaua+k4OjsHlObqDDA8yuPzV1ob4YJVJ1kqUwnHwWMTleXWzdL8v1
7IW3fC3YJ5x8XtMNI/uMatAK2Et7mx8cBdslm/xoWLoDAP9IwSAfv94m+3pGEphp
yPiS4jWf6w5zJdiZ0qLErAb/cbZNxdEl51uAfz3EZzClURD0advtGpHScMcdOt8j
EY/O/cKc06AQbGmAci+jWZ49I4NCG6R3GfLyyMEeeEhBBRF6DBohTdZC99PtiA1k
VFpGinwVb8aTuW3d2Lej/ZkRD3fxM57dGDSPjlZs7qzz3pAqdATtOihBe6Vxnn3J
XA40KsBONID0oOQ+hfP2OTy3o334i8LEJZ2KeMy5TNl/0WDPpLxPfn5SJP7r/5sE
rBUNiBXqZNt1W7IGfmW+Sta4hzPYcdRO2pOK/mj5svFKJbnuGI4PZ3NOoSPXSRj8
7AJpWqVNzM83siBEEB1fxmRzniTaobecO76BUtXddtWHd5Yg8SaA7HvzHIiuw//P
3/MRzRN2xlF1+cUHGURfs4lzgPMOsTGyjKzqmmE/MAWX6UomUfAykb8KqwASxPry
dO+Z8HUhjWDSgD6iMxs0X+D1ulFQ6yCIyuOEipDqpc5AzwxjQXO5BtvcWmv4ze//
Tm/j77bad8VplMFzRp6uAO5K901DI8usntR5CJRtNjuxsoagxl6JMwvXK5ku2htV
6YHZm/V073dKAfn8NmQP1DeHc16rlxlUDNEH2ihnb3qur14CmSMk/dqIYiW15y0R
Nuz+Mt6zjeg4argqP8REtNMEsnt5++6BspsEFHLO1GdoTrbauHVcyvlpBM5xenCm
qx+E7kiykFM/aNEiJ5RGrTdN76VAvj9+kVPGll44nvGxflAmjv0g/NyFlkMGVEFP
6oO3reIv+vmoQhooYA+Z3/drwxuEZvbZWJm9GP1yddvsLFo6vt7L7esuEOvWeweD
Nar1TvODkLZr2hLEhG5zrH5akNuy2ReTeD2ElqhzT3vJDoHZxR9nJjULdvmZLnAS
SWBNYu5fYS/XlqpejjZb33oyudWjSmpb0A6NeBLX1jK2RVpSr6XYCUUyXtLwWTWA
ugCwx55Mc0V292dBtqJDz/DbZhB78uMd1PIEfPPWvnUrIi/Qr3BqSYi0d3m/GHfE
ktXIyPQGacIt2bWsGwN9AvX3ro1xNharyUw0/Cy4oZdMBEq1vTSNRO5APO3DANwK
LD+niJG5lK5fyLNs2ApbVNeQWxQT2ECch9WnhRixwpxlxaqMzGYhiuWzfZAkof8g
+oCYVzuBWghqXW86r0oKA3O2FtDFg95p9toacIqggHNi9JuZnxxwRdBCqUP7lVem
yVRz0wSkao70wO0wYNNxOGLzw9mLk/ktIhfte1Y3DQOI3YoG+aV36EXtMv564fcu
1o2xShyff14CSrpo+1Y4j17ovojFYnKcggsFgh0KM0S0y7KGfcM7N6IaVBfvNsUd
f6eI8fUe8czs01CWZ/MokPHl0hVdknM94uueJ7+m1tb9shaGToz24mPfKuP/O7Tm
qkE3AF0RfGHK2oENm3VI0E7qnpfNQVivMwRj52aBmd1JQkQN8xtQfrsIWtuY88FG
JBvEQnbr5N0kBbqvrI3XCfM0OjYYbGlZVaeKk8f84V8b8tnzOkxJA2lC3B1afLaN
kyFVzRPq0a+7BkUp8Mg6DLloD9+t+NCtaVs12LdpACjAHuC2hkKut03iVQaK1hmf
Y3p43fzSwz6LfwkZAbdMjlX1m+JMBFJOIL68mpDNbgQe6cRkzwCwGlWYZ1ppgTWj
SR9MN1vd/JCVNd0GK4Nh1xiYstBu0nOYwKtA3L7AHLQYo47+2+A1hwFi0l+riMbe
33l5sSV1Scc3pw3XLlMW7wYod6ZNbJZ5PD92KOUy+G5o/PlJHseAXyfrU9Oe3Doy
BPDuhSCZZiq52furFjHcqAvQMkl9NLD6jpj/DBFpGCI57pWco9ulCtgQUt6VRXub
Ns9dlqJJMjtuXIA/6ghNUXGQ6qjBniGK2W7cBC8FttNlZMpdIbx0nN+jPxi7yE6Y
K7oxSEwiN0iZWZm/0JHRU8/oEtGVRvE2bL47lKLNNTpk6pSRzUVOl1hXb1qHZpSp
+5ha89rCenEJctdnMa/bplrm3ITq40ugR2YZD1qPnxXTQD8+314Bm/Ia9Unwr3xk
y9t1zcJ+emyhGmGcZTDnqo1NJvO2lhulxifGo7C7w2xZcB+7AhwZfhGMXXQFspmr
1Fgc65mQFV0AA6edinUB2XRFR8aPb5hU+Sc1E50trvi2vmizt0SlgC4YE43GXr7n
UigRd0Wd/xO9y1GIb+Lj1kKWfB9wOw16Cu/aHLr25Sz+Dg4DpceKUD26K3YTvTn4
rGQLs4oYgCXXcOtVtGtZPlnY6luK2PgWonSVsal3HflyBt8e4l13xEJUwP5irbXv
xBs9DLp0i1WdIXTs7X33qCc8VK3xPYiNAXMbggA3Gsmx13bZudTBi9ld+lqQenPQ
p1/5iRRodq8vglKlAA/I41e3a5490bFy8+ot8NCR/6eTdEXw0/axjoqLVOnIffMP
6vN1IEER7pFqEu9iC2Kafzw/p5lpTslkgu0DLQZogw2slhfsgKpRm0FyzNuq0nAO
8K83q/4dJmBrrZFB/gHdmlq4q4RDf8T8q8+HHHSDwXMgGkwMvrCWLJnWbzitEGue
6FzmRd851MpAjuq0qT6kGVjaKDsLyLuhvFC7sIFSBKJhoxkBHdlz9GrQgMgmJ8vl
5vi5xhHCxJEPDT3zwRkmjHk6LCUivIsjNpEwNl3kn/PxqlQmQdpHvoCUXzzdJPB8
lIANOIWg+BU8bufHl2w6kDlKuBlTPus5hZvBMlUGdd8vfLpkwrDuDHd6Jg5bk8NA
HniQ1z7AihB97u/k5H1vIWeLKmFNhYSF73zh+U/C5aFJhQ46wGvEYG2ORohCki0+
awOAkWFdRahvUe9p8Y31Ow5HDqM2G4a5wQ9IFeyHp0PXjwWuDKtJzVxcwYFKuln0
SECFn8kuQnlJkSX6WNrVABXBctf9LpZKx8r/8XPkroQTn9eJ5Y9Kd6x9ZEvj4ph9
x+CtIbAv8lYzzkjqWL7O/OSY7D4Kx/qDwmlaVRtH1kP3CY3D3e64s22dYzNCNOXE
nvicxPrHBRV663kXi1q/KhbuQiB85gJ8EXMqnFNiMVRNNkXcB4jnG27mzJ/Dq5Wi
33n2KTSvUTogBDHk2XhjkkSbHrOyFGXPGxjvGw5oixas5MiS9mKmV6/Djq5Q8PiL
8wpKIRRblopps+dSxwUFBS/uSlpG/a9cGsMiPgQtneZv0sywfiYZomwb+5XPTj6W
QlKpZeksf5RAlzIJ9wnFE35u+6r+dQklfMTANeGXPgQTJPgzNyl5Nn/UUpBNW92O
WIEiVG2yZNYg32FYLvHxHQvP0Jx/UqnQTpTIIzyzIX/65q/g+CxHSVmpGUTG7nWA
4yU6HF+bZDa32y34FNlT6WtRAkfjWWPxf/SqPZV019g1SpXDtDJXUasGb1onuQ8w
73dNihvWe+o5EAeOiHnHb1AHIW/pRnAo2RoXlIgl/egXI3u7wrroNy8ye847AAEB
OOov2SBwrMdva4y5zGimu1PoSZJotehKaLw0PLrNYDKVkzBVE/DZiwmJ2n+491fU
sV26KSR5oohLJqBLJ9I3KQx2CjWAtX8d6L8NpQUh5tK9LHNoUMmt1wXNLdhpV7Vc
Efp0ffI9eu2yN2RM/d/7QUOUxxgndMulITPuo8yGeUb7eS0/Ke4HeOq/wIWlGnnj
Q442LIBd9N8/0LGYTABRHqOhUov4PSQGygdz26fLsSwZKWCGxk7k3+KyuZcHhY+B
UcLhOxFgAiUqtk6e7XfuxEW9A2QbT04d2Sg8kyiXTIyPX1huSl10v7Azc6y1O0T8
5+JlhGOo/rTEeQ4AwVoI++6MXLIX+n3FzXZgadgVMQHKjrxjlZeb7X0v1GzM9XFN
nWQubQWPQ2nj9Zywzk90dP31QSTL+Q13CiIWwbCbOjNfl5G2Kzj0ttrNee/E4vab
khlshmpYNFuTxjbjDkcpsY7oRdsPr1eMleDbyx2akVV5mRujTsjhu1K1JSsrg5Sj
MXTB1MOxsB+/O7dlcseKNKta1Vf/FyEmFFfiKjDcvyZz8gISc+eJ6hm1OuETFAso
l0PEmpK3BG+LPnBn935BQ0NU1i2neVvxYTzZC8QUbrYLTfborPHOEXt8u28JCS3V
2YJuJXmsfXNy/D4xrEynob697YXoPHU4Cc2/9iPUdEkmOXs2MupwpuLChHarqU8t
EqgoMGKzjR1lB15jNfWxjdPqHUS/UIUPrnsspQoxTjv+VX7EhqMGE5DIAg5V8RBB
j9BtpUoRlkt6/bEtpKJiS43D1KO6Lvwl4f9P/KyOzUmIstDl2Iu4TL0hBosNekUJ
+6BcyLWfnt3aqQ/XuFHzeBXVOVy1NVvKZbb1rGDFn4EvEBTUqqZIS2fQAOAtfnWu
xupoxStqtj7Gp2Rcpu/waFRJX7sGP636Ggcs5nclLTSbO+NRGZB4Pq+JEcaD+CMg
fhx/RiNfhjO+O4G7bgA0Lt1QucxBy1yoxN0ZwexT+BEtEhyWCe2ke0xrNUSiR019
HPJc/5ZNSQXQya+rcZCe31ba1Aw/9xUMf0wqbOz/+JG0s6N/bFDqzN7R6qHsNJa2
QRtp+nu7Nym8uXz8hYawBGHNPLGcLXJfaBYs5QIxDdWQzay6txakA2QQ6PeEs/c+
xBeBC4zIPs0yJ8gAHREt+kSu+f7MT6YHMk2XNoDfpl+OVWgUrqAm4xKANg2EBc3J
UhB6N5/lHoqVuz6TyKjf/bQYNOAiOZkbsr95ARCSMMz8PkItbV62bs8hyMBS2EuP
y3STGSgg27JmqgbKOs7cp2DHaE7AmFDbpwjpsnG7QD9IIl8djrNRAR1EFyCm/g9p
5afE4BupudGQNc28XjZwce6smqWyNQM2jKtCuLpl0oUPUchonIcI+ltdDhg+Fdbm
+TeGM8eJF/2XI2Os4DKjaM1tbikfOGMk69SW4bqBvlnphD7NBY1WgNaWDRkMT9m7
/VIXqZAGIkjI8uNc6sPu6fdoAz7WYiHjAY/rSkz2d54ysR+GXjtP2fQ9HL2imVI/
9ZOLKZ6frmHb3DMwo7t9RmXj43RSKb/hRl0g7PqwMh6DwiMIDWEkDgdlwV/AukKq
y11yl5ki6J+1ZcviZI05sZDlGZGMeSzIi5bgCtjWDpIhDvVD8Km+4BwB/IcHyi4v
Kydzv0OZvBL4Ke+VZjdOSDxckoCrnKcuqUBmHgyCC2DaCbv4dLRHJXTzb13weCAd
zpYokeXjEmeVmz+6hRb2yodgaYyyedhrbGNFm2mKuE9cZ0Ia3oOFmXE+n6L+Kb5O
Ft7lrPRLB90lo1Y2CKStRlzxLFI4PfJMFl+wJTi57OTVVLL+EFX2M2wxMZrRtfq6
1Nwobfife9XI35AqsMaUwFKkWPfSFKF7LKsY1gBFPjHyQGhrr26g4l6u7TDHE+Tq
zDCnLdTpM7cLgFaUwqRCCyXA687ClGgQ377IRHYkE4YEeiX+zk+4i6iaLaSnFsNN
QBHVNtcUhU65Edq1uJkmyh19FhykJSIX0vC1L9k1GgrqEK1iBBmUfNxE62NcpKC+
D1/iKfb7HXftlxIwqSwY16Z7rrnrwBCCiYRKVL6TK3hC+lbiv1wf4BM34+UiQZ9W
myTNeFPAt+VVo8BJRQpF/H9bRMHtHX+7c7bTyzwXO+Af6aeJ69V2SAEVJDCXmT1M
vldFEg1/0+4ZIpWUal+iXXThdHn52MSvbcRfpiXNqw2sWKvCfAcFxJ+jAjL0Vqw7
HJ6tP34gdk6c9c/ZXBZ1NpsmxnWuhRSNsXjW2szLcxE5JGYwXZ4NnIrhovkKSc0A
CxaveinP6UPAu3Nq3rXLQrwRbDIFhjZZRQEGy52nWiByjrW8b5W4S4+M5oE+kxVg
Ihqx5u9zwSoB1tCUCtEH2dXISjZSbfdiQtx/cBQE1QpXRxbDnX6XUYv4XVh8ATNS
A4yE09mwHClYyOBS9MNN8bPYiaY0zrBom9mseFRWoiqFqloU72k1geL4gM7aD/cG
kA36WL1h1iV2FEYU880WyX4VsDZghZv+XoXDt5T5iWOrXLe0x/ZaGbdT7tFQDXVz
WFnWBHKypFU0484eLMZVUKOViOkRJrCHteY7JSgMT2PzLKhXv54grrURqw4mn0rT
dte6lSjKqugFmg5y4bOhalvWLwf3lv06jtkxv43a9XC/sY2vvKYQC5y1wA5b+b0v
+FJbJi41GnD9M7cPRZNeUTkGL6FrOF50QOSF4fVmgzoX+jnr0m2BAeqxfdQm93cJ
fVZVyuEUfjfzvX3bmY6GAOxUKD5c/KJaAnQrYkq8W3z/U/4AqrLJ3H6XURECKYZN
ixQ1+hNEkneNLqAsVG6NyLVKdO23v8ud63iTYN7eyBMiMzr+CdJsHbGU3L2rbcp5
37lLBpkQeXm6NzqWF8/ljRMLvEqLcGj2jGsfqfWDiEwxIMrRJkjOXypX6G7VTLg6
in0T2Ei1/726JcC0Wkkj7+h6h7MmGhOiBFfbX1EpXNgoDASYEBBzgQcFzjwREd2I
o7aHzAmGTwQWkGP2biEg5LFw2eVe6FfxnO00cnExOsTDGrNsIBWWeknVvh/MxYAW
55yzi5psC3WP48RSP4G4M5L1s8jgQKu7MZF7W+zmE9qBX0mWM7Rqo+dvrMmA/dZt
yLWvxdvpFExyl4P5DbNOIE1i6WA6rGZQAA0MPds6O4H4STFRin/h/0JBhZqvgJ1a
pYpEivqRxLVtYiOLVX2rN7UYDR6SBskNALkYK0LVMI5JXPr6fFdRs0KbP05SUiwY
HNjO4Soz1LRBSsGXG+8F62Qimvcqsux8ONiDs4TyMt4T7SiPcfnQ6hoh4Jq1wGxN
t7q1AuJN9ETFHxNdoXynDt7kjiavrD/1qrthbLwf7KbRefPQRYmDG340u3CqCeXy
C9s/hOSU0XbCwt1PZ9NbmXBU9u91m44wbupr4/B8DzlhV/g73MqgvrDoh6CFmPrz
crP/e5o33ND6JKAm1sKH1zXOO7RFTKQkeFwuvlZAoZBY9aF+i+v1c0H8mJ3oQCAl
wUhux6T8pT4KBzDohNGdBOUXu8N/Jre7XRdT1UroRNqzlpJQUc+f2DUwBWmHPWZI
lMplOZ/1AvKfNhJLOPxhdTfSJFhXUoKJ3qrbKCizPBr7vGCNoIqzaFktFtqKgNfm
MygF6IZ/8Xt1dMIMzpEy1GRxSiInbK5A1yIjS6V65iWc5/FiPQ5tDRw/APu5OI0u
hpyZ8GdqeqZz3LRwdsmGM3Rsz2PG1EFY9eSbV5I1sgkW6YLl/iXuVTPQHPhxbDXf
zyu1hse2MgGFKZ06LyDXF1fQrDl9wkrIL1qm2PLscEaORgLunavVhRp8qJAFH3/H
7RjKeJ+6KRwh5zJJx42CWQXjTzrZEGu+7HeWhJmxtWeyf049o8Okq2LZVCOZ60Cn
fqMxHab9qFMP59tU3zE2a6RaoH3RpzTpO2p9jPxLpfDuEUI9orLJKy+oBGyUPXYr
S2ycMcHuudsbfKrhYQAfpam7u0ewk3XY6rU6DephYSY9arZY290saIrGn3CGocne
CTxkpE62v5VJD/NnPELKoyGUADgSKfSYiMIX2OsVGTcNpNOtrGnbe4aPAESR5LRU
q6IHBit+fflM7V76EEFsPyN9bxT5sLcsNm7tWYlvmKj0qkK0LC4UdCVMBgzO2+Fl
yr/1t//RcaT7JSp7A1tD8FrOJukYJPQYhJ4jk9RAp0IPmiVkQceNBsLRNHPPhfzp
ZjVb072aQU8NgPX85FwqXZlPsC6EeaoCEYg3gxfPhQ20VHIv29gHdM9joieaimq7
d3uFYBbGICCh4L4DXg+2jJyc5P2n9kn6ll4uQDRjhkVLkdRpl2kVG5auSIfCOBYl
VAs1CGUtIlhl/eS/yWFA4d9nTbFCANyr9ZIJA+aOHVu08tK/2WZeZN/P802h4pEf
82nLJCtSwmcnt7zCJ3J8bi7DvyhWFj9BuWU66eWIGGJyBqKO2sOIV8F6gc1vQE1o
/XA9ZwHxB+4kry0Q7vxkuG78hZ31MJMRPRR27FGlO3iphlmx3dgWJh8gd7UXigQR
3PDorO9rc0CuPNCnf/tS3+yLiN9UcCxLVGr7zLv7DTazuAJwFYZLGfn/DeaMsDIo
BkdzVMuDvPdkyPz5WC0HPUCGSqo9Ljzn6fFMRQFgkJ6bXOWAu1Pd3QUAreR22F6E
wOIjD8ceVUCCtirW8OP3nhOx3EtCnMgA3zVuaEWmsnAKnfl5HiN+0GQf6q5BYhAM
bjLZVr3E0BTpwPIg8m6Fzi3LoZCyJImRkuV6GhcfsA7SQ+Y1OObPtXBz3s3GDVB+
RbBuLKXGqtvc4bypT5U4oaRBJ3n2iiPOLgWXfFK/Xa/kldwoqIC4iFY2AUjx00iy
X69VElPhQVUoSBS4aiogNsSlnNbdLrk5Qzds0iKIlGj2F1r2QV44kKZHp2h2q0/Q
XJu+Ed4inQROcAdOm4uXL7sBAAHzOQcvB9bHHThbZvn4pnH4HSvE0h1zLCOeaoCn
foM7MR0wTy4hG0nthExxU/43Vq+vdHy3ERd5DAuYFoJ5rDxok2zOeW2PtTqZQa+M
eAOJhWPpZdqbykSi4Klu+EcJJ/YvMR6+wlH/64ccRXbK6QGUC9b0akj4Gn1NV5Kc
1WhXg86HYkbOBedJskgk33Y8z9QyNsqPH9PNv4QcdAcv4y7e/o59frkZAcOwUPbJ
FfqAgtXi5g71GJzK68cv/Dz2v1/mgVsE8nzSqXd0NzMPjEusBmOFH75Oi/t2lkZg
eNAroq9eXciOWkQEDYFkTpd3GAvUEB56qPgshkqVLpfesTGcuSMjTj9yZH6CHZp1
vVsttFr4Q36JzGFjHDWYR3g0UNF1Fl/j77YBtNx3DKtZ8eS480dMf9KJkovTPaCs
1Miv/3u8SeLv35NvkG7YxUwinavbxXDIWMbtE9OPMWuAOomCjRZCEUIVqwy15Ffe
cxQh57n0uqumWbHk1pxJe7aPYh7/CH5Z3RIWQPaXSDoySlM3Fa17MNjQVHec0GZy
DAzyQVBVTFS7UIDcTEJnDl6F9P/TJnz1vCBmgn3lHwUenOGVS6CiVrnArCFrq1bw
1wwo70le13cnDWwqtR+1gzTR/Feehvyg9nvOlvBhsSKmtM/gc4GNsyMmC8d0610j
4OkmTjLl6mTZLCY+9f799uiqLRcYY/H8qDOa/PvrnRXjtVWKR6G8yHX8ey+4noc2
FonWD9wI23VaGspCFQXkvZ4CgpsGyh1p5Gb53k9yNRJV0Lf1uXBd7uehBREUrknN
F5K3stNXGemvl4J5CH/1HKf1oDlQcnC1l9cFXJgDlNJYk/3+PJe5bJ7db7EolsAK
TjIjvuv0dx93jntrqJ7IQCKjihVdXqeLr6gj0WkDCAVDQqw5oGq2PVE1HwBo0PLN
GNbGHEEu58507NdOptvhgoL+spvTvVod8EL0UY8x+hob7WGLOnWGRamfizlb7g7v
WppjNrUUBbfE9Mxa1pVEkIM9wZ1Rt1NZPC8OoxIyPADEp+VYv5gDp5N+hcJCAIk6
qdNNGbIo3PJyEy1TxQqAIVgfGpLHO4cc5RTBc/gTF4FRAVUkcAOj2HWClC+41z6S
hFsLskfD99O/u0gsNcE9GyQMNsFw8dOl9nAECDeX+ZgKDwIPCqzS9jB6Kitczcvc
3VyMNaCHmodg5GCnB63p2/OwPZMk7M92dwMSzyX9Ft2EiinMei+Jl5Rtsl6sCH0x
OnhNhHq3T22tX6BBGu8yDkzB/CflzPZAS2T6JTCs9JlOPjVcdq3WGILO9Pr6g0dL
m7+puyQ8yPSVqhXjO+IFujLdyRPLZ4YvNGRnNTeV98Sc+paLeGt8+LJaZWl9HsRY
O5jmc7gK+fG70iNpCxday3EMDcDPFrfd74krGH//elrcwCmKloYhSGEuvvWWg8Vo
TWAg4Mk98THagZppFt7oN2mZCngJntDv0w7QQm/YSJLoLrnuwnVZB2LRMKYLl7oV
igzlW69xeladMf4aWW5f7auQtSv6JNpZRknIDrZ3e2OvjzDy+kFQDQsDI4+f4HPe
rCmuuugeM0t8Rovk35VMzb/6JQD7hIOCGbNsBl+4NulBzxmZwXnYMdvXvtcAJXv9
T1p4x9hitdeyld81MHoZwTMwzqO4P/0spZ+L5utGBl5kTz7C/f7CCeSlEUe4yTlJ
9Atrw7qj4C3JwFPbVvtD1cqs9UTWdeUmMpkEA7WZPYweq6t6guKa423l2frJrcRG
RC3Br2YC7y7iVU+sbEWDR3k5LQbqRdt7gWeJNg/Lh0akskFnNRFAC3Uu6ffSLetO
J63pi9juDeqNlsALKf//jtGdPu+s+JDVYooImdI+C1YmF+Kb7CFRMUUqOrRVPqX3
3CwwrZrsvAWT/1GNqYlSH6o4IKT4z+ZfVVTZ96Ii5G2yJ+68JvuEjyBFhYSUcsWX
EcCkagtd8RwYc0qV3gIYW0FsU/so4obGW4AprKDzhwg0VKcRc5o6POoei5ljl5B6
rMOJDLd6aJYa74uAmIN3Z5J+qwZ4tYUtkhHY5/HaquU8c1Eq87T60QeMeI4n0WnR
6haHQsPsT4gEHNIYwIbXyoUtwVIoKd2HTNq7Fj3o/IjBK7rjrRvYK1RfRS8Rmca6
ZbVuh+P3cmRmcnVngTBlognKD5Inp432Ew5shvuq1nRpKzPXboJdt9D+INxtxGqj
QG7hxtZ0T6GINMiRLk1fl1qVTV4L+lyPhGP61LIXi1L5JqQKjD8Z3gosZb9qP4kA
kUVi0FX/QKxrqfZZwgfE04gkvY6NzR+NlhMy6XXUg+l95xAazQg8KprnekAqkRCk
H2viJ+D4nKBFoIGtqMtMW0d8IHO+1grWGdkibYz1KLtpaF05JBl2vCEjk9HobdgQ
SUM9HJeEPwmuXFOT+q3BdVCNrJ8H9RjKTiOT8oiy81u7fXhrfCqgFfC/VYppJUAX
gWrB7BpP+lvgLhxNBVG2xh+c7Jtvo6tHxa1OIZW0YdBL+XNbN5col7Ra8IxX/XAr
xZkeEyydSs+D+hkb5D4oXKqLhSFbSBOxo7BqsGdr5QTim79zZcbcNCzSoiJZfmY1
7qMLHymCyuGGVWW5PFwPm/sC6ZWmIE4sL+vzxHh4JKu9UwCE4SzVA2KO6EB9Gibc
1p+orU40tBTEEw/2cIbCskttiZ89X6bWeF5H3RTH0zdWRdpW9O2BzE4tvrNN6fnf
4oUu4wJl9HtjgMPJZdV6TyWptwtdDKF4uJ8El6AMNbBR/lj7AUGsDPzDVPfosr9W
LEN5u7+TmwgzGoz+WgYIBjT4IqbDNnMSJDE8b5nX2ybJ68FbE3OAlajJl8M4wJ1v
jAZbo99mG8JnL4dA1z1i+Z9nk3kSEHoRlDkV51s3Hp1HwsLESeuICe8UyRdkgETr
6uuLHEAdZV/lKbaA7SDkNlPS9chYU9QNIPQA5AH17Zq/eCTbx0D2+b5aIjQf2Kea
ZYHMQaCmHOf97RBKdknuCgjwLbIp0Z1CKjCxTt71x5yrEbZneJ9bPNziCe4Ep7zR
WQf+sBATc6Rw+H2dfqept/XUy0ZfmYEqY1EUHa1yO0v5MtWoJWpEI1JDLKItEdzP
mXbrMG5dYK+IAqtVIArET2+ZUofXGIXx+Tr01cygF4TMx7ZzR4uJpk/L2EUI/CuX
bjejKvMH3HOgryi8rsTCaOp0b8qh6zIS1dz3hLJ8h43pLHmZ7S7jVg68GjLxdG5L
YAZErp0QCrVwhHc8MELDx7rX3JgZjQel4iCMk0bh0sL1dRcwO+smQrsyH/0W4G2W
JXnqoErAu697S0ZvXdmkFAEN4tkXmvWz5oiOva6ZHsmhfDk+Tp4K6xFczNbbLSFt
yg/Joigy7xE+xq5ZDk7HRfUZgFaE6V6swYuMzdu1x3cdCuy3kXtO9cLyl9WjfAyO
ERB6RWihKVeccgjXH7UhB8ckPsyPD6SQK06hfdqw/wdRlHs/HPA07gzigg47axRm
cxK692RrmIc2QJt5as6xoCRPcdXqF71cviItZkElUKhj7Y7dPA3FH7X7HGSgZ++3
Mu2AM5IdD1CoUaZ8lgG8P74Tovotp4POEPGVqeSxQ9Ph0hxrOqeJdR/c2qQ+88PG
YBphDl26vu2q7s57AhtiK3rp7ms4RU0onGXXjdRhGOWU10DxJSkrZ0rc0mb8Qr3r
fZ4c/NiUdBT2YK6SGJZwUuvrfiWDJaIDQlaM0MVepE0rCA8HTsFEKP/vQ9BcfmMj
ugIYDmQkpydGTwKOIf3K+IxKh9/WkSZhSfXldVKp4EXXvay/z0WGArQuV2Bi0pGT
Q9lEXCWpKMghCo9Tpkzn3/R8me++Y2NMXyGH4+HZBXVdZW1WV2NzwWn2kz1kjY4t
IQdG8nas1SLm6HU9JUZNkL3CR/D7GW2cwIeJhIhoxLi+5HGzKiuVuxvwUh6BRLhw
uCs9k1kZMOAJrSoLcI6oAlpNyK94lLox4o78JbdncZBK/ExceiSjjToFTGlMS/yZ
orVJEvkzStrw+MXF05VhgiWqjI0gh39UcyZYw/a6fqgytD1rl2qNojyN5/H0WLFW
U1C67s8ypzZYOfkBPCzYTE1gsy89brJ4EgpsdhCUEDs1IB2DoxuZ33omgjvfqIzq
6NPNnbL7ErSLMUG9TCkeTLZwXEvmCBKN+ezqKqBp77FGxkw75COgwUJUwdyyfIgp
iwz/4KiAmTN6NU9uvnr8Eo/UMLco505KMHc9UG9J7kJuv5ScZM8i7bqY2SqSuLVv
+mNtVb2RRBNGZT6raCvVC4tDMZW7ny/rdhljN4/bjDW8KcLU+YcQMnVqjIsDp6ZE
xTVsDFbys4TBWd6sXIITvzMDH/xt09QjC/+IomM0xJS7UOCGmQZ9W73z4Q3TEHj5
oaWCVyQR6tF9LjKhEbZoY7fBX6DeveDuyxGYXUm8uJt3096zrhGmi4XWaL0JEG+L
L1VwVGMFc27O6MsJuFonUHFhkLiACbFlGN+6ZKFepEFROstHIulXBY9N+NebZp7L
rOlF2YZU6ayO9lo0iM2W5E10U4h852DDW3VL1hTXvKD3muMAVjafpAu81XnYo0Yj
GdCLIaeo8dXekM3dVJNEail5E++fBnc4nw5oJxx2HBQvmrBVSRCTEeUwnmJZqqZe
L9ll1ileloyfnsEjd4W4ysz6olKhI1E+F9DoJhKMh4ypM/ZZ6QcIhPEtgC49R1m9
Z2lyxcE5y6K5W6iAOQT1RG4ARZwckpl8fbF0+58ZTfhnan+qcqc30IxeDOw37SOI
UUQrvIjjsXNeDNHjD+FmrxgIimIojw9SqpkhK0BaUCFF+ZMSE+V9LPy0qwzMHQ97
iiLzWiDC2C9V0N1semIkKfHztAnZ2WUzjZNUcw/4uyaNnMPGiTMljs2QcAIMHCPx
R0WyS7JFjnamWL66oTwzjd9hgBozzJ6A/bIc3c+bdjh1rpAQC4IKhwgVqqNBvq9T
H2C2gdcarK8U091MQh8+YJa2tzYW4jxyMwLVR3BXBIyZOS7zShufH1QslaRp2FVK
mLCWwjifaaFwVithoASam/AM0QDKiAGnZQVFdMsCaGEqiIFkH4i9jvjOslmClRJz
K4MeZvMAlH42ZAuv59KmRabNx3dU4vzg7st2yxFoeImvYQy87UV0glgEQFNRhEsp
rGeCGXtmpvR9nPwIxMGSyjbtWk0OKPYgbAaRjkRjvQ/rwwycdhwIbRabzOFrksD6
U8rdEZ36f0l4uf0Ne4u5x68lmEZmLWh0XH8KGM4EHKY9aHyAySIwOYgUDw8vZXTD
i+DCvaH16jKlRO3VrtBStvDoJMv+D38/smocH5ruAGG+pZqnsBjcqVySUlTIE/l/
xewqFs4gtThOs7E9IrvZ45iZvHImxymjfVbW1+2wskK9SnWCBriUDDBR4k4xVO5z
q/53oBpWnrlClj4nx3aPFI+GYnELL3cAIsVKJBjbZhrJ15wgqm2g2ro9H5YnG1/6
6xcQvHlnhJeo8ofipw5HVnGXG25/XXfIoCe9v8Uo0snVKF/ek+tumBI0pOxnnkt8
mcKOI9fzCu9UAt3Ki6pDz7b8vPByllZt0fQU75h7n0iOSdsX2fFX3tzv2LBydhmr
ajCLOhvfGE3K9pFl9YpBhHlvG0TADPZlCwJbvmInsKC5PEZk8jRXVfD5Ox/05v2u
0URnI+9SAQykvXxR+DRRqfmFS0u/C3oUzgWJzpnN75Lfp9KJdS7egHzCUifGEr3E
II9JHvVzhhXZ0i1QjpW6TMkCT/J9MMZXDmGlIP7bzKxXK4cnVJ5e7eIJS1OOb32M
1VDGCaFCOtDsQjLMluyTluvpGYXNZ9D/VUASxALCFmsMiDTd97qcC031FLx9wM4E
wFLpKE2WbDSFEbyZU6Vh166PkzQMkto82HQlrSLn/5XpVQ9vJgX8z2Ce5XkcW2Pk
3Jrxt61iSVhT98XCwEGsWTvmskw6UdL6kb/0AEWt9E8Tin9mB2UOpLVjj/jwOYM5
SJxfsqDflUjspNlJRIiV31TBeM5GRfTX4IEVDvOnIy1x7XXiTB86TAiQJvwueRja
rDmSnEsQILy2oJkxLB3Mb4SxrYUP73alLDpTt1cwaJ8To9J+Atb+S0ZIzyL/yDM2
Nv4DBcIm0cYoIQ//Nm1PB7WVDklykjSXgXjpNmqP97+RJgr9r224NY8Af4VJcboP
s3SAS8N8+sHuTsWgg3bVW2FKUbHvHuQ9m1jg6guQeUQTz04enqOKGmnjdu3SAdIp
GHkcgyj75fCiukpiVIAzkjJQGw9cY1cUGcNMzLVxhjPb8E8uiTRQEP8sCd0wM/+i
QUMrycTtsrO2UtBspixxL15ILvD+wqjW3NPnuZRel5BIZ94YUECCYjkcb1RbbNIE
utAoBbP8wt3fGWO3nAikTNEK+47ifB0js/2KBmZQ3d2gyeGeAS5QROlV6xDKZEba
0KTHV5zvHZ4B8rAFfupBh7VIMBrKOlkOvggpgKcG2gl3fTU2+tUgceGSArTW7jju
wPBtALqQsMyJxhOEVSgGhw1r/RHd2F8rukNHaWv2/5aBQhZlr645bpozxYGSqpzZ
Kb9tXQPK3neBEDHnDXiwpkfUqtqx1BeaMWpqhbQsv9DzLAH0u+wetyODWLBNnZPa
2A5A6OWo5SgsFTO7Vi1b3S4t7GU4O0UJVhohAgvDtOIS9Thglsu7iGQpo2qL/kaG
RZA93qThojfNdq/BkSlC3cK1dTtn8CieRC5vkYiHGh7c9Cwbvvc6MkNrTXQnN23E
m85znFtXcL+t5TxePivwUX8rSCqFM91azOVpTMIXLS7CIzR+hgl91ypBCm2TndXr
Le2e1Qp3TGYPH7L7VjUTBxlTuyoNNuPB4HoZZqPgZlh5Im6pQDxHvL6sHL5U1e7Q
Gz3lRBOwjUZzoK28zCMfRH/YFqxp1kWNlCSWBBhbBjQ+oIhoV7AkBrKvjj/7IFnt
1IHqq6cUMpXB1+2eR0yyISmVkcSAj0CxRu/x+bO1PDGOZCAm55k9cN1VW4d1wNcr
/Ls9WwP+QjgocfzPLK1e1qGbX0O0TP5uBsOz71BCRneRyVg5BihRCoRuyjOzGcUW
uROSFXdtnoWyMO22WKdO09gu0SS/MmvPv4UjYeO9WU3qRxtBCeN0l7drC0ljjTci
HVB02HFE9XZZhQACHYeLADF0KJvbEJ/mL7ZgP8zAXDGFEwrkytqOnC12RVQmn0rX
b5UO3huu85TMExywWIoI/GgcOtYFXd99CeUWiDspUf9m1mQWFhyKt+ocrGT7NszE
G0sTocWan5WTXyhIZXJzIlScWnDOPJWFY0c/jSSle38+tnn0T4QgcJ+j+yR4CyDZ
RLb/jB5WgATS5PpwzU4w0iY8WIfoi8EV6uInYxPIzA8/JeIfIJ8KbF1OoXCfnXMV
m4vNNvhWAAAoe3fTXriR/6sYIvX2Lh4vX6yj2A030/3zUqWdRVIjtGcLxsJur8r7
0JyT4hDsrmFex1vyyyzVAU1+KdovigQaonNmhcqiJMnUl86dfAbk+EhyjhqPtuLP
WyHrxZoREF/Fr23lktZjGZWro5S/nWOnErfcKHeOL5P753+rqslzHQrhQfp1pNgU
+S0boyeBjDulfdMcQ/BsSKPkDJQaC+NyciIUikNfmH9N8XF0X1Y6c8Qsghv7RvMK
amyih3aysPJf6Ex8bs0WFy5Lgxzbx702QGCOyq4S+QNkXoRX5fOEucQm63jzMjex
7VsRLvXtgRivRWmN0LZsv/Oz2XDgS1/RuIxBN5AUaWyvjLuX7BiMuHLAEcbd5+O9
ZsC/i1TwGj8Y83m8A2vE6FmkprD8/aIAK/9IPESFNhrm3dFSLovTImCjfXHhePy0
G8TJj3n+2RLS3Tqc/DOWhzYSQ3CNBepS8s2Q+FAZNnziqwY7aNZvZmsRSjRfHH2Y
QtmgN0vgApnPFqzT7fE7sEOjK7r7qCRYSVTMUcoBMBAwS4hHAl3O8R82IgAdi2YG
6/rXnjejUSdd8yGi6n+ORyWBw0PndKe63mhfmExZYdcVViPpuN5NL67J1IAuqp4f
qazGZ+9Gxna1mTR7Zeav9grHrBEzzEK4iCHt6Wu3L80z5UbCSk+BXOYIsjieLl5G
btfaEpe6j5xyfqaqfdtkK1KA2rPS9GIc1+2+2KlshGsi527me6Ccy86AZF2TGPXX
UTVIMunC8EZDK9d1lKX8cE43tXXfAHhYzQ722CIzfSaby+Fw9ghzX78e4N2F4Y8j
xUInnIKbCiPMxkleygj13/VWouuAhIb3GzALu1V64I2pX/JLmo6JUofFj3l+rRii
+VUOEMPNYWpPBKWDWzfO69SHH72SqisqYIsXIw4d09H8m+k8xkZYNn8xaU/ZPr6g
/0A1mWcwFIfgV5oq9yo8lHwHHLa2KMr2uLl8SfJv1BD/lp3a/O+JjM5Y1swwSfR/
WfQ3XSzuEjoRnmGBL0mLARTSx/ZjCuR9pzDqsiGhfLck8aNmrylyNEhP10aXdnc8
ZDm7bxH9a6RW14crPoC7g+KrVzCrubLtBwHev5Zq6CDLm30eS6cq6MPagCJ4Ykn/
itN9NpcIQ1pZmi5t3vRGk2LLIbbPEad223Uj/aMEOm/eYYLiKGLiRIJSgmxYnmUT
F8twdfgIuJdbIj2/aPgbUEmZ7d3uvco2Z/05+FvUcpcaUdNBAjIDhG4hmT221a46
H+Az9qj/y0pSrTggG+rzPDYEtf6Y4dir9TwCVueEUHNLPRRc/VK15qwxiH8f3yod
i9vvJjl7742aT0UuF4e5UGAD/aDT7iUGK1j5KSH7kLiks5reaEhZVIZuG/EITbIg
IlOKxMKAwOTTW3FZXNThudiXjSuBdAmFi82nmayAujWYLlEXR3NfUYcWy7deTXuM
MrNpvt/C7DpUIPMkrlKNN+L2YNJ9AgmPBLU3gwikmr4T3qi5uVja+xHMmSA4KE4I
oww3YNeEakFmNQkGBXf0fgVoOSU1hitN5wlCwaFyu8oKmMAqJE89PSV0yxavib95
HTESPqxujJ+KiXV+VBq1skC0qdaZ49p5xyGJzcRncH7xsfWNF0vPMWHGR+lEGQPW
l8nsDxu+tqj12Jwn9W8ccSln250Ia0g5yNSvtTJ011mPnSzNwvh4mjv5lmWu4qVv
ZXXdV/x2d2uQp/u8gkXmx1t/itCMCqmeEUTKNjDUgawJeNLmzIwZBSsT8ejnAsj6
QEGH0VUvOpJwtGHK/VYd1rO1YraVS1RZAjFl4upZN/t495+mijYM5RPvDRQXpeRi
J5I+1E7CakIrh/1Vz4V3yEtpvCxVunOnvM0TGOEuLOblE7lydWHv1KMyZAgGAK8I
oQe4QUn240Ur2ch0N0aE0pgrphyAsLX2RomDPBKAAUURscYtKgO7vXRjMzZOGGLZ
FCYhxaU39D8IpSxtwkbGV+PWfXJ03s9TjLPUsCHXOwUuxUH4cRpScSHwhLc/bwXJ
LBZn4rcVMhJBDHzaS7z5oZhi+djkwZ7b26OhXP/e1pX571mRmVIsWzfrucVLZuLy
melxrel+symrva2xHu/4/Vsc8Szha6fq3o86FsoXOdOFacynW+vYFcKmElkxCbDc
emlZ7M286N1RxR9x8juWZT0Jp5+fzRnvp+I3roZLlxzY3WhF1GgJMJOyAkAx8AeL
kH3ys9+SpA7Dx1RLr/AqMlZdJsRaRktmnld2DJjWGMGOiYd59qrR6qo6Snizfxhf
9hE/n0AwkL0biZ9bTosrdI1hpYyUwtI/wTJWMFNY2OkpskjIDsV19POPUi5FQSab
EbVMOKgZ8oaZWw9ZNO7tfCTHRlS7H7VOg1u/x/7hyvZ72H1z1o7VsuHlDrR9sJDa
npea/Sl/p2w/Op36voqpxT/ZsBOYIm0s6+7WG8mqneDk8fyV1BDV1R1+dEx8wX4q
TNnDqR7T0XIagncrsB6GV7gdEEU5tpE4lD9732paIZfxlIKYEmIUP33cn3Z+HoFy
IsSkk150BqqSjBFlpVEuQLPhRrdwSwzFtyC0UUz2Yzw1eLr+unRXWPlPyp3Tg1BQ
NRCv2Ur1783hB/Anqp0ytaRrlUFCTpuDSv5FspbiKkqB2fAg6MN0HZYtDtSxOo0t
4pAG4fmxGIkLJlaVsQc/KOdw/RXLYN4qh+H6LgUXrlHa8h7Rozs6w76CikaTiv6M
/Jd//w7h7NvACEBhkzRa28heAJip27a6rtEjFmwy/0ccPcuY6nbY0XeAFOiWgFVw
lrr+MO8bAXtOocjUTS/Sei/Cqu86Yr/DsCAIVSjgdZKG2aPkbMHahvRvDC98aeop
cMDKN8Ai3BGFmDEdgos/5/lDoHdR+T6HvqE4qrTCzyYhEvIy4yWOe7CrapCoEgZv
fgmxoUHG2k6Xau2YYlVfM0jPWOnp36oqWusr0p1OcGDrCsmC5610t8J2nvBj05Y0
0bUzF8fai4YbSz6X4c29jw5p+m2TzqLn08GMtRFh/ggPGjb2bzx/ZJfnHS+Qya99
IwCRUP5HXRit+ajHZpCQId6syA6yLou9AmWXRovF8ZYe8Pja1MlpBGfLMEpUgH1i
ISaFODYj/dGyjxfo3qGIDwXBAuNv+nw3UrlGMGIGjb5nZ05vXcn6hRrbdRGyRm+m
RDQ9p2v9X+kVoJ76RNgINhb1gUSyWSn++AmZVB0ykoFgTlKcqbliIYVHrNHX1qg+
S0lCV+2S0+DfArc61dEovEENypkeCriFzYjcdTBwqcpaQqXE/7Rb+OUG97V8qbUb
uiHuE5X6gDQpUWhQHZpbDyUVCo31wers1b71O52zzly5wEPToLU8npvc8Td95M9d
ibdr9fAOpqgoMXgJsMagBa92zcw6zT14sk0H2e6560GXb3oLV5dkqPwBNZsubTWq
lKNJ8zEWy3TU5PNTONCAm48IV7gZzVKHIcLxs0POXzweIgyJltQSwmD2//NNY62G
A6Zd4YvU1dv/0u81TuxlwqlUko+Vux91WIHGS25mC/UE23U9WUeVPd+LxszL5zoc
B6q3EwWqbveXKe3dmi9f/4Nvzm1xf3D/oW5vpHjW/La/HWVCYLksyt4tx1i2yk+u
ZHMCKEfoe8qb91KaEzSBb/BOXyy7uK+pe++NHyneLUjULNhdZaRQsMoHvJQdTjik
aoSOqDUSC1/e8LV698g5z3dJl0v0xyIM67wTNvgr69hevYakSlhx2ZwFXxdjHQ2j
lOCAmMysMLQfavVGfGQ+66DYZV5NWM4Gmyp398ToL0RLByCkx2U1U/j131wbB0U4
CH/njYskcXI6Es2RlJEQOnquvOUUJjIcAD54Y7aXSjHA4w5sD521Ybad+I5O9jzd
dhnM+zE84hwwusAK5ytkV0E5DOWGRvY5Acf/adiy9S9q6g+aYTlNtqTZGuBaL3pe
oU9iRhGNpGMYqa6WMRhBNkdAoBN3D3evIUm10w2I+3BT9/zfhhMObGNJkxH/UlTw
eTH93K+wqTHUnVZEMY/hvN5OIEstaS8PmNuorJdruvwAxvkWHteZIiRwzgr7KOj/
D4+R3diCfHlGJXEtBOJ7DAy3Zj3c7gSKZFgdVPL/G3Ryrq1qy2MFaTVVPd+b3ntJ
Vx9tnKohTYzFxU8jN9JnEQF0gUYMD8bHdfLea1Yzn/m5Q+NMF/LwjUxZ+YmR6gvE
yvgV23xqo9BbyHV2evf4t/2h5xef9gpoJCxnx16SPebB5t/chleblOoNWJtoS6pp
Z+jJSp1D/3UxYNQ7P8OcglXqvaqCJuU78l2K4Dl+YujHrCjT8QLx0PikvuRIxQaL
wakJObTtnCi4CTTFU3bPSKWPX37PAiqJGwNpeykfj2J73rnkXfADluzjk+qVSQvz
Zn5y+Ix9xyWR5vT+1LFWtQ4Mt1gtQkv/trQBEG2QIHo37SPPRw+HYPePcAGo4xU8
zk1elSw75XoA2WF6uUtkQT0QbmhujNgtC1QskkQdYz6NhfHqxbC0MJDgIyjZlzUc
X+cQPQdH7KPBVc54m0j2bhjBDZdDSysAui0a75mZZoGqT3CEnz/Us5Zmu+Wdgefe
Rxbdjz4U2MtvPsodUfHMDshW0l6EWndEJe9WEE4kwp0Tb+Gxhv0Ra8ZmoeiDEf9h
Q5EiUj2wdkdJLkCs55t5yaWiNJsiAMSkSD2L32cmaevjJcq3I3fJwrvipeg1xD+0
5/1mWL8QCHEHaGgYGYymdguhvPxVAzmcNLVACufVw04S+8vpCzL80CflMCxDDLYX
4x+soi5rr2wkFekUwwj3CJ7mc2cZN86m/gmeI6aWWFedmEGV0A0D5Z/+QtqKUYVC
IUR1WTpoXcmR7g5t+QBxJnEtK1qXgNS0tjAwt5zGEFbsqho34Btg6uTI+o1TunUb
CNU9KYnkYUXKU4NhCwfSmSKLUbhF31c9eeMEhBnfpOo5G+OnEExSLHO67ynr5k4C
3Cq3E3Sc9r0kJ6wsp9KRklBYEMmpJDhKBeFbJjsdf10RZ6drWZPlpkvtz2o1DGU4
Qh1GeDY7E/iQ5rDJuZ6dYlwlRN5gY8jIuL3+pmyPV4PtAy0y7J9JYALPrrg1+rsw
ohVyuG8u4K/qtTk79c0nTgf3ECgEM19h/EtMWC+WavcM6IXbO5cJ4averR4UE7uL
WBn6N+HYsjcuu4CmGCm75+BCnspvPNbrOHsREqrPcvOjArmy/9Xi4xPPmNB0N7y0
fZ9mVz4H7h22KdzEROOYtJMNJZ1slu19L67AOM913HNXbZxPS0kUPBVewaEbze7K
A5RDSnUf4uMpjo99XnUHauffOqepb68F6dK7pOkbmapzbiGODBCVAow7Z9LVDKzl
5URPh6981jw2Psjz3MoxUGchhoAx4acy/YIF5P41M+8UWHqOlaFnCY9d4s2z3bxq
E2d5LX/bmYixzMQdz7DhevBTtjObkY42tvsGIkSSQ5ZS+TrPRHG29lxtExECOaFk
ZxJ5ksyO4zfkjhQx1iO+OcXmANmGnsa4+8Pc7eNdnMghy4E00Vaj1dbg+N5wV5l2
OyIbuksNSiD5weUDfU+gdZ0C7X9w782BhmOW3JOrClwKxYGx24tTxObQNqSnazs+
dGBIbxX93kBusmqC5BPnqFT6pZFN+8qOvd5EuTgiFpXB3adQKXSxMPX5EwnRcNbQ
sp3Kgv1ArKFlh+MhB/k+Oq8fXO0QnScBGfOMlTSZUIYU3tLumnTQkohn5dNC40Q1
c6HjydkCtF2iJbdgfyUe4dPaPWOkr2gM77JMPs3NUpZTIivHzKFQTuAA5WE+JOGj
Pp4kBA3OL8XifHmBUr7JyMIgqCY1NNz6W/SsuQAWACY57HDiB2KmGSQEABxtKwvc
HqieJaofhvK6aybbv9a6BmMhNiM9nu0XYfdN9XDytaEtTwpn+ReaoMZoX4EA9At0
mo/4clgcT8LO1QaV96PX49g5ioHg6F1AyLGBR5TCh/A8tRU+7YM3aiFH3Bi2YrkQ
Vut8hGgYfcyopwneUG9KVf2RTP/pZhibHyX9RicuM4g1a24dAerkMtGh7jIQIpRn
z/x4+DmmX7DDyXjc9ZD2jM+SH7IUFRN8eU/LlcKmMaWL+XPiXENoe/PAg9tGW1Ov
xj66ohylCGhluwRfzmwjZoLMiHyEvtva9qA7UJgnJ9C4QHKkqiy5xxH5X42icUg5
C1QV5qJn7ZsEaWF9n2WHJoQ4uprmNJhUuQ9SYCvjXSJNHa7TqleVbJcRnhzGBi05
fVPV2KfjehgyD9iZL7lfEj9u8Zm4ICvOn6f492HNMYOTGnacDZg070T7os6bncAv
6DZkrt7hoP/CCpWOFdpFUpoZPEi1o298k9KIYHbTvig4d6+nyCPCo3TAL/x5Ij08
WA0FlpFz9K4rbyUXqzsjtCbVuzpyONcBinNBDaoUZmdWDZnZdf4hLfbAqGnvcf5a
KBRWA1s6w8/c7l1Im3E9Kz+eVmVHMmWxpGgFRJWI36rs060TYXIDUIvPrOKUABUV
7JfRIo/FCrqiKcaGyb0NeVTpHPjolzDx9Mf37QSS8KgXDZBAv9ioFxAlfTVUVQY/
XZpI8YL5sOAp4P60sbayo0xxZHaddrqeoNaSPjC6c3m8YQlF9ckp2wT46XXFt5I7
tlQKp4EQ1PYP16Tr4muGimwxS21vvkVbNuiB1PgbdC0dD3HRWDYTjERTMdmSHhyi
TqghnOtZxrOGW+67q6kDiQ4JDdER+Il3f2azwOqRfFuVJbkYuTWdtY8J+naZ5/Oa
QQyTDMZBUpgzkHZEa1RDfWh6girDLBYaqmsM2myiEzMEwNi9LYj5aulmyWA17V2D
FlLESecwj+ra4wZfikl6sta1qA5ZKJ+SsOCN2RfmTXVGBEuWunQ/sHzb57p0B8xP
IufXADY2OtMMyYaXw+w1qv6U/VyaTWHx6F76dITV7YLTL5fACAinRkyQwf/L2beh
rexZAZh2kggggFDFxRmfFVgve4LGOZEAlc44a6BI1uNJHg/fTqdl1roDyL/YdZvi
1SMoCzw+dXG2RiCq7N1zwiNlS22jGNvwqTI+WDcXUAR9AOFkZGL8qa3gAu8WKwJq
4BUjfRVEDRJrbxnAyKEngewRtUiqmZ8NiSviTooS62uVjsDOAeeBWKxqrtCzpN29
zxXA2U3sMuDNWGvZGo/DS6GeRAYPGre2+SEoo30axnBLLVuXNBovn+oZaegh/Fvr
b6qWRSFHk9LnFaQHmOyk6jLbYU+//djj/UQrRGZL5QdfRNg8WMvXls56NC2O2Erm
L6OQORam1Gz+Bq4osaGRmlr0jnW0SLsux/znvhXhZ3k01FnoA0kdWTNIMDqR0YBY
jFXaqozFMyU5tjK4Jae1z6tOCj7Iw0PZWAJENMYqAOmb9YGOZJmjJLOzof2o8dAm
oD8kYmyEmVmjIzjGe3XqhckUNO2XDoKKWHGnZ2f4gj5qNoEpoCtU68gH0pLvwJ2Z
Me1hLSmuR6myBP0z7Ksu4rk1+HZSEpzrR/jUVBITtRzzTlHVjr6C3mWPvMmWE7uS
0iFqhpGu7sMv++YrBt79UFqluEuvYRXaEqyaL1pnRsu8iTnfZzGl2e71fiL3MgbI
hIXLk0pH0u2lmC+s3TCkldR8BwzBScXL5ZXYIsDM7tR76K1Z2R2gRFS3MzNnAVCK
+TxEvFri81o5n4D6Hnj6fgCkAn6Q8ZbynuFrhFdpwEzwKDmV+PG9ftxTsjjj4aFK
MITTI7GqZzZtMzz9Ai2uLELgJ9xV9qe/MLI0AA706U69tFLmQV1VehBLjSjYm+cz
YvfxtlN6o2JC9cnuaSgA+tDO2uQRJTH81GFukAkMeh5AlRSSTyCYndS1wy8Vrd6X
qJTLR+x6lcQvq38B3v42MPhUHfahBubeP50xylY4SxrYYf+gT04O4/yLT0O8xnoT
xCEgBNA7fivpSq0ji2rmSMM7X7Vvu0vQkEhJrExW3Q3MClB12EXXj9va7ILnFWbe
pgWCKDXH9e52XjdvwpdHs8zUUCZVS1X/g8N14H9utml7sZMBHEBUcnWQaEfNTcIj
I5DBjihC4e69fU1xnE+JBgYyIk01EQFG2O3cqXcvmIXbL2E3hjonzqykptt/Nb2t
XztBdOECQ/8HYiXyO66qmLz7xSKukkgzDeajrtJFZ3R6nUMXE6oqxOdthiMrJ+Ck
Lp9QXI2MOBAVA3d/pCMba8qpa83xd3BbA1T7dfr2moZfhOWGtrkBhelEiwoDeK0Y
W2W0hUt2/Q3W0FmJ1dzv9hT6gW03XtoPgVtrJObnueeJg7gnWY7IzaqnczD6u21e
zRMFA8b+6iyXaG/fBW842RuNKw5DBL1WLJCQrktCzMeR2fvuRl0s1TISCYEbXqm9
nYWo6zLwCaO7QiTTNG42Mu0SKxsMRzqNBfuvanqZQCPDfbVkavDJHJQ5heMDbOh8
MF5LQeuI43+aClcGR4RnHKol8Kv84lBjxqGWBu/iZZG9m+hBnNwHe4EhbjtBHVwX
cLcBnSVHkMxhyBQ0FDWON/JOedlnhZVd7KL2NlIY4OAygjQvo5oO+ZSxO4q0eHvZ
mKV2uErs4XKKu8NPgWI7vJCe1Af9N1Qh8d2JmpEUva5e4eAQ4FIEKBqzJPzGSFCa
6pWg+xNZSXNJvket4nOO64i3C3vDVCQZmPDegv6D/0Bro2sbxsR2NNeh1qbU+ZVC
wUGIXR+BMMYkT1HRYUly3auulDWud3EdQyAUGodkmNYAn5DTTRnzFBCfTES1lyaY
tG0yACJnTIN3/c5f3ywE/jEwyXAPyag5iUciV2MOBWWZNgOU+392gGmwziVYLzNr
Q5AnyuXRgkCMbo8Xp3KmoSUW1BEJTkfDiCDzHI1HW6ieLMBztv+pR7OQDNwe59xs
t/bkvBPucPLrl3T84IWF4/D9SVymrurgCtRC3c5SWTBOcKr9tPah+UL+8JOEKl5Y
dqUwh5uvaePMpAFIAnHnd2gEUatEaE3dlhdO8dM0vUGpDxw5E3F5SuD/6ZW1gSwG
FP/oeQm3DKQLrZwto4afc0ewxhMffEH+Mkry3YceH1nO+LcE/bQU+8P4w6E+upep
0VULpYXaJrnXLOStUcO35jPrOAAqK+2yejeXBMrQGCyDdFk2H9vH3yZbPEufZ/7a
wp+pkwsvkvUDScf0JzKkkuxZOFi2VZJzGR5RT77/z36sVcICKaB9YTjUs3p5rKT4
BzLIN05E+w4igPM4JiBlVwowP8dhB3TDQZT3B6lpDcDh/o9VTKmpuA45baPyzoCU
Mw8qprgscGMii/a2/7ePnp2qPzWH4pHVbESqkYeL1PBrG2+5WStSsdt7oHSYbslq
mGx9Suklhkjwt1FoiNggFaEQt7gnhNBKH1DY0tsvUcqT0yq8wV8B2zLRuQIYQj9F
8RuPq3K8YP7wL/7oIH1WQWzMl2v9sBMsgrWEhmACyFdGTAzhSdOurSy73ZFkkAxT
TEiFW6ItJGQ/NYemARTCcweivEudNGLyEhRJmGCSwiA820TXeMNX61Gi7yxSDqb3
OWmGQrCMO7864SRhIQ7O9sZubwA7CsoWhxMqjIgefWz4B1xVxUQaze/mAK0XpuJO
rczgiO9i7srPiwcfhbg67qcR921fhE4q7f0UuQ2BaTpvo+GtEzyRs7OI0wcMuFg2
aLcySKbaAem5VCTcDhuswCmk40C4ycAFxntzjexYznxj8PWYIaA2FAvXpmJs6GpU
YM0ms2jOg6PYKmh64hiSS1lZzA3v5a/9k7B4mKQZ8un7K4bTuwGXhoO14Yuelxu0
afJvetcCIXchu63gr6zPgTqLeY5+rXqBEKu02bIlATSRAKuBaAMZkWzwXJUXyBCl
xJVe8kqqM34LGJa+44eOR7OFHaD3GGRvjBMXy/25W6+lnTcBtrgefVbwzRDpfCot
QNFTy/HkdYegEkTmvPIxtEfBNgv0DH9AapDxZPW90UEUBodllxpOwINh/csJrkhK
ORHYMfufTUBZy0uzxaA5CYnIBeyz9XcdD6xVKh+vsD/rPNINkOkYgx0+1RCRHP0G
q1IM8IjNbaEB7+/ZWl1m6MpsAbqL8GY3XqXnmA3O1ZDGjPLXZzokLYmsOnLJRn2P
CjG1JNjn4ZTeV2AOREgY+fq0+8yMHIJdY5xwj2LZspY4rUJSsvTDPYQxC0k+tDpk
dtGgxsyrY1e2ukuDov2AA8wU0B/iggC70fP7T0kUi87kD8LgfGy/A4UuYwplyYC8
/E2pInTnhINrSn6pB6PyqoSjyHgoCFv6ghi//IgrBsPfC/hw++f+Q2wSbot7KOHQ
KFGlzd7cLT8kytRCquxbs3j+fmy+U3GSCr2fashs1tAz+bPTDTdvfmVYjk5LMDe0
gQ4Dtpb0TRo/Coz48g7vqwlDhc5dABlWRDkxEbmqcNl494F3fhQeMNRgvMt7Wd5t
RZbgjItwhm8obeWG7wlky2MaYKfq0nZ5BtCg5TjynQ47stR1SHt4OrN2dh/6GhUg
JxpDuM/hz9zzaW5cXZTVAEaM4KbBMr5GCP69tiYQ8BefASEnm+3IS68022iQ1Siu
xLalshKxUr1g5JnGsIJ6QyHkz3DcMFQCxJeAF5OWOgue2Yg/Enh+XMSOx8zh0cBU
KLi4cZA5wcUCM5tIb5ESiMqh0JRnFcRYE702JJt6sNC8RofFWaZH6sxQBl4oca9P
0i/2pB9u0jOVRc+i04tSty66UOWM9ibE6gu/pEf7I7XPlNu3zUXkbYQU51C07Ep7
eDgv4XKl72z7CNJ2rGbdxT4IxIFJbnEsDnVNeaIu6N2eedcNjoljI70o2TeF2fuP
ZUTIS89x46ie0imSSl2p03JLtwgueUeehU082p8TH2BBCI7wpmESnI6Gkifqpdc/
baacgjCypvs4UZmLgK4IioAkIlb4+qNLdlRVmtiy/ookbGag7MrJUOsLO6xQG3Ms
xHw1ZrzN3vsgqLHs8vGKnKLbdpurEIO2ukO/PulAGuZivrPV2ttO81Bv26ycwwtS
jOstp/Biy+N6qpsztzcwpe2y0ZBB4f+zQcgbUvlAYvM5a6K0t/B1mK32L51ZzGWC
79k1OnP9dUzWnd5Tz7abrraHInpWiB+mjM6RmikLDrCP5RObtB0EAZM83Nze6gCy
TR1aqRJ6DhRyhCQ6U2ahcJestBpLQ+x7m+OrVcMUzMfMvk+nEBqdY3jRyNrrIo5W
x5Q4SVGHxxYvpQsV+Y9olSLqGRfweCDT6MUM5tAfmtWv4YT6xMajJskN8CtSTa0R
RoOnGgpv3AOQReXoG4q+xIOQ2qdFExJ2/Loieco2rt+811UvgixjnIYS+HmCUmE9
+mwlT4EmOSMdOZoiWlMaulnAH8Va73v/2yAG5i4Z5p00Zq9luyxbylJMg1H1F8Xs
roZWk0AvMMjQS9IISsjBegx6DBRtiETr1l8/12W5VSjYfPN3GAu126XxyonYYcdL
jVOauScBbKOutXdAmdITf6nM+uUWoghZ775h0xMK4ckY+UbI/vEzjaUcnE+MHU2k
aAWrxYU3cJ671ncnYadwj8DxGs2PDMj+RiAw2Y/Fy9bWFKzjeWcpG6xh3sB8y/LF
e6gIovD0f1QD9uxFCQYAvqTNYbDvZEjmFvwl0iCZJwetNDZtITU7KlSzhegqkutM
VzutiFpPUjsu0AYq53UnAcPQfErStVVC0cZTQVOufWm+K+J6Al/bom2NLHoWocTB
x6pHP9yYX7zTTum0lYiH4/w9p3hSCFb9cxFm/NELh14ocRdrrk+KYtE3hq7romfS
nuUKq7gaAZ8VgftWDNXy6PKlrEOSJyNuPgH18mfhDpIx54kcRGFuahhZWGIGsntX
WwBQ3aLktDmbT8VNxu49HD7WveQfl4UkOX8jLR1K33Xooc1a35EScPouBlPu56/D
OTRdpiR0KO+QWpWhNkDXnqLH1aRhFhSed3kdSXOsVee8HC3uvVY+BM6s0p5V2oii
pG3BacnI1L4dRH1qR/1VPMiMI+m4QzaFWzicBs8juUTl5TE6fnilXke1B0wvU8A9
evj1V1lSsyzpgp0Cjry2jgYZhhSAXdEg5OUClMH8SeaPqvUOu7J9vSg4SJe2i1/Z
NnQFk2nrCJbbh8/oiHxMNT9nv69wX9MbNwOsjsGFmMZp4KbGoUUSOHF6Wi8h6E1n
e1r5VLpbsH4oYPF41OaZn1Is2J0Z0kpz7pzwsbOXV8P+YGlVkuv0NOrrFpWbEou6
tckSKPwP/MqvZb6pGJCEVC/Pmcm1V8KkHeUXNwWuH9ySTLpXMu3LPZYRgVWZ5tzb
CFXvyCMj00aQS22zMknA1ff8ng2hob6PLY2APYha58m0hLLXc0AXFedn5vuaHLZW
r7xHJcKkxr9eVTf95w+Jd417sNL8Xfwdotyp29xVsH5UolFwUVvxoKCnzL0VuTpR
tQpqfjCmCjvegB7ORwsHplY5CEcXkCAdlIYAXyakdqBjWBz1jBxGsBuk+KOi+fb0
IdbDe0sMRwJwtgNgiep0mrp5pJg60Zw8eMzUfxoOFp9JojxG0StTrL3LH6903Rca
+8kelJQlczvwx9lg0Gz5KzfJnm/XdzD4oDYidlFoYEBIR8ohEhr5uTo+Yn4NMc6I
3u2k17m2vkzErRkF7FRqzj4lDwhOg6x+RnoIzqtqAtqilgIa7/E0XpLJcs5tq9Mh
CEEe2cnZ983JEUxF1mQycS9xEcEImgYFGbPRmTLFEAH/oxK7oKC5n0ETt9Et8xE0
ObFq2ol4wqCh+9ZdWB8Y4kVLueDzkqMd5fZadxgWIiyp5OiIRNQvWCC0S1CAQUHv
1fLEHpyop+Y46CETZdtPGpeF4oG/WZ4sU1zHURJwrmhU85zzl2cpk6fmNKnK5f4I
uejKOWfOB23h3KLqga1adgeeuJEjRL5HiHoLdK5IxYSVWuqkH5HpxFVN3tPJW7t5
g/CxHbpBArL9F8PEa0IArAl1HIHV1l3Lf6T3O19z84iWj2Ze0HpTtVIA0vbUGmKR
ZAAkulsb/V8damFY8EURpFJwZROPGgrK+PNx1JpP+gyOi/8M4AGkeEjjnXnSv72g
1xPu95eQYgNAa6/KUHv0GH9DoN25qqtygPSLu4bnwiDVPbVTg6x48kO2an+dWn7h
LtcgbLvMaXMx8G8Nw/iQbrWA1w+FRLi2bbRtBKH9c9nWNhyjyOIAXLtNWj+QpDMQ
hkXB3HiBVCqzejzfqpFItBDTaeGjKP0Yk5upQ8THwDuMT9OFGK3Od/3szv4794tj
pjBrzBtzo4Qu7o92bd3qtmh1xlQ6mb9u9wxH29hK7ndNSg8hEml9n6mgwV8uQT+E
O44Ae3nGZ1pDivmCdQt1/8LPokq74UOuWWB19OZIjuGzc0QTef6YdksCZiA0Ele1
Fkmkty/6ypuyKqOMCpckoaY99KAcsLseegbBxTTkFWpToApguov/vM3pLXzFWGgQ
kC7wCqlHyv4tT71kSbOWigbXhozdjaebjchFvBqyLRc02aIe+oMKSmTLmRFFJdXk
5cds7eOcKEz6F1CP64RWchriBOG80s3utw2C9t7fTXUUi5A6I7jJ0/VpyZ8siBxZ
XBpwhB1UHlna/OIuRXT+kOzzie6FOGR7YKO9f/rTUWA/cZEZ/Fr4Dsr+DTdMTpnZ
WUEM/GMlW4Uf7QVkzJeZYIqdfb6th+dO5RefK+QaQnw9PR5qwpQxnIBmEoB0Pm9c
bAF3kg7w99mPxXpFUY8hlTqCuNYl9Ic44o3EtEvefudTqYhHRXeFSUKksPqW/h6G
1y37xV1/Ssespmz+UYI9EwPpHjKutkHC2rub6L0zdiFqQbltXSnUQUeQhq4vUQK3
hj6GIbN7d2WLf2MzuJiu1pdPtNXpMK3QMjl6maOLRHvX851oc2YpYyjsGaD3r/Hw
D/qqSX6s0rT2l754tKHa2zvHSGS8PoGz1g49kxeOzYbQd1Y8mln2KoHyOai5nDcv
Q1eEyIz9et2E5+ycPMDd+T6ptD9lUrle0F4TgFvakfYhJYWDrq6/vPjBjNZLZImn
Oq4/wXrgKFnjcvLDXRk6fR7Jxb1CCptzTY1qH+4B1k47hXlEuak8g31WwFepw158
cVilgRcDM4UuD1LKActy+B51h72MlAE+nzjfP9udXpVTvM07SeE9W3E7p3r7wvow
L0tVyTw8u5uBByJZj262EnZGDL226D+tsYMg/BYP4Bjdjw/OI08Fnus9Nq0DUMq/
QxOFeXmBOVJHZYN/lX+ByJBm/+NZOegq7xYuHk3S0y0p5tIt+NorhVY1xbxTyhBg
moVUW5Xj+f6Jjd/OV2BMEQ7Zn1EkdDzWWjm1aZz4TdDI+C2Q8xuFDRMbEcBKFqPw
hPUr9NaurueR47+tKxg8q1MAD/T9ojPxJJDSSwstqg9wXxy3eNBcxpJOwiU5v2lU
BII6kFGGl7OQ1Drw3shNIIG6jtb71kyHHw8uwCxAq1oUot8vWf1daVIhgbzUvfus
uFFdPZr2o0SK0b9lyn99kSfc79wi5ZoWejpzD3As3DBY7Y4wl1ahBJSF2mnIkhMz
3dpwoniyyx21S3ZoYc4L4OpyVz4E+9zZrgnsfoTaZfCoPK/QgHh3Dtg8RhFkRWan
47zaCy3tW5oVUW3VkvC5UFMYXA6P2xLpqenqXxpwvDqz74/dYFeJmw7UknREnHV6
nkZItRo9IzhRiqKXAIdz1zAH4GROHIhKUSvrpL3zeH51lxZ7fR/LhIJK51dhNpm0
QB1qpq34RPg6bXZ3NpU6A7stf2AVllY0w5hK5sjdPk+5XwOLcYYHYb0PCHPjaPWL
Ai9L3+JuDnx0znWN5tXprrfY/0ZFyMI/b8HLl73p7qaCJMPSoXNL6WQzuXcy8Qk5
dUzYh67ZVechjl+zumiBbBk05ywmymAWzLNkSF5VNy+AziTJufkdZc+6IXeJiMEK
1OeFVLAVkVNq9UwnVNIbAaSbI1kb3tBD0jmdwXakrfkGk60jxP3hnaXKC5fBqb1t
HqvESsPWkf2NbVv+DYM75CPW9Y+x+GYHQ00YSNC1XZ1Nr8jcjf4ETo2BZhouZK1/
jmOxgYpl1BHpL9v1IjbeVb9otR+Ysz1OQ74TjL0VJLmVjveRfxw6KhMKPYiu0Mgk
bVUMYAV6TM3gA09GoGTHkMnCyC/SMLlaVR0CmlUd50z3CHoWa8o3uMQLYkFykKCp
ANyUKzGmD3UmzP5tjQv3gF63qMwVgHq5NZhXhgzEcVAdseu6tQ/ZIq0yKW+svDkJ
6VNz9BNu1ffv9n9yQZ7xtTiOmK13UkWipXAQZ2BSCZxmyQWlXAtPUf4m6vQ3LCYF
xZgNHCHiig6hDI0USHA1zzKxlx4XNZJtGWQNjQiFKNLdLUt2SM1NyXPz6+FnXfnk
lypM6u7RFMRwgMaQbOAGbQ6XQVvs5UwrgmRaSEhchLKi4WacXcRTDViTQ3rd3tLY
WnTLk27cpcFINYSsre//iAmzysJW5wyrZav2gXT81JyY7v6ilP0bsEBkihoQGBXa
lbBuFYvSJgEHxnV46PPXibF90lCfyqBkSOgeHrO7WU38zkGCYIGFmdExdoj4QCSS
J/bPHlCdu4spwU8fb7RnFoESyKu0JJJWz+vuGdWg/yzPUOmcQhlK12tzSlEZ5+2l
PHfTJ2RZZmcMRRMT2CXcVEiGfrceNdgGFVqYLsyy8mfOdBYWY88tFdPUmtsu/Ezb
zjlXHChzipr/6fI40Erw4+IQEzWCdgWDgXfwefDWKK65iDc7sQcCcbLaozL4HMuQ
m2CA9LOwjtvA9UJ8Rxdv/3iSqhZTCTSbiXW/dqoh945QX18EhuNJ4fFXwGnBA7sa
lfNPUz/cRhaheDsxqNYWFc6N4PSXLZAk8bzd0XmBx0SOj6zsavkzMcDEV3keziEc
4iL1yRhOuPyHOTv4WmjTPgL9jX6rHIFeOMmQHq06T6X6yqiFihKWozP/bDVlRt/6
iijGyDL/fgfp0WEPMrhOIisVPi/7akXk4x4kBxb0SsjkeCkX39X4h/AwC0BVc48c
rBW70BRio6wSjNBk9+new/gf469C79oQaqQoeTTs7bPVl9JG7BApzF7VY3bJL5hr
0JcI8SkqPgvbSvlsxkzU3mdwd5Vcqj4h0gZfGvQjQLVdAkG9rji7eXM+yZLoGVn9
vUywKd9vPc/5kVCn1aZvmQP40QFQXR6yYGqQFPmQb+1OGv9K09YoktPI1qOuVIP0
QhG3pauZDpp6kG1Jnbd7J+TzmM5ez7jlzBDNbLTT9+XalMEQyme7fVLEPiMZ+9wD
FMFwPP3P5XmdD4A0IYqBrVKUUGfSzLIF9UGxB71MZ9xmjeQ5vlCsHH8kyztPgqIk
6u5r+jM3OiLLBqpJHRlCxsaJdwizm/wimQvA7qfHJbAQP0OLJiS9qdpw3jfi8PCy
ub4PLHDLN994nN11iG0E88wv5iXS2LI7OS3rmBGcKFw1NNVzNpmSgqJygGrkOPET
3fJnzSfXkikS8VFkx0Tv3AvoG/FCS4PRTbD4+itH9Iuzfum/p1H5LE6h5uTASIZf
H2HDoDRAbn+OpW2eTwslRVn4TsayqutExK2mpPLanSnFZKU9wCEjRk+ua/fovSbR
8StTh1s+2gYAoT79wJtGKEiCougLPORfUBXOBcJiWUYfHNY9XLIbLqFzjU7/yEA5
KAQX2YethpNENEWQJkkYDDullBf+76o2xJvMx+cHn+K6arFcIJdOFoV6JwGY80EH
BUzyNEpvIAphuIrY0pLhcr2TbnqBVCrjo/LhJgv6F2n4i3OjHR4UZT8Bj4ORX3vk
Q+f0luupni1v4KoadthvTuUjYgtXvd+5/GOShgfyyUX3H8Zy9thsZFP/crruqPAW
1j8ZSgoRsh2kQwh9oknIGl6hydbc1m192KqCXKN++sx49un1+DPKhLF2KcSfB4Eb
5rPvhhVwNsKqVWddb8qHd3MLiwXSaNXChBVpNudxh7k1E9fN6hcx5+8eRYV2lzuA
uRJ0cl4hcjMxiQnl2Mb1CqM1QujhHgsNEjtNo/10WckRYlBGMHYUbtxwLtR85N14
QnhoPFvS4Sgjxd26wmbtZ67omgTB8f5c/Uju5rR6ynxuPOSu+8GNGtJEjRL9yDhz
ufzbhzyuUftvEQ1nf3j6SyIKMzYuZ6DJsXLbds7fomIg5XvY204QsMjiJ9QqMOJe
hMSxg6R+BBkQK5clJtubQImv9AgKhSDxlGMEKg3QuabgZZJssOWG66MW/4lfBWi0
DY8NXDBkfo4MECVfzyH8GaE1NkXsUd59m7xI2U36oUTiIdri8wgBsWqn1PeuJnVZ
hFWmmR2p6qFVRyGZDIm4o2+87AGFjXSFmMaN7YVmE3/PkVF56iL7VmD3jvkJoxcy
YU3Okd8ih4shYKRcc3JcZLDzY97fw5eHZA+hPVB6MeXqFiFXS77/mNqAa18mByvZ
EYtLOjGSlN1pGbEG3DKuS9wBsr3gag7Vy/BrXdjFuvWZkvG4R0aalKrsCdRTTfzI
K/CW4Ob+clv/NpRnkIG3VZOKPM7gRAxzkmq+IhjJvY/MM4DOdi5Mmaqfqumw9rr3
plWoy+k2WlF9KBV3ezr1TMJnej6f0BiLWqqpm6Iwi+Ds10R5AQxVSN6lYBSW15LG
PpQSV1T9ITexDuNj1p3jbNftASt2nA9HpqIPIoCdGhxn2m3X4bA35tb7EZTDSK6J
bfrDMDRgEySr34RoQE1Ye7lY2ZBruX2uVmeCblXMEUHpD9vt/OC5pa/DD2UMh75I
JfY3xjSm1nNW97k+gmKOlFzMwHWk6fMLirG85XVC/bHQN/i1LHmfIf37/2Ep5W6T
zsuivhlYd2+ARh/SQ9TGirr2ftyVqjwBAGJPoWgIwuqZZlWlZTQ0u90z5CDCj5Ci
74yg0JWAS/TWStmRsBwW67u0jQGo23XRmEOK/1cAnA6rQQJsF2734e3KdObEiiO/
yCOiwF0wcpQle2WHhxTy7L1qehQW54hkFH0zgmwaTZOf96jcc3XkQ0PHu7E1yIsG
d9CfbKZcqCKVWvoToe1NzNsbWxonXdvTbu+1RI44ekiSAIFUmAxLzjCQVPpQquO9
xmKEgyyYVyiuq4dy+D+Sv2Uh3refFzoHIMWm7CSsPahigs6TgLH88E9F5EitODVf
0Ry72ezytb40L/cx0z1mIa7C1LtHKTmF7yLgJ6suCiTERUqmtdx5eZ/co6yZKNM1
HtsKxeR/CsL5G7iZo7SFOvoWnpEQ3RrB7r5nDhcVZgUbhvYXgdWZIawtLUEgS2zF
QM1+h10+tqI75FkYhkzZITTB/+6Qi/OGFyxWxyZIhK5t8g02FXEKRqZbHOV1Xlif
Ndc3zk/HC81gzlF7Mlq0OGLP4X7HcWbX2bE8CZx6rI0aSeDkSUVP1ohim/4yzzKI
Bzu+QrOe4EKirv7hZ8n+b7mAFG/rrC8gRTm3/3pkFlXee998Lybg1xTqc+KsbsfQ
l/01/04/0SkgR2my7s5lPhr8KhaVOeIys12RVKwHOiRhGRfFU8CR3plLRb9jyZiC
CessQ6MRS0tpu57028m7/+jVADJ++iriJftRSVeyf8nTemQUUY0XBr4n4+4T/Jlm
5nkCqV2wADG0rBU2wbxEsPkB3gefwhrBLbUrM7Ixm1DFM7TTS7m2rLWXiZkgTmUK
FIomdWCqZyiTekmgyVsMbvLHQSlkGvIlkiuLTgR3lMYp1/o75lVTY53ZaV/Aqrlm
C12zgHxBh72UQt4fmV8mC7BN7G/OEtgL+l67UzYTeWgLj7+HzSsc4UilbWhHgBR+
BbaNV+vMRxEAbnvrDrn83Eo4vjuBcVkBKP8572Wa/Z00DHhyg/C3vWy5V+SNu73x
hAFQuFYlG6ExLQryxNz0NeAjkexAhepBf2HWgVHa4u9iZNFzuzU6aLA0yWIWD5bm
HPH95CSfBTI5GzhW+fhfQmHBt5DZj21+5Xu1kZSuJ8eCDxVxAaY9ohhWj4Mm5EfC
53KiBMdCZD04Pfq+l+tEjnDPHrkaJ7lDjYKLW5NAH0mE0NKoxMfhjXV/wL1gOjlY
l9hTQalUrf9M7+eWfD+oV6DMlyzvMWYJsgFvFZmdYIvO+2tCX+KmSbwjy/JNVxw/
Rh+Itw5I6QahgdbdNT+JTEjiw6XDb/Rf/wRvvei4EpeBdYiu6WndhT4UAunea5xX
LeCsSAdHNE3xHT2dcVLfsTE0P5oirbA7+AXLOckg7blmFxYzl1w1Rj64yDBFTlpg
wDmsBRXyq5ezhJmkZbne942M81XJqzKsn1pVwtEolRg91vi98v7Xo/VwujjL5Bk1
rXA8NtY6R2hKURAekTfMim8KNTJl78HSz9wmpR3xt/MnCV8B4wcLE7YbfM9k5+lk
EVeUUQ56260B7/w6AZr8Lk0eIZSwL46LGWPXEauOZDfDOz8BLZNJfLgWWwfd1Cwk
Et9YPuFuWASHJI+qziYryIpNzxxYESg07BQnq7CbDRHAmJnVIE/j6GF/FjTkbhmG
UGGGDRe8bfnkZOWymtxGr4h01aLKhF9MqzSJN5cgfTDYXW2kaveaxiIkLwMBu/GQ
20eXi3AERmTozzRFJp+T6DYzQpOuABq7roMlUNXc3Xchna8QRaDMg3bHYbSUbiNR
hGFIvcT/agmOdYJKRPQnElctn6PdJAHyvkyrsxzSd6GKU9x59byGI83wcjxDr5h9
Er1Bjn7MAJ68KNonmc37p9sfucmqcpx69EeKiFDTinEp1ru/rs8fP1SZ3i7+lJKJ
1vFlftHxpl3wBVH1eDFj8znNMGN6+irGIZzstkVzFbrmxGZeF8oXz3PjnGDWfycU
4T3MQFX3peJxKvUSlsYYbp8CkPA3PTqtG6O9Nasm2Dr492Z1k1f1PgDNK5HjKdcl
HCpA6cHEJYubgrhsVuQ8oiob9ybBV5lOUei2t+WgpXZULZcllN/MsVGXlBBDXhBi
pw8OMyH0NzEiUd3I615Vh+qLlo4VzIGxpLKkZ4wn5kWJeBKUvNW4NxyO4I2K6HUy
hG6jypiLPIZ4TVjYxU1mahKcI0u+FiOT2vR90kbfeyz/aIijam7gNuyKx69TziyT
j8A3+fhocegGu3yI49gcZWpFzKeINibUA5k30hMb+flJW36ZhMxxFJzUfvzMe0jo
IyAY3OmicVPIqnkWFHwmp1wkmty/FGrE4hIsfAUEEKsd1SH1jxZagG+5hWdmIoUa
u9enshDkdbVy+F6knXhpfxD5xd+z0dDgaJTn7cSIh52CHgI+L7iV9mrtfiv9owbO
znyshxdeaYfgRz6uWjpNKPH9b8kUO71zD9XacPG2kGd7ZZsSjtZg/l0HjoZ3bDsN
psIqVgJ/lTFmn+0b/5E/iNSoyEvo71c+eW94B1QLj3YDc/Zpkf84mz+qaA5Ck3pQ
1TG7WU1o0CvaPtqz/hvo6H4R2Uta7Aptbabo+XSoghbf3UNLVOUmT5VruS5H7sz9
xxqiL0PeGVZVDsRj7cu/wUlugiAg2q6/+6pP+gsH6kVy5MpmxubtJApinWfU+rXj
X4UENZJKOk7wUCIQvpHkJqMtq+IHuu4NP7qpIHzu4AN6G0/67VF1TA1xKinedxnJ
SuAazUzkmiWqgqIramzpNdIh0822QSCWYCVyrZsq4WTTXJDS73yp+MK2+B3UydBt
D8stDdxdgLUHzbzd/d8Y+heoxZunUJ31Yet28MqeIqMPg2ww0iQ9ygKWdHc+Vx9G
STyEEPKUOIfyAJig16xHPP99my6m+Sz4FezGCd85yn6RJKHeKuaSEuiqgYhiEyqW
E0HawgU0krN/XbsE32hMB0XddNgqZyV7swO4NxbxfPndA6h1xzmMON3CVdtxiypp
yW8RNhrQp4vfSRLipihEYHzcRABFTqVnYmg2ibvkMyp/mgMvHE1mJf9Az4Xpfuax
2YRJ4bJOZ4RIQJraEewa3OlhF/0jJAExaK/l+KFTj9VlZo3l8CnuKJDDw+ewNODG
mQOLPAQSbqO2d2NdzG/xjkdxP4x+v5B4fLBaI1jVq3uuS0APXdFYZrKARS1cFge/
+TqL4nA84MGDV0xDwd8AcGQU13oMnl78JxY60lJDezg9KxzVL9wQBlIUR95zTNaF
tIyM1/7RfAF2BogCJX/dT1XgN+aI8BdEHYz4VRs58MB9CzTCMwJqWwmtgDwpnz06
WTwhhgxpmPss5B8u8cCMn3OZYpakInVDM4S7Iwz0nyib8ulTGpFOW2v4fiABXzmW
0ZJv6TBeIMM16OZC8s1Bj/z9zlWSCzbsPmgNaR/Vy2cCZFwfC9uajFU1nL4jmtra
nJcUQhO8M+4KdJ6c0OGX9F9IHVQOUYvZi9+5XHt2y/LvSQ+mUIVcJ1pUCGA91REU
WpFMgBJv+uz93+anL95poO/X4ROCCIBlBCf3V/YOR9VTZAZ4M2GN4AmW6S6LpGv8
XM5iPetozKP6pV4zH+k0y7uJN8NGL2OuxH+iBSPpLENAb0paLkljeuPQQz4B0ntA
Lnr6Jbx32gr8Q1kdc/qRhFaRKOahf0uHB3NackvqGxwhuaOt13ZcCRD8tBStt9b2
0rw6+J8zYSFBqiupUQ8U9d7VseR0IZdM0gzL6fWl0sQ9ztAp0alVxAVJERIvovX+
3rQ0+zkCyfPcB3nds5q2zw5dcoL80/z2Bbwi19eF7XZUR407eGsmX1z+98jAjnwy
ZnLSJCTIEDFzGctBe9bZI/iY1Mix/5YDjYjb0xKKD3w2orvXM8eVNxNhJYLwaVLY
Mp11eJYFRYq4txJYNJa41DD+yVhEEysMLvjF83UhrkefhuBqD0BplFXocRQ4UtvA
ZMsTLs+ESUX9wrmsIweNTRPrYJhsrnrim6XHyJybzcKCHmaa8QW2/0OYMU4FMyHr
fbvPV+EbmbuA8KtqSmNclqitPUxeqi64GBHvp0GjnGjdLiP1iRhsEKgzJ2xiFa9t
r5+h26+1JjwTOkzCFgB9xSr3Yv9GZER9aiQnV7/7ZHMMTmYC8cY3QdptyOmBLDN+
2r7xDpHdvtjJoaB6x3m7wBVtr7D0+Lq+1Gjxnx5TSmYTfAzzNcjPwLsN7lgqsT8a
Gjdvn58i5p1L8RknsLbr2vrc+7mHgUQ6BRI0u1aVzjJqB9BwIzGYf3om7W7FLoCc
+5TKs7JbAqhISVLW+tCEfGD+xhWDLpnLGRkkaTXMeL8yJ/PSxqFbn239TWQkkAP4
p34i1YMKKHYnouEWz9jahYNfFUpzB8w20gNkp4ty2X13ozFyzwHpjodBvs5JzVGA
4NRHEbMOUPn1tNzjRq07IVWfLiqXobqFPYIBtyr+1F7ZXT1+f2mDt3Dsizubb0ij
k+YBid5I56x2HaOLyL9yUe7cwrk02cjeMSaCm8FCXToPGyp9xhwZTFYUXPDVJcTf
KACmburjCIZBduUG5FZDZkVqA+mpX5fHdWND+VGXmSRRFU4fy9K+IIm6Xsf+GBb1
zlIqRUQBwfp//AXZxR+s0LbEju2IyAstEHSocO1sHD8vKRidOgRjoFK26N3n5LrB
2s2MoZcxADIaruSJ+ipkB2NN2Mzzpl4CbuVBWgosl/+3cWJ7szVkuuHF12aGb5tP
HdLVgOeFaa70/lG6o5TJcLxFxvccCdsMcxavCoN19+V8dK2S81vQ/eyjDoRwa1LZ
Ivg5QAYAtnJFoPDnOn0TdbNjcjBvhnPuaYjE+Tkii5xM9ksclHA7Od3vOnsoc+jh
uSbwwkZR47EtLtxTfbDgamFsAmkt5v/BZmJvMZd0nHx6XNd2NiyOxBR8b6Guvm/X
yo+uJraGyqRfJF59XS8gqySJ6GIgtZMCUTSDypRMUu0D7O6MZqNe8OCDBLHIErWd
O+abdzOncCUzS+L4MOE/pOT3cw+UBYJ3a4MQ8LIoY+WHp+uTXMOWp2274cruncmm
bh7TzANNAaUj4jIP+JpW+JAG1Rhi+auZesDuvTM2dQnKsjDR9+k0PrYzx86cQK8M
l1X3pgtgLAeqcfd9ltFRmgzMnr9mJ3HhwfCRgeFyeeWCRbznt04+0p/20ts5y5lm
GjHVRXCARdOXKBOllhMLR7ZAOke8EPEHCfqKZ7wSWkX0C7SgncQ/SkFp2FgVc2U9
o/ceY8gS3QdMZW4/fkjPd3qiaXObOZLmmVBiHLmMT/pmeU7/CIgnPHFz3bXKOnGG
8/qhFydmn3GImKZN6q4XXbFzaMwq59fw8vTjBCYKEIG/HEX7aXbw6jYJ/WFoftuL
QnqYaUFC7+ggIMOHjZGSZQFUK4DcU6y0LZZY+1ZivjiB8pnpp3TB8cwFoW8bHJx3
O+iDmroRH8ct39llWKkckSJ8t/+eTsL7ojI+vUA9BxBnXwMZctocwu8bz4XPqpP6
ZkTjEm2zq1hKgauUsaAJ2o480HbGinc5ws5mKcnG5N4RL5aRgZmb0yqv8EuOyx82
/koueLPg0AHRAoWyxvbevUHE8y7QDNtouP3X7oC1c65qe6CcLCkgPYKS3VvR5w7H
4m/1ImLFgpMCw9oHuSs9tHEdA1aUE6aa+g93dr6L3lASVYzXDUKOXkAWg23iViCA
MyXvWGxCZ8kZXgfY/rU46wE41X3ZXfX2lizxwUF7+0KyVx/THgUo05iYOSHfcaV5
YNml8bXPSPc4lFcDST/YdS6SKEm5fOU9sLqGam7NjcouG8sj6unk0AyzL3S3WRDj
D1gSeuZu3ErscTPsDeHWgkvjYXxQE4vXXBuNp4ZgEM6h2DfFxyW+Nvp95S1h2mdH
HBAH0NTfnJC0PUPqiOuhkzd5j2peAMlkw4vD8hVdMHebKArYCSd1fmYXHxxaxNwi
cJwXQZhaBIeXTf+SMMQ1QtYtniXdOINH+lUIPHQ0UEaiI1wgTQJYYyPggziwOd5x
so7In3SvBeNazI3ep92CPByn2m8M3snpxAraMIN2jngY/n9gvYw8bNIzKiOZSito
DOIaxcTIzMcSiEfqDNHR491GwXGVyBEPFfZy0E7m1bt2fidgfUIdlZ2gwe1O3Ung
FFrA8PFA1bO7SAgdg/4caG+k16zJ2z1m9qdStMCf4aulyIiZKqicZnSQluz7i5GO
RRGQO0RiWepuETzt2v0JN3SFdt31f5ZZzhErKZj5StNYP2aeKEOI5Zvmfyy0IZoC
gjcFJkiInQYPAtcbh3WeFaRdV+pa5Uo9mKZNTPq89xt7+DAeLWi46FFnzUEychEL
bDRdnN6MxCRsbVriUPD70f938krWet8AncQM8RMWicK/Gd1JlQtAkC+yWY8nIs93
adWCzmFGEO44EMgJ3Qg2Gs+I8945K8MfgOSMO9oEp3f6+gVK9LaA2XQ+TgcRKAv0
9X3D6OjPAOWTC/qrbDHBLbIsDTCMzpa9j76SLD3/jnsZe0jO8PE6d8K4GGFRVMgC
pffcgy33kPNtu9pTiDgdpdAq0U9wKdxxmp/PW+mYmaxDABcjUqUOugkZJCir00J8
naaRTo8uyP5Z2bMMmAkLWC0HFo1PSZQ3uHaGhsO1eyUX/V7URHayKF7p6SX4J5a/
3SiueZyoJBEem5RrlDXfLcTAfGIx1vLOO+dE3nZ9yBlgO/LbQoRdn9zcw3d2T/KF
Vse9aqoGjstM/sPWn2smsWKg7yQ45voVD05NSgXMERrmwu+cIWBNJfw0AJSt8mlJ
mbIwkmHRVUnZpMsHdzR8R/OWcvin8rCJU/Q8rM7xyjjAnvXgcSs2dYSBuaaHDo4B
D37G2ihmgr/RSfUsknpuYjBNNluwg/tZxiQe/GXHTnAHE/l2BgGV51QIaO23BQps
T6FvaLwluPa3CoU54vkuYCXESFTE4kZF7z+42QeTgP4NdNULC4JOy3RxvqKbb2Qg
uXyEOLweLKtfh1yn+Qgg/WxJ4gywB25/lCelOYRTL186sPITINxBtWXmtTcXeJE2
WhzH9gGv9qzB7uwlhlRI8lLvuBesHTDxOYgPzr0c4TKoZlOCZmA1Kfb/TVGfwPTB
okSKI9Vxptl7RNcVgcK+G21rFS4zVLygIFk8COhVNano9IB9FTXOFKMKppXiKbp4
aQwWeb/3YD6tchjac+UbHu7ZnDVLKn2yWH+O6hPFhFv8/d0Lc/TqSUsgV5rDP+Fc
z5gJgY7x/XnDWRcO7BeWP94p/LrdFzUaVF4D0vEIlyKSrXfI2r07uJxrSH8/AA5d
u9DG86QBQBQLkpd5oKWthtqicqfa0/zQNuRr1LD27mXxt4RDvjHsn+h5DpPewOxh
qck1HwASHC/FCEANfD1+zVudBF9987G0VvpifAh0WoUC/JGN7FGeofVFwZY6DvWn
ap6RL98NicFgnsi6z3Bax8uM4soy3oazz7rf3NBnCpEbCafCIPi05+aZuxTu9s74
8TEfNl/sdx3f6irbAwdGvwF7+UPGzAASsYONkvzZ7E2EuWykLcmrYHRI7qeghf8s
4mrnPH5VBrkdS14O66iDVtNNZwQ7FrdEUr2S2+QfOEB4sJ0AdaGpjbxVmAlcL/po
dMv7+KKlSLBHpTH+CPrvDpQfvyosJwV8sIGsbpeN9rztlSGsnh4xRzNVxuHnbdu4
mpJKLbeWKDbogDQSzC+DCyNh/k25urYGj3HI6IGQfxWp7SMiG/TIgCy3AHqi7YTe
CFYFxDZscM9ACAZuGjzhgq4PJpmfjDrrcB1UB5ujlgfj8Lc8wSEop0MgZvlTarXi
QgjHzNqXKERvpdTPxfg6g5qmOxDe7DAcY4uajJCBIBHOotwGNe5H0e57+rQtZlTJ
iRadEZRde3mur/OGNjVe40ACpn6l7NdJbQXoi/xIRJirb380/W+aK8+XVNBCasEw
3Sxla2OY+yv9qomCWbc0Q7WyLDsfgZw64RvElJllNcFV98z1djrZdlEz9bmKN/DD
N3WtRZKRsKepYEuxHOWcTThcFRcGREiXLI8gxpRpmnMYfD1gR0CIHBuEBArrZmJm
VV5bCklsbDRgBpHDbZDb6ICJU4bnJchLQOmvVF8N6MyN1auALaieMUJfR7yFQYK/
7Z/mlw3eExZlj2pjwMt7sFZwZN8sX1kARGxNSyn2KSJWm2uaSf5lo0PMXl2l9Xbf
0jfFMwzp07fLOrPkpDKJ9tFH9CGrpRAZn+jamQ9D2IpMZnWZVFxTcKrogx09coQr
poURpvhljR5i2IeDgYQZnp8fIEcRE5xL6kbeFUBWxc5MvUEfeYumszKA0q5+9yXI
iaNR7Lvq0UrE8+dKB2EKSKQNrXZautEcdTeOjxoja7xfmtFUD1uPksluRGXaxQU2
R9WjubSx/X5Fzvu1rCx4aTZYOaQ0+fCAr5Trcg6/lwmSd2WtCJYhgdeOhXhwTQ2E
Ur+aE0eDweE+Avzc5/iuL2uLeA8zXD0l+oSVx109DJGgYiU7U0A3tlKTlBRRwBvx
8G7ZDdL4Ouivb+dI9NQkIMMNLLa5GgXzxgQmgy+DFg32cdlT/3WNqarjEMGXPF3t
MQUxGNBEhHJcrNh1uFH52pyvaGjJqnJTI8FOC5IM4FA+uG/GwhlKrMLnn6G0FfYT
zzgrpMh2T8dFVdeCkrsdlzhyGMM6iRKzYhfIx14cIe2ZeCn7mF0cAM6Q1ZEShuda
Mw2/kzvpGw0FNIwO8MBrsCsWYIPYdjIglspAt0pAdt76QmBhx2ROa2l6UQm1rG8B
bQ/+IOIMC5oRofDfm04wfETNyCoVqK066Wvhm7ewjclMrckMAqXC7tks/isH8X/r
WsNMk7aOiYa4eKdc/9QKIiV+RGOoJJJlArbwFJ35KGIrNigAu7E49uDcUbQPE2P5
sFKwEf8FmsFufSDFkTHeIDq/AmEOV686o9ZovvfeutwiIrWA9eyBg5iJLs+ZPV8+
zElh9FC1Q0b/v0IpOnIrMNYNakLXn5z1gbSaN1GFSvjwK7M1FDYkdx9GyFldyBGS
El4KbmhI98uBCcMzxJVmRZNxTDUE4Ie4pU09LctZsYrcIQKZBP8XWoeCiZFJ8Z3r
mIsFVklBLDC/hS4rDTjIB69gr/P3pn7ZER/cxt+M3IYoNd4ZdvSiI5MvuG9t/Qdx
7TTsV5D1J+R7OeyMbrQ/Uvwrc0U8E9vtuaqI+oC2Ky3vX2p6niMagiwyNxonLE9i
1105ImWTgJwrbs+v4k+s1yr2R8dvX9rms/wIfri34MYdr8e0FQGfypT249e3rIEL
xZKodck0rtodWbf4+QfSjIbdVm8bgchr4ivIBR8ZQpQ6EfvHm9jhOsKDmrG9j9+3
m7d/PFtiB/QnmcSyIU/WEMacpI9MIlxFV8fcEG9O9/Z7GKqpjO9a9Zh7zhbCWDYj
lKz58CzfxCbm19Kl0xykvF8Hd29C5DC7nCBFRpeuRf0bi7mH2EUuCaCmfLwWsj9r
rtpN05jJcGdpz2niXEaNmkeL/pjP10DjGQjx8efGVbfjFB7vbJ6E366M4f11vzGM
1PGYgpuylyzEYExgAckF3LGHdK67jC2gNrLKe3pag0gggbQIKGmBMvQy1NvkyIop
0ePjWRDWoBAGu73X8Z3H6SKv86jiiac6WgCR5WNqpwG8k+2p7H8VH2qt9yBlhV7k
LxgnUpjOLhr54FKiVoL2OWO8IfR4SAMJnvLHt3r9l+m9KCmUlRETb43ninNBm+QO
fE2Pxh0+9kuinkktrNuOXIeWv3rUyENmrz4wSrHPN9+cvXSa5GqOkq61SswGC/E+
ADxePFb/NonpQj/DD4FhOjFgaoxrfEyv/Y7VBfNz16fB9mTDZlVyL9Xj6/R0whCP
nhNtpjSCKozdJObgxZtpDyks+l6T8df96ts8aoJ4O0ZnUl1raHfqjEsJtFIu0oB3
q0rn/dbR1mTV1ICMUTTVFJpo3r0dc2gE5yEGljPtYc2OGbpMi0Ycq2MqpmPyNWIj
rquJUseOnkRQpxqnzeELUbqIoJQNvv8ijTi73YvRNHcCPXT5OywppaUidDJrW0GC
QMwstPFrOxt4jbOlhTq3I5907nuBlnSO28K9n+zrRogWpymlmlROXpjLpCx/4+ZG
RBftCjGRjuJXpHzzu64mk6pKY2aD09yL6BBadVZfjyG39zRPEQqgJc8xquA6TWfL
f9Uu+Ruu5pEETqaO15PzFUtZ5wKDfbajImKwbPjfVylsiQ14RtqYowF3/FcN4deV
Wd0jbkzY/uMordTf7CKvghF1UbEMfV6AZKu3+JMvzBlhAxrQ4deNnCsUJ658/VAy
F6M8D2OXQ+xTl1Wwg96Gx3ja58j9KFeFFtSUItk4EFHmfDRHQFmmEEtJ8qJEcfQo
zJ0KkCZ9cusauj6U1wGc5wBk9ZUHBWCR1u11X7GoBF7Tuj4YwjKLufsNrlW+ybgd
zodDMYb/oLNW+dNBV016D3FT1rdlEjrGHbvtbPXR9n9pHmPMFTY9b51pyJoNLvmE
4YSnWhfkhNGJlYfTc0zuly1JPvA+e7Egne37aHeotsV0YJm3t3/uBO4dYXl0wq6t
QkIMjctl3zxjBtCWgjEu71rBMnIrP8SdRSnfSzV+Un4IOcQn9h5tkqSCbFdJR42q
k4Ds9MCw/Wa+pem+8kUXeyM8l9FrHYok1NbiHNAYWaPfS8Z6Reet4zZO1P9GeNZH
NVMwriBnwnmsgwhQiguFCCs8boGnTewXVDkV4aympQ4FBmgEOvYw24aK2XJ7datg
CqF8jjPI7wdqRLAf3KxdmUgFrG07WiQ4cv+I6nUN+DHV1X+icqQCenDhkxLF4OvI
2PRHnt1Vy8Av5GWtTvZs/B+qcKspUr838ba8geUZFL5TTqlwQuuDzVLdDKnC+lyU
rZPoe+mSdp1bScV35riHOqGOvMwXgjmaJ3G5FcWhwNDjPuieI03k5ftkno6o+vyL
CHMtjF1eE4ZYAh84rVsDebKnUZYBytREtZXRtQDQBX55ij0KM1xqmg5zogfDXWzf
JNFtoqyg/upy1Q+gvHp1i9faRnWc7++0/8zhhwyqPdTmQXyt63xY3cgmjMKei4Zo
4GwcSdRYFOHqZ6Ht6WkYBVrvrAqTf67OkoV2iu0vFUt57IzIwZ2XjyvTum6D32Sr
islOue+BGkngubtvXSH3DP8aLrep84SC1W6PBkJcjbl6yPZqWXmWzdRBtHVFfgre
SMihMmpLPgfL2bzzITAil2PoDF5WNhqSJCJAPUPme6nZ5su7tXG7e+BR9uXZ7YFF
1+va49Wq+uiswsf+aOzh19E+rUBS3LqOu7ZC2hEOUYybDuVblez+yhS4skUlA5BS
Ijw7FiSc9eGtkzR7wXeZ4TdcEyqnx1X/wWSYccTajk0RRjH1k6rje9LUKBycj3RK
BuYWuwoDCdKkWnC8uRCVkClO1GzHVtOpYQCmK3KQkSwFKMcY6v5ztWUSIZ860vR7
iwDYU8M3/RzBlYlB0SM3H0+di6j7ubJg5T6/dbrUURE9IPXHaku5HOlExoWnrT0c
7rBrJ9BtYU0Awry+m41HqKKurbqmZWmkoOwAelw2vza8GEZuxLlcZXWLEQlYhXvl
8bBFo3BwZcgULDJ/ToZ4uwWE7f3sqODs6pqwKiQZDGCty3+5Qvan4opl8xHXQkKe
dZwOqRb9w2JAgoPS1tcFP05iI5WDG/CELMCssle/3BFWeDawVwvA0LpRJrsxGeMS
yf7bCKVNhzD/jiFFyZQUxQ9PrsxRVHDfKR/Upx9X/lheJ61dxEu1xcZTeBkhJQ7j
mvmdiH6+N2CwN5ylaP2XeXfVqETTmpo7FSckwp44aoyHynsBHtQWwEi4X0zqcVr6
DkOPDlln6JhPOaiMafIMZ43QRueq3CW/ZXU+FR4SR8tdnsJP0JiJf+Ut7jQKzEr+
7Wf47RIAFh/pmukf9VoB0qI6/gQqIJKZg2BTcwVLao4I/ReThLdluQSV4UEueuCg
bJ0bwC8W6mjxyk05/nvFvdO4XydoqMDt+U6SARA1FF6kPXnzm+OnsZSmfrA2CpDy
fw1PHkejLHa3bIKg+1GJeeWAxJDdQCmsfaFdjj7NzMOjakMP3erWKlwqwQAriPnc
MGzsTLg1Gvej39Y0TUdUxtlpBkmJu4ZRV4zYyfeRKU8xhQwB3dmHbyQS9M57Lw+n
yVw+D1tcr6XQmbZU7NEfEzsp9+WwCA18gzmGHpk2KVfo9hxJLxsZCL9NVJfC64/I
DIJ8aKUINaEGxcvs+9IQoEyGFUe3cyNTfanatWhGD0jz07EkRlYKwGEha2vg4bGe
GR4tac+kWUrdmM9wcNNfKfj9iUvvzhuyydnJeBmP9T6g7MYHgAuFixPGH/lKZao6
pOQRLaz3sRJjGjauSAWJFNzb5rD2+1gR6mdfhRhUqDZvY2ZanCewFIzTdHQwwBLa
/lA0POG1t6wCxx0qrRT2RtsKOi7cU08GLfzxiJQu7OIQcxAfKRVPqkRwNxgftF7Y
5knU30PdPEfkA8o++oQptgGjmGvrLcurwXMbtVg1s712JJGgQr1L8Dj5t3RlflGv
244qtQCr4vImDKJ8Nh8iuXyvJh3tF0b3s5/Hun1/bUaPrL4uoxZeJBsxMuXiPKVl
CyH2XuKDxHpE/02r89T0xokeqVLkrhhTS5kAk76WhBnN9vjsEm8FQGSmx3qmRjkU
JhYoVkw43dilJZBOUz99UPnNkPxQGZaR8rZ4P+AeQWDX0FkoTeie3kMzvcaTDVkW
oxQJ+33E8+2W9BocZAeV+T5yJKVuHUaUvgZ4Nx0VXhn86kZwg0hSFh4HyVVPT7f4
wybaHTsoC7xicfiCXrpLbEpKOsWkjitGbr82pI9tgOtPao8n1Z623dTvNsUwuR4R
XA89LcONxxS9GbmSKhdCE5cevTsfS64FPC8Md2t2l7H0BtEojg5PzUAwpa+F1OzZ
fec07hMvKTQ3lOCLqKq1t5om5AJLY7lPhqwQLytzTBjV4JcrxKZ82prtiVVpbznP
YD7rF8BvVW3VZw3QNnyFD19Q08OUBtm4fXFOEhGZylqXvb4LLVHze/5gEYHQldvX
l0TBPKiYa8/QP80e2kL3KsN6ZV/IkgcwFop3lufQrxpkvwl6RdurJqhX+cERPpWK
Y/X7y9G8MeKK1eZreOPxIEzvDMBEMa9Ep7yTfNfB5AobN1+kJ6/4auMAsmNRITqh
Q8GDu6v3P8E0rXRVUhX7g/yA9oWosRADX2G+DMOj0bTkHIgixxz/Gn4dqkreG0l+
6gmx6wMgIJdU3791RoEYNKgZ91RkkizCYvyMQoJfOjBIq49xIqRnOj1FDAdMCeyr
s2iD8bu1xHpG/MS+EgJu5miULXpV+35bVKBh6gL0hbxRKh+kJoDKjyb2Zt7AWEUm
03zU9VAiNA7eBIFPnu5qpG/00vD4iyzUhSoSaZfUhZVQNS7LBxS436n7jS098jyq
QapgQw+JxnPnhY24CZr0GkTiBuu4Cg6I9cJUUlcNJrgizI9P7U4dWlbzpxCFZ7IE
tGiOTqHbhXeEtP44dJOMQ2NP2Xs/8I63w5MAXz1btbkHjvxfhOZcnyPNQdc1g3UU
kQVq7s0bjIrleWp414OB2mO3s0osjcWx9Ba8iGNL7LJ7EAbzoxFmv6cFlYyCLPD2
lWOTUuI7vUVRZ5FrQCfV1Hr5goBqIh27IU0CaPm2K4lTejcFOywYwH89J4P9y8tM
H58izfzRraxTGDZ89vTKiIsIHPwLY9ZvNa7t4GE0MLicUCa2PHFioJQ9p+WzCWtW
W7n4l7ikyG4/L9xy+BgZXQbxcvvgONchrjcFnn3YzS0VDk6IerUhjodaESsAyQ9F
tdbER4LxUAYZFTt/z4GASMyLkjCadAgTHnDpljcJaMnaPGVpzkZG9ZaThglt1XSF
7ZfnmELRXT3fs/O6yvQSRxCczs9CEOsbLL2U3APJw0XQlbNRVcyFvkxRheAXOX3s
lDjy7zpENuD7z22pIPOYccJQtnD6IYye+boaSQelADcT3rbLY8S/OGgRot6DzSA9
FEdoL+8zsv2L+AXGPtwL6Kzd5zIpyf92hQQgbELy4K0Jfyfwzv8k0b5cO8JMKcFO
SZEMKX/xt4F74jmlk5agf7ESH/ZfXzuvQGgpJjxCA9aICSx26shrXvxQUsO666lM
x/+RRqKUhxyrMeJ4UXHYIc3TT62mTMl1sW8EtJHECX/w7VyG8PX1IoPP1mDX8Ul/
PpYeg2qxui/DWWFvgUwlSKZQtJh3ckJt74ELPmBg1Tr8Zi6RBi5k1+Q2ssGBrEkd
kroowoBv6SPQ0OTYZX7u9k7wOzayl6FJkNoihXucYtAZ4ou3693AKVrF/UsDdOZK
D4A75Gf5qHGJKI15j5HB+vmiGx9fJ4FCCzFfS187ew7x/lEcdn2UdIyOAPKymcLG
LhOzioRU+ChI+0jvcQeyQDF+Q2+e3+U8tKlJlfXYjMLi/Cu4hLpmHyMNuZReY5N7
LYAzYoENnOkjyiE31oBarKlOyNxnMlHL0Ht3vfKrXQu6prcinMOWD5WT2dqFEZ95
oqONDmH6tbjzuiVdx9MQokWaOSkyGZVeatihq1WpZTTyTkVEY4A2d2KwAySgl07u
UMvjyC5cV9yV4pLvhdVYzugBYe3gfg8Uh4iyJMSu34aSrdoUdOCXG/rukhop5Bbs
AfnFg96KAoOSFzVIGx3CAHCRmcI568MYhof+6cDT7VQWhddyeZHV+ulEEmdBvG3z
aIK8Id2PeEf3ise29EtVpg/un5s/Hva6TZateCyiJJVjU7uMvJq4eoewLYPaPWbL
lUXxiuU3kyelkrNiWMq79SbyJFgZynAfhFV5FlZyvpV2SspIZbGr0E0KH/IUI5CI
sqjfw1toyjwwN3OY3ZmuYfPGB1s5tc4ofLNpjT02EwvpmZ2nI5PLjwsyje5hsXvA
Rb+b0dROeWDpuRYLFs4CAerbD8vfCJDjG29XqtiR0D7K5j4im3+eFD+l2GJzEwjK
BjKkKFZA1i+Su6wBnT2QksTdoz1sYAoXyRMoiPKDYTzE4UIJ26Ttock1xEHjWPkk
2vIaBJlemMC2FpHgmDbPxOVkciZUpmOFMCX9ckMuAKCkMWbZiXsX8bqMJ/qaBJLB
yhmWH6R0RquxUdJ2Jy9XhE4maSeSe1Z45wRX+wsCvgRGrGoxI14Iedfs8Kqg1PzV
ABqL4nEUb5E6aCZIQH5GgnrqRoiRhmKMpw9+32Qa1W5S6oLUKUsaIki5+khsvx4I
OGhimOk6lfYhvZJ0O4JESUkPIsiK2zi3/8fwcjLyRSW0+zgscXOX7nikQfZHrX9Z
d7kKJ9moXubnrjiHOnMA3EzTd6AJ3K7KHap7FuaCHXm8Eg7suCqA44tE+qV2q8XO
FIayEi71/IOZhYvF1oLrhxXNuCWlP4ucaF82U58eWGWrgXKFPCeaf6c9J/LCxWxQ
i4D8rIZFmTZi8JaxysE6vw3NYmR4MomAT3oMjRBo/qTEy3a0iey1XVWcVGWo97Ck
XH5PKKCDyWuLxLPLdjKXVfOKAVTj6/L8vuKZOJpTQ2AftcT+gTwboaGnv1TqxyWQ
aEwlGqjdLKKRdrDP3Vv1jBoHpiGTGEXjJM29w+vC248ks8w67jys2jPtnQE3Bhs7
c94oIhO7Ui0WPNGHjk0g+N/cK/IghqafMpjEBQZN3u66B7LSofWVRzkV2QVYpprz
LhkUyXYKpnRyLf48CZV+Gqzega5ZOKMxJYe2Qy2tJQM8iNcVv3x5gPtn/nZxYdsM
8m4ljHaw7t61SUCK4ApN1FBFvFtTMhpe1vgpzkNUpRj9UGLjBEboee/YR3ePL6qK
HPMtuNONSmgrQFMH0o6n/SWp6YoPgykCBAUdtUyfaFN4GeU4oRa6qNJmZUa1ZXgJ
+m2jujOZQ4L+v5v1DgXB7CRA739xZUaiMDmCe4jLUU0P5xWfUwrzGuzFfVF9Y72f
1VE0XdkzF9ZzDFu5g7oBHaYkE/rxxJLmEGHRy/8VvXLpcuM2QYlbwPBJOXgz2UhT
Km6WpwAmXeg2IEoByPnWzCPkztRiVUU0q4kGnW+fehNUt/47ewbOMYjso9AW+2nq
a3kZ/sT5lxHOpY48L/2sunti9ZUb1WV5R24DyGpAYCdTKB+J4Wug7T/EuRHEVste
AAO1e+KMlJqsGvOhNLGvtZW3IUnP5LHjXuJ2MEBb83Iqc/gE+ywVR9A9ZpfLUdXS
D64WQz8LKJZ009Hxj7z0q39lcWxSWHRSHwkCFvf2ZWWmayULzaoRln6IltHBNNBv
uUyfFbuNc+pc/etz+m7CE3wVU5bEdxYhNh3xDE64ZWmJeN3ji7QV1qiik8f28tBt
ngfzWJqkylLb25p2JSClwv1MjwRf0ZzU0hozj4x8rxcFsxAPz/4OrTZ3YRo3Oi/k
kFVUM8xNXZqUDiPBiw5W+JgLVfeDwsMKOv5mMUor69W+Bqc/TyeWOUdEjwDghcPz
BqN4mw0CtSEFth//m87W58EbR8Gl8eJc/IzjVfUcteWRmSjzzoCCWyQ1jXkW9irP
9VpzG7ZkE0IPtjnTtNGNSgdfaew4wB1ocbSCS79zgOaTlLdce/xnH0VsmTHMScUu
xLUpl2N6p4m+fzoa4M3Woqg1/9TrR0GdVOLhmFV7O89AVQaIH8omrwh+SkTbYHll
xg3aIISwhddtkW/OAvj6ETRqi4f3UwA6UOFfYsG/tyPfMsPTZ+CXhuDACX1eQC1d
szJLYmHjcNRAgLrpP0f5Eyl7u23gJ5MMdLlpKEEiGH3swvTUHpDL+7h68myfl/zv
LyAms1K8R0Rpc20K3Ck3GpWWWMG3d2CRKsCa7Uhk9eQs0qFjZ5EMFjzk8qZl0LLR
oqCvT3GZc95uOuxP3dTJqZtD0nj3TgApyhG5Q+mMGxOwHiU6Z1wWI/qV+1iK9hrc
E9XF+We19QaFcZsVenxfKZCWAiqfRYQCXDwBzh6D2QmEJIIvNqS0I1PoP1m8dxrw
KLQmMxqdlnrLr6ayS/lZyKcypwb3IVc7T0/o8qvxUmWxFw82BQanShQRS9/hwnMU
PaLqPpXdjEvzDw/xa5Ka/IYCRWSw5YmgfBMxKSozTXI1KYrffJPqope2SsrL40MO
Ic1z7EN0S+oflQ3VPbTb8iT9hLMDKDRbzoIwLjuow28AbB5TUiOZesYEN5EDP2Hy
v6L5h2srhYM69VE/c8LWl/UpcVN5dRu94j+VTbspfx0uzDFVm+RQUQeaPfJAOiZU
1KKFOVHxdPNNmorFJHO3DT8HDKvdJCNqWeQ2CPxh5VyUrp96AdWU/yDa+pr+cVRh
hAlzt+Jszgp5TPi29F08eZFcZAqwULIr1+poLEj4ujzfktnh/i8CYNovzkpaRGZ1
7s+fmxhjK7redh1ugzyVZT4WV9x+LbewXKmw126inUcHKQH+R1qegNn8AFsf5bRU
vxKO0w3Ajg0iMCdm4iYpab19LukLb1h4oT3x6Eok+u6+su2+VGOnuNUEDQlPDgW1
gLqQ2/ahfWFUU0Po0pY2DPueJt8w2rdZwTDxSSgCWxmoflWgs/TBkUsl2VgeSRSV
9x0dgGgTRWOMMUKTWbev88q1q9CLSj9NG2IR5GsZeTkq+cDufcupw+kf8n2S+5FP
sqNGrkyPf6PBFfVp+cZfIIj88xZQm7pUHpyJzL8bhybLFjvh+8tFhfrTX5B0qoJ2
6HQ8W/L3V4rA84+AI5OtIfwh/qmiML8cl8D0uiDdYlnbYzZNjdVNNByBdF2JDMWI
Hp+oGd57JzmhXXLTvqMEHQQDlHT/izDs5vd3YgeJRkZhdHXkLgWb68qBJkJ9O2QN
Wa9LuvyQTLFhSOwvAuOe++o/mW/UXXmO8RDtMPdN7IEAAOnDAbpknZxPeb6Axy/j
EkSB+3K/q19Dcdm3IoGXFfTYa6xv3hvpucTlqeOyEl5cqzxGEf1YsAY4D2OCw+V1
VeeOV/zSgC7q6esCQpsvXIWwmkGyFOB0rzAtZQMezn6nLTZL0z1hsJixtNHkv7x1
dDkF79/2w41uH2CbpQggmVkDhxzZQQF0NcDaUfcC/SFm0HDj/x8o2JUM100r8niI
t21KKaG9uxOpjOCBgrIuYXE33DkgfG+D5n+77HeDBGCaFLmGJy4OWLyApCu9EAu/
AuXdGKmO9FUddXZhgklOwMQ978jeOibp/7dMGtyAvj+mPGdQYYE2qF6fxXlHEedk
HwvNjPKILqIkTQhmuN1jc+zONAdKIjk8gDaOJCCnKXOhj17JUo2PtShqQTi9M0AG
b3RrqWtLDM72+SfEc4c2smBU5bHmOsXb8cuAu0PTxOg0Fv1gcIu6O4g68YR8TXeT
f6dZP1iZMlb6Q/K2zzQFxoOzPu8x7n9dBzIG6WXms09URx2Zg3WIpdycu0nwbZXx
V43ul7u6bcH7n/xey6PwGVNIk4CewuaFVSvZE7WaQ9o9nvhuzriJNkqUKFgdEgv8
1/mltg4JuSUAMyr0BQ8lSJzE3B2hJpLFf4TuwjukuEjtmDkRwc92jLQe/bVadBZC
ZV/alEsR+HrAgo/TbANirLXUx7fXaBds5dOH5sRgQ4AjVQbu8ckJCARNXvlWZu1m
V1hrCph/YHdlVmSvqr/pqiEoN3sC6nlnmtKIwN50lnytChkhSv2GdegQE1WctJA/
74/X01+h79iWvP9DEUt90LeiIk7cdX3eWazjn0Vm5Cww9eEkmok9zOW82HOrnR2O
FFqvNtrscqywf+rhliOKH8iXry1KIErBE8mbg8nbjghgEnPghNha+8UA+htek0Rl
EF11yXrTyh5TUr02K3+yVclFTFboGVJj5rFaMYsbPX7UuMX59kJxnFjZnXLpbG9h
mAkCzn5Gd2/ZfMfE9in2fZG5OBQXVAVMgf0aSof9GGlQOwDxc4lOSGRN4VUG4cPT
pIxG9+Y4/4ZEWarcpg848B3WVPXRHdgZLLH/68qtv9XlqQ0x9GaIod4KR0l42AG0
M0ZM41wVa8m0CRBOKu+BFwPhyOBIVpP6WGKYIGzoDmFPhRVsWV/ssdQKjP/UsQPg
kPHb/XOnAeO9QEO2QohomKd8/k3J05vZMtQH6XZTUv69R3FhiXgn/TKafd81/q38
9sHtF4Hsbormsu1Iij1paVOnHRGj7dvSrV17qkbKXiS/8hJ1mWcLJIsSru3qZ6T2
H6GfqGFUS/0uQEOAw5YS1CZbjrau2rk7l3bNyKa31Cf+es1z+eouP4USGqxb6Enr
ifjz5NpfXdkcKycbMUDtW4UaEt8efW8GHBxj3ZZc7QPesCcSiwACPJuSJyRKKDRW
zdwz72ek20DeoaTFqlhlGIz5y2umzB7/JyyisSGBKosiSxpZVj7T163RXeDfUA+Q
JtN0XPUhLC+ZJlMxw6caYv5jpn6bTOpbFupcmezXeCSUuNzKtQUVJeGA0WbslTI8
4dlCwBz2Ah1KvWkVGhtuqkNMSkpl66WSZZgq0qxxQVeFCyYHfAFlyEcg6a0myQbQ
wydXqOAcax3aqWx3hNDF3I3LbCrbfL30jIFSbamD/vX/ckKk45c8HAxId9WQFa3Q
aO/lpE2a+59mGnuGEoA9n3eN05yeNkVlVuFtejVxf0t3pnVB0+pSdiV6TC37JOcj
s10lbjKKd/RfV04HRhuX7zKhm/je8jmSbwX5yaC2hk0d5PFr6jnQ92kjqGd16xjc
keEnnMJpm7ooKEsNWHKs06kv9uEouwT8PA7njetg2Umr+t2yh2V4ijd8xbJy60YU
GD5NybiJvHhxE0Mgmb5E0zcOsCDVAl21srU4Pv1O4Oy8P1FDuOGmDiV+pPWvjnev
2JTwLmAfbHXG4nUV/hn0xFa7qaIz8Zz6HGDjcieNkvrlb8zxKlSxPvLCwVxaCaUS
85hNfjGPRdaJHlPrHp4awFBFpMbx9GuFSosokW6sWElLjVGTBrb/+n3xmRM0dEaf
YxYohfy/qAwy82OJJuMzJyIAyudaowNpVIcMHz2keizgbkAJREH202qiRn613IVI
6C44swxapZdgENFK7XVd65+YcTkBdBkGTmICNEnY0XjUYP64ndJ042Bt5QqwdaEu
v7aYg792Ua17RO5jujWHqFtnRhF6GqiQC0nhJeitUpOEITCI1zjyBvyD7uMvy13w
G3/GrrMfeGpZlOSiDCY48kKLFcBQ5dOENJ5+5XTFSkioRaRwjLCm+AAZmXW7NMsQ
ttlqBz2gC8hUJ0K9FRZxcLq50y0eJLS18GsJN5xEZ8RB8iI3OScG0yxB6x5i5mxW
Gw7MJ0jkH8/cYmktjsAGx101uMTYNKfLs/QBjvACZE66vsA/SkO//APzYs58B5eC
6G2LKRpFyiRMEtdUPcUyxdudf8fbsueYz+H4/r00EfelnOvQgx4Azb6ntyfJkEqc
MRj414jROF/cAGuatx5a2cVmZ+mw6BZDkTcb38clqz9iFsocHLAx7aOCx3eYd+Fa
3O53FCOHXkBTZRiAro1qxGdIwNAak3RQbCAQNU1gmCFVrx/YTysBr8HwAxJ4Zq1Y
VRVVJJaLY/CAvohaivRsI+sfO1c0BVsGmdjY+nC4PO483NpnD9UTx5Id+8TSgUAb
cPlHMUOBm862P8EX+MxGIXHEFFBZ9UvEXqe/lQy9NkggQfy7w7jVwGhIiDNlmYCe
ta1ZfGkrLrE0KXqWzSv+ieVM/QJ4NM7FmYoWV2qMsz9FwGWjMgbL+PbOhgN5LxLR
xthOAyWKvZeem/K+6LH2PhGqPfZujilCIlK4XD+AeDLVF3oxc/nDgDzksQIMG4Xa
cy7O9Joxla5MxKubYWJxItbsS+7eTP0JAKar+PNacCH/gNQKiUaKFyj6AtOu1Q5S
Tk4hyOIm3bI6G/dezEY/1680CycR3vQaqpza3I8QufXjnkokT0tG3Sp/lxA7UPfX
nekG1n1d1QjOP2r0SoSVS0VHXUvyym6TTkUpUdvJIsYL0JLXhu0JRD1F/SPpHC35
+FCMjjkLbKUP8AXcs/MIUaVpby+uxeEQWWfxe/xKy+Do2V+6KjyEg3UV+QrHjCSq
VJoKkEcMrISkKa3H4tBQEYHkp8v2pW77BtIsqWEnMVyCY2doCBuq/iHfWbvOC9ra
D/6A0ylE8n1SfG2RSaNNiDXWpvWeip2mliqyI99xvzT2J8iPebQGDroarqu/iJqK
Sgy2am0sBFrUbv9juyK2PK3Z3Yb2GhYidgb7/aXaYYcSUsA8ChbyxNz4AHSJM5wx
kCf3YAObwJUvBBtg2Xja4SfP4Y7iQJD82v0MySsWqpXOuKfbaWKJ/Tas/tn4Jh3I
OgYz9Ha7U0YOMtEn3uhDWV1PROQ8uxJmCP4WVwEqcZihdXpvxGLgxhdjDEdah6uV
IprYW8V65ldyHpo6phVZJPhD4qGH4DpG/8HNJwl1Dqcg8kOqYq65y3ijFVfNXZQC
OITXn4CnP/l/S0a8IOl6ti8Qcsfn5rXHk2/A3QqIPxnTCYzU7Ux54DxIbPjOJPwJ
cHSdFHCDAaDDut9MNAKgBporXNQW6E2DVSeo0XbxRNElzdM27lLMgjjfVhLJz/ZE
0YFUO7c5x57AnuwxbZj2R2xzoH4ttxc8rKVxyt06efwzLNBiFu3H1WksNRy59CrB
WFEw5yo4d/tSwicp/hSzWQjm7qEYtmFvyX6oMYiUS5EX6gHH52w21fczpJH/IvJq
bVPI6KfE77mOOw46/IBmp/e9fpHrpenZnAuU6F9ez6pPNWwiOm4TWe7IXj++BuHP
9mtbplfd0aJpMX872DQYESa4TfX70+j+wMHQEAmEgoIXEv+pO1MFkRS2JgBaN7Jt
kemaLcs1FHYJoCcNVuOkrPmmoI0r1bhcXJDhGRL6ayE9PDZShCfoIi9dioeKJPlr
YpJBSg751RlsR1eARWuuv2NnojWmQHmQ5N6IFTxXlZqgJlcbxY5Nib3C1QNrK6Dd
bLdSToBlwhNf/hYuKQJV+E2hKLpprXM0cSl4dUk+kac+bg/PwgXKhNVR8Ts+vnbj
npBi9H/zqHjenEqRgVqdZXVikMqyGbd4rfxlqd/mykVhte7RMvPmbaUstFajnymx
SFE1lWvtzv8brMThqKOx6EzFLyu+GRTvdUxpeMjhdxk1iqVXNrAV+jBuGsblqvxf
fYbnVmY/pHLjEKf8y4511+oZUgP+rDfRWgczeaUsmcYYztYATNrniMrp31B6qLiJ
pN1P7rYPVcVX+JsG4mNsrPzS91f0KWw0syVMu4Ns5alxacBWKnABkoQs0FckoIRQ
032f4d9+pC+frChCRpTpTh7a3tJwqXqA3nw4Qlgmq9ApQPjXFEo08URnEDr422Oe
lqyZdhTXl7Nx81wG1y3Qq3UrKZW81pAV6fEWzrrfMmMjLQ/5l5M3REilQUNHGlCe
6OfEvpLAt0YY3Kg0qKF1cw3bstaVC1WRKLK5vxdA7bmYRQNBYHAUabMCjoYjmuHu
ZicRIFUp34y0xUAvtO1sBb6EEMzaN8Oin9Gp5BuF5RuDBLeun70AUfH6fiPKlK2C
mU6RDeJm2NmkDcCFCsDY5aAr20frSTG4+8NJPidVcaQRmt7SYsIk0aIKn55bDUyp
4QRLE8F0QaUJzzc2B0/9kckr/8t0K1X/kUuTR2rPTWgM03VJMX2xTQgExv8Ajbch
Z2RtvFw1akrs12IiQCrDWyzPr7I6jjUGFfDFVrGSApFudd5sLMnWzs1K3fowVUh0
+ue8Uofdkk8yF6VGCoDd25srmmQac/pE722BNPvpNiBxkKcfw76XsRDEqbuV2j9A
4o4RnWnz75uJzsTuiVp7k/8RoJA6rOOCC1UnRmJDw2RJuKWpqTx5s93nkEsZHFtk
KFUYA1YQh7NZYkXT+ZhalNxyoXzVDxYVBYX3hHx/7+xbZg5usiFpC/nYvG8EofZm
Az94rB9QDJpuZ8l5Zvx7AWck3WHH5K0yAU3YS8nGv8wdY4dJxAGj4JJu8RgyZLAP
FKMkMFX4CXYZLV5Mh5nT2evlSmHVDmKKsIWZiKV8TsDf+onXfO8gofLnnno03RSy
OdUxCl1HlJYXWVooETGJ0uNPKfFKCB8Br4ch9mZCDNT6ALDt1GU+Y0muJs1sEzQK
4gWuGTR9GDo1rMZYJmdj0o6qs8MgdRj4Ia7nN4rYQLEHc92VE0nnoT7/tBUk4jcw
ZZwZDYIwWO+zKvp3Ic2vSrk9lPhjGSKid48717fZtzBYZbiLVaLZvhUeB/gjNhDq
CbDh7OKP3I3qZ6FhfzB3c96tnT01oRx2W6cTJA+2PsECKugfaB/DoqRXpuvBKoO/
gWIojwm5EDRPxW12PoK/KeK6zSprlzzQdz68OM0pIUP3QfIhBDeICswFZ76XjEmX
WsbD9AKVfyxF6yBLpl3idxbb8nSCT8cpRznX7K5+pCAXItdTn5z2m6S3Yk0OkiLR
P69xdYXt9AvkdT9fHoWJtlTmg0Kg5dXE59mWvh/gP4YAWobHxU4fnhnohSsVqc7R
rhq93QzioW+3A+0rS7H7MAyEeKDRmK7PBvSZONOu+E7/rnizprbp6wfYgv71zqzQ
JCImJCPv3SULaS4jd7cWgdcNgtQG/O7ooUJRA4nSEznv5JVgUBPghEycxBIfgWNp
ufzBFSGRg4cAyXkMivdXsMZh19iyv82yFi79XC18NRjJ5/yPyhbDJjCEz2kIHPcP
e6yok5sLXQ0lVQTWHtfOBUWQyMBF+JheulzNgCk+snoTDhrZP9wbN3/upQAgklMw
EAbEuDp09702iZ9hmcbUTmGswhO74RgfJNtdFcCYYbQEFMcJhJHAVkm8/JVsPOw6
FLy0XOxCUmadOpqKHxgL1kM6O9IxMW9Mvg8u0ged+cVBL2kKxcNwjVLCBtsBsb/3
DbKwUEbXMGgMWiOoDf6sgm7Gjt5jQNozwe2o36zXOiXVOwwmt7FmD09bGJcIDeRk
4QA19Es5MiCnOKcIC0HcZG2NA27csFg5plO6ogNem/9HtKFhC3G584ajlmJF67nn
Ukk/OtaXgjvlsKEgugmBrUewwNi64sD9iPBpaOCy6kzyylAvpCh7bgAwueOSq66t
mjoZs+ZLXy8pZuP6ZcvZhxBKmOI9Os9F6nVIUoP4eDo/Df+8YV/DZ8z8IiWhLAF8
+l0BQm1tnSxtJ6dw8gUxARDAMyTEoNffCZ1rrHe3I+hKSisgYGkqRvSeDxwvFcam
3vSNSYnjFDRUp5AKX7QKL4G9Six35uh4Tbh8oxjpAPlCJ9b3jwv/cXS6Z7RspT/t
WpSzo/l7YDIx4dRtPCEH/RwOZETZfrIzEfmIzPdl6X0gp/TiFFZmdro4ecCkI9eF
ewOTsNBagV/74nSspxtVuvvrcJiinUzDoh2pnv0wlAFNsTXRd/cr+YRC/cbNyTEJ
eUja5ID2DqHtyofXF4CBAeuM9q/xIhjotffkHdHVNkMrBiEwfrM3X+uMqxqiBMBg
pbZNK6AzGTVh8CqVE4C83C7FYX0SlK5+lob10xEEQKLCWoibNNAOlVYk7oOPHfyp
IwuShxrk/4DIBcB/FoNh/vbtRXWE1H+PCEPUBsGcNop40NNe/hZ9pT/Gm6DWybR/
PIDLEBxglM+efNAMBuSRhmRxj04HEejZ6RSsaKDpEJ0Q7l4P4TKzlZ7SyglG5gSg
UYJfIb6PwrPCIMf7rLqz2xzgFok/j8QgLfeR1NdbVDjZAmzAb2TpCOch3BCSkLs7
qXbjDyKdmP329yHSl9yz/bijK4zS3T+JMOhrOe47DPyW/7G8s62+cnEaFPKQc9Cb
ENWyEPPb5IfRW0+OndqcDS7KTDz2RjZhkp1Yvvkeh5qPH2D/A3qKzpr27DG7EPpj
QdhsHWCzr/vq8GO6VBx1kEg2SfqwPZsm4OkH80POZpVrqqOIQkTNjA3b/kq2pVGW
1RfQsketHXL0amYXKEYSKTsMu6urHcPORdIEm6+HCsCpuVBJ5y+/f3/Bxahnr8i6
kWDAUp9R0Z/6B9bKXukQAlWFqA7ecu6cOg9pneqwtlNWsD3NyXjnM9M9BZ7oQbB8
21g8t8Tvu7CIqoJTh+VjdiFwF0wGrganrimiW5HdIJ0soV1wGrBU2N75Yw5e9PJf
PBGk8t+SRe7kkMJ90eRynazOT/zaTSVy/hPA6PEvA1k6PTJVNWYZ26IdC8v96dzi
TSaeeuGe4Li4MtHC3Big2OeHA9uIuA3RwjUluyl9R0rEj8dWyBfHaGMlOyH8ipBI
Y5U5np/Q8Z0E/rMx5SYL2tA5lYggSQPlIAt6N7vzEpJIsO8xy+lzBV5+RjWCPuXC
HohW1lB1FI9fJkgWEJCkAVXBGeAfqLz3cgs+FArTmKfQUhM4+DNvtBed99gXCxoC
0yX7sCCZMWtdWXAjGFV2oSua+OlZfW1Aqhal9ldWTpvgYhKvxeZs/O+lJdmtuxtL
G8YfXvbW0p4/PvRFbDDmX/XUE4Dutfgv4as7MEWcnk11h4LdLggm4pX+AGw8Q87c
5S7YPxuA47itLy5cy6rPzMKMTvsrIpZXurXS3/OPOHnCw0yPdR0S4uoJ4lPPJ7cl
e27p7/RVr+Y7zQJHvw2s1McT3XFR49mGm2bBRbkkjosqirUGelgg5+I9R91+P3v7
Tqp1zSlgH93CL04V3KYhGpzVBfzab9G88c6SESgKcXsEFEIzx7ktX2E259LbjB6p
K32FESd/c+dfND0WHjYicYSCGfyUlgAxEYMKkhUUMNND/1dg9e2ngD0rqPt9Udo0
gLS5QNgsGK/TMArR/CudOEu+TYbzyU7yeRGA6uvTS538XeGc7KH3b5dDBKSyX/uk
Y5DReIgLVDxXOtX2dPpOjtiTrvuNdWB4ZhtcYY5m1584DJivvTniW1mAE3TzIqPS
MsaH3CGN8ZJRrLj2DrBhAHtOD/C8PgS7zVkNjQBCG6FxKsTZUCJ7yz5WO2i8Eefl
nc2JN+ApqCG401KJ1s5f7ssflZrcngEwOu4gzyiIxT/ruzutxLAUqsG2GHb6a8kV
c0YrjGuHILN9ByT1Trp4jIlGF4bAlU2zwJ3zVl5uJmf9H6A5PTdsp1nJNSgsSuHF
Lhf3aCG1TOVlJwPnXZjiv9r3gOH0YX7ScQVSDG8UprG8j7tNc2MmL6VwCA8zned2
F6vdyBscn/iBw8qxuUDryQtFbD3hvaHDSPLirvaw44pYhgWNErEs0QliwAhtbF9u
YNhNhF3pBxXk2sEu6zNVQw/TuzckSn6Wobvf5blVbPhoiU81/Ny9MZOW+q8oRUHS
ipblkVg+XuYIap7/+LUsSfFCEfr9ogeklKLumGZrT/54tT8i/dL0/WtMdLp/B419
a6H+omo4vIwYXcIBy5WN0wII35hYkYj0fKwynlOI868MJREHccDg0uuLO6aepoJP
lD/H97HKamyZNG8dzeRsvor+K2PaAW9OlbYG06O2MXS7ZLi1wBOWxNJkflK9Hhwc
nAB8xPQBEqbg7UA2GJv/AaGJTJ8JibTW0XdtYjFaSs7Z4+64Rv1HhVlE1ons5Rur
FNieugu4QUvIk5S6g+1L+//NPH8blETU6/73qJzRBiRb0+CckKDGOwS2ouESvK2r
ThPt6publkkBX0JiA8e127mPjhbIEhGZEVEZE0dBSCzmwUD63VJ+HGZrRDUEdi/L
0OLOhvPax/s5I7fz0ggobeatfix6Wbc35K+5gIzEHmZblfC62LjEFhSt/4xmWgNg
uaB5pHqU4GnZtFzjwZFjFqPlTMr6G5GXNIetzksIh1sz2pMOY6WJhzGFgd0osE/Z
ptrFFbBTVt07kKVmWV1/3tfXSkVBUY88q55VcNYuX7MZRSY6Wvof7prAUwT+9qmb
hy+STNrsn4qVmwhYWX1HWk9AGYXsNuBlN/Wv4ufWXpUFjLxiLZfyT5ZY2SKWPuzH
cz0Job6PxHoebQ036OAuFZ02atu/+KFgRMaWas1lG/XJxKb70tdM7lYXbmHv+bDL
65xilDgXzgx5pbGCSOPfbcJnM3zANEpI5ro9myNnxLPECYI1LU/8wwPcaa+ttWmE
v2REpzfjsMvVpqm4wzRKo1iK0nP/0cWSoOYC6GD49DB6l0qrzeTZOU6oJIO9NR4z
hT+8KyJTlh9dfo/31y3CWG/YtPTp1MWWvmTy/MYXAMcA53gILHs0SMM1nJo6bnUU
aRH3hsF9PryRRDTrfysjqXBRnUVTbAdZuLTcDAF9rS0mEk6fA5o8/MIC/nrCvMXf
FPafrTN6GqesI3jtcHs9Kt6qt5I6CRlvj9JUKCXz/DGhC+dk6eI5/fs3gVb7T9UN
UX9AaMZ5VY0hl1arE8tRVa3Zdr2Sbhv7gVJ7Gv+jaEpfxde/HXg4FvUmBBWmlkmk
zTbJNIkM7J6aUBcUYFB0WBMLf57ubRma0+Wx634DinI0M7o+6SIaqmuShOmzefUH
jYpc5+OqlEcTeyk/P0iHJJ/CiQAd/juP7dnj2Z/Q7kiEPvs0ks4TpXEnu8ptRQ4u
BYkEyeTt6pKevpuFfX8H2rh+O61qOt98dna0ZxcsP8AM1R2xqvx9rD47VNuebe95
9c/K3gb26pcs4UUOzoQuE+ofM1oWpys4h5InuPmMxNXBwstvuI688oIXBJVpRWoE
Z1yTaNfKO7AAKe5k5knO5ZPaIIcgjYu2DJQ5Kv4F95zm3HxgIQ9f4Wr54xgPM6LA
oEXLju1CRelWtHPShq4tL4/pDUk66TVtfLHJeF4KwdgXAKPlOmLxTtKte6jmx2XO
hMBubv/NPfKp1aKI6+Iw5NgmzJ+vFXnA0z72j2Hfi/o74fmodFpFBqKnUnFbrFpu
vYa+hgfXbCZ2Tq5714z7GvVdKqq6Jddj0ojy7X28LAokREzZOrujwO0q1O6L3gh/
ERjUBCZPeLGMyk0jX4L3Ema4boptgDbAa5AVx1f/5n8WhFeNyYVg62VBH9hd1Wt5
sYEgkmx/76jjcJQ4cda5iK0ibagLBrWB2nyMnxKvoQLNGdzl621zWfVweu43AWiu
rnGJzCGfbGiDBTLmdoQjvzBtl9yfbGG7voLY1KyxwykskjKFYPdVn8TdGFiwxdiJ
ZRMHTjM10ScZ0FzWXoY1FkSbAcbis+mDyiAwVZh5gIxlFsZgeTkt1uQieHJpnSLS
a3qCwIvTijiwMNJnDjirxjVYPyFxdilnxEHYfUBVFZmElHOZL4MepdPnQFtRYZDF
zETECTCGJzHUlFIENfGhkiVoZtJ8IJqnWy+Xc0Ptyr9w+bn93a/vW6MWh7AJ59m4
9WRtdSft03rMXw88Fafy7FuTSylrK89pMg6iZKMUnUuLailhblFG6/5bSb7HVzvP
eHSxi4sHlHU58h6eXpkIoK6ezO7Q+M65OZOxBZ82crhyqkAWdqq49mlK3quxf/TZ
kJFzqnfxwGtnwt35jhGOYzpinJN5PW0r8RoAc80x67MJTWwyji9Sotyd++vIHOKt
vMUuZ8r02jQox0YTtqdX6EYytqOlhlXTr30R14l98StF7jvfC1nWWvutKPgCVroB
6bMvVYABXTHAYleaZxC/HDZKBH4nkOM6gUOUCUXiCdjuypYSEit3zS48h2rLhoPx
MIa2oTLfr+OI8DuTlRna6Z06qq9+fP24YRgYjsfbveKb1X0ZHzQGvLLV7S0LEaB1
6OH3cAd2dwEIDHon9LwnvcgjRxqc9+Dja2hFQSKC6B8kT/3OJwmFEVNoyZHWDAQH
N6Dj1qMBTXhXAzoUyV5f67Wax2cgpmYQrslLOJZlJEDDWLUfjnJ7ny9dDH2Vkcqq
K52kjCYg9nnEQSkugQTWkwnRc7z+vA6aRnuFSMjPzEM61nJ40ljcw6sRTv8LwNh8
yVPEI5HL3emz2S+u4HCCEw6xtUh7J3h6e2YavOIUluVXVphVWYKMqbvZNTk1hwIj
ujAdEeXqozMtWK6PsPY5fZFk80W1z5kBoICDuHM+D6I5pLGaLYsm02Yl659MOTXM
wfv1+0FVG/DNc/GS0Qc3Mk8Xft30OBIyxKLrMWSLXUIHV6mpDXlOtsgPRkYNPUEh
w/7aQktybe0eLg8MpTErVa/6uSLE2HPiSmaAMKlEJefonQMt48zNv2sKSZ/voqd2
dbJulJy/NOuyIIDslpXtAqm9lKe5Ww/167c4p9rSMJHaISGVdpBHCWN8zEjTuIAl
QVETJiuR4qx55/F9Pw8pbS3yHKY0eCdgWKdIsmP8uh7pPjwHxnSCrGSeQ83G5fx0
0IgGo8ZqKvKK/rXTAXd0jJ7CNkACK0fb+PdfEykl+YjXdPn92WyM93fMli54TLRx
mNgNP8wD1NNyWUpWOJVEDxV3HMo+jm0MtMuYQEktiBO2NEML1mYbXvizxFeSARCb
0vbCQtIwqub5cjVqgqtpvUMZEohcynOW8V7dBg0c1ZxuLlUbuX0Rdhhoyt1eCroW
TxANMLFmeuswdvBxmmMN1q5t9GMSacwTSNVl6ayxvRYtO+AzPsImXu90OoEwVHiU
SQv1L/zxhNbWvH/NZLMf7OvhzOGgG4V+2ZxejD3JkTOnmkAAI0RhBKMdAvX1KIOL
UNHtZnuk938/wpZ9ewoBe62yzmsAqBy+cmpgWCwq8NFg/ypyQ+tWzimRa/Qs9UcX
nLizgN9Lw8MgGcXFgzX96GZzoAUOZHiaG1ZrDYPlUwCIyMiLxGQ9SLZXR7Wy3++r
lTe1BEzmjTHfbLsaEaTzChEJ7nGQeQU6yh9XcsbruToPODW8ecKAKNG/ebS6kHf0
2lMKOoGCQ9hMZwmD55ANPEKFF5CbvaPElYZZODivS9NDXfB04jKKouicyJTUWMpc
GqyTum8KzmxPB+K+lqW9MwWBJ8wTsf/juLgBAc0xdj7JjoWaj82yKLNcoQdXX8NJ
BprEIAh8oJNsyurF5jpp6YYK1jNaAhcS5zWZ9S1bXy8RaC9BGzkKW7+wdEGjFEmr
dPF0mZnoof8CIecegi1+ox7RFGhV8Y8YWDdG9CNMCMk9uYRicl2IIqgq8QR153hq
S+qptJr8jyxoNt4zc5wT1v+31LX161wJrvderLZM54iY3Bls937qBqjUphKa4XPo
efrh1ek0wh8QiOXGj5YqjUh/N/j7B+2tpsbGApxBicPFOlY/GXiQrhAIr15VGrPI
rOcemC3dpXGK11u75O0fcs7JTB8VCaHr/ElJzBmQ/ohkwcjOb7xwFqD8b3Fg4dt3
NDfhtb0ua+//9hvlbIKSRaldhvhx3yKRiKVYSi5OjPVEpyJfBNzlnxvgnzNmLuRB
biazhQSIEt7gnTBlVULWLa+DlB+Suqii7I6eBbr3i6uzWSy9UQEJ8QdsPKlqlPtW
GMD1/7jAE38jaZJDxgBnKvBrvtwZeDdx9An0/HpZP8wa2+JkCDZhagv+S7mrwS5G
I0QON2gABMBlnKo+A2V6mNhk45hl2TmFgUw9Jjm5aYIfz7kouGhahDQTTsjcnxq0
Fu0jnExL/HXkKDjgeXnPjA29zTUIQAnt439kTw8kPOtn89lFem9ksRyn3wc5BbzR
M/N98ks/xaFE1RgaOrp0hH22JsrDegXVczJDQv5+PJTwiMazfmT1qj22l0Y1gul0
2zGvWRUcb34j6HS5F5m1a+ai2zxPsODvv+K9Le6iWYRDCP6wKqxKoXS7Ovil1C4e
Gvg7NDlzOnlXBTD7FLQunB1okbyyK4sRIk1Gh7wX1NsplU+rIe4fAHyf0oMsf0VO
UPW4zPS53kysTIJ9xZGufMjYHVZ8Tp663TqdUVTHpiqrKrOvyYjLA2MXR3LGwJSf
3HccwDLNOXOkfvvGsWzC0K+2GXCFNLJSWvtlbcUZ6FIIKfvncDBRA9Nwx8QoxIpF
p0Gz29WPVh48DKydNBQL+sBJTu5r6ujOmYpq50CiPNzisRMQz0IBbNzDoV0p/Q06
v1j5xsRlZ73jwRRWKzXxZweMZWVPsRRV7HCyNNSUUFEtnB/rHp7K0Tykt+1Cv379
3gY7hxRXdzl6+8RMydPeSGlfeugGlNQ1qobdC8cYFVnAaZX+7U8OiR1Qdm+EpE+A
6Hx2TZW5bfjZmxaegTqXXL63GLTBupG7wSA0lbthLrhG6MsCHCgDuaPYlVKI5K1t
soWItFvgwbjReQi7/gYkqHLzgS+q9CG8bZSfaZeCSzgHsGIZ+m1Qby2epMag9X1T
sjfk8MiXDgXxcL8zC4qBrsJXfRo5foPAk6HM2fHcDEsiRo1rFzhIkVCg8RnBkbRg
MhNtqrMi7wIyz6FniXoeJJk4v9OLTl3A8VkRnxG5B9C2nQq4IdIgWisZmOq1R7uW
fI8IlQiRIu4XELYznyJZkxS65W8i7W65FyTdhUEi6zI6qyVkULOSzU8Sb5cJru3O
CQOe5XBZZgYrpH9HySDaEUKCOnzNuPhziR+x7QBWGmmr+5UGf0/UifDBTP0x9odu
RZhtsyzXGc9uFBVmLiJEJxjytAPBlSVI2rsAm09SooINjMc6wQT6fsA0l7nRzdtf
AfH1OKrf5AaY9DcbV8jyyFIR7uV7MZhBcBA9K6zkTwINvE37YC4v5o5kZ4RRTIMs
CiylRVvBzdeenyViBbxIJR046ZpqRup5JFuNkdvfff5s6IcMATtjuboQUsnZ3+K6
E+bMCpQiuaV+D94A9w0k9Hn2tK0hIVoyauRquaQiExbw3f0TEeUmsX2iRhSP9Sm4
USIfoWgsSJiFUVyRZn7FgXl11ophIoXMN34pKwCOH6nSUE9eZafthJimI+oV0HNP
DcwXdNjmhhVJJCU8sIZoL01lDD5pZL6+BF/jOFk5ovQ0SQ8NzaR/iR4zVGZNkft4
P1wxLembDHxjF27bZCDVv8lZKcCecv8ip6JV4L5tIXDE0reNYwzUZ/bq9IpCWhPK
zsRYohNSGdhElT0lbNhSIiFBOHJECFF/xEkldT2UpBy9m3o8Dn1TtkpTpziLpNH1
gWWlCFs9fF5kzxRNHyvcyehDHqf+IERX0sTmQIxTCwZ7G6hvbfauOfyOZwCEUvCY
AbHkpDB/104fAIkFgwwNGyygI0PRHboq/MYxFwWoj4gpryiaNntmvD30rmCCEPRw
1sshrPNhBsbzzBlcrgXoFNpqJhtNtLl7d0kqYn68ZRSOWhXa7OBG3q+0kSswyYc2
yY6YqmdC5F5nVFbPY9mHEi6FMALSSDG+U+D3w1fqBoAJ043qsnqIW5FYoC84uEiC
2giupZBGQ5v1bOm0kBU8GGnPromGV/+bNfOeccwAfzLLirGho2oMAnPTg0psc/zV
nH+tsA1ACFsgfDmzzjB+NUDqA/32R+NH60Aaq2U/dTnCbWX2f9hlX2aO60BcWk6v
0Hf4OXwfj8YKIvcATYe5Bd/p1O6uIT37pbyoeON9IYSjqwh88pIi9M8NScVa6xN5
EFb25gFHnBjL0usDwPJwusf2dr6rJEB/TLYLg87mIWWwyJsXq3LpBo0jQ7ASmgMm
t4XK2cZ4zWYIlZhitUzbSYyua4zdutKPd9zi1mRuh5kuweCXV+lxZq0vDKWB6COq
Gn8MnynvvGl7FO7A04UoTRQp1oz4ROXbQHfZgx2E18oH5HW5xXJcBOfnihuBDV5G
pJKD+Xb81+6h/uMSw+lztN1iGjmBk+n9+DKwBQeg27qIG9N1B7CJbXFgFtV5NWlH
MymDCLV3ssHfQ8NLsmMzVHZRW3OIgIklFLQGgpwIrhZWtCgL0WW+vOJdxklWMzph
h9p1FRMl2NLXvD/E5wuzkUvf79iVDjThMe6VMd+kRtKj+4B4InvJ59vy3Ngk6s5A
vwoneiDWUlx6vZOU6iADj84fo4e4LWaubGjUSCpOBkT3JqawOw7zbvdkmL1bvWFm
bPIevpEW5Mz/fogGF2A2QM4OZ3beSlfj64HUru9FlHayX+7QXDTvAwe1Mu6MoMiv
b3mYSHYK8YBeAJfxtei4kXRxECq7PaTMExIRSWsVqYwReJYb/QHBdTvDpquD2A2b
Z1APkHcs+VRbb57efRMN7fGGi6exBh3UhUCN4uoI1we8Ml8pF0QxNdwdrIs1NIsc
p9zS22AhV0Lqx0B9SXTNGML/v2qk1Lz6qxWuTlA8xSngO8BgQGCa163dMVCDs6PL
40FY8tYN0QairL4FFIyHggQ560alG5QwFIyTXApreMGU6nhYYik9TnHgeZtRve0P
unChGwwh4PKAcZEoBdZfhEYgTPaTKIoNudrA+eL2Rm8DpWBn1HxV4JLmG4MsgG7b
E4ADoTAJhg1RrWO+JbHKqSmq2GrF3pR8Qr1LRTz0hh4kTpe40COvyrTZrCPzvBac
MCbcDvy7M2AuLgC3dqEgYmreop4P9UDCKFRsnXTkIOQgBvEBB1iIQB1vyEW5nyrP
AFONtnMHmjptLu+T18gZ8g//3Qys9Qfya1zs9WmrA+uc5C3HQwOolhTSLNK0ojTs
Hpv4rH8xoRLH2ksQVQLWusmSjtlmbHl2sjWpRQ/e1r3YP8DZ6lWn+wAE7ZmSqFuL
+bNtauaKVhxDpGollu33D07m0yQamm0l6LriyWCfV7cQ1YURyvGXLImQgbivxA4V
sCilGUl+jNYh8gkTRq6YZ/5s74HE14i2T9pQCNC5GQVc2QpKNQYxC7lgUH7s7fei
2VAzI1l3Fq7/bV5Z0SU3W2ShFbZWz9BuF3Udc8DYr8w5CUBRfpPzmRyEzUM8sIVN
7SMQb0hLoeesl7GMLS8qzAkNaJ/Faw+iSpa2l7yfNjIxM2Owk1W7UT0sIkCqqv9C
OdELTTzzLoLRDFvL2Eurnq7OITAGOL3B9xVEfmxu+12o9AFaZtxlsvUCSznz3Lyv
EE7TIbIPP9jwixhIN4RibFfbGIz0Cp2xBBUS0wcv3/RllRr57D6bRKREJUz6QMzb
gwiMxckT0jG06BFkwN/po+oMgPjRx0hYs8vmezpoecHPZ64tJh4g9jron/NL4SJc
IkYlwIvUDliKh8HqtqoSKl0EJhaKYw1p/7+/2JiRmmtPUMHWAaN0gPMvjz5MGQ9h
+tTARspXzZqrHpo0vggGogFbYbV8gpHo3WlrGETxZEa8DT6jTO+gSiMs3hdQzCRp
YLaXi+j1eu+PG1HQWSWfe00wv12+Cx7Mn+2DQ5LysFEzD93aeF4cQSVyy3w245nO
G82N/anEY6BMfej6loHc4xhUHxzSfSGIBgrTx5A3uyJnuuBzQG0wiFt2riNlyH0o
M2qeJFqEjzyv9YnnSQ5I1/YTjqGwOz04zfHTKXyynXiVOzCOsq0WRUuw7eZReK2Y
wyMrqnBuu/d8ZPIcUAZY/kU82zTgdV+0mzTfUbrmuTYFLRl2iiDP+dgAK/YhA67U
75wnB3md7pxnpLS8xvbVGPqPf7LziBOzDw2wMlOie/F2H7+vJ3/f3FuvaPyGJ46z
vHbzuzhd+zmbOJPWppLgvZrEKc12R6H/o6KdiaRJ0IWxl0ug/8GBgtbu8jdnkH2t
kVtNdcZSlUZwxngtI8wBYtPhSux/b1ddTSV9xqDSuAPZK6DTk5/icLYbpn8/fcq4
gMdAKBTkfQpUGZg36ZVgw97O3u0aE0wN3BwsFdfl63rn+Umey7INJbAI9kSjNpp+
rYEwijDFZb+ps5en8HmkQs5F8Wx502JhCOahU5gGqrJD7UoE4qLbY1A2v2yIgtRd
2ui+sao9sbFkp7ZhFRaqXoWszmyswqPgSi7tgmbBgc8DHYZ/3ui2pUW6E2GiYMUr
JO8AebNJ1Jwy8avpFj1ihgmAISyxMTwjIObrcw1lRj4Y+aN8h+ZvjpDTZqftZy/c
wXnKbF7JtJHzTQylyZyWgtLtWnnkkQ0WknW7QUEZXYI3sdU9Bk5iQp29Sj/NA489
u7gg8Kqx40/fS2IvS22pkwMHI8OGEcSCcDyB8yy2kjrsZj7IxT7A1u9Erd09gvC0
busY0IX06plvzizV2AzS3oPK9Om0e8DFXUB+s9Jv12lsbBV6ixF3jpXOf8LS3QTS
ZngNhbzcmQ7RFbUde9QNfLXt1FOalpRF/NRJJxMfzwicdvLzXNB25eewlCPIIh88
CPrqcT/u/jwxImkNRIkKkZu015EKlUyOKH2wkRYeLyzAtI/VSzpDply27/gGg0t5
KMIpYmz2fxM+0fwGeLVI8PNypZfSGwuExllBTFgSnmcBdTBZnbCodPSG0TUIB/S8
PRNMONcHDFaDlsdZ8EYncn0mLze1sh4K+YkxZ+IQ4dr/gjX0kpUtSOhJY0GhpFip
WzAmh+XqR9jFqj1pBZ4dlB+PEoJhmgihrxAceBlOqZpSEju0NnXMH4qqmDAmNufj
IciNz7gdkFW5oB8tl5esT213C5FIhURXFIXoam7pdvyN/m1vgNuhS78Ewrix12w3
Y81JbVwCe9oOetENvbLbATsMBgmZMHqeQjjHA+eR87VHqzAbcKSFjaMbkGctILjW
s5lW8JxOY3psoixbDJZc4r7cuFruvyjC/oltMYgquCnEK9dFLvizYyFat90L+JjX
XbJVhQTm8BLoTY7c3Dw3udsLYwmNNsuXcGroTKOBNo7N/35j3ANoQNOlDNWwUwop
w17LZqbutAW2KxylslQoGyLgjdHm0T0VY3vXF5rgAGNM7XD0+K1p67MDIKUkOq4G
zuEZ2IdREEe/xbyo4IPtopB/Ja8Le6XrP3Aj00WNSO5FLOfv4+6MY76N2By1jC6v
1klmUxGmn5/nA2a6lySmS3FRXCnLo24i2rzEMMST/lPqo8dK6O4zYzwjPJ5z0A7S
HSimGE/SBYdBpKgdtcYZi+ojtRZzOzrAsd2ZkgzVDRD1jDGTis7uE/d5+FF7x4+q
Rtz6gO6cOB0AN2j7VMhzaqc8Ukfdc6Qh0p/YvZTqikTJdhS5pst2oyIsDjToLli3
Qpa7iT2BN8JLdhAn9kt9rGaTSWFiJEi0NxEtp6OVu07huesG3slZY8YRnZ4GW46j
pqd6ETRp24iedQpCbC4Qh58iRsuQx7QIPomCMudc3xMrWgMzptizrlEoalOmCy3Z
rHq4WqteCu/U1RKzCzYUjBpNJ5r7E3gxTbmio8AX16OMJ4sg1ibJM/o0ZPyjfVbn
rNnUg4s8JJ7lWmzXf18CNfz4A0dwqz/SOjyIhG9aXXRQcBseaQb24KpELOl8u3FC
5Ku9FtUgbBVP/ZWZZMg2YSUPP97jM2nz2RbvVY/tR87gs7cAQVTxtgg0SSACUQBR
OqJ9w6z9EO6BEOpZuKsXt2Ezw1NEf7hM7zYVOs4Ac/3RRfQtJru4Ye7Fm5HZ0HVk
lT/Hcy/Pmz7b6cCmLmGHGAKHzb+JLX9wsRAfY5VjPPaWzeKeWesdnZjBneLjpN2z
dCU2PhmAZls4Cjc7nET32FzddDcoNBlwcnzHlWuqQd4NLo5FcgCR0a4HjLqH1vVF
DNpbPnPYE5nE6HDZDTfqzZrX8V5EML6Wi0b5r4mVlM4ZcB+YiJ4ciDaNzteJjmHE
YJZp9Xg+1Cz1bpc30fOnQ5CrWTsh1hN01I/JET8kgc+iRRSFlit7ULde3hLHWvop
vKvEhG/TcUjjbWMxoM1aZGaZvUIygEyAwWmRebjrJKSBf+BDCEcLsLO53PgxBtBt
EBkkb0fcDIhguwiz+sRzUmvr6CpZFQFVG0WobdwtUPYlktS6TIf1hHlN/zGeypWE
FHZu8sXkbe8Z1KeEGSmpUTYdz2K2XFpOjINRDQetCrDVN/4ndAW+PIRMFVVudEGB
G+o+hLQnDGwsNny9MswtzzJ1Sz/hZJUJiKyD9mMaqNtNdpGVGgicyvXlvIjRMCTO
AavhFv+KMOxMieBTqXeHHJaef1OUuyoEeoyeknviIcLRD7Rgyq18doXIOgNz5jLT
RGvxmbCSPJaIBi6aIfr+X4HM46JyzrSb3BnH+wfMz/kFwwwu2rWlYiznShT4ix2o
WV+UBFeWk6LKt/DG637osZ+NgkXeVCHvPSjK6rwdV7zgPf1JjVFGFw5md0u8w3Ms
7JPiDXge1CMB4INYeNsK4vZtu2utEoMHHYW9tG7AIsxs0e/a04Umpwrambu1HTj/
9W/+Gtbp2n2coTuhRpVMzcs8n9zIeCnYg6oQnXITnvu5LmYG/Gw+9Gtc83HLTmTg
SWNKWKhfxOKH/DnLh5O77z6AvwqcsY2FN1kcTp6Q3b0bxW21ChF0WcO2jaVI+zC1
mMAn/NvIiVngxODlQtI1PtC36e5hxy0IK9gWFi4WCmm6v5u4HCyiUi7RnaY+nQrA
lNth7VC0GO9FORW/VXkzHzQk/HZ34yLlsyXiEbMNwwylmcfOZ/YHg+NBVJjFEMNq
L4FTF0CaFFWW1ocxm8rPUKSi56glIjLAoa1sKzm90iG/q60SJ2xegdGJzhY779qa
09fg0xKQzoKDwRvv98l0H9xt+7qtrkuYcM4BStdhFQfWOwbtrsJBrV+yEzZPOrsF
2EjF7Y8OPoifzYcaBuyFw/PaTWQlpX4tOngjFogVG4W5S5akGo2r0S3dAt85Fw0C
r0KOnJGm/VJ//dfqpzDjmxz2KzMNKkKrbaB154e9Pwc5NMsxqOfeWtdr1G78w/EI
MhUpPpG9y+JwAxIk+6Lzbn7OSlN0FKIkewBtNT4RHAL1IFXntNiG6rUT83JmkjRb
ldhQws0hbxJLk8d0m1yeEAxJpOX4V6Fb03BsB61/6i9gUSQTAkZ4yvYnyL4/9R8X
RqIAswB/YaADaOTdUSxjRRT7KNrnI6XVMq2ABg3yVvTyoFzcpDxCgpskfduGaYJO
MdYZ9pTBSA5LOwisQk1uiDHDAbAb0QARTMGk6DeOT9rYvKoVH/e+2QkVSnMFW7ey
JGgcsFJMIf7Bxf6WkYk5rOMTpIV55cNPjgfvm55IsSzktF2SCAmZI7fL7zY18yQV
IwS/w7FQSDRpJZDC+3czb3FH0w2GjbNKAzO+dqJVhcUXREqeneIUGvCCnOAMfcdZ
wQyMI5jc6d90vJHUXTXZVyBdeLXSKqdUZx2BIHcKM746VQdqvfW7Y4y41p9JhpHD
AYt7CWHZtD5fAL0Q46vTHy5gWNBIw0Rwo20p0M5GruM4gQxC0IQeT0iye0SW3v4p
0AEtLUrVD9Ari8wnCDJwsYO1d0/+orY3a5cpESBYwGU6xxI9xtl+rDMz7v1OLeq6
GIEQwwtnVwdotdUybWPyrSExMC1RT2B/CgrYp4tlDau0nDu/Vgaym4mpDRr80Oia
Z7h/dzw9M6116zYoF0g5w8lb+CcKtpFuQWKtz8Zz8DB46KKEcLHKTJdn2HfKOzgT
9LHkLNIczs6n9LhzsQuOOKS7nB/m3rUt7vd5qcsboHGGEWWFnl0kEGmDoX9WUV1r
7R2y/mO5pZAXqSdogOzzyOUjn2/y+Yjyo5CpebTWxVy7Th+sMcqEmPetKLqyH2nt
QU7YrZyc1WSWUxwI4ZyldlGA8NW9VRWh3/+J7YIzpJPDuaMEwxIc4oQFHvTN2L4R
SjvZ3F+uH94nmHQmGxlXVTFO4WHkHRf2qJCiJptM5SsnEvpZsgqUHOlLTWeC7OiV
zQjpYsm7c3kft0k7EFBA+vVx682tx0yY1k0QSkSQIBk3lZCVYYMzWQQ0LIZk7p7f
KBhfmUMH1z1buIM71Q8wCWHBQY/j4ysC3gg606y4e9Or+EmMw07y1GB/7usmCM9t
aVgoTlwO+zoBX1p//WwGSejzVGCPZBDoyXeN3IEQkOKJcCyvhLFbSt0f+aveZA9K
pGQD3c+Fi0dkERKHSsxyR5X33g58/WQQI6FP7Iv7A/P32i///hfySx866G2vP0Ev
CPY4GeVCLKcyLQ65Ydprmn/kk80Wi3H/LZtmepRm4bs2xxqGFG/ZLg1ZAgubtKEO
vL5GDxUQmm/b4Z7Bs/HprnwOGDTfUKSBmIER5fFEW535nlld6a5QRJHwijS97Dp3
weQSIrKKqzyyeRVGI/79yhn4YjjKjY3fgUly4Dj9+eVzrxlbKGh7hV+UTbVCuUr4
D9tnDmljcbnu4SVacwYixe7gIe7dsSzvw/a+yA7pWl7zabmZ+suv57rGfczj0GnK
FpP4Zc1SV7nmKfI3Da6d3umcp+cwi9Yk4GPRF0JouaDqB5d9Bfgg4HdUsYPNkK5e
ZXU+ZfJtkrj9F0y3+QwBEnIfMjJ1CEvib359HS/t4yRXcdlw2fpQYiIzlVPFXyEy
b8qh2MdK0lbkZxESS7eIc/kX0+JkoWS4g7vacc0b0YKwGsi6uTAKAzBfsZ/DkRhR
PgyWgeYqLn2RLslgdMBSEj/15pOMawW3OMgOsgaR61rEsmg3Ba1291XCL/Em2bYz
3uIoSzVcWs9uKelliQsz9peDFqNvumOd0O+xPvH4RRnU4Rpzl03QtXAYC0JOzNHY
S8zOFa1SYIk5MXJjCLOAEKvLxaVHJc6OHtynUOdANdR6QLgQoPsskymko4Hzwe9Y
cAuheAXQaiBGZ34dIsCJ+R2QXs2izjOpPqTMwvBl/Q3XTqe0q/7fNy1hYZB8RrMj
SJWG8zqd+CrG0PmvnQ+ZWM6hdiBKmt57KaEXKfdFVA6+ljKjItbq12Qln7obG2sg
rOudqGjlCDDEfgwMUBgmJT42IJsx8gJxRm1CemvraCdvpOgUUm8vjym220pfko5A
TfvICUjwQV8+EMdWOspPZQc+KV2PlOLEHO+RZ6hv5bCBk5X6XmwoxGJ90I0bBuDb
QccgfVgi26Fnt6aIceKgsB/Qg++P7N9dRXfH/n+K3lHVco/wtvR7VAtw+dy8PYzD
k6wycpIo8lF5Vkz6ek29SXvCbK3eT8QtFd73OXzn0o3szg0rleV6SMYsFM74SGbS
lKqJvsYI06pmJMEWoXd/Pw7jeUwjaYSL+LPu0aLQTQ6kc88d072VotGFJpMAlbWP
qB35CAlYrd1CHmLacT5JquTyjKLYwy40GD0bswH47znMHSnevCyigSdYhKRACeiN
cNrkTyaWBUpNcICeK9C2pRSPtvplc6crPzzgL//UCOA5iI60iWLllkJSmpF7Gss+
LBmsy/AFTVPqKK/9oCH3MxN7fHQM/3/CVuifmCJOciTbTXRWMHh3sb7kjcHrUEus
hV4klEMOE3yyZKhNvhpGcQtziOnKKrpMnN1Aqg3qLKi5D7sxKl33uJ1XNFC4SJHj
miIOTSJ5kcqp1nWuH1dMkxyH2BBhsUaUaNxIdzvstSAwuQi9C3Bshmzu5pvyVZcs
dI9BmsiSkflDxcC2FaSaMxQiW0bqF4SEzPePeULmciwm2m8wprYnaXxVWGYdRjMR
i3dDNlfcnD47gV7hHSEi6R+GK4odUAStha825YekeyIAGfkC2+RPweVwfIyL0/3B
hAnuDqOloNOtdmBlMhLR6RchRqOJx3B1lRZhUlufVJURal60dw0YHs8fxDGyQNMt
CqjPCd4kgSNXN3Sqv0Br0DEBfQuXi1LxBbNSDbjf1LGQ0xJ0Yv0hPZWHv1I1HlfT
om19vAr+qga40pmWurnkHpuVO5BLhFcQ4iHed+gMgqxqb+XAMyd80OkxyOUcYevR
pUtrqwwomsLISMWzFmfIFABEuDfJqNExd+8mXohSnHd5FJLKmSQPolADODbz/UJY
pd5h9hyCN3L5FBOPZgkgDv9ruVCAYr4QwlwJWJ2pm2PskYVKxreQOnFCx4HtEhcC
MJmpREzOG3D7qq6fcPJ+PedDT1Q0Y1AXhVHPSUBJ5YRGgaliSxaPx76nAdSSNSxW
MnY/NJS9Yv7duk6ZOfGbN3DRCz81KXarrMdIFw3DbNv7x69pAxa6RMUZ8qbAS2ix
x+8JW1iqoyUSvj1t/nW68d2Vmo4w0ChYqe2WdBrLsTqI5GX6rBYIogyrL5bf6MUY
Mjn2Y6GLijX/4dxttTx3GsjQJC2pxeFtjaQCxmwncxFkViPPm9EAbknEFcM9k+Hv
7FkBcceaPrkyhIPV1Dj2XQtuHDm7GdaSHbbyzUq3f813kOQhl6R6jwQ/B1dMx9pU
OjyOZiKgl1GXWgy6XIN8fFT0R471Brr6CpKCBtnu8HaJFWD4F2a7UJ59PW9IMgl6
5VNYXhsMAIih0dqYAKYZgvRZ1GhvjA/dVRY71zNPBbYWSYz0PwWD84xOIGo3yU60
UvPP+Qgmpsh8XwDIgenfmOSfVNCgZMPu2Yoaq6oeFdmiMZmWuXgll+jERN1xnRVe
jrmMWqjUuucM+eGgPDKPMSvGeg/qo9zRPwrhoIa6sCOfvvi34fZ7J92cRz8vPNtK
DGtqt+7A0h5IQD0rNlg7aodnmS3wtDTIJluEcucjyAVrk1ZFCrn3nrRWsFp/lpN7
l7cSgU7t2eZh+zUAo80N6ga0qvh/DSPGQ0KcxLnq6vUCDLNN+znBywLjsMzy2hlH
ew8zb4Iiwmns91Cy0VRqHdZiUv1CI/82zZujfQepmUnDpxkBIDwbwHNeEp1aQ6lX
CIu+GW6av7tUSnnRUruIEjp5dHxQ/10iio6obkl157LF7VgrEdvrGE9gYYL/KFUw
5vrkqgY14mlgzOCAdtifWa1l04VUfhSzxDIqeUqphy7W14oK7XNvVXPOhdDXCxea
AtHwJxglTRFhm9WSbX/k6RcLNRv+shbws9mIbXAzQNCPssgC/FBKdaf7FiQQlXpi
sQf6OcSP1dKGSxhHvtoFea+RtMjlTTp30S2OFHpbQHSV0kVmbEDOys0PxWJ2zzUB
HqV0ktXoaeARnytu+sqsBz/Rm4Lih/s3fw0oz4lToLw+QM0BV+E0X+b+FAoVLzCf
M3ANCCxmvUTyeaVj/k6Zh2ML+3uuEvyokwj6gTvViO6+m89tK8JUIDjtTpsJVdsE
JmUwfvDTVjiOQ1ZjQ6EpZx51+auJkqds5RzemrbVRoF43NySMRCVIgIARxfwD/Kl
G/tF4/xnfekoRKTP42Gr4vvEwQX1/8PbZ1JegZEhvqCckIfQv+g55MaCbUcXUO+C
3hCWwGIreFa1H30qlGt5uSxcsd7bRa44D6jaV2rHMfuzhjmABUqbsgko4HTIOZs5
mD0uLXps4FhqNCYzCJHH9Q6oeJkOEEqg7MX6iXGCkhTJ3Xalu7vJoqyHp4Lsz0cw
YaFOuKS4F1QZvXuaZSIlOQqqilboV4N2cQHT35DwUqmr7zu+KRlNtS/+4ujvkuEZ
2WWikmEH22s2fYc5lP3K+t2RoyLYRbeA2BXL8EoTeB5lEFcIBDx0e3hPAyxbKmuX
NvBylLx16joEj5W/i2sNG8MgDv5nU+LvMkQaJEGnA6ipGINLPJYUZ3qPdE62XiOj
X6h8PKDGfcZmxyAP/kJQSi9q4RHWGLkPw6QdmHZfHFcMvO3sALNzjbpEy01eeza4
i7QcncxXp53LQr0VxwAt5myFxjwFR6/VaTDfJ6iT4XuB8oLO6easYxC+5DTpC1ob
cLkuSjSfP2Bb1lDyzl5PI5Fbb/ma52/0ICrkO90lybpw6yOSLVvA4BCzTGPjPiUH
o02SJQpdsp0z9dKsxoMMVazW/LFWJLlV3WTTbq266pwajN/82+YoKC1nt24HW1TJ
uNsROoDBsBruXir7CHPKoL6sl9RTgofp+4lc4tYffdjIjF8wSKmak54243oDmRXG
QmmO/kWYOzRZ6SjOK3+a66T3BoZInHg7oMV+rEbakQxC3Tda1nxitTCfSaNldJ9q
wD8qf7ubF15yym7F735FBBL9yfBCocioNoJZ/1lsGO/fxdfG/tY/wLchqqLfwlY6
rRYOqbxcuVP/ZXWpGWDiSiP0ft80v5Xq49MOgOxbFazUPyIg0dl74k5nEpgYzlPb
yBIcm2Kqt1eQi517jbhK/3LmDZTgXAU3XLyp8hccm5Ut3GhyeJQ5rx7PR9jMhd74
OcuxEdrH1KfXYEoMat3rrBzQlzXQFAjfhHmCdQsEZ+ePZ+ENmZTqQKfpCgrXytbh
KPu4RVD+UnfI2gSH1TcRpgYzzqvjERIpq022o2qoCh6cFupOi8P3JW53a42L/OES
R3M/w5DF90403QQfSLakbwef7INpy1qvZ439PQixQOMuOzK5wxs4aQGnUe10Kk8M
LO80X4t3Xlqdc3fbBlg6SibVTLHB8mAZwMMJaR+kRsQKiqbsxvHWRaM/YeHJZm3g
PY3mQ5vdEvTIPaKX3e8x4D7vUwB3N8pGk8I8Qacu54Mj6gA0MnLQiadkypGK6r9p
IU4HUKVufp9nFDxA56mqXpes31KYDvg9fqnx0TkgA+B8N6ljHuMErASp+r3EyCEu
krIkhNiIcTk1PfI6fEcTX/SHEU01FTSKn/ZgRPyGAdheuoMEMo4oYyCB/sf1Mofn
9jidu1MixeevacKO/wL6C3PPbBgqfArfn8rkzVWRIb6PYBym0LTTN6dxdt1p5dbl
IeWiZJJFL7UbV7PEjBSluZfxxSgfnvAt1QcqJheHY/6syQq+LZGz+If6KgcCElER
K187TF7UotYWAqtE6mojwlA2l/G5nyNNWCnHzYkpu9/ohWsaloczv3BTvSGgngaT
epKeXL072en5K9muqPtD/z/DddzT8j5icABcYE8oKYlON5tzBSIgP1zKx7k3dTiy
V6T9uHpervW7A+aGKNAlNIqGty+nu6wRZnhpcJf2B/pk+Anqg5a4J8+UKdG/PP75
/my6SU2Oa5FYsROq8+ZfY+gog31EQjiz3oBne7pUvS1hcBnHoJPmTSCJKT9chP09
xSJ1k8G/Q5ly1/nd6Dc+rI6yyfw3P7b3T+Zxc/DOAhlwVC9t25o+MAICp6xaG5xz
klRUObBN/HJo2iL1YriMo0tNk35H443vOz2qaI7Y24p4t3Wo/+E5zF8EtzCi7XE8
cm/mSo3+lW9EIPKN3BDEVSBqCMphcUR12J0i/JCvslXB2rbe5zc77FKUQo2jgEup
dFsCDWCSKvF1Co8xl2RYHYzjG5BEq7FwZ+oJCxRWk3PuS5n9O6zwkaDoqXlaQ/sG
Rx640dg1D+4/osJPb0Kd863eGd1BNkfHWNH/lQFhZtA7MZaDnL1oWKErlv16wrJq
Xs1V3skgp0ihPIObC1k3Q5d7/F4Gl8d1wuxmatE+wNOCo8RLyzW+XiJa75dnD3+j
r9UkKoRvoUxA7b85asrVujBAjRa+0XZS0YFuKbQb37gFr8jZ1x0f28fR+IEZGZ+X
hfcVHYeG4tkjE0pey6lbsX9Yz6UYYXf/5hj4/SSkJyoWCI2YmvRPKO7fIHinYXhv
MtogdtdG5cxLW54kXPlfIhadbcZUSGYdOQyN8oMIeEGxcihEeH9Bwx0+zThCnS0G
1dZZywhZuGi9IPfCHjjMG/LsH4D+iMNhKtFX/e+kC8TpI9n+U98VtNQE6yFI63C5
foYSZ16gmmSBP4Liz8pZrGP2/CSad2xEonnSXXxhGeC3YVtenuFcdbi5ELz7XjQG
vLz0XTvkkpXgcKmub9zW/bDw5/Wbi05LT6UuamwgviwqlRjA0un2FEfcb6m2B5L5
vwH9Q5ULtOC6dTpkhAmszkqlQVgC+ZER/wsNL8KhbH/6nn+uYjazA8428QmseIl7
cO9aPryc4iKgkxfLTfEL9gY8BswNWJzKHhLZFbcm4DpBCJsPMKor6vIv6ghbBvVB
DKs86gDEYtT0ONYX1o6a47UznWD95Pci1hhFDphIwrqc0D60pvQbpLYTsTpb+zJp
v0skdLHDNZVSFyUSIUjSTvPP8nALc9ddD0WR/bZbF4o38QrIbAndSE0Ktk1UJ6E+
6IRbAQVgkJV7tvjgrnpGc+SbBLky3SF0/VUa2MJmvYMrDsgHFbb9JVUDF8oP7JvD
6fi8bcqE30Xdx/KfDLgLj+Q+Xj3KuNfxN4uYjtEAt6N9+BpVtpEXUX0BzNJYOtp/
s1oSsVpC5FGU3j5TRI0tHOKCBJYHYbAjf/mrs/fJBvcZ9+gMovqZUzBooCUit1GL
GJRa+5gOSraBIsugzkQNCpMJIASNVwC8zi9hqPbu6mJTMc1qCH6c0dHRUJmqvCoT
qD+Pi9CjTZylErMV02dWug/x32p8TITZuP3C+KRzl69nCQ5Qq66lggPUWPHt54wz
FFg7nXRPU6i01vMXte+U0lW0V0was3EyrS7S7whX+p7D8TV4E6edSGZ+ZykAdPv4
KFSHLnL/rabKSjFrJdeweMhBFVWuV5NU0q/Wji3053uay9sfvb3jpdI5udsA8gYb
WbsAsq0eq79hRDGqvC5fnuzUF5V0FXO+QzAhsm5Twqlsu+ZbdWgGgWfCTkeKRBQr
X9lINpRVV1ZfItfuBW86l2oLwUtWuDdBSmmEKaJnrofVT1e/OyHZbXCH9VGzefwq
J2qowT1Nk72WxSeD/7caJp/oCsVDU5e7kBsSnqRkWF+CO6WPtdDyKrIBF2mDe/VF
brGFsL0f4Xd28kQikiEFJTZRA+WlZsFj0pSDHCGBE/0KGyArfThBeGhDYULBDaQE
bO8mWG8c6vIMiSd+Y1T8Za/kqJDgGtz/jdL6e4UPlJfEJWnglSR7lsYnBr1nuj10
Bq5+kKAKZH3xR2HO5pgx3KznSVjcm1zzhUYlhEFzKt1B4FsKmtfz/I7D1JxSLluP
rwKbO1tM2VbghU5xCPtks8+suUeb1sCR1cmQ8cjw/E8OduxFFbyuMusc/dtAXGqd
BR7zNoKl8yASKUjUwmr6aU1jaGw3tyswFn10xvLJ+U7U4Li+siyaOfvVjeACp7kn
+/jjyU90z7WE8/dHrQtrGeAZV1+i+EflA/owArcbMK7ueUZenPjLIljY5HqrvH+k
dQlxPBdEJKMdRnJj5OvgshwBaW0BskSsQSMaHJxEQW7Y/a2qyPnm5EfVs93IMx9X
sIPtUKFcd15KSujKDBYdY/8PggUu1DsRFR/2ZWMABFJInX4zb3SLWKvCjfB0kA/c
uZo7ypUa32fgRr4U/TDVGkDkThJaRyXsnewLXhPAnSQvC/etwGTA/5MifhSHkuA6
y+F8ksthMMpu9C2NI1L1cjty8SxaAQcDk3aYVmwTob+mmGjc0tlH/J+FEBtw93Hc
UjzMUKLJguo+c7Rx9w5DTMKJvyIyS+T0X54AvqdoWpoeF3GXMeVzRBgwAPZABn0p
iFzcInOcBSH8HNzsUXWC2xIrXMuLof6Q5KZxuVIGaC2NxxeIaDbm6bcaSnauta49
zsvS3p9nKmtv4h1LIpqASpeQOsyAZuVEpqIZHk3G1mH/iqH0M80rGKcT2lRcEF4o
Ck5KsQoCGj6Q0xDHA2leX4e1oMogePJucQ2bgPYa+T6X8PAotDy5zVulVjVArsth
WKLpPiGkg2CAf+FTQkeiPmEQMPDEce1Lvl09tv+6Y7qpCOcXg5Jmf4ylshw6cal5
w+Os+H0vxubG4uFMGITbc2fAlFonVn5h4hEM/pVzULIbAyOwRP8xMwgd5IeCxLDm
76IXvbqn2u04cqz/VcFHler5HUCQVm08AS+QWcWGUh+5YecXDnWXoAUP+wYvcaww
xIn8TIXscF0xeUPjHGjiKqV+E1PM2/ttsezv7GxYBkxTy565PPNI+TxIdWLcW+/W
TXx/QSIxLjVfrgU75YFt22AOkoPJA+DNFAm+a7/lrZduxi8pwRfsu9Q8243xR6Z9
J/+OrlvEeBBMwD+lEOoCcxAf68cMKKcjMiNnGtVgteUpDQ0FYSy6v7OAXL0y0bFL
wTFhqDR8xW39q1oYXjyWN7BZa40ZxkMuMt4DodwoRnfg5AAFcIaneUgyr1YdZJUq
E+x1dGAbh8lnnPhTtTkvMHYcz/IWO99uJsQyHkjeBKakdWX9mySd7kcw5oPpWF/G
w3LmuLZaRtB6DI6eI9EtRQJHDvl2qFXnIKb+enROko6Wy6m7kEIFkM3qFyyC/fNq
8v9P5s/BqEo8OD/7T9EYoR6czR1aJTk6cfYl3YfDNJqYs/uioOnGXe3vYDC3c419
+JtZHBF6fuLLinJ7t1nssf3zpMSZl6fzZFWdPbRh1QayU+rOeTXdvE4N7kX99R57
81yZlwVNBTB55bBGG3QPTe9prpd4cpAjHZJT4puJ3fJ73SOzQZM1piJBQ7WhYBh7
hwn+2bLkxktfgmXKxWsBLGz+MzylGIDcDT3WY93Pg91Di1nixhk0SjNXB/yPGUHs
Yexli40irj1eY9iz6FLl51l3pirDCIG5tiuHfZ+FGMuP0EBs6nIvgdBkdUL+R7W1
w7yjexkzO6zAUVR4kFFNGNqX26lxc0G4X0iIw6xrogxXoTiVzqP3VU/vtMwlleh5
UmAKbMgrU/otfXWCgnOjReL/MFni0GGh8Qyv6IAi5eZBSb2aSnqZf1CngqQmV8H2
vqR8ixZwQXX8I7S7OW6SIhe0Tfm0tRtOiZjiq39igKp22UFK3qolgyinugJcfJuI
0GkJBsIwrD/82NOwCxMqnUrljiUWbeNoNzhSpSg3gpJonPN+wMgPpOpTw1myCcCG
0XcKUD8mE3A6SsloeeiYS7tHsOa/l+ABU/nWMxhO7gE1SjkGL9GIDyb96wEAFefY
quLNXr3c4G7iB0BZdpsqxZJkBnMJxOfnGMWXiKU22iuVbNrWdxyBX151axZk/T7m
S7wQ+lgWXwzPaOvVAqMajFaXFXTJ21fB5nHoreV+JXbhcK1BCAHVxlhxXva89UpF
hlwr8f+evKbNvxbzI89kIq2T4KKsHQk7Ek87qw4f9uk9a98l9+XxX1/ZgNKcWzDh
Z5phqZ2hwTT4gPBFR42ULqwN+UdjnbXgltEFX5dZZx0sd7zN3lsDbWHPLEQ04s9G
thvLO47pbO+kWTS2TQC2U83Xodp30mEotXzYM3c46sYUtvbspIYNLO5ioR2ifuIW
gMfH+YG1GDi4e19VjHo9ypI46WogxS0F8EtOhvOG13YVVvvlw87AZFuVirQkTket
hsD9iDw25sDBLbRxyb97Yl78+IbDcVja+yPYqZtx9qCJ5+DvUhXXF6bjCNsIf98g
FWczAekSHA8oGV8hPvK0YBqqNusTitC9UyDH4F5McCjA/JS5E+TDYaH+TgSMSVp7
C7v36ivQ1yVob2g/N3X9sEb01pvY0MEy9D+ALEibgB/Hf+yZKV6XT1YMyvfA+XyO
IhfR7n+H4IhLzzEb/HRVOw+O48OaVkIgdAUDtdBoA6kZ/MjPYHM1QWWDwe2BxS1P
1wtm35bIM7h14D0B0s7O0/SMQ/A7sSU6w3nnIraOIeevbc2O8PGAIscE1tk3L3f0
Q5go+udzrvM2m507fKro2xtA8UVWbfCsUqX4ZqtMplX7bPv4WnZmPYqqKWCCPbO0
Sdb6oyiAFVbcY0ZH0aHz4VMfqUV2ycsHpctNsI0c3zHljtVPPa9kaSkVjVz4rB8f
s0S0wwF0N9MtlcjwW1WUSalREAQThkYAQ8hrCq/89hLmypc0jHXsJNOHjL1JMzbv
Z71YiBvmL7IYXAMEMOgtqmlEKyETS7IlzXTp5/fQcpTRDaGe94KaHihAvYB2oI+Y
PmQeqcTgIL5eNUGfKznHv41BWDJGYEYiVT8nkK4jbraQLH+1lKWdGf4UWwlA+vPp
Ii3Jw4XQBP/sN3TQSLK3pyqLSOGZueTdmaWMHbg4jMgjt2iqLSgiBbPaOjW9aGBq
IKZUDQ4AEHBRpS/HP7f9Y+q0Cpjl5EHztUWnxKuG3A1qxRg+G6AOEtva16qXNS6w
SKDYLVexFwc3BUD50eYVKtcraOCUXuKoLIEoRxXAUcbe7LlsXRhAhlWAuVXI0Pd3
SDlljX4GvGTlFyUVMg6Cw2+ql/yAOucntZRJa7gB/kNqCmCy6Qw/39JaL9gjNTt4
56OMbSB2wKCJokyNabt8KwkkfA7HtUgGVpXx8pHuXddDMDXztVqSB8nd0mSt+q3U
KXcODE7EKjtAJkQcbYAQPM8Ph1P7p64/WuPlrVwWC2jYn2xcHt8t3ENW/kNpCnwg
R9WbRQ+OBhLRpaCd9P0HehMFpAZmZv6fIMTPMTCON91wVGEE/cvIyrGnu04G1OUo
AjWIXPxGa6h+q13FpzUyH9UavPZaEb5UG1Llx4148utyWYWzKfAfGbCrBLF4KPuY
fBgNl5U2l/IpTrSjqbQaoyDQqWzGrpWSIg/ulopFL3q2K0ytrrKfjiXmlNxSnU7b
1ctcVg49V+UI15RfL2eZ5gWUtkqRl7432crGgRd767VkAPqOmeoNsZy5sQfrh+4z
Dt7a5LWyxTCtnO3vRErSriOBLWnhWZj9fG3Y8UaWv6mGj4Tn4peJG3muKLlgir91
72NvSAjF9HWANjEY2E5qnIK7RFuS8yKElb7iqOU7yq41nORxOSSJ3vP6CTyVblvv
VkuIzJzP1v6g41coAWCfvMHD5kpPTBSeB75F/Nz75zcqxjy7vCGA6/o2T5+WrtIG
BKX64ZzFRprSff5sJipM+4PuFaqjVYMrervDXC4MV9m/XE3M1EBmgyzZLZMUA8gl
yEJDNQ6e3Sh5wD+5gjdy2lZWYmdZiR3toUNfJmys/JgIP+djzVwgvcbdmqted4GK
b9oDXBSyqDJKfvyetlv6pGqGoVDM2OQ7j8E3ZeVtmKlRuQ/E8+X/ABhmGdSclbyE
lmb+x9/XIFQ7rLUDsDRnWxuD7q+0ExGez+kSE0Xlk5CqWJPum/mqmPtDgqfBsUIG
AGWcDfsnLBvsoBFzQExQOcTr8rJLZoNzm2p+1jwLpJLPJs6LqHlpizquKmK6/5xj
nQjDyE/2uogssID/xxuFmkt8R9wYtuu4NZECziVwChffWuxV7+0JAFXnGtIWs4Kg
Y2jDhpx0yt2AIabR6tv8qAya3WRaidcMHWuqWormFNEBsFWt9C6h+B8A8gkU1yJX
VmE3UgnuWQwUqljodki37eohehsIBUpYfQ5DuYyJL5lI6N6TwCxl9iyuipGTpq4v
ZjUaf/2m5GrYAlFKnwoOdCgInXLXOf0GaDk83YvcfsrvDg5U/sGg2v24d11V4cej
v1Er6Bs6UBKMBa0dmFksFs1EuRYAKwrMQ8M/W0imMz4Noi3YlkPUnBHunhzg1YHv
dpzVAfFQZCyPJsNkSZDsqd/gO+1Eke3yfSIT267Rl+qII4xZZ8vEB3MVWQCoPaCS
YeSiS2Wo9Nwy6bwoBUceIOkpfbGHpa7ioSUK4Ji10b2ZoeICVTrTKoz3oRzn01aA
PdNV3WPkZ08xfKlBSzYlLHGuKLDx9IzjQ8o2FnrXFSZuP/K9YVJOQKr4YuSLCLpT
nPSz0HeC1c8n0yRIi4bsvCtqvHnHU0Pakc23whUfoaVrrvVhkV93D/dQx3uSmPUN
r7jielchi6LQlMoRXAerpyxsmaHSEwuJuv46DBzgbXRE2jedvXNXio4RjQLEGlFW
bShz9TpNQ5hnuLeRRFjFPKBPYzqGWuGAnB623dGVTBT3qhWDQBDGazWu5Lwa0Nvy
3TlXSGXXa7MuHBuBrAdGrwfuBsUuO2TmQk4NzPkcG+6CCUp72Tow7GuIE0Aes3N/
lA/XtfjLr/4CsVraZgySbUHjeuQWs8+fE7kPy8hKg3CIWpd0CT6HclNH+5dNTKHh
yapsGcjGLL6bp/+CnLXomoxvpKu43FtrShLDmw4oKKLpmWAyJND6I4pPfWki4x+k
d4P2jy9PPNIqaY9HoTMjeczO7afz6omwYBpkzU4yri8nFbID2O1SNvT0nR5evnJA
hwZfdtKQzKYvu7z+rNwpGAokYoTdjuZYxx0EQWiGJ6VDUvwRGdCNbNi6bZW4DDin
fjd4XL2IpKAP7g8haoOMrb+4LECpMlzExBsNKH79nKlclMshtaSIEaOjdlHkiYD6
01tB5wDWPIBchadndeNUByt+4kIlZNoadZ4MUIdw2dVFEhlwTmdBF0A1L8Gx+RO1
ICfNcD/FRem4V0XD7DeTG7KBKQhE32H9KUz5F8mK8HRFGLlJAKwWpauQr+EtYN5+
xS4iebQFv5teGlDgPfNa/c9dWA3rHL/IBpeIBHv0daKDoJX3kbkS9yRNEszsQPuy
zp5eUgjGPO0hRWV8F9pQfy/5DXoIL4r/bsqnXiehTzS8ktk0NLqGJCG0OxpPut6K
BNRN0aVebGRNx5MbqOQnCAHV4EYQy22CyTAUm5VpsrQ5V0wpJx2VQiETB23Oq8dc
urv2N8iy1cBN42cnVQS5TZAngsd2oQ/NmjwGys4ypcvRkhT62JgLzvKR6kkwgDa7
CfV0o+T/jd6mKeHktenudI43ISqAsUxjvebksm91eDpLranYMefQGtkDXG/slKpm
serPMlXgyf8wJgUM6fcCxb4OlTTpOjeQWa2/T+R1uTLO1Ntpl+vRFu+fAvBBZqWg
VgVJS6iaZFzJn3cE0+D0Vg0N2Jb8Q24+If9H2a5gqF0ymv5eYXJQwAfy6rbjT2f6
YztDWevGQCqGaTi04quG2OUZmG45SCGUZEnCNNThuRLqT+Ze9EQF9RFv5WS0Vgmi
R5z4/WS+ueL3i1MRFh8zqti0i/g/hxDB+f6nL8s5iiz1xquXjzBR5XZ4OerjQeua
Yo3tROxWUhRA/P7LFclfsQCxzlZEZW4aRO5cQtq8/2+I+1MIJpnmRw5mPN588sH0
YZh/5P3ftOBNX4k0CE5A2XsNBb7QfsFhulJJeKCf4OJFa9HlZh6xp5dD2nEWw/1P
O/MvZLTCynIo0aNRFYy1a14W6yN+i6/nQgNloy1abpv3NHPWzJ2D5uO8KwpSAHT8
JVeLpQ9LMOwiA91KpI7GvuaMZraHhfwA+6pr7Tewks/mNBHrMo2NEpt/Tu02i6z1
QGEmgc0y0lngPnC8iJH2dAFmzMu+y9YtKjq+SX2sd1uV2kZMIH7fX42n4DitCQol
xSWzajQTzm5SlN/Wpz5hGaGc9eZY2O1ef9UAqIYUVMZX/CgsEIwjb4EMaBrEfZu3
T9pot0YHcs+HsXp5NawcQmCImO8gKcweZMzRzFvomeWZeKaOOBcVB09Ap/RKTCRD
L0W/R6DURY44f64AR10/C5G4wfzxoUGXnJTGj1aTR592KMkEmiZYEtuK9TKy8g62
G+JrCMS8nC6HZqIA57IwdpLPtfZg+or1f6XiSlLM/7QZFklPkhR8XREt466noLqe
KqFe/d7SW4FFtXqU+GwKuh/rICYwEaTarWh14mlAFYKESE/kaYQcsDnAnjlaReNy
J74ZXxEHPnOCo7yage7f0NRcDVB88qH3Zlq8EX8tpmTh6rNsprAEy6hN/r9T8D1h
81X1714ZVMU1b9bKnpkD6hFeYm0O4+hjeKWWTYHMvunYQ1mnCplA9gEqISaoZLTK
7eko4EMghHcu853+FK/NHUr6fuecvB1Frd+UcICQ/rqnu/HBP7Gt35mN+XFRczA4
5uvFTFwOThVpRRThy5NlyEqTw9HPTyQEp7t5wvkphwXdnmq4mfuYKsCAYKjOqjjm
b0FmCK7PY5Rfn2D7MBJ4/GQrIrdf0NgPEyToXa2DH2PHZaBzvRkkK4RvPhD7JT27
zqGcIQaQd3wevOBZ36ccWV1B7FEX5gUy8Y9Mtsf0P9eOkK21KeFimQC2BGriRWjZ
kFYRfXPXqebvzLnL3BzpNS3gfdD2M9eLuBmw4IciLTE3iYbiXl2MGiIPBEqhtfTZ
vfQFcKkic0NbBctLrK7BpJlS63OTkT5mGVaNHD8vz9g0XtQ7ZqL30HeSTx99lC4o
eUKOSfwNFAlm9pHDq1Orh90HvFKJYG/yqJP7R0Og9q+f6qGkmPAui+IH37p79Jv0
sMQNHzqPJIu0wVX+0K6gr9Kbhnkui/cX3paVbYS8WAOXBDsGTa4lqplxsc2DQdKq
xoYHCDvjf6j7WWG21l8jN3vhSsrcS5TU/nbU911+CXBfsUhvs256DWS0ab5jaQ7N
csH4SUIWGTNn47yRm1jMFYoA1tc5G3ubIC66aWzGMDbYrkrdvxxh839vQ+vN6TXN
Woa8eSr7WLukRSUJV3jzGWPlD8eA8tGA5+AHV3AJUrR8iYywwk3gTP7NIzIj48Vu
MOICqXY+uUBuJtmJUhUgQKfUmgHXVbpRYGjemABRr+zqJ+mG6q9zaIl/vdTnYMko
n5d4IpuB7B5W9xsBkDEBkDwi05QlWEztR2C3Fdm1a8nCXUplAM0NUCzUtuL0YMCR
GotcEBnl6Td6BcVwCWr0xCVI8ELtrNwvlCRx7r6Ybko20p7yMSltO5l/hIR+joAl
aJp8tYzLAd+mAnElmEVmemV12MOukyvxLLOWK+GBvjaxLfMpEFIqxJ5cXrNaO+Ef
PIOhS6+qgyHDI4ognTMuDi/LXZ52ki+EkffTQXYMteGqzd5fchHgy+S/zWBlRm7v
d5bK37AjVOVwcXTyQ3+fLxVoZljG7WosgThFPoLro8MdowoHxpgBGKTy06jgFjbg
iX4ZuyJVIZbXeaKEDdMXQNeXVimB4nsvjfK6AzhP3rvXdJAzeRgAQj5Rw5ALC5Tn
YI4H2h8iN8J44HlD77FMgySIKHi5cHxIAArmDIagiPF8ex6nZZ6lKDb5kp317UbO
r59FpRGaPA+ABB2kbVRf1u7itnULNnxHRpdlWgiMkJfWTscmRm30pLimxpD9HeE4
7XuvgqAi5JAR7f8cUf7Jdet3Pl4JrovVZeKbHNITfO22xXtBHwlLMx7EHJm3UuMA
ST/T8lVTFWfghP8OpCfrENOH0tI8Y6JGgu21IqmH6LMMByU6P7mAsBYiJ8WcHxev
Gu2xBWeSVCy2fv6kipCLFXluzQ2LW4GgTfftEA/hwNNkUmRmR3zHXdBCF/SfESeK
EH7wcPP66aAxkdSHofBfEgq2y0RjXbgMm/Mnz4cOU9qZz6Vd9EZXhaUiq1oPouPw
bgHs42kbwSsXUjbht7N0D0Fki/heg1Oife6Ywp+Q5SFdby3kVE1BlhXVMDoTPDr/
ZGq1IjF5mvxoGnvUftDCv0VGBVVyqLvvqQwc59h0UkiA+hinb+n7d3DI5269/KI4
BuqPi0bdogIfxSJXzUr8Z0m4zIoFtG7+eh9AfbgjxSnyTK6tkLYyuUmWVDt6R0gl
1BJiiLBJN1JFx6ayopJFsbSLOcDgTR5Mz3Yojl8GMAO1ZXWinzzhXOb7LJbCOf0R
tMvSqCS8LMFCgAAYMyit65S5xXyN5/o0lIZYHsGXHX46m3SQPIHkA1Uy8hawW8Dg
AJ0vv/ML5ed7PRFXq0ZEy0tyOCuyHYPPYA96oEOlICdtOa7mmy3HqX8Ls+o4JoXS
eScCJAGkR9Hex9WgF+IaZBBcdawQ3yu+X8j2FL1IsvGCes5MroTbg9NA5gl9WV4W
e9b5pzjqsue+z9AneD+Qb+oAvoYM+IKLkb+BYDQDnTlS2RcwL9qc8/R8cc1dP15d
RuArXnwiptwwypW+BQUxrTcBKUtUxjqc1zjCcvCfpIwy6StWgy7AeWxsG6wWAirM
Yzoau3NbALa+IjBaZlR49Va6CYhagFckw60wF/GDhZgdXSCfFxnPob3F6TUeEUfW
9fpdDUYNvGvCSFdIUKFDG/Rdo3ZYUaRGX/zO12P1ESO3QqLgtFJQ4AHiCTXR+7Wa
B5puBVfR3TSrC7jIhx8R0CJk3+ZdedytsTM9sUjgWB8B8Dy4Dq8PJkiRchs5nCer
iYpdJUUp5LzA1LtNOV1g8Arv3aBL+lgBEcJpM+kRGSGkXmGtD1MqjqxaLf7lkDzB
L+eJ9gbpvO3P97+GZQvM8SO7JXHtus1Se3Ww8Tx5vMCpZCagu+3GfdX/fAVNVrWP
QO883rjbdac7u6dSLOP7bvik1FZ8TevDcPESncGm5y31ettJ6Gzo9W1FZTO2lRkD
oMdvA5r7kfzPlRIYb+omQDUurtffJjn/y/s4he4/GrJw/ihZDnJt1MyEK8YX5J+Q
FOw/t3Sy/qiZyfkPnoBKQHaEQlZj+i8vmdOwpfbnRttwp++m0bJS17ENAUw0OOf7
JUl7djsCVKgs3mLrTcYRBxyWJ/pMKzFKejSLrZlDdaCUu+EO5kk1DJ99uVBERGxM
KIB55wB0OAf3pJ62jmtNc0zPq35twJ9xxkmGVJnJ/Bq4L6P/eVFlxor+Wn3KGznb
BL+jK9RMtrMcg6aOfa058zFd3upxicxP9iSVrq3Bl7r7MSQ0oD7DIzsEjNTrfMtK
HfjYk/uKAJAqDVmGsnKlv/hQj3wFftoHv01Nata+yBvMZ0TSAmSoVzZ0jJx+jmi/
01vRNqlzerT4bN9ypQxFg+pBi/3WAFsnHXN+IrZhwgAtNW1FWayOx5TZbZEvAjOh
fDvfWm05LaOPMvIvWQIZKHI2O/8HZG7WB/vyScroV+5kjdumn7c0Sn++pRQYhNds
gcQKacUulglsDRJjDZeX/9OFzJy/3VdCB982lcMlycNBWU17rxewU1femkpfM195
voJe6M3zT85wh6pSmfdMm1XYakDNuthchEB6tyPN675Bm5b1Ai1w3DqJdV3k/KoL
90uR1/PbndvujwEyGZ0VBf1Cu714uvkYbEi0eZteG0W5UofIqNMFgF6vcPF7CX6g
+sdOGo1aP1y1+F232a5tZ30XbcT8KOI0mf79arfy7VCAlQfx61hkc/EwW/XkXfC7
K3u3TFIQtSn0tTw2lfS52rXM+Qqry7xRgyHr94D6MyWYsNsSG9o9MRaurzvHjgHK
chLzeekJDpS2LoIgDFeJJswzMNuXZDUQDbKPTPNKSDZFk3r7Hb6TWMfPHkdxH18u
ob+uKG+E1+cHmUU9K6rpdMi/ktLlNQlM8mD1ghNO8KFoxdgWZpm2Uhfw6lrrCgpY
dbn5M8Gu6tS49DAP8YRXWSYqVZ5zJNPt9BD/FwEFBt0KUkLB3iKZD3IsajQG2cLw
d9CrhjKGqvBXXHdACepYxtNVmfBJYX6ACJWF9kcDHowVlxrO7Og46YuGRSD8tyhq
3mSkkVBQiatWAJ0HvJ2JdYXuYdjfGhlRteC94ie2VUzEZXBuayIpTUgq/KR6irdf
W6r7VEGMIeY+8rj/pwI4dYdQP2OZGGsf/1VMi42kh+s+LCWATWelkmWO3H0diFot
WsX9vtaUcBQ714GmmThnnzyBSZaIAQPPUjv6K7Q/e6wE9yb5/MIw2bCJX55A0mFA
dSWj0u167PpmJjfKffviKaYdNlFOeJI+mj7x5er6cJXrKFFSu/TB4EF1tryhWXZO
tMpcz2BSgZ5P0T/2jS+59W+OLS4a5k6lxeLPX6AmCjPC4mQ0pn41CfWdTht2wORX
JOkY/bVmjvqqWeDeSO2ZPNAyApN3g5fdI/v9c9QWelO9IobyylMc8vam2gRd7g5g
NMn1Xbo8QE2tU4YAYMdj4C5ienlAG/1E4YYsTxOFJrT1Ubfqfe0yJbvA6FSFxBfI
t3yLisVtFDxWnzCepeAuNlWr9fTae5FWYzGAKrssY5K/AHx0UnP8KWGcVkfqa+Wj
DfZCUt6gJMec08h1NvtiJeh8mOKgkr9qknaAwE3Ocmy2it/wunvOJ+ka+m2nPWO2
N3K8mDZ8zGvB3QX3peU7HMJRfrF6gw4IHgw+FGT4pH6hfng8cSEHGRnk3ZMqNM9s
KtyfZnGLcNHxJkQk0JgkO3gMynO1aCHVYUmnZPWD0koPSspuukXG3OKD9hVwLguq
GMBLHe2g2pXRTYTjkXzx358VcRssCmm1MYH7zk+XySQQjBtJ2DxTVD8GoSeXJ3jB
hSzcG8r8HtlMvkNLqq2av8VR/Xn0ukcIv0Sc3+6l3jY/ElLxB/aaYwXM0yQJLtfn
DiCPPIIvb5bH9UiaKkZ/YpMTpyaSzpzoCAD70Mi1bPgIQKBIIesin3TDqnof64jC
MwtwvuvBvu/2c7fo9vFk/Mf+YqxW4JtOXCvjK7EZmqZpsVkRBfuTbtzalUoRpelP
Oh0IinzmvmHnCyKeDSGyoikx7mBBwSGZTBQj2TK1r70imPwV/woR9ZpBu4a8ozW6
ZTLXCi9GwHB6gB3xQs11cJ47B+RfbdKHcGXMTBI7BJYRxH0ttBueEYYphJ79tXXa
C43DDhXNqAHqjsD16xcKU8aAdm4CkSWgeRLyfW5OdEijnD0RIx9QZaldiar1xuFZ
mdcnTCk4eN4nsbxgpngP/3cX6WpJPdL1QeVhQPuaVa4P7mc+f8pPx/KJPFLqIsiW
YQE5WgNo9jRwpkHuWFZDJNjMW48qzc5aXOszgYo0CKvVmS+5m+rtDXTQPStwf1e7
Mg7etWNRDZ0HCFjP3ExEYKEj6UHawygPh7xe9k2i/alDGr/oSnA8GieWM0JGa1rZ
CeJHgi8uMllb520w7CfVDL/9uE547JZtdl5Uwa/eeBxLN27/PU4sZRv8u04F8bFL
aFbMVXw/TsBE3AH5triZbK0mN7y/NkEkMOfFeGs3jKOPuHjzU1aUFjl9vbIsWm+P
8tKeM/SUEqqE4zEuSzMil15wQPm/kuordVmG4g8l9NpbevZ+WIh1Zer6084ciJTA
ZyYMadRaBSZ5D1N5BlmLiR8rL3duG1Fq1ZJEusXRBHk9e9g9ca8Y9hQe5rA8cfkW
jzKKY/q3P/ayeoDp4p+5j9xeGwTXgdNpt94BCSV97pdduM2O8usVpyU1yATdXIkx
TidXcn7pa9s8RLm0obMs+vsMEbH2N0l0ioXe3rYfSLA7sw/D9qfZFshcC25xfnYC
hcaleFUlLJWg0jEYruy3KAiLw6JH7fozN6diJ2gQvlnCYlp4QihB2jiinztglYJQ
ZEXJLyEWZyIGlqL9f8x3mqnoGBJf1BaqkZbFrp5h46XKrbeLBMtk7Plm5jWai6FY
fpzFWOJuQcTIKOGQ+boJoN3sPdclRenOyQJ/yJG15gt5UUk1TPFtTvTYVgw5XH4b
QRnv4T+8E9qH3vVaFbStspo/zqspOj3SVvMLoH1Z7Ll+g3VD/5TwevougD8DgSr8
XJ04UzLNIwFJO4B/zW2uCu1zywkDmkcohYEBR7PNGgLjRjqC/B9NZ2UQbxQPjdN1
GjyVZtz7nxtOmGLDPwIBuAjnUS0EobIV8oPP7Quv77WkHhisnTA/PihEfBZOvaQb
My/vXa/2rn0BoT0XEQ05PDof6/kCK3389/uPmO+1A28R1pftNMrxj2Y/UAnr+Dqr
rFt88tMiGcyWZIjWlZDIgWPSG/ltdK0oHRqIKb9b9+0olIYoxVlIs5L3Zr08uoLh
5QVUaO6V+Y9vcZyjQTjZLuZcVMad0/Nmh32uIUEwFveLIeczQsHyDSlJbW3S5dxl
C/2jUhIcyYA4pNsDV6Uhnu8SSDAeQBk50bCVNiparpE5RS4JUTJFueqTGTgo7nm8
FB7GVUdI1mz7d+2bWK9zru1lMrVqHgAbK40YRNQPb0M1XppacXHx+HwH0H4snKXT
Tg2RAUtIyLBPWwvTSy5erPI/ntJYeBy+0jSdk7F+W1PdND4e5Enm2zwZm/tVl23H
YyQd7nhGl6M5mubqRHoqvo5gOv/brqC0IlRQdsTaLqNi+15fzb3m4qBvwRcWKZTo
go5VI5p4ZRxmdytTh+ZMX9QfhJTgrVBK3odafzm4qLrVkd++S9XsZTVTM4qWNDHg
+QQFfp4tyByAZvTVxhBQtIIqtRilsxbhJ/zs8g18uumvKELJjJzK0VtQWTWiB1zq
trIyxuQL+jmWHKBVvkyvBXimJrEwNbW6ZWI44k+Wiq1d8ophldWVxnCtcqITHCFZ
jfW8dsiaEVmhQPYVVmX0GepacvsEtWC7mkogeuhTaebqtdOkxQKh0hxmXJYDU5/Y
1TYr5rZj6/KSJ1rgag3yw/jJoAFxIlDDi4lN029OjGaJoQu4W6jSDgxMtvbWubfP
WlhrTSnArXlb5inct5m0hGur/jvgS2Ab0dp0f+sAryLfyu3rBnB/+K5PMNo5A1DF
01FtwxOXiderc5AD4PzGWcguLFbm13G6eZ2fPQOTT5mFxvtU+K8vH27n7mi1bYJJ
xuhqu5cMDNodG7AkRRH5pIAiwUomQ9DMl7cmO7lazJe4PXBVstE56oEQa1Ac+xXC
A0zC2ZggPm3m+IgQl+Dp4w1wHMRcPW3z5JRJvLtFnk8T65Lx7ZwsGYouZndV+Sr8
es8jcXUwoM033OsPTmLuv8f5gr/wMH8xRe518r5l8W/exCTWteWli6CaMP1aNxw5
pQ8mcOsSuzieA/klBzStHERLYYwVxyqlFVe3fK5ViZmdZQEHoFJ8YzQyywKKn14Y
DErAg4AH+5OKg58i7GGDvIBlOrHlbWaAZXvYltcqA6+qPMIbeyvZvekpqiWdfrqH
CB7UimoHLFaE1QB+/6pQnICDSQOVAHU/JvMiZa+gvQRQB+Qe+4jfOUBLx1ExokP0
kf8e2sTRo6/B4JrsPtLGKUZRp+7/RBrv+4R9CyMJUwtjDdR0cERqRKJDUDpXexqs
FIaxRbW0pAaN48UU4B/9hYNMfccBUvfIER4rk+FAqurDH6ZTXGkLlfC1WEfx45jf
fIhfseHTqJjJExmyYp8aYMqrBl6QAGnd0JmUzzzqO2PD5Jv/k5xKGDtLhYiplReY
NbAAfT1mM/UiianEvEqxoxmhsDwcN0bHxwk5wXgMaaB7ayW9JjQNs6+fDpa1f69J
Coq/Mv2+zXUvtmK9VEKDlpG9P31848DyV4E7y15IExVfsUcaJjBtYAXV2EqTw7h0
UMVAbVtL6iWvBtN7iqJ5Gnp2HKm2L7kqh6xOuVN5CRvlX7DhWPDao42XTgXIhbZJ
jtiW6OxASfqBh+wG7+cRHYJScT831Agi0NItxOHybB9O2YaToU+1WDFTDB8kPROz
xtRFrkMqqIw6QjCL5MPx8Tu+OSvm2/yDW5GqQVTsahMJMaeOZTyfkyDNyrVw86NO
KgyXcmoPpecQYTK3liQcrv7nMU9bGh5QOtV2ZCiltMAlwxY/m9cJbSzF2lMY2pPa
XVNbYGBEHG8AJs0is6N0HYko3jROS8U269KcqgUFf6RDEkiuykyKkBZqYfvmmBAV
0FdQmONsDCIM4Ktr8L4meoSgwHWUwndZMM15m8WBv9tEJZYLu9wDut0VE80v97bF
0PhRVKb1BDkzPcAYhJWWUfPr/UzeQOmKPSW9L6GdPE8zzyHotvPHJp5C/75JPFWR
2njFZXeg/tppMO5oEpQXoAKG0tJRSJNO72LvcMr+f04Vpvp246dbeo5Jde9OYgEG
IsLsLGh6KTF72Jr4FoWScawhanB4DzgjTyJNZ9loLG5oq/rMgLCWLdmUtvg2DT8X
exJ+6TRoO4Nm1WYLfzpq2Q3oqysI2EGnAXDRYRyTp++UWxsbawTO9Jj/Jdz06bJu
8zQxBimEUw3ixN2RYsmzeGG1QQsVFZX2GWIwSxTA/SUSfLJzqnEanxtXZ2Zw+QZN
babA7eXiuVDwACDU3UxxdF0AVXjdUEds1zx2OOphRusW7mU2UvjFGyhZTgcLBD5r
xMT3JgSBykRfFZVedaZ6v9n86+/AwH1z0ebfrltt+MagTJcHLewJsRaSeiHMqqG1
gWUkn8Vc4RVHSNifdpqvewetlsDKoC2ZgdIG6pILMyYY7IRxpTyEzTKcknIUcU/A
4EgmRPWh7PLaC2CJQrOpgYSO5uhhX1Dp6ygw03XGK6vfWK+No8Dtp9SAIY5Eh5M5
YHlx05fFvSad+2sze/I9JKt9CbrHS87lYRzKvkd2KtS2wEPrYHriX16fUtFe8Q99
0luzui/1L8e+UlOMLDGteBlVHeUF6eedkmV7W8ubvRMH1FSrunfNKuS3+b3W3EmH
vnkMYtu9DK3QfOVDS2OYtOpaKY6mConW+mNu09flG+YUJfcnzn3t+6K52pg5U0l4
T77sBvfiKrUvZglgcSoTTTVAnOJB9ExA0L6HLBJR/iOckTEYGOEoFUAU2jtjteli
Ye0R9vQeZalJ8PZVnRombeuDdM75wsq7rh8gOzWk90h899NJlQeQ2q+/qXj/4sZA
aIhXGP1Sdu058uBaY/oSdXKbg06kJwzd8K/CiJzdZ6VKR7tanRM6WG9bFETWrmU0
IMLdkBvr495lBU1FSW7KD550QJOoNSyEGp/fXHHNwbrrpN8eL9Zsg6DAo1MkASw9
eJ5ibjTiaRP4aGdVtcCrN9FFI5Yx6W/18vD1VWRxzuZvvykmR2EAqdP6Hs7S+Zqm
r77DuXXR45KpvD7cY4oFKPfWXApK/NmpuQrpNMBJSfvnydDbQb7n2sP4tu/YHyNx
YzUUzl4fVBuSLDNZN0lebgjX/Z69bhTmTSxnK+Ks8hSmP5s7GUTJCcLBvexpnmhG
mIF2StTx8rjBEP3whD2EvZm4ZVDfeGC1V53h2ojLclo/BIa46lcXbJmm3wY/tZ5q
mcyeDPewoMOFORO5CmJNUyrYzJCn3AJiVTAeU7cm0JFQrR7ZzH1Dw9VHYSXdUCPr
jRC7nodU9bkKbV+7Zz9tWmJonmtK6wMGQY8U3ZuvVr+amCEUzZi+ltl5elPlPaj9
PEweuK4p2rb+DNx+84VQ1KoCMHGgRErom6RMF0lKrg6aPK6IYB2tSbrAMMrVr/C6
+vH67pKJXJZOqRnrham1iax3K/bk0TAuhv4Kwex9ieAx5q4qQh3eKMs6NRS2E3Ar
zD3gi+tYEcp7C3q/MLCC6WBIBJQRVMyUr+z9dvJ3M3vM06rbgFUhh1wG63t33aLy
ImmESeLj6jZyt2jX5ho/foml9ZBqSBANqsEnPLT1c0Jgg7WufK1bRj7zqEAnvlhc
gshivy2xqMxOtwVTnI/qkADba2siQdsy/jscQnDCU3bquehsXWcyH3065MjOYPiV
x6ykuiTkfhU4rAzz8xTcDhICJ5GRwffiNEj0TrsJoSTRtZs3vX3N0m83si+WCEEs
OlDbwDqno9/D8aAr0KeEzjr6E/YBAPQKvA/Fx14gYJ1Q6a1A/f1tOis631mBGF1S
A5LNW3KG0YAqSW3e2Qdb1Ea7GtO6nnVoohLvc7YxvC/QGtScOHYgx4c9BkozZBid
uhEE3drTM2mwRA82D4VGInvMMAJIKkJnUO4OPvh0qhW2gi5di4NuV9vTX37yCZiT
iInV03JzA5hEGPeJxxG+YrORii/JLbTkHhzO4DeK7dzaNLzeDMzpc9aDkR8Dclqc
qZBAXteAlabFhl8nbDL8IkKImJjU/3RcnLGML9w7Of/av1hpTjG+WMDVL+Bl7W2K
fmsd59f+8WdbYu1gRACdQgTroawFf+cuv8thQHQe84tXjdl2MGnewHmXJr8+2h4Q
FbXVYqXce5F74RZvMv7advYLFtwAbX5/yr/8J6vjtVVGQIbMT9fBzh/jZjZHwyY3
s8eif8ialoXaP0MKi7tokNwCefPDEXvwezpMHMXeNLScsaM6pNgK6NOihXPBxq4E
yWJ5L0FztDrFpvJo8TCKSpCtlK5nOwUC+y6SnDZQQq7PTHDFeSjqIg3dawy1PPlg
vvEDUVGYUrvZ0YddzU1jnBsy09ga1KxWtUVkTMb/bci419cD1Nu0ODk2VExJMRE2
uQOZj6jYCB00hLKrJc+gLCoLG4lGtZmpTDNt51tI00IyU3rscgA92ckJ3nC3oKXz
Nffp2D7BHVrkJhG6iBWLT+lqVvh/AEpBs0VZcmJ3+9hQ6PuppzcNdvxvYbX5WD0i
mIiwyHYvwTSego8/yveTFHcmsPWlGpxFzNFCTrKXn2Xo0bs0GVJD1bh7istYbtbV
2ICp9bG/RcYB3x9tIPHwbb9lk0nIq9F+mYEGllHrxVv+PhRUGArhn+cugBtp9vrZ
lJ2lQLnDJt1La5KGF65KB+PDooRzk06xrSDVfNRu2sV591n/uY30XFlNq73XxZWZ
GrYh8sol0MAmumIrv4lkle5r0z/mFIrTcjB1Dbn2SiL9kuSf5PLi1QQM/j7LaMz5
xqA2t4+90pdNDp21XSmOE83y1/b1AhuRikBD5bz7n5bXcv0cfsejJSAfPKW2hUHM
mB23ZK0s3YESyr3glIx89Dt9Ts67bfIUDgIsYjVMfPYEAqOSGfpw3VMKU+WDWYsE
36XatwLNOO1aUfbCj7xfApTHzxYIy6DGgZXDr1G1Sjh9QJA9AWB9KWgyHFLJUeH0
od9e2vzsdHfMF7h3XZyoD2tqDFF6EPcyah1vjykI+3jFpx/qjRaXu2A2jpXNE56a
lDbDCqHAkNdxy69j1tB/etV6IkpdGFTJwFe2fZgUKeiJz5McOu9AJvcTxTxwgF0W
fo7dXafg60pKsv4jJUQSOxAUPiJ39wrLi9S7UiVMMB69AwaecXz4UjPGWT/2G5S2
EqZg8mF5qmVZygRq9jBqJEiPi+lKKytKtwu7XHNwRcSphrsZmoI7ay50lmc05Y0R
fvCYf0UvNy5yiJY66BbcFH44V8E7pvuSBceUjg2GBxtcXSK4Z17Pyk0I+PfXhAsL
mltBbg6kDJTJ/9he+F71nfjX9MVLtlEDT1gd7F58FWsyuH7D4UNtWHTWx8MWS92X
lRxHG6CMe356Y5slbVUJNNCbbdsoqeh5shQIQgCb+HTOi0B0rkQqFUroRMjaYK/r
JNFHH26DCuiE76NnSFCm+Vmby+QFy7w4EFU5plfDj/SZIgeOT0xN0VlhjZKaPQp+
533El8hw1c6OXgSRZjkscvV2Z2XfERUQHj+4uAKOYsoZm3Nr3RwHUJr0YN7T22o3
MfOJiTwzJ3h+x/dDiahvAkJmvqt0fK5XnT2xRxf0agt1Rn443DOIkb//6qSXgB6D
WMFafMm/YwWLUw6Zwp8hpSVvSfrAOyC52Ojcg41kwa0Jd+6Hy1TyUr/3hcur8cbC
jx0Kj4CbECGYMMo3g8KO6ttDmXhTuFjfycVL0PfZZDVd7kKrCgnq+THD4u0rgVTU
ZKVR9D6bZLYr+aSGFcbfNcS9Sl377yvelXwTBFJpKZQq4hwv9DKcJTppCf2l2TYJ
PKFWEAQtYDNLFzJcMorogDrMPQvGMyvSTWH64707G7iSxbs+VFHC3fIim9e8VS3l
/sTl6qVXX0gq+2OYJoo4CYBM+O2vwJWCmELJmB5UTYXovzlcTWOiLCdcjbIaho99
W4HKrhDDHlQCJ4YLSkUxX1YdyZJqS/CgM30uJRjT6ezrO3WWRmon48pRo3RtTh+J
EMPnXfahLYQhErqk35J6VdxRVxvgv/eZunvNQ8Kzpy1CrHqvQtRiEW/OpqkFq7IZ
VxBdMmW0Co6stV9tRpPZRwoK/qGZLtQkEQNUXnz5n9djhRyvZwPx8XFexec+SA4y
hdRS717Nn1W16JzmAnYBq+WTNV60udqDJ4GA7Xbc/mBC7tAigw04l+B8ON2lrqlw
ZlWlaQ4AQwqMvxhQZ83RwOnYpBMOfYvDfMqze3ZT5z/8VWWk5YPBMpCI7rfNdfKK
XnQ5SFw81niV2si9RlLtcLutrZxAdXTZBkvLRyTHpgFyk9ohA91V4b98MLtT3a+k
S5JE8CidfOVv8ApJd3E8gZ/wDud/laufuPKkaOe3filFpbzUN60Qe90N3Pck1Lsy
roZbbxMrDMpW3R1vc94qJlr9UPv0/XI0ubsJvP0DldfZ17u0fDgSUkciWpRCrY11
PrHry4zRRnZTu5soPQsqWJU7v93l4Pb+evSvJ46z+bdCP4HpeWrYG7VNqCMMsHen
O9WqivB0uIGa6yiJ6MUUwFzzjxfERp4lk2Vm/HineAp45HWOJZMrflZB7siQ+Ri+
bNfCOK1/u1ZkKYNg51eTL77BUNdOOdjqFwKEj/5xQgnjmY+mG/ZaRVBu+Yd4vlzq
sOB675CjjtRkHaaqHTEMVSd+q+dHE724GeGlTu3nyx0Nfra6HR6ZmgwZgUdb+fA8
dyWPKNmCmTJlW/PUZ+ZH2dPjqtcZ0fxVPnGqDv4RpfeAwAVUjAnrjga6vFUt9QLg
/60yevOUyvcxQ60xM1qbU+MNICo6W28BTyF0fYb9lDPY/97Zp6tSDppI5+n/R/zo
GqOeUen5nM0eN2v1LF+vTVSNQzFphLBFvxn7/cTatAh6N3l89TsZhutYNmLKHtRn
fAN9UgwxPUp+PseZt31IBMhje7wjTSLZ3b5gqYllsZKy3RZ6XtQYkSm97Jb/i71l
KXQiEpErFlKwz1JLVDCnq3vNR3o9pzIJtZQ5D16KJLvCsF1uU4L5lcx8MKpnNvOm
Cq2sEoSjh3+svCvlSoOorEZw65YKHOmvCHjsHlD04t7lMVcllqG/wNj16TCbAS1b
kvfIQdE40nYh7Y3KT2v8ObK4mGn96WMC9s0nJhvZOKjpQwr/hjJx3R5Sq1nl9cKB
JbZVmRhIsEKk4I/+gN6Az6dkZhURTQqT5KJFR2vFlcPsE3yXJscW6oJuiPS5LaXv
XZkLd43AKHb//wgmAz8THendsZFjVRwo3Z6uhMy132ayYFQz4IsqfGhlNMGAuSs1
IqUFo/+iMl2+vVpN/eii2Q75CcGAmxJ+kqQX3Y56dSVLTe14AMSn1AT0n2xOZQI8
kOtl+XRvUPVkTFrBEmYrv64pdbLOKuJMrT18FOfmd+5EyR2+vxsrHRicoLuVZ+DG
cfDtPcAozVO9t2IJBvwslgxcm9Xujk0KUN8Ty6+OX38Viclb2WzQoiN8OK+THlfE
2IgTZYlZ0egtumx0DOtppK09Teg660Yz2Jvx9ralAk2E+VK9qM6AfPKLkPQFcODz
B5P89OX/urHe0YhfeIGVujEnjZDwYdcP9lvdYTQpf+QOR2EzK6pt0t9hsuiqhtwu
RlKsab9H1gxY7tz+mBnxp14axyShmtXthK2hTEETLsCfQf+5zopa8jP04VCdQnL+
haJZRh5u19SPPfhBygIFWCioVXDZIokWVpXRU19X6zCockiCgYfAZ5EKX2r/6h6U
g6ZsQre/NzZl3kyG82Hg4NnAh3Ae1C+CxdLUWM+VNAhc1EQLBeXErKnOnSFSnoqb
taQzuxi80d/nG5Ase5sbPliJ9DiYfUzBIg0oUsPcZ3d8PPjtN6s+CbmxSdm9Mj3p
WbyaPQB3GCAwWYDm7t7FBbddRtk0z1GNpZDis9XrJL5Npm/KfRFslSxv2iykx+sk
iCvpt/Fx/8yB9U4SOUvWtF0E0j8BmySQKTyGBaP1qao6ltnyESCvDPMegfO2koHx
s2QcyFX7v+o6UB2Hxdczq93tJ29o2ekDaUzv2sgKrg5CU/QEgSEKhLAx90bk4/O7
lV3wI2vFNpyOYa3YPS95YIMzp7gdr8byGaaOa9wy6ez3O00Wq+cC/AHbJPKV0mRB
OJ4nIw8IZYjBHYvaRB0bwUzSfbQg2HNPl2ia2/ylvuVjGYX/S+NW9wgc8nmeDjvw
3S14UtSZXZSC1E6QEEO2NVuhe3DJZnzgyHR4yKEXR68BZbdTn4x10huo9AEsesrV
5qHNrPbiDq2iRB/Q8xm3uwgWPuu++6qIyv2YDYna6D/HlbpHNNFVJsNJHiCmH/PH
I2hmKy5NW+P8ciIirjrsdz4v7F30PZr3lXVKh/dNdPH3+RzYAxg3+l4XIH9MBm4B
eyGJnabXjADkvZD+IjjZ+VLBo9ulEyFxvrgV451VePn9t/PmU7TrDW7n25Cey5az
3VSSMl6h/COZeZ8qanImXB2jLn7Pak4qcGmOpdVwdzKY8o/MrM6tzBKidJxmvGwn
QHeDbVqp+x8wltV8ULs9oQoZFqtCjB13zuGSYLOqmsgjNY2mr5br3vPi5ogcc+Df
BSBmCmBLKSBIhOTyt5MYvyWEHOOGwArjMQeW6oWyeamAVQWr2u/BYT3Vc1seLl1z
Lh8lfISBgiEO/ueJ30LBpEvWJuR9AKpSkq01Yxj3aTgy1SlvnHK9kw4xsxIqMrHH
eRRoLGABy3BScPN+QYQC3mth8MSnYp3WGXiSO3cotq5/UhjB7kMzqz18ZuUdJaGD
Xc59OrzU9T2alrOPsE1/Kt1j/noQ6rV1e4tGGyE63CK28dR6vsrGnxHzgNqbE5dG
qotVEG2cGf4PXgmKOD6Ey7cluNxVh2KyakGmd1x1GpJnwfOf7l4GdjL/mCrzuIt7
2A6wf7f0aF/um1q+XVAxDeHyZ2/p32egOMFmF4Gcg6gGpr7KdkaDFSMzore+ATVU
UYlY0v3tYkRjCrlHQ00pjNpiJzg5YW10YQMyaJ4vpD7jQ/K5nBJE4u7cH1/jGhbw
cpBSKEbqrgDWkjcNmgnSXCU+t7CwEENBbKXOgREdI2SrgAp7F1+pV8Tuiu1U3z+U
5DsDeZAUElJXh27ipw103ZiHVxCE6jvJiA23A17UanmymM1QhF+5y0zlydlzKQ3v
K/MBYMv7Svp9DmCVytJ3bYBqlpatsS997sNBZmqa5o9NBzp6uL9p9eDpH27wrW0X
tdNxnFwV8hiXtvwaw3DDdaTwcvAsWIm1cIpPWwDaG1iDEdxH9nN85Vz3I1DwT+ji
FdUgnz2q2ZKlR5ffnJJhtXrOAXmuOFPoNSFa/6sSOokRa22iHhErikev0RduS4m6
TQLIV6WR0C53novc5KMbILLbHdWjmS8pA/T62z3XKJmIUEabe0Y4lIOTo0E57pHZ
UzZOEdMSOCivj4/dwfCPPmAL3azfZvQbXQtyCtUlHYZqkre/H9UD/UMExy7VXaX2
yTyl27Pzg+9Kz7QkOviVsQ6e+POFi8mRtsT8ARBMW0vsRTWhfoBlSmfqfM8G6Kww
58ySEtOwmt0aPyDj6j7GLPQM72VuL+BPYMJVfVTTO1cdNVAnGOTiHodHRkUM2reV
EZpxMIezps7r9Z1yRQ7xPfj4oJl8S+T9If0XcCh02g7UPG3ajKIkncssZTfP9nuQ
q+P1xuqadhfR0RmplBcvp5wUO2rjcLMG7uT3Am+diHctc04U2/n/xkGg9aZEwbwM
XYLVAvCTEIGryOEexT1P50t4jnMusoORiAsPmgy/Sa3L/a9w4kOaN7F8d1nA1VBk
UnfleCGXbg3bDY9gl+qPbeA3A/fMptzjpgjtVSh5TBrgY/8GvnwjD1tuz928Wpdb
+ThyoTfUKAUc+Ty3w32yX6XhfhNiivlJXoUzjc/DYa0DQH7tEST1pszlmE9hXOJ/
a/muWq8F1yOGmFltTRPPa7dZHcQvsjIkJ4wj/xsLqtuUYsDn7VwEP0vkJUxt6JjZ
RGKX0GuuKZXzN9GFX4mX0J0DdlflvFANIehB/5pnmD8NqO8EUEDzIbrD2x48OaLx
bYQMH4CjsUb4b3rEhX2+R/A+n9tx1vBChCYotOstAtzj/HJa41Ues55QZj/vTRGt
5O/YnJlxZxhVtf+hFYQ3VdWgwZQDBvHXYU83vq8SsLoT2BHuyIzx5rVpwTmx10QA
jebLZ8knrzDb1CM8QjbCSfCzIMCF4rXERGOwdc5zGjUEfKa+nIBq69bbRzRG9UUT
pyZjjcs7pJEpLF7BS3XRrhyrg/rfBgLJqbP3f0PKEP4tlKRE5B18h+btmoQn5yyz
j15XH1GkvsQlrPNB9wqHcZN4r4zg+iKYPHbFH0zHRSwfEIYeDjjNG2op8yN+kell
+tQkQavY35K5WJWAvEB4M8pb53f+MsxqnXz29u3+E+mcCczAvX6Db1IQ4HkcKV5M
Krhmg2QPi40LWfSeH+d+3NXXDQ8TvMdx2UKA6aJkhZtgtEwbEriG87+ApFD5IWKS
+bAwTMvkfdOjV9MWi9Qg+rp5xKjTor+qplbuOHtW7W0y55PdkKNo3CYn7EcBl7g8
5Vjngb6SfwNvlJ9Ac5NTtuQPqV0aHWMSmRDdxo0nQsxoMrXjhLuS6eoEa04FFO+n
qjdBpBGbhBHgdSDvViTBKYRbuKEcJSYJpAWvYJg/Rvce/u4Rvm3CvYn1IYV4YBUs
pKcam+siN9RemDyg/nLHPczAC2JlkQY24vRciVa4s3/xvV9nqZCuBLzuekU2a7v4
rf3+2N7ePolgvDEpOW7vHGn/aslGvZzrkVQuLK/ruQB6+9Dvt+6QszEaIHhpq7Eo
5PGG5gvKrjTsUmhHZR6KHc4tdwwLAVlFrxkXLCKcmDswQVh28Os48ulfgn0J8JfH
NdEMIefNHfxVbdBtm86SDuBt0OoYBsxQXYpc2Jd70NZ+mmITbM/QEXPbmNdZVITq
jQd1lm8CbtZldvwUT9ikBbfbmgbgcOqd8VvYFxrGJun5j6L4PZ8cpqElMVfv98sC
iq2WzibgogP/HFyevtHlDT6C1mIZnqKQI7Q2lxorDGuNZfuMXAsX1H7KDq4mHfem
2nQcCK0Wekjs5bx29gqWjcQhOhYac0hJzlwVEWiXUTBsNgO/ybtNVJiZ8yp1irga
5WvX4tMvl5xMRsP8Tl4XCrqfwt9hBR16Mcaj41SotKU1F54wGyVG/0Vd+P8VPhnd
WG6eT6mnz89PtoceJvSY3L9LXy33LuWLhg1u48iGu1Ar/6kLaQ9ngLbBOXrftTu8
aTY9c20adnrEqj5IqwQJeW58XfwvDTbGfkCp7q0PS6NiuGPk1Fw1LlKrD0ZOZnsZ
WuqS55O/reN2bUziJLt8Sk4moOqv3R6YJX6Iu5gRaNkNMTkgmKsFUnUqA7YwCwL7
lb7ObnGhwX9MQXPfmzNauJrmLy7lLFIGdLaSTUjZziXr5E5ArZbllzYKz5JW3YKR
pHbQdGdLTZH9ZUbnuXf07+VZoSuPyuPNik43gTyM1HeRTey19XiJOgyhWOLXpNhd
hbAbOrWkgmo++J2aSXB54sHPxzqqYzGHERBhdRJ8tFmbjrF9EsNIVjlnhTqmEVA+
gYWlo/ihLKub16UyVNMDq/3nvvjv2qJw8N6az5zvYxp++V8d64gvnGFi7/ocpC49
MjDTapceQhPkGreBI5xWonFxXiSs+JLQ25n+1RRPI3dnQnrj6O2yQVIV0C2ezlfy
awuI9RkPwu3YXIiP5vQLBRqra0562xiozLvEFRaZSLCnBVYjaVJRLz0BAZ6/xYhm
KzfrkKnVNTiUv4b5o9YlxpFu8XHg6rZz0TSfreczq39ku3XHJNaY5YSf8wsd83Dr
hJlBLOvvb+SuX3w7LUYKIzJun5f5QsjJ9tL64Wi8LYEfl4zOn6w77WiXl/TKtfsy
z9d/AE1uN0PGEm3/6VMSiRFrYPzJO3TecNcXLntb7eV91D7i19PMdGb4YIWYZkqx
/kyS9mZan+vStlRngLbgbODR69jcCyEY1ewbYHj7oBqUR/OS/v6qxhmFBlArjxWe
u5KBIbSqHTlu3Fp88YYX72pYWb3Bmo2bU5k5f7fUyU1iiKqunmabGgp3gXA5RoAi
JwMJMcWWljbc/Fm7dw1uf+6UauAbLe85zskm7nAKinF1lI7SWdqpiqbhn/4YFnG0
1+5wP97DJ3UTvkr+4hxHlqRWCCFwxZqLvSzNYNDRv2fNBMD/6AGxfHAbj9Gy7hnI
wxLS2frvDQ9yxJykse9rHsq2vMPnmhfdqS0kJhgIPzWuNwDrBbIc6Y0ZdGnKSCBQ
qUVmBPJjLZSGLYTuUREL0YoTlNDBCYkhM4EeuFjpeyyVa4KTRuRejif+U8RvkRYt
O1vVjb+mdazSxMEtp+FDcBXZjj/z2ZRuE4cz4l/OtQA8UqbmHuojocs8IwnsoSm2
MonPQUdwvQA10AnZgLuYV0CKUPAJBpn+JzxEf2imeOynfTM+u71j1iLNuGcY1Q7Y
R1LVEL9P1rSWgQTP0OxlJbH/Hp4qUm4BICDTklCls3ys9aNZodAJ+3tKcoljCoDK
8TkuwCOkQ+DwhbZ9WkR4y8Jl1jnFMH/M3wQePrNoNXZGSkF1BMXjQhvUY22veNf8
eqvptKFMfdFIO1EABoLf2nUNzVqAoXjrZiFdjl/k3TbHDiSgRxbIv9wxELZU5AzG
UXUb3ln2dJkhwyxgeVxmoR3ijlikoa1cn/queTQ1hjnWcObUKclRHPlCxg32SjQP
87+LVjpwCfQWkNMDhQ/2q7FdtyGkiyEsKaxrv4Rx9RwwUPx2/924YH2s9iWw+0ej
MxXmao2BZPd3YmOj3CP1OlFxJ2fZEUfiYjFueYaEDfvSq/2wpYEVM4IcQlvo+xpo
znc+JvoVTLloORIzZdJxW2ACPq6MPMoV2qzRZXdaSHNkUNXLKKql41+FRhp60CFc
1hyw7b3qE61OvazmNJxAFTqd4Gp5KmwyvYDoT9GVs/2rFAKLYW08RK7byuKseOxo
X7YksHMadM3MCfA6JZXlqZSQj6ZpxwW73tywjxE9x9b3FP6uPGMFWFOV8h8O4o7C
IueNR/h+drT3b0JpAzYuogtg0WlF2NTdAu7kIABMkrrb/jCKOW3xaWzpZV5yd9ah
NrLQ4RRhwPMZ7EJCGxFqZk2R5FlbPpPFgiAZ6/73vRcuk1q/3hp+PEjE1bqTpGRT
jKDKXIfG1lqHzgmwqApXugTV7wCioCghba75xIY8bkX+MYfAAB2n5JYbmUITx1gQ
LzHWtUm+L8PabOqZFbEvIl++3hj5BbsKI47Txl6ysCUWWQS+vL0ovKCJ9SDUko4f
sonyWZp53iTy0hvsxpUuPpBRxhAke+CdrIQkoGzdTnZM9DITCKUekUgxUZwr1ojX
G6PxiMYXAxH5du0EmPcG3SxJqasO//s6+WN2rTsd4SCwptQq74Ie7MeQzHHg6KPY
i8V1i/58vsezAUjDtaWXe/rEHLzIzN3YCKpAgmyMzaPY1Va8aA+RK+J5xWLWTwDH
mFS35KT0bg6/m+q0TPK7NXHcyo9TDc3GMM+xA6aBu3qBdKz+U2TZKwpfZRKF2tJ6
CVFOT9OKbcMNBXNFwQVaszt7tApRFBNG5qI3c8cI39XkbleNtnLskog7QBoHjQHM
viPy5CebEOtdcTIkJWZGgbebvZ+7Fv8/9CRp8ExBsUVTAntBaZohXL0zzjjaf43b
3XoPJk0aJ8oYdkJKHQNm8n1soRRhUeRBUrmyhetTtvnfoDA62cxQmWD/R92wqOFo
FyJJMT5vAxvU513pbJSF4FxkpetUTpoT8GZUyQnVThIeUz2Hn/InlujOxFoazzA9
/CC4g0uhYSM9yrZz4Eqt+nKVja2dhr3vs+NBAyrZTvhpzYoCe7rWkH102bFGPnic
czHKFwdQBmgcW+xyDMktx3zl++/yj++XaD7IUjebI2WpPfUklTuospuvSAeMhRKV
+t0ATVv/m7wEkrqlf6tWnbQE2wuTOqmXq5V8ck+p7LaSnlTmD2gbhyrz1wOkB5sD
yP2ddNLqLWNUd+AqH0DoSdaFCqhj1fb4Z0eTTCYNzZaEgyUbVXeBCAOEAAg/dfap
q0LodYmUWahNJfepOBSA4WftLJzmWCADFmrI7Kk9gLX5JxbVf6ZWMi4Ke1XQA1dA
srlZNxuNo7LaWee6T8ZZUrE26Hbq+00jKlbNlmZaVeJ2gaMSl1d9hvCmzHaq/TAh
Eqh+ZVJDECEK/uQi05HHkPoACwR4XJhG20Xmspv6XXQs91u9jEBnhYYyQrWMSgw4
RK/i+POv8whXm1zUTflSD12Q7t1ChNT97D8VP7QR4lZb258AWpmipW+SNB1PNQwg
/PWH4JcbjQHQYrnO7q0Wjhv2mr/xpJcSOD9yjkCuAhk/99Ie6IDgj7LqSqv/06QC
hJkpxOifJf5GuL+43xPdHPN1ysi8/n42TS3rOOECSEDxpUCiUoLVSCyZWPjLZ93X
Whu+uInQbemjcQa+025uBnwZF3gykz7BQx1Vy8dMsD+e4VSfFKeIm5pgwiBtd6JX
ggWMzyctOky3JTXveK+BGP27B/1qZCcT2Iix6//A3ndAf2IHBFzKdrOIIof/M8M5
NM5VkG5cpl6SEFFs68HLHuQnE3aouggKigTAd8tHaTSKKxCsOFhK/Hznfk1/hkNu
zV98wfslxywOhU+DcreqKYV3PH8YxtBatg8f1LG4Gi7GOoXvAtBaVrHX4+CNrDBR
f09APIXHICnwtOAxq6v797NTzbBkVoqNXjEBdHO7aSRRDIbRh9gf39s7PgQIdHrc
2uv4dF700pl1qxrO3FnTwyZS/cxGyj4lx2Wv9P7hqZbiL+YXtBNWtvF43C7wcBF+
rQg8jXM931ONAhMnGhaCjitAOCS+x/0zeaax6HjcjcmSIkUiVzpaF0QrPn5HRRo2
c49qHJWyuAqfQRv/uHkMjVzl2EfkzQ+0Hf34dpg50n/AITnhtqm1htynkeD0O4Jp
jzNUvewTHm2M97iZRf2OpVwIF3hXY3yOq8NE4TXBh1AwrTsO91FteGdt8wQf4Kax
r5S0Psy0h7KmmY/4DpQhBsFDWRv42PDitr+ya4VCcimW6Ltf084xgcSvdn31ZufC
vSUM7+UnNTsgO8zXcjxdNQSLM69D2JFIBXxvEmwPIlJSJEzGDXcmHp+ofEiFRcvJ
IOGfwEOXK9a2yxjt8CgZXk26HNHcRwZTSnJh75bE6MaueK56/AjE3XO87i9tKJAw
kgsGsM8WMkKXuIcM2kzSJQnb8eKYz7gIa+THJnf/4TmbIQQcBgyaqg5IcMnWp2Yh
MrWe5cYHqhhzgkSbcSSvjM88upQwhGesI3Wxrq9XxjY74Guvprn8GeEo8desAIJj
Mz7cWquUplOMrs68+1IorLpTi9u3/UcyLWrZ0CQCnzbgrP7B3E5CRvvCtfW2NZnS
i7CluKt+S1tXT7mBOIVGHUtL8B7BR05PTV48ZSR0y9TJio1jdOYAmPOh/PaHBjan
TxQkT9yv5BKhYV1F1rnBMPF7gKSjTb5rvAuuidBJbfinJPWiXWB0edd/g6hapT7M
RS1GKNEndAmn8LYLANDKPWPadwviPXoenqq2uyzV5u3ChJpAHLd7RYCPK5DQbA4i
+vKIBi6gbUpknTU8kcovvwatT7XNlbAzB2VA80DPT9YLTJ30tjz5yxpmdLZaUkKk
cHTgHOY/t1R62mN1CWcpawPgCZoy+AU/mPa8QneFz1CiP5FMjNp+ZefGAXMhAmpM
aEVvmDaBMCRF8jUcQWleVhxBvREiHZeJMbk77ig0lc1YcGBC7R4jUl4Ody/9cAWM
AJ+Pn2FPvipJwTd3MGCciDuLvDJ58brxptZ2FpAeB7uKkfkPtOTRu6lXU2HXOoKQ
UMy2jqvwPo22ILSafc0Dn8BUUC305n3szhofX+MQbD2zs0QowFd4lZmM+JhC1VVr
5zKDGWQ4o9YGU1YS3DezyEj9Kil9ZjJZCg8ZQjS5nBoteQw9eu4fXoihh6BAyVpK
1v23DziR0rgHQYuJRIBPePrfvhawhyOXUw0y0XCbtcgraA95QIwhCihGYLKBy3Z9
zFBXFNKylBczJq1N5jid31LDHmbt0IrRNK4+Wa6IL0R8uehZ/8vRawHgxT6bj7iZ
xTnDlCSeiMnZrBZB5Z74c4fzaY03TaXc6M6+ZbibCFLkR+eGwJK+fYzrRf33ZCH2
ZcadRg1QX0eHlivfls+Q3nNI7hHiFP7florWTXWPfNlJaHmcJEfH0/sKGWTHb3iD
JdFnnWtPt99ghylJRfXKBAozbiemPLXjZhFGN50UZyOtexSloCBbtHi5TZJuD/0G
u6KL1OZ9/vSSbtgckGojcJ2nTLzsIp//GXBwVGweMvzDPLw44xw5WtoPaeRBh0QC
/78ZLvREx6tjL+Chtj56Uy+1Hzw4SN7bWS5O2SC0qQQy2yzQLKqKOofw5eaDvzRM
f8xcgVauqLjK/xGvmm/5/WH6H7GYt3EVjH7NNTo55wMcrfR3ydlCp43T3eOU9lDS
sXmBod4/i352A7/Xzqh7h/fCtOoExlX8+Tau+EbiNTkaEQ3fahrxGC6EnYZkpaXP
23T2rKWZojtxLofRKlcQy/LBIiuZ+E7eYJCdB2geiGk8El2IiR2p4GwSX8TZvkxb
qYhzTvx1OYvoMk63u8yLYYb3fb4ifp2rW1z4Ag0i9K3q3iKOTjWzL/nPHWtO+KRw
CqHOXD0M3hj0eNtWz4hucxnb40UCF4sHt8BzOqwx/oZm/p46HTecFkOJ8JwQ1axy
hCVfygYFQUVTbiW5A/2QVlEl3O2xmipDF91BrlNE8nC1fGiRiia302s2Ktr0+3Rm
OqgqCOJ0k4Eep5cOfGQikpTLyu2iZz2QfQyWgQ53amC53MfqMVhCBpt6UGd1hxuk
c2qfFApt1lO1trurqr2X6DSD5TSij0IRsrZMTObF++992xFVgsHS1wpoOxbxPVRh
R5rtOGD4nx4XGZMufhDOUr0NjPYowxEHtdEJRlNZbIZeu2YsHHk7EguIz/habW8O
8qhhZ7L7cFUBI1f10qhv3UxrJ9k47lrgfH9Tso6H3msemiCiZSu5fQtJHqYIbTzd
eBwT7hV2mY6WKVGPoyhxH2OuykEkAmzOGDDdzgUtTL7EtMQudIxgT3ycsPkLx9FU
bLKBBOhsfeh385hRjyRjwdD/ytZ2/Yzvg57yKMVIXWkFzY8Q0VJKeLmJLEjvzL6Q
Al4/NzYHRWIqszsevvFc7MZDPGNXRPEnEhbTNcU8WM7VghW1Z/dgBxQteXH5Gn0w
Yh8DdMbMyIN11feWZ6pokdstsiTVeJHYZZkdaJasX6H3fFy6oXS879GWAcYqFAzI
9kh7aZKSoRjyHNwqhFAJXnFA+jPm7Gsk1CTmrECbTgsB/UZG1AlKSKo/J/uHiGKO
VbUQCmqyG5E3JHnXxyWWWdIJwj5I/TPUjZSbcAkaQYdrc8JYwgrJ0Cf1N7c/E2HO
s59fLS6R12HPgwPdcP+BHVBU5wHmnCFLjtKhD9apNZUbOIoW09tjkFfKsZmUwJ3c
PNZWjqKXRTk2tM6mJBl/HbSDGCviyXC/IC4uNZbXhqYQtIHYEHkIUchr1XeSAkrz
UR3dU1x0GcbzfbQtNedHolGrI6LiI63i0VwEzPlG6HzHleI7VHGQSsCntLEdwHva
VTzC4NzGRmIEki7vHA0nwdqwEitYBm1d1v98kuxONs3KzQE7791HTH4D9+W7h8tj
ALTt3zqfOQHJNjxKTA+/u3aU6yU91e7VupBVtr2XwSUQ4u2nNQQBqa1ucNP3x2M0
yYNzS9FbCCQ55RswdAITW82REOyCt4aBKXEE3vA4T0HtLwhlTsGkqe60iNZBIvr2
xFiPn7zbQsX1QBexsGH7Pr2Q7EP64DTsGyzIybhKzkw4dMLKWmmp6vcAtDrI6+9O
2D1oXAp5eqMFIeZxElROmvLnJW3HdnO0ouTMVNxZ4gtfSRPH9t9uhbBsiJbBBX00
z8PQMRzH4asYGg85obdaYIobddxI5iARMsr43gEqRZR/ALVidkzZ+ovSDojtt1ey
jDtvI0dGmHJXW00RLKDXKOGT3H0f73IrU+6XV+memToDuR6lRU4kFJ6yvEbwxjej
ufp6j6lyL/047E0xZ3x6/HJUZKx/WrMmW7wRfxk8mQwlNf8y+zUlRyPzwfTS5bvA
ykHMFA2Ys5KGdAc6ml6W0Dt0oXD7RMaNSZNKwmBWkt01frWyRA4ZUZ6NwG6BB8J0
RcV7V6NAdBYq+0IHF0RhL1xgo1M3JQrYhkVLq7yJTllmZkFOZpGdj4GYl5u9NfNp
JDpwy91HgY5wCtzjNZNZGLAboMnbhERKTth5Vq7D1JFL8qcrng1nyAG7vinAncOq
KP7DWGD1tPxZEQG9IX0SjYMp8OZzSqefWAGpOWhT3MApUJPropyCt9sjXpdBsN40
0+YKPtD4gpAaK67G5xA5tEkNWDtITwXju9ue9bvtITc05yCnLuvDaIdJV1JffIrV
3zavFCLt9Xz6DERIzxTNIaCqbSThI6LnnQzjlhSJK9/GRwVgxk/5CSVfwv9rig/G
gT6YaN3e3Jwxm1Cl/VVe/CKpEIW+LXJbbvGykMPfykYdyRENJT0HO5Z4LOuI5Z3s
TzfwmkahDqCZX+pAYakHH59ZSMXAURPM+Q36dGn8mwjknwJ/PhJGG0ACrx+U4k6L
zB+wujrJUOme9jK0AyyyQIfbu9CRTQ9IQD8AnxnTNNH4f5L0IcVZcJJCpVJIP37o
W5ReTFDOYPGwCH1+GAKGagzRKYjGnqZnKNBdk+g/CEl7G8Ol2vSOnnIrC1sFXcyS
lA7tu15N88VhuIMDPfJHE4aOlyVciaID03mL5JfuVMyI8w3cI4KUIISY6RS28jDs
sqfOYgiWli2uQHlqfqdHUAaV3qz9pl7kD6NEd/zfbhpBqG9Hnp7LoyUBj/0BcZkW
H6LFrI8CEBweo32wSOl+SqHQHlKhu6sc9u3BqRx/Ar0IJXIdNLbILi3Jpub3GMJm
Js2OxL+WOBhc8gRaw0PFAIx+r4O9uQwjXrrmJlxdQo698gG8DLYjp6+YmslxfMI6
sWn3rY/+SQY88NrI27eaICQ1daIu76tC09qTN0ldFixIobuy28C63jjYcUsUnOHt
pIiaCdcO/ZMWQud6AS7rhJceSv/h3ZWL1UAFwo0ZtlqPNQJWjtxkH6gYOhSUiVRD
0b7/svDv8fI+yndNvUWcnhEArLrSSNWvLdamPPLZWGMehYS9bY/NTnovWxIEbct7
+kuU1cu5weuFa7ZmIjTtiFCLMQ0TtVQ69yKkL2maq+PTC8Pnea0c/fBU9QPjaRx+
E9+ithKRnytmmV00+H5NmYzfdf2Fne4nq2HDo2v7+OF0SPEdgffJ+kPzDAzorxxe
BbHsAIMUI3005O06yTfU+WNWaNx9jJKwKfS475qsyzIoSkkB+TQv938P5S0AaHxk
Cu7mgKwUYFJj3JTZC2yGl9w8rkQWUFDlGJTXW1fdxugtBSHE7ti3rFleCT5wG/Lf
W6Il+XQZ7yhOVMXsKoYT6a61i0iaNVO4VoUVcMXG08nHFDz7MJlci5oWWarh2p3x
SBs5T3iZ0pCqyMzeD/t3MYSDEAottLEyLgp3e852VaFEWKtj0U2+p8DY0mcxpR3H
F224MMYZXqFElMwuvhvZIeCOF4CyDIh+f3akpGlzmhgXMJinwwRlUtMPwtEnvSTI
06vqQ1dQj8N55JQWx0vMAh7LTE4u0tVponkip542Ulh+xzoVALHV0YiVwiOUFVv5
A0vjig7wWF2lTsvaDshH+yCdrGwdkBspJ3dBXG6hQt4O0DmSjfi4/firBKbj9I70
+63IUa4U+4u0/RAhR4Sj29/LfL704RDe/FhiTHMWOf0P66lU84t+/oJmNWmtf01p
KvBglgT7VFBHh+DdTg7jZs0P7S3bP5oXKsgWdQLYBlzQFOse64wDQ9ujC4u5dx7X
s0GNssx5ujjMWrUkPUbMVAkF0HPtRKynwxyWtoGDj/mrGt9+NikeE/LP4pCFXkZo
OgUH7pzd+meYFI62mq5t5sy1xD6OkaXl9YpUs31XPDBfDMAxQemmNpNc4+sIuOqx
rXJPFGyuUSttBsCGS2cZ97dG6mqTf8QSYXC3hhfukEcapE/19r1IBJopj5oGEud/
1MrTp3tQjedr/ra9aT9prAaFVC/02+MUAKsuao3BeSbRDdB0OMZPCDnV93blmj+D
X+HbPL9bRZNUh4x1ZQfHSBAiiX/q9ZoB5RHHgfx74aH3ok6L5h18ymdJ9ubbuzhQ
+jBHsDzrzIwS2BZzj9BHYvsYmpjn3Vs4k9NGCTPI21rkMDXjpofmJHJm6YgNGaQR
roj9Ffr0bEhxakJWrvHDlR6A0oWi/0Tg5nBMUKelBsT71DFBXpHbpPH85CY216Zo
23YEkvIiu37f+ygcJozlPl/JnIvoa6xaoKIrYqf/tn9BJchFiY7So65sBOvvSQ+m
7SvrCkSWXARX7FXtElasv2N/pTBEoaOFlRrgW1RAV0QH6zIie3du7D1Ich2Uh5K3
3qB81TwnKcCtAHMSrIi3OgeeeJudQsx1uAXKyn9Q22L4RjYmP67TPvLQ7XehGFC5
N63cGZwgeFfxRuVCzn366IhulbEKToX5XhlQ/wIeYsCMPRTBUPPKTrXW5MMpygzN
R0x2oOCzSdGKP8lo8Sktj3OMRG9iyJ7nOhVQBtL8MpdGjAKtuQ+5jIQJvISM9mW4
5LHO4OlCpNe/bFNCsq5DT53dlv0tMj3dD1vcmAcDxV97VN0cdSdvpXH015A/CXqI
S6CDsFVt0KLGi0Df8t/I+lvVBJ8Xl33p61pAE+8mQXZ9ZRFyxDIcBxHJBERqeAib
dGP+E+CRE1ao4N+2UyIY87RsqMMNS03LJn1fo9tRSkRyFzDege6FBWq/Vbq1wTPv
j/iKYRAAfNQchC/hTzNixKqQMcvGwzEbw5F0b5V7QADKYRW5Wtu64+FuFWf3A0s7
olzee3q2WezaQewjukPv/GhsQcgknSz4fZF37QBbxOeNlRh7XPFnwumnFJgHEw4J
l8UOkPfx4OQQlS/qMPBSR4nILzeyz80c2W/Ml4BJn7K3uy39OkEibbDy2Cd72zWO
D18dM4kJl6MIxFLL64twNpMkXX7rZbNbkHwOF3EbSKamXpbmg0tgOo/ezJ+bRSiw
vNVi748Okh46RNebJCUTbCJGwI60GllWeKFNs5C53J8pZUuG82XsJmS7d13SYdCD
Vm4tX4kFyIuPgolJ42xt3e4k3Iy8BDv7A2JuU5tiQCobXr2n9s9Bh/GaPmBOZVBo
95LI4eEKoIhgyGKHeoAjFqW6oD/EP7QkTiLS8fkcv85D685q5eCl/6+6nDMMZtDZ
QPPgIN6ybBXKvt2PP43wIYj/fK3k53PGCY2cI6MsZog20ShijQhVR1xgIx5T9563
x8oNXTBxPOZfHxM4HDLm1WLiX34dbV5rmtlBWnZ12O0XCvyHQy9IoguvFwtKlTrI
Ht4fUbSSGJ1d89qwhfXFts61P8p434arR9GIJYP/ZqI1rhUjakZyamuVhOLY8Uye
QfMRQW5oIPxieq6O+5CiwkYtpdUCnOrgLCJJ2HQ42frCYs7l2+EXt8RfwlRrjnk7
9NhXbjHftQautGyBpY782ImQeYGe+l03If/CMfACdlkqZQm2yfkxaiZUejkAe72k
1MW4mfbi3trXP3inf0Wvgyktpd3AbFhDBgLAVfYJ6jQwch6h6DDua6ndAQSccoLi
XJHHLO2drudMV7rZGuSVdPsWEPVqDq4ErVYknongsokI3Wz9DhzY5Ogw+sCC4S+Z
GSnO8b2IfaDTBxH8dgu2v/0wtpBeK+FdsU4/lfQ5htiExB2HMCEicqIeaPYHp1xI
+18nWsQZxep/89qUgDGXNky490GijgVYNK81Cc0Vcf5lLczytmOveu+sa0XB4mvQ
60GZPezSRS+I+ij4auNtLKHu1tnHYXqSpeb6zA9cRqFhskyedh2vVDigJZ9v5Pm9
hQSvrPQhtJOSis60tC19uBXi1Cuzhkk4EmRfidI+pBGzv7FxrWXJjAadBAc36n7E
xr3HfJpNpYN0tEH98uzOO7h7RS+UtoO8yrG9TEoH37hhWoO51ckj4+7IaVQHDMUm
FuXdP4RR5Zf7zwUcw5OwY1zsAflzDX9mLdHdL6OouUMrK870Q6nToNbhrHlh0XPS
GNWdPk1z94s6smxalqyf1W9AzWLK4P0ASpT1QbPhqkgVV7CQpHsV9QcxaoI3Krmj
XrSNOlPp5fZg0V+ADZKk2TqHpf+lIuuO43xTtWa6P/oIU08xnvWPoohImBVBzVQH
bQRVju9yklsd+KN8OjD6dmCrKYQSG6nAEyZSfs7dMz3ISs16A97PEqrkviDeHqi6
o+t1IMYufLjmCqLWTKmNgqh+GqD6hiSsih8zRzATgKAjP3tywD/SQSgHbUKXvVRd
XMIfbY95HuPnkRXWxVOlhEO3SdmB5VfuBYD68iYShQ2w6CjH5Rfrie7lnJbGqbhg
2BO5xAjG67h2rTqBX5jxyGK+6OV3zOScgZorAym6VfoT8s7xH8607pb8NYdkos09
oWOp6+pcgiwOTtX7OajZ+98/J8xsUgue8WLlhCimh7lJkX9g86GIuAbreB5pQD9x
EnxWEFWcN/Y4Rp47JVioxaXWpSXlCLwPgRlPBO681AH13+snoAKcgsyqVRWLQvQP
2euDDECl3eSqgYVTySkMOhI8CR0uj88x8h3RXumPg0zp2V1IdH/lkI8iWL8FJgD2
1XtzIpAvVZcJu6vw6K+ccSR3Q26Q8vXU/4HSUMSBMoqBzTEV9Y7tSUgfkhf5u2mu
9FrkDFoaoGCiyHSaDQXM48Lb+/YZE8HlXmjAwdq6uh3ah2/tX3BHyzbOSS+lXNvg
/1dNROtBEEV619Rm6jc7ygfekGErULX3AQ/+wqm9NaVkYWirqA6XguYzTcGYfKHS
6yLRzozs2OlAcX9+hTfqR18iqb6fqG2nHrVzkXMDlmpt3K8ZGduR9eMyQ8Qvp07y
d/p0Q3osPiBgRd5Y9eTepMHZhDomA7V5bXIaFGDNcayCy6ySe1WOkYDQYGjm3P5t
V4XjReLwJB9ItfrU/W/QuzO+mHaqnaqzjIr3YsRyiWeUL5yTE826qPdyZ2izo+rA
BQkvwYfwCge9aOfWYYp9AQO3xrIWjpF7DufEqU42zmIZ5QjJiGA1Z5srmn50fw6E
RMek0WkBdlfhW+j12pSIlMN9anDqE4db1ew+E3SdREk/vcGfD5ozy+5SXNHmlty8
6IhOD+LUAovIccapThGPVNzKtI0CnV/GgMLcCNpUhz3oRjPdFe5nwbR3G6YbkZU7
Dbcuf0yKdQMyp+iKvBXuPzcLHxDWUkHFb/KIl92m/Q0fWxaYaooLwaI1vT0fya00
MxD7thbfG/eVipygaOS8Za017UZMCLNDAavlIo+N07mSv1+R5nPWYc4dJ7TFJUA7
Qy1gPOvIzRcfBmXMpfFEsR6cwcjQ8IVT+aVE+q/2z2rI3oUk5ql+oas4aZTdFIWv
5pNTIJFlbdiZX7nDOQ4jFWrp8eMYShk3VLJk8ookTgZoDOL2dTpehs9aJ5ywCerI
6L03I/P3cn3r84Q6Qo3zTpz6WPY9A4e+OhRhZwDt9mSHiwmTY3jPF9M7uhxo4cCz
i3xXn7UyyNmQIuiyT5g7i3RtpNvNsdU7TsLHtgoY7YQdV+UdYIebEv+kWRk2rIwa
WCkm8+yJDjPE1JYQGlYosoacaPN7vJwKGPzkWAbIMVCKq8Oglyck3jegOBgc8S9F
EQlcbuxc6UimO7YjoW7Y1+ksouoDXYfv11RZquqP2m5eTlbB8EQzXQMYZs8avWgt
wzsHcIkPOKUkVqtbPM3lmj5tzoE6kXarwEAc+FLq7zl9awZtmj2y5lwN+rHayu/f
d+3tW6lC6yF2stojX/PJ61jMgbmmM9xh7RPRjvXF7UBzXNy6OYBPn59qNDBt6HoE
YiwbpswuvfZ3PNYD9NqFWM0YND/Y//j1cLEtqWD2AyaD5P9+p+UFQncAzcsonDwh
2zPEtMHsaJPCcHZs0cJrioaV97ObyKCyBHj4IKzOS7FbcTJ3Jaq47B6ecir4B9p/
YfcJu+v+sbA36d8vM2ZSulJuwZhomAI3xCkp1r3rhDnPuMBlA+B6YastHMK5/ECB
W6pbcCCUxenDbctQ9V+f+kEY3cJ74AAyf1qVtiHhAEnnwEEk8qybfZ4xRXJa5f3E
gLnf5rl3avsiXKaFl8Hqb6jaNpScwraHVYfh6IPxJiX4l3jkmkbF1aweRtC/amtU
GkYPFdimtlQeGA8y2oAXqhZmz2KgDBRbs/rLf3CWFTIs2UA+LmyMeWOoHHCGPypu
Rp32elKGTIgv5vruriiuuwI99zIDKRJvq85bXwAE96IYPCw2qHzlmUxAK/km1JbI
NXfa7Ljzhf67FnCOOMSBRjJsT0c2ntP/QXdRAWViIL6GzMrtlLlMY7t98e6azSkh
yz7E55Zk4aarJVCk+UCVwJ+XirX9zYEHKgHEI8hRI24fZPbQ6miPxMAaa+/zE+/u
Eypuoem+ARs9oe8LtTcriDF6XgCVsId8/kCb5hgl+9j4WLA+UxnLklFhLyVwxj4x
vOYcfbN1Sc+A9o0KwgQbHgfCMQpV7acaAe0AgQEZuMUhB+y+Au3RZsnUzcc3Apf+
V10Uw9LbpzUr4RrPNldiJoVoRrLq2qJ4qvJ0kWywUL3Lmc5YlGlmx0THNR2kx7Cx
JeNuvi6TbN+BpEvmKscCDsq8Z4rf8dcdJ1/SJQE6dld0xEwxK4QHUU4usdXztd9i
wRRkO89wPpVE66zc3TQ90jP/2Zqw5R59YGw3hCqr/8S4P6mjwBUM+xH+OrFt4jTb
LFurs1SMSHU0keGwdytK8LlrtLhLoH96QDNnuYBpmyCMVEDVmiw9OmCnw72opbjh
+UlDMp2Gbefmhg8vSUNMiZ9xlJU5qhZmc0iPksN0jtLdLML4Q+q+pxj/2O4WNLRh
AIK/+yHdE1pxDOLwYl0bg47FHq5JzHVHiB6fk3KDJdZBxeL4u10V1eJIEKYy6KLw
qbpRWYd0ubH0d5rjnIZ/xmbm2s8CcceaNk1+r0qI9dpNd18qQSnn01TsndiPxlIv
9XLfc/1/VfFfdGKLXo2Ti7Hq8rVs6+VKhAT+o5y2QRzW+UF6agW6UP+NNrwVfTyW
XdH0VbUzq3wjY9tV1VrqfQwjCPQZa8hoQUzRZGKPc26JMXrdn3U1Q40N4A6pPLEm
MgXqbGsIhZxiNpcpRBmk++axsaM7XwsNqnVMx3HeYW+8MJ7DJoXx4UgiI+GjfMsc
w65iwuHDSZYiyE9KWD9SfT2ANS3oY8cUC6aKgDHo3hrmuFC0wVJZah5JHB/IoN1c
FzP5Dm6qCj4e2GUsPEV1EcPcICnNCeTPvgYRVq2b8ps3YjnK60nE5kQLuGasFYUx
GQofZYEWZ/4+ZYWYXM0joIBPuk7FlVVrqPLlLHPPC9uc7Z3R2HpNllA04zB2/Yhy
QF5VfHDbLxL4ePJGau7sqyEzOMOwPajosq/Y1PEkg5scW+uWjawqkrn/os648CqT
0POsyb1r2XIhE5EDg07UtFe6RXiVGjCQj7wbHtkjurZGIIFH/iHVQH0HZXzVhu6t
fAcHX1jn+GwrFVmFRloFH9luL1bjeuiN6rJDntAJI3PvfADHW8EdiAfAnXHZetmo
ktMCL1PTPkVhxAXS/pJh+xchW0mOfavuZlWiw7eSbmr7JduAkZemfdb3JKwOmpij
piwDAwi+udhcFCCCVf26I3aavgOgFZJHRcET50qfU86IAzBWP7hKmWNq8eqKaLWk
JVo1uEyo+5UZdj4rofoSgN6zl/OXRhwPbV3eUWkZD6qDZV4bKljUyIyYI6+ZHV++
Hclx22VacFevnm0mpXUW7gfHfGvJZTCZgqXa1F6Kfs8qSOE2tOmjePXHBPyzHWTQ
MSo5fIAbXfn9Bd7nncQRNAQxZhW3/InJDE8DkmoTcw6XDCSJcPXQBbipNoviJFY5
EhyoArQ0UuOXKjZjbqqDZJMWIqm+AkX6pil/Nakm6IXDyejmdzAwUK+k2SOLq9DL
0jBu8xcvQ3lO2ETf1ddTQ+ft9h9b/s0+Gdz1HrnidZsNZY0eY3YO39tRvp/rJIOq
lNgEc+NN415owP+tdkIqEA/rp2oVJ6MBTZM6/BNv98RpuioaaydlFbykz+e9pepM
1+mo1CBOYPJfS0Ua1qyowdlFUlCnHDSk8ZHYYLnGtbz6u6e+EMdFaTNnK1wsqKuL
dwTaW5TaTeunuF+eew57CLRz0IVciPLmSC/d454c//gvogEjMffOssYsXB1y/agB
YFDoXreUH0wy4Xo4a1Okrt4pnBtmX20m1741CBzeTonA5EMm2yOif5T5qNGEuEwS
oirrcI/giG1x5X89RlW40JhS9EHB9kdN3q8E9eQs4RSVeMM6ljrfplfIO9kmhwey
XwBi+rccnXoYr09klxPEMe0C7IEBnCQGJKNn6metKOMmdEBWncwmwumToXNn8CLe
/lDR8JSEZJ/z0htkZYJ1Ng8tprcqVOp7iDVOw6w4kABoNO3nuhEWUXa1/kjU7ryD
0bhPsvY0eoSkj1qUqKqoVfQKpimIYwQhSF+peRC3cNecAE2koGljIOciujx2KzV5
6YoYJCAs3XKUl2V/LnGaKO/N5OMMsqKsPrQi2iAtp5OI2FoIPpH3s0mpMHyXiUWy
iguLUxbZ35aR6luRHezrs/TvFaAH/5F64ycAxyTKVNvGHw9lmoccsbXm4fXtwZfb
7U30Jiv9UDd74ry4SUQlivD/Yceel1ZkGzUqOAmG2NTXLSk8MjqUoCrlNpOCshmG
vYTwl5+QDys2iAexoBKYLIq8bCvPyOIzoK1Gx3t21lTCPrr91vusG3mc90N8TS/y
BiHYtRbCpXoWKFgv0eAXjUnXNVdNGMgvJCEmJ30AVQxXUy4hn1rVxXzE9E6qCQy5
OgZgHHMK/IhORNw3APo/DrErO2urYjij5HKiYadYSyb24LmblCQ/0W5PiMQdOEU+
RVE2qGGFlkrposg1LFrKdS/W9F78MOAk67sjzFT33Qq6lEv61MWwgomWDiPLu+jo
qHsrQhWJV4btFDRY+fSGBxkWQonw5vdsGQx226J46BjHK/JasS4NNY9SVRojU6mN
QnPTgTARMNEPX0Jg0ix6ekyQZ+nup1B3gHSkNAoNhu4pkShNusDeYOgjJWG63pR6
o1RBMznf85LgyGEwHEEmXGcyVvBUi1N0EYVVuAvpzJl0Eec62MiPscXDTcTkZ6qi
sbrDSfdd8N7Zo//pPeh6X2arCM4MTOZcYSfAN6qjJq92mzWqUbQER9Po9WnPQnXP
lYkBWm52O3JV5WeJ2nL7D9VKF9ttXh9nbg2yYOG962L0DqrJhfhrgkmruGxLjjOf
T1X/pXIYABY4lz5mYnVrYk6BAuF2SQK9igcej2brAp+4+3MT6eBl0KDzJuFOqeYt
/KUKtoOSud9NbTAdo1FzScO9k82OHcIehSHmFMCTwVoRRoKc+dY7OX3PcyPaJaMP
I1wxTjwkw711hqLxY423vaa2DP2Db4GdVyXEs2Yaoed2aNd2KIY8CcUWFbS9nX4s
FRe2hUgk2Nywp1W/qholjCY50EofE0AiLCtWL9ycZm0ovtNNeVVLvV5SQGcTgGhR
oQQqcvRIRwydOVrW3i4HFt6bAjUfaTFQuqR6lufrzmGfoaJJrWhsWuxK21pbUNKe
cHzItnEYTBtDl3HpEr1245KUv7rnagWKigYH6ZGGJgvdo+Ek5v1zY5JH85NaECPy
ByfieTGgc8MhuMVZ7qC49B/EpFc0dSxUf1DAxmugsOIvxYVOGtl8zTbqg1+GWhQE
Vp29DLse47V87bXJ0sA5VI6k04zYxBATv4QM4dKPjyOdUv58KhqHoD/n+UsDQQmf
FvGURdv80KrcSzwjE+4O+Rq+iy0XwCpW/owjVZ/Ddq7cRWJySnxHN6F21udDfIti
RPeq9LUBIY+5dcOzk+yZga8j401t+Hx0d5dFdXD5E3eeRXYJNFB+0bU993QJ3x5/
WJiUq0iDCYI6l9zjONcOLFWxg8Q9Iog3CNOnMKaHLQy6K8WmojckL9UPjIHVNkWF
0/Iegd41rRgRPxFUhJCyjYMtrqSSNfhKewL8N7ovHROEcoxlzEY9rFu2cm9UItnj
xLjIVAOrFdjyqCoHfMk4kzv+J3kVBay94pJLn7OBW2SWJELG2QF3Aw0ovh0zg7Nm
7BYi5g/YM/xhAoowswQQVOZVPzXtkM0Q+1GewsSRI3g2smkibnH4Z1nZ5o2lF5VW
xw1StcKfBMJAGxkx8mT4zq2FreuAxDzT4UuvFCfFsZ5y4kI6TFY7kvoYPsInJdz4
iR9JroYdP2ohnaedE6yw9DSCVQGI8UQxkRHOfMWbYavOtrS5Iiw35STP393YJU5Y
QwCBs2P4h4VLdUSVYFDm8A8nWksIzdUjeVvOHe+qVMzTgdbs/TAV5I6MSrKuakrD
EYpspvqovKrFZzDs7xTBMfrswmQ3MJ8Kvp4pR19xw36peoxsL/qoumxPcwZuiFUg
GVQ6F5bl4EP1vUjo5MvO4ubHb/4rAH7pBVsCAx5aqO6F7ciKBTH9V8f2gfh2IE6S
uzWNNG6Qi++fJ4pR6V/1qZaMc2da8b03PSk0IdV+lYlv2eNyw7myooA7piY5Uijm
eh6xwJaBTLp14YVgYdpZHW18QnkUrgsB2lOdO7wy/Wyf2lEss/p9EeTXAA1W5FKq
KFn+TF4j0/oLkfMdNVBg9OxbdgxiV90yEedm6VywMfmfqw4hnwJPN/uY3XuwzXo1
JVNNEyunoyB0bdGSceAo9TyZKbctljD7WMHmYvK0At5682uUeaGUqsSkPiVmlgRB
kYdnQUo32mOtlOxNLKNAwfbuCYJuA/h6vMY5LdQlzoRcdEdK9U3XTBAiZvLWYOyF
g25X7xtIsSMaN7lJQ4Y3EpjjsEKGSSps5w5p6mXpGdTPsCuLiu7UMAQsSJockc3O
R8ID9EB4Om0my9CdU7kCTj2hGnA1x9UBlUJ5KRM5Cxz51FDSG9Z3x84BqGYbnR5n
HzM17q7wDiS56jD3Vk0Vd27CZSPvU/E5NJBcJIzgL42Qp18VECm+xdQ7TFfOJcdW
FJkH6vsAvuYgWNpPrIOUhYcg4vCCF7pHjan5BihmBxMDvbbyNrJVeX8jJfsQOeg9
tMEB7t7f2MaKcQEOXedMhI2NSHaGv4uhEfxOvwJ+CctcrbXn0LC9kJXyhLVJ6IUD
dinN+YkzmXwGEeydbPfDgYlL713el0wB2I5UWZsA5UeGlMH+zg0wdEFmHz1Nx58E
M879Ri7C+em6NYfoDTyS4Qwi+jJNSsxIwe5L3+Pza3AOwCOfAAUdQGRfpYhFai9Y
/dNw2fM2I5i9W5bn3OJXDTlMg4s65nxtivTXluPvm/0ELOVb4bdPs0Xpwioxzt4J
dsHUDVVBOR5F10P5nAlN2l+djlt0eFmC5hZRNj7YmLTwDwU+1kF+oy7kWXutdAv4
V7JmneUqPyByLgwWQ6Hu7sJPcb+qwXuv6gLTdGmkk6580QRBs6jeEvOrOBZKsdK2
xHpMDQgBEkEpQIY3J5FR5mrjjztJmp4SLL7DPKEEbD2ktWkyX4cD7evEvrzq61Rb
Qq0R9w2vFbswKo0uny8oauq74tAjE3A26AZgPG2ENKDoZNUKqKcMsWvuu1dLWq7s
dVMsJaEEVs7Q0LeBKCQUzRUT3bA0RH76ozUKNMzUKSgsMqSgI0xsrpLEmQ4golwp
w2bJAc7A10d02h8ypLsU22QRCfsUsq0JdpNOxBerWwcA6h0X8fgRqBOdBkroQDrh
TQQHKn9Hlt7WdBsLYn+XyvrnGs8p1+Fqz2B5qbWLwzinx7mzLM4fEM8WSYPQ/fb6
2JZ2c5WNk24rP+3noLT3nGzww6/WPd96JOc990jp6373YnH6AQ5U8/ot4XFVl8LQ
vbxcerjO9YJoSeu0577PjZpP/SV3bZ2PlLjkWbPZoOKmn5x6hfCynkTV3nGJsnDy
WHOS2yG/NWR8+799I5sd6RIhj5I1EtpO2Fh+9P75tQvN2pHSFMdP5E0X5RnLQKYi
GBqfdIroe2nyUki13Q6Sl7XrfCxq2YEiSG8PCVhJyJLLRr5Bj+NPjshED+5mRFmf
W6+nlS8ylrbm1G0/2NDAY988oaR/D6lKNNuLPXt1R+BOBmbM89jGVm8UY3vZckNQ
b90kYy8ma4nnf1XKpCpNg2yvDMU8LPoyktHxoqJwxqm+HnqW9M8ZBhNZBEq6dCSC
eZ9cWNEHEjYT3yZcSAM5XUi3qJqZHB8ODss2KS/rf84ReISGveMNsMi1iu8U+tVA
Mt+G8iLQk/fFAKmt/kGWsgA2a7ViMbDh9Lp98pe0GzdusLkZSxNqs1+xIV76XRou
tT5k3MBPBue42ZOinkn8G+vUt3vaDeW8ciFM+uKBatpTeeTEHMeMgTzgObNhkXdb
0kp4sij0lRYrccCKmp8zqehn8sUxEH+ydBjGTLdKTwgG7FL6GbI4SXqoNz+2fvJx
jy9N+krRhMdEofaWQxj5pEXLvKCEPSCbcH8CEloiK51dhrE183//brWqwZBM7rtU
1matwtr2Tl0R+MFCdzwJdJR1vGvBhQ932/QEQJGlDDsexixsqf4fwMnjyVBDr9de
51SWxNOQ89t0/Esz6KE0gt4+E1vIS7aTFIhZSZrgGoqA8RQ8Ay+n/C55FsUo7zwX
RhWHYsF8ql2y2dpVaNEpX02YUCcdcG73bXm9Gp8t3IsoeRo9AwFCMX8m47PaHnS+
f4KH+e6oh09PXKQEstV3IE2oBg3fBylwGvhudUokB5oOf/adEDtY33uz0ZAc67tX
Hme3SPCo0fZrGcscjSatVvfcfGhI2bnfeH+Ly8SFt5Rrpyg5Uyn3fcb/+ADFFsoS
IMQvz6FgpGX34Y+RyOzbpOFCotlF7eHEHKbNNlvidgJv+S6dDmHSIkfPTwRGGWdT
IBKXhCjmVhbjqbSxuBCOVWxz1tsZx9kxPp1Qb5R02AoS/AOFo239wAk0tyhoQpwp
6cFk7M+NYp8PvX8HWxMU9Ad15D20ypJVlYJBxrV169h2vtj36xjr3tFtGjLtIEIF
ioLPTJC27Ifc2zd21LV6kJchWcjNHfd0RDwPrmQ9ly1mnFaQKoWUA38QYiJnz3SG
JkNGuLObm4D1j9wGklx0QeQjuoRdJ73MB8nTgrTV9vNsAUmaLXJtBw0AzLYh49iz
MST087T76+Zjqo2gHzE4MfUrjHoIPhRrnwEPZgYe3BeMlNoFpQOvFLbmBnFi2vp5
Gc+4Rh5NQZMkHfRvWdCZQlWpZVaPCafpZd9EmJD6wkMyWBeglfD0EzorqllBXLUv
2QPDY0vEP6Zw3rT4s4NcrjNh9fV+U9TUu66H+wvisvIzyiCJESv4GwxTz1d0a13D
ZAvNiLfOEKaEinvZTtHKjf5/2Ehw0uC1g669/lIx9aEaTSXegr8yqm7JfCTduv8I
+RNLYtttWtW+k782QPpAMLRLnF+g2HnV7M1w2pKDgQl7XkPIucIdYflFlWPnOcjc
v6XJIPxFPu8Fu3zUeGae/8ngWRazy9fMQXYJyf+tW9Mr91DTL0TzTOA1VHFjITw7
/35mSJY1FiijMp91mJc8kfS5mN8uavZAj/sfX7TltWIHXthE8Af3vFGYkFPK2XDD
MvcZhRosUCsCygnaALf64qGQ06OOsnd1Nf2jogUv1e45Pu92i7oGHO9Da8g2VtKW
C6X/FDaoqwiAiXcTwz9gtJXtuOC0whG7y2RV13SkGZ83EkcF6VrqYgYVsdDSHglw
awXQ2fL8r4rvlYMdCf+Ij/DpMeoM/BU5iUJCPWo8huhtq4xh+/WZrGFZ38l7tUPE
C3YfqK6Gn25CNTwYr1wq1w09bWlCGubqpg16G5jB+6anA0U/AGIsgqwbmKWMhEA1
3iBOiYUI4Muu2xkwROCzskAKul9xaHnJPdVguZEqrlQEDrMgTa/yZWdjctT/G1EA
Aj6ng1V9kljL4Fg8DlibW3DpvmYmoCumPqQH8f0DBdoAqGK0VxaKRSPTUgAIoB/a
+HJD6gsRIFVVQzn6zAJ8FswVZmOYOJy2jpb8lXXqtd4fjugF5+NDjBpj1v1XM3s8
hkwzlnC5H66YnJqh2uK0LD0spkI+bFTCtLf6z/Y+ABBy7TxQrc7RI+jn1PKSAAMs
8s4jV3yhAIKZWwuy+/JD2VooGU+DNd2dRV1f3rQ9chH39rhWTX5oJzQ7FniIr4KZ
HEGtycQXkFF3cfg1VOuwV0YN/iKcn/3ul711tusG1F6u7lkRv5j1GikNuIHrap4V
c1equl997jOVaK8S/aoeR1YfC/BURdc5DOTZpdHD+8RhRG0CDvUO/e0MsPEkL5lN
L3TSnTxhrRAZtNvMxOGJSef4wlrOp9C0C+8E7P0RctPNK7jqgl1D2rlqH9/Vb1HC
q0yFYg85bTgS2bO1DujlDnHS29WyJQ4NZfNrzrNjn0+LH97gLZA6Jz+hb1YHW2ML
1VKv06w1ehNR892/1gc3Pbuyla9vZHaPfYFLEAyIlUyZNtReI1RbGZye4Eg4eoAr
2O02dAeh6DHpbVV5hnPBPzK8OvemNW+OsaYKJZdT6txgfN8+wUc53ba+L3Fm1VHD
BiilhogpNIgCxggVqApYtKWth5okNC3NusRvBVQVnmLGFWxc8uVCtDB7tGrAXYI9
WfmqmxRcv82n7PnXcbKdQmlQ25urU8y0svJBJUMpKEFYAKn49d+dRV6mUQebklRU
EeNDmCWdV3Op4ZJ7jLA9AVW6/9LHPllASzsRLrzFExLyx6XwcPpT2PasNWUcDS7G
Ep8/cN+0HKD6TX4oBe+exSjHxKXj608Tj7Y0f3UuuSlIg3a5X4vOCeqgyyGE9Dyf
9kSMVzVmSM+Ylf4rGqSNAaGtanOAedMrPM1/LZOQfFWT3iiScvWVQ9J/Hko0t36/
L02n271WJYhBYZ7lFFyve4RVLR0DAR8fVtWvCvh6jI8ZmoA4TROQcHgGuaGwAg+0
YoxkNMyApeI7r2RRvIcZI8vwpnvo+WhNfsJd5OWv16+OSzgsZIc+N1cSd6mwl9DF
rRSfNtxOvKI3N6aT0HLXa8DbwYUkzfTIhdutyHeKz43y8qYdJrWXEf08JT3pO01/
T2oQFoY97KQzQ7T36cuZYGXkY2uVdpOF2iXF3FaoDqkYDmyic07HNur37nFwK812
0/tWW2yHDtS/TlLjc7X67Ao4ko/C828fk00fPME1sG1HTuMZ/9Z+OrUD+qowvFhh
Z3sXSmRA3sUK/JV/xdb0rJ3+eKEi6Z/TtX1tEqdzzPfFqd2oyVwYeR7ylCNg4skp
eFsY1j1sgxfe4CvMUvaEfYvewVJCl5feO3WGtBZ/Ttwgy1ji3g+/gjegXm9B3Wdf
TVSM9LPXKmrKwfJBrcTPgDq2mr/f75YAMugJMH1iA3NEEM+bErQr7pSfXoZgOPzX
gp5sM2mwJnh9k8YSBAolxpJQmzPpmsU1FoXseyJ85hWwsI/f8qRn6PQTo+nkAgWr
gE6iUyunixraLUW4JMS+GOwLWb5EbzIpOnhgJE1nC35Nx60vbMOOHJmz8L9GcUMy
3OWJt2RfpX0Lxe+Rh6LWMHhcRo9WFMa0QcuvZ6XonUfEz/GsYMKSZTc07L/c8A1e
BzGX8Svgr5x8nyFnlTPQ/4P8oX/u0FpoHw7J5D6y/LsR7E90wcnFFWyZ1eihpnUO
c7wFFNNotL80J8twPUD+wm/rBfv3Hp5IT4FPmZemxdtHx+eMECxgLLqOYB+5FyW1
6E7VCWt4FV6EVgs7dNGc3Ka0gNuMHQzsBKdxk/9vMusLmqY+WhM7HcDadEedFs/2
C2l/Dxqh7FNo7xHdahBZg2sl9V1ARZouBqPKyN5ssK0UNpVnrH94UqaLigMoGj37
4czapqAar5OvVtv5lfZxFC51UAx3O4WjWBjsE3mzQBFVZ/pzHdMscWY0lNGtt6A7
NIhHsulgvZMsv1AZu2U597rVf1vgO3uB93BJ5ZAdYurS1Pu8BEwD+Bi26ttJWSCR
iT1x5Vc7qaCV80JC+BbiUZMlkTxeCyS3SfyC0wxES1sMUEf89SQtJl2TzvZjg4AC
Rv7ciTIkH5WalQWBvbimYTGNIAhXbd0ltWuSJbBf1no6e1SvZHK5XCC+vQDsTwaE
7Hgw8d/cYx3pIC6wXkYnzq4brD/4udN0IZcO6/RHYF54vDzI384tesEQ7fYG/w+l
Ff4ZazdQot/6dtJLT5B8dvkxWhQ+SPpuRqABO0oJmC8Fjrp0WRkDSgH+72FZg4lW
AWVkOuCYffbsHKUAIfa3TE1ShrAaqhgRwY4XCGY+aZKlPyC7kwPavx6NyfpxqAYJ
GuR2p4ZowT8/1GqmES1WGX+vt1OV5JDtm6gpYOeCLH2SZhTNzneQf9cHHpzsQhnL
Ghz0IEWggjFf3v33qvyliTZTQgzk/mJ4DpZNDwNtsBkEeyeQJDGB1KAqC6qy4DS7
YZoMOTzAo08Y6mnZOQ1KBEj9mx4UPVwQSUsYlbaugs1VfTqVCUUuR3NwZ1/zB5bC
teFRdiQG9EdWy4YDSS7sXxKnzOmRGVE8AcWxWhuRyonsD85R8iyVgXquHxYvvk3H
vYUKOUkEvMFK9GvtKWqNC1CJnqNlEZXUpOCYL7hnbYqL+INXkV9KC15A0RD3BE/M
0k9gIXxlgWEliN4880PnC48e/moE5mshadKbI3ia5tLYlMCwYO0RqIOnoUjIZ/xJ
52bAHKRguBqwgiASF6vwvFd73TUiO2ZgJ8BdZL0PChn73gXkop4wVL+PAHuBxmT5
qGs2a7dlmhBVgzb5mhLmMRa7v8BZ+YFg7I0IYOLUJuzsbfJZDgnu3bNmGBoGHNHV
7/p8WmXvVQQGRu6J0HjTrAD+jpolgUm3u+sbS38RqTco0j8MsuAPeevocTr7Tcxt
JXE4+khfWQsvIDAf7I5zWbUqpg+/s7yaDPBw3LTy4zGTTHytQo8OCOMIfQKiXHxf
xApmpgN1heTnP2/fGYSW8BBEE16FLOLeLlkFMmE4Dlp95KbCeisT8HNthMwcw1gR
ynW/khiIygXMaXySw8M8r28NSlnAvMuq6XKdGswBCoix7/OkAD08mSNh+3TWRRVc
oM4X+6Z2OruGgUk/SF1VoAD/FElRjSyhIdag3WijPN6BjHk7bx5wM9RJu8+85fsU
EHDGW6KjLsFvMYr6CfT1TIQOkBQg+C3/m85FoOQjd40tj9uTNz3kWYCqqpFxlnqz
aLK6v47XPRQMsSpo0fRhNtTs4L06uxpBNDX/1z5vghPz5l5EuAAnZIc9qQC+5lox
kGuer46hrUomjkbGgIrN9Rh8YWn7uPLQtXizgAQzEWYw9+rmp8pYTxM+OvD1scZc
mXmTps12T8qOU8SbIgX6wgUJTtrcM1k54ctr+g4I74GTd42o/4jjvKrWVPH+q1+I
DDKZEhBprORvO9lZwNYKp5UWA6KoB4jqQxeDKZbBgPlGD2z+RVZaVhz97G8XslHo
dq8xAaHHYM+nvzLfNnkkVtpCX5Sy2RRREsjZT2MaJAwSVfAzj2EZ58MpTza7XAgM
cnf9Bq4vVv9ZAnNVEZy1wS4Uj3Z9vkXJu+rmDCsnHHRtw6aPsxs4cG5Bv7nJCGWu
IjJ8BYZ5PqzlSx3Bu4PJC8d/ZKZNR1+JTCfv9xEZXjnVdXMxJ2KG5f7Um+iN+ahU
vq8Dvp6O9S4j1sXUQR4BAZ/nV7bzxNJYXSOWIzxpZNO/fsVX5JYBr83MIS3Arfug
+aAp2+Rd8gqMlc/dTiS52MkInY1/QO2A1VHV9eiui82gZvsUZP04eAh4ot5IGSrY
6Hw6JKmxCbWbO6zdMzV2Rtz+gpMB5MX3VqiexqYpDsScUbKarDNpn1E2SrewgG4d
6yOfxlvIxOKzo2qD13+PFZ/GIUyu+8J8pcJQ3QlffvWxzrYL6H7EZYVHaUjimdSb
2vocR+MR/E8NQqqIOsWHqE6ZntzsgUnII0Ckaq0UYdyr68r0fgv5u9uALsyM2SG3
S/gKkZY3McRMBR80wmTdGxeuu38IpjVar4/1Xg1fInYdCTuvw6mc54iGRmYXdPSz
rjtL4fOfuJ3DHb6Xw0818vOWss6XBPqrUXFrr7uWCzJz4qAi1Lk4IfHgbDo/QIXA
vew9OFwgNFtnginsXu4NgWLHspJCZ9azxx9VHPeAzhu6te23fu/U9yA1Vi3GpTPk
qYo7eBls07ov+Y4Awt3oZagG2J+DatyJMnJA2K4mad0crGdjzZlVZd3oMggRkeEU
jxj2rzEt7RFK2Yp7Uct49SkAOxTvs6eWcmcpHKrjF91COYbM51x/JPHllkqpk8XI
zeZnoCUfJe9Pshu2Mi0z7rt9ft1kVe4KwTlUHoozqgVCiUpIBKkZoGxDR5e5X6qQ
x1aUN7Bqmz1Km7fECQNs+L4GlaZrKxSY3WGYlQyyK4kONnFeUd2FIEzf5HhMBKdw
YLrEuXtHZD6bYQlN8XvKu17UNh7qcmnX77ReQPBJsuXGs+fK6pWuk6Ge5QHH4HY7
7h42jfh/2d2bnNjtMssTooExBKerpZdkIfEzOFoZ61bRaJDmuDJ5Ek/WVsuFq+O5
7GMLxbsGMd2Hw/F6+Kwd6TY6UjGCXSsn7phbZ+OYU+X6sLHhN5ChOn0AIGo/CDS7
oC6+vfIyxrDXvAo/DsYqupOBwAU2qAOo1iPrC5r8GvA/hou/DlwUMofpaHqqpkPd
xcgR3fFL2v1AA66SMyaCqeNo9GtxnHl8e6QLrxyQBZrlEKzwDAF+BE4FbBchKEv1
bHqJruVH5jjXwg/qXsDCfSG5JmqSDTCPRMPlNMjTMQvsOmuZWQv/uJr989TYKMXw
zar4BlpwO/evqLr7F4nnrWkE5XCJ8QRuO7jegMc/vV40mZYNv6itjWxgJ2adZoEv
6DW0I+gHUBWJRzxM5xICzEiC6UuO5vpBdNNllEXkWnjCqoumOfJTkucmMXLNqC/E
M0Y1Y1iOJ44XUb5Y7km3dbw/DL+0AWEkHo14P+DX9Xo87Pqc3K6j0/5yL2yxlB+c
U0ZFCLSqleXLteHbmU31dMulXnx0BgTxleHjrujd5FD4wm1eQqvRGZUDUREPCzAo
RETMX/h+nZ6pJLFwNyGTP/J1dUGaaE2UN2DZDgyxNlNyZ3v24J2T/4jLxgWXOPI9
nQQDfsImaUQCLiUGK0b7X4zL+hrjT2uNjMCKM7ye1lfj5wSLJ9N4qwThDTBkdOn/
k1FvkXmUOx8XeaqodRylmcEj0Zxb68O7SCpxBekl0L2c9yNdKARYXGGlnymMSRZc
+fZQsVTfzslNFVgEikzKm7djgnLiDSGVGILsNFk0QfiITWb3YC29/z7k4hRkt4Xu
e71AC0Whr17X5uRkJ/4n/qUk8tQagXqaLZI2vrLJVuCTk7F7OwIrNwoEjAdMGsbH
NRAdcYPpj/1Et22CkOsKwrDkRAQYN0wE+TDL+SzDfMFuB9Mvn7gKLgZUncx/EXE5
hcAknPM0ZnNSHgxsc0s43GNwqMbf/YRe4Qbe7Gue1M6IwljhM25rCKqqhOzmBNrT
pCeo5VJEmS5xGjjHhmVWhdbAtWNOtoLJ6D/mdpZ6PIMzX5JtOYZop/SoEtq8gMOD
hIPer5Jr1NVaI5X9aiZ2prBhezb4EEGj10DRKMhzdVNNz/kIzEccmDcE3kFt6j3b
+LrQrofCg6oPHHCaR7kiqKsb1EX4ZaaLIYa6vN/vkbG1aiG2jDFDFl2Dz721jAQv
nF2RbrmK0U4dGryReKtpUJ8mqyxhfj5NzcvPaR+jxic6aw0tjxQUxNC8SV07uykO
ZdbWX6/Ed0SO1t/TjJoMHMnAqx82fr3IfE0LHrAI9Vhm+gVC/Y9robFbJMVGM63U
0vciKyO2JwcPS2KDw1M1b2Qitf24FuTvj3B9jzt/JpKxva1fo5u8b95sHljJSQ/j
MamdU8IiantoM+jNO03Uzw2po1PoacybK4f3HGrRkicPsin0q/q85xwdP6HG/mcU
KWAMZmr9ksDKEvegCnIFBWtkhmucT2f/LGkYDSes5ELgLBozBXoo5kYkj3LGoFWb
yOKfgrwKnokaHq963lQDyLGep/bOL05JmWFMBZ+P8ojhfWJrxCcVp2iQMktT7Uyl
zb+rCjOpfFiP5WVrPF1HzKvR9J7nJOA58JaEvEbrVBsF67rqRveLW6b7jVm/NhTH
CpjfdKadpjYcYXMS5aQoQSD1Mczk6ZljPl6XlaB7xgbf7NTuRJoRMxnPS5HSeAeR
oBKluqFK1mIZTfhpD3BLIinIjw8HZv49cyt3O+4aQZYL95ruCzXRpkC1wbjKfp7a
GIqrYG8AKGSbpbSPZfVCfFV1zDCnoHSDa73YbVQox8BA5vV7T2N2yDXIgV8x+nop
VMjNvvNNHyDJIyQX4nYWWfPpu8cfga3f/L3J42fSTzhNORM2kKkrlY+HexFImgxy
j6/zlIkhJUSiij0fHSRDZ9yvGSr5/Ck9GRQBgcLiVFRdfxPq+T5si6Wmwg3E6JkX
n3jqDS3rlwiHDeerpThaXvYEVVBHTckY/w7OrzoIO694y6fxK5Z1o+MUPfxq5EmB
UvbFcJrJxv9qFy64xtEViKvFiKag/yGVBUYrY7Go2QKlYG/5DM4zvOpzfjBqnG7X
EbimO8qtyyBwh9LpRqMXVO/WrBkvtyqmLgCDJTdj9dglTeTrlYEoY5GED4VcaGvc
EwApCA+jzeN4AFV3JF2VIi+f8ORrbD1K89wBUfy612AVd2Klh42oVLHNOBf0BDLV
D4CDIZZ95B6XO7pgjL5Mz+DzrzvPskzlFpR2h7q7pWBni/y9hZghxBh2pF0+DfRv
OqLIeRhH/wqNTVGJtDVB7Ci9oMdBkKfn2vdF+4blP4Cl/2hbPHusxtlIOQSNs4n1
kK98JpKc9x/WCjHm6GBy5zXtsUcObtlfa6qVp7IfBHkpgxeGo8sPGIDsn8jUN/Iw
9ZDbgoGoovcaNvSg9itHiRTQqX1QUmO/PphD+uEffwC4AHnSBglcejlrBWM5pCdf
zfkWGV76Em8WahQ2qOIyrapUuZ6iYwF0/1qKcNBEgdqXow8oT+rY48kqQpLv0WhN
iRGaoTxB6n5GwRRNGzK8fReibwhgo61XR+RFNW8BpESNvrT2GdiLpZEJVaW8Ep3d
TWICAEesK8mMwVRv1YB/BkCGndApSiC4+srTAjaQcTPlgpQlDJSbboSbELUhNYIk
RdJ7nWibg8G3j4rgJdF7ywDZVkqSdAdHXtrmlOJLaekGehHgVU8G7kScH9p86T3v
j+3zEbuSZ4SODnug+KDRCTfZ9IyLcGklpVqjo1kIMCmHdJO6+s80tFpGAWaQWjX1
aR4SrhKTh0OTP4hyJATWXYSFqRpAOnEn27mtUHFZfl4/yYRCPVJbb7InejDCphkL
Cvl1vLTQ9V3Cr2buex3tnXRXfDS2RWMDVb9/jWjUi0NRPMAynURDuNJ1tJZ83Rrl
9od1DODpFnRbTgoflAnYAYZPYFrMApGOGiFr5DuvTceGArRJKMLrGsYIKziP/ee1
y2OiMOQcOX8k3TH61lmn4tKZ5Pm5TkiqJmKxcSjGAWZZ1HW+7sR3VNozzmY27EcU
fC9xbyY8kGvAEcMgDI1bv8nFzdmbmYAusuuZ1kOXs2+/z9KdiPBkR6GN73Boql3M
ah+gB7WodUf8xkKv6+y/yUn4xXC23LKMrFmlKg7ams1CA7vcKKexQ/EO/PdjsN7g
4avq6P1TmntRnyDfAMwLdL7/xhzdt4BHaYwgLy2a8l+UVA95jeXAc/cU14HZSi2X
LbeB/LeU+Hbwdd2i7tBhxSIezU8oY3Kh+MudrzgfGRBu18hBQ05zxFpCkMO59S/5
q8uOBbRZTqbdqLnqpdFdtxPHN53tfwtwSAtPp6hrfrSof3HXJAacliY7bxhhsv0u
TDXhotQE42nAeCBkxLK8fJbYbVIw1qjhT1UeKbmOdRUI5AJO289E5+4pujqvQZlU
1RniA78TYhICcXEv9zc8dsDB8tyLL5GGGaD8wrUpwwwKfeDmRSeqPA/cSjNbxra6
Ix2sgqxaYS/64xawuNGTPbC0rZOl/qv+yW7FH+V/+RtM+0mW9J2hplDwnNtfsoKu
0wX9e4YCFf9r2vBCTdko6dEw1ypGS9OsgXImTPIEy7YsALRwSrPEuwgLLEMWFq1i
aOtOSH2gH8MB+v2HxcHelyH1CU+uOoGPwL8sByY6JiZl2d2qxu87OtDZc8X9ukNT
Px2umagCZmeITBnYuy3+qjXT2esPdJUfT4aZaIuKBDiBZMloybKa3FMJC/guLTkj
ARQOSABbfOcdV/d4f2bTyMgSybTIuTBh9jum0U+WttWpx5Ed0r+npVyq79+Ku2xY
stYTIpL644nfr7ZLLO6jd7urlIKUG+sWFrN3JJEovEoGwGXhJwGl1iLp4ZTpIn1a
ForgBSpVzkDjVYL729s4nElU/J/kpholsAQJKTrXohj83cBs1IWPNchNiCXrem80
NE1/82IWncGwZu2+SNf2NBzdOltIjA4ycSF52NSHI7zjO3nVyyLqkTw+JgHq0jTt
3JHysepRo9gNjmUjNNEMIqfRyG0DblgZis4r5bLirP+9E9v1LxShUjhyytkZxOJJ
e3azG+Ln0SNXwcVEdTmw9SHKA7fneLtRZ+EtBYRrwiwcF9tnC694oZ8MZqzC6Okl
y4CuD7fjsUy46AMKGEZZVcTGf3ryIOKEg6zcsnIz55PNjPHy1VlcOwSvxVIow44w
0fh9j7FtIzAB/Co+/C9VC3wvLsCdJe2t4oZHCt2CIgpD2OFsEbWQUGWdDYl0jx/P
mjus9ZChcB4OfU4dVBXfEhN5kOGFZf9yNJEvyp3PgvkuZs+O/PzB4t1wt/DCjlKj
ZL6lYcyR4kP5ZRl+NmgSIbp4ZJe0uSd4IP6npZSYsxVPBamTqxoZSyg/RIAlkzIO
DW5dT6fjgu9CooKKtv0SOwWvZgGxNc/TwTUgbH01cy0VWR2+o1uNFClBFNnkHIsG
cd+3UKOAtcBvkFpSUzENsddm8OLToiKJNLSilqg2ufP2TYB1dsRxpU8/Vh30Iikw
xyPXtmtckGHNYJF3kQKnsnb+gDE4qz4/Is3+nVdgN7BjUMgRbAoNT1RNgyr8ljyF
tr7FWhai01nWHVWKrUJ5iwozK1Jw61xisxKSJEpMChKCM6Qzu40hXKSC/a25NB/V
kuTblzdnVzfgYUdNFqPGXPkilRKZkkXVMpfaLAjZWsllHRM8f3PNPVNJBJmyLmHH
uzwSC4JNWeKEqomkqAWjrU9PWmrDBNBcY1+3zr8Va5r+TMbq3fLaqU0Rx/8c7QES
O3oc9V9Ean89lEikrVQ+ukFPwEfoqhgjflhHwGMpc9FEvzAi8vZrAfRqc1faEBwF
gTxxhzH9M0mUtnR+qgBg1ruHdZbCGTlwYmyg8frTmzj4SdOE9HGUAB/vh+q3Kwic
EkRWJM27BRxUQ3ql5etXV7fldTZLodzPT/TyK7gT3HGZqF9AN0TABnpZwQsrIFUc
5ZeHCdLR2P/4OSoC+ADb/kA67XqOKi5B0vMg/c7JxyMBjlDoT/dlDcHItCd/Ziwk
/cW20pMRj0o2Ptp5JtYDKGqurbCoUx7byzK7AS2AaW+Rev4PoLTeIJ8ZvFzTVE8O
c+gmWClqnTFamUWJ7M3BEWJQawqntPapxeFdv5iqOJq6tj+A5VfS1AwokVPH/dr5
6vzri/0BWUJf4bX54CHfodP/1KjlY8Xky60OUdH00WYn8yyPmCyL3CZ+lO0A+wEG
KTYACgEbG+lle3ZdJVPNDtAnYeJgEr/c/2n3ioraq/GE4IhqSkLSf8M217vVr5Wt
3PsU11XVvaipui4EHjQv9iowsLudkNik15PNWTDsMlJY+JRjuXyTFcegje+zt5lN
FW47vyWDZjSGIKH/huMjVHu9xHMIjT8cxS2z1UhTpwap3L1PzAdyYsjMISeMI4oP
PVI/yGKPn1+YArWYQekYZIWJxlBYZoUP7P1+WFyM5SBAu0eHyAWyA75wAul2Lvta
UbbYNmvsDmocWP3e9KduO74cXH3Nh48tIipV2rfrPRoTP/tO0DAQK13Jw0JOM6qe
w0lcC8JhC6iXexBpDzM9/DN+9zamUuGBGQgKj/Gd/9banBMciO3aizJXOjyHAcx3
NwGb9eruS1RuT2RYj8iOd0G9FTeLKfUuoylnkwqbAJpKEnMFO/+GUWnoUVqtXZ2u
TiyhzFa0LW0n+jhwGr7NydQ/DRk9HE3t4tIJ2U/JqzFX81arwJXTeLl1Mxf+2+/L
A5tPFcKMzPWxd5hd+LqoLVC5c82W5x3GLDd+6vdJ9WAJwcbzeBngZjzLTZIqm5rx
4pEdFIPkSUKJdwlTKvisc6SuLkFWGJjvE8cT2KfLIoKlHIsUwsjaIIwq+EjvrdfN
4nk8LXWMbdVPSf1J6G+nMByR34wl3I88JrqVJYKL8Fij8gIumsL26USYslpSi0/a
oeyIm++6gQYyn1yYUHqeUqdmv41zHzC1O5WGq9HYvp9lwCD8av5eEOR6iGAa/Gws
cC6LL4TusMTlJlcE8x1siKkxPgPBfyv1CcZYQTlWAvH5JiSr5jw1S/H2im/eBSQm
pryRqs4wiVnEBi0cx8DaCLh9pZDVq8qYnj5IbaRR6qmYyCuWhRsAzv3JwCjArNhy
PBf9FsKgL3N5OHiZFQZvaW/gzYx1TLzOdHJzarH/wTotwu8kWBfcGTGxse0TYtGp
FyOy8KhEye8qmr60regAbEMu/TV92fVFWJp/Dj43xRsPYZTFga/FxvzXZc3OLJFL
WmaUZJox2vV/tuSpFhdVChrLbrqxnD1WOnZHSVmjGoa9h60Pg/v/C5bFd+G5zbW1
WUHb7vzMwzosI+JClj3IP4xyx8fScpZmnFjc19M7Ya5096oorXO01rz9PWdqvk/X
la5TCW5hNuMemJUWxX4dRY5Mc/YnAKxgOEWos0Owos5WFPRqEiS7Vgf2DCf9eV7F
nXSBI214mwIIi0x2sq2cxmOVI8hN/p/K8IldRfzdkpQHW97nnay4U/orFz26Lzhq
rYXreb7LXg0Wa908S7eTFYOGY8pxGqgwoSz5b3ekJYWrY4AUpTDgr9NAOmxbOm5d
DH23FE4gGq4EXMaXMKfGGq9a8UjQTa9qKaCrAH7dtI/gxyjspEYToXNATAdAWfg3
ZTKxPmaOpFvTXEXezEvHwRE6rvSmhkkVZcrP/zBkl0s5LGXc1aDMm8dR+w4Eskbj
EfIRxiwX0nYLbs2Odt0Mt1XanaOxwCU3LdrecbehIl2+Bh6y7ffpQcjm4wAVlrko
EBTxIWIXN8cRvHre0YBkrxEH/B9tATQNb4JcOjFCEYPVMDSHn7pzpCJbXYrG9Rr2
rpBkRMyYx08dX7YijzCFaYxO6O8Mm+/lIj7HlL4bVyQPmJWPctGwL2HjOYJBPSfA
+m0Phk09lLGTgpkiTYoKZZcCWFhTNnsQ57e7nwGNrM8KRtW8ncY5KX9W5I2qjq1U
qI4urBh/5zBYZX9BPzgZnjCOXcNH0D5Yx6xq19WA4d24xh9U+JGnS7RLrniM+Sjl
6T4EpiGUNYodcB+nZ47y3BtXhgLC+gWjmj8RGQ1qqaHEBMnS/TyoRlhhqfZBIJTf
DH43TgNwJj7q6zXKov/CTe1OgnTVAzNrCY4F2pN0uFZARrl8mwKg1SC/D7dHQjnc
Waf0zda1klcnZr/HilEf9h7iciO8uODmmw51kJYzmkjqnPpHD5pgX7BF2qxttbGK
XBDdLN4HtQ86dTJw4BDnIG8YC+J7K7pC6pYkxh81W/GUG8rfg3VSLG+uK4DJCZV6
uKXwH1mQeRxxsYUj+cOitpH9nFtYvEAjGrjqR6olG13Ktx2vVEHKQx13jLRufAld
gRHphiGvmZ4G09w8KcpFTTzaufsyR296yTXy1q52PCdHnbVU6UBRq9y9YHLeIyL7
bQox6Wt4/udgZh35+Onn4Sbqgl6j0Li/sUKwQsRWzAQS01rbhfqNRFfAsNqgFWn/
NI6+pYVj0P4X7x3ozYKCrSktZEhLoBs9YOxf4GyWlYzSOBHWhAUyyZMDKvE8J4HN
7XSp3FJ8R87QUenIf0HlBbPs7pOl2oGN7De6vG6bH5/0wK6fQXBwQLHmVkCH+c1D
vnMCvOgVGRKmTroFfUY5m/mhxxYagBAnIkaOuNiKKYHF/Kbk3jGjOcf8xHmM2/dF
0adpx7dxZg+rAnrc5H6aeD0ClpwK91Cbu0U6SueUi+KJFXpjM5jK40GPnSXm3hbn
XLQ/i8rNnrJvSZLFxNnPD/ORGXth13QxUXLAJpSp/7TuVJKcYWg40u+PN/Dt5Nzi
XXIiexcGeclvu0NmwZxyixsXF8cinj81ABlY5J8z8i0agbp9q0zcyNXvMgzM/Jwf
fKDkuj9irdP2h3a1QpMwZW3/eqxA8eX7rf7V8Qhu/bXpUTOKVS/iuWgv31xbJ7m2
6Gnwecfq3s587lXyh778aOMArxPz+GVyGnNPKDSVsKghokQVnRhAnj2L+sTNvr98
KG+rgVQDGhwhOkL9xi2xxlQzxd7rnROq7gThvLZk3ykLx0RA+Rx4C6QTDkaa8M+y
NEWNjKnLCBtQ6faujXGeAWO9Ga0u1B1T9a8cT3sz3d8WLkoMxefDP1b/bEw7hx1Q
mQbjOANGd+dFz3x5cFDc9ZiK8HpfOrluZtClz0unIjczptdLy0DoHlxvTkE0GvE+
tAua2XVQmGfW/6JQWENXeEhuMDNOnvPZOPmeahazxyDhOoWnI/4IY9R7EYVUMb8+
uY5hKbq7AotOPD7MK6Ru0K46C8Dq7PxxjhXt+qNxdtCoMOEGrZwBT6Nz2WchzHvW
HtV6GoL4Bl9XtJmS3K8sGf6T7EIdRXMbgv0rSseIFRu3vsf5fZbb29zvtf/IjEYv
UBRmtvU18OTAOq3zlYrr+V+9rG4gvpiKqkbcDX6/fjf6CxypphlOStsI/PX+NWi0
hnM3q52tQlCZ9lVfryalOfzPl7+q+y1735Ivh9qaDhzqk1XjMoGF5v98oRM5F8OF
fjDUDGmXf5OQjIIPOgn0N3JLZHFmFfJQzb5w45SoVXBAHRoGWi0fsN/lANCj95Ho
3AkrYmQCuIV35Ul6U3UOjV7wycMjczWnFyIOaKnH54kl6Cgusbug1/b5dJigb/h5
H/36ZJ7dy+B5ua98aiAPo3IYxViIKD8/UAxFpsWj59Zs9sGKxKUcEPxFXCUn8OtS
nqLsPXa6lAAbo3GCpJe5wasJ/HHxTJfkXgoC8Z91/PRAXvdiIXG3tT97WJefUsMY
L3U+Xo72NnT+3uGhh2oNaYkQ8sJkVcrtxXkJ2P91lBS8qF/n9gbma4Jy5rh+fDQ/
bqBGv8vjnwQwp0z19t6qfX3hEdnTtIqeobYzUIJaoCmKrS99VwvgpdLgUZES0Bp+
cpRybqVKZ5ic31E+D+spi8ePMOrIrw570W7I8WwUYO6nL+LvvvoIOIDcUoW2HlfR
XdffCb2AEi9aX6FTIWnkj+dhCB0ndE7K2qXk01RZbSZxGC+3RUOcDfzYDZkFcISQ
Sltg9vFUxNtxt5QIDECkPQ4+JKGi8zte/sZq6CHLcbXNhbSONJqle8qap030uZW4
6WonxhtGqQ4qxmO/4V0TPcF0TWBQpHBwugkPmN+Z8LjaQMYkmzDEsbRJUXB5FCK8
r8PxJhLsu9sM/soQo4/QvmXeZ4XL3/8Iqrmuc/v7EqEjtoDiGK/2UsacyXWWf2gQ
upbR8XmJ23757Q/LmVMwRWQXPVvA7XAhnGcq4Mxaooz5GY0f9ExkX3hZu0ZnQBhd
a3pkjVSzQUgJlWtWzp6LQNZPFNO4K/yBS/Zb8Y/0zKhdejNAyJ/k6sZSWpG5tkZH
W5m9dju/n4J12qC/OoqFks6gshoPw8xzWcnN+SNp2h5jnUU3TZId+x/x/J1NuFEJ
E+CCJRbzENqDNE5XgR/diObG6eNqSf0wA+P2zpNe/aBlEPda+0MoqjXAsExbWkqn
20JmDqBfvcqiu5RyIlYQ5xzOaF+cV4MRiGlerXw3UMhw5ZX50K7YFAFGw0hg2GDT
d0kZXb8CyoCNDQjRwuNoUL5ZKlgWTBo7AD6pDIK913zSXEhjx47mR3J1lWo2qixE
eGGxwMPco/J0YWauCoWWw7dbqerlSsXLajD3k+VfhiivxwfvO+vnspo37sR26qG0
hnSPdF6JhlVYVuT37aLrSuHcKExtwEI9nFiTQO+C7A88ETzA9V1D0LzhLDb7TEaY
xX62gdK8EM/5QqvzTHe7tREND5y5BSl5lyr/5JUcrNbS+fjkLXDPGpFM8v6v6YSH
ReO1J4wedMHVbzVfaCLpUJkNDVcpNlPq3nZ0wIArXksPfD7Q0bEya939jfGgI8vK
/6EkR4J4S8eU7mghilG5D8ntRh3AGpamQIGU+IY5DpENSEhvijjIin7QAfzaY/8+
frnAodavSzVeOfPsrfY4Gq1wSF8dQLQnLDIraZJKro/pBJ4itZbxTn+euRWlehRH
CzZc6kUjGJDYZrp82KDbuqO4L0OS+0R6/rAcjoFPACMhDyHsoOlWAioE2kU814YG
dMUu+F1NRnmPW5cdHgSiLsJkS9opN0L7CESVN8n3KhVirEL7SbCCRbhb1JeZw9ln
fjP1/AVfgM4gID3gEyAFWdS3j+uiO8bcb72/Ky6kP0rPRJn6DMJtFm+tIWRIP9FR
VYDG5bO9XWa3mDsXxQY8aEfeup6sckqwt8uuFM647HULySfDPNdp4oi9YzB+D7V+
1wEPpnfKnlliRi/OBXlN8wmJoTyUozLJhKYqeie8c5RyTt4MtdGo9sRHzwFbSUlc
jOb7fboaGFZXST/go02q/ajMgAciLaYdMQ5ln35uj9AOBW0ZxT8AyEw8YD1caq0L
kHXzbtZxKNqz9lpSes/NtQAn6BnBCg6tLa4x1eBnjSsa+p8xzvDqE+0EJOOGdvIL
8C4upqGwNCoHWokDaeZ4Uk4d5W/1EPmP8yGWM/sBrD2p0MBjhI2/M0RNCUZvDDzn
PSlsRV7/SfYNV+pHowZGVQ5A9HRQ3d7Gq17AUoXyruFf5fmal/tLUY7UTmVTirN8
3kW4ZrijowFtReOAIiH0iA8hkreEwqa1kSTVDfAIrllmy46eW0JCWicJ8GYF+7eZ
KZcf4gmnAoHpsLpbKglefFKmrvjnPXaZwuQp3XgPOOJ1hDjwCcoQrFBqXxge+FEi
O3iG+4uKUen2wGeSrg7NGUQlsE5mb+HzO8WDZfX/n5LZj/DHnw+J7EBbUf4ukPXZ
e9f8LpQA6AI3hoEuiHxyH6Fv4OqpdEkly/QgByPPkremQTRWCCHxU78jq+TyR/W7
8Gu1XNArgU1jOD3TD1jfcQnwwgrRIt0uT7YoZK1myoM7qbCZYii/mGAQq1ASjBuQ
5KfRuTyco2dl52nHqOmzdOC1hLxZh4DH50bOStTaLbozgzCV/M+hwD05Lg5jE5yD
DLRMdZ6XHAWI+ECa4KrAggM7BjcQU8nqV7gotBPGCHdc9OJz9rJxyCp07PWx9vNC
fKTPB0NqMvSz27UopaGhyasCGQjP0nf+LYAdraIBf2/JcdE1fqkCcQ4haKlsB3Ea
5DYke8ZdyN7NUwmQqaqjlDKeruT7xGpB+bF++ZZMw136trGgc1FsSBuGB1ANtfPf
Qg4NvSJFAqKwKU51C+qGxNUUzjyOnTX3e5onIeBMJS7fJsYJooQxl/mfpgL+4iTv
I4ukDWtZ53/gcIAA88TIy4PvMXhnI60IPOVOlFFvexc2IXMa1cth7C6vEtrnQQqY
QCB1aoOa1sLeXxEw0ErKNmzZDjkFKo+IcATF05+1557z/nzlYT4WPWO7eAB0d+MJ
eWVM67MMPDGZNPs6pyS40TzUCtuM4boUqiRdhTlWxpW4+IUJn0QOiP7erdJna5r5
Z4jDYFyAiU4cdA+9hvzp5Oa/FNUno8D6y+4NSpag1Z6D5v1rVqkTtwwArInwkvml
8kJBhAUlH0xRRgM4yXAsLac8ohW9iPIjA7tiKjpHFkoSPaL3imGE7IYFBllqeuyp
6FbIy8SPiY4p37Mb8Nu+ksZXUDyapuJl0+HmSusyLsmwd40uPrGjgyma9Z1bLGBb
sOECaOgL8xDb2oJaJ2RYLSPuNRlN+mjEINod380QfWkjwHSVmyNiX/7cjFsHHRbG
L4uf3BveFRv8gjC+SoJ9Emu0t8tlfGKnKo/RUczTYqoIhKq17cjIVgFsSMUr5EIg
hIlIUS2CoMmFt6egLSulM7AiZu4O3ASHumWNuwZugh8FhuBu0o2JfpIDzHaOQeH+
uRC8jzzwuUEsdQFYn4yI+LRvkVTOVIE9/1JTdzS/5odETVbu3t/lemaVT+1CBqoo
b/RyRv4bx9OiHeMzwZQM91T0wubC8XXZTmulbHmVmUE3juDUUMfMMBs7rRHET1Kl
mNGIyXaVdCCPbxtMzvRY7jAtfy+vlfF9uAOHxT7eA/Xxl2TE1+garT4RfxeckfoR
G+VnvfKxad49t6XEK/RqPBY7IpthjB4wrBxrDnjyxwz1Hy4sqIQhCaO9ZbDuSMTo
JvQhiNi6IWs0c5kI8K71X5xaibqyyKmLz7SvltxJibkLgTZL6nN2UE62EiWrSuq9
KkSJncrG2dRGXTtla7QTYbShfP9kKurLagMiN4PtuU7TWKA0afxAAuYsfH4lscFh
iZN5H9yBxRlfj95PUa745Bztx3G6ucMDpdTCOp3Tmv4vrD0VeHzMvNxqJC39rQk1
ayj1eFNerU4Wg7Ho8K0P204ASkyhu86ms21Jvt/54hP/y54RHKEskRJHjHJkLhyw
TYXcvT1Fu033z4amyzKMQL1BR8Jomj7LJToYLYjqBKOahRtg1w92zWhjJUOak79C
5RV9Vj37wo581VambmmaZ14K8fJ3rmC7mIkB1hFO2/cd94Z6475+d+x4NkuEpZLN
n9XZPvjhnsbfBo18+qCyBA/GCWf8vOdHXtiPTphoAYmM5y0RDF7f9AjGYmEPX+sz
cWkZ3GbrRrr/ukmN7S4tdAceefdhEMJDwfElC7zx4bkQ3RIvlqyqEIUHN/YgoGRj
3FLlbXyAs4yeWd4t35b4WYaXn6G6xYNnww9h0Z7nRRnahZv+SK5XCkkyZ/P7O4Ml
eGdxWUJfGKDYormt50eLtUHx3uW6k3K455C2DmL9NWZG2Vkd4GQjzshLQSY4Q9NX
lTFtohYtcRXJjMJIeNYZgdfbB4NLVoLQ1H6Fszb1PNwHoMsTNnEjA6DNy2hFX3Q9
on6DwAOAGOjiTUIbrTxi07fTXRTpFdWIYa/jI9vukiFY2+e7CHIT3HXoRYiRAHEl
Pb15aqy3FfKMlDmy979eXDsZ8lELugwd5ifGVLTCSCbXFhOiZtCKan+LPsJME943
47tLSPkZ+Bu8/vW5I8en/qp2h98UA8266nqp3hI+G+3ENkeb/n+gnisRyJzPM2IU
XKV4Y/vLTL7hnbaG9LqCUIxWAg2rQmUb6fuLOnryuxMAOsxV2lsnCmBWdLpyyJ/q
xd7VsnJUvMt1GqZbvhZA7ID1E5hAYoXM/WZjJbBKr5tp3rYtrsQ8kx0AGRaAVP+S
UpqV2a4hbXtydhb3lTcc8NukV9XepCKtw1fmCKgWuM7nGmrlUKoW/1xFcUbXRkZb
LrTtyoN8DQ2hrwZgbWQZ/yyke1bUpbBttRtNwRqH+R42ETy3hm44EvoZYCooCu5r
78E/njfL5OwhrGZOirKCxoilPmF07DfTukOBjIUgPqckAKOazSioadOxD54BBYbj
Mj9hWBBUVbL7h6nu+4qTuIJ4qm+8J2UmxKaYszYoq8WrgZJxOUPc7lvYpBqWyTxA
cpy9quB1s9Dw5P6V70nfPOgBwDgCBaESZ/mjend07h/e3AQ7YHeEiywYiug4f9GV
r79vAGGYDBGqn6jo2yVuF7wLYJuhODJf1sVXI+G927FpnOgDmMzTP+aaH81tDXfW
a8dw97edDvXHzISXREHDtfDPVKSJXvQwUmtxmHggIMI3NbSyxtlVerXcAB8jvGbf
ONutVcSBcOQFq3PQMiEJg1K9o6BHCGKWf7nw7hxPgWB7alenCbrNyNTXH2TN5uWs
9icC8eycwXdIjvKqdltsUzOFHalThZUCY1CCAAMhUpD10MihCk14PLfEd9d2yZFK
D4YNJG6bYX33H1HZ5Fr0H1hawk0SEmJCddcLGMJbDEvngRH8j56BPYgO3fBbvKTW
WTrS4noBImey9nQ695dw6uVf+IRURcpr5nEkO9UseAhXwqGmB3+MCdGIQRAk6wd0
nAToGAu8blZhpDuow6pvoFsqJEaILQLz56o+oiFEQC2L5Rpq3KKAIRUnniwT50PE
Cdr5R3wpHqb1eHmXGiT+TqwRi4Gant7+QRQGxp9VqjnVRWpiivNDWmf8T1bnnypR
lxpjKIXkkQi14V4+YJlCWwoqdGyVV2Kq5kf+sFGw1KMP5xAPbyOjI0FRo0qX1bmF
8LY9yWFFvlteO4nIGP1Ol3lRbbgttcV1uJRBNeLN3S+XMgqNSmLSNTvusqAXCyTI
4czi0pDGrAJCHl8B3bzPX+nIf0YRIhnSSk197eSk+HboHiVW9kbh6yBfOAeJpoDy
HFJ8oHF4q3Z9wOg2CMOdPKsiNoSY7/dJ6GsXiPAEcpgjAY5lxqINYZPyyci0UfCy
gqeujqm/oCKszSZiPrxzeHdBCbCDhysxTiV3Rjiv64nuiEdbLuxaFDy0mpdHTnbR
13/AIpXQ/US7W0ZqzhX5I3w6ztSn0wrRccGMPg5BN16sFLIN18bxl36mdRADOLXP
6s4nuDy93D+TZnK56cXYxkBsuDMD6P7HXxBkok/fnKwk3Sgxdtxqgcy3qiR8I9n6
GM+XARP7vneEIkXKGCXG0BP7uWGBGr63y4XPQ6fAr68kEMeV1/uQYsI/GtfMFwGq
WFQv/OR9SJHvyn1WQz3QX7hpHblhKWXPvWVbIhgW42K7G4C0RYGRq8FhVswWSVvw
b0ESGC9sP7nsnQIaHiHbLpsuce83LhHKZ/RsFDbACfHIFcUDj+zlFqVX3RzZl15L
Xv3E3K4q9GEr6A+blCayjOVgpv2dErkOJB/aUYcKDg6P/qcqKvFj53gz4/ZFsT7z
14UlrYSRdkXhkIAXL5CH9S/cfOn7sfDatzWNwQioRca29qC04ifO4B+OFDkRDfU5
bwY6DqARU2soY3DzOAbR0NjqiOnBjSY35+YyYG0snqA4sMexxRBitdKbFcLHbgpv
It1OB5GkrAJxpy+4KWjUawjKUGZc4R55TIMIS9YssjbkIabz5W3U2l7iuzU3tYDm
3XoxL94owSV/iNdWuIUgQ7fwyiy8/5Tg2/CTZ7TPUip0Na87zdj4l3f4cTb+LRbf
JqdCHQxF2VTHVTPSYExPvDRciTn7HgH3A1kmrPY/X6DzDEDnSc5hbxugRK48luCG
H7eHLnXBDZdKV9sh4b2vsK4oKYJQw/W4Qb5ffZB06uFGQVExYm2obtDwMEWzHCqJ
DnRYBfEJAj3/beVAafdN2kZQEJdO/K5174OL3tkb96XskayS09rAKW47nojLXW5q
42hBz2Ou0+qFI5+g4f0AGrXptm9WDfFRmU6gVcXAzjh+TcTtX56sW5FUv2pe6xIt
iuWVIlyTfGyzR408TcIFklIifBkYdxyTesyWy60wlLuqUWgNR27+35Yzj69BnTwy
sltVyDXi4G//CJgKbqZHgxKgqf9iq8zZnvRYepHLHbljV6u7qgQhMvCEF5Kdi2mD
JHxMi4M2FHg6JIOo6MjiMsR9x4a0TsjTNCS2dV+XkN9KUnOwby+6tH4O754jFgfN
U8dqxN7Yl0ZSrltju/ipOF0CfW3H7wbvCmE8JvYoHw+exJuB1/Ajv+bDN01gZgwU
C8nV9EyLuileuMEMDGAbHydo1up09yH2syERYMlbtR2FyPUCc7rgPHyMhshXt/Fl
vvuSTMMNRdDN3kyVUtdXeqj288i/ptrjT6InvOTxFaV+ffpIWeFXTfUb5tAL4oJg
9fgAzMyuJigWf0F+pE/7RsOvksJFUqnlCt5mw/S4M/WPmCE2rO+gYFliH7TbyxpP
FjPddigTGhG0bQt1j+O7H+g0yXJBUOwmLP8s7qtVrALxoZb53d/U/4vIVvVeiyso
VD68vnpP3czm2IJtebyB9Y2Dg8vf4D7aBMpYsOEvOt103SXFZgFMefKM//Zr/pvL
Vx3VE+VRyOcMbJKfOJi5D9FhFALixFjV5T/ThCw9cgnpCd4MKsVCUgKTt0CfJf/X
JiZ+ui14CTjzXoXYU9HkfNvak5ANIi5YN15xUJGpXv857mpbdIIreJPC+YUT2lbG
BJ2brJn5857rep38DFZyTgQuuM7lP5LcGs7Dbuk/vDIt8Uj20fpUuXmsGQW3Nnqw
uOXxoCUiPcKJ282iogVwU8GROYr6GSEH2aQQtuehKTqk3+0woaVlKtxp6+560wBW
qPdEvO/9GJdYlhNxP8iPbIXXu3KqWsYnXX4Zm93eg2Dt+pfCxLVmqaEn7YuM6UW/
9CZZso/49h9B3nu9iyxj04eT3SIjlPj7pnnfnOQ1x+dKtWrollLn0ppwgvAq9PEI
Oktmmum6TS2jhN/WMUVzRLIOaPtgLKRa/wNrni/UEA7uhjxWVYqq2MJiEGcMEhVC
dPaOSeffIdK8B3wYEnKPfw4f2HxV1a1LakyGFd46MzEbcDyhGPhWFqVufhteq/hx
Cq5Y3pMKH0b13uM50gI52dbIWhjffqcR5Y9siaBK6ULISBas/XEBRj2f8jQrITUh
bl8kv2KyAKoJo/pKH/OwurwW0iGeEl+q1iDkGcg9OOfuCwHD9mzP7u4DDlw1smc5
Tm7ss29D5n/kFXC0yz4A972EaXo+LBBJ/Npa3J+WcPQIYPkVLd+XTfgkmNw8QIZj
t6tDfrwkQ8E61PqrBUxn343/8M32d6NvxMxTnfUjLi7GYfykGYt/CAV4S+Ye8Wjr
pj+CKrHNWE62muw8rW95bR0Kkq97wbkq/Muq2HDgi3tP8OCLS7huPhK4LBCqjzou
bf5D6zjmcORJWKns9WCwRpXEj9JVHzhjPVhQyYCVl6jUYdb4rjW1WFCsEAE+Jynb
DNj997FZ9OUHTtM8Xr1nYJg0tp1PTtWzozDJOG/vTBWbaeVtI7ZLhP7wgkiytXc+
PTiQ4QVYi7pmxlmQiGYhC71cUGAMeY8IgFV9gZJzzpgH7sqkAI7cupFBtHVuFZdb
JXmQgWQXf/cWi0PzZB/IBLvCuh+I9N/hbvIR0cTDuGs0ZpwE1eOpS//pFjMs1ETb
JgJYnkPSSE6cLwN7RxKZ+VxEWVQe+jdCA1r9tWTqK5K7IxBxdfaxmHYNSkoGFx0x
rEUf4UEKu2gTLSVO4VOSG2PEI3hJAOkukn3vlRV90n8nrlB3VKyEfK7QhALdzd9P
VRh4Bu62aum7EM51EEILjLZ8qqrRQixLXN98Atlz3UjuohBdhP+Zub2GMgYF3Lo7
UKp3Q0qYlfrGxNMLbw6LdAP38iIVtuKd/Oxme/8uMHyLjONNtiAUD/avOBiJFM7K
kzd5m33spzaLKpBTPlKKwqdLHjVYnTd48s9+Ec0A7ky4kXwQM5WJpP5PSUWSdYsi
XzWd33kb+6IMxR9jxV/miei2CTQlLyTiGkEq3vNaeba/xArVwgz1hw9FoyKwp2vI
5hxDQCIOuEADX6YmxzRAtKT2SEevhQfTJ9e+zfl/TPA58YIQhAaOfrJ2MKsRxHPi
spoax4BIbhQd4Qn2xnnQlZ+q5NUr3NKjLOErVyvaMu9seg2H0nI4vCBQk6FBA1TS
Sh4gUswPnaMAIXwe3vMGP+iaDtg7xBub0G4XzxEMSLcJ8CjSJcOfTSUCsIjGbuZD
SIpTgoZ4/+Yh3ONTeEKWdZi4ve7MH0CKGkqQtnIVcjfor+9aoGV4pbzT+cM0ZZhu
uGUzh0Xc+XsgWIr1VHCDGrOJGKGEB2p+WguRUtLwX/39Xu9Ozp/vUl2jQpYsMyho
n2DONwvprReqwngKdxlv470lrHCEnT6s42xUKvXq4SUcHswxwJAACqtvP1ezJyEU
c4lBrDtL8IJ8SRWNm/gp1hUWz4DhYF78roRca2GgkefbsDQIIwqW141b+gPXDLke
WN6/lFQL6RHFHE4s4ek5p/+HYtRtY1ATcyfpG7CZWvWlpccm30Z5josnZE32+c8B
E+yoe8v0haKqzokZMBryyVkkZkV8wwsuErqwHEUmMbeEBDCYb3tVqdUsqmU7zgOy
JuEunlt7eNDguL5dEDewc//miqya+oKQshAyyYf4K/fZzIiSIF/jGW99wjkb1PR4
p00teEGJffacgEqBsVNTP+BwXmUP/jfol+RMDnFvasI0N761W6ccsGFGFwdMNHso
lJ7zBciqWtGZNwqsz5PyQ0miIBNS/8zvVOD/eUBjfvEOmh8WN/GpQfuUvLuGJLBT
4Z+lAXBSv4ZmEE9MwyWPiaDF8m9PFEVdNErniSRNKhfvo2xvgUX5wA0MieKjILbG
bYYmzqmK8Y5XpSxgU2NOcoVfCJjpmfA3MlkJhxWHsMTUD/QqJv22qpyalLQjhr8U
srEWKbCamnFcZiPBCGS3gg5lmBDnQfYlYc1xkNDNqylpb2Hv5bIfJY/V6bEpFLuQ
nr5+d0t0PND9wjTTF+d5zwUCbXEC6/T3jgYiTgLHDSibCrvwobdFzcSOfZBQWDsC
67mqRnqv0sS9LMjsERfus2jnwWlLL7XT8iEzGhe/B540oYMR/sD/TOZNi/7qyb9f
QALEDM5oryN7BonatMsZstEBpDEdynZEmMC2bZ5eSW16ZRWTDQZ0M5WxnFEKrNRu
pkW43SWcLkaYcCkBReYzHfD7p7ivfd5GTkqEQzUy8PnHUvAF3l4eIrtzIC8SY/tr
yog5n5DSfGw5VIKvKTpGfR+Yk4ODz8tPZeQ61uf3ZVoLNCf+cmoYTS+RHdcM8KW9
4CIu3BLCXeSqpOiKtluzZlZBnhCdfbO/o+VrCD5UFHbRdPznTV5TjdaS0/I6OntB
ZBkrsmWxP8Eutxtp+59AMKeq59oOSLqCgefmvdcOley4MCDa+Vo70+1+Q55vtrCq
s7Fz+8Y0tIDBuHbNylB8U0zFIq+XEwJbWgEROsA8+m6dLNKzN7bS6sMGXB+6cFpI
5TXoblKk4fl2npMGbaJmyKWjon5uq3zGKbTEsw612L/YPhxig6pP+ir7UnEh5XWk
4qoumyx6A0n5SRqTCCoiOopqeK8SWc0bMPgaz29tnshb+kN/8Hxc4AEZ5h8KNU8A
89d3aakZtWczjCCxmdLYYRXp7bzh6y+NCTW5fHBMa2+6tQrAcrVZFHGIUqCWM6M/
E899g29bMFddExR3EYDpOUezdhTBdPUyLGJLHMrZG2obbXxF+LrcsOAas4q3Xugu
yP6X/CuUmo6HpdzaF23LDx7kdGA+wpC9pbWbJaRt/mz8pFzAN6kDG1W+KsgtkHjG
OSaG1mi75InDuhv/GwDmSnN6EDYuSXx6sAtZNYFWRVmgwa/Omm9BbTCmv4oD5MKY
LVphFr7POc7WmsEKHJQJ6zyoNBlHRxgl6fEQLk8DH/Dq4SNcXmlFhGw65+LsjF5T
OJMYAz6E359SnWXGZvLsk4JTSFP3Fjm936ExHLgKXAeF4HS2lYN3s1eir5RLgx/S
EZQZnpfrNurNmOt0eqE1KdNYyW9Kgrya8mF+m1vmUvHTnX0+suQydnovkTnGkSWy
CCmPIoxhCaTvHNrZfcnPH84bB6pVd6/fWHGTT7TszFhkX46371MHN0J2tW9BESBs
80nRNHMDLHfR71EAUy/9q0BRguR5hWH7GnjM3Q3VHJYcEHjXTfQdpC3JLFCRsPAf
yt2yrs2utxl8Rrl5YRZbQmFwtiD9mVaWXTGHGL8YCtTubsNlzitT1ZiFggydaC9B
F1S+HvHSFXjIzI0hWC0arSVG/Apo4ZnV+AWMJkO/7kJDPxdFlh7vXeIjPifchBTc
jFqWu9H6EsNGobpAUIZ/ZoGaCcVu8+A4MGLDWRICuIAgGvhFejYPkNRKzMVhgr5z
4pMVZQsdoh+KduvpXYxqAQr2EWHmyEqPN6ACdJhyfwajg71LOd7Cx5xjAUJZAHQY
hLQ2w3J7FsjX6VK+3nIfIQXgUSzcDzzFAxQl9uSvYYQKsayNpBbQS7t9Htzk6a3P
4wJU0TDaGFgG3Fpy7MkY5s4OS4BRRMXvZ1WFhG+kCp3SVUJS4YUFjrmzycGiPXPj
0P4HXVAdMKEziZVBcclfAbZGScTWKo2EJc2YqApTBx5Otkofe2ziwsDVK7J9JYZ8
rlD9OAECqvpVt5pBHhI3E4bjh1kO66L5ALbHvme9rdxHfNXOsEpl2Al0GAq6bXM8
xPgdV4eXC1rvfotBxPWOCXGVx3HIPQLJxjG0ywbcz0AXMh0v+a93rSIx4As5wBFS
3n+GM1MCAzI+ADueCWTIHTOY0ICszl1SQs1gSbE1WGZ5c4FLABUL6EVzgRl15Fbh
dq0Q+4WERfUstrWhKZOGfV8UGE0SKIYwJauNi7zqOESBaSKeG4vvS7anuN6ZqamF
/IQv6zXjy16NFX+Rypu5KhoyeZfqCQSTE/eULj0Q4Flql9iLRKWbVZXRj15VhNaZ
YUBt0NbDYLKXwW1GVOoIeGUlrtMlMaPWGuwN5msZjZG7B15S1E5pQsguGIeHAyCi
afjcHLKZWJiLWej0pSgfNK09FtH+BzXhLWxOxttS+2mcX5TvM3SFr1cS0o5/QKPR
ptPt6Nk276gOtCFgFLYK/L3iJul2CLpHSVCpyyFYnZanYhyS0LFZBWMhreW2nd38
pi7bKmI3XVEiaLnevGhQQK12bgiQXbY1dyVaF09Fjh2n6LbQwmvy2Blr05F3cWLd
3jybatAKBCojQdLtQVVEFIViltDZHRTLF3loRtxC8c3kj56Y2QQ1nPVjLZ/4b6kQ
hsaw6yinAv1g3vcxr6/+ecvPAvudNz+azSGthvG16qWLvjOd3YlnLxwcQGRjZTFZ
3VyupzuvTNNzCUjEi3/rdTS34lfjuuYoLmB4vUz9Tkj1RPCPFUB5Ha+Iis0bvpXZ
HmHR9CJZLvbmW9Te1dRdO4a8/3QMqYgqkdFsIN7iabETZ4pzOrz/S1gH1YhG6aXw
M57bMW1xfnkI7wnQZ2kgs780G+eIXdcvwhia4pbeFmu6nkMIOpjyZFDY7bESyc4o
oRgnG2+BRN4O4M/KZolaqa0o1Mzm5LJoc3jIT2hJDyPw7oFjwKGoj/LRYZfsEkN4
4Qq5wQHsjs9O3f33aJMX4+H/Qa3bXqllG5R6llv3DJeX0p9D2I2iAiWnqto3Fp5j
AIRQWOAtuHrOI1I49IjIVIor7Xlvg5jUfe1LiW9T+jiYfRfQfSUx1uZEcAELiG8j
5XPoL76QFev7w+s8QJfL7phy3TWrM1wRVqvOe6CA5kvKOyO04iYKznWbOrFVxE+p
MKu/At750Sa2lNr+aVSPwJZHOlKOI6Xnvqb8NGZoI9MVU9cAX7W+20rtA5kCm/Yc
RXC0nO+ntgTSeKm1NyyOyHa0++BHdzmK2iUfUntZJpLBQkUBNVW5QbgPQ/5cT+1P
gpuAjL5OKsTVVwmnr5uafPP7u19pJB0wrLOTFlfA2RPGkbU35IugdZok3AmRoaqi
Gk+yLH9Qp5JM5OLD+pngmUnG4GW0kgIbq7tmAV6dnSG/QE9UVDFkSr4G3lHrjDFQ
4XE7onv4bVVdUGi+qHZ/niVgHZrUdB2cSvk525DLkL2qbtiGKSIspbZgXrL7xogP
BK//zNchZsxJzBNn5XPBT1KxY2wBFnJn0JzkULSuIDBL7/mz3F4DXOD2f+abrBvT
CspmDsvehlqBsQwYYcKdDa+LOwmUgP0UpvTYLGDKFq66agkSW8tGcYDo6j0BiqU0
vBseqf9OAKCRdQ4QPaOH5G3QOrqVArxQAFb3UPd8guZGIeufUTWvidRp51sN720F
XcVzMj0QUbzjEwtSztRnY5P2x0vzIUSzDZL7Mpkws9Y52hANGE0btPeP7vTxNUB9
n74x784l+LbfzecWv2b/JCguIPeuTuF6W8tkw6zSMHTTuy1hPF6zO3/GXcd7HVhS
2r2GfoGGtwduknxMJV9E6WrsfV83i3TrT8D9QYFBTyd9RfvPmjGXRD8NTdbDak02
Z+DoS+Uo5ChVfej6YWiWkNAHNbPOCH7norTZYf43SV9jnCC/c7/kLVA32oruoAxO
4CQpG9OV9mUZnqy3QXafrbBsWq0guzzOpChjhODupbgkuirrepnJPNjaLQSEi8Xo
IjZRPeaS0QbtwglwtYHJgBftndRJ7NyPNg7tkJJC4IGMwrYyXs99oQ4hLyVL+K8U
U8b69E/PVi3hagz6wEorItsWpEpoMbEE9qvhrm27/IZfcwTojuvDaX/SDIB/0vqX
JJuD7LU2pljG2Mqgf2aTWRNIsDw8AhK3QEAbSyjdC8ZnJZ9Z1tRe9QbDXbjDVsII
OrEbV4WaU4BrYLqmnf1PvBnagfUmykWD5T6dMNqQCO+8FFTRBgX9ND6Nr1kx+jom
dBoVQVnu8YjwmPXELUdNvGgnZbcZi7XqGMTyhQx01Ktg5CMMoaN76BX1N5BaXxby
KjrrDyv4SIUTAA1jI19ttWGfdVBSuDMBo/Kvvu8FItK0FIqtnjW1xUEaLI7R1/eG
exClVW3j/cgZbKA9MyZNGTkPRuE72IVsIXB/wwnBsdsWk/zSsQRReaOab1p1KXk6
TSXG2ncOZpe7P0CbBdIL4IsMh1oGi3Et6Eztd6ac4Wj7nYvg9ABJzdqqAyPmjGNH
Ar+nXSQWrTaz6tgDUhAZ3T3DRpRKiAl+iVRH23VIu2vt7BVFtBmLi0xNVPbNW2Sl
kOY28hSFSxK1RB4jcbL8GtnX4Jxq1f6uuXbOQbUTNIE6G1fTUNgIb4sNPTHD+uZJ
sSOdy67GqqfWhwivrPWqp0fQM49gSbHngRv5XyNcRlyqkKnabqAnOisqVCkfzgj8
WUYEsrEYKFm3XL+bsKUiWSgSLoNDNY9WKZUpkUEEZ1lyVWWVX9NEFNrJwMJSbyw9
KydyHnbp9qCv81wGrVTV9phGG1Im5rPE1t9H5AyvCPfNKyAOy3TKZL0KDI+OTrK/
UVuHWH7tf75teCUE9BhTRAsbNyGStJX5ySc0dSfTtcpoWsrj/qbzMiBGp5bvuPho
luokab5qVPghy1PFf45W+A+nTVS03dfvItWc58acSrUQznWaX1d46QtDTj6LxMkD
ZrIQTEYeNy/bzTdfhjJxfOIUQhlwXTnIzRESkCV8WyB2ERjjcY672Ool26AE6H1s
iBrYMCZNLsDxXaCNof+bD8omHOCrwNra7DA1L1myI9PxUEiMkwIfXcMscKPEePiK
a0NUa/KXr8jWYZuXco9J6vQm9+oNyCgo5FzKV48EKBOWkrh+nWLdwoZb5LpX0KlI
+MCzvlso7UVicWbs8YcmGAIIbSza2UsG96mjN6OxH0js464A9Gk0ZtOO77rkH9oI
6ooskpQ0akG8MZyQ6Ri2tsk8J5RFk2pH8aLOH3s3bWU5Vhh4xN64UbM1oqPYuyW/
xYbE+LuLK7tbiP4GuwAv6jzmQnRbLdQSmAVlVQLf0BEW/yrjQtVOcOKxhtdO+N7t
nRqv0t64hXZtoWwCtDSei9BBC1NrMMdHY9Toa/EQkwogsRmGxEK3zs2ZAUKPdNEi
0MK2fh1g9kbNIABzmS8mJNzxUTCLCX4a2msanc2d+3vKCOTv3ooRfQzHnLV1xnVz
rG6Q/h2Il/6Uw+r47q6fvpkLvuEAHTz9HypWzsA22FcCnK6Pg+Ju8Q7Lxe826LQC
eeU/3fQSQz0YJ5htzj0MZn073O6HYqhx6aoI5CkWNkqV1cmFKoFeKIVRHvnSzuJu
XJsk2ZgA/exdKOPXmdq8PcfaMnztAUWSlEEMpMeVpMN3eER5eNPNgFZLNFm8lanJ
SypN8Ri2590uR4KsUNmAxEkyVNoJzsMJxM92/V91q7Y5aZofn47D8tZ0W0Ya9heQ
/oSOkPQ5Nd5Uo5fqGHfzPGzTUABJ17QZVlplkF2IvbD8EKKfpg9go+2vyeCngG1z
dDn7fPq20jb+SQuq1BnHLP7rDvF6lwYVefbBLofkZ+jXDey826MoKt1zeIY/aDfb
p7hkJXtfKEndBw6+j5KhGB3wZIoGJm494cEzpu6yzcbBswlSzvF9+oQ1opowZBWx
fNXOWPnvUOgy0MJ4zqD68QaezguJlExMJ0/yFpcOdPFUpQyChCLtwi1ZSzi20QN6
i5ddKP3fXemdAowuwnAyr/b/OrE3av2qGvKmthjszruN6K2luze4gh3lr4ozKGtK
+ty1/5zaRIuTZSS9K0MqNdUEfGOqYgUzdMnth/IQFtmG8OPvkl7oOIpsB4RmMc8E
JIf5dje8DtkSrNT4uRsIzcC4Znx2xwgQcggu5BuH5RDzJ9xcakVBtR4N9L99YdCs
YXg0b1qEWa6YCJotLTvAdoRHXjsNqg/qg5CnGPAVOs56dD5rS6MuzoEv9ejcx5vx
C81aPW9lZKGKiFGq7mYPMF7EV9mY9ReLLH0qLXY3vt9NPCwlEsg3qy3HjyzFVBes
STXlDonNuQOoKu7L1xfvEsXLszZi4lN1x4Pno5kV698gLiNWOr//T0VtBjs8EWVB
eb3KFqDjtkUKd6nlsWSk0xvr+XP5Qv0tHMxjElipOwOVQwDxSZzeuEx06VNDyv8w
yM9rySYfoXHyxDEr5ISjpLDYa7xnNEqWpIVKHMlQQkOtZzJCLkTETtAf3zcTRixp
EipbZWocUgfYiseArkwD+NB9kKwadXkiMXGl3TQKzREAdDvmNWUACyVvU3VBImcj
RVN2Ui+ChtMb1zw+bkPBj82UrDUAGjuFH+C7Ph37XJmLgjy/wb3NFkA4f405mkRT
WMBq76L/rx5Wx087dNxLP97/DUFqsQ9QCG52u4OqQnVy+LuKPEMn270jwxflceXE
QhHcwnQ8HnEioscVvKX+QWRGI+sG9sxvYc8ml+FCSDw/PNNCVZ1JEUB25qVDW3Oj
hCCaLI4qzc6A/jcVcsI9HQiez18P0u3zUhE1CPp4v15kG/dUmdyfJJ3S6cIes4G+
kdlfXmbNYDVI70cLl4NIKpcB7LiC68lyupmMQ7fx+G37WPtN2yYomL9IURoBVusR
XE/6CW0g2zA4EwWA6KAggPU7fBrVj3DOZ99qpyOD0OEtWl0NGqJnatqb0YoFxQ4q
uWkk+pwh3mUoG1EY+Ngo3o7IMRMAOO1S70obBPRNFl1omwCiqn7FtMIu34Zbahh7
4NkUzAuhFlEsS7rZh0C0sAHn0N87uVKvgSXezizzTS1MJXNkl96DKFQl1rlkDPdx
UbTP4y0QmEYSp14fNWiwthPJpEeeDUIDZ6V8xmw7NibKiZPNjUMLUuro+bzgHuxt
ke1Smr0yslPAaeXDnAgyJsyX9KOmT6rK0eihjDhq5DH4XcraCggEtM3DnPj3NsLl
IkJX+3bFFmmLFQ8VnUqZcgNByvMgscf0h5DagFZ6Fpdtt1sFg+HshtWv4rXP16CC
P5cWdM45oJyYlB2nKio2zAbBmSeGEFodrfDXxjioKJPvEu3C80h5lxFKLiUlYylE
5zvdmg1WYUqXM073PqLimgCiX5DDuO9aDUbqk5FJJdMvoQacfezbVo8IuoaKJVVA
mSvm2Vn1UEEZaWUY7Gu2THiSDVOKldW0zdvwyApOiU19y2zSCYmLKLfWsz6bJ7jf
nTrcDWEV+3kFfqbjcLviTc+EumhDt6feva9GtR6I5OEo2QXsrGKg223Zuhmw2zFk
MeHlZM2ZK0RQND/9iyiKpYy08FLJFwAR2kDaF3bPDbXzjvilZJxX+CAk/X2zYczN
czUk5e6q6D9l6LOUcgUHE3u+g5DG5ZJMaDJTlXHheFxFbr4a+YLtO6pO7tsFk96c
56mC4GRboGoXqvZYBRqEkuGZDQu5SpIy3yJLVCRkFLu8J/FqQiEaj0HRp+0GbEkH
iHSxq9KywIKfJ/XKVl5vneNxJRrsXRilDcfPp2gMnNhNs/TOtOMkx+mcWky//i+2
7CXnXjpKqUoyR8o5SNahOcdPn/cyNgiqOUed+n3FKwSBCtpwy+i9Airc+9X4jTS7
lx2F8HZZWjUI+Xmr5paY+qnqYZSAFvWJRuxBb4nBWL0foGL2zIqt1By1OybxdNtL
ZWWmw4bt1Vss4siRgyWBi0DttjNeifwlG/IgUTLFAzNkytpMO38Cn586hN2np0I6
DPrTDcUcsOI2A2zMWPWBksiHsW2bh6hFejFYc0Rj6/7RN33CBR9e86LQ0t4W8lFE
BiA2llZhYs9d2BHmF4Rfl5wSkSdkPmgATD76SV84SB3doVoYVCn8J89UpFr+G+hd
+j7TFyJXt//obNknbapBk1DjDHETbxfz2ClaWo70O7LgVw+Ws8of1rNDRX8M44fe
necHk6xRWZTSpEmh0wheP72jXyZxRmsi7v3VjD3jedeqpMPFrSkQriQAU3ceK5cQ
gPaj/LhAcdY0Le9WPfPYFvwsv3cjNUA8lBQBb15DkYQ36vpmgirvYzS3dBNqzVe2
IAwcUDkP9vU2NcGBt9Tvw0K2zhydJIPIh3JVFpNiTL8xpNy+mTgndODztwCcNslD
zZ2dpY4YeAzPnekTHLcPxvc4gs5qvydq7ancc5NSmvXTP5pPcBQnfGlOBI6zmdwv
yBya1sH59BfxLLzNbVcBBjX7QWh/8CJvR9n30WF76jy9ClmPanTz2MLv+PNUsOh3
2A6pCxlBxSH8sIpOC9T53UJ9+0jVB+ABQ3dv1SfBKq1bFJtkh9ympVx1oSgZIy2P
AeuNhYPqXIcmJMFTVj26DUAjcvjh1EiNuV8Nr3uQd9a5nqzSsVx/JyctwfgapMRq
hj5foNlLrOtTgmtM87VeuYsPopKvuWb5Q3sJGTsvAVjLnHkIbXuSBdneBDJcVo9c
BYV/HJ+q+WGcc5mZ22s8fWH7re7CoM4KsaJdxvJAEXyZe8GORvMjhmj02Iy/4IRn
dcnXeHhJYFZSDZQrvzd+1OaivBg79b9aI/JnlnNsT/E8q+SEUAx7VmJBHEiOB3rl
gL2JNVMMTiCduWbjn22l215uEPiOxc6dehGvNDJ3rT4uBoXAI8D5V9D16m2wxU1R
hzNTaLTXPWbI6F6zoEk0sxlAM4P8TyQBcQ7AEt+cTH1/pH0RptsroQsie5G2yHVD
lZIxfx8NQ6u++rwsGsYMIcML1u6VSvUjxEq50IqPFeU247qZKTEFAmuYqZHQ44Rk
Y119021DwaYZJToyW5wMBGh7MSHDsSMbHhqI8BHcwGX77Al4TcxUZJseZuN1MyUN
4RgQaqt5LtHN5BmM4y3ObZ3nUbEXO1qO7tDo5KxPeKeibyy5/30JF7QB++doz/US
7vNYyVGxV1wuKzd/h6Em2iEzL1iPG0PNHaBfIoScGlMHAFKfsvak+AG5jqUrMeHf
jiY7St3m3tmSVPBS5H1oMWrMV6ZQweOw3ChV/nU9Oa5ow+VuRGu8bHZSBTGfgC5F
tGsuFxV7w2DoR7PreMNOP8rgESto5CcY5AyxiW40iU469DVEo8Ik8trPaw3A2ra/
gexDTdPOw9FHkgkuVcC2LBWh2p82Izai4VcVQHmKtRaDh1YOXKI1acpjGN2l2HBa
ms9tP+I+9WhF1bfJuo15/7MMnv6+VCAaqjlmsKO2fViNm/dwowKyLh2sQAN2qlUn
OCYAv1wc0fZ175L7+xCw8k6lgLmYsZMswp+OOsm+2sv6+8Aoc4hkDKfhcRppNvin
LDwoAdiAHM7uUgX+Sx1VL7AadgZYjwedddfUfH/mFqGVGnxOwOqWjkrJZp7R62ct
RtOjwgbpJlgc/My3YIA17QlWPXfgGM7c1A+bRrhkuqHdXBqRZ0P0CWEPB5GXTQqS
ZDHV4uTA7dVNKdgOSclsI2fGr9SnbOzqpHs2+acXb+VF2uxx65/F6t7SEMYPME1o
MArluiJf+8nY23iXh4XO8tAzBZsSpj5354HeMjKOHzkjLIyXrDN07sKlKbWRg/3T
fISVXoRxNj/+m+7StPD06CfDSN8SViPDxobmtt1UvlZG6DB9R+Ti2RlAMNEsEuJA
ODRFdWkEqtQErYGfdkyB2yulSzVqqrzwgbM3aFoC/pkMrLserpD1cTgitu+ZIQ57
l27NbWjQJWsR3qHrCOwoT+TPdq05PeRlnXUi5ym6Nfar029SFZFe+IT8k4nbODFO
Vtw1KxKryb8VMZOzVUdIZ9fxvyiWqpkznFFPO96pw/RKsDVVzh2N7FkM/dIURTio
yecCVSWNMwQHoIfZUJUlKHcHk2n9H+vJeJ/lW1No5iIG/U/9qL1y7+IEh+jCRi9Z
RhyLvUAfdKC5bAUM3iSiUmYsLHm3IFejPhI1jDwSYO9QtrYDa133/FIVJ5f7L/uk
x5tLB6mmvOG6+TV5ndmC6CG37Toech1HU/HvBTaGSXk86zr0qAnEooPBM7o/eqZZ
HkelfcaX2XNk1rfjZArQ6nnRy3nlipXbjIsqxJpngCdghU+ohAlrE0sVOJyudGAC
w+hAx7Rfb2NSn58zVfdBqKYXMAa+LZ6puVz8ht9AySbmkiA+OY94YQanP5ifd4z4
in9ekEIlhIOU3p5OTAe8LW+rvFRVyBCpzsV/+AWFBdxCyVbi7X5gAWGjjQu2pNa8
vt4MUM4OtUGjhZPba/JBcxQuKtlQpXSdyQEkE7ijI1qTCwKYFQJJX11QOKg2L7r7
CuSdnn0/7Ib51MiU8gaDMx1kDPI2uJlF6i8EV330oHk0s8ocXi1u+jFP38j55z/l
5udQp8BBwcErZiOWo9mvvLMD20NJKjp+jYRjpmohJR4f5yQG/9ewUoEZLol5aZil
P3g3xaTsHsa7oeH81jSuKe8V9/zmrBkuwdYA09TktHcs5UNqqVNEsZiOqbaWDqot
ZlQ+qkZNjzOlBQh2TBC96B5fyaPKmXJ7D4rEJMmBFY6rTOSi7HrZUQQ83uWKSxUg
Zg46GX9m/qa+Ld9LrlHhaI2uDGMWP0cg3t/irGf2EWQL+DRSwqRN6Pr+61t2b1Jv
k3DSaqvWKQZFM+hELlLeO2s06IbYM5SfghWrK9Vnx2drGowkOuWTbWNLQTOnrMSo
QBYiLg8qmiX/iHF4dDN4is1UwzI4vQnowiE3LlK3kAduvZMbowsVYywZCMgeeK9H
1FLzMb1WuKtJsk4Mxyus+3C743RWyiGdC569rRBZiSYrdsmO4JX8ZnBYntK1rTZD
9Gf2IyfnV+93YxmXdxPahcxYxRswuF4Ketc4piAq2NvCV7PzLqYXqiXoAvo7s74P
kp0TBDthXwJCgI+Zo1pYTwr47nRU91QoHilorFBkhj/MvTV5uTUjwj4I1pgXt5bx
qwkDDFj9bYv2HOAGKG9ARfTdC1xBr11+vPuPoWabR7ZFmb9epGCibmDlUyuNr7mb
sS5yMUaAF0HL7E9nkfdl3oqbtvwVe1QQGyKfw40PtAt3mNghpxJEj3P9EDpIHFGe
Ams+tJA3UbQ4+xg3K1nLw3qFGDAn/7YFVy9wB8J7IFUGxErlmWJYPljLpgG4uYL/
0365z+uvka4+HwbiAA3YNnq2VrjFoksvP6SU+CLSAJPNzUI1CVa3aFx/rOqwR/ZV
oA+btEU0eVIHj+kPUA3QKyynDPpqLHQahyvSOruEP/YvH8LstoPje5O3Hb8UdRe+
I/RxHxsCyawS+EYreP6aBAgN0CbgeKPAzm8vqrclBMlUWghj1f6fV9k5+NAi50eb
rs9NBqVl4LYvghKNb1BualU9dxfkOc9gaXEU6aArGiu4iwW+G65kvDGcdFBLwtQy
VJhRewE8j6X/d/Hgy9xA1lj773xAWxOonDos6bFjfdC4791QvnSrfW2UwAGaHwIy
2nmWKPnSbSjxZWEM9WFPX9J4acmTU/5sz+L6yYn0K7hR7hwLh9rIqwyGDWGnMebZ
jDEE9bGszY0pnZMyrQ3xSbPfqLPKQpxLMWAcbG+ZeKmkJxiSrK+6Pp93dUI/Iee0
U3oQSJ7yGOX70FCZOFesG7Oi2jaNx1OxcWpzid9RuExD4gj5f4wnvgBdeqUNRCOv
yWYlW0PhaGcSu0h3oWDRXQ2XcyHo10bbgFUispN80KnN4Hkh7RIeMqll8Y9AYiBC
T5f9mMpN9fO+DtCWqr6pTe4dFBAdY7ys5t4+i8xDCuJv1xgh9YoOEmwKWrb1Qp5U
Feh+COpqioV8VcYuKv+Vf6b0cyhcWKaq508k+mRfC8QPpjYbPxhtv3GEmtOcIZzk
PJ5Dh4iqS+RtHk5sO30ENd84l1u8YawPqwlzT0knbImxI3aA7cz1Ttp1ZvZBrvw4
gfS0XG8R1jAt8dhj6I2BkIRZEprf7YQpLCe253sfrJnleXJNWbnAmIsLPXHv6xqu
+qpTxnwZbNs0uSDoGjH5WpEQyCi1VPGlzS5EXDcz5tg/e6eCvmCPT3pxzkfxGxLk
dHeBINwIPOEwepYl0X3VyKaGz3EZLv7F6/Eda7B9LeMRFU8EU3z/PLXjgmSkhaT5
eA1V9kmoBLYb9lc2TuBvuk63tkdTN4SEweIcoUV0A8+hqpIo1wE93Ql4vcRKMDa1
YSnPR7kCy738DTX/KCAUsWVV9FKaz6cG6bPk8NY/q91RdgxugRFjUPasTivOH1IK
w8iW4/x4YVE1eywmKKock3S2Jpz/VfKqGGRczJ50/U6SWIO5c9Vy1XXyjpI1n/IW
0EIRQ3tJED67x1YbUuD8n7CAdL5aKk3t8wgBFbtktC5cnuZu+IBL6uTlseerOv5M
d2X+9RnvN6t4G6gNh2bXAFkw/5eCdTs9s3OMlquFenA1awkQIPEF6Dye2woaLgCj
idxi62poV6T3qo4H3jhbodr1JmuIaC3gn9Mj4qN4RAIKHNQlVeLvaKLAzWNmt3KS
g0lABapoaLr38gAgMa1ELaGAa9OLSXX+G5VW64xhfXKej8su3AYv7UgQ2Zp9rr07
s6PssVdcod0MGcElfs2msbzozTUv+lNciYV42asmNhAG0ZUR1MpASWWXobi4Q1CI
D69sHbh/Hn6M6FaOw9sLeW6eChC7/Yh+i6EMDbP4Bx6e7LkEeW/HY03TtmesAAz9
/6BO3iHotqf+N5/ZVsSp2d4LEEhXuCH54lK3Teov3RYEQRdM2EjvQgQ5Rgj97Y6E
HoRirWxKg/C7gWJEx5ANwpSfUVL6kExlLUKb2JYLCze49PjB36Tgh1q1mI0pE9mb
GNe6CG1kGmUF88QpnS8NUsTQcQi//258hXhApxvhNJLDKgSy+f6xGvpHNl0mgjlE
egb3n6XJdUFE2S0f6Wc0rilpBy1/6/2nmha6dly1zSxOmFfxUmsM6akmg2Dz8WIZ
XOhruBv8tYC7KS9TJ7AwECEVaywUrAosSgdANzPxL7adzuRkR9e+R3yvuEpGSDCJ
TToHBGFtDLy07gFGxhPn/XdHutDhDu9GGzr8cv1Mt4pd07zIbz+PNiULqKIryMfw
xvGhg+I1OBThPZMT2DdND+nYW8iSbzRhi6dbRMU/z5V+tOvR2g6prhvljvbMHdtD
fpDDE80GensQsCen9SCMuzhW9FDJx7QA80EnS5/Ja4i7YLJSx6C5rQvHQhsIw1ru
0JeZLWOqTYnzgqhY9dJbXbHaK21jTFlCcX0cZfvI/93DjIKtZ1DWjVTl5534lpBf
kzGtuCnfh3Pe9R4WzzAoHI2t3iCTJnuBT7GGISq6STqI8DQD+AKS5Hx/BUwCA+2a
AL0xovXnJ0IlJ9tnHCL641x+L/I1/C8WWnhPETLX4oqE+hoS41/afmkh3aOZrXdU
yEcSetIkplaqKjCztTnnrJaeJOqRzO9l6/xa6aq0ihof7NUe3rQJya5pWdEXU/tI
+oVTIhTKSXb3e3yAC3ZKW2gT9ImmEPwOFjJsOqChANE2YshDnEK9F7rkgg2DiOtQ
wUFImBJPMOkTIsDfxMo+l6T11T9+L01VvNCtOxgyRDq2LZgQm26vW/t6sjD3/s/P
sY4ez/lZLU+J/vxcopkhPRPMczkhYFGlSx44qvP/3HErvx7qi/gSCknMXC02bi9j
5+I39uKrOF90HB9AFMMkt3jxxM9rDZJ3C6f864jUUcd2jyRdqes6gR9Ei2XE9+Kk
DGx+7FJ19JUb4/cXMmkEDlOYOWsGYqO8U91IYzVsqFUAkD9AwZv/CB2OpG1f6A6I
8WU7NnirpLf7Yu+j7EElcCyGkIHQSNK/dEuEknsZeRenA/cwzL6+uJ3+xF8YQIjB
wjbWLrhtaLzVZXjTaO892RXxWB5DXx8dv6Pk4EptGAcjr16P2fbzL9xGoaqzXomX
4VbsMukAuwsW0DRIGwntZvGXKvt/7ENKzGf1obKK+z3BgnA8oKCfBk49KS7fTcvp
5hM9xRXSxkSeZ/Auv2Fi6Mkx7CpQVtWDWEP0l3+caLgQ6GlIXxXCbIEdVJ24Ho0t
NJvdVL+vf9VblKwkuYww8xyfCiVSlyQ6VB1GiVAYGS/UyI6QIih4qfJUBZeNovu3
Pega9AfPoRMsVJrvFmS157DjNL1/Oqdbgktt5XF9KsANAlNgs8P9I/wsL2GM9//s
KoTJ7OyjwXnmi/n2r2yCVzbeaeyG3/omiwYT89XrN6nMb9ylwyH/Xr+eNn0gAzJl
/S7YtnVlei2HeDV9oPb+g97XzQhYPSGblxDd8xGcotxMjM/j0SeXlcE1LC4+fNRC
ulonIMoA5xqsdxpz4ENkK0c0IzV0m/kDKUfcZ/bavmmt7zavsxmolW9CmlkXFhcM
Dr0q41eWeefd/JaIkfhRCgW3+bFi3p9f8AXdiAfdTOXFBwSGsBZyDSYg/vxwXqhe
r/2QwYNZpIlI3hnO9dTzCSg+zB4EXvZmEy3Z//DLYMoRAHv7fRw0ILUXiF6WmRrQ
fQq9yGDPNWiu1pfKteimBVaqb2CAg56NMGtRyklH9iOc+QRpQOAQK1CUJeWQ6tER
CqppyE/Jtdqgmk/E18a4kPMk5XcHep7BIEjYMmRN0bB9xZW3IMaGBnF4qeVnHjmJ
89kuJDJhtMK94/7s/HPaCCKY9IP1A8t3iwpe8j8vD/osUmpXysmRHp3L5ildUOD4
wZC2jz56dtJsvogCTO+rCbdy7v0MFsaAaY7hIb7aytJP4JtVrfWhH6aDjLQgl1PH
Gd6PdtW2DTcLEIyNdpity1MtyiqVnehZRhMpbxf/hocFTUESX2lBZhN+APaKjr0q
18MH6bjbFs9K2V4ka/24NjPC09kGOyxC7y1uN5l4ns7huLmjdsVwwB7q6i8JgFwk
U5CW856waSUmCdHYtaE+72OGwiLeuDBF4uvfzOWmvCxAFsnIcfRJE8cADhDQpY4L
tqwhSV3P89k/u6/ZxsySKIiYsaUs6nE18Dpw2epxBqptlrWn9FSRh/9ELa02FDTn
cI1E+Jpk+TWHeZkzentmW4z9VfatUV7f66d2m/zT1TZnUo/nnL6Ox2uUoPPQNLFe
oLtPij4LlAhp1xn189ae+wgVpBhLeoq2Fup7ZUJ8f1uT7yhgbfQFGFP5icxitdz+
Jm09LLD1rA8uMTTdf/zUC+sCGfEBxWhLiPZlS+SbbLiE341QccCh92+s9y0LSPLp
P+KZXsRMK8KNZT/9tUS0CbFvjQGqAn8GUFt60YF6cYDsYbJx39OfDVpu+8cJ6DMh
LGB9XLbjrjtCO2qHO2hwB4Oz986YNo1X0sHxSmDlDI/zPbUwst7N1PrKIzHVIfe/
yJPiitea36cSG9JqLK6HxGIbmBzcp+T3Xq/G+glvT+AjuPIF5yYucD0ShxCvDUHn
hD1CEpaVa8AAsxchoIMfRFR/7Wn5ldXhqw4jvblUHxPcKH6CzauxY7aiwwLInqe2
gdEhxW4Oj/Iza5Y2tPiv2LrDZfGvVyNcX6Ipk6gRhzYXS6yU1Tqyh5juZ3YMbdVE
rCwZePLe8GZHF/egqDabAfC8k25OS/M+7vDvTEDO6t6RZpxVknvp9j1HBNfUMVYZ
U73y1eDbnSvNSKhMqUKHOU+/DIQUxSGstXFbJtZuDfMOTR7FEGZHzsrlV24jTyD2
7g2aeo5lI/XXmtQbBT7ZjK9fpVY3McC0hrKV4XDnL/hhuDv84ySRPsWSWQLskiD7
4NJdUJQtjHvFMwamjlk9hUzB9GaMQ9baZO7kLt0VgDnZdEFAAGoe5UjZCERnKN5T
rND98J4ayngmFtpuFGwK9C8yDghrB2tOLjmTV7jvvjEpTswpsODGH4wtN9LqQala
diFGx1t1serKKPIhWpq0Kuhjvu6YJdSfhcmY+Jvxdt5qCelnLVrnbHuRDMa69dgq
l/5fEvsZPs4oG6bkx3SJH5nofZPH9KCTlwtWZPZdXQcyMbqgZxCBg9izXgXvsbRd
NICJyL1Nk2e4iouoGjaknSCx7FGcpkhHRvJLpHR2ozIn/72M8uVIMkbYxjKTGsw0
5xbe/DutuFST+U1g4CV7bSA/dGougn5IIGaqWEB00w/QB1Epwm8Z/DSXpUEntFu/
DWG7dZwudqi6BgxUo9X7fqilThmxUUkoInB4O8+E2AzOfvxCTd6vIbFncGQIWLiq
FozFrN6pdDmgdLtlYUueMDcB7dZzs3t8kCAGl3O+4JBKan6XgWk1QebXX2ZRcdm/
wNn5IaXQ5rwey8N1kN7/LeOlk+On4Ur4POXxEpncwJrTdbxE/Bi2P5rRRfOrkRIF
0j2QBewVIxKchAPTjWCuf+QkaDO0QB7nT3iXkSd67H1HJ3dkTHXWRhwZgcHE9c7G
evda3Eza/uupMh2aLc7ygtmFHx1svog9o4WRDFDCe44TZ4gXW7XPu9ldHMLSUvuz
LNsqRAKk1V2aAB+ZDkg41a6wgqE4IMyFXHim3nEF797MBrT6ljK1pcYuiURvxKiF
t4IfGrWx0j5n9rvLdYd3QVjTK2kKDi1qyV7FpIAtlQQzxe8DCHFgGi+OFAXb1x2S
RJgnggtRvS5cKQGzdE77n29RlQdfhHVp79ta+Ik+MwaiDdmw6eNviDgCn5gmR2QR
q2owewJnPnDUwL4uZJ+GeKLg0hY0vBAFn6Sa6RrIWxKpjr6AmeV9E8z53BhAixmp
CLj35LDei2Jy2Xjea3pfJewZzGp+7oWL9eVLkQUYcQUylDPUvCQjFVAUvuz/snL4
B0azZOFGu52IaLyMpICOm1dZYott0r4jkvBJTbSnckjNWEPfIryaKH7CGTNZLscf
BvGB/zdO1mpz/dawBJz4KvGfC1yEkkIA9+X3XrEupDLoMV4y225o8e61FZ9DMbGc
01y5kzjLca6z8dZmPTOrCmzNM4Rqk8IWUn5ZVM7VD31+P22msAWhNYnq+HafvCiM
DF5kaq11vR666HY05bICi1wsujOR44ZcFgcAdBeCI10+Acu2DiBAhc37unjFKHaG
czCxKKF6zCKhcRUqStAO7Kfyhp3o+pnHgC6dNUvANqm8JXpHnyjnFAFe2J6XAlpE
ANdUjx6/4qat2enpv9Rg3lN0LxhtVduxZXH99rzi8s9Qxg6F2ANjTzzE8a7W8YaT
O3KHg3/Ej1tW7dR5toNmi55wfA9Watn4aU4hUeEThvB8s5hPbL4L59a6CV7oz+LB
2jH4HvkOVFK4b5UQtT3VDCZVOfSbCwbmDZ61iF6l2x/gsiaTnLGrFqjMFQXuwxvu
IZE+q8838Cje9+lQzo7cRQVkXG/C1C53BSwyplnorl6dq/eUx8W/rwERknE5ucPb
8P9Y/trFYKihbroj3akyf60vHo64vyMHijZtKhUkVYlemvXmYJB59JlqHDgST4Qq
YoG9kUmImu2IAXCNeGwrAN3E3baLWIycgUDNhHa34UMrwNudHnVKT6Mx/UJP/h32
nmxovJqf2suuURLCmrbF4ssbSEEbZlboBQVxCkK6eyZ51I/yL/cygY4FeIHqN7vp
mkaNkk+WikF6vgfaUfxvMM+ziSqVGMHrvnWpPYIfQI2W3F38oxZhhdGJfNed7xGr
S/bUuw2ra+thfTia7jdB/MkMUZeGkSis46WZtb32ge+F4BOs+W44osxSeihB73KD
DaMB0r07bNAEJuv4twfhTiwzm+qF2AkM09nDNdVIsZWx3wgLq3czCRj3r7Eu65vV
IKAclWJoyrt5eiBUNb9mNwm7NOhUr55OzbjI+Aj30XUX0sfUApofQxIs8wfYd0Il
suguBSKw3mHo3WbGqk9Cw1RA3gQl8cjbBCoUGatwgR3xH8x++WEW4Icwbcqs5hJY
N2vnKPXFm6ni2ejZMD0oQffCZ8yJL+lKQi0I9FTChBUgMNgbgdUFTYRzvOMLbUgw
7bG0IHW+VLKWQR/lKMLwFPVs6dOxOEIkVLyrVBQUYWL7A6iFBo6yfIFx+DOzV6G2
H9P2wdw5mh+ryyPe/TzMojhP9GQ375KvmP+0xNWpobkK0WxrE09EbF9bxtWlUg0d
Zr5jfuMoOII8yboCLWJzlEVgXeCqQvkXOJZPvGeiUq869mtXS8pp/a2Tk8Kqd0NO
lHnhm+1/yJjZHXDc/RY6GxFikzvPE76AuG8m+e9rzlIrrSriCrBdd2TTcwjTeLfs
bricV4Do0CK809rba7CrPKUird6C7AJWrNcEBUU+TtJqJPJuUYkPQAWXsRCkYhz8
WecLKFWa1Z9V0hAjptwuKMQlsq7OPz59jPnmIGF2XovvAtdczB0qpNt7CBoipNMF
9ytDgqr2Stg+wyZ0GuT9LFQlY7BpG1DlHSAnp4C7GHHIuMLY/AGLkFB7WuAIxWKi
w9eB1jRvJJeUUrgltlCz660onKoFqUTIB9KqCPNfVAOrG69AyOUVMfoQtO0AqpgJ
7IKGhFCYFeQ05r+oRUWZU5h+APg9MP0xhFak5QJGPQr9LH6Xa66UCFUHW7SY4AKu
GjHxzCd6AxmB1EB9sZrs33Pi966Ehnl/U77uNXMhRlaK4tvRMoLB9E1NBwKHUYzL
luz237aD72tzaXBH5tib72QS9lq8kOt1frUm6yNpSAZAFhqH25pvTs70qxzaTruy
teeVw0KoyqyIePB7M5fHa1w75W6rd8sgyU80iL1b0Tir7bD3Qee5HROt/tsdcXpc
GlYnhZFO7wlx0GCyUiqCVz5mhVLm+hM6gar3tWy4IjpN6wJQlSYwNU5zAbwRST3a
/6JAPMN1onosEKePEjQDSdX6UVlNbZcKhJ1bnsFV+ENSu9EFK00P6ZdYYDQH1/B0
PSHD6nDSjSjl1bsqxKsj73xe/InsGO/lFBxdTkmdFct0tbd5uw/L3ezEVq9ggDY/
CB7SWMk3dl9KHLkRp9o5jQcoBquivIxyx5Ax3HJ2FW3EltNJtCsI1XjEFGoRJO/r
qgrX/BTkW91QRX73YJ7d2cROexnjpd/mAesgWMAI3yvoa8y9EjSY3BmqU+F6ZU3t
tmSjDxIhp6FJFg94KKhkw2YxSL8NHNVNVMil2RHzRfpHSLwCqa1eVNlOiUBFdNvb
WlIHle7gO5Q/Z1FddnMy+SjJqpKV0YnZm+CgfQpwIpPUIt+Xq1kjP6myzUee7M0y
vfWGRGXjgKDJumnqgboJhRnvwDrKP2Bxm9qkISJ9Z+MQJDW4KV+TQ8jxss7TUgmj
0fhJMk6qgTfOXATMsaJTEP+4voWMVlvFzmobj2WGnPQ3wd5HHHJ8sjaL6zXzwGUP
VhbgyWSzco9M0nsp33TFJfwCnAliPZ8BcEjYqQi98tcP2J/eWxhxoMb/ZodeHOFV
+94XRb6boBhgIDYwVLqvTu+/ZkzojD/GOL+hdQxU7WCCVa7WqEzLu4RdjWtitRUA
axrqSfMpOqL4d42MZ/eyHvi4VoKGinxFjwViDBE2u96YocIrup1O+J2S5oJexC7W
Lks7HGipe2weyk1h8wGbbkOogEauB3PVh8XT7EKtfruSynly1tnXvFZWbc6TAGnR
rDkBdlsHKtscFGh2JwveeMm6nXfIbNcS7He69FSkMATQN43XokbIbFN2FU530bku
i4NYg/615ziQ0AeUnoKYUQ3shqSuh/ERpnNp4B47x10Z8l5dkU7KXJdC09DPAjyR
/xWlrrJy+v9ra3MtjqMyI+eUI+DBjKlXu+U/lQg16DZd3j8ZLvGcfF4HNmBBCBOU
LTiatT9x/EMkbIIK9k//K4dl7XmVrj8KucGvUsFwJQ2FruvDEHjCpAajxRQdjnBC
lhYYTmyJV+okuLmkZpIIOcKLH+/AlJ2QJ5NtNl0+qLrkpf8pEsV6DUB1U7MeWC4G
X6nBojn2FDN/zE1mrelR6mu3fYpRqPB0BBgM8S1V2oBUeOMM9gqJkKQ6kNcursmJ
tRlwj32DjUe+ljoknFIP5G+/IfBut8m+xh+fnIluHLkOP7jVznPSqGm6+bMWrbbT
MEY6Qr40Fau007PTN1o7RKC0LJyJS7cUFxk8bTwk/0QTayQfuDaQn/bXoL8ETf4F
6VmUvpokykSgo4NOFlP1XQHJPsscJLlMqr4NHxJ3A//+AsSC8/UYmNHNoj/6dssz
6IePCGjR4K/AT6N7kNGuRkJP30GZDz6IuKvbn8tV74zOzaxoYFGmjYQGN3vDppm6
DnVKnCTFiFbJI0HdahW5IonpPiu4J6sbz6r8djQHtFEQvoCMWvWDRJ9lGGJxUHaC
x3uvTpWtzdKbkYerxSc8ajcEVclxc3E8UPQmasZ3T7e3qriUryYqmsVqHYufVoI9
FBxBf3UOkiOusjX3AGw77Ft4BPRfwEDjzwWF2RWo4YJSQ+h2bC0xlbLe8L/NEkm6
L1Sp7muSWlCIpFcDTDChRnneAOQqL3L/lbcY7E2Ie6lPeJ5JYnX4AP25CcmXavfN
8tw/P/i9cWwrP3AT+HA3ZvW7jCGbjsjzFOqmjLfIjCDn1H4vOojVKKUv2jY4vCYG
Zcq+XG+LcrZdNicrGebzv+FZxT4anXLO07sA8qb5xx7xIfddzW8061odqoX0SlF7
QYqDzfWEm6T07elaqJ9RXFAAUSuO9oeG8O5/ehqK8GT0T8TcFF/mc+U4aE1yDB4x
IkbZvnFkBwMP9U6S0qljKfUrQkhG1r1TaqhshbXxXkoHqsq1yDRA+iu8PV1UnSRN
dSyO4iJ8Ozr+74U2HMbNGD2elTbd6W5WGfD8IecO/8dn4nvhwAE9YjYVsrWmnl69
mx/AlAiFf9ZFUero444UdqvhhUwiySl2sraFd6YZl85v5O4jfH/Tc08OOvKidcGo
EiQlUQecbMHECmWwDqJ1Hl3008Inpcu1e+GRHOhb/MoAEnzMTc96qu4wFyO4oSGM
sgtPhZiZdU2xII8zdHpPdeMOe2c81S28hyNa/73ROuUW4w1th3hMAlA4QaGf+8oR
UUXE2Rwu4d9PN3GntfTK/Ytuqd8Kv3tr+a+YMOjkCFc4T4UR/6lTbXiNpHz5QhkY
F9yRmKEmIWcmyBDheEbJBXpvS4PAVNCklQzcDQyz2KGYCnEGi7DLhNZftqkHb8+r
k7X1XuT+ECAwj1YeiGJty4xNnLH/GNlHgVKNVRN9/78obzV/urRunRB1Z38TalzX
hE+4w1dXKQJbCN56HWxXeaRZgEeCDNqwMOA0lhB73+CCR16hZarHqNWvkzdtkzwk
vgd9mQhh7w0lyUkeZC5Si/CsiiqYDjLR1rOWSOxN/v+zt/RWaBJ7nIkeR9+ZUfyc
inJBEdcC4y0g0f3AhgIdEDLfKR1ubJP+DLCBqwWeOHoxVVnDOn3BEiUg14A8f9dQ
nbLiBJLFc/jPxp9asn/Wwz/KxEvQSlUr0Q05H3XqiR6ZpGtJorTaZwLWa5Cfbuq9
EG36l9BGNijA4WnuT+IyMqGNMKOF/IU3ia34dH6DFL7NiVRrErIKKe7AlcByiRdI
1uitBncUlKF/oGpL9lc1YiTTaoCEv+XO7pakghG6ddTa3qnGKcfZusUTxlk/uaIv
LL7PGXCm3+LuMwc4QGoWdeqvEVTarpniBMGtS1TDejsTz+/UBRI7C0/lcSFhl5Xa
Z7dLeUd/Nhd+HT5S5K05ra/NETPWTZqedRg6RI2JRCriNcCtGk2bMoc06IgDrq4H
G+f4gKW9TVWvBgl6Jk6zt3lJmp4huVx2IZnv6MZtspWAU5KHXrbi5nXReWVx9bua
kNyKXL67UfZdbuec9cLjwBR/aciZ30lnvTOT25HqcCZCasI7XXeMx9CJ8Fcyys3W
WmeW3mbWbhmvOtW+jzrphiVHmqvGg67SY3sIChcffQUkjkigd4x/PzTu5mtUKBWm
RXizhJXEe/X64+Z9Iv1Iq/RJ1i7HxRYkyZUVA/kvaeD6wun5Tz0RBH3BeChjBMy/
N6rHBcHRaA+hwy0KsBjYLaE6trc7jkLEvYKtzs6fRtqGslvq5Htx8DGazOMsDR2j
ZWtQzi2c/2xcOzBCw3ddiDUxlzpYf5OAA7JKtaNwpSkNiSe7FgonNiXg1U9fIhTB
T9xoCqm8SrF5apcoR+HfEvRKn0tD6YheqybmAhL1QQwD4jZnGpZGqXhETrzirYHD
ruv1cqtQ18j78xqcaExp6+hSJ/sgwFET4gyuyM38bKo1Tq7CmFR3Jxd2oZ36hMh0
zfKnYh9Yrky5viYCG2xKcfprE1pcyocD0Z2MMs1pfzsvGAS2iUdVu/nTWZYn/ZfE
XOESS+Er1OgUqWXOLItAoC9Wu8MurzRCCMIOJI74ZKXTrWoghWgnu+I5/MIDesbt
mIICoeAdITcZTAnAZLQiIby6Fs8KJv0bLbt6SWfjDxID3pIAkSRUkQHm1gm6PbLl
K23QN8L0WjXryxxau6OYTxBvOyZP1KL/BTyaXSgBoeHd3ks3qHQlbCvv5uvAB2va
K9WfwW+ssy/c6b8J1kloGTs6pAKQ7Oof0u1hM15L2IIYvELSZxPuNpJotKqdMizd
MjEk00eE7eBxBGGABY1wFrbOT7Hhd34/99Rz+7Metkav3oH2zQjpZHEtKwm9Xz6F
rnxseYd3wzv8gnxzmvTd3zNb3wHB66wo7VB9bK8ZMLNLJy8SmzM4hUutld+SI4Ql
tSZ3reBHDtD5Afs/ItrqfgVCf5nKwp1Wlgm2ghT/qt50RG+o7LAvlQ5K6XFFkhIe
+OvVl2zilC0LVtaqFJ/f1SPLO4fxQpRn1f1E+t29aj4BGiWb/E9wVem3usrysb3V
vtJjcUZU6PVIjDuUNR0kQLvWPIZLGaFILONu1eEI9pFbmHGAjKprZSC04Xb3brAk
z+pZhM+vrkhkQXmjCwyFmjOXaUryarDwqZqMYB0zR9jhHJRzcJYbnK+/402loRXu
CI/E5WmhnrqdUZvPqlUemTG07FNMfxT2623dXRBWdgNPlgJFN43N+gipxrvJwqVl
KKNiBV8Fkhjr/7m6m06HyxmmJD/aJbhhEuyIqOtg90u28duxfb6eoiWoE7KMfB3V
/6o4G1OwECzUbg4udxDD8/siAOzQmuY7IQb0c0Mht61JuMG2W+O38OHMChHmNa3P
xrbj832dqmkFmsYokI5FXWgDCCvz0ipEXmdwVavptQH+0YSRmLd2axUVLG35UVZu
QURGZlK/fCiwBiHB6zvEF+ogcFQnMNvLiz/dxvgVI/lEjpJ3vci9a0uSz7TZV2Lu
MXoz6fXZJdCiYVSRl67fvyEHKLM8Nkk55Fy6/OsSY8Pu13GNSIKsJG9+hFdFj4Iq
jbs3rUYia+ouRMnNuyTfxyhHE4adbFkK2hf1BPp5aMz/0OH+Hi5nx7ohy4z9tAKV
JqJHPDChHkQCNZM82tkZmcxnfw6CYX8DzJQZGhZepFhw/nYpvyX+Z95or+YNeL8z
72ecQdp8nBSU+XI7xV9pywvKxveOIO77KsrHcz6laOUPrJZ/ofFz7EYTpPnl5fnl
qjcUhROQUC95c1FaJy1uhMVUuFt3E0vFfaJS9SRdsCMxXQavyip8B8MDE9shES2r
9rmH8j2VJv86slUiYf9kQfp5q1KCRvrUL8lKRu/XXEN85+IgfHeUNg/pj7pMzcjp
YCJxAoMLVwvCVYPS3OXDlQV0jqoelVCVVpQX17YgNOrdQZVVgdAVHp7gAhpegOfH
KSOyyYCdYfVdD+IjHWlYpTtzXbyEKlisrpGKE522jZCaUwfZqp8g0D8/FZf8s7sX
3YunnKK1jva+SEtCIxyM5KEAuUriPlA/gW3FdjzyWjounVxm2AWKfkn7N6rBMS8A
VtRQ9+IGBW6a8QSgrtvmpOUb3cTkD7eq0haaJDW0ljt3td3jybj2bR9+1Hf0toII
M2C3kE0Tnqmxpt7RzGVx/rsL4DQKuZaRQ7fDq33KTBKRBVB482M/7GNQukLYRiLM
faVzw0bTu+usZPIZWhXDP2faME4auCZBO4clfH7NbztUkjh3HuMiqwOFWWDO1PjQ
qcnp1K9r19XAJs3r40de+hLO3ZXsXUHq/TILRVg7Ya638bBISh3f483abKv5RekS
sdb1D2BQ6wgX6bf6nZIg6SHnn7j/e+DPeWKGAsvI9owgG86DIR9EYyCtrW+CCKrr
fFwm5ifhDr9jvAHWThOtn8zMl2BxsI1Thnu1acMuRGvXTaU9KN3JsRKOyXw3fxd6
mSAZFNtpEpl04HGCZ1egu7AIZvSXr+TtMbK9hDHYXYqhkRBEJWbZ9JuBKNhEIHOi
cwQWphQFidKF78La3SIDefXVlp27qZejLaw+NM7uzna3TiCcgIDI9BsFhHx2onZI
eVd90Jf1kpN249ccpbLqdwCUEIui0gwOnOm9pC5aXIH+t/8/Kb02z185rWe9NOEW
HcRhswZsIOvXyQVUrJiaUDeeawaRpeYhcE32ybFae9sSXEoW9l1nzHxH9KMg16Ch
Fk8j2Y/V72+6JxFfsxjsm6vEbCxMeZKFUUZ+AEVv/yyvdWfE43aRgiD1vuWnfZfl
lgHPlezgLKVxAq/WlajiTrnTncQtYnyB9JEIWqvAhmLN+e76EcwI6eTsM5h+Mu4M
HAYcFleiYpDPrpurBVjAzfnAoipfghqcT94uxXPEZiutcrj+qZFFQL9lO5IEhZQ4
RRrdcr6qC9PIM/7bK3eWEIQQ68oNiroWV0zEq8hGERhAVJvGEDLUqWd77DTmwUzx
ENU6mu2qHuGEov2rARu8H29EDB65zTie5WqfkuH3gQfAQVLJwW1kGCnOwyLj8bzA
6gFKl3PEieYtFCh3pIJYBBoR+1B2TaKM8KGyDqskid5wJJKM9bE2ByFlYwmon8ZE
H/qz8Vl0GCrUkusDjWPQvvLVgz4akP31EOEa+kMew5xO165zKuIINGei01ypNqXZ
DsrR2+hGwdNYJjzKkXx6zzQjojNBrgSyBy2OMt+fOny8LBlr4Cv4oN0situfYBgk
qQE9XPGVKua4dQp0dbqTdRfTJMe1jhDkXoUeIVNn83Vi5WqElZpijXKOU/ikXH43
okuRHJGyLmUt4X1dCtNofznjhPibpzgzkLM+LEhVVXAn/HNKlpzSd9jPcVP39B8s
9OLtzs2GWnp+OgqF45wTOPQDNbb+3IjrqdKCO2bPphmubzdPDVZdn0VHd/7h17Ba
b+QO+eszJv5gGlcWy5snj4Gz1xNXZEt+yzPjWFlN5rBYwfLY4WM2trwgXrMXlP85
dsWf5QHUxO13J1oo+6t4nStltUgQZDgXg0htRCM59kdP45iLDUXR25zaqT3BE4Z3
EYb0Ym6IwFm19aJy6PhXIQXGwPj4lECCIFT1kOVU9iyEUhvF2ZLktXkYBegYwUQ+
nZbGNDuz2YHkJWiSndZahy4OcYn2Hp7zB3VCQ3TN8j0YteXuFMNPviVjVyJAlmGH
j5JNERk9/S0HiX6I5qUH8kq0CEaD2sEQVz7ZdOIzNyATYXX+UIQ+JDWD7a8r3gqS
CaGnha5cmPVEpKsLpftYX+U6Q1m9h5E2pAwl4Hj+Lvzo4tYqjH1vj6QncQSFwMyq
VLm7ncy1iFUYIIG+jc9/MqvJo+FtDpXrIngcWxf839VgfxgvbTVIK3Who0qtf+S5
w0J8B2lnmuQN/C3dlaDpz8HlQT1TYFeGQVmIthTZ+du7DoGr7+LgQemEBeC4l4J8
Wm0FrMkbqX9UUV83e8gY8baaeHJiMQVx78J6uPj7P7+wBykjfZdSTYZYpOa3oZ5L
WeSdnEcLi5WUkhtOrpWaMHKM0wfS5E8r0tu+5HD3qeZMEEcFO95dV+C/Pac5cM3T
Uznu6jqlHXoMNcOrzIO1yeQ69N1LjryNEnrhHt6R8ivInuNC0kFa6fGfNYd7ruWe
Plkja2Uc1qVLyW5KXdwbrN8KD5rRsPoisG1QQCaYvlu1/NCET0rBLDVCMbQlqLfp
Y8cGtWt6jtHfVu7jifgNHQc4qo7/I9aPt2ltYhBknubAvj2z8VQrjIcvUgBIWQCV
88ul9UuQAgukSrKSvuRdjeDOcrd2yAaQnzZ0r1pwCMsbFLXlczjSAbTCEUQoUlcz
lAad2lG5a2p+xjEWkVH5LxW84mmY4g6KoSSMs4Ei0/HVM6BnXwuxB0VdZ0HfRTa9
uMQfHmUeGqMz7CZ83NX/F7YXfJI7dmW5dqg1RdxOhfapR6IJf0E+3fAvHnM1SkCJ
gzJd7SxuhpRGKPJ6kRi6enDGOvK/mRPwyjWT/tTTbpxF+HV8/qTL0LAQz1F5saqA
SY1UAa7GVbuLLmVN3Wx4ByYcEKfvZzi3PAd1mdMxTZ2ShFFB2PQpiWXKRQ7tq1lT
5TT1xegUwRhx19dVQXIgHfOMFkn5nK/Elm1daaR1JYolaSY7KqLTV8NiepgH2T0D
fZ+5Rzqp1cTk3WwtqH2Tn04egqsbXOAyzamTWOQGrEa5q82QzOvjZ51/u/ZKwbQ+
/lGIb0r3eKqntYBZPnTp9ApiHvJTtPgGkvcyvM5EGq6Mf8LrZaQHmwicJLb4lkNW
XXKUTA18TAX2BDbe+UV5viR/r8Sxqhw+TjFuIN/p6oEjq30ResejO8ayAsNaEPPl
ehpj9dpYIxYqoI0PmiG9Set0Et12vJGnc2CDyAc2wmvt8GEP44CABiWd7NCK2/Gj
j4+uZLaIwNomVNso4/daGG0C0RavjgVtrYz4EDrEWMpqyH5QtgYBApeFqFXj7fov
pQiRLPAPX/DJ3c0csmh8q0M7uBc8NBuNWN4JpvZnByZS6MeWTlm5QtVyE3dkA98I
til+338LkbeZ1OrjsmpzAKWY4mSO16yHUTCsbQa+EU1PI5D3fPrV5nTW0n8GQ1Sj
ZERtd4hk7sq75x4y03d+MOzYOTo4TmwQCo0Bc2coGMJgJcZCZ6gpzZLrctKTw+YJ
eFYnr55C+4b8MZQ5C+qXCfi/u8mxlF4Qg1/ajQ0ne5ndN6xUkUiFCdKwGDHNuCFT
48BoNl5kgmd6IhkRgDsVB+Qu7oSSv+UH+Pbc4GR3pXMWmA/PrWm8mosYd7ELvDqv
bBhGi39FZD/HwvLxyYmz0hn6uaoXgGFpyXxYtYNADu0g5Jq3pQs4sQlPYZoVRGuQ
544B+kR/C+pijtvgQ5IlXzQ+IHKtdZAgHGSdqWLvdpme+YUV/Q/idiGDPQDMxZYT
q60PxFac9SjSdW6xoz635hz1kZOXfEG20BZE1cHegxlfami8uku3reHtgEr6FVo2
jjCHvYDEAaZrJY07SNS/8peQ9lk46GJxkPVXBh8lOiifZfdJ8iznbz2Sp/AzSXgz
gIV3irkwmvaqVVaA02S62HSMIywcbhywXG8c1t15GVGwFKpA1C+/ta7rUVqM3bQ3
SmanMlx75cuxxKkEBHeclbD4ScFndtv8vbzZbw+iS9vqzi9oPL+dOzVqTUXgQOrg
27T/mtrXb8+Eh7tuEVmpXOW0Nh7TNBodjKDVWWCz9JoeBXKGIBaoCTmlU0DqqGl0
nTk0tXv/dNasqzE5tbmHahM7JMHGOOglypDuhu+Eby6NVrmNIHc4SXFf7awowqgA
FaL89Kdz2Wb4Frvyt/kFIP2kHoithDiPNIf9IkGkoWPxUwRbvP0IfFSmoJbtjtQ/
xJSkQL7CgG6Pd0Nr1tI3gDPb+NNTacBarR7BOfP+bonRmRIQoWaxgCNCFoDW+xSU
yeDFpJLz+J9dJNUp5dUmFW/SXr9O9+KhFg2Cgv1OeV1Sux7RM7+8Q7wExaaNb785
ZXMaJp1hnv8zlWvLBl6LnMM/TcVEIDv0jbZbVaLRH7JuicJfAils+PoGpG5ZDn2n
JD4JR6Ca1ltKj6Q2tOcl+P1rz1RZFwUSwZTc9M5Hm5the+vQxbL25N+VD5hnb4vH
gtVeFB6GDD5y4M76vaS4hxN10KtqceugLQ1YVlF/Bevcy9Nknn9CTqt0jIEYzcz/
i2DZwF2JPz5pM7xJTj1aNL4AssCpzBEA/VzvCtvmL2tDIa9d/jGu9P8x8gXg9s9+
Pnwp0LukA7oKSb5pZuDDLMBqxQ9miJqAnogRejpFr7ZnLBkLXtlZ6jrVMeS5SkC6
q4UBHfXZTHYutqJrLVuFSRQXQ1h4V7BOHlAsBrHfMsU+O+D6ohJMUvd0ulr2aRo3
gQdb8e8KxxOvHwRzsx/v32HEEzfg7waurkX0H6Ay26hLLBf8qL7h3xPsVLFhtBR6
JFd2DWSdPehgMTYBpgqBa4c5Ov23qAX3D4iivIInjHSbtFDF6eYNzMYIY7L6Q6YZ
0vpzXL2aaZeClVzj8foEdmxj9vONCUid0lnhYaBq8WWTQ0v/d+QmNSpUUHUP5oyo
IRwdiOjDK0u22O3eMboPczyJZmrswRk6WJwi0iWgDktp+AzVnCmuXwSsIMkFnUSz
qwXjiSXsp8XEwqGyarWd4aWSKGpQUDKGbrpx8jEiAKezpkIc+gZTjtVwPyu1F6pY
qSb5RYuxk9LrxulIonOd0pbT8/f7npLXoiaL2p//jcjkViun4uMBkLtaAWN7sCnI
5la4Dv5wT5FX4ajXjOgEJYok880BgBepxUOTkOPPZKyr273nc2rwwu5h40nIruI9
dTbU2HMLFsu6smXC0jqHgYfvFZrh169nXKp3nTLXpi9y7PiVZ24KcRuxDat0F2cq
lYKm1IwLeSIjHWmWazbZ+QQP53QvBRD9cn/dQYpivmBtqG2FuUVcHFbl8KCHBavP
Inis0XUSljjoHMQjaGMGy03pruTOfyWClFD/AHg4bnaIGMXyq6zjbVedGUcHyVp8
5g3zsMcTbk6aeOYg5vP+0XLa7YfBMVE2R0Z/EBKvmvZnfQqz/LPjFJFRSkeUzmSE
Uv5G/mpCYuVp5AYpVqt8kOb3ctfJNF4iH0FZCKzItucv/IRDlF6dBCbifeQLkABG
Pi6zF1HD9T88g8ffFSKFD3Orbg+pnMbWpemFH7I/rAntcKMqbDok6Xa2YJzXpba7
AEGW3m8L1xhOrw+Fs0SnAWs17HZONWN8olVUCFXJKdtQtJkXDQdZQc0Dw5b0ea5o
UvaRDRmFG3/JH3Y8ZXEZI+lGH0UiUbf1a3RFop0A2AR0cXPM60EZ33pC40skgqee
8mWuAHBlQIYcpEaYA3stUBqwRi1doek/LpPZ80r5117mJe7CoB5Yqu5eclvSRiw0
nUPSo+THB6q95MJPm2RVLBGKxORv44NzrYIGBn2+jewczcPpwqXRyHR8DNeFcvtg
G+EVb4uueCWPxYpfD7F+F71k1kw/rUVJFiY969sqrexaxNJcOLy5dz9XgklVlZ9s
K50tHH+PAmz/TABTEVI8uSsf6xDkWA+GrouU5RTk2aIxItzTGdObIqy8dGqVALbr
LDHyAAvlB5cGmb4S62ItDc/Qmuplzf4XfGldv81NK99s1dsj8ncZmAsWxh3uBL5m
9rpoGxObpkCT8PavFQTSNyg5xhErTi041CpCB6FN4RgbCRD3wrK1/x/PV/53nSwi
m9PJOtKScHfcze1tVG6Uzz7MQ6yrH2HMbFO+8aNuZ05nM7ilBspUFmj4eERRPNRT
89op613vtqrJJ6kIhAbuK4IAnLVvUk8lKF/4JljTZwkkplhy1llrkGwMukPvfgD+
HFfU4Wl6fcxkTIvLsT7FVWRS63k4tmObO0PDx5N4CsFHVlHPS/8Qdeqq/JhMO7tn
FBDYhfoK2bguwSHGqTlbJfYchvNIL+0oEAvWaigodCUEOSUW9S1KytMiITk24B3m
9gNP0QXW/wOrssmrmyC+g3XaJkhKVap1blhIeDg2Eoy+okWGyHL1MNm7eHhdCp8a
i6wK2v+QriJNrRnN30iyCVrVcQfBkyKKQtttIFnxvxsg+b4QDqeSVh+Qgx8GizuH
sFO76Jk8cPXlYEdQuN68C4flQD1Nx6Gmve9iacXjfxTSFogDTblZXcj3hM4PhLu2
M4WC18oer678u/75u0uBKFQ/9CW1c+HFZDBTtyxthmZQgPllQoz5hLGLkL+HdMT4
15Bs7DhtdB/C9eiJF1eI7cs4cGBnVkAP9nckdKxJupLaOZ1iNDytJa9o1JFBknFf
I0Ss/L09pXOOJsLTMuLbCq7AWGiyT2M5L8IuEgzHCWK4KqF5rtmzP6DMwoHEWQkL
kUbL6aD/eVKNj5HZgjtc24f7mCMPRFAjnXOrvdnW18CFW94978p1YWpiMDzwTTvB
7U11ILTnDj27C7jiqytf6R2RHFOuKiM+2JaEKvbkBD7xv2N8L+6zjfWdBC3386tw
eN0qzlKS5X6yhlPGHnkS+OT3j2jn1f15F7hfWlgpQcN5SkCSPwH6g5mVpXWUdw/M
iHLh7mt7zy/lVBWCxZSC59D5Ar03a1thClv3qu/rN9mxcD+pY4f6si199KNRUGa9
E02JNtpt3XQ5w9jJvT+bKUtvG620S2cjukE5KOMnZYwhq8UphJDDfrjuIPN8eIVB
aTwTnOmMFNEt29FSCmjO5oc/q70k+lAXCCHjIxlJwFFr0NFtmeWXZDlhmhTYZDk1
EsHRAGwqLwqkjplV/G1AW+HM2aCU5mYVGs9rbEYP3MCRxfn5zRj/lsTdS7ZfnoGy
8HZTHDngJu/+5Y6cNOrS7Ql8RrLkLcDX7c3DHtXbLk/hI8qutNafwD9H1aE2WxE0
co4yh7WjvVpGbBlHgG446VePT8CuPUHvy8OZvirxozPuIIIzYMyM8OaFKTYolLyJ
9TcS227kmw4wNFWNT37XuiwFKTYeQqBBie+KKNUofBJu0RzmiY41d5pkDdiBcUj6
S8HSds/k0wbpSvk/KgDKKe/sUcRoURfFyTQOOGJeb9T0jVI/yevwpNMqLc4+YV6r
Azz/Rct6p/GxmqQLwuCxZR1u7c0za/IbqOOwv+9OwcsxcDDwiJaXbj5VUpcp8v37
8+aQAu2pHCjIKbR6oCitOEubG28+uQ3GqxSml9L/OfiS2/o7FgnqJF5kaTVmk485
ICAzJKs4xC3+Fxtp7B4LMm/BbEoG+UbNC0eiKKfG09PCOGtu8LlZilSS3/LhBaWy
bXbkzECk0pwha6kGPdGFyd7/b9Ts4+pmTOyr6bs25G0cEonXG7J/kNoGygO1N59Y
KjGLE605HyMTylnN0ks/aS7VEAyzQRQhjvAsHNJqaoizROHORoxMgXSxamS4JO8W
3gLk90NC7vHd61QzhYj1feVosRazU8n9GfDaFl3BedZEoJIu81rgxwLD1EOUCsvt
freHEDXKu8q5mT8kuq0vOSM90t7xlEfRnuHLzs4iChDfiqH3U8yAVC+ZkN0/n+13
Zxr0V/ycOrvFNQU4plzuWSHsOxpC5IaB85WiXYXoAhIoULq+F4sHsfushXW6rAw+
Bk62ffIcyXoinDiF2rrgYyos3870Cb3uyuiCoc1XtoMRi3HoP4xuP4UIXwrjHEuc
Gi2kklOAG+PiTiUi+7EjRjvH9q1w3k0PY0MfJVUqv/ThxSTOJhAm8g3SpWDeB276
nTliWzHsNGmO67IkrMxg/zWIPB5gDGTxSGZGxDgZoIwUKjdX7eaUVic7ZIg06cv3
48ePVlb7TDcC4j9QQFWCS1PSBr/RQPbEN+mozqAKfXrTNhHwRHOhIMBhTZq4qrNZ
Pza3MdEr9VDZVGGVRZR8f/Y7KfVsZfL5qpHcTCtz02P0JMyJSp5f+bSalFWy/fxz
di5MQZktrCCKn0sFPVpIJkbVs3PBlhZ9gawUru4yVvSgLsBDeqYLnRgnqAMeOxEg
nz3bJLq0ItK0BQGSpzsL5zJgM5e6hdbTcgT0gAb1NSKc/xecuTO09kX+ybaVCbKe
UbaBYRMEShsCeuVzsu2ZT9j4OfG55dtvZSaW7lH/H0bDBeHZgFI7Pk1Sd2l6nGGj
+Y2OEAK3gAS1sYReeqBEt+nBtajQAUT9dxThndK85LjeHBtL+hX1VXtSJLHhNZuE
scMtNQ5ahQGQtPuhXUtSmHT20Ha8o4S2ucpY+d/h33BWC0+GKNfyu+mqRwt8j/KR
DyA7bWmUtDB2uKXtVurVhdLqJ3vqRfgIo742fvQvLqRlrmmvsTlrfUCWZT7qS660
upE8LaP6HnP9XguI+4d4Kn0rvOKOL7QpjoF4d8UmwEbKjRB2Gahvp5n1mXfhF6wj
udVWvBtlUz0p6+L/geilinoTygVIJmHG2rVl6Cl83OIn7FaeocqkfZ0N1AEGhSrt
NECfqftBvzGzYThP6I/OGbbEo/Q31AT2n2stKv+2PkNbNBFo7uo6UMUAYWi+UU+h
8Y/ct3zQYllXvO2qM8ZZy1bGqqRbPI4jP1i4wiw91EdVSmk3+Cqwj34B8Apkb+4G
fyUCTyJH/HK3xuDZ7sc0ijQuWxtG+270/wpiThtGLdAQMhNhP661tcNlfkIhGFNZ
j5UyzfWdknigOaqBVgJkLdA+Fr7SMDA9Rq4t52FI+wnNyf9bOU3BcamZ4phL46Qr
7FFD5rticLkInH5XCxMuW251yCtpgrmJf/tkEl8xGIsqOerweWHS+PxPWDXbSlfa
XTr0czVEB4xWNcPfXZ2sEblw2TyLNCjwHJvXF4I7f9m7+HWGE2z3V6lqD1VjwdjI
5qRD2wuEMQVA51aq5MijCiD3eNrn3rlHa2fWlrnBpCI0cfYTA51ciTFHuw9v+d9y
jntJWi4gUKGI6GrsGzVbPmuy6yLic274fAhe2xH2jkB2g3yFwTRcNhlEfbf7rm9y
XQhs69gIaBV9TyR99L7kmWaab+ze7fIHj+UNQ9KJ22K6bN+l1pC1hybdxIrMT84f
4a3zHwU36JLJwqGD35l9XJpp2+ZwTbI31jYDoDvBggdyPJXAd16Sn5xH5rm5HNDQ
iPPCc72hy/t4FF/tr5yWNDsy2ATM3h1mbYxb/u/dUrmmpekhHY+ylEXSoYBGCTIr
ZXcCasZSZWvZnklxdJMnuK2ONjuT+8nRmhpg3F7n7ViChG/gdTh6BSbhdXQpq12C
nMx7LcHX29fbvMnY/uV7BEIG5V/o2Kseghbim1Y0C3+tQ75FgSDiD0oZaHTkT9nm
2zMUzfWEe0ajtsjKyZ64AxiQlmmV84DkiZFbpwLFtjUW4H7lCIu3mqF/DvsvMaFb
V1QK6vtTUFZQQINFfn0m8cCkdSj5+2isKZcBOc3+CFfNDSNfsh40g3LeKnkCVo8q
1iuZNx+dXaUxEIXJrYTOgcVYc8vz5R6vtpCZGYG9zo2nIFsdOa1TFgcQ5FUMwp95
+Po1AJdmJUOvSY6V4Kg4/wP133lU7UJPFL4sRfsEdoAo8WZRkS4zWsjeV9hD6Jko
I8y1+XniXIvuGExzOfIV5jYKQ3LT3oYTKMjejGwVtqOwLWzjKnNyyVMy5huBo08a
WiFWO0hZ3g0+NPwqljjXgPvpd84VPrWERMdgWzG9EYnBX2G+ZA79a+/3FvtSGJZa
gao4N6CJ0sLLa/l+/EVzpBSZeCihB+I6gHSvocAxh3BpgR+4LfjO1tRTz5nHgyfH
DdM/Vdti0isEm2D9nlPUihUx/SHCbGooH11GO+12gJuckQkKinrat+szK38k4LMQ
cTOPgsYJWU3ShAPE8i7IH5VVsUWwzGwiy/9WrcQOzAIGdIOjbcMhs4S5F94nFFcx
RGu9OhInFxJOopTnoflnrJNbdK7hVmVAMUkTNhy2c9firNlONgfJ4LaElr24ROP4
oOqRf71n2lVFT+NKD0gq95KHMLV2Ahdj29cjdVAU18idgI1VoSAKVTgvuMl9gsdR
O2f0vYPYkPs0Ia76BycNCvR0MIZ+USD1WTU7BF40hOmDbdHQ6KXPxP3Jx+yKCJ4a
YAdcEWBM0lvLqlA74nMvYTql/m1lCHJ1h+0S2J4SbDJTSLBElOMxp7LszKok5FYd
gsa7Tg1tY78CffiFW/UyVYmxozK+LfYpw5RPcLwmj4BFNRnJyywmhilHU3js692s
NjSWJiIBL/TjHDct1K1mClFkAhJKpv0X1M8IOD1ZNNM3805KgjIILEpQXqDQ7c41
f6XAsZSUmGoJ9VhQ7MBMjAvTo/MR9RKDYa1MW2rEygxlboLvQSZC9pVZiNxj1dfo
Pn1ReCT2tiNaFtSHv2KZZfAR5RUJw5cj31K7zyuOF7CWfBNQcCyMHUafyXeuQy2k
hr7VWb2n9RIe+rqJcn2V3LHeMuZ5yolPGcZC1n89jJF+G+p+kh7G0lcunZBS/O6i
ozJxp1StgUVp/avXlvB80fTYO8oS6x+z5KlKfIPKqUZcv17vBXarEg9QldZn/vDe
TlKxBpNC5D9U2HRHDefcEzoDN6M9xH1yS+omCeme31pRfMt2DSMH0TC1wcgkSho+
etOlMIQ5Rv+ImccyoEbNIT+j8PNfhvuIqPIWFKmMAqI8r4pweEExULX4SAtk7syQ
3rnRhkkgEMCC+Af4ZuzG5oc68QeUlN3d/jlTOnx5wJUAcyn65HlsA6814b2DttNs
6g3Yx9laYx3n7L9+Xok3Pf4U4PYd/rdoBOZ9vX3AEtQs1yU9ywxu/q9C7pwhdd3N
3+ZOc8CyA/xDenI2aD5Gr/o48EU2HzqAHkot6KgtAyinv8d5eljMRdOPgSgE9jdy
Ag9b7opqryWRFligqVCUr9PYXUJnMAZTY3RgSBUDRJpUDra8DMFr8kVnf1tO6hmN
lOSZececQdWBRLaf7PTMoe/rWxW15XNsSUCRvKF6+wmq2/gcqAco7U+iq5TzlEN7
ExZ/V0GnwlUpwlI/Io++ZBDDazLR9hL3iWKeQjzu6L7mGLGeoq9aynsifF8Zw3hN
HJPWIja+1cls4b2JHI59xgePRsyB9fUvDj/93W+PQp4lvyLMDHPxPDOD3ZlBFeTP
nP5QaVJ1fI5KLQJ3wMUKMpelR0aKRUUjgVBD10pznOaRkH45aCfHYDv88JWNzqE6
erc9Ow8rZrPOgJva5G3zRD1MxesWeYhmBXtJyKJnfka+7UW3uzYSJzi9bOxRo3oM
R1oj2uwZAHC7DpDWBiuWy6oKMski13zUwBYyJKf8FhZ8DNDYbNqSxVTOzKWHMR9U
Pw51+EkS20/fN8u8cji2GhZ/efnnj+jyQlsJLl/HDm2iMkhI2KN0V2AI44NyIV5h
l6ZrqiYI/D8TjDO4pz80ILzq/TadXdUJBJ+R4LnlX3HW3eyCor53pn+EzUE29r/J
uVNdxbidEA9I3YUKeg/51t+zh/aqeg7qli+flwddxhpNkvbEPdr1hqDyzDmPhYza
b/NfxxDTZcIy3beNm+Yjt+DwB0BZa7KkSmadxPpN9GeBEULkTFU2Wc7f6BA1br3M
lmTIEWMKIQ82NVBJKI7ADg5toV2LAI3BpRqzjrfRqv/35sKtMQmW9/EmyvQd+VeM
Srqt+bMfBMt/Wi7IoHBO7vrcOap5WQ2+sjFI9TTy3mK2Gq8b7WD5Q5CtsJzfbH6o
XufzqGXOVpLg2/N9xdK0hUKiqKZiDD46+zk8rSgdLvktJdxlgD5AnyHNOIUpKnMj
o84PVyxZoMUQxNEopRQo9lsGUOvEtauhDUIEqT923hBt4UUSjCyD0CWVhigINwLu
6xMg2Vv82rtZjvPvy6M345l5qzJNen7WSRkWVawNKe1zGn0Vf5a2AtwZlI/r15PL
uuwz/WbVnY3NE2PnWC+ZSxxVYo/bzvqayEIt+38FB4YYP+GnSZ3jOSYa5c5GnY4z
qshU+guUmr4wafkb2WEvLym0dDwrjVaxsNQSgB/lckpRTr4wRzrqdtP+O9+i1sJA
AJDPpQPHPu3dOQQKHIsqKQ6joYfO3z+tro69g571D708wqVYedC0zQmqGZX+s1e/
/lA1iOWFh4KVba0M92k51u0e5K6UymZNloD8fbuDS4wsQDIqIydsFgfZbRPUvgcC
Fvi7/CW4Y+YpZTkHoKt7b+w6PZj9qLqlij+g3c69XV01SGQ0sm3cOl3TjbACdxS5
ieMNCr83zMEc1O1awVThIZhKyfF7Z12LOg0h3Z2dXMrUC+CQkqIkJjFnB/8wN9y2
BnoX+We/KtqoSMf+396VPfXF60+PYEv6auEeKH2D3XAF25zvRFHXwZzuFIsWT1qc
5tTbDi1VW5a7yCdd0XeWCQQfXBrUq8V0eCt+9KSwnE1u2Ex5EeNrcX8eJfOrum++
HWzHZqbtUaTXyibGsGABlOf7e8OqQOlgq9YbtPjpIFyqtUj4Jpms8TXJgdbUekf9
jvzuK+9XrX/UWGvNcljD08fGlNKPXPcicqf6EIwt3+AwfYj+QtSdbePXlslwu6P/
BJIxhFs6wle7Z1EGYOK4A1v42+eiwTRzqnOmZmeVejXNs4lKsb1dolWImSfRWUrM
qJqA74Ot90u0zy29iQFXQxE8355CF+E/mmOolmhBW64GF5BhzpSxRQ5ORBVJ2b1m
dCXtHv3kbp3ZocxPcXiIxJhVhw1WvgyhgCWRsKTQM3L69bfVXdC7rcItkWU1TCGC
/4/1O6EmNEFvQKRDetvx5dMzmBm30wL3hunMXfN5HHnqKR4HKSxpPQq3Ty2VgdQz
GgKL7q3U8XdCPQ9xDH7BK7WUQoOzD2FTpOwqSTN5I4URvrJklNYT+q/pF9IpKMij
9KAUZ/5x+t+A6i7Ph1PuZ/Y3+28oXMo/UlqGALQF9Kri/RV216ilaVLItWejEAgY
1WXXcH91snvgNwPldIM7fLo4tOUbJScn6Io2oWwwdlwi5NnDP+j41CMZR/9YLP4Z
vvqJ25peKadSvdr+qv9/BUjImRCxdWtOerXrI8Hpp8i58YtQSxYv9p5PBkGcwFFx
xDAzmRbySRFOlPE+iBXUGnzccXYfMgtjZsrOIBP5Ttco5QYEbIKQj7gSAIrPbQo3
G2Z3d9VOSYMSPiW/j+J0qLPrur2PJsq4wMGEvA39VEKbfrBJ5Of4Tod6454hQIsF
dsCE4nMTshqwKsCa11tNLqjgHJA/FzL9m4QQqWxnNrlxt2ISUbP8de/Gcf46uAxU
OR+suu1bDE3quqJBSmpvyUnRdeEfpr/fHWbUgUgX6d+k+agH1xy/KiePSNG2NzYV
DYXm8mMbbtMiVIpG8cepKZ/KQITzPi2U/O7zwwtP3Pb3P2Tb3r2LEDbACbb621s4
nVDKJVCPRgbG1XYvU+j7RwXckgjvtrXbRYnbgcrROFaTKE/K2NFyPhbAx9LpTc7t
xlACd4TvCd06KGoAP0PLR3HcgZ8uQth98dX88ffcYJ5z8UEdn9EcO5wJjeH4bGTu
1k+NdbOcz7i2Rr1XX7oTOGm7UdKiMaFtGR83XlJdzC9ADuqd/gtUYaugm7rxRcju
f6KqzeLBw/GbwJcdPgZR0du4D9e7Gi/V5x/POutD3XESxlID7ZITUAu7bQ0Syc7S
ZLqYIkVokFjJ7+rNFvxrnL47qDpyAVlFzbKTU3oR0sy4uoeFNIa9NRVasrQe7NOX
CSv4P2EO2WWMp2rzbbXdPWybQM3mKpKcbQdqyWVh0SyfV/yc/27yXVmQwv0QyfD2
XcTwpsvDxLJbojv2w1csX0ceYAnxRE7PoGA4JzoWkzO27TmtvyIMD4F/kD2VFGGV
eqyYTOZNIFony8D1gUpEubMl1GvzAZrdnDD8cxUduls4YbpIzbN4eWPbIvCNP81q
Y+r0yw+tgkvf488KNroVG8eqLrmNFmjzjvJ9XsqmelLQytBu6cI/7zSNdhZg8rLF
bgsnkuHXPX/PMoDO51R0GmSQUHMTvs3OzdqeW5yGNSifibpODAz7KHY/mKI6/vWl
EOF20gYcP2BMgskHqAdzf9pYUPHeXEZqll1wBd7gcWr1J1Rg0LwQpOf6jRZnlKUz
4mkQSFkKdBViYJVxsF8pu13K5hS7dM/+9rxijilVgEKsd341oYre6Jv5ilxoaL8u
H+vdWueeSObticUMOomdohWxNGidLuzbs0CLBjj9KpQ5MmgHxTIisS+SDPuBLw//
sCVuJ+t8Vb2uzSjhXpTVI4oqNPTb5q7miymild2HvvY8Caw8ajszJIC5ufm25e7W
X+aDVDSJZ3kgs3GuaqwkzjKoBy3luxIXb4S6bpsA9jX2AU8whjntbNmnFElJPI64
duiueow/3Lqmh1p6xEK6mZZc+BeBDqbCuR2Dqoo9HAqaz+rQNObgV84Uk3Vn4o17
R44dQ/L1uJ5b91nWf+bumMGDLHz/JOaMyu4KYLNro/E7FY4Q25UaIt+q9ExNjtyK
MCsKcBesXEI43sZA6JfiDZn4PmKxW57O4XzRNdEutTsx1B1/cY2P8f2B0oZhV03C
RPgRGZzaCWutHZmC2PT+iLS0dwI2UCYXFK648tJSMTKQaILVnkOTZVRLnPHcXiGA
A5Iw4K9M4WB1+m4VLDC63oOOuHF2xiRfMGLMl9mdQzQiqef1VKOfgxlX03VTmIRC
B5Fqg5sN7SeZFd7AgOf0+nDlFuxNZmotxtFN6anCg8yQXxW9qEFWdAa4u35upODL
ubWs780wT6PySLaPq+1NGpIzTOQbxzAUoMMz39vb7UJI0RdI9LlKreZFFAb32KIF
3UPwVDONKsk7aS1iinDr5VD+mZivfDHciTYCf9kWIhAuEvhgSa4kSRURfvULK85O
892XWlyy3mZfVUBIzKgpWGbPyx78lEgqNAUSaRhZd0oI/S6f9r7pBxVoJNF8mLKs
fZ7MrT4Wl8UxxKCF0lLjzyqvuQxSQQCQ7kOcB/wtifieLCZl3XbsAGBwVFeo19cQ
hT2H/8lCxlb6ea9Qjho3XL4q+VD3qL9TElNPo3PHHsMh2q9jnP48ssmjXSKrciJy
DEU4ZZXuk2lTWEA2amE6NwAPiqn7f5fuUB+xfa7T9HcP8/6EZCj/U9fwjsFp8M49
9v9XgpjC7X0IpVHuyxMXnSLkPC0cet7O/S+j29XD0wykXM6KK2/7xDz2JzGQvHHM
t2CxCFA/Teh3YE6nvEKP4NmVtwxbVmuJyQU7h52JhN/R9UCAvxkq+Q+x1dwP9KPZ
hrwZmkJf5vdUWpiHcMF2R13SeoxqWCmXnede6VkPUSlhq6QM3eoPEFldI25n09He
AHg48NsOrgWOwzwgJG/MDt4gpBLyQW4IRNwOzf9tL7AyCcSfkS6ORwJ+TAEwjwxN
HGu1bG+OcHd9SD7ZNPnH9RXs7v3n+e94700/HRHGAu5ALP2W1d56BwFGAweziYtM
B5tuoXIrdSU2iqfD7ukKaTdBe8lAFmsLovgsYh/3TecIkoMcKdaW7KIf+oX90Db/
Rxl9tG+Fv7yh4ihul2wiZN8jSgyo3nDWg6EvRZge0SKWTmfrbp8s3Ml5fRgSXpTC
MBno7/Q+nNyHLa2rxpjZ8icxL/9PHNbdCAQtoKd/mRhsbdPGA/iFVIDP8qNHIk7d
n2S5byVpJYO+V8XsKSm0kH+MazuLTIph95/IiJZovRtXzev6B2EILpjZHD0RjMDp
7RW09gJIGC2k6FAslACnnRE+ipCmCQ9Yr6LQoBN4SG1/naj7EtGSJDhmeMkKEKqt
ri/5sgzikq3cxm59WlcnkSIHZrRqHGjoTh3aQzah2CAdZfWXu/h5hDqTGpdgLQHQ
g0TGShbsLPzEeEMmVQGZsgiy5xmvhLdEUoy24MPOt9r23tFP/XtafAGpiBMZhhZO
y6bALGJUA7eVYi/TnbHCdhkm9k9+HjMIquryuFKOk8sPNxJtqfJefmwpKnQBn/+R
uQ2clo7j0I+uk8V86SEkgeqodsBLPbqCM0PN0cprwYxFjonqw9WSEh0w9HSTiHq3
vYbOUXwqQ2j4Myu8A7cGklElfdexJ2nC+MAJKWHPge2bIc4uy5kFkkDuQK2WiVHh
yJ6ChYcj+eBu74oWsJW8XGHCe8Awv5aWcT9HEV6H0n0kroPstMLx7OH1NUwXncn1
Bse95VPPInoG5M1S5u3K1aWm8t+xHPbiEl3IRGMk0hg8LC88nBOWJjjaOsQAFL1+
r+bApKEWFpktovXeE/ey+7oq+np5PbmCQQXBzCamG71LMkoOEYuiBtzba+iB9aZ3
vfoLcsXTkEd81tNrX8fCwHYbTg58QH3mbEaM30PxnDnc7YdO9Y2kVvdBtPpD9x0Z
i6MM3glI6RmLs527f8kG3W+FrJVfe/DofrG7vViB+K4RZn4CAklem82RFkVEzOo2
5SGJ1PltmxHGyZx4tfSRIdjNLrcYKEsRfLSQV1nzbgVg9B/Uu7FLy6NT81NAvbxp
XxpeeyCTXEBv9gOQtV15ncw1F+Q0VtScsc6Qf0CLXvIcfh86kOhxfO74kxLv1tES
WmlDW1PhYbnYlesI69yFdQs+19+5RDfLdlC9/aM1D8mCP9IfDdY1G2L+nigyLOOd
+p6DEDoumd/5qW/+J3OAQuSUSAyFPCB3kqPWm/ipEYP/S08K/Em9QiYTPhuGGhUC
LGP0Bgbp9DIe0UdKbXZ1jtfcqKo4JwPpAVZRNoE3lBv0YQQ5rJp/s3oWLWqfKGM4
YQRwbKMBnXmnjCalIWIFlvndSR2h/FS4hWyf0/wSmp9Omr/+XjgEy+ji2SIw0kys
uRr4Oe/HD3NFHQzcKorqcZxow1ZckrngS3KaBerV/F+FponrpoGENp8vKzzGqTQn
Gg29UD46YR8mVr/ERuyuEs/QtOhkukaSXonb/NzYY0kaVFjTUQ8Uk0AuRKMgUSKm
MqlJz5lEPyayFcZzthGxVkx9xYkJYLQ/cpe0EbCDBVBwW5xc6Vf2z8+ldcB9nh8B
4ToJgx5SPgcMJCiFvHv+OAcp0HaxLmFEHhFoRC0x9VP+ebH9g+O+0ag0ism1K/7e
itXbDufQyj3QZ8ouZhFHidN61QW1mD3VMDjzD6K3paksqyP9FjIreqn+4hN171h/
nGllaCoZNRS9PN172axKE6zlYiBV0Vc2Xoa+7ntJuqbVHYzDPHVo30MT2/X3UtIE
lCx2mDHPaE2bq2TXzsNKl9ZC/Av6YaM8j55IIx0tyUNXFhd2uPGzKbfVOPhGQmnh
/Ah/Rx/8391t64s1y3b0hQjTt7lHSkRtURqpkrYcfmCU66ZPu/xgEy3IwnMHwMUV
ZcyrMs2KhxzRXh8HpAMChxJZReDRsZKrR/OzltUaWtxJ2G4xYhBrKqd6DydaXGnP
I+b2FwEjIdWwFYP9OgUnZSeM70AQDfCfyW8RnCXrZoSs4hG8Jq4hQmYyJPTHEQNX
a3eOQTDNj2d75ZA8NfkgeLFr86qw5fz7SRPcYDJwlslMuI7bkdGfRxs6HidtVV9J
/e8CuV39A/E8nldX6232ZzXyFQFDz7BJWXYtdhhAxE9WaoSjPIQgoTrhIbF0fXsJ
/DzbIkBd6wJkSCDZFPElkizJJ6epMy+dustM9lyvqDLnpZhQn3j8y4Y2w/ykl2KB
vqW3j2jx573s6yWzn2Wxr+bFNuhenTRG/0fk/V8HUr8LpOK3ldDCiAgqufmywVa2
AysUH6QktChEd/szBc44PVpYKwSIExv1P74IRs8iChW6d+4IDeWCKChm0Iw3eNyQ
+yvuwMVJn5Wyk07aTe1yiCEDii9LBFq7zoGLxo5etP6YKkRdwFY5OqK1KBYbwH29
KOHu1wO+odVSNn/RiFReLo4Sxu9ovP7s86XelwjbyyVNoDzb75Zd77MgnxphQZRw
PoqyV8Jmln/JrLTsiQFH0e9/nMFe+O7XrXZwlGyRgLE02rB1UU13OiswDTPT8sT8
L/e0YEC09bX4Wguwvoebw1qikzMSYJ53KpIf1PD5LxRs0ItHw8UvnO2tXyUSB+mn
wbYB47Lmn5UeYTN6gUPgq9dY1Q1Vx+XDqpbGycnGS3XmIu7fTV8g8muc2nM1Pikn
sawZQXGd8OxQsyTSoWYhIGRSrkClstc0xrPSwXWLkCoCCD1cgrncYgkwdjIPBd7J
jtXBRf9cGDkBFZzAiL264GqugtkH+OCryeOnUBtRvjUg7MJIRZIOvhz7EraUDNoD
g+e19uDa1yqWu16NLEaFxRvzwJYpElv8hp7d7EoUv6mgHll6vMPW9d7zG/2RWIRz
KLorLJHsMtxc4bINKJzqUlEMnlYfIckTOurKtmtGcu3XSOzghFQlIdYFxrVt36aY
WQuullQdbz84AblZyewuqIYPqlKpvtNrljXSB/dlu4v7JX6gY/fTz+xedeg3AX1+
d87zS5Oq7otpDcZ8Zh+zozLZ+a5fuG46Pld95y5uHJ/nBGUrXwRnua2byBBIXnpr
XE+AcNYAW/NotbU9YeRaJ2+/7FPg1S+bUl1vazhfmdCLazywLtVsJiZrBCwZpUSp
AeJuxQohgVcT+gjEW0vod//FMR7N9Y7Q6cTFmBZdLSN5rwRBkMQHuNXbtF/Uws9A
5bXaH/+P1VR9KTeSYOZuoGXuOMYf9yHvb4jhJ5h2dCaHUu1MeJCqam5TMyLBw5wf
crZsU2GBqJfrh0KIYtJmTM/tIr8u1mjRwCGbD1zM4IgzH1HynY5kAHpajDnefqyB
GHMV2AokigcJfp2gA0OToEeVcan1wTAGCo1pMtY/m6PRUZXUT929tCyE7hu/Yufi
5tp7+Fk1mQ31692JzfPaDlGkAfuYcEKhslgOU66NwLLKjZGjfJ8+OLRbU71qAJau
TQ/RZdO0NPANG860/MU6q5mmdt9ZelQWnkd6APcjCzGLH/ycEtxLhNy+Wv1Y75XY
zvkFedtnQopgF/TRQHv2oAkT5nmPvyiGCHXqb+YUca1EVjUvojalAtx/j3cguTCz
i9EYjyv15mQkl0WVssgyqqlGctPuBgcCGmgJdG9uJnRNf0QP6LD+M9PCNh+teHLp
hF4EviL2Xkee1FANa/3NjFmEYQRUSDx7TnEFTG0g9rP9k7G+P9KMqWcJ6dbFJGtZ
ATUfeyzAixYwBW2/LLVgEQs83+4uAnWxH0TJkR1GHaqB8eNuf2MNRVZQ6ahpErNG
YfI0iZZ/pqiqxC2Oi8AFUuc8Y3CZR+GTUkCUPuwwJVCagkt6FXHXqHwC5MEymJBE
1hF2a9+FhmzKP9PHeVtAPMERoEJ8kIjZ053TUPJ1V8DdG2k0EvsOfmgyFFVmixHA
itXHNpvwoLFYyMJa4HnwtYfXqDMyH2GraRSPuaJbXE1S0wdWvve/8g7WBCWk4GHb
uHFNO0nrWVOQDEV2yVDBq9QXiMnVvkCla85GeCvKK372uo2kua1BOf9kX6BXMjH5
LIgYpxKgznt7UH9UJx2c4sSh6du5EvwP52gPQiNV/Hg06prv90gFWRLVj0dMRIJn
eus7HjorYcSDEF4h+V2xX6LZEwFPuVNqcRSQtE/8HSC5CV/kB5nCokAJ9yBiwRnm
BeTxGuVk3KFLETrF623xNsVCnClfYEuYFxWIcL+gSyhrI6rMKtdGhL0RFciw3m3v
fKBiwakUokYVp7gFeNRvNrn9iE30CUgFGoF+ahGBl1P8wAm5wPX4/fLTkSH4KGjq
cbbZ18otu+cfx20pqd2vB0ERI95mrZAcslnXUinxcgllnoxiy5y1bc+7Gm4fXqD0
Z7onBpfHRi1xHSi1kF9QF5RM4sDvQTLsAHC8xzbTz6PnUDmZJyXbIKsf0GpYI9ns
0iBMKrDk4BDcvMC4klHT6a9+wjpVLjJt1WU86hyMrQd6uSNV05rUuMKlMyS2jfW0
TV0ssfS7tWVEcARl0ulIbm/gbrEGRoWbZKmSXyR2f7BXuDcArfndw6Qr/45e+5io
bHDIiAcYzHBfBKumKkNH3uRXYWn+xdH9jIU2nrLxpU2w9ihgWycPi9nNYvH5hxHB
LppZHAGs9MbF8QvSJRy1TGlPXtbx5jj3jSgj7tfI7COsVDgeXYIM1awSgMYKWfdc
qEr0YrPS/ZDGgEN5PTlYQWrQpCxcj+uhAIexIv+bAqJfutYXWBHf+mMmdg2AYBv4
d9Zlkj3GTtnZvKUVmmgKZlwLI781q7wDwprRU9sTgGnUSHgBQUEaDhjzwGrTtUUT
782wkikMP+vbCVBpwkNIL7cneSQ80I6mMQXO1siZ6igOzJPjqq5bCGokEQk5OAg3
YhzCvhMLMiOSuvXf5VnCK69QSAPcDWB000finjRiFaD2YxeZ/Z/gI7wgWmjUvbJA
BLcIyPuZE5XpL8nboac1AqaoPTBVCxCDPw0huPpW0bmj9G049SoRUmU9mr9bOS0L
4aNm9rC/sykH0I/u6kecxzQKEBgFXwLDKS95+UtLZMj5dqq24uGjz77xdHIeI8ad
zP4UY8yYx4qegtKfS3mWCHQOLr+vjb1MGA3n8UkKm3gZS/LqN9P1HbHJNn8f2g3s
/0SWMh6MHc5UVe1I1FwvzuWsZWvN2aKiAfCZg334Jtej2MjdQPN7n7dVZpUVD4Wi
VDLcOLRtoMG+FeznKth/0Sk3nfrfM3OAUrH4oJmQlqkrbh58pR12BCNdlTBz/Cr+
kM+d+OIXLmbQYIRWKifRvjvNdYXkjXcXqnB3Q2rRStbomt9fLkJp9T97g9kE1Kgc
80pJHuNWGPNDCNbvYt/ZSdPlSo6Ily4A8SfN+xjNaP/kNC5leSHlnJEBw6J2VmWK
yjj4SDmhKQZ2AjOi/FsBIe1PunETGNxuiiCYTzc1uJ4TnqqUdtMFRj6rz96JpLqM
Qdwca811VMVQk72ZxED4vzGIgzxX5MSncArPjpz992Mqxba89UnCA6t3pRbyOVbk
fuj1nbNhPgcihAk6U3WAi6561Pj70Ud9i3vBzI4LE0YgcMStFf6eLLNcoyQc14ub
YZ1RTRHbLRkLub4ck+0lHu1SW7fHgAi0EDw8w/AOTwHTFO1tHI64U9a38hCDjgDe
GOYBmjQCkVAkxPrp0SFThU9sUSzSNZb4dKGTrSbLbkIwYoQsGS8CWJVrEZryKaTI
dGYzmTaADWzWZQOOXGEvdMpf/gDi266qStceB/d4q9wcbR6GOaMOUrqSiMgK/ihw
P358HJVnpCeKOyiiNlNSDu8VJ16QofyspKC97Bet36WJTYiYxELV3c9TfFSzr/r2
Vloc/9JSfhYHNrC4DUOGlnpw0pQGulCpCGOIHxqu3ksXe2xzd1a9qmwQhRgdMIFp
zviYd1tlu6nheuZstRH8l3yOhL+q2l2NpmciWfJPFGBJgSwY9meWOGMKCkwFxTyX
4dsYqR/tSGUfgZwpV8l9bHB1X4KuxX1QqCcO7bE9E0bibU6MqCxf6WR/mrcUWvm9
MvlRo3acT/Giar6RBxyfAb3LlZZPeT3bERHnIispNPqrIf2xxtc6k+yAVK/ymffq
8cUV/FKVIalm7S4x4Gx0OBLVNWY9jLPW2YedhTeKL1Z3G6BPFVd/hQ/cVF+H/mUA
/EUfE0yXq4YayQLlqo76Gcf8ZYnjCD5TRA12X/Y8dndbRFjSdRzXFm/u57ByD2++
LKLs6Zwuie+qvh0G9ssGG35wXKXgT1qIA+73FYHCea7G88NYFgk/QZLaEpZyFexm
LCdKZ7CFvcrSjbphlvHFqWaffx4WmnVKimlyn5tSQ5Aahf9uAlNQ7ddrnQCpdSeN
vpwPFQZAIaqG8LmzNI4cYxAU/lqpKjsdI2w2a8WxCuJjd5i+umD7q49EE9JvEShV
Lzeydw656LXLjM1p4zx9nFWfP6W+N+fnSfv5qxqbkyFDLM5iAE8pR3KBsYXFKJZU
HA13eU34c0LIRuiyKAUKIsMa0Qjhtlh2sQk71g8W7qoNJS0zqqd8nC1flUDz/kwG
W07XecJpS72FadMPzFhDS7qv4xpLolc2dRuUwR1Ku6i4u+r2eZBee0NitlPZgjRJ
qTNDs0++01cMyS0cCg7pXAxOJYQTomZTOtrPKX+iffZJphGgbE+iJJX3wLGabQw+
oxjCmi1HMhV/QvaZt8kATd/NSnLXDE82eZiRxl3MXq9G5C0/kQrSQeM/53o3rSYG
u18yfQlvz6f4DXdg+h8cCsm93GcOSs6W8ap3gj51w7WNF5ZbdPv2iPj81hnOSlUo
AWrqgbmCTDLqF7mjGRJRkiDrWqG/qRgTvW5KNrpT6xwJZ0Yxyp16l5R8t/gnSv2Y
iWv7oK/h6r3UzLgUPb0mSaxkOzOG3chEZe8aBwG6Xw8XISq0/vfaRI5z5lHVNkfj
e2F/GwCa881dB9bjSNhPGZ3H3B0KECpFgQ9UOb+1EwkdfsA/xoABN5vUn+IaB9rg
LQAT+TTUduiGrmLmmTaxNcldUN1+Xfg9Aoxth+jIUODVf/VXOm/Wcn13TcAR51g5
MF93m/DXkiCRnuQxfLLNScd/yFoasY3KuGyppb9M2+/BviU7WRwCFMBtqJfR3rlb
sJhTEK3E/m30Edv9Vbo0p5QPGsWouXeDIatS/QyOvxdAWP8iBKMhIZQrm6uPi8RK
QREBGKrAG2t5qzvqb7Ez4YXVG51huLC4NttrPqmlZ+Ne92Stk22FHtWqPEmLqQnJ
3NjRKM2KC6fyP2tmtUi4X8Fj7RlhTVbog2GwWoG7t+0LWxzUvVPA97QDqezIp7w3
W5fGELj3fblWrzJ9a/Tcep7+QKiW6n4C9ercjsm4asx6ICiX5UL9wj0Z7ELLcApE
SlR4f2zMBnAChIhX6yHc1fFQoCKl8RF2z+0JkTBcjG4Udod7IVMZkqarKoVPXnAG
GIPN9WkrWJ3FKuxtBDIrR++8K7n0sQP2+zcD3MXR+LzaCLe0LdYmnMFvrYbpP5VE
Mduveae0YgBKSffsCWu1NfuwttIBLp5eebtNGCcRW0+HjYwYhGhXgGMcnXcdwfjp
hw5F9Kh+usfcx6dS9s+lvqP4nvgop4s/LEqkU8e8GhuEpMgsp0B6OCiIR26YhmLD
O+Ed7S1RU91Cu2l3B7H56DcroPF34ewPmUAWEAbCT/2E/7pvkJN+92MhDVbRKQhu
raJycamW7Lvty5XFeE3Tot4LB47O0+UOVaqM8n/jO9i2mIvlkUrJyuTg6iyxrC0O
tDvS+gRKk1U8y604o3a/SipDMPIknZI5rY+v0lm3OWFy2WPQM8o8/9OE5DgHNfG0
j2pIMHzgbQdoUvhcbZ7Dvkdg989E476OtJeM4DOaXXh5LmwaHyE3ZVZ+1rbjOtL3
drJpfItUDV+/DHfFUOoLiRuL3D5OyHrBTqz2E+h3xmmQIFOllQHuu5udEkKVPmPA
0w21y6pGUVAuoKddf7e9YJ4sdcDb4B4AuVDUKRers9eEsDOIgUs3iO6s1lWjVYV2
TWbKcK3ij0MrNeoVCYUHtTRlyItC0WPTjLimI7jB9Q2VgaKhc9akUj09HbJeFC4/
i9lJLlRVQh0tTyFIyFvy5FtQCk+4xU76KCIik3iuWXqP8JD4dExxiEI8NPTebM/9
DKwxCcbmRN+ov9Gpe9XqT7jjxM2g5pjF5yRa4YoRsPBVwKCDUbXu5wqyupSLdo1j
czCa7gTI8u9eZI9MuW/U/hIJMPaLVYbwNgG6LYUCrVj/aTgRxymDaQWMlFlGEEy+
gfz4n0KTZCv/CDx4ZJ/60IG3h6GiMPCUvhdEcb2CKXjZmSHn1esTdN7xw0wlUbfW
i+4JKfODyQ4CrAfbPe2coqzX0LcN+1x4U9u3jJbohwxG1o3MMKYaqwiORLAxPvRl
pVuF+shedgh7hlGARjNMvBnPPTgrbqmyrxzIiw9xLdL7dbLTjrNkiO0LezO4Yg1/
1P4lB2Vy6okkEotc2FnmbPyAORZ9skZqO7V+D0SOC9MN0WlP55Ow3RkWKvdEucux
9rM/n9U7XKYDv6GGeLgcaQB5UahyPjoFgGBRK+LtNPqkCG2j8vh6D5I58XTkcY92
mgYU41RVf/SKNVbj4NKNTF6nwryWnm3ZZycOL4oeA7x3p02RmVODpd6AaYSJg1Vm
rXK46HADzsS+vlmT7NjRYzAvtLpM56abCbx4/eU18kjnZF2CkJsT5GiXy7qFRLgc
PsTgkx3+lFb0l0ppUuTnnX5H64ErX7TQCT+CCeIqx99ERK5NLqvgZVrh3jEGygn9
LTF4KEggh5M3ADMJGHl0LbWFCKpsQrjTu6zvuB7zrSMFbg2pN5HRMsZEJ7c+yLrb
qHkkTP9ZdpRWX2urVloMx7ZIMH9B48RRvwdThg3hc45Wqgc/ot76rjsdy9yR8qHl
W7QaZB3I74EBo9y8D1uPdyIokeg0boX8iRiFSdabIcUxiBH31jfLqKGQlkOMg1f1
UomcSFLSpQyEO9oIjaO23+Rpnbpfdx969OpOZPXLFQBldllRmwL9SmfoqrH4vobm
EqXq9+ihAZc7xqOPtLYJk83RQD4ICGm0lBhH1gWniIVx/pOjWFU1kVBaf3VkoXGK
G5wVwTlWxiPAUD7BOUyCk6PWsF18EqDF4VGF+E7kC9QJLCiXs91W4+ypqjAyGMl4
KVCRsQ16T2YHqgpQiO91g0weqmzjaq+/duljJ7hmrwFqxu5UBbvUqhQifJEst752
J66uckOMSVQwBADX7dNQgt/SsnQWCtCrLd++uILSSMtTs2ePqfOvDCXmcvSwrIAY
BXG3GbAwm4ygYqzcgzx/2XPegKpqMxQRQ+dENTC1TjC3hZR3AIJ1+o1oJF69dmj5
FqOEZdNKhKhfcvirT0QxuckpkwuWJS5BHGBxOSG/9Nti5KdaO3FavF9+QbqWNsiX
LTIgmzEetZPcXQb96nU1zdPRaU5bDNPkUyGCxGObgDpq8FuDxEyHHqw8g9kmiIpj
ysebU9H2wKrH1smXTxWyL4BqUNhqvk7WBm17trCIud5/20QPS3SJEf9zwxRghvWu
wp4LPSpgnq8F5oLqNFl7bjDhvLkzpuXOx3jxBflU7pn9BKO9/W2Lak150qvl5v9P
iuUxDlOdrkv/e0kCer9RK0Dshafwy6cAvkfrxWhtkjZXx/1t6GwNiJb/6u21HW5Z
I5LZqfjoY/cH660Hml3mjfifo5wIz3JXDQnjRwFWjy0I+0HEFOUG/p0OctTp/uQm
8tvP4qr0PzsazXGfcAcjbpZlioKNsrM0lc/3tF8xxzYF5inoRmWrk3o3FAg5gmc5
5JimIrBEHLm18YOvwdnWIRbI49eVqOYVDoSRNOrbSi1+0yti+P9LL9LUCpq4D0QP
qdtFbFimELo8Cp/mAZ8FPGW18ZLrFhIzLTwg8bmW2rEuooWOwydYq665yH1PWKQk
YTHo9nZDieWM19vrvSOk48/yylluDBSHo4spNDTO8s8a+J1kCa5rfIeAW/0nYQhA
imgwc3yKbEPByBara2/BrP2Ft7baq0l1p9kQWdxk7ZqNO4KWGyeZr4tVB6gruzR/
fj05yaBrcWRvryy217Ce53893fZUwckrBfElOppuS561m6RSWCmRBDWLwgR7Hd4T
rgzpbYQx8ZN9aRk6VEbyvC2Tj3KfweryF1NL2PD7NmhpQoDyvI90wVYPdbW+y4Sb
AW6Ef4hOrpGKyy1Da+iUyuc7F0MdkkhMKF136YHxbL414F5b1/fSyQtgOLis3/37
GuZbxzRtvum5OHjmoHxAnikGu2wTCNi1nTFNOyuX+qKJ4gKb1ImCoAthK/5RkavA
Yn6CepNgSHLAZJV2oi1kms5UV2keongeLgTaaagT4CHb0jq3O2FGBzgsy1xEH6EW
gKh3WNrryNSXvMAIOcBV3OVXntx+y7kSrwCKgeCrlR5kIAFVjgWLTgNIy6Sfia7Z
4mOnui1H7/V0dylz4vudExs/NaVbflfCrg1p1MUrEPW1AfcEiFQRp4+BtiHHevbc
tzd788NgRL4Taw4+JZufWMKtd4TIm82gU/x1vzKuEfJn22Dznc3MmG6me89jlMhK
zZoNu5T8w5KqqpZ0Za52nzVkJzl/Whd0sVmDMlmkn/irns6E9sPhGeQY5hbDRN0l
9IAK+Jl1RVVbCO2pFBLNzl3hFvp3nkK9zDy0+gMyCJY12L/vDH8AgjMI7OFaRwJL
VVuPtPBmNDniWDVPYaU+zbU5akGj1fDScto/FfXsEP+Nzg5GN7DsafR6hYW71SVo
Unt/F6TngwISuig+QUhW1HH9I1wgruYlGAngN4RFHHEeVZz/XbLI9yaBp0ddfGKp
+Rd/LqVSZ/i+ohLQD5MNvsIJsTljAcsXhtRzvDPymz9RKrBonmN1jFu9/eGHQhU6
SClEUnbm63aCEWpTOY3eedGTbHIM3/CMbiiEMAwcvauNZ7QICpzQqnohTQHTpIWB
0FlNchx21JyRTrZJt7LsfUE6OCTaR97bTJwtnK85hzYlyvLyDeAFDIAdE66eO84F
c2OPiBA04Luv6e9UeYv51d87lCrsb7qnyLuu30c7omyYymhBMksX9qFAds6JYOSY
DT4y/OazZi7cjStwJJ3KNCfYadX7/1TCfJaFY6JIvv3jw+NYhrbv0GAS3jgnhoIs
4/sGTb9RU54ROOZrY2N2TSNwZ++Cs4hurhW+JkGDKnDlXSJg71FFULxGd9faMFvK
cAnH72RpoIJEVob9OmKjUYmO6CHYydAqQZ6jx9yedEOwAyibV0TEKEQDFA4yf3PG
wVZNFcSGQiHqmw4a6kmmhb+6XLoACeS5Sc1tiEnXYqIy/CfkplB1+419j9xMLo4K
agCF8jj5SU+hQa6/0KamDm3kPcHpcCFDNiIZGdbyyjBiH2O/4mjTAfGPZS0Q3rLH
mlRtLwY+4/SWLXsolGJ3W67L8D5yjHy8bxXhXP7+VqdJRDCQnjAQ5ThTQ3G4fnDr
utOooTv5qnTbiTlONePQXNr7OY/6n8JaqO0qrJk8PRXtZBtwKpJ25cryMGhm+sp6
I8IS6XzcLJrTLzx9DFZ8bf6/mZ90nxyMVZ8uGmvBKEi93ylywwEmg/9zpG/1KeIw
grQYOgX7wpRS1V+/JQEuss0zp/qaNpn1OqyCdTHdqmU/jYFqRcwGem4imRGzTNh0
7bZyoVl1G3b+bgntaYMq+fUPfG5KI3mStjSgdWAl6k1x/Vq+NSHFPNujKhSb7PUp
UCqib1ztotvXJ+V512k4CPnZbCA3vdKgi/Mqx/Ze9/DRSvi6WtE+tVmtXYBWZgPp
yApIcoaT2fiNtESIc/YkVDIuMROYg7maNREyer2SqdJ1AadxRGIzkYtG/sBBc9s3
i8cR8GwHEvLUYhi+NlUUZKn+Vdc9C4/rM8p8AJS38FgA7Cyo3FIFTwIPmKb8sHuh
1PK1zGWltVy/iUFro3zHbqvy6MiiqpRAMoZD0c/q/uWZ+lif15hRijfBK0fMXee7
mfDNbofxsiPCy8+RPo/Ebybi8CrEPCilmh3twhQWdT0Bif5DhZy7u72rPYnB27e+
ion0LJH0bMIPaqWCCJZbp9UGB1uC9VWFConpc5NYIXKqmDF9qVW4dB4dM0fsjy9G
AZuzSxS+76TUL5bMPbC828r6GcX9Fub2lp0Nqw5WWSwegXpi5buv1jtQj48nBG/B
Wm1snPpJnR2gBpalD4L+Jyp2jwkLMyTCy19aPcCmNtjxQJ/TqaeFlWO9tXqUybOM
5JLJtUs5JTOmjVcFDnr5drMgTZVbmkbSsXGigtHgk5CWAW5QFWVJkt3g15k6298i
P+vSXLLks2FRWdGCTt7coqRIZJ9kIrrTvSCAo5OJlXVhwb2nnDiXDtp1HzSQo7fE
dDQpBQPTIwZzCEcf7Gok6HcvZrBWt7i3QYqUrFb0HZ57jCsRoXyGBvxCpASaHcFH
02vT4g33FwN4NmEim9Gy0q9JOplc+w2ShkOKBUv97Jpx3pPWn8loqfF634A9r67W
5ixMUytKfGGTV7BVosY51qOvxtl5wv0H3CMhzaPnO2uZlVzVz2HVf+cKdxLO7W+I
q+LTvd7HubBa51q9qsLCaLex9vr5CNFE7H7AosLbC3ANHJ/BFjsgSs/5I7RjJZSa
VRPXhTUp3ezdaaPpV5oXi7Oktgvy9N5O6k+3X0YsOoVvyoIklcabfV8wivhDpfMb
Gy3whqgOPUDvG/iq0vxt0H9iSdeBNL1Rid6m0goCZs6Uz+mEu+ReanADdSHnnRRX
4dY1YejytFsKPFLRjpyZqnYPd+DKhk3pXI+uqBZlySgrGp+2F3AvnuUPImfGFiJF
+xc2kI2xjXzpzQaVSm2UTbRVt/sbOhZ5IxlMQ3wfbpj3FBdXcMn5Cwl8gi9GWHZN
ELXcn1xjDYCG8/bYlg3+nbHHzylD835/NjZNxdnguWx4OEib9J88GWX4YT7US27l
yx4YatpG6Cdx8TUJfxTXjO06DFvLgkF1+TYBNQw2IW++5V5OpAXITded8WsfZI3H
+o8h9K4QhF3w1ZR67ej7CBj7kmD7F9RK6TdPhMmBRRnx8xhMirSySF0mrPtttKKJ
MjTWeYqVfrPwLVNjXLkEAztqIbMeNstBhsU0a0aQMsbeVRZjrgG2mjEkz4Ojui/X
DNLrmjBxlzfUOlBilrEQAND7Y1D0C78oPKvl3hMGJgH3p+TTgVTwIYoYPc2RAJZP
4QKOkTzAbbBZuRAyiIAkDuorXx1AsFkXxEgTTLAGDB3+S46OkbtlQwT5QkqyWEYt
bgLj0ErYd+2Nz2ttKBEcZcsmPL4AIB1PABqla0K4Gc4Kd3U74qcLAlb0+srsuFTs
myWSL6j3OWH63nNSstA26KYRWJm+cW8v6qpJkTO384YtuLjDwyLl3UNLGkJOF1bB
LXVIqFN0dqGwwYMy+PvP9DKhdl7sQcb/ZDLYWdPbmRh6MwemuGk5mEFVDxMPHWCz
bDR+17ikLJkesf/eGZhxoQ/geqdmQnq4pzJNhmMa+ZxCwDzJ6LcxsQMV5RTQvjJX
zyoeBZHCcboklwKJWLd8NX0XLunf6yihcqY+e+BXLV6gNK4i21XGP9jFWbSviuOE
wSHC5xBFLt87ujDdHWWNfQP9m4IMq+BxNzdiYsr8bAP8XBIQCtDTGMlo4EKAAIR8
xabl6HsBzwMFLaZnb8ElWkKL8/NUmlO7U5N0p6BxaN6I9jH+/GsBTvenCwG5Sbw1
wZIoDMeG8BV6Kz4x+W7lLskqsHaRd0tCAnGMHhZMdI8aPUm4pXVO+BXsZZ3np7ID
MU9Z6OiMZEP5o+s51MAQLGVw/UeT1otlUN1bScloxqBxGzTPI6s4a0JQxxRcwGY6
iaqWYX34WkyoyGFeeBj07WBgboIJ2Is9/B2cPCK1qND3bylm7Fm3LAFBoCuRL5of
WQO4/qb0qn+MgetDM11cIE95qY4tBvv56NxGx6jGgxU6G4sX0vQ1/HJ4MAiFAOOx
f0f6qwPvvtecCwqTKAh9dToyhk7I1wjnHmp4bx9UUQzOOr5m5K+cWZDDulZo5WqO
HETFo5Xg6lgnd7Kt+Oe3yrKEL5OHSfPsHfm78c1quvguW68V00vo0E8Rak8WknjL
/kgyMubFEdMIKsHmOtgxjMrIoca+Cae0TepkzvQ+MyDI7nS/zwL3DmkrFb5YAEML
F2m9mbdJbHowXueQUIjAiLLYLg/oI/nCI4o/zxdBffn4tm265H3eYBO9FXOiyKdv
E9tZAcDnqdwemT1oahAxNWaMgQefOgb3s93jNmtaZXXqHY8bQU2OcoGD0sI0QMOz
eS82PuHuxDtDOpoSUAZCACXsIUeHfYlnNXsa6y2xxAZ+j7Xn5aDtW/Bgvq3CW+L0
bn5TnTahUk3hkA4RiOgECCS9+YmqJflHARTFD2RuXCgbX8iy4JaH0i7vwapccc8G
aPUR7XN8xgPNFzfcUyIlh8ZpXzmt4O2PL+EJg5X4L4PaE4TG9Qqt2yYZ3ROSwajY
6ak4+VnilOdfNrU7GxvvZKvo7Uw2Rf/FxKrjkCo5gA2qpmDo5L0gPS5SSlHtEqJ/
PQ7F0UOmVN/ZL+JcyxMZh7KybfiM0857LcIunDo0z8AY/GttF18MzOSiQlmfhvZj
xaNF04vaSpet9ctQ44mB5+ktKpzBT+pzoU1FVU5FP5gfcpH9VTHdQ3Sgq84m8XLw
3gRRbHkqUQD3zmSxEDG0mMXjDgm/wO1G/MCRcedHJhEh7rTpCzyaJHYbKf4wYb4z
dqH2hNqbS0dqln24ys/9WOUgNyCilbQcxSBZAqcmlWVtNg7OEPgfilH8WDo6U5K7
iSbMEoWGVerL4eXpu6eotYHmQ3hcIPvQQZRBwbzK8eYhTB4JcwqRB7b62HBxqf4q
857fywtHdy1Lc3GKqTd16W4+jo1BtX2O5N/DWrcSFRNyYbrjj+/op7/vC1u/4xHL
v65CqrdnOs5aSBfJ87f0tmyM9N3yQKe+aiudQ98AgLTJKNRkNzRqxfG0A4iXDb2U
addFgqIjzpC1BzBCzBJr7ZicXzlyXH7ewOLrE8mTa44hr79KlWw7J2LzDn/nn3tS
zj1hpr5w2Aoxmsvl2WOaJOz1NcT2m8RO/1T4+Nmfdo1ONHtYPkD2Dx9nrrwaBq38
MlMchV79kH0po8HL9J2St1NwKVYFheafAev3RHegipd+syv0iO4lOAgrxW9sH67c
DQSuMETqiAMXA0bZIF5U1QBcqb2K5aSVoFYQ3uGchKQjeKByZJN2Pjv5g3FSakmL
Qq9k9H0tePsIIQnxJ/VWlZnsb2ta1G+2ThyPWbqyVxX8M+kYMSqPuBCNApSzFxcF
SHSnwgq1GH6yWBJFNRt+ndNuRSeypNwgX22paIuwp5hjYpGP6pUIpesqFFtiyzsR
dQOt75ZLjVvm0NvyIjp8laWREadSA0s8v7xSQXZbR/AN3gdfJLs1rpi7HhOizlvU
9+tL202I0OrLeuybunH9YFdQ0TgboIXEYvZDuUVGLLB90DtFdJKwTCqrSNn34XQu
vHexQp99KV6aQKoPREiWfG+w+KsrieK2Bu+DyKokDW1bhAwWZUK5TB/CE0ZSE9Mq
sZjeCxKmobGvNPUui/i5pGlXSZeQfjk/YjSchR7F2uKqd8yD/eybo2yq6vTgrHRT
bzvxGQsupqU6tA935dvElHVZA8YvZndDysS4HP4BSBpYKH2H+GQ54MiPgywPQQHa
XTUURq+s8hUkax3fjBWszPPZKzxbH2UXeBz3GnqO7qwY9aNY7hN1mJMGpHJw8JfM
S6N6/yoYVJXsdiGreX4DZsfd032qljQBLq+FrlcWCqhIgkXHmvys2Mqa0W6VZzM/
jtlbYMWIwjVtXhht/UVtQJXRuxBpC+qr86QwYQ9RCbfBa50ERNQyXDVvp0Lpafin
xLUecZE0hL7770uMVFGtQSJrtJTkznbBMwB0cW+Rc8opb9+Zm7nD1L0/AAENxEqE
1zo1JpxM0dt/OG4gbuqAYpkn/uUsDga3fClJk7HqZHdb5eBPC8DzhTMT0hCe42HK
f1Vsq4m3co5eo7dRnpFWSZKDen6mjAfni9lABThZsqM7xcCF95Vyo95f2CrkMUun
mkK5DvWus0yxhhYKmNqVC8KB4Lp1qbWTLF5+IUOCRgGqw4nZy7Vgo2UIBuPW5yyu
SwNZUZMVZ12O5z4qCXq2pL0vNCkaijj89Q6/dybaBB3whiO3gYEeQx02IK+t3P0a
2Fdi2a7QtSxHmJ9VdLxpN+QLeJD66Ea8nBZspbHOfmFjTQ22wE2ujxTSL8xjljNh
61MM5SugmmJBeetYazGSdpnu18h7F6UPRysw5wsc3Ka85wMG+7Qo39aiANE1X/7u
zyIYnl2YVq3d/ofYEWk0nniZC0q9XYzK+TsTy4HBk/luOsLwgGfkWPW+1W5mMTLY
0rje5Mi/vwgsoPxvb97qn3Y0Zg66sNhj0b8nwurmMtqu2y7rIHw+zCWJHYMPtaQj
w1RL1ias4eL6tD9zbJ5LW+t5Vq/qwAALociPt3inRcSIxYl41Vx4/Lp+yQl+tIrM
weRHrYEE2WNd7CHFRZq7X4AbzF7qMHdgHo2xBJBUO0bCH70IC8XemGIsSSBaY2zi
82wwyiwgcdSUJkfcM2EYymaCjgR4yAJhuEZcu4GXLEZMyhJCY8hrO8gxQRglTkaz
Fg1esYt+MaKavn2m85KfMJwWELDrPI63t2LXZG/GUcbJ4C+oPMe5T6IhfXKr8vBA
LTpx2iTghmhyIk+XOHeWqW8uBwm1Mq8SpLrs2HkiJ0PdQJAsTVYThRFESBpO1rth
ZEr4DkGHsLWSe6phGtvJkDPt/D90WgnjiJnjY4NRozK+ME2TITsYz405N8TzXHYZ
CBXlXQxhLpI7Req6anHUPwBlh/+LY8iIN0wt1gNDi95/mi1uhRAKW2CX2XvwjXSb
kQklbHKkR1itKiZ1y30fYFf93WXYpzbWW6shdnm+DD52Oq+dFXZtz/1qkqORyWf5
57jA5yXsriGntX89KmU0yZfbN7FlPq1Uvqlz+trYWeWcLmGfpcJvI0jKWftaze3B
1KHR00zXehwIMoVnn5kpdA/+yoq49ksWOKnbhgeP2di0t4m2X2WVRpzydd9jqyb5
fESrPn5ja1c5RCCvAXevoEj4vOrqsql3cjRUpPW8j+6+P5jGcmXlP03Zg5PT8+bV
HHu69SwM8PYilr7g4VGkNn+jVB9aVMDpZFjZ30ZM1CAkmGxX/0HkQRI9SMlnFnEx
IGiVQtxEW1ZzphPtSwKTbRBpQfKtiRtE7rBW2euFi0SyoANTqWGaihU3fPXzqAeC
x5Xqzk6dNTwW/H2h3nN0jOJJZO3Z8YXERDBmKSkRpNN9QqjKXZNPecZ3g8Wzpy5W
md4AvxvjK+HoDyXwcz0ejWCUjsoiDJ8y3I7GU6k5GxRpfZ8dt5J9ATlVWfnzUJ4G
V6EEvjGRfxqUlmNTihQ8F/rjC36JJAJiLjQ6LZyPbsI1unsrUvqj8QWusZC8E1jX
BCPphUZ6Bke7kKMgEsY0Vza1GiRMPnhkh8LKCwmy2rp7RQr/0qtXVL4+bnxJW7OL
mN5KqSjYPG1LjhYgu/fkQs2MdcR0X0vaJNft+aEFIpOPOqCS+OhET1lNC3P4YPuk
tszJI09q3rhVDsKiUtKx+EkhqZIeXakUiYAXXKdXPF9TvqVL5znAqDI40RXbKE1I
AplxkXGkDjp9hyKd71oh5kTTq6/KVBmJF5sFZngPYmFVWIHWPAGRdMYCZq4mut9c
5pAtOQ2YXKUireCCcnbuHJwaBW5j08IaLX6qPQRzMoO8aXkPDDuJYQ/FIhL8C88w
Bo0TOVSI2fQlHbsMXU6udMlsNh30xB3zr0DHm29ihTIOxyrGeUDUqOqGbxmLqJhc
+isPHm9/NN+ztysc/lCRNLDFe6FQJjEy+pmHTyOI5Xwq/BhzuqkOK64j6Umcfvi0
OxSDJb+cKnrmqgEMuniZLOyVLt8Ydl9l7V302nNm23RX9ShmQp+46jIGdRB4sMmj
7Xja+3kJG8XpXhwhEUl5LTlFawSAz+ENNBM8YgvvhXLnFcLSD0MApQjGujtJuSEu
M57eDSPmX91Id8gOtJhJQsZgx5qtK/2CLMmOPBhtc56TURpS2YGQgoa+nUNXxJII
/LLb8Q/GJn18a5r6Urn88EZmky4SS0/2yRqtiGABsxlQeaIqvi8WSG9EXb0sLZX2
SdzX+HhDD6hkFb0uONXfV5zA42hbqdH982IS9DxYG6P4ijWo73gT0MsSJxq6qf/O
0S9r9X4bYybcquQXkW6Aa0S++fLTeLn81A33aYZcmejfg9ei/+fR6eIMpZyoh/9z
bqJwMUYkGgfo+dmUP/vbUY8iF4j25FtORSr121egqfPfTu3p3DQPz7RuX8c5CwRX
VT6vHtRjWGVH+e4J5Y+pq85eptP+X9Vke+bIx+snxWkpRozhrDZa0bi0coZa2QSm
ktvinZ3zz1IP4kg72Cgu+S12pK6ni303kXlhxelJTuCu9ePBwhKeJ2xGwx8vwdK9
6BIm6Bq2kjxzEgx+fSkciSGrJqk7fDmAePBsVvYglhPbiYI6Es/iO0pILmsimgii
bQVP7a+g4U9nsJI80Wi9JWUlevKMHPy6lTTka9i0hs5GSkXXT1L5EkoWyfDdQt/J
9+baTRZpD24cWqajU4NwmbK3KFw812gr5rqZMOu0niFE4IblWpppKHXnsEoD4kB/
TjPQuXgFCA2Fr81ONcVV2Y2lZXIl9Qepalc+BazD1NKoPSmcdhRbxE8bTthRQBlp
Apox2j/yZcyBeeDMK9cxYOK+a8O50EiuIisspSAe3n83BSCUQAbQrGDU80XLGO9d
xRjWOFjxk2K4uNbYVuIDCbJJYbzs22eWj0qscwRZQG8omDStN6xvyEk916fWfzB9
ntsKPra4Qu+LE94IEGciQLRaPnRTURp/7GE4TWXKWgTsdkF+Y5eYsnVcpNk1r9Ys
cXEgGXOV5xgsS8lyiqJ1T26Oulf0UB7rFC11tR5mVCwxpru2+P2bfJoRoJoP2pKy
HrfMQ/6yO2I0NKQcOJvFhVt6uKYuLoiMcPv8CQ0EsZYP+cjbdeZV0rSBkSco1Ye+
tZk02MUkGEy9BwQP4NihcAq7o8M9Fqj8+qorn8WbLZo3dwMIR2pHKAlJRB6CvKd9
hf/iatmpLOof6cjohri8g+weUWjaXF2xwVAh9FzEV0qUpCimVCUw3xvCJCw6SWGV
EgWJCYkywFDpORbSgIUroidlOnSCf3steKAXmhSUHDAI+qiwdzNl+l4qt5NBEttc
iuRitv4IOp7MZtX0TsGniuCljwVjt86PzBB9h+GcdMcntOr2DtSWt6qS0yyRxWZQ
AZ55BtkiT7pIrQbUa+IPqLDMF+S+7zOfAdxVZX+UHcgSey2tZfF/kI/s1E6ELXrj
RE04TGRT3THpwvywGdTD0DzHEtkIP+XUH3vHwBKFcv58FIobwFN5t0MxVpQFWjYi
8hhebur9FFqQgGK3FHq4Z62g1/vllCZxn4V1M2sjnGS7/4I5iwJsSGib6ArzH0tn
WL0TzINJ9E49/1r9U6nIG/+MRupfqHE1Wa4R4/wV6g84TS8Nb83Oz9qnkAXJwNae
0q0/sja8hgdngwIQIbgCSYwSLr+4Kcyxkaa7gw9gkZZnEBWxt6hJiKhKo/1lYTZA
zUQPT8diXDED24WQYPlcPy3jr7+Qxkvdj3zamp2k94eYCS6KbvxaNSOUSE8OwEUH
+kEQA4CbCoWRc84HQ4m28H3M32jWIPAsYbAolebwAFnDk9RuZ0PfRM86dgh+D+qB
6mVymW2+G8kKIY+l+hnQRUVMBgDwqhLznyVhX4MAx132EqvRr9xUUfnbihJAfIWS
0uhjLyLMRRIHAseGbZ8q2OLSyXooibYhBMUtaFtmQmFrLoFQlFyDDIiWp5RNJ1h6
2vsw4QmLo4zuaRUOUIP+mgBSITuwqWZCN8ZchjXnu6jWv8gjxu8uxLNrXX7K55sL
kSMiBzaG52maeBGBeq6vqq1ydgsAA36y4bMI9fnKTBaGtyQXV9rWqnQ7Jj5R7Lea
HwxbTv4rInk1ANt8C8Z5tt7C0tmyo7xGEeAGHB2fA3VTAQQ6CanFW07mJ7DbKUUS
O+GYEvxZFZM/AJxwsFjHxtQgMx3zMAtsD+Vmt5c/dxmQjR6QoRSzndh/2S0mkMcR
vz/2Vhfni6bMyRdjgk5b+im9hY12lb1N9w094gFdV44aKirjUlUZcRJqvm2BpXEx
CWvZ/pYX+FQ7jVh7IrTazAuXgKWbHsxCkmLxSi2GT1xGJsYa8KeTHCr0DzRqnwKk
3Wr03o0kaM8aEmR4A8e7FBilkWrM5IZcGycI6xwD+FTAaHIXPiL/qjQ/NAbamUH2
kTWlLQg2KP9/vsq0nBhIJkCHOdSbYwyODvkiQK3ZYvpP41P5dDvtttuCbZ7zLecS
pZnMdKKjS8h5o+kHf4lO9OJ0L1241+mkVxDZgM0LzTUeM1asFGph3IA+VvJDjWaL
8vWCVxcadFQ1aSQM2PJHTbPucsF4mSNd84HPQGrL1Nb/q5CNgnUx9tpALYNXEvmR
VFsqMHFFG4J23skSeOLKKYP5x8FEn450glQFX/WNUj4a6kuYI2+Wvkhp4HBzk95h
zBmNYAWL1yXfGtZxwaB8MgoYRa9hWhn93av78rfcdRKZzUXusC3wgODsAm9Af5jM
EKK9Ca2g5O1iuuUZqf9AKwysOsKwVLE+oSKgJjERT10LBAghBr9SPQ/bN9wdFOs/
/YbbsILNqyipXKV5oZKnRfKdqBdGq103LMAfHetSUOEJsuoN03CkTepu4tLf52LU
AJu72WmjlQfO1wui5jVg/ipRhZSwJ/EkIzUUdQlL/QZzCOED+gXo82/Zgduph+1e
SiRzJtzz61w+aLlSUzY1V/tIgqB89lnWL0zhU1qe+7VvhGl00AMRJVZqzYnfezeq
s71aydmKxO937trzbvg63etXpyRM5gt9ykQ2KRkh3+i8jS7Zxmw4+FPmCBUaqWQl
vle4B2JAET7Ofba66Wt47OF8vL0Rc/8qCSALobCFKZ/D2TTm1l5KHXfovpxSkab3
vcuwGQFLY2q/CNM4OKGC9H+tmf9mygClkhVEY2Zr2kWeVxY2DVJbSFhiUQxSKiAP
0RQXRDTaCJHLkBCuwQlIBR0GdpIU2L3ARNZ/0yd+AFPhDS6mFyxnu4lUYl2lMGoB
AlB60GervUCrarDuuQPI+UWTpArlhtN6K3OIqTlK99Grs8j9Et7r/7B01Gl48UCV
nnq0NF5XJmh0hvedWLSZBJtv5/X/JAxCtxvZQZAhnbnwwUqEqldbhAlLgoVoje+S
bviOszYyH6OISMeSOc4hv/yZomTNmmhGWjR/rUHSU5mTXpaHFbjHItCFcADLULuS
jwJ2l8hnAik2psyL90YlTG7BCuDStbMsotYq6guhwW0RzvP7xXEil9QAnRAYoPuX
fh0qu83+daN6xSXovHBLHuY048UDiYNGSdK8yk/EWVJjxt9zOO4bszD3KFuzKpV4
wSt6ctNhDZoowrBhWxCLHkbcMEjrFAfaqzgERzjd7PMJCvyr5Kw+34sWlw3/iiLp
bBjRgUQqkJVf6gvnBNq2+I/tLSpJKE1iu8OGQX2KQKhmEhogZvJIMo4VcXdjlKob
HZUiDKT+8BqJo1Nlok8tl/uUPxZTB5AF82VJXUs+Dcb43xUn89GqEnpXzg5RD1bv
ANMpnI2uBk4t3OThvwHH4ATEVd6ujDejDXPQAN5ic18H8rfAQCy6RYVzzNxbtNo2
YThSaVKTwOFi5vtHzNZCIp46PCS7YtlAHky7tLRi+aa85RMbELfJcaJ7YNuAnBbj
DyoVT0VL7N7dlNtcALJjt6VmVqyOpagViYWDu/ohNIBg7iHZFQlYUnL8DljaTyU5
MH9Zx+vDOv/V6VQYl5DmcNFCLl8aFr3Q4fGNRxfb+XmmiVkcunWvn/lgSuZ54kBv
pMpRAJl5cadnF2NZV2Ts/DhnK0zEWeIOjekXZ/bjdNDI43vguBKq0NXYNv0nnZuZ
ZS0OkByW4yloa3GsIFbB207/UoeVcXlG0SdjGnd547xMpSXz9hs2pK4YVNNc4w16
DV84/bY1zj1FYo/9y9FnkZsJAJjhpE/j96lPVlUZY1XaD3DMyCpKk9KPVfAcJsiU
zPf3ItsNirbGaUPQEBdykenWePSQUAxU+RTp9GcLGlP96RVw9rqZoNSgESATALkN
9898X/lhjtqPIkWN6Msmhs3Y4iGvYnVEmLNHwsc/+lfQObXbzURWUqKrgmby02sX
qlQE7a5CdK7zmwQzH+f0h2ftSz+vZ9kVQR5q0iD3i/MfoJPb1WQxxIUKRAZ4R4dr
MzUjRIgBFjwnDbm69/Qf34l0MHcj60BKU6Al3IwAKRRL7WP36+C74At5A7K+2pr4
Be5MVYB+jwTdnlnwUI4woI3FIFGPbxyi65NzSeUb4zkSNnPS3uibzWFN8ox4Rdgm
/b2tGOnCf91OkxJyhsbSAIVdTAjBsq8EKGyOrn+WlaitKxnG1l2Q7YHDBY182tCL
mubXL6/vd0loYNtIpg7HKJ5dKuKSBqVP8MkyFnIHGUATPUmIFG1soQlQPkpvuqLL
csZd18ags0QXsT02ArpFih0Edt0X1PIDJSGkxnyB4v5r6Uo24AdZxVAKTntw+XkL
F8XIfwd5liKiPrlDfRh6IAqBjbFWqJTtUOb8R/7Wvrg1OYrBAuOoPY03z01PswTF
LvN5ldPDpO0CS3GASWZ4KwVXcwKbksX7DetwnWJwzACbJ0f6pYEIrPVGzkxbVxih
OpBFvfMpLzqiSM9Wpx4RbajXsm/1WGCzNx0eJYoRl5Pdj0f1MG1HiMb/dHj4KcRx
9iIuBnZgjym8HNGtZNJSg8Q5jbSfPzGiOAYDciYuzQu8L0bfPCRJSncarroqmK1R
5HSqSTOqrMs7AwvYEeeY+YctbH6j3HaPRAkAB3KwUUmDld/n45i/Ouxfzvog6aJF
ZA3kPoRSITsx/QRMbPftZN9FwBdmiho8hp/0XWfLsUj4iYRjFSTsRTJVsRwFCEDH
dkQw4X0Gtde6ZZGcG3ukXxjuLcGtfSynjzt1cLIzrx4jqzXV8619oZfcsevPAOSw
jFtaSgOcR3uzAWGHEAQUl1H9ShU2zt43zwiGx6nfFpCCGwglDWUOG5kTuKbGpMJF
frgD7TqcJAHSb21jQcedLs9EyG0lFy/OnD1dIKhL+66POYX4pqMT0bmq5C82XZk2
ggZPy7e6yifX+3fR44x4R8qupY5JXIjxfx6FLPaJ2WWJhwHSG8AOf6P08IcNp1Tf
6FbQXE79AOidOZmAtx3Drv1gABOUXLlk8ASZH83snYkCocOKrLVSnQhjIO0hKLoT
2FG8TQ4tGSaCW4eA3OsU1wcLcfmxJZLi469agTL5kzwZnnlb92XZY0fvZz/HFn4z
Ax6rFApgVz6jpWh8MahLtE3hVH4Tbz/VknxaAGdYNha+zZJfKrg+k2SKCTp7Z2mM
HABmrD0iR3eOXT6kWxRbXun2E+KR8dmyNyGyy62GNZkQ5U8ALrNosySETiFVSVXi
cqZDM4UiVBaByBTBjTMKNyf9I09SLepGiUROHolveJPEzjGmkK9gCv9e0joGHtJw
VVXjEJWJ2CSOqZ5WjAdInEocCuw4AWyTHQs+VuHpIlvlv8MLcTwsZ8lDwg2xxyH9
7sNv6A3JI1imcyA0SWjyxhvuxL2BbbvAnxHyzly8dbqPLZsESoZT5L4bMYubzU2u
1/REPzKZw7/FUKKZZnyUErmBOB1H0WKZsxwi9grmgKtd1XTE0sUx1WlUq2Bwa9St
xMcbyQJ80X9j2T2Cwam3PESMcxQRns1VWvC9R/KzQMRx3CEyDeXzZrEgK/DLfWA5
FErfCm//KtlXmyYuN1gE+Ag+ui8BPzGx/TzW2EQvzlteKy7NmxGe4JEhJjLqbUuT
XEtETTPxyZzOSGv6aMhNBfjGLUB8c0buE63z7KXRWHLw5T0TeWrUm4BkGWNprtbz
wB4aJNYFpZBQEy4EBJcG3pFwHfshAf/UfeQuv2zxFYDLDr9YrqSR0v7g7vqTnAKF
N3ZMmU39Qu7Gw5sOXhA77EX59sS8rsL4pqWpWuUM2VaK9k3GII79Gxxkt7oFhoAP
c25WO5o5+m3dqN6cqG8/FK79HcgGb8OPI/fEHk+w9UM2OTVw1vbZNAn82/+hQ2kV
r10nnlYqI+TyvBqSQqFV32O5SMBgxUTGPxTmckx51QujliY+uPkQbQ7JumOazax8
3WMtUb/9er2nWD/vO/cPyqqnDtIjv5ohwFDRToe5ig/F51J/oPXgrpygXqdVHt5y
TuQntBe43A4smpkxMyoT/fYgyJtgBH8tHZZg3mydofJ6PIAHlvMmhiAs76zpmRkp
fX4MKHt2zYlcQLcryxA+SP/SO51g4pQrzV2Y0KY5nNPS6C+zQHtXGE1oCUJ/CC7J
sVYqovzUd1/4dUzoujVcq1m9CjgdQT2GwuJYqIh/0ZbrsSqokN+y0G58fWsZEXrT
xyF+n6PfAG3aE4m3xWKF0GIBNqC9pg+v7mSdXczUMccraXPZuWP/enYna7ZCBTHL
414ZSIf+k4A722PJWcQY0631ngRs0fQ8XOYvjb6W19JhAbPRU1hDEc6JRipbjZVh
OQqR9/RFDHcxUQGaGpC68SBIbjl0A6Dx+ghuEIhKV9ka7BKeaLfVACD01HuyPhsP
0WdFywcryNIBIAqaoqhYCMiR2KBEqvUpvS2TbXsPXBzsP9EzZtqWhlMgbsefx+dY
NrsKpnh/KlwusIm6grK/LikcGAc7SFJN7JSVmyAFnqQFq06r+a2Tc+L+xMZC1C4y
oZEBQ8oy8pHtJqDDdjlyD2Plr2GpKfrGpTINmDjRqDDgt0+JYAP5ofTrbuyNVDf2
0zsBNH6B+tat5YOQKAEkQ0RwC2U3roA/GCyq44tLm/TYwrtLXlViaITmmrFx51It
AqqyxjJTtCV9m+c77E5nLegpa0vpfMpB3XfXqTTK0w/iv4zW8ac0u74uEqTHcrzp
dszRaQouE4M7EFr5qCi54F/5I8RLIuF8Zs+BctTpU1958heAv3dRPXLm7Ds6t/gr
S/5JWAY98n6q06gt3/SXJnuNG13ntApiXEAYRigupQgLCG1bMOGBgIXxJqMKwMi9
DSc3jU4IYL2Cc+z6KRdTjK+72aCYfrU4f6wztxkidmBGlYfyp86WC2X9KVQUH+FV
vXG0/z3+KuCYsAdSp6tQNZq/N+mHUBXh1ws717IfZ7ZHW2KUFgVQ9EaG8bRNx7XL
+1s7fqLhvME80QStpn4AtIwPcLdXpRtGARHwd6Uo8isY57Bam7ez7STMUZOI4BLi
0c9dZxzbzAFd2lJHmneIO93L7MuOsZZyRBHxOYdRuQBP7uk5ecnYImBFww4T5yn1
+nTJDAHmd3wApczGZJpmpc1y1KKZNf1YWe/8oc7XLu28HKCIQzN1Su6oSKRgQaRW
ygbARVah30g5X60yD1wfHz/TYMGI8VOHahTqe3uRhRNn0v5xFFwfRsTNXBtzwt4j
rlEfpHNB9nCNHdG0l6DbVbdmfXxeqsA195Cyx1lIN95ZiJXZcY//WO+IeNKE/s3T
ze5E7ohOXokB978vcuQ7gmwrXp0RzwmXZcfQmGPySLqkR5kIKEoeiWM6fBskZLs8
/igujjRnWKjx9WAoD+czQJ1W1Iqiha630wimgvVtBmISYErRphUjawQcV5uhXsdD
9I3FUrgTV32voemiMPianNbTap0JNdQRhjKA5uzUJiT+uWJJHEyICF0St6pSbKFV
izX1o7+qL99xCOQAPYyzLC11r6lOrPXwKNUYp/DER/c2SJL1mNWRbECWIGIA9sQs
EbYWbnwtbEbg5B/GOrJJsDatQDbcgsKu4g8c+6tm0jCCzuunmsuw0+ctFYnVAPKQ
iOr4+Q+jZ9OaugHmgPRZXl3RVxoJhKvlJpMMlZHR+x5ECwDisv0cbIHHJFP5QaWz
7GO6ao9gtmIVSNadHaaZAVqXTB9d46oVyt5kU6T/X/FtrGiKhU4QNqRpVTSAXjmd
PfBMvqN19Zfe9dDMWjfFM+ti3FwA6029pqa6CDh6ScR/86AvUixNLDhPNVBMC/gv
kdMidpbr/tOVKt6uclwEG9PQEaZfgUrBax1xEuvNx5/XYb4HyV6v7nIj5Yu+TOXW
Smm7nd5orjQgq58zO3INiJtBpwmzz5YntIhOl7RnDOg77NK7C7eTMtESCxuo3/TG
dTNtkc174mCDJ0tasqsFr8q5VZc8TFlcrgM/oedKuAPBlLaqi0eZ+tO2NyW1fWyh
dPwMAnel3i8PHPYD30vJdQsxCyN4PhU2dmMNv7jjSJ3njEZ6QBaA+h7MXsYVJzsu
ZZ5liZC/LQ7p9T0FJOUlr5Slt3GuNcoKH6Ld+d/TBTz1065yV/kvsFNnezRyySWB
qmO+pkV8KlXavkeo8gKU74xLoSqmUjllKGORHAL7rMX6cjlJFuK/bQ8d7m2JkYok
7AtNeyvbbfwvFCfnDHZ+0oBDJ0yVNgKcLA7Ad1SsMSKgSrDwnNad4o9IY4zBVLV6
b3jQBIwIGKsaQMBMYIS0LiZYVQaTB2QWRZULl5Y7ROf2LD14osMohJkKCuWmcvA0
3ZPUajpZuXPSWyqbEKIkWwerW+FxZspRH9LbXdYuNrh17XBds57g0MUcwlijWtTP
vCRXJJ2OQgCbGckAN3tT/qP8LGkSs6TKTCWlH4m1YzaAwKhXj0nKvcv8R/OEVvh8
5iGdvqHXzXUQuZGHCdWmmrSQGC0m/jGkAS4Kcbe/b26dlYHzMVGiJdw9SiZvF0Hc
TXwvQEdpd/pCrLmHq91rsh71YsxRPj/SRsiYLa49B8bLyc2RtX9413fvD4oFDEx0
BmvA1EVTGP9/pZoix334291o5Ra4ZyyRuZjdfMyX02NQ0vpK83R+b7PCIgYs5GA4
4zT8wboJQcI8mGzZUcotipWYeEM/D1ZzYIFScd1aR82824aLSXr3cHe6RbEsnRO3
UWfB3RIv5UcjCa/I9Ob6AZrJGP4C9XDULlE1PihSRhXAsfy+8gRwUn3Rw0Dr2yms
oqxBqaM8kR2Jvkjp6vATyQ8ALNpWZsN0HzISg2+dIOOYcWezxyAqrMsw9rvWIRhW
/X/fszPAT75yoidxqSzbuQdGspxviRctN3GjKizmtehjBM+j+YhL1rW/34KpINky
l4CNihlzYLXzwXEp8GDp20KFMiECCiAb2tSOAIbJ0uvs5fKY0o2Wy1QneWTPcd4v
hth1Sa4YIzXv0UAZ/oURt0RGWDZX/emnj2viu8s+1gtqvOWewQwJdPV9/LlbqbmL
k+7HrrfPeYHz98ssGHdlXolEeJQLt3MKsfWo+5FbzJ7R3EmcBX4AhZtVo9twrwol
l8fMd4L1AykZpQ3Qz639jGuyzIEbiEb21V5I/Th3Wj8AmhbqUY0Jej0CmCdDdhp6
UKBsS0v8tARYNXtrxst/GFJb71evOyqEEQa7EbmSGrkTeBASUTZ35p1mxRSpO5Qj
sP+q5NBOjEYq1aILHJFV3yDLmlHSzs+o3odjaYknaCCJS1d+le460kfrA2Y7Vzej
38EE/cTqcp9c33XE8z8S1RAdZtqYM+xjoEvrwLmSPzXTVYTvR1H3O9OBU4ZI1D5u
fryjpCDGXo8JZbGmT7Z/CYQPSpSG7JwID9xOfrNi8uFjYIu2io/pezqTtXgKbx72
9uYHavOX+VBohQvMXFuVOJtD2tTJWtpTn+7VLWESEKw685mXkk/CFLvhaGA+cq/Y
z1IU+/Sg4CDJn3grKEvpI+nGk38jMoNT/Iabo0ndTJR9wwpUt0UDIGMtbGa1+OYj
TvS4ofvmx2ORDQX4e+f+ndI4Tk4CvyT2cGUP7y3+ZSoorqCo6wJ2BAlsY/T4mA0A
FmqVHBGpFtsnUHrFEcxldE93mdrn98U+zVd+uJAfrYdXkO/d3CTgFXEO6bzPhnCX
5wlG9Kz+KgCQ5qdy1J4FXmRmonAQD2ixpwRSmm26Y6cc9A92R5BoxCjYppi8GQX0
E1o/uxle9+tUP9tWOb6hna7QSwJitnwNDM58nGg9kvNI6JltnTboNkLj052i2Tfh
EMdtMZEPGY/wysn5QTHQK95Y3NYxWpIBdez//wWZ54M855u0xqmIplukv57AdtN5
fZLpThSin1AvaXbD7XnHvJ1IhHV51AhR7ctUUxwI5jKdzKu5R9dsmMNdOZ1RuM/i
9pnMbwx4Ce7z4HNpLr/5HMfqDUqjWFlFoVGeMJRPojnz945ArxxYEThYNJJVIBFs
nbA/ciZJ7RcKApNlb/i/6FLlL+tcNMsf8dJnCPwhJsMCA9wG6Wfv4TpdoP1bXVCy
AmNFvgQDCDBd6qC7HoLOGUXqj2vTfbjVG0i+iAfrY3JNTxobrsNdQBol4qVltBaS
bVi4PBNsFCzH9E1mFKW3/8kp1eJRtZ8/rZH9Ma3ZLni+nbPwLmUB70R7A6pMcnM1
Aits+FLVQ2lNi9LrVN9xWe6zhQ7ciB4aJYEn0Mzj6P7DJBEqAhNKP6h8Pv5srkbv
afkw+ALfspUGBIpjEswF6sYUFqEmXWLonla7skkHCd75kwqULQ+w+ddacoQSBo2s
FZLdFbLZoSxYs0GjA6f9mi4mdDKTcDi3k2GzNSah+xoqStlEZhqlwiO6bhGflPdJ
Nejf34O/Z8uvcH6X712+jdk03pj+l78BXkfJli7gU+xhrxg7J05iqSNjgKUzaSrJ
trAr2dbjWQ81iQecZpQ3Vdg90sLdeKRlU7l6V+RnvMNtfvLzxJw6sjE3p/pAGtAF
5ksqdZlU73/u2L5w6JaQtLYm+f3yl86yU1euhY6Occox+gEHnuwCq7+ZHW62FCiK
7HEFk2x8LrZuAtzA9OANloqDfpODaMV1ivVPKYofWpkIdz5vrecrqv2falP/uheH
rktO6gpi2Rz7wXJ0w0e3sz/FMOaxR93tuHxOkTJr/PCZF1fUDJ7di2+RB8PTsxF9
bXRqInmtmHEcwt5k1J6ZurDMX6LxdNaT6tKp1VsUlK2fd0stZJY+OxE9jkMEqqYs
KozoXvoR3NpP/hlZHjJpUFvG4KJFszxG4b3ZJqLADT9hB2ducK9N3MeZZWgeVEhO
dWrGJCYWOyNyPIC1dgi3GNIhlJyhLAAlaILI+jI2ELOFeWmrlFJI5PvzUqW8TDgn
GWl3z6zoqP2yGNAagqr6g5G4eOWJ8c206y5BUjhcUZ2WrPQmCRAcssoVfYzhyvs4
s7rgaNTVZZ5d7hJPrJN2i9B8PhU0P3MhE8ONol82kZrdAmZjqSs6Ae+/QIPpzqU1
pOnhB1iaLAlkhm3NzcC+sA5Ns+T2f2bu1PrFLoIyr6f8lrn1VhoTRNMNNTkkY3bF
vWSRJYrZdlCkMt1ytbHHkenbqzLXUAV1/QhMm1P1zdlHcba1aAY5/85S3XxpqM4L
8FJQL7H3x9UDWSvKzROZ0RKija9W6VwnYmJERRppMNZcuPVErGm9krFO4Vo/Ra78
/xbTHM+wCuQPRUzAddJq+5xIAAn+XO5JqEVI0FTVKTwqT7m2S92Pw+b4ni6TGRd5
dyaDbeya5rZtMxt0hGbxVLOUHo2nNLb5yTXHEyQJG9wBJNQAulY8UwruJumFivFD
GnckpPOkkaA+7WK5aEYfJ9kP7A4HNBtkrpTGXTZe0NusUfje23nKMm5riRm+zzUR
Hdc0iFYVCViIXLmtYjSL/btiYz/osG7o6mi76uaC5kWPyOVRNtihV2dfnFjg7/1q
XaIXSES9nyR1eZlbv+LAraJoT97pduM1E+B8r4cYq5iq7Q/SL5879I0uK9vFMZ0P
pCz1jOK2pl8QWduWDTNV6Y/eEpVZyVMlsxud7JRFgqnHJrxEn2HpQtXnK8e52oZV
M2H50h28oSOglqip5t4TJWLXcfrNKYk/fn6/GTdXp6O1Grg1BZrSn3cuPvBS0bMS
s043u7fUXtn9+NTIqh6Yzm4f00FEk/gRYuc2pq3q1MXStOaFMPYcanEQl9WGJnRI
SZXJiLRy1NT7nW9Mou4uo5qu1J+2JqYiZAuU0eHe6EmqpnzBWkonY84BWmP0lEOe
SuBwiOMvHvOtYaudCPQP6X0O9Pp6rgmSqSzatdpOTyJAv/F5e5Ns2FI9pSVESgNy
nOyVjqDcyFBMCovrvcLA86YdAOX0DinIpm42UfL7LgNmCcJaNHGYc1SHC7I7u2Qk
Icn+0ZALLEFfzQQK5gbzfWEJ5UCu29g8PSb8z/8EShSUiwcUxEHVJRYp+Y/emVnx
iPIuXbbYu8YVUYqQ0JcZ62WN0tvEk9AOla6LlVWk86t2qfSTEQjJ47p9eWoq707L
l2XeFQnJ6CVssxOiT20ePgMBQibWPozeLehJpLWH9dxWUSv+K8clbKuq9YZHpeKH
BHnn0PYD7u66iiI26v3BlYUSDoIXtE+skPCmLNWx879u8swpNJvG90k528WoAmDG
HSwtj4AHQMfNKIm5pfWVic4ILIojv7q3xyqmnsWFXvKozcm/Jk9+Xt4H8NrR7GZp
LEy6gMZqYcrZUMCDLV3UzeTgCOMYogkJ/Y2yTt4zSXKvwD/RB6PDc/g9WrxNPgoD
bA0I+TGAQxgMfwSB5MOCEgdmHm1plr8mnX3YtTY0ptSCdxON8WrjtZyozIZ67yz/
e5LV4rufkdrg0GXTwAiwmrZP1qQse8ltpD15CgO+jWBM242GUdeSTpbmuKTm8OnO
7+y5kZgWjwQVAoBgLvGaDaxVI3JXg/unwyRwhVe48qi8+Bn4F7NtK72T4hRkjnoQ
QQy2/9Z2yIDrUDhzIcghFI0ROZ+07MPoDjZhMgyvMRCyxplobhtgYEgCpYxQdrLl
YREiLau7MA28jZSpvZpur9Z/lTFMsUOqQTVufcnuic0aDeC6boEKGZ9oD4Zu4o6d
8hQI/ZB9lEYaJUr4R7aMcyPrFIdEuB3rEB0Jyz+HULEyFolewq7CUhwCJD+Ee1U1
j9Z0MLb5ZwLgo5GX3H7P/atxDZLccJpLoE+XUjLCcMSKyTMt4XizmSGbQTmj0bEZ
CTEylkHCdo2y9aO8o0XZFfhaT/E+qKEssPFDz5v1/35FWUPqtE+F/GhoboCFD8Kg
YL2MEk1iTund6TnK/leaBp5PwM7tCFyuXlZSYXvxboRtKzOBjB3JRyjrPJzoiC8t
BPPVbnjK+zqVqi+ox3DvBiaGRT1JWHE6+pePKeUfIFNY491pEHA7ibSQeDteMU35
bUnmZpg7qK5q48J40cJheh8ZdQKKQ00BVRpmROZlWU75CdQh8hVAa257cSPT1PKy
PJEk2QFyO8PFPMpA8O2NWpmyELuPaVJPJXJXinrJYC702wM7koi4HTETU+FrqgLL
nkR6+z4OwKWzZO0BobbQTewFYmG6Yf9xLf3340n407DrYEcnndBA8q3qy1qceTyJ
8PJ9FKiSxz4s6fRnGs5hH99ewa6GRk0t/V9fiyBGJ4PCCNYzuntcH11yNXQt+9lv
KM8e/mORv4YfJ7+cGCdKeSuKcGpfwDROCnHrmITF3yYCEtSJ6zwpf5V5wGPF5elX
2kB4eywu3ZpJJwj1em+oOvQMU4vZlMVYWO/OmbUx1XEEFGV4VPkkmbCh2B7+mk33
P2o06MmGv8aDJH0y+UwjUY3DmQ3ynhhX3gtLTtiEOM+TnWwOW3o93Puz2IP2E3GN
O08xMUtJiE/JIpyy8u580gralaE0reCLuxcNJfvdA9SkYxosoHpEmS4DU+nthR9i
YOce0abTC6V4E3OF94tAKJW1dRyiU1QGyvOPwE8YK3VjR97MQmbkg8fX7uLw3tsq
UyQLkuIgCLzxqAIdXiLEIgmfbdWKHGAmUC0qOzODOgPux4WA7R8AXLBwRLCln1Xl
MWdi+14OBqA8zM0uUUYvyJL7L4VpuLSawkZE4M/IWqxoCvFf2RV4LMb0qNu3iOEz
+ulZ86x5sKs01m0gaY/qIHIg0IsU/2ZZI5bl1hyOvehWIT9zXPaD7eaQTnHl9+84
Q9qDF5+LQBJsFyn+3u/pMVnJ+7gUe7eaMG6RSQe19gy7bDp7/Z0TYl1opNW1HaAB
FilXpdt0BCY9UAL1d5dMci1aDf35cqY/higTe+xduW+qeUwKMqT2kOsA9fC0zsRv
YHbZUBoLknNyEFBLgjOvXJbwIikx2xDOTjHDgSm2gZo/CV5c5xsHd98mEvVwk1AK
xv9mqkQetpV2jg6glPvB+XpUGz+ogiePPNycZVE+EPWkTKwas8qhZL2EPY9Fpq7p
BV2bNXBoXc2Wy/bO/4ehBsegxZJXb/19kmtAk0aK9H3I4Zar19NbTscitQm71U6+
BpLMDhA/4PdwW5EoRsDDN04Mrhv4jfKSJiniVh5oD68c6bCXb6Z4ENVSALunpJ2N
cD0foq5mNdyfQ+jX1ASP0K7Z/DmsuSAGUV7rqG/5WYN7d307UzBHgCdAo7r/FQuQ
EapJ1e7Snojo+UHRDwigybQrd7MYBU09bEfp0KHfKNqYtnaBlvpXb1muPpYdwcUY
Zr1F1277vaJo13TV8SRY6GL9Wn66aXkVzVH9l02C/wVlNu1pbhT/1nm5qIw6kqdK
HsHI1YTlRsF54rxDJujpaQmjrYdgO1wJNA7/jrbHCO0WYlJN7vSt3ghcJUrO69OR
RxMqV5AtwqD0RlPc5q0qsvZNyRSVs3ORwHJV69Kmhy8AWmsCeNW+JMip+mxT0So8
lHkk8Z5L/a3R0h3duvHz7LwByCaNEb1eN+RLIqc6klo5fddWguvqrJqoKl5cZjD8
5TVhgCRmb4OALNaS7zw+kwpk6YlsGZuNxPp4UL87pOV13m2hSK769OcOHr8w1Y/1
CEb9xWAzH8n6HnkkHGg9D3dXCqiLHaJHe7OexEs96vvu6bgGnQh6OEiiIdP3pcqb
z9/T48SWn2s7V1jpjh3PDUO3G22Gb6QW59aLq3jTWT37d+LtsojxPtdER0t06mbE
fXmW87lq+zEKCVNr7Mn91697ilWZBRR5KW56fV1PsNV8ZP2ToLRpq7tPZyxpR8dK
ESxvf8ZXgSVboLxA3Nocn3c4YZmL6WahTzT4QjoP6vlaH7XgUQr6ehwvPDIw54bB
DyvwGFPyMjYZOqLWKyVw10k2ZkfV5RZFPYi195s/Qi/h3233sIGQUB5uedO2iGGH
b1UXfVNQf2cDW+hKw8hbnubNSATUETo+6bNqFlz8aulH705mxTi8ivF3Vof9gTHZ
utf41cYK3/MbALtztf/xlZhua1YdgdLzR/W3Yxf8j63KaHqqsR+eSN4/Ktsyac1Y
X2BEw2oMkPoFPkWQqMzS4BajW9W3cP/JzM12oz+CcKkOMXjLmrX1RMvtVl97KiCe
ohYMtxFP7Uc3QdRP5hT2xOy+IoMNp6btDGk7m7xvQNMi9e4dt6+HW6ZJgNXTU5D1
CL/Vf0iDN3yAOsts9gWe+zmL0EEVdGAp5F/PItmMZ4f3wB6j4ShRGTlgBBsOU6sy
wwRH/uzpKpjHErm1/8gR/VqQD6qj+MfY8HP37MSVSZjE6vkOokk+YYu3xxQFP+HA
sPsVrqgBI/J0DZQzBoF82mUtQ69fYooNEOoFqxLD66/vVfOQYPQ93SLoMv4fnm6Q
xY4gwEGMRknDDId3XQJDfa3LTcd+zMAgP3uk6VbojrY9ZZCNG0phcfBODqXib993
4ZI2uGmfrcNltMdAkoRAArbK5Mrgh37XMby2LVJruWniiVr3I4GabXN1QFHg1dr3
uZacAnsSiyT5bBt6jz3lAxEls9NKJJsILzXHBb/Xn1eEdBzV1YMhZ93NHbp2wYTx
jHZl8UxXEPjddxSLFHukwtey35xyUdtDKEWybCRF6IE2Z/vxUGLrueseaSvVQ2gZ
7KgY/1qwPv6RsfP/C7vnIbRuENLKwrYSDLu/fRy5sdWortlupCvjakxT7H1g0a4N
tJNEXoOu2E37NLFz41V04+kH0lkn0Aikhkixa0RdNAAyv/9XOW8Fy0yfphg/3iCp
AeC/nwZq50Cn4zs1XthT5g1AhAKb6FG1d4SFv9BdRafe6UeYDTpt416fBEdraPeO
feu9FhyFcK0Y2iuEYBVqiMe5b44oqagpNAHbvOOxcMLuCWh96BjzyWbM4Uldxo7D
GJSdEHeD1B3SWz5/HKNyGEjTklANscMBWPC8DOYb8JLA3abZhv9I3dp7T1JcNclJ
VB8L5UFDBqXHcy53LY3peP3PuluivVX3vHySg+CzMPm5AIOXNDn7Rka5MwpobR0A
jW/zytpzjKshmpgmON4LY1WiPtnr774lVxMKDQSH0EVKg/JDI6o84ovDu1x0nLDj
PWTD+5PcWg+nuN8LKGsRGMz4Q/d9YoVjkmyLBfOaPYO5nMyLDAVyMRe4u1axYllh
YhrQcxdS+d52NZhAO8TYv5axPB4kt0cZzlqs/6f33z7BtTvijvTriBQ5OIf39N3T
9badVoHSPMgHvvsAdVYYqu9Joop2zA/35hchOQjYURYFxiOVGe0mlu03ADW8eite
XpVYyi8Nt/AJnpvKQPs7dJUM6ftzz9GKASoZUd9riU/WRpb16cTQwIIP/RYNfvap
BhYKU+GyG7+Gs72B0L2Waz6K80xYs4Da4VuahRiptUsEEcE/FHvJyn/RQU5OC7jF
bJEXOiv9RvWGq6e2ZxMqKC9uHj/TCpXsC/SkSxp23UsTXWoM4HdsBaGL3kS1a6NP
nAu2DEyQR7LvlDro5efBrMobP1cb3J5gA80/W4TFfPYR8omsWmdDWVv/ZvmtAjA/
0l6OA2LNoaCeO83u5eWRe5gaPxiYKp0yVQVF2cQRNYYAc8OAfI3XSaeLqAtk95DS
5foDo2RqBXATIr8q7CV3yG7SbAf516H1mZb5o+eE+VpeD/tKZFyI/0eeMeO2QSWW
7oTQW0QQDhX1XISCtpfr5lNyhS2ecWUVFkeDQehS0x6G3hfy8BhIjggLxMeMFq5D
seUzUiWLqih23mirgt2Obit/tIViPHwjkwkZyR2JW8qsdxCrbeSqSuLj5E2alHQ/
W2NB0R+XLUZTcGRlJNrKdeJgSfLyJ7R0x2nfODDFRA0xRaE3IO4khE37GFxzHHb9
7Lm8scO1aAJWvdBJtl19bKtBEQJRskH6945KdSxhYk8W7OpwJoO/TBHKIw7IVIW3
oGK+5Yh4ySmaCWOfKPxnxcNniObU0dXmVyturqerjlsrMb1R8Befh8OkoWJrMDPu
8v3xU3lMiW8pNwhMvhG6Fa91aGl4PBpuim6QihtRewW8OF2MmvveNKS29tacrbVL
au7aquay8/tQSDr3qrzvHpPKzO4WhyS0MIStNXTbbtaAvJWtPOS2dJydIIB26aOH
C1HKt/buprts/T0GZWzNID6Hnzf99CxpZ6pUFCeguw+9aRhOOwjU73UIg0oPC6kX
gAtTgdMyxiVzRCuTzcFP3A89gMHz4oz+Us7zEVWT0o5Hx8b9V+wKNWnM6Ow+Rkly
k5JLiJ0ljp4mGn9GC1OP8WWhxACvJhGgL//vSVhxJmLXYHh9udc3Nudry8nuI8Zx
LcIV5ufDh7UCxwm8UMrs/cjDsHeKrtm2ae/c161xlbLJ1Kc90mowGYrq3dL9SOPA
XbqCOv2+J0C/Va3EW2EgMzh0zKoA3bLUyv9BHMLtZ8KNzpljiDfvDw9D8IHUvxOB
4VzGDD/yuSguTsCZOUKhd3/IdSLx54iMlXbu/ABg/Dy97iHOExqOsLOy/OIpAOJA
8b7v+APicCoLSgicNP6kk4/gt/uPyEeQ8oKnglvC1EMEmux8u+BV4Alh8YgJIZCk
MInVe5spJixSpDW8/tNUNDnaP2bFwZxYXq4S4xaPj86jcygX63SlgDzMYRRKhFCM
4i+4AI3farn7BKY1gWFYRy48+1cl/7VNkjaKBOBF1hGBLZkYuuHGuAkah60ppY2n
cavnHigeFJYJocHlatKEW88qiz82QnTFttUkmixEefEbJyi4W+Qqc806Vs4ypR4Z
+HzDCV3WoiaPDnNrgDrhO3CQQtAzbbK64OZt9nnL9VHrg1C+sEwzF3bEbetxmf+l
9kGTCejUPBmPNbk5KDPJJF6tQa5O5skxDp1cHoQySlBqKc+uTIJmpILGOdqPCBPF
YXkUf22oxezkZG3g0hPVi+sN0X/AnfHQ08cIlLwLGR27s8Iofy5LKDx7FGIl8Flg
H4o3FuwpPw3Q0SIxXLe3t3gGz+Rfmrz/k4o56X76ri857oq1XYW1fk/hODrbHbJC
41gt0RpasqFmyhus64T33B4KA1kZ54JFuMZIlCL0TOJEvQVagOGMzYHrH59s+Zp0
PWVmjrnngUecdtB3NInbiwP05+t3rDGhmiIZVc/2mvUJqK/o01Q5i9ffqGNvb9Mt
YgjcExlHoktvD0isnCpDCUdAgWMPjQ/tiT1v+Mw+N1MaGR5qyaV6K/dYxlmq1pkx
iC3IYuXv9niMzbhac2Iv+Nz3CMWk/ZjmjIZ4jGJAtO24vtboSv9FlsObCt4FCKMk
M43VTHku71JIv2ZpMiWLCKZq5RTm5aZ5U/kk/bk+vSur8G9NYg5nwZVlAOPN/oNY
TMGWI03WjeWraJ62H1JzL+9sUKfSlFGSTwt6SDcDbQDya3U5OlVdCJ01A8AlrQqA
J1FDKd7tLUTRc3gZRxFwtieH4rIOPBYH06sJXZe08bpBPvonlDK/N7hDWSKAFS7c
wC/zH6RYfcs41ChCpCyghKSJNpv4QkA6euwOJEw9nLG99MyaA210jicGStlie6Zz
keUA0gjLPZnUDmWzEQB4Oiolr2evnYj4kHwKPa/e8M9vjAaYOTlVvssEaLNlPTAY
lpTJ8e25zmf590I16PYYolgxqIAZmm39imcTo0ckRea+HWBicWT/MP9VRZ5wWbyo
Dw/O3raLMpw6G2fKd9CPQ0pdP/8tGHVDjwDf/nwIRwZJVOywBa/6kfZWPixs65eS
3nfFeEPnclRbIkTDbTjuMJEE4jO+HPDtp3MtCKbelUooZxrTU7Kfou8cjgb0wYWn
PW7BcORFTXzeB8QgbN7v+9y7ANBssn1nP+A46mQvM2g4vV31J/dkCmTkFr4uIwa8
dqFtCFmeP5K7PBGbrsDiyoilsvsJdLVMv635AxGKqG5cQoyMvDSnpxKACbKyIATM
AKHpD7KrSbzWfbAgQsYlzj+GH//YPiLMGRqjuc8G3NyP99lK7wK4110Ga6y/rdgD
PmznuPohsOH/gWhuzGJVgSQSrDXm6LM/eQvATJIUkZSC4CefyXxotUlC1iBxrob0
1EXrOKFPcKW33ciZRCNbyWoSOT6BeDX6IBZAixa38BCCcmADzCz++FmoKjJBgNn7
3+xaLOOsDH8oW4UIXYXNxx5XYGS29RMUdh4qipK4hZKPnBbVSFLqWtCWCrsAa+Ik
AQmkZDQMOeW9sDXZJBJRqQQcdUYDGpmlDKi6KlJBgFpXek5JVQ5NFj9dhNRCFIh+
+kfsdhFOqqfAkvdbW4Yuzh+IHxlma1D/yRZIAExVtu+1KtwzXQyba/97Ms82MjCz
Psw7SIqHaCPaCyZ2JzVLM1LMJbnr3B8C5EUSCiAc3C33yUTgNJA/XhoonH6VIZUz
XbQkVoESKAgkSdrnNpvbIYn3nVQt+exkuXFC5TFlWMvn5miLD1EURs+mPnKRBGxq
DOOiOXYgg2QnNQu/7mN3bNChZ7GU7csty75xBA/U1WEeblQUoMwqarPkPBr2LHYX
tSM0Jkx0n0p3k7swQpxK+gGJ3rzp4+DbPkmmfC6e2+ZIbANMBqObnpwd+4zz6bHj
p1hYfjobWcPbJPAAZHKUtQxfH+OQcFsZXPVoTlSnxeofr4tED+bGT70s4ohegNeK
BwZvkoHDCrLX0TFp28GodF1gmY29PBevp4Yi3+7RBOHVVDikuCdbZN1OGZCiQNGj
TdMV4OaHNE8gDSgrVhR0+qGUF/F4XrwVlshcsrFxykSiKOJqXW2LOgViQ4bZdPQY
XRrJuroQZPnPlo7/KoPdLxlQZYxGtcAOqBjDnwOBHuDvsgweYpmCRDJLj7G1WFOw
yfWMgUdCu0cyRKGsQc5bbpkhryDovCmGvcbJGvJLELEPG0QMU2M0V4KculIeU58Y
fKaxcRoj4Cbcz1hkvNPZj8+yJfocJVrSY1IceE69LXVGg7xFKWWsAFl4pnORQxLM
iOagsdZRhEEyjGj1G6A18cVBe4MFEYzp8uwgrQPFCl251Cr72JEQ1gpLYr10mg3C
imFJOuA2JFzKfNlNEmGOdhWwfxGJyJq/fscPVLjt/Y8UxRjcS5UqBZZzYTTmdlC0
6fgwJYtwG+Gx4T/egj1NAXMysw8hQuRfYekd/IIWMd58y0CtJq0wSctCIr/ARWCB
e5H3dvq9hWriCLF3TXJXQ3FFKvkDvVAy69LFRypDCEDV3eiblt/eEJ8p6XEtZGj2
fCTbgWlsT/vadqvSDqagqmDBMLpyVjhechGAsihIT4M/wBAXLwNT9LuTdnMkpw4I
+vBa6MQlLRkOyre+c4vUu+IpOfJajUdJPeHiuDhZ9ESsfGLT8UOJqh/quHiT6xCI
P+dUsOVNAK27B4FHf3YVgewt46mVUNNZAxjhvV8A4yZjC7sHRWnN3QvMpw7Ia2J7
8aSmnSoinckk5CAIR2DWHw9AcaBbGxby2gjM5SHsSq90XjQvFfAzrphu1jTwPKro
pcp6ru63+4Vt1u438Igql5//vPm7kxvxxSo2rE2QIH42jVfJPsRayMI4KqY76Bj5
ZSTNQkxIThUOc6HRwYV5H9t7F3pqbcZ235jqNbGO1wOsAyCzbDWNgfQTNKFPdSt+
P+s1gmg4BGDQpaHfYmzeTapZTBM9edZe3CAYDx7YJI2mev4vgmKiHGuEMs3Zm9wt
UrGK44Mw1FGyabwV760wyHKsaUvD3FNoMvupkELfPQ8/hfEVwQuH1Z+NQRvpQgQX
8rpWgIeOch0c0z79I2uxhN+0WoLZBcPHTue/XX2GydWUs/UZ7YMZrwqQMRVItM8X
vcllQHQoTIoNwC7QcvfklPSgg/qg8iGDgsRVBQ55VR338vu0wYqj+W3Qko8vz57X
fxMq/DX/uXrCLLQ3XPd/w43vFchqAAvqOikQtPan8+Ji3yEpT1BjDD0xw+j3aGyc
/H7nbkBiMzPFL1RoAd/ln9gFfT/gpz8YqMIdQBmVcDT5yYGgHgBdayK/8KfIGFUe
PuiaeSrtMeO8wbJreF+vvoLi38Zw8BXSelldLiaWJQlZpAaB5Jw4Ead1wjW/B31k
8tNNEOxtkbzutNvLz5t9iJK6XwxQgwfkQAwse01pKH0WLg+1zCLp/8ifqtl6uQdr
/nU1YnCZxLOymcffLBG2l5/3qnYlKzwv2E0ksDcO74G9iDAakXcfr4Buf1nY6CQy
wZ2xxv1ibIw+JOdxxW1h+bzI0ZMKXP5oyBgu/dbQOxiHuujFizxkiwjgHVqOol9B
6RYBCKTcxNNvM0YNVcEBbYEwCeI9Yq3Z3C2NDSSFgS9t/xdOS5hXzVdx6wvWzHZ9
eyd8FwG/dv5fX/6h6dTglNR64QAgWTk2Mid5I5U/kCCQ9mpFhhrJ6HabOxUNpVmP
HaG2fBm5gVJpBnU+zrvY91G4Hla9GF9CJH2ggvBMd9o7R41iT6oemlVYQcB5SjmK
bhec5unrkMsM/8RDPD4JJT4YB7XQ+jT7LJ/U2gt10EurxfCBmXVRPUcfNv3XiDhD
oWDS9aaHbuDoSK1yJPJii2coIOE+iK157d4221MvQkBvd9nkmdvFzksX9CoUzgNe
g3a0i8A6RafEuTB4G0esv19l3QhMEMAmuYxsi0ugJ8UBdHLoHq1479OCjib/PGl2
bQTN/dQzddU1LKOP0IOlabIbAwiSYrS0Ee7Ug8u0mv+oSNdIpNsH1G9qw7zdlj14
Y6TCKaSaGRaTMyHv58NlPEgc1aArR4CzgXxOxGZy5A41g3CjVNWqR9l8UaGFtjLq
n66AkNcMCO0E8mtb/RWD156qYJVi+LGLq1GvVIdUnOjGpqFENaRpHfgYOT1A2evD
OdBxSkQ423En+uAg1B8YQ+3z0pIaGkJT8roIlt/d7KSemGheAhql2I/UOfQwJ9FH
DpHobhrYQKBdDWetzR9xvfHQ0Flf6mOWpX38zUZ4Avxl4emT4FQsrAx0+GUfx8Zc
lK8AfQgOezdRbjdw1e5a9aG1dzOK81XzBjKO2n6ivw6EpK3dIaOuxGDnn9JGZ0R6
/xiDOOK9+QDsu1vi2s/Nu1NAganKimFD+AfsxoS3DXzotvAuTdqQPZiXg7QT6lX+
HE1D/n9d5fRqLTr+XGkI8uI0A+J5WGdwWRRELt/XlZwANecupDv8CS7eRdifSN4/
LsuCFEh+Le87TuRIGZMjH31lOZJMrBZFCyqIKZ2Z40FMsmSVjHWcCP91/0hEtIOk
NjnTYryr47Qg+Cog9SlHatl2Pf2I/BzSs+Q8Lg18+tPaPfa+9SwjSWK3BOjvb+BS
2lLCyHZqLjKyF8QOZct6OPx63+94J6ANNki30lXbkDprcQuKpnq5vaPM11UQzJnA
pix+15xT/ZOlysBsolE8wm2poztCLtTdM3fXw9pCqBkJHYtkcXrf+d2+0QoX+aq7
XaXV5h9Fi6RZNIz3BjmAd8QyDWAv46jMHZ2iCn86QWhFSLeGg9c3hLE1JgZavBh7
CgCXh0IEx/VeWApc12ucHahhOJQbX2ldLXI5/rGfTnPvaNlZzG7w4OuYmZmJVsXR
fSLjjwLPDhUuQY+jVI0ihMZxDICbRiWxQTHMyxwXwk8n78pdC0s3SklOpTzA+Uux
+0o67zX/FcVykn/ea9XtWV1MiNEp7OAYwBaExyQTsL/byb8owZcrntcGfB4d7wc6
mtMZFVaKm8dHFmRo3PmYSxYFvFb0fAECwVdrfhr96ZH6PieD9lji308rNk8dz7M+
ydOhoJcEOjFh0UdIG0X2oitc/VRY1OxHwG7leKdxtciy8cvsQoRW3D0csuaTPTpy
eRcUz+p/5fA6ISEdhYfDWKI9jnnY7xu2D3x3UFY0Z8g2T87quB2tIidIS4WxbBAT
ynSqXb7gtG+X6GvtJXrQM5gseoG6ls3M/GzcE3Nvn4ERGiFtHvgyt46GFBxRP1d/
wamGqGO7XucMMoMX4hBaUOgLQN/v56XrojMD3xEpM7oGGt6qH+UYp9I3waZjNokX
fC50WEaRkz5HyJrTqO7pyYkUUdEKVyCnYK+79cAgEXbukGAnD6e1cQOtVC5saTQR
96lyuRAQa4ttU43eP6p72XIstAiJUsV8BJ5FJ0rPDJafUTctbpG+6pQhlU95iEqH
qTp1mg4sLo5Ub9JAaNoGLeEqwYM6AScMg0VCd7B8Pov3LFBktnEvoettoADFM5Q7
pbziW6gJ1JuLeetBC8UJ259UCpFd+DU/dpCSx+X0tphVnK4p+8V0D5DTpFtvYG5/
hxFIDfNhaQkpeaq0ZFEVDNV7oDbmpqgSDb5dUtgFWAuGT/BsrE1/sqDaALj6QpZh
uBYe3APDkmAdFs4M/6S/rDch5quUxcPtZGTBAvK8gklWIYZrqqKP5OH1r6t3yTFg
XV9IjK8QqkR+ebl/43SuCGiIPFPQ49psnw+J5t5oVHEMxI26J7usr5I1s+mdPS7o
26ipNzMbyNJJ9OWiwLpmWa4jVrUVxtSObGQ7lCdLA82Ygw8BdWpeRdqJwg+vuawy
guTdXFHT+mJv/HEUZbonldYGn+uWcTUl9A3xQSp/bkru+8EdOwvYaHON0eH7cgs2
hyki4asR4yECXD329lOfSBaB2cMNsFuePAGufpS9Ss+KueuPh9FJCNdrDZznXfiV
PnlO3T8MGAwPdLp2sPDBxQrva94AkVPUNDAkXlbLnoR1lvxp62fxsMgu2xoPJWwM
ebB8mUo37yhoBlQK8vgk+/IQhfgRU9/azuskxVoHlm1U8orNpn6etM+wn6jpyBrY
E9nCuvuoZm5wNxJDkhmZEyfiHri+HGQWnpeBxgH1/ibWvmT5e8nxxod5l78exdXy
MuxgPBmt5epOc+zjCxLDQ3ELoPftlbV8ZfeNC0sEvuspQ74lm0+X5YKtHpGozznE
G1CewQfRY1Ln5ferSTjtThOWfX0lZPQI+iLjt+fCmH1ihaDjvLymn+t1M4lZL2vN
rZ71T+72fgiLWXMNzeO5Wsa6NUK4FXO/eLPrGZWS5ruN7RB51Y244al4+LYXlWIw
Ekeh76GiJvNZ4df4kWK/nmB2TUTr10KQx1P/aZP8QMJHzUlyAfX5l9zGp/OcLoGZ
UyJX7oVFyihMvmxEiCKPGpA2rBIaP1EsyBKn/mBVcayJtWzJF+DTwKCl9hN3Lcmm
Zuj091F0xIRcezJMTBQf+nFHiPXfeDA6E81Ya6IAlvTDhV21DZROdB2X8mZ+Gzs3
fnuDrZpxkjzCh8zyny/VTSmYxOIZzg5T4q3MNm5eQKpjvBUTGJPIGW6jFuIZZGXv
eVJ8hfoT7rrtYetBfCa/8X/Iqxpd4/sN8QEEYdcaYQMWRggWSDkVlaqVcyVuay7H
nkIr1r/pOsCfiRZbdBTFMpjhUEmQ/yu8SGG8UQk+M+1vGwYR6EJzCHMeNNd1AjPK
634eZz4dSKs42+0XE3ShpLpc6AmuO5H58nss2Sf+uFVFz+5jYy/hU0LNUvnoDBOo
cMJkZgIxgkP6f+oEnIau+kK1AO8+0xj3y8uvPETLtQGZYJJ1VYGu7298n+S15GG6
U0ZuylZNsIuZBJRQctEeq5a6wEkIWq5YvxJymbbos5Xvt0dTYjCOSk5xzHAqzatO
tWs9QQz5RBWdhwBZa7YQ4OM2TMidn6QwvNGKgW3TqYU9TOFQfQBJFjjzcylCQNM5
ybDtE4BYS67/jLnTG6Liy86g4Sw6UbQfQfYhYYoOwvU85alJtXmkigU4SNZNjijY
iuO3LsfPQUjtG4W35e8vnSdYKpECb/YL+NBdmMNOgmoPGldxSlyTm8vLKyMKLf+R
faqtCZWk27d+av9OtqGec4V2/QHP8Ajvxl1Fz+dQO0BvdBieDf0N+4hmipOpcraw
dwJVY7aHJ6eyxwFdANPmsraaKtf0RNQ0wvVhOeONw89vYW0vZT1Qxvx1JlkmKVEP
PsGsn/slz32TitkdooDgh+G05gVYzxV/UzyEz6tGQvWP3ST3a5GDoRPvkZVt0WR3
cgC6iRhHRi/hOyPZDMTRVHn3OjSLx+1CxnLWcElHC3W6OaTABlvuAHdJZrky7Yy5
sQKUNEItWK1dvkxFzZ0LLV57NSSuGGUTEUgXh3vL5edsJxCwp9yXl1/qsAcFqfDq
4j1Oo6BmoUEHSj/k8yf30tZl2PuzoUI+vXMRwu4ABMfsopHLhOyEEyhIC2RFvHD7
aykl6oiUUxE0VbgwY7zv9E4+npgg9VF/Qi7uRN/DcNYwdH80N0dlAQmA63S/l1rc
D3hL6IenBHtlPc2FLSwMch5+78n5oIhHGlp7pv4TyRxv1wHaipuPbvOTRX1MF3lR
Nb4YIDJhTztXB82hH5fACoYHmKNn5gcoUKdj0nzs8Uj7vVujXD3WoaMUZT/0hx3j
F/fDu5jGWW+ckfDX0S15p8ucZ1eOT+JE//UBWbq66486XGjlHlmJC2FeqODKNs5w
dWSHZONzYZa2laRLSWGLUQh9q/SnVhlvs5yHhmT86jAYMW0kmjDsQ8+aZMLeyR/Q
dbZdW37e+SER67zx46uTdkaletMkhsZmwew02PxYqltVLln0aWwNs3s4h1e0Jp1o
m3LdW7h1b0vjDzp4/LDGyTBpA4EcPhnEvpu0iovkfjhhZcq4kUEhAS/RVsKBWl3E
cF61kpaNZLcG67V/fUP/kYpp54rm3bKVsbck9cIB2gqOcOZLfX4h4QeDjUlCxMaE
z3t/zw9nGX4JkKMEJvqWLZriY81Yj6BW7HQmuESv+7lcBdWbZF9eZm8JItAxJTpa
+S+i9WOn8CMPU2VLjAnHY+YNEwcXvCN/Z0p2E+T6kbT8G8vDqHUvGQ7Rj/QArMe2
WAsXFzZZjIeOJV9xiAqa0NpUEnbEffopArH/WskZg+Gzx+v7ywS8tDq3RDLc2jlu
qFk3yTy2g0IhGnQwWqZ7vAFlCznnl/Uayze3z/f97FBdDHsgjVXbsFLueY/lt5tC
8FdlI/OHYz6m/FgAg5ywm98gz8yauEr7jWLg5b5XTjanZPuRB9qgdgdxoHLM4bX1
fVaFG7kibgYEZAfP0rd/EFVUsxaaIcQB9gLnK1Z3M43m3PCCPF/Lz7oVftEnvdLn
34gK9GJmz5w6GN5dA0QWwD5DdgIDrlZ4FmsjlhvK+MVsJrLyDvu8AhGVxjt9cZrK
P28AZ78zJhbu57EMDrx5zJvI7U/XPfphbSjCZDiUbso5lo7OFCZGpwyG3r/Bib1u
l9E7TVsez+8OF7i4feSLSuAbaDjVXcdb3ikS7k02Fpcw2T4eLrlg2aTy7clFojqc
mDUfKDHf6ZnC2M9rO5gkpDXOYa4Mmbj34YI3fbjYIDHMk64elCryMXthnTCAxS9e
q1nQJ+romEmFKl6qvWBWwYxDyXd9myRKU+BnWO+ez4q0T/y2RZ2Ol+UcGN+M9T3y
0mPjFF4CxwBefIh4x/0wlVv3ZMD/s/7Y50KmXQFiKpyFZuoXBeX1p/GF2YZymjxi
1Y1LtpznI4JeWgJKlfAYa3j8gwdekcRaDNaZgdjrEMBYdcTQ0Z5jnyQZx1u4wrW1
ZNa+miqzgRmjS3f5KZyCVe2R+Vk4oEd9vlo3eWcMG+F3kZk3VBiILZQ6rw4UD7Su
iVlEEDK1VD3C6Ni8dYR2EY2kSr0OzgPtpWFSKUFci2wGXjEqguOHERTUHGbx1jur
inXNTvw4yQAd1mDrPSbxfRfatA9WWU1hArcDRvTxBLJ6Lp4htLvAvZAxVFgUNYyw
CtBDFGgqwQ7HTgR0NhaSEgnGpeArGMQ7lob6ng4jeCCoHG1PprTKADdUYDIMTqn4
JZciUwJZ7uKfbT376XzIbkCzqi/rbJpkKJmOXwJm8UTotWd4ns/aL4PKQrgqjCZn
sES0+eoYG/6CGSveU/uab7O6VlHLs9eB+CmAMqLLpSd+oaQGByvlhLKbfl3Fw6Vf
/1ZbkJVLZnc8YHz7gmvHoU0WmUQwleDd4brRBc9dofPfZ63xIXBUUGjuspbv7NA+
5vY9y8xhb3exR70h450ROhuePSSZTeVttm3z/jfv/3HgudFMeWqquHsI3McxNE+/
Bmp2uiUxtitjusaXsFONfWvlTIHSp2fEqZuwdYiYaKAecbW19WoLB5m2hpIDjIBS
1rjx6kaBMwmlOxKjOOdMkWRuagYM7izN0v2VNMvzMP7qzwGoqKQHdXoep3gq5hWj
S1zZjhGMtCLGOWsuONJDvSiSMuz7TygWsSzrjULB/ndvuRFA7ZMaHrLKLu2b9PZ4
ahB5fiXF2vnYbpYF7ZOcStGVcvF1gXZNaFMGJ8IRKFLeNt3W8FNJCtn7/ghZKelv
sUSAT7KbvFqLMdIu4XXSRW/fVsnUGCDr1UOYbnoEfJGu7hwsbhyewa9bOmjJLUxR
kJyTJNGiMuc9PY7FCatWMTMbLxOSIXhBkqlIgeqf82YIr8UAJRfuY3ssR2ownFpa
L5G+J5Bw4Vfrgs4QbXtfh9cRUGA4klRStxwKH2jX0hFvOcZnd+9BGW8RH49mwOob
nBalrLUpzbSSb6Oi3voEulkK+6Aw+RmIHv6AFrgR7IKX7f/sGaOP8/hfBkNytCji
4GdBWJuajF4CsCXATBa7yoF3+o8x2CfAwe5/jdEZ32b1bbsEd1Z+WZzgsf1536e0
35HB1m7wj7EJjj0WIip5Og/SX4O1EW31CS9FvjaozmixiyYMY/xhPoGsJvpKLNtb
PIly+UObobQDNdFL2eQfVd5cjdt3C+OovlfsYsD966327tif+2rxmyeM8bvpVqrt
ad8NDyeL38a+agokWOpC+zoJZFF7iaLX9qNOv2g5YxwYQXv1guPuuxZ7Z2OvSfrE
99HN6usDtId8Lz8qocU3c9m6YyCnI4z2t+1e5ucHCrI3K5FeHgRE7ZKzeeeTFKvv
x3HRiQFeUVjKzucnywcMj59xIHSeJt2bGdENFn+maJHda101zLg6NJcZkFrxuR/P
a0q8d4DzFgkWEco+YcCRFHJab8AvK55nxLXBhMz5HHPKpEj6zCtmUg2N6ojWay9R
Nk72KQQsycfKK5eH4zLdhZPBoX3FjCV5AmbYdJXCrO3f49gotAe/3aDrVGpUBMdg
VAYxjqAb8j1hWWmPhtp0DAcKA+5u17yo0lrRLzLy80TEtoA6te3UqDE/pqkgB+DU
EKma36b8AYBro1I9QhEOALfYtkd4J3/vtuwGJZYJdqxwd7mO+UMj11rZ4r+mmX2X
ceKBrs/rgnuNrKEkMliIDRe1K0BtbI4FJfHB3F7pPSQwHUiOnKJvFZpenBC1FZs0
+Tq74vbKOZ1ev8t3GtlKoUtFFPNdTEtpXFkcDb1AaGJs0SWZtFSgCDU9AB5zlVzU
PEewHEa+kNJV9gFCT47NjlEIeWKZVVgA4JcMz1wAqKViZjvYVaj12BpPZXK4FUmC
KWrMr7c35E0NVB03F8n/b1ChOXEVfWpn/DKbG2+T4iEqPL/JRszGcvpBnJMl9zuW
ES9q3U3REG624P8IGD8kzBRXrycpvd9VI625OUsKu+Yq12LDPBJwo1mCnIP+6PJ3
8mq03Z3f2m0H7U6Pt8+T28NS9VzECArlGQgeglWHntc85tiXV34kC0X5L0GTDuop
DakwxFurx1N6xzurq80lZWaU4AkWuJFwnjnUSDI7nn4cdncn+ZgInXigWsjeFknY
6iyxvgVxOOo+7mk4a2067onW1xFdY/Sb5Dz+0Fw/8GdpSjULuV8eocv57c9XuiRT
Jn1e/lBu7UONCCjmoXqyOBSRUsxE6sv6ptJrIH9YcxqlO+0caqPkqjlR176IT0Ly
G+JUhkkQ39HMMwybhjpiV9X1xeNwEpUCFaN+nm9voBhe3+iWR2jaNHimKQoye7ZD
eufq5MWST+c2gXmh36T87WmlesJSZA520j3OSzaKf4+q5ZWBzQh88pJhC1JTQr+T
/h8UTOFZ3zQgookTV3m9NyiAaqRaxrv3q2vpyhXzEVH37aqhmtFBuQBHLFckvShs
nHLUCAm30YJW+sihTyAwyjYynD3gpkt4Zz5RqXWOmY6F+2T4zcEFk7+Gxv/c15qg
NtVU3loOOuG3pdNDZdQCnn7NoYS7v+kgfh1Gts40YG9R1LFxlccBxFfeLx5TFO/0
+xO7E0s3UcdBoS1O7D1zolDFhg/qVRKJir4Sb9hPJfFSrSefHr5BkJoVZUrQNNSX
ilEiizVnXF4OgL8lkWcA9hWbNLEXIsL1Czc+1aqH/QtBSSQ0NxneCQI6WD94oKHd
0fc/4CtBJJnmnvI/XYbvgCfAKTCgMBihJtvBlfz9c2K8QktvSOrBnyXhU6Lf3LYZ
4h6idJLSSLvnpzOUa6VzcK9HkVHfx48lQtufWBmzvxzugE+w9SRN1dIJjDY7Jgf7
F3xDUJDqOq2+EWQslqz5eldtgr0JZmAfhR0lbbwysxKl6vF8QPR1RtaazpFP6K/u
VqQkIQfwklRdohx2q1TmQaGoEC9BZJNqjF2UjMpkk4CnEfuc+AUw+u3fR28QNPMG
+FIZL+DBXzd0YBsKgNlHDDr7cVnHVHKNpn7EDsooyKClshZGNBp06OI7NLYB5ntM
jaPpTUrRII5zAcoNLZUxUk9kwh/lPwPDYu2gPv8AdN6oaNMhCfyYS0idCYNQhNsm
QFsQkznrkosCugfGoiojTaw89Gct+U7kcIa6lDOWBg4iJ3f6FGukCcbyNEVGox+L
WyQuNk+17zruBUd6nBihr2vwXcSH2CaRvRE5c25b+Lj95LD01LuYv+FR26bPIENg
YT8IM7561GPpPdvHkXFvi7FTtAahY5JhX6mIiCF70h6MkNfdw3Ey3IBMg4bODppe
RTISlHGWQIZLNNMoHwSDK5yRQlLA/IxHS5559limSdK/lZ4ukYMRKA4cZN5ZXpAD
tnN9eCbd8/kQl7lbOz1RYaZ0/2yCp7aIHEtk/QMlEUix560I5BgCCQ6uJ5sWROcU
PRo1RpTmQQqJfP75jcDMDUfqFRoaXU/VAn76A35zaNSrym7j3WmhDe4IaTSKUuFT
ENI3he8qqR6n47dS2Dvc3g2GhBQLM5sVMzynHRirP0Pmrtm7Cmjw8h3ZkC7mdMSV
4LMuotJga8A5bTeCEQ8+x10nqq2uVNkd4yQ0SXnXCmBqt3aU2rqY4N8TaZ8PkgVO
0l606Vfd/qaNBqL4asQIh+2j9iR/7FISxIuAUqDfxQzFSH66OIDukuZ/15urEV+Z
xrKciFRdlI6GfunuxuE2evL1L3IqL/xr30mFDEB0On9MawT3W5rSZivJ7v/eWnBj
LywFq1AB5NkIlPNsM7R4c3Ej8y7e8+01UibhNnnDuPyF9E3iXnsljmPcw+USXj8/
/MvKIpP0uFkywymdu5nzpC8cdMdhkLjYPOFQlD0FYsjmhk5umXSu9QbHfD/yRD3v
xV/tJI8KRsg6R73eJzlVuONkwPSqCR8mQedjl8rAv65CvvhINpB7ruXcMS0hZMCe
VAnn4xDuTXSWK74xkUdE0dSRXo/BDxtu33+v+ciN7bRfVyK8IJMsd1JNsSoKoGyx
x/V+/kc2TI5na8ujA4meg92D6QW0MXjA0KYP9MjnJlgv2DrgJ5x9D+b++7MDPtHz
qH7pMSrX1y8f/7gtRR+5sGCA9zQGVFncOI0VgkswzxIZkvmLubc7194Fwfg57stJ
YK2XhhV93KwS4T2fz8u1FzzRrcKCmSCKm7RnU2CLa7vx3t8zYYX3kDUx9BskeFNL
L8Sb0zCcpUXRo1vVqLR0AKJk6l8u6q9/XLxHenyjBAWMZ+gDwiCCURlpJOkgwmzZ
+z8/jMFjQevcZnMBw/ckCW7A37/CaNLrax8SRz8Um2PuqylCDkZycPfBXsO7AYWA
XCgO0Vi1DjjnDfio6jnQDaq+7C6LcJm3tfEZcP/ZMqOGtAy6/k5rxiSGavRnFjYy
JdnESr9Onwx8sAzSeHv14nB2gqKre/Wr+KpRmt5oNNFD4J8Y9ocuWotzWEoSj+78
csgsZFLYjAhHIi/6C6ukHLr9E0MEfltFNzo6Ul/BVlfSVd+fP4cbfn0+sFGAjSlZ
uVxmYxnWCLlxTa1X2/Ov4gYDy//sMGaFuZ1EeAkGYeXuY0BlwRC+4DgnZr9yjpVn
iy98ZG1J1dY6hislwfcGIwXWrpHdd5O/5eVbLkedsVTMJuTeiU/H3sFGnOrl7rUa
ObTwgq4DrC49WbQ6zqBSegw9NLoBhk5hREIzXPVuf6nmU/M6uHC9pnNQGDIEk6X2
zCCc6IwJuLgGmbf2unO6fdvn3uCByp8BihEpkApea2KQ4InXTpPe0LoIOHGJCwf/
M7UN5SNLENd1f3i/JHaP8JXaiNp4PCzHELkfMo3sPQ10sSLRy1NwZgR5nCno0AvT
Ul2n/OFC737kA6mLM4XRxwvtzssTjTEwqMkqlIKwLTnPc5aGOfrrmPGqU06JLPxU
5ohCGbgBTbFMClSMQSfDaM67bd5lq3CMIERZRLH++KWilKkzH2FLV+gl0iv3NMyz
xjGHPB6tqTSqIRUy2g9Ax92uXffMGu8xh8zGE+00BE3GkINps3law2MbpuNRA0Us
wwbt4kp6vj4TVhVaPjvK3DGP6GrmIUne+dEevKFDA5xlSms9McraziQvaFNG7rTg
16TLuL0oSpmwKmz8ljuyg2NclnpAZSuPIYJSVzFAD9gh/uFALWpmOSuOBWRbhSvH
wnZC+yrtshJGDQ4fKa2OrBAGTNnFWZro08ZnWNTZYVimHWMc8sY67BZnCcMwrrqn
AwfNxI2DvssM3ogT1CE5kGzJRqWEfYbskTxWDTiwrAKV+iFPpv+QKjYKzMch64Bu
fTl6MGV0todlSYsuCWwSVzRaliSb9c0ZCTlwjq4tt19vPmbUrZjzaR5HZeAVmrlH
bRKnVPlz9mYoziaAkHx5XTPKxOZBiXcvP7GRMif57xCKfe3yRh/EkM8ORNM0jxFU
a+pvrD6kA7soTYG4V3tAGf2GY7vaWr0ezjwhSf9i9SC9GMwxAFIf8gySGKnpmSkn
mU+wBen+zHm//kC/oILiCmaATCF/IGIXmL6As7tp4rc6ksA2qAlM/Fz0ajwrpQTl
vepES9Rpxe7FUC5UNP9/pMXMNyegl7Eu3J3WL+GEMKK5JlF9IqnWr9R3rrwekjgM
b9BeNWrbkCK8Xwj/pUGNuhA39N8bJW+2F3cfCskGbd+d9CNJ8z1EDl4rxmLcsel4
ftKwAiuuiS2oEXO8oRZBZaYnhLkgn7I42P23HTGvtCxwQepJFQWoDCCrkPP2sCy9
fWfZXPEZun6BSz+W3k8KNb1nlo1HXpmhHB8sDvTkPw3B04RGST54dfabkVLGepr0
IiHd3mCY1CJ7pYAQGWu+7JIc7I+WRCS2FDtQp5Hqf8Hg5zzBdi+0ff80SeWGX4OY
3bH8tinXOV4B3D0YMaB8x/FiJ6T1jSpmSsc7/UeK6QHqJPFSa6WIaRU6qmwawnjR
F8H7w5jQjISV0v0LlVRqVfC0Vth7BioJXOyckJzchtM+vnX/OtNDp2i2FioUYu4n
2AhMizt6+x69sK7I0D6snPDI+kqd8Qyt+FUppEn759mKnKnUTicu59+Pm6oZDmna
6HmMb5JHHiL2NhFTdIqNQXz1/a7HB867UmZc6Fn/unRI4M+Ek/jyDmp2JqC3s0F6
oBQQaf0QbG2le+xYmyEBzsOQyMCnh6EiN+liz1pPUzdhR5E0qzMdzDgLVHDOm6WR
Gpkovjc9orkqnjIVNehQlJ2p/1NLAHejC5MnDkPXOoqgaRmcpAX+hvMlyNO+wbOd
cU0hXWO1dzBw00ZtxTnMJjTqADyq2aNleXcJd2wdGP0k4x7J6uWcdx0ObR7fOPTt
6CE2Cs0eV3e0tq++kFOoaxH/JBGn8XhN+mVwbWaYLHVw1c8CWQJk3gf8erdixyRI
RCAMxqM6xFuyHDiKpO92bjHit6zmDNe/48bscqq/Up+nvi7EcX4dUrLGvaC4IymA
DXqwK8GeKNvlaHGNHfyvYmEiGVe4YkNObnd8zSiO4ffHCUKcB3g/DjhjKSR88l+Z
w3Px1D6JVV/r62FJwAW3N3UHcqCZdfy2hnAfCC1q98Sd3PnHTPuNe8iJj3BehKus
f80S2Ki9UKBks/FSm8GALKhRmICUjpiiCN6Npd6AxK1y1+Nma0hvM4bjHWGgKewz
70u/JJ3GRohpyZmrVH47XFJoYYVFP/FZaSPuWd82vYCjDF1BN5P9S+r4+UURLt6P
pXsV+8R9YfAcwIrE8sg52RNGRwsAsBG/vtL85R7THtKT1SiJ8YePtslSOdvlsHAv
aZQAMQz26MfFKSm7Yi/lnv/W39fSvAzVUebaz+ykZH3O3qUjNiCxrCrTXeSH7gRH
tXgHrr+BI8IqMPtUczCAL52gggfA2bgrFfuo0PdDwouxXzy8M/2oMAchWyE4Ck2P
opB/sRvw3DA2Hjtvt9WGN9S9LYdKlv3mfcXXMBWu3GwfrzZomv+LZZ5ixf6D7D/o
FYLGTP6WUDYx/32JKqG8mGI3Bh2aGp6iC8zo3GZNuULtW0gdqabibnfOsR8E/RtQ
zWDcDDeZ5Soe9qLX19PsmMInDuBUG5N4KQcsoD1Nx9Bp76dzfuVM8+vU6cZhb4E0
5lDQaMAF04x2A1jiSa1fKSngGm8KFnW0g/DP25UpNa0XNK40rinC/PWJJy3emNCq
Esqdhfq4qkXsbgN+/r4r462g5IwVIdQpIBp1PqEugjr5/wnJ1dCEvjGloLMoFsmg
+12SuJVfIdKZb5QBcTqYgeu5lCF2nKt+3pG6xHm3IrfVGvJgrgB3Zddyw7157TQr
aNP6ufS85myTzyOXtF67vofANShSJb27QSokZZfW7pgKngpgi8oatyU187CDTMhb
RHTSuudSbuypTmYme22sBzSEnYN9fIs6s66uj1osdida9lwGb5litswanFwXohBN
TaP/Bp2LdSRC8LkB9lzlo6zW/dXdX8XQr/OFknj2pJmpkMsNbuoVflyZTHzm602Y
H8KMR0t5rbsEsil5bN8iOmf9EmgsYey0rJ/SRqrX8uvd9NsFCNWNlqCd3rYjG4xi
9Bb9+W/FnPhcF63e9vlgC4M1WH2I1e36WT6XkCz7/CrWZQkqGbdJm2KKzdHR3nIH
54l9xkxiP2VmoEhTbF77bzwnFH7jrmygmxT5no58LNucwZgT2RzbaK/K6bFMgIJN
PMOK8cFz7WeUgFgsFf7n6lmmvtmH0m+2iTOuW3Bl1BphUBYx7kxf6B/pLn3XHK1Y
VwS2ed76CwQznAQJVzS3Z/kHssBygU7FOYsyQLgBpDrSF+XI7tCXBkAlsPB86QMQ
1oja0brL9O1La+JbaiXqm9ks7Ctl8NWGY+zZY/sWAQgB81pp/6yAvqczg2JBOdi7
C4fvgRGpF3qQhPEG6aIQcrcNocSwz6fsiOFijsl1ZprQx0Alt0ZnbeG8CVtzzQBy
ptO/tS33uYa9NNzCj8f9pKCr6aDBOfFEpbOHUZtXZa8j4azJNfoW9gRUndkgYvKq
YaYk/W/sIHcbPix+UEWXGLtiNwiTaZTQAH78SeNdiMa6kvzhKDMTfDlGSYA6/gf2
gnyhtSjSrhbI7dh1Gdvi0y3sFYTYjINjE6cU/0P+L+fE4oS1tG0gvOzQcO3d86VD
lu0fg/E0PcGCEhlvvAFDYH/qvphTN+chuVk0xgWs/hOrh7Lt/jC0McmdGSnoe8DF
DL8OxZzKNEZF5x7hzuvWBQeUz6fBFqnzfTBh5cZGBu8wpZPH44HnTExO45YFAP9X
I5Zwxbv8pyHKrgXsdJTZGlM/Kmb1IojwOMQ/CReBmuecajQMXE4ZS4wakS1GHBR7
odP6FYoXJH83CwCr+iVJZFX5Y0t/Sm/uQELhm8gvMRTu0bAFYJK/p6gXYsSvSBis
pNQ+HaLWccCkEr+cjyQ2yJTGv57yTyCt88DeqtpKMlNdodF0TDRUGkxHzESVCN8A
OrTN0OkONN5oEiXbAM1Dfb8ILwLHgQO6UVJt13sH0soe+0L2m4jn082MNJec96b1
hCevfe3Soscm1/Pkrn1cHxaDEF6Ur+IQve9nTKeP9U+Ydkl5cd9Q3kwxHxPS+uUA
YJMD3XAeg2PYcdfxQZhL75vf7VZhAuKqi5NGLTyzKCEqIjmhCEUXbN6V4dzDzA62
pGBdVUCdpjGLpp2itE22dSFhr0uYOSb2ihux6DW4S2q6msz3owUyepfa8q+21Cap
TxZyiHLlCCjO8/h7CXWn4CjbqQUOhUPkS7NOMdrkkVCfFwjBMDaDSikkGAyzuAUT
w3Ea7Vhy3NCEE6HZOuS7fxM3+Q0jMGq6r19XjPiAfa+hiJohdcbmzFidNBXHG3Y3
rBb4QporO3jL43D4bWuQAm/sFObTlrpJD2G092ygw8+NlbXll38HgxQJftDbA7vY
ZuStrw6hfmyD7yixI51xLmxuhdF2WHdY12M8Euk/l++/y5729meSIkaskNqFdhi1
FWGGuSsbsK7QdM1iOESjB1ufSovIcEiSed/EY6VLsXPDqxzns31Lc9iYmzfZXr5u
Yo/xz3A+1i0hmwgzUkCZjNNfyDuNl8D9HLOZRZkOc9w21iPKy352H86iKAkgwfVZ
jQQ7uKdMIn+9aGrlhvKc6SG3QEmxZBbbeKspZdSMdpH58j/mZ0FgXwL1wyMMHftS
hiH6edEV5rPgf9Q9YkUFCSxp8m9pen+KURexCJUM8KplZtbgaVE5FeYyZzkFWIMx
rNLzK1UeZQf7c3Skdemoiu7hQZSopcX7S76ZLht0WcMPV7aAp7a/SDU63oeT4Ni+
Ojw2d34cLcfzRyqFNpMWHtO6l2EeLwR/XDT8Y8OzMRTU3LLHFHxxrI0VuxbjtThd
pdNDhB4TI33TjqfMsTOya/nJCZSHiImKARJcFufFO8KRCAzSFCwAlyPCfXR7mSw9
gmmh/teW/jPTDEBWsCWBUuz4WZ8yD/HZIijlrbrQR2oRLbQl94QipwPv/OjxISK2
6lve4SXCuSp7mQnaKdr/92IxltIiZEIm5BIhB1otc/GGkx9p8G9Ii2n0gCuj0n8h
FKv7wel8N+N1XmIP3dD+66/GuRZctSnJNtjOVv/hpVQQ5+TgeASxEuGMvEafnz03
vmG0V6zZSWrHbB6zvzDW+usSNvkElBlL5g23YQ7Q6PVeJ99lrSTvNXcYY17fOEXi
O1YPRRYo1QRISgg4ZYZgIQ1Yl1xuPaHnL/ruffkEexONDo5hNxTRK19CT328RtmY
7I/ls+fVYfY+CFTfE28DSQRKAK7CN9B93FoY+C0B/KWeCHmQygyAGs9fg6Pe2xIN
B3nLDGHCa4JFEGiqFwArCzjzYDFD5gshnUKXCcUMmtWD05cvM7ghVWq6eS642Tgr
IHZA6XGzL6USEfDh9wrl96/TIQRh1f1D7+30QLswzg2OiRfbOK6ZKB9HcNXzFiOF
/S9Ix0ej6K+/93HTihQ0r1j1XSIi56r7rLSvIpLrKxurlTqlNnteJ0gufLTO5TLt
Uj8Bd4vwXoDQKc+EfilZBctE+0Od8m6WUPPEPP7XtShwNn7V54a6HqkprzLXhBZ5
nbIleK3nvh0PslbFsSPXDqJ4q7Eek/OX+BTZ3klSGBEezePsOyr0OrnxSaC8MF3V
lDKzcr6XwOJMmLQOjlPt7KdCejQ3LynDdB49DumduIQegsQqRq4+KW9SPGq+Ojcr
StzgySn1ntl/jEMm/ugw/8+sH87dC/fYFHF6AAr4G0gvlD2nPB2PFaeSeYmy3lXd
PqjrWT860iqI/DeVVXBS+I0wZdXa+IblEqotygrkONn67w93o751ZZ+ijfk4WDN4
bfr5nkrUCjFZoR8Bf6uj8CDQXT6/O8zu5mMmcv29w654XZq2I0ji23ioUEaRo76v
9gbEbH8w+nPiH3DtEzpJ/o+AKk8OujZGPS4wCQIIbShuowCXyMlmeDcBioGsmKNO
njWqb/+OL4wkAHjWEPMnNflz0B3hZnCn7ENYqcbZadY42y0qUikIKLnPZaU5I3sO
qLxGmDxgmDZThHmDTppGZTlI7xWqcSWMQ6VVdnptoSfzHf9DVf6SNcLFfbk2LY5u
CjP7AXgUN92Xv/sXTE3q2SxnOvN9Q9IVzyLUj92dzdWh3ozk5qtbE60e/NTzsqrN
ETgcdGExeOK3rCOf+Ug/ofThgzMkpUYxRu7xGCwTD8EV1gGN+IPiYNqGWQhZqaV6
pcwrtiZrYANtLnOMlR0fdNnqC6b51IWQ6s7Xuwrv2Wm0U2ZVi4bGS6wC1TsT3twj
VNpzxvnD2pkCxi8Se4Ujb99O/9sBFpfd8OuleBwrfdpeD9m2X9dBioFl3W3vJdAn
dCC351YOTgZMvvesQsTQ/uJygAvBf4OSP8+qMWsU2l+TxreeAyZIUb3MXL011Toa
XSAhRg4iD//LzAXOHIohJBO11x8VDmq43tUCUlo+STdTqUVwI/CsZOMckb21Drt5
MVtADsJMgKRnfiyf2fZfhbO/Xyr8IH8fSltc1Go6dyGxiIufkZfCbzpuaxFMlt59
07OY/TLgiQPpTjor2PBhxv8LGBnIjCIsA8rvwOypSKaub9mLfaN0yqTN1MHX+xgT
jB6Zoo5q0A+/eE31A7WE+Cz9wIQrWZdXKG04ssYXWKa6CIlOqeWahsKfYBPCSmti
/bnqwlHzu6arJovpeaexFfwmjqadJXgIJqQx/bfUUpuGUWzwNcH992SkJs7je9A/
nI94fH8dgcRUDL2HVugGwbW5VzA1iSCNpPv4HsPNgljHD6CCWvLw4lmFucWl6s3q
g0Pm/knh60bjHG97UczZUNgwf0GOh9WD5P524mgxcgnZA1Rq/cRznuB5vvjZwBie
gpGmkLhb7NfQdTNIevYEew5rl6AJB6GEecGhVBPSSd3qMlHjKS7cjbYwvJGLM6Pu
cLn6H+R8XXJ6bql1duvN9xpjicT2pLODC7Op9GJXZ6BTv19URzBrZeRhnRJaQ9qL
yzw4WMjYNQ9TF07/64yA8VLMr+OUFo7a8ium88oX5qZ0HWUs2nDkUyEQJGd47sDF
Gm1QY1ozcabKcA3JtkLjmFvGsiFdNYMuguVlOuEoXdoopoBsr8dIsjKdNtSX0PG8
Zfbjb7Ze4lncfuNOs+5gehWhRfYlWlFSap1GyH/SjD9QaGABkis/3qeXLopLczQI
OSqd8U7sncVtPfAncIOcZ18jVVGDzEjGqs7AU0NiQx6ItAox3bDzvS4eGF8PAXsZ
ApgWIPD1w0tEfwtdJuATPC7K3HW27mZ7NccJODKqFCFVvwVd2uR8yQ7K8BjbUu51
u3Sz6yjjm/xlvCB/KSNOXDWDPOm1OKifOPSfSDVLyuGfmS7G0w+iV6sYiixuhQ6u
0l2QwfpfpxBe6sfFota3p963oiWGsiwnUdc3LwSve4bHOOP/z1JlGqkQOpcJMO6X
5MM6qik+ByCir111fesE3FjSiHw6kiY7UXw9tvkkX/WkE7R05nNPx2xasAWyTAeu
EKBjd6EAS7dpiONh6OFQIvXzkZl05k9SXPeIto8GJNhJppeacXD5P7IGo7D+q3Oo
0zttQYSAuWIH7fWAKGyUV+xk0OgYZHBaMZodeT4Hso8Zxg/hEqYBGIV8pDzoq0tU
ZzQLY5teVrGuiL/PacxEw92WFgfSJQnGv2hXN7v8ZDoYg+QrQlJwBIo8dRPYTjhK
/YY8z9QbngGABXghABiUotZAtYVXvTmgeF3nJH61Mqg54R0DcsWV2/XESXA5+jIm
uvTs5urVsfiBhB/zeMISwcSKW0rw1hS0lNQE0vGaNKGxYquAtvN14USFiNIcsRax
BRcC2upMf7kB40N5OOgfAbRFD+sJPeHej33nkB4j6hcNI1//6Jn7x0EPpdNZvXFJ
Hr1b2NI8gNmEvaJbfvZWYe/Sayh7fB4QTDLq5v5nWwNNz5fA91+0s4X40Fx5dkVK
syBYEdbD7ZQBBA96FPu8RLSB4EeSnAmBeVAdTFXWlwZFk+5qcw+vZhblv8QXLQ7q
OXLYO4tLXTRYurM/gjeMqXsRbZntAdF7A0v7k8IFtZ8Wc476HtYv8qG7f8U5KO2k
ZdtLyPHGUyHLjZn6eTl6EATpnnfb6CHHyAoNsaU3OlSiOOlZYWkhQrevbKIOca6v
B7TheET6dqV/JERyTPZouSkaJKtUmkK0K4z1N3CMVrk8qZpskM+ugaQEV8mMAbMl
pjCfrG99yW97hhyPlHqkYaB14whb68jAZQCk3K7FkGNPlcxYRYvp2qzlWP+ZBbFA
60WE7+rVbSms55oYJ9IQvfjAcqIRkUzqkayjt5J2WqvAnArpwJMxVRatzdnMQaeE
k1eImvE1BJQF532TjQfyOZK63Qpv1NdtVUKTi3a7gC/nh1MGKKfRQEeIc/jI4S9k
N1Xqs+MOAOs0vqVUr01j9V0qawQWzpRVMVTP31QMzMa0KUQDJGNygKz4NzmMxuIT
NTIyLfhLNzqyZn5/W4EkhV/+3l4sLbCMgEI9KaKSCQecjy0n4ynrsfK6rLrO8ana
NL3mtUiN3qZfqABt9GCJpJcedC1Sfby5yvn9maYJzglsMAhacFOfjj+ZIIumDErg
CDfgjjbE8ECceEOfQt4m4DPdtOVMxFPgl+j8fNZs7F3SiprC9CVKnBw+tFEIwRHe
rPvP526HofXOjoGEg2Sr8XD3lV/Jj/o2qxHTyWb4PllGOBj1t8WrpCbdNI5mP8Qj
9RBySeoDRyNE6Iw+Jz0p57RY35owv7IBXntXMIACXSGAgwvHoxmQdjqnJe07pbSP
wXb7odpNZDy3IzIgHz46XwIiGjJlGFbzgjG7rhO5tJ+t3jPaq6I2dnIXe5mKyX27
VD9aZh9052AozVpN3RSu+afj9H7NsRdxB7cLN/LwItwOPdzHm22nlFuzxwLGZJmu
AdAI4xXoNkobCDkArNPPskEKSMAIddDbvJEUPCbVaafP8U5erzwua1MFItZbwuiC
e4stOhk0UstHlj2+mE4aHmDUDLaRRz6Mfxr1l7V4BHlg+YkNYioQuZL6ASf8bzqm
d35sbZ2lstKW7jciHmB2H/dpthSH6LZuUwCiund8+qU8XXMJSQnBRAp7gVgX1uZ7
leJMgtD7epTqcMbLOtX1/dFhre+wRuZr3gVImmfQsmfCrSUHrjkQ0H4ByoRkrlrc
jH1uCiOwAnUNJRsyuibAPg4fVCoBGkEp3WbcLqVhBtwyH+6p+VGXDDd6rhqH4FUs
u+GQBjy2dQfSJqk1czgxVhdmETXQdncFnVwCWP9QcGezmI77E8SWlPN1E72DaWQR
YIn6orx3Ycgh71OdPlOpen+oolqwkrLyMtIEQgf4NW5HCsSEK2fKHSiMajCNLGJV
Hej9qEaLq9I3kK2ZVKd5VD2UfLb4PaM/yjrFlcerR+lM0PGkXAK4eeGnyT4QruPb
+lMOoupmCaD8g/3Gm4ugVDSDVQyxG05ygvYEi2GRwz7mH16n5oapKrSbMdxoL+gS
6QU9oyrzsoI8viaSTuUeVaXvl4YxdfuMs6E4/b7Suyq+NGMMo4xyDO8Ng6XAP4TJ
/2xAgf6Ku9BEVQ6IzykXgcq41jpXLTnTZ0x7qLRbplyl8VfdETNo4mK+Rwh7YTZB
mv0N+/D0y667sZmMdS5rxEuq7mmpoK4ZMJCVhOKPHqb4g+ucGuYAFZOB5BsHLNuQ
3oFk92L6d4x/UH2P50jGCeNEST77e+NZPj7U00gZvvGQg5EoO1Zu8Gco6lkoSR7K
OzeOPn7rVVUXt1nyf8sydC4iBc5PjHjJfKuTVn02JqE4JCJ4QjGX04jJ2qfTvezf
T8jHyZJsbO9Qgi5wLTuphqZajyTXz+5HpZIccgl0gizztrJOIx8Kb90LcfvcyX8u
kf2EFDXuL+HIuSubmm3FbJ63Yqh9GO1Vlk7EvwJFrDr7EOIEa6REJDLPzsctv+Lj
280jAbq7XOfnttXY6lJ5LjKdGT3PhZo1oD9DrZHi4FbhadVs9iIuBwgP/Jk+6oxV
tLjwVrsGdXmoGGlh4M0MfSEyRP8gP0HL75HBklVrjMsA6qJV3xtir3ghMclKTB77
izut3oynB1kF0aaoZHusfrlDW3AiPkEeKOW/dr3liAmqjgmr1er58bX9pUV42WdY
4tGCj7cJd14YdA1Vcj47oDL9if/AV8FpQwM51Qq55J0QDwvkhXYzToVACeQv/mn4
xbf3W5+tNY0PIiIH2QcU72c6xQXxAoSc5BKBUmBvC48w4T7MSF7X59vNs0Q50qvz
sCxb/6l/ww0r2pPWl19sYKmWyKcSKd3JOBPmN6Ad7FoycjxC0C4fdSJTEakg3wLV
tZBoCJke/j3lYUlyL0aej/lr/aWCxfqE/4Jgs7K08XHzXGo9Ke4Uhxi1Fqr5MAwX
qD63r0edfdewJVJiyYeBbWByEvqZGzeFZvS9ZjSq5saP1m4iOFnkBLx2BbJmUnRU
LrAQIjW1TvzZNd/niQRXSn4rVN2L1vHRQjiskW0G29ag9eQHzQkL7tU9jijuIZsq
IV9GpTkhZASRXQG2ROozl4x0/HSD6DvaE8UfuBAOpPgjNLXSmWSCWie9yoAS+bmD
326McgDbt/hAPkUSzZrAVtmoBPr/j7eGglsrNBrOG4ee78oQi+vGCD3AUAsWZtsx
0ADfMB/NErJXB/YZBRkDKw1eHCcrwP1xFkzUQtndwCg5mnTQu9sC/VgJg/DW2vpZ
lzFaMb2+oCAiO7rhL99yYgWk9ZC7Hx9dFeKgkyrkoHgYrL7Lf3fLNNBAofkHv6AF
01T3b/QUK4c1RdTwc/SyyjXnJDkMQ807jZykJ+8gW0mmbGnpLQdL6eEZyuVrbcZs
byYJ5I1DgA3IHulbILKI7ml7jKGV1G4+PH5VBtkgRaUiFakeHcllJwDKQaTuaO50
avPRSnapL0Pc9wCnBSkhUwFN4OC4XOn2UL4TqGvsj+n9+e/RFA/044v+LzBf9za1
7/QuGzrQ09p8ipxSlVKnsys5iVvnrAMzX2VbmK73TzVjyCRjLW0PUlWXyETKFdZ9
pqMrXx7G3vJ3dzci2CABYJ0YomTKLJUssAIh4ZY+rlzTIXv5nriuB/uc1TzLILAW
r6HK7V6Rs37WIPjOX+mTnpE1QV8EdfB5YQjzqe8Se6OjFrKwThMVAX1dDF7u5shy
3+VvLNyndTrkwl/mngn5TgtwhSmXZyRJzZNRkZVO6Msn/cGV2E1Q4rcFgViE00yD
KaJdLsgkTDHY/on53YO0TNRUG1iUHN+EdEPyos8McLwlvxNHM5U27d1CpacAPHwD
BIV7Zh0iNPGDm6c6BwI13CqTodZu27B/RM0wj2vNLaHwu+4eSqi8fOyULftHyvcK
4PTSsWszFqUjPyn+Y4kqR5pUGABup3+7wF9fKqj/ayVxwzHTUhHp+n1xfqv3y9By
EWw3EKadSk87BE6xFgNl7MiMSiyNbTbF8/WlJ0ToAnUq2gYT6eGoH0J9XHSJg7MN
qKnvHSBZqQbD/LwVqC/N6KQALiwS7YnsjkkZZECmAghbGU59dzw3JBmnhOlVJsXH
eIE4OPFaQZ/yD7HU9PosbxD7hAB+pGwBgMCCpJDzIT9hWCKL5aadWXLae08YYmkw
nyzI6ufq3EORfZLUrgHLoEwVNbhvBE7g0sz134xWFCLBSvmZ4caJ/+8Uv+lcIBLl
BaSGD4L/lTfDom4VXVR2Nn87xbunQZgMIqjwX9G/fCPB6MELBAMqKjDZU4z1xpA4
X6NXmWHd9ppPuTP9VuaWqSzSWrMT+YegqLosqTpaGHyM0Sw7zne4j5lXjtG0kUyW
NMJlNOrdx8R5s3slgKJVuL2WabXwvP1ftClGSBeeIrHbyFX4IlMLSsP6HIR4XBru
IFThT6OUbhSd9tvdXi6ziM//DVKrNlSJ9xyUZ3p5umwMNouNmOiFCIR2tUhAbhCI
+xI0Qjd8Z836Z82qdb++M3WvW2OdxHdgV9EqGmDROpBllozVyayN9PrTmTuQSmXP
LqhezRTWK8q0uCzI6CEvFARTFVwmnrjxsSibWcFPYE9dTqf2RMoh9ueo+zJv6jk7
TPoBhEAmRnr3R5rOErw4j4xybzCczGwZDQmqdS2jBg/jfWygajV9iZmkbMEYprQu
AIaVrAMZwN705mL8Exo/NttdAta/ySrQWU3rY4g6fgiH46sLZgOrrDGVlgQFhSQ1
9Y+ZN+VDZBzM/6ec4nz830b9IgaL3Ry96CsaLxHLS65oL4eis+adSQtIcq+ATXwg
vKK2DU/3RSz5sYJ+3e7aWrNxLs87W6vJbQx6If3mp6g3kAcqwxjzQPp6ptYcDmkf
jkrrpXiji4+mE/NT8ujf1jmIj+xIHBS9FgNksqqPChWmPypC+A3x866981qVDNZn
LQ+iC//JmisJO+1OqWy6v6evw7ZS9zKf70vLdTgwRIXPlhwUrUIH2S8r+UfO4bVl
PUpajJq1q6HSrvUbeRRHqW3d0Oi0KVGFLGVODLlQudzq0MyPtE1sWeg8A8JNeuDQ
3hMWdqKlUlYwSRpZsSII2gE8gkDR/3CCUSno5EPHIQv4DCc0QTNfq3yBbWRlSkFQ
VpxLtUw67K3xDZMCp59ZA0xGO6h+fqnq8WQ9rwxWJFhgy7V58rTuvC9c9s6LQI6z
R0GG3OdJI2mlXFjl0uY70WM5plTh2oJN/JuXL2zwFz6fCrY622dvDjsqs5aHeZWu
8qECIXSdzaIjk6wK/aZrb+9M0c1bTw0sFsyMC6EHj46wJnIEOsa9Z6bEAbmY+a0l
PjQVpbJ5pAaoemlCso24p8U0ukNXbY8xlzq9unld6VNYAV3g4WzNZ6OhsTq1pqMB
KFCQznfgd20Ui7FyBDLDMCPRQIdKCbPCp/5HrIjvNAanU8VAgvDOHhl00x/jVAuZ
TvQhOngpogXoD2Cd1xDHb/TvpKjOmBFGMFlwNe0pHWJA159F0PAYaODnhb5E99U0
AmauYzEm7GrN0lLLwdm7fZbbkyutalz3BsSVdnFds1mDggAwsg6QOA7HnfBAwb//
5NRuADXplsblLXM+2GiDb/QpocnVMVjqDOgE55NfxWmeeLbLdFaMj9i6YYfAcBnW
RZsfgljFzVvOVuEQ1/X9acEro9dvrKDLlU9GHPoeEHvICxkXtcRDIV1Fqej6tcRr
3pLDbM4jJ3YTZNfzaPZxKT+AcYCiC8Wq/fmK+s62JXmPAft99yzczsLAJNoBUtmK
CzvCiUmfNou4to0NJXeyLJKoMBtfZUaryV0+6Wecr4PRoedmXvecgMXktp0B9iHe
FywDlz4QYn91y9aFo1w9gyaMIAfHJqnTndtjrtJ57nE3IRVWSinLM/+BRVRsevSG
AQInBkMVOsnaSnKh0HimikhZ9E4/1MQR/XpAlPYMCci8TnAic6Lp+QzEmKL1AbMi
KFYm6AzD5QZVSGpH/ZXxyW9/Ok1VGNWaOpVMxBisQQ4zy6uKWUyaxqFbR2qAc9Q9
uIKGJnL3QmQqECyybYqZNqXvyQ635IkFnvkrKBdhHUkESAdUW/E9fe3cUtEOsTK1
gkdPWaqePLwMjC8AyekLQzgZbSwNG8LSjOC8O8ls4xpneF+Y49pc3XU3/tXmfpur
rMXWtcv2wLk2RW48La6WMy4II6W1qiBtCPQDNnunWafOakLGnwMqsxwyelhKnRWr
QQmnz7kSQDL6iH8PrFG7KOsmINa2/aSp0PZiNsNZnsXGYeCu4mSKuPmTYFeD9DaO
NcjHexXzzeY+4/Px6IHzt3Y6oB8kCGWG7So+LOugY78w+HyqVVaA7tn/lVeBoa7M
x0wX87UC2th/pxCZKzs9TPWonSKGbR4S3+whNU3D/m+6lNUqz+J01nSUuZpVp/sZ
cmPD8h0ecrw179AjGS6dMXJxKMXyWnTQs9zAfWBxTonKiqx+f0aoAWlpz2b25iXR
jrIxN6+wXuj2Zg//PTFJRB/QvL7t8EOvT5bPLtQ2fkSbJAsQ5Pw0gaxxB3bUx7Rg
1r0RP9FYbQMFMFGKdllRA3m8BxjAaa7zreH0h3TpxqLvIUyeFY90S8mYRcJ4S42Z
luU8ISpmwV37WxgBgADo7VrL34BBDLQh2HTKkX1TQNPcSRGlXAbGkVt5apORJt3W
g0CvZVsBNQip1SUp+YYbsgrwRyOXC22T2MTKw0I+DUvmWiOeqBm50W7SdUtw86QL
/jqWk47SOkTu1rAoNKSBp9Fox8r3NzDTTFDnJpbnTNo2XrnP2rmKpIlz0xTIWHeJ
7LitiGvX8mKOKyXI5SNlqxyer4zgQexSOjFgPqVFCzzZYGLVvnIM+EsdmR7ZRYLK
y9ImTCxR5W6hONfGzE7BLJ7dSz6aVHcSEIzW3MDYHhqo89ED/4jQox3/QVJDayFV
M/cAhxdI+oTlNQapN7VOUjnjPydK9h7ukOO79xJPtwxcfNUop8+cEFHp9grPIiYj
DSmRL9sKsT5Xa0RvBqiyqmH1SiueSmdcJwhE66lHy+/IdbaGVMkYOpfGWJ37qIZb
ucSuVPOcagvZtVeDdRNxwdyF9oOTB9vkwS+I5W557hb0nSNZ5dl1T2XGzE+oCD46
QzYp/w63OxlKUtnI2z2Gpn25JFhXNeHPPszfafrOD+bdCTxDp8SGR7xZo1VbMCyG
rpQjGapJLBlol1VkcgXrs5Aq/kEZhn5kILcULFXY/tYg+PYSjPgB7GEzjMF8aqoz
9nJzQsOKX/LJTOnyz11UhrY36Pt0IFXBQbu3eStGChMBT6xG1w8SDR5CqQdbM4ad
C86R2tmtiXdglyVWDSBZbajTxFUXyQ+3EsxC/k+/5g9bhsg2a8SgFR1XUA/uCwjH
qJ0paY3lMcKxQyX2mfIhODnLh6EdzRUOjTqc4Ed8pi7xtDxzespG4s1L+A5CBqZF
mzBmfsVH4tJNAPxw6lBEFqEzKQJS97UgYT1C2ACucEV4amKr34dfb0rMnjeC/j1H
u/vN9uMsPnFE9zW+vxVuDIks3pXewIFTGKZ0jc5OAuyZh7bpL48S1MNttTW6dl0g
4eyLx1HKVgKCZCcb+zZm+5zWrO8GI+1cJ0aVIIuw3e1zIxG4MV0WUhaEmcPd2eIZ
w05ubHgFwJ2uRCHbu81q7bS3nkCYEBFKmkzjR7aMegOmbkz9H17XKEZhP91UoO3z
WOSXdXnSrmEI4zB0V3topTKHS+//tvAphcu7L4Yfc1V86kNmwIg2w+TdA0xDZWNl
hHnLvxZP3+jhnTlOIVc1ZeNkINGdxIZnAOBR0ZJcnw8O0nC38xHxo0ROVcr105jD
IvqaNzgsGt/qKWQulbNhYnV2jSwwbq86cRh2K16kwwG6XYFIM9trShDLJ+c6UdMD
pMPXimjSdD6IrcWTL48yupox9musRljt3SCdK3tfdVnOTk101Zd8E3YV/h7Wtp1i
mhqOO8xJW1qaiAtQZlbcSU5p9HhvTni3YELEWIp77Z7cz/vOrm3Euxs35Q2iMjh/
uhdGwkkBxICWzqPA31J4PRMT0HJasX7GXw1J0n6zegwSvjY7jWvrmH5EavWtZQtZ
bNLU6w3w1pDhlmNHpnJ5ftk3NySeg7AtTUY8jGyKiTpJBTnvqEBNMsJhMR7HS6X6
l0MYtCGgU/MlgX1WkcqZ8yw98rUk+T3L2QIRVzv2PPKtES0b9WitKDTTw5YU+cme
ymuoGnl7lpjxfRuf5BrUJm5Z+/aDsruVZQfYeJULrgzoJpxizHxT1fsLD9z0RPP9
PbY+Xb21OqFiq+VNL2Zdz86RXGHcOhf0JowvbKQEdch1hyJXbHqbs6hGfw1MmMfR
Z3Q2Bf/G1HuRHvnYJxkCX5fV9Dmr80IxSBu8ORZT+opz+WPso8J4JU/AeWDpops7
xyI1w9xQGUwdmWwRsIymBSBkYl1LtvB5V1RijgaDuOKI3ntdahrZlw+kgwfhwjAk
toQLCCaH0ELu1EBIoMmjrWHgRN0G2VOIMYrunEAkijflwfh8a15rhouIAMGW5Hl6
a4/NPd8DGvpF1/lRq31VrxShZM4w4a1bhMlKhnZ8zI3Ke/wY3/7FXh0iEAlmE+4q
P4tmHhqdZ+Vz2XCfJBpUQcsldYI7lW5g7vupBZlkYK9ovhtVNakKDq0+j+zf+56/
b9+i4AI1Yvl9C6s3IOSMBp/L8O5+KlEQXScCCigEMZdG+VRSpOq7MOsX+9twU4Mf
3Uz+R5bSnpl9l134l/RnJJfkjn28hq7cO9BA/4RPPD/5sUuBGR/B6AZ5sLAJFaSm
3Hnk2WvJqTXs7huMnihH5vdgPOiju1xSo+K9WDG+3ImBp6ij/CgxxTPbHgp+AoJV
VkmKYyLxumUCMiXO1DJsK2uRcPWeIe0VSnvIRcEVKjvhFtN3eUn/K9oqxBzvR8WE
r/xPeQDRsrbSUgu2QPLxdbcc+PmMJ6Ey7zRhe/iugWDRw4ZBOuAWFx7kBsHPFoZw
fG5XVDFU+5Sl0T3posXizxFBalx53vOpgfy75r4B0BzphSTtiY1bZO1UIKBcQkL2
fBBSjeYdwTbfUgqniFQs4qsYXiC/h3L4Ba/Fels826IimMyCKNanBo1Em43T4WYS
pdd/rzEcId/kMv45DlqgyOfZKY99dtXj0+lmYi/iADcVAnXg3YyfCLJ8qO2vyX+1
hnB8rpUm0vdGeTLsFmHvt+bR7W8dtdb6LTCC8DIqsst48XS+FIwDGuD+enGVfjRX
CZiLugZGxxCvGm19ckeb8JZv1kCDqvUr5V+Eyo0jp1RZjjuKxxAteN96puZhr6Q/
xOVhP8lnIsYf2UHG/54okG/ww+YjZsNyf6LTGC0fdrfdI3XbkI5CHmswG2XZu6aO
MHn/i6EuoAmhSfPxCpYql7cm1soH6Y3WlhfAXX9snf5aIDUwxOAckboSRYJirsQY
obClB16DFrx/prTKqPZByhxcOoLyjqZEPP2m4sHLNdY1sXlaYuC1wwz6JfvVLVnU
FJDA6GpTUALByZWoOVAwHAgQjv2qLwPKG9nrETTPKnxpyTYwTQoPUpzRbwzdkUyU
L9Tlfb8MWSw2l2jJkSnG83RvyEfmOETInMMUXdJzyEyaUBMnIDb9O8bpDmmVrl9H
D9WulymzOm7eRIR4+9uDr3rh1A1b6FNTQy2jkPGWMZRokfXWVbnbQV81A2/IZqGI
ETLNacvii0Dfkz+EXD1PgXWNRLGf9WZGYr4Ck0u2G1qvYIIcDgv7Ion/tIPG9Q1l
jUxJRkUNlOJJC4xyicTKw0ou0iUkGGx6GqZruTVB+Git9dqN+MFJJEEDme4OsBU+
VSJ6HSpiC950pYif04NRpOAbSnxBZ4c9nx61LArEStDQjfJBuSYyB4P8Qg7wqKCy
fJm4QiI55IjGNvWFAXXFjAB3/Oj8Ndde8k5bSG0SbeUViVewJd3dep9Bv9ZqSqEf
NMTsWjJujE/Yggoy4+WvBgllkQI8GW/Yq2FNWRVNrsiC5Ibt3M8vUav1PybtxtR8
9FZF8KpStP5XsBhraXyJNS30yhd6dnkEP9z7gLFtysoVCwuB1cfT1dPOw8OVRN47
W+yYXYECxHEyRt8fb9McCaq5zX4GogPwKlaxhg+K/FTnR7rfHotP/+wIz9vbUlHU
tOz+e1GFtCMJwbsLogxGtVyL0eFHR196PL5OjI6GjtnkxIf/28n3M45v3Gj74Er2
/YFE3FbkjG1c5VVdZgIPnCpmpJ9f2z7MQftWW30qcHX7exOzNwh5IiMUPN5FQQkM
HgGfRK1vdNQE0PJf9VoWVhfAKZ2opHmSPZ6b3pV8qXzZN/oOiJSueTroA/sov2R1
idLSmVGw/zT0RaFRoiVv+7O+wm9BPmw5s/uPYJ7djJUFp9LyMAV7gLdIGVVKiIfJ
7gmyWCAqC7jvERpIKW18M9WqFjVXK8AUBkgFi32He2qqUROTSSiJlZLGxRR61lfC
dglagc5wD+MfowZXHnbiKLRVAmJvRiWy+A529m3e5M5zHFoWlgmGpGh15yFpPs/Y
1TRQF+EeuInC4E3nto5u7IR694HA7tyKwoIw8zV19cCu73JjBS4skuU5AbT/Oa7V
eXw8wBgcRkmq3qKO4EvppN3Zibf2PKViLpPzZVXIEehlz09SLaFuY3M900RZVQ4Y
O+/+MVEEogA1xUOcjbKBVhCEXnUXd+s3p/ulteEqgZlT5Afwxm/NSKqqIlz7DeUI
qGddSHv8r4pO5ljyHTcSX4Ns4Xxu/qtlP1f94CZtHpM11jixnb2fkANlpYzvxCQa
0231n8A2QkJaRVYEOxg8V92z5L0zzrKcOYUhbMrYmp6ceVjxNczHKslnU0924/WK
XQ4/OhfI3qccPYyCHzMVJQDhiuEkSOVVxL/yqCbs7IQezlbSKzl8UVEL9KFgVm1t
Yj/Y0UViqmzfQwVRW09Ami8KMf4fe/IzaSjcmge4m2YjCIpSKkQsl4YZ9hAGL7jE
+0gBN9bqKfa1WHDrHAVvpRkQTiCyvEPBhL/6L0io4pLczrXMIuFRrBfDSK/I/co7
CgzWCGLKxAEdYF0MHWjIUfiTIRpIENpTaiIb8508PUgpAmCpvT9NccrWVHBm4UjR
u8C5G40IJzeuIdhmMQCsgHxkR624ESxeVS61/wi9X5F8vNVYyjqM4cOTs6WgeLyt
Xa3cuDrc8LfJVNGM1hy78XEyKJg7WfoheB0azepzfq2qhwhbVtL8af70WvnBS8yP
zreGPQut1WU1UGeTCaAxQMUhRVCv57oj1wgLa2awW2sazSalBVXv7WQMxPVf+71o
NLEm5ELcOxTELkP5zpA1JDhzsHGjTcXxLwr1mYHqT6os/ZZQgpZkhoQzLNXvPCRv
rZAGlsVtUxROVl0RqFM0a/jTo7LMsKVF0jvptRFy+fwFIH5D64JOd+3FI1uX7Db4
Vf86FD4dxoJLR27Jy8Hfd+kgO1iUyugoXxupI79+wLkbayqGWhAYnQmI6VFHz4F2
DYdFx+Wbid5O0Jl125JWuhyO0/O8IwEe3PSIzQHv5eLia33SAXgnvY1Q4QY8x1ZP
g3qG7VR14oyZBqIPjvraCUKL5FnE1PBaINhp/VzsiQ3SSr0zY44Kgy/gof16skFz
b2ElFFdqQ6ecH1hUmopGrCJ2g+X4+RkQ8aH0HLwJVxasOb2sOA1mbPg+OhhQsw7P
zE+0DSBd4bLH1U1DRhaH38lrFoBPBPah6O0/npDUxZYopLi6+Lgi44PFSIV2Nuqy
NCYonpERSA82xnKYZq9xTPzAl0/XQk5LhRdm/TIjGAi9eeYEpbH3eHnJHWgp5r1a
cMTSakLoFJ7q8p/qjZef2suY9Ht0llvNejN9klPgcrlpOako5cR6gMx5Gg3y92UZ
FXkD/IaYZN2t2ChN79n4CRRIRmYbMj31xVp/dcEvOrnzLw9OheCRv79XmdVyplRV
XMxrLwnJzdtBU4ali9T6A3PtXWxfnJiPHpDDOZl44o4JAdRo3ionEo+Ci4HHxW6w
MEpup/ovQ4uV0v8NOMLo8bndn15DZzNVjMjz33Vu5boOjS86fj87GQxa92WSGcNA
TdUx5T61c3GyGYS/qT1s1tbz1knIJ1ubexsgs0A4Z4OKONLxjHodhIsFh7gvkoe0
RfqvOGq/6aI8UMS0gDj/+Fzfyw46WrXVrI3r0s/xIcSNN3oHfSZfdeuNibXxU5zf
+gpY0zIALSIbS9zB/+Je8vyEwNYuzcX0sL0WNXv1+rayCUcfjgbfbDu3/1Qkglr7
lsU5hjpuaxIweVkA8lOu0hnzZj1X8jEja9xdnO/94pLTFipF0VIR38ES/0YNujJh
WEaMK4WrgKAXenKP9aPNOY+Rk6K/7hHTPClvezAv0YlweZ7y00wsyaPhxy5VnbcL
rYAMOMNg0WNAqdU3o6hvdhX1Y4m1tLJba0syOpN712gPSw6InJKX7bfOz8PRLwVm
+PDmfP8FOL0g5zJ6IkQ8rnSLAggPGx4WPw88nSSJFo4B85wHBZqehPtqzYYs204K
VY0jArEVW7ZmqzFfS0lyiD2cjyUAt3NQaKRlPBhV1Db4gAgxJlysWgv/n4D0Qmmm
cVPuK2QrF2nifYgzTSwD5Nhb+Af4aQNuiIr/NcwhnF6z7zfvTcsuRMu8JzeJGRaN
qH/W9Bz5lvExHzesXAxW0aAaIBtNjZ+2dt9YIgQU/nL79aTTW2wc/F6F6bY12s0m
hPfXQRJQCcORUkXUC9/AYO39v7KmVUbZdyATN55+cU8ux7QjMfmYekFUAP7HOV0N
4B9gG+YqrNMFwwX3AF4s69+I9HnuPEvsGNRZiRURub8vZxTi7wrp4m7wV2Ey52uk
EyB3g/j5mc81fWnQK0KVOUxXvwr4Xc6JJXu/EXtwVNqTe65drgwA9FbQ3y/4H7pV
4N48pwRsU5ZdNsB1xtS3tjK3Tso7ZaF9fSmdM2cgKq8Y0YiC6K19dqsiOsDK+U6P
qRlICPIAEVcEoGqBRfWAEUv7lf+kaNl4fI5+peY/BfyTCkpbdeX0pX+ZnE/DVL/d
1jZN7TefmkHi2up/YcRzrf9L4JESMgGbeE8ipP+83aKQaUsTyhwf2CaZ6ro7HtAL
bPjQ9YDi5I5MZeyfpTkxPe1EELnRU8m8knyT5Xv14KsadDNgHxiMpyDEhroy2ZFl
nJzbZWQqNa940NpryzFnhRPbR0xbCSNhfZ0SwFGvsaODWbwaO1kWSu99xhPhOL4t
v1lrNO8wljx3FQZg8r6McgSd+fjSq1meJ7k3Ei4oN88aw0D9EJG/RFscHUz0GeJu
m0sPidEwLZLLC+1zypTj7NuyLglQwOSxgr7z+yp+jxZRvxXobgpSYXrGujxo3WM9
rftLeqJDHVrNaR5zZzxkKiQT6ZthC2o+AREJB/9DRiqT8DWUKJpijtWnUxMe1SJ7
6wN/LZudI8FHWkVgLTVFRZzSBhiuA4tCwS6DaWBMMxgSn0D+LNegGj/QHVIwZF0Q
cGQBypY3VHExRTnSGc7UwQoXxwATMOx+2eAr/B4aCo9LQ7pvjv4INmff8y5A2kWx
EeMZPY0Rqs2MXHvHlPTyN9BRgH07zMGfmwkgBRwTHkXp3EDAc42818eqDcS+cDAM
tKWi7tddPLKwMXAxSn/RKUXW7i+QE0YlV1LjCKMI4Jz7cZPSi+DfyJ95IPm6d8PZ
fU3VatphqH124O0CCsfJqVIEM6EX1u41VZjYvsRTWjXLsYDlwVm+MiKKXYdJkxbk
qafm3uAxY/t/h01fr0tpINhyHwP7g16cS6L0NmR0+bZpOYFCbJFawa0tXXzboUfl
Ip/KIN/0Y+29t8kXDNkrgH4T3f8/vEAXeEu6c9fbkHHdM4Q4GSe9jNssiNRNUkMa
iwziSchLLdYSinxx9DHEeix8j01py0JBVMRRpaeFdizv0N++bENa3/4O5UzXvkPT
9OYlygnkEtsgBRxitmWSmCBtsvVAbyOgog6fmQJ3s2wuCjj5RKkdMrYABrdzjg6t
HyQDKf8rdRgm/twS2BxOeibj0EI0ru2WmVR057X8VgYpJATrv6pV6WBfHBfGB2Bq
W6xh/b6O8PtJj4rNyM5p2GQFTsrPR7x1rcaWLsbZVfufmasLD58SoSBeCm1sdWYp
F7RiZ340YWGEkusJWtv6MYqLbiU4/OSjNwxxPtGX5Xecrr8fijP9tWmrB2yiAVEb
89jgUY0gmGYJVL+HjNIrEU7P9Tpt0EunIblSIC0wwdSx/b+POSZrEk1u2IUddWbj
OcvyXs7py3tQ9pkEd/L7oFE58Q+OLCXLh6zNbfXUXvKMhuhPWj3rZ3nhkVFUeQ/6
UdtoFNzEATLIIASnA0w5DNawTfCV8weHEknu3BjsngfA7bRzXnG3wDr4CJ4LK7LY
TpOgvgGysETZoVTo9s7PU2fSPUw5ZACnmgsCTfT2KK/kzCfW4WZ7YLzpFtoE6x5Q
VbMhQELInPgjCSFMwV4nMswQ7Y1nT2m7/tJQiPdx3p9HXvQZqDNwH5yqo7+XGjw/
tv5yekBVnaFUMIIdD8+8u2XMALNaHVvq5v//AF7+wScc8tiLmYUthrgHvO4w8wc3
CP8ZbO4FeL+96ZCNBTpL69MUrj1oO20WyTEr6unaHPglJ2d+updGRPv+Or9Cnkpf
vpdD68+TnSxo4Sqf3mm5d0UHoKkRiq0YrO5jheE8rXCTY0TGuwMabf3Go3G6bPT5
rrMnfQ08ltqhUociloqJaB7Voa75pv5ILZiPh1/QkcQ3/ffQvjFxfk0w2R84lMgM
m/iain4XMxwnLLBnmY0qe8ZaZUmjSQHkqlR8e2anV0L5dApAo1QYfall+qeDK+F7
fntDYHvSq3hzwz5UiGUJmVtyu2vkhOXqTSHqb9pZ0msxfG/v0DXQP/k/8bzI19kx
Ehf7HJ13mS7m5F/y8kuEjxoC+U+hSU6kyp6A7e3Z2YkV2CJTdBw3XBmjn+o+gcP4
DXsvwxsN700tbgHX3lSd+RQYX4eDjDHWz03roDSn9Q9TQEU0ltDp8I1q1OkSimGq
ggjbyxhLDpl8lhSvDtHsOAwQ8HZ2DFYQ+Pyzbx098Ut7VhRJmib+BsbjRCVmOr79
HuOoVQ/n9yyTK3G4H+SEm/U0mT+tMbM1F4vJI3ugQO6Mx+m5rc8Lk3NkRY8k6mJy
4l7b3EETQ2NzTVh23aWNLeG3HW9imdCn0NIpOs/mK0rLghNTHkG1mTUcEpinxWlC
0C1Po405Y1Z9xxZCMauLrqIECBjO9+ExsqlO9fQuiz9aSED/wUdGU7NDWEKyfczD
0Aoi1FzLHZxit+3zTLI9VhtBR6WXhhO27Ac4a+oeFdrIIOqixu1NI6qMHSnTYwSD
scmyLIbJdHKJr55TOQJe3iZhwsbwEMHDAFmNtLYPvvArpbUqfdlixRrSsVSnEOzl
+U96B2cywS/TwMkFTfj+0DKgKXacvXoA+Re6Y60CKXtZ2l1u7css4XVq3lRIyBvF
aGARQYU3/9b4nj2JH2jmITGD/QZrOqq5g3SrF0j7mppFauuRNxNzwF+cN/GDNxvd
R6aqY18NI0T2xxi36AGJbKMQkDb41XFppkyexQ1xKMOqzqySahZD6GmaHp2u8JTR
bvnnUiKoLtLU+LwzrhoVH+RrMsGfkiLr9zyKVbxh5rhLE/eDr+3ZcUMOQU94WEgP
Hn6rPk6Q2Dd1nc59Inrf0XgMZqRzZoMQp0uZ78JX7htiBGTzTA24uuisLt3XhaM1
SBdzDERtX3O0bVLPQDv37kfpeNc1+QliEmUt8NcLoqT3YEfJaGYM5SRqPKzlGpFT
TAiL6t+gjUw95g9L9TjW0Szba2BZv5efU8vwtXuCMG454dtZvNqTCXspRPZyjohJ
be43nJPPCnMrGCc7tmd2zd55jYztqGs9RrCT7vyh+vLcL+YXehF9Hl3Pcrsn9TD1
D9dZmeY3uIG4blt19MG1reB3aHU0bAyFUSrq0hx+xYR2pRvzakxWQA1iYcIcXXjm
UD5c3cc9xlwNXvsRPZ3I9yvDdB0y/QfflcN1smLuj8geZN0lQTzPFXm7Lnyd8SmA
/hMBIvmEVT3zYpxrvDjBsAiXomVhXISaP2viq2oDzhK42+BjE/YMlz6oRG1GwRG9
RadE3evUBzGFO+jbqbC7JoCMCLosK/9Xp3o7g/UDnHrFvoN3xVovALdNcj7lZj0y
/cVSr/QXlbNR8gSBBRId2qjsVAC1hklmToaE/UobwrgoYP0o1AIjECNUK7piK9oQ
hN0HEdx6uptSd6A5LE8GR/THe7dnDFiFJB219FvhovJpOYgJ/rLuRpqixMsRGnwy
uh6QDvFCYvugPxoS/VMciVYg0W38QADe9MzzWS02rDsi2YOVPvfWJgiXUzR8i+D/
YKaDJqGkVtZtPNTNqfKE5BPRaGZaxbAfzDicFDVYOvrlQGqhLJ/BB1t9bLy4SuMf
Cjlhp76irqs1I0BOQHpVmXySpUnGY/38RoBojzv2etUqP9+PqDICefrAVCoEG9tK
ljlgpVrkqqxzyBXnASs4Lo0NDC3stytWT4/M4ZugxOe1YS2Pz24JN8+z6JpnEZE8
zlExUqiMrIylibcxBOhI3hbVsuQGGBEcimdNQO43zZwSfnxww0ELmRnoylEP1Ysf
W/iE0vSI/0SNYkRtawg8WrC837Pj1Z3wsxBWG4ES2rbHtADvLc+/4ClBLi1A9vua
K4yyoFGnPZzyb9Ip1reDufL76/V/eJR8IKzULOviSNbyxXKLHM0YHQkjwa32H16n
iPw6dn9QZs+AVM63f81cgGBUmIOoM1qnJ4y09lB4tnqRItaMxnXlfueNAJcs3U6P
i0HD5+Q1kRt07/76v2t29saBajiGlKPqJY3xWtA0xMUbK3IyP/xt/6cFXg+TzZAw
phUlKXhWQ2pVrxRMzrWdftSGcxtRpR6UowDauLWxGQkQGrh3qXiDNpbjn2cLY6mj
anoyfv5J1BNuCcKDt1GfEHljXMmZXMZR4CRQwyBBRQQO0gk9b5jWSbfc9MpseO4u
n6/gxYkf8zGw3o/VeBhjWb/gqnPBTkXpDcGFVhJzpCbA3vR6pxNP4Q03Zbj3Ds/C
OOYxgnKovTFFFuKMqPst28f3qt7kk2QgEwU8L5hWZnxldtcA6kOnAlg2skxSXdfO
GbXHG0Nz5Klx5GffSMiiJ1SalKbDqYRrlO+JthicdFS82z0YzPRgi9QGOH9JbdMC
QmfzoiEbEiQ0IbmPDOAewK1je73hXSrdxMRUOSGz2bsrso3fc4QVov2h3NgD5PiR
Ii98CuvtMsEpTIvHoobIVxVYP3JZxMJTnZkdXMU3lIUPkMJJVfKwEH77ExUZGery
pb+vPIRvNNXffDBfuTq5ZzB05wPkMfz7ryk02JRilSkdbhP7awVSvdoSBrSdg6b9
ZrIQ0faqZp1d2kRVjuLIGnqOIhhMpqQZARmitboVr3aA3aKUDlxx8vnJBsSgIq+4
trDmG8itds+SZRRj8Km5kpCb5U4WZklbmvE1Qat/XS8Y6RHM4Bf3E9GaQoB3Cgbe
Ji/gztYJnmjbFCnpZs0CEaq4YnvgtH7dnm8IKzwounZJDbya1PT/I29YB1CUXeji
EKsXW2OULwR7J5QhhNNoWGEU2REj4D/OigBYk/5Wt3ZoUHeadjd4s+QGFwOfDcQw
QJj9MOLmAd5hiVjfKYRsQ4SjUx/wuYliRe9nIQ8nb4iNhcZiNKiqQb50Gtc2qcYD
2iodxU6X6/M339gdk1RPIbevFobclcGTiyRdYKbpXwSnHEr8qCCyQ0qQZwvPd51s
rDyAVbaGwRM2AJq4J2vrkkdWMJEm8WjAFyX4bSrv3cws6pfrRg7pOJj4pExltpeh
JQqCRaYPxObJweQlncYphjGE+e/xPeD/zvDMc/ylJS3NW5FK9yKN5qe/xPiq1xv4
thBe71cVbXOrHRVfMBxQBJx4cXXywVgjF/Ldjb/gyDp64KLh1QuVxoY8tvpuaWyH
+soj7z1j13ieyktU0TqzPWY3C4WXRPHxkGRkl9wnhB5/m+U1gMgiU4wOn4pFDIp1
x8TDOv1wv/zf68QPoWbeZbbJQuBmZNh4ax/xUWoPksrDTkZK2icFu3nfBw7IhnhX
01SPMK3ppRIsLnVTZ5IyIr7k58cp+DzvENXDG0NLvwveTUVoIrOoi9507LYiSB7K
qBrYiXKc6aYKm9/sLSudh1B9uCsTLItKxosPyeCKBnfhJQjVWz+FVID1tLqwiOXP
FrDEYH78n13m9D+yZYIIghgYk7o+gln+DXQaW0ip9nXScq+VrWl1trBJRYbl28vE
ujj0bdPQb4J8oDtGNKYmZTivg+mcgOntUUJP9AxHAZDbC6Su0vvijw6uciUeIXIC
DGPubs7tvh2IZbEu/9I3J0EJ0vm7YxcAZx4QyA76FksqP5eRuOV3s4/nUyUnXWGp
+EQn26ApXiXSZYPYeWPiScNRwGdTjriXQnpRnsiwfXLbzZztN0wX8F4IEvkZKvk0
sUTH2JsreJ0tpiUzvv5HskMd/OWczYlTm805Xg8YnRpEStLIvdf/eMV2+mZvg3jO
gqWgKP8GwdIETZuX5Vk20QQfle+PuDXpTR1Yz6aucL/89kV1ExMRNhXmrTU6W+bS
dKTGGQcthfVtNPDueFIhMI7ppPkTbelg6hgbvnajn0jUy0MjAf8FVB3OIbchxeyl
Asewzgq/3j4vfz9PgUX7CVKoPQUkxqobR/YXReTzcrPtAfYpsnIq72ws9wbl9/Bk
NK0+kSvRl/vMhNFsmama1G09+0Pz7J51T05ron8xziM3V6dhfo6sP2L46q62l2Fr
DAgo3bPbIC6pPQ0tZz/u+aZQhyw15kSbpOE5P2BInYb7SeZ4nqWMidIkYrzPdKHy
1F38Hnq+PbVMNcCei50q0GOOOsLYGDYl3mVDkDLaSbzUzlgEcURfSYYJCJLI1b5J
QpxQ7LcaWhrjPm/OeKZcK4sW1BUwYEgKxK58W3DPr6nAul2O+Hx/Me+ilpzsW2RT
21YmJi52oryuiqFFVp1qI/awn3hvGwlwzABwSYbMjDkgJglC9Tf8Q7L8+Aw7oaU3
nKMhfjwuBsu+zZef7oXJtuZVvYBERjlI/BoJ+Qn41ApQpqoTIGzwJP43gZeRA+0f
FrP9kF5B9IvQsWtpfzqJzgEQK3r4E9qexP+uo8qIrsbnK1raP2/z6BXlAukQ5aD9
0B4Q8q8pOomUoBu01VOnsm4R27/wSPdl6VFFl3TTV6JVFEeqRFrPn9RI2m0kzhOx
s3k16YEHkpkZgt42nAKbqB4vvz/FA/8DNOicSbnOlMTwG0QJ8u3Nr0Fd54D9jfTI
J92ZPRFJ6OvP4cNmn10uhYVJCx3roEV/md0bKRBZBHKXrL11RMoBH95FopBlRhtV
CWbYhTOiU/Al0J1pJi9RaUHS/7GbQTEn53fQ0hoo0rqA0sbnZlTK6bSgx1WSECI/
HMlIT3OwvUudRqrv7/64YvgUo/ltgM4vZSFqBAas2Fjub7+hwvHAzxEuMblLUEaQ
v0yMoLaKAGJ3YTwf7gC5HsuSj+4xYLbdycyKnpASMuShBvSAKD5Q6J1yhUKBLJRN
j7o7qsQCG3FhvPNQXQVNttcwEZG8yR36jy1kyRAp/nT5H8xDUIdBs82gxsZIbdTn
mEQ4GAi552MP/y9qcd4XEy6hlro46ydLhopdcIta37t4ezjaFF5v/vtH0yYuMcUe
QJjzkTCuX0Fyw49q6r1nirtMPW/41LBmlkqxHllLpBLQO4PCBz9MM20V/JauyNd/
SSCQ0Y2TDZHLg+8ieN1M1j7LkkN89m4YSfedc7iQud2n/67NeXIAnY5Hx3dU3mJT
CI7j/sHjegWRLVMVGJHHSLIRL2e9yZOe51AVBaan39UGIXjTSKnpa/q4hzWvKvmh
dZnRdTAdwMsRnKE0w5YmINKHUFPnn8XaJWFwO00eoJhgxI2Z9Q6mDiTAZO2WBFCI
DbBPulO7dkgof9D1cF3YP94D609LVvYzsYWbZea74X8Lq+dCD23xwFhkeGreoDzg
MHOx8mfHFHRZ4J+b41DzSIRik2UOiKZO38CzLODXToR1SbS2qtvolfDMspkWlQRK
WM8A9g+PUC3dcJR+qwei/VrUs8hc5/wyar9hwVN6rw7UKYsf9czbsNUcQaYq1O0z
aW4npFrRBDPUk0F4ngUsAHsE7ROxjysrMyVcTdVf7O8MP8XUwbE0M/0IKxSknium
nKA+v+UNzAClTeYVUNibrrHdq9MYl9wt3OJr8B7j2GplFxZg6B2CI5R55MbYP+g7
yfTRZSIiDKrePv8tna2wQQI7uUEaaDsgtCpMXi9deshqh+RLpPm5PWCPI+4PSHSh
2t9Dy/NKEqdj5e0sF0D5IP+2hbPwpPyMMwFuk5rJkqmLHZQMfsDF8nU9AQktdKfQ
6CtHse7IGYwUHJziPDQP86zHFj6OCUpHkm19pKnX3EHzA8Ex2F0Mzd6wzaIL60j3
TPPQ2RR6KhEKoOxJJJx+10REvYSfqXCQi2Z6FNEW5Fcmwnsk3OAfSIF/Uer9D6yi
JOYMVvFDRpGqni2tFz98bZx/1dV82NKUv0AKChqyp+wUz3VpGe4VixJuHKRSEwr8
P9yk2VrfYRtdYCDvod0hRjvBbJaieIoc1Nz3nNt3qIi1KpTDI2VzT+JDNtPh6xq/
YtFb/Z3drRsyrXhGuXWqk51BaHe3qZHUWruqKkae85Jfg9GFPYIVtg4+uznSJ9IO
UHZbYgonqI4PrSNO++e6LAz6bvywnpZpB8hw+3P9Vg0eZA7fprQp1oNu0N+yxxbs
S5Dyjl0ExmrQyx3UQ6Jrvdq4Sahj5LCa6oaT/xMqh4dtCVsALsVwU+QSVq+Dm6zb
SDJezwJMKWlyY90p0wffXI/tg0BAf5S6h9Xu4xzNd6sMmsacWPzAHQZqXhSn2nVZ
+BrbuYV/75o1I3uma9rk9bik6/n/QmJFo2BnaQXJmO7xZUaZQzi8qO1EiRELYavg
z1QifWj48MpeIA2JaHRo2oCFIKG1k0cdkoh3YaoIQplleO/dDUOAV0nErdm2X7sX
09OBF8oEpZQAii803lEC2N2bks4Ck9tUtrZBFkGJRUEHHTCLh019jSVvS0anrDU2
fhhm9xLzh1yMbFK0mj8r4K1MLjO8A4yw2uPWhXSjaZb9mnTISfbSIEsWQD1bM2Ox
QV9EYVdDKT3wkPuOQAdfZ6Pf2zYkYjfTorWpkgz9BIWo0tZp9tS1Sn4cZrxv46rI
deiFrQ2oSKGMSO1NqXzQtvXQJbe5SJwZLii5rErFdl+jItTXF4ZVi3Tlkm7jVA1/
q+6N3PH7be2sVE1bOa2BtKz3smxSgonebYpNgCE5v3q+qj774Hcm7kA1NXwZ2b/d
zvgmFDb110VQRGanFU56/CNWyQXAcv3iVRIwaw20ngwhFP0iQ9Rk8kdMxcWJ3bYk
Nxuf7lqHDj+KU7mF/nJwuuERXGmEw+fb8MBNIYQnNCjLkAj2DJNBGepRxuY1/6O7
Z6e9rVPc3+wX7Zxfwh6USXsNQkxxAB27qZmMxGYENX8bRP/r+mkxM52jEALZnRu0
a8UE/otMrQ+6EWBvWEqO6FcxRLpnG6jkbG4nuDZWraInNTCXsg3YovPVZ50AsPHL
VkyTDzM5cikY/XdJ/qRkPcI8rnJLOR8tfawgufM78CAK6H9CGfDHWQv8tCjJUdhr
OnlMPBtfkHFKkrDx2uoDlcQPh6FDiY6ua4ZrKVFZCi2A+Lao+XKTc5+LxFWe2wje
0P6Ts3xU8xtgqXXeRViuvZIzwLn/xmiCllV0rb0sI535SlDJj+yACX3QjFh8me33
DVYLT+Auef2m7JegA2v4swPllSxteH7YhIZfwnU+HMWNXTHzkYN1ETq0UlUtFc/5
MnJ2tv0jXfJ6TmX5eIw6zKMkn+zwRo6IB3wWP+fU7D/YAL/yR2JDZ41LFrhD+nsD
ueMTO+rmoI2mD2x7wKPTIjBNzze9MM37E7dGdT7jtzr3vGeO/0VsMWc3wn7NBiRr
5ax+wQJ3wAvl1iVyZDYtU+9QNpvjLmd4AfaPTpIRD7rn3VKJLpEJEdqrDE0JITiZ
7YyxBiXmuNfX1NZoLkZY8kKdU75zdYYGqJ6/ljCuyzdxTjdwZw4Z9OlB9s4aZPHf
O0bdS/LM1quaAo3LLNLVXs/xoXCiMun+XEAm7N2PaDz8dBIiPTEtQzjDPGqUOZKO
dGmjOaDWXuJmnOyhEM+HU2bOiHb+mb+11rIULFou/gdzLnB+p/zU3s6rmXuHyx86
NXyNoijXVKxp6YTVHCY+WQsvzsfUov/JvnUsXBXPK5pR5SykkYugo7hHnkmN4EL1
/bQErE1ua+PNSJV1ZaR6dWN8xhwuSip3hSSaL27pgj98VDTfNqE36Fjm2meZsYls
4Js+2VywkW89U5Ox74Z0HGN8tlI/9SVs52uexAb1leamniZfdOSDEhP/zphdJrSI
vMQMXhqrKIDMkPzc0TROMFAB0RkTCv3qXIVNu7dansXtaumoEqM8MSR3bBjysKAf
dYapZxyBwtquO3rEBK7H4DpOciMiE9zgyqQUwpB1SyvnpbqAe/FoahlZPDhnaRQh
f+abbwN4w3CSgt84604KhyjoqIfSPOIUWI7f3Y+/Hw78AxyiOOKR5/ZWD7QZuKhv
fm8M0xolnqD19q9iSEP67FXvUjTMWOD3eFDxzS6Y5wh+hUCL0GeXBGJynOwdp7Ft
w5fv6MpT4KoYLXDJhYlwQvUFlzfGuBV5o26gbT1L2LZCQw3Qyl1gd5IGOCz253Ok
fbzocC3BOp6TvbBp+pzAK3VoNVetSxAPVeKS62TDTJ/U1jE7PFN8TQYqC6C7pzI3
28ZwFoJcabWdidY1h3ypV1HwPgRNBdIHLcoXHHQpd7l3almspyoaZkoNSmt/VgdJ
iA6ZzoyHcoR6obKZYhHyO7Nnxwp9vjO80xWgvf1+aOe05/peb66O1ilXnc1fBA4F
zV7BPWANlbu0G/hVITrxEdPnwypweXZaCVooAhNfeMDd+JB1ClpbAdi1xFWsXW7e
Edga/FNeqYU6T+eIOEc7cnWpmzm9GNfl7fd1FfVaZoCFkDhGbul4jdGDwhLfy6Lb
Nw55JjsUihCDbiMpDPKaNjqrvPXLFa20TPNIDxS1yV7eyROhZRGeQ2DmgOOPjK+k
BgAu5Pa/2s4u3iK839v3I7cPCqw6uxrOSJq7qe08o7XBBdgdR95WggieEmOUYSK2
TJbAtCXpHdbdErhDP4RvjR35Cfmgx1KNJaW4k49PwAZ+1MFRFhNgwqfAqzicj8UL
fLKPm0POxelAMcKs7ZIlUYYTx0PaaMCPp+RGJjXhPnk98wcpN3FV1Y2CvF3K9DRu
FfN8h/k5XIyopZMfqFvs5ZgOS92yLXU6co4gZdXnCfhbK3VNSF88wYlyQtJKot9R
+qvwwg/5xZWHd/yvkXp+Ew+zQsrZi9P/uie17bBEFj9MyyFlvb00N61rwAepOgQB
w2M27YTS7a19cnb7b4L36pH4fiyVBp9AwLyRf085oR2TI8MAhBxjcrTcW34LRvZa
/6o9sfJx1eqsjsrvdnquTddyxSsRLqaYGQQ0+lpEqSgHruhabguVb68QgiOlKDAQ
/raeiaHWiDRymf0SzVJW2xNwstuE/sGMoQ5GrndJGsa5GyoMwK/Rm6KanocDxIzM
wkwRAJLwXKNImRYIbaraS+4DPD7Gq6FMusgQ8Mc6b6ug3mXfewNigs7/efj/s3MR
KU+FNd/n/qDTeMGoK58Xe3ZtqfBneGhHLZndeDOiCf8WkCo/vNn+h3JUH71SftNu
OUd6ALkM3Ji1WTNTYIAfKUSW9DTqrJX5sgyPbLkn0/BTFgbyzw6bQtwJSfHwf5Xh
D2JPIBCoLMqULwmT5VBWDmGVxNP52Z0/+z6q2Q/DYTkXP4vvAeSQQAtiJc6QxVPN
GWC+hu9zZBMUO7UsxrsXqnM7T+L47yM7pHNe2LwiwezzeUS8mj0SSphArOga0egr
eSy32TvA/+pOdV0yfX5H+fJKKFCsMBWE6auw/414yi0CW8FDNirKxnhxOVVq9ouR
jXSiz2fD9rZlYoqOCOh/5hPvKiTqkWaqafesaSzUCTf0CcxUQZZTbSQWxsKJZcaa
iXZZy5Sqr5BcPmIKfmMhpJYV5kP32ozU6JHLEHACwKtlPRTgVKcwXr1gdRncSSf2
dlro7UbRRch9aa7hqoQPICodIIImyKQVfo0/U+7d+u+oHyRapY1RoKwqbmhKzNOS
UQiUnJl+9xdt0oAABMrXnmpEbfgJwjAfi9vyopbCOHX7lHaY3l7LtILJhR2wpd8x
pUhlgdmltX4m4HYfuvTpgqpemUaPkkbtfZOKPSARjLjpymsPhL5zDjrKe67iPCYB
AgElqezvEmtWy1oQ7fj4nUWG6P8M9mqOjO4XX0VrP5LctHe/CYYDLTYoei0pGHog
7WnpclfZfQzNo+wHabFK6BLyiazxGreTywpgyUDMQVV/65cCGu0Tt/RuzF1AXJpd
QwtRLMvAtfBkmlsUkAiKJpneAX1hMqiSlOxLdKYpovUBfniPZRq9jGLMDSSf59Is
/6802WMduTidTi2nMw5NjYsjgi5ttvGRSPQDZyPpcpOwCI+oDJA1vP8F1Qsk30yP
9lkxhDVeG2KTMiPdI6tn+puslfp59ksRCMwYXCLFf004q2CbYHCVz/KdRdxkuV6J
p5EBiO8/a9f0zkr7xRmpiru8mDy30YeQ4RNDlMjEULzAFN4doEVmGQk+RDGr2cUM
ZulAfIHDyiF6Qyaa3rXSDXM7abk3vcRZdp3qwg4usjGGW82qI1sKo7coEXce8EPb
q0WLxnwgCd9xjyZ+O9a+zDJyuJB82mQCx/clMvimNf8eJJs+O22Na3gSFs6y3YuW
JhMkjS+/LTEuifH6c79jRsX5IR1O254hKvkO5QOiDV8GEA4JW5NjVo6R8hJwY0iC
GxyhRvXxcfe26DmTdhj9wZW6CltQ9QGnX7Yz6HLa2upIxcC1VgP40BHbY1Unsn0w
18sIQJ1rcU7EhO489s1Rvi2BZKEUh0eCkUxXvieNGGWL8IWXdO5yyuPt98A/75tM
Mv/FaurumWYquBzWFqpu2E/AC3KkHNo40mw7EZ21HfHRXbojwoHgx1zjgfxqJ2Nx
8V1OwP4zBV0CbccKXQvgY/VWEkHHSHCd255MSES80ZhRzQQsuYs9fnj89DbdnzBn
nBmZIH9C1hfGGs9aX9N6dW3aYk3j+pVgqkkEoVgU6R90HgbwfXdZ8GiF6F6HMPzg
6pEoX/VkHauKaRH9XOtaIfXydSXzKHnoa5Z3BQhYlOMW88w0Ou6EiEe4ZSXVeYuw
kI9RMDSiAvsBfNPn8MFoIacyzuSpP7e0ZTVU8uXDc91ZryshnAmPFVEpLWAuf/gx
BFyZTlXQ4UJ5QMlaGAdWQqFadfXlp1TU2680bByrQ+bLmlR8UBHTQyv+G7fBan9e
r55mN/51HPqzvkGc5cQ5G2XTHJY61FwAXJ5+VFr5IM7IfbBeiCWOBLgP4hjgfr1V
8VzoXChRfsw9G6fykGWIaoHiR6dojyTQyzw8/TZygZiGItswIqGFQh/R7XiRDdiW
qrRh5qtPqP6zy4nsa2jSuB3WirVACgDCCKW+V0Hwa4bxuX766YtvZ4cI/fXZY9OI
6HgpHu85dsKUSgrowWpgjpk3HmC/abODEbm9KHLA38nZOnPXQJynukdhJ5CAw7GK
h7Qf27QI9ogoi2e7aYivjZDNTAnFSvgZOtaVOPw6tWTVkSbC2CZ30iaHd/FV44El
GwS2T6/Ep/hJPf4VviTcyZngmtfnw/4UK+hgcGkFZjj5c66tfXb0GOpAXpaaOLkR
ge7BOb6unK7uyoSg7zFNjJzhiOmbRQcdQw3Z5UHWFDKqpAT/ZLhcKorfkGlIjKa3
24lGSxg71stl3/IwSU8iPrQLc+NK4WRyZeWzK5ALo3XpwwyrFWwr09e9ZC468gL1
bRNiEOat0Eu0fjWnVmsWG7jxiflVUZFxd0PdqiRxjbLNpp/KeoPh2IS1w/3104mK
qSm3xxaXAlWLXCcnzL9ZEBV7VduoV3euGTaLGth18ziiI//cmPhRBDe9A5J2iJ+g
fVJoRD0n/JPN5aMH9f0+ikA0U2xHCZKfgahNverWYOsQp0W6XYCNqwRLl8+8vp4x
mzjQUg4WvTeVoaJFE7q4r+OG33yzllyKVNB9af3QOoAICTOf14B7iqCyi106XQ3O
XmGihintp9QR5lgli2iqB4g906sAzRFK/v+nlcvd7Nd69GNaN8KKD6srjG3Saf1X
0XsX8zWxFOm5SujCrEvMcG0aOw2QtBzugXDdRZH6LRJY/VKK8m5VJ34SW4ZUSJuT
EPYFi5radjoazCG2t4yKUr5vxwA64nhgt1nAhGMJxiKhowZmt3zI03x6DOMSGVdJ
vcvPP2RvRtSOI4HnSuHD51C1wgaJKtRBWV8qbl0yZxpW8PQ5QJrf5kRGlFIMIp3g
xT98mXx1G3hCw4cMO3RxLBo+saWkoZn/MCA0Wp2KLABavV778JpmE8ccgvzyH1s2
xcfiw37aYQ4H2tKJRtkL3k5I5HhGoMclQZFUHpP28QvVonqUEr4dfo0EFT/Gk/e4
psy5xS531dWVuzHfCKCmHp975bBFy33KvMzVkf9HTFoKqtTdRHjMaxStxr1Uk8bY
YX0EN1DQXPxmkuiN5Zpq04Fs/khX6bvVuMUk+W2Qo/Eo3WHkM2Vc7KPwHCxbdyer
efpYSKK1jpbOHjbr6XMP722oENYHZeVkA5nRC8QEhNthvNeh0d2bI5BjIuatmwYY
UVw2jeM1aeikGTZw42upzyRpJjPL6FvIGDf50iHffzBDB8obEFuqCkBxNfDz606I
+bwUXOjE+cBJ9GDjnHUviB+KCOXm+AFDODRnJGbesGSFzjcXgXccqZsxwVStwFXB
7U7+HtgiqpO0mEvoTs6D2nlPUUnYXRKAr2kOJ3c/ZdPMAjBc1kWOzJqlv0sNb4sn
EQy9kaijkGH5OzskhOpiI2WJpQxvEaca2rkFPiCZYC7l9Q3RqLa5+PaThdaGXbfh
5qC1ZFBLpMglADmbPzQ4N8rK+D5HSCWMfUcjL3IDttPJRxagkkb5/BEVDKJ1fP7s
BRSi+FpatpY3rhHqupD4K4baswcU1w7vIxh3T7VMFtqpQAUOHpHVXzKCh3dVBnKW
GyN+qTWBkJY6tk3YvVvxMk1HVRHBhns25BHk3XwP8h7ETt+19veq+/5PvJ0GBA62
FX3UrewmLS6p3PWVD+OWq4gqA1utJpdPdCfTwPcMwoQ4hCEuGfaN829CrM60gCy4
1CYWegtP7leMoZGe+fSNr9kr/OYte7zh14wdL33+6xbbDfA27OLOZDj+VjOsbSwk
El6817P87rqt22zexwavC8fSfCCGW1Sg/IMAlyp2KgjUty+glhN4UeZBTY54/NGf
m9grNB6ZMkyfEN9wMpft1/GRmxi61Lp/OnZ7o96dGF9qAXXL5gy0ICDMCkK3l30z
esi+Tg4tdQBMH2CW7OcvPc4ODp+ojdGlZlhJM/EwVGnjOa34WV1vE2k1VX6oNRS2
ZCQpu7jQoJDITI1ODD30hH6JEv7FnaRFbjk5q7SXIAvwxZU5HMljHAEM99ot83Yj
rWSh1coWf6LOfrdZ5NE3XqQbJjoc9wS78wfBx4lE3FPvUvp9K23kWjYl13o8Lk+g
N0wbz8XMh/WcY+AQIhqQyE2ZmzJi/rEaImtWDTeqii81TIMXECQ3kHTymI+1cvU5
sl68+1/CmSOvSovH4YRbv+RUwqH1349VBHbG2MKYkFYYruwDUrgPQwAZnDtiRbHS
vyk2BMMnR2O1cEGlEn3blsU5ryLnmRVOGwj1uv1JPjEEtwC1djGKNbz6YL5vbFm3
CEvsJ2Aoc8e8r8G6UkfOL58i8Eal8i4H/ENvKyj9cAjlUX/alFFhol40moyxdjV+
O/UvsKKTAFZwwSG+y+LOBGgo2PJTwMgKBqFBHomhN0wUcIIMONBM8ILSSRwMA0a7
cg+l8HAoq5CpZF+3DZWhJOqUUct2s+VCiqnuGqsSemJl09KM4UFRDPO81ZuySVeQ
/tT+ERrkKD7LyvGlyLXgAlXY+NPcUzxr4NX91ZroV/XIo+JS2vN9f8/Fk6IwA4Wl
I7O2x/WGLOvxM8EKAdyB5BNyZKlWTI94UEkBYUacXbVKKwzs67snzp9hCadr3hfy
r1nBIxbybgzQFn5q5sP6KBomqXT7Jer3nOgmRHsMHyHDwgKKbgrrqKJNIPIWeUOp
YtghQylgS4zrl6WkEuLHg4bjOzjCNByojL1Qix+ZD+J1D+w2vpvOtjoYW7OMraN1
6fBnAkr++YDOnfgPsMzAsT6T/2eHkfWdw/DNv39yHJle6uq6XGuKXzD9l4iGZJJ+
lyEU+7n2Dh0vw8Rf/CYqC5ifyss/Sdl8P4YuBsqxNAkqM2FdOtILyhxKFpunxxWZ
MHiLcTTzMEp4aoJ/wio0QFxN0lImpXVjHgPDRAAVR9c/k7wTjV6HxkDvocuzwpDR
p+p13rTA84IByxdQjqd/MeBhCXEgAoyJdKY1ijRISzIUxz8JGwjE/YXuU77H1Cir
6+GgKsr2eVIZmAJOdawDf0HH+TH16+Brrj4/s81Ep60oUz2H4ne3JK+M1GvM4vCn
Jtvzui7LJ2VvR2Vjw2PGFDNEYeaatt34VKZYLTWTox4YGDjWJ3J/tb3B6FFlgacR
rEauMdQYMcPF0nkBGgHnU1/qlXLNesjn0IgoyYTYdYgMbdJUhc3pbwW+p5UPCZBr
bZ5l+vD9N+d6QI8R8yWBMnqP9LV/QCPoCKEbRV9FEeI4TNXksRccK89Te1J0bE5k
T1cxcj8z0vixKOx3Pdf7NYWa8RxK114pfvqrWWTxPeM7Y3qIK14ykSt9nE8TXxBX
Z/oNMb4fXfeReiO1jvyQAgnPfyzQPppfAOg8Kyxxp7MrZepfS/8gpf839DCDBNpH
8kaANIcjOica3D9YewptuV172ePOG+attK3Y5dqc96UNIgVI8fcogUlLPEHD0LVq
dNLsEymSvRV8nE0aloDsveLd5YEl6b7YN/9JAAsE57mSFOkQBSDdyW6AZMJGYJeW
nPhYLz0Eme9IzT3m63ppwxtAx+ACQSVm72bA8oNcqz1FBEEcUk7ZkBhPLSTkj9ns
abXCANx7YhlMzCor+ewfW7arz3tzeCHScG89vt3t34SMLg+AG7tNEmihYRlwbzEK
5l7aEF7Yb35MDs5b17HD6YTcY7zrOILBf1UhwspLuFZ7T4YlByd/eLs6B5R5W2Nq
62k5OSc/Z0LCpDwyr5whQOOyRPm349RQnpjddMtgepK3EhoyJ8vq59hncsOZ+K8Q
iN/IELCOp5fm717EtshY3UmNhHk6LCDZq4zP7eCsql30Xookipm7+frY4v05Ef3Y
Jww2r2Fmfk+bOZvtqGkY/VPJMxCdsWHjhaAQbmyUzYYSARn+3T5i8fGL03sbLzHm
s1yRCAN47XMR9e/1TGJRzM9Z5GdvYO9/muRbI8gFmXGmAZhCw4kHQBotF/x6bQBR
xbFRiOeXKlpVK6YfaEr/v6ASap6VyDBOslxVMf94jTKG8lhErjMcY7VMCUhIe/8m
dhQnac4NMRnmsvV8vYmm8WSnmhWXInhJ9wLMozkYpkWjQ7123BtsFGX7BuOxi/pk
Xzcpl7/mGK2wcA0+mmdj0KLFAV7dN4gaIKempTIhZKE2yYa3P6LJJytwDi6hewvs
45in2KkJXEMLQySjehOt7EmK4dGbiMnDw/MtYWarqCwbkQCNLIrOI2KWZxEtoQUm
8G5Ncmedto+jealJAgmpz/Ur/KJ8xb5q6PXRrvkkth22NbFeiq1FAApyvBa8Nj61
a8PIbhXWS5ihSCnGHx+x9rRXzkViAoDZvztgXWFGlY0eCGZVopx4D43pw0xqiJK5
9wdCSctBcE20ytaNXd54Vvm+vwcwEO4+J4QG+Ohgg+68bYKnYqryecRWwhNwAFTy
EvFm3cYVbuWi82VVSC2sIJEQAuoUHfSqSWNi5FyasmmTKYrRrhWtPc2Ghme+duZB
dyYUlxKhhqKC6UsDlCxy2lvJfHKSvwcDA0+obuc2sN3RQvBiPocXeHGI7fuKwMvp
Cxmz7m15C6KBA3anSWriMTzI6b5I5t4EoRNmsiih8qibctqAajU6qeDpfE0uOLPg
DgRnuTkVRqW7O2/U6Za4jWsMQK4paO/e/N8Lr+C8NPHx872UISnR2tg8lRT/JzMz
9zvS9LPvGoTI2J9LuYrm9yyazVKsjV5dMIw2JxCoqRNv8btH8byeA2Eut5r8aqfa
GV5+nP6a31e1Co8wOKJOUgwRADYlmbc0huy2sonxgZYUfpkv52FBW+YNAnkHy/qf
sBjFu5rKqf3FdOHjf89ORe1ojUymw23HifvzvxaEXk6h5e2XfHOVbLHDxmpj2bEx
pyOt1AUk8VpQbHPWYfbrjiQQwAfIexWyakxJrR6gy0B7Nb4bO6P+92lHCZWx0UYJ
Ztow2LZmxlttwGkORwBJmATRLbGWMblZAvGmWSy1gdW14PD/XC7GXzpYLmGEPnuB
7bgoC6gyZsxiHW3irVAHLyhAyOqnM7KASTVGN1LjNL+nTAnxeAXvC0VpcDFpuHqZ
TYtPU9QzYBR60pR61uxFu1KYIzPNMyc43f7n+NaF+3oXTyVYrVf74YSpxJyLUY6z
y0cVzm3rbeUrXyI0gGAfWBoV8s1oDSNc2ifHhFvz7SS/eQvkk22pT7yGLCjY3Vg1
QbsVq+d/ieeHlpCGZX2hrrA+Q8/LkvR8Sw0ss8/nP68Mf60Z9C6GJCoHM3mNC5v7
pCm4OoSsqvbWO7Ntddpf74ONLM5736pSvFJE6EH81qDK8QRjSjigiIlnWYJIR7rV
GsOwlacQI+pmaZvcXkeUOhylnzu6jLfFO5BDLS0CICXqsPRG18qnwmcZ3+KsC/9+
Zc62WmPAH+7OhpJBgYQK+7IMpV0RxZJUtW8DoSxYrDp62IL0DJIeZqqw8vNqzYZU
RYNAl3VE5NXjZfmW28U6OVpWSHRmbQuMCR6e8pS4u5bwG9yySarghZGn2nsR+zjl
/V2T0BRCLSG8rjmiiyMjiwjWSqI86A2fOxA36i6H/N2mI2yqw7DEciBCq6o88btZ
Psgxf1j6RtAIFq4lX3recpEoICEolTxNGPXyE+0EPq+HT9uQtSR9RGP5lgWXJ/fM
SaV5ucgkqZhqrbD6erdzNfoeNibkLPPOraU7a7DMcREIr6HmzzaJOR04C3ermu8q
a75oMr734+sNcT+prtMmp+d4QUIG9+4i7ICnSaV1/GoiDKHvCUP5sZVmoQdPdiS0
BkOE9P3Lmx80eKpYzMnZ1R5y9c8f92mJfUE6CIJEOMSR2G816HKxCDsBr0l8jon5
X1oWVk+EqcfVVwBIZIQI2nD7n8JEdzJytA67Yd1Y4tJa0V4LXoZfYJALeCjjGuIj
3AhBsq1a8kB7OGTjTvoGRduQlmZXLcnCNtcuhT8gK8vvmofdH1rmF0ZqOpAinYPT
xOTvIopTLN7WghUMgoTTSp6kx1hWQpsHA7PtkWxbQ5gNiXyTp6sCva3MtozTywHY
R8+nLScqepzm2utlziQeul8IvUCB6E4/EmiNVFB9HYj6UvTETyYKpNr9ANmwTxT5
AFPzOE+tlE3jxZd1Gx9ovvH67lqya9zKiilPA/j7liHvlJlKsbC4cl5JTQEG3L7r
XZE301zoOPWarmJNHOcrgdJSqqYYVvBeW8j3uK3ghE3OEuoMr46wb6Bwt7l6k7kW
tZe2mFA8z8r+UtyoLvN5iFg2tcL+aEbXTjqmDECAeOgXRwDU/UNi0oDGBOsOTUjG
YLkYHGNsPrg/fmEnTCD8toT2P6X+KWU2iAQQhmLD6MVEIUSQdkslSqTiqDqBQyXD
yeslJes53Vu9PpR0jprDpNruuSvHjm/WeBrOgmcMwud5ZI3x0VTvY8FEXNXwVQ7Z
3TcprkbThZvVyDlw5jJfWt9q/ROVA1xVppbRl2X4AqnWu7fklEeI7vzM9L8vFxmw
bFwrIfvhnwvBOlNu8AOKWW0gPwKlZe5KFwU2M1BbwgMEO1ngChQwsNp+t4OG3j/8
oPyLm5xdzPvEmjvyFyjqE8hV3z1RuxO1Ix6XTyhwwWl/dqvmpMShCsHuiv3xcIAJ
9wZnIKsUH6YoGAMHkhmNYIjaHNLf/hgZKsqFBqltloG9kTVb1ZDGnt49BHewIgtt
mgeDEEpvGcWigmI2bEXKGNlbmpsy+v3Zdoeo2w3qJUZT1JKjOATfR6xPlacIFeg6
DkhNW+OGBZSQrJ2NLtPSjP9YDMpfiaeLuFX9XzVgi3iIdXNmyfDGR91rTZ9YDt1o
V3f+RTibHcoJVl3PFAqoE9tiuTGptwnJIUVNUsL/mC42K3E1hIg6Apx7opxpwRYV
9EcgGRY4ebtDTRdcjCyzYDNUI2Hn7gyzweiB/91PcHGx7DdkrUIDOm1GrzKQ879J
khs6T2yOMpgmG3BbiXIDiz6Snm9MXB7lorJ5sdVVR2hs3GF9/fMbqQs7QBBm3e9a
+2j65xK/67NwkPRRn+e5j5y7q1Lt01bda+A0NXP4+6poUM3PrikTkUBiem47SfDe
LKgDVuxJY3BBm8G5S+T8jppbVGs6McJc7wgafeq5xOqJ5Yuvub8SK4JLlJ/vmEIG
pAu3EsMUbg4duJYSqlP9KD0Dc02lMGIWRN5h3W9c8dpmjnnLAzmuLR5Kw2g7Ts55
nNzGJ7QQTDwJpFEld9unC5b3PPjB+4etr44H+NJfeTt21Esvrgd8rNMyiYUOwGeO
N/9zav9jJ33zG1ta+DJcQUb0JADC3zUGe0VxqtlcnnDermH8mOSmqbH3BnryUWxo
WxgKd2ngR7x43585yIfeSHdIfv29CkdwUg6CgFT/VAfFKla7fKSNGawZ1+9Qfr/W
esHvuvD6fZijcdIzPGTJodk4E4YaLhxqqyKdOokw5g1YL1MzGYcyi4daKQHrp7kg
6nd2/GO6NCw6aOr/1GhtvHuOYSn9dkRKioy8LcGUCMYnvba4iN3pVMKegOFcdL4H
g5T3gEah1MaQn8Sh4RziUR8KVbFmwZLoh8RgHGcZm9aisqePCqmwVxSBjhDOGK6c
k9KBmkOZ3WZsMAqxy96egJMfkAKPxiPpiqkDTsLRDEoUDtgF6a6XZBDvJLNimkci
mqGO8jdhW0LyZla7bpTh+Dwh2aFYm4EPUkrJ5HNCU35+DFHmzM2jHy5R+JpFGYQK
Vs8aummrm5vRUXfkHk30PhWuB3OYg6wosZtLNE8kK2QHf7jHwgcEKn7bYEv7eiFN
aa34wc3NWpRKc0iP/MM/WJJgPaVHMpQoyMJEr1Wn9MLxX06m2MJ0d8rkYr0m5oy6
JgkQJ1fHAPKkEgZeF++8rgss3LK2SwwvQ/ZbF+RayeHkxmvD2EYulekENy+8mgeO
4fx3EfKgjdZxg5XNjUWFacygIKi2wZiw44VRNQ6g3GlzDQHeOrD9kzC+SjTC0tsR
h2zPqHhAB4wC77oHdo7L+RME7aisq/NSb0vz+QbPvY9tDs6Ia23ci8QmdWZ0FAW8
LhjdPEr9dkO54Ej7mTBR5GvehaJcHUDXEE2hCuyunrVgVf5G8caD9JP1IkamyRWu
blBOL4tE9oHki02FIZgLRezku91l3CnNZrw/Mq+qkw0aZov18j4eJ4TI7vBIRXPx
cVrd9ciEvGAHQweCuE23pJEgfGuHCeAzIK65QT4MvWCW8lcTA2z6E3Aq2EARLoOq
SLKCmp9ssunabnsh0X78i+E5WRWvWqCsHlLjaUt1RyAVRz5gpg0nbNzVwFP4rpcf
Xp5MN74q1Fa8Ix7EjOelDLImschiuVP2hHErUNzDvTNBkYj8n/yO9WI5qfgxtGtG
IZGDRMtTYeYqMxLYW9B7Diy2jjlqxcZgtUdPlf5KTFtxiVzkZn8F2MN85s9Gnu3I
5MoXNc/gqof+142SEyHpLj/LqDkeoXMB3NXuQQZ0FbY6hq9F/9+wTT8qVousQvYA
JVwhhHL5RwKq3NTgcqS2og6itxFKKZZW2iiO+YP1TcZmPbKctF/3gwW+7bKGry9Z
vCFp0Nd+WzgusjE+MXkeE0o0mOmbUyIHUzTw/JjDjMBl5Xr9k2uSYdn/dIq/CGLH
dHd9FpMFy6p2HqXwhznCCj0A/aDS5lqfKob4AEeGdzVt8O57sZ5yWwbOYVbrCbQA
4wJY6el8dghZwMVMZODKOYLn/gKZAKaImSuA02aePIhBBIc/dHSHmOlU5BWO1HKt
DLw8GAUk1mIKvlIAmq1gQKIvKfpct9j8gnciNwl49cov1wJd5XE62NoJ8fbdDTe9
eMfw1GbLq1L0uSK4Ipnrnv2oxTixP/VO/ta9MpdMRVBTfzopSH16IRHUbFgDeVuy
1JNwkRZm9+my7H4sdASkaJUydB6C+Yctr6SHjnDxTWI37Sv6BxucrXDDtMUCCEya
Wtm2Qh2CePSFJmge5Q1CSvMayB4Xi3SYPEVK/yKyZYnTof+Jf7L9gAECzOMfFpCq
yLV9dGGdoslnbJ2OO1bHb26rRF4D/Qxv9gK0tp0JGtxFJwboIhlz2qaaDVwaRlQg
7/w/X3tuKSlkF11aKhL/edWa7y2ym7FCIk+oMjN6tur4N0LEhlVm2OmsNM65W3ds
kYkgfrCmlHs9QcukUrSFCFEtC6FdXkIkRdPaU7iFstWC4HHOBG/4YwkYwqRE2kcN
cTFykZi/FHJ67mEIMl1b6hGVR60sIAvqxPMl7qIfCB39ajD1V79W908K5BjpgqWJ
EMVHoGKNHDFHd6wCH0Qh2VkfoVUvcqrQ78Jgb37GSTTTQaIRowIkOrcQLyeGf1RR
1JRLz0+6qs3S0RCtiiRZkvXVPyib5S7Xpc82QGFrtbiAbZs7gsiE4lfF5cAORQ6l
731NDc74SV/UInBXmxuBvojXl5EMlJ6dC/rw2l5uKdLyVx3gw8GkEhcx/WxnBcG3
rkV6ibl4BODox5bqzIGhXc6omgd/JpLAN8EqjxLIFJJKhhje+btd+dFa6hFGos5i
JUn1gDwWMCf7xgxW6MvynGyPYF2eqprqVmVcqXxQ2/Z1YT8SYVzEYPL5bfQYduzo
oS5Rl0qBcECtpMEEfgrKqw0jcuvWSCEpsJmCJ3Nv7XNhLu7bIPK3gqeIlRBWNKCT
qfjwAhhy+8bpk0YOlelSV8SRJTxsEh63oGj988V+RQ1O2ZXuO4LskaRE1wkVeTEf
uOaI69qotwMItd2vL5PuqtBxikEvpDXLRr10KyhBzKai3yDhnUes0HBvh+S2hdly
e1XoNZyJVKAVZop4TOUP4LrHnJ73FToM7pWlRC2Ex1MjF6D0CfGSvId7ieEm8j/r
u5cYHGQl6w9dfL2s8ZpGBQx7DrL3KS9FEi+1BQ+aL0o1YY9GI2ZEGFVRTr0ncT/u
DtwhAGqRQV+EobddlGoehudLtAeJWZITv2pT2lwNhSG8fFK0uPDRds2INS7SjtZw
2acBcPH603Jz9s1OB9otKSiu/iWSouD8XM6mjofmpQ2kd0JAbTes9k+rYg46Cylt
vK2YN8aD+iBRL83kghXXtw263Au6Mcmj5VhCDylJjdctlNujGnfbdKeUmfr0Vb6S
sCAxIMH+zPSn004CqiwwEu+6OjaibG9DYgN+ByGSTWtO7HogY8csGssmNBEaHTnB
xYsOClZwou9vyXqgdSGzWqUYJT/B07NmknG6aoAmeYLjrGAKE8DnFtGkyoGP+i5F
CA8tJqGS0lyPdB3YwagBS+Nav2yathXTYNGAbfRYYEupI36JQHz6aMrXwdkco1RJ
H7CSEFykL7UMtPsEOHZbkojiGBaGNF8QXlOxFjYVlv6c4SlUCR+/XFmq/O4Radbq
8T9KLiujPf/GAREglOp2xSyjJd/7jhnet59335MuioI7QUh4xy+0V+qdZCFYmEYS
5OhqvJikKvLUhC62e1AnliX2AkBABjI8SDXhhSiT6PKe3kN0SQ2f77Q3ThGxka9V
WAmpU4eOyurNU6wvM4NgSde4U1NvKMLQcM3lVS63fGu6XHZXKIx4C22R94o0xAbY
AESrUVluo553Ayc4YGspndU7f0jVE2TFvOPwK0QEo74GrlUDyvqDORvNQOS5OKj0
/Iy2EQXEW0cPfHlQJUXyNvhGiyijKcoOypmmGn8K6JQNUdKR/4OCtqG32ioc4S2Q
gxySuO3C7dNfUBCIV3U39zqw1lOXQrOmrrf4mudLuOzFSxefxGpFTFyaujRcmGqP
KDDYQ9kjHSf2GQmWWxvQAcKC1VywCaEN6g9elIfcwQXvvT8k+eAqGGG328H4vmOA
AzTdwtlxNqiZ7PzP5avUZOH4ukYmo7HYbHD5sKceNcqUylJ3uHSgusT1I3tWDjBU
AsICKTHmDLwSLSRQ3PLI4ZGCxZd8L0xuD8N0aT0OPKgvUIn2MiqfqaHZ8SJfoHeJ
uhtSq/Vxbfkg9YLX5S+8gCViZfdlW8wzxsEZLmPhSqIuma9ffkotmrAOGeCLAbwV
LNk6lCUvuni2fMMocJA6QV2RW5cRAJYDysS1soObEtcj7KRiCtiiikd1BMOcN9QO
qxOAzrwghnXBkErSY1DV+FDm+h/KEwjBWCxoPHlam30WYuHt4SS3hiuY8zG5rLyz
qCMhv9bAbBcDC5abxJA9tWjZ1aIgIBYaPp+ADFlauWOE9zQqYrQmsaf3vb+H+rzS
XUDSY6LH4Ku9Xrrx2JwkQGeWZ8cE0O3FTFFDaVGlA3rSkBtL+Hh/Ld2ppQX5iV/7
B5fpKEMBqZu38BtNf6AWohjthPgVTBNNPJPb/CpfqktlQNuoVuPt83DpR/kTI+Zj
oIm/dfz3EUWevtUQS7kzVJVnYsWwAzdSVmmtdpFp/JQOKMrmEBrdId52gYvEcUvV
YN79BRmCNeE1/RYPQpKpVQbJh/xEdg8eyTirV7l8BoLwzATsbJuVpOIYgIxembg4
1sNIjFFl5acIRakGcw7XaMvFuYGZXDvQt4mBBwElQW3hiHLodlYjfpoImbKs9uCX
ojQPetzeOdIJ4LW6ltDI59RbXIl255pNkit86KsQUSVW2g7Pspb3KIovrFS5QIOJ
cUwCIkXgaEr++RXY/VWo80d3cHKsnOdNqEemUlH/9pYTxyRLU37sU6r/fmAGxxGd
fJowsKiJuYVnsbBpWuNYc5KefoP2BvjSrf5sq4g/RYZfLKV9XH32/hYHuPDfgiZ/
3iA04v1tCeNs/+h4i4uOht08L1t9Zd6AnsolVCyqGWZ5cEK5D6MrM9ShCy03ygBI
9wWCalW15O97OUAOQcrPWoEF5gqKFIFisW4rCwulHp0ShvWTZMG1gQRtlmwoNmu4
ogw16qQ2GmkI46BEIav1cxVm93GXB6vtZrf6Ul7G0tuLL4cgZshMUQ5CD0uCWiID
LDTLU18Fb5vHss/N4W2KBSS9mZoS+mFgJ5fC2oXh3Dxqkujy4OrP0mYkqZk06TUN
wqoEDbNz8GIsk1/A8xGKtKR+zAuOhGX3MBp5FFGxMRzdYYD/f5mzJYBaCdapJR3g
wmDY6H7vYuiQ4dTQWXEL7ui3LdDh6PhCiz+NR9Af4xxKEiW/MT6gjuhHnk+41mSg
vYhe9RDi9Q5Mk67dAaIalej7y7hDKPyj0enujtSrsKobckq6qj/uOoc73+2ymzDc
WItRTp6vwl3MyCW55ZIQdbdE9+KDd4WjVhHyJZeJ/xqTxTiY58ZldY9Luex0gKoX
k/c6+mqVzarYNUO4JhWexX5Y7NBFaZvgUGnCFlHjUxk98iuRe4LStzHh5N1kH1c4
GbvHS12TAVFqtA9njH4TJwXcXsTWbQ674DCom+ut1dtHkRkrRioHTJ9kVf15Gdql
u9Xp/XmVZ0r92t1No9uJ+XkDNdLVMgqfn/l2W3bNFqNr/LgUb90AeAMemSyoZUsY
TQNdt876Ch2wIt6Nrjgl8lm2OwF09JRcNcqXearPnY5lEdOy3Scgfxb4s0VPAM7z
y/KtYRbth073pmsV7KUcM7V6W3nmOoEF3EII8lG+P81TbX4W3TuhnFlwNkfDSHuw
ehQbC3mGvlUN4UzI2VOscn+GoWaLUerjl8f6Oso4CQpuVN853yTeUD2y8jRdB6Mb
mC6FC+HZdjFBqSapXLkx097s956fgqsBBoVqX5AvPGfmfyVPdlXv584BBeM/Gphw
fgCXQDq56PBW/pw2M3/cv74/pasr5aaCeiJDBg2iJhDbkuB86XPh0+j1elYsRVK8
I76r8WBj9TIaOYVRwwjDth77FxWqVKRTqqp0J7r2dbpUBQGBBuTUq/FA/LLOIo20
opiyrVyzQTq2kzIG+9bCvcbMWg/ZH5gaMw/MVqHGsTEw1r1Gu50VnxycLIBoG8My
mlLokIEvgcQhoIXrJoprdiiJqydB6qJ/UUZ/sAJlW5QE5OPCkDcUP8/FNtSs9mmP
TcmrN8VMKSh3CVqokAHkjmK9Kw6mevfskGVl09qTt2D0e8IbFmBwIEPWl5JUwCMD
bGMpION7xW8YZSyh0m1sqQ3AykdtCtItZgXYG8ruoZpFkCdzEWLUA7YqBVSBt06r
cr/IWzcDEGFgT2rz2ukxMp2FehmWIpEgZrahekkn3uQqSTiPVmPPzo+0Jb1gXqmr
bgKV1UmTdckWP8XZ8EUGh1JTjmbdOqZsDSVmWiR8MW5UZD/6el8OPy+2eLQh1pom
mERvFpvRftzi4aeE6x8U4fF2gCUpYEr4wGj8r2snJCMlCt/9+mJmxxZEWbEamjL/
daYkhiiA8qHdYs0QWNMI+kTUKCQI31lX3TWI/+sR/wuqsLFsgP8FeVNXTqK0Pi4m
Uz+tQpj7KNgxOceLid3XaCDaPWw6i89mIBSfls46R3vXHv4q410dwdX9MK+k52Qf
mC62Zx2+29UES+Kx4kjIXElicEWJLj/O4eETa9R9jgd2E/Ns429ktjQSssEW425d
Hu5HjsAUcfLZwiprM0jSTjH/scmXQopf6nEVoLI5UHKu0Ojp5wMwtEAptnFBEs94
MDR0XzG5kTRTYZ2/9TkVlHRJpGmk7AfVauVb4a2gha5Ybxd4oGP4GBhQ4nb7Bad1
MNPOcSC2pl47aTlfSR31gFGXIe+zhsZxagvnRelFRsGeF2U5FoTPyh9RlDS4iEIB
cgD7J9tf2PeL1e4bCLX16VdMBkZjujFQu7lRdZmz/lBud2KvfvKOjptjxs5KGOVP
/tquBO42mNHldYJ4/lRprt863kYy+1qq6otse21zFNRxYQ1KVSBLCNNi3WmI8hNx
1loKy/Qitsgtrf2RCwroaR7zGFSgbFYzx4DcmB63JsTFPZIiU2ScTs/gd0k7ZiLo
BkM7WhoorFF+UgnKvlvZchy78RFmTMM7ln0vlqRnd97IZ10pRVA1sHMlRuv2ZvyI
F3GjR//zed0PbkVPmAEPvMDqMgAgKr3wtK6M26u8WKwrLzhO9FuLjWoyR10kZYmk
ZnAHAqpNyhq1CkkkJ8Y5ugRkOyPT4Rd74pHiDMthrdDkHNno5Z2CmxkMd5ChtnBx
sqIZu2IUIA6xvTerkh6aTJx0N1SNXe42rvo4an03ZBKL8O9PBxHfGDaculO5nQAZ
81xviPDoKNJNKjkQDhXvHSkJ4QlJdJ1YJloKNnK+dGa33FFIRW9KJUn22UYzlEQI
zHPPHcYylEh3wpOG6zr5WqP4USFk12Oa2bN8bJ8wDG0OgwtkdXWEM0wZ4EDmPHDc
Km2Fid750JCrRqqQ83kwfcH+vMVazPz7ffLzwVFGUj2eEW5Usq2tIoT0/xqy69zf
SrJeDqY8XfiiuPwcncnHk5lpqYiNCIckmRYPahOyG4HQIqn5uip2Zo4zN5vVDxRT
tO+L1u/Mro0WTw8auE/kPgBCVJg5iLhCHogutYUGhApUNWN93LXj9Vp1kn0Q2F8a
mMHMLIWeG2amhCP1+mskINgZ4byP0+XCe2mp5I+V3D0qw7S1AilCii8SAZUF4RyN
qfxVlNI1o1c6MTxu2xgoJkoyjnHhiEOvl77KByvooVGSnKcMIBhAIMaBNyXvptmO
q2p5bp6+LG+7rBqZ68NyxaFkVS0oUDl25v80JG6z5kPByqEmOhWu2x9pmmnXs9nL
sQkyzCXFNql9W4XipaByoahmP0bWW4fiuGiQQpm6FEhkAeDOfpL/P3yNABu+5LGi
qjNEEzlvxReRG5pJ/60enhPOz+TiSPqXWMwo2+HfmLvqgNZJ8W4qBLZAqb2j6SB2
tAy/H4WLEes049bPBe0ZIGdqxzpovaV+ttkBoFIDT/MzcCEfk28FWxiSxR36rlvB
Rq6EPNccz0Dn67vk95o6NTX1Yo/hEmkI2efv1iZsn4kUB5e2Wusg21qdbjse8IUC
8vvqx5ta/44ck2pQqtaxeFG1lBVGBWYzLX8Na7I2tjNrfVzZ7ZB4+1Nb0HMKRHv0
BiIXVWYkVLLm87TbPfFVdxh/TBboEZUnAzWzXqiw12X7Pos3oiOgQ1jch33KkM4L
j5YPFnfZpTTqkYR/4h2f163MD8ztL2tSc29xowxnSVs8HOleHJ/4dS5QyaBSHhZP
69SC3GEN4xVK7eJVyK6dB7SHl1BQNg+hTlOqhEz9vqZBhyn4WdgiO9Xjh+AIl9Jb
ggaFa3w7uXJx7qYkKmXR8KHQr+5NQewy0EODqmNSTJQzAcgj6/InFr/+haMvVDrh
YpM/wlGvvNVgDfsA+1sAdIv5n0Lcp/T74gw4tYqwnRLIL0q3bF8Mc2mKJfEeRaVd
my5eRfmbETkEdOcL5dC9Fc2emiSeAkp1/0nHxPaMNpL9kyZ9sEhu2iotkosqbIVt
/x2qKJohrSgsBXb04Gtl/a8kFgBYC3GgWMnLtnPBsCiLGmOKj5LgwtxkWCXrltye
dXwUl2DA4HBfrzF2YN95TTiUn/OxNp7x8kkz/65kf5v9qYR7ao21eG617Df9N+xo
PwzUCZGKfAi9Lxd1RqgaTNp8AHwaTPyw3nOvR2rOwJauM+bXIyGAkCVbzh1KSblW
UqZ5yxBnpn4zo3dnyMaPvus+8Tctvm5slTWgh3uIgz41TVvIa4SMMOT1w3q3yV+O
3WdHdAsOQgktTetMLrOd6z5GYsCIMXfFt9d45I4Pz20F05wEl5RwZsMAPYwV7zY5
/htnJ1DqSEKdce8ByP1ve3Wel76mxQ+gA2eMBhs07zJi2xPBJzyTo6j/UsL/AjfR
6fI4o+NibQENLvfDjpzy44cMDBSrmN4MW85a/O+VP2VKfK0CAu02QLPwCiUrj4MV
P3vN0XRtLT2Xtz4AA1S/pEnFou9IH4up7XUtGiPZ85lCYi70hLCMju7rYLrPNS4F
//3CMrrgGqC19PBwGf8vBdrnXIr6OC1dMdcuJP9O5dS4qYfuACeqSPz1rSzg07dx
wYKKWSOBbebK9kBmbCIl/Kev83wTXRkHC3wfTe6DzgbjFav+3TpxyjMteTsexhnU
GrT7xMxkYZFCl2jOScyUHOKpbNsJGnqWWRCSNJUnGCMJvsL+KRYRCoM/OynkzFGc
yuCqPuGPoydTpWs2CCPFJxGNH6BKpo308FbaTk5nqNP6ZLSV43041CWc3XuwZwIL
GMZeFHTpq0T8/p6qLZWkua3RCxhyS6pDkiBX2O5QVWIVv/+QzWMgzYOMbdqqArrM
kK7YTTyBsytGjPKzyp4k+n5TbYIGRM/LcScQBz+bCn36igKJr+2dH3+ezJdw/ms4
kxN5m0xJDNuMDyt40pkZIic3X3xhJvLfAGeJYz3QEJN8HWdmIAY+1e/YmtzAmWQP
pkAtpd8xhTQgycTymikFEkgaA2A59z6RDrSkGxI7IDCV0IWoBLKU/BJljyRiCn9i
RF9CjmjyMex2VkSY4SVHpjRh3q+3h8EiBVf3txo64ByJwglRxzR6DXSFInfZsG6H
O6e1io9qN/vG9dCb14jx6o5fzlKpUxjKpgQy6CZyiwrGBaxC9IFvbyhLEq9/BW0R
CWg1Le1hMz18DuLdYz4P1OmoG/zWO0LU2Ogm5Gs2yxuZksisZHxm+WSEp7fgJx6C
9Jd9TVvNRWw++DaeEGkMTLfqqvygQP00zfvVtVgEU0sQrXup62iBtJ2CGu8WQdc7
zZW7H1yyXY3LVUd3214fber6o87yllkHnzh7bGfDDZLMLXygwUilfZAi46+eTBiG
Jh9M//Y8YifX0u1sfJk6U0/pBSHdShIT9HE1/VrHJcQh22pLsdDkTXq+xeTL0Shh
RRFBR36tnfajVXSGzORFPJx3Z+oi0k3DLrH+gXHeu7+Njm3TYG67t9eWrWOoSNYQ
TWpQfFzt9f/sz90ryATq4nzwmp4rzOFJzO9WzUR8fAy9z3WBj5F4i99TZrS+EHqD
4c1ACaUzYzqpoGJFVY6uTLLwPoYayLTsxTvSIDEmXevxbwfBHRt5/3fu5/noWI4y
1TRez2LzMewcOIErR7eSam0cJkynr4wpW65DJ3ZVsdOgNL2o3ntIBnA58osy4GIM
W7gRhGcCAIlh+Hlg1XPfoj57xCwNq1mSUjnbufHaBfD75NMGAyuDL/V12G2Gxkro
L+yjIOU/HcDuB6CMzvuiu9V6KCXN4Ft+DSjiAViB0Uz/FvsMetNoimD1AvYamdOp
+HuwJYUfyuPzgQfaRnqjM5Td+8bHy2DamsRCX888w6gyPCxUf9ekl5V3rONcDQNq
9mlVmLooAOMPvPfK/9agC93y8CU6hoHunDMDqhcuOOqGKysD7qlipOga1iqP/4nC
hKfAIUZID0XKjDWYPA4hRHoMJTZUs2wRMbX8KuIVVntLiXgnVaEwv9RVuGdBghlV
mcO0bNZl+/N+CcnQ8h/GleEpckJ3GoaWGlQyDyvvNied4t+mZaGyuHRns73N01Hp
OA0smfsBXL0AGqGRYEaWpdaM8S3y+HHfn97RxDAwX9Yw29bkY3PcISUYges1WlT4
GyEG5AjHYvxPukRZhnaVwwGTryjvwgTBrEcjNv6bLFsItI/4hWmvxFUAcVfwsFn+
vjCGdRxKzIYAmq580Ggf7RbPn+yXC+khMMzoBgjRy9SHksTh+krPyA1bSxC94qG7
R8QDS8Ft09zyExZW3oCmo676ju3iH46pvZNUUWHhxDDmVKKlqFd8haYjMpGzYodi
Q4y/4nA7DZHmgbZd/fzvym9lqADIq00Je+DUzPxPTxY4wqxzZo4CG0zxSI4yGyYt
DZLI3s/rxhtMK1C+2q9iv/Z1il3vbD8JhF34Li0WwK5QQ5Zs+3zM/GcnBP86y//N
YQ/chzQQPHJcL5JvXjQFqIVZvSTQqWiXQaBI9tSjmXhZn69OTsn0IDpblfFQb0ox
DUF3shMdEBka/s73P4QTxEkX+D9qNnhhR51sKesqZ+lwhW/ID7Jv90TCO4EDYbu8
3RzQiNmghxkvNYgMcVMh4v2fO0nFi1CYk6PVGiLIbhhzcq8iSlZ3egKQFKVbDPRh
hDoQBG57dqCWXskSg96VrtqEsZy/ab1O86QpCIujsorOpSQ02ffUXZnAKWo7/C3V
kyLTfro9RQIMObXXcFf4Au9mpE1Bnf+AN/ujbpuhcweCXLG1KNIwhUul+eSuYgxD
yjeDKyGRWndsKVsYKFucJYqF4p1blROy4eORoPx6MqPCGjDPq580ZjlSQxuUseOO
vKTGpoISccAmHQECYdR0weqfdGmmNFG99AgIWrGSdfNvOgasfOhs/lGmLrbh0toO
upVQ9JpEpDw7dcV7pi5bQUUOkCo58H6tg0+AdLCnlhautEhgLhxjubkeRaXPUdPm
cHQVCYr6VhTn3vCFrfozPcEZP32lMIY755taNnTWNS5/o0cJ1Hr4ip/1QyJH0+ky
e4mafh9jlR1yLqCXWCrXG874o/BJL8msgA4ll0xv5CS9C6MrfqdAhR3tuz92GLS5
DK2kg4DYJtbgpdBVOPnfP9D0UbOks1o0rbqTX9Ryhj0PZ6sbp8Hnh/RrE1h2KH3/
A5rCx4fUnw2ktg2S9WHAftt3siQ9KNd6NLlNVMIHb0/3Y6hghaGEgriz6MUAgOha
/35UEB2ztoBe4EzVm7Q026k0KoU7YCF/wz0gRvIPdfAr/dX8Jexpuy84sjLjc5AE
ipd3tsDFkoN1YCRHNq8eRqVzM84x+LJUuWvxTm0s0erSXdvm/4HKMEFsBNQcLZoK
xARotHz8et4S81/ExqXVJiEiLBkgScDh5UOdK+g9dVTM3SoJktlENtLrWVK+r34P
7rMK4saHQiFU1NdT9n1VQhDagtmvh/TgjvTU4ZEGlXmMJENKqnph2m1Ug4k1RYJX
IPaOXGgWgIW/lz8OAgeUuGPVBN0SFRkXna7B7i//Yj066OCUsCH7F+a7A/NPS1pz
1qDVIOeFpHoRyAaS+tQkakyh0BLDKJ8q2+dTTZvEWRAjf2wO/XR06V3qYLv4eDhh
BpQFcCNrlEPWH64wuqTAix0wrUUWuSsLc+P/JiEt4pS1ybH/PGK8EUlA6LoWVV/W
npP7Iy8bF4UsbVE/tmmxOAJtk+4TOMEpQphuOsB0vt/taH/nInbpVewmE55qpO/s
E8wt+rDLxmKmzel9jLjLKOCaqdApEhuioDnp62Q8TbDI4nLn6SCFib6iooSL7dIa
GLQWPQk7XJcLtzoW1nOAhYcUXVXzkA1C1dHczkiGKvW3Fl4uBfaalefovnU8dcpO
A9jQQh+ltfa6e/eG6NNlEtnpnoegMq6CEyTRifc/9JoKvDEZY4SzBxIAzubJZl9n
7/o4ukyD7/1muxwUo4oO88xGeahkndqz/lEGpnxKiHXncmvSFkAybP0uGVvGw04P
+V4aYNbY1/3ljPxhjfbcEsUBMrgCFBfmgu053l8B2D0iYkkTo4GJSs2tuvm7ssst
yLgJTm/4sw3B77gdEXRqMfxM72+8pDiFKjsarPC4EV93MANNJdsbscN6O5Empe6K
zaSqIMW+qKO9v5msruH7ZI43CDCn9zoaV0iD35YpU8hc2qwYoOFLyIgTubRhE6j3
ePusL0OMgA7kyChUL0zxyp4oJPyUDpgCjN8hu4bB0VZGX6MSvlIwoHYLQ/fr8cJo
jDB+mIa8NAp2iX6NUTYShjRe/wSAWcVsB49mhGB//aKOd08U4vHFKmzAq3KACdIg
UlN2/mQBcHwSexSq2KftLPgy3pMrDLVABeTgn36ISdnVnzcShTd+5ZR0NF/6DQ/D
8cIBlPeeYkwKAEUt2buloXgrxpGJGDsTkedFPNvXD5Dy0qJbmjn+I/JZ29O8cJKt
BOK7dPZxn+WA5QJoUDRiXr06Vlie4UfeLGN/QcFI0U1NIVOhTgAoQwQZz5Ob5bP/
RscZloKecxEkjAQgdTSxehJxjpGkODQiP+ceGKB3iEGMI8DWdvT4liGyEa9npDut
kZO+lDpLP85wZBquBVDYbKwFGw09mVuBbueSLXUK7Wz6b8s/t700xTKTViNJUYhs
wRSOte3kz2WazHNpqxv42Cj508XwbOTSwTLZojLJUyWEqSXwLYqa2kobwsb0wI/j
g5qB9mho7/FAyaJ5bo8lf0Y9us0yuWidhT3z+BVfqXu5SEogDgcMTLpjMM0ZDV8O
GLb/RapC8duAI7sdZmI8iqRnZ0lBNEyvh1BtXPGkOAryw7fLVOK1eXB0lVB320HG
ZevuJDFIU8JoXltwsd0VrPC2nVrgFnEpIBrnxaZCd0Otu7phzXuF9NSqZ/D/BO7R
zXqe4ste9Z4ufL9onrAXqaUnqJMSY8z4WH4aP7o8kNJ/xQCod5OeLsCmbEF4QyE0
qS3GB+2Gmdq4pZ4VVKv2+U3WAuuXsaO/DaEO/qNxtrWLCuwy5Nsqx5BkQFDXIUJ/
aRUau98enULyhjOdd0UrM4M1qqly8XRoMjFh0Oojf/8m3Lv+N08gUXj3sfa6QSSK
cUilAnq9B1yfaEVlMm42obxlecWjvBK33HeOUXFIUcuUfWN9Vw+qvpt4SadTzlyV
J2CAni6DYqzmmf7dsp6970jcJi5SV5gyQZQQpfrrN2ZTIWiHpZ65wBDM6Vm48rw/
R5rn122cEU1q/vtQHzC4HIg9RjNz/tLkAxzFQutdKZc5IW53lHWPu0RK4Dr3T3uW
EU/93qs4Apss0OW2B2FQJhO/6IFwhusajHvSWpIDYpIXAhqwVAjDY3gAFiyKEvNo
+7iULrNrDyNfxSOMMrZ3sbc/S4Pb6OdO++k9lUDSH44jhB1fmsOST4MgEEBK0kPV
Z1i7P2eVxaK9bC8zq6Dlx4Tv1qKWIx7ZtbZml5GMkES54IXlVBXNE1+BigRUIwaX
Hh8p0uZLmR16DuqxwGc7K7gO1hRfE6tLp22toOjVQ7FjUApIGcwFKURxORcrxRMF
bFB/7sQjU2swPXjeIiwTa6d5a5JESO5FIqlMxYN4Uz+BUijU/ZHpGKaEBbXSjGrk
FJj2M3TA8D03Ta/qQXh+Yp6mOuO9g+xS8iFMeUmaNqxh41ALpT7N4kl1F/n4Ikt7
Wmzl96AVP22z1Ndsm0FwcYNOsnssNwo98PII43jmFbjWTg6k2QLW9n9qkpf8D5Gs
V/zLWVTMg7Gm23j4e1ws1W8tYZXYa0syRb2+XcpbIrbhFjEYui01Sq8ChsfJmXYz
JlhT8pK8MkPD2VLhtBQ2xq0/5eV6I5t85pgje8NfIAX4ozqMZ/AjoW5M8MKz4fas
a/USWVRvjOvpCpzQK8AMLuqpPb0nV0GXnNgWiG4uKyzLE6MpxoJKYxllKOaF+hGd
XESukChYllJbMW5yPgAulZqm8GyVZC2vCpfez68eYH8BGyOI6AhZYClY03QTTm4t
gQdYsbZh3lYElsujGsO8jWyrjg8V/KSlBwy432NxRSZgAU7WQmXlKEp9wrhQVjAD
1K78oveK1/A0bieYMzTPpF9vQl+LLnP/6++f5hup2JrREfm1vjk6ZqYmjCQ9inhG
6YRDWqSZQMS/S7+D4iv3ZqXfX79aV9EgLyrCuFqO4NMkSzwSBDer5Ix9FpI24u6p
JbR55yNLCnWEY3L6lQFxq6gzjgW5cHe72v2grnRLLOT8B65FslDYK0davJGPPCZs
FlRK0yYxFwgrYNTCVCZX1T2lu8KW8VtI4l2PgOLnbus0NSxZXbUBZSdm8jZ5BJYx
+Sb9D29VxcYNC7aQ5CG962m5CdbY1dZdkid28ATcz7bpPi9GqImFmbDZlu5RabWo
kWR0stgWKhjOCoM5fyS5UIt6dx+YHsur3epobMxTgHkngyiwL3aDyIyrmTzupgV7
F1DpNxd16MC1iScXAK920jlBA1oMmwJux8EXd+qFRKzJ1jY8Ncm3Pn6lMD6eEMPo
+EBEeHafxyzSLoaOCPaHJKhbkYnxkIsgabncybx0Bla36/swzuJ51tN44/jys5JL
Jhtu3KVKkR1ec37ALfoAslpFUeGMuq/Flb2MSe9c1D0cZRKYSgwPj1tALc6pIWiv
XXjFT3vpVjpLmNRH+RkmBgB0+wjJLYWPz8P0GCYKTfQYKDImbUAbu9bsMG5PGsbL
VG9mTJDy9yTAbKC6UipYGzYdPGx5itTZ3fozR6Z2WoUH1pN/8zLqkbYPuWslI9zU
Toe/lwb4ZKQsPlKX4rn68mT/ta6qx16jKC0aC+/HUQia6UX4bEPi4Jhy5OdR2wCW
kArc+Qj5tKvvtpFZ8bUVoGSBXuugAPtDS2q2Qr3mEd4ASic+Wnp/Y7C/sG5ApQKC
aM2r1iK1LncjQIgzMBqdr125/9CvGR/WyXlAhn8FBAsQWmRQbo2uVVy4lGho1Qr8
Vl9C+DrSV/de2IJSJtNynhq+wpfGe3qIT0qI1oiHwWelEOFW3nPEdg7eofpQRE0T
AJ8D+xcO1XCkQQ0c7q8KQsRwG3udPYFPn+77C8Gh8VHq2t0TesePikIRKtN5Xxi6
W3XeTVrdh2oVoROO8nVqUhxwccX/aXqS1oj5wxx6X73RESsq7fQGlad/0h0m8/8a
IlZrxQZKv6LO8A9WEKrKXy3O9vSB4iYUASZ7bMfv7a7Bfa2Q5zh4+q44usy6jKHP
kIAaIPgbxRY01mQj7pZbtK0gfvAFyh3TybM/iBxUpmJDWBLuVtvptErWOM7VSaYC
D/nJLFaRvtYlpwgeIBbWRRX3JkEPtS+p0/+zkZMqWw+F80atL3tzCtlvkUvoOdtS
tYrenJCd92ZxkvW0D0klTzP3go8uVHXtbMMpAJq9BdbcCQp9DMn0TCL4t0/MLtZ1
TIfnl3luN5gJD5No/nQ/xW62iUWfpokQnwbrfzPuIJ4I01yzfim7+QioLbgW34Ch
FJB4Y0UYR/MjT29rEXuI9e44oR7uqJFK9kj8aCjex3waESl3sWu4eDMzOL7FBINF
PAJ9J7h0QM5f4/a+DHHntEoNWzEBn8W2bTSyerrD6Rcu6bMdPgOFA0PBxK1CPWEL
fqdurr3tsSy5QQJHYAAvEFu28QSQwaSDHrMTyce+I7qhZK2lsm/tJ26R9XepRvgs
0irTvC/74ISyWqqzHWybUD920WOq5htF8w9lLUgtrkz2sCYPSTuIjw379eiziT06
PenLfebe7kQ+4/VC9rZ4lUvn91Z+goFPXxqJ1ZB8u0M9yoUL7AYbMExcFcRx5INy
n26l060FV90Ws2G0VNhALXD/wGjylAY/tPKyxkHlu7XToSKggNBdEB/ghfJ4ttAE
LUbe8n45d8rD/ALH+QeCcDVHOhtyuCW3RBFLYv1g/trYdhGXbOl2XeYncgTSvKx7
DRkdYJTDt3zkqlKUUaIXboMi2+lQg+Srpy1MVO16x2fXajw3KXyL/yM9O6T8GHoM
BztfplS1I7A2m/0/dEhnQwMLEPExkuXFA7byR1N7zcd8grFd0UhkPtr5wsGUb8m3
dXd/0yg5Fvc5dkpIGAyeXJ9vhGclhiC+4oeH048YzdCfFnPnSkk0JjskdWf4ttYf
I7TcdGRNoUU01a/kvSXaDnOrs75X9pF7I2RUCMX3orclh5D42nq2TQnr4pUMkjmj
6JcX4cmZNT2e6JH3UCyf1dKJVLUCRPHv6aqgYouq4dLbF1ZqkAjLZEEJG7FTY2Lc
WOYoxbOamZNDjp8RfFeHjlRFVQx/kgIF5/ROHVX9mDTRknUfnoNOQXCH+bGonfca
2xR8s+K3ne+769+KgyU58OZJF+2yI0fauDQN6P9sXDXxWwTBJjp3pvFOAvTs84w+
Dt7XLR6GatpHHWAg7QovuhKTZEX6nA71HZuy8mBP1NaS2Z2IjCaudsJkbYfpmtIl
w9x/ZHVJ/HWW3xetTC9L7LBqk5kNQEHszpD0/tbvsNcX8mTq7TY8p3XXQBjzXdWB
PRrUCelqE7kR9VDovnjfQsf6INC0bApxptuHHJtJaitdrXOASykvlSH0INvkiibK
HurC/7R4GZ19gk3mXnOvIkQ4OlqZlnNAScHcNMUBJ3rUhrjYhLuVilrtEnZcNKGr
vqKHGTjl1p93k6m/mdn5f0b3ZHb+cPkHvrW2ccMxT+/I1jAqN0ZndW0/s4v+v4Bn
iVcAS4mllwX/cbNC+nDeVuXKMk6lJI4XPVUAM7mArZEjDBOPxzlfK/RizHbP0nrZ
aoA2QSyD9vB/PQ2l5lsicjo6ijU7EpnqIrPUWaVLiXcFGJ+kHGYNvib1h6jYfWgg
xdVOYeyXCZTkEZfr8uupC00DOQo6jLhHVj3sdLxIk5WuOEaLmtczzfihvvluZfn4
dAmEpdZ1NEv9PRpFrY0v+S2AMp4sBw2KhMI2dtx0mvkU0bgmqa+U3LRZvEt8hspK
C6NZvcSt273G72wKJOjEOsiU4g6gT4QQI4/wKfe206o+oAtCKdI/TRke3xbog+SK
Ume1Ms/SUNBSlbExCpaBMrlerlkEPkXZtQ1Q7DmZb/qo1+AkKqS7wRtdGQPW9fw7
KTfyYjpE2DK2jDeq1SEt/mxAYbKZqFH6eUDZpND+9oNC4gm+12HBpD0IMNVwMa2m
3yr6XeYGlZOToqb6L4zjFIuuCQy7HddBqbEI57kwzKXCzGRw7T1IRsI+M0uHCYD5
U4Md4vfnE1fXTyANGEnsalHxqzIbiSX7ceGaOkkOzo519mjDa5swqmDZ2K6/ZtMf
w3feFXRLhYKTZRSGhCA8Fu4a2PqDPaOfp7MIz9XyCn0h8Nmyq2kUN5Okq8giyQh3
IOBfmxwHGx0/xz6J/0ShqVe2upjceORPbx/M4Q3g6j7IYPezseyb7NfE6U/IFycw
1J1JRmVmqOltrq25JuMa3061vb8LDtqT5nsOadggREvWZNeGnkVFkvTLuRyUP5UR
Bi8/D15tinnwaNbCmnt8IOH5ntbpPcABuCd35sxFb8ruQD9P4v/QVM/bd+swqLtA
ImJl5AM0UnMUmTg8miVM6hz9+QdRWliPg9ebNEIgMdgEG7dE9asFQ7dS1czSYZcc
sh8mPagAomnwSpGU5hxMADNGkF+5MdO1aZSAdCv3He8ZgwWrg0UCxB4gAjztv3iM
Mcvw+Fw3WVlMTJV5fry0X/W9iY9Ky0pY7EheC30rR+lcMdvAMpU02U7Q2nmo6atK
9aiDayUldN5jL2nDe/Wpa7Gd3ZPMCjFGC1NbR6wWXAoyP3XqnVUeW+8vod/5XlJZ
3+gaYWNKUP9gEcf0bfIjV6Vc6fuU177AiASBi2zDPUelRiVGBqBH0IHfTAVPaOMY
Yklb47qWIfSb8/TnnoCnOiCp1NYoZheyZexDmFqbW1l7C0/MZXL49h9x3Eiyi1Yp
vvAe/9p5IhlxRhmiilxyRQjjYAIrM0nNtWiKSKDebYnnGwUBfhz1BKsEFEFK85Xx
1pv/UBX48tKXf3714Ja0GRNAWfgXrWHBIJLEk9TR9rfmalXNOv0tkOuv/2Hmz3RZ
SN8xSy/Itv77Sb1Xi0cZ5WGPyknkHUKZchFU+w1W7Lkp9XoGAqTRCULY1xRjjj5c
HGSJpj0/n0PnLdKfIX5bDlR9L0xFajI5h/QFFEj2HAO+mxS2HCBwPCzzKC+DolSk
JkwnjZwvYJLYHCSPQ/zl3/j2jrxKhtJAIv0pSJQcufTw1ubgK5AILnnoR9oO/YLO
slzWAGlY5CuM1+jU4iKd+03tjuBkc86HWS+hul6o4VsSOi29VCncQi6hzFwh2FGa
Cn+4tFq2ubz9Ku3Lg9SeqJRH632mdqXMld9EXx6x77xpM8T/srj3DMnVgg73pZIh
YlHga4jYPyfp45p9NIj8m4NQpbQm52IG0MSEf6+tKNff52EULBCxCH83Ve4Q7sww
OC+HgpKzTT9e3z2wWnyzx2DiUFA5mnDrUgPscxGWPlt8wIJEhV/sl7ql9s27k+BZ
CF9H+HTHFj9NqHGSx5uFYqfFvcDyjxkNEMobQpPWDMYnugnXvb/DrIJqF3Qk9tTB
LZIuELYTBjG9F5BdcNmD9YIcqIJto6noOHbgyNDtDT2C0Wa2Sa41T3TDKw5AFTHm
Fee62iecpkjB96SgX2UrFFHYgj9OqnV5zU6B071UyS4ksmmJuXx/l2ktJJQmDhn5
C11HSuFb2ZtUqSTG8MLmCM8jJlmpC4EULgtqFoOdVrzayWPHytXhBf0MHp+rDsFZ
9ZWQ0+QQgUo6Hda6KKhHAxEfUnEiTKR4Kq+Xxk8M6REdEqM3t/GpPqpCkel1fi0b
Rx7tIBPD26iiTjv5pjWK0KTYTN4AMnK9VLStTYh3JkeUb/lpJ+oHW8fhozXgbNE3
JnJcuOnGteyy841NFja5qUcQMAgvLE7VUbopWRDyUXeoWokbdi9b48xSmWGzb93t
PlHOaSv4TIj9yWhqBHEcnfuQHm7jCIUxQ7V/g24BSs2S4Br5DVw+es783iyh5H6W
iu8WFQ1dxPMOypUgwonvaf5aZBd1bSsIlNdbRdPSKn86IvUWdciRI5E4nHOS3CLk
MqJWj1EDyzRUH4v76NhJVqX7nFwWhVpZxvVA5CpqT/lTKx2kFG2HADq+27bnGqXI
9p+Ix/SRLd5TZP/0VERtYNM4OTM/zGV1sAJzMrIt8Ga6cEbopmBHx+jzmaDQcTAO
gle3kFKtfdY3njgHL0FJTMV43ItZq6Mq0h8OZgoKRdnuer/30+82Re+8oaSIsd80
6Siwrxf9ecGzS4NhYZQJylWygbSdESkGMi6jiqJEiXrzFmqb1+EsfsJs3aBgBlQP
NHYXvE8P0v7f8IXUROZOhCR8EvRHgs12x/a+9zFGDT2FYgnhFq03udeNAmc5yCS1
JOead7RwxAGD2v1hTrBZvi9UcnZex+OwDKSNpAZEwvdhqvDgNXOcmHcAYqqqlNIf
Gmbagt6KYUSrzHZKBbgKxbxn2ddEPT5xxPJBQh3CWVxLlNbCvy0poUEUbEuBnPhT
3hZfVkAZhmKMd7/f8M3QpSOtr9TValNDD5nOBQAYD3W9WzQb94CDZ+WpM1b2XZFS
vkJoxGLUz3DwDdBjnMpt6jTj6f/lYZMaCyiRv3dmPfHqK9MHdr9lvKvWA2ziLXof
G2II51BaifZShyTfCiyOG4jDsNavK1h7Q7oxRpTLPRfORFf5BfJKpLPkry9BycGx
Z50XqjlAE5N+q64b2k78eF/AWBF/9W82YrYKk8m1/9t3FcdLyiiuSc+cjHMxOwiV
XKEntoD02diAPjIdNRtRC7AywP9JIb5QJ4QQJsoDBy0C54/opvD76609h/OkjwKw
Axy73QeMF0gBqz2XIQew+xtsMiUaWyxyFHsSOTF4Im9KK1IPuMxCujJvn+EJnDuV
fe04BB0Y8MB0+K94fdov+GC15WcF4tySk9RidM9HinStZrpVCIAx4CfRs3HUmW9Z
x3SjyjAC3CknBBEyE1xEKe+b2iikx7mFJCrzUhxwG1kfW70XFmZVORIKo0nLOnoc
nDBan7G8VKa+VUH9b4VfuUPelgQzRJnMnkaVjsCCvZctW/32487Q+X0ar8lBEz7D
nfv/MzrkOQDtc1ImOD5vD5Cr3AcGPvql+EkEYFFl4NHb+tsEr2QGQTVYiXBLnUXF
i7yW3ZZCKg7jC4K9ZBmK9KSAsxgHdqUkOFLYAKiZ9/itAyWCeQ21gZIXDZtTNrii
RqWuyhJOl+0d/xPkqhDeoyloRJNc2DUMMWksLrUWpxiNKDW3dri2dipt6GynW4ho
gCjeKawEF+kENImGLU9c6+ThDgv1XssOYvK+YoQapsgtEgjovNQOPIS7N111lb17
YhKgKWAxiWIekVGBdHC5iPuX5jizh6DUXrumF+fAk3WSwCK7PSfaNbvLYN9vSyr5
MijqnlgrhDgnfwUJprwWa4oVsFuEyjn7fENKg4MAc851xYLIZ6i5xzq/vTF8V/ev
01J4X6XuOCFlUQ4b/oZHPzalL7GDYokf6JtyNDc/b+SK3rjuVwWksMlveEU+KQFP
PBv0ViV+CqTvSKqIMccn6tqttf22Z/0PWZrr8iKsfwMlyET4AQQxd816v9MLqEvi
njUCY9kOU8bin0+Sey4ulBAzTPFgBZ49cNocEGOLsWA18aZF3HbzJNgRksjCSve/
l9qWOztTAvCx23SGz7XWJMBAblMAKtO4MgWHAHpmdBGfBdKewgo8XkDh1LXiDbF7
QBgaHcf3bQuHBlhoR6O/9qtUlUL28yFrFQN5PS7XLOaQZKvJg/iGNC2gECvKeHrG
dpr1EnodLHS7ohnRZw9m9QjAgisl4Rn7pxIMjRsSITY3FOcgpt2Loyivpx0kdEpQ
mkqFC1+21uIq/0AEh5Y0oZca+YFgdnG9eV/OgDq0PNamoFJnQBc9vIdU7PB1UeN9
/l0M8vSA6iaGP0MoHLLFChsZxbBVaeWUuRk8XLZEfw/2U3n2UFFMSnT8PXcBxzkP
N1lHWMEj8Y4QgxID5e6DHP8/N0klem5U0MCzjUJog1Gus1F+J1lAJp2C5WBlgiO3
QsVNJ9+TfOqpVcTGRdmGVJ3skBvdrVwsHokC38McJURxdp37Fh4xa2dKL22JR19V
ODsTXlcpQVq+QnYB1N0cwtUcU66TORe/8+lwX90JuYt0F7D7WhACJUZC4I1ccGbq
Bwdj30kAB9lkkagC8w+grMvoMzaAxDeW9JWlgVm1nmc2CejbxaoN2aiVsC990TKA
HfKG6pgATiKmYJU+nxJWO+p3pSMJkprTOQQM3TnJrJINWzVbQ+84Z2GI1IuwXtvj
mNQsmb3jMTbr89i1E7xRxB60F3wkwI/uBoZU0VglWStmcu8PiO/ih5XihZX+m6PT
REHPwLcelXx4vaik+jqTNor930U0rjSCOoTnUvd3miTFFY+/SU1RTg/Le02a/7WP
RegWXkJyNT5YVPyBHcsYMsWk9nXrkFAV5xZ6tKjTRdHA00aKLnBKUY17u0/whSSq
gfB1X3/0yG2t+VI6tnPVkJGta0LQR6rtwFjrIl7NPKGzsVjInFEyAeULCQLl9tdT
GPyDo1yi49po+44j2KtLdFuUGN0X1ri4Or+XQrg7bXQMYg3fnEuHTtr71rVBj3AL
tY+qRfxB9tsbbbb3JQyQDbKYZnQ/+gcCfjBg5cG5ZXxvTdqfc2pst4a9m0Xoi3eU
ijvc5u0QYNIHQeO9HikT4xu64fkJVqqmRG+w3x/LeKxqmCKy3Zb0p6jV1OeKY11K
WK+JDifcTu/X5bxfnWn/nh6Mf8GN8D5C6KA6uAxYM/U8+Y/NEI2Ld47RSSYtIQjY
kpmABKz0+Zp6fc92AWSY1GGNhooWYqLoMS47wQugy5vAmP4yLANq4EXEy/p7HoJa
ctiOzZA17ccv5KTy4LBxd/f7H8VfyZ2ha5eIDdXUCvYaRZuyDbGNrRJqvSU/EmDC
ZHxbvUEWE7rVBPh4E3JO1rWQDPlnZrcSukqAvuEFl97Xw/o4FC6S4jNmFyKgzPcW
va4ebc5GkCLM82i5oI+zsWSzzqJyEM4ahFoTyLwaszQcMaHPC4ngiU3TJFhXunNi
c/mqB29unAMZrBdtRhQlWowFf5UmxWErRk7nC+VEo+pXzHxEu2H8ZechB7QWbbjn
hRcwAg/2YsaWLZR2ML5XYNVn2vyDpARWyNv4D9YxWRqKRbU+um00UWOgva6oix4A
B+ITxdOosa5hwhi8HYSe3aqsOhQIrlNtOIGz8L+j6NKEU8PvaMQlL1gYpSOJ4Z7l
/N79TFU567da/9VcmWkff332XJNgsbFv7sMH56xYEww/9wsVV6SdBkVOKD9q/CR0
itP2Q0/xc9BFpZpWJJ6/2ciXzW0KCrFIpgWwPVhb2bpCBcF+XFrSwfHSk6zu4n0X
3O8KO8X/Ha5q8Yo63lmCaEjlo+TSKrPzFzXSe2QwbiQwEVOzwb+h5LvkGOAfvRW3
NgYWJQqPh2Hwiom8pjmyn0za1G2+xQZ59c1yOFjTaMy2IEDGuapfWCAc2NpR4cuK
/m97HJMzhzMcVJ6dL0OMjhsbm57FVdDWb73pOkvQS7l9+CUHGcVhF8ujpXRrvkHp
vDrnTLVLvnngFVZhkU+IJcYByhsgs8wQvqul6VBzs3i0awg/WwhGj2tW880FRbn3
dGd66m46p4RR0hmtF4pXs/JwEVXQHrvLbnMervw6dbLubKvMZlb1405Y5AuPlvwg
qgtLmC2nhKRftkyXpDn4jJKFu8SApJNo1WfU0XjPYh8GZijz6pcNPLo9n3cB/EhF
8p9nbnzC+64RodX89YYaOsoYCCc8lUa9In2M0LEdHoGYNe5HVt5j2VeyK0FB+bqY
owSXM6sRiCth8q6o6w8dr3jYOmJxRjQ92m5sxYOutpHFI0xamfDJWBkyZzrhi2zX
39ChyrOxqgVvBk+0MHFOFw/6lsNRBw3swLQD9+6TLkg0hXA/1fTQhmmoye51Fqa+
aRXEJSvwa8cfibCHBxRzvebcnb2Md4ZJZCmCHtLdjMf7CLLfOWve79Osexklsa/O
jbnrdWz31WV5oRt6H46heLS0GwJ8vKeDhBwuMWutAbsdPCFqQ8EFj3Nl5+PwOEx/
RnBC33yQcTkSMo12TAWxr+ckJFERnaBz8jI+hDSk8GpPROw0wIr4jQ+EtQn6R6Xp
9mnm6A2OvdeZ4sVac3mXijc6JW1vZ2RdS9DuUR6pzm0bLGvM+0lt8G6Jq/N93mZc
4sfc0div+Rc9NSkh1Ij0Ar2eVJS6KLEu2Hkgtgmcc9SCcoghVWzTkYqOIi5Zn5JL
r6zsYUPEt6uPngn4PX2OLbapqS3HMP45XH7oC9HJbRtCC2YaRL1DRotS/glQTMCl
t73tN9Piip3QbfsJ9ygA+rmr/6rmugpnfCwaPO0vjUU1bjqdiM8baXlLOITNI+AI
ikkBvvDwEthEgV5S6ubsypKz9FaQ1R490CtGqL8OOERtF2cFuW/wRMQSAZzr/g3D
b6Wx+0f2ySokA47W7ewiBtdewzjEbo3lP9T0lr7O+tmjncisxqmuADgbDXEXlRb8
x4sYfm5VcPqw7lFQfU6PWmj428hAQb3bMvBK8i5swlpI6rOKZyQ7pKc6MOF9qKae
TlvknR0OySxFxYv+/H7trSLhIiV+AwgjD62wWP4mGAvciKj1PqY9t/JFfOkI9MWd
NyBPW7Z8Cd7gTmngAaXpAP0mVyJPide5eqApQRI1MPRmPy6W4PdRFPYjGukpeHWv
SGEKvr9XxgwskqzwYWCqmd5oo9B9iYAu8YQavqxSpLiH7g7sgK4/V+uPsG4TTyPk
4b8f70FsDBzByO4lCzXObfP44RWdqGA8L/VTk4k4ZJMqBpcH1R7anxMvfGYT8Z4F
ZrOlQSv+XIlqWdBRGVRUHi4bXbq0EtyuQHzMu/qeIADrNgU7gAcglU8m3w8Hoebp
BqA8kn2bPVRuRulP8sI9Z49GltkMelKveTl1G3ChrGziC5gjRYb8wcDsfsDaeEmk
0g/9C3X14LLyXyxKUmfsU8Iwh75DrcXLfalM2nkHZ7DyFHXupsL7aQ82Kc8SKl9+
HOdl6tTwsv8+RvnZ8pIyyN6sr/hySMzBU14aApc2eDLKjZsIFplqWbzCFRCLh0Lt
mW8s6YdYAwKry1s29KdJVRodiYcG5dcVJvxAoLH6W/AtpMAtcoixTCPh27tKJMbd
NQlViOidPqVTRuOGStp1laEq6Zbun7ruP3RZfb7DxLni6ENSN/fc1apQRd54c+HV
NTKVL8/rOs3vYOys2NYofXfv74l5heUtDy/wbdxUrcnuVVoyjezOjGOMj6H3+n/l
PqEA8aUxZnlBsQV3BUvqorsRnqYaIKRgWkJ45+QjOjccuC7HHIQNUcAlTfflDtzt
s7Ul5+CNxfdbkWpUKFzCHSEtOUxeurtl2vOdIOUjaaDScA6TYNVhhXaa01EJON+C
RTDCRSMjVOBQJde2e0AykOjaRPi5sk80QdTkR3Lf1ntufw8KvvIJNJ95Eircu44V
+aQez3abwtGa9SVKBvjCI4cPS54EbV5Wodwuteis3HCIE8Oa+m48wDEQVUtjENuy
u84r9WAXwsBUBV7GdPcY/PzUsv7lsUngmBqI92MakU48azL78uV0NA0UUU+1GBbP
7NtR78fMX2DH4GZMb1pHfJA7bWeYsr8HAIKI/O4sARjv4MWtIxNWFroZV8mV0Ej+
U8O4tpfjl2GRvnWY8wmzSoJxMSppKgVq9ZZpEOKn+lYoL56ScOMfH6whWDgPOOSq
lV9g/WVZ300S+l3xoNj/z5pHLpS8dLHDTbVqxTfPGz4RjYYKTjDxB2LfgapVZM9S
nplfa+asDWQ+L5NBMx7sjMxXhUs/hfNiJKDJGFs71mrnJRN3mTGAQjZkJmMadnPY
ZtJ36aTjg7pCVd1ReJr76XYs4NiecHsE4VKP7PDR2/Mh9pKSRTblEV/dcBJ2UwV4
fWYKRzG+sWbXWJpKjrqVSzt1yD/YHl7magW8vUkMxxxZ6yS83HGvN+ngm3dDMsD2
n0HBGQQe3m8fIqdikLjk7pr5C8n/WMknCJU7yPkwj6KAhvYjqeGddxbaM9aDQmW6
0cfJqwf0o8Z5Ox6RskP/8nDor0n/rkP9S1UM+zRNUw97YfxzJpxT5kZtppI8Ch1A
sV2TU3b1NO/SofDi0PmzNWxGnCKEWS8GKYzFv3/xhG7q2sNxRogeNsaOp4yiV45F
hCN1KQidseQRRbOXkQ5uyFTSDVdLlcfX0AqZH7RyZndN/1xkzhT+XXPyThIyUrA8
mpqBF4KzsG0iZCgWVfLvf/F7XAbqiU9w3oxh4EuD2IqJmvTZVbXL+t89cthpIfO9
fBrVpp5XuBAh2FOQLNL4rsMLTqtefEPfCHOndxUi54+GdZgP4H01wj8plyp4faYE
NG7ojiR4acEyybhi0DBZELpEO8bgL6NExqmEsogXno7R7BU+A+Wqv1QAClMQ59BU
ARq0wvmuKWTwgJdm6/xyKR4EtYMeRn8+URw2sXFiHLxJ+g3kZa0MoV016KJSpuqM
8srqYifYKSYq1f5n+PXKSoovPaFqLIvkMnx+jWs54dTQLM8ObzjLOVBGZ8gLZ/oP
ap8y5FEChTkpkKvAOJlpCYdc4dCuzNL+4oVqAzfhgpVOmqTKHJfAXpBE3Vd4A/5p
e94RAQ5Jyo7Lk0Ydc4ixgihrBfVCIG9ZEJ0VbQamYelNGJMmLXo2IcBThzh898Ml
+kKjkHBFQQUqgVuGGUA2FZDjDmwWZagJsg79Y0of36534mjKQnDQ3F4taJGzJUtg
5As2oiMY5YUh6M3LFY0uiZoWyKliJvUXNtC6t+QEbf+DCE7AneTJps3yWBBVkcR3
hLadx+/0uEPcPxe/iKUqpgDhYAhWB8LV/qnxlbN8kA52x/9VZquMSuAPuWRD1zcE
V00Bv6eIS/b9PccpzGf0FWbz4t4UKkPd3hNRQWWoSFv/DFCWNwwx7IyilTyBXw83
ZfYvgqA2momZ/PvY6iLsDSul+3no2yAxW0QQ5HjuYHJkk4vDRR77uXT9bhrZt/r3
87a7w8iq279gOLMfj++peWSolNZDr7vvbFZtGX2N2Z1PfautKPgqa28wnBc838tR
1QGiTa2kZvF19b38HG1AFcRvqCPMfn+NSoWkf2Bn3RIWSJ5XE46q1pVpe+Yetrzs
3K01EGUmpaMt91g7vQlP1AI6lZObqzfn6QwmAWpk0m8fnfVc4NzrXPN1c41H76jJ
AuZrMVIAlJnm/E2nP+MZTjwruHwaU5RreX77YOuO21z/LSafjK+iWgit/8Jo+gRK
07uAM3HuB4u14IiQT2KRUolL+7PeDMBGg5LVI9utk3Lt6gSGaOwe3y83a2LtkKjE
K93r1wPVsBYzzZbdJpV6zJ0YhyesMvGb1oURkYYEFBhO9fG2INqIpequnUqPbM3k
Rwa8SyeHEANRHfiuYuj7QgWCYzJJd3bjkQ0z7ILXxd29sdZRxbi7JCuDMWpdWSZD
6QyIky2ULA5oCio4DzWH0nNCwXTlL5sdB1aSQ+Na7sOCKvjLDb9vvgr52OO4L3KO
7yB/BqT8YvHt0YhDoDGVNVJdwQGNOSnpX5ZZHFYqVcLhVB7xuFZLcMDauZO4fz/p
5Y4KBDixdBVrF35kEO4EoQT0Tx/3TvZJyYuIPvjgEB7hVuFsa2sNGNFdRI5kTOno
pxcunEyeoLoAL+TI7Ll0uuxP1m+DTZcEPn4/yRvaJ+V4Hx+dwoOFLLNmhKck2dVj
0d6soFshAOIgewmtmuCAs30Ruadq8Cq6Y4xrgWRnKwVKoBqirr0p4rhOfndF6A62
PPi5pEH1OJoSbLNneZg+LjRuuW2s5XNBdbXbuECm3Kp1FzyGzstNjqXSVqm/yCG2
rt8ukxFGEYAZxVij0oTlI0NOm+4Vekqv+JXgLdNMEhwRyQROMSdICse5473+9zb2
dYm6yfUOr5JvjdYIl8J1ZgZB57k4dHdCAidLMGkoEtERPKrQXFIfPtU6HxawHIZ8
cQNh/GH67LD31puKZnNmYMiK0GFZff0yY7ZIGG0kilfp1CJXQ6XUo60y7sDUBOPW
1VCN/1LX5HIjL5W15sd2EHAMwNIhuLDwWncHjn9NjsZ6UbsNZngxIAsJTSShi1FT
rk4Jhu6XwNm89tVZAlde8GBEp+5PS/jVyGwb9Y4DpfKBZV9RsFoFyZOUsDeGlcUJ
8ypj+Zf1rSnkMcEzlg1z2Tc3Gshfb+6Oj0MW3HE+DBxKs77oh4EFv8ayInFFCuy7
I5XyYpgAKYR9oCDL+Mk/5SR6LIgLAUQrLM89WzgbBt23f4D5b87a0ikQwiFUaD+A
S7PBt6wbbI0/L+sOkfHmsDzpI0ujm/ay7RyZshpeIaWoctOMhT0BNBn5Sk9RLnmj
i7hRFKXf4YstGlN4elmyIciIof1DQLOxDfeTuMr6sVJDUsXskYi1rZTPtE3fWPvS
2Ba9+2K0KtJpgfOgJ2ezmdCjvm/N5zjMIyyNCul2oyG12ta61iLTUzrT5nYdg0xN
XNfFNY252IDjBtxsuOlxyIAElmOJ9njFHB4R4WxXD9q6ImMe386FO4q2qXE7T2/M
SJaGQ4T7pjeTXHZp2tJhxCC6JjRy+7Jautnor1Nne/SsoVRtmQJhZjmeDU3J5vEt
2/4+DJNn8gsWC40r9ToORlcrstwKJI+4APldhgfd+OWnyIc1/qWpu32NUl4XDqiA
e/d8BT7zIhpTGVZg/zc1dAWtl4cm0PWfMrYbWW4f9eJ+QmfQRgIA2pkfT115bOz8
5xgTjSwpBqh5FE9eKauk1aA66yA2Z5vjng44lfMsBcIp2NCtY8jy8h38xlds6LJX
vmf6OqF2JagKOrgp5Ahp5OTAcNDtH1U/WHMgSXkbyCZOsBTmPkbifxSgq5T3R0um
riUR+D8t2EGH/x1scgAuYe8fimAi0unS0C9Pb66WrTdTMDo2YLeb+9iZFlEXaI4U
ENezIYsW4J2lgoztpElx+hjw71QSUExNfDkSx8jugIUklVGenpUgNY5sVEnwygLa
StudoAF28v4rTzvRbkKxDwBA3a3l6QXXlxi69xzhjLV7V5I+FwJgq0F4DNJOLsAR
mN9pkMqrgv4HNCdHWsc/O6sdb9les+5G53bT7S/SGPCTOzj1fYAdbN8Qqw4UjtaG
Qob9nbS+kfNfkaClnmKZthlSO/m4kCm++SZFyLV/zgSQ1MhRl7Qnz+PSs7qqINzm
XN6inwOvx5CdqwVcuJigAMh7/ThVk86U1ryle9Dcn0+TDWBysYoFQFa/cM+sCUip
5t3KZAKnplZ3Hz1nUmAkJeEYll3VKzbeT5/TjqHfuOWlOIw1gNiIZ57u/cILUpJi
ekUJ7KFykkCVAG4lzSHrBYBKbSM5VEuLmFX6CWLMAUesPwx3wVjH4N7Qk0rYGn1V
yPjOLoNISWB/fXDa8SV5vrKbtozw69y9ht9jxhDPXodnAnWU5FAv5DAS0Libf6m0
It4sSK4uzPz5NONZk5+r7BzzRyCSIMAevG6FtfZHJz8WqhDEw5f6Zdg3VBN6FCf7
OesDnwp6uYVwCufamt4w35LaOuVy5sFqPaQGeimcCreyDLHUqHktORAoL8iY4p0N
/uXAF7NJcBIaFRpBOTBzkMj9piaQ06FMcoJ1nUutMfiVZfV+6hQAi4sQmDJMaGvo
kZNBKdvhSo522I57YAHLUdgsINApu15rk5wj50kgLcRVdtxcmmuGfaEz5ympVuEc
BmdCMQt0BLhIsJ+iTisP+A2+THOv+a9QyzDNz61mwruL8/PoExOXzm3R/NezyNs6
phvVoNEa1H2XByMqSe1eWJERi76Qwua+M0zGPnwQwaELjTgnQ6hVx0nNOsevanLo
Gtnb4W2XfKhvkxc2SpzBMpaS3uhh1aLoWUn2quYCF4CKoHifqC6BlPai5hOuEDyh
fZwUDQCJsUyNoEiteTQAV+38G7uhHLq3/6iCKfWNI2dZk8ULUXv5M/aZbK6u+Fgy
RWIakxJWKapn6i2el6bMBWRA7bLM32V8g940/dbPEs8LBTzhgkie+A4Zct8r1FF8
BJzaJ3Tvs1FP1XxKrrTyN9LVvRIDp79a0nqhlXFenz4QvR+vn9SNb55ekFxNfE48
/4rD9+QC38v5vn7DRbg3HdrQZv0Duz2ohO3n905rJxxp0nT3cdsgTQMR1YIeysdr
cLz/HcMs0dqNLerGtaovXYJtIw9vc7p/ZZxtG1+iF3eB2Nx5qmvvij59/zwgNIkM
ddmTAkGlXop1tnSeUQ6pzzqH2wIZ+ShyW7bllOuHykfSKj0xZ7w0miRvyZYfOehf
nZAN+dLl4mIfAbs/ly6CIDAWavF2v6B/wf8YHtyONAVMweimTRZG3IMeZbPiz4kd
u+IKGDTccvO9c6afpVGUdYPywMylUo/9ZMP6rhDoJb9TUTOl9IcckD4iiPXgdIS2
L8nzt91fyit81dqnMiyp5uhxt2y3V4RXKlVDXBm+rReo8RgVYFO3V9FM3BmYzFlr
0M9S9CqzTtPe23paj8ExarLDft9wHTzzp25xBTjEceWbINrf+aTq3+p2QYGTkAui
u1Z/5AgMN6Nqs3IbYhyfqkdYx0W99h1OfT2CC67Y5NdcUUZ4s5A2ZJOm+B7xtb2V
qoYwpsmfqOVguXOX7nUkYH40KpzkRwgLFyVuA2cYVjUG/p4y3iTYDDWCA7Ir84rj
kT0R0KVeDplx1IVvyy8HQS4yhrNomsv+zFvuU91+JQ28SRWuWqTjlqsNX5CCMw8/
bpl7MrFVwd2pF0PiImFsohzDk3h0lC5lVL6UFRTmAdJgR4+vMFOQEu0EwMVwHxPQ
k/Kp7uVYbEOhsYuV6pJ0ZWtGl814J3i6Vzf4NklU5wMzcPNQ5/W7xtrMmZfvCXKR
5/8CurlZgcPIL4Mxm7IvlcAqjhFFXajM0lrQH2zb//ZXLnXa1zqiV/30ykxU4jfr
i2q6ARSznZVpjQe0GBxwf98zYwX5BNWUh/Vr9lvs5RUGXIXmd4Yo0SILnWgi4odE
nn/A55r61SXe70S8s+IQLVmJZbq6IuxwOOiHTpEL9Rhrj75X8nkuuuWLAw0H+HRZ
P/bX4VszZpftAMchhYXkaSz2UskVlZfR5R/tJ4TeW0664AJH7e4A+gM5E6VjPWgD
21ET3jUGWcQl9hPrf4JEIcv4tZsBY2sxScZ+RCraE0tWS5YOxiPnHVEBrWaYJuTE
sesMQeNpr12dQv0rN9kKJuGhbw/LiMYGQa4gYm8QBPWNWr+43nnojKCWu6jG4Y1b
3w1H/FHCn4K7h7rPkMVO5IYI15dAMv/MRZLf0xqzPSoqE3STB5GouxyVX/0u93LD
vGv0qWggu9h5ybuMEYOzKonIpusM8uM+EK08txJWVIXp3sHYVlCU8wJRSErGz3Qy
7lAoHkZMEb6RC4WyYbFP88Stc7xSStgw0g+8jB+Vl6H3Oe0ctu6XkEz0f1lRdR2N
SPaAtMRCddWjmbTOJWQM4hy7SwimcdZJjXDz4XhLqZspTeJSbyrPWJjsRPVeA446
zaqdC4+bIJgBCrrlBdBValznH6XPVoMi0oCS8MjXP264GOJ3kl1kcVSS1brjvT9f
SLtmzUNgShvrb3xUiIo+feXDb5rqtYXqchNVR64i0AgsaSMFeXulBBZlmrMzRwgR
oy1rLFAfNFR3IQoUEwaAfVvhVKHJUFCbZPQF8VVwscIByLEE9Mk/KKxZiLjmkJY8
qg7+cSxgWUwwNDkT4XeQgR+YqtbEps03dedkLtMY76Y6EC6r+6yzAPTx6rNnPNBK
v0HXi9mRaDQj+ipLtLxk+1EXAJiC1zos95TskLe3AJTC0Tn26ZmBNq7aqjcC+faw
GwYorNKCo/Lu2/y3W6WN9fYn7uMm9JYNijyWjO9hpFmp7+e24u0n8FeBSYNFMLWO
0uZD9ko86K61FzYTdIw3bLLDocRxglmffOYxjbmk0WePR9UfRByt52bh5ZgoIMWA
N58zjIAc7aJo6gS4sT8iIXRnqhG6E7mYqUEgQrY3ygpvndZ3hUGM6t5wlSTy+jWx
XLk6f+EC9f7SrZ5g0a/L/13tbl16D9NCZ8GV8f1vpaPOyhG76oOVr4vSSERWbJXu
Y0xF6q3CkORWq/btG31aPlS8ZD7lsSLfsBpC6dq5+M5swu5YSdVjRlIxuM1G+ICC
LfhrCJIii0beIskwzPxfWMLlJQE91WFUmLL4IHfih/b5I5rNEe+iBiSHXRgO2jKd
kTjXQVT4ANrWmDSupZZoVItyAVU9bO699DeRw6276A+N8t0lA+bpxInleOU732Eu
bDQbjGPlPOg9VYDFQ0LseKO+R5ktgxNdt6fcoLc8TScmShAawR7fUM9ZCWwyyNh5
DqR9eZEtIF1aUHsAWVE1xDku86zmcXTSuvLal6AhMxeDyitUM+QfKDwDKlXR7FJH
uR54M0kVZRKl2tibUnf3UCvJugbkGhJzbBYuq/FZvI6a7MroUYZEXZ4hwyt85u8i
BHVMTa14MZlThkqLajshpilB5D3HGO1N5hXk49HG/kt9zvoQCrs8jb5YczMfHTpG
erd71h9qXgAPRi4Cyf7Sq5rpQYHmqdviuO1sziddSNlr7TC1fo7I3j0hpXR89euL
Fvz9khnNhqTYigr4y9OWva4nXmGY+JEvQiO1vFlBGOt0D7Foaeff++voxRsxFvdb
Ds21yu1Ga1LjqmiIrtzFgcRErB75Oknn+/w8/xtB4qB4Y6Ay3cIqyugYYq0pdPyH
tC99PRp5C7LrEWAa3NmJCIapFDVSVgNyQo6N/wZvjxHKQjpqMaj6SBXkKv6tboda
utCxveBj+73G8i9v+LjT93pKr63u5Nq4zLFnVay6wFpqeQJi+F3MHvVz8+4TFrQn
umN6K9lyBJO9ITcFMTbV4thGQEj4krSlTtXKf4fjhvEI3lOokHhgTo4bkGOxrPq+
/c+pJKJLsxnj0CDHfIr4E3guotUab24GQPdsjk2z48f3GsNeg7SNjVHQ9QVBTZD8
Yo17HEpQ38A/uq7Sc9RK66Up4XOK0MrDtJV6QmG+usrOnUt9rkjtAO0JV3tBB8nO
uncSCkIjkebW7DOo9Y6wI/q+B4xOKz99+v1T8oeEKrPCPU1mqECZltYkc2YpUBlW
+7SSfw0ktIsi6nSZBh50Y3hqjyUIUeGXOmrT/OjF7ftR2e9xbOYe5p2mWQbAyhzS
SYUc8Uz3/WYXIQ/pWISoJ+YUwIr2gtJX8DHpsCw8L5DWmJE344GM3UGJeiJgEmN5
XQnrcrw9pTEwg29K8Wppk8GpWUlK/XLqRrCPJ9ZCNyM/iTpMWcHvZlOcXT9HEZdy
4Egi4W6Exo5AaD5BdBsO6veWU4UgOdeu/CjP0fwTmY43zMCzr4R2c/AhWaJKh02n
jgXtvjxtXLDhDwA00R9ytgi0anrEKNn0gGn5BDlSH+Cv9SUtdlo3eivC07asdKk9
Yyuunlv5u1by6BO1G/Hh90gr9y63cmWI1MgTtjQNFyNzyk/81R5VkiXH/74gDnXm
dzkDDWYIObCInh6ZfPsRl1hiGNf+IeEO7kZLvTsAXmRkj1fYEvBuzhSoj9HBUvO3
SHcLdLvmThZHLj+g9hKWh2oKhltoJOv1l4ASSjkT8hiDAFOnsEGvy8X97PwkJXaJ
78/DcFGi+O63s75ZxyYvl1M54GlZiMqX4WP2GeQGOFwsr+uD+9SAAlhFiXY1IZH3
9mnP+kB5rulzOkXTPaBygnRiFQHpgekcBsuR8l9qrcanHdcmKgEQ5QHDgxZ4cmjf
eanW9gtD2kEOuencvUtMPQM8HksACAvb7UYT3ZD60+nGMNryuQC9WQwMnbira3ju
Ddf6LLqpQYJpSN8MnJosQN75+7+wtbvpmSdiBD99m1ltoF/4nDV1pH1wOUcX6tsX
CYyqv0f/xHodFYvVhbTXswkl6bexob6ATm4iVBI3p6qMY38ssFMDOAimVysHUJDF
ahHJj06fb2Iu2D5A9ramcKvfd0ILdYMRSlfCg8mqNGTLTOEaybFXFBbLqd4QzfYd
im0ol33JtLaTtb1TKeWyOBnGCUO3PYKDEvnw1TcycWpB6YVv2FQ4dLg/G4jSo9cT
mOcaHSnXUO7wg/P8zsm4OxW7EFozysvzUJLoWbYGXl3dLTbcwsYfO2unzR7TaEGB
0hCqb/nuIMRzjvTGlk3xqWhHBxgkFYl4HuxFX8stlA8Ppp9ZJCn07ujiat+Dl8EM
ZIOvDevrJl9SqU1M1eOtRdI5DILwroyiJ31o+I3Ypyl1llroVjxgnTDatSekDsCd
bQ3vOJNXFjtSwTPKmg0auznXpcqCWjvTOTHxCmVvCZqebLbCTK1VsILL61Jb/jBw
cesqXLkdfXzpYPAHXs38NwE3Myn5yVypDEbOjgy1lQwHeHaICT9DNxg3Jxn9JVFQ
AVYi0rJBPOksARNBrfx+F9xqzFHT4WJk6IbbG12zf1rIEgsWO6dkvE9rk2U0g2h7
bcJJyeqnhj+TBt6h8lL8eCoFEM6ka5Oi0cijo/1X3d3SXhIHCHYUMd2VWDsX1IXi
AA6AO8cOQa51bPiWPU5StfYhazkr05/rbYxrurrQ/zR5rBEjSIPY5jySMpxAHGMA
QwR5bsE/jxe766iVLgfAt6MBbpHK6jQeCQJSxyra9d0OUL8T81QovD38FLAE038c
F6C8RbC/1MTB6plDx/oyH40wviwO4KlB5tEEjLJhvJJWl+2/kfwskGSNsHLghxmU
rdFQFmBPkGsjeG15ncpN6gf5I6M0mQO4RKIx4Xa1pXOrM3X1BAQdwtgeViSz91bP
g61QONkEb2HPkgtwc7OBtK47K9emEQvE6BR5uybl5qDVyhzl1URf1s28qGFuIXCO
oGuGSYJnlEXy6xGMY3y5Laand1O23K+B38oS/1QXy+0Ze5zciyAYeW4VIqPdxd0x
y0cWBDm1CGFO7O8laXqHB5GTB6mwFIcdTUZLS0uiMK+WO2COGlso3NCv7wGNC98C
FU8oewHaoHqPHOZbcXIQGuTwddb6bSIaLUppPV57+dSNmhAfEeSl+WMgPYa2CrdK
84iya3jVKDVS7xf3B1Za0J421t/jEA4SWDcTbnHwb9XTp5hLFiqEWgplKwbw/NKz
sEnuCeHXn9ijUcnQdATqQ7efJd+CaPwLUqRziJmaTGyGCL2wffs/p5O900SXoy3b
A4KoolzevVid6vx3v2TiMtPPW/xdutFGWhcImBl/g+TYNLvPAOew16ECO9Om0rrr
5GZGzDx9ctqqcylWWXTj1koOl3Uwy7fx+ZRSHU/QzdM6M2+SVkFr7Prc/SbKjlmc
6yAvE7O0cMtWsL1JWyWb8AcBK7hShYKgtTzVpq4CXVgZvgiGNOGCAoEDA4Xn9wiN
gwmTmwDJwtWlYp09ab8QrbUdeScPgpWNareEHu2dAn8ChuIfrQf6Q+vObWgjBzBs
i8tqYS2bJdnVZPzlf/0p1iNz9p/q5mm9w6odqRv1b+Q41ntbb8iibUHP+98LgQ1j
KSn5+u6CZAvoIOpg9/O2NM0m2+ZfbWF2cEfPRGu1NoyoZVpVGy+3z0Q3HxmgCaHr
FMrVeAmEDHus+2SZYAvnS9vVgnO/iWTZIs+yXqRGYxB8zdQJnNvoZlbraZJog+0v
M+6uAt28jTDd/vugnkQhFpetaFx/ubZXiDLGpsI2wCqjwnWUVDGGOuN6wMhb1poa
+fIrKwOC5f6/j0Hbmf+IUsXnHErNaR93nUbu3gSWs+YtgG5InGMPxD6oyqH4gB5F
KMwR0G1C2suwpV5hTPTrnewTBAghvbc9d5qAwc7FjCIWvWbxGBgAOJMNZ5EqPfh+
C3azG1mt6YhiSh3fLZoWTieCg5Wa2NhSyy69d5VlTYWc5m8c+p2XURVLG6PBht2V
bOxNiTUTPi0iL46aAd0JLRYdrJPxDI1OTB86T6+TK1zN575tAnHf5VBDP+wloUBc
cjE6tVfvNWt5fGQAJHNCOh/KZ2PBF6kEjNAmS0VYlC2HvLmdoyufvRmzec55stvg
pyYc2LN5Osu01n+yvosc/Ly44YTKQiI10svUsqKjVZu7D6CBUFwPLATOQ37O2u1O
pW2ezRhQiT4Wtfmlzs+Kxv7EjlimdTrTVzo8GYgzc0nG/QuEKZEWxa2qt04jssPq
Cz/HAMmYkc7JU2Hb2smdoet21GqbtsZhfXpehdMi67A/HozaXr9wqnZLIoAdyWeq
4TwaQJOcUvUNybnSFxA71/XcEGg+DQ5wLlyvRJSD8sLRZaV5ha9Yhd8Q+hPGrj9f
rnyHKB5m0YWLhEZljj36AFhRBlNYQFgjAoGbAaM5b/5ZC1RQs2Ry4gGsamf0cGii
dVVgXkekKMO4myba/c8VgvqasR6ic1xw3rHLJsZIFGwhhOyvvq63roqD2Nod7K5C
nqRIzcXTPK+MZhcRK1OBCiRCQWuxkDf31ghjuazne3UyBNhP/SCZJqRJboq+EW00
7Cf1gCuS7Wj0moIbD8apgXdKEBJd6MmNCQyHYu5EODw7CiamDCG5Lgn414uvV470
CNfnM+c5Q/rismHbJ7NdcPWY2F0BxYGnGSbpy27Bcr1AeuerzLVxA9ZDPkUQFCas
Ix06Zf3WlH7GgYxAdyFTwgOK00RGsKw+XrpKtFASBukkcgHa9zPrKT8nrtEIR49K
fF+NmraT5qCFV7Kg2lBQIaCQelAtSV45bHtwzjA5XZBSVOcUIyEUmqzBK2f2wjne
VkBpHJykA8llihGx95RtY8vPlVYvn+VC+NX0nAads29hT18U5lMTuRY6iwBTJSP7
YoDYOlUzq0hTQHMDVm7qvR8+FP8i2AntXdkFLyOQxigZZ2/v9D+gbqGM019o8ujn
Fi4nbjKanQWPxHctH+6I29MGTlzHTfV5q+jqJt7xFuF8PLXCbcwDecopzhG8kdmF
NdMbEK4m6FylULVJu2Gg+oLcRfNYSSOuU5Y71xCgoupIANnEZLLYd4ehKnTg40uo
97iAxHU3zsK8XjZRNgEHWJSPkMyUVySPXbzo/B9G8nLVj9lKxp2oEXwyyXBEc8Xg
dcKEwy1WFhC2ICvN7VbzxdETUXCRqspewkDANq4YGd+U1oJEgM0xSQXqih+IeuGw
KemgAj44O/7JXmjldvIAu2uOYSNEzYQorq0wHLFzGUyzM4fCQuFtz4SaM5QtU5i+
n5DBy+DrjAQybsCPAKnpALMivjgzJgaWBtijMwxBW3fMxdmr4D/RpEMTvh/2P+js
GLSYIEDTFIyNjUbfHBKtMCzu/VZ2Jffo3KCtMYQFKLDk9b8hiBN9KTzA65U58Wha
2bZNDDKd1PlbWbHi6ZS5DJLTQ+eEjYcljCRJDbwb0WOdeGJoHssa1pI9HylBUTNV
pg3KzNSCPOMyNboq589yGYQWcBZDB2qAqjXJDYWxGJOwCp+JIbtYmAlQ6s+Mcvkj
ocbVpdn8gY/BdpraMdG5h6LX3U3j/LpfodYpnAr4NBITI58obQSNwHm58K7DlBgJ
dVB1SdoxLA7D/ykdCT0PWefst1FcVuyiJNVE4oAsS9JuFOY4SPjeLtKuPyzUWobr
OSn+ZxG6YwOaixmmSmXl1Ry+auhzapdzxRMWOXWcmTlDTZDxAmR+6jqQKQf4OWax
D6i4wr1J8tOD4iO14kiRoWSFMlxpfVQpPTmHLtak0ZgdszG4qqHWKBjt0X3JKcSM
6vNfDGya8uW2GMe2VcKRWysrydYR6X+GIyvnUkje0IJxh2jVO9dr1/1k3/tb4zjT
YM6ezxJ7r753rs5ar+6727qmmZNmBl/CdGnXBcVUma4FByC1vpEBQUWY9VdMjIJX
jHL3+D6pVLAd32G5So6tELT3DngNbpzjGWLWGpJegpfgWa6qzG4eUJ+Wq/SxlXtW
3592zGhM9XxefxCwDZIQdJph30JqsX4dt+/0VaOlp7OFpNgPIiqh3rVngOtNNFyW
jJKJZBZzhkbmEidu3tgzQVMmojWxzP89yoX88mklRQBfdLy1jd91Iijylg5sYAwD
SDnqXDx1v2MxYu5mP3NDK/s6lk7J4qxTMEXw+gTlIiC8NcXjz8jPPJ6uj29BD91P
OGKe8mrGkuoT7L5jEUFSDLg5Ca/Cuch9zG3TKcm5s+DESONWYd8Ve5GbfqH6TA9o
lTNRPvXe2MkZ9+bBZARWXmXSa+8GMzL6au+xG15DWZU4URiPiGuzzLEbo48EbXkc
xez3MS2po71uCrUFOA68FNY670texbwmlyYELPc9k+AQGuVBo13UD2Ar7FXvTzCQ
Nbba6Cz9hoArTeYdmo8hAsb97e26wfBKj8uubSFTwcgUjJkkbZ5ryXe59tjVyC3y
/6pxd3Ny13zvF7VFbGIVq0vVp377oNWeDQGhFkqpPAQaVmxeF3agDkSEWkUpuoU5
2sOUuYiHAMwPdAPPRe3IDjbiwtkqmisx7GqpWibnsG9LQR0wcphoNL4+xLlGoXrg
sCVIoRFa1urxQYtJCO3AZP/WY5WcEYY+M1z9ftTqpxLBVUJI6oyLqANV9j3jf86b
SO66l3OV8LlO0eSxPNpcjkU/O8Svz29/MGtxDWYm+RV4Vf91sa1TjmJ8CW+r1n6Q
ONeqNn4jZiVu/VqNEQnppRmUgDER1BDtE+OzrRUWA4guiadxB3X3J7TrWzQ9Bjgi
74y2NT+iUtrZjXwgYNdWfAN77jaFkWvh+kw311mX835usia6zRsgxUQ/a46bJeS7
x5ff5UpAez5+LPRJUdJbio2TyucSXA6I+fQ2fhO6y5PTe6XbQ5MAbFyUZap6+LNO
vEzj4GOfrxY2U4d3Tfo/eDSu1y75pXpEHhyDJVdBIxLiLKqITlyxuXLn/J4ApsbM
XbA79/+RyHOwKiuQVgZfibGcEiSZM971q8VZ9X0WKPP1jwQZ/k6KWSXAywrcCb6o
EN9qWn/cRkHQC2cQvqyASsypcMv2A9iA8bgXZXdfnUQCR4hhzMxLOqCrSbkQ+pOY
x5hRssHi/Ox6NiuEmOCGvtnSa/e/DxRkMaaUjFqorQPkWa1hAR3QRrXCw4dRphfP
5iIvjbHVNGouKUwfom/Ar+VcGG3Oq+YBc0nOd+59HEM4io3SQlGGnsNosRVNn3bQ
nGwcrdPTP0V6Ks393jtUfLtsKT9AVjfqjsqfu6HxElr0kCappa3RYd+2b7JjmRf7
7s9WfLSBxhL5IKXp2j2JCnHclGlM6/uqwkeqXLv2aS59JNRe0s4pReATdO0p8CC9
sgqpztZisUItywFtkc4pHDAna+EB41Z8NOCMLNLbdaMl4iFPEulG62W+1gg36o4h
NAshjpuO6vTaVTkQgKV0uqz7iNPC87c+c5l5Qd4elctA8lfizU/AXS8LpuWvkMa5
87TLKDOEjfyvOcm8Pf+IoZYWiUkB7CUilzC7V5yQgJZxGxwMWa6wKSNoJLjqB2pZ
91TEIjyXzQ8s9sgJ76X8xeGKXPJmQWqxLkt1vSg4+LujopTM3OygJ71R5+/jp+MS
JwnvYhbogVt7d/zcoMtxSHs3hCCkoQDBsvuLCS2fNRQuWavx+LyQMc0OQYHdhNt6
p7sdo0GplqiiBp4Yl1e7Uf7+4ycqFb8zgssXdULLC0A/Oh4g8hrWqGlltA4k/rqV
qFrJezmI6/T3Rek0yRTorXTAxgQ9knIhNldFLKdmMb8mSIHvYHeSmidhsdgwfdHl
/iUCD42nbLb+ttjf84ElVX1flflVdQm4AcXk2OeYh3KJDLCT6+46WxxVyo6XSGuT
9TE1xBJA4bimCvF6Y6zBZgiPBTLaFstME+4SozoiD4CXNwPiKujCuA6b7jxgerxP
rxWVczljt756kDtgO3JAvnUGmz9piK9VN4PTfMKLGe/AoWKcxFHusPmRupb/RtS1
VF5UPMutnV06vXZFCWK/JnnVQAazFnG3IMb7YKtGabGhIM9GxbxLfwcufDXjv2VX
wSN5asd8K7Mlpu5ABFf29d1d/I+jcJertrjRXr4m3LK27oSbQhr4hBZNh3+qUsI4
VHQGHAfdwFRnZ31Pa10E3G+0GiiGCsn7Li07U1ge89ouELYlc82ql5aUvPeP6eyw
p5+OpOg7nWMFMhRrabOynIvQl3hh/oxkobxcCzc45smEetZJ8arrsG+wXSCFsx/h
fMshE+87+aoCWwDhcRU/WkwU8yRX4jXC9/IHGhoxlHAwmXS5SF3PBRnr7ubHAO/X
LrXBfACd2EAX5J0dcOgU1ZYW4CVlLm35ly9rAgCTuJhbJ345SjyhgbHTGroByBIz
gDMtCqJDSs7nU7LAjuRIDLC3B+wWY13uV4tYB2yAcOc2vSwdM0nyYoQgj2Cht2wi
kvDsmDsClgm0q7GvWjKc430/iDEmgLxWlDobIxvlfendRfvUh3bASqC4hnbhHzJ4
9omVN9xcq3ezzD0VCMdo1Sj0s3fWnAX1fzpDCndZvO084a6XUyoMRo5wU2msg656
z/2h1rksXnc8KH72/6iLdu2aK5kLeJeBbSxkQOnVUMA5P3t95YYpf9P5j5xlVStu
KpyxoJ7qwcaNlsRu9PZuVx+9xZsQTNptZnN5fUd2B44emUOMfeyUSNE2VX9tgpHB
H1psLOB7SDEguQ4kMuvk37Y/0nPXgfmVeLHMHRK+BrFToj/NiSbBV1yLnCaUNBfE
TlH4PtresPPKKRcfdYs2UEQ3OLcfS1D8CI7JdF/NYZhbeVWj/ijFCk3wAifnYQ3V
QUgmwHVMy7QJ7Oo519GDLxvDXwpVPnBOw0OBswEIf95Sm6cJz1uIzTsExvsXe0MA
v7dROVGfYBDjcuSq7hJo9rNDEUe575QJQSU1hNxvLSVx8FH9Sy4Uz5bufZ7kUaNu
ClO5JFnEfmYJgmfaEgwH8h48rhFn4ZkG0V8lZ6/DcFjZavS25JMaANAUxKds4egO
gHQf86n6gfdziHGAZCMp8Z5IZgGCmG52KUNX6QeVy0JjYGdE71Aa9bq1KDLTYZW2
Cd7R3doZomf7JKOY+sLivkO6HU26bS+QF2PAfuDud8WngkIXiAB2/D6vFi19fJ8t
6E6x5R3TseUy9cWAp2oeoNpW2bJRYGY0Ivr0Uf+URx5I/wOtdPz1rC+g6mmn3iT2
TrQ5U2CLS8j9L/6WxKluPBvYG7zKqlSp7eCjl9xmjm6eGS8W68IqvOXeVpvoFZLs
oxYjqok/b1USPq6CmaF2iJ2Zk6Px8dwoJdcyb7iqHi2zKpU6U48WMSPgwYYqzaNG
Edzr9Nk8B4PaWwNqof7KlHBc7dCBQzO4jkO0vWKxs8VhwZSVQgmcQyylHdMVIVHR
11heG2x5Yz7oGC++Nv79jBqFfI7UCeTaM6iEQFYhZa+9BSZKbwiYIxnCdBELhNak
qmeug96MpekvRwnJtB2136mtO3SbNQzX2D/IJ6zpt1VQCVIQcHuFJvRiMkT/c20m
ZruJgIJhBwefJs0UBhAFpy2L/BCQowJSQjGO4QrUGw/6CnfmkAsoKmLe+UBCvARG
dzpg9hLyZDBL+7Jepwc6LMhMJAMlspph/eWlWh4XriU+mnLlQpEytmvC4m03SdIY
6R7d5ih3gk0tj3LclaQJZTM5fJx35I2EfRFU0UkewTx5P9Sdn0eXCeOsaOeewW/E
ZvAk/8zWOl0WXiAbOknKGxlRzcEt0Z4zZpLFQFlbavtuADovuZvjFWI9DCTEj4tM
qdPNRQVnf7guO996cJwmYZzZpnx3W6rGoReXNsuG/G/oZAhj4eBojoRH5Hfkwk88
UuuifwkPgmxEHQb0qZ7aWMDDaCbrZnMruBeByQ7PpiUsegsHy8NOZX9Rb7KjEPY4
JVfkWT7LElVzIoPVz6IZ7ps00HJ8Y5DQ6tTZpq7cS+SrrKLrnMkQqQXlTY3E8on3
K9Sw41hbuMn+fS1pOeR91bxIQlsB6kzaPr0vq+r5rvBVjq0QesIw+Hho3GW4FvWQ
Or0B3J5RsPIc1vDDlxkoL0Cvd0hCwYFnT7Q7N9QyXUV+I2bVWGqheKFofEOPKytR
u8/t4+TqPmTXYIgwQdIpGhpf26yZz00gPnTV/3aL+J01rKgKMXRNx8lmu9WyOyR0
hMnY/0wTSMntv4CT2MAYoU7wEjXicgpOw5j1yVj3CFqw3Np2GFmTngDj03lqLt79
dw/InZkDA5WmCH+1JJvQUs/vSTcSfl72hfg8leUo7pXDhZR1myS/3PoW0zjJIaSp
R2RcMpBa5er7U0xGpMH0IRbL6dMeHQHY0Nys7UaXK9n7ykgCNOSj4ehijm7LP6Bg
ucG6+CL05C5e9IQwcbZ902fKayzYtbzXsZkfVReGlLi258d4l5wLJkAWGkDAIC8F
LAjzcFCz/CKHY1CatYUiQY+PgIvF/zFBj3DMel9rrz7/f+LW4y/lqkPmrxacxfty
t5jFu7avKTV71INDaUXji4OhW3y2GzuuG1CQ+W3T2VpB1HOrIe0oEJ6ZU1n8AO07
Lo4iYreprASrBjPKPsf80/Y4w+X3I7dfYSp93y9f+f9CiDiSSmEHtaafgvJRAzmY
Z5brjvOKcWrc/4AD3Gqr/dLrY8zt90Gm/clj8BSJZdXyMF4n4sRyVAVNM7V5Tzro
DrrLtsBTZbohC5XkEhJ5rjmYZIsyiDdJUHQZBC9x0NsxuOOrF7g2U+Yw9n/NBsxi
qfQ/BA3jtleXLXADR92NIdaiF4RF1ZI5uBx3NXIXb3LNxwc4ASDMkbqfDS4CuEdv
6lPCkXt8fyXZ0oPUcdTQ6ZjK5Hl7Aca/x/BLVlkuQCIWOnJ5hj+uMTc1+tq6hniG
hIgvm+vEyhhO70P9GSBbbJpMGzDDPHaGU/DOihRJqWaRZnGjWIQAsLHYPDWXluqU
wCu/KY3X7kxmqOMSFCnf8BxFTA9vUKopgv7Bm/njO0K3pq0XXJUY7s6bkOG7MYVv
g+5ErMYfZvmx2B/F3f76HmRlu8QY5ZR11AK/yaH7iHqvjQLxRqCztENQsqww3bfm
ePmdLXvKz7NGoOuqaYKccW/twMENtEA+jihrV4Oc0Q+iIsq4wGhFsCni7YUsSnlc
n/FpHfl/+SmpVdlT2vE/zxuAAr+8dpE08p+mTnnqSYkZqOw3OcOVfXpVwEAhqOKQ
MsJT73/hHJP6Ro8hqOEnJa4ZZSE6UctUdoMhjOIrn5WzoPmMASQUhn6+c19txkwP
kt9nf8ABIdYPBDgs6moat1huaBDH8Mp3B5mhP6xa2fIttGzv6EmjYQd6SHuffAHN
fMUz8KXiajaGthgxLnljlRqwBJpHceku9HFxcF+VKWUTYUS6QU9ddMpAJTlDfWe5
ihqCKG4Hrm0LTor5GuwmlWLH391elRrGrfZ87WvEzbZnCh69IboYCofTuL4NKfyX
0ii+iOafMHtrFHrJhLyVLGIvLxV3JOfGMfx1DaXFMYyMAyDD4QJRwxbFJ2p9tgoe
6J3BNFdr6jAahLKKMNiUzHrB8AGO2eypbDbO9PQ2+MuH9oiQRFCy3S7EzcDvrdRf
fgSceAxJkcUc/aVwPWRbXmp0dBpxhqzxn4UwduVRo6DuFHgHXc97ADU5Sr8/9BLR
K7UBJ4EOvh42QP8CrkuW9sIObSFHrIJbmpJ7gazjXhOngBi3hwy+w62GKSXYpRAj
IcTmlXTDBwG22nsq6SreOUFsYBCnoKmN5IrbRJsmYO6Jaenb1tFMfTZzqgoY08si
CWw263oI9xPRmj6EMS+gHfVGvLEZ41smYiuaSgHgsXazC6U7SVJMg1SEeNUjTsxW
of9AKROhkYUYGZ4NDzL7xnipuWqHy2YxnLZ67EYeokOjIg8r+kB1Uo3tkwhbHynV
YEzclyj/cIBR+//3p06XUmQ4CeFLx56kiP6G8RNIoCWCkSVd4VO9fi4mzW0M3cIa
FbOdvt/cwpC8aihV+4iqRZGRBvR1N7hqf3gJtdikJX/rQWx6FAgJaDqR14m/mors
9pjhs1Lcfa44HfxDGiDkB/CgCT6fPalM1e/pT19izExHYRR8d3ubNaRacBW67BuQ
BOi5G/O8nTCZsOfizwEZ3K3RY39QOav0tEbyo17dceBC1nJfVpa3ffswiuEZpnh4
dfYhAFBjLb0COMux6383p4ZwoNKk4fMKROHRoe4nYURDER5GQjFd/yvpwZNw7FMT
T//uR3o87GAiUXuIAfYuQx7TvJQeCUH0HgDAsiFUUaw55Jn5RZ/EbkjfiqlE4TVv
HH1vRwSN+12vv+njLU57RlYDJ/uSc4+SYrUzZracHC0kbLD6AO9s1pqa8Ldv+6jH
o+1u1zJBLA8GWtP3NUQZVffhj7fHjj1oQh5OwYvFbZMgMkx5FLvgkSlQm2Qif1aU
TPboIAWTumR3oryepa6eEN2rthpCDmU4qLyn2vpTnqWDtDPMV7uRPOeXDZ5eMOKP
u92qs+rR3V2oDgfqJyP/tBLA3gZCTTAjGDev5a8A00M64DLa9ZL17RUmvv7j8Zg3
xYJsF5sDS9D/ePWQAx6iYxQVrubqZ5NJ7VaoaXnxZniDFlP3QW/flP3zl6/NoWOO
BrRIBSeui/1TPigvu68hOGI3d+LkJcUJEhQpUZ9dSG6BOQ78N+nz1NMHqluVLOR7
A/XSRtq0tEchwU05w9hfsV+YfCX6WH/ZugTDYZoUmpGY5U45teUhmwr1nzJWYLKv
um+9UIFQgeTu4sH5Bm0fq4oh/AIjl5wJTn1VuSLgm9zhGofagQylBz7ER0OmZX5Y
qMI0Zc8BzN9+iIQh/haRXxOVPhWLGpoxKhKaFkRQvd2A9665Wuf1Pd7vruRkiWHs
05v+ljJDQxg1VldEBETMmQTfPMuzpD1GlJO4kuaDv6sfgfnsN8ZZDoFxsLd2GSx1
CaIDZko5CB7h045RYFyNcIHMiDWhSM0XjbQibDkN1NGvrAB0/eReNQfqWOJ8sELx
Hxi39rEASNs42OL5tLnZLVNtuD0QLsyGneoMSAmxsKtYkP19gWchBlcXXGJ7S6MI
bZoMCOdz4TMWnemD5/Et5/6A4+OGfQjH4bFCXA6WvTign4UVTnD0UhBvvQLfUGDA
vfXpGjFsgrMZWutotN9xNSC34gIVUfTprOREZ38spT6LB89mVUvJ0qTXUvJC+ENQ
HB7MHTmWBXW88B+pRM6tqfDLjZyXUfv8chFQTVJP3oexLY8R48LMpOb95NLHioCm
eWpdiAnQaVkdd7eJwISCZXQEmGW82VQy/eomrqciiRR+6GBev+KlVxSQSLtZoVm5
vLcpUIx/BWOlQPbVJtx+sO22873tys1mcnTpnGXU/p1DhHWliznJpL4dC4/MJOz6
yuRpc1Mdr6ysP6otcc24/C0LsgTsusgtufrdOzNh7Y6ao8McqsQef/5vbA9tQiag
4kcks08XRevB7ssJyQsvD8ElEvajy8rQ9ub+QGw4FymvGoUn1r+dtHsOOejz6sgw
YZCvLxqGfKedApfejv7hisI4vP9J8AYmtvz99Cu4bb3RI4NkT+d+RN2KfsMwno39
vZxLP3AIbZz/tM7t6DC1/axZYzyfomjsUMH8gR79LMvSHq3yP9Ud/g3yrAtSRb1J
cCNcWqkd0qwryqX5JfVSkvRCb2ew5DB+97Tkfijq0Tt3cfGTaJNdWWO/o6na16pi
Psf8nLVcAjSZOxMRMup7sCEFgzDtltsvJAUZP/+eg9bRZb3A6T2ryIvjApMmh1xc
Hs3VPIG6f5MkRqN+2GxsLz6v/Mpvjvi80Y0gHIXBE3HJcPktNCgsvHXUtquL5Q4D
aC6zLt+vXoDB1QDHoGiUE1ScbuOaz9P36r556gMTglvuKR1VLvuyEDSnhK/z4GJO
YFUhmEK8+83XQGroM+NLmSZpG3K22RWPG5pZFrSweR1gtBlpfj+6LOTQ4XLLbjnQ
kbduK4e4ub+ue+KfAc/KretkCXKYJSc0Y4VBARTvpdOO0wSGuW+5swNqkLoPcbz1
mZgBdjrkmN7JrHYPeDDpZOPhaNrunhHlhS1syh+m+dn3ZnBNVBPb8zTROv804BZ5
9fFni6LSn7/f56L6tyyPqoPr04UGp30BEHudPnnQ9tJwD08WKfrYTfyZUVAvHgfA
UiaDZPwTUMH7h/nenaZtLAOVA/US5LIuaauWjENW+gNbO7GBFWKfd/Yc44X3zpi7
lrhmF1DmodlYv6C7voq/8Ou4xK4x0HgZt57gcvh3ikTYahB/qafNTDNtQByvZYw3
7JqECVAHx7zWgrTrTmVDbQuydeAAEcQbKRzlwaWKF0xZQ2Hl4FSf3gvVYvHLTPaM
6TXEPKAn8rUsLurr6vgIg3O3a33ux1bi86h3i0EXXJrSi055vnCDtAwzmn5qlKOm
HMDH4fRsbjaxGxCbpBAZYUNPYAdjNOhPGI3I07xi6h5QpJoW5q3YIDZM2hFEAA9u
5spa82qRWg0GNTvwEWoKgy/BlCFP9kZloOCZzlzvzygXwzqn+N34ebVJ1mRODERY
RYx8CDrnhoCrT2psR97rCfQlPGfmceSBifSCLvM1jW9PStCPbB7/ZnbEfNx/DBw4
t9TI86sg5PZDtgkwZbt4mowaybZHyyUnSL6LRp4fWtJiqk2CP2AUwBZPuQug/Kpa
OlYgxh/9EERTURQ/U3NoEz+ZdOFK4cfx0s0l2nN+EfvfA16vRhGz/WKHIpCPPxRZ
xrudcheGMVwoethNvW1bJHNUi/bhsLl/GDVw8Vm+uWYuWpBuFkw7SusE5NBQrFiO
FFtNrcKSeHM1D8jSUuXrTZiGnrQmqcSWRNNt9uGxiQ06QqMAp6GnfkvOBQ5F4/r1
VgxRPEOJqy35xlXrmO2O4LXONtJGT9MFYkNxXZ+W12e/KEpaNUANxVSXchhkaFzL
I2Vvg2hzbsJ10RrItGrxfcDeGIbXvy6NQoXRVDP2x+w2V7A/Rd6zbYJB0pbwakzl
gcM2Wkyi9euGDho1/s3pTZk1tbcJI0PuCVaR07JxVO17+SArT9koSnC+SH/9ikqp
e2lk8gV8k2rDveXOh60APxlCkKkx3b0tcJX4PLKXm8ofbCeWIvcc+RA8LaS4CWEc
uNpAQZsVh+ZqiJDuiQXL246DF4zNcs05QHtYxNocculZYshzduHmN3COsF6dfpE7
9ZbiOPy6prFdaACK+GKCDJsu/NfFwoBqglH6G0y4407h65HIcGOMkqBjKHc9gEv8
fRS4WGnNl6GjlO7zO/DW2xrxPEY/wqKFqxES8xbYvqmVZ1Dd6GGKV7QVMfT57szq
AjDjmmuBTOuQRiiB3NS4JGaZBXAj2WuvuX/98YubUt7Wkw3B7mxVeduXCU5BsykN
JjgpC+yIBFWfvZCkh0nT/CTr1+E3nY534Yr9jSBYyPfPtr98k0YWTdFbcVRrRrRs
XRe2VIldylmei1t9fCIGuK1w1a173vl8Lv6QxQeTPMKQ2mcuUxXhtKOYq3oIxZ5a
/UvTpNVEQru692TtLnNwE8WFNmV1Fr8Y36fgvSMlXJFwgHqq5dl2UGyMQIor1+Gt
BjG7JelNbod96Ua7zVBm1xUKJl0uymjlboFwNpJaNHtE5jXtei0ebqX2PC12fInE
XTOzuL+PU1D+Kn6+P9j36DcN5jhYKE5WZ7h3zWpcz+SA6UDQ89sPEFnl7TanfIrn
77E2n9iZpNflYmwGFZkaRj6ZT4GvZmZFAPzKZaFGegmf402Zf49A7NpefkHZGOn/
Fylv9OPlx/S6ATkITKNAfVBFLjxCVMTjCeyFjuQxkvv0kI3FILVcTzouDnEJWBbp
/n/9h9HPeSROf5zHIrWrvsm8R2BSsDH0CFgy3/HHXlHSQLkvF+nP7FYIaHf01Sr5
e8YKqyMxLp8Nnl4KduzLAgwKaBJfsf8rAHfn1GI3LHPxAM+B+HUlm2egVIH0OQZR
W8SO2sCjVajXuV7Al/ma24SKiL3hB+vasW4LHxSYlQ45iOl87e8B1nqfz9deWHoA
0p45UasFHlIba4ie6t6QiPpgIXBwItcqODLyNWaLcWr8yry6fDLGUIDWWmRNRNVY
sFVS3aN/jYhzIXzejza9Vtt7aH/GwT+2DR7p0BbK/Gq52JLtoO4fbW4qeTobIxff
TDBlfAakwcKeXy00Q2RoAeJNIExnO6LG65lVMN7n9+rcsTgGI1AzZRk6FuLLWm5g
nNuUAH5l6wkJOOh7/9wksSvy35FSoT2HZq9x09hPXyxeTAFtV9K5WqxtYXAJY3Af
YrRqdeV13czqvC8MH6CcuWupljNbjKFU6awugKDVUMmzQCaiM92FU2PJ1IGJWnue
j83gLSpJPMuYmx/Q1uFTPT5Fpr8VSNcKjv4Xg/oAo5m1xiAJRy1RPcDWzRJTOXaq
UgrkCIQaM8UslWlMGWKhAFzHNUwvfdqAKTDF5WBjsU1m9PfiUrxHTH1shugv6gaV
f2FtyWd+akACmRVr6kmK8BBFk0XwBvSsJS2StFrzcEz+ChT2UgRDAoKBIffJtCyj
2EJ4SiPG7yugXfQZQnpocMoDD3d6VsMXkZqtQ4aECZ2uxba1mExliT0vyoXWdKkv
8TUIZfCFCq7o0QTj8DXpF2pUk7ryfWcy0oGnYDMnUDqLnvQXt91+uMkhalsz1ZqG
75TFwACBsgYWFPmCGHUCNf0JHiajSu8wjxln/gmNRE6sQKN/yfQ11n6vc+lAd6uP
6gJamB2b2HZDJHFyCLa084QdN23eyIES+Itha40xs1Bsa8f9/GURXHobuR5sw64A
iKZJOftNxolzgkFffjWbUXlXkGDnHFux4/pDlmZON6zVrM3cXfM/UiLn42wlqPnh
PMbywzwEHFxAzmiOeSRo5wvIy3fcE26NnY07awwRHRhroDmPOSLuS4NMt53udnMT
wOua/8YLhFB8C6FUt6aWEUHutcAnm+kVNEqN9L3sXT1afvkrOHSUxpNgdtItCyu3
PPpLn7gNDZMNUtDnHJRE+YgHTT+gZnTCcC1XzUomo1bvMqK8eHXdLh3ZVvi3YOhJ
/HSh1NaJZA90KGtYUEYUw5K30QiKHDGKuhMgQBiPbF4BJIdO1DjMpIfgq/SFuSkS
DXdWSyDRWl/60YzN4dq3ytvrzJ3Zc2pBwgx42o7szXGobN1ACV4x/mJ1va/iq8BV
5mQisdPJT1HauseMgFSXRXlypqNq4K/+kaWdc0WBVKXjF5XXCNBYXwyezxO0Hydf
ib9Vi1U8S61GLXbgOV1E2AQ99OsxBkJC3qAlgjZoZFB8f5xuwXlHQps7f/B/j0po
l2OhN9JyPYJXJBTaTeoZbc2wlsk3KI7vuO+CNtGc1g5580H9NvTsCaOp7iwx3LZ5
+DjgXlRAxEhmIpM24QNoVIBDT3BbLezNrnkd1CQlau1OgVVT/w2yX+U+QC8CwFwv
BiCPZgciOcMx4qpKl3Fi7nAn6BjEh6Csmr9Rl+/t40sxwJmEUlycNa+xxecxxWbW
wPXwBRUuKUNVYL9bCGBmoNIRmsf3k7U86J3cCKoVSlubRrjbOT8Pj6MNB53QRTxU
31rO0FHazKcQEsbZJ4UtX7c55/s9ieMKz9skEqLEl7dXpt0nv/FNVnnHGYMFVe7C
o0RSwWYqgGjo1axs4QgPIlXNc7kQEoMoYdxNYW5NaQzvGTGIoBS7c6s4vhhI9zES
MQWS5E/9W7zH8n+vCWphI8weS+TM/mgzXbH1nHInd+Cvvyp1PlK/BL8JSakMh8HA
mL87XF4/89sEB60EubqNc3RIal6WchQF0xt/c5VqLf+TvasLMNo5n/cpUX6LjHta
6gKPdpJxm6kxWVPs1c1keO6pL06IwtQ6xt6OrOos8jXKIZtEwv7vaZgyiMwpX3hx
jvlfhWyYrr/vuXc4NuHXzaTKkhvRHns2aujFrnzRPLT37HdT5+MjghQ0IKuQDQhz
24WaGD6UPqtVuO1z+TXgpg1Ik0rd2ohosudhSnvIL9+il3/Wo/OAsYR4SHqQjJlF
GeNJi5KJyPRKNuci3PilBlpCGSiFBelWamyTj1LYeluu8pcMBbGO7vZBmJo4ZMeS
IBCoIS1gKJ3CHkJSzamgEKErg08Ujhx8HWS6jEZghBY5M0h+eLXDrIusormzaSTH
noIwR+qm3lqof1fUUlNd+Y+ck75u968jW+mB9NAd+XdzYZEo5ATLTGxhEjnJuFXN
1QSUjdR7BjK4rFrgzjumexsJtyJ5G3HxbhntWXYFSb5jfkNeHJnzItNa/eJjeoMz
fSRPnBFMNNHt5UHlcqJGU5CPryHm0UJoOag4jH++BTqcFbThcHSBFSnY5X/0gbmp
D4hy9+oG63gmMy02yVVzXH5ShAOC4iPA+1rp7yEKf4GWhyp7sFpBFOxJceDgQ3XV
ZVqGjY5S2e4mqJK21OXmik6aQJXWsRJAd4P5WuppAz9G8X41pU3WBK67RvIlotbe
RiokmRy6CG2bgHy5PtJ4f68RoiKawg61U+umcebCJUZucqldXssCipgFYKV5lnXE
VxPWbNDzDyPS5g+3+cVOezSsAGJ6/Sop4+yWwHyzKli5GVHj9uxA2xhaLs75bMht
rZYAxGbuxx8K8Pc7m3TU4QOrUt7cvHFkUUhBY5i97oqk7lz853N7b+m3emXpaTky
0+g2NFzlyajcG3FH4dTWnVZy8AJvlW4yxBVY2vKqfeztY6zU5uVs0vY4T9EPDo8h
qI9hi01/NtRQwfk0YLEMUWcqEMdI2PaUMFVwUxdwqjmQaVugcYLuD+6OP+j3lzDq
VFmlkIWQECffJIaXE0YhEWiZ9cHchrQKbXKRbq78LNscepbCnCyOAaHyvm1iWPwL
58a7AOBgXxVxXcGJwux5nJpbYCq5jcbxP/2vF0zb9WOCfTFKs40tull9z4nTA/sy
v58xIxshf+CmwTwDZlSrJ7Rhcgui1M/WWGSm1oJPhZQxSta7eu94Yj5EzGJUQjJI
SPKuNbRb6txe8ZINnWEK4Tp5c++OPhFHGRMd6XPnQwxUZZ7eZkZoiTxpz0LF+Ljk
gA2enhW5KUPwr3QyhT49lv9xSbg/zBQGV2UDHA+kt3YRe79TuyUi4dKtJrNU3L0A
h+QjkETcgSuqEgoZq5VTsLzZzx+qoNJ4fBdb80JzTHpWXTLycVJffRobHqAseC7S
1/APuUo36IDqOetiT7HArQgsSUwsmpb0Qqeb5bNlqJXyUzbqRmIpHs4W3uMNGkSW
+vFSTZI/JfXcgz9PUXOKErLNl5R3naWedhuvjfxACuodIkvjCh//yhyFNABiN4kc
rQH2oe0yNZjGHgbbDa0UehuGNsj+iYLoZ6JJdQEn7V6a/VHoyYxgnoINX44NiJsG
boKSLLDgLWZ3I0hSGrbfQKC6idnM1JTU2boAT94+axfVDp5zKCktcgldefy5k1Kf
Hciim9O+Prn6wQIGeRfpf8wLCTNIKFYZzX7nHzYt7x0tqszUj6DXtIO2jW9kkxPg
fNCeLwwQ8ZAkZXNjMjk8hFJxReohtAtHXfAn/qxMb0WCMKBMHtKeyq0Cg5jvVfUG
m0BwzszB0U9xzQYDtyqoUKfTqsJjR6PgcYRpkALN69Ti+pWCmhuTaDxIB/jhfuNF
E71ZzUv3wSy86qCzIyM+ywoDAAlzOsmSnnbiMD+ncCUWhYQ3yjcVvxEK9nniHjto
S94Y5w5vpDvYGI4uKNUt8x3PKYXtcP2tObiEZXne+caWt9xKAYO8T0lveXPuWgfi
AKjZD/GwOZ7E/o2/SJGpP6luy+BY/8u6FFav04vgGc45hHvy91UhqjwSZ9aqscpd
uMQiMtaq4Qj+daG31drVJkcW/P5L9hi3Iev8DT5wwrGRkcFXvoYSMZoWoGLNyYC9
NNuYbqKO3fhbfxxwiz0zp4Pw4n9zfmVgdx3wlAd0guDyYsPocbAHPDXQy3KCvlkp
/QmbianoOugC7At0oikJO8C/qXI4djekaGzXDTM4AHYee2OWz5gSxEUxF+nlsQHy
jtKJtABHobWfVFvOWWlug/j9cKbJR8Vr+PBcnGrFUe/Q16XDWofXcQxXH7lv7QLu
yRWyhjoKovAigwFgl7hVL4csHdHr4miazo01Jnz2BP0U1bzioXp8HyBJz8Y06Y/r
GzpPY3YsiJj1EQqxVcUjTAHpBWCdpeEtp6D89ctPtnWl0bxXgalh/EVGDDq8QbFP
UGtgtADA68Tjo/FwiUCTlbwK/j6dj6a2xxqEy0R1gPezZSzi1Mgon3gynxvAMSJz
y9VqAqFtoozu3cPyece6bBWjf/EolfvNxPgcXf9O5WTTodkRitL/P5/RdyxCEGK1
3J5/LySf6EMOF/3bHVhLxJPakPApmSmVZ5KTZEYVsfjfU5eOtFHI1Ix4VOd3jUDC
pgip8i+hyGKYMtLPGyOIX2MjjrsCsJ0C2NZ/Wf/KB84f33m0ISH7T0/YPm7Kl3GX
F3VwsxzqjLEi17fjU3GlVskSlnpG0BX8+uh5kplIu5YjrYHOVaSqNNBYcKPkQRdI
GE+0RTFB/RIiij+efzQl55xFdNTkohTuNHcV3pRDA7Lm0HznZ14ZWk8ghh+lB1W6
TxejCU9xClevWAiOzgLVLSCVCEa6CE9pa0/4uryyXrbvSeuBdD1oClR1waOJ0/pk
eXVWpeaEgaQqOwExHYCXyNe4mY5wS6dGofc9eEWgneZQbekfZlvunUaOWgND4IB7
tB30H0QgaT4DuAHR2es1GfOwtD40JI1HsiTdmAiAzyPS72Rqy8vpnALa01nRzm5E
N5LSjfYNW4gXnMfYDPogpcGPOXxbRx+H4fIOL6qdB0s1yU7vS1WPEuckndjTcsvX
W9/WX7nsmqf3+3JJMQlCL59OWYaK0rPirOfB7wRqvVd5CrJ7YeN/1AojIncBg63R
p/o1Qhu56yuT72f12wb/EyrdKhIy2NZcgfuT7vzClXUX1+qNXWPwhX3EoSAWUY8S
iruVcL8cIv1Btpi4OIpXAHN/CTk/7f7yaxPD5uqz7n+uuOLs82/XFlKxH9Jh5naj
2M6IQZ13QyS77PbOB5M6aO+GUW9yzomIbyzXahk8Eb1j73h5bpH3A5Xltd1dxZRx
vRBThejFWIM8/MkU8F+LHwnWS5SdQySyxldEMDYc4zngF5toQ0gpFGPv6cuUitrs
p+/vi80Rdaq3Ltbh7n5xMttq89ShfnlW1ufCccQTKcRXwoBAOSg936+V14mJmixb
lrHdmxn8fgNh+TFkQ7NK5o2jpOjn1UehdNtLK7YkjT0Ji9aYRMij2gU8amYW/pOx
v2T5s7gMY5oZu7PgKCPnZ9eHdSj/8+dA8XggowBRdQnbkDeuOVo90em/K9RKB5Xd
mE7jpCMpE8Ul7Dgcx9V90LIWTzwxKWXt1Lt+LBFOsD/q8MBY1o90peBOBor6gG4L
mpN452UmWV0gl4sCzPwiw/em1ree9aeAKv6Kkl/hnutjMpQ7Wao1eeueS7v+IUlU
+C3LAy9S9+juKspwMa0Q68ormsa03fcUkcIdO/xgzLh2pad+QZK3ILYrlU9/5yZj
QjPW7LxiQ0HPRlR1Dh890Fh623IGOxLgJW7C4TevOmf8Tx3o6g8Tg2ygocKQG0JW
a/VXKezxnGs2dXRVuLlOUSG2CTKdzR4EoG2s//h333OKM0IpDfu4HCx+deD67R8x
w/xQHpOmfZu96uqCzYfEVDHthrwY8s7ISodeij1GxHalWSYu9Y0wiJw8VGcvWXF7
YcxijLmTaMibh2Rt18iweRibUvrW713q+bXndmFlFJUagk/Qgmy3MSDoMg59pLCG
e9toWBIfbx8u9ehMEH4VLZtdBs2gcb73LXzQXddwcf0VIobsWojowQLzohMOZZcG
9dpSa8g/QpWqkWGxg/bj7BcyxVlMCxY33M0KVpT8uNjX2ZL5Jgb50lGj82rBy7y+
ChxON0qBUQRz/j97iKrQGMlgoCsCukcfKtDK0A47apJVo6ZC4ZWBC6cau+nhNHuO
g85hMnv6ZkdC/o9+LRi+PcAOEDT3BH0DnuESBcts74KYmZN6uMEHcN8oWuiEgUAR
HAnEVf1JdrH4narOWIrE0IFFfMHGLI3cFPmPII8WFafDbyxTDBw/reYfx6ukuUe4
VZdOB0N69YG1/XcAiyjpf9jkPD/nbZt4BnRtIKkqNQ1EXNLphTAq4VDeQCDUvQ3H
7O2cl7IiopGMKFp9u9PQkh0q4bApR+QME3xEMMnJWDiAbq7IAzlKyXSJ36IaDdkI
+ijoZI+K31owWudYUItWGpJtHkkpoI8xV+8sf3zH0wCoaBmjBiwmD0lqiAEH7dVr
t/5OYHo5mruPvbZ/oKDugGEObycC+rS9MHLIS6IFtRLjvmUK9sQ/2FDPPuPLDRLt
STFo0y7ijhkj22LTGCNwvxaffY0IITF+RjMLWRyE5mW2+N1PXKKFbLRw/xpshmnY
6Z9uHFB/VCVKZbFch+E/02pbdeQI2oZ3zHnIEhsO+6MMqdWTYHP0iYsLPDvmVzw9
c5YDM2+7uOg5HEeYbVDvek4zFrwPIicWYbzMudqLTsAw0xYIcSOFHOwp9YXoWkUp
XZj6uuKHETJBpnKFfhL+ThSmpDiy3MCAfSJpZF6kCz1ql028GfO7cnLtxzRmX3F1
7Qof3EvPv9ozKrDukBUnHn9dUevMPnMZ+EJeV0shECGewEGdyAmeTtXbuG/VcP34
JMS2L4iU7F7+6VQYafQv4GXqFNY50wlleUZTS+WjHShJCZw0QR/lCDYWU2Jc4P5m
VNAduDw0T3yUyD1X3cxOjGlumiEzd9uwbXZyFm6XlZLsujlk7YYHWmrRpy1Qv76K
FlP9DHYXCv3RnNJsmW7fCRs73jYaKYOnpZAyg8Xl9FlNdSLHB93w4OK3DWdh7fUl
1QDwvhrG7EgCA/7YE7lPvNuizTefESA8eUOiQ6k2uVRH3EYwgrKj+WStJKk9ZBM+
CygnLuUu3ZDWyQpjMz0Qb8YusPIDpuUNxgtkakNsYUA0Xvf68Fb3RA0Fv8OIeY9B
cZJjJRgXZFNGKRq4gbYkCc+UUExH4dUzqAFINA3h0rVJQbJqrlswiG2d4BoV/u7n
dEep2l0/F4/JTIzmSMu37oyPHUVrR8VQoIrbpvCfrvpGbcBV5EVnATUB/SrtECQr
lYvrJVGMuyBmFLZgXC0op4aQ09h3u6I+ccQ1mEVvKAKoPpbeYTKdPcKJNDQr5EnK
840/Ef2q3l3NzO1LpjER9KLPdrEGMbe26ZYlRLyGWW93VurVfo12F3Sic0+nYzNp
YbaBCHOdDbqzqsHY/rsIMqqL76xuhTI/z2JKMV4Mt6JfsvgXiyuLw83/KJ8il2Y2
Xaar9ILJ4t3XD/s4ZomIrA/CPKzqT0U2Gw99OAGCu/T+Eli1HF5zN9ki2xqRYS6g
2YxhiugEBYyE0UtgY1XrxanDaY4UWpGvbFsbWtW2f/fJCWvSATDiARRENT6nN4Sj
5iqRee4Xm9ViUN9EhzdhTgzhFd0m/SICJgIc1qJme75brLSocR6lb0A2OfNJREB3
KvIOXSwl4o+VEhpMB5pBdErbZg6ZfA/3vzZuMH9xhWKXd0yHv5GmvHrcE5gv4mYM
h3mKMIhALZGW3xxAFWEUjG7LeGyTK9/wV1uC2JDaDGj9gJ4QHA4jzG5g90FMz2Ta
OvIBLYDpoI0j2ek4msQnE+BRc4286DF4CK88AI6oAgloWRGYTgTcUicxe5UCI7/m
6D0J6gPYPlzoH8/OTMvUV/qMNhDK5BwJq/xA4vbPY/yKJHjZ4Xju6T98JPAOMwNP
29mvBRjwWaGc+35tVnaedcaDz+2FWEVkhmjNLNN59gHt4qoA7QLegeR8gLeYRvRf
N/K7jBW7I2NOoRReqvGO0YqGK0omF40+aLjyqbQ5u9CAlkrZhs9W2TsETwfjSrR3
7wE+aF6PPYwXm8qSOfRhw+zbHPFnXiibl3ZuoYzXvrO/x3FEzfakk6BFl2cm6rWB
x7/jE5A/xqllNK0spRkHpwXX3bwLTmrdS/g60TGZbp2pCFo/Za78YEAHAAHC1ZRR
+2grV7hRqmyFOTWHkEiQdcXWulOsKlALT/0F+HN8s5cx+P0L8D/MZNwEf/N1HLnj
mLyo2UBu0wOLqkJ9y66XzkYEFLW1C5BhjKZu0n0i6EFMfyviJEagRpvL2AERIEks
tDmY2vVqzBprqLTQyt2x/qDfjFJExUmkhM/XRjG7/5KEghwAWqZl+ptdSjhU4yxR
QqG0+d7cGSFMQ5w1Gu01pcIEh64UErDjr8l+0n0xSg96fGDdCvpaoJaqhVFpcM9U
MyrzB7wCSQ1QFhw0B+JEmYB4fkirTd1D9pPkzgsAR2E+RaOyXMgIHfxEAugR2uoH
lKthY8oH0P7l5e82kZ/ckbWAlFCdA0LJHuDrqQLww3bKMmiKnKmwbl9hbnkdTwhe
rx9QqgR4YuasGdFo0JItq1lCLJdFCPwo07IaYf/diR0YYO/v2+2wgLvOEecIjEwq
xD0ImXHDvHWD16MrWgL1ZqcjSRf3qWtLq0vi1YOBnWTme62j1EU3EVpLc7OeVkFG
IUUjwpa2vIFNkJhiQNtKTGHe0jZi8GYP/KhtbjbkI4+HcqHgz/5TwclrgfxV08td
7mWC1Fdp+enQWbdzGeuWFwGXv2+GA0c7oCmrIVODRoQUwerhEEF4yIGBB4Sdz3Oz
TO2Apv07f2R7K0YpxMvXwR/E33uwgHbq6rYDxCEahUuiW633iatYywh3Wc82kSvS
gGtj86ISpHd/1h4WGo3oPsDebM+ZYSTvmMnoWP0zKhrFuNi0IABJywMTC6eYc4MF
+0YOIYFkr15bQ6O2/0hTI6aDnhw5UmVdCCI+YJXZq5NOVfTsenCP37EowbTXWAuY
Hh3apXGckuSWAT3FPl5/A4+rZoyLq6Sw4O73W4C4ux+FHdE1Q+6clnihlEEzTcxn
OPNLHhkvt016JLphAHK94iscH1gOZTHWCFRkZAZSAMJGqM8ue2FOD1U0mQV6sjes
FkD5sddvgG9C9plFw9ydxiz2ZRWYvbTaEoxYKy/ESoQtIUaOoFxxq8BPwVkpNbMv
b+aXr2iVdSPLFH3427Jn107kBZ7CqhWmDQ6LMJG1kpAdIcOgiELwon5+rsPIk7pE
UOAy75b7EF7wripoVS576sDhoSFYRHxmdX0Xp+JNMFLu/BjJ4IsAiZhvf35aEhRv
wyMEqSrRuSjDQHPaz73STirFI+xbx/WU9TkqDxKFtKHfRmzl8sKQ/U/I6jAm/L03
yoSgcFbUsMkTOMZhq1JmE5vNKM3+nSpuND2TaA/d1pEej+sWqA2kUPW58BXvYATj
9u9U5sc6rW9QNYTpUXMnXssBfNc8VCDC6mdK1315azAS6Qm4tM3yIm7LuqAZjvU+
wCA40A4Rr4b28/1CwC2TDznYWf5O6PSKNQiwB96UDid9vkEXpdJ5S6PzAGt+C5y4
OCU4K6GatnU9NPh2l+/c0pb4Sc9+JIOUXiQccyksrryo9NQDHbaOXcUpWP6rBw4E
CPfQBc0KRnBV9ItijXmNWSy9+LhlchqEgMCXDzso3u5aan0JL89F3TLARd68r1d6
ZR1ZgJ7CqCU1snf/x7umEuFZC1rkq0bNJPLG1yBassk734Kr+iX4IPYexCtk9qOC
p6+STGDhNHxIro+zo5x8wXi8QlUMYW65U3CKcjJLOTlYkZnmUcieXjLpT+cakNQV
Xn/8yDm/i8CcWxmH1BxfCFBLZCNYqtZVGESLCe8XLnHfQzQpuEQHp+6SoxTSdUsn
JsP16kFsbRUFl2InpuvE08J9g4re1bIHd46OyzhseM/EJaMF+ZnRQfjFaS9yixbU
Pctdc2ERPL9UIsUIuo/FsbTQckdV71eGTRlESTZ7HL6EZ2QollIRH5v7Ub5CuW7E
HZGKHjIClih2FJB6dKJqj4wxYwrZd3wNJwM4fJLm0e6noyRA9nkZED3cxchisUpW
67yZpwueOrNb5pF31t4sE1T2nFgLeL/dRNTPKCa7qy1vkqrVmnZrn1yicVpqh6RD
MN2QMrGirUfub3KFoPHCIYbRbcrGB4R8N+k56TOH/LBPuiLCsBUpnBdegzcTMYDJ
KjdpDXi6RcEdAG79KucpkHl37iKmmbRtkLn5UxJcAsnQ7sb8kcX2RaQCjZhmngDQ
Ja/PrDegxET0eHbaZ7meRhjMbsDTicpBfrNlygGyNMIthrSFp6YV3yazlTgnnwbo
1qUsQLIvp3GWj8pt7USEBEwDs/zTlNAcfRTNCC/JtaWNaEOe2Fl8dRICYgzbj3Q3
kMD/SBods/XGSCbs1e1NgCu4neLZCPZrKseSCV3v0FsNMkaOARSoaq9vhSnqJgt/
fiy4qEN924mr9mZyLHILNmtLEc4lUGSV/B39RAkesJr3AhOq+qy6tXlPF0IgMcvh
ID7BdVvnUe/NTCRgP2V1qR3OORYY/dpesAi6uopt1A0J0/OHvUug/Nq20CpS+Efa
M0JSMFsoj/NFqrRwfUD1jI4EmkvUyi1eZtwY9EP/PKOUvJDsNfVQTBihYEyfjBD2
ssTC1jVRwDOsMXJFnGCijXSGmZm7g7rRnkR9tMANCPhXwH8g9HBm8digDEmTff/9
RdGoXZyyGv4hGbguPXqbnbwX2Dcvpxhos8U6G1L90aOpS6sDqlsFr10mszsILduS
mcljkZgKEb9xXXCxmmA6cblPkUUYrX/tkg5gGS6CrixKpusvLJi6XigRsN0Hkcrz
3u0z3bNbTFDfxqDgAdGv3fwDEXSbgpwQxTnlQS7ntQ0/xgMjYSlwLNMxvqlk3AIl
P8mi6wvfa7OXleWXKMlRQlRIDOW3E6KuiS018ulGf5j+oG/3dO50m0VlpnavqiQs
J6DQJyIXpOmS4kWXfNqzUhgyzWWo+bFPLimuCPqE7wHEdw/Py1PN6ZS9dyXmyfma
rlGKaH0sS2glEfOypQMruT7UkUDXzIjwUn1DTBxubpftWEWjHSCXg+Sukyy6t7aB
yEtpQBllE5DfM8VKCGusHSJkgvqVRxuP8NtF0/tvr/fy4s/biBNF74ZIRBaoc4ZC
nBeDEqXwKKWuWjVUk7TY2DvRD9BCgmHc6jor5mfl6VROFC4Y6Y+8KKm+xgaZziZ2
tsIT1cWZx9VdnPwfX/Qah/ZQZ4spXdnVqRV8bIwkCTRpK0D3Hot8GMXgoP5CBmJm
Vp5OKs6MJAddz2ciTtNZ9THJ//6y9CKHTmVuUdn2bCKrHXxSFga8NYR7UOdOYjD0
YAZACHSsVPYveDntevnem2RFZCZF6QpPGkoTvSj8BaIbiOkntYMW4eNM2aGdlqAZ
FFcO6wtWhvrPUpbUbEgaguej/MHnEtSyUzNDZHcy4VEY480S+UFOWRAC5U/A7lHO
uc4z4puS2cRDsVqDnHsZjnaLnMgCQnXIlNlOEgcMbxgHu2uYzGaES9Tlx0Bcljg7
lUdnOTpX2w1Owc6C5sEUZv2kIqWCUeyti31atRSbiFnBXgSccyZIq/o56oRka42R
vvn1VAg0f0fFOr5wyeGZTyfrb1z2GM/rn+qxTQ+a9A+VqusGXcwSDzI808OIxXkX
r0tTg2QIQ6PjQMQbOs3k5OANipCYVyirJYrFf31mcb632/kiJeYMJ+Yx8xQxf148
JS1shqpXNG4F0+2Dx3a8MGI+lscaTxY8W9gVbMB866nYGXkXd+jx/0EH11a0Rw2D
WAW738mXQlg9eIzjeappk62B8zQg8BNUqu63tz7Dr5FY2xdLAzibFT2Y//Uv1dgG
/axa3n25STCA614/pvh/DH2qVDI4qvYMMKjofpYh13ffbZvZaA+S+kdHNupgYCIF
UeJFA2ACCM25WRW3LaZ2uNF4DNIH2ak8h3ExYNxhf3xtDio/4YE5yrvI1QFKlCkC
kCa/wgm94nTwm+sjO7D7NhMMta5PvVElktBga3Y3LXCP8UKk1i5XHVcajf98Tl9r
HSwxMIvy3YsJpy+GLQCHD48FgAamt06zPKCnesSRtfrrchVQz0h2USk1KAX1Xqyj
mRRZgLdUEWKWjgs7PgRn0ZUc7KfIbwvEPMJjrm41fApF5Th8mfgHhxfJyvI91TlA
6MWoH3+F4JY2IJiY0sgs+0duN343Ee6L6rEV0fta9V2CIEIPL/v65YoJQ37EF6CZ
hH9c0+M2Am9buhzBCCX2R6qyUnsv3VjuUQtrPYu/kJljR3k28BwfTMTXBCPSqRk4
R0wJnAzVhxpz8wup+umMkjlsuEG3SAWR7Pmf+8udP2C69+QFQCLEYTPDmrSDHaFT
xhok2OCNCY8R52ZQIElj4qAUfH3H9tYPP6g6sGWsH/J9bpP7rsoEHmcaNBS5AMzK
SjhJPFeY0ACV+WHlQIbjL212+8K+PH7HJr6F9tAuGWcYbtr/RWv9rh2GdSb1AYLw
VQEAfCMWhAsR/mbLFUf6ofS8gGi7ZgUVQ9QRL8UOapApEsqbDKuV5E8MFqxM0tdy
kRo1PtcZYrmwnOF7BjV/DHHGd6sFl5goG8T2k4wTT4C7rSb6i53PM2wzam4xNCoO
Ph5HLT96bYNBVvbYKDUKl2ID/aVGvetBdZrGeCbV/oUjM5aLCBM5EkLm3G7nkZw+
uJFYkelWF3r0uyViP5FxgKbLSSc60jChvWejcWQlfp680ska/PAPng2n7ztwHY9C
42z/XsPTJ6pAhgb7mLyMtpY0b87HhGIFttNRvwc97iOIyw8rLDiZ7VYnm4umMqMP
3ntN1T2IPYr5RttUw7c/2eQ6ZHB/nP/T+8EImke3VRCoMfCLlgzaPHilobRkyP82
Zs2DwkkM7aKvGwpp45iXOXsEp08RaoKBA8WxACh8a3CNeAyv/rtH5kElMt+R9636
wHg1KpqUw+pG3zgkeuUNFwSorSuFhz7txgXcX1mSdbnZ2bZw/lEKGKeKw+JgZYsc
PlZp50OkVCPim/WUz/vzj9iJ60Z2d/jaHaUXI1Ju6RCUVdU+mdvVLlhqO6b1vijz
wCEmw7LopmSOfAjS4d39JMrTE3U7PQoJVwwLIqlgkQAGewEgO4xV8dJ4Nh4SMWCG
8rYDaoVLYnhatcMA9L1aSma50dkGRWdfzuRF1ZexBSbKS3kRrnBO6KXFUIsTaYQQ
EwqgV5VKitHz1qch9NAKXuGMaqDXcCzwMcfla/U//Fs/KtHqL/Ygu3lXubfRdk0Z
Hix7TfMUsXscBHgv90TaP7Jod9O/oVwFj4K3WU+FqnH9gzdavxFKfdk/TGfw326H
cY/+KRDBX0Sdjiufpjxo65hX69nniNEQFMmQDxSwso1+CqKtns1PCdo/jR73nF5v
gIZhJqFazSq/cHrJtg0zxvRLCbxAjS345MtWJCFkhtnepHeVkv26qOLZLF26jWS4
dI5cV11KKnpD/KwltHaWaxxgKK9lItWgXpqnZLmR2iE0wwBMBKThoSoQO9yiylyX
F1mt3OurNqdR8WzqNj53Lhv9w9psBcnvBTesPhozujFMZagrJLs40mB5oLVwzbS1
RQCLLigzDvBgxqlriHFJT1XvEzwEi6YdGHYbRZs2OsBHMSdqruingHqh6aR648Rx
PFh93NhB61UKpe1vfrefkAjOA84EBMujo/u1cl8/7De1+UAMX9XIuwXb3tgF5j7n
wMOClhaUXbo03vw011ynXPCFWZXhnj3vK/Ahx1+3mM3/iWKVkWzCd6DObv0ZgEi7
ZrMYlArWlzjalGowZlwX+TrBDl+OseT9OHiIRwciEYKhhiTZ8Mm7eraMUhH2iB52
6N2DEAaiBOwunOCWhYLOnqNs2zGfImUeUr67h6R6ApKF3/gvFeHBiizafOgeL4lf
8wafLqrCi2oQbALpHa5DIk9U4cHHX07GUxJ8FwBHcCGbLv5aL814oyX2dcc4whNF
MEN5+n3SlkwoOuZMQz6rSHPHW3DNhYlVc3tgynl6/XcUcAgueaaofraaIEE/4ked
8jRQWZ6cmP3Uu+BfIHZ/SBsx6p4CUwxjJ/ByZwARJ7bBzUVdU4WE6MeT4PYBoQAh
vAMQ0F+pe1BTH7wFh2pl5JnKFK+SzXUQuyGc2KM3QXofDaVOV3VYIxJ3RnZ3fmMp
0mqg0G5VSG1Vf6S4vsQ5Ry0MbHLx89NDiyc/ITcuZoFAuCJPxvuRiCH/Vd0crysE
9DlcFiD17NdPUr/wqnI2AfnMWMKvM6xtTjbS14nN9hdr/vZpJXRIG339nZNCLJMz
LOV4cmcoFql7fKZ9fC0SFCEMnmz5XJBeahdUeOohxIa2afvhftMb2WWSl/8YC+uR
qgCvbg7PFvFspzwUN+FBEWr+Zg7MvHLQ6c7WIE2dsbFxuAtVSQSG+AsU6jATYW2o
63D6Rn/IVUOvfngVpAbg2gTdPmbzKnHhqkpyBaYaU4eDTEsjXIEOKslytytORnld
dZSYEoiBn1D6fR0jMaFrWmkHeZOj8s/kq8DjuncXQpy6hKD7G8x9SCEGxms11CLu
w32C7P7n52Td0iUfAtOXNf37MfDUpFtwjZFhFREbJxcUtK4v8yy31pxk5cyK6Fdj
a8L3eaYKnizjgwqcL1xz6fPQYkGGGnaPphbut6cS0gOs+FyqzI2v+87ABZnM5eED
IDe0XZ2a6aR2f1oksHwVOpynsiYCp9/luT+g82oZqODD6GI8n0fCGm9QLMy//EKv
BDFmrVloNxgHHxZGr8gw7f2GKHp/QcV6fxg6DKRh671A8BnkEYKb5PIWH41SyMxq
Dmh1YaFmdrCFE4Aw18J42Q67rw1Y1xZsRM7SYgrAoiIaL4lCU4uDeRYVoBgsMFMh
d+nE54zVd9VBRtfIt1UsqW2D0ppcPg+4JoHb4JlzA5XumdqD8sbPl1g5Mx02IAKS
4fti3pZLGjkD1qmZUHD73la+9kBfoJ5Pg7dOYWXBtpipHLOZp0sdJRIKLMhn5u7p
xchYowKlWF3CVEK8MPIQHQ8/tIaC9IwVSSnY1EgWBJU9zbN2H/QcZ+BHeFkLn/ze
ONZdM1Kto5afEpOse0jfRPTAlviRmABKKK1iwkAUB87veIneKQWnlVh4eo0dkKci
2LADWtg/NAQS1x8lZIi0kFW/g3x0c58WMmptnfMyNOM6aYT+80X40dbcuiYFt0rH
nefwGdkhYl2Lcws+1OQv+F3QcQNbqI5OTuYuWwlqDqLJZY3Cx2NH7GvhkO+Rj669
ph4i0SeQK0zfdCxGiM1ND99yl1SSPBccmJcZKWpqNf8kVZWYlDK+a3LPsTBFQqtK
QhngtXaDrRBBvJGkTll0x0LNalKBylhJPAa3XDCNve3g3j4OTDEROWUgx9OnP1Hj
2295+C9Ck0t/DJx+UDiMX25HCawwNE/o08w57Es3fZA/10puXrhQXO58GoH5MFmx
FEFKPgT4Dg+SxycbyNH1dVgK8uZZ10MAGS9NVjmgkyE5/4A0NOMxBDkssiZcTw1I
NDlUEjRFbX+SVfxH2CNpvceKsJawdCRLYK/CmG+wbWNkaKsSmOZjMgRmD1HMcqSi
KaO9FyKxUd1f7ZWl0ypw7myQnB5C/132bIGkeO8tR5gFqxUQo0bHrXRA7c2CEvzT
rOf/A9sUYSpgRPQNciUQUkxCaMEOkFQZAX/pCDxZsQg0vr3eFQvEqEtn4APumGVS
vzjzwGblYYawY2TP2Ab7tNeWJZo/h8JZcR5smXdAhPqUeDRf/VX+xYDeOkH5tMKR
DAGDywgT1Pa3rIn/RlTH1E6dhpfZ6BJWnngSHvUWq1jIhnlbHQktPkt+t4UjeOo3
DZpGzeirZLbihypXQPC1qpBOLh4THeN++vVTwUmQoARgUC4j4SFwxFp+VA+1AsAd
2FBPfDkYScD4ydAkoviOZVv7zHSBle0kUG6mmLusII4xvnU4Z9E06IBPNhZr88am
+vtpTo2IQLixuXYRCLd+dC0zSxLPvd9k0ZCx2he92hu+7TDIP9Y5O1KgNWJKPaM8
oNWhsPVrwe5sA9Y21LYfNfMdZ6ccPMaFdvY4SZhiDhcU2tBkkIyqzWNhHCZRN2t/
Yy/TpLcwsUmyuunumBd12ZvQNZZh5RXtVm57RxQHyen5Z927b6bDxj+QizcL4cRk
Uixk7TwZN/MSJ9TRztAeAIxMQemc6g3BRlObpVeLwu7LhgAGD4YtpPHBY7MgHQ+V
1ojlNTw/N/7VpKtTIqog9ka5J7WtwdAIjklgLbnNtNSLrYI3mBQ5DbwQ2R/MgO2g
O1b6kNjb5juPqyvQGM+H7JIiWlb1piY4W04j3sOdqzNyk1ERHUarCqEd+mHKDExa
4HnTsrKNe5f3ny6baFHnofgnk+upZT/LkHuLQgt7cgtsENIlgcybHiDjKOxWZWrh
7uMthyX1FBGclZQjNYB8YiIGX8d7pfKnKdNc1Uan3a7Xc3CO6X9ipm+OHcw9YGYm
qjkCOrscQhSWVSvKLq5PBUwtFEed+isyYKHMG2w/FMENdbAv1z1FVDKsorgzJByL
S7a/Tovp7ghYt0F4AZqV1BuaYot6l2ODxU6Q2NUsAAl3+z0pK32PUxPUq+FW8uTp
i0cj44iW+qKTsGGhkMQtC/sIG+lz/WbNNE/xEIlJ0NvsVhrRK7myE0kZTBV7WePc
qrRCmiH5DV7Wg971kbU9oJ04lrSaw/CrrxPcwAaViT/7TpLePz5pD5wrRKkp++Kg
M3UCeF4gK3HkqJ878ti/LmhMb/uOAVz7P/lje6AtBtONUXOL55fjkw0DlPp8Hety
YxMZKlcg9ctbsp6CUJJpFX422muwCxHxHXg3iLA5zAC1jItVEAMb67K1h1mCsygp
c4bI38kPTlMI93qLzb9EVSWoKh20d+KIybvJvhz1Rgc8L2qC1mfcmxFOJtXxy2mv
XpVxXjJMF6kGDE+DXpuYwTYetN/YM18HrPfDASFOuq50K63QYu1doGmeNPBX82ce
QcHb4xrc4bg5SrSpz5VF0WNBhd/wpxlJssFyDXoMkN6Jzun2FlsmP8aG80UG0sQT
08vzMWBYTMeRHjPRPXy5iPw1Q87bbTN6BwsdqTmTg6ilbJhT44dQc92xFXzCDYR+
+5yG7D3EUXd/ejVfLX7V4KngxNdkhoGZDXyq7X2uAmuaq39j/Hil2MCBnJgICyX8
P5+BJGsQEAx3TELdQm9z0/jQEps3ao/FH4JISYvldo7OWFIUHTCuNWwt7JfNnwf5
Vr6zKPUK79qSDeCLINCpRpqiOXhaPfpcpwP/86vIAHF6VL4v8HFaqiWybGcEemII
8ARcfnPku7SwHI3KrURl+TKSNHygicbUNOkSBadrraWGp+q2Wm1abaY6QVOgmCQh
tnggKqcp22skHjHxz0UHlyPlvQs4ta6S8ZG7A13xeIGgT9RVo3eTbzwLB4/2AlL0
lJHFc1AQNd/+jgvoYio6/T3YeFqTHieZYaZuX5JpX2imYmqRaVZGzpSyVv7p04T4
0wH/tbzou+7f+XNf0k0Vvt4x8qpNzTdmluIBxYcV0j+PNdw81zaSKWwZfMTcLAsy
J8rNAPWBcam78uwzv5iadiKgtYtXZwhRLehz2RWNX2U/3uGlk+G0nj22oujKJsp1
IYjsTAlXvYCvgu2lZsKe35sg8b3vmwDIZPqboQ4EdPzdKBf/ryf4W0MzXYF+JdN0
/PbTYhL5ANaV/TwEXR9CNM+PuUlw5RPKkBKXifeFeURb2eATJratuQoxfDHnIdYp
xvOq2Er/Ngi3AZ1djvznr3amYamAkYtDAjxR75lMICJB6rTtY5UvHPjC6n8AKzSy
6eOHOXXxDxGOo13GJfhl9CbmtIe4FYkKARyciQY0oR9pQnBImsaE5HJww6svxd0y
/pXIiJ5Rr97yn/IcEVyLt/be8UPMRMbaCMVBjgr3iwXDbglEa1J8ws4uTIGfpSOh
yImIJY39i6JEImM7miRVmPVfUfDOke0a+t37ODfVAB3GnNk8qKR9eVslimgXu3ZP
doJJL78YCLw4Cz5TTrabSyu01G0kJVMetlMxUFLiiwpEvcBpqyByB4l0uUUZx/Pe
z2JFs2INFYKLNJsRDiOY8Ora0HZ3wkguRlsvjPZF/wZFYtnjZXtVAKRciWYlMgXU
CCQyHdbd6FzqEQ+vO+s72gwqhLayv/TzFv3U/GqUuXByelQZMb8oFRqPnAZOTE4u
mdRQREDzHmcW1lE17jzgLaH+UbM6ftBdM8GGndYL0TwgWLecxKCMFIsK7G/FVnyr
AjsBdeBoijjT8UqMGrr99KK4Teypg/TmgaBqmU6htGAEc+FGjOAYc9qXTN/FzA46
alwzeZvwbzpieJP7M3DT5IoxhP+iztx2zgltFooQ71bRTsAMoRZ73lPLyKe4Wb5X
+3nFjV0H8unKZ/Jwkq7kyrd0nuXpHaRFWun1EEiJqOZT3UZqBex0ZzGMDDdo/pvu
DYDKR8W8nDPBH1ixjiRpmRkWdaKcoIKfUoHOeRnrvTRhn3NxBr7+FJAD92sdsZbt
n8osu7Duz1uwAZAxwpyFEPZJQfi6JDX1ncEPqWnMvLJ9p8HEwHjzu37nfZ8GRcSf
YcfSjoCz7GdMfL58ghCBcet3SyosNCyPzPt7GfODmohgWSZB22QKr5GrpLr1RUoo
u27eDDfBZtJYWIKyClYpl51fOKkopVH43+HO6rG0VFVKgVdsMMAkm0ijXmMVZM1y
8ILLa/12T5f3Ah1X8IJUC6hbxcTEWOIY9revFbrKpFhHRPqjdQOO0p6rGUnz7/eh
p9SNvrraWvmD32c7SwkvTxoFjeaFhacTY4/FAhSSefoKL3ScuepmuLeyt8+HTe1k
rsV3EY5dr57RJlcc/YR6r3tilRMxumNNllm6gMVwOfl2Jg3iA3PpGIHOXR5OtoL9
m0i/d+T/tOm3/of27zkUY8Ao+uzoOV+bmKNFHY9jkVl6FsG3L4KIAmku0bKGuOmu
BVn9cPpjq6WDFwZ6nyplFWI0tddIev85WTSJ7h+GXSQ1xCLp0vXCRIK+i+ZqbD4a
Uqh8nEwnTydQfHf68YxTV0ABVKljcN90Cq080kcBzzM6nND2ys/lqbjF6BHZFwd0
TQr9oMp4sRsVOphnOjB3D+/+xLCc6qxL4Wxo/9w93XHbifx07ar4RNxXZIfAJlhP
ZVK6SmDIIsQKou1t27cbmCpNcHNDkH9/6K8En0HHfe4AOkQ2lghShr/tNOnmfNOT
W6MlTn1FsOUrlC5H2WS0kB4tOcpFA2cJQhsXJku2cHrs/le7OAbWOX6cwd6FsiX4
y4+jfdjy0DcetsbPHLuSOfXqNPY6LY3y7pBUZmL/GpvUDBWzfc1HE4uL5i6A0JQ5
bSQZeVEJYsq13jR+yu1hKZFxK82PCYVyHamMgmP6H9ppeWMcEv1doZUbERwLKgdO
zMDDSpObMVDEaGM3IPEUbwDfycRHu6M8RQ8LhRFYBelDVhbfHG6lctOCZn78Knbz
e7YGmj8Ob3X3cdZPJBnhR9YFKynoGJclbzbDjjTLQvX5HP7VW8SnBWchhmlcJlR8
kGCa5Q24uhTwj4EIJhkHX71mcvYc4KHqXHpb91+Tbi9ZmWRbtPkzTJKcMfKt7j5a
U1SVKQobHauHwSCuG9vCcWgjZxS+qImbbQg2TY/MBN/S7XB6PGX7dl4hELPRcqx2
nuddBDSxNF/YZHNaZJv/Asr2m1D1XeskOO6mL24IGgx0hbhukYvpf0sGlqVbHOH6
MkFrTQPoQRY1NUuOhOzShvaGASTytwm5Kww5/yOZpt6ZlpA+4nZppHTCVjMoEDp5
yyOReFpRNN30ZIKB3zHiKfs8/VHjcv+qJAyz531K7vHDnMJX6ft3qJbbVdSUrwiN
LGNLBLwJCErYtOIHi3IFPr/nVw5zOGjAo0sPhUGLBXoWY6Fa2r9mzdUkX72IdiJ5
bnyTZh7ywy1mCA636Y9YnfpHR7T+332c1A51y4YcpwY3Wya0rmaceTxbQW8sF4RP
yAG7HeyNYKk2fcue2MetLmtnoOPFEt46PABrgd8BU1yGJ1peKLvxfL9agLW2adQO
DBLqLhXDIuyYXRGkjmuMqPEO6L5FJjCl6aVVAnT8sCfj/EDbBN4KgJfWPSxFB3xf
lU1UMUY9YFAAJFPnF22YLSOynha7WdYHvIJe2a3zQybNZloaXNOSoSwkf9trllt4
4KNMt6vHf8YkVZ/7jAI3bsrWLT27sNyl6ZkQCWC47+KTiYhkXtgE1PCRnGACoZDk
7YW3Z9hOmdEURP3iLIhAgs/B0ehLcZRXjOl+PpEfYw/1E95zdo0XmRhL3OdT7srz
9iZc02kN1bdB4YnOHvTN95vSHImSIHl+dUtoPOnoN8B33A6dkKQk3VWqy4+L4Svi
3sgDcT5H1FElKrQJyGAX9CcbXUpNYiehRzXAMW5wcQbnP7Am7LnQeKIAk+tgG9nk
F8CULQPB1KyDM20FC2t8ZE4CtUq3v1Fal6K8zbPFxlmlAPdb2/kI1gUz6GFfifHV
Atd5EUnGU5utHL8PP8UYh2b9zJfgafWbRZXvXRmJvLqQwK33KScpNU2Vk8kO4zA8
WA6tlZqredwoURa/k1MbJmDZie1CPkJXfkhtXJcetoYFFPSMfJwRHX18kSO8dugG
+7DwmY08vAhdej4stEVGrynONcrl1bi6Rm6kq2R5PyVx11aw86r1MVmEvkU/F5wO
X/crQbCVUmHtZF+O9Xeka8jtJLIZo7Bm852Lq+EvLJBBspCfKC22zF3yJSZHMWui
x2YPAK1yzkmlm/eZylk61Ezqt5dZSXCROlG7OI6Kpd7Xh7E8/bxdizrwkBrX9G6I
hq7FzVFJSZHDLNDImnVjrhjgGgDcvIhaaCLOrjRN5KhY2K2r6a3cypJEQzoHAya1
ScZbrVhLR94g/mA5zNWCaLt4rsjBVuc3ftGBheYXm6ZhJXRlE4XZnh9eeqx5n0wf
qHEELgnhtPebycIU8yWr9Z7UG4JfnNrnB/oAniXdhzTn9W0M69/KU219hfWLJ84h
q43FcYtbRw8jmwvpeJFPK2PxCdCbI+zbYOi/HfLDGVCDVxazPO1cUiT0tpHhI0GZ
CqKU2amb26vazji9X41lEvjY8zAInMiDzT52RZUKzLY+z54NWb4siuwGMQFn20sq
xHcHBeHoc61nOmcQ/MNU4fi/Ik10cxHm/Walj4cdJPXknrZKyjtMtYYwnKh0audZ
8wPJitri5uerY3JHNuuS+CTf9s7Pb/vEynkAUkIfg26tdEuBIANdGu6OsypHDZ8a
ldnxGEZp8eIfHeCDYLfjpY2efo5hwYzNbV5vSrwbXPRKWP0ki/83V9Vi9gsPuaId
vPYIucF1SbcaB44Vyop4U2JG6RrvRdT5CRR5MyjrNkawA6NNMlznFOmSltOnYalY
caXvz5rNU5X5TrtB8/+0oyB6GS+/v6H0F9NIgsO2INkIMZCnO3X2F/j4L6RqwcK5
rRGHcbF0JN+W0nO1Ig4NSa9yTBSlu0q+fdyRotwLmbmeAqwKLVvqqtfOM1x5jZYj
v8j8lHzkP0vkFfIw7Lj0k2vBkGNht4OrerToNuQxryYQcRRp7L6U2+rOD+wdT0jf
rulJxPOquadP/vfxczjDXrXV+Zf/BE9JME22IlaUCvXhC7TlBABBT0s4r7jqsmS2
16Fad6FZq1jMMX9C/yKzHhSkBsckz0Sj9cZphSM8mhgCwqjDxNXw/p0laWZkh61o
yMc/+41ImUpU88WjoLHgUzPwqFYfuNxPSFwQD9KXlNgR5N+XHObmLPDxt7U5/+bW
/qVevG2Kd7rH9pRvoql705dUPDTOjmNUL0F8mtibU7YspG6f9goDGJiE2N85eHhK
nhipPe5WI4csATjQQztCkx5vsCUEdw9UR+/Qj/AZ/ql5f3pwgQF5rage+L/BIu7W
JLh9a1hZCCi4L2rGuwO/uQXNXd7fdJSgyfjF0RhiEe3UZTGaWJD6jz8hIC2W1rq7
eWG/y2cBNhI7WUY3+EP0qfQlyI61+HpOYtxcma7iRbi8Rsy/3Niylsk3VZyPbfvc
2qZjO6CokHc/J2u6MAFpo5sZnftHCQvab2aNZW97LNpqUL5oF8ASE91o+temY605
B1ihAkzMBlfT66dCxQVOyumrEEawOvLQNGDmf28dhcDApQD20zeJ+D551mhvEtwK
kUFqE0piT1PBU5T0qb5MlTSCOwWiI/dgW8qzqwWZ+Eo8c0dCMkOmX3QFVxur3GHa
X3Gfy5RoNKfokpULPrxb5Qg7XzIDEM3SCoRlFumHo6iYWMeYwW2JVjeGkrSIWgSL
DOTMM1zxSA3Na2Kr7fNk6CmMf6FVAtwiKaf2OXCc3wjrXXaiOyiG0TpVwUVRh0tm
x3nDpBOpPjmEHJav7ISIXHNBC0AzjwKGfTXzMwUA1/baUvop8GMLiKX2x2uKA/95
AK4x6C3U2hZeJ9fTolFr6hxd1oOqtOXP8uFmaEEdeE7DJrcV845BufxNGH+p0bO5
Qu0HA8Jg8DbG0Zgr12B5KnKASYqyjcPTgD02TH9t+2nz3tdJV8RdZDxT7ZlrjzlM
ZlNUKph5qEOeMGsjfwWVLvkTvht42dfwDvyaXO9AGN1uXpFR5ErDtuVlftacP8Yu
k7WKsBKwzW7Lcfc4e9R1lTQjxteCcxL3hbtq6kxLoTCBPyGctXUJ8VKrh/Nbkxo6
d8u3Xvyh5lF5OHeJZNN5ycTnPgcT/lJhHbUX/vCmWu7Ev7YfiY14emTIrFvo5eFQ
XA0p5uNh6rpxCYL5XtAJkV/p2C86aMHFUM07AbQBrP/sezzbDndqt8T4+5nZQF7C
9NZPEcoIbxJ3ExB9VjQGMoxoLRF9RMvYwr1MNxjDVFIPWoNX9Je5tbXYg9a77WkF
m1XmAKe9G4rzIC9Earaei6Ovl/iFviBbWdps9q/9imJSkAYTDEhigBhyjjh6KrZz
KiAmdG/Cmd2n7AfYRk/0uY6iybNSgtWp60QYsNekTmxneymdprekHLBiy3TQgy9T
hewuITyEw2LzErriqElWOzggw33c4mEEV4NREBXkUWXfYfDShSqQlf1OO9Bfsvpr
A0EvGwcD1GomAX/wJVcIGiOgkWqszSNofj7KyTEMvwo2xy7kVuDCRmV9XPjMvW+B
MNJnltbS0zSbOFe/bPAJH2Q3sCjYK0WTqXxSn80dXOkxdt9EsbSQQmloaE3eu5yJ
3dOwUybg5L79f3Orx+Vbd69+s8yRdyxcIp2zh2Iu98yp0TItvfcvS2zXz371BCaV
s27sRM9vc0NXkiVZSU2CuuBDwqzEM8F0AAtghinISgROwfDKD6Kd3tru+xvKe2Cw
ZVi1Bp4dIBdD3ZqYABLrbRETagsrUV3zfSgxl6z4Np/oa5W3k0G3rzrr1D5pBDRr
somhBzr3A4A1egQ5PEY9DCiMPa/830036hT65JrfB8loFV4zjxosyIhtOaNoet6k
cT+mxDDZOuNfYQVd7IOTZermuFxvjd9HICkYVM1CpuDBwAz5rZIWiZY8L2GtqjXW
6uZQSW0jK1I/QJrw5SyX+YOgcvXwvAXr2N3BpH3unKj3LURanPVgW6JKtY4JNubX
TwKjOIAKvtbWuiyQaEPCStf24W4dccY7nlwty06ysSXMMFvkaV/RP4FfnOcORW9/
1dzzqFn08f7rZp95P5pOwYjzuveI4odFGP2OahLCD94SK4islp7NE0IAshMrrtcF
4ieqsrNnLTt+Hkva4b7Sk2cmrGfW3aTjiymM9N0Q9becaSBmngTZGbSh54Ew8Erz
X4sEdjxX9Xmpzq7oYbLc9Gm7vCi/DEFFXsJQumu1IZ65hA7SILTNsCmhFfqkUmPq
LJk5R9L9EMDD9Uvlx47hycEwjGqNbyYDtalCtm+apFrn0FHjyvD4FuY6nuWIxGQl
DON/RgEwaMHY74T3RPrTNM2sMfYK6CVrofuTlE3C3Qwirg1gFaikQI84tSj4q391
oZWYXyLvxNKYn+rYdd4XQ6GJ77bZNV0SYBcHOu4sHzT7DA/NOiPTTfoGFRX6UigY
cDsLZNw8j5afS/MXGgBizIU76XFr+tFFbAHPbCuRGCroYOVZ9oG5Iz6Nx3KBlN6m
S6vh2/XHMJd5IzdqRvKRoxRrE3NCvsQ+Rl/QJ7BaKD9DpG1OKNE09NJJ4HN6/YU8
FBLkBPgNjBbgM3vCB5EeZsplkScdt+Ojj6G/yM94iKXov3m0wRJTczwN+X2H8WhG
KtSn25p0yLTqUY6P6+V2JtnhSXGR3JNAxU9WeZLFRTUQiamWYyEcFEYFrM1pwM2p
NMlSDiL6nKigNFopY+gnQcOprXC/YRiLlfa8xI6hteRlPY4MhtpZZbRDyEQBqx7a
A8ncdNKfcuPuunVlqT3xQaxbYBd35nHyWXloPbxKcI/GEwi8sSGX5jWoVwgl9Zf3
hhVbKjiA8rO43LuNIzhw6qlg6M/zD4bpd3/y2BH23mIpxis+sppBYS+Fltvabwv5
zHZyo3WfiRfKWUo0xveViKYaT4oPqNcjIYHnamCgiEDT/LXK6hd74J2JuYTi7E/1
Z1D4GAaH1LAQzeg4Si4ehBLqMGY4tl47y3Zy4ZsJ7oeb04iKH/qguwu0AtmH6d9l
VYP/K3F1p5Dcahao+nzrn4VXiGTFkPNmvextl/0r3OgMmTGegQVjsJchZTFq2rKf
1s8aTT46O8DY8AOFMe6AyFnOpg4Wjm7frBeIZ86H2dtIeVXH2BCQEFMdD6if5h8z
YrQPCfLtmonGwYqG2nHmS3yxDd5wE1TtYgshadozjM3A2Kht6kz0E34n8T8F3njK
rlIg68OGiyEm8TjDy11pr/hl1xvBai4OpcCFyBUyfmRJK04FXpLdVWm3KQjzdSkT
3p1jwk3rtxI3KCF4DVGGVCqyJRzE9FdTBF4r3WmrGVWJBFlBnJ0WXWwaKsIQtF4O
hZXJ+DS/FCLc8SMKZ9bbIy8DCh+RTMgrOwnOPEM8qpv8iAVMDL1gR0VjpmC6jfv4
xBJcWt2gk4fwAw/OlPUVUgNQJTaWnH5yvzVdEDLOPziOth+5YTeH5Aze37Yec8hi
keYllG3XuF1OJKFVGe02mgMawTZL1KYsChG3E6B97Cvq0GMpovZKJqHMOlDnf+iz
qj0EckrlP3TfrvNW+Ypnaq6gwNUNst0Qch1ycjvxMl7LudOYKuSXv1hyxdS1HNNG
Q5vO0if0yNy95Q4Hjqvh2vlkbaJGj8VoI/TPqf3PfUfPmbeQtVzWGm2YzIhIsr+e
+mUxOvyO1F30mDbtxb3HrASUjYeD/gan1tDK94H92wBdpy5DK2FkUiX1bTDL+bN6
SfJzh5xul6/LeBBXea2QQUuUL5iR+z3Kmf+EBlCHV76dEQ4oL+ugJsQbU77s9oFn
PeXYhR7d0UbHXgcNrj5um9t7WE9bpLLbFt3HfO1vy0icf1KqVk+VyL1wEffkUDLB
M3nwKIgpTF+Edlm8l+xpaRY6Gsn8avKxCFDrxmhGglaXUbZQyApXePyykPHwM7TT
wUz94ScQFejy2c+UMmwmR6zdLNyjaf50agS7+sy6fmLIWWvGgsBf8USfKEVmAGOu
sxDXbhi9itooKpnbpjTZ46CuaI/I5AcyShpgZMLGsSp3T05YsQmkXDSf8FZu19DR
1kfuSnxCqX8AC2yhjUZGA3NkvtnVPXWISx0QMTp4KeF6aRU0HSxtS7IEXpY1Qlsq
JQ0zZ+67Nh4P7JJDuUuHSggfmqxrGvtTXkDl1eT7JrV9zj455cJcu/TyOCX0XdIO
P52PAedI6w40CrQXROfJyYkzG1w8yav/1T4dX9pbRR4wlk6MAm4f+Snfe+yPJVVP
4q724Yam2m9bmAc83e46b+cHijvKoO2FYmGCnpHyVXorcL3YVUz9hAlNgEr38b1C
RbJoVWtOp0X4wQbHkqDgE5Zcgs6uEHJoXSul5D53nEEO5sVtyPfkoCBCCcn7nDAu
MLZc1tyqnaEKShc5cDyoREK1de4NdpY3PaH+Dd5ePdOG+EZtkkwQWO6Gbw3Tmcjv
B3RUvNXUeoEio8whyX15tO9oTEGARM64CcypRUxsNqi69873pPq9fVtpLdKsp+o6
9IE4Ln2yuIn/O7MuuW9RJ+EPTFL5pKOytgKQ4L89YFbMZXIHA795VYRcwATaqsfF
oNE1DLW35GRobn1hrBJY25x4Mp6Erf8IGzRz9zfaqnxq/28Q+nYQvZzmoi087Tf1
5XMMSJXuyaw732HCaMdtC2w/AYmoxbxnb8Up7NNvHUnAJxPkHw4fxVCV6nhhvLAh
IgVmHi9iipw8h7UIqms/KwP3XN3ysJ7Rr9G3bBKpeMcKQHFThJsVNA2oZtpIKaGI
MM/RCSVei2oJT700RzhWS6vsTlzevZ6Ym3+H3IT3n3NWn7nmSc3cp9bZCPNSqPlF
Cyt+5/pLGnrUFpBQQwOFo+YmTPfuLxRscck6nS3FfEL2Zg38BGtKNacU/4AtfzXs
dB7FYo2aiq18t8DufdsKYWF/On7SILI7L3Ja77qVFazw7CKg0aMU4d2CmhPANEzg
IhUdlp/ZFEd/+pU66rGS6xVwuN+qxMfVPFJiNP+ksAZNtOWP23Mq6xY4oDhSC7DX
izvi8iyPPjU+zO4R9z+QsvSV033Xy4RV6jwxn2hXi5ALhomyxRbv1qYEdWfV6kV4
Q1GZ3NPml68Bym8+Ve7TTw3J5FDVEr5ULLaSLXQcfB7VPVfRv+te9Irv2iOJMYWC
2UyMg0GsaW3lh/0u0d10iQcr2m+bocXYaX/K/YrY39tlLAnZ0FrLLLyTJ4qjK2Rf
SiWRJMdoCBxs0lmSY2MYcEaL0JV8qz/e9yUOV9vnmniSzq9wGEGc0AMhEewMJ6XL
Bn0SdYgY4KAvsNPseo+dVnmbxAPHUoGBOZ8/6SK5Y0oQqAFotRxwvD62tZGDutq6
qom7qewHmUbHC3f6GlQZz9/MByLkQbwjD6NoZ55Ta1SlWGPamZMtip4VB4A1tFWh
KzvMvINy8gFxJ9fYajJYr1fbg6p6A9e708ElCX282juSVA4P5lohSdHOJSjpvHw9
WTRIOYHLzo36SA7t0sTkm9ZRnecgptrFteJeSctA6GUyQW0MSoqJ6t47RuW9Z7hB
eNjW5qhoHgk8q64+MH4HVt4Tl2r+SztZOhnI2GXD9i90h3P8K3ZPvqfXPIEEJ7k/
mf74V8ogwX2kgFKFzf2JUwjMkd/ghdDIv9Rr9G/e1e6CPjSwFSP1hCPlj0O14q42
v0ZU/zxyIB13ARgGw4vv/BM0M3rEYxLx1xyU6NrO65eeA6VYlqVpoen8mExTyk+D
8oxt0PiKvJ38HuCuOaj2ZKrcYViHsl2PPk4m8ncQLTcgrWgHnVNaGf7rta3U425c
ZlqWDcZWyWRqboi/dQ3CgBHpemXSgqG9WNEzHQJTz+D9DILfzKaGbPYDESqpsSmW
br3olIa0e3wFD7RB2dS39VzKBRe7dMVEK3NTmAR79k2kJILQdZ1YhrypUT53KEmV
n+Uh5Dc8iZLmnNeJICFwZqMEfBL5ngirjNFJVae39+wJStxFzgaTiw6lkOmnTYnV
T3jHtKa9sf+P69V00aHiPmgYxVyMV2H+wzU3pyUi7GaSeCtqSRjfuqrHINspHRGL
IN2shIuRN32TZpFWLYTLbR66dHjlniMzkr7iA+3GkxWnQdoaA4HSghEVjTqBd1Nu
2spPLTi5OG2Y6p0HAzI5fy2eMSfrZVYgMGfi1t6VJ9nHWrbX9GvFOLELSYn03S0e
WgZsqvbK1MCqVZtZuHf7A4gAg7WqkYFALL5/DVmKiqizGEYbffQdafR3LuJoTOa1
eNo8CN/xOGS10a4DpJt47jC6Q/bHW9jcxP8KgUXzHdLIQxyUyOokXpyoMTkRIGYJ
b8eAxYCIDE0ptjk3epimL68IepG7IbEZ8kSABqABi5+sL20Fvzc/hG510cSNzGjX
4yjml12viflLZCtqVJGV4mMPubMWuP1k36cphoH3R73DhZ1q4bqL3v1txvlnS3LM
4bsliEIoYaXUlK/K0JtpUQQjXyz077NK31NqnYDzQsGhaMCqJyk2S8/aOAe3KJ21
9JGhYtoo+YRRA0D6gAYswzu5jS/1fTglu9zon7QweZ9airM75cyNZNWqIlJ+IURk
5uqOPEkKMjyc9ESieTTkg2yBa39pwxahZtGOoI7cKT3n4Lvjks9TJoIsOw/lqvy+
o4YFZKnjB5hfdKJX4ye/EknQg8Sjkw4rhi3zbp4ZbrWtluMU5lngEy4qdGAFu5Qd
NzZ7TqIQ+63BR/eCtMLumVTao5aN7Oflsx3kO0O8/5lpwuSpIcbsa/ZiMkwNxW1C
itNlXc+2lACXsGkBZfPrAXKHWetG0XZObiMoz2FF4DdPQlAKyBmfLpXvvaVAwRfW
pCrOGiF13QXo5b1MGXdqmMG1MbQqk53WyKFYfrY6DnoJgHbfs+y3uixW9bkKIu8L
05jQ8z3APfrr4ax+1x+1DO6UCGHaX0j3Hne8BjU1r/uuycO2uwCAM3/MJZhisWtp
Gpbue8+jsm+2LmU4dZv4xHWATQbkPWUo0HwAbkHQI1IG5r4qFd8w2PZlmxDn0vpx
VXkuQKCiG/+RpQkCOtJbffcxvRtBkTNqm4qjJcCUV7irDF608BdPc3e0tgNajyZJ
YL5fO8ITeTke0Q0S+9H/aXvRvkTEJ/eq4uDb9kjANHs/zZzd6rsDcQnlN2orpJQT
n5knd4627Az/7/cBqTyyhckh1ygXZeRT9EE2/7W2J508/c0e95quaeHirnZ511Tf
7xKz91Q/pFU7U7sOZlsMJr3AencmosWtyaEd+hBFPxmWOaC3V3HJYaShhjqIisBj
2k49oKdHoSDErMdvRfoY/Y/eP3XIljYCEjKpMvotJIFDhyeg8TOstYrlxXz82/2w
rIIk4IaSRK2tc3sIGT+eyUtgpIKsA/tvHwtXPYA6YLOfXYKzoVQiPQu2hF/c9B1G
mFHJuFhxJLfujv4+xJ3bNV2gNrpkkT4Hy1ogGMHWhqq7BUQdSYZIWslu7jCfH6t5
kTA0zkHcuiHHnx+xDOSu0FtyFw4YU+2qE/vadU7C+p92mZUy+aM74H8GjLl66LuB
2eeJMmpIkcxHEHihS+kY11mtJgShqRf9M010AtcHAlOBMtdvKvvvnmCu8G1P6LqW
awVVv468yMyfT7E3S9IVAN9HRAUknfnwmD3dVWnTYg1QaZZ3ZdSC2jrTWCMMjaGS
CKthF0ggflvJIMjey6aRCelxkwsL0Du4Ah0dHEPTFHA7QkdhCQg2BjbwQaljZIoA
2qfA4pnEAiC3DWdo5KNTfYioH2H908iG6OswnqQUww7OFcswjp/0nebyfhDHOx19
ICIoT3nYV5aAaD60rCgPJpINd8Kg4NXhRIkNIbJToJBDYaprlZiAI9yTFpNItFt/
roRoLTrzort8Q/xC8wDMcxnT0OR9q5+NWPV+/aqueIWZF00F/gpVFerW/7U73+Jw
XlXvSil89CqPDoKMJC1MYNswEbhjQluzsA1Aea/4S1bFQnSWjGO520105wtfMmxD
3b5eMazI1dqzRDAFi26pXvvOaa5hfssUE0qAx4q0rYeuDQvMiQKLXgxrdc9Z3Aks
GdgPg12JWG7l9xa4yFjv/eFt2URPeCVaT7Qpwtjq+/RH4q2CInCs5nUs5+arMg1d
RLDUzV17xycm4pLYvZ3uRv+bWcxt69UDN4EcrPlYF9iB5fL/mJLbdxLoatK2vqNa
cwf3eA4txjmu50sL6QSOb0zyJHeGCFVhCRYdrTbnNrgZzRErOg0i08CLl//rv+4u
ZyVAU0A72BAq0q2mNf8ErwP6TkNuKREbFzdISiTSff8lS3lPKMPRJmX6ZRyfC2o1
OxyHOes1vnuXdVJpeRkmCzl5dPxhDOpiRfENGOszhjybULMZ+6h9acUJJ3UAl8C3
lkHY6YB9hWyGSGfckQ5I2ciIckszNRaPIeUwCEGKOTa6z/Nc9rmSV+VgKMgMNzsi
ofzkj7xrE00TYJnEZ8Zf3gXAbUH6fNleHWIsdEhRszsygl2TwF+LVzM8L1GXRiIJ
Zi7UiZutiG9IZjILpaxUUKbK6vk1CnInUFCZVA6ahxChyZAiz7gMkVGYKSCm8NtY
J7jyJ8x/3Azd1etb7pB323mpAb625dfzuuy+uJOQZJ5nDNYuCMG5SvSZf799q6BL
qE0uCfSXifB5bai7pPcq64yYpE0YjZawzMnSL+g4HUsmgTxjoR19dE1MgJGn2ljZ
rU0jtAurtK2YcLUMKmmJNBugM7hAn14Io+JWutYXG0EXe7Iy5bVRYvQg6/kYWmlR
VAqVWDqld8u9HIwF2sFwWN1fbFyu/cFF96KKu34Ij7SsP1zXRuw0G1VZSEpUqLnf
YEicOyLuuJmj76xqrQoaCqlQmiGBlNl4OhW3ghuNVSshl9G1lNefCx5qKPB1JNdl
QVwqmgGzwqHAMg+yomIwbEae191odKtW+bgo/tgxdCZuusKIdPXOzPlrppfL07gV
HrqCcVH86q4S3okdefGID4ITQtOJ8viZSCncM2//hpx39/N4NIdwpoMRJVNkcWlR
NIBxzRFECHg5Z1SKrC09fCgS1IIpwDVWD+R+i3SowFC3+lOT+x9xNC3tWzZQrhW8
jhyckg2t9z0L1KYC9zIzwe/bdjw5+xtA7wwzVN86Ld0ddEM9eSAy0HQkxeBw1T2H
ZHD88V7hftz53xBmG+kT2N/sNzHJaaD1QQaI2q3HrxMi4jPVMgRaBGoYPnJ2hOwj
VEl7kPPZ8HBgwZ69ntv1CQQLH5TCKLDPJ0RFS2/Sf4tCQYB6Rn+B/uIsFSJZvnBg
b0mf6VuouBCFXzlODHyEwEjvKLew/kh37q2DI2YC0zssN5GwWP83tMgJxwlPyzsC
Xr5Lfog622zMXbZuPErxzxEensKbW2eSoQZnx3YccKedH3G42Qwslcld4wvAqXS0
+WERSO3vp9k6zMvzFf1A7ekm0oD/p4a1KKDBQmZ3IZkpVvUrSibdqgFaMkIJhUed
fCk7kuKBAyXtJGVQBVd4/TNU2OBfF3i/TbmcJSN1WU7Pmrrganzca6QpNcKWmtHi
EEwT7dnwomxPUm5U1smy3W5XtaVi/a37OBkTxDdXHFECk0innP7c2/YDKI5ERnmO
5MDmI9kRHa2olX9isTS522SHp/+6lhvhafqbucLtCx8kzkMvq+M2bqebM8SqEHus
VZxF9zudahCOy4JoUA/DdA203kfXb66eZivvIeQLqOg7ax11iV98xJ+L0v6VBYQ9
gALNxM1GjtJDzZfsVkf6PWsoWU0KwpSaSuTIqKi56dsp1p6eiZamkorld0uCPVRq
vvnqtPWvh0cYt68V8DXh45LVf4WEEgLZZ16KCHlgAr577S7bs8EC4/4jcLHf2Y4A
sWQtq2QTuAZzpIrnXUUU827Ly4BAogQswEspXxDue319CS6KPSetGqgAX0UK+RFL
rJaYREyK5GsreEATZKSMAj8a51diDtvPyYeLKGm421GaG0i7YWUT3YNeSTxuliFU
uey30gDmxz1vJ6zrtThMb+w7EDWBmqIT6ylpX4KnsdGsC2O3Hst6xQqyKxiqqS0E
4S6vEOmKATsGchANJwH338rO9MENTasLZziT4IOxJ4BDJf+1WI5WGcL1qwPImG0z
1L1hZySbcrM545y9pdoFi2Txc9XpiM6J5QebgUrzRqVppWVIumMfZ9vJTt58Yum+
clhuxL9vNtyaPA8ypQnHjOw1zZRuqkOWpGzWzn3wUL9cPEIwuy6+MduXBZ5xmoG4
JerhdAA5GNNscryKLsA2cnwqSFDY4qNFDDY/nS09009E6rPbb5nF8m5UJYEKYxnK
NCrk33wGhtqMTTLO3xwC0rEw6/X9KwqarjUVOoxBaXNocqwgVY/hX1FMazrByrWh
doMMbBuHfbEeSMvuS6Wf1n9EZ73A0cRpJax/ylpKn9ynmzFQqdFuDBz+4P9MbWsn
c2hutzlRaoqEMtyPSwMc38BOhVKXgwDnezNKmalvYtSJh+egwSyMDNgMUCq9SPtY
Bmyx3zHehPTVqg3DmQ946CBcydC+8uCzH/KbyObJIlTj+c37JR/lgW5V8LnvtifN
UMnnPsTvK5Qjhqr3Tol9Q1n/Y1QZa2kglGiqmGzwg1yp4Av3F5PRK5uzzvrpNlB2
SaFxv2VufWIMxUDiiVyIwKb1UJbOwVbDFlS0dYY0jyJ0aW2huKK0K2SVtFsqztWf
cd2VnmwTTyKcK7+JmDP/tv87AhJiqVmX4lvFCcnOuBxaa7+dTwYzbPv6F6/0XvtR
8z2myjdZFO59rrhnxONw/AtaYaARpxh3f5qZhd9jxsk6LlKQfxUk68gWYRJzLrd3
q99PPY9kinrZskHGXIJycC8CdhBN2t9wNbuQTtVXRugFjsiYCt4sv5UNPE5VcN/9
wKjfJCtYGmDFSmU9aWvD4k8l5x6kM2MoyAhnVlmE34M3kBFjFr5E9gN+pEKZujMn
bp8YUuEWDmKgxyz+yFyAbKPVjrt4mW//dQinbmCS1iI3l3llP9uyMYh7tjeijZmt
mudvKbpAEIKtzyTkM+D1yStHaQT/79R9LYt37TA0NzAOQA35vq7EihKcRDZvfKZ6
Jx952RLGdtpWTeiBoPgy67MDtooaIiJyiFatSG7eeoy+lCAmezajg2loLUY5bzGK
QQyVQ9sRzfx6W7AWRGB3Je8+8gI84YW5Apew2LLZ0kwn8C0ySua2hm9bcuZIOk7W
JGeE+iNuTv9NnNYWzDu08oc7a3J6xSBJNtbocRmlhxxVC8YHGEWH6emr/mPL9jqM
cEKzYngrheIrssRJAUrDXOY3HKw8Zry7EWF/gIxhAmyWHISPis5c5GyFf6uEeOAK
yvY5Lw1BvRJqvhJLtRbBrFKoyYRCk9+SfugC+u4m+/5b2WkkkK73Er/0YtRufx+0
QSH1uf6K2UlyahbhK90sX+BlA4+MWBiqnARYUNteStNNBxbCbmQzBQCbS98lA5lb
9SSjE+4CoT3Z1p7ckoVCcEEXcxi9GbSc6t3Ap4ZjdxjO4+j65P9dHpIRGcNkwEyf
OdOVzRTI1VbNVreHxH7AKp96/8ZG3SqpOSzhWKAfXpkJ2QCF6mv/EecrGg89wU/X
auVgJXfE66NKvhrNW5dgJEEiuD51JgmgfJeqF0+Z+FeUorlRtGDtluYjUks0YZBj
aIsC1MTmqOR/9kza+x8VkZZHfWPydS1nsWdE4lNuFvRgbYKUFVvK/VTsL2YpfEG/
W5WiKEGE66KbPxG+v6eV0fAEXa0M3f8iDsN3AYF8fLuHut4ur10wGCMx4VpYWIcm
RPpfO1x8po0FKeSe1CzTQ5/JZLtWqQIReIcG9dzVhpICrarmOPKj+VTWZ7bsB3m2
P1iqSkJn0A9nbVb6fLW/zkl8a/JVsoAUE6IAW5k7ciyoXxaLj+x0pwAr39+dNaQf
Ei0Wl6B97qbUGfrHkFPnrGpmoSTEqE5440AknaIQyFATGZtUta/J4ZNLSnt0S1cV
3ZpkDcM+2oXb2Jzyp6rTH33qMhang83mcSWa+R3GKH2mLNzziDNm18FBuGGHtTJQ
16zhAd9vD0nvwLs3izG++oqGpJTIcFQVKyi/C12VmY4ETxafTo54j8bZjBKOffvO
wBzsD7gAiT3Bep0KJ70GzswWfuHLcRWZkEWm3AeLaXlixdOaAJcU8PZsYRRrEitV
PZZA9/QeomZLKPBbTXPUntEPJUMMBw7Dq0OEQD8W+vWFKiuaJUxUT8E8KFjYdW/w
8tTLqmnh5MCFJynngNCVRDOvPUCqEFhGrEp9GDLFnWnwNuhHOOhCMZbkN5lvXHuN
aWee/9ufgO4TZcFB5OPwnI7hupiuYtiWRMCJF429SgpjFp+e49TNQn7D/GSE5E4K
b6bMXEm+nQ1O01fKM5blfqVK6V7CwT5z7jLc9vqYghwq0FDvH4KqtBMvFWMJh6I5
j4tj7jFJJXbqG0+wnOIfGUqlQPP1N4oIyWYN/OP4AIGYdZDjuKd+MmLwQIpXZZqH
2SaRNse2Md6Rl9pWdc8qcr4Zf7sNH6gySP+MVOKBXnPPg+CsN5Iq7fYuXt9XR4+1
/7q4wbI8+qMZe/e62a1HirSFhb2Jo8CZm/0BGNhlk9ibZL2i+LwhfO/iSSFpXOX6
NJdqx11uZl2RWLMWHsUr444nWtQZKfuXbt1PZ0/8wzjKHbwgLP9AfaRzyIKVNeY1
4lvb6ktYaGCllY40FhuXbnRXYrIaslM/QFTdhWinQa00Dt6BqvqUcA8MBhfw3dJP
AjU1LezVSqnq5OYA/IEIlXYMbI1y8DpecEMG8/trfYXDChAocFkMBv4zmGGKnEy5
blUdDpTlLsNlSQGkR+uFfr7uUkyf5kjYjkwqF2DtHtESH/UAG9rJ5h5HUqHkSr5Z
VwmR8Ccsw/jNiS/G9iQwZ5UPT2f7nYCNujdxffVP6BpyuR2fCuIVwoWfy7Ebql6J
dEfx/K3RAz8zc/L8LC3dpa3KHsG/46aQKKxvBjYSTL1dRLWp58B4zuIJlWQHXJPa
0cHb+q+Ts+hkhFtRGILktt63yur35TF8wuwW8JQlRrtw4HlzRPe2DnEVmaVawMRg
ekOzJBXEovvcXXLiTgO9KKEC89FPST2CmyqmS4AJ8LrUAwR0U+vrJ+cOGZmNwNFD
KKavmRiEyjEMd4HBauQ1MifB8U3hMaLyqSKP0RiDdg8GP2BSI31Vg0OEvll4BPD4
r4p2ELaDUYxcmB/M5bT1wY6Rvfn+YGd5vL04IB0aXelbaM8FIxiJpcXhXdAOtmkp
R9d0fOVo3EQvQi+AedQ47OEljR08r7+0vkvns1U9XcMBcd0eW9wmStTlvEn6yBAM
MqcLE+MMUMfMz/3qlBOhGMzcKmh2/16ga5iZCXiQtYl75znZvYbzAhxdkIPer8yI
n/YGLjrOUwKMEGoB0G+AGbHfg5BEKIy+5tqTgKMOFuyEzLF15IFrFwXDoQ8/wAom
Rxvk0OzfXkAOCnILOncZIyDmzzz41Lyc5A8jKQGFEHGtPY1QOo7aS4oZ8VXfJn4D
h8/DyYd7ERWDBEC6YiXSNhTqqUbVC4ZqTODMo/njoVKZ7a3ldRSIWz4kcekp04gi
eHKTXhT56lQie+9OCUoW3XazLKjMoj6Qc1pSr3ltgifJrP06OLc17izVq9q1jfyD
4BWAmFBF1Mqw6uy/BzFyNR/PzNb770PjFQHyagkKc8KH+P3KQfX86iCmdEvtTCh2
F+bKEHNTXbXkXBO+Ij1q47fslETY/1oI/5ZkCZDeV9eip/vMfylRQe3hUPeVID17
z1qc7nPFkER56Cv7Qcqh99FH2EepdfORhGLG6sN3MZHwSa6wlLFAPYRrt3w0VoFg
jj10qLQGtMj8bwAK4etBzXTRG2fqs9JnWKtoIz6o61+DTxvaGNcxrIantS+vTWG8
eySVZFENjHENkUcGhZg4Pe1kxO6Jf2a2K69/6rpp5r4P7O706ml2PJ/NoTlZlDJP
rNRd1X7DIGfERrxWxPS6gVc0bP1nog7muL9Yvje5CBwK+j8gXYz2Igg52UmB22eF
fg4NDjinVBH7gVpgx3jgNHYgo3lPLw7zt/VCthQ69ZfUHCbi1dSLfU9f3pTIutH1
zAZkc0hZH1Lb0TmyYMW49unTyJLJoEo1fWn5QymQn/yEi2WSNnyvodtYBQeQ05gC
F5YLQaFfvxYnSA8KlBsJIhsle/eHv0HEisqnlPNaoHraxP/jJIfQ0TnvvAzj2gBE
bP9E/Df1sUkbyw5leAMlJFnjoh8XKKh97QDfwcBb0fi2QyNn7ytGG/PRmI0jVVgM
MT0+g8WZTMyMEq9E6ge9x1fH+jtskKQiUIdn+q939vO7oppnW0SNGwOs0gn6XhF4
Y6pFvmpMo/ujtdZrlIxNKIvIl1H4WZUBCIRYLRnj/n0N5ZC9IBtC2+PcqqvLpN2B
tY+ji/GIBb/O8+8R702m0cfMngJwSmoo6M6cP2EWXaCGTJtOdUo0zwJLgkx/aq2z
q3HbIPAwnaZtJ0Iq7ECD/vcD67CRU8sMm3HppZwr8yc5XTc1lnLIJoux78JZoZds
CV/t19+Vy8xM5Xk5Xo/s/koC5pT9K4FfONs0tvWaPbCp99AV+9Fzd4hanyAllwQp
tGbrhjB460cUibhMUxedQn1b02bBelE5XmAMluJKLqaMfEvn7UkTntRDgr5ro3Ka
6hYU5Ajpi644drxyDmGb0lgtdkfJaWfONbI5VhV7AguMK8mMPqqxkiBvSPTbiP7o
6QPsHwTQR0zdNy+vjZovitaJRT0utfaX4p55qry/4rVEJdIdwg2BYH2M92snl9l0
yeOm/i0u+XQEOMGsw3IoiPXLpAHuTgPtUuJJ2aDAaFEUUurGeovfWRUChIpxlm/e
kM/HQIVZamzdmO+xZmhEtAJn5xy/MyTDyGn99ZWynQil+S1PjECc/m6of30aEWDY
A6wtapBWEzFRc7nRP8Eauh2bswBaEvU+Kq3KLK/yxw/DfkdfrYIAEa+RlZrPB4/k
FwsGSl8XMlVpRdEBGYPIKstkfhcU3PBfszoiCAxgZEfr9T7q+6nDXND0xKUGkK72
hNTymjLCfB5dqomT9La7zbASECjllFiDeiGtHOXfRkOmwpNFOrGos0lwIpX7JHri
0lQWO4SSMb1mvyZvvYFJhdS2rVQOMCZo7AkDegpmLvGWH1ovI5NVZefJgJdo5FUY
vbVdcqNJlGTEnRdJZ/I7G4C1ZVbtp5lozS1dfDOYOIvpjzNwpAWakU52cu6pSMeE
otjTmIfCeznrZryd69qD7RPBZgjk38DRZmsFHDYv7ta8I5A/ptxA4lFF7ZSD5inU
jxIURJ3KcI6g9XOUGhUW997YkrZSmcf1mxvc8DQgFbQ4K1h6nUK5n6lqHhy8gxqa
ZEE7J+FEUumS6ztoqnycFxYMoJTIIkmhxihHOy7zfZpsV6Y+r1DfjJJPKle1nqrD
fchPG8VyPDif+wvx9CGRTiybTbL0oIMF+yQFMHeugnk7pqXc5H1UvtP+EIlZMLBk
5eGukZlqUBS4mubJDJRRXS0/AATtFmVUKnPMgoFGCVU8MrPyiYhltyX6ZTkv8JbT
4R4+wEwrCCLLT8xz7XlSq42JOQDy4Tb0yIeUywnpHaT/YgF5sfnxIVDregklQjrj
9iJS/2q+Zobf13OyL9TCasM5glSaOOChHQlsF6UmavJ6rU8Gvp+bqMTD2E4HGfBg
S/3FHIWidXyPcqyRvhda86MuxUCyk5cOQZoRth5fhwfIb9mMrfKPp/xalFrpDOyV
kaMbcWs1O7ImWqoipxP7pQ2hsrzIJi0maWlOY6jf4pQTS5l1cHYyUiEC4Ys7wHdL
My4FpSu1GM5gWuCVLmrCX0VpqxA121GSb6pAdoNX3rjs2pWQzDRcT/Rlxi8tDsfM
mqe7Lwa19LHXfVEol+Fb3lDFBgvku+onZgY74qxXItFyJMCSYkC5d6jSgqeVmO9z
l0R2bOIsi4TO4z75vrzeN3Uh4VPE2lebDqWYAeE1RXZBUGCWhs9XFQrh6Lt0ORoN
Fqv528gHFD8T1qT4GGFNf5I1h5XSmsy2HRiiSP87FBh4ZNhit6KbHYlSLMdZurV8
fxphF1n8mn5B9x8JTYW9OGapTBxDPgMPLp2Pj0WirBHj4Mx9fJCrdsGd5xuT/xxn
+MQXbKzeqMVoyeqBOhanbALzmz0xFz7jn9iYV0RQDHjIErr/6fIzCWPm6aZj8eNb
YllH2Rqox2QXce+e4MJTLq9tHFoj0ffMvdbfWj8s44W0tnLRl7BWKRP0Aj4hciBu
o2cJk2N7mxgujcPUBPSX3EK9aWbUqrMGtaxa6lgnw2f+bCqS5zJ9m95fZsg4j6Mk
Qcu8B/IpIXZeOGcgOkZwQBrM0y1550PSl/KCN48vqbeBJgdsGdu1KI+CF35Oz7rq
Lods746kqUNJvLBdtHkKnv46swRuZmhA9MKM86CPImFu0rPLadCTf66KXVFSfdl+
pe/QUrZmWZl8KdwRFXAonFho6EA26Z14kykQz/F8321v6aDckkcncSwScJV1S+xl
IkaB91qwb2kip+2Bn562MIel5ipHbXmaNtIH73W95Oyc7UYVZP4zpjdLnjNwevdN
IIsUmDJeERQWiyPK7pcxaHZ0zuhdqm8QSd8xPjdVLQS0HhpT6tGwjm332WK1ziW6
9SqkhVMdQSS+WK7FqFuKXFPp/L7WucCIuPSpjmO4vZApcyS2/OIbGZWbPcK7qYYj
903HMN2hjfgT8BahWdsM9PMTJlgHS7K/zC/mdfJxCmMHNRaFVGXZJTyjtRJp6II6
+P2/IScyP2TlmsrlFsgwd1Tpwz30AVPO5pzUEF7YjhSUwgGzniKZry1pcDYzr06j
/33Vwjl5e8dXuy3fJ/UaVF34EUVgArxSsRvaC4bnYRtlVUDdax3HZPsece2RlRS9
jrdbKt/EljdfjJtRU1oFcLFiernYO7d5oAiSnmPvS9Oz2knmmhDBE4GAQ09KMi6E
hKaB4YRmMtywIaCrCHpi0Nq7aYJO1jUuvHVtbVE0kAR0m/jKjINYMdWx7FD5W7jD
DmCrqEgKcgPs+r+lA+WCgjroEQadls3jrknLuftlsIn1q+uTQ3GsWh4WhjPRfHFD
OYOHzaK9vQjcfos+Lh8xw1neLofzkUqCLH1vmgRiMlmRiC9sNZlmZ2s8SyMePMih
wSw3AatvGWyawH4gOyED0Bj6I0Xb1PB6PdL0av/EFzFyKdkf8+8gdLksF6GtmWVC
RuCZxTyWUlc5RukpDDvXPnM4dWTl3MqUCVlhWDpfQnRI1e5t7Uvtat+nJJBasiD/
g7R6oM+jXuIHnFAiX32bd+Y5sAZC1u8JgmnWGaEZApWsQq74n9hWHjGXdAtcEDOv
sbIlqdU6ru3DODoqaj71y5fdziV1IDpWSVVeaW+lVrQMtHANh8S7uAdPkoAxNMAE
RsuexGr8IT+sGL9BuHhPg7ArLElGAlMIn1d4VERxBWBmZmI9apzm4Y/myK6/66pc
5It/C/lbB5WTUn7sqjmeLX1EFL+M3FvpSQ/0RdsiAOT8kGuJSLjQaMWZC+lXaabF
72TtE6A6h4xGwi5KmXgzryLJ2MNRTqUzcqFX517N9OKIuPtUP5rmorbiODxch2Pr
40CqFMziFUUich9wG9+CpXpn5lDZGdaJ7upUCclupnjIYBntsA0S3BxwWyxT/wi1
i93oFl80vUEwCQXAHoDs231X4w7FfHTs/f+NfHC4htCnQCQp6U5HKJrJJ/pshNFX
9KjWcpcxrlZHdzih/PZwLoUq6mQYdkv8Diy6DkDijRXavpop/F4klTI5NjlqmAeJ
RxfHzcsjB4QMLidCgR1Puk0h7YR/JccGrCQTA3+fA3ZMJRqFiLPVpzIEMAAfvDda
2He//52wqIDLyhIL7kQWfBDYGo/95YJozx7JqSea15kh39Zom1jWmtT1uJJR6T2f
z+06TgraRl7LCwRNlCFZVYS/nBBtw5mcqcZWzxSS63eQK+1CZT+oeBi+BMGUXjDM
ECx90ccLnV/M0ZHTJ/0vTK/hcgfbhnxcsPFEXQQLrIYKOnypKFpUdWKqzYRX5tuT
4nSpuwmVHfiWNkBZQS+a5b5tLzCv1sA8jw2gXo91LniaBeeDA4VBOwO76W7PNfRF
QkgGkbi7nN5iNqIyqUokrUfeSVw17OIIoLybNBwO24PgwpqO3RbgUr2roHTq4RV1
+ivrhR1uSZV6fhuEp5hfUlj+pZFe+lOJ0+JlfEInNqvljEiUxNrUe1xlMTHy4xS6
+CkX3NTx5UDcE/D9I35KE47b97IUCg87/v+Ai5FX36BZADCcq8yWacz0PIg2DGNR
O5tw5pwaY7sVoH4Rxnb8L19duWTodW8+9IPyMAJ5eOaF5kNslZHm+N/5qj3Kdy7L
JyPA6eC94AFOwmzkaQZ3MePozgkD9RTaf8HLOfUA74gs3Zq0MGoZgcd/OAZ2oOAg
AqQXYQ1K+G9CRiqpj6Lu6ooepLxEiScmnyzaMu7p9eQb+RgDniC/Hi7pjwz/jx0k
fz7bu622jgnTWoJBsyem/gxa2PGzZ+PJEHDHFTqD+e1e4uQFws7TrndHDT1OcwYF
1BXtU/UVnIeTZh25unR/jaFYjfDKZrUi18ItDlLv0WeglMJdt3W6Qyz6QN3/wvTa
CA5u5V8kmRH5BKzS5TYfnqMwk2DhhArcmrKVjDbYyG7J9K6JhawrKI43dZrrhw7V
uKFpedrh+A0sIeJoxCseniw/BAR/voHrfFXw/DUnSlAi+37OXL8fd8kMCwEwz3cT
yNrE1VXasoVbeLIBpjK7odEZ9C4qhsDbCLWdwhuD2HoyW4xP3WFk0c3X8yrF57Nk
fQH8nYOOQae4vOsIwflgij9AfXQ8XrhwEv3EwJPRCT9tw8p54yW1438oBmaOdo75
5eAgqNOIKE+30sdiX1Q9tMy6lsJrcuZYKm0rSuRC+JEiVb+6T+FoCZy57mnMyjQA
7vRFUZtqZ7iQ2ySytTQBSjGnFD4enTXyXLhEZ8AWdTdQqTb2GogdJHUq+OQ0m4zu
NmYAUZIFajFPX3uwt78UNFD21xLVXcfHVh6o8HjMb8/IlyJAVly+Pwcm0nq8YrOv
rFhI7YmlT2gO4plfBKWI8dnIcBJnnYeESSysrv13vIMeMt1uZQOiOp0CZo+T16D5
gHGAH7IEA+Y0y+t6lS5i/y03hT3iA5fJPcxmCoTZSOZd4FG5rHN5+WFHKorWX173
OfrV/DXXK2LFtrqpbclF7aau1KZhifJqXTHnYFmHdALlS5KhsD6P9DoVbES3cL5m
sb05GcbVSswDIebaVp+ENS2V1BdhP5cLm/MZooN/OeETtOhiOhqsVZreGGt1n1Da
FrQihAGLEX4r3rP344zPJWlmwWQv3wrj0J8mAkXjagB3fKnmgIWw1/Sffnw0dYFE
Hmv7cN1mcQmiF+Opq4p5G08jhmOCXxDyoXL9DJCItBG82dgIXUB3/Zl1IMCNSZvo
m593pfbxYlRHgZI9bReTbSS8rlelBwXeav6xeTMwuCLfFxCnNvncEeWJLrkX5rEQ
DSqVlaUTI5tnbZNSc/FH7dDUNjxuXxzX5N2t9R8V4UZVAfrO5vIZXOHoRyb2XaOK
yzcSReLU0rDvVn8bgchoOzceFhx4bzaj3NynvFuiDPetvO/ln5Mw6tyOJ6Q3+0cR
IBV3zT5KjT+nf5P3jUegnXFnopOj5sncE33ZZDIukXhS+keQBSEFzKZe23x0WfL0
VWBlXa+dYzyJvh22N52VeH1LsNdboWXCoCPm8q5Q33kS/T4Is62kBbvKSdWmH6E/
ZTI6RCL5i150VkjRIeKUETwq6tQGiZjW+gKZqHmAuooj/qSAe6h9AM+RT0WSkxzF
t311DKowz2v6PXmduYmUXVNT2jnuFDG/fLgC7ZX+q/qcZhLoy2sdChkP+pwyVwxW
grUIgxNxmZ6zP270Rz16VHAllf6JY6iENMw4dsZSuJaLjh5jBeNzf8Gsxk0dj55A
vmmaLWc97k1Grc2IWeWtXf8uBsCE6/vB8Vn4OVMDJk4LgzaX3ZQpjChMRotPDXJb
HiudGq3KrrRgc81V52/4c19pkM8YBSXUKAM+kTboCRNEzNHcDDbpofJcIJPk49/S
qVTrm66p84fMfjLr1DghkEqPnyjwjF6WteCSpKOaaxjP2bE0XHkSL0QyjWrs+Xei
PwaYnayFlXOM0fAnavpAixX4Y1DkNVeIVq6s5wcf4vAQoNYkT2+qZp7xVNrUp7EB
SkUldxr1JyDrJAW5PTKwFPnibPfKqZAQZRHL5lOqRTfaEAPGZQp5gy/2YSWToBST
VPZ4k4CjgShHlqoL+V4KlzJzaVnPsFTlq3gbW6KJDHsgMAriSaQD3hdlM18sBYvi
4DVHSrWz10+CslMmdIESVPfWhURftfe7oNVWVfCXNJTIQ3DA+sxnbFs+3oMxyOtt
g5yCqB0QZSfdJj7EkMzdHKR7r/Zz8Xf6iNwqnoL/2W+CSwXvXDVLdy58a5jdJpyg
QmFmPofYUfjl/70MIBNUNs4KshaUd+gA5kXLKGJ0Y2/Ud669eHDYwtTBugD4hbmj
ByFAtr5dN1oeyQ7Bipft4ZRePTqJoZc7ztgsOPdWgHdjQVe8jIOnRx2Z0YHSauOS
tBtBiUm0A/wD3rdXJgcDoDg3WfWJb/9zVkAxgeSaRT8n1y5aEizHsz+DLbRUnhFe
vxC56gCVp6hlhnleVUtdRBB/ksnohBDG6GQKcIuIG5Sl92HAoKTyCvMcpHMRlSPB
CA2JnG5WOVdxjlohD15sIZTBDvD05SwDjRWMNx01H88gUIG74nIvu38PwE4g9PTY
suNP9eOsMxBG6O5F0aTbzm5/b5zjpAqFGIbXDSWbyZ4YpXr+RJVVLcyHgikxjaoL
4APRAZlFTtltpbGUBZqP59/rpFkEjtxCqwIZQUJyse8jYPXgcyLBvarW3sQluyY0
gGiEpbVjEpSgEtVg10/vAvcANMvBcNFWjox/NikIkOaUKWNVIbnbEovMo2WzX946
VVsDyDLpVnB0PLvSQQVFP369czmzZRl4pXqHzwPNgI61jP49EEHxGljBC2x5vLNf
9WC+dN19Rfu2HELI82GXXKRQMNc/lQB7zVPRN7sxvXjvFSSs/rd/iU7wew7QUERG
zGnlwMbdk6XAyRWmDzFENStQl54QzLs1UBLS0FkHCuJEifB4XWhXpbweRkH+62k0
OnnIQ2A5sB2FFoO7N+sPoGROy1LkvNrAk/O98cWVYQafsQa4Woz0+r9iMy7I85zx
jycfH/FkNvMC7P35GYoRmERBiqx0L0K9G5P7PmNo6ExmQnnMYBGTX9EOumpkBoFh
jjaBYO8LEm5rT3/KoB8iRWyce8iWz5sKY4biUxhEJ9JxjBSwhJovejbs99KPRJqD
IvZmBjsPamUdy+3Xr9xB93tG7Ft2pQZJdsEU4VErqg40y6LW3f553ua/HiLRUHrW
HNGjPMxjqpz88v1SHY7zLKzNtJgN0FGkMnzZhBr9N+qpAD5taa5c7os2LniGiSgB
OFy0k7F6VrJ1Rk4XKVCJvBX3ZY1hEsYLrhxdWFmT9LE798R/rvruXObxonzH1BJZ
LXQDENkRCnZ4HCmGkuckgHN0s2kK6Oyf8i0MWcECN1+rZUPlSm72POJu+/5lJMik
SnnIqB7ejKeu+IfwQunCfvyr+dROHNxFlC8pKm+c6WuHDae2JxckOmiDUPIXyoFl
27LyghHQCl1RaYa85bnqpPfTG7BkSwnuH1+5cF+HlF5XwVA/vFcnKzk7v3ppTfaz
TXPQ4Ovmq8OrbEFZ7TfI3wwLqyqo4gC825ld1s+EpNKSEqAUkgFgJP2qC6wDW0ll
WBLeWXsiJow2M5GS6r6F+ex/yNYVYBK1Li5j6d0VcTcFhu/KqB6jjflzYdtzGP+f
11aehFL9fNvWemQvgK5V3FArUkwN4TLf/ojcGiQWixZQXlmZ9HYstLkHbXSw1vlW
cMsLbhBrvSVBsMjkXq2mk0iRd5/cEG+l/+1nf0xPSnqQNGkNN+7pOMOfzVnZB0CZ
3HCBYfdSjnQ7R9CLmOluib6huLLTPmXO0E+Bi1imru/BHoVv8enFBbyXcFtMQHaN
YFzn3ykxdppSHqwvw/aBTU7e35umuZMGdpoaIYr+cVoooWBRYUA47IFYQn3ewYIW
A2fadb4Z0/X6m9kGqSpkYetaQpDVOkFJJWxqdv45rMkZuftIZ0efIgl5h4DdpQtR
8LtpIx+240LoY2vKVlPkKVIwx8NlQcf9q0q2BogOBUR/deDs8HdrBY53NFAvChxQ
6plSbd1gK8SLkMatIA1d3Ye9LO8gXjX93/JEx8/YK6JtZFp4Dq7Qkc4/7sEwf4c7
xxlbBFkMW78/mR8Blq4ORJLdHjVuiZfbAFR0T/DAganVU6FoZ71smjjsdBC3i+jj
cwqMAKJWhzBAIqzbzW4ZmI2MC3l4o7LiCOzHyv1Iq/Vd+kH7qdpsiU5whUc3NTUI
sBVW7ENaJtKC4EbG6yWmLTffcA/3lp4sUQSSPG/lzDSoYvpFUXBkGugtIaCNGQW6
XyHM3M4CgXHaUoJbb/mNajODyIvbyY9Ed3ySAHsPCQhynJCKQD1neFB+QwJmlz9K
qyibHSFVK8rh1/qzmQw10oz1D9uq9KXWmUb6LEU8pZy34YcIxfm5bWicNN84CWae
B+51O4aw03shUbWA3roafLWlUZ6QpA9feVccIrk2vLXtZi14k9RoliOlA5MMGach
V67sNHOjCHY5TUCQEGdRrXnZcPbUi+JhsOCEk3+pwEThavMbakPj2cjxvDiGeAYU
rfSetNqx6iFYtS6Qu7qgWjuyvr4RQsPs6Y5p4o4iwVm0TrFd5LWwpqX8YPCSmF4e
dHPVYPNdIuvsIZWGSqenBahAQxjz1kI/2Otix6tyVl7nK9gDKJZSt40B06eEHlno
MkXn1ERhkpOV7lYAReLuTYjYCrw1doMHECxKfR77hHd52o79yVVJfk+1ZE71MRL+
8VqogiAuUMPP47JxSVcSoKkxMXT/0oyXC+W5bUOaD0xhgkr3X1sneU2kiBDWQ4TG
CHV6X/1G5p7EoxmI7VHvxURKd7Wha+2GFOnrYqQUBNS1L19/IXbPjQvVz1BuUsoq
47+Brlp63wthD95cN53xoEUtb/0uyW7hQ9sqRGrpwjKJDq2bS4APGweCb0DeKgbA
0gUcNR+/6cpk21e0ulhsyAH/Hj7Msri1033yML9wlZhrIgRyh807w4SpAE4V19Y3
kwdQK7Dwu5ER8Pu0FBZ1P3csv9+fDrSh6hYU11XYclFwkfm4IqlJfJF1WfiuND4q
hlb14W/5EQrkccGwhn4ZDkccNSnHEFNwNjuuEtOK4/9q+JLjnXi5HgtD00AX3Gdh
6CASdoZDf92cmG0h9IytkhPtw0wxz1auU2zbgETL5oKQWdokuoaDb/5a84bI6Y7c
RdUCHOMkjZo8pvPSKmPlwhphQfjBtFcMREdf6luqrchsCwhmnS2oRzOJmwo4QBog
mgigq1jmLubnUBJNOj0upQXsKgpxJ0GiDT6Tn84akz9czRZPx3+poPyCrbS2leIv
uT6X+WiDsYi+uiREGAty5dplEZxtgyjoXXUGks5NdXwZ1JzSKAV5mHhNopegKbuf
WdY00l2NbgowmzmhKc+gjZ2YyOOirfk3g9v0NdxTIlkjLl+lE6ItSBKoX5OVFUmG
q9imynkdfiqjc3wcM1nm3A31Tm/xvf3xUCn+SW8WDlfbAFpCEXZtY1EgwKczUxwI
d+KsZ1WQbNbwRltRTeguiZ2DfSZ+sEqlCJ9pMp0C0JO+5JHjWvlwiUuEzpW/QwEr
TbMuTopr0Zj14KLBv7g/ZMMJSFkjp5N8BlHgezsXJpb+zlCgPg3epDi5BzkBgt2D
KFVw/ISO4ZHh6UmDKLYPqRjMNCKYK9z4lsbe5gBkNfBd9pOP+pX4OOHIx2efjOp2
RPMfkyD+PbFseGNL4fufXD98UVbRYtDcyJjO2GvGFdsIr8SJY/TVSysc0fOfgnjr
Je3tv1g0zU4aD06xWRugnYulmUZJIk/QFnjV0Mto33fVk6pS0ClaEAWmYYIhfT8g
QINCKUHZKfWK99p8+WjGc0FwT8uUkRmOU0dPp/NBxN5hW4qkaqyY8pED5GvyKzzs
FqKPf7iBf6KQIFQLkj7FAhQ0SQdRREgHiDuLQLdCKzhl1niI/sBA8llqO/nBpCFB
A8KN+USo1JgZfCKXGvQOZq0yubHUXwOgaCWtA6m2ud3i31BpShbZBlAjcjA9XHZ5
6KMchtucRZN3VN6lCr1vuEjEqFSCzRvAqzwHmBws2rlbD0PwqdyC1qyVaqfyd/7U
GiHJQ6yUiYveW+/EQT75qAQ+gD4xKUuIVQX++QKmTgS7EPZZeMDqzedLciJ2/CeG
34FqTS/GT1oLjGWE/3QjuRuAOo6YAyIwi/abi6etQtmo4LkyWOYpoXyvilRyl4gy
w6fdj3Y0XKDKz2wKqQpdEV/ldxorq27C4ptJMqxH9+/uINKvwsSQytvzSNm2ZSyA
TD2NeWUV+LLaZ+VCFS5e03I/RaWO3EIrlu5iHncyhZgZJBINTLxgTIEVej4TZiiV
x2Y0MJZeTHbJ64DdpEPCsBD7ouRSeHeu3UijFgYU6cJNJnyTYF35+8nOARlSbP6K
+3L3kKZTzn2971JVS9Gsj6B7WVnGqIpeiOgPysZdpff/aP7v05KxNMuZM6w3p4RS
0BvAckCXRWdrT86isrUFeV591TlN8/+stnElAHwv+EKQX/d/3X2q0y/sDOfgAxeS
LPywvFD5kW+vwbbKc7UFWm895Ppfe3RJNshiMsAgG/IQzwTHoj3RNnFCjuNkOXpX
h7Slm9C+P5KM2e4Dws2Tc58qEAJA43WkWThmNRfrvlDY7pxf76qpLXBs4L2k0sTD
Z3TLY7j2pd0kHQwrMymiBogKNwC7TN8Qcgf6+mk9SkBC2wYqFUgRi6Gro0Eh51DH
ecJ5bzuBsPRhyjvOLkVr0vXl0V2S4uj6vpsjwzUS7ZGh3bX51lpTQ9AAjTmSpODr
3GlNJcR1NrADKZrjpWJE/QSpPZn0yaJFIU4PgA1HwizuMh2k1kcbJH8wmG7mMBGY
UcdOO6aW1HS+o258u6YTc7dkHcyP//nJfMwq2tOEb4MVN0FUSKOpSqOjo/8Tfva8
CpESaFIXgNaEhcmGcSaXmRG+8KchINHZJ4LRdmXbPKKF9Kd8NyRXS+g/M5xKNNwe
oibXD23NBtW2YF9c75cynWBBFWujwNCIjl8Kqn1p9x2SOpsH3f5pO0CE6sevoG18
S4TVns+kzqYsSQvR5EblhBhmNEgaEo/G9KXTrBJEq2t26DGLGPcKgtXDB9w1Q9ux
vVQ/BbmM45KgHAXqOcQ1FjhGMWLz0uYPx6vIq/HQDmohxk64bSwf+mCtDAi6ne+2
IAV+XZQG39bnDheo9jeLvdA3qwYXjQzASussB5jJN2Yn7BMfRMllQxo8K/3mJkXC
kb/xXv/MlVb5gGFmuZdtIdRrOYs8C5g7IDXGeuD6GaonxUhHzRGS8FKJ2U++AFT3
UiJrWMfYGmllkBCMxYXRzcbC9sU/ng12NB2GDl2mmZQlFNW9Y2IuhYHW+AalXsrA
0z3iUo0wlc4RY83n4D9zFvYL0BPa8xGuNRITUHOR93boPxA/3sNVuBRgt9Wtl6rD
YfG0Rc5hKnb6MqA5lS8zgYpVM1ur7yHaR2if6uv+HutbyhyCsJbkQ3Y2OLp/YQE6
R4r44FgvSp205s4A2BGjKhhYO4dv36ZZAG+KW303gUoZwURT0fG83yhsUAtpVWfz
vAbaiuCu32pv0aGAmZHnjclig7zGgJgfqx9vx/U+XA9sylSfQXpRysMTCRZYdKir
fW6xVRxs02nNqAElvT29WqdsZ+x0lkahs/TEQgTkWT3QzcJ6lYsi80MwMWfhRNh/
al2K2cznr9bOWQy6aW29h3mIuReKeRq8wxFrGyQO0SWBtQO9vY61dlI/j0yBrAbg
ztHygEMSXwrM05EZTS0KvTzSVcRdvbYvNAGfsAPYqjmRMOS/wVoKBuhzTNTq3FV0
5a+Idx20yskz7bA7C0BBn/izswW7iN2JUcLee+wO+s7yoocrDOl/hIHUKCHY6ae7
49Z9SVtWoZvMFzmxad8IxqVU7PxJ45s6Asl+b0BSelJxl7CiKwK2wp8BWFyfAEMi
63BQNc7AigRP3i5x3omnGRN2aZ4yG9L6ME814X93vP/6WaWHdvE1UZmzPo7uuNTU
nRO7IHiLEjgS8S85uR1ZomXPN1yuiD2E4Iaua210X7LfVXBJHln9Ryay4R6mpp8B
kjJrAAX1bp8a8ujz0lWwufk7B0w4MgxcteMpLV+Rp/bm3aQuWGsNdhos9ygHuoTg
BYFhg0CE4Bzzfx+wVm9omPssao6ab45dp2B/QproWSa61tV4/3DsZsNzY+pmLmBi
t/N0yFG1pxOE9ppYJ3My8WHAxt+xAYHp5soI6TfM5ysaIP6ZxnycMb/f9CNcDDNJ
WqSTMHGkNmHiOuVoRF3+7vbvG7I/ReB4CORvdSikxtO/JFGL1DpiYyx4e3br/vh6
g2h7AcIBWM+j3sftZNhx4wuj6Cmd9dRkgAp/8Qyr9g5YZByzG+eWQrAgwnD1xcVY
0hayAsRuccou3L5UjX+Zd3izRWXLdTziAao5liyr+htqzM1u2H46MBhxMaeUXa2M
D/Ezyj3B7omV0IkpBvEYTFhR0jyGgxqMDWfuBtCWtuWJxQ2cKXeXxuQ4qHulJz5D
wMHhQcVs2w13cU2I3HfZVadPP8+wMJoQ0vrkPN2VcEvNA95a/qSUdDCd1o9buKqn
TCNLZp9bj4LuPdeVLBMvzPKlSMV0Cink9gvzeuzsXici9oB/RBl2apTKuAn5Tt2j
LKWw3ycrebW3c9CJAEXF50hJQtU/PJFES5ATP5737/cs+dKqKi8zUG1LdFIaxDEs
ouapE83bfu+4MI6+QQPnd9e3C3xZyElM06HV33LuwadOZZqCt5e12nx6GrzrEijR
jU7BNQShGiDqHkJtnGvNmn0gUWw3GtG8bdeEUOWvDTeT2vYoqhlfb50cCGKG3vOk
+r/0CkwqGWu3N3Fj+tD+XaAVfPovCTQ9XtsK6fn706WaRF7nv0g0jQI+do7G15iT
uWSNXplVGEQh+zIY62cBr/ZQosm5Hd7XFIETR1luuG2AyHLuSuLmAkHw6g/HF8/X
28iv8KH7LG0Rfg1UmVTxj8uKjE04f8ih7NeGA+QrH7fZbXfywSbxy3steX0P0cvB
k0edj5yB7YaOXdlCtzUb/x95yRBXx+5OIXgdrwd08VPxqQzlV6dckdkJojvndBnz
BolVB7DXF0zQvqbc1jDtJlvOnC5tRSigqdR04XP+DJqpBDqoOZiBRfDYkpoMmyZZ
VsuJez7r6fXw+ymF09+R0CSWRWN3hVuCG+AuB1IE+T681/QIGc9zPziIY53fPo5U
Dtkom+Vd19Nq4sgxUElfLovj396bv8g8Dtedu8mAj510g2X59J2KpVSjIfk7ogVW
CsCdUXs0jUTKfWHNtTt/tF3lxFEpHEKpU5dTqp/XS6fKD0gKz4Q5e53fFwRaHwKg
Aa/lZdz2ahHXTx4s82BjgDHR/gtyEjQQmrbMqQrtJBTtCdZti/3T3krYLqdfY9B7
vYlUNq6D1YChuc1cdBxoIu9hzBgbG4pkxpkGdBuDdPY6XGfwQcSDgSD7eOxC6D2D
mRFm/HgKEffWkO7XDgf3YbWac84iCScJAYyuc75dtW5yl6yxCTMYhV82fxS71GO5
g4QG8qBfL9Xg7qJOyvUvMSpIl+xfX4M09Y/aT77ym9FxZdLISHyqhme2vXsoZyYo
V5/5+HAL30x6OleEBjTqX4QEV3rI5Ub/XNeb8d/tCtxQ1t+mjmk7Aws6HMWWiZVc
JQ7/af+NOEYPDOwr1Z59G0RpM9LJ1CYrUDI6HVWnhKPbQyZTXWQihaBC0OmZUEGS
cVgEnDuPMRzD63ZI4qXxs1fzHUVqC35AtmiwZFnuuvXs61+btK+LDgbYaGn3UWrI
Ii+QBb5ca5xBtnq74T7VWpdrVNgh1cntizcrTL2L4fPy3WxjWksQ1KAyhMLyBk8U
5+Ak+Y3kp4a/Uf9mwseQGl6nqfxVBAhoHodzH+YAAPg16qy6sULhoIpD2DfVk414
a+0ozvT/vk5pBHVh5FieOVeTS1n+9EK7MlyHoHzszHL9nnE9ycyL4+VMBbPzSNpI
3T1s8XjYNq8jCloPRqnGTr+fvrFUP+t9R0FOhj2xtSKU3fY+kT2O1nfETi4qW26y
xvhH4Hx4wGkooRQLDQV/XMIjxE93UdER8r+HJU6iXNq2uvoGjhXkGz8eWid6YyS9
it5zL26lHnyMWeQfGNO74Q3MVzXF7aymU5xbTh6j3BsQppcqnlSQxwjzUhiHREwn
8uKlU+DJsdmHmvpMZiNhunbD6zHb/Cl8vCqse4LDWkGD+2NqrWRSGYO0ju+AYuBD
aWdZag5jynQYX2OpYyUwfW8f43dzOgtXyNLBKydpe4q+AecZJ2DYzvGoynIb+gHz
jTwO/E9xhpfLhv5AgJbpINGOym944hDwGcayS4FGVsPWHPAObgi1A6JWKNC/gT8S
oTea1U2tbLIbRbPltgCvV9kNaV9lcEROntSyQ62a49BaYbPpgq86ZAwvYkDFMktk
UdkoPEhWtRDifm34OzzVVn8Moqqm3DGNCCYAQKzjDl1vzhRMvEkl79VuWDSA8LfN
t86epyddyUtVImx1HaEz6o3slW03/ciKnJKlSqJeJxDqB5TACqUHzaZEcfg9GQ5D
Y3Ju9E00Hl5Sk6IPqbc9Tw4O1m/gMF5oryndhYyuiZd9LiQFip9CHi2uG8ZLxmBr
Tgc8Z5WLkUHv4BNAgmX2oJ1s7G+DUEF8ceuFqe9GnDT+/qkhigRt0N/lg5AqIqq7
oTBysMRE8deZ6zx28meDIVKw+Nirl1MFCvGiXFZe+3WTREkGiCg2mmHc0f65aAfW
aqzUVf2achF7UnA3Kl73IzMtj/OXDmiSlNBRcl8H9A2UY6gLRa54jYJos7vGbEAL
q5lEVVSLsYMu2PSZAiwIdtHOFJSTxqXyWTPX6Smoac5xN6lpP0v+lPA3gr0ggYt0
rywDho42Uj7fC401uhUq+/nwbnpP371E4Nx7KjWbG805KwCz3DvT71OSbI4XYpu3
D631b5uRwYJVYNXkwQFcZQRaCqsyph3jbtTklD3+wg682mB/RCGEu3gFD/OMxNMp
fyrewOwccRIm99Mf8UKZuE0nQQEj/KS2qkgExZAwqPa5nIkT91HSSj/LMs70rGyh
i41SW1B2N2FeyD7HjyoLdna/8/TeHFZ0n+mvs28mByJP0CxRjbuUZ5b37iVcRkU9
CKlYRK+2o5WAkE+V+wEYzrTfz/Mk3J5HSo8Q0vay138sP1rqLH5dj7AVXgDndG1R
koKwcYpC6Tcm+wKE3o1iuv2mDvQRQTnfJbleLmXGIHuuj2MVguBWnMoEmEasf992
w7YjFU85f+3gJ14NSC1bIQpOFY3Dh1ilpfvctm/SorINI9m5i84QewCqOIDy9eNS
rl+b5mLoUx+DDTiWCl1S8huNXC6dVkJ30MF84M/buAzaIL7B1//Ug6Bfy0LgWQkY
60rcXhnHDMiIWIFEfYIoeK8wxvk8ymteZN83E8//hqbP1d4+NVsBFZvSn0aJPUqO
Uxnm79b/GCSxNwaBkDr5Lg2pY9NKTkcYM4lP8H1/RyKACtcewR684/3IQ7CZxpN4
F34YQC9FJYvgHVUQypslQWIxH64srhUSQ2zTW+wUASNwhhvx1EsOVrp/8i+dgqTF
Tb/m4wBqvEKMG+LTEJzial3nvPqcAqpslgx0scuraLT4oQPvBm+f0zltRzGv+m5R
mxAOlwONsDswVnz7yYHs3f7TDjJxQRQo8EXvUT8u+RCruh7WpAu40/2uNdk3YxTe
GcrqhPGtCs8lssltPIdfuS8yRu3Zu4GyAMIvckaXhIy1pmH19Mf+RQ6Uv0utk2Aa
N/Y0A4NeCB/3Aa2LmxyStOshS62mrjejzjYpSIhG+aCrY9RSbAR4rEJj9iB/DCqy
yk/vj1K1DtTbFVi5TkO+5Squsq7Y3lzozi1H9PCcsTnKcGZjMleCgJNI9IilRfa5
jLQ/wne6Q5E/n4a+OsORUFeLN0k6C27ssW/IHRVA0N5vnZZ8L576si/FuX0FGOYA
EU4+duC7y3sJ0ZAdQx3xJIpXF4orDQCDFXlsKs7hwxuLEc1MENEDyCNORic3wDCo
O9zJSiBxbdH9Zst2zYDpkPoVGLu3zIsuVF+J/MDpLbwDjCCRi8Ti9ld7DtbEXaKz
EDEfbXnzX+Bkc3yX8XfbpqWIixySuJtc1WNim0IXJu9ya0BVlN89ml2DXQrgK3jH
amMvmEQKXU2kXynkMSmnnqm4ukDh+63OOqzOvfvSI3iwhwC0Pu4i60o29RAFfKU0
LpWWuQp8m4fTjuNDfBSBseus89z24uXBOopyd6DNP0bgMDHgYRLfV+ttLqI3oO5X
R7ClZ4ysFiLsl2TTu5o9th9oo3HbP3QlVE2kYjhmsHPss+y+xko9KS4qIIPKqSsN
on3Tuqm61HzENuS1EKdYpceYBogVoGBO+WqLgCUENGYnHG2EutvAn128XWxMDXEZ
ThMOOuBpfE6XLh989uuwFDy+fOmPNcTDwfcBn7uITu62bqwxhGelnT8oYj1tgh8B
O0bT5pJM2UEX1eRzsmCS4mb1399iz6jN+Pqnajrq8ndDQ8Qh6e6DopXly77Gquun
5A09WNggWxlc9ogvgd3Dde3MzpzaJ90EPx7ztol+t2Ve+Fq5Hry1//4ggraI1F9h
wkWViDA8Mis4qlJgNFvSx0rSWJdd8Ac5opQBT75/rbMdqA0JSquGSFhHFt9q06zl
Z8dtGjAO0hw059ebUTLgi5ghpiVwdDqeeNWns1Df7iGsELGmGwhh1ovNrNVnNri+
kiidaxpftc4A9pj97UVtkqHhIhd83/4J4sOCZApaPN9YdHcJ4ftw7i/pp4DNCxzt
eSNoENWRlrAVXbrWOrsr2rnXNMGWbkcpecfLLoAG/RiiMki4vAYTMS3aoTDVXgTV
ufmIhY8ks1wrIFpECmRvZKleEXKZaLTTTdqfxYuxOC6wbXAisEtvBA5Ean8vNKzK
Rj+D36wjUvgtD/Ob4nHXFFGoVmGNT+hHFRjBjtAgsBJy6UbD3EN9TUa/+rmdIwBN
VjF/5Jk4p0XiB6CAlLMit/eOKxBHsRMsykGQ4B8AvhIrf1BUzaXvPIpbI3GDLzlW
TGrOfS7T8R5he+eSotf5ln/ed4GthkaZjoN7wQByT2sfY3rOtSV2Uo3ObghL6W9B
NbyoOC7DJNdujgI4yydwYkGrBcDQjqyKGVD92Sv6oHYpjGGYIaJbDnM4TkDixrjZ
hh91mfqaSZE2yB6aJWZi6iJxNWJrvh0VIKA+Imsxg1ha9mnCxBgE8GE+6LVRkBNo
rESx3U0YAhJoh3nR9GalTqcon5N1EcSchpIBfRDDcWaPRUHDEIP/ecG2NiHExQJ1
MTHIKhZ8v5F2tmQSHgiQyUEmdEMTpzwtrNhB5lo1sngQpyy2K5LutsuuvAs9Ynun
39er68NLWxcKeYr4O6QElQHJZaK2pKoLfHqRfwg34b/FDVTOajpi0ieZ62zr1osE
+Mc9sJicTqeQK2iIDylUAVO3QuXqBY+++5vUKffEC7Ltz7SgYOvF8xGu1boxqi4s
/NgQuzTm2M28IPl7j0jPsew+0UsuQIhe2v4rtlBRgr+PwQds+bd4RAqZA1nXkf8c
9kCkWcQq8AOd5dqdMtfRD3eIHhlJUuDN89tFBrZhuzCrhN9BxaIorcNF/Gji+Q4E
O7w0kVc3hzXV1bmRTCYNk/BkiDYE6SEoJsMCl4imNsB94QfIjLjxdqt+z+E9zJb+
Zwld0Hbu7oLSYm2j7VZlkBNSOJ62SetRrvuaICBCnrAtTXXicNRDLtmh5gTAJu7H
0gEgK05x4FQcAnoVTdGMpEg9pUKom01pzQFDcEoT3gr6KfAGTKH6dvScAT3AiDfs
sSWXX4BnAlEHj676LTqqphcHop8tCm8N6+V67Drsy5yRd8HvEvD3mhKdsOZQjrC9
J4LlGncL5QSOLVwECXr46CRNjXi7NHTBh5GB1JjJVlEjCHeoJanN5041jyjmkKXf
R2rxcmyaNnUKsDuGUAB38sRgGdkvZcIXNkH35Y3CjvpcZ69ffOjMbhpUrp7kqrjK
ccpkDjyyEaivd0azDqWw6/wQX9SawYDgcT4DmZTw971LTV8l/2Ve9KHYvcGTSr0L
bJ7NLOdkE7PH9PZGZjZLM/H1Jv+EzcyydGS1ur9EarDTdB/FfVyasLZVvVQqAhB7
w5k1ZugePTjeZ3oBHadoWOhkXQbQ/rl6YQJjdhHqkJYUPrY+zm3cZMdiE8yWNNEF
wo3Bs/mZ5iQsUTRh6Vmh8hHDfdkyZFJblLq/jfYl+SRijgiVtyAX2pOxG8yzKzcv
PMaeNsLZxNf5+RYncK0qFBpy0zS4iLqLykrgOp3N/m3U7FuFR5dQvx49sVGqGN5N
roen8RfU12XVwZsjw6T+H8sSGJNS7+Qb+Rcw3kfQ5/aZz0JodG3FbQ2TII1gU5m3
oUBhIf1RLPOCsvk/IBIPueoDbCO1HVaLYUF2pYy5ET6yJA9swjCEWvCFq2cpKwEg
ltApg8KEyZY4G79oJbFjevK2OJmRcmdNoZzDjNCW1anQzo/h0kF6b+zgMhlgqSnX
kLoLBs275+zgF5VHfHnd17oHJ3xwF3rfRM7lkhS2K6A81yGeBBun7DGQuQ5LAoa2
bGNYcdvinid+jrIGMKUPUGD00P6ayYrSOzaswUNuNwmtrq1/kbsVzDqughdr9E/X
Rg6Im1aRGD0NWZmUFurkY5emaDuIF20mL2FH+j7k5VOqy17FYeY+OgtTiWTF7+BH
o9WwC6dUcCjuuE7uBfCont8jUd9PKsdm88A5tvNdAqL+fG5eR0DRYBrfx6dFsD0x
dh2iPeAlo8OuuscIfSNhhOz4XiJk3jtqd6xFdSjbXdWahbZclh+royqJ7GDaiKYk
McFp+FPf0dGWvoU0yRbziOCKvCx0PnSm7Mbv/I8yiRaSoFvfD8dCPJ75XWq6GE8+
IK/bL1TXgh4ELQybVMzMhSrFmW0IoJuhhz+jiY1+cA12CxdfcQbNBVWwaZ1XDtvv
H6h6VvVtQhf2MJ/8re1sWd9km2sFIRrnuKmupq51VxoZ90JrNMQx4gR1P9twQvc2
9rm7Z6uHgMVLBMUjbWQmmyrtzqHH2IyjLej8FxJQOcDWpGR2TP18dwrXLUUawrZ+
hXwUw9Auha+QrX42R6j5GM6hS1hfUs0BMbvKTKxQtrxLcEGcDebRm4cS5M6IgYVJ
t+aFUx6JqtE4CA6l2ig7waEJ1VKPpsu9uKPJ2eqcGwa5GeNr0ZOz42YF+Y7IiBsr
80iAzTmY8mZGMDQcqjupoD32tr6gPPjvBa/zgsow1x/LtF19FWe0cb2fHuTBYOQM
ZhmXdxNV45BU+gkr1+N5pu9GyzbYjpLRa0FI7VzaYRTVIRhHeJL6JO2jmQPdzsJI
32rTGr11I229Kkkh99sRsBX7Van5mLx/DZ0yMYG9BtcxTL5h4J2+Y5qrXXPuMzHw
Heg4FztC90iUq+NzJd8dZjEE4vUkhhas0FSpQZrh/t/Nc8oFqnSB4CWFP9EF/qrD
Sjza/rsGLXn/d/gEzSgjrCIomd6KE/cMKYctWbzUr2dggaRF7TmNv9BCz94tOQrM
WAMXgXjApTzny4vN92VJPKhJaRAHc8PHR0AUzpujLbtPomFM3ce7UGa4KRl5VHNz
hsU0Hgvsx/WOFH+TXrUAJFHQTvuOFhN0QoBREDgrWn38BCBCSUDpQ0WBVU/Al/C0
lQQUcztxaGwbX/6CbMsqt6R98MzTyM2iGLIEekCkhMG3E5WfZtS5AEtXUZ6RMPej
schoGpu7swYmlxo+XBj1wGxbR27UM3xBQwXKmJUR15Hh8+OGf8CsG0aCpl1s6eiP
nykAEwqBqWiKPdFu+JPQFbSguI34OmwaRu2atE66smv8wAtE56Ljg1Q9e3cxFDKv
+hXjxZ1S6BNeve4roBWdRaggO+5ZESe4ff+rfbUAAgvMPG8psAHvfhYTT9ImjzrW
ygTzxyhD/ae8RkkuLt+XawsI0xeuPqZDENqQgVA9xqu+YZ72xnrgZfYUAxtP4KMc
TwanH59Vv1q/v+wxe4QBh3YsmP9uQTT+TKP3hh1IGUo0J6JbooTS4ndrLbgjFoCJ
zh7xlgeGJKMk764uYkQ6byAAOqXdouuUSksoFwFV1s5ZpRXu4QnPK26zRafAviPd
5NqIYF9V3CMsWV/UBy5MS70QnhvCfr0DA274fVB2EKDXnP5Z7zG1fpTZJKwbJZp9
Bjdrt7uw3yscxO+AcUipdYNWbjH6dBL6i3njisowPdC+/Ae5QqC/nHF/2VT7ferp
C5/xNZ2gnBPNfdMYUYSzZjcOrQccR2Ul6Rj33kcKjmJo9Ju1BxwCWcqCQCX2zmaS
+BRS2Nr2Cgb0f22eluvCWGHYoyJ9P+Iqzq/m3IvtF69oYmIloQvb0YeOqY34egkX
CBahttJWVbIZtcNPfLZLOF3zhcZPXbcB4GrpBZwSX0U6SKHiwNiIk8GdsldSySNI
KndPrazrfsJldDFY+cP/M0UaYH827VEnUXkY54DS04XXL2zIcD1bia7npaTmUDW4
a3BBOF+n8ZHyd7GA/2FomHTN77rNyFQA8hlLp1JfRZqGR4QjZFF9vVtjbUVtGhb+
kVVC62922MW07qPVPxND/l6LpqYM9R8/OdrMNJhqddOkO+QOB6qqMxBYvN7JnI7Z
AHFZv5GVhY7hBJjSeOvrBM5qadBOuHhSmP9lm0yAGX6AkUmKHDa5gmMYJ8DqkPsr
ZqZMV56Dueyugq62yU/1URb8jdSBHTiQ+vc4Jq/3h8S+ZD1GCcexEvwai5uZagxd
gCTzv/VtgWSvsCD0z51x5qHTC8LFKm2yBOylTqBBF1iRIZtX/8NUe3qwt+6KoLaf
Tj1B/DF6X1SdDZUAglRPk/OSxFtmbVSVcGfDdmDs/GGwHu94hheknxYJy43tIBkf
TemKExE7JHX6OE51kzSn90+S1j6yFag4CRoJXtxG9o4D570vqxIph+Di0scH0xzg
0kgGxHwdsPoNWN/VMu326RJjPWQAiPuEd4UfZPfNUmF0nh91UuJMeoxNed8j/IzB
+INn68/fVqDRchYOYmMWXcjqB6Fv2/tLggC7BLbotbD/QxAfr2ZLmtj2zJ8CtOk+
SjlmpyllTpXVD/PgjofeEfshK8pbpmWO4aXgxcaXjfW52FMIV1m2h1ubu9dDItC9
lw9n3nfeef3KBZSpcC94xRvpzVHM5OU/GMtBiI7Jd1fpvEGapvnuC6Rv44fEs/l/
sio9of1SEHQ/v6JPnL9slSCGCSVEZ9MX4F49/lT7y2G5yRZp4XQl7Fs9fkbt0ZvM
Oxz+NhvwY+14UcriK7wEKSD/fFbAErk8XZYiswUtknTSfh7JT2AIwTqVnG1Fj4G4
Tkfh3FGTjwhnTV+YYjEOSuX7iaBFxTEledphsd3hsvIW6o344uuIg5r0imFKMAIw
wbPjC5xvl8g8KeSHHMrhdczfUePIhcPM8mf86yH3ca1ABYrh1VJhLkDID3KxyHKP
iWfo47Sj9aKo+9ok8n5DjwXBSmgZzaZwd6WxuQLpmQYPIr+zBUocyTYJRvldnV3v
DILxPCzKGPy2MUH2vPJ6A5ZzJj1Cljok0i440l/8JQUslvH0ZG2qIYVPFxueRqez
VJ+2SCHMzXHiH3ijMiKAWVuJdDQ2eJ1VldPb/veMnt8wXdnjsQZvPQ/mTLmvKBxT
qdOVtMKR78X4MSwVeoZ0Cblxrj6uqypW1y+z7dB2/IuEBv1shQ5JxSHQmvbSCRBQ
sp8y/gL161qlcdICySVBs5hsybHbx0xjMy5fDOWQYiWghLH+lZ9aF3+y45l7gJp3
VHsiXtk7EY4nUBiHjE92Ls1ktCZNBbJGDZGpaVq1xFMXYgX/DS8R/ZBJdslrBoML
h7rgHuuOvxNCo07uKpK+e5Pl86CaN08fvrTnQl5BuHFTXzMxmvlgeMi6k6I9Bk3+
dYLgDKT3FzgDBtnbM9RKDtNM3+53DV6R3Kt4KWrIYxy51ngRWVCqXmbFppgAzPaJ
UVnXdDPwYulpTW0AkGOC/sEUvWd3Lg2tZTr3DZtdUpAGmnUeGbeGxnakNrP+uaaC
e9M6YpsDzdki4ZF6RWE1q4Aa14vicoIs0L1LBDelDxZIFtRaNvslscPml0Dn+m8S
GsL0etz2rAIeFGTCmOOthJJ3w7xQweYWfa380AE15MWDIo+7jhamt9Na5DM11vPZ
3gpr+/eA1tBLkG+WuLV4G51O/SOgD2mfgpRJe5fPX3qLzVObHRkdQVlvwcrWmn+z
oa4Uh2zsUjXMakyz+nj/1DDvE8RUiI1d9hjf+53NI6XolJmP9ulS8MUxLzHWB9hM
Ysh8EM38zfIj53Nm9+jugYwmkYpf7izvPi0aYz/AJyWgmOZeztE3AiEUFZnKtZjv
4KGuhSyaTDzXQSToPPY6+dLqSK260UGavyxBMChugZM/P51RHeuEzyF77tZM1iW/
Fuoj1/eyfcSpJoZSvWiUX+2hC76wRB2Aj7eOqIiCCjmqKXgtgDd4hQq3ZJXiJPBK
cQgp39LFRBhIV3yz+bkWVilfDOFX7/HWeRqbMiXNQKYUyl3jhJGiVmUTwCA8siIW
pYbVR/FIAr8hohd+2XRzzN6mu3FHOUNIcZjdxRTswH19niFyyUM/s5Ly6U7miHTk
mWfFoRSXRn78b/94/0SceJE4LwsQCKA7ZBfEViBiB3pW7SzPqkjet/FqXJkDjsGr
f0ZznDZ/oRKpDrA91lWQNQ08o05mqJbu4RSAq6zkPOkozC0heWCkJ1DloED5l+XU
Hr5Dv8SjLhhwr0MRwzD2g8NgkDDU3X8CZgnIC3+mlUW85utfIimom6zr6kMyL1qt
PIu8eS7/76FsHwoXFJ+1tzdC5/z0lYziKCEui3vDT6rdf9A1FmiZbQhzY/cEFUu1
rhLLwYc0k04eRScyPqZHzabrabOiAy2DwhLdxf7e7sYhPNe4FIfND3adLSzgutCF
1ZzAXmFzxC2U56NIMsc6pN9wAFz5mh8/2DW94KYlLBqVrjUImHoiwJQ7Iu7hmFn8
QM4J5M9w1Ls2N6i27Hkc0sJponGS5OHR0mYx4Rk9h0L0Cr8fbICCTIi9hHK10zko
TEgpq6+OJwb2YLqT99tILqEzmAn2Cu+Zb7uyAzxBdOGUID6yOPPZq6RyLWHC6c1s
R3w+PlOlagJDf/NqQvrMhs5ONB/vqmvxbe93b41kO4p7P9WHaUUvA95J6nkHQdI8
0PhnsJ/kluU9Qm5uuhylER/2JCypt/CxXdg+euH4BAX6QgKfHZG2EYh87o6TuyZv
zk9zx4/ut+r+RM1TizLmgMHv4vUANxkphXvqsXP1YJUouRnxjsd2wkvtfLXuNJuU
stIISajGNZFN9iXkarsbA8TntpH1ALlg0QKhPGZ9XlYCbk55crUHVeGM9GYg/9+9
Kpspf6sehGyj2+ayZbIGO7Xt8MXLT++9TPsbEqw1PldsNANqsQuoUFauacHrA5BF
qX4oXqWkGk+Ini0nMPoflt/AZsMHOvYa90DmpsyK5DhCeWRw/ByXQnmeiyhCOYuc
9mAGklckfMyev1mODDwSV1KiLnC+wrm9ZwNrAaa2tEBZo9vPRXpeoDISPgdNSsvh
kAxzMeFPTqx7aK8BjpT+V1UMBk/mQYqaWYsOxbZbNm9W5pWCETpAHRzS/TW109e2
Kz0me0Ln/2275aI9S2hTnZxBL8etxA3CoJ682bAxjlzx1a6b9IbB28nM+eZ5ZjfP
3Lc2hwTi6i46NfdaVEQFuua+wQEDR5LcNZ5ba7W0r/x7rtXnh19XGn/0RzAXqg22
P6/ns/GVXS0CYhglqJZNmDBrNAMiYHrxguxPBljd9/jyDNdq4SN3Zzk3Yd/QFS5K
/VSJl/5/ldlsCDN6yUVlR2Rlbf89nsIf6HE4/5kxr6enKrvP6nDxbZPxC8C9N+xO
yYj+OsIInXcFi/360c9LnxQvPSpk/6c49YrQCzPqKBJYQqtE85ypyFG7qMl5TM2/
dIV6hijNavXdWazazO2WoHkSRiaGjhVcuFQzgGr98xC9Fl8oLmjtfIikia5lxdee
S8IK92hgxE2KImASdizApgBfzQIyqZDGGCkhpMo0UYWC2Lpyj8gql59i8DXjdLii
Q9xm6IYSZOubGdryZzIBzxWHwPBocrdIIeZvtRQcw1mQCBIy7zM0SFOWLZrrOmIr
EVAccExF3jBQQo5RrrX7nYpdQZwpguZUKRcJxT7XEkpsMSOReNNNRJbq1kh7iDUn
kY2e+6M3yuaH3xwo+R2+s54gtXOiMkn8a+0Y0Iynk+3D9wxDhRPvb/t5Uuf6KGUd
WNaQoASSFFiSGnQlbnvk8uEiAkzvVcn6xfiPs6MQsCZ4dMSSiRwnOAUDm3CEvR+m
xEmfvWiaaY9JC5IPDl7GSuej/uysrYcpY0DqaUfbkLh6DJO0BE2bICGSP2TJHNZ2
CKtjm2IXnM1Pxf00/44O3Kerl8qUP334xF0+vHZNPy+1bNTpq9Iqn4KV/HmwfFXk
02NuWGX7MJp+cSLAyfipbqvVh2m6sECMfaUQFc+9HVzJ+ER4nl9hVsKfrSXPl/t/
kdasM5VTSlb+GP6vWJnnRfJiDM0dPtJv9hfpSXQzNT8oFe8h+SJHDmeIiSXFiPXk
SXTuCttnnViKdxqgx/f6N3+Aoo89A+KimZZIVlbERV6ZNYO9tWaOyWv+C7shIUI0
206YMDxcZtDAQESHPisH01CGgu1oeLd5CLUEkoQKYIegnTykJmlPQ69j1oJDq6WS
Tk1CWrtXoRifvB7ERpWoxO1m6EZ1drckR4fMQRaqu94R04RtS1kFEeAy4p6gX8ym
7oGBph8dNyuHCzUbnO6Hi9kjcW/W4vTtQnJNhU9t1pUCgPAwqhJHUYrElteTYu5h
uIshCYByMocQCeV6n2KZ9aOaabmiUgP2ksKAhe4Z85zpQVsTUBteBBSDb6MP4EOw
P4i8ek0jxeWBQMYsnH8rvgVNMkO5tMwJysOCbyxeDqj83QbeMsGjDhkVEDkcXmDk
fI1R3kPr7mqfjwMg2Qu8XNeXaHzUforxWHJDXdqm7VI1axdOZKQDvpf0TrybMKAJ
r79gI2vBVjKDMYgds/alppwBav8IkUnaldPRw1VhQu5sx2j1RypnLYPal7oOEgqC
CrOf/Xc0X6ZVigoU/TSxXBAYJ0O05X+A2XQPrSEqV7+vgiGqgbSnV+4ygeFOHjCX
MqLWLmnplBT3/Ggkblr3m/+pFMdVLrWxDrD6Xau85bUnfafcOWn3KyeG4R64qaZR
qcAgapIj3JmaJRvxvL6THrXmL2dgaaxk8VbjLLOZDKkCjTKo9Nj3HNvQCO5aE80G
9QWjCHgSjApCnaiQg3R05gClbtehbpxsQ6yvZF7NHitrorqUsMyvBKp8oDWUWhqE
Z/9axXNRbIGL5eP8pzHUTnz4gqyCI6fPYnoJ+9t2uE7OR6qlmbZ7JNdxaAf3RPZV
EjmwdvF1P/h1pa8xI7DMCBtE0mFJMKB2I1G84+bqTt5enyI4wo7I6nnEPJ5n5XM8
MskG2W1un/dSL7mypVEEpaoxvKMSdKwrYwgk2TrtwJdsY9KEqkBX2ob2zWggi9z8
d5TF2aGdzQZf3vjuAYa12ykJeSMvCb5FGdrfErkUK6kHCbr7Ce05NgVdW3US0Pm9
35kk/BZzR29mcgbyQ3PC2r34qh3p6IO/GP9zJngU+IS3mpD8sYWhFlLayLw4nc4t
CLc1yNaKG5Hwwv6PxcndkqfzA9XX9NUvezSpzHMRzZwFz/rEht/bTsQDHGTUSmKj
rJOeJHMovqTJul+Wbiieozar/wslQqNU9/irzwfKxNOErtzkd9LO7EUBntEmRpXr
zT+pTLNbVbHsN4M9sledXWa/7qF8vlGkvo2M+12vXEfyzmTpE05hfY7q/MaOIMvh
J1aLw4KfTdtlyhcADjH3vAKV/5qN6WRG6zeyXGUriKMcu5saa1KFU6WYNL9h6HdE
AaafJU986e+EFsHeuSOO9xXdsMD8YoAPqFjAAc8QeiRuVUbyjoriov/kxcejE5vT
N5LrRMaTdW+ZrcFwCUvRPkbH5mt9YrJ9e9DieXbLMkyaSBBsALGSc4TJDmxWPzW+
Xd9qLX/hXn3yIGlCaD6FNtC2CWWGFlOxOBijSyVXceQAvmgV8abPZ8EKEBXj4oyi
cAF9DAZMk0M/gNuVk3IpUdxXhc+UOvmH38S6uZXE+gE5B/XLNM/fIw5jnNrK9PO/
WkYUmlq70NiQ6kbGg8EPtCLpRFSrfP5gRk1SVIjeWWz/OgnzRWsDqSIwaNr1pjar
l+L+uhNuUzj91CSA3F4+It6E516n7xnCJ9i9hUI6Y0ZKZT1JNUNl6g/8GQyWKGe5
dLjb8R7h+J0lvJvXxbAUhVNfGuXmNXgvWemJpXnIDR1v538dCz22VKFp+dYLq4Jw
TJ3lFMr74G1y9MEGl2s3k1+K4qtuc68kg0Fmc9CX+9jyE3RVuSz0dbZ6YlxE/0Ts
yIXGfBX5iEiJmWE4HnSf4Y9m4CmAqWZJRJHm5LOTQb+Ov+2oAuMMghVRteyBkEbY
D/0/riSmVt9C2145f53ryMSPmsLsdjRusENe9txgx4SliFsBpL7xf3rYdaCwYpae
Js+a+vhnJ3j6MvoEVheKrQqILoIMmXfjWnX+tLfYfw/tNVIXmwmRe+Ic0p4PQjUf
4lVumYbn9R+NOthOHJX9KlOy7tMTeYzq61SzeNqrUPRdtIhwYN430SPU5bz5NmbA
nIvHvGNw26qc5/1iNffhGhW6GavBX3fLtfG4YC3eYQff4YcBRCPjCTXS8nAq3zi/
vXpfsYzBZQZ/0Z0Tm6A/Gv4SqXEbGGld3soq3AATg0YHGvwEJjSwMhd14hZ/1S5N
HiCCkNL0dbN9vGoA8mo1U9ImW6SCGXfw6evedW9H4Bc/WuirBzCHqNS3C9LURX89
8Q6aWmxvDhD+0F544JutedOTBPscljlhPXj8+i01MxSz6AGynb1tlJjoPTJ2j+ma
4OD2GnQMAkApTXcJa6GJNb/SFrjLW6edCV62KMOA0rVPnxu58bROKpuPjhFQBgNr
BFDfFtS5V1L5KP5ZhVTwZl1OhX4zIVx7QhBDdaAD1Xl7mIf8X5PVnLZ5EFGCNi2f
TPUl7XXN2P+V9omyDen0pru0HOopdD4VCHM6Qg0ujle7oF3L10+G5VJ73VgWdG+U
AWSsEIXpahctfa57K+8e9Fjl7cw2TmmvcWFEYA88hDVVVf/fnvJr7BMK+0gsIdEj
K+FqLflcI53mpotSK5T4/dZF3PVEaRLnGbAwOFHaJoBak+xYfTMkjMHNOsYNqAkk
PjjjlM4ktLR6p51EBoXzSONa1NjqPLHBLoawwnCqGPYev7FwP2Cr68K35KKTCY3g
9J91SBy63V2L1lKQfveQQkgSaQPD21YXO/3c2YZg/lHMbeVDciyE07Xehw8YhhLi
+hBAwAMBox/kbh4BlB40WTJx2Mt2ARIlO5v1TFg5GUPAtoqz6RWr5IK7ZJyMKCky
+6tSuDZIOcyCCkvxGxmZDQGAFczP5WihpFDDkM3o5GuT8QUyvfvf/LWaWiQaW83L
f0rvIcmEkB1FuqPdy+MVl2/2Mso8HcMdvdO4Kunm8yqZmI5AzeViL1Wf1Ug3M5Ct
HMwXQqyKXGOKZfs12MtbyHe3aBjXtivcU58pOxG+a0hXIWIFkfnv8JhkVcJYWY2M
aP+Bsq7bXZp+/yDqyRyDFvQ8BZ426WP8YYDBQkwmVO82fhFonA8Zwi0378wAGo1H
Rv7sF1zi2Xjj1wphgTlmsOoKgvequHom34yFHUHzrgaVHimLaHHjQ/XluI2Pmdiv
ucWQ0s4kjgHhZ4qeKXbFgrbH4gwnIjCTkdfWOGZQfLW9pMlH4fs0coUBJ1J1lLMp
Reoz6A+6+fJFKqf+wPz3MvcEXMEKKmCjQuxReUe51N6wSGL+G2i/3vIZJT2DtQEw
9QDxTV0tu5dkeouZbEoqK0abc/HV7JomH+tyhF35hISptTSBfeKnwWd2t9veN1GE
Hm1RKCld2HLdYl/Wtp3QDsx9WWS4G4LAMVO/Mtbij03V+BqXgqQqIMBuXbS6kifJ
37HNTQOHqm468yLVCYyOdJAu6N2IFnhtAEfdKWZp+W0h2bX4fz2gJ3k9pxN1tuYc
518AUqCQZV5taJ1ZGgQYJnYQJKOZDoDnjpTVoubp781shWg0wAW1WpXrCSOHdSvT
kSksfA4UhkdsZeWSjnS/Sr9j0q76NXLOwerul5UlfSn5oJ4WwVn04I/vjJTuHBsu
1KUW06wqdkaLZL/Yt3Y0qbzP3ANWgI88XQgqwFCs5pyfiahRYquQGNykkZuSsajo
cgNXLhxtEHYDnxS5DoANH43D39a1jnbW97XOgiXO9gpfDY60DQ0A4PYd/y7hPPlc
hGHASix7fPcDPSsf1hVxpAoS6Fg5om37idyCF2mtutM+IwMVdMS3aGq5XdaTWC49
x0E4m0SDNLBedE5qL25HZNBcZvX0UhN/8TwT8mV3Oza6tqv/7AjleCAmBOQ83W9p
YgR7NXMzj8LqbKTrqH+eruwit/w/KNJHI+gJBVQSXAW5KmdCun6UkGUKEFPJG65r
nceLJjB//hyeXErwwoR8yzih+NEGpxxp6+VdGPuA8Ls6fd7+QKNsWC48yczjCTo0
2C5ac5IcApn8W5Esmm8veFN4+MgyB5lH0Wimz57TzkdpAf7Vls6RS2xhZCaYNRG7
CLxB320m75PEOSxSV+Y0qq5tTb1CI2LQhUPXfq4aAKGOKjg3iDbDoQzCDzFhUWIE
lvxEvc4d4kjitKhA926X/hI1dLAkcFiHM7FiVIJymw8zfbFc1sXbf8naXCjnCltw
lhVKnhT9Ekg7W63zT4J65WWKFWr28c4lgzWTM7br2Y7Mc1x04+CVexv7jRwYzBuK
XVlK2HJh72yCbCmXD3M6zSnL4Y7zQNTZpoO/ruv8am71dd3B9tWKZxhZru+ZvVuj
cbbBWVwr2TviUWBLT8sXITJExsTxIXkpateTb8Ti1kUwwU46R5wWnNee8YJxzrTD
Eo4e+d/LZQFGj41xv60crH/KSW1spGWp2W8NBaffEPg1qFLjFLF6wKC0g9zE4XZM
0h5oDx5jEiGuW8N9107v5aszsAgqKNHNlF/urcyFPVI0RsBJrXRey3jmnOC7VeNh
0A6dKDm9Y0MlV1dRKOuhl3FQARGz+E1D1PBmECAFQNhNafEYGsVnacxhrMmelgCf
5ghBXMOP8cRVPaUQdmmTWLycX+NGrAOqJL3u3wnnf4ZHUOmoNadX1cR49XuAM37P
ZwDMhtnlQlQv+rXGgFjaElFGgwCHWDkkVI8jM0mF7PQBJjJP8kZBF1mxyDeJFk0p
1AMxBBy1prVvyKRrPbjJKgA1L4jwYv/wfvn1DcFBhsdsItUdHOkdmOOC7JYXyuoY
8UxUGklu0ZyHiIJpGlqxh27Emf23wxx3X3oIpuaBY0bHr88CA5jpx1vzy3ieygkh
l6LWNdGpOFVEdrpAXXgjGQjXOeLX0OdSAmqiFAVdYacyeRh2xY3GrQO+99AJFY0g
Ucr0e8hPeSQwVCxLTyloTnv/6q6+o6V/BBSaFf0ez15pzuxj+KeoV1lRbbniFDP+
L7Pgu7KN+fj/NhKEAH0xvUlIs7E/B58CtXhZEmFXTDoHrtyswEb+9luCURVHGdrG
Sim3QRdFGgIgq+pFFZEj45s09GdDT8V3PBl8ccb9H51cDC68AZxG2ZF2y6fYVmRP
GSvBCIZyHMcsp8lPZ+kwVzYt3nMiOiLKouTbzxKMrVbu3wrv5t01liRoeontpvDn
veG/raZwcCswjQ2EgeeEMeBTiLPq/9Rh28cCdTsfTlqvyH+LU9m6M9Uizf66U6pZ
5TUtyQCfTYuaajs4oq/ngSini6V89gAcevcF6l/EpqE7HCN38wRzXig+hYvx+ha+
8Qb7cL35r+VNSE+dv6jP1p1roVtZtPzDg0cUGuvcNrt9yd9W+OCgcTaayR3yVyHx
RQY1+VQ8IpZr58+JkFsyw51SPow3xd0sLauZ2E6X67m78b2I3oVwlrOq+n8snqkG
qsTlAzj3sNaRwe+ByzOjCAvnW9Gt1w145Q25KBXffEduTtEEjSxxUmQ/MNqsbHJn
SNSdwsFCYVu/tnNblt655x0jZRjlOoM2CiDB6YVIvtLL9saW6XAaC8hg4gEp/r4s
EGLJ/L85yeCGhrX3vqsB06QPxobOOWNseNQGgdw9EuE5sSqxlu/IRJ5eVUPGYc/8
jdi0BdSAZ3GHvPWjTpY4KIjO5tG9RbGFDwLoAUsR/yuINbHWHyKIXCEdoLAqE04/
M/1p+IeFTURpr9Smiw89EHM9r6yGPO+ovoYrkpuboqSbgrlQWVIJTzo/UwNxtzI0
HBvySjFynWMvqXzv6cPbT0FB8vm+Yzt/J7oGNLp/jZf+Pzwqp47wOEo4dE5Mvwvg
VkpUopIAb4VEjEtG321qgejC2WyPhgVS6qrkpyQ627NnCe3kcn02wbNvZ+9QARTO
oynbb2gK15qcVmmNMpkFU5Bei2PMqDENs7RiZolNEtVAVUEhKQx3EMIfAG+VDbe+
NL03D4qM9a2lniDlBz3rTeFP12JCf8Jbm30OV+0a1TKsM4Wx4aL/QDIWgaEdhs0f
w7f9iB8BqZzWeJbY2LcLKtG1pDD9KUa8Gy6XMi2nomXFHkD90rdFXacFhID4NHRh
nhEhWAbMqqeyFIvT22FVgR9taaiHXkCfhD0MI6nbx1IOxEFu9Ji16e1kY8p/Tnmq
pjAXPIjz3DzwGlYqrqLXhPsGkjkF+YPj73pkdwVPH+XhiepxviMBD4v7qRAfognM
XM5vqRupU3DTI9TFt14mZG+ys2GNMnF/VgBlIh+vp/Lv7hpEreI550jzAPE2hLrS
nqVUVFVcKXTqRo8TnX6V+wP2Jpx/N95D0pprNy0slmEkYHEwdgPVwMpGOMvT3rWG
zV7HEbZnbNghjbOF/HJnyiKx5F6u/h2us1cxiE0XmDMsWKjTeLInAtK5bPMzEltB
EOL3XIi6IgUDAn6vFEi7aAn3bQLkPs9Pws1XRIrHW4+h5oKlum1L+O+yOs6f+90c
Ro6di408xDKphBrouZ/FHxUAwRvfKRs4HRWOE43Qmsy7sjFf9BQ3v4uaS0uSqvrb
qXotG8FD9KXFyp1qoff0oc6h/anIM7A3orWw1laiDC5xWzpEq+YTjXXB+aRFI0hv
bgL+BLFihbZTfWvpk7jAgN3K/Km6CcRYZFom0de/v+9ISIxVcgsHaSDe4Uxtow8V
0RAQOzk+fndbMwWpplCjCNBYqKDGa8bkqWzL6pYiDqeqqP8gpbm7X0zI7tRUOqZ6
IKhU353DFtBl3AsQoxDs4FkdHZLCKmvaoZRteN7bPqntsSI0zzo4B/gPvSJr06aY
lmKn9fgag5MIQhrqT7s1oNJ8T8qPxdn9WH3NR+d6fMZA/G3n0MlkD/vYms6r1Ww4
SjoWNdIglKkWC2isiFFxDXZsRIzKuuS8Syhzraz8ieEUacrAhwPUvhPjCtmDfJsC
GiNNN+9iGOmyxMR1IgqIXFu1jnOkzvg+jZvgjZuBWgOTLzYRNjIdOWyeKS8NU8gu
IISOCC7YulImF6SLUWiaUrFQXe8uznpx9PE2SBiK/psCsu9R6OcK0OFVUiiTXzTS
OJ4UgnhSIcdY8odh4N8Ty/GfbAQt1qafrop6aN470LDuYfJuxrnZ4sdGig54vXYJ
UBsLSRRDlblOdDNCJ09BNm+lvo77DfpjF3dDgr+UC5lEB25z0Fxb4dhP5ExB1XZi
M1rhY0GXaRL9mbHe2TqRFkXsndNWIxtbsBzwfD6oj34bMLOgIq5m5sE/DY/q8Sl3
JN/my63GyHo6nDvEbZrfnhrQv7ctcEFE0fbM6uxGoByv/AErWhifJvTYRUy9AFRw
MPfy55mW4YkcAZpC+EZiqMLw2lXCALRY1Xqmjt1BLf183Y2bCJiQ1K0U4kNpCHWG
vV4v6D7cr1zyILJWm7RzscVbQemZb0qjezDkRrhIYoc/4foGTYSQ+LD/OckaX+OJ
tv07OHbFmfPFhmd4RtRuKa5CLr+bjpHXjt5C6cWTSUshJQz3XBSCElUsq/nH2cpY
UZTMIEzq1RRkitjxj9CFYRwdF2a3P5IHgwjcXeUsJn0EThLHa8pB38BWqEJZ6LLI
PBRN10UfG9yNGvt91cFeone1ncyAR/oZog28cb5nHeB5njmdKLJm2hH+4ugV1XDM
wn3KkWiSx7DNtC3pA3s3XUogvo77tbhYsTQ2UBsPGisgG5POA+4ZODLNj+y9+Afs
xl+9bluiJ5Eo3SU6EOe8p7fkpk3oJGLxRVhdxFfTe37N/ULQPD/L2hWG3e3iqtIY
/r8acTbL+4aZvrPNpDZdsPxa9x12B/+hxtSNEo87P6Gnb/Jk44MhfTPeivVK0+b6
7dTDlVO5eAHNEyRqztyqCn+8MVWfbAhsYg2oNHxrlqyagxVbhEaXvLa0sBTDI9AG
JwmT3v3KyXazu/tNWuByrwaBZduuZRdcnhYeRUQqONkExwXKO//4EWI+hNTn6BL5
BepeKqjT8c/sAaVH2YgEQk/fwOVlIxSp7SPSo7MuNpP89bVGnD6lgbPRK94/jZMl
x6Dyc2V6vv1LKi5CHUJiHP8jxdsi7PFkp82/lRklVlk6XyN0tpXfpTQSV6p142NK
LAUJEQiF82DaE++jewHXft6Blly83HbLB99VsthOk8k1Fkb7PCmALvIFhl/Ir9fF
MqUmln+MghD7V8G3T4Q4LEjsjYR/0POlxDQYUawUZa/Sl0wuClV5zvdhI1B+xVUX
227XsaqbVumWKlTVAqvaK9kCruAjl5aqjPFPFsAXgy4TewWYox+BOyDlbvG6cHsX
v8q/QjLrZvngGzvzOxNQE6DnYZAeU4bYDeFpAbJYrYjPmxs53uCSWH/iHSxz/q7l
9dyClFwF9M6xeDAyA5puzOB/RvaegR5l7r5IjpOC+vgmjQvHZTxJIpmP5kfIDC3i
+v/Gy4pJBGVMBcRNKkoxeBONR4cK7T8h7GqSRmCfh9qANwGRjHL9C2zmHlLHp+ZT
MGCeqw0bvHviNuAlUUWEUIhpcQPl9j0enTYBzc2zLla5hsK0mkGiqrNWNdBkHaTe
mvC2geqe2U+XsocMi3fbPSqYmTFVcQiBVqdJwLwYLnUODk9pdBBH27MXOk4btpxT
SBKlAU55UCfCH0FdYPX08aJC0P1LnPj0GkdATJ5GDBdOfjlVbaU5zdM0pUQutErl
/6ZEfFHVdPKAcEbsreWNnRzADUp7nnuK2KYe54yUXCg3wLzyLvSJK6V5+F4hBImF
6MfwHskiGKOTP6+49QkFNZiQrxI6XBMxluDnE58ccziFKxPZR+v4qIs1sDuXRW8r
Lkg+bgVEybOby43EMY6MHmAzO+lLlHhe03B7DHknvRcZBJ+oAqS0HYASSQQswWNc
WffwOP7gY2O+EddAhzurKfsUHSm8++EeFkO/OnWqWEj4SBE0z6beL00AYMSb7Er3
oK+nh0z2T1KsUbnpkqZdir9tG3hwDpZQAfqgHj2fTDu8d607Kbn9a9OQDKLwkVJ7
OPOlRAl1GEo4TViULz3YShMtqvT8ERlBcAQoeoHY5XWkeVXrlz7yic7v0YrwRR6K
oQLgbn5iSwngq2WIkJdflikJ+ZA0YZ0etN4N51oBhl4Bm+KCJoUfOI7Pcajf2ZSQ
BjTmViSbtCFz226LCjQekbtso613kjme8G6s581sdgaSU101OTjtJGnpfke/nRul
BsGuDNlLFxMwSALhYF8A23hck3uvo4i3VLlM5z3BpT/znuWE+4odjJHtfU9kwNcW
DbwSePYzWyx0B3MumtsjWBOFC9gACR2gWlkrz3dbAdSBAEJWZ1dn+VSRPodk8WsJ
2s1qx1RB3dt77qYxCMU1E9PnotVdn/XcSZ3PfZfZyt9xbXKnCL2vNT//rIxvqzPi
BXmhGMod5jV8bh1+DJvfhu/7tGtmPU5xrOxTkqsEIO+tectCCcOsENjfpdvgkTQv
rV9iFZjcgJ2pqVM0jMs9n6uLy732Cbk8kSdosxx2urml0bt4UepoMIWzC+Ad9YNN
fq8LMgulLVUlwPBvPYg/XFMvb/SSwN9dvqngFoxMjyNYMzVRO0yevTbGlKe0gpcL
C7zyPwW5hp8TE6k1x0ogt9+I31Gk5d57HEO9kju84A8OGlAPBrS/ZG+fXrPxbz5e
sXY1aVRBkjlHdvLsE/hJ/Ga1MvzzAkwDJ8tgHhJJo60w57Or9eOnmhuNqSRGS9B8
h8+vwQ45+Q08w16c9FiCuz4E+0qtCiUqMlD0rAuZ+sC3ufndd59EoneyDgv5DKeo
woK+JfZ/WfWuuli7B9vl1igPRuDQft33Du/MP+9XD2g3xy3rHnym8y/1XnGB2Dn2
LRs3YZz3y4NJWLHLlHA+MM5ZM3eYdIbWKQrkQCWbEh9DdFkkBcROhVaLVsdBqBs5
R/dN810qQVXXs+LgGCRSxzGTaCORIAdHEmlaeTCi30n/LqQ6mqQR4XQKtirbP1lv
Af51jOpbhYmEH6/K5p7NlZ+kaurcZLWht4RCMbHcAwsruoSRzGlOENzBTfFCBUj9
Fq52PA8+KfaL+3f9LSvzucXFyqPBlNxGEUDA1B7l7+O5PqwKWzXMWEkKKS7xmicE
K/j7CHMgydVczQTi8DAHl/Jp4pTE2d1c+1aQap2NfOiUFvQ1wzlPnK5hPinkkvq3
TO8+V/ovFt3dpMKOe4xEc5b6u/z1VEfiJW1b1kVr/eAFTDarAXQAgFSWOr9DiByZ
oPgT59hp6+f/CTmF4NrOeXnaSYLQxISziMt86Zcdsje+eaz2lXVDVuCMXbBfNpB+
MEb46PHCq8L38mbN6pYBTcfAx6zKIShm2EHErX2szvn1xSZDcsJ4k07VTL10iXu+
Ut0txL6qoXM7IWv3bbMd0/Ek8gOZa0y2nxxqo/Rq1iq2EWszFkgLOFocuH3wtPVC
yyVgXDqSlbvXmw0plzdq50/E2Ady7sbf/BL7sD0VyWJ3+MzDYZuTdvIWQasn1js8
PY4R2FH/3ihJi8iKqHGwGF13HrUJYFHwiKk7+GvSLeNyWQQXt2B0JSIARDevL4/w
TgMomvZxB8EyWrYUzDGThIqrsx+og5MNQvD3QoVWDG20iAzkZtQ9cReXAMhOUaGz
Xsw7RcDGgamGLEjBGlgFs27UeGRDj5EziOVstGiRokOiXRphoIwki0+DWOFSGq6/
3qM+XOFDHkO442bhB6iCXM49WhQ+zJEOeIHJdlof9PQFciZUACaJQ6wliS7oFsix
pI5ahemT8yh340zbK/v5KHGx4wB2fQTc54hdSvtflRat4ILcf9CqF8oXa00cLx6D
MatbeYN+/WuiZnTn1gAYRpJouVCK6FQUNrSIRfGhzXdW/v027oKTTi/sWw46Jb9s
/xhgH54egymj/lb36v+G5q0KZGmmAMdufyDsFRZZaQ15cJ+OM+3d0d4wKD6gsrKD
SbT79+Qeb9WKB0POGvbLyAHIXWASkNI7y4TayGD5BvQeAnOhVoMRyuTVP6QFz/9I
w53JEGQzUBH0Sbd+4EZApg4vnU2skdgNbIAMrnXszzrdLsnv4xtnymufRQdDtFcT
h0rJpn2ZIpojk1AX5QINAYdlm/olo9vzq55ZF9jtgiNz+s5FaDpOrL9cTq0Skq+6
tSiyPTmunTYPxghDwhh/X2K6oOOEY+uQKu4TSAWnfLWVzvvHCIott8CqNMfmeM/8
nSLY7XiulkUNnOsQlEmw8RH+yJQVcFEPIRZdYt9c5EWLvPCJVQIY+MXfoNnUwyJ8
IecZuGlZQ6x/LXXOZcruizJ9EqGo/uYQwB1+ti5RFPvgpRyVcJrtCVS2E8FvhE+d
ghP56GWSt9F11xO8pZY5Yr/oPQQMCnvhQEtdgfy+uScuucHO0tXFKkRXI9bXmUWJ
t6YoDK6lnOIpAuEUYKUblHEI55WdvHbEMNDVZaGSG5Mrz0xB/TmL/ym/z6devyC5
NxBa4MmqhBJnutn+onY/OiIp7L1n4FG7Rr1qnzR0PXJiLcZq/seNYA3ha3I/E45u
xzg7SSDhQB0KQaVVx9cu7CiPPm4A/t8l4fh9O6PkrsR4Q9oqc+tL47dBtEeo0sJo
Dz/JG5/BR815WBoEvp36DhrZaUh9bPMWB+IbZL2DpZQ0HnK9qsFq1r/XipjHdiU8
Y9rx4JjkOzUb6cSNVkfA+fFrtPs5MPXh2IetZ1oY2ZZCzxWBvwbOmL1pTWvWF2B2
yCi0OTLxLzEud1UHdaJijLbuuVdlWyvQ7rZd5UKvxQ0o++f5XmcKMzVrY6yevtSt
n5Y3g53C5c5gS+JZI49HfkZdWurx4bX5J69EriJo59X6CIMv0NveLuHpaO0VzHWm
n5eRuJ8Q6UTWTvrGHM5zRDpgcH3ApnPDrUNuq11FO/1Acd1cGhkVaIxG2BiOyKze
P4o9Lw2slKAwqC6QctvObB+XeNgCjgzTVYYZYvnUmoGXOqK8cJpdLJmhC6FtXcVo
81dtSEDnrc22qlhosjHW53wH7xP1VyZL9Uo3UJOB6deFfpTYHMZxvjP3oFEyEngs
+cQAk69liNdrPkWF7h0KcPCYHDXf6a9fl40YOT22GIEKL7bjb2NTYTyXo36mAsDx
9oDlndhIW/Wljx6LxOsSDCs+HLL12z/qhAIHVT1q6W/jnyTJwPQza0bWY+KC4Ruj
AeYZzXWMRjPIvdIXYd5HENo8j5CtE7/h6V5Mn1zVtHmEgRvcu6o+gD0UN82p2bJJ
ixMpURBxKvAZ1A+Vw5H3rBpk1jPWSNCS+boZFf5KYtZWPRGQsuFl8PcjFC4Soitf
4EthIn+KUVr3VmoUztuSxBimokS4F6D14djx0I75NjI367+sLnB+AZTnpidq32vT
KUFTqa7+TNLNno2o2P61DHAWjaPUMEMXq9/GnHT0lxbLIi2qlyfuPnutF2/QQe1e
U6yPHc4RPs+q1m/oebZkSxyifM6PPLzEb5/A4huAGY5lIcgq0R9hf/pAqBBHR5p0
th0NL76f76jI6PWh8SCK/pCwApW/DJYsRhS5PwbESOvN+XV5Wj+4YCO0uFAry7o6
QxFg8wXxo++le1x6jvpI6y6WlWDrste1+spxAvDNOl1QN4hNkH0JJj+ovkq0At40
uNPCTvtGzQIuI21A3GWoWf9kAmEAx1ksJtyULIUpQnMAY0EbSU2OybYFoW5G8NzJ
2wwfDt2zuYR2zZPTtn/5G3IOuD8mLrIdHgQyImFZn4PWSkItosEBakQJzXM97nCb
mK8c+/qXC5whM2bbnYLXyq7So5zKfsGe4SFRh6U0fmnc83ozmk+eHKL8msITc9WF
4zW/e+JK17SG3IHGqoN9e7euJXnetu4KUaotk7R9now9c1hdFY2+6ULAyd7/Kdez
vd/dEQ2syKurywwpwkk/udS1XuzUD+QocBiGkqfgsoAD26v1h0oVZjJ4KS7Z5xIL
P9rSASCM5NEoF3ZTe7PMF0EWo0At15poQj/UB9Y80MuuzI3bCJed2tULfCMa5bKm
wKBifMDwocCgTpet1Dgx4L4/4tvwPrYwsUb2rLfrM2i/S3mxcv+3sa+P3MPJMn2q
/VN7ArKNS8IcgUDoOlmo4Bd1GycT8opf/Itiq7HcALjvB+r8XbTOPSVviWAOqfpt
N9jeKYWxlI5bjxE4ao9qgK66N99BPgde3NIqitSV367m8Oam/oUvjTtx8e4XUgfO
ZzFBGDHbhhUPpJXz47kSuWAR/N9SpvaL4LkI+/MtJUHfrGNVwdySRFmZQuG7lVuC
8dO86gC+vD8JC87DFi0hynW0p8eyrMTDlkh4FMqTKJzNdDwFw+VCT0Y0OA8EjM9D
ZKlYtJUbw3B1PUVofxQ4xwjnGbRRN4W3WFjX7X5JnRoFfW6X5/dUJqoxBPoCVJl9
PZh/IUmvDCEh//eU1jqt9sT6jKDJVNLHlQKyUwRuA3Y9ov9yI+dCv+AFgctIEGAX
Qcq2kVMf+dkHxn/uJSGtacpWHtFe3CcfIfk9/JPNpQai6dCx7CyqLWyOAa/1hymO
CIjygVSG+OykUdSZB05DXPoe1SRwJvFIrNRRIQKBuA1ATjb6FIX0CQGetzASsr0C
SYuGLzux0VZTGsC2hSnx9Ei27Wlbg2hsxNddbjk2fsQZ7+00LL3bouKl8Rh43jUw
D/eb8LNk+uliEmMamQaMQjAy1cA/csV5vDkEpKcKkeS4oOj+jHIWv2D55WidQGt7
iUsynoAJWcecFueWHI/396O4QBt9+mIuns0kZExy+jR8JZBZLaNkAuQoHAIi2Bja
sGcTjLwEtk0QFhD9ZSYQuiyRpdjHKIu8wMcXW86FKg4aJe6E+6u0f6LwD+23vsv9
cDemEBQ/WUIdmdx6XLX2cYWuA5eDR7PJQB0UFaTsUspYVlypi4C6CD6TyyWMKZ+C
KmIFB891PSsTGHa7eVIu4HlbGxdbHi76e6u6h2/rxG/3P36XR/2ltXy8BUQBu3Dt
yt18JxrrSfdiA0V6RTwovPfIleTr/0IbI/0sEGaXOUwkXS1L9RwFKSI1+PtYWFeB
ntsKgrGKv3BfrtE8P/X5J81FoKJ6EjO2GaEwS3Da0FPx8i927lJoIoAR20EJUn9R
x56lC6H5GB4gKTCD5x+YapcEFoOVvqi8b1LY9PsTFDPQ5MN1irLK6rGrGxFYFnVj
4rI74baesaggZQ4OFQUd4/H/PPo8Ws2Ze8wJrV+Fv0vqzcGfKtmv5SjrmxBoWMQZ
KhBkmXlZXJzmcgaPdy2ZX1rTZHZ+mkdL8RQOSbrM05yvkZqOAD4bX0y4Xmo9G5TK
Wmd5bUsXD/JzEvMmc60IjpPTCdSTFcEaJyafxCUhQ/WFA3YLyvY8X1dtX6rfUIY4
TsYDSdGV/mFgims+u+zPVwwSaQceOBCE81UK6ALOEPkTYpzMS7jSE78Bg6YMutLM
vwuB93INPvl8Vh8J8hhNYFmZ+m2SPiADWrWBnWu+hpfsqHW/Wb02UixzYienFS15
0MLYLqJJy27Xc3rsxP79qsfT3+I7gy7nR6yHq8nbanrA+he+BTA90CJJZkp7Hthg
a7iZt3hBIWqfr1AtSnJ7iP1aPPEz/zng2nZUyA8dMtx5WIdw6QJOMSEkYhDaE5pK
s107APYNcJ+S9Ez9yAV1CFndtfaqiuVgdt/WSnbsp1/1vbQiEGM2km2C7lcWdJVi
MSM+GGdd0m3ZB/9FyjBfImZ1iOaz7f0lcLuLPRz66eRaj9S3xTA4dCr8ZaXA00A4
Yi85l+tVYzEhwan78stCfeWKicpGqRfLrXplxLKffhV8dQzOE9pOHbtp1lY+dvMq
TTsAeRsaMP3sKrcLgfmHDi14B7Rfv6TIYVcjqtqSQ67g4IpXw91OM7i30FBs0Bpv
0tVpzray3b25+6I0AsvqCiVo/emW1gKKsOf6BcteND6yjIRNwbHKM4e7pybR1nuD
/XzESGPmjkijgexOTATmLsG9JWrP6ZAAE01AxkRly+1LmsuaPVfCbGaOH5KSgWTy
uQdHVsRdDrrq+dy4jz0K9xlNKGyjSywDMXOKMiu1jKqIOnfDxBR8CRV7nbY4sRmc
IXE3RCcDSP/6SZIfJgRBa/W2Zokvv47UT3q7MFvFNFCzyPSbkTG/RwcnonxaJAIv
Y4t0aswpFR0+w7pWKHFyJ6SZTn8lsMCjs3eovmE+FxdCG8AEKHtmD9hfaYPs9JdP
W75Ut72HDPoWY2wHkTLJowVi9/dEL7Lo2X0hoH8wl0jvt+rs8aIjM2p5MThnHUX9
jR5JTszWAQ83Wf1VT19QkKNjAvDtt0P/bFXs7wNeFi2AqcGefn1DCDyFDhhLWAne
4V7O6r9F6CMQ1+LVWExWWMN1blV+B4okA02VWIzXkYzJGvXC1a8hYI1FKO4m/dhh
gRjrCgMNUChB2MSO2TU+CKPM5hTmNvADRnrzvWgeSwm8J3vOeSd8JZI5rkW3PXEQ
LUYW19PDT2zCbvNt6VmjBS0oKTV9RKrmyUcv3M2KD7PH+piHcuqt+yWX1r6tVbVe
44kTUruOxk28x+ga3InKp9RBK0j03nzRzhStdgtdbz80rPlrLIS4/PpOuauREaav
4fGbiSQwYoMrZwybyczcdbv+tmj39owdcKGlqWDEOSuKGY7apxrOQ1TOC8z4pu/R
3+uQ+yASOJcmVuEvXiWGT1jW8262H5bNAUS3ADs4DWDz0hLhYWafEbUnYpqq2U4P
H9tm79NJsk00T4sb0X0OoVxBytUC21WTdSxoS0F/BRXbl8DyIEWy592U2C2NbMeJ
j16g05OGLxrv3pllYYAIH30CxGePG4P2Qyl1qAmkdUqhclh1WPtHAebyG6d/VbcL
WKPQCaZm1VM9JQhdYd2Anbam9+Lnxgl5wA4z2+t16HWmLbAnVO0IxsmJEPDRphuT
24+gmRQtqhnGxY3Lr0Mz0eFGLjJGXenc/ygfcOVjp1OfMMjsNFW2CkHqg68SKfcE
aV5dKkA1GfDjrdbeVNwywjnaZyaC2xDNUSJIrVTBWK/FHTQ4uwqZQZYP7DDSzbrk
Subf5q7KpLWE8zmeFZTqXr2E5H1jzkyK3vrtEfi02AZRN0jtxUJaV2ARjWm9HDlQ
UsA4NHpBrYy2zjHK1K7FnL6fpN0tEX1pd7vkdl+Tw84crL5Ri37aXxrJDTiNjGIg
vpJ8Mh9sE76SMxDLYncf1MdbfDj5Ka6oXLP220BbNC87FvJhTQU96qmInr648oeS
Hk0Sg/ur3OiPA37ZTB501kaI/rMlkIrTKT6kx/tAuKlR3zY7BH1JwbA2cEeG4OxL
877YLLNmWN1KmLZZScccuUJW74hJyZT7cSjX8u08u5vKdGrV9vM1PYqxHmW8cxOQ
Eh5rv40JjUzw/zn2d+aPHNpDyurTeWV8sHSYZlHvtzlkA4uuANdioeBNK5NwfCfj
mv97aOF2VDEB/CMonJLKR4M3/pzilfjmcHdfxJWJu6zFFvmQITZinjlCs+eK7VWn
QTKL+wtyS4RaHSEQC0z6QR+9BzFUxrTe1Fg6nWruhQmgQC348cP3u3PumCqW3SCx
BTi4wC2FXWk76WitCEaDpESCdm68r0PnvgNM4Sgl9EnP5krRI1wb2ehYnUdD/M+c
nu4cqOQJuGjrw7L6idop3BiCBA02NNr75c2xpNp+7Cft4bNWwJZYNEdHrziWmGxs
qhEPd5Faj0ZkdvrUug8PaiKi7g9LXWjGRRn1XxkkkU5WgIYwqsxunwI9YYjuthZx
UeYnnxHFDlkedLQ9Y7KxeLi2sGruBHhQEf5sOedepilrCFGLwHfbRsd8bnZkAi+E
XlKANAg2Ci7r7YpinkF8721r+tCvcV1cymkohmI6KRYb6kIIxdu1qNpYOe+WN/oR
pU3pLSh29L3AEt2r6EmrupcCum8OUNHJR5D3EuJ/qrWI4KjSj/WXGqf5XWmI+yjl
lN5IF5tV/7DuICS9tiMqyF2BS871BvOf6avOu5nzAhg77OlOhs7wNRGDb28ZTVmG
oZJCAI1zNoVJ2+Ysw9B6+bpjhMO2JTmIf4EseqtL7Mkp+8MLqqbncw1UfcGqElVr
HQcR6x79674TtnqdBpwEXjJNgdYQpBjqXEhEQeVsjNbwO6O3yA00rlUIfr6M+25/
YcURnUzE1yXXqMV2TUrt0dMd5stTwV9XF2SgrNUKMRwRRV1IR3fGm9x2PqD7MWfo
YraoHaa+UbxG5dyiAOMJSsyED7sqXkV6GB6OA+bQthjJLSK8A6i556QwYx6Fgxx5
MsjSWgBbO6HHCaqlmQHWpTBJJ3OQ+1hcH+fuQ7x2QnF0QG4ymUytHvO0ErP1ANcq
n1kczjqMxfyC1FogE2mZrlZalzf9x3SPN2WBUTyzomoJ+VfGUWVPMy1b+aeLwrSu
VvFQMaawMTYQJiAH3PmzvKOs5iIHOaxpL4zO8Aba1KeuSy+Z3do5iXF+YLKOIxvs
EvA0OUdG/FDyNRpQ5nmscgf6v0ZpIDlFr48O7y2T9wKpjKJ9oBx4cZQRmglvoAGv
uKDGXStIm38YnebDvG3WOALZD2wwSj0VYejO9ebWTeUU2lAi6y8hHIjHHI783wz+
7LMpIYpLvWAc6LR7VZ96nr0v7j25yRA5e4+gGXMnLMSwNEWUWW4qHD5609EMLwRk
wQynS/dXBl9DxoCJt49Jm+IpFrLiRi/79YIJf8mGGK/tHmszYo+4IpmT/oZnPUva
cyzYBA89NYWe9kxO/2pY/Vtw5yZSdPrZctTVhQ5MoDqU3aM5SNgWM+FtdcnKonkx
vODaVoSzWNqPhiHMxYcmowMmfNxHcKf5R6+6jfpXNwSKuRXZ0gOvs/VeD+jU5KEU
I6aT5pue7adCx0o3Rzs/KnObW/FUI19BY2uKvMxHuwzyxCKDqLZWg7goSarKM81c
CZPsjGAzzlpgB33UlkDUD3f7praKqxJKjMlQq8vEHCUSmDrcTvXsrcFiTit4Mb0/
ZuHKoSN5ZcTYBcUmNb+/qfQDUGOwOimdr/UgBDkXboxfTK20Z5KFz4LtQtrGc6ga
ROYu7bD8fBG7FKF0Tkv4YZLyZQBHm2fHk8WZryAinzITPENiAdyuGH8vhD3wsNAv
wcszyJUme8meQBT8L+k5SsxVhooaL5F82J5sCJDdSVtlqpOd2Iz4/QFestthkq+1
LbOD3bUMQZoh971SkLIlqgR/N0m78mbyiKjyTFfya0CePsgHn765T96NULNb2s56
hAbCPFliAFsbkGez9pXmKR+/51gplo9T1z5TKT0po1Wo8j68aMCQVTW9eX4gjfGX
ESK0UQw+4/9pKb713PZciAIkq/MhByN0P2tuCNUbJFg9zkicU5hpzzw/8wfd+Kz1
RncWkk9AJ0pEqNFTqul7Zjo9wYomr94/l/XehMUniyeCj3JEJE3DANydzawu1YzU
DuB/CY2Gi0w9SypoPrxxa866rf+uDfGq8kAJG1Gm2LbJG3gs3ZsSEv8rRDLEqfXV
p6CRl1Y9XFe+PookKaZk8Ij6Rpa9s0cTBT3ega7OAfxFMqPKJCFEavqOQGGGMkKp
tt87op40KubHgPnhJt44eD81T+1VemjHX+iA5qmECd7t1+UcaxAbqIh/nHwSUXdo
JGxPxUjE+z7ote0Dtyex6Jj4f8TWfiCmaz9fT8HhkvrZC401d3A7kr7Ou9e5DMIU
eWpaiyHd2u53/9epnsZ2bMs2UbbpGAId+hjWQZi2lUSU3ekiiFD+r3fDGQYORKbr
F7ETv3jAsxOYM162BBVW1zW3i72K/1+x/KR9DlQjdKRUOODsDIcNb/RcECIvJ45W
CizYdC3jvNmkI5x3l8RtnlEq3zD0KFT3l9v+++O0IVscm48jebvWjSIkaAcTiFhl
3w5N4NlJSR92qaoDvU8uS/HXoSzwFXDAFUFyRNlBUBRyH8TS05/ZwP9eD8JUbzAV
VfkJmSkiEtZGuLmysz3f0GR9Fa6pGm/XU9dFfNZa03ooCu0ITkj7m2Z8+jjnC69M
xzhpDmOCa0ehy7sF5R49Ryw3jcJvmegZM5kTaoDblhiJUlaO0btZTraWXty6hlTB
TkFGUWd6HbhdWxrKHtjJal1vSZXD/pj3Yk1TDCxHU6Of0p44FGI0BQ7j+rWvOslQ
8eHpoxerThWrOwbb/4WxhSGI+u6PRQgOmH7Wy/j2Kd1jzVXICMjpQc8BIlftOeEU
d7ZsmS0Ccn6broCnjLyaZI3hs7Tt47RtkGwS1uOCdYtS/FqYRW3oAziTlOGv00z4
CYHE8xmuIlnpJ7bcxqAd02n9fNrGHJ/L6hkjyDm9KSQ7eTcp3KoyFCs/LoUfkXzO
ZXoqzmLXyEEZSwVTnK7namoexu9hZADUPGopA/DHxvpYaGPWgoSlfc063xJWpC2K
7uf7Vwo3b/CkA9X5Jf1We+SG1HBN+4cNLUyHtajZsX3wiBI/FXUH7rEUJN0rkfLU
Ef/ldAnYgHAc2EAuPI7JceNvKdmwXWv8OSKQA5Y7zR+tbo4uEXOsV+9nxQK9e4Ha
0pf6UvI2JwI6dRpZftqT9yiC5WkWKshmcMEdBHMRIQv49Yg2KNhNhdNKvEZ01LEj
hXMIOg8K3IABqt5vkamSiUtkyp8gycWcWgTOVcEup6NlPzg5VkOgswqqLhxP7TSf
Dp6QNu7ll0MoIdY6NYUqoJAnD/5XPOuIqMzJ+YTUuzFZC1CZveP1zqyJjunx71Sm
ChHKVzgxijqsBjEn9fuyJsaQXyevqdLi28WuGCRcJ6FaiB6w2y2NhGbGfFNBp8M7
HNW7ZsQi9dZUsY+Bpbnx4gWOUFzd5SIim05b+mFXdYkzu3emGRjxejb0zEwJ+oUK
55QHqBdZmolGV2j18ruhIMrXAgneDxm0mIQZFB0JNZ4Qd4cJY+T4vPVQe/vSvdyR
7lofryilvUM5Pdudrl7wdQrbMaXsk1kenRfmVV8s4UvixRiBUUH9c2RqCQUZETi7
L4noCWWwZikcKszWFlVDsCmMPdEMyjXARZsosO5KOFhreDBZVdXd+IYdjS4ChG8n
ubbYun+q//wWo8l3M+KB9V4sAYIV6nIY8C9Q7CK6lBjbHrg4HlL9/rGY9Ued8nPU
4ZiFxvWC8Lg2yGbCCfXxbN01M6tEuPv1hbm9/a647nB3bg3k4vT6Q0VbalEs6UnQ
CvzoIBt1k+aLZnQ/yvkI6dfp4YbVQgxsxErGIafW6tVM1qRO5WMqKgFVZfdyyHvV
E2LOhiNWnS+K86FXEi3ylozOjR88VaPbdCKCBXYowlkVjGIhRigtObErdVXNXnJi
tKtH0/egx9veN7KBS5Cg1RR8huMFXLhiENZjzHY2ZE61eK60GNSs8mFYtsDZlcbS
lPdcjPfUkVTNeXos0AHv8ZYmoxIJXWKB02mvn729HXFmeOTahPrmF9/xJEi1yAw+
DRZI2RBvdEqnvxMqBYLWk13Lz5FQxCuOB/1ncB+FG+OkiCjU8d5babPJlE0McCLS
cS0hdDl5tK/X7tD5nn+GShPikmqJVVt/ia5rMjb69ZRC9Et+vaoX/09cVxJ5aFhz
Msj97GO0CQ86Xw6e2cZVnocTfdJ2T9mQC+oqVncmJDBQyhG/gnXApNg8fRRjgBF5
713cNqQSo0cEOI7eicbp0hNeYA8umbfVXFx2A87VmXaSktH/GiAhM07fVlYIbGm0
4vziljLQ35eugliAgjPbX3HzXDiSThJp1SC3AEVFgT7FwBfBZozDif9TpRO4HAhM
5yNt5aukafMJjLKiCcpTrra577KUJIuCdt02gsFmAhbrQy2Hp8vh8pucJPOapwfU
IYXhviSgCZkFAqtC7zKWIunqsBFu8J1Nzfddhx1SVI7JsXqDq+HDBiTmWCX/20R1
LtKyOxd42812pEgtPOOA9VOkj/uSB+JpJXMreSX27CZDGcgbWOkek6aApgEkmH0C
PZsKpfgfQ9ZGRpz5+iQfMBWe140Sf1+tmHbIj7Qn4c/3Xkv7dkp4oUWWL2w4AJVe
rF4noyXMsfhXvZwQzMOCLZ0Tcn4l1SqPqhN41ot9vdJqVfHwzEFZgLYPhutycmxV
Oghu35DLZy4Olo32PMrUMaGDF/b1EK72vRzoZ+cZv02vzMNVT+vvMAvrkECLpoeo
ToEAHPWvQe/zypq90Fj/swbooh2jF9MssgvnnqTrkeYqSeyZqMV6aPPROtuKxmNP
96+aKi5hLgIApcvHk4VDxFT9mAv2juKkwaGXNk0fTR0ofelhHi/ew/TmWJr0a+BG
t/4hE0QXfKKfgoJGIHVoM2Ggp/YAleyGIHmYspIalWzKOemWNFaQoi3txBIxsiTa
J4sCsPQUBRbAQ+ucwCgBmH1D57tH9XwOAnQoVgN9hZTS7voZs6FYmj+H0vbyiMqd
ZDHc93WnEUmTRpUqXRHAx56NoA9Xi4YeVS9ks14AHG1tA9ia/0sgiNZ3ss9CjPwr
3J0+Zjg5P/89iMVFRADg/mFqlLgjFpRRmMMAGNRZ+46NeDb674fxWJw+QBqEd346
EYnXeVx8U2+KjNidnh0iNNflRCYPcmujwbJQPf8pHZM48Td+G6LGboWY50kds7n1
v9/pEfp1sWHn+Dloyf8ZXYO9PS1oJpMlTuOSkEllM/dHQAd5Q8O3i6aGDDGk5hRg
U3yjJyXUMUXmUw5msdOG+B3BbYI/61b7cdccD5lPX/A5AibzCplAzust5LqK9NeX
LLQ0SrWICU6IBCumqoFGnj/5gUNYKZ1VS82ETi0Hqqoq1Pvipn17j14JLwUlroKv
bCETc1Jk9l/hqNzXn34t4ZKQkZy5491CQO5lBFWNRGFK+NbwIutKs2oo3dVsFQFO
4kNl2NLNpsDmFtvTfPSLY61RHWhh5h41sut/7gyaOsG95Qurk6lyXcITMCrPyPhc
es45LugPGYyFjljKJcEhD/92pPA7CL9OUMANWGs5r2HppVTSKVeFjQ+fbWnAb2AO
wz9uK3Peg0QfZ7Z1SJB5MjSP+pCEfr1+yMkdNYqHjsW/SUlv83/CeR4Q9PlOl5Zc
SJ5AVGi8Ji8P/YsGkMVqP7WNBw7EV3HsOWX9kez/hpRUZMe9f3YWC5MdXodycEhA
q96c9v4mrAIGuMyaJ+mdNy3uHw6PX6X3Mn9NeavqLX0d1PmG0YKYX9eyQNODT/Ib
/MgjRyBT+yVUtP4eyOagjSN3Fc8CmmOsh0vOJw5YTBIk594WD66bSvhO7Etc0uE3
Xt5zrOjrq4QXa9tc4HWRrSJxFau3HglorzlxIlIhLdTk100FkUS/1jyzlRCzV+Wk
eAN4l2iLdNWw3HdhN8rXKiLx0M0MKgT8hmWFxbV95Posfu4puzKWPgo6gwQuhHej
PLt8RFKvLxCIdB2/zWjRKjt7VO3EgVRDDWHGf1q1qbfFuVupdQJLsUh/jVYQA8x9
HZSaKDHYyh3OE9s20fezY3xYxYZGKhrAemIwVd812dKX21DtB8BF5eTAK5W3HJMv
EOXnZ541dm7BEwfxjWg8dSFprQlSE7iOXfa4MT25YJXV5DNDr9WcHJQtZQYFJb+Q
J752f5rpP97v/bsIqBZ88EqAbtmo7chK8f1p8TDlJMomKmGHHZEjl2xNA76xvNun
xVtyrkVjRIzRpYakmkM+LDo5DssZqEgxmYTWncmoD4+A7uWZlY6Xrr2Y4vjdNpF8
GmjaaVMqWGKBfv5a8rvmTDSI1yA2N3gy9vTdgaC2s/r2rkHjeQluYdKZ1SDXDmjg
vdQYV7b0GY+A98+a7rsyfGkRCfzjcr8n2ZpFrSaFKr7l4GEJKKEvCvfM1/yaUOXj
Lvw+4c3kdIA8LsW4bxm7bazHFEURwrvMs+lc1rJu8kTtycHjbSAPzflYfYQoEgOt
jvSLbnDw4UalkBph4NebYf2AMZXvJ8AdPkBXHXaHlMrUCE4Rp2jxGui6RwBzvNXN
+kJ0LYpsjCUA0LIDbffal6ZtJy7QWioI+Uj4DZKKBaIcEwSrzZ56Ps+xaIjYKP61
DKyobdR+wyuXSvzNENJk/k5j0jKY5CkdoN/wX28TldNagN9yVKfttYDYcDF1BIcD
d+PdJnyahuHTHb2KJhcfa4SaPryKd0A5mcKfjn5oGHfbS/aNjtyw6aKsvzbWsIEI
eCTQx6pEGVZNzHL3ZXdR0puG26Q2pj2HUeHEDoMy7P8tWoQe+xfeDEg/xg1DL1nS
vN8Zbpu8FpUZX0XAlQvpn+psg0fAg0mMGOAtjS4UFYNzvDY0ewcxtk8CO4FaEYop
9iPRKbZHQeZ2k90j2CYwLQctwLXdb95NHIc/c5DyyXXU4nx7kwlGApXMpwRh7z7V
yN/MZc3SkwUvJqKvGWx+l3DoWN1+Ss/x3/YLpHlJixqEGVVY5EsQO0eGIB4PfNC0
fG/bTn5QKrx/Jq3yh36fa1lKpy2TC4NMYW0tw3rk2qWf5jrnfIxVRs9u38jrnJIT
2bZXGEwrbC+Q1goJtHNxhf8Xere/XjOSk8IiRjFdLVmrGW8l5SfbliWUgcy70d1J
cnm6gy2H1b9BSkR96aqqTdBbFGZ7V5FnwLwoeIMMmhGY2qSz4m1LSWFKXutuOQGS
E3sN1S9NdA4d76HU1fOiDq5Tlen8NfLg/wTe2IWOoxsSuUZMVv6GXwwlZF1FnHnw
TeRIREUWLz/9NbZO0jMKjhVE/bP7+kLG8RlRV36gTB2IEFfJGXgaVXekguavrltz
Mwj0ML5HnLt+Bbsa7JI5YIQImT8jyxXg6s71CIUcc4znsF57qM1WzFrIplIDcnmN
p+SJh3FWAHj5cMUeakTwSVViMXPcX+7Tp0q6Xeq3AkCzAHl/LuoYa9DU/qPKZCie
Ul2i2yKB12BRymRcf5+p/KhNYEXu09WH/HsSHTu0o2K8QXzjJ78SURW5EkppWHr8
qpajDR+8WfDKbPDsXW/mFQ9eT358IRNMhd4Ow+S22kNCSyAkxH6Jy6XBhfCrGJcz
KS2S0bNh49uOvP5paSt83N4CMNY6hjjRClSsPv/CFK/SL5IUDWkfmmAE90S7yNqf
Ucm2r60WKRjGH0bLm0wSUy0g70qX/NGEUSy+i2gq+OZC5f8B/NcvntcKIVJHws8+
en3pfVo1OmXtKVY28h7Q9af1LQAPxg/I+EeeFwGa5aQ5/1btewgszTCXDJaUeibm
SvIm7o95cTVHWnCoegEk8k9SfCiu+RyOx7crOKmBD8Qp5F3jYDY19FqO3yUCzq/O
cYx1B7scnUyxfViqFJLlk32CcAanBztOScbBI35i71cNUR4N79UvPoreb4gY3kxo
MH/eibRHbt/qvCHfRPPbZNdxEYZCNIcQF4Y6hAjo3BWXtvFo+nwQ3MNii7y+spUl
qfVHGtKg5lhqz+LV9l7h3jnC8F8n+MBZGCHaBLaZ7crtiL+ZX/y6jaJN4D1xo74+
X1hHgGC7IlElcBMN8TgiPHR1SjyUzhK2Tr5wpOnqJb9VK+OvdXInJkcmUDK0A/ru
MGWD7vx0fnyk2syVsSEdfOPfhH8RLhyd1iLx1uElbHLVoc7jUlx8FSJT3jAujXaL
wzNAcotlOKVaEvkH0j4gsUiL/ll40dCFWIIPMRoLtUPX2li1q2V0w1T7tS02tm10
fVBOZyU+TXW14Htx5TekqRvudTbDMJ3Jxb1+vfl7DJEIdJ0gt9fRSLGj0KUd1ZnL
SnrY7LaRbA8Cp7f6D+JyXC38f/6tK1tquyDOIVRvjz81dVRYVOl4UxOA7U7j6hgX
0jPXOSwwRGrE8sZwG9+j6fUKNoJlmqEMd5gA9syxX/36PRZo8cyMNJJ9n4dRlVX6
fgpP6WH5gfZkdeq8F7lJoe3hpg9Bw2vZNOcnfN+ugUAp/gVQQ3g+jQaMvPRyqJdU
2Cz8Re7bQUeTdVOOu68USVTY1Q7f9GTgRKG2ChNAT8dQgYF95l6Yoz6+/+uM88WT
3q0H4g2uVOtbLgwspvyYdbkBLMKMXmHkzWpAT3+MGA07X7DDer2WhsLEQR9rLjGV
LvQiyC8Ah9fknLCHTG+yPPk1+acqdYmgwPL/cqIuFAk58W3EWSzps8orRbKf53kH
hIqvM7c1ptFwCmExrYRHmot6BH5HCzfASRzl90swGwTt943Ev9njbtHyacpsdXEI
IIhTc62HhDlNYQMhy4aKMbW3LuVGnO/YKjxITHuPQffhEfDtUmXdeShIrC4DzuXz
gRlq/Ljh/ulNYBt2twihFHqkusX6h5RALvjKNEEDWY/VGIxUAxSsfiqYAAtWLGJG
CxMoTvMebGBDIPTfs1uaHUArAzTnLPyd5b1UnmbnsF42Ok9e0w0N+KY+j/j0ckOz
0D/eJzkISX5DDAXDX/yN5gvYhF74lNEn3PDYTtrxhwgQgYq3+BRIZ2iwqOJ96LDV
n8OZ3eA3V1sz5Oe8pPK4Xxgb67F79vo/pDU/9cKHG4QwBpwDeYFyqhKvCOXTdZ1B
LcE66Aswe6h9oAXC3VTcJ9KHe5Fej3smdh43zXs/hWhj1mwOR7QVZo7lzljB8YN9
lXHhuF6xg6n826/IiC6xvwgjmfZREjQxaWcKEK/vn7fnrjuaAG8IfM54gOPiYTXJ
/AcxNGPdL9a3uXBY2Acv1jyBeghB0JHtrTTlGZ1CJEnz94vz6hg1uGPZIl9njz/S
OdytfTbGvdgYPQkuStN7sP2aH4RszVMZ61Rl8gHl62947NG7UmU4iHgw0d3nzYPQ
mwH65MY+cGYQEGgNX/1mFk4tuAMV0k9m8kRMUPEoAsw76197qvT6dYx2A8ETSY05
eJj/JkfQvH4G312kZNrT9jEiQU5rwwpfimYjJQfQzW6G3cLVs0EgIAR+50P/Gw5x
JiSsaBc/K56h/wvnZ7EEJgwEdCL390GuIeQfYW4Yl9R0l54ToSC4Rx6G7dTuynMb
9/aWkUeRVGYzed6K42I95XLn2VtPC/eqxIcuxsgRrjyGQDGcGyrGXgCngefe+ORp
ApGRap/+f4oJx4H1N2iKVQakeOVXQGsTMR7CrbVfg9NkNXUJn87HykJxAFCaXgce
iR2HUT8S4zbbfcebFS2qoFOnGi8fEWMpv6r2Gz3voM0kWCa9q6HGUCws/ECrxxjC
SBD1EbAgJbShAGcUoC+UbVJPFSbxePtErkaFoZ+RTBLAfL/Ovexy8QAG0/UQ/BFz
m0v+9RA3RexgNKiOef7WfVHwuYZvb+FmW4XudlCQMsm9SqvPzTR47fCykYMBMq7s
vJcgO3HNkbPyaVqhL//hbTFOynoeFj9bMuSIi0qTzxfYfpQhQkq/xQ94PBtF/feZ
MV9zjblYvKK6XsW38d1no7vmPnF2yDHdN7DOrjn+d9N7AhVt+6l9s5pG272L8vNx
sHNfAeAhVO2cNTR++H8JfqzTlrcASgqBJ+NINaf+iKJpaFWEtqvsi6e9ogEz50YE
8Y81uykWp7Nrnl4jRYqTnxI11eiK9B3RnKm/oUKfOUODFLwPFhp+MslgtZmEpTri
9AgRdQynZdsMqclcedWAzF+e6kcZjOrtJRD9g/t5oq6IFvkRtl23bG6YqzQRPkS9
hdx5PJ4FWeGVujaSZmMgN91DoqASXbOqwPL4I9KHc0aZ4VTeFg8WkzW2+H8LcGlv
4K9m3DQQv2RzBy6YkArJxfarYfGmzELjk3b6JPJKsRmTyU3xAIXDUD9txGB4J0AT
i+7vea97zPd2tB5QzTYymB9M4ykx/aOb5T3hvzTL48EO+SwUrj2uZh0GxKuECKj6
chpH2ngw7988Qs2zWiDME+4HqnlkUvp5yyzKRlJw+6cKxS2vavp4VBu1fKn4RYUX
RbWbv3/Hd0UrAjrM1zJFGaUpJPaGGiBHLsB+R7pEGjA4AS5i9GKlE8mMWlG5QFqj
5fjHpTVu97Tx1cvJca9l5Md51zFVZFNpI8P0t+EtsvXbYP6EhzaQVemKFm8iQEb4
HT8FHaoQsBOzEHSBZ+Nw/OMunc/GDDGIaGwVtjWqMSXDqxECyJaOUE03WpwFqfBw
/vVKc0MxefcOTOexxIoLs5bcBNQcF1TYg6gAQQmG3k1eohRh3WdzyyTX44v3nEqT
EQkNa7wxIZZ1/Spoz7r3ZRKqq7i0+9/etNOe1qRZyVBrw7/PcOD1hyDC6jl+nR9Z
DnihEyA0iiNhXzQLda622BqCnNLFdo2hfNbpzsxhPz7pg5ULQQNuNX3+f74M8LEU
Bxx4TuBVu6pFZVwYpRRPGnASgah2+gc773d2MWv/9L7bWkb4U9UXlC/SDelpQeZs
OV3mk02TD5h4AmCfkddhm2RbtB5op6pmE70bwaypEM7ayycF8Zg3WGGgn53S3J+A
CXJcZUacRrt7b8fAVjRZeANXSXZswXQlBey0ZSWBihqHcrj2bJqp5Dlf7k2ptBxR
96F4b6ZF4xIwRMMcCLidHvZPWVhhQBRO59eK6ijg2BLo8P47H3f/tLGvJhRDZy4m
9/vR2dDLV/bXqf6PvgxPtGbuEhAMMjwKKioBGWbPQ+20qgWX/ziy1U+rVSU2/zi+
MmywvLqDSNxHLDjQzKPYI8arLR/aI5xYotk7Wj4eLsSQwQyh+DREYzQomyaVsuxm
P4Y+aelqtwl6lu72Kp7in4o9o1LiAIwo5BDVBJkxKpkD9vMenWOTHJzzH+FdQdKk
DfviPANjf5qHltJcyDLL7Y+lk/8BT+8mmgPs40f2CJgL+MFpQGFBXRdwUHNA4jmv
TTgiZsgfSfw2mwYGCgq1vF2EJ5JNwse4E1gw8ItGnM5F98uwfEMUBOr7t9ZKHsf8
E3t61qCfa8vN+EgZ4HxlfTqtS5Rl3IE1aVQwPe5gmmdwFsNaCvFtFyPWVS+siGOY
dc8YH43QTTxLNwHHq17oJfIkRf6lJdisN2B0aai2/6ID2TH/TrRm5VdXtBcHcy3U
RTRZwWOfZMq0w/keomRecV2NenHtvuZd0cqfnZXBR9ns8sobU+iLoEY+UiV+4NfM
yTZ4kUPPFyQOirVpTnp9XAJV043dhaGr0Z7Cbv1M6L3a06gKEnqGc87item68qAK
ZvqhgKU98QgXAFXucghW1niktKIV1AJUR8BVpf7K6UUcMYishPzi7r0DttsqHnX6
FR3fJ9NOtkP3fXLRksbDYXDPoqS8mNO8Ipi2+JLFXGv8CcdQVad+Ei85H7tvKHoa
+qIYMlhrINF5Yydn5dhvZz5iYr1n7XYb+ig2WiuDapb6zPvyYKle3WraVsaUoc56
WdUCO6LXbfWMNVUvp+as0IhTdeb3bNs9SvyxhtpcC/OdIEhwkADEfe/Wfd0OS5NM
TANDAJYdYDddlGhN351gZem3MROaPd6lCnVCxtmeadOWIAvIPLFBIBhFzYDLkon8
O+GycZfFj8R9sWyP6S97UmleIliT+ghnSVpxaqlwfuo6xpU4py/9QfBu238KBa7e
sStrgBICjT87vjj3qYyzu+VZbz1jlTDWqA3MelB8KcKHNRnw3Gu1iDPNNr9N0EVv
HDKxWO6lSSyJk4eqHbDj/Lt5PrQpbUkEWS/wmp+i7Uf+FHVGur8qg0sGHOR3BmXc
ndLGWHTLhhGJQNnoRXHruVUNsAelydy3dame9RTqACRNX4tkZL0hkDvjryfRjBJh
7eXCvzYIG4AHUnP9u7bJBGdG70EP94PR/ClvE0Yp7LuMdt6pVHh5h4OqV8ao2/9W
77JShHjDVwAAJ1nczK3vFsiUemUoJeFvVcBKWv/UM2hbGOXNZg44n5b1GH8Ub959
fPs+qWAxyWvg69npOibAAmjf94bfumEOlQqlr9UWfn7uRLKiaFhCbPvsmh9de/YU
DXdjdKpQ+m7bCNFvEetrDoAHHM41j5+Buc9HxvmLkivgzPGWptclrtxRVb8tY0D1
+qoS4hp30XlP3tjpDU6En5MWn6fEum7bt6drkibs+a9PFyIHVfWPkjUrAtwIGxIf
SJL5WRqaZdjFTy18dejvJBhyuAiY4ushtrz0JL47dcCnRVDk8t/lfWZWwsRp/IK1
AgaFsVNfUkyRlhTEMnJuRSGUJWdNBNTu6PWb7IdkU+jEJybSEjuWVUJy94fyzS9s
AunQ9S/GJadGF66yX/aEaqIbiQfcvGrJUjl07kok5WSS3nZSvQBCxw5rHQBKBVRr
t7OEenZQMGlGloOXthEn8jeWkbHs4H8hNTVebg1wiYYE6AIdtrWHTt5gt6nLq7F9
FoPwwsUyJcJ80EQ1jhpFa9i5CGq5X+GP23ktFTVFj2WqKFAPsv1824jJj1Jw1/ad
gD8mhJDwLRHWEM8oOiIVz3/tRLTlA5BmcbrXTKVrdIP0cvZFruMjMwXXLX7927uZ
lqz6xKTjrexgeYl6KqTem57QrP1JlHY33uVuYxnNHMAfOUGWs0sqokbjyb3jHnLO
YlfLcOxhqF3/5G5C/kpTKxqnpY5jxpSVyQcoZpzR0o0ggl/6K+6WrhE3vFxqUHDQ
PZQoCD+86MXQQN3SSofyUEi6pydS8nz42T6/n/DXjv7t1pTVRuaG53/i+WWhFj/D
NhraiKflc90DtlrO3KtKBe//vrMUj38wPRqyGSbyWr+dQ69Mpa2LUeOrubaVsiAn
PZdePyV6T2DLQH3XOuinokUCAmrHGhC7JJYnZ/Onll70pxI3Fli/joBeHjOOyQtQ
gbsEfm/AF/yBdKxmbMgzJoTeA2/A6eicBonmgUN3jPwVRnCvwadV5EU3favmTSBd
V4+Ne915kNuRF1B6WCZ9BWQNexteKQ1JJuJfLPB8+NoPi+KhLWmMKkIRZhQepSkr
k9PZuUpihxqisLC0daMH+Ah7JiJwIyU4umKiJzZz8SltACeady+fMPfy8I+ZHO0a
0m4aeov17dGoy7o7srH/qL0OJBe7achfF8f2VfAM71nyc0onpitm1GCpOrAcaq/T
iVStOOUMs7FDA2Mdpwfy2u/2hptSl0rnuDhZ1Aqxa0dxksq6eAFjPLWJi6McG29p
6LGIiQYLW58P2THUgd8ri4bWYVwuO9xrIBYTr3DnySi6LivNadOFDCrL2raJEwoh
xoPyXtpRGgYQ5Q91q7dADsqj3WN/zs14BRiOW/X5j7MahVK5BCmtf7FNDNSDjdXL
jcZdIItZySU8YxI0wypPrtfFUvWV2CReCT1l+0CnlUEDzaNr7YGiC+q4gKa2BhHK
dd4VEuuoWxkCNLPmTAa9tmpPs0qB+F2h5UCU66cKJY5rzuymOz5QnPRbLwGLeFFA
o+xOgQtVemEZPiErZA/Csa+jixeZyPBC1tE8HkozM/xaWIDDDzH2H42oOW5b7kYS
ZRHUoYVfc+4kvOw03EH0F1Q2NBPKF3UcjB5DXZ/aeUuDxlNw0jj90q97n3ehO+jW
nMRTi9loeSTMJQKosko2kNE5cqGJGkmdfXGtYasr4ie/Fyw3FAl8sTobar/Mj4a7
tA1rvfgEWdtlMU1+dzn3jiw1bpbnq5zqXuLjcJzD3ap8BPPVce1r2LdW+qBHIuRl
EAV/DFFGW9f67fruoy6QtKlJw5GuxLueGNSE8jC7YK0IsUBB5qAhcCPqUdK9gymj
TUjD40wQvO7rueohGoYL3E8PKjtovT2PDCRiVNQAaOUE9QaX+ZtexXWyplTdoVJ+
2NNt1ZcFIWH56Uy9ldlBg4Wi2zFw+/K5QExVrk3GidKhb9Da4D65UNPYBqn/Jl+P
kj7dpZHzzr/6oO5bxJpLmms3uTCR6UNUaw/2qPaVELEudA68HpLzOBEbXXA7WzBO
5E5BYnAa0eNU+nSAFFHqU2I2C1D3auTjzFCv5rQWBVSMMf05XQ+gcpHPf+gL/V6w
Ulc+rAdp8PN+yp0Y64sW3vrociwvdksBFTsObhhs8Vn5CLJMqLH2w3isGYWIQD77
vP2yrsnHka5RSYPcn4a/JPxS5u34RJLmknDAItQgEHahf12TzYDcTP5tPY1zzC01
hSnphtiE7+904po7RehkZJH8cgloGGAXAYXGDPD9vpQVjX75/cwm3BZNDm/95zb/
DfA1J5YYhnvMp2Fm0C4n7TLMfIgc7mpu0/Qhfi2A3TxRvpvDbDpCjHxeNUR9HUBJ
wmddQxtearBmE9orSvidt2VWb4ztTFYcxHTINUyY4XDFY0Mo7bKGGyXj+ksu+m4+
lYzNTRrMI8ONwvTkVO4x/C1PJno6hcMZd91e7+YE4gJXltY0BoU95TKHsCAn8Y97
EViCLv8Oa+0vqdrmLKaw1nkJxH9suL086PzvVkb/SViqixYC396whvALThTQhXo5
hyds7nJQRds7eJW5xEGNnkwVdMSo96ddgFwgueNAMpAkOPV/XFO/sj6IjR9zJ8mq
dP3ozfs2Xr4vb19Sopnl7UndiuzaebunbmO0sc2t91z1IcOB8mQQMRVoc7mM4Ldb
lbz3tCJuJ33xol4lznVZQIDjzVAo7ACpwKBL/ioCoNRNqOWOdi7aba6urIPviYd1
6nxWVoaiAkIZdjsbHuNWl6tE26MslLy0aht+ds0uc37V5LYM57byJeFeW4dQFV0P
WIqbmLBg4IZzsmkZ8nURcd0v7v9yI+4R632JuS1BMBIq2MIXLZ2d833FWu2zKDcU
UY/RX2x/kRKiFq6uxm7vpdiN1vrIM8yB77eY4J/aJSe19ArYAIeEkd8JLcw36+1v
ZjS3+bvb7OdLRKHRW0GOgPuJClD6QDjKUOZBXvPhkClzOjlQ8MR+Ih9elntm3n+S
HfeRNH0jMBoBQbDREmx1clMe/0x12q3KPwMVDebBSLzgPrg/PmDhf3SsPytjoC6O
5NwVQrR+FHf0Bzl3MXRZsSh5LIPhEaD5+ndyXmVMuxuoevr4bXrW6d3an/ZXQecG
gLfy6EzfznyjFJ7oL1mn43o2iHrJXsj7nZ73QnvNZgPqC827HqD+xpPJlNJmgT9R
+Pacnvd+8oeCEcp2cp9q1b0aXYNbPAs2Zr5uXm+mHH+ax1o8xGUjW4Y9G5E6zYKW
ARHnT41JyuPsqx8cBCrd/pWnPA7SWYxXlhjspbkNQtSh4aPQFZzcqveBCkC7MHrt
mDIR9X06kQKE9UkInwR0kTIRdG7XO2RQgXfDh+wPtDCTUI9oUO7j7th9mcUiqNfb
+W0N5Xf47EtGqnidgg5J5sL0FfcJqSgRMkfFZtFdCFj9Sm4Jr0PFeW3/oWcKdV5M
BXtItbke7OQbJJJn4gCOc7an7i3ln6WGQFWeE2evmrDomcie+dE14T5Bno2EV/Jt
ls0//z/tq8RAETlrXwk0BaxW0qkWbk7Yf1/sY4dqAKqdi1ezzqSv5PZRulk1x35F
LcZA/hF0j0TIRCekZRM47J18zhlCDVt4o7tcaZwQVakKIzYY35n5zy27xnFvowRI
36HgXq0BlhtorHCiQyFwtNa/18X9j/ZboYWw6qrGNwSzptqqgOAcIWKfdGab+FpH
nm0j4gNjxFMlp1CX0W/wAebs4HYmG5ufwkjUSADTgvOGaIutRitm51DJB+3xwQSH
mG7EWY/pyWlNW8UkOmvAtn51euePe2A9s0ciGmVhIXx6XVll3Kosl5vzrvRYj3qx
uj1RgqMZkjtk3jFpEbWkUrob7YYL3q8ivDQ1PctDOruDiYK10kQSx+FdZNnC12S3
f7ftir2FrIcdXy02oVlty/wP43f4jHA1btGEjsvoksX5rLMbkrLCy9SVeszAPU0a
P7lqy9OtVzpdkdiRHi6r0Zyy4hCbofzhmZgx9zLZw0BJ/EOWgS+Rj4lwZt7dCG8g
k8NidOMZ55GPyDD6qyhGpXiiGHiRAoYJRprzzUEYwurBld31BOMVhmXnjZw1QwIq
RoZu8qXE3GLnTFY3Qx7Ok65k9b4sEBp8C50SayjaxlDDtOdcTGqs9mghuG1zJHvH
CpcvZF5FdzpXOLjHB7i1R9vbksOBaLcXjgEdmE6znfIXvKDEMXNZqdpYWcM0XqK/
WaLCLOGQyq/0qGdAmpTeI72zOnMFyVXoa/8xOdQCpEBSW+MwUxecjVPwIJbR1P6b
wVvj3GLL+Vp/pHRmELBzsY+Lj/sQA03C5n0cwmQza9jP3Q69OI//Nqpc7fy4znT5
hTPdUDTTZ7jIRcyCvGhhckTejUJ/doVpRmhWGAtSuEZ4zi/yzelCtqJUZnDGxBCp
MSzTdjyBxUNoTor8J7zyAUDXbuB3RObcEzG0DLnUTB+CuA68FyeOZoH9+yWNaz6f
Zq1Aq7JT0f6GobefJBL7pzuoR5KVBeLWmQccUS3Bk/G0KUM3LbdYDcprchMQXwOa
1HPfUAF/kvjJTu08TYGX7pqjESwhNbSN2iEzy7XClGdUEHllH5Xz39Juy4cDNVZb
5nV3qh2S2EqhfzO+rfEsgb1HKseWm0UbTr+lWJg0Q2nCcwrflMVCbzf4zMj5vpKR
kuJAqXpmvO0E8oDzsGOHVXM8yQDNYiQD6n5NnlJQ7Lg/2OraZK7ddrWbfJ1ImVka
IQhzdybrnnBM36odADH0gaGY0fuhFUAhN0Ny6qtNIFsYVmaFSmeBqqamoGPQCX0B
dzZXEbTV8h7vZoUN0NABRcFx5qXwJR2YY1ay7SVYof5hm900RY3fr51oC/+qqz+D
99ewzeL0pxWfRYfTYLRjGYf8HDqgno5J/zQ88fjb5XToFwk0uyAb4CPwDadcao7M
ezK+sVgEwsuVentB3kD7B6mvsoK98McduVcsIvjM7d+ZLPkhVTr25FaMSMaUlU9q
tiobzWoCPtUHZQvn/NFHbzy12O6f+vb9XL0G0ZYXMy0NoaA5yjfQjrolcqwemYux
8ELzh51RCRocKxprGyuBEcZEI9hkx+nJEFxINPCfCjEcQo/E+YiY/D8RyAat2AXs
rmPhOhTYx2if0klZ9kcgnWHwxo2rvDfoLaTsxu3b4DZsADp4Bq5jbLNJgVJmNBJ9
Goa0hXBlnC5IHM1SIKiJNbngxtZoeGv2/0AfMQoj+WVZhxVgUYKgr85eKSf2IYWL
v3ypt3ie0fGrMoSng0VfKAZ8L0aJTAkpF3HUKZuKsnhc0oD4jMjZHBYfzo2HsAYZ
cmZKG+TPIe+SC4NVDaIqtQ+gvxFBKbtXa6+zwNBAv8Cbz0poBnJzhwp5+qIQJLka
bgnhxWS3+QM4HSiF1N9fAh+2Mn0uVu6VnRPec5KTz34CzUbI/ZKXu9yx5rQveec4
KUc8Gkk6wk1q+Uy1d+hioTm7D/RZH73wF4ev68mXdrP/jroNTdo2ODdKJKFQOcT2
PnxfktO0H/+RLdN/Zr9n5aMty8OTX3FS3q3FjoaRRMv8ndtMz1NeP0/TIqaeCXEZ
6PYrwNpdal2YT/joBYQnybcKNBeTk5s0WRqmvQOliOF5p7d3cuSWyjgiVBgY5h05
pXyOjV4BLNRVnn1E+uPgwwBPqLNCIY09pAJIje59VBwMyCyK/Kvxnfk5W9o45xNc
FrXfFKOuErYkG1jIbq7lIM/L7RlK+oMugjJM0wKEz57VNVlWiSt0nnJjB23dd33L
KSdn47Ypv+Uug/4o61DY91XOYXiIHM4JhaVsDF7upWp5AQaAEQe82DJOrZRmyB3x
rmq9PSKGYO2ETACJMIREuIQqzouYkndFVO8fbwYm+GKGcf4k842PUOqfOoNuYsZe
VAbwmDoAper/un4GTk7VJ4iCId8XK2DOUjeCiwm4wW7f7o+D9qNf9o4jxLfCJvNS
EKEeB05j+atBIW/BDR6/oRtgkjtt6lez4RbE9x8k6rxfEstyTTCBF+QvaaHmTz4B
TVBxpRO92oijWCW8VupsDojQoU4zhUOXuMOglv0kqQaZ7gf8qpqwtihiv2/zzQks
dUzfiVCikvlcnAeRRtOM4K0X4ZMzHQpU5jXkaXaGM7PWyd7MGD9grLCbXilbq3FN
7SxCESZBJG3+xxMG4bUl0H57ec1XJ0LhXHJ0TSTxEXe0StZNxmW5B27puC2TNFgW
ipbvfVk5zMzxa+f09DjzDvSqtYBGZCWL/hamPSqst8lQULBnVX/mgE+lB5wSfkT7
dCxwkQyxKA6w86y7LcVvZQDmm41W1oiPV/BAabu5WLIdGx1oUTtEJ5EXLtOn0krs
XojFov1jhVdLfr6LGKYqZknXZEIvUQOFRrLpYYkJxzWh6z58J/v1jgCCIx4yDPkL
XgvCVskpUw2BCnrAFQhl/98Vh6ADvEPoKqDQxGTzaCRB2l3OyMDH69sFjFJrvcQY
gcGAZ5QkKkjSR4LYwe6M0+Z2MDp4gLu277K+Bk1ul0vBBV7zW+AhQZtI+1H/Adb0
iFru5GQnKhs4DGf3yVeTxciMPyxHVIx4eLy0xsx7rvMVQsX9TSjSLNzrfXKeGlNb
C9oU454YbFeuEE/l8KqgeV3SNbsVsygAaT40wX0afZFCaRrYe1zumDZ1cKbheM82
qVj+pMcjpbBwx9Gy8AWt+GbwjedYJ2qegHYnzcmfCoenYjcdCLCFWFPEj3WRJd5J
PsZWu/7fw4C4/NUUtoI6Hy6hbwMOHZlg2vfVf2Kq4mS9VC5QEyz7AIi4vQFssU8E
ILZQgARAWqDb/y4WNPw8O8gO9/VDLla7nufPmPvRJXH3cpi9ZdSqNCFNvMktNyEp
bZTY5a0GYsbYT57WHUCaXUAttW00soMyR7lU55AESE+IPjhHol3eqQ77aQ3mhLzK
0dH/psP7DUNYgsZs+AhuFuTuOZJfu4Xb5KsxV1q9gbo/qEeYKisNmtXxu8DLIsuC
6rIXxbX/IAZy9Afe9v+rK0QtRea4YL4zHi59rC4BZl2UafFGUh/5ntxZQg9jtT5E
SbmiBFj3109ikq2PEmYJdEfcpNrxK4Pqcq9J5YCb4e+IA9KjTcjYQuCFkfaKSqVr
klt0KRME4LqSJibUii0/kSaJ0VKMBaNMwfm0ZpA++/HCpSxffPOkHmG5GpEk70Cy
Z1lqnIMKnRv80nf/8buQ2/liHsBJ0kPIhq/g9lJeeKLKo/T0VOGo9c7efUo5rRng
ZVCkAN+M04QjobTmzhRj6irjXIZr58zOqRhNXsoIldkYcATLTMMUFoknQfNKUWQ8
OLMiCly+4Ch7Qx5+K2MYVQxq0OBxMQaOqzE+Ms319rTCT7NDEKmEDb678KkoTg7c
zDVBqzF5oHwls/0rs00D1Nhc3G3Izkrbko0JcR3PGe4o2+nQYHBSwrGmwugm0eng
BrtH1LQmXkPWAJVSfIrHqajEdbxFr2eSRNsMv2W37TWj8yGttyG0HIs+8s35vzTU
nqdEVVHwS5fep1ZnW8atRu2JuAEA1WP4mZ/NC/H9fRS8fONiPO+s2Kp57nbydU2e
zpfihvS2/2Jx3XcMXfaLQjZqpcQfeNJGYG6xBJnepRVF22dRGTrkSGpayL4pXnId
ibf5I69/PqfjQonTETO/VqlGOAM2IUUIo397TyD5BOOO3/PYYNI8nD7jtJJ3YnZN
ZqZhxKSV5ktXsgpD3Pd2m/S/iq9NJ3TY1Fptp5B4TMBr3fsjtEDL354pmVdjpWUr
mkiiRRZmfWVog81uPIfGlGoVducrC/L0RUaYPqDhgnhBCx8gnMwsw2bKg83jNRVF
8po+J9+JWEZoAJB140NnpTDe/Xk1d/nuuMMQI0/YeZvbJ7YA4T0bgJ+Yj0qqagO2
JZvRtMp4ERf/0GUG3y5/6yYMotFOgx1a1mOwuZAAg3/X22aU380RmV4vNof6OAJh
1CWqrodGTv+0rKqHnmTG23lFC3f5h5sXNKXM86NEW0ZOKgtxpP6wJD1r4Opb7Ekx
+9qcAzsuLYXRn536yaSRjyyNL8Ybisk6NUW8Kye+qVxgWcX3kTBK+npWqjR2n5uC
15lpjEbiBz+0Rqf4R6WYVdH7jXuMZw3TpMFXwQ/EtqlZGN7jMfb2Hgkf93Cs6rXz
X59/SOJ13VnDoSGimiA73qgttgxzTKOLdwOPty/ejQ4bVyFy75myxnQJC1xQFUqX
o21NlUz0albYExIWVFikJFFAL0AycNAKTzfTQcuIM2rrXZYSvomOM/TilpDXJ4mM
48cmG0GjmhoAsIP1WoGm10IN4nQ6gaRYaOUo1w0jH0LaZe2M3CIhUHReZd6BZqa2
PDuSsyNq03jhZHw7dU+MPLLZXk+2M/Nk7HvCbIWhsq5HOXZxpssPwDfqGE0wNso6
0jYkW4bKbJMSDEjfQWsflumZwpkgAVEf0i5MKnzvnkBD0d49LueMY2EHb+nBRF+p
r3vOpNTdp7ZlCP11iHxLsoJ8Lvean25YI/K/89ZewhPSjWb/THoQazwZP5PhlCtm
bgtsSpqR8Xh4OiFTgEX58L+kdFZsykOi0fFKw4+VdGKRZur5BQbuf2blXtD7Zr08
bTE/hvzaY0m3kxxuZNhxyAxLQ/pEXt6bNsHmxEa7K75DjiyQUZS55aOIGzFgoXyA
hs/aE9Rh8WC2XqxM+djWnxsCGdd47K8Woz/f2h2naFjwEskcLG6UzQ7ucz9BG7Da
BQdgj/UZMFURJXeZVHp9vAu5unY2Y8e+/AiiU+JXwK552jwL2l2MD8lG/HlKQ2VX
DyveznTJPamn5A9BHVsv8Tv6KjplZpDRQg8tLHHpQgG+a27tFUv2KTkRCe2+yLQ5
cUFTB9ovhQTTZ0jDWVmS8GGdVQbuAohrIpwsZKSypAiF6jrDM0EHLwvlvcPDODR8
MYtkEwejj8kyoNQReOCklzRVXZOKw3O+WuGmPIR6YLVm3lN/NScIAW7A9qOLZMbH
jzMGo30zhEl84D6qrzCGzOTLvtvrAcc4feiSOyZV2i/ynCtR5zJTWB/vS6IKU2/t
Q+DFpHIzKo9ekRfx/tzS42o5h7a/C01HcXZOJ5PB/BYye2BcvtmYtZNvs1NmENkV
5Rz3rni12uZGZ1W9G1ztOKWhccFdJJkfY9gr+hL4CuG3OVPLJhQJKqN7ZLOkPIjE
tIvmaFDfY3O6SloBOy9gf3g6Lb8DARae63OCkRCS3MzgCQbXA6lsKQc+XAxdVZ0m
LEXbYzOIZVdjzkYugXznqv7sd0MnzJdGOYA+VHrJmNvKWNVibDJzUSwOzryNxHbt
xSYnWAaCzPOS1B6VsIZVDY3fRRCV7GIHtT5004wLiHEA2fFdDozgc7/jDAImQo+o
y+K9MpULdU+FveMKFuAe8rV0oRf3kGKYR13Nyvl/QzJnXOhFPZFfjsDcIzytLmbf
z1lIWPzq7AVMeQw7Gsrfjyf4uKjlFtUPJxSWruEflOkA3/BdtdbU6nSvscPo+Wk6
yWgQVUGdVleRywQMl/Jln/dF2qpUSh1khhyJNPKWuTOvi1jy5ult6a7OoHT4u528
Im7EOySdSc56F5DBfeH0USwmqDsFlpWt5iSCW6xK79aaYZ4zNmxcEwcB+w5mk4JM
BNjVPhdTGhyVWZr/iK5PKIRGmXn8hvb7/AHJwphlxBIfda2/5JtnGXkOEU/QWtPB
okCAT0qaKjupH5uafqcw29MTLJh3c40IGiQuwq4/wSMRHJS/34vhjJt/O0u6Huhg
EnPektrTBCAMwTk3Zf4DJJeI7pL6ck535VujbWYbqRyaFliZXG8uKgV1G1PgojUh
QqLGqo3TD9s7KIcxfPzgCNy6UCgHRL2lVw5Qn8RT2UCqSluKMaagvVNzCDzy58mS
MynMbaJwi940ECfZoEsiqbTx2M7GZbXU3lYV2R5gZ+hZUcfpFHHuu+gSA69jIpRf
jPv92Pgwx2QQ+o015rceM2GUC6FBH6c5ENuUK9c1zZ1Dgjxb9tQBokAHVfjFze8M
QCVvghK8tQD6f89IwCm6kNgoZPb9A8rQsw0EN6nQACbZ6Xyfr2fwujufWpk4VDrE
b3Bw23qsZx65Nsvsl9BalXOdMdmND71/WP4c4lqUiToehjhuzT7IwvlRSwIFBHUs
amohg6ptvbjT8l/lGGgCkg73whXb/vvn8UKyCanB88VBkFeKdCqmQdYgoP08KDxl
PAve+0hGNs4zITimCN0tPUIs/UZjq+YtUmDy1QMPah8evM54r2DqSgWzopOyiuY8
g32BxQXkD8+Z2/bqzDzJb3sGuT0aviy/KD57AJccSwSj97pusdpDgNwo4X0u6Q6b
QF51P9fa8QHMZyh41ngHSneKSC+rZvU9nqKjyw7lwg6tnXW7s/+MrLjLAtuYMvEK
rukuUOfT98Tht8Q5UQjEyA1hNtpXIOXzpUF2GMs3rEwbxEJ5NmtErJ7LZ+3qGMME
LfQzwExgizFM8Itjn8gOjM5D8RN9maLAhFYWZpwVEQNOKr8tXzF72BqApUi20k42
W2B78MkSRBazsZVR6xXACVxgCh4k/uy0XX3HAPcFDS3ErcvGhhBiAzfTA4IzKQER
R4zVftLkYLGIpyPFCPtiRq01lW7jzPqAAoWVGJ1G7lwGsGzucootnB7r7+VfrXqP
fN+6RHVbS76gdpuKQlE2SO51JAogmDOT9leAI8w6CNu67hhKG4FfDS2woCdyaYLO
r3cHdCwHn0O0b2ocgIBqDWT/o8/gKL/QyrUM4SSh8tkvRyt35vkyMXQUIpjuN1/V
EahMRcEcJQPzDgM3Cqg3WDl3S+h1C/Ese+UJe8GXLo42pgUE8Ojj2ZS0ysrWQAij
DwVJRrzTVRdFbBjSXbr2ke3o5DmvyN9UCyIhSq/Ug3bh7LLTM1B3LSXvd1XGf0qS
bx8s/5X+hafYSuWsDTLciVfCLrZrVjPP0JuNIwXfN6j2ouPJcyMdQ35NAn2uVFEI
oTXsBb3bKsjsdm1RKb2iBNDEXs31mtzj8BNqjBbscZB21pUVFwbDcvZvlnLVxPK5
s5znNLOqI5ifCY4B8AhXGz55UaYZqvpbBNMVX0/sVsBcr1QLODbuWqE46Hy80xUA
RDeUqMk+kN1wyrGdWVaDbe80BMs6YFk5nV5qDOg0u5WkyeVgQA66k4ONw7CxMoqo
uc3Kv8muQ37VPvAF5Nnr4Mp5X5l4MR14hU3HwrhoifNGuxcwbx+k4PZd89uqD2Ot
d1cYeaXf4BPNekGvG/UJgBP18YA+9v0BL7WGRKtNzNju/GdxtHWzMPS+ioyfEuHn
lu1cRzLjZkGCw68xeIjZB44kqG0HnjayFt+cl1YWNcTtLZKqLMFjeinBVHcFPPzR
LqL144CE6gEFAj4FZVFvDs8oOxLiaFoOhv2uzLmMUE/Ap4L69lKqGe2D1lGLmznm
EWNecpkDg/dmI145wVM7woi8ZtGE/nYIH44yinJUx542pay9Wza9ahoDBQMqQfoa
M2XBAv2YxUYE4NY893P0xBuj8RPhFY4NpqGeqvMk/rLS0GBbcrLtMxhweJYpD03e
2CfZSbaIVszT4Rsn2vJTk68iNqAk9FDLZTxrRN2PkvFEbfidzc8tbKlIUQqF6Bad
sb5RLIJzmXT6PFzmxUqh+hh4hFGuNLTamcgmfQv9w+erBrl3JPHPJWY5wAcDez8w
Kd8iemCcjLKIDLjuXeCezC6dEDX7NPCdudiLv1BXJpp+CpZAvnrDd2VMMElINezz
/zTkExps22FbysH9YoHRVJToYjt504Axlkhm80O8HSuQjXoD01PinaICDNJGfU5h
nelq/cTnz4dF/CK0g0WSHDf9F4WIc78AQdBm7WzC4Ec2mfPjGRW/0tzAAKpMCAG/
xs6sgUsjdbekAznybhYdtllz8qwOJKy5sw5gINHkBXs1H8JrOpke71Et9dtfFoc+
L6sU2BCxsTU/gdoM+SuO+Y3BgEB2T3SRTzBClSOxnedyBTb2lgoVtcsC3Fw1+ARb
u1+0zlUTQeDr5LasR76hu5XXnROgiH7cYEVi3DZ+382Z2G9YQ89bl60VPg5XcUiO
WIzgCtdjfMONFv2TPBXrZfxg7IbpTFtixZYf25OGqnLJ6MKop2SXhWeVqkmy+J/5
chYa5JUWshSoxNxquDwHw1bpxALgPUDoQNRyCWqQ+XrkovJjlHrVjOmeISWRKR2q
y7n1AzUASvQmKbl3Q3ttqCVZMweVPBoLd9cSp4AHVPo2t06mAyiwrBMwfASUHzxl
Y8aG1XLYGHtb2oHuQk2AOfm8aImrJvoTO+LwU26YK5gHhyc5Qb2/BezId+CXpoZd
tGkBq73IVxJmstmnezUE1DQiKeHg1JGEEann0OB1XUD5+25/vUYubj7lhdSzXnFg
8ZxuzSMARmen2rsJ1FHNktQ1ZR2xrY2n1lIAgnTnuCw3nQijqky6J6SOOKO1muEY
lGy9lNO2SGryDXX4Riy+rvwm0selwShISq8b8QXG1YY/ChN48XOfZIcXgOrASxqG
63QeKsjD8cgVk+21EgMgEo8IM6Xrv2ch/VBCJ39qMx+QfIYICYXziOeyV2Vv3sS+
6dDV85CIBbh7aUyVGHakJ3OVYfSy8at69S6ugurk0PnO4Qzb/FvIVboiwrwFxDIJ
JTY0MMuyOrjfw80yvhiDAIhg4bHeLoiLKblcvdPzQSl8qanhj0W2FBVj+XJNboF9
E0TOmoqdicQv9Cj7q/rkGZ17GtXlWNCaiZYj3PHbXjKkZGZxYxz0g0yPgfY1RDFC
WTxMW29xOJ/9SDeODdGlroa0StTD01KdqqyDR/MmIWNsG53evVDwXp5ASiemX1gH
AlJKy6WcQXUeOuSBVuPPZ7i60+1coN2uxKbEsx1jB7F2xzGcB55Blwr4vLNo8skp
24xz0c45elrgJkOHiXq/Ic2sjY1+oaA/85adp1xIqhJiIE3qdOKYRzW+NxwweGwg
nPGVrwyHrmhhLorYtVR0z9KfRf8W1hxkWORO4BcsVQSTlUluN+yorMNp19uY+NBn
we9LEDSv9sWgp9eU0boD7/y1e2jCOoUP4i3C/FCPYzwKYyf+xbMdKmVrNZ70ZQTm
c0w31fGaDPFK2D1U8/On9YIuWq0H4qnaw971TO8bOOWkwjgDlFP4cXz3DCDozPqM
lDJyaAPHcLBttKoip4MaMK35b7GAsusI033jvyG63bdIYBIWvwCcRx4Ozlq/Fd1z
fSraZKsGug9RVY8UL2tGIKpCzUkB0D/vKIf3Iyhmh0k3kVVkcdEJT1N0ec4Jyc0v
19kgcwrfbYaOSXsnmX8gw33+JpIcI9gdGOSiQ4kUhLwR+K/ywIvyKbUc2riAVxkC
vw4TIHJNB/NqY7grYkIfAtCVztVKamTS3OLDc+dbUdWhKXGkzTRRomL2vDUL8Qu6
040h9pjt24lPhZ676dTDnnR62MTa5+dt6z4J0n6wALyGkQ+n+r1Jqv4yGzaMjLMB
8bVObsyqL7V9VGCJwXgqmaaRCHVSdI0QtjXnFbkI/nyMdw64p9Z3ScJhTNWDSAw2
Zi9kZqReewgsaAqX4+IOIXncDmMxqEjcpC03D9RBV4zzbmxKGGiwqvtzse3eu6I5
UqXae40LB1aP71UoFuDi4TuH/3NXyyPJaXTzTvpbxX5cqmhOFWQ2RdLABuYrvS1y
rHA7h74ex5Kg4s4SB3iBosNvoPCY4lip0Pkwfu0tnUPj9zQ1c0aDLwjMn7va+MJ4
KX5whlhHJ2ZIMR6FTxm4gGc31Lh6HMw6YbK4nptQhiVZenpost6HODWS94lAFcYR
ot0rtHiAbwLhBc5pkJKFPWDBqtREjxU9/+Rb0ZUG6pdrgsViASQybxOfqSY3GZZA
DNr5E+ETpYZluIID5ejXeriqsqWVL04v7vuAVITd0I6X4b9g9h0/52C9+bq1cIXr
QL/djxHiYmw0kB3/kE4x9Zrrwzcjyof3Af4VDLVsUrV+vAraJ8BbwTk1LOlb/XNN
SOUyclgT4TOmdfR0N4T5i6kVqxty4atIxrkECamT35rnSmWP4wNrxgOd3jef8FG6
d8wKoyu1pVviubfsP2FUGSxRR84yn90HHMoxx2COsuKmXQsNx0q2dNW85RlcG3zb
1IuISl9Woe7DDJ9L70cJvsH0cLfikRVJlQDjJSl2SsOcHBSzfadGE8d3YPRPcuFS
IMnz8WRxN0gAlmWxiH0FeFYNhs5JEWZgUJQf6ADy75I2pYEZC7VSayjjpXDYAaL1
I2mXkwpcks9gZZgvHQA16QkFif10GKMvDoM/tcwBB5ofib2+arQjgtTOhOKbgDAj
NHAhwfjuM/DRXPLkk8arIePUzhkQ5BlKrFDyxYAP0TD7NDFRonudBgUdbpDfCzyK
OlatWHWVV8US5+K01uzFGuf5xxQauzuoNf+gFoc24ZOMNg4+z575AJ66D0hC9vT4
Yrwj96Qx+MJQYg1ozID79qEOVys1zm1z8xz88sgYqD4f/u7AvOs+AZbhj40JWgzH
BhE0vnbI6NXihNsAwsbWVSXyvwieOjArw1cCfDwcKzWvxGyvODcX2HHKKz0bWnrI
XYHpzp5IgqNhR8QJYwQlGafikQKtiDWQxLFQgmF29evBXk92bFFw8goJ+JATnTQX
HzDMAf0MopKRSp2lYhEJ/ueA3NeGmIsrR+WU7mQT1j6J/bUrgi0rK3pb/O3vFrKa
XvgreKUt77oGIxxVLrt4xykfebCkaXTq3pfhLScXfbQYZLXMGibII+Mi+Ln3jF+X
lNtDDjghhZl4MEx0xKoUibIBrbm4XbH0zkt7cLfYVsN4F3jnM5h1aB7M/6cMHH4t
3zHbOktqSdPAUlbb6+AcTEJANRy4w2qSjQ3Se8SD47/c5Hg1Pc/C9yo4qyojRBBp
zYEkE4K/5bhFQ3QvJ9XWJEVJHOBHnkdFMhwe0K9aZgLn6z7FZiM4QdhhEH9Uyree
hFN+FKOjzlcQ60xizhpSBBjUYfLfUbkgCce9PXHBQS3eDRDHGxyVJh5932EFDhkd
w631SgX/cjwsRHqXkScNQIqIhXWurB4clsXBCVV1G0yKyTQHB/DfUFFF6Rpf5Yqt
tkH82diYq1Lr0mQYujXcbn0VUrExhGhrSGHjGLWLlfby5VPRQuZqRJ2ZfVZyYnVT
kMJfWiCW9g3dm5vhDOeFM87KXmQ/VCYEYMVVLQ4gblr9NnTQ7goTg9jpgxs5jUKS
5+gZprDA45Ed7kNf4Tf6eLH+db176rIfZNWzktrk7Sul02kyYPQO1tiN5g+c1dCE
q5i6f57kP/Nn3pxhDB4DrgYMlrf+0WyGqklkGEXdYvpeJ98P+aX0yyhtSLnBerlj
K1arXfn/Ka+QZKFRp641BhWkv1bcBfYVD9ptbwIWCkx2pvs8Vp8s1FfSNamzYLIP
VIBiYG50A0U5lnlipxV1sOURSEQ2QqfRAk4IJ9WllQ8PiQLH1tSDbR2chtoMcIFp
wiDkSIxwz2r0ZhAc31lDThhYfQSV2mMPg2iSH6ULO0kKkWC1CR2661vRf1X8pfCS
cIwgAEVAoCYUCORw/Mn+dL9f9a+ryV5SUDKOhV0p02XY/5J0q/irNqFFlB83DDf5
/QVATVoeFI2zH3vNU0vT2wuxcJhid4CxjwohlPBILOnqr356Xy0qopLZZCUjt8rU
nIUkGOfsijEj13Xk1m72B8aaFRbmcyQ11W7FuhiAcCbd0y1Kj15ctqTcWFmVQ+EP
WZ4riLxuEOkJq3A5wHAqRgPtGtdz8jaq6w9WrgbUSt+5QYqXWz4CV78GFnHXBR3i
ioQkNCB0QGlqIsfZi9+P/MGQMg85wzQ2qLANnnbXd+wm3OYyiS9ebOh4JCMa4HMV
Y35qZIgKF0vLegnXCrKZfSjmu3fB2uwoPXZo/Dt+ih/OYG9fD9ekm7wv14oOhQQD
TG/djEtSeBH9b6l1vJiGwHDHaTyCfVnFPVDFbjS6vufdZDuSjmRPeuIS1FaTaNZt
VlHIHtu3y3Sz+PBCVwf8sD7YPDddrXCoGxr6knatxCWBgqLetkwi+8+fE0b/LFSJ
9Yxzr4xo87TQUi0g8izLzmPIzMqVRyA/f22WULGKgqP/8BcpMsLEEvwjtg9cRWK1
AzGH+xxPlJcFIUCTvQZLdq80CXi37lEtbYGYTsEzn7d0+8oi0Rtnn7GdunaGkjOB
CFRaAznKmMcJF0D5fIgzy8p44xYpeQ64VYh01yS4se9pq80fBPBIInpIjotKUrzt
NeXMsViZGNm1nxHaZlPYqTrvR6qiEbZWlyYv+tFBXu94P6Fa2UlPRIzHbsHALl6h
NYhuuIX3WDW+thqGf4wonX+nUbiI3s1Q9JinzKg4Xyhd/XwOSLL7CbizpVbV8/8z
fDZ4cOPcz56nGT0lU7xiVtBymXmEwG9av7nispHakwzL3AVhGc4s9Oe1rc7iRUE6
+9PxroQOJX4+kHCuxfcvRtqQL+4Pl+QT8cJG7WqJAyMf79Ojd58ME5rfV89n6L/U
NcGDsMGco5ShzybLPPDrfUUgMsXNiyvB8btpzlMXqumoUnc9VQvJbHQMjBrW69ka
fh7p8FxWvYf3yjMDIe7eQVWInXhTNsvLDhbhT5ZDFmmTHbLpAIhLplEyXa2i/6JC
KAnoy5RMkdaJCQA/2eNQha4yW2Owt+Cfqm9BAfe31qskA50WQabZ2D4+hY4tISZD
o0zi+QplLJ1uFiyRDp4dRgaVwX6280lE5lFc9rOLlejAlpJR/b3+eIAOFjUQ5b/l
MN/9SUpRmUXd1SB4Kp+zxwVtz1FvlcV23mNTvC6XZ7MjO5keKvIOBIPDzUaMMJvI
1iM+SBEzsYoAxMXM86BtHIxMd36oixsRtWpYpNroLAWQWu6BSiGoFnThjHzIDLAK
N88ZPGbV2Wpn603z48brZYKQS3n7GD7dtMK8xY026HYp4XpxNmJJMjnWraBtTPxg
0nSvp9w+jsVQsSZLKS52absUWv7Vi2Ps4semdCH9e8ta3ttw1gnAqUoIQyYroMhT
l3A6ZSt/OUW9nbaBiWG6srDP83/T8nwtCLxt+qUAYHb4sgsHYogLmuIeWukTXE5U
C5zJD/bWWUFq41mjAhTBo9+203FW79sIqnwuuaoHUMeeajGUNdz2TCRvqsIJohZB
sQTqGdM4YefV5FB5kJAG2u48gqTe2S/eMCMgQk/yzhDW1hfARrLtx/h9zOTh+ttf
GpTiJhU9UUHB4xyW07CWUf+RU4mcvBrEkjD+F+SW/p8MHBtDBtbaRnYJMAdp+mdE
tjCGwq1KNa3vn5szIFdUNt3MUimuCmVYpKjFYKvN9TaNuC3wNV3Xufj1pRxPY0fF
GM4tMm4tRsSOnMhNOa+HIrrA5PIJD63SDMEEYazpDAxH5zbAUl5Ycb+FT8cD1AU8
rkvV0chFaCqgoutQiklqjQdol0bd7exK9rmcx28QzYwLScXZgTWn+GMwAQn6vdqU
QHpfgIlMu17f3BA9cKQtS7+Eb3IrlNNLhYWJV79W2eq4Oo48ecTVTpL/iMmoct9z
cJNBd3lePigaisq6WLFrkoSSDGfGERzpzLNOTEQ2qaElRAMiS0JxPWcY0tQtfRLe
gEZonVX8RDaoF0T2WzM+LIAOAnxleGh5oDVCzhxpyftMunojT+jlaaDFJKJS91Mq
WEhJudu8fmY7Qhbm8pYOtJvwANhiI9qfzf523NZHMIse1hPW9MVkNlwTA5Frp9ij
E/qe4RBu5IeCrQJfb1VzjicS4nKOlyb7UBjbvPmia4qdMFP12tASyBG/4F1YWDDq
LIhpBGnV5dyuH4A50zfALeYwvFtWF6/jNLxbEtKm9bMZBo28p0RPXQwHzFMuq63L
2wzJdwCpy9r2kHZ7N4Keoc82jVU71/oFSd/1HZMyUBvBXmQCYeolZ+lR5dvAlQvA
08gHqQHk92mv1J2p8P7UTrciGDjqgE7d3Q3hekXp9kioHsrvQRmK2PuUnO1mmHa/
yBqAIfs+6YQuEiV2Dt9GFjhs5v7jk+iqtcbtlNsrtA+NjFVbVkzbSIl+x2ujLAPI
QcJvB8eT5GyXZ0Vme7k64QEoBaxRWfsCn22f/VNKdkO7pIyD0u5UfF72cWzPnSG+
Dh1FFnn0eMSiThCW1BgL4Nv3EqwQghrnXEuRO4MLcyzb22lsijXTdJ/2ZQu3IU4c
S+9xQOvHZjpKwZJUr+JWGYaE4ZI/zZaGBKJ6k6ysnNxks5l4SHPpaCsV+Atru6JO
XksvGLoSpwc1WcaSHJJNVtLBA+HDhl0s+1mJqTdTRwYOLXaF2E3VDuhmVLlE07p1
unglt1QNgcgHdJWMFSwsHX6FMiWn4z99ouvqeMrL4fs/G/RKssdZe+QqvrsGwZSk
OEuWR8HXWOxFL5oiaOrnERCiHkz0R+41U/5usoMxoIi5vJ/gBJyJjziruZRsx0eg
o58nc2+VYRu+JY1GT/kxmdGhbWoaL12j91EV8i0IE63oW9k81gXlyJiSLmEBO6Q/
buTYS2xhOfgsrRV63e4huhp170NBfHDfyCg1J/CXGTio0o255y3fwmo7YhdPYs28
mVtes7OKL0ocwcEuG8WQLyCFCm3VcR1D2JMh3ViryO/5Ynrz2TFaqK8iIEZvbHrc
8HKJ9vri/x2X8r4x/oxzFkJbc6Amc3Nz4lkx7A8ktYi1ebDe4Wpy/CNbSW/FgHQY
r6sq+GkIiqHnRCDSSPXTSQ0Iq0i++YW9Ie96vLdi18O+LN65lmR3TdHhKkVC2eCU
u0nBUuKQWkRVLXySwKT0Pckwm2WSEq2c5GDepVhKKM0epw8tqRkUXEkR0cYEc5HE
PG6Ft3/oWi03S7m70uKP9dciWm3ShPb076ZwLaoLEgu/LvRk8dhdeSVjzW1j+5ZO
IG8HA1wWe+9nFSx+audtVrs0nTAbM6b8837J20XkiWac/9HZT+11AkLUTEm32Vak
xYWqA5M7yaPiAkOEY9ljEPj4dX+EaJZo4sxHx82IHunZSRzSyVjZ9ak3D3sG3gHT
O98a00SXKLwogipYmNtW8X/MimjJ1mcO15cr7TFh+IOmuzW5iXln11dZIe9BRx+V
xSY8hSwK9fy5Bzpir3jV2Ep9UY03Ki/uKIOhcpNuAIodB6VGST+CDpbukHRHOZqo
RVwqkMh7c/fcj6LbBijaaWIYuSnHmy0kfY95JlZZIJd05SwwqS/lWQjhhKSxi1JJ
FALpSi93E7iew49CEe+Y5Jo2azJPM7qk5biltt/fWl02IRxsNf5vdJscxOP69A+9
6u6X/qmxrqFEm9vpEUkVqpJBVorhfp/MqXq3mDgrPwMAiibkB36bFskfkwJSNRaO
b5iSLYrnRgHJEzInmoQ8BaXq7OHdBv9/LZDXD20TiTJIk6feWyuo0dSRyzk8MYwh
9QfAg3aqPZv0yuDlMJ260kGqJcU0I+JqRaSK7ODg0u5LHSHWM+5/ls4cM2UuTBf0
DvoyAjh1bojmdJ7LG5BFcEupbu6YaU7Ncx7QHFeFXabK0j/PSC91WMrH9L117tXT
Esvbl45BPogzNL/TdTq829WLHuj4C8YbyIVTFS1SlYflYG85kuLMhbZl5k4r9eU5
Vl4ybQOVNvla0gjH0vS5i78tTpG1PHFKY9LDjwClY68pSi6cl+ZUdVHvj40gvLp8
nRqIEfD4B2tGkalqHopq9Wz8aA6O+OIb0+NpaM3vMun1S4CmYhvmPfxJWg31PA4b
55QXXMmDPQoOtQgUa+4SniLUmZtSWcAWMTv2eGJG8/kXLxxfxe8EvuRHwfjWDfvW
K2Q9P04BpZbfCDXO5s9O/VoktQ2lmHsQ9VJLtsvUMeaK7hnIdHx/WT12C87JPsAV
3RnVcZqMY50qt2LMeRml/dgPb7vfx1DHbUjrhWpzsJsAvKSIds1xGO4m0PrRWI5m
sucrQeJvkzzK1Y1kp2yvrJ1EqxTVfrso2Y0uoRbcysa36hOPQUOUHvs78Bi3L69m
rOW40H/ZbGtEM/UjEGy/c6weNGDFcVlPjxxV3Snr1LoX9KwL+gJQME5oEJ48fmSf
PmCH5tsVoRBiQDNHGBIlYq+KCLvBYEMUGGMx0Dh+Ve75U51LiLAdfrMLPo9259KP
JecMcKnvk6IWbAU9jVLOvB6HRxicP6R7sra+2K6Q2Mr0Jpjoj7FBZ9ZsbURVRkwb
pVT6eCw3MO4hPJTZ3/a/gJDE9UYtPGP9QjiCQxCR7UD8M4z6lWNrvdvc2ql9m+Na
EfrTCVbpgQCI9F3GCIxqYFBqS9fBGgIjxriAoMgIDdwtbYJAzNICy7pgXc7s6gfx
YOLjLkypgI8JaaR7fsXStE+DqUC1nUd2tw7OQzAlKaU6q/oB4p+WHNSheWmI1mYN
ck0BkRXUIPSAnyhZ7y4QhW+4NcaKsaUW1q2BXpyIvcojXq+ITcuiUA2/RLnek4EQ
4PW1BRRSnBvFkb8rekf8W/M/ysLaaKNp7l9vni7ytPpLkmDCHOQChpC9PysieCM5
PlBVBCr3FLRMjh1r6x5kPPEMTFGQTftC6TXEwRjpN5ywJi9vOdm6auGWb++A/Jl6
QAbzQ+Re4J3Tx8ebkZQWsGfGDgd7zxkkCW39wmifmX2TwoL5UFR4Y9EXckS6aGVF
JHQcwa3RWbmB9Sa2s3tFZe2jYs/RuIuxSYtvJPglB1vOQdeXANrmVRoAtlbSecSu
7TuDICvLDTCDZl5DqlBGOxOJbRqGbZ3KvOzHDFFGKKQyK0DQ3Y0g7J0v135EzoSX
2YY1vMJrTLmAeRlMyuQbxLg/3yFGu56hoX7qOk9fDzFGdoFLMqBqK1n4to8Ylnf1
PNK0wq/Zh7GLK4Ip6LSGERQKJ0UOqsX5DLzVgHlU6I1xJroWv98/cKleMeuNrF8U
JmJsb/8jaOIgSafrsvFs2WVHsg20NDwqezEh9ZbbDtwExp/k/qNGUUNgX73MqozD
cD3/2xI41ehOM1Uel7s5ylQyNXrUP9k7qwg+Zx5t9FlK1qagnNQNZ/ZFStPPJIhU
7XVjLXtThud9MPiReNKUmEqOhil+Qh6dd5N+bXXyP4RMmgHE9bJe854xMToB0ef8
uGiEJe1NoTC3NK4Dc/WjQfOl/qDcI0ZhF6vewDh/0YS1dmVbwDu6f9FU9+OFyjK/
Gnp1p5tUlO5W78tHX2Q23t2qMLj7iqGFRvVXB3v8MZ7v2NPvboQkRhycJLsRHsc3
szqyzzOE7RQZcj3vhF6NgB0XZK3x1rm4FmLok7Dp6/F3m33CfDBr1jeb+nsaBKOX
a7K5Wx6nZVU2Wk1pwMevpMMNB/hs3uJLn3riOgbbkEAY7cZKmx41Li5Ik6Nvp5SA
CkYZWp53AlY5FVQ6uAaLZa0LaMXfaJHikCpYBiAM0J44vS6SjaUO/reL+zz4CCtG
uh7GQlsTrIcn2eje3ZXuSphqrRw/X1nrh4bHzv7LSQAWRyj+Mr09vwFU2NSXKsSP
FdOZNn81JESYZM8buM7g+DQbtHG6k9uoJsZgZQl5El2RP/8TM/p7c4KXibyCMyj3
aVlIQd9IUCkYGKyNTz4WGjXuqoEWBWC5rNQ3j1rb031F0VT1Lj5ZOqPYf8H+QMm7
0n9GQJQfdWfmHGaPEUMueFBHFvOmTQUvrg9bkK/ef2ZpE8+p7MyX9q3x44KLuOx/
DBe5O35Llv3pqPKda34LAVhB20vu6GuTOPoVx+0ooB6PwZX7I29oxCCf81AYUcx2
ewmlluCohXMlvJHCvLeQHnQPdY6rdyYt8B3jhV7BRL8HeH3aJY0WcwGOigPQVtmC
JAeWpQFZ/LGKr3Q1nzV36mZNIStOOFRexLKLXoJguJjPp52uuSjxZRS8Jk2GJ1jQ
8Kpp+xbq8BLZIWG0tkxe6u2MJMvpo9YqQfAut91hxrVZAK6Vi70BamD9op5L4mwQ
GZ0c5PeJPHE+ohn6qam6szNwIsnHq+6Zvw/tbLL8IcadtPQmILjzwPqhs2c/JMr3
MAxOIS4gsS67cSCbZVgo6QlGbECkiGYuN5pCeVsy3FSSv71Oa9BcfL+4bjNBTW1x
d+dGOuMDxawz/ye5qyFb8Lizt60u3AAgVIxhOSRuGu5fj4malD4bzaa4QcOxzHY+
KozQYOunVG0JlJP11g6DLZFuVQR46ODXdynlsD+wXAy4cgU/JmDhlIW9SAYa89tI
Nvj355I4T+ehIjn3zQSV1zqKq/y9WT27QKt5NdQY1Z3YEBwiiBNClDNuGMq2aeQA
//fUkYYmMvI/ak/rMxyKNsO0dNFLXVixdamEwybw3Y1MzYdPDFJJf3OzXVkX7SpW
JfZ3iLKI2+JG1hrQDOnzDs+An3jkVGhTArg49DV8rJBchBRwka2LRfb7aUHOI9Ax
9heuCL2mkK5nmABie07PEhDUkjc4nPk3Li2oYb9l7duh1rrDmoAwlxCYjSDZaF+8
oXItFNn1leO1sarDGe2HKo3EqldjNiKTO6PZlvE34MHYlNF8baLsb8N+CskPnUlT
0iIZTK07pdItUjQBrGeB1jq+seDk64RY3fciMC3LP8TsS39rqBQ9/vCcy7FMqA+V
df0liaWHPvy0Uq+uSBEtFDPuKeW5ViOaJguD6e3mjZ+2WYztOd+BCsvx7fidGl1G
LdEFhreLUvp1eyjOn+Zi5RyXVGvmhIOg0dQsvHvfETgi7Gnx6cA/AwTsCmg3EEOd
CxLoKZUktX6ZJF8/TWxPUh3sl7MYrFqMdnU5OYSQpj/eDH67H1yk5V20PzwFBeLC
URC7z9xC1WukkBdtYhrf8UDJ6xZ4w5LPA7RxKak9toyCaqsas0N73kCvtYqBL1cn
cMZ3Ak518GKAaeE5PDfhET6AbHHyOPljz3fQA9mhXL9b8aZrjCNG/ii/n4S/IXi5
bUOiTBdSdUHAq+sKiXHrbect9VKAGgM3/Ug6Eg5rmp6hattKwnOHAbk7k09OIh1u
8w+V/EKc8x5h4fosYpe8AnAu3ZVJI3vwaoOn4mqTtgHLozau1F0SyYzF+3O1ruX/
h8uZfS8Qo4C+qv1PDLYeBBtaILcrY6GsGltWOSDamsesaO+fD2tDkTK6w/3pEpK9
N6suHnszchtID01sIZ/t8x1Kv63PaenzLrZ/TbpDuSyP08995ar+b2UOftw6Feqr
gqtK7/+7EdcU10xTxz/QGHIeDoUpHWdPHX1LjYHRf/ib3RlYTy+6ah3tCddrraWC
pxZbOO3pkVd7qYXVwb7+a6ExSgyGutp+ZmVsFpJ9NeW1I60Ch6BxIYScP+bGKyC/
TkOG0pbCHUI91glvUpePRd8k5X0AJCiOO77drUOQ4uRbHgslmHPr+hTvIwgGhzeF
Z/PErYEp1qquMmsZxA4nOGDvd3JPWmRWZdKAOl/arVQ+//jIL4Sdvwty1ijbmiuI
bj60bN50jhUV6ByAukq01x5PO44KGDiGP2PZ61rGpkigt8ZacYuwPbqYnNhQwU0W
9A1QC1BwOsUX8UBu/Ge7+u7Eqn57wIrRHjHNbar3+nPuHw7YPPnGdVt+DI/B1QPQ
C36X/vyXnY0glNQbscLta6WEJtlKhesS8HYEyWQz+rCQxTx5i+tOUQB4Zu8a1AbG
abgn6qDbPaQ3vWWmDArfVWqEvHVOIDp9za49sRi4vjogdmAZlaVkgVfP4w4ZtVld
Nsx1XDI/EZhKjrWjUerqp8odjbqZq6aoZySZhKy+PONHW5X6NAmmdCc2jhGO1y48
JbRlNNNdrmQerB1meOQn8187Czkt+rd+kVlsghLXgzu49cW/gDEI1YnEEGBRT+gJ
sK9fhgntHo5Yckl1wj/BIABzon+ABxnYdBVFB+zg1zA16d9xPFuFmKUUlehAQyn4
ji2oehxDIsF3sSaXkzlwHiCnalPVteKA1JgE77F9+ZLqup3qFkJP4KiA7QTskN5P
w7wZynVRMqES2yczOzH0cyIxBPvQhr5twLorVgAbkBtw8oiS4UjA3fzeIbiZibUz
e0qlbLjpqbxRc1IzLLutaSw+UHzMqBmOqt6P9pVKy+29P62Lya9i2QABMN6C7t5w
E4hw6iFXXn+g9+RoiEiSvpf8K1mZdaEkjJXNww3amlJ201DNyu2C7naRtC/TyfeY
41ntowW672WjTz/sf08v8Bnx1JXIYojI8XERqKldkumig6djn7n24bTpojqse3ar
W5QW9yN+k72GqTX5RuqZ6gh4IVpppDpLoa7fw4msg1KPEsvUA9DUzHH6ns5qUQ0H
qaRuOfAUA7JISigbKED+9KbDCGN6/zkIvw05xDcAisrR3m4w/TT9iFZkutLyDtAB
sz3AlxAonaMD5GLRaLoob40M3KVMPizZco3W+YspJppZ/ngn0dF69i20Gw3glHf6
gnCYKiFctM4rg7PgOFR5Ao+did/K3TYFJUj9n0dyIl7bmdUstmjfhBXZjpnE+9sc
e+dOi1TbehJtIXY+C7AWY8745BpTO1muj1Bsl6veUiPH+YSOMdoUhbo5QlrFNCJ0
c9+R8Sr4AsF7i9kCFPBVn48F0kDuvvuGZKfCiAPmllOFAJObrY7kezcH1QEccqS5
NExcLqgKNfogH87skDIuj8Abv8BeQ5yXoaKTRETrEzEcLns88FVxDncMGsFP7gcA
jreVcOyR1dcluf6iN/axSsJ6+EY5qOgjUO2cOhVt7BNBhft44wHE2sOebbG6SLE1
v6b4oqr3P2nVa7axo+f4LLosvJV2KmmGsB27a+aQyIk90PVE3rNHGqSU2wElOfYb
3u0b3SyAKQ74NxTjarytz3OO8MEXxLbVUcIIctjQhgi1+TSpLv1TFgTXykbq6h91
h4l73XgkRXskJc1zdF4E1jGfi8bKeUkAbbBbqpgFTYPSAj9XxcLHuvCh4Kf7wI92
pjRpx08cd0gWq2GHexmk+47eZPQyIeadNAfY88ErQcBO+U9ohCMvi+XHjSckSplc
Tu8UuovjyE/AQMDDYvZbL81VBZYoSTrv5KBCwaRhXf5q4d/oQ9Jw30eCmiNCipq3
IlGD49Vr6pcfR0MkG5UgcQ4vhWEWvHX8TD/TOtV1m1/Qxb/E3a2lXB2qzuHt1NaX
dX9xzXreKgovYmJBtAdvbqGgaWNNue1wHQ0wEwAGWt7JeO7CZ8ntqmPqgb4GgLUL
oozWJVAfSjkj7I+Ki3WnrVWsR9Cnh65Jc/d1ArGdT/r9QFiPFup7Tm3lneiamWVP
TpFcMFN5LbmEx5xYfC0AXR1tWy/R8iuRjczLeBOqb6NNXEYVIZTn5q1UFhtt//r9
VpEFewoXV7BqdK+uyvWTOiLdiNnb4VXp/YAywc/BV7cadhfMT5T+yTQzTspQ/IAz
7W1KhZsQ9Z4DqQpIaDuZ/iMAbzX90/Ln9VMQuQ0GbVa0fdOf2hdMzqadn/umuZpt
5wxuOa0bJVosbXFwctra/A7qEaauBALhJJGMuCILOIUfI1RQ6r0XQIqcPkbH4y0V
43jCns/pcJresTu6SBLWjgTH7P+pkIdVgFx4QzUH2/3uUaUxLr4wPuqY88SFF088
qOqpbypOd/FPw3bzMvBgvKMuUTB35CFVowxwt2/mxdGIOM35a1rvGlSE0BtmXGxs
cnOHyYT3E4k4rJCZkyFrtdYC8B8WmiEfNrogr6kYPJteeYXH48r9BZ9MM82vu3n/
LDBwRqoM7W2j2gV30f1tr3Uo/FalcvtZURoqhoUczl5bGdCC3E47cuB37PF+y+z9
DUSAZsNqQVvjncEfzZeoIhmHHpij6Pjyoy6v42R+vN+U7571eHqcQIqhyBBBzMYb
P35PZRRGA5+pjM8g7RRw+0C4ZKgSbKQhUv5cyvQ8gl0YtHn9GB+GoJDp6GaZOch5
xSX1v2ho5xfbhO2m0B6l0ZsEfatv9FVKRfN2A4bpd528FqDm5GfFIRe4ox/bNwzD
APGFDP3+g1HBIR2PvO+Y2OFNa2yRKEQNLUixF3p42lNfDkKJ9WaVtCnWYn5D6TeX
NN4B3X03fMqdaVzg3HDpFtcU42rHMXKyBrdFUozCff4lOMNWCAHSFKVVO/mzcN2+
uXd0tpEwuEBkZRAkgEHM5fNd6f27BeJ91yXCmAkbRkQXeNPws9vKHvulvNsXY5mX
LJma9CLB24micCO0PxCtcVsk4WaGs/5WkPQl6ca32bp1xZH9QWQWtXhb+2hrkh0Z
v79XVDy83v6eRV7+OLPK0hkppFp1cdQ8Pr+3iR7+zRqTZEbLX3yHgrZRDex7K4/4
LRrn7K4F6i2J1vvxQMYz7iTdQh9r0nENH0d0p2ih/jOFSXO5Fk3x+wvc2o5C+Z21
ECoPwvt3MGB5hQ1SDuV8MOA8Yh4UECCJPY9J26X7A9++SgyOkq4m6ZHIaf3Crt3v
qOyr6nXkKK8HD1+fJjynzx/idePQG3NO0T3bb9tl8Zg7Ef66PBwB+7PbqEoJqjBP
pOF/xefeArjxOXqegJ3JorI3IzNCil/yRb8OFZvGg9C0B141nJ4H7BdyoFhh/oqQ
h6FoXQRk2vqk4mfc33XWhuXap9LIdAGiOUTh9QubZDnKwjta9HNCjDikDz/wKj8J
mb0OUM8MebScmjqri1z3P/j1J+N6qXURAibPjUNVC4DXtQMrjK5VdP5+Hxnrnjl5
hpoPAjsTTmpSrueVvr/oC3cZsgcBKcbiC1nLfNt8xiiaC/xfYmotfG+6wvq7Hj/P
w8XGQeT84l8cAubpPU1EUPq5aRh0vddfCuXlKxapdKmpiI1JIEfGwt82l69N1uE9
zT6N/BdnSW2t00TG2LaJbeE2BWnq0NLEtmUMovu4ITTpLwR1WpXGB/OLq1uXW/gM
0JQVaqMrIwDppED/aYJIqgfEOhyi1BHMku3PMCJIp5UtmApCf1aIWuryuZDLV/ch
gbaZV0zUWsKLkHroz3vRv2TgKJykjpIXT0Fvpf5KobVn+tgQXvU90tNXRuwYVr7I
WfazPwPZeHrXKSb3VpsPTeLydOpHt9MXxC9L17Few44e64wx6jowcbK+36iXCsW2
gBpcTslpaT5cR9xDy+BjA5HFGrXVW+6QP3RzapUZKyMPJyKueJztr+iQXNTvKjsE
vrlH9StbCz2IlQTPby+CQHPq7hS99okvlu0Uez0rBz2ht69AOzUEZ1Lnx2VWWlRW
gq1q4GbSxxXsZB2bVq3j1cfav9RpxBj3wSctqCid+AK6j4g6FhXZx+crEumn2k1y
aSUdtG+D7zjCQ/xQBhC0m+6FzWwEk7clZ2xA6CFsz8mkH0KcDbM+cM+qByewDLCz
lrRiYILiAcFoojvYJ1nvRiPgUbb/BgrQS5bmN5dZNMl4Nh3vKOF9Tjn2aIv1Y6V1
obLvtf6kPzUxmOom5WIReT6Maf8lPdTVd6ziHz9TCEVOhZeQqvj7xJkAE57A+MQX
rwm8qnRN24KcuZaobj9MxxC+lelZ4+S3KCv2Vj348txhYelmfM22IjTBbVmQmOhp
Nq3Z+UcfCKVQznHWyWV05bRBulbTuGnYic7nUGnvpeqV1bsbjyLMzS+nkpB4o+k+
6E+1flaZyuNWRxz9uXuQ8KD2VPIS7iRV+jyYnIvOO5wEsQqhrB54Z3aj27WPfUHU
9MEHpyRQJw+UpwMke0iPC85CxLn+yC4OtowyRMIK3o00st64jCFEaGeba1n6eErP
/TWHjqTobG/O7819ce66ROAeOY9uDoQzgDNatvQ1RvbGrepD97ucC+X5Ntw/9xio
r5Tjxy6lmij/YCEx57Dbh3vZv2qvTx+iX8Egxt2/p/97EZ43BOWWTFd+Qg6EX0JC
d7Yhfp72TDulNxs2U0zR6k3KwbDOsx0/pJGAMHIl5drjpd5SCyUQADIhH+0Q3IQ2
Uj17Ngut50EhpQtYaRB/Fld6mlJuuD6AAyuZQ+nOrrHt/8Zmy2Ur0pFVP2R4zim4
5GhQygYLDWuBJXhjfg4i/BGAXxplR1Qk2Aja1ms6dybGXMWmD3iUNGSgi9pd7Yyx
haPIrkEoy67EQVNITPEv7eFl6MDYdxVG8+QxCx9V9y/IFzuN+0X13XJGlS597oSW
Ge85Kl//U+tvh8egPXQ/HkVGE7Rzt5F45I+4xyfI6FZfS2iaq6VznxTXn81lZRBl
LVdbW4N/Eh+1in8cRaGI2JCJc7wWlvxvfshUJvxBI8B6hNYgUSQYncWYoJoZseck
244HJw2Yx0sQIvRMebNOLogeOvByry9g4Qq+LdvY/NLqu1LfmRaYvBvc2S7VBQbf
E4cMdFE1FcZDcNMxWlefcje0NmR7AMXdnxngkEeiKU1Gf4QdcHCUiGESf16EwNfY
o6e3LiRj05e1qK2p1L5Vg7+Nn24F6WkerQpBPDxEW2Bh5Fsn1Azgxq+Gp/DMrnC6
0AAS4Y3FINeWirh9pvI9TGBE9Ln0DPrA3icJup2IwMmRPAC2xPHmkamV0Yh1AObA
CpjUSWNwDxkdFajSCOM3mLqf1ZWb5reIsUd60tQOaTFSdjkwH9t0Et7dw5EFSWMB
e3m9P3wOJZZAC8aZi4cEVcJ8kYZpUygjMh6Rg2HLi7FHmNTrZ43xeLA83ddDEhAf
XEJ8fJbmTMGDFnFTbT50ymUl3ccMl4hYogBkUuFaD+3GpMw9b2e5Q21h5KaAKFue
05ZA1CrVvDE0qiZES2bF01WpREOfbMSgT7ryx7pheklksKbjxxyWkkEoHx+ene8a
ankis6QzqTpgCu3wiIhwQO04bFUroce9KDgtMp5JGcwjWGlqWroKR/GQ4SzxkQ0l
p8cwBQHlCGiKa7FimaPRw2Wnk3EGkyjWAxQq/XXAdp4eHBn773kOBbU+tRphr8xn
rixvhn5JqthY/cJXidWmMY10JDvfsUcDS5sfTyu8rcXKV5GVQtjCqOXnxtjoBCUo
HmTqBp717XqIbkZZRo75eJcO8KLuQezcePUTolZ5P8eu/PCbVPaOsI7y6tsrvDOE
zlpFKCaBS4gsBdITVlqvNrOU0QtAiwgSQOqQilhV8jrSCWMvOJcLAW2xZnVA+1P6
Ug6xYQuw9Spn3v2lWvbs/OW/YdXIzvucxZURMat0LXKAHY214qmW2LuwBt/LEsfk
4hI3o9bHuBVxAk03TbEm5pudZHdWy1rfXAnzzgVMCFgwOTiJvY+LNPWzbM3y5ua4
jq5gE9u17K025anJ2xvPQkWoFkuE80PzaNEgD3lt3cLcUL22cagLJ/+bHWgHVPhM
oj8O8sv95viqD5+o83r12z9O4bMmKaiKzMmPXYuqMYgMoTTvwZOS3yHxJdEXoXL5
IGjF5mi3pxlzc6ipE1qPHdHXJla/F37xqIyTm71sHVxWp0PoVwdTHIuddt2hB3li
8amFE7hgrM7M0lXcStkOlxYiWFiK1lEKxtGbg9gsqNmvHdzKu+imR+qRkJuI2yzD
JgcajIWMU/ebi2VYIixbW8J25y9QvTX17wETCTh5N3XA3HLufjPSx2+AdJu2xD9b
OKYT3ZJS04Y2rBRgSplNP1q0z7YkfB7JJwqaI00GHgAmDPQkg0ovvAdLCNs5cVaO
6/hSYOxSFWfmuz903kcUBqBAqeSnmWGwXCYP9R7fXbd9Pl9FeEB3G/nJWQbsMg/0
qtDHrPx+RagLTBKGkuKbHASX3jq2sNdDL2eKGBfOaAGemZgSqFUwFvhbeQ1t6ZVT
Ql1SOsgW9YfK6bnFu/nSTvpt+bKo1FY+gwbsoyjleikG0xgsBMRUHksFyOjW2D98
I9HRmmA52dE5dcXmCjWZNSSUL3qVa5TyWrAVNBy5p1v9fMb5zWMquMuXkvi9QLmn
rfvLqamxaSisGAwhPxc0uHPpTghLcZnKphCFP4s9aLDxufcyvV9/ymJ46JNuqfmw
lg07YTUEHuDFxv3Jvdtllv4wImwuLZSMRcctzSErRVIiXcZRIDPlFm30fc4Ngr2P
2Mxh3Z2rsWWG8NoFt915xPw7CaW7gmmsg/b7/4VSmdQJVQldJzUQ+PV5x8lEaJbe
y/vEOSH17Lf9WAu5nBbkfEc8/Mz0whZsGRpiXvv/haUYXdt2IGksDZPO7SFbtTEa
A4XGusNtHcGWo5ryXSUoNXmx/hhsW8idf0mW26fWSP0BS2IobMyqY4DxtexyVOq3
ft0hn1M9hk8/Za0k18kUKvciHM4PZdowlQxct4gRadWIQpkd+wsZqTDbYNenos11
/0nVycxjCAYww9cgJdw+4trUYeOnpRw8TC+1aAF6x+f3KvYRqCKItZrWYI8JYL2F
F1j40KxP/sUAjenR6DzhMI2xeWu3F+TF85EtDPyH/AQAqIkbJ2n9skEBdWHCoRc1
zcr80G8bARvdldVTSwQoKJQyQoedWGGNvvxVjOtkCUtVjBMuFu4T5KlqaDUDlFDh
Bj7uGjpWHoBJr5f1bnGJM8pu8pZxkqvptqpuWJAxihGThOo3mg8C+4du+JcLFN8n
hxJ7206oJP7itEegmnTAy0gQQMo9MkT7etSifPLaN7t9NO0M1eUlr8Mg4zA5tgp1
8hM6XGkh0bxpsARLUoo2yJG4qJxG6z8adEQvZrmCV6cso60aZVMImj/T1/Vwdptq
kOTloxJCBkRFkFqWow9mFXOIKBDimak3TIWHsfmkqbXjLE9YL2hKN4tVP0c5uZrm
EnaJkNHVTq8K6bmp9S487xzlpme4tfp1sU+dqsqPwUgDVpdQ9Cl8CNnu1SLEBEDa
5alxyJt1dPDpmfSVJ2/RAttLTSDis0G1CLQmHm5vvgeVU1TPYQxYVo1z3h9cq5ZW
Psj2MvWrW7Bv757gHzXPO6Id/erq3x4Fkf5mOtUs0yE3MB1YeZQikVGiUzAsjIAD
/lTTP9jschRHyNESlB5UK0THB3Tqa1NLW+zFCm9/j99rlekL7NWxoBqocqKAEuK+
63OWWN4D8lvMsYj2mDOaSnsL4GwMwCcdR6bSjYji9EidKIExKvo5VuUzwcF4qXPI
CwdzAsIlJMW4N7jyZ5Z7nGCuqVjQ6bP8o7yf19hu0mko0A597Bu5mKqdrMNgJBoq
ET+akeTI5WYYV05xKPKVWLZoXj3K4HW/iBS50cK5kbcOWv5vbhXi6ev0jQ+Y9krV
FCHNAz/IxII0F3prTsW1q43gVBBgimAEQiZyZFguOhZhc32WqV1Faq21h6ui2lyi
HryDRi4mSUgQ0b+itprUCud5HWwQH3JxYMVLP2/tpqpDPV6aNIGGHLB7f8c68ZWT
ZRh+0lpK5QMX4jDCLGLQBaKanNYjQYb30ldz7K7JY87bzylHUqYbFdv+2Y5GUj9M
6uG/sXyFyrKYoHix81y/67ksR0eyPGYPVnQwVEGO3cjnetpnjCaqP0h80jj/UgK/
z1NhSb1niyqyt5yxMxc+ppggXQ/I8UXkV3PbTHoEKEUNd+agRAZ8lLTDGqg6nOYt
UPtjbgiHz4EwevHJj0AP5b0OTJUAuLgzPqntoOEHOcwRJXvO9P4iau4IX4lQEes3
COun5ccBVzBpi4YYsSA0udJAv7N1fnjdJIoukSlKmj/qSj8eqkSzGfy62Sp5IVMB
/8TBh5tjXX2DDBhS9rFtuVEUFxHCT97Y0SQIJPibIIRdDj3QVqm6LeZSg8xphiId
q0ZNZpmoQ8ldcSWVhxwurF2dy0tzuGZ505KbHjc6AAVVTI3dtDekk3NI5GMWIcmN
Izf9Sqes2CYrLnUKtd0fQr7TeV35c+KXt5Bp8Jdvc9x6xopHavblf2EXXuVxsHAn
Oel6YUdDhKwuCEudfGnbVwYeCdlIlVqmeMeTQXz/djCBGjkJvqtbH6YyO7kautQ/
jLm9TIA/zTLi6Q/bcQYXtcgk0OPzTpludtKpd3WxDT297ogsAoNu8+j8Fzn/FY5G
inBT0rKykD7T+2UdjBGAdqEzYnWhvfzMNgWhpdUmycYj5N9cWMsDFmLkgcBpnaN5
QEUKZbpbACozTzrJkoBVJOqV79N2dV0L7+jKdE004R+locri1mkq5PHK+mIHxoWD
j+s6Eg5S0xiWfTNd0UrbWR9mIhSEerUbD0twMhYTEr60xzSa9gfBmG3bPVrP1KFW
VcAaL+wjHu6W2Ik7Xn6qrs4BOVe6DCFHquQ9HsjU9iA8eyDPD8YYoYtla13nhXCr
lgvtR5qyNG/Qf2WeABAlv2i5tWaDr/oE40k9GEl2NHvrL0IpMNoU4O3+waRYDxN9
z5pPRjghf49MNNtYLHBrhCz6hLpeuITnDrClKm/BDMyQgIZ3OgvCP4f2/8u7pYJy
ZUiuyJWPDkwGziPivkizPB0vo9qtrgjLBRleuk+xPbX3nsdUQKENAG3dGAOWqX+d
i4nbF6S5eCqkE1Ev9u/hCKZwVhUfqUQrNKpaUAJ6wxSEJ9luiOmhBuqlzoXJDFWj
xDc7L/rGEmHdLxW8Rl+ePhB4P96jw6O6+ubB1Y01eU8CwbwCd8wX2t7ucniHhpzw
6rVXaGycFb4RnyDZGCus3/OJLiB3d6pP0LM6JCDpP4kU3AX4Q4ecL3kvF6nepK+4
91qlyS6Sk9FwlTwHjbFJgxHDvGaLB3v+1oevT2VqnoQ0W7UBm2v9mLe3DCwNJ4i8
mV2klqv6MpyWIUscqadW8yF4k79NRE2K84gfN+4+2x76vm31DHtsIhsIzu4PDAaj
hwzEXGOs4hbQPXOaSdo/cMHh5OYo19zN6uwsCvgsIBsffAiWizBBkV2OLEiA3oPi
Z2zXgW5FMW2afWf2atB64bgmq+bX28EKSVUPz4IXS3m83lLEuBcWjBrBOO9rIUby
wcRbXSqWdib/t+NnrCR5OHSx3El0eSdhkClETWfH/U2vAMa4V3a5y7PiUw+O00K5
3UgxI4LZa7HCejyQIiP3ADUdZiRayR4+hqR55eovs5C3h0w8rVTcTLCCWfsuwP7Y
cg4m0L9gWxinTGRPT/m7vKXRYPbvckhFnG2zrkVlGgXao+vcjLR4cpwozDcolXqf
Igx30KaKjhIRcArZJxrFBOdQ2aZssGWPm9wTsLAfwX6MJjmCmcyBsT9faoUx81BG
WVlM8oGoy1+SotdQwoDdL1x8nQ69l+LVVhuAbkJR5krVxW07bAH+4C/z+cjrGZNZ
F4AcNqxEzyY9DACUABR/BJ2Tcw03q0eSUiQHBtznqTn04zvpChubH2qvu3UodRRi
n4I5W7BfzWzIOKkXJOs+UQ5EHRFGV7vqzLVFb3cP9ZC3ByNE9oFn12cARyE/0ifN
cVPxDQSKteojo97tMdMnVffo2RGQQ3yr7D8MJwcLRXsvSAkqBgX1OHMvrVD8bi6A
aSWlaLBMPJRP1rqqo071uZCeJV6KnRLqg2xwAUhfbeNdcKIrHSDM/XB8U4WGFLP7
0oxNr6MzWCa13P7CRA3hgjM2dk6OvHsAzhEgtPrX+EcMt7d7QcfbtefmdtoH3Ofx
rTUkx155JKXY6qmVnUg1VD67bQd8SEv33MIzD29fNGTE4EhJwMnrDEG/xc0u6u5E
EH0t6s7UbmcwCoBQ9DX6tL2L+oiGbc+wwWN3JmyNO7QzokrjuNb2ayBTGCFfqz7a
1Neo0B6P18OdkzLHv493VLLHA8cFMIe9LWJpFG/odC/YAVgledAgp8K6U2aOq83P
htR40tQlExn09I7HpCFGh2ZYozcQa1wpjpER0YFr4FA6vMe+Qq2W1kwCR/0O/y2d
F3u3kRTeXPIiHVXUydYSXpYgc7Y4Bb0xjW1HJOyaN+mubye+o1607OD9gDaam/MD
58MCdoMZ0eVGCqF0vB3Qhj0NHqztdia/e0Lb5xq9C5lxdA5BgZrtmicjEAT8jY14
Li7JH0hUkTHc3fLa58p37QyMYcbp2zGYuJoFEou91lN1XRKGzE/30mMlW7a0Fc/K
0IM0cMjKnj5C8WRu5A4nws0r2WNmwo5ajj76LnYqG7IYcbW0fpEhSxFW2Qh1Iyv9
dUgi2gGoB70eT0T3b73BjojBWtrXXa7y18SKDUWohgHj5YSWA9LYRIizrnCc1ZCP
1PmX2IVrVh0vmzYL5NANkdbAK/pusHdmCD8gocg6eVgfLfzGMxvNfpuFnTqX1Jf6
ejn8r4nzN4aad+pWGJU/bNBnixIoXMJuDgVm4qlAFQoso9JYootR6egPa4PIh/d5
B2AYG+ufFhbhGHkaoIdjq/CRxOzaW3BshxVQzLrSAxR+5vbOD0RzegGDLx0ulYrQ
NOonI+2cswyyktcWdwXS53SH6lS1vQrh7SBCVEw9+PlsQ1WOG94SjJ0ZwLVLpURd
5A0oWa59q9gfmDe9XeNTRuYCtzEi73wfdRx79KN/6PaLE0/3SHAy4gU0eeqx3Ayf
7sR3e9fsbSjM1ABb0rGJRmyRzLFnaXJ5Ji1mGKN3J57GIsJIQifx9V5wFgsAYh1l
e0wl0Gv4pGW8XvgB8wTouuekaArdBdEEZ9J3Suzom9r4/irJRI0PC1kwZh3FKjTu
gsCfwEDvUsb+bQ8GYFPdFL9HjP8heGKB1JlLewrYoZAVjTADTItqoOq5TyO/7NBg
TUOBNQ7H4V4yj+6x9S/ZLt1E/na66Gmx8Bj++oYcVSZ9ikHH0+CsO/LadE8l6xAZ
8PL4/qN4bM6JAXKKWxt1c/O/VPXF/wvp0m1ur6sx8Cf3Zun+pxiff1H4nXWuVS6O
4eqaJGH5Llbgivt2KKjdvnVZr6OPuQVUvBPdAD4Nwl7xklcdn79JQKmjmkK486+s
Cisc+nATCSYyrbCQxxPiGt5CU7ts1LkefIzOPC+NpNAt2+Jjek96iqRyDjDHWj/N
OdtQ7R94SxrMRWUq/5t6eFpvN4B2k2K6Bj14Sf/QSAKWOiJu5WFfgDS3Xynz1vKo
TYkBJHXvBkURwlcWJEBV5PzU0Lc85Zaaxyc6coxKHPFBzWZhb5xDdg//c8+c4+X6
aRUJEqduREfIebigarE7HZ9eyyCC2R9gz9MjFDQKdATjgfStke1Ozk/5u1Ft+tr3
mPLNqcDOFWsrnizdxCLyvq9WeuXrVG++2Wiy1ysGxcYxCoBa7x+BncVV6ouWsRH8
iU+J+Ap3K82AR/AGv1tnx1LZlIwotCxoxaUHQK1SsnYjJGv73tVOGfNDrdVMcZ+g
L42QfvCqKyKTVwmEz7Maj4ntwNLQBkSFKjEF0LQbZCoc45r7Sb0h+zEDhko60i4l
//BYJt2GZPAdfdarYAMdIo+yXuBhyErUbVJZeOU0OfL0F/0VhQ5gEUEsLcx8/aus
x2MUr0HsPWPXG7VcSE1AQtJKUe68eZ5dudGVyxNp+UwQttpKdE1e590vG9KFomYr
ZH9l7OEwqro2p9LYZMSaB2vhkT7jmyjhAdTxyor44CAfOSsmbEimYQkYk8iOA/a1
J5CUlfhckjLJnRYmuxbvsSSdkmWkb+ZA4edhJTvg6SLMQoO6c6joNM+eghC4bL3U
LMHsSFsmFzI7F8JYnmrNWAXhdOnRh6ZVx0gAGUBv/fRJCTLbNk6NefXuShvgCOgb
WW8CrqnskqmC6u5n10+qLIS1sEns5YTGHZkjsYnhRhzwt7MTwQW7qZnLa2UKu11t
ti1P+eMpmtxbd5lsJYSIz3drOggUMT/7zym4SqfEZu+nGWC3A79tvFODcKr7e0aw
92/y8zL96vFvD26btAcHVlAlGjjQciqPrkPRZF9M0/6OR3/v/lo1VOUbWBJf6E5Z
5zQv0+HnbzFmsOMQ9U/+BTUW17jhVUqhK+lYJyHBl7uKQim32h8VMmNfV3/U6GOv
wnQMyHQJ7mzJU7bgrVA1PTLkDXgvDW6AadDvhct8UHGlCV6UqNf2HAcB7PN8XdYR
khWFagt7Cq7phUdqOQfp03+BkL4UcDzlxnAxIrz+Csr8/OUY48SsQn2NeIC9bGOc
GpJsHvEgp+0pZ1ZRrgZOnKsiCDv5HPYd14h1vQnjrLJC8khWRR9b9XE5kAEcVv9B
L6gIGVfdNv6OQ5Ra5F77X1ma5dNZiQ0e+A1zU8WQ7gMW6UDbzSStYVgaJhm92Tlt
ZzcXS40WM4ukaco8LQE8TAXmG2aDe+Z7SbOgoSMXiOTaIX9VaTbJeJvUvkBU+fgN
l77SMBovJAIqJeixykrO1FYN4I21CUcQ3rpUnQABESu2gs4ivWxU9coYpUmbG+ST
Ks6CYUHHbbZG9eiaYmsqNwBQXnkmtjpHavdeDbJljVo83xZd23rpgN+9aPS3uihF
wbeTaw+RAQhO8PytlC/I0gqi4hy8Qc7ETTRuyINH0gjhDauy74eDr+XFHxUNxicW
gQoVQRoS2sKaXzhs6DSugWElb3owbMOpRnnd1yWHrYTgNBWFFRnkjgeJD6R0FVI4
AMLExJRuW6RY3Mse5k9IIbp8i3OWHUNAJ9rrpXnrIMX/gYSx5nALFg5LFVzv9e/0
eGQ5T72SyBsj7f3FLfO9M7E1wTdDGVL4FYpgaNxQTNWQ7qE5ZrQ/2vLuN5iKZzS0
/6eGCFk9Mgz5T7QxR9roSvrarZnUyhTDxnKjjz8yLAcRksx2iBGoGuVZB8L1dI8P
TZT5KJk5NnJwNyC8vIVF3LTmngnQvicMdtl1TNurz/mni/dtgVkcMO/6+WV6kDRl
fssqLiHoius22H7y2BfieOKIJ8anJ4nYhmsDIau0RkLYxtIwVw0pvcZQoN2IMj3y
gFpvD1AMSCGbcZVWVMgr/KYNGw4dUz7+/xe4oXzEAECURUv3+yPUZqCV2ZNijlT9
im9GDmDfyrVOTfkfvR1xg3rIHFLrzc7IFTyn7YtwZZitwrPKk8pE3PwvQHCIUNxJ
eVSgjAyFwlN+yWqE3ScNAyY06dXsW/KxiiCcgLMrlxqIIzGaLkuzvo2tWnmRMslW
dwYZ0A/ysI0ahfpA2+VEpEk3ijUPAqb6EEpOwS0wdeX/4OJFzIlFmlbXAGr0onRI
yyc9aSScqR6WzLWA7t3Kavllj8Nl3yfVqF2Oi6JnpjaIbpdr01tkVH+MgqHeoJJM
PFn2ELvmtzwC7VQbqAu5dKPf+gpQQhUyJfjQ76Id61G6ip/ZXGpnw3Jui7tkU7ca
KYWO5/2+aE7j5ewr8a41PxQGpAFs75k7OesyiMyZao9tKnRJFzKX0yJFdygklMXl
A0bB9n7E+Gjzoi89Orc5FdbZsc4Pun97D0R+aaPpOZhICxNn0ZvVfy3HEsR+8q3+
r4ZjHdyGAeVzsArttmrq8/+K++Mrz/5Sk8WMb9TiBrXQqaV1I1ZP6LH3ie5tGaml
lhcMs4CuiTw6Vs/6bHz59SflHWnDWCFmY1DIbggL3l7o5Ho6fQRYZYWss5gN2OXj
bisKjy9QmAg/mXdmbOn0tvkgg3/7L/tt44t7PvAZ1WcixyLSQ4He6OVvMO93u3sx
MO5yHllEkXibNGI6jABTHPwztxP3MUxeN2OeYLasSoYvBBzEHw3JcqUbtlhUHry0
F64UWaAtOda7/DsNAIs+hZtz0PXfoYVoxasAuLbqlYbMMd3AH1r7kPwg605l/IIJ
ZtgAyGxtFBgrNb7Ex3vLRPmAi1hhP1Vlg6rWUt3+3E3a4bTNuBSJbjYRv2/ASEpM
TnRDfihcIeXQyy+osIFn2l/ufs8zaG/iiOjT7/Y7DII6rbnNfrgw4QrgF3qV2DXe
XLWr0DEoeiYfOgBpXYbFx7rYkj+Wzc461hWrLzap+dOzAQMRPo5X496Qxu2XpK6D
gwaCLuhvDpP4goB017MHeC8edKlGy0ni0CsdKb7cVWN/V0/9xNf+1uU7wfEs8Uco
cvBLApCaR3t1/NieGRY4OlbQ47Dj9zDOd4tgKSfaE+uQbZfuiW/wTeCCSeUBTGS5
TozudHe8P0YHm8Ka1MexqVcJImOboO+2a05vvKNTwZWZxQyKjxK6EVNpVto06dmT
x8ULc0h887wNAiiJYYV9cLuXGvzsS8U7aOi4TqVUPClVdMrajwjKXBu3Dt/Bmg8Z
uAzKHF7NbCltq0HkHwPVLZ+H/jHGNHCbnOXbvEOWIOWKMwszN1a8+kSJMG0SCJGV
OtjAGqnuh214q7hWdWkymKK1prKu4nqgOI1nIhISd+XF6eKxg0/42gKMHKjiWzQD
8xu7qrWsGvhjUyBO2VKWuoZTGcHr8/7Tzz1bn0jQ0yjNGrNd/yy3agFMwbF1CcxI
peR8iph25No3bshUaA2yMAvIYF4Wx+0hRVQICvTF/7UOpaYWTZn04Is+9paHp4jB
91MkShgCsdD5k3LBcJIc6BTxJ+9jIAHzsiadxk6bK3YxgFru+Cx/ICaLw9JraXiz
GvDwedY9rFvlDGQxHFDbRfh65eIeSP+uyIhcbZM/T/Dy0IvzK72UaE03xd+NhNCX
L4ckbgw+UQ+sayEb1OzuWV5/OiJXGC89duJp0mFOLqaBjO562NlBiw/28OFjUu/T
ekFq36Kp9w9vI6wWXDfoH5R7bYQM/EPKTdSuwpnbm7GV4+a2GOfXiBFnlxa/Ugzq
3/S3avv6VEItlZJHz77w7sClXCAUWaFrKpMfzDRa6sXTHGudHfaTJYZXmbZfSvuN
1T5qFz7U90Zzf57Ua663K6Nv3xZgeFaebh6Fb08Du4lTo15n6esBDET/1kY1BnxK
7+DMNzX+SaUHC7PwuQaTegoYt740R/tjq7y5G/V78FMFl3zKBstPadpxhKsXRquo
zKxdATmuz3ePnE8kDGUFvzp35zQUX0iHKgAQM7z3F9GONaZqITycYsX2xjtBuUqH
WiQZkOHxNa72lipm/TGhM6REGuue8lPQ2YTie/PnT2kah3hUtk4xk6W5kqMNAd+l
nltaLDjqE0/Q63FWEHT96BszRctUePtpBoaaVb4gWeNO2Jpu112+0jPdXWDQcKGv
srOEB9wti6qtoZrT8Lu/mJ7mNEnIlclNn2Ukfof9qmhd3xKy3mqQ0M21oGnIPCmx
04RN+Wxfe3wQfjrDror7Cb5KW2CXifEkOtP8yuv5z7C4kI/BbO3xYhwBm4tQr6BV
Z454aKzbyrRFXmYq+tfpD5xc/IhyQlscTlkLIIueI2BrOaWJiikupZcO6fPIVb2E
dmHtYwVZk5vbv7g3ztOBk68wQodIkDuv9Iu6RWRx8zY0X9Z1cxD07ntxZE2ceQ74
QFdaUzSEPAmzc6dZS/qev57j3feX2la2yqGYg9lXbI0nlJEks1IF1QXW/IzGNvtg
E6ZhqaUCmLYnUZND3eb3I4IiVSuW3pYBFVjG3vi5tylO+2c28zaafmHv/djolmm6
TJgkFesbbQJf0NCw8vgq84U5zBYXuJf/98wr0gewx7RZwFqJzOPZNJjht/Mu+kAN
vAh9DO3dghwGqnYp8me/JeGQrCD3x5m6kY/a3NVV5b15s3AVtt/537h65WTmk76h
QttnwK43VzIcFYb+0fdTsO39qykMpGKovgzF3ySXLTkYdE1Nb828DKfbA6oS1fiy
A93iaWw6KsJj8iTzVegp6PavzOJgUXGREBj705/c8ZND81Arzlh5bfQ5/7ijXl4/
fxIfx6D8dxdICpF+x6HAGQcl5uqdAcQiQNcifmsR4zJSuAxlVY26Xpy3Uln9ZCz6
pDsYrp9xSK8cJLF4glfFQ1uaUS7dFCEssB6D+OXBSUv2mjqzpT35QDctAbgvA2e2
d7Ti5N1lZa9FO9Cjtcsl+HBNtBYN36lYMG7zYBj6HhEGbuUQ/QDVDaYWsycm5MVe
FVhvSIBbV6eVpcu0jNIARtFS8RKTEQJTQt+Psts617g9n2JN51Z6bcHMtcJIzeky
XZ3FUcChv3c5BS95NIMj7N7n4Kz0aNNJBgBsdHpsiOMKlAMB8NWeJaJYMXqIJ1IG
Q/WMQJLqC1eVYXKMbmyZ9FQIheQONdsf1tdHhGcAB2F4FaA2oxZHZGeGpP+aFvXo
dMffgdJySpXAfIuuTL3cLIEiwlJQATcTDj33wrKAsW0ufvQ68plb3bNs/wlvJfYu
/ADICQOv32h/P125ydDPzWQdOCLc6IRrv4GPW9sN05+w/DVIlfejMkpU8Lk0fVI/
VK7xYQ3PdfKdRsWu/1/oZgmJ42k7qsKdL3juywHQrsAscy5+4lu4ieGFtZT/bbTT
AzgNvNhsm/6Qes0/qD08i8Ik8lxTcNAQKSL8P692dTEbBBzJYTeIALGkzHUFG7sK
QkpUilUk3j1+3uh4/gEvMcTJqCL+UUdBuEX8kR2Eregj7GECa6nUqlZ24SO+kLo2
exjlQv3ZfZ00cZp42TMssrcihISL08guUgjNGS2Q5Z+IbnnmbJl4f93F8BIaS2su
YYZcMNbouX9ymlRCtB16v1TZeE5fyEup/7S+5HEIipR6xNyZIRq185uYl6oMBGx6
/PE8mrW+dztGNkjirfpybEwx4mYXGPgYtUJ58mYyRThqCyx/5UybCYU9Zxzwd3sM
I0IvpfNV/HyR14Cu7cTZu5Vla9TcYO6fMWEEHRdZ5qiVUdKkwM0US+S2o4uRQg5D
PgWFY1zbzjePIS1+6Hyk49esmV9a8sQJ8093rLs8Vh6EguGSH427kONnf6HogRQR
UZmrmUHda+S13REQlK95z8ZMHh8R9ggg8AgNtnud676HJ57D1Bd7369ct9ImqIEW
YBoWt/XL31uRW7y6taxian5yc0DwL0y3ZbbpZ3Hike3YRm9/xFXXYE9S9yGXEW0v
/IsY7Zjxl85bCMiYNfRYZbS/Gh20qI0zMNJkH8vgOI8k2uu9i8QJeLT8gZ/cKODo
g3fmkPybfUj18BjWZwRrJHu0Uf3Wt56CoDueKxbZ1NyhX5Q4G18u/+BQTDPecBe9
oxYBjEy80Ws3bZR09rOv6NNi1pdxrrLsOTxAtcjPUUL4zG6411dj9J4AFFd+dQ7n
u7E6u0J8nmv0yXbU4LfzIyWdmBJUobzS7tDZJ2Uh6e956FgTbaBcoPM36DMQWvdt
3E3esecCs+Lq62YYuHb7dvBl9aRKpF0wfsd0VuewEKYcCJcaAa3jg33dowxbX7IP
0+lLE3otgph/EpSNQ5gsNqXiLl9CbnX8XLZshtpfMCUDSbBSsQoSiekZy9ja3O6Q
JWRJ9BOCO0pmPnpzhvJLpLQDUTacPgHxKrrWOymatajyOiT+FnaO0LUlcjrCaX/e
GlrfzWKC1j+SPr0srq822NhjcOZQRFrwMhrHCpBF7gdgH25yAm6G0RT+j7kOJqBK
hcugQXm4IAJOf7DGvUYI+p8J1Bq3KFpS25kcW/6+kDKkdhV6k9IaG5/6AHkyDdmW
AdEhfXSaxg+EmrfnFIgiRXDdefKEWe3cOk4Acy5qtlbnETwQZphOyaUa/ZNZvW5b
MUeM8+1jsH3dOUebbqxGibbnAtyz2vx7AtvonCfHx2Ca3yp8rOqWgBZpMqnYMAZY
G5KKe02xOvg0GPXYD8wjklvk9p2JIN59Qyzy10ah3L9zcKwMHE9xbrEiyaWtzC10
zdX4geOv3ikVcqPpug0kKnSlWvZMSMVxcGxUxIloJydYrfHEmbKcis8ssnHVfCES
up6P0zXQWON7oITCH34vA7Xr/WxuntYsF4iNDQYehif3RjH63dbpk4cnR4d6fPTh
d5gwIuZuSTWCKtHp/lWTXXKgbZNvN4E9WVHLAw8cHWHgXA+cEZDZUpARydJdZlL5
F/AZAXOmHIuowHybLzNkyhS+iFt9LCE+6HaphYSJQDfZTvWcJHnOeYgkRFDtn+5P
RULCQYvhOba48/BB3sDahIQw5lPT8ATBiQ05gflgD53T6h0+iJmIcsNcuuPzOkbZ
90SHgSWDCj6ssSas9xIinXcWDSEgAU4IF+pWAJFlm/cbFyIR2VR1vqkN+n2hDAwJ
b4sIFDYv2U7JI5uiC9Sr/BnR0j/j4jXKdkQj2QeUwCffwNJi6/ZucZH3sGeNLoiS
xT28RU4QkhB0n+kKwBOepRD02eyr/So6f3FMQliSA3oYqva70bBpTxrQ+Op04f9Q
Ez77uOGixMXLO+CyN037cMmbvlBAvvWV+KmfIocD469DuBvG1ZAYwA2JTcB/CqKC
ObNGWRG1ALVm4Hhbks2MM89svWLaXUc6kTStRkOmMlKExRO1kWcZSbqIucEFyRn0
HKzpi75T8xtSjDL+uYHnKeIK80ks02Xr1w8yXFhF5x821MEBmgzZcXR3TX2iEYj8
fwhVSks0Hk5ubhds1sAdo+Mr5du0XHehykhsfeFi8P+CesnqdQIWxRRZhIYBqjuc
z5xoSHJpW+xosE2ChXTU7su2mhRT4g4KpSGr3qENGwQZX90lr+RPmpoJXliN0N9s
8X15bWylMxslfPlsuwJ6WUyDx3TusvsfsDyNqWutdBPWltnG8Mpww5VkNasSt2/F
fYw7j89dbpzEYQ20zAxFm8pTB1YSPalfVzFICQoWZYY+vXCFzlvl35PZAd1OfiPF
j9JPI7iSp9C7CNANRkIPfi8SiElrkqI7pSLhadnYAqywIChCr6hIVgFRaZwqPzRB
iVrcLjFIOEikYbMYC1iWHa86TUv/tJto29+DBZEDgk54519zbxAi6XklU/hM0DMG
wM38NGhURGN8k+5HF5ynbBkmMx6coyjEEUYuJoOGoKMfiyh4b5B6guXgjTJmhlKx
5WCEv8gcL2zDiIxwpwOd9wl3tB9XZ0yN6q7eYo5tOgAbYrd/hG34+z76Pg6sTwSy
9THKtObD1bTcu7ywsGQwAAdSy5/bii8hRnL9e3UXnORPAGfBDNO6dvxbDORggiV0
P1eCmTT3wKuumaOi+ABnu+3Q+tzqcJ2b56wteiATxEwYTLzqeK3iBPOjtynkG5eC
uNz5JkPWzDlsShiir6B4PK5IISJqCe3tA4UDhkLRC/HnI33/Fl9yzh6jnVMFWZ6n
O6GbffUjdEGXX19R9jrh3eZ7hnr4LAL38gY/sl7ai0fOcG47w7RGro19JoynzqR/
dWCqgVpFD+7GICPf49ftz45L9SszxBjNn9fH4zohRDkBNEZ+V98JhSaILKzJH9X1
arrm1LXI6FXAaU2dk7n5YxUN1eXoEvWoahS6/+qV6CLB/XZIJp5FLlw2yBDIIljj
YHyNKH4TAqHeELfbdmDNt7F7M+9IowfTJ52zW5ghPU3bEugMpYCBkigcoc+fVzk3
4KhSqCsJyQq4P70mGI9zllD5NvYVs0O7rz19NzaaSkaDTusqJGLEvZf0y4jzZIjm
b0Tu/a4CFnjnf23yrxNwkuf8YYau59YqWUjWS4IvaBp5UgHJNM3Vi3yqYQ76ia0a
cq5s9X4axhmd2ED77o7QOqeRCI6CBK3SUbJoaBJe589A2kkjEyOEoNh0hDEjTZOZ
G3uiTrWsU05yPu9MPjT+Z9D/YB318Df5Zofh57Rde7uFgpK8/fOgQ7Vfq2ePGT7g
yOFiKDiAtfBEDA0YFYWuDUSYEFTo9chRgRVL0La7tLZSRTck/Mz97C0ceIYtK05F
cQaGxrZTg+4WIhO3vmDdm0KvFU2N256hTyfqiMN38nQlGLW5ushDUp/hJaHqqmpK
9EngoPuSR61X+sxZyc5HKvO0NciyCefHaoCtz8YtO9UMgik9jJhdpVw8bBlMZnbl
aNOSMhCGoClz8GUNtTsZC0lkXS9/2Zpj/TwCMTrMC3J8nQvPY2PST1bvRz/wbpzS
jgIoK2b9CxhKu9oZMAsPj7y7bErLDjErhOfsBx1otF1GKD+uaOV6ac+jzjQnbgp7
SHSXNhc9Ri1ERf8txKNn588sLLE1QyKQhsx+A9U5HFP4KlVkcdyQ49mB34IS86M3
RtJvmammYCs4g0LZqL8rVhwVL2YzgpJvSYHkDR8KZOWbHa96ScJraGy8Oq1Fjyde
SaVWv52vStMked8JaPbjR9QFZvyGQ8MQBaf2luvbngSF6MvQsSvaGR/aQM+Fa8tn
X71imMrDCMyPCbS+5+N7GYJLJfiRm8gwwMwq72q09aSbQ8I4FV7EVs9d4UZHKRmG
IWMY4URleKWcza5OM4/ZkQY+knBg88ivhwJKujrZKOH7iei4aJ8mdwjU9F/dOKOM
wpRuXY+5Z7legVt1Dzb6SzIp7PNmoYG34BBl1lOeKLoLIGipNE8YVX5r9veDO67M
l14L1aoZQJyaASrL5T2csGL1Re8LbJ5yr1QMV6WKYwQU7ee3vHGEp/XG3pyhVQOU
hwgL8u/bKmo3wTF3zrOK7it8oeK5EE5oLdMyJ5eheXscKmznvmLvxy9ucy06voMI
lkgd+VaAcMBANzkDVue9tMaUlnC0ceeJFDfTPupV4Go9reBQco8IAol4CB+GSF7C
0kH6sZC/QBE9OGC9nPGBunmQ5Nt4nyr460StKsdBidvgstJS6IVFenxJjy6xHv5m
AS9B07oGeaZjH3O5Ii7504AAt2ToFNtUyndZyloaLBduPLf27wcTGCG7ixyeEUNO
fd2/tXD/GV6n8OYvriNebJ1oFipOcahj/sC4ROqGOMuF7MMlMPJCDeUdElbIPbat
Ft2/6ekQviQetBR/eRK4E61b9pIwV6Vs1g0oL9y2wx74DcM5MRq/Z1zVPYvOq48G
mf/LRrW15rylMftvG1W98gDN26ydZDe6rRGR1D5Wcd2hCVoADE3zPlrSmwIzxUYH
VbaLE5CdBe2h3LvuiURIpMcviy55q96BRqcEcQ+2qaKsfXlxji40+ji+aazJeo3e
plg64JhbC3XdliZ9BoVUcBNLe/XAfa1UUQ3CEmtuAvhdw2WGqcWrUwKlJPtlaG5G
QmtECLxrFlbPxikxbxfmkq4RNiGfPiDjkjIPlmRzlbtkxivTX5IviMtQ4/QpaRA2
3SmnehHbBSKZca9qyI49yXHHeGQREzITrLQnLtHDwIAPfPX988XXvaxhae67ZO8S
szDTIBgVufku8fYOXQqTKK1bxYNVgig5fKjOwKCYyWOLf3nIMYknZ4tg6erZwxyj
IOJkXA2tQiZpzEnih7wuJ8X2TCwsiGbpRbS1S9A8nPvdaEo8V/h6hfIVoY308Srw
o1XAT48BMI4jTi9LYFFcFcuqR9G5MwsjNFEgy8ZFwAdO3+VmFdviNZqEsO6jHdkY
p3aN1xJ5QptCz31T+llEbk2vcWsGjxeC0mh5LjXqSluxohV+WOmY6MoMChNOVkio
Xcny7J8GK96J3WPDTd00byUVz8CMyh9fngnNdeH8RhorRZ59WP0cRwuy7iQGqJyv
2Yv6YXYDaU2crW0g8sJ2g35ENkUy8UyfhqoMwxI1I+EiFODdg0UaBHMAmlZl1wfq
rNimmUUvo2ttcSQtQxgw7T1gGvvHKjxJx/7GlzLxFmLXgIAQH8iegMzd43Pf1CoT
acIgM0QrT1SKnfR/lu1Q2OmQMcRDS3tK6p0MvQ+QWFlP9353p1iMyfIcwzG6wGy/
ReLvxjWcLfRVjl7SQJnQ0KENOFoiOsiDHkJZPU6y/yrwWfSwXtakEGRALDHvO580
c0Rduhx5j+cbVTcABb5CUuFrDAmEjLyCjh+iRCFsPC+qWq+mMhyXp5tFyI6xtf/w
TMom6PLJ32Vs39QY4cr6tXb9Sj6RZT6pq4B9VWeE5YCPFANdMHiheka9Ttbt3re5
nZomrfh4KXk3wKirdFRimupwuhq/wjKv5wxliECuoyMX5OovAAEmCsAYUl+y496t
qHW9JiXb0w8PQwGBCWvDHLl9L6GI4YVkENXRUzdCHE6Ev6ddVoReMEdXzAxOlnHo
98UE1k6c83TqP+pBrpF2vKaG5bjy8QPa6P4/rYiZhjbrc5XsaOlvBhioabdSo915
eHdlXhqkLvJplrOmtD9Ls+Li7UDv9bnPcMLVSDTGjio1H79GQpCOU2OYNkf4e7om
yj0Ga+sToVD4dDPwT73V3vGSeVGgPBq55b7KUcGpqaLvofCr7EMNjNRA1+d5y/W2
mklm2IdkRhn+tQGLQl3Wyc3Pn+KqdnaNwl4OTIeykga+0sdN29vb6D3yYT/uzmTv
ISVAbnkQGtBLXN3VHii//anmfBuzWXQpdUvRuz8hRXXCg8MILir93J4lRpDA1QKY
zg8Ft78bH/iFcjvBgrgenr1phsgizBXa+KFK089P2EzsPNhpV5OL6rKH43Vvw2Kb
aDZgHv0NI+chGAVWpbR2Nhz5OhjIRLoGTxeJozmIyiNJpUWeSIu5TlEjvghDVsr1
XVZcmTz9g+rZDzNwQcJMPmIOdK+oEv5jUmTzFy5Dtl88Ixjgr5UvXnsNuoPt5vfu
9QI5Kag9ck4zqiW7Aa9+Ehs68SGNBdn75wz7WixeYk4e5cIgR9CgGD/viiyytMHq
QRJ94tsClFDD+YJpLRaOPavWxHRq2bzc92hApaqnzS2zv9rsm7aBqH76NGNsLfj1
1TUopUn+3t2+VsOCkNGNA9r/JVqY+K+Q/gOAopmgoXLBgvVbIvXkdevE4K3dlrsG
e8cNG+dxII+h7gLuKLsNxaPV4XvWgD5M7OB+GU6TFT/GFjuV+UTeQXRDrjtQG2WD
N/rcqWERvDIQg/U3lsKPw14yqUY8YsWGKXo1JDoCRn9fcCqhRSFMDPU+95Cau8A9
/N9fESPnKxjN1zrbnEr3gEvRSBQ1fyTgbO84imlrqbRPlJYPNc36lWdRbTbHwTTy
b84YOXesdvR/+XjdB5Pq0Fd6ev/XJWlbZy1/z9lRfD3zo9IcVWnlqhRBGa0NJVAk
Kz0VGPj/7Cry27tJ8HN56kS4rcGawByAft9dxiQWCQYeappW7Y5xc7BIuxzx9+Ja
X3HDxwvNuMETGHIjqte3XNcxxgH4I7ETfs5biE9V7zJCD+RnWzaAX0vTGmvxV4sr
KqBuOk8gnV0Vqnv05E9HUpP1ei1YD1GybwuMuMn5/vpDve4yQ8fB5cRSMSlekXmG
famUAUFcjBdjeFt9y5b8aStdmED3Ne/8VzHvRFRwJ21jkIR1HSAglkV5p1RlNS5l
askUwqwstylRCq0rFkHazmFyq5OglCGzZB3mCrrZ2AzQny1qntliSVkEvO/Sajsr
yWEg2gu5IGX50XEudAfbHhx1y9BO2yJy7nOOyqkYK4hU+WyQu5P+rvC7cSUfKdOO
uFgEJ0P5k6uD/2mhk40nkwNQKugvSwUYoPCoecrLzb09lQaW8o+cBCFWa20cbFGc
FIFRtFQlRJ3x+c2Esxu5k3/Ifrsjry46+PsKBqmnP5stOR2kAJScBMU3Ntwp0r62
Av3na9pNCwboKxfTs9acZbCvlTL28Sly4Ml4ub5EeH3zwG/LA7iXTHn8KS3ASzXZ
RJfPkidbbU4RBCDZvD6IKGpu0ks9FrNiMdYGOZKPThPC0imDMDv39tvK/9PQL37J
40dt9pyhxubV8xxGAVseEEp03h4kQRnqktKxP1Tdg8KbvpHCi2pAdedPOq5soYFl
0NXxgahQTgwm1KyGwoJI1RqoFikER1CPek0xyNDsQ297RMtKBYO32UdK+Tno8cRk
VI+enXssN7xK73NNriW/tkhAy/w6z4kAvfVNvK4N22xwsTeglLFOhg1BW/fiKSDv
7fu1Xg714aMOlp5Y8KiioY+Kuck4wBuWYht6FPSgEDA/8wxE7iwNzpmliOv5kRF5
+HnXuTWrLXvH26cKy7Y+bO7S7CQ0JEo7xImP7jVZh3cSXQDO3aVwPXkbwnYN4wc/
yPXkVzWACGNzzVv0TpRSJy8iacew2PQvk4H5agyqO04Nn3JmuNMEHmmnLm+I7/x5
4cTFMVUO64XAOWWl86xUlSXvJww/ShCKJvzLcsgrSIaVxQTDLiyyrUy3+jFP+udQ
0tBZ6jHycZ3QTkE+5DwvsRjHhZiEKHT+4G8RxcPParBKnI6EBHbJ3lDglGoPCfky
fx3Gz2EuzUxr4GnaL8UnGfT7IzL/Qu7bOlPNUpccCumPvS2aoFYkKQafOs0+R4T4
2JX3Nm0T6PwqdbeWj2/F9642P+yEeHDHUDUddjupGCzoQCUNTjuGcdV+VweLDDq7
TYdJDIAb0jXfIZrLxO01NODqKcdDB/jX3vbqHUyV3g9T4ixImdLlUnc/UBAAECBD
wqp9gjVsyR/qJVCr+cyFUlJa+P0cbGzi+H6lQBE8FTg9PtBFPoBK/E9ImQ15SJgT
zIINYzG91J/ROFl8xpCFCaPahQNPX13YML2yrDUFPsD59mAkWffp/e+lJRJ+D+Bl
QlqvKMwD09Mc9/q5xm9Ktg882HGnwuZQIsbB0yiLxRCsO7ydsU/xrSxS0MH8/CYR
/eSZjYVu6TpqYcEsLZP+4/lZa9k3GtuG2hot5+OuTp4X0SMEmhmmJGUbLdk83HlE
5NnJ2/yeOEtw+S0zTOJWgvA0ldOMLD2EqolL8pW+hkgQMKTj+ng0v59F1nZAjlyI
eJOapjnI3ZmVEm8SEsNg2SAW8K+/XUPgwrVH3PjZzCxjZMqLwE4W99nEhcOt8bjw
ItAl6f31bE50xnaYmP+P2orZWsq/WeKjeqhg6xejK4B+C0vfrnUD7LpVm0vvNMsv
1tLaaOx6AQxCBYClf7ajLbZLYysPNgDQMu9dD1BzVTllWjCMO/KZ+qTDS87fGseD
UIcXggZdIbJEA4OphF0BidFgb3QMlWDA1a/iDwR4AP+PRsP/lOTjpxKU8gaI/PC/
BWVtuIb4CkWXz11InHy0lZJNrrLF3NE4HEBNxK6kf8aW8LyRzTPFtfjjLmuK6hR3
SqLjMmbK/Hj0BvuK9JfRSpc61dJmS+OfQWk3jZLcvYJVpU9DSzvvSz688IgVi+Rf
aa6L1d8Bw4mK+8cWgtLgw2jT5uFGOZ/XJnG+MUE8ZtuD+8a35ZKw0cWvlcS6BPak
q740UkAhgm42fCH4xPm7HS42HJ4hUXIy17QXOlRD13h+x0dRiJUdlaSflLVQrulA
dpU/nImgBDkmDp+kQe7kxIgbi4BxxA2GOYOJJbcfwfdAFAnSwp8bVqwdhrcF0Kq3
L3rScp4JNkRNixzWVodBFzpXiKjfk2R/NBKvMHtwHd+NE95WnkZi09FeJmDm4yUy
5cPhjIqfWw+rIqmoYNEEChWnDj9MXVuivjYdgG6QYo7EJ3bSAh62wrCrdtSKCFXa
J+1nfLGOS+tGzjOMqFwH4MXA5cJvkrUuDzavhO46rEi9bT8QKY40U2zm4UydHnAN
2wmG4geqmKlTFC0uFts0ccXcIRhTJ//klpZGcYZ6/AewqL66WoOoK4OGZQjsM57B
EAhnL53ih0n2sCW7JyoMbmg2yl1V48JLdmN98DEfYURBu8naAZgwaAdx79RBmpjZ
xlPHu9ObhcNTncP2sL4PIbu5EHTSd3Noc8GeDZu5agoFMEyawn0fJRJQdz1jmLdM
jFo+/EQmWCQ1jctSeECEfNyUBI6Zy8iEN/1bleiS+dpo7ODzActUug3utf3GFgiQ
sJvvZ1SgzlWJGsgiUG22BRgeV4W+PiOMhXmUvRTdMXEXqcxx66N9XPKhYIK09JKv
I9dsSKWh6Grcivepkmg2I5SF8yFvPhxn0JP+4vnsx7yzz7XVUfi0+I/imt0MATjW
4ljFYI5DwmNxdPNV4YdsQPfYoa0kWdpDY9f6HdTj+ZyfN5xx82/JDTJipnNlozLG
pjKdkT2YYcNPyeSdhA9C5GtjVF/WAO3cRVfT6S/BrskDqEm7VEljE28pFm+XmEmU
hGs/dwYYZui+AVDEhKQ475AHkkO3rzCZxBPECGcvI3KuWg9CRq1hOF3JwclM0jlL
/yYu1nMJB7lhl+EZDPInJftIbbU+jl3/h0UGlfSVaUEqkAdwOZM8of8ww9PlmWQO
+IOqEZhgaS8PnrlSfIt+2fk5yAI2PEeJ2EtPdn0hG+ng976RExBJ934w6AH/kusg
LJM1qtbwxZZV6HV4nbpSlQJY0mDM1v5Oz9meTSBsftSpOoPziUtIz3lTO1e+9ybD
f9qeZKaLHdLLs1auHkB/zquyZdEyOrbZJRRMpMfd3Vd2YQXpQucRz2JD9ppCVv62
4KHCDGeNUZsFrvsOtmIPkoEPhq3gPd3xcg9/bA5TkEMI5VZlxLNlgcW0H6wsref7
Ry7ayPcBIY5WPzEGgUnL69xxCmyJoL5mDTUuigl2yXQv7sVVHbNoTFGZAZFqXzCb
B98NaxeVw2znqzVjVz2wkmtJPmAI9RqKSNQ+3QKf+jhN0aHh2HrxamyTrp2BN0Sl
EhnhyVq3Ca0Qn5j9Ucgn2ssZRmYC6/z/6ASU3lKbRrDX7MiihdMvLTRIEMLsFzRP
xIfQIa7ZUpl+W8gL4H0Sdbd6Yb6+6PSLBlFdFDkPob6C3piVK26oselcTXQ+bgGb
9XQ0EMho8EXUnnhoG6gPKZdPi19iqT0bCEoisOixXxhk3aZPEXOM+CeEk0SfYdmU
QYic9BOXiorgAk9CTkv8wg1jI38Masu6NTfGWiqPi8FPNFKKujal6kHr0bQ+3/Wv
/mfPkj7HUT7VhjhpnCc5GcyLwR8pBbJM4z8keT+QmBP5vkOgI5fZxfo4bvFZioWH
en6AycFC2muIcnsgLy/VKYPXmeMoPhF9p3SoGxf/9gb6niCRUm0ABmjX3cgPf7gl
MKmZYaw64n8osbosG6fuz0FuyCtjNHBoQ19wCvQZMq0kZGBkA0d6Eh7Xz85PMh1C
++g5rx5hpZ60qvjfPxBaRrwRhDZVawuzNAB82L8OZcHm6YNW4V7p3SClxIcZqy+A
KcmMQtdnhKA5L/5WMjgb0fyBlueL1fFWh3gob0VIgaramuTIW4w17/yU8+Okuo0n
UFedeqGTSt8rKLuSTtZMrL9uXUyGq2MeIVFjgf5GERC7DDjLy/8YmFDA8p6/RkuE
pFsfl3Qt7sFv8Q3CYFmRYkZQFoJFh/rkLSJPBZI2qvObxtQihixJmx652rmLRJjy
ur2QzZpbv4KL/vFaWqFXG7yjF3LrsKR7D1HIAYPHQ8xou6+wQck2Fr0FOtgtl8xW
EyDF2Qblox0xGCpC2YsTsMHl6UXMJ7+0pl9z6Dq/gaWK2hZGcHABTO5LKgiHa31N
0OUe1wbmdfTGq1ujhEOQEpfVUmHeOfdQObZ/x1aaZtG6tTuZVnmGMH/4sZOjCyAv
Kv5lFOa3NR3Llr+aJ7QPmybg0vTeYPajYMV1uMSowmniiUlQfRClPh4ufUA5sQ61
ZA6K6zjtAkTuWgOm42i2utpWVERwYFLixmrf0O/iltviAqnlZiLGnKaPdtMhGmVv
cjtGujusWr3gcQnP/hE9mkc5IyApSbHC3iEPoMG1istvDUkUUp4HiMLsaIlhgG77
Xs/arWO21MNWD+pkUUmCexYUPyH0Zf2+9XhRajPeORfdksqVrz/ktby1l59iN08b
tMAJWg72hvpKgbdjHYqUxxz/X897zRiRMaXNp04pK0RBlBpP5v2XDLIzmddDcwlS
9k22eGUCAms7HMcUkxOiSRimp04o3piRMMO9eMZNx5CzhrrONf7hgp0IMZijRqC1
5WUPmjS/XQf7Fmtm8eQWAOh2iahU8tXwc2EAF/SaS3ey60935K1F5RcFhf9GCiOo
xY+KMnYwxEbOBmg9ha6gotd2sz0H/Be+fwFKGWZRbIBOWALKuASv+yjCD3SlOVyP
T8gY0XfgKwSKJ0wJB4Yb6Slu9ChoX2PB1pu+jMiHNYVXqeiqiYPu20PJRixWBvmj
7ZVt2lC9zbBpTGuS80klD78PNUEKhvAMDlWpSVL/6LaN8+lxrTHQUVWMlf38n3bX
PQJHK7RKHac+HjaNd0d3sA7qAZcH5Fd/n6JsvLPeT+iS18dB2SSGirPUATv/wSRj
gXAtxucG1/DABHp0kqYT4PftbHEmKItFGO4xH3dm+zJN3q9HQtaCxVscLh7t7O+A
10KevuMrm9VY6lfn9UNuWrnF9fuuNoY4jNP2Oaqf15y11bEIuXgQdWCTO5ks9Cie
Ys1duD55SnhlP7cfO7adaMTTQjpc9eZzesIQZeNBGwUKacUxSiW4UlzSkHPtH6iM
aSt6mavnQR9iVT7YNPB2iXZZneHKJIDpabfTPa2KZjnhmLAzCnOxbhYZfV+LEgNX
84jqquBYe9LGvOBMH/x3sY631LjSABfRrOmVhZDKUZwtd9q55WN99o9/d4a9SD9Z
DxkZMMHQSyE1p/IClyfDH699eknK8ukNNNgf5+Du30b0OFMLCEFMqiz9YZDftqZk
DpfPsDA0Him8f2OqppLgHcSsPSefLCFo0DDk2ApPY38Q6VQULEpZFsRb9T+uNIJM
XoQzDfp3AjCPSAJT06JNQSKpzs9wf6mVviE7pRLoWUXpaseLmPymO4jFJkfX/aXZ
oHSKg+VQb5XaedkNIy/AxNZn85xFt6x1Dio21A3bfDACSElMA+vukXwWOjDW4E6c
DlkcfqcJbRS7rrSnh6jkTskFQjE7dDxr+BjrYFIU9oLjuPJqd6E9bYHv6UkcOjIU
3zehUrodczoWV+z/7BkoeRuKFGqkVqpRKlavuVkaXSqXYl6npXFaSQsMENUKyAbP
laerER1VjcBH4D74IVvicLjaWHj8ibbtjJNP+JIUjBbedFO1QuvWMwyVL6qmftDZ
TOqUeDnLN2UUulYnkx7ROEzE0Sa7WQJlflv1k03c4mWsWQFWSSElBNCbloZuVDET
2Xu6cYDYj2F6j4kXzHTWwqU47mzLRdo2om1RuOTf2fwo5iQDB/wEIPJY0BtXMYok
3c+KkINNDYx+Ppd3IWby4+Z6b0le6YoWJKj3ny3awbLn7VMXxYU0Bn0jmJDAZ5Rj
d+2r9zJbCEFnchymgiyofKdepPvJMmCblMueaShzrJN9/JZfkMK8lKLcnOadQciG
J056fImfb3VBBDQD50emoMyXRDEt+pcz7jyuw0MrW/G72bCayz5nMJm0nwLoLi0O
FXx5c79bJq51hkX2k1SavxVUVFwa6qur0SCw1L5s3iYNj1I/ivbCFvfEmiTz8MoY
MuC/QJsY++2GV5ypaMD4qbxb7w9IhRiS1g9ABvd6Ds90BzxOZ8C5x/jxtE8n1ET/
gHsgyCg18tBTe+G7yAXEjKSLSQ1RjGlpGXMqDTBao7l+WmdwbfnTQFQTVv75+XRV
FDO7Nbjdjg0pUbOJ05brXfCDC+rGRN+6DgWlJux8hQduaAdoHmoUXPPlZIO0wi4M
LINqk5KOquRP+Zu//N9AwKQ4x9uPWO08k4faYM6TNOu1w18HTcO99Z6yARQ8QOag
yFCyanIfpCpC/kJ1jRiWge1Y6SxYyyNiBOM9INaE1xys1R3p2HYkZgG9mhfE51Pc
VQFRrwf6aIDUMa8LkoGZiR7ZuUdXP/ls90EDl+igIN2tSr+RJYsEH1gwPVUJ7CEd
p+FfGeerUQYtn4LWfEFDoA5B5FhskNMDsQDFURFAACwXA0D3o+TO3uzJPyt++iRX
qIgLrz1DTsDRRvVSG4or+9X5Av5+JzxBQ+7ILwoj0Tn+zw7MpaXFa+BwLmWYnRrJ
ffF0YQjrpyNWFkTrYmA9IXe9SoHw1HEtMQHCNZ3Perv0rkgiX713UBo86NfQ/EmX
fRq0ps8EzMA6njhyVt+Vw8RKE/mN7ziyAHlYAbRHHkKKrRrqZUbgekdSYIdCOQmT
eiH2c+LaGW7TvyZG47eGqwq2aT2t7Bdy59LuqDyZIotyfkGA7DUtr+Yh1G9N38ea
zvy8TBiPzgDAFAcLvFOK440MEmO96YAAP0XbQjy4lFIzEytKJAANH+fX027A1zTp
IFa+I6OLxJ9Iw4M0hQzJh6sw9ta8nTRmd0BewWjxTKe6KF9bsmmDa7ZH0/p610ZO
AmSUrvW7Ex+XZmp2pCjehMVZOaTmopzc/YhYzCgw2N57uvM8RrlHE3hf53igi8La
9W7Q1BUlz4Dt+0+bAB/gRHLBf4eK211Gaa6i7qNBUYRBAAcAtb5CqtbdAeQ13xlt
sBq9qrEy7kNHnQyreSNTwyxmaHIlkmu0s4ZHhFN0dt+pybBAnxCSTEfCnaJp/Vuw
XKIN5AifixtBXvImQkYtxY95mWxuE4yn4TGhmiE8JqIEPVhS5gkCjR2X9fC9wBIj
cN78VFq0TvuvSuAlHljeOhdepR/B/tNxPhjaEjsqRLFdcVQHAmDbUkey/tFgAEhU
UQYmRj3D2oE9HvgVE2x4ebHsWLS0rs5+esuQQfAYp+UYidROL0Etebu+BRaPCh4A
CtuqcN5YcPE1NYqOMTiNta9aM0i4cuXQB4Qfr1Ki6P6VSTvHbpOMeW+IWY8uyGVJ
WWuST3Ne4we4p+o/cgq7u5RF0mtGjOcisyKfbG4dzranrBLQDPUxwC2Ip1l62zD6
f71dUnVG5qSSWJZNNfGz8FON6vGoyMH5xjAyGluyDDUgXfUItLF9HtCqBP7Hn/oF
FYdNL5YhTDU2BzGX6zglI7XzSHK/M4192n6IAmNczhzWyfX2Rb9snzi8fVmtODrZ
39+pKDb7eLEuyqqCQP6Cch8lmIOfQCkgKtjkifO/b0UwSnbuVRkYyW0hPXmqDB5Y
QcCMQArCc9WTobgGW6LzN6B8ThXoXyd8AN3g6W4suI+qxjkMVJMNzSCDilYjT5wo
iZl1+z3Fk85JBTKI16hlZmKJx+RZ/karP86KuiBdhO+71OszirnNGYkujio7DZkZ
cijW8D3MRUuRhGIMNhMRTo04QYm9aW2yYL7eCn8zan6/la1rsxkheq/R4Xdsx3gB
csBdLYYBxFcQe205kTv3eEWYHRMcUcSS1ntjPasGgKcTxxqdRL1jWReUvbwEtoW1
ouhT4hkkydfsZKeTzbvrUYoTx/DyUcFzf0KuWjhkwCMSnrQBd7dqEqCZt9Ok4+KE
m5rkmhI5UmfCDHnG4IglNv+Ay+c49RhFRpgtpB0YViroDpBCpDu3yaNoCHywOSxX
Bo+imuWHA2oMXacz6+jfQDLoytaCgwwszY+ShVX89BfieuwTDh4/0pyHYCIno8sq
SrFLt/kQ5cRJZqGgylFU4bSdVEB44dVohtjYTBBQqCFSJifhPkX/jP0/RAO/RadX
5A1ShXXfDUyipOEr2e9gepwVqVO6RTUcSKwvuRet7Odtk2mnPC/STai9LiG1y5PM
CQGNC/GOwznR5KT7bDaJQ1G+GT+YoZ+2n3obbzGVnIkA4bDFccMPVI/ysbBx/izg
svSbq9GatoiyFFQ0oKTiKaifGip0TlIKd3/Bx6CSFOnS05JT+wo+q29M46EXJNJ/
YWwnmvWB6pSrv0UM60edgl7xpQZl9AdHW8ppo4hMBTTg4T6C7lQZhRHrq3Pi0KT2
7Q3Jok1AuqXYLohP8y2YUVz8GlmzpfV/Ojz9Zph3DO5Qfd6MyWyOpngJlWr962H/
XuqyvV1T1reY5mvqZmv+DRUENgofG1+fejrv/wDFsNe0sMlhiaBwwhDxILZl48+I
p6QocXggfjeIhCpbOiiNrB7gDYNShrbAAb3qA2ccsGE18skzMoV3gV8/RTyGLBCL
uOH9XH5Fyf6zXeSYa/SM+ZUAUtNxuOnSGgNPUWm2o/cu9Cu0vWSh8KzPqHCOp9qk
JogTNq6KLjqeCklFoBRwk02s1kqQyrbV/5AbmBYAP2zAeVIzSS6AiglPYVnwhAqp
SbKzOEV342Tijs1wJi7WtVgk5VUMrDECJh/6i/h7Acfol+APcEjQ4lwWsoxfCUKi
vgw73P26xq1TzD51owTNIj+SitYBOQgPYTPAVqhAieuOqi+jLMFx/ewdJ+Zh6+0S
sPHc+PJf86vO2SIYJ7Q81CsjwB7ofALK+z3FtxpgVghxC11zusDusPUiKVFHVIM7
AejJKAUPvmy2pZB/M7ir6EmjkhnM8603YKBmLtDJFOKOIHhfmCq+NCCJNb5QFt7o
PBiENOxY5y0JZWVyZc3+6Cw+8OHmSDhsEsmh+PZ42ZjitWPeIuA9sDgDlpa9Nl4q
18hvE5qIDGJ5U3wRdgQbzJg0CQKzy519eUnf9OZMoaS5HY5CvF1lxzBtYeIBnN/d
zXSGLjD9IdvKv56ppoy+9/iEhtswrVH6s1ImVIntYqMzycD3t26oHsepbSmp6Pe9
Y6oGadbmNEQ/Kd7uFOsDdAslh2/vXHbk8ImOIOp1WKl32asEU+CPdpe+lf9FkvvB
7HT3zrLmQopEdPnuCxLKcfD5gQ/WLYYG6jnzWkIVSjIVzsesFQIB0cTuABPlLZcZ
mtSZJ1ZRgy+mipFESb+Aj+sL+evQmymiDVmjV8lkdZj3rpPHJ8NKnmtiOf0DA4+o
YFWvfgzG30axGK3AZqkA6rBTGulMJHLjvFkFuBx52Of9hFAnReU27qVbi18h/zxH
lKHzj7PgYD31mDag8LKbJWnrURbQKT1kVWR4M1bCtWqRIrZr0HRnrFjpcl+96AnY
MlgWx68J9tNAIKqkIIwznuvjKh07qVf7zQrrYmUX+MaijEuykUVevkcwhXIF1AHQ
qcStJfjvgPif5b2+g9ibk7IpqQdwuxrvaGPuYPXekMVG+7qMxIyor4ENT6l6XPMw
ZvVgGVvxlGppDuoQbZff5hywloIt+BySL+E+ijSvVPz+osKO+3LyCEIJ0tSKU8dV
DTxFdT4JEVUJv4+UsxFSLL3y1ngkpLvCZEM6YSm/mn8dEvjEq/Gb8nETGiyTvfnR
qU6MQfwMkmUXbNSWv6JAnhP4F67xAzpiB7DaU7bpsj/I01uSz1mIig+iwOPpx3gf
GWblZcDYt7wl/efuy+MaX2hGLK20FG9NOBsqdJJ2c/EYBA05STkgRHHbxD0p31n+
kO4btpsGJyPrm95gL3qQdgEsSflcaHN2sHR8i0OtfuP8LtfWV8Q8tH/weqvC5lBM
zdGw5fC/hupQ24mDNyp+D0L5yI5XbXMVffXBrzMfztLzm4cr89nYhKYmOM4y8Flz
ij2hF0hkgdUSVv2wJoAgIX9Mnrybx0aGu1GaxgatUVwxH4NDq1RodtLE1L3PVJu8
AoaStoJwO+0LO/I/41ksXEqqn809rR6B+XUD8EU5l9wxvDS7Cl8ykbU+JFBkLzNC
RL4Gc7RMMN4puLttkxCYQqrvvaUp63WL9CjMEbV/At3l2iQk8Ci2MNdRuoCbiMvk
9zg5ai7Vdg9WLNEmkenQ3QaX0LYVH5zscZmXB4dNMGN4X0xDpCfd2mXUxKyyBSUM
J/n6/Z2OK7rJ/J558dm2sM/dk5wG/dxds70KLt/nwmUhIWE0sBmMxlYIaVRHJIx2
NsPA0SNjqvEKLU0j7/sy+R3oYwkLQgX6qs3mchtEWkjtHbuivtH4eKYgSCgyUBYq
gnJ/b3nevZZdWfGY6TTYo+zh8m98Zcj1T8VM8c09AOlA9oV4qJ0dzzyuECiEt6gW
VwE/7oxUyEK9VfHNjCSNMS2+mIQR+J3Ybc2C984i+msGz/ITFr7OPOWcefakYz+O
UxMFEunePzQB6MN5TidOiWZEDPnWmRTSAWCAOc39hDK7wQkzoudLh6bmVSf32zN7
S2zixjXCx4qP1Dsshlp0DAmuV9DygUUWZowKHsnpGe7XbHkKa2QjDodRCYYEyIlq
uX+I7CynCCcWVEMLsSGaJVZWvrP4+c5r40sO0+0rpCGU7icALxHYSSVW+P+8xwAJ
tPcQs6vc6aZQ0PRWrjPGP1YznKxiCkAGdxGZq42H45TX6obJJZ6oCDjTvPedmt1d
Q4Zoac8ZHW2sfgCwLwKFwI+0UPqRO2uqejnlmwdSlawj4q2FVwHLIBwVno6yq/3d
oyPJJLrFQrD13h3fwufWwlscsEMIO2RF9fNzUCFKGWZ2c80dGnMqq75NhPRkdbBt
RBYh+KqusCnt4woqT4qc5fS7FniJGMcJbUYGLJSGrt/DYcbqgKAg8YvHbZxuZ2cJ
5EYPdY2aMuHqT9esQEv8WksW3hNflQTYJFEoDLJsERBGBsJS5fJKPZUCXn9tRydd
B4E341JuRayOYgRwuIf5M/x8+51gB6Bo3VwIPcJIl4TSZ27hYEQ50N6AAKGvkReL
2x5K7hge/UIVO0z4R7bAyYrT9wJRiK9IGs4nYtNTUG8RSsc8EjxRIkIhBlvH+XyQ
11Pwe+5JMdvrs0VvUFdazfNqbBJUpK83+8AYIhpjapMuI8p2g1s3EGx0InKkF1Nh
VhhZfUksEmeGTCK47xYFIEcVSn/Dsn7IuJW8YeTlMI1jb5eMQDsvphEPii5gksFq
44u4zHr1Hwv7kDSVuc4T1ZvhOPJlu5ZbAPXgGFykiIz9UnpAwoO9OP+e1nmEzazR
8VBO8bm4WcUQTxTOGBp/yTuUjXlcYGj6B/3YqlSaMSgqjGiygAU2resBYAwg1zVp
Y10g0DLBcKaleJ244zhx7/yk1rcxztziCOEj3xzoHovVVljmGaPourSPZdwSQmlh
2+Y1FdFuWg0f3SVObLAKoVpM34IwNuILnALwP2iki6i9aHx+I5fv/1AuXbEvBhBf
KELuV3XOQ04dPaMQd3gDQaADgPM0F77cPjvH2T5QIzp+UUvvoiVQDirFhxABFkam
wCLJOX3Vi1YCvfTXsBZzG1kfWSAmxRSY8hH1nP/QdDJVHr+61RP3wkTrDZE4Hcw8
uWIjnAEGfzsokgt0PmxZqET3S7i9BotM3lrY9SnovC791j/zKGD6Y12ctLQFBYw/
gzWxe7vbb0xWf2dWrTDanGB/jgp5eQinwgdc8vh4ZLkBG1KYQq+aCYNaCt2GEhyh
/ZqnhmBwRtjS9ZxPae03FITAJPYk78llbAC7FMaDSL6mw7FZ5fVTOrketFa0X7Vc
LkvipdOKGYQc7CpnIKOLKPmPSLSCu8FBwGfVhlBdEN2CjRYWUR7UxIqSa3LKZAA2
bLBkVAdf9eRHNskfO4L++0nJ0TTLfjxhvAx26QgdaTU3Pdk19+lMHMdlYkJOA3C1
NPv3LIrH6Ep1l9CmobOLZDPWbpaBMmF6didJO0Tfpy6SzXSKlAGw/wTBr/8vRj5u
sHz45/vRyRxeWiBk4+J14N1PeA1rghX3B4wue65US3kznLPZBK00+Vrso0sZxX0C
FqOu2IHLL5SeSxaMb+j8qcIhT7oiwiddw09ENLJ9APS5/yCaL22X4O6RmdLN+5J+
/5gqAp3dMQxmfKsQR86NRmHI7vXcD/qglXii/X8nbe1yn40Wl9IuUpwToU2e3eJC
FcmbN4aoIjiD/AOOrIH6PFrhPakbrAB55df0GjAdbnRzUERHxd/N0+EaWO/rZzL5
1FxYfuA8SCR2wbxyPVby9PE/wLr2FGsKdtdZ1MgSfzIm04r229WoKE/wtvni2uLu
CvL1Pnr3k1MKErlGefjP/QUm//b1quD4zn2llrjBzNp3ClP504/uy7l/lOeRa6nZ
eCHTDOfRvRS3bUnhGRS73T+EynQCqr80OFWKlxLQ4qshlSialW5xRiQsyv+3282z
NCvHjkp+FZ61W1pqedIKbMgI/TaggmVzZm+nGaxuQWh3sTVI/peHIpx+EjAaA7Kd
RMWQNHXmDQWx7JbHfliLyAO0cPTKEyZIB8gajMpFPYizj5bnl1GtY4WZyPAajq09
yGGyNjfFddyej1Clyzk2K+cqJpxsKbgUx5ARKgI2BTSKIamezCZRpd0RML7zv4TS
b6zwrDP4sxJ3zXrxUr2O0+4BQXbJCJxRID9UAXmnwCsYu3KrHaxtth76DiDKA5bj
QlMylgfVfze6jD4gWt3a6G/4E3kBk1tzR5FvOuOxMhaRMq5YTIB6zrpFOWkQmlPC
xfr6uNZQdoaMoboga3Q7dW7+nmvXH0VahuyBGqULzdh82jCOhbNMcZq+ls8zht5G
K3uQ4CtuXYqhhtzz/cmi20La89ixMc0OUO5gHyKbp2B2wzNketm7Lp3RJvBNxWCf
v5aTcSIeQB1Wg3paS6v2LDjFkAXfAg0U5+gHCWX2zzT4wKKSzPytLfQhEazvldYp
RZOv7Ydl9cjjjNP+Fi30Qz5lSHLPMDR1oHAdn2egilQ/fpTvDYhXuerYEjE50m+S
iAceKDlbtron919Pg+q1J/UJX4YiQO1ouJl/Pjr773O5D9xAEkoUBwnHgYmwiNO8
6zQ23LaYKK+6JPBq/juvdqyutayha4zctE7tmV/0O5yBF2I9BTZQSKzo+3cF5cLo
MhPgmi/yA6yGYF6fURVbdS5zTCDAosxGR36Boh72VAYdhEJjgHNpJCM0mPpmLO9j
r2uEYsWLiIkwztX4ai5x94p1j1p8TJfVvpw9wgYs4rnwS2Mj9RXexx9GZVN/qdAV
1J1yewqQJosvG7n0v38BEX8gpdtWgKQTpBAShzQ/mXvX837H63Ez5OG+EK6t/tER
DajRFL4Yb9BhUWC+7Z24V9LrTLO2BJiHnL9EjkgujYauEEjahEb8Njia4FQ1E8iW
eCi2d8cCXRsKWpBaGT2bQYTYLxYseDPzsWpPHhl9LSjeAJU8WnRXsc+eYq36KCPO
kQ0iO4cklY+km3Tq1yc0s6FrWweZ31fh9xfd+1Djv94IXKTzjWYnB0LxoQ4XZeMf
Ck/6k0mHN9pBOL/UrneDjttinVLK7dWEkEvuFZH/Qj0p3jiQSSgExA1BiAQAUoyQ
2BGDyUM+vCMNpVEuijzEMY4ogMal7id+jKChpVTbyGJxQnmUAjFL2Xbzw5F/sY4E
MvhwhI3uyy1ZcTv3tI3SUIi9svZ01ZkIwyXRWTxxcNrXz3rjWe7f3I3+VCcSrYUc
WxMAXxgAzkRo/jLOxHJYCgYrs1I7dm25qa6b/EHx+ULZXArZ/CbD0mbk9m/wjVkI
+r8yLFyjH+ozec665Kbt3fHsKq112bKEar7pSrEnuwEBEybU5MX4F4pXmzdpSWPn
G3rqVufBxri0Db/Bg7Wze+oLfQSaNOBTcqwSatjvM9XojhLqZaYBhWOOthMIaZ2E
XE5H/WDMGJVSnZExr/GCyAHObmJ4fbaPY/wFYXxobvxRFFctgu2DJtUPVgSoRvZ2
I50cOQkd/qluaGjXvN/hrpXyMb+HWiM8KigF9qvQD8U76Fbn0JSGinB4lIK4wU1A
mZG3+gPS4Absmoe25MOhimhWDuIc+ks9DCJY6C18SyjeYtAVNlRj87FX59H0A5vh
pZRqlWaM0+KTsBaByrG3lozewg0hTjI/6K6gwL+PHgcY3kqZl9GjZ5a3ImwBfQr5
7p5lYS+TDweJs5BvQdQ+cKqyJZsnzJOMtZ85D1ZL4Oc7Ad1jjuOD08GdVnmUswqd
PVyfl/1Bn3a65s8mmsmvVLoxu5Xk5NNoIBLxSadIyQam+lBLMVkHUURYTPkaodGU
OGBcZ0unexjn54CKTBSB55leFjn0ufdtBLw9c2o+z3DJRrtxBIoBryfdqLNm6pd8
/lBSfv6kgpQ3UbZudhHhqa6Nvm92copg+mLAFR/9sW8tgfUtAtSFeTdbMr6L1Wlb
690NIpSBIX96tLp/eWD0YiZgHFQWa2qkMBNn1rNeRimCnjcCf21td17gTEXnnaLp
M6s11/r0Sbah1t82jLc9hiLWl/3/0zQTDm1eBxLRhbcTdlGP82mxPxijOrNdNvTZ
i3XyC2T7bsgk8dyYkuoB4fGe2S9+bWRFhVziNFjwUw9CXXis7IJ8DR37nZiQ7O+n
Aqo+cmKDRPq5yypJfdDl+vuw0bmlM4Tj4mTD63nwYWl4I0wSFvYjspOUR/hgHX1h
G2YUIorw6auwKgpZ+xKNvLkPhptIjU2c22mUr/9ntshC5RQA0PXSpeiBYaNoYXiB
6NGGwrJTSPiGUzrEINgyZaY0hvbu0+PWT3ozjGHhCZo46wlg8qjZ01/bdlyu628B
YXDcB74DhBqkuFX+XyQoJvMiVD7SqmZWtycT0+nPgViy53O96k7GKhClj3X9MMvs
KGvau16H+9Mtc8Cx/EXPCNcHqregrkutr4M2SLsyV7tHmUzGhlQWdtPamkXpQQUu
sPS4fJW19u7qxbVZaDxr3HYpEt5a4WVKplRiUmr97RBkRuPLZQDhJYRlV6U1TmpS
Fo9klpPz4Y3CL/uO/gt/xDHnkrLs0/d6IWD7lNQGIjyGvJP245ROV/Dh1iErS1Cv
3e0U3hLPbUFaKrJzevAAyQ0zZm643U99oYyBwfiXYIHgSJa5hCWgexMII9h6+c1R
yQpZqndcYoXdQyOEmZieZptq2yykg4IlinBvTvk+z3uv405GiXYMaFoqJlFsNbWs
24UQn8De6EvQydvDsmmUGCFnk3LUwnYqjc3y6I+fjkBUHMCcFePv9BVfssBqj222
E1vIMALI1F3fyrf3A2UtKDdY7kskKBOZp1BuQCd1SUqHBRPm6tt+J39hir/sur0C
qFRIeRux/gBNT5fC79dp/SevoK7GfgcUyueAjMenN3wLLAvaFmHoU2p8hjLWRiKp
pJnK44d5/E3uz+vKB+5BidmHzggbKPR/CMbO3LxCzuCrdsAghOgjMKiW0KPoivA4
XSZREkYk8Aw9iqa2mi8tS9uGHfPwSJ7avPcM71s6qc21iWjFuunZ3UeJWmPB1+s0
Pz1ybb3vBouPucKbLKUV+Splxw7K/JCzilJFwer0dkMW0T3STRJZhtSjz3Xzw2wu
WzuUxGnCZdWaviC9OmV4qz+nZxtjbaOy/bp7aAHn2DGwkk9i1luPQyU9nWZaPoLZ
ZDTX4iRvoQsjqwoH4+jNnbYvsVnpuAAJ9Dg6pDPcEB10sNdJLFiYK/mSYsLDCD3Q
fxqEOCDbiEctGfLNptJxJbCocIAHjJVFVeB33FP6aL1BqszjNV9kIrE8YjVtgHGv
qNG/z+XU7jQOzE6pmhojQueEN/5QVHE4HJJzwrR307DyizkLUpFYeLqO6rUb26Xf
cJH6avDblNRxPceoBP8zvVNEHTHG/M+jHrXjS1X4RraQ5EudIWvgDfZerMXh03QH
32NTx5y+uA8ct2pYiy7tEZwv3mb3rBTknXOvuSqXes3IEFRrmoalvjdp+gHNaUB3
eR88YHI3sCDYujXbEkQTpPu+FwdXY63LlOzJQJpCoQ27GakHIBDODtOjeTbVEgiK
aFeZ252EjxsQ4DYroth5voOneTlfnCve2nbKlxFLd31jS0/dGRZ/1FlfEfndl0Of
2xdx8KwMETvUDnUPxYnt5DtcIzdsA/3kTEBg0m0jmWN766I5SlaCCG2nhXV7e5B/
06wnrtG/VseQzcBSLVGEcLRYFmYnuXDnw5kUWXdndCX/GXKwCQVgzdlpcV3PbOU+
WPc37r8gAwtRIv1LtnanKLYNNgrFcxJauFOBFoleo6lNKONBnYhSrgogB4XvZuxx
idJYEpVV/4jk+sYwxrWJHUa42CHu/M1P6oVN6tUUQbGnw9o7/Cn59Pu5CB7EscV2
5NsaVdS0NwbSFNEWGDyeMbtyUixQvwF6do4LjrqJiH53o5xObFaYQmOiwurzUfsE
5C6P8d1mWxmnHsbBdYT3D5L8AXNIioLhh2hDOoT7UMbmONOZQ3K/zE706QMsLKV2
Ak9ndvfa5/KtusRAxZWf1qu1fj563XFa/T4fKANmSLqQ7+3JVveJrgQ4gVEhsq0m
BDNOhWDaf8P1fe1TH6WVbag4Ax7Gr38CqYR/Ug9IFbANdNnFWd+KgBeVQPWNHp/P
jDFYMRXudI0QGWYm2s1SiLW4bs26qCCajANHdLMUhltngNGq/7CAH+OUuib212bM
DSYGRpcV5SYAOYf6oPKNBuPRiZqsocdstNtU90RdUESL1xuSgCVMfFOcyhilTcJU
COsgzFF/UbjF3ccLNkpy0nvCiAZlvDb3aYmb/gl/CxooqNerc5Ys4pInB8WdN9eR
WVm9uJ5lTOEF5MWR+EJwQsKDI8X6o1H1Nvq+c4YhRZ3NITxdvpRiMi5WOEKksalz
JhZ+sTexLp1b3i7ZaJEIzXCOG5uLpIsRRPkiyp48F40kZJR5UdjGJ/5Y3PHjPi1o
l9xiubV/IFC38h36CifnYcjHIzcLP5K896XVtVMG51+bT8QJH9s7S63sKyEYrBx/
eii4iZ1Jkx9EcC5keCjQfjramniddODnq/wE4/iVXWb0MGj4+fV8gZ9h1KE8oCS/
SVpcftGy/cmidglCekPp0LYpOj1bIqCmsXpsp9Exj4ffFK1Xp1hzvGvdgWZoImfb
gGjeT5VSLafHku0p1L8xX0n2zPj1FWbZvx9Ka4bO9GZz2qQv+hZfnDwM8//xsYPK
A5DeYx9tnZNnWO8pePYiTVi9J5O5Kpjr+BM3tcgeiHQRMSszTjTgEVShzq9/ei5j
5q9tiUcxGiACjTIIz+MfpZ1W99R8T4xtxvxY+bRaWDK/WBEAngoCECjikIDfVCwq
EocIKnJqSJLHO5unSABZGNYsg0n16ZKAkYm8wzde3Iqk0YgErcStWuXjV9+UC7Gq
4dTWnv1+UFJyc/PvXsOrajYaN3JsrANMzig6EtbA6d3ZPwdpNRwW9MbvnrFZVZOC
3RcovJgHLXTEOk26vzryllEm5cTHBqj5C5AWCyuPxjsG5pH96joKsk+YuN6d8uTc
q78wSBDgkBuz/NiSYVGedn7ZLByCGBqSySKYm8lptx8GfUtmbU+rtkeyIWJIJhXy
fC6+l9FDHNDjidRsjCENRkw2l4UwjyLPJX+mp7r0gyibAh8r+5Gd9WuofcTkEgMI
HxeYfUeG4sr/MjRRAUAKy1cutqUwSPZwAQjd+4fiCcbIcVMGHlRFmzAmepoP69aA
t4KoBRhQ57cuu6/3zyYdNROV8vRHKqPzfiqqbBx4cxyyLA1E3jdwWPFqLjgFvBw3
EzjtApWFB9Kw5/toGLjaSCXOqhpKw982GWEc1E1f8YVf/1WVtEeQB8C1GqT03GWx
qTS+qbJVBbdXCiVqPURwvvDIARx6P9Gk6AAGIs/xZY6E72LB38U2yApllr14A0bf
9NpyJTfuXVRgj7S2kfIrk3BQ6iEFj0Hizi+DFZQLBUDP7ouUw6a8Mv4MEDkpKw2e
jAOsMm+QhemVAxYpxHMPoDBk76EpYVWzJolvOxdNhWyK/DYie5bzgKhH6TggJTmg
kYaVpqfOZlJYelOyK0LO2tThCCUkj932OMkkDZ3fyXa3LoThDUWUiFB+ABQLzIha
AG96So6i+zYd1wIoqk7j0TOZPNUMQZRFAtJvKO4ULV4B5X3BttqYvmLhv0FqAWXp
u236+gUi5t3dmJo5NmlqQRq5Y/Rw+PtGWbt9rQ8BhfRxcfkIQwAXnlqknNmX9IXj
gn7t6LMbTYylsEasLSTRMyJlm22BFIz2q58FeqFVK0wt7VhKfjbg+iVXgMs0iSJz
ceSHYNW/sgT08dnPeQ9uE7ts6tLNYBWgGP4d2LyknuhUHUmafBWHRGj8rwieaO9v
JqYSmiabhcTtyC+hZsAMXHjMlfbnbk0yLTipfrk3DgFYJXqG5EABvO6peYhJO6jk
VNQKdbPsdG1YFP79dI+QiGVYXMPTX+pLr7Mc5BnaebtEPt7+1ajF7fn8fczdR68q
Jb8/Hv0JUUk5ULtDcvqoj4EOw6VPmsiSf7dru80/s4jhzZqGcda9jikVPNJX7bM7
QpYRi25QrDqrC4SpvjeOeLtdV0VQsCSCTnv7gSiXdsObQTtcPxM+frZxaOQ4hd9X
MSxnW3OblleYvDYmRbO/57me6jPhwwJDOaM/UsRNZbNsqXtY8bnrIyYiXif7MQjs
MPuuCzzL3FKBTJ5RnXnFiRfdPYv+sXywd+PuhPooZF3r0JDLnSkS/LBpX15qNs67
CkSXpHtJfBE1EUUUWTh413+jzZCb6aa6Els4SDAlng/FHpBllOHCL0TzMy47Pech
Jdzfu04/wVEfKjQWdA+v+ZQdPh85k+EE/PoYryyPu/KEPgYXkud3xoymgvHoBl3B
CCwS4eoQTiVMMvte/ikX/EzzAGb2+ZCxqjYEwnwtCXUdw3V2CWlYD2MjiuFsivhB
rn8RHyu770wWRfzMzMIlcy93J9R99JJTHHaY3nRVVhWWhPp5DCWCS1Ic4xi4i8PE
/p6j+9ifm2jC7p+gsyTN3zdQAlJ0nUi5cloP2Q/167463LedSFBOij+edXwmyCyn
KUHKx/6jFdLd/0E12uSTXumQZ2GDivIyxifiE9Q51hGcMaBGR/9hYOgSBTYGEaE3
M2CPlvbJj7v9/lQUFKhBzXHi9B1x8qFQHsv+Lk2wbj7LNfMnhr0HPQ74zzxHK3gK
7W2euRM0ZYpXlBNBX1Ya+b6iKoSgFz2pOLgrOQeoya7aSpbNbjBXdQt5oBq69zPb
F71A+8JnSsG6nsqhAXrhSrRF0+77H9nom08fwg/IsbbpstALGarcDhsOazHPnLa4
+qmu3n8DpCetdRQAVjnetLCWtVTOu7d7GRLDlFFv8c2kXOKG43Dt4jOJy2sE1k2M
hc/4eqVTh/g6nFwxURbeGFGFSirr45FiR0AomuiIJFFXXQBQUcAd/2Z28U3o6Fst
1DKgRvA4hTMfCO9PPl7BClV6K8MC4HKNFOCL22QPDwEaT8omAMktK2aeetnr3PCK
l0uEutIYB/0tE5WwQT/tXIPDjmP/XFeW/Bmz9t0VktvfATKcLBFI/xLJUsGM7MfI
QWSd1KXS/UEnUsJdjqL5y3j4Ph+IC7x+mb3dXMifQxQ0MfL89SVcM941LU8qFUpz
oTYVAv8O2LavRrGesdhffsYNLdwzkHloQScAy/c2UB0otxueUyOnFRNPGzQGjzoJ
1FG1sFBFJ0oW6epRk5GDkWOkO401YmBkrNJYHeN2BtEvyZM+kMHJynIvoIzlH3Wt
8nAuxRWTQ0CO22sOFXMWTpD6XlqYL3D5ag1HJawXi24KjP+xzbeaA+2UBI2vJw8s
sj/p9GGVQ0tRdPvwygZNiGRZ+8kWj9x7rSYKmIeW56mJK0/61va36sBKIw2A6rQ9
0gumQPlhVjlZkqJ1DKz3+z6LEJi8bigo0Yz8+9/hH9dsKjo/rHQSWvWG2dzoQGDy
SUcl0+PO+2kHb31zr5zJkznE2ootQlc3JkqnfbkE/9F3otRsVufazsvwCjXCrHcV
KSDevgSzV8bMMi0eoKhO5uxuBUlJPRg9yNCE3T3iE4UaU7Hxy9Wm9JxWbyfA/NUb
++OLUByS23QHqNYbMn5ZvwsPa4C0IaouvMdx/mFmohaTJEEoaYrhr7v/hWh/jnlc
c/Y6bUubnHV0duk+JxVHtemc1NFOKKV75UfjfIGEDmAHqB6wbDk9M4f+rgHMN9SX
QIItMgO5D5UiWSSX1uMByElyiTgiw6kY+EB2E8gv24trH8Ycw4z6LtmyBztTcFFF
ayatizyv0FCXNtQyVshaFodawudhYp0PgtzV+xAY/6CcUdVjRpm38bqNa7peglMN
dWDxE/XZuazWE1/kAE4LZOyksPveLNrGlyamUdUHuQJz+FGnXTVpi3y06x4HMJDi
rFS4N2drKNArhJchfS3j9kRRxRmUHM1thFl8i9bmsGrX2STKPGWjXQgs5w3YTWKE
0TOyPN+S7+A/yEOi9wrMmVd+QL6414EJ9al/qYJkTG5O4v3fAx+KhE2e78UTKa5h
Fa1Gs+gU8MSiciIgFD5KfigFpdF1phGuHg5hduX7Hcgq37cATBwbh6eQKTz9A/lp
6kyNYl4kvfTS8SroKO22kUuYPmfWpJ5KNBLVJrS/zXh++JmyhNv5GV1DjCXfVF+i
HS0gaDMWkBmo3FzZb0Ts/3p5VnaoXOzYOnyyPfhJCyBQizQbyUa7nln99635qLbZ
2dvBvYKGQCh91AhhpITcKiTYD43iMvdxXcVAZA7iKYz/ARyQFinSArzYR/neYMYa
k5miaM6GqjXnRiDhrTFlvKuRhhN4WcAtQ6f0H+S4QnxZCxP+3cCha733PltnwFuI
cEogDPrqJSHDe0H6xcBOEEaf9JW3OFkq1SkhsGPqR0KX7d504nCPTMY7rFYVVQpd
rv/+mCBxtQ2X21tWPLfLxEi+W+PXnsUZ5eLIqOpeGBFGalzxZR5qx/wIBb6ZLAbP
7H9uRrX4lL12iAdLe5mg0KxjYVx9QUNaJG7WwyUVXByVYl3N2AJ+1WLtimUPJlhE
Y3VXCt0hsSrmN7zWCoxVWGRH0ioP6fWjCip4GSbiQ/ujlTgu2anzoGewVdonMzDk
jrUkC2qd1HhZa4D2+JVPqQ3VU63VFGQzAmEhhZNrAtmOtbM5g2rJsMqf9b3J8tZI
HwApPG0Z789lOJGO1SJKGR8X7CehxvzqQaSkP+xXlAG64vb1thpuJjEHBmzvCh8w
pfZ4eMWNtUTzkLxDfRxIRkxDkAOuUH7C/MMaqtghqvxNJoCOfyC+8C86UjuFi+lT
cygubbdUcfsiQ4GgpIwbmM0ar/b3LI6DdOWq0+rQ6VX0rFu0xgm8CvCywKYx+XJ/
cQ1p6j6AqHzGvMkhor5B+7OCtk5xHoeb1IA4u+ZJ9+jpfucvLDd8UF3N0IE5pibW
EdgFwqFYidXtrTPDQd0oW2+vxnDUCURnvcrQRgVz0XO0Uw6yWt3yKpGM3EPS2AW7
oG+hlxLkm/3A4cuftLjLccZazCiVQn057JDzdCx667TqhVbj1zH4EqiQQEjoi/mK
KIK0qEY/mR51bVQlJQ+oDfv3Gg7i5jimiqCq4DimYNFEsCZc1UyAtbcTs8kr2jK0
Kbk3uS6nela2mfaJtVeH4FKBy3Ml4P+BlPdJWQVU4l2E0D9cMG4vmFVTIcEyfU6e
xV+7KIoMkxQlKQXhBx9zJYqGLU+ax4Ned8VTwn2r4Q9LsrXPEoA2L8Bua1TxQd2O
g91DIw0DyPpIV8jyI5HYW8ps3xHtilxqfFu0w6Mb25M+KFu9snYUF7pzsmKmM+tV
/xWQw2hrL/uUN0NgkVpstQVuN0eGcm2R8IsXdrN7ovjkqFDenqYlP0YZc5HGF4Lj
4fzsFaMTjW8UFiyJyZYDb2CF9cgBvorxB+OtM87AueK2sFiT25QAU0hWUEPRt3BM
yvGCiCEHFadMnvcxp9ffo+I9s8M1xHX55ju5k77ztjPutx+wTZWirZwNkOR9jg4q
ywUnc14idQmY736XA0nVwhjNnGV2VuzImss1VaPrji9HAJKJzwCicRsMtPlSV4uX
8w9gQ5Q7W7vWIYqNfCJgyE8CdW2zlf1PNz9Y7UaxMrHI7HAcYPUOQtxs1E/N7BG+
nqTWxPX4dh6gQow38eepswJ4rY537bzIQBgc5lKciajC9bKmZSKVUnTl7wBUI5BQ
7gkHuH/Cr5+TvxWTSFQoB+HAQb3eY9WEZ8QXsn7vX6Ef3LXtXX5/kVGWpPkdppTU
isUB19sFBDPZGbAppR2mElobiMtefxA5R3MGtTALhl1GCJ9fKz0+JzZNaEvcgqtA
uIM0aBRQyCYhJvOBlKrLi4Py+GvoD5o46pom+Kyvl1v2UR+G7sMTT8Hr/aRlOL5d
5ylktq8nGQYgYgyyX0Vz+iYmicOH85sVqSOr7mQPKT5TbgQmSF19OYGr0y+/aEjh
UeSieSWZhcKQANCSfl31JmFjcAzEP+agVO0lGlu9vT9xRPXWjubpu7NroVLzLbOr
rWH/H6F4gaMkXgn8xpycPu68oczv41uwd76s1Bw/MASVteAbqsBF50gc9S83BkLB
qUOH0WBsLdmakq7gje7Mbh59EJMCpGZeVCGwzNx8bTKTGxKXRoStkj06wu+sn0hA
qzfLcVF3/Wbw5FErrE94FR6Fg3KSr6fuZy+kiTpPRXt15u9xfX/ji2qUxKUNI64+
bp8YR1SxGMDA/VwD3Z86wQ9RnOrx8UAb/433f9cHpwkx/tiTbuKxNuKPaZTfrnuj
sa13mhv2R/EaiskCgnT67Rggd2J3kK+Nn7zSxTGnPhmEaYdUVHXqLqI5qZEJaKSC
xQI3VmQaeQbBmv6E2/mKQuc2vtfhExXgx8LbTuGI32scw0U+cAaf+CU/nzw6Tkq6
ZqPGMC5OEuMjOg1rk/zarVcqJGrIZ+appZjiH829eZPEM2pTNJESTfr+knI7G66G
DXYXWORl33SeebStCgPmGCkesIreWis64/fCEYNA7Nm/zQ3YkpzyPZtI0sptMCEA
9kn+SuPLGHVHDlZNZ/1g/IOf8OzTXWs+FIrhiPd/Do48ZsRsZcnSEs1LCfPBGepT
OJ8x185vXaPqOGk46vifrR4PonxDuENEz888YdHFD+DNLRqxBHSjeQDidDXHAU7Q
YPTtse/i9g1cVr1/2zfDxG6ePjZGA0qt+WMukM21DWXY8k40Ag106HfJiFPnoM1P
0AnXWJf+jMnlpKCxlVeyCsCF09SivW6VdbiuflWK722nMFnbPVkgPR4NanD53kYw
CBQOOyRel2WaeTLwwnaQyBmF7ORrOF0Rsk7QOENv8G1e7e0iaB33I+XkD2qGJVZ1
qU9XV4RU+Y85842/yHRl8iayyXexD2MR9+sAxJQW8evTP2fcaxiCPWKsJENhPfb6
gMYFJ8/mJtMQPnVwuTdatl7KSh6YLDFEzOlIeL2zPqYkYIlzpiE+p/QV9N8cYrbE
Va+s9UZW4CfTf2yNEjHobX7wScFbGCWUoFxSNvPPDsZvNDvKTUtsPB1vqdC99qs4
g4wkjjHOQOWQq4wDxbYrDI5g4LCC8txh2OKAwywSHo4J+kgCsxxt6rk+PluZTLK9
hRvE8sRzsSLB6+orSyMcJlZDjsdXLoz//B0jN+N/1mGpbfQfUEc1lppShj83cgt5
ajaK/BmYsNaaFKOUW3ATFlVkFpM2IHzyiThSEBNl8x1s+JTrv0+tJA5Xeww2Ottq
aF/x+pLVLc3D8Ky+XkqL9Za6bkFG5oYoI/o6TDF4ge8C3dAH2jr73taRHafKvAdP
tz3NREEIpSnO5jZuG7wAyRbIsrEMkHmvVQEiViuZTJVooleyeiPTJkclTUfOQy9F
gl7tpPMEwNJJU0Mh1Se7/9EsoEjyqML/lacooM5hkoZr3ND/7F1jtJXo7WCT2oDq
S5Cg73VaZNcOFB9dh8vJMUVBbJp2aWlzS6RgbBhO0YcDL5GaQ4W5oP1sX57u4pyn
0A30xIrbPkkCeua8AJCxrdXj86CX2jCrvjgqweOd+x33fQDXzYDAghq0M0hLmOSq
hjF8qy8Shr2+CPO+9lOTa5s+co3urNqt2zObS13e/h8wdz84loVb1Yc90QOkK6IQ
HQoqS3FntTTbEghzG5EB3CYWfOtUzRHeAdUZ5PkVfOsUyvs5sdUsfmtyy0+fUhnj
NXAM3J5tQVSn3ZFLWD+cI8uSV10RSizpPR17C9zKkfr5uL+ORXhnPbUgTG9DFoa7
I4/Wa9YUSizLHIHnpo6Yv9znFeW5zbTF/bAko9RJClkdoH+NbSdz2M52yWyAx4jH
T5WTx9vo1zM1EZIRnKjUvcJACmRpq2q6HhHOSj/pJj4Qy32eX3zJbrqJcl+l5ZH9
Z/FK6Z5MEaDTxjnu1zidOtVS3SWiLUdPmFvetgD5UD9VRzRceeeaKAXDuWplXKR8
ecgX68lf15gi1Q1TNlugAO69RLmpwt9t/RhKOY8lCfQeHMrRN3qtLJmmeKDvbnJ6
uNJWGy/AofbypM542+bxsI49Q39UhfFDpuDYv18KwChiIciVBuoRev9iB8p/KxH6
uwXneAFNPlr/oQIwoupeB0cDtuqDRWV05e0NrY39YI0GdE4mIi9wsxDxkkmlggkk
MqKY50zDnalAmL9KeZ1jBJ51YsMDWDYpbdI18sM3z5zFHm6eTJwInVMBqGpv65MZ
SMMCaFivwvCUqKSsrPPc7CM6aEJk7uSiT5Pel88fAG5hpTF2ktsBF+ZgSdMMh9+o
t2f2AKi3hmSu8DPcCDDCwPkRKNIxV6UYCaSM9DUQCtXTas47Z6W8VszLRNahS4Tn
yP6dHek0/WYvYGpC4Ot9Lgdc++dMxFpQ6OG2bfllKJUZYXgOXR3fB853XEsHaHf7
zC6eBeJXlZi2PcS0fbK9VfzNZK5wRecnr7YN8Hbc3NyUZvfed3LgrMlpXAaVl8F3
nqUY4PyBhkbhIeBO6WBV02x9hym9rMx68T2ReIrBX1MClPWuYm/Spxnpi553qQaJ
x1cINAAETejZmNp9M8OMyJvtHY3s/Z8TsHKOjLy02HEvDp0dfI8Yh3H8lqKAuOF1
DSF2rb2RPObe8leNWQX/P0do8r0S7+FNX4Pm3mOFUvooeRJTxcZb8RZm/ug2uuDm
NxuqqcgbqCS/r+Ie/v6b7PnsMuyOw5LZX+1g8A+H77eCNjF7FbRmdEWuwIFWgW6e
amSRrsQjou4pUcjh9nvA2QEgv1SXTbTC3ffsdyLARxgnMZcqhhlpp8DRDAU6FFfi
GvrQdew56wHJgEy67T982tYq+BCL0QWIlqvRxXlppXvd0n5n8Q5gW6hYa8od+Zag
d/GOQPxhPmVKxDUVRxgFGF8dS9RmqB7Y+ua4sD20GXJks4774UPjS6ipExbLYK2N
nk3HYmWofBFLID18K3vyZiQZRVa0/Auw0KlpumrhuhsSGwNaGasVOh4RDtlOAC75
443AJOTbeyMHtsTsugx1P1p1H66MPojmUFk8aZc+P+1dCM8BKeneLT/RTMYQ77+N
UNo8VFvFTsP+0J87WbDEmlG4gIkuiQJ+5ATA18vV4E1D7uBn4x4YIK2qg+NA7DUL
WvBYFEQs4cerHCzYxSbyEjTjSYjgEZoPzlOWPPlmKNKmuf2Q5IlcBqBwir66Dadp
ZowpI2nTWYKR5Pz1sFblYxyXtNUke2VcpWpvLQouFH63STnBvncNLu7G6l/SNzy9
LiyqUY73PT6RgMHTAMLx/Y87BFd6VPFx4w5UHAytUlgog6rGJQrMFRbwqcRsTErs
l78zQ4hlzw68DSTUFMXFoub+R4p3Pp07nnG33raNzkNE14UY+72bhAcF7h8B8q+/
jYCYZZTmBml5Y5u22YQb+s+tRcsbiydJZ17BMOgMjI9W4ttonGUndGZuejsj926+
W+GUk7QdqK6vMmJB0VrooxeLKMGXkn0TVMF3T8/8z3T4guzgEMpZ9xGjlvDILOFg
eVQvnWlQ5Fuzyp7t8rsPhAHNKNLt0xpKtV9D/NCdqEVF+q731/iIzBRyEJmZBH/0
KyvbeUYcRDCayvIN+heoXAd5CrRzb4LTm1gjWrDM8I8zw/NjD32/y09Wgt9v/gdZ
YJ2HOZbLXaXACJkjlnZRGTKgGw10qQFYwEbB8RH6iryEShUR+qEugH3467Gjleog
PxhOwrwo/CVFvYXlGOg9gIHQNm20Ns2nMAv4YfdZYiOWl3TEKi6Ib+ZpvYoP+O+D
ExDtDaxqZKaxYwCoYEwKjgLrlyUvEzioM7VQX9o7XxKS/2t13sgYghejwYmzjETa
bT39cjrziWM0CKd1EQS487FHiW7v3mlHy7tf2Chz7KglTkeYW2qPEQxZnHl8WfvM
oKfazlde6a35UnmB4/oF8ga+1sii++s2APwhLDoBoqqcpTjh59WkSYQSMSwCI4DF
FhcTu8pT5Q08AE7Wc6jfU6Z5YLjPNq3MDd1f4xJkw32iOyRNaV9q5WvPglHiMxJq
A+VJj86q+GfDtP9Yl2KxiZt+PWTbLvBwVz/JcjNCCtO4IbHbV054qLc4GAdY95Cz
VqI2tQepGJxxLzvvN/0X/L7wnG96ofcmDE3z5bpu9HlnHUlmR5F+etK34Ig3LWi9
v3Sj1JAQalc6UOsesS+eKwLZorMwtX0Sq7NtHxf3+k1Bp5HBbIpWZAIdnBhkB3/G
sfiyOImUDNiyAzivL8Ejucp2bv7763NgBtgBiLVQUwe4hlmloUczxEbukNqR2HZe
o4AkM8vucv3R97jlu8OzyJpdNdCaX+lgOOB6tjSUWnTyxqf7ujYBCJdWB+F4IFkF
hH9mJ91fE81q7XzqFblzeq8mweTN4+aDBeeECxt5pyuR0VC0cPRuG+5U2E/Uwy5P
e8Yj+tkTxXThgCC4CG8txUDTuWBktsJNlbX/Mxigbb0iazM/24O/0ah0kqMLPavz
Gl/L4HGb1IDHzk2FaOL5rX+7mUUUjsvoammhpnrSsQ0U0xmYNkIWHquWyxQcdNcC
UbPyvG3KCkdplr4a1dtpLOU3gWz0mk7BO4B8xeOokjK69vtiNcPoInp3JVfZIEhs
aadsnlsr3uHq1rXwiHnlJhSkknppZVp4ot/hqmwG0uA5i3UbqfnxHt5LbVUtj/OK
U5m2tKbDytlmxut7K2ZqLCBRjOasobLCHd1YHzTOPgtXL1fGrSQctcnnaosDEP2S
tsDAirQjZiQ8Dgq04FCx2plsds5RgFa+8HC1jR82/JPZ6iDBGdEONkq/ZGNzjBNT
c0Qu2excziXUnWaNN8Zue6BzbkLQcwCmtI3vqOYxD/sepjLCEtmMTDNOo7ygaUT6
SSBxT2PEdIL4FsuSLULYj10NEPaBP/BzjjFR+Y/0GMmkbJUjoQcNlkVrMChxuQO7
4orCLhAa16M8rAZ4avG/7n4iiUa2YLYtNu7NNOXJskFhM3pIvYR7x91Gi9zBLLze
JZe3nOK2oBqg7pdBUiW1TA0uAsTMQ0YbRfwFcNw++KQTf03BDKJMAqJvUudgBQpM
AzrE2Niw8MiSE0pVR4SUO5cuAFY+HbU1ycZPWfjc/IlXC2r8TiajeNIAIWDA8fQA
aRcTJX7EofPPDrotqWD9I9khmrunrO4Cw9eTb8brHy6phkIfjUgPlylenjrGm1cm
7L4eHfKFkB3CB0yi8r8HW86luAI7icyQe0J47azunjT77x/VjOlSSMalColbvm5h
hQwsbqJcTG8p17rTzjfOLq8BIB2EOmOwHboW4xMRkV1vPMyatwrH6S3ajHdxZPUj
bjt05wN33U4g36MAZHsLjobBJcWUPDPGrF1PvWI/f/76dT7BdxKD10yPe4kC8pas
rlw/2iBd7sIq8A6/su8KMfTgO+E4Oxsqt6ED3vtUwFtZ8+20t25q/usTBK6GvDkI
G+hBZEQii6poG6NKU114B1GpS9U39aSbkjF9iea5j9ktmLpNqmeX/4pf+gZxZRnr
lRINneClfSI5M8+nn+cxclppgI6RjeK8N7UHciDoYMff/i1wLXyW7W3rY45nyc9k
5ukm1R0zrEXB4uWsCuZT8n64lCuTYZuUc5D+ouZt9zmIUsfJhekB34MlUcXW+7fT
b7PpuOmtSueDzxFH1NTM0VWR+i6RJWFIy4bN/v0wopBQ/qUUVKiAuC+uxi3N+DT8
LdSwPx5QXwAvcfOXTU87pakdgGHJQQxw1WAZ2cus02NCUAfgI8cnhk1whpfNIToM
JtJjjZWLAmKGJXXQrHps09ftoxyEsvUxOHoQ055LX3vT9NSi/3byA4GNirdGxlv4
pKlKMxATaTbiGWtrjrmqe0LIJKd92prmPg/BlF6Ru8/5v0C2W2MnEWkQCWZ5p9CS
hNgJiR0qXmvGrebqso9gMTjcHQC+8sg53oj7z5C581s7uCr1qNgCEiQLOEDcBfD1
kMcm30o2NxOy5LFP6117ZP31ae7Xhs6tXYPiiRTCTy8wZ1h0n/zwm+v9TjffebNr
hsLmj7MBk8PtO9Ez0NNA7dpXezQ4cCQPn/0zCQAlRgE105rdyGN6y/PLJX+By0j4
alDMiB1XHwSbLm9sLW+bSTct1PpGYKKymDrFZ29Y20fiUaZ89GZJvJYFKezCOJbH
ijfRaHXVejgzqLokabrFuwzMxqcoWQ55FoC98AqEuC5dOirh5EmdMdy+n/Nwio+q
ZnzPIcSmq1QY/UiaoTS/so5uItI0j92dvJZT1ZfrpiargWnRmvt8pBPlLLOwCxXq
5WEp3UCkYXs1xX5JmcVrBrNFtipvsxMUYmlzc2/aTlM3pQ/wZ0/JYk9txYI+F8XU
FA1jI+7kjlx5IRnQXRqzBKs3IY7YWiCSMwa1z8BCCK+Lv12YAgkrggI0eWii9gJb
wpm5u4XUyji3I/OZxOAekaE85nX3FW8xHUNEu5QQKxt8wDqhEeu2hDokXeennxR8
hoFVfhrMg+cE5juRjUKJL3oOlB9yPyzbbytjVLIK04v5tZsZ1860ahIbc6p0LEHf
qXoMvUSIHGEyunZnY/xe77vbgmOkL0lZVA6MVxyKOVToP4hr5Q/W2lC2R7ITb/Kw
olq3X62pf4jWarvok6zcAj5oQp7s9uQnV2nLWBWK+3JN2Jhp+FIvSwgJVYmKCqWj
Goo8gbJL2NvtuOXlPx0D7QgXsbw2NfNTPbsi0iVxhbNsfD466LkE/Ucx4jAeAjK9
1NGN4pDvOHdDrXfcK+L3W0xiS5FcfG7OVdiduA64DxaIMHGHl63VRVb+tKEU5W6D
GJHkbh0NLKD61J9+txnEt5BKeimlfACDn8DMv7iNR5PDiIiwxs4Q6Hr0ANjJjEmu
cFghMzkKHlJ6MFxD3mAVGELAL9+sBlmmgy682bWxePE8VpvdCPcqup2dX8OiC5eC
brOYNkHEF5JS6gJDobg7B45vi3Yjuy5OiOc95lVptmqMPoUEKaL19D9CHmEGfkho
tGd/ZWSJ67dFPQhBKIo7saMuwWrsg4HogIZVjq8oonYAxA1yo7Puq9m3QpHNu/ng
68HxKEKhf8BMfO94My05Iybbb1SdHhBAa5krQJRcgMrqPF5N4j12HPdK8yXPguwv
IwHLnDMkBbXkzXh1XtT8hGdOHeRHGiCg2lzJNYv1qQBWeyoO0Q3LKHeCV5j053sF
OAlbspRa1CRVYU3z+IiwbxsSZ0YUkJI2C5fVmQVan3fHgha9OHzxG2U0NVIZEj3Q
ZWsZAK4C9T4IWWN8HnQvZNwJxNNcxe15iTAhT23TknpmTVWYW9SNED/D05vZfJ8Y
yP6KRy5662z3f71azKDR3NmikN/R73HxXZOciljk33IwKR830dC5U4lo7cqVDEH8
ar8s6AF5weMzJ/whMT2eLwVjR1/KbdZGSFOJvaykuJv29jGl37q3e+w4vMYuPHHg
JroSOFgJiUnIuQ/Sl2BRRCjdSW6Kg+EWS6TrAKMcQEnbjTba9aUKQTqU9RsruhMV
DjT62RHNe4zbLQ4ENTAxC+x9kBi3x9jyngBP63ecuRlfMViB6dxhO+W4phFnMuW+
YFFSMkDrf/q1nPxiib3RB4iiWkEdNppoFDd8iZX+FMDYAFs/kSf5cWuT9lqvtMSy
USUS9te9peiA4lBZs2hLAq3sNf9RMBHH3Xpy2/1JZDiBqZNcYa8haEQgqmtYjhFf
AV6iJbJuSK9Cdx8fFLrXPVoZkFeFWFs4hqQlCVtUjwXMIyp3QP5DzsR4koZ34QC7
SHcVj0KDJgxJKYLs2dyRbWcso6xnAb2RayfxHmo8qZnMOrX6YI3nwaOlDZrhD6eI
S3eVNv2ANGjVbN5ic7nF0vaxHBNVJ+GecLguLER8KSqdn7mk2qghyNSyEn+RM2/e
B/SRJ3HY4ZazhiJ0YppHyr2QfrzVUExJtH6/rJRepMUXqZSpq8q/8M6dN4fSZhYZ
vXbBNgXPAb7mrlA0Lwy7kQ52hHuBiDpuEZ38V4zUFCaI7CQNNWiGp9jnAXwA5Tdq
6gXqS5Dz8Hog7r+Vg1fI7GklaLGVuho4axdRt8Wny9cJ2KcliT6LvulphD+CnHD8
KVDAtH6ixlWHvcMeAT2ho/ciauFbHxMGvXwW/w3ovqZ4EgO5NBptk/WYVeEKZOl1
yE6iOefvPCoHmMdEYHwLpCttk+oVHIQHAxZ7iIsG0MCeUH50pYEEU1CTIF6/0dN9
4QHPjvuTTlfdOaBt66dSivZtI8ClWjKBevY4cNmEmvpWboej54e/2AKY7BGdHbsD
CVvTJgLEUHdtS7QlqNXz/BfM8C8wu7+Nk77Wd8qu++ee0FdZG97p7n/QvCTVOZle
fuOo2eG4rp13RrXycTsCjA80k84y70NtqR17/5n7bcxjIYYtrebl+ta0W97TBdnp
7ymKa10M87lBSKa4Qmwrp71F8mMNvsj7t/vE69/ladudu/LCN87bJ5eMyT2XmqJj
40I7ynv050YlovwUbGV2O+XQCiJAaDWg5Oh5oPiZ9KOvhPzmRIesna0pfQyD1J1S
gF7eghQ7U4Kefm13wEmGooTkIWhVld9w2Bs937boy44L3mmt1Zykrn2oFwePvom3
4X86MjvSlA9hV/0GZnRBsAynvVIWSojUOwmb6tByYrlIGo9bAiJIE//P6zm659L/
lcj7uWHotjfX+7CyK4xdCp+AFINiYULzdHKS7wOJXZca3080g73NPEncmRLQnd/L
Vlq8QOSTASqsHxe47sZEYCiZZLC5cTwdwp33gu48d79z0pJH02kqAW97EQRpKn6L
q+PBvW59mnT4cp+N/E1TcKF9YKdDcTiV9IlilPgAsnLBhcBTEXnmnosRvO++9iXb
oFuJkb2sxCoe58g7Ye8gfJxCqcPJFDYzVhPvg6FxUGgf7Tx2r/gk4QL5CnVDjEvt
ywB9Olgl7qpase9aN8B/XMJRTfdAN5C7cObUUuitOzMo67Zx0oQeR5pVymjMSPJu
yVWKC3TCOM+Wa4gE7F3wgn3BxMV47MYkwj3a/d8lwTp83Haf1A5a0YLQHXfTmu3b
upwTnyO3pQbc3fgC79TlDr7hNdyG3noHNwIxxRVDWEXEMc3OVSFP7d3hF5nBQbO6
IrP5xZ9UWbYk4rsLrD4W8EeGETOdTPkxKb/B+gMuwCzSRcMQ+CzUtWKoH8FFOzx+
MM1xIkEZzBl+nLGm8GoTRylbjMDNvEorvUmzqHiqzKw1BWb230DHuaLkWAffh0wC
iIyGcrsHgOMa8RBEmV0/Wcwku2tQJWHZrPSZ/j9bMDR3Xl5isHSWZ9QH/0cO9qqt
zSz0DYc56wZ4Bl5g08Q7dAxDMvHvIG+RxW5CkUgzV756Xm1TjhlhqMKG2ODQx2Yf
G5ve0/P0K1HS6nyrhPsuB+NlCPh9x6lcFc0RjXpGB9EHUeK6rEtllN/pCxA7k1XJ
gSDospdQ1pFZRcYtA52aIinCzTgpwAHSUpo5YWkm1vyoxAkG3ax3/eSJU+ZVKj98
TL83s6ISVjKehOWoxwCysgtRQKoWGkmC+si9zWvyWbzCsygDka5c+TzH9H110iDO
2J/TZwfhy1BJZUFya5up59u5JU1SFpMX7vjpk5R2+Zd11EmTy/2rBbYWzUnShf3x
V4K5WD8XUYe4bfsSXC1pH5T+9cZzZjCeTGZ/B123F4ZxV5YwDVSfaSGeifzkyMGC
sym3B5dKolq26qSBEH0fBbCZ0ZNgOiG+rRi8MlxRcqR2lnlR+HhiVg0ucgwDUdg5
+Z7EVtiCY2ZQE676ihpBBx6ETjlO4GhaJZZ/k48vorISZE8EeVc3c8NdUqqjzFbT
JgpKNrEBFsnBrjU3RfKJ3P5ihQHUtVC8HarL74Olm+7NMU3FsFxzCOGGfCCz+A2G
vZYgzu62e59B197AHRxThO1CU3QukzZQzLvpZbGvFq4/hBLQr+6ybIPlzo4bInDp
fD6qC0wPk3BazUoyaBYiQTob4UCRdTvhBYlr64LxNi5LsAJcX9ktHbdSRcjFljqD
iOseOYwD5lg33eNJy+kkBrQeM5EOTFAzmCKilnz23VDSa+HUbFyuiGCPHuIC8Z7I
7EeqcI91EiGtbtw9Fluvdu08CNb03WINEpEDr7BNGzi6avIleagWmtn+K3cYfgmA
n92Hvbm2RAoS7Z7YOEd09zytulUbxX+5aurzaU8MWbfn0RZGGPdz7RuygxqU7BWc
vCwaj6IfEklFyV3GYfU3otmxTrv9FVvzvejJ4/9/3bFnNMkZzpCD/vE0Ihjor7zk
On06lURmF/VD1DJOJ/V6FaMGyVinmbLIJRGInSmttx/rTl0DNcdAdYjcF+QNpn5K
pZyrK0n47iWYOzeQ34/dWNS34p2ZLuCU61W0zxqR8FGrmvuwXNkBDuT5CMKoC6Zg
9bdmlTPF1YVOYYsoJISCxYjU7mAiR6ksQsEUnu6GlP3tGY/wAxlkW0OA6oxMUk9c
xoRoAJSZOkAlZBNIGyTkz4WmPHOP6bfGV0J7fXFWwNNUGAEDUYkrEqKYsKfETnnk
1qvYISr5GkTLDRdG73y++rcILl3cpcnhE1emiR4wqAQycXtVZZGaAsZKGVlxZPv6
2N5jp5KgRYMoEA+u8oES2z7l0DP+uXp3l4xmQoyDPVlFEMUpM0aWkIUOssiteXc5
HKSNayvKXvJC4yg3zpltn+8BSmFgs2OofCHIxOWgb8aE//sC6xbiRCrW2Wuwu+92
CTnODLjVKjj9JZz9wOtbwy6mzosioDEIFqNNRphx0tMYbv1cgAdQoKMmBujAp9Xn
nV15dIRx84j7j3cTNcMV9jJHD/pb5Wk/P5RTqq/4YeLF6qwZS2EZhGp4e/DnKngh
wBSTh3aI4nPN8jyFxo/fantuZid0NKfsBU8g4zc/loOYYEZ7S6v1eZxH3fE0rsT3
KBLmfgbzi0Oaiux+XHhhZMxFIorFEBVYFcka88NejIowhbzrmX0fTfAXPxi5W9Ln
oUxj1dY3OKBtCtnZcfZaBSVB8pnLcJ+//S9cdHaKgvo3smdAPERgaae8VZ5jCWgD
+2EewEWJYjHyX3lYNGuC0XEfKHshGC2Vr/RQmdnFva+X2q2iPQMCUkUhHrubIRaX
r9PelS22JiL7qZzuPFiV6rWG7iIbhFv5NjhOChU7VSPPWgr6jegwMcAaBthJkjTe
HgTsMaRgIRCigqgXed3OJv7SVjN2+gO9w8L5V+NReXV3dmIKTKyt4dZxYewXEh5E
DTRsHe4J5ny1T3fEPEhJn6tdL6Aj1VOr7lXpJtBpacU+bM0NnpBMeyomZ2WzO9wu
P3JR14P/baWGAFPLImjqlG5k7jTqnFrO58JB5+X03mMvH14uJf5NKK9YJusl/ZCP
75jurzdESdOYrQcWIsQXh6E8GXcy/+5Ighga3LlvZTTT5IYuplb0Fr+itcW4GkM4
dqd9/h6m92ylMoPGwDlvVWr59HMl13m7RIdj/ceKS+KIeGwhJDj7exUcrAR8A1J/
5kfp8Ny4gxGB2nRYlV+3t0voJEBzTP+2RaRx2LJIfcQL8jmeGcBzPVvGBcDL39df
kDJ7lpJeNH7eDGpLi0G31YL/BeA7YTdyrZRz71N9QXqucZuhqb/NVsXV9puGXrox
Su8fwxIZMZ7fBMNJc1th+x6tcD3/En4y58ybSMF6Mu0WsLhJKQOiok6ApDz3PHyM
bffdTZndfyYDYhR+B2iqA2smguWy+5YhnBnv12AIQSo5V/J3bTRL7YqjY0VCvPIh
lsLOW/Lru6UJzrZ+VJOQraSkPKZDZXaY17n43CO50J4CeYToXCvz89vEpxsLdOH7
S8DinalIULQBf0q7bAJ+bLxlHWqgDAzK+gHqeVvMXPLus1U1rsCMhv05uI7qvwms
IWsGYq08r9fCbPxrpAtVyImJtXLq5EgkMtZi1KIPjxlUXUfSKCkmIgJmWRcAfM01
Jwmz2nfN+WRqqLujzl1nXmSF9ozgwcsOYTXIzyMBuvCF42qso1qHBvql6udKMKVJ
GTEzo59+dgQ0ZAuIidECvONYq80zF/7hUK3GVnCjTlD+Y7QCPOBW0/nInpIJbI7e
dl9YY88yQh+Tws7GaisoyKG65bJjOjajuZqclCnjZpBAaGGvJTKE2cZXGHCDnMhU
ZLEMHgKRSi1WSdDXh7cY05vmXx9dTYNDo009ATeBwnL8pAh3Ys/mOxqTSuWu4ZCp
pe1FZmLlmku4Ne4d2PKeUEO4LWOIf8K/K7n6YZhSjULW4A5dG7q73aNGo0Nk9fN7
CEpKrLpuohkgwNJy5qRWpwYefJsBw0tvzmttHyG03TAE9J2kMx72+eXfksKTldwk
qClkHhzXCmpcMXjULsW2sSXbFPb8gsz+gHLVvDjaQEFAjAif6qUB5HKm/6ao6kZZ
m5o+i+glsio2rTxgG2GVJ+y2+JISCwXv6pCk2KTLKBMJY/Et4bsNe3hzvN+a2Cox
SpRDZ9fqxpI5gaWSk6j4prHlM3rlK1Q43WYIJq1N4biWAGB7WSN5pFwLkyyLu0tF
RF3icqq8SJ4324APNE8p+nZW1Z5dCb0NEpNuBVII2gyjxGJm7KMVU07t2OFz4SYo
rQfX2IKOmS9FXFsrKmopCZ0tGI8H0an3MXSybQG1Wju06L7GHB26PphZxPIG84qx
1RXQ2aaOiZhk1dZ6uRzQqVlL/kw2QHgLC/pmJoiDB9tMHmUznbh4PFua7cw4HJpS
e8VT1JqxOx9rW/ympgm0sDhTLLEpjdHjVxeX9+91QDgdUrO6ULC83aS0MuzLzEv0
V637LMp+GhfX0mA1BxbI+wdfVYGi/3VSZdrEKcGk2rZ4mmztoEo5nL4kRga+wHUY
eCqoASaPGiW4+oZ0qSkLJ9vStEbxcZ+CvX9DzHS2FbhN9z4x+l2/9dtXqRBO9Xxg
/aHMd2deWAYouBnatTPYoEIY5NOpQ7ymCdhRJKKkWVm5xVPY2Wsko/kHgEPF/5I1
ZLsmeMgErUZpxM0vnYE4UvvrlKbow/raYsBSv5sgCtvyMjHYG3XSMOASFv6Oxmtc
gPKuiafIMBzXX++/wpnI2d90tdDUISLEwsU7o5OnR1lAdmPV5i+sZAQPPJyndBkJ
gvpZQvALGUlBXKn06lOzOFz4s4jzAXJDA8L/OGxUSFCsEXMVxGiCNvgsLBlNL8ov
0fRey7wqObvB95y9NqRKU7g3a7fikBl1o8ffBScUktS7PKG7T9HZ9kbyyRz1ESco
3Kp3d7tiArhtPRzcVM16S7lgvVNiYKSqHXBIzYM0Ac5fwO4O+qNEpH/uV1XMK4Rs
/XYsiHgYOOAUb9jz6pk1stWdoWDJdoTumgNSc3F0lf7uYT+ddGdlt35EoEbG1TrU
Apasbtsb45uFVCFy4uu8NhwPy6EKTkB3eH+8eybtEoDMBLdJXlRskVI/ugY78D2Q
O6k9waybWckfERuOGyyt00FpmFpWa+mCKv+aKEF+3VJjOVQSgUl8jZUCHPZec4sr
6IViThhSivSjbFmrlLElz+7fhOPEhga8REZjBKwLhxL343CM5lCC14qsaaoYtjva
mPmw0sWhciCDhHgD9Phb1sOdpeZ3wAJn2gTpd4YPidyFbQLSaVPAR1HtY+JYCFed
vVXz4CvmYQ8W9pmaoov3aKCdD05MOdRo1dbcxeS86G3GSlTjXpuRhel565oW32gf
0H4BJj1/UhXcD6Cs4GrDtI/50OYZvu95s4zxeP7dZmGhIaObr624Rd6KMWEOwQVh
46Ht2Mix18Q3nMQNuh8T16FnWuD0wiU9E6TeamQuSumGN3MQo5Auk5DmX4SPyFUA
XMvvj4HlJc762Jzj40vvZIA8LTb32zSZvrLR3lpuOVxWiWbTXqUqiz+Oae6Q2yio
QitafvC3lg5517ZtkAtvrzJFj9h68zP3qmkjBjjmW3D8PaCZ8XtURfywZNXWgvz3
g03XqwA26kiqx2EFxIMINGBuiR2fH+yk16d6OyQtF4t66fK+yWlFdD9L0wUBK6Qe
3VhLSirI53t26aRkXDufOVd+wqI0vuAo9gwtlpwXLS79V2dnWUtIj1ywf7WTAt4o
ck8pWhCpFcjdiaKMjguPm0SPGQdD+TkEYBbssheT+zKVHkAWETK5F+Y5vSloNdmq
pGiuMMryK+ehl6eowhq7SZXsLh5KrQdcNUo3uUukXHjJyRVnBtkpKxYIAOkwSae+
HseDLpdEMnleTaRAPiq49+jCwSCSfgkKfUJPWNbyOOFompijkeAbMLl6gj5d89xD
zUMuFvU1O1Odq9Csde2bEtQ9MOlFWe+6OVqIezwL3QIUnU4ui86g3VBrvhV7ZVJ6
8G5XPghBwPSbJkzrZVCOtFjFDBVh++xtMpAf3Ukl/WcYT12DDNnkPexU0pg+iLml
Gb48Mi0Pd+BJSeRsugQFZwkAQcwn6sqn95A8++uN5SXnjRDpUS2XfMtK5eq2oTMO
KOXwfJgFN6sdP0Ar2kWAaBEfi+n7760/w9rzaJUrOqfNvPdWb+46GzSKbO8Sldg+
zFxeawa9UtvgOsP/PgW7guii3YgPiuCEC8r9Uf4IX+rGF9uSyhlYN/CUWdCJD8DL
fuk7omI0JADODYfo5wGRQe/MXFPltM8xikKQeuQlnD6JmGvROW07s39xUFb+KsLX
dCmQqPlBRHW/srHE1ICWJctGN34IFAZ3rGi8wEONGG3yM0PMBwbFYRuGIXGPQh9a
62RGEJVXeIDLM0XgPXeaxa/YOdje/X9nEZPteZdp9nd4FFdxoU849uuUmOaW1jaG
qGYZNNaatwM62QjJ5OL76ZbXDYeh9rrRIwrbEgHJ6PZHZDgcEJ+WpILj2GsI6QVC
1KT7BmZd7LDk/legTb1XWyp1Mkm8YQV5CmpBqDKHAguBa9AsIaM2NYRn8cmTSRSG
7jwhy899iMpr7i6NijFg1me32oeSxLpOUA9IgVqwDarfRXr9pyuq3Zt6u0hsmkqy
C8uzql2Uprh9prh28mCYBB9ixNU9pn3JgcQGrjN+lkv2ctzVGUKCxMJ8wib5TiMJ
dx6xw3g9smNk4a7PWRsovXa+0OCnDGt0cVu7f2ksYLhz1hA8hkXi1+PqgjugkXx9
b/eCjOWte/UVADvXY8C9/zCrkvUl7ATJCkBDEvFNsq1Wp3CRedqqnzofr7hN6aiD
Cfb5HD+i8vAxuV29pqzG8EOoap20V+4mKcJTZk9QzB2IE/GxnzPucyyCOTFE60W9
/XHoPMZdKIgCCLjGWb5G8Hkf+A2ia/XmygrT9rzrm1e0DH8rfjCiBdkE6qPBudaP
jmih+3t276IFWk5DRYdHl5OfqJQ73FbhY6iRBX5vyJbaQiPFxOK1mr70fJCcGW75
OlvBtO+ZYEKwy1leqMm2MUVFxzwXvShm8PdodeCWUMveNKbc8lFcLHp8stNK7eph
IapGH7P1eZxAXB2y1EIZvTfljr74HWKbuP7dUHypE7opLotZVXZThzAC1K8I1UM2
YtbcnledUxHFT2wuMDi/yRB/NgDvdKO0Wnlv0Z9ctAbPPXmnG7m3Ze2qJyo2TxSX
HQrzPNMQItoQCBBSAN8BaBL1g1OkxWNAZ8DNPix6Y4rTj2sic2nVVWoJgaveeZTe
H+B1paeAWe9GgJCghiAwIruaHD4g+Ok8z2zgguMhTbH57JnbYLPSbO/RFsN+drAC
CbeB9e3jXvy9+wqvDCdIUvpHAO4Erm2MX/eSFfNo+xE/QvoRZx+hfSQNLLMFcmhZ
b5nU4Tq6j0MIhUEs/b0yldHpIJBP4Fbaej5smtvt0fC8R2HT0LICFrncukWU3Vih
Ae9wHaXytmbLDeGZa9cdc47FSKFkQF4R1Q2Np2uSvaq0jhChyYFfwhEpMgs0w90r
A0YGACCBofg2bsCIhETmsOSCW6vTyTdHuW1zLO/i0mNl6DdeSo7WzR1OZTURW58Z
j4V6EMBHJhEA00BXUEDgxegikW3bSc+4HF4nzmxWDtxEzEU/rMGrOzYXXuWPDcE5
3Lv/xhgNZBRbzRCCu1qYf524TkwQuaqyjktO0YGyk/4dt6jfcwl5ZsECHtzMugZ6
aO2/mg65JNT/jLTvDvsj1JU3686zze/lptY6HnY5gGEdc5uLw2sNMOdLXKFshlNm
Ivs59oiUt/GLL/6RnE+tx6tEQVXbdqR+s6gEFhrBq4yCEliu2unaqzNTxqZQ+0yI
gy0cYJUygC89kW7u1SncfOElwyDUQKoAmY+3srw4Nx0x7UbT+BE1Myv0uj20nWvP
+89jXyToTYCvUHNlo6Q5brnTVdUnEjAjj8uUafEg/2sPEnLnqzMp9LfbGvwuBvW6
AaFurabhU2Zh9BuL4c3x5FsD5XdNw60eqdizjr3y4fAi8Fggp6K4d2Tz9OXa6ak0
1DqLRTuCTnU3D5JAK/Bkh+Vbp/pq0mRiLQlqy/yf94scIPtWSw7OU9kAmghReeNt
sKbiVOfNgZzc7EFM0GS1/To/Pow1+cg2k5N6VMtqpEgJ0oYR+Dby6iyvR3GqMLm4
takDm8PKHr3BSqCXgLll+95vinTRaXgVqiS1+SXQfzQbuGiAcBgiN0FRJSv2phgz
A7/isHOH+6vZ3Hm9cCM3LK3XuLdAmHd9+OwSaM4k91fjMN3H9ie3BhQAgUcH7OGs
Wxk3e6IIxU3DRGcVQUNn3SONR+r/qleN39iBhJIcEYrDPbQZeCQttvAsRntdOk/L
Mxis2WPcoVFCfSvpO8e5XvhoTM4r+ZVL4Zdv0WFVkA5m62ousk7v4K3Fg1cyFgyO
UqUpbwGrV2jybQTlYSHeyyPLhUC9NNSsa6dxVSqq9Ni0AzEaOqQgEq93PC3kGdsJ
JZCVcxpjaGMcxT7hwpcxnqDn6LBbfv0YI7gXaEE7i3ijlGVWDuwLNxan1OEJOw9Z
lers+vCoMuHdUUQt7O9zzp7uD1ZqzG+t8+adjJTu3nsElr5hAaAzwciGuIGlhuXX
j2w5ApaUlnLRebRhHQOkHkY/qffV30me8izih1uoabt33dKNU2fFeFNlGudEPuJc
AIrFGivSgJkbKVXX68nu7RIq2TldZM7GkBZnUHyKR7/mkLO9o56cxJeypDiuzWj4
w8ulsRb9AQ8FkJVAE7fCwvMaobZVCaoRKV23Z+Ymat6ybCxBnsFDwTBQbrwEaUZG
SEsfV/tzyQhsyWKD03hdALqGx6+fBh069Q3p+4Jjw3RAabk4WXOIMFi3OHUfbRYP
SJlyDPdbDdE/IkUwakiDdK6XEB+QKJL1/rj7SVkmPdQ4n3pGx8+jTkgxG4dHJ8JP
4neC4weB3MmPnyEV9QXTfZKMSM5WQOO/sNYDZJ5PpSOg+k5NY3iKfKPuHKnYWxFR
h8soCYQ6mDk2vKDgVoAlKpiuZoRp4k9rqo2iDwbkhIc/ISQHG9U+q7LMCoN1z8At
fK/eiqRBVEd2OLP3Ufpaghn7uDq8nYet3hbcXgBR6hLqX8okCBrlfE6yUGE5MN3D
72jbUqW2eg1hX02THVtiHR8aUQJ6kBK92gyrPgorY8mtJ5JgA0V/5fSODKU8N2KC
kYAs8Vm5xe4WzdbBhXVGCBGAPB9ANJvL6F4QxrVNP93G3DlfDILassmE0oN+GClt
PSRWDONFcOFe2HLE5NQjHU1hUlAXozJOH7Pu4yOTgBvUsfbDHS2T/6TTq9eNKBwa
qqz0tEMqrboBJOMUaDLCJnYmuUDalKYnVGyJt06tYld1NaKVVpxh6ut/5l0ersjM
Sgl4VE414h8N6EHe4syQ/WeZh97yZCmdJriETHTsJsv3lD/fs2I/Ei9erZf1au5C
n1Ra+oLvXRg7+82pNDhha9TdYZXL/NAjFSEyOCoqDOwfufi0flbXhjJb9sphmvuK
CYeRWpavGfLRlKvKqwCxAIxzw24k8p9LqXa6JxO+q42QHHXl9wV1IGqD5MlLOmuT
9v4KEXi2H10jytpArw7yH2jwcFZj1rlXFf2puu1iVKdWcq3tv7w9Mnb32iXc1JzW
p0bwoO+GnV9318vgXUUXCCHVf1KKRKboWukxOx7EC7wHMqjGCK94Y7XNfu2yfvTu
xn2PTZ1bzlFkVD16cHTUyTGVGvtepLZPy1WNOraljlCCQofrkmY2xsYc9B7WfsYe
zkeZaTmwwBKVXGSbO3QQVJ2pnMpUcCldwPxw5yZ0+uGR9hRwgxGv0nxr72a/DLD1
j/orrCjEtK/ev/ugmRl1uGJfcF0j/3zRNY9/oYcYI0oLJrcnvarVLRVP1tkcPcpH
E8P1jjdk7Xv6pgV014qJqtYOOvHYuRWxSA9MEw1e2Qe82go9XMoUx1slfzQ0lzGB
4Z41U3TSAP0jfZpXZuq7EyH4awl8jLzbF4ALoLshQOiZXJ4796xgbe+NuH1y0Dnd
SJiDubV3S3Uot7+ddFpTterUv1YEWv9wPcflVx6Jtmhy4uPXX6QvW93RTe4eKkSt
7PzX62FOH+BAmt4JrRwnpQKDtEQBVu3xhLqTiiP2kI1RRatS3U2Q79arguKwhqWZ
dIJUKZ39m1O5JY0lwrqAGXWiHg75DUI9ucdJNlkzjgSfMHcKSP9JsTZO+bSuv4Ae
qPdb9p3mkS7FqP2nsHJFRPR4oQU71Jh/OrhYuZXGWm/mT0uaXDcpLDu07/iI3X/3
zYN7JqH3a1di8hXR9pXTfB2ligpLL88SUVePs5rw6n/tHnOSN/8iGvWfbGKdbPm1
yOwcYsdEztFqLJWoYoE2aokYkK80EGhm9SJZmYuz9Y/jx9x3T+C5Wm4RlRBL2eCY
9VcQEExtB0Rdfme0g/SyRgcfTpZhHa1iIQMPhfAfWt1GFEKg3VSOrEmo6UULQobM
LIT0IZ5qy/twFuzOKjKpNWFAn7pqHpKUKwOV/RAgdFP4p5/S2phQOb/WGDbLGg9U
GUv2OTnezWg6f2jbARa3Kvu2PtFxoRj/+p2qWi8ii2fvP08flFw5rTJlaTd6sEod
nCe9I9B+u5XtRafWnsvC3r4g3d24/80irFFidp4oeaeyRQEr2o3bB9zeCMINTVmh
VuEICvuu0W+j7miU9uQyk6DgU52OqBeoaeCy9LYkQlmeIzzCW5LYdAkyjZ0eACd9
fATfPlHLQnhED51e1LayBT8CLQ5rUrfiJhU0dV9VPiUBqjBvZGZz5gOJYoJVJnDA
6F00Jlo+VftEUMu1LOkQYbDQze0jrBsAaY4JL/iwD8Dd+tP9NViurOGVmoOlXvfA
8hNUSdeE5Tw5MMsm75fkb0Xz8diaw9B7x0Urni5jenz/BJZTPwb6DtAUeITrCigi
OH04oLeBnE/ETTxGsDjXr6nOEEf+wXuSSNHCiNBJRz4JE/mSTDH0lvuV5CTO5aCW
otMAivtDyjdeecIH/KaaSoEOelH3plqerNsFuNnEYSO3i+m2IAjPqXuNdDEQsB2r
xJMhg9s9kWsiz9Ou/PGpOYxcVGUC+I1isHg1CynbU/szfmcBuyhJequsi8wSoAuW
YZP+ajFuXkHU5IfX6TEcHVsDdTGNI6a6fCiA0B09ipN5/bvZvnqgo+nzRtvCpKvi
NbKKnybJ4UGeG4FFuMithVxmvVAMhJNcMeJmPPSXeVitz8EQD98XyQspRSgkU3lG
Z3fZ5oR3umAdKPN2KkQRrI+KLcFALCBEFMh2M+b/Fqnupnw+77bgen8t4r4zAQET
Qi39z+JR/9kiBKU295jVTMBbG+8PgpjCUKLj+aZ3ij/WeCFwV1OaONT4/CSvm+X8
yV7yDzNIwHqn9DpYH0Y9FgVqmpgO2b9W/OG2bbL8qjtxk+SyX75WSdl7X6OeG7a1
n9Ld2h1lLOZZ5SlIdgLuafQZJVi5BBWkHwGS/NQQ7dclHcePF0OT5HyZCSfWdGPr
A8xY4IOsytXVr54QuwImGOXv5siShj0PO593DLqvmk/833RqoJzGham4RuNETWcQ
GztP22++tTepBcGlaSGfIgjuD9Voh55/GZMBdyk3emfE1k1LjAsy0lScq3DHremI
7Ik7qiGI9kluWlrC8qSC9vYasF9/545XOmXjPT5NApSmrM2scAxEoMHDL7p1Bcqd
/h++79jUsVDjr5JiA8XZltbwtuwk21j/ueucTAZgs/VtbE8q0nL1wLyI0Q4I+qzQ
9mdxUteT2VnTUwiR0622RjyI3BqAoKEnHsASm0obNcij6n2L/VO1BnSf/WljWu9o
AETB8WdWAFHvGxYST0iubw3ejCvTGVG1nvHuZ8wxaXKyyFAdz7Ek1jeHO/Ymtyj4
n8iR5x84Ee8aRaKiMyPb5IQDCM5w6suByG+LXRJ15W4hz4ZSfBOl+NiNZhI+/Su3
oAtkh6mkOlly0ckQvt6n8LbhnKu2PWDz16xCOfti787mam2VGy8BnKb4DPkCakkM
NL8zom/Sl5P1XVO5xfzayeexir/s9HX3OQ4wGjnlLGtwMvtYA2qf67zb+BThwlsF
LP+HUYRqfLxba03unEqKPD4aE0aF2SkQ/C0uSUWouf6dIsnJtGVm2rz75loY+V0v
ike+ZA6Jj7rl6JyDh7r4C0QzeStL87AVAP7JbsHQn3Oixdf3ili8FM85vvjQXmq8
5HQinsixdIBGKF1p4jQ44KPKGEMm+b7pTUXbDfdnNxPmQcViDBGEF/GleBy3BKci
s5A67Iwb3XgywksFSPnuSfGeHxYz6sErT0uJhMhM0+VYAp3g5yVPicXriA/i2AgN
gStJ5WlOzW0T7mTcRj4vfF2q8l2+bNIj48IOlX1K+GlwjroPsWIdrC7iIEFOE/3U
IjSI21MH8wVqtKssB9GUiM4hpBT5A0GxNjpZX3wpZmJvk/K8m8uWmlytSVOW59CY
oyTAs3/HSBrvIqZz44NhNZstv2zU8z13eZb6IDjjFpA6gF9Yd5gcXwqSQNH9KHgO
oUGBHXvL7yyhUynBxuf2ToWzSZXBzDDHWO/Sayve2iPx2ia2mtZ9jwqD3+78zzeb
oHSJNcoyJMawfZMYDACN0jXxEwvsJ/ZQL+3yZO4oNdBuK8aCg5ImEyNUepQE2IXu
XuVSM1tjWzYGrBZ1Df7pniWQp5Ahu1kz+fsJFgDY5V+lJLR/AtZT8vklJlm7Trwb
Ecj9a3siPbvLdADkr2b8vL3HowNmhN8a4RT2MyPw5a21B+dmPrRJZjnllxZm7Ryy
Lt4GhGfE0pDfSH/7sGHB9K/Mns/PJ2aHFyU6XBPpSTPbl/2MXtc0xCqEQMJpwH6y
svhlSR4FH6nr8VQO/DGJjw/JO9WfjCqdxfn18ZZi4Jy8o8KhGc4VRffysnehx752
OwMxqkSZnqtxVExoeci/dawoEc8vLhB7rl2sa9Xur/abD4+NIJjsTrGE3DGO7Y8O
lE4R+u/B3I+WKt+ddhfk3UaDhqyMiGePawRLr7VVWuAdx/hPzxupaJGC1Zj/K8kE
vueJ5zyRlU3OhDq6DMv22tBsv6wtRtgbCGTB9sDtWZUO7zXjHj7IWqH0eoN5IImY
eOVuQo6qiyJ9lbfsH0OSvQ/8Ys9qyCvo6t5D41chNJ201lKlJ72nvHfOfzvoHgba
91aOId0PyH9u9yS6NUBMTKko65ssuP9b9amsRUdLsE9+mdLJ06ZpMtML2z+IuAzg
P8KpjKyJ2ME8Ij+aCSgG90Kksw+vmaS1pu5Vb9S565CY3fkNASgBBycREP4/aWtM
SdEh5Hv/asqgsx+9fISPt66fwY88iIs9tIkX2CqvH6SuFMqgLl/CwXW3P285Btkd
I2xONS3q12RPHnX9hfWL18i10WKYA8D/0e+4rpXA82Cfjh3cSu+YWJlsN/v80nG0
rHxoy3jDlMFcK8Z5JlzjkoGY3cyTe2iw7DgquiO0ge+xMr2VWmvpQxDjc/WNgN0k
MAAXxknbTKWVJ7toxR3fRLxYY8T63zW3X07ULhg/y6Q+LgOfkKIzD0z2+zkpkIKx
W/e6X/ReOePhjOtOkaaVeVusKUc/Nni9EzNSz9xdRY3DbRmFcVXyi9knYCU/0Sx1
ZTec4if1gxmDqhPTkvKxRjnh8H01cVqpwtwHbJvnOm6VnyvQ7MqVS64YEcMTfh64
J426Wzm+aFlIHRSD4XYjr8ZnU0m/mEmw9xdZY9Uxsp65qHFalwu7P+D3KBG4oC8Z
Zc3SY07EsZYKon2GKKwhY8VdFB3ar3Xa4R8UvlBTxEwTnQ7RClav1XLtQr2y9PWj
kGRJGLjDTec5MXfXJogGwALim6hwIoBZ9x0Wb+5tue6KnAGcr5N/1OHnLCk0hTpX
pr7yw5UUl9QAO1LRYTJF5dXpprjlYzCLzoFnlbXwzTfqFtAkm2Tm1GMfnPKlx5DC
8/MbKDoCEw1bSED+Jd2ertggRXeUUC2b12SjP4PNTsaOCdMEj30ufwV8X/2Xdblz
6HFWCDLaIvu47gI1hlnVmYJHEcc2Wdqd0U9OoJA23hFViAunXd0DxZ2g0377BKAC
vF9Iaj4my+cwIdwgcqH6NTlWIZmdc/LH272WkMy1T9Po10NXZCmEneg25EjZus6D
vYoRA/zkP43/88moXb3Vx1WyBvlBjmReDl2rCVsduDpVYIxu04DGTUPZXMT9HNW6
sLDG6PzLdUTy9KPZKFw8EE0Wa16Qtjf8uyIaGTIKPApEPtkK4r2WBH/lf2xrSfbx
OpMluVGHZ5JNVATGmjMIAtarfzruC7krWwyOe6mINhj6wqMOF+eJdFNEP9a+r5np
ZJ46dfKDfNgDh39GFa+3IzfiGJCKjxACPwyTOF2V0f4gEQYc09eoGRfVTXDbTY1w
XeS3lp4oCZZHof4H4lwhR0oNnDi5NQz1JRpdTECz6szWRr6RhimoFy9g7EyfW9LV
ig7W+k+J/GzCwGE62M7qIIdmG842XF06oDvlS822Ozau5PIZ2sogk5D6CsMvk0eP
I0iFWAuMlttXYhbG0a7pPw/sBU+zQAJo7tiuFMk6waJPz9U2MCyOr3IiFG6+uaXj
e5yIOr4qpgU58JnYblddp679Dxgv0bt1dvtWpE+8va5ItkxD3o0toUmz77veLsq1
Ku25NOo/i9q16L5CDu/PqFEEPXfz1zh77lCFFJR8B/Ft1s+M0dNZ+eU4hbzjUFdC
C3jSiirUqePZAZnEXJ8NBrmpLcI+FSFehN8IBWTsElOIqDg+a11xhdjy/yfjE9m6
NnPh+yTm4mriOX97n+tkMaQqm+5vh7nJJFSNQ4fbSKbKGvduR4spNAURcPxqE+KU
AQgEg+/86MjQjxIOZ9zPSCF2WiCD1hgBd4tLHlECnyyxvCigFKlD/ZJXbK2g2QFt
TCyBVWSohoAKLPlMFNBNPkcN7IzV9d7255JUx4bhLCA59uUmukR05MbnVLn4KOo8
RvsX+QZboThwXP0U5opYw//Vvc8pwtyvrGuC4IXs7qk0k0uKwj/MHoZEtyC772iU
BRL2tOruDcr/DOo//SuEFlVX79Tnzw9VpGyA9OpgwouKwuxnxU/zHhP4ceYJUixh
HV52CKqtIjGPPEgmbDYrwqqQs7j/UfmfmgKDhyM65c6IAlsZCUGgmx7YAFNWg4Or
fhwRbXeUSdoTeivEoxMiUrcfcaJ0N0E62g30z8DxCLRKOk4zHILOKrSkqwmS9zKN
CxkOtbfCd3D+fDRGhoBNWFMkPzw6XUd0g3w/UJdkzsF/SsuVAn0nTK8rNuC2w33r
kj6dJBWELZrMYfGPI1PXyZBBlMMYw8WtQ7ejw2F7w4kxU4CoL6r69mslN5x1iprx
0q+E3Ejj04og4Ex/xtvWHOEQbN8IH6WevPiZ+M1DdPg0wbN9g5J6akSS+Q98lPuq
iWFKirMSIHJSJfQNHrFZTmvj/y3ckZhjVKPnmyKrCoBaIEvOwIDOdZmA9fL9HlGA
/reJJn1/P+LYjbwG77H7IFv8Lz31g586+w4JWJyB9P3eaUcMV0yk8wGBxTrAxb08
x6W4DqVUREk+0gJ8ksdTghs7DFkle2WUA/DJ9qUqVT09iWg8mOPpxQ78C9F7LZ25
VRQ2kdpzTgKOspwzLUCNuRC5QqfB6Z9Qf8PGNFQm0zNddnMdvxsatzBn1y+fYNJ0
hBdaA4cnG5Z1mEAIRapWpvFQWVkb1zXSpkDTG2hJidrqlHtNzslqA7yey257hWby
tsFZd5fhlizPCjXmFy0LR+vYLz0tE4MFYo+qcL0hKTJUHuNXKF1jLPh8iNVx9jup
954wr07TJduQsosXpnJKV/nl7IyE0NpKHWlMcy/5t5yHm+tjetVQP+6/fjekZaKe
92Y6Zq+ebCZSwfRMchj1uEJQ26iBE5lV64p3h6u27e8eX+5eLaetVYqZEenar72b
vaPzfUucjrJOrg9tA2sRBnwv84EkQU4rLH1ld5NKzkiOIlJUlFDKuAlaviVbOigZ
Vgv5adl6Z2vTn6MolWKcaXjWEi0sxV4PvFcXtDPRIHEZ/rfhidZLG8qreiDh3k42
cDU05UOhpNQSSkwlFVp09P5xi4bmjsR+TmzOgcPijR0T3VAfB/kT0tmHE4v4KMOz
tJh3+SB18ckFnCWspqE03ex25jFbrqEYMgAYmVhssu3w734FCFEy4Qlay8Rr0rF+
VqpotVKajAfwOHGD6tZG2s/9QVo/k/gOPUCSRJGcGVPJ4AeSH5c0KuOVjaaVgplC
R+3QisRdDNjtiqzjtm7f/V107mm6bzY/pOttnF9WbvPBcTzokybVnjngN0oEWtuU
zgehUHNEKGrLQ/KvcPvTtDSwJtBB+txBoOsHm1MQioRmFUFq8/HdAEZ7WC99Hvik
SJd/186zBex2XyXK97CvwTwrDqVRR/9OMuxpkF8Kj2+EisIsK0JemEkcK/H4b1+n
U+be5IQz9MBlfJJyxteSzaevvh6H8eNv9r/o8cQUK8Ro2CiP3DZw6coxXWJqimYS
F/yOCR8A97mLfg9V9QZtXtRzgiQSpNQJY3cZIt+WFRgr8MVn2QvakNDunNMDNMlr
1Gw/B8UmOw2TdjVEpvan1XIWnivi2JxRDiFkwsYUDhwwb/WOKahk30jo7euarLEo
WWnSNG7sPb1mmHrNuJxmFB9p7V0dlrKMG6UM5mfMaY3Yoemdiwh8x7fkcD1ioyro
T7DZOih//Q4GOwFmXxNyFYl3ZkdP/SyIXFuiA/WzZ9tLe8HgUHbHCeXIvA2k50Dh
h5HfNuYmXIEH1MTKBDLrdNepqlBkjRbIdVQFvlh6DqQlUrFyuO975d22SKLwrtU+
9qZ1dFRhKu1J9CnNIOqmyxiLbZVVCSBRfrWcYoduOgn76dNz0vYmzZa17yGJjEgA
PjuhQppkKLNTAL1+JdPwjuzwE4Q4tc7BpW6kDa2mHpIMPKxjhSJuPk1NKiam9TIE
X2Z2Fo2104e4iYYTeyZ6V00DdOYBwkfVUTbB2X1017mvO6b425fyqoqnBCfSQCcn
p7bWOvBWTO7LrRET8TAvqbx6upZUmcbCzEwwgkBjls99Hw2ine/lJMjFksWcNJki
n2i6rhTEvmslyH13WCp0QE5fS5p4mPSwoUpcjz5MbWI1FDHKTWCzQ/Jig3IAQRTQ
0wwnnkezYdjOJbX7JQ5zl+ThfOTPsrGQMNeIhA7DRg6s4GQ7N7w2SBjRbuUHsY8P
sXc5j/7CdFvX9QaRgfzvk/ch9XLY/aLIt+O94gHz5mTsJ1TCN0dGHDXbRkln3+BW
SykgzlI6RhoijUM+mzpHE/EXVpbnS0mIe8DYCoPCoArZALvbQQ1aJeoJRLD3YUZJ
vzqa+anSgL0Vph6i2n7E//55Ho7GOUi59bllOnE6C9cnZpK93oEggxztJF2wRHA5
wSQB9xFtbPOyJWr9A5jPXoYGJJFnaqnJma6RKNJ5i0Bf7RuvyxeX0oeek3q7p2oH
SA1ri4qNc1dM7e90MHODE/5md+rcIGbOHuMCAwDRJ9RoO2BifINpfJ8Y/M7MVx/1
Vf80xrLTJSqTgpNcBMQUAYlMuH1LTAq7DQBtLr18uYfKjcEAg7l4zvG0SbN5p+Bv
rUSEk3ZSWlSM3KxCqa3D4tt3I4ZatgwcyKvTm8fjZY90SoXjaISGdmwF4RNFVUO3
xwT1BsXS1F5gLuVAxyK2s2ngNvcdDraBNheEYTmoqtsxqkEVCT5Z0fG19qkva9UR
tUKhO4DJyX8Vlvh6zwpxO2U++Wr2unXO4VVFJxn+6ofNy6iUzdX9atNJX/fu4KOq
FdtbStL1Si8gjEsHrjhHodcXgdq10eZ8cAfAUwYKMAYugpoRIoUNMjJowjMRaJy5
nxBkxqKNGj0q6czIuMWhyfDWS+0DWDrrZqumyhKZg9P2qrhcNJ8Wi/rlI8qagSUv
xdNn8UuJgpGmMxK2S+NId7H4lbVlvg9GuqJ/5RlJM739+wcGoeIo4pZHrilMljpq
M23MzM1v5BvT+Tz1b+yJMquHQT4EmcaytbVORz74zKQ71jzxGtxnezTom4W5Or9r
sfQigfn8KEmGkBLizRYzVtJNBap/zQInq8vNv+HDdIMzFW/rrwRlhYjlvbfNBhCz
KMFkJcXalNSW4c7gsumhu6sZ4vQgZ44JcN3VZr2VJjK6kiX1RUc163cmY6KLQw+c
WRp86maQqB493eQSf3afVqB+BOGvvxGOdIfk0WpnjHx9qWjTH0GIuipivk9PvVTg
qLaNOg8eVYC4QopPbLmjkxuT+4QhvJqZzSYH5b/XDM5AgsM2GqFlhmyRbQ+G2QzL
fl8fwP/oueuX9VZhWZ7cXzeYmgPpvpLoY99dPR7S2M9bclzDIzKQZXe6ja0Bqu1i
htPDqhHv2ljqzzshgho5FgPmgc4pUABAqObexqZyLDxfoBG/+hqo6SMkE0pObLvv
vrls7pGsoFxQwUNq1HNPOIzYTBR3C23bPdHfjPaUDqDPxB8J3b0/0yI4XsRzQ/JI
hrf8uu1z3RfaEq07ebX9AXBdQFq8IBBNMyb+AO0X2O6R9Gd6rtSfk4MSGZzcyRJt
tzD37MRd1iGGVHhWuNJkYv514jkMejQIybUlW3fIz1DcCl7Bgo9WpusZGKXBlcDh
+MVAFq4zpxYPpsMxF+nG33HGBKgGtYJr9FQAwePN3vIeMhl2aelsgaNSqjlaUQFG
nhZjXTkWvYujCT2+lnobBUWCbgizcbXQ0C/QdmZgDqBiOC9bJ+bmaTzIwlmmqoPd
YSL7MJOfGLVKPMw/1Nh3vbvQTVGzY/OsTc7RmgVsiT8siOzhR1zQTmENnKSoN1Hm
ew9bmdMYYrV8dhhMSlqWO/l6HY6xvq1LmhRC7IfoUNQVLHvQwfCWJr2HXxtCWEsj
DlJ9Lss8ZGnGSUeGW9VYZ9kBa4JUwbPRzu9jPGTUz8orX5rERP/wiXgWwiqMDdr1
KieBLRplhi6AKkujQgfjm8cl3KinShYCAVhWEpSrFXVYRg9gTWHgjd3slaTssjNo
XqInfRS6oA+a1uq7ZnsdT1f95lnytdh2YV4sCN1prY9X612DvqAdi+uFrOVnmr6u
M3csR1Ya9ZJrKQYZkep4DIVYZTkYgV7m8vegjeqly6TuYP/2keFr4H5glGXpclCU
LRY7pBNocM+jkoEl2JoWQ8Ch9KOmo650TYBJXBdhJ4x/h64PcYYrgqfNiIlpX7kI
hyLZJ5Kv7ow4g2WZtVURDM5okyFvOLT2ZXNS8DllMzx0oXnKQalJAzgXwI7wCV1W
SvT/a+rtuO5lCLbgyVwJASZ8rUSwQiVAdrfp50yfFThIVChcVFbfvR5HQq/Ph+bl
hWFIOT/aZ5nd/81ObAPR0POMyCs0bXNnYZkAV4LRCynFkrnZElQQqnE6tTfW92xy
Z8jIrhnAdb5pAg34ywq74nbBhMAmGWM5ptJ+aBxHQbE9RxGjqGVL8R62ddFXgnhw
1rKg5y4Ma7p1wKBDDc10IeL+9CWu08fn4FNRHt/bBmnoBt2AMjDC4+4IBlCl7Hfw
mrqbo4kHQoBMkDLNzMvaG91cRhrbkFypbUQHxVtTJzBVjLqh3XfuV7dtC514SIK1
D5AYt8g3MJAZqCSN+IYuJLOiG/pnMEtrMyk6PYAe0CuhHGl6C2IMG/HjEMDN6XkQ
vlr0Avp9RKQuvqUITLxHBza4WaEZ1p6z4G/K5iPX9xUDm0L95ykSlN+yeS5iB0Ck
9XP6Tfj1mMKSMGjN/YORW8XUX04qdsdnMeIMxVgaF0pkT7BqUCjrPBI7wT7FCSuM
7DCbn/oTc2W4Cs577UCgI+j8c4K6O8F3/PVsJJ9b0jf+1bOmhMkZgccJliuFoXBy
ibfGiG5iy5P9jmK9zE4QTIA+SoVIiYzeYEBau5a0xCLnlIk9rLqOmD+jC2pfRVUk
ntc+mjpAe7P/x//6OBikTzEXE24ZjyqsBeVeQbwHfBZ6w9GP0Nay9hPd/wONcbf5
HdlUKt1M2JXehMvWVECs7njV9YHUKGVVKmQ0vy6wj/owwby7i5ttXo8yRW4QaFsG
zJLUHYGQ8YWZUz9JEWJ2K39Uqvhvq8Gcl0m2PQNeGZTUeWefFtubWlFctdPggLrq
kUn4Qui0vr+vGDI5wJAM3FrbYKv4++Ntf5vVy1zoMcaKH9ISRfRwtSfJ+2GULEh0
vm/TiPjpLSYTSq2hjPhIUxeFIBKsFc39xh0xepNFZYYnLpKSHVOmMypPsgrBI6Rm
LSrgTnzBcYXeigjIKl+NkNQD9LClz3G1gICTZEkRWeGjH4svPc6KB3spWHcJPIGt
WXYoQVo84B0GF9hM3GHO6Y09fUpRN+JOfQDPoESs3kYC4s8mBNlTfDzg7moo6+Gi
PnuAcXs9uv3VphQgAEE1+ezIL+VT/6B4RTrYy/lufDRuI8a4ulb4pGy6BGelzwdG
kaIoeJBbOpxxkR1qnj5hmLpMhuS8pfFJHn+GKGxg3A2XvOWHMK64D5AcI5n74mxo
RFWdonWYLNLCcw1SWtq/zydhpROR74qnZwfHVVNgL+OTBRre6LhjOvr5dJvm1VPG
gPFHa+sKbjdr62HWJgdf5USHSzsYdIJZhe7vsRajQeHA5t1nJp1TyFP+Tg6sflhs
WqKpTSBu9YX6v3T4wUib3rY4dIOoVBsXW+nIB4DT4+lkuCyQn55y92bIb/iHNdNL
rHzkBfEIVvkYwn8UAR5f21NRvga9k9AJhyRb0gRDLjTSpQUzWOMd0UscES6E4HeU
rRgRBulP1bRQE+e8eIwDeP4LL+b6vCN8dwMOvJeVwtOuaykY9nayjqzyFpehMlOt
C9WhKjtYdfz5GKhjJmuAwH2pPxRe/lTSSctRPNn9NHajV48ajEkcj1uuFd+0XiJm
x3bY/qlMFUZW47xNiVHth1LzRFroH4iojBoxl2uFlcewoEtvFz350KAml8t/47m8
PijWxutO3VilI3UaNmxwNfBxUUr9igY1wpXI6QkPIDANGwlCMxxCLAfM2Y4yFipd
56mQCxVW+UUIMAz+hdtSiqy60UAysceqS5g9IMPd1idWyTtU+XffHUOCpAvRpbi1
jTS5kneMcKfNqpIHXxDOOpKcK2+Fxc2fcjsRDrQdIodJ4XzfO0+qDUe4KsWTtl0Y
pXeMRFxtCEOjPSLFK9wAdi/ogDAPkoh2nSb+L6vGFNvtylziwlZA8/vKnraYe20W
cXpRRI3oqzhnaPVj6ESCTASAwbHfktbhN4nhOC+JVZ6KrMNvALNuOOfX9Kme4IYU
19F3qZ8konz3DTgNziYpKuLOYAn5Bo2WTIARLaD+7gbVuAt+g0bak4hV3me+Ftrr
yW8nkdQhiaSS95R9Ls869WYnv34UILlFuHRI8aa3OnaWAZCmKoHQGyUBC34wtN1u
nZyuEkLnsbVBV7cDk0BjBt1Z7Qm5amJ7jcaGPo9hzwd7/44UBvlegUWV0CJDmZF3
WvB0HRrBhH45256lOWulapv8CMgAydI/C6q0syaCOCgvfwYuyPcAWMP2CoI0QryV
eUchrrqK4LSduPdZP3DGfaH7g6Q13PCqN9fLeSp0qw1huQUCzGYY0aH0FoVIhg+i
6VDeush+zw+c6biuWmpjFtt2YO296ExJts46oy5LXOk94v2HwAVh7cNMGyKTNYIq
hFT4P7ujrEo0IUsOm6+uATy3+Qynfl8niHyKz4e9TgcHiKfZ+6d0f4wbEvLapqGZ
M5LsbtLvxnS9p+mhkhRxDi6rMthHry6jE2pCZ5F4SA2FK6D1ShAy5EhU6s2lK2cT
hA2Bkq/xTEyHTJGekpmoshiV+OwB8qq6pH7UfZk7lYkfRcGSaM0tmBQT5ZU/avqj
Fnjj1uiM2N+05B+auC3Rqkx8x4omQrsa2vklZGJJBBocu45Dx/TU5GMEt1uiy66m
LMDJbY8Jceq3ALT7zn809Jq48yh2MpPVx7YWJVJwNiPVU3T5f8cJ8kAw0NDG5zVl
6aOsEqD2J6rbyNlAn21o/+n9UsKHrI6+vMvAy/ZQPW6gByIkfGQ4YAACDUuszK+S
bVoYGjTuG0VxsFyqPeITJrxAMcljfLOxR1H/GgZQgRzZuG6xx7IW3iZfi895vMeq
SsMNikyk9ryLREBWxTucB7gmkdrCyte04fiitE0xsR/h7V2Ha8saWhfbOZ7BxRvm
dT/K8uadF+WdUFPfxbtIWNj9i3jZ5+XyM8440zrx8wO2wXoi6DRdtOFFWtNgKhsW
/ddN3tHXHIVncSAFwm2+8fsGodhagOWQ2azFyRlI1O3kbIr/3FLLZkOpmvhecMut
QRlwclyNIfz6IIt2RCmlB22gA9dSNhtS5IkeIYVAjOF3P082WpW7xbDx3BT7dFwW
FYh7b02AzWBURMdyULdKQ7sXBv/tUYl0ZnuabQZ+4bJ5mYd7dEi8ybB1rTm4a1TC
uTvRr3bfEACChOx77eEiIHE+BqqbtIzCKdy9s1RP83PGjiI9n9sDfeilH5gbP5fa
U3JpkS2+0Zm0xMCGOIMY9Cnho0ZSFDihYmQW4cgPh9NmG5jiww53a/UpzM6WYkvQ
/uF6mwZaoT8LjkFA1e+lJTuR82Upyaa5db/OOsO4z1yu42WD8hC5ESdSwJaHrh6F
aIo/KT4VhuZpxhZgFJYru8+Fq5odnhQgsO+3ExSQRfU2Nxhe/zuxZW5xRLBrWTlp
amC+t4AnLkQT14doO5+lPKeAwbHQ5ABHjLqWex0HFYErGgyp4exz2G4x2226IUL2
pQ93GHinMmuIroFRKzECwPlvf/SWkdzpq+i6eZ+ZJswAZC0/tIrjHfg3LGuoFkJq
HwiV2J1h3oFW+Hq5aXZNBEMi8qaKlmKwW+TLtaUWFmO90B/RsnyGO++pJWJWSJLA
ueaXAQMVjYvuenLSma4fgnaHvPh//x81+8UUBBpLmfAOon9IU6M4m9wSLFp8hctx
vXwc+0W7krynMcxIXFJEUVwvENOAdPlE+tHCWajdhodAeepeR+9WC8K49hTRj4LY
rO9R/b2Birw82/vUENu8UPNkqoqf6YUKe/QznvacDunkLrRQsttIe8fyMBqYeds/
+I2hEa+ahyjgELg08q3zQyuA1HLuasthBAQqBs8978c0ro13Ls7eDz7Ta2YizxXW
cjPW9haBtbmLL0LH5JafqNcZZutl+K3iKqlTc9a31emoLtD77HimHawiGNj11su6
Z80kKE0x94jA0Mst2RjjJoXQgXBGTqY8iuiKu6On4/nbKRCrnDkKoljGQuG2cajJ
pW1Ekgv/BkMDfJuLsWdOrOyJbZvJ1koFaA17b1K4q0y7s5e3N6gIPuRapRjFAYqz
uGdMswMlEiyYUPGBl3vhyj6wc+QnX2RnonyyRgDT2WmcC/vepKg92KrYVmYlxL+X
MQZAAjqAVDDQf0l6wMxSJI7JVSzp9VmYzFRWNKvz63gK4z8ROVWvBXtkVCrfuOK7
g11/Bx9KAasxL5h/3KYnF3CduuQnQE9UI4EgOBAUlnXHqh8G5QKInIvsB/ebSnzV
rBBt9ZcEtUn/c+Z9lUkdXzOZnAXVuOc8l8p5YdgJjgARiLpD1kiHdBVjENTY3qVP
s5K+VFLjaZqVYJWqm0se0zDC8a2rtFwODyYcjaSAcv98mpfaBL7DajpC8klPrwr8
han8fDHJETwm7zFxKcOCXk4Gl12xdjfT45n0ZqW63oHOM7rPtEf7JQGrpuxoP9f/
Gv7KnwGs70KQ4d0EQ8+kMqtG3A2bdTXOsrgddOgBimMKD3Dl+nSuRTek9ADZonVN
SjlKKGltmVo0wChEQ8ypf8fOUG65qTZ4Igfkjl8gPoTP2yFpDT6/oJsZXAsiiyc6
nqz4lwjLlEaDqFxWQV5WHuYnlqiPSA+X+Ax5ePhHQYfwZg8fy++ON1X7tdeBUCcn
5t4bPI1f7S2YEYuPTc+dLA+Z6CdyLUSbZfF9ThQrD73Tn9BhCJrpLEuVqaFQY2nG
uDhMsF1or4RBElejdN7o05jGoDPJbWzAE64BMd+Pwh+anhOh7LtiKCe+7x9/Eaf1
9vcHexB9tW4emkHhQ2RXlZqRv3W8MPLxMsNg8uRZDMJzec+9qKKsIPk/2FFWX5RA
/zLNX2etZOrN8zPVP65Z/RmCE/DjHhkQwGMRWFFipSBhLT0EhOLwhoz8RFt0ElF8
IqT0kdg8X9QvKZAXLPW2TK+FJPAMoGwOWNsDi3ipZwDg66cmE42jsYG0N7XoG2O7
UQm3bjLrDkcrJubW8Az1khlmAVLunmw9VfLQzMR86wfvJyNaq9a+PLFQor/xLuqn
gxMgSt+RbrDZAkHYQWjwClcoovaAQHB361AmDE4vkVy9Mbktt+0sADTMGNHmoAVl
iFtwIj8wGX+0OuaZP2SyCru3gSDHVvWYPEQHMAD7vdh8jbrrCuciSJr1OnLGr1UD
hLuKKFBBJDYBW4VAtgnu6hovXXxbcIHOj0TGrsywgxeR+9l/MPHwmd15iRhQpo1Z
ArjyhwzWXqXSHy9lmH/du41RVLF4xbQZhVLM3sREZ8Z1XAmybZ9M2oXSAyj4N4z2
awS4VPeny0A7xR3bVwbtYJaXiUe7E9tNYRQKzjc85bZANfaWqyHrhTTJyMPXOnfj
qPT//wGnJBM1pa5XXNzULWoBdtutXY0VwOg0Dt1LsNqoo6cL+k+Kuj9dEDn/eKMA
aTDrK6+GNpV5BcDd+w8ndfhxyV7H9o7vpKyPPWiflLY0oslUGObjo4i/x/fzlNAb
R8PZKM+eY7zBK8qzHRNa7s7sV1/HjIIa5PskYvD/MOyq/sJ00/irSmOnCHU946Ca
Vz5OU9mNqwRP3XLB1tP6s0AtzTBscMCWFTVeLqpO2ue+hvFlucG9esn3yqKb8QRY
tbxBKHICI171b0H0N+47WErn11B4gnDfTht3/G3X6dXjYxIbiLnqZKjObAAJ65Qm
WzVWNxVTUGTZueBlVaIycLuyVDs2Oy/gHJvdxFcP028yOF6/UIuE5yUATkAJQCzZ
WfDk0Ol11ZmXIb55gnjx2hN91PPgq1sXXvoe+NL7w18b4buN9UNAHWa+9gPoi6cP
CPpxex1rjHd2s0tBvNnI6ChuK/P20Akh4/x1+ZSKVZlSztkcL1QwKOT06vy/oQ+H
C+3Rpana9SI/WFZONANciDy4GJS+T5Bjclsp5tq/WRHcSF+ebeaerln6MVJbW7T/
LdTxqat/zphl/o5H0UhxnrCo7iZEQHB00Ve8tX3zp9XnkbsBcdJeYH20RH0ZGL+t
fFgRCTGNW707pZ4dMd+LuWFphG/JS9Ch8OYCAjzP3hXyFzzzBXAqOiPdRxquscA0
1LKvJXn3P8DPGHAeR4UQTn0raGHp2PPcyqxsT2FdciApPl4of88d4ov6m0GZmgDp
yKXhRccarTchGFQxusROqDuWhO1T30MFMiWDlRGnuFbek8y5eh+6dzWlrYMEUeJj
uocTQv9gTMSJYlOjySeOs7in2+ulpEFvFWhMy8DsbsMeUO97JR9Gr8uRnxMYIk57
HIuenyu6HQAUUP/xZEa+43TlDA6X9znqhI4n+/0qdB32ZUq0A8/OE4+w3nSY0Vsc
BZypUZeKwGzbEXs3j/WEGQ39Be1pKyPRVHY7GU+569OCmkYudqAr5R2LsSKkhYBI
ZG9eHEHy+xNxGzNuUZO1jA8mrWqW817rIdOCWMJzhZUuI2P15qAhy1h1xDvd9k6w
GEIXzx8Xo9L24zzbpHGHYqEmXqIweSEi8uJw0bAwk2t7aRY+CWiO8FKflbFTbkpI
adClr1HV1IYrQBom3LOITmPQa8WkheSw/QcDGRDPRrZ0Xhjh4TBVIBSQL0Ic2D6a
/Gqqtpua9rHVWPWcWfMwITp94g0q5/BxMQKF4d2xhLj07nyfcHbrNaU+LX92hK98
wUK6Q23i8/XjtKHj0UnXL7+aZ1BobM3FfjE/JFT3diZtHUtozGyEr6DBM2hyp6/2
VSv/nqgQVssalbx/9Msu1B0i23iWdi4qiQia4PkHCFkNQJ2QLw/h4LZnvmF9/qAX
HBBl6xgdNCUQOlzlcUV5L1otKPQl0OdLAwOJ720vQEwwJbsxkn4foDy9Lw1PK0aC
phq78ioN+wbIAkGckisrnoS/WvuYxZSFNf1CwAleHz58i3ce4DlPBGXtcG53j0xs
O320Qovo/YSrHaeV8GAKKf9bLlPDJl0L1k2wRvjRiPRGowM0zMVnwiT2kwRrlBsa
4bOu1Hau2nQiLzOLspdB5D0nkKwsZKHNg3wTAImgDLGO/etnwKBJZry6A4ZFywvr
Hpk54t/sW4OrnwS6bhyfV3XUmssaDnRLKvE2YMd/1u3U0h+B+hlvabsJveCBHcJo
xQE2+jgzapSRIdoIbHMI1QzRL+VY0aqAnfEb2KnbgTAhtbzMrwx029hdGHFeUp7K
+8siZ4s6eWUlu7YAaH+8mUC5t1/aHkm3/6tktNwXRqmiIbXYIVg6SwVl4PYVyXEm
I3lu9aoYw2mZEkTuPLm24SnEZJeDXeCTeCAC8MctvdZF0i8MUdG9F0oG7AEdhfyl
ViH2PUW5T0/WHHxB9qA2eT/yfonX5hdXiRVZGahd0GqC120INWlKZ/P3FZXW6AzL
F9nGysd4hDqh+Rg2dvT4GdBZ/AWT63L8LKwhMyVy+FhwJhB73dXL9ETp4IsbvR9Q
Dc/Pc4uEI+gDU+e9U+3Zqrkn88gjSqrDAZvWsArSEG34gEXxFqyhhB2BZjK9DCvg
kbnxIIjILE/aDqzhl9PGgdbhP1XHhYl85PM14pGY4jFQGQvEjVusy1EoWAdFOZLc
Jljpq28LaoZbpgUz2rBhX1P3Qv7idzt+DxnYdf6KJBGYnJslJvVqGoFd1YXwvDKG
sMYtFAeu/En3WZJhITnAJWYBP+WNJvpKsY4SK+g1pXCPYyahXCIA5iskl8QD69RV
TLvEiqW+6ThO1jSFqCzOnyCTTzMwr1WT7vjmSNGNEDHyWdKzPLnszPdhclOeJHZg
/WB2vsaXigmW7AeNy/EE3fyVNWMovczQ6Vq+DwfQ17cuzJZZ6vKyH2LCAPLTRw79
1BBCOS6t13Pep+8ikkGy7wyYZ9nvxYtYcUnSm9b0AFALk8P6Fhv5DKwePebrIXTj
aa9zKBp54ETWAK+j9wRLyCzM5T0bYHfJME82xOsZfc542pVCYn5com0rmiVfYk1d
EZAzsky0pHoqEBBHfAGPw+Jdc5Qzp+YCxJzl03kMWZ9rWto44yEfOtZtTSnI1oUQ
fEfC1910DXvl2l3GhF/bX/TUzJQqYtIUeiKkX3qQ3NeuWTHqNfv2ai+gOxiHD3G3
9ayTLTwwa/qxAyJ/VG6yTZ2hWfZ4qDUIdPh69Y8ad5hAhG9Zehb6BSGcjU/xy5VV
9mN9QM9Q8JNirV3AsItO4cUyIVCNysuKAJ+hTeOUUVhMQ55TihWdQgCh31+bmLzr
c8DMpmRU0lbpNG9FZIkHxEhWICWXc6WlYnrMcICFDWLA6kLvEX4bdZDfSSmVFsD7
vA2qOPCsTfvFdgOpKr58IS8yklukg7k1j9jnjvqHv8kSK6rqqfQqMKnkcQb0UzOq
fZO+nYhv60eRJLTj+qmICJjoofR9MBSaIxc3y1BJ+WVirlqmVkf8XiARhFUpnK3x
lKBVo2moT7YqBA5G3BtcqFiSh4Dk1AOBhT5oBjMr5bkeNfevd76TWiUSIY05VTuU
MXW/bnkR/v2re7FZ5Xj4OCNpehfP2CUYMvZJI7DyoUZvyKWDvKfCrwkHEQGm5Puo
irMmIBPKDjjGKXni5G9vopp937Z8bBjHS3EFjQLMpNyMAUWzoPPaxdl2LmU4xXoC
sHS41ZFSaB8C91aU6zfe6vf0kA1pKAmRAk2XwEVctDcnnF5X1rN2x3y/zoyXOHCO
F2UMLQkJit2aY+IiWPblxUg051hMXJdYhdXmEWG0PQxWWbuUCvf4IVOyvAU0ttNw
EA78xeGeTiODc2hPUCUKFA7a38owO8mlQUmuwnUMNEPmMfL46vX3gLkWjm6rbDaN
pV4FEsscqkwQTFDf9WZ4B/WMQWbRLXqpkZZGnfmO1q1vam3VA5yZIY6biO8jsJAf
VmZEaGVhxBW7lhbY0Me9TtnW8yOKyJOF1Ol0mMuDENePrAGu+riiMzHbHfYa5Lpe
5dUh0NmRdVosvcAcGnEtEmOR169L2Czu4klvRV/1IzOCbiUMsrunhfnaLn0hq94y
ZSjfkClTOkKRbSDBlXcHyt7fm/htU+c9MVYpNyaYgUo4t/7qxFDcb7x01XSxc04j
KDb2wJooKQ+x2gkGBLZnegwP/GvZSuuP6p1s4i5wawO2blzzeX3UL+4hwLCL7Ll1
unFfJvOlgRMabIZfoe8Qbv96tNtMMYtBQPovjgJBF3O4niILyU5tULCl37/0P3+0
ptdBuhgXBbSQcQuTgGd3Zw2fU3g7KdDRc7AorZnJAVqlRMNufOtR3hVIRqHLnSxe
iwUTe8iiEGNejQk6jUQOWVbGcoAvk7oC9dmL5D0VAw7mK2tk1FUZQa21ZgVpDWOt
SrqCdOKW8XtlxQarCuxKWSTEKvAFum0uPyNjWrGrvPakZpspIaZ6p9vLQk3GTcOs
uKW5xCeImug/Q6XgPYUudZhV6DY83oqb0v58doPeFY1sNYvcPV2P0Q9SMpAfi9MX
98oYv3oXfN6o0UdL4YzWN7msFP68WTJpmKBcpI5dzwF6HdcXH4iWZAP5ZLIlBGZ7
E1qunqnjyNQmyAeDxAyH3A4xIHabEOK15N5OOz8dspSCvcumNaFK43CHHyzp9d7f
rF8iHObopM010UAwapLohIf0Rar7cjvlKioo72BnTdc9zTIj7Ra050JFfZ0cCEm0
slUPcjNcVdlLA85V/hsEcEsFMOA2qw7K1gAqm/JLnitgANLG51DYwe4FoJn4gWYj
e5aohKq1DCSHkSFRV1q8BhtNQq/ixmKWqB07L+58992tSsMSHtfAqxiR+7reA521
+rgkH9v5+a5pkf04L00GCOx3Ui0hq3/4+CtmL8jFMoXKmVk4EStg6w4aiTi8h/Xf
Ky5gaLnQMeuayHiAOvR1yKnvRncLFWDu2YrQAaC270OOnlFRcrQZeN4lOvjK3rOH
rBZ7h2iIIhp/27gEZoKrMAYy1s5IvXQrX7JP1719NMS3xJVB8efJh6aJPOrgKNqP
RdnuwVJS6FGtU9ZlPKm+DXr8LJkZ63kJ/AXu/h1rZPtsl3Cc0+jrGhApPLvdHt4K
79e6qfYHKJfrx/j7067w5xvLACa7RCGk6/7YZSAzj+CqjRrXQt+vCLVpXEfgBIVZ
QNs7LE5XpZn8azdurAi+IYZ4zdGnr/REeTQt6+3b1B0J3CgxsOT0tIcffYuMbT7p
f2lalupt/FpCsHe0pkPxVB9s+THxzU/7y4WzRspzK6nIHLCpqXvIMZvyci6g010O
2220lMT18l8J5OBj/rBmvTWps4Mn+SHvxgd+ziklyMVErDzBULGg2OuT75ktYOpP
1CQA6UY1tJH/LZ7wwsWIXGZalbT1nTUKmHCc0/acrr6OjkDpxjFvLu+N8AWq1OEl
Dx/IcBkJTTTaIPMvT3oUFKQts4Pzh+4F4+Qf75mZg6lzW00+JlK7HrCRgJ/7NZPM
s5lJ5qBlPAHhQko9Bn4Q7f8hS3PPLIrtRSeGPkyzVNjZ+djm3sNcS9uCL00HVfbZ
4gI1gPDoWfyt3UrZZ1AkDgZUKNjztAuhGXKNgoABh/c8f1MZVoKTrThEtcchTpZG
z1CEgadNZ5lbJaJ8I/eJvn3GGMCgOfwhMVa+qvEj8zqZStf7yACyf1NjRaqn40fD
DKsEw3Qd5cgU18M28ZTpihGQNI7tJECGRN9bbNB19pZdIySLhf9bOiIKez9uEIuW
YiGPO/aomDWnA5cZwm86AdctyAcMLQuuni8Cw2TsubkTCpEeVCUW4jJiz2RfzRvD
J0uf9Bdt/H9NJPa7Kd35V78Kr3I9FCDQxujctVxLKk1+XHHpiNKKdksGxiHcCQtZ
atgJKM4YLeijqTmVomObmL07PQ6BqzXQIISid4EhlSRiakuRMK9SDkI4a+xXImWJ
TXnZDsQ3ibWDGmvQv3WI8BICdxZYeMOSlKk58yblI7pVhZZG/jsiCy2GRu2CG+PC
jzXzBvZoxsRY+7pPDle8oMLHSD5TZnt9tzhMlD+3wL2SlYTdi1Fl2QVtSGcK+Uf1
sJhuaEYjDTwk/sGi2+76pxGwl0U2Cg5ZavtHAvyu5G4CS9Ta6eN73e6IqZypbeha
WQORaL4egGi6Ewe+SBhlZ7sg6EQT7Ji3AYWUqHys/mPTOrM+p7Tfv0EdbKGgRGNO
CKAKz8KtrGSZkkSEr6oNcbS8yNj31m1/6tBQ10rLpNTFunOezJ3Zbf6ChyHjV0cb
9vA8YldeiAK2J3oMfJG74G4Sv+1oY9WvtUrKQqCliWC7MEzePTJEoaCxffuhA/uQ
jjKG7PWMXmyEw2ExwcOXGV7C8ys+EreaVS0ycaPHk7hvJrdYgxXJG5La2uz9Cb6l
0M9eVt9c9Y0iIJ7X+OS3fMbdb7PrY4Hy3uGhcT+KSwZoT2jbCYf4dwuW4gnGZaos
9v+UGZFrhjyJ5nrdEOJKCjw/I9YEMFxObnA6lLolJnsBA6Fy9mf0PdRm5n6ZlZ/2
Qn+9cB3zDzICAAHRNZa2rkxh0JFAZkQRRf7LYgXGiqZchWn/Cf6bV9SPBXp7yJf+
mDy77V0qYPbJ+54FZaTJKktHz3kxKigLFGtbSSZRWaPFFSm1FHn2sutSh4d6apjf
yuuPSWZ0KjPOS/DFt87sMARd1TmJOOXByopaWF9cNHkyhXyHMxn7xhBIH7QREC54
WZ2avHM5yLU+OLGvytVPrRulsJspSjGhJipHhEAYXBhnoztSt2BDZ1Rc6B8+wyLn
x+7EFlvJNlCDkKKX0lsA4AK2T/yoabYIg76GlKP6kxzQPC1b6j1blwtqUzjujqbt
NDOE4l2Qu/9pCtij9sRZRYNymHpHCuwzBam3I+UWiibeIaAap6Wd93nn999NaM/P
kyo2oOcjGmjC3oIg2LhtU0we62z3IZ2cK5T2cGIKz/o0tfjZ/LTVqn2Jgy64svlR
QMKglEd4J2Jj56A4us/OV64/CRLftnV2o4B8VOAUXTu0B+OdHdACgQOjivPfsepj
KuljcCiqma+7iRMKITgtq4bnBu66ppCjUWoHdYHm6pTNFs8411jGIs5tcTIur+SN
DLoZrMap7Kj2xPh8lMZCyJIdkJapIR3ebIVEtFVaBpyTRS/177LcxjaPADoJjcw4
TqIrkI9wt0wI7yG1tkS/VKdEgDvUygGWQ+8OU3e0WMXgMHZ59htsu3DCphwhrtp+
iLHzndZ5mBZmnBPGtbdMBHovtmIXvf1BdGCKPIyNtC7hBQgnUmFOU/8DuKcGKIyW
kevSqYnNGiHNjVXIMFQPxHrvXBLHMKhQ81yAoAP31HdQECS970OKgBJxyUBa7gCe
p3LWkydlGFZRNsFDSSRZZrJ8GuPBALxIY+DviZ1U+1KQHq7z2sB85GkqLqAJ1CUS
5BePsxVRFjdhF21NR5Z3lWV0zbe0HTS/9UxJS634Nyp2kuEL9TRL8MNByFXvc/2M
thnFAt0ZfgMrXes6yWfzHIXy0dwjF8+oRvMeoG1MJc8mp80CBqUxC5HWouZaBCyZ
2UZpFXY/Ws3qVaF9WPpGEMmkQDtdwNgyI0JmxJJpEAsjYZqupbajdqu4jEn5odCy
54E0MDl+jiWX/lNspjecnjpqOFkPw3+CiOVhkLa/jVMsE52HQhgShwy0f7pwYLF+
/BIG8wSg11dg5XVqKjlo+jZboez1UBxsVsuqAh5hMkFzYOHWdZPDHJ/aojS6Otf3
75qd9ksYwMuwcgY4XKl54xaAnOUPHwGUWBJPkkEI/L837zRF+Je3Pbo7X1EscPeN
QVnEnvE5St9+Sa4kY9hkrks6XFmI1c8E/fJqLNwwQqgcn6QSEn66tirdgUuru4+j
+l4Xc8ZK6LttvVQ085kLXVX+4ptapMCuYJGXiXuKVTUD4zAFJtW8edQUexAh5N5c
GEJK5BqXyjw/OpW0ozRR2NaVCvfZnq0iETa960Pv358zghAVjxS3/s39nZt/ZHON
u6buZxbqzLGxcOl9PvdkSPCnbWI82fnc6ZoDx7H1fjLfRPLCCDr35l5GgHOzRWdE
aPcfAS6+Z/nN3zAWp3clh9Tx1Dx+u6pHsZzK3FL9i2t50TDUyiUhz14dfVgKZt9U
u0G18Btze+K2gPNlP6LF8yQVhzuV557c/T3gzSladrtv+yHb+VDV2C1+qqzLDgRV
GBdgBq30tyManjMvtKH7UZGfg5W/+EgE7TljZI3NJVjKazWeCjCCUK0VChQs4gQP
iumKw1vCSpBsoQUOhhAoanAt/siPkDuJg1k51wia2FbjIp2xZJaq/jTozETb1Lfn
oGfUEjDPR+h7L6dIy9JXwXmuVghDSRC4W8f7NW7kIE6gYADG7cVY4Wlas/l0jdBt
zCkqAVbn4t6HH2PDnWahSjzDys5QBOiuwIfq0chD1Yhf4bXAz1JQoZ1Q1bIznR1f
Ei0zGwSK25ClpSocqi2LsLCrBihz8z4KO763xvgndw9shpsns5E1b4HoqoI9+Kja
ILOjZ7iiAfJ9bEt1n/DbXSPy5no5WV74k33uD37TtnyMSY5eh3tCRzWo3iIBByfE
60jJHKwoXsLgPPdu+jX4f+hAyj7zTw8iSSx7a278aYbKDj46kaMUf/ehW0YknTq6
rdagotvthscEJLZuX1Qv/BJ6mLBsACsKjVG4Q9VP5ccrOikR5Icf6O44kWtuKXLx
sdbRBKaBCQO9qAw0TnfMpMBwiQNlZjmMDwurx0OrVCE0iv8OXIwJ0VdnwlXBIX2Q
OJ9PhoecDOMSBvTzAD5zt9+Xm3R8pTWFjqh5O6ND/wWgIRC3aAjOUyarvJSNSc4I
JhVnoYctrZ77INTfI9MGa6LBhYNlwA+HANGTEVh9Ww/ZBtZHwen7zrFX3PmhPEMn
MbD9DvPqPXSIprORO340893i/shqu2vrCoa9vzmoOM2tuyrFfosn3X4d3PJ46RQT
rb/2qDXZr8R8yGK9+p816C/MOe/4L44UPKmuPjJo+P3UyvEAgaT6WueBmYXoB7Kj
QM3VPgkeXsMcwXEi7u9owSgqmY8A68HDlRDo2Yxxj1cPus1VgG8Fnqb2ZIUyue2v
9AePu5liWQ+UQBrUAkN4p9Ykig1wMyL6DLx+1niomZ/tJS8OZN6AMy8Z3xvnQ/bo
TeKroKm4P86ArkXqDWK+R1o1h/WqBQ5fjSd2YtSBIYFu7LJvb0mEP+/bfZca3s3v
C2vRWZv3OAmMGuT8t6/aybm9BkWBVFu1p7TChARd6Cuppe53BSZc/Oyzr7pbKevx
Ozgop82uuGV+d/UYQVt2RIgt7ivE7g1wZRzYooAkRtiAwIFBAulfqMd1G0YMIebL
iJjzhf+az6dEJCIUVOoLaAxNM9czup7FGoxj0L4zWIwgWsGm4z6igZAp/TV/PtNW
4gt8lGmteGlCdSa1f8xOKMGjTd15beeiMVPcvXRJTAoPH8pQrT4qVkh1VsIcebkz
jAdqYT8Mlec7no7g8PBEul5UK3NeDk2jkVMpC823o5M2Vvt+qrDicI0O5U5lqgEA
CmUCkYhKlPloItRhVpRZzJCNlECupxl+FZi8PAi5mSt0a/vd5E8v8ppdvuEP8wre
fMAcRr14ypaK//BohSQOVJfpqmWmaBp7VtL4W9b2brX7EMHDqYnmI9tPR0X8xjSP
DE74LE9xod257DdIB1Sxt0K74W/5mbpux+dT7OdT/1KKACOoLbrMv6DS32va54fc
7KK4CGJDdVunDcaDJ41pBdwzEHHZfWf2nMe28HrqTrnY88QLwUH0buSEVuTsipoL
9XZAA6rIA+SgXyDg7OWRZgWz8uNFNwyNiz+gSC4y39BB8su26i+PmtBqm+tdsRkv
0G2B5krHhr3eCsYGNLEuEirOrzxm/3lR9tAzObFzxrsojlZWuriTGVgr4l6Hnbzh
6aCH+RMETjipzbV8qoEtrOpjR3kCcq8XH7hiZFxHY6eqMDn7IwWab/UWpNG5wRix
UGh8fYgFY3OkYLxRBaXNPn25DjI7S3CjwqhZy2aBxMm4K+pPJZyIBH9ZUVOGiYp0
xn5HJ1RIvb6nhKor6IrXhWWY+e9+wMD3ZxTk50d1dlWFi3vQH4tqQErsOp/zEizG
hecx2Ah5qSH6n5SNLg00BFlSlTmmK075rxiDEUCQ6405h+thFtJsocFJ02iC3MSK
5U7CsZmU2+3cANayauH44qG5Ta3lBXfWsJ6uRaiDyRo2H1B432BjuvZhyaXwbjg4
iwGA63y9TXkY+37Mg0crnW9yCxqi5m7DBNX7PN4PdBGMXQKIo3IKTU21xRAILEJ2
9QVN5am5bPKMo5VGjzh6ei/CjNk7ID1iw8JS8uQiciJguUMW0kW8CYjM879BAJi5
J17eu5RqmzkA2Im0iiGEg8D4NUucpMeK46mNeb5U3Ph6fAhbx/a0/9q9w1y1U9JZ
ltMlooYZmIEbb0OkK3rjjADRdzyxG3/i/dCg0xllzd3iheBSPU0aTcX7oNcWAxVK
HclhNU9kcV4y+AR7SWSmFT5XcIYbSauXfqf8I4RolmdfwuKLaOevMwAjjpRJU/VX
S9Fv4pi3uABmSbhQ3qZ3xaMkQDd46/xPAMaLxgN4Ko0uX5IgDaFcAUypl4Ja85zl
yoku9SXqCUoRy5RSqYEfWF3ZfOP8Un3y8BWL8Pb8cjtct1qYeZXKBaLTnWHCt3V5
0OUS4B4tDLmm5T41e9tbbq8ZpPGm+gYaIdQkIAb6v1Dn2t1otN6rYBbKogT6gDYb
JjBGuXZlWTviTexF+UP5T93pN4BnGf1fVDHz0QwwXCcb9gqv57+9vnLhjpnQ0juf
V7Dn4yYjccBvAbFapQSXAS61JemI9LYyxapw1FH6m6jsfnhnaoDTsIiT85R3NKra
/qf9WDvNSOLFaqcGpWBFGtJGQvoKPID4FzD5bAhDEQUcCUTvWHfxfAHNii/erfjg
heoUj/iXflc+p0BX3P+sQpsE/iJiKTUzMwYzutzJRz1Z2Kma/Shv92uEU4dlFgyz
mAfAYE5uCl/DXN16urKEYpeuqrrlm5DSUXmdplkbyw9SFLGypx89mneFDnY1HcDt
fb5JQ7F1Dzw457U5Nl9CKMe2tvE6d4R4mtjF55AsMkrmdvkvn58R2t1E1o74DORJ
V5aSdnphfAxl+dMSVs7YznVtxmEvR7jMMBs74iNLFxDo+TJw4sosHdj1qrTHY6xr
ERMzBRVyQ8mRNk7zvfidMSe6rqvLz7AMSEhH2ZE+mPPL+3uDA1hXBG0lFO55DJCb
og40ZTGlpsDQplhI17yyZ/Gq+VBWJxcZw10LlZ+U1m5ZrEixZFn6luW8fFmqaRUL
8A85Yp7l2yZiAhr8mf/wvnbXL1Agt7fPo1LXmPcIYIqrRgKRlYZwQxPxrGNLPUyE
O/x0ZurFcGHABeLMkcmj/hY+TTuWZk3kXZzE1LtkYkFj27ON8BR4Ll2DenPdXkgf
igAJqGhMvswVUqBdZlG/LlP6gf2p8SkA/OCLeTNk4syMJnXNf1ooghart+XfB93f
xfVszU/nf2jDnUP2QJ/eOqwFY7mk/VANkZ5U/fY+wYW6jmZt+9PvTd1qfJVU+kAR
hlqqdI9NauFEF/rVxRsBkE3ZQvO5eyprK0dl28Ign8775BdD1XJo2sf+cBhGcemS
VyaQE0b3KTCRL8qGtnU6bJeWaxqDx4Vkvkkqiu8eROlGfGSSfyyVa47UDQe2tTow
1oE2OYMfyckfRMQOSkL1kS8d0dHkqpeWlc0GAXf0GSe3n0TX+tN6W7cxe0vtkSfR
vwT1ixJTRwxhyL6UeiI80hmaOD2k+gbUl0Q0BaO/q5kucrPLiicubwudMgV8JEOZ
S/qKJFjuTKzIwuwm1TBoD7aFotu547B946H9vJ8A8xg1Xu7ygyetyNDxdMYmjoE/
g9IkgSClqXId288K4VcHH0PNE9lCESdoAe7sy7aWS6BVM297OMm5gWg96RLA0ZZi
V4rPa2u6wcTk6RQub+GYhBwEQSZ/UPfXraDCL8GlDyQ9MGlbkEKJkK0lmfAQAWkf
2h0yTjZcaIDIVll5Z5NsZYC1O6SnHW6vUqAFCzqzC02PYr7/0co4qFArxHh+i9SP
tQL9wiusVWOe5zElgiQcNzcqg4Mm/gqhpH59ONuCPGrMkj+mNve1hJfSQIllgZ0R
sZp262we+2afrstk306MilQCwgBHScqpCYSYvWL2ES+/XI2YwJ1StE9/k901d17l
13zXT0y2sptqmdyaGhX3QtQl8ENjGmnP7okJQlka3SrER/UcMeu/WE/Qy1J7UyHq
K4Ac4wN7kLX6WF856r1PjLPyip9waLCHKIVIemwqED8ppQn/ACV0zpQ4TPhACSA/
KZ7+eIoFhhpnqkmugKxH/5+HuiSjex1GGRIyBD7RH2f/Jx3e59+vjOMgJvwbkJaj
rOuAtlD+2tBfoaTCPZb0wrJlgfBNuw0yo2NBBRrI6o4JDLT/uXW1mp67FBOn2LdV
e2oYn8z3DOXlLRZRGhhQH08uriUZo+XiMUT3hKW4Spb/YTRHGJSO/INJuCBrkmFu
aQcIjTwXX7uSv3lFlhURVFOaEKkxQmREkKGDU5EbhVqZl2tkOGMCsaNrvlQyh11g
KkvnLY5A6A3XhOoNcZYh4VG8wD1O2zESUfl3fLtrWcP5lTDmb2VNNc8R+AE34R8h
8ri2nxQAupZh0/0dSsfKRBtDdY2troZ+pbJOCodSvoXF5dvanudonw4CdS9AqgBe
Xu0gtHOgPqwJ0G7neZaBlUMQKRYRPZp/fquBU5FB2UnQAY7+h+mDzNVtyJ3W92h6
JUCMF6089s5QYegRD7Nx1EhHqlZj6CAv8ZKctM+C9SMvPFjp7xrb3l1sI6Qr2+lm
n1YcA9d9zDcO4Bve0HCvQhRjlyWFm7/YZ5NqCYEe9Tsz10IYabhmEMYIeZOzMHP8
8XIsH+NtdsbhCTmqbcEDfeeHMD0pe4HE/qhiQVwHRkAZYAEBQOnKQtt/bJhlMf3d
DkUwKsZ9sDowRidipWZqaePyq1d13jLm2crYmDbxwDCRq5IFtdXpRFo2ypwzkExs
s9J1w4DJcU8pI217xrqOgZP4mU3NQiqg7R0T1pswU++MEFGif6fc2NABGoPuJvr5
imt63hsTCy+PJr3+gNLRpKMny1bnGDfH3UvlijiG4FlVZtNoXv/UhqVRRGq7mrHh
ps+WVfAvTmquTcD4synCD0b1NIoTUfCj4geKnoK3TrW1Ho9U6sl0VCBsEJBtA8zz
s2yZpNuFXBNJSO82qCKDhydumFq76QssmOS8Jvgn9jIyq5QxuKzUCQ9DMi8TMjXd
byGNRxYo+CWWSa9En2jAvlj8aJmTbc46YhTzcm7saOVNg7BaC9xWQczHrKpTRbmj
sJBJPXs9B2pOXiELqOAKsCRnEflm4hwcOfo9PMrXQ7fl0CI4ERmYK+RMIOAxjTs+
SsHwU5Ai9AsojsYJsrXm3C0kI1AjCX9PK+rYd6x6fV5VodOGq34ZebXUfidROp+X
OZJD8Euy6JYJvyjQue+vPngAPL/5DwpowPfmJ87FVEzgk2UrQhOjj7QcVjq0iF/K
mX+l22YhMeizr0KEOZZhanulNHc4MbPd6f+HAEaWoUC7DoJQ5iSzoY1M1TJkURkT
5J3unFT9ZJ7BztH0QzAQeGfBtkA9doBBbhz3GbX603zFECiZxiDuamtL9Zh+OC5O
VzJ880VhYkSxhZgHjA5nOLowIVv7BUFeU9gtAJk2kH0l4EdZIrR2Y/lslWk7SdxJ
fynU9fM2iyL9YfVR6Knz90wJc842dQ64uToyQptH8Vjy4B60n/1F3/cHpeLmkHVG
gqSdeeEEBD+4JQVcOfr5Dn5YcTaFEjntOcn1dPQ8J1rY8FPD1i5g3anEbiDvsUIt
L3AvDqEr9x4BIJPWTBRZgXeXzdLE2QHka1o0ZowAvST8Kqrnl531UzMGQ848d+pk
T2b0LbnqsvvMiAyvSNeuctqgUoYQ/00AID5oSY85c7sktLeHgyhJSDg3R6fAw78z
UjrDm1nAo4KW9uM93qVofkvolucVEx7tAoo65nkOW3tovbGa/2iM53bqVUhPclR7
B1FtB++K0C35DcXJ4tx4RL9r07O6k+B+gTfAUGhXiMz9QSf7I1Q7SGifbiVL0MUP
j4jkrRg9VpiHxpTnJhgOkDfFhZ0PoAYN/FiZ+Em/fjtv3j6p9oioLOqFhtbO0Iav
aRtX77DjvSwZzO33Kf4V1MLOOUTzLGH9L/sjhmU4QUukWg2mdGfH20FAF2kgUGdw
bMsieVAnag5bOs/2H2CCWLABNOzyxXQWly3lEUBbkKM3Wq1xa9G09jZfrM6EsWNc
u4oCMJo9teXt5LAiyw0xS9WmSjsuOcwWzHmkG1B74uKmk1T6+h3gyvnIK+8PCFPF
FrbagPhpulRc3TqgeUQihJ8kAL7LeSOKJproE6XTZthdtnH0EA/wBFrluvtjncMB
XKKl8RTjIAKeHKPgMXAs6S3FaVAxRqIm8P81V9FBQbgcNnlFuMF9nEQEziTvDUko
z4XnN2PDJo5MXWBoyRSQcDvc6fpddSl0wRjowRXK4J4JsuId33KdVMTVDrRaQTLw
6YP+Ryx5NZd1demouRb8Cfkf0arLEDH+3rmw3Oluru3mqsdN05Eklmsctxz09yC9
0axepgaEtmUcVPnTjbV2cAHq6Kf6o1T19UN31RrxdLxi+9v8Wu7DTh11LXvLHuo7
FXgNIfTDXTozNVume9ZRiOnEvRteN/b2rK5soWZJVIfjLqOA7dSq1Z2gLUfFpHI9
7Wpn8LrZ85BF7YdqMKnpaZevksmR1hKJWYfORaU1aLHUDqCC+b/m9Gfx7KBLtgnc
Cx1/A7ghrh1QFJnu9SHI7XwrCjIndJGb9eC68gdV5ILu+LjaqbnMYceun8ueDRKV
DdLNHmPfgnicysQWIjB9opSf0K/jY+6n3puHTux6ERh1DJbYxTs+5f8QlqzYlK5M
wEfq4hwmxDacWDA3ebQ9vl4HKaYx8iEds9O0karnEuwcNdWGsOY/8g4aY2UwO0Io
9FfmP0TYgJ8iX+KiQxMewfpdGrIDZ/VtS9itQrDJ6TXiuEtqR0+kxkNIzzkHQtpM
2dZF4QcrpERbsGrLjwGAJ95+0n42+ZLAt8nkQyEgYI9xlMO6IM5Srg3QmaXM3Dp7
VJ1iouj1clLwpo2/wo7laEqzrouwewTpjxt9DdEnzHpGItMpU+sh1LQzsl1WlW9A
mLYLCKJbyi3kjM8AnSINZFfrZTCnkJhsvzgs3DyzpjUOzoJKQAMmkxr0W4M61xj2
+/Lf4VpUkuyZIUn5yLeD0Ox3+GoUS9s6291ORmoOnlNIGwbSeSkctzEB9yjhWdaD
J5EP5rUL82AA/TmCwcJvBSNswNlYPF0mvD0IshTGixL9hKnfbBS6wObvIEgGxISX
VwDuUexFZsNB7q5WovEXcNS2sgno7988brPZhvfx5YB7vE+o6NkGCt86u/GnpIDk
LImcgMJsysiRui08tIjI+q7Ms95ZQvwPOB8b1SN1eD7vn0Txgh6VIfpSnXilWU8H
2549Ijwy/3W06NGiDzX9j1c/gnVRWMeUg8umMATDeIfLB4TiODQkWz5t0hH6edLj
dnRtUNifLSvQSSgZKevBN5WCYQ4J95Y3I2TVtNc3htcdCbC/KyKwhqLRpeMJpmrP
Y8ySP6BPD6hpOfdRPcv0IfsvfGUyvmX7hxoaO7zQM1gbmmt8OZ7QF4iWTufadhTm
Vdphbp0e4LoF3FSrhyPlpwyiPfigmQPAiYPDVtkGtTIF4tGgTkF65LHrUfjAz9pC
w+bTkPZLcS9YwMnD2JNMg+R7eSpPR720cMYbRpfslwzGOfEM6k5LHa0BH1nldb25
YTGM5SB1Ps9I4oqlcyRWHzSKq9n7FrP8scQmFhRpgZ1t+K0zyT7AFkezO2HRqeCz
O5UDmHfiZYKMT9ni3ssSXv+tD1ZUi/ZjOvgrjBpiaMWPaHqqr+LYCBccxZw+bVnu
zA3RoarnQA8vABilgTRt7FneJkEGuDkHPv6iHWQuPNVKsKtEqQKD2GGQ2rw/dMAd
FpSo1ubmMgf3NJoRRV8hAmeL5KlZ/b63vviVUslkRCwVpGVyo8wN1eJHakLhvERs
KXXmbqXwT4qQq6u2vRA6J8Nw5kagkiRDPNiX5JMsLZsLiiqMX/xvmoTwPqTfdPHK
pVcKSrKPFcn9fXhBLOXTQ4xmvKtLbpXA16Gg1m6TnT5U07Zl2Xk8bQNfJPG+7BSZ
4CY1Ih/36TQI+ZjozInBpkuhANiyZtyyxtKjnUEGd/vMWZCAt92NHXK2bMA0BhIf
I7ni+NhQXqbIQzOjWvDBGyoPytzp0b4wJ6LB1pob/AqXCiheMtL5I6T6DZ0twiew
qmCy4tSfysbekQoPuXAifAp4A/i+myD9ZsYdQxO/O3bY1s/VjKCcOc7Ijo8VDjNL
8lK/IX8cQxeQaXGwIxm67m40S48ykdqwx1TDAuKqQbGNsNAnysq3rT2NWMgROUa0
9QkN8OPAro53wm9zacLtGLrWZxLCVMrPtHXWRCDbCDdM+sTODRnvi/lc4X4MVyCL
4L4h3EGIcvYFCmiIbMwYDq/1CHwgcZC03G3qR6Mwye9858V8WoFUN2XRSJkZ9vYa
1X049caL62EM1hn7b0jhV/YP66JADis8AP8s3Ez3MuqZzvEOw00/NTC5FbX319vZ
LBkazYYu8sntAB9K0NcnXvjfNn2FZAooYmjHRqaxdgssCVB2seL4+KAMQ77JCvzQ
CAtQK73QB0E/5lLdtW1zyT7XGQoUBp70Klb+meB8BDr00koA4/gIDncToYfwL7xm
vVryBfkws+/YpkRX/rk/sH5z5bRng9W9F0uwdWbzPOTTvUgGDclMLPuOaYwFtVHl
SBN0wJ4IgIeO/Vbmlq90Qfw8NPXeEBAhBiEOYToN9CgjouonsNnZ4ixg/r09W2ij
02bL0/svhnyioL8R/pmWf35yt9TfJ6MKL28l5vmiFVxqkgg71IWSJbL75eR3yh7f
AEBrPKHxOKOUxw9mtBZ1uyz81I6aAKAkSu4F6wVX5cF5z1/dOG6HRexnYkPUd0r9
nOZTryOMPRy5dZMZUVLdUFIL9ekzSv6EEXHmb1aoMgZsw3vfOdpAvwnQsHEJDng2
lFF1UJCImNpF6OCHmB34+eSueOvIiWbXaewGldEj0jheDF29AflD9V/YrHAgyzVO
XXZRMs6ydB2F/Am/Id7e8mxXxypNYylVDnvJp0uS1hk/nrdNFIGfo3K2/8AQ+u2s
D+ZHePF0lgaIPXjgURwSeBdijtSFukq8QntA1c7QrsDf7tFD+Mr/6cAfQcf8JU5z
gl2DQk2LVbEMfSpRNfShT66eeH1qNll91p2xkejwFRfW1bKW9Lof2oQOUpR/0hQv
d6hLi0kSL+a6SgI3rFOmr9r+3kZI/11jEpYLZeLkCViYQwpjZXHgWzQDeomlhjXG
JN+QL7E/SQ3KYTSYWX1c09toyuuKaI+8oW20kYlZOb75uAuhdCq7dS+yFXN4ZSWR
ok2jaSeMgLdQP5pGatkVi52cVs48UGfSiYCfMZrWrIO89MZ2PcHwF08BRWD5eKCb
zgY5hdqZKJaCBb8icKxInkyeNBA8WWeekAzTQcHG7IStWs08YKJRnc2gjdeKz68w
xPlCAH7HkdT0VqKQo1V35Cls7dvTzZFvq6B1Nr4mpw4ujYWAWLGbGmJFhoX7kq/n
Dft5XRJVE7QSAfCQs4ip4psICc0ewg9Z4axa/jI2rMXIXeNOGmBBieWouni+xqA1
KKKeBBNxAUNFErsE5af75++H9gO0L+kHTlvaOb3+yEEKULhpMsUtYe+Ylyi7HRfp
vFK6ienI4CdZbyeC2iNj60rNiT+npm1AYlY87i6HBLj7YaJyaDs75B3wFNVQvpcB
UbFYsRB/YzRVLHg+6hopkqD7gtYSKVaqAtpFpBRt5PX1EtydWokqi4x9f3kR1oVe
LaiGAbaJuvFREUpZQ4XKC09A6m+t+kb7ryHtos/FmE6b5NaxyMpA9WJSxNPPIEGa
zZpMSZj60epxzL+/tYMhA9Z5/ttID7lLLtuU5Ig2Pc1iPOsAoFKz+4/vMZvpc8AA
mJMHA1FblOhmWP3ezZQ8pDZL1WoLMliPLgzZUzc0X3o5++D1C6M5zp6GVf+F/evE
gm5/y3obycni5d9PhgWtdxko/WoeX55XM7U0RgrGF8zLtsdm+C4roz9dLc72ryrB
cxkft5UeAaJ5No2z864ZK4QHab+ZUUqTW08Lv8efNnEnal8hLhwX+/0ug1VE4B+O
CulhzAlTWdJ0qknk2nJwv/3mC2jDLd4tuD+o43jJNdm4dDI1Qh/bPmjRXd5l4TxJ
sOH+DWs+t7EDYrZ4o0pnFYQm4NmADoPzW8jGgw3jJ7f84LMdw242cBiYVqdwxZHr
LefPv/OlY4eNwcyiUcuG3BmVHc3h11ccup9pnmJwoALahiZTdWXoojqVzoxz9XVf
DY5ok4tVZSbrjqx2q9xzagliJ0lzX//607lZt54ucLPuA5nBsN8VOcVNLSO/YV3v
R4RZDCFXikpNEtPqEJEeRUvPT9GR92dDKycykWsuRVN1tOD0IvKXQlVLY04EO2iB
1YmV82hvX4S6/ul/L/UAzRQ996fJ3cgCFwPmC2jvFnUXWb5F3ToGUiXTLCr8txcj
Pn6oa+ALzvo4IdwszXq1GeT/tyuNMICY4B5imXHVg5M60wNn9ws7rP0/vlhcLtBR
wzNLjPvQrM3rnLkVwyQBOy/qFdeP5mIAVIjVesbkLMGtT/pf4guSFzNZiYx4NdBF
6Nl0Xp4j6HIAITdt51GCMLNAIqlbpugMPKTsyjRxxLW/UILHy/q6pT7OrSRdIqn+
wKUpFWUtCg6qD3Nowq/+sMtSQq7WgfanReRucZAQbLOV2HJlXulOsXi1+V1+k6no
ZedSxVXP7iRrkFi4GjinALzJtn+adW4uRFOi9K37gkBFwns/svAtVoivhq+gmKyR
94Q2sxSxa6CIXZ2iMBcjGW0TShs0J7sVelKEISFCrH52k1qtBu7Ugk+Yl7aL44KT
PTK5bisJKDzgdIm2du9zLJ9lFLQorJkPiw90kTkVtLHngWQPoqeeRUs43TUnYlvn
UPOakgKbfK0YFwkFZ6NnHTMAeR6aeyIXBdp0FvlM+zTfdOn/+uk+36GvUez5X+GT
GS4wmwktlXqYyRbVZayhTUeSTdH7dwgiXjhK/iW7lFYaMHwJN5dpds25aYRo/+6X
GwFH7Uo+3kDxcxRLi4lbg9ep3GIdV0bXV/ih3/pF9HVSCftrZ69zxmwtoJx+VLSB
6eRPoegAuxb4xg+yrqy+QWFyPs8rcyzfHd4nEcsJuqBNL8VpE19q9ZzzVZH/GUpR
zMBkU6GhUPAwG7u0ff29m3K+WZP8uwNzLafGsft9SJZ89KuC3P5DQnKVtQEYcZAj
F97XW7sTIMi51jESTvDHsA6yqylJIV0FpRl+eissf0slWBcyBygG1lyv0JCCVbhK
norJwj0xjKjcKVkIZtPS3s+QeOcZhXsNpIff6crXIsUu0clnA8fhBC3W9JDt5Te3
CK8/+ZnUIAUqWAIppGf3O2XD4heM7+LmK38SPW2bPBMKbk+W4fsvpV9/IRbA7Qa8
uMX6miB6xoSIirgI4ziu8GMkXNKqpQIghkoXOLIuux2zonoFGGAYHrkvwrqWl1ev
gDpJ3tLeR2ayxNaHKUCT+xLnZeUIhT/E7vftWg7YLkLqM0KaT+7A2iEf4yt+2PO9
vQSXel/OfFVPxb2rdaeBZxH6UKonGI+bvPrhCsn8mhAekuPOo712wdnNjzMdTx/a
ON99DV47U9nbqmI/FsnsZQXDxFDKBgFWkHgWZQj55H9R+nCYcV2++4JemKX4yrgh
MQslgMLl+mkJ4djDT0wE71IXcCDIQnS+OG4sDZ5W30aD2LgFta7BtXBWsCjEEBxE
tFF0dIr9QItLZC1HBcAXG1ox5Lc9foDsfBpROea0xJB/WBxyAQ2sLQwS1QNzNS2L
Yrk1K3/KbjoYJDqGVLaGZHSh5W5jC46p7A8WsfG7OWSRDza3KUJxqsgjy14vrqjg
a64aFTIedcV6wDAXBjbYr1s3/l3HhReDjQNblIdqT0Ai/b9TJWJG7gm1OcRKE0ww
7EmUJerD2iXvD4k5LQ8Q/Idxf+5IDVoS+5juPGlC59DzL4YUDZs5V3CSA8A3mib7
W9QNfbCFOZArP4LLRdOdnyA6mAKhxvLpeOfxkXVNoMFEaJdQ/kxXgjhQjBlIlAm+
Bjxify/hvUzWD5aSzVS0sXZQcbtPy5tVkRmIPynEFRVsOKSX8zNX+C4Qx6XGLXPO
SZwkMxvvoez02hX9fkEQeI5C3zlxuK9v1BakoDqMotqReYr33MHkMIXBoACKvNIV
1QNR7x6KrzB4n23RxQXFvcSqoRw9D8Ki1PA5AEUV/7FBRNyzjjxZ9F0+HWu9EPkM
hx/l/Q6QMzO5hkFEXAgqL5kdn1k9lrl1vuOu1CtMT6uR4tlOw89hLHeA0QPoOooU
zAymN0Nk9jB08Q/w38dEAePyeNxgNdNv7E1c0R+u1bSP9p7a3JwsKjidz+P46aqR
mwIeDZjMYq9hUy5T0UmAEJJzg8zhrimKUcPTofC4LsHcY4xAqixjzvFWhGAHPGux
tHNxAWIIDMHnZjGXhfDrGG3I0wH3Hwav0f4oJov+EA9ZpJR12gXIhWyF8B8+cvTS
312/cesJ2K/1mjViWi4XKze8nQ/K7ypCQHS7koYc+lry5gVKVt35VX41go7IiBXo
ZZPY3trd2ldwseM7BOaLr+Gjf4XohZBe5kWr8ji9j+D+ZCx3bq/cUKIHJrq3zvZ5
i0NRJQ9hM9Dg+JBA/iNSH3sR2iYj9VoRQ6iV3Zl60DcsrPH03Wz4oSRwAPi+duVi
+XBnuBrfoIfmZMswQqpry5i4xe7X1TuEBbASyEuRySNP13Y20TV73ZaLfYQF1ddF
h2iPDLqkhktQ+0mbk3xiCUJPCw+HXft5Q5EZmKXX92+csfdd5+Si+U/hCI3rocI7
gRflveDfD7OeHm37xa+XTTPKJVm3aThQ0aRVQlzJocEk8z+JuGT0IiS7vlibcl6c
CWdLQKPCId7I1IhBi+bJK4sBoCFRQbXTt9PWewlFIbQsODhr93tKqtj5/Bdi4W9V
Z4dECdrmZcJFxINEIplHD1hKCMobVqA7YkfRY94Yv+KqzqBJz9UzKHmxChLlniwt
aPY+4ADANSJ5oammoU51QVCE1phRxeLEySlbxWgJVsqD3lIUrw0J/GrI2emMlGUj
gs9oWg58O48tx3+Lt4WP+cln7IvLpELQ7TvXmBAgmAnQUbSzFvpJqUQ6jWYtQ+Br
gC08ULRv3Igp+cclw22IPzVtEQ0PZOIheiSyrnlHCHowe8mBd35cqxPB0fwtNnEt
jiHTuVdRZkx5K6l1k0JDotXj9Whunk9tJoTx68ArWIzLArjJRMLopvAAiR5uJLD7
G/Sf0aJhJcWWhGbeT1t698nwjMMlhHyC8bl7mHoKCouLD3KEhMfZKTzFGjLHgNv6
kHVXoOh1hybYxGsVoudenPXH40XUy5abl+xpRYKx+SlMHr/tAFMj0kKrR1ytajYX
nKtpBU/8Xhou/QupQaFDa6Ed45y6VEAgUUTvNFXVM31sbISvsaB7NbMd07c+R0Pn
4hVCNJ02srrSxLSJ3pHHwXM3tjcwjF0TvyKvyKYYpNsormXkvised2wr0rS1BxVk
Onma2tRKakTUHPVAhPv0bgE76Q6R/HL/pozs7K260E6xjkUTuGRvU1ILawIv9rPp
oapy2dTo2m/cnkf2qz5ualOpIyw9t30WhACtgg3qFHu/dyaDKS1qM+pQbiVhowa2
/ctC2tRwLjUrOmoJ1gIBxIGv/VVqewXReaWLt2mXDyARrazDHpSWYzgpQOzngWIe
EA0iGCHqZH0CuHJrkv/aYAiK1o2xHyQkZb/InD5m8htDfg8DHUtQTTazMIXBeoWE
47el2hzQPAgjakP0xjT1bg0UZLqFAZYRr0WwjY4T6/k/3DkS+fCcsapIdny8Gw8g
q5j5iLD9jAk8kDhK2nGlieDOGid28dX9fKuRuBSdqYlP8EQf8tjV5hBkqnptwKJ4
MPdbsjVPdOKUdw3gL9jpygF1H+L8bMAfZTVfslIVEHKGWj4/1EYAc7PBSCTv8+q6
qalLlq/qLhLx6pkdCP+MGcWo7OziHkbBCriATfwpv2FxQ9mlwXiG60Qzgzlx0w9h
/Bl1pNPrFIt7iwwZlnrz1lVD8JN3jni06Q7NW6yAD7yaihIpyCtNmymhhc/w/n5e
kuMuLe/OMvFGPOL2GJNpQGEV+b+ruLI5xlFW96dn77ASLef2OIICh9FeGl/48HC+
xsk5/Aq6vzXR9Pt/e+R7hs19mgy3FzvhvNXuRx4s4UAmH8YqP1jJ6OuXkS4xHaCo
id6brMPkwt9jjwaTcvbEnyfN6WKhJHUTf0VMIhHk/cARsPn9l+cpncmzaWnGjh0z
/tf+8RQllTSVJKrdJK59wjlc+MNJ7HOhBwAQZ+hVViJySc9xRf800/1/IXX850kM
ECR2e9g9Yhr36RBmBIoYthTMkmXa6ABfwE3uZYAPIPVapXD5YJi8foxJ1kn6c6S/
RozjRwEN4elr+Ys7E+v2m8d9VFolkBjdLh9d68jSM+PrzMKg2f+7ebfGxmI92Vs/
7UGMaAljkjT3JWDtSG7oySGnxY6n6J6onYF3MdCPUnM47V8TpABdtm0SvjUmqRTo
+7de8qI23sIZ3gxboYqfw2whz409mtgQ7DQNtibzgzOB0mpUYex2QaBu9GSPuu0a
qodudl492iGWVzuP+E4i5cybXNl2nIXNwPfyp3t9n8kAHEVmEqYYY9dBH29+UuBM
KA/MPtk487vFdA5zINLE8DV+HGYA6KaqY0IDa8QXtkOaFFFOoLBaFQGTg9YKJopQ
ngio0X96pVc3ILUL6gGE+Cy8H4Qcy8ZJVjQMZhb0cqSlwnjeFTn/Du9AWtt8bcrZ
xbnT0Nx2GoWYSz88mpNsHy9zU3/aeFFV5Ham9a32Lpi5qQrpG/MWYsNo/Apyba3I
PmZvSm3uEvV/c6BAaZ+t6UGpIgNeLHtkKu+NRFH5/opLGYIjC1dZ3/6wSAx4chfZ
qVZQ0Sau4hFgslFP8hZrduf0T5PWO6lDucsyXJz+94wV6NjNs05nJ+/HRCC7x56R
kk5pae9voNNQz31EV67wFm6qmQ7Rjt8k2PO/wvOjIeinXGtN2X7ytjXDa1UD7aHx
MoHrRsed2OZiLnJeMcd0PyKrmEWAZVm1wGvDJw18+rEiLw7rDmVEhIz42kDw5Bs4
HL+ujq0wmz8/9oUklKavh1IbQsspVc0R308CoOv6W+gXbz4BJIghoAMplRXDDbnJ
2VLVMehnKSiBFAoMyHn71vJ9Ch+DTOViszoHYnJ8XywbWQqbnUxPN2mZSKXCsyUK
VOpdKTM43BIj5+HNy+fUbZAQyEVWHZuHHokKFlUFMsKXZSVRIvvMDk/YWDxwUx5E
CkJXlK0AptWw//NGd6n2J+yEgXw8nT0PBYrKWE4GOaFspwNRg3OmPG2ldUYAqqrA
yGyKcj17Q/4s84MiKk99sX3OCXnXa8j+7kjUtrqVLyyVa5dp+JhuW+NBTBT/IRR7
MIqOZXNrcvCsGb5ayYnaV5rEa9jqalo++XjU/RB5Efma9RYf0+doXKMKiYP4KokS
aTgYs1S37ptBZqAWUUn/pfFn3xCIuX9sgGVYRBL82XIisV7uUpjtTe9i0UUY5RhB
tETre1RRLpvqTWbzAcUeHAwpn0RySiD1ZZ1OPzyRRdbL0kaDOQWPqElkjKrsqRJB
9gKbkIZM6IB+e3ttu75hZhUYeAtd9v2FwAv/XN6kjkrIsXT6Cll2ckVk935ywvuJ
38UCj1cuizuK5qK/x/EHqwjsOLUfE61IdpIlTdxbQMRH0ABp3FCkMx/yNgkL38ta
pI4z4qq9tc1irXIn7CDKuhbTduWBgrMNDUtXVg89Mu1yoKQ3lp3z3PnHye2cNuJe
kHIBqMhZhzVCNfvM2zem9m4iK2T0AzMLYymN5MVY6RaWk/ICbJkEUSzRtP11R9l6
HqF07DQkj3GN+ZEHrk+dhB2rcPAqBE3Cf0jTD+HPMTvq2wR93mBdiUflzUEdWmd7
eTEn1y4sNfvCtcwzoMxmqIdOUVi4d8wE/nQpxfEPOXoT868A5N5SA241TmUTH1xa
TN2AGdM7pVsu/xbwA0XxT2Y3zXNP2gWW1zOKMID+iV+R70A8YctNg38+UFMZn+fU
JUmruHr5+pWZs0R/06g/4LIdOWl2KVAZgp7onVdnVjVvHR64r4V0gckd0NHtFBR+
JA0zlREvY2epzf26uS7+OARF1+968R0jy1d9BRoPlf/4m6heXbkHS40rhAOl18R3
Ab9u/t/+Drc8hjVxYw/n114sPoRE2WNol4VkJHPwpw657sWRosy9P2svYlBNitkq
wvB/sWF4ZyE7TiunFb6WeNRsJuqnM2RKPOv0b7BCsvCMcMI9QqdBsCxjK3HfEhlf
HPh5SxIut5XMoT2uVf7PA2TUO5pYtzhVmKgx92SmRQEBV4oNTMiT3agXyoJpkAci
O541UtaihlNhF7lB3G/mikkOEl00u72wPWA242+SANaZQP7LhVSfNZ9UcAkFKfRa
IH3sGWgvTwVELe6NZsFKd9E2Zti6jP/2lSsNFmr2ZnQ3ZOFA0BvoaG64YEV4EU9+
nec4wizXoM/YAG4L73w6uJmI5gSdKRkPhxO/f4RxQoVKd6hp96Avd445npZ3AC5l
RHWKHSelIaALjYfuKY+qbKg869UBw6l0Yd058qSKtXspYIH8TGTFmSyVkQtzHtld
JXUmN697cjEtpALGoEMxj4iFATMnwetEe5EdC7+tEDp+rPDnzGWNZ3XD6OJfXzG3
af6dx2ZJY8d8tNwiyJ5di1JKb7owDAqTFQZUXBuC9Kzd/bqdw7y6pmZLwRQS7xF9
qlyvfEmX6z/arr8gbHK0iW6ypZUNBa1roAozwqx8k1FIYZxRSO7GnXeVRwqjA0fG
z95l/aRf9ZwE1pZmue1pux0cg9kPfg+Zdy9++RgBc0UfaMAI/yUMEOQbnxlzqkn1
/Lc89bqnjqNb6tc7Fpknrm5LfjWZX34DOYULETF9+rJ93xNkLufw5GJFPUDEJaY/
sVHn6sL6h+7cEugp1wejzvmhefub2QUVHgokpiHP11YqvXYiGxfKfMm+tFG8XlR/
AD63hViXqVcE66PoBdCrletYdpjrwFU7BNV/5epYtTifT49m3r+K0k/QoM+tjrUn
PHYCA1q+QhwOi9c2y4Q0MZJmICLZtjH++q7/XXgjpaqrFGakM8ES0iKZ9OSxlGiP
L+HTrXxGUWs+GPH6jy1oGJ44BDYeJQg0lmGUfuBkvETCwUyoDNIK6cnUGZjkW6PL
6aUYs9JlQYEnP6Ndj7yZFVr//h/0CEoIbbhLUZAPAyVpwQ/JxF0/ivs61xnkY3Kd
Cpcdtp5Z1frWyC+eMdjV06eZX1laxHeiKhSXXyiIrJdvfQ8VzyuVw2TKvE6uSV4Y
GjUF7/q5gjXWWgzmzCbbin2gOQSluW802CW3lLtwPyyBR4gys+Jdsncsy8wvePjU
s7UHKsiKiNDEIsDDxTQr0AdrT14Ab83pvmC5cLs+5vkN3i8Ow5mt6eCWF2Ave1rM
EyhEnQErBigKjoDVL9cJpEzwg4w3etzmn672mgQyXcE7u4hKnjs391ZFhEpKffrb
h+KlkmUlljAb+Ir2XrJhx6jKZAcbxDmmuZdDGs4jFJQ3xTdMRKD8WHVnyAaHOgED
m5qm5h0eNiuMcqWcJNFbUncDpRgYFCRN0B7H91PjZ58E1KYlB5qkHigvDDVwxuzz
FnbxxRwCf6G0rE1Do0dCMlr/o6DQs/KqKeu7zY10lZK6pSa/1HoB+wqgTh3xzBpL
8JnG3wyCzAHpXSzL3cxVzyk5P0meb/OSiGhiidyN0A82XwoIXE4Vk3oI5gfSE280
oku5YBEPlBhNSozGA1DHmMYsS1P2ld1uIJgGjzL5OrcozOoY43vwxDDAcat+9hkb
yfDgxuk9WG4HIN4sET/5p5iuGNNVv9Be4AGG8xU3xWzxM8eTA5pGmncBFrpLxE6Z
uLQfcNly7phSVLSC70j96n3yYBayRqQvGx84v2DV5UoOYx7e30ovcPCARuVxCciK
D/v12Y/jJvSIRdVUX2Idwz9H3bbilRJJkOl5BF9/mlLTL1OFqgfxzenzl73/1eHT
haVwXmhbubAPBUHfAFO32FGj4ojXozxpNhJ0ujMPpydPCrySr6qo72CAnnPcM/8n
Qssk1y5Cof9wE8p2x7PUdpTg0PMLFQ9e+VGbmrgXnaxLae6Sb8mlYTmgpU8S4Vw3
in+6sqh2QvXgVV7dQWW9kn4TEwjjchPAVc2cAPyWU0RHGKXM9K5SCGhS5JT+Rc7p
RFvBVQEhONP69QoUiiJmT4g03yDmRNXI3ReHownh1ScePym6kqHM7czlBq6zV7Hd
YOcSLxxQ00g84jgzl9umFvCovdjlpP8mGKE3RDQZkpcNdJlBVFVQOMzwJYCqOC+A
EyyA7FWeSKUK1bR4nvVEkhIe6RyKq6lHdWHuvHSgajyatur8VU/Uc2gYX2ngBwJd
KvpLLDn3P6pmYP0BaBrqxJXxS7bpmoPBztxPY7uBd8MszwrbsTNk++ngasEGcyQA
/2DsS7sLwdoyjyM72R6LmMencTUhm1aKjMXqQjtAP58D054fYZDBEFa0mXfsOzkL
7x46x7G2G4dUYTtk52f3qMsZOONkSeo7cLrU4FopeCndCnaRQs65NDiZ5lwb+Y/L
h1CsGUt9kMQmVfRM+1l2z47N6I4j3TLyaIu7HLBf94qE5DLixqi1LTKvW0QZcTA+
fTLZ1jQOqMrauRFn4kl6im24rP3W52vLLfIcx8NzAcSPMOGZN9xeM/udRQ3DUCeo
WDBqvMZtPBh+YWPBw239cqVc2CqkPMXfZCNAsa7HUyWCzEOH0j3+okv7pILffIfp
N56xEt0I3hOjjNtaath6c6iSF2bx4Jgy5S39z+myrx5E3hueEYWShiJuRlvBcBvr
wLTAaNEegOjmVMJ8mrDKHbp4Ez93x3wV8XhTWJ5s0G43r/ky6om8997yOixm127R
dleAOJxzYm2t8Om+MqJXTlYamKo7xxpzJwby4AcqqoSTFk2PLbBTbup26Xi/FV64
ZniIhY6eVmPjtx4BzqrGKUYThuQTXA+ShAX17ws1p06MFRXHYQzSeseHuuG/G7up
U50YClO51LEJlgKwKLSg4AQ/wRGfk0pxNS57oXZnnUZANFdSASkPhrC0pjf5dy+h
NnYfSH//g9g+iqzV8HAlGX2RoevDgfKB7BZ2kZyQYTRHdSoc38WQyRNwx155n3gT
dxqvELVH7Gb0OV9R/w0B0yJcLAZpfw2CUIYqfVjXv1P+p2xqlzzqdwN9svFsOjpD
DzEU+ucyMbp3VRyuRo85mTPhHt+GDmBag11zmcjteGS0uyGwxki/Hc/PZ01YA11P
I2xBTPIQMQx4edwRqKazpcQeYkOPdgvedK7TNJACAe7NsW1UNH+3h9+N0xXyByen
RNVO1KNOv7Qj5qwMKvcUv5g6ES2Z1pNC6P3Ho3ujDnjEfH06QNWJIUZQWXqyC08R
2KB44ok5PBhQ4ulVQkF/ccpWR/fnhkq7013E5yUlvnVZXvz655uDw9N8gHRQdXta
PH78ygtgTkFUe5vtFznAHkEcDih5zst5/cvktbUH3wcPn2ni1QuKV+UmvnVFerLo
RmKVFHraGd4dzqnc2yt1u1Q/ENflkDivZ2ZH9JrC+pwKGE10CzFZCswUHH0dFlb3
Cfg9Ebx8LwaI7IdAHfMVABF356X49AgevqX9YpuTbukP0AWeaUyqVHnUpQVyjAWp
Jqv/vXCLj/5cMBtmvTqX1T1bp7trUtn3hz6KgwhosTPh6Hh0jZwxCACeOBbZH1rD
K7N0W8ZIns7Jmvh2i1dCG7y/MPk8jCTxwM3rz6JPsy5PICHABHeWmZaMvPRty/5O
Gg75o3jKccW0ZMk5FP7I0o6gts0pdUuTH6JQJnd/0jE8d0JdOLB183q774SFzpb4
qn2m+gkL9qXGCTChhzM/BNVXVPjTHAtikX1VZZqyznYSic7B5ZeKaObz04/pcz2i
YJg54GumnKig/0ch4P5L6YiHsMPUok5H0TopPY96qDjt8qq1NXWECEdJohqIa1gY
sLvrc4y7b/l3WkW160tK9YpqAw5Djj+r+lAWH3wYGcOgcXjrSu1ZDRc6E5Pzk25S
rI0sQxpPpvZEjBbFX4Loz2PC//cugJ+v75qXPw4LU99DwuI3n27AOUyr/Qs6oUdN
80RQMcYQeZeqQY+HeOoxA9zaGHJ37fMweUscKXwTXmV4+e2PMJwlT7KuZr9KOqHO
Vk5j6V4auKKlaU+uRuLVv+w2xhzoo313/sGXU0a5LV4ciTir4hVzWD97xCHipOgJ
zWQfMzKhUjWgnW8CwojP/Y16Hko6R/Y8h9ETt3hoHA5LSyPt9gLqkb2BGw2Sqlfv
9x2a+yEO/yems0dvp6KHxQIU4bOdNPCV5rdIrdxO+tx4pgRIq9DF5hjsOKei1/q+
q91bxJgcOQzaQWLGHAmD3XqdxBfq8Ra9OAibr0D8V07CZe3QGIqRoHSVlaFCbFr5
+PBooVyDCpWKwJyohHH+Al/IqlT/37EbycjHm3VmYRw95G1N83ZApNaeBRwWDzGh
XzPTTYfJPka/muYypxdCkOEWle7sngIrG1o7hvhZLuRA3s6OIEOcl1SF7+QtVzMQ
3P25VghjLX3Z+K/RnwbV2L9NIzHnQ1R+NBYxaswnkHID4ZPfqcYF+rV+djZjgIxs
4XQcqH6tUguJR9F4TWN1z7707o/czs0WcHcTRW71JxZSVBNJD8y4nlN1RmZC5oMb
sRzYm8HR+2K0MyZGeCiVWw2rpI9rzXQ6TArJxcmYqrbPcLEsS5E62I71ktSROEui
FWJWJcWLVF9vtQvW/O9Q8esHhNnOaksDJ3xTlm79XMYXEIMWgEQdsoXx3m2h1pAA
FsFPdPkcKX/HFWVwhLfLSk1gMxQgzQwzM6RPRq+rs/Hlqz3QloaLFiLiF6uLx3CS
kPnFoJ7DizA/kCmGrKgUp6IabPv+c29F1t0+9832QXcYUZAp0x/Zww9Tf8JmU6p3
59rwjfPMD82vEff8tQCNNXmdTR3sIXUYw/HHK8xlqfh9Xqns43j3U0wjv5dfi/m2
dWlyC3Nd+ituB9ekkDQwOtKHCpnfucbclltMbrUgi+GIylLLhRT6uDaCQXncyfMY
VnBuk28frFSiL+j6CAW2tTC5MRunADnf40DqtXGzqSpqVDJTgtpo+t4MTsR1PjtK
mjllMBBK8yib7SchRtgzPazUFX6Ne5//NnduQTl6ALGRB96s4EwLkzQyz4/7GGNF
Ic6AfGMEwmCs1iwViS0gTQP0QT35nX1hQhSuCqc5IXJQLhoy/jtMx3TL+Hi4PSgf
nYnuAGsOIuhulH28ktK/IrisLwregXatTtFAO/6GdripxTB2ZXE9Xva80JbkBOr8
cAEYg/Dtqkw2OUP3iZdtdK837w0dXxdLAWjevg3LAHCme+DVSiKn13ZdZTfWMOzr
ojeQNm5Hrywy3TPB0LgMUTbmsjZOu0rzmZJcIa1FufucS8SJmkCJw0n7f7KkAxpU
RTyd8UVX2rAMGcTAgMrOuUkXaAWyLJDOc7D0tnv6ZpVAyisLJtQ0q4TYMqKvQme0
4kTy6pToYQH5kQg0u5bBjvxHB7O/qq1SN9TMoR90a83zLXxeMP52Nguw3hYp850M
GZ8INZ+MGEMWqNiuecQq7BfImG/gyV4Eb7CO8bPhpUjvJMslsAX7Yb5E2ESj0gBg
gERK736ZnTog3dsoqZDo3ch45l7gmsRS2I2acgldyimKPr4EcAYPC9afa8sut4e+
+OsDBBJHhBwxVr0jA4G4TiuKewO73vnSPaeKiAxQDIbV70POpIpkEzntnx6cqRGd
4W2BcKLrEspCFT05SJz+Kh4QmLBDQB8iF3tnJfdmuEeOp1ETfsj4fi+NMlJxkLHx
M1YotIRI5u8TNKWZ83KkqsacLlGrHWNeEqOmumTejVyrbhJ4Oo77ixyJZPYWeQ/r
RZLI/E4g4qkNtWH8UdTPcyKW/LleARpgDjOGyEsNI3vG6il6Hj3hdsHjkK7AN4Oj
fTVIS7vNZbt/zk8H5FoL+bBbM+NnWbUbVGVw8XVJJKaVmhuk5lc8SCG1oEAjaX5+
EgPuLs1TYwlEYXEMoXeg1vrgmDo73jpFsFBi1KiyppbTPuYQGlVM0/SQTOuWO37b
L4m2db42N1srZABbJxvw9YlMiNnbWctQ9K6BGeQX+pKP6GuQaDXMM27JVSUoD4Jo
uz1NuLoz0x/DepW/LikiQmj1GyNJ8IhuAw8EyHZIz4t+Ari1Hiog1+MzAcJk9YJk
sXMnD3axiPyV9gSZH5TGHtfH9iGKCE+IBNwwtQFnUWeTUuvkCc1j8r9kK22MBS0v
Yx0wIIqfDl4IKRJNQZQEonKY8Fr2RjlwiZrhu1tS6DYPi+lkmMhorstIxBtJCjoJ
z635rRig2U70g7S9FVOOmeoYiVlS01F2UzyVV8SxEWPn+wXVAcsU0AUlcc6In33i
VPFYS1tbdWAkYELD+OuAgYSrYXqmArZeMJvb3l2shGR8CIpzM2aXoQ1Wmg/Zgene
wkFAq4MhIH8YwrPe2eAc7LGNkDMPIx5TkivuIPpNgUY2gm6zOT8F7XAn28Rpa2iM
e6Hj7CsgyEs1c7E4dvOdaeLpcziHIu+clYFQ8UIBZwBkogvgf5lX2YppAwrBdpBI
e16Ee2BJRPGW9j5bw0l343WEft7sY8TBVnYBd/pQC58NR3wb07VR04kMKRDTs3Lx
M1ljrdU+9MDY6ZCAbQrQNWCamfHxosjvmVTOxqko0/KW57b0wEB97oBq4gv6wbuv
IAkPAaYqP5qVRYzbjgyrg24oJ+kd3xOwmkqVxNODveSBUppNrD7i7lipHiYgIySW
o5VLGHWxEW6D54GCUgMWaPcZctlkmxzvAnxoe67cpcMGwR5x4F3wdxfyEarERZ2L
Vbgkb/P9oLGye2M7VnQWsGse+OkTfS8MVyTexaM9O0Y39DX1JHy9G86qqmMimmFO
+g8MP5GPG6b4yz2CaCi98hrEiyphdOLJN2OrbPglH9LzJhPr7GkrORKmFtBpG+dO
znvmI5ArmE1SUWIp/sAu3cqFmW2p4fzqTbpT8e4uBF74E3k3mNOTehXCSIhUm7R4
02fskHFBJgqlWBEwor39KSnvfkO7XNc4Dk1i9CwVbNCuWFMLoYviwKmGeRoAA/nE
no0x6u06FA2N+HDucfMj4yEA5GrfkIkcotllQgW98SsA7+DmQyn/owS+vSyy98JZ
2z4G7TxFZNXgpEJFbtkdgpvOqkiA1kDvtOXIKLi1NVrV+5Om2DovrtY6ycI0TkC2
zgmhfgKtsXxzncLdPrxglcic6qV6AzpnPSmdWCvTEn3vpLLA1dzTTisGA5v5x2jJ
jBhrqzFTFuJmR2bxC/ipTVwOcVC2zga2xjX2r5bTLVhTtMLNQIv56s20iTNC8zCA
CwwylAxvMPVjI4CtkyZB95PwcrTr77AFMyHOJN1s6NtXSxI9K+z5NYqCk4jmGKUI
VP0XU6hfS1z9NhSmIrPJ38En5Dcct6bosVnaYOvtKLd8TSSgv6wS1CFTsTt3KI+G
qN5NJlnRC/i4SE5TmFitCxvsSSBxvjqMmllt0M2TYvBxuAUe7ujGYNS/IG9C58vu
WvRu+Dw1LHKrLSMIRNT4JJOVuc0Dt2+voU3ymE3i2n38Qs/MHCV8iKKEK55KBhwo
YZ8jjGQAeILfLjjWXtpJOcWFwRlozzA8YWf29rwYH+R41HKxeW5DroeXKvbY3tav
JQf+H36yTYkQrAhtjeN2GGEDJTqZhBLuxHGCbCBJzm3GKPEo/wfPLmjKlXoi+bZO
Ke2gHBM2nVSBHAJPih30K+aFmH2M7c9v/FzRG4yRkk4YqzCkAHIz1kiJdvsg+i6L
FPak2tECIgd2uoyfo91xKGngznDcBlYDXx4vXRAIqATLOSCmMFM5g4/yN8QpfBdX
QD8CRofaAmssa7CdzZxJRitpbWuhzQscRseI/+0i+V7wGtRTjvMF/6o+8DAs99jw
+IMMch5yGPtm1fiZEc42+5KK4D/5W5zmCllf9HoATe3mLqCfI+EpIkh9j/aMiWsU
Yw4/p9jZVZQDw1gtDjKgoLFD83uwV+3mF5LqARlIEDzFRSMng1dC/18+sSGciNBA
FuR0wYN/UA6R0STb7QheI0uDzh1Pu/1DKvgy6um2JoSVjU/7hibPrr/I7QN4y1fD
Ha1OYffS8xH2U/RPFzCLotQbDdinxeDc231YiD4029xxWc7s2O6Zuhq+SyiZZT1v
yT6u/478rhPN3KRtKeDi58yUHrYnPGmWfC8eEy06PJy8fMP77N7kkhCiM9dFr6cR
uQ6Z+wMewxHLdbYRd83AWMTAU2OJDPYD6vVpj9hsKzHkFMVmCVhsJO4302Df78t/
wn2ipyuySUu6wyIRyJJGEecDjSzyqJA/RWs32edJ3sR/ZZXJ1ebp/NksMAnOtWt3
DoEZjzS5tBY0+ppI7DgkA9bfIs3B7HwVqFkC1wzhL/FXTKS4kdBrpV4EmrGI5jzI
/f3SbIyFB5Tv3jYYxR1ygpsNjpLvKehlsY4A9yoaYAH151wYqGB/O7+Fso/F6vyu
cWkKd3SyCVCHfgUeXUiPFK6w/xyEBXAoJWYOwKTm38ZMkAKn43MxsnjBvjA2wT4O
IVuaUUhEYKCVR7cDFVfEFyfIjD/8O5CgOoicLJSoDc1uOvCzPEr623VHm7Gg3y78
jSFz8nbjt0X1y9J7lZhDDDOsM9F2eikQu+zf2dkeD6aIhjZjGRDXFg+iJRl9MqCt
F5nOaML8oNS4r3UJCr/T8ENBH7Ny5jNi389aaSy+nMVqqADGVu2dlEaJbNciXiKM
8/jcJMWjIi861Rs1/bohMIEKVyE5L831Y49zmqZxsCjSYpAuYxfkVFz1SGjkDUpY
JIVUBOw7Tw0uunyfbDcEVAhv9QYGAFr6sOrS+84kRAhc3dAYpiWoOndDfj9lxwBy
qoVDCcgGTPwqZnYRL72CA9xu9qVOKlxydcmyYyb3w9UYyZBG/J7DDnPG2Gm9FLjY
/5SgNwgrDPCHFLjb5FX/PSOq8CWgF2RDjOfc+FCy2aw3t3WBowyJ+d5YQvBk/nG0
RPSAqO60a1bSYndl3rSLO59/0tkRVPMluBkKckChPPqXloCUlxu0HMIbVzyZEP3w
q1cSU2U0SbWmU2J6q4pdAgbjDSMQcnqA8BeJJNoUqTqA93szLGdFn/awzNWRLdGd
2Vb+vaHU6eQsKCNLUuiQ/r0/ZRGyEzVFojD4VpFYDsCAYUsh/s/lsZL3qUtq06Xd
3Ie+gpwnSUjLnUz7oD8E4nBcPfTVRaMuO9KdKheBn4jdIQc4GiYGd+MTpPCnq5Sh
L/z5YWs67kwD/l5sb8YhylbWiayTiuCEkFhaggCmPm8bMjiqTHucyA5A2u75UK/E
t+3S7DxLhoK6CLKmqnbRmj1qEN/JPyY1wN3ifpuZdH0hJlnDObMF78DGqo9dXSgu
P9ufQlL+e0Qk0dI8da0o1q4KWnOWeYxWwaSniMQAjOilM0DLOzdR06b4x/KgJ4mC
BLlLYdO363QE3SFIdLz96KolqO5Ef6M9kyzA8aQtzsX3b3a1pgjLMy0mHxkIZgEF
tW+nyuiYaelxIjzAcZhO4/EaA4cWUVHOPBV4YrWIdevuD05gTTd/PdxPkt4SUdCb
hb826h5UgltvZpPiOPU7ljh3YryulZO8Ev1mjiZQnf9p6OSc4YkakmuKVBbaspuz
toFyUo4uiurUtEScrby6NFiYgiOeVbem13W868vk9BKRS2DU+ri+aryt/7Elc5mW
oWU6Xa/Lzl4o+rBvuDFiBfpKzYHUk17cvW/PcpXbl9PfV/KIdTtG6kXrK7DIg3YW
UUPWFIbS/p0Q0XD6fbvyQooWcumrTfHjxdj6Bf97IEf6wies/UkDC6cs8Ol/aR5Q
K/8XjkiViHO0H+V4plUiuiMetoRCymdRIm1TJYKKPfBtZ6h0pMYIJLmzNLpuWMOU
iFPF+xaWc/1URUeLVNrJ45GPv9vpW12HcffaQ3FpDrh7CnGp2BDv0rdetAxfhI8e
9Jhimax6hwIlQJ3+NnkQ5YSRTH6rQ8PYpeaJxj6QRBqu2ao2SvrLhr4V4sv6XMLi
41EPrr4tpUEgWnrfYeoLN1M91x4D+gDJ0fACLk0jF+DSdwVzPsqe4nDtZEuHLnqH
nkw+qzcA3UGhMzl+a6Tyg9hbvfNug+NHZ02WpXD2FDkD4SBPHmTBBo9Cnqx38HD4
qCsQj1vwqar3XKAZasJ4UULfJsshfRzKV52pAfvqpOmkX2bZajXSDSuU+Te/yHwW
6PXQ7wzok/WcxFCYdMXRj+vPeqrB6VzDW76wDD2BduFtpU6IaALX1diVngprhN7v
nagR8dHlGDlkkP+VuTG74nXOC7n0MtU/T187qnyliCZsXd7UIp9A8HIp4mv1l14/
vhRDzaEI7Cux8RkZuakxmwSRmvSHOGbRvYa2Mg8nbUqY8b48vXZ1wBOjpmbIoKmf
MR5mSXMtSwiiLmKR/Chm434sBrJm6+hkjBowK1vSULjq4/dUG1SA6Vv+CyOMI2Sn
T37kHt/nplZQsM5y5YgeiS4xatNfzwziVO8+aNdEO2rtFnoVL1ruDFl5SuwxNsO6
zKuIlkqm0GRngo1d2+ThYIlbrpiodYb5GxCk8Bw4p5IRy5SidYI7ZxCDzB2J0wjL
bsenQAx6MSLMAqFerruptuqYTAwBRwgyNaUdQEStMfVqQngBul/sbBGZfOtjKDdp
XghLKR0idWV5V6coXaC3w0ns927uMt12Xk0xNTvLlz3KemKXT1xTI9D0R83hVBhT
jDL5a5S3Grj577RtButq3TvsKIBQ2zgYczbhIvQ4vTMQdZ7WK37FqyYkUP7n2arv
crRs2XqXq/6mhveTwkndljetF+IrEyyFMqAVjtSrCOLChAe6a7Vnn3NyaquiuJf/
ujh7hcWKJcqZiKNYrRxvsPS0otfh66H7r3lG2fsd4GXmLZ18FXa54ykx2gzgvvfk
MrlDtnvI0lubOSUW/Py0Z9h6flS7j7S8+ggHdLIdBNUiWIUTTy1qn+xLSqKMKg/u
3zq6vA33IiN8rWsDqztbgcVIntEaSFMmxM1LH0bzlYntTh5M6bGK9OiP3vCuHTya
TvCGhlGClQogH+M4pONeYZ8LyqnHWQ2WBnMAmua3bx9r3pOWOFjZY6m1QPKTkcUr
aVjZ31HJ+GtMtGekOaLRVhZLXHdLiiJB7eW0XfT42Fs2C6s9smpYwvJCc0rTwU50
sta6w2XtbWirO4Z+LeKSSWjG8iBk6qiM0+OIyilxg1WJWShHoymuI+rFY2FUQnut
UMaG8wSp1tQ7pERZWQtBAD1EmY8WquUspZ0Z8vrsvWPmTaoyFnNuZjM243uNirgk
emKdwTbODlBf1ow2ow/qb/OsWRgjNXn4vHyP0aodiwR18mS29hg+W/gmze7lip6v
8SBEFPY4XanzGxPCEb+tAE2C6sU/rAuqEhBNDfoDMGACLIw2U8o8sDNydDRAHOT8
iTxzdPGrXZzAh42+Q6NEA2BCD9PbVpqMWySXD+snO3Sc0gf1ufpRO/iuhHL5PpsC
2mozg+BU8/q2QqGu0c4qlUyUrTVjMMjOcrtqIkQFfCPhJaZei8We2TTesFpmuUzK
4pHDvE9JEeImnrrZ1JxInqVXEER5RMkGYP/nG26201Rf1sRoQhZBxkjxklrtThEj
ffva3vaJQ8SZOlgf2DgZIPfn5i70m+Grci7MD8LgZF1yU+LT7uJC3mDpOjuuWI8a
IJYglhPUPZDEF8WiWJZx4J8G7QZe+TUCD8TJvFaM0X5ej0jtcC68k24ijpJVVEeZ
4G71/tf+24aa6+MUnLMnXkFF+f+EFR3XUAGrFGOJ8gKGYsNHi7ZyMZ9GNCjI+8+9
L5LtWZKGPDufgj1DD9NgfD1qz+76aebklqib3pg0Um5S1S6c7ELCNg39NH2/BUJM
6521hASSrUfO1utRJsbPZ6jA8mnOd2CKQe+B0VoZW3l2G8qhlm7XhFJjClHnbFhD
H83UMLzdo+++fVw5v43izE6+uDfBrItNcwKFckvvIp0ZlvGM73MNF823YyyGTBaa
P0Ge2ddozdXxzTionyc4Y4rnJqLsH14dXwAKrLlzMIWTv00Vz0djN/U28pFomQdz
AIQiTxSo90/H72OjpYwGEmXZV8UVgPezi/ZQ0ZbMNaLLG8Ra6M1wf21wmd8rxhmG
rUnPxaqErWbTjpLT7QH6Njs6PeWvhg4SIlhoSNT1Dzq6OCLPV7dz20DU9sWQv+oi
f3wztyZKQldkPcYOH0CaCfDgi8+1GCQNJT12DCHq++gBMW2tzIlRezd3Ri3T4z63
1Dr1TjdY0GEw5F+bgxc7qBHwnZ8grvWORkQJg7w/q1LWJCTojH9fg26Bx/vExbe5
Xq7hZIDiHtO3Te7HJbVDiNduEWzmKo1aoSFQwHZVSUt0UtN1BKcc6Ydr+9Pz/xro
gBBsiqUmWYVcWtf7jMxQLF1TteX5VUxYe+2kVnfrsYckiZJ+iGowSPu00pWqLfRk
yvT1d3yBCdyt7c5pdLfJiHLnmyySSmpO7S7OqM4aCvPWiB9a1kddDlp7pDoH/Qnw
WVYHLvvfVcV58zjKyCNxyL5CfQrZfGeQVE4/cgA4jHM3V2RQ9iOCtW2Uyy8pbea+
bFmxJp+2cfutnYqzgDd4J7WAn61rimYdktDTK0qOVkAzO9oMhS1oHYy7jqyl9GaF
/M5f1HB7whrVvrt/9AiLdt+HUdIlsHlZ/Z3pjOukCoV7Om6It88gBS4wWeI7TUdR
/qHGv5vTObzeHRH8qYZwr9ZPXkNq8oYvHKkRWRM96sfNilv1ss1kEmRs58u3Th+o
K0vbQxq6WIYCsLpRlh/Uo0ebck0XV8VtdelQL7ZqVDwHT+h6tRexzQ2cnLCSkBRx
9H5o6WxxIGW43g4dovxdRi7rpT8uwdAAVTUXym21bQocxmn5WHxzyUt+kWuz6EMl
eJdH9ArlsvkdWXJLaE6v1YKyALgP3VzQar1GzW+74LowQVMZxmfze6JpYkwKFClt
StRiY6SpwN9OejO2qWoPmFKAaHUvhp4wa3JnHMf+zYA2np3VxfCTOi4q7I9zh5vs
sFBZIzONkqGsolhJMzue9I1XMLeU7gbi/cktNu2mn7IfXPdZloixcc/hKljSfqcU
Grrm+pZaxDT7AE6hMKDBqnotHDxGFbPVwcrTHqWCTU38HJMr4Qc6rQQ9CKh/kjgB
7Ww9UKBN0I5svpY5PQxUiAVLgiLBqF+i7ojeJw6ER9dV086ePEXMmEtALWDStn2d
r6dRcXlXFRqfPKwLpk0Yrk93kiNECR4FfD9csET1TAA2cqSTupU3O3fzq2M2IHMm
orgGSAA4opNa+dSZygG2TNDg+Kgqf5QseG3U8fcn1CLnKxQ2K/4Fjyq5Yz+KBXiL
M3Jds4Mr6tmHBH3qMLXIAHwGwQ2BjwMhsvQzqQpQy7sdIL6GVSlIqZlwr22MIOyg
Yz/KFEtPV4yWVaNri1Do3MpGuB9t2n1H7+ccSU1AAWZnkNObV7xn4kw3dJ9zTPdy
w7EI4aAlRr12MWzmyv5kWiZ/o+1ZpAt50y9eeoJt0+fz+Hr7yukykANY0b4vWa1C
xx/Dr4EAw6O0oD3nYCYq1fWp3ZnZeMegx8dNQ2XWovr2Nha1afBORye76t2uwasW
JvTmhzxGsxFaIg1fz+GaeEdxGxg1aXG4xqL5dMSx2S6vjLu8ZbbYW1uiflHFzpqv
JdNcaXyJOCwF3KENo0NIiQdvDERIutijwCMZvzkGXEmMS+zqXZTYJvyUVT1G8dnR
tsPKu4WooY1iFcz4ee3Z9RhH238whtkP6gD+F1vTT8zm5OsyLauwLfvH3/Akl4iy
hQxkFjQH9PjNXHkiZvMMNliG6E+qBzt9q92pmSPdC4FL05pxEwF8Qi7/B03CLG8E
8RM6iNwcB1DHJheqjE1zjh2fvEMPodCuXgPY68QvuwRGIW7Gw2IjxrxhduOBalwG
c22dUEtkyGQdp5ZTB4YrxEtZ0eO2aEfyAkUwvpDJYRHBkwWwFxUNytwC1xsBn/r2
VgB4HlFNSSkxNExMVrCJSKTGP/nwlw1FxPbrRQxajpl4Fx8dfghz9EdEbiGVDR+8
ns69sYDVjXeXSdVlLxikRNW5Bz6pZ8yeEL3YRxM7QT6e8Zycw69XQUIZYVIlRhs2
BmHaHA84JWcSEoPQOvQWP+LXHvR/3mKqQACYc0ig15vtR3/lDomiOiJ7mcmwiMNQ
TkeqPQHGIrSlYCe8abgbNq1I4mGVtmvb+bSb5yzG6UteMdzJolAAdy91lJYQbca8
ukcZ9Sah08ET6q6BiJOmaG4XaAkwV3YD+rBdpTGl3LKyS7nc6c+DYSIlvX/OcF2M
kcgiIYd6odxCN2h++Ehnd0b9ups9Kqx0WkMzEp9MWmHL64AmgMd5wxgxRprtGwtw
G1thDnF5YcmlUMZWST+9cW8BcwFEH0JyrgEj/lAyAyPQjDq67W0ELB9HkJ1aat0G
ypht8HEA0bX4X6NtCu1ROeWd1X3ikiG6hJvZ9lXRrOxi+xIdYUFHwkKs/YsFUX75
c88NWJhWTGUMC3n530naEY7UA5xE6zh1h5o2n4VANNC5EuoOBD0mAzRLp+Q+xOhC
HNEqmDEVuiuzqL6i2wrZpif0UsrSK1Nb5oxQM0NkO6UWuDt4zXcEjBbZxdufPpI8
A9zOUxO+rf00whMEb+Eu34Sz8UwAIqGRjIGMLtgzteNr13BInBNMkxPw4FMLpYCp
o0fsTpGXN7OK3+DP9ZUiRa/mt0dW2uYK1iLkh/nZi2guX7rXOCqVH/p70pYmkY5r
ZN9Ym8tHDI7x2nTfU40pAXpKspDTFYlH0Bt04rbGiI6gVgsrmZp5w00lWYuD/GEc
bWYhSbloOatUS1yatPQ1hp61BipTQPgBU/U/c1zBqvyhKd1g5XQYsGSGsfwUmsyX
jETMPjCG8MzoHXWHXRowtj9x1MxLmMCh8oZEEcuApHJrrnj0nXBiw0zNDf6ImaW5
ndH3r3QT1JQcz9Cw5qNL72QoFEp+8oqsAretULSqZoaLKsM972KHtN0eJIAmiDik
ZoHqs7L71sm8bVZHYqvH6KZZRTSe1ss/Av35FnepMpqTm4BbRwqy1BdqgRndzZM6
9C4pBQziIfelPzrZqtKqsJKyr3E6bV4VktCYhY3JP+cDvutIRv3PSkvLVZoonb09
mqA0zV7wbH9wOf+zX0Lwz+TVDib6XRegTTUuRzdXFFvCUx+p+ndj/Ms0IjEbsxiL
znWBswJwsZKR2J8tcrwyrzoXqiVj+NW20erL8PcCFvb7sDJJWHM9ZZuNDlkeiJ5r
CKOQFaA8OnCiFZWe0iTQ6Gt3xe/d5W1byP6x6ddGWxTzTL5hHAqrCcby0B5kFuo4
fKKRsGTlaQD3paRDptwz3K9ZuIig1o5semtfzARRnZJ8GkgRPf07tIFqO2DmzdAy
WvibjPW8TDRxsvzWsCEMsGxC7opDYuGMFJyPaJMijacxeO9Nd+kott+QuthfdMR6
HlR71ibgLeouv2TVnCn0ZeyOMRmP3HZnQg8qPxR+HWSlJffT+rVnlw9POYU5d/F8
0jsUXo76DxzF7xMItnZp1/vP4JS+Y8SmZU1H9vlozrcpefmMDnYtD+H5htEIvKcr
4wh3pM42j/b5GbSqgHrj2/q2u49xwVSjfgSlVkDAdFDs2pcOtES4iY/xTQGv2alD
q/R6sqs1OgQ/v1kBKBEzinnUMMy4pPpW9zzQtjuHarmzatWpgw/AmqpImYzDFva4
qlhLNvQ3yV55YMvUF5Hk6LUAmb1OM68pvMYjqZT6+r1cs/vUql7k4dJxCTkccbTn
Ocnj07gSNdfFmq09i2W3MA3jWVQ2BLC4uIig4iXH2H/yaJdPsvyLNQEptl6WU9aa
LUvWiQ46wJikeIoVoPfO5zbo66cvQV3SzJ70cQrFXzjsFQCVoH7Sk796mwstcahN
CmSn4ArG2svR+HsU1ER9VXbvyoK/iXqi3M+Op3kc5FZrpWhJa+czv0QN+HyOeV9v
Qi0Byo7ZlZhSAeBjycsgtBujqTi5PZhiCtZ62Ke53024QKWFkInyTeyCKLbmAXa+
E1/BDL+c2q/14qGPURQGTIBGXO+2onDiO+RJ5EA4xo+1gh19j6XxR7+UwIK1GAnJ
2kjVthNC7D3oAYHJqkB5l6eap5RgLieFWAjpBk2gjyFMKSHn2aw0p7/C60SVojrf
fsh+D/YPdBHx51C64bzoiWW+eVSloonLYQkYTBKm6vjD63AgZ9Zrik1VKorYr5hg
b05wruEKAWM7+bXG94FLqsF/ZZlEKSaxsGRGZxegHwLyGyWZj+mt7+fkjgTVKRMz
M9fbeeTDgg5XxP5qPp9AZd8eepXOWXqUVfxE0hPex3iKw8G8l+PzhqoPqrFvekSu
48XzGc3C/0rNeqKa8M/UzpWrT5jY0nDWrasunVfg0SZBlFP5STFtKHOMFu5ledST
fSwgIBOYyeYKJdLJUP4gjrQ59GCihTCFoqpLyf1nZ8iccJWMHb5pUqn6L7i5sKbW
vmQTjOTkfsOibn/Od5nv51S5L7W2WMtvLeYVDHgl0OaT2s8/4Q2KAmP7vdNHGgbe
KnTz/yQXgKJ6YerlyMHvsx8ffNM0TP48rZ63q+4NWBM6eyCeNpoOJ3ksCAkF2JuP
0OYHYDNwuW6Xjd5d6tgR2gC/TZJVkum+pHDEGmRedcDRBOC068YDPB/h1BiaphTA
5j70vOvNCDYHVlP19Em6cGGCXLj16FSFSsyZpUxKRwvMBoy5yGQqZL5kC5SIXTpT
35v7EiWELn/ANQZQFCnO72rqMs1t29WBrt5wlSjXMzeBzV+5Ix/m0Ixb2hhPQ1Vr
IiDhCbpqlcJIILB7jR0GgjdbydcHTbzi1wFYW0cLs0JiYv+4e3rvRCDHrZz3M3Vj
U0uwLqMTEOn5WC2jNs9wjJ4GQ7hRxv1iXSIPeXYYf4T2DD1hewP33OYi/QA+6TMW
oJ7H7mvCdDRqP6bDJUqJO+1jsjZFuFwb/3v4+th8aYi45M4is5ykA7NYKsCjpOaV
x2/FsWBl4WC9lKFD3z58YIXPpnFP8thUzi7hSU7pFaFUKWT78TKVbKBBr2Pza+8b
lj63T1gFF1W7AlCD7RboP18QZdEcLOsUlNuq65QWkVV8I3cSUCN5nafK7jotaXu4
wVMVZl6WfCxmIJUUq1RicInmWZ7p5mqukgDYIXeH9H4ninpBgBxysnSkceKGAlhJ
yXUETe1fv5RFisNo9dNQTWY45iFBjdZFuEs6qatWuC7jzEcHBmLZ7m3hH4DcKf5+
hDpNS+grbQd5joU5elugCTXAdGCQQ469HgRMjknRt/oXwE4KVa7lQTGOC/JJ4rgC
xx52gW8g62bNx/zKJMguE3P/oWs3LZWs6qJ13ztOZC2iG7SkC0aIlyXinRwHvPFc
NzqMjKtJSQRMqK19f6extPqsvrHB+LPlqmij/Ehx+NT5a1Fuyu9AU55xPsCR0+SF
NNyPwCak5ZDzTk6FY6lEkipoeu/xbx315vD2cPJcvccgzqQhYFpHF1QUZpJXiX/F
3lwvuNssoTjPOr3FCrOdKQVnBHJ4G1F+BrldGJb4g/wyPcSbR3b4zBlMfUxOpQLF
OZWbQYBuo30zStVSW0zdFZ5kjE7RBOolbWfiz8LhAgvEb6JV00Ujm4wb+XZmMP5K
zto0S1VyLy9i72HIEHyM+snORvimL2sDJ3AR9HBxuT0Gg+tLIFIaRhmhE1lVOUEq
ypdxFQbVrz6fa8kGKu0wyyd8qpwEW9164vyQ1egQIbCa9GUKMGYG39lqTzeTlERp
Dua/yL17qraKJ3+kNt4T0xecz1ON9ziupw8FujTmKdU8jChVFHWHlVURCwEhAHJS
/8jpS8rFp3Gi9qmov0OnNztIQ1HueEd4zzlyKoMeQ5Z3rkQpAUKDS8+FK/mP2Ymt
NiTCvXo7h2DGWv9jKvchvqVfru+VCPLhHRiMxTD0EwqzPOgdWRMOnRXJrJBFnFRS
/AkBKcvB2V0v55wzlXXHYscFAC/Jbua+mqNQLpQJKlGXptD9XbwdMZCuslGcYywV
uq8mpGvsMUImPIEd8VLfpxIg/2Byy0E6o1Ik0+miN9TJwILLktYHbfcpAZuj7Odh
dPHKVXHegIPPe+PpP0ZmoDDiVvrKSka6rGeq5bLVUdy3NkbStEGrMRWXKbqr7Oj7
vqSKndH2yUoHUsD3DOw6B26sS5RRq+8Tgat2OIMCNv2btazv2/3/16cBtTmGQ5La
GBVE5X9dD0xOxAZiU6CCja1w+oVcI3RgJO0Rqp+0L7AHO7uwXArYYnSClwv6PMch
vufxC3Ecrw8BpNRs4jMzzC9FLsr45F0+i2cRNPEr/VlHllJ7u2EKfj7uEy410KGT
/cJS4/JQAaSgIKEAJnuZP9An4gddb1p5qpfRvnBuV4Rop5BpZirCdUafi+JKz5sl
JLs9bve+wv6eYO4SJk7n9orNCf8PVcIZFWp8fidNSw8RcJytN3dtxtxJ1mVlDhpy
5OUmn2TIq5AUYuJyxCOIAo8DC8oG912fAr5DiVZK+yRLcMKg3yiopn4BGrrAw8jC
sxdaoKg+8rs/Y5FjXo0WsJykBizCAZac3CSNGj/mJszsUZtNcCfmErxyS57vu9AO
uhw65lWq0OiIv7gIF2YXQDiL8nzJNyL/wgXmgKSwx3fzbYHFjEGiesICPz0R9YWG
JwlJbMkP6D2Q0qilyKqxLh8FKol5PD9ePh1EjfMYAKv2FP3EstDQ6AAcChXrcWKs
AhSoc77ItmJgEmT6g/Lh8O9QdEV3WgjNZtVZOqXcNxOw1Yp4z8/qXszRCh/jcPwe
nmkRV9E521Q0IwsNtULcmklsqEUWuo+zbaIHVe79v4YJqTe64fLbb2mrXFtDzOvE
LEZ5c0h8JLaQbdPTFvTBFf3qDeapHtFp9Km/kAPh0XnVKGwJZiVJS8Y4PKfXiAa9
cXfu+EJDBDMjrddx+7v1tx2QFSzmFvpKuK44PegRjCq+7abGNbd0M+SSp+fsI4qu
v4w/HZdExuQsUFvnlKqWT275q5K9T9HiK2OF/mQjBhqlcbXl5TEzbAKiOcoirjFG
xVGSp/eC32/yxdSg+0xAFsThtAozuo+rO987+XFnMRoksCyPNWIjKXswRs3OqOft
/6xMioI/bkIDR0isnG/l/Dd9Bz5penIDL8a+AbSt6fm5hjUIgfYynCyMCF2AiXPQ
j/2eorCUfl4Cn3b/6F5Ai9THtkJswZE4vyEO2VkYCMOQAVg6Id68eVJSpQrOS92x
eZr9PX3UDRSHPJgQ85Qf+Hx7jr62bG6gvM5HXtYdpMi1sZtlShXw2OvV1gVoUF40
9GMsEU12et+jGpVw6Xfjp9sTLp71nBp8EPNtyKGpz8Thqy+usd8cpCtJkPk35e+o
Cdw2QMFtVQFd/eOF3s3gH5HPsqk78ZoExavCtzJzszN2WauLl7P2XkNqpZpmOdOr
l/RSQuXhBNsPudK7DL80EnH+qJuMRo841A1Lxa+POJFOYg1210EOOMjqkOS/nyRv
MazfiJ4B9HGqxFm90aGt3Tm34VnYBWlhXkjVY+/LMpHKTUO5KBiel2LFf6fgCxEv
KUCSaMWJE12s91xLN4+udZO8VOGuY0sdOzdfqoXHSlaEZ3819OVBhwXN2rLuqZKV
jaytKIzVDZXC9vJ2aLbGgz/trODYJMg4LOM5L5EuiJ+y+RPeNFEVTYSCAE6PijQs
dpf1LajKbpCuPJtnEaxw1LgKOI5a/0D9AKSjgtrUjEo9bn8Qk9eC7XwrkNzAt+Jo
Vwr+nwruC87J7kJvVoEAsyNTELj94YAkEOWeK8RprxBXZqjgTlTRHvWnMJ59aLYP
6BueIufFURU1ppdplUOWKuXsV5EhbFhymlnlbENl8aoOSKGBQ/z53u0BwiYnXbh1
rJgmVpc6mf1DiVe8QImUs3oxdjzUZfemsFMPCmoBLeHWbinUapGIyWt54YDiy7a7
0rFEpTX5lpxSe7MT4D/NpwD4w4Yqj78Rh/PHb+r1NfPhHBdWlS4T34HrGyQnHLdU
EpSO9/8jumB5urie4eYhnvAumcyA0kcgS5QRu+7zqu8xd1Dy+wM6aYjhO400CsDQ
lDLWjHzZTDY07YBuWAcFYUna4xPZlTxC5kahZCiU9XDiv+6zwna4DTKF/kKqZSko
5Y2ftivB0LWr2Bw1MO3tkKK5/+C3I9EnuL9Um2ST/0SQE338SGELyTZBGeh49Ffn
Mq0BbiEfucXbtAWl7l0SwM/F51wD7G5DyxL09CPUkyik98lwufY7O8Sfi4X0Zj58
5zLRzgiRKdgmVOTMZC+goXX+nbGLcdmEJKxwBwuJJQZGc59r+4F5MkiHfcVirZg5
lEEalGT+w5tjE9J8tGPQ66+18BCGTC+lYU8rjbFG5z6vXRgrJKyQWl5O8jtzPFKz
dnY+RmJHJurjcHnHMlbudVc02Uv6Ly8AgFrfcmNUULE2HTSRY8HwWeHDtEhFUU+Z
pUIvs8WbBJIWxmodH3Xhbl8Ek4GAI53d39allyppry3wBJsryqy5bBDqMnE6Vq6H
UFHJ1GkYjZnSy+3FYDzAtLJmUZZ3wMzOw1FOPNzqR9zfCSWkSTMtACneVAaJvEI6
5/8TGaQ8d0Q0BVg8xe8heFKWrOQ4gJ+j4KZj9sJFpWlZ4wzQzTW1Z3RSThUz7U+X
sT7KHda4ej6rZ380rbNgS9EryTWYH46RJ+Y55gmd+1Ds3BY7+50+unTPMhL1YZ7N
qYS9LXwMceII24zVk0IpBrfg4UWTFhH+V3r3wJBSqWQLudN8gpCXNvgYWjbH1YYZ
wV0/pE4T6MYtgEA69GHRB+T08x71O1kp6qSCZZXBAFFDruUiFlUH4VUsUZPgaH+G
KMmQOY559KyyRUQ09hRZv0Qwq1abRkor5hJHFiYXKdq2tzhHZQ/Kg0fR6XUGnf6x
yLTiiqyLnc+T/x/oZr+JfUMRr7CFtU8eBJcIj6LPiCCb55r8/ixjVdCID4gis0Vp
BgvXFJejKF1riFFWkMoNwbMVaSA2F053M61G+XhmRlQMleGpgsR+bGqvNyn36ZeD
24xYVcrT0oJIJqdsxssfekwGgUxfNeCxG/9D3qJevJuG46wxTtpH4jlBVS2CQ73H
V07tH0zM/dDIHTdynoVozK/5Uk0RZgjZND/9gON9tsdiJ9tf/05hj+Mskw7MwIkI
JHcfUWwTaNI8mEh6O+YDwQkTrz1/8oFm2/6/r+TElHAMGPvpMLUIFC9IwXCNsQcO
/mpYPF+owS+qy1IXATHv9L0d4B+Zn0l/UZrk0uHUv2WZDyU70hhKIr5MoOVPLl1U
rcLqwsY9K2/QOhYLGrvHRZwMmf0QUKLLuORz1h3Az3H1/aJSgDCEmwrU1N+3QmEN
CmY8a8dnYY5p/wJyLiLktYzf7l7AVneX0mJdlaNKtNIzuha3/qrnLLUYlBp7ICUM
R4l8sUbiNfY2hoh+0GRBJP7cFn/p/9LmcV8EmcT/FGqCLk0upjePgp+kWC9JCONb
SXxGQMKN5T6P9/rllPo+OuXHWkZYEDddVZpZQH3FuDgm8vNSslVTy2AVHesj4M3q
G9z/2mzkvHOKMNvKkhN8MuZjmXT6yGV4FFQhxlv6YEZYHJuR5K6lxKCw22epV0kg
r8VZH9XQrWh7QHpTWKMh2IxHmqrUIi6MFJsRn+bufnIKrwwQ4B7wYmI15ErBW40b
MpBmqGwxhO6hSQ9VIITN5Xp2UWyn1w15eeuRgQYss7iOetWTIxZpfvE1+E1BXKty
gizW4OMwHrkq3KdqBbpzxCkVjcSMGSPBBT3KxT94jYdzPtkkGtc/5LA8wkmzT+yC
Q6C+xTR4QRMV/gbILk81/vdfZ010Sa7ktzDvsOBRypjsnEW1lNGMpNUMUu5GGpNK
nr03WCOjcjueBTGTHFCmv35WtPSIssIkbissMaHYlbXH/s2+6nWN+v9/V9NZNB/W
sXvxa/cLfvgqRcMmJw+L/mhF1VVHhfKhbggUbJnthILSca/BOzkD+19W2n8gl/g7
al01RR8PL+btut2Fpfy1tRKhZLtvK6uCDgbIiUgZ7KLkYsETFKTHqUSUUwCE37c7
38NmGcV6qqr+b/gcW0lmV8oL6Rmzhi4xzWBuy/SyWUV/xHyeLMz1y0UTXLE7RvW0
8V4b6DXTU0D6fA84dTHTB0D8AwE8clZCPVPsChQKwDexeb3yOHu6BpPfXEuIGHhJ
YS7zwfhJjz4zHL80gcOzUqaxhUzGsKQ8EEpouPvBXTaahZzanK2CKQd6J+ds1CqE
2H9XXFugjiK0Tx6XRz3hiMm8w8ZYXa7V8BDBvYnZdeI23fEnfcNlR5KmdzOyKlWd
L5CtN0MAM20IkQnMqppyqNry2jx/wHxC8jXNivU+1kcWUcMoMeCSGTsxQaLfxZ5B
UX8qfRrIsMyHXiNCo+yv1/9doXV7KLgyP4UqlxLZO/c/OtH22X/ODE3CZKObM9/p
ilEWwg6VE+b6Phq4KDgLrzV6k8DERRs3D1O/D8ppRMYSvqDGGu3zBL8SBW598MKj
JYQC9/Z6UfuxCLETRAPM3pennLNP1myTjZtIgAFZADEYXau2kL5NgZdTvoeeaWdK
irAqCkhIOkR0pxbSuDJBky3MyXB4SkMjas2D+FI5/mjkS1s7BVeEuW34MarAZpsx
zjFVZ89OkWeh4NjiHskfWFMQuyLFA/aBzAzwFPOaWDRKcGmuhjlsH2XORPp+j/h3
0K/ds/4wayWkkAmoD7aBFN6+qlgsuCzzj3TpDjDxMLZLQQuitwpg1Zj9lSvl4K68
Qo+QbGQOv4u+xZuA/FqtBoGvkBJhuvJ4UUw+F23RWdFJq2Sx4gsAxZg1Hc1E5zfY
alWs2j3J185R10juKefTLl9xaQdKQchnvFgsihNm0NOKfzmogHdogNBrGFrYq//g
xVG8pOm99Ma1UM4BUFlA8re1u4+og8N65sbSlkUPDKuRk6ILu8GAzBh6ImDoIkHS
2ed4KUZ0DhXDa4s55fVpMdXCJqPpEc3iqzZ9Kinw++OevWanhSRyMLtPqw04fI7S
evVfsCa84Wpe3qGLO2Tsaw3Q7fGttLrzqdh+owmE3czaNR1tVexdtWBXYB+KYcB9
8vQj7Gtz4fui+sV3VWMavzjGBXbIARkM6vr9cAsE6jkpLwXz9c8zFIqCr6Kvwb69
AMO4NC4DYxKyTIrazNDiCiYGxfilsbIHDl2MPhJKXGkNXxCBrNnM+7jCIlQrHTBr
hJ+3N+0l3Hb87s2uFrmawPJJzRjKZJ4Z6ILzmKcgJZkGa519z9htjcUUPBd8LcJ1
ToEF1uYCCcWjkFGMlzsds4lAMkvb0SphGqdDbzkSInGib/WtP3UaESsj+Mm+tcRs
6+aiyI2bbvW8eN1sAqpd8gTCoYH0jELjXVOYSzgKX2/MIHp+ZVT8cnOfjkCAp4SK
vuhiVJu00HI50IOyyS0GN5Ncr+GiVaMgyuxEz8HveBKA0meevCtBR8Pk3V6EhwRp
EPynTIPAsWHF2zC3BPOhCWrTNoZ1h2rhFhADwp4aRFFyzQ70Jd6Cy3XCorSbeuoP
xKSdJ49TViU+goEGLqqhSHVxmar6r7o3r0MCjE8l70TI2iveQGZVftqXOBv6JK2R
UOsIdcp3Ea34ALQz2HLKpSSZfHVH+g4oD89vIZyrN7IHvmo7bmINRVYHGmNJMb+W
w4/YHiMpL9vfr4CUpd08I5gstMcDfZfWyJjAp3vFDYrPEsJTDXayhU+i5/lnPwp/
YLnnpUJAX+/ysS/TkbBsjPmM8mYUDu5uNRaBThCB3eZ730WfQdTn5aVs/xYNr5PA
N16IEPNXf6MFJrK5d5nXmGRHrSz4s3cpGZm7OWAbQmCiisr8B1csDq+vfV4GUoi0
3KarAf3GElOK+Km144KhQpqwGmxbod9eywaAEDN7lOdMG1dPbMSbb/PNudMZbh2m
WC821u82uihvRRXIhRef6tWGBgz7nVkCcCGNvCbg83LBXOEiu/yxMX4aJcQxIkuV
l+n25gBl2l1zEY3L3FlGVb+JGhFzePD6d3UBFoM6Wv5dzLEnP0kk7ccKqyZ+ciED
CuHnAEQMXHKsfCMf7ToXTWN2kbiGDgTRhSC5dw+y4Qb3Vq0nG5GGehJG4NYkw3gs
CMLpmDDU4/PFfxV2sBpxhPx54X550Z/OVUQPPI4wvlrOG+yG1t5foK40K+laDqQt
aNB0WcIgQv3qCCGxLcOxqYG+BXYRwUc1cYCp9egO3R2eKj4zNuXgpl4kVyPLNxEM
SsUp0lqY4KP05JtdTU6PmWa46Vs6nFolJEduvO7mvnBw1wWzenDtjcoQRZhbPGNB
SVCrzevy1+e9kGh5xIBSpL5d5VBY9Hw98dqXulbBWhyfDKENwecp+okLxXIksbN/
q2OSYvoii7J+C30knTZe5Mtt+yjIZotYZIa9GeOZVuSPf/52Un5E/PhIqLRuo1S3
v7Q9z/QvcRLP5CxE+yXEdRnbxiw9MuAUy4GdXbKJV2vR3eOCN0cC5dVxGiTSwHBK
N5FAPscucouM/tMU+tYgLyJJJFeutNEOnv8JUR1gsAcbSrAqRs+2tn34bnBcUMk/
5ugjKzb2ma/h5kGo3TT4ZO0ljXtb3lEy/OkLEYz1vCu0RUqrueIdmGPZsdy45vsY
ABWSRbIXtTZXYaNnFIzwDFBk5aJnyAwLrrtAFFkxiZYqXUL6KJqs1a/OnXxzGbjj
8KiRlOqWDn8hk8cIJrp3erlY/4GO13E4A35ll2o9pJGvTDcIvTAlUMiDYftO4zzg
vOMCZVkle1McsR7hz6PYSBk5x3mj39Og/ds2u6qbbCe5hF+aoiMGiLecy9kTI2qu
Hk/CLaPAPZEd1SiZ/4d0TreWJ5AyLWzOIaDK9QYqVgGhw0TBg4Aps/sOiXYIlhfX
Xc/rcLpxNU9/o6ytlzMkbohlxBfUOuMdXksrFvPAnftZzSY3T1BtvH2Fe634cgUH
cTaM+ZwOeCQq9BDTIv2Yqqgb3AxWVeerNvTOOfNiWA4EGJ1QafRUNdRrUwikgD9O
u80O73YnGWgy2bmL2x3dzUtoaP5+hQmjDst2KgvqahYnOCAtMkFSDK0ZtE2xtOt9
0r2NSQX0cdTlyhpsb28eQFvuztOI+4rSi/N7SM7Mi2zM6SkLrrzXn9J0Xugd3++J
cuKHg3yawubnQnhKXwEMtKd41a7j3ffnyvYfA6e0AEQJUqOoK15vgqsxFr54J0wh
cLz1c/E0eQzAZlPIBeB99/cqgpcyIIxR7+OYgYY0+U8tU6d++jSeusb9B+23e7I+
ecOKmXITNL865N2LOrqtxhdE/+VAe6CVXtXTg6AthDqb0M3xVoTMPO/edFaq0sNM
c+KO5gixsWUEwDDY1GWfuGOl73ehvlmwJrAvKQfnhROXdjqPh6ilOjwkn0LDcyO0
u62ogOLH6Za5EgPvFrQA2jeEFO6HjR44MVnQguNHlXuKZp2Cp58xj2zGWYbBfwFm
wZEaKyKOHyX81oA/f1u0faJn6QvQTk42U4tHD/w9AZftSYVyBvl1fpl/osMiuMU9
qy294qkEdhKaZC1tNJJdBpGi7vvhTxddvIkxx++PM5TpbwvQ7MlEfib9Tt0/zXix
+BOTLU5sWQ+P0AxLfbCyJN6q/VmhCLNn05WEai1EDSCgEda3RuBHNqfrunkqzyve
iSbsQvl5adYSYk6beNiVtRs8066JhSHGooLLx/qzdDaeabJInFjRHOpffeLkwkHe
yAK51PxlH0P4SZUTTUMKhlupZlFwfe009SDRK1KM1txmJexhHddyWMEQtwxThL9X
5GW8yvvk66ExvZa4I2gmcXPFRfum1BqcS+nR1+zGMk/25cmHndSHQXgzbTtsRdwj
1HB3E6BKMY7PdImHKM3+b8xh5tlHG56H5HWGebm3UpqhQFF0yIjXV2LNqqKhRm6U
aX2UxZ9kwOc78d0QaF/oRSAEVVvlqgTlKkROtbOUck5O5KUnUniZ4oZ2yFoFR+z8
6IsHWx6kIw3C17SKFa5ruIMf8LHGkCpNAkGsEtk/bYdsykSB7iS7JTg3NkiT2vNI
lAgK0fl/d+f4s+dikoOQCMK+kJJwxd0ghCPTp5QEnGbky7q+xi1k+znMFNMEsiGq
MoegJB/QqOCxJ+QfGhqBeBjUsrK+ZvLj0IUeVh/xha+adJoaDap5PCwoVK6wsp96
sMUgB4huxgMBZFAwfUXw5U1WyijJdi47WVn0EBTQrVJBWsXIOMfIRqK83PsFbA7q
YXY2YidrD49c3FvOnR3zXxqM09IlIrAtA73rFlqsWad614GMMu9XX8Yh/L0HGWvv
l8u/kQ4d797Xqm1IYG1nY5UHB3dX/dGJof+beTXfG2yulvZS3F/hhHYQ9yfQbB14
DTdAgBeCX3Fh09/WQZXHw+n8H6TdjBW4aljj+BRBzzQ3+Lajg35lyfyR0ylcRedx
R5p5v/Dvv9BfND16SEh+fX5C5XlD+zOfvI4QBE/PhhWCBKBMYEjTpoLWg5dRdDwc
kAgzDlYFwl/idJbCyqigjsvViT6pgzstUpNcHWXlvYzit4UE80pcYecSbAkGijs9
do6X571S3kUJcXD4P1QAXCTkVfoXVoZKgKkxoJI6Ceyos6tgfV4ovQ2e7WUNa21L
kU6a8LVQbJqeiUhFz7kcOdYo97ud+CkOlhvH6l2TBIUymF0kD2+RCR2Lhwd6pRs+
yguA+XPLQCmNyR3Pnco2EEFHlywzmC5LchXdjsNZFyPTQw0SaB/dto696yKQ5Bco
fewmsNh9oe+MDhodClB3r5xx2VlZSFwb2jF4TA2Q5d+4yUwpuHMbSJXcdqJC7p/3
9FfX8u0xM4/8aYUmnOo1ihDuiZCeDIl1DTAONDOdwdQDn3IZQOJUz4hhSUCzDiBn
IHIFscUkxYt+mr5z5SbVdLHfsF+eC5uegMsad3nXplsFgpSZTn9nNNo0aKRkJx4N
JlU/pFy5RfN8PeGThEFJzQNnxzKTaRCaqSUx82Nhj+2Afh7fwXVrDBZj5Zj2Ix3E
uHBsKJU/bpV1PPsQVWrBNNHHVCAX/yzdpx6z88rZ9H9fs/dfNCpVut5g4SD5uszZ
PQaXJ1JV3dRs0160g9CI29xlQSu32UobjU/oUjfIdCCw+Znsb8bmXhJH1p720MGe
lCA/pgySiDVBgII0MCJnesidfv20IZYoEid13g6QXl/6WBQctdudGZNqewtLmrFX
3niP6dPy0aPqeRSwLr+YPwY8bQ0uvILccuEHktJnbThU88Cdiuhh7BLxCuciFQNF
RDTrmTZnViBC2YfEDRM1mtSkxAgHyahKaXvxMBAz9XWdvQSZ2Fu2yPGjSgRBQLSn
CJP3FqigREHnIq3XlPVOjEUi4B9USCcD3lmL6FV2YYQw8asb2ghTRsCFqTxGSNNS
oVwzhyae8zkCaARVjLHwrgAFFbkWbZOU3LAKHypLFSE9BoSJ1OIVDJjnKvU34Ls0
QpkRA736ZpDDtHcZIctqfvIDTK2uYFEC0Fis8ejPqhGiCKwgPM/G5/p7ecO6xa3o
rQF8izmMkxUIWlqqoAHfO+axrvjG8sHB82d4SP3H/eGeHO4/ttgUjZ0aOhh68kpu
OrS9nWJ6XNLph8JR6ToHLGBX3/z34YXdhK5fdlFBrm28kA0ifjBFmWCNTsRtJ5Bw
pm/eJqsFIvmod1gVkEEZShBrPW51zNsbvaQWd8+pEkFFE759Nf/C07MzrM3u6DHF
hBbKX/L/bgDNVKFb/tAH7AZY35GeUotPli+AwDgYQqLaDOWVMKVpHof/NvkZs7l6
S67Y+ktIeSMUYiGSqKk6j+H/poiuxpCg0l8hpNYkLePNWf4YHFPeQEjzQ/4e5fLI
2ffajpR3IztKZGGe7akPJGBs1NIQ8viVsH3BNDklRk00ED+gtmic7SKJQs4Be8tV
3FpH/j/WUI5lzJcI9hkxuhM9Gw8wk0ST/VDLstTy8t2l+tqxvBpqNXesrFzpgo54
dJ3kqgNYagjLrkRqWDG3fAfApFCeOoYfV+IFlvT5eExQoOq1bsSbQc6ojQ5Mb1b2
DmrgFgjaaJZx3t91NFBXHKNIcdox6M+zeLJgNYzh1DK8LYSsi8mBEp/aIUuIF6/D
VHFbaeIgH62K7IVUYb8XNa9Te9CGIsQq5A5t/ykkqCttAckt1t2fl3O7zAJ35zJy
bdSI/qWlX3X1RQN6T+YUAUWIeKq1zyvHR8CngSGqhffZku4wDSOqQ2kXi9b5/XwZ
yzGFD6+vQUPhNGTmYTh7B6hVWpi6itasK6rNEI0CQ5NjYNCF+PQB7ks7yE8lPXhG
iQr4X/xNFV2r6pwYlR9zg3+niOWcfAXKGoCZ7ItPmq6fk8i/XFxX1XWHAlADJI2x
djZA/p1pXPWi07mS6lpt3sXXieTfObnYDi07DxG7Kc6CM4Ljm00nBIBZqL543nhq
/TAUzom+CBfa3yx/u1PUgsFFjWjXPGBRxfm3TrekqKoJR3tyWJUshSEdW4QengY7
H+d4vPTBaSmr6SHwmHqRyYyifkZyOOF9nvQfOgPYQALIDrrCTgogVld8TyqkzoFv
5TLqTWMN5kp8b6xG1epd1Zv4H5aWcEe4mRhAgxbDN3vGX2PYOw5uMQ3H62Em3X4b
cOyPJVbCBkENVzod4Grb9kRMEozsSafZMMeFx24hjTQed5/rmOmNVMhSJ5TM0t3R
7EPVpNrnT+auNNVgBpbxuDk4WdmCY0L56COGP9MSe6AlmHhN4lgDXHEOi0lSeMVE
kj4Hfkvoxp4gYkXwM939fLd4/L44V/3X5wQYPcH2HWY47UKfoRXbUHl24IC0Spsa
mEoLkmwztZtx5q6hBBLj/XyPFKbuT9Uzw1utllSNAy3LuLrcv1Wk/ejnCA7RkkmE
B4MPjv6Qjqtt+xB0XMYPe8v+pa+yAT1JiGMnM1HLwlVcC1H/3aqlHtz3N9Fxo+/v
bYFWVpyNAfb5aBoqMXdjUCiNKKdZVd3zk9MMRAr13NevgKgu99kqylnKbXk9UUr5
5FIhHBwZBqief0bPN7iZiIzHz64RJlA8FpPfugZYJILXWsjx8EKmz/SUpntovgDh
Jgrxyc11C/YnYclyVjVkJf9ClFKLDiq02PPDhulPWu9/v5ITYmL7X0yUYKYbu6VK
4CpdQUrecP7Bhp52FeHt9qQT8XIBl2QVvNfs2OJHbPYbJ5+Nll2U34Bu5JUIqYy2
BE+tKB1mJS3c6MiyphN3m+lAgb0O59/jz9isDvqR+JtRi6J7NQzrtWv4zgNL+x3P
di5PHa+Ib/TXXTqPtA2qrF093M0UVCt1IyjvJBS6ocqGVNbsyXhjjNi4nicnXU3H
ARiyNoysGzomUDzcXDJIvX21jJbevXyPVw9hbGjBrd7CZN7YVECFHLd6PNlRiKIs
OZyAdG0KFOARiGyDZiBTe3rRbobTCChpYRk5jq9+aLaZZu5gN+BYfN2mXOyNhIEQ
IKS7bObTmHahSKON36z6bg46weEz7dpAT8OcB29TaFpfvEea7ynFlX9mGCiYikob
EFefW/M1BbmGSkyvvBKr7Wj1CFsTuAf7UvGVdLwlmV2PlKHwDgFn3Q+VIzxHUjmw
XTHIPAf+jnK798+gSEwlsKAPueLhdf4SWMZjADwrWi+oDkRJIrIu1UyApzuy582J
I9BcZA/erxs+KuN+55wI0HCruoz8hW1wNpxSRdtavwEN/VjggmEhRdX9GF+K90zM
Nq8W8OftkWuwNLQq1wDOcBAfEScxFvTLbWB8OZguCW8ibWHXQo86I7oyrMo55kx1
G0cGq79Lw2xxfOntmVKcM1NcHL3fS48TQpFiwvWw0T1BoIloPfHZ4lD+E00PSbun
bJ9lhKJGKK6JEK+lAmvBNiIdw5mKhJ8hnjHObOieWe2J0tcWkZaO7ZQDbjb9jWRW
nki0hoKB1d5xwuUuES0jvPNMhONr82TTzb+6iP8gdmcf25NEssGBnDMp3v251/qy
47PGOakBsNfIdfJwr11F0u04pKAyB00SN1AQhFBxFTwje+5030Y6vREqwy0Vr27w
j1CKDlFFtUVbxtV17A+pnyDPNK4CmZKxytH+s80oYTpcJytiVEdN3qt+aulNhjrn
fY4RtRrwsK+bKRIRcIud2nQ/XfCYIWGf8uHcRjLpaXA0phLYHNXzaRsam/WrBB2z
zO9SAE6ZppRMqyAafW/Ermc1SZl16njcwyVPy/72xQNizUrBgj+zfO0gjX/X8+fm
OaghwMzDiQwo+oit1hu8sdlew/t0Sfswyzx7pcoriWcaEhBNm8abRJirm/lLkqiH
U1s7o1Esb29j0POh7gqG5dBeY8XtysyRfP5E7iNlXjv7RQSmUwfDeILfYgRn8GKx
f14hYqdcTo1+nsFXL8Ufs6fEnDzLR64Txnx32SehiUfquM7ojAplwnoIpZwTky57
EfNI+3eG2iJDyhdfXfmZYrDlP4tT4I+8KjoKZeh7Anl51BMHZc5IlEQVgaLAZl7r
g76dZxzINeOXyvfV3GjsuBv3qhrdh52R6+4upb4i0Yt+xBt1jSeHJ2WubD45mtTY
8rJBY/8cAezMIglhgJOllCp/V5Gdf3Wx3IWTyEoaoVXBs0KrfXTXnawG0p+76mjm
pFW+IkiTOzZ5BLkL7NEQt2l09w9D4wrGIl6GsflbidyQ+sBvLg9u+fzol3WmN6WA
Z+1BfoVpE+UqRCADh7f5lThJsRElZruYDfm7sM3epFUaDYCMBq/lOTIld00CX9jv
n5reNKvKNx2I0OlPN/GlUYsOdSdfHrZB8hFmVN5yHLrh3QmdQu/p81lXjbJPhzG8
ROeuU4fvfdceCWg0990FAmuOx80t9ywwzWJiCv5702lX5eQrJV0SaOsoyFgLwOgs
2XlQpPf2vvcKjPfO99zbUPaIC7ZiXshGa1+j4KF+Ec9P5MkYA20qC/nSbeJeoqaH
v0K20inzXCqDAJC/vdi+zUDPw6ZiC5YMb7/GBsQVsII4Oe5R2WQ/DFLd8ROaCt/d
JBzZFCzI/K2CdINArV7tfM5r1T64kd1fkk6Cup1Jxzqzh3DWdPSCrJCBTl0dEYqs
stRgzqbvb/7xsGRpiFo9Qtm72Acp3i0lP/z/b4sOva9P0riQ125+LLLmyynuNxrp
YP3lFj/Z2xcrKQubPKFv33XE9Pxqt3voIwiOi+N06nY8f5eCjO+ib1xzL7XpPkp0
TRveg0lpb9RjVAhLqIDf6WnV6EIdCf/1XMn70C1GTTITG5y+Od+Tqa2X+EFLLJXT
V2RbOU86IBMZtgPHByJbApMMwZVnNNzWZROfPgQ89id0wuTuVX0R71tacqTldKeR
H3+gxN5SRlNfRiKiVGx/h2gqThhDB0bvwW+lnPuxitorwcYy3A1Ahm4RcSv50IiA
ablqTlrARy0IXMxSqSrPBZiWAqVeQRL3pwJFYc/9ZMg3YtaSmgTnNEsef1LXO2YI
QkdYEOMnQGsVM9PEJhJrj2hNx8VSyIkIr1+2K5jOXjWOAEFysm/SHybe3Ro9V2M0
RLxwoNuAHLt8nsVD+KfNRxFLBxqkbG1ojSn4BA0bXysRhvt1m5kS6wCag9eCGFI6
kvW+5LCJHjNN0HOJf86qkg9wlQbV4WywKbz+ZJD+6LDeywN9Ugp6HXPafN8vy1kP
WLCEPqh7q4Sitgnb4Rs40RwRmLIcNQbB2lVTIG8/o2208hOEoLGcTHB5ymS6RxNI
+GadSGOpYfxlI4o/L+OV1GztW2Yfjx3AEcuUZP/J66okjiK4bpuEK33kzdh5tHyF
jYrsTPhuJWfKFRfgSvfhYVv77vvD6prmWe0JW3cfXdSccvanaU7JwTPpmt3BKjxr
61+yH8hhy5EzeM3cp27NfZHKIijp0w3PiYkrd/+znhpq0UwotArVGvxVqTjylgkN
MIY3vAcMSxczVVUm5cRWWgV3WSWIQxS5BNPIFahoLoSg2hGZ1Ij6P4j+H6hxMkbC
U0Jp3AlL+R/OiGGSdUAaxE6ryDv50pHs2SgqsBRxkqssMWWOeoqo5sL+QnFNlN7A
FIOmWCOvxOgWKacM1WjegOjtbrT/cghd2CmKJLSuPoN3TZm6Y1lAtAc8pC86ya8j
arCL2bu48XxQqXFyM2Qf6ow/dslHN12cvGsRStNZX9dLm+mKOwJm5DllgEwPRTPh
+ed81U2wP/qtlxRmVT/I+MkXverEgewoQY5Kkg6mwxkzV0rMMFsG+bhy8NDvkAtV
VX1Y2HK8dfnBcESkRoSt2QHpie0SpI/V+ZwVI2Sgwnt6Fqwao/ziDCBYXd/ybAE3
rMw02SXw59WjklWqDE4RDlEC5I4pxdMKtBUaz8I4ioL7Lm61A9Xs4PfrH6XIKDcM
Vi2eb0Qih5RQlL/L3lDp+zV8PYHrZX9ovAQbaRPmTGvxIh75lqIMfnGMRD/zBUjr
nBm4ejzVCU81zU+5x27OELjS6ry7jw4BCgZqkX6XGUedArwmJ0DBMIg+K118ngAz
o6hs8DNzQVPtN11nhnnxpSakV20qroPKSm1qDv5CRHD5HXiGdSU6euDSUrU2jpsi
QQi8qKrVZoci3+wxwx5dEDI8WFJbjSfARcnp+25edrg+LhV8skrdwCOuuIlptH5t
fGf4Cav1ccdCpFUNse5lIXVu0JG47G36t1Dnn1zZOf5L4atkzXvFKg/XWjVTFLWD
58SEwX0O9cqGKhBElTLHE5SxwWer12QEstlhEuqvBLrArlthL2U/vkmI2ujkFo36
84O+A0bXHMJo2nrVfd0vRu7K+02EFoxmMo/3ohjMV7ZBe8K6Kuc7NZJLo2b4afyU
TLmbzfdowzyMhhg/7b5KYYf+llel1redI6p+eUUezKymMBKsQYU5tW8DuzHJhGSd
9LBdvbG3ck+6fXnun3VpDsaCpUGpKQK0A5xaLQlgRDWrJgq6ds8/ifzb8QsjXNgp
lnSLOOdGMI14cOh/Weww/MFprznKQ3wrTDjOA3Ppcvk/mxJs1VNLd+lQZWHDi4NA
nBw/z1+FA/nHqucvTZLG29RohG3k34n9aoJnv0u5Jo6u9XbKAiqW2+rWt0h61MYC
veGHfbhCVkW6yo5M1pk+0FVfWr8Fsizd+zcSs1zq/wVHe0MLP+RX7zqn1MoTjwVf
KyOakTGfxmobEb82LfLDwGLfv0zs6EuZALkfpvemjjrDrIIWVynXACGRkGjnPnKc
ROGiAg2T+xgSmdk4Wii94w6pXnssoCcSWqalHJvmOdjU5xG7zyghDvlRi3bi2jqd
2rfAVeIh6PtNxOvtFwJSKqePh8CX4vJL45P1GJS24J8B1os5gKwrsVkDcfDO0NmN
XRUsUB5chsMw8wl3tPW0mgARKjoTs53U1fphoaE4LwAuhU9jxKIF7qM44rR5e/pR
fBD7mJCi0f0PjRyfl4KX9q8hEx3D0KdknurRK8QcAr2Fd6Klt/Z5x37EcmOjWiG1
FCITVjHY6UpN8ABqskMDOHxFaMzKFEWG6+PPxLNBHG8EFLuU7s2KbXW9FyqZAWdB
mcb/NuFYJuqAPbYfQj4rZb9QCzYxqYNZhW3uaIQS6ZGLPW+Cckh9NrjNdOSYyqpP
wGLtrWjyrHgoIYvm3nrI5+V8GaohvcZNCX5kSE8Ry2Z12vkgE3RHD2dMuHPwYdwR
3LmlZ81SviMs3C0dAwUA2vp/T9iomtEsp8p2C0xgsCsFMMRPxXHk6dPdDztChXIQ
AjwCZrmPNUeCBn4SVD9I4hip5SVghqBF2Y42ZQ34KpGDEwmKakLWzyS3AVFzbJXR
8Yrh3E3ZsN3VFfSuhkUKKasm4HRAJswq03f5lw01/KWLY+UYtwJ4NJTXARaOidzw
a3hO/Jhv2SfOcEhJPM6CSo32LBduKr6vtzQwbQgmEAtHpfVwtaUwWOB+0xorcAg/
Ok+YX7fvRKO3HVz+A+345xQr96QHeOi0XXQbdCORRNMEJJFawH2Q+9QLFt5oCdnq
Yq4zOammobcZYPgjnn4qqTS0GuMOwmgwwCQ6HrcsWSihp2G+KTYHe+/acKC6mGVo
7tenyIyxvlXTshfHKJvv9ZHeeyRzVlONWDTGGqNZiWAr6WEfqQvlrwxZ2oKfuS7C
jA3e6nzYiKb9serA2EC/WIdUqUoDPnhrtHj8JtDvQuw6hCDI26lBPAp+/kUfbxwW
Swh/SDZCanDdalQ5rq5tzHg9Tk1iiAl7p2ouL0AUylg2BUZ5i5bSMXxjPvKIMTwQ
oXf0fJqVe10/tp1DUaWJUx7awyC26odmajeDBZHlKbVGBKKh0klhqgQWEEBNUc8u
rkZqcImA+4x+8SpJSssf2fwtADwrYuPqhR7NW9MH686auXpWF6TAyFF9kSbGP0rb
gXsmjAOXM1KCSy+k8y5HKK0SRNu0BvGbzrMrWjPiQzUg0TD9/+WugGpnLV2j8OBk
SSu+tlp5aNXO/s01d+dOlJoqeNkxM479cSDHeOQIRlyjMaw2pj9j6T3aMrQcrvRh
MkQ6PAAPnASSyFVnnFY3FzIqMYVdOCq2P2cfU9IZnZhsvojBGrVL8iBKRgP2M6sf
2Uf6ujqg269LosOLkmtUBLF9dHd4suED5F1/722oIceS5A/ALQYB7uQB/vABokud
5ce4WLcue1CHQt3pPa+dFZ6Sbu4dZnGodHbWtYR/QPhfXlwPH0XhFK6t3fj/qUlr
o5ZAOycslIS3lwQ555ooiTf33aHYhsPnjjlf0s61mtNtt+uAoQS1ZKlB/SLkImr9
tYOL3nqwJ+YFiuOfP4uUc8F01yN1fjm4/LJZVbTLO2OIkuKt7rdsyNz6VxCgJm6O
qtwwPLmgzjPEXTd3NrKXVGNtQx/swGfR0dm3ginpX9gaOsJ7yYHJskcHfu8vlqce
/nDBkXPZavpm/PqYAbxETpSknidEqLboZCegm74ACpelGacewJxwK0l2xOEm5va0
z1YZL7bSGSo7WqM0QCHeTWNq12AyL2OozOBALjR6ZulS6JxAf3d2KKPh9vfTDapW
2OZJpOBrqoBBGWYjB40S0hNqSFpHboKkTMkLKUPK4hyZG/7IEVSjyabXqP4BX4bg
WhRM5ngPw63GDKs/dH/PvdDtAyryoyDZwX4V3CnOqlozbBR93eGRiJn+HTs8jTlF
eYo9WG6kdBjWH38+VXa3yTE37lDKtyv3hIuglfFHKFx4B13fPN/+QPMdBwPdef2/
opE4b3UVn7rEty5bUA69m8ynYwvl5UrNPhcjx1LgF9jORNBUE98B7Bd8YMbiHz6p
G91dWDeGknnaTtKXkhvZ5eJRizbCGuaNavCnAchMeKgGSb/XbP3bZBfyBu9540j1
k1NuhkqI2DPpyQ4DMhUg0ZUJNrxVru0zzmEONmOo3CXWhH+tYKa6iEU1NUXICpdz
4wanrQnhEc0iomOFR57VUClB0Lvek4L2kJQW8iQ6wQ2xLrjjuULu+NCwxE7I8e3K
Zha69wbdTnoP9yKQpFUrF7yOUQZt5fs6lQwdya2SFqhq4H76JSF1OSAthPDmN/BQ
hWlotq++j6af+dQehcm2nyjeOaZhQoVa2IabPFWo9Dbdmr919TSoQFXDDfUL+mHc
s4AO33R+dMEl48upfWtktTq8cn5daDtD1Ue9jkawLUJc9b3mWXTAer0WgiH6Mjm5
ZInp7O19oW5VoM1IqqgNeJfUv92YwkGCHkdBKGdWA658W+u9xPs2pOuKHaZGqxYd
mJ2KYoICSBo4DsJ1WzlhvYcF5154t2cXx3wtp2l8IS4W97wTxNsZ7TpUZp2lIyI5
DFYMJrgU7+YnquosYMUHyrBvPUp5MHpnrF1HPigu4DUlZrb6Gi99ZmUQA3FahS/x
UCidqi6FEq/AivRGz6cgWaRNME4giXz9yj47ti1wFMQy3WqK5L4jacPkR+qRRz4P
FJ6ytNZTdnRFc45Zg+LSwJ/hf/zelz2bvp9e2C2fpWY07psKu/2EaiyPXyARlBJB
3Dd++RRq3urBfArZ44lRw5lnwKRKbyLGcit8zxrazvWzIRsFjYtIs5IJSEoVA4KQ
ZzbJyAc76/+Js2H7tuAep4TV2N7vEWRnxgnnkO/OEuByh+yijYWHi1u9oMSofgzi
HVBcESgj7n9NG6YggllDDxwHZhmTuTYGG/KWN6OAync6FPBW7LIbgVg5r61OF+Vn
+UGZqQdoZ7O+qbY00VlfIg2H7huzl4aTiy+3VfrNubdxtM1zkBXV+Gr/sf2Gx5Fy
VdE7iESxPD2+u0m4Mhe2599FKGX6skPXH2uoZ4TtuQxKMwylqBuEYgZIrj79hfBq
B9pypT47LdzCIL7rbdfw3u+bYCm3f5c9LvUe03GLLzhyajNwFRnrISDC7kwJ5Q7L
Sw3o2kkR/n0Gy+RRMwv/tMW/JQw28N8mDvz99FjVbQgwpe2KWC6TaLiNu/NBJ0bo
Cc9ONpI7f3uCFwALW/i4RHcfWf5XUfHctB/5/Fq1WGxZ4NZW60+A+JcjXZ5YhO3i
gxBPzAbV4SXSXrATjLnZDyErmT51oskz5dn2KMhGgERiXOkIJqbGWMuuUOc0Cdqd
qf/gqemXa6mEc8mVPNQo4V1qynB5XQ2gD2u4RD7SRuVUtAHwH4BjVRanZbxkJLEq
PjAcmVz2BSYHyRFRwKEFcSNaxLhbfc3dAE9o1kEa+bkwo4FsQlIO+ShwtaXQQuNg
xgu7B9/VH6vXWGm0WGP8BWgOCktKdtfUE5+j0FhChIseqK7k0t3xTFnN24pHDWBt
ajYoWINRJNUPqBRyuWwp1nBXNa/V6wMzZfcxCYUgw9KcbTRLAB1t2sofYDb+MD7Y
jmcZa+loWwhPPXTj1n+y8UJsae79MJZBSsPKTFGsj9h4lz/sdQgnVg/z5krTbgl5
jMVsHwV8LsOXpkxzgRwpax4YlQiI7WaC3Hb8ce3kSR9LYAmY/BpTWa1Md+a562Al
ZdAn+xiaih48IM5Ueg1qAnDFaMdKI8+XU2LGT3e9wd23vjLy9SrKSyI2F9a3bVow
POkQm8D0gwl2QYbfr8jIn+/9deLgCfObTv/Po5F/aaj6uqAVBpmDIDCLysvrQxAs
5BSXBvwOQosMHDlcTMRN975qO6wblp08TLLAlTs/MBCEg9uFFNJkS26RfK7l/Vo6
U12c/W6YLvio+gophxNyFUKKI97MoS5eEUBHID1LaMKGox+XiBdM84iuCpMIf1nX
qjTkSFmAwrgP5gDYexgR1/MMYMnU6K2u5DqMFo8bxDUaBN2lqpaWcYaY8tkicETi
rsXKNSu83RIWiozEDFVARPhuOXZpWxQtZAOhRfpjrbbyQ8rfct5jixbIzLt+aH/h
L89H7mYcvjv3ZZDHMUWdZ+CHlHrRYcj0OKFz9OWY/j60Fl3ZzIpDxvA0nhvUUzOQ
aqgNkWcezu87uVNhF+aA2LPY7fGEDPCyZkQfiO1AeJZjmihoBm6PQc3IFIn8SoCU
aGCISI/HNLzEPlo6dovnVChahW5mfX+J/g4TvIu/KqcpG77GgTamjLEXE9MS/8po
foTzQqn8OloL2J/rclm/ykZzc5kfFaUM1gxsLv7GC5cTnvBPJg+dp7AYChu70b53
kMWjWs+LbWaaDsmdXUzOIHC04p8NVPaRI2JRwUoL24lTb5n9vna4E3wR1HYPUrfl
ygPDXrWNEERqCKO61WYOhT5RYykF4UyK4k1MI8+BovF3hFzp9CBgMWUm9DTab2sp
VV/d397u/RwexQxr5aK+dzAUeRpeS0GbSGZpS+9DIzXe7zQ7aAyqIbtD03V8hWs5
6qWrl1UrLXtLiO7Hvyqhgwwpr5xClwRgJZNGvSvnZp6kEDg7KJCoivSfvCwqdVJn
VV4FTFlgVjfpQYz5cqZb5oPbxNqCGKvCEJD1o2U5uM/mk1s3XSnrEEaljd87oN43
cAB/H6AZw9l40mPvHJfnl9HCgRuJ9X1Hu16rNYc850tbpr/jNKpOT9FzKGYeDeWJ
n1EeFq3AJpEkU/WlLSpfvk1TNdRw/XpBN+6FO3rNrj4cX7Uccpw07GZrzA0msoLJ
cNm1FEUo/+AzhLdKarUAzi0TxjG/O5GzkwR8HA3XRpovcmyiNpfuUDxaD3vOCBfr
URZ8H7S7ZlCAGYnuK0nkuE1/w8sboRau2ykxHqpM7luFMR0R6b15zwjNSAKxrQOd
oaH0aQaWQFLKGQ9ZxetMTDX1IRNHfMaoHqlFS/SDEkwy9qGHTfSWFR1hLDbmYgC5
vd6hm0h/KhJ0vHKlH2pXwlNUbs4MQ/XAPe1mwsbTgoAiSVlyA7PJ8ktFHXPio6IJ
UYlQAxv+pmY6lKbW+NX/d5d5BkXo+ZvVhBL7QfWdQoJYbdRCmVkc6OYepkBEbMhn
iIy19g0MGB4mUc9wxxqIpBIEcN4BDhUGrEE2jVXKxryXKEb5QZpCK3WrdoA1xjg7
kI7WdRSQajug6JV1oHsyrVlkDFYRsMF9Y/teCMYPnXo2uNttuDFzyNuIbvtOjvPz
rVCQJtJFHnwNAPGqz4K8WCgqRDO6S5fB0ebaur7hoD4EgxurlFao4jzAJOahUSNU
CtMPr0ODGhpEUxQ+QsHFA0Fnv7bwDqHj6hHRpIzurpBgRFEPE/zi4zQKty+7h5n3
PhSe+aQhLTzqJ8QLreP+/LwaEYPprTyGHQYF74xUdh9syjlCxfgfDK+itX7gXSfB
b0fHX25meE4yECyR2LZeKTzExHQ/8a6wqjWxlTiv338FJYt0//ZEpJEcvlAdC2EF
LIO3rOJmDFQN3EKWd+KNsAnyQW7P+M3g00dZ1gqshA+296JMJ65MyCWfXMTGunnX
xi+ATGkaO0OFhrRlr0pPIVdDGOUXwlNiQTG+qn2JVYeyuikEDGS56atAJGaB1sTI
YVX+mN7Yvry5o4pcLYTTQJMPMuiJ2xSaikzGW7TaW9yqXd9NSM7JSCTdFwRTSIFu
u0Denapwz9Xe17ueoFWz0aj9owva7iRqrDBWMhbwhGHC5mURuojjhKPGJNIDP3Sq
6y/boEIMgnDR9pw+ri/OaOjhvxKGs3v4pFz48vUvq6dFsmHnEuoPwHza9qOECHys
KKisTYZkliF/mpPyBwGweoahN6efCClspXfvkITK1mUxYTm5UIZ8AY/VMnQVEvtZ
5O27kNW9sPMs8rE0vtkU7jIPfVbHkoFfQ/OD9rm0ZJaSfIFKZxIXuqPSfoME/ZSc
WK5RN5QVz0YAChrOjl2aQb0SS0kvXZeAkgBkUYxwLPxerg/94xp0PezZY+2l3wze
kUapfyCQCbsVmo6mUqcPqLdSMVkGI7KZqmwtMnAMhBe6CD+W1GnKDc9gRqIzupj4
zqFUidRBzYf+ZvPrboM9r7IduBDUZbpwfUNdWUKIJr2KHWPkmy9xEQ5GNxoOdT4x
2YIkMCWcVG7bxlF0rOG4eXjYeFgNA8y3A4vTRuTxhVn011eck4lQqAlrgjxiT1cl
9F2+4Yq6soXDmNJQwBGJ+QPVOJPJfJjJgGG2oZL3UwqKQ3uuWbrNXI+Zh76cB9gm
Ef4857d34LmBO4/N3i9ESlYJWMvC90XunFx/Ddnj+gjTi3wh2gyFp92uJca8T1pK
wUvr/KKiL+olmXojDEaB93UwJJnf3dm5WMjSSdRbqP5rBW7sDShf2Pmqgp3ETJZq
tZvHVNKZY6pLZ7RhOruyqA61cuPJkmxlAEwcEugat4nIN8FOlMWei0DGAI4qU5ga
zAmys0Ha0ritgFqFeKXTQS4gHh5AUVO0bhDWCritsGravBMAUN3YgWeXSkh3oxAp
WYiFhQld8/y+bxdx4bl9EHABgxA9/Lnr7ECENCcbQfR59Yv93cPsNqpv12PSWf5I
mJXlBGDazQc86zaenhnuswfAwArAgPKbVtwenyU6+ZzLAdkCjRZWjuyqt2SeIYwp
WxOS69y7MHaS13OnSxrb/H9GBnDHZXlgT+wDvUyzdjucAL0tBuREf+R6QRSizoZM
pMEiGJqkQWW1j1U0xZUcX3uzoQYXbhMlQKWdFMnZ6Lh8FpX7qC2nv/8jZo211Gc8
8SJcLcuAZT/n508lqErabH2wqPRzvDBPny7xaQr/x5P4QnimcwuXmAYhZfwPtc+0
7NSt2ywSzzgHx93LpN9b8DhqWmDJS1CWjlNIdrjTHe806+ylsNm/x8fvsoyPyLsH
8MdmF4u9Tw8cCAJIG1aKXQpEGfAreN0BTrjdi8lIcbEFUCzpdONF/j/OG2baTezk
sfh1gdsLnzPyfuRsB9W7+GA3qWN1l/kO/YXkAJsHgo/u+daKt2H+b4pcEMM4oRcV
weOqa0vzaB7GdEx1gkgQCb9/ktKWbLR3P/M8+OIkFcKO43oQSefHcyuA98nNEBDK
zePG4ALSl4MglNVQGGT3E6/shhAJl2TFD5rGdNMGFPMLoyEy4kPONYabWiKLpA84
oXKaH6PlwUFdxLmLWNjvS2pBZNahG/NrtQ6v6H8yNAZ4Ip/z+pfdxSTRJqAbpEMa
8A11z1VVyiGxq+RkAdCdrLno+eiuA6WrcaapmI9pr1R8YF804dMImvl5iR+5hofQ
IapQ3d8v6tKVObM90cn6H+AwcHyFZNu3QgKd8dBWVMXWt/kv35tnXW6T3lhIOuZO
N/6wCfzxvCbSH7u2AmyVC8Ap9OxRzAVRNfuonCiIHz6KOelUdgQbdsE9AisaRYNI
448jASBqRyQkQPf4pK476B7oGGzhJxd0uQMTnYeGudotiMdhJ50RXCghIkXnQhiX
42w5ot1Q6wcV7y9VUgW2WaQoE5pOjqtMdJGaNsmJiuGsajtpKYF8KklXBYWVXyRF
9F82naTSYWY3kGyiOA0EcHscX1n80TDXFcJqSDCrVmcpk97y8Fir12i2zGKGGr8/
DZKbudsG7V/TH8Db31Hycz6/NWbuPDgZ0p5T/aZOMMw9dEKH04gXxW79dVbrUOjP
KefA3AA+X3/8OLvLpmp/0J4qlHi5kiAKpr9116J5SPZPvhKZ/fDPxbr38PLRHFmr
bpwGMCaw+W57IupoMX+1W+pBYmmTPr44Zze8xT5TPgAqQ3pE5/uWMUnwl7Zm13dr
LcU/w2xziWvbrIQdRFSbE7oPC/EZ4NKpuPTgVXKM23fw5+QLaMNEkzEaA0Hw29Fo
dXjaSb2hoVoRJrgu5OB82DbG/MBvORSn4+aodgPuISTSFsDW/iJgf0HqTjM8bgpQ
/+LCqaAWDTSnUKONPbIIREl6kLgYZ/kCx3jJ8EUmRZYKkj/9Nvst4wQ0gr/578hQ
INsTbJ5zfLmwLp9XPdATpDIaDxbOsM5/qgZEacCj6XAMtO4IoAsJC4NMXPJYjZ8p
Dv0uKHd/QbGZCTvms5SPYowwBFg6aoZKkPmDHbdpUUIGRVIkb5Z/FEZWvbn/KvRG
+n/kbmD1MH2zIYi5Mjvc7yqJ9pau8P2X99xZPBU7iWkv8czDsEvONhWW9dTK1+hk
W+oDxy39wVk7te70+L6yxfhSTJL2KD0g3Kyh0YkRg+GtS1kA+BJWgj/pOiGxGL9w
PEOl0yll3DLi8zUEDFPi9iBRkJGwVMg+LrxMEOso6oDVKhY9N9EnHrMzz3EUd122
n2P9+vOYGrONvlsWAlV/90Up4VX5Et3xsAnEMgxsTYc0gMQJoS2Ii+F/OxTHfbCF
u3+QVKO4o5Y3/ZpxlYQW8qpSYqpW+XeQZhLbOjcpYWIHQjE3+rfnyhPKkv1LyoLO
PEIos5OdmaKokY5XbKs7owq8ii4xiC6fSyzzLYz7jcgCg7V/wMj5Kxn71CUGmZXz
sz3Fov1OnhgqAvuMXDUgxl/kvY6LH7A2tFxf949ToqbkD8m6aCgerlunxZ8U46Yh
4FyTaEbAva2XqWK2XllRl6tPZ37ALqTMQDQQuLebOb+PefUn0lLkxYS/MSAj1ZPz
oQeAX0uEoKlB8zUb1u/pHnXm2eOs/0cw4ivG7JTTr7hhrm4mkQHulvga8iLAgBnM
uZPsDRtI2h5W0UsPrDE1X8kmlomd3uIEPGWWfTZhsvSK7nAx8aupcvqi9nhgK1+r
A2Gm4LkXJDK1iIgc6dcD6cpJ1L20UfAh1heBVskjggtMtmfWrW5Lc10WC9iPhPIC
+W+iqx2xCcrJDk9c2V/QIo++4mbCkPUsK9IqZBR6ePSCtRQJKA0vzeTV6q+cZQQ7
upEfRGzBSVokqj0zdEH2BYHYfQ0Vk2EVfag2DR2CyAmWg795afCxKv3nX4dfQLaH
5C4rcceXoTLj18+P0niESc62sDYu3lk8wmiMlUh3/LYc3h6UgWzjMy6cCFq3yclb
x8nv6lqckLmMKOT3LNyLkwsf+4gS5vDnUlfNeQWg25RZTMKRCJgNlDbgUydOC1Sw
mMZE+9R8mnShs2lPK0Dm7HQEAZP5hfKiRCz+MIZhsP13PqHxBufF4kMmW2W4P320
YnI0zwJMd05R4xRztRxYvMwaXoAkTuYPkFNbxDje7w9lVdUp3oDLr6MQjwe+FKdd
AUL3LUjGmkjelh/YDun0oVHawU8Kebnxd9+lR9Cz423/PNU4SSYnvg7RLh02VL30
W9BCr5poNBOoBRUoGnBmMIIxaX3lrd9wdUzNUpLCIXkTttoH+ur1Q3q0SmlXyIrd
HPwBmpTjpJacCvZksciOcm98vSI7ZEaagd4uzaEGm/WyCiM2unJVtkwST49z3Jq8
lNUPlm8T7usfIzizb+diFzHwPCtZXVoQQsHNKpSvIVJeo8WE91sYZLEyP0fMmnm6
EarUjHqVWiUsRfePILc1hVwiGuzIRWWC/R32176yzbWF+5N13NnvEjugVrvZzv5L
tfsKa8EubWbMbnthdYuaisdgQGImCJME8w1Av/uCiFKKzBQ50yLTLAOK0NuJC5M5
3h7kmVpfKX8o3A33x4xqu2jvn+S5jVfY4fuCNm2GHJJwZGZydHuvWulOFuJt8lNo
sevvvbcla9J1Y0vvUjoQ7BgEh4V8LyPJNiFMBLkYmQf0Y4x3h9RmEMGEG8y4vC1M
3IWhXKwgUraO3X0yaOEIddQ+glppbZiuBzd2p1d2R0jKPZd9vPfnONKgZ/v/O9te
kDdaVJUJUlmbRHChSY4VnV8Zta6529nzwQl14AYQ8urJN1lE0EdW087zrhSMnDJp
b/deKw/peK3d7ozQHw0zlmcPXPxeNL/eUub9wYbwj/x9yaAxGssSdeaEM0uzKl7Q
x7J+D7G1f+s4FbBQyi45YUVQZ7puztK+TiJYHFGtCsx24CO/762Gn3Vs4Yja/3Wr
0fVhtVf6GWm7ridzGDmKU0kPz9PBcG59TBhTcC/iQH+B07tC7udSaCLL/iIDfEkH
VMpofC+svFIDIvoF8ncs1hVF4jwbEsv4hxKFNtEpn9MqG5SlAfE9i00xqwEEMtXG
KjL/wgB6MQ5+utGpoh6YGTKUopz8wJAZEy9caIhKcOcZI5Kvy4p26zAzgNbor6eR
TSu223TM3e5obPWXP31kwk/Ah9mpSAiMT+1O03tp2+WQLj7k3yyIkA+fGw28qxjv
v26sQMILKqYpM/ecz567RrDZTd6MdkTNoAe6T9z2iJMPd0UreTMyRvWQqLeW2fCd
3m9fGuOwQce5ZP2z70i2vj1amhGE1BzULKmv5sdNhmqbrxhitWkyd1aWP4v05n73
bK8kjTq8LcOqe329VCU+M73K19/u5A0vssF1WqaBt2PO4gyJOMYt1BgdLvswX03y
sG2xpaVyvKmB3JbG4bUe6XXu+uctMZ2Yz1zm4+s8uYg6GdkUAZb3P95xgsvffmvF
nIa5W+P9AyS+TttASpmsShDM7UxEOI0SFyT0bWRdHJNEij+XSwAWUiM/ABemybhb
Myt8QUtScHpSGB/rFLUyocCcgMsxQ0sEjTYY8spELXfQjIbXNbFWbJ3njpFBtInm
Tc2gKP3L3bXzrw90eXMplhM1phLdSi4pJDNCRp8NtFYubTH64ioUWBJutJKWHQHb
4zP4m2tcOalWJMmsocIQh8KAyXDO7Zo7X9yhRLJLxei/MNaikMhVWbmiTjWWPmRn
23b2+ygnvCKvECLPB1/SyuKyM/NmQVZj4ZzBn5M0mn1jURprXLkPcAWaZL2ger6O
o/86/g3f7PFr71dcgEaM7rXG97+PjFt0TghAIx9BqKJttC92C1FxU73SPJt6gY9h
xg6WtXZgL8fs4pfnnl0bD0D6ykPcGZMtMUn25v2UBArq76FLkyGHdQdt3xOzY5IA
suBUAb5kcUyZctIM76szBTgAZaIfDVh8rcU4Q04HeeW+O+SFLhBWPnZml/CA0SOr
f+9Pyz6mbU1r3/YoQmTZCIbPRoP+R8dv+LuItmMf9ZDMq0uoe++nexVIggs82DTQ
H2aeSOo942a9t36TdY5BYGqbFzmKp6Ndr4aUJmoZKnqJUHuRzeA0cIRiW3LkO9i7
EtysAGG1sBmnW0GyGxPrXuBNgnSkP1g0kpMI2bQU3Jnb8pN32BYQXcNBiB2ti5m+
vjC1mblg1+O8r5oIIfCo+cS2Jd2KLQND6sbRuEbGvjzPRumcQd1yHmZ9urNC2VPS
lQGXh2pH+UvE/2TE+nQ3GjOV4vQy+E1A7I/O51aQT1vW6SG3ntX+y3yunuVpwSzu
VtfVixeYe1XL86qmHO6csq5hKWlucsJ55Q4ULEynjCuOq4b5Af5NIbmVQ5ekXPAS
IUGEIPKPChsT9qWhJ8X4GL3eRo2CIMx/rHXJoHta5NgjBM5+N7vOzG5s3tl3IpOm
R7BbXJs3gsU/XKfpEBXAQzMfMuLKOOQI7dCe5yCWfZAW4oJf+H6/nAMak7trgmaK
gY+1pqTZvPEU2s6VgNeh8H4Y+8fubENNrlPJT3GK+TO9WtROzfG2PsyuSkAWkBtH
ohnhUTJwoHdoxPVZf6erWjqV9NhhBrFuwv92UNOLiCEkD9e8MJ4IZBEYaRUxfBdp
1yvxYufdYiEeGoQH4ic1F03V0c0u2/vXG9kOz6WF9BnzhI8CmEzwobFsNOMIIw0A
MnAHTEKJwC8zmzYpHhVgtcOXJQkg5G+d8wRsUzs/qnreCmYDfXJoLAIsAtU76GMm
ePZ2r+9dftwxc6kt5gQElDUc6ZJgjWTBp2M0x9kV1nJ0lPoFTXrFRr0nk/HtM8/A
2Z5PEzeOtcicfBK3r+NmTma2b9xccjsKdNZEpVGulCm+T+H1kPYunvQ57gNxahfA
6wqXZiugTMnGiK1byXowrxDDNdXEF2ccVVYWIGNf2dr+riJAv8yMRtvkyrmZ3Z61
vjhv8se7slOz2MJ9DEL8HxFJciq/YK6lMnx7w5yf++W3Lkm+5ZSQNu49ERdGukim
dtZIiSV+cMJN0uzelKZDr1oH/iTJjp7+GRbra8VaXkaghKvsX2ViMI07e2C3a5rt
U9A1nKPm4AzI3p4IIzZa78XFxtFy03PFojZk5rk+CepCtCUVq6PpHnP0wRZbVVcl
u/fMZZVPyKoHL8RdwYgvdw/NQUyPjD+3JNQ8bYs8/wXYee9kk0fOHQ63xhLVnL5w
p8KuzhZp8Q6hOw29jm42HnFE85z99QauAqHiBmhFFUH6XEXpSQB/hjW1zKIm0cNl
xRajZQHDhu3M0VUjPFBvl13QtkWNvsWzFGBH1jAGGuxZeHQ72vmDieAXlpXVKKLM
W4US7buRFf2z8pQUArxQ03MgADtQ7Ivt6EZIK1MK+ir1b0XOIG9s4Eip4dH+wsYT
qBun5yYW85npwiKt3WqnSy5dcl6361wNHdTUtBcuwzfSCE+dwhjr9uvgKi2BAttg
A3fX4FMzOiNq3h4JDJJ6XluTMLJNjLVu9x/R3dE1JRs4dRzugU/YNMDaI7jbKYgt
ZyOvc5Pq5QOr35ImwD5/F6eT3C6VkzfbOHKmpzclnKYwK2hftBTm4U5VWA9NaLK0
JE17YpFj505JUC8Up5Q6nwOInX80IGr9vMhV9M+F6m92t9Yg2Yb2TtiiVLdCVjGk
5wcZsBpgl5UwBleIDQ5QSmjurRyNQLqXxo9G4+AGCtwXTSVVg4PHD+wVSuyYkhMB
hgCfQVTvnAcYVrxdYUVsZFYrfar7d89DGuQnPXZgaktTddARyQIXhlYwM8AgwcTb
qKofoyDuAK4QPWfjAaLl6dTvr0udumDOl8J8iEym5LF4wAR+LeipZzD1C0MTbGbq
tJ0CueEVM3jxzEvaCsWo7dymvj3U2V4BW14Beg5cINhJu+D217bhmEtd5QvMmJKn
6oQ8nvxDIcUPVmrGPD+lauCVEpxd85P14cpTOH0LdVN8C1XkJz1dO1TqUoDkmM66
uOFnqU1Rpa5Jf0MLuia0OHLZwHJIYqKhS6G70VlcAYHeyiekQTvDnjiaw2wbSOQ5
hDCCI4kCCaqDexy2nfnpmMzQeGDXVRu59jnyTUzBoZ82K9ixSp1B7S28hBjZ4eP6
msCZuYEZAZM/XeYKsZ9cjh2gOpAN37DYnRUP39+qIKJDqexzwRLQ0ym4L9+qTH5V
123+4MCqFKkEtM5ON5blKwxySW1b2U5RafPURQzhs1N/0NoWInkeLPKG2Mr9Kqvp
pDlFJmtIbt1ibfdfRoZGAzTMsWqQw0MDSD5q+Yg1+52nKFDO6zVLXomEGDUqlGQa
NyP30jh2CCCaRPsw0DD4BVx0OF/YFaUDm/OGtWXBJFPj4aPd0M/AYSifU+ctZSUZ
GuDhl9qLK0EWw5/qASZWSMncWAdbrm8D51Rv8rjSqtvNVAP0fpOlXPFEbMnYC3L+
D9ZVcRS1PFt48O6oPVknhJuqxDRLoGhjR6xmnztWZgwv3Cl4VvxdcMUHTBspHEQ4
ldU1WnSZgsNr6fU3ggplQf3oBbeNJBzbiHwNFW/JFti5F+fTIaEtx5G93o3DXFzj
/7R8LUcGImJra+fKXgVyaATQEr7utU6NOggSbgn7RRNbA/oDU0M+400U1Xd5MYfo
LiDXRSPtuaLwbnEFGoAd0bEUF9gRzHtGBmSrfq65wuB7dbwwNgXyvdOhR4BPoq7T
I1ig5MJ4mRXF+f+1GaS/4F3eC3tiY33vs/2V/eA5c0qYn6F6HLTAgNTlULfeuPlG
NlTieW8ezcf+xwZDTrx3QDFI0PnvRt3jC3fL+wNz/pp1UxwIa1vLgGrLkUlJpfxZ
VHhDirj2/xoOkY6B428GWwDKQC1hQMq6Zla8NdwF94xPcVFn8GH+u9gkK1nRhFze
4+q/wiUOyKK6EHDZXp4QsauhS14Nja9etcPq3JeTxNQggM/6uSn5NZdR5mEqO3h4
Y+NcwPAedv8QqNnV25ETn81pkb+qdUDW5we0izUx7nRY/XJIXrfDxpxRUfS4Lj9p
SKmQzctazNt6lKhH2snFqqOcW61vktA7I4s/j5I3MDj3s559uDw0o0MFEcGfShmu
H81qVqU7O33uTR5LII8bP7S6SYEMVjJD6NX2AuxIH3gdb3t/jq0NcAKQ0SWOLnfM
0UwvAWmm8a1rFTcpfyWDo9ydcxaEHLNmWu6obXj5gHKTLvYEvNNnzZk9+ycJL1De
74UUuFz9ZtE7aN34CkaDJYTd5kD2FBvatN34NJXVjbdUjiHP110G7HmBDVstfh0v
m9XI7kQrCD/i0yNDFwAHbehr9JG7pcU60sUC2NThLDs5AltXQRFYNrMlUfYNrx8A
OFfkZ0JXxFiI4HH9MGSUbTId0STiloiYv8eF8vfvMDcmOP3C183DCjmS4kSkC5gz
fGe3SM12xaOYyVBX/4yVSVejWm7eovFHQmTxql3UbpvsKYG4+OysMWJxbQneTIkM
JV1mh5svZqKqnnZzGLFLRUpb2Ktm/HmUnGOarWkdMkPV+4htjaVIOcoLJ8sDiTuR
jGExyKT8DzaM/Spy64luQj2/6dvYHrtlSUKKIyK41ffzOmHle+T6cG0vM5/NTM6+
ZVJx3Jy3aLwA9Vha/R/a5CuN2M66D9h4Rg5jSu7+Td0AjkLYjtYyVsG4jSYQLYaW
N5nnTlzjKIFTx/85J9zyN3ZsYat7e8fu3MZfHPaRoL7dyorHw9b4PJ0Zi63Fzaag
Qh4PCKk4V4cDd5lC5MTBRk+BbH1p0X/t0rFSfzX8PD/QKu+XgNTRVBNO10VRLNq4
LlaLpa6PkObK/gfu8BOrdiP/Veba74+5n5mNBnYk0E4PG8yL3XdV3MBH62/tZKqh
zIRdmPVGx1QJbG29zstQSRh1P/Ck+Y2BRTehM5tZMAafauShz11Qd0sZ9eV8V84Z
1PiPJ9c1rsG5qsLEWxqQFcgx2JnbCTgSm4iyNQw1GKNZjIO0kNSbUK1/lMVI72B+
FyxsrHTDRt+W+qorjFF0IuPGIVr1Oyu3Gn3pFHB/DlgPNigj0rfkNy7oCX9IEzAi
DjfFLiyzmGVpwF5gZfuEXJ2I/6HYimXRegrEqYuz7u9Vrgp8N6j9PPBq700Q4j4q
YRGsM4NLUqm/wkAOAtZqelJB8ltwQmGMfBfvb6asesdHciZGA4k5yhi2gVw+UiSj
2h2AiUoH4mNqSBUwqbxzlkcz5JtkQ+7ULiY2zmf9INziTTL1LZ9bjA61GZK/KNlZ
bFyzv/CwriirRqhQAilz3KQiwTqP7dYh0gQ55mjaj7u0bwvUsEOrN+h7rszOxDZE
ee7FfjQnCuLEwZSjEXc8JlXk1QwfkzzN2yG9LrdBjZLNePPYBiWxE1Ejj5Z0hArl
ksaLB3oIltpgmcIFtslm4YI/tIdSyODpSZ7kes6frXKLFuEfMYF+0mDXE+Iqh46d
o/PxQQzo3SwJv/4ry+qRcuLPzNUYHQby2tScYxtiu0qwEmnPCzhFvGf4Gp33Lb10
l4GaNSEVN/F6mKYxAwQBoXRVi9IZrebWfk6Dk6oiJaUzw027uzidxGoX2asjcsAx
HeMxMnV+noeff4JZ58la96ebzF0czHqtYXtqgGJQh9tnyHqjXyeBiupiur+oh3Yb
OPcVWAir3YFGYhQIhM559EwgqgEmGJMe8EpLzoGVId6fTyiKKUt8AIg37AdiZEqA
9K2tJ5XCavKC+QqAcPImaaLwdiVPubfmqgETuiE3IzyLbuF4+wAEq7YKL6K+g1by
NVnm1bFDXfZ1yNzgTd7ad6ieINnk3wb0lQlm3/RES11Lguxs/kwfgQ7ll/NnDEfU
HVVvayeZzEY/n7pkAWJVbfQ/8vfsTfdo1n6qgaQ5LxkuQBuXSB6osa0WcaQTfJK7
B8/p/l1c4Lq+/HVBfiXl1QCskz8dRj9pn3RTxoAIMvDPbhWiW75yjIPVbirX+bVa
JT7H2lOMrFgOSBh8ZxiVxzuDlQ//vyLaG31zrYtQVyE8I2juVARnarWo++MCHBRI
D5FTp3H9Ecx4ft9T1WBzs6OVm4utTKcpbew2J5BKSiMRTyD8lF9idBCLGxD/tLbr
3swJtuEJglWxe8OaIHmGyCl6hA1ixCHAEUvUMg4ZNTlYYhVpR/RBbEhHy3bkyLGU
Y6uxV28ORN5e4f1rVpNH3CaVT80ehSeCeMf0F1hA8D7ybf2ESWjHQn27f6qjHJIl
b5+P8G0Ye0z9xG8f8ReQU2qzUA8VZop8r6Hlcg8FnzhNJI3FPdzitdawQEbSDe9u
K4oiKCYOHvAKkuak9pU8/vz42WT5yYRKZHkGUATOtQQpEOkWVrLUmqLXxPBbYq00
KXaX7yy0HFNvaKAW/nbAgrVFTgzWUtHKQKRObV/qoTntxkmrpECLv/vH9DbqQMIZ
EJy8yerf2BwXTmsXI/OX1MO/WMH1AXXM9kHS6REjAis9p+UASRBScQTu1Hvdkuv9
0jBlsb/ph6KkMnGvPEKbDu8oslXmbgijApV/CL1kMqgNLkw/+2KESvyM9uk9RPM0
5IFfDsBGUaJavd2d50IGJFjxYChdB8LU1Idv3jM7wWGXCSz6x8/Bt/rZ4Vj4HB/L
ncSyE75iy7O0FMBjYu3duohJj+EI9+E+NSdpSGPw7zMdxxeQ01mAO+kxoexHWFQO
f4LrsTEPhJafOahIAVxHcdfd7WolnaZ32dLvgjCU/wkQFyhKW0ujdwFcOMK3GPko
Fgu1I0IRGWGgTm7A9WGin4yqMJeIGLNN3TAoY9eQzm4tzhDQCtpeRaQD9Y2JOLVO
ITpITyOGxmyDInttx4JE8LZqAXvvAEo0I7HmnkgZ7qeSfKnpzzrU8n07oCjDo9zy
D1kfnGjvxklOoaAwiyGnnXGvNhp3PRoS+HbYtn6dPsEn2R9QtiaRI69DBtkicUKv
//9/4N7RC8IwAAkKGjuE8K0g+bClwxVbHodZfvZRJ4PhKj/yVhnmogcddgUOjcXM
wAC1t5PS+s9UAcXdWvMByehH1jEMSjfrqdAb8eLq6HMBwjDsnUy62nDtFqJASkzU
++5U4zOAgvTFpazD8oa7WLH8xO9Op4xHGAL2unzVSUb0dKYW2m1NJo7PBFJeRFe/
mq7Nyk/9nzwez9+IIRiQXocHt54nStc9Rsl5cw5eWGb/3PRmoJ3r57cD/Rvd7Xsp
rgkwVTwhEdOPPKY8BmFeEKYLuHMMY3hjjC/YwlGJbmQrOMNJW8c0+26N70X8ziI/
SQPLH3Uz7HWUjz9id2COl4Fa/181epZ9gTKtcOrV8zpB/L24QypEC21SzL4v6/xG
SopQNPUAdz55xpj7aqfuU3WWBSMS80dMfb5gZYnmE4y4xUC6yCXFDhZKqh803/Da
/NczOWR6erIg3jmIgk5le1NDRLvwa5pjPkzesUDoAIscGHGtDfEwrtLC119P6TZJ
p5Lvm8FhlQUQDj7kwyuVtS++m8DCEzzCnkP4Hge69ujqW7+zQcPI8gp4r7ETTP/d
O8jDgcSOTyd6tNSfm4JO2yUuvfZL+RIkQMgxgzWpPVrePgocQF+DBJss7FG0nPZN
xlYxs6ivxJ8WFZcZGf+yuSWiGb+T0aYzYu8uIlhMyKDFMCStuL/e+lvy4e+gS01f
ojdm/yUAtGHQGovLc34R33TxshIex3AZ4mhTgWLqMmIg3Lnuf4b/txnJQ3kOAjtU
46gyVLygpvvAK6Zox1keA7Gq2IJZslAUMgPDTfjw/7T7Ve8Fs3EGAa/B9RuvEMIR
8Tjoq91wa+agxOFLVeIq6++30yh0vERu5JlJ5JL40ZnKRLRwg4ORuv28cR3xmXk8
8eIOw+MRKxkGX0yVIH3y3+oUyZO/Me8FLNUkxs+VMpv7tKBeQEZTH+Ym1Xp7+uFC
qXvL43xsxS/4nBNx58h5xsoMWsI2fBk9xlm6fj2rkJBbgfzR37VdulKCYt/wSX9R
IncFPRbbsWyljVZeYaMyHGAWdcMcKVfzQkm+rxRaKzVzIVaCwmAUI6fIdji6todV
ZDW0jm0I1gqlKlkMzPMQZQBZA20WpewiiMGmB5MAB0Uvd5lOsnSCtA+G+m01z6WD
K5JkYsUy73nDgSKEd7cPezgzfKu3Sr44zEVEHqA7OHibuxBHUO5cizp6bf3vKlrk
eYxZjtfhxRtkoIFOFbZlOeUnvr0cx3LGUJ6chpGh/1hGGuo63mW49x4XsvhES/fA
ZmL4DKNciNtDv6LkSxjhI0CCjgQdFrDIY78cJokBnMJE67+0Qr9C2iUX+sJQbsx3
TDeYcAzezavKsfdxkzq26onUhH85RamxSBrktD/gkzFnypogNMLyldCB3yRcXdb2
H6G56PCLE9/RvaISUKi2zPTjcPRucaixd8tebOI01XRh+XPQE1AeaCStJzfjuzP2
2Hbkvmzzr/GPXzAHOJjJ3niQuKO8Yvp05CNXHtiXPOB1lu7RiT81ggFQxIQENgag
nzvo4wUhEAc+mNP/ugBuUIx+aF96y/R7b8f+zVrekazpe2WBRgblcKniEfVMJKWu
CFTPo+pzbFqOFgrQxZe8/ifN8nNuIziqCyWl7sXRapr9kGO6ytYXQLC+ACqw3lP9
UtT+8pG/UUb+TUWWgUXzop0mWU2NTGKRSNfRMd09ZYGWZGmhbmjc/c9BZh3iebdY
rGxdfb/6YZiqRUTqIRn0F/NBB1qRw3D/LJJZNPdEYdc5+P9QxX8OliEw+ayRlpJP
Z1fFtlCjdyChd5tZq2Y0gOW4+KQxwl3JOQ9o9FUKYw3s/6mj7qZnnMiqdUcq6IrG
YkLsBMltf67vhNsiZvTUFWTupNpxTqAKIPRvqhBtjT+HFZYUqACI9cK0vC65PqLG
N23qkSG/cqSf8f5rFxAmggfsv70TgkWhLBSYCdY3wfpFD9gI4FdIjXoC0hpNqftM
podY/nLfcBA7XkcLEaWE2WkrizvyBxrNDjZ0M0TxMLkjPdE0LjK0UjKneAkqoaub
nJxvQyzzgcDic2TZ4ad+7LLRZ3EpFHkboYQxuox8IIIIZwFYmtt+/sj5FXc+Orym
XpOG2hwIsqkVKoVG1f3sIXlcl+f+iS3QeUyzRlO1zKAP3wmeMFOKhMpAwyMwNrvt
8W7aP/yBhk7jd+Qx8YtBbDZdBWCxgYKD4wdRT2BjgXXo5KDoXeOs9/+r2CZcE2ny
1l2Z+PKmN+49TqEWxgvfPWP2+Z1fWOBi+X0NeCda9pYj3MTjCJyPi6uhPBN3cRRk
5FCJ0XlCgXeR3GwzlYWIQ5hBbu47k9FqOjnRuULmjm8QcR++/HyridhRI1Hanxcj
DH4rUsMMNnZm4Cp9dt3iCkasNxyMEPRsp2IGKqiTRKbD1sZC3Z/Yc1OLHXkjHnn4
bUegFUEBzp/E659CazcwuILfEgFRm/nvE5+XUoXDaYxU1/jeRcB3uCELSbFzF7Zs
hJAKz5H93zyww9+Bg68587OLCGX+NZ0fpTj9bwHTyfj7aOfrbIHLX1UbIltgIQHW
n77CeIl4AEiVo2d5T9kXcz2X+QeMmYGi387kYRnWAPGJGQet0u3uFcVrkLAfhil8
yjNCoEM9a9Iwt5/8zBPnEuoBnvK41s7OAhoSp8yEwnZ2KW7O6stQhLzVZ7HWDfJ2
qZf7tQN3UAGIwUArRbdd2X4c0j2tCCKTGuDZ4a4dRywQB2PS5yV2mxpR7XyOvcEh
ZgGCdwiqeAdl3plgxc/3Z8kuWUQqigt3zgv131Hc9fYPc+9QFI1XKcZZS7oU9i/L
7nj545Zgw9j2SP0xl0xr+S9UZfvaSMJ6VbWO2DhOYi50VL+a6KUIAW0nPFh7Wm9c
rW3Aohq/K31ccZV3UK3Gwr9N4e10+HXjljoGMLVV4IAOq07XaxllE82/cLtmQsp1
JyAIt8FKbhSHwB6nwgkGAPhoQkzJcVh7/RPliL3sKIDrbwaEUwqbdkncAGWBPi0C
9P50a2MsGINAGnJkWhlXnwR5oGr9HVXcrvSLaerMBcp46++Bx2hP/vcCnSeFqccS
PLRxwOT7PZbq4bD4yun/XJ2VdaOG2D1dQMV6hUwJZp+4YPzs0saz0mRHNUVHlie1
K/GlnaVGWIPKa2TbSrg0+4bNpkEWCX6tXzDpptQHOnCyPvo5x6l65fkDqpFJyykw
GdX4Em88MrAEnAFQJ3Vziu8Ucikwp847GH1ZAIi4kUqPXz8oZYOhE1aoOcCXFXjw
65C+9Uy/WN1rqNcrFcmqtJTnkgjPEhY3PqBzA/JjL7P8dpjOJX5wZD0a3IKRyMLT
TQblWYqNCXE8AtuMTTi+7mpf5g4TCuHWog9hTmGwqLTZjvAHbiJfpPPlDCqoO7r/
hBps6j65FAW5y+WKqInS3LCLA+vz9LF94SHA0pjVZl2T2TM3uXfAER3qdaE/0nZA
t0KJugXTmYTEifkw4m4rzAMGfLOAQTpWdr5aJlPIggSKC9dMqOOnlMiS7kxXH18M
N2Xr2wUg0f/+kGppIabye3qpo8XuCk4XbYRZby5IbvB1OJjfs+D1mnl86ymGAF+K
ocBRYbmIz5CZ1X6DmYKy3/c6kpaRL7STJ4PyMtkmWtq9/16nh0ewlp3sjiPaLadV
v9B+sUADX1sRgBZb3Ih17/fkpj7mHJGodQp4MoG9ycj4OkZ/JjJeaOVJDv3S97NA
s/3SsWMbV9vOeclDIzZ8tLln4k2cggNj7Pn2G/m9ddRIfUsGiB/soPm0/APpXiXL
MVn0PoEKCxuauhnGq8RbGm2U7Oe8FldjfH+JMrjVnssuJYYkzCe/nWS+Z0AtIqvF
r+uhdyGznZB6mlCb8HvxuQwhiPzY/BXTYYd3hw076yrnID7YjsE+TcnsEXfcxIjF
dDDDrfFGeRxKu7ZgCxPTz5lUkCpC9lQr8cdCh4Nk3I1UL9Gz7Alj0v+mTXLdVYFv
nIYVi52V3k+n/dV68g9mmb6z+lJjdasjyZNsmFfa7xBGTD0mnGPaTqtx4HvibJYi
3bHaFCx1VV68Z2fTOkfzzh1TKgYxzYaHrf03msHF4I1EuSa3rYAKBkwejBJopdD+
OpOcmKe+dSTFip5KYFTEay6ZTRiepOhGLec1rVkqBelVFzrgcdfJP+kL4LePTx1V
WdQ53vtz6cz10wyYOKCJ6SyWS6r+iDmb1F6BzBQ1j36WD3G6dUbKKzAu3Ri51k8J
3+kdI18XJOPAneesqNw3woQ+MrwiUQuDolJKq97euWct2F0cIpIONMqz8uGWvXx8
lihEEx8iqimUgicrmrQ83xXPgwTqO6kyoHfMdCNBM93NqNqSmmlnO3r+3QnIKrVa
X2j8xunbps7ZnzcNprKWlOC1CrKSEWPgOeWhxHUU39MdVOidhEgyf/RYpwT6I5lo
B57ECEcGIGKhNZK0nK/0UnSX7/CWUEobOQtEUVqjZVvmxefizX43ILD/BAMd1EYE
IDJhI6vJaWBzmb5DXvMDbGdsYJe7deGcG0KIjLSTTCevmge0TlBeIaRo+6YVn8s0
oRO11XwC4PVBAQ6k9YCKJdQRdbQoQQZGOuSomgqCFf4XG/TRYgrZgl86P4Xv33PO
03qyqkMEbQPPo6QUyTcXJj2gg0xII8AnEmZh6PEt5tb/uXrW0AgOpu6Ya44ZBfRo
EQIBya2pJLDIGEuMfTjhLzFKdY/dtfupVOx39Cnsh3yZtPdv3JW/79naa3s3iTJw
AKh4RYsii/9hMcc0zEirMYsmdbmb+6qVTXSU4dxdkZ302lwii0YIUpykmFdvEQeA
Te3sWJu5Q4GfMjrwwWUEAU8GrSwDOhxWjxtXMen5FWU8cXjnSnh+J/oXQiWcPZ4e
zTcKuRbDhfR0MeriT5+QkvV/dl5LXVGp19EWGMkv+BBcME+RWmky6Ee9Q3C1GHW4
WrC8feZZ+0uo3RkUThMNLoIysMp+fC08nIn74+gqyeYRMGll2CPw4yt+a6KuHybG
KQ0DIa+NBmyP/caVsPHDommoUObhSaB/wzBsOGBzSxUz1976EBdhGVVN9R/+1WAi
NbWB/bWN2Ae7m6Y5uM3Ude8fPnnC9Xvzn+oKzin0k5xJgSZshHaW4rbELWADPqdW
GltFfZqZsv4Z1gkP6LzAOWHkjkd1xGUbctmjeVrCFF+wKG1AnIuo2kqa/ERgFOgL
VA22g1q9UKIprU/kTrtaLgTY3hMW3mVXfIvHYtpaX7hUmrFVNJ5S8aG3Fv1MPkM0
rry+rwR+SbaR7tWHff6XKZ6uw4Kc54Qcj2FjYVaFZQIHlYqfQfrdVUoXOCkFT0Jj
rdnRoi1gH7fARE8yb8NMit116EZBq6PpJjpfebgWwsM1z5Y+QVg7XdAJvNq9Q+zB
VBlYqXxB40EzIR1dJOR6pjd9Khem3Rv9uT61FUWpo0C7qD4fHk+mn0+R/SjtMrMw
AAa5eZxobE+ADNEY1tD9Rn/XnQ4KRVaf6bCAyz6j59yEnXZ322fddUegJMUafRTL
s02VcKPwmSczGWjIGSD9pN/7xhKjgvMDSaYf9VKw11GmPiz1Ic0Wxzfada0Ayu3u
2mVad9la+mPPIBIev/sIA1How/7cmjZjcVtuK3KQCto0lcrbJfYKk2GQkXjvoKwX
dSTTA0Sy4Lm0zB+Mik4C/k7AucZLnIkx6NW4OOBDdfhzTe5NVcUfyn8x4V8CcCxB
Xyqa6gWIy2mw2YGZUOLSqVn0j09t0BIkUdTsX48xCLKakOnHSPhKMZZnGBDEBdZq
iB2g3IHrxfEoSc+PoFWIbX+j6EHGwnwxXZ3ve2uxlcZ87YlY6oaofQEJDJF8O5yS
xTUySV1cjtpJkjaFHV/JbDaLVMPbrOcI769Q6Q4IpUucAAFaEflEFXztQK06keNE
ZymlEhd96lolZ8S6bTFH2BO5z0hTBSXqh1seKObWN4JqNP7xDy3qpNM3EZ8rZ74s
Bn2MGwqZn/0trCr+m6416E3X3oWJ82W7shRpTOuS48lydRDjWwH9KYaPbPlm0EHg
zqrXj6HzVkNavygVoJg8pgSP4lVs/dTq9UxGCPrhTVd18gOcH2xw/Vrf3z5v9aeb
WvZl8wNboJ9Lh0Kz27aJ3KiOtXySNt0Dg76qpF1E29Wck+WCtANCgEOOVT+21GBU
SQfADwONAiErHm5AmbcQPySE4TrPYNjRQzK4/pL5MLilPBYJpcGRGBz6j6ESC+WP
II35KiABrKvEdy8QjEH211N3NaMRm8hT9p0cdHmfbVDwar/YwzyXc0TnYZ98LPe4
ZVZG0Jf1nSkknIdGCbOMfDHDdzzLdsDshpixCdshInFi5POzOe10BhdmzMn/7aWv
/N0W2gvPaU2JiAAmaXIaMNtTq1HLTR+Y9Ae5BKIb3q6ENfpcR2J+abnyZlqnNIRE
7aQFz0y+yYYneyNYXqArHBiBrmNeS/0luM3UZqalaYoxul2L7+JTbjp3BepZb+87
2P2Ku9uJnmZZEgw+ZRUpy5j+5tWsGMpKrD2H1i/grmVg31bBUu1l7/qAmelrGCfg
rzkFYLZ8U2+S6NaCe8+CNGmWWrtH1YNyr+l/2E0P6yk3DuyrtjNCPaunwhYMepxg
SEeyFvgMtw3wQXJ3u+6vH1BMMB1PXFadu5fw2TSALHWJ3ib7ULpLU9wTj2sAnf5l
UCFjR6P1shP06ZZWKeQE2ww9O+qF+GPUtuqVzkVK8Zo0B6aoAzYfUNENHLNVhD61
CpAXcT42J8OsYP2Eoj6kyBuce5sSDf4HV8uDOkuUhkb/gC74zvkNNVQ+aT1Lre7/
N4jLVrh3X4Egh0UWHy5036zUA4V+oKfuzvtolAkIXyQB0Mlf21Y4frZ5aCY+XVwF
+Q/0wwGBxoaALQarrz9nU5Apho6pIf9e7NoB9b/nIUDoigzQ35mMz+hXVFyEjtSD
xzWyPmSCelAVzzjfR4KxKiGBefXehyYecXAOJfcaw+uCXkM37oBd+DJ51Dcjn8Eq
5g8WORi2h9J6HVrOE9a8/RDC2GneuPRdlz98bQNp2rhqcG1oIVEWYDwQhwWk3iPa
7/ROtFPUu1IqVPztdhNzpOYKW9B0lbJLvZVScSFoYa+q9MtUL3wD2iTShC74l+dO
c1E+DwmfyxNnU0XUdpC02ZN2UcGPIIY0adojJnefCuKYzYUyL+0iSQgD0Vjmy66h
fiSMHQanTmgqftRpVpKsGcTRrIWzzCRkgI8XEH9uxY0auWWVrkP96neAqeZVEd8G
DR3QXNagl7zfF2Zf8j0Mm5sZnxQI6Cx66d3mdTK0ilkwW9D/oqcucu0qCgKg1BvV
5lKiCdQYb0ji5ALoTTw/9QV6ahBj/lg3659h5DP0sIMXXWl3jCOkpvkkwFqEtIFr
v/4PDxuaEVKLxfFVy9uta74BQscb++uLJ1xfpUIMEZJeiXTUPJj7lXL5VDifVc+r
4glfQ3HXtrf2I6o/A8NBGiaCaopEHEupsmcO7K+qEOGXSWpu5xx03k9SibbmX8Fs
bkR7BmGg6U5cvJnfyD/Fed5knGJmQ+C8KcoVh9mDhzRGetCoAgowz00i92XVZXCE
t9Aihbsu+EbZvH4csfKKJfusiVWVLO8MaAXzcEPzgQvTApAECzgSHhr+rJXrJUb8
5YfQU7NF76o6gY+I5K0BCBe4/b6y5euYj9O/Wc4A/uqgrHCCc7O/Rb44SsjHLgqI
MTShpqRKkPlODZYeuYsETRU0DqIDPiKXVek3cY5rdB3aczdwibzIkyRZTSjh7ay8
KjIlH9rE6SNNlFkeTeoyVjjqyU11v9RJizEEXw97TrNLiON/MuPHb+JWfRCli5Mq
Yvlplu0DCgIVnLcaIeS5JzHSshcwRzaeFywI041tkrOAQ0nt9pLqLOUIltEMOTPR
/9l5qQOJY+h8s9oa2lRvkZOUopIPN2mmfOC2r3rik49XjOJGystEhwafBw1CYAYk
H6MO1/8kmINlarkd7T0WY6UysKCbEh1dxOa6A8+iVgmO9xI5Qg5Wh+S8hqT8jb/d
8YvvKILpEEfB08Mb3AiZknxXLfdiJldhru9/EirUoqMBkKqyyrf+9Flukv5C1Ob9
5SkARDNwgmzNdCEXPyPiEpIvZCVorR/C693O3uar+23RTitoPZHzE1bAbN2C2/Mq
nR2IO0PotMw16jGuTNmvcp7vs+EBXfG3SKzg1Ypo+AU7WL8JCTHHsMpWt/RIgn26
iYQIXOKNvCV6rSrdbae1cPBdkbg/VPnls2+vCmmq8bbAccXyLVH6FLbrkwVQIS08
yr4vy0CDyqnU3ZSj014ZZD4JtHHrUgB+bJzp8h1sRCVGwQoYY8OXq8Fp+n0msSNo
3JO2DZOOTEvNQQxCU7XGPHOHruuW3WdPLMFjhoRuxQGE/xSRoFtT4F1Q1kN0Ech0
+9lL0lUZ2IYXJdgMJWR07yqm1hRJt5qKwlF33UTWHI74w0GVRMh/48Bg1/m7FEwl
WdcKnH9OTPixsVzi//1i3VyyOuH9N5S5EJd4v57Ls030sgWuJ458sPiF6irdTC9v
RPFQPX044f6gSeJegCiUZ8hFEOFo4APdpSSupUVfcnkPZheiSdiEvE3hi6c7bWy9
XJwVzhfqhSkVh6RNqVC7acbUBj7/u3RTSfViAc8p3wNd7vlhbKVwpA3vmPxHMR99
7MG2CBKR/5A08Z4xJNlbe+Vjlj1HPJAh6KGecRBXA9HG08E+SFQHc6I3gZFd0cdy
S+FF0qlXRfEddb/8LIezv2bf9ryNnt7RmvJJvEkWbW96XYlIPx6GgJlKCxu9qy/K
JWE8hWVVzAPyA/GylhZUsnu8D4KPbNzFnMsV8GFfbv/4Gza5QuVLL/WrUdpNQdpF
4Ui3WhJeHvqs8zvdrQx/+P37uuold6tBlBv8HmIEXIU4dFn55W7OAcUhrxgurXI7
Rs408bLNI1DqMJXmQKRDF5UVpN0JnESynHrftpdVc58sdf8xhS49MSJ/Gyt/sWPs
0mCCnZNJFTPB/Fmtj8aNS97Q4q/sXDUT7LSdIW5lDA33gly1/FLEE4p/oT1hTnmU
4FX+8GGA+GCLZxsh/JGP850RfA/zF4rKJoZ2y+lTVwidewCCnz+yzqWnZfhSiKrv
DcsmN1iYotx0TIx7IbaKzwcqMVKj6hcWTZmjAYF81Lacgyw+KBZxj1zEtJem/+pv
adw7YI2xjbfZiBdaN9xK39+zjsDnTquzC2vzphqnzJ8QkJzexd8wGiwvfOXnyTs0
Uq9gc7mxXF23SiOIdxYqoz2VbVnzxXjOgWkBvokwOKaPXiGfWAj02IUN65dQ6aud
ud1IIfivXsvnt+uOK9iqPhS3sWMLSrN39cZ4VTRlzjTh4gJbHbbcwy++ms58BcdE
6U1AAlNlqMb1N7Qm7B4tGQZ/TtYk1DVZwhIqew2avwtJfzCPZkrCTkhVsDRdrSO1
kHfkDS6jCtWoy/cBpC7WBSusLAo+UxqXAKk0xnDYwmv3TZrORiNtRTUdmlOwNlHR
vbL6zgWxnCvbDXE/BvtB6plJph/sPT4h8bCv9Wbn3CTlXbcB7PvAc8Dt6dKJY4XS
4pec5Hby7ALBo/dMV+4K6J0Z4wTJI5lyHga/SOyX7witGqR8sPz6psNj0PmjGOqb
fq6O+zyJ8Cs5ex1goSqHsWwEOy/C4p4f9EBVVSkFSfgO5hw1PUhl8LZVxu/Yl9Z5
2J8AN1DwuZqw7BSdxLJoW8WD0lduhEWwsF3NGJNGM9TX4wt07f6vRYLxbEJeqJU0
822NjSlnmIRHdxl0LI9H0ryroZhfcIoGWuPfzI/EUd9B3uzdqPqUoFVuBDbHqiTx
/yYiaAC77KjbBTVeoZTc231dn8a+h2w+p9rsXatJe5t6RJMd3EDoyuuw19AY2JRz
yy0dXHMELb4sifgvKOk8Wndd4SfnnbOqThBw9wwalCaE2BUHfVefAewP3LfyCnBp
cSxNt7t0abzVVEvSwYohKusaCe9G8kdkIvJ+9WHJxZFUKatnnK1RImbY0jVySteL
bnmedecXkOhDCN1ip6EHod3w2+PnZnzVdIdxsPN2E/KY71Tp1uL5yX0qPwiRkLTJ
JdhaDEPMC5TBnoqMgEhaLYb0tijmWWFFeTh4Ph64vM8BelSELnTcxHIPnHEOWiQt
cbO8HqbdbjkzOkgztseC04TVnR8u3Vx0sizQds/cdq+W+NLHEkFREIlurS6zorus
LMGw7c+hMsDCgL675ZQ0gUEMHm6ETsbmcmyx3i3KmBTcvz62+96GSoANyU5Qq+vm
HlrBiqQrqZINBgOIeXyCMZ+4eqNTnOD5uTwOgQscUON2dcoEHPu0h9HiYVJz5WQm
Jc9b/ZPaFHtYji8OL5WejFWt35bRG/qL+jiQ17wbFqRuMQ/VkKEAxhCDw2XO8yGz
zuK9Kam8NWifPuM+6n9k6yPW+S6Ylfi+SuT4Z0EGUiV82gJ2IHFf3BU+rwPxCFBX
Lo/VTVcMsu6bRk/eGo6b4XEwzmJh+iBI7mWM7Q1wYbIScFGr4uZwAJ8DdiNyG8Wj
5q0N+zQ+v29OGyPuQ/SBpdZ/t8F2jPhMLxv6BnV7O/9k2C315oJ/US2tXrI0QSDN
f8cl6NwHFFj+Ldh7glRAdUv81Od3OicG37zUn/1V4W9rexds54FUZ01aa/Dnq/1J
T+pdXylo+tQSjIb6h32dJJ6se2QKI9Vsru+awQU/pmsMa/f07RQN5mL/B6ryZB0z
HSM1oQoKaCQclt9u6TsYTbRXnWsxQVxdpmAu5RliOMu4dvqoFUPT4JgDLGpzDvdO
DUO5PLeX4barIRZIROMv8CPFpsmD95jIpipsfgu1gSTfAfzBIESD2jqseeK/fITH
zKpYwONf9Ve7MFuo0eBeLWJixSmJE/LN9cdSOaGyTNfyUwFG3AjwauAubbv5e8zD
eSdg28LzChZ0x4Vql0HixhgN4ydmyZkLU+JC0QWdPc3JNTK+IxF/52dLyAzNLLCA
/9hc+q5yGwgYdTIYzZKD+8HILEHZuMT2kOkA1YAF3tGrwGWa9p9BaUDOm5yqul4R
J4vTqsauGAhZnL4msmgvQYPtmHvYjvc1LlfvBe9NkM4QUyvz59JhjuB2mdB9/oc3
dsyWajxYPGJdydOSJibJ0dvAStaPUyP8Z3jjvMGnAZ84JxyYM2ZgDnEQt3bbAVwi
4guz19iwln5tL83VIoDbgtRfKebc5i0WLKzCjOD6q2i4uQGq/dyDo+y4nInPt2E1
E5LpKXI170C1E9Ov2rlq8JiaKamkJa9yBhHMeVPdQzR2Juqaoi0XwdkQdcUBne8Z
R7Mk6zooMPWZe/wMQJT+pdYPcW4HoNydGhFT7Qx4jjJfjz5iRAemKYoynU4cFSmQ
4ZpW9PQeMyJKbXf/Faf6G0omwd7pKsuvX+AM/g6zSFJrZ7RmAbQ4rEZJuq6M8oCT
ZpDHyfAdZchykJ850QDmk9ItYDvduN7alDNTkFlBUNsb8ER6jOqLNFBNQYjQFEYv
zamT3OMpII37OGCyfUkB7rEqM8pBf2lTj+Jla9HMRTdQXJc5rQT23sbVGqN3EfYc
Fi44dAKVYumyM789yBQvN5qDrrbwOyk3Z1ify5sa+HQVShX1jspKtkg5zNpM8PmV
KoCg7uYqPR7dNsw3lsnVQTWOhobeGL4ZqxVMmYI1gZSYxFgLW3dl+Aou/E9FDNsw
gcIVXPQd+UWXWfl5POucpJF6RjsckFBTjGiU/Bn+QWq385RCyOZgBXajX+914UOb
b6eOcaZBCUyZm0iFMeu2Fa8A8GhQlCWxIEjKelx9SAH3TFKuThAOV8tbb+n1gM88
+KARQHyaVYrZ3KPvANxGOyWjT4UXwpLCMmK9zPo6CH5Jk3Xc6+EI3pif/ZwfDe+N
lQo9vVLya4xA8yVaCW2jm5krxH9dFJOdVcCMOKYDlrhKucvdnKW6mc6j7bzm4PcO
fNV/z2HcBbnlxfcea+MXVxHqBU+t+2BL+dlhlkUcMwlJ9o2NG+XmXmDYZbi9COik
A1ZlLv1Eudu23n5Wz6NB5q06TkjxKMI2ETkXvvrr1do6AfiIksU4iCavLRAqfLA5
1nFTY6+4v0IuuWGfXYA7Wh/QxKW7nBeq+K/HnwKYEZ6KXYza30KUJyMIYh9L5dVx
g2AhD8uxRGeACXSXkH3mI4iFJR8dk1CQxzwkWT3gXGtUCfXaGLKvlxZNEt+uxpry
NUNbwjDonhMBC74ZOSCC7YZSmkFFAhXkB8us8UVJfsV1sXE42cKlVkjk6jyrHNe+
LgwOuMsageOYM7yd9RZEkbGR2qCetAC95/n/yA0TwW4reLcaM7KNXntekCADu4CH
YBDcFrKZ8zVJsQ2jJzSYYXZHhiqYrpP6yhDfN7NXJc+AdpnHiYwPgpzrmnMyqWaP
Nc7En/DAYE2kKSYMxvCuRpPWzjYndEcWPLF9TOQ92WGVtpYQiNLIc8HewtAK6dS0
AuIha2fXrH3e4irvRiWOLfIARSZA/wVcSuOxrvZMcXzb5+N4a3cd2ODe3TyJBdY/
28LqT29F/t6ru+XJJFIWz4NnXNMLcCULBmwrsBOpikPEOJELJHVX4JxqOk1zpgGr
nwEb0iViFvxRUkC87Uzxv6FlAGYK9PG5e9BgONDn4372Q1XXhYh44F98YOZwNJ8K
fQfw2VYGTwwNhdRz+n9t+GDROIlnYp3uku0/lemrc6/CNGIq0qm9qi4ikrF/oBrw
oTqUo8MMI929aH35g3VKiyNENuWqh3L776G+Sn9ph2JrjZmlYpU3lpfTMjw/elZk
5q+xvH00uGDXiLTTW6FTkl3KxZ5U4LfJpXBOpOPN63H4QZsJJIRYp6lyPEgulEuz
AtLsayft5Op7VZVKcin/s+ObzxdrZrtFgSJqvvKdMxPUhpt9Xwoi3eupsjhwtqQ6
hEj9WdEcZ/CuxIncQ6KYzktVyV++6kLrWs8Pr5aEbV7QRFshRdCvX9x6BlYeCYAX
ZrLVBu26mLQ2ha9Kti21KHTu7sFbBMs1c33yuIxCrTu1OTz694l6lFljgi9XflmB
7UUYRt7GP4wH11+v9BJDv2jvaMnpsU6gF7JgMkKx6HCOSh8qeMvGvoLLSyouTPY2
C7lcAQ/vQpHSsXINJ/t3qzel3mbs9b2kNkz0cyHKfJEK1aER2J8CaOeE7YAz9RTW
RRZwXUA326JeG9iCm1fLIhWguKZFl0KUmftC0WptErEQSN3c4cb7mdciJpIUUqY6
BJgiYcsd2WFSWGiSVx18bEZf2WXIAj0KX4T2S2DZSFsl1ADgwrhAWRTS9MvSgeW6
YoLVBxLPnyawfOMvb0YGFWWZ2luIibaQQmq5N3uDR0Vbu+bxLP6uxXpr8x64fq46
kL4O/c8zb3nrX5ZLkRv/SbxigJNt+QWBD+2lD47sjQaMZQjNRoFaPlLAcIhoigIN
rOTCK+J9Bovx8A8VW9R7V8FaSkKmC4QcAhUm/ygrbYuFCAG4tpN7WcyJunDc4bGK
B/AWLHFM/mTsNGWDS6dAdI+wPnKoHYEyYLEx1bQT4eVC9msQ83Prn0iCxSFQ0Ceq
EnFNFmb7isk8F3CPMnRaY3ZLwJFcEmwAcwlmxMmka/jn3Q7tInwy4xRhaDzCVlt9
3xaczlth7PFG5HpU7Ni8026gqvgCN5QKd9bMdlK+TSJPNUDsvGEWXUZrYMvNmYZ2
QYv4tb7y0nMEqaKJlblW99IOpq8bDG8cx9VGYGULdWKOwDWlPz2R2C4SCYLXed8C
P4YieK9bzTFAdZxn81IjTuDtiKnG9kL1UsgXDVZ1ZR+yKZKcz/2biHYp5m9J4wIh
8WS8h0bhLrUTsYHZSU3uKQ5xH+IM3oF97lE/iA4nfdDpQpSSK1BsehBH2Rwu9tv/
6itQYDBJ9G0IVRmv3V5yuL7aPuWw961JF8STVxX7fF5Eocrafb/zsPawzGRytFJn
MdSVT4lmCLHmR5al8kPd3P5CPd/24YzaEOouo3AVB5c+RjuJIyqRFUwB+HnHBzlF
+NgqcsjvM7eg3n9SuDZK3ICXLNR1kX2p918cDsNpyPLom6YA4ruk7u6vQb5HIzbp
q9lGAIjGptXVUwQS6mUT38jT81K4nfC+2rPPptAwDgBG6nruJC28poX2Wws3/8mv
g1Xnrd0krb8uzbe5KGrfbKeHIzAdtVr9AlurqjGjren5O3/Fx8bOooeCxjgGcxVS
2d7pANGcNFFElHXNmE7+Qu4m9uIRCvKXt/kuCyLoaYUvj4443I9Q91yQWz5E7JwC
DT7dmeWxU8Z67HUZJ3y5QJ4ozuhr6VmkOSzWOSRdUNzogz1vwDt4tzZys4G+ZtRp
f8EcK3UwPoV95pL8UVmO3u2Tg72G1kUyn9P2xKPXNQobL9C+m4xxraKX5HJ/yx+2
KkXKQV9sDPY+w1CKEjQxSxWiTxhzjobch5RF11tBfh/Fk4DpZrkjtPt/GBHcikaa
IeH0Fui5aqNd59I/LpQDv/lXo/V0Pw+aBkXXF5elasaTds2XjfYmOuSi7TsuELnr
Ny938AbccqQTf810nxpXIsBEDBZYO8app2nGjqd036g9Scy+vCerztfKYn8d32Lz
YLF19JtBMJiEhgCaQrSInJbwMUmmx9frTODWCsmdmz/NnS/+QvoRAanVwZkuw9iV
QxEG3Gk6f4bxLXP2VDaiEjPr74EcBQeUC1t52h93CTsf7C1LSHgO+WNup8FybmOJ
6P41NuPFUih+84mz6o7QfcTzcf9UJAFlXnYQgeEWEqoYy7JziAW4NASgQUZkrusb
cE53oou18MF6gSPE8+p9DUjw5r8/yF+TTWFH54jXZxmXIwJ6YQqK75HGIVIAjri/
Mg9k9it/mrwX7C8qHlXZ/cfMPy8GrPhBwUt68fA4loAVt2S3wo5/AEOUMymeb6mT
uqrMlBpokw501CTssMBYjz2BM63Z6cztKUjuqXszVNT61sL0nL9VBIAD1uBszbQ6
gs67gplaqitwU5ywF/sPxiSTH3DiBMRBl6IVfR79Pdd1uxkttkaKwmuWBTCUxkgg
4NwBqS7vFxt191RIzEzVpjo3BgyEtW0DakyE6Vw6VUfCXfapBNubZZ/SdWzWKsSc
6ij2vTyEmQWjs6o5nuwueO/rZwJLjIsmqAmmkIIr2FINNoTbalizUyNS4k/wrrlJ
RuTDM7IzBUxeDa/pnHfRoQHNJqbL0UT59UfAE4Ldi5QCPMEJ3A417RYH+1rrIUc9
tndxe1lzSfXN72tR6vftvU1qhclRTZk8tio0kF1/nViYXO/Dbesg8VZBBTOCC1Fl
7X8d82B6uB1tlwifKU82WX7Cx0aDfUk108UMn8XzFH1ZXl8YSOCwm5X1YiGyRaey
rJ9xOFc6xuH2IdOnY98QGhGqPwxncyq4GMRIDex7OXHn7Ck5hIKw4dX0Foobaz4s
nAnETIIFhNTSvsFaw6v9Y1RdxW/cB5YVScEzHRrobNGFR9vmTi/45eCBtLxIRSS2
VpFOmGXcVVyAmzcK75iqHXCP4VNE89U6RRy51wIemAMhkOXxkWOCW2bJX1+hm5AL
NvJoUL0LP+G6EeSRzKLcBdm6OBApElL3SUR4DhmKrkCU2x27+Wm9HiQn7Jhwh4it
kmiEhO/qwx8iArFZVG1e7uc/Lu07IPle/fc3fYpxotbkK4dHsyYtk7wQDapgPvJk
uvGJvsjUKZKVmqgH6dwBGlN4TtTawtGOolKFGuUWOTk+l2qz2u6rrTapeQrCvkB7
tQmapx81ueTtNEKEl4Pdd0Ec/KSEbBuXePNqS0mXN9FV0VnfZXzxHb1dFmfg29Bd
DSzfKGLb/Oopg/UHr/DV5lxkHBVPU0mDXlMEFZ5QqgjnstaMO50SlsgUvyDKFt3M
N8V4qhqecHfhkp/CjTahYqspfjpCUBHEkvkMMO3LHZ2z58Euz5AsRm9T8ddB6rWI
jNXCd2Ru/EQNFYV2M8HpJBd40eqAngj0KuAM+lCMYHBME7bWaYmcz25lPL72NUoG
xN3AqTHrVrLkEcAfx9AVrBWDMKpNe/7TBhogFU2jbwC6HnbrgUiK3UCtc65qVPum
OEG++CS5oK9FjN76ftLlL/QV+m8Ry7jK8ldDi6qByTyMk18Mh4LOJAXxzyY/D7kn
Nkr+lefbkMqUd2eSfa6XiIOrwbXd81Mk9IPXiJgat6ULy65Pcs9EyApAgL2m5KLD
YnnqntHGqjJx2+DSInwVrc7Oa4L82jpwH6oVKhsXRE4KzKts/KV555ByNPIhYGkN
ik7OjEyYEIZYmHaM5zuxCz9e0H8g//nH5H3+fU8AZnwdSc0qUVSA9AKWaEfS8DlX
vrLMgtV55PxQwehzFnlK09/lkxcFDSdNKPCnaKtRP7iWcbUWbgJrbgi0OFgKt3qD
+xGUbCuiErzlXJhojq8A4h/cjaLxAPtN4bKHGke6Pjz/Ucbb3yVgkXvluHmfpXSB
h8Lz5CaZUkocuUGlzLZ3V0RlosO8n+aAFL+pkNHDHwNMEdRPG2HKrLSiQST9COJY
f3Lvbw6IDf6uuSfeFqCseXWKGFonPH1DF9TP5ymCtQpNf2nkmmn8Al8pcNZfxjH4
i4QVzaDFJxsWjYB1Xp0sZ8vhyqGAv8oYN2DA8Syzo7K6uVPAiZl2Gz1Z6gU85EU4
/UN/3YG9GdFOQFBuI+Xciz2hb8xDOJb6NldQ6EspyT03S/Na2nQzWhrsU1hBqfgM
q4txwAC/Mc83m+/A1dU/7WELVruot/yN7JyMkDVaTFrk0YYGr7Yrjy1NLv5Oyi5E
FvYszKtMBQsgAfUYj+wahNTeUaCjLaJNYD0LceVTYRdQ0ArGlKJIL4IDpA1dKeZ2
X+9F9BBG5gBI22M89iucUNSn1qV6+D5tLE+lXo74D8mkKnj9qBPEyMSZC/CESsnH
fB5yFWxBLv4hwt47362pVbRAq/tlJ/oW5pHh53vLptCwr8BGcb4sW+DdNGQiBG6I
ICTGbeok4dlPGuODMoyJIM8SXYlqj9x46GCT1+thvWn2/JCPuCgmWDOV7gX3PAsK
DEginOapgU1t5cd+Ypezi9O3WlcRaZB1E40bomXnUcVLXT2bFKYcg4chVjIVHu81
DDJpX4zAJNTT6CS6ZMnTbj+H8snPSPcriPjxQFkxXjQ8vSui3jxFuFcHlL3lmJwU
0bJX/K11WwdSEdt3/8dKAzAWD030oljLxE/CI4eKnyxxdYyrXzN/jyfxSVDuK/pJ
lzKh7HJPD9OMUfS9urOJObkhHHw7Hk0ZheHeCZBgQUTOeLSx1pWl5lMBdZMVL+wN
iO2BJK68QcTDLDkET2N8Y4rO6/Qx8XiZmbz2c1ALUr1qLA/ZFNPYuvmzSIRI1Ddn
m3e+NMBL8YlxMQZtdNNaLPqcO8A06aK9AduM+zvxndAzAo2Fa2U0GfEVQIPPCMmF
zyU4Pdl+Ni4wUucWoBT7gjHvVZAq9AI/y5NLletLjVjfD0kaDqVSBIGOdtMdXIf9
5Ml6YZKSlku8iarI5RZAHWIyZJUVjTM48iCS8gfYlgmeQjVZOnu3Va6MehSNSb5s
+I09AewZ46pOPuzhQaStvIWn1fSv373mQvRYmWjBJbbu61Vga5ozn4WebsWABshK
CjtuAolra0uEqc3lWeIA12nO6CenyWQ5FjISJ7YJfRAvnpH8GAJO0ibh3EFFJQXi
Hm3wUKpgL9NHqNvenECocpV+HUk73kmleIrqKGXsIDfxFFtF5Q7fVbY6ABFM6zw7
Ofhs8H7xGDlSIf/8wHww0LGSTHF6Ea+AZ3xfzsBgN3wd0nAJdWnVVvub/84LUL7D
aruBg28Uwr88QlMGy5zujtFFz8PjtWXOZCsaKjddzZshakce/BFk0e973Wus15aC
8tGQECPLtjGWRTeqtKayrEc7oDVFAFlcDkziB531/EZCozqISF4XSumjGvmAkpbC
Ak0bm7RZ2TailRMU+Fp7sUelkztpQoQH7b/47c3A53kK0JrjPCu6q8RfNilavSTZ
jQZWmDTbSEG7jwqe56i1lL02AsWF/xQ4dv644VEYcTtif52ilL86viIzFSU3x860
pNgX4300CHmAIZSpKH7tO/IdCUSysGlS96y3t4PkKtcr9PuQyNlv4IS+09WlTjij
13ZHVF48U7dcOFZIQmmo/wFFi5CwwprYM9pzDYjBekqHnuDdzAp9lpjv1vjXtHcD
Zkkslcf9zclHVt2ZXpV18+LdG2CghZF5YyBUwoyaxis/tsdEXSYyryoe+1Sxbrvh
hrCTxT2U7LQbkASHr2vAdy5bAzwdaQJGNicfjmaPuOMAV0DuAVVeGZHEoaZeyHf9
KBVGK4P65gNljVTvmZFlywzKZ1LyXNR7un89DyMc4TAODPZJr2teM3VRIckuyh5x
jsisWKyoThsXloTi64rGGL2TNudUPsbNbYbg3M4u77xLTON+hyUOH9hER76HMwIf
oFX53pQzgp/FJ3vKJzYiTsU+yw5rLgLEhcg9qrvTXIAhXwrBgVL78XorpO/zdvcJ
fT0ax0EeJrH7O+zjwoel18kUGUqth0svsUNxhrGPFiDaUphFZd0NZW5T6Whp63hL
tS5rvgH6MbTUq4qYDGFFuhX0LgbzLjnA3MLs+kN1XC+xHfbxLNRUomkLUPCQAr63
KuSgjpR52JfdLflfxUvEblJU8h0hqrb4jPHQxadm6XhQZusDMyobEU0xC425cmYs
W6gGnANUik+VYqIPcZ7NPa/ZXalAwtq7gqvKQqf3a7jJ1YPqwq7MISNfqTKBRl0U
ZTEOU/BIu+gfl/Gu+a742VnrFvhXaJhf9/bHDCYm8OuHQScc3GA9YBgm3r4elCvY
mBvPSRk3reOLkkcGVItCAhzC3Ex2gvG6PnkI+EeT3YDgMFXA3niulqLx+RlRd4eE
jdi4tbisG1AChI0kk0AXuFMBtakVeC/H0PS0GCPyCLD7gLyNea+Fwjnr82mXi96m
eHm8mrhBvXM8AVjMEHyR1mVFzFgzJHN5qAikKL+DPWMXwUObvnY8yIDJ8t08906V
SxeerNtEhKBOuq+yl5cKmNOE3IQFPp7MNwD7oCJxazB3GMtQQGcPvf3PUmX4/aKa
oL3sqMWaME3P+NSy/t0/5I4At6SxTcjHNpEGQuoTTwdMojgCA7I0EBxEre/rkhmH
JqsSwWzusqM+iKZoUS6vMIrNAl2VKhn+qBN0yFM1TVfefu5rH+C6BCLLY9s4Vvq/
+t8MLrmUiwfuOVosbuqX7ZYf3L3NcjR6yi6ZWTFdHWJN3qjmqx/EAgR4iwKqq/o6
jJySDfCAtCwS0Lk9/Atj9Y4Xkhwfrbkv00TAqc0kP+PXgRp5TFZBEZL6hz+4Yx/j
I3pGEyd687qmnTaIxyjsonN4TvUtWGMu6TU01A6xXkcWYZvNjIaB7XOE/wKqRtNL
XlUT86+zfMi8naG/q6YFFEO/iDGeU0dRKi0Fcl9FLYIEf8mzsBfP5ZfJaKeD5K4M
h0FLxTwvhPmFMbc3iat/I3iFzt0iiDuaXj+odjwNf03jq03h2GgKA4jvGqFDrR2p
AfIcYadDmAHUl03lJB2YuDWy09uVbKlZi9xuC4DACMR6D7e8l9ka+XRipkJs1vtD
btki2kRe7EZIK4WthSoakiskxY7PznpyMndi6THodAe7AmexLCqA7yrtTP5nYqZq
ewtnV0X2pErb61dvNq98bx4dYw1oROHQw0UGtiv3ck5yk+xyc4bDU8e7Ndjq2Xvv
MzCpS+SDFkWVkRAYL8U9jjZbfw6wGum9RsuG/mxq7bMeKkja6KafeiP8tTyLITFE
T1tRRDQbPZETzNwZ0eibzVgM1XFxqLYHsNW76dGdytXgZhyXKVHZg2sgqEEs9ZIg
ucLZF0VHX2c+3cnIJUpgIgn0+2nHgRcCikDytDjLEodpJVhgafuyLBdfuaRM2vbl
bMEX8Pf0pu8m/RIpDTOheu7kZ68PYPgWOoV//CZPyTPzRZdfXmWOqct4S9mrW1MR
vYSlYi09ATq4rGmidgY0wVr1QyU1ucezRfn2VQW/F0Mm2GOVk8GCTc/Jf3lS+ZUC
KsmF4rdiB9bxO6a6GoAszR5c66kPeBYMpw4HVxxSLcPKYGpggSjykGhFmVfDGLDJ
6cDmp/ctb8gRwEuAoiUKEX1FF9ZDHI0p0AX2v8JJNBxCS+du/Vf41PrcnPp+lKPw
tfRnTz9tv5t3mF5hudMC25yXxvOtpUfvFhuMjLWe97u8vg/hniE7geuDn9CWlMoM
oYjDfhTJTIbt8cLDdAjORAlPQPEfRcLPMgs8Rw0IvyWHezGqSrcxtGOwfVOcNVk/
aQY6AQ7f+R8pg96C7pgdB6pgcswYQDI5x7M14b7nidv81W+ELDW9uKqj4Ebf5Aab
ksNFPv85xYA4b0JQOtdpQFOFTSwpYOEHqT5HMyF31OwjEJGOrkbev1ovtrQCcI1g
atER8CDtqRBcaGihj14j3VSkMato3yK3GTMeqIPAJ/reSUdgjUecT7MIwgQhWer6
1gGrw8j49jca0yaXzRQ3g1+6NwZiTfSG7OX7d6SUXXx/hPKOZeluuLVIdfQK9fek
zIP62BXiSqGChnLpxjGlSx0sBuAJh/aS4j+0m5k4C351NxCe0fcgaVgEgs73b/CX
Djt5JWNYXeYxB82J4Z7EhiMzE5peeV1z1qGzRKdyMDLT+y51cCVoQvFURfZ2t+oV
aU4BXCrUGWiR/BlP5pjKwnwKa/asrO4OChoKE9eFJ0cfSGkOs9OmKlgT3RueFtFL
nEZBTKs7HSAkzqwWcmA1TIVQiUCBNWu3nLpBAh70wjFFKweGKGRhFhD1qMk1MrR/
DTDmY5J/atngnnAOVm/T3cywv7RX6KekU1AxjtcrBByIpAlKni2okcf1Db6eCAjf
0qTkHpNeqG1EJ/MS2YeUIjZXNUbVhGgtFjsGSXT6P1/UTxyVA7po9E/zRDhey+wl
vshCoMOk1empt7zytYGZbAJhYGAR13JGy+TyOmkNxYGA6oUZG3yv5AipeWzD/gtv
tT3n07HGDdmh260PBPwA3Pc9sUJFqT3lkEmFFD+Zr4ju3sX7iJEzhks8PP1alZ2w
VHGPE/TSyHJogJrvOv/Ccr2pR0ehhIWlSB/KtncDJ0seR7jOlrYhxlkpDjjr75F4
5Ots2hdnFAnjR702atUIv+cK1vO6XH9FBxCgNtfJfYMuj5sjT8fwoWJdLCgSaFQy
ndFOB0PtFazs1NI3Qr1bMwEjbLEnd/Y0xQCC3tt9hcUoDrZeHdHkMorJoKgqnoue
6Pto9u7FHRZXGcykfU0M9WHw4hYYDiBV1/OjJfdsWkKjubiCyW4Ve8LCBY4Id87r
dcWZuxIrUsZXlaiQV6R3PucmhSyvEBMxtsHarXN52NLGLOBYMCOaKbbdjyHUJhrI
hfc0uUKrls/bC5lw9AXkU6r3MuB+yCemxnrPp+xHaahXZKQ/HwVY8P/r2cATL9eA
LLtOVi9ZqJjU5RsJDvyixQyTEV9i+5ZZ7hPhBgbZ69QFUs3Fd46LztAAjb+YBRVc
2+phMXRv5ZsV41sHoLOPIS5BJyNZMOH/hjjTFPHNa7WSRzEkvkHkF30Dzk8+G+lA
qQ5otWVb7Z9w6DS28kCsv81NT0Vqd9pXDF/XU15IGDLSsevf6M+i8ZZEeBSMuf/5
zbLwhB14cHGpT/+3mL6wna/x0OKLS8zWbPdXU6ZlS7KlQarSs+3sy6tI5R+gXkKy
lYptOEKuxjTxo0ViS022FJ5i23licxU0A4hMB7+MOeWZDwJjW28UtcsC1Ed8qQZ3
TrZAsiAQ2HI50pQHwMzFUZRTi/b7QwQ5u6nkjq5H0NISldVr0XYP3Kx5kDGqJlWr
RaVb/hyG3iM0m5tYcjP5W9D3JHzoC6PJapKswasCCNVlBZids6SjfNIlKtOIV85d
O1poLDjMwJvyI9uASNQ4DWecbmvQupGGTYN1ExV7TM5vPZBbTy3OjBXBNbQnIKuQ
/gslXCsvdz3VyTDn1Fih2ySS3P1Nk4NetnLLm/izIPAHaAWz0uE/M89lfMJktoql
9LeRo0OgQQ+CuCxbs0xZPrTT/zHUzkroSu2Z7kk5LGHUhPj/p97LFNIywyc3opSZ
XRBdedfTsFRQy++eW4IVCxCdFvKew4Sqn5UXGnw6egqBGd2QetbQExkfv7N/2pG+
2J1caQPEHQK7lve4LKjjTJiy4sSqdUP/tBU46+dAYx569Sh5Srkm39pKTUi5TNdK
KwhV78+DGvo1Tfut7iM+HqN0ggOBi+LIH0yqw8VT8wyMq/1NmCU2Hnv/og6tnH9W
h2vTPJKeJjll2HFnGwJ9QRqeNDY8R7aG1m3o35L4ihog4ve1MCdIy+JvHrcmcznT
zNKi6yu3cRYttcAY16jyy68efExzGWzXS7M33dadTTPO4tT0RtNyLF8gj2CTmNPJ
sHCOcuOfxMrBuf5+Zl2966m+TkEHYLmNFegiNEQUXutn/Z6iy/JhOM+F8QN7YTei
k/H4kxtRLPK6PV3vk0coptmviwwLQGCwcmTBdL4wgIDmIPQnabx1CzjlcnATcJjb
zszpSwjgY6fnCHcyLgpwPUs6/Z/Hmg6rIqkGQTBpPj8UH6COa2rK78kCB/Xv09w3
KPKKBHvBf4SSMMvFVpZ3thOgiEetZVwMhmxNuJ5lR+mvfQQCTR9vMlQ4vqX2dcGf
YxkyGpSoxuWHdJH5/3PK5gzVJ3VztUO0s7Zr8jQMJJXPEket2W6R9sFjPsxw0vSq
DNIDlcZ5z6QTkcRiiF7S4zQItopUx7E4U0935kOC9TtaxrMIVfebq8/eFwF7JY3O
EACFzmKzU429f8hpAU4Uct/XhVvzyLk2juGske5IO+T2tzAP2qeEITR/FU0eFPo6
aOOY6kcrHoDkrX2P+oYr+0KU56AAbHObhWfsKa0LFyaNEQobhaypIp6j0seAFpa7
DuR0e8gpINeIIvhJMHIRGv3eBktwWJyl4wuBF+AKTTbRCyshwTg/WA1MB+FV0LDR
5SVPtUFAkVa0atgiDnkT0cABGbHKvexO1StgIxlEKNjOuciGV3URdv4bt7KeDdq0
EoP0stwvYQynAWWoeoOmBsGcgqzL1jHs5LIx8da/IpqGlbRYlSJKRaJiGuig1SBM
d1LXgcEXKjN8q6jWL3pI04OfG9wRi7NoXkoe5tl6czO0BtznS6bc/HW5BSRvZ2bB
+6KpCK6jaZvPpP6SOcXyhJNp5zqIWyzzdM0si7jsTTCzRcSbLecgVZQIQRGhWwC9
GMpCMdkx2y6QSBCIDCaIx9Jk3MdOk0n6hw5TSdVH6sNx/Rg5jGWA8lL+1eIkSJnV
0A8iG955KmVWB1nOOwVhLGv/8v5FNsGk+B3eOuo15Ecwb9/u7M1hnJwHxaG3QvES
/KCPHnB4Jm5fge5PbpOBYSB7sxXxx8iXL9KR3Pblg2IBr2RGk3MRCex/Ro9ddaTe
9Y0b8HjXZYa3+OcunD+NCbmwOorBS17af/8YQrXCFURWeHaE7WGhDtf6rg7ffZ/z
1a6xLIgk4sLu19hHe1QyfDoGO6SwXFyyPJ2c4kD91wnEHGcQCqJ8c10CG3GSQbET
mVsh+jINGdbD66F3/flOmE95bUiT0xm27Lm137oix3akvx9Jo387moalylXAHox/
s0HF9b9qjAQY+KknEcw1rhNBc8Fg1vnh0SIpQh8c+xwSjohv4HeYdlqFOu4bbqQX
DUVrziTnvWlNNKfYbFIiEPBbKjLMWw6A5d0c6kU4mVMih6oeRm+UepfFPYs6HUHg
/ZZoLtN5LuWPNpTl3d1UqTzrMqBo1ZjH7LhcUe0RJQDKIDoAHqv0pmK01qx1cyyV
ceNHZkWsdIT2tDkjD3Ctj7bdDHWaJa+E5UUEWUvZsUSUeutPUf75lRGLImvQEw2G
rBCZmgXBtknEt7eaT7wkiDGZ+ytjLFj718wxQHc0TrJyNYoxXUoBbLvLScYH1nmY
LsJD2FT6G90EEFTnuref0loj+gR3EOMBw33VUI9tFFLhdPpkP98sIyZtTGXnMeQY
kYTh0VJBMmFoDpxiJUGCTMELyCDDMAiPs3cPybrwKx9AdFI5pNVC7vJCyqvN9Nv7
NhK5YtIanHLQ1NnAuqBrUDQTLmQFs4CKIOkpPLPwoRfykKbB9REUvQU5b5r7I3Rp
cQ1hz4HohQ374q/4kgp/2h2f/0unkJvelhNYz0I+hcwQ1c9My7/1p1QdQp1KDmXW
UKvVF/obZEFUsZZJ5HZ6fgW7XsOgWbV4IxAD+8yO4fhX28AADdwmlEiRiIgv0YnI
iGEvdou6nU/Ae87kIcen8TfNpfktKHj6+dRSQF/KXl2lb4LsG1sUGiJ3Dh6943zH
LeJm8pefn0a7lEFQtHfnVy2zZ1gaVhMH/s1yP683ud3e68Kq/G6hiRoT+C9N0EtA
qZFs9c8Gq8/wJMD2JO4v5lqf6jQy8sYw67rqOY2fGySf9d9l79qlFf8HfYIBF3De
9MSnKgcRh7VhphKxW9j4H/a3ozNNZTg6dm2+sVjxh7q6pED8brV2xvLuKcqRSWkC
W6hOQy5Gr1WZ4r0k+xGoHMYh6hMt7SfAT7QqELCyQXWgBxUCiCHSSR/lpkx/vGPf
pGsGJI9/EYBwci8oGysbHqFcDlz+Pvt88+xi96QxEiGoLJgMbn4jBVvR3+V9Ntww
0FS4JVprEP40BStmFjN0YSv95f/sJsW7gGoIg3VSKiFn9XXFu1XDxHzzbZmhaR7M
pZTIyKTyNzaYq/lvYEY6AvD4Gdblx7Flt+jMUmjj5uVDLrPCBSZRd+sUSAYG56Vq
VOe0UCyB807UDXC0rPb4aVEtP1d4bZOMZJzlBW6fScSUoBxoVs5To1lgzk1FeiTs
i3VK2UoO3YsJw046dRlC7Hhshy8av+dt5ptgPjinJcoK/XtwbGeKv0nFVQjd91N5
zdYLryFhM8Nhyce8nGzqsTHU4kJEPA7dmH1fh39FEP1boEih5XFrh8sK90Tk1CeT
TU8ftg+qITQgOb82d/klHInPEV8p6+pk+U5xu/lFpqrPgWjbDIzZICz/wOHrMqbs
VN96q3OxLWHx37s2a5ctIRVLkGz9mBjpcnD9FXQVj1bRvVtLtzv4Vafyzbd0Svvx
SUcFXiwDPUNgu4nZcyXtFrKbuvK3rUxj1DPRSS2ym1VNiNXF1PQfyC8Xxavzgi9T
KyaZK3XTHXO966hW3eva6ivl7iCE7si57gogQaPKpXOfddurnani63jWGZJMTy3W
10Wj94xNU9b8SsnqMHEOiJbhszNJZa7n92eSPTP5kKRZzjIY3rnXByT99QpNiXwB
pmnRT5Txv2ErV1b/cdd3vPssnrpKSwwl0iOAxgKSAgCzyTESEOs+bVUvPZfiaw/L
NglnQHhnOvgT+g1XJ3G2AGkdYzsk32JRsgJ27YAym+HB2/fqWdxBLe7IRQTvUn/P
YB8RwgCqXbDTpWTHJJ1YdUBfg8RnCR3W5CAlxcOiMbwtosraqoX28UjXc0+KVFBv
4kph5vwuYXwFTPekjr15UTAjo6IvhyAIQpve8l43mXpAUozNhcdfQ/5i0X1T0AxT
JXSjBXqgvKbTUINWSOVBtBMzZdtE8lLtUqAEGBED2RbOawHP4haDl7PI9UX+OQSp
PqSHLuO6JraVgCTJuWpqwW4SrPAdoqOYh/cjvUoQWPqL0genh7RX7Ev963faV/MC
Uxtw91bCsMhEv8Y5nlBNHwcPS4SRKrbWVF+ErEMw1Kp/EJnhFEHaY8+SEaFT/ziZ
qpsHtiXYbdhZsQxSyiJN9pfaMFAgSgD5AnGM6CAuQ0DNu1cU7PUh71t/akn+aoAw
Tqd3nJGLBq+cxl4XY8N2vt2OvlF6EnPmGSfhXYmK1VSiYRhjA8yh3H53ROy9cLJn
JgT7Qxv90G+ryv9VYy5YiZcZOT2eWuvEO/AlGuUjHc+8s9057dBLz2Bqh+YO1bkA
6JNMOlhp3WH+vPULgGAHX4y6qqrbOAWxRlRWQJWZ3wkSDrCjCfTeFNgZjRNOt0W8
zFh3XEMnANfQemfEnHxtLXdeYz4/PTtHIn+u/Mz5MuS8YTe3cDzYkpScoRBG5GFK
e1ZlfDiQqHedegZylu9Hj2lWKe/S8lKWjsyVn62+IIHXdbuAJuLFC7CLgX96Hbd3
rplgPlDMAlYynyPSuVV2ubX17piKDZwuLJWg7quuD7OwEc3W0XTfAM2FYF+KIMTc
O3tpHaieeyWpGky9zSo5BZGWs99Bp8I7t2XvcsCxeKRLLkW8KYioumZIKFXNAwhd
rhAQNiwE938pwagZjhgoLPb5UvFxlFeyCU9iuUa2ELTvpgOCh7Dt0oCCUrwX5xgG
DonwTan+QsTbTE0L36lrnUtKFOSDgEN7swjVsJ1WsrBZ5L+uuLmZXiMKadwPiCsD
rdbWTzEIrKluOr3S5zZZyqkk8aL9tYXC8NoCRhA3ids+Cn2EZ5irp+ZTOqRU1ZOU
Qes9ms3rxuZTVk9WX2xlIE9WGgpr0vJojC01JHpkB1lDaPk/tIAjtpzTaB6vO2ts
zs/QPgAWASmnjMrZCUBxCoBaCGS7LE20ogGW8G6V7LAkGckRQ0wYOscXmiG3SNPk
872QLBgfHZVIApWYTx96B644r+meH9ZWAcLMnAh+O3ZfMvzf8167q+X+aWSXbugV
fBaMSJUROiDlHSuQPhs6KtnQT27w34tBnQDqgeHoCTvMgwved6jm+66Sck66u3Le
NphAmAGMFPUY45quTziZdK3oQc33bKTN0sRrWawagc+BfdRYYyK0EXwyjQjyAg2i
3CFgNosPsDfhXkyVgEk28tX9z5BwIvsT9znJLt6DjlVa4bOf4kK2wkGzDXFqBoHj
FXZrYtOay3NFYxOYpyx1RVe+QXqMJo0+nEma4Gqc/ImIPAveFB3dNEAAl4Z2n/YY
QlubGq+C3QldWGHAaQbB6kpHnd3yuvi4I03VQ0nN6q/yF+F66qz2bTaD2v7LmLg/
95MFWiLiH8nIi9kv7JGiXlj0JjA0DZe3zOQe37T4A8KWss1ukn+fJm/sqdAmoH4W
ZbvUztHOeIHP+TqRA+nZeF6gTOYWMLH0N56ncAyJ+JFDTXA+6afbQHRfXhh2kGMz
8evMqYfInbyPrS2kAdlo6ZT7XT3bRE1bmL9WV2hDyGQmmb69f3Tgdea/ihChq8jQ
b+KCEqta0rHpnnIyLOvtsMQNvg9TvY5MiJ+LWXlaAZhrcIEMBVUAughxUvIolft1
y4ZqeN0sEOeQumw8gmpHhtAoxenrm8HKHPwJvcFeinW0Xx92YGnJwwCSnp5IXSUv
na+lQL4NzC20MdjyW2IecA4OhlLFJFChmd/NmhsjR+/w+XWO7Vl7pq2TW5epkEBZ
17ovS65NCBAHfEQmSJI7j/1+MeTkYWbqvDePUKr5CeIR54JIKkJYFJlOqiOoryzO
T5au9t/AXOXFkIm9I7mp1wVSXlZYp1DhbotMQqKQMFaFJ+c9NsBmARqnDGOQIw5m
uVy72K1ZoPDxWOcyS9EU68q+9UBdA1qNLQ+dWjKpS2DSwmaMOkHuHYWwa5c8kijv
an5Q28P8L70ZkHxF6aTQ9BnPl4aYNhpz7cGsb9L0bTYHJHa+FkLHhBsGoZHRarCd
iiads4zCWA3wvQIsrRwkXW9OSAtMCIW362G1kk2ABD8XMEi+Oq09dOqZJJG8ADQL
3R0vSEy2Qs4U8s7IXuGITZDwg/faEDIKAYu8/WOEbKMONieWiOvVN/7gxkL+Iq72
TkUzOh8G7ikubasjRNmoqwPLYGtvuFSxSsRCeTaRyEjG0J86jSOwFMw0yuGgHPoL
0BBbsf7jA5ukk+OAsWxpx4towJC1Si+kSptKTvll8fD6+KtLpC0tZx0JU2dCSoBM
RQqNwMCTHFFJgsR3uqa8t0UBs8EHkUImt1al+xPTGvtvBnLwAWlMEfDe7cAeRt9D
zmlzrLxtj0A2W8uslOo0Z457v3maW7Cf4TD1Sy+u762EGuJDnKkDGeZUOmohP+33
Dr3/6/pkHgT4ywMXOPDFQ1xrHsMmf9EWQeHBrkhra9LewE/I36wisiF6Novcd/ip
VLO7KhtxOIUUuHrDOmj3eod3GENEj3yDsYQTOWPRs5f3EpUnlDxSoxIcxTUyLq4I
8Q5PMksW+RvZIcV5y1BVGwW5Z3QnBkrbAIy2pqR3zT84HkQ88U6pK2PMaH+SaJhg
30I8ydudg015ZqO5IhIQ5UYPxUUpFEJRW/oUIAY4HDGMB22qKnNkAnOdpNogR7Yo
g+BSE1FDLG9HMoxLGcpEPEpyOE/5agde4GbuiPBl6B2A8XgyLFh0/3anEtSjK/E6
lJNBqNm6d2m2UcJ1/v4mYK+P/FBtJoPKD6Fh6PIlf0Smvvrp4mD1riRQ6tttJmCr
+o7ubEDt31u6qv8hjvvgu3uZn+5ea5/D0d6YsVutq7be3N17S+QT3C1giOJehqpU
UHvo2ZWi4/AdHWxF3VLh9MXuqlpgCzOlLmSnIz7tCjLvyRHj4rlDI8wMlYqxRIho
hTAlngoS6qsSn6X1/gzPcHB88gT8qFxtBPwi1zA2UBBlPU0kcq6LH0IEwHQrDknL
DRdjt2N6ecnr8qA/KepSLu7Z7hNiwrNFhwte4yb87DQzgIc0QDu1y4nOKa4/91IH
k9jGQlmSth07whZlw254WrD1QjCXUOV7KkYgOo7FF1TPJ0wuxWUofNsQy1Ew9WBC
xGGIPnAaX1+nMBj9rM+70+THzGpvoj1gPS4ZkZlQwANiRixxaR9pqdUqId/SAvz1
2+g1HXynWVwARL6Lo/Hp2395K+k2191PjcprePorh4mdlh8Ta0Shv+yhpKm+FdEn
CZVcjD8i4jhrHNucGElNTZSOqr/7szZaM39gTxOuEkrHGEcp98J6WZT9B0GzZU3y
Nlohk7sxehRqTP3+vmg4gP0a9/nfGm67WoLvNjcZHkPUpzWrkQap687scveWcvQn
wD/ZPJ9cJqqmxv7sTwma8LoXIb8+fIYwXIcKen5lDLknLyaQ3NrhkPPTbZzt9cSJ
vBmUj1v7UxDSRl6HZQ9VYNzDvDX3R8YHJ0kptH1xtmeqyWNCAZmYvQnViKn0Ph+e
GB1gAIeaDZFFx3LoM2ujmZpVmWIThw8Q6jiNPY2833tyEFhwmCIqwOAll3M0CVNx
or4MIrHdWBUfaxNBRx6PFhn2qyay7sYjiu6byQzd33L5ZvC0IrAIdUGGb/yyflqt
Z4xRpNWLN0fssyWoXQHQcYh0Xbh8exKTjqk30U6hn/ZFLIHVH1Vj3fs85G3JZK+e
k90B2JeG/0BprxjN7oQvRfNi1keRIZs7ml8//V0ADBgjIpzz63MDyZqykJAtub+U
Mro9J7oF/baM1d2aLnxoPb8qKKFV5B0QawcvsvK4z098MMIXXozCSsCRN5tDtCZ9
zYGn8EDY3zntb63GIVWG2l1RHQuvlveKkcUXhBq3AihbXcwmQQylGlmGNnA5QwhM
FlCkoPlLLnx9P27OIBPAWj4e0zeNrXM/1QEOi7yq5Cb1lVIij8sTYB84y3oCp+u7
BFSEeIjQUMhCJWHSRcRthvkZ5cn3wO2LtJ72W4Jy4ypJhViro0NGd9kLw019VtdQ
VAHFSYbRp6qC1Xvs6Gs5+GSo/C7npjNSlwHg/FXJ0UHBlvqa8AEEnURRHTfZvd/+
4vqWgIqnYn2n9PQF9RSgrPTfSvCVCz8koAbyz21tRphs8xVu7MpVmXKu/5TU0TFt
ztEObTw+gSKG59uTcCjaq1E1LVpbGgs285qZDB+kes8DDQBQiwUSD2jey+nuJVkA
9AQQDeE2PWV6KYg3bPG5gg0xc4Of5ikiU6n/vPaA782khXlhDVUo7haZv4/NNo99
tIesWHrVpowTWVg/Nqrb8RsCHBeGsjuRQWKc64F3x5vSyfV73oGI2KxjXZbVGiRL
5FvkCE00BysrNx2jQzwwzMdVUJMvl8xkyGFW6e9rqoPlORzbYCXGQ35RGbqLds7r
3wS6+Gx2ZjtJe2vgGxhL0yjeGbXQZ2VUgp63LqNQEFrQosHWVq3k4TTy6rfRc/Yt
8IEB2ceqOulzJ3g09VxULwqXIiFDWhYEWehQHQ9T29a6stGQ9t0Q2o8CdfBxRpOw
uiYc4GGf+d0w3UAVm96x+je9igcuE55dT8F6/15lKJ7Q5RengFa29P2rdG7xWwLj
JaMk0+ICWlb+ZIRekye6TJETMiMhAyGhzonDIGE/DF1UtUGOUe+aJkcf6ML6QLer
veJl1tVv3Fq/WbUzdQDkWpKQPFWtY5PPQtvRmDEQGCQpuSUTKk2a1t8CakB6sC6Q
YXlnKuNJqeuYF+0qprEgcuH/Q4uwh0tFyOvmz3AZur+BDZ02JBvocX4yOt3j+7RK
zAMGCiw07a2ZD2AyIcFXAaSUHDR2VbIQbwnSOemHekoiGKobprHVurpjvagph7lf
xETR6rj9a175EHygW9L7wqZM2DdvYJX5iNIc++wqjCd2ZUmAPhn9NkrQ4f0yK9Nm
Mg091NSCRjBibKKYq+sO6OI/iL1Ue9pc67DsO9cPbZaEdDYSoiQkRSu02wdqdRP0
6Xn2RIbv7mC5JsT2zEkETq1hm7LNCIX1PF/4X/nGffMj/ylalVb0I8KflGXRpIr0
cRmOgIuqHVHLHwqCANfonMYcPskMcfft2BFd/KCwv5CZZTHbNcmsiKJIXyVxSPJy
G4yBayqbWDNM2PDb2Gg0repaMqj8nWP4YQ1RGS55QSXoxrdeN445y8xDnaEgdzX8
ehvxlUANezQ3OplDzt9XuKw/FJH1L/ijhf6vM0OHJs0VpX5UGn4nmFFe6blr688G
wKmt/joD/l5uFw6FF+y8b6LnCnwQMaeUl654ntOuJse7LzKo32BKvPSDYQvv5sVE
evBoOKFfcMh5I5im4dGcDIghujHPP6wbgHmlAyGw0q89M3W/mVFHzinSG5dNNGDs
2cUvCypodG4tp2I9t20NQM+VJ9gnyG65m+d6h8C9n/vil88WyN5m/Bcm6Wkh4rpc
OsxYamfe306BLydpuh9heliYbj88f2C1pFsAMU9/tbzxJL0s9Zbif/R31A+3vho2
nP4gaSnG8FdyEEKWEoAKmZNDfUnHweLkUE8tiYnjyhHV52xRpCxs/OoRNkKkmgZ5
Y8o5gtNwI4SQBUSZ41VVZynktJ7uD15ZPUjnGcdjEPhe31cWEfjjqs1ag69GWE4e
egzT7jjOlzTzLarPAhdyGA3DJQorM5VaJbCXITkHODT97KeLhySFbeR9ejqxS6aJ
bHeutkLeP5fO3pGTkDYxOEpa3F0WrfP7gZQU09C5erQcoed8Arp94l7t7kEZXYVe
WiftuwEOe20yW1RApE9ABMUEeOUoARnFKyu86JSjB4PZEbfjU+NERWaV8y1uQzBh
nVDDyogEbHRcDdWoZZOrnFeXlgDol6ttFUtDOGa3Cn98ZPMX9j50G0TrGKL9V/fb
nDWhH/4j4vLb+ECRieVwgWznaK4jEyB9AUC1hUaUDWWzat2WfM2nTk5kv0luX6KP
qXf/biC4XckhLBrxevsGEw8DnuL5yE0WlShfxAMcrjmv//nW9xxlCfYz4gz9hyi3
NGAvIck2xF7Z/yY13FL2OXvvgK+Lnk6+9oFuwocx7qxdQELP5V53wpPy1QmQ1XvM
GLSaIUUB8P3HRZN5LG2JIo6H78QMRwicBkaK17DhDknJWrLRy6fjGDtuMUDk3dJU
uHF+OjoKBhS2eMX/DKbfE/3tBEc7nn8R6GHAhuqj/mljJwYlExRhRJE9hWhYeQ/0
V0GJPvsOc+5RJpZQt7db0lAUUVJHToAPlf4NhKBEZpRHnD9HssfS163R42ek0Ilg
0/D7YK37GdBdChiMMZs/3gPI1k3/3kUovxWWg3BjW2GCK5pICCmKqUbvPnxQ1txI
hJ5A6RmGhOqO1SvX+MAf8MQCZUTnkNCit0BpkMXvlbN1FtN/S+9XONntcJ/IcGpT
VHrl7FVcgG9OWCdsupDQeW8hDtGmyvZYA6GYkED2mOWwbJttGAgay/6o48+ruOrM
LzPISB8UwQlSA1g4u/b/CLX71Zan+cvD+Qj8owQkEDozRjnjD19eZmAJWa2YhOeb
tEcHucjMHzpdEXowrlX5v9nQkUvSQdlSxbh6kLpU9UNVPLlyEvtpc/tNgrM6BinL
sHpsxj20jVuFQzaxmbCjSS+C3lmCM1de82PWUPzi5C2eKuCb06KmC8jJcgMoDL6h
ZIouJ5sifWVOoiOIybdAKafZxDzcqK+6ET7Ba2O0zY3pxhyxsNCENPfeue9gmXok
BkZVhKwQPmWbCroni9oC1pJLHb7JFP3FHn4mbi8cRbQ6A3xneEF59Liy5EhOCpIa
uEn70x04/qY0EsIPGMj0x4Xf6CSr4ug8W8ClYfwcDt6hZo3ZtsMtFhG+D6J9gXXT
cL8NMjlSR8V9JkPIx926TCROYeVYM+YjvxzNoXYZRBvdP9WS7iNtlYbEs7kha9kE
97Y+6UocuJq0mjn9QuEmtcALlbCCd5LPm4GPZ/cgmQaCSQxd3g9ZNsHFqTMnwkA0
qoeaOdPfgd4UIdWrTJzWuLlapmfPWq8gW9E4K40MrinLSlRwo2i8lYxwCOv4dkgL
zMnYCiCU9VxgTa3sg8maDRamBPQt9SZLODuaRE/t5dyCWuzlYwMQfmJ3ii+EF95/
aa8tVjGXyKQZtn2vVfPibGNG4B7QT4+zfuOd9eNbrO2XtU2aWuX9e2hb/9By/tig
MOHefRbr+yS3RWOLJILJpQCZe8UWhSmxfK+BSMHg8n/14WsAOY6Q9gioc/7Q9vWU
UQMVf09+EQTNudgBNnMDs5okg9x8hAcB9pcBIe2T22wa4U1qk8ZmxxJP69B8f2rC
FDUhygePY6qXDk6QGq2Pp8N7jIGTksCnhLnGCc05DPniI0+zwRZCfRVr5dgeInmm
EggV17+T8D51Pzw+BlWizAQmcRq7UxJsqKsTSjayDBF4EDDBUZW6R27dUFKzgI1F
2qQ/KjDxRuJvNX/pcba5f6x6/Sc2HPz1hUdd6aF2dG64ZST+6myDZSu5hM/h2bo5
aMMpYvcXHIsxrzgQatFIqf+ReElhWXnS66Kv0xa8t5sJEqoa/JCfCObdFR21X1C4
GXL+3J6jnKz5Kt5CaJMBOLIO1QqIxa7haiXF0gomEH3nUbH5+RfZbgbUAhJsvMtC
lqNWcCZUmFV/cMM2EPNbX57JMkiIrqXA9nqvEWhJrZ0A+bMG6oYmhYqV1xAIJkgF
OcVmVxdOl7QQvSUFY+f5CesoxBhYYccQgY1lNY3iDhbAuhogrmcsVAM6kgNnURUc
DNxnJUTyDfwhNhNCRAW3C/UnVD+hZKCrO7LJiAz0S3DhIU/xQBeVLfQrihTnuAjC
c+w7jB0XI91rACgkrpj6P1p1yXOlnfJPw76yWeDfFsWF4Gev5Ck084l+9XK2raXc
EUlPZz8BFr2nmHX6i3DB6muimbNzbCVPSnZ5ClSfL481+qvpgLXBIzHv7pF1m0DA
UfYFq0r2FQK9nrWNk8WRTQb3TRRXjViYLJU/3IZHtCcMZmb+uEq4Ne1oEc9S8XoK
NeZpIjNhUiZoJ9sxQsXpv0cOThUyz5CJGjuS14BWCSLXskzA9vYoiURlmiG7u3Np
yu5/NK17i2Tm96fAH1rtho3laa3RVt/sfI/F9Ml2XlJ7S82F3oQaBV8qsmUWdAnk
kTzy4fLovAS07tgef18X4oqzH7drNBJnZCesLuTq4grnoDbZzS1TfbyhzI5U3RHx
Q3NdeZT6l3adqjLfZhc9/L6c8rYVqlRcLEVNNvbH0yPUrIimQA+eiqnV6RG/eYb/
Fo7GjBrWDJlLmSX1LRpRNhZM49P0IORN0Lkg8PqZGJhPEU3qS6tWPySZtRwuf3+o
2uJmDtrM5yev060RvwbzrergLg3Fk7g9r7xKFWmC/BvKtS/waIR8O8Ttd4A5J/Tk
5YnlX4y4iX+8da3lgSUUJY+sd//r4VDlwC3CdPVwseTaSDBjUebf7KTtnmNZKkuk
lSxcesplIIC11s3Qcl3IRW+YzNpIPEIXB88skKKyLbkALIxcp46FUSvi3aWfta9e
1tkeemchttI45SaN8/kFQMznSqOPF5eUBZxInD4okt4MBeZsPr2TG6yBUqXEd8bR
jjWAWs+UkMsdarkz1lgmTYGYlsxgwMtoTXXdK5VTKDoQjsiOT+p1SbUXKKnZVIFf
UsYkVhwFmse4F7lWYZL/p95FPc2iykMkeBpp6SbvsycsgEv92e0Q0a3va4rproUw
4wuFPctobCDidD6VL2sRMl9KnD1cFvWvPq6rPmMjjWe2EzDc9KShtUUAb1c+x0mA
mPYTWh73xfy71sbFTe06djuN2Zg24ayY9sVFCdxpUmiH6eKiaoxxseOJzwOwulNp
aIlkY7TGJz1HjJ5AjX2CF6qVNsmpCvpTgXMYAKlszlDJejBAkbGoDKiKwVGStHmb
d2EEz1yZCNq0Fu1J5QD4KU7CzUB8hGkaNcWvmOvpCPq5UHykLfDhCHoZnMhNgG87
lqO7nVt62IgG9V+dH3/FeWDg0+3YesyLaedLw8OcEzrHI0KPsR8N/a8QfHSOKa3a
qOcP96hojaMPbRWNjau06Qo0GgaAMg5PAA1vzmAs7VJQRtJjEp0Yg1xZJF0oO0ww
SOFU7cLGNcYuiaYU+gXndxSkulRuJMv7AWXwGbc45sxtB7li+oBr8ZZknPOsHeis
eJH/D8+bJBAhWF5WmOqEnTkg9M6g8SDamGRmhUMmne/MTzQ3AcPI3SGHIf98sSec
0JkDQoetq3NU1zn/HcZDK2sI9uaWp2myWes+0JE4Ob9Hi2Q9PaxApJK8GvnQ7hWi
nLhx188l9uBltR54U/3olPWlbY3GxGbV+3nW6VpajBT4sSbdvSL0elzldxgQ+s0k
pq1nH78bcPZAT4VJY9cyp2hiZxjq1YVJRJQd5PcaJuSmzli2U6XYHn7yFPB0lo+7
/dqB+OJ1ldTfcrEE/GrXdQgA+WDT9wJoQ2qJa77Z+bQOX7YfZnCL9XkcvhGzKx1R
sQFl4c4vKHKNeZLhymci1Y3jkL2TUEjwqDFg9Wtp8eG8NjQWQSbV3aC90IYSSSTM
rd61525gEVfZFo5Di27G+9n0Fp+H3Lt9mmRHmJkMe5NHHpfivB2CdsO4/pFYuSOo
gBRQB+fv6z6eqHbN15H8ve6TrHtpmeKaQyctQBjAXICCUTAvXJA4x2iNZL2bLs38
SmSPTivKyD0Vn5G/vR4QwG4FkVioSjdaK12WiQHWKUnTxko0+ch/VeOtzM8PgHCB
QiIrY5funL5Qle+8tBUcVVBIIk8ifNQLXfyml6s0v5lyvMomGV6dhngR9iCWHJh7
v0OHL8sXbrp2snkbXhBYCqbBO15XWw7NhvjGzn5Pk/Ed/0j6qRVzJ6m/KVA860r6
ifJvQkhrIYvGH90GqPK0C+AqJaIs1Od36u0k3jShsP/Dm12in/Jxji17+Yfldpm0
2MuBrJLyCaaSofiOiAgfJhBrMpCs1vtocdhjW/ZnUiZd4l1NKJgdaIEUJavHe4i/
AqsNc/yq8NEtJnpO6eaQTuIYX/x/dpOsFtmWney9NKLnMDwqtD6HuSgWZFAI9JWy
RpBTqSG+4gqE3rghgZjw/DGzJbG8xLftSuDeHH7rdtRKJyO6aP2k9JA1GBkx+VuE
NmEfNvRTSmUFMizqW0st84lYg1KUbGKfVN0ueekwMtvuS++8JtpSw57JzazHzo4f
0mfkon5e8ScM/kBG9rOVTxXkyrHJuo8nKz7PguB8C3nicr79ZkNWmrskCVen0EFX
HrQwj1j1VWES1XBxWQRZc7pQrqLqqHh9iyFTm4ku9QtVLVkctp7DiBkqQnE6gjPQ
rC2NAUB7g6MMg6nDv9uGSl2I2fhXMEtuTLDEKxq3CSYvGOvyqgm++5EUp66er+z1
cgl5C3GmyXxtBzu4UE8J1ZTurCX6S80iXlR/Nw1QkqsB/dCVhstsoVGsIVTBq5uw
lOu7FjKYr4leB/u04hlcTcyqjP0dkKKWD8p/LkTTMiE4/v67pLrhK/ZN7ZkFNoK9
sCIo25I3eB+gU/fpQk+1XqUnnl2ALMYfb2dJsO4bc7NymL6eDuu6TJ75q5h55t90
Kuw5pajRwwU7Cfh2re/wYDsV1dMFbvjAdEI/So23nBxjLdMncLfBbNnpqX2oXsJu
W71mMhDILU9AecyczddCVYsW+GZnPwwgFVmTllfSL9hPV+6EL1wfSkukXw8d/BPG
dalCLPvjLpYdlpzAtfDCiNMRWmxDZH7CzLidPSAiUnZRTVtgbTx3JrPkETn+fOOm
7QudaH+WUtmMtivyczAK2TTyk6aaEkN6IUInbAvqIVO6IgZkiS2dLgrId4V/kXKN
b2qyl9CsBDjXkMcHnbWX0o78knm3YerH8jTGpacsLP7lx8m3/fPwp/snslyVXYas
h6B2c2wRZuSoMXnYUVb2GoZ9Pt8hdLTz0sxb8bjkOPe2lJy+5k18UuREtFQNdKP5
UWnNumk1JCsYjJFcuMllAsrTxt8jUtUT6GNfy1ecKfiIPkPdsBp4NbgqDjhT7lM9
7iW3R5d8M44DBPIKag+o9esXwr0AFjgY/MEKg5CmxRN+4IySPijs7OxruilccGnk
jnHCCungXxQwckgza/GiI6YG3ggPxNIzDW4++yk65uC+giqxE63UnrpVPHLaz89A
d1XKFei5HQZ/5kzf+Pi4LN94jr5A3YCydEZOKqu1udNuyMhJGGse7duJvOvqbcQm
gihExv/TRw1c8uaLGuweR15UxXd1J2hOQmalu5i1DuqY1vadt1zsfF9xNVztpMsz
/2P4zVpvYyxjt/uibnTgFyjfpRakqddingyZvnHojnKBg3KZDmfH/OEBiiO0yHpt
RM2kycYSIeUcM6gpMiQCMCDSEhR3ef45ix5nmNsIFxe68mR5IGXFkyPbJMj8Jyh2
TldeY3hmjdnbu/RDBIsdbRcZzWieN3PF4jC3lI8yD109Rgkk4hQjshoV9jPuQoAr
fb2N4RTamDwK0ePInQItONSBYB9YqXujHvswTH5B7sHYiEw45NtCbb5+VYgSMcO/
EyGnEVvjip7Wpa/O6srldUyLWzChKYLA0v0KJbe4Nn+ffvlzCWzokIIgLvKllQiN
o5HSHEMGQaOjprB2M60PuXPl9nv2XI6cVjqG3E2hFngXKPL+lV2JQfWZqsr9Djiu
gxhvkZZdU7c1PjWS5YyUfjbroFxvWMiP4QzO5QgLn1rZ8jlQ5TxqKjWQf7kDPCQv
y/7+2EvOcpo9WEIl9FbvKR8GrXU4wjlhz9aggDHZ65SFjEifwtDraqI/xL0BX5ti
TreeDLheT4PlPiN/CdoPaG4lIjf3Ocnz2CDfads+NvZfAdPR0qxzqYaSpXZ9IbxR
oTXwSrTN4q4JNVQ8MXFY/goEhRNuWExJN4s6PCcj9zehmQJDbYg05diD6s8AlCEx
O2mM5VTltyoTM87LOLgeBE1Ykr7Z83JxBC5geC+UDum8gGz0gXTqVAqXpSndKlIk
eyIjlcOymrrwUMDUr2xMhAvbAOneVLHlrANIQPWylflpCCkVagiJ/zeAnNiujSzD
n4l/VUm3K7sLTmPbJvAotJersMc7vLEyILK3r78PoB53jRcACLlLd07LQ5OMqz4C
OQmnGI91+bvIEMK8rsT9nc1qCt5aMcYXXkc/jcGFzxBvOB3CJ/7AYQ6TQBGXrlaU
sIj7VKHsKOZi9zKJ54IQfeNaY1NVjRNSavrOvwv50ZIirnNCc3TyEmPA3j60vXCE
AEmMhKIcraRQSV3GIimc1I1oHQg6bHQGT5luqJtFy+tOK6pdeuMmtvwjbgVV1yb2
Uq6kCJdZf3pcJYPEj3dzNyQGmWuAhQP1Ya8ejIQjxeN2BccaAnhTjWHaPQK2ReqU
u4dviTWPL0MS52/yjAllBpb0LKJDvQhJfuHe4DstrFFTFIVLurAsYgob180wpUxS
rESxNOhoZ+4rnjIMhHz5g99icc2+/rmu/0rFk75CKkNsW4TIX84xldaYAmPyiHrc
WSZQ0neWOxhObyDcZ5avbWBUwGV8TDSg4gSu/Akg48CoZ0JOhVcD6kbdMcVaLaY0
HWZWrtNBEQoh3/tN6JvkaGh2O8pMAYeDLaczRS+ewXJdFc4yigjlDCtLl46gzFaa
bc1Zn73LxWpjv6h5+MkTeaTyTA8Mn/p4AlyNrqJffWzKB+ZIP/THL7M8jdgJOG7k
h/TN3G9sE/jUJX6kiClFYbxydF3RUEFpxe24sK28UH5yl1T3SyIeMQlHFNEf6q4S
s0D4pPZkeLNSxB/yPi0hGvBQKCkFuo26XejsKLu6N17fax2A+QsOXX1HahKz2oGb
y/iHni+HVqjqcn1160LRxE9CCwkobBF9Gp9ZvcmMwDKcIN0aowxrVTJlGf4F6+IA
Wb9VzSvZGqM5abmmin6PWQom05imbztvUhSrIPAQ6nax/MNhnsA/QzLcukO1Nmks
VhcpdQnO07tvUvIt58FvmP8WXDR9yrHyd9gEN6MZtEq6hGvTgB9Bj6ZIpKUgMUg9
wisQhClaDv/gXun85bn5M/Tlxe6J498N9WdyAJHpBbXd7J0Xs3+C3Xv+hORWxym6
hr1yAHuUeW2z08Dn+6V8bYLKZBOlok4P1htDl+1IdJodnv/Gx6MXkOE1LMO28VUT
5zc8snLsOy83GYNJeRLyTmMlqvsTidpHp4nVpHdGtVCBYnWex6JXwVqvQRIUcaOc
3CKPY+dS9nFfAi2c2og4o7lI7qeDYtkrH4s7IIR4yOi30lbq8H33WbmuaZSl7kO4
O43qd9tfogBAmJ/eLr+qvxNVRTLGgrKau5KVDntMQnIW7WvwnnGZ8LP0zLfFjiDQ
v8rsGZsJCvTx7KVFLB/2nd9xQxuDQtKEECoY1N7yoI8BZkgGk1ReOcz+nbTMG1eB
rQwBfShGQD2r1R6NwQ6rIMFIGbEiBQDSrzAHgwI/tczvoeqX6OIQfhFTbWml/0tg
9GJYlygGsCd6Je4QafKuTJKie69ifBx5oJVqlT7jAubTJMHBNHLrNjsdCqQmW23o
gvGfion92p0jmmGSnoF6jvTZPlojEmpkeqP7IA1TwJIx35ReSi+mfFfJ3GmyAU0W
hlzXuQJv6K1bkmpfKVhon1EuIFKIHJbjQSVgqHgsyOST0VghEzwCSOCEj+vO+Apb
8QgS5LNAIzr7bL79sFOweRf0Z8DywYS+drPpl8UZ2zvpkFdDnUXk9lUf5GQKv+od
rn9hkuJ2sL5ktwdNXcc9llKVzq2GcgCYY5SCeY4QfTP0yi5h0t/Sz9ru9YwR4oou
aDvJO7Ia3tweT8c6NQOQDRQy1J6mGfS5aFIcGyHJzMr/NA8Kst6uEdsLxcwNp44Z
pfteK+q6dVnOOsTuORUOdgkmSx6ixhQHrkH3XsgqmHK/AvJyF8zkxUaUlzTIpGyN
r4ttGXMMqiP/w/jgXtQfP+DzggBq8ptIx79bBZ/WMlyAw+P+nbaUw2dLDu+EmK+x
E3TVRRI9dZpCk11Um0yYb2BHXuNbhNvoH9ZcWQ1uLUzr82I59n24cGSPF51SCLZH
fm/zL09CqPcD9rBPfNGwKR/OVV542//4Pq0ZRV9Nkif3mtJq8c/iRoU2OtDc0Yvj
ydfXL974V/NP2XPXATcfIz6uDGZcso6IR2FFQ6m1InLgj1xv3A4hq6vC4XIlX7db
g3S+JPNMpE5WGMcVC7lEws1YFrJDARBKPOapAPSZp6YZZUmX9aWwNap57lklG3FF
/2zPIo2xVGeKvPQgdi9hG0/AsURusV6mDErhRi8Ct3795wgH8ETKuw2RHzD+FwwB
WDsxYzQJz8Dd36tlTLc9v4zgceLo7qKYNFIBgPqvuNmbn1jjsSMUYSmV97pgpl2T
1YuV7xx2P1wgYw7nY7AG46tAVnSjX6E4oFAbGO3MVmsMYxviYb2Pvf5rEeEYglDb
WbTZWQzVx3QDjcjgBlyj1ou2cDa5FZcIbpxF+GfA25QAT/6n4k8yFx8OQcxNJxOX
M44z/VcfmnCXgsaQMCMWiGieuU1ROyEsvEk/Peg+hS/5EEyFi5TIFK7WJJQKEtVP
pPR2oofazGKikTztZiDceSteIeN5WfUvOyMXEAgwRCWISI9RTaDs+PsRRAOOBzCv
xEswbxFGNI37hLDYA16pozuyH9mStTkggNMyY4KQQ8IKZ+XnSoRHPQBoj9V0jDWj
JJ32LAcmcU7Tk9uuS+3TsCKMbvnefRuqQr1ftSxFeQWq48qm4H9GBTaOBDxzZW9c
i0YYCJeoFuXhkZ45egnRO1Fdb4FjldudLKYN8b1T4p7IgadKhkaRi/zK2NHb5RCT
2dzFvJT8vTELrgNsdpsqgT/PqpVg3O8Q4+/l7rVi5my7trtuvEc6jfPc5oI+v8Sw
tGwrm07iFrtn1lAupn4IIZAN7B7d5X7x98ztRR2D7wbf70UD3lua5aRREltIW+d6
HJYsMd6j3jX2ZYIRP3zKTAiNPMcx3sKD2s0dfQZm/KZFN5ClPKLdR/BaR9H2s90c
+fFVqBZyUehJk3nTeuIjg9Gk6RvtxlQlUYArpdq1azB0qsU/W8NzzfDKtinkpvLt
7b+pMih4MSvAd9Q2bGhS+gAmxoR5zHWqaAwaX98CZbokNUhoZ/CBvQ9SAqwcMZU6
AGvurK1ejTzARHKj0y/4OUckhm22Gcmo7SvPiGDICoewljCrgRGVmMiCOadiK1yO
opsPyiB6aO5chf1rLvcoTz70njOl3+lbfedIGVOhf9FkT50w5PyqSNwQiWohClt5
yyGDMjNDn/BlrG257ItQZDSgLQu0Z5pcgpZUcOQZzTuVoPs+6ttJZ97Ec8UR+jd+
SQmlSbwfM1ehsS/bDrL58ZddhMQf+Tqr56TXjmnnGBdMjjKPY2SHyzXikuSfZnpF
QKHikLD7Sxjru/Ac/VNCpBJMkByeY7sN+UoKA+PEkOEL1hxhoE8ao/hSMVqwGzM2
Hzdf31YFcZ/yFNrRYixqIe33oroBovlkA/Li4LM4DZ5pRg9FW0Ey+UC8SCdvRBex
Li9htQBXNg/wj8LOBNFWwKrEV4J3+gO0tF+lNwn0POJtO5B9wllgkoO2bNQY8Dwg
fU5VqVMxtVu0bvGSPGcTFLsmxyZqA3bPWO7JorOzLZMLHEQMOlA9hczwWnvlQ2+s
b9ojILnczpBb8TRZnBBHHl0WT1W4LoTAuYqeSq7N6Z2uJdSojGNqKbziVeONRJ0n
Qq3Lms8Dcoxp6j4ycjzeIW8aBkTIQuSaVJgqWZWhRlVJoQ39POK8tvsg+v+WHE5N
kbUByqKqAlYvFkY4gnF1rpBb/Oc2824gEOhDs8uKw4t6U4uOZSoZj9p1Fef6KHoz
54L/i1Yl35EF+oFM/otC+K7QAQk5IwfzIxHe1mcq+KTQm1umreMpP03NtAtn8d1o
EkE7i8p0v8quFJnnO/6j9aRsv6QDsvLIevRSm6TE5lN5fL9byzQqvXGrZSomjtqC
1Ig/Q7nbieJnR1YMia/E5Hs6vjYwsF7JV1lSUeb/zKD0v4ShgLkeWPgCkfanPbvc
yceU/+lyH5Osu2zljH0hMnmXJ7584zn4k7uEXTJrJ7IawWYCkZwt71aEworxLwTC
mfPQCV1VuS6ehGomwa1oGD/ebPgcdAifXbsPTSMFQCPHzv2nUEUYu32zA991OUiS
Tr7W3Lc2ysIJEdiXLRKxde3o8GrFFoAiP8eEGKVKmF9c+RwMT3axxY9ePjpnLLaJ
zsonGQFdj4QFuPy4wEmMkAK/MHzLdr4UytVARECNjGE1cN3hr9aRxAUO0mmeRaKB
fiJvk84lAKElbz0h4gyH5MKEJmSdCA2fg6FtEBdytTusBUQ1RKkpjsPWfY2MGhrr
gh0pdUuj1um6X/vMlbQGOoQT7PFRoRMeJVXMKEjC2ZgmwnpiYK1ildEc5X8S3G8x
IJJ3cnINMy2nQ7RIuF8Yt9WW9QdzbHPQAThy/2VKXZi2WeUAYLQHAtw9UDvOBjwU
mwohTWmfssq4/SVuiZjVJ4lgdRCazMsj+45ME0epfMcajifM2FhCP+UxjJ2dfa7Z
XFfkavecDyOO1lo+8n074H5rzNxe2AJ08gTSIkjVZKHX7WPwUgrLNsWUT0etPHqL
4YpeB5dtAChszSB/m6jhtTtGlmcd7Z/I1cPD6XKr57bKYWb0yDyCjAPjCMlmkJv+
vV/+/ILohRf3PjkWXy4nlyXWxEH1pDTTE28xVpxYnEcy48B/Ntutwl6Sukudionz
89FDBSM5B/5N+Ks3pvv67bhaN8l+CxA+U+oWU64dKZpYuImd4Y4KBedeCQI+ginJ
ainPCW9+UbyhNMNCUFjQmZCJn/SBrlnfK1dNne0mb4Iz67Bbs89LCnt7vWQU5eYX
dAvX/kmEOl3VsBOOr1RVZ5uvxRl9mIw9U4PuYnCRmPjWGka5p0OW67Og+UI8RTMa
1a2Hx6Stws44+jXInCJulKVEnQTMy0OD6tjfYM63sJLzFsTxsElo5HOMWu3BwEV5
GQkr9JuubPk6jIoS9XcjjAvUorwT6hCT9/fbg/7Ipso7jOyYHQJYpHRgQnbYCJM8
FS33TGWZku+7qvc8cI+MBGKim5O0bL9BVXXDv6640uxSh1rfqkdoh9EzCpHSRTHJ
HRJOsVS8mCIXu8j0Of50WuDWMNAODrXB7Ndfg8oELQnwwDyY5kfIo+kORYWLZBM4
aBVGk+3dLDInPBjJHHNlOXmltAxtBzbnHIJ86LH1YND8XyFyIPWAqAbkPgQAx9rd
s62un9n5MDXRZTyE76BHWyzedXs8vMQ+z98n/1W9uNbwlsAOOH/HOaG3VqKumFEN
soV00+R1C/xpOvE4L5ja/sHifYJ/xen5zgrMSwLgx+U68qQ1cTgO20IUuEc6vVmL
FVvPChr3cIgBL/yOGAF4YproBWJWY0G5pFWDcertpkuASbFMU+8XYYAcuiUrXKrj
6pVrwj6x8urwauu09FOeTKSrBtPKmy5/GFmKLyX0N14HM3Jg5RMaylPb+TAw9Kt/
+VZZgyoJ4loVR8O19+MKmCjv93NFH2gk+eE+T+KW9ky5EJlL2onjrLNGPCa1Zamj
SmUHbq7gOqtmswsBGvciWbavtZpWCf23daICtI8zGvUH0zBwgZAOvnwbp/auQW5l
/aTUSp4okfIkjiYMUX5rH60gUc9TDpdEDEfW3HNoIkZqnUyVJOvrVNm9BQg11HHU
0pBI0sLUi4knjMTKv6oayueX5615ejlIJRjCL0MXPUFbo1Xw+in8O7uuS0GB0sXM
eZRCl68RbNm4jHRCiLzsimmC8F2LfYlmkwb9kIDv9vkKTxC6FVioXjESvMKac6pJ
CSdG+qnvkIC9RravCjo/Ky2idHo6LMh82+yDcfiUpu7mDkabZvbb3OmxUoAydfHl
WCAi5P5AS8MTvsNVQSpINzVOIUXVJtLiYp+CtsVFmUau1GwtD0a55Fk1uRQZU3Eo
O4tFYuoj3LIoRQ6WEjPRMh+t6r/IM+ttsOgpSQ2QrN25MknUMQJ/EjbE3svW2VMF
Dk5URadlOOmCvOKe8kRV7Qmu9RgdV6qWMgYMXJnDpAQGLYcUPTNcXf0/KUi/yZwe
GNXa1KgPy/5AENBW01kUStJ3MaOLTHeUcLn7T2Rf8/c4vjHbxkmPpN4C8JLhSep9
+bI49/P0+fcLUXI2I21BCEP+LVFI9H2DPkAnhXEMqKmEdIJAxyj9n5ICXbfab7dm
Mv8oLU7xeXTpNrhKw1mwVsRWrXcBVaj2XIGwVna1Udimw1lFm5sBtj/i0oEgC7G9
9P3qRyyKAi3EqViZTCApVxZTqHGuAFFC3uhmxC24d+uthjyvrZbykk9QulripiZ1
QQTpMbiCuM3uLaBYLSKVTtG3nda+pq+NvGGXhOmnYe495HJiSi1IcQ/OFid/quRQ
4enQhl3HL9ujVzAAtjgWLVqWWtdaEmxsKG45nnC4tOeD5AvLdzE71uAxPeFX84aW
P4kaA2SfLCrMInzFf9Xt/LcDCCi1/tcIxDh2riH/j1KfpCXVigsAWXlKq5oNmWBl
EM8KtLGZgNVaSjp+zP8dy4rAj1dht0xAquFagyD1N+gqw05gqMcv33d/QPiib36c
i/vLs+jKfgD90iXsaPlENtyc+CyBc2qZM+nQJUAC+mFLxDnksEHgCRC/eRIh75Jq
0NE9BDmCuPnJCBzjw4IkTTzEbFAPWI+KTNfg6XqOTnKRenKEgp4r+JqXTFh82Dko
zva+nq3mmBIPqhuB+WoxHb8DBG4VjGjc9da9UZ974MC/0SPC+Bq7B3UPM0llqI1p
2km2OAz518/O4EWuDir9ye5yO8H9bxU7h3uG6tLDRGBamBc6nqyZ5iiiA0wXmQRg
I/3MFyeZvSNysNaRClWPYAu7/dA8eoFPjPi6G4P19334MzU3OqIvdjDoIj6uWrcJ
IghLhN6nlQ4MXSBiMItCKmXLdc1aNn4qW2S2Zlj/J5n3nelmkb3jdhXUKaXWU6rj
/1ym00eyz13/nGBdEAgespYPd8Wg5I6yk8z+KfLv0Wbwzu16pEJTSUJRKvRJngwZ
lRKhB+bRSyD99A3ZK0taO+nUXIpgDPwKVE90HO24ObQqLmgTXwjK0Vrumb9GzGKR
WaU+S9CplZFh4Qyy8sFSJtzUeSVlsqstWsCoAIUDiM5n5itxVdgm/dinCEUd7Ulm
e/ydRJD9e+X4fmZcfV4LbN17PFgLuUdOqKRASx5Dtkg6hgYpF/pPN89u26LvLJxS
lzQ2Ruxst39x5XKZs/F5ikVvSyp5j32PsX8sv4Evsl2QxHBqskbG1kjoBJbUo41V
SoX/FLfo9S4JWFtbVdfi/ZjYwcN8mszTq8e8J4HAucY2SSh5J8x9JmeNym1ddmDi
a3Gm27bM+ndFnyY7GYnsZ6lMYKCqcx+9rfhs1JjSQnzvD7RDtTDtRx1qOdu2AgMg
p5Za63w9OtKlWL/3gdD8nCU/RmT2y2wBOc37kLKwPew1dhIqtMSmLTpGKtOUDPjZ
FvGm5WwwGIwgyELu9PYyyynJ2xc6gH7lf500RrAsexusTsJl1S6pYSN3ES3C6f3q
4iGIo/PeIBhV8yPtDVnFrqeiw3sZyXb1oNht/x9nF/Kfm9Zw+T5D7LtGv1AX3cDQ
bfWHyqvufsTmt0INciBuzbQeiYDZvnhpvdvsbxdbnhwm7T66vJzBgSPNnT8E5ViP
dqFbfYNXwto92iauoG3eYdq9NlNX9pwCOzPz01kpL597NYRXPFyQaT7RNvw3we7K
CdXA6Tm1Dl9m89MSlqonsjthuiv7zRhifwbCJ55DQcqrGKkK60cFF5QhI3iGLr/A
fdqyl06y+hKLaxPVt/3L9J6S0PmbJW5k1kfNOCkQ7nnDTPNrEnohP18qq/yA67so
9ZGQgYzEnp6dRsH1PdjdZ5vAyp5JSdneBfSr84btww0XQu4rjH3IaaI6oMkpHgzo
es9I+zx/559jxf2WXMBV3FIxB9nUzvjXh1nwyem61vBnWAi9OtIcvFeJq8vxzEJH
GxX2OZq2N/iKjUL/fOy43uhagqVNaBcEyBcAn7ErwdBQS3VLHpogNwJwLfjtdj9I
1RELHVJgke4MIRk51lEiCMDodmqRycP8XeK5j5TPvOc+Se8W+63NxUHiUsuOLoOY
j4/T6AVxXPOSCKGVCLGPDLcuR70hWie1ql0oVguFzwqdLbaOp95T/Qo6111RDG2B
MbspfzRAQDge/4Or9lhDMuXfZXXmrVq966L6mNjvui0Qc4IXojAi8+L+7VdMxlNm
2GiK3YPx416wf4zJYwiS+tf4ON5vcItWzk/dgse824qyIvi9lrKcr1T58MGW8R2a
f9FrGfkA2gIuOBk+stwkeNfKHCVSCjRSpEQORu+s9uHgQP54hEHyPe20BgYwRPp+
doEN1odsbHZyU4pULvM2ddwPlcVhBwYbiUDKRpTIQkhwDkVKCY9LpxLf185Qt4wq
4VYbJtbe5KwAhiJtGGsVTrzPI00ZhLFuzOvqLRuWaJQWZJb0JfVosDkzAetGRCQQ
gnrr9J/vDrJyh/2u6URy27MvPXl2Dh7kJLsEeWSaNjeg1qaLypG02VdlYrlzHE4n
Lhyl7xsj/Afa504pahvaj84NCWN2G3Rd8i8/55b2vxza3dmZhs8iVcBUBm+CfKFN
fwn398gHr6cjNCLW2VMuRtN1fusJC3lgH54vzBSTzi+DXDxpEDj4svUe/VIKkViZ
aIQ6HnTjA0Vv2KT91XgntezZ5tsKK5+jFWL2Ab3AOFTqYStqtNyxmO4+uTJt6fHp
guVsndUiEOouDNjlumKoYiRmx8qymvx+SVxTIVXfj+tHgjM0UCFKcl4h2xoa81E9
7oWM+mcRuXk0VBl/okKifR61rrA/G9KLTW3R/mtRXfWSIOi4lhUrIcyaP9vBXXMo
cBEeJPHP0sNDU85ddWG1XhSxkBQbEIvJBXBUmfbC67tVBk/1dmFba2B8lMIQz833
/GMzV5eafpveaRtJKtFdS2hAmnyXCd3rQLBAXHxcnilU3sjfvNK/+sLG5POu8fQp
v+5bTaT4H8615SCO4l6BNzNOupyFmuGmIckEr7FmqvGueANE49HoUtQE2kWRbLTk
VCNq6uebwQ6FWU3vhVKznTX1vs4lQkabRZ1xPDjS9SnvbJbOoZc38a5Br5OX0MRB
et4aXtIJ6WnKe7a31cUKWJGsvBn+hs6O9awmT5ozgZnColFl6NXlIbaf27h0fh9p
ovI3jef26EFEHpnvk6FiSA7fHRlVNsj+oq93MWICO68oMrlSF7byP/rvOqR+4r06
dIv1u1pue3pdkDISVE8vYjZz1vAJBU589uk6QIdzg/Mk29yyD2aGJ5+VNEgV3sKS
N6Jbg7WMsH7tLaCz6eBndRbkmbSBax5j7473q1pxxp5o3MMatswu84r56Vjv3sAo
weRBezCNIcfQCE4pZcwdnmUoQimDizwOprN0HXmAwnjh3deHhJwoWRra9hM2NW5U
Uou3atJZi9wCNWxki+LMAV/WEUDas57lAigQ8qxvSHYUkQDKY/EJDwoolfV5UkoR
qYS3POY/Si41Y7d12yh0XeabMn8W/8QOgZwaVEZEZxEX/bjXjGnjg71TVn7ocmis
Uw+5ZHJGy/62f5KhXvi2fwpNJR4ZjxL11+EY/5v2/fl1tL6ioVDYoQtzuKTbvj1+
W2kVLHVgSMsFfHGbAwm8BsHm33WKFz4FNnIoVAZXubbZVLG3nP0QsGs47WqvZFyS
KQvcu8xCxkBq0xHbJTFdhtXpAwdf44eknaZLOf+X7scgjS3OkhbirkFba9S7gu3f
Mpnsf/o6yNXe5Cov0vdl5z5jun73vQbCqGRj2FoXedFPRVi1tXcAataFnf3hTmlI
HrBNPOpAqVKNPykDoybcL8sYrQgoSlmRLGmCtFYOX94Wy4TLkG+EtBmdJfNTefQy
HwmGRfTQGFBKTJ1CnAYnBsmfACwYhS7gJLcPSqZsFD4Lcytt5krPdtQqMjanW5Il
Dn0yrKJrQygUfpKwNWjfIZ5pb/DRr08fhSLtw04AdnYh/Kvv+PXwUI3ycniTQCdj
2m61l7/+qx7S7wZ6rPSI3B8yKIGLZcHVHKXM1AL7osjg+O2IcqCo3xxx+7T5nN43
xZzgmNyt/+j1TdNONdNEqReXgP80buOxrNbwpDmaIEqsQyQF402dADtjt3PUi63N
aUYozpdYyXjnetj7jXr2ife0xXZprjPEFqcpMN6hSH4IeO5fKOJT9VpoClIM3EEA
4txy1vl+lPboVP3B7GZ6tA+7K9LHEWQV8/75bleK6fqnQrq2toSPgsGcoX3SXEEX
yaZM4w6UXxWKb6NZRrJGtmWaweQW4F8ltDMLVTOWHzgX2ZZqQ4AxHI1fNc0tlLVI
P/jm7MqCG2EwFOsUJzHrZ5hW7naxueMDwtUpJAWcjdOOR1zgMs9Tz5fl27q6NySD
//KFnoCwb8SEwkq6x32nLAIXai+s2kogY/TcJzPc0cbNDu2fkpTa6bjXhSs4fvWH
t/PKKKcdIp9tOppnGnDz7GgJCxatRqxcRCJv1Oiz2b8WPWaMQClXCdnu4+3oKaEP
Ac1MlA5p07vG6R1ZeecVObWuAGiVVRsK7S7ZjCldIAWunAihRNK3ePhkwE03Bppe
YPWCdYTfvcrVAVjxzkFSavvwLJOtMvsbH+O2TLo18g2s5dKz794ZzN9862efcZWH
RIzmjshfQbaOXdDEYfY7oeb6UW3DITbDpKw8cC4JT17vM60E8God/m0HD3WUTXhC
IDuurXywB4wEMSmfaMl9dL8LsuLAVN6HwZvt1zC0mrGjZvFzMEX6wz4KXf745nsX
Qc5EQFbED1Aa4/bbh07NljBMiztWUtIe+UhB9epvDNBpuiOCprziLNWRMZRbg9IX
B86ufMNZ8thhqeQGkSCoMW0CVtjEdnJsNnFAuTYFqoJRLf0RUmFWqtbOqkcgmtIs
NHrrKXFDoSAmwVWAWEALiIhKLA7ur6/kppgurjFcfOhrEyvkN3z5Fa6B2RwlYsTy
ZpWRilJtPGJQt5aTbEuiWaDwAK10LETY3hUgGsx3bls9LEUAyDCNE6FuMMCPctD5
DPABP3g7PreS+Yzh2NRpdP8/w2gRfuqXWX2OuOSzZBZ2q2BO7z+tqCodmChnRbvc
rqb7qZNdePYZFnazFfL1u+s9f/8d8vtrEm5RXbDhYz0Q1rcs9Fxwu3O/SN2jrM11
uIk/b2D5WvXImucclMcxNT+h7SgDjR+C/wurr9QMJGE5Slp+ZD1hl32A9NZOcDE2
MjHfXgmMLgfoEtXwUhiqRT5qMAodi0zq5xlnUfvzmuUmirdRtzsMp/2933tfwHoy
I9d9ekhyJoes14U/OCrFRM5x5rVxOsloZH7Ms2jj2xbkMw5Itxnt/mt917UdZfDz
NjWG5rh9f+b0OpIZIwztAsz9sbXh5YVC1HS4sGBwwoBmiottwVm09vk8yAODW0yb
cWyWgQpKCLEGUGn0H4gXngxTwnC/8vvDO1D0kkmlUF2rFiA1zKIDs1knElU8hydi
sz9tx7gybgMdW7Z8T0LukHocvLzp11QUlDOKB3HVf4uaFOVVSNmi6v/hzZT39tFX
2cIp0/ir3P4J8FK/4t0A9l5xURhxD5piQVmp0Y0VVD2D9332YTtxpogIuyto8aGS
HdEt/Z93f4l6Hs8OgjwtAlcFwiSstGGdk44GmG5RxvCIIYAaz7Et5PbMwiaK3jqi
yckuj9EF5RH41QAIHSGlfnUIEMlg1G42LfZpYxKwpaOjpBrpBGCFdAj0JPKHPdY6
bL0nxkvazVjlTERsnlgQwrCPR/cW9u6wMfRjxyBjtLeR8NjjqxcAyS9ZyoJCgmKy
ZePiIyryX00k38X0zDz4cWgDo7U6CuZvzCq5zfSjCB0LPoOrS1SUtG2gZxC2xAvg
gonudgBzLCJN6I4+A94wj/0nYLmeyWDkehL+5vitS+YHhNeom7D4/H3aBKSRKY10
E0M0VJJ1p+DbzqWcBnmHCLPRIv2y1n2sLpkb5QgiHFgjfXWZk926VBXZo4h7Czrs
xxXRFanjUlorbHWvUYhIZt/fZxn+GcgN+JMuJhgVxQK3wB1SajvyNLLmiBY1Kx98
VtQfIUNAojMj9D5aGwwgQDpdGT2yKIwirlYzgTR7vsLgE4RRtq+akr7aXpFrfvfg
GwWdeJVaSopJS20Y6EVE5Hkfc+NZ+KAqWEnKVUudAD0R9bwg/X08kAVmQPazZQQC
OU0lYxQlAZsm4Xk0D2eC59FRXjDzHDhrFJdAUzAXq8G85XvvA3Y4cJCNWwODNxz5
EmdyVsX9/t8Sf8qo7HXH2uDR6mEiuwBh4aciaD/DVQKrGBVpWE1kVY2clujotUij
qkKAFcwR/ehKAnt5TF/c2rp/xOrBiM1KrsYuksP53wSK8uk7sSoCQ//awFCSbRk/
1vSOxibkw3yCLutawkshEHlHwf1pLKTgyxBja17fLK9IGxiKSPliLxoG5ErIaETs
kKqBjXfGnhqjJfT1CYQHppsz7yEn67ucP/xH4BwjrXTl0gujdOr2MLJERb6NIpZI
V3hOXuNEcRW3zs/FCpedi4fXYkLOhzURbvaF3cWN0JVELQkLwMzkg5CTgpTt4lH+
bwcErfXn3SmJB3SgZ7udy8Ws+PUZcLL0ub48JZfwC3cDNbnmrwXOExXriBG7dEjG
T4vlPiRU2gdis580oqdr4wjqvfEvtTxqFeIczan9lkwewu0PSkrQAKzfzALw7+dA
YMv61tQp0X+g520IPFFf1zEad62ZGBNhBt3RdjEAGK8I+9uzLqjTmCV8I8xb+NAp
HcVE3o2rxH4iOSZO1yjJbhlHCJ2jtn2mcqtvKH5JXLVVuyjmLxmsgxrd/gi0mdEw
dgWioDCwMQ2gxQF/y2Awdy/7ZEW2tQAfVaRHFSsvjGxHx80XwSodpKloW8GM9RrY
l+oqGg0e0Mi9+mg6KokchE7gk7ImAr1Ee+xCkl9C9tiMryUA/Uce/TiRCOXUm7Oq
lj+BIDCIKNu4useR6xV9x724n8NC3f1VsOWDjvyiNRzeaEw6A3ADM1ufDehrLEmt
anf6TwVT3Qx01wysvllYE4dTVsJF1NfFqVd3jWjb5ijJg9qD0FxreQtmSFJWBta4
Fg/T1l/Rc8YpEg5iDpTo9aAY4lvUGOZ5lxHAs4iJWiMi8sMsbXxrZcFuVhZcpwHf
MXne9LPlgUmnmwqETh/G5mc7SRzHlnrIw+yUImrv2rj2GiYKPBZwPJ7XqDI9hghM
XsoEm+GR0sM8jU3aEwj9w8m2F/SYHPofOsD+2XtGDRIUoqTOUJTSjLwZudEsojJr
Q9F6L7gNWm+afWxFvplHfS1XBULkU8SU7gwAUz2VzfkSSVGmpduekpTVkDDAAQC5
0VU5cA0iVu/Iz0uJcRm+pce3TWCj5V9REGrnCjAA4Q1t/mVDZD9I/6oavHEeedUh
8G6Yjz/LupmsKBL8bVRlEVvrvGl4OCB2Tw8Wooa8MUeSLiAxkak1tD/0fnOssLTG
mLb8PpPcz4bZdQiwRjcNG3SrbOq1JpUXz3AP/SpqYMP/LAHO/g/mA5NvtcsiffAx
H5gHY0ZWBHwfmVmDYlx1eU/v27g5YVfX9lMYtgDd8MSDSQLIVV5K7H0KT7hIU6d3
/pmgsSA+upBSOYVsg9FjdnoXFFc0wodMx7WnJfcEfuRS70q8QIejfGH44HzD5guZ
pWEVbvzpGVlIoLtKMP2jKbAOiAAUrOUoe1SIaCFEg18Nlqy/lwV2xX/UdMQPOfib
/ZPpo4BNaEjLrukIkfikpYiBin5t4Bpt0g0JQrM2eNSF/WuHQ8NX6Oc3ynBMwf/f
c2VGZhQ021HGxJaDo+u4/GRwR4fm8zBm2rX0LCKLatDc8r131QAgMAPrZr7HdLt1
l2I1t2waZTn9Kuj67go77HFT7qrlCqCtDFqgtp4xAZVL2h8Jxgv9CbFYBV/I2x0E
yCIvftpC/TDn6t+tq1uz9mZha2LqsVl7O1m+Zv+gjFB+jCYQ+BTJzDqKtwxcPbwQ
DyflGbozlb6aqxGxICf47sop/uvp9yO9ENWcSaFyC5Hxgtbf4R/h16jxQG/7pmPO
cjIHTpwd5Us9XyaZWStTayO+0zLh0E4kB+e+tcGC8tyqaC68GA9lYTOsDDOwMcX9
5MV7LO4T4FphMGfs5wsCw6pbEgG5NDJGZngGH6N9g6s9QU2s7zpzM9YQAM6ZinJ/
xdisxoN+yBh3J17MSSIjmTUY2reBRQftyOwjieC15Oa/P7tAlCEE7YlGGu79Z3nK
L37LcWtu5EohJVw5qHDNUz/syKRjJLzUmcGbNhyHZUvvhoR3qpzAr8h5wEV/2c60
5QrY7B7QKhdfvLdereuNspygY8BkbmKQbpqf5J7WI+3tvBXx1KTWl7zD/N4zwUXY
b9d4bpPVohG/wCqjwJ1kcQBEhE67YWb1tY7zN1pMo521/6t/2gSSxccntRc1N7JO
yNdVSpTa323B2f3j4ti3p+ZdmdNE5SRNyDqT6Lb5JBgHHURF0hjmLsWc51u0kDV9
1OVq3/cghJYvuChFaev9+9U8n4gh8b1TGlTxHIEJlAHUaZ6/PIH+Jc3/qcnOIgh+
JhSL6fYVORGSZRwY2y7IaucQJbvFbWxpKIJwIlVkJ8YeMSn99JG4JUD8nOT1dCtp
pa7d6y6f9n8tVILJUDCRNJ6menSBxe1+GF7VlUJ+a6YLhMY5EFpm7WQf8kaiiEvA
uc20nUPujv4cHIDs+4pe92UYa5KOykCh7Vvl6xpDnehppimAJlTVaztidXnXitKd
0W0HQ0sY59LLFEnj5UTz2XAFNKx7Ed8vnZQ7Noyx/uOHN79IMfO8EkL9xechiJSs
sdXUHQhtMdKf0CSeGu4QN0CeYtikO29sp7iUikgTAZDQg83CRn/BVbgUsqyQJOG3
vGNhHyJauE0BjqQZUIirg+RRRTg6FE3DqsmqW+rqcHHS0gxaEd0vdDBiim7JED/E
vw+EFmwbDh6Q8U59qVrE09kh6mueCB4UxCGYDE7nc7Z1Gb1bQWbcp1R6BKl7+OrS
1RNC8EljJFFkCBHAh1+mlhhXJzgUwBjRM0+kRLUmmRksymtyR9XD14ZL8i0P3j15
HAgocfRdDGHsTj2f3Eey+IQjpXJQOdbVuqhKP95sFMjdILW520o6ZLFmczOk/pJ6
7OPBVltAXciJbLtT1Fj55OJh8+F3ndcxmH9eXZAoRcRaLhKYGoEE7hOrUKH1MT7L
tFGOFmjKqdCQRwMkF5zXKJsZYNdt+M3IVEmHOopAmm616BY3EUHeeOih3IdJgt5Y
hWE5drgUQOK6iV/QgoJN6O0BNv7OqAY8qestvf9xXE4SSaiQKXKheGRNRSbmj7tD
4hcb0Bmxid+okc06zGimOryaAmD3/yDQjzaQKeG15y+NJOYlTIiVoqHqav6N4o6Y
/icZ1j5zaxcYAkYcD3la6fjNqQoVvGlcXbgq0VwMkSExyi/FojLrPsOJc3G4p8VR
qtS+NBpSXQXkItZsV/sq0yAg68sV8JYB4dYayXSryMZOT2HPpmshoEmcOP5bt9yr
hpWsaUIu4bZ54QauhpjLKMMtbPpJo947gf0GDfdJYh5di/l0OoLE+t+l89CUryH2
wLoqv0ZEG+SlhwSmTJrqmzhqJTo6Wop4ZiyfDWWqohIhsxffQd2AzMw6U77916AT
ImOwBdMffv3df4ws0tDNUBFlAAET3qShTg3GILK86hOCEZyR1KLCB4RB/JaWwTuK
X0W5PuGM3Ob9lgnDWGk1HENCkREab29IhnFEjfa95B+XJSrHrrSaTy1rRhH8U5ls
5ZjEHuTT7jjebs2Ffv8BNauautUrYeQqXkEkDki0Gb1ZcLmL+bh3B5dkw40cFAI0
UKE9nXXdrQIw1k/Ifzu4mXDH1g00E7ZWlU2SsJn4gv7pWM0/zy4UUnWT9LGuW8tw
fUKRHH0WfUrjbbrbmbTNGcCAI2dCygAHsqS3APg8wDF9U3urxOCWcjiTeVVldQBs
Jq1o9BuRgGBReA3/VS0tt22dJFC43TF8I6I9jMBaa7MrM3cpASYtk4+EQBAZqIhA
nZZVuHIWgTy86MNccqvR7OqVeRZwyh01LE2X8H0Q2LN/vjw0aGFnXunOpBbcDncd
bpimayrvCgKqIWk0j0UKfEt9do2sOZqyX0jAr/z6dftwMtanRTr8cLagrUqm/9ep
qQg1rgcxpO7WLR1lTjH/yFrZXtC48It3W1V+hcXG+4fd/hp26PlEoPr8bTclzdtm
8uoqYMXYpuycyAwSLgp3buYNy4GtoZRnSjE2PwWEBYgqWj4o2uePioVChGTjirGm
3QsZ9DlwPQOjtFVOj7UG1mwq31w02V5dG1wsW1iS9wi9DWm7xg8plwiAN2fbT3Z9
c0U27uf6jAcZni6BT1imQSs9coUGCCemk3jg+eOh6lGCR38C8sNfejWJO6+Fnx0U
rPAoIz/1ZtTTgp0LK7Id3d4d1Nevnw+avvshl/0oenoBo1pE/LFAII7pxRG85S4B
I+BQ+qejLi7dEiu6rT/uVxCrA/3/YkFDSOG9RL/fQJyZBKOAyk348s3rUCU2x/jJ
jjAtnHioNfcVbFdpk/ckn3PMBG5WZNMx3lbxwee7OQKZ+02C1x6jke/LEcjt3QKZ
uXN691g76fYXz4RSsT03AdFevtmsHW/b9zNTiBikDjyS8ZWyawVWPcb5DB9oTyMO
OLfT6G+I+3xR0t6k4QChYuZG5ZaKGCgZCg1Zm6FYZ97fbED66spuX8j3RFI5/oVr
Y18sAJoo3wmxSPieFrwnxUFhE5EvFbemKFg2drxfEP6jqGtoHoklh/yML6RrLdUc
16mpNsKtiamDmto0Y9LSn5YHs58AHPZAjuRs8/AhFzbkUGIts4AUz7uUwlMA0lZN
Iitb4a88JECEJQXSSrcTYcE86uth+speEz98lxeBRDSp/OmOmGcCyFzIoWdS8MeF
qpm38+V8oX/9MkWUgUbqVa+fBnvPzSGBi48uZaOUGLtYwPToCPEaECf02L71c0oH
Y148HSgggHhZN8om6GrVC75ocT8pv0iUUUZ/QUNsg8JqCkj6l9xhPjY8GXN7w7Sx
rKj1DDb1Xio35rEXuHFvawKv5rt924cXffYv8LW7E4uDzGqOF0stxUVZX574v81R
M7pVaDAISTCRPeK84mURVEqRb3JyJW7k7ksxQQER736HxkJlNJcFmNs7PGk85cat
56RsnVgKCLec7PuI1cr8HqUxVjboTgH95mn/n8ocC4pqfkbsqkGTK9oWJ/7ZUHWX
MXSp7IciGSiyWb9kGmf29JjzGKuky4yeh1Byuf7ADSOxnLJXHOC+m5UoUPq0wJfd
7GCGkUNpgvCOS3YzfbAj8Ei7BCPzLbGjT9MkO6GLh5KnrE0o6CyprwPmLEXpQG6B
I61xmk36I2iPpoCC2ATi57wiHFXpHoOx+X8QynjBUpeb1Le3EDCnOZP6TEYSKnNl
YWjg/B3glSVrGzAqodQvzQZPnji+I43sDZ+8m8AiMvj7kx91apRoVC4UjHeWonbn
qeGdNCByHobCIcgpTjkokk+uEcAwife9SglE/sqOx4Dk+40D5EidKftxHr2/eGc6
j4T+uO92kxIsbSrTGcHn/lLCQjzKiQ/+89h+2BnQyEKh4fDx7V5+QhbBHRDRHX3t
7c/dyrhc2AFpmReW2fINoTniv9IZNYFwye0MV4C9Gk4CLOz/Z5Kq3DnU7R7xxJPZ
xu47qG7zCYkRLLoxO484I/JpX2l7tR4qYgRun50UjDeEfNuJMPp67wTRZs3IgxP2
eedy/DjsDCtWKuG4F4ulCZ6qVT7MMVXlzsFqIWie0SE/wsYluoO/PnfqqubbF3pz
QNRY1HnVjeDbOAcAL9KXSFbiErJYnD9Eoi8TwFbsrmPOEBW6R6pdCbQD/LMQL2Jd
+Sk/5UKiUeBU0idn4SIWkuco82L+k+6+Udd1/PU3oOPFGy38fKDqbxgQBCjIZg6l
c3328iEH2gXBGosv5VggquyptTXh9NVNedndCidoKnp6ajoKVPJOz8r5hTPkAZ7g
+A6BBTGxT/OndfkoPuCqBtFuFW3hvwqgqrIB7iPJfW3ykzJHTeYmLj5oLUZhKHeQ
fZIqXFEJ5nfoymmAsL3moQ+WbVRON/tOiWjrkSjEYz0fveWcGjPNYunzk2W62yoe
73PpOcx9TOoBZokmd+Kf2HV+qzLHoHXLZwzKxUNyYQiXp26s0ze/qtNQ/9eGsnSP
KjMgEqpQelrfP8cpZsEezAy1LB9A+wpBa5j+zez6nTnqLhSUmoRB17N/Nkxl2gG+
d4f6vR4/4wMK5pV5/Ml7srZOHvyp+groKMfcYtpNju3XqU2wgdhzo/wQdzNWdj68
6p4pGVBwjhnbUzC8taegveGc+r5k4q4ILDP/VQI/RMdPQSFMVk8I5/uAY8UBHL7P
H7tNvV6DgpwN5GZKZ9uIfKK5Ke5q64x7WaY43T52I5fc/HTZ6XkxzDH/DHUCAjSB
gorVFgbdXHv6YLuS+kH6yQSskfcotnp1LofHOVpBOSdHxiRRRbhHddr0D2fToj66
KvKFEMroCvw68hZCEM4REaHLMypy9qepLa9MpW0LiwFzH5kLHgYjij/StmPCAo6v
qzb4BRd2Gt/wabbD8UI1tFW5UUqMLUK7+sKANt91D2OO69cvxYFoOiVhtQ2npAkn
VlkeVtLR99UByQomYH7jykIBJ/Va/UsQLD8Wm8VwdgqVOUAOxl6llgzS57aUJ5co
mg9xallxiYWm9dN4CCDZxh+MC2b0HDmidc6B+IqJ19AJWWLgjUGHk3sQDKQ60gdi
3gy/91NM7MgHshdL6k9QraHESieCo1U5KF1IhRejG48nQdvUfecL28QYIOFVB54d
LDr2QK09FJ51zcC06e6xtjLdJqadbucqD5YZnmqg10+kvuFSJHw7h7PiHRRPS4YA
vMRin3eC5AdKHK3ILjC4q339ZQGPlePDGHScCS/oyWhN+JpiR4irgrXu4Aknde5+
FJeMUs2vKo4nc1HlujKgOx4JE2Jd29JVpn6xYSBDwuzMv+9vdLsdpXP3mVGi97N0
VbReXc4VC/dZNRItHNF8ELnI/zNeXg/3ntTNmcsEvLIEzB5/xGR3JJ/xP9OwEkMs
J7b4KKsS5rgCIuTyTwrarC1Mc3ehTGeqKfyJQZR5oC8tc36BMg7xw8Bh8rGxoK6Y
b3G12XJ6Iw6Bs94EcuswVSm98mxCyAxYpM8MYXImO+ywlAHap6l2aODzzf2zSNJ2
hinwg9q1HWwP1is2SqGzAfvQkInzUWh4SZtw8f/laLKl6gwlrTkVMCVKjamWiC/7
S9o8ZQdJjFmJ6pK1RW0iV7rvp0oo8RkFTKnALv4l3TPwE8vZZr6BbpoILQkQ6UfB
zepGFZFsp/eKwj21AfJwktZykYYs0qIzxUZoBN7HzNKmjktpjD/IldAP45Bo4vfr
JwEBGUrpISZYiRfcckSPqHUaPpKofO62nz+7MCu9C72rHZfdPs4jPu8Ww1FGmehN
Dt+K4bj1948gfPqrED5iljd7TdOFeeWYSFUSNBcYj5A1i00BA5b0et/Weow2xF2N
FXMbDxRDuE/OBGwe1SA/bUx6k6VBs254OEWN/S71BL+un7tbYsiTsS97bdBL01gE
gNXqom+lnjKfvRokBs+3+ZsgzKiJpE8hBynguH/L8uGwO/gAMnPlM3Lj8vOxwwuS
dPfSkpjxCjgt+ayuBLePaGlWx0An7JpDBxyLMO7Bpugn3/OoSEeGKsBZ65NdC+JL
M0/Kw/67Dhy0E5Y2MSND0HHGYEHPiedmvurF+43X0OcVw6u7sUCuKv0TTrdcp2Ul
8FMTDyMsXyI4ymqN4CRzllbMDV+G4CrBbToa0z16sDu7NGykoV8DlRuUwIYz3TwP
XLoI+YMxzhgzYe0Vf9MAB2YrHUk2t1NCDYGGOph3I3sVcgZ3PFjEZLc65tOZPOW0
PPV0HpyhQKOSbVbza3RL9Q8TlcwD5nEmyZHxIFwnPQLVSVMv0NJvuLmS/LV4VHue
oEk/T2kphpdiw7HkJzC0rKd5JJE1fwmKiCN2IaAIH7RgAkqD0VYPRdzn5UaGGO8F
OeK5UUt3mocFfCqrwAtWJeLF7uKve3neUacPf18yyGRrFTiiY6h0briXusmOW6Im
zBJgQrlRegP6j/tqQZhNKpg9dLZA70sYAu0Y/CAxtVHceyN4uTvvj5y3zQf+CIht
pz1QspFknNj3b8KdAfse+Xikdl6NAl4ouUoHVDr76bFMevisBhQJmKMCwddP4HfC
QRzr/J30x1aJ/dggfwulGyO0V48FFwbQRDk7+h67l2z81BCVsVVhxj269bikE8SH
9WrCgTwDRUE+XaUqt01Z15Yazf9vX8Mxv9eOvRC3wIoU1xDpuD18ptFJgJUSlhyR
HS+q8TAQqcYYYUOSvYLGdawdf7H5Df9Lr+hmbgDp+tOk+lWo4vXHpNbFUqbw197z
ge2c3saOtMh/zMTi59e8mI/WXk76AQI1/d/qiNlApZGsXhphmRIAKcs3zwnYqgPr
yxIq5AneIyS5Zed0FCmTXBbYfKMQmA5ZxTeAziu2mFxkfeyxNDvpBCI191wODQH+
6kqO4iD5k1/ccGlB2l7AyBmZmTKIn0ivgwqPw0S+QnepPZjV4xAknlbx5sMya3BC
VCI0K/OwTxImU0twK/v08CWNiAclXMPjrN/PyTJmkL54znX1gcYg5N/pVpPrWdVT
XgbD1HxUITh/FyrU0iPLwhJaR3B6dRN+AGL2/qoFTwEJ8kr66m52QF3uYTXIuJfr
5Ft/Bv4OA/eEa0BGh6kV/yG7Gyf0LsOxuvC0xKkEoWoqnmftXyGDlFVuvJtrNpJa
0dz3+7L1yDl6Aq83c57t+OgtOWtfwCNle+ZJDpMRXh80D2btBSTT90aOmA1R4vbc
owdJfmp2gR79Um/tTD+7byinjM1+g5SHimcwYVXR9g1uKezcUzliQch89ASP0uRV
2b5go4wKFSa9cR64KVzcRaS6H0hgdFQCQfRvbLaCdyPj9u96lNE52layi+9N2de4
uI5529yRyb34z9nFoVL9q40UzNTkR00fswSv3dv/wc137Y6LuhPoTGBefc2FSAHG
kiSN+u81fB+32SYPoIOtQcYDOm64EY6a5k7Lovl8q2/1uySYMSHtGxRIcf5p4omv
3b1dpB5IQHG4T79rEScKf2mYrwP/GwDL7Yb3UeXleg/Wqf+PFPa1OjlYmLTzvCga
GmYsot6FlkjnPERXcHWrlPazjWukIHWecUuOR2u1jMGBCG6OpDNjQ8qidLCVAAoE
1or2jclpul/L7MGJh25K+0IpS2zTDwFR2nVxrYKVPAmFNtR/I2dfCzNHoYVpC2mx
3wfiEIgMgVyqAe3DLIt/VboEebeB9wbNsSx8s8DF5AaSHBGhO5UCqV7dhfHzGdgp
Ya9t/MALBe3dxG1P3ljIsE1BJLT1N/1X/jZNcNTm1g2NKmIYl7IsThbpkK2XWs0v
A8Btr/XkM7lBl318ZMMIJTFd8kZ0IPmrFmuJYwFaysCHdG8zlZhpwJHqChB4dG9K
ZHNLJiuhhLfifX6cSkoqYgOfmCqCMMvqhcoX8/gly4vLWLqIv/G8Jt57el+9cyvO
T5JwrthL1BUeLNcjgyVOhb9HzzDdjZJmG/qtzFtYZcxr4AI7jXbhejEtk/GYGeQ7
L4ZX111hHngmVI22YXI5kn9yeY2h8geJzoRT7ffcMNM8SLjIcXPyinJtKrnN8ecW
pp/5GLYe/qli7TUnakQ//rWenc7rjb4ENs1wKdPWoSDUgXHXdr5KKQt34xz1Lyzj
jn7/oWm2micIJQuQkHXW3ae+mUzbhxrLuGKlN3In6bVt2gVVrhG05D0aOCAQO9/p
iz77Mzq/ASEFeU6Kzojo4nIzIv+WBSIRhGOoVDcg6jo1fMZFJnIVWVaO3ZdlGRbz
brrQzLTElF+ws24qmY/Hu0xXz42lIPwV1DtbhBBQLQiOBEJj+VK543K/bAMP3qrC
Q3J86/OZops1eSwUf1ZidjvNtOQSvuvkKoEKcfIOQVnwIWcuPKmzw5sN/Qh9X5cF
PN0+3t1kMRqS4AFmetGrAexII21/n5xSUz/gAJu/3Sis/kUtKG6o5mnNHL6XyPdw
8+jwopKVSCdT48xVpLjs2zcIa5TN5xFZMlR86XZ3fypoTzjJvKKmxOJ9/uxl4CqB
771kiahMsnpU3gMHEMhdLlWr3zVk0oUjYmT3eM3C+x1ZxpQ2Lanl6tZHZNkGRZkG
dhMCtRcM4VI5EyL2kYDR99rgFN4rWb7lkp0ZJdh+gtag07M5M7s24VFNIAFABnR6
MmR5GKCPyVQSKPbZ0BZbNLDshbJgQ0BgHdx9ASrmMNn2Hzeb5sKlH5PsPt1vA7md
ypZNO7YGYwMfh4WreqbZXZg3hqn+YZkMRCR5L/1FqQWca2cgGILIOl2r3MIMnaAz
AHkabPQ64hSnqeyJ6h2HfVbX3r90sUxm5NH87P7PvZsswoML73Mk8o1xArkKxPIx
uwuj4No2xxLFQ93DhAM8uy6k2bxUkp4riFbU7AXkhcNM+osZjwNsq0LNToY4wmUn
aEJw67HrOIAGuziccJuW8DNWykv+WYV69DwN5AqN+cuSZ5BM8+KoHPnyEHRrHqKU
InXkGdk9M5GaAnEom0egLpPJ2ywkPrUlqT1wHMwqj/69VXYXbRMW1z0rfJIozZAB
2vZjPbkO6oRo6Lhua+hXlWxqxk9C3+jxnt3yuQXrJm/iIannE4dqM8rb2ArqwEho
VeAk646MqfbxUvJO1VTMNtUcNy0UgnkY6q23z3mKevCte+jHp7WqFLOE5qxuOQuw
XN8Z00eBYSfWNllkn5TjDsHvbwg3STd+wbZU89kQZeBURDBWZ2SAPlshGzzxEP6Z
/zqlpVaBB992OAFiF/VovGu3oi/0qLSw7OH6nN+jT62NDyllE10O0a7TTeLaAcba
zMB5SLsXz3cSCQfSfk6SCHcAE2kHOHGIwIHX+kcRQ0QKo8oR/YKmDjQdCLAeMDPI
FtGVUDmHJR0/PxVypHRpvg4M4n7MCvjm9ebNVVc5o2hvNB1Q5KiMtxAV/7ukz5GK
wfeN3QKGb8FU1H8j1vOnEWMqzClcrTI8HPujlr8a8lnSxXD54qakk+YZEP9TlZY+
As1WCHDi86ay4ViS42uwQEZEfVF0GZ3E+axasTRxvxv67emTJzrMh/29VIyvdri4
5431B3sNZIwbhwSqON8yr54wdFzA/DIPSgyHMV3AMifO3efbZz4A4B9jcNPJgxwD
3drCemS5AJV7oHtpnWDZAptumROPFe//xY0LmcMA93XNM5ywmCwfJHK2+t5y2Vsv
oz6z6/AMAmJoUC+3PmYNPmiyd7w+nEsXwl6STRWqAA4DVNbgdvL1R6RSAvLHenVl
AJGkYq9RCSabaOhi1aQ/ZbRLgGIAX5LLcWZTq73vPSY6w4kimlF+2ECjJe/FYyU/
f+whGjODnP0upo3N2b5vECnVeE7d5oICz05gefLrt7E4JTlCabvdOH6Bhqtnh25Q
VQnV5lvhXIcQVBDF2ntxurTyXMjSIBo048gBOiJI5p7IC/HMb5YFb/7FmlTGIBlj
TYIJxlbXk7l5FKLiDi8LbBFG1TtVJN+q8T14yrV7t2DToe6w4rnfU2GVuJMx4v/v
BP0awh83MsfqKLipA83s9tEEvhJR0/38jD0sYRA3ZsThfKaX+lAuzovWbvWH6IDZ
DgWyZsdoXbmxO0ZkgkS6LgiUvgYCiZD75gz8HrtdSfHc2Sa8KOFbjex/+5iSiN3M
82uFsGBCLhKyOmcHsxKHAYG8KzQzGUqyg8XqWeJz5jDwby4bIZyeqCNGWCWRb4Pe
Ob1mYNVd0fk9mA0yfBXLQYqek54T2FkZOa6MpZUfFw2mTOS1iCdNcS00fl9GO58B
BXOT9HFF2zA4jUvZY5haVPgBDrqGPZan/Kjza8T2OYXd0WjOI0qJlVjIxpeJhhF7
Hmu5WdApw2fDFKGs/xVM7v+KTLjcWIYWFFMDCvfQeW3ohRVjgDTvD8HL698UGn1+
uS3pNEhRoaaslbEPlu0bCuPzgDP8qw4nRqhx29WMLuKfifQ5YQNBVmMOLO2RVddT
Q6yvsDSMTTUUNkH/4QRSMYaN/cih6z4ElTqGAPIzrLtEkNS9F3nil+5yiYbVx0Uk
cm0/qU3dA4B+KOCptSvNcWvta+quJqLYzaEv5lU+8O7lsIK0zPW4czbR9V9MdyaH
2JuP66eCSf6QvXMzM3Fe7PnuuoFIqAXtH34L+xMLI3Q4pgvUHJgtxCxyU91PvuPQ
zMC+1TmLcjtNeuErswBNVDDR4rKTu2Qb0iMMXO8l2tS6eErAd6/1OKJuEoDkvSUj
Ige7PBgIKZ5wa5EphiBVXIOH9eyl/RVwAE0Loapb5JtySHq5NvdoT8rlUIsOoD9q
wmvHO3db/3HsIfbc9+KrGNHn0HQymKJaJMUnnMv7lCvSuZerXL3A+nSCBmj0CE9q
yESOkhdcdeKYkwzL/J/nxXdR9lIOW/Zk87+fUvVoXt1PrZovyrkzcG9XU7fxNes3
6EiR2A9hKVQYql8Wy+8wSsPuQWbN7R5rWqJuZHG8kx76Y+xYAFTe7q0c5OPfh3v3
26stjQza7S+tedBEd2nd7T/i6wz8oBdilbmMVNcqq0qSwCyswmagsrfKh5APAY9E
cSana3xNXH2OdaAUNFcg6/j2DwcgdBJ40BJMHxi1s5hRpmBDaNfGf38uyW+VmHun
bYly86QlZ0x+gAvuKuw60u/teN5pGhEutLE/0wdPtkCN3UaThSMaQAHxUgxzwFK3
kY/zXrXnkEgUp/iUPGsAr+8YOvWC1TmZBLJK6MmpQ8IIhyYlB6K5f4X8aQZRfOQK
DoZh5faDQD9xd8+c9n9bUilSyzKB9JacVf5edN8FdYRDG/xVT55aZIiqn7daUugj
b4xThqWtTwBEITqi6CfnQo5NA3cxgLnL5+UuIv34av0tbwqoABsykNBXYRIZ39ob
I1rEIy9SH08QPGIsPQSZEzIlLtAADC8aK2BaSQ0XNbM8RgT6EEb0OVQw83dGFxf7
0PFP5Iv5LcQusGz+gI+ei/Er0AEbfhqItrIqBwCO2xdNv5qJgOnwAcOk8q5hqH6H
S8inBajGIX+D8ZhV/maLKBnxpl0HPGbeBOpamDHNNpoXFc0u3lMdkx86wugXEd1B
sZZ0kV2wQHODe2u5YqDWQ7eUydnjkpmjAw5yWdO5s8t0tG5SSJkR+cjtOMR+mqlK
smhv5+rc0mQsjP37mpOgwFLM0cibfQdj1xMx4/yN//E8D5fGB4CaoVG4beMRFHPo
cdy22zI0uK+QV0UN1+s2FDoCTPx7wCJhQZnwSTuoZDMQ/T1YeEjbNdPfmVzO4M6M
aGq7pYI/Z28nUO8jZ4L1hJlk42WzfR8J4nomqWvTYLR9qLejdZyRO5OlJjdLjgg0
5PwogXZNSjnkwy2MEEQ30xR9s4gb1OVq6s44y0PvQkLPk7b2LDpUY9YK2TWEWImU
cU4icafskM8cBBgljj5W7JXfOuMoK/ktuC/I8BW/CLBvCo7QCF3YZlu7MZnpGkrm
JtGbB1EpvETf47JGSCbwPKNWMp++JSlCVk/aOZmfj6rQNFdxqJ3iR6II6aJZn25b
QUcCxJNhZKaQG9dDTlajJ+LhEUNy7gAi3rhh7KE+ul6+03jTAeZIP4Y46CFCQudp
1ypOplFUf7jknQFffwfe/j/yJgTsTMfZ5+WGQxbJG0wuaeOxzGdXYZrFyJwSUDDO
pug6rDK12td+2m7rxPnVC3RSrEUmNeDRbqRWqRwlu4JZcu2Vf6XhhvrdDixL96+w
QCssSlXNwYJLnKlfBsI0dv5cR5vrhVGnIFVY9bPWSNWqPv7m5/VyLE+GooPHOPAY
VjnwoaZQtiY3lHgl4JNzB/EKDQjA2UiBpTU/U9j+JT0E63MGW1Nt8eyo0Y0WyTqD
3uY6W8gBW7HU6MFHtYTsFBIf5CRCO8BWtdMjzj570xVA6Ub+XFNONXc/CqX6vy7s
C10z1tMd0sIrc0w9aWL80n2xLQlJoI78d6RECSkmyeHUcdSZZhtKav93i0cS8lwA
z7NZxSlC2ThwDzrSU+aIElcpneGTqNHGMa0jdbX+HsbcYt69rm+EW5n6KMSuU6Ct
SwfcQd/paPNbUezGcULdvSZmvian+hGVpl2hA2aEo1WX2daNpQwOKr3+WFvn+6JP
e6J1C/7t8FQS/O2zqkHb4d581SXefECgQ+aSBblSvocFx9Yj6GG+mH7KwRW53UFd
KOR6kE3Igmo4e6S52ObhXkoviKI4UfNjo3j5lxOcLtx1+a95pU/vYmlG6S4kTuPW
yaZu86d9uA1MlPWoKAWIm10/Fu9NHUCxdAbfo08y0c/cF840Jo7J2C8WU+KEh1L8
kuBneOLATBcqARNwMhGDUrDY4cWDXGR7PVObw3Acz8hMUl6zDitGm6G9IgU48zJs
JuzVE8jP/BXJzJrRPhHZrqIMNQosM7xwI5a/kvWb/rViCnKXzF/rLtEIqSWnvhne
eadjUMgzOLvZSbNrEmudUhHfNDGm+OEcOCzprqtiVrmsMiVXc/WS9SofEGtOs0lI
Ot4Fz1Z1mYlMxQh7rEUFW55wQTEC70oT4JNaAnsiMqYkhkyTdWh8LqjaK3qb+t/F
TeCStdLi6N8pknFfuXUjInD1jbwyLMsl/nAbtXstgM776xI5Pp577h3Zi08wKxcv
eoQVeqBmsYCOOuAqrdfD7LLoAAiUmCKpyj8SwBFn+yJCMEm+6UnP/9y3QvSC7gvd
hztri75AVJyp//hZdQnOyrZvMdpZsf9SHdGd65Nj8S0ItozYTpM/BDY4P931eeZF
sKahFPm4qxkHVFKGjohmrOKSX6TQw9tITpFjK4EosqGpNcTveMQWJ/VJhgFSL8k+
3MLUf6+B+sHWHi9YOTY9XvuX2MPJSMmAzyoHSqx5gedS9hXeH/I01yjUiEgMqjMi
mJEHFPm0WwTGjCCH1kHIpZzY+c06VKz/v7HAZl24Nzos8+MYYtlp1ypKDntEGEkL
DgbzVYJ3p75+Zs/KtjgI7moMmiICoVXlXHBaG/RBcxtSU4kpix9kxr19rIJiVQcX
BrZgpJdptmHvXH4A9EvNkKReevoEgbGxssxVjzbeIdH/hN4Gy1Y4rt91RPEDDcli
s7ZcWXmPjfQ2cE69Gi3ng6tZUzwtg+QQN9ww4L1U5FDHUTc00stpUNBh5BgNV3bT
wFudu/6oNYH/l3QUgMacA5jQJcKKH3eF5lxab2drb1fSC+UkEbr4aUIz5hKvs/Ch
88TDu8bfAn2IKLlZuJ7nxN0l0VqnGy1CQ9ctvghqpeuUna9TQl1OyYPZKGb7yNpw
QKjJ28KgOeW0nD9R/eESK3S90vzcmKCNfsZkjBLhrpmb3j6ZfWB6J+3xVLq+zotX
O7yJSOoUI2H+AIHHhK6Gfv2Su6YQXIPoTuMRuX1Wj6LKK7O44dclYi9CGNotz8Iy
xw1l1Zpy1mFk0B+Ovaau7TVyA8l4ea1I/6Qs1Jz897mDghwhMMlP2ldann6roO7j
CPJzatOGU8jpfIwgof2dA2lOzhqMV3U/8OzZUVvuTAGKhWJm2gco7/rXtYiUktLM
3zq+1EycOff1CKqjWQvXlv9X1h/ir+E1btTnHFvjmRpZOJWIp8JS8jj6R7iSoEHf
FTFOjEXKXCCbYH8wxdq7do+i2p1xOlGzXGjsvw6yQGANCcS/sORvaRKRdIlxVkZU
7UYDTXa6Tsom/ZReatfOyHAWTjYKlPf4QgiPmEisWFMNi//WS/urkDrthc2jBBRG
F3ey0J6+NlORe8hnSDECmuG2nix/dJzIcYJQ0kCbr4SUISl+rK3q4IhbphNr1nxD
WZ4dWE3k9yHJ8aDuxN1xc1HCIjM3Ho/VObwSf4lsKXZObqilvVa8K+n/Dbhz4/1k
EEUZIkUzPo3ppQ9F8ZXZicf70S2DK0v/R0Kr+Rt0vRxhyQwxJJOZqGyyA6eKYO4J
eDZ68kHkMeeIRWUGZsQxP/pPY5U6t086lOlNYipd7r7v0EEB/K6/OLdqg1/9blmK
7UOHuIc9uojFEKpIKeg2dgUK5VdCzzr9or5Bg/1Xl5ohpG7eMJyTxeNOjcbtgDRB
C/iZALWDdsmDm4eLhKZDRlPCjQElZwmGEc+6nb/fglCDTWShaYt9eAgmwPpusLOx
I0QSh8vK339QEvDZpYjoPqIRLuzHoZEYg1iviIIRhB5xeQKyLT2CKTgN69m8q8tD
JvcAe6C3MUwfFyP2eOBRp5tQYtQlOO96DB2EY0+kCWl+fAbAmGwj7ntI5EELg0SG
yi8q4FoZlOG+3et12zuCi3ZkxcdMvm079zvxzqNZAncrO+nJaO6qQfQblZlh9SqG
GcLRP7H06+0EDWVPTZM4JQU3DnjBQzd89CClVoIlaXDBxw/ZQ9cPxKiagzm6Q2dr
Yn6Cw02MRcdARh0d0dicbd4zbw8yZVhy9cDxZWCxS7aAS5W+cdNSOSru9CUPmh3t
ioeyv2WHZ7H/j2Dd+IcC9laR+x3pukXw7gFHXmsV+hPBORjt6eOXPehJNApIx/33
MqsBQWqTBLJhrCzhfpBSvOaPD0+FdfLLXzbAsty3fRLuDw7hQgD+VW0sF0js4t2j
QrCDkkpkeU62IBdX6soCe3BICoLqF1OXeBG7gnDcr2amJQnJRX4omN7pUcw/uusf
eZZ3j4wkLfJHHhdamCJcIiRxqDtAqayOp4lZmTc69VFBxcVqHlem5/axxdv/Zg3k
TZ6jLsEzbHn+Q3yixpyW8SBEQU1wPD3mdqXtDEP97koqFh1VwwxaniU1mlBcHoCz
zFipOU6raLdkgoToSrLZC968jrf1NW/ZHr+y5Cvk3A4afr0vHo+b2kt9IAk/2tju
mmFqFYVwcFGQXoRdYPLC2DaQaEp80zIZYko1R5cqUkzQuVMUC6PqxTrqrE9OccQm
CMVELmyAfpD6Ho8uRbCgdnCaPN9fRKrWyAjddZMU4hSH7S0pD1/RPm7m2tHQx+kW
mevdLwz7GW+SjJxau0RUxbfSTcuPX8egAkHBq14ygyJxObVi0btYkiRIpL4uRCvW
nDjr0uAdcUK3/9ibE5CkhsGisRIa7ylvcN3X3uS4+mcM68iIXqA2UOPfXjALyoHa
IVa+iX7iYERW2YMAIAY482ipF4bKk/QLbMjHk5vSC3ldARTh8glXcoO1G3O2y4nw
wLPFXr95jwNqz8G12B3jfinnQn+Wf01T6YKSZmmgZzmoTkOyGjn4Koru3j8cuaQ0
q6eWtUM78o3XkiaV0Zw6gRTKvYCw+6/oSY5dKpDlr76LnIS9FFJIJvEVgtKNKkK7
i66hANQLlMHuhvwrxi3UIInfvFslSTmTU2NqySOL9TnVqEMsKQF+oQZRt0zpICSM
FnOItnqMyGleC7F+I3Sch3RpxI77mzQOFzb/2GgmbJgv4OJxKsGgMkX9A8vCvPJ4
6Rysd642cX7cg4VXC1gpPhfqzZjMf7ZTtwqhNaVoNv3Yw8MzabU5Re8pNLpTPhh9
TMzmf3QW/xVMKkj4tT5xcANnWgI3aFbtZe7PX70cEDFGgtUC5J1UVWNHBvrKq5cE
xUS76NHgbxhLaiR3ZyhrxHzhdNGXjvUpQBW11BXUIsGC98/nuBrPTUGuTmyzrx+K
Tj1d8f7ZctJSJtCMtwqojSs/Uqrvaiy8dmf/xbVD+ztNijIWcR932RW8nbE1ia1g
BvMix/wyI7ab8pLWycAL6CI9dqYT5G+6PXSbbk6DuR26iqURAPPGUrTmXJ0+79GO
0wIlgKa5ZcEZgg9oZeJ3LjJ8f5a7jjir06tdPQLWwWrczXeRQjQMFcylzvP5r82g
BCBiek6vkmJrx6uw/GJbJvDFtaaPdkMJ6rNCk/IHLLY6sEg9W9jLbhGEAjhRZO73
CM36+lzjjcziqUVdLL3LvZGBSOgv6DHcpmmlIKz3i2x3qXSDUwuUcoshEFXqTMWF
Ne78UyEhAdQixlZxr2Ijf2H8YVjlgSYRTgaBM5IBlXimt0DF+42e0fxKUh/BGU7+
/ZO+YxjmtH9tLayxdiJb1KIRK8oipImDCw90X7W4Ty5sHdWFtHuFAlyAj1oFtVV/
34JBm0Ehmd1MJqTGwH/wWM9z4zuplhob6jxjloxXUVH3cKB3zCxaorJGBRFbyflE
eZ4LYtotuOj/5oVos0Q2u/Hd/tc4gh3Ty+dEHQwF208B1iJ1Ex23K+RNIAtAT5UI
g8woMhEDi3rpcFcH5+GpqWGCmKkzdOwJZtl72Ik+qVC50yuKFmtN5A3qAwtyoKgY
q+iAkYwkf3I49RjjB/Fc4/tiSj+tmITpo/Z3t3vljb3X+//izZLMbpvF3Hb7KkEm
/ebJ4BmFvhX5ZCll/WoWQWfK25OO2YTW+dSRtcxT+NAJ2vKR5Iq+uJQEX6xnIdvB
lIiuJyEs24VB3J4DIyiAyBgW+dQdIIEtWpcioWau5iNCJHe9J5/xDx8wUpRKBT0E
ngcil0PUULVtorOJ58+RwOvSqVOk8JNqo4FyhJ/FXzusQP42SdESyctX27o2P7a7
rjfpRMGBiuNRkh/ccPSKuj2jHjq3dxR/F2PQspV7f1vSjRLc8cH5vugz4y959Jjm
iHSHZJ/8Nmj/pQViKpRd3W85uXKEhFjR63XU3jgX46CG17NUg1xTeSrx2hjrHGDy
IIC/9sKxsnZtELPstOCarooUi/F8kaWGmNk5oYtOz3NUiASOBcILMYrCYzIEj9uD
AUKP+smcxps6Us7SLIPuciWaBF1G0u7fLzgWTU1GzL0M+tTiN82qpZ+dAsTuJUde
3C9SbFweex942kb/uwMtZ9z32Ddy0bKabQU1R9Lrc1uc5rls2TpSV98YRtykLlsk
u3XfNnWe1OqkbnOVUbhh1eF7hYUJVDjlZrz/C6NfNbJjEIQM0yn0Hzm6W3wVe+4Y
Ub2AJIADxD6MzvK2jA7/TmZObypW2+UBu5N9VP+QjI4W/tnkxwIRtKZYO22E7Hy3
jQqKJJYLmv+ZN/3NWrIEc5r+nNFqj0hd5TnDa0YBBbQAAtjPyWdtdKAWNjhM3zSD
J4DVnlsyc3oPGzj4paQc615CmBdcektbxmHfM/w8Gke0aTl3mxcEcNAAWotASllH
PJM/l4fISkyksOC4WmdnIJiAgUaofdsi/ViMNoMgvSaXdHPjUZ6LX151cNj/MGHr
BqWVuHCqul+qiDP2qTcHBr8vlI8rs6npPZ8sxkNHRd88wAlywA8Lc61OOAcqdBhS
nt69zzk1gWpNtORqUw+Hv8xWlSIWYleZz8S+jiZwm1XCK7gUYqiZQJ99iGVauw9L
L4wlhKdlyJ8cr1GKNBGwctuKDXp1DLEhSh4sobTYyl6Abl07skTbQuc5CNAhnERx
TAXXgjEIF1dndm2TBYPGahuL4sLBMChFr7lTMwcZZSAGfS5QauFVZ0OUAFj+zlBI
0kzZ+FUkmUUFP0O0T4/8QNtV6iFz/OXkVOyApTcbeOLstvB0fmpEWVaNUOaOfpZe
KztERCMRIx3kaT50tp02fz1SssB1eYVIsE3tqKYMg7gJ9aWWO7dxW8ykUshGR71a
8JUITRA5Tv8ghTiJO1RN2QbOOajGFwwM75uM5QUuIvEqOH6N6doRjXS+F1Jmy2gE
V2IGsMoGIbbOyHbyouM6h2b0CyXL0YrN2+vPUd1JOa0FY8ouq6eiomtqCYUdrpko
y4GqCPWR/tr9mjqoa/LWat/FVnY9JaJ9rC1rWX5uPvviH8Wjl9amluHkggTfy5c5
wz2tGpRDeNDF+hUhrBBCAsjzGJqbUK0bMEbpZBEfENt1UByW4rgQYzwy3PL/W+EE
i5OegjIcleLcoZB2neMnuRq3bjVncEG1r6qloGmH4m2fx6P3t3S2j+oGMARejFwq
L9AAjrQZ1xJR+VQO+bdt5KvPwfknSXY9AYwfQ3E+JX6GUzW91gTc0O+4zMuIaPrb
Pb3kpipC9CPSkveoTViB254D6l2m9BpVD8Xs9kXFQUClJIYIlabzlHhoJDy2brIY
OXHHduLTuzVcjJc0mHcFWg/3XXhYVoZY3PobClCRb63xOfpHFgta3aZHRh63sz2c
QyENcxkmyqH5m3GGRlN8PaZUg6+0lm+QORm7t3gc8UvgQ9tKGG0vsmAJfqnqIE/w
hc/BLGqqP+pH+Ophf1DKj+tDG+4Q6Axp+K2o3CxwaCTRcJSp+8NsORRks2hMciSA
dwDCAsZRv+PO6NTBb15BCU8maLSNpCJ3BH8zqGH9Qbl5Alv9SnWR6RZ3GCxYDIRa
lZ7N290dBmDaChf8lM4zZt8+odZwdjsi/CpfXTJu92k40TItqWCogqA6c47NPuqi
yuy0GqyGAa3MInSFeK6wRr0BcO4f0GXkMuNZQdTiHh3nSmVetCbu5n5qFuKFbIIU
pfWAW2hEp2WQE5wbr+z36C48XS6m8Q1WDY3BRY8NB4lXIfhf3vJC/QGgIocCyOH5
tJd1appCV3h9BlFCCaE7iaBSPgA332AoO6JC2vr2IssTXW+gUwgv67VmZapz8cNM
PFHRzdvUctmxLSLg53WCeQohyD1n+1f2KRUFps6z47ij9pXwkD+4QzXHoIj4HMCm
0d7Coh80o39sWBBQphWwfkspj5tniJDt0nblAysR5+MSQPBrk8wc/mDutvK9MAfv
FUmAc99KAL1kNmuEZ9GC2hv+Ty/IC5O9R7pSVWnXKAcBcKs7fTYl3nOHzRR2ncgl
Y7qbjdsx3ndvPVHP4CCiirF5y0oxUYPmJG0pL7kchyhwg+Dn3mSzNZqf5y/aRp2Y
Z1xK7+T/pRutgMeZ5ZgC12eJIBBSrvJ14BIazo6X7DinwScmgobql+v28dJvq1bE
LnpwKR2fDeEZw1WnAehw5gnE1AQ3B9sgRmeEr4NFKYEELrCpy3Tq8OHGS3WS1g/O
OZj/ZJNxaVnHYIqjCa6jEIpo1vZGkHtfUSAG0asr+9kOEPqs4ih62OwVkykceILE
Y0xbVfxTT4VizXD8KDiYXYsw6aXXy2K5gZCn/SMro1/3dJuBSlQdyzSjMtniosKK
R65EvTXbxKrlMjRfrveDM5ZWwNoqxX3TZdkB6zSD62XrCbYXFoNTOSJ1VrxuRtT2
0Rpmuj8OKjrduuOwQbNO9NO/b4CpU+KmHhZ5UMzzBeAopXAOTYBuL75t+TGrjVQv
F0SLIYSffKlteSUcUsYWGqlBe0OV3kdpoocxbm/r1/SLScY6bXh8OfEmJc7sh2rr
2LgqHv7/GPmvdLQvieoimog4GAPJyLTFzS208eJNf5pT+2WPFbpGJfHYlIvYXMiV
bWiHcPHTY8it+RGgGwt/ia8R9RsqXoqxTMj+jllJ+xDfnyZ3RKTN/IaO8LUDOlTU
J8HBcGb/prLwL+UfSQj6pc7q83p2hUj10J/MvS5AWBgb/2PmGOGIeIgRiiBKX9rI
IXBOMzcy0Gcpm0GQ++EM/pvXPUqOcyI6yZvw28NYpNHV6UKGIXYAINMS76W8PA89
H7Uu+n65sKa1tB7YPXS57hH6PzJ2H2fzrSGKuYPVSwbfOgsIp57Qe7y7qwEr7UzV
9rPUVHPYpXs3M+5pF9Ks2EB/+c0WYYL7D01KABfnsBzzPY0THhqfHjP6DY3IGWI5
rnM6IkWjBoBTtJ+BQfRdvz7fYAVAeI6gmSH9h7iWwNhit98hNbJCD5VxXsKu7OFX
UliGCO0Lk/gdMBcYRXmR4qSkttc7bysqt8L/j3k48dbj7XG7cidFH9mjpXrNPkVt
OJyJhncu1WKnWtJsrnATP7WnnFZCewiR7TdWo4pjkqq1FDTTUxiWtlNo1G5EC8hy
CAPBNZDw2Yyv6WDjHe5jUtfrHL3/IBzyK4x/9Ggkl1q7Rko3ob9UXiWcGxdAat9w
ulWI8eGTaZg8U7rXmo0OpT6ul/xjNvryOslRvQo8jJnP3y2pZ+tQR08UxVeS1+hu
L447e8vpLcsc0XgFIVuqpTR+fsXj88FATTclY6tgnNZR93zeCxcCgCofBrJCKQL5
RHM/XdGGzCMIbUCF3kGG1nVqG/qEEgyJTmxKaF2jR/O+GFhsP5NjHSrBA5X8z9px
8gvRZfpPSbb9oR3WTwCNH5IPbvGKsI08loSv0BefkfkP6ADJTpGFRr3JKtioaNMr
y7HKmnKiatNrWI8QYf4sSHE1aHyd7m9QcHbg3ZeGurv4LUO8AikzZCvLwC35xdKe
4nwIMk//sevR4G8JBWW8qqr6BBriAFHVWctRkpVlqxYIL6r63Lwj1bSgeXutbE0V
OBzNJbi+8dvmifpkBTeAr0TLkocL+VftPpHAVAHslujhgV9RPAxuokRif58VdsQb
uPgfVz/DLCQ7JIK2lH6QM4gMuXkcrRObWCJREX+1ZnWgBfHphGmoVIXbO0doDsWX
jUGUL6q8VkPQ2ldDE3HX6J+Tf8+aEHwsyp7SmPfJkwC10MqCPTttVQtPpdxMzdzF
8uCPyO3/KNXleWFWrFlbmx2VtvS26QdJZ825CHqRPkqpz0CYzDl6/RwjFM4/LAh1
J2vOwPg9BEat7WrTOyLO5rHvR9XaScljWf+75pr9DfJSRoPYD2lgw+v3R7l7wzVW
L7k4zh7C32bEafrwLTysf/IrpFOT7NIPwjjO08BTReIXceyjWWPgSpWyDPwCUi3i
+Q5/WIGjgFkYcC+yxZ9ObHDlxJa6p/owLb+BxMiZA0oFpzzbFsH0RdgxgFmmbwrB
fncFSVbBz4CsHmS8GZ5rbsBjrAel+jKYTmRpa00UBmM0lnCEa8vayWDdi99YjTxc
Bdmg0x54llndpxhj46iGi3qyBj/mqImDnGDsUe3CnUuI2T2vEyNtaDHbBIv8Kogp
SOWxm0CcfBh0o5QbgyezTawuCvdwr2Nemr//BelRVr8ENl6yXF1ZkuWZj/YT8Ils
sCZ3ia9pPqDza3zcSQQD54FKK+xwMdtAUJ8lqPZbv2hfxI+bGbst/uh4DAQcKldH
67IhVZO/sY3i0rOMVFbt36pKfGVZeHHXqjiKf7JNWdf1Lcg8MTHvtpAqxx3K8893
BVdq0v1K9YVs9gvF70YGGrpYf0FXDNEuqvl+dufAwf5YYDzyoCQw2i1/+2sE0n7+
YxBFJBVleM1QHWx9P42JoL2M2S7tAzLb1d7oBXRCaUNUJI5HUAWpb1Bu9kreuptL
UtUtYDpN6+AGaGWR0HfL1SXPDaqBzuqC4Wg5DmwzUEUlhg0E/Ew74ET+80VpQ4sF
Yn4e7t6ZlQuU14aoWBpSXcShVC4VMr615Qnd8NUmqAIU3qmg2Q/MggMkVJzRLy4l
aeoBiI/GuGzh8l1VIBbT4kBxyG/FFJRoqq1R9cTtOxW/rwpUMhfapoNi3N8C46ZQ
ty/i09O7lR4lDKn8uUyWWSglP/IDcgPRyVBZqgTPIpoXZmVmzRFF0VsBJPmuEj9+
6izE67v8zKHOiOBbAI/EkkIS1tRCE87xyYKPWd+xCVyuWEGR4aV/L5azwJEsjD2u
hJevUzTiGxidzK7IkPaITVc2H6QkR37lq6sbMBdhMbd5l0e0Fmtcs2Ry2hpf/VOf
ibqi9vzT5Mpvxm2taijrME3kmrkkQLRg2yoggIqw/FxpCCCyif12rAcfXRWOjiaY
2lJ+iRzw7v2iwEdi13VNBahjuc4zoCfBq2RIMHR58SKrqZgElXf7MZgERKaGve3l
KLY78rCxFN2uN8JsWlZK5ZRNJfqOPKU26aJ6xZbvqSOF8dKfR3AckMrT8SRC1h8z
zvH+yscs+XYKZAvE8J8EggxtfgjX54vle+qR7d0LF71ed6ktrPUF34kphowjJnbp
dO/ROyjcCLa1Zir/iNsooMyakPixx6bo6t7De667me2VyERo/htw+r0UnSfGlQla
qwUXofRBVLWDboXAYINFgfDFUROQUTTCkPl2Eps/tGb+zpngKT8wijad+3Hm70E5
kmkulWOeZoZI2njMU3p9iz5RW1D68Ta8sFihhy89ddBM/4+JbaTx4/5SrMUK+nVV
7ct6QIKQTl+aD+2CME5jDnZpGWw9tynuzVogHi44UH4jjnN7iV3CVd+Li2NFIk4f
3CQoDXfSV3IHJ1UDz8kABl5SdP5jwdmgZ54bWruqcI9ClhhEKo/BA5RxdCpBo+I3
AWKmQnFqrwsQ45MHxQjQZCg8lrT51WdAjMhlnYF3Ozg5+t3tW0y4DBM2dCO02pEt
JNMaPfKMeGIVwhs9+QvmEqUXJ2+XQji1Sr+K0z322AYod4BtqacXl96yjx9lLnH2
LJuqBuAuvGKvrKBzUNJ8e76r7IaHjamjsz1JpYXOPVQF7I+wZ94qIxOfkrfj8fWz
6xkXtepPFl+oVFYKbWsZGRexEZfe9J9e6vp0E8rxzwzc2HpyNsBiaCz4E+F+BHO6
W0Ukf3dZeNxxSsMxJJVsYOMDPbVF44pNXav2l0ur8wspPWYFXifLCna0mgTvZQyz
Cm+VPuFWKDe5CWtzmYFqHhlPLwOadn9qTvHCnABV4lDSss2rkVBu6ptmOUt3GfNz
JUzAtgCgQWf3fOmMnqKsgB0+ekvg4fguGzUwU80/Oh2mGWz+G50q3P0OwPvrJJrQ
oGp044B8vTqGc2NVLAXFKXeof5gMz07mhKMkopqmLEEd3buJE0rH1/hIzZ3tpPDj
uvDhrkQ0E44hgG9Wk7FVGd/0WBbU0v3wkesiedGre9/LcjT/v4oncJo74ENGmwWL
/NThl5d9+wL4ZvTsXiTYhkYmDLP20JuFTw2nOq3jl8+xGsGbXJPgj/c4wxi6b0Uj
Say10gk3b948YTEdbvLcvF++xRKkhjOyS6FpomlagxvpLBPWPYT8nwPZcRdVpGwm
FpxLAdM5djaaNXS9hlxEfGFkrKoKopedviiaPlCM1dQk2ITLwn7NFkbgsPMHqYOk
RHhV4jEZ/sNmPTSdw4CdH21Nelw1Fj+/d8BTcWeeP9e7rEwOafVNVPdDct+Mi8TX
0+V5NQ5MSC1sADviB/6VEgmJMOSc7Jo29NZLyedzjLN/Vi7AisBTtIGGWWay4wjI
9ukAkBtwM755wyGyMs8itYn9j5cnwh1wWK/26+Iqq7sGE/7XDX9KWGEA8UGHHBCB
VDO7LeUW+ifL+XtTBE3IuzzBZB5eUv9nKwcdntoZxpGDL9D4/+CR9rVRoDJljV3N
2/8rINZSsyH+Q31Q77G6UVdFIDlXXzmLHOz3e0B76donsH3BaLf1atzAj7XZGIXN
qLDinM8BCf1vToqKS7pu545o6WoAxBKYtLz4fAJR8xtZJ4MsBx9OAdhjR3lMEpwC
qKay8w4cmTs8ajmnbjvi2iMFktQ0ji4XiY46iQjkPT8TFXUlfRVYfoZcDytr3dMn
xo6iVJxvIvKdmhd+kQpN1S3gpc3P7hJcqvJFMoRCT3QhZorPqD5FfbtndI6dVDb/
ErsbubSAMgacLUmtiAqT82TiKglojIp3kLIoynI0jqQmOtvznIfP/yDTgxJR9iBX
8VJj7q1HqlVAcF+f6g6yEfEUDm45V/6m0Y3d1cCpRX/MTOPvl9/SbMSvFeOsW3o5
XQhH9Sq+fUPgi51pWyY2YGCW2XDhKPDM/Aizq3qluhjrurMFWuQRYFpgTJ3UgB1F
dWCaJmGWE398Rc7iSihwxVtwAf3XpqVoGSAELFvli9OSyJ80A7cBW3jqz7TRVFGB
oroOIlU7P3TjpbDAV5GREUwhnXFyaYR39Vtz785ysW/U12E6WZKgpTi9MQ+cMj5m
eR13YSX0rM9fQj9Thpyidj78sc28aviKYTmsaiWakeXXgC6YGmeRSoosjKx2I98p
D9bekqQFEy7uTRF+KvZ0ttqTqZ1w8rmu5ESB27RulJy0vbhuJ+dQXnAVjgoGnXX1
jgvcIYkFVn7gQ7FBvJV1gi7E/AHCY7jz7cpJZNuNYSot3oaMDqTMl84p9BtCJ79j
iwte8X8wEesT2yiXqVMlF2bmxuTfKnfBRRsCkmpbDGh45Lyna32SmD5Mg1wsnHeE
sNHe5o1NMroBJiDYmmHfgJyJN/X6Q8S9rvrYjREKRT4HOMpwBOmmMN5qpzm6DMb2
ni3FvsWCE3O4KExgNZHtrbG9BEQApgURsiniqDtlsjFwJbzE3E3wAXwouS61OIap
+leLcBFijhGDuw4mUFSItuS/1EjJQgH6bdXUGI/Bd5A8OksGW3YZFPyeSNm8jQ3p
ngjMjW9pzNPY69XW5oCQqj0i+FSWJKWTTUygAJMBO1hZnxrq1agfrnhJ2s6UQlIZ
cn+GZrC7J1BMQMzO0R0HX745xwF9KgNUgLLnWszMc53jGXcz50jUMB6F1O4Pcygv
rdYPFRhkePLi1HHwYhfhZ/U0emoOdNxotRHW+yXj2OfQgNB1uPYJ6TQXbjVPF3Le
oyDiZjDVJ9lxqDSjzM/u7S337R+qfoNw0ANGzs1d8uwI9PEFVa08QH4/bY8xDQWv
BSXntlkipgamUuas1wiCMYpVq3a7QUeT8H68SXAIiIY31Toe6f/D2qz/yU4zMfY3
nIR1wgD2VrDomsbFkSoMfLOcofzg8TjzXZcMes8IpQoq6+RsSXevBnToMAO2bQyf
hDoAPiCL0jI7oYQqF9VncDG1hQyQhhN9rac4RrGGBq7ojGqZf9OXnt7Klv+Yljwy
1F/7+UFgHNS0pERBThOS3omp8tRtaw9PrKuCgt86XXwGIW06b8J87CUIFbOVSa6V
hRcy5A6n9J6YdlN9lqGPo2kmSjx9+YQA9M2KSp4Xg/3d9rM5mUiucQCZLt61x29k
Opevdel4Ira44KpTmApVvY6gcbqUSbQh3JmGuYQXe4l3MioyfIrZ7ejOZDRHny/S
iGtryAqV97Pv1ghAd9ELnY6bMXnzamgU3DEQaKe/jocggWiEAFP1Z0pEcRjvKm9l
CNN3QYj2BJ1dOs4+ah9y+nfAjtLZxBzsfr548t6ndMmQxXLw0jwXMMocDURqsmIX
YD3GDUdPNjZe1N1NUjNEwbOlOmcm4RHm3UOwfQjvESdHzMYsHrqiJM8Zie+gMCY3
pJG43SBgoj7778OkL+3FVT0pbT+bnbypNOj2IITdQ4MKU/zMOV1RIvRWQYUosuTV
nIS5pdeljA4PN5n9Z20MWqPq314tvE2qaiZXs+vzoDI3OZ6EoBY1gvSr6B34N0b4
6sS9E1RX+kX/pSiInaOJF4FzdnO9t2ZGSdzK0ZLSr7s5kYlah/dM0qwUH7EGdAoH
u5VP0rZplNuJE54rDRgo+QbOoKo4nru31/ebKvFOU8Zoq20QTYyiYDthrQ29BfY1
dnJuAfPIg3ah/NzVAitp/LIGzG7z8/ey4d11PbIrVKiQtReD25ULI0aPx8pHKlKf
glvOYSibuYE3OZmwocfYnvvuQ8b/pI2D1yfiObY32KkOdjRzAfQiLyks3/efzuWS
3//9ynu/HHyxHVAzdTcTJZ18iLSGh/fOyXJFg7DexMN1/vBZ4WV6lWz74hQaia2W
EGH2kZ0k568PZDjqdj0OXc65LkB16ruA266Nq6F1AzhUjCHrnV2Sllo7BmpQ73ym
pjesYRZmbTpqNOXkPvXsy7iXgtLbk7QaAkyfqM3UjaGa6pQg+H132GpK32P4Qdjj
dgnQJP+BDr7V1wO6jMsgYeLM4PYs5Bm3RU0g/Rplm6IwU8a1RbT6chPYsP1TjL45
YvkG5rupDG+Ndfg7K1XNCTNtVgIcG9RM0oLqWYflI8FLc07dKWIFLRCPiOmUcSYF
U+b3se3wPaIgmJHD0rvqehNU+rkGUdLV8NzfJm/A8F14UcyOmhtOWk+XD1ncBQCB
ayEXwMhlQUvA0yVN5OqDG2Dhvko/5Zk9R6355Yn2db9+Uw25iM9xxNpxSlGIpMoh
d1TCVRbUaATrOTtOtJXVtkBT7xLRiDHsYOCfnGUVXrCPVtDD7GPkSjRv1iiNhSwA
k8EsPc5s97bMmTOUa+a6J2CIMHM4tre+9C7OcYGRf5U1tocgKYXKGWci776BnKhc
0A2ui7O7CwBO/B4Dh7OqzckaKQINujl1TOmPkdC0Aq2eqZG4gzlpeHBSlIz8akPz
xW6tXbCx/uEj1cdpxfU6PwXy8oGZbrNZ0fQbs9TMUzDFQYoBHYAxF4lHXjLkVrR9
k6G7sHRnSf9W/TrHx56/pMnZE4xGc3Hk3/tHrUR7WmcUiSLc9ac5+O53ObiQsmqU
JJjacArpQmeEVdQeTnj+5mGtjc0osvmAqSaib6/BJWeGp2cE7cgjotY3gpzknHj1
pp5s5K6AMtgb+vIPP9aqMg35S9IntFozCJ7E1nOuuodHcvcRnR6QHbqMdgpFi9CF
EvWfJtpZpOUOOSEl8F4ef/G39qnzl7G/cAhLqnSk/Rh0qDuDyAAUYkidkFIs7B1o
TnPViRPp6jl67OxaArfYzs4LKx5zSYxKLvP58zB6AsG5K9OJkeqcgy7yws5xTX2w
ydrt4zdgll2R57vsD8In0RnrP76p+POV/xXHp9pmchw52/5iI1LpFzQEYBTHiZmV
3tzd0hxRI9HHnAdl8y6nNxMPXLjUeebFWekybdrUEhBaGcK6uuTAV622uDII9wLK
0mzmobGIWMr3iDsGldWG1quFmwNjbc7ZiRUAsR7mFp5/aFYRWZZIyTaii/VFdN/I
Qxvqw2vqSfSOvX5BK9CwgAsl9dU1/16CpUxaWvdVuPsDRl1reVAhqXPfVsIksXc2
O4KO56qlO7/UjlIbICuy8TH4S3YQZj8frt2JEh+jf4RFhab8SLcyBwrGAJrwCtLh
7FpucoDUA+B8a33jFia+PbX5+ftiOHDr2qFPMWSLxCwoL4A4oUaORa0yclzMw7iH
cN6vjdktbYltRWVNHUQwfqxEE2jSJ2USlPK7AMTGdZKr0CpsYDvt1IaizIDr8P3e
GWlb/TGauIxtZFrQB+HQC5Ben2MYtgE1EAzC5Cn0jX4C+9oSAH0qNLjJrZwTUQuR
fVLjUrRBREul/A4disPJXgUImDmEy2TpCLEqAZt1PbA2lc55N35Ku15OJ6danTIC
FjoRBSa62sQVenQoYrCC718W6I97KOQmD5DYDJskYIjmC9OECJp6YNNceUk4Er9P
+mjAOGJSiJOsWmOC+Lvx79s9G7sYP5JUuBGnfSaiyHDTmbGBVzEbLJRtrGYfrBoC
JdQJNWQpDkavMLmfkoz+GzUJQ8jOwbzF3XEIrJUCdUb+jBWaoCFSgplj40A38zR0
1/dHa9nF35XhbQ0ykrFoJuHCMufcVgpKdYTJOPd0IGJwo0HTFezAgBVgsdyvHN36
a59pU87tY17L6QK0fOvbHBh1dU7EQ4U1eRDLo/knIGVTWpHExdk/Md/t8LAq2FBr
uDLYv2C28bmWrgmrwvjnCMg8rSgoNtot2PQ8l48YKccEkUwHlHt1VWX9ZuwpRUTa
1Y6Swa/9dZSlqClgo3zUC8Z6wj4z2TAMX6UCAlMAseSuNQz2e5pshX8l/RSf/81F
RplAeVUBz22yQp4bnHsbQe08xXHyFG88YHf/sGDLY3vbk7FKm+BuMSucsGuGWExN
aM+KDMAxwvJsfRzvJX7aeR+9hpIcKJfZDYCD6ZBWEzZM37DvE/H9yEwMQfhrgmXN
K+fI5DPyePtJIMLAQeacs7jSGi0UGTb5yETKVgbUStdvvwzODJXyLFQh9XUmykCn
XEZNhET59G01rOvwEng/i/w4EqII1XRUPkImbSU9/twfZFzlAjYkVKYxvgCb8eG+
hm0kBIQC87tQ8BXRqfeH8CHVwIFKx4w0vzW3okPETAu/+DdUFhAu5guZywGtO/J2
j+L2h4ZuJwQHc8XxKaaZEGRM+8rz9srEBTma2FQXHizBqMkzpTID22EH5g/qSZ5h
ZyqtBSp9jm/eLv/hn5HgZfBMPTXiqG20zGnLZYPT5tHhuGQNSlCMXfJoHq0sPlLB
aeJpewpY3eJWsYOHjf/Zln/QWQeTJJ0lLwsDHbWxzAY+oaqXvkTc4uWj/26FYAoD
USuyp3zvl+V55+U7hnvmSNSC9eETMH6L1aKs19EXGZd7+ShiwDJihFuWLBZrsGvr
+rgd39KJCGVdinnfgjzV64vb/qOefcjlv7TpXh9xbFwX/bvh17uplsBnsF90jWaT
mETzgSHpDcH3bCV5fG3Dp0hwyjgg7QXuGQiffqMaMRnWpmqq5F+zWsaDN5QUGmtN
gNrwOU0EZGsntBaFN0HzpQkBfoVaok5ADCZYN6w+TP/PgeB1lAhn2AeUuvgYSgc2
VBLALbg9GDB5NiZbMK6NCArWzHZTHVdzkngOsN4kZspKk7OBcyw7kKuI7Nuws5El
FkwQPUzmMGE57LvUgrX0zGyFl46BZlHeJku89PajpWCs/2Uo67GFx9Ap63xBd5WJ
RuwDB7YNGE0VxYyOpTZpgKx8S+GivNmvqUiqQ2jN1FjoFuJ+1CFLpE+IDOLrkBU5
GF2g/Zb085MiG8ELgOlFkHwxeGUxzOPXNNnoycQ0ZBuW0drZSqVt3McXztsBqn57
CK4Pf1s6oX2D2Q6kkwt9GvELecH8BailB7qS/Z0cLyFw+IHucV/VH+RjGluqah+r
CMrmbDq28gJ3LDApLok8/8evOjcdjL/rhKdNoaX6lbHlKxUAP3081Ei0s/QaGcyr
LhctEhcTLnfaWnGnM7HPX8msFv9QWo1pXf1Wr2lGDYzyRCrCx9LtS/5jU/WJgClE
50GKXR273Hv9UoJ+bzWkA8Mz0XtdqtC3MKjzJ9sorvNCGR2hsbbKj+TD6MUp5UIj
3B4FDknZa/89dMgMul6EPhBnYCFod09/begO1Cxv1ohwPcecS4oosx3Jef20FjYy
WyPE9Ely3SorIiYWelx/9dc1QQ48/yKQDOHpS65v13jrNBI3HwvAspx7oer4OS7j
39x8kzlg8yJ2T6mpnBW/iG+Ltb/rwbAU29YEM7sBzG1pGhA2N86REBmA3+J2VBBP
KSc4150SM9n/p0jm5BIQFLSdJe86E+xc6VfJfTyiqx+nqh+J4aIXQBN6PueJBs8w
rxpWucrSgkJQ8hkdPYr+b+ngkXSOLU6qjhtgJUP0xt2aVhY2EHncMKxiroKVoBXL
0SMrO6j+R4RZYITnqCfFLVDRLA70qEHOzGB2rQy9Z2BBW8wNtqVUlB7v4b/7bJe2
UyOxVK8a3dgcfR25AmZVcRH/8kT1p3Ffc1WNpNeql9kBSFJRNh3ovkGM5jcp+ROd
xwKKY3MLgJLN3qP8NumScVXyQrWGUl2nE5JKuY63Zbo2vqwAFDivUJQp4yNNRgX7
LH+VUHqLGApwXW5GxN56ysOrVZXDIDH0HxXRCkQav+c3gVwOVugwZTLbdkYvwCNP
9l5JyC/NK9f1hRro5yF+TNRRBr4b3/97RZhJTe2pKWPzpUK6taZJA115rLCpeu/o
QQI8MC8dQxnqC4eNgxkj4XVtFDOMRSKpCcASZwWyOxqYvZFtxtr698vUaLxemKHX
uPvfE/ibXHn7/p9ju4HJ45JBbucjuX2DlwHqMZkdkPm+gio1MPhppn+jmxLhIZmw
ExPEKHfEJ334gwCFyXhhlHX69N3BBVZZjDOUkkYL1YtaTBR9CnRqzaAg6n3wJJd1
4CIdznDzY/td9U7RSZGefi4QWVxiv0cIYJzOEzOoG+0rL4kX02ekW69CBAQMPGDZ
N9EYMKhB6l4yF6Ah+NR9byoMY5oskF87s+ZIrq12pSGa5lsuTJ/G/4KzTlnQj9gu
N6nyCt+OXPNR2KPDxv3ehhQ+wbz6mt6XFiFCY07YhWIicqgfr69wtxkveLNsqEPB
fy8VIrXpjc484D3h8gjFuKticMQM45jHkyPgzYO+/GiKGlo+j2pc11Xokv3U3vOR
PuAppo64ldJIB1WsWtAWz95ZW142BeGwRW3LDvsCbSmsa5l4yieYFce9ivf6wkCT
DiyTub6s/8NfDcR/H1HAQedWkesXMSW/Yv83RL32BKKdYYkDURy1QrAtqytfaKay
r6D1LJAvC8SX6DRNHGQetA0bFpM9u3devTtsItexKoPZKW3XgP9KUJycs+/mbyul
k0LqGVe2W8iFy8V4FZYtAiDV+zYBIUeaV/S/9tZWhB2HGwX9ShDadj8lLydbvpfR
CB1Q2aarxVQ8IxQ8Gv0dVmHlYfT3i39jkeN7LeI9BDFSO46FzDHlPtL93WWQLDVp
GxNXepd/GTQESoZxln9kQRqrU3SeF+BRM6hNllpdTs6C/l/VleImfxhE6U3O2YW1
l/+8zzceaoknNQwyoz4AsjHlGcqRhh+B2m2deKg+vbGR+GJ/1qx6AJ1416mDyGvi
JnDfbnD4VT6Q/ByT1jfjHvf0ittM1NdWw+g0nVt7iGh9+zCehp/zopz5kcoUdSeG
EMScr7imTM/SIanZz+fFQfYkbEFIy9bhN0EYRYlTOxGPwsXgPgZq6PejuL0PYbbg
+FQ37rn6N93JZzcvSH8nEbzut9MtYzIJrYI69LmV3mlkMhc7+B70//eKvln6jVRH
OjEJy2uACZjmf5AOPvcVBZ4fIhO8Rg7C8oT8T9mFBNkubxQnI61WAdAbj0gwFjUP
J9RyhoLbEzHfeqE3XGIHSRNxJ5yOC+mtfco1cgceloeQ2s0yUxqUTrjKy+BHbkDS
9rxYsgjpl5ZgVJ8IgDESc/4pWu2VPkQv+CcJC1eUBMFJ6Yq5FB9dj0+137vrOw2N
Z1JXX2QQbXrs4zichy3w78o/lQ7oVVRgblBOVx+k6bZAH07e/7GcQImCSQxrwSEf
nH8HGWVnJ7YrmGUf4Hakc6x/Sk2gC3h4DfxY0h8cyMrqcV+P+3u6l30vCZz2UgKb
NH6FernIhEhXsQcpMbeM4euJc623Dej2xKe2Z6et1yVK/M/z524eO7HIkyHjbTRV
J3bPuB5Q3GZ5gdQJIKoztJ2oMYtjFaCfzlvnLo3AJ8aspyqSdziyMrl8uT9qh8Z2
fT7bquAXXZ9qtV1pjpT5Q1TYtSqpUBUuK01Sf2VIk3O+20qFCisRC3wY/HNREHMT
y+gPRJKNxGqwB5DFbUAhO4hvsOcTHwBRezuYTNHfl3GqwMZezFHoWg1bOjVxAEHW
R2eWNC4eNcr2vSz8JD9nxNSOvyu4XAnLJfS4oeGA5c+lop6qDx02Db8UVOGY/4ax
CDoAe3tsJw97umaDU+oZcuGGPPtmXPMKMak0aC7DoQoIPy+fcetKaeGrp46a0mNW
2KmWtif0Men65KbGh3VLff5keF7OX4iglywk1yIkS+IQ4Gq06LkEnO1rOS17oyVV
AN8Vz4ELiQTd3IRQ3BEb9KEDlZNcV++OfyG+vxzAOcgHZrcQdvecgHbAH+MJlPpN
ngWXU6AkFyj7k935H8cm040mB5LRsq6DzcCQwLF7gjn4oQ8pnTNdlRRtxDIR4zu2
OaByBn6NGfvC4FsoSttNf9aKkgrdHrO+DimN7Womu46UoKBPMfS4tUfqYyPt6Jkw
xoDF/KNFQ5FzFASJggFPu1+kKyjY+cJQGgjS1YugxNmq1iRGALqJQlWNpQqlOxmv
6p/UR9q2ZjUaGCPXVGPsZW+JLIziLxb7dQi5gAOhe6RetJeQVOQHXlp/NqBbmju/
l0wGzPpYdtm0yJ7/CbLBkFISzDeH7a9DWiW4Uid7XHBtO3x9HZBpPVHHIt5PXw4A
JBk6UFKcuPI2q7r+KrvCjegUYSuO15qjhGvs0uCHjfKswrkLcjt0RlQTNYtJgSnx
04zfM67ug1xTaE3/MEy9Xy4qrKWMYMCwfW82fsfmY6jgUA+OUjwkd3N4uYeMdSSd
ncMzxYgSeB8hXrpa3OBS7mGtaeJ8gDLcLPD2ROX8gYT5qy+KGB9mmIxUh+4S3Plm
h9CzxzrCauOKq+GUK6VOZ8cy+U9JoTjbJ0WvEOUv3PlES2amhjH2WhXJrZ2nyuTF
cO4c2R2V2Zz1TCOFFVLGaspuPF6JDpN+O2wiVm+pxrIXrKF77Rkog7N7jy+B12md
FCcVNtJWfEW5KMI29N3mw3snZvanAvK7igg9UzHvQxuxUOzqHpdrTs5n8otmDw5T
txDKIa+Zd/mEe81aeXYQISrYYoTwtMi4GPDyCt1d9qWAND9skep/7j/vjUvPbnl9
J2Z5hFyAu30aWBsHmatYk4A5v41YTBo+98rKsdZ/3GQBMrs0l/cxTOH5VhEVy8/f
sJ4r2JDQtvrXZehuqRoPWM7/VQdZMpViULandOOSiboF9+ueigv0uCkINik1RLR1
ASOoKCV2KKZ+m9mf8dwncWVbrZjHbXQ/+nciM8G3rNRPO1zr23nUYLRuPF3iR1cV
hMnvnvRArCjcGjx1X9m9ljobb0uiazw+VXKAS9q6fR1hCiRFHkjltS5HxOEdVTZD
EM9eMW2oC8elp8X+GcXbzuKqXzgqSPXDb2HqHTnaEDGmHwT//TJMVcMjf7bGxlGk
Yq0n5lxEaPkNj6emn73LrByI+7+NyqexO/i3WkZqB10rO8qfkkYyFMogkkt9GN+w
aSSEdoNosIc7EQ9iQzHBcD08EEZNTQ7qK8wfiFyAySR5ElpDzusZAHiTtJ8PbjIz
du/3zuJxAKacag74ChMJmbWLtDYxdfymt2WJfGZ2+U0uWPGj+DHuS/J63EYmD9wh
pu/ohsULb09jlciMM8GoQZMzpZKT+vyVhkC12OkWU8vSp8SMmP545iOXOEsNs4AI
RPOn6CAopS9+ax8omKKweivXNnOH9zQoxh8BrPjza1MTVmQvnQQM+rMqDPqYF217
Nzh+EV+UsdQJAVyru9nvLG7NV54JH1VNZeN4sgOvNkJqk/68b++PXiV5ojyr5Ynt
1zujIZpjhSDUmtH2nTwmZmfq5i+GgrLZQxGnXtZGbKTEqBBX+dcBGZriiwYP1GG2
RpXtGiQgKPVViJJfSCtPN1pbptzLwT6gPHr0hd3ymIJ7EYPyoj3PfXFd2MhxWX5w
rAEnHWSaI4Hmy/PpPM1Zdlxv9RhUppDty9BfPBtTE2gJpA0IZ3EjmHTdrpO3W6Yy
QeUMIXnXmbvHpTeLrDd+W9DAUDIdid39uTVWQz4xi5R7kBwtJoFp9XlG2eNbItaX
blPwuGjZJKJIQBmoT4Qogu6PUG7+NoszxRvfZrqEdPaEVnOUVQT5gTMPQkL2YI+w
VlKlmN81ynlLGYtM+dah7qtOyl5IYMq+xEhX1RgEqNqhlsOqYzvl+cNbZQsk0GAN
KGO5JnP+3zG4VIbXSv9+jg11AvbLJ03M/YtExIN87wu/J9Pfpo+MV0B3wi5RV7sE
AC2b1rD9Ds/bDa5DxAE3Z7UuXl6O8KJus28Nq4WmPIp+MJoK35l9KkHOGUxngJKU
PmzfKvJdT1/BxDVGY37HPhRvN5SJSNkZQD+p+50x1i03unjDkmisrv1IVSb+s3eK
rDn6f4rw2x+UVXLXxlqtXQskELRPLBg0VKzsc7ofZVIOOZldz3Gxv6AoI7g9BGUs
sbVUOG5k4oGNQIVaTeZRYpkhBq7bEZCIfAIEpUcuKraafeFT3CwiMlAYSrW/W0uA
SHRcz9WW0xCef4NYL0Culiaw4lOGmS0QQrOxk5n8RR0Z3UCxZsC40uKccK8rF6mQ
RInC/Mh789dUPcMHx5G1X3l1yTNYj+NZdYpgXHJk2ISVhxpbWSNLV1MPwzE49VsU
FP4kFdSEHpc+R6FY9UXjstF/wFqUjTDllqE6Q/bqu+1JQPWEeE5zymM4qlKChAPj
MUvpOs7YMT6aRv9GoT4Fe07FgdIoYWoCAoVo1f7ACDTnlI92414H2pYiiGUSNTqN
y6jqyc3gC7cZSM9/Kore9T0V4ExEun2Isqwr9kmJAiXM9dmq4w7aqjwIHvgkPwKc
sk6LdB/GCw+Ps++Ps9c6Vw4L+CdVHPQHLnfB78kijxub48H0Hs0IRreUpRsbx/sy
bnJc+foFC+Ok6gxq0zS5+175Ao5cpn/VYQCNMl8oC3Sp+uspy6Zx7U537a6qqLax
D/nXb8I/tCG16JwnQwe79TWelOdaYaEEaWYjFuJRHWB63OdjEJ88nSU5XkGvALt6
207Zl3C7UroAHIIiR0P6H2moX7GOOTLN8g7rJOr7jPdZDsADMO+1Z+ks2zf+gj1M
Rp2D7OmZKcuyHQFygXia+WAw3pSP2DqspHStj0mQpYBt52un43Yg8NaddfYZ5vnd
cRNce6voyxJnf6TAPxpukI8VABZWOAbJBJJUXRg3/cjv0wu24jsL5H3Et4nNS5BN
JWurtAoP8h+xnx0T7w7wd5KbxdsOZVih9WSkPe4iV3gkt66CwyjeoiiMUeTjAbVm
x2PUXCfyFVZSj2bdbHLOHK6nmYEj/tQP601EdBHC/wt9oHdWh4/YqPVdlt5knJyb
3mDK9xDEQFWtKAwMIswBWsMWyZWzSR8XnWmoYDyR0OOTF8d+okDgo3dTuMH//nK6
MJ6I2Aw7XuRN2ScIs7Lrmics2gdQVwYd5ms3cLUYDvN9mN7x7rspvyqw93bZSRT+
rPdbYUvWQNipqswTuXzhPl47hmZMDRKsfao3dzjyZ+Xi+bEV1rZ/YCCQHueVoMra
ESmc0a0CgKNwzbIH4k0dkLCZpowUCXHlwUxlOUGWC3JZpN5Gn3mCXG0KN+3EjGHA
4x4IXqzbpmSMslVCXo1p9GiLHv/BXcDfdkh/k3TUddzOFeuUsy70JkhootHzfV5F
KYyY5oXzwmu2nWn8AO25Wen51fKsXvyfjqwp1rbGPKhIRwoYxrESF0MNQ2XgsKtp
+hEAp2Rj8MhwLWkK85v7DXd9PPKRsEnJgS/Sy/lHXSva7yGar5urS0rikcT/CaUf
k7Fp1k4I8pdVq6oiEHGrRX1mDKinUXERyFG4u4pFqEPQdMZt7jHA87WQpy3DfZO6
CVFIWGc9vBRhKUH/MW7uwISHu1gptqSN3ZaIrgi076nupTkwQEhjSCl7h+FnNGZp
pnl7/rmy8Hw8rYJNoMNgTxQMOfCxOmdiPQfWrsAB3Uux1GAPfWp/GIosdCrpXMh1
OtR4IlmgoitvLeyCqVwGcrnks90wJwRLiLV71Vv5iBfR4iYK5abiwUO/zlrO05Jv
OAGEEj49enE8XpfUwnP/70EINrm4+x+mI70yvJpFrsAIhtb9kgzcORpKbxNJ5ATL
ylTqbRAz4glmj+jL+iJCciIwuIjJW4N5VdUvv7Cgmh8/jqBj9PZjxsOg+cZCxfKD
9E25geFktX8Qsz9/c5338BW0vUI9dfWob7CLlnRiDit0/K7fnfnOs6HaCGgU2xEJ
doLOj/Rieg6t/8JVbONLaapWlTaHeVhCr1YWKqMs8RoZJoVPr3rm8jdUPDQskTsi
gKGtImoUdR3Mpm7i6jPyE/dozsUPnPNYPpDOWbuJvgCZn8oGppZatnZ5dzko8HYY
8kRa4rF+GbINIarsCROMcNHjcsZTG9+QOXzK/h9Imb+irKS+JBORT9XU7Rqc3B+G
ZF4/UhCFpFpPnSMPS+EO1XMnuJE2ERJrssK1WTkuQxao6/AXxYU6gCpMv/Bk5AA1
c/WxeQ/Fk9AY0G2Oe/+KmL0wbzFpz8fbjdEt5XODnvEIZZMBQ//RfNI984v11fe8
Kbp5GwG64jECWoyieRT+c39chG7jsbPcV1/F5/eFIAc1EfJwIyDuzQtZRwymwyGS
FBpoz3Rh2dlZTtrKtu6AWQUF5X7nBpzkrhyrC7OWwKjrIAZ7+KGpWSZX3HbG3FSe
NgCSCf9Ks4AcOwrTnD2OxaxnKzgC4uVBtv/ZGSilxykh6iEhr2mhhXQJGzb9Gg6E
TotZJWsYUwVqqDrk3Ca/kuheo/L8KPm1mUT1vOD6AOGkxxJmT+gxOxj/1NUi61o5
Llx1qegC0MiL1vA/8huwzXuQkNBUgoHtJzA0ixr0eXUUxhRKe9eqfLbKTkAMmfee
yq3ckrZTS5IWOj1LZp+e3NXPelLTsQTwKiz52T37elFK03LHtlR011Y59+2hfZZP
Mkzy+DKzvf9QVS7Sl4otblhdZxzxmm9eJU+SQXvk+9+ZdYNR7DYbroaAw1+RN+Sy
7C0wccDRPPdddjEspppa/qjS1cYCyC/zaRfdJHk5cpKUaVP8qJEbInjvhCFLNUkB
KLPbD7VmASMGSJtLVl6r/CWVFsoFsSXveRNlqah3jrNxnQzYIzz3mDJN9f021UdY
R5HNY9IIFw6cZiwb2qKrNHK8c8eyNKUMabVZUiPgowrXvUVcSwGmUdof6d5bGq2Q
xhXtvQLGofXZThsruXQQx33IcDSmbPF+JJQB9RgByXqCa4qiGvHUSj26/D7GF3Ou
sd5UeO5XNXd5jKAbAhP0NS0RsLuJj4K4OM3oMw8Zq6nMcvnZ0d+5pHcekkZ8DPIM
4kk3TRXJtVPZcb1a5h/IlaFJMIY43ZsTbHaO72jUBTaVEhsFC8xl9jE8KmDZx66Q
76FajWqpLnzMYL7wzXWLFSvcgS65XffW89eHV/Vl2TIVfsyTSyLc0GIF3ENiWbD+
IRvQAOA8wCBn3tqy78ieLl9e8bJXvfpJQG+CeNemD6yeVg/TcaPk5ptP12BZTJWu
YuyZCSFoAAp9ag4pzveTRUImJXWWOlz/VIHPNI5pCH40vdNjtWP/ZMwmAkfVIoAW
lm8tMUhDFKbX6NqRKMsKp3ly54FxM0GXUJD+b+l6O2UmbRlJWdFh/Hv2t+Z+jXpr
K0S0puYq9us1iJ1XqCRKH7QKnx8ha5VEGsVTpnh17iRlY3lul97JhkYFtXtqS2RD
h9PDcpkj9sJjoMLMScr6aJsmElYc0O/bdWO/GkpZDc5LQzH01s7YCKJQ6cu6/MBS
mTOW7GCBWzNv1uIhGhYDNkoaAX+xLyUQdLmjxK0lFKAxosI3n0rfz8iJRlZ50ssn
YOiMpw1zuhJNyGX9lJBmRoZblmmvkAopj6GynOhFOLsYFBpATpgLmwRv6v5ksK4e
fV++0f4+m7O5UU3+S7hze7jkO4JQl+x+JBE71baDjv1EnZw3FGKOZmGycGlevyZI
pNpMlCmK2InY0TMoJdFMyfBhwCx3qJ+8yhVNHv2WezzTYeJGFk1rRGJiwvv0FaWJ
jo+XLss4BmGmzSOz7e4k16LfnsJUMruVHNtDx09CQq9VFjaKBV7KlD7Txf3sxlsq
jfpMGthcphvYe31HhP6DCirdfFEWOepUC/AWM3QLv8FCcHsqTWYcVgXR0UV+vSoy
KhyQpMMlcYytU1JQlIYOc2UOjbuk+9+c66GjVn/M+YRfoZoQW6e5TlfU2WrP0TBV
M12qlWLtoL1vz9Fcdslaq0rV0LoybMgh32h8DshkQgvQX6RzHwUfhbibq9mJ5f+7
wyo27Uf2kjz1s+/Nbq3j1MbExCTJhgEQKb/gTQqpJCYd8Q86WvR61kP6gkzMB4mR
4Hhdt2q6FOx6n2oAhIctZrUsi5zXX3HgGYlX4Lq6RkanuHssd417gumGga88oO4l
p/fYL8q7ihvillgxozNfQGBhbtcwc+ZmrDnuxMsNx1S6dmD/sN0P//rFy8cox0fe
1rixSSRbYW0arzfD22PkDdL12LXWPsMLjCBvRdIJyRUidWhb+x8caD7gOfG6TpTQ
zQjAeQH7tHFgLeaB5eCjiHSzbKCxka8Qe8m5BJXPvFh5AIDzPZcNwsvXEGfhDba5
CTMSE0FsHTAhiGmriWxUftqAp2+Nl6fJZ7PNKv7kiH9YDs87qqNMTLF5xyOZHrLO
g0hgsUEeoiksm2O4SkYICUaYPpN1nURZe7HTRvERcGUuqw1QLmxmOEH06o2Mk9BN
byvsmD8rwn20wHM3JZTDf/+/h5ntcpWmP/kwojz3cCkmqU+7Tp3mwngH6Rn8xhUu
gV9SSIS8chfHlrcBH/5JmGXtf481FsBzGPGqVEwTePxByGfF0IRIwplrssiI4aWF
LWCXHolypS6HwjVLOotB3UrnhD+EZkndOlsaW+f6/hyuxqPspditM9RBR2oWYUv1
Yyaa9cdgSQ++21NU5aWeF3vPLppI6x6K6kACaNWk5IHZs2lZ0Kh/S3G6xuaxPEGs
rKZDC0f9tlqDkaNAWdJ4m7UvhhxgjJd+fVJsCLNHL+SMt9a7u4KG6qAYhvS3G9E1
p5+9Hlft9UAElYxQSfpKlsyry3z88aCO2+fxxpz/PD7f2vMgr6JGF6lBImtCci04
wx3TyAi/t8kWqTOmYHX1RR9LsxHeWrOMlrkUnf88eYiGqZ84LqRRw6/Fw2W1fPQW
d6NuPxTFVN/0yB4R+gg85ATDbwGG5kqvkNB2YmFl1ITgvhe2vx7b4eieJtwq/zx/
PUXLTbgPIbG5u9JmIvFxXf+IIexB7ZZs7VThoWs2sFdgkjA5aL8wxp+1nl3mkGzV
9vXaAmp5jzmmWUEm++/QX/WVIzR4hso14zgZrTx77ECX9F/pwl0DTIs2QJg9IzD1
xTzMGbgemjjgwxOHvxkWNFfotkBOxPyHfjbF+F/ahk68zOD83fxGrszq59Gs9gQr
/RTGnxxP1OaSpnOgbWQIUGWEBO1pe1bNTNUN8p3jV3o9z997c51iTswNRIx1oF0W
kfF4ruSFZ8ZjjgeNhqFsP3RXy2G/c35AdB6A5bYV98oDrMQjF1AAfkreZtIILQZC
kuo9wHJ3ZlJpGdv3uM40IMjeSwNCxVa5WLw/1QbDnXW7HunCQi75CTnaVEairDSU
7AHEBFxh7jU/Wk0WB4t1VcRtwwHwUqsvzX83CsGC6TfKxVkZgxP9Jptt9k69THjJ
dcHQJteNpcHy/Qi0/6OvgZLfK7n0U3ruAanENV2asUXrn0VO5e1GB6yATm3v8gTU
nyihFY8k/J3DaH0bFJ3D4aH0cVeg33EetA9bA34420OPsrMHbia+qoIHTXJ7xDuf
kWUe28tIzKmKdE4yz3m6ft984OExA8H/2feIDq23NLiRbR7apdbw4krbZoCQWZcE
H6D5Cw2ngZdyCEzM2E3GUo95AxmrvHWAV6Q1+Wwa/Btw2H/n2g7tgAF9sci45VkD
pwUWeqRzva86czfwtm/XxiKXANa0XujZ1pPiOvAVhP0O/UHMZySNDnGSp0Z9k5VS
1BKFups45yV2P2TMBVScugHSFOWUtDgv2y26p0xrmuOLYKD/d4FwQBQKlGVt7Fas
wLJdTs0HSUWQh5Hw1BMJEFJPGAdL3cXZKCaUAZ5NnqZN3q8rGq3WWU2VKlAiwus8
9DqxO4PHReUacMbFpOMIGKp0mBjcWHwzrVKrXthVeV/3J9wei7b8TmCIQnABuUgJ
l2aQ112dpIzbbcyQu3CN1NIJX0ZF4PSF+LgkR2flNgsyqO1DQFqrDez00RIZhqYI
DjbegZ9bBtZk3n57hCd5RqU7jTKRj7Ba6Rrzk/3dcHSlwy90US9T4ylC7Sw8f3F2
7loLWRth9kCYGSL26nP1Ksa7ehgIVjqwpJaBh7nhYGK8CBU/mzrF3gdKCdtUgRk4
QwL8PnNZlZE/zHqIzn+ci8p/YVC5lE0SHnginQsOOLMH54B8C/8GMXndpPmawTCs
5YZ6obtrD8opOXDngOs5tAn0nb7weqdnlICSyHh4lODkxt34MbNIITOrBWQ+9Y5w
J22zgSrLY2c2tg3bLDIQ3ub2XJzaY3/1oRn/OAzSy+ktyB1gBpKVwgXyLS+nsHzt
EuWke8jIjI75wm5XJbAfeXq2SGmTJo7/VthtgHuPG3R7am/+XrRBt/vr+dJ3FLq3
ldoWXxoSOCcXC2tcOM25vQLgO2ThCumVVy2P5FFH1NPTCEQSI1kpSrXTmuxbeX0r
0nE7ChTNOmAqNZwnIH8DGC+XTF8gHf2BhQ/V4WfIF3n8+EmF59wsn/d36PHtjbfl
8R+kc39p9TVWswmnNkCXoe4coYeBE4mKqzMG57lZC5nUs30Vp0rRw4Tj+tbO5IqT
t6jXFkpW8qAqbzpkiNJrJLClD80uXKW4zRwGvAdJztzuMxzR5RrpBQg7R5n/W/Nf
4xgpIrXr1DorDCRPpn3lEZ593bgk0zNwVH8EWoU21lhGjQK8+YfrbfhZMU6eR9hy
6xrOYBgVBWlag4xwuhGTzjjl7jQRHOgNHNqK5Yn03+QsxojX/4OQomBCwI9yYN8P
k34oNr+aN30DCrgNpfKo2ORhfGndMl5WBHB6g7L8BnQUyr8/tpHNOfARBxd2hT2b
vCOPceuGdZxxizbsUhFJ2idDWTtakzUK5T7PctbT5SnrQQluYoqmGp2Esy9XoTbv
hdXENJKAxUbuzHWXLH1tO+IVRmKSbbh2fJgIY7PWQO+8QWetW9DJYmNUsqTH4fRi
TEJumpGd16s3yzbNzw/wxTQ/cm7SSTxdW1U67Hof5b6IWj77t5yFVpDWKx3k5rLR
gPjiyTTORB+CTNyMygy+kUagYNQsPmUXGkx3mVPjX3WzDAaaSpRDPFfrKvnccp6R
8f846ydQ48cQxYlk1L7VaMPqZwsnBcjY/mvKfoF4Ujy2fq2xQY5DSrUz/WZJJ2mL
jbhf6PZOm9zvUw037c2Jb7QpnHIFnVfrEDymgCk6wUbnd2CRMxeFzTxleWUV06ud
9WE6G//ZqGCyPG3IxhYbL8pyYEqnSSco6VNxH3qz7PjwSYRwsQAPjt7tWqKFBP+L
Fxgndh0n4BXYYG2OldcvnVkGcDj1ONFnupu7lD8hChPnv1oDIdXknpF+DOgnoN8X
9ZKQOKJ5odvC3NdN1kTVjGLwhxcsX8sAnr6dAvY3nVmmTNLG0IaO9FupZdQaLuW9
vRAaTlmBjN6w4zAK0iOE4frknDAg7+Gy0laSiefDWAOlq5axPY6HBXuyF4qx42yw
1+k2ohUu3q98cOm4i4YrDxurrfR4e9bJI4wLXm7GcXY5sWDIumUOqmSVH0dnmj9d
m2tHy3FardvCy5v5YAFbYcAzcqHB6EyKAKhzc26di7iocejpCoh1gpQ78PzVU33h
12nihGbPDqELmKuD2Ze5jzIAoDXZ2V/z2tVP5uNljjFIWRbG49y6e5vIbXKrDh5h
bY9mbCpATgPQAXtfM94KpoWP7Ibr6b89sMJXsnmHMOcVMkF8J3wuqjzKQbY2qNhf
nufKUELBYG4pqjSmdGuYnPdNDObusBojGeTVEP9QKIGCAdMDagbt6BlACjrssMcR
Cth3SWIwJxld9/mJrwWMJi9CJSnwDeoxs1BkWlHh72Cd7ntAqGWqrlsXtFRYUVKN
5SeOm2xSGyjEtKUqDjb8DxW3eRhCnsdY/9stqAYDcxDS6ssMbDaz98WjhukdU8rD
kje+zwfvJkHdP3hb3c6A4pKZoOUlWnwhcirDKz+xPQZVKurHQH277rpzAoLo2zab
j5XgKwCuf0h2bx7adqmrYfn6LZXINHTt3mddR7u8WninFhujMOxjEf4ud8NfyfFF
SrNKqvgPhOvfVQzS3xHBO5x5lh86zWg328sZd+6GkhpXxEhoCDW4J5qBvDzIheBR
11tgVQy5xi3/iuPgWchE6H8AeXH35Q3MyxWUaO6uJh50yJvPJF9Dy+cIp9imy6Gk
ruFzcIyROzfXddTQSUXVX9whmSxpttjOk46b60ljpy8oEfPaPzQmfEQ1Fcuf8389
Q5o/1VHkwHu8l+en5+pEUgNIhQ51Jgz89LhPv99EJ56K3hslbBddZW+biolrNTvU
q5qZD5xkm2yISD4a2ZCgSWMNBYYvCDHBRa3poq4Y/FCJCFUo8WkmD0cZ3V+T7PP9
d7rq5HVSAfGNxq+FaucXdHRfFuZ6o+m8ec/ie073FGKpsMEO4CPYd9PcpvrAuoHJ
H1btsElHlsJ9OhwaJm4gxle1L2nJSm0RACo4fg0kW3kUA9lWXFfcAtV+2/ob/gRW
5l3uTCr7Gz1Lh6+p+dnqOGoxqb9SVJ/HF2IOo5QqFaIG31JFJrabdskUnm9inAyU
NGXaAGPITxcWQq9kysFFdWtk0JHH8biat4nKV7bVRbuQncoNmyBFZ32XldpiWNSX
gEVuI0rxGIBphn+bRNDS5uVKtgFYsZgsoJjKutU6N/100UnNGCnj60QkPNDd7CTK
PRRc6ZGID9Fs+dsU5idwyX002bwKhCXKrI2j+1lvVXSnKiV7eZ87gSHOPe5/sv1X
AUdQJyeA8rGm3z/FIsk1ACOfhelOc7vxjc9FzMq7/EddZTIUEKfBsYB317tAUkK9
/Ct4rOVjSLjInSHGhSIcka7L1I3jA9RIYeZ1ZSkST2b5Wr3YqRNEon4ZncBShUAK
XqDISqOCARYjacidL8T9UXnQ8dkDmVZFGXGZc/JOK5F/kPKjdvr+vn5AaySLyTyQ
HUhOhQh9qZknde+unmAiMHXxDn/688UNMRbQ+zZxksiW0VNkAEqUa5T/Qn36WUrD
mn6SzkpwbeItjcXj0P6i+GpdF/1hKKWVVQq02bkcqmxuj6B85QdvuiYG747IDIaa
wwLO8MMvVzAcEFUTc/7erkUwPgkjQ34lr0s/Q8j4qpjDmP4V3+v4EcM9p0sOcVNn
8Kt8Rg3CUJxyHDWCNQ+5KIe1BUFSHnks+eHi70I8+Hft12vHcXj/Xleiu/69HEXC
0/cITBntXAXK39tKcD19Y2vrqhHpr5dRgrPN+rK0Nfbc75l4NjM2M4FRSYHTBQPk
UwS4IA5OE044zbTvl4v4vwQtKHsrKvrqX5IHJJ43wmS6+Ngl54X11tpSk8Wjbbss
D64f75a7yz4ulemPkSEeovi0Cm62djgzn2bBzN98AyA0vNUYuc7mYK6sLuyXL4Ry
LuBnMccZHGb2EKIOgfDd680VjxC4Y5CQCgxj8ZKnj2d7FRnETWuXiZzgy8P5n1AK
ZWGX/A58jC6xXIDlZ/mqfTRId5+3/6tcFdbYkB7CXzr9D8pRxiF4CGswI/7oKfDz
SdCdkdlyTqT5v30CZWJn7CAs/t766kGJSnmxZ5MHghYLeWPxTNpeZWoEUWuNwkLp
G6PPdJwMiP62XGL69ZedEWZBRM7ezYWDbIde/yW44N6TFOJ4hMZZHatQid2xJjer
WY9XJ7d6xK0t4tEcRJEV0hdvxOJh+L28w/ck2S5+2HALuHsuV8/Y6F4BWKa96FnG
J4ISrBRclsuEYmCnKqS3gHoO89mG6AGfNW8m5z/Daa7ZkucbkmzqgsdEA68KFS2R
QudvO0Q+TtGeQ4uiK3aBJLvKq3THwRLZBoRKOl6HCfC0om3dt5ldqhvHwV/Rfoha
lvlVgASOiw2lGKUjUOtoW5Ue6ZVS833qUz+tiTYg1/xRJn6YJ6AqCQ2LUQM4OiUp
NcS37Gsa1mLIB85GxNjchyUlk6R1CBmPPMHvUdtpVx5pIOzPisLOL46Qc+SXe8sa
OhE2W1qsG2zou6njhcIQht/MlDNXKgBUXh7Gb84DOY/1KUzUeC5o9S5xJ2zqwLdH
pwyIfHNGcuB4vusvv58QcU47lBxfGC83t4Ii/BcygetZsPvo81g1fNjsXYCVKZ7O
ZtbTMRQFMHm1z02ZZupMQdCv90dMVhZqASKafVGAq0eH2/ZTD4V/bxYn+VRf0Uw5
RUIs6g5SWfaSYrsNTZHPXzAI7Uw7dOHrPhZHE7xaAxftZ6IG5okAIjdlIvrdP51q
giiMnjnv2o5XLLwoA4qFcDcBfbUHOsOW1NZm6w3GF/bBCgsNO4ncT8PaXYlhFMYi
EPzCKdgrydwY9+n8SMDXblQjBYMpY6Eeg3VJgelKJKdN41JCXtZxZvQZeFlm+l0z
sPCCWoKNxAxVYtiyaXfdYoa5R3eKPGdYVXxbZLZYMwVhuNIm8FX6Hn6ISD4eUnXe
Zj2o1JGiRuvPSyuIAjEJEYhVwpK6sHJjU7tmpgQ6GjA5AAbGsG00o3nLbH2jF1Hu
H4rSUwc2ps0yjz2vAFLBJzjQgVW0vf16NvrRvTjEFaFE3HGt7/nnt+SC+loOt1X1
Yf0pd+2q/MqFJ0Pr+FyBo0R7RCpbh+wFl2ZM593awL/vupkPb36QmvUWb9QfxD1D
ahm7MQYSAoFK6mcgquQmQKZfClSAsnIguIcuyVVns8IO4M79TMM+g/n/QG5ybEAW
PD7VAbwoDVUNMjH4qGvrLDjVoZG4+ckENWDwtVGjGuWPaAFbmK4LOCGbK9C/j3JE
sxJwi0BX/yL4bnD6ET8l5tzVQb6YwDucLyR0X+oneZD+ZRFIFLPmdVM5OtL7hYYg
ZN7bNsqAuk23I8aRuao+GiIlc3sO0QzjYCC2iNbfKl8J5HCKqqJnlI+bG6hpJrjO
VUIbld5g5TmabNYX/lK4jZ+1IpbYjvtfwlgMRuiVp9xYjeG4UnkyXNfOoQw+SI8u
m8sDl4tlfdGPU23PZTqNB7oP2IYzX7XUcGQFwG0YMHEaoRgFcTzsHk17nI1/XiLO
9WL6d9l7sETzRF1YCiUGVar4cqZbq44HZvq7rkc6TF4fYkKd/8OE54EZTUe85ckA
L+ZsBX61TN+vHpI5eU7phrSPmGPhtBPbHHbztGsVHIOL7/EkyTFSvXuF1nYM/yvm
+kgFYdPCa0OA2LnOdqnYYdxrMRxECQQerLwksKNAW9hNQPsjGWQ0HkMo06JT0v1f
E+Qhajd749VW0L6K6QHvqakJ02p7XBhgmP6X0EBgnyuqljHjaPsYrB+EOCOPe3wc
Q427FCV9idEeQECWQbnbGkV300AxG0dW1gUA4lWjJkfjy5VerjgoWT5yisOrVr2+
2EoGq9B3s9MZgEOqAMESB1I1lI06xWxqfThIRD4MBWNiWTJXFLNuxL7hE6Vd9yP+
IaOWWTNPeDEfjSNL6u3rfB05fzjchi3oSj8Vy1s88xUVJsVNDxk01aTzFu16C6Wi
Ifuw3X+r5MXsCJwVChpDjluZGiEr+xz+R1q/bpS5ygcunkQ8f0ACH3kqqRMfMPOz
mvMpBZLdMlOWUAiyXhgyZi4FZ5NbkDCTu4JtYkcs0bVhNyyIV6A4Obse9hTA1c1g
ZaCBhYCayfwvw1TQrezZiZoxK2pu0fp1fOw/AWbrNMGLov6dv2YJErZ34zVk+qTU
lxtF4qMUrBTuG+eiiaBisGqlRdVo6DXE01puE+bU53ezytseH+5jtldLZRQDWkaS
vZfg663b3Zj7pZr8ERq85XxnSaDRHm5FDVFT4lHYFhv5j+zA1dBbEE08a2gcd9NO
K3vGL+G1Zuckw75x6ooiJmun1TUjqlJyO66OOQfEI6YLOJIUQGaJfs7Z4D+1UuA9
gtlVLt9AXx/QB/GGhjDlI9JIWnpBDCcSJpicEakU0Ajp5NymoSwwN6QRyIde3RCA
02ZcS0KYg2eeREBuTpecQnPgDBzivhl4MdttIQvqHvmHLKHq6lypmPUH4Y1/g1m9
jXOiYi7KoYtX9RS2i0K6wkdcP1GQbLMEKR+YEf4I5HJF3CvjPWMv/F/BKlEt5dpO
EqAExCEKe2CJ2xT7DeE41rD7hXVphCy+0kT17s5Ed6qrIEYlDlX5MrnUYsfGIzZX
ztwQelutPwsLltFMLtEifra3PyjQuGH1tYWYL068dz+5SZGtWj0rnPX4VZT8jScv
GT3Ke21QLYMMPfWMfdKJS38D+EHh4Dyme6JfLVwT292rgaDoEt0rDhR2O/rjmsLh
T3G7q4xtBELIO4EJBfkeTeZgtJoD67QiW/ANYz1X/LnOnycAnxlnABjYAWYimS2Z
vusnmu4p8/joyLVMOXpkQcb3K5RaBYe0FsZ61+uZDV6YZG/QyJjOSAIWCrhTWUYn
zfzW7tWp24ZGHiLV9KWqUmf32iQwQqpEW/NeN+cGYbHMfaXe15KQwQOU+09ECoq1
nSTyvBFvqGM4bE2YEfbEYU3k1E6Km8t7dxqznMid1R0vWU1CA933f2YxHv49gQBI
ibRxLU14x45Hf0qa2IzmMdAjwqGMgsqzj3wn1xEaG4Hn6Miw9jH+nFzXXRKbOvIF
1dXfpxJh+Vt35ktliapDw517heGnpoHLu9D8jSFgPAQ8UDEgkRlpz5qEF5pRUHhi
9x3FHNU/CsjJX3HQmWa3PG3mFdiSozmqQDZOZ9a7RXR541Pkn3pZfzJuPynkTxHu
+snu0id3hKY+EZFDNo+VebbQ29+P26Zd2+eB4CuLbQbX/xFl8pk81iqOpglxAcv1
gxQ0tHMmEQ4SybeSWAiEanKjI1sa0wCe+HXBx/nzjCimozED++AdnM0cR9WamxA/
b7RBSPbF1WDinfmicfz4yKYH+6gvOkYBVqWbU/NJzYO5eG98os7ypTlmyaGff9ji
HDM/AFJ8M0DZ39gYtPZutq62et8aJR9EZ1v02Zwp2ZWyfMelE/laa/oemPUX4p1X
mIwAjsLCmzgCSEMa2ho7eYqwdCPYUZVW1XQEejf2HUJwQqVjZaxX8UYwE7pNHQVy
OMbFyA+HfU11kEDVXMl0MWFNcOuGHrHEmj/zTxFYEbjHdMQPqNYPsjbSC6FnBkHa
B/HTqmRCvRGhFlvO5Rh/vnR3THsmb+uug2ckRhtNafm5+3zi83ga3kXreAFOrakY
HlJDcHXo4MsU/Siqh1WVrO3nUKpACBSBSvrYYauKXWYkz4St+XtwjDkLfmgH3Io3
/kx6+inxzDrUp9s218WpYHKbc1Z2mg4KV00/VR/V702d1eL7vYeKj17Fb6568qj6
0utiMycEzjM1tyAfsD0DiJ3dpUkV2EhOy/DggdRg47mBtCC6rFIliX1WvgZEUxxU
ok4dpGqX6l+JYo4eAhDaEprbpxZFRevfQcakXZ70r05sXKLb/G38dU6GFBSecJyM
fmlgwWGrkRp1WYGvKN1rniySHdfJILuAH0Myb7wi9g9SR0wIFKhUf4puWlTGhbc7
zc4hBRnFvSWpgD6H5tSCvDxW50SkIv+KwEjMziaB8CYToCF/ycJksIV2oOs0VCmk
X8FleNMRLcqudy1wuh1TBUqDTnT81Ps5oBal0Edtizww6QFd0VdEjZf4LYjX0Dym
Wn3S9TcgoltfAe/L1VAllPjGDfW8iMnH0cT8EPbBLwx9fMCTMml//3Bo8b8xFLq8
Ddu5QmJF/jhAPY+FP6wgop3zel4bgHgapMZl1DA4PK51sN1eXfQj16SXdB4QMZXa
cLXtm1wr3CsXgV6Z7YbbZCAw88WO7RDWbQcxp+nUOyxDxC+XUzrhLTypA1p2xaSF
7p3Or+akxp3w3HpcfDeWRt0/k/eJtzhDWi4rbjWKTG4Y6vhlzIoYsH3eEkEQzTIe
xOt4KI17Fsz7k9+p6ExiHGZTUE6aPatb0SO1KRsJxoPYy4aAjGy3FZKW+1gMtIOe
2hzqtcMXj4Kj6fPhEZo/sI2EMHzqS6UJH5XXiysGcx/qZp9as+Je8v9jljZkzcHa
LTvyFj2lDiv4JgiSZQPgoLTgUNBEXyXuUqvw3VfZ4YrzuT5+OYo75s03cw1WvVNA
/iCf716qFtUK2qm1NYseOswUjUrtH3liYhHZwmM/cIX1YHjr7cM/LVnDiW3m4MEe
ZwPlcotLaZ+CjjARr2kpy1fPHPTCqL1fkA/OfWNXaH5lLlfCPFcTyfU3nZJj5GuP
Ne5TcMoATKGdqENUlZe60QLzrn8anwYwrq5wsGgOHlsAWuLX7y3fjwDIwx1WVUiW
5p71Qqd2y0QvriDxDm/mTCPrl7mHjMCW+9wPAaUigMaoHcTGM2L7VcpUmfiVU/Uq
yE5i9HucdTHNBZ2UoBcUAkDBBmmhpgU4SwH6oesXOTHKC2kzgOAobrLmLeneaCCZ
QVR5VPUqitpHJv42+bzsUTPxY3TNPh09tn7zVEFQzqzkoS7NKAM3JuZH0rHGJy+i
AMd2p8SGMwv7KXOWZ4p31Lw0XRB1GfT6pISrB9SW5BHFx1bDwjB5pcqb2obsfFlb
eQ4swEsK4Dk43duKsaSYmcfu94hit/40Nu0AhnDNFb9g/6RYreFobX19x/MmyZbC
9ackC0abAUdojPnwWcOgAkSt4g2tWnkGE1LdB8/OvwHkyjFYChTeXU5HClGmlhNU
IHeHd2xxKTFUgMPOI/NGmN9K8OGTrQgIZqExRYwO3NN2l4w+2pFqpnLX19D2b9RZ
ymzJPNAFKHg127NQERS0C3dQiwgl2qrB4aOX5WUMmuBNPSardU82uSVYbGWNYxwy
p/9fEuTVNx3/YrflEgQ4H0g3BZvnZKTBfTHfVkyBZFsSVsj30TwcJ2Nwac4ADpCL
afb6J4uclEUwBkfFA9Bk4PokDSNuR0eOxUChhKc4X8M15gagI8F2OS7Bi/ljHZ0K
NZJDyCxhNw6lXkvzxSpSW08QMY/51/kg7HdeIxQ6ymHIigZCutI1zbQNJ8vZ6Tvf
f8nhXAM/205q06O68FL8zD5xeeNZ0UUfylMIhNsb1cG5AmOamlKc5QOGNCzC9/Kn
3HaI5mrnn5FMt9yNyYMQAwr1cqVcl9zt1FPZo/uIPvlntPr8ZP+RErSeG1nhgh0Q
BKAVHGpFZDaGhIoX2915DIybGTE33cVeeR9Uw4PO1hoiudb9wnDB9JsdsU5VCVYI
zgAyigq/UwoReArdohr+pmNiGlxvz27oaMZVl97BCcp015DT2IilZ2uN+ShZaa6f
I26cXHHDPC4+E3AIV6GmybA26xSBFaT8VRj42E6y4SDCNssOGtFLsU3vtBantCp7
3IuozKUD+SHt7FUydp4J1n+gGJOyHkF2ZJtJq4g+Z4KsPVU98sD5mQki3emJuNQ6
/Kqlnh1J9vgmjmWVnLElqSr+n6G7bhJJAEisMeVvzG8xL86Pmjucn1ONioKccTN7
20Bi0hUDdA5FCo0eG55BPJ5NeCRIKAEtztk2nDYT8Cke99mRtmVTHc+VJk+iAau9
k+wmIZQFSB9aUuxBU90EW8Ie+q8/LE5tYS9Bvq1iPZRKgta39hEWoANcgVRFyuKp
5SDUsWGm/t2dwpmu5f9CG2gEChzsC0dy7L1EDxDAkfFg/61Oydhr1YKr9utUA6v7
5v6yOwTPMLLHzgta3rTLOh3FpFx64LUus5xnadp+YG+apjPHZxV4+kftHhM1OZE0
e39QaeKhE1h4odxVR9Lh7Q/oKcE4P1Gs9bn54/wFdfHblGTHl/mS/CKJHpNyFqm8
IZTf+lrqFXVe6Rl1Y2q6v6EW4jug9tHamooHaw2OOBy/YfkMgG7Abr63Ggwe3rdh
IOJd8Ckzy3jHmwYVa29N4ZPV/6nXZvX/Wxo0F4WTDWpgtiQ6B5TDXwI9tznGiM2d
gAockawqVWXDzaAU2TRscE3+w3mEcSwb52VlYQTI3RnGpat47eK2xsKxleYEU6ke
R2mapB4/7JS0apCgZzmUmMCpYak6GTKVYlOhbHrWpCTYgSORjiY07djWlvV+pNFb
C1j9kJWXiTV4aVkLfiMb92WKhjDJN9Urn0sIS5o7E1LRhfPPkTSZ+0sCYPNld7pq
BGY79V1qIEIX8K9fbS2595EF3PSbwqbRsWCRvuqZd9zdEFtonC7WuxX2DDBxOzdL
19aQSUcUr9UnqNqau4QkQTnn+hZoW7czw63NEMU4iPYpHx/vBSegkBhHzO6Ic5tT
GGrr+jbI7uP5q7Nnb/oWaCuDGoko2WtEjnk+Z/7J+AlUdhkAtsCUXR8zDkGqqcEl
4EVVppGkaPMVkxeGMtNK8rwc6d4hb+VYS2AceoyXM3H+Qh/nawmI4Rgbky2VTXU5
ZYd9mzzptb9Wfo34EfI7GlDk1fW/5tuD2+CNO0sf9IfXYR9JTf6tmQK6H8agNykm
nBT/C4GSQAtZFvQfDtmYV0XnIpvC6PGC319+de6k9fDK4/kywB72B4W6GqBXrIzc
NQ3DcUdgOBmp3H6RNKhishp33hfYg0NIgdirsXAsrLbby7I8/61aXLQNiElg1izq
OsMOflA5S7kJ628JbvKU2M77XK0lkumLD2yWbi7SyeB/OvF2IUwa7e+ljS/cdHAf
nONtlqpsLY3ejgMfzRTmO2spSVmCb9Mo8xAbObXCYUqLZRl6U1X6VU/R4/WHrk6B
UpXVWvsUmuj2/DJNznLBLuTfRDaP0eu1H6VMNA/qDdsMPxM+TFKsYaIpfHzIJspp
aS7RPRj/v71hyzMpAFpsI9QdI21zPVI9Nym1AKAWSrtCyNEUYcve2fmCUyQk+Plk
Gtn+z4wgBmWCRMie3yFWb/OlyzUObgkDzPhrqeGphSCs1Rfo05Z5rxu9VyNL4WA8
H9QBXCRpdsj0blH9UceeIm7Ddqt549oDiGENnqR5zqpqP9uPAsiL2+pRNgSz0i1L
/yC6rH85z+WCPQDoS7FVrg2scnZANk+M7Cvx0SE1N/s1npEmQnI9l4gt64QzZljt
VO1cUmwPzArvIRIga8BIFttMg2POjbejAy13kHJ5y/1sCY2wvpwRPaM6QUiMhus3
yPyt+xhqEIiML3s6JRV1+4R7LJeKKMuKSrgKHoyBUjbqz9NgiBDzY5gjW5rOK8u+
ZM5bonJLEU+L3wqFzOA+DQi901L0M8qCTYoV9o8a80lhPM1GWQjp+zFK5NpuLIFM
OK33MadhD8SxyAEXjutsbf03/zrOU2CnIMOmeTZDArBfpE2zRpEGk5WdwhzM8pv9
RPGCz07BRvP7GV49bh+8iKFLnIoYIROqG9yDZGNjDkI6tNR3LBUo8U2yDKDoCGFF
Fe6AVnpTdvYFrqlLqEDum9dP2DcnGzCnwqz/GYj+8ic1/kGx3Jueme9fudIZgtJd
QN4k534JBpeW4QgQnUn/8F0sLWDNFqV7EwnyYsErEzE4pbohb4/KX08Zk6tqfr4D
6kj5zHMijWnmJhLTw9CZ1eeAPAHT8I2K2KNO51toOazz2RzRm/xHN05zB00QvVHC
2C/2gBX7jGWqpFE3wUxNvDmQac42Ajl5laxeJe95a+DqNpcsR3loHOXmTWTV/tv5
b1FNgkq7H7mvM20Zs7Eom8cQyRZ0exr8noPs+D/BveDuGxZmkrHqETb8lSh2cUeu
xbsvyZDJRvtMAOMjQZJXkyKkiaW90HWUY1tlbTJNPRi1/paRAPNI19tbins96E/T
PJxIZ5ralOv/B9ggHZAC/lW9/tBrgaMWYMYcj9V6Cwh97z2X1APQOF6bLpVMtJW5
0Rmy2lU0yZtZidrIKmMXK2vqtvwFiP3yc7iNEjilzJjnI+BTxZYBrBDvsNjcI1zw
Ejrr+NmBguLgs93P3KxvsyODmltN4IAnZd+NtM3PlUrMYRu7ys/a3eNYZd0D5qxK
ILIBFAUGkHuXpON2lXB3mL+K5P0Onm5M1LjdRYTLbsX3Pxms1pxvr9/T98nbOCtJ
kFYrZ4JyN+yeXmOZgMr5ylG0tviACAj1KsqqBMdQSPi1UKUIXbpkoMpFRDzuGrtu
R46jaNWTJzRX3871XzDa0JBUkeK0hyijFhb9ksJzoUu+37un73Vn74FAd8EBmbjv
Dc+whBUim/Y+8Hcx+07ZsOopSfzVEekES7zgGSA5qkqn8OEl6/bY9wNJquNIzywQ
ePTvRSTnbDz6ZUog0o9fSOAu0Q8otG/PObArERGh/DLIaTB6DS5xwjVL/OvENI8+
G5G13KR0bVMQu4ohrBamt9wmVczIrPrBmlf4K+BmijuTithkHy3Z8ub94f9i4QE0
GUvZlyRdPvD2SFqjbdpTfDLy+s4I7QsVjdEbxDWC881ypbjfGkcdtdkWm2vg3JCe
tPso+a8DvC52CZJb42NnZ2tUKDyIS6uwln0981wc/JpMKsbfp5UYLohIJytnfZYN
Fj6seaQeancOmv40/+63OttV6ExHH9xucyD99GoWYB4bzLGj7Vz0kUlqjBM1soDw
y5RTiF3fbhKnKuXbYJRu8QtN7UNO6dEt24jkPYA0yehjyVfYfg3+jRF8iLNjBZk0
BG15hVSp8MUaogmpDeg9u+lnaOI/XVFH7Nrrddqg1pSN3HOT4KeRUT6wrUp9qyDf
CeeUDZJloxcsNXX3j7WfHqS6CgeF2rn+MCUvUZDauFI0eeV0J3b4xz2Ug3/sUwf3
3ndfN3VVwqk3PnD8jB5C2gyLPGFdWZYndqHuZo/1T0NWpIQFo+Jenu1ulVy/GjN7
ScGZUt7URVtaeEJLFVAo85xzVSUIxdCjx29T6VACwBz6dRipxagqui5dFRhFhb0t
nkZLAa1Ucws1bWWNa0v1lyP+3VtxEoqEVwy0Qgj3U1nCEwKk/e7nYITgzMrn/SxO
S1Kh3rpqDaOPeTav4rckfVPHFlHwOVtAh4Msx+mRiBLmQiI48hZev5cRAUSMbfvO
UVgG21C/7zSRm6Xw4aM3+2RUlqXDch2rfqEcw6J6tLKDbXHESD3hGIgzl4L7GN5S
Eo3rbm0tFRid/DF/gu3LqUsf6gFFJgEdP8wclmP/IdMAApSCAP+ZyNBFf3yh0zA8
Gady+YX6rdmdhGRLRBPXN6TuGeA3csdKZLA9rQ9jtOiG77/FlqicEy4EdLUR0BD2
y9Cds5HZX7WKH4s/XO/hUF/DvNCLrxc830XIpqezI5GcigFj8BaTLjrAnL2KGZMl
F+pi9kVSwLTXDdCmTFJBfwbLQNSa2Bul7QCPdhFk+AhP+uZDXdlOnsSgUODisTgL
ghvOSKWIRbjNRf+oT5DOhVPBeJwC0bJDTEGGP7xm6mTEagaBnDFHVA6mt07USypg
zmbKSbD4ERPpW1ff0GsgjiiQemBicajT0BidaV8/0Z6PmYMjuV99ralWtK6SJyUb
gErGyVW5KkyPW3lOtvtOpZ+RAdpOGucskDgcOZnatbKlPVzUtPD4R9XC0aD6b7mh
PqbZ5fFCR6+7N+hiCUrmayeVmBizRe3n6kEd3H7vOrM+o0IHJWLinDjsqx1dYAxJ
BVKQ49SAHaoTw9M58M/j5h0iw0F4KO7vHx17rXo75W1XsK1MEPad8HOhPPAg9hV8
7LwpRDAMjkeR4+Ngvz5TH3cm2Eb8goU7OvbvyHKtKki52sRWMToYXWO8zM1cEy1y
Tm+2rW22jnr+PUWC1OO/YJ8CVGuHxXZq1k1NbIA6dWyRaCCaxm7oam0h+GHE8FQH
1kDrc+vwkViuHY3DvrG+AVROkRIiY4pV/0Pz0svBBYT2/BfyIqQJzUIFELTT9lK1
pnIAfKDuydpKsKLrJB8D1AZ09ryj0inpC00JzGn3/xcwPPGVVg+Vy+DZt6PMYSvy
l1f3c/JiM9mAwyZLXr6hKsAqB6tnd/dRg00M/7Jdp0vNx6DscbFNWhIPYwOWB8uV
vSi9vOsRjmPufikwOSZZCnGDpZd1AEJwWTf0aUw0ZPT7+QL5x0p3facrmniK32nO
kypavhvqoT9W4Fi/1oKFOgMsBi8UmMnhTb/eN2RZcCzwTAp70FtEOQCsXxVKb1M1
z+VrMi0G9rzf76a1nZrEkX3B9TAvplqhw+96UAXnQmV4qg2pNJZrrQ3opvP+P369
olvywtgGtPt3xa3G3o7BcS2tsggzL7SvkjV90CQHYAeiKq9FtgxbJC+T0KmFkLzK
LjqFtUw1Wi5/MUnG2AP1cf3XLPbGNroQVP0vzwPRIqnY0EUqizDWqqC/TW2V0gEN
/kNE2nwEyQsunmmLzPa1kR2ZAIZISfZHkAZnv1inh+gv0cPeKn+SdXz46SVPKjIO
47kusgm3oYKBHi0QmhCV3+Bpb+y6w9tB6iVsnO+n+8+Ms5bvPBSG/2F9D5P1YLUL
7vaHdWtUPtabn4NIeVamhgIZWBY4BlOK0D4vfr8ClWmjjzFrYuShofdb1wOC3iKa
CVcnhmEP9KSH09QcrOOzrqkhb4PGBQXbmwSxc40tk73eBwKmHPlHSUMRTjPh7oIF
wcd72XiABfnL5ShQGy1Bfcvp+1g41GHtjtUVxMOKRTD2wbUPeKIrt6meN2Esjg7E
HYpTOWmhtNf5vbOEFUXoTqqB/xwG51flzPDbijvO4cPRGkosXoeBUzBPnSDriZYn
yk5+Ue8/gwA+T/YgFXozv2LT9+DrExM5c2XSAi00bQZy4cQbCw1HgJfr8FuSuZCt
bMM6Io7n9wGxwfC8Bez9nZtYpe5S8N5qKkNkLBLxtMbIztkaRHen7xsxw6bYoCBJ
hjIKHy/6rfwdjlGyHBe57+zcXgldCngsqwqANsU2i0V6gkzZWKwe8VaKKmpNc/62
GTonFBX8w2UVw2iNkefNG/mk+uCtVzpxFSTrS0qTmjg6s554tQiefEIA25HAURNL
Yj8ZmnNFlt+ImT6XmkNY/VXGnnt3QJGrtPq0VQzxj4exW3mM7C224lgZcQbQCJfg
fLTsuy9YbURdBH+E4DUZxOVtxiCG4dakAy2eykpRQIIWBpB+pJyKylByPGWz1xaB
jjuwPbMLAXMZ2TitJ7+iBnesEkEEGKzpqWDnn0bosbP5tXYZStQR0ssarsmYjIda
yMwHVfZRvTba6BFuYsgZ6SFVTsWR+JP2STXmzVadBdssbByRKNejouTNvFd3NyO+
HcqwRQCipJTpd2Gl/bXcT23jBgG8aTdjmyo2CxziOjANVBH6ROQJVdDB35ngWYQB
Bo/q2WH2fApDs3OBEfF1xphBVbcp6nBchy0Eccj/v+9pWU4n73AA1s0Mjmb5P563
uF+0Iy4mFo9ZREzvlzk/lLr5JSa1SLWlFTSk/CGq8INZqbd7pOK6F9lL1cxoqunX
YyRusbiMogYP2UN6LWbswkHQyltobNUQrhZmHOoPtlJtEoIIfTdF6JUkncAbSAEK
zO0USfc5qfynpHuiI4iiVY1c776E+YuZWQDMnWUPYjx9TaUXg9g6Wb9PQOLUnr6f
4hGsNOrFC4Xxmz4PXWDa8Ha+vM9oHZ7IHs5az4uhguxy13KBFI2uPVL0PUzyQVZC
IfWKoVewJXp7QSgu4S3QuofCh0affB0/6snP/BAzfuEdjgNTABxGKtlr3YIe8zKf
15X4VyIKy6XC/y8nYkuGAtw7xOHlQYtvGAU8yTV6n4t8xbUUBbH0h4Dcqo25HfN7
YDogZk0BoEYb5c3j8elaMRJjZViRqckn4ghnnUbfPExewSxzWYhem5C3CR+x2qbR
2zqsHH1UVS6fmO1WU4RiehLmTB5TbyZHKpps2BnqURgpCrxk96mewn1S6kFXUCr+
grJ1l7H75UhSfqe4mvjNqOXCi//zvLlri7q2ctzXV9HfU7+b+svA94JaLJiwyKS4
dIHm9Eimzx+WqDhDDbMWzghF600mEGGt/b3ALV0gJNRIUwZnUkCk7qP2ELzx2uWx
GPqCnXkagzSpaZSVhioRuDdml+whSrEwssW5VtFvf5bz84L1oURc5CIeTxxrDHsP
y1wyhSJnCF9e6XiNFic/9dzozl5H5E6jfiXil1rJx0qsSL/vhoUJLxE71+tUZkuw
twXfYGQlmoytiVIVV1lg+m/2Xk505vfhxp7kOycQG2xlzb/7mgnmXUnz8kc8FHwE
MF8jnG9w03MgHeu99DUp2681DdOuyMbJOKpyk5wia0dtQ1F+cDltfz32U8gEiCeS
vmUN0ZNFK/bsjSQmJuCkVleB052He4AZpQ6/HfSZ3HwqXMjwft9pa8J/mxGjd5fG
OKPa0NYGyYYM4V3y4+0IoYQBRFOJmcvxGwOb2zKHe43K1s0DHrCiyKoZOhemkali
ohFD2hJaxPljJBe8eoRZrZ7mWBfhuis32UZG/nAVHyNCkOSlNgt2XbRREUK8Tert
hsQhxHon51LcuOy3hn/qftiUBIc/ceuj/uW8kfSHIYOujLdRcmucpy4ndX+Md5au
7kQPq8FyXEJLRjlccHHDyiQkoJIDXiU8lKveGzV7dx/CY6rsKhm8gzST46WtWryo
2csbB3cAanJjhJOOyQUkmsL/Puxk+TTmhZV9GXwZvWk7GAT+4IYyv6qY8JUn4yEa
rWJaRsPuPOsmiwxZq24OKnMf7O3bgzfo30ivNFYIIpi/1LX3FZzbHNi6bXvtnGCQ
H0cBroq11n+U7Somj8LevIK0K6NLeuj5W84J8drZ4x7XF9tCpxgqsP8m+gYUHi0l
lJY3PaEu88En8P3w6QN33W38hHVDbgM2GV3rNO6goVSUluz0HlzlJO/3FdbMoczY
L7GpVIn3kzXoKmami4CJp3ZFp8NrMabQfm3XJ2FWBELsmUNRP62pHjciFIu8EJJk
H0OQ5N8HzKlpXwzzvow3TMBvB00Ib2r0h8O5PJeeX+DOhl8ZW0IdEm9XuT8fZvYA
fLVWTdGGFERj35fFoHLkrJrwGU0Pm6fJfoIw3Q/sRIa3Cl0jvnRbvq63pTjk5c0u
2tbhE0FdAwEOyj7HLn5IaeCskpcpJh7lPqLK68HJTFyIlSVVgbGdhZnVEO0qfO69
Np0b8dXJ7gFT1E81W0I+Vl46jpZpBUcjrQgf+yIhjSvbsPxfBV5TrqbfWKAWnoV4
cL2D94J5jcxM/eUGpgCPInvkXQypMexvdEGQdG+SF292d3hc6uFRxPES+Me143DN
2tBTlps5Azj7tPaHBsR5oDq0r3gkh6QlE14iybmF8FSuuK2q48q+qLGLAZSwlOWu
8sN+gPvsPcfarRkpDXkdK1evWihwmZ5zev5Uxe46na5ZvqLesuqT6siJq+BoDS4S
T1q3xsJfN5miAGeHg9+kqcoIIuxLbO4A5uu2Y0oiveJwmSb6HxRTb5eapRgP5ue0
4fNpluAfiYvUVUOrXrJ3Na9pCnUVXSClzgOLsjsKSUNQeEIbuQSLLy4CzqDa2U6c
A3VsKRlt7iObmBN+Kb2QzoWNUxVZKQEvyXLLv/cB8oOJ6BsFRDV2kped4cKgofyS
NUrT73Mb5idn4AV06M1y6vxilQiribIoaY5jCMPJQuJsNtd8hTnYjnsqA/pQMOSu
K5zeKlMe7m5Xz/rmX8dTyP79kej/ZSuQEvP088xbV4S348qcJ8AKTR/rkSuupbax
FH3ckhUsQCsMXe5wXkClSredHZEACM5SPasDXdZwpRglDZa4K63UrDKXQ6j3IBwz
y3TWSxB+2OW5NoavAIBiyWfS2/5g7i9Xf/JkW3CfllNYBGNcbuXYTr2NBLkavsQh
mCjFuTLY4au8LZ8MGiKWlDOuGi7WPgpUsFevaD/8tS2oYr/bNe0HUjTMFTQnOw7i
DBoW501NtWDf6pMALrF4d1c4q6FtunvQphIn93BCVe6+1XA+ttegdAgSatnXeJs2
PBIBiVnn8oODTVQsRpiSs5w5xQtP7OOZDevxYCUyF37piXwNpX+stWMj4ecGvhWV
QXoA7uaCaC8lMHHRpb9Dtn7xHNWJO5YCxAs3oty8y0MzBCmppGszk8E9j03Mqd2W
Vb8u8aN1d1fPvODwgmY+fgNhV3T/4diDchuLEzkH5g4l0SorqZxcUdurT01SmodA
vM0A6C8TTtzK01nZZnIJbAD3y8bKgihkJkreDfHZBj4HeS5Fedfn6Uf7n486VMOA
AftMLnFsL7N/73ypZkFesQepmaXvPXK7fPj55sCEW2CQLAj/tAfVJ4OsWWSo7CqW
jTrImMDKCM4w7z0FYKwcgHFIgvYusaAUhKi8Hh4Nt2UYptLflw5ycEhC41RDhnhd
T27hejACQ/Gbjie5yf2cnDf20m0jxG8bDLGZ2bKut81PtxrtsQ3QVwIWyftqecRu
dL/+OJVYObgknDuowDf+5kOrtiC5tJDHyeLOFTFHkdH33kCSbI6Bs8+EJGOVXteI
bKkiTxi3h9RdDfVZWcF2Zi2Cgi/s5TGtjA0d3TSpTj1agBE4Q8YV8OusJzHyroiB
vTHJxspUFdBfoTG9ut153gRD4IJFj6qSVc27Zyybm9WS9B0/GNahGVLJfNNnDYkb
KbdrDRB0BXvN6DamZ/x5/QZtzgjDtAQPZeiwI3pQ/w4Bt9DJX1WgWWN6LhscP0bT
YHM7O/09yZbHDxc4aM9vEWA08gmQvnMSoLo3VRldbXWF01+lK7bFzBSRU010IO45
EQ+nsMA15teuNysxaiaoqw4su3hkMuXhQtapNGshSY0n2YE+XvnWxKisqc4zSV4Q
+X1l+rqbXXNu2fxAJ8Yjs7E82KGmYmmjXuQTN+FixlsTvvEideK5ssfWqRcL1WUi
rsiWHE1pUpUQ3DIcSSBZj/JyCikfxgt62hXfiy1u67MFBn01tr6vAqccKRnBfLa7
d9T6XQ2cgjX7HaRP88Sz2516rodV4y23DPzLxG4fkgH7lXYCygI0c//s1SgEQhB2
GFYVJXew63l8gxN14JzooenkfVXFsArUZrDK47jtBmfkcK/63Z69Ny6GT2QS0WAD
JPMJVakD0/Xxn5v1W6tIX+DRfNM/f8UVd7E7cWM6bVFurzQITfKTmwXpOML4sHLs
3gfUQ+9ksd3uaqn2zL+WGvQp1A8bNKzl5IR+AMKJyL2cDFyYJVLkHCk75+6bPAB3
xovgxj6AmP9YH//KgQrY6/qGPhhrdzRlHCF5t6JL1CrMDnqqAgOtdFgCs36R/w1i
UOLJRRvBSfCXybWo6SdrwnI1vn7nyYZJn0fZZb4nO+rR1DjZiaysJXCJGFfB5l2R
K6aFj5/+rcXyT/QQoEm3UfLiAEvb7Xc4GzdzJd3FPzXaZZCUj/ZSgcfYoqGzczME
gTpZ769UIqfcxpGgv9zSfm368Ft5Q61NitCgGPo9LhgE8oD2JGzsF8nP6YWxjcaF
MveBA8EKgtRpjp/b247A5HsM9qwctC0cr6PtrO+tE6jjSvo0G0wZEo57Z2c9p/GC
MQFd5wQ3WiOErZ6EVvxBGDYTKpbDk4Z6CnE/PL5tW87KqptKErArq2pGpM8iGbcb
OZgahlrvF7siaB1UBTh0Oksude1IjP/bmS2EFZN1CcaH44Fdq+KNRHF52VdTh706
pL1iRuocRYPaAcwMY//HMvOygVNR9pVj/HqXjT/1OnUuHEMOmGLtWv8uWsA/lD7Z
1flqFSokiuqc04+GhH3d0kH/qJEgnsGPBf4Q7xet7z9M5d2zG56IAHgABEunv0/N
BywjNQMzGGqYX7vXMCQ0L9Md6KxZ/hL0FJomfrb2keb6caz1lb2g0bKkVoYwqmjf
SJa5Mn0I01B30nB7y6NqxkydqLfJ+U4gMYbT/grA/tSZXFoUBASg3uzMCid/mk2J
al84bdrDKLDegL6172/s/QJu8C4wMkocSwYXz+lwRIfTOPeg69U+aQPDLmoZnaX7
LSD976MtIWvjUYUugBLEDr16BmdBQXUY/0rqr0XQVTO2iKue3wIax+1ALK/zhCtC
xFZUc8b5DEQf8F6ce1Qfq9tMIUn3BcqXNyqkb9U4oosvMtsOQnMEhbzeFruPEEDl
6huCUs8KNcMgecI+RrzmVc/MNuTi/FIp1uEv/aJvdFIjrYRVq4nh7mo8EfCU8ih9
4Y6l891l2rZJueZUiJUz0TCHciVzMTKuUMLt7LpUbLGRc56gfj6q7JUWjAwYe4+t
fIr6sfRp/a9915RxXKlS6+NMwrhRHDJLPH+TZzEZJ3uhJ8XV6WKd/6JT444fzq4H
LOArFjV/ENeE00NInEwIZ6eTt7xB5Bkk4OPFI6QiVmtBbkyVtcnqIai4+p1sAsRp
QFl11NU2I4zNAF5SX0NUeg70lZMXPQnAMbwBWm+yY82PSr6uouoTTE9ddRSardaE
Wp1cTZP5GsU4LfiYImC2fQhuLxEwlusKzyxIdn5Zl7h8i70t27kW9ubmZUgQU4ht
IU6fEslQE2mGvzfiz/t+ZBM/CDaXUgJbrOdCl9KBSrRTdpHUfaNlEfgGYTgj+J02
ojGZdqrhiolnwalLsGxCixyFXflF2iqD3IMpHj8bLBGH5AZ3m0lu/fG1adbOYOIs
tPT6r8Z7sEnAbZ3zFtYkK/CSfPNSpCBq2o1v/LMd77Yy8GzYSswrXTl/8W9UPx/h
5UT/WG4pxBUwqb7gn5YX7Nz/+vbY+LiaI1pE3IA+/x+Bi7E1y9CCFd/TM733Afzx
97sxvT8GvsnVYfi0IYinwxQpfjcnIESxHJSFx7SkUD2VBPptIGufAMFchq49ywBv
dw+v9PLQIfYQywJceB1vkI46M0WZs1BBVUKRncju4KEUOR2PL43X8qzM+ZjhpPqY
Tbo7ptnOefrdQxa7WTQRqMdmWZjsJX2UfndDtD/AQcrr8nkyctCC8Tm99GtvgohS
lBwAzJk1x7xzhZd2WaXdmV0Po+2SvSoF9gVHVoI8KjA4jOEXhiVhGv7aqpr5FmEf
B7lFRsRIRtXOGOy5pviv0ZsXCOGaGhfbKsUH6GRr3cjaAuW99k470HaQMLAQx//x
Yfl2d8/yeFoNqSHdlhNwazQYvBcmp+8VuM5apeMwkTpsoPQkebDgzEbS3Fo9jRab
uirRqCoYOqyySt3c0gSKBVvsdkpBFtVeVr90n+9h+SEJwJlgvL7aRIs1WUminw88
gw3WRbuygKfXIysLEaQGicDlTMW07MW06vKKChIn77V5KmDJm4TRl6qPRqd398l2
eZriRGnh+ZPLMLGgSwGZVkysr+KIUrwyFjqbI7tFN/i2N4gMRootbLTx489mddm5
Qc2ppYT7tMjq9tQouRrwvrig6IeZF+HOdYsFZp8HOJfIirq1DOpHOx/kxkykx7n0
/bugkYIEuCM4y6mC7MnVwk4s8OM5unYOGbYpgr87QAUUaW4tOeO3hGvOypTFNfW+
xT6U6m4UL0a2xPQzADbyATYEU2OVncaSmS4GCMSo6UmsVexRfdF6sVfmkFWtfZo0
gfpSAWhNKnUKqh1evsuMXNBROdiJcvZpaOXw9SZdzFqVqynBHNRRdyAFB739x9D/
b7lQrN5RvoBbX3XdhBNSq2oheMV1+B3AmfZqpoX53CnBb6gph+kJ/tWb9JG4hJlT
IkSxSK7fBVj7rPG2Y5cVgyT5yQcqUuxDjdvR9szO0koR1UbBE6y5T+GhC9f9i0WM
Uh4fKHUgY/AwERW/4/0VVgDrUP8Jx5URLP4pQAmTMhqZzdegJub39QpzAOErupQ2
EuEg8MOe0FQTZrbglaMrlx/O2LMUWv/N7cQ7o7DwRH5d/vFZOZvCmdmO28jH8ARl
dZXMcaswIS8GS65oCSY+6zmkDxAfjgXiR8mgcD/b4pi+xEIx2vtHNVHuhEavWANY
3UsSFmVXFcuFeEJmr0u7jFRgN14BhIyo1cGta3JMZ8XGABt3K+8ObCbKB/6zHOSD
JLRpJnbkTdi3W7D3rugvlM4A1VdHd3Z9MIgUJPe/ocgXqGUmu+NYCJmP02w9jOEw
AeOXcyRMzgulHkv7qF5c+68GUwRqTfRgF3gNrb1+YiDNbp9o25xxTHMeYtqSiy8k
7trB2S10onMGO3v9UF7QY67r2gyx7OKh4woP+AKgWIZcZGEH9RDrjE+VWrk1PClr
0mP6EQQKz6s6Jc2b/xHfExQK6LYuxePeNkvDnzqWAAe4pYNwwcPHwGAwJlufERwO
drDC1+AbmwDMta7Q3qozKlpImmdo9w5rtqJ5QMbfmUeK0mfnTKIJ6J1xP6ln0Kee
VgcLbXSuEKO1rpK7A9Os9QVuzPD/LCSUlaV+kQIV4CGq0Z5NN1AEQhwCTpE3PH5Q
2v8EKeorZVk9YpGxcWVJFfafLTpeMqyiSl+scccR+G7gjNO22aywBfFN0SV8jBMJ
LvG/q9G969o+z32bIpWLoidfC0Gx75l2leQDzA3b1ki4zBLg5epOtSerSpRow6Q8
OWA0/3jvRjulBi8N8gHW1LtCRrc9XOMM/CENHUuBnMDrFRcIRove3O/Nxt8cQ/1J
v+9/Bbe8xNsTC5HMWSrqeRFeWvxjMiYmh0mmIfqL0eMIemAUoOD9uvVpAIE4i8wQ
vr0gg/YQWpjigw8OKI9nYnO4i4cBkTWbogsYi3J+2nxFs7ekI/rut5Ka03TkabQ0
XAkYO4XRuKlrvozV3S85HhNdjTm5yhHul5yTQGpJgDePWBrP2tx+RfMgNhylKSwQ
SOVKyMfM5raOdXKgJUdhCpldhpGvbAE/ud8NWfnyyAklGDxkpb3oNxYYjAD88II4
QaJV5W8Z/mVZGAIAyBgVlmGMCwQdq67f1qF93aVt8eKFKFLqmW+7lQDale8r625l
KN4bp/vOhyH6PqjXBhs0oFxZAa/GenfcPLl8Kse4HBatALE6ILZXz8wBY++yVj9n
ZRruTYiTIreg1/rVz9+yt9qQGGm0dm+SIyskP7hhDY9eAhSrU5E7PmWKF1I/cxaJ
bHP0uIi9YsYfn/uYOIAKoTnKji2MlIo6nwFmUWt08LGoQ1Z0SDJ842eohRxGcK69
xJ6NCazZBdfkcl3qE17S1i4ra3YZhT0vdv6yJ89By6lOTNbdmE7BzU3rnED9wzYc
VB+eP5Y5IjXuvic8ku0L8QXUWawnwz4DuatNPymk43qQqghig8wOH/xvn4WXwb0I
5gBELBIjXuL/bl9+YS794bW51GxdBKJnurIdLdeQHg4JOg18jWzGoV8ltTtnTdEp
H5xsA3HIi1P42pRZk6oo7RgE8ddCM/xTiztHcVuxq/MwqGmxdf+FkSRBCCPLG0S9
V9zepxmfegNmyKeVCb+Ri6EHSOnFp2+8YFVKI9fvfwp4HFSWoqbWkql/aFH9kZMc
PB1RV15GceTitcydsKwTsW889VpWXEXlazzYP2GCP2OaANUUBZ2wq/jTq+76tmfX
q74x0S2hZydkqVZc8ycdrp6y84rPHwfW8EU4oTt2yJg6+U4NyZC00cZ6ykwfS2U4
4B6eHH4AP1ev8TYKBCfbjZmarTj5EMTQcFoilSRv12y0h6Oc31BmqFyxvcQHHQrU
G79cIBvQDkNTwBsCWpj3mkCdHJptbaLf6UdLiNk5stWShTkTBO0Dv5ILA4AkskH/
G6dbfL54jUkkyR50uwWXyG8zOnFb+pypyVWx8FDlkshk+S5bkl3d8LTY7GYSi8JC
tPOumXzj2HtjEwp7Dzo+Nnj9g08RNyb2alPchVcNlhM+tl3nc81Yfg+XznHzF/pt
imLLk+BiHhJhzhcCb01RTP3JPMuyeDYHPBUMfAyQ55wCgU7IGuxZEC4TZ77s1GX/
SrnUTjaZokYp+7SGqsJ/SbWX5rUmHy+TFMakVXNHS0U2Z3YmIyTqJsiBLkxM6z72
JXjjK7a1Hl9zJRmPNm2dvt1PBWuBspqcy34KmHkYJUJA4YPGb5P8QE8l2ubpVlAH
ir9HNYdw58CAl1J7idX074D9il+Y/adBtZ2/ZZhHsaEzsPX6V57E6QgGxoOQwlnY
SjnZXLkT/Fe5gqeyfOQqECsFO+r9X9b71Ma7jYsDvYGoA0VJzgS6CIYLJaS6G2rY
qhv9Ah4mXyKWYk3ADBB1Rb0WDisBbFStmI1COKolmoQBAsZhwoIRAdu5StDCGeV/
giGvAewwFP7kT5H+dX7RP7GWqCy+/ciweI38uInx5L1N8fXIhasR4vvGrco2zzdV
RC/dL5sZJ+VIH4HUB8DHGv9Uos4UchhcmUHO7e1BGhuL/fGoYnxYGjTNFeU+XEP0
iH2Juo2AjPJv0RUZq30r8WoxaPBllJ9YxfT59COomuBhBzX+eZqCT3uXpIQVSRBu
fKMo9G5Cwdl4kxYys2TtZRvsKZH/TIJ/lKswBZOiBy3s079OmNpY7CLoNMWBFpKq
dIBjIwvER33aaBqbZ3yEPBt+9gbyqTo/inL+kzznMpQAK/NCl85XMYr6JFXqTrLC
ulkxq31eyWSsHITlI18cyWK3cMvlYPp5ycgU8koMX8IPMiWSZns7c7f4zdSFGWkb
FTLa234A0sKkE1D/7YoU39elppUg/WTsRHsquZhntI/OAdwJrFtvw0jKsLFvmbKp
6Jq8yOaoZEAbF6oQgR+MAivWaZj89deovDQS6rgZrX5oYXx6OCxpW5+/yoLGmd/E
q/nlTWE/eauJKB1VnjzxuS2rrPe4LVBsjyoZK5eKes4AIeoQQaRFqJPHkCQMjgsP
T9NEk4Pg9OAKRSTY8Tq5il+9By8Gia8DQ6dAZhfaNFGNAwD+x4RgN64Bjr3MOLET
6jB82v9dk4TUGj6edIXWIOn7G1lxkkoUO3a1eQSU1aODzz5F7gZ0o7wE50/VHEpN
du5E7Mcnr5oqiayo5s2x8G34HwNw1/e+qkmuXCOHcy+JTj8/HgHEIxxzK43Gb8zk
KxfDYxxDX9IKDIXvMPIEqAe9LUmRyGMM9IgSpAuJD1DsanCE/+UPwy31CltvvuqR
GIZMksV3yvXLRKXzuzyWWDI1ML0hRKrJUpGWwTqApvoHqNf5ra2+T7a74nYMR3os
A1D2QOH2vEs7Ha9usLLKwYlDL/HC27+D+Boxvkbx8oxVygRXmqdt7LgCAQcEyNeH
dkP04z0//7fo3W+n+cnSRBs53aQGXwXQYRhLTJIzOUIZ4ogmO7BH/MUUODui1+Xx
+C5c3+h0n3F/LQnAPAnUk4OvAVb1pbNN/b2WgkHPiLsKqr17rip0BzS++YdVaCZe
b24A7LRQSybO8VxVquM27mzFvsagFqc59E+y5nMBsjuxLw99za0HgaD+jm3pCEQy
9ghtM7K22DGdeohxvL0Wnh4Dbj8SP9EHl6iMUrHhYg9KR5pQ04YSq+C22d0rG8wA
bysZXokTV17KlTv3ZSKKjkKY76yIedeyw7poxKMIENdD6GkxKSwo17j6NuDt+2GL
wqGfFT+RnBwUWp2ulG2zXzqRSHTO3MXBjKUCmB9qyGgW2OcmvrIjc/9jaguycIVe
crp8a7ePDbK75yapBxJ8Zj41/MqfP0IS5UMXlfI/cB7BNpFqnnnCoRTaKWTUfrr1
8Bye8b9FQ9QdCw3t+2hNIJuTx/bC9TmzDLoypfM+zYntB1y31sK3GMPKRbwNpkPC
ERuatph+r9Y6LqjFTZ6O7VILXLYxfpK9u8BQ89IIZh0DFAH2o6jfcrQAE7/B7269
PPrA2yybcFcnvTplxdvZjRjQMhxPo7Y2+QN9aqtLYwCMRIEc2d28ekQhafvl4FZb
+LEhffa26J76Zl9kjkffwzj/qNPqT7mlsw14N4nZ5DruTL6E4AzhkQ+e91oOsnqs
Uw67X02BdV9mlL1+H4BkwlDU0ouyrL/KOBetsLyCBwpE7UXgF5DYtxTux8i7k5wy
E2eZb5yPm5TnYyTAFOtWy29g+KGxbeIB/KABlqrjRmoO+MQYZv4OvLGAfpbxY8GH
B2y+exBQqn8R4H+ik08YDZHiFKSKEk9Z8MrEdzZ1PIZe0HgymUVFWXENmf2/eCDh
/KxFrSyHBAcOD6dHjzfutUrUusUEqpvu6f+YIm1B+awNoZoOTTJk2KqvReKBhzMq
MgP3y6MDF3haiw8iaM8sjEpJt5MnJuDRGtylw5L9eDJMhoy95fZ8rv0EmS5XI02G
Gid/gi70snri0awsWX65V+V2kD9PnZ9ZfThbRbA/wIiYIaquSzOT27jytQrODjjW
2FlQAARjQrwQAEDPNFDOJ+xmzhGbtU+A8kiGElvrfM53YXoSHNFY6w/peaPAPOCb
jcoqGbi4R/z9c0K3Y+ybuPPFWRnwtwwQm7JaOJzvif6DeIqX2zBd290+gS9Nv9sF
jqvdoeh23mLnW3ekbSIxyTO1CR5UOAetA13DyIKFD8eEEK2d/zrBGvVkt6G6cWyT
sZtbHcxgmIbkG3QLOWcfin9L4dZ4c6mRz8pWzTPRkIXeeJjb7YtRrcaAs/YNIAnz
jGoW577v3KZmpcAYItpvhtng1Hr1cmKU/qmRaQbK6IWpd8nJknxhPus8FO8++8Z/
mkyOPOoAb/FfuG32FhqEzIWKgoGfp8llNGQP6+fRu8DHBk2ZMQIywuDUP6YgRMf/
dK9d8HwXpGFB+8eNo3qmYszBeqHs0yS7PndcL99QA4ZeZZ7lUeAN5LT8Y9g2S6ro
AJ6NTOemQQtd+qWyPQZf+2Rfj6wXmIOip7Fel40ASVnskHQcQtYEE/XM3t+ysBQD
J5oRFOr5ctyhNumgh1GMgyLG2+o0YSZhA211wfJ5aNHcYCs6sKFFZnlyx0RCLJY7
8CmeWagiM+d3f/MjtsfesSzon7vjABPDDPI1JNgju34YGfw/mMcqn12waumERjQL
jIRSWMJS1yyJwr4H6BvAf3rNIxyt3vKZeo2zB3le6VQ2l+SLiX6QuMCFf37SY9Ag
HjsenBOA+IqXnBCnR0VbJ6BBTBVGqlyALPeeP+Bb0hwHOg83Ajo9jSNE8sQ9SxdW
uIcyG0OQvccwv6VV7I1EZJ2JPCyiWg7mCduqJ4mYEGGfuTTOCf0xLfz+AaNhsstn
hqtmBm/1ZtIEw8J4oxXonlbkQc1FIxR7MXodtMv4gBlivK/g4a4m33beEoiX9CnG
GoyJ+OnwbwJQY1O5Itd5ZMyyi3O2c3PQd+KM3K0EP2usDMkLgtRsKbhbAsFOBQEd
nqjWV6oEKraE/f7wCLizTFJLPpYHrFUhev0IpFVs09OTwcji6M8hKAEzyb0qXSX2
sN65dfNA3hEWg21FoaxUgKl50P0z0ypK4Huw6/ePQeDlYFA1kvvnAEwpuYWStBE3
g4Uj+btK0I4aYMQ5aQwiGNYmbaLf6HyGpJVjr47wfNzXe8rIOtRMyZn2AXSDhnKQ
lS1SUXjN3mQxuiQ00y6YHZOuYp2g/vPsLnx5Tj8BLgaGYYLvyWN9FbBiPyBGCl4G
hHN7RDtujmv3UTL91j+wEofnHBUeGyvkvf9SJjfKsCLyaz4gWksuJo12SUDkMRmc
ie7r+0XjjP4pOlXRyKu2Gf2RDMlelrIM9hH/8AM344Tl/+CiMPbDR40JUN+pHw5z
beYI+bivmiC5+rSe5DRn6RW3BpXFmO4OlZ9oiESHD/F3eXOuHREvwCqiFBGoz6Cf
5bhpLc9UC8Bjq3jM5HTnX44p5n/xLECWfrYa2WRBcnqKSyDvEK6Wu4gaRqvKCXB9
ZvFZoSrKvMvoJPHX+5eaKH12yPLd02yfGYJWmilonMeuVNT68XRkNIDz9Bx6oDO/
ENJZ7XBezpnXZvCQ9Oj7WdFWUf98GvYESsaWJ4dN0N11U4amn/hU1HRcLaFGaMPh
1jMQp9Cbfm4BcWJBBCZ11O8j1rKZwYM3nt4KQaot5eOdnVrzL5sh43kaREzszmKW
2vLUD3+s9BKLS5c6dRKqoXjKkFvWriP1ef9S5ohSfweffx3v0xhLEAUp4E6oLMkD
+ferjrWrYXFqfc0eO2YDH771PPiJ9Tz4ojJWSECH4feGy6GRbC5qY2Ltooh3b680
+QvS2H5pLk7nq/yPqIh7tncksBPfuchKx2Sb5q/UuJZaIwAwAzGUUtylcC6l//YT
7Krh//ld/qBq5IMh4YDDlCxcfLKpxVIvBXba3LPrfJmBJuqdkKtjb8EFLOcXL5m5
c1W7mgdp2BS8bqRCEbTcbs/aE28DCQz5GeFwmxJ/Ou5VIL9kRVtu5A6PQV2N1DsU
gxd0pfTvmMiBnbB1fTVyHVWLAe4LabrCFkxDwTaE0JZoPD+XVCgUC2ny+Uuvue7K
pC4JPBQ4RtXDtJFNSSLUt53kyd3PrVqO6931h7stDZ1fpZwVMqUxcYOOWr2WdKHb
k64xRfdofuIhVc4L2Un60cdRo+e3KtFrUYfVTBtV8+T86L1T3t7vLrQbOQt3pZO1
lhcvKTLv/Qeb5I+LAchrJ9I6JGi/nCe6Onc/tW5oS5Qg3bGeormaBUHReloGG3+e
83ccI820eW3QMypIAL2UdrhmoE8c5WNtcZB61FnFgaE2iR5pukAybooSpANPCgi+
HMlDSDiDwCbCPLnDrP6SM8DFuNjQ2p957wh2IgCITV9uDXDXZ3vKcZjZ8SjJj1r/
lctcY+fw6AEe7C9rbOHouFagyyz02PpL2d/yutGLF+VAB6f1t8ajnR2TjkhrqhYi
bC7CH8SCB12V+xg52Yy/ZsbtdanA9r39rwliWoJhf28lWQVWD0Ip+ld9YDBRNUeJ
VO3dzsqYKHnb3G7GhGWcDuTxE8SxKDSSdvlQKDqiNTuzB8oDUWp4kRMenvlWYnj/
vStC1aWQ69SK87SBv/C/Lvc+drRe9MKPA4afX9tZtqAipv5UCB+jrtWOdn7SxWZ6
UaxxYFyTmhz/BAUKlWoz1WuP1SKxWo2EQVmfZwFk2iWjj5Ih0jhVm+l2VP2fxGz1
c9cUFRoWd5qKNcZIWW7Hgm0+6q1RHNKc+Sr1D8pRtiR6Wmwy6COL2gi8ffhrcfXK
Gd7PghRnJQeo+ZeVqS3eI4diqvTU4UPI+xv9HdRHr8IKL5slo0Jq+184jJjdbymS
ZwiMyoRdE2zR+kAoOtG3ZrNqN9/V82tkxW5jwsFsgR59GTIXlvXC4mQzFCK3/Srf
u2LCp1gSbjtgQ11jork84dMxmrg9HIo/dJ//8BJXY0G6uQboBtqbh3Pfa8SWXycI
GE1aePyU8/S0HUxXca1hZ6VhqjOodBZYTNywgXfcwunXrCu1Q1v7ZUIftdmzYh5h
42uXGcyT7+h3wjLiQgTX6q0EmDOlnwXoTe7Lqp/wQZcU1keOFpwXsBVgL/bkeJKA
xNwI2UfDWzVjxwFFxzz3lTrGNfyYae+u+kMKbXiWbQgi6OVCqLJ1s1DIikFgrgE+
RMUCus+ycNbxSCHvwBO3S9tlSCD3KVK7mQWMWtg9ftEh9tG4sVc+libRan6wowcT
BpahEBxZ5K9kLgA7DPl0qS99uz2LxIRoNXg9GKkU/COiI1oFnGnFrCB2WHCRhVAz
r7WFUTZLpzqfdVJB943mKFeAxLf5o5qPDizU02m1j3VmPMEkh6udApjlc4F8AJM4
myEq/DQSIqQ/XC1s5onMMqcwGWauV2JdU6RIolWvQ/EusK+E12CQya8JIDmyr8zC
Hu6IIdRysCMR7XmFrRATK7JWM1NIPaNZBPeVwRiHO6Sos29tTw8PSrgThGQnOWmo
fNJL45CpuGygVmtp5cjr+XLGQpmw/YaA/B8GfZV/qTs2AgnPjf0FhtELRzL4nAwT
qopMROsB02mtty56RVzg5xxPwl2wf22oPUFlgJaV/1cuFpJpKcU+c6F7SlMTd/3U
svcyiiFQQ9GJhOoq0pbhDKxAlzGGSskFJTS+0yj5+/7ZSqs5Jo3LKnnKl4dqM4Bv
/uREH0w+8j65n67IBwNhaN3Tjuz+GLnPy84qU9NvQVVBBEaz5dOOuKeloxTmoAbw
79pzNIsIMnQ75SKyvbzq2joCsRlHA/WWgrxSOkEQlF4EnOB2+ESDZ9hUGpzpHVkF
AvCuBbuu5FjTMnjkKYaxymxOGTFYz3rW7kd7X9ZCBlFSA7Lu9z3lC0lAlyhKNDI5
haDCIW943oaEWDKI0qHViRs/iQ32oQ2WA4B+OGgDGX5omLbGM7uqqScB4FCodeXO
l6RUpUGyHDFztgdjf+2o0fNtYTzaW67XEZxul+1CDGJekueQ5vdnclBetaNgFdPQ
brSUWCVjaf0HDQtKfjlnMNuK8bhOUQ90bXMLuh8h2W+7IOiMJhTYd15hbqZxmph6
5x+yTmlcXNPTrKcJtaLeFlSTtyW6ZLP07lDTmDNImg4B1GjMG4r3EUn58l9ss5pQ
X93MeEgP+A29f3lmL6YU+idyBFY2zewXWxqKBT0LxMVxNrlBgi8HB58spnVYCqwO
oBfz1A25euQPE7sPYBtFfnVWLo9Uy1O4vmlaXjckHcByfznnopmppxx+Ja/LB3cX
P851MUi2yMj5qCjzBUyW7HW+Ey/7wOcESY3gulApsOTtd2WwLQQCeL4JmOM7WW4Y
PNAGVhwJui22qwXjIfmjpb5r9P2iC5I8glL5bcCGVY2NrSZ/StJST3Ls5XCorTdi
HuGvdDPVCHO9/klJUFpwwAopc8KXgWu58P9v04p4VzOayUTpSxwekrcxP8lF+7H8
/aA4BR0Q2H7XnyYbgiCy35TrR+3pP6FAqbg9mn4DKwWPXLHz/r6fvG4fEAzv3tXg
AliBYquWjax6gtbFrHwC5FIUP0A1qCEdPS9mlv1BTNykxuCQHpgwugC+8/ZQdSmH
7QsCOc9PM1B57/kVqmvSgDxPQcfZoCXZSU6rat6PmsRPNqBsd7I/9hjaOKsh/nnE
hkxg+YCm/6tqJqtKTc9rN2geKu8q+rgIwNIq0HX92wF0xJFqTf4EppnCv6izIsSF
vn1r3EBQtfarbG/VmQf3CLC1csPDxb4KLQ4zGwqlxUrHbc0d/ikaJBJU9LwvxvlQ
XaFMzXzWLZB4n7uzNrrRyFQahgqqlRXoHHk3OPqKqeV2tetiu/pxuy7RHFzi+hAi
1Ct2rnN/WcZv0yl7ccEiWHNGrV62O8h/5STLilCfse3mbQ+W370llEaDLOzsq53m
trQcTgNXgptT9UlXhOw6/JF8UhnSINvffTrhJtsnOcp5Fx2CvPRHvyDZuikjE7Rw
11BuKyoKSIFJ+pMg76j9nCbZNerySaZI4Wk/VFuvmVHFzw/GYDJbHjrAezkwlmzZ
b42810UZg2twWlVEbJpoQzMPIxcMoU1oQfKDxdTYaIgTsdXlKlAIq/8Sy+gfj6CW
TJY4WVSuxLPywltgefMczJ568yDDkZIO1ngdEUZIqH+oc/LH5XS01rpuWn9VXdUW
IMGDNsgDnTY1hME4dy4TzNK2//PuC2cOllbvceI8+4gwoZrJmZw5CaBLubQI2Kx+
mbKcnSAQUOsZx2fFBkKoTz7g37ceQGFSN7ioGCficjYFLCBEmK9TCqD0O5DbIOBp
RBqaCa7zpxEc5ikukMGuRJmOCN9yQuv2CJZT4WDx0OK9oWnVYNgLW7/T9xGtccQb
M0cyRO28NhFV2Fxuhz78F9F2khdfsK3qT/ghoFdg0424U7fa0MtP5aiduZZn4zjf
27PxhcojJfChQGjy9VlxpxEdoiBeQ5E5KWMk5dO2tZI/vO60bWtRajKZj2xEClP+
MXlwAtPuG+XHcpG60aUxomQ1tSz4ow9H8hmv97vUn9HfSN/i2akNs8ArPQCslyff
OtURrR0XuHLpSXLZVVwBU81//w5evRhl6E4OSYE9I1rEagF9ELpQe0uEfIBSlcsw
h4DKY9zhyruItwDrWO9LdCeHy+bKu5YSACw9nkB6qHMv8mjqlsA4Rrx0PwJg8gy8
2DBY6goO9HK7cOQAMpOywv029PZon0EvoA8h1RBcHh80HtSCTJygNho0diMceVE7
8M1lCa3iO5qfOhNHkmXZclF9hZllntunpOmJC07ClR3xPd/AHRro4o+veFtGfghM
HOfsDeazGxqJYNABflHsNHaLL3T2pw5qE9khzFRJce+9UhvK1Fru7hSP586EgQZW
0CyO2etUnWIZ8lExsjp+cBGNi8VA5Geya9VOT9/LaGRzapC53e3rouwATQUHyTMS
urdeweQUJFe2mLgVcEtw/dH/bt3SFYIa9NHm5uHQJGNil4BoJRQKJ3cv+ydCyUYv
IfUsEiYQYk6HGSIOdsIBvqUCJH0T4STpb+4VoKuhM3sad2a5YFcBFobjiq4GS9eo
9DxP7NsgeLmFHDQ4rlYcOXNdwf5E63eEhfTDLinjLcPVpAjhQxNpnCswK4M5XdZa
sOgbVqO/bw5P1x5Yz8sTtUpbmtUdCje1zQnAbTJHsCPlW25yxkT7087fiwJXQCzb
uXRkwtLHekvnO/qkqw1ey8VJ5lj/7+ExGqrb7X0Qz1mv4j52APo4BJKhAwjRY5kz
RVmcQDl1eYt7nsAXmBWcRIQz7PXmjhlZBbkXnPI+2m2vVz+FdUVu5jHYgDfOFEgg
Qw0KNzFheKBJCN5JSTC9NM0zyp+qL+2B+EmVYs+YhSC+Hi3RuWVSiP1+xYcAG1ri
/FYLsutSIprUf33JHLIfSdmtRbh5euWHyoKrg0EXuUxN/+/HLkzFBBWBnM5VLGwt
LWqXm29QlajLXd+XNqwiGKauSH30Cj0F98vDP3KoJZ7F5RdR0CHZmqE0svatnQvl
br1hcePWRg4n/sP6SDFBCpN5to2b1Nw5LwZj7fGX9BXk7JL6Dd/8SDf7DNu1r4rO
ZpIG/sUBupxQ+BFMC6L6ErV0BEPlVhHXpEaSmKSLZAtBE0utzIvr7g+c1GODLhMg
SwcpnEckT7hhPYaBoOLSecJ5Md7bO8GJa4xvqlv1UWEAXyOYztY0vzZMXGxXqLjZ
+m6E6R8wj9qy9d2HXG5CfZUgutTdsij9Q6w/QVwKMNocCqADZzw1QFbzPshxthfr
g+K9o+McSOzV1t2yrSiOMaE+qkkxjAPGBlV8oLIGj+GXHV4rdrTiLeieSBZZeZn5
6CEMhp6DTUsfc2mzFfWje257BYW38ZwVGVxjjzIoMrndmcV/LGjaZ+v/Wxfnb2VT
P9GkLC8NS9C7+DTFXOkanA4vNP2I/VsQiaSQMaPPQJ8K30Rl9aj95Qxtcrk0EzpY
A3TW8Y97ceY+uCXeFwikFHBBuw9vNbkhBgq4hhgNjXQk6zIP8Zh0sa17T95jFclv
P5DyomPRXiKRmAS1sp5zqf5V+N3mxERFPZjreSFGu/lF4/OQV6IT0ms3OWOF5N2f
vaAXNhJRePfJ1bdr1hIde4IS/VVj7ohzKr75I1jf9D2hGRVvu+tLEQizITo5lwve
U9B0pStoAAZ19A0wfSiXD0L/nKER4VNHFgZgHwrhgkH+UB2h5P048igbbEJMW37O
oplphIXmq/qKy2Ma45DJIzAcSDD4fOL+MyIcX7SFTjIL+4ay7gIguX+KbC52LIAd
2XoaExATbP5Z6tFr4JE7ZQQQsaGkHQXUkou6GkMutIJNkbz6dDz4J6AD0VhtiMaH
PKo2vks2nybUWj7N894na7SLuSbfDuOTMybvRG9mkv2zPs2U2JIdADTJAFFmYCZ1
2QCf7UifoTu7d4g/LcIoSoRyQeqiTsUfHkUElaIv+UrBcOtaNMxcTLnUy5gLaCFv
EuxQ6jnsIV+ATqkgw0704TZ9/J+vmXNS5DaodgS0QH8xRgX5ftlw3WMwP+t/F16L
WQkSlg/ZG8fGMBxtYC7GAke+D79Xcobe6W8cIDH08OJGPA4LBu8pPkrlwxTB6MCv
ldFMGDcEVk500MVRwjV6YhqVz3waXVNAKlEVwzmANdmj6+Cz2ulzzHN2rkK741gv
OE82I3k1wl3AwyN5bSGYiLp82buCXFBFhmCuTD2KlI9EQLz1Ktc7bdFKAvHqeRly
T+TXYkCwX3e1tiNQMYFWkhS5hcpTYRAX5lfA6rmL8U9cSHwrZTXpqE4lBfWYw54V
kIE4pJ0sHT7YFHpZw5FaWDKhc7AiZLMTjyL9yKltlu2V5IaNzrWXt2D5cmnmnJkg
D/sfz0IYZtkIQAYPfI/lVcijPsgdye3IKnNIOwt7DecXml+hePdUibePukgcA8ZS
pPbLaMJllqNg+3yUM7VXEA6MhjlQo/09mFDVpmk3RjU5eecwtrWfmptrILLTeL2F
JfGdbYgoZsD80oBxQ0jQwgccdPZ4gLWxpAwhdHSsSsUcZd6qVU/D+EBw3+s9pf9d
hnPMKn4HD6d6l52945FuzObAQSwpbUBeW3SVpUV9apISUonO8iUq6oSpl478eGvl
heya54A98aBl1AMxmyHnbEhRqvwPfQaJntAbtaPmxJt7/sfEJSs0irwgLD9sgrb7
st/YIy30p8tGMnVI3ffLpAANyWdt0lEgTFugSp3/P97OTrDg1921zZtz8u75U9pY
gUKqHCe4gisaULZYo5qUcVCdX7uMERm8Kmh8+Ok+9Z4tzk/rMCThUrL8Vc+k8KoC
uXtOoFzkOX/uhpesE9881PryBxkvlIuZT7Azin9altWKKcr9WvZG0M+EBmrjNfS1
u26xhJwChTnUS+9rY+mu2NsWW9B/8pv11jvZS5ALV97JCplgt0T7ZAVHdvSy+MHW
8yto7FB+nTdcCdswEK2+Q9RQDac3aEdft4azvgEkHflakihfZBCc5P2EIVhGOvVf
RjzybxU0gpdjjNrPARdbqCEMDnhtoVX9WadyeEXFLdzH5nlkIlp+phxcXIHVZr08
e91gjaG++RLQVQe7So26XohLQgeAehpMt4a2M7TwYVWOwnQfMupy0c4Dq38m3t1w
++M/ByZn6foHV4S6ck1tk8+OvMCxJfXrA0/MoASKJ0nIdR53HIob/LEDKm/rcqzM
/cKbU7K8lr25Ax4QKJVbIviFzf1qS55t6FsDnvog3q55mhyvWhNV+1juHm2ocXQt
p41P9rM7xdiMM6qnutilbqqMWuAFSJEX+iFae1A8WkVapIM7hFOliPq4PuRZn1Ne
GlIXbkhTn142nEJuTbqn+6SU2P3GY4ZyDWb0qFT3AE+Gfp6T1MNz63nBSIzstPAw
5hTS1XQlEDfQ71DhzXwckijDgiX9MU0v8QStL5Qbdret+oRGyLcktSd38Ue/jyI2
MfiGuWopKvXxGmh8xvbLqW3OlV5b/klsnIdlH50mEEvMa+9C8ukiS8g1V9YD9j5k
d2Cvk5oAFCjit/rxuT0EFyS1vLmHc2lE2ifsVlmwt9g6dIA1wRBt3FLOdTS5uWhY
8U11KkkkQMXROGp8VsXNgjyg3QNingesmD9HavaShtXUVx4UlMbS2oN/F0euccnJ
1u54F6CQ1DH+q4jfDuOhP3Kg1Q2xcHLtC9tBRNshdRFIheE7fbkXrXQvSsHx0FGL
liF7Yl1oBK9RIO627Y0DRx9GR/NH+ug5MdIXIOeSODwUPmiUK3fKxvkVKLvittO8
A6ir/ccug0aRUGCwok4Qv3wQHgW6dRyzX7BIL4cjI6C+jOMhNoHgZr1hIMpDVBxH
s163QyG+z/H08RYneisJlKZbuFa2Opxbhj5JW0RAWhcGW6XCFFIahOw4aORcJTOD
tsoAFZf5mVNkYZaqvb39p4hLsptb6AFbJz0XE/XqdAnsH2hIkD/nWyga+T9Irhdv
b8raNSsY5dW7/ZRFfTQXeUZnnHAiSzMWpkcJB2SDXSWsxJsIu9nZTcsxWLIz4/3z
2aLy6QcGMoRD/iTK9U4jBSnVYxUL12oFZv3YTK9HKcx9ToZVfjoGxRoG/AlaHeZm
q1fWrglT0dRyzxLQE/xiDCNv2irzOb4x5/vC20KotJ6NEWaYkpGA+PAOpIdPd2z0
8/+llgS6f9dCr9asVojz69EZt9Z6yEwkiA09FgEDOHo93hbgaG5ILtws8RqAIQDP
wCaRM/ODsN3xtcJruSo7HYaUL/qUEIeEZJMxMI1M/evz9yJphCHOkp4X0SQPluGC
RLf2Gpiw6SweIXF/9dM1sEUDFU/bG7Cef4G68GVqJFJzb+ykauI2FnHcqwsKDC93
67pgY7I/1F/tF2ZmqT9l4iUY3dfO/ZtY+9csG6YYMnNR6vQo64sSuc15ctRr/YVW
pGHD3zUVhLETGup3jmvWMr1X6ZyP/qJ6UzfmKuR7SGiR8n6HWLyA9+Gai6GovWMC
T5N+b4h2hK5j8b+sUv1mj5xewmI5U/yj2A0yZuAdiMyu+qjQRaU/Xowh/Kd1gThq
IyBYLFI2DnnrIeu11prHqO+KkmlXqd73s3Cy+wcP6ze3SY0JMtQEkRvquNCQZT5t
k3sSIdxQRuqZoIqeDrlO3ahHJU8ueAw0ntJXiN1FZFFOVn0ydwX88L+dC2/jvzUM
LkIJvT+OkBUCtQsUZ46GAfOMjGrBoFVs4GcV/URhhzS51MNisIeRV4RieCZtua1w
tuFEbTopruqdw4Z3lTvDQffduM47tyfKm02+NF2Pm3FEowFmR+DxlKAVDYDh18WY
DJCXt+qI4QMk7ZUN7pIzpanZd7YRr83uzW0yzA063wBP9gaJacykw5ypfxCKfPDH
1SaRNVmlSJW9QNy0Eyum0qvS0rWLCDEv2Nb4w1j9fY94CofPxSwHHfxeLIrl6OHW
jymlyJ3Yw9ipDqjQWcDycc2yBV4fzgG1DIUeWKKPRVvrruUg3D18WtsiJ2BZi7nB
Wq3k9m51hIZRGPCN/YT8jpcX8KWsnlSq5QBW7vPu53rmwZJ9CjuUx3RSzt2+aubq
KpS9nSandOjJEKu33KFCgOnGIyLcWSW9w+krZvHptOTFK1ivir3o40fenQ1OefMt
XcMECu/z1Z5WTTSDt+2dahMLfLPlGzkkw+92pRDqPW+3QE8fmIQfCt0OyXz34fW1
KwotErmc7jAzN5bGCOatrgwyVfm2ZHO6pSIvCfRdfUZnI4s2Vmx36qNAbW/Tq3kW
acdLiW3Df4xoydEgiswf657Ldr3JwPsJp8zsug+1IfiXpnzXzqT7Z8tJbNp2qLYs
pIipBW3FhcA1GDhQmtD3BCeuTJ9/NTZywQtR4cFdvxISlro/LndpadmRt8T53qPn
uxIWziWDxn8MQwa+st0+psVz+FFG9VMtCX4jAgBoQwNN6nJneAoWVmvMVaL81ROx
Si27Aqs1UjscGQiOs4yJDg2kZTEKvQgwx/hcSkb1o6/vTk3Q+jrKezMUAvmFJru3
4aUVkVTi4sZULQ7B3JQK98UIrBjkLAMpIiIe98m2zU8jprabGV0Rbr/C7StazLlk
CayHDGCtEYsKPOoJOAB3NEc8ODmPwJpcry7CfiD7oze8ysiUY5gWEJIhSj+D1s7c
aZPdD6JFUykSj4WS+DuTTG1b7FnTbEzrr58LySRjcqhOjpHahshDAbDX6cVCIjTh
wA78GSaqN66dv7slATO4bNiKW1gVB1lkuatjicQbx4JUKxSawZD9vE5y29IF5YnL
t5Wy716J7g/Ve3GjfUCS8cHg4xdj51k4qHhuBsGB9DR+HWQVAAv5nb2lWDTJG7KU
w4C8wfZIPO6K1JLnCGIxMzKNXNx3mPd7Y/bCcJ2VfuT0rKzkTzAFQP76WPSSmH6z
BEgIJ/5QAfgbTGrCLce9/gAKv1GeMri8+zbO5/nhbxveOkQ8MWYaamDi7D2pZTfP
euaHIDesuWNaQk+2HQBveE2jqSJ0fNVEk4XvbHa43+LUSusrTws/qGiZH1BpNaOZ
0kGgvN7QXezQTFqRQSBi4GYuH5Mh+G25m285/fYXgvhm1SdrQmUrpysXiRvatTiP
L/iEas+3BESNyzFN2ebqhHvXdpcA0Jo7mdNQPibHPKitrKQ67G4crqv+GeXznVn+
9yPVWiU9nYX6fWe9Iqq8EUVrq90TGaLlEOfAT6NTcOszJS+zmZW5iX+7t27ghFHh
AhpXQvuNRdDYUVE0akkiJymx4bfvbS8FoTD3F2r9EOt94hnOOTTZ+gJQ7GT9fZHp
HKlzuCSewt5hhNDr4diYg3OvO+fnTEY+su2+gEK0J1xu+zEj8MZ/qy06mZOQ/4Mp
lwTba82UYpNO/RLBcmQKnbY47eD2Mpm829+93zLXEnxUhfB2yVAr9+uY5KQ2rhYi
dfQCFWALH+u/9UsDX2PpCK57VCdEL7Fbn0FPUICyOdZqYWYqbLoRDRq+Cymri4vI
qCj6WeC+kdCiqoqCm7/E6yKnq6LroOtO9kwJe5fOyZJQx/VRE9mwOnZbuUuMwS+O
i7991Qf6esa1xngRNdQqiXGuNhGjwjo1yG95BwjbcQFZoxNWSkUm59mi/67UkZ66
j9BDqmiXVWCYuzMUigW6GTZ1uPVLxV/fZkD+b8zTZrsUcp8UZO4gt38Y8O2mdJie
GmOslzP2JORb/7pJ0blESssLmVrQADf48rVL3pIPPnDvYOEVOlxRsIqrCoKnTY/V
zVUtP2paVx5dYoqr96ucQiEZEKnh6LLKa5kw2CT+rSjLDB6ofQXhDMER87aTiIM0
8NfnMpYgsphlSTuV1oZbs1BbatQzieFb5g30XA+sYzWefjzPH9PcreN0OmgeVhBr
817WvrUbF3fipx6ntop0br33f4iBBbrTv3vcZZ8asLfbQwYIDyvrDtzJudfnS0GE
O6LWmka0p5dHAJQ5XMQ+3MTMU+oCFlZ8TGeS88lVkOSPR7R7SJBz6CWH4q4JaY+U
dkJfuIZWc/WMIkv/dbfcSXa7QEnTmEgQphIGiCED52++iSMvM1G+58MyulklKVdU
S1ZfaT4dqnQWOh4DeGxqifEqfhS8GEzpFICnh9wxCbMthPFGVYvMJ8L19cfT1PkT
O4ngYCwWmMwcqfwF+nZo6LzvB5bgMp9Ked5yoTbpP4DHccYXYdBRQ2BKrsfvstVC
JHXJ2xz+lYDvmZ0u+EtR+/qIZXCZQPAuBs0cU59WwAUUVkaJL1SKM5SGz0JPYYKR
U6eAs/AErwlUaZHnN+fBxj1lPELSJd9LhDMaMPp87mNxL+moZo5GZK08cquiaJC+
B3DVq5c/P0rmgu7y8/fLCHDUJb5vJTncc1qLDP+C2bV0rSuphS7WICBqgHMxf1Xk
nuQL2O9nro0mHrWVFtQHumzM7uSaETNGFOtM6GZs1apG74qym6cfyGQ7GuMvAQhq
W/UocpoujhYrvJ12/w9zl942MwvN+kMiTUGvgBirHl/WWInGsoepKR0uGYFCRo+x
V6w/ngcArPTH4hLnq/oB6yWyzvSjF/WjKc/TnQl4wlRmC/qvGzCC/cg69XUi515m
a1Eg+jpFnx+za2ovDdJd4aykL9uI6HW+UzwE3z03AVIW9Aydh/4Nld5P0qBA5J0K
jEcrjyI0WnChHWhwBKpYZG3dJkjKitCewTj3szA3dhWtcdpksMg1TY32j/CX8I3/
gnchY+oz7saVS6CG2N1P/Qfq20cE5xuwWJxoyu0bV4w9argf4Ai1ia+t/eSr57yE
CDozuUqBQHxD5LJLiQA7w2kIzy7+HNQfmvfb7wTTwksg/arcJiz7gJzIMrs9Z/Wj
hgdnLyMsjHbvayJ/jBnJqmBHU6TCSFxhjGKO4M7FjC2LyODDEy2O6yfOBV7kczAf
q8ZzfBbbIbB3G6VD4YaMPv49+/KfoCjDLs5tce6IHqFf/W5uElWYX5uNiiFwWyfG
5YJ5xDTa2ww6iSv6db/pnWJZz0IB8F28fbPvvI6nktqgVeZsIk/VVyt0sTZB+ZlK
t0SomNSGE/ZPFJ/EJSrLhIVEcdkQtYvpGAy85H7mCSHvJMK0DBBpZJ6JY7VS+FR+
6cMVfJ76DsDpQVLwSHK0ougOeh2mT6z/7qz2vtOu0rGP4YMT2OcjUJaQw1dotuAP
Yc6qiCceItmefX+OvgMoqo0Oc5iCtpwct/iN8iDuw2YCFHWDUsltVP31YcK62Mcm
uI4P+5XpS9SkYcb8JOQbBl1sIKd6ZLM6wwGGjiEXMUDAt2rKh2AyIsYYlJjoYWuf
/uzCHUpt/GE5DWy7QfKPtZ6XSoiTRWTEoTJpQaVvoZumKONV5NMQfW6DFYVm6tbK
5JQL/R0lCdDoReEyerpHK7798zBaGUK37+fJijt5q+YCBzApA74+Qgjtbio229UH
XTQ94u6ju1rDJl2gBJY7PxeYnQFCYoy1cQSgL3e+ayMWmcmcC4Njm0SUEFYSEQOv
XyekSNTDuvrR/v3pJpXxCA0Dy0oPPN/67n6DQmLHi0QTQETL2sEwYhA6pKvnWMS6
uWg7r6z3kvawBmtlS4018o8xGkfcuSq8s5hhuxI54NwlDEsL0ePCmUEk8wXDvvvA
6GQw+fycCvAGGbLF700aKTah+JQpZ+TEOsyvzyzgNz+bZ5xlgqibQK+1KoegCduc
lxwfMarwzXDQ8f+I8HZxk2K7I2fp8O9FeP0diEZJRxVFaJ7CPNB9xBK3WlSkLGoR
tGbyxRoc8GayciaWczyfeGmLYSjSrwSGVCIMs6DvNV7+hvSjFBOQTMamwnmBooCh
Kk6FzMx+Dlp2ylCPDoS3Mirw2hYtTX53oy10/2YX1uN2ZQwuT8/nabPnrcEKvW6b
3/jXhHt6cq9Uetg7/tYcDdfmQOfSytQ9Lwd5IdhgeFXdfpg6NoqmH06bbSWV9llw
jW2HyOxUNJV3tbAvY0QiG70DQhceZWkkH1Zefpx19t1xHgx7pEBfKyaUs085BscH
UuR6Nt6IIlmFwT5UqFTIyk6GinVP+FGTRT8UIPxlRv2nf2o4oSH9nUupXScfwP3K
CGtrAFNj/UGGScfm98Tah53tVKjDfyxFM7CwvgVlr0sMn3J6XJKWiBqOtm4cy+FR
EZcjIeloHJAxWg/Rh4n/fW5phZ8BuRRp1EDLm/jsgTFCwAdL2iY8hGWEaQBwqt/0
+T7RqjKKc4mTuqnw0WRSzmlH7AApS3kgENcwrn/+0tj25VENIHJkAqXOsZrvnNBq
zCgF1qtz7ftFEx///IUFZwCueHbg/erbu9AvLUeRmb6rnOjwWZvi5UPzdIDJ7Pyy
+ZRN1qCRBIpA7Cv8oiUsk8DQ2oldJgDlz0LrVUihq4cuyBxv64DSNiAFWVukRDBQ
nq2mJDsUyuOJ7EtHrFo5x6z7vlLrtUmREGdov+u2pyG+zarVHvUJ4VteC1RwAAud
eMn4wfVdKlLS8MN9OpDy4A/BQhl0ZF3LAkRuQOnWE4NcK3jjlHo5DV6ScF65r+ha
czcvSCEfS101ctzOAguATb/quV+RfjQfUnJEu331sEJkRKkNA0FjpqRqR4OqqWzf
q64Uj/03x/tzOsM39EaqwS8gCpbKyN8luyQBL3GzCVWWNAu0Dd/IU+UI6NDexkQz
hVRyowGbb3mCFKgnfMq3u2GisIU8gdmODwv6fVO3jrXNt6Zkn0sb/eg4LkQUg2Di
GCgXiB/LNVV9mCd63NNEUmcGMBKuy769sth4GKMJbyF4q4viGBz2BwX4VLjsWnE4
gAnHf5a2ElFtk5jlRxYXqjM7CwM4Ch3sQeITasJJ16lm3Vvroc855iF4vM47KOM6
/LwBZJUVbfmEGdVrUwbtEWqyvZAauvHskEkbxiMzf4QowaDxF2q0xAbsQHgnrMKh
gKxr5v8XavHgSZnksxtuI+RDGod80YGSLt8rSzCm4E+yCo1qJhuRSe/7pzgdzZ1e
t6RvcVJs666yMOgOjb0ou1p/zuMK4JkhGFdfD8XKSUHMJ35g6f3IYDZO88jpn3Eh
dWFpuI9aHR/FEun7XYPpU+RFfX9GNM4HBowgHOcOSlpWhVrINfHkz4vcDA+WwoSd
Q4Mq+tCQR4tU1NMx+GSRejCyYZpb+l3/umWt/CzIbvaXESPgvx2vDXKJNjJ7W/NR
PUPhwirkRqgLplOwvDaoLMdwAhGf8BUJ9hcDtBHlYXmlDsWVD9eY4Ih1cq1AWEZl
Dr6SqMpvDRZKSBm0Nwg12Yd9FR3/1ADjZgUYx/++CNnE+P8K+lD5G9/i8eGu+95A
rdH1aPyJ6icLomXlCPQINnS1Ny0f6Vxo6E73D686Eh0BKXz60Z1cHM2auHbKpAlS
2G6DJSbl3qcIm86j2u3xwuHRqouZN0D3M2LT/mDIte4plElqKHcp9DJuxmMwAI0c
3B1azAcDiTcmnmQxeXDohp1iKLRui61dmrHEKoG7Q/n9L0VXgUaMCKGVijHIeqwV
24EWuF35XP9Zwetohg5jz9NpFrnFwzS1zc63RRCRRfPHldehtL7H7ra5/wOBKgWu
+A98UA7s3qeFcO8CsWij52TXxW9mQgm64uGUSEKR3OXV4YIrw7qfErfTpyb1nYVz
f5OzUJyqS2rYwaUzNpLPKebNBCCCI6S5F/i4rRz4drEfsYzHxBvBIycDmkJr21+3
JNP0dYJgK08jywonb4VNVxBJtK3zUjqd+j+kuvCuhChRsh9xwSh9Un7fwNzHFKUM
atjB96Zgl8GcNUBpPmy54c4MOCJLemfHiB8FFv8HAiDfePrxfvfo8AKMTBhyzvqc
AnysE3p7i2Uh35AkCKvH2xT5gY++IwZGb5iG/dAip2g6tqZTKOR84ku7VsDO4R69
7o923gkuwkfS5CYrP8LzpPo8v4eIMVCFd6DeXpONElXTXFchfY7ZhlNCHBKw3fV+
zBiopu2OZW8x7MFP8Cko6VdRd0amxYjsyZnoeQ5Z84+vInLwSWpRVN+iEN4Dxgek
m7vVxlt+Qm8xH/SAwk/I5kKOBb7qL+weBYLjHSDstkOIr2muUy6HB3stIC85jLWY
wdxOWa27na6Dlqz260n95Zxm0CcJjEnEDCIKAzDCOUAZfvzrQ0fklBae29w47TX1
Ug2/1HZ2Nf9QeYCKQBgK9u5AfEh7mE085BLAiBj/tPWTE3Cqgj4aHzdv7YewrV1l
r5613AgoX8j4nPGwFS1CTfY6F486BgoR1Pi8rzkrQWK3fSn4Yy7rrU6rtBR6Wv7j
RoJExOltnY/2Sv4VKxcA4Pz1f71MvDkzdGN41jn2lDtJGF1mJCBGVN2YjgQzX9so
k/ljTkAjqfa+o5C20H8Z8rNmyDpHG/0koWKfcjZxLeumEHXDG72Dgn0bZiysx8gf
B1LoQ7wya8i6JCsqLf1jcXjGXoIcu4CQqvj8wEs3FldUWK6DZWlJmGlQf12Dq3nb
hDhM970YaL/91OKFsPHluXgIuRnblOrUMCOJKiCjxJstnhkcMMxeyWeAMVcWxFiT
MVlxs/wSyse+EQkPxdaNAcQoA2DEptxuzAkA3J18vW3gFXeIrJCeZJ45NEQ/Xf6R
LPhYFgiYTihmvEGg1VgqxLtKFjLWEjJxn/fRZPseEhsAd4Cjpiv4cHNFfoFcEX8q
ydupwEBdZIs8pivXQ42F6+Vrj6PERKkn0J+ZZC0IRnZbDSVC24cVLMIEZzNBXVN3
Y8KJFLqacdFtNZH9AgUUZ1XJIYO03FKVNBl6+9FUGJURiqdL2uCu2B4ebascwUK6
jo1zg3N34VH3PwLRqrSexbh/OLTPUTex/j+AqzL1K+7cHdx4OnQVREPmP2gfYQTZ
HdliSC0btT5TfjB19HefwmPsYewdiPoNpZbyXcNurkaNmm0Vj4UsWaU7CBbmkqGW
nh/xsQOs4zuNqyQN/uRkHRIR1xWW7g2opOWgm7wJlouYlcSMnKmr9aVcWLeDrbRs
GKomBF0+NlvG+zHls6SQ3PorpvpeXONA3bOt84S8W+vfGVHI87bgtgtIW59j/6j5
IskZkc0tlHFEaLkfOd8GfMZnlfS1EY03AJr74qaxIIoV6W9WzuaHLyoOecgV2vf+
FiI8if2oRjUuy8zwJFJMp+woycSwfKion1dHg4Epx11YGXtCab2AJ4vZedl5sx9y
gpK5XLEd7A4gkdCofkIv8ujBRB9ria6T8A6Ddqf+aILG4cDT7IGHTQnX9AcV6S1I
U/7mOd1RyoSfaNfNPholOGl2J7zVH/yvoERHUiKHs3qAvaGpS7hn4ApVrgIBahBY
yOzQxUjpIbGvxiJ1pdzKx4bcNenmiMxI0csHb9Y5c5DTAcb2T20Q+ZTXltDXHJw+
4MP2Wc7fTFP/P9c/VjNMANPZdo7vAzTvOPfZkn5Ek8vh6Xa8pJ2FZrAYMkpAdSRE
nEEmilOs8WZpG+0THkPAS0GPrusqCFuUEExKWQdMgKsdS3/kQAKQ0dpFzynevbw/
LeMcimDrAPvDuFiSD6KkZ3xc97VyNJYeZcV7UB1+IzSEDXpPAwGgjhutMi4mRNuv
pJ6zkIwQIBZiJiejBpWVk5uD/l1odoM2oeHYZh6S5A7yLAmHeQwA67IuQw+iH8/o
r3IhPLNfDrMRIrmmOaaooTqPWx6zb2gBpVRMNZrX1eM35G7uxMpjbm2pphDYYa4Z
uZKNse2BA1Y0ObnHZs4pcG1FgFvhtmwKyl0MOi3qvtfIj4kVYSgUI1FOpSh142iH
4q9JeQiFKC7Jw9I/4R6qaS/dK/tPNQhhu8+co+Ud3DZ3QTyPrcfMmZ8JfV1HP4dM
MMrSLhT4sGqy4C5njdGYXO0izD/uB3mvM4CoFFpxuxQtr8PRKX92A1Hp4ZBc4COo
dE/5++DWz/P3WJ4duFvnYg0qEMktj3HXvNWdPK/38kn2jphZzTgZuPLk7SjZm8Nb
Ps/wltT+k3+xhIcEL0zGqq3b1WRMnn7Qj0zLrNtuIp3BX/3gaPtaB3NSuA08ZRiW
UgIw89UeapPM9DO+0lYSMsbOTaIWAOm2M8pCC9Ce808iJmBict4YllsxKsqNGFPP
XrFYQ9MZ1QkJWJ+vsp5u8WogmD1bZFNrWJkymclbIcVCpD0SpDMP97moi63pgB8e
O2xr65CITbOH0nkZ5gEJ5TZIUGK1RZaCVDP2tB52dHczkec77ufIurCakupOPtxL
PK+a6IZI8NWiipksDPZsvkkHIMVbxUFE9RUzJG9ylmgPdzJ7a4wNN2/HT0OhpvQR
RfmCgkNEC4I2vvi0mx6xOF5OpnJtn1o5sQIANmzPdH3keRFehA5qoqp9CHuFetDR
L/EvTqdbNHcCxPqmn1X6X9NCDbCkAAYLYTP9hRT/+1QY0KpGUn9xhwnVvE7sYnkh
PUpDaWYpjChspTT8oWTp2hf5K/eDxQoC+sohB8YMwoaQzohm1CetyI5an1Zg7ZZ+
5cO82CZiDqXuHRfIQkNxS4wnOV5Qp1Rsn03zNcgn5ir5lxIY2coxG1AjxPxdmPUL
stzIfOQzYY6pbw3Pw5cq9JkMGaVFamZahU0Oc07cotff0vrVV9/HBLCkPhRmGZe/
zSUpvAOVFvlrvWQj6Q6WD/ujaTUpE6gikaQr260IYS3CopFnLeMFsRA/5GfJMt7k
rZQST9z8fdK5FQl9iAynUaOaugPGEwEc8+vd9qtmV7gHqnUgrneVQNPHY38C6vR/
GhQPSXnodfSZR29YXfa2Fb/+B1uJSRDO4nl0JD1RG1NlMyciO5l5XJ7WEse/BSWW
4TdD+Uu9HWMuD/nQsppP88ZyEWfY01IIgKn+Zcoh3I9V2ahUUu6/hs80k5fYpNQ7
9JaLgFnrn89z+DEoTJexkkuGhrCYXeLnv0/5wdddeVQN8sPe1VSxC8jBIt6qBEX6
tpDVgPYDNAer7B7y1VHilrfi4VPY6y4Ku1XZRibOX79UZ7in5q5CabuhZ10x0qth
WBWTebDOXHXZXVtG1lalpfllLC2apcISiow/dWCUaz9exUul0X6ZaIpG9sDqc1Lj
AKPdQPb2KapBvOOhKoiyr15R0WpAeL5w5bEX+cwTGfdqbtT7+jy5TL7ORbuMrk2K
gjwUq0hFboSqF1N3RqbvKURztMpzDcGSX92gdnnCKXv7Tpl18CaWWfjYN/AFe9Wu
WZH2xjfb4WExQBtS/Yb2LUMlsA3iNHoLHi65ulTZtIB9yrfeAas7B3/TJ6iF5Hhw
TJ/JbrSGxP1n0ZILviL+tNmO5fvvkPh2UXD46L1JTg/LU1Tnwbg8AmGzmTfrhUGs
k01HDSEN4Z3i4MO+zk3O1LNBMyjXpT61vnZxibNXzm++sud3WX7Lbk42Gz24PcJO
lEfIoQqSjbykiAF6Cdvg0dV7wwBG+Q7yuvGhjjwZf39myMNbnxXIyut6NBbuWj2t
Oe4qS7wvW+kvBhnAOEAtM6ZAi1N6nJlX2tEgh8vp8AKPWaRlRb+OyyORR+TcFMvt
jugG154moqyCDlVz+h63xUL+RERugGYL9vvN0RIb6cBWqk2kn6db3ozyTOOb5Q4N
0XwhVsmHyX7yg9UMetrihPBbseHJlPvxBfBGDOM4ENGTSUZ799BxBraMn5E+8Y/A
KMU7e87vA0oA36+p4lQ2foNRCRp52mPBTwFaEY9NzstyLnMHSHoHM51/wGdtRgiN
kvT+tLsaw7+qXmzp7bXy5EFGTKu8siCOgUVMuKn/Cpjf5//LwbrYGIYRU0kQ2Om9
b3a/fm7auCPWoCcZ4YBI4LzE5wKgpkPG+C4sMXpvVlSGZ+tTpC9Vco3Tk/KM1M0M
SJ0YyKfdeLDMZVswuiAUkPZk8uTQeZtq6oxVAWS/6j3IfLdQIqIXiO/X3ybgMyG3
YFso5LgRhF+s8ChZ3Ycc8+sQ57bpKvFYa2P5XSqdmXio1AmrgLUsPZM1vOysGdAl
LbCnA5vfJltloe6W/+z3u9fJLPMoeMsF/uYuVqt6alOCCzLN9/8ZmIaQ85wXlvJ+
Tx7ac4XVGTEriWFKXn76C9vBxCUnBT7i2COL3x8EJAnZW2obCty39gWtrNECNfVM
bk0QKOr2Zb1m9zKaQfLUOp3kQqNL1vrtJk3B/KsGRZC2QE1MXlQPMWGf4SPUS3/b
MY1lP6JDUPyDd9J8iRHnJT2Q6ppL0f7b907E+ZGqONYlIuFpyOKfSAdz9fxr2a7J
a8AgPkGtAd0XBiaACScIyOE0E6z7OurGt5XUQOv3Cr8gjQAFtlV2QpyljZTaTs3H
DInZu/qqEvuIzQQnTNjxp7xEGksgpoRFtqtbwi4nlig1kdW6c1PU5uQ2dunwzay8
aRnKLlajf5r0Ru58MffVr+q0XYhwmATJz9s8exfIkXULVfA0a8SAEZByfB05woiP
NgrqAl/hnTHQCyVeHCur2Gmef2xa2xoOwLrpVMcVA9bU3kpQ+oE6ZdJqjVHnZYTm
L8Hpewz/GW98/ucALz/UZO1lvyy4Qof+lUEpE6b70ZG7h84jt9RROwLhkFomnKpA
FJLq6TBgfpZeD/xZkOwU6iWC3c6hCszwBvJx+nxNCrlTN2VYX9bIIXYzeflPujFa
g95DYeAkx2+6+umf6W6RWde09vzZf3MOf+KWzu0FuU/BgxMUDZ8Yujjp79rWY09J
4RikHKRrRdLPVzlfR1hwDhcNN3d99I07PWmJpXhkm6rlL9JmDaJ9zRQsTGu+v9Mu
XR7Fs3lv7kwcHQjymPiCsN4YbpjzH74gWpHB/UoMTVfWdMVV1nwEFwwaOLWJddZN
bEIhe2WLBHJFxWL92Yy5iLPS1q1LtVVjxg1OZIzwu7k99AdgjZ7jvX1EC0BSMJDK
OYnM0ehKxiqUbXs7GAtTbKN9KrcQVK+Xy6KbHcue09WMNpjfZd8l8xlSY2jRd44M
n0NObqgbzCTa/m/ggioCrq5y8TRXW+X7Pr2m8dOsQNc3olKNcMQNuDdA+ZxCWbQZ
MuqXAyuoO8F7QsJjQOw3RLJ3qrwc5bgWuOiGKyxw4+1PqyT5+Y6BRWubXPV6ZLJY
oI/9FEEweRDuxQ8G/KBQ4c0CxzDVYo7if06oTFtqZxYEjHBTTMNhwz5Cw1GBsS3e
8RsjR7gWHkOpAuvnnkeR6zZlAhfTwkVcLF0PAF5HDBTOr6kH9CTwfqxQfH4WvcNi
mNS3cRt+/ZzLSJ5X7qSTBjr1zFAdq5pAc9mRzY8BYof2tob9eWqyccs5TwN/SNaR
H5CZ9IgdOTVCw4T9ladjIaUrC/HpQx82/qGOQx8JqRA5h4xPLFH3YvwSYLC6TTwi
F2v3b+hC5nbT3gO8L7kZBnFSkwD7hB31ulFjuc0nh+DGVGMIMuodgSXmnZFpPJAM
bFVZtla3JPvA+/YeJtFH2xkR4xgCw9BnSFudl4jT0fKC0kuUddw1c1MIU0VYt3xo
+uC4P76qyiQKDa+xcbO2oTHObS+jDjAN7xukgUBeDpGQ4/xnypyZSZfGVnQ8T8we
ClRQnzuEBBtmskt9yUna3GWFoDQtQ+sUk5w0SWxnPQ6Rj1nHsMy7FvGr4HzGZfUo
ha4vy6VnKbuJurRnchGEUvxKCWg9//6/VacNidj67LQmtBs564ehDytOS+qBG8S2
ElFx4rVEyly4IGRva4+mG5kDvAReH6zRqM080N9J8pZ4kHyxVLmCARVYfhcFfQ+4
a8EMJhaS3rv+UtPDOTDjI0U1GTdgN52GijR1wAhGVwpCKFOInctfYixHzSdf+Pzl
XbeykjXmGZKD8jVEMaDY+xJiURF40Z64Qy37V9NbzLgzmdx4IwG7yjWMdOavf6TP
nt7KKDJ5vEwhxtuEUJVXlmNIMPhaE4rW4hTbl3oANO8WlKUeqsMAq3fUJjYtXWu+
zD+srhmuvDNfPWBateOS00+fCyy5nbksFeL81piIWR8aEkFKwSi8rU3mA2qqlqUJ
YchHD5l1uYvpMOR2xvKA13TdEzbFPBZorIhQ9CDQxJO8T/omQFw1MygE6X60M0bP
P9NteTkI5oPwCjhDMD92tyLQf523Frfu+1nybhjxMo4JeVcYecMgRfz6uCYBiw97
Cz+YBGuZrE2cMWrGIPesflt+cYQM+5mCiCZytg7+5HgkXJ6B2nQoDA5oG0Ku+hWD
8fACkqYO7Lg7m54pz7Zh9AvPlAG5vWUYaxjvNYaJJu6Xw6NJ8pU2cZdn65+kgt6m
7ndrLqyTUsyH0A/x6jTOwqqGoNv3FX8YQM7yLGSZs0GwE+x+xvHHZCzx8alSfLRV
sarQlLDRsEULPsIHBf/HZqNhqTL/vfK66sBA17J7CzgnBFBdSKavH6dENgjp1WJi
FtDxThoWzVj4sldKltVsIDgpmPC/XB2dSPywW/YEd+5q71kKdbGNE29aLSffm8lc
ZD9KD8LZIG0XEJo5I5nGzyiTs5qcDMrZ8wfQZ7vAcRF1p+dWEt29j9ZrZcyrIb5X
m5kAYU0mtpr+H/MJmT1P6ZJWE5SGTmBmimTGUa+cgUXq67yGOFPRbx/asY+MGk5N
jmQXB/tnuSfAEd+T0tJf2CPXx1MfupGugm58R39OrpKNOZWzAjWH0yoBsUySG55X
aE0iBdbnKgX6aGeZHP5Pl4q6M5KY6O3bKhO5uj9JDxA8onkuJppbUDaMKXW7Jubz
ACRT2knd4toWCWFKzUkYGGgHactinexFh09iCJtwQFHn+92zzW+buPRotUxoYuh3
Q8NQcil1wkztDDRyZwE+ZHqhqyqqd6tuyvnkaykbGvrAeyYtiZx89cIkirYQervc
pIC0rMqrFYmIVUL3pF8T4o7Nn+pLdo8gNTzh1cSvcQxwLTVFa8hr/FvCJjVlk+Ub
v1/NoYfsrjrJQUF/feAlaTzUEYQhW8Ref/XeGD1bWKleMP6rW5sbmIyjnoSlfmN0
PZx28gVEN+AQuAETggWIQtgbj+QRVrCvUTTk494lKTjn+xWOIcDAuBBU5jWtLuT1
CVEE1hXbXJM26STRUvsywpXIvZfUw/qFVdVWJHQsDdz2Oft/VCkpgJMI5OsmHKXq
WaS5i5rKixgE0CFhJF/ppluKlkdFxaxajkik/i1u/QlPgIDCfIFIVguO1vnEmBHa
aC0ecjtMBjVZ4wrBZJwgugewfxari1EOZw5Wzi4pyz7WzNHvGR8fK00rfIEo2LH6
rQaaw0dok4k6T+mswvilOtWhdSoJ5aPCsR966xH43Vmja+hIXRzZauZJ2eoWu7S1
zL+0AMIMnPLXFjfpgH2QYTOQ9LRMivs9s6KmBSVysawRZdOAf5/hqLA/Qlto0sqL
WyDoOkWUOZriiORMuN1I8ThnHP/y7FayvlDjScCzbsVsCjVaRDc82m1aGPOtbL+w
530kC7kiZb8M8FqPrgoWEd5ogbI6reFsFKIjvDXwr/ODKgxcjPVeRattZJoZ/OH0
J/Mq3hbk/Echg2hIxLGydfqwr+z7kkS6sAZJamTxvPWSUpSKu6sGvnOn30ZgtYP6
vc+eEN/9j/kigmspwy6/kxx2CBsOsgqQOWfWEQmMRJnbZQxtfIFDRSj4U45b0Jw7
FLLRfpk3F+nc9aYNJCCOIi9DIUPkuqGFwDCU8oAHXyFrwWboJndRDu5BREiL4PtD
pP8SD4a1+OzjmeJ9764BU6jdLl3XVU6bfPRYteY8N4Qw2bo46a/Cnat1WMa37+Ny
qan06EUH5w7b5U3hj9XHdpUyV6XO1UuDoDlMUYqop2qX1vcyVTixdUCy3SbLFKNq
ACWr2rBkFGhgY+WwdjMcAXiO4KowZKYq4Gwo7qcGr8NZl5wV5pofufvVtO8+7l+Y
MaKzuLcowusvCT1W8CvNtYy1DxvNkHqxIrkLicDmjBlfqdyk9QjPYxlcULGIJ/UH
HkAvM/qkRU5ZKlNWPkRQ6utAPL6pmAybm8eHUNkGfFS2E4L4t2rwjCfQnBC5SLsh
I6as/Hy0LIa9m2MJBdOujMnde1Vr5v5b7k+jCP5ZBZlyFC033gdQ0Km1aw6igJUV
2EHjvwGzzH+pDr0eXJgb6cXC0VnNtwfXhbTuf3+FGcSGmwWxxpQHCb5xL/zpmxSM
VcYfe7S92R+GjOYz9IYB8sZtvxKQsSewq2x1HjRjvq/Dd79681C+EXarkZuBpSDt
k/EpK6m8mevwDw1LMzgssTUY8/rN2m8umnppSON+bHwbC1PqDaj2YeY8p2Z8jIKD
wLlC7DeKL9cbkdB0Ly9Q0vGlQNKdHO0AYzOSLEgyWb9vMAhjH9yIaiMifv/B0zLi
fC+z4WKU1mn2yxqVHWxiuLf5upQEDorqK3UqFOygOYH4SZs3LW2dHUR4z9S9kVdk
D09EVfDDsRQP41xVwZPqpdh5UiLRZb8jEIcYlqakdJLqtIaRx0I9MR8ykDKClqDd
BzSOMP4KQ7P0DTNLV95LJoHZZJIQqGlxxAY6lTKiENQtdJI17QYUpGm3J8a90vFm
xYdPFSdH1V8nRKb9jEpZBXK04yINLXN1V13LnJI0nyarF+KKAZtykc7Ep213v9IQ
6G0Hhj6kB78ZFqGk76NlonYZVBtjmZLXh4eBdmmIYQcpQObmJ1fnzzKH6rEDuhSN
vJT1+fIU6c1FvMTCyz6MAIO4ReDo99VSWFvk9URl7zyrrGz9+I7Ko2megonAl0Zf
aZry0NxrZvSMO3Q0SyDYeTBqYFcYCIBb3cYAViJ4D3ZEBEIkYxoGxMa0/ocL/0Rq
zZusDZpYYWp63MnuJEV0b/uQBbudS5pOrv3D6fUbOyGmJJ9K5e2VLHBzc64Vh5TR
TABAAsoSip7uefVE1HE1/48ioqo9SFiQPcw+eDCWvwCwRkJbEyAyiU8d3tHlvIPt
ezkOEZE97uIz0Nz9br7WOid4lxQLSi2cfLVBQDAPC9cG9yiF7K+9s0vRSE9LAwU5
Dbr2R5TEcJ5nJtROl7kc0X7hvi8S5sVg8e4dBCrnBpyIJz9atqM3x3GSJTCaOqhS
HYlgnBu4EjZZcLO9ruc2d1pt4eiUG09FTt8EBdRzq2MnL9uVOqp7aVfZ2CV1nErH
TyuP8WauXRmd92k+NinpDVl9c7DIW04rh4MpQO+yXLY5QwNrhJEH7ICHrDQMSRKM
2IznUSLtZQVwJqUxYkxNA8HB/usTdO+iJqNDcXKep8cHgN+OY6Gz12Oi3Tv1zXYw
GAj7XsCjj3HvlHuPllWDRb82sJlG1xGhWEPGw68RPfHMt7Z1Smtr5oV6wfYS6rh3
etiLMC0V5Re399gx6f0ZDgzQMfY42pOYs+u4InAM+rqg+6mIhyZKboyRbXCwpZH9
YMN/swO4WHmjO+/oSjbw+3DOFrvXOTnfrUtOKt2InYO3np1f8RZjhhEDku0JdbY6
V5lWDs7OSJvXUHW0sUl65hw9aAiTs+XRj/CioXCKLpMkUDKDEgmCIhEah0yP6SBC
TzftOy5qZl3I3/CZ7e2xnKgQSOJoKduwSAMpJ3dIj02nTjSl2knLic9yjbycJE3t
7BNYVvZZi+1vLbZ274dDu9/bWRBmxvF09aA1Bb6DmY1j8q4SE8CY0zSC6cx+wcfO
1eFFTNgts/n3OO34T9wLDpeCwAKhR7rU5bRs2NgFWrHrlDf9AQQi4bxsn7EjmTvj
/mknuOrTvTzo2eIabAUi5hiWn+oPLMatiFbP+ArWSDz3hZeodfSxvVMaQ0fvnCFw
lTIsJxJDkOt/U9Tzvc9ZCLT7yWYfkbc0FEZOGH+y2oZV/LGFohY03DN9oqnVZ50Y
Hgttm7YNmFwufRwFuJRTdTadfpc4yXCgvc1d9LsQptxC2EbHQoUMg8zB/msLFxgp
r5voCpEsqHypzCowdZWCoWhphi0RSVU00xuVpxTCmvcG+M+IHNN9fJOtRU9pBhmG
sXSNfkFIaGbBhoZLDUw00EjewSreqX/umVUVmRpqH1uOUCfPd/kAQviUb5gRmWnA
nJoCubhoxsRUegzrGECsN6suKV4pzwAuEBpw0rMKvReH72QMXHWs7wMA1zeXves/
gl10ENPXUQUmvoZXjOLuzDQL3sG3F89d/8MdowSHk626fIJlQp1oWqMrep9T5szU
i2ooQVG39f9SDtcg0GrhkyVTaspDx1sri5gx02SluZT/abh0OFFTXAVfPr44b13S
OEmQKAonSNXQnyRpB84eXmKEjs+/sYxShv5haPbK4VOnV1TO61uaUIR//Q4huwOv
7YcKs79MpEibH55UxnMSrSlvgvZ/7ZUi8Z47d+ATUbrmvPzatLaipoahZ9uENItf
JFFKKTAhm8jNNZsUNj3nR6GyHMdWTeUtRMuABnGLkSzqT80gf0LGP9L/A8b6Nf0a
hnBWgVepmefY18mre03F+9uVhVcro22FvwmQpLrULhIBWFMa0xw6xvcvdwu5l3Lv
ctibwqcBqm2jizdqn0HQcPj4pDY0pY6hzBtQwQuoB6iRh9W80elxUInVgb1jhYC6
Q3idxPDlATcPkPZFc+4T9KePnnDU+ytaHshwGgBf2h5udizgbXLWdu3K3Xn1tICs
yWQnPQ261Oz1tipOCTORIsNACv79pNRdgHP8my0zqHHknowNDfn38DMXCtQ5XyXa
mER9RCn+YeYqArbpwSVF2AYj2TnU/OLOM3TZo+dhCKwc3o4bWXp1wNcVmzI9MqQ6
KjSly+KMX0MIvL2AQz2wEK6SpPVkVVf71O69jQyzEE853TS/teBtiUiqIjUD9Zz/
MjxC4OFlOcU3fTeUW5FhmDMlVOZoEEsQs623ZeKUACjISKHZR6su1BeJTq5fo+bg
2Z/pTAMAvN7gn/OXxrc0yvDEiCvsCo5AohRySkqnpV/QH+vFr4iJlLreHndr6i1q
poWbHIp37YQk3z9bCCDYaYIjqksWfAVQwrETZusQVssnIRZe13HTXXx4MME8FDxz
4QjTCIWHDdudcIdSRV2JTH/vQRybdh/cWyizII5MFrVNHeq7NwE+KoSwu0VwybFQ
2jJ/oF2DS9YtRPMB0GYi7ApNzIjf/We288Q2uYhQkE6sXgmM+yGLfyD7xCspZjrw
9bCRrz6HELA21LBHoDPVddEj1wRMK1rLO3wpkIu9nsK/Tmq7UHVCyqbV0Pmw/pw/
Wp0763/NqGmhgDRTJQhml1SMFaHpblCOo20s5QAvxceQTLpAVlGmEt9zpXIZdmrr
N5MGov22Mex/rylum3229olC3YtHH6M2YzWeF5QvFHxYCWL1TuCAZMyijVipd0fq
0TYoMV5pymgxQ4lglvbBDKoZqWwTM4jkEh7r2XnQhk8RUHePIzCaFnN19in5aWL8
5JjsQbxUHlRgQpHBOTjgTW6j9rrJQSrLXM0EHxKSLyaY7X33RzgDu1CONiveIvlt
p6ayOdz/Kc8nCblYlKHzpaOJXAXnuyDKFRJ9SfCoI08e/KrEGFMRYKUS8JzqEibs
oELnGKN5ZzdyWuw0wf8ccXJafZpukLzTGNF7D/EIT/UwUnLSaw5Drx/5ug5P3I7v
5flIWHTcnPPTF+fUvL4nDBKe8R696667lzlCypbnXKHiijj5hPiq/to0iiBoFj7W
7s61KtgwMhwj9DMYz3AkHJjX+PXnNducixB8L8LzgXNnvB7ybfoanDhyHYwDreHq
guaDz9oxomsalABOM7LgNu+WgL1nM+EG9aA6mnZZ1jY6hE7dLAyCkZIOR5luHOCX
iaPBl/jNs5IM5poTN34TJf+SeI+ow6D2eKCE0uv04sDJ2pRADOpDYykPFqtdJHHb
npl3lmdFoBXpHVNaFY6KFjf9rr7cvxxNVr22YP45XnMx46RDZJFca3g1PewMoxH9
eT9w3aJvv+JUoRJPFYx6qUIPp48B6gyI0IKKKgnVpsWzr1SaQht6S/0hTkdASO2t
HZCmkpAde5Pk0njXZK8/VCVUp/BkVEkiUOkESnadXj0MqHv1mf6D0/KaDNhXym0N
9a4r1HNzzUiwpU/dC0w1zup/GAYg3Qmu2eC2a4rJiG/+FfjWZc6xMD5ovbTeXyA+
wLYnO6dhXurmFOVTACW0wY1dez/nv9Cq+vPL6n+N0ijneQEq72jxl1F8qC95zUyK
M+vPnUNJb0POrhSqvv9+5O0FyXXSIB2flQEGShob/0GGp63YZkd+Vb2KiWxLiI8P
sSOkYMhP3b18sKR0cCRY4JN9QzF9zu1OA+hhTadtwsEmKCgXcFl2Z5afbzct54Pg
tIypNl9By2E2Q54fl+tiKuQKAYsWL3MBiLSLKm4j5Wbp/Kc45xRPIBg6szqBveNM
IqulK0Jelwlw2cQBvkTU6NYBbJX387EsRdYSzMtd9TC/XFNqahKxlYqxA2gI8cj7
FGjdLrZUSxGh/dhi0IN5aPDKKlL6xS3JCvwIGKaxQHOfaDO0KQLbcxf6Bh+TEaYV
/AKtggvnqboHNFesc3m1bDhuRGJK/k5LmPK9vMfu6F9VNgBoS8bUqX2CxIWG0WXL
SVH0d3MHKcClnx5V0OnZIoV06QAEBAmSJ6+glFmzNm40QHhM5YuRayGRZ3C7aY9e
e+HFO9Q++moA59+GW3IQhHOGSiDk0qkntq/sY2HTKrE6zB8/UTmGXvZ6Vq4Nzmsb
ekv2ENcIFc0CUTGvMn1+tbdxV13iNgX/8C92xVBm/f/j/froLWymERN+Kj7qEv5V
4navUliKA75cJ4A1lY4nSmCKxQUHUv8xigMEaWhscPTWPxUiULeh9fU8Tk8zwLBZ
L0J7Z2eRqC5kIjljA49323Lrhxg6E/RKYMuDZlPNGpyWFazdgnLv4yOXf9U2Rzin
UDAdkK0k4MKt2Ju/ZmHqJBB1cQMAxTkthtv2O/0wTIAOpJ5LwYpSSk7QX4+Tl41l
CUp6hT62ND75UeopJhJC0m7BByrJpOsI7Cu6HAd1mSNXalHPhvbZMcwXe0+M+1ID
tiUqw2d/gRJkQtn0JoJMpyQlzfocI7h8Agnvh+Uwqd1GdzW0KFSPcpJDwnTMPd7c
8ioeA+o9dIWDuZSB+66o8hbKjqPUh2jXi8A5aFYY48E+aog+JxY9mO4CQICHVlzw
CGYowjqVF1wzGK0eEPonZFJwS+ucApv3wHS7pGR6o6aCKCxZAykVBJtHgm928KUG
Sdh9TRWYtXukzEaRUSrC2yw2ce2wgZ0b6voSPwCj7wY7nDRlEw/6VQ1KlhP3+mhH
qNKxA+vwIW4I+MpE77X+/m9JLm6ydPc3sPMgGpku1hkie7eCn2v9+6NTwng7DoDe
MFswWbycJf1A88qMPEsldcoU8laWJz97ySL6MBuFYuM0v0/c8o+iJ7/wBVi0uHBB
PJXzXzP3nnBDtorydHvun6uFsbJcQhSGZKbAPT7AYzQKDUkYtgg3HNUGyktkFzzJ
MBmgrWiT5eytYZW2GvDSK5iBXty4noiertqyvDqbSxKqxNwRuyzlI0w7L0jwtyFK
ZuKHKI+1nQ1AvlW48cYbUm7xp2fe0KR0hHWtwYAtZrqIPsNPTB/ThJ9R5GI+NHyE
bFrmPgpr35g7kllpwCfPN0PkFEhuu3P3L29npBl4YyH8ar/fwuDRuARSld9v/cDj
/A2pfiLBRUL0/kbF1o4fA1bFArmbA4RMlmnxLPezyTfF23km7Rbd0qzxCYcEtqBE
VvhTk+AoyOT1AezN58Y0qGtHi9zX+pdVkSHFksSVo8ZDTxtw0yVUa+tz6gFbBWb4
EmjFUOY/DTiPMjKyD4OWqexMehXbi1Vw1E1aoPQ10op8WpH0DkZR5yy4wh20o3C/
hG8zYPK9Hg3NitNVPlAbPKRF6AwvkfkuMjfnr/5piwK5IL6VWheTn5AB7Y0pezMi
w+trnvjvuBN1lcBG+ac30qyYo1goHpW+9T5ouyOeKiFslxcllGSp0tTX6xw9QGoF
cwMa1rwCDH3fmN3p8pz+HdD2UzsiMxD7WWSELzrVEDXt7UwmI7dz6ZgnFfp2atv0
rM8VSgHqD/32MMVMePFTyg4tZplxlDWLxlfLmzfCJ5C65vzJjHGgAeqQWvJePfkm
Ndc9uDntNvmfZYL97RREMRgFnlaBumtGfZUF5fJJB72pLysws6lXGm61SDDLw+QD
xLyUViDzXi4PvZjpA428jFR0l5qyRCD6JBOpbuJuP2qk4GN97m/Xc+8Hp0b0EV58
ijNS4uHFXf9MWpCAcLm1mSXKQgptQTUDvrA6P1EBtagR0eCG/4l7MzCRa4UNZ5rK
h96YahwNbXG+ZE901jU/EwTkb+Bl2nWq2rl6bnJQ1vHANd8n2y1XjhU/QOmAwntr
AZtvLwAq+Y8/JUD8+Rfs48bHDpDWVfIZL+mjNZPD7K9GoAdp+TnEejhkBIiEYqLI
dZklORa2XwVY7owAp5CLTKcppZ25YJ9R6sYB19xgY6r4eUHF3vOtFRZF5QP4tglW
Un/FDuR6WVC2k7Oipdv5tlas8WeedJHL2gud6ul/ZUfJ/x/HdxFVxGqJxrQQ9eeJ
+r1Xxp1SaH/izafd9aXmkNxNYVTXjc53Co+iA5aN6c2/IPrx3mzL5WhzVCwDdxmN
qIrwSoy2fwcvAfloZjN1Wzvk6r2noOuGyLXph42ewCQzsAqVGqyzc+ymNZRCIoOZ
rRM96zhL7ofA1xiMkPIY3pPEbMMqKBMhuaShd+8Fa6vfPu2sN+StbR3C76nvHrZD
vyeFYCJsbLVMBYdycxqrq1GsYS3oSt6PD94roVchzJirTrRgitj6jZm83gxa6weV
zOMK/N/rI1q3hykY8EYQHbvAvtf2aXYJuRX/w4wW8STb2OmOMxzOiFLu9Fz+GLuJ
7aQX7f1UwnhttlBntlfidnRFm7gKd+J4MvX5wPmdcfiGPdqQCOO6yE/yBk1pWAo/
JfGiSkuusdrq7PDDRAI4fas9vnWRruSP2TR1LCuEfoxGr4o02u8E1LK/mF34Qnhx
Aw+0ic+JS8L8M9HColHkCUMoj3ot19x3Xl3p8TDSo+ulRCRgjc49mb7wGMMJzfCc
Zi9VJvrpt7GaqrHZvXRIBFyuhoLzX1659r2uxa0woDz9qSifu+dYOk8eBEFpjY2O
rxqM+uH618K+Mz2di51IKQ9XTMiwlN/Mcv9Yo8+2tc5R4N6tV3PiDdAtym5MiIaQ
PBVwWGHUcJ10BK2X+xsDD2MzB/yetFSDidM8+6/LrkX7lU+QNnYMJ6/ao7z8lCrv
W2TnbsnjhCNNYp2w35XzltU1OrVveESVOnxkpiByVNhlMv2WI35cGc2rQ2eukbEd
6X809Bhvyotc0whx4VIwpzdlYnx/58+7kS2Yc6Fy1pG0K07wpE9vd8unEwvyy05A
SkI5N2Ui+kFNGLsgi/heVnYDipYFXCVOpJMZmnVatIQGVMTNUUZEaAJpPQkytGD+
TfpWO9Bh+Yef+mTveBWzv1FxYHzpz/kpcx9qr+PYGNaKjdBNlkDQTNHwda9ZOfa0
HnqTv23cpqVAtNtRLnUNYu6TBxfGTpb/0sp0FhEhm9gkBF+SkEADU0xy5UtctonG
HuMM0aSYeUVxc7sWOXNu4bw0XT7KHngEY5CN0sNIv6fyI71QAkRpxLt90MJ4pEhR
cK9babnbMw9xIULPMgHI06tn7BiIIf8tno1JxCydoaCwfQhe4r60QCvfjhvgBm0w
fgF5TKIA+ZqFD2s8myRrwBW/5lU/E/c/yJrzJsSfJAM5Ub0Bo+hofGbpg1q2gtL8
oyNUV9F8BjdcgxjiWm4+7oJXZfbadjXmtKcCTfpDr6yOEpqgGM7Wgn3G6OmzKecy
ZPHCqQ1pCVPt5ex3xm8IvuLD+p6Bmn+4n2Qm4+63HVd4We32JThWf4Qb98mGBGjd
1no7R9yDZNw6bWuqkTZ2bVx1BRTOvkfttOUKtQEgYbKxaqv4fnpGOEHdYueamQfI
CZ7yUKDoJyYvEPc9pl2DVsyD1bzsXPopCxtvHARDqw7GKv63v5PWQIe5L/Wx98Bo
JOB28n1w9QSgtSB9/lZJB/JCqEHF9RsEsQjOcrGuv4fIUqJ9GZmTg6+nJNJ9FS4w
efR8nsRfsxE+pgp3SpG907wu85vZ8r4sqtUIWLCMZxbDAvn//Zd3zrODNu5F64iP
Cd0gm7zWeT3b8YtiCkyo1kPUDE4i0YxKJRXVbE0rX4CPZgjj13bM6hikpRO4dlaw
cKJzqB1Fu2rPQH+ZUZYlbeDILE37QJfztpwAdASMWAU5fmacL75AE9/0KZUhzrOT
WNa0aQG5HThZowZXFBBbxu5DfUb61MsNYdvrBvEX/Vk88ZNsX1XWZ2h7LJPrcy0o
074EN5qFZSl+up70XPqliPaKedZxZhD+AROvnK6NxjjmpBtGOiw2VWYx6whGf8Lb
BpLnicJFKsSiaKNSJ89LiaceDmpTXtkeBcOlhAS55tFncsUwkIHpKbWRQzENsjPl
SxHxA22pEbW6tcn9fUzN8TF/O8jR38fD7FWdWMYqfXK8h2RgN/6j30fAcppjWKyW
tih9iQMG/Vrqv0u+oTpotfyouPjl5mCLM6l0Q+AUbhTKCVyCYhAWqRP2nkT+TghK
i3EoLzCoa0C1sVCwL3Q6/AijLky7GCUhj+LLsWkd4ISAinDIXCOqkhmYbqNGQ4wV
dG9VOKNQ6Z18u7e4Lr1AfX8Ct+pBw9buVNV9V0sttjEoDxnWR7Z67H1VTpA7+0w3
NGTPrkutYmMe6eo1mfrGQ6zwUdsCiu5HijxAfOTMgqkc57rGgCc7jlNCi7Wz6hLj
aYhvQlB9LAIplmR5cIpu38oXQIUp/bit/KGr/lyLrphHtb2JY7yrWK9LRCpOOSsL
lUdCIqqqg+wZofSmMFXu1jbRKEwDRxGsluyzO+wdriGA8/3hvBuiGfiZVAnF2Ap2
esrWz6KfdwCTGDCQQamXN4K9Za+20mtxJaEYgGWSML5PzjJ0p+xcisqyY6ezU+Nt
Ut1+b4mZ1PhfY8OZLCdNHmWukknC+nPmBlQ8Op1pln3gN6cIxN0qutBq5i97ecYY
nvPZOqKNUYHz661gYkYkkE77OOxaHhdinJr/NE06A3mZ5h7tqn5Uq8/BOhseswfg
j9Z5YmtDF3IGer7bkmxqVK1riyZHwHLgiBzqAy2NsZ9GHKPyId46KQsSAJNiG2aw
0stK8ykqzrVTF/p5Y4wfNYha6dZ1wYuaBq/4plMihhljOu/qOKUxaMeokktHiDnV
rtAjLlhefopiLTuZKR4HfDs3QmbfDUdIIxqrctU1DQz5zZP+y5MfPGfRpwr/MYeC
AbNAEy7vDJiGnOj/YXoO9S/+in3Cn0rRK+QxCmPIfpzIRFDoT3uqjDv1GBpkVF9I
UL6v/yHIMBIQKcMuElhXmQ352oivrL2AXsMVNagRN5E3iuPoAdOj+ReJYBXV2nDc
J7MesblQ2758Ifw2QDiWfDUYx9S4eBeDG68C4F46OwmQP9y6d8OCk1HY3v9w1KXp
UhOZoGGsU+hMlrgqReakQIMdLdHMD2hr+a+7ieJcM719EtGyM2Jx5g910VjYOWR+
xN2GeAu+r8srfxX/yOyEA31MfRt+HkwUd0yxH/ZLKAOUrRhKwd96AafRiUUkmpkZ
nAh7JZy8Uv+rk2unUzjgJOMTbbIKonUajg6ZSk7qKFrdI8Q6I+iaYJfznxFlLVEt
cP6fYaP9x8z8dsFg0kXAg12dPgIjBCFJmDcAcDF3dClizC4h4uC0FcCIZBCckZx7
/9ytDN2/vunv5WiKjQcZ+H8HTPWZONjFkCipm6q+WJ0TvhNZQjK1iVSaLR+9d3k5
7aDbQ9W14INAcN3jsCfO4KpEmysXI4IlTM0ht1DC1vVvt96smeaDzB52DlgDD6mn
44ktF5kVk6az0oOF/EtKzxd0C0O9RnmXlLVr+jNa0f22RzD5x+o5oyuZtqImOtWz
o3iBi/w+yctDrioPoE7YLp8GOMmcgQfpS5E3I7pXqusA/7LibiVSymtFgYe5z0vS
o2pslbQEAIwvp2TFFBxvVu8/yS5hQA2J5SRaJLnQC/DngD86A14Lr6xSrgAx7TIH
qXwJGR+vS/g4EhupC4oDFJOfQO7Uv1//yVBuOL2Dziywd1qRIzJBNAsrjgAYsWvU
YuFk/aqZSiyMkolUdn30S2VR5LRazhpZI2LF4asIYjOH7Wgs6aP26GTgHo1LPHzq
a4sNWzA1XfgnwLDuDuwwEO4YYmrLZxRJ8ZVw3EEii6Zi4bODOd17evtT2WIJ5far
vh7fUAaDIT/23QSdc8G2497j+fY6skLkCmX8+6BAiXENcpUYij+LCejr43HzysOe
6bDf9pl4FGqSUPYZORBPxV7Oi31G+DjRJzXGyB/Y2DhkVHoM4M2YXimwwLMjoSTM
PoQOBfmozdUupY/pMfzCfPYkoGxHhehmKk+O5Ne41xcmmA74/akwt8S5smLnBOiF
RMVofuqhDfGOKwleE1d0bTS66/jbVIXHOdZURBxBrN+8QXwiKS/bn7A/WwTN9mKr
2e9COd89ErmGGVBRdqw7nn1vzcR4mjy7/wT91n97uqaASANujiUJ/yKFJJmJ4Cbw
jzLs5ex4VPw8mkxfF7nJiuKqq/2827H2+Xixv+q0XW2WZqaPQX5aIlUMlhJlnjbZ
NZ6EGgLmS1+WN02iZnIUI9/i3n5y5bqeMElJgb+eXYjzONS2YScSXovDbGcvY+59
LVuGfPU7DkiIub85e5f9eM9AeiJjJAs9PglFlV8mfswr9pXR1UTQBxaqYC7lBL+Q
oSbAyLWti2WskEOtbkm/FwJvJir0YVGNp8LIbKmmBWnNoeuSroksX5YPAtwD6thv
yPwuJi8B7RYaz8FWBVzhLIvawft4gwnnB3fK/R0FIpu/uNgnZHM2F2eoDnx6kqWe
ddzVjF4tHrlt121+GbaBJyKlTZG4A3W9CPoZogPDgHvN2iaJoc4u5ELM2P2B9bBY
Ra69AzglZhSI7iaLL0oC0iRvjcTC2T90lUNfIl/+ixBYnIS0XDlfxMqvcruUhe6r
4U2NV62sNGDGKFx9VDd6rAuOrJcD0W7uTR6ZFfWnLirLJ++KUTk0HpawYUNr+b9R
TLo7+rFiuc4R1lhN1mXCm4xzQNcjMq6brtYHikC0ee7lysfAhtZMoEIV0bx0sK1D
w33qUUp3Ykk3zJZBcQPawFWTKsivOYtml2LM+E5L/6eTKA/fsDhER8wKb4rLw6BA
7kX0EJctuLJGMScdvs3OIhifR3UIxr1KeTdqG5hjUoZNpay+aMYYVkPrFVTuZ7bN
ZREyRvX0QdnTwjf29ut6EgbRSIboc/YeMQgaV6ruoRjDCDb82T3ksLa0Ehzuwsgt
uNUlYVa2Ry25FJi2B6ISZBC8F6nvN2xKkNCt4xQyUbKpVol+ddXghLvv8s5XfeQY
s82CPjB2lyBEjFbDsHpYp2ChJ9u61wF2KkQbW3VbBOAOhWv7F0G6BVsBJObW7n7a
tw2U4lurmBWSzLFlNslQ95Oo9WK7dXGbqoeIN49RS1I19YdtS6Byg8KoKKTLRBKt
GBSTs8ExKDCiO4U56zbxjHGB+vzzzlEMII6qTVHwT0LDE9rGqzO6xiQh8OJ6+MXs
JtDtsLnZrwz828ZhIxF9teY4sHecS2aa2dZyZ+UZBGQech0Upw3JTbPCUOsj5+ma
1b7ohzicPnydKatSvPqsF34db7g65VTuHl9b1x1owNmCw4KaGImUpjkvxT/uf+Hn
NbNUuBlPpGTqpG7c1+p7eA++9TRmgsWc8ZNijp8v6ovHSDKLHBGKt7A7UgWYGK1T
5G1bLc8Ih1zoh83b5Z1FizjGRtkjjFaHJhDhKoKP2hJEoCR5TsLhdmXl0fozZeYW
M45UcuWvHkd2pdQJ6MJOLqP8kxppk5eQ/NkJi5k/ZSuCN/7FuJqr/BNL7xwabz9X
wPBE9o6NnmJVQ9MWgcYAduAB/VYqi/Wl5EGY6F3SC+7x5+ApBYBqWzL1bvCx1xj3
ZVKGj9FfRH0FmfOUNK9Ss3vVTOOViqMDKDC69TUcjF6I5RuElO2uv3ygdVIBSRTs
9ZYJO1S9nRQe/7WdHaEDWkG65zGrpiscYWKkz4cDTY/nKETa8R9qldqqIQMWraZm
46XfL9eIw0S3vspz6nqaOEFO4JUfaOI9JX2HOkxo8NXZEdxslwd/Ztne97qQ9C6A
rZ/HxWRtSHpKKZTbo0vEFGIYWmbcFFPE8S5it3iIAhCpizNmJBD+Pm4yNjN9GT+N
6jizMb7KPukxPjFQb90RB4TBeBvZqLpp/0aZ+/4XQ/0TKz3J1QBiX25Cgqr8uaIJ
ZHpeDcQTP614XqnKC4rqAvjd7R5KWRqeBy0M+RXYTUs+4v+ioCuSrIMw+7IZYZwU
vNLir+BQgzRPx6bDDxOOF32Lx6n3YhLJcw6R/BaluzZDLebVitVmOH2wftCnwzR0
NvgJJfShMLQH4TglsKUfXz0M6AKYGoppVTBxvCOlTItDafMN/LsooQQldJeGgWO+
U7d2xRsJm08WV/OOtaAMl9duHaWpK/YP+s+jMpHv2Tr+WCTSp0r4Yf5fwBL3z/FS
aikuBgttusAbo6HRW5tej7UT4zpT3C1KA9urpKed3SgjRVGzlzeiSSC0ddpMuAsK
6cJHV4zXf3QHw7FiDA1KK4ECGgFzv+MK+9OjeIa/SYZ4Sd6jtXW5jdUSUDl2K/Og
f3yl5CpBjfihng0Y/hpthuN6gdqz7VTJq94r/ziyzXd1+De1AUzmlLiTD9P9l07A
NOrbbzydtl01uosI7uV1V8+wS3PL/dKk4Cr9YSRrnL8qdC+XscBAUKAnu7PgW+CC
0zxdpWhdJMYLtgsl15vhJrjnBgnEZvYOpB8NoiYP74FbJ29g9gm+cdytP/RBO0Zn
EqywDM1cUBRs6UXm3PsLppuKO8Ciji/vSgRcyfSXNG3JDQTLMgq9XuLgdN7ro5A1
RbnbOsJpJTlv3etnnoINxmqnlkwEvNWOWpXuXy2cBuDrTcCGWCKlzb2MAgEXASs6
C+vDDNP75jMPzlX1MCcNeyk+DVVzRnAQkwNLc+uvBqlSJlq9S/4zPtEKG81A40cl
rybqlLwC1iYL21IjSUyaC0lWrGwCl8dxtQO9ypLjt72UqStbIS8IdumwTIhe8MTz
iiyBR4rC3dWoE9k+E5GrDYK1jyjM8P/j+rJuOMaZkchRq3jh/II1ZgBtxYJdtmpT
XWsn8pziT46hk8h+dVgVuKQFsEwkIMbpDGlOkOOLDdWCLCrKuKvweEQlPjDMez8p
l6Zl8ST80M1JmWzSFK7as8VSxClBzuQ4rLTygG15tk8pllJTfBFAD1ZqbobCXyKD
5cNTskw9SjiJVqRWibVTcudkrnR2FuwdMZ7Yp4cCOXZRLeIbphMVFCB/FyDji2gm
5HbFyVpS5SwbIX5FR22TvaOoTGDi4n0dfEqXQJBI19HaBlCGuMilqbQqTC68+EK/
bSRYdApiRZGwmH2d4PM6Xoc2LjdiMDYJ2rE8mRWpAlYlQ404tuVl47+2+m9DSg2r
WlFnjKIXNeitIpcTpb4qIbntS8wDY70Ku5OCbfwcwTS7Ry+s5n1ldX5he5XpCcyk
z5uw0NU/f3p1NmSqlE8siS1XgsGKQ40///wUw6MFOi63+nWkR2zPsHpmRqtBpyyX
7HKJQUgCKPt+5G14EM0AKKa+QsGytZqc4QPdYPx//qGk03dmwwvZD2owbHTRBl0s
zgsQwrRmiJgidbYCrfJ7oGNyBhqONRVfmeKQM7TcI4XFaxhdBNcSAfLOFkktrj7k
Q38OIbR4mgz4GRvw9aRNlNLVIhyIifED+yVMuP+8EqZJ2PlL14u0ep9nCc2VOwbt
vY2aBhvftDlkvYJ0ouCAk0KrT49/7lmECOFD+Ki+ThWaqX9hlyX+7v39JAk4KlR3
UIiDfvM/ul4PqRgyjNrcN+furY9NW5iUjbcFPImPKRZlz+p1AgDM+WbfvIW5ZIfR
r0InhBRULndOm6gMyzvnNL7aGNadb8I9SXF/pgLrBbZu1+foCaE55hUlWJGFFFh2
UEyCRFyyXB4YwQGAYLsFTtlY3eiG1hzJcdv92flZkRPJbFrxqMod2eto65Kjmoo6
JDTuSituHJe+t+Uj30SA7jxoAHfdfm1qm2KjR5+Dtq+lALV+POpx/AHBQTNm9e7n
DtQCd98X5ttVeLF+ABZrCJe/V6uAcbBZvtMu+QtEL5VG16F4IUndJjlWgJiRZL6C
fXocjP4SpDGv9hkaMSw4dBSVpWVfa/lCnJNbZGv9cI4y8xY8r+Auu1Q6a2eyZF5d
JNQgtNmRyfFGuJbne4zmPxDqUP6npxnto17aIvSDfh/S5DR3TnXwmT0vLkCne1N3
PMONidt4yvV2LIwXLP5Uhrk+MfMzQw5ygFHcYTD82yc7PwMT1aul5jyjMHkhauk5
hDPJFtZZ7d8/S3ourHSxIPP1FxIgdvnmW5L1dmmGtNUNfdiVKbidA8Ju/IFCHOmE
YIOE4mcPA82WXd5m932a6HR3CWT+jKhXYAl63YrsK24e18r1L0dq5cBtXD0Wf3it
iHDaBbux+2oBgOaAvAFmTdB2MI1aVTFT8LOxLKWK7KUgiFHKTCjq/YJnEyJ6DvFc
/TOWUl8lgaZz+CoV7tfgrDu7oiDlRz1owzOJISvvpZ/62s/3EbeECG8BB78lptLK
q53qoDI7K3+dlLURo/YFQbkoTB7sDoy824HaZRQBlDISCWpHczmD3qi7OLirzyKs
pzgEDkZEU4r54PJ8wPxoYldAOxWYtClr+F/oQPyYpPB03oZzw/yT6c9oeeJtnCJf
7/S3wU8rLg0CpwrOAhmwU0mdmcAndvRtHaQ6QZHjwAQdxCbAm5/Gy4kF6L3slWSB
Ai/yIQQIMqsbhQu/RGtfeXd/aPERPQJqN/7vKMYQP36I6PoPQlqFx3IS+BrNp6aL
J9QkhfdF/9QsKkHrUB2XxSvrgUWDyBlaqiGr4+qrNHMOw25qMrH4vortdC7Wt0Rt
YNkLsch5mdgxPIfufRLYCoKzpUaWi9N+DpENyTDR6Oeo094H9LcPc0UBEKCBTlS3
WijqUgHBkURmpnqphRp/zKxq0jMwO9kvvWap72sNynBZmlwu7ON2bod3O1SEfIDv
HPVMIO3iKaLbyltT7bQY/UwNjC1BmeVHPYS3x6eYX3umsN1KhyJQGNuUqSDbBTaJ
csdnOZwNgeJPcbkuH5kGRoSSuGIq1LEIWNdsai9kpvEhhdN5dIS0uiu7ceStK7F1
Lu/DtVZR/r9UAPjwdLTWXg84kRkRiH9Z6c1KKSLxQx/THLv2g3cHcRjnAKhOMvgK
QbzEHCvKZ7OJTxyknPnM/QpH203zzCGWneLY9jvD5+OspvRWG6kMIvhLXyijmyYS
eqOnc5xPNH2XMe/xLufpNE1OnJgX5MmNtov7J/epMNyAkevOppTrAdCgLIdt7rT8
hb5WQWRx23vRv32gI6yXosjsgbwoD+NRDi7hoOY0Bh5GyLpIoUeqKDh0SLzwbhQh
dr1kXQ84CYtNMEJ/Fd2RYz7sAvALC9Ha+MA2PuVhcQnaxIQiEhQkGqNXQYTond/8
xoIiqACqNR3+T3w/9luxI38pVIjFkGQwBwbJoy+Tcae8aFd2q3HhEWGBW03K95jX
I6I9ExSk0M4J5GEPy/6wRbrnZpL+l0Y8IlD/EOffg+8lpNF09516BEwYhpdml3HX
0ghg6GIIBGkr4fAXwq9yfI/FAcjbdPCX9YiJ306z+Efw4v+CRnsPRcytpjggf+qD
dTxAp2pYfo2N7enV4qsfc63PRHj26W4/pZ25yTN1OpHid2BYTKGT2NuvXiHRaFv9
4steK7J8VsskD5KS7NbbZcuZoprVWqWbfVWedUoK7cR7tfyLwcJEsO3XFpguUBM/
o3GlhemcZQPRnT/iKvaoS7xcdpG+T0sRo8TxpzT+VzoC3d51zF1AX/rlQo1NHyL9
yKgGbinfRNplYkf1tZx8FN+BrOXO3yqyLWvOXjpRaU2z5r03PCLZ2Rs+aRLKQuEy
aKal88QEhusqmU0Yi8tdzxQi8mhI6G6w5cdwCTCmiOsPpwh8Di0IHPq4aOg7gB9s
WZMteRRScaLL6My/foomqmjVrvQOjwWMnn38Y1xw6QVh4JXG8tY+C4sWDOEMRFIg
kXTNKJxD//5KZmYdgxDtazJ43T4XonsFV+zsZ244aRRTZrzQr4ZGp0r6gNPpXaDJ
iEv7vbzWfScloU9pXyiw4WXLXJMR1yed9JVeVqEjIF56+24Mnqy+ZG532YEb64Ne
VNjVnHxbAQqHcsD+/oetSM5D1LO8CBh1wFXeRjrhq3RUCb+wbmhbkmAjModymbJx
CxIzFXzP/P0AFcSAXnMSPW9DcU+yxJcB+c7Bj9fQaLQPbEJUsiOWDWj1R7ITxs0y
pZQ7FBC4A2lAuzXMw4s/umi4ldBDHivTdMDO87xGcE7GQhAeqcEknvQflvJR5PAB
TBNQ5JLp3jCO77YhUbFNLb9SGzHhLNaD4N3acg+DQn/ad6bZIySXZ8Xf/N1AbEbC
f1RegpkIM9R6/2Tz0HOv/Cf/DNx6q76oe3s3uNzZl5PI3Ino/GQ/nvAycAWMZQYc
ZoS9cCFFu8EqSJKJIzX1Jxwkw8APih6cm8v716N8ppNw/u/q1E4fHtIObDRV4K0N
0L5z5B9+j1PQHxIRrL02wH8shOPZZ4ALA6Z8KOcbpMM2fs+8WkjkfRkWQ1xnpy4J
FQjAPz7jFZ/JyMpwf2cmFKnhjAoVt7RV7pLSmK1YJNuceOmrkmqlfB7/5mk3xJv0
tiF7DN5szJkBBvFf7fqp09Pyif/XYVqBljXRnm7zktToQYqD2BAQd/1tDXOx/qXQ
zPCmwa/4Eu75uQAqTyNPs1k4idZWlfUtYCwZ9k1SEFd4SznnqPx/j/6ZvI3v46As
+1R5cvD+mVxg0TgnWc3mTNchMxI+1teY7t5wEJriA2aFoGBv0TSoZja4LCyTKh7s
mDsgnwG3LOcdS0yVB3KZ35VdKShtMVdV4uivKwTc7gLBlzZq3jcO4bmCKcpsX394
vEbnNQH/hETDS/It8ktQtFwXyQs3aBXeNvcG58O2KqWkPmh+6HYqn2IaOnK61iUo
bSD1CrCXjJQoqURdHMLL2+v9tUvYUA0R5B3iXDLu7IyYKkhGjK1ktt9r9IxTEKlq
gZFr1pGj3+Ft6A9ygw7TdZuE52HkqiS0qDPFxrBuFU3WAq0VQWvQYQAYLmtqLtjj
sFYx29v4gQpXLdAoMTwZUXanXrlvvwDxDFugQ1ZE6A81fkK3OdxS86/ookY3nY6D
0ZmBoPkJQwizOGyFJmQGuphaGl0NJcHJ9IjPlAj2y3Km8rtj/iFJMfTtCLvTmRG6
MiVuTB8UI54AK8uf9JE5yF3+ttg2hB6eZmDN5EA1h2F42WVem1PX8IcXHmZpwv4k
KsZOsdZ6p5drdvE8fNob1Y97IrPZNXlZhmylmYmcwqddQvD3RbjOO/RUxLMWEBoQ
9COxy5sTUndVRGzCCvJ/RJRTCp/CJ+Mxyi0X+gVeL/FtcuqRdWJ2q3vE6ZM7x372
Tl5POiIb1T4gaprZqIwxEUTcSvXsboAOWcPR7UqWyYg/2gR9Ka7ATzlT5rv1v02f
rE9B9sSRe0YfrwyUYF4RvIpVo+Nb2+fHP3vNWNFpTUlK7XJfDg8sxSKAwq2BHznj
phiyS3iTuqPsctvUtPCmTpmhsYoCSd9Md+Ka6sUtUkiwlNuCHZV/1111orACgyEl
zs9nFmrjuF6KvN3Goblugh6gKtwCOTYEm1tuVuD8uN8bo4PTfAru499OkfmF1ezg
ww1sbTgZ92M4kyzT9admGbNN+74BvZmgPdK6S90ZKx8drqi282GlgkqMrOSuJaR9
roLUQ65k/Skn2lTHVFtkXx3clyz3cP38evN6wN6CPi5crQy7zWxDZPHhovt9B5r9
zx0y0gwhytULSv8x0JREp/Qp9MOR+iDwCE0nPd0rdJdhFyb4AePRz90xewa3K31y
ZzNngAoAbJsdAvI5KiRR5MxaLqQ6ngt5YB8tv+0fB7O3iMvqXc0u+opmkBzf1jy5
8/+RBVD/o08kjf4474v7Lcc69ZN6Z83TizfNh/aesta6DUsybopgNrFuglTm2xUt
EkTNhn1l3Nxu+EZYTcZjWE+VG88sZprThYEaOwdQWJwyqHVWh9ZjumR6zuymFF0o
z86kDa3eYL/ijeo7PJnEJA27NtHlcmUe7zM+Pf+MZS2BAU2UcSqgM7/TqpS+VD5k
SQTW0TqwA/DTIwdeSSDjZQomPgF0r+dSAZFxpozc8x+Axft0BnffYOd1h33qyGvs
sb8D28pqC8Cb6et6Ea2UaS2lGTRj1K9MjfwUvfnaqaAsi+ff/aKIcCqDfohyMosC
9cIZrmPSQrl1nA5S4gF8e2rB57yNbrWPSvDn89nyT6czhY6Obo27jA8Uo7xzDOm+
3i7Bg3J4QQgIvJgL3WIg0kqDjhTNw35M0rlXvcomvjcY9DdwhLWoRo26o6SzR7Yj
qM+Br6xoO7MeDwKTnVWT9NIsn61oTtjzk4F5sIJdkcCvRFQBeGVmc+Xqn0fw8WqH
CdzHksqoRCxYLrtfqaoEKZ6L8LuB4RETRqZPLigUGFAClSVxL5s/KhVPKRdaMRAR
7UfqgiOAkmf4zFJua0CqDAOvF4XgRchwtJs90DlL3ei6EEcaKdN9rFSA5TJlOFNU
zz/QpR01cZUYrkmMnhe7I4qiY8oTWdbs6/Ff4AuPaSoGPyTscCQC5gjlbs1n8E1h
PDki+kWhGvdyYC8fVp0TXFxX9ERJSNGZVcOau62vAZN776NAjNE5B16Z5e8pWS1y
Xej53VAwsgPnVHt6BhKVblH4XCM6S/TrDpoI8ZT1/umbvGLqZZ6xMbEXSxJ6DVS0
6NUfcRzBhE4CyREAnyTKQwJ6AZVj61wD0veC6kjvQ3FZJC6tuzDb1+dPyP+LYJAv
qcpzbyaShxP0BpYnsLJZ+DVTtrN4vua5KBnHUe9opnQaNd/3ms3drlxr93amL7oN
2CY/o4qi3X7ZBZ7mwqtRq4/vnSxj61HD3XPzDzgsgmO/h/rFEjOJK/biG/h1sHD0
t0SjcJP0XA6+GMmnO/EwobvOzODQAEv6erkRaD8IlAoFKsa+O7ZtvtbaHF7d/cTj
mwt4DJzBrwW3f3WF+M7jg3FvQPf4FHVznY1y/3bu5/pw5lsbU2vkkHVDt7kH9ypt
Pth5J8IFXfqPCbR0azN5nXg5m4YErOo7y0dz++uUPvoLh4eItgmVrVGdfzN1oQbJ
ocRkslLFDWX+SJldoAOmjUEw+sftXXgz8+Em7+03pvVtqlKczuokjwq3eh8JiPrk
hWQSXgegA0bOuA32l/9DWixgVyrw29t5tx4liXQip5qzJsJeyODz7qROy1N6Dd+P
6Y6kKoVkANVtF2YwXSkrpXDElQhpHjK3oiys1dWd1XpUDxVBdY7X3OuriJDJs9vj
i3zT2QgcgNzMGTE5UpAU06uAP5+iZXdli5M3JY1Ch8KTwPCWz0cc6I5KCDKUDeYG
U1tNmphAHLDO25VbcuHw1+9lYXOvxKmRxE4GTihim5AlF4itNgUfLa9R97xdiB0s
S3q+NS9nQnDndQRt1stlvxSlLRbrdR80H0wRXOaMCPM951ZFzFEtaEOrJ6hi5RMG
rxDPKrcJfnpEG6g/dbCWlAlamV4UvTYo2wLgdclPhLO5RHJTN9aQwlrNXRo+8h5e
n4vdVjyIz6Vk+J+L9mZXwFI09bTxLBsksEDgc6CDrUplM/efF8B91SQ3u9/aosN9
mXWRFjCiwcdRoV1W18TD/Itd6PkADzXTmMet9YSmycV2M5uWE1ggzg8u4B3mxOmN
tjZNvp8pnkq2Gw3aBrtCaNlyplnyXFEAWPGi4L8RaUNwU++s28y+6rynFk/8V/uL
TWeJDLleZOEg0d5f+jdOGvVAdwKGqPuNc40Hqm4t+Tge5EG2flZQZBWQo66mjwHG
iXe8U4CDphYv3kWBQkd12xVoWeLUwiurCkBoQnnbE/fe/msAvLBJcTXveh8D08JK
1zfUKsd1W9LZ8gAQ9RUusUjS9fTvz9oup10eoRClDFFGTMqH/eh5l76QwakUEhMu
LYCVHAP4HSrwq16/9doXcM+Z01L7JW4oBNHEiyk5uHwNlOsj2HK6d/kAA51vo7HD
xNV1cwP6+T+wL2hGDnbBE1WCGgJj5YmIK8HgSOdFJSTruAV9gaz8b2dRkaNX/4NJ
qT9v/pDwBYHWibdJPcVrYO4R6ls0bMvFCGw3V+F2geSDnELCwvGhRSLXla8+bIqc
agiFPMs4uEvD4uT9VuMiuX66hyGvijCLvDCgNMsxHVzLAuxBypYtJPLcLDqIAhv+
RJKXZLuCAR0tA3Cjl854C9oE1QqQ9YxJ4HfUbQjbygRCv3GWnOtsa+ppssqeUc1i
0weO4KYJGg5emb3BUlVQc4SsaKMIyXS8Ikr+fO2U5YDrFdw7WP/LH1AJlrO2u2wI
CI6m0tstQZkO8d8iFSCX/1gbwG4eJ9n/P0COJKEeayM9UKHU1IOClbQEa4bPsdI0
C+ZNSjlSb1lm7X5pO4Te5VMuDzzW+oUWtjpnt6GcZ+gydvQqzN+vlRPaTptMvIf6
37moYJw0t93jT451lc0eVByJKDr+knI2Q21yKxYAJ5LA9OFEAXpYBKb131VFrzIF
LBBse4Hc+k1X1yPlVh9SdaX7SolT4dr8ARPqM7oohtuU0MwWQ2tw+tqpGdOkD2BY
NgbGMOIHLBZyHkoA4c28VoSipceeEbQqFc3L4xO/Ayb1ZUL1uR+E7/ZQ6BTApNop
KcJ9D7a8IBY8Ry1W2Z819k7v/mGW42ma73LT5iP+k0Ln6b6/6zCgFv5wp/34UsLl
kDdrlM8AocKw4dnuihXdojyXk/RA3aayeBViDno21plBexN9LmpNpf8fmm5bSlly
iZuh8inZ1vjLSMJuUlb3YmZgPrrKOg5bP+lZRVFXgwx5CHARSRc8X9PT4+cTAUp2
JWRXVS/ijJuDjjfgrClUUEaXtNK7jzssGKsj/+PxI0oJXbsqPmrEdR0H/n73tkNF
JPsPIbe3T/YGHYHudnvJB+NVoQQ4xe9Lgixl3kBxLpwZnVYVPNhmP+ZWZlFwNcJd
G5unE3VSOWJsh3F3G7nu362QNGtCFlF3U9mG62SvKn3KO0cAiNrEjYEDyLe8933m
xOS9IVSSKX6uVVsEn3gJJtc001hV7BWAP2xn9VELPF3WqnPvzGEm944W/o2fww+W
rpukpghdlESiHeei2P4fMFOEmLQrRgGUoT9hZ++CCQWTvNAJP0wrbtoB6YG8KwuG
mxi7SBMod5mTCkA4b+ntMnBDsSWWl9341FHq99ZH6OTl3wMh2UGNgQjbPTY4oYvL
L90MkMM1gzqa6DERVkWyPhF8M4rh80fkY3WMHKBv7MIJg6VIRWozQiEn8vViCGJJ
88hvyeiIbTMnTieIdypHMtCaSNHZX0Afzt6XWxNk7JENicHyRJArgXcOwlZwCHoa
4B9CRbFvvjbOtkBOV5NtdciUHBvB3T8yPDzToOYXgFWCv8pGA51r2bsTJ+jPl8+o
PE/3e3lULxO4nLVspnZubWdazwduc2mNR/tnlBs+gHeyo2gLGshKo2rcCJaO2rUR
UHPTB527wPUFIhQ35Ckq5ny3YpAIR1snv/ERN6L8vMyUJQ36j2arEO7a7sLeHpTq
BsQ4U14xdL5SsIdGg7wnIjG4ViF+i8FfaCdewjfcN3JiBBmaGdinSiYJ4+WHF8Gt
9B2PA7Tss5pAKD70DSNIFZaZxDNeyidZJm1N5VZ0UvIl+Mla1/Aka+JtZj+ef8hp
fQ6UPIRuWLxdhO98XUBKqUIHbUINW2iMPiwOAKdAfwFkwm1KvBY76SeY3wd+O8W7
ESy5Dr8cwfOsJpP0sLTkJeAJLoTBMazicSoT+n9F4qlTHjVixoyGdkj+eeHE1GQ6
7jbSzJrjrj0FkQkbWWvQuE75FYJoW3xvNPHwRgKOVxBBfAz6nkN4JQOe0FRSyMUv
mv64QuJulMpW8ubmPMxgHLKM6kB9ueV11t58KQDB/Yk5wRSkpcZrdS/YB2oiOW5d
Z7OX3YdJYNYVyJq/1ifrt+rgbOnnYGpG/3gWkkQd7hCt84u9GI2C+3qo4yt+oSMh
5sdnh1Z0E47Mg8RceVO58KtKsJGNbIaGg+fXQSNc7Fa+/mjPc8Gt5xbb3cr4Fgnk
AplG8vqLn+aoo9pS8WS7Zlcx6NJXwXWSuCD+wpjjte8+NS1g118KZMS6sRpjUi7O
BgZTOa08RxbEG4iFo0gPHiV+vgrUD4mQwnAxXr4NNC7G7peELKUqFF2XG4HQaxaM
SzOT2w2gK2xlU82rvPYXN5xN8jmnKKBFFAeF8mbLWl+/BgOKAkzox4YRiIfLPbmQ
tD6ZlBJUEiwVyL2PQqSYcdGXYXomq9oHygAkLajuRtlZq/wvKGtwAw8Dm70Gi4Su
9tNfR2kTx+HMQGNMTeHCHifqVWYYReJFQ0VeYBb/JWU9rmDCrilp5WuCUnps9CBP
X4Cec12IAldf9PyIi9ITRAq11v0teDNTEIwSk/xN4RbFjHWbQM4buR/4Q8bBgayM
qhd6w1yA6YxuJHh3os1dSeoE9U+WK0+ZmW2oI7kcjc96m3r1bvxU1a9aHniptZ4p
ZTrlBp2RRf5W/QFsw7bCsylhrQA6ikLE2LODuEWIB1HOP4iO974h3bEoKQuLb+74
Oc5lWxbNMtFwAFijWqtpa+k6yINCQUDQjQcKpctPCryAus8KGnt6LTJa+XuAAobN
GYwvz8sT4jjru70fGvYABWaNSPizD5R7hA10CZ0aiXPy58J2oNAt7ZFIDWX3Zuv0
sWPYOtWMe3jLY3/X49+7et3BwavlqUXrC5kpGJ+7LYUo19lqrLOPnMLDKrXPgVe6
E7aeeQ6zcrvgMlrO7tJRcT4EFDlV2s+AMBpWVMLgsKHwqljyAgXJYbq53YKW1w05
i3PG2Mn81WiPHfFkRMJ9F9mjeQcbNJ8kQ1JRNh4nBqj2OzlxfaxAz2L+HJBhY/fu
S0SG9SFRDI+f3+IYo0Y+DsMYKGMIDU6gquaIHXYQ7ASi5hcwcEAXPdqkbyklo8ii
8QFznUEP+IMVUoI0Q4Z1lIUJJNluFWRShif1qagY5/h/+8Q8pyntb3Ie78ha8GxS
KS8A8dVohnvc+irzGfkSAxainlF+y/OEZDKC62Sc8iCSZ4LLNCCQfRN49oXpGThK
rawrx9TjAqyqBzNa8t8MFAIM0kaoiMHCXZSj11xL+CuzbSWcZGpfQRQmdDkVYbtL
0WXTwaPwwyNuPYxYXYpRLnJKdHcuZprrcVaJLfmnCG0gtbniTGqdJV+4ZtUxFcAc
/quavwrT92y+sVec4+z8PWf7Zn6KOudlJJzsEljO4Ul0QhZS93DrQwFKAE0DU4+J
IbmCTJy/PIadZhCgGCzCE2TsSTbOpYtwqcq9B3hfbUuFKMmenL/7f6L/0QESAe0a
tqI7ZQcXva3i4Ue+s4am1o5mI6kjvQJVy4omLdPwgUMAm1PHG6AeK0J4s8np+4xk
piOucY6gbTwGIZTKVb2mYVJi3s3TjD1EWPWd6BRk/JR8GkpbT4W1qbmOId1khyfY
WU4J3evEqsjn+VsUCcwP5poB0GS/LEUmILaSIh/y8lPlpuUF2xaylY5u1C73xjrH
a+XFFv+rbis//DNLJIh7ZtAbQt+UZYsH0hQ+rJaQfhZgaKbS1GKYGKPWnFkquRC+
7dK0+wJ6t5bpGZOBXplfuW2gf4ZRERE/Gqa8RnfgoR2cIZOSWzD79joT+1LOdo8U
/6TPdUJY3d5b3G4IpfV6zvXcdMrp6a+ihFSGHWdsVowhsRimzKXhL2bRZlkPJIWl
mblzIWM+ERyN+ihoXysW5YarDkDhoInbgGZ8ZvY5zy0I8ram9K24GL56KHB4/0D8
nBSqEXD3WMwkhrlnapxCahxpjrw1A11pUVB+cI2/2ZHdzeA5NmyXQV6zCRvMzYA3
T84xPYNtfjModCRo0GvtA4TjMIvNrdD+vnM5HesVxKKFjXPPzGqA/EIxJxS9O/o1
G3LON3qnTAjmlpS9ibomIVQ4WRxnCLqBvQrXzi7k7K3v8ieyrXSVByMYKQDqdvdm
m9PYNONRei7rRcZTHHVihPgfo7dH8I+BKvpXwfkj5lMhwzg/vmf2r5vb8XSp4ndv
eIdT7btv9UH6rSAVYu/D9ECdCtcCuFb9YbnDyWCOHnuBAOpd4KB/4QwPbIgilUbv
0FmXzIR1h3oTc0MbYNgMd9vFvkF313tE9v24JihTMBAqHWPY/dljDOvusm+w4Bi0
/bHJ9BuwHUADbmepF6ZiZS4POEdAkekVLNLjOvu2eGJuLb/UKj0QLov14ss3A74Z
QBP3MJqxmtCAzXtYZEbRwGoPBExHvbO3DNqvAveaXrhi6Od+ibk9Z0jiGcGzKj8O
lfTmVmRAtx8gfUEOFUVFOFupcdW+zMKu/hPdWYEKnNJfmq66nGdIimWGysXaCxFA
IL5OqxG3HtH50e7Zc6hr2yGfawVkALJM2qFPe9kgbZcSHC3mLy73EPd7pZ81EIy4
yFn2Tz2RPQWYSVA2GRqBbEkwDDQ+/SE/t8fAawfW861YjVsz57JMpZF9IwX1XarB
LTYF7pcvycDwkM9beS6fscrngsymJAUoODN20z+f9W2jy7Lp2UzDJZNGfQrz/9Su
6MUHgGOVUqx9C2Q0pnVHlS4irj8sDW+vpUqPPlbzpkHyU9JynjLw2WNJlrCNoKTk
i8UspneTjak3oMlmNNitnnn8UcNs/bs4/Sc1LBwyqRPgEbzSqeIa6ydBk1dXb0mJ
8L4DWhCre86d7RLSA8jngP4ZwOYB36jNLwS25i7UjANkDJeyQ7kTARalvIdF3xKU
mO/xGzCSbVTa84E3Wng1HOVGNgm9PfeIQVdXhugUaq87W1GdoXUacKtXy5cmqkWT
vpRcvNSnFA4xphbylvt/LR99y3rNESfZajARqkEzvQh3oJ3ji/4ktkR4/rQA7j3a
d/kHa7f8wdEu8xpYkjmfJVB2EnRUQrZk6dJaeJvVCQrSNvN4fFyHCpkUYU1O4nk3
G2lkfMSec/7GV+8YpkRLBhPbdbGFPDtZs22xla0KbZsx+uhuXpJncmKdjYV7BGtg
JbrtImKeXAD0VbVDMCqKKfpGmbeCYT4qnUBPJ9D5NEWrwfDiLjvvEUTHi3qpfcMW
yKMdfxLDDOxQknWa30QJDCsMpxTI2i/9MMWAcGOuViOfrPtni34YIYUzFAK5sEad
czZWTG7Sys1Vcm20nH+RigxiF5+MhMO4m+NgNlQKo40dxH7Souu70M90/WrPB8gH
KT5PIroCtTnuzJiF/StXE6qIS66OiemExMvqeU66AMIZkLQCub8uP5Al1IAnXDa5
3VFLH3GtuGxQGheGnkseHjIHKN8PqSELwbKSFynubhl9qnuqII4iDYmTgdMeu27n
Iwdvo2e5OM68lO5v1etPG4VKHZPn1d34a2rIR4yr4D/dIGofTpogM/6iJ2RgAOTb
bT+gJvAxOshQt2WZSu2FObJ1+kr5ImEiCa6AReR2FZdBeAadfG7aM9kKV37xSoqz
EuWwgGz+/di1J0/fxvwzV0L1J+TmTnHjPUwYcSXacbWoywvwYBs9r9iNH/yFpqQt
nZK5Lf3PTgUg3O7lfPCtAoWD0/qLvk5t7DYDSBCVTQIOJIXem5psxN4UhHCN82LZ
2fm5BEOkT0fomLeli1KkDriAvwXjwBSWYpF3wp2XN4P5UVNvOSW2wc8tfwsaW+fP
8kk8tkWwjKcBubJwMLkes0BVpR5m1d43N06v/gLfvFKAbZct6n8CkAh2bHkC1h1K
xQtw3uLwP2Q5AqfAsZLn5mTiwm5LG+E9UDbVyZ1NLW8GLsGwVqu5UUUnOVY+Hx0E
yLWfNtE3vsrU/irptPouyf4TaBvT08Kh+o7yrooQRQSU8JWr4m4gBItiBCX7JGx/
xopu/QBL+obXwOOkPzf1YnGkxu/z7UkkXPQuIc318ICMBvzzaEayAShSA326P/8Q
3tq0lIjkakdKaRpEb2GNQpMquM4t/azjHxJ8WhiJP1xvzQAKR9SSvULlj1gF+j1v
FKAw7WTcB6zUlhTqdSa+xMxJjqtNAR6nwk/4dv9Wof/NDoKhZd2iCnyj4ednWiI6
OCSFbOFUTAboK/Cik9qrb/d9JXvMLMZhjpxahB0EuwNDQphq0nZnv1n5gbAYyB5I
JVFVVhrP5uqGMIppcSP8guEJyRH81wD+cCxzhuq7TNYq3/nX6o4A0cU2eyztR81D
3hT2uAsrCST++HrH5hD7L+Y1RmhAYTkt0oNJr5Fh0YvyCM2/cBLCOlAJM7V9sjYW
I1IpxMoz+QDUyvp4rEKEsRvFtGZ60zerosgJh4wUgn1jARkCUstpwgXy0niu8dCt
ou5cuKtXPpTh+5RG/dUoCVePABPD1Lo0XMkxRKG2gKR3V96Ea0LJmfsAY/MyHehp
caOpLcPwNjy7Oagm8wmFPATF0p+aDJ0J14Ohh57jUeITpv1sPzdC1e5vMgqKylWw
bDrRAETflG9Wz6suit9nU685ABGk5Jg34T8c68fl/GP5dZA0RCNo4ucxf46eckmz
2+TSY5H2GChl2stOg/FcWUMSKMtt2mipX/HtusanlTe81/2ARZEmrW57ehgCeEWY
YP7+Rxp4OBHj1iS7/ngkvyZnxGvN8WQtT5kCst2FT075Hm82P4kuZAu9/1DNMOux
UF1+rpaQJORXHQWw70AC/ZGGB+04bEqRSbbbyvMV6PwWor3PMuk/lSKNDnYdrC08
BYgs5q/cBkboWBnNT48k0WUHPuFdIaQ/L1kevx/GySD0hgcCSQxyLLM6xkms567m
0koeccAP9PlRC3buzmquFhk32/cUFUeWhM3VDdnkbJX5oRCzb9DF5Mkpg2q5GfgU
SUGJsm9LmwisU3VHzWrhL3VqXG9A8ylpHWEOP28O2IkNs8jJzpyw9vgPlLJnyImT
PpSlpO2lil57BO5iPZJ0zJY8FR+uNbKTRdnHdE9SL10OthClen7mUHymRDwLFO5z
mIRFuCvyOKFLuH5XQQUKPQZgH0yWV2si3ac+sdLVZJwPBne6v1+a/pyx+DyyquGl
WV3mhA9N6IjG5Es1ogF1uFewmH+/wB03WQMnCn5wCUQHAfn/CgWTm40crblAndYP
EPOBedg2BEnJ4ZVmv/8gkLzy7L5h7wCurOXYsEYgPgbZBPkNVx77+9ZCpj3nsHqU
Bt0FyQqdbtvvQUcM4pRjVE6fnJVdINHaTxV2Ya1WX/QdoDfCdbtk5BLrIcHZ5jC3
sIOKUFHOKf57Agt6VgfDyJx0YR6j2LC4ckCRNzM5xP3mxJZxgKWpgy3mh4Laj3mi
jShwCsXWELgh+2Jn7MsgxODzS2bsssSd4Wv0ZL7fQG+mveJk56G2Yjg1pgBLNxPJ
aoO17tuwFedZrLrdPVzmzh1NYkYxaTCQ1ah6lHqh0QTmF1LUZ6BW099tT+zA/qsl
CuFobvg6eRR/zj4Ep7sd3v+nQyIDFeZ07epl0m2ho08qXgOunZ9bTcJgOpqwldje
EPi6OnRyMccOFRKsJY1tMENRDY3iOQQ72l4pLHwIVftv/R7n6063+PaeSv4jGEwO
NJLET5sFVsmT+NYJdb0CxBTUn2EPrvdt3b4XMkz955CZbTnngmY84JlMt2qFhNJz
39ZQ913nf/vvDGpAD/54BvxbPti0yoZ/2s26dDkj+GCYI7NjBg6vPbI7k8WUDo/5
9mhV9dAUByt0cceAooWA6UBsCPKgFAinhMMu7vDjculR73GLLvz8kJmXDl1MAlKj
c9LPw0AatCZzO9najukuSFE8G5AVJPm3TPT2ZLwXYRUKetIXjQkHfyQNvZmvDiac
vzvzTnAEHSWOVTzzyKk6pgyEa5aL3f0zVx5UMDK9QllJ1utwPsvkEm2LOj+6drQp
Lp22aBEY5njy4DfodPtvFfdfBKy2ulBIBOaEtOqZnofHYWg0yhjRV20m8vWymkoV
YRNDbQl3LDKsNnlf5OfS1eDJa/FUYSdlXP9slVnVt8bMQj+6BWjnLMho+bbJwRgt
/nheMVFXQbk4+bY1use84LZolAcNTf/8WNoIu0zfIB9pVLsjkfS2xjJmEpec/3QU
yznLAifegbq3XZgna0ifdN+8tOjitAYN6+J45w9L5pNKKhsFv3CPV3wnaL7L2DHN
/E/brICe7lYibD+5k+4kMsEkbw/eqjyfd6kaoA7jySCPWemmkoWrgqDjWovOqzqT
nNlgsL+nxN3V3WsCjAH8T6v8Lzzw83whcsZ51IfDW9BpbFJJ+sApBv5SlBmgqXU9
DSEpcDzjlCFNtG+3f/fSRFC3PyhW7cp/72RifssacK282OyNhaNHJe6D9Zb1l9VM
kaX1Bvsi/pk8ZBDjGJZ28rC2IpZdzW6zvspZaOBDc7DXPwF74Otc/LynnANr/Idi
+iVHFKKQlFr+yOeB26/mB0TP1fF4LcQmlGtczBJc9usbevGvai3onz1NghF/yumC
WeOLrE1LdAR03zkEgQryk3P+PLOKGwJNQrNrmOudUdzI811GJQBBcOor864bpHfw
O6+4NkWf791gNaCfxzJ4x/P/Lm4jSiF03mhMZX6LQS272AQ+Z5y+geCHMqxk2nfL
XNO4qFEyZECDt3ugL6D/oVarJ41uA0oC9xeUKyNl40o/S7nKFMGqw/Jdb9dMGDXL
QzxnjFq3QMGh2wNRnmDbHDDwyKUnYgiLJabXqiT272jIsf/sbQ1gal8TEA7c7o8P
kYNT/4vKCxtFLpDpxuE7barLWCXRauU2L1+9JnP05TvG9wURptDwQQUFA8KAIJYl
X2Tsr2yDjwosastWf2V/P0et5tFc5cOc9StRtbXsD8797ek+4nfRYciJsQmnTF/3
DBXFdL4/LawSlf2msOdjKt76yZCH2XgRn5eqayO6H8HTC/F5dv/m0i/MUxj8i0nM
Ck3whyQKkuuYRyww7srPX8xs7nG1OqdKfjRmnqJ/kNw0dV0IOtFeIT1sg6mCA1EX
M3oZXUi1g8ukB35lWxB6eYccF9i3G2f39p+LkSGgfjXXVAoSaBuyNehlTp4QOuwL
6O3VJtb1iBHs/vFv+ab3lVuXf4fORSGulJjk6LtkTAuwF0lTca1sR6Ou4jLpbVMK
9Uv/Dj0hyua3OJ8ABTDnorXr+ImP65+8xet7Xaxeb7vRoibZWb/KlgG+JkiSbMFp
90fcu+fG6xyqrlRNriDdUmZqgHSoZ+U1bZeOu/qE2zj5PbX0VaLx3GbuYqQIzhP4
5BiKgwJgck+x+8nCw+WzA26zk5sqV7opk5rKpUMKo331fWROnaedl84pDROf0DS6
xw6yiIgVz+Xjpa85qj2p8fuKkk9aErdiWdAVQ8699z4lJtmW6cOY9lxiPfD8Aujl
r4T9nODNprZ7Lvd9tBlehAlBso8g8c7VgqxLIok0Ri/KlzzK2jsxcfUYdvmeeQIE
r2j601Jzf4yyvZldANbVGzwPeqQk8o4ftRf2rt8q+Gk4A0suAmNO7+dLL/rt1nVp
fNXXQkRneXwqbCmmot/2kQlfkSqSV8OgkeXw4bGNzLWFoiQfHHX2rDaKmuUgDbzG
xARYNiPDsnv8sSv8+ajT2hta3F7QnaiA9RuovFVsnHDwjBsROqmTO8bbNvG2+HYQ
hQIm6VYNsE//meFCB8SmGe9gAnTflZC1xvocAaI2TVEon7t8KF2oa1pYrP2nlIGp
NMKSj7q4dEYeN+LfuyFy6L5FuHQi/Rr1i9Gmg9ElX4zQJ7erJoiay/x35sp4K1Ii
YVmLEZZKMOnIEyNjaL+1WARp0wlVEHh3VL9K5fGW2HjUVCWyFiJqfsmyGqOdc/4Q
f4MwDFQxoqB+xQSLjYdw0VJp+eA+MYoFdwev4GG0KzeOfHqgn2XywF+8guiSp1BX
Kjn74xLGSKjczGmktCZAtMifboeLbedIwv2rbrea2UxJCSYUPzpE9jtNTBaEVRhq
T3xQtkYKbFwPQ1qHxkKXhbZjqWwA7fHJhxvAqMSNmk2gWqt6hohVNmyWWjUCn6FP
ndeTSBZYgbWLRDARfyAZYkx34cYjWX5zMnJJLrbwrtmQWCQisCKAg+WzTwSdLsVn
3GSz2XIWpv9V4JR1FyWZ9/BRmz4AY1ywnMtZwHxBGy6meYAUhPpjkvkzXam3RxQC
4klcI7k8Ogj+Or1lgq+5DiPLBEuOBFoe5IUwGkPSD4apVgEV2eySSAAbu3fTdrhu
oCVEyWoKBDK+84k3gQX9Jv6PByqP2yNcuJMEDw1xxPcTl3ZxakbqKnytFG9TV3ae
vpMEkV7KCGfcBL42ZJcKWSoUuI3ZP4rUjrH60cIdA6agSBALoNGOv+7u8R9T4BGu
tPY0u2gTSMIm1E5ZoAwI6OLUgfgATlA6IOMAqdevHPdUFVgfsy352Isd2uymmthn
+gGCkDCHbyMil8KxlIHviSewTen0bI+rPQY2d6OVNUFZacL0iWUUBRgC3GCDXUvt
WlkXfGIsNfTILIZYg+WiBagtnaMUZH76Ffkf3U53HlVfOMPHXrW4lQKsYb0+Rvbr
hWWlK+D+Vxzes7vADcxWo9WsNLSCVTCA6+21BK1P4rZQQG65vIfoMbwgpDTwT1VY
4i5MV3jM76VyyxkmjKlauJwPfDClTrbWIB/oyJDkvQL8iuXdTHAflctY393mnrJw
gcFE6T0Pw+0Cb68qOZ5jZcVzU59JtSQtiIMt1ydhTUlYk628f1RC9dY4eVxDrHk+
7YkAxR6j0OwYPB3aazZm4btvpxjv4fUQ9y/iaFXcuclT0I+Wr/fnuhlQYCCO/wTk
fZpF64zYX9ylL9A/PbmQr/05+XIpRaxpxrOr5KWqSSmFyw8AZAnC6uSi3qpjc8Fi
IHo/HbXMBL7AUtpit1rYIIiO17LQdjX4XAIi9DoBdEduuGhlbpJMA2NdZOTGQu+y
9dO3YGVjJGF8QvUPR49WHssOBpA6QTnBNp9XYuvARHjH1RTTD0aUSd7OfZEJn2bQ
cGdk4n4pgisH8pWkHalFZsqySDjsU6jP9xaecTeNxeuxu/EJ3BBoqHsKly6QumJT
tyMkLwJTa8fySc+eClcGCPqc8uTTvFNLNb34bgHo/MPnawjXsa1Pfkxv5cCR/7Pa
WApWevFS9kdFMszkJlxrZFexSdMzjX8bC+l9Sy1xKziYjQCCGDBTsPrDkl8l13dD
v3oosrUATamyg6wIUbZd9hZ/R6tyWuH9ZYQSOGHo+FtiteQJJ7KlMfskcgOJfSCo
7Lbq7itzaJH+biVtTu3xXUrKuzfgXUmMk7L9CJhJUzUqhLt+eRUKt0iANcQaYGUk
LOIEtloq7e3BBDvrdCdNbFkZ5Q1SXMoXarEGKeoCe9jXSNCDwIlbV2e4gOH+7Ezn
jlaLPYqcTfZvSZM8dPTFLKqiJYs8Ch7hJDgQFn/ltHNfptHpWTBJg9RScj4PDmnq
ddEtqrxsQ6tWwK8bNf0gA42PfXZFbrisbMp5Qjwh3gZG50ZBvVAJsz2nJygLH0Lr
Ohr7XJGQyv0diZt+9QxXx4IX6qxP9qTH2HNuo9lRkwEoFFWvHAioaXQYkStkkACA
DbY6NhXmNyDOSR1jtKRz8zDcfTqvaNbQe48TWoh4DfbyTP8QAeEjmWZgFe/w0U0I
0/Lx0QMt0n5pgGlLOCY1QfphaiBOiIF1oS3etZ/ZTqCAEX23e/1V4H+s8RuAwujZ
ukZkPBu1dGGzkCboigzH82B+WdGhDjJqI7ARK4ENRMvpHqzpp7P/cfCcPw6Hpvr3
+jnjApoyLjVrBiCuKK5Lle0z9w/o9FIFj14iMNQmUG6gFpBPR7cywzUectDZl+x9
bvqory74oPrWMYsNQP2PYOkwq45nNp9bZISHqkBdQHJDk821rkpf+qGhuY62jQ6r
g8F8n/4YunG3ennR7EjlnJpbrBO7qK8J3jfh6s+UQ131zulGQ1UC65KBAzqgVT1S
x5BlqRxRCxDrRLcK7p9sv/9aDf21jDRWyUKbT9QeMJhodT5GqicznlPsW4qskSgJ
3MJzBUPRP826d9viIhYPcsp6iRGrIV5Ul3FlH4uabiPp1tFeNdzzdVrSpnPnQh3P
7mjVlZoB0Khi9Wik4cvQxTkMBGizDIQXszAlMXbgCuBDIeO1CsKMVh+b/VC2MfsG
XDpomlnvYFCwFXuh2Tc58hnEcMU/llcPgLaSmIGJC5YILthq0Sk+NRwnudPeNwRB
Ub8VTjsZIysnCqEOFNLQK8RbYjKNELQIDnLK2i/MiYAxXl+wsblo3ycqzOiA/Bpa
N7tCUen0O+AgWB4monVoxXsddNLyd/3S4EQQtmcTxrRN0EWVhATnk9P/EJzZrOGY
ogBHkWF4VMr3jSxmZCrQCdTMb9cm5aepaAZ5UrWPRT6GCPe345FWAzefwD3GGdrN
TBHVz/o4dJajkAe5vUwgWu7KYMjJIWTiib6kvejfPW5OcMRaSpwPPUiWJuVFCIhd
5xTYFNfx9C+O+KDMEIWms3FTlLwNXnMAV/nG7RDSFotlHQSoOPSLRGkCEwibecqp
67DcmN3fEzTeIL/v8PH0FGkr/+9m5XNPGplz+BlVk5r9/cDI7702xYThx+2lvYXt
B1u+B+Mq9fG1Lwg1okCEcNjW0DILIlIfX2ET0Q5aTEWUhdBGVb7J6vjkHP1PA0Ie
VcWl2zw/DP3iNcqja9ObEBBuK5M4dmuWbZFNGVJwTXQVpGNLxJljwxFf4+BEdql0
Zs2zIRrvSf4qjqgroOVRrQcQ2PC3YebpQ0ZKszj8p5LGrt38O7G7834/vzFcML2A
bmvOk8ROz/AN9gg8R33hHTrdy66gRlmBKG7dMXAVTqD9o6VJuFYRbdI2nydV+eXb
0obhbYtHgHiyN3x2I+vuU7DVall9V6jRPmvwueL8qACVP0OMh0x4HUIaAC1h1940
TfwDpJ/DXhZQuVJK2wk4cH/SXl3fl0QRtAdwP0bKtSOS7oEOlRVi3Tbu3rfiGDKp
ClIN3xWG/vC+9aN+YCarxyWWZ5o8MZ1ob76JGQi5N8rneu6FTD5Od/zWPnerTUm3
ZTioVJLr7BVbZXb4/UIwp+fvmMtEnsNuXjooSxg5qSJfQ3WReL3XVJw/m6ugHI0M
cKdIHJv4NMXAOPdQLoYlxwPA4tHXl+LB7cEOT7Nu8bHGPhLcUEBWefHUDanmcwAX
kk4culUAZtLOXiPV0q36k8lL4QrbBj0YxfarSo/dafnkYISQgfVQowO7whsp7EUv
VxRrtpn/HGUjukGtDyyUk+4Isj5datDXQuqM48Y9V1FrtB07g5ExsyhRHa9n0/fB
RvY/SkDQlctQfdQsAaj79GWjhsnaEbjR+5vTxV9VMvLVLYWqStoFNkaDxCyqjvTS
oFNvGW857nyWTFpNrOzfFeQjyNWKVLqeBu3Fqdx8Pq9juEQy3+aj8EiC158S1aJQ
PH6SgekMxJbxu7kyY4dQz5ATzJJ9HOjw0uEYHBimbavXjiNGr6m2z+eip3HV7h3y
1fQREgs7JlTrl7w3CFMvPbwg46vb1q14Ud4wUywPqxs7B5FEVDNemVKuk+ZrcGu0
vDed5AkXt7Xh6k0aV2a11ZLJEyT7WpcfDNpHwuAnXkpU1XHiVoKGY6xlUv6UpNdP
NVCNmp7QsF6IQ8Gcalrqz5o9RHXGzOuai2cTxD1u+LYp+mhxxTwCFkT+ozP4utkO
WZbc5zdeWD4xm3GmQkalPTGkbWLUBihx8xJf3EV9vhqDk0OAKbxFiB730PjgIHmt
3XkHU1SD7mTAwHaCfX57bzeQzco0N31Yb3BrEjhjQBI0ptoYe7qKDNybDrov0MZQ
dglQA5Qq5n5YaKueRSAwQQPE6tchxHbD81m1nSrAdnu7ImzXQ7q63jh8AuBB8HhJ
WMrVaT+MrztaRnoV8lKRKL4HFyTEQUnUdwIr90AElJ3cc0JeCqkEBzyCujinfIS8
o94vSY5nz+QEGVMO/71xecNAXTaGhZfqduoK8zw/b16sEL6NTF3SR/LmSPvw2k5G
0vudMGgSDqmDvhUMdJUZyEhfWGx8nDw68LQIkjnyhpD9KEf9e5m29Tk7fuSG7d3f
kNGhhT9fPqMsBL32eyULH/Jy87FBYqzGsLp2Ze8qJDWUvzWfMXBzE4cVDKGOohLN
sWqOGXbNt9vMhiwmj9jaOsv9NdAnBsBYm0+hXsZfbjuxks6sxj/ekUeh6xc18KFP
VL91MLKppoe56Ko4hkGVxlzigT3G+lNe7/6sso+u2SWaNYEdUgoj7a/eFn8XdSmW
SZQG4lJrnUtJGeAK5aXZVZoWubtbYdyP7Di95KA/JJ92U9iEfYb3GpNl55cx1wmz
uh/uCyFHYrjO4wUUU064w+Fvn269u4eFAvuvpi1tBBtt4QeKnoHpgib8pvZVcBC3
275wnzt5LBDcDYk4V5wUNqKgtl99ygLASQBwyBsX3npYrDB+PzRhDFBYkrn09OFL
auhaIZSm3gEvUQMgforQIm68krOQzmvfydJfSjlXIyyXNugLn6G6EN4kvukIzJ0O
GvmlofphWBYzUTCg6xR0T44U68oY3ZhcMfp3FSiIjkEpcZKkqnReDR7n6WwahV5e
FNBQa2RRrK6wsdVULTTsd3sbyqcHF7Ot0QYRjTa3H1hFdoItviNC+wB23GwXfw5L
8oqB20ZSS39MNo3n28BsdQW9MqOoJIQebvEqloxQ8ObWyhxvfXNNtd+hlwHr+sMG
s3Qhlol86izpPkgT5QpdjGFZMvj04zivYRnom9SY6WxBCCSFc4mpG7n7Bd94la1j
mX8e7BszJF7A0KEQMr6ekJMhB5bQ2XZKy+6hzisXBKsvkvQLfr2aIWaAY1m+J62R
YRcklsa5v+CLuIXaPxwRfOKIplfI24SPSFlh4wFOpUn/G5PsVUvwJXMRr1D63IF/
drVOUz63VgqDK8oBYFAedKcKtM23d0Xj9sooY+XnTcIhmCGet8yqHVe5OmzMHWZ8
3MebW0QhBPxMH9vvLtZP9lfNEjwd8mSBjwnkXwxarXnREqYaj42+fYwAldKVHKu5
arrOhjtHXc0fczqHiH9QAoilnZ5beYeJHoIoLyAHXuGvRQwdt5qKquIsv7Jp+PjG
doRXgR30/7QKrhF79aM1HDtD5rtRSfVRfX4Tr7Cn3UNfo3aUdmv4y1AlnzPVjHYs
Q70p3heXNWtBt3gYM2kLfjMc1Tjrb30CI/2DX/lKIAW7f1Adxyz1ANeA+k5i8F+A
/RgFTpsIGDL++2ivzG8BMTNHrQglO3ANbdPHG/ZJGGi/v7qbYDm8sVlmQOd8GYJl
yfQ2gED0StOyNOSnW49sRmJsSQMYyFLGXdKqvw+ECbJF7duiM5vVpZLkm4nnUY88
9wWJ8q/5uZqmS9X3lGoTqVV+KcKevYrQg31hiJtJocJyJ3HAGxT7FMcApn8kRupM
83fI9nrtzJUKNeC36BJ9R90rBKBnIcKquNi++sOHzaaSsEGyKo4xpaWdZcGGgUov
gG39z9hdIIPfwsTcEQ3rUdDX1YzElUB2sghw35/wdL8MgLrzWXXhoubmnqcT6aEN
LQKHUwENXaze0IDVM4iJsgdiDMwFVpO/HCtOMqowasQbjB1KiJbiO7yG3rvGN/RJ
4qMLKLVeNRQ2q/lxxeCIuv+S5CnzpiLVIiS4ZlAShxxb90IlatzErsIvECKYvF5k
qDRplNvEuQ8TtSpnN94AjE2PGAjcCPp42Mu+7LWyp3jZpy0LTb04JLwjrlW35rxx
JtzZgObkYIrSn3MU/tCYeRj6CABJVYljscNwWcZRjoC+jtlYalWdoTuJJ3RDlPqA
DEJczflbshz7vLVpVzI+YvdErd04zPG56VvnWmqFo/5dm413tuFHf/3zX7bFE8hX
WhdsPG+U+iNkya9L0F8W0xfpyjYXg8EydqVEROaxT4eKAJDOoKwlWiDgVL5Sgx92
0Had+VDuZc7jszF9FxGG+yymWkBqTV2hDsZkuqvi/rcoX6IRAFbLOwlEmOJnQSdz
KRKFSiu5KV9kkk1nJLbLlZGReZDjmPWQR/EMIpW4v5UOyeGxvGvqvTVYFhEkeSOu
6FFkMhQFMeuTF65+wk1PTlxOl5Wgugb7Y3RNwFIm04OKmHcvpjBNVXEmpNHJ+avS
wBGiffzKCFDGthES0B2c6vLEv3qPkeERAX5e3UZ2SfweKnpv8fL7siJFrYiBGvuM
Ec49+Oi68pUl1wwNh1roSz+OrFrRCCJkwzR7EQI7yssSquYxr/cqp6YlA7PH467S
XhahZqiix4OJ3YQS7qtAMjewlP0NalBarFoSOD1Vr04cObgYsOxxjye11HmlEWOj
FfxEpWmTsJNDWtYUaw5z0v7FKI1rSzKhbLvQCL7TTONTgN9uE8/4zyUktc4yXoDv
xknhV4L4jM8f9xBzTfMy0qp7WgJprmYrhznBjPPX9eADPOy+W0jnpSvKTeiL6t3J
17hgAth8hdrZt6m7ITBlLKkVjQLdcBD+b/JSIwECKDt1xIMSBt+Fe5Fs1Ydcnm2W
xOXMsrPDu6XA7PQbYkoKP8BTUV0G7o2fs7HRXbWRSlxoaIvbs3i6HO+O1NIG2Dpu
PzcKCsXyl3HG6h8Yqrze7YYajVJixV/+scUTdwhIUrsYgY43gMP60h7qJLO2HY3n
vHLHzAWXCfzvjkRrq38lkQivi2eCgTjFHAtsigqH74wxo8pp9Es8WsPvM62/FXS/
tSMGyDoBLPcsqBGEtpQHZv8oFtgJmQ8qYKd5KbwUUO5drtpeNuoVpZFvsS/GEAH+
aXpni6qDDTV9hQ1elOfZOmV2pwJ1cZeJQ1Tqvl++PQS5d5c7o8aPTMmf507rxjQN
8uuB8FaLzT2+LLPPddJJPb0Q4EL16WPguYgOREoxOslCRjusM24I5u71tfH7FNR2
CPO2D9Q0QnP549ERy+sBc54/We1fKrriyxcZBZYRjB6b4u71bXJJuzTAdvfnM1Ln
uuocQ3eoEt7jykiaWUb+o2maur/MJbDXofwYeU8wQV2yuliHU1hhz11U+XQlRfIz
CX7Q00im5Bvo46iDxNHzzoJ1nyRhkNugN7hmA50bghCH+JvjgX0D2C4GaqFEXnGN
SUYbuwV3ahnQI0AQOYrmaWe42pSrsxfWYrGQVhchf1TVQqrI6PZfjP5epLmfGGma
p3vXS3kTaK8yo88q+dFc9zwKVIn2H1fCpmcEgRT5RhynGrtL4sNWa8wr/OJ8BjhI
xdwqPLHogY0qhiGl8OFfdpsyOFcqXaCvojgDgaBz6Svdwz93XL4VqfwY5iJCnyPH
B2ZcxYm5tab0xg70IKgOSPc8S3oH9fGhHhpQeRl5er6wn1aP4UQYEbyVq+cKTeP3
T0dX6yIgc6ABg58193pZv+pZ8hoEgigxyFo6ByXaUo16OFa+Y329PAegITrGU0Qv
457QYUEh7HFAj/1HNSzJ0jiIrI9RHAdryChW1EpS3qvDLeyp5NmLXXDJgkpLRSZR
QM5FpS2TaKpKYRVkqa1Uq2ynSoAH8zlY007nJLQdFTHUGVyAYsKP2GK48Gb8B+hk
pNJQ46QQNM82s8WSwPOrlmAECNboMTrEph5xDeLs+4sjmDTVjNlpHvjOswCyoIpn
HAaezP2y92zHya6X+fDOid+OOOgMGQjosqA+AvUGm6eygCQKUago+8I2shf9Mh+Z
1Z2ZXCO5mn+rTWk5HPTTVIllq1JyrFDq6xSi4sEAe+Wd84YRKj2wsA+EB9RX69ac
H0K8DjHo/aD0gzYFPYdRVh5Svh6RxcVN/scx1bcLVZ77SHG7kRnccF9RKvcDe4CH
edpfUXqyUTtS76zvBhKWRfTBEmtsfXLAxy4ns+vq8//Q48we4gEm4vs9sc2oHIoh
9bS8+OhU5qtuppsvVD9HSwLY2Z0vTFb1lzZB+5sZAtTw5143GrIUcDydjFG0iCEa
sMnYlnkXv47bHeSZqTrahZI0O+ipUbPyANBGf8GYJwMVdpop9VJpzbpXGx6EA15a
iknINHqzfa/e0+rs21ESakofTJeK48HqSgwFBPoAxmqx/9/g+38loV3DYJn/wIfm
AZhKgWWRInfGZfW8fm+pDQjmimyRjEKFvptf+r45NgGroDrFy5s7uF5Z9He1pExN
htweywLit8lIGbm1ZYmfT+j45FAJd60eQiCGbBGA0Yx2lCUO51QBOjH+nz8AhN7G
Fpt9vHgWvYSUow9Qu0+jJ0t/mwruA143VvlZiUINq0LCHl10YHRPw3We6MEFkUY9
hLKWIjpJS6NQaUOiBEADU9Ce7dryWQKZ6qIasWGhP14EciYKKuIISxO5fzqLgZIe
eKPP0h1GqqNRY3f2pVpgqtTKTcM4tKuYud/hOQN+mJIeO6hxVpcpDXKbf2lp3UcU
kwgeCWlc2DFhHFPTtNVAU52R+zKXJLXSXwVLK9TnZIyJCA0Oa8ntn27exaE59H1N
N9vI+qFJQjnWsWy5dDbxIqNo/5D+ZHrxhbuooWiRtjqnZ0U+HFKnhVP25F/XGRvW
U22VNaOch8VGyn+8dW97l+fYTEhQJenXE3G59HCFROgY+udh4vKoY22qqwrkcLf6
T89GVVAaREoe+BGqGE45wfYex2ogsGK64Y3KPNR4ssgnBnZMx/rU3p5wVfi1Uozu
0cSXx+txTfqvhaJsBljrJuuhM6/hLFRAobgwnT0AP+26XgZb6NeCnGdO5+OAE9Kt
ubnGhsNhqIbIAA/N76juUhtyDLiYoFXs7U9L0xSalZhxGsrA69RLMpamw3lbCcvK
j71qB8K4HSBLYjK8UWvv7kIhZEiZxhQcE6mwy+LhD1tQvnnzovfodLjIU2KYiAhF
4evWQaIpPtMOPwO15qg2FvyZ2TLbLMOtLh0lcN9lWFNke3uVfi9sVxMPUnBUsURa
4xRBr70deqzQoG+RWVvpPYF92GehlcA2gc8UNJKNNDHBuAdf0Yz1SLwUCzN3d/b2
i4EBtC9Ds0ZwpdckAaLCjZg1AwCxz2lnXAD/7C+w1/T8r6HsbWeM49yh1jCRcKCx
3DgHDMAHCg2LBEu/x6G9cLc6uADy6VobAtc3KB3WD4vjAmwDI7dCLs77ygW/uo0O
lZAYSR70IY0i7T6XWtg3DBwhPhWjhmXBecPdyqDoKue3zbKc9jQ+f85cVW7IunbH
PUgEDJgTUrQX5u+rOrx+8XOoShyBu8dH98xCctVhhZkL2VdaBQzf/D5uMUzRNnJV
PeSNYsLX1N+FidijSi2svt+EaLjFJ7/eqGlA8fxQSvH12URE/jaUt390O7wkAHPy
2Z/wFvpvASJMzTJOQhMvLSnyV0rI5A+D3B9o0zGr05wfGKe2XAYgBsuNl/h2TQNe
e0JCUSNMQubzRxSnWsVPqUneU+vkqbfPuUC74Rrk6M7VwOFdxHBLdlP1+2eNMpd3
RGOJ23290Xv6uS/yGUOwFwZe0UTU1b2ErcMa9w+Koo66296/qRnsz0pWjzSjsPuy
O1m4QcuStF0KYcs5lEorUul4yT53qiUvY6AepCJwEsk1G0jS2eVUV7pp5Jgh2/+w
RRhjAroX/B/071YgKfofpwOIrolr8J+MnCthQAFygbv5jxVpsd0DfUowlXsnaEbq
HNYuKxIm4iE74khUrlh8CHeyb9I9hKoYgNRkcT7o3Zq9H3EOWKG53ddl/9oXN3pG
76GWG28tCPJcf0M6e+rF30RBUVmEIIX5fbJG15R2JAAcEeHmZVlva0+IEL0l30EH
AzJU0JsNQP2y1vEQYJw4Yj7x0myerVtfbr7bn5MHp/y4EbmaWeGPt0sPwjy3jCyH
aHEF5v7TYUEy4eQmDGHz75tuHz6P1EChQWXMga8NJsC7FKtyR3T9xKHACMbGkJyf
lD6RDZbnOuwxwSv6dU+XmmX68KpDCr9d/tRGt44RGsD1o7Oq+lMca22YU98EiSNn
n1QA+YOY3aEIb0zcAdaMFboBP27UplFpTcsj+akTkuJjL70KTrgDZCVPupnHJYUM
9G1FOcBfZ4nNYqvXoeynnnf92fXZQuyzlQ6Msp1x2O7jTSm4UDe8zWNV+hRw6zEL
Z1e6U5iRyll5D2si9Jzpy1ZP7oisK/UyEqea/m85MbR3c4eKUeQQmIugzQ78EWYw
AmZAFlrVspS4YyJtxJt/60gxXgA9yybsd3qPqiINOp9VMWjhGamI/duKh5SGvxnx
UAfQ5Arz+uo0NjuA8GV8XycPvc3ykKoCZ57SLdNoYofA730cB5xUN77pcy7M/Uw+
794EVNChFeJMMai/zoRAqCP33UYdZxL0+TURcnVUcOEsezuYCqIsy+dnLKwPTB1f
YN8WTzUcF9HF2YOx9cBCTmoglyhPqBPfMpMMdJuFoNzg6djgGRtq3MdTE8IK2k/2
n+r6q6qCRNGUgzeRK2IxzivT5Ubjz7T+EX4BctMBUVh6VAhs9qreOqPYRb7zByX8
AbROXFn5cOxm+dyQ3ds2jy0rzk4E+TJO/JzScikyHMRyk36AakL1+gr6UfdRK3V9
VFrkOqiFm4AJxrcdYM7CppWKAylTDkCaklkAVaqMvfnQoocEgGsotEZc1Za6rDrb
f3IfD4R7vgjD5zjhI612EidUxirQhJB7j8NmyZaw1EzSI1f5QdYR0GZ9zX5pBrDD
Vf/rWR1r4jT5d6VrvXl0r4cRWx0nKAnf6hrKbpWJVIIGVGVdNFX/7acxen2pLQ2m
5KJ3c58WXay7G5NJEgZ32UL4QeFrnE5V2/2ZbzzBxUz+9EUaaG1EADUyuSpoJnGI
mYV68LZUoth2tx23+qavF7KA8YHJ1lTplvi3roDI0bOwTnra/PgifZRvH8DIKJuj
H08mEloU/AdcJTGzvkgAB+GHw9dUgTUGjRBo+BueYj5KX/a5PI7KbCMWh2PK+1ym
vdQbhk9XSKU7SiRcBEzGKrCLBGRoi7+HxROi7UpJJ2ALnWoJQ6E2bCQXCXSS1FmQ
FOKHyMttJawDautH9SfoNCx0DUDh7R76I6ASbE4qyfws43ACgAgfYy40YrbnNyR2
mTz08Nq+aL20ZvkqmnhRkIUqaYaSk81f1jgSuOWop8qtNu8OduQIZ/c9Qth8dknj
OcsT/QvDMBY3WIC7MTf2YLKDJuWhQXZH4oYF4bfrZPJVJMO/AJOwLB8DdspoK75k
Khm2zFzp4OgGJdUOQ5kvn+kxT1r+BXDEK6MgCke/Ss9ZEY4XfeGCTASMkuC8lHQL
j25xlPylkkiXjJm2B0sBfLuumgHzKrVQ6aFZHgg8okPlnTM/EQdji60bfnW6Q+0z
Ace7HiWauvleN0ldZYtQ2WAHEvdNeP4DkxpAQPH9ENDPPm5Stkgc7Z/JaEkW53BX
iUg5+7SpBd1oqLMqHEYdKcdNLC6yzJS+tgL1z65oXkLdtE9uz+Y9g5qQPnoZPS4P
MMfRlAS+vduNTuGTkJgJuD17ZYb2e2Qj3EKjLSO5ozBWVY9t9S2cGjJ235igzDo0
uiAkZadBq+BVrn5lVwrRPPkOWLvl0022vrDgb1nbZhBQJKPQ2lWJPxA+ZE2mU2t4
hqiT8fymPE/fSCvwpcWCxP93LkOdraZnsQgeyJyerrFZU4fgNr4ftIiJLk45EM5Z
mkuRH/gOloWAT6FeHvmsl/ZbT0cgJYh4tkwDzv4ECPfn9Z5yywqTcnIYdd/exdWS
zEL8UnJ+GXGXTRHcjFUiQGdHaJCcwnkQCcSNVzfUTQV5X5gTkEuKwVRJ5D/+6vOP
LjZTxBW5tr0iKPYtySRS7AKLQyDJfO3wVHjPnI8A365wMCnAWEIAzSUedSN5LVNu
k5hRFBicQCifT/g4dBjvVkwlFGcyewL3xfsRRIxiV5NGRKUInFzCEHsjwQOgxrQO
1I6iB+l5HhK8xTJh5JbKZJjSZAElheD6iF87ju+mRi5J070qu/aJWnUlHlt+Morn
TH7J2u69wZAXgXgNWbat1YASazHLpsoSCdSqsG6z6PD7IelqRan9ilSfb9pQix0q
iCW84gmdX9ThAhawvOTZLpWwT/QPRiMIzv5Hh0CwBHCyOerTt5luwxbBlpqA1syX
XFJMv9YMxdEP2mztwAxmJDfyoVlUkHtrHwBPQGH1zEJP8/BkLLtSdsF1ajOTrAPO
U4yZOSY6OXO6vca2sfqf+H/dN0XxCBKvPE7CML+siuHQBWKWwTaFIFGdk6pyacCp
VmyYhaCa1A2xVIWjcerYatZ1AGN0zPaMl6qg7tzbeJWJwqLDZcFUk0nMi+AaxoTy
SdMSmfqFQ7fEpI0OCa+GLPQrPAqKF6+wqEYPBOUZY1tEfqN7+8UVrGN7QRhbizDt
YpMg6vIP6PxWW1ziWBE4pYTDOUrfbfCoMvVyQFsnIGozS1dz2vqkv4BD7ePDCJuH
oEbzdqzwbucpJMg+CtnNl8nyX0vILAe1O0pSFCB7xrBRtDxEXbf+4NvJM/na+ZnL
X0aXCIIuF4m3Qqi06D+03Qj8jpbujdczkVZqCacTAczcAzQHhYJ6izXfrzyX+2Dt
0gueuZCIES9VRHItjUU1d9i+yPw6OoxamznxwEIcviw0aNYtjNyhpHr/i9z1EWMg
lKRWb2FbMU/StrKsZ/wf/17CNeMJlAu1lUl+GcEheAEKRhvjkZt6Y1PJrTihTgz+
/nYmU3BemY3OSCmQSA1yWGSqIChGENeWH0VypqnC2QH44sDrB3RfFKJNOaZpW6ea
6fUUSihPw+gI8mIxSoKONmVzYH+Pf0LfesvJRFxHku0hH6oznUKCn40xFZNYItJn
Q0kWe1ytzZ0s/Jq5e2b6HsucVntWYkwMPq8mh4vuCQvn/lL5ZEuMOopNEOwjQ7rV
zURMF746/aSD9c91AA2EoGBiUJZRfLNBDqotulvYreQK/gAyt/yV7/RrK4eCNNl9
d9HoNNgYJo03/uaHalJZNYRhFAJhx7xjcYcRH8pmYql/1YV4A0IUPrWbzKJz1pZN
B0S6czpGy+VLbMZ88gczqz/RZcUCLqPSX0/awxAv4AlfMnOjYgQjod3PwLhrisG5
w2BVNP4HEZt21cH5eT/Tfs9JLCFQE1okzBOmoNAm2Wl8c5WFxGLO/qVMawPGExUk
cM+OZJLObAR7Af2D2xsVKcaJ0BC/0Dod9DMjw4UQP3GZLQt4Sk5hf7kA7Yn/DwWg
dG7fNrfbZVhiDS57a7LrvYw9tvZuaVQCcGAK9dthz8rIqez/nd3yZVfEsp0Z5DyY
jKAHwvcgu0AVsyBQNmmTrzQj5DCDILvzBo0FsMOvkkeTyc1ik60FYdcdPrqPuL/w
ObezH0pvxtpgDbBSo55ufV1OgfNAdWXhjEX7p83OCptBox72F0SL21dFb+uyoWHj
zZTu4C05WXkGJL/pWZ40lwHYKaMQEulPe3wmGy/oa6nAH9AESfzXnkRamGGtIhUZ
1C0ru8tMjmOfQmIt1uMMCiFZES8+wZGwKRyFhagyB39tMDbTyf/kaV2sqXsYplOW
NALfHjkZ8J+nZSv2xU+rZp7urUvyW+S4MDorN10Gy0ErUyQofdNjc8KCOS71ECrx
rfdup+twE6JWyb9IbSlCxYa9RyVDbQTQMZlihnRqeF2R0oWd+EgjD2FbE2Ih71T5
Of1vWHYVf+i7lZhKPbKjZ6RNdOxL1h3R3nz3bX1BCBJCNaNhLfTXpceBA6un2zVj
YtiddEP20/4ToSpnAXYFI7qfjI5du3XNSazkZlTkxBc063oX1hP6Mv9ZkvMQ2YZo
zvv6elOVRCkbifKff9tdMFsRn9sArfQkD6tRfYwGilcPrr2IAxTWE+5nMEfFh1cI
zUMAQXyk3yGsi49pzatht1XFxuojhBHoJIe7/9ufgHb9eHGPyfnOk4eH+yfj+0vl
of85r2Wt7PnYiMYZILWHnnhnWkgWSusRVqhFxkYNcNwzic52xMS4kMk2RwNzCcSa
KFFRm+v/9/Bl7MAC+KWc3UYw73t0iF/R92AzKb/FQ0qHW+l+HgiaygstHzD1Mwhm
oTsQw7fnslF5xQKGWJzOgTnjJ8j6IYISfIraVfihJNmcaDHy/EUGCkwhTymX+8jV
Oss8qqM7QBLHN9e0W/LKS8pxUEALDBR3pH9W7J7AMcMHn2AqOqDjHe+8FPveliSt
gV3JMndUuT/Khj1HzqUT9ty+VVwXB+BzPuTQudRDvlMtbSMZ+X/LGznQ+QWSaFIJ
6mqqysjcp58V8is/nBza/DoZDmqvGIDLH5pMIRDdPOFAfDPy8sDypaYYGPGVlnT7
BLdjlbVCv4YUyqjRix1i+/rkYG49sadyLc7NYlrP4WXl8q/MGRLunwh/lunQ6adr
RqA4uDP6MidfAmzquhEuv3MKsE8LRZmfOJm3cq1a/KtbTcFeOA3T7iS19auIIq1N
zvr4HxOkJm11YRqoH0Ykj/Mm2MNPJMHeT1/Xdn5/koD+EU7TTH5SGMF5LThTaSDB
NrMJ4uNcCisqdpEU18refSpttvncyR0xYi4ZQa1px37uEfqPqSqkiuvzCK6XiygZ
e4jZYLYG8ftpVaO+M9GNt5xlx7ramrzuQha3LIpxhdk1aVBK327uTwuiF2Jt2HuY
NPUTsxVHV/BZwspLSfd2ynXFdtp6hNoPllnWHfhMBOn6LtB8fNyTOB/bWvW05/hE
BTN5xqaXcTKeWdz6viTkNfg7HBNtL5JbM1K9wYQTSmOQiriobTiJk2V0BEmiD1Om
oCRBxwvaA/zK9G8ZxDOCldoXlwfP90eUZjb2k57W4G9F/e0YjYEb77/T8Sr0xvX6
Sq9Cm4w8IM2s1nbSmEQ+5d0MbJqgjisoROc0qm02JmDWKlyjHv1smkSZg49WCzQP
oNWIIkHmOzySgnBqh+Vifwi5bfrEJgt4m7Dw33CbBj515ABYGF5AcJMcEUI9HR67
/hoVJ4H3ByQWwQrPUz5WP1rNBGHebG7QMmmPmZ6jZwH8EQM/MwYA1GvZq4RJHlAe
vTau8yWBkHUIkvVF186j6yKWSTSAGfwStTXkxuedgRvDY+RiMN5ecj/SiajaQFzQ
TDKpiP40tqdRkLVY7AzAIgL2xNEAHfFaZ88nAd2P9i8u3GcnX816hLC0F1F+6+jf
y/sFqqc0NnKxlhAgccTJG9D72565Y7NZmH6wFZIlj1fzzZmJ/ZGuLXJwh0TvseQm
ONyncX3G00qyogJRL7qz7k3I9EE8cUEcuE4juCCXxJSGU0CS9wIy2n4JmdaIrd8I
XzSP0hPqJLG7tTDi/UEOICDUdpkLECVXKNu31d6yM8b4vE48FGVfhiMSw5ud0wRF
njK5cUR1optvhaY/YKrt413PO/r3FaASzX6lbSNOx9baT3bKfOoQwb+sdK8bOO64
UlvPKSC2gnEHgoRaaa6mc7uJ7GhQx7mmFsjO0vagVsmgt6Wbo42i7r4+x0SXB0Ez
kZn6K+unUSiDZMMyvdobsBvvc3BENOzZrBHYme+PAmzJeZKJl2OYOjvexASdpyda
7DS32SBN5RQ5lpfG3VcqdVe/V/pTk5175vk1cJYLnAqkizHKgRgeabvW4NHxLBQo
DrE+niLTUjc6kgWk9iR62uSz9Bk7v5b5UyrMggq5sDGVPkUNpmIkSnCRbi+fRqxH
46NRNQQeFQL9JJXlJFALkCCmnq9lCVzvjeUvLbKsS5BjZLBiRcRkokOEG6VanB8x
qsEsV6e3B4vhbjZKY3r/rt3JzGraczepCOWpyGzbzuK65GITETnotaxkPMMLgcQR
hPNVme9G0KpcBglJc5Bdy4Yyku0p1WJLthmi46fC3PlrnFUfIp//3IqNyowSV3bY
fdNTn9/zGsCS17VaWalNmzRN6wmDUcFYaMIqs/uifdpq9Nwj2FODSE0IPvac4fv6
mPrKwicdtKlgXzN5NQDsO+gmZ+Kw35a9Sk3pEBp5+Co9CAlcCgwz3QfCxrf3vcsC
ajbtCkv7Gjis47TivSEuV8Uu6tn3rJYze++yMplln9Rg6iOtJPzIlyaJnC1D6/Cl
lOkJqMB2DDAdMKcSFAZ6zoZWP/bOkeL/GI2+rxfsdMNQr2geQ08uHZk4tnOLSObi
jkb1MklqHx79mIrKVVGL6DHD9XWv79gHwoXsHY3w8TuXZAVRBlLcUjP2kYrc66Tm
t7Z10ghaqC4ucG/rQYQMwkRrcyXzBKrdeQc+N8379MeXZb+YMzwYDfxp5UYrmssS
FuezJjnTGuOxqQiRp+kA1b1m+Wqej9Dh3pPrci9diNHLwsx1QC3ZDfVV6sCRkw28
QhX186S5TBZpr9NsjihWxLOIPkRp+1dSnl3KYzGHRWwyLRHDcl4YgEbjvgAfNLPm
a48QWidg6RjpEpDFHNbuVHdJRPR6AWaQTItYRzluTwww2xlEwExBKsYID7dvns1G
xeYciTV6duKC0fe6i3tJTyvkUaGDVNTCLcQXgPVj7YAr1aiPB4aG49U4M2XdQgBD
2s1G4b0Nfa6sJkp1y+MPeCRD2f0ZwrNREuyCjt9+ObEu8cavxdM8i8jIKF9PhkQ7
bH8EtN9mFlp5WunouVQt+wgG5DHXve7JofPDGIMwCKt8aZ7mV4eH/Wf2gAA+jGgP
i4J/55ZSvqJtdDQKoNaqVLmyeHwBW2XZI71Q6nJcynb/x9V9xBfOHQrfVb7glgGJ
jiPhoQ3Ce7RkyY1yIohF+fQT3XiUjeRJkhb/8Pbd49sEgBQ/Y7oHsYl+p5IQ5GyW
Fc3J5k3tAuHCIueB2PaSJ3Ihg190GLjI5FhGYpmAKqMwiN8wcGxy9y2xr20BvYeA
HSzpQwXzd+Zs8RYnFW2vtMGAoeeizYF9J8SzSBsW5vbEh5eVMFlpZNKluG7C73pt
ARjEDMgEiIXw8yNcLhGepplooVbUbre7d3B3fUvGlKiSYih/7qYaDQdobKY5k47B
gakSMxjgZodwBHoaXfayXdzOW9gIncdnW+Y9w04DtfhHea+sM6C8z/BCwy1FRHt8
5z5fquo1em5zL6VJHPUUOfNL4vNUOSyAp2cIKJ0aBiyFLwsdAuUYQgnPJQqLs9qv
F66XLXYH+30ixYlr3f6MfhNy0lc03UH59mp2b2CEwqdsS3nHPipYCjSRhzjwTxbj
GUwS22zJCaHMMRmVcgb2Is7eigzOF8Q8+60iWuBYddEdxFd55JF6iUYq1YtJnMZF
JV2C2rneoXozV272/a72DE5tDkxOOVz0AQP0aO/nY/alFyI0C2fRIPxfdzAevJmk
0YPZCWYKxaD0v4Y8ZQDiEqigdAw4MYiaQV5t8RqqrzSo0ley3fbFinA1YPpZa63M
2s09L2L9dHzno7plddHDGzRoYmLPTsdcpV24+CdsLHuqkX7BhUzSazuXegYLo2HU
5fUVigs/IAcxEYUkTYQwo4HzgRoOJ5xLzcszx6wLmNqJ9uBkImq1Y892fDAtKoP3
q3zitYZDKrWZQV/I16a5rfmOOxM1WjBUDXyUkBJMmEDkjmZVG1grBRVN80rPept/
2gCp61RiHQjHIJgeV5Rt/yw2h4kBODP6LSpAjbnbLnPsvts0oSa9MuuH8ghPRhgE
B3Rr2Cp8k8Xvhf3W/XvedOB9qf++KBupY8o8VRAvZS8qGwvOzhVSoiwaDDapv28K
sq8Dle1U5737CtR9I6DEcIrNRk74/54nehL3Bn9/g9qPU5tb5u53VFH58R9LrcvD
EaWmyZPwpP30kGQ7Ia2wHHLsLRJvqZn4/6N4OK5VQMtU9AKU0HRYleQK1wNp/K3U
CGafLj+xW0TL5wBI2Ilk4XNMVlXcLs3SxOwG86Jf8aHjQ96yswGDXixGO+hG5k+n
8pzxVRnjmXdabaHzeSbqdtkiExv3fcuG3bt4qUg3Ut45I6cC8fRAtdbxKlc6NAyj
QqFyhqaqchBd4OxruytBZmensM01fyWbqkkCCYOjT7x4sSTg38vr7WVj1M6vAt+X
yEnUWXH/xaQZNEth9sX7sBwJxzvnPx+4ajfgBoSAIlHSsEIU2hTu0YYS2o5rw6Qr
l24GBE+0F7C9ZHHb2oQhA31j1Swkkz3w6hgRyAbvtZD9EewzCj+AOG64mwNuhv6L
3i8vwQyjZlypEDwDuiKFcf0WBOa2tovXWOxiMeXbgBYndF97wbkEn0J2V6cya9qD
HBnE846M7OlQd1/kPgzxxcpPAq6lPppw4OqrQvVZj6i2GOCQTXrR3lHcebNXJF68
RwABLV1ud4vhaemHECmUNSOBeaHCRxbeA4SZmJtOR7Qh6wB8Ru9t7NELCEOg3R15
H1oe+og2uTo3WSOdOGk3K0uQp+MJrW1A4Zgo7LBbxdrOvS5Upyb3WC61XL/JAWdC
FSA3GI0pxN10jq1pzp6yfvenUqrNp+gT74AxwhLuF2ynBld231lII9Kh2zPmOm9s
x2Gx22Xp4wWgXessS7Yuhbu4jC9CfgvsPdH6E0sDnjnGhJ2H/KZgdc2ep39AWKxR
m/3w+jH1RrXGlJni62J3eCgHlA4XXRxLH1nr5anPUQNIh61ZdxU4ki1BGEcxCLqv
KuWF+V7aJxTvogv+YnNeI4KC53wHUwel42i+L2s9Tns6jDbCGPfXvQXHmNs0FHN6
RX+jtZ7sW4uoBKrEaNX3k4gVLa/D9Mb1W+nYtH15O82tlc2I4Dpq9YFxG9G8/viI
CVz++1rbhQQ/03pK6baGRkRdjkupLH+40hqF7ilHHs9+ihFywfye03U9N/vrfD66
RHaMDzhN6BAJSIIxMIYB4wj5iRqYtONIbiap5S302Kk7kDOlZ19+vSprRH3DKWuw
+GfoXvcuRCV4cRLZzmWGI93b51efILpPFdviayECt8G7uAyoQI7nSCRrDDX4P1vS
1Vf/ZdFS/WXreTioznp92SvE4sxUnn8dGI5fJe191r/FS7/qbskmRdiPO9fuqcAz
oXPZdOHhALrFaQnKi/FP81fzC/nue9Z8wmwlIg2n1CF6RyyWONpjT/nUBIlEak0/
GkkeT2zh0bJUo3X9+sjHdYGr0PXu/GeZ/r7Yh2qt3/CReyHNDW7ErauI6lv0fSkL
xDq9qJAO3Dog5IwbYQv698zkjQAnENksksOhT5O9r1BbgYig8gX91yIsHAIIRrIw
k/dGA8Gk6dxPJRIGl28yvV0v9WGFWuHibwO3AUGMVJJ/RoNG2pwxMe2FzsZhg271
5U1DMpSfj6A+oNiGMm2Fh7IDq78CHpAu8gqZidBexd+hCzf1BgI2+ySagD6CEIYQ
Dkd+28Psf4Y6V4cGt6ZEcne1nIll9Lv+szC/GCqLEbuaE1paW/wdSyEn2NSkqfAo
fcOhcfauvAifvMcFalai51UZuVY5Uyi/orQl1EgZSM2eG6kBSm+V1Z1fgWCWW03s
q00X7kTQtE5S5Q1qfNbMxATWGV9pzCfDzfokaK9HXrmWn1NM/k96w5lbgKnqc4ik
MumNn36Svobv1a1izTTvsjeyma0rMkk1L4B1nQ/zZIDQ6jCLEZwzboG9xYcs3jTL
+dW0z2kfcgdri2Acfbo5nIgViORRktcCXfafLrXRTk2Get1dOdH8+ym4smktQY+7
BNWNR9GT3MUGXGXAW2Y2TvK8MSRSyWr9kF2pwukeT65mzU5GRNGvR4W0PybtKfp/
RVmjO00kKt6UrtbU9oTVLMgXCCmXTA78MgU9phvgD9gWKE1r6B+33lHIkwlCFWXV
pvmaZWgFbejng7Zey6Y7GtvsPhkLRzUVsgxTLswlzk7wB9KKu6EGUCTmyw4fPqhU
jvKpwI+agGtaZL7Df6c56nVXELJswtbEKj6QTSoiYaQnpC31RgdNTEBAmRPKLcJS
jOGtp1dlLvuhjuFkUiCoLyzthSaeo5BljnVBrAA8azkhc+GXTk2G2xS48ERWsbMY
6rcVPRc0yqg3SQ+epJNbaHIKt/m5E0394v+P+cPj2J6sXWt26SoyzvN9TafGMmOE
ZSOL4ZI5Z0mr7d6f/UIjvIPJ5AxoZs/sm6CcqwHuJ9y6lqUMiIGz0Lm0GFmKimWV
hviWhKHIfUYb5RcQcPaKwUGWMHoPR1Hx9B2kC5XeEiglHpAjLDDL0fMV+eapt+gr
+FBeAnZWVHFRRjRlTj4aGx03rpc/WatZPhl3A2kY9vuBLVD3TqPcxNyvxfgBQJ7P
SbMMcZYKZhASn5+YBwUeJaZkSroAC8YBsTxI7VdsQseVcEm4HKrXq1hwI4zxUD41
Uk/E3uJBXGcOXQI8srRFcirbnzzbdVf1j6NroyrOwY84h5wUf+EeU+euvStJpilC
vLlnCUrCFZbcUdpcBUJsgDxsrJFKBCiaqswMbIuoH/BuMtSNL18Kt3lwps2g94Vc
Gj23zeNFAR4GHPC2UhtSc6OH3Uc3/MkL0LFHtyE4pt10acSoQQL9+tfWcH/hPjw3
xG+0RViPSqkebPNZbsnIZOVh/COcnB017xTAvLaiNZOQUKE0QM6jsko3vpZL1uiC
gwleQTd76IeAOCIUpc5Iop1lsCz9D5umrxgLHf8RuAwN+buSeVNfdWOcBFp10VCw
k8mVLArPkiUuEpZcc0zxvu6HXt10/AB32GFARQqaZBgOxPC70zqez4Rs8TXVYtdM
0sshWpsMneZyRJ5adyeG/qjibbegv6ceI1eH8OBqV4KlFRzfWCaqIQJdC0lyLb+i
o6o4A6l0C/T1jokZTXnWwD+u8atpB9JQ559Zozi2MHwMfNEVSDzSkUqSP9r3dywA
ngoWKAunEU7wksUlVm7kUcdxO9kdMg6x5GNLkkRwaZsbspVSKN4H6UfABclKJeSl
1peGWbR3zpOBQLUq9npahuMsiIomkBNcWNI8c6z+5w46cAANMDm2hx/wb03WezcX
fRhS5Q+6pRu1RTz3AFMILSVYcfCNm0+WTukmYD6VUEZX9i22czegVXs8WeNs2ClA
S2XdxTJ8VPLa6fv6EiEvqEbN5I/dOL/xAposOW16Z0x2DPpPGnTD5VIOJ2/mhWMD
0iCqH/W5HQ63UVbogHDrwLlokAIx7WTLII/OyeK8Es267V6GFy2bhu5jxvKUShGW
+OhR8PtqhDjQLq5m5Eh2X4dn41AA+1+MOybYJwNZl7Vy3eJXU2INgmRQUcWzlxgG
NDk3VygiK244Qho7T5LDSmazIRHoz2e12+UX2KZY2VAKGLHrUjQTrcYI1YkyME45
YC3LVZrMfCtd81uj1znLR5fpw3V0hfeX3qTrVWNMn1gqRZRICfrd7lPQ2iHf7nOC
ennk94E8YrGEkIG0VLrnnKGQa6bZK+OUp/48Lmo4qb6JGVzz3Ci6+M6IhXVVGCPb
scpfdhX3ohX/xebjBniKXpLShCW9jZVznDa0TKOE471E6Vxhd6o5CfWNPU/5er3W
DOf+obntFQy1AmTATc1I8isLQCoxYXH0ryZTr7VcR4Ap5Chmt3ajW+1rx0l4q49O
fXsyfgyXVWwyrEBuItmrUPYaeaF9vdjYBjdQah+6WmF83MCNggPSBuZUv17wAomr
TU5hQhjOkF4UaNAz2eMyDEdXG1d6HlUYINXD5U6Dl1JT+ei8A13d3wSyHzVUyWgw
GQ1y/j+avhhbgVokz7M5+Z8sgWJuqIy2u+235SXf95rLZypa0szGCRLIycbaYGeh
0hkQUbTKSgMMA6EOwPC2VB8lf+tCTjLHWgenx7gztuHogqTRu7Mem/UOph9lGasq
Tnyh/ch/wnZbnjF3OJuL94va8XG+f56Hoir/PtmF0CZotLCzFP+9wY6We1KXoNxz
BRUb3HoUfe6VWylavWF7Km9kxW+fmHKmLea5ZN+U3zjsNoOCpAEFMP3hayLiOMFW
YYEV57wBHKVcF9h9ABZV+F+/pCOHEGYY7rF9OHfR/vr2/JvbdECB/M9hZUTzp9Al
Wsy9W31Wt2nILkN8Z5SQVswgyttatbfBGbaanTIY2/4Vf8MxJBNaZyGqRRNLwmzV
bgFp7+xNnrB+2xNZy3S2mJI4VaYMmE1ygZWmsYeNQEvojpiCwQ0jMI67MFdnVa9M
eaacZ7nJcdO6D/vT6W5rUStu40big+R1XS3vCPycsW79AfzdiE6Uf6lpPexTNO8V
C244uQKQhwRe/OPWsPG4oWh7uXU1cYvhvTI4WrXWXJR7LRLu196onJ7kJDqSi1E1
Wd28HCMOUuzkuWeyhPv3do0DSGlM9h/THu+UZ9R81EbmjHcbmHBe69FuSKvtkSke
s3DPY5Ip9I/RsCm7vQroqr1eXcEg9AtEG9mA6gZU3LMqpu1yA5VVP7lK6A1aXQ0V
FUjC9XVCa5kR+0a7ryl2FfmdQN9PWFTT9WT6hopTCj48mDzRCGZOTOQ3QW4nO+Z/
P7JS3P5UTzlsy/Ci3qKjx8rGgSDiubTsIEuT1TL++lnQ4sPW43/jbel1pedtJHPm
bzJj5LK6c6s/qA8wXGnBnrkowRqL9/mJnCLybSt3R5OCU5VL+ZdWyQuK998lC+K6
8u/ja9xO0M3KxNayjWpaW9FZ8TIJdWoRpxIPHVDvniLDYgM4+VGvJaJoBOmtLfKO
ujF+CL9+4KP66ZiTUn6g0Is3lSPtqy0RPDQrESlGRoKHdHAAkSQZez2BWzrG0BBf
lxdh2QvM+oqLlfu9i4NKwrHU9TBq3gZVzoGT/GRQIZWbiXpAv6G8A3v03Nw42vUo
TaCstQTS04B8Klf+oPukvkxgrU+utwTS6Y6f/4tOQnebwx5utANXZl+ojUGbx5kD
+IZaDkWEQyp6KaFskR+Pt/KzfShYVg4wqt/p8hD7HVlDhI7JGebmtrrSlDtJ9H5g
0ENE5aVM8WRlmGNdcMHAiXjQwiLjBi816jAT1L2hkmZuaFynBKiE1hXHRwnYM0G1
htG6nr+0C7CzmHnWbAQPmO20Kh0nAw7sCx/Mt+t0w8pE/y7ewVeN8pmv6D9h1OKo
AS3sazBfG6yV6if9NVpRcJusynNmKPFKgDbi5tAae37ACOIJct6TywYA7UtWkgTE
gxALwhJWy5llVoo7SXCRAJDP1MxJxa2xmldZlhPyibhgpk21WYYNgirzQQEhc+QH
Aj8meWDASny6aOZ37/OMns/YFcXif1R4HXlnCvxVMrNDInrsmIsMKQNE2Kh7Vw1E
jhDVzHKXuI6GQtFJqWaEDrguM2UxUkXRbIqGyAZcYtGEc3blepf2gk6w7ZH9Z6tw
TDfW8/3b6Fl8mR+6CcsrtByIASMGHXevE4wJNZQNmI7Gq2qKM/KNlwRE/C/LBxnW
SQlAE0nbOAt59ibLe28CmiBEv8DCcGgGBIwq1KvxrY9NPlgLjY/+7ukf+awu+Epf
VZ4YiVCl8ij4Lo5wOxZP/PMEP491gbBnA2vlfNTXwE0rt6D33ucl9vY4V6IvPw5D
C7lp6T49TuAEs8VegLvENfnGfhQTBrbqwztURQnJJZzqNBbZbUkbcv0/BF1hzNOj
rsiDYn+XGejGg7Kq/ETmYLt/J+ZwK309/n/clVxKJcu1x8ht0+I86Wj3bg5B+goB
J5b4aHmLvZWehSPq3CLPK/D/qdSGFqrs/h4u1wleDoPo0ViDowkEfcKrUN21ej0j
c+7xpw2CZWI8m8CjOXr49A2HU3Acdn6CYLBxyCcbTzu+GxvwM5AKBFdXvZzw2sdh
cD0NG6fPt9c92NpyHbaw/W4JHm4ltJ9yBnRGg8/yFz8tzSU2HnRTiYm5DYQdwp4B
o6+LkW/xR+9z5uAZXIth8nQDXGx0Z5yHiUZbQqXarBlnaxX4LfXRxoxYv342uNX0
braPH1CSImk7aHGqIw5SNfFNB/Kycykxi6efU8HJN9SSZMTAc9/jMqtJuB5cynMy
ZWLFE3ELC5lussmtrtO9DsnqhUii9+7/ZHETMmFB4ePk7L6vWbRkUoqYvlDu+d7F
gP5eOyK0+wOyNscu6QEikvdMvmp4TchA9nI8PnpK2x/1JpAUppmSB9lTdSFnjMtu
MRYV+3RQHhJCwGE6Ml+II4nP0zG1A7eGyvGQpLO1onnBP8vkJIYu16J63brYAZL2
kjajFy/WtUASwGuKLgd/I3OQIZvftt+1889siz7NFarWDTf/qbHHV65qES94uOr0
ouFfq+GkrUOB8Tf3qjdnEMzo9jbbBBDZD0pUwIv0aXXmc93ta+cWripfmTQ19kCq
iResRiTJGluEjcy8bcdSOsKjG5+ryTh5PAF7OjVjrJ8Pg4TrR38AbfsZkOf7X7zL
9GK8w+vlEaqi0bTTHqhQ+vvEkw9sYkJNtXKHOrzGgy6ZFfen9ysDKsyTP48w9XVK
7kyTduh1hmrik/nzI0G6oxD0OVNyn05wQbIbA7IJWgE1ODNxbLTjsX+fKToiBqZo
Zt8N9x5gFFMPVQD/GFhl2ZZzbKznsuXtXEHkJgjjtOJjnGeYtW9czfVKWk4Mm57l
1IINfzYV/kHFCUnA7NC2Ng9EY+zxT42VQZqVt1tMFgPiuXMQ2ipDqO7Zf6xzUIAS
uwh6sPCElIEuOkwk5srE0aWSgeyxmMK8dpKGuuKOnhLxakMRzwY7YBt+Rmg8oLvv
1RyTziGWxcMnM7dmD+/L1LAS1PLApi47nm7vQOE6YSxY6Fpaw39L3urr60XqPmML
hqzVQN+8bQZqCUsG/ZOcl5Ka3yQ76KYeUZob3hOfT8Rl9bWHumwhDwQ0PC88UBE7
ILQOTrolxfwp/3eVxYSHIokJzil9OGHclBG9VOXiufA6bFxjzzBaM4DPr8BrH/6n
D8CCc8tScrE5XwG/+OblNCJdC1SakydW2P0x1KwQcWdT8vHt9F0GmDTmlTW+bkvH
6PGUwcQ+BvCDDleQ2wALUqEix1WOMzfUnNtgCrTtErCs6fe/R595R3ZQLqnrsQYg
eQGXat8T5kLcXPwamBpq9oqUniOJ8jWIySay41xnd3aSlTwB5obQgWPDacafeJ+v
ls7C9Zq8QL2KypsRHi2tEcUj5BDfPFNJnbnAfqnFGk5LT5J9VAEWLUtYnKxVHNkr
ybtxMat9haOBRcc2y12C7zz7oSdrlbW3ozK5uSJo+XeYbSPY8leYp9kkMulCMbZi
U847QP1vkPLf/aWSvww1vrI3VZ7f6QYfz/ZLFSUBYkUFNuaBZnPGdr/OKVRQZ02l
DBRTqcEe0Wbx6F4KknisnKpqL38Btv2Oo1L8DW4rLs68cl+w3VLiLzFsDJx9xczw
jtrE4PQOBAbWYngx3ezT+hwz27X5LfenFqrbY5FgiciNFq4//wOkhecRQuJPT2BM
iHDGThBYYN3SBviJMtTF8ApaBtm/P2++QMCN19dp4nB7ZSvQNyHIfKGdKNFG75DE
ELxjBhWVZL37ah0/E3noc8yPqdLDL90Entzv11F0XLf7qZ+Ha46FxBRdDh2tVPMu
niGETxz8kYsen4CHDJ7narbiQcUM3TtEclVguVE6EKHqqJfeuNC0hstNjZjuX4R7
OOXrHCF5DrZLdQlpMSApeX6BFicCd1e83UVpKfE3jQMw9hfj5Vj7DJp2E9nt9t/q
IBv8SU1ubHufASP2rHMg6Cru0p9NGjqrwnO3DUrmr4AcOUBVcwO1gtp5VGZn3TaX
SjJiIJW/pGe4pv5bnE/qa0bpoplpVGKjoKHQUl8yIvEcpntejXNFsrVDqGq92KVP
7qjeQw8TmtPrulGrdY+yptI2uM+hDFZBC+qV6tgvmP6iMJJS4I+hUcdpLpYQDBd7
ZHoEJviOUwhrqjJnB6zc6ycYa7WIPmD3ADmiltokT4HM0oG3MTaJPfu3NXY1naom
S4HBHRGWJ5AYOqqx3XTA+ylcxUpiPvCRnjNRWA5ET+hf7A+zuBNs3fCaN+v/lcuG
lBD+iSmNDNnA7Me00UMgfMEBenv6qO6aEKlvhJn2ORgh2SZWqmB25k4Ol0Fr9WcH
c4wLAsfBbSFUw5321cGlQg+1eQa6oF0/v7jINj/nmcWq650dia1IuPSal3vPIBxI
K332rCE8VGnNwkTL5GN0Yp5ehO5QKqa90IlDHnUaSz4YTnghMQpStdPnUOxlLaQQ
piyf0iNBfGrvnnmkxnGTB+Zk2F73zNJtjaQGx+hRHh61m0DZ5H6WsClmUCbGsWIy
HPOv1aLBhmbKYjtHcZJhmOxgpxiX+wmmzUHVKbRfhKILCStCEPkWLofFciWgogZ9
/ax2luNqS6M9sJw8xFRivjNlQSCVfzkSdM/7yJjwcVQMoBeaHsqP6Uw+TXWUcx4w
5X4LHw+AoiQIJhvFn3BVSp54GFmNVDlXX3+1ehC4M/y8MRr9riaU1qCyKes6DAIX
rm7ZgobJA7OAe3EoP61tTqGFtNPk2r4OxfPxbIrw/2+8sGenNqlLf7wzHZosIYik
uXMvIP4C5LugMcRLJYOnFthXzga5eLPlhP146S7D/9uJ4eeZk/Jb6rVFiwhy53ER
SozpgxXxgkMrSkwQllg/NfpD5lkRhOHTKH5sERhqdAIAHsksKosCq9g8PLl3wHDq
c7HAncCHpkrO+JlnFh5tt4eVld1uiBDTNxMb+LLVIg1N4EBJ/MzRTMxpCIi1hVLy
UXSUPxHZiFh9bh2GkZll/fmZsIRkgMClTpFhccv46AH+xV3UgAAfgKI0M/kicoCq
sUJVZluy8jkPZaG76EHzMdNwbvBGArKpvdUZOrM8vzchc8cm3vcmxdMN8GV8aGnW
4cw/SDg8e2acXBHBGHrTy9lw6OO20Owa6Og8VHYnCgNUVF8dkM54in1qjkBV5MJN
yUGXbA1ddLDWo6go3wtttqC0QoRX+A15Xqvp66VpOLyDIdDfoAIMjTgQ5MhJjWqA
nZ93Nbb0ZXPxYKnZLC3QTx4/Roel+R1LTAycsVgEN6U7S+uz00jRxaXNi9Xoab05
OTR2AyBzWsTHLpH5bnYUdAnYKRcaN0M82v3DZseWLYei1ivG8Q+obKHfF84mms3Y
sxE0Oqgo9rN/LotwMqvu+Hkjz4Ynw4Tu9DyV73xQAkEJqS1ztCS0CABQtHJFj9Ay
hdyqivjRDxclWpWAL3f4XKpIiAD+eiyFjIw1Z8lVc4GhihRKP6uQun3/3o4z+MqS
znp5YkkcUyZjFnULHdAbWwI3IvfjJ/po47Zvh1d0G2h6kcG+/7n1UBbxOAdIKag3
ZWuucuuVC/U8oKDkIVwkYp+9vVF1oxivA0clBwgRkxAZHNVa0ea+mzrx+sQyAhFn
VsVyYkIdh1fDcEzXM18X0o79378gFUcU7gsAo8wlzOWUcFwJVDvg9RZY8gUdA8M4
POxD4wkzU74mAL/wtGTMyMjNxZYL4qa745zK6+1Cdb9jG2C5I5ZPjD63KaQ7pmw4
vhmH/UxJEQNdfAAOhtm+vTJrqZK5FuxX4txe5kOuIOwaiV0P6qGnkcEpfxxq8IaK
dHODk9dUC3ujDdOzWM+vUySWIehJDs34cmH3dpuNNoI3KvCZtCN8z0jbs0SiFnzn
3AvWBT2D+OCZmxr4wVTqqhPcpXl72vMZ2Er9PN0eMXJXOnuKyrAvIB6pic2ItRTD
JSSK2sgVbHvKR6fipuDOslQFmXtqIhAwHHbDS+reo0Y+om6svDJ5BDE01ZH5ci2m
Dup14akkAmaFmrJTdQnJ1iMGGwZB/qwrPHwje7m3tu6OI9XwmdwPpU9/slOzpJVf
jHJqoANc1c08PmQPu9ckTuim6YFVivYkyRh6T/gYbfhvideOuk2HwAEYcUAr50nw
qgGiHLCM9aSO4jRZCpUkp98ghib8al1X50uH/6vgqBHDcP/PvKz3hKMRMv8V4ZTJ
sNI3tyqgpgvVMZsZ5dCusqoFhX4vpmRKU/3MZO1RvUfLgmZcvry7JQjw4iVTv/yk
J70bsHypYTM3dKpy3CEgzXqLBATGPu+joRFUS/Jpx2tn7r/KwFNHKIUTBymjU1od
8NKRUjuCOmBzMmb2KB37DDwe2tU5ipoMKqOuMR0WFyRuBCnGaWniyYdj77nOlICf
guXF51z9W55yMGmzmCvIP2JMyOlb/pE9X/7cIgjspzCwFw/GvOz96UmdvkS2RoC+
3jscTncFo/ctugrhiIqIs131zWvL6UtNqPawZMImArdQD6Rrtk2dugvr17S7NlQX
jm+ox3k0TuMxV0yynUwIawlZA50exYn11HoKtUS1ZkYlzQGZLvYChiAJrRxH7qdU
BFKZJUh2OczWAp4Eo2ejmLYEVj3aCiRFXCcG2jrLK20q7yB8URQ0EAp+dLyHbG25
vxnyf0i0Jf+4Hh4LTpkag+Qj6itXi5yEfTerBfmWEz4NGgRQh5JHJSZC1OKfeY4L
LIuL3s8AE/BUcndsSbZUIcniaqXVZzKRs/o+pS/k+2WnuDiiTgYkb7TYw0bOsM8L
qxCbX5oKgWV0mC/IoqaKXtX7mLVdpIdeHKYnPnAfUaWFMH4TlXWPbIadupa2qEad
pAv88L73HAzb/ABr4HayDz2q1RkWXGclVF9/WcBaaNrpRatQQ5lvrOlO90tbiqXA
14n0VN53fgTxOpUG3qNVi/Cgv7SxiuEP6vtoq9VuJlG+HHO9Q//sDzUH6ABIjtZ7
EhtL01Tydh7Pm2RyyQ7r36iqSC6vM8iiUQHS68Y0FcxOGFm+qhN6K4QEAPcWOJkv
/0o44ShTvl8UP6DxWQeZ8aZpd1IUoQgTY+yQRq3rIPGAiDePHkYZDsFkPCvxmKJT
aRWsIRiEOY8VAd8GDAl+QhImvdw2+ao1VGbT8Uu9KrLGgKFNvOeix9HtgIITqY2j
tRI1ShQGiUZzknTPWx9wG28KBFDD961Gh+inULBgQ9W8e8XvWnpopd2XO9hDb+QE
F1eJwrQDo3J4oMVSO5KiEo/ZPZ3O/qyPPVVmp+At4Z+8cWSsGY7X5KpcRcuRef+N
tsyJZH3pwxnPxmTJZEoJYZa6wQkH82UJTVD5Vu9la0PdXuKTgi+pUdZ66hmfZJBO
TLAF5XL8n21iQRVsRBY73x/kEpD6AVv5FdA4mZ8ZS3kg9Ts2XanA7efmMkcmtqbt
GgKgrOPLfXtOV1xUpZNly8xKH0N9P7lF7r1JaScs5ffFiHEGxE0Br+LtXZJR6a8n
s9AykuCeh8rs0sNGgFYY0XDjlG3p7sxcHY+qSQdFcKqjlGq+kPstq0VrK2sdU3jE
nbpHd61rxCaQt3tDzc+Om5u1txXcmTVm6CrPsjvnXHvumkTvYoV5n4s/BZ4SZlQQ
GpdOLux9O7QxhPYTVHLvXj6ZwlEgbycxNFF7btIRVXDlHK6mzF77oJSjiaNn0cTY
wXv+9Hn4U4IcibLA8pGNsaYoLi+2bm1alUmipnnBDepLGpfrq9QFUcnFmnZ6b4aT
AHzf0CxQ5ZCVAIyBHl6d7FQklek+4UWvsb7pi0eYSl/sDNGnLP+DvlWfPzI7hJ4J
ef7ZNXwo7g6HG/87NYi1FM7sLtgeXGO4t8TQZKUGDk9vLAl6dq+mthZSi1bjtxiA
LSEGZCB5SHE73eSjIi9q0DpseOHnGLkI6JEIlBYOqvlwV96OI8vH5to0gCGtLFWN
uEX7F5gXkhrobJBB1YIHQl9N5oUB+VtQfyqKIVp7eh/2TKec1865LgLj0YJ0S242
4qY1iKFWobIXewpHR2vaeZJQO5PG+ics/C4RvvV4TnfBFZo/kXEz4KWKb4nYc+AN
JzOTmVgPmzdRW4LoH0yTxququEIBJ0+FzUpvvOgpDM2HHWSuf14v4g3tud1uH1K1
9xzuXZvt8lNPqBhYY26ToUfWwoN5Ou+u93kA5sWQJhZQ1PaKBCA/qh2ybnbfk6Fn
nNczVLKEl9i+5Gumc0F2miQGL7J/F3KVeipXHyQQKtQ3J+8RJ1L5UAt6GFXY/8OL
BvpItWhY1DvggvgT5sUXNdAIinowGcuefjv3RNQxfvuyIUMySNPj/dT7WvJjmlNk
Xb9CNuEwBkKGK2N1fRLIPCoCFoTmDQwWb2vpugVsxPDO4d8CC07gewfZVCTUQXaq
jrK3cwpIxiPwfUwGAe129lv4kw+Z+QdvXmEB8nBU7BFhuO1zwYwiHs8HigTjnURr
GP6cEYReSvb7b+2dRk9XStWMUIvPYzwf58LRZGsZ7jaqm53sRSq/MjI7PILE6O7D
wV6gmvZoD2jBXikZr8Tmji3ZxOSwFa4vqN5ZynkzzR4lpjbcEdrao9Si4LF8OY5K
A4s1aLsA1IN1IR4IEozz7rvRkm8MQRr+MpSmV9/6S4s+9hTwBnO8emivSxeBzf2v
0847A9KHtPtgb+KAx/Ofig3AxObGk1+WSjGZctCjX21OXOLIIJhphCFrbKXD3RhT
YQKuZ6yoai0Bm4RNKfudgGhPUT7cTksdCv8jxMeNeFEqsOCXZQV7J+B4pMcZhY3X
qYXnzMwtdudkwkuRphFQw0j79yomgJBIj4A1EXVfaWaTl8S73Lri3WXQU1ZRU/zn
MsUOHI2lDgbM5NIgKZwjkSxlvav24yqZ0pq4Qz00CQMxrY3zGJGn81KKyakkI+Hm
f85kE7IxxRVB6lx14it3vu3uhAQgGU4Wd5K9pLF4pHMjBti7jphjaTooAUAYAuxq
uxB/SyATssjysfkMOR1QiK++OixaMxf8jPF9HAJatRje5i1X0WKjOIjwgSNd0rd2
HPwyYTa3/bvsIqowwYbD3DqVmW2nElOpKVXvmswab3y0F8xDpANGq5+slNCDnngW
bIKwrOPs3XwvV115JK+qv82vTgWe1259bBt78zDNdV3iKi1auoDA5paHpmE4Tibx
yzywo81PfMFcNjN2D0XrT8K+Rac74q4onXOHh7tJneKuNY7+pqJI12zD+xb3871b
hbHNJKuowiP+DbGgqeoa89Y2G5U6Y1Kq4U/u8QBPTE+Mx6Za7DbCoLg9BFB3srgI
kglvz8M7G6AK79A1I3yqnbQ3xKFRqmmNvnoz027uVY5BXUPJapGBwca0kVsh1QLc
JAj6tWxIPST7Lael5QQrEEK8P+2mY5haBtqdXaAQMI81BLgoELg0asccWMUeNBNl
4OsHmnmzrHm/Yz8niaAsLqoK+HsBx8s9hrkvghBeBHVQ+1JncoB42P34ZsXpYCVj
9nUo6eDm6oscy7AaU+NTd+cqaxn4KWaI7YXy4slKHgEioCR7KGWwPe6gqjNkZcj8
/cqrEs3NYAqwced+hKAnN9Rlrpzdj06+dt3c5X2P/K6COmJ9eBDXY8YtR5H/EH6Z
abpKg4NosV77o+ZbJ0Yv9vRAvb+oQzSHf/sILnfAbT5rcvnNdyyK8+JNHn5GJIU3
ohxQ/brnKDh6wGVPhJFvNno7uNosmeHsbrjWPMrjXfQQD5S7hni4Z48/6kjU3YLI
EzlYnmUuGmUWFhbtxznhtISovxy+nGWYw2DO1+QZW2eUfgH2P0hiR9Q/65DM4YYx
GC9R4+7FNeaUQCVUHNVop3yx99b0w5Zf+uRukt8uyYiryGuf9srtuj/W7/ohJ8tr
/5lD7W3CQuriuZXEdmiW+wg+VQn3hp8b9bneqxmQn/5QCBWMj9HPYxiReR8Cp8Jx
3cGosmHHH2YjjG6ttZTTjWZkKDCXQnNKtTrcZDYcR1YtBUs8qoUhvZY7NTPBaZ7y
nbCD1kYdbyIBmYvum946ENlGMAMSCEZjcRh0us/y93F1cg9p8pmvUQP1C1QZHvkG
MMVA2nzmONSrf7e0UMpPgEF4tL295c6s3a9ndANWyjcJbHIzqXvp+qhch49xSVRs
Mcy8s3X64Rpm6oJtlDphGXRz882N08fs3QBddsxREPXS9c5gkqivt5GNYlijHQu8
fhzpUST6mzOauyWF3oNvprAupBhSKdpbHFmnQG67BfYyzrDLMl5L+Wl1PJKwxVZU
yIcgnk+q2TGwBOQuQbKsE1kAmIOozvalsoLWMoivFFwdF+rp2vrijRoxKmriwnPN
ww8m15JB9EEtU7L51xVcfERDGxUBmkrDqI3YI2zlXbLNO+uAKbjPBOwlLulCBCm6
Fvu9nWIXB/CIYtRX95nqbiEq+djHhcC7Gn1x8XyNK25or/VJA09H4TahDHV5YPvK
i9vW8eqsMVGtR3DnRU4Ue2Lp7oTDZTqMZEFIevzmLnglrBiUeCSn3AccwG3JXfjp
ljgSCRYc4QT7FiqhzD4wFLpEUJpbzCyJgKeX6AiWWGfJ21RvqZJaPgOfcG8J7Ok5
A79lcoj54uGJyUj5en8pdX0vGPfcclNOs4gdVkAQa83Vr8LpVcx9Mi68q4Q0Gv/n
Wmv0EQjKXys1KJjcLPEdSFgq4F4Dyn8/M/Q67bW26FE2XFoNKK/bHJPaqrqONPnW
UMKMU7+9pyQwAio8qbKUWmSkPkueBFkC51Rvu+YCScaMlNIiLUOTMZRXNa8a5k3y
g28yxYwY3Vivp1Nh7yZDZt0D5gsuGPu0ECxBwolsP0ue6xRd9gh2Q5/ugKJo94Ap
+CAV313BB4T6YkZ0bFDGlSzoKKRuyjt/409nOVk3Q/LKqQU0WRjWoUQLUDbPFYv4
FROIs+nyxuzII+3dJI7nrqr0/R55iizCugysnx7HreDa+ynkQOVek8b6BcUltyoJ
ch6/EeQfYJodwdC4xx5O8OCZ8zgxpzIaIl7Xsu4JvSC6TGjcyO2jHKdSkP5Dq8ap
pPEYj0roGEjKGxGkMFvtY/Kt7X41pksYAYeEadOWYA9g7Ui58u+xldazXvT1Sc9/
LSOFpD+Hej4WNibS7ZJj6qYv21pRgTJlwQydj5RULhoHN+fPDpi14CuouPKE2HjN
wy/FItxtQ8eN9s+IvrxtqClh3RGwQQaVw0k/EtwtVXxHLD573vrxHsb34qltCUbU
RocCwZfpQoyVpGh+CigkR4HRzyGXXwOGoL7oG+zZc3hgcUhNEsHXtijA8UILye2V
t6HpRh/dMS32ES0iH5DWJ/blnxqqj5clYQg+K3xrTcZOH+jgwhCBLtcM8I6DivGk
U6rZKFqwglsF3++22JnR8HR0ww6N1kpUQj7uG/+zgCkcbCHvI764ga1TTUpF7y7o
7SQrtmphOHn4Fo1xOSv9fPbSioVf0cay7x8Gl4YC99Zs1mi0DuU8uakQy3Q+nzKM
xZJ0BmBTWC9rcDLEz40SWBN4pGQW7PVTD8AIrrERCSMfgOZ/gRhZa/6PdYD9in+f
OTusfLrxbVbvyt/QOJp7QqOylnZ73RBGZn17DZ3j34RzTaKvK3F521vGz2s+uhnR
CCVve2qB2BB2U/B9X9f2QMyX1sW2jY+sLP3bi7rPCHsOlRS5cbBMituiY+IhwSc7
uZbgO2RZomk1+Spdimb+nZ6I1A8iAPC2UR7pUVBmjxdEtoqqcqfrXGZUHGkY+E0Q
92rp+lrqaQu51tDiTWTjxKVYY3WcBdpFrhh6CLlfDoDHJxBxVs+EvCWBw3l8sLXu
Biu8iFz3dodo0qYqlOgYT7P87tHSOzwO4vCynVOeCWmKMXH2RZHDc7gTwHX4MtiQ
bknHN5xAHUXJmZ2EpmDInT0SilKcijm9BJIzncGULOBBKuTqQ7Bz+1q1WvktBqIq
ALiUgKdr/sKML2E+jVoQxX5q0F9axMAXIL2kl81jzQ5PSr6uXlQDB4R9r0YKpA0r
EEXTPGDREetZmCupukron9v2nzmq+JqDKp5M4GKS9za3hCTJe6LGWkrQwImWZMld
eO5K1qnHYm2iyGkWnnBKQfAdqRoevKZ1yJg+6l1xV9z7ogCAMign+p0ns07fN6zT
whdwRNxPW/Jof/HcvhLLENT9Njg153RjRMSiBQaTlbKcUziq4Nn4WNGxBJn/mdQo
cb7r0ZTrezsj2IzNbyPVQsDea8JAkHOCce0b7VCwk/ce3hWDCJVglWdoIODAosyB
gnx9Unz5qP+Pn3CqbMQ9cDSwsZ9n9wZvPOoaUx3z0XenYvoZy3bKFeIj7d/zFXeo
BH+qDbEB8ELzVV590MRfaou6+Z7qz6hjtEP2ecdJaAL0uFfXxu2+Frizp59/qTXb
2E3zEiBpxsMqfhzgUO2QftFVuKqJ9SWByiMQSftdkF+D+EP2v9vlIAXUyp852QYl
ysOMXjoXrZw+Sa3c2Fntycz8qN+FZ1ZkbIvY3ZYokGBXnwDe1ubQSi0PfbD1iDMJ
va3azeF6Y+IX8q+iQ/X5n1kwzC8/V1clwQqMWxd9IJA6LydyoSYSI/Td4Wb6uR/Y
K1M/pj9F7L27U75eYnTHzD1tN8k4xs+6YUVi+VI7JMUOP8ax0Vm6NzouiEg1bKDx
C3FMjzuqoeHN0xq4MkqgtOO5tyXespdflmj3C982KTMsyzOF3+6EFCUV3rRchsUO
Ekbzq2lEKxD/8BSZA1iG9pdKCZ6QK6qnyK3i/IpChyj3MgttrvCqC1RsIuRG+Pdl
eWDx2OB55aapv/dUQNNM9cPl3cAZI6xF+UiMWtQyOdrVboES2U0QpXcHQaOjkuGH
5DRMsCiDpvLdWwizFxlNtN5Y1lxzpnmqab7gvX3CfJrfBmYkMeKzXvYtswvpmcCq
X+JC3Qo4/4BLvXlIbLG7u1sYgBOJ4FgzheaYSzG9HmX/a/LccF+527ZfYqtkOy92
j2y5ZwK8M4nmOIkfbhcoJETNVUn2tuDOIPUsEfIEYiR45+D8jzJNJNy1ExTwG/cP
+1xON0xwzw9/8X6UufJcJizj2y4/Pycnb3vQRuku1zRF980QU2844CeLKio4Dfc8
4/vzZ+kvUPuXTpRouPVMnS26M5u+KRq1X8Hz3YfU/ikPetLbm1d3gWfPQ6Gz2wma
rOfWb3L+IVD4KL8sWW+DXM6gscPAspORs4GZRFctaAcC/9D95yS6DhUrRQvN6sqB
DKLVgqPAgrgSv2SYQUCn50WnIZ7rXo5yarqlPXjvonkYKphH2pLHxwzIRPRb2YdA
tS8RUsqD6zJVhcC6krVygPG1qhjH/CN4GLedWmYlGkstqyCEk6Xi4z9dvK/R0qdu
P+wnht51+HeNlBFAjatN+LdyfuVKPs3i4hrIeR1UfOF0dAQ7FU8UPjzyx4Oy8abS
/7JV4Hz9761GBLZ4vgJqSABktIFvtThjvD9UdhuRswVtXzpv6rl9plov6ePxKX3e
kcZDaZzJANzCZvISrgzWlsTIbVxdTi7bgzGnEAaR1JulUc/NMN6SANkRY86pGCuC
b8zww6InYIpE4pcWAfiHF8k1NESQDmYvm6uAdgolwNP1WPLy8FVxTOkl1lVD1BaP
q8+SwtnB0rBpqeDgjCn7GWDdiHgcUk/iTESbcefuVjusz9+ccUIUCMcnKgi4HFd1
PrgYqr81Zoma/7cd9qTZKfmyspK0oPbYT9MG/ZTUQ7x5LvHifQUqYV905rkC5xHg
HJGDo3RB9VlQOAKVIAk4Mh4uu+S4Tv3iSC/EGdDTJBofxdpJ+noq8iR9nTn3iNzd
JJT8dKOVLZZ1U2kBYKB0yhnw7fgOcQ8I2TAftIrBepuw1cduy0iihFtJabLwRe32
uDKLyKKnYO0nRo5RH7LAYOlyrigSfvC/zbmUB43zcS6noYJ8Zlr2wpAdqsSu9PLJ
P5vH2DudRiWvMh1I3H8mznOhQ8T6wXw9otWOBUsK0w4OWBpAC6OW4bus+pzmDt7A
KX5FEhO6S8xiFbQmnUZptXlr/FvweaXlZuNUhDymA41aps/I6hVz01Sg+xA6srYD
TYHQ4NxU7R/8nhENWGNtHHXKPwSasfu/CgG3pJP9vL0j5oenekRTr2ClZui8Ni/n
TAlZX1E0HdWLfuG+GL0PD0EXSibHDEWv64Mfjh1NtZyEAj1IaeflHcqm4p6G6q8k
+G1YfKmp88I4GgMFgfkfdhNvOR7QAhP3OPW5I4XK0m/X+o5bLsM9LEjZwteTG6O0
yvB5GGb9a6eETwC+cX4Z0I4upnS2meGIvPzyd6xvtweJKjAFLrAjhAm1f1KtYh4e
jPuA6M4F+1UQIlXnB/m3ACSm/q8mHixUfyzuJbaXUoFOhI3S0n2cK1l1n+aZI5zg
ztBRb4gDlDXDpAfX6I2xKV1TTArCJ1LX5fBNtJpEKz67+PHmbWgW5je05+GMvqpB
YWQYH+dRHrp3AP/goh6SQ+ywI+JuMtxgfGpJ4wdn9RZZMKunt/I2Pyx1F4Oi61fp
z9XmfNgn3lREya2UA+x2hzdiHJrTS1KEslOulbi03BMaH4EU20PUBF9m/GhDKbry
rG22gdukGvCGqib/5s74U5fsScOGZFKAwLRBjjjP4UMEfKLHniMxZ69tIkSRbEGY
dz3wg3HGHiuR/H4Pq4j2R03TlD5cy/05SSGN1NPQqB9J8H4lrnU4iy0tYSjFYPzM
WKrWX5FDEefzvGSSlM7EOfitSuDkR/GqQ0zqFwc+FPZFb/6JjpjGdBFd0iXVc5gr
OM6+rgqvbE5YM7vgyBhIh+w67JJHr/9u/gGmSl2PB9ki22fs7cBOTJhnTQOsQoyH
TyTlj+1ZTu/OTj9jBBSYd96Zag8lnHskAZD3s1BgtHM5dgNshB8LOhFTi+WBWNG3
yLA7a8b2iN55Dd2dJNcpL8Mio6OW5SX903jdXvb4PQj0aHFjaZYDC41FRPbJC8WF
bQWYSBk9UfEPXCPT3Kuno3+Ze31PeHNko8HcrltndK9FfKHHmheaAWvAA38HGqw6
c2LQcdPbsajO/Qe0C7iEjcyqa5HktiQjhsZRG1E/mp21izOTDhEfMWRSu0u7d8Zv
Hw8XK4l1ItVf/mkIwJ7niCDPaWucFtMRFu1AN2gpAOn6cil8KYrOBl99GwXaCIrT
JXhxqVRckYwLgvf6mYvoAdue1GAePXOJeuWxSuPrGlOqAxoa/wfe51OK6VKKmm/G
iv38K6oNogb3Md/O3DGCkkAGpFaX7MQRlKmI/y/gzNy9/PXGvsz+Wk68/QdrICp4
XibFCbTAIS9B+NQlobseZC1iO98iRMnG8P16IcCqlkZve10Zma9NCB7n4m2OGCA+
iur5Iw515kxJYuidC7sUU6pNMYsBOw0EnBF7OCA0kBc8XgO4HOU/oScL+r67MnJn
R3KehGaaFUSccXGCPpIxzu5nvirj2BZFbzd2NajxudTLAVQMQCZbenq5VESa5vfr
4V8I2V8DqKA08AkxRFz+WZNggXecSKWSML7h8rxaLlWhIz3Zm1hE9UQPgTBEFT7M
Mjlf28I/zG3ka17ofSDgfPq+bBralRaJLlX0i4xuy/uBidxYCVrOEcB/KFqe/4wO
OOfKm6NZc+Ge0Z/VD//8o4WZyX5RH7izpbyVf+/HRE0KZfAW5Mzy6/0k69POUgv/
U1s4EHRe2DB7gHqVKSKonOVFseR7S5OVJKcE1cggRycEqvwi5KLw5wTQgGvQv0wB
WYS0UBAT6t7QETIW1wWv0JrmQ7qeH4ETcN/6XF27yvl1I9PiySPvl0Q/PX7vDyVf
+4SkqFLmFVFdi6zZSgTg1BAkDF17Cpm7ujrMt+Zh+NldZ9ubjGTP45KXOay0EySf
kU4KNFoR9yQLNBawYsl1JefQbsVTld/yqKO//urHhJ2wklRORdqJfWSj0yGs+x5p
hnybQONSd2uW0CncBXDVvnL4vBesjXRuihvyEYYhbF6rFQukHSUuHnQ/BA6RtCiR
M56cnknrc+wsqWpr+p8aLwfzY4sp6PHMTgS38sL6EjnW6ljpuO/gxsHzXCRosmO8
ppCBZkEhZKzJ6wwA7ay9QdRqJh2+g5iZ+4JCm/cYliO2xIfmEDLFOZunveLaoLoD
FmJ1VJfEaZTRtDjbhAizl3K4ygM5HpYYSBe1JyqVNQkua2IppyMVGUg9H+f766FI
Yzt/N/N2HkVOpUJAXby4HWNVsdd9jUCAnKnrW92rw9UDYLX1/wbuZ5k557CqDg19
JTTkvTZhGGMakNCXOf9b1yZaEkz0R6KxvNuVnIaEDUmDXmBpFFtLqgnZli44W0Mv
MftbkjpoBJMJJlpVReNuFhBfMSkDX/oiKiBdobo7HJqYpk8bSm0OQRwPD4z7gMue
vVyklsHkT2mMVtxuAYsrOxrNf+Xkj+q4BxmOuJ3Zjj32uPOniB67uZcMPnbQS2+y
5tzDhSz0mqwOrIdYu6LWiQdyvEfuCm8JmS1xQolrCg/iaRzfWT+iaJqrXqpF5BJp
p9chbQWmW24uAjE2VcPtXtbtcmqR8+XK2kZwz6irIHIVycsXC5R5od2YRkjklV4O
Wt5mdLXhq8p4hFS8zpXFSR7qWEVEN/VXJzmpdC/OP9C1khU9mj5Nc7lvUUircCTl
ecxNteAPUJP/WHLZDUtqHV7zwTIuHoKZkVYq/M0SgPbYAtnNoXx5SzAfAzNx1BUU
FAhiaCEb2ngdVwOjn8LX/aomVtOFLxaV+KDCpGUWmTnFWid7ClTa1FVpu5auf4G8
FEjwpe1++jRpQUcOyIyRHY6b048Z9wEkrb2cUVXglbqku8lhSZC0uCvBFZ2Kn5D8
wmK8RG5t7OpKEaz59xF6MS8kR2ruT5/HomLUvNsB28qAo/2Z9XVDtf88ZMtHp3/E
tUZX685EC3oldm7PX9tVV+5gk5mVWb+KFWr071lGTJQa1N5m8DgmLhGBxrJzjPMs
0i9QV6gOWauEuA8lkFsTcJb5xNX0zHaDit+zhzQg5ucdFgu0+MNe1Pplo2mR3VjY
hziBf4VnPEyvCOWNNGp8jqyJQy0H8jzpy9PWvkoWlFkV2P6NkR+J8bD0IKPC+V/C
y9/zMydI1MoZQ0RjYQjs2raWuXTFZIwtz5Ppj7KU/3kOeGq4dmHEq/E7IM2HfRZk
VAdA46KQOSVB6yGGHtDx/ZCptPHmSB2PeWU8Nx3fDYI/m4J00cL+IRp4/ClkR75N
nfdnH6YUBPYp8Kwy0L/CnvK44eSMehDfz1P2DLzi5XIaMsFAXLRJ1zO57wQJh7Og
5vrE0Tbx/RWpd1YXJ9JHFevUfVpyguNW2r/96PkrjuVmH/+QMWk4PLlpbNpidNDJ
Jc6VUOZ2R6QW5wLCpqSMrMoxEuDmWvYXgc7pBq36AwB1x6iUFZM2cHm2dpn7hzHA
oFUeLCle2s33M5RMgIbpjcMcfVdE0PXy4By7TDRN2cxqoqnfH9Au70xS7J9xlEWi
x2IJwazbaLaXr31lg9kbwUxldTV27Z7pCpSYgW5Z7iMyI9zEynczzS9ZpPr30Huq
QFShYj2I6x9alC54qkWl9e0c8ZC1QScbQ+BwhRQiis6WjvhsNwS9DemkjS4JQfqN
hhR/syxwpdXIdPupvURJ0DrZ7MSOMlYCetpVMMxpj3AEb7okwL9mFLnQlVHEik/a
OLRcj3c2Ne8z4ZwI+UWeKo95Asw4KoaJGK+T8+M+jKdNJ9dEwJGsloV/QNi6Tt6d
SxAMTzD94QY+INNK7alxy2lBV2ZZcCcT0vsu3Fh3KX8qk5FmZpvglvUhorZJg/vD
Es6i0RPxbpFaQkkQwUzqjVst2sPZkzR0cgjoxssEnSpizLHH9rR5Nc80MnxZl/9W
xGrt1W0vdtC6TnrmY60E+MtZd4nrls3W45w3rOBr48GmxnLYGwOzsBsJgWcpSluM
udUd7Ws0ibDvM00o5UZpH+XNBbkip1J9V2RDr/7VBN8eFS+CgtRqY2J1+A28X2U7
RFUl0UOCG9zR4mmKa14ykwi1QzB/VtGiiviDn2ScnkHCnvA9LadeuA+KPltvEi0N
ETyWg9E2vsjNYKgXS6ITFoe1/YViCcHZGXfJnIl8bJA5cFkiROTGRzHMU7p+FDr/
k+Or6IiF0hv7XUigmC8einbdKYEsiz9kNZVMFTJMhCo92pZeOGDNwfRtybrp4Qbe
mRgw88Ss+ijZPBp8blGt9moHwS7KcKBxHm8w6XuJiFnnp4ylhA9NmMjJr0NlhRDg
J2VGsiLUdlcYhRBverW236qgNQNZL5XsikuvcTE5iN1vDfylrazi25goWI4DocB7
NiWzfCjaXoJPkn/ALW21Sc9kNq1WRINJvVjTaLM11o+s8uJ5h61ehje8hFG1kUK9
xCkDcfcOSuCrqGzYfCwE9yFUjr2G7KuNpkVRXYp5mx/QvrfBPaSqL1dzF9C/6lYQ
u/l8BOWR/7B7w+g6eenCgaYW4xSzjiDjot4QfbbkbbllFai1Dpm36RW8rY72J8qr
+M0bTdB6FV5xwM/iK8lCWfxyRv+sD52RuvUulP9UBGgehMYP0NS7wdI9I5rocGml
e1xhcxI09J48gScGoUXFKijKMH6AbhUrUnq6p2z45P9v0sT6E66SnXoVAKtLTg5p
aRS/ef89+RX0JZZpsQW98nB2j7MI7oDCfej56cK9lRsk9YTPC4kiXVMz+0GOQytQ
2QEXR7WEb1Bk4e+nEF4Xy3rG5pXud0ggIq5GM9otZrNmR3BtCp+Q6qRrpcNYKxKE
BXB6QqozbLntNAR4Wyk8kw1L7q3UPXFUK2dae9uX1pU+hA87DBSKES33VDr5RdGv
hyIrMa3qRQ+ZL15fxrrT224/KyPidXsuQhQgVDNWctB0xFgtKrmGyMvPncbgo2Du
T+1/ePY277GNGT7W5URw9fcZxNUytvBbGGrJeQkXfSC5fI4AxpmuJAzX+HKauVFZ
VqET0Lrl3oTrJbRvpMlWRXkyN+Y7p3hmpuUzZnYNQsZeOnbKzlDPQtwRCf/GUlz0
VGp3Rml4g3yC3TCyNxA7GO31beImt/txnplxpeMesCqSke0bt5gy7Y3RwS3vo7T5
25yoHit7TwtPuUKbbW59zZv9eVi39xGs+rRfOqnkM4/2tSOtC03+WNjRgNx+GY5Y
GPlWJ3QpcAX+YFePqwTFHUKBAq8dAZYjXLsk1iY5L9cPYHbrCiKfHUvrz4k6pc0S
DEU+nIRWxLOE8WO8jgjQgzYK/HUHt91gzdwDPIK4stPjLJauqTP3Q6zESxOpNCdu
MG6zD500vhA4wg3pskKfk243TSO8uOUL76hhL9KikrECL7TT9iNo6Juagd9MAFnV
vl5MF+u4TxanPpcaL/dB1VUKUMDyFr7IELBT3q4RoIKnSqZ6IaNMXNUvDJyCoY+T
jjE1TDioHLdHiIxuUwYcN/Dke4HCWyfer9D28peHUuWAv287bFFMx2YHvudlmtKw
uCMrskQrIYtCyGiqFRK2RYbU6UPaQdzJ5Ex3jMyQOX1VExJarV112xJElVnWq/8s
vG8O29zkb7MsfrMdmOHh6TbcqWoDF4wX89gTlmsFMROCWupRdyMF5aDcsREyQaJn
dpXNK3tDmYYPGfNRPEBeT3b03euYsXb7ydilctr8xU4fhOS9LeWpPRH3Ha+/ZID3
NKuQVckuqqCYNP+V1XuLr4kKysC00Bq3YXpPP9NcjQMnLUC6gqi+Xr1XLpNNvNyI
FQIogzhIUaC9HE3nnxLdz5C3R299pxrDsWVV+3nU0KCzK5G9v2XIxEa1klo2yov6
UBMwfC7FSrxY0oLM8ZxqSSOjxpQ+T/Zwtnpdf3kM2RbfsK+Fg29n85xLK7R9Zqv9
C3blwgZ2Gt6Lz48JCRrV1RrIL9qg0CkTaXxHiXDr2r7a8j4zbphABMITwZn6NWCQ
9S3qcZXkcoKA3vuB2Oz+NqSuvMbupldiBQm6U/lAU3Fb7C9Inf9M6x+lU7xnpAF2
ToKp69S2qbZnIxc5Nkx2twuMJBhac5U0Jd8/SAHV9MHtzIUjLQk9a+d9irpB5esU
uCYI1amM5D8w+588QWG038C22+lVpDmXScwDyoccFKeIZ38h0SYcyEFKEEQm/Th6
4auOkasPOp3yKYB9WoTuT3cq/SCzlksDaMOW0R1xApUwyE4p/ykTWWq6CgzGDqbh
rdJBJcSO92+PIgaBkDlPE4thi+zr3g9cnKR5qgwId4Y2o4eZwWYqS/woVtpFNTWX
VAgw81JjCVC7clFCxwHqZVmarwZ35X1bckCVNAM/hxOj2iqCeUqEcOia1vdGKJzz
M2WrtjUVpfBdXwIJXfZP2cEsGwAmgFx15Mj6A81D/aWVmIe0JJEhJIfmw2kibaki
755iGhhkCffl4jLCRDkb7/tl0LikRTIjTwthLJLSlF9WJVte00lGtDuvW/2Ge5ph
8kOgGaZfwi3ItEBv7Pib7/FyLDjrRCp/g673lNZ0RU0VuRZGYB3DgE4NpeU681I6
SuEBj5a1h6vWjJ94gcPJLoQekB0uo0+hlDOIPKvdnI7b3iws0WbGR5ZG9hgCP64o
zrDnmGn5E97J+XYxPVKLN4QFfjGQzaMwdyi16srm75ohzr6PbCNHU/vVBEJH2Cb8
mb4nLlZyPciytq8IL2P8T4kBuITet++jhN6qwrLFAGkMFaPiUPv7sKDlibwVG/pZ
NAG1nfAT3/aItxSLfxKb+1KLvLPGANt733nBMYz2l6Nh7aGsARObOm+73MH1xkZ4
Xu5CTLOX+bAbGBMhkZ96fnnCMz+lLoaJl8duU25MTtPToAppj/VzIKVMDdFAj/OO
r4ln6HtsHP+IP7FUb8wnsirqDMEuTACKtrc6jZAQSxRWv1VAZ6u3l0xTP1uCgILV
kyGBJsAuEHcGf0Aa/tQa970ENAOeZwxoX6hAEUdLF0cD9yZQZJ0MI2uiZdP4WYuO
bjL8Bq672GFW0qUPHNFRB7KZ/IvOo8d0bWyJ+LrKC+LEq/NjrMGYhVGv5L+q7LA8
Y2Qn9QU85dT15e9jvlZ3NW+p8voGsRqxmK0XtPw3HYdMT5/jADEgi+AEOQWz9jn7
iXpzPT2DVVjBvZl4AIQt0J1xDJ/gPv7hslLY4gQ7LMBzf/BLI50CZd81Ud9Ep3oW
4q7Z9eTQD3jWTJP43GaZS0IajFgm15MxWeKRdf23ElfmZEJWj4FgCkTB9y7y41cz
kXpQ+OcFK5hH9my1fzitaBeXyFSdpJzsVbZHVCYanEDQGP+Uka1b2Uu3HOqZA24l
WnCcMKCUU1sECXXIwDGbop+Lz+rKT9H5iUklsCgllpWtqDCrpgRukkpY21LfalFW
3JxU+D+2/MrAf04Z1XxkyAVCDRDOhJwiotpA2w6tbLb1NpoPrHJcP43JcUehIkhs
roxdo9ALlsNGtB8MyitqQWjbNsZ2tPOIRwZcQTQe8YpZKWM9Eg6avfP2pF2DluyX
Ax1ZQOMgsGXBMBt9sUcynP1SsdnvUpHn9aSV9RwLWWETshlBX7DKtLc1mqsL1xcc
1OMlCNbG+Ruy6yRv6pcaVqggVXpQVkZG1cTYeLwv9fuZU6PggDzU1RDGrMWvX7Tw
1wMBgNH0sg+MOdLeDT8bMuKimxc3bWF6lXhjFZkT8zR8HIJ5eIK798x9mQHkab6j
YcMScVVYyigBY0TwiCM1TYnkG2R5b5N1Do8dPgSoEL/cpj0zpv/CPYGxS6r3VQAj
5xjLwGEbv065J/vvZ1XC/xG42GrdiaekecL2xgDWlVrHU5rNoUAPH89Q/vWWOtwm
QsEunlerJICryRpfa6VQMkzLaZgohnZbK+D0WprGeEAu6qsPkDELIbfXw2NpCRzR
TnLqGyF8/Dc8UHnowETIwRQKdHvnuG0ELsR8a89OinH1JBf95uzVX1Pin8lOLYpJ
olQDKZlzTrY9usqOmBr807UTHkCActZncv4apRxSF26Fk77MKw9QfiXi1lquZQZV
KcjZkmBveF0uoE1MrCNKwCHo+886sLEyVVXvqVCq1uNIBDG58+nLHUhg1opX7ysu
UXgI8vlYDqJEbGGrVJAiJ+h3yoKEao5ux3FG7XG79phuMxehm4L0uS97u+FPK5O4
TGsv06IjU6aqSXQ1pqUWMI0RsyL1/MAYxQZpdE1Eea9fuPWhyCoR0af/BnUGe6BP
OdoTcPK6w/hKrYTOxDMFGHqy1C3jI27piTwcv0VOyix2309p3wDzSymhBb2guGLN
CFTUa0n90zTLZHSXRY8X/U/4NuzVONSe19Q57DIUZDY0qZvcJ3tq+Ze3ByIsspuB
qiti8nl8a5iz6gHRQ+3OpNDgFPXc6j5ZbVl0p0DhOQTHDEGoK6MUiTD2CyicqQZU
SYtQh21t6hCKmZyWQ6BgMyude+MBI83XP+yPD564o1XEWcsIM/PhOJCAJpEEnjLZ
yJtrgF7Uv8uidGSj+iqE3m1PrRuhEj+7GJi0EBISELJnjhPk03dpjQzFP3gON0W3
l2mW1Pt3DfqXyEgTXum9cesmJihITn/BGl+s8LRhsqBEtj8q3A/zTGvogCdHQ6bu
CyWb0VrsGsYYYgDsxzbh7KzfQuPy7UZijHIEDRhhSZKvbxe6iMIRUvp5+RfAzimh
cvI2RUXaNfx7E1Vva0gR6RUxZgsIM1OCIabPc+7ald4I6dPYXw/g7yy8kPa4G6gR
Ytw44nJ/vDfe7KA1S0I5lxA1dCYoJivaM5U2wMD7WqBinLY1mG7RC1gczHz/ZyV2
6iHeOh6/3t7zkzmf7aGq2HhXRe0v+6mFMZUH3NP4sqCvp3Ev9NnrdvRgrjAkEwnz
BNXJpa4jWjqKYEhRaxjNhLzJv0ABvCEz0yKtry9zBYpxv+ONAQfnieppc5vFTReO
mF/uediR3uYVUwUjlqqHsSazPY9N3zTWvW2xivFECDsu+UpM0FdxDhDT/oIHUt7l
1lkFBSNTPVDLzw+PjGMfSVTWDeZUK0x65NXx2WHPuIyrclwf7k6pCURzG8Mc8D+x
9bbE5urstp1WwAuelB996Te/lpxnvWpT7+HMoVrHlHxGloKF5iBm7VXiKV51fufV
cF/nWPu/hy2ElgBqk6E2+tYUSNcRz/XMbePMCGq/9dkz6l/kBvwIyCabrmJLtS9k
KVNirSOAdNufsbnBpL9R8Rltjg9IlzEK2D/JAZ9I3c3rPIgh1f9iQ8mB0QUv2p7I
HAzLyRVEdxo6nDRJU+YLCqLUpPX5RAlq1LuRer6i7GuBnEAfYKmQjo4ukw9530Ob
O21Tntu99M5tJPGyOcNZHOoovtUjBz7eFWGy115u20exMAxCkJXqRfy6MRr0dTQQ
HsUtk/y6wA7kZolW8dAIKm2ZUWUWWlO1U2mkZr0V0YMQe91Z8I2q/katMGuYYV1a
P27oQvYgnO7wM2CNZbugrRFUW4Nmo35uNlMS8K9nVESGSpUreNzTKWBQRYfMmSvs
ah/EGQsR1ox9Pyar0QnKf13aUQhUdzNzr53SZ2qOJ+fU44jaliUk5MCNGOWdPVjO
fHibkw6/wwGRkoYUwIJJgOsTywCD1QD97nqjrUwzehrwf9FbIZwYTSVdidRT2Qrz
PbjOq/777RvT6sM6x0v9xQR4bVTZ0If6rDTqiavoLT6IQ0y1iKNsLKxp1pTZPp0m
9E2qKsV9cFOkReRpqWVwv+1rvZI+LlNj98gNyaGO1AMufbMdsxy1p+cw1LHDaVH9
8UBJGfcwZQVmOcOniBCK9vlk/SY/6bI15T9FPNzGojOHV85eTNN0ndzWFsuAEToR
3pQd7LnzDvqz+2rIcxNblQWDpSpuWwX3x+4mSCsMOumZz0q543fizAjO/KKaB0jO
ZY5EEYg3ZtjEpb6IwEwdJ9q0vF7YfLQw+peQorspRJbr0NFloRBwnrzoxYIaOnt7
JUnl6ee7iapU+odfEpu9y44mlCttOk/HjrktHT+1U6+tXUWHAbIoMIznYIqqOqlV
3EYSplzxcTevtTL3yUXn8OP2OQ4GpRsmA11nQ5ajRNCVpfMGWrY6dQyGXsddTYzS
ErqOSyXVPN4nPEmrV8joREdA+6VMzhUAuI+jY+LQIajAA1cV2Fu3eWJx16khj8+D
W3QemXwozrFG8TlSLfqlFq6gx1qTHj3KabUsrJairpiTYB3qXPOzRpa30mLEGZR9
X3uRhuTLhjawHQhA2iwTKdT2LGTlJzXGVZueSXhtM0bCTWQQvQjLUP6MsMg13xhE
jsRLic7uOj3YuKPCc967IyUUBAvTp7K9IQ0tjAFpbMPzeX44hr+I8GAkqxTfL4jy
SLCDI4Nom0PJCg0aRResy75Fu+dZy9m0Vn6kWd2xAoafoEU3EVoaJFhGJmffFrBa
u7PMeb9/sOTi5Ao4JBS38eW5zWgfpbURBfXBu43CJ/D+QgwGw2D0OSTYLHAQZHyI
MqhicZrjzIKoAOhuk6cC5BR5iGEDsCR3VrahRKZxYqyur8Zud0zUjEcy15HWJ8n3
avpjxJRT5xG/PvZe5EAoM0Aw15YkyPxbZP7eO7cZp+VX2UadGlXSU4r74KdGyh/+
33nDhRL7qNTX6hzORXl1ByfQDelZJOEHpMRERN54nEmYZJfDtGEBB/OUrnfSoqHE
GYHufGMFlsv+J/l+WhzEXWaGTtviVF/Ns9bwBm07fTxnThtj7kPG3TKnaouJzgxW
sJNnykDWH7L5wBRkhNND1zwX7q8nfIByDiv9ZKjqdzuPda/MaGoZOLh/jKrffHAC
FtdPY2i1gpyRgt8LkjcrV8KSX2fMGdAsq68jR9I4hHMKy7xzj5xbeLF+OQAV/Rsf
/Utz1OGtKn8lrt4spbFdBlNsmYXPRdixUuDECDfDWYGIdTH2s+GVN0L+j+or8BJR
HsY4Slncb7aE6+yEbQLk9AuSVDjgf6G7L8pmwOqafCCM54ttBM3OjAqPbhhKHOXO
XQ2qPA32xSnqKcs65WN4gQAtvMEGYApPE02QvwcDFh/9zvXSk3Zl1/kJswXpATJX
aAVBCoDdvVqm9+pnGWn7He359qHvUNsN/llf0qSQfKHantiaJRFN6yGnQuFrBDCc
mt/dXxBqiwr7bsneP1dmZCp+TJGQc4uLLFJpymjybCLwvGxmorZkQrViA5zK4/yU
OeFt1q9XLTFrYmfuWZICIIQb6v5hNbtniQVLgtoITlyaY2pmgM9dBiG3AAwvpo7y
4Ud714vmUdaUuxj4M5MrAiQcq2DkVftmTwHkrwaseOzU8XmKi7kx9wvW4w/o18CN
PccYKbPYDcK7ZDK8GIKLc9dSQb6Mk+bUxU4P7RH5BUx+5jborDGXHHqkJhurs3KT
kZv5QpiP9lGx+uhycQ+5U7G7IpAOD6dudUq5NxJJ4LsH1tJVUZnYGMWmqzNEJN7p
uP2Cy7uGlqOG+VdEfCkscdBIEyuRBvA9hPqWDSL/hLUuGfqm0g75fC1b5j9432h+
mwTYSE2DeBHIqf3IKIv3IRkDbxcOoaxDo0PFwVV4JCz7hyTMV+F0m5jKBdRMOHhM
4myYy/JMC8oe0LfNBb2wIFIjSlH7+tGKZisMfbNGQsZvTR4FPu6/gXuzowQo2ARw
rLLdaQ7GTMMWctJC8NJTKAC8A2euwY/HBUxhdOLGT/Vj1NjNLAMqebn8e1icNHPi
mlGVqlYrP2XJrXQ1SFuD+j0EO2cKF2kDqlEQFKuq5p+v8hCI8eau8dW/fQvA4Zgw
0ueM1cg9HsoIeOmHYLY0TbUkkg17zjebGl5at3fajvJ0e5IBxam+J+jwsD6H0S3L
22r1MBVo00VP2mi5H/yXT5L4Ret5dg4c45Kr8grn0PSPbFIz+4pjlDhRyBCu5T+y
eb58TSDAIJeHJ2fJOvbSfyafLetJaokm/lgs7IezoVtlnhRN2IB+VDi+NB9BQq+Y
m86/hvFhwKzmz0OtZkOAg0VenRP3BmphVUJZCRKoqlFKYujJs1TRZwTjemT+feas
512223QcdjCPyGB2MGgRssJoEFRPGkpqVQ2qMinB0Y49+dW3JyheENQx8njKA/mA
rXAolpc4FWntk6mL1xTKBejERP85jCgZ0A+khaoEEKjvP4rL3Oyg9tL4AmxAw0JL
9h2JgSC0Qj8ok4Uw4Aa/9YEJIgNAOQWHJ8EynLnjk7JAy3CZCyqY1866Mwp9Z4sk
N3DVyqhjAXl8J3d9fIecvgaotQWkExRVc/oZFxdDd5PlZtDbmgKN2u6SdHXg5+yo
t7FjeorA9vv6uDpLAHeqLJ44vfjPpokrgPGubs21GUtaltRFOcWYby/sW4LUZKDQ
/mf4d5VucmRfUTY7i311oX/hZx252fNkMbvN2ZebnSBeYr8L2n7zFUJ7iz+4fPNM
G+TKsf1f/jG+dqsiFDFoL2IDI6dnQ7K9n+6e1Px3gavdiofwzEmWjQTlZZr5J7yN
2e0kX7yRqj/uPkAykZW1SlAaFwm8J8jvFGlX0baqOW4UKXKDFwmf8gQPEY/X0QTG
7VxXZhwSxY1/rU06MGg1Y/GKLatbGFX6UKgB6CxNrD2iIFSaRJuFNDQqHZXVHL8y
cjvnZzGmGKTHfuZc70L///6QMNIIT+hC6Kc8aFhCmaYdsRtO2EDqf1qKd8M9zwji
u09nzdmgR0+FQgzVyPso2ZsNaNjL3C6+m4VjcXZHGNbIZ+P+YPt1uvJpIPJ1zsXs
H5cev0CkMvHQ1z6xDbUD6DKltKgZKfyR4KzUAgqJvQG6gJeTnSenY+TkvzjpG8jL
66vqtDFUqBGV/1PFyEIAa7CDsP+VCWUjaNGm1lYrOat8AEXIa+Tew3vWPje6a9h7
dRNyvBqc2+ZQtEzpeEQfRURbrs4VNyhXM9KWfjBe4L+xl81upGwGO3aYi9q4IxOI
36zynZnN4EHi2QkcPHnQuWQf3It/iwfU7+7kA2kJWC9Mbyktqqkhszf3BiTLagMT
JsLOp57QJegNgAaehL79oQmVK0f9XVl/PM3iD0jNskovLKbLkWgvj4bE6Rm/tsOi
2pBqo3tg4dGPaNlo8d+Mf8+KhlPVOCwr8KqQQzk6KerMQaUOHNhZ+DJd8E+ZVfJp
XpYY6oZ1GVXYvZ+pLxNuPacaCouLvBTAcG4i8/RxWBVNGnFGNhdwPqKCHqNnxxLt
6wMBChF5Jwxx8ReE9KYPLJuHqruYrsF23ZlKSkt/4xH+5wONBZv6NdkZy5/z/eZD
S8KO5m1dcwTlGhOP404dAhUJ94zoVUNdTy5NXNMIxImpygdp18vspsgh7Ld1FcTO
voM3yppEO9UbBOd5RdGZ2QkgrSDTEyMjhNC/gTbK8YW51rRfxV8aq08jcNgUH7n2
dOQfAA4CCdsmyfeTNSupPHdFRWpYhUeTWEqrYAPu68gHgKg44pjZcBd9qWSQ2qkH
rLMgCGf0vDDf/sR6j3hJSFs5jXshY05ndkFA8fs15UesyS4C4hrKXs1bWEl1fSXU
91bf8GZfXAx+uOg6VGlRRIy5OM6GK8L58MCdgiXzA6Svsa0UHLyjeQNbLChZW/n9
HI1nfiPkwDZVb0G3L/kiCu2HCWxXUv8zgh8A9ZTewQXbCVSmjUrIRJHEJDzMCzZW
YS6qzkYkWp5h29ELJ3nQs/jPEDyQx2jiPDcJZ1U1IqEJyUDAY7IsWjQYtmmhBz/C
whNaq+AKb3HDLUCqfhoxZ7zsP30omhpFbIDReyqvHkFiPruhXqhd+fCZFyfOfg00
nZyxc66E7uSb4H7b6pJ6FBfuGM+8oklAufdSXGHYfi/hsx3rFqrK0b8wc922xud3
6lxgFiVuYj0xvg7THSfvIPGjJjPJQrOu8aw3vpFCgsDFoOak8HsdZb+Uke0puIEN
ZbhoSa1gJz9JsYx7XYz1Aorf9+mRxYK1WWLFTioRzwA8gIP//p6Cu9wl3kfeVauT
FP8KJ5SUlg+TcibnvMMvmzP1dAOsS/1nOUV+oHnxGFjDXmIqfYhZ2MjiY1A1HPP5
GhkZbpddj3PrB7Np0xt0N28E2RP5P40gDEhrOD/HctjXClZ62C97nHm80A7ENJ+h
apIrpRqk6w35A7rdES6F5BktxRoJHocVffzJ6bllpjYwKEMCQ555+SCXE16QyaDF
RzY/YijIaQVc3mnPQgZ7/cPMmGj7rcYjG9Q3v04RgF2RuE3vCEBCYHmXfPL4UGRT
5MurTf1rKLbuVGQ379FdsmjIQOT75NdYm79epI70LRDgh46mK0umI6j0ltrOY7mY
IxTFlV846pum6e3A0RXqR9/s1honeHVpi36SA5UdvXOWtbi+2HjkQE7yQcSiFk1r
/KJfBcXU2MjOQUPNxeTgHissqkNx39Csj/Lsv78/X3TEieXAuszScvwtotxE+FTZ
b/wp1bRUjmaBtvkuoqq/kMZ1boQv9njrHuhIUVBRCgbpnq8o1yoRxjFMnEHIs8Yf
CEZOay++/FHYnI9TnWmf8CEiojm4Xdl397oij4QFUgWQjpsQKn3ghrB1Khp6B/+q
jqHEYqY2Kzh9z/9eZwLDGeYfG69sgkOPy62NFh8eyvXTPWTwnGh1iWTsCeJ0RGX2
EqcFo1sz1tR5wWpPdPnPKegrp35DQdzJIgSfTEhIlfpyupJjP6DUjXvLk0ag6tCJ
XucnCCt6Vd3z0LfQA3j3HBgo2sn17hE73BAJUhKvhRiugSB4qAO86tgG1PEg7gfq
D28eMm86s4Z0UfUojGj9Pw7Fd0ubUcIuXe8IF2Y+I1xULK2RoyVNV3xcMgyP3ii0
anif7g6IwcYS+9f3H356MSd+Vw5hCEfnoCbu2Dnwoh2eOzx3BKyZqTs8bTdc9A70
Fvw+T8Q6mwjh5xiRKNsjsu5qPElTh6jFV6M3NLGF1UQ+nwmmjfh8gY1k4jc5FJs0
0GgKOUSoGlAeXLWIVdcMRXgjb9fCoxzI80QSAsaXIp1tN9ql16H3366p0sdgvh0s
3tq82M4CAJgMx5qkzykWv90eqphRwC2FrDUEs9rotpY/xXOpMBan2ZCrirpMR7x5
L8vakTiTtPhb6fLyvoolZLqWJJryF6j3UILBKUa5t35bVcuJ1yrZVs25lAhNf8Mz
2r6uAmlYz5uGVwoaydCga+kzMTnPRj9H2Olju3w3Fniz8G93Yd/R5BCqf6gjHwDL
sewj2716ZxISESIJTzVU/ItvDJP+TW8k059imBdtAvRHlpgIUxrX0B+ZMuuDcJGT
ruDIDkdZQ1QGwzEKItXzA22KBqzXZY/3sG9mc3ikMaWaP6Enszoxd+PUoEE71xC5
xQO3IxQXpDTw288YU6PMAtyrz//3Q3X7b/K+kA0++Q6vuhfh13xE/LrN/jhtX/KF
CQceWQpHBLSEjiDu6jQZ5uQFBMgBOrxYnWPi/fp+6YMSMwiLanbbyzGiZkEKFIDg
T3pNDjHIejWH9Klwl3R+1rpmCQwK0S0KOLCJ6CxvfmYsNkDeWiBFMBkgMR5Ndthc
XSGwkBqnw5SIFkmGYCoW9czStehE4mfRjUhIMY7fayuzwEeeAGeySnru2tbWPHGr
QUvvCAp7usnB8fx2I01rKze3gr/Xa8i4fo5GuCggXkVFxNLiR6bJypnGINOKiuye
XwqNOgFdIUJDVlPQNcoGnlScpetPYv1d+94jjqVQpSxr1CWCpIWD8OpOxySXPJ7y
hq6hVW0qngKxON8LF+datnRR/P2fpKFd7NQQVMryeSh8rNtf2bCJHMMtCn3Z3fAr
ldrdWQFoxPUk9W2/KIVenLoSrR/ShMF8TVXD+j8PelaqU/PfvaR+YGcUluWNNUsp
zUwlnZ28BiRxtXmtNGyAt5cgISGR3JC7HurdB0qMzZ8GtLML+MlNaoWiIhwbtNCL
xiaba6MXTO9TjRjC0sxjieVIzlBJosM8UKHI68QuRg2SXijz2XMyBXk+gwkcVPrP
1izL0y/uRAeeEJf6Qns1sb0wgBBXVqPC8+LI5wApcyvFFjfoNIQm8cyas3Yib6f0
Xjg4hQ21V+dLdOzvUnQ0ZqNw/8gIsAkWXT2EUuWse85kz8vJdO9PQJLOOwKJthoV
4PyIm4MxFP67vvEfAdmM7l/QHt1rr0RswTi2ClD5AyfC4hDe5vejY0MoynJMwAgB
ESht40iPh6ZvB0sOkZ9Nf90wmW+ebexd/nGixp3OyYP1CyWOcnLYeqttBq9DUe45
SpDs56pw2lBbny08iAcfyHYNH9Lxhp2vsXLaFyKPE7ZL8BwU5s4CkR7mSmSsZuM9
W6sIJnQIjdPoO1j/pdlYiLs+fWrP4s6UNrFX4hH9gl8tIrOnrSMwsKD8exdPUttJ
iEJrvK6eXvFHQw4cYY1z+nQpSezijffvTvS3u8nHL1f8iFAwtAveCMi8YE4TIJKt
NAgzal1nTparR6wBG37C62IM7f1R86+fVtn9Bb3ikmghC2DxHz35eaeUWYlyfxAE
NRkWz/xRNs+ze9y1nIiFYbS7IZRyoDMVJGJD5eqm1cXZ+hrh3zcnlYs4hw9tqsB3
W6Aju/GWzVS8bFmVKLCEv8yrBXHYnxsFu1Xu/1Jt0k/8Ir4n2lsMFqiAjd8Q0clV
HXMpTHVLuOqgZu3WVHAo1D7SZvzDKtdXp9bu/XHzuGn5fAtkAwcWFvq3QqlhYiz8
R74c9HXydQ7JTFtFacInocgjP7R15fB/nGfvu6nZJ66I/esu476ObZd//mYM4ysv
4YSaVfF3odItBOVdxBID2sA2vP7bByyBA28W1Y0M6HAPsou90iLTp3jjpxhL80wG
VaXGijFTovaAN9VsdgAO/z81KQzE1uDJcpNcei1u1M7UJso5ZEhXNmtKTyMw4ku2
QUWGi9R86JZ5k8VcRBo2SPWchRbzvq1jNsrhTXooyV9Lwa+ak2lTi+GpThgxH6K3
b2wve2PyeeabVFI2OrsBK+Rmbtyp8Y88+gqyDiHob6mFpkEiUtxSt8oOnT9jOmAI
0pm0AZEOdsVljOsAepn+z2t1iPVEJstfeM+EMcWjJaywtqqqHwHW72v/5yODT0Q5
OjNr/MRb9Z46Zink4qykoYDo/8b3qJwC2UtAZSr7tYR24FkRLkldTNahN+uYS/OL
NTaghGd7q0zdJRc949TOIzOy4/YNF/Rlfoi6YTe5VSPHOpuK4LPv0iTKoPo14gfF
N/6i+Y65Jwkzev6Ccw49TZv/C+ygQLWIAB0qMlp/36kyOp3RTM+NTb9wbnfSYjJT
JWVWyDE6IsRZ7KyP3Rkj08t7wepE9zfeI9p085M96KAwRFwpSJ7wd0Sy3uVIUakW
dBFuMObbX0AvZ2gi67sGmUjE3EfATxNoP+31je3Tk072M/vstPBEDjhtTdaswR8n
SprAdv+dsAF5ssNaYWkaDAPb8J+Vdg3Kt8w0qpXnJBVpxxuxuKvHQEWck7mLukr8
nYTQfIFVHMuymf+AX+0W6FDYjaXd6JrR35pnu+BwYv0OfsOFnum/tlBOq84lKcOY
tUhp/QBcx/uCg8QONoFBkYFphECT5Ea/ioXg5XOQlksWT3FE3U3Tyaanhnnw81rj
QdiM8+I2xxw29K9vQx2L4xBQHB/m8SGczEY5pLUtRSiL4GAht/Dq13fF1KPqCqYJ
KRSGrq2ib7x/9avhYhwHL7zpndrA8rEg6F51LTFMFag+uohFTs3WbBevqRRZzcUE
vYSSXV8ewHkURAqICDZqAEohTu+KZn4YBDTNDZ2yKlb8OqA9N1MhWTFVNSGaTzZ6
Dyc5F3lqA/5g7tVHhY2+uRHB5COoQCACJ17A813lZAtHCl20mSBJzfl0B/sjXsAW
QV1diWd3OLc72T3HKFbKxWO703JIVUsQi4b/7+5TM485iW0aJtvLbaho9P/m09ut
f+KRN0xUysndtGGmuxD7PC7Ma6A1W8J1VxIe/Ed2Kkbib8F6LZeDnCktM/Eg9MLn
FszrvEWszRZRy1qkhK22ZLVtPGHEb2ELp8zRygjaehfqfsBxsE48Qo1h9lL/DKVk
aN27PNOK8g/ImWogL7MzD1B7FHE5Xa5LzNZwUjDUcAySMXhpBdXxC7LapiVwIa7d
DoD7aTEnt7YXNHEcTmlRom12dK1War5czNTblT/zoOHPkXh89XVeYmM6fpW+ghsr
Z9JS2ECKTtGJ/SzyyeGSzZrmU0lbddTW/34MY/ynbvON3mSrcRIhAxsqhyejLerF
vcqMLtH/WJVJVDij2yMPwEQ3nFxzaHd7b84avq3hLlL8Xelbv7NzsFiTXmw61ZQp
jz7+k0ImB8lVnyF50nrZ+euHVuT4zQbb1bfCie7csAwMBN4c9csS0Dws95rCeEDO
Ssj4Z1Q6BiDHocBaNTygKgy1o+xPLhPHy9RJpUYx2qm83nQjUW0BvQp3Ipo+UhY5
pdLuOTx2bCPYW+oPoR/07aNI5XiuXA0j2Kcg0Jev9xFu3sUmkFrliPmVza2uG1Zr
fu5tNRYbcuxCWutOBlwU2hhhQ+LEjlM7eRck89vUjsaxFjxPqEnl27ueXWbBSsfR
vjOCGKM12X3nMAQsVcwDEAfv1vJoSRJ0yT71NU1vPW83nqilg7U9CTwCdNedBEDD
Nv+qW72lNj1JzNNncdHBLKrQjzKk8zNw0qd/hLgr4fyIYFQ/NojyHlWJ6JxOfapx
QHWqCdl4at7EF+/B0gPdIR+l383nVmkCeGjzyhKyZs+GR6TRcaMnC4eyqXyhPKlm
9cJ0FS2THfF0Lb5y5BsoABFAgvHzZkpdGL9qaYLRHUDg9UNjSWaSCFdD6pVTYiKk
JJcW+e9cadrxD4lCvL5yjuN/A49CO9UEHN0Hu+BMYOjFYEMH4BIjRxOOOJvAF5KN
gEdtnV4d/DIcdHXX+EtnHOGNZns3awva+IkBqUF7RSL6rBFM2mH3jhaBfv6eUFTN
6TweUl4ew0drU+zTQsTP7k+231fS4b8jdwAMBnRTHM8njrNQe1tBJAgwxE/OnbK8
RXipA62No76JzsFXVbDLBZ/cC2/wIedwcN//bemYRh4MksTaEMI0F2ByPB+/LQ6x
GmpKbDmcXIPzXZ3emuuWO/RPhrDEUlSK9TENzlHB919u9kxQXA+7r7nIXlBtAEFe
JEJ/pNRHneuww90KqTOesTuMNTetKpwrd8/bLk49t+OWPL9R5YkuNiDWQNvUCaiK
Pl3ug81xCGip4tB+tlC27mpNHpUzGJKD6UmRdmmFi0xK+e6jGR3qAthgA8khxcCq
SjoEfsC6vYD02STz+kuaJSJgJciOhwR+WlkCzP9EjVmkJhpPaquvXhDIcRkhf+E2
dQrOHxqZ8iqIkpUmdAB3ZtIz5YEoc2xN0HObvUmlyaZWdZDv0scuYovpAKMrpjID
3T3iKacP22NSbWTBn6qKu9+Rl8VZdCo4X+XuD2AgabqDuY67/wYysv+h4k3O5iRi
zO3m9yShE8lmNih47Vlt68mhSDvQZtGg6jmfGUWn2eVVn+MhalSQ9MBnBNiWi2G5
OoFdFLGT7GZgg8qL7OiZyRVreBJoaHSeWrCAGjclPifXMVzu9f0onxo0co3FjkJt
LBGZho9ZkKn9OL8bVJ/piPpHjZj/3qQIFaUt66jEe3gWEc3BAaeoKyeqSip7g02H
64smS8N6s2nT/2HOaBY1iGRnBKsx8jskYDl+RnOpiiM8JhgLdP+B8Y1MKkXJ5/bp
RUryfVDoJoEKbg87KRP53Lp4WHBvyx044wqS+4tP+4Js3s5hJ0YOoZW6kQwNZR2v
WiMYKfZOmG0m/ZzHsRzioaoFuVtD0nMYHYEUYNIojFloBCTRUeH9qYH96QY1lehP
M6EICS/ZY2PE5x+k26Sc8Kuos/aJ+Zonp+aEGG60vVMovtkLDPTzyzFMCjmkS5Fv
kbl7xIXuNx4ed+n/OXfyxrjubkFkrE1qnbFslNYar8P1U6vBlfsDV9xFl42JWzsj
Dct3sFkRH9HnzT2HwJpPZCdiJqrs26czGLwI/4ie6PAM1y0pLp7ntQR8nR3X6CBw
dkafoZWZB7KFIrOKUhffQjH8ADJigax36T5qdB36nO3+PrmV39mkVdVamk548SDb
3Pl3t57Wl0+erm0czzVtb7vAjnjFS9nsL2haKDc3XK7T0QJFu7KCX1FfzBd/OCFy
KjPtB8coHCmwn8oPzNeci7y2UpYagBChSei7EfNWqC5HrBTFVBvtyYqOISEE90ur
r4FdkRVJKKgZb/y0uYvxKFEe16Rt5E0ytv1QJRtzLikk0HrYshsjtSYCKVD+sOg9
ZnUY197Pu8hxr9yLSqhVo6igjZpuAGfUxknmO0QDI3KaucU0uRioD+Xr+UGp8ZiE
uxrhkcIltdLOIUHIYBoExXXp/DkCKqXbEuhTQDguBPGl3pB9oC/oKQPGA7gF4ibQ
o4R5I34/Ns4rTfVWaB2XfbNl2G0V/cQtT8mifuJoXWIvygFMcmUAPADNWIRXS/46
s4yL1fI7yxDKWEc9mt9aqiX+qh8tvywNvg7E1D0u3S+zqB6MN66Wh32w5EvJkvp0
cOwqhFqF76hcSINshrq2kkFAZ9cCkTJxMGSRiuJU6hKdl9OLs+iMQnId2Qp62U0U
p5kzjqW4Isx2x2TsngOgUULY5PRj6HYRFC2+lNbZdciIzdkjgJ7w0XpJ1KVTQlAR
qZMukk4KaTSTPHkhWvIpADIsMoBMfNn8epANgKV+SqZfOzx8LYpZvHXLv3XoiNBy
49J9oLvxVZQf0lq3VbWDfFyG73EKobhWOf+Ye5kFBTZp+VrwFxSkRojOrjVi+eH4
usXN9+YTNNnYK2V8mvYEI1X2f2pr+hrGYrNqpqKDgenVq8r97+qTPrG4nXDxsq6k
RXPR+rGfwRXk//kzSVWCaK2HV3Lz4zEVOLI5vgGLirGNuy26metIkKkRJyefOY+n
q4h6AoZ/tHo8iWq0ZsEQaBiro7KHcEJJWATQ/RrkuBCG0JR5um7a03I8sw6wRscY
hkno5FZ2EYyLecBdGtXsxz/RuORyQs23YE5udiCjbNwJAE1KYSkPEPv6Hwrkfei0
CQtxwMLs/x1jiWvILXs6EWinvacRVr6HDShzuqt6J5I8XIPUSZswQe9XLNsgTjaT
8bXObuS3CvOuZtdCFHErY0HG7GNnOeWIn3oRdVqmTE4EzcCLaFrVeR92c+UO8GEB
Qj3bLKJJ5fQXdKhwZ1lFM7flpoYmQT9iQIxm9ZhPCv5f8NaRto0rpvqUbyseSdz7
5mdIIKfEQ+xnctMmuvmQY8NVXDZXWTVb0KYL1o5v2AjX3RxvnKm4FaZWzOxiKyCw
2ynRFUKURfDZjGzPklIDlSuL0p2xsNNPWxEwdzLURbtFGF+2O1ky1kemHVJVUA0W
DT5zz5h9LqSMyK3We/dsQSn7zD4nhm60J1U4BTAGP9+9Ra8lcDdaICt+SA3ZKqll
O5cZ3efYH03GW6lHC/UZKX0ePxxr9+PyGYaEizrTLWhZk79iL/DHOVwyz3VHqpwr
tg2d2mg9bED2vIKmkuX//g/6sLc1qlqWnuj0/z92C1erniBxk6W33nRGCww18Bea
M4Xv0NaJLjR9ZU1hIqaGMaJyC6odSEz1XtRThi5yort8GGfM6a1K/QwW1Hq2BINg
6m+WdUlBCecrN93UhtHBF+npSwi2EvEjHCxNbU9+i4AN2ZbZhIIJWmx3O1M2NmJ4
wjuRHUS9Hg7uJo1m40PlZShW1KTpYK1p3dtVNeCQEJQ+4KyrnzCCVlU3oaAx04A5
b3EnhXrPZKn2rHXO3rcChCgR96JWkkB5eDpVB/KyHJni+7G879h2cualqX/yVQei
iz3se/SGlPrMSkXUOAKFTrOVa3Cn/dRWjSHDtk7McqdMuZKDL7HnOs6JiqoaKEkb
WqlsYCZIxmVr/pB9ZsFD2zCp0QBW3NgiIILY9LE5r/rnb65l/Pevoyt3aEwhs8Db
e13EvBP8EtBKF93pHx2x2HH4GMDdafaBC7s4C+/CsNjA/jj6z3frI1+HE6CItpaV
DAH7LoAZEmsZ4Qb4iw0n0UKNmWqaltgZyQC9gXRnZhSouB2SLP7jbNRL3JtP3aGk
0bRdYpUYMH4FyKIM179jeUmyeH3eEOmmtJNS8hO8CS9MRw88WhcNLjAxo6mfOqqC
t2/MJfsY9bEr6uEopJo0iGLIiwNSt2o462lu3ubH7Jk26jM44dy7JHFLk0ZRTe5f
ljId9FQAj9UoKOYmEqU16/Oak6MCLyB0B01ppDxeTubfqTHEY/3itrje6nSMWAgE
/hu/LCm8IYwARObLUMZqBtfADV4b+wSH3kJ5DO7xWtfo/IJdWs/RzJyDathfb52o
ooKl07VN5O6VtyypOvQptHRbQx2Yysygquh2f1RF0GlCjkVA/FNanXCDEHmHQBWt
pByEO6mioND89O195PvGUfQV2vpwftIuVlXE4RigCV7p+2NTedYjmjAcF+upmJmf
KIOIMCpu8kUI5WqLO/M3oCCQPC6UuFdjUTscmfRoB7V8YT3Aeh57Cs15W+sOCliA
aQOqPXzcyGYQOw8TB8SYNOVsRHG6zHk4DXU4q9Zv6fkkD6LoEFOl3awh0Vsp9fgf
5huO71hc6RDbwR4svFdwwohOJoWC4kJQ1QQG6c+jEoQZ5Fmjt8ZQXxUVhQeEy4Rx
Zs6nY+zsVpdNHM1R6AB4UyflkSyrtlKJ3VwxaR4BBfTseCXPw9L3at2A9dOT92Zm
b5tpG/QvBiU+m8lfSeZxh35CJ0MxoGecSdml1rA/xAgoZ+3Uy8mKr4d+qTVqd41a
zS/NHowco/1izNYS37WfonotHX9J1OOmDmub16hw0rcgw49Y4EvI/qARUh6QJ/eP
4Dzwt/C3hp+lBevpa17jCvaBk/qBXfcmQtwaDFqLkLUOvEBrrQXvFu1k8QiLWFUF
SXDwFM/rRM5GOl577L1G9i0oVDlXXYKjiIUW1IxK8A1rd3E1PU6gvfFERTfKE2MZ
H2bLNIsRfobEar8PHuTmAbdUzo2XTjkdS5ZWIYwGSD53w7FmN1pvUOMoSfJRF+H/
/l9af8Jayp2bQsuj/g1WXY4Bwy5dX0B3bKghzX4zObImLxF7nLP9eNWu3gc9BSFT
qCBCaVgYUlpNxoXH8RVoHkHe/E0nreeR/lgcEH+8xTcsQwbqAO7hDgqTC69IoGEs
RmraLyrwksHUfLykx9CgyjXFHtBdijRB3TEiA71cZKEWA5fuEzfHLYuAkWx7Ovjv
lvpXA923wv3sGgwA5Y8bQFMzSv7edmiRkLdNH83xZ+aOAzwYIsMzfX+XijJUEGmY
gnEtO7rXuYSnF/YMazBvTQLyUwFDYeiKdMY7InIVBWs5oc6Ly983YZVQwdJCThEb
HZDh9rGoqNSZjfuKOPAHdadZ1SWapNu9frZCmExFfkUeOTNpX0NG9IQk7LHmzdcN
VYtIiImuD86EE7HQUeSCNieNBvjkI1kCUw0F9iQgjpCy3gOPe0EJtSEiHXGKbgLE
RBWiG1nTFVkJaC/RDe9SAmZdMFitmELvDDQF0bKAxFSdYdVc9Dwr3mUE6AjCW8ao
eA/9/ydyucbq022tTLetBj+zY7eUMpGChxi+/mIjdft9KOB7HpjbQAplhwFWQdwe
l3jNBybZIFUGNT8XqR1J00qdz2k7tc+tG3D9E9H3BQRcLbPR6z81QAU8dM8wRu3S
XtaJbxr7OUWO+pjz5sLilsNCF8ymJr9wM3DzOoDF0JQhL7T0aVIjjkm1Fw2fkOj7
j6aR3Pk3vN3IX+bVm9EcJY/v81vDQ4w1a+f3jCkMMT1BvHsxJoWJq7ifUoSh0a/d
qBpUJnSwzmAdSsqfjywitfmWkYKzuTbgz57eSKQXOGUD9It+HjaPkSn3eXbDmAv0
8mVBXS6TIZLL75tdFVJpxEV0JlSvKSvemOVl+eK0UMMsmXzVPEfWhwTc9LcOs5PK
Dus/B6lTWP0pJoYh2q3OWeAbHG7BsRZfn75t5Sxd+8pQYVB1mAQfatpR2cvLvBX/
Fgldkqgsl6fVa8Fe8jdxOeIiyIpQ+y8qBxA/e8VHhaR3pcXOheZ11cUTO7n4kD3T
mQgq5BBxJ+YTisbZqaSJGya6WQjBV8xt4muCqKgBLCL11SH3GNVi4muza3E7zJoi
aTBwyasMykwNwgbtU1+MQVYHXQOXi5I1hHwzov/KiPm8gO+uSxCr751P/v4CFNqE
R17Pqc4xqOfC7Cjed6744ETjSbBhtPaaGv8pDv4lppiPLk/DIgqHS4Lpuznbp9Ku
XBzQZLyo1Kx1fZziOFtFtixXQFrVaMqBwPn6H+pMU/PmHtVpkoskFjWAQxda2Jg4
8MRdRhYRs2SrOEJ3rh7B6ty87G+DTuq243WmJrgzXgfDf5YXg0IUvUPX9W1UfcOt
TFJbyzugkStZj9OxLj+OY0G5QrZfncj1Eo96/x+r1U3M5bo+nMrr9+aacuOW5F0M
TNuT/GGImm0P3kzuxJeRK/bcjLrOZoqmJ30zz0HcqeJGwTeII1SLiQU8avE8rVx0
dilISEgMt2Z3Jmagj/BT0IAlB2ltnZkHpV3NhpJYR5a9aRNp49OxecEgQ/zILfzg
iL7J5QdrwHZbYLKiZQcgP408+crQjBGpLr1QDsW5bxGpRotd2vT8o0Vq/y14agbx
LCr7ECduaHn20NE0PyKKr2lbwRJOccfpa4Iv1DJZyZViK1mdKDc/CN8oLEUwVFM6
TlLqYKMnN+laVdi/n0mrYdcDiIQhXU2sStH83Tx8FdNSvMk+dM6f5tIaRTfBQDwF
1KAPZq7FMC/PX8exJ+KFGuQThOLAHHUlcS1/ldthaJws2+ICH7ferAWTLZpS5NL5
zgX8NiOoiUeyziVf6Np63FpDBivrZzbSRXj98EgP8D7FPXzFVq3DQt3a4cJzTi2i
Io184TF9zXrxals07YgD5H4WHFwSYpTR6zdjj+SWc01fNUiZNUE07nQB2OzSBpaE
Lqjj8a0mSyZhZznRNdk017GdjmA5JXNUPg9lWWsSMD+UdiXw/gl7x21xS+neH/mD
fLvpt/Ur+a2fFaObFMHDug/YffIAW3JLaaXri2iPPhaaTR7lv9BvfUzCzMgI43Sc
O2uhf0PcYcuYl6c2RtxFvDEyokL0y4p333Si+OEgKe55jjwJudBa/OIO6l753e66
M7QeJ6exu+g208Ec6tSVgb3c+JUUolk1AXKBS7aA3PkunWAEXg3frOzHXgeHvTaC
2uyqQHctedVP0iPqOF/HycbmuPF45tNUFXE3QiyBnfUejOGJwWv015ufQffcmvC7
/QsiyqYh9tnNHryXIK5nJzIFEUeFNR3iJtLOcWAmLuYi242sXDq47xJCSDJd4Ofc
7VBp6Pg1AAj2Zp0wgtH2qRwZhrZIVj+oaY7gCZz9BXe4THnCW4OFFYxYVRSfVJ5n
TOZIr2ayM5PbEnbtn9v8A+x7/NKZsQuRnU+X9OUUvBLyayg9jIaVvegMioZ1TbvF
dsPivXrEZdl0bE00mymlhT2Kkh+xwtQk2em6pbC1734zJShKH8Gri/lZp/nhD0VC
Mv6nFxfURiyxLSYER4HSJjfvuctL2X3INI7uq7yEKHFA78BotZZDibl0gebHfEe9
I+/NGBHQPxjXoUpbh8r6sXu77D+ytyvgH6+3pWDL1SP87uqkbHzSfVrbPj8Kc2u0
s30xJDpCFbpP5KCPDa6Aw57ZueNkparWH5E4lD7asenQuxkMomVX04Mffs9iIY79
W1fJeEO8hvgbU9MyrZqpizdu+e8drmkFgdU0Pd3SYm5gjUMNOXon4dhNuUdjjV1+
xLBazUp+bYWZlE7+Kk+KX+9d/A7cp/hygs1h0tdh3SZThWRSb0UVGBZhBslz5jnj
ZrelYqWQqvy/we2LZTVFmeeTub+Ryf/u5LZOVCoZ0+qBxVo3K1jqmBv9f/SfFXuv
kIdIUjKTVro13LciY5ezPBkA4sZ2nmzHMpdyKMIjdNJa/1Gw4AWyPptmmM1OmES5
O1HFRby4n/Z9rrQms7kRvFkXoIVakC8adQarJMw0ClazY7pDGIm/aUaQy7RQ6Y5Z
m3ao0C2ZxOOaf1t5ScJl/040EEtr0DiovtOF28p9JYEOUz1JwsM2+5Uko/gRDm8q
SYg7GFXMstiuCA08gcibDPhq5TLvkpxxceW60Q9iM41NLC1Bre5+RGO/YBhear+b
htqppZPAqAZAil0jBQMbqllRxVpCoSmUH8m/XIKT+oQvdyNI0xm6xxxG5aClMp21
F7tLN6Fem1p5BZh1jzJt8zD16uTBpzDoIiZpaR027afKTS5dVgrKslmle0UTNJNs
EM77JKo2UKyY3xF8Jf+JGZ/KpIXm01rvi+BLNuRh7sgHF2l4Urr8Hjes9rvwqq5H
RKASr9YrPHQmIK4wnKNj29igVMBGTECXfDnuBUOmP0wG1g4fKSqQkfL2CQG9d9YG
sfqdpz1k5XWSHLVmDroq7DzkJTGe8A9AZGmfqP7XZr30jrPGo15tzvaAiG3pLveu
trsPkflznprQEC3/tqH1KnvSBvUZY6YXzlp5Ghd92pYVVUtlYv3CLfZekzBMuPtT
wnMmdJmsX3ZJABkgv7tKzgR+BhmbG8w2UXww3CD2f/LM7FMbesol/Sln6JGC+BGx
/XsJANnIHkgfxmsjPB7U7gZiVEz04vDkijRUVch65fpu2bn8XbuZkyWW9G0DRKxt
Blq9HyiQVgQ04BlDF3alE3V304MbWF6cGbuT2dYm4eN6HOru9gtr37W+UDM4snzo
OiA27Ay2R2EDySqqG4ay8LT2WjuFYdllfqXDvyeBJ69hM8dJkN+7Yc5UTVBwRQT7
WGRIsmzTFg+Vb2mHTIRfZ0F+1qq3u/ru21Gsv1ISywztJqG9rn/eJK1m/SvRJ5U2
JL8qqRZ47ITAaT82eIODuiwp+YzJFyvCaCBeovPywLSLTCpflmanKYAEPBWlj1Bj
hn00b7bqRdQk1HX3oILDezhfEnUy51Hi7JykQMpFpePpHRcJIxEvm5ioALhmIS3h
9NLZ7p3z/eFInNsULPsRydH0YGO9OIGQiffH4FgeU3hnsAQUMF2O4Vo5Tcgmz6FG
9e/4SpElF3fKJiniplUVwbuH373NIT4WkZecUjYGr2gDyoJlhGoRJqhPUhCI1qJW
0Uo8XvQn5sKJdLrAV8L4JnIQDGeA0C6ogKY0OM/3G4k57wMmNT2X3ifYa8aeXS08
zvbKhaBmLx6UXjrc3kMTSnDzPUqH+Q7XfQ9wCHCLx8bxY55197PvDdZCqjHOKd/b
yCxh3kkY9/gGF0TjvCmxeKbH5cmCuBjfpyXso5aaF8Cd77nl7aFINpqwY+IhaWq7
pObq4lMJv9oPy0JLaBglwlCRxxJXq/k0iJzRahVXOGY6Cf/4OIazoZgX9Nt9a+WG
N5gc7qY/1yVb0ys4JO7goSdFgFQJfxemRLp3FGfjPZ5k8O67OHVttSCyHAHsGYpG
giuAIzeGmTxGC9ghyC7BnJX8wfN0B8pSIf5Ie2m0sIlq6T6coLVjsR3pNV0kLlnM
tNFKjDgnEfZYVURMamceiiT9yT76zwTfVHyYhyux0ajxjzot9UqRmwvGvn2EANqa
miCVdf/QDcfxG58VK1FiBj744nDeRN6q3lgcc88h/sly0YR8spqHak99/EB6ViA9
pzYWPHq6eZTU7T2plwRYvRyyQF7E+EWn0cbYVK4tZ/5I6GffDJ/sK37fshm7TFaK
metF5j1W1wGBpvwJ7T3LAoY9Snz+oufRDkGUuPgVMZs13vgHlpUvj3SbS8Smx4zC
FiyNlofibNV88krDyvptUKQ8F6QL0lEHK1bQQI9daAb3BlV95bjM+BCw1SH6/zfe
IRNwd0PAHLvXEdRt6OL+UIIGywNlaplBNLFVzge+OjQ//mQx9eqesKCydo/DziKh
M0zE7tRPglXH3AyyJh+KW1IY2U1XnnojRAPvlCJsurqgfAM5uuJwEJMxK7Mhrvmt
6jlzgVhq7Uts5mvSBkOdpIAdMhU79w1G9wy9vKvr0hX+Onc/kUQiOebcJGw1hf5P
STzFVkDW4/YpJB9bgH660n46x85MPaUeLRiJ5CXB5YIicESmC4fceFAZOID1gYA3
Hkgs7ZQySM8+bQT33q6TeioNUC8pVxWF2KoattGgFvl3mq4fKov3khUKB9Mgg3Ta
qQYoe71Czd7qZv5iGcnia9vcDbbh6O27rQAyV/HM8cm+Gk50ohMMbBbrjtfVV1l+
zZkQ5oqdKLFmw2k7kpYg+8LJl6j0PIZOSOHsEFExi1LmmLnhgdc+DuLQyzm6Ecam
pweA+uI1IZ3m2f+KmQQeSpSjc6LQ9AEZZzGS2qmHpIvAS2UWeVh/xcDt4D9/wwXL
QhpwSYlRzFOas+g08S83IeokSzH3P+GyqswkULbHM8gKdTxiEV4FWgCRv+0LE7Ml
VtPIC67tMeS/nF0Xt5FCb+3gIMz3NxrBZNdtOjOi+avxKmHd67UFGgJmS51GA0In
7xwKCfkNc77ulakroZlLXBZblzvkwKwIOfoTmAOCsb96SuzJR9eFKRAvd+YeHb+N
dreB2lhnVxdTmY+SOFWSnA+dlTVEe6JjqrX8RON8/4+BMuVWZ6TTmRBVy69g/MTq
n+QpDL2ge6h+PGPeACFlmtcXu+3BwvdUoSyFmWN4EN2YlnmZZALDzaNleHxx1PH7
hACohpLdqhTexhtLM8Y5ZVk3ch2i6HXkwvarHwdVvXRkGogdmtFPcGbfvmIVG47k
s3cFRBiO3Enzp/dDbdRKxC9+3skLTPXAQYRZ3WNFpTjaeILMYwP0kR/O2Rp9Raq7
AAiYQ2Pr97I6HIGCVsRcy15W6LZBlD78bDGyMalVAv6BE2qSZVMAnH7Xav5fWBUv
uP+IldfChSZEzi+lFGuNXicU0aHz+n3++VYAN7E/wyWUaE/aT3LR7d8dam+tu8VZ
MfUC68MOrlnbZVq5kiBre+zPqMEITzMeUOXTgpfu6oC5Qk/28w5Uilx1PbpfNUO6
XnlQV3xHp1JZFwb/3kIvfFvnKRmx7WYQ91LR/pacrjypYzwFFufY1I69NwH29atY
XI+p/kdwMJHuxlqty43wUPHM6XTq5w3cwsYdh8SwSjdbrH6ACS24jLs+SDEWeFW1
eGfa/dBu5fNmwszyIk1xv0VhfmHqF5Ogt1o/tCCkKKLezwpU7CxARomBlKPna+3K
YiAhbTKu+77GOgEESUCQ3vPVp8gSZWyNAaiXWqqWGs8p9Nj2Hv5AViF3OmK2vn4M
LsDAD7OEhAqJq5uG526xjjuxfMbMirw+SoUAs3/wcTomPFolW7GYZ2CyJsdGa1qa
1yn0un864wL6wP1J0XFZiqvvK05hUy/efiZt8+biJiTs8kv66WYZHShPyaL6Q34m
FEwkpizytD0x4bElFY4kIv8BqPZzwJTtB8rVoPj7FgTbAmN8aOY0Tgb4FxJ3TmA6
PNkqvgGKW3OwAmLVbpPn8GRsyTpqPQ+tJCsatv1lWlSyMN7t9tZqL3I9AAtpmQ6Z
CTt0Wch6+MNsmlQ4OZyTV7xm/W9si4Ax+MP5DlBlPqzNG/v1q43WDms0+2OTmEcm
z2OMG1haCSskNioJRR7wczM+0P+xz83G9GdVS+e5lohGq2w8GptFn2VtflstGR02
teb3dL9C1Dkkz0oLBBd1m2apKqF5GuqfJ3v/cLQnyZ6AQQ+FfTxzwpwH8PYytXwK
xa1Cz/TkCtAyMzL990OcTB/8sTF4+tQkQbqSTFzZuV3rnDlHeG+uXXc7JZQ9FgOF
l8jdIFyALaohPIcp4PdZyArJYTm8YXC598ZOFr++BKWSOXMTirHIhBjQCc/G2ORx
CuEtcdGR5lflsJZ5Yl8o//vrcbduKM72ym05ZWH+hmQ8Ic8mVPYh2hfVqgEIPppw
7dWIwa4YYPKKjeS19laaq5eUY4JFw3SoGHSOio4GulXp9W/AxRUB2DfhWqbz+0Qs
ZVB0/75J/ghOF+geugn18waOV7RF4Y74dMHue2I33h3lbw4H/Vgltk0YxpHSQKBl
awI7fVESGICQeMe7hhdEcH5SxXdv2cTxQH+nl+oSxjeAhV6isQzB8AGYDR3qemSs
VKtg0Ew8IltpISZCumJ9RQf+M98SuYvRHNeMA3GE0P1gPLTWUP1SYYh1yJu9PCE4
n6AUDKq23AxZ4nmcEdqHHQJTclGWSwztvzi49E/oXwJM11xrlJxGcxFYaEQ1uYAS
vjl6PtgabVN2PxEZmTdOXsW0FHn6EpHzZQWWVdzaFePt+V4p4/C/DLgV+UTJDHG+
9uLEY3uoQThDoq75ZZpuIfEu05QHecFgmG9sYcodXymcCSa1bcoJN3ZPX50xt9+x
TnJMF99mQRyQ69etsls8GnC//XgI+/WrcnECIK8Y4o2X4CPKWz1QeQFdNbxDCNCP
HHISD05PIh+MtJkWUVsAg6xXqDbG8cyrGjJU/sW5kfbwl6jt0GznscDt+uzrrcyQ
UvhUrRgH6OxwAHNjdJ2LPN45OpCMAA62BpmizVQB+shw7Ea0VGWkL97EiHciCDhK
IeeXNWBgcp4hvcs+JBliuXiCOFqqz0Em71v7vNdwjBXrgxX+xaL80RaGjjvnv/W3
CnCXIhAan/+xSv7hMDji9c/uTc0369os8c5bKwut3fGDVZMuubb803udFgUfFx/W
0OKsXTncrjot0HUVRrmqA/CU0yXqtCS1wspkoM18B++iUSsvH7xm6IMN9VjU13SK
sN2mLOrZpXm1uWHeyb5AHaAz2WuAHyjCsTTQqwTiemD+IhNf7Gn20IorICdpO5wu
BQoxpJ7f67qnvlrTngF3z2c7bMpqpE3F6PsKexALfKPi2rkGnG5H8bw1nbJFMdub
SsZlHUYCxf2QIkhKP7y4zrjje4LjoEk1q1Ehs/RfgyRy6WQvMcRh0mICrOsLtPrA
oFw7H773OnkHP9A9AIU+oCXjEJw97mUvAvo+8peCFmM2G2oLKEoYBkqH12Mwkrhv
h5mDQ4Ai6ZidiZIEOzsshIxg2wr+B7jUovA1X5ijBTo7Zox8dJ9trd6Wx2c+gX9h
ztQm3cM7GL1cey3JRgHjOT7NOXoSN1+b2bfQDQ8Kyw5wYc5eOXzV7CM6f/x2NFEK
mwIYDIn/q6b5dTjLWf+dKdNY5s07HhOrq12aMHfu1621I+ZclusKuPxq7eRIuWpE
qi4fcZ15i/rgGKX9usut+Lfk4a4hL2G2peDkQj3VShfYpC2P4dv3tpzXYMCfdVQT
4xL2qzK4KvUZ5wRgJWJo/BOdaRNWS48H2wvrFzoKt/B4xNRyTC9c2HM3c920tgy2
beWNiFb3pj+Vl/DBVmvXVxCNHmMAqLrtRz9Gb1SbLyN9q42bPHQKcEEn/T3uHAPn
dM/WWNqjNbI7EGhRoYkQgzTdu6iMOBDFcvAMg6Z1LQNeGLXWiEOKRZrMNFFtI1xT
sYI/+cAU2wN+FmoBAWQiCmf/GY3BSZArPhNB7q8PgUBC6j34i7YJyDQeU4497EtZ
Lt3mn3kpMiNnCCL27AZHPKzu+7ux81DEGXhCBu1RtQUQfBKPl6XkGS3ovvMGN7Od
uQ/QR7LjeGw9+rdAArDj8omDjZa17rzWxZOI4H1nOVwaH3djlbIJh2qgOPoC5mMf
SrNkDewB7vGF6kiIKd6OY29i3OoqRe77r33z1fSmT7a5U1jxYDCVQcjwZ7UwawSG
KSlshfgfsHPxjtbWZ8V1tz5RpSOrYcoJZ8XrmxPQQQKWZQ/GiYum3dUdsvmO3ydv
PmKHhdaOnTwTHTWyBbCHtrovicogudWDlFYZiuASRgTzMNs4psFgLwJW5KmunINd
0r6cUAXqmq5QOoN2tgqW65/YJCgwrsM9ZWF1LpThzQwKGJ7phP1utgJsw2zF6S4k
9C0yMkeHBz8rKTdRqI98R96IYbGxG0DPs+MrS2clj6P/QOYtp21/z7FGxVD+13Gl
0bJgQANFySZfy+T0TsXvL2ebCNjyBA44EHfBPE2O5mADsfkT+EKeiJonF/4wRh5R
62GFL5pHhL6RxFHw15a9Rc/7TFa5gkTYtWABmclpKa8kU42T8PKpzyTdgZy7Uy4p
1A+zD4qVv6LqBMi3Iao0BLUvUjdT60eWIU/gc4dA7buMwa8BNHJZyN6TnMwHdUBg
rNv9+S3f3N5LFVFI0Sy/GErSq+CgYfo0ympD38NqOvST52j8x/Ljo5LigDTThqjH
DbjQQsV6uHYeab8XQtYmm4SceRNT8BIYgbzr1et6Pgs+h59dnLl3lXjN4kOKhel/
LL13eeeC4oMpTf46rGlE/E2GJYM0uXzmLmnqNUEBkrLpc81jdN1s4SxgxJkbZWhb
peZHGuh9qYpShbbn4AvxUBjsJlKXOdzWDIT4989kcbCHgKEt9ufLLN3XT0gLHzrO
RMsdZVnyhGDVYZ/4NS0AqUMZ58oiSeILwybc4GWHioOrw3lI2MdNlC3dAbYX9dVC
kMfFz7+fYN3iP/k+ybkJ7eBBWF869khp80ADxlkcJfyFEmtYsOgqQsUkioiGo3JR
oGsKhh1bAhWkdZt32qqaNSCHmwaUpIW5ZZ7Inp7fmrqQxjnf97oIJHVSbLyx4rRq
qVDKP5nGHiEAKU1B9HnqEl69IIB/sIvJufk/tUERJo/yizcxtpqGbW7rA1v5eHVI
dsRq/0fapb8A+elL5dmBWX26P4jXiM4A++BWjIIt8KO5udkD3TeAA2gzrGUVvqVk
Od27t66mgeDn5WpOQSgePQ57JtoUlytZnHQpV7RWhPhRpRUSpxzpVWchh+LNAtkn
8JgProOw4YJcDcmHlTkdQabWl7YZ7bajF9JUJ0zSSnOpsj7SV7raIMoAbPqtBYGr
lt4eDFeO+BHKID1ZjgKHRLw9Paa+QtvFOeQzxrpQTPag9PtC+1mZe0oZNAOK3zgU
3RMHm2VZeeRT8Wwuw5RIhmWqKq2f9/zuhx+90WWIpyBir+ZIEkL9XHlQH3ONUCTo
2QAolTnMWLbRLiaq+N5T70P/Q3Fg8/ftY3HoYT/ReKzAhiNOdcG5CFxwsh2CpQu+
axPjmjZ9gy6EBTKVv7e+6HVtYyZk/Bn+GQySXveICu/jABhxt3m9/azkASHUMxLB
NwdlrHCo1TCbYYSsKmdGIN47MF+6hON7T27bDdrnqGV9890c92c+96Zvv2NC3uko
HRymSWGK44fop9Kcnbu7Sni9JA7QxrzXPjMG7/yqTR4ki89TQRnwZl5HnGCP4KtJ
9V3QxUI63BqOHbFXuMbYowtgOBHTIXsKU8vRoLw1W+hmr1wAsfgyU4XgtoYbnjr6
7i9lEzKgx2KSFKmbdfx3RRlgrfE4OYIGag3gv0WPxbJdqRZlmoGjPqxL2k9Elqs3
PIJfOqsU8aDhjEqVI0fxEblhIw8tmdr0jYK0jnJT6P52IsRMzeNAnTmaGSZLnk+f
P8h0au0foL6oznJc4wMpfCzeU5W6KY8vhyf5+/WBIrMfQmy0zp6UnBYLsabOzIV9
7YrfbswIAYiSrppLn24hRGy69G2gw7vz9jDCz2RLb3nDEbxW12NCpzvWExivLCrB
tahv9MAvXzQ/DiLLtCJuPQQv9MgFk2iFBQY39Lrv92wS9i4aPfxFyXPxDODel+td
0tZdpey8BhjOmQ3UoCZy5a9OA0OetOQqFHxqD1710ykAfAnYWlpzgsOW/HUeH61M
/Vuti4QEWMh01DDEEDY12Mo7OiS3X/L5TMRBeOxIILA38/Wp2g71fY3SKszJt2u5
HdJO7N6u6Nhu/BiVEWE3RFeyJkmiDveekiBrbDcpYEYFIv/hE3N3jXkY/TjC4GpQ
fY5Tdkc9RKas4FYdA4yIGveb3tDHdlIlRfxcoc5+MuBuIXC75tMpgOybg3Hz2grx
gv3+wIobxwqWvNCz2MPUEIJdAD9Cbl7mQupZ5pgp+NQQPWRnLqcj6S+PmwB30DaG
uiRFTYutirZevP02Chdckc/+s6Vvp/OnpajQfc/NRoieq5CqWI0shxxf7g+KltAP
7S98/uclBMg2aKmYXOysqVUKrRlNuFJg3r2QblI+P3glIPHpraw/AmYb06kXB3Ig
XtGB7nkfW3CVG7wvcFKhkOJDacSjvHxVw+7Zyh7PveBBsLzXHmk0XYEUvapHT2xe
5Ux2RC29vI7oDV6DCTpd+d+HjvjvGV2k/j8R9H9r/bwEKkzoRnEdlRt0a5SUtNiW
S6YWD/9lg2tNCGOxo0fKj7eRwAhBuoYsmzaFEi1E9Iqxv9ilGJdj0g3ii0Y4Yxwa
RnRBEYEEwDlGnEQWLZb6AEWhrrvrmP2bdnR2AlNw12NM7HreLeIkvt8uXBSWG/34
2rgfe6KqwFTL/cdI9K8d6glWVAo1OIJswaWgfl1RucPVch2wZ3KE/0a+psCodgnl
dgc4omDi4sGOay8GHVuhdWH80y+rId3ds9oVv0eIpNuQVJRSzD24ABzdOkOLJl7K
54Q/sI+eWjOfulHBjC+zIk82rGJfxTJ+Jy1y67ATMcMqxOo+u6y2L1xOQoFZrEYm
r5esn3BCM/zioUnlUduCEBLWAgoneiYUjV/DORNEp1FBwFsQa6MnGFzQgxxHqvUn
lgbbHf+pUg5JyopF1ALbzO9kdXFMFMGJExiywNPuQ45n9VTZI8zcYXSqCy2H8x/W
EoaHhjZANfIFH6Dhmjjd2cRxcSYS5o8eeglKBp1KqwT6t3TNjAISfwsMzNSLu7F/
slb5LAFyOY6xLAxFEoIOvVE4kCGUVpuCE6/xUfhKJRN7qKm5ZCRYtNFMy6rmLD77
8gBRHcHSm6Gexomz03JLiwasNvPnQZO6HrfrEJkFfrQZu6ZJWC+2K3mpYPFVHWB7
MmVauT4H9lEvhV1UR28jw4PKJlS7dnKmsajbJm61C7NJT6gl+9EBs4crhFLrOAAZ
CvwXMc3EuN8hqAa5oPY01NDQ/aXdmyAnKnFZ21pxW9FbwG4wsKFTFSFzkTk9TUAh
BnMB380SkJtYAh1ullaR7Zisp2bUkiMoOdneXAQY4XOx5x1Jnyz+/1xAaN3f0eew
b6vv73l5uDBoGiDafh5RtV4hzA6+wKjTCUENP1fscG1Ychv6Z1sNbm8c/7m+dcdD
Y9QHjn6vIu2G+0HOGItgVN9l9Kac2NHC2GIYRDBNRCdwM4Ua0a2+dGP6csMkTRpd
xvRNOhQbI0Bn46h9QlhBbsMz+MKOpWusAsAt4iNn6JCqMnA8N759iE2+W75mgOdg
q5o7K2+IIb1YM6+DK1psYWyrmLi4xMmMyguqIlh+hMoPoLzXHVYZMhYKqwDaq4Yx
1LMB/mdfHXwcv5ZfnR4mvM+o80FukwkGcPnnHsgAL37s8lYT8V/pCBakPavPyT0w
9hj+4/URrTS8jy+kk/o5tYYeZYd+7zdr8rkO4DJMhJQNBJBUcOJxj7vF70kjcgHi
hzY2+ENii3vshc9xkft7JTXE4VAZIzolq59GRMtBmU3a6kXvLn6yTQbsM+wZD251
N/lsmK/93U7DkRTnjzXrWuy+6RJ5hYY0zkSFKufDxU6hty4WkskiiEmp51l1nIpf
sNFmgdTY466NPCj63praK3dHXjt5n1JAkjWQRYfJzDhfz6Np763Ukgcv+Cf6Rs3I
A9nlFsmZkWHx15vxjYnf9RuCUMUeVXhKqa2fX0TuRRVxmhbJSUt+nlGcyI9kmgKX
FuMHlDTP/u4dqrWGOt7/QnjzG9aWVHFRwaNE6jdlIALCLZMWFWLHvGhhERs3na+8
c57+ly3I4Kq7WQy2PaC+bw/EMsbIMfAYgcSJKKLASQ6a8hNfVI/krJn+uQ1N9INj
GaIYw9iSb7LOfChfBh9/wHHZKRK0XhJQND+zHHhIykeZL1nsE57eY7qPjO1MOO6d
jMSId56paoOpbAe+3Zj4hLt3rBfJKtO2SqMtx4G5ap5KVLYcBWs250raB7fDcTdG
WsK5HSan9mRlEp6IW4Mo51DAd4TvaSGboUvPGKxK+Oin2ftl+dLmSbR9jpj46YA4
00kWNYeZrz9mcivddEPDN6b+BostWkSCSHr6BVWFbAu+7RT6+IVzVA3m5uEnkW1k
MAvZbb03EoQTz86rwXVIhUWH9+nqRdDA3s9YfJFIlzz//UZVnOfxPoAggc+4YCZH
5TwoI73iUXDkki4cvuMexp9RPivt5xkTonU4rc6662pb+EKyHW5+vyNXoQna6jK2
c4b44sumytjVIoSf1P6CyIAKM2vJ/fooYcym4YX7tT8TuXgFX9yYToCbJ1/CuRDG
UV3K7GMZAtxi6NozVOPGA0O7iP0t0vJlKCrYrMRBHTtdDGGOzt3dOCHYJLa5tugE
zWhTtdUwY06EQJklAu/yBJWNyDcxk9V3iPNyCuz5ZL7VpljUA3/bKe8BTThIV0vz
Q8GeSY4vMYocML9iQA7uIs22xuvLTX73hY7PCT+CeleOdjGsO2kBPg6LFbLSoXiB
grwooCk2ng0+J3emAmXL+qY3fMhwTEXFdivfLhIXbJ8VQGj2fHIcPT+s7e59YWHg
ww2EjejkD4IcApwTyhwwNw5jtWveklxsBJnnVgqpp7utzZJMCVOeo8qkPIW4lwaW
Aaj9KPAJwwo+whRXAzXnrDt53+0MUXnEGmlWvQkyvxh0RUi4YqcyLfcqF4f7kDvv
pLzQg5jHkmUDJFjJBEf0kpzgplmf9ClrEvdBxFviuRwtwi5ZVBQekH5BUpoY+6g6
jXj5Z9yHxgY3kUTgW991VOYJpxOC3devNBF3nYq/1h/gnnr1IcJ+01sxcA0pKPqv
X6QsdU3YJvj38vkj6eqh/UI+0cLjXwWlDe3OY4kSe+CZp/XT9TCngPnPxLoEZ/xg
dID5b7uvfGACbUGBiFiRF/NoB1Sf2Ej4u+Qgaxo5hErReFuoneCt7/KDPUe5hPd+
g+o+W8AJ0lfx2oayq9jeo2GuBCUWr+HomxIldlrRz3IRHmtjBQIzYzMfoUq/V70P
WQpP9y/tnFrFR9U4HFOsoS7rAP5pUkAiMsYz6h5gNGyTvz/xfsgnEubSmtkCP770
wnLdWOx7U/t7rqpuexmNq+rNxP0DgZCrj2aqOZBjFfhp4iQ9u+XDOpW5/Xs4JW9E
AdtDPAaZF39dvBVTi2QeHm6eZXNhWQtCTqFSangbDulhM0GOMHNWlFWtSnA3fIYS
2zMgt7Y5GSZtYE93U1JNhpU+F3PACtG5qVylyrdGEhAic6IY9fV2A85J38QVEtKg
ntlhjm+jA3xWdaLtUe9LMXW063ZTkewu6oE/uMX1cX/2+B5w38Qr052oZoPyAOes
VdcVcCpmeVy1tnbIivS/f6r1UHiB6NDosaAW3u/E+WpJC9Zg0tnDCYx6J8kw7gsO
Yyi5iHsHz9AgH20fVw/r15H7FaDmjZzCEeJme/71LkCqUfbDM/24my6f65lwz5i4
1ZcE3i0tUKPnF5FEvvXBdcETn50Mcb6Z7IMY8inlXl/ra59Vgm4vSzGtm3e1RVGL
h1hCEVfHHPZx46DtbUF5XlnGvTHCVGuQVXY87/6HqeftXtLD+loa8kW1k+QB4M8+
fFkGRs0AzYXkc6Wle7bofzRBM/zz1TBwK4sPT/AHsA8keZz5RIyQZckohnevC9Rb
n1VhC7f77Zkdttlamc2v7UN2/bFzoGHMyomWeGAjxFvTYw8RbPIlG+DQUbXDr4Pf
fC6fTVv7/Pmt3+QdsVIbhp2rHVkiFvaJW0ozkgM2qb6MgwKIY3wtlsGqhR50QjmB
I0S0Ywdgi4SgD/IndrvG6R5S1NrOeV6sOSZodoFoVvzGsDlyvPj26VRo/JBNVXdl
3o4L6F/cnOi+bJ93FYLD7F7d33NWhC3nnc6LwrkedUJyLC1k2adgtG3nIkswe0o4
KoqAPLjsf6BIdwUAEVO+D8Ngrp7/+zn93lsk3as/4JOXpPcLjv34mc1EGTv0Orkn
bi7kxZF01wfiBVW5HSOPVLr9MiHn+Qx2UDevUoVQ4r5orzlERHfJzKUNvLu41iDz
5v9Ob1xJIhrYN8bST4JYNe7GecOC2QfAUzWVMCuFRWS4i9cUlAlt8b7O2Gbm54rj
zRngTWcaRJd6lJTn2xLz8eCL7x7kvYfE8SYVOkTNR3Xp2r+V1Okl/NREfmugWs5x
OxuTSEZOjf95KPOi47lZBmf6m26XqPnI8foKB5zciTGXpCIyk12RaohsaOEDUN3P
v31LzFk/hJpnwueux1oJYiRwLXQpKyRlKo91pcTU+iFhgMUJFULVpEjNaUtW1A+B
lgqxsgFdvBRVAUmcnuvVaXbbKCG5CLDYvPeAjdciQsRLkINYkyUPeCyAMKG+IAC/
JLvnmN+9o09Fh4ATlP8GPJs7d5xDgijJxyVNcObTqzMUwJ9ashAqnKbcKzYGzOfc
jwCbmt8nloFeDGTf+sSvGZ3+As4IMN+lobeWrxIAtXWI6fcUDxiuIArQj3bbNQHP
Jeu6BejEHWqYD/cxzgbzvN2a70uSvF2hLTtbISIA2csZyKI5Z7F+bZUd8sfe66OK
yBBUVMlDwHiU4XV6ZxSo+d5Wd7wEv37gWFoyo/O7kJwO6ePyq4tVMso0xFzq1s46
bryfw7PcxUPpRx+SrmbwbcIPIzS24AVWtZcXhl+J9mFMxrSwhLTAjISsfVRMSed+
cPzE9yrEj+QY7ETFxh0zv3qHdsVuZUEsvR0pdPbkrFheNKCvSzysnU3TwRbIzhRD
PS2N5BgrC4IYJfZIpSpJJ50PTUgRc7YznVbYraUUu+vSA9vDuKpjTbWB8JAwH8al
rTMe14A7zNmKBMHG2xG1wV+OXdSUshSSFwjeYohYczaWBX3BzqHOlrr7+XMGlJ2Q
IBYNBPJDNBkWkq7wuSJM3Owz1SVNDoj6X+zMJ9EJrwXIFk0P4vTo28VI8FwUQqHV
AroQY1rSsADtVeVlyYCJl0x4Memws1+8csSvDNrrfq+l8BaWOxMGfnNeu4OD/5Hp
1IsVqChN3YWybaZtXnzeViH+LC0jVeySHnPYWvT7c7lgM1KYsJE8QXd8Su2foRmr
w2c/imDyv/MRK+n+etryX8CWM1PIyO5WZ6Wl3zNUMMhUilFfm6Nq2yoYjx6Azljg
W1qIJD2C7M+BKZibsEZwhxEx1OXXVeqsNZ9oYQklECWXbfZNfK2uz6VzDGOOoD9y
JVnrtQJsh15gFpUT5DCeoy5jRMAqSw80ueaYBXWwDe9d1OBPDpJpPP90msgEB5zz
Hl0tFck75xMy5DOYn3AmhPz1ATYI2gQAPZ5CuLosMKQZQVcHbQU80NDw2x+nQNje
HLXV5xC09bZ+rF/sxeGWy1ICPEflr11AZMhjfh0XIB5Q6UzsntrTZL1RfRFo6Bcb
6Y4m9BrD6sCAtPdlUdSAjbhZNXxPlqIVUpHRzPAYstI1Rs/7krAz+6j1wSUD5BzS
ste5S5WvAbWltE9jxFpejCkFoAMBy1EFau4aU+TWTCS1ADWItU6w02k0JTV5AJ8C
mGtR0rbMid+ELX4Gh+tmqTdCLJ/OhHxYIYVsvPjDDsg5Xh/BNHfH6kxeH//Fo68W
NbUWy0xEqhCXf9tZoVH9OMC52Z2Fz0q7h6gOaU2D79xzKVvQA7M8dRZFWYzJzu5V
hcNc0/kVF2ryE28jnVrgu3gq02JDTYwapSy6ZKgMmWf8fqEJj3Ns5StiAJHfCpa6
20W4XkyqpHs27xmy6ckLnbeONwjO3DCSQsOC+KVt1uNtSzmFV7ouAN1CLRHbHdvj
6BSUDvfGHHeioMIGpuCFXvok87ztMlKAZD7liuvgjCeGg0osfYxuFPO7RXSJ0dZ2
jqTGQpaRrVdz4MlM9H7RXo9fBRyMAGuEkmNwFPeI+ufgW9NsZE8rQb3Wq3tRCwkU
BCm0Boz65+bFLaFU14ITo+wz+p3NPmMR6GWalUtyZYapgGhuGIshhhGEnK4mhdeP
xNbNouJWfPrW6ve4mJozpAPdiCV9VEhumcitN+zcQ/Tj+Y1Kr3m+h8QK11EguJXq
0m1zcNof8Ko4I/lYg0sy4+wm+gVhkLW3H6RP/kWQCRIRi8JJLivHiv5edFGrjnuv
MpusHOUf2xJs8zTI6DaqFgqwwOUqo60/HEMq69iMbkr2iPp5bQWsfqVZs3AWRGV0
r7VBV58Y9ECSe4CVof4t3jYf7FL/lTLywrN/OyzzRh+oLH25ZNCR3JEImEHgjZyR
k2gB0wr/zyzMbM4yWngItF6TYyPCmkIexDuv1v2BlPaHZIMgH4iJxkTWjAyu4hO2
2rU0IllGXRPEz3FKCyyXGp0cxVmCBJabmIPd8/nvEQBS3H9zQKUynVSknDIO3wOV
LmzWC37zjHvRUJuUfLK4tL4EfWibwSYPFCncWgC67ALFapVi2y02y0u6l4oItWRz
2JSMimLTtFYuOihkWce4rT1i2ivKdx2rIDslVo+KoqOIMQ3Ek/sYR82Dd2fmj0u8
o7kXzJm/m/sL7fXquLXlwHHxZnZjXxDPy0+yg+xUCDH+wzbSTTu/IjVVTb5AL1Kr
Wju9UToWAvUPOPaWVIG+WINZTwiVpA4ADBi8L84z00LFSwpd+LLkwS38rCuiRQxD
iTDyYQ8g0Hk+p9f/vJpslKlEAuG3gZHAPmZsMZk08x9xYzk+DpwVyjT+siYjmiJ4
0jTdlDD0e2z3+MSZx+c2y+ZHzOSM0uF0ilANXxZw3gnjzZfLdTJTmKruHCLGS2uM
RKXlTcaW2EYTBzpzC5d8/iNdP6gFAmo8EKCgtwnaec0g5nKBknDEiBVr9rnW0Lac
Gm0qIEGf6/wcM7QcTDN34KQtNv3S/Dv8jLghiKKzvksGWB79Eh4Zm+5bNENc2XZ+
LiRYzWEI5cdzp5J3/oeOfSJwboofo5GS6hvRp+0mlHSacfnmIMwOI6Hcr9iCVUyC
J0l5x/Z0mccR66OkFAR7VWuvf2gkcbzoezhMlA7OZ5QUo+0d1tvlGrAHNr5HivyK
0GiV7MKxUcv2T65f/LaXSuvdBLkrelDiTuSKgL8OWbOx+r4XFUFgt4qQzKDRTHn0
MLPz7uGdwALK+YwRVEyTiyEzOlULkKp43mpkRQzCYZRxah/9ckHcl4TPHK/8U6W2
ZwT7wnC3ntwOkKUWHdZmju1hxF186IDXS4ooVQZvdQPCljwXPoacvVmmQlZcc8yv
CpUPX2YaDdnEDglnPECd2ikIimPwZHomxlMq4uOc89AqICYKH2HoZ3Cs0/jtBoNA
yVnGmfnv/sC2QA/xgG56Ve6qVJ/Mznw2CM8KHJSQVV/qjNFiY1dPX/V9vLwLuWoz
6F5R/kBP380UNRnkTpLE+zpR+uJ+lxhWDeFiWRyn76GKfRmun0eIxUYr7j6xrwHD
wdaCeyk0AcOr0dwOijn1xfg4KKm76G8iee/2Xp8pfGhF5TawfMi5LALoLL4qqo2k
hET0AMfCUj18sPIo+CxgoV3KhigpLai4QdPpxlF9wj53O7dvVaSQPGilL7Um5AkH
eU125LgQ3ED2tc1T629vNgM4cfLmD4u+4iq4KPr/bCR1blpLamdLLjewsSvJnUKJ
ZG0Yqczed3kJc1Wj04Ik581YXsNNJ1/HfusgsCKjwBRKxLgnLoRG+FePH/FXM4GB
73tyIItqN1kl97i6fr2cimeW/79gxOBIGJLFZsuaazYRUVvCvPmzm9md4UpWdrEv
pjjedT1RaIcHF7xQPbrd1lnmLPDvRX1kyD2Bd8Cb3ZjJCe9u/v5YawgX5C6Chq7i
yqhtxBV3e5rAvwn/ioRgbBBdYtjTQ1YY6CieMGVWqZwuEqupY4LeFKJtGb3oQIO4
algtu3QLUug8n6XPVBWE6Dxrp3CwDlQc7Xk9ZoLvMctITlnEuysfbna+pl3zjLwa
25FXVD6fZnMEM2MehxjUlaG68y1Pv11F02cS8GIoefn7q48o5Abfmm3xJOoXjxri
MAGftJ8/hL4ZiAs4/4HyzDKr46G507xPR1A76Cly8e5Z1OOdc6yO3jI7lSX/mCL2
UF3O2K12+dTQroNBZlEbRzD1mlhJqRmvh6Q+i0Hlz4FmmcqgVrVLdn1nsmSe/YlD
iDyIAaFDKg355JlOvPx3OnfBtNxG23uMe/MgJV9ujcb8E8Gjki+7av6RarvTa7B2
K68NB+PR7lEQxeljzBU5LBOCtw2a5vXce54MHhfKR3KsIOqU7nwi5GaPzeh6+gPt
aG+PtZomTYd3PthDmYAMPfqBicquGOYJEEwn8IGOnt8Fd24xEReW7SqWAlWGt0FF
uRW5b0aaBAp+lE0R3GqoR0wyIKkFK9pWQ78O3Qe0wMM55Fmi97Yzw0H8j9qzR38a
/ghgpwmuZ1ecHgC2CXejMpzkoTzwAjxVNDP1EDwHiS2vlf6O4EQNtS8qI79jDxVE
9CXKfaDCoT2oALSkqN6j/0xGMXaoAFb+kXGZH6KF229w92mFSOKpRuDGGiyTWhwS
JlT+6acNr6sjVF8AY0Za2pf1VZS3+bHCP9aCf9YpUNWt2IBlIWrhBjQ8OO9mGfKJ
0nGfxRQIBi0oDei0WVLeYeIUcslOomKRAx0PvIWgv8boE5WK6k3RIHy63/LQ/y7b
fWl6084Oxqlupo95D+gFUQ8o+7IrAxpfvxWRZzzebvhju2rbi/Bt04aIBGpYjyGV
p9fdYIJg1AO5k07Gte/Mhr895doyl+F27mgtbei1kVR0dHVjWsU9W1spH35CToUh
TLXcwEy4N3zFEE0CD5tnHyvuKwdmhuGfY7tbjK7DnWIprCIH/5zoSaYfS8Cebxs0
mWCEIIj1SOkva13RyWRBqVR367hsQEVLz8J32gTgPDXXO1Mp17za9J3EHgCRqE4V
bT769T9u8XfQL9LsB/VEsmD7WbmK/eMSlKVedGvnUruzahzdaA6b+N38VWaVPPJJ
wLjo1GMyNRz3dbxcfe5opullcUdr84MQ9gGi4s8FBtobsVKwD3RHRO0eMUlTReWo
NT/6X0WaKlJMufLKGXjmtZBt2Ki33oTutIGt0CwuRTDYnFNPdQ8QmPl750xwVedC
7enfFmpiFhVCpMLyVhpPVcEbWkStzqsHB9iPX32ivlmKrSnmqPamf4N5j24lT67I
GG0nbYXoNyYmNzolFhh1NcM/trOsJnvUoZHVKzSctVZ4W2dg0kK9A9LfLDrSf/K5
QSs/ba7P942Z32q16qYFDnP48ItOuEfzQn0kUWLZRq9uRuDJGz5ZsPNo9Y3itPfI
voCatJfoiWpFuIq1cx5RHWYXjsYqTxDRsJGOih1RlzOp5KAOsD/MK89O7CzZ6QzF
vZ7bD/PqosqFZk/0t5UbEkXt5ViUmebUzQpN1MndwVqzkWJCSU5/bm87nj5nxqe9
vg07GFWHgHa/pHMQD1LSTB3ZGGflfdtl3Km7bKBnP/9cxRn1Qii25ag7Ik/KaVdv
2XsSXOUHYEbe/oNEbeMjLzp/nXto8JNz7NzysYc8yFAvyKVHkgN6vgPw227O7UqO
Ef4roZAzWt4JmUwLDh2syADGYGjjGJQwUF+2h7ASbRkAkdpwc/znsse9bG53MuNf
6/tYBzu66UfOvwFIGTcBv4WsmcPogM7AdzGnhw4V1rYsbzyxoI3+GPBBhVf/+eM6
Eq9aojw0/ty2fpA1HbvdWxYl+vEqG31bBZvIDWmVsbpXXT1E0c7U9LCz6V7xPpCJ
z1Zk1O7wDk6GWZBjoGuBdShWGL8ljVOKKBYE7KVe2IC8qXeWOgJUswdnB7s8Z1hD
a7OW6P5BjvS6BmKUkUJsg0V3SES/ZxUCwOH96iflNBfafoq9eiX2cn2BHbLtALQV
K6/b0+pCTo7I12+pUgifVqVMIOJouAvWtDbidswD9YAQ+u6z9rTIqtSDO655T1+m
fKERbBtNeaF8NvQ1viGlj3pKizQL46JdrIYsGS5IwW1NizQb4NITdpn2xZOoLPCo
Mc8k/jTOufSCB6p/XPAvG6Dz11CucM5WuYwst8Srg0KRPPhD2fnU6bwd7I0zPhdY
AY3OgJj1WNyFnkoY7SNg2z+AUYBkG+sLBIiPLM0d3S/aPS3/kgIBa2HmDXC241r8
X/Yt17A58a8SwZbo9NB9YcfYHlkqBzQqxLLJaWBh4aZ/RjJfnm1rxq5XVem5rJeC
KK8P5847wRtx+P366nZvhRtiU0UHMRQTCT7yUd74GJI2+NkWfHSuzCY0oYv0YEzw
a/Kuct6+NLHD8x3FSsFp5jUxOTCfROBubg8u4BW3dk+cADTkbSOexKlRCOMjQM4l
awNsSYxTIcn2J5gsnwG3G/+vPUJbQ0C7ppaKQxLLXDQd80KZgw+Ze5OqnZMI08SV
WySmpDRUC+qK1LeI7o4AJUMltHhR7vXG4qZNKlw62J7JXzFY/Ffz5aSyrsa0SHAE
XT2JwcF91wLgfmSQL+VgdNwtlQzyVHzz3vMQM1DAaj6z4hlj+C6m/Q3XL62y79ru
CuB4oYIHVn5WuIbtJWHbmgkYWmm4TAnNb0k1+qdemoOSUAg4+xFKDopiDOMHUpoj
AeIaMSQaRhzqInMVE0CalYiT8VccsVWrM1MtpTCT8tKEk4Dn6ExwEgHJXhXt84PE
jOBfsiUIFL4krkIxNEGsErtfAcFKfLYjPGmSOMkqXp5A5AALEaqohV86+8PbIUII
rQQvp4vXj9hmaCaNtcnHUQ6z/+UmcdFI6kaoVKiwWmNO2rJJ4zbJpdSgnnVyuw7F
aGkkByKutLdWvqaKrSavNH2uOn8F3nlD7EGfWMnGshjdTIFfKDtvLpoYFwV93FY0
yZIk3BE3IUXubTnbSWeT1Y55gaHyGNq9qnFbkNDNKmDbL1tmx/R8L5SvrsooQqBX
lDtPttIQ05qt9brWZSm8SNKSISMOmoz03IXd4cFDKDmOvX/kc2pKIu6yyo7AJVFV
Sce4PcZAQUTwSHtBRzrZCklZklXeMAgKsvzoLhhQoIQbc5WPLWVGOngZLa4x1q/c
DhYKl4StsZEu7VrHE8sGKccXBc0td6H2mrdNEHfWthkeia26MCjIM/djCeKRKEJp
7Y4I6YuAzSCjnFxptqvTEYTAHtkOgzr7tfvnpinne3SCJkJhPAB87j9DXp4/clbS
gXPeQ3zalO+UZ6g0ohYj9WdRaDwVDIPTb6PE73udl1GkGBjJtDNHCHndah9cNl0q
eYqBKtfgwhV4sddPHB0/IAGKG+bOifzBXiAG7wrmEwZfKUJPulD0kqgAPFoM3MK5
rV1+Y23AccKFLBGsPdx75WQVr0Ah0ReuWIvB/YS2Lq1+o5u/b/SZaZhSbeH1p3yg
9exx4PkoJ/WYveZEv8DHcqZDGQyypLLJBeYaLGN0E8mxCOSaIzK5F2NWZZm6X2+m
pF/utAAJYfQs+Loj0eAvJsfIiIoeYBwihe8ZnsQ7l8nnB4L14OvfSIQiSL2EK5IP
7U6F7WnkHS79qe66qhhkXRVyIsmtXgk7h1WLNGdCB30RGmbRDju8AhCRZsai4Wif
HnsS7Q44lW3Tfi3E4N7LHNOdl3JTgtTvT9qJ5bWBB88iwiASauycuamKhGvFQSEA
TMjY9aC3c/KQD8bjdv6HpFKIfeyDSihUKx6SbrDwmaJDXcPg/bCBX4s8NjKPcvPY
MGxSKtjgzm5pZ2FPE/XdoqknA+phY2fB8UuosdsEHOGq4lUrbnOIvrG/Sy13GQJm
+0hViAS77152wazHo+yZ/KE5ZZ4onk/c9thzjoyJek4xZJDVoYbXHpyGRz3iMwCv
SZdWmPUHiLvru8DdmH6+7zKypH4/cCyOSxdLGrl9AT3EhmSf2pUsSxgel9WPX45n
j21Vtgu9Kse4gK2nfbYVgUyB87SBfprKnWV0t+37mKkKBZpQbkGygkoMu1vF0Qeq
W8/Tz6961ppzDJndJ/+YT7yxOHr8bZzitOMGms5ReKv+1Eo25SQT8eehHOAWmFog
KYbWby8QmXxQt+t9Ml9hpDbjrnhoOCTHutP319gAYLOcYwBlJrIXWktLh6cdtutg
AHRVqFZsnNmyXTNBSHPxvjEu/faBnP/I+hokl+8uShhyOns2jGyMGeFWtBvIf+Yv
awrG5bYyFNRRTMdSUMH53CIpX6Hh+2jrtsc4bE/xAb3A8p4HSqztM3799vgD2cuu
ULJCZ+YudD0uQ+Jtfboc4xgYZt39TFfZoguFCIFs8VimkEqXi3efq1bIxhJLB2wO
YAJtB64XRvJCSFuSwCV27cBCAmt9rorPfZwa/L1q2scxx5675ij+JUlP57ektPUS
9z6KcZ1cA6tqD63VIiPU8sP4HikOcpSwm1MFwsxdj8cLwFi9cjAONuO/wf1HHmqQ
xjLmI8JoxamhiOIDEGsp0Dj7BFgmIbGRbQOQv+LXgFuxNFaeRPWITItsQbdAfD4s
5jAf8fRDJzidM31KzJO/cwtARzn4pjn2GqtOWfqZAV4+7GC8jRhDDig/VCSXQMbr
dKKK3Zde9Y8zm0pg0xFrq+wFHf67YLPAPbiu2gCy0leaNFqw8jU0pQqSVR+mklmS
5GULEioJHl58W6vQyM/y6CVsQ0HmV5FqDJidMOBWtfg1+5qP5XZWh2SJIqcKhax1
3zIQZhkc7wVJljJi0TnlSuoRaSbj6/L9DLfFYjbWWx8JAGAuUP/B7ZNj+FJW7lrS
fyGTaBgumCjujqyQcEHeEDHsquNwosFBmPQAsDyOgqHKCqFy8qPTr25rexZB/N83
zvhz6IinThwZ3k0Wo/M94P1ouPfIs54pZREHuDyqCZgGv9rZHqLGqk6aTEYv3q1t
d2qi7IL7gL341ddVihxWBlS/VzS85Ojfq2jiaV+UyvXKlkqyEvI9eN9qS0kITWLL
wm/P9bcPxZwDv/oEzhuBiOwlFHiD4DG6cOjjGrxxDKFjAygkj5G9HNsmEU8pGpBU
bdPGk4HZbMv26EqiZ4Btu7QB2u8ijsb2tm5Ezia04eukc1mTeceG4xHFXOVrSmR7
RsqdqZSUAnT900KP4LR6r4Z6uMyE0nV0tEEMvN0bUVnfDF3zXLSQa9uuvE5WXOSt
uVhQjfdmDdMS2nUVu99gPoawHyik5tZM+ja+ipIKE1vXG15vu/1yHE/PkWaNwGO0
GVKgEdpndoWBF2z4Abd5svm+J2dV2DA66FQUMMkZVPeBSPbyQUXETjLsHVKg3g7d
N4NHXy2Cj+Qodh3qH1Dh0qSBYCRRnMuyLIEbW+EKm0/a0mFFsuz9xGZ0VkY04Hqq
Cr5jMWRnu9Q38HA3FpXd+/VMopyHpunuIv+v3nt+24XNo4ZgwwxEKATH2Kp5jXMl
yBPkU/yvYQhcmWbyZ3QJynolf9IrNtyoMyr7Ee+2mBvHykb2bD/ZAnpECCCOguO1
BkvxFMikWIg9VeKZBujx+8LWPfnSXtIyk5QR5eoeyYhpxp3pWRBp/337njiEwH81
W/rPLxTkIQYQbQEV4grHd0EcYc0ue6PH+iL5fuANP9t6Nk9lwwdJI6qilO9o8OBc
IT8300C5R5t+azzcHAPZbKnXoPrcoxpmlwvTUnp52vV+pwJ5Ox6mSWaqr5BGhppS
b9rtl3EoH92xllpoGfqM7Ry+x6H6gfheL+F5kBzYchGE290VzHTpDhlPwUthRNQG
89zOlFkcJ955fDw0c+Jdwgzwj6RRyeFT0NAgemY6dMrjLfQiDZKv3C73DLAdwjFS
Fi0eoPDRyZEAcGpuJ9zG91+nckJ2jxm6nGmDqwT/gtGt7V1x3u3CovPZ2ESnUo37
L0sg0x6GXrBs3ud/YLEp1LWilMZIgx1kkt1Z2RNEDUkK70cQas8XgClkjYVYhLeX
3eaXBfdHRFxTjJqPxeB/5gCRGmqOK6ekKgCZxIUu1XdlN5JOEKA1WU/GaxSqFWEP
9yq3Ah0flO4aPBfL1Q/ToxoBDm7LoZ/SfJw5W8CuRQNahHXykFrM0RrZD2fj9Sio
4idRnI1JaDpvptP6FF+O71ruxk0LtnY3QAkN0yC7Xbr6KCY2jLXOeOvoqkC/JN49
6y3g3RUm8KF+BZ6jXF/DtK9aPOfRk0LHgpnqWRqqz5hfdFdcTJkS9qa5X5UM4j9Q
NUw1XGjE6FDEkqoEIzYgHzWUdhO2R1W75UjDtTmb31px61PuLqJkzfmwXlr39vts
k8+ButSbsU9/Zv16prgp0iuAz5TTYVq3ou29jAMpjqCjDjbFPP/vpu1Xlq0kXwy0
cLCEwfN1icAWvqnzd1CyqgYD9UH+UhLPQgkjWx493V3eQSMabzRquE7rYkHYy6aX
5M0BJq59EOPYPA8pGn4In8rQV0bFtYQdNfypN01GajTGxXXsVuMlR32riIpQqW31
t0dFAfyZsVlObXrgO7BSU7NEbbpYqg8OdgBoQRVhRgBGOyiAnDd8gqIpxlh+952G
f7SKrolmJZQyDhxEZjF/TFFPVgYKN4UKG57iMmKNDTo5DGtHU/FRV2CgU12bHT/h
s3S7rE2GqyM3X/XrmFP0i9/ZcM33F3FWnFKsa4HUU4XnoU7VZRfEIXgdumMjCxg8
UQ2fFx0eHU9AJtDUxWVhWC/OzD6Pgtq34zALvhvlwe6M3O6vTazf7LgRAruSpkiE
CQCD1PF0eL4nM9xh2oH25JiKGxEkcLVZCT9nW9BAANeENZWGova12XlUegbuiNti
zzSGYoiNY65UMxO7rT1j4/3IstabPkhoC0Ww9rHaQxQbaBu+g6utkjtfq877le92
oMvo7QFQvJJ01Y3K0J3SIZiMPVC0HgvsN7lL84HN/jv5IvDDQvQA8bLUjTvWv/2Z
sEVN8jg7g/U6Rwn73FRWexv/JWEay9AHun6miIS5lDp4OW5VrKhDBF61PxiddOSd
b6SkT4NkxnLpSTqdLNTptD3/hd6Lx7RsFVfd/xRRIGvHZYY5EXiUG1MKz6hNGJYX
hWGk2K0ed68ByaZmifkFXl/KUKQHuflCn9lU87quu47gGlD8QllbIsRsS1+xDsYe
FtW+tDDd2D5Z+CnHEkUvm7uXcSw4oCNKyE1jPlKqMQj4x6cerCUWy14KkrZKJys4
+nPEfxT5ZzhQOZVFV9TStkCq28MH6Zo19D/vsg1wJM/ZjahgiysrFHlBlq/ALpS9
m7FOsP+ETl1sJHE1HHATOOI8cHisWXYRFWougsFVC6Lvtue+RmG/mwbnKFU/fQAm
bdE5jnZY5b2hdjqof3xILI59ksulCqY+0HtbW1QgzfiwfFY4+T27J63/HRL57SyC
9jpBZIwBDpKxATk7FrTfA8hExo+rpJbZdZD7RApbfGCBe14kDU8T6loQUdeJSpEn
I/lJV4UAfOe9VDKcCC8KapAAT4xYRADnxgS4YNUM4oyeLTRV3h5RordCga2n9zua
hLMCQVKB7IAPH0x8fE7j67qy9MUZn4X0AGDEprIYTW2P1WPcasdKYADUCNn6j8Ye
rlqRw9WujounvQVfAD3YSDCpi9+LRSmKlWLbPUL0BO1TbgSrJ2n2DrGD6nEJtx6U
CKNFJmaC0sd0jEfyax9QZe16zuBOLE/Ol6JNWNifDypnJb/5O0VRgUoyW1GTMogM
hiHZHu62uem0agBuu9iwSqsOiOLR78hwtpB4l9QtmE0ZstF/1r1Sr9ZvmDrLgYtR
qzkzSC3y4CeXC+okCPhtLm13UzLJNV9x/xagxVbCP+fLnYQZnxDS9hLcAO2RynBd
s8k3wKqM7g3sHmHXUoeH2AzgKsECq3SzflryU6VGlA0j+t/97OlCji+TChqvpj1K
WirT2L80obojecwy//+IiWL5pkg/73TrKJ8tu6felzloTaj96fWi8tdBmCR5B7rH
KHep0LNdHrMcnys+qxd/STfP0JVTrg4L4E9QMdI8w49zpgwaV1NmMyDGEpDYagUC
zJtxBwVbeS9LXleKZ8jRoAuhAGlxwKSBblDhkOUmfQoQ7wSBM5Al7W3sHl8dzkp7
yx8WEuFzW80VtfCvGMEq+g6/zhdyXSF0i/fKLAhaTuUcdd310gbX6FwK6y8xtxxA
MZ8xaVw0Uh4nFyD8hBsDw7QZ8LIVilj6senJb3OwcAcpn8kU8TCyz1lKnGUOVO4n
RATk5wR22RlIGCbIYxrWIA103KoBuo3fOrVxnk0KTahvJ2/UXqjwaxsSZo0KZN9j
E+WPqHVVqauZEEvn69U5If5WpLKEZZTCo/y1aw0CoG32bUtZyhvsdaVWL7/JHrlX
ItNuvH0WAokV1jz9qPKn+JQlOtoVW/jMqJ2rO9NKFro++JwVGlJkQ6lShqZDw4xd
IztKlYCuCAVouhuNIjEmr0Kq1C1FRcIk+fPPP/D95lkuh3G8SkfMyJjngGKWS+om
uVfOeCLmamvJN5MT482KH7ihuuz+5+/BduYZF+AA6salWbKQIIfyfmYoNEOTMgAm
ZV2wwyvw7BxqVBxC3FBkkOoFm9+Z94KFerunomncuytxpTnhaEHHFPPvn1bfaZrj
WoU5uthfeyrHOHpcHkGQNEzZRIPcUJzGWiRzGW0ks/K38xb0Xm9s2rm0ABDPtagR
Axe2XzCp/zS3DesNeoJugN6Ih/VSZxU003sSMKCWfuTVzuYzsnn0YqglE6Yk6II+
EKCV4FtgTVktWHNIb6hiuWZIV05RoRdhtvrI4R8n8JrAbpvjuJVY18YjKkCG/Cpz
yWiMGYJohTQaAC8t5Nphxyg+Ks0l+wW/nMCx6R2U9pUe0noMcWKbKiFCdG00MM+T
CdRSGp2xemJkj9djH1XwwOIGHAtt7A5ue4N1JpQRC+sWcpMrVZQfcR//7lSaiZqs
k0spUO1/Rup+ZKlfaDR2xdIUNv38ep9XnaauOsYvn1HmCd0dUn6d3Dl53TzTaJVb
tkFB49Pel/wHERhB4oy9IJAiptZeXZVPm2MB7WocD8pVgTysJYSIrcgv9Ewap2Bd
o4rxJMW61Zehvt/EJj+heRDT96Eph1hTeQr1mn7DwW5BsHZEQDhDmpm5IhMIkKO9
Ks3FdmlkHM7N0PLJUqDZ0rrEmvwL7zD0X0bEQESfFvu8fTLMXZjRyJKOh5RAL+QJ
XF89HFZ5N78b71eVYxcdg6fv1wEAoheQzsZqiFSRc/g6hDgBMT/DdiivJI8YP7xv
/AA/VuZ5hq/FPPuWkfroklydWVBCT3hkk1sfwFecpn+0zcx3MIpHfuELc947kDmb
J0fawkOlPSdfk4dwrhJIIRxTgz7jgBIlOAtxYM6pMO7dKlz0D8zCHW+8FqDhjdag
CZhqFDc6JVd2LLMwu6/QBIA+6V3NB4fRPKCry/WJW2bSdAC2vc0DOTF9up3N+10S
qrn+qob5iViNKtTYPhLQzE7alPwRc2+4YLK+EKqVpLGNZeM7NRQqDG192aXHmhjR
XHULURot91sLxhzwVw0/4N/J1D7/IU/bto2vxweJrntcw7dxHgcZwc9aAIkFUyMH
2dyKrMvYZQ1CP5VWff0tZsWU0BelZSd9h/4NF8X6jiZ3n5Jde0dot2lidZj8wEBq
eX9ImrWQgozSF6rQyzsPWkiX03y1r9Z5bTmxb5Cvdv4VcscwczyNUJB+zuVaZcnw
5UwaRbYvcC/IeSwrux5W79yRLqKYX1U8tEhZ1gON99Htt9ETD8A8hwBRfeHf70OQ
Es0wrnTdGa9JNTNHaGarrwwfQlMDPIYOQhehomnrEmiAJc2ZvVW2qEWxaXPhQX9Q
Dz+k9yxAQ596DDp/ixMAQQCfI4o/Zv5y39UNJPKFCVXdG4/Z674E++JGTAWuubjY
2HlKY/ajDHOHewlSOCZbxm3erGYcTyMDKTYOxd5U9Z3BSsGEFk5YSJb78OSJOWCm
ER8Ta0c2jgH1xRVcGNNdzU8q3Sx//Ewt76TbeFX5WqsikqwaGTsXYTzznqziKkF7
8Dui0Q3VC3STwMRgE6aezpFti7qQDJMvd6dJnrrzqOX6QhM9HnKFkIZCoQ9WAYhG
iMSOHJ+nJFrjgRCoChblQpxo3QD8j0A2LTxIxUC0/Lg0gWFBhwXiV6g5f3kepjdv
6oPuF+oEVe5bT58cU3k8PgdONLebXzr59V7ARgeMz3fg/VmYl69FH7JZCqNMPVMR
rRgww1t6A1OzQGCdNQWh9WHC1AN4NApTnRHHekiEjuwPcBH4FbjQqjLrXSO7F86L
6ctueQTHVvI/HVZp4Z9/6Th6s+xqdeqybZDzZ2XrPZuofl+6rMh/2DoHHTJEvNVk
fIHMJ3ELaIvpQjQHu6HZEo+jPeqdCfVrLYzcQgsSVnwDBDCxcKo2o3xEUaI3HhMf
SY8TLI6qvB8NLkS13O9W93QLB3MZFbkzNL2jSzZtVsnjxPgO/XzoUjMuJLjpNSH7
WsHnK9tldHkQb3TOS4jJDyPBoszZbd9wXPddUxRHOdRYXWBrC685/lY5jS71YRGg
1JhWWI1eO3uB033Cbpy49Y4+f7Yq9sw1ehzsFkdEXHwyhV28C9yPk7B5vrSq43Nq
O959UuF9hFwG25KCz08DlXWlDaK7ExV/kch4lsdi+hdqSKHVNk9uJ+29kvWVWS46
MxI2j5qCnpc8IhoUUNbz/YwyElpMmHcgsoSuQxzSMXwTScHOsGKvbEy4e0KI6VXQ
Pgafmj9b65WuprO62Z9E3A3btOx1OLnWswen9pNvf7vdvY6R6U8hujUFSYCBWfZZ
NK8ukJFUfz4Jifnrg1tmyGQTYn62ZyVv9xaXEvUSGdzqLlrXRm45bgRbudUQK2aa
mq5encnNiuZ3aVArUgQWyqZY+Z2PktqPLCZ926ck7wblABIPiMmoj+j0OgAVeZ0g
y9l/2gQUBRFQWN8UEslLYkxCMm/5sraHh/7ja3CYVLs+rp7AuaEgJnVhJHnXgKwA
bOVecqsHKQXIpLSziVeCDkHqAEVzwXWjux9Z//SHFxjcomNcrUef8KkUqT2d/Z7e
qhnatlLzhf5sckaF9uy2CbmuxzTSB8wjxs8drRjvUlYOnh9ZvB4BOiERMp0Hdzd3
PQfj0hIAaNgCsHJoDCjOTBW+qXdGg8ThGQTP8Qkcvyd/MDijYq/xhWGOj1L6ukOM
IgMxX1ZkAbUIRwj2AALp2j21CaD6j0YK2Nu5zbHb1b0lcA4sVC1kegTVnbZ+NtK+
l7TuuW29JpvOil1lBEzq/rj5mcn4BaZF3hk+zmiD8V93ALjuet8qJ3WKENHK/3G+
5eHsK0svxVspzcPUL48IVrJ71y4mF6d0mK0nz7FpuU5jy4C+SZ9G3Gnq5qWREw8L
qQpBtacvNrfKrv3Hm9fagckLyMtDhvFuVt/5ifie7SBzpjootsN+A5DyaYK0cuPW
9jGhGK3sY+V2j4RwW3nVZvq5HPhhxurZG3K675YdOFQ1mUt0lL+wXR31xOFzbh9H
QcTLS7869MmAevM2yCUSgGuIZjKwIFCa+Z2VwxN7OtoKZdVWV/cW7zmIAsJ8TXSq
8tXCtLKwX5fRfLnWyCtgSBqvR869Vs1h/uU0I7cxeYwTshuq+gQGcr8h/DaeT6yK
Un2tj1dhiXK0eHcAyp4SoZmy50UdlzGDkJ0jhprEi1B+6G1+/LRNB3cDBOZYad95
ANvSYTxFQa2vqSUKBdT75lUizdU2IjokHb5YqOgMWu+SKA8WYkRJLdSbAKHyas9a
xgD3pdfX6T8TXUb9tQhMhZofIrofjZGqljNv9N5hTpantr0dvK5Qnbc268AU67xO
7i37Ft+wlvIZin3g9kLE/3YjNq1ONs8wMmvWid17+hNG/4vevC7cIHwIONd7XPB1
vaWcS7OCRxh1f0B1wy/A9Ia9fZNg7qSVgON7Hwtw0Gw68mvvsXpYz4EfXqaMKCoG
XTrkmmEjC7RG3Fss45FVhBfJmUmvpj+XDcn1JCv+E8nidZQ00IilSHeF+l1ZkxRV
X+E+ZFVZoND1CvYikSwVRICDqf/+t87+Thg1oXQkJZw3nJkg4d7gAkA5juKbxs12
HSJMDUkCP2mMPtXNzNIf+A/mcDNAKOaqKhPXqPemoXOBBuejjZqijc2RIeH4WVre
ANuzMK0Z746ACVPpP6w5//WK0yvv+NbRtM5Z+F+Ysp3rzbkh6iNoc4CarSVY/0rw
3wRmO0iUPSBY07msgzfAbC7iUBP3nQl8pJx7OHjmw3f/cirj2DrWldIsqCXP9Ruo
zMdnIry0mQn0yPhKYZFASYl46SBujZN3rhQYRMoHJ0WUo50xfDMkFaZkvmCO1ME0
uduRDMNYnFvelAPLo1qJntiZMFh627kBaHdXPiqDatujRnMaWOrStrazitszPEhC
IHR7NIZD6H0QOMXvzBa7bOVIWsa60TH5VbvCCKmt89a6C7ntoCLSy8tMaR46PVfG
fsLxJ6b9Awz2FWKoOXJOZptKang3SzKke8AaVoWQCvCk9FX4mh3hyu8KTP+U9YRK
kJGiT027GbwoHEZzTNvVKYShhpfvWiw6W5xAonAL/yBK/AKGS2+ZoWKtcAlCGhUE
QFuXZ3BbIWRQVnbLmpXtgjJlEa1vuX5NJHDqQ07wVRX5QCwpkuiKtkao5WdVWg2z
WdP6Cd2mO5NsxBVjNGcjqIdY1WszLAYlFN3xSGH+e82qzyeHMHvIXlyl2jUPeMxG
/c/nu4oaLEUtWPN5r9rZJG3mvtTPNi7Iy9BMZ1MGC9m0+q0AZUxCbW4thtHJj8JJ
iA26RPA+itGAhHonY8JBIFwoayRWiytL3E/PQGEXOqSkSMV/DyRO+qPl/CetEZ4Z
lFQc6frU6iEqfDWEmNAzNfKpGZcRjLjPLw6mKUZ+A+9aeJmrjcIxkPCa2ETOY7PA
6U2xEA6OPiPQI50G5XrwyfzaYUwOypuEodJ/A3S6hTtyYntYSv8/BdIOvmILRy6M
tH3TEZ6LyQHwlSaTqzjzckhCLkHM7wd8LoY0fy2rj+ZsxG+WI26SNoIxkTurX3J6
BZtPa5lKfDrwrJdYyTTlLY4FFD5biayLNNgXQLjV0f7nyFDIy8b4oEvkgHGV5Rp9
6e8qHtk9apXT9pnKAsN3Dtf+QKMFDyaQUz65mVZiexPq7dtNTUTo04gyANWZpPmg
z/zzcvwBUJHX6NtDK3skBVJklaGRUw7nBvY16GGPSf4Gc/z1P+JtAC9od2xxnW5c
n/zPBpotFQG3LccnnQEiL7OOHdeUskerQNVr8jBURHBIxlGNL0qLx+SgDkwuTbe0
gYTN6IeZWcAimfrtYHMebDny/KTL/UJB0+xpl/DNmiohiYVxb6sjha2oYRT+7o74
cxqOLGDqKRf/n4BCi5TooGr4YEghCBjkzVCdrU+pcWtV7wg7WQJmafh+MuQHtHKs
i0dxsDSd3yz2BVCaxdAShoUms8/SucAt5WdQX0GQq4OcW0YL2dDzWrz+OasWI48X
Ijd+rQxdJ/kAynbW9JO8rbcTxM1BW3eFinvY3z0WfxThgEPX7aLQyBiPIBVVswXV
nsOpG8aVsv0NmtAHdLbRXjYJq5qsmozMdmUkHMrQ28d6Qfou7Sa04UjwUmRG7DFh
ma7nkoBqwNiRe4tinEh7rlfUCJxkRb3Px5Wc5nD8NIMhbmGqDwTrdFL1jsis/rRW
2kYnz8ZU+527L8pk/XzDlAO67hrid6eAZMuB3bhBR0t1BmZIxygaQcrRdff0JbnX
Uom89guoDHiN4JRCy2mTA8fmI2xRZtHmhSUc3WOpf5jLYlosaewanRIs7spG10YC
Y8wxUiJ7CdXBjjtoqyd7RsLptF9VMbsFXopOhwBKcjiKIOVUasjKv23QB8XUvL36
37nD0xoyBRLt90Ar+cw35I3w6QIfSEc4plIufdtpQDAdktURHzoaxHAUPLmtsZMK
uIL5PpAZVvhJQDF31yU3vOQUEaL3qACUgSo3UnZ6lb9iRLQB6rShfWc3QqClY9H6
Bxm/Jp4syEC7lkyVD3IlPxc0kinLV0V5jcs9dpGClTxQuuUaiYjqzacaFYEXaROr
qv9FUQjkch0kzfEEDNyKlQKTtgLX/szZy8Sk1v+0WxXPp/khJEbiWckofHjJNblm
aSVqAu0QwqPwvquIjDoE2OyA2cxsWVMB4d7tZyiPgsOJsTiX2Hc53+LBdxX2mipz
f9elGgKL2dys786Zgry7IGG4yhQzrB4QT60LbN0V+qnVGj3aM7Uq260add1l1V09
uCMyNQfQIwVXcEvbt348YPrKtbiQYB+BmOuujC+DFE/olmNdWVWXijBep/fQuBSh
4x41p/B27tZqPcnUz9Um6XsiOEZkjcH/ve/mcU6dWrIbwFRlCmLD9aWw6EJPcZaw
HokUjn8IeJ+CseHStGxsnu3QbuF5SUxtubbqfwF31XfmEkMc7RUCub9FxEk1wEgd
3mkch7OjSAqnjW81HznYd/88DXSuRw6/8SwtCeCddZTua+Uhyh0YOOBsbFu3jJCQ
rzwTyywvH3HcQJ/3eLT+eTGNsVqoLCcqrb931RSdp9OXSZ6MQSndIMgW7XvXRFZS
mrniGpVuN3QkQUw/n9oRfNgT28R4mmoH6QtnKr1GE2tQ/LLxoPcavEnnUo74DLTs
TNafVMx1eRiJnphw0OWiaiuxCFanz7LblV6atFpqFchTrajl5Q961Pq3CDuEe/uQ
ep3cznRGug9AJKJHwgWJ/c5wEFoRwwKoO3NE6PMDYWd0owKZyH2fp+K+V2+FzElw
eajfGQTM4L9NoKRYykVhFsLVCUd1uyMhnlc6dewV5V8N8NxWPlLKpPZmlS8pLf3V
q1kMpYUN+BtsFY3t3J+SW/bB1qIwAmNYnUOpolXgV6PD6yJzI7GaCzllKzXNSdvL
avTEy6PFY3x/9mKBwcwySgiCdFiz+WC3+4VPLUGwGxuL13/w7rX+qBrqLd1PdigG
jMjY4VkQUUuZ+G8LTX9byaemRdB2jg1ZODEaDRcHOqfw4Oti+uxBKNDcgA8IdGrr
wWrngtEMAOoUdokn3fkjLCfB39OAgUzaIv4F/MjisQIELJkHf8wqCuLgfqItP9rs
zzJPImE17Mpp9RE7Xbv2vlLvdJa4T5uP4Mv+g8jIzKBSfWs6ffK5RaQy3osqywQh
EsjySmxDhrp/mmgZueeVWdTRW2UyfjlZvkYhEf48o9fZQjsr+14nljuto+98InxT
EOTrQNlAqrHVr1jZ8LaNqFnwxpHTPgZ82UGB/yosptD05GJ7mQwQgkxFdsqYyjBi
/PgGUpFZXY8suDRVnxG37Ygg7UtqaHqELLHJJC+fQSPYu9JJ2HzMblVhhfTQvHlh
U2YHh5LYPk4f3UwiMSbYkEEEXxKK9J1eSge8WgNaBigLQYsZAU29MMyl+VWJDlzp
LSbyfjBUCBEwpQRoux+2fsT6sCaGKwLxguWQr/aswNGt1Grwo2Qr33XJks+G6yMt
CKxdkvL0QmXVq9WddQAUNCNN0eCnjZMJ8vFI8rT7QmKJ6xqaowY1aPToh6Tqa/Pe
HHCJZtcXnuFHFCYgprtip5l9w8OVM7Z373NYI8/I8w6tAMTwxbL6COeHGvA4C/8E
/Su/BPmVGnTUf8XkpV5VE0pi2F0nM5yuFflHVqU3ICHGq3EftscresXm68LYlNxq
EWyVFcwZG3oZ5yeBsnryxWuXPpYeoO75e3wZzNkkBHD7SFfLYeOt+24DzFF0Ver6
3ydDwzd1nggFm2at8T07QHApOhNGn3mlA8V4yui3Y7ptWRQe8eTvwXuwNmqZ7kUe
yD+Bjj7WbgfoNN+CQqImxZDQAByID2iOEoX1DszYJsO3xNMEZGs8FsTTHVqZoPCA
jUZsd+jOyhBumkFemPSoJSnV6hDR8SlmyRB51IEOr25Qx2VjK5OOkIfxehCPUrkp
TI9eE0bePn0pJ9yl6RGxKR9OcAKW5ExNRw0ciSOs9mGYUENTKbhLcX7GSF321RRF
6DXMJ5MLxhztaHJuWDbctFAUn0O1JHBnNrHM6TjKlvEIKauFDBn0JUT03xaxberJ
3B1n6h62NUi9u2ChLbK0lpO4YAVUzLolsc20m3LBtclrlLYzvL6mOXR94wVL94uL
+mvQ7oyxMImrym5XOV1U5PMmmPok1MaKAZ4DoZwhPkdlBJYSz4MRIELaWQ/5fkYa
9fdK4BPDj/p/veUlefwpN5ES0SyL5Syx6rEe1Uw2HY+JyQMU632ehwvStIHqCtd0
6n1pJoa/+hWUiRVPOe4DF+dFzmcZTvkZr4+S0AwdMZWkzf/kwZCFM+DusZbR+P8m
xtlL3gcwVgMcQBYPStP44/E3ljnH1ewtj9XCg1KI5bh2w4ZFcfkzjy9XFnzxFJWD
QsJqPXGPtUmlmnK1djht09vkddlpltApFWwRytzFbhVHGWi+pmLz4lO9cEzhY4+N
syivJjfSor81L83ilVZKHpKp9egGjRv79OrsJSADBuNA5m2Q9e8YIrINPHKvevsr
w8YfP4M94DCHnYHBBRfN2F/gXUEYJ6jZFShzGRD6UEmGKL1L3ZZicoAAmypmSkxq
e2kRz1ye6RTzSw18isDjD3qhuyyLn6Oyk56AnfFxm4k68cV5FXhE5c2h+W9s2UYo
d+WNXuXSsnRO+yWmW78/ILeuf7/1KPpNXNDXwXjbJkkTtef5uEauWghkggTXNi+w
WcJd7dn7k1GGNKjb+Dp5azKg5VVfTowVSlvsgFV9skvfsyX5xWAExjyDTWIIFonT
q0SSd0OgWcO4HBmW8nlsFJe9key0HxxGpIYU1d7Hy1RpFFbsVn2HpontwIrhOGbv
hqnF4P+0lIid/T8qNsgICoSViC3rf6+lrHud7YCVNitwVDPLSM6iLFGsES7eu9vJ
fNMNfwiYIAr5mlsSPXTxk6F4DL6w/qxtI1EQ3TF8UQwfdVsBOq7d08do+3CG4jch
8IBLgiVvUS894g6vX+yOyv0HIGFtoWh8uLZwtXmhTCb9+JD0Aa4SsHcVfyycY0dC
yY7oxQ/doSFyymYVrzB2PLxKrSGoU6rG6ctFj3Cxhh+Xfna7NKKH2jzYW1f11mG9
xQKlR7vBTNFtDkgHDTlZdxAjOTXHanAXmbbna2looUktS0uhQdYfPYXJCyD09CqJ
xyiECp1IE12GSpVOKIS4lfjePRmQK1VXIHV18rXGRTvS5ZIhW/laKrMb497pGCLE
hiD/cguCo4+YO2O450DycNi+sktBpL6ValuPV5eZaOASP8Ab4YJ0DpqYDvolJil1
aCpXcboK2mKDuFYUF49zevylk93VsWoSZdEh38xlF1+K7+sy28fnpgXRW8x452wv
G7GeWQ5rz65j9KlpSDS4HApiSViR755gXsI7AQq5CvckZKisttTMYSNrluOaU6Vb
SeKvlTQG9HJuBmGY6NvIHH1l/3HDWL8qjB+3A00g5+ELHeDm2wlXtj7pCnzd286A
9SYbrrs9oTAdA6XCpt8U0wlg7zoE2cogr8+Uh1eQpEKx7F5lb3B8nr3E2Odwc/Uu
ciq6KxbNfooJ23lEEHBVHRurrWFIChTkeoldai+EThwPsOvO6j4qltb+XHJvGnp9
kLgWr/ykPu3RGGfAWZTUbGp/Xu0b61h86w/UzfCn5ljBi1rwtLY+aXViAwftEouU
3QIbnCVQIH2X9k0q9Zh168t7ALvpm2HKI7N6vqdNuz2VJjjimF0U9CcOd+nETg6d
CGnsUgGHhTnvVLtVQ2OnM29nIJt/KNl6zK+JxKdOJ/C5bzBsQjtQmHVxeBnTP68T
9LO+H2qXVYv0jmkAeUXD/uJ8PKULyQl51JHTJ5gyAwn30nqLax6e66v/Z2lgm3j/
eBI9mqmVnw3jqengeJTctmm73KOjhrH+ERwVfbUzYZ6JrdMrK7iYeEY1M5lWKFB1
t1jM97w+iDEXekJp3awUuzc57iaSP6C48m+uhIf3vdFgyspFiE3rbNOe24E9qbb0
+XJ8KrSAFMZDaj5VnvYMv11+oKgbIM5ec8cKS77psnxC54fWM1AR9U2odMehp63T
U2gGcATS4oxfYAg9MfPRzYcif2tWgQLfA+GgGeVOyN5Kq+rNqG/M1COxrBWFsOhY
NY3zR+xfZGkeVkQDADQW9DHJx4ItO0uK80WZW0aXl5W2sg/yr/fWmgN5bhaP30tI
s1iSvxeA/48638wjGo8aBVm7WbdnaylP27ZVUmQUkWbAc1vXP6WiDzsGni3nXjR0
CrKVioWNYBC/y+xfOtcIX9l4xVyCvKrgtQ37dv2YnvdJUDZSh5R82gSycA59Ftnn
hEk8L5ArxSe4p8xqXldVHYtHwSGCKw9M3+8wpD4fkAZ7PA5l04f5h36W8wnjtOjl
0FZlLee3LuRVzkeR5fZJ1zGCgPpEw3FW3Zpy3J9iDksGnA9Z8TQdTgVs20C2Jq8A
j0R8TeKwZqw/mPsl+fPuf2RuiacMMNekHPOgrqdLxQpND3I5UuHFXxENtCjdNBXB
Y3z993Ugosnw1HHl9IBp8gwr29yFcqeDdc4GPyjXjWc8Pm4F+t4ZbmYELez97yqT
oWa1EgQTuxGrEaZHEiokWxSdzDFNuwu4Vx1sJJgxqp01/biwJ6F7Wgj3bHFnrpuf
pQv4Qv0dU0sY0cND815YDQ1KmVpgkj2w8eRMLR0xc9lald7bj6qGi1P9LnfEZN1n
mWqxZvQUxog9GaIoR9gj6GV/L2Ajf+izXKxEYRiofXFMbM0OLk4g3S98VSG3E/m3
0IkTU28Zqm7dWrGvmRvqTk6QCWyaJptKV0L/nP/GL7slWpUHhxM0CJnSlLiPlIsm
n02NVykVr99O+nPJIYW6gzG8OQR5dDHHgtDIPvwT8p3tBm/iNpwut9sauwjUmwH2
OoS/yqAE6/82toUaMloK1mRY1kvXSJtthjSc5dXUWpLx9sWWVnnDCaiSARzDAoZ8
/jQhYTzUGp58rT0E81BCJa40RPSyHIMyhIyoujTQItb5AgufiDEzAvaTA/QH+aZY
Pk3tGI7iAQzjWgg2Bj6Y5QBVOke1gvaltNM04kLGg0SOPfaba+BKIJ1bONzsaXj5
KjWjiPCNkN4a2jKVntW/xlOZzY3xwVM8ehjN4vauTrWHqPwjpqCbR29ljSxel5Y8
/TfQ2RVKWga2arluJsCeWngmJc45RHubvOHhNiGF+bRdkh+I3jfDaiSoqXaZkpyP
DAJLpgtt4eNbjTOLnIkzp2P0obKqLuJHIhmof1NnPekv/P70K0HRCY28u/THA2H6
1bep8/Wd3mO6INdxhofqdzdFCD58sNhfoZx+Pt9xehMZQ0k7DdB/Q6/Sjft4SmYv
Y5Pq/1DYU/R95sp7bnSl1+nwZAEgC+WvTU6OTOl04budEb9pqwm4SxGm4ZHPER18
0XV2Am/1+P2PFnv7uc8EPCd+lzIs0FFEimYWIwpEI/vs8yz+ZT/GswwzmoDJHrZ1
UKhww6SdO+U02XDyg6yPJNMnqdCnYISg9eOIpcoI2SHZCB9jhdjF764Lad7wS6nw
YZ0KztAKllnqshz9WgpFSmFztaWdoG7vU2f5lSv2nRgLPRiRlAGNwzywPEMklQac
UgftEUXe5McmmVLFebf7A/FdKneBsS9V1O6MKbeXBNOlb6fY99EFeMxyzkt2twZ2
cEP/QXm2XA2Xl647KXF8I4PpnWpa5LTUy2nQfYWEdDT733e/oCmMTgyKlktafy8z
m0He9I7uRJ7uJ9XSYIlsf6BIRo0ShABjPZDnh9QfZIesPVucHQazQU+oJZd4UlA/
gau21PqKAqr+uCWrSzM+hBkVwnY9+XW2AlU9X+FwsXfNSq2swff7GvAuzBDLrK7z
m9aTTcYbH8gvLgcxyhXLp6/j/DtAukOaNeeKQfJ4OcedeGi6dc5iQY1tE1s8tsVG
kkMMQqb0jlylwGuaomibzs3juP7jHal5QckwurvFgiauGYzEgvnTnaDlcVnQRUGw
Ko1V0H0y53N1QvSry6jc0CapqXOdTyJnBk9P54Cm7kBLrvI2gAIKwgwYinGwcVmT
zwoQMTirhjkxPPR0PJz8cuOTQuK7neVq1MSWl24qFBVYjoQe3ZWEqO4JXRG9238X
EZpGtJ1nLz8tJyIKriso3xoY08tRVo212pXYU9Ox542+t3L2272he7i9KIZ7rozw
L6+4J4KZaQss7T+nFBN/6LSUdHd8VO2wfve8MvJzUbtmNbUMXTKQ+Expu7wgLyDz
vzRRQ3CLkGYkKROJowovlF6Qw/gwEd0Swy8HpWGMs8WsZZG8VjpGYDNpeGgEsy71
UxFdqmQvTGaIz8H7sbeqOJi04hRgQttgm/EKE7RzhapmR3NDQ+t8SNUlTKjdbAZH
16FIum3WqYZSTKzwgGOblL0K1DFCzVaGFDb9ioPb0+Lg52vFkg2FvDE9y6ILVwMo
PnSMSPw0lWFGxpSSDWTRJ8qf/+nLHIEZpRrG+dD6wYyKzcD87R/xQ1xMmKcSoPSR
EPtk22H6Kjl/Ripo6PzGOC34sY4AnvZKsEW8pSO1rkqRsUBX4AkF/2+kUQQugIHf
Pr1449dn368sbBSaBjHf2Od1rg4jcS/KMEpdev9XNp9iITgf0KbRgYiGWnQNHE3p
ymynfchJLY7FH4M/FWFzGtly3YwBST2BHRnF74GyLERRGPq4vQ4e+Y/hL2WRAf84
+fSW09y5zUdM7Y0wj2WIesv4gpoFOI1FVIb6qnVbqw3zBtQscFRK+PHHmCNR4NA/
a9fmI8TCjcnaG1gSwAgMZhxlSiVF1lzu9FRvsgBuGR+/TTJZ3WSudopqemcuj2fc
lf9jZBQX8kPG6mehmkZKnlpB7iFjV+btltV7ex1MIRI1ViUfKjj+4SHt+uUKBMzh
iiqRj6Ok2hxEZrLXlGKOFOsR6Y/adfPbFB97UPezSD0oJt2jfgAYE4mXUqstZh85
dyRoiHjjhF7+HVcZOtgwwi2LSETQALRGZNwEJU/7ynLF4gRSSa7OR14PRKxO0r6I
7JWeCOXz9288R5io2b9t2/7gbU3WeOYPyDtIaiYho5G45Jjk+M7VT/JgdFCwBkrO
SRUzUbQfka5a3dJVyo89O2xjq9JHTJP1mC384vvWLX8nb1mOPSMdQBt8RRIo17x5
KkSlSmqVQ6/wjrFibpDiMnrIqtX5vigxZ/DE82XSg+5IquHFw2N+SJ/qeLegCUiL
E/cAbnGCYRhK1QdhxNGjMXE2ZM4+AOFEmI2nG+kfw4P5+MW4SHFryB3BG4CIW0BP
XK3cxnUWdTfQjZ/uFBPbGZnsB16XlbpAujC9hX1DtO+25KLCMKusGnSYQMPV4rNS
kvBLy0WngMtwIp3bnNGqlVFhset2VLlI8G9Z4WJcsLNbmOAjUIDwrA/FHRNNhiPH
JMMzdnV/dwLWxDFrd8kpwoXn5Pf9L/oCmKoh5GVaCmDpHVl8kxQBsDuow7/lAiZ4
YdxgObUoxQOw7dZvT2K+UNDBYZ+3Dj5v92ajxz0KRwnPnH5Nz/alxEVmb06r56HE
Z5t6eJVnmnAsEgnh3XTS+SXx0Kfe9y967ej0I1VD9Osft/RRYWdYk1r0mtjASKf8
qVtATf50hjNMoUc6ZykGUzILouDWjx0t95n8XIKA0kqeobTyqsq/ftxF1mI2OUmF
Kd/0HUs1ojuKt5//VPVSrc4MEWyKFFHYwb8PJ7O0lk6mibRJtCqwb8NPFT/RIAEA
OyLREUbyA9CgNFPEQ7f6VixgNAjLuSs4C47AHqN16y4EjIrqJCMcvq6Asp3Yzo7C
emT52Kud3Yl15ZzHZL13m7PRo9KQLqEyt/aHWx8O3fG1JE1c5r3zl3EH6sfnseic
0mnw7q8gZO+L2ZaxNM5SlLFqp8u6tGJgACUlYMRPIL8h8NS4ELrFPm6J+o4dF+Pz
r/Fu/yRlUrYel4rgFfB4WoERD+psZqve/rZ63JwyM31D44i2WUiCfrJBYYBn+vy+
GpUmHgb/21R1NPmTQHyV1yyeMyYfw+YozJsTS5FxQjleR2k+ZGxLo1qZsfhgZDfG
WdMOvA0TVrnZyLpWOoIWZcRF3uRjMASm8Lh9KwULg4ENBpoI/YXTFZH9W5oC4Fbw
ea2qr5wVhov0Ry+53d1JWh7KQuG6EoJCqJ1YDYOEHnQgUtb+diNtYJUGE2tbUTOs
78HfHiL6aCxukYvlDtyxrv4FqhNz7czmviB9203avDWfB7CqUl8ByV0977dB4UsK
3It9lJToqXsW99k/bndcHR6nLOfQmCZHo+oPKmTxSBBTibPaVgiAWVfF8qtDe0HF
aqsFpHmbP06sd49v8s8L1+4Me8yGR7ZaF/XcgCuuwCQJ1v+NtxvOiPbiWT1S4ui4
YsZRkTP6PmLP1woWl+3gAmjkTynMMp3vc+dgGo41poNbnQfjQNJWsOWswdr43dlO
T7jM3LT8Z1f3vWJT3EDL5lhJ0LergyVp5KF7yY43AkUBnUHWXBaMOW07iGP5jcgl
GqznoNhI1kZHJtafPP8fD0oqUlgtg65CgEX7fQkvSzvZxt5Nn2SWbkXTminKhoZO
2DdeyphpEwiFqx6Dk61tuKoS/ybM0N2a7JRX2XLTrH9hBhPw9+zasNZZRVzR9BNU
Et9XF43OflpCHKZEGTKVT29FIh+Kbg+0DuvmDjzfTUGnQ8dbKz08YrUCx7V8Zud5
4FjIfi0XVtMOIkEC12U+YwIPAe7Mupr12sokFpS8w+OG5ErxKq3hx+eV2jh5BAZo
ABqiBcDJiZyQRK4UbZZGgfs5udGLGUZT6TF06b48wK3hYGmb+uLVnUyszzA+RZ3t
83ZnyS6lBJUqPuDBvGbLX1lqyTrWLzqPhClDpCRnnbAhQG7VaA/nqieCO+HdqiBv
hywIdfQJfpf4uRirNabL9gC1N2fQRZGSzyebssXAsnE/TAtsCJauCo/s5wAZo6Lg
i35YAvg2rRFQa2CwSN6HX7Xzy9RQFcT5WrK7buiwebBcZpHoFDcg5Q/UkLLcHoq3
sdKqZKc5HZ1lUBvl8N5+ESTSxv0BKFxcG8xBVSVy/NYEXcoaZM/6nK4+7wP2YN4l
96DKcF4OK/OfWIo/8FDdH0klkFVEPH6OC86fH6qhx605iasHkgY6D291cHBeZ819
jOaIr+Ue2laNbIMUerl4Te34B/BAgl/1w9h1ekID7SzKuAO+snXj6ZfdWfmsYLlJ
/Xyk3NUXDCheQr4/jz6NRGJs3Oelw1Jltlzht511582Eg+0wiI6BkD475jz9Zfap
r5N9wDkxoGyfQPsABVFQUFQbC7gRN72gqQwHjDiGhhkjldF9YKnLD/cL0v+ixLPU
rVZvU/v7rfh4YJQ9UTqZ8wPJ7PvVLmu4QhtblWvrsizKcuUNtNYhNJEdQYGHCEgR
THtL9Kjn18xndHFrqGP/mALvsE0gCOg+b6kIYMRnCrJrpuKZpNnyDCDaLXpo8xSh
bkkfLwcujyg29nPXdv5QWsoC7A2lyt07kINLvggFWJahpV26fK1b9K5kKJTtqQCB
AGktryNkzBvZu82DXImoDbT3BjdwR/8Jtu+u+QUfOE5XxFNb1lfbZNnNm9VbnbrC
JoW0sHh37mSiiG9bnzbrqkBgQ1O6Wzg4o+FjceX3iaf6IzLu5rUIlM+LleKOD//6
MsSIfqSQhfmwhfxXiRwGy6mCwkQsSthavgcwkSoQJPIvOuGpE0P0P3tf9qGFApwz
6EkIiDgfVaKG6jT9vd1UyygMgbybda4MsTIGLfo5viqdcXSiLQB5mVm374OHrtBW
jPTB7Fo7Xw8Yq2mbf6S39TXHoCpkP7EigNiKCXd1d0pyTjmq21hgrzbPVnXDprXq
I0pd2KvJ25h95iBg1vEj72shrMVZzRpuwN/ZkJ7skktGUkRZGQyqBdESL+26esTk
lS1YO7efrfGtYbJ2VYpJpIsCsVcDBCpzvsxnGXSekqBRlXbyWv1V6Tvzy5wDktqq
hJGHK6JU88zjyVrPjMpeGMYeCBjrVtBn2bSUtjCcr/8NTNkvgOFf7ygQkgjSxMwP
p9QCuJzAa9hecEV2hpaxxB512psXGEhFukUz9m9Khrvhf8EHhWzw5Z6BSYKpwUTf
uU2ZtVbo382J0epBEuVuXD27a7TB6LBa8EwquaDeXB39gQGMkBLhhCLU0nz4MxeF
SGKWU39nZFS+JOHL7vAHujUDsNjA9gPq/g2FM6rukJ/OGdFd6TcAERh2DWQov0Oe
PbFVIOCHcD5+fFoMRJEUxR5+5LgHkv59BHJiKeg+5wvaGoTA55rM3mr4Komv0svd
PLFp4RyZQMY8Oc1M+3AJzPqsUQbbwuseqqhgEXUxgsZQ8ZlaAE+R1/eNOuvEchTy
b6gxe+DqrqOZgh8OicUNJPm0tY/q0/V191a5kCCmpGO4sHsomSnt65lqe/g3jmAI
upXXlKsBAv8gMAF29lFYakNkCytAGt39rd7q2jauBA8Q95+gc2rrfeJRuAbP+syd
8DSw+FM7qsVwUR7t/E2FuMnAootRoWCmjW29TGXN7MvjayRCtk0c4MyXsSf5nVaI
HR44Wj4d7iEuaK3VkiQeIhp2wHEciv5YeVAHs5leKFpX3T3qygTZ1QgIekS6RPgw
KsBfrQ4tSeMaDn0KOKJJ9mGXqsLBZzhS1C6OpdKbmCUXPVth6T16Qt5qFqqEFPxE
zlnVILkSLmSTqa82cYTQQymyNq5dO5rdTEY3InBiKaDH3qrtIFxafIlHAO8mXVX6
RD55fYKs3uKHQkYGuHvXKEjNvcoA5Ava2adOmigvrcxsuAFKkrs8nzDrr1R2OqED
72mO2eg0Cqf7RU/RIpeGRB2v5cMMcvdBBo+2EZ8Y9EWYEcYrpNvBQiq0Viqu+Kw+
hYfgpAZaNeoE3dV9hGR/C7z0EclTP/ihfW3HgJMCAWJ+VzAfNej7jpN60UFN6moj
D89jQ9qml/+tpBUa8vc72W6gKfZYsS6L3ikfp/FhpsbedtzYt5h+237J7CFWHoFb
VQaG53S6cGNI1XCYZ+q1WynGaVT7iOVsUQfTXVBc6fwx2cORZyiBjZMRKmEBDPtS
C+zu+fqrZvDVb5IZ6+vO6nU4/QBGKyniCaKp86CgKwWGvu7rqG1aZu2eXBtMYVFB
JLRnpxzPbLnuC8K2ihY9URmAUdoMXksquAh2ejgW8c4k0T3uH+EZOdMmIEQSMSBK
NkmEBy02ZwW6u0BuHg36MSb93ARafDkN5w2q+GPxHqphkoxboeHJkVeDkRKbGeXo
VyUecYavAqyCo9NwDdBgf6VbNAeex6EpDOZk2W7QG36et1Xn4kyNrSxU47tzrHcC
ELAphTYfzYqnDAmqteQojmtj1Vl4UKrXHC6UOL2fxxsve7Sm65yaK7F3RPTMz58j
De+MtnFVblgoyAWPGMWjVjnnsVvH6OoKXlAoyJz2IeUekGMs6pzcJmg1rF9VBxfB
ehvlaqeOMfOW+4JaLaOT/BhacX4G3kGOmUj3b2oPGETQWfmoiew8fC+GphOlHcj5
j4d76jHZcEx9MHml1cTCGR0UshxBfEpoiLhwE2z57IoTCXx3HKYPHpFm2TI+Q57x
WtfkIi0tNzpv9Qrqy6EZqOWWM4dwfWywwIY5PxTPVYURz5Ntg5zErTSV806FDDJ7
QGPSj/42PZYTZZEck5jtignaLiEPleRT2Ktj2rgjV6MxYZZcG/vlTKMTFJyFXoVR
h9SOlhx2a2p2loEea7niegdL1Q5uVfWV/0KMlJRIib/Cz24YTe/lAp/FLPWYNP2v
NnYsvbihKMxTI86AFNI9XEqo0yhjgPyDfkUVBQXMYuAq1OI9167QRCPUm35h0uVm
TI9J8N1WnhJWnMEslv9QM6PCSAUOZ9vqsUKfEEyDGIMjKDx05i9YbrWyL2EAkcfn
VWtBWlkjbjWc5QTCrQRKNbzWvpXK/RrERNXKE1aSpT9aErmXksmvP6U8D01Km824
t4QyPYxo5mxYXdZxg7chG4McZX20LmUxiOTKAOPRzoo61tjUp+dkKAtTxYlPyzXg
p3fiRD3TCTECD/uM9bM4+AQISD/hAq1sNZiwFE1je+ZkQuq+F4mnH9XcArr/ydI3
7BUg2OqIjJRnKCdr6fp2GacDDB3nlwuZVzPTBPqBK9e8qOpwCzYmUGJlASVSIOOK
Ip4STqnMK/Dl2JmYLez1YrQjqdbiCOsmjjzLq4MtL4SNeFsToREWeUAR2oWOX+IJ
Fhia3CAFJNNS/sruJYsRIWN5nDMSffFy7+Qn3UIjIeFhNfhAZ+C/RCU5EnlISiPC
1FUWABr3g8ezrm/CcT+TsFnoRIYTrk6LgJOPsA9p2xpQSJYLYPOiKauq+GPRe0P9
lBQ5RICguz8N0WeO7cFsIGYzwqIOZa/UCMZy0CUPNUZ6+HIjCQW0DEIK251j7UUy
Wy7wtNWi1aCwmpwUlvUcQqj/RknsVFlZVJMMxsPjbLjdr3ewD17HXV2bL1hTwcT0
VPvmfJk0HZ4mlxc0wFvuQXQYw/VG2Jg8KMrFBOPNwYxaLrWyvt0jIuuvVVq5eG/p
sY6ynXYlV4mDvZJBSQkOHl0TB8lBocv0JcNroVDqrBn32+Ff0r3/yJsjm7Nz4VjU
5yGkfF1ifDsPmNZKGG3WwMRv2Kt30/kZBHLFQK3R/m3UNveFJOxZa4uvFYXuh2LK
mE/GkglP9lRsFL6BhjB9uGoo/mAgdMnoLcNX7c/T8MhZ6K4ys2JUf167kwwRtyyI
GBJJHe/TbItYSztMDe2vnH6m2/ymb9xWVTXDlw2U1YVDyiqIno3/t+CHi2N23Fo+
cVj0uDrn7i8gR1qyPRRn5rCBBxxJ7c3glA/EgD88hK7joC0jt4hgMuWctb73E62K
A6uqXhgKagSeXqahKn8eX1aOIG1+wHYE1+lheLQSRGMYEqsDrEU3xB8xcwzGtVzn
hJSQax0Wfn0TBc9Bs2F6RgRLIdiSEL4WXk+tjsUOwtDKE7yDdM3RXJRJcEGyVNG3
USx/gRwDQGOQs3ChWOaDTZXe5npLH2yjLOUQiWrgXKCCTUP08jQDNrDkS2tpxfjV
gFQ6wN2SIM8zxpigmFgS257WiXapfCTjDh7zM9UlPOz2dzchGqlVhvuePebQPfP+
0pj7jNVMewgCknfF4QdOHMSe508X3PfCPI4qQV3NWMh8627JotQpha6CAH9X/i9r
xzJ6eCCnCZMjwgHLDQB28Ce0Jp3rEDuLCFzZBWSRA6pS7ej5eKszl8Lnvz0eW0O6
V0ysBnmrvnJ5C0lVTYRyf6TZxqsz2gIu9jA0SvSlB8X07Rl4L+Us8q+vRHnl+KbZ
3+G5m9NzxWCK+sD5h7JU8G3WJRbw7KppNUfCpP/nyzs0zD1cgNTzNEWTYcjnnnpd
uJXRNmir48EmGqnI6/LYauqHCVeoSBIs05wNwPRxbv/6v7G6pplX+VHl+9Cq/Bdv
bRoyfG/cUlC7CWg48PCvqUhQ9fw5/IN2+UISDTDe2+QFN8QU2ujtAWPZJUCKw6zd
Dl3DmGzubVx9kcPpfuAVBrmwUuRhAp1HPKJiPlMpt2toCKf1HOp5V5MB+6M3zcem
JGFe3zj6IK162gKbkWZ4Wscc3IXqe4rWTjtrNDyQa/OwIJwkc30ANqla5IfDr/Gu
dRT+uLbSV2a0U0ZtmU+D9BzVAMMfEtaqZCfTmCV9QQbEuWqbvVPxBEf/YjgFa17m
hbEVo9RzaWw+Yg0tIIan86MrGHSAjlPSuXjNxhqoNqVg5354X3qCHwkUV4ucNFEF
A+0gUHSNN8fhGw8wjST0+IpTwFvz+XdStAWng1QKK+HLuTVDUCr23sxFkFqofQ9l
XH5ShJebxBaRlVFG7vu4biQL/sXel82FDC8qy7/PLFg0CbyfJPHK8ZY6tCUA8wvj
bpKIMcsvW8xgZRskjKZDZD1u+7QarUhw58Vkx6q6zgVhcsmyWnzCDEG4VdW9ozBF
CkEsj/2qhazeYZuStmhzypXCWw4hFVzKS2tonAdTS0Arun4RcuLGL1PU/Btl4Y8r
LyXMFLP25B+V/hpkrVl3EFN6S0QwDsjlr5MVmoYs2dcJU6pbD9ZsYGDzPAI+i5gF
WaPGGLE2IX75xXan4/wRmP9kv43lpr5mdxJlkJusVHj0GxtyyoM3VLD54mNg1WCO
RhDo021RdTp+zpBBsA8B9IK7QdRoCyJPQJmNb8rnK89HS2u21+5zO7vhgbxHoGA1
iK6IHh5RSuNdCNThGh2C6w6FCMMtK0JLIVpSMBBeBxwZ8pZNRMxaNYe/bDhL/oLv
PBZ+YjLSQLBeaGrr0NZwKfED6tPCNN4XBUnUbWGfZzb/lRTBXB/1Fero551r1KGm
vkTkp3V9jGXp+Fa3PbXoEFug63UrhGhrNTup/SO8MNp1F5FS/m72pbinNxQ/Mq0c
5l4cNOLHLiFg1zRAYDZqs3FRewtJ55U/V8inH+Bz6o0I/c1yeHUe4bgH/xNusqd5
hPjFTFrJLfjbNxYHdPJKACbCptzZ297GqDI0GX54DH+gKvx8DuDXpzz9ak0zmvK/
E8JrvTO/3W6Kg0aByiCa1cxJT/wODeCkPBU70oeuzV6o6i1ZZV2tGX8n+hZZV8Tr
C9al9yjq+2sGTXnpyg2lpeet2xjQsEcJ+C7xXZKbEoEulO/XJMpVMvpU9wG/jpFv
wxthT/xJuRGCwKG9+H5HNpwQ5AfYyCHJbKgp2bwLhhkhB/+igWKKtNEBUUyGMUvv
SjLWyW4knt3UpOPfRwkrQRkg4oFIAJabr6WGEbanrbzBFNS8MVWVyQ22LQHnBuAX
K4UT8K1yzeZnORpqt9tq47zB0nR5cb+KGiC3a0rXBXiyFWA2uHayPeazIcXuzW07
GC77qXTAiCPOynxLWVslWgx0Mb76Kb8gAzhS1U7QumHWQZsL6X6jJowNQrNw8nlT
MX7eGDMCzUKZMg4FKUimwfLDHDeRIgF9WZy2UgKLzD+MjigcF0fzPyYZPehf3Col
8zD6VQZ9L/KQ/GftrkNy4juiFdCjcznSJMIvtjt4PeZVykoFtSBt7rC8dT7ssTRL
RNrygrx/GH119Bp8yJ9HD/gTx0eRE6gajEgKJxlzrXYvi4avwj9IaIKaa+1cJU3x
3PyzRuglqWY7kYfxMdutNT3Zx+t9qtHvCYXqNKb3Nosn8eHVtuBn4G+B3XPUB4wt
HrbHqJwAyRkONhpTl7RQQPWWEs+c65PZ2iMFNMccwwdV7vgSXUsBBYhlsWDYbbCe
xEuHenGNL2wNvmXox9OHOxChfpTwFCy5zh8MZynthD/30jlJpyP/FnHznNwewwjH
1HihsHrLvgDrVXud74qGRNakxQ+g4/bA3LGqGu3N/lbBRihMb6If0X9nAxkq+F+3
PQcaYVQzetqy9vdp74nIguS6J8VR1UPudOmcAO1GA6aOu6U++vROttNXGgvcSpFL
RdDUpOxJoIL0dQ8Vv7NPVwTSnViQmhEq79HrzI3egfR6Pjss1deXTGiUpD2p7DL3
k7QyM+I8unjg9ri6BQxdiTwaAERLs63aUfnVARHypNdgWB0tA37zuxH6KbmVMWJB
bAjOqh/AJjmKyHr1lhSSItx4U45LNHulp8AMohb+2AM+MPPqa8WNLA/94O1GaWNh
AGFyj1A7AKLnA3qVbHidcW0mbS82rfO7gcksepGvnYZ2FSYWQ+yEv9JSFY9C9gp2
p6VMWkQXQK7HGjdwjK0LWmwagdWYTmJzbmZJAxQ6WHIh9qJg9M1zQkPV4Ne1s0Vs
mYY2M6Irr6JaGWvBmuxhPSkOXF8FW+OcXrMBeDtfqMpNRlUvaoPbB8TCQlsWudSK
Pdcv4e9CKH+7BDPbKW1N645+XCSRemEoHmkjHWVcxJdtovY3P2kHIbQDsOZ792dg
qVY+weUh2AOIriUjmDQFVd08ywhdeyOmtD3gnfD+XfMCVKQtCwM8JYhakLVuNO13
7p7+SjZs1NTS14VpmBmj0g7Q229Pdybl7MLOnOK7G2U6TKdKgT50NHhVgumFpQTT
ETF5JY9bzcXjGLdIKqAc+4uaFPMPODgRU2kZAcMHNWPleLJjloiYlg1jf9lou5rb
hdpsS4p+lawbZ8HO2cgtO7N883i6m0XK6Pv4eeo+SOmq+AnpXZBEvQtmMUtBg55q
fcNTxlNCT9c4alTGM0ipRwDnRX3YCXSVPWALlAUG5IBzyv/wGnCtZH+sJk9kJevX
41n//NRmGzNXDjl3y4/FpQvryJjz9NTI2eN9JAb5JUMOTrphLtRlUBRirRN6WZUg
RXRek/kItV2qNSc37qQusQ40wZcBZhTxJJbL2q1HBPssKU0bm/4VvR3QNy8OGSBB
/5+g4lywXi7cZLhzXrLhbkWEefhAbXRmIKtccyQFuMZs4vC0jfrPRyP+nsZjsJ7m
nfRcuVTquV7udwqnIv7ZIOnq2+xyR0o5erRpnEmzJ73o5keZHuk2k3ZXzhvs+gPG
euszth6KDFFWVdvZ55VjPkPOCX4D5NRkwmkRP8OUBf7q5TZpd2PJ1zAehvRGO+9n
CjLP7xCgfZTucbl8Wj3ZuQI7zgymgvk7RJ5r1vlQOXUsgkHBx0Zdik7ReyXRu3lz
hW6VYpXO3as2NnnBAZ8Z1yhQ1pIsrts/2wRjmMXxfWZKws7846MJ37yl/tHCX8XI
olGZ7a41oRvcZ17Rgfc80pNTqtfWz43MrmypU7xRtrGb7pXhxKmzIfOrDT8J258/
/qPOvd4eSqIY0vhnkx9vYKMOv0mkgBnIxgRI+NUFSlE2apg07P9bm50BSk8s1QEs
XmDqY6uPqpjZ8vBlTPzazvdHxIDug2skkBGFgs8jtfLN7ms6ovQHl3XgVKsHdrEk
NwMXpTUFnEahBYr6iB9EjGXA//Z2HMGyr6E1yka8i6jXw/L2xwCgxpy+lhr72b3w
TXn9gcvSCZ5kr/3q+hu12LgVZZmkzVAgewN3WhtAA2VMCAi8K1l9nR+deyjX0a2C
Kc1ZCzH+kliH3AMR+y4iVHw/+9PTUc3bIkQqYLovKEuJu8OpgVPL7V1teD/XGGd3
P7zoY39ubIN6eR6SsTI7HdKJsS0joTWvaBam4Hhj9wri+VySyfB5zmPgB/+Gp+VZ
WF901hH8FkIdcGgdVYgcS/t+aDpQtxWICAZrSiNzPOWJQtl4OYgrNvOZgVALovKZ
A54luIZoG2bLiQ82B4ZdOh42OiSLcnQF3EvttSDWV9NBWAg+mawAre5DKa2sSuTF
puiL65DV1n+XF3IoLW8D2G1bRpXWUcInpl9sLzW+6/R3BOj6OGXT4OGgfd20ozqq
4gn73Gn/cjO1QZ/cJnfQzWqvAB5uUnd0lCY+Dg7vK0zwhOatwOuUvI706D+Jv3au
dnON3Eq22wGqhnmrT6HqppicZ9DGF0ZqYw/uH6lZLpsP7LK3mMvbNHLrlNbwSFsi
WtM0IuC3WNy5RCB9Q1AgbnUxyW8nE1TuE7HTKw4TgvIKHPA9iZZFLS+qsLw0hTVK
eOA5o9G0TedzjMuMJegVZQ5BuR6yUoeznleKE29uXYM/Y8wcCh5C25kvLOFp1l/A
tEcZMsXbgJKWtyREbiZeSBl72J7/AmtTkLtIWLCIPtfp5ZRh3hiox2hqUEXKfEwM
C27NKjZjyWJNyhFNVRaFA9W9hSfGGaeU/TkJ/Z+O6aF5BxQKB1BDxVSwLVZMyLsh
tlo24ZGhZWcKL/wF89rRnLCwYeyqRSLq+litg/1J8UcZFwn9/7EjVpwEJAPAu24W
cb3FS79IMQZ1WeCECxcpwXliJP/3DpEzo6HzfwwAt6KGscdip8mL4UUCGRvM+ihy
7CCrv0GAscYvx0u8lDBWb08y8SonPDNOB20k3VNUwmq8rIk8ZaqAgFD8DIXcTNX1
1skbrNvqwY4GV4xjyYZYhSFVUnFuN7fXIsdVqYU+faOs2p2t/rlCcyWdt3q13Pjb
w8IEEJG3yFQ7OSNkblGQnK+Nsl0rx/GCcde7DOD0qWI324puOUDKdi9hJ8HsYc0s
E6kfsk3/48kH95q+GggGgU82/Jyy11iFJGOKa/eUupajqpuVBPzG4CMMX3GWnBjz
cuI9wc+jY0oMvtqk7EnrZbycMFtefp9APobBER/EaeY/AWBvQs6fzTiYzDRFyurc
vbuXfPamQ5QZGHZ68La8Bvc7vhLVnriJjHcADSnRytxvf+CO/JpOXO2/ogbeTj07
LThzVgddEuhEQBlOy4e0gfGU74xN2FOZn1akIUhwitD2f7GNZQlFZQOy217o2hSo
BnIgTcNeuBxbAmLAKttfjwGRgr+kDXUnOhbBnBqJKkrQ+TATAVNEBVH14yAAjyr7
t0nz78MSulGF/RijjWmD5s/CXxEEdnaeQ3uZXd9JjJRwE1tc35Sq9liQooaY93oz
BP6c7FAbKUQt5QJhhSZMcTZ9kMWOMT4OKQtZclIMA8pKDqwXH0iXYYmgzI6a64ks
G8T4/UOK34d9KiZJEDWjb9SB+kMdbmLDrOtN6pKm4VWSWYcyNq8YMpmOhR4YAT3W
iwSWy8g8NjtSs1MxnPGooWhhLy+jDyAlv/gmPHiMLeu7POwVufm87JZ4r89Ad0oa
9jtkxTsEsmD/1MvvmzA2YoltU3pXjRIhncTcuyMgQeQWzXfIMvM8+oOr9A2wG+Nr
3PJ8nrsoc/uTa8hH+gV3gzuPVWvy5Gr83/E8Ypph/nWa2lDw0V4UXrcEiXOiG/9t
ojYkLAoPpRPEV9pVITo5btihl5WnlWx6I0Gtsi6lWVNvLdi/VDIIff07gyxNZC+d
/TNDGI8ll67OuBJ3Tom4AR9PuQdfw4rbKAljxw6MtCM7NAyyyCv5iVgtY4gg54Wa
vGygiZQi4To8MiXYK8dqnQ1amSbIvNmGCpc12mEuFHATDI7dkHToVrpxuMKdvkXJ
qpr8Y6YQWo8BGp82UnnTLdVDEXBvfqojGnN1UmZk9eZmUU0fnbeCtSysRyPMUQGl
EEQyUNlRPDNEAJwi2NFeY6JkKuT2EhcltRPlPpoLh4K4pw9xj8SVhwT2wnYsdoIF
lPT73CDDXVvX/EvJAIAUOvVq8fJGcKtVkdll28CYx11tT3L53/5Cp87GV+JExObs
PpDPbt7HOXI7uDHQsCji7MuI2FxIJ1ixzjZ7LS+yJEZRUeM/QHSPSO6GSfUUkH9c
YvlBCFYHmQTYPetE20ypPsek8QMOmfiwbuiP4Ip+TqQVGssPnPjuhPAlwUpmSP7V
N0WIhOLl9f4mdweDfubzAayiICQCPwHx+AeYQGqggdU8k5fQPH6kNDhf45ISolH4
M8DSBe4GZ09V+sF17RPueLjqIzIOwYUogwxevomBKlZQZuXR9Y/xmUg2CXfye7FQ
oZrXtTCd6ScBjeVeD8rRSUQO6vzmOcFJzubusBOCpHFgZV3d9VGOOggWSyE7YJNX
6OPQAW+oeEOzuKjB1RI0Ly3ULdUM2gA3tBjBNwdiD6gXxcQEjY5PyAfsD8zQkDxA
/G/+8RqSbyE3NvZslBRgoCH6DYmkjctcd3d+iqwG8lUoN/thdSw8H8X4f4SYXIK7
oeqwVCXfBp0nzF8qa6PPR+tBAAIFKTtFXMHaTcKCh5MGnpQUMQz1DDuJLgoJTa9K
ij6d/mMcNuFebLtHCuvchxUMkpfl2nyQG2hJGhGYlNIj9kwdaBmWuHiV4d45TeAD
G/ljauE5R7A40U7ZDZgJW9e8AZOoc+PfHGtAqKYVDoVtL3dvmYVa1zGJfiOdQDBX
iTMixDH5ohQN6emdCpP5NvmDQCiMKWwEvJU71enHpHzGLcdHgx/gSxjFW0cz9wui
9xMVDRKCif4DTaNxsQzkVApt0m7WT3pwSD8jxrYGZY4RhVH4lAy0Mvv4/epwOz8l
VJXEimi7ewysKRGmK6FNmSlB81D7nBmrv7ciOoGLIkb0HlRIxNLa+zmqr/6xkFlM
bixN/KEz+msLsH9DdH3wC4ZX1v4xj3Ul/xp0Mi3/nHEth0ZtPyWjTPPlgXG0Z2FU
nBih5p1quLlKnodghqdrma2Q0SLnSFuurs/Qjn64+lm1xLxw4Rw++sslwqWV2wwl
PEQZOfbE7Sdm9UPr9AFmqGLqFNojLwK7KhKuHe1JXbsKAYec8MyjqgUNUsxdU2ls
2HOaBFvfBtZk/6dBAq0AA5C+k6iOafsYQpma+qubI7/0BoXDZNqj9LmRO47eIhCo
L5QLm576QYgL30IfilmcI7aANUJJ2KPoYYZ9f6Oto3hNBduS8F211gQz/cuEIR3L
N6qUqjm8vTO9spZDrH49OBGVqpUPtREt/PNJCuZzV2dxTIxvhIOSWMdn54Kf2xrp
uEnNUYzebwQVlaghfIYrmF0/eSwR7xAa4vISXuog3miaC4WwsJYLg5ClAOpfLkuB
UBlZkL5pD65WicJI2oUAdSoqZ+tne+aF1QS4URjcQHkJRbz1RnzUXWPbJvHT8z1p
VHTl++VLwR0LNqx4LVYS6pte7KCTAPf/fZgn3zK4IZ6A6E9deaed/Z8h++Iq2NAU
3ykkxl/6hgANvlGMR3XFaUFd/piT+nBSvatFiwWAuEF0rJPcC6puF4CCX85NCKtM
FGv1DVZdoLS4wO3c6f8SZSePt8W6UObDS30tH+B9B34TXzk0g2K/JFa7udk+dbIx
yxfsvAA+oC9Ul7r4yDMCGkL7DDdfl9MwJ8DtVw5SPFBMtKTDDXpxHnQpOyhEzHCD
yvUW8aE1XVKZcyZyyln7/Ws6Kk7cNV0fq8XsFLLiy4v2xlGQGPH3l1RhPSONtqRr
1RP2KOkhTqQXAORE+c/wW3X4ul/gPcJDB6ibM4/U+3QQpJgj0HFv3Hv5tLTGVL84
bynTlDLKSuu6tsfMOzZLKT7709j8iFy7Oqpst1ihD7rJh6rcHGPetO/oV0la2VCf
qgxmjbu8OrrAE9xshv4TqepqQoUyQoQhOrbTBVOZQvessAc5+53SMeaE/Hk6O65r
IGy3SL5XcFrD38MqMF7LR6HIDJcFWWf9ZZ9YHpTg5G48t2TEdGovjXiDPGI55TRB
yu0pUV4MLctvyfo3QHpBSIY0hsqVIEaP1/Vym7SKNBz4dWah/CkjZi7AG5Clbagw
JgQ1xth8ThHDKrOni52wlvFzH+KfFRi9X6jkisI2uSvWxYyNc2ZgQvwJK2bYIp19
JB/japHqDhWCNJ3o6DsiMUksUoFtysprMy4125772YX59MSlFOPzS8jbufgN5UjN
u0Z0xUg3lZE1xml3y1cAqVmNn+j1Slqwb6pFW48oOdbtNxkRM1MC4gTHQRhZZv3O
m8oHzpdzezaVRqt1x+RqErysGbzs7P0cF179QxztwUHjOO//52tbJMF2PCOdFyvq
wxfiqZm6FmRB9Y7tk90iY4kjsOjGxEuB8C/xlqmYs9V0LvPCzHaAuILZcwkNa1Bd
a0oBeYiKUwV57jGqURX5usGZXEeMvTNQctX4Wa7y2Nvdu1fi2F9zaFjjhrDUNzPM
Z5JnPGM3LD/XIAf+9OeOCtKAfrNrrGPffDAeiWcJXeLzG60ef/XXtiH+I9FiFm48
EL30hgEFPCgC2FsULCQ7CnE0QwfXrr2hw1Fk01XnFWNRgwVVOuVqZQ/8BUitzI6e
OP9iDSc4EwlXPJ7U25RdBGu3vDAQPK4/BafJmyf9EkN9dXr1GWXHCGE6gbcpbof/
kyPoFJ5WzMbX41VW8mFQJDzpaJilYEYQ9q5xNbqL6zedh6aUUO/WAixBV/b7U7ps
N7yIJ9Iu/HKPhtHUfhocJnh8beMPhSXeZpBxs3fidOST1IGjXIyOHc8Yur3DzJ2j
iZNLRxscwsDupAiEukHiIFq4Bd4qoIBL8B4f1ocqhHg8ZLqVA52SL4Tjy3ncP4ns
Kx+t1HN3MvIlDLgz4ZVnkywOv7pmY7hMg9pCJyYxtQiRi0sxvQ4jceJDZfF2VkEm
MOjujKVSMFYwi/ZdxigKlk/CpjZeP2GIPZjie0y00ts5xGfPN6jLwhWp5eU4ueMZ
rQXd3OFbahlpq5lkIZP+LNvOJ9UaPAXhPHkMdJZA1XHynfWed+uAvSBBP9WYXHx5
OxWi8EFjybDPbEMtC/v9g4eJHukIrwLAkrMPnZM1gtBMtJ3goNiV4+fQNuEF7ggw
OChs+1pjH4u8IpvC54kv7OmYx6gTEcimm+ay9bP1qvGjnT1o6d66GlWdaaVMhLKs
ESPO60mE6RqJwJ+tSYd9aa3bR/DCHz1phSy0SKhCz7wlmRermgkmwG75hOistWtW
DiQmAyuoKrVk+XVQ7sGg2jJMtAJNiZ1s9vRK8tuS3c6SF1cwRcQiL9JBSg5lxzSt
4XA+xMSvrOk0/R8DiECWV0l2rrVGa2IJCF48XD1DIRaVZkiYaWpJxgFP4vMKQ7QT
AtmicgDJmyLR2rDndk857CnRxygsUiGVHVTayarp6nFMCcwGePHqHtvu8xcGcfxb
RY7+2k4EAtdmVCv7Qw/NOqGa+s/Qy/7oo8vDG3xDykUfW/QM/sL7as2IOpBNXiEI
HMP86Dzr6U1XeLTxAWNMIlVgQ5ARXsbOBjkMaA82l17vs2VSWPvngftZAQbVzF4m
RZInPe/DDwSiWwoFAYFCub5rw8Rwn/q3IX/Gg4ZHzdYufN3qRVHKVaD9HcBP+1DQ
mZGxlkgg7Zbp6199e1WMaB3Bk69ex3X0z7SfgwefpyO5W1OjenjcveoVrwbED0zq
AxgrO+zY7rAE66e/Ipk8Xs2JeCJ4DSIBAoG0VVYgDuj6Iy2+L393iYnes94+ugAB
cf/5eO6s63XTOcSFuMMDUy+Z1/wGQNfMUxpxf5lIEqIDZatOx246HD6MT0wkDuVL
rYUrWFzFk1kqrWtt6wQK8Syk1X6GCJp5VlfqElNEH5TguZnpCF3zzggsP3A9PXXm
waZU6g1xGCK5r6mKcmXBVVpRiw1H3Sn3d6LkGemIb7knkSIZWPogoS5XXjlt6Yeb
9FZiZJ9HX4lEVPOLvQrajKQzhJYY2Hr4sAm9S1D2QXprBpuutaoTHUwM76fcWTpN
YplitEk2BfSNcBvXG/MwMqms/y7uBLBg4DCa8pCNohVO3YkGLPSEMoNGX4hwaeui
WpsG4aKxb6qg3/EpoUfZvHMnx2FWx7F9UNiGSGMzD9/qSbtADbf1sId6TZsWjERz
2c5emuvY+TLmcaUu7YV9esaBslGlcTS1TW9Ze5oXk6VXt67zfPMSUeZmsKQuo/Ia
8KR1sU82XJuMrWModyny7mnlnAh+OoEgtiGbYptNVugqH6UE0CNcmz1AEHccOa40
kbB3bFr3LPBgnneujq3HVHbDU71jjGiR4zRFpoTfD1oiW3nnZ68rhL6IgZYoSVbK
kd3NINHziLzjXPYi0lblg7VF4As8dX0gUI/lybU/Dgyd/ca5HqJWfo0Ip+Q6gDVH
EF2Lg6u6UTkG+rZsV5LDmsCcL2ptmzquTbNqMvlkC24NmwwRQM6NQXySmqXaKEhf
/AxcGo07wbGU6+SA07p5kRYQQLm6DoczGzoaRnvqQQdoZR7OPEtNMAPt3lgPneTc
cmCO9UToh1T0oO6MvyM1w7nJIjjmh+WEkvptlu+5YZ5vo3GLPoqCu1+hVZGUjcKt
UsOJgDV//S60dBVWpXbh3FMt9DsS+vaHHNCltKLgQU6YyxwxKmlzVbBFvzvrrjgT
CUhG61QGwdgMK7hWw7L6Z0+53IXnEuZySszoJ5XAxJba5PINaKYtKBrgyfH73/11
D7Q8600wragLcQX49kVaynHDn6bBIrq+WR/NN1nP0ubC6LZp357GXfr8Rcyh9qqo
HQeeGH1DsE2NVt3prb8qz2eEDI5mF5j04jugwHUQbei/56hzNJ/Z8EDTvhK0JL9z
s4fG1EQKmSm+EYNhZbEoRTGHd7dKtm5I7BhTkoEojUsWcQoweR+uWEnzG8OFfI0/
cf2lcSpjGemfKoWWODLjTM3OENimFIfGcESno545RIA2MLCax3eKKrtE/fKu0T5/
1jD+U3EQqES6V1AJUfxVpAQDAq4QcHXB0Dhw/H08j0R54Upjh5jemEMrgfGKGE7Q
VrUq1ezLMebPFj4Uav8TsNtr9vtW1FdyHLEAffswWf6Ee7oxcvXBh7wIrldVbZZV
nkbMrzTlumaIFIyNz5cZhiQ5k/pNfUdsRorpPykv0OlfEAJVmXo5/W8hxDf/Em/w
kbwBKcMGvpQ+VhEjZymafKM1zRf2xl0/tzmaYWA+k0YQmHcxU5nwYEILCqIFqw0q
fdbPCs0CvGkdiIfBGizrZf+1utFNZnNPEfDRVRhwPSmo2olIT4czX+e9IeicjZFY
/7g4S2/6kN2b9Ai3cKLWzUtSmR7yHvn3gYzzspAbwL04CtonrnncuaJoJbg9ke0m
zMtFbJM6PQN4NfFkr99T9EKNer8flDKGP8sBFHAgTNJgP4xBM//1m90dmRlE/opb
lx+tpxUL/pIH5dLEOvDdzqDGPcQAMhARx6RSaUOFV+YSZysWMz9GkBu1nczuR40a
ZpDIgUKb+zdVSLA35EvhEeYyGUIY2SLsmN2kRWCLGkHpGoxOqQbSyogUdjU1Gpu2
/QTau4OsQM1CTvBiMWGa2AnC0s0saaYn+KSp6Bb5LXMwpsjFaIVmDDS7K++TkwCu
unDVxz2TjRUYL7Dugyvnu7WUDAObiBwewZC3I8sTnxuPheiL7EjuLz5E/6IQuyIR
rLR7aDnduWlq+LrthzHAHsQxs5SLqDGtosoFyJg8UiibJCfatXYOJnubiprJaASw
A712Clr986iOgaP9/CgTjvn2jEZo6VKKhpQUjgtyqgAZ+Ewl0RR2z4dYeqKmCPf3
bQiU0e7TdXKTKwWwAM+wsstCXVN2RR2vES6tGMdU/J6JPdxHbMXZXS9+wMXN+Z4/
AmJZ8+eO0am6NZr+/f2InjqL1U06PGaLxXfK8hoFOBR5ONLOiE6aO+bUAAqvWWFM
z5KbMz0kW5f0fm0x1t9gxUT8iM9TTgQ5iQB0GMCf5Bhnupsw6zPkFuCbwY7MuyVj
VlwewG92ZicVK71xMhBaArWjimzF7WB58cPHwog0yB8yKuHNvXC56DUH7CGSqMco
kTcwlExEW5vEErU4vyiQ83CJFweT+4PcYeaXqfe3+mtoNM6a5do13FKgdjXe2Wg7
tTqNPHZXUZkWzHTA/FOp8uJviqWQtfdVkxu7NEyrQ3hx218YyRACjNoblRLsvvnY
Z6Zj3C7hgvvrKqOYprgsWidtxKL5Kg579SXQRUgil9o1XZNRrDHodxtl+6Mi7+tr
jnXQBQwThkXIVGpDVrL2032VSAbImrEOPOO6g6Vfrg+cYlpZJi4tN8QM6vjPwxtj
YQZKu6HFgkvplNSxXYMl4uXiZPQmAja1JYWFG9MfUgpqjPuo5RGGMyD6HzrNioLk
RJdUZn/CwLlF3TGqmo6oR6WTIbSynYvSYFRjaDGvVM7yMvL+2z9hKCHRC7Pc+0AR
BD6gzP2b0ILaPRY8xXBRdxuhTd/zPZyv+GoedKVfta87dUuXoVkXjWx/O84gWC/g
mN9UEBgEK5KpPYk3rN6pnWKW23BoiqAU0CTB7ZqaOkuHuQMQ0Jrn9izLKU8wI/Kw
M62O8BwkkCU8fI+jQhcSqQL8TvyH9NH6kISAdEi9jDMTdjW8GQXDnQ3XO6v4Z7Gr
rzR7gUBHPgU2WjlgNELj2HztgODgQqpUk5xhXUjtegtpjc2ObTbGyuvTorcDg6O2
jouOYF3MDvlYCr+GQVouJxzsPwA/13vAkyINK/M8CF+AjtpNT3A0vj/AiSl+vGUj
twQoRorcAtAbkhhgOccYjibuJK75lWKscuV0AcwdNbb2kI98JCLYe5zxbfa8rgQH
nCy1kKCNTqvzv5Xb/kgkmrGVQ918LxwbNhVVn6NDHcIBgZk81CcTqEvRzTnxHoDZ
gCs6kcUph3/yGvjGfhZ9kmsHdJQXzMlNjv+s/oSq0cHgX0GV03gLuYNXFjt01EZU
45l3k7yWz8WE7OP9H3OYBFyIKYgKc3JXAfY7xSmzUJP82XzwJiN1WiT+yMLVJPAF
En8rZK2oINVYumam1y6/2YiYyRNk2e1OKl89CGBgHhcA0qAn1p23B9hob1AMCvI1
XFChPgT8gv9dlKLjt2nO+5eDLtk1hFcJJxwnZAwLTh5y08Wb1SZZngYSmgfRzTGC
Pb6qVZReB3da6Sg3M+dqHYuI4hn6iAd8xfXVINziodDvZe+hi5pP4hP98uzW7KoH
q+VFnA0m0gHgtuzU5WU3HhykmU2Jqs5qm0B6QufZILUYPlFlaUjesGloYIMfUuUj
8iiXl0dLsrCwNXwdhQEhVqRXGbDHrCFmVovr6lsrBQBlgni/dHbTSx/1p4Sjxh4u
n4snqPhdTc58ta6EcWA9aszA+YsPelqAcioBqNn1V12pPwNfaGNbriuh7UeI6DpZ
FSw8tAWfCwAkTmzjQKfSoh/nYeUz+InsAxtquCIOfGyfb6vnL7HegCAFcH2n8zON
YT9dh1TQpJWa+pNnkgN2hJdcjKmcA1517bj3XWzTYXl61MJqeOVIbBjTgndezrEN
KQmabskt3HpIrve6YogXPrZlC6XluKyGQ0PS8+zQqaE5cR30tFJ5clEr2bYnawPc
JWP2bUnJiu2Ds6nNrohrlzJvUBF0CVy/x+n9YgLX7j6DRE+vbprb7U2mEzTDQ2ap
pKpXbI44N6sO6M5J34t4yZUZr8ocp32csZwV0BL5dn2ApSuDbmvToD2DWcUiTHOg
4MDXZ2TICMGxIDAeBRioRnYeGZeDOFmCoEyaxHZztL1hVBccRyYp15eRyp1bWL8O
9mu4G9f9ARSD01qtlLQOrq079yMJieWlspUuO3Zo3VsWacTf63v2WIkZ16cxM+wh
JgSf7jgMhbcA8+Zp3NTmVWBMK4BP+nb4HUHacthtqah1f/+tEBLsfG5TTTJ2F+LL
DQ5IPDnbBprI94uPC3jnr5okn0EYWBTSAlmlVBRHurBR8nxDN/QMnY3mUD2Y2dKi
1uLyb+iLWusWnZlzHFyIfwkWVWNZc0HdQMkxqiifGx8qOy7gHlAjaCW+0r6IXBP6
/Np1cMUv1VSMsUSV0RXoXMdlAOHWN2lIS28RkqbrLVk0FifzTdFgZ61ye2PFzdot
xXmARBlM4J+6U1tGuiE4LLNLIkzAJ2xnwZZjNJdO0WI3ednKcld16p7YVnlThB/Q
lA8jD1WST7WShO+e1p0jmSC33FAf9QHgPgP6ecyhqnF2mu2NunY0wErbdU2q9oYD
3Lb8dPX9xGhlnmasa92DaOkxnwpHsHTdRo0N5yn8Cc/FcJAbXcO+U6vnAsov7Am9
GgLRw0gFhsRHF7sMXnoy0W+nqC77Ti3WOxOtyDlQ1IdzrOmr/fXk744wOS2zc2D8
pVhSCemQ3cu8sWQ+c7224KNRjFfPcfvxCBibx1kTtf4EEjz9iD0jXF8mHYRUCm/3
VV2ENx5KwlVDWb23+HzVt72Rwrd75egOgGONb3wo77xp+E12dVlIHcbpMQrnO2zd
jCCL32ApbtRAs4eq3Q81jF+rk2e5Brvq9m4NWrsMSwAvpjZ4yBJXHU2jN65UAKrB
88Eg6r9pJGXn6MPz3qTMuHrzRAQ0g7Z6YSTe/W1mf71z92sqKJoPkTrOMq/XHQnV
VGo2HlqMMeVJ0MQQvaxq5hx9tXVvubr5LfjB4e8D/uKVGyJGoUsrg4tWcr8TjNX4
1CYXvkr0FVmZKc51Hc+scz3lo/ChXBkKGPZrnGtFEyfJKC1n0o92hpLSiYxpS7kZ
1+T6ZCRC7B7Fg3/soxVfaJnmXkhVcVEhaLyUhIxY60MkY6Yno5wR5vtgPI59fDH/
wUGbZZ1n8q6BOpOgNXZ3iEp5ToZIfir0NZCveQxBbKuKskx0BIlzTf7TWg9emuNS
k4/q0Yvpop5h9xr2fyzn1U6Tcx8LRdTz2K5NE1VQXfdMm+GRB3GUJRh9CqVSDRPQ
byXq3Fx+6TbsygXIqqYRpw3XY647FeejCFzK0fSOiXLnowAqTqIWy3WGbgPOWin5
kpsuRO05NQWN7x/2qael7WjYawTNmTIxg7EOyDzyJWiZDVbVDSwEIyTf7I1h6MLQ
XlQhLtLufXM6VcqnZoVYFotk1LM9gdE46svwxA7HoK2iTOOevyI3hCgQmxfSkkk0
wWlz7DuNNg4TMtK49JWShiBX7XBcPRxVHycTH+ID8vYJEJNYN2WQjlmOqX67wV8B
KeJBjpr92l/STOsjAwRFWDbrBCh8rMbsULcJqiy9wlYj81hN07UUHvl7paUrTJHI
9oa6lBbf0yvz357Xx6qYwUxEE9hVSIDZS5HPNPY70lpfVK8SwFvAifF1vNqeX/nz
rhAXZDHgW8c82bVQdGF1TmPPInEvjchUZrqzyVkhEzMgPF/patYXY6TRkJUPazPL
HKYiHvZCY/o0ciU4KiZ/BeSmVzigsXgaA9EPnToAs2G1Av/m79OrdnXl8uWQXJI/
BrSfp71NFcERXyM3GODUYsK5X/aro7q2h6qPaerIhSbwY2VVtx9ikoiajfNk0uFz
9pk5juqNgFke0NWjF+QHX1Ttete/22DSTBjrU3iMfpBP3qIdEGctx5Aj1Gnf1J42
8DlIVSKMOl7yKegifVp6Pb3ktP6DijgoBlLihlTWSTQa+xYspOUsnTD+wi6uO/je
EF1MW2xJKS/7BmByvPTaYIZFNVHaoV3jinkNeQf36NolRnTFa+zXpgRtyzO4TS+B
/BYRBhRLO8rOwjyRACcj7D6UmyKaoDt52KE5TRE6OB9RKC+WhE7hWZkomz4wUj13
SFjgjkSySzowbGunxcTYwbDceUmjRGWnEwXGF7DAP5qQheM6aoTzJWRc89f2bfdh
bBHeikwDQUXtTqtR/KMt5Ez6Z+g+IwSnafBYnoDiE9vtBdV00XrOtOPGWBZnwajf
8zKBwbcYSdvXjjYTs4pszid2OvCDZ1nFp2tR5fWZ4ZdR6B0xFK3aVDh39CFVeBU2
GGkOHofV2POPSKy+SsyDOMI9rnHXjZ5g6GX3aWsPwLJ+ysCsgx+5Zr8ocJlwm/5c
+f+dpXHCe8+Gp0Ud7AYhTnA9yADZq/38YNRlkUD0thnEW4ci0uzHwIV6j2juXSGq
dfxxhujhSkPsNbcoon8TYJbNjjy5mGefk4H9yta6Y9mpMaeWXPMzffiWOKiX9ssK
gNCuEHIK4GxWE7EWNnQxPC+uxrrTO7Z8/bhA8MQJDhBJ+7EZ8C23LNTci2pcjQWj
ydCRzJTD8wbMYH+VZ64BAXLkgK/b2cV4MTc060O76XD9hU46ZgKgOKSnz1oXFh0Y
GYfyaqljXgM6DOuEe2EW0ZDu9e4I06Uof1CkaGEhu2eb69h//y/XVptCU4sI+JPT
qTlSqArOnygBSxFESUrrPehp3HxQWN7c4gHchUUZjC/eP3r8E+KFn8HUpumT6X4M
pJiCaK/jlMcfevN6WQz4BNiu5Fy1AgXg7yD/fqg6/gJTpCChFMWmKIuvYTxrqW8C
/WKuIlMbN5Mq07kV6nibCJ2euWRgy0QaNxXJ/6rcvYC9T93j5586Vnv9j1hSIGAj
T8VlXQdWBbEWRx02fXOHLDWxKXlxn4rG4VlCQeytHW+i2M0Vp6wCHA5ZMphWZjfW
zFjOc56RWb131qoy9gmjmbYuIf3+OnNWZGhmORMZD0qJh3pLQi5LBYe7FSYDX6ZS
8cgggfKGAPjH3ufK8472N8FxlXViPnW9yqOJJ0O7HmKZOPGIb3E1bWDCqgXCbUYm
/ZoU3KYY77OkabkjsGAaMWHqoQO1FXsZjb5+eh4QLA/gDqhtj1EG/uZTCxsK+gB1
yaVOUl1oxaPW6pErf28tvhPQ7Ssi3jf/Ty6uiwLdbIzb0+Uo4c8vmRWEoeyMShkE
S1mECZAD8zYmu0UMPLrspvYyLCbWIfzQ3G1+Yo5JMNYN4ebGpKfvqI2IzyfS4toQ
g/0Sazr0aBWQPpVEULuNoFlEl/N6v8dAo0jCVDSO+J1e/Lgiq0AU/ohWAwN615L7
yEhl68nKavuiaEZJGX2kVijT6KhSnySxiGicLHDtY8WkoP7Mu17RIzne7BYBQG6U
VG+X5JCYqYfMwqHAwxq0KAEc1uevQvITfbcLLKfm6KBHErsM6ZgS+XueeNR8X9Fq
XPHHZxYTsLpfF8CaPculsd0TPRAI/dn45+hOGxBm3hxG9xOG01EJyleCnTyOCKw/
usFHuJFZnFT+KztIfQDDnd6w5/d+g9C3ei2GhScD6ozTDXuBKciDap06YVS0O5IM
oABy7psKZAdXNevIi1W1eSG7JSXWdcMkV63nbvuN+w5iLiTVWEPBN7u7cFaZFzeG
mun7sBiLuewwhmwHAKxdxyvKdpGEuDmnnvRunimJWIh37I8AbMje7FxMpIDtfgyU
QWVPqEDGgYqaN6fhb3dKLC8wP31diUGApGq/L5j9azOG2k1qNNZmjvYVi9fOphTN
1jXN3R0GTkT7P+mkJOX3Edsk8OjBuKEefzGpGTBHPLVEn80pshIEIjfIfJQuAzti
8+vE3CC0OpMvFsg4H8khGLz25onOzOywWow1Jb2uvfLutE5O9Kt2AOlmc8f1klA1
g/GgE1c/aGUNw/wZq9bdi3dMivGBeHW368DP46rxyVY7t+6h/yMu+xD2JGIbOdDY
PwbEqep6rzoCnQLdsO9Z925O+nlqSWyHXbCqKvrmNpcRPLWMiBqMX+7EC76xrZJb
kmzvcn+5U5ae/BpBM8qmdNRA4KhK/75kIx/Hwd6ib56IWqGz19wxZL/BPsynZa8X
5IcbzR8IUbG/U43sEOHUdN2T9U1Y+rJNXxnnCNKbW+FkTBkF5TxHgbCL5o1MNkpI
PInZOmbOdk1GO/ljuy4upUJs/Q8oJW4EUF+4MU067RCpent45MoERURU4eUiadbA
/vuUAtZ9JdbKtpGiFpRwVOq4hUfRPNYpp6fCmlkwGnVbAK8JIInlFx4qenaCeixk
hx6gS0XnsyOljturP/KnIRVOVoAkguawVJ8Z0gd7/JB2I7XRquT16un2g1y5lQKS
/5w1jPwq3741EPihRYdyFlMidrxxFKUKmwdbRKGDikaxNPsSNe0giMLq/gN1OXHC
c2VT7hGgbzbxgNg5UiePlyqmL4uj5F2+ZTi4WnwPJkhe+j4VMVBhy5WRfp81588q
/z74q/OEK/bfiLdsxi+NYNsoZvmZlp8nENPrvsxF7mg5IRSVxvexbvKWgsRZwLhI
OjdmIBBv8bthnyYYwERXG0MazT9qkVhFGdMrEk/9SnUrG90alahCL4fqx0U680nV
xoTJFwdL2TNwRTy2MmT05/XlZMI6ik+ItpI4RDJ9P3flDLJNPjXutaiXrU7vvF6C
xobac6w145z3lFu9UATOyan8OAyz60wmQ51mGt9yG/Ig8OAdX3df6qUSZI6Im7Bq
ZUjc9+M+TJEVe+Fx/jCzGGATbej4fLynMb4zrK1KZ54fNanOE4iRnvjjxB3231Dd
jLAWdLIz48WHYv+I+u29IG8Ez9Mp8+kY6JSzBQ7lmAKJMAapgNeI0PkZnjjwzIco
z5qj5X6cTp6vamd2Tu4K+I1PFPL4RkidrddpNtS5Fd8dLJ2rsYu/5h+iUMx3oiPT
e+iycO3GJyXEEe6UmtpgMGI6+O0D6HmsxKdE4ZXrZUzIoTWVOmHO96vxbVnb2rFs
nJpw+OfCI0xDFOS16xRKTtJn6CYIInXxxbfT8XziXa+UdWm/gXHMhPoOlQvagIKX
5fdQUaLwzjdrbE4ql/e+/bVa6aVZewWXD3sb7uI2tFHgLpjvWyi5mt7upy+svV/u
UpCgDsLguvqn+fqfVV5t40li9pxV2bhFFzxUcR10HZ5oDb6lIzE7yy+3VozGIEhS
7oluXRJLisd2T5Iw8xjAevuHl/LC6WM6+5N9d8BgStpl/d7E7YzsqdgMv35At39k
gi9h0pzsOVXF1Gszv471BvxZHbwwgp2v3LunjlbF84T7NduEubD52xZgekgzuo2I
OB/dK+eFWlAFViqGBF9SfgnqHremiy1G2RiDFFbs0RlMyWcEotEqLmG0Ppf+6NTI
90uQfukFLEml2ymoENHYHUsybHai3QaWbLNN7+1PdVgvZ7c15lSbQQ4YLVfM83Cj
WXxd/oG85Xpe5n3kGe0eEoeXPiF1M6CK+dzgQ5OU+CGzRdLob8WawjkCq2DVpSeS
dGizVRV1k/jIVJUJ9b3Xk58WzsMocpS5YQaQfmD6sXpjSrW6wnTTb4I1XjxUEmMq
QqU6ENilMMbw6rpIqXRyfQU4XiF5xETminPgjTqdDMhV3BEIS4uG408Tji2K1Y9e
8ifrxoQvQzni3cRlbulsy7YunC5sWxbUmDxxQk+Lbd+s/t04pSR9zDatsLCfMFWz
KUINOoaTtOD4VWxtzGprMV7zUc0ugbatHcqU/wTaIWuAM5465fRI4vrCUUI2kjxy
/3bThMDhvrE4l9yyBGM3CT6zei9p8rQtyxgY8aZA0udukob6giDNQDnRFXXLdTK9
z57t1iOmS1jXhZK4tAqgcNEwz43ohYg5SZztUIw4DwrCdmOjj+WiQeQnk05AhUXP
b+ja1nROB4wJRKjoof0sLn29sGeX7d2KFTpjqAT7AaHEFX1MvmmJ5JwJe3cfUkPr
aVoqjYAfopx0Js9VWm+XWmcJBv25I3hRNaX5+TfSX4WxZonC+oIw9oDHvT0eZeyC
SqYv3pd8hW01L+2hU6lHwgPqUVCQBR8scKZDjK/+ylXBS4lmf1qPrHYMfcfCwgyK
1hfeDMHHBQq0r+e2kkLLP6yd1BW3bLdCIAUAudu288Pu1UPAwxrBR/ti2gQxYn88
gtfAWZEK7Bj3nH/mAPzGJq6/NhcA/uZtteCH9fijmcon8QNNKvzGWlG6b1+7mpQH
01KatLzvsKBV9V/bm8lsHF4r4fVK0nX+Jpe15rUODWJ29KTbDZLUwo4lhNIAHM+z
8Ks7SbotmLCc9X7mrssd+wj2QZVkAOw0tC1hqVr2bra+J7qGFdgd0Tnog4gH5bSR
fcixDendpTyJhMJH00hPTunRrYaXL+2CFpqmLOZaUCdRG7iNEyV1SWcRDpG1YBh9
uv+jYHF7JBgpd8L5XnWBJ82Vz45DDCdE150lDnRxAj9X8rwQnIvpHnTMdkJmjIQ2
bh+CUUl/6Ev+l+jDS5zPiayztpDGzJCV2U7r+Zg0OlsTRXiTRdIkpikLYKO7Mk46
73A7oXx7O41zm8ofK60scvGuxx7xQY83rm6/T0SxCSqnrqd7lIi2MhSCWRAxkcXQ
AGPc9PR5W5TO3xTiFzav6EVRqZCG64iAuVmlBw5HMdZ7jLDyBT3UJaye+5YNmlTi
sH9gvcqF3CWCnFGLWVzJag++NKcpAZt2llPTQqe64ZlqSN5g9k1SQ2dk7QzoAWhk
eGqkBo9Jp2Wvo/z0TC+Gia+MUmRAW6Vyut0081DzZBDlFkH8LufgH9LGl9RdKesH
QiAL79aTDU/zHBg1NWb/BPYyk/dA5uNXvdOt1Y3NTP1GdlgOzbBxBy3BUpqDQFh1
4X/mHJ6e4K1Att39CFN+DUoo+sIoeN2bty7WTviZ3RIGD3LlS8DBhE1xALREOFdB
52DKw6CjjrB06GuDkz40YEyfijiFlhUlkylGzkV2LS87WzUqiQ0kepd5HwSpJxOA
5UsKF6tWtHqb1EgC0xlsgOlYP6rESoZX/hq4puzglIq8zClFN6wfA7brYWEWPFIK
949glZsvEu566ZfD7urQG4NCU2FlPksNcKq3IKSoaogK+iHz1yD/+75n+50F3QRd
GeFhbRPQ8iiIHNGUT63i9Nb44tzrHKexQF+PXiMZFkg9fXndbiv6jVoUoIOxpyCZ
qM5XIHwDeypKiwnYlA/SMu5+5zKmekfBryDtomxv05NZ+TpQYUtZsHoqrWe6txiL
7lgdeA6d7wqhFl8eT2AQrE3OmEm0Re4USN7F8fcWS0OvQd/ylTG7zzqkk84W8/oz
zWZl8bYop896TCg+tXgAqs2qrH2U7PvvumS5ZzRjNcwYmd4bv+9juekVq9ZPLKoV
Vc+RttMHuemIHM8SXIRaSkvbryhwpdbNzD12nXrzxcTY6qa+7RFpuOEJDcu+fZcO
ibyjtUnR6U5/dmdtBPClAz2q8C4bN8VwS/cPGcUVwRelGtyY4sfk2Cxsz1j4ykmt
eNlIO3EyP0X4ElOENDKfvjE/3huEp65X7iKLKr9gr3G9B/o0CeI64ccGQ1z0LDNT
dfLlcAv/qSjVWxh8QBmu+Eb2uva/2L3YVqWrQH2A1s0lxjzyVlLnA+KN+QJ7NdVx
J4i13iLMojPOTqETitV+wIT0JzVvNID+kWA8hTqY7aijN65SUHzqteNCxupSn7DK
Nqh+sqZbrOQfKTP9aHJbT4U1K1kJX99nkkZHBMonw8Uph8lVzgJ6o5joD2YDutcA
9iP1RFkc2mdOeAzhZgtHGvVh8UfBYBHbSXjmnSymMFS1rXKgM9xjcXaZZ1Lc3IpI
5H3DJcHGaVP7KYhpnEEUguOYbtffDyD8Po8ukUtjS+juUuSVqFUGlykUWNnP9Asp
CTa6R1atZkUWIUlI4SIZo3Ip5+eIXHYy4VxfINkVFQfC+0V/AD3mVkaXJZqjwnje
/GMt9vFeUfql9slahyXNkwCNCxiRSZQQ0mgE/NORMqyA7UifHB0hL5Ki7I1OOZ/t
ekAvau/Gc+a7cYs7cBOScLWvIJWhxlmsgM08hY+KdtcPAdi2mcBIhrOQc0W7Nx6G
FG+exCgMbYBNyfTquf9KSISj0Zc4PLoRHJRIMzrNc7s8dV1zK3SvC1CI4h2SWMUM
ET/HO4pm/4QPVm0EpTZ4SPhSU5YLm867eBIXC9SKtyXYe+mVa4rQ9qO1TwtXfto0
vTRTkWdQ8ZD/pMNMm1uDe9w1freG+SQsQSuUhsTrEAbf55LibKFNahYST0sA2oX3
jH2WwkM90eXmDNGQ0y1exvCdF2TzXmYRa8eXebCseZg39pfSbd746v6cpNnmDy8h
0NQVsekaxTbFymCuwLTerMMzuNAr0+A9d6GQvMjWPzD0m6HDJoYENZSDHioq4XlK
Bc0ShH0Mpp2R50hrONKnGl3TGd2FAAK/hekNvK+4OLD1zZ0PBtRwiSEjL59CFxJ4
dr1U0EtA/YpbT+yz7zoq7cKyQ1Iex5yShEQsbiLJrNPd1GYyRaBQQxoj6qHJ1f0W
wggImu+oSZ/QnuHwN/4tBxGpQ5LjZbangvCHrHAdetTu2WD2V8chcui82eVqVTnc
Sb+n+rSS41ProlartK/CvCxlTyb6tWN7RJm+0FqsFaSTiRPWcRFFSKKKS9LImgWu
h5SDDffmYo+h79YClCJHa+OdF+Dv1PMwWBbacMZgLSRXRyS9VV/hzpHWWioZe8iY
SKoSRIpUcjQzFrn2UIrYetaIqHfRm5fwH4/zhCCOGouJzK3J4Z8AQlevuAOUfKXQ
zMdKdTDqDNiQ6ShRMWP6zs77H8/RbsFdM0YqBNZrzkzOzq9vyoux+36WyKEyj6IZ
HTL9N+tu0RZdurhFxfhi1UrzbAH8faaSh+Tuh3Gg2fzkIFAXj14BJJyivLGozuOm
9eeYpEqJSND52roWmFHk5Nk599eVT11n4fxwX4nxY7ccDoAm+kh3dT2L9OIMgNiY
O21uw2slCuHcPQsjqwdrTsvaEIJFVKFnVCB6FLJAzgx0d2VCC+OCizG2Ztc6FsYn
mW3bp3GQFcwgg2U8kMS4I/Ireb1FeDIs0h/FauZbB04sbIF8MDQNIHBut1I8iGyc
LjygjYM3lwFO4xk9y3WwEcY9Q4Gz0PVvDiGCEqp4HhZKDhSf6anWM8r9KngXl0ap
Dpf+IrpdFloN4fGCVFI1jbRWXdEtCj7xHPElmbRYbdwy68ygoG9wdZBUR+tSpa6o
vvMnt+YCbazwmVbTXBMit+rofsDtx7PNvjQH2I8u60X+yByfQDrQFUiOG7MdTMEO
wQwXFWJuR34IYKXcU6WgbtqZc7SgkEE73R7hT73gjLfxQGu6zG2iMFNViNwtGXYn
Svft+VRWifgNDlC9JHcBQGr+vqdM5JDTyXUifEqKa8SLKRlmNLkelc3/SX6nlAUd
k2O3aXjKqXWyR1lplCKgpil+KNKWcCm8rlD+Tnt+DHBgHNJZT8SK+sBfZi9ZEp7Q
RDHC0SWOlfDKiY0W6YhdrJNKkui/gxkqWet5F1vkffTrNR60xK+4ZJXkQkNmL6cU
cyuXIbtlobinDNF9Nl7h6JCCjDROrcijGQGnBlV6mthTy+63nweR0GaAcDuJxIqm
0Q6XwPGDDLSXTRX9cXN5DoZ1JOXw7IWTj84VXXEHFwqssKb5UvihsAO7ifBJVN+7
ZVwQ5KJJUGN+NkrMsonT1HKzi3o9LFvaXwM0VZfIfCTN0tOaIQGM4bTGea+k4hz8
1iJp6t4rWa8NI5imDRHj46ZaiQPaEUBJrVF1Bq5bON1Wk6vB/3M3R86nc52Ufeq5
/+zu121RDfFhJNwbXI8HwX1nVYiheCnhSzLCzCGJ9dFMQGmBwFzthm8R8PRhE4rU
MhnQkLSkAQSoMbdu5aCMdEUL7i8Xu5GQmcHLymSsKWxM7hnX2wBSKX6vqJzk37cp
YEjq/7rPeLEzh8ilzVVaSYaYh2lIsVZiiJ/ZeSHgeRvN72qWtBzoVIQ98txD3Gt1
j4aaEXQfWg1qAuukcYGU8Iw3SmRM66Gkef0iiwqEvhk1xCQdfUnTHg9+o5InXz0I
UjO9L6Y93An8CsstRzJDrR1/+j49coQlwmlsIsVHpw/63dOenQM6eTEP1MKvoveJ
RtwHVU5wF7CyfEqpcJ7V8kIlBAB0qlxiN1fRppMhUqUL1iUsIur2c0t/UitJkhzx
Zi4fxnmRKNAs9qc8Tbh0cuRFKBxT3FTPaminIlcVsHirbTSwxs1S1XRFLuore46X
M4lsuKpYOv8ONo7zqIlz7Fy6xFCAD1J/r0dBdLjRdyHFL72vvbRsP5vIrrj3kNQD
YfTz5rB3BWs64fJv4vMaBD6AWR6ozZXtYOkJ6Kd6EylOjXYkXUuHfd/UqWf2BepD
4URoErqmlHOqmtoMQwiQJIjmCUtV/3HFKGxwDZjYXv/f0ZH4rrEmeauUgdcX9U1N
I85eTCb7vQXtcq/FoVicX+gmTdmw5g6ehf/AV3qh3GEfrj8pK5YtdnkHVhycCPOF
hHWqVGG1iFFqpPrdrIOQhPbYwwAFihVZ774XRNMrDF1gkuZcj+v3zZAI0xwEJe0Q
rVVBsQ7Kw9oCzTcPE/HZCGuLAYim81xQTEyk26nd1b/gTAGpnfWGBkfi3s7TaSbP
4CZqfoIb1Quxrc9occcFiuLjPgQtIZr+v/G8358gB0Lh0RKsF9KFzMuzLepJtsZ1
X5wfdN/B6hyws4xh6kOoRve1np8l3v3Zk3SCPX7vRgff/wf5tXAc84vKYqOVx/1Z
Cw15tAK4o6yTGM9OGXx1JtNnfrgg52kgsftlPDh9qosdFoKqoK9chPsfaI5T46pz
MBLhm4cAEBRJBALBp3Y4xgKQj+COOOrN4Q7K6rF0eNtQfzchzJypt68YGQyz+i4v
K9FEQ/5Vhc/rJpq0Ou/2brnv7XPQ5JezO9piOXIYmtkibz2GTr22zqjN1p319H1G
7Dt7YESN/uSQuJ06C7B6PlcZGzMwuKamCD3R9uPvFR8m2joQvjO6dziGVHvDC7/s
2+tifujab4wc9xJxvAyH1yuy5an3dZrUFc7akXEcTbHMKY8nSwgPtM16HFiGAu3A
Uj4jVQ9fQEHun8nmc7Pvv0pU6Kwxxo8/z1kGDAWX/Oldm3xVfeQ88bLPYhUcgHZl
Yh1Y5SE2MxzYz2CE/yz/5k8jmSerYLUEkt8k0dKK6QqnmbsY77PtDBX1XAyVUYzm
KliQHO9opL96lbGusaXolW/ViXsT4AVyF7cbY8skIQtKNFfKyBHeaiW+lTL8+Uvk
7hFEuN26KBwYuCkH/z69Nd4mmN/CW1bk8DU5CgmE6yb7iN3DX+ip62JGaQsnWnDd
qLY3BSNBWUodskyZ1lCcBLIewmq9Sx5fmflG67WBe39SIzAdvp5Y7sV6PYAULaPS
RUshMzPzI0HI52FDaLmT8L7GX/MviIVbMSbgAX6Xw/KSAQVIseoht67xAoKJWv1Q
URuPNDVdqM0Wd/AJquiyS/MWWa6+1tCOenQjuJpVGSrT/sWHKl/gNwd4HlAnNQxs
YxeESkuIVMsQp4oxEFD6gKw1n6DZ6RNn5x8zfOBG6lClmEdUvXFBsh/WjjtbzSvI
z9+AmDbMPFph0RhBJF9VftJviGV6gRUpGZGwRPacbT3rIM7PBtGa4GN+5GgSWMex
i9CeGH7lDyQWpo9sYznrjo52ywbaVLnLqZIPaT2GJ4ixN5ZAml+qnbMRg/sCAvb3
RsJghXvGvIe6qCK/U0VA9wNsuyc6tPKC3I5OAGozgCg5ppYCgc1f/CdjNeT1dw9h
A3s9mxo45avXhvdMDS8ow9ivS9i3OHPfk/JhR9N37LrdxPFzJcA9UrKlOlsRoBJs
Ip8KL/ZPn2ytOugg/4IRJ42eLg3QX8KQlOzWFldzPKMxx/uiAKgfok0fVOyjk8V5
5iyAso1jgazwKR1p02jUnJbZA7Z1IqRKirGSdc85CKQEuaWOcHcQjFutiRZ47UJV
Y8fyRPi2r2UNHuqEkbHFspgOzRAxgyBCn+WYWzajy7kP5TxSILY3QnjwSLpRKVjW
qTFCEdf+5BAOtp2ECVSsdsuPSFcweC0915BlWkELSLPmVyX0t/fno712ehs53UiA
OJ8KayVptqz0JtYrRMSW32CrnEMkT+4kwnrJHOoI/RJGgVH0y+RWlv+ANnQLKzlk
lZnm4welo+T+cmRXrAnCmywA1mJyIjJb6AedWlsvSkiPvZfAeqaVm4jMt9YYEfcA
opwuimkFE8RSLS8ZmXyaOX3zoTb5H8uAZmBPbdOvKDTswdhi5ej1qnJEM5fbJ0F/
IStOOqqGTTScPQdaAS1ZQoRKHcxxkY/Qav/K7ojVCe1bWa11NTYKvuHWsJn0Wdy4
kj9aTIvhS7mxBxorBC5VGum0ztJDQcigf4r1rXynbR+iWtqYmDvJfOKvQNpAPrMA
+ugyVSmz/ZjezwN8B8xjGaBXG4IS8ODq8CheogsiPQMxDCR27dzve8Ml1AoBjm46
2vOxa7Wj3Lbf7t6ReckJO8GFsatthmKuk2iixCMRFWQJq57jsMo/MedXA+B33MZs
hk6QpReFOYsPr/4D2c2R7QKI26vvalq4iWcnBkjc7uWd1viyXarCDe9inzXncHl8
dj/LzZ5pJzVNngQKV3Jue9jgQMB7CG0H1HqSW2h574tp+PJF0Vqpv8hiTSUwZpUw
Rl/9K6y18hNITusnyAjMi0+9wCKZJxn1HnBRbP1SVeWNG/B6lJbElkqHlMe2Oi6t
XC+yfitCiXWsTb2goeP81M7dmD3PH65A1/TuJ7ejlO34cwdb856svFWX7I/VI8pv
o0n9Bs49kNtk4pruSdgk4Z9U6TAtkzaC26/7QC3I5r6E4ZxVGSsn/swthfJB7oqa
CbjbibkiJp3SfVHDI3mIbJ9ZA0zSd7JgEmVF3LIaItbNuk4VCu7p9xzLhpffDGnY
SP8gcMK9E5xJjaar1e66UbZn1+u0VB5Suva/60wTz82U922bpZAzxoxrD4fC4Xj9
D/iSCX7QFRcBP8GXtRXqLe5oi5BYHzwnHM/Vc++8oaZnhcdx+9UM9hr3RUBQzFbt
Z7X3pzqO88vRu5aOc3/vbChOc3mKUwkwd9aja/DIGtnpTIOdhebnW9GbknmjzA28
TNbv/NznLABaB7i8wBZYjSP6StW/cQqxpYW+3w32uYCsC++kPTOfWl4Vkyaq1sKm
lT3gT/POEt9XTw3jSfGW+BH//lwolzEEcD6QfAJEcHcW9ZHsqFIAs4qRO8VY2QCL
YY2SJFgUIUh144sABa6yZVt3mIlFe0jhRAZqPg7QLaJAGAyqYr1UY8xNxAchLpz4
yD/vZP4ta/E7KkReesupKo/7wWnNXT57sr8P6GfoiXUwfbNAg/YiroQlb0DPsu4j
x2p5TIrjah5lEuWsCTXDpl4GTaSH3giMhqfVjiVvfkxIi8xctxT8vOzzee+/EkDL
7xtuefpyjpUltDR+RkAxicqjQswi6AqmMuUqUCdYXZNFLembEwZsVwew1a+kq/2M
27cGUQwrTpRk9k73LDTJfo8S4YqmsLWs3HvzdPUPIZFDe3t0/+r9/f6WPVa57ubE
n23nHpwm812h1OTnOIOrt5FaaVZkE6XxL7l9CGQ7j4FLxU42YupbH6r6AEzgSeNW
5iXMWCDHIAxF4kUwUb7IcaRkHLrL/Lnow9VeYOqyOKPAD9A85qVqo2iAPafq08JE
sfTpmRkvnH1tgRbOjNI5yJqWZOw4hqhbrFtmG/4YOev1jCCs23v+GZGBUgJL+ffc
YUzdrTN4ae0H3a1+L5jKoR9HJEknoGdrwsVqXvW7jUKaKseATMV1o6WYr/CYq7tl
uuWCeknHdC6WweamhipB9dn61dn6bjmuv1S0QqSThr1jUjAx3AimmvTJMOLmyes7
a7En9ETjmFvlg+qjeyKfPtkUYjrfCvw7EZQCcIKIwstMXMTcGGGkP7uuGxfoZTGP
9TmfLMD9WkiJqSC1fPGnSVJ4ENK6Cq27Blj2cxSfOfGlOFojsGmh/h6jQF/IyGjH
mn6TtkhfWmf2YhEeym2LHIVLLwdsOxWA8GAKmALrXljUJUEc19TItQskvlUTcqjr
ycEgQbPGZb1EQ6sNl+dVBfJ8ZwXysbOJtQXM0VanZO1MgATqUV4ZKCAtxHSDOA0J
tfYEbGkkIBpEWoMDkftyKf4h4X21q7EwGo5zQGrzaUDzKo3o3Im9L5lPkkAkSfvJ
kpI22yUTa3cHOo6yugO1pFTJ5vDSIbb00ic4eLrs87ZFdYqafk8/heVp9SjZYz/y
xUwOcLCEwe4n7bbOwoZ+5XAgWJc095UQoJP6K/NFVevr4S1P8c64cgtIZceN9IjD
/IwE8ZplLVRMZVadP6sHsqf+8DQt9rxha3vmWP0ZybIwwsY3N+dGnFpUAngzvI5c
7zeC+o79TV//TBKfgV3Am6hbFyifNt/5OFUhfdVXr+aDEDB10a0DGza+gkzqyJIr
4aLseFaEcoq0qcdY8RESaA/A1ehaaKKeqW9HqAKjTeLm7xow8/0nfa+k2vOkEfmI
VNbcuFH/TI0+iPq5mSsr81Mv/QzUbXsjwJ/K5zByJLv9JGo2+8DgWyTp80kQKQwh
dfYqlve8FWimMuu7aRO6Dko018GBs9MgLVIGBAoOuSHzNYHbXKbjYl2s5v3w+Gk7
VJDpqp8+2NL82XErrZSKmSNazOMU93Du5uzAMl1l2uw3/2uyeODTBuoOZJ42eAUU
De0zQGrwsXYHG6cADWz/mQe6Q1Vyg/2xQEE7nOtMSKxT7YRveB5F6BAsh1DZzv+F
3IKKSCbywr52vYFQsyhriVVmMs/jnYUnpe20EuNwWkbSuXvvbvXx4SuH5ecyT5/Q
84KmXrS5NmhQTxecry/hectDCSxNOMQkgf3J0LnZ+IDI2MuY9FnohHaURYxur8oc
ZWb0NzfkpvCXa6rrQ1o9SvcryPU+tXEWJFH1LsXDBgOF7arQMAVG96FMXMqM7Vi6
RuY9EGyIYjsho7sZ8dz5N4a0x5CGCSSm1vk5gX/At+j8rUyThItEIjfUeqpgbSPS
p6z2Kc5ooH+0Tt3qrmkNOC+zI0KgZbU/aFh2ahG9lu9yRj0hlELnQwLbAOPvSejl
jAyBTXkrc7q7bm+y8k3V0BLJecmMSfc9kRv4/BUst0tiTTJ806Jm74bNfJuV3IK1
TBP9+/GtzS9l5Y0lwvjSMtgu6DAGsrQTGHXMAaWzeuXVB0+ApIIKiOkwsJ/X7RCv
GZKfkaSoOMsVQY3IYaG9KAx7AMpFda6DemTLrRBgR47A/Gw9FmEaW6fq8UNaGEyh
pP/shjVUmSFNhmn9leYm5mhWwqlTFBXRhuaHire3zhFaDD2/+Yu0YmOBzs0WUPvk
WLwZxkwydCgrrRNXlOKDgkAtAt1UWxEcQncBlfLuG+XeBjB7OEJvf64RHe/SjmTk
xdhwDTJj4/gJga22VHOcn8kA720XwrWHsQgeAHtilNCY8KI2lJnutZ0T6/3LJbbV
S6/1eFjMfVfG+jnj0GZkrhFX3tkHwPt49dHL59x1Or9zbVyZy2C0qPh2attc8POm
dVYvyoi1LSVyV2dWJDsq0kdF3SfUtK5oB3jS4oVbqG4q/n78WJsBLqzGmSngb1A3
dFHecmTNrq6gO76wQwtEA3HMBww9EvcgBvit1ziLQgcFJuG9TQQUIbQnch/VFE5k
GigIJCeYnZ6AokJujkREevQQfzgJ6YYpRsXKrRos8Du8+GBgFNI0Fo49IWm3Gkle
XsBNgp93X4asAhNKjs3P+DE4Ll3onWTndR/4GiG2j8IcUcdXjU4EPD5UCa2AmqMM
yBvf8Ez9u4qsQQOqLqUq+3AQnXcB8vdE8qNYY4MuVPdcjodDU7k3yryelXcLkAPG
HMMg0G9srFh2uqhtlUE2SKoG40lGqNrUvz7ocQhinUyC2/FlRY1NJTTgM5iS6TfJ
IKlOsp75L8jj+ziuUwH3yBKDmJFgyVp9XyRsJppgLDNnhSZJxqbEIUwoo2n2y/Qf
nEwOh2wVSb2ilzla4O1Vr02TngBRFGVWCrAW2NRYktzIZYvxu0UT6VQ3JiL5CzKp
5C+OJm6oS4xfue9tpOAqKGIvmd4KQ2SbHtUpcmpxMkdX/glrpIQhTAyCaMWXWRjD
qxKHzzw5MKvhpehCdCYLishMWatPrlDYk0HNbNtQePLtOx4w4iMqALm2MsVt8qCB
4ufERQCDs4fQTM/DsTPDT/nm1IrW47ZkCfjsUprFvakyTVr59HMovb/Gq7RL0WJa
PKaphSbnf3RpMe9RL3LKEjrrkHzgYTI9GHXDIi1wZrzn9+bDJTeCmREqj36UJj6f
O63W8No/SCYV+kg00aUUTliGlY4Y9KFpIB1wOs3Zm3UkH5h7B/nY2CnwIxbZabh2
B67pbkGcbsJDFThovs2ZPn1dCA7+jKsOPwtzr7iPsxn622oSp5n9UWq2cc7mlBX/
eW3ifoQP6fnNVHJwqT5PnjCFwszLq+g7yr+Jm8hrsNMk2SILN6yW3NgrqkCNq3cp
1E+pFN8SpxZXK4RsyQBfFED+Kn07FiPeCN3QFqw0Af5eLVY/eSYerxY7/QlXRgCz
SUgw9E0beDkwjUizxKWwTY9dxRSodoZa7Z3AcSYccnerwiuUqq/Ru8r/HoJ9IUs+
TYYlmSva/sBN0KDhJrI4/CQpyKNptZaTCE+9RbRCi/vQ08umJF3rvtJrxlu4vvQQ
CRt9xLfoCVajxT3mt5kfC4hf8Go5XaDVxXo70Jld8yZuaDd5yIvWmFyqkMNHrPtm
x3dHMrlvxbGsUH0ic1bRwuCkPZTnqn4hJf+Z7nmsMgK964zlVaUkqZulUSw9pgPY
KijmVhEyOX2nB6gyypkgAbzNF1izDGWBwcCoFd1ohkPn129pqIr9hS3wvU6ka9ZA
ZdJ9IVVBNzwIgVg4D3dAYMqzrXquFfKBpJ4h8E6ZCBBoiopMDUwPkqkTgUmrrwXB
CSkmiT3huwRLWjQ1SAm4/Tls0owFEZNDYE5UJ9CDwFhR9lxmF6WANjbo532Rh+gM
2QG9qhft+HV8R36jJuTRcKbiVOSlxDHz1oskpw7YhxpTXqd/yWEMLafwhkgF8Xdb
cBuAj1o96jbzhANd2sKkz0O5vNizAnwp7l0rSAabdqWGY/722t09WNzl5im9wXAG
IGZdpFQtdOsiMMePgH21uhW520W1bxVpyWT5g4FVDAaLptoEWYV1GpP042ZuRqW1
2U8131XvczbG5kDtOLIaye+3Xo0CB59BYn6HlWwCnwz7zz6vUQe320sl3RMtG/7O
bjkFrSme1Nh8B3jdsZDrRxwLG1Kmcqn4+vlBG0380lr3jfuw9Ym+WDJIxLKcP0W0
d5Kj/tEYfhY96yj97fBrozN3L7V6HoK9o7HM6UbHj0MerzppykL0l7TSW+6gSlns
DnD7Ov14Nsj6hG/LM6rp1fURa5MHquMy1GV5DMvts0sXjor5SDQ04Vzgo3ndgqGl
dYu6kTqXxDNu38v2bIJYtJaY3+k85mDJ/S0Vri2tbH2AALQu8zKjnTukXW+rkqo1
7iSKHBzUD2JXoa/6QydwI1n7tbpTlKk+rnB7aGV8GEeDpi3uhwBYzDlx+FMCWTcw
b73/1y+TZAYyliuiMNGhIt9kYCu7u1lGzRnbYzru4SRlvbd35Yc2pNJF6KzRNUwf
qyH5K7xjSsI47Ber0iAM7lwOuJ8zISDV7DVp3JzTULReS1kYzVr0oKX/EtP/Fkb6
t2GIcpBtZNv8/H4WcbLFF9kAUVx3tHspmuIaEl6QObYasgzfSFpcaJHEZ1g1brgV
LLqXDQ9pMKSZbDL+3ak10mEp18sQ2d3V/NexbweW/2/OFcOjV4YP1CJ7R3wZXZvn
eZRE7cW3L5LoMS21t8+T8Le2JZ0C9rcwMdiCHiQBGBJLgF/AtGNo9k0v5Q93egah
4kUbSGV32CJr4swmHRlAzo7lb3zHw/xrCvwe9Tbt5XgMPGN3Dk0yRNj0+09bB1Ba
SuVKDbWcBqkZ0KeeHKX8UhmtaPYW9/SD3v8TX9oJU/hlS/Wpbly5nzwDq+geti9C
UPSY+2P+SlmbNbzRnWv+4zSad2sZ5rgQpdyBiaJ9leboZXqoOq4eSsWtR6yMN/JI
HhYf6XDm4Zke1rIkgdQOpCfhqW/NVvT7tcSNzPj21tl8GCtIGYWsRkCyO83LtHM6
1/HOC5bTUI5F9QTnA2y5zhrfb4Cuc6ePas3A1dI/KLRdmfmsSizCKM1zWAKbgudF
xR+esleH9jpWdQcVZLsA/MlkFcZLhkpuwIRnV83SXsbBL9UHqhHeT1GV3PrOoZlP
m2YZiJS7LqOBVUUkl5b85wfeBbnr8xcrqmVUSsuv4FFKg0dXnw9t3zfXHtmLrOAm
gMS5tcf2i9WepY4CSxFrzWrw6WgnQoGyOTUpTUBDnAwK/dnPzkBKK/wUdZCM1nKE
haghHlP78ZiQ0qYndRuhSpREnaNGL1/AXqV2MogXCJg4mPLbVlIFPVWswLONgFBG
8Dygk+WwDsD367qVdTjvLVFxLyVENIP8okK9tZS+j5Pd35nr7Euz8X3xOKAVQ3ND
/hsJ+CvixiPkp2vEuewvjtvrXYKiSkzuDi7eVwZqglBWwOJhPxPuHwZrXY9Qw5mR
DWpTScmhMFgcchiFSpH0/Jl7qWGbkkxTnIcnlB+262LKpGMV5aGEiSzNziTrEySE
ezDqhmBVwwQWLPaN3YSA28KXCpIt+q5TvI29WBYi3NXT5X2xnBV3JuvivzMNv5My
QTsaFhvW347jzS3Hq/bkulaIa8qOQaPLALpTNUpB2ZtBm2X+Fd2wsggTvfU+u6MV
UzWFLbmg1eJ59L6bgJ4HI1LFvQWujGZwj8AXoXtrMnujc/sfatV2kZwE0IDxZK8U
i4iXTysPeUlzvvYVljjT8FbdmHzO7wcBPseWt33+BjtDW39p+2b3BOr9NqknbZWy
NIjYK+oBc4A0hIMJnZc4hkphEchWdwyFSy1lE61JO0kqmCNg1rXr3D5wxopoZS+k
b3KmKXkPUjEY7UiwrKPLWG5qwP6+TzW3vmXsaHONHQDzjmMpb3QAVfIcl9t71s+h
88AHV+rx4i5lxi1P9LveOWE2g3Ivo3pcIj4cEwqbU3bDmsII+/C/PqqFv3oTfoCw
SBJs19bRQINRgExpLX2fxUyG0HRKMUIKnChEa/7sIq9qq98r5vUuBOXnDa1rGV5s
ln9owCfY39GPJV+Qtinoa10Lg3Bb2fnboRUGMVrbLBOhV4lnHEnYu4stBgRKMf/P
5RKtw1cUwBeG5DIxA+AxpBt33Pg52WLAKSS+aNnX0Q+8vr1Fey0NQw99iCB5BxD6
rz51ENcwuqY+Uit2LHsfLDx1iQQ9OrER2fw+SOr3rVi093yTGdxTUJ9DGFoHEXki
65849UVGGhBQn/msIvWhNrTwByCYQW4Hp6dgPStrnux2U5KcFm3t90yCrzUf8JkU
SDqeme79fWxHdm3K0bRJzZ8/IyIkUAe/1ovFePT3LXlQtWvPI26qion1+iuOEGKh
+aJDB4RAWjKsS53+dLYuIw6X8nXkPOW8fLg/HlQGyIuU3oj9qdGnRAlGMyaa8g66
Oq7oiOULp/WzUH/+TLijmr9knFKDHkayJbyFzm7+ZYNFJKXVySqOG6k7slAtdd/N
FrttVvfwN7VGJM1HTD8Dv9cOs+d79ImVnrw0YYUUv9KdymN8QfUJ1JZsmnfrckNZ
r8A44LnV56LtCjec9csfBcMvLh8rrYN6hXSC37HkOLlIx9gvnE2dTUq762QSig4Z
0Cpn00Mu3H/UWtr7FATi53eyvy86KF5ZwGiGuRicskiqYWnstMTYTUvIeQiCVIBQ
q6Gk6sdAHbWiWBGU2+OVo1gpgNsOGAKGEYzOCbTG66buRT4mwmq/D9XFy3M8k8la
NREht+UuYOPRIFQY9N8gxpMCj1gDBeMoWs0kLB9Xw/2VpoEVjDUExEAKXXvV6Zux
QLQZMkypXelqmJBtzDj73rZtvUh/yTpLNObn0807NV+ceAf4QtxQgF30yKGmaPO4
/nqQAjImgaQyoN2uk88MXIx9M1KYiOmb87oA7hhzoZWKDC51Y94PrIjg0lcF0PSn
dpsppkFH4aZDABU45R2/PFpODKEge+WU45Mc2dFCGOvLwwfZB7aNw19pS4A69oWO
bXikTlsTz+k75GluJaEygpSs2AWsPevFOE6uRcIl/jZ9XX52pAHauykx07330cuC
E7jLdThRG/sZSY5wWJQo5pioC3D+FsPPPet1BIrlfYNJVYMEMek0Js0NA6bZjNWy
u64yU+9LCEwGoZgnk5HAmXEoW018fLd6vTcTrdr8C3BMh0EOLIcrmImhvpJcfIaY
2ZyvFpIvwrOdorfs+Zo9fGt7nhyLRdXTHS1GUYje4/hUs7dIbtT9GQM+iRbMXa8b
/t7Aemx/k0UAHDyin3Ve3kQYPErzV/4q3YfD8XJeFxdoua8aUDZsEzXNK0wRoHzX
tixMBJ3M+yRjCKuJ4B0PUM5EBKJUHCJGtksgUFA80Vo9/gqg5KmimXQRE3mbqKLC
2hBsawShAAgZ0rwMp3GHropD/RCoVLpU8qnRK606oSFzT8ErlMJnwdlNOEaDgGkO
31KiNwEtlWElkf5IKDIFJAFWvVZUEojnxcv6XPuWS7f/JLLE9tWNg0ExE/OXf+gg
eND1UcdLLkrEjC2gXvZnvulWTCwjwxl8lPhraT7NfB8vljpw3zKUerDAiPSMvmRu
DuMYbvoRvML/lyPS6opGpLXMEMaUSchV6IRhNarMMyYVJrixSlmPWpd+R3fdL0MH
d5VWvfh8WKbmd11NYasr6tkkU0Qaz91kcwIXsNi8scfZenpVVM6TwyPpP47EpsWG
oQ0gRg5aDfpPGE0+b+/11sWnbkQzCvjBcnDGUoLIqGi9uyDKaxgVyhD6+CDtXomQ
YlKoE+xOJCt3A3+2JzK0KkgHsfKlI/N0vHZsSb1ZGw+7lqqix/xBf9/3Zqjy/hdZ
HvKy/K9sLbJzcRkTtBv9O+TaMYQhFQS1rWsVhVBcqet3twiBgXVNS0RsgZqKfTkE
K0srdJJkVBmNqWvyrNUgaKemiPzL8BSsjtd8Pm+T1TVQ73Q9xlDzMov4vLNIppBl
Ey01OIKMExR9RZBsafTB2HHAh7suQvT2bouoci9TQFEpgEj1P6d/f+zSHm/hCiDk
MKp5kxizadnsQ6FBJEUrWmIA2eIzi9eZtIujK+Wg+U2MFbTvp4HXFl/XIOER6QzH
gj5NhNUC+QEmlEMgPQ6eAX+NvQ73RMRx2j0ymZoSIle3mUrVTgpBrgDvBQWzHzIr
jFQ4jNQfLsnyoeSppPyXyioiAUhx//jq3fBVRvEEk2Ai4EZndUXKeLBhGnzCM6Dp
SG21aulkF885dY2gd8Mml7AqEbtwiekyc6AeTZimmygA2m9zVotbNkivKDHygKYa
orMKN7nD+RWMDbw5dBhnxlK3Sj2w1zQZYfVjb4wCJFbQz4deglEyu8Oq8bDl+JPW
oqi2jxbX8Zz1ox1Z6pRyOexuaMMHJhN6fUcO5EJszr+cQuq6CxfNOy20gg3W/s3Z
wwMF0KCDtxcwHkPXN7R4dXNLiPjPRI45QTzXC2s7ZChEO0DAKrBsYMas0P80Grt6
WeLwcG102qo5BW90C+6GD+ZhwHAvkJYtyg5Kw9OIDqSSz4M5QGnPlqt23dKPZ08P
Gjz+muP1Y7/HEeiNC/0fvx8qepPh8BzFUHQxGcYKTBjnzBY47QzKSjsqYSHHP0hI
xG5n/a6m4WLLu7QjDv6psVnRWIIEcAO2ij6Ak7G1L4h4YV+GzCCMY46Iz2d21xrD
Uax1EcE15QnwhSanafUrBfS/+W4k9EbeQNK/Fi9ma2Lfkq8VVIiLq0opim+jWtaD
54CxBMYR4AMIFA1YNajX7G+4NtkQQIrD0zKtYTadErS3tzGTg8OFIitnwVhNtGdF
YnYCy3fCIzzSip/fqkXP8XGoFGVkN05EqQ+oZHER+g9cXtdaPFyVDaQrWU6npUNo
xnuY811qxd38kU9I6ndiSlIqMYMU9lk4SWOkaVWKNLaMcWVJT4dqArqybfVTVb8+
bJ2+xg6IkxdejxtV4j5HhTOwrVNern/b/4s3SwQEITXMaUHMUgjQYzBEe2X59frH
yl2OD0iZCoxpF8jTyygNBADZDQyJQIrUPlDOTRrtm760pRxcISI7g1YhaMYVqS2J
2jVpPl/IezoUWainNeyPwNNHLnJidCk3YcgiKrhNxcyQhysUs7DEoS8hwwrWTaH2
mDDidJW5MwJNgEd3E5G2FkGWcExbxLyKkDcD+EipR2cdvl3QbgXOa71syznBw3vg
SFaFBUlee/ovFk7jwqf6EwXHLDYM2GnQBFVGrFjig5DNy/14/lIdrdGuBDPnRsNA
9JH++jA2AFpsnNIraWhUBh13xAaRD3RHBVmnKUwWuPYh8SjsVXevYJ8Q0y3J9XGj
snUmLExTXOiyXNmrV71MoWsp+Si6sPf1hVPZ1SLpVhjdaAybY2DP0ZMn/kVW6QBf
akG8KoMGKvZFs5TLOi8hoGXoW8gCOlA/iBgt3yVGszWjZz/NZsNSE86GSdW5hGuo
MEVCWwZH5cml5LTi+PFwPvIjQ4QeFk0wtscTxIWoEw149MG1Tt/IGzPHK50PeZZf
XHxYrpzh9/5bJKb1SknMzAWM+Hb8OIYofRNWyBaIMU/Ke9PB4uFFi2FOwMhGZKYj
L2CSKZb1BNxmHm6U2ln2ubEHJGniywyAgIJWQz1HBinUCn7Y37YOjIoQdSVtzNm7
/f4xUm7oKh4ilst1kDuW0yPNAC0Z0vo80wBNCxNF8cf87PwqE/WZFsjjLoBusqbR
F1sUBiML93nEOhrxicxQXCnLPCBpcPb1nBDY56aZF2lL6OGiNIREOYJO+JPzdUms
8b13hFBDETNwP+K7/AU1yLg2PbxWvCg1kL97XtKqG7feSIwSNI0MeyLfjM4ImEiV
YPQOZXUTKAMfb/stjGVa7ZruZzBr5ShRZE7I/DwdWguADNuRIBFF9Fr2QdIyM+iE
JecLRwrcTwtJouBB0NNBezuZaDtiU5QYcl9xqqXz2QGfidqKCjp6/KR+8kl2WJRP
KAgpaL6pChqIFgS9kSvr/P2FSIjUIsUAXwWQX03nKEetSMf6Vpl54WYjR5uIh47t
/aRuOOxeeOe7bS3GNuR+Q8xEWJn0VkmRAaRx4ucpuZXN+xsOrcb1sPCJxk6BEseW
3bDHFAKBAIGGoTrPoRjtL/SIQVwBzUQsQu+0otjVuHzabGENiHe2g/IaO17p+Sys
2gCvWB9lrXWRc5oNtOUI7FIiTZbmDenWhbWfkinsgvsf/EJApTWAPe1N+sUYHESb
Zmg5NXREe9T59mPk2a66jeW56XSsSBgFgRLFGkjdkRH+yWBzJZ6Jt+5amwvwvgh4
tFCoXEU65HSAFiIHbKDhejz9hE2zQqOA8+xGNxuUg8L1pFIlv+jiGThntaVFlpSs
kTeo09PhiJA1ZXt1koAYBE9swzeIDEEM+YgtL53hm9xQwnbKaGCx0CIECPv7V+B3
2ISHYyozD+hRDH/gejgnYEIdhFQ0oP4aYz8ff/UHTeaXde1Kw5+kb1kgu2M09wrw
LqvzXfLDrdTZq2pNpjr/R+plWK1ZxHqU3Ku5lyxWd1mJ1DKUwO1eEQb4NenBfP29
pLqbSusofGPKc+j2qzs/PXW6hQUcGPNZSYPhXFDwwmZDbMtdashxnPVUG0POL9Dg
KzFJB7TTjifYqaR0J4ossT7YNE9Kd2FkuUNlqqmnajrdDpfZ1mW7UewGJ2bC3i8V
8th8OaPozBfZ7XwgEtMnyQCsCb2IQ2GTcD9VkiZZYDDC1wbA7pCbn2WePsh2OiOn
raEmC+SmMqkLBPJqACi8R2boTfWCBe3cjiL4Cf1k0Euncltau0C+TPR+kBB8JlKr
mwWfThFTVItR3nTXgo2o/QGVBEy8Y7d6Yb6SgoCpJsCVk4qhMByEB7N2naYil+RT
dvXoteuqDIBhEUN40modJWsyo/Sfwbh/Uh+aBYQAdc2qZyYUhaisoZieVWLD0E4h
DVu/Y5VlEp+vaMO9w6j6IP/Zk+V1ypQztpKJfXNK2mMQ9ztw18UFW6tjThk9K44D
CCBx+A0BWhVql+fTDW2Grazsry7lRWeBrbApVVchmCm4nB8sg45VvjW8flzqHrit
FfS7pwHlJW1OTBUkY8hCa+X3OsJu09I8dxFtU+vrVx6I46jDyMe0dFSIYzegqOIo
+MiW/w+HUEn2/bIxUd84a8jKa3/RY75oiCmM35Jr9D1SkNkDxBM9IXmxhmWMvi9h
uGo3ggt9NMLh4CZUpqsmY0RA26/+FSogHT7UspsvtpV121m4d+dSJ8to4Jp2JMYD
7Sl5Z6QyaOArkF5TawzqAGUPmAsSQyisF7cQXq7VYGfwWEm4CElZNmLh5ASDERmE
tb9G2zzfTNjth71IJ+HXZEBuwuIlhdIH9p+6BLhv3Zmxa8fe/itY8wMu3XkA3lv8
eBCHAtjvQ7sOYMzD4Eu1vAH7cYg6OUKInwB2hP/0jUd87u7kZMycidka28OpBW3U
kaHfHvDUGpj5XNjattE3fs7v3FIgaS1ffCNFq5hPnz8t6VziwWLMlK54Zy0A50Vz
WmOQ/9Lpl4lnO3VSQQIUP+CUI2/nfe8O3m4eRSFeEOujVpJX/rCrT1xc5HvitQk5
V9Ao9HBIvg3su1524Tkppq78HVFD6HgCF1DI8jLQICaXIW7N+4FcTlMUvDztVm3Q
dmRilqUGxz/kpIRoxCLPEXQeWcBrH2oELlok/ukks1nfY2fy/A+MYs22dFvsSLV1
ruYb+Lb0EWwmZ1EYWD0kAkoYdLb/O433L40FM/p4AfBYXPAIh2XZimZYwOxcu74m
OvTawW1DBxhxkHo6LkpHVHVlTaFxa/DRrJyrfiq2lyvRNNTBX67Dm1x//oG3NTUk
/XN22uxuwHLL0/6yUjBUNIpeaUCCyrTpvXsoxit1y2BgOXRoDdC1x5dKgqWjTPFd
FA0/7BhREjv63Hf/eexcnuC9XRE/3hcocuWFdmZ1QmkKkkX8L29PSG3r8X3Tvw96
Ufl3oFk2/i447ckV4I/0oZQBxeC+1UfAxTZDhRmMtvzeA4JaBkVBDRR4fNG37CLu
gXuE64G+sUkR6vkrHItv93b4Egt47PTGCHw0q3CggjmAfccQJ/Laa0QsjwOxO/jD
6O15lH/dPoZft6w+BMtQlPXcJ/gH88lRfQ4txgCYoIDU1ait69Oa2h9N0OTuYt1c
2Zi4RDa5RSNKkyDDw2WnPwx5KCmt+D3OSwVpu9fRpkk1/+Tlrw1sKb7bTMTP5JrC
I4LrqSt37qw1iReRNMgfy6Z6V1ZFXD/9HcRtUKQhE1TemYa8MTeL3lbbZhYWMuP1
jUc3F1iJdnhai7okBwNVMLJ4Nf+atAa8JqywTaHzvQ49TmbwLNr7V3XAUuH92xA4
Hi0KrRsqRfquiPLjlOaayrM2t0omvD/ORNZTZA1Zk4AmP35pOLs+4njETHyfMc6I
yGJJmx2lwmclLW/RMxp08aoDLKtejno5gqhZQZ3ArvI5NwW4Vhut4RYr5Y4CfRfy
K4ZWqG03+YJQNbdR+F+q0OtCc9uKE/Qa9JeobFPffUqPAGyJxXxvgKFbjZ/m/pGK
XOwMnP4Dn81eoLyjutXL62giGzinxoKy5KU9BPKtnPTl3yzTQjaMM/yY6N/Oyz2c
R7OCRBIrQZPGWxRyAhal5xM9+M0dSXmJJWafcQPPq54oM27AQLj486Uf3zQyEt62
JCg2M4vtSwByPdBAgOZ1FqCJibKHmRhE1gb0u6JFGO+NHFVEuS7y33Wrzn/sGMsw
d/J2QuRHUHTidin33q/kM/KW8CzYXxITLrV1AqFQJDU56vseeSFktxdHO1qUzdNd
CanX6p27EXqCVnEVNep9eIwm/e2fUEKIg7ry7jyhtIP7P8ZcAB0UcIbJmC7SYc19
bMgK+GVe0psD2NtJTmC742cJuh+iefPtCSmohCmxKQUv+XY4gsVMkwU1sPmHui+A
+02rYszA4XK0zdiD2sKhqOT4Ao8lt9B7mDa3HbRA6oPv9QWyN6T/xhKvbClMUqgd
uRUR0muFnJYPgphFZdTMF4Cc3qJnLa26N7HNI5LUQlsBon8yIXPpz4Oop08mOYfr
YHZgQEi6A1bcK4PqMO3NnRuopWl0Zcqg4tM2cwL0DCSMBoIGJzlCN1Tmm+uIjang
rPHIgvQxbLaTgzRrl73Msje8vPbsEqFTlYlx/ZRgiiBFnekC9P4Li2d3YmZuDI9k
FvieLbd+/iDavUJMZkO5eMYITTXDKEEMVzuGQcdANR1FMadrmJzFRggwBlqSFpQ9
NbpzOogOgA5z7eZaN1U5wOPbQyJLFgUnZu2hcaEe73Gd8srx1c7R/5n+cDsjliw5
GsCGsjhcYizrH+Pkh+2tTQCIEyog17pTeu6cNeann9vAn9Or7zUkUMvvX8Z5cRvG
2fsTxbnR2ZUCPdWRWay+Ictf/m+8ZYAUxI7B0nrpDp0XmRxIT0TePtYwZbSF2BwI
O21U3ulc1KJK4sE4cpYTlUmMHBiCtBFlSK5KVTI27s3VlEvbC4nEodgarv2ZOLod
UHTlcd9i+i4LAZx/ODJxNPC0DR6YFpMXspbHpZCnqkBTFhCFA5wn8Cv+uMRifTxS
qhY/+afjA/kN3bA29lKu+mdRcO1tliQBER5Suiojy/+GI0GZyIFASOvKsgqpgTr2
3fMXMreeBC5J6/Gwg6ukbmc1rEqs08SQYGU0PyAZCEMAX+JTklb6EYDhjuL6AxWv
6j3JknMcKtCBP7F2uL6vfEIdznkuxjWs5BvqJdzov1y85u4fVem1VKEfaMEpODcO
sDyP5uhLEYxZ1lXCnC721MufNehWRFsM5U7zdHG7x7mkEmVDKoRoz+cyjHzf80R5
qmSOC+Su5v89ulAEutuUK1NSZYWE9Pw7nwA6GGMXP907BwSQ3VKxWDlCv7Sb/MIH
2xq67e83nw/oMXzeOt83tuhnJtah8YcTJ0XzJJ6YcoY5BYyp30kJxGW1zRR3rSjK
nO9fxNyBOL68yJG4zYEj27sDIb0KlV1HX2/SeDE2qVMx3iuubMlvyOjfWGHE2p0b
k+oG70YGRnqg1WHT0CUJsYp7c184wRQHDBnWrcsNcCyyh11TirmGsAvuIEZyyIBO
ZW8BEOkyYRLFyPLIII0SBLtmSWzcWVDAC1YoUY5XwmYzCzACsFongReSHHHzKLYt
V1c/LLsqLG2uObdOlOc3BR8RsN+6nCzFu5XSsMM8mHW1MuuZjM7eV1BLFssL9DNz
eSQX40XK/PP9st/9Psmtladb1TxnxhVZmVxSqH77Slo3pGV96z5l8N13PtnjPLJc
JFeNFfRC/9ljX+ISCvvCNMyXVjuZrrndPycvqORyGVEbwJD7LaiHWdP7C3bo12Zx
7oizeOtU1167odxstN3a44YU4FfxTehSi11AOg1D1ceTfeIGPUT85BGw86AgpzT5
gWAuMRj6/Rcps6M7cOGO32tMgoolK8XA0ibzOysYuM90kicMT46BggKInjSkWUFQ
VJsV7KDpZZUuoROrjmSzbi4YMryroP5jzlT170zoSPp2xWUIgyUMVH2dIF9UHfOe
9Z5m+JUrfvmSU3paXg5eZKb3+iHLD7Miv3dC2ch8s5BnQifGuKGJVViXW7ninQs/
g5BGyXZGgDTyZ9oFyKCQenbdXwUvhrCgobRgTmNrsgVlAG/D3FvjZ+vDQzSKrUVl
rgFLL7C2Ffk5je/oKmwG5KuSPVaLRIONdA7uK1i1qMws5dwO+jwGfUnkVl8LZxeP
io8L3Qm0hCVXX20uuCSCokQGVSQZwQ0oiE5XADgG3ACW3zLjK/wk6tE+RpvKuvyX
o/eydcxvGLpGw/NrQiLbBmXutwL4gwV05v5KaBdIOe5dL7m2vztAPb0v1nzWFAHz
lzQjdAP361D68nNdadVc6AESrf7s/cT6jKy6yt1WxsNkPKldr9xFpgbckGp+xJRn
VU4OUfBEOnNDWGHJXW2ReiA9h3972lRNqg8SOQI3Knz3jrSgE7pYYTEXFqm55SaW
kOk092tXjAM1dJYxVB0feS0SuF1+wky6hOVD5W/EqBE+2ECk2W8HAM6sWP8i54cn
0IsGAYFfl0W33F/u4yP+uMtxCejD1R6+9DB1Jn0Igx7l7dMMlWH3vryCg01AmSbK
FSVAX008mmigVlR2IHQbOXqVo+JjT+ovd04POhOpgEu+4nj00u4xaR7+Hf5GW9zm
hRorepG/4urMlyHlkfJK79HcJLzstoy4mvO1TVc9xE17bcWDd9yfknf8HHWuJP6g
35UQIzE9pMsJzMs3U81sGHTXoRoriPLMvDY6pr+Yf0O7YOnuFThp5WGnv8DuoYqj
cVdpBE0ipr/b1OOd2iSE3Cw2VAFFYvuxcM6CzPzOVQbSgmyr22fJ9adPzTXKy3QS
fay7qbsWJ837ObYR3aVjq8mNYYmeM/Ud3C60+xc+ZGYaNS8bVqGTcgFFaf+3Ibcn
ryi1lwlg+jzYGHTy8Z81JNDN3KauQywjc/s9cX6sgWIBU95z1IwfgR1YyJsiwQph
7wNF/SnIFaZEE0AEVXLwOaiJlgjEXEYJnXWu9CiL4KFIcyMXbPOjHrpra18fy11w
lJ+IWrWEDBd63v5dxe6k+HEGfmxAdpip4vi1NBT/SjbJL/orfY4ee7CPaQq370Kz
FHKQek3ihB4O8hgZXxax6OlY9mdFwHhMHNRLUgGR7MQSNGw7Ju70+vo9itO/m7iN
vptt4SRpqHDZZk5584kZoErOYscnxXHPrdW+LaNwbg7AwvK18uk75zZYVaLZ+DuC
VbEDIhrxd8snT6USp1n0bRt0vJyngC/GEQvAGZ9o1I9Jj9qxbydT0EuBvbfBybBx
ehzy99UKMqEYN5ApzwVNu8LVJXMWre1vI/P0TBtuljSqWlQ8O/xeYy+bN2Oqn2GC
qclDaLAQ/NGTgHLKUlD3Mb0E2GMDvBlQIUSl8lVzvn+UhwoORRZhk/3pTv9lmnGM
0rKCuYuORa0rrigCBXas6YHUB0tKgSpr0pQ03usGa998Fm2nVJedavGDhYnyD/VY
c7Hs98D+DvNkC/l48pKm5FyFTEfAJB4wd3rN1GP5mIhlWyQqJRNT+a2WUjcF4glG
tNwrQ7Qi6H0+l0JdOshjV032fkKjomOVyiVxFHtgR3N4UiABkUyZ9jG+y7cn72cm
moHQvztLEHxvSoQFIFIl8UzfQ2Gpz2xsUt8gH5K2nt0FCf8W2WNXaSQjtPihOcQE
ZEYeGREC3cAF9dWWHRB1A7sC+BpvGyo3WUyI6oL8TdkaET0ecLgg7kB4ml0fW7+n
KIEI0l3QnupBCwJK9b73oY780hmnle8bOWaTmEYmejjU64Zf1cGHG7n0iG6xX3oO
r6fSPz18TAz5uRC87/Fbo7IZMs8Cua3nc1gjxFO2ORAGOpWG/r3MYBc8/6ZWCmXj
0DAIXZL7ZdFFiQ2c/u9G4VgCtjNew2I3bXvqXSoYTjiwqb2dyKf664i/bwn3+HST
aQ9bheFZhodz2v4dX2KVjlBaJUubIeS3NEvKZ7TDeGv4lcX2xiREwE/mmy8BgHH2
gW0iMf17PWhtwnoB293vgP0grxCIcYrEwj0JD0tAoIAmgcddnYzTKlmv70TBBQxm
ATdU4hzuAmb7XBfrqp0AcLHUNjllpQK5f7U+XKnrQRRsKklFOK4liGmL7xBeyFkp
JYcwiIjuptn9qRkr/R/qt1JPBvI4g6UPiJuaET89kPFOcEWuL5YTotq9SHnZZ26u
J0fBnYIjxfo7JmixS0Dq/kNOM+t+5UIPE03N5humRhS+bIbVggHtVRtIPaFZGDh4
wPC7IM+ocoe7XYL0atA+Hk9hrS5KCttzs5jVplhvpBy9rxoQ/hXh+aDM/G9c8pKd
WSaJ1tpbS9kNqAO6NQR/eIfPfi9j51T86AsGPVudDy+3xVPoc1b/nO7ldRlzcM53
+GV1rs1l4V2hn2BljJTg98MqkwrjNwredYVsqIZVx154slQFEWSKQXItGqfZD0w8
ogzfIdH03L41im90VylSa9XOERgsG3uF6hGp5kkB1cE71bWea96gHs6+lOJPLEvz
TSK7eWVe2zGYYdpC+jbhxg7C5fLqlBdhcP/XxRVGjZe7s8n86U4mCFVLzUIZL42L
HbrTsRTS055RgL5kUCBjeyD0aRh2q/mH7v8VHoooMxWVLuY83ht56lC00Qlze1D8
iJPmVTNNqtRc+EfTO2IWaHvTWXMEDk1eyo6Wal/LZVYa+mFYZnnj99Yj7pojwujE
bzYjWhJ1NhQ9KlddyVTydinTPthcMeBonu++s6uC5kKDY54CWfmu0P/bWkPmITB3
9ho8sbirzvmCslvlJUcb5y+jhO/P4E3pXgiBFfqx8BYZmbVrYeqt+FFFRd1Te2mJ
aGHaTtWXYN8x90o82aYAxO12yGSHaqMdx6MK+U8gIAuKp0xQpUnrfiRJWDTJhQ1o
YBTo5FIEoFcvr28ng1szATgRS/kMp+I2NXZ9vEfKfbC+au4/gEwhGventoRA04fJ
nfuUFXQDUa98KTK8qvkZgfC8bhwVgE/0aEl+uyybw5OMA/Zu5Sa/o2aCN7V828ps
y4V4Kn6pK/l5W7YtxtQyGPm8ezvxyy5EM7Gs2F9yWzFUZHnc4vwx5Xqpesnop/Kc
6x9XA5GfnkBNH75wsjtOK2LHTKZ24T7joTt1yLeH/P3cTQZehS3Qzz8xdyWu90Ow
+lIRsx3oqnUzMKtYZU3nXx/+KfiT3/kdNLTEvV68g9WPsNFJA94GRINJ3XvoBhh8
H754Dg+Ice3vZ3xczM5/laEdtiVcsOb9JA8rOq5Ev5L5K9Plth+g99IKJHwS+7Iw
yki0adX6TJOjYXRQH0YAl5959t6kPjV3vV+t3st73ZTWG8k7inXODKqXX4OnWsiK
Q0T4pJ2HOxfdRSKqEDOQlBbhFFVrM4raIS3zsBVyEV2Tf8MVb9HDWwnBmYKW1wJi
1Fh1vJGA86TbbjJgDcfRq5i3Qic+6hyCJZudIJ+m+Qet9+3sLzTo/pO5QrCNjHdN
LvWAiAacZsHE5Yg2C0YN1jH2Za+O+MRg+7EL6iOb0N//9VwaqxMjpUGJ0r3ZwDHk
C2Sh7lsuaWBCockSG1qkjCuA84djDPBjrdFNIXs7GPSW+RCi2JHiyysFdlUzZbb3
jA7iR00k/zddhxwuVCaKb3KdlivIpydJvzfhuq33HQBBOeFQlQM0XMK5erITgiYm
cv70sgzoZegICylPA+uKzkN7ai7BOYM38vAyMrBAZXwtpUBcIjNfJKUSxibFSYvE
EkIVTwsfBNiRow9ymOLAwoia/Dbp3oxTvJ1C73fD6zP3+dJIkRQiPRer0VeYwpng
SPeOe2XCW3BM6PWfInJkrQMht2ysdS2rvIkmqX8Gkqv/kPME6+c2mRVv0ieEllBP
DPd/BMrkLRwDwBPo3IBQjBG1u68pBtVsAZtNnSRofCSW9Lp3SHGsn7tegb9CikVf
jVZFm8++fQUG2zo1dCXd6Ni/3Rb0jZLorAqLzxz0Bctofm9Qj8ZGEe7lVz8CCZ36
m6AHBI3P9zM7rxOXy70GQZYJ9ZwK1Xt+UV/jINHGMz/k3pBkAQxqCYZNzHovbIyn
FE3ZX+MAn0H98nCmB11uEItpxYyGjVm5atVqOlzyhAd8Y0JThmQNVIX73e1FY9kw
N2o8saOmuXs/3eOMFgzRzYmRk870QyR613yRh8MV5nMhrcpTAFGvUqgHvfYXIomc
8fKxP0T9p0ebvv1Fy9xIAE6pcs5Ld/ZL9Gh2VsmrzRUY8ufTdHWnE2Efea9QHTNR
XPDa2Qh2LIaSWwjE1MwCfcsJ1USI2PVURj6uH+5pCaml0mhOlpr8EkpQzTHOjLHK
it8X2LuVm6aGGHuUaoqYTetNSA1xG33yetcE0NxH+cwgfZj8knAbm4sOs/cCS8Q0
MtwGrR3rBmvV7UdGkotoKCSvW/FTUECBnj1HwNW31bMYquK00GhDy+41vshV//ny
rvRKKFdZSto8Qdse1FLjzuNltIbyBN8MZWkOxxx3okpNboqeAjWtDjmdmvAva3+W
/g22VoWXcyXJcpOlR49i14ZJ9ymuC66YH/BUU36QdYR+9sV6wfHVAIL5ajy+A2pE
zyIJLp9+SkN7uqp4d8pl9wBkHXf7qRtTL9qbfmyAc4wR79qSiUbPEM9r0+KSjcwM
tibWos1/OqOc893SWdkLUcDLZiuv5BShgbB2/oyZGrPwgqkkK9Mn72y0Tweimixn
TGaNoogItVeyZPT+zcqv6yjinYQI27RP7xnFyMDPcLiKXipv9i7/IytAnhCZg6dJ
yrc6w+RtP+wh7dhf1dig/iROODN7a506J/waOM6KOn0f/s4ABkTLq/rKUqhacsPM
56I1LhYzhZLjpRD2jaAF6gY+LsR16JOb8tEqwfzikF4kPB59oDStWrk0K0+2TY+L
ZyrNBwFt2cqiaFMLmFXa8DmtQwW+C5aLU6xKhSaV1+7hhym33ictxMzJurN3a1CT
gxlHRyAQUryU9CctukTR/OOxUfecm10/L8O5MvZhxPKlSTknLheZ52GuljWEOJaX
fKXH7gOEoON5UgNSc44f/rdNz96jImLEDIqYUcxzgrgU/RP92DSzKTf14h4cNhbt
X1ET2vE5mC0Q/edl4EdtFm1Ixax1JA5pqNd9sN9fgQ0yuptQPxY7w99CapjWDHUu
nlLS9lWUSe/ZCp2YjIcH3uJZEEChRsSuqAaOS3nGh0DEgMQ65LqcSj/uM8+OPRAI
thO8PwjrTNdTyrwPkR19RtZYSyTBKb/NZAF114rcDu6/KQ5nJhysZ2Hr0a8QY7JF
hmm6bRXKz7qe7JC7Yf4T8OAi9apWSzeGcEEs9tI2TUOQora/f7qAQi8mFI75i+AE
Ef6u+3xofjiOw8KEPkOxrhHyMynkG7rdiJM/A1zXAOPHWAWz+8cvNBZ2fwunVDdT
TnlS0g356jM/HYmtWf9aTGkZL+Divb7zAZtmixXv9qPl8At3WcVz5ckkJstzaB5N
Oq5yPTqj2dZjb8Wu7sDnYfRhRu5J+cvUnJF1dDbZtYuhMrQHtnuK0Rvt3spX0kF1
XS/Kj9v/K6c5uvsJ7WMcl7Rh4LS2/3uey/yoduUSnLHBCVUmsZX4DW/9bL0A15ux
evmZ7T1zDd8o5vzL2n1teLh2aV/Va5pS7y2+4kAdpDRJzxC9YQPTkwWjbmpQAsuJ
TD8rC+s2plMTHgY9eCH50QpOIQJO/JoE1OYtOzDLL/QlmjBDLV9vjhoHdEaSRy7W
SkLiFGOeAN7eNP7HgRbcdIYE0Z1rDx11/1bpfvfC+5/Trj2k7o6HxgUnZ/rPpbN/
0wUaunq+bLWAC5MSGAoUVwHlu5aU0ARQtlr/biXRAvE2eoQ1syNKnpWe+ROUqDyS
ZsP5257khexR/Ddwq5fT/XgpZx6HpGaA3U42ShJCyPwAB4MOJsrnPm+OQSnmFtJV
whtJ60A8F9fmiDGPswdPIyJvqjh8VBgbSafEsDI3S3uowyEV0UDHac2W2Mxwl1JI
MYMQgWswEyl47xnIX/YtkwS/TyHvZceXS+a0R092aRA5o3CB5Qw15p1j8DORihoB
riOD2ReJugDRD6aF/D5j+kzF6Xv1WKdadFWTx5PQ3pvjaRwtiNYtm8CVA4EKFjzY
tkxCwtLp2BzNI95x2Ms4Jye2GYJxJ7cZgOt5OcScSZAXIlP6cQY8VZ8LlJWubg2E
VePnIZfPdXHsJST8IwWI5JIRGcH743BIqrEcChU+IEwHhMVEZh5h8iHw8fYdDtAi
X33X+iHlONI5bdya8arEM2pA5IUHzmtgJKdJJCOCh+EN/wow+2zEngntWTuPc/Wq
D0we7tjZSDWB7ERuIlW/8+YFEKBKmdEXHsnlKBiCs9L+Bk9xr5DM37d95Dsw1+U4
xBlea3+Q99cmzDA8HR7yBpcWsJbJ45lBhriBWSgelL22vfvnV+u3XwdcyzIP+5XV
r87o0qtm3mR9cEUMIh72chEGwoosBws91889dkDDp3YkYpuxUgWuBjFZRmyfBiO5
XikzyXY1zADCOP6IeexzMl36zz5id6pWag1mVGkA3kgz3MQzvJOgx4uPVT8UWy2f
ouKp6OZeuAmexuYJlrQi6PW/CmWyd4Oy35Q/wcC2IOnuRZEDsmrZoqj6VjjGe8Sx
NfZu2t+E+r6c8WQb7pS41Y7F/BA4T3dWE17xiuk8zho5BYhY1Z0QW0UZEi6/Fk9/
83TKJBN2ZEZcB/WH/5yuF2aPiIwy6ddcde5n3Vw/zCUIZ+ZEbutSRxR2JiO6G93n
xk3WyPjPZ8DYDs94G7zbHjt3+6QYTfY2tsBxPsCq+XjxCU7GwsNAvfO9Pt8mc2eA
4dFv1PCBfRf5YqPQiY/BOSdltrFRkQYsJp7pAP72uoRQkZzzwRI9p9JsdMPYV9z3
IlWzB3NIzP4u9QusOy9eZdqaT9nzqejtfyNGHLE2oRtWT2MilXc2JXfjAt2jH0KX
mzNsqLkcX9rY7RkWXFXnIuCF7rMrlXIpYXJAfVxjMissTZicNfSUYPFDNRKC+dE5
0/wE8Rjag47xcFVxVHlasaq7KNQ8J+2i/hflxdDwgLj5NNdECuS/xv+B8k+d2eHb
GCzT/Uq284lbexCbQ9MQSS66kFyM6OSWFqeCUhoD71JPMxY7h10OHkY9oKPselHs
Z4Th/AsgzTAtwVMI7xSpYaWQ8ARnjmqxyi2ktpR7qmcej7t+EgF4OS4+isjFX0b2
ZNw146vO69u++pTvHWLm511hR9N2971sySV4j8NKnIk7gxZTMSyCNnxEJYFKQVYk
FkZQXVzfNKMMt0MV18tjIADm3a4lNMfbBGWFHWsa45yfBPr0Zl7aj9tMMa7zzOTX
WmeAuyMDAQgFPBqIRNETwAlJtYpHFvEaLcE2Vz8YAXgWDtp28dc7HjK0471U9JwZ
aIMDICUiPNAqe+rjOf1NIJ2zocnRl6UlZej4RyMhfO2Ay6c9DxS9hszNrrdO8cDO
ehEQL2QjBRsYYT2Z7qNoYwFeS7/mnlpOBYEwxYPUFnq5ZQxV6Sa+IRnvMQU8DQq7
Nckwn1PrFVnUckQnLqBa+3dCgGYvSKXWP3fT64QU2c67C+Ukcjxdie0G9h/fOa9K
U0x10ur0DGexNoLNLC/agTUM2bzTSuBh11jPe5QDsB6Aqr2t5G1HN7/TY4+AXS4Z
hMjHiN7H7V3iWwn4GyjQ0DhJS4K/M5ciHYyrCL8+MVExfLC/0a6JwOidJxGdnBXF
+2oYc9wEaDM51RRaM9UDfLcPI/BarSHWMz2VmKfrLTyfv7uWf4z7wMVMrwEsM66b
sbaVClfS4cs/CVZswUHflCBSE2LbGwU612uI+93bmc7/FMEaGzVAIq0eoJNpT4eI
VsHZlIDkPOsLUxZ3+M9nwCbajNjPfwnEZDJUTc9zITJtwkys1JqYhAl/I/MFDUVE
qFR99LZuUM1jQFE4KUWb2I/m1zGtV6YwKwt5R5iI/hDs5oLRNld/N9m+3FxG+wL4
Rj45EvswfJ4lG/tuVsmXmSzmIOnCsiORCZS97fWNw3XSVDzLZr/o/h/efobeVyA1
r0bYxF60OP8mKMS0zwltYluIXpMgWKkF6AwlM92fE/ajcLbjE/V2RT/nmnKaUDCV
LLWTQaQjXzur4seYcxvB8K5INeWfDZEDjrNeb0as1qWZQKzL7EoiXZCTXucM2BBr
cbKzIUhAvPqdpGmKoP3xTGm9KEAcOs8pDEiBSMPGfF8E51uu7BUV1KhIc48iyBnr
wwhzCk8Z++p6hNbR3MFT2o37F1o7XoK38PA3qUGWO40U9KEalZPtYEOOIeV3OVrX
QGVpZTXrf1xKVZi4fgIUjxFGDfDdN2QtuPOLNz+HsTOGIuoMPMgarIJE3RNTcHGC
dGcV7sR7c24A4nIY2wVDJwApRvx9bGWMgRI14p1XbpKbQIQzS+n5sG8ALDkXlvy4
3GslHgV5VVRF/Q7jDgn5NDHgnwb1wS5WVPaIcVxdbgUFqvjhTvh29kT03oDYB6mg
LQ7cZYFo8QwMkz/JqhEqKdVO/gV18omegiRdu91F8wT8uq8E/29VoCRWxGPqfs5Z
glOMMXJAFbPM0qSMeEePSFIUMUlOzAQ+lyxitZ8c1waZbt26e4jLBuNeWQW3irQz
skq/d/bgA/mFaYnCTXR0SCwTq/8bNh0O7peNEszzDyBG4I5SzQV3umsKVYhL9DBu
DsClDCc4mQy6cZWyjqPb0Va/lyivcYu0ta9JD384+IRzU/TtjsLGRO5ABjVoA5Cw
pACa/vsdEhlqTEaatJRclPDLpRz1LcVIh5xcEv39y656K7GEL+WAuJzQCCr+fpYZ
fKw6Y4OaAWACPPgmTc2RDQQKfWFNZGZ/kACJ9DMpRBq3zqFIlCduOAR6XdF9osMx
3f3fUXxHIO8ZlVcsdJ+hR+rta5SJktTciPSbojLEA36PukXmhooS9oQ0n7wmY6qF
5sLudOJ+vtrKHYq3Kvu3+6BhupmBAxtB9pv9pO8PHqW2CiBpoF8Iuq0Zd2LwiMIn
2fOWFXv3suP9Ea5c8GElVu2/FYLjM6dfIyiZNYNPk38990/cZ6Fe3Vs9qnH1Zzh/
/u4PZUfxRl334qcgQll1efadZZWXXBEFAV5voiCxH5g7YkoCSNj/abTb8325rsdx
pG2M6RJASHFCAQp/PAttACghhxGcAvWe1C0bKfew56wefmGenAoI0tJAZWAKl7Sj
9Xf1SNaAHQmt+G3F22tv9zwWR2x5ckY0+ehgUaXzUqlN90A+zDuAppsTPB/b1ztK
eB7JuW0t243IQf5WA+lB1cMWY8xNDUTM1UYKcMRs3JIQsgSSEZoRxAMuhhXUtScr
CKL6EVynxKeHFYCSeZo4X6BrGGynpiG8GNXNQcj28QPWnSTs4Mxm6AovSoqa6/NF
qeX1V2UwSXN/eLhs2EEcWnuNPiCBXgB8cq+AEk0dzm/D49s4CCHrOHT9ey/FWPNo
kSkgYaf+ltxI+eJskIntLbimm8W7KKW9RvUk2bmZDD3Si4LFY+7iyG0rSYwUiOjV
N7O+Kqgpkgk2VwVm5wHmJG9a66IvBMcgXCOCCy/42G1lRKlD5JsXYK0SEXR4pbAd
fKRqMhdm3D+AFenigboZaos1C6lFL1IBIj2ydMLREV+rhfyZ25ozOYZ8Ziqcwr7X
f3lquO4jyMk+G9i4luAPL2aEnqOXSiqsQdQRfNEW5Oe1UjP3DkqYBH7i7IjUL9s3
SMX0+lZ4xghr/Go9tgCmBiqV33OqQdwp9Usy0xokx8iDrWa0U2F5yavb0QFk8Mr0
dijQDgAK4/AdiElHjnSNspLYKjil/OVHiNPW3a2cqkOPW6gGErmB+0d8H05o0NpB
xkNS5mfni1qiCv2IK9cfrX9L5jf9Il7lC4u1QMRgrvdAwMntGWm9q2IeVnoo98nC
Q9ezqFi3wz3dkxLpNHLmRC2ydfVUi+mNo3PZvrJtfXkhGqNGTGcsKuV/qedGmAvv
yRyCJEMnS/H8yz7JL/bQja/GhxQI5BY1Q2bOlQvv82dElUsN5uIY7cwmwbSQQLzl
uc/SxKL6gZw8tlg3AYUQlxNeHdv8dOgjjyBSDk6nB4zrnWmZNHsizKF2OMeVrcjY
mZQnAre0ow6Gdf++k0OS23C67q0Ykvicm47vsM4K8n+qeQLw9ckZdXTrEB0NNC0y
5/xj7G8ytWLQNFVcVn/xBoyngN+SuHdK5RS2beUyPrciBGytafEwl4BJ1n9Yw8EI
A3dBfYmIRW2wE8peJbr5FFP9PCF0SeqSWCGt77bwf+RIXHR+9yKmaMTU6QA0BEBx
CvGMdi1nuju9mbObt/fBg0AzdnVhyXFsziaMzFmL+bc9a4YUA7ohMR0z1KzFFGgx
DS0FPvtpPjNPxMQEMBc6pcHXRLV4KHyGgPOTpb30AgGUusMsVEyMy4KBvm5MB2rC
aSz3oTiQqyRGjVsWGYFba2+QCFczxKGydPf3B4ItnPPHb9F1dY/hZZmCPJHctc1k
P+ozg7VH5O5nab77NP2EQBs4aU6SRm4s+cfNsjphj40DuyAIjTJBWKg450qYGYEn
RWdj1bREhqCMYW/OE/W5AvRB1jlPCOPO9hKZ85Vt2WNI5fabQVLbusQ/N+3w3PA6
ZVUy6UBU3ZlP/ik0/HUesDeDWFSroo+VqkjJqasEiS1tuJT6ocLBNwOmcfk+zEsL
W/KfUHrEZJYX6H7MIaO/f8IRPRtFDNwISsAzmw3Gl+KCMtyKlXR73k1AmmHBSbmS
XC/HpThG39Tr3odXWMdcWPEgzDVtL7Hm35EWi3ARHslkhR6sQKDwkfNvKj93Kkof
qvQVGKHMOP1kKkePXED+gvLn/R4b+75yLSlGljR5tF8AEkL5bMERLPT43wurOfmF
tTJ+lK10ZwKbKll3yB5wV2AJeqMxX9E3MAXGwluw+eQ56jVsCSG4jzhWc/399kAz
AoxtJ81UNF8mSMoxKlIa9oULDO8e7CvbFjNjF0EvFvQrjZjiBF2CkC6ABHvZgrN3
mUDy7XMIVbjgcXW8oX8FCIw6NW2YYcQR/7opr6syfWF/z85nhAE25vksd6l7tztb
cVoCnu/laMFbUNTnaAxDRHQMPNLMbuNIq+/MfcJLOdBCVTnpu27vOOvcHBQaUoWK
ZjxFt0N4YMWBlXMyPGZePdmJH6mC9oAqITE3pcchRS1FOcUNEQEJ4sEbjfyriYbk
t5o4HBd0W/6OJFHt1JfRoA75cMdkaoPvO/3D/QPEQrLn/FTnMNGZue7iyMkb4IzP
XsibX+ikJ1aUpAu2SJzxyrdJTfZtcWceC585F8q+HSjx5Itv7yTQBF5I6LQPhOzs
iQuPBvdAtpHhBO+Qh7+LdZ3n92/JlDCKuGH1qhQ8+vy2FVwjFZgiuZqmnsEFBn04
JT61BE7fKxFqE5SMjl5So2MZwkV0qt6Jg8+wWhRf3+lDp92TTxgoVUh0LVzOfP+6
Cmxkjxttl7pz6G9/iKkiuuc6RcEEU1F3EsdzYdsOTxTOj/l0VPdM7m/53iZymZIu
bURY1lKMl9l8+2OHSqWqxgiG2P2hYZ97PUrtQYa+OaHdzxLyBAS5ntMycSOCf83V
jWsOuWLJAJ1UZlXlt6e31zRqRE2iUAxFtbMnoslMErjQ66+YiU4DV7bJues8JyxQ
976qtPZPEid0q9mDfh8BPc9P4SqTJCZIRLvsxC58Hd1L8Y8ukeixlLW6no6QVLk7
QnB/4MFR1jyav4rvJzuyWKSi7vY5GF5DJjJqsbKjbNs+kr1A/Hmn5/pwd1/0/zWh
ckH9TMqTer9ss+xYaoe5NO6o2/lAuNk3Qy8l41yS/M+Ww+VvKSVE5o0KW/e3H86c
7nCu4Dm3YzC9Qn+Hk11ma7iD+byar62OlSHy+ZXQP04ClwhMB01yIoy8Fx9tKJEK
mkOVGHgaa+Q+Qzdu6PWqZV27Zc4zIdxa5logVbPt211B4yMzLYkI+zMNUxY4ipkp
0ZjNlwLJ88hUp5GU0KkD7RM4Z7xYTX9PV82QEpOb4ZkX1y9vaQf7W0Xv+ZwoYEkx
q1Bz6ps+4VYwSQS6lzKKgCjfitA1u4DZ2PqzEsheM+Tbu1sDdOi65gYBWb/WIKFT
DHM+gZbOEqSaw95DeoHPIyTMpIw8yuPuo0hVpKpbi50641nvjzOArhszktsZGCRi
FwWOkGA3JaozvWet4gMnuU6/UkNUsJlG+9OvEm1XJx5epvDZhwcX9bYkmo2J1QRQ
eewpK3V4cB4dgob0yXpcZlrK/cVlFbdeo+V4yoE7T5dVwSHaTok1cWhrvfPDT3Tt
BZOdhVVYSd7YbJ5KCMw3FOKqvTUYEEmK+I84QZjKIo1wrYSKzjrdvrj04kuLm4H+
4d8DdkoGpnyOvoANABPB+Ig45Aqc/8Lyf5b25+vgQ2uWu8/HzlB7ItgQZ3Q58w+5
yRVPL71vbxVtA1o4D445H2sfQm56NhXNlj76TksdulNPmjvwSC3eEe1r4EIAA1cF
iSeveJhe66mFZbobFp9s1JgFrjkw7YY9plnpaRNpG+pGGiJaTVSikZ0gkfVoP1U9
SrlZ/vf2lFq2QmyxG9eqd5uUomsVzLwSS+7A6xUNhDaEpNCqGBs1qEaGDV60wWbk
hlwTrpuzX45v1JjCiUzX/XTER7CxVFevuXdTO7DvzVfxsbP6sDPsArUp6KRpLkc9
aqWsBFn7MN4IcX9FAshge0WIKTy5UvmVIfpEJmY35eyeliIP6mdCM8BxR3+nlymn
xuSz1fA4L5DFvb1JupAknkvGUlxwaw3pEwk3tBVhET4dKFAR9ebKlZoj/Bg7CVVT
qRllxRonxqgQFY34FGq77Iah+YC0e1UxFNsd6pGsr2PgGaVggQEE6Q5yNVCR3AQb
HgBNkKjwndW6VeFO1VHSOW9SkmtI/zstIgGeDwGfCSYMQx8i3m8Y4rA42f01RK7f
qSw7l25oPER65mL+pLsi3ga0s7a3C63xLV+VVUZeaG8bVi1yGzdm6/3CjbxXGFpS
AvfMKBIpy0co9vGG/fcLOGet2CP3Yt0IgVBdZhNhVh+wTniuCVtBKVgDFLoA60WB
fACU9aRzyRBwVxvqIUPzKrRPEx+VZp40lWsOXwa4ziv7cn1K5i1yBBTPC4BnVAiZ
uD2K0SE0UyebXj79cc/BoPqYbojb9UExrd+sphCNSquXnKoqphNrfDviNWEu4QXp
2TIrfaHX++TM4WR4lcN2ZjFx4DZGKU+5bxh/srOGjZ9Ic1lHZ4WM85sqZk++IHCs
KaV79C9EVu0tS4rBKzs6B7nWBsucFjQ6QYD1OB7URQNpOZPOZ4tGB6sYZnJZA/Rc
/xciiqMGObGAFR/CwYWxWQpTSnSV5rghtTzRfZcn8KW1D9b9P0e6BWDHh/o20T2L
++JO6+qtUOceY9rHNO8pYaJPH9ANIZgqDYWHQgwRzgcP8lV9rTUE9xbLLopyCsrq
W+GBgpma+9QEaYYyS2iZDoiCRT75lRrIC2s4s84zfP/Ix7vSZi8vNZKKRcuGzu0Q
A2BLgIvSy4+nd2fgzlEPBB/USeZRkt9QMmb4/CaMnI986KnFKZj7dV2N5a1Iqv6l
/roXPWJ4eIQZLgzGX+6iLMD3RWWejq4qB8Q/WyfIf2tkyfaFUHaiPB0eaaZmlOlW
B1ZFdvu0iFMAkj7tatLqWX+B54IpZweFvjZpmXPBP3Y0tIDlC5DWpU0ids3rtruQ
cR4fBtls27XmuY2aTDOKOh2j74dpUqFtGfWvok0/Gppiqi9zJYISPrDHuMp2C4ZZ
3w0h5b5YYlmOyQ4+T+7E8cJBxeXad8TMdMX0/6+w0oe/69kLHUoyDkzWJj3K1LHn
naltIz8K+Nnqo5yJS9lS/Ts5FJwbB/hK7hmEG4KZALQFSWMnG9/sXnzJUtBXzIBv
m301v7nMR0hrcViJc8+XRX2KODxXAx7y+/dCitb4oefUG/dK8894tjvzyWYAGYqb
OlXCjgD8N2g9dMe3uCPuWCpQJZ+C+tcbBAlc5LAGmqoL+dXWYHpULIEfQwuY7ILT
flJJXf7pzKEvQuctRzGBDwKC3RimW0kFL14QaWy0AA4/lQ1LOKwCqIncFhrxGS16
cP2jcXD1T0+z+5LAf6H6Q7ib42exZvTmnaSeZwfcHsQNnOYJT1py9olPIVRTmIYK
aeQkMU1q/Sc4eiY94KKa1nNkpP96VA/Awo70FQxgMjlyKLOdoJ9SJZa2pUsOPMh4
CXAZufoLHuJnrUnKLzZ1D1Be1gmfiOecwrUepqs4NgMzu+yoBhdJS2zThKQJcn1g
+HFj5cILXexB1NdIfu1Jh+7kXIRTYkk0QWF++yw0PBVk7xJvL6eFrS8Yoka8sacD
ektbmKkivYREe4KVPALNcifhzgEXvEILuFEQVDGaaqkRqxtLYjOgQRmYhyD9OSLh
IDKmh5ymbhd2wwFThXovnCsfSS0MWMP+DG9x7OpO0WvJ+7TiCaTJ9x0I+eHYusrg
i5I1/URypvWcY1Y+HDAiluu9GAZgxor1rzgODdIYLKeu6SZ18J5u9mT5Rh2ZseRk
O14M4PEjsGRwO2uac/dQdFTRiGquIfCuDF+QUWWfpfnJJoYzKjxrpAsy1gbr75er
qwfG1c4cVIhGsSxwwr4InRVJ9I3i72jtB6PhvVBtusvH/kDbPnLwNsju8xKzAKGl
5NkVJubAaYRHmsZdvkF+q4QriKFeTCG0/ZxPbLBgKKqALUFEytHbQ9DUE7/gKgV3
UCQDPtbUle0KXRDsR3FqjsRkHDaOC/2XbTIyqLdacqCLYiMhsVt4VZNvFgsaw3gC
8hKoa8Jjo95emFMpjI0ddmOUoUQA4RTAQb6VFUqICugJUFy1Buag/18c9GQsL2m8
NGIcmBY+6N/GAyXKyini+Se1ixFKve70wv6W4KvpAzyYRHOEC5jydnlHj95vUg/R
4v4OpIm/3qKsxSxSX5stYUSn+TSgCy4qu6CD1XijjP5e10i42BFU/h0NuzxHH9+b
SZSu+sL0W+z5GeLFaW0Y50rsu/iZ9RNaVOgbC+EHvGpMd6JXL9qjNHMbhx/AY+ux
S1986PDSGRI+AIUOKfVF/SBEdX3e4HLlJXWfFHSTe+SCz0ujxlDB8Hnu43ibvP5Q
sR3Hjz/6IDZ9ZdI456PGiZYy9c3hIAPk51cDiFaNA2CUW02k83IITdr4jHU/ewM1
upmCWSydfV4NgrZMmQ1SClEBkHLdBHKSq4kQWFHyh1KzTybX42uFelZz3M0SZ97R
/uvCeGLGCinjrd5+1stgdepfGBK9aRIhf/aXt08jFUV1cLnMfWI9pe8fFJ8LDP2e
wONTQjAgvoW4Y/NGzMQlYc9sdOzw86+ttWsI0Tz5L3wDqYDZEYzpNwAbPWviwrFa
YMJoPy/K3iXe4kxKCl2JlPhEfWNa0oKJOkjLvKxS1e+lZXcndocp+2yO1g10yjSQ
g2IWwdD6CiShpWik93YU4v+Z84mg5FZ0gRmlICAIMvEq/aaK7F4WQMLnKclrfvkd
raI5EWpZUYKGnXsMiU+0kaM3+izc5/zoB/HInf4RX34rs3C3qZmqJ7CH2A2043H5
F7iMKhuMDE/x7vrZBrNSuhBntbJSNRtqsXvAkYZxAAauv8CbwnrTKPN8lSEtDzvF
Ao3zFnZ56AuFPP2XF9fSRmj1/x2MvB5r8sEluweBVHf9hnyN+rL1xl5tT1RO2KV+
9TvL9Y/lLJB/K1BqqNlqkkqByn0iGu5MUHwZoWIEiiwuj4GJJrTEl8n9WHjTlVwc
ty5VHA8H8qNxANQqwGDC1xbI3iEhA6yZPigPObDMf1kGImn3FCO6Org2D+X3zMUd
b17VlE3nf/zmHmt2JE/tkzfWAwDqY1f52RRg5APkgMANKNv6j8QCArC5kEm0dT9U
juCypBJw92bW2cv8QWBIYUl5sf1rOMg0VmNWiLLbF+QtfehiV6LmPnRcDbK2wVIj
/gemj32pzQrnPtW7S4v3ueqnPHZ+yPafTa5pYoO2dCffTQE/fMrMn4VH1leK8sl1
Ckh5ReAmJ/59feCFqLbf8PEYjqZ4/8Zt99+H/GDCbta1noS27rGDRUEewXg7QHFp
dsUxErodweJR5cl4/6tbJeXQOYKfHY34EVinNfi1SMr8O5f+K8OiTlE0BGHUaLoo
KrRYIrLhJPo8/9BRlD8MXtXGIoBc+BiXeQy4mlpLTR5xDvzcRpUQsGP2yKg05lGV
JMU7eWT9RhipFH3myuIey6aaifWxXQkU0zT6RPwUDitzVJ3E7m9FQBvgtzI0kUow
3I8U8xLLxJVQpU2EW53lyrT/V6irEVVeCKCADJQxtTUyFzZ9s+t41BTKEq/qkM3/
ojA/wW1Vsr/16f3m/xQd8SbiHxR8BAV7HIIceEfpi9F28GSY7h5+ElfqpoQJzNHt
h3jC8TJP/XOQALqNF8yl7vlmBV94ODmbj9LgF9PI8cf7eUwAYgcB8le5655fViZQ
62/79NumkqmgLkpNUNd2U/lW/mJjB3y94sMt+u6hZRuczvlqMPl5AktovBfZ8895
n3cNLpSFSaI4eU46NHIt/s3AyV+Rmmd7sQEi8froLfpP3eaZpBB66OnOALJusoUz
7z+xV1gcoXZmqKSHM4l3BO0kPnJzcH+wOBLDRSOgolqB7kzj6Q1DhnpNdzr7ipAj
b0anEQcpQ/oIMd7ipXj4n+lVsZODR9015F+ffiID6IYhxid4/n1fVZZf4yRAbWLP
/8fYtVIhj8BBtNxaD3WCVqUslLnJ7LzCsLZjoHjHl8u/TxosTev6R4zrQHIYrHXk
8j5hovon66UQ/MiCKNCXcokpLNz5M79XTp/ssQn+mbAkq65hejlktIuwjl42XRHh
nR6d323H7xoOPGy1VTkGG/1kH9intYsYAmYaBJSbFUNAtVndq6iuRjun4igNYDJC
r3iGd3bBtFms4IdwXRn7c4wjipV9Qd5Jro0hemtjpl0u94CUrGem0boEjul0nerp
Q252Jw2H26bs7HvqPpqMdXapQgKgQVaa6gr8vd4QPbc7FqtNNQUSPYJRh1ktCoIn
frfRAaP92YIh5EYTiU79DsdGcPcvoIMJJjez4LGtXI79G7UAVz/e2aECe0tjNB6j
6huaS0JhqSmdoZHS3K+N2D0GJFV0sYwDxQ+50rtuUf3CpPXAKJgsFAiGmbqlyyCf
sBPWkXmHdrgEiBPmJlT3Hsx0KlL+wQHH0kqt+7GpXFgIZmRJvxHCBokNpC9Z2V2J
o2uUrMujdmAi31bDn8jzevPqMmu2ACVHS0nlsA5Pc6u+NyX/aeVRKct2oCZTVlA0
TCheMtyDDZO+xymN3lEDP+g28cQXIheG6H9SCYnRHIfot0kHbN0bLSnc/enxt6Zm
gh0/e1jtPgw28Tuqv3OOwsQs5b8wFrLMkS3n/z4TVWraWEvKfP0ywmKLfeT1XnVW
KtH/etBYN7o4yAOVJ9ueZhkNtnEwfepy1QZpZ8ee/EvCgkybI+oEZaD/WIn+Mn6X
IFAAhiWlNURYr1YbGhVai09xDki4oEdjRHwTgkXSuusVLuzgnbz/FiQiQ7Z9At7c
Rn++oyTrnFi9KV1RpaOq+3enoBajkA9VWPbpNJqZP/WM38D2wQ0WcayyBMf54Pp3
d1hRxgQFnrsI2j4wz/NQEZJtStYuyym3J6VGQukYJLpNcd/EdWANbog1gRUthaei
1lZJ5RzEGYJs6QAP/JRgiUoCfTPNBvHI/umV8dO5UtzdkzI2pz+EYUmN6RYN0zK8
B5fCBO5YFTO8N1hE/32i8ZEApCyh8tACQVmI/To4eysja+RcXh6XJV+A0zkP+S+C
lQ55fgW/4rBpPdl61jM4Sc3iKFGpMlFJ0B9UFazbutJVzpcGWfK7WOaNifQ9UTdp
BctubTzZaZ0BSnhAk/9G/8YWmoXZeaZfb73/EbdgIFkuaSOHi/w2i/XTXcRDxx1r
YKM6w+c/oAYmZBkgvOyLunAbcPiRVWTL8xU5zfwbcTRL5bMoR6l1jvQ5vIKkUVt7
i/mVFm4+2D1IBiGCM0jP43Pqp1hY4TLK1MribsAHGW22xN6+4ulYuVfuI1omVDDN
qFjtuFhhRJr0O3zDJz1qUdIJItWGTQUoeu1O3bpF/rG+Qu95FX914ZYkas/6K2cF
gAQ5baEw8DakSWRJAfwQM3axNzQZHiUfLs2h+1kLrolTue5ky5JJoSbbwEvkBiO9
FBr0PXgkO2NI4hzU/IgxDbDfduHme3GHm93OMtzTA5FJFr85iW4SuXIXwpBOXuss
K7aJNa0LOex1b2TUMhG4vxvhz9/VHfhqQZ2yPEJ4LluGXH5Y2vL4xwzHqUYeUsEl
oDo2oe92ZKasVPGLAZ+mXpOLMk0GcYJd7yw33BTseWI+R6ZiQhfcuBMd8fcnEVv8
KBcoVv5w10ysyHSmCiclKm1BTnY5UwwNdPKNazYYZrlerOWBuOC2hcOzSRlr+MAC
HSyhpNV5V51xpZvjksU8eL8iemo8tdHLpXdtIR04gsLXPhyhujKlrZckL9E0gPcP
yAeErBsa7X3hjKbI6jxvFOURjAfaKtDZyF3BROTLYv2nPe9Jh3VJBhZm/YZ9P2b4
zj+Videl6rLAWW7RfhqUHznY1ElP2z9pP1U8bP6jNC4FJHUh3Y0PC3HpGwch8yfc
vLqyGe9RZznjm/KjvEr9xpFf/OKlhl+AmfEjTD2rTYg0pr5DqkcXqDWsLNmOf/HG
z7aROuwC8cgvo6q9a0eX0DGP5Ffm3gKCC2qN+sraZRaKkFMBwgfd0OsB8ybjb+WJ
UEY2O/mFf/1H15CJohVDUboRZ3bDP0yvDu/KA2x+OUUDagzLXmJu8FL+bnCur7AF
KnHRW+AgiAy0IKsepUGrInF3xnkf+L1a6G8i4SWpZn97cVQJtacsm5ffUJO7pZpj
i+V3OENAWvWGhu65qSw0Cw0fLENgUX1mNf5V2t8Uzx3fVGVIGJMtJXZbmiR+RBCB
yWdHCMOdZVluMVCEgA5zLRz2UVcXY3kI+we+8PzS6SBM4rFa5B2o2AsAKIcVBFNr
Ch2xeXIvY8xdkTimuwOFkPWKLyYas8T7Km+wjlA3d87QqUAT7E4v3Frevciwv+6X
1fOaDAAp05hcteLHGGkWC8ABeFEY6XlBCSjr4qN91qeXDv58bJ4RVFsRAzavfIX9
anfJliigFkGE5FoYqlyzYOPaXlWAdhcDeRjSAVCsBO3FYW7BzgZ80a46l9HJ8RQf
ybg/D1lfuHBH3AIJjGL4qJCgCjb9kBqZiZB7fSRklrqHjnaK3JmfK2axr4vbhdRO
S1biwqi3xHo1PQsTOnekyQoGEpg6LDiUyW23tLVzEiZbWkEy0LpTAJYchHR47c5/
VDNKNmWXu+YrxdwAWeSBfVN5Ur566JqGNnplwbwbHPdRCKlNimZ38KvxcpPNVAa+
tzkRvV1BWihCtCwcL8JrXapQ10VjWn3ufX++oeTwAX9rUTJeqKb2idxPo4qZlnas
bCyw9XfoWxOBPpcQlW5FBi8f6j7ginLHZSBzu1LPVABrZiuYAg75hmxIhK74Ud3G
hfL3G66JFDUZKM8KMgXSy7yB7jxy+//GlPUWKngytoMbOc/xcue178offAGrp6Gu
AFlVlOkyKtin9zuTCo+wjrkE90U6+RtS//o+k9lGyNWjVNOHLSCLPSQveQgXHK6M
pzlaanUmNhFilU52hqJQTV6HICENIUrTQMWS1whZoPBMGoDm1Lp3UhI3TOkCW9iX
YGSmGw1+dArWixwdACrnvnbFBionapuZ88cE3LpVC9TCcXz7azPtFSmq7Ryj8fhD
u/wxLX1uUSnDo7eC3Zlx61KuCw4QDHngiLoXhsXwFf0ImoIc5F8liaedHwmQ7Upn
FoKfgjLxH6gDINKYxhrK6kjj0ocJ/NJswglyTH8uh/W8UFMKJBd0Hsvm7xHWE0WN
Fv6CzOunj45fZqelvozBm4XlIiBfcKPjZms6D+WnjTKcOf3Z2+/MYOndtbRYs6C5
XIZd1hCHtftT+agv3O01IuebDz9nqkJAFUzgK28g6xG7wUNRp+WE7ru/JcjeRl8P
/3F6eUUHOHidXYJe2uQjXxWq7z1gWF/Uzfj6nRX0EQFjcgwzsCwb/dbz7H5Imdcy
NCiWA+T/1CAiilznQSIVTj+r9PvCdCuhZdcSGNpYHkRL67LjU5V3lx3NEcO5x8N9
LxqsS5MqfrWTjqLitJWaqTbmV0b0zDU8EH7oL6sZTi8D3jdxSsGrq49dS/rNPYYW
3JSDlAWRaWj62snp3E8qZMEbaiKR+can7SHRugEgtPwU0W5JuYhCWelK1/AUuv4X
pPsvfacFK2H9f6vBnSWlAAi614NDsLZUvgu+fBxJXz8wjJP6kah7TnvpU3cQRm8d
VgPrwHCSXIHOAD7VichWT01jjvVlRdRS86J86H5WlKIfugb4vFvIDCsk9gFZGMtx
jUMtOHW7UYOwF2tz6ySpn8DuhXnlztkCwsQPrmkgSXKBojThHlMsGbSQWD0Dcw0k
Wyh5LMlb+ImdHQ1i8gc1uK9AE7XbyE1jRt/XZocevnvY01EKOuyqefoOQ+fM6l8g
9RFKONbi60ISD5iCF9brAPjjavhIFeCxcSoT3J1y077/+NY1Q5cLTGnUxV0Wm+RD
tXS2/AuqHYV86I6o2I4ztxy66pTj8nEOvpiM89WuJs8vxIEEgJOsSt6CPiiS2kLF
MXKApScMed1V6ZCY8iC6ebEufkTo9xOaif0aF6CkUGkbPLT+mB2pGKNKXqvJsQ2G
9qlP4CxBHCyg5VsDmiWIK0HYlMLRDV0/Ars94hd5EXE3FB/lzAhXAUWsR/IAbtLf
nNc9UM6jNlT08SZ2xJ632uOfPsms+6/+gjMhCdjOtv8itx2UVKn9hifEWK6kHoAz
yQ2WEsBhrnW8eKJb+yLoEveeq2bHGEeebt3/BZVbvSa4BZw3Sykn2hByaxrpJX0D
PC1H2B8r5yCaa1ARQfLiqsJG0ElkZBJvV0Aw42dd057ix2IMfv3QVwlqvDe3ygYO
/mBrUD9MAFJnp+AZpNlwHFJJsSyCB7l3pepnNtx4aDOxBhfX0XwlFroD9htnEUaG
o5/mhopJxMoegAs1uoXO4ERsPOx//IVVFreyzrQWD943wY14iQCCNbpBgCdAwlAd
4eGw7/TjsxBb+1FVsGBOThDRHNQFIb3MRQJ/Ihjfi+sS8LBm0YLiuL4oMQs6Bzr1
unHazr/V1MrEWooyiUkH/XQwMmMdKhvrBfODi9jG3Z7BpcEghzt1S0Zxuus9oUvb
fBvnhCHo1j6GbegIOg8FWOXJdJAi6+t+qriPQb5IHVCcnmkJwuHnCItY6pi5NS8i
fkUrwebuAh5hxMto6eMv2qzhytXoHwjB9Mru8qr/lsD0UBRK8ss1WElH0LKCP8dJ
4X5g95xKAiY5S2dmy64Ms/AcACdnaTwllQ2rGNAVFpCS7mxOl8ArB9pl2NBQf6Is
bvMmeY9pX7SABWLMe5XswYvaf0Kvmm692ZRhswGnk5Q9tso1AqzPD4TdyOIz+Obf
LxuP+3uun+DtKwfTzp+zEOzjU+lCWm2bvpYbEu3Zcb3n5Pu2Eh1On1iZQE+4UrMk
qjGWOF4ZyWKWm4lH4sgACClf8t0Twn7Vh4chdPr09SmKoZqbTrmpl6NDWWk+kyGP
TJJm+yV0ksGiaYxys6NQ+VZlpA8RPJznQo8w1IZiiQqvN0H741Ak/ynrfRHR0pxS
5D4+UwIX3j9S+S+2iAWm4ATB2MdIcVcnOFUtA9pB4U/sN8Xvpt6m/+uRku4UFBrG
VFNByNdJHh1negrC4Gj+0thyMVRbAQEaupNzK/rzHWxrE+zTUsQ10N/4nuar+A9X
rbkX0vQTFy9dkUU+eQICimFVYnIguLjGbsd+Ty0GxQIKwjWgn/9Jq3JLs1UdPK3c
r2X3PlKGDSadqADmvrJejvlymI+XXyXR1eBKmWSfjhCmXWxQXFGCGNGer4WwqiIH
dncC5iKu/Kq/TUqhw/PUIbfWIKYOpijrXsEbZwtoHwWG0QUeUd38oFJHb5f5eBev
aGzf327KzhSxsobXrSkLdjAx3cSNmgKrGSvzZxj7urPIP8K4+UQh5OaOkJQHJB2o
0jy85j77g+/EDElPkkD78QrE8XkaFUVWDa2prKp08+Fp75nxuJlAYsqTqCb29SzC
k9Bibl0w3I7aLcTwShYo0VDpT0GO7XqE1julq+VkJQ10B4gXzefZOHokyzsqTdUE
Sh91CgxtkPUySXjt63jZStqAjhA8xg32KDeVRfsBOBodZbCCIscCG2DcaHzqxzpX
pS8P/Pu1i3Y4Z2UrUdFLpMvp38ZMHayVhZ5qfNBbRNuHekXWjjQG5xMicfAKROxq
QQAyB5r6gq1BgaQFVIEaB4MnsEavcJhB0yhc06g1VOpoxi7uCTgGsIDhHDjYUG1z
DAzn5ktcHNXwHW3KH8jAuOilte/9yCAZLY2khx3tQ39teefgdhcipLKuq7eYEXAb
2Pi9tfPeQpbvoWuojvR1DAPfD6F/q5H6xMY7XHk5/rL3Gcqt6PtaRfaOeG/QbZVx
n6RWMEfUiZZSmVBSS2x2wWKKZyvLa14WOwUP86lBN48jUzGPy+Y3WjCR67DshE/g
6OpZR7xCKWLgHAbXGVrfqj6ioZv6j4wEsirM2PqqOL+h/qJs1bVwq0m+6tXFh1yS
H1bomGB4zbC1NOQpk14/370kmgwYuYp6DPqBAXIggOfeiHj3zgFIeOXyO44y+gjA
yR7480I0BoyfwevZOAPw3FVj9F3jv9/yZfr/hd1RoAqGcWm3+EjLlhOFz2WwSxuE
zkTG/WajFtNvgxlKthNPLFp6KOxjbroLr5VoXCfx0QFA3WTchXhfnDBSXgCYyZuk
pHwHbe+oXwEkmxPB4ZLd6pe4MKkrVt6qggeOh1tShGaUSHddkrDcJrDE939k9ula
s4abkSBRWguK3f2E8fRKLZDVJuYk8Wjlv+vr0FY1MdmV56TVFUeIG/smpfMapZac
D4cOedO6SyPR5SCSb7ojdmBpyl8FfSAk/Va5etdpYJUkwZiy88b9D6SP15S7A0SO
DEzxfUqUsp1I0uJzkqO/hnyfRm6VitmyerG8BEwGRG0zRK/Fz/rZ4u06Wnwo3BLt
ItAWG6eS9B6kdVHNNGz36LoZmEn89Z4zOARXwRumGNFe18QEdTcJOdTn/DaZlr2C
ncy0Ld16Vexokf/mXeYGzqmeTW0z8aY7BDJ2PNq0ZAfukLpbu9LyhQ2sLstQmMYD
wXh2D1zBWHq6hMg29DAJ7Wy9Ic2yp/y+VaEAzHy+Hxch/xIKcvOvZlgtC6olLXGF
ydQNn5pvAzQbmDh7F0Sw7xdT20zgtzMz1HqOnCePzXqEWuLBiAojCakeFQVH+sgI
SL59H1v+DaFCDlvGyP+FzzwAKzOIZcjVdGlOfhnxGG2MjUMwjiWXkavKDE/vVuU7
3dj/xa8K+RGFsIStdi5OQKGJrZ5WdFsMqKrf1Kmwi65zsH4cpo4VNdBJlX7APeDM
ib/NQ4Ty9XRrfDcz8mXVPgfg4ehAe2xpdjXfWphUyuHM7lCwSpn31HbK0FUYM0Mh
uYisefvFIdiW+pSk7WdquElGXlP98/WxlZK1nkWWMyeC2HM2bv45TGHn4MH+EVHa
hRrWrTf+I81fimPLlq90Jkj19Vc7c7mtToo0rM4Pyg6S8tQowD5iQ++ncPSPvS5S
YqnOjyvB8ayKNQVdd7VJBPvW0UGwrkOGYThLsVXDKEdG2pDtwnbuo1vEIPZVTLb8
VgFPFhC4TuTroGB07Lac02x1UV6GpzS16/0pnsfbVYL6K1FHY5gbkoXijMWcW7xD
lwOElRhbQovzqDw+H4HBbB3gzH67u9SCoG2uc4w1nOVTtyvNKkF3eoS6rgnmANBx
Pl/Jol4Gcd9pLtZ6/mgdiDt9u8BXzFsLRlZVSuf8oPpDnqFE2EYMsgxLxXxIZIb6
ym+yZ9PHMQomKml0cqEXGKoF2EH6FQwGtTlJSGUm2AlsbCpLcvcS3JMD8E+yiSPH
MwZu+fMt8+4ILqSKN/ZWr1Ia3/2og8uewh/uR7SvuAJcK4Rk+ofDfIkGmlDtXb4T
Gzi53mT33KdTZKktO15qtnUoRW8XyPI+RAWQiSI2lyOK0zCG6xdB0EdSJQdNC6eI
tfYwsjWrebZx3Wp9j7KL4HRoBQbAE2dSFRkYfS4sJTJGVyd2w6dbHdx48WYtAn4m
YSpSIKY0tEY7j1M/VulwCUghiPSZ65vdOvXZYGK+r7CT1xMNA2m40jNcVLtintQ7
aMF13HNY2/CisubF5ljq50cTGw5LWIK1KizTT2kAINSCIk1KgV0ogObUmSr4psyS
2DYSc2rmNT/wnsHyIvcXIGqI+ipCSQFoamNhZPBxNibYs+l1x1dQTejSQs3ZA5ni
+kLXMQU5ab1qLT9Jnpd5WK6vRp1ZUJO1OgUqb4X8v/BZ24jSSS9mTqvvrdmx/VsY
OPs/afDNrn7Bymmr3RZ2h9H+XH8IXE1yjVKMQ7w0BbpDw/V3F+kH2DLPjYhyqy8l
A5qmv0Qa6UB3C+K+VuRyYZ0LGzl1ONyVumZ7n1bQrdcfCWVETYzwVFBIDCsxTlMC
kiA6aIABtYv5XuzvGhE5CKRfTBggCB0OpBNSuxUITPaaZGn+ncdp1CRUt6bYo1QD
8xTaxHTEL1TCmDwwh5STJjh30nu5SNqIH/V17nNImDPl/p2rcX+1Ep7415IhrFeG
63/bRuW29sBZwDx9fo1Eqz/xyT9K17ih0sc6BoXbl7X4DXVe7lXnnMPgrW2xS79E
CtNo0qnntgZztM50MDzNe1FCAZfld+kKQE9suqS/da7e8aDqT+E8b6b7nV3M9rli
0RrA7IljZbQl0VZj8tS8i0SGrMc66euzEpy9kCQ4BJIdTzI6W/nR6eBb5HCoLaJR
SwIUwaM8wx45smGe10ftFeYWHi2yAUbUjPBtTxSWtc581lN2MDQWKKKQ1da0YJOd
CIjCRzy/ylqGDuoM9sF2WTxpth7KhoLUfa11XBoquqtVjJDneh78Lya09zhIfgyg
Y/pTBHsHFZzK2SAFcUmtfBGPJfobZMq+Hq8pE5ksuohRnAD80X0yC6GbvkyssUYl
oPZdWAeDQPP8L4XucRTuMPKcIwQB+CcNcuaixsN2Mzywf8uSYcURK2mHzQqtG3kA
k7UNaY0UMn0rnr9h9030hc4LtNhoRvCrx7tcuKnQmWGcJR+jXOBmLRXfib2A6ez2
CKJn7944qKXoZkPYmzsafhMRb2rbtf4PmVfRuEnZMyAfzIJQIAvnMOMLhXTdT0mh
oNwPPVIckXCc9N/10Mz/0ZbRuKEIOifkRRQ5veWS7sdwcM0r6Hd3DS/N0xWbDjcn
E5Szl8AWHeTNcOy/RQqKd7iTKGMRZhtvxMEaCIbA+ec/R804GCxLMbGM03XfTm3o
OOUVCuI15KTV70FKpg9W/tinR5CCkisT/2A9YLV4Yul8wmH3fErD4wE35Z+EvBOO
y4Eo9a8dHevHwEAsX3Vn4kQ0hjwVM3dKPp4De8F4/lzuvhg3LLN7nSluY1zNfK8O
NXB/fTO9EkicULdBCOmUVAVPOiUGV5NuXIbuD6pFma5BkovjMGI3Mzg4NbsjK4Yf
N3dXP1Ou3SOaQ+dWdAQdyAjK69rvt+HelU8d/WyadiP6G5Ts91IMpy+3Yoz11DHf
nTsIMMvaGYs5DTHT6QWVHNrateNJy0F3LX2dyI795F8y4b3SBF7LPONzYilzjf5C
ZSK8bJ/rOljW/b+uDsKtbxdPsiSRQariuy4RV8F3lVJbHL9173ZKj5/uTC61aNBl
A/ML+k8S/G2+FjbZTrlPzcnqmr7SsCOx9iay83FkU5y7sckgHnwN/wQ/0/za3kfa
gIZgK8EDhUajwwpG8cudhFk75Ee2e3ycMKAO/FbblRhDklnj/20TGtImT9zJMj8h
j0PtilKQFxkxBiL9vJ8iAwDXu3hHaxvD4ZDj2MQvKMbHMkw5wKYjHVaY8Ki/vpjv
DTWnLUzE8U8O1MHSf/MZCAOQDHL+utAiulDwEJs3lz43k0yCuNKE0Wjd7oFAvI7E
ZcHtaPlVnC9ZTjn7n7qriWtsl4/xh12g4YsGtgUlLciOwt2LqUriPo1qdoBhctWK
GYKBjQxEn58CI+kz/mDJYD/0KPjurNMZ2gkAPKd/SkXnCUWn2zd9tiixkKzuz67V
U4hvBMY5NXPisXmLzCqeRo5Ep9LRrnmQrwr4oGxoBj9ISJvrtPOBi1K19GkhjEtP
CxxKGu/42KgZf2jcQn4OCbJr2YASa4FbGrXL5wFn3KeEO+kfid3BY+wNt3IWifEx
1FW008tpE5VD1t/y00Bc4/mt786fQ0ZiIF+nKOL/VndlAFIoEyb7WvirINYSXyJV
RBrv8vpX7T8mASygVznxvvRXl9EjrsaF4pkoffG06wPltVbDFeqfaAQF/PLrCASe
Boagy6uoL7xb7MTGS42VKXUQLsoBQa7jT/V2O2VjOW0UUXr/PtbaZUImmtpHq2H9
EVJmNl9gveGuISlmirVFx5AS/azc53P9r66G/He90haD7pYTwjvms0A9G3TgvtIg
eUPnlhK7S4ErDTSOLsE/OZRj0vMod434mfIfAj6KAysX5QAKOUxPbLOoZwKAMW0w
K0nnqgYl1twE2RyYCv2UfkDnEafJl5h8bWadmrXjPe8YPRGbL7KaYU5znWh89Ovn
TFTwUpnsOST8jTgREcB3uWTdhLSzkfbX5bDRX58/80wXlwAh0vz1kDonFACQx5Gp
vOJmM4EDa8N0bNE2CEtleG6zrF2hmwVi0/i9oAQA+nywtA3JLq7/W0qC9toQwyB/
KMD8bCQ4Ttmp5Cd1fZhJpNGfrYoDEJslSi80WUO9yNsPAeW6k/P152DYbyiCZ/x0
xbb08t5VFcY36jxMqetRLqOcgeIQm6gEywoPclQxf84oQVzq4lv9lrHqm0tQZJau
KHZysuyo3MfUyMB+J8hqG7zf5zZ+6PVZKaZLIK4lJyQz0P1cji/BxnESEz41CwoQ
OEKrz92D8pguLQS6BAKSZ084s/GDohc43yA2Eb5SgJFvUVzoglyaVR9aO1RAC08G
xAF/8NegcBg00xbL72tLI1hN+uLAQlRkaaCRk7qpO7Cn3nsSjgal0ZsldJKYWMF2
NOHl/jf2Y4wpvrvhAlLosGzl1cNuOcTEvLhHXB/Ad/v+7pJ2J4aq6ubdjIzFZ17J
T4jzltez9UfBOCHnJzD9ofiJX6Knye9uFa8iWCS9e074zM4ZJq7MgbARHNijzzf3
3KOzSrEXs/XZZKL3MgflbeP7e++ssiCqIutZkU8KGyxuJ2khdeuyr87deqo7jWE/
Xe0JEFPhlG+k8/WaTxNc5Tm8TTKU3N+c6Fcj2iFpP4mg+krIMhetfyUtOcJ1Z98R
4b3ue5TJrGYoMOj6owkGRoQiRyWWABhPpKzAFwOiDGVSeYGg1i8qg+f4H/9QjBsC
0Mex0egA2csyHSBQ5DF1EAUMQJEqp8EdT11yOz0YZ5hg/2xYqUvIxu+Mb31vlx2v
Wl913bcMt5mMxufLX4BGRWhCllXHfgkLJMFqr39KpTcF1FCicmgu2wR1VUJRkL66
ZMPgA4SecEwneSKC1WsVmGeeT4RkYsqMNntG8hRia/+sWwa9rsxUilIZNmcJMZYU
hbR/phdt958ENBHthu1H0rHTcuDGYjuR4f+6SiGPeDBDijpUjf2rKDcDfGDLvc4W
+n/aOcF++5nQ6tALO8co7jAVD3l6bbT0rjDPnPoz27scCqcR1Q1jjraU0+8CcPpi
Y46WvgXCk/oQoytbxtUfKtAfqx3caNISb48ZKkrTaIuCSmr8W3B8i9V6VWBED6RH
TTjuvom+XqXks1UTHU/BW9gdUg5j7WEJCLY0j5w8LeJf09c0bljS3IM6V0/wWUAn
yBsPZnbUC2STpXVizXhqxVX9N/kwKWbf/2l8ZR7/fedAAJYxBZuUOms8O1mHvhCl
RA5BrRZIJqGJiY8EQn2c7bZe6Kd/tWE/FdY6fkbTgUQvSG+ADSKMoyEfFN1DPqTT
5qbQWW2h5AXF/gAB7vY2hi3LF5i0sHCkhY6aqKTMwRysDoJeOsDCSk+/DpPG24u/
tcykl2aZS6DSsCqQKlCVX6b/F/3aeVqSD0J87SK2yDAsc36J+Fti+3qmkb7p6zCL
Zqy2YyqdntQGLNTgy0X3C4uJmNUtoYX44NbM6vj+iP1dyn3bYPRoYTWGA3/3LDSu
peJ/j2Um1x25g+SGkb3KCH3Pk+9jdj+iLsoxlrHICxDiJQqNF57m9CD7B0RzAt0B
raPBcjPiNVRQ9eMy2Yqq5okGcRKZKfLxrC3Qk433FzbKizDjAZpy2gEbeoMEGozN
Uq+JATDl61aYmEgXgs+2iPXqiteObQgttNdImQsNpYRcGISjEQ/xgp94jb5XLlgc
BxzrQxwMvxLURxfuhriPu3PtSUDyf+Mf56jKckdMAokCis/ahGPt4OpdsE0XjUd6
JuZB2NQaa9R+VF/m9TdoHHXZpSFH5rPOGdfuVOMx4OYPENj171652JfKVwkuPGuJ
w/sI6mFZNJQKBzRYuf/TjGJohiSctW2t/Um7CtaMjyiLu1H+D5uRgEGhf6tHvXxp
vSuR/wEwDek0lRdh3CGKDDmqj5X/IIbAuPO+R8BQbkAqM3GC2HaRdY6LDZ2xmWNC
x8r02Kwv0slPgRPUApkZaW8h6W4ntf/dhptdtW73OebuZXRoIX+RF3kw3rOfOGSB
EXTSbgaTKNILGo72m9zqaFDbUoUytf6iO/qZaDBYdo0EG4o+HWArJ22DqSKqbr6w
CSP7/44PMXPNesHsgwMCNEH1m8V7gqCOsZpwOvNzBog27OHa+h4mlT7DqOwhXeP5
sj2R6R7i1PO+Puudw+LFmXEs/gZ+SZ/VNYYK8aJQ/XWXJfDbtGVOs100ftqsLA8p
NnSF3p4Dq77IbvmQIVN7rnPRqU4W/4EwC5R32kcvNtji30o28bDHkwYSfj+zu41h
Fw43SbwQ0MNQ/bvvZIIIiBkq+Ev5wIdhd6MudIJarw28gzpzeDfhhfSSDifWymZ4
sSmhQdmb4ne7LgcMtXLYBFijUAMjJfhKKTVbgBCFKvgzE34L0bcKPHYSMNSlayHa
NSr/nWpsEfvoACk5EXVqH/wQ3sKEZkw3pKeLBBUs2ke4cQaoxdTRO3V/ACZ4LU66
nRM3mP0HNsTykFr3U3/A4phg0mLauLcgjdqfQok+uXfBaA8PPFnXNAZKkhTuOxAE
Qwfd5MC74hXCP3a39aXZ4G+mslExYPq8Cn2hp8DiP5oMfAiM79nChrY1vVRjtxye
W8XWxJ7mQLI4fW+AVgwlYO50Qh+ZaDmIn8JZ8lf0ito7oeqDj7RQJwMxAbeFlXZi
sKDmlrdFZdPmhUYnw7SVJKk8fLzbvZuD1eAu6fcoZ9KjcbfIjrRcJFtAAbnfbcy/
lpwY8a/Ksknwo0YPurCKVrU4OQS8EkrS16KlLECwykMPu0QQsvO5Ep7ZNfccwpXS
JqBZEjnlDzRBLYU8qCwY6OJ+3YNpdTXC1fVTBjuKK2W2kEdrLN579HAQlV7zOm/C
4H1a4FxC4HlDk3M5vdWKEqU6JITVUkcyc/ZnpGBLjqbnxOlsQhMXPvxuzLx0wdpv
dg0k/ArnSRXGPEWrjev4iqfXwLPZd1Ju5q8VlX19IzcUKVedgQsB8IHplOtnaLzB
dXBgAXSawEu2wH/Qi9SCPXw6sba4f09k/aJoXJchsZL9Br2LnOOOzqKvOIm0jjDE
X4nNsFvISgzfFuSRYabNqKyku/chLkXovPfsBnehZmnvHcg3ToU1EQfJ2Kg5TpLi
Y7CLZ4y8AUk4o7PlkEFkF9ASGUyEvOKa/2tqX75sya6heoTPzavCyMaLAQ6lZChM
wtUc/3FbcFkI6aRTfL95bDDTP5sI1s1YXUIas06F7yAQMFOKPd8fWk1evClUzkhV
S/IWoJ5EgHpuZ3MH2ZZqACfxIy2Fh41BgVUsHs0E3N94DR11G5J+mqL/O4rhrNJy
pzsnZDPJZLIRWkQakCKIDjihNh6rV/yIUCFKgVWuyGOUHmkzeJaz8s/yYt/M/oNJ
VlG6b1df5IhLdxwKDIgDNprfeFR94UlcCy6FHbQIt0KKi7Xpif9+eL5OQ8EgVEdC
JBw/bAHtjqUnhc1phNXnlMJAVXsXk5Usd7BVGdwR+J9XxApyBx5LYBxBhineMJUW
Zv1YuZsDhfTvdLgd+eB4lxI3YOCFnRzZJ59ErrG3GLu9K0GvL8RuB13uhIUS5YhF
dc/Cf//3EppUkOY63bpF61Dxzxn94f7gI+n6Ax5W7S7ePkI9GemstPdQ03ptq3Vq
vPwx7nRhmrBiv0susmI9Iqqas1jgmvKUHWaftWDLxJIfHQ4dQnf2EKYHyssmwJrh
ZBC5y3Mb6NZPzVHN84DQrrlmhXHKqTOLjeGz6jgYpIqt4KIvMn9zoRHnZWr0tBD0
1PX89PGDbJj0WlLtGjPUB7j8FM07fQx95b5Rz1hyXa4eRCb7PBYXcbPd1pfhHR5M
r/66jMmFL/F9Q/6gmuYHpnpqE3eOvI5a6L8JMpBm9VL2zdie7dhCMtxQHKxi7x71
QWpiI+ReDENzx69/JAiVnfhGI3lRD0hhIWtGV1eESR6Vq3aNJGAdiJUOSiG+a8ka
z2bKryVRnFrqLji1f7dm6Vf6RLg2gh9BzFlQ/QECyVjL7lBz/bQCz+F0hqpDw4T8
0Fpj87y+ONPrdZtKkGWdAfF5qrTR2p7jWiWIeJ478tWq+c5gXcozQ3CPKdEuPK4J
uP8K/2hiq8g5g4gLLZFyh9TX5Whrn5Y+hpqDTzx6zeDljj+8G28yK+m+Et3RNAtl
K6Z5fyQIaKBhwYKzST1c7b+9U+2XFvV8G4PspfbtYapEwtaiw68Bcvr9cbj+DTwn
puXKhNah/FGAMCPrNaHH6ieDqLziw092327oz2fwMt+yIGtlOukZOPWf9vtQsv9J
RVWMiW1r9tJy9RcdaLYGV7N+wcVKFA0QnRXoTNBqt2ugz1PXUN1pfKgR5ciqa+sl
pzrT8LtgQYuLN4J1Xtc/7lhJOzg2sdVCaeZwRi+S0Ebrm3Wb6lM/qTU1J96nee/1
6U7RzmzceWgitTZZLzGosS6s3b7RxAUN6adKgsmjdj6jJhzMz4MKxXgd2eeAzc7N
0yPKDC3yK7eSF9PlUPpD1Z/AEJIXnv/0otKi93O94bGbRNjT3YOsBrkoE/HxINCK
VJ/1aHDSX6ACRDc8tZ4Z/Wn1+uBiNccgmSGJQfaz1PQR66KCgqu4OZnZeQqFQG7R
mTsTNQ2itsO4QwLFgsMzoZEYUfspHiYHZX07csBDugOANnd117JkqX7dCtSVsyeb
VX8FatE3wsxQ5PcLCAc4AsM0FNZbGjBaJYZu+vhrOEQ0fgCWLY/+fGILTS7pUviT
q/j3lkdXSrgJQCO0jwr6Xi5XPfEOoTN6PJpaqP1Au5FP7ZQFuib89e11UwKuC1DN
qxRC8DVC8J8PXh9Uv1ofElsDK6N1FQBaoACB99aECBz1586iKwcqLpSdd7MBc/BB
QJHQBm9q9RZrp52bKr1WRIlPWNH/TYrCWInXyxmJa+MUGHrgmtFuvYDH7yQGFbfx
VWNHaUa8BVFUXgmiW3P7U5FVq2fTmTomaljvWI8Af6umK1zu8rFCHsREpTeF+4CQ
zvTXyj08hs3G4N79rJGh/hLQflWdkfV+7nWXKHaiB5ai/4t3UrgO91sMzA038UE9
pnntXjjhwT/4huiheapjtXMCAm2xOLPWhPi/9X0ruRqNSU467Y6ZwUuRdPunwIHn
d5JhDRoYbisQDdYwFV58D03/HAtzgt0P81NHuk/yGfSZDJpNeLmCD/FP1kb7f3c5
WfV0uKCLyef21balArMj0z2v3cD7AkSzAcjXrUCcZHepFoPTRMrnlRo9golQTxH2
YAKPozGsu3tSgswac3nOm6z6ZGO1AIiDTl1wqKchqu3VH41RWcMOoq08K1kkewqj
qMJbBHBY/zTAZJlyyQv60xbGq4eFeWDfuRWIyIIMn7TtFI67mqGqK+B7MPR163Fz
9U2fBqkSv6dtInmE1sIARru7drV+6jVsIxQKXHTjHVm2uGY+XbObWymF1cgAbTib
nQF8yZTpsIG29ilVSesfWSwpi7B3SgBxpLd+LbwTinXFaMmgx2i5VB6KRkKaRQP8
HasJ9mxD08iakTdLX+r2GWU9xhO5H/m7kL67kp0yNsZYOfDXkGjfj1FQX5UoiLc3
uSnS3KIXKzPSTP4SNsOBDv1i/I6h3PToSozdOxuerBdp4wjDDx05lW7+kyFGoarO
OZj+swV+f9T9cbdp49XxyeWBQghKODyCZ+CpPbZUEq0SYxeXoljtq0DtL/pkHwfv
cllnLKM6XVT3O92Ac3m9dqOXbpTukRrMqwidimO36AhENluMH1Meib6NnO14T57S
R51VrNSPowGfRhK2lEWEzLwzeKS9jIuQhHEDlHwnaSnrNHH0ko9/YUDDEMzFyaFC
OMvS4SOcOT8C8vTnlpQ0HHCJIHSZSPuL/AeXubaNTN1h0G8bVoIg6eVKTGlkz7NA
A0ngypwPrL/c5lxsODMhzX1cLX7FWiPm4GUYiG+gzZCjGVHchLp993NzUvTD2c9S
qXc4bNTBW37ho8XNILlIxZYYwUBlfTnQAuyBzKZH1gphghKng+Y7pY+7jtPzF8qr
jgKVEeoKmV2lGPewjwm3b7LQIrIZ21hWFByl4cgMsVODdubvQgeC7xbW2lQpaWZL
PClXTXx8GaKLfn+BIg1c7WhgIsForlQzPhbLVz9/ZlOoZ2ihUY/ENuRZghA4XPEc
KThWHCasZwoV+HgqupR5ntV3bg4TnhFR72qRcBpzsL7YqobEACxeWERd3zGgcxY6
G7+G/mhl/G15FP9J2mbW3WV4U8PXOx5Bl9BfCC/qYJOkzUnTjdG2+Y+aI0U1sTvn
426Bg1lljRJWQJtEis6K1QDNfPYR0D7VBe0LFBd90BHTRn6by2lPTU7GNH1V2tgG
Gphx5DjdKMRMiQJmdv1EfioC1NM6B7NZPy5sM3l+PBJkJZbPoX1bGWf6+HjxUExa
3W9n1YzVefP+R2jHYn9jxFUez8KA8621qnV9d16D/pChQH1smh8nEaHTZ+5xjWA4
HTB7LF2sqG4tVHkMeZymk+81DzLG378EhcrdtmYWycgpeLF2N3MsTqGN6zYOj3WL
GMIwvHtJZYpSBkz7ehYxQhgcubGTZXim504XPA1OJwO6OlB7Etd+BaRIlgJHhv+s
kCYg0yFDLyIzwblC0aRpiuy/yB/OSbMaN7mnvLTAUaj5JwAJx0AhML6JY1Z3KXFE
o8xBNtZcFMvXAJE5GPjRMBooUkwnFxQ9pEmPJUGFtgMqgjWPG0cz86YkTBNpuOlN
AvKQYMc3dQS28Uu3iXMiU73ExORHvN8Y5aNE1GTfwFpHozOBkINOMqyvZIeQVwoW
H11eoR+kRYdguwltznp9bmYym5fl2y+WfN2BkGW4UIi8w8T7pSocTq4P2pmKqoY4
IgiFfWmM3TeTpO6l1tN2kURG3gnwPWmXbMl07Kziy8MqOs5IJTQnGtahL2xGp/NS
9CUkLGcRr5LQzdrdJGrOT2Vzw9mQoAAcZAKmETahEGFym+TccyvGBA7YU4xqgoJZ
zrKISjd407E90jjZgnPWocfMOUu3d81a7+gpiaNHKAo/fN5j/Ql67N9St+bbol2W
srWyYg1K06wL3OEmcAp4rAOe4h4SwdTSIXn7X8ChIMRcRhjv0telXkWK8DmbqPcF
x68ZY+gW4AAgPK3DkswjcoSu4t22Vw/b9pxLluBXnhbHmxHGpwRswRoS+2SMUJU7
2SY3sqtagA16bEFNsi4D5LkRpqrNlja1y/hbyMnwYk9KYxJKe0Xoa8uM42j1kqeb
I9P4GrUKXYtFSUAFVPmb/cSsfLi9OTIGdt6CEImTHOMazZdFHpAoPPI/rC3eVCIf
wgdjUIpv3yZX8ndVQN8AvTYWMNqSPp8Ghdh+9sY4PYR1afyX7W6ZEYag4tv7Fpx4
kQnsLlx0R2NKVvQwvYGE8IOGXgYXSqzJYiw5WsTWizFwHiQBwNe64fZ9lo96MKAG
d+joZvIqM28eFA4HruQZVLSRdpJuPvCPdRUSFmNtmn85N1+H0lemFyFYGi6fy7gi
wvBAvOAsBLtyhnBWS/tqrtgTZbPGpFZ/aHFYLR26S2VznUSVjdYIsZKvMPX8ZQZV
wDdB66S6bxpq6meGWaAhWS14iQIBt2Jr0/5b44rA8BKUJ9p7gCQg4dNGi5RPMa+9
XX9dgCje7smlER1/k+DsfH8/PT3DnRym0/otNTQpgSm+dXV+ACqHXD8TBE4JB4G7
b/CseSLpB8Uwx2rDBHn5MHxrVg7u6r2vtlEp+7n6ZBclYHhimp0TMAWbgLLzMo+Z
AYW3Cb5okJn3US6vmBBnRTjd6jA8tRrlExdz41oz+4811XQdS+NlbX0jAEWCtdty
StWLB4Ihj3s7aj9w1nHFe700wCn+YqeS6H7pnTcjrmvhb2Gy2En7p0nm1yYATxKE
2+uncX4mNBZysO5uSQ5+O3xMvi4C1mYrKSNu0EkTvYSdjppdoVgKB7rL5x6hJwJd
AfeGgjLknBsyI13diGMXDP+A+myMnviMSXmEMbb8DV2+5lNQQALfnSdEqxQR1S5J
VOUB0thyGFE0klnKpAYOkEDqBrDljnjE3DH8LuP+dcFeUgCpEZeBb4zlCLWGelOc
iLtnScd6QOzlkpleytdPXoyQDfUyGUqOPxqZRycfzKIvYzTKsiN7JlWxUjDN9jFJ
sXlhtMa79Ume5XM/lot5qGpB+bnQRy7eYUOGS5+oYkxrdUKcFffWESokA3iII9mL
QZkhHEFFwGoODWcadXemvobx2lTl5/+W+LHlen3lGy/SrbxTZMoYTlqdZTf5zHEA
uo0mdVdVlC99eES6qZa13aAnODYdtLylHPIuy81Lpuaumr+p+VibeZRrxbXu3eFo
UWz6UAF9yM4Dcv2FjHoXe4OPrRPwxNN98yTkC27ye8x29HP6cf3HKkYvMd6+emGW
yqsf3H+uSyvwz8RtaP5KrU65v7fR6iyhNn6Fihetoz/CvaHWxkMxt0Ec9pAQ14u6
zlAvkHIaZvXz6MSyxnvvsZvVX6cp9oCYFkNarv7rVc49eFkiRnJ56q4omL0kfqox
TgeFwA68NJARU9KLcFvehK75Bqd3gmyMF82roYC0uF3UuY/WRJ5FY87sthv3M50g
QwOWm0tKWj6I/Sbo1qMjAY8UsuzId0CcdUFSEGsByHcGpdCsn7zUNnPUz8bJpkII
I8OBI1s4MBkwS3yntGvn9aqpZuxf5AY7uj6DxMu9oGrRIMmAFvMtF/nA0HQ4Oeub
uWzYpMMPr0XZZFH/aGPYdpspZMyJEHXBkE60QtLxd6O1PQYKTLrMedC5gvVRxkCr
3SL/kKX5eYyEMBP7A8c0WA3Ay1MO5SxBwwiS09LJhJ9KkdIzEHE7XRCsRNOaa4YO
h9Q2Be18YXJSJL+Mhl/P5UwyQ8gg1wqKuvuOsFejr4X3RKm5nQw1jCvsoJctUpZb
3bv2Ah4fqIAiPWh66+n+gfJJQvtFDWx08Eov+fLj5grPXyWV49uSv4+rYeRGOioX
6yh70wwpL4rvRhxUWsoYt9FVvpaLkD+32yeX9qlftCzeKnJi3WNwzD23rhdTo/0R
UySxSuDQLrgUWnr/mhdr3ttUzBeb6TmmE/5ej4t41cYiXGfgrbd5LkRCcL7fLl/Y
CLUvfT6+UnC+LuMGYPkhvnm5j1B1O6cpNolUeRDvlKUEjTHUPISMpx7sBBfn1MYd
BmcQ3H/0y6s5053CXEn5SU8GBLtLBMOe+t11vgRO9JVa2lhxuQxHLgB9gHg+/tiU
qtZrkDMs5MJpTyYBQjPyfK6zcdjgucZ3qF3v1whVafO3O++Vcjj6O42x7gHF4m3z
ZUHRhCxGu2VCPqmV0My/MifQQRxvn66L8T9mNPq+fEOSbWTn7qbj+BtNpCQWOTaR
cmQQCg0zYCGAJiSg3p1TrraBB0Ck6jX2swnJnSN8QEN4Vw2FsJMSgcKyr6PzpCZP
z+JqtBT4QqiWJI/6FpyHD6pdrerevBX/EAXA05ws27ffvorXcW6GWqjhDWGtKdnD
2nj5g3h9na5J/8zxSkdMxhDwxXI2/dfcfV0GnW0wa28xJ5o8jJPNTWoTm8gDcJb6
jkKtgOwwgzjJyPIBpuiQFydlGhjhOP7Qj2NXz5KF0QLA70G78O9SwfJoHQfT9i+v
Ntl0tQjlgfxjROCJls7cczDxzP1AqhpVQp8xceq4aENX5bMzrVq4YUfuyLkJwU7U
9GDaZszkPos+3VeeQQ6iMRS01vXgPGHjETAvXQyHV2mgpNjAVn7eDs39H+0oje2S
rUQqHqqehsNzA4Y8NXXxvDUD8f3lxWpBataasGEv+0paBzb3fspIkUw2ge5LwLTj
rOoflzIBEZS/TPfysZgBzAItlGbwPWBmQxOlNPVNG9CAHk2sads85MW+NeizaGSA
3bsZDKU/isI50NdQ6mAaCaYdESwcae0gj00NIrDnb+RkpWUFRXpiRwqaGkwujefA
9MztFnXwTZJ/d2w10u748QjnXL5pz1t/Knf/0omt0nRmsrM7NEWAalwekz0Avv2Z
3lPML1Q0EhTHku+E4njyBRViXUZygtKnLK3TOXQLR7NpEpMgXtbuAjt5DtZMVZ5K
FjCwgxmRvgJxRZ/pwS6f8xqCAdf4va53BGlGTR1Dsy8k5tKpqvV/4x2N0Xd86i2p
j9zd2ADPT75QOZuqYL09bbFkbBao5CHONgcjTcs3+Iz4shkJd2V6sJBF4hLfBqBu
yknwVgd/BhLIDPMtxxJgNRzKRmXzmNoMPWZWc3oBpEuRpw56YdZaznyHzc+LHnfh
hIBRJVkj4EjAT8uA+Ub5pRqIFmS12xhRXddyhMfErC9SE/bPHmuUAi87jmCEMg64
Gnh+n1NKZ66awvEWEM87iPJFbTcYy28xoCy1mGti/CdyKl14pNteSdDzRkJQr1lk
pTfPo0pwTlvQgMoFACBUmMXgfNKog/dZbjClJun1n2ubrm/i3dx5AeWPlT/yO28J
i5yoQWZpulbCpFqILzWZ7IHHh3CwTBeD1jqqprhIe+utuRHt7Yuh/gmvJ0rS5Lvi
hvl2gLem6h9ubHCY3vVreVU4HgDQUe1s0G/YjdeSDm+C8Yus2f8jCY1ISQZNYaci
VTnf1oZzsIikDG8StdGM+KKCqqbtyWO4A4YbyETrF1SdDTWI+eNoSAhi/Pa2O1j+
nFifiWCgOhdqs4jlxz/GBaDoTwpjbuVONXA9ynIXvKgpXIIvYsFPZ2NEp5aXgHtN
rNP3/D30bJdHdnm1SfNLOld79UtFWMJ3lI3ZliRzT+Mrz5rZoF2td8UXg9fDGMY5
xvxpajcTUPgbJOumeertaBFN7rNNG6A6sevfWMssDHPCTwofEsXimAJtEyFefXev
UPU4O8kyaBpwTB3yVDOCRZMYQjwE9WecjK2GwC8jDOPGzAJKq25rGEwDwRcysCny
rybzt2bu1x80eCJEN1/RLDpXXJVu1CzeeSO++Qnv3DA8uluHTsF5kqXYrPTkjYEQ
h6jDTl/gOnUKfVGUxvic73xMYZINQOkxW0yU3L+zbwtK0IpdwI/k4VynAhQc1qRE
tx0YqSU/51zZGn9JG/dfVTfHGaKzRq1o3o2iEmOv+VQJVQrvuY+kg7T6VZfSdJaX
Sjfih8znIuYU0itdskl49iHV/F2Rb9B4AkhaF0ZVZe6+laWcvfKuiqT76RpZWECA
DyweVf6NsSITy5n1Q8DJrZs3g/Mervf9hx/njhMX+/rm5YrzqCH0YP34RaSMn3dJ
EkgqsmDrRpyIcvLvBgkNsJfJN9sPEtSymUiUUihO/Mn5pQGA7+N/PAA6NF19mAUI
UXWHAkZYt73hptuqJBnjhHu5Sxy87TPbgcGbTq2Lvhk73GHzRb88RYdpLHIsZ9YJ
HA6/KK7VfhbTLgMDLAJPaW4bgcFp8TjTu4PIHcxVau8xpMe/zVj+pOUqU4SE0IEU
3bX/eptmHuxY5hP7r4yNMlOB2OKD1OqM7+oNUFT4GrjeBwHp1dNyUB/Qmi0NC+eV
fIixDpMTJPFLEQ9mVpf7pOg6Wx6mfJx7IOEP1QHhaARETyWvs2pZQ14wamwM/Pv9
/+reXHdv0rgEEB5GKl4WhsfD0BznjyVh5wmY43AiJ2Ns/kS7ywjWo1+p6EvP1YA6
39VVa1/o0BUcnX+5Tqk7FB4mnDzGFUK3rXta/X5JZMBOl/k9Cp4LLIu1iDprYK+z
DWMcoloI5+GhZhthg4cxuZb5MXI0BnQfjMMuXylFesemWat4ScVDeABlVFWSuMnG
XrXbDe+uFuHyFZh8yTPpORjj4I67ylcAJNErw5BTBZo85+FO+U0n5aMvqUtUZzIK
suk/Abu4LLMA4dNKz4mMa/yb4JUziJsNHmnasc1YhFbDxDVchRo0i3r6A7wwkbh/
dEp6E4r1olQrB8usCU0VC0XsDOTFOrvIe5GCS7d52WL/4o2TH+sPW1kH4KRbM6tB
lJ+MBLjgxyUnnOgtohlncaBesFozljFv8c+FaBTW4aRsFgYtkHQphAyVDB403Qsj
iwEb34UPmFP+JztIA6MIppIPIG4ZkNeUUqkE1jKjqq150zOyYnYS40l7J56hF16l
NCaFqWnTmoEzUpi9YtP8MsQAeExXEJELyMmqVc0WlhOoQwPfYLFwPnazk8QiHGOz
cFRNoVt+qFd4jr6xs4QMuSBrctW2hBE+1FbEsxFPeKxYCxgDBs69P6yKNYYkkVaR
/P62Uk2HomTr8Ejnm8gPhNZa5lSnZMOb4HJkt5Z1/wCo+WATdN8LsrhEsn4SKw9+
vprLEEoTeFQJONUGArMHCp9sk49MwbzkWLr9y1YeVL+bUXp4xKqC04w1z6nZVgSa
Ppmfms64WddfKgHxQnMUUbEwNVqPrYDLZtaEQN5m3ln/6vdBqh/PY0F4WpMzwPtJ
Rb1EEOBAymPvjj6Zlts8gg+viL1k3GG8P2MvWsjL2RHn88XnzA5JVDKpsmphkh3+
13io6T6eZL5Nwd+5C8nQjLc9BBAklm6Frp5+UB1d5Nc8l2u/otXmFN14UrwigbhN
O8+jm48sR/8nRl5QYASY+TKYpmULts60RptFLjkjpeiB5ubgiksuRyv4nTVzMTPr
8bdDCa6gP+Ums1dzVaR+NLYyEzK/EAvSAA8abGdVcAF1gZgHP7PRbvmYGsr90UBP
QYXpPYcXAWAhOqzzAoyJ+YQ2jcAA1IKfhFYXNvSd+QNrL0Yx6KbgQ4NxpNe6c7HT
eKKiUD0NV/uV0pY8UNjk+WJddtfoXbj0pZfyqxM+uFdeBhRHWH3KG3UJi1E7SZ4m
IZG6xjnUQz+1qQt82Oump66vfHeKM3LOPUx2B+vHuTfzMW7pTv1xWNqvMPc+sC/a
umQAeIaysOHYkQ0Q/GbBK41//t/1C2/3RHZiMMPmXZh9VPncrDNa1ZnDrxBFUbG5
O2dhmqMs43+Q0EFRwv2M4J3B1azSy0SN+TNfAdLoPwQuBcI6ngRFDbkfnXJcWMEi
uBtWJPlz11XilHrLnmZ5044sXGyXjko7xktDE+0SVahBlAT5mhxT5ML+ZqXukh1s
qdiFfMyz1lvao2g5Q5AZE2B2ZDR4qdMQ4dMXAjRkd7RqjOadtQfo0JcCIzwuPDIf
FL2eTomc+/L8ZKMNKTL9XMVL7R22zBr7Xv25KZ4ShH9ibMqfevyMCGCDRCALqebS
W2j4nnbM7gp1TFWo77ZUBwyqYBxwLiKGcQ6hKb3icYDBk9ItuuC6sFDEMcHx1p2s
EYyh8fcOHBCwoj3z6wkAmeCFL04b7PZAr17RZ6oTu+TVztcDFZeihR+yTi6mDiLl
y3V4Av436NwvB3FHU+gxuBqcLzR1w4RniL5atS1lWQo4NkYHxPgv17xd847N7dSg
lkkRl3KDBQvFjzQQRCS6YxphGFMKo6WGlASDTq2aUQ71CiSwdOa5GuYd1/uqXKny
AeZ7Jqa0rDmPl0VucY+eoTL35D/bY+ehzKWHU+nhkIWgv034/kvSrca4qkwOQBxI
5zcuMzM9oC/Y6BVFYeWKYvDSj49s5ZiqasgGkfsdlKEaUu8gJW1AMxMnjx8k2B4B
kRRj4K+QdBuVk7EkP7W+n7H6962A/VNZ8r+EJCxQdmkXrcz9LEZSAQBBNI8auGVg
N7Zk9YHG9Eq5Yzx+lAKdYyzDI7YOQiUAi2jMwnayr/5msECLO47wOYofAKF71EhS
iANgV1KCtQWK+RlHgAHq1P0vBGgPlI1/draRk0MSkPk7YVMZ9sKXUyoqGY+N5N6s
RiPPn2FBarsOmyLxHKeQDl8koWICDaHoGG5tXk41pscO5f6wUccfHb/QdeDZgqzU
ryLbJdk1xlzSLT/StOviZA3e5gZURV3Kc2OjRPVVDYFXXoOpnIVArPjGDF0miYrk
mknqg0ykmHmWcIoQ9pDGfxklMV7FJtjGuAt6xYwMw9HF63LpWOOLAdUQkq1yTKwP
AHTR9qLSN7hbb/lU4qFQn0McIZ8MUyFqYb32Ka6v2HbeQaB9EPe+5bKJmdgvA0VM
sHvBYH44B7SDvVtJpAvpwjOd+3xgf6xD23EcquuRZcUVPQBylXs6GfHvazYeoVFQ
F1kWDNf3prEgvA3Ahvp9jHjmG2vC81V8VZPF5ajVUipLh4tq6AFpD2qB2h1uJbB4
N9ljlUoqmVYK51WRlBQG0Nb1BtfkEyT2fRiI2rohUy6oax4r5a1S0CjnEog9ItJr
nxGaq/ZY1XQIa/9hU/mOfTJ1n+gCg041RQvjfkIzCCNbmKHIaE7jTjDaRqWevF9A
tMwzzOgAjtLGY33Yb3W2YxT3Bba7wOFEnZU9YzKOSeTvSGmvXlfbs9c+30RR2IOi
gRVV0Q/6dd7PoBXE92OQdSs5/pylE3d1ysEwtbrizpKiRGBkf2ymEYDBy9CDeAM1
3uOEFWBNsE1Um99iyx/DIDPZlmKBza+CiYGsFhTv2FHKkPckFQ4y2/ELZU/ei4k7
NnbK6dsrJmJUDDEMP6jbSVD8yeZBNjbDxXn0DafbFO86fJQQd4o1FY5sWVkBeoqa
Lyt+GK1N6wO98UZuVJvHbl08M9gxFIvQhOTHU8yu6/pkP4uNiV7qwIu3vp87bwEq
as5fAGtn1zC8Scgpwal3TV/nSwoAFueZeFBUYlMYnKbs1CnIyPSJIvllSAYUWuk2
LTew0fkf3bvnmNJh+gdqKCNXcU8vtd0XNq4rABDfvsHpi+suihzmJzX8XWeptDpt
8WgY5WeKap95G0aGZe3y2APut1LnQGRJeoz5RlINr8alIlf2f3AUguWb4zu19hwt
VtZLwzmhlNVTeF5RvbRpEgqB4OVY0lsO+QdcFz14fwhxtS+PyKF5ddnyoIauWg35
eu6r5S4uqf6PsZnjktbpEeMcSIfOVomOP5Nm8Tm7wAk0Kaupi3Q8V0qExOyJ5Hgd
XFw8GWfa4Ow84RtN/eykiyXrxLWSx8rEcKMWfNoW2dVR7BvH0kDNQ4Da17qygKDz
R+6wSKT+mbmo+9uxStxVoSlIEi1HHSwSUbtS0PKVTerDRboacNA+buOAOcik2aGO
2OI7heMkbb+h6d0kZlrTEx0OciUB9AU6FElsEAJ+DGzfjHLcoSCTe0suzcQJI/fe
doIlfDzyEszHCtEkzInx8EP6zFbsKIZ8X/C3Pq5g1rSWtvJeJXpLfJjRcplz4iG8
Ci8L5ypjFoSwWAA+cf/b1WBjx2qAPjsFZBWT05yl11hkFqCLPOEBqi9S7lt4dman
rExhpQzrIu+87onPPNzGUBoDkG4f/a9YUwVFagM5436dzEH+JIGYfxGNSl6FwXaI
JYIvH6NfzI/xAEDia5m/UxujM5Xhwg6wGEF7LbsJamYb5HSiQPv0LU/HnEw517CI
YDhKM4py3XWOqrBjZe35RTDxewYZ6vPW45Xcwo1HW3r+4cbYMRWfAkI3LFVk0o/W
A1ggFUDCHeB3nOrn7SXnh0wGrvSlg7Mpyvt+/5Rjv8Qge7cyt9DOG+wBhCQZ48WW
k/6EKMdWyZ4mvAbY/HCLbbQbm7Go03KDnzIu65XgDP+rddtiumtvQ7U3i5KKRgC4
ZQ+gPxXVSumuRcm9NzxMQEupiOdQ+2m/f+PHeXNq+fZKQQqVWu+PTboibpA9saO6
aZuSbM7wwkyanzV32YcPASAOb9VmE7O3BBaoatua+/s1hRP8gtFzSrXEef5Humv0
WcH9WpZ243gPgxkzg6qC8pp3WgAu/g6pjtrFc+S7OqzWTf2duX6qk5zV9pObr5wZ
ZBzQfzEfU/8nCXWtterXPMojJtJJ4g5XR86LXW1bOqe/NBTvhVqk56cLZdH7sMED
zoIYW8j1T+ocysCLAR8+aMByL9pfTZgz5BZpQ6uH8TNqHMBj6F58S3oN9ZKIAxHs
taQwdyiWJcR+162X0qs/lhCqsWnXlXIfxNLj24GFSAo5c5BAztmvEq0yjLve60Ye
cjRIeMOB/OQSA5+vnYxlIMAm4tXBPInEYCx3lnbEU1vC6B359nwAdm2Rs+Ii4exh
9aPMlQ7/HQjCEU4dlyVzzfdpRSO4LTXXB+gPmVijtHCV0ao0jSnSSoiL5uxAk46v
QM94HC5Ma0V7KdaU0Yo4nYLXJwspjzpqhtxbPiJxgI6tWD1fNVsRI2rvKx5epEdA
kF5x4RBTpu+0GLRI96A0QawGnlOtWfgNXEgol/KfbRTg4KV8Nbf9nt3AyR/rDFvw
1W3dhPXqAwqsFQi//oTDZcCtxud6viY9TuiDVsX5DDkXcwZ9eXzeFevOmZQDHRAz
/KPhm9o8Fp/AKL+LpKwKzGBlnE7SXrLpebv21NgzrBngsP4vimzOc/LFqzR0s2fh
Sn0jg+BZC6ts32th7t3Um4zYEWXDj/lfa6FLK3qJcb+1KpxsO/A/iiWWGJhDO5fH
KXtQVNiu3JoQC48u81SRhD5PPWbkFKKs02Ir3/c6UZD3bA4Qxx0hZsgcApgmoEyJ
7f/9GYoEBxgx59xzlw20tue4thglEQ7ewrRAd/btSNX7TbonsAx2e/uGFUi7pHoo
a7bHgLiKvWStvsZZTG8PhxnSkINs5zAzzGYIXtpm6/hOS3ZIOhJzz2M3aAdDqPSA
uNp06rkkbuLgvMqM68GxKQCTFtD/MNqBHmzhLotLjHpTUS+EBlshutICqc0Wwl2O
vlEqZdRoloMeFGm3lKLqDsC/elch0C+WzOoL9fFpezUTlqpKGwMFJ52MXoESDUvb
VUrCOqr6+eQtI1FOtuhpTYr9K1lZHMt2HSH6MrK5sq/QFy64+T2DihiGWjO3ZIUB
q+Jjsm9hfW1CjKAePQ2QcLqTb4L/1APkF+xlPoWQXqgIqXAGhW+apJX0OSMwL2jM
nJCSNU/R43o+tPPRMkzjbn3wZGmCrJ33VK1R08tpn49N+KwFbLng80uuEJZ/rzTR
WGAf3mxiksSK7bjxl6PUaYa9OXiRt+sUKAJkHpIokugLM8Lfq8erl9lNQuU0TS4U
Q0hIvD52KFSqg+kg/BikvWJQL3bCNuWsUsTm1ri0EZIJNlefpcUqX5J++7/IQ+7O
IG/VNv7R5TPsP9ykxy8VQTcVCA6P08aX2GgYaITCvtu4fzcycoUmMNrK0XmWvghR
ql/XWR7QO4WaU07TaDfioI9M2uaC4zfxZ1culM+/P3lWxZ+Cgwv4dQwwvzCB8qpa
o65j/NGUCrtCR1sK66/+qbwRhVfYBVBHmIum7jj2LwPm60sC2IReXErwKv2ru3rw
tmh5c5cCfb9I7ZNy7qFa5cJYxzXsKDeLtNSlpHX05G2WTxu6O3zqWngpNN1ATrE5
LT30nmvciAqFQ2CrTK7GTojHTPemxGNr/SPNfQ292HA/ZR3bygAmcaEbpNv9Y/lU
yJAnqRAS/cIEtMnWXiVz4zwawLwWeSoyd5VKYkRPIq4UjPnG/vQuGrzjxys3nRZ3
TQFqCqXDGnzlIGmEnASmWgPq1SI6dKystPynJPpNE+mRcudE5h7EpwKC7WPSJ7de
wzIulNj9xmwoEAhdG7C1qASWfS8175d6bxF0tdJpIppVtMyjaZ6PxQ6FPjQNTAwO
1Tkuhv/2o+R2cJgfe3EnJUTACbiCeby2LoZ748GQu2l8XPnMEhMXsALt1BhjHNTe
ydLkw5GhIW45Bp4+aA4EPAmcLru2dO9lDOEfLovv75H7D01NfwNEKW/rwU5Hq/tw
BFcFcJH5I12AFYhugIna2LSDZ0dnDySNUYHavjcla/ywnHXvkCmBJ8JwUCPFDTbs
BYGhmuYSIqjsKjxlJeG55CvIDcfnrczKIFf/zN+WZ67MWNsDBgxZ8c8G9xujm1fn
gzc441DkTGmsVNuCFy09fZaG53jGXt+mhWjtbUWByGX6hANkGfXonXEcCgX9Jcmm
hT+gZAS0mvRh2qbYGOBczMF0uXW8VerfO/b4Dsqnz72tPNalnpQeC9+noJVeuM3y
tF8AF/lc0AI61uqHoLQ2p1+zC6N6UUbG7x2xWpivtQlVB19FkkesO/+kTOxoKK2B
u4wrQbapoQOqjYZue0GAgRKwJeYzd3yGLihq/Xe6YeNRw7Luqvb9hA56FuCEMpq/
qfbAfZdjkxYC/In4gfkQwYMeF8UdWMCdp43csyDWllj0CI9MKedzTtR7k7rkRvVN
WHMqswjVqIWhy3YSPLTYwgQYoTCaf3KGcT1lePIFlpxPJztPMgPynx33Wvo9GN9K
omleDT33Y6hBHsY+qehe6D1Nezs5Aq1MHSDo3xYuokuBximttd9lrQl/OJua0O6F
aj3D0raR6bKr3TaEKZklGI1FJTAlIVeDRTAnGEqYSC+I6B+WmAIUdfDzTMFiVSE5
dvKbxgbLuQEuV0kEBseQ3P5Dw6IVKaZkG/0nK9LsaJ2Nf4vqQz7IhV6d5YdhWkdR
R5eMlhzYMtX6zmSmx0NGVzvw5scRPGV+EwU7+FOUI2VacB2BNdXJy8G79GZgWG5t
rB8KGIb/CYCERMZdpa1FZELDh+37w+tOhgWlcwzSE1HdVvfoL9/qhY5lM5PfTD3g
o5WtNd8bUJx2SJl9n/jOhbepKQB91BHHf33x3Tze8NggwQxqL7INBu6bxWDiRt1d
9ZKCYoJdCR+ZoXEI1BMEYbCfwD4FHSJsM8HHf/0EAjdop9CvO5NacpuaQdPfk011
jxpJf2Kds4UMktQ24Wom7bjfzNA3zT6Ck2McrfFaB40t89VPDHauJhpZBOUqYP6w
Gxm1H3SHMip25jylehWODQ8nNt/9w2ouW2kTN9JjmanbX4T6RTuyEwpBju9/lBPP
03gjVoTMeAFW/v48Koljc9lX0EkEAcKaSpvpORvZj/FFNwe9B/IoSLsILuh77naF
UdOggMFb22GTZMoFt84H7aEYcSOhdtG2CJEBbtp6XP1NYuXb0rNTi6oD0zjBC5DM
/BZsncw2h02v+4x3v/G+SweAy1H/UbLWwu7TtOrbsNfX+NMTx5/Tswnl/Yjq/ao5
M5UBR5idmjfsLVS8zx9eSoifJFx+nZ5USBKvQ5XOlF62029WHkM0jQIfuapnu1Pg
1jQlM/fwYwlNncU4Hotlz4GsX6SiqYjRtXOiKihsQaf5lyVujAKNjyMXaqfm2HSx
0/uUEM7gzv+7GIERvhzoGKjSj1bNF5v9HzvCTuXJwxcLo+phffGpR90sfhifW4OJ
P3nyjnnvHT+e5VoXDRvNqZ2ZWp8WcG0Vd6sR358GvJnjPMZVXalHYwTyJttuXjB4
eK2gNdxyjF2MkMvxWyAdugj69cKvZDn1SerBE9q+6S3bIBl/PY47ZR5OwXfXAWs+
AmI1hDI/3Lp0b2tpxhAi5LKCMuAT8eJX2pdCjYqiZfsp7ZuV0GBzYlQCxRnFaQb3
TMrflljTKoFsG3ajbDcJtdaVi2hVEOeNmaow4s/D7JvHSp8+ZZpuhB8uGPstxDas
xUViQc6hISY8+EjVAukVkqm6O68pNOc4xHiIthxx0GZFF7sudtdLoa6WJG57/lnG
OurAvvWK9CmeuAMF5+Dwixk2023lViL4R/yT7yVW6ysxxLRVHtQt6w1cXbAt3TuL
gB5zmxlQiEFe3Rj7JZJBh0NgyI4LMl1LESXoXRnlUc+ZuWDG+5tLa/uMobjHb5nx
HgNBkK4kxVAFXABjhLnr/itRurwnUve5lELbpGHGAZVTPk85haaqvetv1iWXHWRe
AQbbe13FpS4Co7eleHkbQ/MYmumivU6GrHbVLSDxvLeqGO4t/6uFBqDW1i6tMpOr
cHKily8qpcsAJ7rbSWS7LT1HQAhWL5lNtuCCGusGECN+plT3iDH3Plmznj6y6YAP
xEOUb9yIDZ33ZBo9PS1rSzlvTtvL1thSU6y+zHwwN5LsundRlwwrjArzb/1/nPY6
GnUOVBoTPUBzigYzbJ/1NS2KITiczDa6B+p59GdI09oYwsWXTSF6kJp2QQLil664
QyBrJgzWGWFOE6w6Fsam7ehbelEafhFgYeE3fvXF42tMm2Dnd8a7VEb4Qhs4raxS
zG3tIQgswLR4IewBoW+VCujqhAJDtbD/2sYjnHGoXBc0LRTLaWKMc6A77W7lXTFz
qSzRTG/W+0OzdMKz8kSuzo42tuHjS4PaWl2rB9kE+Wo+UMLT/cmjDjG7T42lH8R4
IBV0Xnly9qL06aEk60N7zDw+4pZ3ZGWvCP31sAi0nKIV5evdtqx0Rbx5PR1TUKQZ
72hFEmTqQorasxCMj9QJmXaZ6mobDNp9BBJ1LsK/SxnDqYu32JHUUk3aYsrfTgys
9vBqMTYheuXhefqfs/ShWCtji7+/dOPgp/8lLzIAlyzlGKz7FqewKmyXxuMcmQIN
KDtiYjghj/QVSDQEES8jHYrcYn7jFQNgETfebKcrvyvXhFVz+5AYDfVo/l7Mj+xq
2/tjxv38RFAbgioMcnb+rVnZC15Onzm2bx8Vv4HakTPRlmXp1DW9xTS44GzyPf7G
D60UcTXBO/TQRo+IHscEKRJC6iOERSi4FjFl4CDbc6IZkGgUbf3n/yFZhEUwnaqG
nknY21k4GktV9zg4aQlQY0Ht4g9tX971zaeIkvFcryVGisiqLSP1j9Ei5d+qcqcI
kHMF7/WSUCDL6m1ryGJAsUl47C2rFFCuhkhi/jq2vQVb4QmnAggoDsmv3culAlWj
qaCzPw4aoeHPLWIDselwVny/CLG4hTdLJLEGJBiXj8XcgOr/GmmVjiJ9KW2V40t8
P/ygnY7/jaJgKJss3aNEBtMXZ8eG9Of8BRGLackl2HTBXKAZi2VOSCrQGDFZFZ7C
PC6+iGPiK92ndh+U5WU2a+cvf+yRjCuEVWNUvAqaC1W7DmeoUo5XHcc4jJ6w0nKu
Ppg1i1+XG9jBWpbWu8mN3metKtjsAN9haCQ0QZTCZHHnO4jN4ig+wti6WUijNKiI
9UegWO0YdDbwFhK7SNIzroVTXdkU5v6lPS8/VojvjJBKGNgwBMfsaT0gztJxflnx
U0tzCP0Sn+hzKvTniROsn5Bn/t+ZFL4i1sQK5ucVVgYRec7KDcZ4qE1A4py9NRgM
Gq+/g1oVKpasRQWjfobA4+iswMYaDAwX+kP+lmTbRuXwAaEHjWZbq+6vg17SKmcp
5842s/eWhkGPdX5Ilur7UusbSkmNKjqSM4GUX/d/E3ncY/pigx8+gX5vZD1gECtE
w4OB6eHAalsZwrZx34pR2jjoyuTp9I0ZNrkXgrS6ecSO0rJV4wKPqwI0wWfLR6oP
zjEYjdI0ePfJlLrcsuw1XmEKNseA0hwEe7chHDtMdLaKNmcYkvqPS5F5DjB5PheQ
3rIzaIuqmpKFT/ALEKCL8gaRoHdTcb5JIGYWqkgDrNNP/TqAIDabo9CjJsiXG3Vh
maYKMTKHOy5Q4/6lHOHHCiC1oQv2xU5ir68cVbcDZq/XIEoZudjUw2rizBgUzmAt
fbGZMh6kWH+nk62e6enEq0R9C5yZllEtJkWUQqoqcQjfd4Zq0ZUQvpk/UY0peYQa
FKLv0/J0EJOW7HMU3XQ1Rdd6AiFEXgOahCwOOz5Rzc6lwNNjtDyzEXO6Zf4xjeLQ
ARg/vL+mP/ghFu/H0aS1fdk/OMb9QmduI+LYnqzv9/LCdWYImywvBsYsk9HxaVmS
BFDnt563M5UwxJUR+eEB2JBylCaMK8Xduvgh4wWMhWwRWYhhVLuCYBaDgd0AgPpd
dz3AZOi64glkm9FMdu7X3uOeCiSVSRQ0S6FK+1GLd5MT5WwD4Dqk0sQTOUbyzTrE
lJMBSSjjCkx7ZbkYLST4OVKf+x32PTIgNsL3mS9MRh6KV0qmDMeMNQysfyxmzuyK
I6mS5eiyAhLPcMkAXVTuvao9438hCauGMsYZHA6TrhcKaNa+LCussnHG4gUTF9C3
YfqpiaqDoTbA4exF08B4EjgSsC1XYqW4NhT9CJc97m+X+866rx2s0/AXtcbyFUpc
CBoSPX/ZD7Nw5KpXjVDOi1z+UBQ7/hdLWDphzQKZUK9BgdrqcxnrONTeDn7gr7cR
BETacaPjm6HtBXH/r9C5gDQM//m+QrO42NpuPZzZ+2aicVwkwqmbrLjeC2H6m+xp
IIK1/PZN6dspb6Ct4zkG5QW3feVjSy5nNHl+BZDvGNCwfWyxjylgiNHB3fnty1/e
XqvqmGnZdriShiqjCyqCc+/f++obgYVaMt6saJN9gnf/iYxjncnlVfJrgUFtSQZS
IHB6b8N/fUKex1zq6CfGaacG2UOsraEK1ZpJB2tGgxrLaNapeO9kCSISYJQnTUen
HaHnDijuXLQcKpI2J8HSMRNBPtWIP7nyTEqf75Lg3234xNQZBciL01ESCr1wLiR4
t/RakhsktKt28sPmz3VQKuvqj6QBswFEplIy/eePHgonRKHGdhMJG7OqxB2urJOh
U+5FfxI24QM1Dc+8Qlyh2Kd4a/JvDkoPJlNsuVE5c0Xjsj2S8TCQzWYTMITy8c5k
02eHu1hrl2QTbPL+ftoNvpjuX2r+rqNyQt5WnJdOqlCZzhHt7qlhWAFO89HRKXmM
BiZs3EyBdUSKE5bYa8nXLv5+BdltBzvtWqVqQm2eiYLByPWh6Wzy4TEYUYG9cFns
AzrVvrktaTz6REkHiBoKSOT3hbjomeoyN7XJ0jslEVOiLOpiqyhRrOypz03Bf0VH
IKsadstzCYUs7Fhv400SPt4gBe3+6Dk8b6TfjIPZmLyExbxXNpPY/juf64ESoew6
RKSZ1VZ1vdh/BcD340qvUcjqbAEB0unJbiP2J4oCRJl8GT5GONrirdHauwkMwzuv
ch7E/e15Sd0EGtM1/eFywGt7/QwDpCUZAc4zn6th32ypjD/qoxteKxfk0TRPjP8E
naS7A1+EfyDhF7tR9vVYmNSGrOhQGPqLsE2ZKlLRunUgDfZX6xuFumAE0+Zl+gEh
I1wQ892mbD2DFwxzI8yebJ602BxTMhBLNnnL99uO4EcXME+UJ50udB0fY3yPBfga
uKeXWfLtzfR58ZaWUw9czzICKbWJ310uIch/Rhayoh5TTp6WxcAynqel35O4a4xo
vsntiQUxGm27gL0GpaKzuJvwG+uGbjwGx1w2/ea1SGrPy0LYrRZ288Fcrwjwht7c
DDs8UyGwcHujbjXdUrGF9pqxnCGKUBBA+x3lya5WfxLIVlQ73LUAYG2it6jZAp4l
ie8WB0kAASHCfOXgAmMXucrrfMcmvLhYrT0wEuGjoSnRMzR3v0zzXr0NclCK0Dor
YNyDTLjBe2khTLIwxQZ/9b0Y6a9wvW8HS8fFvIOYIoP7pv77w/HLvj4sx9CsW1EV
R4gEgE7Uljh3N5Ckebv9xJQeMjLEOvvo1DHCLSv0dqaCLcfORhWyHkGDOIBnfPck
Ifo+l9p1d49XGJGPTMBv9NYncppF+W3W4jQ2kVPUTcZ7YMTmn8f5vX4kg4Xmob+Z
r4AEtFGteDLG+RqkKPQbFsxF95JOJLeuQl7NZT4Xouf9B2EM0yAeGG150urpBZC5
ldTbyqw7iP7DERMCf1jhO+KZfBZAHTXzNhoiXtSG6XSpGGunNKs3QV0gnQP16WuH
YVFEaDhz5sQ/DvUu7fdIHAdOgC3ph277XYWziyGddD947av/EjXcGURpEwlhWrcI
edeXVjGkR5pmwytXca721V3XM2FILrXaFidSf+fVslVGv2fpGzMYghkq7asxf9aA
Cv4F/GUdAH3uwCwvP7CFjdzX7F2OBbaSC+mCTSkUU2nNSSducny2NfXho8ENMx6v
wc+GVGeFWdsbz6WR0xfo7bfZDTWWKrWfFDXl8pYg+mklHm4ch33bEE2jfzlgMXWM
HcGeqqVenow0J7n6EbYvi4gakPDn/Qkdhk8OJYsjvzKoogr8NCl3ihkzllzFfGJs
H3OYeL6MOvGe8j96G9KigfT7WTDJo0KoDVsWbCPtHS7WiehJ80UaQ/3qdG2EqP3B
dv1yi7pC+J/LWX+KpCwvKFyaRG/5jOZjmupWjLHAQwB0MH4dMHUpexL08kzn2Shu
LvptF872/leRgEXoVeW040rls4EM8irgvp1ccjtLgKR8a3tkAUxhNv13m2RJN1iM
+JQXIUOcWIwibpQL3huszgJwx29oNR+jO/OYfV0DIBVJNztxLBmy7odYFEMyLsHG
5Ehee2LzGgD2eVxzdn3mWvJfso4P1IXKp2ejYYbdra2uItZiAGZVrDfpGY49hdoA
lt0Mu1AoAG4WcypXbVB6UlR5zAo0/CflGBGaaBuEBBtbjAdjPRhvvnhMVZGIKwmb
YgheX6+8v1hCJQrcLMgX6IITTv1U/xHcjJ6EHabqdbkjA61qgKaQbk6wAMjQwugq
lF+RRXAJyf8kTPEuDaj3N0ti6KULdv9Nx9XgbUzSTRJbFoYZ9Cgo/Iuk5Cs0d2HM
HuHCVmDSzLOJwT78LH5Oa+LHi7EvILJV/sg6mc7T0s4R4M8ah8b0alnDYajYr3Yp
BYZLe0xIzqTfWJXue88dDYqpyX1EZVNgkwyBhUXxIF9m2NCYAPFTfd4doeLO/Tfy
2Rhhn224Y0nwP7gmM17bWLtse/6bThCGwRuxjFDAARXl7sLvTICbj/2HTECgcUFJ
7Zfyt6npogoqt6jbuhJusO+qBTrSkqesrcsxdNjkJUStbolO96VRNBHGN85OJNlv
JM5LmHYtHsYmsZ5LiSWJOjUq6gWatIRsaMN+UEXOpwwsgwDjE4gO66zZF2hXCbrA
a0g+fiE+y8Nza6lm0C8jWgqaQsPzE2uQr+ANLyzgCOZGOHDwkxZwR4n2Fs4Wqa53
/sSHvGj0O8ebPLUxJaDiPKRFI52g1aXBdY2bn0/nboOru3sEzcUfEAXAwwptG7e0
VpCPMbQxY9iVZPf/rfsHsGVHBR423o2Ex4ISAKl4sZCskR/24z3b60ns2LRgptpC
FutAo7tDfIu656YeeR7XXDacuhyAlEl4PNpC0eHWcrUf002TMJ6DOql22f65YGl3
7GGq5yxTvJsQnZhbbtOo1UBWHGCtY8zsKKqebzQGybsLDXHonhFB66bI2w9xp96V
b37/kH5spWaCV3TEQl8FcIwjDx7aSJGGCgwEOymlAtVAcWb9emuKYgkEjd1hDOkH
sAWCHc0g4iEbCRxFKX1DgBWDMQ7D0NJ2O0P1gS8boh7s3OudgIkU97gkOBOqE4Nt
+N8LX6W8Nvksabu0EnEJGLKiR0snno7QdQkzaLpGg6/f9idsPvdVhLsGjX0F5aNC
Lr6j4Y72La/AV0e/dSvRRVlSOO7PoMBjuJuUgdb9On8HBrDSAA4qfFyeg9WFaVud
dHSJYnjio6iLmCs8fWp1rve47lomGHmaU4H0nVticCxAUbvpgv8mLQXohAZU1XUp
6NXjGnEcW6ecKXst55ymNxBWM3Q7KsrNl1gg3s7SDg/7epAgKD43X+ErQf40EuiV
q584RxI795l9LjCPR61ni/vf51eXTE4YyNp6nkvr+dbKCB8pGUiuhMcNy8B857Bh
m82Cdx9EASi+v4FM2vL9YVBV9vhtE9GzWh/Rnq8y0hClziP3DToz1po+BXAvleHs
OZdhI5largq7CxgGobd/uRj4Ym1yqd0gSdaOhXIAa14lg7P5UeTK3Xhse8wxX8M6
tHwDgOF+VKC4MDHHPTi8hGrmAKbzTV3T7V9pygyW6W6yrD3odbQHI4enY6kxdpNN
ecQuX9d3gIn1XrBh7xB9356nE37JigG7Z0zzHpUkZrosQZvvUpztAaq96mMYD3oL
qtPZRDEKvxMysBhNHmBWH+SwzfIHk2vCwqk6Csvepk3OztdtdHesFeZO5j89oNtJ
N6Qf9jETp5p4nfbdIeZqQOx9HS3VqoOZ3Q8NsyMTwoIR51P5BuJNNUE9Q39qxS4j
kzDyyLNi3j5U4xSWLfrCcF/5fLs5OJhdYcC5gOUQoOD/oBCXcfcAKLq/v+09PzsX
YY0qfEkAjQ7eR+cXNmUJyOOwX5oNlZeGPvyaf/zM89j/u/RA47DvWnS9zJ1Jgddi
NgYdofV/rMeJxpNkcJ/fRXv6ASJtXqTmv8wJKLhfgPVfLR9eH/P0or+/5H8xz+n4
cQyahWLnUG7ECubB2YVkai3hQbXFPzJHo/Ne2tlJSDpos1QGzVAUyprR68TgW4UJ
hAjag83+XiBtMY9NHz9Wl8FontiSIByscoWP6JWjbATuuW4ihg1xg2MHC1ao/vtu
8usbAdg6OCS4Y/oBdep4Q8vnoT9V761ZPYbSKYm6KSQva8vZMpWRj++yrTnQmwYt
faGyPnkeDbjmBzR7Hv1ULR4JfwdVfR2uEEuMXlBdViS4PQMLqZZEjQ06ttXoBHZp
Ap76kaztuVzpb2nbGno13baW0WdBg0o8TnLpxueIk31zEWnSll+mIptG4H2b4Tc3
wL1bkdfu4hH3BIGd7z/lN5htcTcWnx/dAOmL0fYuIh7lyRmGSLS0rec5itnFqiSW
ocVDVW7RVetmtllL3bOmEDSmkrX0LyNEaEF/nSw0qL9sZixyiSa4v+ujVsrb6Qfy
MK0PaDfxNvXKepUZ26pYtbWQMticMoWdnrJE/DfJOtwWW0mZc+2zFVe8eG+Hr9mT
Bwj5dFG5obs+dY3k+cflv8AhNHYNxRjz2zF9XCpof7ivQCDG37fgM0RLkCBe3Wr8
GEzNzI3NHIFS58TRQGbI8WG4w05MGs4j0YsU5PuiXJ2QnYUwTCn8NZjnvzJxlugN
Wv6WILltwk61UDiPK/0eTLvsAetSGf8nowZZGFmLuDiwjK131Roepz55WM5A8gSe
kX1C6X8xtpyHLlNgkRwRQeyGsC0n3M3CRcVRLcGMwjmtSo4VUhSJGvdDQTnX8b7j
GvPVoW5wG6lLYOhIDyvc6TYxEMFKQHN+ZgLPXM6RMXRJDEy3/07deqU5yUkAIXS3
NxhtQzQ4+5cTU2wyAnysIAAxSu/jngxvJaOi2ij+4Rxm8NebZkntBCmmNwwKQfz2
OSrqkqOBB6D5bLTBcB2jwEFTjhIVebH3pwL0XWl5bY6AYD7M+JY3IXv/CP4GU/lO
uuoBVPFAzPc0E2ZxDXmFdzc8mKd2lORnyCOJxg7nX76HVDNS0f23ULOtxnzSusqh
RscNsUG2wHzWgCIdKwN4Pxj+t5kt5FpHlbe1/HxzLbcMGH35vIziBPioG3jiRZbI
HeDdxiFBRBspVD0ptThxjB9CGZvyQ04tCM/IRL4D2oPhp9n2uXl1HEa+zhxIIkgI
+SzG1ErMAE6YNbMYzecy3I/6PDr3AIadlMiAiEcdLrpMlpKiuecQtRUwDQUUQRCV
zSt1pqksWKqXCTGnaJ5vt4B88t6iU3UouilhrqLhCuvExrrGZ64a4LW4rn13UWxl
t5oAAhd92UWF3k/a1XLKPH4uGpNobsKHw7SJNaGY0qLNfzh4NcDPqx8f4IaCZSof
ucjLO/2RCuWbSLEw+KVUhaWNzITLYr3Crn4lZfyyH9MnHm8T9D382h0gNBGeEOM4
WsA2qK2r8yNJEBtmm90YAQUfiKRXYiooH/RE+Kc9TxbyhG/xiVmSjBk5/Las06mp
fK8BNXM1ya8y1w6J7yDD4Q507FXxF1nNnBmY/5bSVBgbUdT+6c17kqe/zgL5krjH
ccHcTVu+0Uj8NYQHM0Vxgc6ZH+KMavBtAO/8vpidURC89crgEUk/DSUyU6A8huia
OyXkXwfdKc7RBCv6AdW38zgTW7prVP5kfaTxeLQQa97AwjQg8h50L2mxmukU25K/
X39WG2NNQP7/CpUdm6OSd0H4PXRr5bptjUamAWhWg526e78SUgKkTGo2puDm/5DR
REa1VodB3JcVFcdAbkSOWUZP0GYL5g348AfMrSp7/ij8wC+Phzf5Z1CAnNRKo831
BSCp7LpDDt1oViNGaY6pRSHxvr3k6whJhfgicIhVDNs/yBhWwG5ghZic+mIu39kh
xuJcXL20bcSLwlzR1BIj0TAlxX9BVytPymUfy2X9hf7pC7/PsFsMgfREBvVogeD5
9CW1K1jnP6wv46FYSrqIBesPSKNQJLZVJwcU26742GNu7x/9f01ajjmpr1dYcleh
MVLgsxYk4pjQL02IvEpBhWSQkkYK3qj7KwFg/kHlWkAfHmN7sL4EozI4XKM++BbY
HsMYTPeBPIoL8w1Tm2HElYSsGONgx5zjocquhT+DxpWmgkKTcLIMF3ax7wnsB2G3
jVKziZ/XBmvgMacOKE8jAEORTOD+hrhq9VLeaALFBc7TvaY4WQSS/0SgcwzIMI61
OzDguVff8BLIycTt7iLlorMzEv2oTfDAZO8SFRRM5h+YwUfHovXkQYD882EpojOp
dEMzkC0AkSCfq13NkaLmXWOBL4F0V7aOzarcFBnTr71drRb8AR5spQWCnMoPQ+SP
gc9/diaasOjfTr/5u/USEprtCKS5G+OpNMahOJE2wIUNTmggtxFWlkV9RVArp4ER
4JF38tvBv2oPjhboJKBav37XQEbuye3TMAt4JpQfiAJPToOmUYm637C6QbD7+C2R
PoyXf8bvLzL8GWfnPlv0XkEl5HAH+pe5NCip6rPb3fx2lkjJeCOSor6epUm3JQq8
YPjFyi3BRW1DcFGanIjw1rnUlE/xpuQjhHKADgJWusfCDHTYk5H8kfsSuMq47/jO
7L3PtGXR2StUd1flxH1XtMsRC2zxhasaLO7OyFec8dVeYp0nv97FmdC2ZKE04TH6
OWPJHRBRNUnUSq+u+Rg9x56PDknovLrA8TNs75rO43LYQ/31g/Kdot5KsmzSxJHR
O77fqvgX/7r1SwsS0ai86tvZiLdJMcn6NOgCvqQoimv2W2l/Dd1rwquZNpNT0Hi6
ud783aKuTcOzHGBoXmU0Xkpupf93X21s4+8Cmq96zldADptGUe2RV6l3cm4KN95e
WdGl57NuFS+71eTGOdhurOYJOe1UjF+FyzCV9VKb1V9akjUyWG/0waAeTJLozy6t
IYoNgwhVEf+N1zMlm3dcBZkSMH1LeGWcyJv8mOQ4eJ6bC2PE3XEPviSw6ubBf5Dv
LHJx3ltOaIfzpcjqt9r3AmaRYBfTbs/EZCozb+www1jFOiNTrqizC5iCLkOCGdvB
vLwn1oq+hHukvjfTs4oZ5HIM9Ygp5/7YIxHMV6xgu8AXCTrH1/qPa0qzK6nyR8ni
isxJy/LZYEMHBbta02sDH2+ZVYmFtEbPZugBmJSlGbVB4uHIfPXc2jz717NhFHwX
UZOdkpYcMXvI7g0ZuuCa9J6oYsqYFRVdEFPuNF/5HI/TjHwFmO6mh0PT9nPf7AcD
FS6INhuvm5JekYl1+1ObIe+8yneM8kW5uprKlS0QjPfV5UV0aIf+dvxpeqvOfOYA
1QZ4JXyNscNnJ0c9i7EOIqzMgAXZaEBGyrZzNjf2sABTw9r2MANZfJ80oeiFm1a/
ZdtHJg9Qux815Acwczn9XFy9VwldXRxG2/nJr86YHKhMNZVvuvsDdqAb0Rox6KNw
9BC7i/neNXGzk8F/xmc/iL1/w8De/PIfdhVfr7bNeKEbwcUJhl6TNlxeAcPBKydc
dHsg3nA2+rpRzpkcwBXRjKOb9Vv5BR7U0LNhTqZ7ruyq803y7PWKwTWnMLAgTbch
sjtKW/NiRNblRTk45mnC92uM7hhdIpmXOfCy0EH7Ey/XyMGSX33pXrdRCqP0yEUy
tVDl8oXJc3+feH43a9Ki7/tVftjgyVjTm8T8YKNinK4gXIytAEb0qHK+U35W3xZw
X1BD0Cc3Lp/ApwrLzgB5RstqayV1NIM14uB1zEKuiLJaNISuFXXBd1KKlIbU8DKA
mto6JE7FVzWclQHcQggpHpb8rmuZICNtRBVdlxn9/P0vG4UWATHTef9wUYhHBC72
iWcAUp+H1xpGtFf9JuIcFuBjoiG7a2m++QkFZbLsiDdAMxLzNAFbYk2DEga1hdr4
TbU4RmZrXhYogmHCSrSlFxINNqB4KP7IXsMOLHhQ/gXdOPTNKH2vGTw81SoY1ZcV
vSlNVZtcoX44AhzgrFBC7q/oF9agoWG9CGvn7+fCkocwctnkZi9cUHaBxoqwvyP7
phQbSLCXE2yz+eiZiIsZn3tciPCfW/rUVCvg+rnxmKTvfMcjimE7fk6Z2BFXWaBk
Nr0bPFngJOrDEzwg9ehI7wwE821V0k5fr0wB5iofNkKxCnJaVHp5XfPX4ZFdnlnB
dxqKeH5+Z6QblUZRJUp6aiBQmi30N8kzUZKV6lZem2vUsfVRZNR91o56qWARjUXn
QV/l2D+LJf2YzSdUPOrDk8nFaB+bulwGmtYU8SRIMU7WGeWbr5worv1tRDittqFb
9zrc7debmvzl7lavI3IDaoNUa1djdANYpT/JR8KCEp3UlrMf8MxQfCW+gclAwxTU
A0Im8Z8QccEbhLHlImlz4NlACjCY+LO2h+v25fNikWPxO/ejHeqqbR3VF9T9EARO
3a7x+x2TFJZXd8ncYPbnn4yoV5JCBK2pB7CzYBfEw8/oWH7uhC0VwSoYCK2CaUf0
stStPEffyj/zqq2MortL3/luf6QGYfgvy5QeHPmSxnrWADcuEGb02so+WX+WI1sM
b3FG+h7IyuUASal3qlA3Nbh6MPeSYKPL9fz7BrvzvciTRnjbTnnWdzAJtkFuH3kx
gTgIi1hH8VqzK+sDJSS6ioQTZjycQofcx0/qHjQKpjF/esIt3aZIaLy59QpoiTti
9gDQ0sY4pRKhFpc4r9/A5qEp+KUypuPDNYk+B+sQwCvZvQOEmvIyjIn5q0+hKugh
HleEUC91q+ecQctdoDav3ax/A4u95qoecxW9X9J1QJeZZa9V6qE5Hy5a90Ov4q5p
c3efWD3CWnOt7Lwle6xRVJ7XfZA1sJPZkjgwp61VUIE3WcbtdtCI4V1fTDBkuXAm
JeKvGNP170diYNEIR7YCXd+ZFfa8GV0V28deGocAGrmPsOiCPsMnKKjgO4m+g8Or
Yyv8sWodyF5bGwvn2iSQNdC7GQ31tMrGh76Pzd0CTtEyTR5ELRPZBrxwmudh7CCC
wvjkC2B5Dsl5HLm2KHoSoj+3rzw3dg1Q6jLkFeCQv04iVSFEnceSJG0Pee1in3GO
rEpfhP5qf+MW3IpfZAOuIGwyCVM6W55OIOpKpl0D6d7rtverR1S9hQJjlGbDBJA5
7xmM3O77L12zFG+T6FbemDp40Vl0YiTZe4Ta7/Z1z7j4jFXerLYwYinTh1PWM/vH
0QA7O9evgArqisXqGCFawttP3LReKOh+o/rBgIVszl13iOmLFAY9q+FOVxmsFPNP
3Qxjt6S85+nI6BgHSY2QEMdXSf0x9kyrYVUNdue2dIR3HFeNKmZObx/OjIQREpKF
e6c9Yl4OVIim2nGtftqVyHvg7aSeWijFaDV2dLisDEYYZ9z3SMsTh05BGj3aYjOd
hQD3szOUs/BwgmKLJ5zUCX8Z3vUx0cJ4hRC6z8Kizq4MMCHVxM7y5nawgvpLirNd
1Hgxi+U55tVFNrmACTfnOcrcpFgRaWgC7B2TEuZMDTVNXECKzMVjrtVSCX8A9hWz
xPWHj2IYVRTBbdJoaOq0pPDSRFDn/lYzejjl4d8xIeWBXq9haHvbZmdP/fuV7etJ
LBA+Os/wyqmUqdZ3uQLzLbC4TSd0il5SyWxAtf+R3rlRH9b85XvBHkmgUyOk+iWb
ptCkmoSJ5ENrNA1rUt/ueH0hZweGzW5aMtkSaoHjCTmh/ZE2l2pDMi2RHFo+ZRCV
3gVeQha8BNUVvbx1BWXW5KiSfUDg9MkoKWY/VaeGcClUHd+8bVLjUtp8CZRRyD08
/jPSLmVsauEh+kOtAXAJ0N6m0jZ/NG/YKw+7Fzyl905AjkzFD/WdkCsiW2QNfaIR
0LIcoMgyG56sdRupCuWnRBHT3/SyOftn0V3vD6NGQbg+Ur7xLSYdaFYLDhi3VLjj
ZnraCRBL//Y7NlXLrRfkMedFc3f8+s17iO79Cki+fyYfU5f0KB28lR/kOtEGdRgF
AAJllhB9mcveCFg9Q8JCy2UTuaETWXFwufwR55r7KDXO5n1hgIlLcdUTQ02u+i6a
aykZFurGty4oLkFBXavbO5HAdsRdSx4wPGEg//aTK3++UYrhrAh9L04ryzfZ8Vgf
dxWkHE7SAPtv8N7IF/GSk6IlCznaEongnkzgawgan4yfcsTJinvWXijAIbTdAmkF
1bl+CAdKogTsic1br7PI9JUCT98IVWoerLLb6REzgd3wcC/iZKYpBGqbXyJ9aUib
TSTDObyq3Ja8S/wkYF5WHUCg3ZxJchnUe2W3N5XkVsRjVdd0oKf1CCIfMqJvp+Ft
Lf8Mz6nA6o0bx/7E3KoiPmrp7HwxHUqzdbJd3vHmXkOFrHxIyKohi0iejwOEKdRb
+Rr/l+H3tMSvQk+FX/VBjjFRj9JALkbRmlg8GAZDTXh8MNnVyRANKr1WzCT3Ppk4
ckICAuJ+w5MowvhtTlk8ugx8mNuYxY52MlpYswti0oTYEIWp4zDBETbUxLuejATy
JqQiu6Kqh350DeDOMRJIPEbjYU3Y0RF512o0HJ4Kcrj9TRIs9p/J1GNCiidOjLZ3
4KsMluAyl19DzKTtSl7srdOS1/OO87cG5xYPXk3TPxkJWpv6CrHQAlCXFdyUwi6Z
8yYZ6/PKXlODxP857XleK52D//mh6nvFRR6ui0DIi/Scv/De9EZObSNitcU8las5
EwrSOCI/KvKSFme7TGGsy5bZ1tK7JC2+ltHlFeYSYa+fxGrTP/r7/DhzzA+B0ZdK
xsmfjpsnXJZ1NKnsycBcbpP3wsWaWBV+TipRnRgfAptsZWFtgYONGpouMGSjveCp
Z6Ra5F4Jl49N5nT54Emr5l0VpG9oZ+1oq7XdwjqnTvemwIgX4gBiBqLP7/PtBZfk
cVgoZsRZQP62FW1mjoh2nZ9TCK4JlOkmnluCbiLSJOgiLwNl+/x0lmlT8daocIJM
oel77ZTwuJaDDI5MG3jRRPMMjl92qZ3JprGWJGWEd3iogUo2v3XvHS4VVJV1baYk
ljkACTcajOQ8L5JbRWR+JNCnFalJzMXmsamN1hgly47VKK870tuRpYCAsaGE+OHx
Fe1Prlf6xqTzU6+Hpv3bzSa2z4ODNYHUhZL8HEc982L1l7av7loY9AblgyE8YHGY
00GkJAf/cnvNxVFVfJr48HqW8caOQPVAxh+if+7SpegrpO7CqyKO9wQCwgo9fMNO
eTiKV862PKTNP7tYXLvzfPuxk+Y2xdAN3xg5pg6IyW4y1+5HFwa2pGljzNI1DMza
d9qnLAfEJF4AtVk3b48EPHRRAv+WGUnVcafJBZUR9AeBsI5Z+OioBroVxtzhhrLx
6ujooqvQpnYuVNV92AbCD6+YmTkHAjyKgjdkvTetYePo3cM7MvqDmAY4C3ENpaJZ
UBaLJ0ULOkh43esxE2XhLRys/mRYwjA1l0g6d6X+ml3YncMHTa+Te97PrGTeKkFr
SYfbkXKdk2beA1u/36UGpRZS4jKD9kDpsDvXzabnptGFOwhRdVQjBdbo9vziQCCc
re9ovdP9xMCfCi+deGt930tR71OWmzhZgwhQ7ObeiGVKt3ftglx6VJxsNwieBdpJ
oAVo3dxjVOH+8xvW7ZVcFn3RrRIP1bIPjVEUKxT7A4XYLokP4JdHcQFpgbcK4Vo2
EuNJwxy9IvqT2CImG6AUdpG/tHcJl/oZfZp5UjrR9fW5NP+uDyvo/C6hFF/AF9d/
mEmAgNQQ/Re1qxlUFOM4ZoySs8AmBtzDuTWFuJMODIFJez5nvTK40xTaXh0Dene4
pSY9yvSICdg3IIYKFGeyt7rQMgIaS+hb3K8pwLNJi5jGdeZDlo5s32H1NBxGxN+0
IHvH74qd4OhyIWKwhcUtD8a4U4L4ZmyUEDvppPau9qVozjzzibO+ReqPor1fFo2b
asbJMiuPy3YqCqGJbzmJCuzuasGl7l0plS8DnW60htk+vw0yt9IUhjOi8ZRpfuY0
dxu1B0WnjjPa9b5VcaKL6hbEfnu92CgyFBPoRGnOmzrI4GuXQYTJTvEpFUD20ZPX
yrkH/4YtUYngSrdMz+OgBdOsblP6t7EE4y/QFpTnrZy0ui/2kmjWqcFfW6jfp15e
5P25QS3CpJ4/TIUuI6hTgxsdAB3bMUVLdELNXWgQ/1HxXfO0qkRjsSY3LNoULwvt
NTnLWr2ViVY+4gphFhJbuZ5FYNs/kwlCIt1LDT6I78zNbMDKeY+akUri4sBjVmFF
eD7uHocBfLUvrUi+dNlZAmynCxHzUX6LvEi1AAW/Qew91rtd/O0kexSLWS87B6QR
V/Qqhm4YMD6IlGgVtF/rxBM/w2LGH3J2xP5px8pwpO+jkVtuSyaQrShiW7lEk4ie
JHh3RGLrri0wS/q/26ikYu8R/ssiL6BiE1m+t81wS1SlybEeimA/efrsKzVolls2
dkg7EmitnF7M9hq7dzbfN7DDFsU07o79AYc/1YHB76z9Ri1zADchc1UDfeRNh0DY
ytV6DDpDO+hm2q4iJ80K4iMc0dmEp6j1R5CiBhoaZFgdnxEEq0AGPQfJMMWbf3r3
nF/wm3swNQRIWoIXrcm5YT2qC7KhVint5mSJWoD0dCvtv7fPtMbf8s1Ta0oitoBt
7n+ihHWlhVNuyZYegsg6/QJcVpb+/qvpkU/EFmuz18ePKDPwmhiwhCz5TveQ3xuN
lTe5cx1c5A+FC+rzgYohfZQpM+UqB3G1yTHKjhZKFBSIw+jBV3jI6FL9y8nYqtxU
0l8pixVWJuSaiI6wD2F2FLg6XiP7t5akF9LwjyXrM+WaCpr7w8T+E13XrGqR1Pb+
JEOT+aG0mFc8z2AM6Gimmm62ErtbKukp+9+ZvSiTVSCmTBJ/lWNd1MQTpTBywAU1
LoHRS0sR/nTAddy5fim4ReUV6+LJiQ2380ovIr23qIQyJrObix9May1kjB2ccnLX
WjNp4NenIhVKwd7Q1DiFSsMQJEXaZm7nZbmZc1Szd/iV2FsWIbD7uRK4ZuQIkU+m
RJfaU2rIOYccXxbuPGE/vFeVqiU5urcfyf1l25h7CDmPnSahlttwL9l6GeMNghZr
BLoqkNkutd8YLzannxOs/jQ7wRTJCh5rXruyrmGJcoGgFtuq7a9LFLxK8jfjv/eh
hPqd+iz7qJI0QKkQ4wXGkRrZmL4Wk4lY+aECxhcNnIPRThdeC63oDLcHIrJhrWg1
PVPIX9iiMNDAvqbY8gM2H7ElfpcigBRBWKsGGOrfDAgJEGDV9xJA/9Fn5h7tln51
CIo68av9sfGZljzWGGuJF/wzxfZYHig0VYvbT/e96QrJWAmgKmFf0YMx5aEFtsPt
C+KsDvCJFWtHA11XTWAzmcd0xyq/YrGkzni5iu+Tixh4HOz30mmVSPO8nTpCEbyu
0iYNPHbPC6Zyatx0ZSO622AR1gGMagVMP1QfadOAsfxipLHjnC449dczzbFavHl5
oDWAYVn3kmjnbo/AXKv/bPKTB3VPmuNb4DEWBX64RLP0A07kR7doBU57XZav3d7F
+QGa54xEnk3YrL7Jc7UfaAjMZi/UURNi1zk6yTzWq0UUREaNBMmWAa1vz2fhHWTX
IyI0nl/03CSV7VoqhngnJ79ZXJcS7wdNuT6D6wjglDWxFAKwCFLZ65mrY2c6/Sh0
YgasQS/KzhVJBSkGljYrcXbq9FXGbc9DZlZZhFb/41Gh7EL2fKr1Bq4dUg2T3pSB
7s5c6Gq5ucbm1hoWE7Ha3/sM0QgUJhHF+cs+bB9WTgUEadz7gJPOAJG5aU0mq2/k
aJ0Wgo9BJYrGsbAjTYfhqnfkeLNR4R1aBeZh6p4/WKKTYbDCBp2xzpoqC8q03KVc
RY8AWECNiihcIs6htNFam37OB3QkZrGyMIIEzsIFMp0CvAbQIevaYQhk+f4LTnyi
2fOjW4YnDuxfrgbOKi9KPi81IqEAmqhw3hjQ+G1T8O+kPrOQ+90Bu3/4zp+0+Hq/
bwgKV9z/KqSwW2yQ4etJq2cmjsgNSnxDPe3zgtPLe4duXbN9ikFancDjP+OSE4wU
aTzd1o7LkEffqeAZdrGADBLbKa/BIJMsuai0qhmVkv8+CuB5qyapoHN8xTrqRSpx
hosjl8zrFtv/0kCTUTLEFc6ioXGl23/ntFtjuOycTl9HcQADoJwrEeOnPbjuOrvR
K/P6OMC7R6sqsc0bw21jBZadCm8ge1y7L2MCt62+QixsxtbAB3PvQOYyr/Nm0w81
Sz0CGRl127opULVuqf6CtcnxXFd6VtFoJz4cSyIQwSKS4RKPN+ELUqljW0jSlycp
LcV5sP4mNZQ3MaEOrzM/WzDrqv6lkv5WksR1vhGjsDnbGBGu6iab8xJovu5MijSy
a885KpeOc6N5MO4PQkVqA89DAzM1fgx1IMVi+NOSfIk2+BDHccSAwLUVJD4KVu7a
2RrUr5z2MipKBy5s7lBq3d+GEOn70hNFCuNA1sfMClGGI+GmPjWPeE7O04GMLte0
bJo7+qiWtpcbulj182o6pccWrErytuQcm8COhXCdgyZfHARKcily6YTS2/8r6gXr
BA/8RWravDofPmmtBC7KxD0Vm5uvpzcMmq/iMOS2GrtNJzrNA12qKVWQbhptnNMX
QTlOL2mx4oSjkXr1MZcpM+va9m7ekNglIAudmyvfKrVh4rSa3ndnxvx6195ew2OI
6A07/P1Jw8J64rD2G1nWXEDwZH6FwwyyIk8ZanFzVLYziSOFmiEst9Z8E4FYQNMx
afdhL+R4PGbc5ytW2jEZfyQDDEuIbY1gPa5+r+wjCZO3jjmSsj6tk24oy3DJY7TU
gAAxc9fMBJnUvvnIjgjwMMjnBxuuHZpAS+lWGoP6Bt2ez3GIC9vykpNCY977UnEn
5x5D5x1hGz7kTMWVQTTUziVJdb0v9ayKG9iZNYY4MpLY4q2mVsmGuEJxxByLTbAs
x6ab4RdlFmMnKxeMkTf4bc94pruvznb/9JBz/hVWVIWuRkmmVMhdwF4RV9mbyFar
8j3m+/eRiM71pkDL9Lue95WnBqFTjG2OfU0jm5+bun1U+Q3KE/vp0D1F/uq4YOt1
gU4biqHh5busjVUBoyNaWtCb9tK1UVa2EFePdioNg6JP91AHTdnLTEU8Usss10Cj
4mTcc1rorHQOi+VzsW+Gxsbw1e3UDz0zYdbaJ/Ds36+OokqhLs8kxef8/RDiy/kZ
QFueKzgW7YOIA7+mI71diq9gQETlg0Y5Sr1OzjoPFx4vrvT6El909ZnaXRNuD6NT
a3asev33jt5X9WyrkZpt07paIBTngIDtqwEgiMuXOXm1UNMPylPrY73TfhpOqCbL
fmNeeCKnD62qYYrrZ45RLImLDtHiJTmP4MShX3g/DHPq6OK1UjS9sm/4KYhvoOrJ
tvKljDXUfGXD8JyjkaJRn0KPON/rpNRzpEECWYAsGEONnrf0XjXz9RyOPvSrISpW
cC2aEZsVcFpG+5U8o01kzCEoTUPBiN5/LPITi1oPQg0qAdqbn/FaUBD/h/+2WBBo
R+l+iQGWcFrKAZVFiPSF3bT1zosM3PKDWKdqX1SlCcAHMvwKKHdoX7t3QXU3K4vQ
oG8llsFl320BQJL7LpoaMuyp3rUyN4P98Bq8UFPhqRYRTnA3hXsBMpzoN1RxYeAc
RAW92PHbPH4TVitlGu9cxWlVsH4D1eoCcGOsYdPcBHY4zsq6PqjjMBqOrQoyW89a
tQsEfti6WMiJRBrZAtlYiEiiX4GjHKJEHxL/Gu/ezt+QVZCOkS/E+a1pNcMhUV6/
uw9j5eWhZL7l6DHT8trwefhw8MgNVub/qqp5YAGl+SmXSgBTMLe6t0Bz/dQjRKvX
28G/w7P6GVKmgOWCNRV6Mz4XZQZbcHXJobjJ9wd4Q8rvzu2R3u+Re9w/a6SC2PaA
kL05CHOrYMyX4VKjYlX681suXEPxt7RovPNhiBsv0846Cg9V6BmrkMLLiAOcioWI
vC0GoCgegNHQy1O71L5xbih3BwpYliccjQCKLnna0XwBEb0Khad8EtI18/g/4okB
e64PAKzcqxTFKZPsVBeyDqzO1it1Hp7sTaokTsUN4az8HiqmLiVXTg9zHX4kFb3/
Z3/n27BU7QTX96suVzkUDh1oCZjDHY628MqfEN2hdWFtehhBJx3qeSVdL/4DBfzk
K/DQMiyQyaRtfzTgJxzafQjyLaYtaJeDH1XJjCO8+lFiqQDRTLfb4OSvmpgugyJo
bzmsng4acwCD+TLvJmy/mEYlp6+iZpvX9GSlQxNbXs5zGfgCwf8/kvM1QKfYHYWF
sX1fuaeYCJr4hxI2if17qTOOZxy5hhrbjznQTuBm7v8y1xRC7ki+IaGAtgV9haln
+DOx4sIO3BOp2WclszSDJGJGxSMiXVLfwjJHHCPgKZRT3/FepeZCjqcGzAuN5DVA
HvS6z3WtlpMECF6YNPZyCje61SbH5ITdKsKBGNCNlStBUsM3Igj1CypxA3ocrntB
UthsV9MYk5H4bbdtmy7tB6PS43NkYeBX5pF+mf9hJsa93xuN4xw0abNNjG9eRwEu
r7bECcS6YlHVCUf22EsK5OZDcBs4SZq7uyn3CjbHu9JjVWzRbto8diEmRrHId5zg
JPMLtKxEONM7qD1hNfQNC9aHkK5VtUKUV6idUSE3rJDCp3TiIQWjCWQONzz4pNjA
DEbVDAlgaShnxAkNkGeQ1B1yVCEoK9CDijDTDQSwrZ3GUayKHZS6uUh4bex1gbtq
1UGMcZjdB2BcP2FU7LU7rb+S2LNcQOyEjAI29h0/ATEoEizjsWG4P2mY6bKZBvY7
8dwg7w+CWy8B8wFwm6zJXMLqLADyDYFqL4f/jxXhj/2U4wbGXkVFm+Jrj4kfEnH/
9gZhwRbTgvQXK3GIOqaYrraoDNEqu5FYB2yWi55PsBPTa2FPXGCkXjIHWMQtrp2G
yd1yjDVyODNCHI+30+5qOSLZIEo0XtumckAQ47TPg59zqVpjHkmbH/5NE5qcWJRR
2ih2DqgLXRrc2s2XTgeuZEATuW2jJ1XnTE3S6HmOweQgH9pSTN7ZLqCKVKMUF0b2
jWl9xr5KQp7eqrw1cfflJW44o1cAheC/n2CRCHgq9/bGrIuVPaP/MHyES1Vtq69W
wxPfn3xMBx2X0+FrNa1hvz2eyiE+fbFRRb0six/VrsDNFuwGNzM2LtLw7nQOhBWw
/7a7hANEW0f+V5inICMYXA3teyQEPKp2T3FWiTMhM68evYjcIFkfK4wq7eaVv3ra
3x2UsdzvmYRm9TyRaDo9jzvfHSI/KLHjJbfXB42vRZuXYchB2utOUNwpSpyZ4xfO
5Z4Qr0xNs0YeJCwSi9SzUKZEXCUR7AVWnUoey+GfYp8J3Bp5yzWbU2gRb1Ouu6Bh
yX5yp4VJekTScOZLiMDTCIGYGsc9gkEfl4uSNu+zszaxGxRa5zjVBYBOvOv57lwQ
q0AQK9UvPCNQJ3XoTQd8KMBkufa032bYUd5yNIkUJjPSJUM93Teed97QpW+OXwca
LlipvoPrTsbT7y1cnWulOF/KBHA5QfZr97VUrAlmVq1g6jHVRHZDbSLTmt0ofxaZ
KADWOsD9llRsdhzHShIvBspzmCHshxOBE5gGT81buEfApaT63X0l/wnhWm4Ymcg6
QX47BUwx43+Ss+on+PVhTe8A48p8WdJLCG4lVPBHSaNF0WF5BMl20eVlIGjmrg2N
y3bqmS3kdHjQsL0uxtD4Ip4H/TPX4jWVJ5RS3si3BAKNj2k7fjXqLhvZBesi50eC
LOw/bd+MZeLlV2gl7avwpTj4HZDh2IPj6JoLrhR1jRqK1Ib90fsTrTmchV9n5OPz
4gNVl0D1ETCD/QIrRmTwf3eiQmD2H8Qs/84hJYCbO0hm8N10EpnwTNGBBQKYWd7/
03xjMakZxjqy+M1yDpStpyz+QnHwdJ4hQj68k+8/ZYRJusDAHzEj1JMrC7808S6S
j+oJVpkaQnoKyRqWdm3jAgT0HkNV9VQTGmHTp9meZZGOmcyc42ZR4vkbrPoL6bKG
77ZfWNDb8SeGcqpj3tP5aZ+Wnk/Ule+5e1v0qbfv+kfrCBmhImgJZquvjdycCc3q
QuA25tiOxy0OoQbihMvwqRKy+18wb7th2wiXQKllgL66uQ1dIyKzdi3r7lkXQ0sI
B4eA4ODDpU8JlX62hcvwWX0Mnd8Vi4bXxf9qLXuqHRwckACzxvB6BC0elolhqTaR
yac1LAiggkCILYf1zmGeEd1fNX1ydTbD+fz9onYHnqlKNUnUel2n4TweCOb3pgQQ
6/C3H5uk8u+0f16ufJn04jKN7dPXny6sDKw3IYTHMixVCWdbv1JJQ/SSXyIIypQR
4El/KEKuFRwZ/XpfXW2UGUURwt+EFFuziOuiPFZ6aOqS5Ic8ix+eJ+KpdYBPeNIf
xtn+JojOpGl0d4Dd/d5y4uuCVKOYY5Da1Z+h4Nta1TdyvdQsz2+IeLINPfpFkGPh
Oy01tt73fqA/cawP9C+e8Of1PtGn4aAysz4QChaZp6vkKTz57FnDHgge8mfI6wbc
uHA/EGkRNtf9Era79Dl7rPmh5rjV1uF8gBsZ61n0YVqUXL/9c+6nQru7rDqDSjOR
otdFgIme1xDYd8eVHyU60i/xRrcgGMhYgQsy0L9uTHPDg6IulW86BPVZ8X7pZKAI
QGxR5IPmbXo8s2KysbslC44he+4UrYaN0R2oXzPOKpttpi4e3M8Hkj+Ka7kBCjlO
WQ8pHJsEZrJP9f1329jV32dpIFEfkkmEklHa16wjYuZ7UDVSe0p8/01B/1gLAmSp
MsqT75HmyyCTFiAkQ/uT9Ks7aMoSCWZasIKNeF96+OPGvifi41pLjHVIJXxo9HRk
UJSm2thbMsPuNPlVFM3OG+a0bv4q2ONtMfA2xhN8CG0krG9mR9E/J1tq5G5CKcyo
5/EC8AVzOc4CqruchySoHQe+NWBVkmYCXO5qMrVKlN8VU6eZAdZMDdN4ZxNEvWBQ
stM3v0Hx0nOfXHnx/mYeplBGDP5ipmQM0aPu3ti2kLCLnfQeABJI0Gh8AFM58CmA
cSq9GpRoeOjbhWr77XmTOQwuIf3yXv/C4x9WoTG0x+pMAlncBOodikamdySLnR7a
gytkL9Q5iiDcUjRm+C6gka9sjAp68J4GM1suWqqhDhF0Z5txabP2KjYbkqzBXwvC
bAfOAGRV0zwBk6vvc6yKjz3/j0AVBTVJjsTzfuz4nEjs7RF9CTO+53emdu5pZVO9
KO+N4TeW3KAPqjnQDttq8wou62ELqCLtdiXFoejve+nkOfJXmnV0wH2e908+7OIV
zzl+qV5C7pOtJROuGljKHfZ23SgtOxM/XHvTbHeUpkceBmuEx3KDPhls5QK9O9zv
fGqAiyVSI7uBDYZmuZ18lgNk1sGHEq9yFsyVG8thYZ6bt0sYD2gYFHzddhyMTZNM
Cns15ztfmYTRL2eyD0xVb5KRWWsbwFYrRuSxP0GZvxSu6CVmWrOrpbj+ZibodpLD
TeB+1efAbsCOutz6CwRDfoJF2pzHBmY2MOaRYYOCSaTZjfRSXWC1HfsRhwsQH86+
QdSyrpSJrKMDxTPX1aquITYXPCS7Yaini3UDqDPWSSQ+HwNG3FZGM0gQj26jm1bl
QBajL/mk9RJ9M2sKDSUhCCqaQZQV71h53T8HqvrXcc9RAf60LC9w6qpU2wc6DzPd
lLGhx0XRagWWAIHdIC8Oikar86K6vDUOh7MU9pth3McbhgUDq1b+qF6mjleHmg1t
9/vIQ7XkB/Z+aOoUFMrtqRTc44RfGKx7XKlEhOeR+URu7K0piV0csjAMsJF7nvnu
TOYKNGovAHYGn8GQc76akyFKHrmTfKZ+ILwEpKSzYUgnsr5WGfrj6eHEPeAhp9G6
qr3ndL9mI6ledLZEdzuiPN0VkcyhAiMBRjkY6mpcEN1i2xrNiLTVkgYzrzs5J81t
LGp4bAffSfVMHhEHFqwsRzqDkHC4+AcsTpFSziOQ6DenrRF9hdvEiq0V8SfHbeaD
qYD441MzyyUD1wk1kmtM0Z5N7mFir3jWERF2K7Z62B3JnI8lDnI5lUzdDD6jNxXQ
l7YmKoz4heKTHmNpzjln06sIfxz14O95WiiV4jFEklWTlWzKjlWka6s0Ag3B9iZz
wcxUx1SwSoAv0Ox7EhxCvqyKJyzQBTD7T/ReMhNZ+qmdJObm53XXKs5a7qHOo15M
9YenJW3WMTVR7Z2J0ZfZ3eqFdlEmN7z/3VEFHKEH73A4QIGuUCm+K8BNXZ4GyccK
F7jb506Kl06n3e+gmu84Xpu6TI3jMFfkFR+8fX1Y4CIXRLgH0WGkwolmQmm5Auxo
jpGLFgRv7JqD53cJfXKvU5ZkAiNlu9qYI8aGCFwW+5vgMEvugxb6PYAHoYXp19Hq
dZk1znMfKWcmqa/oO1A1M11M27OWmK/mcMoLAEbL/rVE0Bbiw2/KrQDCuCPyJCWE
9cI5dtxYSIHVmMsUKYdCIIsADeOm329piBsC/oV3DmI4NUb4RqFBLy5+MCkGunda
6BD3JwiC4e0Tmlm5AnrxkyWmleva7P0/O+FfLhwPG3t0U8YYXaqetqpjJ3ji02Jr
jymCZHEJFM1Y440bIoyjQspQ/zVHMO0CALQuPrYafmOm/vlmLfrKFjGPPjSz3d4E
jpDmDARfnPHOTfESJR5T2aO+FlWcrJrWkvBXkhJUvLKqajkjLmpd9SU4E0k510CK
D7w4ZlqDTKWmlBLOIXcPTq2bQn6AX2+TvDvoXVGWZyEj+XFp1qRJKt49I6gH4Fzb
tIyClJ5JOPMXH9fJmMNtASbTiWVeqP0zuW/QSeAOQfLn2qo5Lh44XngmqifnkXI2
/1dHHYMUxf7KjZCetiZSNcmm/tLL387IfUwOE/4MRSZLNWF2yZN+W/aLoKcxsiCH
Wld80cJvOHnZtNlv+wdgX9xMZkXPcjvU4eFc5rvADcQFc/U+7nVaivY3cxiiCnry
GwH8zfvuDCP2T+qo83DUsfTmhy0ae/3NBXHvwv9wKdsPKO2mnYDIANsgGv6A/+CD
bPu/vEXBTfCnM/BfDsoEnT/HWHMKuKRRnVTt/3Eq9h1bk4GwhF5mIHLDT2sWWIun
U+c5haOSXZyP/cgwaAk18zylDh/32qiFF9lVuy+J2AmgBrQc5cVOVZgMI+H5bjwl
NPCIYvdopJQ93GpMrc7mn5I9t5s8GmMMMikEB1oAOTBnhWUjPMLTOVel5AEXmWIi
fQ47//y3q3K8HWeogoaQd+lH+TbD1dI/TrYPIBP2KEusLRORpxffFUD6DWwXDpCH
tWLXn0ryV+puR+9HL7qLOIFscJe/qSPg2d4KB9I4i44fS8KgcctMZjXzenbykK3h
eE/tp20CpKYAMw0nFMIZBNHfQ6hIXEeWCf33nDLyeUR/dB0z95cH6guV0LGv0gvv
eWJzRFkQE0fcQAHL+M8e+LwgkSmikDt1+6oqRj1uKAMFU+VWrR+JksrqAs/fsmZl
syQA1O2dvgb3FUhTTqkPqOhz7UNY4iO+wYE6K/UKtPFWJRlw+w/cwWWTVNG+ajUi
GirlKUufyI6ZbS1PzvYmpaX3KM1zx0bwbCdiXWGbG9dfRyLJH5/AcJaw0v0q3D4E
4AMa/BZfVEUmpdtGGEnYwyAG/mN+4zDrmye2T9l7kpzlJCi5VAG4Mq6nbammny7G
bpXeg+djUmMRvgx8YT/7EcxGVyQozaIQRIphRJHhs1pTRLcrlnE52U582VEDUYYW
o6xQYnbYR+79RDseumr4WhgyR71SwDe/213h2UumsnNn2of2QhqJJBS6VYg7FzP2
KXlgRi2pUIXPxpbTJBcskZrKvd3eEtnxWrWR6PIMXYHbZoAyi3DoCAxpKitQbaDX
CWd0eQCBHI9JqSTFB5A8Q5j9waVw38slrHeXwB7Q2CsAlY8fayKA1/2Xv6dVcyoJ
b78XbHRPxMq1q6SiRgxCticsY7NS0uIi/4y1JEmUKDHVBqmSRdOWqP8AiT57pCHs
3uHhbpeXG937UAZLAAhEzo+gemgbZN98nRL4fnoHPl2TDc9EDyiqwwKEGu977z8P
YGkPmGHroKzjOjKECvDzu90z0XFtVNBRXdpNGIB1YMWxfdQBfFk5+Fxde27fbkxa
1a1uFxY199FxDLRgCsyJA31lP+Qfi6McknTihLhhyZRTbc7uvrlnietZNz0wMONG
ZVWf/AO0jlMJNas5LqQy/hqmghk5OLIYVGDoWpAPY+LexCjY6/HVneexYybhXujo
aOcoic8wvhVrDfLnE/jSlBUVxt49Vgd3h1kwxNT1XsMxdTvroV3HH1TwqO6ADT9V
zy+LdVeVVE6b3PkxyCyqDPyEHPxgGgzKnWlOzUa8Uh4KwK17nlhQThP5r46qdSPP
/Em5GBKDkr0EHkfDO1E6UQJ0P3hd1p+M0kuLOseDBXEmPjElMXhpnwert/WmPmb7
driqCSwtLq6YJp6FT+oMFe0ZYqMFqMyYiugqpY2o6tPTC1S1W9pu99j2+utiilTp
yDYJ1pXTwTzn1OibRGwQlzbKvkzAZpt8Pl9OSXLm5OpPou3ew9wjP0J75x2b8MVa
H4n4+CASuT5SPEp4P0uJywAMnyZdgJKKP1jyv1O/kXGllAeZujDOfblPhLlYHxHT
7hUfy7WyVG3yG0ijkCvKELRNtPz3L6RncvxekVT03LrQcZoaSUKGqzTU6ZuvcQAm
WkqY+xsj/KJrY3JOBuNUTfMFrr0TkImBQPR6Y9qYmGwYhXfTa7zIGRV/unKY4kU0
q3foUCiXi0mTqHHrReJLRd6WCzpy+jghLbBJFcWhQfdkPSutultlx6na+WLm7Rox
xay1UQee5+bVWT0RsuzNTzEjyMZib6ikY5RlaE41kn4kHR2VLxFhYzJg8Dn65VrA
wDz9VhDF8dMqEirRstF97aDo5XT7p24oNWSOI682x1XmeeMppo/ZEk2mdbFiPlvD
FsMnj0lzjVziB5vOPb3Oz87IXe/QXjZ2PGHe5+mqDQO2SobOv8cDjnnfXYm6zUTb
q8VIfeqKcgYoCrewfAYFhZi4e6CSjllO+ma025svBFDKoZrm75h7i1GdDD7Eb+gu
ghTTjtt760zwKWl0+Rok8bzrQ67Sefk0njkl8Ezt7eJ23kdmV2B73ay2oeq2ilnQ
uBeeTs3x5CjKFwTFMKcdP3jSA1decZwkubdMSG3iu2Lytt5Sise5ZZvFyB6NeOQu
0oOpy/c6QQNFMdbnzutIt3BjGpzvvEWfy1KzcvS40ADNRUDleMt3JZz+HSOHtKra
Qy2DXQynStjrGpmVHBWzdzznJ6QrFzR1aFCCTaV0fvFFm0aT9dKIcAMK80x1QjrQ
b3Ri5JT6rixeNAoikxgv0MT9bbEjua6BASwW4rngz2gBuj5CxVleu3+QgMTkk8w1
ZTBxlbKQar0kilxW8WJrnUSzDcOeAJX+TuIAhffpmiPQXQSSv/r7CK4xcgDO1Vph
VecOuHoawFD5PTPeK4XPUn53i6KN/32XJc4sGZU/uVFAZgsYULZfbPXvX7OEnHvp
Gn3PsJEpC2CdViG1k+UP++V2ugFUS6Knze+7p5hHR6HqUNlNR8/FyAwzlVGIW0oY
nNHUpbuno4lWBjDu8YlrUYo8YuBbxbMBpulL2jFYDQHH7xJ0hK8ze0H1NMgnKPxY
ZmrBOMHFa8JzgyaPjFU6WyR8L1NdPknBM7Kmy7Yoy9jIU0UBqv1eQjfW4cWgDSac
So8cUlVasvDNaurAMpl783Aq657SxfyltY7AfikG9VDdqj+ZiMdxY2HtJbKsAxtV
C0NPAbp3bIURURuyJUEjjbMLt9H59+DJz4CNo1/1txd0EwbiwxzILV0BaUkqbBRD
Qmv0Lq5KgHantuODF6vWg1IIwQzLNOa0ySOxm0kG+H21rVdphNE+2gQ0jJZXsMAa
hBHFfX4o2Rr4HsCbSF/B9lUkGQhk7zQX6wIQOG5YyoVwY6JX1bQ1R51qY99i1MAU
0LDoPJ9yuZ3ehIM7XdU1Qzk2JbwDUvjDuS/H/e2wWLz8XloA/0W4zrwd2OIX9CMa
54kaTBD7hFBSHH+438fY8wykxfqU7t3D7wbrb+39ydfAsqF7m5a/9go8cjJPN28f
6tD4+eY6o6j5pG0WgxJM1a46Eu+gogOcmjtvFk4WjNd6qqSTjmNtpZQKXhqPjcPm
NnyO2vpbUfmPMuQFdF8xHHadjbb9roeOah2V4s+x7sGFxxbbnBDbCurB5WpHdXhr
V23WMb2aTtTpEpTjy6TRDi9QNKZl1u1Yfeuh/z8+nMjeWcXU8apKZuir95RrNONW
2g3vRT4deWz1oASLcgaP2nV/QAFZA9ziY6PNUn5deg02S3CGRaYW7Z/AzLyzDnMr
eLHtGPotVIcGEXEATjiYmfmxJ10EGqNRyrAZHkaZzfr+sklVzPIlPamIi+Pbo1Ni
evhkU6r1A5hz1iqiDmYZd7azHleJlNswdWBinWjhonZHoyqN64PAt7AKfw87OYaS
sTU4F3yfRjUGomLm9Rki70xPRcN3Ru4uunOwyWz+1tMo9NutVEYgDbTn4tfBd9c8
0bCNreoEcdBan/Jn7UidhoOKJlTPfJavNOPsAWbwFPTtHYQA7h2FBUEUUuxYL54L
7iOTBysDKoXnUK2aIEDLQMZuTojqy5UHepF83vTwDCpXzByKRUxVJf/pWpjPF1G2
fEt1PzGMseJgT6YbmDzH7R03hX0GYCW9XH9eFq3ZaF4ihSh91mH3dkHLbEJtvNdd
Zo8K0V7RKnN+vWvBbUtJP03pxoh7tijCdd+Upf+2s8FMFIGLXtqd78krTFoWRSE7
mpdvmiFD7k5hoEWvTehnPcyX7QrPZBoKaOhNwvt11oWNfnSoxSqbqHgR/3SPUmnP
3Rsx/U5suMIrIOg4y0s6yo7qaTUxPN2N0qgqYALVtVzsfaETd+zkMLl94JOQTy9q
s4AU7emBCRa7ZqACQJVBvOSSluLPq7rOzpdZaEJgqKa4P+hmQ8D3KJ8wxGQrzS8k
0ZVp3UmsMCbJ0UbltM0/S5ny9hqcrN+cdDAp0qmcpMtqy3bKM/Zc4NQsJzNmfHKK
Ixw155Q/KleiTkCITm9JgKkjhsHOsyrYNUBR+DxU1VIc14sxwZvoSonwMYgvpZLP
TeYISVd6XdC+GcLkYDJyUGXcI8bw1WlsWuQ9ClhcJ0aLZsFSXxm1VV869BteDWpM
jyvt+TpA+tyyRspRV7luA8aeLx/5IEskdJqldaHY+H7l9Jz2tZ+4ZP6fVMLURRef
/t4T0Hrt56ktu9W6nu71FSA9o11wXoJ/6MlEfztOIlxwuiV58prefYBM3Dc+6ooj
NQnjAtt1yQdbLyndmQVQQYTPMEEN/cMtjCDgk8DVzA2ecooiBhWm7wBD+Jm4X7LJ
P2CAeOpcZd67QRTQRTcqBV4qAOY6kdu59Rt2v64GcHXpfDqiEsBLwGPrwoEI1mge
i1hx8V2vypaEcY4aqY752X3+q0Z4Of/5mrDygzMyQhlJGHHMgeb1s8d+DR0GuDTa
q8X0/7pmmCKg1aKWDKq2ZPz8dq3UAPUcWF6ajuJA/rrI8IGnIbQkQQHOtxaC7ixH
TbVyNO13K6Xxkk8dDFk1L2msnToyS9Y+eRoCH8dMI1jX/ixx+20A20IP6wq+UY0I
1uSuMfI0PGylXp9l823WetsXwaVTh9wXEuBangX0uufAChZxJ6bji+guEL9stc5a
Cb11kllwayFiqjLJsNIywboz6BaInQHVrxhkdOlFze0sRckqtKfmTM1mABWzcyoa
zSt0k1lBnXG6D0fxEg7RTRsek5V4eA3SDduB5kiuFCYmMb6pR05TRbYqIlk9AobT
wWSglgHp1WilO+W8LljHEb7+k+ozOXep2ov32q6StcX4hDcxA/7w7hPyCg/e3L4z
m8nqltV9/rJq6PKAJJbPYhffNFgHbeEmndoZGvGt+Yn5AZ6lsRN6bfoTRo2is6NC
BZy4Sg/TLAGyJRxnNZOb5t4b5OXbXlb2i9nWxiM65YxAIHXUDO/AXZaWV1CuWe44
PLIVhAocqf2Fj/foJP6220soYXSLBwRPNHYpDqO69sqpXZjf1kfwtMcRmIWpoJhO
er5uY6Z6mmICNPgrlxAsEpKNpr7fVbYzMpgCQtnBh42mQuhZvpUOLZFYumDs/Lm9
loKXrDYHJlmqb1nSahMobq7tbgKXC8HUc0/BumnHSMpUwRUzGyb4MahUJp04ME+u
P1hxHr1TYU1lLMQdKHRc0BFvSCtfn3EEmPvvDsIeBYmYm/67qgjab2ZX8kOF+HlX
zcHp6R0Tl0gE3r0OzB3VYRRNidtnrPek9Oyj/XK/C81zjUZtWB7rNIsfb3I4QsHh
USLemrP+hkjksflgPM7xW8/E03I2PQSq6FANODSUXD8HTBGV0x/cBPe/5H0O9jBD
dvFuROQa4ps1aopXA8W+acqgVITKC506A9HBqeY7iFx2vel/da0A9E6Qiue2RVlB
7dak+zuvTxvkK92DEb5phW6EStwmJdwGA8nuMvs9C/yNV0LvIXSZqu3rpkBL59w7
jsFhi/ATWa75DsxUzqoKBiged1kTY45qq/ntIkQbFpSqc/SdO5WmRPWxn36FWRWK
zFskVL8qtXE/NetancaAICFzQmKM9YwQMtkG20DptpmfSVcMVQVrbNvb9cmlyHJf
iCgLKbT3FLrGDbF8QwBkefTa4H9eyxNo+DiFsc4ImEBsRQHmZOyuyA4b7Rm12caO
jN0n9RU8a1miFx9K69Bv78TfhGr27zI+/k9kepqHLT0/jUfFsj3luldYIhOlKuPk
2S7NjY+JGA2dCOrJl8LzwTgUIsaDLCg3wTlL87sLXVzWZup7DgWCfThBbzQSnwXe
WAmDti0t/oIreEi8MzEMiI2M0RheHK1GXa69Z+IDCb0l/Tcx8/hS1xCmvQc2u1gi
2GIreLCDdmwW5IuSVXdwvYcZ7q1FazH4BWpo+fPjGIEJwy5yMDKcRUJGAgHHdyT6
OLmIRRfoBeWuJig1SIZNl9ZxJhm7tgXmTUm4TLXd3sDtX6A8hw9/r3/I+jAhgIda
N8YOgq0u4dC+0qEK7zJpIj5QMnJAfFAFUH0+Dls55o5ATv8bmB/12yqheRLn4u5g
gQ5xx7ehdIvXW9bMWsJyNucnfPVSWatiXUJdQEByG0X6xjAK4+9TBLfkicDoSbSQ
+1gzesUHHCtBK6wLZXeTtYW3x/jkY3lr70rJNZdGUopPtIf9H+RHEE+ZHDayM5wl
21Ms8ySt8PpQ6Few5mYxeFvttWMyMvSlVrj3m91XW9aGpHnlvHfGLlMDeZCqQmod
WsF4ruxpLXJvlQis59YDyA3WJYWyNf+WudEfdlFO+TPcsm26z1QXkBfr10gIqLiX
l8jueZbI7WdPoQDLZuqeZhvmHtpvtHfamTCCwrjwXs3QaEJx4BG7kQrA6yhZmaIN
XOe4vBHMh3OvaFKWzfMrve3gG/2su9h0xpnO4VEMXg6+TKOT4w45aGI9qmeb2C0k
hchKrLVykxu/3V5ZZYT0Uj3SKTnJBv2++YzoGp5hy2WObjLrGQ+14zobfx7ST9ku
lNetmDMPu50MKPvP0bmb3MESGkYP3QYD4gJWrxb9ZR+daY149syVIjTho1lMjM1d
uHBKsaaKk22jhrQE2IqLGpv5iNAA2aTDsCd007cv6Si/vbBP2+6Pzet6AHv9yF3l
QmGH4ubavA63twIniBh8eOL3ZYNLUXO3EJK37wle9jDN7orRxNiDAzxKwxBKeFrP
HCCmafixwfWBiRsrNCNSlEYJ+pMBNGvI9e5AwD18XmFiimE3khSVAJ0seTwT7Fc3
FLWvMce88A/5w1yraDKzZh4PkQ5n9j7VcOoeNvSojVvFXR8F+k6aujSwjuZuzNGT
TmTnINo23iii083ActW0STQiiV+x5OnZMi7JvqepKKfBT1AJrL38JOK3n6YeAuif
8uBay7rqrKoPBYcTbfFc5KCivyud09e72WQ+lh3hjV/ig0ha+PJuA2yuSPaGH3ZT
BVqDjL8MEnRvFEWF2RpH0xLdqCYPgyQEa2cDfei7LVBfhk20APcIq2PxTTO0BnDV
zBjxHbO8zgXd93fHIEJaXPWsFU+FSn8JXPMVBSf7dHGdBsCEfBDqJM4odxV7dWdp
UsaFM2CYi6FOVmefplm5xLjXa26nmQXVwxFoA9mNldTXWbXXdyoCXbhjk3nSN1pB
U3ckls2NL95BsroGfTmXaCuYJF2OrLnTi6DHk720tf2cXeP23+Bb5olQQYfxjUv8
aen4qvYelQ7sF12lG67mq/tYdWTF9Xd0isAWGPJzsqANXvHGIobEywMiLPvJ924o
Cjo8H79bdlMuKdAzIBt6HhlO+K3GJrIpF0jTsTa9IvAHBCvuFJeoFRcQkDNFtk1E
m6gFo5Ssax0TzInO8QUU1QLVa+RtXbEMjUyKjri5dGtzd+S4qVlWnr2DBGICtU/C
cgGx3rUSNiZJPjDrV9fn4mf3AyPboy54943PNa+8/3alXpGb7MUzdbrUlsN2TRG7
0AepcYnxUZU/5ryy9eEi9JutLgimf2OBxiXMfY+/dEDQhbydqtVLSzKcOysy3Hn9
ee/F8zF1OPlLigdAAOrewrHRdPawVVghoxvpMIlqpLpbWoJ1CuP7vv2mAEpTbZpC
cLQUaMcD2ciaBo794Ge5wvDWhuhV8fkoL0It5vZj/5SGE4Ka7Ou/U+kJPOkab0Xi
hUbaJK1uZm0zlJBVsbzzQqrpudRv7bbvHYQnaTwV96hZyjEnC8/Z9xBTuBsVvJYi
xhCMlnhnGUB7q6j34wo62tJCWC6OKfsxfZgFoTERQeuVcPxo0xBPtCHZ4eTOEWZ+
WxEr2jvPOVEiF6uUjrTsDC+1i+6/7SjW7nqCuJhsMt4/dVwzo3B4ZorIre7qibge
Z4fX/Y/AySsR3XwNfBmGgOmTp/fYwEVT7VPo18o3ruywsM9ZrglywoQNFhcPnnw2
P+khRJdlrA+JpV7c2cu3FnjuWUbGBO0BhlilDDtX33P9J8GuntWg2aHdtjtf0O7O
Taaz/zXTMBZF77l+7sBBqrhBClncZKp++MfnD9GIVxSzkyU5yBdUSvDTe3PbVV3q
KpLj7YDO+u60qxzjTqIvFH5bzJqRFddnypc6qWsqPvRvTuod69v7NSqfKtZCmg8h
MNoOfg4gBKkUR+gvZ7tN7Avlj+cigsYYj1jYD/TD2vParb4FnBLteqfJZOXRmv9d
Aruffc2uQEFlE1+LMaL2KyD2eI99w/dOZDM+CLm7v3HOwqF+mG9tRZPx7S5dhBgx
UluQQd3Pp3r2vgJzaNuQJAP/Ht/IssLWa6h9D3oZy2c9PQc50jZi3gt9CZRJKJVq
r/ZNST+mtBLxuoqC10gwkBKIkONVibYZll5iIPjIWMEVB+UO1Dm+8/eLV04V153k
atonTy84UATGXseZW2rWYm6uokCagY61NtldbaQVa+yhLd8XdLWJYDpyD98rq9Au
SfVtS9Oe/Ti+D5Ro+1oldF0sW3rlZKLaYuuTJ50yx6XUwBa1D1GyQf38OWj2ZWxS
MVhvTsS7YEjwHhqMqP/daJW5EtSPJNdDPL3X82m2nRl0pssyuP7dFx9AZzSHbTfB
32PWTRNLpBvmIRGxIhddoXyPU7srvwIFUdbO3AbrPC3mx+3xj2+GOj6hv6WgHenh
RdwKPITxIw4AXL0b1Dla5wSRsRkNKmH3zwkK1qplLIZhv/URlLzoXBUc4QclrLRd
b5V9RhMXsNdYldEArGmKYwtmAUzwq2SXdDWbAFlw8bd/Wuz/aXIpwAR27FP9g3Np
1kJvuUyMTIvQ5qFktcfmnLDYJnUZfnrrcDYuQAQj9vlP2lACx1zIedy75nyeHO3i
NWAaeeouwQ9jIQumXUOdkqV8Do8cDNe/WKvNvIR6GY3/sBOWRtdEd6sJJVBvIumm
zpg2ONcjpdIg9jT2k9Pi1RwvEbiKxqr/MGQQ4sd85WGbU/1EWxThRbbqMLbUtYhi
OcBTB6qn+X2H/bxbBE/QpvFc693niRrVmKoPDvJPCB9iV9buTO1PmyJZDdxoV8o1
k3eqcafOntlSw+gOAlQN0sDz/6aK98LkopM9+JPtgJk0mp83ZsA/hP04N80E9wop
FdwSnU+l19BTjguqoeGaqfRe5f/cHckviHbPT9CckCiyVb/Ec2r0iRCXhsGuYDuJ
j/I9zjdjA8FRBokov1Q3itLaAx0SKuP5Ke8yYyBb71NYmOu3SqbOChj9dvh/3AAT
JhxP2LuDZbexGEWhSA2jJt3tazL+sFMS9oyS4TC8/A9+tVW06oMD4Tfiq8tbl86J
2YjQo0OunZJm+VlkVAbNORzkGEgwh37PAV9tPBKfVqS+5w+wumMMBSM+yO/LgTH0
byuw2PH+Lmto4kpBEoyh3z6wMSPVX483lnLi/UR1qxiJvOokt/GgncOJaxUjb++W
2WDkGkS+X717D+m65XOH/oM+t4BZercEyjTGN0HAYGR3DKgaWjDg0jWKNyALi2t3
xrC0o3ym+CMKPVl/Erh1RGWRDmFIpqYsY6kMgcrDvsEcUKm30AcdresMllUVYuMM
BiB5zPFWP+QY/pHZUQuBUe3YjqJJ16L0eLGnhxDajpJ4OLxMxHojLZadye9lPIMR
fHRSZxDfYgBSjMe+VI4i4Ecc0tkCC4ZuzQBQ9/wPqci7HYReR2vP3cvGoCAw/zoq
0HABW4IGN7LkWqjaK6kYN3chHjKclhiDpb+Ph/UHp4YYCNcTqUMDyvxp8o2dtRXn
8EOqj/KvkmpLslupKj+BFyl1gT5WttBU/w6UDMrIV3574r0maH9DvGllW99cTGqa
xkD7sYm1JtQUv7NbOZHEM2uLQvimMWKRn5LJtc6FG0lAboz2ZORR1NjQoxyJI+6Q
jNLf8xf9Tw9KodZciY2vPeAmL4s9IlLLBwDJstVD89KxO0wC9A6t/VpaVCYmld1j
rWaGpAMLG77LVznHBQ4B3D7GvnG/3UlvOL/izGpPBoUMF9rgDDNJ1i8G9rhdiDDT
A2E9GMd7sbfU1Z2+amhjGExqJCDxyrSyIxRTJRHugTXxpBHvLcPW9prwGVx6nXvM
Eb5tiRn6UzXA3t7GUh7UWDrpEMZ4/Wh5LZdbgJqjlwRQLCwE18n8mbl8y+1TRll1
hX0W2Dvob14rWRm25ijwv7DZon66jbEh26QJrTByuzHXI3Ftu0nDKd3ZXY4Bbn0J
v/8fC7Hqgid/byxS2c9Z3Os9ULGHiZ2r7E8aQSJDn4r6IlUB4f+q3JUXoFEXW/Rl
YYwgO/gRzRY7hOO/V+zP2LQPFpKEXP/zYJcaDTdiKSt80YTQBMTVmMUQ6jhnsrCd
h/okrfPB7fx6zxMNK2cNdQPL/d4skz0x/7ZRoQCx3XX8RbFcEFu0MilagXo5Dckg
79963uttLZd1rfyEdFPpRTKa28QnOv8v3oTciXWR2XR3vX3q4NxNsvjajo7HTGzY
5+Mrr6cp8cdgmjq7vO0iNMfwLyufZ5TChbGexeaZOOazsPKs3+CzTw+GgNyz7bKP
F3UWKZ3bIje4xvS502HdsdgXKVe32PS/e6rhy9DNLy2Mhc+HXryh8xev32CnRm9Y
mdz7GQpgOgqKs9dUbaEXtqT82h4UAkgBICqtYe8yKeftHjBmu2wp8sIY3pw64cXz
cOsVW/mCiD8q1Q1pzEZ9BKNbnKmbTIioU1IVwEmuY6fXm9qk0zdfpEjlVtPgNyFH
TvwEnPP2KpXO94eeb5J5Dzu7mBhKGlYTBJFKcwFwmqJ2Es+plR2ZdDeajbTkL8uQ
lsVMW87i8rwd6+0WudzNQ5GTA1bHnMjXgFc/+iPvjNXlITpjnivStEf+SbDjIWBJ
7kESAw59FQC4rKy/1juOtxBSnegREYpJQeuFqEozVXQAyFww1I7Xj3HWP5lKDvJF
v4xlQ6yhnJhPBdr+dnD/ol4p2452E+flyHllFct+L1LemZHi9aPniDZj919+yYlf
HsBKeD4VvpoIPrYkblEeJwdrS/u346hML+OyD9qK6FMSdVH70t1eChnAul7icmV6
tq6AZnqq52b0DaE7x+Maxu8wAh1rhVfOH/IzAGUeyTwPQuJ4ZUk+kboeM2D+5nk8
gNq2ahdffCNO2xCSeC+cft8oI7A0MkyqmiRGOn2hGE/s94L2aP+q3Fsm0g+Af0lL
U8/IjAdJPCDcpuhPeX3K0MD/jyXZVfE7oeHa8ywJrZfw3Vwhsj2wUqw6GbAyPo/h
wyClEiZXgE0QGu2L4OLmdRDsvL3HM5lwNtoDs3WbWTwwDYXnZM4xaAJFeJN7Suh4
wwUizNA5T7OZtZcc0ZP3uEAbmKID3Q7fz+nATfnMfekuh9nmUh7PEuVPQjHp6YYe
3Wzc3kK8CrGnJpzmjHr2cgCaSRqgagpDxnIoVAPHwwuvPyT4yGz9ycq5pJV1xBop
5G53aoCZsqpapsw9VVAN9o3onBrs2eczcobiazmlbeXJCVjJHa2Ix8JnzpowbazE
2BOJldsnTX0PLdfaLxM9hILhU2zt+Q1/+c1un/Kt4KIgoDdvWhcUnxciGbQTawwG
PacP53ZWzWOXi8GFu4c2PVJc4hNMkab3UkA5bJwANuLSbu8U/WHld5NxAaBdpcDM
uKZa2WIsuSA2HYw0CM60Kag5R6xsF73esh4PFrrp2dYYONj8CDlSaJ5xQcBW+A0U
h91SKzBfKfegl48FZb1kJ8LZ3CpjQM7SkyxWR2gzFjTq6sBogv3nOC1U0Dq7Y1a7
zaIfW6mNv6lUarkCjG+7GgWY2/vJeDkQtrMB0t875IwQDRWNpjurB5clrKmdBBDF
Ls3aYpJpyUmmJkckFsU/UyghiYEnbZmZzFDw4e6yhQM4XuapdRmlKFMk2tk/kBNa
r9+pedm6hAAni6xFcFhhSj5bYfoui3ce9ZovdHamuHzm2ldis7uH5PAVO645Y5TA
ZXUr2xR6FxlfDzngm+dsWRVFTGUTr62TUky8k770XqJzl8dZ19h0W0RFc//ljtnc
k24KTPCxR65hMAkRfnwZz4cTzifAZA2wyo8L56AdWUBmP3VPkMPKY0S6fmAuj723
bVPZgex/n88zDj5twFVzTohHaRMlZ0Vmz6xOEH/nWQ2Y1HSp7oSyEUESM7ndCZxj
NpnN4USK4ONyYBFp/BHzsnbHPeXEHLpDsK4SlOvDYEgR4GfLRl9S9hzZxe2B5BTG
0lPOOWiAAxY/8JpFTmN2y6//QIvvhD3sUmlvu7cW3XjWGdv0jCSiFEY0EdwozGVS
QRlw1iOZSBUg34JMQitobUtt7u/ZEHMW4PQS/d7MM+4aNozXa8kupDTJ6ezW3eUl
L57gSdFho+EbVlZqT1F8SYbQWJRD8ESXxwzrnkvYr7dwJJh2sBUf6czZfEFGNXN2
bcZx/aC8LqAjBs98tVqAV9izTuIGft/YbWUFWO1x9wiVGnkO+YT7qkJvq1xoYbSy
jFRrlVrgK02cHW/XXz+xET3Sge88CK/+bxqQmvuGVY/JEvjsF3KrgbGIzXIGw9zv
JQcMg5fJUvvWYErFit5M12hbmufPNFo1iy53tmtxsUfVST6sBIEvF9Efb5ulhAOd
Q8tJH9SUwDbSAbV5epCiw/tZPenZYekEawiW+TlYOrgOvMvA94qQGP+lvWY28J0D
4KJoudr/8HnNXC6ZJMM7xuTITJYNzT0zxCBWUSkzyIaH2HJQUp6pWrDATsGXcPY2
NpKFz9DOTmtUhpezz5c72bncJj8CfZCMk0r+X/PEXUU89hSnjxNgdMaa3SzYOUP7
x/P/uHW8H99levvVk0XRyWBx5mGG0RJk2fGQIO40bfeD+lUzEEd12BFAyj1ymaK6
rmAJzMWtm3ROUGqKD6higlHM47e1nB9yPtsdQsbv6AHofHMgd9A9GBt4ljTS1SP+
P1v7OsAvblfzI8hlFJoQgtUnUpDO5eJWkH1PR3ovl95/sPuuKloy1vFK+z+bUuiM
IWGDmO9EM/8YOWKAhuxBPOoW0D2eNdciUydlC6XfbhRrqnDif+13Z3f14blUAJHe
+KXA8JHdK+nY/OK+dFXr+dQ627vkpOyd9s8Zsn2geuJxziobWeiCyxyKk3FF750h
NXh1eUZR8TbbGSpzsCVVUsGWseR9cQGqhsSZ5rdVtXz8oVEI3NBR+RwEWFXl+e15
5zjBPU3PBO1Hdfgi3psdtLTrVHL6jMU/IiNMgdCJa/HyOhbXlpWXspJsBncTXYxP
Jk9KQDdyULrMWBuopDbXJqXaxS6UcWqu1OzUHBZDinVJIozXP5JBBMDgfgA4fhAq
m8ag262P/VY+f2Yb7rTJtxHWwl0URQwnrWPJuzb/CLcy8Ljl83Z3ZhQNBfRZ0NQF
AjDW+cQfMnxJzsfOJevdFJGIFlPOzNtmb3I6KjzvTrbogs24DUqyxRYUlynd3MHg
oEyGMGBlq9onQEqPyvrVhLDWhbyC3BosRmQ5rM3Kc9XfbmWQSCXS2jwxOL9lakmV
odVJgfsPWV0a1WfXHJc3Ys9IcwWF7gb4Tadk4PINam+ThEws53+mjvyTabDSHhpm
5Xjxg/avRYfwDbGaX/LG+uYuAwjwrr3CSecHGQrbHnu+SYjf6zxHNhGzRfU51pE/
4UC8ddYzmaOqP3+O8P6kTi/nZR0/TQvtwiZGMV7FwhmywlXoKLxHflQVffks9RoT
Dflge7zkhHfaE0EIzeKGTw2gy3K7/m66hQkq2eXjXjxVTDow5qrdKKtYqV96ZCLr
yqTnyAQe3nkayaFwJCDvSLOAlFc77YUrPIHY1MORbB5Qr7vpYeO6aYKKj/S5DDzi
kNph0ozgSCRbTKyHpA/AQyQURb5/hN1NThxAMevd+m8JzeyJsrozv0ZsZ4kxBpRk
c4mUwXqy3/u6iRZnrnF58q+umHAw6ze3c1ZCiOIhcYb91v3ol/DgEo5d95mX6jlM
KLXAm4cN9yE0Fb1yiIzD5nJBS8NTmZ7GBIGWjHzHqPSSOEzMp9HWovaoJ0sDuOhZ
yWgv7aCw9VbBmHkLXhGCFz9dcb5AECrXak5uGBdezoKsOL+q1ToWyFYebd8txdmc
99TneGgQ+KsBVOtccAunbKADtSdUvxn/OPCwCQtYSZIVa6gWY7t6W5bGrD2TsO+O
t9048a4J0hFV57tOyMzTu5qJqiMfKL0cjVaYBckULIg87q5V3MZVB9eXYNHnymve
+dbL7TAmauvoaykV3/47f8Srvnu5uZYTUO9tfzX/P+jhiejiBG6SKF2+yijLxZc1
/n15cVl1kjrSm0yDfYA5ui8A6Uqn+qHktBwiHF9fkyZDnzajPZNjXeW4242+DLoM
BV1Ze6IHBIvP/9T5989g126WIbqDkV9uW/pRsZuEf9r8a8gXJSXkopNjEaLIg7eq
OKGUvwqN1C7+JP7ETjLiKdVlP+om0ZRWzIS7ugF+t87bTVtSzPvNzT+5XF49Jsqi
tT6+ihtG7y2g3gR73YnfWbW+torZR1OJsdExwbr4L/U+gVTDcVI5gAqOuFzMoGe4
UUKcHNjFTNqeu+kMMIAU+wn44VI1hsZy/4Zn9JwZmOqWhjxPIKgjV6JTaPiWAu1Z
K9eaYE/DMZwijjnCttccKIbVZzz2lM/1boezW29zvqwn5ZiSeNLbGPajHoc3wGSb
oHlkcgnsZmQodyK4p2owNXUD3O1cvX6kyQ8SeyCA+auMHQq7Kl+GhSxfCv9E3hfn
5+icTcEOLOksQpRMI+xnpOstlof7wesBmAEuVwDc2OFGp57Tz+M35nvq07I50YOG
oXaJBCifqik1bk2Wkd8YAszo7dmyV6KdLBTIsttJYan7cTtShN7Bx3B0kDP61T8m
avJAYEXtcf4xtXmXYp9bYc+Y7Hak/W91RyoogUdsHmK2IT/MJ1Ev9qTeL9m9OTNA
s33rNFYFeP3811yH97zHeP9S1DnAWjoWWn9Y3K/0bYn+zwbqoN9rjAzZRKleeGK2
UO2dftB3/fipW5aFB0lX97DJfdpmiYn9r2QAYXCRsJozfA8QE4T7odd4KEk7FMov
vvJkFeKZk38HBvf2TPj/fR4G+16UZ0NH59Tk5f8ahpu0EORHhoz2dVUindesaEMm
Ou6SLv5LLzuhOjf+ErRKj44h3n89NZqg3e7X4FmhpfKC15QG9wcGVzI2wUt98kGx
0AVZTy/dKnJZcDJfbY1Q+M9jcW9mLLLDta+dVBBWQav6fi0KdbMhzO4ZeORpuIxr
mL9DAFO0eWDweFKq24q8JyxOnywcJwWk1gGrk0S14AUqSYO1QEXh3rUNkQzBw+wo
8rvtHoeaP8bCnmHnVk/Eh8Zi4iBNKskdKV1LF16fD5tWsGlwoCr+lGvD26venAkS
JitE82rJsninzWNbn/cb7wVNm1bsf6oEH8M/yZMjHdh3gW7PKg1qHaUSGzeYveYw
MtUVVcOvUO8XZgLVwSmqZmH1u38eOMupVnljmb23UxiwBPcmJnkGVB06dfLgnvmi
Q3CqHQYimHsEfDz5+XGf6uvD+fVtN4yLjfHNQYhQtWJMhDVdx/kmbmamKQs2c2bb
EPkVywDI45PGTM4NbKvG/qnEjkfkaFFa/81bYIdnFpVjv/nQzlEORMY62K7l78fI
Cg0L1e0YjBMUfq/Py8hdhX9g3h1cfyjli09bZGd4PKivJFgH0A8rb0uduUERNMtX
x6YMagvZ5OGd5t6wdv8/G80L0nfaZNFpkWXyexGKkXdFePK/OrLTRh5dXnA+GsBk
BtyMazpfxs6DqFif+Ci0KRWOpdJwxL4AADL0QKBFbc0UIJMmQoq4oqC0C/QqIRLb
IGRCVeYfikyFqs13YXq+y6x+01zbc//fg3cfjrVGgIP3luWHf0roKSUaLc+Uz5Em
WLNiN4h6bDwbzcldXOoUAH9No5pNoLsy4+duesKre0y7xoWKHCUL48WL+8XeW3m5
JrkrkqY5quzWIbyaohOfp0Uhn2YqcG5ZPRLEAKS3ZG64YwY+hEkrn4xbgDTiLwr+
nlZYmcGAo+ZaO3ArUdla0KPuyXUGJjQldA8MLNJsCrnEfZerKnFjqd9e0t7Gt05z
gJ4u2oo6ATBDHrC1Q8YiLzuykz4Mj6NwgkWFIW0NjaR77xDJxXkJsSuItdaTQk4i
KMJnzSnKJUCGwm2DjMdZm/48DFC0XYVVFkFCcg2+bJpMLhiAO2QuzkXXNxGdHnbh
rDDFD2EsBIo9k1We4TwhkSvpinE8/v+hf0oyv5NYeDdlIz6dKXy7OXZCOnCPiDQo
IySGUJ8qPaP8Rzl9wnxzgNJUktpPw5YK3wf8KeTusxF2oCZNAUpNgqa95hNhHdSS
iHW/jO3aNG2H0/mgz+yopWztlfV9d4m4rfyAuvD4AZtTT9F22zYYnt7H3lxsL7aF
iVI1YFCVW+T2rfgXF9eg6CUa7+7IzVtAkDfwrwobU6OxiTb9F0Vza4REVhPGeCyL
wWnlVAL4TJ4fdfNy+e8acg4r7zx6QT/rtSz4wsajArWg3CMT7A2q/d0IG3H/08bX
hOBmebFWfI23HlCBltsbQUuInisUjCt++sh+FRc8iSRECVS3UskDTj571kPD4UoI
6ZFMZmxnwGVGVcrg/X929MGeaCnfDVcEXb9VcYn/vlCfNdzk1VIKPLJTk2Ic9IOw
kWbLJncGRu/BsKuOipTxp5798sDDGpp0s7GDN0uN0/9Ko7XJEVN5yDSkPXiIStVP
KYjesHvTiFwFTv/U2FZn5/knN9dUMLWBGJHAOQ0L8yKTvg6dxkltMZi3jfjVc1jn
IUk4FYDVeDxT1lljqgVGQvqjcgz1EZWyOKYI6MFtQUnhBC6hxiNgPEmwukAit7Bt
/CPyBPxnWXmA39PIFPdFZOjRgNi/Z16Gt207Ba8g/2BjxdDySKWA5ylU6tMd7QeZ
ST3dl6tzL5ZmHr/KsNsX0LFBQ/0EDGWbbfAGe7MzjpDjZj7y2aBEOJPktXRIENxJ
Yc1XIr2N4HlmyI5OuzAOE5HtSFcRQGGXn9qBzPSPUePiVPwz7R8Pm4qd5Av07GzK
Wfci2XumRMl14SQonios/Ad+Qyr8n7nfGsMkpjnfFx9/elLPiwLWzlLDacOlG1lw
iWy+Ryojw5L8IJVTdo+gVqH0ys4UdxRBRg6jgsQaBIn3ihuzGj8vTSIRvWZ+xocN
NOX4LJjALfzYRUIiZBWcV7cjHwfT3dZ1IrCmdF9dkeSYc7Vl9UfkR+mSNdnPYrup
VspNlwTQZPDGkmcsJBIKNvvXi7msepGrBMiHE7pBHJoVklHJmvPzK9tpkTOTj1ZP
mu9mc7BBua8CxK7LR1f14ekKAVKERllTfUCmrf1yANrPImm/Qjxr4FguJE5xSl85
1pbdVCsGPSIfZFn+Q4LnYUoOQhBm2OzQo7juDxlJ7wBQPLoJB0BozobYn9+PZ2lC
gD9rF1/YG9Chms9LiWODNPMmqrbCIw7j7XhrrY75RVpYj23vXklESNDOcPK+tHjz
qsUgqnCH05qveiW9z48xNaqU7LazYSwGOUcz90tfn+Il7Z1cJzcwkGVZLfzf/f/z
8RUndN0OjWBcsRkxpCAY4YGopZFoF2a/kGVsoMYkKgToauoRLOHjMEvkMTMorATI
BurvmYbqLD5nohk90CEq3n16hr18tzkOzRJsmK+uPMoPMwDJ5+pvR7YqvAvZB5cy
ONuTQJiESrkRMrPzRmYepNCZkayySM5VY+fToACNoUHDsFWsRudPnWusIp3+fdg5
8/KJKkFq4uV2QsoFJBpERh0H4DJx5hGuoWJb57CKjCpmBKgwm7dEE+P5BmP62Zr2
Nkq1isIbz7Ej2wKBEvL9vdaiMNq99Sw5vr012GR3tvyDfVhkNmHSiaWn4FWRcfmJ
Y5ff/LohAdTeYoNOpsTw54bLCaw8GZ5g2MuCtexW+2qqwUHM79393pTrrKwF+KE6
TspqcLMaG980iI/EwzNqBgQEkblXAA1c/aw7kbd3exeiYMxnRQE+RtjgMCqL8tjs
aMyLEP2xDKLC50PUo3YiA7Tb5KbLEEe0bm16nOcBk9+oQl5/AtptU6X5guL7X6UM
sAqO7d1UFyvjYUNXGxlXZR1vX2wDm10YaM2+hQ0RhNnvzfmT3TY7CWMhkXQn4DXP
P3XaHwXTImnNtQoQnlhRfDgfipClrUYqttV1iYvUWyIKyfJXfbhrkBsrD/W+m4aX
HLYVK3gd6fjKw5SyqNpEaZpsaMcBVITkNhqaVAmyuGIc76Zm7ZacZOGIZvP1qAjM
HgKlfd2+UEMLSWdTlZ1wYv5SnJZIH8FIRQ8VLLB621MOyKRV9MLBX9V28ZsLg1Z2
x/wvfA4l3brjgtGQUW205YxHc8hbEsyUd2w77fSqdstGhuJvEWu23f6uspYDKQJI
cD8OEAhchzDrdmWtHDy9oHqlXm/NryCk6+0eWzuqPHN/Y04JW/nEdFmz6TvuT1CG
di5L+T6h/WUpijXtxUW+xSJaASJoXbQwNFeSnbLnEtdeZO75wgqplPYNLmy/rzTm
ejUrBUXsceHxBiNvzQnQ+2hRjn/M1g60flveTzmIq1R4e13RcOHfuj27ukdB6wgB
PH0KvqzhPSmyOze1VRrH//q4kHbqxrTHmx5vmUc5uGmUPAWRAbemUfz4c9nKne7h
ttY6hMdM2NyPc3IGSW78PjsyAIUCGsclshYqPODvpZIUyvRh2WsdLDzoRUSZJJ1c
MAaWnQbyZeyu2v+t4hG6oR1iJoi26bbRXDHt8wIuxMwNaiEcHsvEgjWN6WuVu/qW
ZLGIrXwJrMqtEe7czxVobeL/1Q+vPxtGWZ3+Np9tFpjmex1kmJ6HX3Gy6kiblkfj
vqXmnEPDLjQ8/s9sCVPlCGfMb2FhSqK9vhxuXJiQRUInbix5Ep4FVOTk4iRRuS8k
7dwJ09LWRSkoFYxDpTzKenEFzBci+6hFs6z4EDCfkQ9FjsVVg8SxcYcbWVtW/Nai
lxmE9BNkRe1UdWYFN7fk8qKT1Dc4lwweulAMF9EQrUnm25yO+X6xLEL4gMeB5A7Z
K4kLX2Y5v2vyTwyKK3IUmP7rI8dc2hPN/YB4vHdIOGp3/bmHtFxi4T6xowgRtyG0
RkhPh6Y+Z76lrKUPRCRiojvxQgpBZoh/1Pj9euzhH6RwiXRXZOslRbOYjHLnBlQO
A6B2m0X85Y+gQXzhqAoH/Y0HVKeSPVpL30Jf8J2KdhlrublM5iG8rZhFL4Js0HTy
BmgNCi7VvxLoRKYq3g0DC9aYZbQ32e+IpOyVLP7wD+lbxji7sWCHo4t8YqM0LKlB
51DgChj6RhZSAo1emKTC2DoQKrqI04T6MVbQxWh0Ne7R+1CsoERQnpHXCtGuFBjl
hTiWqVsLyaO6uPfDhepGtSgbRfHJ2DQgGDPaFW/jUR1Z+A2KPT7z9fCN6N7dS7ug
r3CXQvuLomwLEp2m94x/kOhmvRWnRHBBaZWH+uLDTvB54sebtNO6lFC9zEYUQltq
xyePMcr8GmiCGW2iq3kAPgYgxnywZK2iB25sWYtJPRAFpEmRg8MBIvkVRaME/+nr
ni+EsCXwIhB3Orxn+icblVVgmiaeED5j7T6aLSzc6RNkqtujVEqZvnjdibJuP5KA
23R/pHCj1T3DaC2b6klXEOoactrCPToujTpuMh1rS9AjPGXud41U43pW5kFF+4D7
qwx+evXtZnDSInDYh3UzQuN9jtUf1pFqTwEFeaDv9m4helnLehP82iOTrEZbn0xf
25t2J+FGWrUJEdnO9PYJkYgUC6QhsDx9m1J7Szx/2aeVz1z7M8WNNr6lSpm8k38Z
SAExAdtyvCkxcPb01PEUrwx7iTdSpzUZHJz+TbPjkKz9KZgnsAVqkic8xU/1XGPw
l9PfakmNO2Xf3Y2CAwOvwyC3zF9OKg2iEYhpwGgDdF+k63I9nzyW/b+d7vkFaR7V
5IyPAG6eTFJvmYg31dHd3W6XdXzhlCXnNdVc0bkWwYqQuVLbM+SfEfWFzX3tvG41
kxYbPmSqXf5zQxxHj97cY/DpZUhcNVXu0GzTBu7Rjk4X5J8MSUkJfishw3fH1mJ0
xKCJoH6NMsQ6TGlIAd053e8QoNf7AMOKOVYy9gqLd+1HgZICvfebEeibqaV7ORl+
7EB29sd4BWysWmDg/d/tx2UO2yvIHt/KuI+0/ngH+0Kh+fqaGJGy9Y1uk468Vp2c
baG9djrB7jmRLBLVuGUVnkuIAB6D7Uea5RMV1YdP5250ZzYQOWXq+3fd7GeVYBnW
tdAPMD82SHiW++IjYccLWNNM99s0fIjHGn7T2cmLj9fgRiqahAD51NCIlJN7uiWX
VEVLY3fzNLYTYQNO68lu+VyKpM45vXDuIFlQYXSCQAPx5+CuJP+0Dm1pVCZ99wuh
gq8QsPAmNHFL8bXEtodb1L9VbfWnl0HelFz5125P0Nw4TmenNNbfZtEmPY5udgD/
cZKpHEzyO3qOwmPRsrqRz9krIfkKXvNZjlm+pcl7ZrHuwOZV9V0rfVM+TCyWkXYR
y9kHfDO7kIL31SBO/teKhfWW0pWdL0uzNoxqeE+NmWrOOmzMthIkZp1C9eOTiYPd
oH0QZR4gr/nINwo4oDv52+yTfcYT5eZkTTqXZXim4ZhJQ7Sl9+MA/ByxJ4Lzel84
oN/WfwKe3SzYDFuLPmUQiMxQUMm7JN7snr0dOC8xSdfauE9CGRvh0fde5Wlt9QEw
8vGQweJzDhfYdk4491MPFETd8boH/Cl+2t/e5jYajNS+0ogfdYwL4Px1COgcuqC/
ipfciXmXkeHPIMiD5Z80Igdjbgef1UH8tMaIz+vJ5Yd41/nZlaehfEDyrsltw06n
bJdpHnaRtKIJ9RvXMAoiJohYw2LbHSzuXaiwc1b/vg0naZiIiUBRqTX6JyfOUign
B4AnQjgS+KKUwyB4J758U/TEHWUujNQPBHPps8QzbgUJ8iPpyT1Jvj7oaadSfwA2
l3H/+omCh7G7lZCpwufhMoDHGeHDinc7NuhSPAO4jIhVMAy0sPsVea+oNzSrxYbA
l0XNyQ3zy+fdkJ12zfb36ZlKsCzmrNtOB0vpEM3ty/K1FcXvSyOUYhQWbh2qbc4l
i6GlflKw3IgB+w3GRSa0+lBXQn8T6P3ttxzoAFju+O4PwGQ3FvaJMigfNFFvaomD
Rt6EYC3qSvWFRkB8EUB3g/BStWb6wV/g/dnU1WxbjwLqX+JpmaGZAF29cW917M4q
jF+8p1JO/wnqUkRamo2+ENoFjBTdAMVTl2PP/N0Ysj7Q6XCsdGAgulov3lCogmjS
E2b0wE4uvZe4mSiUc2xeA40MEO+6mMeV6sfh0lBEtvu/BCrlA2RMsNnPUFBSj40u
pH8SZ2CSAod5sXigmpvWryFs7aaTSVcpXAaDln6wcSHFCBmZOoTvaiqLAKz6hVgF
EBeWhzjzzA8C4k7lv9lzHBfq85wWY8NATXL+wWwshNFUfEkAVGmwZmjEb2kBrTqe
x0ojnXC80ZNMmTzAuoToegcr+XgHIahiZQXRrFOXNs5nFk1HNA4mfRNERo3nQAWe
+b4cnnNTaVY+uR5cmFCpFx2+XPwLOw/EudNeGVV9JT9vBgVrzGnu2A9MEiBtYpna
kLHt14nzGv13irxVQbGkyiggsLDNeelk0kf5M/heOeIpSIthVPlGKu5BH/lqhMFr
/DIKspT7pH92fqeXgNlDcLlS/wEyCF9AhLkO7byFBndzxcGuyOLmKlsAXHDlMwrB
tl32q4e2swznzbMoQrcobH8jxbJ2NXTYNO9X6FPNwBTrflfATr8pNwTe+HflYWvY
kGkC2583XbtWpK3qA/coHVX0byDBC6A4ZJRA4X3t5WEc/cVzhkSrn8u1d9V+7eWn
ICa6mS0RrYFhLQibQkFp8GkfGjpKFOAwWKKNgUfWes7ygzZ9IL+je8EKHGuKSIpx
gVvZMUx0z6VDXoy32MX8puVFkKoYUZtiYddEtwo7/TC+KmWUXk1Qmkv7so72883j
DLYBMQh6+DoI3CQjkJ+q8CbYVCzEjX4IQr+hGZm3tmPnj1w5mBa78ZLthKmGumPq
OC/alEmfWqJnSTBMMjsvvAB9Hk+kWjk5dIlhaIJmikQzaxhvhpFOkvRxgTqq2pZm
sdDd6LMQyKZHcJWulAti3JcwY2VRHwvN5lvDcSEiEk5tXeZoXJ5hqhDHLMlEfd70
WW2WlRh+8CtX24KwvT2JhGUNvx/89Wf66YU11osA+H90JiGL8YXh0WHAYE2KFe9L
yDbpRD87L8RL7IHOBmcoy2Ai38ezSLZ8XvbDXqd73E/Cf4/d50ggZ9hZlQ7wN13v
oY32/G70xHCLweWHP6FkFNvYMEKQAmq/29R9LFKC9Gi/eXDQpat6O97ag/DN3cwG
u3zeWWks8lvd9qgZfKPU+gw/XbhY6wQ6QJuW/8hdfUJKTS27gV1WmP5U2PHoc1aP
T8qKFEeElfqoBgg3OWz5VuEqO+ArSSFMscO0WGiHS+43b3a8N0EvyaptEk2HO45N
HUL1Aoyo0ZYMcbv2hpRmuJr9iaHZJR0v40FcP2SGczxiATjUYnMzNlZUhUURMk4v
+GJJpzhdEq0gq5wfifAoLlKht4IV3X1jJwhB6lshTZ3SPPjuLwBsdxJ07vBiyl0J
DbB5HOSqlxnOIO9vMPAYkFqR1tuxzDAjAHlKZ47w6fkvO4tQflIGUEykFjo5mhsf
j+woiVrnR+T+a7+HO6913tOtcNVCzZYWkKOaDOv/ydGDMzlbdrvW3Ti+QwRlJ9wN
VsHRuDLRlmdYpyLgywEj4ldyCoyaEu2rCzScoDshcq4ZtNDkYM6Uh6eg8pdyk2uu
+GGIPtvk3jFsC5F9AFn4ik0smwJ5RZPNPv7f0dIjsSij+o6oP684wv9ycaBZyMAQ
llN2vk1SF4qkA2NEyHFm1nP0SKfhXSpVtG5yimyz7Jh/W/k7XBkiJQ63rqchYjfi
4pJnzIlDNNP4JsrYMV7/b/dwzmjaFrR+gNuwqS2X331he77qLeAYT8L3cXltVyIU
pAVm2C9Jx8OIC7Tn/O1VEXZxJ18h08LIpiL7vD4mif95fx3uL5KaksaZ3hKPceoI
85Sgt10EpRpSsVMUfDULRatjlCfZNIMrCwWFI1Y4JrKr78G2JQjY4AMe8W1TxqE1
ohDb74Vu9M5q7ZTOa3JGvgWRwk47zNEhKxm/PgHbkOeyw4WwhjFbO2gWOPVVwcQR
VSfEhfoFCKp/8srhDOMKlvI1/OSXQK2pNI1QPuzNYM4qNNV5EztMVyqVRj0kzwks
dTZJoGK40FqDQlQ0E4jhz2XmLXwWX5fgKPHu83b4LsxZdow5IIQzOa6Qv/bHdF5C
b5q4PHDY9rJxLDMQPd+hNpnusVhkPaHuOOdBqFbXrcM12AMgZvH3SoYEtiTduTnm
P4LIa9URKRLiTLEgeUxKoGfK0evoPwKp9pe9vbtjPr05cLNiyLMwCUG9PlOg1NAf
wCrzroQ3tt6I6gP9U0ypJxc6LHIfnquicsjAbs2mTMjMgiiJV+/CslBK0jERuoze
YN7gHffNSRwM58yM435IoSTL1IALhnTc6C0XLQoQrLqOzWAzvSWjT3kQhmNV0buC
QsmlPc0GUP5zPsnJJ3UEo3q1uQqAjwFiyrswhyk0JBwZtj/1e8DmTW/ASxC+Ny/p
xfswxfBOeOhLewXvoXSqICk7lTZBLn1r17QLhSdUXoAh6jjsfgPzI4TfXsLcd+EW
DmO6UPzUaMPni80ILg3e7HQRAaQs0Ko9WruCAH/WTTzflC/2lBS+1sdaZLjPDpDx
38Nq2tHwjPBhR4GtaMxr2lUNLo+HfQMNcWC9v0kqa98ptVYJEWx+6CxDqXMldKwI
ESNxNhRZVPscZpcw6YJkRrI22Ns3IpnINOJY7HOkuxsB+rG/EapIAWvTLYO7122z
/JEBYYhcnNzOk79LaQYSuMXHqyll7/BU2KTa7IHGL9KXHSDVINN9SEl6Qj6tvfjV
3H+TPVkmzjkn2Kw67c0eXWVYABfqJleP+ZcsRSJ/ht9i4Ckzlkjax4tnxLmSUME+
NkN5bIslvUCIY5rs8OBXIsJa/2YAlODXEW+x/j4jMmtXEFrzRXbvK9PrNrXCD+t7
cpzgYJKxYl4iyBn79jwbhfQ/Tcxhn0X+q7U6iyQzh4ZT99xBqKEBk4PrXj0krD9g
b2Boq0SftqgFNjdgl4DBSN7lUPBnIVjxqRp3ecg6JrQY00xAGUdWv0BwItmXLvxG
qGAwlDjgv1ehcXX81sN3emhx7KLtvwAZP9ZUwkh9EY0JxAWbUrmaUJy4GFZptnNa
xPmaDcdQiNMxDKdOkqueAymuPyzGqNf8dHYNKyjyB8cncc/3sIDBdnBFBQhoaQD2
6xqPhol8lGWdBxE1U+xw7FnKdL2OQgpcbnC3xlFbooGWYq1wlqtnisd+Lf582r+P
b7OWiyyLdeKDDg+SqnkmPZNienFzAodboyW5aOePl2c/71WJQ7QilGK8ePtr7/MG
1VtcR9NaNXDG9vHkYlJWMYSdnv38WdA2BZwMFYxzhpf+k4cz1iPdGuhPya+6eZ/a
/mAELjwUkJ03Rc1AV1mb4dYE8U4uLdho59kXN/lMBI+OhsvUAo1iv001XOZG8MTb
219ulGF66h1XQHUfCTF4SvEgUwTJBoEUYZdOBxeIG9pJjIy+aohlJsI5et4v5Y3T
dXHu95EcdcJKQwTyapYBi+O/aHDmx9lsAL5WoxnV9k8LADJgqcAJzZfOclBK1LuO
0HpsvICOW8DHvi1GounV7oC4ucUZnQrKi3YVyDDp1Gw0H3U3nvW5FQIXpM2wJ9Gt
QXledDbemKP4FUybyX312z+iwtyPnG9W5wJvldnHDc5joqYjQbbn7hnLxWgR/8FH
ExkuwCNAuYiUK4/1Aw+489F8h6RRNWIorQQiyKi/lYdoqKibCv6/wumBX8vxDYEt
L45kOTvv+Eq9iWLKhBLKRURYh3+0yySjEQCtScvelMSY+QyCzjGAo9zE0g2YR+6o
mc0lYym8Lhkb2KxslmnVY0H+bFIxyEBdtlWDf+e2EdK+NhnSUdCqqJ5dfCp/IvNB
nmV+F2S7yN44K444k5yQs7/AfAyZoMJRlvRyJAsu8/84JvTR0w6U9c0SmX82wRkI
pTRl/CmNEUwlAi92Bw0cSncXks+a3JEx62ogDRywQrmKLMGQFSF3iXZ8yEDSuSBo
62uRCX3XTagUuEwz+CHuv7S0EMx1KXM0/AQ155+BlHupBeT7Bqt2cMedR2kS7gfy
nIoaNBRZxXny7GLYuRDmEbGwx8j7HS9jVxjJfeTZiA2c+W3Mn1vwcmCPvNFr5iV8
GMCJPTMEixsNyhg4n7YOjYEQ1jhC9C4PAPFWN3+9BOSpJYcW1YU1SS09A4asfJMD
2LQFjL5lM5DnomQCfglJmGnRFMzJTTwqhJE1Q0wC8xV8hwSIOpANY7RqTSj/zYeZ
sZRGkSWD7h4G42ykFcQAwRfa9uAlhl525NGBJ8Fcjt8O8oaOPRWWG8XsdMCdAOE+
O9ieWaeEL2f1IQFjxB/VAGoZBrFou85NjdpVI0EkpcyVfzc2rjZ036isyLV7R/aD
nXwJurpUr4xXwEKa6QLJFsVYJgkj3em0MO4e606G1McptQAyyHXP7pAI1pJ+S4fa
yxNTBXVki6hprvGylYWk27kLEgJWgSev/TXthK2IDzJiTGEQRpDDDhA991yUD5td
ppXBZji3KJuEX7KybIO08hJWGcD79vq8ndZjJ0QQJOJnPLPryXMy3aiTYVjPkrKx
Uw/6Ag9CrV6CAPxygCmGiS2heDSOjDsEe2/LyzviILcp6nmIwW1QPvTAnBcPyX9G
91CvPcOpz4iqmIvft2P50n8wR11P6UqSZpsjmYv0B29sDJR/YjsGwvxF1m0fESnE
2xf+N0x0Tb9HoLed6KbgOEyEM2QKiRZH3Y7nBevfoJ3XRvdH3s/iLy5sf4eymvwJ
eMNHzr2RLOZDn6Kn6CxuEoAE/RYKbZcf4jJcsgPIx0wIOjctJIyKLnuFLhkp/Ny7
WD6x9gSzRmF+JLc9qNi0Q1V7qQ9+CKhDhB8yKuRKnz2F872YEm4409mF2WrAhr4i
n9NUeT47CXcBhzxQwf54dwx8uTggpO4JtjMXc9I0PR8+5xhukmcQ+5McKVWILunD
ENWvIlu51JFmsb1QTSjqF72JMMN6Xu0mjAfNPsSpDD6rRdK3/MytRe6VRU0yhMqE
tUGlvMGfRzFcFOzClmRFv/e2sh5TNjcRQ5B3SYAJ4/rFWYCCU57oAJW99LPPYJxN
dWDSFsgyOOytTc9XR6Lxe64GAqAJPepV11Vs85BEDcgN9vmSAKga+FCH0TG3hLwE
6lgLiub6+Mruj9wuSoDRQdaAT8xCTVTpr3vaz0uZqd8Ev0U7Q4YUyNEQzwiBMs4g
yQEg5pZpyod3TRwM2N/EUg4uwKaat2RuCqExtSxCMJKx9FTWwt6g8o/NgAWW3v2g
a09pWLRV3S+GbXmm/MxA8GB75680VyibU3f/uJ9TBsc/FRdq4Vjj9ai3vebZ2+LA
1sww2tkZuPa0nIXXzOPVZTjlSrC88Cl8lYNuHNWy7gPMgzsKTqPGQv7ZU4dvn4lG
MfqP6xHO1HaUNWSroR7stFP0W2YyKX9LZBKPL63a5HR5snjQHBZaufGQKVKBq20K
208vUSZBfTa4r7DBc8OSiTK8W/X+nQwAqwbDEx0uBjBWRO+pZJTnFjYcDR8XMhs6
gqwHjUVRpXICsvaSz8Ia+Cr+2LmU5nHoRWOzE9G9+cW3wLNbyY8GP40mP4SuOjYh
yZcW5IK5iBUKywq8HAH/0ioAqzTrB4UR1ZPAksGUH8CjtqY4ih9Hf9BfrMOcBbbA
M0G2fSfd3kmEMtmMQtZWs6A7p5OSSPFskw9zQ6dI6rsjltH6yINhHPw0xhmqPb9r
NzqmGrTsmLLekiw2bkRkImqdYIcN172iRxkfWnLz49VftiOZ9YTFMP7BZ6f9v1oo
kn4d7CxGyTB00dvk/6NgzRTMZpK8yKYKRK76MNUiY2HM9jj4S4CCjAXAV+MGvLWo
0atT/ZhuvmzxgyF4Jlh0DQv1S9kbN4akwIXrnSGJtNiShUvc3yR140AHAEtk931Z
Zb1ukGSGyB3fgSSgrZMGMLGfMXn7aeAvD7XtjBMS16ovsG0OT63BXn5xnv9m7aM+
WBAR/IvRJISRmH5J9mAYDJa2F0FyAD4/oqCP+tEvCy8aC2d/qqJKeS9UkLUpMMX0
eoY4qg716iHtEhZgPnA0/+U5Defcas14DkqGU7AJqkazC9NXskvAyuKshtJRxVvC
m6EZpUoCdaUz4QQCCCQl9fcDmDANPWnrU7wk9A1FQ6eDZkapsw6aNaV0KVZze2uB
STx9qbE7BbAFk5JBTLGX2O4XSAUAaIJYrNbxkzL/0XozvhZ5NbcbpdghyhgmB5jp
GF0qd/DWxrbXKMhosvZmaHM+g7de7HoQtAYyoO+VhNgQ0fNDiXcxRgRR7yyDNjeh
jvxFRKFwQVOBzgnJ7lhkOOfPw6Yaaatdx531ohYca8IKmFj8Ku+oOyzyePHyAjtE
rnf8iJSMVH62KBTAbpjVKRGWbEo9G90tzS9Q3Es2K8CXYHR5N36dwF+F5lAPnoT2
4ctnWuUtIZMIirx4ITWaLywt7E55hTKoKG7iKizhjCay8AyPTsCyj4ZFG7ppAC4k
39ih75iMavbH1qxvGtpQ/raWIRr0JXgtETECwj3oszk/O/iVyl3nFze5myN6yfaX
srqOD9LzM8RKQPjh4Td2eeEjz1iIWM5dcP7akjLl/VGZlKZrT5GodnH9xxFyVOgU
YKLiVSQ4bxUppxngabkiM7AZ/hX2eFCosxSEuU+aJgyBnQ59vO++klKbK9IFglLc
8TJgSgJJrShQHYGW+rO1GsKU4tSrLyUrIQ9iFs97gQJq7YPtqhlhUvWDuzRH6RQB
COV6PgvlocqnbGMwif3T7dd2L/JHQWPWtuBNo3Sd36vZGwJPrf0LZBsH3WFkGhvi
RfJjaKK1bI8Umdvq9t01fSNdGjbVKO08ZmoDedu29BJUm9t1kImIHC93OFNg0uVm
uPP1wQSJ5veePkxIVBWFeZ7uu6iTlKQ4b8LsT1TcPuVWu9OSU9ohEWKShDs07QF4
mxHhRyst0G+gCeFhJs4x3Xhi1de7tsaExFT7BaSqnoNChfIZYw3ChpxKbjs5VTvN
1IKJzo+K65avYcwRdhH21WUouUXTMVGRH9bo27CEGiV3dDjUUYUFEDxZb8u9n1uT
Qe4++pOXwI98hyTVHjFRvBrqRjwJKKM55jpkMIScPzut2qWbQO4Nr6pacQvUGrQ4
EkS4n/D/7emqGCUkkbtirweO8mvzXs7jqwMdSBoyQdXUyizO4Q9jrFS94aAlRlW3
bV5Wyq/qGKfKvfHNXeq3qtaF8bgFZSFd1G7K+5lpHMqP7VQw5PnQPbZ7BRaTXsti
BUAt7D+9VdDIW1s74DungmF2JkINdvXJFhB+SqKLVT6WkiVo9Mx/Gg3uVnZ7AvTm
KFRB6t4bP8Raq62cgWSLBvvHmZZSkqI58e4q80csg3fBHVm3/ecckEVUTusNWj9s
RalaYjG74ApVp2qK1C2hfbtSL11ZuiHcJ1L9kLVxdYxeFbKvM+2h/nGCJ5gtbzCc
owRx7X+1mWv+7XHNmIsLGfZYySYX7QIH6bUqifqYgabGxcfgS9sImBlIbyuUWeyv
S7mI9xSF2zfALjpRXyIJBWtG8kwufcuEcjCrIzysO1bcVaYmRDqx9iyJjlqO4KRH
tthmLonaDJr88S+GcjwT4/xwWbkvYEgYaG3Awbl1VPoj1djgmYNJ+y3bbFSgdaCZ
+TrVfWOWxzjY/z9VzbKWdlswBlAOixZEZShHcCKyev31UyWOPr7z89HIqNwwXhwe
a2fRubjmKqnkihNS5LMQQy4ENX36yYVi7Bm/JHPcsC+OcnZ/yhWcG2bGQiyO7IzU
AkoT6IGEaNLiOf3AgUfJ4XiquC+7udeVC//fcq4DyT4pmG+8qYlsIkEC5xQHGyon
HmMyPBELVtak7Zj2LY9IO/+R3DUkIUotM9jfRDlQ6et0jjqPlpYuT12tXhw/f48P
BxeZ8F0c32vsw2CrQp/w+G3AWuLPnpcMbAvRydOq0Y0ynyxW0xzDGeZginFGe7aF
BiYFTGY6ZZg+1lEsFpjykAXr2ZZvHzxWWCSEZWElE6g5+aaudQjHTMXGTFeMUUir
NuZomgcytZGmPEHljsxiAp0kYfwWDu90YpTLZcGh6XbxCtrATqu59/g5QFFlGgql
ZnW/bDVQKaF0akajZrY5V9uFcYPHt5lIbBOw0a6EYOogSGwUIMZqCq8U8pO7qi1N
S++/dC4FNzYWapSSgpkDNOzeM6O8XmKSlg+AjUETR1ozztn6Zgx06/sSbhQQ8ohb
rg4JAF1KDtQKGo75I6SnSgZMeNycPm74od8fu7TjfeDOTa9OxLMpq+pmfRpJuIMy
1+QNPQrZJWEmON8hIiNKoaiCukwv84F2zehMhCwr0n6tqoP1F8w8YO5A/qXyw8vA
QXycA6lmO30KMyGzKkyaCeWjQmJJw7IvFaLLGLDKDfqDnN3FChiIc6ordmEWz1vK
Ksw52wFX3/ONogOZRTYZqkdJQ5jf38jNurOzdmuXYM8/2DhAZSQx1QS00RymNjwF
p9a+3Y5Kla/lpwAQnlWmxR94Iark1NfCafqrgkiY/tog+d+DqmqHf113mb72fzFs
9QLxxM/eF5cyJ+k2jTwqnJSbabmq5GzvBYdnMUajis2ZNqoFejbQRP9IXrbKUr5T
NlxyfQjIY/LHbxjBf8No+LkPMevGUVEfnNm5o3AvRtx2CPFxVgFDpckrUbsjkIxn
spbqxTGYMIM2gRnKFyRyY6GuUSUJ2fcUFNfyVJbjKMirRW2T5psF7vTj5TA2/d/3
a9hq6vS4NPbGzuW7sz6h8rafJD8h+IIXz4hpmMY/ejhCttt8/JW5jx+CXiSE+fsm
qhgQBDvCKL8uXIv8tsVOlzhCAXJ4+ep1d3IAroseOcnBnXSfFQDqELvuF8ACZ7k6
JF+s7eO2d9B6n5NL7/CD/snHkqOVEG/6/69koXeBz3q2mpChEPDian5UhEWZH4xD
BGPtB4Lab/3XpPj76RdVKuDLRM/x2+dHHPeC9rAxtTyvZluqS9Wre6xSD9wkgnVu
5maAH3yQZv8WfBqS5d7Euflq9olF3fE0WbwTMtkskJtt4rQB5qj75bXCWhWGmXlo
M4OHOKlHTWU7siiJhbPFi/BRCWz+ounHJ1Xf9T847b7NG5XTMgCDbJZBdoGYVB7z
xk32WZlsSkxx53VfQ7ylUWL8Ih+tWJGDlWjbjcdGu3f0oXvCABhGULIChXuuP2Rj
Jg1ZnlSO3OFDQJFmVv+AYDExtQZ/OyXCahL8tguWUC6EIgv8lCkpicEZ3Fvoymsb
bC+J2HTifTBw2DyfjT2Ep3NWr553XvBx9KdJxA9DtRMczLER5/3DBOnsswf2adai
o8yyOYIW0qdiHOZHjChyzPbuZf1f2LL79Kr1g0bR6chX2P2o5dLNretjfG7/NWto
7twn+onqQOWvoHY0Zopt+/FIRr4rSBmR2lYbE2cVuRsgQpwF3mMfAuwWcEF9nT4X
b8DwhiC3LQed4MHgrtQ0Yd09BKN+xKIatYt5I3XdJFBpLypVTUHSi+51wvK6Y+48
9UVhndWKwxDh5LPRz4HLmp9RVM2vz+vElBC3SQ2qx87YKWFMwEx5t1SrVvXmbp1D
SMYCjXjOYJKvfODrbhDOBFFRupJKRFpebHrMhZG4zXEW2wok8HexQIwUKRZloRxn
NPwTAGv5i80XBxmMpAR/iyPNtPHEHzgze8UKkWUVhGQmV8mju2THFPn5RclH+X//
NHCgvekZTvRqQJuWjfGlF9Yhn4iZaYab/YI7qtAVxswTbZtFJVmCElALS5QZv5RP
bQdPOHKXIPlCzmxHHAdoV08xbXatMLdPPgbfp+GdCzZweU1PPj3op0PBL88KqiQJ
9swpQgyRwTpqHH5p60T2uy1sz33KlQ+pINH4kNS1kw8q3WP3aBjZ4FvCWEBOhPJK
m9zOVl4PMQ50GOD+QfFBbI3DYQZWOjrlw5x7AMdJesF9LcLg39qcd1A7RAg4Hn+G
1+Cxqc8KzkupH6MAt7OSllVzgJjSkdU8YG5eMfEmF7RfQ048WEeYpCy9TIKjGwTL
7c9HbWpvCb58+vBkWwBSxyMhFSqKzoWKbj09UN57RwgVrw+NNmflZ+UgT7gQKnk3
K5SiYdvZJBVa1+HkR785+7EZGVBq7qZrNlAbU/bONtq79pPQ4oASWM9WAhKjtTqH
+G+REsnit1QmtNWVcboKgP5g13XK4ocjjZsfotyV+0bLXsOM0gUYJ+gxZatlzrJN
cUDgCIBPt0s7IyaZ1ch1JfySVxfQpgKVe0o1vr0QH0NsyNkUwHSwhgRweei8A2z7
IAPDGq2OwNLAIeZwq0Zh1rLZOQKqQHkcOVPNwOfJRP++gG9EzWQG9BDsC3oCYGVw
m3H1Iw9QUec6dtN2s13as+nawhYrfj+OZ6hhT9IkW8GDDCR4HXenpu4ohdbDjxIY
TLSOBSFjR5rG0EBx/uOHZ3QoxEATIDko/YY3lJmuiC41KYSm8ySq5+CfRjv6vrL6
k/L0DQZ/QGYSZ7vHbuhAdfN3tk6XHEp+Ep15dhGpuf43wZXfY0gP2ywNBcBWxQA8
BWSMcjlK0h7VzQuRMxPUbGkPwTShzrwiAPKclmOUz228wN7Y4/SaSog/uwcYR00s
x9TEkE+W/0jM+9f/SamU+zALa5HjrE+lCvENZKhz6jNnlTiEtbw6C+G4cpvksYJV
m/lYhrOIHvg3CjEoaPqpn9w8Aqh+AMPl/6ykcnwenYwnbhkr5tweRhH8gztZuroJ
78cGluXPRa+LDSZNtKy86mhpPInPc81tnxBV1fnMOBtcWbQVpqvhFFXw13NaEtAR
Gzps0gwIvlnZ+9L4bcRNN6y3UT3uUT4mpEcg/PB9PYD3l17LqQ09b+xZ4TEXyWcS
1UmjnSzjk1zQ0RCQTGnYZyH/flaBcIp19RwSNhXKS7/glww4nnYF9buKicegKWle
RKYU6QsDq44bzbWp0Mzo1/MI2awQgjgIZL51m/CMCKXYZ7DHxwPWoZ9eVrv4x6ht
Y6A1t7luZ6sqIrHXINW/4JRxrV8rLCOTfAIQo/at7kTSFchcBP8/e7FEQBa94gZl
Kdc8pfh83PeTto0jTeOhWeKsPVm+73CMbXhs20zMQqD3ALj6ud6mvyWKjKNWp6+j
VSJdAiBm349RmKWcYZ6ofQ9HbzuHJ8M+fisiNi0udPbQIIlbINO0+NEejGPXbhZ0
QHfaUPzU21QKXSZXZuJON4C+ujnzMsq0G5G7HDgK2JniI8RQCKlkPfZPl0w+d3S2
XiqQpET9L718lpainF+tyd/NA0Ej4J/V3XPCEqZMA7GlzBhEUMgyfb9sQW90Wp++
+OFLk6hesb0X2u7HGHJsseY63050sVdJvNJfXHiOs0iZ+VUsBnb+5G5OJ3+l7bGU
kEL/hVXv+DxywOuo3H/GqTKWouCwjTnQ34GCbWDoKa42boQepElnCUMbNQZDyctI
mdbRsdVq3j2raOgj33g7jbKWOlYOsiolC8TNSmEeSXc2FYTM4qc8hv3IkPCd0DmD
SxbTtxqEVi/MOogD9XIbfOsUO29YK+XIbTZa0DCoK0z+cxqN5s3fBmLtZBl85N0n
1Gj2Mf1bgJ4QElkVVxSKnkdGqu/rN13pzb7EpX5ITNeQyNq9aP6IzWWMLzjOrBdU
xpcDnYXQPEXDntdv/DGZlBSHwpCLcfkVudnMfY7pfdhKAtL3LbGOdy5spO8XBiy8
zQgRurn8pnIESyfsSubfvl6ddIjRPqfCNJnyOObcuTb0Qs5F5TO1x6LxCkrdsolq
baA+iidGienMQIsKRsdy6rgLyCj6OKrm28lfcvrRumqlLfosD0REtKHtEuAOKz7U
NGivlcex3/60TRUOcOphurjeexFrF1z+bWX5KDGOC0mkoJFxMIh0MYCF6zL6a47m
LzTqRGDC1sASHTSSIWM4kmOMHIXNFb7oi1ynIhK78v97SKuipEkct9OvhZZPfLNx
3Xcq6NTXbQjk1u5W8YOOhTUqI9LFJXYIBuYjjIfXxMCR6D7USMztBmE84pzs4iSc
/G42X8PMo6fV2NCUiuDffmC3n7qbtlFgfnPGVby+JQ0NvseyJL5O0tnlcX1dWHn+
635jTH982kIGtG8zceQFOQXZ3Lio0W3gWnj8XY8B6Mm+ETmd1l5m3lh/J2maQ1DO
Biy17TqiHFH6ivYijrTHA30Wvmp/pmJzcPbW6Wc30ic+xq01uBASbJFP6G+O/r7h
qNi6gyXKqmPqKHKUVCmeD+Jg7034ygEEHhP6X6T+H8w31YBNYjjUKKylwNK9KiFZ
D2MJpecmEdA4EkwhEjvhQb/GsjOObBA9Ft1fJU1osw/FaBU1FBODodLCx86Z0usA
vZU2x1xMI0o1TgP8V+XhFcf5NFl0jhc9BtZINocL46IohAOkPi5lZABR5A0IeFlg
ZSTIjZuDq8/rdStReHYt6naXSrsXBo0g2PDNcWHy8mT+DR/N59WPtKws3Ij/jES9
+LmY1jdfWmONIT3HJUlVTGMPA8Ds5a7B3DQJXiCMKNzkrwSNRQwNLqQP/59mgAN7
RETUBJ1tfiqHQ6jlOHY78tGU2m4Hz3tv3oNeGiSWwo4nOWJqUCz+rpFalTEFL55w
JKG0BTCp2+epxdLzE4bHZlkpsgaLzZFvjatpJddWjA+yrD7WWEE10I4NQdPbm6KB
sZf3nxNG2Y6Bhs8gr00zOEAI0zvhr4AMcJS+cUnBHUY4/ksTF6svu5cd0LNDvUgO
Xu792PNr5Jc2zrd0+yWZ0AKmaiKYu7aCc1b2v8T0CyJyMcSKJaozC7ZYjuiqxAq5
dM7KlYT5BBCkD+6HkyVu+zr+nVS4FAjMIGlciJg87ocDp9pfvv4P1l7LS2dKtYl/
/HEyJsZF0wfj30+uMz0KzDNQT2q4vJtAmZS+ExkO09/FRuvbnHzdmlCGbw4zSDqX
VQEctZ4eH0fLfSeINXMgMF9aTO0cr+Ilr+MzmqNEoJDgOOPyDi7d3OhZbWc/wKk6
6pMhZHPMsul6/C4AF9nhAOhyci1VmYGruG4MUwOmbDM9N7kKHkKdXDaHlhMtoBXf
hg2TSAifUfyI9Kys7ytd2YlcjdctbaJEyemPWRFWyzCHxtLQJsQPo9IqLBOUJFc1
bzcSgTi9sa+9RGUaZv8lFvdXqCea2HL3SKNKQkBXj6UU87qHumVfuJJoZSpAWIXE
ehMVUzXfErTikCVmYHFMdBqTi4CqdLcyzBlTTxkdY/rOiz4f5FXsL+1wLDphONqN
Ms2Nq6PNDJ0UGyvExd4aBEh86xKVaamWlF+m1sSS08kVjLIDvBKmt+4hZE8o9xid
NoNioaUklzwGcmp8nNpM8Qvy25ucjxWL1Qrk3PW3kn87EYVkEVqSb52ly5du4H9y
NCDnrWoyFWZSJoyO+9C5e3pjS1z7XVr4Tyu89sOdn45Hk1akkmjVsCKshY+RkaIY
oolVwFoZlAen3qdzxGvF0YCzKqR44MnpMKa62q7GekBhbVBzRsRFJCrYG2Ok5gGr
hzFPd4SlPyRcfU1KduFdYDVoMyUUdhGyX5WFT8Zhs3bVMGXHdBPdxrh6MG/Peerp
nB0BPRwRPPoUtZ89r+fqfZFDkfN22osmPXPnzcysEvfQ9sSW1tNN4VRt1iwxLJUN
npl7QLXMqcNcxgjHA4DR+L/v7Zs8y0m/TTjctn7Lgri5UnRsmiXBgxEOoK4D4lq2
6317F/quOMfH6uJQqWnCuCqmAWgckw5lOmsuTizrT97dhxBlktgcS8VWNyWc9GXH
G9HDZkDZ077MTuGTFie0eZx71nGrYYbgINcbq784msMkBu71xmTtxtWYUGxwcEXq
90LRTj6VUWvAa29HvddS2egC/KsaxMbpBGLF4kWyx/1Z4DJDfSWMXl/0tBbU8iPB
0GYvXWmvg+SDG07PCOEM0oJLR/Gbk6plyEHD9Z12CTcqDsWPpRcRp0IId0oIfKrX
2/mvcBSl2QFqiGWYbH2J9xCB9RXvAFmD55vOlIkWw+iHaFDJ44lX9A+8f+tjKipr
5h9KgKjbE0Uhnc1aHrxai5hAvdtHyaKxxz3fDioludQCmfKbO4VvRpD5Bo/69jQF
zSB0/+7W0i+WXmVqxfhGNfWo2Ixf+gU8mwScIyRp2GwDlqgDFyDzn+WBphf3JIkm
r0SxcLmhEbVedJXsUYjcf18go28JEVxG6g29yCt1DkA481PoeLeevP96pV78yZZS
5nQbeIcCat+rymkMHWclMTJ06fhS56c0ysF8qYL+YFfLMJm23AaSK9WxxuaNHfgE
qW1l53dtK+LzMM18xVAfc6ALIunJjlfewiYWlReeJjgZg9ovAXFyvhUTuDdykIxS
0GMKR8Cfl+6BQYRnU88c1Qgvt3qRtfEZ3HGcV+FXeXs9+NTOVHktRyQMARqammDJ
WvNLQnlePzyjKldP15x6b5lOYznG4r+5I3CQ3DMHVOe/ew1lOwCCFO9oK5wbK2Q+
0oPs8vrlWm9q1IFfInkYOgyp2R728rJ8a444heKpVYqw8E0RrdH1ECoBkQdEtWyU
OMopS3kzm/tCMjibkPW6mg5cBGnQhoTeJ6TEr/nLY761terbaPd+PBL9RbSEi8vK
7To1TpozZL6RRzDnkC+xnqJNP/9JAr/MtPav91hQxwAuhAO7/HNYhJaYwH4SrvKR
/B8xTsxoMXdaKfp5VHQgRU9fe/NQxg0Wy7ZZRFcqfX4bt/rSRqE97+kGgw5iklPq
mZnilA4MQezJZHCHDR6NLitnNfakhkRD12Y+CgREyGtM4pXUgoXBoNSkPsF2SzOn
pFHR9ZbLZjYJtHsMV2eLBafrsyAsHzQfYtZSnoGRey0fbwCGG5gDqEsj52atdePF
GvqWplg6bjUKLGZaN/YVXKtf4a13zoeS+QIegF6IEEN8ga8oKP+tFtu2CrADT1ie
lBjWDxU1z8huiLK9lcs8M15w7FLntEI9TU8UDB2kY11V8FBlJEmJ4UFAyIZHLfPY
cYhuXgCBp1khVcNtuoSJbzI81XRUPqR1knCH9jKb5kCXKd8lZKPlsFXsjLFJ6BnZ
kGzIdJfDXXroscFAn+KuPIZMWS+4nFt3XO6oDTdauP52uf3lK1OCCDsuXlFiNc93
IFonWUic2dTjg1QwkEN8aeyewfIeFB9fQ1r9ecwJOuoi007GyGJWMDood3aDkm+P
vcqJtz39monaCvfWsBDnZ5GhBDqnD9xGek7v12EcBP+lfcUW2djxGDtUoLqTVAa3
42z3caf5o+cSvVw4OYt/eDmg6zUWcoEPMiMomsHUjrn+PTsh576FDsCcn0pLRzKo
q+c3QBy7poNnBLdnj7hjDZZCUr25Nu6CPrWTzGzQuJjrfIaWNtw9hLzt0npQIAi9
VaiAsZ0iadWXpSB6EO7WqM/0BAJMSKVmdHa9MT5YCkSrIMxQ40apdbrGOpeqxrC1
JZa1aODD0bZy5TkV1lWLN/NXo9l440CkGya0O1YcbSCaDX848KOHxyT+zmQzGOTr
EjYZ1mAZAfnrF/B+fDf5mwqNVDocPmobx2/pWELb9K6uodXtAI2tZP0g4hn3lUrU
ejyC71vsK3B1+k1E2KU1NqItQgXcXkW2WefEKOHAS57312xNkvGtOSsUMVre+tnJ
58EmQKEU8QFQl+3PfpmOGu1nfwMAiaXqalUsIYA9HqKXhc7R2DLGRJ9bDNCji7CT
fFuU9nTCybtDWJB7WBpxDGVx3bx99brLq+AI3aZ5KhRrkF6QDn7r1DCA7X8PD+0U
h2DzFN9qnqItWQkmF8xjMP9s+p8ON0QdPsSmLq72SvmYQ5UrNdXRcAsdlvoWUYgU
rv92Cet2CdJTNllE4W0X5PL6cqR48MCMhcRVvzW9FxJjoOjXkm3XSABko1dmVQ9/
Ry5XMex8hv2dUgCH8DNwUKUT+Q2rHNFOxCX8wgkZc6J5lw2bfZXjw6X3rGVQQtZe
h/KumsVimI4E1RNtmlGBgTVvgoJF9XyYUU3NDm/Hy+rOhlmmYnnsoEQrRuytct3x
ZZ8Yc4kfIQtkmN2frhqSQhSFalIqjIiZ7y68p6N6y+CI/iBdQuw9+oSOURwzfWaO
4eZn0FThs3rhdj0/IuFW+Aj3m3w9MzBsnEEFlQQr7342sYlwlFpfA0sCTsb778Oq
IuKCrgWedv472Hx1vFfDIxB4LxrNsuS+ctwgHAUvgHufebZducJ/xqVtkgmhn2bX
YOaiuW7nGSh5b9lOgEAI+9hTA6OyCRiMTcRBqtJt951DFCvaXzz6TCjA/drbsxEG
zHAlNUDzvIWMsaOnVFQ9P+S7e5dz9rUBMGAlkpVmoMBeUpXNHZF9l1FVIpnwBS/J
xbFD3tBPtRJmb6hOSb6kXriQMpI5QKM51PZ5Vw6EtA5/2P/GfLdFW1DB0CO3GoX5
g9yNqInEKYh6P3GxddBuhQE8jsR/OMF3OqEX4hkEpPXNLB9LBleDYAlanEHgNLru
j8NYrWXYI4WKVRzCdKpLd0yxoFG+XqY85BZ8y6tYPRyMqhLoSemvBcCvga4uLPSz
FoLIkU1/ciKrkKZo3R5vGvDd2cb/I7DDY6uSLbfj/KzHJEbAvc6vVQc3CeR3lq7C
j6gZRPmbhTR3uCpZNhgUotng3dVXJ/7B1g2aditsdDIPvPkc029Gy8IiGT7ZV2ZJ
ftzYpFTt+pNqLOGjRgQ7AnTsXFjf+yy6WsDOy1Hidj8tTxCcQTW/6l7AHhP3Ubhv
NtYKkepncyuiZ9AOx/bOrr9QZwBLozjaDGwl20pBUvuK1LmWHhRg1WsHWSpxdzE8
5c4T247RGAmdI/XBh4WX5h5Q/VZoOAczazkQ/3BjVA74s6M8Uj8UA4OZNNJTkBIt
7Rnm2eMmSaa4D7jBx7WTacb/OTuL/DXOvMU6C97OyoB4fIynK0BO3SjZysYqYyZ7
uBJKcZkj7zViS/YCQEOoF6rafpDG0k43bJqtHP4CYQOlE6XIvEKiXgh9DDalmpxj
yshixWEBWsy57Um3PLsMqCOHerFKnhsRmEy4l9NLvWnSepVE+IluIZFdh5zdwKHx
OpV4mCPs8IFVcDhYJsiE39cfmGffUFcRgrq5+5ldI4FbSXy7BPlkMthc1txqVloF
gmtvifft1A1PaJV2UhSYQZSeGNduH7f/bWa20q4LrkCSEju7FU+El4MEYt6/n9Eg
OMBPyQtKAl0VEANt/eAcMZXsSRWlvJ/HxZ6bKc23LTLfRa0Xue3AWsbKcstb4xgN
JVPNarK0GSnIUixJOqjCQDCqdAVCjo0bQDYrifngnFEiPKMIAC+LzBgim6Z7a8dW
dKcErYCS49npMR71i4khGAkqU2Lz9lvknPmxT5nYZGBPXYS8Npzq68GLtOrCQN2d
8/mbNQnur0eTM4icaUEIFWofsEHPLWF1IgWgisgTk3YCIdZwOMkDKysNGsHL1J0o
gXbtZf8oRX4p40+X2myz+pt2XTcywBrjPTIG1U5YCnsBdbvml0hx8TlOvW7wxjMb
l5tEPmzidbGexCq7DNLs+cr8AebNgk6bcYmSCfAsDFnZ699Q1ecJ3CPul325OH3I
bAbDuzdwqmV72Fm5oCYfFPWIemVbe8EyczxAYUl+lDHNx0nKBKwGSOBZoNv0Y/bn
IPeXmpIN0hrknMudt6opc/zTx0+2ksYkPKtt44X3IAPaDxhaaaryWk32yf1wdnSQ
Y5woRy9r6s8vzqhUug+taleReuSRrqY5Z4spU+tdyT8ewADuKSEiJxJ/4QVgsMXL
B+xOkuLDhi1+kFBIjxYd7ORh2kn93lnX+uITwjuctlfga/uxFYwkhqoAfiQroTjQ
7Paa1oJ/VeFHNcPTxOBpWxCk5PaUbBUCDBO0bLSY10+dvlKygDEg/eoCviTO0kgp
TXQoAvYZcjg1wxRc+nyxq56BVSaGu24biT/DsGwtwM7ClWoSjdQZf29u0uZPBbP7
Y5bojF9IO647XyrqBlvV3Jf1MwKPLKokxBZGqpT4sCPGIE5ZqFwVz9TTiNw4avN/
MCTS1udELXUlVAcrJF8KIERCcUYXhpfQJ0tn0KC80BI89PDwYwPpzWHME9298A9d
NMxWTkJm2myFu0PvnPwT/wwa4kUuNRQzJtQVw1we2W6mtiLi9jwoABRIw5ARDCom
epJRUiRyC/eHPGbRPJ+mnq/Me2f8sIzcGiHETJ2kc+kIR5XkfcfH+iuFkzO4DJhN
ZLGuW3SonUYbpXt6JW7okRy6fH4fkN1V46gEkuqyVSarUcoS5ts8PzAUZE00H2C5
jRT8ZxaQaOy4RjH9hLVS04kd5yiqPcPhvp0ccFk7SZyGnOn5XMpfgXOaqgQ9aPgn
OKXdOXTxGJDdS9R8iiwsulJcx3mKw3hcmg2w8Ja+x4Dc8Vyv0IpxXZjWNG3tD/Yg
RrLZFWlrRYFYJ581SVZ6ypJDnnlr8xBwc94+sFmzzuMyXG8CFaUR3FIinIJ3jrnC
NyurXY6mJrIJORvtVK56qylQtm+U3aiI4DQStOAkOEESHJzW4uux+Leg7g3Wt2vN
lq9NinbXc4QxIujxbDLfMMrLLsc45ZTz0jHW9h8qF/wB1EhYwlej0Y9BSmSJvwiQ
otsHqq8WxphXKbCVTFxqt1Kh0ws7O0DO9t94Wn4RgxaZNMCCPFW0K8lNJd4zjbaL
b5RQwFguezRHmTiqpJn6agxU4IFhb+5iez2xbl52VxHVrBy/9K6RTyd/LIQmyJ/I
DKDsYlUv6m/4P34K6Eq+3nBBetqCBV/KGaDf9H3KWD4y52Xj4c3nvzj+frXtuMqf
DamqQnaW5fyQ+0r6f+ANptz+w/hOV2FuKJWehY1AWLm6VMqsgZ5FfjbPaOiBMmfT
C8wV1EasgFGU7KMxyUWIsReO57Tq2VrdJxzLr27iLVospOzhQaTjheBu/M/ncWVC
ZVMUNoOuW8o6/rkXEK87CT1pP8gseUmnGqC2kFJRX0wx6uLMapa2ujpzF0MZFjQW
RAaP6caTkn0HkusvQjxH/Ll+ztkBkqXorubIw+T/QhiNv7hqNJlJ0ZhH6Rb2Ht+J
2CVfQtnIu0+gy/tCaGXo5YfY2pL+vg0+Z8cERJZTD7mCItxJdeAR/N+sBKkXhHWN
hK8B6ogHwLthhlnP2PKDy1ygvOqTemBeh+WPxuCxT4H9Lz44rIJtD7hdg6h/xDcb
H57AbjQJI4YnvymXn6nErcIWscd0WPa4zKG8N+7o4HAY76S35rrN33hAYWE2/g+A
rOrRAcK4Pqj5ui/1G1SHe/JY87UUwR+3atx5a9CLay7p1ZN6jpoK/POhZjjF9e5Q
4yMqk0KNqNsT0zuXuO4VeVeJC/J0r3Kv5AYBtull9yBzLGmRrk9ptFqKDx+M/hWU
MbMN/cH3IZVOoa6fLklHP3y70Rmr32vQwkkhL7NU/roY2qnWHnvJgdnZbKe8kllg
k9FWlJfhKbCNgVPdrX9Q+Gu7Vr3hMnDcbvu7QWYMjkHTEN+NiuE/yHzDd8jf1EyT
oovnIZJDfK55TR/h/J78XWkBmdARQUb+U/2nVP67tOxDK5pFbL9YaWVji9RYZ5rC
viWKaQVyy/GPdodxk8sSVBZmtnx5wDwA+l6CpuV8l4K2iIDbYa5T9tPgsgCcoY7W
KwI1Z03F+N87/di/9brtKPvKaHDrK0fg7S6woSfYOrSqNP+dienYLWyL+lVrsx1e
B6AA6NTMuAW0J+eN6h7zf3RhS2fBgooyzO/uSmBL3E+RlUttys3pHN70nfSTibR1
IIDarGLApDbcvlvpQ97459wpFq4AdCsQdNVojxgrXI9wBPIFEjoTi0eSp7ciAZCv
wDe71eMsPNTnj5gFkRaFY1/2pvWAW1WxngqgGRl4iH0OKx/abT/0IZC/gdq6UMga
n4+FT9tPeBSK2fH4sVpgpNT6MFb5UCm+5GH3Yd2Fw28FVpMArEc0QY9ECLXB6G0L
PYBw/D15R5l/uFSDvJrO4Bz5JCvpo8AKaNUHCopuwl9o9aOQ0INqW83W4dpb4OfU
i/cgZ3U6NNvt4Qmb3mcKUJyK9dfC4AjDBveNmARqmZ4M27mVPhEO3aLffNmlgou6
sCUbrxl6OSCX+hME6VWkbOGKT6J+Kz4l7fPV0qKvUkVMvc4mwIHSOywk3E+eOe4d
W4AM6sZW4x1MCuPSRPg51sc4asoiG5/pn2btH2g/ehqHpSnzFFdWcte9Fd7CPCTW
PCxpu5JN5PWh/ZB3kK+h8eQugJRjpoYneB5owW8Mgt+NqpZ8MvTpc+evdQHsbwMN
lsw166NIdkvxNF+hRKQliPRMKdqjCH2/MZTuMMQ/UlJG6alFd70wq2PnplKwXJYt
EIV6Yk3z7atl0SYMdlwhMMKfMprIt4fUlkq8OrFay1mNBilNEAMkwVA/vdGuH/LC
UcFi9jH7M7nY/xgaHPYpvxPZqofae0vB8Yr6BecEGCX68z0nLXTEIF4rQHxZpy1O
KI4jExe7DAeRsjXgnv7W3yeKaHqDEfV3U2chreOasrUOngeB0PoTFsyVDk+WWPys
AXGsCX+pbXA1guKOsUu7Yj5BES7B+UIumN42DjRAJ2il9WtGpiwWMdWhJxcZo9jX
7YBiCXyO6130jD4Db2+kLViRueICJTkDZAcH09Mx4STZw8J/N3r/kTMqJjbqOUb4
MyJ0IbCs7ZHUZEJbyihA2SQZZxzUx8Bz9U1p6+O9oSuBlG5GoensT06S1RowEA8Y
GgWu2+uM1KiVNwVv9tfeoiiXSHiJkpcjYau3cHL0rJKXooabWyEc2qWbS1rBOshd
Jog20Sic9lHQvasHo8HlkDJk9iol0z6Au4YbmlfROUcORIsLzvNsg/wEQBUMXXlU
N20mJSLTWNLcnWNr40Q+Tgcavl7+sXFGTV5H7h45OeaNyuZ+KpDx7c/E60vh7jj3
LumhTsY1G0MSCL2aEJvfLuYQoFWZ6Sfz9yL1uSCT/EnMtYnwaT1ra61XpxM7oMp7
3drfeQjAJJ1mEDFAQKbGtlt/dbnouCBX88DzVdKO93V/0ecqhu+hf88+DWZ894u1
6rZeYvkTx26akBhSJU9jfQ91R07GNhYaF/qYRre2Xa/vBpDHVx2W0d3gCVdYfLwA
E4G3wgzMh89r0TxVmBuy1snYf26QdSEgsfVUyWhCnMxqukdNzMuSK0YdwQHpOvB/
aXuMl7hY1+bkUYcSy/SnINoHk+AxOg4XCM0pIz0/1dlOQbxO/9ZgIyleXZJaghIh
e+/vNg9B7AmvU+qJm9n6h10ary0OBMhY2807kvGeFIboR67s88GCgybI2VZ2KesX
qsC5FVnh2FmpfdJtx1I35oJgAt6DwN/j6sIQzV4U0OffE6OsFlpgewWS+uKWUffi
0bQN15m+/M/Neq2E8SrV0QTEz9nYXoE/zoSmE/UZ+QetuuxSuQMSTBnShxvXbngM
HpsFLQvA8frJ2MwMJsnnsgygiS8dZiddrMnjYkcknIddmyJJJJ5beA48bIF5IHI7
XraRC9HoCCPOGtiZHDELaLzNTJBwqfqyDAY+rf8EOS/VmJSc3oEFJjVv6CcTDThq
xUfjDoDAtiMIg51cEr+WXH/DpE7ee1X0KWVYDddbrVRkGekVL8u93ROVqLZmXN1K
wHR/p/DznmDf92UhBwQyL4TQTtnvz16HZL8OkZZBJBDde+1/m4GEntYqZg4LqguB
yXoXviMFN72jKhmOKGTKy+pbyhUI1s/bLEtg4S6NnRm2wD0kFzPm18XmZvrc+QKw
aRKrCCLnYmGeShv5meRGghuCa2GGFR4cq4/YvvTJhElQk964CCY312pd8b+AZUOz
hUacdXPRqHfV/dN5cGpkpceCIBxorfNUVkcStaEL15Z66w93fSbm3hP6VbCVPaTI
ckXzEibE2lbFaGIEpvJ105TaW4PX3vhIUAre1SZgGctbknjwOCNebO2qLJ6H4tuU
zO2CsVU/1DxaPzadCCg5fSMeFVelFxWZ3m4nSmFJCS1L7Ih/3zR15Rv2R4p9tqgS
u6GUS0cmxThZaUI0eHvfPQ49gj5PioZOPtGlIRXyp2ck2QxvVgcTOt1XBl0IxmAm
3S/9QGiU28CD5NJPUPElOep5whGhRBvM8ffxCCbiAyChDCrDUnUGPDguwj9ZvoCl
PY5AJJdbDCttdSmiZQOXVtLEfyrCPdfy/hGUNGqSsPU0si0kOS3Ro/icaH5PDJ5S
LjVCWpXA9Ep5uxD3ototUNMYeGM3zMKMf09gzQYyugUI4mQQ97HRpiHOqOrsOsgD
4LiH6m4pv/Iad2GOaY5H/M+kF27fUkjetiGBgOdXfAkmeRa+Ki480m0hFqVA/WZs
L9eoiOCKTi35tXD6QA4CWtK0FsG3SlTqScaWIkR5ioXWbmmgHI3K5RaWytNG4FFe
lfQ5ZDe8ZTe7PDescsxbTLJ6FPS/4JzciBIajq/FTW+ofKHaBkkCmnIXTipQrN2O
se6U7Q++5VQmVe3xqIQF0LgQHQpcPLgTcxWVtkJri0qV41hGQjri+KnLsKsl+7Bd
cO/0Ba/3C1lMV0b5ArC9bHdo+3Cb1o9jmKcJxGYoBnekZCLQIIgwT6MIJhrj0N9x
kMsfjtgQ11d4LflIaTzpY8HV5kA596zCebCHfIYK5msGtedPhOzuhbhnE43c6fC4
bid4aNvl79sGwl9Q56f395B7TFrDX2XYg3WgJCK1FrMgprOKaPdtgButEzy4vEhZ
7p77Cv3TkCR70UxpKiMGkBqrxhirkytFzc57AVMwcbzYHYQC/aW8vK7DQQHPqEOe
ZGCdizDCc3J06WNbzSyKjH7Q/KAducK/3BXYAHJVzNXy79ZI9BraewkoiQGZjY1i
CXFmTP5JW9nivpuEYZSOIxv0gZgg6nJFQvy15AnZl7JQ52rMKAKnES6XyQBJ0EA7
JoWomnJ3LcXcnBS2OiEO9GfAvwI8AZV8lcu3J5TmO4Hp1laLcuGobdv53PjeZCf7
vggcKtyy4Jz++Wz75uCGb3AyCyW6YNnF+Zauw1xaTNbdRh4/ayFaE1VwgFrkTwAL
SnX3YIzfqmLI612e7lvd15dovrMN6ncxRqn6ioZWSnxiOwXWEOVuVR4U51Cghc9A
jL+eg95zyDGIoPAIyL+eRGGgfrcPGvwO1j2nGBsyqQ30oX8IoW1ywQOtZwNT3unb
Ke0A/VMQwL5ZboooEBnWjM3cNY+xO0v9mf3wbaZdxU9A6kJXwyb4SyvAPM4qGv8M
D9mj0Q1u4ekLvun+7SngbMd4dpWDVSeVrcIEaECR1acA4KLQlQi2TVsr9S+vg5HS
khGH7U1hf7upmqxdmhpXbEtHEL1OJP/1wR1e7aRC8PGvQsTx886hgQGGc0aGviHO
Y3fX1TS5ChkVBtgv9lhzVqQY5HjDjU8+mlWlxv8uxViNGtZBcF1+2oWz2O7MHePh
JwS+2D3DKQ+pnclaDiH2ZFtZaVXLVRqC7Vjahk7CVtodMTBCWwlB5VqNCpmYhrkU
iOofgN/wE4TNloeedKwCOHQMDjwT69+nhuO5JdnpApH162rpv4dbH/u6phOfc/FX
DtKKkXOQRIkoHSdQl9JjX9tCrNn83Ui6Tj8kzB7kdjSF+RXm+4gPo4aLQywpX0Uw
HngbczODft9SdqMjmlZHTvhkMFyvW9xrZKRrH5N7AO/Ee45W/csd6dxa5xzUSKse
7ptzecuq5fGcOBxpbN3Eu+xLqW66PMzBLJnyGN3+gdLhdlMTkH6TOltSrTLjnLuF
DRyZ+CoxStzGWxJ7COasvgolqD+cx9QDeC8fW/qKq+VqnGnwn+6VUwWQ21EQmwLg
PnraxK5+KW2zAS4oMfPvPJ3/aWpxg1Q/DYS+wlzJWvZ112zg+DK+2Z9f3Iwv7iWf
EOIXXX5BtbEMKRbXchd90Bb2gVUeG+SzzuEOMUhKL2RV25+y4nwfdAFxNcaDpKqj
ErcVNS2TXK9Ba5Ihsy0Z0mcaKDcRNFsKXvUCNzAf79yguyjJ7b+6wVNCdV9+biEM
EbzHLhsS5xQ2oKvJunNTPTjS1ceup0XxXu8IAOdpkPMwkRg9ytn/Sek7C9FP9BNU
KrlBzeLq6dG0E87mvMB2h6DB08S5NFAEVXDYWEaSGS2/gFmKfGTUdLNBj0REY0Ta
AVUOIuGviVJOR6fuo/SAOiV+k0yrtLQgRLA2JhUBEz9w3YVEHWKMK5kuFjqfUUGO
SIqmBFMI/Cb7nNZTnElNhvEyUYUcIQMnUVSXOXnVuGQHVaHq/GhGW9/cg4I/Og/Z
4YumzVCWdmQ9KAOg+36SpWqyD3wtqk95XqfgILJwTqjPxHGE4x6Vf0LXn5Jl+TXY
HrmobOUSMyW6UIDvp5sGicsgwCgVoXA5txXg+N7C1J923MDrapCLFWVcktiFYSHg
CCWBjSH56JtPgmH9ZOM05TFmOfum/KtvIJfecodjFZxHsU+Ff6pzocLhglV0sxdp
tDXqjkQplwwklU6KblyBFhXYa0SnDg9mtRikcovSLn7Qc6Ibdd6lJWkW+5mLr3bQ
GVrOJwMNDJkt4ufMEBe0Hym9lzmnNCHwe6l6zAn3YRrIN3YyE3mThfL3G1DJ2FGy
ebzQ6LFnNaZyZ6XgeuMcslmrF5cO3rvdgtlZBPqb2+c3DX2HlNZijlxTuIHbeUfu
QnDlTr8Fd72G2fzy72LHd6Ff59E/QBhSuqJiWsab5u0EuaEhFLVO3X6eQ4YDhmhr
HsMV62Rfp8pLySp/Dkz9flBWI37f4tzT8sUwnGrZj5jqMu8WFaUCM//XGw4tzDzI
lp15X0pZ818GD6bSBCVusQInNf3mRkt2EfsYk2+CvJ8w0bIm5ul4Ca9AluL/FqZm
YHTsz4G7kMXkretHO9kyax+vCbVkyolb7WyANPcKy9V/RgBMHbkodTO/S511I2Wk
5C9XCoAD0Lo7qQd1qpcZjEDUl5+Joutg4AJv+8jHuOehXkuYHel6D6XQ79p9OG/U
i9prvwCkj6jBySqtw5jKTaXFhGVx64zOb121KjQdPFuBkJRopppFNTbqBkd4aQXL
4hoC1T2vW2PfOXb+dWG9GK1VWCm3y8lrHz9LG5qOaJ6z5hwnsOmAUUqYtZ26T8WF
UWlUgDUGmRrUhgwcVPIyI68C9EqCFZkUPd4XcQ6EAmV8fLBSubZxpVH5S+6p8Kth
KJQtBxfPtZWumsjppPasu+T1D8xTSxAZKBiZdukiqAuZO+hx6mj9sDgRS6r46xHR
yPWEZ7JS1ChtgexfO5o5jLpMo5bjsovtizF8MqrcYzPlcK9rq3boa07UWRCycBxF
4TdqddXOhzsrVEX0ZPzU4x1v4UoNJ0KxWggEEzwluNln03lUVLw+Kpyo0UHPFLPN
zv4tDkFMIuR/7EC2dLGdV9ou2GC2jmf6CNNKBWFW7k4c4uSm/0+OtgxBu1ramOa9
+G0Vf86UKBA9Sjy4qgvc8WV3qwHe/XovZuoBk0Cbvr3nNp1f3x7O486RwB09lVCH
wCV2RareZF6+L4yQ/jjtbrV3RqvjqaQzyIvkJiWyS306taHxEsDAtEVOSsKermQY
hhgWXFkEz4GM+1bYwl99oU/lDr1MUZdAPTsdtO2dCvm1lCY6baFw5I80u9fLePJ4
XUsA567ucVmfrgSRvG6yIsMuriPvVjfBgzN/Qe6EI8n+c/UpDoYtNcUPqOb4FpGV
3ddJ0Ebksq7FX31bKBShyQVhM8Mb4GM8QvaAbSFdjfAlNp31In1s6P8h2RSuGGy4
2aTyDd7aUYMUeyLYWpv3DRdROFTICRFN36nS4lwpew2zAcq7i+tS4lPplS458yGx
Wo9FU3y4azWejsJ+xgUQ86bSu7XJWu0hpixRpPVCLP4UVUjQtNwuC1ibfeZ1ILHZ
VutX55BT0efVIfKoki69c7LRAhcqMAn8/zbV9teZWb7C8vn7mUQhXoyCTgmytzEw
PATFWE8JM8Qp/punL5Sstkp2QcSeMPkMVBj877hFZHf4e3k8AHKbrfU9GKe2vuCV
/WgILebbE77fvWDJ55RRx6hCnmvN4lcq9O7TuRecePXBcGw7zVVvXHyP0OoKQbPl
7sKRajcgLlICrUeWLG0I7+22YgUO2ckYN52qM4licFiAOREHB2ToOsv/QwdbDRQt
1A/6xJguWgshe0R+Vsq7AIHo1P5o3APLxN+mdRxR9mfPwv/ppiTTHPd164cQbG2c
S+6VcNxporE/0ultnLLZFBIely7ychDQtETG4k4GN40Yd2NtnI++U+OzzfwoTLO0
gkBmXZ1GJKg7vBTNTSRqWj1R2peTutrSrcuCDOZgAWE81q3GQZxeDaWA4ofk7yv6
bnkw+H0Lj/Si7iqJEfMPEF4XF4F2TbniNm7jqbeezXz64wF8Va+SciENkSu8w6R1
Wa2TVusmdPFgbenW9qFU9yy0wJmBFacqqVM3lSXbu/qdW7RsEEY5vuWo9CsReYio
q+8l3BxdN36mIOK1ABXAKjqA38X7ItosHDzQgeUgy2BE4w9plm5oWbFG+56oHmsz
2fYmdNgtvTs/zuCxphQN0Zl5VRzPC3hyFQ2qfNRndVaP8dGNMMBXMGA/ts98uXlI
x1mvNm0RGHVZQnRhBHnRC7r1qooyQrtwYHK/RyF/gYWWrfnnig8dc6VNCoIvwhJG
8RSkEKkhnb9bVZMjGrMvvqfy47tpdaMAfx6uEUSnszoJMiGWcc5N3BqO9YSR+uON
SKPcfR2HXN4+SWjlyQ+TyGi1l8+K3dUplsPIf1O3An8WPY1BMDLjV6gikW7vdm/s
BVfGvnz7KVsgRb/XXc/2BgSHxxANEuR+hGIlMMtZpMMSBXEpVhB0Lzgnht5kwuEA
HJLl+qFlG52MlVveNIdNfqCWAF0LmHZxUchlOdx4gzQX8JFsQ6uYXra5hOdfUF2J
OJodyr3SyYS0J9M8dN/zHitY9VvvGDnjvidky9kTUuv1YTXzWwqC/bqZXxzc2xr4
r+u3wt+CY/CzcWxDEjDh92wBn0quw/Eo5oWnDczCeIzQbwHUwJxQnIN3s2TA32I8
l4xp5cp9dGupdQVGUEQo0Y9Z7G6TtOzY+1kXdM2dDI9idQ5zJeTsG4NoNIWZ3wJM
9Mc5Dssdc75GFJJVXsr1gBjsfv0Dl0pVhwnqufA4VtvQ0oXVr1Id7WBXiKj7/1Wm
X/l5HDFoDLGHjd/0+XP01Lhw7+tsUVKFc9OXFATW+Uk97iu0407XaBARc3PEYurs
/axy+APE36YLcH2ALa2rB1KlLJmRChV0vSfqE1qUhYbmzusZ1C4WOV6N8TV0reF4
pOlR+0VQZsgjDkckCQVQeASZP5WMsCNe19hX5FmiBiceNa8mTWt8WUFh7fLaoip5
u+NOk0uZK5tzM2csZkHErKPQACNtJL2kfMM16HazEcZM2psnmFJl+3r42xBFIT2V
QeKHex1eOGIqVi+Gtkt8mN0k2FzVU3fD6iQK6LxnMpYdP14kWK8YkotyX2EUwstp
firUSGYGsXQCS+dvAR4ZG49c2YyPMcrZeHyKUWAfZkuVOqSHt6duaNNqAiIeqU6s
3jyum80GsEm6oHsq4ogKfboC6tz+OQnEOKw+heWAj8ipcXu3LmIjZf3wj6hDAmVm
0W/4nnwPQAJOkrHlkEeF49BeD61FskkJSblWYCZHzeOcWU+Yf2xw39qWwnEnq/aR
9wPukxYpe6ZyY/9Mlm7z7n317K7t7+g7bGgpOGRX5w4kJom5nmkcY3qQRAxOwVoV
QJM3E16b9Yd5a0b7sk1sXHV4bR4Gyvvbdt53fXvsBX/w7bsk/au3vCOcE//2j5J5
3UO1ltA82gLZr1kcn/YCZMq6rT6SG3ne6FwmPLnYuSbgSdZx/Vz589Opu87UIFYq
+Ei+SgVZ0UbB4BIbe+6uEokwPyF5ZNHEjVUKLj5S0npHSM8p+E59+BBkD8blE+H5
v4+QCT7zGfpFJE4XdKoFLdr//KF+6xcJIQjxGIy9ShjdPYHfn0sofPNtBJGgPzIx
UkCWoNk5sPDENo+2jW+rT0VyoHq6NtMfWUtdsZcBuV7LS+/wZZaKj+nTJ16+AIC7
tAVhOKf8sX0VjqF7w2AWIQnHkTnSU55BNw0rSAQMxec7dQEdWFECuZnXaYG/zz0l
QBZjn2PpVcjXcl59a36T9x5Xh0RLQWlCZM+TooRyJsdNTjAh1VLC5zoEXej0ZGt8
UeOxdXZjixJPNgNsSNFSoMyEeNIz8JvP3ogQjlWVDwQNxaDDJh9WBVT4nxzcOCs7
F8Zx99ayXQVkW+hQeI2YPU2So1NYuFfS0GYJoSqE/x640ZCOofucLglG8GiZxWQF
DJOAWEXvoqbB90Hw3xONUJzbfDR5aTyh/HVEUJXhOlzxntSoWidtfJXrMFXauX2X
ABiUiB7wZQBz0yi8J2/HdtzL/vsNJ3kwGCXrwmVru7rVAlwkEXBGwboO2oxeQEqu
hTnCfJoUrUbM7dbcK6g6fc8yugd3Nl0SwOUBFch6cYbHo2EylZPRD3t2yOSpQ+Ag
36hWDYhZTWNTJClNaluIMyVfcAzEH6yiM0gYTMNhrWkJ6I3Wd5PoQIm6hvbXDdMi
bwxdRYKTo9OO1vWMBHA/+zxHVxE6uiJF6+Ac8MNTG9x4DjOjQGNcVoHsUNx9VUJo
BkbZHtAajsTF0mYrNT/ms52WS/JXbIapFh9r/5I7lZDOg867SdPeVGuFh4p+FnzM
xyPfLxhpP037jzxfLldBVuHbRmfX/R7+wKRNkcchza0+3UCOMqjhxxxbvsS7S51H
tK0vd/QkkzlXVADi+JhSW6/TXjwXiHRfaYogZpka1ftcfHBiaFgVmN95qomzseCo
O/kekKjgieI8jT403yqECFL/Sczg0D0gQ/4l/k7v6ADwrYTk+9Z50CD2YGBmBxGw
tDDqMwNDS/jBoHdGSz6t1QNzoVgykPeEYW9hhnnhCWQvxtQeExZjl4uIAatUwpah
uugfTQQpVDJSSTuDju3WE20sGJjnQY74CWPFv+3ntvHk2w9MWl/EmY3upKAT76bi
0Z6U2n7AASgth6rUaLAxZp8onMM7V5Ghu43ziL1mY/mnJWhJFO8ZyjDBBPN90BGH
OAs7IKtLZk89n7bMGOp9U7F9HmHK4QlFhKVu6z4i6c3Ob9e65yHOWRRaaGQrClak
AQMdsV/njQkLj1P0WZlys+VfgkU/MXgIKKu2elLmo8vfS6bQkqhfDhp8cJiWXBox
TQYihAn5PUKNReeo+7Tu7gyUXHoctXnZHN4tKaCMFCAOBFt31gvjREkLTzxnuGp+
W0QzX0hyLKxpYEj+hkOYqDnNsQD6NhnGEqOUjh9QxwQ0d9nyZpfT1SPZ0RboXz36
xg5/nOijmhd5I55f9J1MS/8+PROG5xcQ6noFdOqqmhSInbjPXfOxLRRvTNAdBm69
nLzmUqSMkfQ9v2lsuW9qcQtBFwP3fDBLOS3/ZMtWvHE5biA092r0Hi4+Hw0VnVQA
RIW1ucLgLIr5SPaI3JsvW3j1b87NXuJBOsH3JjMt9fms+EJz79gdVHfrDehhd67m
XGfw6Gwg8B+sawAbissqcDCJI7eVrn2NOJJfITAhahbNdMKrG+Ju1MuYil3M6IPH
uVRyABX6Ma0kYJPAmB4yJfiJ1ryc0ynziqHHKtwXib/Gwiu3kGjLUw/tUoHfJ3Lv
cL3TRw+pz2UTBFvSHQrau5y8oMXvxWyp2K56Mw0X21PSTywyn9os9+fHAFrqI/3B
XTsIPz7nM+q62k4kDZ+QjqiPTZ3gdmjRrNgGjf2q/E7GoEbaIBG4/IuyFDr9odQx
PXUkJ798s5qUBUK52VUkBpYa455i6AJ/RjcYj6fmPYy9qGIusR0rCK8PQ1udwYHT
z7USpJftXPw7I+cBz5KS8ZwIBLed3c40PlzkasxXrtbUobPhkHuYiVeTmT1dH9mA
7yFY2vlnY7QmVMOzGzIq5frApkpc2TNvzHhWBPxxucJ1xffSdRWtu6jOOnvEVPWl
Jyn/tw9MG/y4+gZoi9td6S/pMogM9JUek7AKidPDYNWAK3wsDBdJ6epDqlpwHf3q
P1eaJskNB4f7AgKfCGvXiYRSe5+9cpQ/Kw0iXHIP9IcEngeSSgnSWWxKQECoqV5j
g4K8ccZblR0lp9Wu6IQMjOaIOCGoDhnUQKZfVCNjnCdhH6Q9kqimUt+JPvsGEGol
BIycNyoCLhxiyqDrw9ge2KrZPxYmCCWxznm+Ik9+SsaPn5wmrvyCmDKS9dEGpSSj
S4wIpB1pBHSqTYBYHKUktQ8NyMeGwTgVn91kxkKDCbnUDGbU7CWtZRnfbUgPSz+g
VTLL68cgv7Mx+F1RDnCj7OaAsQ4ZjFGSV8YPEdh3isM4HGww4fMWTIoczlVhgyLH
tLRDbcblOrH1uQrn3oS4HNjg4QsSfHg+jyhlY1Rn2SinkdxRaCUoOw436c2xiwQO
OhKxD3lDIsr9L1sp/YxDb9YPlUtBiwDIv43d97dYHan7rnT44AKqsorgw+draUwT
V/qIpYto7iIw6s8A977a97Ug1N/cnzqF0a5zP5W3KphBZCA9PzIBiQhcA0EALfVM
BVRdDzLvR5TLhmfrDWTgS8Ysu+jgHfGd/15H2JWN7drWtwiVModYF4ZizvFN86nX
uDfgBpWsxNXh+GNgyEVhbMOgH+sTEb0Op+Tv9IzsQpR+YkuoIOLEEw1kSzPtZfA8
WGvrHyPjl8LRsjSeFhXbRyihygZmQAKVIvmsZY4BnBcfvpFCq1H4tWy1EPImCCAG
9LnN5SikK+LPF3bF+E6EIn22xZacrn/8dHkr4FM1fzt5Q14kJiAv1b3ijo+77ud7
VRUMCA5wh0uJEchh+Gho6kTU+5h6ICy175PCzHOoFelYVYLA35EKvLqXbQ/sAC5y
8PMt17FG11Ppdaz7zOu4hjx0v+4qpndKbQaSbbG1BiA57I/9lY9SZ2YkB6El3jLC
mkojGlM1ye1uALC+Pwagnw4Yth9BDd4FJuF6N0xGal9RWSzGcZzsblt1c3ozwJqb
gtbk0Yh3GbffB06GKh7uO5Y8fgfhs8mdYN0avkN39diEMcj7g1HzYA6YrerA8HMa
6X3voFVVbf4oylTRQ/4TouSgE9QBtglwOeLwbrAnKta4UybyzJCAcinx+WPRuCJL
26hjsefLNb4GKbxM0TdkrTOeMnB9eM+D+8nhk8NcclLFeIQv9NaAtbJgK/ZQ7WYG
LzwHVTBZUeC5X91dbtWpzIpX23e27SBOCiVUSSjC1to0SuWgPJcQQTIUhgoMaZWc
sYMLc0/n8TOUnS2yGLpaZwM5rA5lMdZE8Ai080HfjGb+3MzGmylmz3D/8q+taYbu
QMuzFdvgCPL55hueQHQQOBYvoGw7XXj/jkrbjS2Ww8zwmXZSxmN56tq48pMd9Wgu
psgnrkFz8Av8xL/aMvqx/jFi8ddsbndlfYWQs2BGDNOkiso5+4jgh90MXoCcqqa4
acOoCEuMxNgi5TpcljjVwB58hC71jEJyetqevHLoRACdt4q1jeP2Ne3eGaq162Ec
4ES1yJhtyG/VgmioX8gkzW5OMLdiX258qJqVBFS/drMKgcbjCibZslrASaEwQuVB
DA4JEQzTok7DEMDi9Qb9ux7bhrP2U07pPIw25wth1pv//12jLwJyTqERK4kSv9sg
atCh3yOfK3QnsxaSnhYdEpX5sXR6TfYL0VVGnoYLO0hyUrt5yFQzQ7Dw060Bh3nf
2T5HAGtz9zEV3GTC413blUzYe8XfAKrVFK10vR0tMnxTw5K6mbnOdhbqrKAF5olE
T+rvV8GzMlIuK3wtk+l0KM1md/blgoGqRwOJdj6N9HRif2auZRvZH7Cn1UyWnVcz
HN3etphvqwZ+gmYDp0ceC9BOE0XfAOZET5XJsye2W9y8Rn4EUleeakocsT6BaWDo
/f5YLVKr+PRsxKXUDlpbUeOyj7B25onECQe04aMjyAe/1DMTTLGW3XYZZx0uiTJb
ePh0GMT9FIEanBTb5kt1pDV+EYiMk/M51r4aidxthR3jJCBN1b1pvYbj9a/X+5nP
RF//MQ8s22EOAJv2/ZGQPS/srl2QMYZUb2WTPR2qlHePGJdJY57tW6jg5p/5qFM0
x2PSCav+fKWBXPVLDzqEkXdscDK5Ak1X4l3ns5T3LbdseeDGP0YxpXJU52rTqDlf
SvbtSFNuuxnovke7NyhGE21RDcxuvlKO+Ok6KdfQ1Ntv0D7N+Ov0nHHXQYEZ/eaK
WgSwHw61B9hgTyn/wjrhykOMNyAcwhOS9y8XQKXXPzUATrWwtqMEzrwyXPSpgPaE
zRaFbOku3C2mWatUOH1PJB//jU/WrnEjC3/+36HguC/A4FcsHgH1Q5yDkWBYeqh7
VP4ytsCW1d9VSZPWuGxHqzHpnayrBgQdfsG4kUYkVDBHLtIInmF87bLO7uUQrqeW
ar/MApNHngzRsFkLOzKru2mFajrvopflMnnSWfUQqlVnY7mI8Lz9+GXKFg0xCii7
5ww9Ak0IaWOpBTAHXyu3AaIxOrIAGdhe8EU6ni4Dj+gVjDfodsOEfGmeUQG/kb6J
csgAKKdPDRLWPwRMK7vApBX0Ec8H0DTwyAzqDzVVEoUnFk+lUmur6XjxS4klbRLY
+QDDdBC/RQ46DKysXV7cwwjVUQrhgX62QaTnt6a5peo9hlIhTAoFwgQ4KYbEk+mi
E40DHg00vCIh3ZjioXyv3z3fUccyiCo8o3/3Dl+8PED+ao6UsuHwXy/uTjf6WBvP
JX1+NHtdX0/g8FzxJhZ5j02axhgQvlMG0p/QXYL13nl7e3VJnU0fnf/9VB2CP+E6
42ghtmcAboo8+0NYWoPJE2YqyYg15eRmJE8qzwBMLA7/ZqFoHrNTp3nYWOuGM02b
Oy/Qx0XkV2nVEj6aKuMe6+WG30NochX9mLVHoAeXnSyEgVOmJANeNJIgyg5L21TE
+w9PQKq1eIfCfYsbBOzM+UO8SYb3QGi7K1mZq4vFRu9AXUscZeqaX9INCwo44s54
OXBw+5mulEmTOEhTxXxDBZ1RPQwr3OZB5eZDopHeaI3EWCCizjEJ2g0UOBLa86QI
iJlhcnP9co/rJfvvgNskiOJvq3LCZUAUgyJVWbr8qQ8VQdBM465UDxbujSBsNmIc
i87KrbaPHMEbtK8WpC9o3lLE+sWEyrlSRB6dVi5j/cmXiKHuP+6c5+eE3VD0jcNK
+zCwwlOsq2Ndf8Gu3ATXt8h1KUMUdorDU6e34aSzXUqANz67m43LLAKBjP4GUqHk
tgOEdcD2yMy8QTW+y8pCQd5pSHqJBXeY60j3B/fLftuW134swKaByO16Cj5xryfR
piuV2Ddw6nXta90FPfczF5dU6lD7/5a9Dv/GjqU9K3yHDZTMYtKZ1wks1Av+BaZV
vWDhOOuH2z8KmZ5PFhNxFyeqladVDxBBIPXDNT1JN5bz0RkGifsy9SdoJNZg06Ee
ySlZdjpPi7OQwS/9vgSOzobBa/kVahxTOfc+qpkewg8jg3Sxa+eGTFabGfzMG/Hz
shpSQq7DTSWlODyOYxJ+X4bA6RL9qL2CSkrgwzmcqO/YFnesAXkE85i+P8xL0Qao
FRc1GudBqoquWMeKvarHtMTK7KdOEc7rLoVdXRaesmKoHFSRImQ4FfWBGJfElKgA
Bl3u6APWLFn4wrq9DLw/laPbobEcY8qEcjHvYQGQLjfLmkV9ztlJRUQgc8kbcWsy
cXH3XOQr23HY4QcraS/r1Rfc6KecQ1TlKRkmiqRjpofyKf4CfLYB+NDNKa0cIvy8
iAvq4c335ka5Typc/u3E0VQSX5GXI6s9CSKtyO6PnBAEo4ffj76IA+Y7g0O6Hy2+
OnbMInNByLNEzgi1qhX+pf1ivZY3/VhLDsoqpeAyV1Rr160WhHow8wt23IdrY/vL
6kdt7QuVXjtSAo4mA3ISwppIE42kYGfoyDlnZBO7WsXXQEk4Iei9IUBha5GeGiTk
V+no5UPF6YbcyTrUeyzi0sTxL18eiNeHjJBagyLEEkmk/AZz2s3QQ+MwKUaKMZO7
jS2u8RwLP3UHzZYKXVQT/SR/klvFpUyEDrobJwMT1cSu8tNqYbfWICT1vIzHFetP
C/JohrY/v23UpeHIP954q9Qw2iCQiIkrZHkVjHozIRPdPitCzfieTQj4HNF5eHid
sPvWrAVMwj+5sOsAoVkAEIKMqnZsaAQv+XRcMp27whUZrQgmVF5j9fD4zu3d6b+g
WZXiJD6hzxBhZ29gPJuRPScEgW/tOOQREKOzvhAjxfd5WUYbfF2dFcv1wkq4DUc9
1D4n5R5fEAFL67dzSdRQBxuFjWqW+jt5ZHKFOTmh9qlmKlP6OIxSd2gCPR/XK6gh
NOHTygpa7au9TJmsuquxexPlSm5NoT6kbyZ7Ln/w2foFJsiq3zVXJ8KcekykTHke
aIJId4bWbqXU6Cu9TER1V80khI339uts7uKycCS5izuFTZsuzQUBsGOCKBeamzGH
rMC5A/D2IYPwu5kfQIHQn46mamCiGnoPgKrOC8ZBHQrz92Wy+0B+xl8xyXi1Kfer
k1VD2vaZJsxCEzTWY2rMPTfZyvDIPRnmd7SB/L8HLwzZ8+JkNpyaVuOzYGVhGput
Wzw0xRE+mkElHQTqgVsqgUINDKqNMwSz1eL4u8tzJbA8aCr6T1YsivDW8VV+Ej4v
PchdEKrLb039eLKTZ4bVCARJXw0tUf7YUSPJ5bF4qTUc6SAF6t7nhePHGXfWFifc
MES2yvLCdsInbXHc7LDSX8Y35P6vJqUMnanEoJ8nN7uLI6y+++UKpZL9pqwdyTpT
6vfI+GqdVpy9o9asAMnSoQWNnwI8AzS9eqrxRdW6vaJfrZevaVatNkS06rGRQoGb
m3SJYhbmfbCDcKtuR0XCwIog9pyvPwtjv9TFmgMI/sGRW7d+muFARGThXPLCGMgz
V6rG806i6IbMZ9hCX8Mgejf/Xn/P2uLTuKVKsErS0uO9R+iFIW5BBwUjzYAYU/a5
y9TO5PObNGdrCZJ98ev0e2980LUTE5r3CBM+aqGIG8kuIjEDtghQiT+afxrKitw6
PGEsdArIANMHdSQCkujBT3VRvrmw96hNddkBPdEEVwBQqzbcHNDmM1v6xX/YotaA
qSQiW0AQdEtlC/j8w9bwXREbhFiVMOj2bIN2whRC0NDa/QdxztbNhfy8lpe/A1SZ
b8de/fQq9Mw5RrD0yACiPpEz87ggBNVHpC28Xx/EkpwqNU8lwipEI59HT5h4wRd+
GFkJltcf3yuRxelzbhtYahwZV0iLWaqD92cpG4k1IpTmrA7jlWlcrcGz8Dhxcbhu
pB3Xw+sCrRWlXnasLsPhdrYiSKFkuXWrUjUFfIqriZU79GDnNsCYZdoXCffUTJ56
0zzO8lWHpeWt35PYP6wdHGWCSPaj2p408K2QfUo5070SIHWOr5CDvxEywfTHj1Qr
Bmqs8TZN4VQxVu+a5l7Zhpfn3crCoki82LrCTEENlUKIBq6RFTNzgzRgsLZVrmvh
CXPXV6hj8rdsJpShnYcGftOpH8zlcfM6KoltvAPo/BLUxjZZvhvCoV0AGjcdEtm7
6cl1n7xzAUeFjYp5E1dqAdDk9z6UQHCb8NuCGaU9gFGaTdlpCxHxDXUWEFtzCzD6
Z/Ahkm+/Di+tjH/UguE1V8HIfQ426xox5g9iXwupt7cS2xJQo9qY7IO0US2pgaPd
JIY0r9D42TfC6nXmajVlLBeYmzL3FI5XLwtvWFiNFOwmL2Omqiu2TkDgzAuUP2gN
i/GaC4tnNgdgEQ4jcFIi6FSGGXKTIkYXmejE3i6WhgI3z9QsVrY77cJ0Q41iBxXb
kgM4A28SCxs73WxBb9rv2BGkaxIA8/Z39tfpe24ZGW9mV5jtmiq7ha9kFnQ8mPR2
vljQvn2UhkFcdC3UxL4Hmw7QcNRexm74+xsEek0Ver31sMcY9mZGOL/9xmIf/0ak
V3JuMeEgckZf1eNNkXfVYsT7WnTSit28LrIUZzvn3ualGswevHQVigeymy1W/eSp
4joAzP+9KtcdpUE7X901uhj4jNjLjirfx7WJjyXOypWoADi33HSpCcFhJ3qaAas3
LBbotExFsXrFLXN7VhIeotoAKoem/OhG2Y0nBui6KcLlq5BDSlESJa2l3r+ZKfjL
cRKQy+I33cQhMIlH0ej4tPCCIinDdjwhnSDDLpBrzNHRPzYblmGrHs6ikKhiMzWR
a6lMseAwlJJCLet5Akgo2HTn9LQiS4k6abhao/KSMl+W+eALpQahwAJPTgwuYSZM
btmptKdXedG3lL2iQDb+nzEY9BAw7nBmV6EVoODS2Byqu6TAUlEaRWGLW5WComWH
dXCmfVraDqtnBZ7vPQoODPw4YN9x/QVhuSCw9gGRIUfIGq7HUgv8mrNGWka19cDK
4KTlxNT0WWUpcj9HxNhYo29ZIn13thQAmVY1MbgLyjYn6gSM7+f9VwFJNoelbFoO
NhQjbx/rijt7kbHQI+DQGXgYwZ0ldNoq6SX+sX8+agvr8mlSVShKyiktX2iS/lFn
Us8bXIcldl0ZoScQmXG2AkqZtqZMzL3KBj/0MyoXep8nLY693MgIQ4pOFAGGvHXa
BfhlUC4yUxMHjkhWrRTfELX9iaZk6Yx4aN47JVSgt5jZcV4Glj/Knc2WyU47SZdX
BtML8B8wPAZvPjbgSphc13EueI9rheADhYRNcG1XqtygtO3C/lcRdqc5sFt4zKEV
FtQXPlg/wnCInd2tKpVRMtjPCEn0vU4tmF3rxytnfmJaZX2A8s2l9dWv3g+qqCBM
jH3bTlCRcGsx4LtqaLycfl54vTjtuy5BL/bWSie6J8cEmuoWwjFACgqKPhc1ajeI
Ul+YCoZGyKPygoqUH7NDHhQs7pBkJvjmMPHdsK5eX6qBFmCc17EfFkTU4EEkE6o/
SGvq5fRTA/Cg2suwi2WTjsrk5XX3P2Mtt8CwSMza+UqChYv32Z6A7MozduvAIhMj
ViGCkmrcTrVT0/Dm3nHBxsGd8WiecbwwbsBfklFJYQfoVFh7NwW8zeIGYaB/026z
Gc3txlNs6fn7F2Lp+uEo973JMgoFNGCGETWeznAXuqIZUKLrjlLDwMPqGg/t4N4c
r+VFZuB9n4J+SNqVE/vWbTmpz1q9O17gVnwYO+7dPzMBQQFOwMhXGMBFLmr4HTDC
IVDR1zc1yHXkOVBsol+QCQ0z2EBybh0dHl6Do6Z+nDsFhPDng2cjKXzVSN0MIHW4
NLZTM5Mree7+gm+VqgvwwN0KbaXlVqIWi0jim6NjC0r1Ne4IsGvfFK8trvVvCh/R
eG1uTcn43Kmks+e9HrntWS1laI9Xzw54AzCqH3sejni/uXZX62mPVpsGkzrte0wV
yLAPj0h3gP/B3h5FZ+wV0wX+5Ct1DosJ3ID3sFGAWQbat8uE4GoJwfHcXbAuiqFm
yQ/QDqL89LrZIM/ltC9ZhtVPeQx6QIHzMmygz+TGyyNEZ+OFCP+4S+pyBtLTvpFH
gcnCUxkdx3/hV7Uq+J0+iaTtKpW7lts4hBlzqBbPIZK+2/6Dcu+yPJMlDEgcfIOv
rtIo0GFUa4Jchsn4DR3imfQkUZ/1HPxtAJue1vblF6b+n1C8bIO0FidwSEnriGU7
09KZ9NtjjXVgGryeJnqvRIZ4mfPY0DFfxtMxRE3W4LfVRBqnNhDe20dLAGOnH4bT
V7HafJuYlxDDA9Cke7zOZ5sSyaefhq8tHfDF4gncUT5dsgV32UEvoC/9025+xdOK
4ZYUQKTvvbMNABzhk8p5+r0SSfJGRE0Qp/s3qgs6Vz75KCCPuffG8lUZSsk/k0GP
Kqr5jLXyzmTYjA2TyXG6n0X5E2nwXNVVOzMks92k1PNxkkig5Fu5+PhT7lOMadgS
CLloW2BeT8Le+ffYzysivhkPIRtRyhtGswWJl8ErfVi2tQSZWuHObQDHbUQBhG60
VDf14QNqoFor6naVVu3goABOOMVtItrigyS97iy4ldAMXh18OrvYU/nEQgutk/Nn
NIPLpJnfssPAJ5nqPwBYLAdP5kvDN2/5Zb25uyuolw13YuoF01a4hXYMCULcE0OW
HCny14DL+UhSp3aQIHv9ufu+xKz4bWFtedqoxjCWwpx29JWzS/DnOx9kMk96bU5s
wPD8NPU829AZHu3ilW/vZKmqgqH+4W9yautmzoTnbeS/GNw5WM5s6hcDOVpl2ARb
XAeUX1wzV277Djan6LQw5IE/Ghr0cPiGKeDEsjJD/7F/YaySp/JA40FuYW99yPYM
UpnO65qhmR/o0S4A87hwjI/e5E9K80jwMi+Yvs4ZGxC+VEJuyJ3j+MwmrBNSPhoK
Krr8ppQCLK5hXbEUu5nGMaT+MTEj+Pn+EAGrbqRxFMTwbaMftqIqKCwJ+gBnAYK1
eGHEe01gfiDqoGVc4BVEu9jGCgn8vfCYCUhE5eD6+PjR/HuHpSSfchu7XkwAvm8Y
Ndehwzt/NJ2u73785rt8KzoxD5JZhRxpV/ieYP6htdAjFyhhCo+/a6E82ENsPhq2
uGeZce/NblZO7PPJNmch6LK664QTUmi7rQtAk/4mp34pILCQNIk2VZNXa2V1onrv
4rAy1E8nalHWuVE1ueOLJrod7Ci8jwLe6NkYaIw75FH35+JbTHE6bi4lrkqit0WT
mYc73wQfhvxZOY71s/fyXcBDWBHVdJUgp6w+91NKIL+P7RQ/OB40HaC+YD1WKCJf
95R591Zi/MbQEQyCL5EWa/D4VYRTTepnbzwhi6nGTdbpwOmOAnDexvYTA72lJImN
2tVEbZa39G5OFieX7DUlqSBYfFhf2scoJ6SGQo1Fc4msYQnEDI/TUbbtDxwnKwdb
LgA8akypeAemQkGUgniWZlmbJUQKq9/lMtRObHz7fEbV+tmJt8pPahfEph8j7+Ef
l6mnar456krwYmhUvdJ07rkLPzQ6jFGh0SXx23sW4qmOXnyqp18UZ/U659EE/fDz
7VMkz1aj481eINUuXY7IPKkNl3/1WDCKqYRsRzT6jH2xWp/wPf7YVuudff3Eyjy+
f2DkhXTkZeKKJmME+p5Y7rietIjgN1s1kfywNBkSdhsH+fNXquDy/UfQCBOqAhJc
nuNT/2MluwaWU3mAkPJmPwBmGG9qQl6smwl6cC83uLG703KuFyrUuzojd2qICilN
M4xcbvOl9RNWMH82bme4UvtfZxg6f3dufzDUmVFWIqLmco62TTa7R4Da5xJrrBzg
rgnzLpaqPlFLPklAbso6hksIngnJHZrZQkklrGMqTSfWbBTl+Ping9LbrnR9KD4h
wRRUlgxaYiaX0pJKRGSBp+anwAHpeQUniZwBJIFmW7WyFiAGTZzuqfuc0KIHnEqo
QeylHYeIq07PgYC/zMngHfRFoMvXMOK4NinofcIjONWBB3ClGg3F4CuRl2SvRs7P
urCtC2WtbB1zORDhy3+n0KXPZ5dVRpauAY/UpRWyWbpk50OgdRxVyTA2TMVKtCCo
ivFhp3EOb0NILXP6cSMuTOOGwbZRdN+7+odaB58xjnouV0S9VzJV3qfVzAyMF5Wm
ENIMy8oI+VeOJQxoGCa8lKJrZIH+oEhwPKpIXNhoff7hNfA9ZxYg7YwkgS7gVQuD
Ymo/7cMWzMxqHhqoVlU6MxPlKu7JEvXrO9XMHyR0tifXVtIh7xdIGNVUN5XlkOLF
eXMu6X982/4MTSbrtgZ2wVwvIl/zeS83IdCPMMwXy6Mz4oGEAzwbG/LbL1DmJcQt
sRCOgRDoMDBs59wLbVTPLQE0x0MhAuR0E7OpBMdZodYIeZ2MPWN7sLvIk4j0lwTU
n3GQ84bRluZtntZf/rhNSV7oFqFhf+UK+M66c5FmJ9C8O4Mcw8oAL1TN3ang3k3u
D74zgpNnoqCiH8VeWtoVvCM8FBBxfJGQZLaLT4TM1g9bvPiqpEoyZvqYgx4W3VCC
Dxi9u02lJ6jIj9gBtjyVVUStWMCqrjCBsexLqc4j5FwOS+QxVuXVDwQRJoogCzov
ZMMeVT9Fgf53V55PNcb7M/xgkiU/dxJRN1qA2BEo4o5mSCVNmvkQEibQvJyeP0Th
bE0dwajmcUEho+X73hYDXnT48o8t29oJUDSVLl6dTvc8Ogx/JwiLGmstasABGYbi
CmW0q0HGTagRjdu6DemwT2A2S1esA2kBoBfb8WPsqeHupjGr1tXszv/3wD2KGl8Q
aRHSWMgOYITej1DeXy8eHdoFQPqers05mBw/+X/HzpagABF1qDYE60tzX0Bnz7he
L3eLOzfCjyRNcom6njHhEHlm0NoPVbcrEpMZxiPzhbwRF+mFXrBbqhzlTwPxqeiS
aaIqZ/aL0j6YTCXk7L6Gt3wQm2UJEh/bTeSCZv+OVbEnre8DaeV1DQkEQe3bEdVr
gzuS30cfp1QGLXwFkpeMPwCt2HDaR4mVMfwzcjbXhsiO8QraScfbd4pOu+Zxcun5
9T13DCg1AGe8uUWZQmuVEV+CFviJEVAReqQHTDaVFDuXcLp+KHHpMFuRnJu51UMD
Ns+zOAP9lLdXBT1T5nt+d4JsNLgMLNnH8oKV3IcxtmoDO3fjkSqGcTmVo4c9qMdI
wsUj03tkULOoPjnS8BHgmcru163sAr3jCR9RY2X4MdeA0Q9/GAArYS2aWJ2UhCrw
fxt16DtFvCNxR1DrJHaNkW6C5JAI6Cj7lbq7ZBIDlFkYrObG8dQ/TR4V4hmQH+AI
4u4mLTE9Rw0mNQI1PzkF/Px7dbfgdrFpAiZtoLatbKG5xb+z0IwmCFfYJoeksXCW
trOmJVKyIWzpCU6XnEeqwSJhgmck/RJiEqzb8APwfB8fqiPvexQFyPgi2yJrVgZQ
MfyXqbWDO7JCGkW0Ky0g9ZwyJUQAJboc4Hp9FozOKdFJZGpu2hFlaFa6fmPIVeXn
2vVys7o7tZFNNYnRQvSwa6cGukRa3kdc86mvusRpphtQYIgXGuDy4qCPZP1ItpOJ
wPMYdqsqAcuIjllO3hYHAX8oZApANZxV4CDwMmHpVVed4bz1anjz5Zg6IZbKc2PX
Kt8FhpCLjrVtFPObzSNK/nHp3CaIIsTEfGj4tSBNXos0OnR/oKUdWFNdReArO15I
tL/hgdU1qbayJBohW/Jk1KyApUTDEMoUL52HtT/tJ3xrFGmxiOVDJIDv5ce5iTGV
a/cAEr3AzrYd57EEgGmwxVK3vcfZy1+zQ3hmPlpB3yw2V5tn5aSfX//f+WEv8nuh
IQ9spMQ4ERJu3NgLlIiDkeqJtG8X/18Z09IyrUUUFqamBlg6xJLoEqwut5JidtEk
Q9sVUtglnWPO538bFecCL3gjyt67YZ2zbsoe0Zc3ivD+35TjNV0cZ+1aHjx/W0UO
Xo+FAppyc0eqwx8pBbReMDPm6UopSVoHmhEC0Eksv0xvfk5csprPLt35rWOD+vRg
5GFojSA2HPrMWshf7wxW7+nCrKEFp//HbDCZafDsJYJl8yYJA884V1rqCzWcmD7f
7ZdP0yYv1L3EDy1A9R9SOA8qGYDB7K5u+9ExuGQKgzmeOoIr+jvqA43uwaeRZpfz
yISYu2oZtBUGZuRf0m948mafMjrsIuWQuxMKijx6dWSuqWFo6ety/SEkM7b+7KRO
MJnIifTXV8XXOXjcvSooKEHxGOCPAHAULkt2acowx0GYZoprXaZwk0kFcNDFFt9R
LNFPqsImllHyvneG874ZAVfY8wTc3zIXaXRJk538USMmMWqvGbErt3M6VaRnmzrb
LLQnAdaudcbPYBdf+ZH78Bs7WKNQUjlbpOLLTIJjLHIGIeoPBHIxI8H4LQtZTF3d
9vKPJmCZ76CYsTMB2OwwC/DUzEUTt2XcYRqRg60hKTxUmJTPM3H5DPweJF4rXqcm
3s30XWk594pJAm5yrg/1oFBe5EzgkEuyA7XUnLunmJGiI8qk8RHAXJhVhw+6Ygqa
zF9/IJpUCgzvlSxoGpNI28hWxU9HexwxQwoRUIXl8p2YKwzsvnk7IgpUB5+DN5Fw
I6yeoScWnRrPmP/TuqWTdQ7rOp1LIq0gk1YH3pKKMbq+NJhm35X6I9IxvNBUx2VB
0wQmFaQN6xn1FnVQ00nyKj+I8GBPqCTkZg8vqLwjG4d4AuQvlapKkRWw7dkvSqpC
13auueYv2S0SIuxiTqA066B+KaYsBFqEQxaEmpKuMlIjdi4KgX2cy0+QRpjwF+sQ
dWpLX8eHLNDh3sNQVU8UdWbJAT8Be1R/+76U9asH04z9MaRnUNHEjL+4JNfXm/P7
McJxa5AsQlSF/TXBjBZrd/+yPRFcxv5QwI7/8B3IyqsbUrLbR92YvZwLrpIBpQza
vVwGUx6iqN3gVTSegXAI/UtJjlSWFsIOezGC2pUMnZB2k8kPzRGTE8Vos0u3VGpr
nEaVtvi3gEM/zX6FY6SvPbKC9eLjEuVf4uJweJ2DS8JaRnE8EBf78NHN4Jn+Cfc0
3NpGlx+vCA8ZJSCRIEbVsH/DqV90wkNm09THp2qAsCa9A4PqNMvHFGO3mHUI3OZy
+Ln62w8dWz+ja0Q+qU8+htFpVvmUszCaKrW3dn3wQ2WfNyyfU7qsKOuJ2tTgGijA
ZQtjFVloFE9Wm+IcemX9nA8U8GvIRq0UOld0qUgMc0MSak1wLKt+sTrkHqQZ8qbl
EIelFV4Um2g33sF1QYWAmb+pI8KR47+7U/Xvm3bGCJytXzZ47rLSl1Q1S3Z+imgO
MXTF1vPNpsjQ3hA6bG5ZBYO1/iYHG1O79/ip0QjEGxXyVq/JawSlWlo/jXx07XX6
RohwWhueknkbp8C3C5ezcA76/rQZ0b/nCk+SNSXfS0EMoFq2NTP24o/vasxLIHu1
OWeJZneOHBhVTvrq7vKL3MaFhwe3qGYBwQcFhWGtxVHmu8yexo9FrNoCWzC/+jGO
hg/L+oYfKcr5kzaFzIpCkmi1bmDsDpKtXzBlkDd1mDwp4YMqaH3CSGKHyxbkjbCN
rGbIvysfE/pnSGISzgP/aEm5352BXv2PsfR2PIjPEKevttuE6sD/atEYuaEwqcgU
S4bLMuzPkvpDVhohy5N16c7WRJQF+ZjxuuwOFVL13vjNyPwglwBJZTiBDhMOjaSD
X1ORXfoc72AQJKjmTivVfsK5bs5yW8D8Hs+TcXH0kRsglgM99Rf4HB50OdtS4r+m
wgop6E1UN9iQ4/CQ8T+DbbMTv9YWevusYRc6GqTv7syXscvLnVyc5rToYXvS5mCl
wZ8LCu6kzeBn6M3Nc1u0phBv13CZonZFjJcI/N/BXPY2uT7CtGH79XkrpV0YFLWm
6EjPnQY9xh9U30Qwnwg0MCqm80vv2yZOhhASvD2qffabxkCVZ3yrpaaPpH2SI4dO
T2OwOyNbUrSgC4c+S7y94zz/qdI+fv4Canc75uiX2TjNy+0EC7WMl2rH+h/ISOA1
NdbJL4I/72g6SozkcC5FC2LfXjog+5tPHMn+gcYCG9VfosOXz/ALUum+QGJyiQki
CQd5nl3o20VGhd+z/87r/Dkw9M63ZWmwPkPR/DH+hXXfFVMpeaPvretTMrUREOP7
KXZFdatoKePulEXFqF6SYP2aohw+wAl/oHLDedYVM/nMioWGt4CusYxNypB8/6+Z
vaq6fYQvcEQ7xhWARGuflZ6+mmoFhYyZyJ804JJX1oyXOXcy0wQlxzVm9BPTnk0y
L53IHZIPSs6Juuh6U1YyTuPnTCLovqCpRPdqtDgqmyDK0gSYHz43Q/Cap240Kb1F
Sp+aAFPT87xruLf+Y9YfVxFlSD19f1cpm/268jJvJMOsi1IU0mbChnc0Zeu35CdC
ABBVKQ6QdtTSmW7U0CdoE6i2pw1KE/9rRBRNx6ND05xq6xegIIpa8T9Yx/GM3YL4
RcFjYsb/X5ww0s5waATwH8bnm23uIcvwNNr8x8Pajp5aPodfuRWJwF+lKjLF2kDG
FBT8SvliP+e7HdApE472atAD5slM8WvmeyMaYg3gFqz0vsfeYStsObaLuXpH5S8L
GpRKi8vqgDCDmHbBI5MVLrGthP7CIO494wiKSm9nmJhy9fJ+orPNxWSamOhV07GT
GvC9axhfIQQFNXnrHyjMczOFAo+6LJZZw9NffYg4eSrIRZSCFM9bH/H0ZRlxyoXH
C/BZYphKXd9xJAdFNG23tkXc4HCnlNzFnXevOynpn6YJVn+D7JA8j25ucjb3K3HK
a6ty2Jv76Ajd7GrOU7YwxEGil72oEY4eHQLlRInYQSVA5MS8ZcFCaZnw5PClvxn1
dvt2+9+HtpeRwhRjCXH3PbV6HAxI7jBY3dpR81qS7GQXtET5Gs2Fv2HOfqM5kIwr
yDsgd62BA2jvizu902jfTVUb4j9ARG/Weck1Nz6WujaCMhbXqKgj3O2cknUj03Ta
KWym5k6cdFINEZDOvB9vgni3CacykYvraBeonzgPTSB8SToX1/a2sYKn7YELK4MK
XPtlzqvg5nfQVMfsZeH6p4F3QgXmo15q5mZiBirDLhx+/4chAxeDdUt5c04qrCN0
giSLWhkOOMFbfpHGEtsMWMOeFfVeVeDTMPnZf8cdtsSd4RnqeATkPRUtCeiDBfNE
t9azgZ7Hblfv4XneLOeUIoYxGZZeZmG1vVBw/Bz5IpZD5kp1zmu/0rgnO+PLl05a
g6ZAP6HIlofzsqDmg1CEUzdExsLQ89UEplaw3/NmT6fib5LFoe/+BdVVLE9Kq6So
lNnDCeR1RxROVLyg+IsS3pAmLNrwNBQxNoeXt1r/4QqjQsUkLMeLZmJc3gNXdAgY
4qK9vfQHIcINVeviyjE5XNcjZxxui5BUKQiuB8JlcxEgHoMZNNNg5IfySqqTsLWo
Cabppw0WraLksFTYYY8k4JjCFr/OuPsZj/Gp/l2/GI2fIvRedUB4AdcI+FpDZtJ9
QT7NNKEv0Ho/+TYkKl+wYTu5WfAcrE8SCuVOSl6EqkkxK8ExcGT0xY9m7tZ7dsRx
SoIqYL4/otGAzcbSPs8ambHV2Z7PdgwD1bnnSQ5X9Ara7rAqtP0bjSMcypcKt4ZZ
qH9vBjCMAnXNaHoAoufHioN9aoX5pkx1zNffPH0oiGYcBwQL0qpsY6kzba+/DoVj
pNYI/dyTCIHL0ypJYC7axeXFTZRTlRMa4LZ0XBGHk6j1o3DEg1YZinNmHlabWPTh
9a93ut5gL5c6bkvByFU9kYzXS3RT9+z9xXTCBipzj/jTkDDg/VyIp5gX+Axcv6PW
D9PHpUQUQkUtxh6jLp8JxjbD3Fqq5QLxFcXPVwmV9uAjC/MyJMDsjX8uMyvdFS7c
exbN0QlhU8RORjSfm4+xa8G4Ws92cyw4zJsMlI+Cag2/QSbQdwv5QyZOv/7lOlG5
SP57vXdq9mMpx/jFwB6rxMPs8/5YWiijIrvSSrFzy/ihllAOnrop4QMBf3bBXUyJ
GVNQRp06RU9IhkDSqZOZoB3k9yNT4M321RTYT6z7DUKuzUWdhB/rBWxR1Yk8hljO
B8GfzoAYeak8vVIY1yMCoTneqn6SV2p4eJCi6bY+XugdXu5Fj0SC8gSP7jHNTj2Y
exWhldLwb0lOnQRnfR4jwFDmen08vnPeOowL+ozfxqON8ZTNgWSJzpHE0ie/HGM7
TWznDVGGzKpUZtskxH8CF+BDqkWkbmJ1FRH2qqEBkQLvpvoP2VLz2jdKzPcGtzLf
Gb1GoqiMBp++nygYhQGhB7IjwDR8drNv3uMYlCf+/mT9UJEhrBzP+ouQALDOUqTX
FLAUd6cBnEj0MUH7Gb50FTFr6d3yxNn8RTSqrHvB4BH1Xyb/w1DoYmKVdHcwrnBQ
olO5lcV550eYWdC8ocD9SHeO/u+V/EHmLa5n5PUCO+xMV2FpyDwEyGmhNZ53e3/J
dJQGMebPBPqsUyzNLyGNZh4K82BIbat9SDlkBGxI9OwEgpiWfHsxhVSnfYFl5Jvm
cWBDuPfLYi6JUtFkH4SG3/jzXATbKP5xVX9Y/Z/xa2YxIRDoa0oa+0fipPYClaVM
rf2n1qSwcvOHAZA3Btq66cYEemg8Mw9ATjfWmfgrg1wnXDEfXUJnqMQxJDzkuC71
I4sUukwNL27jC/M4mYjjX3cbD9b1utJD6PMGNAX+7j7NuRebRoas2ICsnQwy5MIP
tlstJx25fdVxXoBhL2iJflozbwmsN0xCFF2I3WcL1lVXb6beNtCBw4ATuUksz1jj
77dgQBDc1SHgTYcSQ8iguY+Le2DjPVnhf2uVec+VPobjC3YPYv+8zL8RfeWulZZL
9/tjPMysNzRy0Q6cJXgGx9dspdpvcMK4QUokxN651xj89VwD60qwVNJgDDGm3oiU
T1ehbVxsxl1YcfXWmWpdno++ThDo97dXBCCamDSiY7V3lMoycK2lhQX3BIFJylIo
wFXQuLWopG1mNGAe62t1qzYU4pY1GgHUmpFsDLduvWexDw38BgG/E1YDLbYvtq9a
A8sCus2KI8+k80+YRcSEs1Vy+HPr59HA1zQPY553AxLu8NVT1fCEVU7Qhrz8MAC0
4SyLCH1Vm8w+Y8eB/qsbzVi3NrkbcRaMwwhHxwFEuyDx6iiWc18ASUpgiWsR91gV
Dyf9WtBpbQl6gVRTTmrtHjVq4VajmQ4DQNEvYgEPXBAXePiFf8ZifMICAaoDHJCV
5TVCa7H9N9s5H8IYEJinUFkrZ5UVhRFyhgi+IASPK3lBQeYZPnTM0yJhit/F7g5i
5j0O9buqXOuFEWpyUMDJqGQJcxSaVPK8WWjsUrbKf7xnqB8iefFr831BDjHCa3D7
ERC7aAJLt0bjyYxZj89kgqXmST8tkAfAORsNMy6bJrw7UGpPjpFsfKTHQHxFI8DH
4NH+DyKvxoBaC5KGv3PGqVj5c2/TIYpfQBBX4is/Zw3m83YQ0UNgpsETsyjDpTXB
fT6qJLpFOIVxJO6NQcMw8PHR9lP9tjSplolBJJA7kSj2/SKIvxWzJgq5+mF6tSrS
gR0HwNmisHNzm7eJf2x1TQ9LklbNnTXBYAQaq7Zz8UGbcANI5IbIb5aYzkr7NSsm
dIhgne155ABNVofsx+CiGsVeJhBFM96lEqSV/8+RC5Tc/YtT7POwnGLWtxj5027I
uqb1t0QsuSwBoFepR9N3vGDrGwmTTyUMxWHraFmT+GBC5eT7o0nxxAwcnSHWWBD0
XIKOhU8mTN3//R6PB3lNVetImxbSyBvq2thS3S1l3b3OLZJw1QOVh5muFWzMegN8
Zz4pEgffdII242OtMpO1qyzZw5uZCDEWjbvJz0lCghrHv2phUjyLyi1rIuHI1gPr
h2aEyveetStLQXMYy3ZX0kleXTvP0WUubnKhk1Z4/OLuzlobF9fexge5E2sQ8wW2
PA+sKh/FhQs+j+M2+Z2aT2/ZAL281PpBPyaEBNeuSzZY42t4dbzcVEjyzjB7HBKJ
7+dSIW56OyyHRsNh5qILzzhqasQciLvYZUQ9sRXNknbiweicFDasdmbyyuOZWQi5
jh2N9DAB7BYMHRFHU3MhSuvLQE0TFfXRCqSVlxk4qhTwSae4ACINKWN+l/VhYz2u
WexSZX2kGU88R4ytvr/N9WioPPd87uCbf4ATMT0lBvpnGTYDDEM3TOVMb0LI0UMZ
nd0RFcrUziTYGlgDzD1iISKrDFzUr0mEuX8YTFnOfd7rsN0FwCghf34S5tZtqj/q
Vv9brPKtyLbOmWByz9Bzky51KvyIJgs/ktuXtQNy0r1E/sWDzkAp9wZBoUj6EhPO
WTUogoufhyWMm4Ful0K/sMgATir/tc2rPd6yajofETfyvz/hKVnaSfRnN5977iTq
YVOA8zQ9QmcjsLz1ajvuBvK2+AWTSeJdHFTi6GbqsHJJhmntpE39cV8n4tZtOD7W
fSz/VdWn9N4RFsGWVYiC0i2O9sI7ogepDgUD6TP/9snH2NtHMmueJCGZ5dgNNIgG
rC3JlGVHq87q9dRSoknt068eC29vmR0QMN4CKGnJWe9M4F+mC9SIb+nVfmh8DioO
et7NoxCTYGifY/xifMo8qRqKuFb4zllUhD3UrwFkjPftyo2IONhS05CC0Xm1h9BM
qV+0hAKhrrWzGLaQu08zhd4C9tkdteBmkm2rJcjd/uDv4L2uy3iFQDo2X1pPpOAi
o+4s88qktTfCpHXU5xStb6SslNGnkoM/bJWsWVtaAc4DnusLNrEl0x6M0hDIHbbc
7SbzHzj4d09CL6LZ5eW6Djs81dYC6ChXTqWELLw1+SPyP0byj4j9GNFYKI7R5Rdd
dH2Fct/gUESKQd3g1meQ+o9x2AoTbact2KoJvlldSqqfhuzJQVPLug8l6nBXSPNv
1ng2OF+2+qBJHGc2RtKHRSFY2r2gUVYEirgTWfbRyBnk1l6xnJigmsuMqifSz/hn
BNMsqpngj2XrL9G0kGGm+fxBsylummpcIxpXuCXP3SFGeHq8jOgVgFKQbIxnAlVv
fLRLvt8qwIndCy4WUN6J/pynMdSuij/D0vNae9NaAPah5iWBkquJ4Z6qnI3KvgK1
Gxm8LCwH5VGMdcthwnySfk354rh+sttIHYCvh5NpdTwcavVzBbj4IlNtVKMACnJ6
ZxM8GCbzWQmovautoYfTFxfO4CGbcKlGYbu9X4NsKKJVWIoz9cVvVaRcQjEqCyq8
X/AWrhUEkKewZzbrVAFz4tDNTnKWOVFAAELR3TCQRqxLNOQoWSwo1mL1QMnovUtZ
otwGHx6LQn3u18tJAXR51z/YIMySZvKUyrbLbDpjgvpSXilb8isPnjQL+ldRPVRF
ebXrjT1lHcTyc4WoZznfcOHy0pCYCsJThQfUPrvVb9eRrzz0afZ7b8ogtdRiDY36
qZ05qzYVBzU0jwLflaC5/zVxEG3fVYVbdE3pg9NQv9J+EPmQZd1ikhJ3KqZmNTMM
M+xqEHfl3GpdCj66AKsQVJ9vNQh3khA7+9jd8lgRa78lBjUe6k0WlwLB79QKYqgd
BDmj0QUfisRrwZQV5jn1fEmYq92JxE/JYI/iLjfofEPKvtUi+KzKPXHIXkq7izJ+
ftTY3GrHkfzM9cItw05PeQCvfo45rWRpmD7YMrccqE2Sui+mtIMEKl3p/78/Lhws
OUe/NDGzqz9HcQHM9xi3V2+Tov7/GO2Mw3pduOSmpVw7SuPBxBY1NP/plwTFbxxw
p/XVQoW9JXS4VVpxyPVwUTRhr2Kzv3Jd5Bfdolx+N+/VPnZlZC+bfHwV5NAXzJJv
iSKbG7psxW82eZc9RdwB/62a0aCMMVdKUw70xBrNzOd0ITsULkDEOQiZB23wT4L5
0LSop6JwWgMFSp/7TT2O+VnPPqrHfLzuaHMX6pdZ8iGnwmFBbPDRqbk3KkSdUgSG
Skt8cawDoLhpNB2D4pV6ndk5V4SekhQcgYv7SUxPVcI5hH9NZPLnpVe+POM4kDLK
QYaSgDX0B3JIpflkto7HACmM8fBegYqwbT04SAWwqLEoTcqrkthSsahMYpN+gvPV
Y+JIJGCf68sb5JqVu23nJDfnjo3LjgzFS0yrjXiFpscnR1Wh7YaeKV4CSnTu6hCc
fxeeQhg6v7gCEa2ztl8fcCV4hx1uLiV+kMcLhpIqjy7TKIs35ggkUOlURbVWPDZW
7QeznafXeDT0NDpupgT0RcMcigqezCKBWbQMoabyObG2b0dF6MctMbLafMxZRyrA
l2Ktsb0lt26cbyLgHwGV4lnbrI2shL+2DU+ygOzphoSPUtExNKYRIgLqpaql8Qvj
pMH3eOkgW0xZGZiIJGGiNZK8t/XDMJs4MCT9VDBxZG232T8Nd4vtCpkg8gH8zoCX
smNTQPOf7Ky4QREJ0nllNPqkWMBsJuMFYPLVjwC8kzDbzsd8HTURNo6TMjX6++5t
6fIPqVEy9A/RDB8+MztUN4W9UWn2mIBmSn0T4ajbwajwAb8tM+fPlWdgeLgKtTVr
HyL5B7hsdbttAeIzuJMAVwfNyyrqZ42bX6u5SEmy6VtK6Cd+/2ahAPUZmVgB1FDO
EsJsE59F6rWEapLEvQduh3rkOWTVnOfLbTqXtY1/H5VtDruLunap/YVC81jNe8T9
0kvzzhN0ezyPsgW1vE0K2hI9btJKlXmIiWYXUW8yLfVu4lg4npFIuuJ4LXL1NUWY
IHFqRcUpOAdW5uN4Cv7HHwrzcvuUseeuYMiK4AF0Yv/w/8OiLNVDk+iYSQJI7GOX
ghCrkYpMOyX4wuKd6YFzeJRjPNX4KSy9IW2AaDx9ovs4BfBxQHVofis/nYwYftqi
23klpvlLC2V+nAbLGXiH9hbLqNO1uTeZnZzegOaO0/J92roQ2hCDqaCZn6h5QqJT
O/d88NZiy0R9dgqGsuOXwadL4NFjLYlzr/3NoYCnHzSNJrOnYEXjWyt6isx4YqL7
RTMlhLY13C+5HHuju75rJkNCXiCGct9SV9zHgC4OyusMl6jSo6aRPzg4fVVDG97H
RgwrEaQVL2K2EzlcDoq0wPVePSWFr735ozlu969UBNaxj33J6kdRzyLkWypbqxYG
Ra1+qbs3SEdkmoYR+bYowlVfQf+gNu/v8jURzQ9XykO1eFoxR/D8ToeETxx7/5F+
+xmQLF/eCh6jiN/10nG5iy18FTicIRfTovhDQZxXWRuOWwuIxXBzKYRPkqzB0K8W
CR57icMjn8dksPlqwWssT0NCoivmvrQOpImCP11VBM5gTa+xgzE3Qw429aHjwraG
F8bHpJ3kyHTvsRktWl2cOeRBiC7hMfTKN3hVdmwRE5MzieHVywDxrP5oYau523cR
7DrF+Q7gzjMLE3P18ppFi6LSbHoc3mpJfyDJNK6sNGB7bzTbLWwnJGr8CAC7IBxD
0j89irIGtFNlWJqAuRnNmemPAPYbn7x714LAk0y7Hovq6fOD4dYUG1qT68XByLzE
4P1VVonr/kv4o0LjbbKNXoUtSkLokbffwFCs7okZrrf2+oV8HUC+zoD+rxqm8bhz
uybp2i7ovLEXvK5mAdVl++1x0qEyPLSaG3ya2oulwrYUYLX5kuLVqzJCbXKFA735
OaC3qi503jCQOJoDhrjfY1MCIZYYR/BU/PkqFaHceFwxTxyOdulTdIr+gBLf7UT3
E+a3E6tCJHeJTKSFX0570wTWSGX+CmKg3RWIJ9x4v7B30yc6BuUkyLdhfyGxXqdf
rWOhG9va3qn6GUE6bINCUhe372mnvhgSS4+8eu3ySJQjNBsja3IPLkMQ16O7uadW
zmOLay1hD2iKpxG2l9+E6HezTJKOa0aiINfBmdmpDA/quDtYVg9FGElRzKRIXL8o
5kBX2USOlY5PabMyy/excerA3fwK/szAd9ly8RVr9Ety16ZvtksEyL9lApKynmBZ
MUpZpryZsGlpnBwZuivpMQOfkoctp9rC6m8Yc5yYAjy7ht4vAzi2e7efsLTLlr4v
jquTswykDrxeqm35jSQnCGuxC/Jb1AFgC5YRnC5bYvaaP+qerU+w1tc6Iu79rt4W
eDL9IRPmQ/sNr4P39u2BryM++a1T60BgI2G+l6VVuYqrAt31EBy+zfmMRYYYHpSs
+cdTCb6zlS5SdS2PVIVsuW5Orr76/VsGKvWenPO3EOLu5eY0JRL3MHMqZYursD70
UI/4aQdw2hSlAWAoWYa2lX6HlQrzo7JVaYRWr5wT5aS7QYa2R2xuv8lWOfej04Ok
3OPSlaNrwBHCKqryzGvtPf8m2PZOkz6fsfM2Q/pXmd9mdjTD5pLcUyKRr3xVIOBs
XCD632XfQjwdwED/qU5fImpTWWWRoEFtO6JjvJ0k5R05+lUqLsFgTLIFuHEeZrEo
1O7vHK55xlJLMYCgMWp6IYZ2Dxqo91BFHFwKp9VjE+jXW4KQdgpU9yr0yYLrVHzY
yLF6ngS+KccKqLXpPzVxXf7xCckXnlIseDb7iEJzZVmngR1FnukLclcBeuwcfG8d
8mGOSRswRFu506suj/8wLFsnKkvlDfNr5BUQDTubISlq4rfB89a2qhtSueRCFO7S
9h8ghDhK6j2usswdkKIXm5t9UNxEx/xcrT+bX2QL9eAr+cU1c+rRMuCVyZOSl+qW
d+XEezVKbCt6C1UwH0rwSSesh59G+GjxyaDXHz8bDTZuYhjouwAvDZGWN+ejtxSh
qZUvmWNjqB3jgXSQXUeSCZ+pTr4o4fPmNfsrM97ImPdk1D2L/lRkHPNx/8Zmw4o3
/aKq0kB2UnusRHzTogmh3RJFt2aJIO6bqQEMcijJBEe+J/C3IGr0U1NCcsjx7HFH
HgyDAKj6Zz5exrF9LjShOE+eL8Ik60dhXnh943zm0DS8nFnF1R9hYBec7QwoBhbF
2acMpT2z9hH+7yMPUoYu1YFmoIrn108R3hZtcihxJZyawKNcQfFWmfKC/L0hPhAl
YknEJhJ/qKWZA2E7E1enMeA6s6OE0Ny+9pBiSA9fLxNozvXRqABoN9cr88lga8jM
L7QaePeyVwIzWA24fsiFIXbO2eK9NorkAtQIpvjTxvhYTmgiKa2NtoZ+aZK//Mxm
mxjGIhFt1hrjKw27ah5/g0d+X/5vZCo9qO17fMG4xPVi9HRE3a9yBaE2Z+zk9pR6
9FRrk7HGK3DxdYMYprpSgXnkO119VtMLOH+6bFgj7Webk4+J5t54TVCfFDLl21m4
0lDo/0nnN+corgBRdCEFjc6VEHdyYvanR5wkRz5KSPbAg5bfpaOgtB57fG446ILx
VlxtxxxgqpW3J/0GJg9Y+A8xXvbvQg3VbTljjlZMRegVeZDqYyKB5EbGmz1P2g7Y
4hrjOAYuLivQZGABKHL1v5+HoXfMyQyWC6WKh1yQ9IdVB6NuTrqDWeJg7F9Ty5+h
B7ra9VXUhKzZRcq4gMGw4+nSTHd66ipLI7mZU9px2ubNAc1djoherssO5xel8+VT
BcEE44lHhLHr/wwVS2lohlX1wpPEk2b62NH1p/aN0lSd/RLhY783vcLRdenImg7/
Gb33LywsmjCmYtg47HHJe8Zw8k8eZJj/t4UhppPrt5LlJgM1doM7kTIhPphynHF3
TZszPZXKkrUkGDF45gnttUL1pefdwSoCxfe3WlLWRhIR3nEkn1Bu9gxfKuZtfvRw
6lfjhMeiIOMmvCZZbWh8k4Wpd644qADPRNpHICIAH+wtAx7BWrV/8Dgd61XsMp/n
P+qKdY9/J13WY6qa/OayDSlW/PW4ADEhZ7MrIhU0JWo/KMUEhVagJG3owiHYJOnL
214fNKKRHanva+j1O7cKYrydX/vLzUgh7Y6TvrnQrifVGnM1NR4luCR8Dub740ji
R8umkq1d2/vwmXrjJve0d4LLUvZnL8dkrcc8+CwcoTc5XyHHYivtuaNfTpGbSV/U
FK8ighG7lyO855aj/0otxEs71itYpThXrzDD6qs3NQNl0q26fMzYSdVpH1WNXSZM
8AlJCalKZBJtxeLu5BQubvfSe81LS4n7ZyS0BAk9GeAOIsEiKXbsBH88XOw6xesN
WJ8NTVQ8VmqUi9RH7wpgcMot1VTDeFj0zlGfbm+1Ht73+Xlwl522DH+p2KV3SZG0
ogSBx8llCr6Cl8fvgvJJPhljmlta1Wqz/eBQzFWIYD7FsSyqLSIwENyNtcMXA2Re
vq9Cl26YRpejXPQ8ieq5iBnUcGBnZhNJmNseLJwvG84MDErFA3r/koL8Ok7cbC3j
iHeti6Yaj0FIKdHk4zw01GlZ6mNXCboDXEzz9nhLgWxBkPKX5TsAOU8nGYsU0wXk
xEYL1WVJp391333Ik9OTjOX8NwIgqyFK/ZBupgb/ayd11drDC+x9RrDaIkjWtDZr
FT21DpF1ze1/NFi55Si+ubh6GJ0yx7g2fUt9ipOe4knfqYyojQt11nPi6JevD57+
Ioiik53W14LYHWHtvPylmoh2MmsN8nLNPl4nI+WalRFK9xRDRNmEMeeVtVdjrhVX
Qc1o3w6KDlbaHFMcJsrLD3+QDQZDFTwcYiPIP0F5Xv6d2kK3M3WtBKIuD841jnlB
HjjyPDLAj8vJoZSKK5yeg+8NNBdrbXG9R9cBk4NMxFkyfcwLMDCvx5lK9Kh+ynGT
O3kam/cpk+YxeCDTpVgyq8x/GlSTxcbcqwOb3WrL0VM6Oj3tWnHXMj3d2BJ/dDJt
Jf9EDjNcN4gCqFeuL4WONF9RXIaKsmXxHKZkKhxfbBEKSa3hkCmmoucUElJMRVox
+02h3qY/x1kuvW5vhSbx3bdqdXrfpTZIzTqRR1hkoGCNONExv/WA23ZwChujJQop
01SrYMcfIPq52fnWc1AjjwMxYEtM+7I/VndaGgSSSO13Ms5HOa2Qfn0+/U8+tRzz
ew1uEVrWIUUeUZ49iM+rxqDOm2YmkGuzYSLm8xYXTIk9zWj+rTimIU5hdHePJJTX
0w3K97JoLeusAaWhr8Bc4IePh/nabtIgjYm8vdQ67Bn3zUHrqGL1CO/Anrlg2JKi
UrgNH7NU7pXhkY1q+mzBjQxLN6Yqlq2N9l039YY21MteLFSB2X6x53adPPzCl7r9
jbZHRYGYVaZahzmZvb/Hae6ZTOUaGB5Mfn8X4XZ8D7Bng6ZGLilgZ+xluQ+O/5ps
A4DRmofF+8+4JZSQwWMZXdTIJ087E+Tqzsuszpjvw5VkEpprGB1VdoB4KeQ7xADP
HeadHbkIaqiNUS1TYfXTkAPyBkahe/Ao9lDYe/HpjBxFkcoFISPqYoPHBllzg7Kb
126HE2Xbo62Crg53lMAn03sBrpWfQFdjCrLIaHvzaPn5KMjdkXfDgQ121Cju5n0e
PH1WJepn/6tuWqkOueHBhlZmnv13f/K5H2T+cY5vMPhkORGhhhfax5lKTV49HN1H
FyoC36MzQ5y7dBMeu1/BC9NkFgpYFDRI67CDt9qCDqkxqvmkwQIHd6cINOfp9gJq
4p1XmSuGQj/Y1/tggo+dRkLdYD1BPZqec0o38PI4AKtg3/2Q9pULSIcjKw0WYwaz
yvCEJ8zYVYajRURo07NcGBXL0rI3NR7t1k9kLPlfzNVr3wZWI02l8/fjfVU8sMF8
+m8lJrFzDp4jAYhznCLhcqqZcVVbw/2cYsXBPSqXWjSNEyb2ukHMM6AMZwf37iQh
36t0SpW4EyCVv7Vfg6RpbDPxToVAq0KaQ4hdmNyJPip7QfyBXTxxCAI66W0yMjwZ
MD2Qe8Du4NZjo7c21SO/XPEh1Yk0YYDH1VB6jT6BJMGRzWZmUXg8bDmZ35+nAM1u
gxJaKLitf2dZGH3CHtQbDn4/2nAUOYeyWQ6I3jR1YnsSIP5R3jTaAG0RCF71iraC
6gJhtzJ+BuyfdB/O0GTRQ2elgxkwrId1P/hr7bRS10EgjAL0xwaFCGxdL2w6e6O+
1u+nGTc8eJuAkhxfInzznUjJhWamvC3iShlWqMzltiM50qsDU292xpmUfergqZ/X
i71m1KiDKNaOVHVUUtSae2mzArn/MYBKLdWY2fojuonEp9/p2aal4waBwgWrEL7k
wHCwe7oxyD1M7cu7mVKRRybEZ1p1L8pQHzW5mvTXiUl4s7Ns8sCGrz5mzaJpUb0Q
b7SCk+KhJsQnzGHoMma212sx4vVOadWdaz9y8VZldDm42n2TZaBB+t1CQRAO9NOC
+Wv2TO7s2Vv8XCobH+fhuFl0KN3AtapVUP53X8fIA12Go6uPFLmE8vli945Fo+9p
96FNbE9SQyOiixm2VDODUCvosJHEh8ytwtbje9oCQt/HkO9XwlxJ682F/EbUhKvB
K4N/Un+xIBGFgSzrVyg87e2DCGid1ZnubQc7d+c8Vfq341krJirLuch6Emc41eDS
nZsR+DtGrmRyYvNQPo+lon4f0e4figbBoD9RxvM4IyXr6qez24aTE4E5gX2j4apg
XTWrtA7cibzKVyJz/Ve5o7ujAudjLiRJIs0iKDIsk2XbsIG6tPbtM9vRJWjm16hX
Wj+T7o1uTtD8QliwozkVeX3LhLErfpUNArLNBpWI5Y4FJJeABt5QJmV3imJ7z/0U
MjjXGH0/4ftJFzj/onSu+XA7NbXLRowU35haZfQFq935wk7gJPlghu5o9NmHwtu2
5wKVUnArR/mATPrdc6fqbd9yWHO+fmZ+pbCl5eyFgbBskBE+u4KUlxUinMoL4mLL
ljny/Eica7ZFSyB/2R1hTHd/nI5OjHxQr7o/jow93WuVRX7IaWyhnrAR43tZHrSs
YeydO/gkCOImwok+j+rMDTvo+MkRD9ZCFiVNXDFIpUxr3DmcfNaGe4i5gs4KqaW/
f9hQR5ompzkMd0r4XLmh/56fzmm/Q/1h4eip1pbiOuPOrRP0Mj2wTAD5d4xlrckO
gpJ8i8xbiH6s87+HrT6p99olURXEeVFRMNsPKAVI7NaRml1uYNflKXstfQI6vCT4
XWobGmmoojzkRFYfj+p4vlXzDfXppq2QIXgz8RZZcoks5Bsors3H6Jygb6vvI97R
rj2WHTcDFseLYdDuJVrblja8SAWmEHKm7LUN8U9gsSDdpg7HbgPWjhQw3vnJax0m
HS4mQ7i8sECSlIP19/Id7ieZAzpftfPhFtVg7AfwTZaPM78E8m/10ZyuX9u/GOpa
+ffLdgLSkdkuDPpWygGDs/BNuceRtpRLSLCU58xUshXWhxPINnjWHHOCWU96gjBc
gJKzcBTxlEnlGmEMNmFO+7806dzOixoQNRmXvYbfX4UmXFEm73kNxk4qoGI1rCZy
+eiDZRc5gMmkDbuMQUUI7q3anKPZvI9vW7Bf3TBgHJ8hCut/dlqVi81W2hiy4JYd
MYt2pb/ehJxrp+xBnR6Tz7r/cyTQYJkAsp/z4PrtOjkHjUJL6r3wd6qkET+L6eLC
TOnxq78Qw+pN7yQ+HXlNdu0e5JBe8kLmNnt1M92Zjb4822GeDREPxGXSuAhlufz8
5igQb+TxiIprJhZYF/Sxt/CAioH44S/qVR96H/bZKO8RXo0TpI5Yj1aCe676R0tf
puxWNOPZyp7oKpgc47fYZBxHYYCqNImnvh+vzr+6Itfd/Wdmsydq5eDg0/jW6ZzF
euH8rRVdWejSNqVMbH7LU/ZVaiwZ/dJCTrZOwgHHjQGjfRdg9szdW9Q5vjWABtmm
hvPFE+fwtd/X4UR7cpcZeixX6vy9TtajiUbezH2NjRBdKZSNhqc2RGc19khKz3Gd
UA+CAFObEHSwTL3ZXsY9X7091T2zqrCtAQnyo47fOo5kjzMy0p7lRk23MHf/+FH8
3edUzYWIi5Y4PS/p8q4UzyRL0nLITtxKnBJfIfJYbcLSxO2Wpf8B9OCBTuzl9SSC
7mMiRYsqCp1HGLcZAETRvq00hXp1J4thVQbM/tdSuj0xLEMkHAyRwSZSkzOVT4KN
vpknKPJn8WAPgr+aCF3BGfsXqCHrkhSWafxGDUl5jSZzpRpQ5/4n+UvhZypNMhLx
q8l7r8/+3dYDRuEM9b3ZYskdWTliaHE/5Do/TKCXf2MpbkDOmXJD3iJsL5+xISEN
idbz9mou33T6Npw2mF7Y686Qk+f2CIPsZfnQNJw5ZHzyRYWF/evRVqMt9Yw+/df4
xdcqsZOXv+gdA/iqe9vdp6VSFQMGyEHcpNy62A9Wtxnabd6gtpmMFjRN/SYuAEwO
/AYHgC4CNR4T7xO2E7nWSle4mmh5yvhHdQCKXtVZQDDhQa1WzxNyZnaCxfw/+YtS
tlVUvpl6vtb8uB5zeCUZE6ZM2mxzxZHBMitqadri4c1obxPCQSxVU9N2xDgaImXH
yCdrYRsbuDqDPf6fWD5IkQChxYLkc6LD+f9ztwVEoURYaworOP8aZh7kkGb8AZFI
WCQqNMQP1lRW7t1zcVQ2CYeFYwhw6HGTl44q8vhSJqUdkVEE9Wp8LV5UT0om4o1/
RdqJH27GT7WnHHiAOO5tiNAi7HTxZpoSNhPUjjTaaLPuPgvGTWf4w8nKqUgVFtRc
/1eDB/T1UjaTeXXd50T90LeVOry6rHkSof03Dq+bluBsY5GNbVWs2wVq4g8fnq7m
lgKjUvFzq92+jI8jnc/UkxvJwd5M4nLC3gk/Mp7UBussRgMOKgmEsyTiJQJiKylI
3LcSM46KOiUeoToKQpTWpuSuMrfa7qJdD9fkMSYMvwAucXvDxIS5wAkz6aBhSyFy
zO8IogAc/GJaRvFtZlgRar1SDBPjKPR6QZClIVBeobfq7P957DNvy84iXHH3Ml90
K/3YeOUB+6CrhwaCtSVd2zlIFsWPCkuk0vM+AKX7EWMxb6+7bsm6keW3ez+DYNWT
HSsmPRHWICFITyl4seztIpZk7ezwk67CxecGlMXIqG0OFOpSNzLkwt63fupiUIc6
BWpKXUB4Vc2MejsvPiT8egnmgbcL+KXc0YGj2X9dpCQaT/OCKhfVFmzhSsHHArjg
uD20oye5qhg9/GOEI9LppctbRg8h2oBwl+Qm4OI2JNBS0TkCRfSFRFfhIpkGhOev
7UwCTdBeposQaooKYAmEuxvelfrsiKEPdwEPTUTBUvsWfKHTX7H0dc58Xc9DIVCj
L35Glfebnwx95fCEpFXgQObt2NKRfG1AA3cRiH97xcrnaocCGvC5MuViKw0L9pHy
wgbocq6K4ZVV8E6c5puPoGjR47AhjuZcc+u9CD465587zFu2MvFy0NOZqdpAtNle
/RVX3szE/AA9sbL19YhGbueJzYaJBT+D5aDXaC28T4SFf/86tBkyd+PKKpfwgGWG
TAMUN6Uq9Vd+YZL4QuaZ8SHZ/F3xfsJE0Px96UhDYFtkw3bLBW0kNpB9z0qsKyet
S0OJSdIGADCYETm3SFNmOex+N/NdcXfQUNH4ocKFn7nqpQXcnTWq/kzFEytSWPAc
bNjRk1r1dlL9KM+hfBJsFa8k7LfA4QshyBOSSGAVc2eXjZPhvjsGJCxpnVbwl/hV
c8YBvUr2hcMnu3DHwoROaX8jiGwms/RKvM7qOAB0MvvdF0kXX3kL1mljHI4ibPj5
iNbrdpVtiqVQ/xo1xbStldw0d0rh2vs0TYqs5T4BNNKbZT4H3PCjSjQQ9I469unT
f5PURizb5LWP8a7mx4qn3c+89/3fqVXeAAGo4QtI+ikTK8cwQNp/ZLbKduxL+3Ef
AR7AC1GNIkyK/LEYl8eGVrbtQuj8S8YO1bRcevy/SaAgEDjtbnnLP19DbK5pKK/f
a9s1U98qH8vIveZ/FgNMXZZqX6fwHKtb5rNnAdsKS7p8GmsRdmpxbEBjTrTCgG5W
yOFRCPdowMer4LFOFW1UjdTYvzkjFLvprCsjbaGCN1sZ6suk9K28y371V5tPxNAg
lfB1XYKiv5n4fm0+gHEGmjnqBxiv1j9wWjZWG9gx9ZOtn06XuUNhR54zI53cP/KW
WLiqg9NrBjOQWJPc6RIijlIdpqcX3x7OUNCCVhcYeYguLCxv2BpmGjT7PYesr8Rj
fmAh4/URkfFHB3vfHhEnmUP6rPBt61Le6RWn26101m30Jjm3PGy6cSzeA2e+EBdz
eKpWUtnWDq8SkFOpAFTPcse/SZRWZm4TOEfiuwcDr3xkLqzVmQ5kFSv7jfMwz+uo
TEInV6G5eD+lCGHwpksg/S7+XNhoRPb4jWhi65F/DCUahAWWvZcmMItsRJlSw68U
Oi+GXnsCbt0Ie66/4vdyVXic8YpWRQX1dIl5UzAPp3DJtsAJrQ68WB5qoZ58FYNw
wlMSGA1Y4dUPHUO4KDYom9XMFCJDgAfcyWIeY4g3VDODaLUjpAptw0PvtZ2nvYJK
WLWhwBUM2DqsCyh8vOVRBfae/OK1/+xYtQrGH//J/xEAUULgqnqQmJwnaaaOVC6i
wCdszu6tSHNYukmICfseUyzalXOtgiAjSRVXKkRh8LcthmV4xITeG2ib6zRimjgy
HTIEYTtAgJ4QVKaZtzMAyZ+vKEUsWR+p/fXjmaeFzUf3L2E831XA7FmUXYvg+vbo
YllJKqdTN/qjhHMiDOsNO/G49EApPdxYXrnXQfWX9SA1YGL2IhMrEZY5hHqcCsz9
pvCxPWSDVkL4mmqT2csz/oCCuK8o5IAzq6VI5odtgT7Y/M63lcvXd+aSX3yTfnA4
A9vy23RKAbiYwe9TzS+TFhh0aJL5WulnAVmLQ/FWm/MzXNMnuzAsvmJZzTEw/TXV
LAMG4Chwuvp+JyD1ar+jh/rp5F4UEe1Fynmpj9rlPezr/8cLEAQJlQXR3DZISu9n
vOXzb/1nsLIgT84scAgUgNZ3HNEqXFligrjB5ZVGIGXDp5g/Jnv/0EKmFgXQhOAr
eBzgwQobpnfHn9tFj+dw6aXwII/7D8EFvT2MOgJpjakSg/8zcUaMX+hMCYXarTCn
jReh8gxqRfSddTAbXhdoIMqKnJQ53tTV+N6/h+d+yy+5nPS7SkeZaKCc+WsqiB/o
x6WYDH5mP5XzukTSEqfcSo0w8ihm5UA54B8DSss4844pgsE/7afAv3IOuZ0b2Ndr
P1sY9YsRAfLxhznyp7YFsjIdyDfq0eUb2fmmiCIM9DDtbb9nURaTvuEl+zpklJZx
9yqC3EG+2GCu+S+OFQsjNKKxY7UFQIYcO+pnbcdl547Mt8xQuaFht9gpJ5QGrIbc
5HpknOt4SSn5wl2O9LCZ9UZCaHFTDHU0jJBlZsTy/3k4s0BrpFP9WwiUaFldlR+S
ooIJf+Xpr9JQAmWcW117Ov0lWkXYa1Zs6Xualyb/TCLWeSqqr5ytIb+bEmxCg5WV
vHkbQMKmOj9UWjTqnU7v6Rzolg4UsxopNWdY7fER3hCgOit9NWVq6JJgsRwPNB9o
99kRYGF3zhbZ0225ATUcGzs7I5MGHeYcmGr4JEALmmNeTrD7lj+ASmOPmjlZ8+kM
/+hdunvvPdJVWtv0k6T8zyVC8p4ZqqwBEPFPtfhQVYCkQtNnOag18hP2f2rk/oU+
4yFfn4L0v9/WO7+hiojl7dSA+CbblSPz/7bBHZrDH0jXkAM5l0H8pGgMBnIbZbEI
PP9kBdhiA8nk/2DyYrGxLTG+4AFTcEuquqZfFFrAi67C8xMoqyYTM6EGpR74fbER
C5tI7WkypL46w3byEXDjG3WlngAbcxHjgFDgo8gxc5J38X3gjCWq7Wme6+L0KHVD
Vll/C6MXeRpqROynp7u+/qsijxMD2DgT8wwHR8IFDRnsIQiTvT+e3UBmSVeZKOAM
6TZpfjo2JCHORvG1XN9n7cOW6I96SjdQmwJXGUtN1IAjcB58o416fOmnaDYMNLDO
8LahX+W3wsvmtzQ/kLEadvfV/Ti+92C1QkMxnxZGzy2p1rcLbftIbqojEwDRHa0Q
CLx2gj+/NJ9Y6o96XeV6F7Gk9jr9gUn6292wAtJRNiKWojeon/Q6UlfINiaXdKqC
oGraveJTZqdMFdGZ4acOaQsuqWW9uHTeFAyKQKsUykc89bKzRfDB+XD8gOpkKt7G
TwC1mKpmolafP6uGQe7xXMz8gub6v0YHdDkG4OBtnqe1njVIdYHbLdlTbOhVMdO9
vufEMqd8Wgh5XOmVMLpr7ZkwMTRwkZMuX0mR8iuxTvLxM+57MUR/yftI+TQ4WxOP
DhexDebxJPBk8e7pgMZMJxDV0sK4OvjaeoIiiKp9UmLyRy/uduzpqILk7M54rTAu
4IaSK1kWDzqQznhRO3nd8EoL/oPFC3iiOthc5ECxE86zgtIILeFn2G3ZB1Vj+s+e
Y0CIaLezTqNX6shIkX++1LyAZ0EzjPIVdMbjxahE0j9TDOaf7Sk9Q/vGoIaQA5DK
ciODb6hALhOYAJf/bkG4UWWVJv2xnPFoTWpeQC8gEDUfauevqQSwjD4krwRnQQ4+
UiAD9UWESiyTDxlpbS0EVCxLgAGuVlQiZBzXEnySW4z+4WAJxn7VoRu012xcc11n
hQXYJ+Ci1AnjdIYVHzXViEm7pTLgpzWlupmL7rN1NKQiuWsqCBWLCq6iEtHa8dBa
CXJgiyG8JOXVJMgT/5EX8v1+FZnbxWBI8jFIOaNsAAq/RjRip8q+plWlEccXSSbD
uR+NAwXvzk2w7obI+u5dgC/rjh102dkQRDXkPAxpbWQiL+idV03GDlrMc+jq+2xf
99CVQRFuuP8lya2LyOmyCTeDudHN6FeDToH6C3xUvydvUpjIl2mydyMopQHI8Stw
XHWIe/hTdTbO+aip/uPr4q/QfDqJyjEoeKh9NAsBPwbUkZ/1nM8z2QpsgdmMnoRI
5WUpHJQX/ggmTGBg6P1E6DdC1PBcYPNGHsgIlCYnrKnre76Q1FpzSp+Qhrha/J+2
x7OuD7qEsRKcF3hZRk2uauDTI2Z9yd7z6/U1Ruz/j5Yiszqi0o/xGocGMox9twJr
aVWeCYWUUuJBYJ66LXMI/6dTZDzW7+xmAwe4IYjIdvFQ+fvi6v5LKE+vJU/bbzGk
ZH07Z2eA+fSOqkD1LpTSuyjNiGFLAFm/OWJEwjOnZJAmLa3vrt+y8FhLWtxDxW6e
7dhWCNV9hPMVpN8+vBOAfomz+P6YAjQotEe11AblfPcwt5Q33n5axDwYjooXea98
wngon5R/AJlg7uQ70iPYmJ7s/XUFGF6HwuX12tzjJMEUqDOwuQl4vnu3B3/oEbvx
oaUF510tvqnafyM+EP4cG4nc//YhuMCPJ1KNDiYNannmPEE2C/K58ATEOpf6dw/n
ODSQtAaIGbEyCJM0SFXkQ2+csrp9lWLwfRK3GQclHIYoEryb7dw5/UIDF2sgju6a
VuMf/lmwHWX/b1lzftqmnu6rGqj9d3WzzSfDdYYI443lK3kXDG7pNCPSRigorozU
7B14xTnnb/Z2OqCDMse+cGXoKd7NjXnV4tJkiNQ/Lfoub9wXgCOrqB3eaGYXftFm
68bkkOPE6v6OAvth7T+ygN5u8ari3jhw5576KE8JDgIlxE35sclPCHWFuqfn/nRq
BAnWWRkUZfeRnLM0NeMtVdFyphz1ljK+N/2DTSHeX78R/XOe9fmjthVViuVp+uFD
KqqAbTqGETO6tR7Fq1p+WwZFJglMNTRhbHqOvaQgihCJoXFicmfOqeHeh7/mu+wt
eRvRxsZ2/P9fMIqmTtlTpMgC4YAobbECGtRr2YSceTeQZWMtTohT5l83mJqqrQ0o
G5XYDtLjLT/40e1uyKdrIuK0LB8gjw0tMeORWR3W5mQcyVBNVs11q0CFPX0HkI5x
SN+/TPaer2XSfqCllmzrQx1/IrMe5U3OtI/A5DyQyMOrFGOPLABYNGLgVCBm4STi
8SiOti3ZSHrhWjJjYF6eIAeSFffddjcZYXuRNCKrWm2NsGbpi/McRmfbFypD9tiW
PYH86BAohO8luw1j/je9MlotSVrKOxLcU5+ce7jGT42c0PdirL8+q7p1nGlUfdOd
gjPSKRLXyH2cLAGWGc1gZ2qZ/9wI7dudcJfXfNHJdeSbkkYe7ZB9O5GLfPIbO+SG
2HkgXJ5bz0wrA3hDl8k0Ic2K8imRBrgZ7hLprhwuEJRsIX33EQ5HFILjEp4AILR5
9i04W2BmQRguwFwbIADUsi1T0ug0QTK7EosrblYoa5/uSiMD+1G4pPrDwD2qfZiy
vdwtA2kzjeBIWV5mNe1f9wstRG+TXDTYZkX6gDxrnKPp4vJybpD/cCBdNS2qHmBc
n9/E+Vl4177lgWv5hWx5yNvHxGdBiyaKLGRAMrYVayoZS4iRleerXzElL79qQUzw
m/QsIjBdBDlOmKkfTNqPsQJbrI51zy+iva9gU6OZF1+7YnsdRp37OaI7ULHqfLRQ
VOCdYGon2C+NDOr9Ii0nDcrtujFz/CiX2MVvwzoW5gH+6ktUvWI+JDMlKJflImE7
/v4QAmI2dQUe9Y+TJwagHtec1evbM8P/VsxUKdjc6o4dLNzg7TypRidOpv1D7O3U
LfqK3xpI6qtbxIzn2dCRXwvJrG7MPPHJOOA+4jQobecraYfg8M+mgTiJItqMx5Tb
aM/gJZevrj8k5KXK58ROlphUvubDsqOEiQuOLFAjpffCUTJyIprAPcOzB4ss6sZw
q+y3T1VA18onbgrSHxRPmzP74R5JLMwU4+w/U9UMF6r1tCelyidZ+X5aVIrghJ/2
AzAmK6lc5qJNdbxQT7QUecYzv4p17Hehh27P6R8aoVhRD1H/e1SKV5E9G1RVsgKH
NaVG7FbFZFqrr4F2qV1/Syy95r5STKjy8qByHVjnqz4nd8fijjuvFBJVkhi3hfHJ
qXqQG3c0CxoLJAjAOABz7n0lQAou4g3uh7kVXlK3x4ONuvbx7sDHYqi2sM/IVcG8
pgFu1XRxzABGPoOKOLROzof5Atg8R/06tZuIndrla3Fq/jqKNZKa8bWEUV/6g0YO
6i7TBU7jznqkxHkoXaK8rf5NN52/h6Ao7zU6Hj8+OsaZjr9Dcx2ULXTt4vKc5Uxo
lpizdGk4fs/nwk/KoasHSwSDcUyb/qHoda0xBgpFmW8rtRukkNVGs1fJ1AsP62Hg
kuz8CoG9L8OtZ4wniu5QrUJ8IwYPKLeMB5AKDYiB+3ykYF09sfcBnnjJ3M8/tHNc
JBZOsLJrJRPiohIvaXmFBeBRnqVsMf2lQ+yhF4huHEZD5KXaMoSyEfLzv6+DdLp0
Hr5YtGJoBwaaB+9vftWBHaRnfIJ/XOyijgVFy9Xqr5t5ZkhfercshOIi+87o9bGP
sHyT3zJrtDpegJRNXaYFJVSPJHQPTG1c/Hgs3mqOPS/SuJDTeoRDtGBUmCcFYHIe
PaVOc5MA2pZUtXi/RkStyjs5ZQNOiCzfGE6MNcq367ZQasmucuUAOlPLRgDeyu8g
fbrcqsPlqxuOLP2v1AWs2SUqAaS/JcytRykwQKrDwr9L1DbLvsGRClZdIsVIaK+z
692Qk1Wqu6w4vos7AzA2oe4QTxXdm8MnU2vj+eKyjDDUrZdaaIGhO1M3EW/Jz6eu
9BtgQDZ9heheE/jUQzzAPSIKLP6xtFNEFgdhVfXpYQEomWrNzZBnG5wdpei3yyq3
EEaU26LoY2AlaozjVUh9rAbMKgBFKr+p9DJEBXmlRLr9pvx7W1yy5xZQ3kEkynj7
X0QTGwJcNA9Wt7cny+6dqBtUwVeO7/lGeGhXLt2Px7C6Llnx9oLcOuU+RRqdCeKc
aw7mW2yboxmtdRbbe5oIJOlxA2j47lhw/Eo+M0wR91GYKZ9N72ORwCRLsF48Mmd6
CgfiSF6+0ZCjlttyIWaM1sYG9ZdxZ9kHq6IUD20hy0BMZ2jDlxkImH9pcE7VENdq
gZqg5YuBSQa/c9LxeB9b3zORL7BBySTFNbqJiwGHG8AzdawHQmalpS2Euk6HgHyM
cSBSBTZ4p1O+Vjkhq7yrg/42Ywm54OVtQMRrZ0PO+6qpGrUhrDBwOQjayFgifDDT
L64jKzlYWGXDglNwEaBOVu/3DWFThK24OVamT74qjtG0oe9WpZQCc1Rx+3fOXiIZ
BeU4iTbaSy+bLiH3xEeEtVNMp4/wYhKCG0dPBiYtWPg+ypmoZS7YNV+c+wuycXSY
TlD66iGFrdfmvRN1yc9XAXhGrrlxc9Ks9mU6+LH8grxXAP2RzqNiq3wfQLrrq64i
J1L3mR7iAkgIbHYGxIpcNtrhe2/b01eTcovESDqkIrzHhyNpfY/5+Y3hnS8NET9I
eqc8q520klO6Rc+y4+0UFvxDnz/wL5ExzWg6lgkFyj/bidiGzDXTAPLSotQGx9/e
mvUPBgNhiFGKq6FKDQkLlYyFlI/yPztVB9YPIOXaHV7wuYs9cTgMOMV5x3KQMYnq
y/tjr3+Af/aHupv84KAteZlwM5A0LiUJx+4Qz5bmpikRzF2mkOyVC5mLLXSBHuPR
xndcaq0pH03hScQOtruYE13y9oNl6PdydDbLs0AMo38ZDaH4iYdQK5lQKvpWFTKm
5rlRzzq1aOu7OXo3u3MsJmHjeSkC70miYqU8AWZr2rlMT70qZrCQqsXhiXFRcAQ7
aF+jsI9oaO4B2IvBFqmtLrt2Bz3QVL6JafuBdlxgQg2xK7TC67OaxlHesoh9f7hw
0kpMhvLo6yBJAwmJsiQVCLMEkpjCjby+6jjk6R5QP1bmZxE6lAIO24zh80xXyFK+
YoHHM0H0QlQ/LsZXSqjcJ7LQt5JIBhvhhPaFtDSQEMmeL+fh8zl2Z3WZ4Ro64ot+
uBb+gTW6iheI7gC3A+kq/vpwsOAbv93ACdqrU4lsfQiWoJvNqyjt7+hUZFq+xdKY
wfbgI+F49cZkpH2j40i95Wcdnf1RyEoNOMCMdtIu/Y4r4uPX8Kxz2ya3h8lMTTlT
dC2Jg688PjJyR7oZ3Aspr09xHr5kfnBXmo2lot0HFkx+HIuE26juby91wAkOKd7R
FDh2BDxi0vgvrzc0sL2/tYOuSjln1VPRqkyx4+azLYew0YuY4Q4cEOE3ichjRD86
cWMdGSd7/K/Xewseul6AStSTyrwAzM4i057RHfAabzeVBZo0smFe904bDE26kVR9
78YXvVrBCCFRtmMCrjK4Nex34L2zAH6S72jCyckI8ay2AiK5pCKs5wVEkaz1+25Z
Tz7J6caib1V9139MgqxRr/fp+TP9MW1XiS7Z9Au85nzyMeHjOYDqWrcO7Lc28Q3r
h53Nq4+lBfzDJWWga6xcMgpYhcRbWIeApCwtnyo+5bZGQU/hyOHmHgd5mfBne2xl
RylzXnxhBDC1AmZqaGEFrpKl+yDFuCx6H44iY60Nto9YUgllUu3d/LYbrGGb8knf
BIMxGHFOI7NIbgNsN/TSyGQ4ts1WT8WhX9fYwLgTOXBQbAgU6xmuGiJLdEgZ0vIF
s6DMibGts+DO09UcJz+leXdmiYdLywxIFyEZjKbEU3MzeNmIstoYe6MaHbk5v0oz
oVF3ZdBgK0+USa72rOwGPdfOb1Dp0IUB+B0/668FbNS449LyXSrKYX+1PNF8X9pT
oa+jeF+IjuPP8dgANu/hzsle8qYxaG1J2L/NaabPYyxuCWK3+gCGUNn90SKa2kkQ
bsBkPxiFQqiMqU2jKdmhe4fFBBJ8Tt0q1vGiXwuKB941Wip9/cSlmsoOUvzSw4iO
1hKeno7kADX2ts3rHqXHspqWNd5hCnTthaoAU5I3LEojaN3DlJhlj6/gXdsiGfNH
VTz8jlTjzD38aBILv5ibPNiSaDIbLuEVvwTtfodPVM5tB7sR6DOqhmvgLwX19eP9
vOZlUZOopj39J3jlFrNuudUYNwTrj1jNj4LPrxv9LWyr6APXz7gf2cO/wL4NiHzk
RiVab/+hPPVT8ioG1fqq/UV4yyK34gfEhkxqlUegrZSW8FA4q4XofX9VGQuCACQX
a3PxJ608+an1eJO5vZ3EAwJhcuC2zbnVjz4IHI1BfHHMlo9g2XyJUdeM4yq1+NLm
6cWg4HjMn5Jvlo+079bHijdCLKmaNsqF43BWpQL+RRagwV8YWX03wWhBt6L5Wy6a
NN7z7SJDFkIByDSNel/hYLmvZARyyjRq7ab4S9waNnt9ZQUWbQmL9EnARFnW59Fk
eTtgtiq/cyCJIATLx/PInaBg4X8EtHP2qUhwoaCjavYU49rZpWDDNXGoy18A0Eg9
YFnTtC0rPJ/zu+LZfnY3/a8uhF/j5Mit49b6e5MOqOXcgr+pEkih06WIvO3Y9Uwg
YB3JW8iD2R/In3clKBBR6CeinsiS5T24RrU2OOD1N/W79lK0Pe3d5xJ0SORHnYAm
+05Md9ZPZlp0OfMk5RJVcQ1jnvVOMXB0esO654RfI/b2kxKwy6IoCTEMv+ITgTZi
d9NIQrn+ILL+HuTFs9JwK1sd6zSZ5WNrCtsjn6h9F0XZsnuPq1kz70JWjA/vfh0T
4Wi2Y06js/2mNfeyUXw2mcCptnwPHp0l+fMB+ju1RqQk/FtT5JKEps4prBTSkgm/
XrvFh2876K0ZRgaKxaEOJp4XFcpk55Wz45JLN+EiExdM9CQC2mzOVeC848YGI6q3
9gl6K/HfbRsA0Lpk8Xak1MIp/PvhSexAeUineagwyThwaJPyJ87MucDoMjQggnPC
H+Kh9CqY9sRlVuDcQ5aBx7y6HbyxUo3cbomjTJkDc7Sw/khfKHdr1OCez096TdED
/74HkDuZ9FDXj5jUXvyQJcdQkjxRKElyC9GYmdb4o4jW1Aa0zKeYjIDRDCgYqHZl
9frn3NbGd+kugGH0je1ownGqVGXeIf7DLIhg/4H/ryAdld1koMv2H+RQ71u3TqDa
Kdy7B5UAvbnN4b9Yxl5/N2wlUqLyvB8gZrnGxL5c/ADH+l13a6SzmQBgBa4Iyb6g
Wy9M8NpBPZUyrHoeYpQv5WTN7DcMDbOXag0YZ4sVc54NcMuTLlPt85LT6jretwz4
pLaUbb/GTFiOMtq9NI9re7EjtOzKXKmWC3OvzDO0i7Pggs8MijeXpYe/2/cWfyvO
N9zKTqor1GKP9p+ZQu/RucuD4kKlXV3v45huP9z6N8SBgpv0F531WEcdqzgCyb8H
wrF2AIpz9fbvBDxKoubd6n27CuNdDRxEd/wfq5ZYbNyK2y66cKUVhkbHS+g4Evuu
mPWFTXYF4gdQzu3yNBwt1ZtRtPiQVt16wR/ujEwNZHIEPsCvCsIcz0gCa5ubjM/6
Qj1DWmuJmzC7tBn9XrSgMix1k0E7QrEi5nR3RsOyG0JTgmuAb+pe43ecZJuwAj/H
hnSy86cFh9/hzMNXYYrQDpZOXBQh5v3TU5EcazNxtbqYYxxNDZkXQ+QvGxgg/C9o
LrM5bsFSxEGyoT/qyybz4dfTUCz30IhrVYxXAxX2pLuipH69mTlLuBVe7Kk/Y8IL
h9p805HBCU7KIGZ8cSZnBwjUyawaMuiRgVsQYy3oBFRuNckKS7YSTzONLRPe23XA
rMySaHwMEbdWbiUb4JxNWldbl9sGRq3Xe9wQxYc84J7NmDqnz99Pyu6CYF8xa/kc
KdLu5KnCwksTATzbdq94TtkL7bVVF0c67zEh0+AwW4DzXmvb6Vu95xoJOX6vcpph
MEnqnsRORr8K/PrqGBgjTIssOv4203mJVGjGn30Pn+PL9QfdICIuU6J52+6xc53g
gmWpmO5cM892NT9cZh0lr9twZupsFw/k9P7tq7MzjLoUoyyUWHhPccCRg4tl/E3f
3L613cLucINkHqEIQUDQGwD8I6f5LV6tGubePRH9lWFgzLVEHKRb490KsJz4vraU
k9HwbMTQpY/fIT7jjQ4v5P/A7bxHeVp90HU/xWPdWKZHLqNHHNdUsMNUl4O6BcL8
9CxRDsDtJxjRZn6ROv2NsbDl1wjb7qTEYFruxOYGx8xpoCYmYm/cIEnoZ0oNSOh2
B1hRLyT/pgcbdneeh7RwJimE4iv7XLU0FiGG63zz/GGuaYkVmZNxn+0G1kl2fulV
rVvvi/V3qPHfHN/3KUWbSkI5MQ6r5XODHl6TlrreinfmoWcGV9SpW1ks+3jvmEHk
ITtuF5l0+w/zSGtAAfySNjajP8BzxnyfXfpaFEhfhpe0QXexx/Y0wip/hLzbGT9M
BekkzUUfHYnypinq+34GpcfnW5Q+6G5NgvEY7KcWGf7g7G2XJohY7nkLetEEm69s
hP2Dd0uqpF7LEvyJ83cW9KqrTs5hlNe847j42DyoFEN/jOD1SpYkNnk7TbnwlR/u
tCvfVH17IGS+TlZF2+2lkpyYhhkoXsInresCakPPAN/L4NZaT3ISwa+TyYigrCZo
aqogdv533XG9TRiXfbbCsPKXkTJRDzeifdZAvDF85LUW3WqniCe/D2TLOD9NNBUI
utDP9Q+pmi2OBiM5eiYALW2neBKMxT4ENKPsGMcoUVan6sIk1npbnFkYLgXC4C7K
Ca+lXhklHLb0HdWDaEyySTVlo5PBqH9VhgrIeGrIWYvwnVbigs9eKmKjtdWLpkXo
y4gH3zZxLOzfJBn1fV50/knXwZXX1R9qQF6BgFOXIdGXz5bm/5YMin39ogbbyv86
KhVAQn/p/+G6vX4HP/FT013A/Jxg1dXKu3Ll2o+cTJaKDGgS/7u62HtwS7D7Jsee
+7i9lYWv2z+UJcqAjTu1p5pKt4I9PNFpLab95hwKWLCOVD6fKQUQdsbCgz6jWQHb
bHIAeLM+K7iM949TdLHLBr8bsgokfzn1zRrLShpx5yhmnRUFC8ijhOwzcc5vtxYl
pYClRCQW5QQEkLN3+8E2MCrJ3pm5LbD2zKeL4REJ+VWOcNVJGU1KWsSj7IaedPM9
1775SJl/h1fjnWCV+BXsCxQBH5O+KC+aqYriqYBG2yhN2Y+kBOlvN8TKqfDJBQcM
D45taa3w8/iyQ1ImZB6fHyAwPzpDpKHdG0mO5Z7hfoEcGtYQVd5FJuxHK25TKNTu
tATiACdy5T/PIlkS6Y7j2y9aMY481+KgWQFSSnXCb6ERzIOIwdQsV0AVhna9ep/Z
y7+K4MYtZ5GRhi8iPmbeuba8XS9p2oP02eQ3BkglHloa+1aJUfsl1AiQvulnnuds
musRQPLLg1tTMgzS1R4hoNAK8R/Rgoo2OMdqbi58ucI6wcKZrFzKA00jZdI4KzSL
deqb78EwY1U0KFGvVkKoIWergznK6sFWvDCXtMjNz3FxsF2jtsDDNgCueLhgNOJM
w1O30kCeBvu6v/Zt0ezds9czAAak5ART7QaTRy7eMvPEJpG3ca1GCjYPRml8TBXB
WILCV4pH9QNKE8yvB3q5i+++kCZnv7f2TY0cca9DYNgZNLapxW4l0O7/eVdM86eP
GsNigauadyOPjtr2OJTby1NzX7uj41z2Rv0H26RDbMTshEPmeZ6DneBT04VvI/eE
ELl08+mPqrjWZIAIHzABfhxUXIQf7OIiJRtwnVPcJXg2+rJxItmtGvYlfyieo0SP
uaQfzJJ6fP/xhN54TsZy8KmMMcbZTg/qbBQD8FbY8031UOnH8/md1POFsPqrMaMy
rhJjSQPSMF1Gy5xMGkqOXyyo0eI2MzCvTa+Nme1XtsdDx1ycBDKk3QT4kztgVR54
UwGSZroGN3N+e+bO2CHH21AIwr+g+PPmr2QY6yqaso7mXCB/SeeTLR6pUzfUVPY2
BYkuooml3xL9MauV/Ctwfd+dUGnrMeBJr4YjX8ojYKocoq+UlgTmNUy0lb/25Caf
2GTk13Zt1Uu+uUhasgur3CK/f53PgOf+wr9dXh8WVYSOV+lpwSjmm6l6aZYsbZBO
4nED1kCdOmdQOn+UnBlRbUrcXbO074YcTVor8/Y8a8EH3dMN5nZmdjHhvYzX0EQ4
5yg0CGaxhKhvEf4m9DvDEGMfQhXtybLfIX29JTraF7nLphFXijhMIW4t3mi74G3m
VK5ICSI9TFUD1QqjrUsDZLD7SMdCGNGQ8+7OquvRvZxVFGhBDzEr8+trkG4tP366
buFxHVP/8fsuM03uwFU82TinOomtAXSKacsVd1jW7/Ml6O+4/4LCtZLEpGy5rhO2
wvv9SkyjUSVDGUnXMmU1bMECznAcWDdyUJB4oUg0lnBcI0qLjYSFjK5zBujwXzQ5
QGrcBGfwUv/smtglM6dtYRsXY3g7A3XsLvlpogw3ZxoFBOt+bgU2vGqK+nZGwyxy
989nHtVFSlfbl1Om3LoBl5SrEv+Sni2ghgpgdosyCD6n/WIcx+IpHTkf6cycObcN
Aq/7iHP+LFvNWlmvQ7n69mOOnIIkTar2sELfyTBLFAvTAkYZ6i3SdkQPQsYEHBGz
fvcXnXiX1Oj2s71ZfbUhJH9Hl75tjlbW19GFr3o5qE1Vs50PkV2X9sH4HtdQI9OW
w4VtSIqThNWJ/PdhtQsExCHzoSBftM+6DJgVyZeh3jlEpxfknzW6WlEX8UldNglc
8LaUB4X+ULgNJdKnI4FrEIJD5yp+NidbnAjAQZD0qJIZq8k74XUBmwCBbAC/Yccm
D0QsQUWpa5jWztWOMRPJVMi36nbvSJGboOO/CHIfafLOhmi29RcTl2kCBbg1BBYO
AMNKS9jRd6GsesMAUikJaHHAzmA32VJQLc5qCoFb46OGW3SntgqJLOJ5w5x4sKNv
ohbN3mOBDE2Lt6SWbRig50BFoAeY/rGKpQkTSYqE4F3pfxB+S5Aq4P0ns4y5xcou
NergALGhEXXy/IBwQq00YshJfli6H+mJkk/X/Kpx83FMJ7bdhDjCRUoAgmcIgZPy
oy/sZtu/cQg5Q5QvFi30xPOdc9ZEPgMjk7J6Wf9iybTQqnKEvnMrbVlseqDs+o4O
ZAVjLblf+FBgDG3kvJQsEZOKDbPfLveNAv1g87IzMSs69mVZpbfmfXNgEOudJklh
oDtNvBTxey03MEc0kRwn9v3+oWg2p6Jvi+NAs3z+/RuLIc/h+0t3lmv1FYm+WYTX
7/AYXoKd8EfuEtCC4xKV53kExl1UhkeM21YswBTEPkxcyyw8ePGYBH51OBK9pA80
6jm4JazRCBSDlzOC/kvSREbkY+tQgtXMmRi/TdTyyYBveOCdE4hThUNkov912AV2
Lx1OfIfH9ch35R6B6mbn0eX4xHxQBTjEI6ZNbxwpOQatmL5OFDiwV5CBRjGjKPCq
9yK5R7zY1gc9w6CoN2OWNQTeErdhEuNU5GF5gJ6OAKCHb9TyeJTZxJthNOsHSk+T
TK2YbMMODvu6UlIZyaO/OuaaXP5Nq4MriK0y14Paaz3SVkd/NFwImhsbDAtEjw+i
u+jOdrBBDYzkmYLr3Ic9C/GfpXozadqVaqUKMXJSTxS+aajXL+/vQC4jS2c7zLq+
L9EgqGvNitSgv27HB+QvelkBwupidso+K/0gAJEvEzNwsPEev3fUZo3fQEqbmw/D
iK5hP/CadvQiAcMKvjzTC1CbEE93ExAXr/zsUNJgamafDRrvwlc0MgfT8uwcDZHZ
xiTHqkrr33aGQ2vrjk0BIiLCvmlP28/15G6zYQ+Qy3KrGCkt36dcoQvX/pWKCjns
P9B90hnXstZcmdIhnMDCHKEKJtKRybGe8jn4z+Ru5zBm9yjrs0R4Hw5YLENH7QCP
7NYWObP+P0xKsxfFN3hqMIuTZaZnJZ3kpOFxw7hg80TNff3Sb8E37YkrJFfRjhO7
45VOU17t7qkqsAedGptqGcdZKXwoZ3sLbagb4wGarchSiJwsxlbs7V19m4Vlvg36
BBancyDSn9jFY1tlKdliQxgpgcv5xqf3Vk0zFdUV4KcAa2bChVb/uCDZJo08R0Tq
mkRJgQ5mx7oXh9tNMjISaciMDiksVhSjBFZMf3VoJP6wkbp8MJ8Gbr5k+MXjZxcy
W4WzoRD4R7yuYTVzBflgaAzAVH6+wrgpGTp8xuXI3ZkJSll8FHoDedN3yMny94BP
/u1jpyduXoFmDh6cuDtBDm+QcYAdLGhUKgEwvhK8MxbOlak1gAXgL/yehBL06/lI
wZdbP9l77tM1xooUtqYgRfp7/KE3aUfWXwLV1Z9EevbFVQLlK9yisvt+wtIwVSpD
peMKJ/h+PUnUSCDeMeD2eI2Hvd2ZIilzGScNxdGwbiDdCeIiz+a07BFxxCHgT2u4
xmc7EAKwJ0Agnp/75IUqgvBUhs9CPJ8v3mlJT/05b5508kEEHt24Ha8IgfT/Jy2u
wEsHDRjINL/cNDOX8VujE7TSAEHHd40yUL/vBaaCotXr/5Y7cO35cOyg3ZK1Geg+
5Bj6rhO+g7xCFZuInDca6CCkN7OlbvvThM8wwq7V5DR9/RaxwLKkkyWS2jfd9W/r
/T2HIUW4gKikSgZy8f4M+qFlaS3Wo+KoU5y0r43USzw/bWP2JULtL3Fg2I6/3mwM
kO6oX9KEdUMyqeiD4RrzT2ErqjTM5cPi8aa6OGufQ8e92QaZLITiOiNbqxeU2pnP
CG2VFmNQ9cVJGToM6Mgjy3m6wsG9Au/cUGsGUN0GcIBjdTl/5hrr7Nv4BLJFNmjX
pnkoXkdkVzgsHSQooln+7AzlsuH6RwVwX8IxZeKunQSp+CgRwWZ0lUvTTjU7k62r
xRYcq9UwodtIlxF1z6GIdiig4Ee6zFVVXEvvpaNJPTOPNZ4RsrAe/oWtvvmMIbWn
2eddxwJ1jQHYYHWFuyINy62+xQuv7FcNujXVSLAoe2gh7FDdptD9KKbudiDbac0i
pwliKRRVXgX/jLATOlzZf2TuGrL/fYDiRhOB+hS+jeNNeOZlRoH09sXZkxMC36jU
LGiQ4tJqPN/gcqdF3JBopDFBSq+nUA2IYQSOrkZp1q9ZnwF3DrEQmqmXKrcT9o8F
9BMrxLyk/B7hE2cBdq5JPlqmUjXN5uyQGg1dFDpL25BPKmLkCPas+ANgqALuWDTB
otDGNxnzuoz0INUJDKG6P/uqPKa+1EK1rwr14L+mmyglauKFsPSLdOwNtnS6LJc0
OUyYN9Dfu1JgusBHRi3+bw05jQ3BKGWoPZ81edP7mlxDdU14hrEgZtqWvXkChz3E
XBxq7bDer0ZBEp3hLS6kBcZXTdSzwnK3WdW9rgHZetqRoXVHWuSuBV47RFjybRH+
zrTHE3X74bJjwa0pHe5951NWykmQ+85iTkK7UaFhpAPSP8egAlFHU/FS73wNPOgG
/A7Q4PPWYT5dqW5g6HqyCIfglLRFZULEJDEWJMPWBvfJK7YQQk6pKpispJduwdCk
PjQl6wo8FcqMJnqicpBf7YDeGxMIGzPNo4jsaVFtLKyA3z5i1Hn/vE/jhm7H4JLu
lq2VX6lGHXoV2jKi2cnki/QesODBATn4NPB7iu6dyh9kxmy7iNasN8+8jY8TCZvm
AMLgkMViODji0B+VEAaMOfAD2nVhiAhOZtd1tVI8acK94oP+VPc2uNnhtSwCZGlP
gOJFjtJ4KaEv1ZMsdMv0Jn46waNFZC9inwent6gCj64EtICAP6ibdNkkxhlPs04N
f92h4YA3Xfw5ocvSKrvMgFlgVGoSW7hJ1k/UcOamrCR6Qgl6obITvRNjUSvngnEx
S4sY29fD1y6fbc7DcTT8mjk7SJBa3hKsipDzZ/ca4Q/aMzs/mao3KQUw9PGYFmdq
+A+X9MkBYpKtf0+UIXas1WuWe52tdXlL8PwSMdueenpnjyjRQMTPmwrLyTq+BTYZ
RHbOVaLF1HV5M8wuLLYOVVwIwSCTFK3ELcrhEywKnFK7j+qMWNY3dXVCvAHAVGJP
9u3K4cvWaak+c8uqSnc9X6SumYHbDW5uck16w/GxBPbA61PxwDt3ua8LgwJkV1bI
3mmW+vv+YxcUz+Z1ufVhwQvM0ZI8d68XQ40QpMxoyht3QXxijv2STDp48k8VIEkn
CncYYnT2mDMGfDgxS+KrSDuUAQZgoYygbo1Ia7+pmBpJL1AAdFqvkciiAskch0fb
DN1yday6yUL36e43w8ssGmJzLRN+dV87ELCsatcLdmFJGiraDGoLXZMvL/YAkWI8
IICX6LAeQUFN15Dgojr452f/lrJoh6sq0EUf9alhILeaJk1WF6jYCjpVMvUbuqgU
/yrdTSMUEH26oZtMh5lVkiRbZv63K9Qs7V6chErF0r7BJz5zLQ9pmWtYKJo5dD4q
3tBslDXpfZHj5hMgLa+ZWCvphSmkyj+ZF1bfck3BJOB8ql8s0FQnoYycyTLwExl9
jBX7n8PLvNI+3H13XNKUOxavgPoY14dQWwwVN2p2h+SnE3JB+6K5GrdreFK0ujZd
Wm/fA53dCldc2DrPZsNw+gY8b0XtRjkxs2k+4WsHE9/OqY0Y1lS8FLbIez1BuADC
iSAhK8mI0RPKU0Nme7K1twKXLrWsbpx9A8KnP91dCIL0OcdK5DBNpdDiQnjkvITu
/VtDFCuC7hd6/Yh4RKKRmkTq8SwUecd3vIbHAUx2YQ+L5+eDSfe/+bPH9R4jCa5C
fbURtfYbAdVPnylR3GBHNueFeGxEo4n4uVXStEmIx83AV6q59PwU5voEHzB9ISvL
VrJTEFgDtyTUSxtzSfWI7flVhzZpO1TRfLmNgU30GfbplpjmvGMCDcqoSQQHFDXH
gckz3dewGcSckXX7PUbzeMeLLmD534+ounzIRhiw9nWsrqUjA+9bDjmD9bYKyr3v
gqIPyigjL4M9jPp6hOFaxYO5LCql9xWcmvJ3i1cR/lMHThfMwBeA2qMI2Um0krUS
m6t17X2nvaqBXzaUmZp1RcLh+WEu7fcN3Er4b/jGObqbbJ77zK5ZdxH527kzZ/BC
xgJVbHJiz+47vaWSDxDGpgo1g9wvL7ver0TI+B2/BfqVhsJVZPdRUrOUHGq/+Myy
g6RePcQzDhXRgQ6T5NxamDVI8fwkbZmSkPS5MN8sH/qhxGnsjIukJQtMImW5CyYe
/uWW5on7BBFzQOwwu8qEsB3sj+jk9NyDnbKE6PrLgR3ZOyZKI/Yds+qUSYMXmu8U
zDKOBKB+XtaZDRL2xJZMFliXNp55WX5A+qWyrlrZTHL+GLgz0mmWIQuNPzuVpK4t
h4fDj7mrCwsWeJcPCxPi7TAJcMl0m4o2z0XFCH6X27YuKXOU8WXGi4Ynu9STxTad
wvlbO/O0HscSUcdZuJZOt9gROGGi9T+500AUqbb4T98avcHdmOzeKLNo03jMTy3Q
mriulePBlgWOyctaspJHkLXzDM8IYD6TEcCykFRx/XMOTQZEItNBqK+Zv0W6XXjh
UGaU8xz8QdELUfXJOVsjtWdKMKUijgG6hOHu+lCiX6r/xHlyFbN30JTyXJXqg7Eo
2R/fT7y7w8ViOhHSQ7E7a4blLJrqiMqcUSKXnnfQYrnWAPsw88UQZ+S/vrsmObOb
+8yyzfAS2dT4gC7kzwKrFcQLZ7kyljZDSgdD6J1Nhx1BBfWW3kTA4OnFwdd/DBIy
ju99XWR5H2SOtaEFbNB5gZLJZ2IoKaWmF+XjCh6E5e7rw+Lvy/qKuux+Lp1jxyBk
U0YthzxogBW4A/711CmBgDPxMQhq+MlCqXSpML1d1z+2raFnj69t4YL2fXbGxiI6
AcIf8q0/s5hdfX7sLtD6JLfA/nEsJKuRIhwNs3zqHMmhMzKmwvvvXqF/gXgBWwtW
BfT1ZBeS2/IwsSViVM1NNxPGgL53T8f8GOWFeZ09beGWC3bV64FODOwzQN7RDgeV
ORv7ndTbVaG8ckJRvaYBt0poP22ri6VloQcDW7aJo+NUjI3aU9VdHJoalB5HruZl
VcZLe7aC31Rg8ZGlSAysFPjii7Ty8PkoRiy1ZVjmMTmnj9VjNPFWXM7MqQcINbaU
VPBt7S3tvmZmDDS28YCJZnjCDBSUtNp9JqkuvwS7+DyiJTBC1d+PqrF4sm1Ffm5k
X9Iq0+OQbWY0B6ozGIsPxiZpT7Wg0ytvi3T4mlPxyhVxkpAHI//Q0N+Yj5LvkQix
w/c69YJ1mqgKWZfMaKxS1q0b6WyOvUVtmmjeXI64cg8dP5J1thfSimnKwfUVmob3
4985diWLNBA0aBrbjCP7J9Y0arQPOCdBd+5UHb0YoKzXCU0SnmfbiJi6pxI9QzZw
oDifw8BWRSSMho8O2a0+wibQako6y4LA2oBZh/rhXZpyBKxLhJO5nzPn7U4Q10iK
9r6HEi3Vafroe8uR0goh/SwW4EJ59oIH1IMFmfCu2w7vjfQqRKpPtmtFus45JXce
OQxrmUq2RmggXzBbfLNmKDcKey2O0A2kPQakjFJWDFgwZb/0pcdqo1p0cocPfGbf
XixumySQ3gDz/ZWbuzzP4lPjB/PlmGBZq7jD7sXro/kDlg6lLEPstbiHNqupiY/Z
ute/MMiEPeLpok5FBosclAxjUyDiyAVP7hHVTUksoJ/Szos2gSQLyUVO+DQVDkc1
PjmSlVV14CuknkiOPovq497ouA5i5t1Dllh/6xhYC0nseiPrt4+ADc7y8etaLEdc
QB4e7wRqDGE/9zVA69uVN93r29hTKULbjTT+xWDpI5kSHSfvN+p8WgixteTPMUom
NX4E0Vr9XWnYjHpLI+/PZO1gNgL4dhBR3N8b2IdIKybr7FfVuYpNhrQl8h1yA3yF
ZIbgbt9SVT1EezstBklSwTTSFvLeuSCogXtcYdARsaCfL1Z6mm05RyL/SWoxWj9o
48hXS9Mpvbg0EGteAV7ZLu7RlTeU2CT55CL10H9mXWbQh3DhtREfweaOLar2DABW
j7HZceqKAf39zFhQSeDAcyWa6MFIRMyj0kMZIbZootgkELcKDTtN65H9843oHNnv
96jjNJRc3V/8CcblsM/hO6eTEWRkAX2CXjc68ASMmKJcZSpu5VxJIGt62qf+IQjT
fpurEphGQ+i141AJCNAG5kmqRO8D82MPuAVWP+XCeZRxLPuk6jWCNxv63J5QuT0d
LubzQ9RhLSDy2jBnvNGZqekHsw2A5ZY2WwFm5q2RlAPpZxHHFHXz6ODv1FqIDi+g
b76Msnq2cPFcNPkHmsoR5fe+fx3DoApNXCO/WwLeOIn2jeU+RJuUwzEmgO75YOMC
PlcIU+KEq2ZZpkcJWdgiUsJhYHdyoYytwhERdLEn0GRXEKatyba8BR4KFamRNoRY
s0HrsQ+HIQI+0IN0u6E9bow/Znc3zhdEpwSzS893UZVeHE6v0K2vO3CWwL8yJOQY
seYuCvr2b+LbAgvjdZA6ym8ZEwM1/0swbK2W+k0Pt76cWIQECCZEo4PF9gbpHCbV
4rTG55+0MZvGRTCUShCcrDcCp5bjl5aEjhCJrmNW9y/OeF7795elIkOXjBjyUnKR
qMzyftwg38Ytc5tBZKb3LU9z62EiP1ovya142bRUTK241WNCtAaYSE0HZp6NWiwK
GUwVuY7EkRI3pc87/eEwSw/7udtJAc/ZQP5mFpXEhG59tmdJGGEfV+YHSSA6OP7U
CYr+IkHEmUXuRAYt8RuvaGs5Y8lCM7tE7m+Cr08ug9do/yLV514XxlEXF7zcbEOw
04GpSFoF6pXiZUI75mfDOfu2RX9SqeuzPxK1C/quUzUFK+czAY+sckTSOZKmqerz
QgIz2HAc6iNpcTMux4ylJyTxkUTufRulAvNQIgeHsfhMO//VXSJnSIVQ5CT/mhTM
EZK+VGEEIhrc+cAS9VEYnHPCB4drKqDoAPzXy9yIr4s5pfO/9sMk9Ayizy4XCl9B
fVICMEKFABIgfv2Zwgfx2L8bZQC5HfLNyH8OhUcZXHm49uDl+cmx57Jlp6z5JQ6G
9NXEtfpFJU5qFRIXMbciG8hRU+kZExBrD9EE/RTCE1MXQG7PcE0mBPo8zPiOF5dc
zyZLzdOzk1WD8L06JhJt7iA0ejXWsQwIiVZSWN+wiqvKnd/yCtRrCFU7ysyypnq4
cKAJ3EtNR9Vb8FjJPQ1Ckl0xJ3LqYD4bi6lSrzZ2BfuA2hY1mTBQT/D05t6oU7Af
jmwsrvH4nZo7/UYigMKdwT5Qgwm/NHMdrBeJbzfkbitVqGAwMQavtgeiGb8WBa53
e6TZu5HQa/wR7+hqGvE50iFYcdHh1RCQQ8q1s95/5CAG7yNfxhanOGr1rnj0CKg/
j+eEvsefYLivJGCevWqNKvXtuAzv8NinLOuWmoXTpEl1x/kmQyc9pYAwqzYeavf5
xZJzY0eIuF+28Un1Q39jj7yQGcUsXAx0Fhd9iWWGtxM5SrNPSHQIWH/ykZCQiFKe
B6yjUJ7/MxRWlE+Y3ayJLUJsx4hoAWxcBXlX8fL44fvhedWLmmSdTqB9UULjdDDA
s4ReVLh5scfHWMrboaAtuR8VyGjlsbm5VjX5ZMtlvR3/mG3lDPUz9iBbwe9wyJpm
AyfctiFQkCmRKlbiOKVzNJp9JkYCIMKMnM/9grKPaco2Ol/ZL/U3kj23s5XO39lJ
q5P55+RtiLYjoA+Ztp5aKjYfScJ0l1Kcmt2uAWBXdXjeB4k2+McseyKtAqNSrp7v
R3FjxO/GpvQrCIyY/CbzfXLg9EcWffv3EzmgsPsutrjjzn4lfydvTZsaQFdX/AI2
2CV71HD6PLi4sDOw+wJGO2j4iormgJPoNuwgcdo4wGNcRjTXQ4nLALoPP/xhZBD0
EriWS0I/xKGEB1ioxTwR4zFJEEXCRmknSjJ7rm8p8zeeFn03dvDfwsNP79BbT/NU
hhpdsOmltj2jpoDQqTHCMlfT7MyRiCLA2zfBZnet57a2ym8k8JOpHEjcMunyBwHL
1vczG6a2+h4XikpgMDADh/0D8jPgyG/TxYCl/0lYPS0qJhS6Yf6OhaY/PV1dbAV4
iQWqTNvL30vAGoyNER6YmSDGK5+domi1ipX0L9CG6ObJHhUL5xLlZiqQhsFOyaho
VuF+VqWWeExA7HhXVtWH4ST+oWePiTlKTPvJPqpicznt9Ifl6sPwQxdJlG9MdNDm
c5J3RA2j03Iaixl9TInb6g3Rc1579dzn7ZZ30X8rUNPv5HeTsLJhAkOt0X7Q2uhE
b5B/nbOLsn+UR4l5ZG0JPPWsia3uH2h63n0CrufQKU4h6g3LYPhqVroweSw1e73w
kZveQiZj0ZNprYarERC2Ji8kMUvcq3Y50m3XGeCL/e7mLQpxwjzuMX3YLKYH7YGY
b/ptCBULZ/87OlGowa5GGeHymCsx4MzTDfoxYsJGQyrS7I34YzuLYROvm5P7rySw
+Q58vbZYY0rzj+YVwph41RH96C4u/DVCMR4fONIb0BRUBjLGOk3kz8jZbYG4xrNT
vUa1LdSyhyvxc8OdfqRxWtOki+ipLKCS4jjO28kLfNc3dR/WxDm/VAAhrsAXJUXN
xqrtmYUx0k9PTEvhp5Xp3J+yrONcaXsyqTI2eSg/+jP0sw32kSJ+IqTbJiBd2u2J
+j0/bo7iWKN2EENP9AEYBjzedkoK1Xq7f1M9YOtYGrloM8VJuaUBd8HmQODeD/hz
IuAcENvpJtOEtfe53WaG8NjUWEmPq5Wgaol8fFe+YVYxQmH8fdQTiF97dsm+iDwm
72oc3ER7E618F2L8NxXfjKKgDY7S7jYwjyjI6N3YLbwIzVpxPA7Rcm7ELUBeQaca
2zjwkOtNz7bePgTOII032mW+qeiHheiy9w21UZhxrguXV1kw+q9NJzrBTMpFsVT7
ycDCnr+Km0sHb7tWKx1A558frAyPwA5HTex7r2vxB7w3jREFuVmJzX8gVa9iyVrf
luA9nb5C6T+cjGS62ARDpexycWLfiPCPmEJ+0u9yxJ+wy3Qsm13iebh+mZUIviVL
PgX/x7kV8D+145QBYky8XxzzuB4lQThp6Cau9s6x0ekTC98iEX+61tu3rt+R1Rdc
s3BMZQJ1rWNXnqM4psqIgZ3sovGqSCD1yMfSUsCUgubR8BnTApzo1zDTXKLngMfC
z0hfIthy0BjAGc7Vo3hsVOdqQKnvKVTKz9BHuWoq7YjHd/cStgflnnfKCVCcs+HJ
aMfVk45EZqFBbAgPIdyWGJj3Hq8soU0DSQV9QvZDIZ6ImCAlzWu6KL/kGWNCywSm
NG7HzVvzoBQHhc/2rt12/68Gq1d4IxkESHPBBZi2wEZcN/O/uKKC0/mE+oPwPMYg
toKB7uj3tqP+uS/+bfKCKBU2ygLr3PpJoOCq7IExAS79UqELQBs20ygry/mPthwd
a5rgyRQrAba6v92l8+5iRuSrRundjf2HYXvuXoIAov7kgi1XoMcuUnJ0lTiU4OQs
R3YFxOBsj/C3lCMMwyWsHG/Rlr/B9EUgQqB/xaK2wUdDKVYrhZLILZNHK8smdHmC
n+av4tFLs0AZTFpDlYCc+oSYO0ayo0E+Hvo2n6HwR5vS+MbdycdzHTOimRJ5iOkX
kcHshvEKVg741G5yc/o94LYIexH/C2TK5P8/+Vh660TdQOXRAg1VI9TvZzUX0Hre
63rOYGSdNwu6D59nlmocJOG9NHI5Zey6ORKpDpIK6A9ogg/0g08gM3VusP3Rz5WR
ARArgQIO11dm4J89MMS3at10AoHzoSsAbbw+yVmRHiea8aZ8PW14KseRa+FDwgfs
77XpJcqbd3VbZSjk+gQJgm17IiBjfXeYcusFiNv7JQDxz3jrLs7bleAA1jAdnwDU
SLKfNZ+SSznJrOXD7eKcl6JHVDuCHBj+mjLwFk5fRNTsKJN491KnHbVdYVWwo9sS
di7foN/yPGSBCYG48g5cLvNLOrSFd9ayqJpEB8X6eakEcMw9Bo/5Ruin0K/32PnC
BdcE4xuskDaUL03xF64SrdBs4FzmT2pudNXkr7FuWI+JHUHzhJ5AegrVTLbx/z6U
Q7NCXdQbN2XaUhSdKUdj8GDj3vxRW6GOki6RXt3PI8q5WthCpse21lKd3Wp2caVE
kiLRJJcCPlaDw1jUOyRrfYGCYTp6pC7SDi/ieUsSbiWk5m+uMhJsefaR7T4CT25J
7nckrOGRitCGwmZyceWmGrEnEguS95zOdswo86iN+/mBWmO+B9rxh5oNoqQ7TU4D
bqgn22wVBm9pyBgegcs9qo3yuEYcIiqTHi8rKMPcqko+bLCTcNGFWZyFxzjyLGOB
rTYo4TPKngyXBxUrxSBeX9b6HSObM3IQ504v3jKzpRJJ02Iu8DVBTFGIraTKPn+8
aWph9g4xJ6XuDtkjcQCkYp/1XpomFsOpl5tR83JDD1YJB5gGn5t5//U0/Xp55CUp
AJUsVm7Mfu3etbLRoEWKBr7iFnViCB3g7s4duB5Q9Ge+vlX1YB1O3kkbnr/Oe6OV
bJ/TyTO0Szu7MjaAX3tk9hv3YoQDWFPmMdmFK5FeVtAe3vCShOJSMvbb8KyqHPdM
nFlHH1tFu/WvgCBfUjZwfkqcIkXv6q6Wf52Mdrs7ks/sZdyddzGmPO5DWMuDKsZM
bDSuoxMzdE9d37jVn7MshNz/NtKkIPe3614v5d+IvW1iFVwJ/ch3RhRaOsrG8lte
pbcDnoznFiZZigQWeWKPoSHQWb2K/D2zFXCTFm/dVOga4z1ncNuU7jU5VABvvB8g
FVRugBUxBJntjaFIL7yaSjljYwGHRsYguzNTKP3NP982VIGQthc04ixHqZYXPbk3
082O2m/YOfD70ykIKsDV2PtDxRR2BtOhk0oyy51qvi+IuvDS1nJSVaZeyoIhvV/F
m6j5aDMAX8CYinD1S2esbUAQ0Av+ZrMkhJDUpdqH1uhyWplPsYHdLFQLwwEKU1GT
8W5PkXLc+3M+PcwAIr7s3AsnUC+6oDOVVuooMrAeC0TPKAUUjJiUbaXQIb/uwNrQ
yIkFLU/vbakkXv2Y2GVqqOpA7aeOB6A5X+snMIBYi5IpnE71THdAsx9Tz1AE3TR3
6pOHcgo1ZVSI9SFK0VSKM0Lplc7koKXiXqu5dyTBLSOub8arhlAtf9gFpG31n3fh
SSgIDjlo2AX9gnoewYnJBe5PVdcAwbvzU3wg2t9m5EBGDXiPnBu60LMJnch5MDfU
11oxn98npZNnvXCCtgmd7uxXACJ+X6+kbhQFOUwVfPyalF3fX/VEbcYor6yboxr8
J5fcTG8R2VEeQSxCtX/mRRUeXI/5vsOp5Cn99+HDAQ34B03yDj0rvPAYyCWBqGmw
SIhYfOa6tluu9i7Z7ekRPSJ8R9NazBRB7VjJiBXEIKF7N5RaeKWYK/5EqlaZuITQ
/KVPUWjBU3fAhv/bNomZa7VOibmzrSrpFtr7ZzyQmblgeBTFOxZn1mEzeqvInuvM
cTAL6YkTuHiMbuIDOglkMjqe7Qe9l31kN38JGVXK3WtOti8mvxz3zbCyelaoBGd5
tu0qHIZ2l9VNa8QzsFxoGhCUbsGIPSa6x49pZ45KimFGnirsMm4eqQOiH9Jabtgp
lQrfh3ug0WHOQURSXML/aIEKs7vpJIZdeKy+7CBjL5pP4sbXwfkeUNHxhTtt/vt5
fkwZkhAYFwqqNzARQLCW2xRuRPZ4uza0obMTyR5OOj+/3TYFE3risAuvhPYDmP62
5QxzZjCJ95YvXPt6iYBIkns96wS/PT2isPvq6Lr6jO8KneBbJu01Gk50iBJM5MUQ
E4BBInt+NKoZEK0DzH0beAIZ0zSTDijs3kNwk4rSHoWXLbiKy6uDWiQuts47nwB2
slYHP7W5UP2DRZvMtOB1tjVESAQiNhPPmAaCBj9ouzLCBxR7XgW1vKAWRLbY5Itb
YVy4ufVDImiL2K2a0LHgyVhL7WBxuBoz/gSNTqgg6oykFsxCTjgcbQKq27If7Wad
Xsa21O6Z8JDte35SGbfFJ5PXo4itOjxtlmTuaeEaaW25VHWLAYVxN8YQmarMQSt1
n6iuroQN9pWTLR3LihelfwzRahTvc7lVQHca9u1/W1FVenIwONVLhu0UPeGCIbBe
3zxYU/UKVO7CDM+BXS6HTKZM6gS8bjzg24I9rIBX9kVvZ+5uzldA/HQHwJTCPCLy
559HiCM6uwr0tC4s9JNM4qiW5AHv1Q0fM0/HI7erEV/kRUkO7WWSaUrGP499BvXH
76uum4iPvgja5tNP7vcWsDCBhmlKhU1sLgVH1qpa10mdFIKGcztSKysHibc612QR
lpvbEuAWd3L7zztCWqYCI1Kd2m5guAAUUWuWVRkLKQh5QVaPS+xHPitzOMV4ESob
BGN92CFFDAdqu6qDcUIHCkvqKtZOv114yf+R6hT8F3RaHO+n3gV49CApj3N8B9xm
vZhoYFGK3swo3Tguaz2cdeTfjNFXAnUIhMZ6vb2PA8bCBVG+EydVoiI/M+HFZmhI
m0A4cIUOv5O1TntXEsoe6qBxA2HZ6AwyR8SgPRGj1NpDHZhfwGFRSmyJQc84wtVx
Z0+2dqrTXhOuiW6T/a5cybZDskUvdWNdxcUXtMRQUbMlh5s8tPHxjYkncQoI8uB5
SCy94aH1xQgdwK6slwMktQMMis4JOBdRxwueJYGlk5MAn5Tagr55YK24GZ4GaRU2
JvX3YVUSGkSufzV5+W7BC0v/V6rHW0msGwTOYZFUmoDc3o52qaQJn+gh7pEh+Uyv
z+7mNI3lSlPVWpnBQwpdPpMRhM+94cpE0NG919Y4geRlmzRBkM3t8Rr0nP1Uowao
+C08DwO6puxfiB4N8f1zCGC38jVczmBonrXql4tFb4ocv7zGH0qnWgtmxgoWXTi8
QCJQ80zMQbAYdGmMt3Jm2TxaJRZn4/q4dGbxuRVtVoxFXPniF15ny/CnhevEc8R6
QVj9LUk4gGoIrQfwo+TG3swz4v4vx2WeVNguzs8yey5p5k5aledidxL5Cz4nmF/1
6Ho8B5efLF8mbtoviu4ojk+34KkfmfVkT70sxHnscj+jWr/MqrqvT7Ww/QEWPubL
ASvF1pwPwqbZhnq3CYm1OjH6lSGTJfKZL5LD408EPmuR3JBFkiEUQHoy1gK2CGT8
bMpTgpl8pMS7X0BuzFn3eZR1/6Cvs+nlK/+Vb5chTzKFX/30EPinzwS3R7+qIr1U
P0IYh0nhybrpHXTsmMkfFzifaBHfybR1cFdoUm6Vt9PgS9+Fo39ETEogZBvCAY11
0YRkgUzvXK9d3lFhkBTLGoOl4hErpZtv7q9HHJ7AYcIyL+dLteTCUVbrOAZUw8FP
zfYy/V+ohptQzZZ4AfBHk4oEk/6289AtXN1dKanPJSU4sqAOUxHKNE+pn1sYQAWN
r0O5ivrdC8X+u1I1u7LOocywCaw5scIq52sfXpdDt6sZciIAji2vG8em/4Q4Pl6M
AZevIfh9yCJzSlW5Cit0rNrxkv7MRj9zGMcZfH/hxkUWlOq5pc3+Ztn2QrRtVByr
JeWsJUIFNdw4w5BZy+CDgaQog1MHHWhcI871G4Up6S0DcNBINVIfVGMrZMQ87ACp
Q82PnfnRY7tR7s7Gyr7TGR74WNu7jyuRqh2/oo3A5kPq5xcG89EYBsgAQvs5LzOS
k9ccppSeKIJrrnMKS/c2mjrnFQ58wn6fnXmmglaYoczblYqFOkuvCkElo7s5W+li
pQuba+4tW3JE6Xg65Ki6owtfVf92Rg5FZWZkN++OoxhpaA7WddKxxSGgjbl63OPp
ONyIJUY16zaqJL1J360NbVD6NAlu8St5Rq+RX4fTT8wCEvcbA0vHXS6huxbaBNee
k6FssukSVQQT8BE7X+AyE8ijWfSzvtldfnOCYfSsHMZlg2m416aGR3YWg9G3HjpR
y5GSfx3ZGxEdcFF1SrRuv9cXsMbtHTvkfaPSGH3cSOi1H5O/MjXeAftZjL0M0C1t
jRlTpLY/XHsDSITKZmF8S4C4NQD/xKq6viHLzFEzDLb6qq9W7AuThpXBTmWHvtgb
1z7EUT+ykpgCm8CSOnQZen/36ciWq3cZqVIUhHExMiyTp9BtvU/6wItSHyik6Ps8
V18F/xn8PD8Xs4I8KE2cfZriWIdEtpSRSeK0CrWTKk6rI2zMDxOnsNnPLlEWrEGJ
+UU/t7IEIfXBPD2IpSidpdp2Vy8bqVCKaRAIy6bmrfVtmafaFkL2w19zPfbyEJyx
F/yBgIROCqAYAmwnn/69xLXW81rmi50MmfM2gno0nNdnvpa4keeHoXfRiHuuKWOE
iYhu8N+qxZENtKpalykYCPQMxgLKWct5Px8T1RCJFwGkshPhVN05PmdFq9Njmlx7
KFFniunMhR6wdrWUziqTCAHX6gzmDFq1dy3PWBxrUIw7rngMhbXBwEcxyBkQhqfc
8wwpucqu4gZII6ztXmiBh1s29bnj5nMfvvLJfb2LLqAW+t388nIbIFlELV7f0+02
7g4mcOIj3+vmQ/wVRE8TTTiXSED2/6YWoidV5D3CpLI+TLZEerPprJcVnkuFW3mp
7iDKZBK7T2JnLZFsTDAKibnJUfbdELfpfEZn6JkwhMQ3D6yzOpYNq09vl5uHQLrE
AaD5rs9FSYTsnwzH1FBXehB2EjNsQ7Ioz+xmEnp3Dswbbjiv5HNN+BVRmjnLmHL+
M8jFslNui5k/Jy4R5S3kNrdulrUuZaeKCFpIYF5PkM7i/QDUnZz86rr5KzqDaFfm
vmF5leFq+38VncTSk9viKYEADcvCOrrTrrjXSwSOT3/ftr0ydZV4sQzy63r81SqJ
AJgU3KXm9AiX63u70/1TI/E7zmiywcHa7paWsLLyt7W7lApXmaFpz8RTX6FEFV7j
OrObs1d6uIwiOOXmoAeEKGeFzEyAM9GIgAeghAeQ+/FoP23a54+ZfpAFG9/ZNBW8
4n1bxSp0LPhLMWfrkXfmhoPFtmEkCb64SrToFchI81flOpoBz6pusSPUKTf5admt
/schj6Cu7IXF63QdQWX/vrhpMHsDUFU5Ji73PWDQEceh15PONS0a2fKrQLJHVn+b
9FMcZBsn7wcYwXTPjJDdfD44XmK1PL7xx2Kyvzmpt6WPuBXV+7loGQXpATk/HInG
M8H980CypYwtKpQK4/A9qtobP7eBLk7JTEODPHymhA+JXj267uOhyAggmJ+L7RJM
tuwlJv2uGAchhMLvaWdOXeCLicTXYai7v4U7oNGYfVKjKJGxUGz3mOVtiI6iJ8qe
64KAAukQYhIlkDAbACptiLcSyygcSpkgb0EoaxlXQu8Ivh+R8CXdg719KUlrh9bp
VGiHSuDnFFIb5iYe8qLqTckm55+ZJt6ScsW8ihhQaULCUVLgiJ0I/eY6KddOjigQ
nXjfpp2bOHvzmAU/ZeeXduCBUAhb6rB0xTlyu9I1bZqfKT105IA/kmJ/EgL9Neba
oNfgezgLnvPlfHl8dY6pYbc8nSGvRFjZyJE0fmYTYjY5yR3iVV88i1XAblxXcwkm
yccL7Y5FGy5xr3mjdBgS2KKl9uONZMFdd62OlNGXikRCvJd14vEd+vDwf0k5fxaJ
A2G3JFDbm8E/uYDWRGfECtc4XiG3LlKSgf1+jkFzaNHhFG4c1T3Bp9eCAGgrZQhO
eDPirbSWfY5naP1wwb6xsYPKkHuppvtk7CyP4CSBuhrLMkbLYXSPixph5VGNJrhy
Yy4/t/T8GGduxFohOWk0REfj3MD7surBgHxdv6NUIQ/otWxjmFd7mCZRvGGRncHs
uS02YQz76sT+6w7DWsBBhXhWF5cLyZl/S/08ysVisFVnMnP1fb17DCQpJkW8hv3l
Zspw+FUauNVQLwksV13eKGm77ZZKUGBrQHi2hNmE18+983tLgZoVX+9LbiFmbLZ/
JaP7FwLliTQVwFE74TB//NIK3VLv9wUGe2ctbJWqNSyZxZ34rvLLD3M0J7rKEEX0
GG0US875ZddT3ECZDpGvid7zr4GjlPsE7Gytho9CXrluvqDiHPiLiHKXDmTDXFcJ
d1u1WEGDWoAzp8kE5lCcanal1k0npvK8fx/B1QMgbntHVW3MAB/cMgkZY71pS6XQ
TFUsWmEOzlxTOg6O5KzlNr4OB/ozfXHa9qnLMOe85PtOtxSNeIVpAMo5iGkkqJFy
K7eqTm+6AQnTwO4hNgOBpW+u+oAx9zf9TsIf0eiBBlaoBJxrnHInAPNyEXhrSLm8
CGpn/tkLUAWySRsYxVCZsm2WcXphnvGPKle9G/bNKMQUD9/qT6S/sOUKu7RsLHRY
e3noY/DfIURxFEJz23/36QB7OobpGtFnTi0x63JK6abPnziiu+kLSQkLR44FVScG
/3dK66or3fJkGsZ6VUKVR21Vy+u9JDRm9GtAhM5vNfeJIcUp/pa+mDXqMyuzbYRh
d5Zj5EAJJNBoQnen2vEeIxG2VlLG3whm4oIioethVnFaB1iiyrKgFI2WY0+BSXw0
8kkNhca5Cp1PggwTSCrMzlqwVxMC16ryREqd2+nrUEEQqlkrGWHwxO54s6DqTUpc
w6E5DdQFbYEtQt3StILsGAXWMpyeO6R7AOPo4PMpZ+0ziQXrzTicvyc5wGXns77y
k4j77Nd5+yRwt8/gboifRr4ViE1HrYfWHF1OaIkhZ3KvjqW0GQlzTHkNsYgr/1cS
VSmWjbK4ITTnBrPbx35pgLEqoDjS3xDOGz3Oey65OU/HdJp1501rwymWXpBmNL9x
Zrf+w4z40nhLbnuPhGDdfd7+RQedff2LtPk7Gz0ZeqvnTd9y6tfK4D5e9GjDJxob
uCe/o5StchnJ/kI+taJyw5aSP/XzuFKnDUYsmSgxFsOisxDuleKFGLKboxk0wBWf
1F66xFr9m0TsmeJHgWknYgWgrxkNiBE7FfShynCmprXx2pqvQg63vzIMArTdr8az
OYui0PX+ZNtqZ9IRZiUkdhGuTJc3pGX1b70moO0Cc9vwNms2Dait9eNR3tcr8m1W
OLfgNkLkaeMbDlvuivnXQTG2UBo09+vMc5T0iBfQFEBrta7e4JbI8hyyWwZc5PmZ
VmpzKcHIk8YO6p/jHArSyW0pkqN6RSOucTRgiu6bqBFgsb792JoJX9nXH2pa3D5s
+Ue4Z7YE50fmtjgqDvDCTuv21je4zSdIVFEuCC4QWGJfCXmOWnGssjIwrZkFmHDO
pIlBkNi8XQZrD0Ed8WX07mUQ7KwDY4c5qHTNRXnyLCJ/RwBevuZMXE8tXx2sBDNM
iZ/xhToH9jhA/rOzirlJ3phZOC2oGfzmfJ1L8TsL48MQYqcK6kdsTKyAwS/rnCSx
QDD8xz438EbdexDk+VqTofWpL5IkKsW8n7elN4syJLKnmEo9XEtEP/gecu+3Hw7r
uhLzf0L5QYryYv8M/GaXCoQ6K1YozOgVBop/aBR97gkZWNyLDR5au+toXwJhLzW8
CJbrbG5tBnswTu+z1qCll2KA8b7OoNbYJ/dZ/DaVvdVOleGL8TrdQLxRcEAiI3NO
eiOueZQLAMCCZDLQvnWQUwp/Pccxb13Tnci5ECnyYRO1UyPXez9uEHbRuhL1R/ug
XUaTAmgreGlGiGKRRFTBPdMzF/KTpbZDB+2LKIi/1tBD+0j0fjse4Ha3xDdeYemd
SRwHcGoGYLpnhOYYA1IlXPL8Rg4hZQDQQHSl2ukjSEh+hNSHRQSNMCMQWDxH2ycp
w2QbmBs5MG+av5TBQxMKE/eXVJ3lWmoJyJMxWV9Si8zrYYmGow+cjLzDGg6smEys
tGS8ywBhWROoUvBk13YkhJmanhRtTaq9MlZJRcPpmcPnNySIdpq0SOkilfOYLJr7
gd8v7vAhqj/mzYCRHNiqiPiKu8boSj5fs5V+djifpQCNNCnGRI1WhUaI0GqjmERK
SsjeZJbOq5M5XrKlGIz5xP9C9wUZ8Ku+aTpMylzFRC7UhitxdqCv9EXO8i2wVBKc
PL711ThvdLVAUkB5FggbTBMX51UCYS52zNcFG+0D8mZxk9hw2bq50SdkDb25Skmv
ZqTjVm52Xn7LeQGinZ2KhMqs7D7yYbdPyDhSpfsLMNmBfD+XtBnZeFc74R+Ay7sx
t1GmgD8o6CpbtFPABi0d6E3S9cfRT+B8efMmXFb8vAOpRY8yxhtspKf7ARgyliBr
63yna7/taeNr1ylrvxxJ0mNIVCV65bw/9UxOcykW5YSvNO6jnNq8XDG/0DfRh4Vc
ftyvGQyKtTMTsZh1kumrbbdPtOOVoDDlhvH1y9vfFO6L1GClt6nbogCOpzjw2Ucw
HnCzb12FLjx/l6DlHWTInV5ULwKHu4zTxv3W61EolXJdsAU5SwpPVFTiPthzsugj
mq/nNk3/HWXstLUK6dWaNIbagKVjPuTNpk7TLA1AETAGNydLZJLwn/Zb77SLc73t
0h3MZ/LPJD/6bfC5nlZBzqtmo7UE67shqLi5Ak2ryhBBeWjs5A0DP30jtsCAB1Yw
GggyU3OWdkTfyIza7+KgIKs3bY4/T8KZeJwrEyMBPKE1Oa3brD4xCW/YMIuG4P3J
rpHdw4a4kRmZs3Wc0rOkVNMVwpVObL2ZpTOkbYiXMKJdDK19PGPPOtaZAfX0+Jte
EqyKeUvbbPk8OKVVXPuAnezAM7ROxoTvoBhqnbJ6o6cVjYI2X7p7wGpZQIKISSRp
1Zg4jrqfj1WHKCPb/OhcuTm7Q4AGytvFzUvjtvl+boH0B60agv/GC5sib8mz6N7e
+j0D/akOlS0vzfUF8Ag1b7QGoyk10RDnAGZ4TgDU+jVYbWRsKPd7lsjYaXSyhCpk
mxENJ9lALSeWzgiYYvmfWxsV4iH6HCEkkbAbznvcJllUQtUr854GXAzCATDHSeFA
q/zwLQ4iBCfGBR0Ldg9lOkA1Umjhko+qH4ofX9oO3sDOHAs4aLk/fjKzwYKOiWBT
6Yx8Vy38yL1Z+b+vIzKBH4QIS4R6V0J10YGOI3vTIegfw9enjjQEtSscaGbQHYcy
tEIolYhm1NTc4A1Vf6fWuyLJbPJmd0M/e7hsVhKu+nWtLGeYeetDEpq9UwmnMqOI
hD15TJszQInRCQNINbKcbsUgbHVQ4Fo+dCtmnhrK0IBmx51ta3NmyTvSg+EZE5uD
hqkWWaBzyVLXMJeeadEhdQllSy0eaY51n5bI9fmeI1nT0auKUmbZiZ2lCC54cXN6
aq4Xet3tElVxj9caEVZQcSLAsc+tf0MkK8fscQxj0iOianm0B3kNxxj37QQOYrYk
iOlXd5cKxh3NrYYFfHGxTYQ7OFheygM+SItlSNe0sJsW79lpvJjqXOo8eY7xQNun
+kWUJEZVSXV4iboF5/ICIBf98Ag0epmA2kJjGAnNWdCIvzSFKMjtQLbo5AXs0j6C
95H9KuwX4ZotBQS5Vqoyor2pZUv8ml/PP4sFjXLpe87RZbeYlKsQEh6rbqudQomc
q8Y3Eq6TKXpcRgSHha1ejpCJKRR2I3veY2kuYHnIglBJNm627axNCIrgXbgV8Qvt
jguO/jds88240wiADIpjxw0Gnxoj/+f8VYDp5+zdCS/oNwS9Ht1Mm0MMDwLv1fyJ
xTyTXWDz56rT+oNXW+G8cmcsENEmQRu8MjPig7eWMYvIBRZzEE692REUW7zayyvT
QeBkuqPAvrMIrZ3bpFqx7Jy2Eomm9rZ6x/DI/wEurMjuUMxIjydJyBYP2y5R8E6+
OPnVeniZGvbHjGPPG6U8eOslcJIIx01b6XCjm3YOM42Uho6qE7ZYHzfBzizc3Orw
eWE1TTP9TfxrQ+uCuT5alHYXj6N1qb2EI8f0om6jj5bZ4za5jZznirp/uBpP4L1E
mpT+tO6GVHWQ5bGlPjYead68qQZph69Tiy1clYamHeIukU6sc3+ChvHe3v7TrE8y
UhPiKSomSRFzy82+kOAnGmOCMxfjQNsvFlFwfcSoO8O2JNclPGyYVbm0ca38nzcu
3sZmDtS8CcAWJ74Ukf4+WCFEhJ2KmbsjPaQ1u/CgCKqYylQSYRTBEm/IzN2W5QKW
x05BxH6JOtioxp9KaJHhEhlhulteagpz+pCqAZ4GRk9M/S7qh8EO+IHIUEGijiAq
HitvZnjTmauQBRo1YWk5y1ZRVKKRokg93sZzFoP9x7+lByoyrSyH5NUnmM8umY/x
EfWUKgbbEjZPtma7gTu+s73Fdduee9egxsjb3f1HP+pkeTLgYj/1de7Ru6oZXQad
EK2gNme44actAMkDQ2Z2Vqxlkfi7t+mDuFkjIRNj5BAn7Pz/Y1DMIxQTmfHvPHuy
8znDum1oBe2eCMLCzvMX3QbypZ9PZQ2+dmgL9ApxoBQWLb+P+N9wWYAg8pnJH7k0
3Gv7+rwTIhvLnU3+Wa7UUGe1IJFJdBHGqrrlYJ21w7SUPCHZ4rDG+rY6k/yjMUvB
ZoYLv+f6R7eT1iw2isapWUGEcnw9xUp396WXk7QCw+jZLjWxen9OTssiSO65a9Ec
IzsZYFwJVGPKVgsvS7V7iDGnqvkeGYBQw0BPW/1rhLD70IWQEV8BpgDTMhMekmz9
Qp5qj8Xpe3n83S4zBaXOZErzne6+AH1xbTAtLy0w3PHK9LUJ2nsGzz4aelG8kgYF
VClIFmQW7wQRb5bd14+u2oghCE6Z6GxBUAkrZ1107SHkbXyRry9Uk4pUamUOT+qc
daE5xmhEqzFiFWzLVStLx+IVEOM7lSAmiPbtcY/cbB+npEItP85jPO5tlUnXurx5
vfRQjtJ4a1CZNKcjtSth7D49zzhA/RCRpRBBjU+Km6rW77u/qdVjJ2iNrL7e7yNN
tB2YhEaRVVg+yuD5S3bSwcdpK6INlYoGDLOHZWzCiFHXNAqLp1bqzM+OcSh7u089
AUwx/ddKZPjMbfYZBvp8FuaBSPL++PlvvXOA1V2OjlshUH6qgsIR4ZwpnJGQYInl
Jq2q/WysVdUjSEARub++gxJg1kBlxgU9UlBxumpbts5EtMpby3jBw0klzOKMYvxg
FU3XNTo8ovuC7jpzNlw3meluhmwDTzFwECz/Y0oSUdYd0MYHnOYcdSjQaBMseyLx
4wPaciAnI1047DjRIdoFttGHUZZ9/j7LuSYQ2LfI3+HS1shVfAiFxEFf9mHg8WFo
1hTmSeavdlN76UYMoyf/qU4wN9JhOk653M3LPHJdNqOLznK/hmR0WzHwZh0WHD8L
AglekXD+5ZZpnNb6wekDUc5JFI9mJf/vIItHq90Jht0W5GULgTaPJQ3RBw1WEFQW
0npj6PMATlHxpPucS0DUHlVvuRM6cXtI0OGlZSm/5YKhQ7EJhg9v+Wv1FgiLwSfM
BsVku/O2qnsOjacZTIfUu/Fg+xMNoo5lh6m+z9nYiq5hHR1Osa/XlyUWr5olVRXX
4/U1a+t513yXuHnxKekLo1ov8uqvBNFdQxoJbYcYXWEn1e+EEsHIFRSuSx7iQdaX
y6kRg05Tc57f4e1tbv5VkHSJimVxtqIUrp2riMz+rndQqcxb6WLBS5x//rqNx+6E
w072CGnC/8xFp+ntEo+dB0SXq9FuZOJJWReOhpcJzSfZ3tAsKMQuvTs+AvE9MOdd
TFVFYVylSl57JgUx7nKOw5Vo7JftyU2OtLz8NdJg2YhbzP3bcZErDFeocXR5kR1i
+BR+EU9zXWBKK8W/aV/4key8NFATYL8WpyedLgSNkyoG0jQJVfj/eDqhiQW9kXYi
0d9eTEF42H/5c0kKg2Fp3aVUpEOENOHI9e7J6KDbuBdUkdaT0lFjW+GLwxDScXO/
NR915vQHH2/bxaHoaTSThX2y3qn5GyOP3qK9a5RMVd6x1zNBrbSSQ6s2ArOhMwpJ
Lxijy/qqkyUoQTDfLXdUUPySPwwJ198okn3F2TbM7/KHGH6vdQBZgO8wON6R8+lX
L4fTprN3dG00SuQbsM/HqOqtybh6tOKx4GB3oq/Z2wNteaFTnpJy8XqUJbPFVZpG
1WzC2J1kJCrk9Dx0ViH322Kxigo66JSSadk6kWYwj1EGmUKguC34RQ34e5tNCFDJ
M6rwtKgjjI9isl090Bi592mYHzcy9N5DbcWny5YAbsiWc8o4Y4Svhl/JrwhqJ6I1
szWRcBVOmbYEDgTQhk62A0TykpY252KglM7pbUMH2lAoIqjWUdDxsUh8tILiafVB
4A5uxvGkVnKYepOAFKGOle6tRSWd5TwVt4GaPthCJAjwJ4E9Qj9oUitxYubpaYSo
SY2T4sboZyCvq26YQezByvpPDaKfoIJ6jdkB0OjYWM58QCjUFgs1LwXUmIac8DMX
hpU6tFNxUf/U88WIxtDYijV0mNPA7mtBGecwAs13GygEiJGvc+QPYA+7IifvvPWM
h83RkidXw9Y4YjJd+yf6Q9K2M00bJLAhfzfC1/uvsbs7RIID7LuRI0rV5stfLA1d
Mwec/6O5oL+SwLl0pbmnWuTr15JQqCOxvYc2EeZc9V4q4RZsLUx92nWksR2wIn9o
6J8z7GLVY4LtvNeyoub3/bs7+VqZf6biya1LlFZtsdqnw/SvaXS9SBvJetEzy5HL
TjHS1nHccbngDJF6n8oO8xFfI8jLkweVMMochhoJ+H9qD4pPalDIRxg60jSuc2pI
UNvQyKLawOVf7DweA8GZYGEseDbGjLsYco3pIdcPzQx4bD9J2OWzt3Huyki9YN9+
lH3Wac3ks3fg0mQpmcMd2m+90Z0mFv2XL2aAGa80L4LyoSmnw3pWOc9VSbF4A/rE
YDl7NO4FyYA6nqE+ad+v4iOliotzMJ81OO5a5LElgSzG3myNzjM93X9508T2Wggy
Wyb58+N3WhnkAd6V600AgFpA3NpmQS9oC1DFEmRnImEAbb3voQM3VqeviMdxoCgg
C//vxNddNH61nwjsLZBZlFkMTBoTe0hoL7hwhhuMA3JJS4L01c04nhFN87xIHthr
WppUnuKDswbJMeiA6UhzKDT59XGiLlsCpWmq2uYj+T5L/SpA4Je8aWLp4TlZTPm5
jwe2TOxCEuP4ix+VnWtLsLDUqrNsMdI98Dij9cIHw2aCtZAD0LHEbIl+wwSBYvHg
i1kJxN8PxyjuC2SJLPLFpVbj9re/afvWxmROTFbBQ6E98otU3IXu3nrdPHUUGtn7
cxlDED9wmiOJfAeJZvlxVCUelwwzY+uNJ7Y7rPfF9v0o0LnkbiHhJZzWDF6bTA1I
GfgH0BfOR0qwHAXcP38N+bRkOAVCEBUUPv5XeQBo/8BELGPC1BkeYfxho6uJkNOX
grYYmbMocZ9AZFzO56ASMx/M3sRuc7OCHqSUISksG+qBBXaFUgEDCI0kH6pP3nSW
YqZwUYzOLa/sWZbAzgnx6dK9mpj5err1096ZPuDv+Ku8Ej5ugmn6Pt7Kd+V+yFtS
3N/gE/6MUefVE084nisUwmXqSpLX83aew7P0qc4RPKBJ7eWFKWU0WXpqoLIUl46j
8lq0m2GArpFD3jdwj7UUdQVruzsXfcVjEMsHj8ezmi5iS181jKVnDEorFGwzPMlh
niMAWSuGDK7B+tZKNhftcQzQAezUSyIDYoTlwzEtN+/rHq/rB0gIHZy2409gA/IN
j6kvvGxtoHjRiTAnvUgeckoy9ADOZSOZFFYd9PnA3vJdipIB2H6bGqx5xXfd9+yp
hdEId8Vz7rQmXMbJ9/wffgf8JqbzEv8kD6yF+8d9pvbWjcAPL+HcSxFOESEgbp0N
mpwFueXhp3rOMX9M9t74hc7/Nd+ultuzkxn2Ciz60SlmXV3LFC8TZ4d6aeg3zl/g
Y3yLK5eRtNVNmId81/RspvFW130RcZsJf0cNIcg4lBbQZ2YKVl2x1dbvD09+nJd2
ruemMWML0+mZPQTYJNb7PaFIWlFi7d+R7AC5W8xgjIU7Wu+h8M6OzBXxbnkiZqvr
8wOo12AyUT36BjdjVWhi3z/srYDq6905tF3LieFipMEn/XJrfhcLrMb8UUQgyNol
N98viIj2KVlAJfS5YUXeR8PBWl3G9xC7JjiolZyIBcKJRk0vqdSZj7kPaBC8ULW9
anTVW+FEcoX/4o6gmcw3eroFB0uuuqu1bp6y0aOWd9dRGYQhv75Lde5xwlCRrwr2
KycTvc2lC5+9WbrzohNWyA0xiEafu+7pDCG7IxMBlVHV8BAynw+PbrWGS9wwV1hR
hXIZMNzZ5G6iYYcWwZfsDWzRNDrRY2C8Q6yw4nLp2lyH0l3BHLgKBREuEEdaPViV
QWrJ38ZoU9hXMT3sK6mixUjhNkTBAcgOq5LlWpUKaLXewTJ5S3V869qOBxnAnqYZ
v15VtjSKnQycZ6hOX7LDAb+79jVmZo70DcC40+k/GFh33RxRydTRXcEcitE56/E5
NWbeOI/fGpc9vi5LXZZf9vYt3A5yW8H7/O5X/nCfAAGKTc/w+TdJVXddIyxIm9I0
8UbfXgHJX19CxdrzZXP0w7l1tNnN6yOWIfsWrruimPb5af8giODlAugdm1nuFJwB
uJZYQ6rYQKpJW9f3rTXUYb1glo8soLDkvIIIwh82r8qLCMdSzfLcdrxzEMFLIbsW
wfReyf1RCLLZBcpVNmaCCF65B0SNxNJgz6uayEetwrtfI0xGtDUUYPYzZMY7tbz4
7c2Sl8UdMTmchaw/pR32wmoOTSkKn5Oojga9LuK7p21CyOJgYKNC1wuUXM4O1Hy8
/gb+lmciagFQL3tMRM8m0gnKcXcIeGbEYIrS7TD+kOQ7OJJtpeypkAv/dGjxTbX6
KsLdlQeTi7rOJr9BNIHFHVIm3khnRQpf7aPGTSz2toS96WQnp6hAYKdO+WE0izOD
Y4Pjk+SrVcUm+cOnO35Waa37gN+P0zYGEPkFFnaEEyBleK1lTLxsDytbQ8Ft+xhC
eTeBKTJpRl4PCIWkmw6coiL9dj9DUp+hjDbTD+fHePJhTO4kW1V5OO7UxhNRAcIT
5qWBx+yUGjZYma1g+ADa+41qEZwQOE+TkMA6sPNtpD9SUqZfYqOdhmJ5Tca3uHy5
TS6ZFue7++HNSpbdYMaBzZHA7MTmpdljfUhSliqyjVO1Pdz1FFeRs/uhgRlS5yNS
xAYA0bMjXuqcuyGqHhdIv5ePZQqSLEt/kOJB7Ox8QeoQHRRSwgLos7dPP1KSE04C
MWZmy1dSe280EkdSH5VFq+jfyc94O336S5LfQyDlU8q8+LPcx8DKGEX8xmXfgRcl
ckUOzT3mTDb3DvvoRLu8BP5LYh5iC4FItNeZroK4B+inkXXpaAKmdB5fHRP/jyj8
bEsrjBZVqFSbOjAHXfFZYtCwjwQhcwAsdc+nJzujy8umM/9YEVH6FM6fG93Y8hER
QWGp0x/9wj9fJXBqZJixflulAzcVMupoZctcp+omYXeIyhMDCSI1c6pl84t9GuGt
j6pA5nckqwX4hAlDS9LoSnPxFnAVhMQpM/G0MU0NRVNQqQK66q70+vwGt4eyaJ3E
GHHhSAXMp00XNV9X7AJtNTwiIc/aLokhwDIJ0GLTUza2lZdNi562w+GaGoDRXOLX
SO137PkzrxOUeC+VCBIDxR+gEEEYJydsDnzPWAdjuq9FNPkwgsEK4ogQkA89k7uO
RvLY78Ovg+zfN45DmJBWNQbq9Ljdeo7rTg7JKeoMrdUFAMJkFah4XabIsha/awlm
1w/01Czx2mby2rLBLqx4YnXxhK5nBaiWCwTQd9UFP5QcgCl7tOlSp1qYNgG/tQaj
3OdT8VUrosqhovErS/IdZtoVMJRx3y34m+/dTNPSD51w9Ge75MYMdialMEKqdz5j
HtPUDBTvlZpphVie6I27ZXjdqFzxKHzXlFz5csujqD5RUODMMS79/IS1+2QqcA26
BcadKstzgKv49HEd+yq/IaVnAaCyBzcM7GVzxdsLB2rVxL4c+WF8kDQvOC2ZyjGV
RV17rv6I+vGtqm+h91rb7n0MyFR0NFn5GDl5NJCJNvociNOwFpyJvokV5i1XwInK
d5nHMbAILdWbUJeHvXIYJsPCaO+9NZtEoDXouFu/7sYyLB+vUeJFDwc/ofhlP4WX
QIgG0emWxsaPs4R9YwtScf/H8anVphLHbQfmZM+DqH19cFW/fIYctzA7ycGfQvS8
M/m0TSLaL1eO3amTuj3n3xjdxTa7ECXrnE2VWiP5yxWWeKc40JztrTqWFPWlPukv
s1kEpYVLYnvBEZw9PaEqZP4M5IBpx5lBmBDO7gEfYf5reysl7uLoc/G5axui2pMC
sHOaWT6jR2xMwRgj47kFjemfg8fudvFYsehEzlDLAxfB8PeDxf1JfiJL6pvJeXvs
mjp1AleJnHsWf1KPJQ/us+rZCepFClMs9SHmDa+6QhG0gZxwkMN25M48QjrtcFhP
oyEwrVDWPZ0fPqh99HD1hNQ1IijqVqv/s4NbFhwo1wwR3dTa3srcWcSTTF3QRkXF
sc4f54p3m7vNl2iWF4m/+PwYYJeUNsQ42mEUHf8zg8ZBIdVVhr3J+qUSGsjtcImB
47zTsSfXMB4qaUghTIHVG0C3P33cnMJASD7nhfh/MRSj/OtrdFufjOCF/LjxG7ZA
xDS4ww7EEH/RmwkG5ksbKZxY04BiThDqfY83jcrR8PIlU8H5LnBgTEuuoIw2PVIW
kkgl9pEI4yChc/SsAD1T7V9VX68l84qAsqP9hZpXxX3w6D4eWD8PPT/3ue2rbd7E
UNGrCvBQvqWhufpQcg03ZKMbE4h9gzpfBQtPtnYv+/mGnGg96g1SWTwADhXp6nbs
uBv4CBjzRrAKheWn4EMXtg+xGFQx5OQ2z8WkCVQGKe/Lbz5jHSS3QjJ+TvmLDatZ
13kc8SP/ErbtnKLAiHnpQMWC5P270+7stKLPBXj0nl9kLEAteedgKXiRdhOvUmgC
mhGbFAxRH9V7IE7RcTTd6k6s3LTdKBZ2XVlCrhtNDj1fCC+ngDrRDRnNmiVqQ+A6
qeVUQPCPYagWJP5ch2InYYKpa5LclsqpxIKAanVPxqN2MjRPHK9rNUUWR7B+D4qn
z7gvgsQpNM5xPZH5CyFW3q+Y3Fb4EJwqSwg5b09slu1FbNitzGZR4PuFYU7l+5X0
tlSnSrnFUNELZ/EyKQdrQfB9MKmd+lSEzDGCPM0MUhGbPr1HrLA9IVTRgmBNbGwI
Xz5OZ6pCe1qlERhACNRdmfIWCsSOFk3i6OkEnDdy5yqAnAACVD29T1xoKyFWVlDL
voHeOT9F6SHfRnMWDVChLjx0AGL+UlgUF2o8Lk5GpLMHca6/l/aAjy7erlNh9fGD
IFA2w3Fc3xXH3YxBqQLMaJbA/TnqyoxaCG6/ACGgIuyruBlizaTSohtD+f6748sU
seS1nHlspe4CupKfeRDf2EL8kgjmiB4I25qhMmP5zh/9IY0y/tQL4mW0YMl7Ietg
AVFVo7kZenmcaJGhYDzX7tkRA4yZMVgpF5WzZDkkM6Gxqh713X20ayLruzmwG04J
c7DNYu3kyP1EyudukehjYXPoQAyKdr95xEjsJj/P6I6tACMZnLGoxsfREYUh0XhF
FsBgGx49qniWfIxc5NDm6lLHG3ZrjnTQoSsPMYhZLGvnmVhfHh0+WIRAaCBpncCF
upwlkMxakF8T7u3MdPS76zoMYjT9WJuCRUxpGxD2Yc+OjZibCWXaEIyNRiS7W7ov
wGk1W4cbbnZ+WO+FY25Tx4uOWlFbiFCc7G6xRQQdXQZ4GfM6QNXtBWna0xYMyCGc
f+Egucc7d/u4aYWQo0HY63M9pbmC0lkUqQ4DamrUM4ncNZHOywScB4kxURXw2AHJ
n5WZyx+Slsll9CzfH+6xnHlCEUZmTPgeoKQQQVD7P2LmTS3YjZZBAvmRnDOCrNpo
3SIY03mvFVUVrf2NCF37WE6WMdyRr57Tq44QHj8gSgkm8wZfBnynD6oiXqFSbk5Q
GIkFozXnzxC0E0hl1c0N7l5DpHajDdpvYYWPOtWcMtyRGFBRLKTnMQIAav1SuUmi
0gW+m1nLiq6/jxt2jOfOy4/lCXqF9QXSvw3aFddTl3hYvseJcUOLoY3JbV3Ut1gB
M8cYtzSHmmTVPvjotg6MZq8Git3khnWf8gUNMZ1nFO13om93TPStDnYYPMcF7/ug
eq1u7Ay/yjI4vOyCwlTtVXbzPsxIv133JkJMdSD5BvE/GaZ+hUKRlatoBpe40P5f
vOpb0+THtknlgUChoiDm3kxGnTYkJYvsypzoSYyNaa8ya57AUtnwGH9o+6EnoY3h
UukfZdzy7Tn5cEWacCKdxV54wiPMR0Psb4gqf3r66TQFPxLiX1pwSSLpvrLdthhg
SunDAS0h68vWb8KVPgn7OgvuPIBPW3SERHEW1q0NbdClLNxWN+w0Lo1Et3Fp2eIC
mROaUkKN+VKb2OAqHe/oDut16hBJ8CpvEm1tMdKRAXnO796ltDT/hnwmE309jYSa
J1xhVLVtvskjrYYD9iB1FONfxym5E2khbO28iN/UdSvRETja1+00LloPWMxJhMfM
00pDPdUmbwmuG/oEhCycy8Is4SD0pwt72rd3jowDnSXN9pGEd86JQEnHTczwPeLG
0UNjQzhyH5W3MlXDnaTDPNVZtpL5T8XYrxIMFawBCGaEmCYBbpysCdRIYyUrkBO3
ZFRmXB/efJR69MCL66zaYE3JgRBa525JW2WUUyOzSmJWOyqQvX2R0If1Q6S7I79p
dMORnDrWKTdnJgd6FgT8YFh9gCiD7HTBhi2yY9w2f9yJGBJcY86DIsO5ZGuKp24/
U7rpWExWLIWpLKbS1wZlX0qgLbsPY7iMikU58yMDfs9sSX5ZKfvmjNDx1aK3z68/
Y5Ut+S4wBuI5iwffAiyGnNtAd1ttLxZiw8vx61HKyVx2q8w+JYxyqi2ezEUCDwR3
P5UtdyO0A2A9cariIlRi9HUMXndlxDbHjUqwVPaN49skZxcdbfYo01hZ17Omxjvg
5u4QamyEEwmtrQ20F0e8S2+z8l8YFhZhVsPnEx4UIYLFtiacm56mBQDu4XpF8Fo9
7g4b5/9L7N0sj5rEzx5kkp8LI/Cgw6Z+fTuNNa0fVHOvaCqBXtBEifez8wSwIHbt
xUIMAYOqXrqYJsErS1tMbcKpstX4jcKn8w6DlrYjZrVn5ZTLCPMXRksA2qUfJarQ
Mas9uYzwJsqOKJQdbtqAxpiRZ5vUBDIMHLzvmSzYA9kdyLrj06y9F7Doxch6eq95
i78iJLQoxoHlIfsyI6OmD3EQPQLvmI7Jh4uDJnvFzRdApTSs0bLwZnsaGrNHmckQ
2v2itR+KSRyWi+OsF2d4yQADuRl6xBIC1uQpwZuBlNun8Td897v88BwFRtz/uk5y
YafsmWEij+82BnmVCvDoDw5MVuJ5EjtrGKv35n/zZm0Umoyv/bb40p6Z7C8ScecB
5uhA5P3KITi8vYKDEo4UxVViUd+OEXncArwk8o/sFeghmJhwzIVK5h7kJnBgaT/m
hNyzRWKkozmiOoABXxnSwOm6At8OXlPt840AVqOIkOw+G1ofNclDMjkyYsEMLA3m
zjODgP9E/VrBq8oDLkRyEXxkSwEuZ+dvTecKeFusa9cqRsHMCNB2Wb62gPaaGRZ8
BKZ4XqTRkAe8DKHzsXH+lJ/A8MyR02Vmkd7I3kCwBOt4NjVeeulenD3G4Dr/qonn
IWDqJqMaXsVAK9TTiFcxx2e3wzE3fbfJ9S7C9p4Jc1ZiA/K1qHTpytCfyMRjEnKZ
S7ZUCZxQ894hbATX57Qqsi/B7g9PDydkPg66r/K41IG7Laxi1ZwlcxLCfkCPCIl+
9I6c5d6VwRMre9U2Z5ce22/NNa7EJZ7LmxZuXdjQjOahWGVFCSA6GiASl/S8IT72
8hOQQZGcPJQLoqqa5Nmy97NiiNuGGDXro/Nk0kQ7ymkQ/PVEBRQhTQFgpAWkMWlM
0QGpvoEUTZG8BcB+EIU9aNrcDKUe6wzCjhN1eq0OW4pRkvNxtmOVbbSu3zUY4k1r
rClRV8t6Ea2JQQlU5+5NmrqIPUWWMK7rISzIMhq9NbgaXFNDSpddFrNpItQPESg1
jB70WKRPlYoPEWLmgBVP/Oic6pZ3Ph2bA0SpV7WllF7Dk3bU7tjcGnzi/MId2UQb
+lq8iFa7k0FKAMpUogWwXLxS1o07fiyGY9UPJipPKRIfng/mG4+0AJyOqatOUWaT
gjsdzuiOHD3Uf2N4/aTDEKbc/c2c+Sq3nl/6LZWIpSFttt9k766nRoiGKh1TTslT
XBi4mWR75LrsOjBfwLHRror1vkn1ATmq2yBCqhcXN0t/tiabVmsNu0zQwf25XrPc
PnhGSkW8p9Rh1NCVaz9atEW8OED8L9MUK+SUZLnYQrvaci6rqOwsJXRaZ0dHfak0
9GPtzANtmOHdpFopV0RayKNCLN1gEg/fUFmgNMPcrND6YkEe70gql5SRuQI6tck2
Yv4/eMR1P99xUspDzuTneEh+5OLvW2c0Swu4GmXYiF/6bFehioJ1RgfiRhLDjePS
QFqNf68HGMeNft/kDOT5nMFXmUhN9xMGszyF+rneaKtTkNzR8FxoIwTxfhcPiq/M
BzcCUlxzgPiK7aLI2YA0rJzJuvJcQs1mwYzHw2g4bZmrOpMDZuBoS5KD5iYAvAAQ
5xxQAuqlZIGLjH16+giE2ryZmBXGq6IpdHn0w7+YuZI1c21hy9lH81VsI4BF6ZIb
XOzNwubwnwoRh0NyPeUyUW2IHNB68RECdEUo2UzdD9jJqOttnQkbbQ6bhx4fetp2
Py3Fhedn0CtZ0TYZWlWChufJnx346cWf2yPhi+wOWUuTit7oYs0oxhIFD3mMoHpA
RUcVchjnKEEANxtQP0fHTc5kmPU8W9duXnVxvPxb7Dde/Ayai+ByvfxGODn7Grvw
92Lk3pKExIjrjwFGXLWs32sY8dadWY1DVOgDgmq9lh2ji+voi8k35FWHDM+CDh9p
pSyhtyn0FSo6w32cYM3q/v28fNivZ07P3jdc8Mhy/5kJXHcuimVSHypCqSvSM++M
B9vzhgwsT67oJZLEx8mU2xlXCAU6x1WJghvdfH+hf0K0jVkUrfkTpHiYq265EFfG
dFRDmcTpNz4lWcsWITVEw/UnCWfclYLPAEdjIzyooz/7TgvgRgKAWiIt9TUVP4kI
1o2psjgdVkftmUSW2/68Z8SICY3cVATUolMl0JQz19w1k4NgMklix039TAITbZAZ
gRHFjBSTyGfOcMAaxFw0bpXlr49LLbrJ+bFd+zQdsKHxZCgbuCLTThd+zvQB42gI
olY+nxDAHRT5ELXg+y4BrARnJp13u0QEbNKEGtatyD7t+knaTxpGYM5U1q79Th2K
1y8QEPHjGACQqWklbTBNasanyd4eDQ4Y2mR28IdSkN03PxqJjzvC2Lso/3i6erw+
jAkM86H7e8sA4EwJ+/+LWLKLgZQcTMDZwj6yYQ12vujTHUlBKHPNvUuC2Nsh9SHy
IoM9QLZ0EhBwF6T7KTyvMNUteXPye1lC++oJSNPbfMYJsr3WtyOHOEBDFRJnRbSZ
vpLGHwmwah5Uyk39TvHgVxF56Twx+DNXNP9Q8Pnxab9116QeBfmP4p0jNI0hl/Vs
5oBxspuKz0dtqWCE7BNZ+WV8OEfr10xkL+gfSrT0/mgVkEk/Rv/z9BsvbXRcAc7A
hhPjW1bMjpabOJPTQhDBwqkvl/G5+qZl9+DUXr7Ba1j3als4UBx15EVIWSThfQpi
gGWdxbuR0drJQ3Ab2abEvF8YkoeorxFC8lepnfm8C4Xpb7d8uI2uZAhA9aJlNdvJ
uNcOUaVCQSGQV2KPs98r2xg/LQ/hXZuwiXaK2wgjFNjlwmtwzAVBiDBXNQ8IArw+
arFyyp21gL2Cl8ts8kEeMNS78MU2yEoDR12wHZw3fY5C40vIJ2X0s09pSWHQaUaQ
45HgEzyq4S+c9ZIP1DLZ5ZIz8GwsyL6jhd9VoKu4mbTZp3y9pbc6PQHXVNzEzZ0i
Ps7F23p4EF+DYCLgZuH35wGI5pwW9xH9L9/xthQ83HVK4kanUrHA3r/MNuE7PTk0
4BvDQpyOt+tgcD1Mk7xLtzOXqtjdAjL8QTy4LvOjri62u9LugxcpblOMQNW6d1Uz
dV42V/wooZpX+ckCWAehpGiyRKgrboJNSEUVBroEYbUq0Qc4y+7mk/h9NGxJ9Riv
aD0/A9oZPextQEI2bT/xaKHhmuH6tqu4LUwXg5IQ2AFG4BATVEvG45AfycmC6mWd
aOO5LxgiRWJZVGuYRmGZ+ycdhtUWCR/LdIDNuW4Sq7Wurx036liY3jc92LufK2Uu
sPx9Ab1+frRqAIbywkn3/X9qr4dHnnKXrelFYNiHHklWm+Se0lix0dUObXksWeju
RB87uSY8DsrMuPMS/te2wyEZkG9PL+5WfZVr8ZOx9T5h6xbQ8Tz38YRwfu+hg4XA
cICvo9BqIPCJVVoaiTgHAhzrIU3KwVsE5cGo1R7RCh+L8Rgkx6CSdU7youpKS4bM
ggVVGXKvbRbHXVxzrAmARlQNZNiBh0mfVKKmXSyZNTOFrqlUEOy89vQgtNgFBzqe
k+xaoHShI3llsJEevi/RHF/qnJC/tn61SVerGsr8Le4oEx55zLpA9UnMATgcLVkh
UsRs2ZXIp5JV8vINpfSxcgHCfd0nfOtu61NS8HCQLw6Loo9uM2VwANP+w0woh999
yAW/frtsB9CDS6U7KrygJR6sRUkpYp41E91FfYy+F/mZp7OnxxJWaAZT7PWiaXV0
z1c78FbYaRdR3c603pyATkTGpFSs4QkLZkbxry99IauZXnB/U87PZ67SWcnfx3Gd
3iVnl2a71yF04Gm7J4lPpksqTzpI25fr6mjsHOTHXLIA2jurN9IwHu11UXtOWG4R
A2O3jn2Yo7Tlae+DYhT2hCBs1KwJvpH/7nFJz66Lt1rNZaWAuPdukpGeT2O2fu+e
vmXhEK6TLnaDsvuy+19t6HtM/mpbLHF1VhJy74AbEwHYU8sO+60V7HBnK3AafNCD
OD8vzSkMaK31YAeIU7hRm+ozhmAG19QlRq72c451fDDW0XZdqSrai5Ox4JXRsb+g
hXWbdoiGxr0lCNtTofBY7cfbklnj/0QUdHifH++UFGODy4PUBvPMd2VN5nxzg+U5
CRcwIZ0lFJZ65TwVzuo7dGPntzmuWJNfNh/mvstJ4iYi0HEGx39mLx+Dj6v7kRXA
1irfVLeMLos3LOrI4/wJQH9RN+bs+e7JOUcRfeFCDJ4fCqKJF3NFGChpTkSJaLjG
JfS32ggp9GnZFdpRu5pHPmS+1Av927KcEq83d14P30FNYfUGO95f2s0teWJk1LpT
RoXYbd9ZwLWKCkF9xRg/u4AJZEj1/rJ3O9lSLa7uKGbU8KFO/GVhtzP+lKiaxzyF
GWeARP3QG86t68bmWDPiaZOgYqampZFFW0woEtndng68Cw4NOajAR4U7qhwQDi1W
fWx5Vh5RLMePlOSj0huYxjMsIOFsvpzOeCDLd6zWReHEVfafFjL+m142WSX/+c+U
qvcsle4bd0G1ak+vosab2VJ7x3Q0/ijkGPMaeKZ+tBWb2YHkq78OlSRD6DPK1LHH
VUK4/OgYt1UFa3uYucRcfKDjMBff1Ul7NzEjnS5LGW+gMG1vyoYLdDWHJJjwmCLl
qVWws1FBI02v8S6G24ykQLPgz+km1pcsKotdcLlM7Yg/jI9adcIY63EzabrjtmGB
BpL4XdIuei8Je/DTf5qdK7Dv/JraxK861fpT0sFXXPmWULh3tFZbxZ7uS+liYYQV
aYbOxUYQCfW2xHgsD3XytcXZyTkUu0ZKwd6zeJ+V0BQcwOYT9CPpOWnJnLIMLuWG
eJRxomWqDkmKhiSAfhzQAC+CNeIw5F4m7juEJh2u2QHRqAW+6iGTlFJYEERyZDAw
2+yROZ+9VzfwkqCFYhfHsYx2KRAaoZhuWCX9hPDP0NfZIqkLKC8OmvK0lYUR7Y5g
YTyGFkPl/V55NLrYTnT2zC0mbPeGVKAnIOkGVDd4kUy64pyaMq/gUN1GM6O0fpny
XlVy6vx46s/XJJfakUBPBh9u59br9kj1UlwgbQ2N4W1zTu+19m3rfuU+lVNE8i4L
mn1JfKk7GoGpQEVuH3mEBb1JChsHsbvTgBZMzlwAV+HVjMICr9k6Pwjl/GrUXhoO
n8zPdnoPcfuyNdxV3IFFtvEgfu5hGmI2LigTqx0B1po9+Hzsp2WgM0kclOMcVzFz
GAQlcfYZNgiFsxISoKjtbDMQnyc6Za4qUKgnwWoYMqs/TZn2hGAIZAoFoFnib7I7
Ub1Kj3ibUMLB0So3ALRYxHP4daFqm2N1klHAOQU57fPqnyeGfW2xIpqgBqQ14rRY
O0nBe9FcofaNVsinHxXj2Lmr5XgXhQUj16P3AdyHFZmucDgsBirBvi4Occm7yiBn
hSTIK2mEWR50babit0p2GFYimlyNFO8DVpGqisPIXO2EvSRB/izvCBxl4RRglMdo
PK+lGU+/WoV41j2jlbyWQAIOUTxj1xjgfeW7hZyGSc1lhsCCEYnNkik1oyS5/LHF
zAZj7entivFJQu2FkvR1nFaHeUi3lQhjSBreYeEQLUFjTYT9B3wDMaL8WKPUNjKD
b5ZYpzaaVEovSyi4lR8vfLhYFGxJQYyj3zQLNtzL+39GdygkTTuAVB/682OmD0Ax
QfTfqycNlo1IcsJsMPwVC7ThrzZUA0hKaRFbG9GuMxttGfQhmzMkyF72F6DbtMVJ
4pERuElmzTYjYXJl3lXgwzTmUeAo8A5+mQoJIzbyRqiANAoFUAamuPIdJBO4PMNy
wzeBObVlhF1pOmHjx81yKYLYCs6ViBNRmTPlQpB7bh6cBvrtsFTIlYo3D+wO8Ox7
ccTXlcxNXPpyEQGBoDJXV2TZ0grajXrdO+s0/ikBeZkVaII5ComISSM2rcnlY2I2
CBV6An6f7otesbLPzgrTOGL2xEqXsXyYBJ2DeIBbH1ipGoppSJphXEkftM4D1aci
q+J7hjGwu5jIm8a/mtYk2v2tXHUvoKdEwTbKfOy7T0N8w6H0QYbPTeh3Sa4qK5mC
/XGG/notNG5IMyoC0XQHNWUVWWcB4+P+5SG8+yLLodgyRNPANn9rQ+ZWOYtSFXfG
vrLtbTbQe4YKRMxfWoDJIHiZeAr6fpvw0VBVBB9hn9lq746jSit34WVVhh/BqOTO
B+wxwAy1LIC9fHyl9bU6sz9E/MxYXpfJ4IFaZnYmgPSVmzNfHwV/lTz52GbbORey
XhGsRSlac4KNcfJFMQOCc8HGTI0t34OhUqKgztJ5roFnjZ1d9X0URMgOsmUzfr/O
6XfQVyx9Wi3nzf33+qKDFmeJtn8QG+2pC81uszEf8/aU3qQ6Q67qQ60qR6jxTH+Y
8+1O35IvvC6kpUUSaHv2krA1Z1u7XEepKsvy69E6YVgQ15LENxL8hjYNgKsLtPoh
b3Jz0a8Sc+8f6OeNllup0ONgWxCPU6P6sGKT8IlGw65EQM1OgMtxsPB7K6M85kJ1
HR/yXCNTUC4DWxI0A5pO2HqH3Tb9FMQT25lMal8JCniy4I07zZB39INer0nlhtJv
GiXIA6HDhtgvnUx//5TtgJ8YfmBXo4yy07z/QyXP2qTjhU9OE6OsT+i8h2JRoeF+
xkhhA0gE5e4y1YszJzwLwcHDIIkXRhQma1HUFQeqXbxAK1rhuKK+tIGRUzutY3Hi
9bbjRHqqDipM6brImRUN+3gFc3KMtTI59xw/oWof9AC1Iyy6B9sFSq01Z3Civ1Ga
BrVmGMpFM1951JZ2xueOGakUH4QOTCnqHtx/7b3KIRrVhcvlbWzKhgmbxHhru6p8
YXKvnf6v3f50JWZuYXcoVAcfQeAuxnm63slRDX0B4CBB7yU95wQEiTDGlNwCeMnX
YHaf3By7ninmEt5iNV1XhrUNWK6w3kTMecJV+7fOEsU/UloYTqejYTHZlmt0XY6q
t00ZWB3x5Qu2Yut4B420DCLnYG3WOnQpHH360Gm7qkb4QWX+pn0k5KUE57ehqGG9
rGzdYuIosfpDi/VH1JEaUeW2NjSf42HiJMMmiKDTfakdOR2881QHXZYdOdtG7JPv
ioTCMOrqmR4IK8v5nklTpg3hR086aK6D0Vf3pzehsMNk/j4bcohQaF9aYIxl9Q8Y
eodjgXFIICnwXcp0qzSkGLr9a0pkjxgM0wWrUG04PSlIVK9pLp4U+xgux8TyP8Gt
lj/ww9nXk+AZA2qzbMGY859zY7O+0M4qTZbvFRqESbICdkf83aCfJBJrbM9nIANz
iw+Di+wMplz4g9wwlXrB9h/mr8N5p0cqipCV9XGZ/x96hhUS8VfZZ2HNei3/Ll2M
nCQKoee6upuj/CtWQLGoC7HSXF3Md2A/K8l/XtIz0xtZqUZHPXuvtHwXeL530A2U
8zCUIql1RfHv22+Na9QABMygvq8PLKlnwXKn3jBtleoO7ELfCENQ3SPIRhms6+eQ
kQLWnLzGLZc+jOl7FYWg4vqGavJHnQVQ4IEgxjcBrhB1G4O8Ix+RU0Sh4ll/HTsT
sNFOtqnyh2WXY70RMxRx9DVfr+sKvQw+mj29AB9YUutz4GtLaCv6zTuKaQaQU/x6
D3OYUvK0Kq48m261GZpi80bfNKE3a/tsHLJIlDXQ3KZ1iKlLGvMfWx2NBURBnIiz
KLizUZLzVQmaQJerkLZjKuB/4wmGwlmmCkn+RE5620PDTe43QL6RW0sMzrfmjEO+
KPvW6Bm1Ssw07voLa+WKG2OJ33gz07uObggVDFaWcGlKw8E47H623H8ZCUD6qial
7fw5mXIOOJGQ1WNRv18yAmEZKcWw78S4W6uGYRj6VX2k3qL49RFuv0vQRJG+Xs0C
SPb2mYqMfFe2UTR6WtYB9/7JH+lHp0BNR9APtrcXFbxr9YfjprkUHF7+L0xsod4R
Ybkw6Bv3c8hFaIJVYojhi6tVAyYsc7JafnP6tFKfE0/5SGfmcO176WokMZ1ryLKP
/mMjwfB/VULHUWcJ0mcEwjDS/s8RLpduekUth1/VAqRbZQjHz27RKK054+AuEGBd
Zro1+M1a2o4ISuv4kBsCVrCTSB+2+zPM5u+yctgrIfiugGUx/gIDiaWt2iYzoieT
ErNmCp2pZWU72aK+AdmdFixdwJffPjiyIBK2Lo/RoMRQ1DNuWWyAyPjxavaI+JmW
MG9tL+Xl8DoAxFvHlJf9zisiN0pTYKLaU2XbSdo2QvLfMuN5gST60DDjg7yOHGje
Ntbj9KeQduolsbg0kUh71bKKUTTnLwsXdaQblfAWhHChUoSWv+56I0sY9Mrtb7DT
ioqzYdsrqTNANCmeMRBEBEDwbJuHrUpZKN6efuizRgMitx3youwMqwWbsw8oJidJ
XJaCPIZE2aKmTgNIBvmR/ivGv+oI3X5NvcboRl6TgvPTxwOA9PAXRveJb+/YuMCW
4VD87bNx7wHQSt6eRyjEbRshAXIKPP5Qb/88+rPAP9RkAl+A2097tg4b/SruYoHY
VEPRY1zGLJrHtIX0o1zTrvpE12mewBmFpvECwFVQrVeoj4hrpPyaKPEDcmR71uk+
RnBvtUv1bNVs+o3UX0V3HWPxMRovIQE4PWH7cAij41mUBgTE0v/T37eTGASbHfNg
U+LL5T8MuXhLANhD39MDi+jYOU5Mr8e3TNN8g21bN2Tw1MotRSvzhFnKxOyp4OsD
zOsP09GIxigp+TPMN2XSOSmlAxOts+4Aa4fTc1Q1kCvXfRxhdZqdBWR4O5v5NzbD
Qa3b14mdFlcLW1oID+7eB+uMXacxsZylTg4RuNo6TPN2HxUO0hDyk3iTAsp2s+ny
I0CR1mxLHQ83NH2A4VrPBz3yKe1TgttZfU+Kxv6hZoGKehy7z7o+rGSZg8G/mmaI
1Th2gOfn2w4siKZfC2DxJOn7FMFQJj/CA7BxdVwIc7SSZ8yQw4agMLgtO870Fks0
Vfr9N6Z+4WG14iXz1zYX/8rf8sPhjJ5mlrzB/dOy6EgFoff8azkwBtQ0EA4EILex
uzn3oG0BhnuMs3zLfnddF5MKVpyzkEvAcd9FbCS4IN9jPCb//EsZbzB18mJuHNU3
LcIlRSfzUTO1WneahD+iUJzplFDyvrFBYzssyo6fIlnJWY1+zTJQd/VOzIrS7T5w
Pdf1cSDUi1nGc+bHPfYnSnEK9vA9W+boOPYo2zZMQBdTTPF1fzYAjva/fEbqwjCn
YAR7eUcijyTAFA8zc/DDCexmbDNvp8LYc5cY9cfPOOi436bbaCuy1sg3E/YLw3d4
yeckXKAVJlDg2oDhY9T7yP6afHvxs/VOh2THS7xiEP5HZzhQYdISVvFNbuBb6FP2
lgUNsy8iB4jNdQLF+UpyUGKzNKGdK3dDhvXVBWR/Y493VBAMYB3OHxDdZlJ18/qd
iqr+pkt+exKB11aqQG69deXmfGqNMgkpY43cFfFF+Uc9jEWTbg+fojIhWrTLOzlI
ExWx+AW/B519fYg3kE3vNOvsIzPmfL1w3oA+HX4gZw6fmXMO90xAWiLLUYSNxufh
mnhk5AMOZxByDd8C7ogUO+cVh/Tl3NhYTU+MxSMbIFNRWx8hM7loM5Q4BjnYgOpK
vP+yDheEe0htKc1qo0GXKRtUxudUq87+eP/Er+It+NLZLDCUwMqo0Vi1m/Pw/cEb
XZ0aj4btuMOZu7C90+bdcwlO8lJHvnr8/UDnkFpsFYyFEaEH/42DWf4vf7aWNlUM
miU/RUf+eFrQ68WDK2ULdy5wFUaulzVLr+ZZunoK1yxlHMBG617L69nl48PP5POe
tIKe2BPu52G1HIT19v67zhIGARm/d1FQuGi4+h9FcKwClHEYELjNuyOerFslgHGL
rQXYwYrZSptotpbE5zz73iT3rxRsbCdXKSAY97k6Or50IHVmwwZ/xnGDgUpLs49O
IsZfMExsMu5fXkJA/SywEysyWBS3wp9f+gqtj/ocl1Y1RmlvYWREGLb+ivRZr2+L
1ZpHXnvwk+BySSaoRNOl5x9mpUDCEye00dCiAYOKsqoTHXYouPxSeN+ERSrEkaid
FoMTO8wstKcnWuTVwbOGuRcOKZstpCLeVWo/G1oRQhfjPuVY/qzXb+UJkd9c0OSr
egeBjOkcWKDR50upAF9i9hn1Wnb9cd6HX/vU/PZXfOjYxqygUHNWzG/BoyiHv9rm
eo8vCh/onVUykDX3WYfLlonqXdcCz1WpD3Ma1Bf5bU21/8xMqnIH6MAxAFb+ahB1
/qthbkx7yDDjxsSmuHbEFo9rmU/+xpk9WMhDBwGuYs4VMwpKZuvkzlsWjVoyu7Qi
pKBZk65ggZ42v1Pnz9fR+zr7IW03MuUbHE36JNjVlz8mstZJEPBBSNmw3ZsNCg7r
3NWWse1ld4D6L3u4U/zFKCaIOo9+lllG95wwDYbSzJW0r7UZQMEInejFQnqb+27K
4RrwGyAHslWCBDBuJKpdMPEnW5QNGIxj3phnIJbSJ3c+7QSBnl46enQti3PvU9wM
qQcLiZul+98jmbuelmV4/Ftj4jfYNof9nFFU9baYqkeTwoc9XtajaNcRuZJqRdUD
9as/ghsm0Dy0Sjzo/Ve4TOn7yyK+JfoIZWlQaMm77beNCIEPnO9XHAMVZnhOZro/
VxgbyTzHArZnBihRcv7VeK+dPl/UpjrthLA12UDo2t9vyCI2lUz33x6BYEW2ODHB
I9hAZIldJPQXoLWoYszaydRe+makuPg+sfuzTUBPGFRwAAjLDz6VA1yOJGlJ5drn
kepES2KIRo4citFnlhWXSSrq2NMr9YciBiw9xJZS/VpwuAdPedjy5tXTV/zEi37r
wSI8nixMv/e1oQcR09RBSVHqEpNhbVUmM80hB07y0vWUj8rIkLDheyESVkWiIaNY
2EWhznUqoIe4FISwY8KCRzIlUO+EsQ7n8zVZEdrTxwdOyY/z3y+P5xbwUzaKVued
Git01/WZzwYGn73/jNhSoeNJHdKE6/5Fk7AccBh4R57J/ggjrsYGc6givsABYiwI
8ju66il067EvbQzUefPYSrStBusR/gmPcgCxGEe2fWjDuGQPVXTP71SRoqqldQfw
XqH9IBZVMJnnjP3EaSnvm54/4V52vdKHWpIQrUaIGl1ULvNXfsTNv5YXos5v+VcC
5qPm60ukerh/rDuTbwG9OHOmRSCfk5uFOngr+EBLMXFyCUj8KWNTfSE2DFPaQZIl
NIAaDgueCCZPgMewSK3JncGhJYtUlJKLw6RXd0jo+zW3uwcVHKfNHHw6NGvbW8/N
pQmLjAL1hABvUu86GtiE9U3RDjXU8cmLiW+6k9abcweIuDCmp0YvXR5z2wVF9U5C
rf5zD35lqAXGba6VhYdO1+AGxotl1828Z0N3METtVKGSTdcuHXkYzKqh1+zznYA1
rNbRnF+EZdCFrEaTRFod+uPvLVJhvO5VoZ54Ihehu/bV6fVA/so9r2A2JW+ugUNu
mdCDcD1rUhBvOhltfgwQNWwVL+Vff8KylCguzttlURuaIBM7E9BZSBFJFbpP86x6
Iq5TQQf49w/tAfxt4wGHJfShxhZLVNICJQGe9MOS1fNNJno0cWNY1RnYg7QymB23
HHqmuXWvubdCV8Uj1CM8AUGCWxCdyizxIp4MDf+ONjoSrXQ5a8TfkPFEz4L24Bl2
HaUdIEyHA8u3nYSq4TcP3bGIoOX9VxD7H3FqSHkXLSqg32uaYJSe7qneZohX0qmU
aIRVum1Rbx/lueZiRNiDwbRAWKWQ/OGZj0PWg7nALjY8PEIqK32hywDExUqQfV71
LBRKt9wcmYchgp9x5SQ5ujqCvknt41zamEHu3Mk3q4QxZaG0JHqMS8C7bqs74sdp
9d9FYDV3O5BB5K2KMIIX4pStmq+LklzgAUWaSgR0JvQ4dSstsmxnVYHHHPnhLsTG
MOTv3ntY24v2yp0JhVzNpL/Yjtb6E0fo7BxUuWn7wR5SkB6ckj6I58FkoWOwkjrg
7AdfjG8g8UrBge1MSMGu5kfbvkNNjzveIkRCuyHLPmMH//auwd3qQp4xrvIlyDzZ
g+JlfrOJNqD+5MxjK3oicfFYaHadvWSfob30qIpzOi4fBxPwHbMfTNMi7XRWdewG
RjxObJ2pPSMnLAA6nWs2Hqz2wD2Kmv7+dbhDUZtLZrIzo67xeogVfPpXu3OB7e/R
fBnFHC5FhKeUhkM44Pu6dZbKle4utsTY7IB/D53hYpJgA5G82xC5kCcoTq0/6TyI
P5fJ1AXIlmvy32v0WFnMfsYAHO8K1IyaLKl6C9uSGxV0SslTYz9MgTwg3dvYtkfp
/CZ+fHkxn019RCTLVZf4+mrmgpGd8m5l++LimLe8pVwjVFb7ampcBPoDMlN+SZqs
vp7zV8b0+vkZjxmaGKtDXAQ/9XSkgglnluithQMxs8HxOCihczyafU4IuUUd8OSh
oAyZobjIJIOi9Oq3I43sbPyYYnTxCZoC1WZ8KRMfQC58VeTmoX/PZMTW3UEayU65
hVTq76ZQXekEeS7ERVT7MR+cySxM/MvNkTJxgycV/ejC/Pqiv/6IIK3WF2eApKn6
/Hqm7irf2Z1Q0KOz55IxZeirHUWfsC7GXjH3977Gqh2xDpOHxqHN64xW9ZE8hRbf
9yDLryzHTX5fipbdXDjjzzfmysx2fSve7gKSPmjIEWpVAep858c0nKASToyOBIcR
UhoRNPzBur6Lo1Gnm/eyi9IOiUA7iITbM7NWTHnF3IOTq46K6QXviLeYvWSpn7AB
UtKZKdzwq8wQk0GIneqCHv0BND1iLlQf6pR5xPFR+gXWPXhtA1j1EwK6R4cLEM5r
7G35lVlY2QDzeqkuJSOuA6fqVWWWFxj7QhBvLkDqL+r9i5ViOA+jNowxbr4xOd/m
YNgToB24fQo5OvrW8nxY1zQ6qT+Kje10FfK4cuo9cS9Up4TGyo7qxXpeP0Jxd+O8
oqWCYSoD4xSFYuvVmBFXKd49vHWlb8Gxhrqg86hW00/0Fo5YBCgeCrJquTY+KDTT
R9CuiIKKDbPukcNuzoEiqonzjUAwfqVY5fbdgvHEVMeksp9UVvlpxTE2uxQIwGJx
jzNDwmHnm+5IjuWoifuWCV7ChN62whTNowu9Nu9yz3aPZZL7Vzig7VcB67YAAX0Y
ATVuaAahslczGpLqImCe9NT/55nvRbGRSbFWWZl8nBOPkwue5EbJRnwXvPtIN3hZ
RiCuOM0i0RAn6t9/TpriKiwTidS+tEGmLnSGYT1WNTzfqXftr7R6vVJOWqyroMQl
Q2858vYNkerExzioSVvCMSk7+R4BqXhrTV2okL9zyZcYnUaPVyTY0nJl+Xu4j74D
+BN5BIC5+J1F+v83FsgPvFYWGF1LXF4xpfRBg1Nwh030yJABS/LBXgzVHJMdo7i/
o1WHE3NkVqPksvOYpAiIzb71OLgHuCLiiD3ROXTf6qBDscBeqpk3w9WXw76G/5MA
7JMWjoe48a/kr8dtx5Enqho/AZyTswXmhKqj3i0YTzwBmhUJJ9JzrsWJq+z0HFW+
xGh5ojwGiLkxmrFa3b6H4f3qCFq8UzvA2qGggbN38n9bx0OQYqCreR8WB5kQsc30
4O8oaazESxznhsAzlvY13uetryhjXihG7+Clw8Uhnk1t2uTPrIXVA/Ja4ATEG9vG
mNFY1uTZxL+QEInjAS6QW1RfJOqP0nY77/HxTpHiObx2U7qxRBgSLCpgtLMjJ2vH
NYNPG46O9MCRNfvmEPudJuRFJ6iGyomnAwxwRWNC8HU6RaKA/5O43xfRXE4kh4Vo
8PJWxrnseo/IBI+KRC7yz0ZPEdIAfJ+nfOYtADSy3vTC//iecSD0CfCYvNimJzkl
bCLe2TgPt0MJU/uNamMfFYEUWJhhnApgOn5w7sUF0y4oMa4v7IpbKOxzVxi27sBP
8Vou9x2de53e8uy2Yih8Tb4GLZ7m0aWFjo77VdgTb9S37xtrL3oQE2n3GyiXnU+/
hczhwSgIKcb/Y/nN2E8mFOAnlRI7YQxShPJzxfIhCLH61//LsdD/aDEr1gL3aNNF
gQk62+8AlbZIQ1cHh0TVfmqe8vgF6lguTuSsxrnDURqQxOq9HjeKsBop/nk3zijF
yQ0rVjk5399PnDlEPB7Xees9+VM3KrDP52xyfUvOzpDTvfUnCBOEhvhHhtkqVmiM
gRn4qShafWTBFsmGTwxnD8CC+W8ppgTt5SyOia010oz+FNyLdZtq5Zh22qS5Is/y
auUbgbf9LLOUmGz/JChK17WrL2DpvRpYPOClHjcuUaLU85f3oqFdkHx4O7G4t8Nn
YRnUpoQ2p385J3c20ck1u/0YGfVgVQSMfMcdhQNXXjIjFeRv/sm0vRZW1EEBiI8L
O4R3zYcXxd/iLivcKKa/chB0NcMuw2kkN9AKlp0QItY9mB7zf2b/C0VcGQ6P72ks
zBNpJ3Sw/9Q74IlxZDa2Nzrr7AtwQ5axypXCJEsfP95KfyvWOK3+LmTI6mRpmP+l
5tAyhaOxikc4O7/n1bk0Hr+gdviMuLf4O3nGfT0MS6+yRN2bGdhsqJn8X/PpCci5
7ll+P6/ql5G+meug0wbf+lsNufKn+ItC8wmoZ1vekhIay/Fh8CeIkqaIsxKocnza
96v66H1pyazS12Jx/LOPVRIWy0A2x0hPjou2D+OeCuDZk+N8aICv1ZAJNfT/PIip
NrnFTV5LeQUe/AxN/dQJNzYJxCLOXXsPWywIiKFKnwGNC0lTw9HWpPzGeSM62OQO
gry77V3OLxY0ONTC1hkCk4SJIAZwZL9BS3ieUZhyYIQcvygnf3PbUThWV+qDCV9O
NqfVZQwlWZq6L7TCul0XGnmau7ACrI+EC2mkpCJ0uRFHo8l8DO5yRqczKOsnjW4c
DkbOvawnPjHWLYEp4r0hzgeJ9RRg+DiEKMuXQxOnNsjxXylLGtzlbkROxkrICN8l
f5MZu3lDoujZpbT6NvwEhTPvydIqqpQ+GTFC1Ot68Pc1FIdUhCzwWTDwlNJUHDQg
o3munZReoM3FAXX6835WNi/Tw3iaLsGtB8PEka99d/eIZ0+L7ACAvdD5/qLMikRo
XX69nJPECRmkCFWMJYUXouN7b0IAK4T3soWFgwpUXuGL8CwfatI0dP9ZxCUd1zmI
ZV340rUFNFiCKnIGE1c12MTCzJRf3bebkVP6BCk+bldBFrGqTsCl+cGTerNwiTy0
Y59h3G26jO+PySEskt6v+rlp0M8Jm0ToQ5aA2KxGXontgFnG6yG5wplx2OFeUbiS
wVT1tJv+AWYkCq3MXFTy97c39X4rN7vUA+uMPJtsDdYC5058t7aK3xnYFVSbGUhO
ijY5M1sK4J5XFKmSN1canZnXpeuukfm8keVb4uD7+RduV3ze95xqvM3tPl0kk77K
85GLzJFdcQMEVrpBvDrXD1C3vcFiOstl+OwXr0y4hJU/hww1OMZUXN4CxBfEHVj9
v+tEuveZRVyy5hY+hkXgjH3nDf14ucBRNH+FxJSyELaqMfU3QJTJnfDNSm8zL8Z2
3DLGIIz2k8XY3gdUtYLgr/HMK+/Jpx7OiT2l7ui4hKyHcQkvT7pz7e0sG8u4X9MX
dRCuIpbQPX0o2qB02iNt1pqAtDWKPIMVpMCIunt/Bg9qpYiNPyMz0yIPlFprw/+0
eZSqa+NNXA1t4UcYD3vPQ+BAqxSXndoD3fmT0J+9NJGot4STF69ag4AEWHT+G4F3
rLJeVqv4DSjCOldNVlZ2Dw+2Lfsz71ztx8eN2pl0HvJoATLZfgrhBeCICwEubLJf
jNY5K0p357NuQZnk6rVReM/alI296k6y1o4s29EbXcf7v87/MlU0HJCyy5uuAiaB
et7PsmxcY8cTHeer3AKxQsVE413t34qaH7IAX0MAvzfOLLeYCNTxvzv/M2iU6BG2
y/wdOwp1GTZ7XnpC2Ruto06Spr5suxnvM3MzzJFGsMJEv+sWxdAcniOx04yCP7PU
ofOzkk7nBGX+Jtuz+KyElerpR+ntlhGLBOIZkNjDac0a17CW7v3iTEaMeoeJs08p
11B4UzbJKjWADp2AvnOWHv9Q26xK4Y8DAG7iNOSpkcWxgwItzPxweNfvfoLkJexP
7G6TKk2/3nfRYF/ouA0WI0qt5THeuJcHxpRc0ClzE29KU9R2ZcWDr91IBqfCRi3n
SLOyaEq8WUdpF/L+85LaK2n6Hr4B7psnO5upzCM0ZpWbonpYS9kyvY4zGjVPJQ3c
HZ2Unud+KkNukfEpgQ8FIkjlVQW4Sdx5DuP+3aOcBakbMmhu5PQjkWE/0gsQ4GR4
DgVeO6MHx+JsKjB1qdfuKg9LF3yEV5JAChyQOpC6U2kA/YwYzHfg5CHSuZ78cQIe
coiaaN4DalnumqI6ZrTmTq4vqENcuu5vZgCUuEhOmW9X5mttLWrHTqazbNftEXLj
EBxtvLdHMBjb3kIRSSNVFZpiUviMEZaJ7lkj/Uq6/Cg6GIjfU5/cdZlXVvux4rK6
Frx+SF2GlFZ2y/NjEWAbU+IW9v2CIo11d9AzTJYOAxDRLnKJT71VSidIV0DsbW6h
wn/rbb0G0cDfg9kOuhnyDneZ9rb07kq0AJKPiA0R7S1f488CI7b4mxgo75orELgP
xhnlA4eZI71C7ih0qET2KaOmDIczFZ1YRHql6Ogs59tOjzwwLi9wmw19QwRPyCVK
L3D+aNh+ctNqBiDrd3h+OUSbCg56K1C+MF4VgSLcyPJprLGcbCMTenZlYRL4Mfij
xr+m+1+3nmv1jpqRuAO5kXUuHoCO/TgL1x38mccHL2FZaeC1bHfa++lLdxi2fBTv
QIOWNAfKl6NGeKgnMq4reHhwiNBFA0ZqZUrn/E/sQ5BoTBQ+BwYsY/HA7Bv3hOl2
BQJ1hCj+A6fa2NCFXhPSjMNp/hnHLZfn+wGDbZDA8mZK9/7ImCDt0YPix5ZX5pbT
diyxUcD7wc+Nai4ExwT4WrOAcbW+65eBVryayhz04e9xoOak6d7HSLqQkl6+Iyun
fKlAgUzK8IBd7Ia0UlBJ3og+NRAw4FWWWkfxnIvC3BVhKdEhGj/rP+yYxCgbM5pz
DAuL+W2MckRikdVjZKY/PVYtm9b/zWjFahZYPXNWWIkjZWHQTEteFq6X4T/0f6Ig
XPGuwcEx9zjOk3QPAFXlPWQuoCRBHzQqRX9tWVksqbD5EL8FUIJWcqnE5uAudy9a
I7XqlMZg3rNpHDdXA3E7SycNaTILgpl9uEurtyn2oBBQ+PcwwU9+aB+eA7dTqn9J
BRkdfsKqsd0IygrLjsg5gl1IjUBZ1vk7ZShUrz4Uz7s/iMmHaA9+m6QVhRUgRwv/
r8HZCfbaz/gnyoEsze9GWs8Z0zVCUW2I+/ObjTwSxKaLvnhI686HaX6FeB3mLhL+
lFowS87JRgefDvorNsLUkpqDdGXfybd+sdzUURLv29J0cULo60guR8qsp1IN6wxU
1CjzFzRx3mFDqTMdqyPcTjc3CiKlQhC/rxIvWSl9Dj7SOJ9FBTT/aPgRTixbBGFl
Cg2uKDZF6NZKZl/6CPqXjJBsTtQpLG7m7EiDz5Vy8lGczb+PXct237ikZ22lbZWd
TcbSi5VKgVhdGiQ1ol7umha2hYGB6SD+R+PMV5TNiTNcQ+fxiZLkJI+BouSAaqa6
7bXDI5evg27KNXVlEuvw+WpKngUlFUjmidWT9x3h4I+D1LydsqoGKKahfM5ts1/h
7z/JlidI7+9m0zfaU1SWxaAl+YeSSEBwxwS9+0EGiyPwuv5UBUJyD6SW5VpewHMz
CWHuEX1hxryLb78I0mzkMrvl5LGw28NX3KCS93iwBkohEYz2QNEFWVWMR9qA3qzG
UVfi7lTqJzWm2hyGZLVn0tNMlgZ+p94CWp0rgPbl8Z0L2J2x6N54mOuQI/ypUtLc
WFYE8OeqXB8QQohKbYylf83gSoSmP9ArAXASiYE0cbLNWadqGOKCSi02Owt/t4/v
HqSG/LkRXL3gfogdExuh4H6yPOvXx7dyxALJklUvU+bCN3mxJ/g9DbDRb0+Ayj45
aAf6QeaNvsxpR4E0Lr/idF6nNj8oz0DJTvYFOD5D9Yf+lrhDuu0EbUS5kUxRhBFD
I+FGQizJ3+p7pNqxNTZPuDsTXdeqat4KbNKP+aWidT+VgcSB/kiWxfsr7T6BHprZ
FsONMXGXfd7eCo5el2XhS3b50fitKqXB5awi29vUZbrIDRn23Cjrah9zyWEMJOYQ
HF6aEZIj+mTKIprTllUzE29dgbYZdNEsxYUfbyS4v4x4LgCadkEeejHFGVgfPppY
aq1nrjtKJAx0NEmygugLQrthhHr/Y01kdReMU58OY6JWROqpLZCybdihle9OS++n
u+orWgiv/+YPDucy/M0Je//Nz5yEvARz7ZFM/wOnYX3/nNOUtrW0MEVaFU5rCoPN
9TzXLhrYV5fBBJ7M1jH05jaEsh7tqHX58UjT0JvLZ/eg7BwZhpBuIoPe/lgm4ggK
KJocHDTfWAVGxqgWBTI1lgfkFV62uwPMCMx3020UWJ6oGw51QWmqQGcgyGwLy1xQ
iZMkAlZwMIef6h1owXelDozLcAW9lWaXz37454Mgk9bUg/7IgawDtLGJgSPsjNUc
ZLdapO5ez57GtHIGvgzYoI/dhaw9acJD8iI6TPDfW4R7KN7Y9YhA9FXLWVFtHYzu
kzYunE2wfblRH0p6g+SGQciIKg+qH1yOW8qmeOGK1+VGgLGQj6VtdNGGRG72DPza
BLxNMbBW1uJLStocnTD4DvQUFVX+2QrO0XXRSlnd3mi4Zk52HQKEsf11to2UwGa9
B8UC5etj07lDZQ76WHStvR8IBwRJVJbSorOfuzpHweNb7waF/lgsX7vIwWB8tDl1
Eo5Qheihv5KgGHzHGiwNVqVBwGFa5jeJHVBHAc5/18mZya+zO/JjgC9tA/uhoqZP
LXpqvgBWBtnafjn85EOU85cnim5ZXmQADCfcq2U3c0Qk/FYecHrEfXJyR81jDe7O
2YrBnT/pwAwC4eqOaRcPzissZRAkWwWzaK01+j/Hl5lNaoipIUw0XZBAtJd5VAYd
LzZs1OJu+L7zKUpCE+BpXRbyEdO4GwWI3m7cZlBinLPNRjYm96poTRQTlBhrMthx
ECE3V7vWje5GBng0z2yPMYJQcZjVuoglMViy1thIaY/dvGtMcd3pB+BftWErg6Nq
kvAnfGwdRyqTXAfAudtoeNQG8NG0B2gBmNTJ33WFDfs9Yrpya2pA/IPilGinujxf
t9EG6BEmsvHubHWAhnPFbVcEVzugLkyePAcuEkqBZDi2ys4FJHL/GI8oQj7jCj9H
zqPnBcTy/bM03qaNUlcNqqsfiyazFmR1o3oFZVnZk/f0k671UJAzfg+wef2SFkJP
hagXsp38ukmbEM2NC3Li772Qr3dXuTnl0UpRB/mqy6/x49SfI49opCnJw0OuBzql
bTnDaF3hEme6sEl2lHOqe4BGkrwR8YwkrOxVSfHPd9FtKqt0pKzT7UqlriaRp1kj
NM6XbfjQFrSbP1l8KlgjwBv0gyOIxr3ijTZgGt5ltgDgfOhAO9bHMF45LOVkQ/Re
3T2ahBwiZ+t0DOQxEKt9dvu+Q84Cdqml9qnjx+0yb4PjZ3o/55gXyXeA5YeZZRCd
XNditwtU3FTO1OIOrRtmVIE4Jxqv7+NRi49tYNt/fndlh1Hs/dEBXArnX+Bq+8zs
cXeCkLrkt9PzsdITG/+xrQLEGxfjnR/olA2Bzy5UuyCe1UU1rZ041CbTZmlaR6Be
mA2XTBTfm8QaQvn4+CAdv6m/d+lYS3O00TftGaUXC+o8pt6YXdVEzrO6uRsevQsl
moJ2xAwp+JQ6ys2RQpngya3Mm10lqn5TY5Wb/hso7bRq6f0r1rsCM8W5R4tbCRxK
7G+IYpHtkspUF9rqr7eISJPl4D8smIjqstxWVzjymoD6lcGcIsNW9rR9U8SO+59Z
VyKe6XWvkrCHju1qBGALibBhiiuRukj9iMlErw6onLX667iK65YavxnwU7q0x6dy
GjkuXyEiofG4cqbCrk5P6I/xCtF/iiYDkAINMs+dmFnLf9pgL+yqgBmO29RswDDL
WxTLMGLjUjl/A3Vcxw7NvpmQfdHgWIJQ6Q/GLUn7GC8715KnhHmXHJzexLWNSwx0
MGjRP5iXYt8tLgFO6hjY6Qu0tdrm0MhgGbuGbGdGFKbRCZLMC2wwc4c367CwmvfA
3C+ZmQlf5X+ZJZXSkCf/n747MWTG/d16zVZWsaE9Lt7QSbOm5U2wob+SmJx3ax9o
nkAdVDQFCaWRBSxTsROr6ZUqOd+YqmzD5TyL28w+dALbVzP6/z8IKzjQ08KIaa72
i8YvfSK0rkmqvJlBuK3WEN3htwnmDYIvRYdQq4HL9Ap2Ai3s2zTV5XGcFB+N0/Ui
V+Lr9pTiWjWnUnglDpjSzYkjMF4nRfauJ/cMq76ht2jlkUEBlRB5sN+TX4hGoy4i
9QsmrFKbHnkNhI3CmpbSg5+usmvaEi6Hm78Hlmgfhb4F/cK8WncDMrXr3yga3N54
RAJOXwEgO0ucQUwAg56Z3secfBYyiak6+jYVNUn5yr01D4jFWVkOYM0OK4DLq2KQ
IHVDNtgMG1yM+2g5xqkPCbacmKP7x+NzPrQFWWs9sg1rMt1N7e6hXzDIcHFfEHQ5
tLPL34O8sQ4H1LTWdE33h/7Hw3G4QNEboJaL2l/NtZSZF8ZEAwhkLMxXFOXh4whY
FWHM8l0UOqsM3sVeVBGaC4HZOxfBc67ESrwNLHfZx4hM5scaSRUQ7OnsiscO7Mb+
WsE5kgpquzEljYGF9u9erBuV4LSAa4CsZhWhxu/ioz5PQVp1uuXGwyFgk5S2oVgA
nwzF2Q6VSvVWHRsBFYZmYW3KbZTZ3jI1hM8EV5kM6+SfS20B+wft8OllwQ7nJMb3
0XpHhY6F+iz5iRYUep2G8ejLZgk9vnshmfktSbfVYdnIsoy60qptCmsYRCZaYRM/
J71sk+Mk2KR5DjOXKnh5q3RM47nL0G4DjSUNHjFR5MXtYhXoBG6uAS02vty3aSdk
QXPHCZ7EauH+e8oB7UM3T87JlX4rne4bOHVSkf8vm5kPLMPMpLeI4pexDldmImpY
i52RHEnGP5EejO9au3y0FpcsXcMwHVU+AKR+dhWucUT4amiYfq2aGR9wZWK+pc5V
ms+wSgoH00mSwxd5f+Zcm+8tjcEMYkS/mhGeb8c8lxIMH0ZWUuDtRCJddy2nijt3
ip/NlAAcCKJRmCcFE6wihr87AuYsqc/7Va+kczp/ocZ38f88ctG/AhUGzxYfxVxk
be1asKVaEfTaen+3CjjjwXmXkcZtUdcOXvwTDtF1NWZbAey2wgfQ6Z5Z0dTY2rvS
34JQRbYAyEWvketcsNp6E7CLrlFDRyY6RkDIojntFNdPzFgYvWhSqeJ1+m9+96TD
TJPef+j0jS39hWlHaxd0x9biRikN+0hJtJqT7OxYyvtUakNIdmQQPrHOp1dVw4tw
06CSe18rupEmMGVuHHwpv438YmcRimnBpZFSmrM0bm3h6Y87mo4Hh4ZLbEkcDN47
tICv7XiNJzJDec03yWJJFke8NEA6xkXyz0YYd6t++nJgEGuDNHoO6gGQs3RLe8z/
+p3FIwtEWbEM3XO1zfLtyChrXDgovS+NayqLbh4E90ReXApIFMLfclv+ENkTuZGP
vcUHRR8+9ME21sdk+288aQMqwtUoU1iMtphwQ7cXoDkc1z3qUXkLz55H9jsaVhQ8
BUfbejGmq6S95Zj5O0IN4KgVzwreO+3ZJ54FlUrTjJXYTs+Oq7FcbizEnrAYgLez
nATK4Q1p1nnSnOstWAc0qHdNfyQQX5pJjEY/tD2oNM05qHNq/7Xs0yuQIPO9S/fy
KuDpdSJv4kbIxQm88U9i62/VDGJuijbx0DR4lqmq8roFvijQSDrw6rQH89RPH7PW
OA0GUwWcrR/56lvrNalGp/9wApl1t5Hu0csfq7+yQHxfn5kE9+pM05+f0dqwEIEb
2AUbdhLQz1zPyZYRP3mst77UMYL/82/vi1/b0VJBO8S1my8HurLFHOh/BQsakjs0
uY/x+iY5gvSMmFItkAoQ54bFXUeT1hvPJu7c8PPZUPUWjvsF8WFsjS9tqaEGBy99
Cln2knGZG+7ftwXksoV/iFC/7IY9hsOvHgC2Bz0Dba+WBoyt63nNtbIK8nejw8fG
yFEGLi8wCV0+bUXkoqFJKPw6T/bi0fMeFHTc1vVUdkvGtsTDE/d4xeIk9g/reSYV
fNvl+XHkV+mZi3o4MEu1hjCLoHO5S6hAV96PIU+CD6StC7vucIIV5ghpiGMqW3SS
EKy/9VUBg9y9K3TIqO4nPpjuOqLSkwED9JrIqU9IP8D6bdw5QyH1nt3XSSw1YIUy
GQSk0IbsXRl2tJDjidjaf+w0XiFz/fmPY17YG/sxJZ79pTK+ouBEyhwMWR5Uvn3o
rmhxEymmbPLVZkZKwdtmTxYAcx+3qFX8HzC0OQHXRVYAq7vtT7qE8LHtA0XyFfjQ
paRI150QWIZ4eT/ezwqUC+wNjvxWN111HgdPo3fFtriGcnWIAJslC8VW6QtRwZwi
x6IDboEDigiXqxDyu7SfmobGm84gMfnc7mc/OYsTKIHC5JLuHL03j7zvdI82NwOF
UK9CrkcECRHmL3HLgJuumnhd5X63wwtYROTVUmOyWEA/ziljOgVWoI19qDzKOV/o
4yarK5rYsim10xseIMreqA0qMhMyHzaqnn4dMeDP780bLcnGKThEBpnzsRYhWv9O
D1HlLH60KlzWOsf5hE4oUMMzEga4YtH/MFpiUOVoVjJhASajqQS3EKPQaR9mGG7B
BzbBtgjGOQsM+fu46e95uG/rEuT/bp6JNG4O3ZtOADffZEFRSs8mv5qdfNiYuM13
hwz9tirONPSNhJoY9wyWykWzuy6jADYRBgHaS7Wdk7GTt6RTvpzzd6SO1HbuEzT7
A5cjWTilMk7wiP7LG7uPavYeaIOWRHm582Z3hMvq6UC+jKO11Dou+uDANbdKlwX3
81UlRMu0M8b6GLCsCdHuJQHHE+2V/qDMR4vkQTecVaKSFxJNdbZtOAcegjFpS8z8
FO3ObIqwTYx5tsfdxZfoHEQOq3AqnisxW+DiCFYyhE3FSWmsIaUlyl0f3NOVi7uN
zvsdwZPhHCX/mdO7iqLbmOFs+KvO4lTVwWOY+4ZcyY9yTOcHxJ8jU5QealTkc1dE
D2xxABqXQNptRC6O8HVI6Praz6yKT2MrLvtik/SG6LDFnzFqceODPx2TgvTn99wu
9ldeX2btCaxq+G7W1psE5ut97hiZzimaAIMVnku6nXIFgEGfijXlnGB2UTHD2S5e
3/GRLRzDif/6tHa4z+MjMLOIY2iQXDdZaNYxWNEXDqYfrA15nclGLjdy+Pna3afv
Y3UrXffMXqo4IxcMGcUZ/c12MdA8b1BoC3A/YE5lQZ0BB1LOjEtrrpNmWO+2PV+d
l2UEwNoa1mHU+zHs6A4CPgvVjfPwFZ57x0j5zxHFfylm70hJFKTMiwiXn+5VeH5g
ZRkYido/SChG2mduJba68cbV7cSEUow1/+kXVR1f5RfUV22YEPninaRfNq/4C+Ts
b5P8M+DUo8agcC70C3sS9GXFykFRitFvmvkOwBMAhILUJrrW1uc8pXg4+iFc8kP2
6QUG036B4zvs0Z1YW/sTQt5y/23IVFdNwPOEGIPFg7OxzSxT8b3SQsMGOMDitzxm
k3AUZPyCZAYaxaxSJPgEpUXwNC2zLOuLSLKy3vCaJnDL5Rpddb8Tl2XHWrJY2Ean
aQ2z87gc9ruEPX8L/TbS1ibpwxDUZlHQaHbinOb3GJMj01mEB0f2P13hS0zhrCoi
qSc3j1MixdG2z1T7U1nnJUewsk7BEMBuGlKOPlYXUT4FrEegBp+iZNoTlw/1jNTj
zqRXHlhus+hlGf2XH43C2veP0v1yasFK2q/nWq+RNEVHTsZ+xDTdZ7v65c2czMhi
RJW4tF7WG29P0GTQvWOJcN7ZVvujcsH8rpkwdQAlZKpGwIq8uoxHvTeBGvdR8g56
I6TDtr/AU3hEKSqtJSvRxl/DUQCLrFJAzPb0TCmoDpZHiq2BFmTHtlxWRPkOSWyn
KZcPNRsN852DeGN1JZTtMl5TkJkwYLKrWfa05D8P/cyRfgXYgqC0g5EgxSbiIkWI
TrelENYJ0VAXHRgchEgsIt+QErA/VRvgVqGUPUfFHC4RognYaAOeN+iCLBJ3yxFx
fuzArDOeePVodzKEgTzrIC1f75ISjPqb9ZnB/yIRMUkR59+ltTytQi+n077uUSI9
pfHdVJH/tMmGU/v2+dGSflhvy0FWSPGEZHO74eHI0/Yx7Ius7jBLtCIH8M8Px3Rr
DfOF6Mj5DPWsV8A0iMqCK4boo0RFh2ot1vEgkiOHSkNKkPKdzApvcCKFc67Cc/zo
ZlVTapsQcsthoyXncaDc4xv97UhupJ4JuBYBAVXL+Nu98+ESrUpB/HH/ZTGdeBqy
3lpzsVrRYo0c5Qc6q3F4u1u3LZTI0tBbl64WXcTsRaZqvwCJ2ZW+YxtUQEWOI1Cs
AszYx1ck/JPs7biPJaa1JQLvoVUrHmTrulB67QcRxCGpWSxMFB41a/cwURtwMDzx
XoScAGVZhe2thdKjbbveY58UNCzX1e5H+oa2zW5rLRCjdbDrZM6c8FsmTjRaR/LQ
EkOHVjZUw0UO6liDdcG5qWkUD+wPazThqOPGqR3q32bqth79BNIU6lXOMeMs+bcn
GWl7M5pp5p/t7hmnkJCvxtt2HSQ5qPakzeVjF3edaN3rokXgOwpIYZPIYSeQXUui
NweLa97sLgPmgtXSAffPcDqMsNoGk+exPxRoojwH2ZM54COn54t85AIvkKcV3mV9
QLQLB+gJKin6o7Yj40Sw22lErn4nAUz7577vnlbzF1TJ2JjFN9dk7dxFLUuPASHo
bxeeIB/9CX083HP8j0cyxTH71lXZ6zKB4bO8MOtD8K7s/WQtkuFPUz6xPiTw0U9v
Vxqn4fLYalF5NS5OPNgFYTX2lKro+q3TVXRCi9DzCo5K087K2eiQx4EROwI9qfdJ
W+6Ilhaic7uzIMFaIJmq+ON/lmg65Gzk+YSuvXlTCfkfQV3imrjFF8+6nyGikLMY
yzwhphwOsc7DW8/TC9+AwPxGFq2+kr6I9joM52g9O/YNuZwSVfO29Usni/kkYuQ7
Ms2ZdOivUm8Q+2Q47i9mskbQxPrS3gXvh5vy8LsZUq6RfpgIZ+WNQwxw3JdZHTrx
AgGj4LIac1n3v7gBDe5ZR5yarIeVwyivSuDU4iS5Wx4cc9TCigKDlzF9YRmequVs
cCQX6w8m2sl5gYmP/5tJ0EjzIu5+exhpA9oF7X1upvOO/ZBZZ1+Nf9yvWQDCZGqw
uje/ZiK3vf3x+qcbcadxlyVwS5+ySH98alG2V0kXUMcX70HlyZ50kLflsPvMqpME
rwmTCFyfM4F7iQYFVd7hU4in3aZasz+xZMniO2Ei1dyrqG8XuavgZaotrWCOkSp1
l0klq7sRqFNnpbVdeyac/zO+ZCxkpvz3QBqs2JaMFH6rbcXaoZFCb+cbDVzgAgFR
6AcKHKlUsAxWKGqyUAKoVFPqcvJk0sYoFUeTMrGQIOE+1j81tkunKGIvcrJ+5BHc
FfxW4MGXMD4MNvovGoskyc9uAEkxSfbgg5xCqA+HBratgzNz06WPAaxwxMPeYj+A
hP20iR++SxE/zKauRVpSfvuz46iTm5O90Em58eE40UzJxE+p1CLL57Mlvl+Jdjaj
PyeGO2Qs51P+LUGItX0/0c5uimzcT5ht4VMfOMTCpnBzQyEmcrfz7LmucPFz13Wf
bk6obSFrPkOIIdPhbUczf3/QPVabduobHzZfQY7m697ya2ALSXJ114W5WXflxgnW
cFuFwiGWjvloaXASKG94FoW8x6OHq4wjdWsxb+Vc6/HnteN5FPE7w0DRVWfXJwgV
n1jnjzpR2AKS7EkFZyiVtkOvZycxqkPKWHxfs0K5CeRW3UheuJ2gTsywGcL+4Pkj
qk32JBGR9dVx3g0OiZeqYIidxjrBly5BRs3yzq9wePWFVPq0vKwNzrFVx0gXXU6z
ZyuDSeQLUZxWrG5LFvjX+bKNuHsz4/DkK3lKbUIGabVQdA/TD/nwV+ohMvQ1K340
CMtXYiDBbZ0DCk/oZPwXaO2Sp6b9r0TqWDyGciFSIszcU7knPVQ0ksDsPmAvu+sz
08a3boH0XHC1Izfw50gxlOb3VbNpjxCSNVByXNrD98HveYc7Zh5zRgrXlhr4Cxic
xp/qm+hDAqfSuQuFpECSVaf5hUcFO7GHx6aiFEpCYXMm/lPoxGSB9BWtRMpGGH3Y
g0GZwBgoAZ5aBMx+H67T5IrWtuRhacGTNeJ4pmt3oCp649q/cpe/o2PEu2KAvQdA
N4NhlAEYXTvt2w4FqhLjuA/7oR/wxBjeJUq5MYXYPNRWjOFKLOUjj+Vj0k+82mZC
cSrzZOzX5E2XUXB/w+PGX7MBGMZtu+UtLeW82TvUJ7bNk+o7hGbXoUVApArNqNLa
irBnlEJZKYOOTiCvrHZujPKGY72lDZ53r9W8ir/QNPwdF7bZFRXiP66FHyktRY4U
td9EKzbCEwPMgBiNuu4H5bE7citndVW/FZziwqJkddtMc14LDn++/GVi5GhRD1VQ
Z+wQT4+idkVnW2V8db6+FALpMzt4OIkwM95/YBOpJHxAuKE6qFWL9Q3WYWM7zBIn
jP4j5rP+CgNRNLorrUO/GpW33+mGSeIilh/Z4bR+U4G0L2hqMR/AXRn9oC3eOJtn
dE2aFwvOaoqzDNk/QkTq/PHDd5U9YEV9sDV5jEefci5ArxygIt1BsEufART5pOnb
UBGc1u7Kl6DQJOm3zLmAr4ZLKmwT+keWfgYmiELz4cav5tHhATw0nDQp+TGUlTHZ
YoJzZzZaQxZXDMqknuXj+JOvHwAlMN/a2lACcWnIh0Yb7CDteEAtlUT+qDEbksz2
FZcxabeyRdByZXA0UimgMfN2jYie5ddtTbL8x/rHXHTBnwZLtrBn7hLoUbhkWztu
kHEqa6BfnxKBYPn7AQTi2mUSDlnK/vq8DiSqE+g0lmcibczA69GRKsDFxrKEr8B6
oeNjzwrLx447Cre8ODW0rgwaxxyagh14MaehbeCrJ6PzJopowc0HDRqkHtONOn/E
8HU73f7A87usGF9IOAoiI66hGgdXS3xyUqE9v28EF4D0g9dBQ2bafD8xozAecOml
2ZO8n0UF9c8sNwTQdvE+CyLhwy3bSQaNioeeTcY7KK3I14XdLntNzr8bnlzBb8VC
rNgiIW2/3E+O68F72QFzSgU0CPMiIGeCi1o/ohFVPTclAm9KwYpGvHwVggphiEVS
hVgpnaneX5ZYW23q6XJ3uM+TSPbchmWAEyu0VR/IRWu05fra+gUFN3grr54if8g7
7WNWC735jT/UKUPlvMlNsw2f2eMkEEO3PnEunVPrJdt0wt3QPhm1qYJWi6M7iII4
PT3HrKEREsa6r/fXDu/kfyFb8WUatClCNA6BPWA85wiCVLEhfta0vV+mpzdngNQz
uWcDOTUTTqkuO/sT6ZRK6Ee7GybblhIhsj3Fe7SmUpawgOBh1SZnlpEckxTv4iU3
xXkiCdJRgmTtrDXG5AhsGRosLVObaqQ6yuiGMxQDp5RD+TTaH0ykDKL+6aiK5Kh5
KZmKJA1P62y90UHAfxf/roBvp3UmEYQGTFum4IvpKHDe5zLBQzQyahQVrfnmFmVE
ThK465O2/CG1nqPiJRjcSGCPNfcMu+NMrXHg6/phkYHxjMVLJqGICZhKOmVNfKH6
O8+Y0sJR9tD2KF3bTVAuwjpAZH81SoDVqU2sbSABRPs3+Gao4yKxw21i8vlP+j64
hh1b5WpafxKb9UZuX1fX9xkiUxh/2re+4j72Q/imj56HR7pNt2F9OdS7Dypq7i9X
CVtrV4j4gc3LDpy/EKVZic4S9uuqR++QCWgYBrBpkjpR25pvDflr2cg/x8PltTgz
UYxudaaLLst7lx89AW2yBQUJKmojfzZDa7so6foy2j/VXMttagdB46abbZISqiLH
sJd8QrrsX1W3lwkPZXnEJ7oxDqcibspwm06x5wu/WFNSWAvm+0F5tqlGcGxHvD1a
+TizM06ddhpzR9BnHl5E4lqPsMDshZP5F94h0h9gXWuV7sOHX6pnqoz+VhERrFMX
0zXlc4xgSu4DgO6wXaGZk2IWjWsLrkus+qtIMHgI/5oKLDvXd1sGXeAfg68HV/ER
8/rANvrgGtCP4HLQVs9e1NM+spJAJJVKRrW4ynpFgFByi0zZmK8cqJZK55VVO0as
4NS1S807zmyMIwn3pF/++Db9vKKn8rhX8lvOnsWoQU3mcyrbCFauwqWj4/QGViR/
0FZ4SehNt5f6Fab+oSXU/NNzYO+Fb/9h2oBHOumRPuBWpvAKT14yUkRLOSEFMg5j
4HDQ5poxxOhWBm/2CwNVP5siYscwNJoXaCUCaCD/4hpp/i8QbpxGsU3VfvacYFF0
nYNfVpEOJNFZUJuzCVr9cZK8UWYy4gykuBgAi/8CcyF7WGcW7KBeIqGH6ukeZerW
VWlu3YRZ09QH1EEBGp4Q0be/Ee/SvITBe5ZlG5+A+QHUHm4Cyg7IVUSZ/MrRVZh1
xtpE7E1PgcZFP9cDTz4xABmcL0M4ToBI9ef8ZH+1Mr+MUMKZ84Ql9FTvfShL/iSc
iSqeKe4HYjww+tpG3yUheFpuzUAyo2xUAntTPhdjcf18tavSKTfFCj2b1arUDjVH
ZYrWXiuJL1DwR6OXtiEE6H848EtVh2Bc5mmAUF81zNkDtVTEiXxMIHOt+65uTt9R
ug/dlymT6U3wKl0ahlLYjdzN+bYUC5X2XgdTTWQK5SbLwH8PIIaJbvqAmut31y+5
tjy3lJmJuFbqafrget/x6sJuteP8UWqn2tgQZAiKIFPMuwKUFGjxCKqeZuRPZIqY
s3heVYbusia2GwSnDXuaQkTB/z0u6u19F6drA0o5vsrzhLJwF1Wtk9+prMzdWPmx
D+1qT6/VyWaK7kp82Lgoc2mozQyhrmiT53DNruPt5F/dNY9iKyREF274NfSffTdm
+PMJ//dSQm1UFl78GiX8aMFUynNT33NPUG6lgH4Ur/ucpIsyCJtpGKj9Y/nIcRtb
Z+iEQY1bAQBn0cbhXajd3nJDcLJU9FTjVYjuS86JoEj4+PwINJlIVQJ8aJrnWDxy
4AJb0UdfOd/mW+dB8SQ0Ta4vSqo33bdy1u1iMIfb1HI6n90Z4AG+QhdYGHcxjdKs
DX8vylpEUxKNolQDzi6nt7UojSTkdajfzakXk09Yzig4DjJmZm9k2Q8WPdO93Y0v
Z/HFl7WcUr4+tDoy4tgCsqth8AU1XV7eUBMT3YJKgMegtilMumy8w9I4+kvdCEDn
pVP269SSQyia8hM6qzWc535m0jqRel/pB+ooh6WJqj9mzjowQhr6eTanZb+cC3XK
P2UMgc6m5rJpHp29DPcRHQvrhfNo6HX8BopL0xjbYroJWxwVtsfZy9Ti0BfgXK+D
6d6GPjwFxFQYDCp9eY/1xuKgi6g0U6qGAINbv3UYCg3XsCtrFlQUi/ykHwOKZEV/
gGUZQiFPdobCPptbd7oUiCy0V4TUkbck0pFcwn/KwgSvxHn3dJ1thyvFJWHnEKIi
kQvG3ptp7CNypZy4ikaNnL4BQC4TjclfOwiCwd23omQetJiKObB7YNcE5hdjsVOl
Q0c+/qrlCnXiN8p2oa4t5361904Jzc4Q7VUBUE2940kNKb+6TKex1YcB0pN4IwAF
dN6bZ3h49G1Wcr5B+XrEbbOV3nFF0b9eXppbtuaBLmvEanSmMtf0beSuyI3QEtot
SNUdxV+3dmB8RgSSw2KBmPq+E889LzuP4j0ijyEq8Irfv4oLoD1+8nCradGUi1nN
fGpjN8/jRb24nTzLHDK6UuRg5B03Rnb7Ai3C3iZts2IVW0GCCgge/D/kA86XpSw0
wk0F66SD8KUNth5CEOfuqK7Qdaxm4bS+6TkymV/DROtSCb0DzdwfNhyLeKyYdnGb
03bvNR2He3ubBE8ce/G8iCLtAkLMzC3plQ4458s2IIBJg5NA7JHVAYLzuMMRNDKY
NU7+aNBWhmInZ/uLjbKw9l8q8yRRi/vDeZAGz8HE951dxfY/0pLc3y0Y38Bx8NXZ
sP/XE0BqShWbQct4mYQ3M7mb8jRzalBWthvtJwZ4N/P9lwnR424ZrSPMCYUg6KYu
Dhd1450G62ya/wfdndnciMTPIJMmfLMB3ny13amkVnVIA+bQq6SYhT5uHW5608w5
FBuULFETBKoCAFW1bTprNumATIyCJTcT3OWvDWZa3JpbwaUaTly9Tp+QWIFYpWDb
uQxMogSo3vaQmlJX7VtD/Tjxan4bSmtyXaP/yAjL68tNUrtMdDSnKtIs36RU8UAo
aqfG2ZCYtl0WXDgCTVWirUuaFnhxIeELeSQihSIF6PTfnQWrCgW6ySWWlaUQHv+l
a6C9YDMx8KHWp/S6a5O0EDBlFdWXHeh79gLdgdHkIp/mmDy9vVoSh0GNziWMsKXV
iOjXGvbyScrZ9ViZVQLNdAqh09JS/nVtyGr3K6YcxQv+mosQPpJluPllEy/4JDac
t5BedErs4uuU+NCjKQpWhj5wrWYlcN7+vDLhlm7mzRmb/2EesHMpx/xOGc45HAhW
G1uUNcOZBQvrGwDLNWyDHXsffCkOpRip6jjtm3ZJgGG+D9lovdwx630AZXQfu2v9
xs+LW9pKmDnXH1yaefEqk9kim5HxSZWklHQQTL12dhqcuLaHRZzib7nA3Ea0GvDH
MsNkU9GIzH5JEPimGdM2RF15tBb0oDKDoVoOPgskh8ZCxF3ZnSR0qXP5v8Ay33fT
UPiYpfFMPdrEp9WCjboVBCbQKjBFq2UxwEJbTRNBxvJfdv1FE3I+ANPXEc5pbzY1
h+JmSy+S66B5IzwCtvy9SMZr7MSUW7I8rXXPrv8AcI9scQC26B+okxPTULRtKUZy
LZeWFALAqLtUCOW80Gttocu5YrUGCm0umk3mGfh4QQ1Vfv838oDCod5d4ooRbLH3
xYE4z+TkyXTiAR1G+Wylgm1INl5410A5GVXdvGtpyeMzkzjFnoOnyMysiQiBgOII
9A7Ez1D6a6pq/vHr9OZFAqGkIWZrsuxb6HGm8DLPs9w5PBnOoNMVw2nsL1l3XzDE
lRDJhNAvKvhIYdk9P4m7U64lhSfQA9jCaQEpeWwffoxq/xbMD2VbBZTs0cjS9O4/
uIr0iqMtGPzkd7C2H5dr2L48U2XaIPMuvhSTeLoJknKfCXJwgIp6loE/2j4cojt0
x6K2Y+8wThae9GqSE7HK2ZXGAr5eV8WyUOJhH+r3cM2QFcknl1b70Dr3iAs1+AT0
VjQUyCZkEG9aR8oDGofrn0lUc7DELRCbFTg9doSuDyaJT1oLEEBJJa5ONKsNTker
c1aj2oisdUSp10UYD2hK7j1f1S/JlF+EWtd046f8scXMbMW02YUpDwXvMPu+EJOb
zErR4B7ooVZ6UOblUAGigOiBH4fn4BbPYg3nqnpGufIp7yw92vh0qxGshYX1LgNo
jDoUfeVuAfER8ECs2MKcNtZFq301hgaYqesW34fAm5GiGyO+FAsUjR1Ut8I3EIFT
RNqypxouxLe+gU8g8g/Uu0K5Iv0rDB1BMpsS4EOoEVB0ctiFHab4KHBInKlmEWwl
mFrRZlnBvB0ckJ9CgYDgchoR7uYY13qUtvkqKm9zbmfxq3gWvNjEznD42l4/bQhl
7BWoGFxJmfOAyDbgajuOePFpYOMOdzkdRC0p8MnXzFUmSZcaclo0DFF0xG1oq7IJ
f7Z+cNoMTpnXB6/KYK7+caAmUt2ia38135N/rkhMZ2cY4HPHjOIzXAxkbYB/mIhu
S1CXBf4I7sq+RhH7afN0NEJN1HJcyjQzxv1pB7rJMWLukkjW414/aXc/TAGxht1n
ihJRS5cNRwo/ho+I4Tuv6cU6aj2/mpUCuhMtMe4ezYPCgHY5eLXktaMrGNeXcmQq
FRDsjveD0+Izk7TK/7HjOgMy7eRP/mdTCMUHZNcq3Ybz6Ypk6RDbn1IbmP2fJnKd
lQBY+yUrpT+TrBTCEBra6hQaTag5d9gPVgkdp2qLR37bGC+dvPli1lBbWhn7qZRZ
rLgZiqtqW5ODKVt2cPVtkdB3J0P+ip+5TB/H4IXqxksx7jNEhoOvc2EU6CCofthm
L6NOxFaYnDOOX5XlTisHtf9wXlVXRQ2lYvEnEdN4tU16VXoj8EgxGR4JI4zfPmJk
WkJlNf7a/42AiKn9EUuRaCKAHB7D9y8lpib1p1Q+fwCHDTl4kpB/7cLTlxmWz5Q+
r9Km240fd+Wo1eXDw5t6c9OrGAf7GdORVR0uaE8OZ4bIVE4GvcyGD4Cx1xSGHcAn
d/A0/u38NSKnC5MB9kY2fA2AOHaQ337q00Kq/oteYpdz3CDb5nOQRovIOwdxURqi
vD3kkMZ6YO6EWWpSjnzdM2bitTME47IsGXyPq40AJm3155YiF8g2mSBYJ3vXS2dv
l8ikw6/Z0wHPY6gEjmSXgW8g6jBadA5R+kDzqixnSPbcQWSLCE+++5edo1cPTpVA
nji3W22IF34NBE+tqOZlPCc3a4PwxWF/lriM34cqV6qVCEYrFOa1F21PkPZFXQIr
NUKFd0gm1JooJ+NOUCluE5QT8CFBrIB6TSmrzZ9qxC5t+jp5mzfDTsQYVlInUd2y
LwebYQxz8crHBocjHzWOiF8JwqqGyn8sGkfHV1+hyZFAzFEj/ypx4CUrERacOn0T
4reaWmteKKsVCoQICtllANfkukQ4zF7IsRYR4tRVADnYDeEnLZZQdFUOJnd/hBwA
n+Rucp4uRl0XyMgei1Hz/7b288SjnAGVkV8asC7/dV81VUJxslPMIsiDdYESV/MU
eUU1QP1MN8HiR7lJhN+u5WtMfrR5/1RWaOc8K5msBGuWgHZW5wgBgULfIkTn4oUn
fvhqHn6BHWtI8OFGu/z8qVGm7kiMuB4n4tZJFy0xm0fNFiItLr5xfoHVSgLiAdE8
Bzl44sxmVnULrczn4Po+2eqbUleIzEm0W/wugDIV1D6XeSv4ZdjmdQBkb4pMuV7b
W4Q6OZ4oh6PQxxqgX5WtO1eplpgyJxKBd89rsH/n/ZtP6HQ3hl8IGrekn068tUgb
Bi7lXRMJzPHqW5PPfVn7V+J+rMScLqUzNvrj2iuAa6DVV5xl8KegqjMSzWpnF6ky
mD8vZn8c8sDNdPjdX0vBBsyVhblk3ZIs4nNPy8Cq2SKEdjTfig4OKl3BsYWWqwja
5+hnRupET53GIBY/Y1PonY5ChnB3jIqdcY/h5Rt/Z8x5ihedE1ASMiH7ezLs5ao3
Rwg+KNUnVMueaztqHYtVOtMicJsPi7fMXQ+0R9qGWicY0wYz+Jqy6KPasqWieru/
t3Q4pr0NevuQD9oeqG4zT2A3Ia9DUb6Xb6g+ZxCHTk4tknQS1tcuPzzF/zutbSLz
FTI7sPqILXyWSmv2eQAJOG6Q+DFPmUrIxbQQNkoJKmWgwLpiq8gYsNSVqvHE4eSr
kaU3NlFHP23g+8iuEo9zPt++jGdUUamWkPzSfG6lm+91M/4zQbDGmWOMpUuFika+
IT2qy9WoQrklRV4Uk2aHq48WGG4Z4HoNf0tDhusZDfbO1OvXpZQhQVtP0LpWG/i1
5XWpok1LqXHTQyFPfvUOqIzZbbD3FboSyFqah987ZKaJnm+dZy83yabLHRxLDcaa
Qu1gHNhkPGPSbc26dMl5qW3nkqw+LAxtGPZ/lIAlMLqOyQtuLycxDnmbnvV2vImg
xzLYZquZH/0fTPKdzNPogrDNzh6wSu7tjD4lcTg7Mq848hVUoPHBoXvYU+GXM/jK
reDNUP/Ct02edJlp3rg++LZ+1R4tToaAo2FR8aRmFyNxQ2enYs3VGiL0XwVYKFE9
PBwfLNXgtIT5Tmi8nTaxcOTghUN4pGGm5v3n8sZcQNP27gdC+kvFtnI/9AnR3owm
FNzOSBuviLQkK967xef8Y5ixI8ubxzCUsPp+Nudosm6AhtdEiqa+FCVQwqN5LH/H
T03oc0RSsYpnLavzopRIcqbxISXa/XPTqdVFZIjKSHumnAkGo2Q8A0N0DVtQgrgU
G05I7CVDSlI312/8IxA7RWY646r8MiCCGKTJXu5I3kNSiWWiRKn9arkfMviEq2Uz
ECr0r8q+4ZTSbVHgGYijVZH5PFwEJwgr84lblHxt9Prj+psUU0BQLdwm4UfLNwUU
QZLVNLsKbLG1GyvrzQcQUCu8AbWhJFmhbm6efTKaBLSzZQlW4JWLhvRGsNRh68sz
ap8c/4QXUDXAYvRxlcf38Zx8dwOFmZsmAHLfvEXakZYBxyTSOy69YjOe5Qqbyrbr
cBcHuEljTAWANa0bmwC3R2tGOB+y5kFKzbQLNYwxPu4YMi4Ifo2twLqj4FZ1HnTU
St0tB51Km92ysm4NZkSC0PzGiev3Bt1ETpdPZtmhCT1G7oxdDajKlmqaAddvmFfh
jQTroLGtTKdjtnOnxQEMZYKcfDR6UcyGLf2I0rsBLRh4hTMoL06EtCLvTsJMU8b/
EBBZSGi/jp+NyFTO67uFh503I3mjZlY7Xi/QCl1GwAtmIDum2k9uXcJBttxq6MtA
Al2GLW+yt0kucJVf11C7panZA8REiaL6woAi5f/qKXpLudtqNhN83Lz4dqdIavgx
L08zraud717wAzqfmN9KLUo9kkABKyerf3NKxiJdLhadcUUFN7Dx+zYGTjGFzS0e
Yq6JTwM6SvJmfle8ka7gZiR3cjUzC2RfYYfSMXYiTcMZbjeSlFw1XjtS/3pPt+aw
QzYp/JEQHiI0/bNZtLLbuSbhpDSbRD3gJzoLYc99CMudFd3i7BkEcf8pRvIqJ8Uq
Esw3gYiF8AO3oPrBeh+uVglTyfSBFRAT8VJGySAOnjw7wWaSk1yLWU2tLViwUvKl
/lTIIn3LY3gDt/vvLd/k62HiteDhQqcJlUcm0Szk5hFb4ZUb6dfx6tiBzwf5RncO
uFMDPnWT+A+nf5RtvE4fQppRnqIUiTulonVZD9NGpjJjf2b6/IOLvb0BhBu88L+R
x3NhlLxYQtgv2vT1bKgIhHDpxgsCUgeWpdqiewTS2OKW0PmX32sgfiZszeLz9jcs
O0aglKTatvTT1KNWApjoFiUoUGHvJd0SWWN9bwjeKy+hrLXpAJNiUQvSLg6mXCQl
/H/2IpO5GNrxSlv7/3WD07ZIOB7Lc2Qebkdi1FAnWGDbGjsbn7zX4DMiM0Rc/+Qu
7hSzyl3piY8gi+w8oE0pPYJSX5zT+DgTPfQ44Aij6vJPh77gQpGL+tul4W3zUGDc
2oWRbsHykHodW0ASJKh9NwjELcPAKfYQL272/m1v1lI+oJuAOmwaYTZNAFofCDI0
3qc2FbIawIlflQfPzZWXwFQ2S49U5WLAJwxzSfao76Xu3j9+hKAPcoqrWezgtOUK
B5/WnvjYIAK6Ze9BAAuqd4uRqir+Xm9pnZIAmdg6rQJDkISNFhsM55dvl5x38W67
7vpOMiop79sqYscfln782YdPnSOo22cK23pYFZhV4NnG46LGG+4PUuNYosK7zh9o
oOLuJ0iI9yzm5MK+FOm9kuDHg9+7ACwmdwvQkla9/HZIdUQlwPSC/cXHMjyKpxgE
c7dld3NWS7zohA3nVnVOEyqwcGjBxszwGg4b3/dEzpfKsltD92Z9w5ovM8J0cUj3
YBhLoAh3429rABi3vOleug6tMEYfpSHnH2cYoeR8BV7i8O8sqeFdC8bC6kg/sR5l
BDf4eVT7uqLLA3hV3zKceuURA2zpCWJ1h21Amu5y36CHk7EPQ2smdP6ss994tko8
8KcMDQnG5wi8oQEJuehxAEBXUv2dKfJgPgvG0Mg9kbBP/4e3f6F4JWOH8ttt7Jqo
sKlv6W6p64MlxyOPYm9ghAnS2gwW/sAu7915hiFieJwm1emYYjIQktHwu2uignOP
btfEAh+7L2wFsfeNADFzvbfepu0aPtvA4yGgLgqEf1V+Yi4N6bppsB1fj+q4wTgW
vjE53MqbdsYK6o7ma14wc54vrl7ize4HKEiALHVA6LKPqQWTEaFQgJKw7qX6eg9g
f3gOvWjsgjRlHoUt8XNNUIgaF5B1XS+XdNx24gi0tDu2qVGlAw7a0/LxhTq7kaFo
anQBOga9SChc3eVc4x7HxWf9pCqwlPLtb0nt1eyhhRPB66yEPfnkIWZyw+Y3NB0d
pVdJbOWdgVvdhhgUjUcRZLVVJ7OJ83wZPugCS2SrxFZU0GW3ByVfOK/fySRT6BB1
/loMRPzGPWVr+GRc92ydWdvwHn3X1efmX5uXf4r2ZE1nB8KWmP58z0YduIDyZ4CM
RRCvHi9STN65IIGwwuw/oIcoP0/J4jLz2HjNrjv3B+cAv1PGAEUu54hcgWqCNknS
KkxSIzQU9/54wngLBj804EVmFjgUmhrg4PuGhsGGuc9gANSLRYgVS9kVuuOQRy9N
md16Kmn/pEMTLiCc+uaeXPWIUwK5f2G37/vxTSV6cL3OwRhVj8qKA4mOVFv7eNCv
KDp6Q9LAKRW6qx7zpCpjR3FRoy8xva2c10yNfVYf5iHdDb11UOJrb9HaGv0fUPOm
hAuFL6AmHS0+mWDv+rEMUjPaJe0cGb6Vkln3jq1VRrLf4zobl1ZS960Xbs1Y2Hy+
q1t3+tRgCUXFBi0KzZvilT9XpA3amE7PnIZbpFs5Z8x/xSOJDzo8bgguaiVnqibD
Ro5HGt9DvyY4QjGR6Iu93NgIfUXsEPpR+1LLahJpep7uBNPpcpevOnql2VjuZnj0
5DVQBnQeqia4h2lbiivZkXFWnPM9Cn+xDQ1j4UkYk/EAzWb184K6bQ7qwdxBNegN
c5ML2j0gXlAsDSAGnAQPyJSgohL0liqf5weaA0qJdN/PQ9fekoy/BFpGzpaRCTus
ZePywfDcUAhWtU1+hovYS/dCYDEN/CWlZVSxtlg0ZDEFUQKQHqwmCePQdfumF5y4
axnGCChMGWEi6S/rf9jGRQcl8iXv4q9FrLHqqtltRkpvMZnpbbocYKvt9WeE90jB
nIbQqUKv1w4ntYAU2Oa+QgF9+jGreMenvMrUuW4abMnQ+fvtTwVQOkQzoirzKO+o
Dy7XWaKmySSKS8sBNf6NlDh15/Snd9POp4dzxLinCSs8cPc08M7XeTQWodW1Ih25
324tyYe5j8sC8EYALZMa+C5ri9/GM1fD4pf7hVGEfe5KANXt2Le0E6p94q0RIfhn
0N8XzLQqjbUHhMmteUHwajzkkxKPgTEp0ebaN24T5NPSh+zT58K2lXsJLv1x/rFt
qIwQd8dKYQCreN/DAVktOT4scxdXvDkDnRyjUKxbBMqnhmsUSSAXdFBhVPXKwMi3
9taoqQ9vwdsbZ/vBt1eKDaCumXyku8nUvEzxpVuqQOiC1tlA0GrhChdwTIgLvDv5
FqI8HMNekfqBgY+LGfcegLMMDv0PbjvLRbjfwSsvqCJ/+hvQzZUiFhti0H3hwfl9
pxZdn4XnJnrQ4RsTgou4zTmIfcVl8zS2Gm4j5BMP/GyN97O1tx+lWwB6wTaw22F8
ilSgDAnXcKxJWGn9188MNKSe39bikU5/5zPdwSK23QvcMexvqSM2wl3KbLcC46EC
H90zXhF47YR+pgediqYUNeuvxFu3Ola67h0xD5Z2Y5JQOiR32ilaOZGLFXHTmgjg
nLZ4hyASBeKQXTAbhOnoVaEDtq94/rd+VmIo+jKD0DHrEtiup1gThoOMKDN17wCO
+ZeByxwq1iyN2uxYk0fJQeyAoHwkvn88qVKgdTyGPadEDAYiSG5l9dGXn4x6WrM2
O4IVkZNDE/eexnbofAkAhQecq4mfmV6Q7amCBgrk+8SQFjPiciMCmQ6UTGVv1eqZ
zNThP485ytdzTuLmgGzG4P1ntlwe+Lt8OoMoqz3rRHq7vKlMLH7SHRl8VF4J14Za
b8PTf4rW3KYeir9Sbujjt2fvd/dAMVzEIaFglgG8vOMpueKQVxA6x/vcoxk6rg7v
lWMACiBIHI2yDPYSVZi2HKtblWAHmeWO2SUqP9bf4dME3QqLR/m6fMS1l+SdyJXK
m7QM82iCYEN3Cub1fb7tMTmeUjaChfY2UEpzlnzs1wLJyRVyvwk7/r0yS0FrZXy9
Ov0chraanZll3YkmltCgTdUYDVFqDLs+omvN7uzMpjHdblWVLvXa/lMex2KK8hBC
JJ1ucFGaqkOQSltmgu++BSAoQKNcCNZU3NvWlno4MXnqBDhRgLP9eHODPLH4BPxm
ZaAlRgReoc5Y7xsSkvh4go0UD8Kw3yKA3zDs5drMxWd0lf5oTKCTN+1keb6UDY9B
lyXUjoadYNQND1RdnHSm374TDeCMfU2cefmw7ukbeTlGL0JmoGsY/8JHXGkpT8zV
eqYTyjIzlwkRSNT2LBmZKeXRk88VQmsNhqhEn91jYoBbDaf4/twJ0KkIzpt7P2JV
XrNPw4cZPWNzicurSDtpYZZZhHRy+47zVrnWFjLQdXPomN7nR2RkRDkdDNdeEiWh
8WPTIT7A9wTpMaNfLz0MzxKuhaU5fISfUy2V6j9vuXwssdJ9ULKCXfkCQPDB5F5N
T52L4WYZ4E7SZQd3tKrqBYYNL+2YxrZh4Fx/WGlhfpUnaGIQyTY4FFglo2/ARwv9
eXbQasxZqUeRQl+ekR6ShONrvFOCcjt7+iRbxxQOSgDtlhY0oAHFk+fKqmfwig2v
lBtqCA/yYu0zlJv5kt4TulnNoKH+sMyYIYgEHhJscS8fQq2Me4t+3yR5+npOAdJg
Y3y//J+IuQTo25zzXG7Ffosdqow8H3g1U4GPS657vCeNjcIH268xmsJXKNGlmcQS
Zi8pBiDp75VDfT+cpCpssTiPGr2KBavnLYWUDBItwdeleS6iUNNId2ONIogcgJkV
ay6a+ET7SwMNiK1h8D7UY5jBrnpu7m+KpW9R01IOSBZaeYSAZuYRjXeyJEu6wGtr
u3KX7o07QMo0og9O/A68W/ubs5K08jxIPVKNcTYHrHP5+Hm6lg3lwmoXXn9Xij6/
NONe0nU1DInh27LQ+XoX4LxRf4cQcd9uWNbZpvvUFLBhCVASlXbOCZVLl5k5eW3v
LZSLx16NKTclWVylFDGiUIOJGY0VgfXlnVxEhOgHcuYpDo5oRUV2C2lbZpp58ZOI
+HKHnd3hqg0NK2aVVTIge35he5JNKBJuMNiZjqfDEh4vqc9nx1Sf9LfbAE54wO/z
jdzvNVxgMT0+q7fEjv9AlWl7O4R83f+1m4R5UJNwDy7kc/7ta3JDEeeNyFUZakNh
nDjj7hnYgDVvQbuuOUbU2PsefuAUOvEft9P/tLUAcmelHxVoDV1KEE9MRCAEScco
qtgwRVCq/b8aTHSj/ORd7o+FlefctzTkOtkRDRa/ZT5gII26ELeHdmSryKKjoIPt
L2MxG+eJEtTCsNOVurXMzAY7hHPOVIonmVTQ2r7JdKnImf9G7W7fdc0BE6/QsDT2
EpmgeJgOgyZwARfPv5g+N6Ni3CB5eNIcEzeNoSqjbebIZKcsdi0LwqNzw6y8+LzL
z40sGLdRHV4gukwTuPSca/gK8HaQNIwxSQhHvo++KwX/7NPUDFYSukaddfG4lPM7
mTl+odPNOVtYMOtwBvy0MB9Qp+3g/Bxce0rpYHdSKO06+cw/l9btfOiW5mTuOGB5
tOAyNtbuoqqKiOVbeikySwIMPSt7Qe8OglBO3cJNJUPbIBNKRTvtTXsCcKNFZA7S
VT16DB87JTaFKdEEZ/5qNWneXySfTh7tKl+ySbb+Mnmq+9k40bD+qeTNisnPYzGv
4MAHi3b/l6yyKU5IKGe7VxxWDQudHClLqwrTb9dvjkAGC2WHPC3Dla2J1OpsEpWg
b4r9tLw/MCr/H8EcFoShRKe9EV57a1KxmOt0XHEE6plDLobnTuVpByYTq0AAneYk
mefzEQ1jVjOCCbrWsd55LO1DVLONXlcxBiS6fazjjQPLFrTuBPzLBWZffTBrT4S5
9in749pW5AK3hwDqYydnKcHyQ3QFOVuUOaYrVIwcqrz68g27TRRQ8j58ZjDAizoT
qyvdZPoqCd5ikvGqKIkSOxwWPnf0JWwHWQ7dSJpC5IzLHzfx0bV6FwMGe/wHWBzs
JD9vaKi8GPLakDI0J5qmGcadkt2E10dB7HAVHq3Lf8os6xnlEySU551AOm1CnXbj
GuClgARq8ZKX1XZcXFRpJG1wGAzY1VHFbbFCVaOD7WTnmEeGUh1or43UmMLgc79z
aSy0j5fxYbAtMWaq/r7v4gRe7RCPkdFXEUMbn39Pq1ntJXMvDjXYRcQX3gZrB5Ys
Pa1MBETIiZ1Nl5K9BRIDWbGmOP3d4wPQ3kjDzhtdtSNjAHdPXGbXQuXPZH6d74h9
axVQAgzmXMKFqPZSKGvBMwuuUHk3mbjFlDQNjjv2lcX1kCIVRmBeWI4wzLwSVk9y
GUq/9MEeVT/pY5pCaHXPNuQSnaiUqZOPxhGGIlSIankEOnvb1Q+tINobcqZPLtfN
i9PJppwF87R6tO5j0VXdMf4zVUNSbI+hb+i/ex+Et/YYzoovmvv/I5vAlJPsIcLT
iYIxbzD5BjV2/v0EDz8UDlh/SRwm81Rh9mwLHCqhT2TXmMQJ5ciads6h/k3QnjmK
8OyeC934fG+fGsVOcL0G7LLbl0iM/wMxyNbqdFF0VMmnSrRXh9TUYSs5wvafxf5k
w+nArQoizl3swjQ3V7Z1E4uGsC7RckL8zCyow2xW2UBihMTQ2QH19j+bC4B0ib9S
c8ABCxNuUpyyhxxzO0N4Psq+6OCn6VgFCP7NJSDtBJxtIIe+gwLSxlodcxZCxxuG
1FKoaElSea/m0p5rGOJykUkWIEmVgN8MC2/PbBFFihCS575FH6NhBm6eN30rDJBS
Zv+G780IoqE+DkedUkBUs7Qx0A5llXZqECj33UZcB5i2bQ71I4jr1HfxnDVczoD5
vIChn5Ftnmput2iPxLG7tCNgp5ffPZXw5Pq6bySbiQeaa3MEOb6HBa3sOc91G1H0
AXj5MTpGsDE/MWrikkWbXV0dbjCvVn60DscnEv7+Hc7SAZ54R29Od4VImlbNooSi
33LHMmUBV/3JEjGr9w1HBVQAgIIzhlZbRZ4BrlqUua/gyOUPV6Xuu814hCjExXsn
4tttqrS8M6M4N3TPE8ck3jw2/BtBWQIE1wSNWgE59vx1yDnJdyff0SMfuHUIXjjx
XmsZjm2kkKjo18LHu+uQO/pCGWwt7KOoBVhFPItkJ6iQkEvIYVwJPev29KRIDMqV
TLC1XYiGwht2MRjJvu2yLCTrOafsLagfWps/+wYe+fPTWJcNubv+sxQuqAy9aqwf
nmROD6NSXKHYlE38dAcUy068MimwAK+THwmrVy3O8oWqs6lsoXQCVmjRBvqmXxgF
rel5wyVYzF8qJ8R29lQhyCCA64Lbnpf/5XThE4sQaIBVHQGF1Cv92InhJmJpy/JT
JOrdkAsdDLxmnfu5PKx149wDTGIT9zvh71TqH11ljyh1GDWS8j4SVGI/nqZotvPl
oh/6hWyjturyftVhxyGNgLtofN/IXMO355AAM33Ae6OJX8rvCIgZhS6r9m2QYd1F
GQZTPLiOlWq2610HBVMPZ6Zzdi2ho1sZrdwtq6CxhLgpgYyeCZCPN2ToH+uzKW5g
cc55V4yuMutpmYYvwosaE3fqvimgnc7V5zXmjEGzcMeWlVdQqybCsS388lZ5eoJ+
WoWJn0gjzZjQyOH11ydOHMaR5pKhH9jrxRAzsQQVqjH0FnMqGgRuIV7lQiuvdvVr
49trmkPT3tpRP+acvxHcXou2rwTxA6yXQN7PMiZhxmuvtUbg6NHvYeXPD+7jSR3P
ZQSmRWLtzKJkw4+CyEdlaZraSr7yRRliSVPNhcYiQ6HMALSH00ESjNcYu5Ygm8NQ
YuzbzCSnPiFNRquenkuLN2/Zo9Fy/cL9cPaLVk9RXKseL33K3lyxJqHpZwN+S/Wz
pQR0MqxAjM1DmllmZf62sU6nTwP4xZl2TX2aV/D9gAuYZvGJYo3+e8qD3NOdReb5
hRRPo9hs0mkKsaNStplT/VFaEj4jpQsh+FYunXcom/uYyDKS+Vuyyjsk3iFNypVr
iQaNV0LXawqtEUsIj5CnCitJp+aq3Yr3RN7m1c0Q0u5xSVrS2IPRVdyyiixKh/kU
1bg22fCx6u2HWyAse6noFCST01k360RcqaYMdKF2yEbCVJUfEbGNOSgxdxfriyaH
g11GEwLMpwW7RUoOvHUgleoqpNSFwQtQJ1laHzZXDucwTfARMS4LXry1npwAyJOs
Gs9TOykZN2xZxGceDMFgYMRXh7syk0EjR7U+8kZYqv86zj6GdrUVtSXerUJ2N/iW
IB4X08EMy7ss3DS4O3rMZYqog6msdL/7E5O7oPbgiSgRpEitudPJRNDhcK+ywGa9
EI4IHh+bKJ+a1bgLqh3bPd3MSHAh/slXx505oHQG7gZxP0zGSA42Eb/c7cRDdkQY
I3GWr+4Tg2os06Hg0M94NAKcP9wSwG+ZQfYsN06JaXNIWtDxNJPIRi8ZeeZbWo3l
LfV+hxJqs+2E7vo1IuHa+UJroNuqZyZMmtsgRV4juu/evu6DpGSd/sUvUi4laTbp
hVyAdno+M5MDsqh/gLb0aG+7v9iHMN3p1o1syhD3ZedmXn4Vej/PW+P63x7OClZO
mY5/OwVh4jikzoQwdSvnaUCPbN4CtP+C691sJUjumYgl4UwN0ZpNVtjLpqKq+tc8
LkBrschxouuSGsCXpSASPLPzstNLkjzEdZWUcyEwf3EGtLLdFC0168Y96ET9ij1Z
5ZYrJMv+XbvSnzje2qYcao3ncgPFneB+vz3td5PcMDPC+IJxG3frGCU27S5rEOX0
1x1jlncJ2EXVeGImaLZAAuAQnj4n2YzLwuV/qvxPjlMksIVUaOIDRTv+w4wmXqIc
yEWdgfZmXKoxARHlZvgaTQkrDNRiBgz2oZjaWOlmDkj8P7KcOg4sVoULCrXjZZ1x
EAOuYlEumt1mvC93SYXIZm4PA6uxLHHPHxHxVLXXe18vVpVWkZqwnQ7jniMNBWPm
WXNPGa1hrcUxsx8cuglhyeZNGMpJHKFFz5zI1u7z2EH+5lsopg6Yn/1GSskx17NS
9Glfe6GanGAWByd+GZTnhlsc/1jKpQTCEYsA6PmdN2jVm4d4EyvlCydEOfVOgarl
l19oShfRyQLj6rXDCMoflL9ho8d9ijT9K0Tq/uGKGdAfoErg71gX2roYO3UaHrHq
P8mMaiVWFIjWQwE2w2H4se8wnOgV9olc+EDzSvSye4JeYwEK4JNbWcLuEFCAHF7N
OPpVCJXvAHEynqlm4db0B1uFP6lMOwAJAEao6NprLpagzHZO3G54fIiUA8gqzh3L
nGd0OBdF1UY2j464nMchnvIkES6AjRmDK/CPOPuPx/keH9kWDCyQjBurdF11o13A
yPyQ43XFLB0Hei824yMg97EDxaOBpnFkGDZ8dJyYCok2UkzfJkQJyv8+UQhi2uWw
EbGCIutBFasuOrjeyhB80QGZxHNLOzISk+qbwfFzRaTtWk3TytNcvEmstYSHeJAc
/U6LAltrAvKdYWJgAy+nzb/h1VBJFtfDf9V+N1NG49zoj6ocemICrGvFuZpcKac9
ZbUsEVim/a96xE0mxbYh6EBimd+AmALTFqS2aTFz0WkztjIYJdEdHY78sgfJqYss
Z3AT1q7/SK9TZqlZKGPJrzAtB3Fo3/Zm4DdJ0o7Qb4cuGkuadCIq7nabfdImt3x7
SQrvVyUaZJz5ANMqhaYJulYqQEfyr7HHWOeTASDPlglCurnlFLbLSbxYGLfX0J6C
mOV3R0kddpWbtFlV6cecSuLmcXEKlXW2Mkc5ehA9ak2AvY+zaCJYKtlRtJhJe9dT
IzkET2TMp5fzedT5MjNzLmsuwUu5VZZxcCCXrzI0PPMxstuwgaB7EQDu/yToT0fm
1gjIcJz1BtdT7oJ/g2PbYrNKdzWkRfXbqr97WJ05Az/VtB5s/kPH+QBERwAEkQTS
APVyvcfbQbLbUC8yLdsTpj0Y7RW6tcjVxfySZZB690tbjLfJa7+rWIbnvZI9WKoN
7JwETfxc9+00RJzj1mYxjWzxKHt158QyE+J8Cjf9TxlkOVYXLYg6eAB+wU52CmCn
QLr31HykXH3Hrt4xEaLpYIJdkT3PP4bomRX0CZzD7Y6ESZG+3DlTLF2arQEFeGL5
NKmCzp/On2eLRGM61do3Am9yvzcuXtpGBGbIPu2me+hfYxm0nWu6eaYQzHhnHBAA
DkGLvv6CPCLokLj9dA0ibQPUk8159qKgZNXQzdw0xwtWVF3cljRcB6Kc00scql3P
bO3Ts9o41tjaCuc0YVb0GbWvSRciQwIuCYhSCiKX4QeeA7dCo3qN/crkJh3HWeDJ
gj7GT6u26h6smfEKIcSxrZLD3KucC5Ou/tuw46uQBg9Z2lrhyIQdZCt9BJ2ZVWRH
+EmqvH/OmqUCdgyKiAQolzPn/kX1zpH0CmH0WpZBOXJ4NE6f6kHjC6NppPLeiepH
GcApAnMZNftkrbCrAQvr9KXambC8aYZva7Hix765163gsDlycZG3x8Sgy8sb6kuR
iKSPKixA4V2F40axJwqpX/jgEWEBUI19tVqys9FSKcuc8/DHMallK1U3Bwp+duRg
zLzpZ1lN8o9d0e/hZf8bRP7Ae9xkqUPyfEHoRT6ZJA+c9+holGowkvSSLiMfxgsm
CJG6ZkhHdnjK83PyNpqj+3e6n9AKLRwSZ+mXnBz2ZzTxKiv9zXJbeADdXJmlt4EI
Du6WfWED/RFDjBBoXxeEgdXrgQQhISqhmrADN28NTTceH90rwgtEfvlj/BjMNbcX
MpXAgQ1PQaauA75QFMeHG1reV+aE1diLYEHqt/WB06X0dDeGbBB0SLryaz5A+DWh
AxoziUk9mXJHdlT2QjOIdJt+ViQamd9SWYt55KfhbnQXbZiuopSVOsULjLjYDah4
cHE/Z7Q1bIuUk7gQdUa+srEXlWW/YH2O59kqkeassPhTUkKJeUHhUjoV4XYDFSJE
A3fy6bDsRrah4Xw2Ex84FBhLMAED0awem8Vvd+uq7woK2DWSGfyxJ1UtrJPvvUh5
kcxGoRnuNuSobfzA8Wc6wdYDeChYdNDFeL4Ury4lvvVHlVtexpKyQ+rRT5M8mf7S
ZSe1Aqd1Ss29LfflLbu++a3NjS/w1R9WARYRrUeOMgG94BLSuU3EfWvBWRtmzeQY
R5MuNpPny0Q8E0RFHoRnC6Hd7LOd8PS1G/1MotvVoSDgO+MO2bwaJfjZENibiHdO
rQIJUitJSwxnMdy246zN5QtKWqa8tm+XWmaTtpzk4VrKLAxL9ouF5ZhMlv127+UB
8S4JzuUsf0k3ZOm0OgzVdCyCI50CMjoN4T0Du/jezjP4mZUDqubfTmGN8+LdkrRM
0OiOyzbk6vbeJEeyPpxshdeMbmt/AY/OWWtlO8BBtobO6wW6BVkWDzyJs+RE2YGv
48NMgtI+GSLfDeD9JBd0mVM+ty3CZcxHfSeQv403UWN/M667x1Th3Lkrol3MSHWW
8w+d1Qm5/BiMjstNSzB04cR5T9hACsMaYChwRpFA/OxEn5yOApnze6V15IEJ7E2P
ao86rKj5Abj/YSkrhtqid/Y88Gv7RiE10m8t5D0a5Ju3CGpoTzP9KTPKWcI4bkNL
HDxYSrXoIVMG8XEJ6uklcxYxX/HLeWnwef0o756L6y3/Ob4R1gMSYueRVcWLvT9e
Hen2YAT8e7wQBJ2HplXGMxPQBHAMXHCXcDQQEko9pkbe3aNAAhIbry37Sk7XByRG
TnZgJNAQq2VLNCaeVAkMrV0VHoC0K5pQZswYhkW/7Bpd2lDi56MgFz2WPX7EiS55
QcQo04arKReN/rU+/IJ1teCp4vgQAHUgqw60jisr67cWG/jYFcpaxaX8/pqGuFNc
1PucbOjk+liL7qqRLFpNlHJK0sWn0EBhMJZKr7kgWU5kanH/pKX1wlfTHsO+2GhZ
rVjOiYifV6nydAYl20x0jMYNMe1dgqTdLiFnokgXP71QtqUALkudPswximUhQEwS
+wRbIQnoCy/F0tgxUDS3wyxrp3L5HBtJmGJLikBip5ZNxdxJJId2nCKzQqKR2LG0
Gsa98sNS+2s66VLVrAznirCo0CyooXfRzIwi5EbGXQn8tAJ+AHSwEwvgIP+HZRC0
iBuuEIkCJV7o4JfknaYaMtr4HuXnK01f6Owl4SQuHcMuiC5i5/xPPPyjUSW7cx/J
QxvQAVtp6MJINwzx00YzqsRKn/dkpc4Nu3T3mdIaNiH3K+n0wrKZYdMFx9wer4tl
LRKAYPwMHANjYj2zGuVOX9m5bi3IfJgxDyrC4HgLmLgqYTxJ6zgJvB5klTJDtCe2
faGAOlE6nITPJnK/Lo4EcRxcZmro64juIZZMbH3xoxW2SD2tiUpAL924o/gnzbm7
6xVjlr5GnkhVFtqu18kdkZP5wOKh/EfE0DilevUHWwx+EOEQ0EelXDfvj1P0ee+h
xABmf5SFlDSobidEWtEdQReH+r573ou2644VkMezNW4NeEosIMaRJOkhMC5vPfx1
vQK5EPZiOlBEhmjwuy/I3MaN+dCDLQiuSJ9TO6RCMVy/fTKD4Yae/gSE2W0oYByv
BSvZWKLsXJKfD6GflBn4s6L9qztHDYbNjaWv0LHmZEfEkiY0MGq8+V1jZHNhx9st
oVMUg2stg1jTFP6nnI6JqLxhZXBp0xd/u0xciOC+GYv7MmPVNmajjP4iMLBVhx1f
5MRqhfvj8l6KKHIYXXbXEjij/HBPD27aR4IsTS5ECjoXTjUcLf8NM+YKQnWZTmPX
1WPxjyZu1YwKR20SurkS1i6dw13pq85QSU2FPho1p4KywUooXWO0V72vvCv0sr3Z
yoxfg6kf28Y9McvjDEZZmBmj4e7s1C78+1lO2ujfQuu/29ychP4vfxtTvbdOn8JV
2Hr2HD4oeeIz2Q6zvPg4FLSQXLs8IL4mm91jfR63XsgC6+LH8FJy7nKzcvHqvIic
phZh3BhZVCQQVBplSzruoSW/T+WrGoDJQ6Ci5rUEqCZFUhC53Qn9Sjbd2rJfiYsM
XPu2t1ej4k9ejVj2+8vLcxpQvjeW85+0EZehU9J6ITVnKrzbxsWhZIBHIAeQLp+4
mc/18j6Yq6MBnTTg+8hA6YEqLNehIibGkY7SEC6FNoozNnd7L4bNOaqLau97yV01
1tRAjBZjd+/FBaa9KMvLdG2NyYwxjFukXzyK9tYWSLAzNYmTvRpF1lq5lZki9yjN
vUes1MliZw6UYZLv8Qm6RpLw62NO2JSY5KBC4Oq6kvsqm3AVxFJO1YbXWzsAzB6X
YVHuRts2/C6u+iindBv4/Rrfo21k+VuLf2nIBoZsT78rjOB/1j+aprOrf/RmCfcY
gu454/ShAxLdtEEulldUpbxf865joogbcH6CrJt+pzyvdvzygNJld03xHLdwaKcS
HAxBwWX6pg41pEr9qf69A1CJ2bozmFF0b0KiwmNL073YEN6o5JFg43nYYQZEsggV
7xQbS6AwmJqX52lB7gCgBPmzhF0Kc0tssliDPPgUDbLr4TQmIGX6VNt/0cPv8Ikx
O5sb0YcLCF/PYQ5CPqhHVxHSLlmftY8uVq+p5FjAO879C5TLibra6ltf0nSpOiNJ
sK9HSUM90kJbgOoiiNy1Y1ebnQGhiqH6/6Y/KVYnIYEmIaxWFklhLYsMBagxVNRN
7SGC8CMPyXKLLfbybAqXz0SUvn7zt4+0U/VPfpI2B45FBS9St/RramxOep1VJKOh
tmdU9Yl7P6Jm8BhssXgYY7w5vIv8i5g5MM+wkzuyZrz7562i/nRVJUFLUnBhkBk+
/ALJa3kgJeSaF4FZeJqcCdbr8UI1UGssaJg5ZP2v5cGnEewl494/XFUMnQ0nG4fl
ihi1GpzZzVwksAU1U0XvNjQCVoWrnWoZBgbpGXQqfQro0SR+/bSdevkRNxWPzztY
+DOeanMtNaJbUafJowp3wKWVoGeBHsRKWPcPFknO0bp+82EnKdI4LYuYoUfLIY6N
tNKDZyMjb1GKYq0VHT9r/dHiGmZx2kxZCm7RYW/WwPk86vErVeEZzkyY2gdBF7Ql
YNx0ZArgfr8XDiq6SfP2SPTla4c2nJ2fRv5hrV2CLjNqzJXS+GTlaJjBKzQdeBnz
LWhZbCEuHizDWBLce0BFIAUPPQvxuML3GPnhlYAr/5C9zNOSx+wdD69MyfwZBDOX
PY19NYhBkD1bl9MNHyJ6B7zGPITJAfdcQxOpvJ1uz42XQm2eNzA6u9rQ5xGX0ZFJ
QbP8gB84eNzOLgPKvBVkeZA58dtM26Z32g5zBGzHRq8vBonFtRnrCHTMwgDKYGnC
PeVhW6R8GqaDgvyeVU4Xpq8Lxd9ibgkfmG0RMbSvJHnE4Vo0g+pHww4Gnd10h+EZ
0/HbiWUCi3vjslITfzWMrgtxA4p6gEqJ8s8H7CCsypIVpuhua6HoODR8H+9/1NMN
qmMnGbwQTx/DNP23CFDqBMmqfX8cCXUJlRRjOsoyuHzOgydmg/vRN7y71X6jZjOo
5Qywk9vsquiGrapzsjUrRmTZRWS++uB3YK+AvBCnVP68xwHvHlz7XVTEN9CB6iqd
m0GTea13Qw4YjYCpEiJqUvwsLW2J8ynVH+4rPCzynJgf6wA9agvJTegE9YIVlWq/
clcmwdGY1ay2DK8bduJG3d4lRfkGP7BrgWvL7+X2Mgae3sJrydjJ0QPzBiK71oP7
YYibI5vop/5wVjO/j+f2fmBeCS1bWJJFEghs2uR5ffoRP3UNnuQv87CsnC7RXpOD
yEMSwwk5QdrvaphFP0ukJJnSI1XJN6wl4MCdyUrmcYS54jdqxTSS/JpKKGi/HbH5
CxehnJdIyN+Ci39t6dOcgqiaK9NTyfdoZxIZVmU0naXzGfwx+SKV/2DsFY3QSUpj
c2OzkBbCVGdDbz40+meoKUf+UlyI3eR5bgUDTnYhCUF0o1NV3b0pudMEE41AbMF0
DVXzOSqmbZWPgQoxEMROLw2CAvZ2h+xV9FJexlrEW9qVrsdU4UUWuzps9PNvDT8i
IYeD8WYrNomCNIDA2m1OW+nZM1D8sR4hTDMxenFNhV3K7NHIaHCgxdWz5p7C6aJm
EjcZ4sUeR8JvkrMX7Tq1OxDr4OR27SMg6FHAe+np0M44lIMuAD4dDMUTWePpqEwf
YOSLmkcG8Af+WwIWJyWwT2IRmfu6wu6Yt9eXzIswOW9SA4wOOh6quuE5izZWkIfD
Ksc7TdDbgRANYmLt91jCPCCT6lL+sqXWuxS1A6aAAUaG7ErQuXYMT+1qs55qq7J3
axAVaCH87kSDlPXzz4qWPYNjvoyYq8QYfJsxGfVvZxGEmfB0mV4ZukGsUs8iDxA5
t4TQs7DcwSsPTI/mPftz7aPHyF5A74rcrxDKKrbvoLUzBXPCscAm6xosDdvu2isF
U1hJnfrk3QH9qhO3JgPHdwcJo7tSQQL2qrhe/vDv0LnSDMBjzVoBmoJ63+g6K6nq
Pm+L3sFJGmrrR1mEKjr11z+jGcxeZ/XJcs6QifKCmXoZhata1rpFgAsU+pMeG5OW
lVc0EFAqqWUosjggPufD1ALx6NXRaPMyLhlcw5tT/ujwECtQq+Tp2Fe+l7e6sFCo
INM5YoUvjbTmTs6yZics2YDFoaRWMoesRLu4jCgM2D8MRFRy5GIZMcMsp1pBuWEO
vyC1JTDkG1LNLce6Vw2d+v5NhkIvS4Tz7FcTAQ0dz3MLjVH0c9f7nXTjcwiqP8Fn
+inylCfh9RjoriKxTBQFhRnwYQBgVLC3ZNlM/RtT/2x5yof/7UzkFMYXjJhxvvkE
FfPvx/uoDtGnGANer7oPHANalyISiC/69KeejuyQg2XSmlqqfajg4csZEd/smXoO
ZVTS7ep19Ax/qt0lisnfEeYAWwCa4G0jcD9NSMetT6ZqEOmRZCTxkia5bnOECYEb
VxNowmqZJA7DeJ50UuB8pDOsPjzOfhUKtViLGJQJ1Ii4yNXeJNpp66ISd/+csBn+
Wjh/hiUgm8TpfDCkz44yMHAFlHQoYjkqwpNlcTTJ/RcdCoARLOhpvqUlEllpAHQ9
0indpGYzJhFhz99dSJ0T8Ql67PocqSMd7ZDhJ4syBj2IP4DxqjByHg6Tho55YCQj
uhXtIonWCS3k3to6NP28ZEWHMaoQtA0MG8iOaIjNwcjFnAk9ur7vOUNqdEliBwOX
s51tKp7CraTBLK3a9mOqRZdq75jAOsDDA7FY9vGmtZTZ2QOpASeDsFI6ivzB2+xm
Mes+DXe39lqjr7UBOFejsY5H4dIr7fSImF+UUye2ki+DR7nFdRFM3jTpQ9oZEgNs
NOEwF62TP2xnRio/dMbP/1qF0i6jZN3FMbvFz5T1aYz0n/JP+SVW2NEFffM7QPYZ
m3uZZdn7zo/5hau8yD36bVdi04u63MDzuwTziFc4uefoc3qE7tAow4Oz0ki1/OW9
CGH2hGMWupyo1lgILLDXLYbI02LIBtLo1nXHkakUQt33P7k5uuieDQuZdZmePGjf
hC5kgJILxA+KhLAg3tNqUlF2yZKVc+/JulWiHmSsuIoDAVSRxV6rZBKgnGKF7tpg
cAATDlacLTS/cAOBvUc1acUhVWCFUrhQHAiBXibVn8tocJeq+uJ79Okq3z51X12x
mUr4Az2tX49w+72nRQXumomy7ioq56ya9qBcv95+6uf1YAjDM+x4rwYgq82zcf2h
E6/12l0QutB7b7uwexEJc+x651ewi3/ElpeA+hRDwTXZp28EplN4tvXwbKScD+30
/7cX0Ll1skj8V+cYGwCMhXtsLj1QVig+yUJY98hbzxzFHjlS7hcLudvHVJfQ+AO6
1EWEbtNLX/ivofYCK2PyS+4xOsa49xjD4RqDwD+Om57jQJkNZJ43cdqpJEN0LdkK
Uto7b8LGKksc0WJT0sKHVGzMybM4b6MGaaJ1p55A4QFC7jd+8pkp1KTp5s2io1T+
JBc38EFhhZzuZgGwJxeXXIXptmEkDnx0Ik1VbJbjT5RzvZ8rX/ENvnC/GugokfoO
9xfuwRF5YqK63oeFm5vrV3Iu1dERzXTC4pYsF0qPTW3G+lzdUi1VTZIGiZTX+wR0
KxSPvsDpuyOoV2GghIGPRnJpIAX4+u9PwpnunodRRM4+Y+c5XilWjOwyA0hDxb4R
LOqwXsDdl6vgibWEX/oKiOI218POddgq1pceSDusahJT5I0f5P/8YryhYpDvClV3
qIccnLC0Pkixm1+Ydfit1qj+kQ+mJmNLolAIrXIbAboY38TS0rHRIrWTqwGWdde0
vjfULFCtk0/NAXw4aTps+RUK0HXbE5T7/TIGCNDMWoCrKA6znlK2fcDhJir3W9Gh
xRJMc8cjXeNbvYCnuPfWKMuvHqimT10v8QdAEdhcb07nUx2RNCm9C0kzRAJIzqk7
TKzCinocj62e//2CXQtUad7Azpk0XJIDglyvXZgZ/NQvtfIZkwKwf9za1DIbpIL/
iiMkc+hnjak4ZEnIFIUbVp7ksrdpRULcFaXux7AhrhSuqQzwbSnWlX6qW7pkG7s8
zJ+NhlrXWoapLJ46PlSSdi1N/dEjJAtne0KSagU5E9hBXdJ3bl/plbVgUO+XUskP
8+h56bjdueaHnaC5dYaF0GhzzKuFN6yBBeyDh/gF+b/p1Nf1EJBt2GQPivsFYkiM
VxLYpAUM6j+y4h81Zv3pDlt3GPfHmBek9UCyV5SIguGMdCgm9XfqENsk8RhnwDQ1
80XRrteIYx4kT6bzHO9Xv3sxImxmkuPRiSRnJvf9bAnPp3qdwZF1ianzCFP2Mh/n
oYHVXNBexjw0SbpW0+S8AX2NGoqcwP46PBnKEipvyDLXLQrGUHrG+RMFm6FGbR+J
EOY8091+4Mb+nj0tt/A4w1pdRyg6QzSJQk4TP6UolnGGoY7gvUou1+ugiyxuiAzv
CbbXMnz94qicAX11+nX5AdyHb444CziyFfhqvyJLFN0nnJmjJ17ZiU4I5bLEVSjR
ZV397mE90sZolC9txPTwAFnJ2n65znlpOvcaWgraONj5/33WO7iSvVjUgAdfvNSe
HOdEmx6E5hXXvUXuE+ib+jej5u42/ml53qji3G9YC+25f84/tYXScEsJCbY//Uev
klMkOe58sXP6MjFt04SxsOji6K0sPOvMEb4k1u7fZqZkM3pNaiKNIG9EeftH1A/8
i3phAgp92QbHi9Eya8AWW4vL8sR75s3Mq/PGtLRYpaiIAeZ8LkmmGWcQRFbBB0ZG
Gzo2kC3VvT8R5EG3YVlT6V8cHXw8Te5Fj8093Cv+OPYkW6j+wq/2UlzNKpIX95PV
LsQ8dVaJwDuioIyqQE5GxvyMhk2A4rss/39Xug+MWL7ZmxxCbSvEIpMQUbEYbTvN
tPR6ptx0cpnGgzMKDc2lTMep78MEIbtdOOopxYxj6LTzw6JQxDhlpW2dz+VnwlOv
/ARasurA/6p7DHRY4uGZfcrpeeuZ1dDE0nsMnUrSn65tevhn+uYio4NmihHnw7ts
Lk/AriLaot0UR2yJ0M4qz7TdLBLsKgJbDFatWoD40v1fMM8zuiZRlfTEOgZEDW8j
WOn5AFyDzsv2M+iy8XP0Qk1V/WEfUbfbEhzj98V9o8fpJshF3UEpJ7E0nHwZq5j9
TFyMNH2SKRVpcR18GnT/fgpSuU/vxdDveiAKjKQ5ecd7djqzq6Aui88GBTVvLvPe
mcUp+iMcchJR51Eq+IW5KZkamkJ/ScsCdd6UsAE5VE820WNbGbTh4tW22Pgr2kfF
tos9KNNU3WfOl06MtC13/YbMprmGaDtdHYOLHvIi/zYew4zGEiW2SpmGIUqMODj5
BiOq3aB1zMEOBIU0eSlXPkSDlIjpsQD1MD3E3geJHvkeugnf3kxT/klr2YgiQRAJ
YiZG6nrcx8DksOMrlgfJRoXoaLLYonaAuQ4iX0xONIXLBqeG5SCV+APgBw2krdWE
YwFo9pZC5tqUnhPXD51C8Q1sGzLlhvMIT3lUPhNmKi0Jn8JOELCRb9Zk/R3Vm1To
LIbqUNTqS9fgF1boIhTSpVKrRyhj+p59jI7s6PO/GUzUeWnP2G198e9AZEXAHN19
U0mkyKcnUWn3aEdbs8mWIbPV8JrEPNE3RwHtMpQMGxUesu/I7oUebZ9+J3i6x8j+
rI9pZwQlV/5aClWVF/p1taLFqrap90hwyNYaF4udnojv0cWTbI/0TIrgz0ftWC1J
7Cuv2AjxhqsdOviISSDaednzgn2BvA4oEnCCEPyacUaNORNAma5MJQShFeUEBCBS
jPpmfSojwBIUEZr0forsQ3TtYG7AxV4dNQBiilinyt5hL9pQNf5AswZcw/7353f7
N3m7QO9Z9adZN2PSeucqXcVodW14DkfGt1dB3pCUsN2SjHeGh+4KIWP49E2Tn88x
QUyU04o0QM49l59/9xl1NlfrDvXdet81MpR/86plhDq4yH2PBowetOk75+Cw61YT
yxSC8C6Iy2OKe0Ysq6yXS06033zBxnjtcB5trT5qzFcy0nBdT6i0/lPiD+dmkckg
P95Brf64Lnd9k7dZz53WaB1K6POhJpTTrpYvagna/dWkwULz0k5O4prUOm9pIq6A
hyqOAwuXtLu2SndX2p9RbpHOZZnw7pAco/HxwkCV5YqJx/v4DQkyeqIY9QcIHZV9
xs6J124BVGbOsFoGitAoEi2+PH7xgdUuUys+yMspUqzz2r26yvynDILT0xWHDz+m
S/hZG422H1Q3550wMnK69Od/3AFRcZVCGnrfaFDrfI27OIh/B9DII7sSiZ0s5DkC
YnomYid/Z3li5GEX9xew6LopifCfDAjHVkuSBM+fd8Az7cMtVWZT3etNafG8GBfX
LM+2pwnNRz+/dIjTTWP9qteGylu6azQCQazYyQvXPrrdOtD2lMutW/hdb9Lxfz8/
6NqiVFEVhKWxcHM38NLYULxt+AjLJioxH1UvUCJCRPHZ4/W3WNzSw2Jddk8D99Es
KQkHag3MMgbreBGzVLJ8hCHlV9wzrDRXTSp9OmaxPeS8EHA7pF78q1gPRFiwuIxy
l3c4yswHa8HZbHeuGdMbKBdvxklBt+7kK3De9nrI1b+y0uFj7vA1H9lpkDZF/dNR
dlXIEG8yqdRGZVzZqFY0DEdPQ/EHOcEbx0WRvKNW+ldbwpxjlnlENQ8yc5YLfsxy
7M5R/PpgBGL7gS5YcjTyjDwojiukmEtOT16r1emSs8aEp9jPihrMUF2Ev61F8cfM
CgxASsFr5I6VFpQz1D+m2VSoaMkww+iAD5ftDZQWUAdlMRF6qACiBbtP5umqP5wF
LpXwqCw3Ugy9ROgQEkTTGCyUnX3+T39aN+q/sgq44CM1NgO8GnyH7ns/ZaXvVyYH
WUaEd7vHaX/AXk/YNCH6hFDjwRLPxqr+X9IJe8w91C4tEJayUF1G6Mo2Wc8oQgVJ
OZAFvXnNdTofRf6CKOcV2e95dQkueYJzTPRRXAHwvwfavu6pubWDvkDMY9eknxdd
qy3qHgqZzJ+2TLE/zMTJMXlz7i5H+cVutyn0nazd1dqwMs/D44FWFz76O6dmiuY4
tidmXV+FTsKkEvjvHWhp7tEgc4brHFO9Pz+xQFDMw+zJYCNc+RlNRxQ5SPfICT64
eARbpl188FBmuDKfCv+D3JHP1lijr3wQGr3eLcNwLMQBp5p7tkCj3C5HOzde0MSy
vWW4wbc0S7ALc/9+IknPJRCSqptQx96m/Jpr09yierR2R3Nlvf1r6OqaAnTIk+wV
BRBCfsQqZFDml+sBr2HEBqwNFIA1XA32Z0yBfsv96jEtvlrEt6O/qfpxHdgtgB9U
UjsWapjZoQJEkWaPe/i0obi5CkNs2JmBSdOH7IEUl04Cz3/9xPIq7yCR1sSEae7U
/hPhXH3t71DEmMagiHR30s7RbqNyr6x4N1zEnsDyZ6cbBE3dPB5qyzDL3YJP2k20
mIaGq3iiKOMwuRjehU1F0lsHfxQVjNKNqebuFV6rpS/z537CKMk4z/ifY9ocaVU1
t8mP0Qblug04wS1leJOEiUBo4b504hn6XH66apBOK1/jjXmHNq7wkAd9pSHTxs67
b7eCHZmzA5FzoRlbwfW9IV4HEO9vpxo31MIh2jr7SIo+eVOIbD74+bHfHxoDluV4
7ww/vsagy2sAlYPbOt/FWNoduyi4/EcoSfnbwGLgUANKGUSZNGQYbM2zA0sWITPJ
b6PgQgbVe9I2/TKMCscqefn4tqYsJZq3W2vuFc5olC1QbyaSAjYyz4LwsYBplOlX
DUjpxhSwQgmit6dMChpc1dWZVjtPXbgSrhj3oUs4FO8UOI27vwntfYh+wlaUrJZW
yePc+71ixV8XhGCYzJtT6Xc5ehrTkmMRfAMKIY0Gd/P2nlHV5WzFDwGtu9aK93BB
LF1aubYE+xcKkV5KKiN2yoOIGK6t8tmo1RrK5e228ByB7nIBEBZwm26HzAwgVGXO
hyk1nJItKLwh13KIomJaJdnUUtRLynDjzLEjJI3dKRc5npdPoI1c6N5PbAjBNl5n
AUn5XdWwRgAonn3/I+oFPhkPios97RobC8Q5Dp9ioO4f8e/ZaYZuN3qFk/y0wpM1
xLzw/xnhSL7wB8X3wMTJYjGswLv6FbEXL2afPZEIJlL3+zuYIYj+gu+d1B/a7biQ
dmFgWC4u1ADJXMWtz+1BOU3PrlxRZDNW3wlxT9/CF/bmCYp+QJEYBPC3VdsiCwV3
3vDs8R6axdOaLXQZiPrT6raXyrvaUiqZNXP9QtOHQKkOntfVb2vESrALlao+CqPo
rlbYnDEacjEsQyUUuQd9lSx+0oAEuMRMauql9qqLuDVohWD528u1Vgh1dnSbdP3a
wXO/gZR74hvFJKe0b/At7eMnwg6rETNUW541ptoTDH/YUUN9yLckcG5OUfQVtvWl
HpcYe0QeSAVDgw0Ydm9ueS35j0eYkutxutQG4ZZyEZMmOkK1Av1tWuCUOIUTWt+A
XWuBtriGl5GqVFkVgihWVEJjDzxbSmDssn0ul02gSp28ocz3IA9DZJLmwRgyXIQk
O95KckjZ8fHm1bfFB1GLcfhoHvgWqm/U8q9bxPkJblUZmtsoZX/xfa9G6AJHO5jh
MSB2/Y6ECBfVYDyt0pDMuaN+X9yy7cnTQLO7MI2BjQhw41wgvvzAUIZRJrr/6sU2
6x6WvjMt5K7QKXmfUmWmCB6IBbuaknAF8ThqK6SJrGstAs4bCm4PgjqWvHcXSAL9
n+PwIV1zIkfXw0oRO46xx8SQUQvu1t4vV2sdLsMvivdba0ksdO7pneXlDYX1viS6
XHdKVWEOIT31leI1g14IV+tG+bl7pBXIWBGqpMyZWew1qRTj54p8tarIQ+duoaq7
TKhUSZoYZKMd0d/PnsDiFtl4vjYW9hvLtJsSCPtx/fjriC3fWNkFFc3Z0d468cv9
y08bQYoRLkS/RRJnzkiLdAboW+wA3vI4X3M0xbFmTJOr4LEAdkY9dK/Wa2NBlkUU
Z5Sc7asPCUmkZPCn+5I5jsrs0HMWGWOjzDU4jVJP1kc2RRexSvt9bhUhGfoOX3Rx
QhuhwLN33EqmjWOD0dizoufsQZF3IjfPMBiXB8AiZtitHA5FoKrNmEdb6kDuimTy
Ku7Y7gtezhwfbZAQzh1BgrUnu5SZMUF1tq7438+MJM3aWcYFjUJp3IbFg+65d4EZ
bk3TU0DEzvcTOkxRN1Z4iWfJOwC3d4piXJ3/g/EQOELyD4b2hMUF/bnwT007Ut4y
OhCqsjJ+4Edq51p1ZUdXIWtz4zhqUbKt9ig2tucg1oSI+lTtwDu6dwVdZIjcexZ+
PtkVlC0oqYoeBwxwPl94ZIzypcM1E+XqxNiVgGkr8TFg9cJyFh8gR0FnpW+i4vi3
TaVhANPwgo7TYsz5vsjxCDEzVhrNW2q+rFz8rJ14Yj4THgTrskMxxgXLCqwbzUuu
QKFtC+sjMOkk9SMDpG/s0Z+xHznHcbQh9Zoiy9mAEQy2lPECupbu2tKJfgpIdkpF
3HdXB81OfyThPd4qeElDXbEU92gJefcTTxgnYHf/kWzTgmLHbJJYiWvfjy/Qqugo
VcUpXtTbviTJQ2gWt6dHUzPy226ILeuGj10VlP64UKRDVbg4uma7gA1NyouJZI12
52RO73FFSkv6BUKRmoRd4/C7Nhc4Bjvh3HzJbpDf3msQc7x7nqGFv7xNic1x4Tne
APhaVSWKU83FS8HlGJbFN1Ic7q5c1yf7qlT64R/S1nloDixp1K3rBYYcfPwLvzLo
jeoxwP9NxNELqwJ5YCGUB2R+hptVW9yWI5QVqXN6UiAixRf7/C33xSIvsU987E2A
F5Iu7QF2qYcSqKTlQQI0ucUyAkuhZl0d18zVfAqZ5bdfMlJlkY6uhA7RkWNdvjzz
z9GShDUhv3klOL0WTUtj1S/xL3cPeLLZMJQwsq7QZQE3yPqp/Z7ZthA8CAashjpD
x51bUKZLNFeS7SRuKGo1VTZxSiTMyT4dVy6TuG1XGwuyOMO6g1LYMWzpjQVlBMOL
p7DKG2385NAnwQVpNO7eCq34WqzjTlJdweChJpWqILHG6EsAw7ykh5GfWiZtoVsR
3tGarfMBx7qPKszLiaQ6aA+XPXookc1hLtLrf8mnMKXV6/bO4qvuE5hriThMEu4i
SYWCH5v320X3P2fi1x9eT1UAFTmlvpBqGcgpErNMJhIuOvFLOSnVc5+dlxtATdB7
4j5IW8ujTcuf7GH4IHhWkGSDYrNG2svUcK+9jEjbvBkDFkgfVPXvoAbQtGxstdLw
Bw+KPugFIEb9eYWPXm/CvsSsMQJJ2Tqx8nFP7g6/hUkAOR7mJN26mNMo1d5njULV
shsSe+ZGUV4ddmRC+8squiHJPyjcuBxNsB0yf6631B5aN4lxLBaAOqPxN/ljTdfA
1JxdD83Rx7ABWgCbuiQLMHeCWtP4Ee0XBgotY85PKekjDO8Dyh84JTcyclAVK2Py
SxbfPgcqzpoXP/nXONhcubxF/zWCw3rKwr1eNz7TZU5QnrWIL3dS/y19TGKgy9Bj
DjJi53V7x555BwJnK23OaBDlEkzE6y7LxxQpp8fWn9G+zGFKhc6Snsh6CGmuy/Mq
L+5EgVt8Z9wCvD3afXU7AOgSUFhYOl1/x/al9+DUHTLAC1i1mS1iPD9fsP+y9lSO
6tiI3b8l++ZxFuc+q5A6j0CC3Sr3KyE64s+N+fGxDICASpeodcYUNUUeY06CwELG
9IHZ6vBNL6s3SClmVrhAo8/DSY99rDpilZxuYNg/RHDbNGixSVfTw2NGDptpvxTt
6RLkNNh6KaWDlwra1/aibZNGs136kn8xOFG+Z/Q24QeCa4M8GGE8jWR3AAD7EUtO
An14XxdDdgqyY3YAC64DlLx+zFVs9h1ewb2XXIstc6G+Ap0ueB5Z3vJt47W4bRpt
/976zTahxQXOcZCxivX5YcJCKlmB4BuAKLxAZCsgSexkqHlEAd35qcUXZ8vm/4Im
yIO9bEX9PVU4w5e99yartqRiwwLwudGNYJrm+GV/4yXRGsW5nxAwVe2hK24atJVl
sCIH4C7wnGq6oEqtwXZvs0/wQI5uNJqb41uZCvVnfH5ANt+q3rZWGRLV71HW7PLB
JY/sqkb27RarbJz7IP3tUZFS756Bzqje9JmCy2XGmXVGOidS/hjqnZEs9GNl1xlM
O53tMtxvwaabvyuY3me4bsH6G6PEJnqBM/uW1KIa3YfP8aPu/CWu9PZAiZIXb5X1
l6bUmDS7+4C7oULuNaxcMZzHvNzxULYB1kQkAJuYH45YziKqlJctLx25c2/2ZiIG
S0Iksw6x5+6e8vN7dlk945Eqdt6GOeyqcpoIR/NNEf+IMh5LRy7HuC/xBz+VOdj8
g7iblZlJQTLDUejTJGVdOfyveogurfppv9FjDfliDSCwth/dLSdjD4IlmFRccj4+
4Eb+X3FUJjwZVFUxek9ow3jvev1u3Kx27cy4k7XoNikEhalGayhjwLN8U6NpTsRG
f9Ckhg7kSUp3S0B9Q3KxZoQLZTe8oeseJeBpDLyUQ0x6pGhGWzwYRAWrs/eF0jic
TdWdFs6fhxV08/KIXshJPnITHlRTbnkETty276BA2NAa10dAuy712nc0yoS83XTr
I1XjCPP/y5BtWf6len0r2nYFkLoCSfjMLvIUP5OsmXFxN/TE6vCATg6n89YhK/3T
RF3q/KT3x1ETesxy45vb7aK770jeWXdfQ+p5BQEH4QyzTasavkC7PB7CLBdgCLaE
yQyJQUkgwaAqV6uh89+4MR6djaYIFEswFu/Ud6gzb8gx3uE7jxRn23TKh2Q/QxGr
R7MFMWCWzE/AfwoYcM+zuZsXoXfyYR8xWUWUyCqhDKEh/snOo1wm6K9FEJ869xVz
GDyPcd2z1mdWHguFzq+lqJt1Hmosb9WVgirZmVdc/rtybYSbGa4g5TMZZgzY4UBe
mftTpMEuYDZEENI/5aG/hoCtdL9enQpaYgKwg5p08ZMUVypbpltJospAfUXgLtlu
CJog33ci0WiEKf4JypHIkBYWe7woL8RpoN1SLiO9vWavXvVo504cqLh1TgpIZ2XD
OByJgDzlXzRYD5oBNOxu0uQQ6r9qi/pO9XMkJZ358FChIateiLD8ZmhZ6vYSVXy2
lkc6uotnfAUYm6kFyx5ckj9t85tKFGfPJ1bop/KXkUyDg8/0Ityob66RB0zkOBfn
XcfgNFqHRZWSjHiDtOFKa+INCDolhMu199ZPiBlx607k0G/vcHrLScalPzIHxIjI
fXOolW+HQvhQQIOxM4EJExIoCyDK1Lpk8ne3y4XL2doff3lWfTTd4qpBDCcU3EWe
0tEn567hySyn1VKxuGkC2IKiwjsSUHCF+TeA3lRRKedizv6mPCv681mYJAUb7KDC
u6VO6hDUWuDdCiqdHkBSTH9hQqHnZmKBqu6QAUc1/wY4CpYpQ+qkxVkiLF3iQz1h
Pd+7orVzRUbrn9JrBuUsYxWXBEgr8TTquWRUSaGQ4J6WzBfXPYZ8oC0jIpU/oKzM
vUfSJh9kOnCGWAN1PuM9NR4myZlChdwot/44IkYB5IIm3d1pBosdKbqY8HS+FKzM
g440HX0KRuESDgtGDpcbbxZt6W/M0qkrShioY1dh7V54VcD9zgLJqHyqUsQeQPNL
RKU+BiECfGn6yuNgeyX0ZTEJMvnDjEOam0lwEasHqlYsL3JUR1n9jtTc0Blak9yC
qfrC/OMkP+wbowZOu5da6/GKcip3ZYYwjqKAiQME/7CiUSUF6scbJOmraGWVJKtO
dpEUIFTFD3X2z4M4PNIGU1bR9p4L97F6fm707CF1CXo2h3bMgro0VWkqMbHkz3rT
KBnnEjPnH+0hD+FNarXLwyY0t61AmuVHJtQGW1mpx2QRBuBdcsHedCT/vhcO7Hn6
+5bPzOzRPJSNhDhntDai0r8eX22rabnraf+9+1ufHn13Vp3fWHMlzSgqp099B45s
lXV9pe2SxSzg9+9DwoKtpQLFzkFtiHQgCqueG7WM5ZwngEyRcfq+64zQw+aUZYlF
H0voshXnk6bQZvuWNFYLSa4mrMEsRZ8BBPtIXG9kpb/mNo4GgeG7v0H6vywcZb+m
AWIU7TZJ+IgCvJsrMUMjRJ3SI7oi62S+8ubRHgBLefePSV8+HoZqRTnr5M65N7XO
ep1KV1zEXCCi5xXCry36ZclurjQNtX9Lqz8BPWMUjwlxqmNN/8ppYhqk31YpP8HQ
hyLsOE7Zbx4rBZcSZkVs1GOl3+rNtn1M43ki6WVvV+6UpmuX0OdNhgGFoR7WwdMq
28SNolubX3KJfngxmijld6+wAvDomrVRUlhhH98eYkGCPQAiZNBrmJ8mdmlkrGys
XcZKdYx/VJK5dBBlPHhp3q40YJOmg/tWfw8Am4E/C+9wQdSgZGxR5Qh3m53Y/qaK
vCBEyDkkSyA2okK5LpJIYnUNeiMYz0cZxzZ5ErJPCnVJJgC6smJAx1f4l/02o3cB
EKshPnbrCSxCahJM+ji7Dow4nZYl6g7ywxlJ1GRafaNpcxecSuMuK2cJHjuIg7xg
u98dwb15sd2NWWBahdcM6I471f7z5RoH3wm5oYwcR8NpteTt8+c/8/02WaNjwI/3
QpUWSnvqyBEThxrC2sWh3j9JjfX0uWNuD8+NWAsar8nQBo98NnQwXLllN1OaIniI
LPdyjProkVGDxezWdKspkZ4iCqb4bzKknVQCJT1S2Df/rYZTNhckV4xch/z/KpZ+
apc9M6SBKNnNZ/0/vBIdQVa/uUtOJZsMM15kYJMa6CR8p0VY7/ywTc3RB9F1pxD1
9PkuXnkRnrFmSVIvVo+K4pjtWr9mJ6lB56KrqSA4qSwp2XRh4H48fJ5zsp/znklL
ou7gD5qTR3Oas0b1KR3cQguk/QsDGzzeqtFvUZNo4dn2GXmbXPAmV4G+Nw/ld+I/
MLEFsmq4yum/4SzuuYNbZ2TkcrtD7BxfW88mBAzyRek6OMjB3kXCYDgajprQCvty
yu6kHgMILOrPGOFh0v7s0wqE5zQDx9N0exiFYXIppuVTfXzOukTKDuBqXRIktyk5
OhFPDkyAxyPkfQwS9hkCDdCo7e7fklHjG+8Kl53lRCw3ci9VvnHDNscVSHei8/b8
KcjORNwK1S647EGlmz6J4YbnWmnoF4q7fSbA85DgouHQVM84VYdkdBOVQv08G6Gk
g0yA6ofYAIROeQUopPCfz5CDwZ+a6sHNmdxOuGOP+VU2F4djoFtfSLevRsFS4X7L
vqoO2Ng3Z0nFd1+jxikA0stixQbHCe44HE4XTuLLkaw98i2BccpYZLTSJ3LCqhF5
dBer5Hncz4tT++XY0bOjt9dlnpka5B46/h1MxXavCDHomKpW/yN713JatW+lny/w
yduL8yp8n5x6m1TaFpJndbeqt82gO9N5Ufnkoxeq50Gu0WekUm1rUdFcZRQNvdq7
7xHhIJlcd/Ol8EYlIGUvG80bMfSeZ5lwc1lye2/szOQgWxS0N6fboCXUcAGnUplZ
AaWcMZCkzhe3GHBexkzupHt7t8c9TI2xh2uVnV2J8HYlEBO59iBigejZziioMcxa
6K0SrF2IhnwYTP5aFToSVGsKrAFaAkaPWJg3gaUN0ccQH0O6cwCWVmBbwC5eXuUr
Ottz0pwCcjq93ny2+Hn8hsqKvoEj8Aq84Cz0d/g/eyKMb/RvjV2dtcn0fbEc2ppU
r655tyx+RhgDJX5+w18N7A/pi7JG07ED2HokSeVFrVjCykPwwiPrnEkYGuSpgDCr
7HY2pGBUTpw0aOjSBQ1EYuRAnkGQ66eX4bBe5Zb5er+Yc5Z+PFGikLNydArvPkMA
5MgI9DaWVgcpJ3A3+vswjon5dwQ4SNH/k+5jwOJ762k1AJ36345EydDQOLRMZZbX
jHBvYe8sFuPXA58qOZSIm1U6Ga7DRaezcDe/K9KpZzY3WFKZNWwcWXC2ufFbnlIX
n5Gr100uEX1REU8yqsF+0uqRBGTt1XMwtlLNsn1LCY/7wn/jIDYhzN08lE8AyY2f
fIJ4xoKUN4IPHsf2CcQS5Dum0bnbZu4l85D86iSq0zk9dX1bFoGl2byUqmGy+Vvd
qIKoAIVJVHdgz3qVZ9Ogo9SV1FMajoY1qvSdpgmB/SrcvP/uHdDaqbCWnSkKZ1CK
0rZmX1NHmXlfCYbLn45UKKezGilITdH+PjhRexkCWFzsHfaCL/pLF0bREKLkxtlL
7zYxqku3FFUsx4FDxlONWD+1Z6cygyn5tCcG8AkBecXUpXxRo8EyqIncH/haCiba
s0dZHRHMudtwRfKlexxoKC9CA61JruIzYeGwwf4AiPsCARbHDWFI2KwlTN1QFhY9
loYmxER2pegR0M+592b0mma139AeKa2DdXvEznVDGF3N/6wM3UvAzFJOw2xTHZzB
AaYdUhbasCaduhrCC4oCOCz5sNF/BrflnieAB0EyKdaK5J65rmvepuTcbEuj8SA+
ZL7jI6E2QfMvY4tzTOIhWnOPCLCfg1zM1KdB60WcarN4NwKlKbspkF4475k2tTwl
wuUVbivoPcXSzzhBLw4VWgLlBm34lZQ+drAE5Q+0mfkdCK8UoxUKC8KtZZaCDfBw
nqDPC6htUzD3/C6F0tkJKdfboZicxWpO9mg8735mWMC7EqqSsNxIpeiauAWZCTxO
GCJiZMHXpX1TFu6sZvGc7roSCc7glmE+eF1su+7+PuzhVE3eFMwpR743tUH4jpib
FpmEumvZ7ppjgxtjXVnN0V/ZgTy3yKCcFUKDfyOvE74t7u7oce6v2enSsWntp+Iq
JNPCfiGy2hYKqwBRQdDpl4PbxqKWcN6xolMdF1bjv8am3jOSeIRu+LinSFHPq0Dy
npCxKH/iEn3Yw8/jiCM9guPMvfXYkBUgcNC2iQwODAzvBvUySYIoOh791fDi2k5D
DaqXi77t7FBmeTsDwM4ZHMLjTPF2lM/GqP7WkUYTlXeV3DvqSW7Xt30gQF+RnTMb
aInRLAGi71T4stNlbrciwY642XYzjDeg69vyod4skDuDpXpiIlrXToKKdejJycQz
PZYNMdTtVHecY+NnBvqQhDlt9BBsInkmwH8kmXzyau7f25O5DyHrz834zIZLbMXp
zCTom+tG0wYlSXG1R1rpsIptSSIsu/GWHA+TB1BVGp8liGq4DMKdWp6dNm+t1l2L
3T23h/nu1mSuAs84Q/nCfkkiFDZwxG4PjbFiZ3vqJwTU0/iQgWiqUGw5h3Ke0XVs
AEvaHBJmfFdV+Ba+IJy974jj865ie+gg/ZtjQmxWa+VcUfjBFka30C5kA0KzikEf
77LWoZ90sUSV1ta+1bJZDNXi63eDBtoiBz+AuU8jKrFYMP2c8Zl1BzPv1I61bFSt
vGU77CBOR6LQPLZb1isHXDuD5thw9sWwoHO62+h6sIKEWMkB68ROudi4XULYiYyS
M5MuLwDCxwHCSuMblU2Z9JpO+YtHAVYzWSM5e4LUu54KdqmdUoi1hqPwaZJrrbi7
wlVrVFmwshOFzr2Kj2rWCYB8PRuJSHEDDfoLN4gqOSnT5+DgocLWwgVZ4MzA3jkn
HeRK/CfIcpSrVdTOYAE47kXbqOB5auKEOQ7iieXfTcpXYVDnvHfZDcHXVjskXHnP
KxwBAWYYf42cqEULjY0Cs/rKZvRFM4cpSMqX4/3P5QmW0wdsCEo8WfoBRP1h6HoJ
075qjhSWAp20WNaaaItWMAXptBo2/jRz+3RZYUKU0j4H21p7EdexXHTZ1IO2rTBv
uveTGIFyugC7B4lEU2MpXeCwXzICtE+Ylsutn30PPmE60YjFrNR5Pomr7qwt6vhd
9C+qMH5kfS0qj/TeDFgSuLlUB/AykJ5kH13lZkOPb6mQRNHfr/6mcsl6CfFrTa8A
9fUaw3z/YJ+5cBr1C4DZ4QVbR8aW54oH0yKt5sYBUkX0+oh6dGbizH46DYpYIcJs
XhmPwmhW+G9A1LeFETNJ7ziamzfNW4MUUgHroWu55WNNiSC+mhtilZbVo2QDHb5r
mu3PknMZ5K4WEE7z0RZuV4wCpjYH7hv9jJcu5H2PWwUH8LlymC0+Ru9na/FvujH0
dBF805NTqUsdvBx6Z09LPyyGF82irynx9F6VaXkAFOxwrTerxsKTLsVOjyFZIs7S
oHGdSwEh8SEKlPwXc0a1OJMb344HL5AavsLk66Q7ZgjejsAQUIddu2b1/TUcYN2U
iyk0N8wHMpAyvLJTii8h/mr4DII+n6xUZ39vJSk6s178s8HawO4litN/EFTuMedg
dLLSpMskF4lw1ak71InQCN9MwiLZ/EK3WTyTdZPtJFYUquC82QVKGmEy2JSVL9/l
V/TLECNZVTeNXfXaVw3oPLl08HQXntZOahUi0gnVDXm0vtqfURnK6D1m9iVsdu05
BOo5/pxXVGBQ1YeWjYtoFOjAN8ZXsEbYVGvegak0JoAMPr9DpGVXq9iuZ9knjQDL
RakJolixtOGaWfhCQHBS3LT9oaKIrJepqfgPBnBCOVIaiik5DhvnhrRru5/xenCP
ArWop+i4ggsVVHIZUtzodP7gum++T9X7KYY2QzPGzUfRVQXSEGA4nmkNS2r+adJ/
UOmT25CbRfwJ293sFckQKjn/q5ThL2PhUbR7FRfNT4p5FN+g36JH19HElmCcPn5X
rZU68HHPuicJGAwb5xgAKzD0lW0ZcPBXgk7jhtnMMR439Pm31vEiip9kuqYGpGHU
go8p07rqRXwOkczIFC9hXE8UYObeNTWheXd3nye1oIDkmKTtsPHEdQ98BJywXnsf
FPTxn66jW9RoRstL2A1LVZAgK30NafZrQpSiV2wUCtcYC/kWsQgKaksmLATcJDB0
m6YfoeoX5mckzRoieu6d9jQ73EXVT9ca7s7TJO6qVPFvRZ0jXgsyKmiCygzPYRDm
+fJYaKE1403AGZgjMFjX8/Js5fnXbW3HL1KuMHE7twj1EBOWd7sYoL5ulqn6dnlR
t3mE9yK/WTybj00dmMDx2WWpDk07VfboTeE2qTl5rRqwmUslUq005AECBMTSLsiv
4heh2fFuCXQEv9dJozWbNDPWj4P8Ao6OYz4/vEAdQKed919KKK+vPLtbMJ/T1d27
BWIXGb1rNrq/RbmJnPJhYOeRkY2JR/rcnCzSeobRRaeBQY/KCYqe4btPZ2WyQhyu
EA2QkXsbHGlQpC7JiGu/k6LxSF1fb0T48+GqiiYDw1P4Xc6cNBV6hcpC/A1Yq+56
Dhf+wXf6Oe0TZ2IGtrtJtBJy2lNMo1pbnfPOIp03wsB04IReiUenadV1Z7ccaLel
5eYuivjacDzujuRRFq9fvjfkCfclKLoeHtc2oYxmmZv1PdaWhNPHDxTNiPQW1tOG
E0nP6MQ8ZmIaJZBF14Je871R688b5Eva7XjYXhyCdeA9tug05jR3/RjnYr+TDp1H
4JKWCvzU9XvQRxhzagxXRronC9pefM1tPFeq8OySPYuDi4s8yYhvuYNfQsdrFYL8
4gDUUyahcBhqYeV8w7AwjeqJocUR6lLYkg5JLkpDYg3j4sSt0IydA+UerOw09tXj
Jz9hGmetMfBkFBF5hDOVMHtCNpp2ja4zkNATPtH/5Qp+3gXtk82dAHkdou2FlF1J
DxwV77E5Y0jUkfW5MMEIIG7gm8iQ6t4jIZNpFxJ7oDvqNVJ/+0cvC/TRp6H3//mk
W03PgN8TO6aI481iUsB8/gGxG7gt13zX2ND9Zg06tQo3gXC0gwp0uQKin+7+PNML
yvUPt5EGmKSUZWg6GR85K+gT6iq4f2HzgVi0OGxknhceYZQ/ggFuzPgbVepnPCsK
YozycaofKGh2LL+Y4C6ijPhe2SAj6IBnFBXW2qFPiwmGvN+BBTGmKUoinSrGEG7j
icUiClzUGHzEEUnb/URwcNQqX19usH2+xlUBj0VOfqylnkWgD5Q9LgGKB9ZuL3++
I3xN4wtP4gyXwlFLwl1ctKzLuVt45GcJv/ixrYMVrZk673NTav/yWCB/4cISkJNx
GoAoszAulSMjl9anYCZYiXlsc6FX5hP6OdySCVZ+743XyA+dea4V9PGMy+FnLlC6
odFUNHCm5xFXXTjpx2m76kslFqfqDzKS8OYU7cjLQgd21tDPyZD3BIygmXMRCCwu
O7JJaWp8myvqjbnggMfLHHsyps8CKr2hxEO83EYtY8A6ci2TdE31oUkXN55Sh0Af
Lzg+TccjPEfvU0x7+wUrHBLFfRGIYodlA2EuwCZ3bL8IWIL7bBt7EOYt/62B6Gta
3Awvx5J+5zhvjNMrccyBowuCrAR4FpyI7zZZmz8K5wdW0jf12LKupruGLW82rLtW
bhYb+C+SGaNfXGRnmOEI6th/ieSr7Cs7nG0UQUfwFQNL2pgTsD5PtFcaQWdXoPH1
3rcCJRvOGPj0dKP9COq0RKxYY2vPEwNVjfzwa81NBjMcNMdptbyOBPaGVmNVkfJ2
GrTkoy9RzJT+b8wIQOQHzb+UjtD338Z2MO0TzHnfADlOUCwV4fEW9jhcGMI/IR4d
/vC4J6YcYXva83HDtCpg3L5JQoKiijh6ZxG7Hwf6HpcCUDpysQNBMOXBQpuXB/1h
mL+lLYjJm7ZG58PFdSMFZyT2OZdS82nK2KQdp9DFU1/NKTp1Q9atVhu8vR7qVmuN
tPVI4u2TmPug3KOzMnn7EE/Z5eXqp0AhG7X0dHU8vWUbHbRAljIUJiTE3LoPf/7r
WU8ixdx/JnEtTlc3iq2tG7aFO30TZSd2y/Ei10Ylppv4jaH+lb/7u1YAH3zPXrdX
Fvr6+uUWMgoaojjkYlRIfeBOEjV6Erk2zyXT+IS4g9m2v6ecxYpFggrpUSz+wQQ3
dOjEl9N2Rry4Z89e90ml6THAkctG+uwMvRgq5micqDt8RMkt9aZIAEqAyztOGur/
cSksQMa0pY9M5eo8zyBgYyfiWpFdaJQiFfPkJ+Db4PNJhEAX7swrr7eGD74uIqcn
SLo3dq9dakZ0RZaH28dw1yMOA+yYmmL4cMOoX01R8hcKlawt/qkvMSG0NMTitchO
ubBE4w5miZL2qbaGT7EF3e2gOK8hX5fkX7mGEv1CpqTYHDa2R4dEicx6uwpGQuu2
6CZ1QOdi7dbp+jr8gPDOh4MzSP1Zck1Uy/EqGd2RXdcC822N+GoUXt7gaBrPllO5
961hxkDd42EZ7GFSeiRFM8k8zAOZMnoPaYkWPCcWrEhu9m4lkFlNdf52Tw/mJf4C
vV3Mr6BuOOoPvuSLhsJ7Vto9umAHv7mWfCp/xoTR/ZlXkpNLyJoXNO2Nyr24XCYY
sI327VB1MtH3xE8I40XRnQlcFDDx4jkTxKOsZz8syZ3DVXmNAAlTG7o75fNVW9vl
QKU1MN2Bb2JVS/zwrUtBGDoiXRntfCXzuHVnbQlFrgUTZl1eZjG/VNey1BFE3Az8
j6o45Vhr152KRPXrCIS/Rr3XreC81M7Z4ok9BjEKYkACC6RaUAtRa6kacEVDslR6
Y+3pMm1S856JEuQoDHMAwOfEJQ6IptGLnWR9iUyaeydfN06mL/AN7G4iM6Qmi0yg
1HbUJyNjPVXKNxRHi/t6IYwd29hd5ds6+MKvC6qlpckpInLtsBwsy4pTzu9s6Iq9
rPiuiga6uhb6CdWcYhzlNzo+wKp0pv+sqWLH+WGPQBb4QLTHtzT/XM7H6FeDa4Vd
bMcpIQVtw7wHkJC+5Ao7TpCbC05I59vokpoSvPh3Vu+Yv6gWM0ztQZkjK2iS4jWF
iU1JCPZJfLJ7mnykDmLmO9EkeUHSeCb56aODUSJ74DEg2cRvyZxIuCxGZdhseAea
YYV+FXO58O7GJBK1Up/TSqV8b4B7MLVUPM7Pm7hoKUY2GOS98l/PA6frD8/wxW4d
MVnP4pGPmCmdWxk3UZckIkrpBtNLn/TK+DHHEAJkwvY7b0Nmo1V2qEpi+cstTNaT
QbJEfSeQE9IS13FWfAgpgVdrO0QGalDwxgKLUrNaT3NCPSpjH7CxyRRmAVHrFkD3
565Cil9XHdpryDVweioziIkf0jhDK41vKctou52DrZy+yzXxKBg0Hz+Wq6zZONLa
OEq6fmD5FvDLhl3vZlHtfYwEV95PHBwSGKpTgeee3Zrgh9wX+wEy9sMxJ9qYYZxF
chfN+oFBULx4rGp1f8LaXRS9Mlx8GkAeu14w9mIFQLBXLmtPzr3orctqg3Brloq2
zPsrtVU1V0Ydi+m2T5cgu+/6BGEmkkzrvLH4AYRc3EThRNFvk79zJP1neOtUBy77
lgeuy6sGR5ZYUeUT3gwWiwSx/WiJDd0XyIRSbnWVo5kcKJ7vzRzh4a5VApVxhk6I
1B5uyM7MGi8VKYFaoi1S/RQtTkVyDGiKLrB1uQb0N0GHi4gxEcEmUpprsPfiW+su
UPKSWyST1XZiY/vjFT8bP0c7hdiFBiI+eNg2VXSx38biNCGG0n1QKVjxDDwiM1Kv
TM4uu4r99ZY302EB2Q02WBWHej1dDl3aapj2UzswXOxf6VYIgRMnpncTnPUk/8ch
hlUSOd+fW94Wl8TfV4D1spwbGUWu5Klx4c5LQiutb9Wh8IHL75H9f0XkQ6BS7JoY
TMdwAwOKMVFClHnqpUprbfoR1iUQEX1JCTK7NO4p58lhBXhmOLSvFs70osEAgCAJ
KqNuheRPpIlRTmmAsDFuxNfZMpRiCDnHJvAI3LmP0ffuxKamZvkpkfgz0zKciSDL
a+wM9rpAoRMbdvM0uIJqKCx2nu/GBU6XSiAgaiTepz1TsLqRlDWJ5nlCTJlc0hhe
FZsCDdgUSJcYDmRtqYBDQv5IT87V9evktkQ0MPlUyCPisv7iwvqPKrArvhse9sR1
wjnsALADmBEU95Xw+JFTcGPywmiHcbNXH4U0x4HBP/wwzDmAPfiIeNnvJm+9wl2O
56A9OfAS67DF6nMHgEnienb2Sjh4p0GUsL0d/DGLzpXoSJ6TAco8e8hOgTAibIgC
TY7Aqstg1h6gH6wedxNapCh9KoKx3UM82C0oJLjbNAikswfXMf2TLSLLJARqhSyS
WDDEV28qe4zJRJIKniFY+OngfiQ92ohb2Uk538cibxpL41cTiwrSJ7TFuP3Ok4mj
MFuR6Mg9H6U0xV9eXTbrfoodTYQlVrPnCNz2Y23cZWUVjefwIhyCr8Bhq1YxxYJe
ts1RrBErr3crrpalYwFXBhk5EGFV5YnsXe+Yt3flQCKugA2Vp/zKP+IHbARux3Vz
5ULp6CpaEtPlbC/J8ZZDpRPOedpu/nrdAkGcefRIJPfZH7Egm4Xs/ehvtsZK5KjC
B8oBmHxxaO1y5OhawyuRcassEDHxMWN/ZCzTEdQAxBgrWmLhdr2o5WKSve9hdtbk
HEerzoLA5EUfNrsXD38ssvReBC+WEUHPdw+aOs5CruqGgFX+3an23SBHXxGEKhun
qIbFgBxMQT+nRHjLzRPO222zUijnXu4X/FxxcjQWCAET80CdrkAlit7zZkQSuH77
0ShK5tzfGgPnHWenapJIenNCmEKExXU+Mbzr8+jNnJgxY2RvcTWFukR7HP/BlM+p
D3Jxk8TyzydjY2JoTUWO6/lI1ulp9xyo48iSo74bpTZ+Bizh0FxMnUJvVWWr/O2s
9Cx7eYHDpj6gq5FGMlDq0ifzeouB82L4WsZlUmUT0U2lVJtn9hdz/zG5lWXwV+ju
lLZyBBkP62mFEQNPAhqkPA88M/cKkxrWOZ8RVWhVKled7HQcObJzZy94sC/KdQv4
0VIwb2mOnwWN7HlEf5XGe55CsWmHtZFRQ8LB0Hs5liGlKnzwksSyqonF4EeTdoQN
TZEgEs6P22fsIjq8d3okaHARuOWoyt0Q/uqqm3TCtrRjlDgqI0UatPiZYhXcoHjV
Ymoc0L83M9Yr44LJfUWPmzUK3WGoszX+0ulK2dL9/pLpBF7lczqSjGJkbfBIz7P8
ksCZLZxcAMpufR26ze+30BkHgpbctvCLpG5FGA3BJF/cy2exgSIitX7LMYdxD4Un
mqOiq4hf0J0ILB3+l36Rk/vjrO3Hc4d6RVgzFmm6d3MwLB6X/03FNG1miBfFz6Eo
2O6153jbFQe4aoBeExlrYwvjZ9vsbWQupVqmhG9UpYCKTYtVQauogUVA1vDtz7E0
T8uSlTTZpKg2UW9GTC+/4ePFuM/n81OeRvKIuV3wsVy/YaWStwqqhdVHq1wdxsGr
koLIHzyEgRXUjbH3JeEFPGjWF7ZmmcW1SV9j8Y0sC5ud65Cb45XxQisAOMy4Dxk8
SVIAm+bmoT1gNEFRRonYHhBkWvkhG9EepgGLCxIUz79uYYuzz9Bfy5F5TOFfs9Tx
lnivLMLDoc/Lxu7HCRb8TSsrg1lAvfb+E7Ke4aiMGOe1S44ru0lYmtIzCMrz73rA
MtgBIOtZTRW48DS+F3u54RCAJkyFfXezwkxiJycuMLlqzNcZ5ISCb7dCjkXm8HoR
F364F5la1Zm+Whl9AQYdQ0iA0FXqzY1TpKVqNUab1KdtBKTIAHQ1KLcDFzFlktI7
xZZOKQeMydJfk6qP2di7lNWByO4sNpqCxBggcnz6q7FebG0EsYXS7eIX9t5JBd1o
KuxvAezCjeAZEjE1H6EUO8orkFQNeOrIq+xtIembUKaJqeWSdZLN2DrY8EG86umd
oiknR4/yLTVY8RnRAAx6cjmZJifHOT8X0xpkjslAAm70mG6lpfw7alLbsf/G+ZSX
WLgRkjSMhPqYE2UYbzxLLEyn/lp7jzu14MD0hB7t33zY00J7jwjYYwLpeB3qIHIH
zMd5l6M1T1HTSlP4rC6jk9PYyd5LKg4ZpKJxN94qaUOmuO3FlDnZrktdzYMYveux
Ym9Il7OxGVApaA0nellTpXJmgAcLF8KvZ+M7jSr7EY7kz3IQXWoB5RXr+u+rzKZ9
jSaUipQ/z6Zc0R7YP6VTAZ3EHwIM50TlrZudqubJyGwaIm5RzrhkaE32fZTpUWrn
RfbDfc+klb4Ay11WC0ipx6xM+Hz7P4wqsNlau9ChwQMGFnybkfsyY1JEjiAE+wet
YbwLioFo7U/Ux4bESO6HSSAMU2/YMebHzGvRP5MjfBrotx5Rve6DLusC3LuRG9D8
Er+YNxEf2YLaxqMpcZsDLJek9hiE6Rf1IwZ8sMydtKx4NNkZnTfkYuPVhmzObgO9
mjeIu8aMTqHeciQW+iYyaGow+zVTOygGlZbB2OE/agiyKYFp8RxdDU+qsDOu5K1B
MOk9tirvdZxlLeiueUQdtj7bTsc8YYeki499ErJNE6lqzp1hNjuQCveVxXr2YU+O
hiTUq3AZrWv7btJ8Kd7L5VcgWLV33DxssNHWyJpuapv9wQlgv/kbrqKr1RTVdI0I
JSlDyhvdzk2uj/iTuM1EfxfOARBywrEGIexrIRyiuY0psnZjIwU/h0kPTbfgWiS/
ddL7I7h/SOeF6h/RKmX4e3ILGA7FIXh78LnKbcrQd32z/Noi3pvfQd9Xq3QLtyAH
9ZNKQP4HyW/s1AnscUeINZcC5WsYTWTUvCgOh0H6t9kd4h7HKPQXdFaph9OR69Fh
kstsBKnz9GSL3sHg7GrPHsdrwf0FZ5WsZZTNxSRvZssHipvry7oImkK0p0TbXJCx
qfLL4gyzOWDLnK1W5SuIwFk7kx8HqZxhd129uqhZS0UNE7kF8knuiuVrTnKhsUjT
IO6/9iCd2iO4FhWOf+BocPvk+7NNHsga59WepTlE1Ug8JjLAOKpyE9qGp0E1v5Q7
nm5WjvsQqj9cAivmeBQCZ+UuOZ7V6R4veLXq9nw0F2cEyNu4wyfsWCqtivqxl9cV
ktnVZg/r/HcjqrxS4QcDFwc/Ne4R3lHisLHreraG1A8eG5Cz1ikCDhjVGpIaCFVe
4/mDJ5/HgaFsZKnqldaIf1HcFK9JQvuCd0UAekC3442IN9Bc7fwrzu7IJ8XfrM8/
fGY/UwFr8pWPriQ7yQQ0odMEShvxx6vuyCDDo1PA40VUZ0UsiJMFLaMf4LTCzaaI
BZ3yBy4oBBJAOrzUSyrkB1DfplsYLBlcr9vErim0TZHVvqf8+B/KyrqeNp6fL1Y+
ISlK2un7QpVKYM8rIWnQxcwXkNY+4fiR+vP1PFPBwTsFDDV1w3ToVV5xdMftUAYh
u/WCvXOrfw0lotBcGGXl6BbcDZqpkDq9aYvuQ5zkD0tufRaX8YF0CggMQr2WB7R3
KcR3rVYWmmfOwx5cduMlqRyoUpqhApPuoUoARVE4tDkMY4ZHnxea8aWDZnXckKIX
R1Cw9evyyzNM7b3p5n1LiwWvEKTjPRC4DFe2P2n0N9S7KPLsWalhLfaRoosbj9ok
AA+J0I1qMlVN84dQT1vtDffv4U84j+u6zcRRf4XE68Rp+K2OqZ2HKNiufE8T9+h7
W2QFkvN5YjhyD3ln7T4NX+vnKJ7MbW/W4mDX7HZyMpjmUUEMadVJzXkSyRwJFQlI
YXNm07MW7yz/CFppSSt1MqOQhM8E+p7ITBbBLnF804YJaHD7BsGh+ookIUJ8Yc/c
0rJ4EFJH7XWIL/WGu7pSULyDmnb0kD6W+P4VnQRfQf2KoaXOYvG+1ZJifRu4sQm8
Ob8WXUzyBMuKtM7gPbErPylNIz0IIyn73O8us+QRYKRENZafbaeB91BrEZEMDyHa
GyMtmwwOs3IIZfiMzI+UCbIzS5HP8by6pnJh0uq6XZCYFIxthChsof+5Anf+qeMS
BE31QbSzA9BVZqSymtM6Y0Cpk9VU9TguEdA/eK0OOlsLBWSfy/z/wWNgS2YMOgFP
c/Gy5xP3ssmO6lQwgDcka1b4T+FVjiWSIO9pcxsoEiDxzOtiT7GrW8O+b5pUJiux
7KCmhuMtSYDe9nSPbj248d5NppJG/zEURDmERmZzU6RQXzUnrwjBnOSG8pPX3Ewd
RcmKcPhfNgoOwKtpKNC+JSjGlJVRxEXiAn0KYActj3+zIEkbprEK1D6UF5lrR4wX
QncHORr/QppkMFKqlZneuedDPq01jCzoKryJEV4uwnuKYEHl/TdnP2MgIFOjOsFy
MrPDjHT19Qpy4daYfWtcLC+gJTOzi/Ptg2Wvi9kNkJaBqXmow0zI+44vMUOC9i9n
kI1Vky6BiZMLpLOUlbbrAjVTzgrfayzecejqQAwEPCOM23/AzqdBaf9MCsPKhyki
OdWdtbEk9pUVz8XG/aUkHcgDCW6ZBxQWh2hvgLORQmxF6H/bg9T9HLy6KPl1nj97
YNoKDi2z9TWg1E6vrr3uGxgIOHRRgShihECzejw+p5e3xcnig1M3CRzoBQ2UPMcn
C+Cqp0a9ZSbck7C/i9fSS7Yg+7tk80yAC4C6lOPZOoQxPji3ZCL57Qg/w+IHDGA+
Zm/gQuYvJeYgjvMENUH++xypf5ajGTulvSBAH++Z7OH0DMVh5/VVAOAe7DLWQHl6
zsJlEswrSQ9LB2nZ8MYcC4z2h1RSUbeucvHomA21mgRgl6JLfYqpB20aiGJ/kkTn
lLu/49m5bj35MDrOso1jbOmLtXuUf1KcZdznRXq3L9xDfEtN1CZN1GYLFWQp8kRa
82SWy8XSokkhpdVH++BeUHxwfPhAjg2SaPI5cDAW+1eHnLzkcmixr0ToIjZpkAw+
r/IotTt1M2k7xawjtnoKm2kN58KBQk8pZg+EP/ey2bW9nif0NuR41JSkjqokLpUP
qjzl5HDKBO6q3c2boTOB1co11nQURdjVnpqlX95mWmA2Fgq3piptEYTBnmbIBCHl
ogAbRnceu2SWqTqD2eyhFV3sgv7IX/JecHrQxNmp+LOrjmumEAO1Q+cv3otjWTYK
rUQX40C+lxwdvScxw/yhmtIBH3o8ZLBTL7yAdHikR2vff+JKM0RNzowGdcN0EzMc
PvYLRxUaGeo332wrKtAv/Hy0OtIQsqibfQHT4/op+Y1dLsOu3D2H3KU1Seii5CYd
qyXUixysY6ZRMRT0vqKFRkG+FIJelOgBAECf5EiUTk9ILe2Lo4y7nY6ROiOzjU1L
UrfRrr0aqBggvcu1SHaIWEVNP938uCBd/h6q4IRe3qza8OtcPMEm+2U/s0EP4sVA
KwQog4gpJiGx/ySxf3BD6m5Ehx/W8Vr4VGviGHtbz/AMHwLtR0z9sxYuUwIgPzGb
ZS9xJiOojWff+g1ggMCsdixG7GU82GLXKga5l0+76nwoJVEZIZA0QMrdXiZ5uGy/
tgQM/JeqBA5lGN0zlfWlUD5eP+KUET9biZ0qhIh7z8lx2vA+9RzEEeddMJj/KcZ8
2rTGE9r2jJuiSbmLYhQMqgq8MlhDv7VsRGW6QCNKQXcf7MwVLsTG8Ro8GL/XkfG0
+MbQ6qTa+KKZ7fveZy1PzYje1LYjzxAk5K/JGtnUOgR51hlBFcSBSYQoGxrB7Sxd
pCBNGpEhidZTWk2WNK6Bw6PDmR8hX5ZBjkh01h1sZcP03SVpFfRoT8LjNj1bpZYa
xGU7UomcWijY3KTXpK50bF42NhpnQcRohttalYWTlxT9/021itWpVXwepRm4+0bn
C3v9+61HFVvPrxacXe1L/53PAbiQUecvdhkhH8mu9dKd6NqA28Du6OZULE/OkL7F
M7sQ4jQfca1a2R+QXT9ZqoekXvds4ZXaWvDeLp3ODRn3CLpbJthiYelIhPomvsip
PKgunusP9Qf8BIX9D6AiC6wzLpSct257BVv73R99N+zfTGk9PIooHvxODcdvO0XJ
/oUC0tSp4+0n42cI4YZFHsTTCOIy6uTOgCBJU+nGHz4X2Pne0vDiwDaQn+X7vead
K7pG780S/wctKdfrLPvQwaNArveuVj5KMOkT8vfwr6q1xiFoZf22Hv+a90rRAyad
K7Tee1R2XqXzobV8D3FdyTVh5tZdB1oh8tvuHvfqasWpcWAzIr0SU2zkvvnuPQJo
6JyW3SOS9adKPyH7u3LSlmN9d9DDMx/1mNj9VyuhV499gyD245qTHn+TyR3jlUMo
nUxlkY/Ic2vZlOTQC9NxuDwImDHFm1QE7x+wynrjPvzIzgb0F0WGtWTk+i5Z/rb4
o6UwqWgwJIyFPFhlJcBfH+gHyZsicKA6XHQ0GGWvq+jdHslvYVVr6yoeWoOHueXZ
bZnASIAtZJPINC2E0B4LsVQ+MubFvhq+glksd0RrTssxARyEcx1lYlks6k1yco/2
HPKOfjJcEjqE4ySKhNIyEYR2VzwcefwprFPWOYz9xoTIbR0H2OxKxPNHuPb97+0y
7AINCEW1oQ0WDTlEmp+O56H7kvS18AXu7QBnW1+EGCGcTvUIWLlKe6LTPWrgPTst
xXNozboddQoS2qdg9bN3fje/oK42bnF6084kgwXZNdFho+TCh6/oEpxm/zw4SnmG
FkVxKoaNED6RgEsBdiiQa5pOgRWjt02FakvfZHbYK9mRStYMb8Q/LoFKk328jUUl
HZxrBXvlwuY+aZysNnQG6m++1Eslg1+HV2sdt7hVmN0w/4Pqj66pwbik0jd3wT88
CTN7pz1O/+ip6bJI0rbWoDlFogNuC43jMhpxkU9SnBvDTio8eTCnNLHXenJ++3V8
DcS35IfPfhsPw8lwyWmF9rPLB8hUWHvTOC7BU39Y+swgRHzyGEdEm48rLovnaI0B
jzsuZYFl1yOsZQy1dsihTaM5l5PrjSL71gy/BdimPc2Nga7KujfBGZLhJi0C8U+i
v/xIcRB0IWE8TjvdX0z7BkofwNjCoSd/+zxYty5/kHZJBCHfaw4ZxPZb5JBuRYPq
rhWAUDQOtUqCCJSwpgsrVx6PT8DhlF3I64kcaI47n6iN9feMmeYcpfvDmPlN+ObZ
M4wUHae8TgWO0WdaSRK7ReKBcRvGTyq2EcfIQGMyiYAlt8CiKDWNXEXOS0F4SrZ+
iNTdvXL6oHKhUirgqC9g2l56gyvlKOgLGLMW8qu/zeyK+jtQF6miTrZMTTBJMO4N
SWShxEPZXMqMPAYufvLkylB4HEn7Tvbno2JwFaUaGDg5kqbR+JKWKIwXVbCllSlB
n+GLkaYea5sidxThUBuGW5xjjznb2DuKP0WHH6vuuHqCShFGxvDEScpyA1EeTEFJ
hAmH7Pb0uhtc+RZrx4x+pGDqkdi8B+AmuoNqhEU9I5QyQtHObNkdcau53NPELhnB
VvdWbYnFTSnec9FB4Jd9dherG5jdgTcJI+PO0MWVfpiQNXwwR+u75JuhSPTIugtj
E4kAQG+29TGbqc1UKE2W9TgVmgbS29U8qkI9e9ANZlSUJzjIdTxyEB3qtmFa0WlR
+fwHZCg9RPbvagkjpG9xEfXCUz5NihjOIHS0AnkCbhK+05q4y/xtwgC/PjGhh/bq
xsQvNZ0OT4ARndpYTF97PGrTfgm59J6TqP76CY0MG1SpYatlI/JKHUHvQXdulosT
Ri8NOrZXtwzb1+6UkkQqrwauyAz0hq4Cix90VOUtKSIrXdVNH/PJHvCxQRNSLE0K
cmPT92RFVXuA4SSC3dUhtala7E8RId5uxg+1dNXpoapiHcZmKMqsAjyjEHsVsOY/
bMIzpuwnBkTHXVpt2TMLdw+vdue14qkYjVleTcEaKzzUpqZjQzgD1Wf65NkJ8Hpi
GLxfqNAkcreqPPhehc8ZC1CTBiqcoE6A0toQeF5HkdtmUL7GMfcUoF5CgURONzVA
EJtZD0sBpksDyLrkTfMTXhPMenb39zyL8Xa8O4Dofzq2o0PA8MqxB2nUM/B/ap/S
CdweXpKgo0eiYsVqZygeE6eQ313srAnlwz5xjCniFrq6R49dBrSHCQwV4TeIdDqr
K7+1hl8Djr1/j3gj/4R/tKARRf7OHCNQ/NA8pzeoznDsC4kkyJEmFoXGPe+jE6gm
ii9bfhht+EguZmqVfaUU5oeFkr4Bg1g7ebhxHbenJwFTWH+TKO/X/F7G9YuP1/Ko
Ow/fcafTDnsb/1Quv45MlnXCNIGySAclxNibDQJcnACOTwhFdC7seYDENvW8HiQ2
pezcYc4jwemv9LPZ2lI56AZQrxEEp6NxLkEE3RYw4gIzOf1XCgw+xtBQVR50GyCg
mbIzihqCHKHG/G24gt0CvQWOeRNzkv4n1zEXtSApwzr+m4o3AqKEDqoF9eKVNvtf
SQQKcarCHcoHoyCmaVnBQK4yHwFO6f9WZCKK8gbptcDJpadLAk6h1krCCi6slmRJ
9Ocs9971FI36jXEZrDMNnFqstRQGT2/2Y8UdSvHYR8WVk9NEX1eHpB0loQsnrB1e
IXI1N/GNs1Xf8yqk1iu0KGbgipQVXVlmS9IRDbtoavtsgGJyj9EJEXaTkZ5DSQKG
lPOtiN1T2ICJk93QKD6NfWtk6KX3aG8m29dbT1POlr5MIlsISX5vEAYvbG+U5gFV
ya2aDfgE5LOYCvyw0otJtu5oONpcHHaT4KP/uxyXW9FFx0NYzbcSW214lPdHnPMP
RZPp5Gg0Xfyn7QngITK6OnSaGPucSATW4vUG7bLNtRvPlBptZwjBT+WUExUn9lXV
Bc8m32DZYXjsH4AGex9T1N62axLuIUSCfgDDWHdCviDa+GQoJFazsP1yNphDaN7f
rUteFZEj2EX7N85kMsM/ZXQgt4kh/g2hdOwKSr0r3NSLEwLP22l2NxcYoUO4IQaj
zfOKkIkNR07N4+p74KHCsVXaVf0k960WCVIiwnGbLA5rNwCD6oe1+hmXmt6Tgv1g
sZToR6sOB9hnjpdAA0zumIQ0ybFTlNdBdm4/TL5V0QMjsAVLrG3a2opbRUmvkFrF
DMt7Yp3C4XXHIsvX2V4mI/89WEASqmm5Z6k28dUt4PtO/zJMTvZW0OkzmH/aedMi
ZPNjpXpx1Pf+RdZUP3+DMoxQ9jg95yvUMfl4S1FG1IimWvKXavH65B/Wp7eOn1TR
vhjcz3zBH9PID2wxjMotSfSHJA3N1OGQr63PcD3bzoO+5709YUbFUqcVCJaY7w/F
dO7UiGKUAy30cwOYtzZvQVoYDT+keCbxt0cD+Q6YNVlfXkYSf/VYh+YFwNNckTbL
RoRNML9lKCSXaIhY59oAN2yig7GzyqTT7GGoJsdbNj/7roOREzuMo4cpip2/dv95
HCQuQfAXYpekrK7SjURLxgim4vEcoJ3MlwVFgmJtIX11ZpMqArTl+TrB00yxat+6
fuz2BPHyLOh0nFlJ6zvDjIvgJb1kTl8vBuR4Yp0FWFA7S3mWPWtksdolBbFX8mUF
WxfpctPwuZYZp19eejSc59/oVVKmiVRWbX4Dponof9QIwZ6oDhS2bmkOva6mFU/6
arIWwtno1Wq0YdiBOAwBziRKl9WD/v21BpquQ/628gZvaJtsYBGNpDOPtzvbOkgV
XYTW7vs5CW36vmZBiACPOyznfFzQXOvlVty1Sj99lROSNF/oc/2f5nGdA4G3fGeh
LwJ17cMrsd/DtzvCQ6Wu1vUkTyQb+t4IY4rGDXMVpc9eaRv6lAv8gO1R5QiOvxZj
xc0hBVaFOQDmZoH95RFEMto9GygVpNcVX6wan3wFSj5THmrdNH4hcw+tBYUylvFF
pgXAHabnudhUCagvVWQw1oQz30aEk+X/FgK6gGKeg7Ei0vBaHpMyA22pwNgiw3xc
rqs64oQoxi4lBS9nDIyALV5tVyoC0uwd2LsJCouXQ+BxKj4zxDqKQ7QjD0txNUf4
IoTcVPlSKArDD98lrGZTpaKoi+ZTf/br7TivzQlBxbqkcPFRXhFbGNzkYocLzk2x
asw1F1/ki+SjyDs8MuNGoU5AGM/C10H5QoNIfe4M+lTB80wBeeKkc49bhmKPElnA
Rwhy5Jk4NW84H0O3qCc7NJ86JULKavfxaq/yCRzH6SybBtzyEL2u9EQL9NotGjig
cp+i7fjdoKq4YYfSHfZMcCCANzkkXOxFhxtb25bEC3GxdOi8q7RZ1h+o/W5zhKlZ
UIwo0t9leyh0dOoFB8JwFHM1f3jXT0OugNHtUQwROFLE5MrIW8vxwQmnQ1JfXL/+
tYSNTucsb3WCH/vCuZARZQwkJowIxHJI5Q9DmOR1+DbG37Mrq0e9LCEQu+Wb+WJ8
Q56XdwFSagd5jPQKIJM8nlWm/zVaQwn42BdLx3/N4wredgu9J/zROAKlL0+AJZaf
G9IM47isEPLZ1WeAabUloVusjMzYF5gx/oLKbTApSf3yRsmg7JJ3eXiomKE4JS8k
b4/9hvFIK3q80vX35SdIXaeSByQappg7dgMeCdOSmg5PxA65V1EDIy8qtPPUUru+
x1vMyKxxqx8FfehRE47O2LCgG7mpP74Q3/Ep131GhRNocUyTL6mUbahbrBQAfmcr
TekxDZlOEkmRZyRJGw1IF9bQZTKKBZ+5aY3+hdvRl5U154n3rdvAOMMaUqtkN6H1
93kixM/sWgTHBAkQdg/cTXRZCNJKeTVqcdL/c6v0GvXGcWnsxvQOvWOxDu/IAZIv
pAdUn0PrLgYo63xMDoyKZoaQhklRCNY3tjgHBjiWzu4PYLszq/m3UaPewRK5YF6D
A/SZb9ObZdHAtxwUZKeL3wUwxVSvspdoqSCSMsVci28FSiOU1m9iOW2krDvf9GH6
sPm+qCosyCn9L3KD30L4YXpZ/RxVVC5r275gzkqAzgTlwTxpKjOhF7wnHZBOmVMM
q7YOy2xCnw+v47NmwrjVJZvV5YkgzpxGlRAa3/XJCP+d3jBaBH+wFnRDsvjLiIKT
OnbjQiQQuFUuD86yPedOdw4KRiGTu+mQ/pmHpxtJluaSbgQcuoWWPy1HdzXFtbjM
3TzMyPrFV7VSrgEf70n1OJtvGyjA9r9xyRQi3fodL02iShiCTQpaH7QNrJVcKeLA
19YXj+kZQXX2V/ZUbLyKtHODeAPaqG9VUr2AnkmXjWI8xjP7JgSO46MxBHxieePD
UetBgKwF27CcWDTTAIvQfBW2n14SvouCMxw95FJhFlBQHoV+1FRMv4UHeNWbzHRB
Pvbk0LU7UPbPyLHMrDH/LQR5GrSB4459z5g8OIU3k9GhaolKCe3F+vSCfriURPU5
z5V3C9VOpd00OKd/EgXyQwyI3KDA1q+GhDj6QN2rS49GVuxlQciHzRrP767EqPtp
5T5jOS6mMYBQiLjJgm2cHm5jazZbGCLbXsX65uW7CtPipPhc+bSVhS8FdL9cNyMe
e2jN08Cj6lQ5AWtu0S3J5lPreXzyNIGJZQNaQt8Z9mxBhYEQWMQmnWuczNKxF14d
NfGs2kbaTWuZQtPsZDX/lghQ1kVsZB3xIImeT+GA63MtF5vXeGMarfVRn+AL47FL
SeqxkBHaSmCBNU0i+YKtqnOL/9xwI8EpOvlCckSI5vGqE8pFuM8/PDPgsIkL7ys2
3/+cxkHZ8uIguZpZnEykZI16Nd6YsFl2KIEeX0X4KYJA1opSs//36uGo5msLJPye
X1b4SfZPTpWVCMVjd+3J8vKkIQ41T1nwja8hGPXyJhjM1/Nja9GyEZJUPdwR3dS3
xYT+q6LRdeDhTzh3cgd4w4ESeZreQAQiFg9PXhiF9PX3k4qxzXyI6msI0hBk+WXX
7CL8hFNNOeh41ULgqTlnKf46IApsMzyuz1VPkh5tbAHJk2SRkQzR9g07tG4ZwM3q
Ril7NFZ9cToSHmITtW/s8RgFKA2Fr/WCoLsR68nvxYOQYEPEdk5K+uft2rHfFZiI
edKhLpguiqUbAWDzML8gmaCKNwv9Zea1OZexZxTwiSv4gsPmhtixMp+Fa0yC+Oid
fVIQj5bYyXhWi/YCz925jjkBVhjUmf6IbIF8ScaAUgxBywHzC2cFo1fenhPnC/9/
gdO3uZJYnDuHmO5J+kpIwCtDnwiMOpvXVRlZoC6h2C42RkpjIKLmzRdnmz429Ok4
VcyZy2zfTSKlwXZsjiRNP1LjOot6GVirkX4omeTCw7lrpiXYB4nbagnBpfQMulm0
FZ91bVol4dTIWfhC4dhJThSe1F13EXVJN0f0eBdHWXobqksjenh7Rkls3zLMCW5c
hMf23+Exjp4zamw+emtWajeRwe+2M9pDkkIUb+yhrX13gcUXy9up6rYTzHIptbPh
mYx5C6xJCrIkbMDNC90ODZsmVXIK+NjwxgXK7igzWKppczn15pLvlWI1wU7f3cFG
gIqUQ9uu0uV173ayXT6MJB7sDDY9/wQ9k5WSop3KonlD9KrJbKf0d5k/q9zRfeda
AYb+YrhYODXx3I7sHjigjaj9Qqe9PzkU+2Auf+HNZhPFFuQTAJbS0noMIap41sRP
4sfu2aK2gozK57CdiZ54vZrcnDH59Jelq3REdB3Arfhd81Zo3r0BrMGwh7K6v/0D
18FfRcUbcBQaQUm2bdQL9GW34LVMl8cJpG7yEJzXFAS+TWzwd3f+sJ13wH3YBsy8
u2Hr8UtF1lAmZs6DYfYYka5NeeR/fNq++9vZyOvEqep61zb97KlTtQgy6a6SDSIC
EZgIkVN8+ecZmfRzGConNmTUI0nWPyo0RJ66YImAcx9FtHUtuF1rBWL0QaxdnbGc
nER1LB/IqGWeDICqAAN/g8cT0reVDwoOhrVUhBHKj+9vnOveAVBTCl/VE1MDEAXU
HYKeVCwsjEgdNI9n7XxN66t742Gs1FgSwz+zL9HnurLMbrKI4/bQJ8IWAPQOq/wZ
OYjbtxx+NPARjZBqyVUZy+wlaIjOq/a5YXaVZdspXHu18q+pfFIwNNalpqhldkqQ
Ya7qF03gMQ+4NQB7ccpIbPZlEoNwyrivGh9iY9NsyEXHvzF0KXW5CUu6DGW5RuRn
O1liYZp8bWvVGA3bUYbz+ODifjlOBDpQsB96YqcFqNt1F2YR0gy52OMVshxDP7hU
2G0e4G+Uu1ToalKsfi2+5sbVan16aVfU02o+X+RhT2/032HMHYHyYfJzj5eL2lt3
vE7sYg3J3KLTQ3DCSrrxRUE6PDAapyiMfFCRKDp4+DMx+Vr4ZinDKvYdONyJV3sw
GzTIZ2p47SHfUlNSB0pHfxy166Hz29GenR4SbdE3lLN0+VTrWW/QSQacH88oK5Ee
ULrQM0HjK9EjbEIuDQVb5jP3gf2bOWvZYxk5pEzluMNC9qXEy4c0BvEfr0WbT2CF
6iAUCsX9aciypz1oBM8l6DtS2UU74sWyckurKDOHyrAkhVaNZOMJB6tIUohQll55
liAyNLC7whPBxtUKkhOkG+5oSMu2oDnxqo9X8dLb6sqCbuQPlv2jkpRFm5C/GNfK
nDPH07MLeMBo3xj08x5oSffbJlzMJxd6uz/hmvBiHf4hdZ5sxXFt7b0OZmSdngKi
EurVaRSMErSzTZH5ux0CbOHDRGyIvXa7MdyZWFq7ZcxAVy8Gg5BplWd1cjQWjQb7
fpoxk4dOXw6/iEa0qYGBNL1J1C/CNd1Mg80naPMm5JOaXPIPJfWa9EEHSivPEZSk
m0EhpzyfdhqE58EVlSFnpo/JYzbYyHiAiX0KRpdyRgP9MetgwyCcSSOxGTzH2/gM
ei5I8Fd4xxuuxzcEBVHf8Yr7Ld+5M+Ee8LafRWfwlAVrUogA91LAbwAWoQOvClxR
4PMbHS0SqvDZ7KHuNOPQgKceN59wBGYVz1JA9l5y/JKYnrRRwvDzleSmn2WjjuwB
cotiANSDcSPZGULY40xvtlyGDDd7gC8CWs0JMzoPEW+lf3rzUicXMe9+p8p1iLMp
GLls0EfcNPFiG+9Kkr3aRvn6elk38hmiO366daZ+AlMsKIcCC219cAXOK1H+U6JT
oO4adbN5RdQn3lUUBGTzOzS1aZxnPmxJAgOkhYTB57MGfRSotHiaXjdRaZZca/9p
/S3Hn1uLKlKxVBwhGlrt4lByT+pOEXK4EK9e1UOpaJ5uFgP+1h4756Z6cMzlKR3Q
i81+fzNjX/kBjSvitE0AOZTIypOLUkRnL62adZdeyXCZ+6zwJb7tvhh4M0uKIOs9
tFIHdbq5eDtJy2Oc0/2XU2wKPd3j9QLWAGPpU13FZJ2g+mJgZM3uWjg7DEzJz0n5
NO8EK1XsGQ+VWswdzloG6Zc42PAfGJzsipaXboCL02ruHyeSbMPKpDGgwTvp6ea3
yg8SPZLRnFpisLutJqz9I3kvAgiggdIT9X/VnJywfxda7BGTVtGHXhhF14xpaEfc
AFm60BDivP1jejwvGb/bw7cEH5AugHWjrb365wrMjo3XElgSqqNLDOMQ4E2Es+rf
2Df4ZltJMNnwL5YYfUg+e6tV7uKyj/bkOAcNYwiVSB23DRmYLqnGlscgLKQj1MZa
AFxSrfjjJwUz8TW8IoplG45wnIHhJDHqSSNJEcRJ01nO4rJKJ5BHkRCUb9z5Z9q4
SWsjUxYGWg/sB4HoRGhtmI9phXiWyUVWIDrAFcjzTz2bUaxHXuWj4qutNvWp2xO8
UWNxyakKFnIOejUATJMwgPDyf1E8HSLBdCZjEXaOfVYPBM94cFGFmb4zg71FPECk
ZJgd3ti9VYyB3CVz9eEbLDoaQIn20bDMTOirFnr4Lps/ZMDWDWzW6KJoWLCk5tg+
k84OxU9EsuVaPLV5KYBgShS68mmcVidwfAcrJRX4lJ9DI71rAzYU35dwVBviRG6z
3IckfOmAnisAzzT3eKoKQ/9eedrx5fGIoND0OnG1+S8sHN1nf1yfW5KjsltdpeQd
PLnsHsyCMvYjrK3mJZfSxsg46srMCXOiEkJD7LKc3I/yXtqIuTIA2oTeNk9LsoJE
nH8CH8bcAJKqVzh1LEQCCTBHA+glnGm3G/VPIB/DKjbPPqw5plza+6jfgVW3DVbc
kGL2hM59YnTtTvQOM6S7yI3fPJtkEnRiPN15xKhyMJZzUksJHOJQJlhx3nnHTbF9
MMo4hFnaLyHERTZPNqGDT7Vk5NNRgmt9jhfBqoz1z29wTjqoJ17u2ATM3qgiYGod
7ZnYTYaknAVOe5SYiyfnWWiRgaE2nxVs36TMxn0hFgJUqHJ7H8n/9XB/wzezzsb/
vtPAecSwDiT0STaYUJDCAE2tVmNAgdC52abR6yp2Nwz3eH7S/q026rIJe426jV2K
/lQWHJlcdsRIMKbQOVBA2SX6nl3istb8qfvwJjPSiLfJjnhU+m8tch3cE/dVf0YS
zV6z0V5HMW179zOTkbAJOCHYEfzIBSt3AOUvkCFuEq8Wv2aCKbjgFSfGwRJo57JL
EFh8hU/KcR6ACZPRHem9TyYesRBXmb/64NEintyR0YC7waKMhX/DC00wX/TP7bR0
lBaLV8fzghjv16fux5G8CuEeuzB0Hy39L+19XeVozl90O/jYxIcjClTPFMth5dft
HiOo9NaRh9lhwmF1ik2MElvA/tH4VNBCrW/H3Kllgjj813RQqnDDOQmBsQvF44nE
s9suAAHXJ+NZ9EPzg/KSiN4LK6b1odKBj3P6FrNI9YDegkTgob8yZpr8hoHSpdBI
gslAmJGwnhZcoN3o194ObfcDzWLbwCo3YhxyRB7bdp2ujMc1QrN1zHRcOAs/dp09
NHJzQN1bgkmtnLWoL8svdByZrJ4wZnQY2WsBurzMGWMZsxDEctz/KiJi9ar+JPHr
YhqxEsfqEvn2wWRdhIEu0dEZeIeT5MhdIrNYnIjW3tzvNGWOyM5SHTexALSpmryi
57x2cJNE7ZfdqVKdaEoqS+XCZA6wiCcmdDIdKLidx7ctdK4RFAdG94h+zQnGpzkx
jNgXbouufm6pNeGDchyq7vHAvgX/2CH6V92dgZDM1qeksOzb75DxGcZsLP1NQMz1
LPguTOMIFIQ1NBkNKweJwHBVt8sOPKDtU0Y7UsaYhJ/XGjtmDDkakclcUALrlsW6
2tUL9FHWYnSB7vUxoTncQ2WeX0g7RltsH66jH6V1NbuYJAOEovaNAuRqajkMaDRM
rGd6VnWXFnsU3Vq2XUrFNxzc0eR8gQsbpX3FLVChhZ3OZI8hj7g675ZaKYVoGp9F
78N7tBENI+0mgtfQiwXypCynMfh/fCcgRv2ju5osfvBwrYtYfCRAPPHQk2FWmBVU
TbQBCaomFEvPBSlYeHOP1NGofHdZ24Sg6CX1zkHYTHSB0PFw8pFe7bmdH1L77Zy4
VBKc6KNXrDnsgYQ1ZlAOEMdvmbV6hz8vhLrsimYJjuCHKlyO1eeEZ9VUrLURHcvP
jYkF7YxiKHXaxZwQvfJLvzS19a0B1PwJfjNiN7W95o8nLV2ufqxeQZC24NOYAFjj
IR1+BCbSm1DAhJ+aZQJcFIAgao4II/Yk3ndpkUU6SsXRWXN5l6D+kuPheICOntiP
vpK2CTJQ4a0KtwLDXr5JuGVf0MSFLxC5fGi9sW75s4xRd1QcWyRcaASmTY82aiPi
qPxwha7qD4LFdNe/jJ/cH30h6UuJB+dQiiP2ZjdsePyI2iQ+cNwP7luV/eMcBxIs
8cv4dM0U+WfZUz2ZeuPdlCRM6YBRThCJuIrizWmy1FENn6KfvpWa/Pe2DZ5dh9yv
m7/sV2Bmc+RSfMu//CG1I5BoRrbCau6URYz05NocPntqRGrfxP8SwnHBQa6wOc7O
cvnmitQ5yl2MZOKNMnX6sECHsBTQtL+R4YIksrLrkH+901o9TkenNQphRVaplZ55
YyQ7E1VIQJb9x68bq7r/s1cnDg2REJ9aZlEyNdVAsJMkisiLl3z3rW/9oIrsckrp
S1diW1cE7PJGnEpJa2gBPeLS9FLP16AN4O1U4vNtGf4Y2Fua2WZk49I02lBM85pq
ubnjdK1596TgLumJgvu0qdr2YA1GDihT80rX8tzc2UwI5EWJe8CHpgbIbSFJ1P3H
KAUJoAaYOCJdk1n81DSYrbGnuvuG8WARzTCNNUEnWRx/+zu7btukmYH+5P5HsNLl
HS7U5h6EIzKiManKWo0JH+aNYtG5MRjTSKcvgO7hoUwm7M+dw2+LAhfcDHZ8ENjD
X08NXfb/RrozZKokR2AcDXbgPUIlXhiq1ibkHGqaupyWsJx8jHqHab9Edp4H2kx3
nvlvFZOYrYRRUVFzYhei7vwlaGW9xIffOaCZbnCtY5ROFt+Bauf3v6Tn2l2qz/L5
W8mAuqOQqUoO8i8x1e2U2aL0jjJwD9z/Hq3G0xwXdObE152FsJ9ahS0H6pHvaGV0
TEyvqpj6WVWxWTmRxHOAP9TAdgozmts08Nz5Ztr7LUXZupm6I8OteIPaiCynFxFd
yXRUvi2jNQNA8Z2q7d9rOZ5EqV+D3F/y85C4V/VeiVQaVizw1YRPpHtvVAYlDrUZ
/1A396yD0n2oCdOW5CE4x4ECHNmFcceBf5vquZqEDRGXH6OCxTN8N02I+d+suO1+
bHkXNzJwtgTReMma5ew3srpS12/qcmqIRcYxlir9jY/fH6GFgR816KDx2gUiG9jU
1HjnTitoZJlgnzaxY6/2mRmg0EbueSlkzMIEIVSN+wkxYsYndozSqCIdNQvuIeUs
ZL2FXhK+8c+xmlpn8zdv0d/MQQStAGJomaSgUEOlXtsNSOfELlaMxWGJnsbL95ly
dm8Bvu5Ts40Lc/cJlokdBE1UdzJlmKa7Gan9mBT51gwESyJyvtPAgeUBVdvlaDXQ
H24RHpwG9D2/U+vVR+eMkRDSgmu8HQJNwgk8BRA35/tRiQHx4dtQMLtvWPuVDqX1
MfSithG0QGF/r2eHuWCaIeS8H4dYuNY98d7ut8stF1r8FvyEeeKVFC3/u/C0kQ3p
ilTYTgx9Edq2js3pqnnVTk/FdApCZ5RjW9Hwf2HZGKLwMt29TeqqQBrlPLec/Mf+
4Ad5AFEcw+Gj2GPFklRJOR2DirGfFQFbwT06180Xm8ROg6rKqlgUR5eb3zcN21tU
GO1P3hWZns4Q7K+M5o7GUWkng04Y7FyrSRu67CsbxP7a77ie6RVHj4S9//Pr1Ax0
C555Pt4M3odyUe7Ren1UW2PpV+5wPuSD/lsjuAWL31EKeJ0915Mu1US1tRyaurds
i/JTXr1l0/BSSF88KWIeSWwQ1LYm9jNvfoxpV8ll8SRFycOBWtyjF9d2lhJIfYKb
13KKYKC7EQIVA+Hr8nPDPoThiFPKfg6eP6zh37HkdzRLnnyHfOtLRqb2Lji3Alvo
ppeu/dgl9KUM7PPbeRZ8AzP9D/knidpXZfVExy4p4Fw4aYkInN0xCjdkFqxAyoPM
zEpjY+6c1Yi8m5wyKaNUYUBxVY8zgyq/7qOMnzJ8uEuh19wHCcszKNXvdJgfaLfv
eDgsPzjaM7nCqwSzARZItDz4Ohn+1Q2kkR8fWdJetiSIIkdU6EvmELObKfXho/ze
4UceHzMnBvGZQ0TM8Z+qqi/OplekQF933PqSh5mROl6g1I3LENz24yz/876Mk7TN
BcEg63u3cT+HAv+cH32d0zSF9KS+sKxlllaQdjFyXWWj+Zy6P0TKNxNTWWRMwvUu
Cr+EJw4Un5t62a/TTsurCcb843lq27U5ebvL+QGhfdPQgdpGIgp/11xLfL1p0fac
OVpry/X2tClmcfO8KgJoaMmaNCBcDdVPP7blLFRzEdv96miNkKm9TRH66veOJHwE
jVKllrzcmdQaXhkKIj2F7ZKv9Wft7P58aezAqMSyzj+eX29gz/QSp8EVrjNBm8LW
z58aZT5vHPBtD9nA+3bqzjnx1EvaesmJUpOSgTk/cx2PmzCl1V0jYSMa4PFGNXVj
xbR8EeM+bYuedeKfylQLVvpZNmm7uAuH9664nTi+WafXWSZyayugvUX6S/8qVUpV
z1mAqR2qzdunefFwGrCnurhKxnV0WcPGcz1WdjrgA5gbqABCx/kJpr1En22oG8Qq
RIEx9QvdRfyEiW0qQFs1v8MJM97aJ1/HahSifXL0qoR82zQ6WTmYnfT1pcHYFoO9
OxMYUOZ1cls1EQJFBhRUzWP/wx0QylWCiOPuFCv+ZJ3VVPDnLxnMjP7yUZ0cT4sZ
APXno+dOdKpoRGPiea0f13p5JwdsO7s+7ud8sEZSx9JKQCpt9jsA5FczWLe5vtb1
7TcTSgLbKJWYLaSlGGHrR4lpP2yICY7wkFE3Q4LtQHPm7N393GPQt7APhdyiYWeV
l6W9TKhKsc2BN8oyNk/r9Aoa3kAHjTwFrT77/8SclRIK1I5hiO8gwsYdvVWz0uEQ
tYUNTvjIKsxnNE2MaHYf9uKIYFnniC17ecRituiGds6io3gpLdLYrFvbQfn65SYJ
BKlCsVQd1cWJEa+jQ1r6PlhXGSfjGPHDwz535w6kHYAWs/+rnefKTZqTgbp53p3J
UeJF3hRIwytgrRgFydvR+22u5ycc3WaSLVkGPkuJIAOrPF0BMHCzzXK9A+zRHv1S
VN1jwDgm5YtXMtbtzq6QPxMaoHMVbV3bf17LQ+EPXdiaMP/XZ/JzkcqNe1n78aFH
8UI5y/T5zf5HX3YJg6dLC1t3rgzKLOMpA0gCv7+FgoPRx9veJSlsIqmuQDnfNihS
dGe6Y87GwnfjMZoR85d5K8SCRBYqLlxF/h4GWPg66pJIqVVa60xQCkvoF+hfKzAq
EW7S+u5dNzVah+FE5FxunMBDVP8rnrKj77r0nY5xzh3G2Vm5L7wUhD1R7hxr+CFJ
TPQBJFBeHpSi64KBpO+p1bfosGDHp3wpSt3pEz3/Gok+om9HNoPHrEAKntUvLtNI
7NrJjr4wqpW2kalRyeCs67oEXwjXWW0fR7HeFGPDUDJQjNuFJwX8pBET4RcNAaPf
j7HGayeMd3VkA6yXbppyRlQHAZifrrMDafpIgjnovvsEE9hGfFlim5sKmeALt0JT
Ae6JQCwZhdIUECq+qt6dS1AjUzWfPcHWydtUtCq8IeTXZtTk1DVQ+I1FnDgjqZft
AYBvpd/iYJXHuvRH0bI0vPMfm0EX+Ow4MZzjMrKsGU2VREybDKyz7fNPurM/lt0I
j2My45armOqoc2JdydCiFeT1JWfXQiXquE7Uhm7YnCsv6Lm/egw/cN4eJ7liP98T
6cZhCBvI990Tx2Tv3TST5dWEYV0aVeZruGPYV/8T1sCMSZdaHKLWgDBeJYxdkbrX
tKje8vNOVwIFG0/seEOW9+fDaet/GhZez82N6HuWv1waNaa873U0cTE7HCynAYIV
yB1++fkTPPTPUtWKHZtdX6RxcxggRfeAsieIiIsAlEsuJFMRHyE0k76iKO2zOTqR
UEZkT7lBpEJhIrgFVM5XtDxhyql3ytg6STR+hTCyyCaWSf5uaAfJ4ED0GgPFsZS5
F4+/+H7XH6MCgE0RQ0j4i83govnVeyoOmngBWV8SuNmPibfHoUmtT5ywyzEHhb0w
zH8o8aWtFydhzra0Ndk192TnUXYh/bzgfAjE+H7+cMBZWFgOUUyGCV40hUz78qET
oq7nVdh9tB8ZXCum5xXz/RNKHLRNC1SwUfPuVXEBUQsnV4/MvCVlGSf6cLNoi9gs
ry63ElfIzxUarN1OwR7rgseeJcmfDNoWR1E6GwSchx7DshnqVIaWJrRweYt+HTwB
sMZihhViAD2lTtoavOg+3AHCfKvVR7P71SPv+qG8KpATeHyM1zMEUwDZXYpieIzn
qiJdCE+Vo4jvPIDG+fg2+I6ul7wphb0A0gB1he3jQTQZidvXPu7hCsVDiGyKBNm2
QUKQ3448zRBbumx/HAjpMis2cWv/J7V4HFYyXQkeKkV+K7nlaDs/ysCTsDO7xwA5
VD3InUONtIu7jdA+42CRD0yUFdECdBvQUx8Z4fZmj4MHPLJTpx6aXrJYRl6ArYFB
fLR4cn2Rsn6KyM6cnR711qk2Ztbvy/4jDw0TPyieVBgqHdew/RPnxaLKyTXxSEty
BUe+3ug2oK2JPL/CwWEILCeLTBn61zYwUptssdZBu0FHVfNJZLQYcd+Q01Wr0ckC
WazsRZPrFYDJDfyElbSM4bA9qBy9/oKAlTJCT0+2cUvGiwAirAirG/WgwJ901hfs
u5my5gviW1FKq4BOODiWTqj2Hakx3H05mppcdqag4Lcf5r6qmPNuWavAM3OlzK+E
ndVv/J8qC7kTwACisC5sEMe6uWOsNM+qYkYYz2H8UxaWlR7cinhkL1sbtq8ArkQw
U+bs+OJW8mARByRwmS8ls5LPNMt24xI9Nn8uwXBiplIAqQxr2f/EfKL8APQFgWYp
8g4tFzbm3zpN4DV1Q1qePARiOYcxMP5Su9m8R4J71u7bbXU7wezkSVwJQWv+Uf24
YV8GCnExz1migCBUN5O5EEaEYv0X9IraWGxYrmMO7lzXeTz2SXgIKPc301WfFnLp
DFHJemyd10TscWF73kGjPc95VjaNoyBUXbR3hC7LZdSXyrzRJwO92aI3V+YsYIWE
0BSBWD8FxXTGKa8m7gBS2SWOnut9iavzv6fvwfljeZI3CIk4cbx2RLz2mr+uR/S7
sGM/gDsh5cP36M1bdCZcLMqL2hIGVJtK6pxt1rxFVQ045qGRsRXRiI/8ovYhsfvw
WhaErGFpbDkCAo0gfsLWLallRJxnUQX1dgl2QJyF2+e10HsxV7/x0dGAvwJy/uJM
hZ2I0sYU9XFW5S3MYQPuNbxinmYfRlrcmYv/Qs+OmHvv0bqoeOFJY94y3fottO5N
TbHeVQlUYTUFbGIgq1ppP6DYD0HE1yPp44mMTdPuAJsWGSRwqgdhOo9+I57hg8Es
TaANY3mEBAMT9mBSbsXIdd+rOi1g6Jt0tfWJ/GnT19wtrYe5p0VpYL2ZRuJ8wMQa
dhKuSHpVFHRUy1ThH+RZzqcUFWYBs/8oHgmMzLwOhZBJlZ1v4BXMYCYVXKhof/h7
PubGC9JLS7c75Xj6407regGKkrpMeLdJuYFlRZIhWRVuD9+fynoDDXFtF430DQJ2
v1/L8moo5/PDGp37N5vPT02EhAuBlLBeoesfq35Kjki2nEMAloB9syJ3EWaT1YQS
eBBTGlwRK5bBwV38yf0deZQrVYtq/VWCcP+tVGRaQQawa8uBYD38JW/x4rAJPwiB
5ZZaxgkZbGWRdySA1Dq5C9fH5NpOeGLt5kHvIXqaFNNLTmZq8soorYjxGkz3s+Jh
AnPriKv58G1DR+iTRt0axrRiExj5sfPc2XZfUuOW362CLPeKmEHNMPQsrmNVeuKs
qUJFRtTUcMfNsK6GX6YNFzSNagIzGPRxqGrApK5OM51lyzKuZlLndy6yIo4xjPGt
sc3v3yoINl8su2PXDgImNbd9UVcJFgnjTUakOsQ+wAykshmXIBKIliyKJTQ/YSVg
4SMqlAw4zPKOsnxja5Vf14KZjWkgHKS6VseS7HQde8otC+9FzoU2dwa0KsKwnm9e
7bOZz3KE7DpSYMOJNLC1OaCBiz2qyg/vC1ckALX7SiAhI0zeUzq6Afo/97SAfV0z
L+LiIRHFChSSwrIOoDYd040AbWnhs6hXuj9iyKDOjxPdaMU80mMIx+PhM0KhR0Nq
QfWn0V/iDJFYoy83e29+R+UxtvrKEZLxI4Ax1eOoSEOwb82YeWRNYaR5eIUT9nz6
+o/R4Vf+tmHqJA8BdYPZaYvSc2s1jCpwu5TRJB/U/zTX6q23Ow2bZRYWAe+5wyQD
ZnFC6kdtBXUUAqIrYXfkLRINBwu2uLdCrmZioFV/fxhBb5FdP3/vXz3FpMbinqNE
1chNUPLLK145hcHXBK4TMuVBULvXbd7zFP9Eee5F9agnbp30IaKtfeffT6xVc4nQ
ALGZxF5VWvBEqzpyemBcj8aQSH+pNBTkUvc9vz95YiiBGev0gnXGYiF3M8WWZMOb
MctBtcHiMIYjXk+GTnCBRrqvT19w9jlE+q+bGnIw1AtJcgGWhHdp98H9yq0IovV2
l9KWGI+8umVokUxtdMimYA83C+kWDPTpar/JqTuVqBi4Mbibhgr1Lh3HicF5oZil
3eAzpAygp+pL0t2QCODiG0w7WWh4KPVaJneZPALyca0qSiAjz5+o+lJf2BdaapCU
iRshtkCgT2jgVZj18ffddlYhfEeNJfz1Iv0IEGFjdfIkOaZExeqDLgKgRsdwjoMW
0ZCz06+3kOhzItv+XTfNeeuPZoiN7NbVXOvR7rQY5z3ZTFwR1+VhccPmD1JWhQMc
DH8gSl107KqISjZ1p6nFMUL2DVlX5rYx1DN/A0hf1s62y8ECRU/hAxzMic1qbvsC
FdpiaeuSAtImFL6Rp/hOSawIvBMXDTExZUvobigNevbUSqc2C0I9W/RmGYyHZYEg
2/IGgnQCBS4qPe8FFxZ+Gl1b0T+0AZCJne2FGsT+JJn3MkfZ+VWcREoKgbdJZYV5
iuGFLrDCX1MSpsUY8RlB77WeZbrkaR+AcUmWcv1HHlFr1mQ4ZGAoCsDiCSoY2ETr
qlCuLLL5HmGAHJx6CRNNMq5uRN6q2378euueb5kRyqpfiWtZX2ophzrrtooI16lL
tnkOnJCK1vJQIoPkOUWqMRnnWhl2lVW6zRqO/uY2QLbRj/5LO4WoCYCGj9PM4CNw
hzpVAzFj/gEkbk0lsllQT2J6MQgJjR4/znXibbHgqATFmvwmEj3ENMo81cEU8O5i
FaQ+6ZQ2zLjvkyGJa9KUar1a/jWSQD61DD+3PYf8uLchY4xaOsYFmQVCpYOxz6tI
J1VWto5vPaNb0Md2of2AKEKVGC1bf/eWscEH4mmnyiBiMFmqwVyyEaXY5V+TnQWA
WHK3riD60iG6KqZcpmugnINDFZuuuhPmpBgXwIxQ3aWesntTBDarsperul4koBDO
TpFNjUMUfX3XuqaI/y0LrL3OqoBRbHw36oRvmen7gYI5YOdEWdIVD/p14b9MeH1z
JvlrmAm6be6AJc1IV6Yv+Quwcq0iSLH/POUIp+9TSVIk+k1WVaxj3ClvjHeSKC4v
FKcFhVDvz6RBk5F7VlodX2Uy8+VLA4xu9tglyvNa13tnAtWXLoo1T3vairvBb3XQ
aC/ia5cruwNcTfW2lbYsAO4jgQQVftwjxDdmLKwo5p/LeWBx7Mcj1Vei6HRd5aRi
IZAN6LmjfyK65KdFW9lDI/FU6NAl+TOJd/DbrALxXts5yYSeh0Gzz/bjadbbOzA0
Na/7A6GBG4zBVuoPdXjqjdHSKgXdVkAvf+h7n4u15wA/IC/TRrEgkLwJBOgxgevZ
5Evuae4x6aT9Gag3bjh51Z9a3Dc9h2ILGqtiNln3xSCKl4KXJfL1CNdQe8a0SHds
SRAAEuoNPqzCe4xIV/kaB5Skw6FA8BpKRSsL1j6BPD6VLIeSlz9bwgQYNHGDHnpf
JptjUBuST6l9ecbggqAuYuCRMuD/2TXcxA56VeBYbKeJ4HDO96bbRQ/nMGn7n4BV
rfwo3O8ta8Y+u1uoYRY0zkFntJ9iVSSgcYIWhQsxlAK5tEkKfLYQdGkDp/ekP3BM
7kdLV+Xc2rmkQTFMXlqUbuZS+8XatOjKqfIXfQTMl+lgkpnL/vu78QcwFWZ7eJ7E
w+tIVAjwLebBEQjrCJLlAOETxUvREhSIKNd3cqUO95mPcyPIKbLABvuof9RDjP61
dyV+Fpxi0lmlUxIpSrXjDcZntUGwHXTqiwXAV0E/6ZVlmH2DGO4j88gUQ775kJD3
hvYRiJbcuy1ILZFVdGEqOu59DRMZ7FJMfY64QZxS1RGHaUsQ7lG7/aEkujuXu7pJ
E5Tt+BkrN2Ow+n1WHCOYGPNg2IWD9IsIfnUubcVXHmiARjBa/l0GwMGztbdKFICi
jiMGsOa16TJpwioQq6O+MiZKtnsFCQwLPTa2WGh2UIwq6xqTtUBxEGTuENvhI1W/
4ohqP2VZOT8issQDa6APHy4GvvKE8UKVOs4xmvIgRZlxM/kDOT+tA0i/Gv5YRw7n
w0GQvsmeosCud71CiRnT3ZZtdOHBqVfkdD5766MoZQbZUsj/r6qirlhyXMCsavQ0
Svi+QYnlmZIiTPNA2CCmmXIacwkCAcri2jBlwJmT5cG39vINujBI8L14usd1aOpc
bbg3mNyD5N8mZh3havitjltawbcGgHGJ2DMhK9ugNYWCmj+0nRcRG1FCFZibBXoM
zPiXcqfoEKlYrC0WsEhg6ZOAfxH4SB2riap1gWr9P1IxvLTXZqGeMiFpwRCJUC+w
R3V9lI3wsaXjp595kmiNurHfEfhH55NvOOtxk69qQfI18nliLlwRIwBtP49+btEZ
AWi1dxPNaHoyWHVIJYm4QVogmZgKDsboXBmdywTYQakm+nhUrdavzqMy5m1C3zVy
OwQZVi22ayR3jzck6GfBQMG5Ef8h/TiQafC/b//kmPszzY/N4TwC+6/frqI3fTMk
1l6Nn/AaGunXZfT9N//HraPYXt0g3IfaL0UXZ5rWUExB43pDTTaoZITnjhOXJcqp
ATqQfol7qP4dcY3vGZgXDylMpEiLqvJd/alQMXAHfTh3ltmzqJbmEaxkVMvMw/fo
NJu/MTnTIqteAw76d4pkV7pUkgtkgqUb3aTqnPL3/zcJT3lBnTpsJxg9HySEqz89
UQE36Ecl4zkO6YMko50G61nCF35xxuiOnA3JosUlWMv3X8/6mkXLXzi5CvWvmrJn
wL6yTEiti2+f/QrqKKVeByfO2UB/r7z66mwXVsv7PdPjSgOzTq1f/8lOxhBG659q
ILgTVQyply0zaha30w+BToX5loJBHQFlfh5pUmtTBTzjloHL7oPB3bU0Z4s1Bxjy
FDmXMTdsEqXDw6xqG9G/zMFnUCwSXAyhfka76cpHkKuqgpFoeBhOHGJciQJAMfD1
EqZp/isAbwnRwPSRAM+PolIAmcMIAqo/z44jKNy5EjZMly5Gdf/9s6BLxyVlyK27
xLMT8CFeymcKqm68XpCegROxbvMjNFqu7nUSMryLsiDy94Ks93XEevB/owIrVbVH
vsGjsrYUmXII/++SnwfIs+tHkpLUYgR25b1FCEnNu2/js3hdP28TKAsc/xUq9XYC
WIgPhXP6w5Q7ESQles4/7j2+wWjiK3L7xl8svAsllMWXyl/wPMwa1IvbwXh+8YP/
KSwZZOPd5W5yB5c9R1+rt39/LxaJoy+se66ZoZ406neEcCaNnYc7bbpnYSU5v8p+
dKpGDDvCO0eovgSXfoWj5zcVykxq7rVmqACXxgk4Rzpp/9I9P0Lpt2M1fvUDrxtr
MIi2Ji+dSeo5tQf4lcHGeI3VS/UpEwvr3U5O5GsMtCgwt9aHDsTdxInCjEGCkoaM
v46j5tK0QrWmaZVOQBmn0BGfNBt9s9Z465aiJfMfQDBTcDgEt14JghSqcN3FqyQw
CddFFgHi6lPdumRisYdRV775UTp+ymFh1ficVdLSKBj1tA3HIkPo1eeLEgXUJScr
5nDQFYO9OVYFh/l2+Fd8NytrAlMuxUQK/XO9dHXq8y6WsI2hUnusJ5JwFBKTGB+q
DWigW+c/7EMFXLklbxm4cbYZZEMP6D4N0ae9ca1slkl2k8ebdtH2k0BUUNGLj1mL
58Lr0tON2pm/njcgmPtRpJGb8RrRvyhcrsueH36z57AhdbMptz2oCDo7uigp2rVC
cp87bFrAykD7Qf/rU11wErQYDVbvOhmk1Y0h7NWTnuXOYh33TNA2RhKRnN09QZIN
aGQHMz6/pnfNHoL5NXwsdyRu5qwIwQ+hEcyeWWE8LdpPvD6PytH+t2828x6jrVkL
7j4qUrmyZGhQNN3wKcSSi3SLrFD5qYeT7pujRD9E6OAc+MBEQ2Y3gVe0F4bhrowx
uMbTWRoDeQm8j1bKrSruBvO2DCOXYYz6p7rvTDvW53t/2oJE/P0A/JjDGqPpWgbx
vxksT8/KWa4uS535dOFYLi6tumLn4MC5nOkxzOIyeeyhKMQ8MhH+OS3HziVDDuLY
Z0yF+gBr+xYH8vL6WHBUOcO0xaxbOZShJpfVjDevPSx6dipFydI82Bk5mLYxdF1U
d+JjUCbSR1HFPuBvYYbntokeb8Tn8L6AXCXOPJksEXeUvMKhRZTLIzvopp1KaeLo
wyzKeQP4mC28BFCMWN4ZYg0YpSFt5nU5QCMbW/N93lVwjhKagnlFZL41HEFr9PmV
vYLnbGThwc3bl1s5M06C/j47MGjBQJ3yMJzVmjDr59HgiEVL1sfsPURzumSJhTm6
GfKufLKLz8bNIrhaajXSwmyVYy6AuVCduevyIocI5fuF47M170KvHvLFBJjiz5xT
9GNOeUjWYdB32wZhIYcBTyIieCy2X3KSIIQzJyUfSPK7sfgESbTLcvqKHZIbsbbB
fAIOSZ3Mdm23EXbeyaamh3rhSora3P8OJTSswSMHLFGwcmqlKPh00TYoiZafYjTX
KuVdsE+k8EaXVftcKnk8i5E7qEMi7JzXcidRnMnDYcat0eU6a+12kkVMcJvyqxUF
wQLtMB23zT0oSpMieGG9mxNh68/uLmVi2NEsW2dZl1r1WWuy0V2zcBDtYyRVQlDN
fWQSZyn3kqYwn5epHDKjpXxyou/5ZUmOMMwwSjJBciAJWqLHCJVBmPTJBuskKKaw
L5xmV9DmsuX18wx6Urnq+dRX14h66dhnESEMN3m7dDQY5iGPdAfB0djGGKxsZwAQ
z1auUrLKvc8o3vMkPPbvo2XDKUuJfLA3LphDkh3cJYPcXgyQiKlzWXK0qNeJhiXn
upJV3yMO5UFT6V52Gw4TSal/PitvQXBr29/zqcMEutwejBbn4lR4AjfdNZ5ivkkS
E+rMYgdL9SFLo+0sBzEAg+MMofhuVUL9Br0AgqIG9gaIRMlJ7a0TJaIxudNzQW8Z
k5asS7pdD2MMOuaWtsUGamQIZ6s0FHyS2nkLhQPqcJ8iErRb3Rzku5GfvwOD02Zz
tuM2rAH2/68XkzQVNWXntBAAEeyViwkzyaho6sQYbX3AnbchKhPWVnj68onVTnhu
t4bloPijQoHQ+TuHTieCl0BsYLNvgnrsvn2J51gTJQquj8f55CY21X2pqzvFNqfh
sXSbLqkP3fbyniiodIDQTT2HIuup9CeNT6ir+b/n2dL3KOZSLOeHSVXhl0Btubi5
ODIXtVe2H1chTyXimaK7iYzTNBF24NNdBvyoakTLwzZWKswbmV/CZ3I1gpyi1Kxz
24PdEr+7NI5cQUBnWWtYebSf9CckvLejZsFWRRSqV2pKwO67t2YgQF+au/tnIkB1
c2aWJD/xiBhO3a0CVXqmdi6WVy+6A6N3dcvw+Tmb8ODihlSdChfiARul1e14ziYC
XF4Uok0w0ttNVtJcb/z6NHLWT3vjvutuDvo/ee4rv+CLXrzQs1y6Ny1Ui2Lzzq0y
bmup51cHtuduNpQITJS+ktfpe3hk+FoMZKzgoBRup3jRnKEZeo8l0pYApF68i1OV
ZVTu0oGBLuxijwWbE70kKGNqueZJL9fh74NnW41k7AEfqXTMugQr7Z2qeqfUnLW4
AewA0iLXht6H+H9Y4gVYx3LUlw5xKRQmYBKBLywUFr/W6PseeePShtfpikysZRwc
PHujeLk0VrCyxkEoZoDIrBXy3f/YOiCCiIxrYsTljG+rUf0JhfJujRobib2tfROE
/IXkSa460a6PaxONtUjnBnvAAgxptd37hFKBF0MCr+UvyW8J0XDeWLBw50Hp7Yvg
hJPGRR0Cx/9hLNVM7kS1dnHjP8qamMHQs44AmdrCb2E/J5kzLhJHaUeJfyudjvIw
eSLqlUS5jzbisERCzVd13+dNLAc2eWykbYNzspHlHQ9+xMT35NbMWMyDi2tBpkBT
OIotpvn0yEkEBmN9m0jpkuNaUcbS3JqZK+fbyScJK8fbd1aTyDPiJD7O2EoqoyeE
XeZg3iTobVELVxNSonbUpYuVYZJyxVPE6lIo3ywO9yPhaQugpWGc5TY38GiVqvVt
8ShFcKUN1Zps8cNmMwDEumObxGCJAfoslz7rPY/bnDd7vbfzi76UaHbaM02a2qq4
JalC+0WjL6gq6oiyZSESCN9rMkWlQf8nSE67WjDRtzap5rp1QxXjkJqTMqYu2pgV
GAq6c6InMNzjttlHu9ABpumW7SdcpiFMO9QO5XUB3TO1fFBtU2GiN24rpISOxTr7
5tQ7DBjq7NBR3AZ2hvnFhAV+7zQZOafKE1ZnxWj1L1repkCsqxAK4WM0X5LW5rlI
QaRG0znGZLR0HzX36iM7JmFpsKE5BjzvNMuKHeBnTTmOKaB7sRNlLyyq33NNPG4p
0r69cBsmzQQSM51tYK2TW+OgF0G8+fhw5M2xTgp1u9ZVNQwnWePPZTgJ1V/cY98r
tkqQ8ZjTz6j7WY+ev3O/HVwUgCuO7pLZ/pIwGsEi9uGEEHhKSBtOTOVSIb60rf7f
CvUIo55ypdZ0M+OzZQFE+Lm93e2MdaV9O8ym+O/dDEcL4r8rUcQLHwDg7bhiBbuY
gwmEFuZ8v5eWLMvGSRDRWkqKD7T9TWgWk11eKFTEOePunB8xiwbm0IfQQYFJVsf2
6zSmiU+TommFbQmv6JMEJqzh4oS63FGwV9RNtkSFL+80vrJVNxrZEvjlFx3xjDIC
ciylg59XZJw5uSUHBeQGKmmZuTZ/f5CCloAPp3VcAoKvfufjaGlDeStdP45mXjtT
rLTvOYDjjRipULEmVq31G2q7UnaAC7ZQLxqH+NWAaNaClME/WkfiYe0RXRvgvyZG
GFiHMZqmUXTZvf3CUVUuPPEAhAxo8i/IM0Yq5fkp4i6OT1BSEoU8czyl4vao4iv1
xd/gYzbcBGtar518hqjxcPH601GFX4+bhgk/iX4apyno/bWHqpSrNZMgSHiu7uUC
Wtq+d51Z6S7v+PrPBr3gXicJH4dqaYCu43HMijpDSG+Kh60hjTE/6d+TrxoCC49p
nkNHCxUdPFuyPhLwvo59RoFg2Z0aNvgPpgzNgSzTaduDOZsf9DG+qj3p2YKhoUtv
cIhlw+iCbuexZ9blqSm/7yrH1jbERrrD8/nnaba1ub2WWHGIR3V3T7+PtCKziInN
Tml/rgmD245MRYjCYO4Ufj3e9h+LC/Cj62svAZPxuGnb7cPyWix6pwyGZHOQppE8
k7YpZBY0rXbmD2Kkk6Dpuy/dPfwdntIXAq7jLoF8+OO0j+NSpmviB8L11g7pI8cC
bMnzu/PlUf6rr4hHfTOJ6eizaGT0d+i5COQDX01XmdMt28UcoYgJUvTAbwP99xTe
hnniCWymhhR1bHu60V3qAjlIO9zL8NvqMye5WNOrrXM6WETTlFp3KvqK6a0HemjZ
FNEl90SCQcFQ8b5bf+rOAOjICSmFvCV5kAXBUuAlW3ch0Yalheb+MX8bEcAZvwx5
V0vSqdxT3Xe4oCFZ9iCoyZSv5/hFpAQZUq+WQH0T3wj0hFaoOSKLECKXKfa1grif
1OQFMTbDeIoXfaE0E+5M8wY46OoEnS/hBqYPl/i0lOvUWOoPm5fuj4WcVV5BcT7L
0PQ6jfDdZP/JQRL9kmIkcabVC1mWnTxpIQpAVUdDu7/1Pw3XI9fb2E7/SCenvUj5
qLQcu8z3CiE56xsGHTEQDzjdjj2o0wSJjDejBrUzQA+ZZA+/doDBT/kO4WBGjOpL
0Fn42PuW1DUhb/eWrhVYe9SfQ5gNG9WmmPZpGrJd/60G5aOnWIBgX3LCZEOCNXad
ANw6GNuaFp8lBaIHeACoVP9ZDYq+bzylQixOLuKU8vd8CGTTIeNrNSOWKXZvtHJZ
lj6vHntglSItBMw8va3UA6Kr9wD6oJh5I1jttt36Nj6G9BpSj9g+zbFIlpVU6ghj
zTVHQel84jFdvQhaXBsOytDIoRlymKxKIZInW+bfccpKATBRIAY1FTr88QJfBiIK
mWqBaQ+R43Q6ntxa/xy4VLeg7dXJDrPbdpyqIC+lo5wyo9/TQitYZA/mXdZmXCaN
ZBYsPwIVfcPNlFHiSlCUpkKDE0S0jfIkvJ9nPKKOM1tjbOhuPHuo6gydD96mSC70
mkgOVNbdMXGQrSduWT4Ft60JRR4TIA42csBmZJk+6fyttokbqV3nLj9lIrnhYM7d
V8cfWIAB6dctBOm5OzZ+gWFwMRPxtIq0BqunY8Z9jFOAKUO4Uz0JsLd4xEmwiIrS
lw4/xB4pd9lrxkRR4aq4UgtR18/1y65aAaY8ad0iHQsmn/6xCJA64CeujrCIIf4q
MU8XUUKpJllZDfsjTIEqc+l4XWTirx/n+0bY3iF0fOVe0b3Fj8VfteLuPPNsqati
hnuwH90Me5iYoaCQdiL0E2BT51VMvwxPvqD5JK7S6vaAd1OcFtWpK6nLWZGpJ8hV
JnYioD72SmyNVbApeVwXeYnj1VhlARzG9QL8d0o0tcqePwzAYepwPi9J2MpXSEcz
86PAW2oHoBgT7NsYWgUy/EM68i5udAh9ZQu+cQoQT7Rm6U7QVQYN41f7ailam6pl
FiIOcQb6J+x/Jo6+vIbHxxkLeumNDToiaUHbzMYMjSLEN82Cx3uvCRy+HtlBKyjV
Zxj8aNOgxe23m29mVszVGMhI2E7wDOYigx4XyMQAJvq2j4cGW2xoOq+nJfW0NM07
ql0I2Q1sKjSxSxJBjC2vxGMjx72LrXjEZgnmQdlfcnJxedoSrhWRQ8L6oHCtffSK
J90vM8RkdJpflmyswZtBkIgISpVMtuOJ0foebiCnBdGsVo+GtbWEcwu5b65brohA
ZVQgtHr5oa5S5jaRAdoTu/s2FSFrghUkThXZFw5XUf/mP0IoNSrUhsGJOzblJsgc
o/Tc/86hVmiwLAEBvddgnDDqOJ5WUfJ0Ejq2TSXxFzXAIQPKYyXuL2sLFzhZEzdF
RXtDrrIY6XXJHLhbaRsgIOqUHmLN2C7umZJjMLpbi4h1u9YtcYZvQ5G1pP1yogbx
Aw06YNjxGK0vBChGh7UU8zexhlrBdFExobvURQecn97O8m9FYBOpy45KmvQKp9Jl
Own5W3wcb6XUGmhCgHE+UFISLYCBQHRmdbVbUgnWEKHwAHcy6IxCWPglJfd03TLY
YU1ugh0YqWqHaYgSsIiOA31iq1ibxAbPXeWJaTQT3/FoeLxKli0RUJek20Wp3JSz
rW/sbxbCF/sIj7z9c66lX05pwncJWXSw+RzmJNSSYnEFcq8gSrkMEJQRGRLpJiqe
Y+IFKEIncTb7cG/G8BunVtPH/twK8dbFOKR1plqAkVSv0wUIUUMeReidoPdXX+m7
eeVlAnOy787aSIRM1+Fhhz9eAf+bG9LC1TYrZRr4imMPDs4cbStqy9Shjmt8TOKk
kWin5ALtvua7VhOV1A1dVtKRLnUzGpu2PQBUWCRWX/zqQKdathkwR/MkV40L4/HS
V9AbIcnTF0DR6F2KqlvSprHiAahlOLmqkV4E5T2302V5q6Lok2a2jTECfodYTvQi
cl20A9uMK9LxtY14LiMaxd3gbTv/l3/ue2Jiiof1VbkF3meqLqDc2kIy4WswA8t/
bfg7th6ogWjwbVm88HJOlrDBgz/lj9evCv/KlT7oC+oK0oWbmfDR6Gh63Z7NROor
uM5XhGLAD4KV/cdD1a1WgAGNzAUFKWKJy9uETG+krJFJTi7NVDz+2hsWNw0dF7QM
ZK8lYBFOLrYGiGWogBV9NrMDcvSgzaxyEaR15UAwKP/jT3quARHJ9+2xwA2lin4w
84cy14R8YTcvlG94WUEBOM+onBWq/VYVcK66xu1quNw3mFd0tNI2xAn7DiDMLitx
pR33AhWrOgJFmjDrEJL/fcFawnBZq3PvHfhjAZdk/ib5fHVmFjCe5hhQ/Nr9LZb5
3VWW77Bzkw+zUt2C3nSZRZydVhOa6W18rWWFgHPp6DE2+6UhfxOwzFeP9HIyPcTj
moskr35hvjoK+lwUk8CLTWUa/wgrfBZ+a+vnXLeJGsmcDYYPP+/tVOY+fFPf5IJI
1Vp0MWV3ore/BmRPhSKGRnGIA1/z0S7gHF9vK8ENLS30oXbT7Vt0vlaxN0TLpeqS
ulGYO7MXWrCC65fy0aE/zyWzSolC7P9aRanaPCn3YPvQqdfmX+614MRlkTpCpM5a
CiuULsdxeG4dHc8VTvQqMfmP6B3NQl7KR8aq+2SMl+NmbiWUDAxajNQY9e0jqHWW
9V3vx0IMyZLWuTOV6PeuKBPFhRComIO71QVtp6IOxfGpj+eJF0+TcuqamzFGmdoY
Uq9AUdSNwC4mxrRbOCanfGJPnjGwpn/7S9nZb4zcjZxYXqxDb54Iy77hLOscOJN4
Ko83UBJpAjbKNVAOkZmJzaZpWfiXmwPG1Hu16f9njuI5HS/UDDSDg2aM2Bji8dWK
vpu9vDJLghRgPMDBMza17Ld8E3XZzbB66Acgxs2gde3xIYaEifNYtu/ykX6KtEEZ
R/k5C6qNvwRw0DosDp1yz4nMgRlxN8rjXyZFQC40k4nJ0mBaynYFTQY3MLCvB9kx
d0HHVTE4gfW+q4rkI5z4U1ds1909XMwXvFz595k5+NjU5PRYMLu4gzRF5HF67+DY
qrAp+PsP1m8Ic7mrT43XRqvQHoSufnm59jxxNlepE60GZ3Kxw5ERJx677eDZkIrr
u4j+Uz48YxKUCk5OyjpQGSU+GpywGNMNW3zDBmrRx8DRTuLPny7Ft3Nlwk1+o2YV
ppU5xYENO2OAQoVuFbFZkMJnps3NrWe6o9/XQ6/hkjR+N8MYqH7s36vdO2PHe53F
05D1wcc1BbupaZkGINcfd5YfCcH/GU6el3y2FK06xh1nvwp790LDkckP7eaBYtqc
exL+t/VsO+d3W83yGfiPa1Glzhi/nzHN3sSoRxKOxaYbLwYR1I4fec1agp5DtgbX
8pp1jEZlU+xMFyRiOlGAR5lMMQCbd0pGYZHC655B7I95c8jm778Dnqu67Co1JXGY
/2FdZ56bUGdWDnVDhdlhweh60+iOuz9z4wlAK8+PDa2HMnXxaFsUIVVk+rh4rXKU
RLaLoOz4QciJ25GWQtsEP2kXuG4gXmewWLflARIdqH9i2PcuaBpGD6UmDq2QZcFG
5yJG4z/aHkTRkg3ldjJgn4l3JTfJEg+QJ/pOsL2prkgm89tqae3DTyJgeADGTpAj
+OMNgd6xUmmqdLrU36WkNsExD/R0XLCgRFsG59pw34pluTSHhedp5PNECeDP6roj
2wQY6j4Zzm71hOEljwiBMoCHxrKQvvmIm/+3hzuF/xrJ3bxL2r3rEposMov4sDfV
6Jw+czeQR+rz+u0bUabWXMoap5KEEbOS2aENClRbn3b7yZxgR9MwUGLQtr91oDYd
FRfjDYA3G6lvz7m0xyzObHzQjTWh6/VnVjvMfH7R7nJp0Wk8p6wvmtfnt+KkngFu
fAeeaVW5WLzWHQHMdQy/c2KMd2vcwd6+gxVJ3fHPrieoRV/rE2kl48tiUN7D3vbi
n+OyWiKLsjzcR/aVpxs+RSOCrXk8/WD81h7WfPT0ppA2S1/4OW20LTMWenVh7MV3
kbe5urEUg2pDMXEHyCKOK7KcOwqNb/w8KIkb0nx/17aQb4uMK+r2dXz8DCaG7yWf
D5ZCgfvshzZ81Wx8s36Qs1DSWGCs3NMKg7lytHbg1JRLCMxZaQJScFMRSVbwd5Qx
rrYj1uLVec4+p4rhbGgMmTBGK6FJ9ePnYZDepqZLqxhPckD07BP/WFKVW/VpGI3O
IA+xgTWI3N3ySsQq1abxxah3j1+XL30JC8QVWWbci0aFaVxzjHlD82eWBMuLQ7lL
I8p9RKU3QRl9JXDsRuzljzD8dP/iM79EldtL1V4ZcUPwySRmVWYXM/219p9T8Jrq
WHKQgoFht1ZojxZawL9/HVtCjGuCAIcBgx+q7rQVUQAW+Pq1Rjk3T+CrPT9NO+X9
nTLfztvtXnCSvyCCSMB4lb6+owk1N3MiaFG3dLWEi1BTeIccZlNEoSyIUH2c8EVB
h4O0omCmJhwFXLQcI4sKOjjGVwg342D9iyywUuGCfXX9fJ8Zv1oS7U/dFmbZnrkv
EzsfdDMc8lEB9sZk46AC2+t3gKx9xhZC7t5mkHDa5CltthYbaiuWZ969DH+TalTI
HmGgqLcLZyufDAr6PrzW0aEPu6B5VRhQwPhbY92Wz1nlAgf7dFgneb4EbzlrTm39
Xejh+ZTezb/2j21n4l+2nWE3HRh4tlS7fDZYTFPNZIPGB4tHqomaaSNd526CH9Xj
/hIGRY5Kjp4bE075gUTRF/gygepfya46WNZYlLjANbfJfn3joDuaKviuEJGWMSqy
1alPQ46blGsPJ5Tr8Quk6j8PkcPr9nIzrkDVbUEOgV5H+NByeLVEM85D66EiB16/
frbtIXz47Vzr6QRHfXYKD3aYRVTsZPHhfRyN3Al0YZz/DV7NqdRHaDzmeIJxpu3A
AnnbjUBBTL+A0VBri7RHa2MPl3xxNX2yxL5zQtvKVOiX2TQTDWT/GytQaE0rZ62Y
m3lXMqA8bVuHAGPfzYphXU5RLerV8IUwfWSsIJz7YLntF5LEDvM5xF1UNxSxNOdc
mjlhNfT4ZcdJVcRaUZJYOp/ZucB5L1+OAOl3IiKe+8gMwt8OhhJy5f9LUjhaP3Fi
v8LRaKbhYqGvedGH4nCq4EPUyDe70xcQObYA5aAgZwoYBEFh6A+ttAaQswT61DUw
+63Th0F6l0wz8ueD/J5H9yvVPVh5I69EJgzUjqmUT/L21KE0jnL+YdgtitVUtx32
2cqTiiEL772hxiqwxdJ77UsmRgHY44MDTvwbcRPi/nQ0t+hY7jlH4Daw2tiYxYtv
CORwn36BcAjhiC0nkmSEBpPOvic/ygeMjN2I5SXMTJWBvs0gimped33+zMp+SxUm
nK25Fwa+mOM0skLWUAsjXJXcAPpmzibgdynwTsbyl5ZPVsGUeeD/wyR93B8E29hN
KwHNGiHLf0ovGWh9bixCdzEre4qicS48qocMj4gh85znpcDOA8EIq30ViB5M//qC
1go1xnhvgX8ga4I7wza/N9iT4ookVrqz1NiAk7CsuAx9XhLzvVXIX+y7bPpu8J3i
fElHudTBNdeNew0K944SooyNkzSj6v41tbj0bucNMATnD7UMU5yK2vVl3GtMQhri
6dr/9472QpxB584spYrbCWCNJo/sorZAaniHBUNeZQEzfMNEGjsqQ9nmZyTMZlCe
GRA9HLCHbfQI/PzE7Y9PG65amqy+hm05vCSKoNCpIxq/WanIAPkN3yd9bHtMUM6N
M0eycZBTUXwPClCXL9d8y+KpjPqp3ihuGtmUxb16HZ2zkj5UJv/oMU62tCJWSAuh
KezlrhggijDxXGje2XpgygVMw7mNKMQb+5ej+tEW5puzOyNnOAaItofRWv4E3dAT
toIiBSv70E8898W8JpH4snMaUUtL7T2DszJrzuMfoorNrYZkSnacBgYTYZokclpO
B9oteQENk9M9jHiHwgak3qvwllK8/18eSAWZ68/69AjBnJuAhmn2iWSUMky/H6q6
NZCIesk+CAb/BTdZ6CMnis3F/SDRlT7QqhmAPxjEb+4aV/qP7YIEeKH2JGPBZe1u
ZL+1yihe7jfq+yofgSHyART/L1a7PQ1QT9vfWr0/gMk9vB/lTZDHRa28QxqW0t7g
IPi1bo6JvlTFwiyjOjZrkcXuwPoqiae/Wpd+jfIlgmEYnDjnR1lSf1/hNYPip9dN
DFYGrZ4S5W85eFV4LJwASOet0yTcxBbLhTAxvmyWu8cwIUNq2mfyqikDK8iA7FwA
vjECR5j0YodKCGVK0jA6Ris2S1OrUyBKcZgPBLC2DY1X/Py/7Lo82QFncR0XU3Nc
inczO22fGYmBvnzysPQfpBlfmCxPpaWFL/W2JLb/w6nbjpF8dEywEFAT3x6ZkUWU
dOKasDiZCSJ2LeXqjP3nLJRnKJSQlaAzzVp4Aid1CgOAfNsBNqWl7RlEwYUYHmU5
dJRIi+B9XSRcg4zQblrsYiPN9ryYxTmk91mifYyCGUrVs2A/IGjfyjs4ATAxzP1t
0DfGLbY/G28kafCFW3rxJfcvat7Wm3Ew13gzJhYwuN+BJ2PRXDArPUOOGNt+g0KC
+E9JlBBPOoaPRfAEJZMFdhrW9c7hcAFyX/hn2yUs4ypw6hoLqlrbgzrHT4mB2bdx
kSrvC04ZTa7v2QB11Febam0TboLr6hM/B5/c/wvbstz02QG/XbWF0pCiWBTX9ZvO
SD19kEed+hl3TeXHOQvChlQ5ZkjOzCsZ06WxxZJ22RYN/GRqAjxosdOrd8pkuEqO
mXnYjUYcaNrkYwU6mkfwGvdg1pPRhd4tqOFIOSH6y9YZR8bStkIEP2rsQ8j2N2KH
vo/Z9jpKH/2BjVCm9CvxAC8m1IKE0iS8QjqpFIpQiwafFj56DOZxBrwE/dTVTOQ0
poq8D7hz8CYcn3D/61nVdKf/0USrRp2s+mxSpb2DsFGp1vpsqtWkkk+yifTO0thG
HHgJeDy1HkUbiqyDlq+jDNuLRAcX5WNP/vQ/vVE5v/DlRP9NUnif6/7MBhdDBk4T
3z5e+Ry0hQIviZSVcU7kjZAyMFvEAwnI2jeuvXYwVpLKkLkTux3sT6OvWFNF86CA
OzBZYfgW77HokXk8Fid0XDTqmMdDS4J14aKfxWMkCh1VZ8BVz2I3fUpVAhqQCHzf
ic5kHsHRPCNfqbbsajm5e001nVVAmqAAI4EdJSBHXKK4H9M3PP9BkQ0zdtuWco6v
hoVATzbdkGbShHgKWXSntznq2+Pv9w1TCu2QbBBbC7Qlj5eEHXxSDAw0Pf5gqFZo
aACOMqdShfC2MtPYO8b/uE1cnIM5/nXyx8595xGcp+UNmxjIe4YOVb8xXIM4ioNf
pVcp7BevGtwLDHX+QyVA8/1uqFo1Yqf+Ebt8gcGwnZvLSJaS+q05WvKWCGstX7A0
+tY3SRKr+fjqWPY9WwKB/EFc6MlZrxqSVMOLrAxuZWb3NzL+zJfFKXTyD3a/vlA5
Uhghv+CP7Tstp0aKzfo/vI8PaPp4Cyqg4xsA8ZcFOEwoFKrfV1Hcx97UWOyZ6o4k
xZz/CbDpPo90Y3nX++G7jD0rpWlBGwOVOgV8H3ZJoAaU5ScoAvp+RbVaMhRhn+4R
ItMD6IUj4xVOCZxCURGQOfJ3QrVdG1KEwdH6bj+jSIbaM7hcM6pIkOPBPJBGYHpL
SyBHoT2PQ5a0ZRZgqv+3FY4K54ftq/rGzotenv0PFJ7pVMJ35lz3iJeo6FRafhJ7
Z7ZgwgKBWFDCSx+KEvKz1LHr+BOehKT9LgQTwryBLF2GW1hJOdkTZsEZbZ7QhC8K
DQS5e5oBuXHJ9TWmJBCzmFKXJsjMKOZDRYcQitHJtwGSWoSMwsSLXW57Q8Juuinu
PHrpE4uILQR7QRgvGEhpVazzQzeZoqqC4GWXmfWRkiwbrg3Oglj9ZO7ro9AynsAJ
ZmFVPaseXK6MSR5JCJr/rQYpQ5hweUkWrUDEbVCHJe/jq9lng5Wb3ZFK7uZqjOHh
q+PyxHwKimTfsWor4yJ8Aqc/6ZeBLxeFiAnObb/8qqzbbznAfilKtDAC1R/JEQfN
gk6kuJ6z2ry5hB3jCDbYkwyitJg4UardkpdupphV+G9znwimk5abiuIqr4eYh+uQ
BDE3pmHSiIoX9+pPIXYzsp4YViJsHxn1z2CpLH0FAped1i+/5b1WAuOWwwIVbyYf
3YvKa7kk8jdTPQyoXTnTd2S7LukMAi3ulncWlAbomn+LKTiUXx2fnm1Ojqx9hLrv
6zCt3ySkk8AufoqGr1K9ucYH8T0UI+XRnyieX8WaBL07QBAMmy/OgjgCYwFE9sT/
o0b5IA3Or728CrYhandAd10Jc6884ol8ZiSirYZIJZWgeEwdY219Y3jf9lUcxzFO
r36gI4j39xza5IxePStjp3tsWE5zuESeIZX6XBOuHveiYAXC2Kv7UVk8tLMYSdhq
glOnjkgEy+gZGW6zPctr+oJillOHEVVz3jgxm76/BQNgvVjWfZabVLZj/gCuCcqT
lAQ0nNvS/fPQfV39hMvIK767qCSSPr2/sHvYxk8A9neoifE+fKzjD96DgiBzmcMO
Xr6FqK7KgO/2ve30B1V8J3CHAIndOLwF2087I6GgGIW4Zbzg+CCDsrHlQREEt6uE
gSdjgWTabOGG90cGNIynuPOj3ioOJqdBp5wbUXWt0Ddi415t2NMIK1XiWwtX6BeW
lskkvsZIqZatqu4pp1+WzFvEopi1m/fcLfbmIOu1IFofPAPwq2uKfM3WXGJY4yfu
QaltLJV2Ei/ZnLKAwd9TmVomFZ3vi+4b3xmzJORH1R6Yx3L/0A75pjL/gL2Y/pbB
gyFDbn4bnZzMJJgQF1UjFy2upd/khc98TEY8SKYBuhAVDQJ8o99gse+ix/clvUl8
7eLgTBy5vO4x/AzBbaOx8lkeBqPBg8AECazGhpDhAqK0lPz/whiPHfIbCmqFEYFs
vfsqmy4KIbffvLUMS61EBO0kQp24qeSKgjpXHPdwFQ/ZV1C8lNZ+uH/R7KyDM6bJ
dw2sFwPQy32o4hearWnhy2UbG+qkeDb1XQ4IYhuAD3c5Ginn+YEdGVUpgSMsIO0z
oXGfIukuK6UVbkpWJFX3KN+FXgdMCyb653zu7OV9Wsf4J3qRdpEJUaTCMVL7Jtd6
BK8LBZiCFOcgM792vkSVxib+sX9SGZaJ+L2iSritFiqBhH4Gvxlm9HgkdxjxrThx
R+XUiLOUy7oGNRTi/PCf7FKcRf30lH3vFDvpdxnx4m9QPucrI/Bi5Q/5MjQFX9GK
TbLT3ek/BOp/XRu3sPoQTE2K1FFMpocaUWXSjcbjqVylPUYWc0JBHICc5EbBQQWi
fdKVBIsd/ESc6gwgnZYIbvy3addxwgXj2+DM/I414cpWYJm2WC9MTodNoZ1Xom5L
dxOQyMgplg14z79UBkAQIjbNjZRyhipTz2CyRjcrpo1BqaDvV0mUUipF7bJuBcF8
ePEgmNuF0pMM/6R0hHuFejy36ysle4jooDW19BtRTXqM1Fvat5JEw3G7Aix3kE//
PttKl6jNg4RTp24eiR6d+3tZWjNRpAyxY7a8asYhLi0xuBGJoJS9iff9wc8QP9uf
cZlOmZEwIYzQQo432J8Elj91ouasbKv3+d/+0kVWYrIF1eBZEt7YMbSJGQhYIwJJ
BjoBNJLdDvWibXN0qVpe6sET8w4V44eBqxvn6+/zStHZ+98Rh/9toZxx+swN1TuQ
15BWBv4CzyGmR7EJn9aflXhXsIAj61SwUFE3O5SP0Aj2/aY1G9SpIJObmwgFjKvT
B1uuQ91vYPOqZtqK2ms7y3NsgOP/pRh1UWJys2gxcnrtyCTrKjCwmPYbZDatnrBu
e+/7arz/Wj2nl7pHOKukJa7Jbpqx+AQyCmaVIdFnRhOpWGZUbjHmmaUClMtqXfhD
XPheUIfkZORd+b+qze6aMFnic4ER1qs42dv8OAFGgBeV9CeY2JP+7uywYteNiOf5
/A7ec3VIrWOgzRT8AWRxdMWXJvn6S+g5N9LqzIEGHT0yPU/6EZ1qIoVChxRZ4QTC
b5LgL23lAJ3QQkJ+vDitLQ0YCqate04dNRmSWNBN25gAC/HfqbC0x5tarZnrCwex
xufp6FUIkhO6n0bpNW4OYW3GEVSqAH8qji85jEYugEiVBUgG6URx2Tvf3z3gnBP7
iqB0IxGxEg2fTpT9fcA2NEG6LspsucTpNZaUks7/F10RJ7evleiVJm+NnSrL/SPu
FPqpyuPJpmJY5sK1IhGgtVa+10MoIDYL4D9sQTaPmFgft/OlRRkaDe1vzJTwBCRA
TqdO0BoiLcir4AgkFSVSg9YIBr+4mQg/Dwl1kRJDH+f7eEcQ6Ffl0X7jwRQv5NFY
Byd+tsQkLkWw7UNCTdrAK0dotfGuSY5Y9L7f9BrBwrcBe65qd6ya0gbVsgzKR6wS
FLf+TQE4pMXuEWqeKJNS+0ecVhdKjlPis6L1fn37Y+rDTEaJywwOoYmqv/YI4Oif
J1MXwzHJCMduoqoQ4Eb+BGd6nfqcb61mdnhByrraYP8pELuLhXxnVhBvRBIhSEG5
rH9OUmlWV+RbopfLG4v5Bn6OASoUSraw6DFthUYXISqG/YoLMP4F8fyWDgHJowPa
AmgIes1xeXeK/utrPak3zhrJVODYuZoR38n4NZNXxkgVwNqBKGrbFGaiLjNh0hQ1
a+MWtUJinJNXe/mMGgGr/Kupqu+mPWN4Qe2xFjpmiOjTprWIMrJi9NT8Kr5Ou7DJ
mvafWTkEfSC09UgTgvOUZBJGM+gQa4gC21piZi3ezenANAhcRu1PKhzVFfJkN/gy
BzitaeAluwe8fKLtItnsR8ws9Ijj/R3TeIX4sv0SZScfU1btpLSkHHbPGErdeIgq
IToXBvHl5P5D5c6t/qGEAhPPhzpCOL7oQrB+jPWGYK28XvmsGLaOdTD6kF5lbpGv
DNPsirIaubGcKwBPVoxoukQ+xdv0qsD3bQ+rV/ozJal6bZla0XExZ0sjn/N/6LwC
l8DI31TSx7TthOOKw64dbJkHLz2BS7IiN9sfg+k07qkHMTrIEO7ZGGgF8x6f7wPc
ghn0FxhtoickQdErTh++AK3fUUUHT4XLigFZTp6mGhnq7BKGp9uKCLUanpU2R1SG
FacvIDq0Jjo4/uzZWXLYlOR8hfcf+iTaEDwlpiGws3muSkYJS25atdsADNbMYFKC
j6v9EoDS8BLRjoWDZUIhPN3Yz+sGWxDiHvj8EXAWGfyWzSisIHQCjTdVBfUov+1z
LqfNHUH45975l/f35TrtlePtX6RiiESymgyc9waowBEHTweqao0Vy1DGSApzJTQm
sE2mfdgQnxQhQOXHHSI15UlkbcFqUp1FhCk5/KmuJmN6AU5cBuZQxTJNnYrpT4Ne
+diCbajyqcTiC53knYDKhja+H7iKbQlrs7c0A+ttWBzUUR+35Iyc4ZHK4YoXJfzT
AfR1S22Y2Mf/IEJ3oJleas6CfE3DxUxHENjtW8iWUPuh9ogBH5FNEiVItzZNYl0A
8ieH6eEYt8OE/elh6CSHY2t5Wx/mynRg1cXK0dxUoydWZRJSWTInKmhWHfkJyH1F
CpsIAV67MWwpt78e3iwaXF2vFRhJCy8dIW5mwApbuNPbUqc5NW8fG0kPJwsHOmfM
C7mWQtJdsztTJW82Qf4fZ0H2mV0Mx2G4egSHMw9K+AoyUvg1ubyCJR64f7KZpSSa
3GawloAWrQ4S6gXc8qDkWE3WuYWL8rvKeF+VHCratszEr1Ms28lcas4zaodj0LTj
D0JJtmPWBDc2/lOF93EQNoIdeQOTLbA8lRYbVD3S9oJhSws1S+9zxtR0gfVcbWSr
Xz0iUrmqZK/Gagnc/LGWBnjEqXiywTzyJwEqCCajpBGot0jeBtgGOAoCphU+B2C9
6mOzhg+YcEegwKEGIO+jbmSht257wjK9NiaR1FTjBwKfr7MHC0COOS5EbFY31CsF
qRFR1PRp2ek9TWHOKxy15Ymfq1QCVQKnUY1y/RNrR6medaO5RlZ9mc/5zGE6H1jM
npWxd8FoMiO1tjEWXhyzSJBwEoLaUjAbpfej/cUG4zbfsY70O5CQmYWbX5pYiBmL
0SMJZxgivGfTZb0n/5kld43TCIeqKCAXkKF0owAEQ3TJNZsIIHMNjDS1+ApXDUyd
kt8hnYp0W4rJnemD/rCVHbS2ZbQJO5n6J8BfWzfIt90ltp/rOr0lQa/Ng7WN61je
v1uLNL/wodlJiZWCK5sPBG8RJxaPKXUPGa7nRVAiwLKftxxeYq8qXzpBxDC/5yrR
JXLrMOBn0LBu0pfE3XPBDW+hGXKRfrx5uEzWNG55MR73jpeh03qJskfRynL5rK4X
E9VTI0DlqoBFqSQjUpvVuFUn7Evfn6DNyU7h2fKxhQQO51Rzwa61lN6S6IMfOLdO
2QOCYmKtqPxgZsEz7yq5iVFXdWRobyaae0s+pB1mXc+/X69mFJjV31uTRO2c9U6W
qbxIPN1/EKh/n4aQA419sAmxwE4mieeqsT//JurveasjU2wmetmLAbZfS7T9VprD
b7IJPx5CTDJGBEZScm/VNOIRzkysuXzGKcdNJRq5ym8vD4MKGOvo0AUU4/VTXDbT
tF+WbCFN9jUyR2IGlifDCYlc2jmiIthpaRNcvPlKGdNo1EBWfCxthBjYyRf86PVp
GwYIuHDTOVfXxS9addAJpVMJngU58q5p+t1UvD/6ePU/kF75KG8kvdPreoZ216vw
pj0Nu8J4eScBnBHQmOJ4XwPQa3k0f54kH7d6zlrhpSjQpaGfXwqbUQQn971bD9/k
e0lqabs8EgyBmpx/rES0ZtXNDdlf+t5GprVoMf1WM3HpmuevJpEa4+cmXeluUY4l
lbO4ZXMPqWeb1j2MI9lkkkPtY0B8oGoJx9hbV++IwbfXQoAbKcgJfVblGmI76RKU
HTwDH3BZnw4lDE4oLHnZGUTMwAsEWVQAU1OBahF81yeXqQEi4RDJ0RUCSAtVvJIs
kTRyz/vaDdFfJ8uygti1U/iJWtLoXY5wAhifjSnB+mv92cBRLPSpTnXDcEYpVD8E
4BPz4yzMUfNBHVl83Kw3vanChTZRBHigDfRv1nV1jkPxKL3G/94Bt7BSpcsQhrTS
UT24wtxMgoVYj9vuldGgUVWOJPO6YmIir3CjHBywJUr+9/miJ+RjGkSqx3mF8pmN
0GUfhMvp+A5Pa9ap4FIqK9phk8O6CqEOkPz2QxdzJEnPtks7oK1O/Tlyaeoq+2Hs
RWjjH/BNtaswk++zR/o7huCDpzpDRZAzxpd8XsnI4hx6TMIi0QNA5+EcArUcq7QP
bQRXEGCtEtAVsJiak5eDgM2LJNoYTqSLup7XcH/FGjZSkr/wHTNuRzm6rsV8jBpk
6PSGpvLNoQsSfDLm8ZN4NLTCPW6k92LmxCKYQnmB29J2wodQ22yl8AuiianwZMwN
AibxpYcYWAHZcF0M+8vxCFKfXfzNPx6PdlWJE7w90xGQxbN/Q/oR4DIXJwWDJZsO
JtNtkYkvRgFdegS8+NNDRQdIDxDNsKsGIGvwRETNXSTu1veeMjj63u9j+tuulXjU
b8c5VmMlgV1ra0imCOgFc+YN7Tq/VfQu0UNE8yr5QV2KzB2qpWRtBUIGAZi11q8a
PlcMuyGkFyIY5FWDIdCp55HX3q6QLMUCYZPJErvjEchOQxaw7OdavR80HobP0yrC
z3PgToLx9qIHt+I7v+0FYISpmXXZyfsYc9uxkTcD5WQ6I/izQW77lIbB306tjubO
pjZCcK+76iRyWk0AXUpEYsbUOBlmpdgw6xfXxLoftXeixlT3oAtAqPpc5+fHRZxK
FKVKObUEf0Nz1ShcD53phtwzmQ4QYEk9auCXNwQvGsQyI1mWI64LK13E9ck9f84u
JnzMWCNhrK8sHMMJGOg3/YfK83VoXMJoCEn2XDbjueSsUFxGmamgHBQ9mBYkX1U+
C1snJEzYiMNXJ6u+yC/i+gOHPqv7t2JHK1Avp4gDaaRh6dfq7ZRORlY4frCqkXAx
3vq28RNCry2G9anmoeszxFwsSgz0Kl96fAUExLRy9FnKammrLXJpPPUGFIS/LJ+t
oHxYiwcnDWpJZMvOV/dXWIgnxciAtZ3vnkMhXR8kbITeM4ff+4tgi/mk/KPR0fsx
trFGxzfph5IJUVf/PRnFj2egPMxiVrliXVFIFQEFeT0Gp3UorwGFvaJtZG/yi44b
tT1pZhZkrrMG1w1S1+4xIq0KEIe+U/giUvhMy8wxdbkUcZk3Or/NvNT/EHEWjmLB
LS1Ws6XJheK7Whek2g4/fKaVvRyFHwx2/rokuLnYcDixoAKzU7QrZKZcgad1Hytf
QlzqNiqXp2awmN5Ca9oV0wGYkGn1EknOa8Zun42qxvvwmikkrzNzGc5qeOmZxLDX
C+lcPhMp1HFTezcskck/T6Ps6Jrrl4FQaUmLkcBXPkaHLph6hDlncc6l6mzcwejR
FyowcJm65rrAKHH4yeIpKvKKPDDcLnxMIwRdFu5fOFQuluy5XCtiaWVgm0V0NmHc
GdXqg/rys/vuTrPiE35JHo/A+AvVpxrGs6spMx6OdU7MG+hWVfj2yhTyz4GzX8hU
ZkSRkbrhH23KTz2kfjXbYjG8pGlg/x5ZKz3lQx3Vdapte1/2LvIUqukaQsPzMoJ2
T3iAXEVz8mAi8vGgHzhKBT5X1jyUCMWQiWjpiEr3MS1DqVxVyCHJGt1Gjq1tbOzg
GtgphhBdKfGucxnOFaN8QTVq2EB6/qRzT5nLvAL3cDLfmzkVJm2XN4ySz59N8tKt
ywtRDfwXD7zPKjSvcYebiFW7gXSVZUeHDlDdVHvKQL7xBzCAjb49Nt++TEBfO46X
VjNvMHEGkkg1R/RRKFvAI7c44B2J+xl6FFB57vqlxpkQ+Z8rMuECyPjij29NtCs1
UTvvw18kvODEyy2/X3Eec67niAP1n1PHnacTnFvKcp17Z/QDCmQ/KxonJLF3MqfZ
ljrFcr6AyU5hVtBKuca/oRe6OyVpC5ZSUxyVb9caTYntIDhpvY5U8rr09Yd4cLIK
ErYZpM/yJFz99GLibWLIqYa4Lnp7uGUQTa2K+zptrKROrRXkqRt6SAByq6C/BkFc
higGQqr0TMtSl8cj+4ABbALrdQyZoOnYO7+GcF92dmNK4GqLCh3dl1m4s8g+hQyk
aLJwY9m9c8XqFopitFYyeTSzotmLoF8LO3zVs0RHzYBZ8Yb52IPENwAAJ7bUyciG
MuYKXOqLDasgbY7/7KFnq/71H1+hhT9IZ5bSGEtqIF55t53tJ+1pbkGubjkF4SLN
RI3jNPFfgVOO8gVos33HTT5bU2NnHBFpX26HOQUOIEO/A4EMSJn5uu3JsZa/w3OV
fISU/nwej5rHJKHcN5FLJNFWSyhAuh9mWHU2dWfnHYi1irCp1Zadfde1wD890kAS
F5eYlYUS/7Fc+J9liQiUWCLxK2i3nZXqekPUNfPc0tbxvdcwHSlFpwNtKmK0pde8
81Wnu2/xa+i/e5NffB65+blkAG/2AaOZRl7ye8IqbaowHF2ANpiRuWbcUSaJLWQJ
8fUSuomnyUjihji3LgI9scrTKKjjy7zItJfE10wIckPbMfZrdulineqw2E66uXnR
tk0lUJWDPS3Vf82DUrK9XehVNa8RBlZ9ZIBQteZdXibXwcuxqvqlMPuYFo4rqyRb
Yym+19PCRt8+U1Paf6c8jdSwNdCjd/4ZPnH8s9z+Qs7j5FxKEV1/OBdDO+BgLts5
0ZNFuTCMmdGtArbAHYkdhZc6LtiTZ+HrPR6PYnKdTRtPbn67yVUJRujn/sw4NiAG
CosfeXMfp8FGjHsvy/dvunABWAEs8+0APra3Vlr5VQZEbJSAy4y4T/SSAFOl/gor
DP1XOPa07qucKueLk5PWgLwsTRTx3R7DHLRS0+/w6UvtWyTEyRVu9qfhQN0YGNMW
XPzB/mdjhEn+xjMKFqnhNzwbKVruM62K9Q9Y5Zb54HJD1tAoCqR/RSzyvMe3swDI
dayLLqHG/Nieb1RNsyZm705DH43LZrInUadf05WVxi+9qefrCf0hPBGl0HV7wbu0
zah2sgAdY11o7VdJ2/VxN8z0weZy0F+4lnFHunXnXO//jiwCarlT5TOxjNw16D/g
SgoXRBf7YHI+zdDWSDQhok/jiHGNCIg9CzFZVhKGwUTKOLMh7otGA5Tg7hB7b3G3
XxZdY32za9oB7VBZU8k0eBi7C13lKHQvnc1LbejcvvTjrQ32KJzvTDhp0Iu3rgPf
m3h+CiyLHIIQThh9mBWwpe+xJyDhHdqtpyr5sfesCLrCWyyviMe7hzEHXlKWuCtg
PEs20MkhGeMhMRnl/nm6IsixAvLqOWrBVyXqpYz0VcVUWstKBZCQntV/xYWUTT7h
W6BQ+H4x2ihR20/fris7JPiLAd5YFdjaZ0pn5tNMZh1MMdZ3svW6mPsVlELM3G4S
2Ts7FQswNPIAKwlq6Ii6oDR6kJO499NREREki96QNJU1UNN9BRlYy0Ym1yFu8clM
6xNF4O5JvmNu/lMgKOKJ3AqBQ0kfjKdp79yJpIb6zDd50sjPmpO2K/bsqS3Vcv8c
NShiH99ZDDotA+8IAddeZ4EvGtcGT0hK1ipSiNF6j/dJPXIzz+EqnU6ccILcIzRO
JVGLZ4P2srAJDI4DZU0Cl3gT/u+Dr4qq/BsbC/G0r2vraJuOQ25i9hqoSlo4ttES
y7T7DlD0SXR9gfHDaMwa21OBrg0+I8Sz3O2GcbR5p0yQtTM/XopqhwxgzSAkNwuf
0vQbm2S1jLrFMaaHQiOaAfhh04eeSiqUjF4nNVjgE4h9+gOQ4/2bEZJDK9ULFiux
0gl49/cB6lrbTuCteeW1aVKOFQLiNyWfjwNjhyqegQy6LhgXtcZuPTXMDiaz7kNM
l5sDMfPdlQ9i7MpVkJVdQOuV1n8bj87nP/UUf1Omm0/7y5MbB1jpAlJwaQiYldMt
eti23loGOxyLRQR1qQxSu3m8sI11iQDBqb9n4a7rAyRVvfQ+gWQyz8eIkEetKNql
rRIgxZv944IArCV3vs2GCouWBDSKphJkIiy43zfZ7suVO8UWUEymkNypjwBfx9UW
cLLGGs1IFzm1QM7mscSZZYn6OQe2T3dFX3EUGQCNQO2/UvG9p1kDsWBsvW3RgJgG
u0g+ecnvkAdIennQlmLB1hnciCG0ivuHXobRAXzV24/2HeVy2QZhFUjDngMBf7kj
BKIhZ+pySy+/4tBBrnxW/1hSDedEUe6EFosNqXTqlEdDEn2diSU5utpdkplp1OzK
YIofJKRw3CitrFwFqb6P7vHBAWsHvq9kngmNeJfEClZCQ6f3Un2V89Abl9WHozWN
FiDxaI5+20k0piAcp59X4c7gcv9aauaUIdGymJC0hjFN3iqxbeaHMuMoWB3TRkmz
85rDUw3hhXCGlMK0bv9fCazQDZnRH30rkB7ISu2IsNkez4H9HtnOpWelNMLSoZMi
MdlcJhWIcgaR7mn5Q5AIzbYbsWir1Cl2GDoMF6C17/+m5Luhyg38j5mLxQ84Iap0
+89sU8ytJnGmRAg8E0nFUHPHFesnBjio77hKJQk/AKstD9mxl86yV1NdQNHZTQJt
+34ffoa/aSAFncByn2z7mda/MWpk3kjFspKkRJKBoYBlsoOmehLKaqojli0H4sqY
4Oll1QcBU1H5Bl8vdZGfhplCEaaCo1uoP2K4N2hmh9f2xQHFBHq6mIxJIJ27vIGu
TJ8O5MC+pzI11pzI2JloV0fu7vea73e1aBMWOK1dq6hbSx8vkmdMzNer53LaZy4W
ip/3dm1iBwfJG9tDdwN64+yjjhvxDg0RKcz8y9taDvGMh96HfZeS/q6lCcsp4hHy
E+RfdngUz41enZZocnxfrTnYCXc2naFgUe8SQoFO90+iRJimQGd5k6m4N4n/8eel
TQztVzdjeSv+vPzQO2h+/M134H+/MWB50RvwUT1o+k3pJ/tQu6FUQQkSin7Ik3+1
4dItxZzXqq5V11uc/AiAqQmkjOlT1OrtpZGYAz0BpD+x/7D86hn94YGcKtjoB5Rw
5F7uiTWxtZuzUjGNQQTOap+Ged+QKYVzoXeXGN65emGP9GyA0h75IHMaAdtepSHq
tdzyyCcrRJgT5E9tArjn1ez2dPAIu8cvlEmf5dFkLHYI0rDcMiIpscsyGnaSJDTP
EVPiyaUMkgbdkM2vrxAVyc+6D+XaQdeVzNiguaKZvOphz9MzfiS6a6IVYtXhk0/K
QkSLBj49hu7J5BSHBPl3byLLkkxWQGjxcc/tFmxVUSK+ZahpoAnUqaTmvwSh7wyK
YrbidaaYViOOH7IBwtKMd2jcBipbly1lW6Lp8lT7VuCDlzuHmcZImnDRtP1oASh6
YVE+hQheXb81WLxZWcP0NH+R1Xn8tasbfv4b6Ma94FYrY7jOFPAh+pSOyI3e6l1Q
vIplc+tS00hpNOiHvgKpMm3BwITEtgkqlx2IxjLCMzdV1xIoC+D7wMNYLx+xQfRZ
QwQEHq/AJP376fdoM1US8pGvtjEsIqtJaxGWnzmsfuxszleQBh9nWBfNQfy7JT1Q
vvPZNoDpBUTAxe6HEcLv3XNwr886XAIg5rP4S5NK3/qmeo1pF4KnKE4nsyMioN80
5U+1knnkq8aY/OBcKPc097bgw70ysKJkb4fvnNoDC0PkZbz8UoKkCOoKdEwPHGZv
xI0GugfUHDX16MnFFyBk3DBynjr66VHfyRUERd1ANzb/v7pD3gRzP7O1Q2NS72Ut
TW3FIAWVzxg/d1zBXRMulxUzXSuAKTLq2o0cn8xun2OdDj1m+OeWiIE56j806ldn
ys9pXzwVvS64GWyYjYepzcYAR78/CZ/SUiqq7mSpdNFQtCkP+BVZ5Okl64VMIfv1
yJo6RVGCt9J6yy90ImdASNb2b2+HvW5A4RF/HoNgeS6+FKBOVj5QY9MJuLwhNW8Q
8YzzEtLP2WMxWaDrvYCN8Fnc7HnONMcfELcBpm3syJCIZAkCsnOta+QTnQDSvUqN
RHIUak5/T9AvfA60pLVSdKOlMhLlKzxDRSe03TEX4TSzaipU0GqRaxtqiS9jw5KO
2YBCOc2qaU1I5zuytnX7ADiNHS8cvBfvFavsaxyHyCXfU1o2G1DQR1IRPeLuTi6P
0ycndVN+1Cb3E57gtvfIxZFl5Inq6cWM9CIR1ea4Gn5dWVStvbZ/546p2bpfYraA
NsIamPyRxfSa8hPzXpMkA7MUPKR/TPOXuiGBqKD94SgxMwsTNAgN+NRZajc8UF7H
7XEMXmz4SaaVL9KfTOjkHHNhPx+2MPTFCxicbCDKjyEvGP1aXnWPY3cbaBmdfAhe
whKdtjxXmpkRnSeg+tiQiypdeqt8BV+oKsa/KURA8FfH7/tPoHy22fT8HRQsSONl
1upPOBwDVqmBxRhzWF37EVd/56jAY2+r3lotcqt4NI5g+BIO6M6T2OAX5UqQVAIF
DInLAA3sWZnmhfLdBx2GcOUjR0Vq4+3sgEU8JCT16llYTlMQX/k52QVxhvjja4Cg
DMW/OIGS730xtwMiq5VRVGjwOWyDMolpwTel27FnLYx/WqHBc+7bNdhTa8PDejAv
J3U6v18prEkgtlckYSmg/fj8SVKdL3moGr2mgan1Q0CnMrPER9lMExNXe3KrpzhS
m1EBGnSwdYI5ig7MXqf/uuborHJCd8iibGEUyjY+hdkN0VDGyYPhqLct+7+F6480
T0DTD/3ZBK1Djuj1CDgKx+n3gcw0MbCA+1zLqKGPW3RsNRhbu253QD32txyqyS5o
o/d+VHa3KhuGVWaqUvhAI0xIOT/3t9GxRRIPni6x+nWngK2ZPzQJ89sdnQOGlsPR
IJUG5MJayke2JzdQ1EP2yc41mI1qhw3AsNQdqVDak4uMWAswCZJ6SAEDJhODP2Yk
bY2vcfXljQBC8pt+XCb2VLBIvBz8i0uwuUvf/xnapE0u/uyWIxBleOnrVeq01wbK
f0F/sNVi/J/LpoaZNND9bafsuvqjcbdqYYSV2pXa1trRp5yQmHq/ezMUd/xb33Yk
vYJ/XhrdUTlaC+O1N68OQbdbiJgX0ZR3GFm3m2tJlI/TAEygCSGH5bBhmU0R1P1N
h38LulN6WeKgX/+Pc5EpX1AkVwBtioydMlWN4A31QlNmEOwvG4jq4Qg4W+H+erqf
CE0VWX/kJDPtDnz3g1lO935X19SNdvuh++DGFhUAfZ6jeLpL298gedPu42tWEmjs
2iOZk6cIY/8sacvrg2L9tkvrNz+cu8Bs5edRCjVX+6pN7tN4mP/cPVu/aNzO4rtZ
jchX1DzkQMORJyJ9ywj7bRPKRQsQ5o6cIGVr43HriTjosX2VDhrVsXgGc7TtceZl
mNhNW0bshDIDOJaCf3mvMv+tg6pXJtvLIYQlLf9R5cK6CmWS6zu09eKC2v7q9M69
NWRs83ssL6K04oBFRQwCXUMLp2TIhYooZCa12FyQNFB9vY8U1y8AUpm7gKf/gSOK
X7/DmT4TIAPjj0c0JCBcQQDw+wAbpZ0rrAPrUVp+qXQ/jI5xsW87HzzWya9kLRgy
v2rZ7zwZR3JARq12Acl8E49QcTv5Yw8/ADTyeCRrvGyvaynKfd6IqUP53QjGutZc
F6l65PcXJh4kmNowZ7WWJX9zX4lewSmVvgyf866GBffHmUjrVhAeEH3v25rnRguK
CJM9CfEuFVFrIkeYBfZ9VLz14AzXsa8QYUsrETkuNA4AFGREgLm0Ls/J0Mzfx5ll
RdwtP6/1H/8FRGz8sTUSboe7xZ0ES84Q0YEKk5amyGEc2nuz7IVcwF4h1N8mDfW6
j/Mj4nT0CskuRfD1Q1OsvLrAc23Bsm3Ol72NErIReqkEJ5Yxa7f8q7KOf/X/jMOc
16zo1+DAoEAgLwTpsQHDiUwcU3HozTj1td2ff3gZ1+3uPYI7BYvfh5IiKxRwybGL
k3NQy0/22P5nmnPYnXeA93vd9kZy+cbQ2EneeEqQYQi58qQpQDWjtrGwjZGPkY9F
ZMO6bpkhDn/QKRVQfEi0C0wY6qdJ1jmXZkS5ouOAzjZW2wPGn8YlbVYaHWSKDqC8
qBcpt/l4xwknEFUazNX+HtjG0aNpb8wSfKmP0MS1lJCCiP5tS37U5XmEc/6btQSg
Z+A9CsEg4jgzjOcyVyXpjb+qAfkdhVl6nk9kuFh3iG5P7H3COkngr/VEIk5TMNtX
70Kk62hAFEC493FUoq5wLz2zgEMzHN9xB1XBAhjYxt9ejjsi1FXAIaTwYT1BRY4/
Srgj2oD3CX06f220z7ZwuYUHqrOgT+oP+liwwE5bAfqSwS/f2DsgUlkMRFo7l/rc
lv9F799mikfZ/bu59LP4hroTRI6OZsxQ6jdQGmyG3wYFrCyul4DYMmwzFvje9+Ks
+iRx6dBnzroBgMn672+wMnkn1MT1+/m19FOSxIr0N6t6osuR8I3IY3wQ5zo3axXV
WyXqOUx6m0bA/AGbz/3fuLH1bH5oa45yWQLLMm5KAz+hxiScY1raheCZOLXw80VM
ieE7nDx6eqvHxnci7/LDQskg4oBt6LMn5y/4XU9e0QmPFmdsPvBobudfStKEozsT
F98/K2ADNNakjdLwCYveSiWCtxQX7QopN4SBbIjO+wS6PXNSrgNuv4ZbVhSp1jyf
LpHaaubpYFNjWGd174ILptckwHHjQet5TPLYRVdlbpBadkZvnIOxTCo1OZrjbzOm
01KAEzRdgbC1frv7CNXKRusFpUGz+GC/L9BAjkzAQMTmkMoS2txmteSg5CeCISgs
08n2wqZgitsR7tyH3d/tMfgstygH0R9vNpRr1MLg4ERaYzpM64Qh4EKfBZpCsU8T
gkfCX5YyfRXvs/bjnc/p9MO+kBPPd4KcJI0bimYjx3Jky+7bF4x/kU6RuLgIh46L
/fXjomw3oQ+C0EzJeUuSV7GJojXJ/YB3/LwW5Ydl5yPfO/gvTlrYc1xAYK0mxnn1
Y+Kg4DNUfqSIZcOhPVk/9iZi/CWeXskejqs9AizMAqqmYJUUKXz6DyBDAW6dc04u
BJS3PuZLnm5hpNN4+0oq56Mp2FhZwP+cP1in7g2zUqgPlHHXiByR7f8PPRZu4Osi
InIvwU6l/BWgfh0+H3/q4WfBdPGn/flasQjpexWOgWBUUHzTGYmAbRj5HFWVu9BR
rMJFhbCft5rAVOJz+6+C2GtPpO0pHO4VYk4u+/AsA4iH8IdnHWAqZP8A1C1aPMNK
88h7RKgZMPvS+7sUdAwwZ/v6z1hZOVf8zNmCxbvOMwHAaQ841LAVbgAGUpMRb3Ac
7L7bPFqPCkOfwYawLlqGjlv7P0fk4nxt2qXwjGQeMYJs1G5pU9eq7CIfBZXIuTwF
WhHkD59r8Naldfgj472P1vb6oqwIWBq9bcUs8Cv7hkCjJldCXdqW41Ie9eSO2xgk
AW5c8ORCx3tetSI58+ScTYiA/o5Y8oYdkQfEODQMy+Y81C6oU4I7S5jZ+EZBmX5Q
j3mdHsnIoAfL2IYBsfMBGxDcX9Ert9pFXdAx3Df000EgkpVM/FACse/ACsPRP8Kv
nfkkkgDhAL8t03wzwbUmT7p4jHpnopc7ZvPWA7dEIuoRrKy1d4paoPh/CXp1IwOt
M46cgSNSNESROwtz4Lbdz03rhrE7MUM0RdkRDEYwP0rO52rVd8+rl2RSYj3dSqx9
+RaywMC8HurW1zp8RXrzSzJKy/gvS8M8vAIVyZxl2ySaSMAyWw8Jd1v0nMO3O/n0
Mu8NUOK98+rw93uhSvtlz4/5kfn6lKpcbyq6F69Nc9ovhZ/CM1P8lQGVUgj7rwoR
ckP7NtNAJjVHRY/uO7JrVobJz8cwCcYphxSlEgvjzJcnhGPrWojliuzm17UzGH7n
NColWpZQ4EidTfYbt/OIMYMi+1gSGYMPTSvm8i46svXWNGqXqLQLHFJqrEy5SPiN
EN0J7wFjo4Fr/LviGS0TXlIqiSchbXOLDg0odkCcK5iliZGn91J09/fOjBfBoY/c
Bv0uVapR1h9hpY5L0onGpm4TRlafkX35QMWzgW8Fv5U64iCcoLHtR2hE0PiOj3C2
sW8TeCQ+TdD7t9LMG/It5bt9et9b/qJ7ZUIxxP4/IEp0uyL8qfFwCBdkLo9oJQdm
vTzFQhTgxQGRJ9w1kVTFWvs7T6dY+nrtGp2a3wK1+gYptN1/TI5lOw1oE1wuWNg2
v5ButNuGJsNT9XKCaPsHHe+A//fXpkxvLev/1MvWXt8KgYcc7NT5fx9G+dYxseOZ
BhNYymtWkpUo42cCOVl9bUxH7kKNjG0+qB8OgU0rR7nXDNXBcWcNiuODlP1MihuS
LqJRYu4zNATsQVzrd+s92TpOqYmDID/vOH1gDYI7c3s2x/vyximCk3JQ5ChvPsbp
Yjxzs8u7Z3DwYEls64h+p4eGt+ClSJqcUC4eHwPxh1SRcJFxLAiVLcBumw+0YsHB
OH9nw5f/UPsPHOW3cENUs+6QPlhaYos47fCVE0MqjsNAY5TTcOI3qsilGgr+K0pd
lJbFOA+B8TDEvO4RjV08/QSeg3+QYuo+j8O5dz3rX6ija9K799CWYzmTJ4CUG+Vv
cJducqpVbB5vhC4dsSfApNMAIuXWwCh3S6lCiFOXhEJlMdeg/fx+qFv/mb4udUHt
a6cZh5Hb8hU8eU98hlZn7qyhdvbLxNQUvbiHwAQCdbiXLizTYTEDCy1norweWC8Z
Qq3+iaT07PO3Rvysth9iBbOSfjVQJwp0t1Hrc2qZBOqsucLi5hP40JGB5sGbxeEq
7IazPwwsE0eFZWOfjhDHXy1Cp35euiue/m9e/Q4Wqcbgs6ik7wrBhneINQjm/2A6
o8KCSS2NaS8KVQfRNMHweGCkz69sopx37DVdbYjsW61okY0NuJBOExw5A8Fh22bO
zWcytaSD82smaAdinIExn4PVZmNFM+JIquqJo0vR4z48j+lI7YDOBF8M1yLQHTx/
d/0a7GG+sVyWoEhk6SXuppaGhmxZTb6+Kzr+BZNeIL4uebFw7361p5rU5Kc+CTln
LFyONbgzR/vfvSTOoSL8HmhtKOjRU8lvkE9PzjUegyTJWp0/80Isc/poOCbAc3Nq
IvlTVip1Zs/5gw9Z3gquKaObfbNp9MSUD3DKhu5OMDsVSVjdTEAhCti5cALQc6sJ
CkqDJHcjbSypwr/hZDtuqYx5DzhuZ6tKx24UXwR+OltslXllO4MFA0E+qbPV+/W2
koJ8Ayfd/C40uBYxEWgNDqTwS6tTD+9wEYXNafsKKStn/DSNVTI2mnz13QyUPumX
w5snDk3jJERZ3fKpSHmgHE7BTZ/hMPBPYfRmJeo64cxTWSFAYP8yxi1mjeDN4tWM
b125laB7u8vTYxM9g+m4/Cf1YZmqPtc8TExmS4lpxVDzolHUP7WC01kMAbN7f/0j
ByUEkCAGqWTlKlXzSgFNXJgHwYKFpf5Pe2dTukYJ/Pc204M0CTf5645ZUNhgYQKl
0e/71+TksZvgltzJKSrpLFGamROtbYdp3mPZhED0qaqmS/ZYD38aUULGpMBLITwx
1rBpF5YfJaDZ1vop5qMMgRgPlielUgDt5VH9tVcCfTmZVz+MPO0ByYOJEI/KS0hb
x/T5XsearuCpAlklsX93Uy48seT0jSXPXol1E7zuh3pCALI7MMHHV47i8H87c0Cv
NWspZFk157ETatffdDc+beBD3z6ZUKNx9orpYSNWTvBUfwHLw9t1U75Odd/TT6LE
6JRPULP07WG1pQb0eCx0uKkRQRfat/qdyMBh8zBMjlbIApfKXfbI3luWhKSEaTbE
JJd7W0Fjx6XGyifE9WDIe/icPQcFGU9+65/4t1mMs3oGW1QvCFjR5MFzMZ4uW48v
mx+LUA5LE1S7TAAhTw/D2E/FwSNhmrLegzIbev0b7zT4aZJbcYFVcLdrYsDMascg
NYLAxtCp+mKd6bHLpQPiSjSY9EFUPH6JnhA74PeKjHXzZZuV56sEhwu9AtqiJuQk
izIdX3tGWIQRvF5RXHSsqbaV7u423w/ZsRt3FDNyRVAvtvCYTOM+4KOp8V2u2YTw
A7sZ6gQZUSg8EwblLIuR3QoeK3RrpJaV0HYLArISRXvcKk7o0v4tuIdTYnPuSMB2
Z7aCsMmkFlXGgNvx8js2BQvMzMo3Iorc3B9Z3qlZD3fSeNFkS1bGwrcBVNz7AXGO
baLDPBW102bFzQqrUaGl74A2gjv3v9A8Q9+Bad0ckWxb4gRCFmaTE6he6V433KZp
FDpqSgmZ6zlFCYe6jflChRTTuBNsdpUI7QN2D54b2kY4wsRx4EtTDuWeljyuTCj6
iTgAQsQ0CwoW9CfFyX3A8dKSa+oWZgUFqtgCAruIs8wevXMHXa43MCTHbUgtrfUK
LuYfhKverHonv4eZi61K1lviOF1piOr72594fRB0ZO9u+uoOoVhJzCGIhJi4hnEY
NfdAVX3xgw+8HFd1kre21M+Lf/liHE1lFUvq7uECSmLuCLR97A5GVFSEOmCq/EFR
gVm6xQTGqKIN1TiJE1aw3RJnb6N0b5ay5sswAtHwUSZpPMK7kqdEBOTbm23LCTZr
+1FzSGf5uCT3mdkluC+0ZUqYazt4m/wt1ERVUGmwO+EeaUMjIpcBp5s59t8TCb3E
2wZxvQYr3bxUCK6NygmLnzPMkRLMKD+ZpomCgCRqYvII7Vc0XGcuYWwinJ5QphkV
gf+36RZXhN9wgk2d6XKBH38zDk7I7vx6WQ28oMmWOyt6GN+KSsm/4OLJSRu5qGQf
1PtVhA5drMHJvvoCrJqDjjgHqfyHZP5T6tMGsTwPPu6RaPbd+MqBWHUI1q7WsyFK
C5lYEI6SgK2TmgPUF1YOoV8vpSeGNmSv5IajwZnKMfn5nhKi9dnlgiORUka437+8
WOz7/zJhFpgrb7hLX1Fsoqf6BLSgRC0tRCaemVe6vS/DjVfkGVlJtO9ZcaUzNtY7
IV0mv3uolJKbdALowoLSoOEM+on//CfN+mUZFbW6g/XGGSDOGVKJjLiQ6Sx94YFr
dfblcg96EfJlruWtD3BCHDwcHMnMr4XP/CIGZK8HR7IIZKHaJTXrF+At1zMhIcsK
0BRMjW1pX+iZKh/MeZxG3VN+IZH6RKyKavTjMLEFpB//wbfMKvHU7BfFmvrMY7fq
T3uRt01IAQblHCzTFhOonRSX8D7SoMvBWZqdhvrT5ZC4Q5XDDw2FWLF16FWfVcWG
FUzHFAXj7w9MlpFoiOCWness9aYm11hu28rdvLcwi6OtyocbFhG5NQZqybq9e04R
/bdRO1py20rEwAlB5k+m5fD2WaI6k1mqcM1xmPyvvlE9dlSvUZGPcH9gu+70W16H
kHDk5G0QeBFn5kWD1I++4cbMtF6MvR9Ffu/F5Yz3lzRp1scEe96WzutbqIMrTUGk
GdjPUr+HkwDVTXuVJTiZpyVcC1uJxU/ya0B52peEmDXJVTp4c5HGBiKYLPWzQ+2q
rIkENrb0H50GZtYbJb7NqDo8Xq0LyB82Fgc4HQwHZMHc3CvmR6kBZjiTanEUW+9B
r8AKdibnPiUNfzcrS6pLoQsZXfN2m4VBL5SzBnKIoBNbDgNKO3LpMCeWQfV4bJZq
mBAbyHrOmeXa5HXBm8eyGBeUkxHyQr0/xDECTrafbrm6n/uvu2209aebZ/zz51hj
6++17kWLen6NZ++oOXFyo+jbHDNMMdPYuPkZCL4DQno7MgnrTeqRN6OkP86Iitcv
a9Z1gnofo7XQEnQtvItGbxv4Meu5tCFAbLRI3Mj6lAMNkMNTJqYYN6PgL8atIifp
ssK2sI7Yr1fX/HnXDnK52o21qBjGIZb6kvIq3zFZ0ZrSVgjr97ct33FR8jtoxoc8
H0SW/+z7GpMsLur/9U9jW8xGiNruNk+503iTIySZWSzsTLjtB5ZclIAXjssEr12x
SZfdaDURyJWfiqkDnmx3tCK79oRBD1b/oOEFNRlNWFd3mF2fWrj4KJZo2wAU2Tjm
wtenYy9bWeGUc3eI/y00wAJAgyWvK5CgCx68k+yv8L0+42yULy0xgAyun5Z6TgYv
9be8/L6baxt1NrZ9aHO4p61VX9Lj4QEf1vrrPZ8fsZ+KBra8S4MhBQuSEj28tDvP
+++XCibZD8vIA+ytcTaXy6NyL5cdbuWvryVxcGorQc56QiUk4SJKO6J0YJgXDgYv
wHg6UemIklLKWWwV/Ye+YOTdcQYU+tKyyFBsd5oXUCqdf7fiOX5EEsaQgAjmBs5O
DihJ34/QhE3IjQnnzp6UR2jwFC4v1tv/DzHqnsEQI63S3RwvGEKUeYJlJEwixmtq
Ove+mD8HiyzZclNEoHrrF3CeOhqYOfaEszhsMzYzG9dcTFzFODbWjjtJJEiQG6SL
ZURLC/jcqElR6NHFb9Ewq2+RffSBzd5feXaTJVds1d683LVKfeFIbo3A3vWhkucY
zjOezx25nkijqBmv1N69VP+QZJr+bi0p80+VJ3o3C4TPiPSxkEGbEqMNE1cME385
7oHzjXb11CkQkoNTpKerHTENVqF+8VMf1uPtgRR7brF/YFdi/CXgAXQEcRmqZYha
LY6g4rge5dztxYx27vrOoehp9MuTVhIvnhjbsfgitg8Oa3evuli/zwg/fhUQhQzv
oeLsARjP4nv6dr4EDvLScLnrdS2XWxDyydvFvScjKPgSnbZb9/6wNkEc3+lrmc+L
Li2t/S8s0sj1iR0CbwbOgWJ93ftXHj5AwMsNPX0fAwvL6i7uM8ayNZ6EhadH54xf
CzlsYlWgZGwWT6tmnPRC2C8uzIqvE/vfi8/oT5zqfIQblCWkA10cyp3F+Nx5LgCB
0XgKCNa78iJ4/WW86+JR4Gk0FoCu3ZuUuoBsqxmFCS8VFhJHxQs5LSgcoQhV6MwT
sg7gDxM4n9S3sYEJ5CQgdoCXKfGb0s+ButBdIpneeAdfWc6rwwZMC1Vp8B78TIUd
F53yvNJLEDb//AQLDXaLf6ZCvsq7jWRC12RghxJaK/8OU953vjOmtfpLK9tn8Ywg
BVsTsm0EdfELOSVhT+fzi1nuAY6L1t4oH0AeMFE2cLN9R2yUjwt7CNJ91f432hRH
jF7do3+IXz8Pxwpy1wsOcnrCiArkToZVp18tsr45e1Cfv6rgBTvfjCMnsoh1JN19
skL+RbGfVf1I05w6mA7+SfbOSGcFaNHyuRzinQSaZF0eXjfdss5MtQGuWmCvuED8
fFwB/4U3wVD+rytLkUQ1I1GKRMhXdRsGTMPevZCKG126RvC80SursDEzCZMl/y9j
CfyHGUOy5niLdgs2zYfhIClDtkBYstMBC2WLcl7ITwqaaNAWEikteb1pmqgHrtNE
5TcvwfWskAgNUiqNPAO7I5ftFNp+iMc+cYfPzAOhU1HyNmSgAMDDRb+6rGweFBcz
amozdA4yrx0DFAevSKD/r97I2PB5wAH6ikqC7h+HFMzhdB79mHgXnSa8vnCbzcDV
f2E8KN9QhHewZGswofz+auOZTkDIpU1ujmFJMJlhA4i9ud8X7OeWEmZiYrNX4UVy
6/ASDKVVnqjq4KOurrZOyaWDANW5HQXf8gi2knkTeR2ql6fDHcaAVtXfwLA3H+DN
5htWr/Ap+i4h201qnKhcCK4+aIfZ5nwIu0F8nCYTH9RCF02UvbGujWP/1pvtxJnM
mEGzySgDEudwMecq7nWne0Z5+1QDhhsyCyti+J4rUC3xToIC2u25FC1zLvb76CzI
tzEekWnEQGXB0//VJOZaKJnRRI/l3qJcZxlumbWRfZa8gurAv04omdM+m72pWJQ8
z/XhRzflHQrxpx7ysX5IBot8tD863DtrtFIBwo9to4q+D6g/TOIPunRdWcnmr28M
YnZBTw7Kluyc2cxUQwXCuXHzXTRHFiTkLwJjSWppmQZYQwtKqyCHQVb1F+DfG49o
28M/OTfv2fd9HJmSi+Jqn3v9OLLWTEV2D0aqfqna4ji1QYJ6G8TAoWl7YoU8KAqO
brsIIMVhsPv4Iq0JS1A+GpU1z8k56kNlQ20KT5rdu13PY7fXVebp09J+5kFD5+As
TFo1l6YfaO5Pvt5xKKUTgKl0+ahA+X6mn468UWI4f/1cx5PVLtCZHvX3JRJmk/RL
C0VcQ79mbm5F9gLMpbdYcINUWZyaoctXxphtHGv//5ypxqM8puFCClAww/9ce4MQ
Z4CJ7iaByA/y5zE+YWDr9FHa3S1zQH5II7nVzzKZhYSwXIFGlE5t74mV99xJN7U9
JKTJSZaiGjnF772woFQy2eloy3nW0YOu/bDqx7V4eHvXbeDHoe5P+nJ14yRKCBNW
yWrFigrVMTcC5xyPU+ULM9oUuyToTMLh1disXVuBhfdQUd+u89ltYWauktBm7sF2
+58VhulyskWc25xdPUuo2NkOWI/o3IQqnoh58hpF9NAK10LSs75YbxkGc1D8iwJ1
5CX8hhaU8vs21Nlp/4GutNxWQqy47Dwt+ue/Ds+Wba74/wN7KgbztQcwh81nXmcA
Lm+abGkVC+NlpZcFuXyNg8+dgRkTfygNrwi4K9lWoZ164M2yk3CfV/h37t2rw2r/
WTU1rI9E1aOz67SlaSKrpFCzkToCacGs3PtCOog2qyRA/VWOA+kv0A6zE9Nj/9my
y50Rx4QI8CdG78ZmT/PkDHG4MX9qreyPoPRb9MkofuWMbu59CS5bEbGQ8H9LIgL1
6dDOLb9rqosf8Wr6F+BHPLtYFCyTf55s5ZHIJdnPvdUNB5E9sYqF7FptS4IZxTp2
M6DisvzI1oBmoDdfJx579EYkIHTyOVomr5Wlnr3dHzOS0gbGiLMCF6b+xXCrLKLg
2LUW+yuHPFtsMt7qU3lynOAw2EfNxvGER1cLb7HxGozQ8UrkHstVoBAgmnI7TVjZ
+BgV4cI3F8qSfms0MzOynVUyb6p3m/ErwAEzUCnfEHELFUHZjO+JzBl7dvPjII1Y
30u2Rnc+Z5lqnb2HSeKAHI4Tg0L65eaJLzcNPp+OjuOhe7V/J24lnNuTstvme1bP
7EgxAMvahjkn3TM2wPGXWgducfy/nziLk5yW3dnCaVs6tXLP6p5Kanf7ggkjrEN/
fzRy+EHGPie41ORvPceUVH8giiVQvyJhQANWMEMGsLXbvT2eAGOk1/Dee218wpuR
IJc699kjYeoF0I/96QDYtN+vrT4mg0bcKpSFIXNlWPv2nRBVOfcVc44LF1HPBBfu
bwgXeFy9fWIbEqRI/obYzYSa/Fko3MM56ZljGkJ1jpIb5lOqOez6B5wFco8Mt42A
w5jDFzIjGK97EebMQDdE6j2lMe7sXcdN7VLEJqu/B9YKwzFp7Fu+hBKrkyCkZlrb
/4cDvGQ9P4+dkE5j/RHBu+9EAo6my84BWHOThApBqa9twKlsmnNryvMmXE5kDOzf
3qltxousVWwyjIk8piVUovTnCZRGLrldzvrTHmzj+0L7pAIFeTXpUYAkSiJJlX9Q
milBHJjhUVlWzzhhhwRt75W3PmOKFBJq1FKeXIjwlYV7Hc/Mj0jU0QTHy7L649+m
j6EMc5IMF8TvmBuU1BgC9v8mpkHf6ioDvc18cUXRRhADPjPHk7LO+eYcDlzusI08
dF1ppx563VISqdVgz1bSb2viQWs/GrAoJGeJyGJKaYLs5SK21+NP7dqlYH4EIEQO
/0KQ7qEpbsLU5pJgh5+yubTEKCbt+dkTk+oMdk7/W2/17yGFo14SeW4EmCC+EYFg
FegyzrRFZ7SFa849D3ZZphG5ww8rJBEJGm6Vw95/AF741QVR9VOYEnfipYYHnG/e
PSAyztTljd1a5WYNcbPPgeFxSds3rleizLDJWixzceAq8J+J9kXaaOXS2RI8EBCW
cJ9xEDm9DXM361lTOFw/RXZOdZscegmbeML/wPWTY0NvL3Os/h9ExleGEaVYdTQC
QVt2vu9btHN/bA546iuwSh/7F3yRjY3g7RrAeIfiqoyK3kpzvaY7CKDF8v30zR4p
wdpOwOcttd98JnFMWwv+jlZJU2ZDRPHDem9kBPpscuIYM2MBpPDMmobEFJuuH7SO
3tv3/NuER9c+SvQrcG8PN2lkYKfJS5lyOtcEtuKykZmCs/rnl9BD6uju7+pGe51z
N2i83AkMfXvLFtYGcKEBFFZqYaZjRN4X0t8aT/1OHrcu8q4dxuZh+v6HVrp5bCOv
tlpWdCRTQSwHW/oJglcgMzrmzUJhgbtIbGurwWXRyhN3jJ2QcO7Wp6hgW8njVCEc
mKbaWGYdDX61TtSq1Ne4rmUIZmAycAteKQWG7kpmupBypM/sQuAS98QG36ixj8oG
GQsBt6bunyORnlJDJWmFu2tCf+d2769EnXaZnTDJNjuSSUaINm8hjKrtv8pIUoe1
QrTMFh6wlJgQFnPXC1rK0nHlVHidVRKk5nqSNXBQQXQGhn/D7WtfvYEhub6JR3cS
yWt7OLUoBKEW4mmgoxyxmbl0y0IOGXK5pv1RU0NWoy0JayjClizT2KlGriCzWM+J
qH/8rBVp6wGPyEtuHLFYXWhtGIpYvk/rFEGo5sDXtIGbrE9vWxMiS1nFXMcbQHS9
HJQvefi67OpzIyMMafIeQ5U4+DUUpAl/GGKa7c171lUeAmnDyia8B9X/NUlz37oY
p5K6882SiPU27YdT96ggufl94MRWZZmauZznQp83/5oNIOLhMt2IoaF9UwTYvozH
IzPm+2841G2swF5Gm21uOoiL6wsEGO5BKW+Bdi5c50HaroiyDhuoxoiAktS5Fs/y
oTWLdvVT4NQqMo0Wb9Ym5POTJ20FTQSEIM1vX09HpqV1lOKO3GSwPFWDq3UP++75
gSdKxgNVTs3QblNRbApCtvM5QiIunKtOlQo6Pp5FoIwJVQyLuGTQINbXCuQyM7h+
b9AV1mGFgwsmQ4dXLLw+lfznFlxjR5fJHRwCtMkOIIoTdozsg1nQgt9NYDOpET6O
gbuIWNmjnwzQJiOUszsthNG52n0J3PSR7pAt/GldrGRT2E0H1s6/EqFEiVmY0h5j
TUYf54n1a2FdSDreLvCLZk8SpsZM9x52VkadMCgizEzCrZc/kz7cwti0tU/QOG8B
a8GgIXiBFWPluduOyllp22qwA0y0tIhySlKO1VNjeQtfIdwjVva5Wi2NbpflyNRl
4VVuk9sR0MnMpOI+vkVsKwzV7kE73kyByEsMaeFoZb+xhfz6R3BOK5/MEvEbSBJt
0mwsA+oA/oakpBcTHlpI4i2D8Bv6snmjKVLGodbnuP0jI+qwNQVI5sooB2rZDF1d
Tm35SM+0B6/4BAYKeMwIYf0Bl22CSVYSOvmGQUKAGDPu5OM6hrmZxua89bo/jWrv
VRFFISHskg3xJnMd232F8sVpmeZciWGEdtTj8UIJPzsdY5BDmHgGMZQ2W07h4+JO
Yf2hbCeCa/8LKNKAx8mlheZFRjaDVkueoQ2O9y/mJX/s0vUK7AVd67VV01zoWSuo
Qva+qLPWI+7i7CDbS4f7nTR1I8RICHwH+aaV7UP8cJWWaO8JW5js/iazqNGZRn1U
JtIq+SiAJ9GNVpAwTn6m7+j9kJH0epRCwKll9Pj9lVzS2J/gdhbFFqDLaC0USzph
t0PywnkOnc8kZO0F5RWfAH9JU7f424rwbHrA7tuc6BktJT+jdTxEmphzs6i5hgpK
w+OG+IwJCeScASYoUgAZq7b5Ur7xxNG95v0JhcQVyd9ZkSP/O09ZbDeHwsHsLbOP
hr9g6ow2X/ZoTW4JX4Ka09GzfMKezdghVUZAxXQygMvHd5bY9u3mZE+nSGD0iCHm
YcC4jj7HviRnd99SJVEyuVRG4CqbQpiqLsv4t9/iYjKNClypbUkCGtfv0ZEYenEM
dGxihgmD0X2QFKgj5HY4vBaM2tqFduwPKbA5MhCCSsrvFPvZaIoZ+s2O5nkZZKTY
+tXJQALv5lAEhQtgWDnhKkiUPJuEeFQJF/rrKa9UtEvrx+aHdrqNythYgZYrm2kJ
wFbgcoaJqWRlT7YkVtFjIRU0AE+cd10t/2GQSwjBzosSPo1/mPgukkzpwLPfbZIk
4/aDfY8Ks9tEnPPmxyyfYXWx9apgpinmDRXl6C4g+N4Q6iV6z6uIAfjiH1M6QWph
nNrvcKQXCaP2uCeS46bbGzLLBkC7eB3Owof6AAYFg14EWLDFov2CfzSvUC7gRDn2
sTFjlPZKpVhhkt7KJgjQBiD4pnvHs1vU6KmXBSXHS2S1rV3MEcLPUtbYxk+iOI7c
gR07Du5aknZs/MZFSumjiAkZLq8Tz5A0ODvjmustKSbtfFG5VOLdFKhjXfvm+FGW
xDelEyOAShLV2CO+V8z0gKEsIRFk6ytD3U9DYM5od939UrfhCCl7hQU72u+KekA8
yIHDCJqto6b1WIFdpLJlZTtQ13dLes1SUKUPMVExe/8mB/j9gqaJAHCKyskbzJA+
ZfYR2+fsjE32gaT4562QDNhFkm/+T4VWrHhEeKrlLaq4Naio2UEsfYu/c8feqsXT
mixul7bD1lrhcuHrjJ3b4gsYdt/c9XVKM53JJlCZJd4+3u++ttD3DLrYU6Yhtc3Y
JEji6HNBnR6OnVzEW0tbUo3PuV9QRQDUGVokiupucNyBGRwA/B1FxdBWQiyGiTgA
AowAyHG1XmNn1n/6qKZc/36K/+Qky5NRAfxRZolQcjCLLq7z/2L7OgjxaLmmvOdv
aczOrqIgVjs5dPH6it7TAqW6/SexL/2XvPHDP87aSRFXFAC+RUnDxfL4GAUQRerf
FvHd6CQL14RhdiYCe0EqqWKf+XyOUHusrQqCr2R5Hrs99GzyGSu+TGA+CS+Xn2oh
e4Ug17nDIkBAt+cf5Bu1hqpOVT+PmhrB08edX8jSd2D0kW4C3zW9fkS6oF0736A9
H1G9aw6Dt/AjxUteZFL6E6ZEgaecDCYIl8S6pD6F8gxvCMmSlJ64Q+nBT5JMrbCo
sewZXl+ETOq93pzQTn5NE/xiqRJkFpRilOwSyEePPT561aAj+yxJsT3F37JGNulC
EASO2acChe6cieLAEsZJXHkQVLu0GvYqlcgTH3w3HEK9R2fv4GfGiXZygSuaPVgD
+LwmQAVAIzNf9GFAEI9zZJSbIm5vJuh80G7LkHvX4Iukl0Ej0O6AQPXXrQ0cJ4St
/KpA7wR5C7ETbte02kGyicv5lLD1Y4Z/syKJqXwBVv82uv8MgJaAKelX2WBH9xM0
YRKqK6SV3dNk/wgd/FhZACqFl5LinveRpxSxArTBwLGbvR/UD9jceRrCCUP2LkAJ
vrUaPJDB1+qxO4IZPQ/XvDQZNLDCl6NuUWxHSDHKHbfgbubaB7fPWN/jpZdgVCAD
kXwmYXFmKUKUjxlwQUv4d/MNbo3Dv3teCEeuFrl4X6KwhFDSwF5nUSWRZ6WNp37X
RK3SzkFzFvrPLMSeLM7DSGYxcAq7u5JL+W0bBJYVB6fmQxCqXTEyNCO62U8k4CEf
pnosKCwo6wGqUO0GKr2TShA788Q9TwLtaMzIju8BWdTH7usLLsQv6iRP3eJDEY7f
bOq6tW6hbggz7nAE3nqjB0m0t0x6MMFCCOPOzzfNawKdWQlLGq/Ny1Xcltd6oXY8
nK6yXsjmhFEHKEx1aWV5B2RtOsEsYGjS53QJfaToIV/Dw6PVuDrRa5ZDjSJvApla
vAg7IAFFGiATbey7NhQOHXLchewZzxJOkigrgUSg+fmEEG5NrJxYlj67bXmlPhY2
QyKcs2Yt6tRGd8rQ1zwdwuqhy7IXwFh5Kt+8i8JlijVnY9JTpYXij90GbJwkMzYg
obarSymusdRMdNkTOKZ4ZBkY9cz/aH7140as/cVl4kvqoCFDtxsWuCICi4hSdFay
eKtTMYWRrsxcxA4v0hju34XWVWoDhJRviHlfZ83scSW80C25DH3dYwmRR3nAOtxk
p5WJLxXah75rK00h/D7MouHJWczSnpWA6aqrHdlIkSVdphNwj1TwGLH6okUA1wcr
niXo0LrUrX/RXkisGRylwukEdKh/a3IFkkh19/kJGL754Lw5kAtOA624iI0eHRQ8
Mu6X2l/L4hOCokCfhpWloaBxOUACaD4u6eKo8j4ezYT97Q2TV5XpAiNCg+54qwN9
5JAGQfMA1/CDYs+GBXNyFa+CyheF19PMZ0JVLsKn7k+fLJ3Q1wJ9/5hUzRf03aoU
NQmSZ7DNIwR7jAyz+1gQQgISviSvQRJKqXg3/OsuGqO+XJjixd6weThVZw+5xjnu
Kgdg6xMoHSlM+7UGQEVyZbbnTPjl6JdSMVBdJfoG/tc+CInL4LAex/W6Z7WDkkXU
3ykx5WNusbZBEqWE5iAVT4ndttdC9iqnCKWV0P+8crr/pW2KNSgngCZNn37e8dy3
a+1mobRjA8eO2MLD5qZFpAF7l94LtPBtBNqXri2HAK0srpsZz5FkLnYqxpWUEz9G
5VMA5oXFURXnGauhbZkG3OrmdHDdqC/mmpdUxg3GxUxC4O5Td9S0x8SuC4flnT7a
o698jDQnF7eG5TwyZtrBhtpVo/CF4p/vngmGrfE87ppNVkQxU8rnr83yulwpI/iZ
FcC9XGExR99nbCdXTsVUbxrHVEPxE85r/nNf2p3DgqPcFG7PRn8xMMxzrDirV0db
goYbKPbZ4l3UY9Mw4nqsFb+8Ur1DxnCUSv8SnQW4wEtzig39EVxlRHL63wPuhcSv
V0D6hOWbKHenY+oudKDKdaG3qBhpvOl+mt428rve7YJv5J+nk8BeHEbHNbdhIVL/
s9u337ElApF8I6HknW03EMJFyNDziiGMXYzZ+agp5Va/OT3C0vwuH1mPV+TrZja9
830xPG6veSKSlDZ8rtpG9Jr/s8wGA0aI2OAnntJ9om1Y2EvxmMtuyvs9O1NchPjE
impdaHtmfM8AVCwGtUTFGcHuf9KM4Htl+b5xHpAwgQZZLPsTvoJubfSxGz2MFBfX
IyeYTJy2xgff+VSoarEj9SwgXitW5VXN/juLv89r11gEcfNsO0nELa6EJILmau7n
tu1IXT1BIuTNFsb8szuBHQ+eh2hOHBzO3q5pgw7Scrd7SVmpVUqNaSpNe3mNQm/i
ez6KoN8nqyQf/9IIRikudCDIltgn4HA4I8H2W2Qm8jtmu3jVfDb3KP1hJtFrkZIB
y1KuJtMXnFQ6KMXscdt+vlkDlZ3Dern1k0YspSbx+3j5YaEWsggr0V+NATvwXuKK
F3ZhjPKjB2EFLqcgYEXYyrTHxrPnsw+rZAbqms4kRbaec7BgiG47T2ZIKTMMQymX
JqF29y/Mh+7pcsZXCGRA3BUnjY7zfdchfkfmhmd8kKoDj97PJfELOxDtxISHv8om
igTojiR5k78DuwfnPmgSORDUKVwGDmptyN12Z+mP99nquI6oC42jk7EoLqvaBw4M
/3CjFV+0JLNwBWMiDTsUKVEel7lry5aHdhcNmkIdsT8/Vh+8Tji7VsGau09NwCY/
3pCYf7SaDpJp/SKZxvL/NrcRmTlrZ3i8s4U3P/R94AncpoZnMTVG2ZW21eMStHA7
i72JWTtRN1SprdyOhp4je1HmpBqTXDMwf2Gos6ePKFVFId3nvLIQ+bKZi/UDMV5g
EwLtytn7NM91unp4mBxA8lDL+ao1UBuOLCtHikIDSxWytMPDvDe7ZBIV/mmbRhuX
f+ybMrVba3FCGlyTYRKNz9mE4oaqkKLvEk2ukVQQwAoSY0XWAn26ZK/qLDE7gBYX
Rb40uAzuIBGkQfMbfMuInx3Q42vrBGkuZ5/5UV2tAuROa4ko8WnearTxNeGEvuJe
HqPGitULAiyIUE+f4f0qrvo4+KbvstJ9xpyj2Cg6dPDPcE/nOAjU2AqvoQvWbvCf
T8UpnZHQlgaNCfLHsdALoGENt7nmcXOkNcxIDSXtjlQyfbOv9lQ2FjySZdJmSsvn
OIFVti3EAMGvJQ2QqQtbZr7Ye6FTrkoJBTJMzT+4xCqDXLrgI9LGDWwmz3KRf4oP
l1E821CWWvCOyxFHfOFHNjxr1TYlUT93IClWAvDu/JeUmsX8cufuTjIN4hlzgXTG
ijxLV+Jlf0K/DaaJZKeWbIAZ9vZVIPZNPLDTTO6BHQxYD+7Z/WFmEQoY4kor+M+8
G35naeqcLkJSF5A+iSsYcvpcV+vqHMmyGWfjEd+27pUSULK50MvFD8IjlQEJAlXp
C3pGpov6t66HCI8GPzC5hos8X8J6wXXIvSjDc2p9w9X23klJHWWUpmqVeJ2NHorq
bSZL/lXxbewCMdzmtL510dLrLqtBGlcZ5RfSc/JF6PCzDGmwCzjjrKsk1LV7ssk1
mvA3M98CNrl8AkYFHqilPpq3OtxH1IVmewgZs9F63AmERuDiF3b4NMHcL2KA4lCU
v5e6r+UcGDaTWh/VrZbxZhzEDbJlXLlhnNArE9stzTd3etx/BlPxuGDZhXlvXUE6
sj/h0tlpBLn0OmbrjyNJ6M3xLj2xQZcwX/FwZiRhf01Hu7W9QNwJYHqnRemA3l4F
jJcmcg9dr+tTX4GCutR+nSJ4TVR9tYvfZhUpOCYAodkWubCu7pXo0o1oNNGIY3jD
Ibx5/KreJAHiF951sHXuqog175YJnkJd7OgFBb828CNxPpEzJ+f49qwbYWwltxlh
YoZSYeJ0OeTn6rnxUDKpOGI5ZbxBHt8aVixXdabNHTUJuZH69gN2gML4hRxFbEko
9RfADgTsOiAy7wK0F+Q8PEj2aWmt6TRP/hnzy8AiygmZaUqxQsXkc8n0Uz+FoIFk
U7IBezUbobOt9dHSOAVpyKjH7mzO0Bc+KBiiYs1PSNG7tvYa9LHfr+cseIMABSoI
SFmxjD1Mza4+Euja9CFD6hrNey/YA3thZjnT2mjMQr1MoXlLwcH5XX3lK9FLfSGK
pBU7Zse23s9NbbhVJ3tfwm4Q+BlOFFF2C6PEsb5QA/UHf40MCRsXmtQV3ak7ef6E
Dx4vIrbCXvSZyfIzKGp6OgiK21NWCNZ14ERGwYEfUj99qoKMy5OrnwVEuyAVeoYK
NdlJeQVULDSOAnhPT7pkB8ZWW42OhXex4rw0J+x0MbIU5TvK4RdfIzs2u+yHz7J8
iMsQydaHlITWUeck+MBU2Mw9NmpSpNWSLZRROxN7pm89HG7Ic9vkM3FbEycEHfHN
P5ZJi9xrK1kR4XHDZatHs7fu0jQe8b0R7IycR4wzWPi8hE7MGcyTr7+0BrB6mMD7
KIeZFoplaZNZIWUmhwR/bJeYffC/9lp6ZiYSnHB3cNIU1TGyEoAs7B84K5L4Paw+
cBCr0OPc/qbUsvUlilB9poyAdthJEiNRMWpVPKVLH2yXirWKAabWAraiwOtD2BwB
NO3+oE2ypKjsc+/wO5VISi7ilXoxi2jfQzvtygJkju2q6Ny0tX1W3EbSl/QkXiKU
gdHPxIps0phdWeC8ezObsPm36cCBDuF7DM20dWfsLY3P/cA5aZtv6xhMYGLUBcSi
PPX9QFLprlFw3zeXCGamDjk46GsLx8+GSKF5m91cynTJHcgUgANeaEBzE68HR+j9
Lg+CEv/UkkSSYLk3jPDjqVpNno5NmoWm95UB+7AO4gSztaWmlxHEHUs51e80ZLPK
KuMpnNR+vFCnWa2xPlR2FSCnIlmXx/Njjz3lEVKVgO2SdXOx6V80FbjVVR3wsZ0w
2Fa9ZTcMmQAjYaDxRMz02hmVwK5YG4RNUIg2UL36JRfc7Za62+0rr8mLXKw44GrG
svp/eKhCFHSOfx2d6CrRCFgk7YpYyvNPNVdgDcW/SvAihXOvi5d+DfSBtRQIH/BX
Z1wos+aNlD0PpY8OJFVRrsetIpcxT3nlHBlJBTyBBpExRaT+H2qPMTb4LqWP5rPN
GhGj9Rurz7WsQpC1YN+/dEwmla2PknF5aMpGaKr/eKPVSAMxumjuZnvU/U69+22h
ypTeNu0t7wDXYC6NXDk1BS2Qn92FDjn0P8kK2wuorlhRui7wLuO8HsTnzkiq9uzP
0SqhAz1nM4pxpHCEH0zMxyp6KhBTU3Ts+qfy+SCezjGBTmkWrsEL4pf+iCu33NjY
/d3G3vBS0e9dq6gAiK9CGTht43ptbAlbYqaAqVXBkscUzKnk+tbnYruO4J+RT/s+
GIqppyOLBYZyuxKsN8Wru48t8OVlYNCAbaUN7ku1trV8Z+3w1RUffkjS4iiZN3uV
txDZGxjsbEEhvozOAwoMt8CwkRMdi5m5oYNldZfl6syRbFsCyWP087/Ii0m7FhFi
QiLyhSZDiT+m/72ibreLwibqWk+cS3dvmQkU2Czgo4rmToEpAbEdFlVJLkUsLWI8
ZXPq7Mc0vhJu56pHEWfWWYjJ/xfzTU36vQ1HYsRTYIwLuS6P/AsOL3w2g04ps8Vw
cY43waZHltHLfAcDEHX2QO6MBgQaq8LZyhmKinMRVrAHGEHRw3zKidW572rct9ag
HVgjust5ntQ+pvdzpyC8I5NrKWWmuA/z5XNK2drjyIqbGPBC+onry/zO+dEHBHYP
plC09AIeZ0f/nC6BkHh9quh+jv85Wlp11cB65YACNXwyYySFPgvO+ltgJiHWriYc
w5bAn4UsM/NXbg2igfEf1rwFy3llnUmm6NcXs0w6+CBn50asSqSLCpro1hwXW6Nr
qAfxv2f9MMDjWvxCTKCthpuFzubANooZaf0XMeYXrEbTUrkYDVxD8f8f89yIh7DP
4+SsLuAE1b2M6Ka/RVl2xWBTkNXJvKLvftsPKgL2d9kPaXzYEICV3MHkPIoFAZVz
HGXiO1i1aYOjtbzQQbELUn/gmws4rlVqzt9/L+/4dCF/wiaiQN+TSEIqlVbgNijD
LvRajQauz1Edr7anmzjoq3dQr76p5F1P68r0DxIVUeuq8Bb20hjS1BG/Bk8KWfMR
8Ka4Q1WSnyHirjt0qFEspUhINHqJDG6eV8rFSjQXFDZmgABwj2Mt+AZhvJMrQ/WW
RowuAjqmVe0/UnpjlvnYW3hXlnfqF3q2pz3ku9Z6LzqRX3S8LU8zgSQ5MtEWbAGw
KF6ma0wTJoRiRx4dOy45uZecK5iA2Tl8j0AM3patYAhjUnjv+aNaGxcuaaHj/srC
zjBsqyQBdNBn+HBiNCqG3DzZHwLdMUvqdOZS6thnNVd0L7U1tJEojW7FgZh1mptf
VO483Znbx2JX/ktROpL1Ok91EsfS/bvAxVGItXccGu2b3Pen1UhD/uMdD5m1i8IN
z8RKlhfESOQKZr2XBgVAbmtqzoem/cjWVgMK9QxUDUsiQ/YR5G5jWWjW3LUhZIJ+
HOeLcUSInwzlk+G7zvthStGJuxaOWEoycFngmlMjamcwVZNyaLUSa9qgm5o6FZe7
NjK5ChKMhLwPDrt3yDTBuO3y6AN02ikh5vfu+Lxaf3kvaK4FbHHx4TPt4O/JTMsH
eLmtP4WA6sue4zMunP35BaqAijk+IpHHEwhupeSlkWR6LJxpK+Jm3eL6EpqgSvbY
0MRwRJ008hWnf+D57RNGqKDUMK7+w12lQ/hk/qlUK3IXuhmTVA8V4AwVVC4z5EWt
b0hl64cbEGmY6JxaeuWV/G/iNT4pOVUmTdJheMGOmaxz4BLZXcR74VW5E9FdAjxm
NjtLSDaxRV5jgX89GgjFcY5oCqFN1UumGS3SVHjuwxI4YxUwuOY7ig9bjmELe3LO
CxmNULX8CARV9L2D0Qqr1AOqHgDw+29UacZFGyXfAymOaMLeaoawtfwMI5ibbOAg
DBf60Gej2XYYrFAeqU+mB5gQ3B/z/tuoWUaJdU1p0TUfyDCXPUlJlRKVuY1NdpoS
OwWP2rl6BaHaQ9418JQyRyy32jnnwg011SsR6W/BdVR30yrMVgSWnuZF1nhxInKC
Rktjm37Mu5RsGPvb7JsgXB10iAvQn68C8mEYpULMSAkYReUf4oOTree1MNnnau3l
MQKSle2hEY9R5Ejx5EyM9O8Ww3r2GBpOMRbxzFxDUii8IcjMp7/+6hkpNGd3lm/L
f77Ky/I1Qj2lGwhPWJKRvk2tauhU3Caed8MxnlzI3HouGVbEoMTKewsrefigCgSa
SWTiKY5jX3gMBwBU7kyRZf2neuNAeTDIEK7r0OFbJQIfXgHm7nR84v68V0Oej3Nv
wjgeZ8QgC+a39nb3jBqxLXQj83i3wAY5deKbUXFVKDc7HVub81kNLn9KDromn5WX
OnF9EF/sf+sdwDmQLKx2UVAjcaI5MPlPkKM+3laL8CwQ25KnI0XCRmOZ6v58dQpG
ZdDWWiImnw1k5OJNRiFu11afkCr6jK9U/4u84uagOBDO2zOlYGcI2swq5vk1Ub1C
Xe19xwHiyj/2S0vuGMTks3b1WDNjJVZ/BiRRNfj7MHDfhMckyurYZX9qHFpn6tDM
chktR7DCFCJD5J7+SpB4CGOsSgjOZOVPaUmAHcRAYAfa9D7+G5Zi9osRXv4+/tu6
VCDc3RgoG6jV9uH1TRG9NjWwCS/4fJf4/BipFCrC4s62Hml9hknCPkMo/gSR0d78
kCiUZp4KnDL8ijGNPaR2JXIWoK8KEdVTgp5foKvfBsyYmJj1aZcqMY0GSo0XsV2R
HJIwOw3CRL2C2KVndzhW595U6+QmxXZwKAGxiPNju3U3atD9lZU92YP38bNnuicJ
SF/wlKgCiAXRAM7TLJFE91BwAeI1NL1vlw+y/337/VhZkERJdPXYJvKTlAvBOInO
dgQb06czqH2ohCK22j6an99LKoBOvo9Ce+mjoD3tLw7rI0xc4avHtzHrLidFff2S
gIIUrPNrzwzCeFJrpdkaYacMo2AVevGQR7gZQ1CuQcI7Ewcdbi3P5Q8CQi+ZULjA
15E3tO8mrXQfR6h69c3yEq8WaP5x8jp8Do4vE/oBolO72BCXrBdeMltK36/3zRqS
DHGOIu+FtDfY4MrAnduz0ApTR36rbmEv+o6Rigjm0oVLLPrVspdfVh+jtZvDZeUO
2MEK19ALebZ9TOuW7caR2NBJKM7f3JnC99zOKyimZR+HqggMsCLwKDvCSRyQ3Nlh
t6WUU9tgo4rmAkLhpk43ydi/+4tTU5UC8WSzQbMoS3Mjt5K57LozoiTVd7qmhhmL
FCVtJJ5slDoByO1Anoclc6azTjlmXtvY13XDJnO655/d4KTBm3+UprW45kIsjH4v
nL9ZvbSmu9RVPn847478LTeAVrwAsK90IYl3wD5t5+BM5WeMgFPYByQ7tNKBIJLN
M2Eill6FSvAlZVLyIfQfELUQmyqzjejs76Nfl1Y2pbjMYRhdXf0jejztFsRzSokn
EpIk51K0sFmJ4minN+dgtqTvOU5mN2wtZ4Q2KjsXzzyW/x/JSA/cUcgvsTQZLsY7
Z35P9ySTvbdRYpCjxQTH4xYxLhBuP5OUMDXMvm5xvpjoTkk2sWtaxGjxn0A+G1m4
M583xLwt0y1alUFCavKdXz11EIQZLa4NEHqcAPMmwmLOO/sInsLtAKT/HKNVOAoq
gqoj3u/H3q80PboqNqGke4K0Wpk4rMEZZjzrkJlJiz0SyQv3ULsJ3mlUUzgxkoer
rDLZua7A0JT2AvVyKCb+VHsVvLlOIz2XBk9b/vkuH77+Ykeel7lehR1fMQR3uPnr
+CRiksZL/Tq6vy7UbA5HONEtV0vt8q8CQ26YqMa4UTMlp5XyjDpuTtqfHxdkSPZh
/y3sO6bsKDT20nCbLHSlAfG8WAEndUudlRiYNyvLqHUqaeMZuRUUXQWi84xVfFv6
ldEO52eN6fJ5I2p4pLCcol34tAa2jCg5VovsV2btWMC+tW0UDKAjbEPoQwUJlYCM
du8e4ELzfT4tq09e4y9P9uFuK/n+8LkC+DN6Sld+uJ9ygY5+fBzuvq7fAFCGs8og
01JwqPxvzcMSB7SIPeLwL5yzWtPctdNIKC3gEVEuqDCvE7jMo88rmKO2Ko+XEMRb
cxXS5v8azcbPqNDdeVeRYodISzum6uXz7IpsQWjaPdBqLxD4sYVhBHVlNNOiwGwk
BfevzVrHwAOpiAhAz3Np3+JyTW9TeCkdLHvCCKPDEH0+AlzahKTzt3KgGgTfh4cn
IFcd9L5YH6PBiBHWP/WV6SJEqBMniwaB21goZEtkLbEWjUaZTIL3nFXRQaff0wnp
awqdZ9YnshChFy+BdEgKuOi/4QQFTrM774Fq+e9ekBWi0HZMjuFLmQiVdmW6IKqh
ajd2VOMfpP7rUdxg4G0clBryU/udY2uM7ht1CnFUY69bIxC+exElk/8hJmqm/gAe
c9KrOmSxdf8XHY5iNWaAla56PEN56a7pL1xgKPsDi2N6ZFEpBh+RykbUi/O6g9Pp
nQFFHbo/2kgwWOqhXJYhOgDQndvOF4IuuSkQTKgDsQIOqhop3UAC08vcrZmOMZGA
EAWFtWxnwoy6f2NnVApBS22wjkuJjDopECH/WA0Oa2K8ekkUPFzNX1nrRTFaYh/Y
c+6xObGy6+ytwWzybINsSjMn7ROlvQsSMd21l6Wo4gNY7mO2YSFLvpReGPgWd5CH
NRm8074Zvjd0t5TEgm6bC2v0iN2MrbPvfgR0RHWkPfii32tWW4Bs8+TpOZND7ZCU
NyIfMjdevrZNAPi5UuQ6QuxNWJEHPjBjt7ZCefoRXYjdXA1AY2rse8h2wfsyk9KB
qr8a5PJVnLxW07Vvq5w+TCevhXNqQxBKm9+YlwF2sBGkNetk9+NyhIMluuC9H87P
FxqzU4w/Cg+HniXsBTpOaEc9w0/Jpr1asKkzjY84bGtUukUgxW3LIM1/ll6mAUbK
/NmOQfnTep0xc52gq0da5Fry9mUabiQ3yWl8GPZKIoDqE9O6FDHiIoHixXfsG2pZ
hVGdpU6fGAeQpm6DfhkNNVKf1EkGC4vKdBm/HF2H8tPzV0ruu4lsMdZoDiZ1K+qF
Ivq4tZOY/7axaV+gn4DKY/UFk3DRnJ5F+hPGbFyiuzNHh6EAfRIzjVVXtPonyopp
7dSgLnxXm4i5LwEVRZYF+MSnuGZeTukcBOrLYKCUojGpWMqrWCN6TSKnkFPSEHkq
UXZ3pqQ4KFKqx0+SsOqEo2W/l2SKJnCg7vLId4JEyLnCu+LP0gmB7d3cKFJRB23j
lUf7NTZlKsCXF/1BP5BQsyU7qNmSUtitNV6MKhDBgzPobGvg3Jvjct8pwiZ3W4Dz
F4GPi+l3O+KJQPOIagYJuvV339bJg27z0Z53BZGcKhACSvHNCbHIiJICstk3pVBB
f75jcRMcKYftweBWPsCZbFJ9WQPQNGz/2L+AOnbM3yHL3Ne0DFWrNENaIyfKscX+
kS+G4pIkJTb4LLY/jdxmgXMlUC7jvMlPkHy8RUUO/EHXACUB0dXuErKUcEf8fOx4
ozml96rQs9y4y3iAv2RIEc0Pg+3J00iBWeFOyuKlaNsvpAIqsP9cHaxj77U2Ft/r
2XGhSJ01JE3cUtn9Z7aZJGekge7hbmGHLyCjvQ/gwaLbEPBJJdmF29N6SQc6GnE6
zQR00HpHnq5l6nryN0X35CQYptr/La/c8RxTY9TlDFZoBig91HbqIXS7mMVNVPHh
cRO4HYhbndI4jkvLW8Orp6fRWPbyh74tzVPETlHlzOh83R5pTTSfphjeJOzouRdh
4tYMnhJxBNd2g+eYPRdbagU740fCiCcYF7nGgYNXvcJX/DVzzKlnmh/UPhyKWngn
/ALRjyS6OvP9oee7kWmUo6xlv2/NqIu7t/ECOkFTKnnsC/hxh4jWzWnTu35uobIT
m4+87qGVSQZXUstqF6qoUKXVDrMn8xsbLrQl6fhXwl4mKqPY+KgrVElao23VBJc/
+sODpy9K5v5KKGDsLWhQdYz99Uf9bYAOxO94oKOBtG0pvWKZTTZD9iMTGZss9DjH
V3pMofGf9m4iSS/DwE2cENq3fagrFLnwYdwWDDZFNZ/jVoxnHDVPw2wiEtgmmUi0
bpMUavLXMrYl3U+Zai/3ZblpkPOg//3qotz1QZVLVnfTsU8iGn8kFW4+dqE4ItLH
KMRjPDrqxQKEEZy0uHWOqkYlcDgH1muE6qlPYgklOyMJgK6byTTaEt4w5zI7ni8o
tIIw5kG8FRufaVRSJXX6vQ3BHt4dF6NiNOjWhuCzvbQHedNh1WDGEHFv7diIoDaB
/r2fjh67NL+LpOsOJfkr9gQ/mFV5a3SGAslb7JUOrVYeBHaij0DHsleGGwAbH88M
Mtbzq6INyxv8etd+/LADYIxH4nHHo7TkxIgCeG3/gN5LxaGZM4TBXX6EV2N+PdDr
LcaHDVXO9Qw0A2SHrqVEGBSsP/ZE7sve6knNnv08nD9pQMfQaDCAy2l8iE6HOorG
te+bSkv2lrn6IhpACSDhL74M4uYb7/9JJVDd63kbj1oM+5yvvgNrsfNACvJfM55R
xngm6I3lLWpb1Vz8CcMY8IlxMzBIHOhFAS3SvJ6/gsSf/s+FSEocecZWVmSvc6vK
83zPE5AtFnVj3e4JwC38AfWL35hNWPK6O/FiKENgssIUjUr+3J1BFdMLrFNlS3Qh
FR67renrd9tNWT15oFEV7rvp7JeC5kL7kHxJ6S7JC1Z/IR9AFWTaxjz/Qxl11xSe
MiVAB8CkVcZhdlOC15AR1CvNx3KLQXdQI4OhfNhkz/9YhPNaEdG8eIEwUe8Xx9ZT
f5sIlW8vddoHAZCO1QPz0N68oTwvFUTZeP8X+HyuE6KqAA2lmC8ZjlH9/drZYQ7e
3YDFY0yYNBhZ8p/y7HGTn48TjR+xq2Yz9bvsRUSqDJ2Ad8ZJS7EDPgAlQDS2qPgr
/LUi9lIrNYfqTF/JOktDbDjuE5ePcBgZ13C4nXdF2/aa3ApFxDPJvxyzgATb1ohc
0HEvd7ZgyNw6T5KDkJdxAmz/XqQ17zZoLtIOPGcGs8AL1rrN1EyRURR5Jye7zllc
Ymm3y6CSCg10aWJLL9qGB5j5HLmafPZAxmQJINDmFXSCajFckWKC15klXhf9d5qM
TwgRMFdSiHRdCPytNQ/S3j74uJFNWOaOlmzvPe9gJxQBp1nIVKzlMG0oxMDm1LbH
xll5isFgoywURVj6Zn+iqRvV4R9OgXrWtDJsFTcKUixgGmVHinZxzlcVcnkWUNXq
Ww8F2jkEp0OBy6Z2y3k/C46E08e9tYtuNNUhwS/YPArkcYDStj2faCSUZ5LybTgf
EeEGqT4j5+IvIm9IDeHxNilBs3z49qKe7dNmqg1XYCzgeOKjJWwqCDgjczIGRe/t
Y9ao36GOE18OEHGHI7n+4F/KdoozUzli4Z7hZu4YDs8zbNed43xULYoswVf13zby
aDG0ceNtoBfMvmgp3kCEnSbuohGRHTwL8Ro1VD4qDfqilvyknUcOguEaruZmueqo
/hRsLqgziWaqxCkd6PuhpApDRBmplcYlPDer80vCq357BfFUEA6D248pM9cp2AnV
PAUL809v3VqP9oif7wtTFCu2lxiGOwTYSH5ULw/b8a4M3oE96py1ETiPvVe0ZAeK
m/r7tJEoh2MkJu9SdCDjK5Ug6Dyn6XhnPjyv8QVfMSGjUGgrXHrshGGHY6jNo4Zt
zEWn5Mhuo9m6+2tmGF8Oa5wqCJgll3HEpFUBCDrnApDyIJ6uSJ4/I/vFiIW9GH2b
MqSWCxMyhF2e2RDs0EOt6ak0XRBmw+BNlJzATv+bnMsctxH+zj7KcCghYzjChGCE
uCVO7il+ScZUKgBEENwvrEro2JcOE0mKH9etFHEmlXo6DU7zdMIKGRLZ9rLB707r
falzD+cjVUpajC6wxNhRmhgPBD6mkiA9snPdFaCUpDB07+EDv99OY0pIL4+GcvOj
wxMUud2mp7yyK3zmKKCzvw9GKKZtloXHpxwhZ/9OYrZGnHDB6K2ALs9PhGGPtClr
k3KZxIZzMG0w5AoiAN88Ris+7/GpNkAqjWa3qEHozE7ftKHS0IWqm5KYUcwGUDjk
UYpdZDWP4gdnhxvj2suyT7kQ5GZmA29xeAT4D7xPNv8bejdNmwU0lFgCwcP4yb+p
y5W4PAeX2adIgv69UAodCdZjA4ILM/4dWOgo1HGdPGA/y6/O1ODSImZwVmdw/tHy
RGrWR9Cf3Y2erdZbz7doHJGCcUSDpjgGK9iaUllsQBS1LdVwlZcvooxNMMrkDDog
voafB6YEdKDns8+MhrDTM+oS6VYn0s9KUdJjpDjQklkaZNXB5N/s/sPm76vpca7z
mPcB/RFECJFL3Zjr9h5697RCxQ/M+GnoV4OQXAW58f71I9k+mgGEA5Hg36mcTqDo
Nbu+cdyrUsCqGeHdYU1BzTp4dyDvsRA78UtObHKuM33S6nEqv3rG8OlO9clyIN6w
vKg13DkW/aWgOgy8iH2ix/vnlpHd5QfT5Kh7vC5pfADxnwQ4agzl5EEsfdc3AhdB
92n5tS74AYYCGKVK5fnkd+R/mdl3i0j8geIPTQCALTepHpIKwbOYTcqrvmwbgR0L
cwb5ndGC6Dlxtbc15lYpXOgeamp33+CPOS6ToZlj1FSFikZzPJ3zugKRFVubZXCI
mLGgnLq5h2uv+vXgtTRWh1SuxOOOLhPcw/CIQ1AZKW4vrNKf2KAOGNKaxVL2bDFj
VLijX8vs0MoTyyv+JI8scPnNNFHJ7jROr9QO/b5jgK2jE/49mehyA14iawjkAMJK
5Txctx7XaNmebgwyuC1KLs9+bZG7vxngDWXrWrs1rlrgSL5Ft7PSrEkWFrkXYFHe
7bYDTo5+BM5MFJfn3GMpKr4xjcpI0wm5YBOo7TAUPcUSy18uQRYPk/EfWWUDNCa+
92gYFbXJvxH3oLf4NGYqVAP/qGGwF7resgfvefA+ezRhcA9gFdiTedt602yUqDCf
obP8ijbqHPiWHBIIALQCHKxgfGjjoR/IwqZZ1uYntOWMWhT6nUAdvVJHnDubs6iB
ctwKiV85MaTnrwTSrbVBgdlS3LKOJIJHknpdl3shhPe7QhPgWo9qkWK5wZPn1B88
9EjrfjPfzqtuBSddalF5EzH2EI128uXYfwlZ6fbVtZJkrMGaXiFBFQJBp+rELz1E
picPvl/O0USomuWuFEflOZA8hVjnpWYJZLlyOnNi3PY1Fwm8tWIUn5hb2vb/UDJl
12ILs9+Yb59NlaDW43qMabP+AEvU7NWDO+ynREtcb59aW1u4VestibkbZlwDl913
1v6qyvFRYA57aGmWeO0i1rMv/XNBFa/DqeMEN2okHokRBXZdXN6gp9ycU7NiAkJc
OTQ6sWfEe9QGFnSlzyFQ10GnwG2CQgVzVfIntINZurYkvm1en5zw0fuWHNaAniAB
phFHzfzBVJ0CCei1wdDxj/gMWCqGoR3nLy5Q4kaNOxQ4MzlGwlvdf/ssuHvqEGvF
uBydZqUPFcHKwQt/5O09ppoklCnZxPCINXcPZqSEfaAsjw+L4PUQ7B7p3yhOEojt
ODfA9XbKaYsn4Y4HK7gFUgTSYnbP1jcLXMvoYiQlZkZW69S0zwONATHomF+QVqE1
g9DaKsYCxR0Sgs0rnyRuMC8dM0uP7taeCFqG0VJ0+ms01qimAnaGD4QXZESAbyF+
PnoiRsR5VJU6SYC5+gST3tx6fbyPLjEDfG3FhI2ThW/rKTMXou0LjCKQ0buhcrvf
ixn3nRaSrhG9XgPad5SkANLDtHkJhOYsl2SuNhmqz8gkO+whuy2vC1L/4voVjWHJ
AJ2WpYbi6YOQzwjKBbA1NnRecrHsJ3xHjy/BP8cWcb3UVfUTn5l59MtZvBskh6HC
47Oi8/3Dxpve3c//dUUgLyI/WyC5jcRt5eAamr/ZyCAdN4BQyc0LJta6XyeHIBOX
pzJQTkJCFV9t6vCASY/DLQ2spsG5n0SMLd+ex5HxOke/4ErTUmarGds+dQJcXxLs
1gJYHxnncdk36Eu2A6eQyZSjaATPO9kkBPnOWGYvUW6MvG9DwPT/+ZwRctwmg4tV
EycfCsyNLrKfeln0ai1I5L0p8ORFdYJrs1dMolmo/h5y609bOcnBfviJ0Aobk/Jj
No1KSJQlNMrFcn/vgCNlPJqXVfdfruRZ4UUEWR4nsdl7TN67dvhQLtofCmk3+MrH
SQ5eK5MlBwbhWDCcvO2HnoLPrbbK7mrMuzj7S8BWEIFLjpu1fcRwy0Q8TBZMHOxm
BqScclkbSJoHk/zckWf+tzXEd2df13SvCXcJ6ftG/8/+NVGXsCVW9NbBK1x5kJkx
kKeImN37kTDRIElBBASE2VR67oOZ+aDbMKBOlvoctT5E/9Y0X13Iqb4UkQphqWl4
NXuHMuzx2/ERV6qBksGT88XspTs2fpt4vlv5c27ioQsdhxm/iGlTB0e1GOF6oHbi
gbkmGBYSXSGIZqbK5mUetDGfdM8GgBQOEd3bcJ6BLrH0ZrUMGUrHS8+2pRVqo08J
EwJNRodnJGcNbxfYc5fiZ64g8mPeK2bIysK0Nn27afnxbwbeOlaPlZlEeXcZg1oE
ankmgtM7GhXh4SHlmZ+KEYpAJoFTPm4Xy1D1EnP56VKMAstvOwhNyjWVDd/V35lo
0s8XCAwuRCANd98DdBfrx7xu7We+Ju03ReL4aFzX6FF20IVl8sGOVd50Es0eHBxG
IHnYJrlNXXEo67TqfMx3P0Nq5YmREG80RzZaAY5Hq7QWSGVi7w1ZE/mXjytCBrge
S24o19fY59C6GmbrFvZgURPcGu/JxaK1TZR+3pkhZLn2CVThHMd64uqBdHRvYuow
UJKZbQ6R9sWJwW/jQ81Snfs+ZKqOQuw0CNvdErM0rUCg2kH7GfWEmgiq6T9djC5w
ChXM2LxrSuUlZIEHaGwujNQ3/aRVYmHdesakFiJrtwSJgFamrbVxZFhQj73QB4aZ
mN2EwT9rIHs8m2folUle49JG3SY2dDnTSNBdQhUTDNxvfJQFjUY4vjw6Hxj4cfZu
2D2DmR9ZLe+IOIczxPV1GWcI/IqJQsGrL3ky3BrmIahRYmf+RkmC+w+8QeX3uXc/
RnGQKxagsPHQY/uq+r66YcOMm+3aq02jWlTFoXO1mjcvv/l17VCzx0xNxWV67ipF
189FHye8pVfF1LCB0OcYVKh3cXQMM+fqNns2pcGDnyBy+GTg+/DhYFLdM4XhQWE9
a7A1MIneILexukLYN7Sh+Pw1knrll/3q67OTwa7kyApstA56zY13z13hEakUtOqV
RIcgQfog0tzb0VdCquhxXDmbfxbpfNAF44zbp6FgcP3PEVlnOGbaMQRWGWLfc7tK
RMedLjv67VhfSzONoKyooFLEeX18TqTf9hfmws+JrKfdKWJdSa5fPWFa8BsFoutW
YYyCEyhOvYJH6RmyND5VSXZVb5xNXRq04j4WtoAjZEVYRfoFG7AQdIU6ieofILx6
WYspN2/lG3qqdmsdxwDJQYRvcesI47GHBhc4EPNSGgzu0LjwX0vNzm0UZxggAwG9
SmrF3rn+3CsmE7DXY38yKlcVijvUrD0RlZHioM3KTZtL0gdXHwbRvRtcMuMGRpZE
y1JmyiARHSyDqesjq2vy3ZkDAycE2oXc8c5lU/k1+U7n9ezNRftm7arXffsyoTKs
3HPZBFkdteXLTZJZH4UrILo+/UUImw0xf0ANNL1WasEvgVvONwQ2LX8wSBFJuHkA
lPeS2tcG398ntZFnJcEO/uzNmL+mOqFA+xt0sGE3DzNMWlc5EP1RB5jCKIIF++vE
m7oCLZEtnYd5Wcg3iz12F5UXjEE5OwB2nO7makTCYKy0w+30BumRonwoqv+aW5aZ
gTaXjhUcRs2bgoryyBWm3aKot5u2J5ZlX1vdyWDfTWttSCxjW0k4jSPrGocqSjeI
ALHdYjxBEtTZUwzkiO3e4lcbsnGz2+aIrd4/+HAEZbKmfFySGvu+MADOaJq/1U/y
oXP1z6DnJiX73/Lm8ryURbCeRZA4kvmlQFWESxPWto2/2HVSaxmhR0ySUhh71+eY
i9GsLUEQBmwkWkoPhvJ3KBHbi1isnzEn4ULF+Kn0zfm+7h44jkgcjGxU+N7H7i3r
gJWX8Qy7ESjAbWsFTJgCxAk+kP2+j+XyN24UP85XrQY3d07yskn7dRXaZZslABJc
7XDCrciOzqBJREgcR03HGjaiMCrN/H+DBTdG/Cd8nO2XaKkz94dvjMwZbu+VSXeK
xHKZA45ptgBQ+xwXB0lNuvVHp//1Kw0sjD2RnRtJ5exhJMg6P038BZeAXRbDf4vl
isMhl/uyTbSGDWFHF12Imn75jqRTY3+9G0vYGNB//mWf6dzaY54Tg7FJXRPQeq4F
9qIYGbYkmptD4U4MgCcEIfgL7agsi0tEgxrdIKI7SCF9fd4LFEbd1XH5mYqzFuhL
9qut+/HXAMS0wWMcK3pnqk+7GGBxS0jWFTagYO7HkKVAMDk9h/2ua08YW3m5J2yz
bhDArj3+Zu72q050cQEHLqB6A4oKmSgi/8HQ8CU1sYdR5CVEWsYCI68QCHJAOdQr
P3hvtdqeOZl68BptsVzvVB1Gs6fcjePAz+ttdcXLi3Y1ZRSfoI3ye5dboCpCPK07
e7GQOEcx4D+M+2xbKiPRlxqyguD2M7JmktIe+A4GP9pkriTfBFhxu5FfCwHfy1Vd
kyK78FK3C9A4n4V6a41sOXr2gg57P/Cw4+tctQU/VV0GI9i9a5Ld/SZqtzig6USO
R4VHqYL8VbPU/AStbbatrTqoP2GwR++xSVinUJsZu5FeyfzCu2spAmclZDEWvETV
YasDsIUk9oZkgDTWI4TCO2IalK/s99AHnYwcCJyhwqVdt6mGZtuLLEmvxaMB7TYw
fT93C/D1Ppd89oEoLd7q0ti3a8fRk1y5f0EPAXTYuU4Kkxe6UODujs7ZgQD7ZKoN
HXbj6Yz5+lukP70atWm9P7BwBHCnCiwBtH9VsjNFGpGMuLC8xGyV7gKo6Rbw55s3
R9r/BJR3jCY3yg4NstcxAp/ONT/DLngBogGrLk0isDLOVa3osflN0HYO8xT7MlZw
ADyfzc1r+ewxo2/zZNmW1RyB0Rwps7N4dQDvGRr9oSwGNguggAW87Vr9YcQ46ufe
ERcxI6PFworztPnLWby5slnLDGTmcV1FKo1r5uTSTnkO18bJI8y6fNQtQZeROm5c
OmIm63j3F7oOrDzUkBtT1QztPUhaphO7wbyFTZwH6DzGHrUOkPbARGCXfJ3Hrujx
Wp2QuExOH8Qa/hQeZog7z7pj4N9dqVkDeQMGkDqmhS0I+PV6JytwaWP9dnm882pG
Irde1tWO+Smg6ESPFbITrZ6741BmUGC6Q5pU3ZxLpkKM23Dmz841fllAQgTiw51A
d2+597jBehmOrp6C7cz8/mSfNuxVQcpJesX++2Z5PjLuSbuK+OMO/FW+JagsNDJa
GH44KJ+mahH+25iTTDSUQvWhn4Jd0dyaHKf9cJsunwL0x1XfCu7RBU6aTsQwqOAO
k0mRONe0CYggNlbM7YWiwJtD9dlVDvvEAzgDDDK5z88RbER4kKPT6+oaPVzwfaWh
ZCe9VftBHO/BMllfwW9fW5Ao7SdkZSgB+10UBg2mrjYGSHT1O02bmonIiFaeO+aJ
+x5cWnU8zH+JsVZA82X7DsCTtiGZMia56eNsrxyehAViEbUD9lIcqXaHJZ6yMEB6
k+/eyOdqkZ1QUoE3CfFAYXuxGaHK3zfZLWxVb45busoIEJT2ke1Keae4XvHRvZiX
+UFYVkHm5EvZtr98s6c/L48KGmCXkmju+qT1XJ1TvwlcZKd+87r8zzoNb3gCigJG
hiiNQnzBxAH9NlaVHqbSWZqjaBsHTVkakmWIr3Qf7tqkVciXmRfex90aM6gb8uWs
H3sU1kY/bw2ccsWfo/Cbr3W3TVN0LdbZzYNO6/UTFI9XeyqI5BACcs+aUqC/MbAd
9gWYTJ+b2LkZE1BONctD3S6bIKP9KojdREMXjOhhX7i5TeOOcrIMXdWrlYLHjBYI
vAaJmHGcnziRZrP5vr4MbZEM+mJxOp+93xY9toEkTQJhmZLXQG+sk2JSxCdOrDUN
i2svJyCxkkvULU7io44y9q+cHlSNHilDWeY8g65Jqw9F9Mc8QI8QHtn+Og6E1pKI
zKqxJMJsQz/D56XB/FhrzTk5KlrSRRM27JYJDhWE8FcnxerVwWKiP/HPzAbG94a9
rHja6OANNmBVudlgMTRgIOPh3KCUPvu+B+j5CPOYR+OKSKwg6FiQM2y1NjszPPjB
o9LHmzXPa5/v6QNbO1Holuneq67iJLCMMp5rNeE6H6kSUhxemxr1PZeAs5Bdci7z
X1XNN2G0lmGRmaNa5zbx+tEhcC+NDYfQ0IlirUwThdh1h+JmZRTqB/IDXNp/H2vZ
b1nncuyCcdTO9AIVZrY7XYocJd+CYiNROQPOvLahXTa/LkhsA91BxFjfl5sSLgaS
Filh3QMICLRw3ZhB8zMQKp7o0URAJ1Dc3kBuVQJQcWd898T+04zGhz2DJvLHTjr8
R8A+3ylM3xnagARWWHdWd14tDhrlE1GEfv2CUTfqssTFFSIHDomHVHCMhpbfN1uY
o34Akj74/D4PnC0WG6jNF0oE1s+sdKO4zKXZPCGgQtGCrZJw+Dd3JAiBxVW8Dssm
zUz6KgGmTAfaLjOF2/QzBcGz+O5BiRPQL04tncqsXuZpzAI9+Fe48zQAk92lNVut
sY0hqILx1AjtijCZJ9ygFs9r2oYbOrGhOd7jcKIyLh4lAh1wWj3/RolxaXvoydxP
fMBiWlslZECwMQml5yNjbU77AoLnCbvikkwvlFuErPxjvqA9FWbotrYOlPGfEhyJ
W28W6G28DXQYUnKv0wxY/1txpY9jqd18SopfIgRmsNCrmffMi4j343ir0Wp43Vzp
5/gu7xtk8KVP6Pao79+LUQLFrn4cRTEM1bqWDbyiRolUVAOZTaaiDGMJZO25//4g
sOmLN0b6QhLGb7+mzhit5ci9WLAqBX9M7BJ3B5if6TxTMHlkqINWan33//ruPYpR
yLQNSYLPUOBt1SuL01O5P52LIbZqvs1qLG/3y0vLj95tC/WaJCvI3DmGKMn3zEZq
umRrLbUWwYTtnar38ABf05j66n6ILl3oPuQEHjpS/FQvDNNFJIkQzrLhhAXQC+RQ
pxxpwPc8HGspeQdmftf7sLXQ8nBeTfPlgf1JHH5i53j3lzgNqlz8S7OAhRi8Gy7p
wUdiRhzhnmy41NbAe6zoy8M/9sBNMThE2TuYHYKlscrZnt16MZaJAjfookzr1FRX
vfsuguFqHmq2OKpmWClsG3gHVVH0z4tBlALAgyZu62KcS7dPxsAygiBmrrtkqLQg
Og5fdNnzbNUrLrqxewWDdLtff/usaXeaf7Z6/r4f/A42RuPfdoO453eahLrBAZhQ
ZW+XlIeX/RYbdBHb4Ck4uV1zXxlhn1Fy4PbBea16MN4N7s+mej84bKkNwG8hbpg4
wmeYh4f9wPs0wFJZWjVUaSbjunZ3qwm7vAd6CisM6HDeEbkyc3omERT28WwWMrdu
bYpquGGJaXrvlFZlyxZ9MxTzL8WEL/Ghpu+QE8VS03MWa3hf/hHa1N6BH59mRXaQ
0wYyyq15BmKj/tQOtW+Wwf7hLqxgJg3xgt+22sroJkLChevjV+QGl1JVvlTYzfsU
NUXajBIBpqv5htBi71DbmqLGv5w1poEs2D2Xhne9t+wibKety+IP41pMZmmMgsLp
1aLl+tMP2f9Ze4clVZPvlQgnsAijzvlZuMwHm1CduWMOka4p00ErFTkINmAQ+CGj
SWY10rxLiYzFdoiN8CXYvG/b5yHeToQCjgGpWIKM2B2uhr/PlBewJZCmsF2+QFyC
Rgxddb+INhqENFxdvfHzhyv9I9ZtfQxmmaf1cpbKNDoAAis3jRi6lo7sMoiSWC/P
Tw9MjxYc2ieWVVDndnobx07FUMaiWdrqbTnTDkfiXGTFbgQIR7CVaz22eyw6bAx7
HQkcw3qLJvw8hTQneZmhJpD+WRWTCg+fHI6BOZvn79uVnn2SBAwFk0/gzRKqg+fU
SHZQ+o79nsQqq4wXvbF9Q8RVAK+Rr4y7PJt5eDBzlBjpwQzWDFkQWylC3yyUVyJ3
B+QqfbSX5VYsRDvfiHhY2rfqI4r8SbN2XydUl5Q6Pp5NP4Ll1Y2fBA3vdMp0ziHW
G20jZfVUaVdlwojZIGFr6x+NmmlB2Em4QKKhWksNY2BtHdxbsIQ1I4jF4Yyy0EiY
E3ZtadKKV4WD0cyN4zRY9v07hvrdw3YRVjKUG9kda9crLDE19iTCF8FHONl1c50c
tQ16fbg871d9xBcAkDsWDIp3r/TGePD1TIuc1ZDeiQZ9YI4exRXDpnTw4TcgPFCx
dY5dhPCkd6SVc4qUZMCyzrz0CX+VSj4Yyd0Wpsk9LohQTiLwBlVzBcGDa6GFGNbm
mK6QYsfrLSftWc4gbsp120deGk3tzMxIKXpCMlH/6BUGBEr++OlVcvBwN/SysIzC
KcwFWb2/y73wTi1Ikor9BX8Kj+6nSQFiaa5KWb8Ku3HiqYi2f13rQVBY9lEryqTy
6V4ECoLyRPxG4a1oBtuTI1B7ZQ8Dv5F5rL9HfFjbIWoburiF5p/GCEpS97/D+ctv
YRJaS65xvz1VFq+YBqZ19xyDP9JMePnD9pxO+dZEEowbqjJgNl1tn/jKH+fdPMgN
kJDSdYTiFD/W+8pXlazKdThrsGXFrc+3Okp0PDpNjxftQbK6y0PXWF3dXxt8EXD0
Zxpa0H37nfP+52IvRFi6IK6UO3CC7kWAnn9WSkAXWCQpisxXe98wVT1j0w2IuIhZ
+TpoKX8e7vaNzk3AuNtPKERRtyblPjXvP+ki5PTjMiUhcwRcAqFI21hCSOT6421c
ihKuqlfQgDNKIIQxHuuZ9vg4NRmWTdZsXdiZ9bLJIQrn3XMIFIxqq0dQ28GIDe2/
8qWSDWo9TCYbZSPc8pMdr0OMsK/2n/WFpLWwNusdrDQB89bN2rd3P/15EQ3VIbXe
4p/bC7AuVD+aQu/TzOA8yJB7jmWCIpkPNVezLKWVRRqfyOfu8K8PxSzySebNOAo8
/TBtSypEH1P7eqkFQhOiYZsbO+twAYv229YzPDOZSSLaCioXssrOwe6AGF9SjQh7
oXw8vQEScNgjtpzI1rHD3OVT8xxlNoPCCFjk3CJSMkp6z+8vcJFtuulyv+s1cByH
YhxZbqEf5FhXJ8lDN7hTH44VBFd7HsFqqaPFSJF5B9vTgZZijlOOS70X4KWy5IAl
0Tgu7F/fKtTgGHxkv3+gMSyknIyIB2XckyGO7h33tLeS3Rx8OuPyE/IqQapswi5H
Ti/6MBAXLXRfpaQOnMvkB33UHGdCG4BUb2XhWDWDFHEm5nm34ibQhPwhSH4HC3l/
S9ZoCOxvE9AfEmya7q0RzBdHb+pl3LmQonE3tPMt7HhCXRPbQIV09vc4mmfmIYmo
hXfFp/Qmi1bmgifonkEC8EofTgCthAYjnJHF0njw8x4L9GrmQ03w30CuvU8W9UBR
HvEeJmGblsupDs8j+xFX7h409//rMW7IdgEuaU1LH61jI6lgxbWg5U5CT9602lvp
dTKlQ3Ru7o59jkheTOX5kb+O9AM5+TwojPPCbtCrlOIyQKZISOErCUGRXgDA+QoC
+ht/cc1o3eniAKnhc2yhpTXon/ljN+L54ug+YYxzntqC/9msstLe8J59WD0/BPvA
8UyTWkEHkxib704nSqvYXwJnIkfGVHA5DJW5cIxNtfRFfZ/ba2GoB6FKGDnY9hvH
jkMmgQxRrIGoA66PWZLuBv8BgsdWY8/E6XGzxNQKrEppACCi7kLdFzIJMaUkz6zO
IxU2gcpK7TusAAdI/5XdZWko3m/8LXh8raWzJXJEgToFtlcZ9389B+iHHky6qSP2
E/xx4PcYMs/agPX2WwlmFSBm70cVlKhpIiDyz9fS9jSMI75vmDkRSyR738iVjDNJ
VFKXL1l39NfuuMND69NOFjHttioERoRAQ159P/21UAdRKUEISnwZl40/9wVULBv4
LirLP6kEAxXSde9bf4YFgSXkoanHtWpeIVWM5Voxn0IHRhkMBSKJQ0KMZJVP2sWB
yB58jOkDKsPR2PLg10VpvjJ6uNILJvql0xcHfI9pqY9OH8VtSmP+/6FGEekcfbQt
xH3MxDfygb5z2Hmh83LRrUyt7ojbWEnuaOkXje/BjjjYpPBw8W3trmuEIP+Q9IHM
aydDzCClQyIMnQTKRj3d/7tfhr/z3hQaIZPhXCDHA5eEFBsIY/a5CipcJxqQ7AI3
ymDKOehwilkFq29YMbdulthvtr7/gduzvm8O+PenzuvFLmsUtJw1GE2/hOAObmKM
ktqlULWwRavAppztD9rPBY5a7PlE++g0zfrcpZbpc//0OX/fPTbcrvJ86+n3Fiye
zmwloZAw5AvDF+f5yfzH97z3rt1pMl3Q/0bUPN33nYFN9uk6t/jM0H+y+tYPpjtG
Scvi+kKFVz9/Zt73mKVQSxoGxn7Rkqko3k4V5SznOElkbVfXbvMb5DBT/pFPgDyQ
DW3AeyMOkjWEwA4tTiBLRsBmjpRFGvDWMzixvvbVTE39RdvdUYgnddCZVMUQJNfL
oje6XPOGeKXwcwPG7LQ/M+9DmKdpi6ZLTfP4bNmFPVsWVIk6yeUZ7OqcNfm/H+WM
Qcoo+qWcHe2OR7GAu/moNJSfBhaQxrVSNrTvNFVdOTvabwD/vYq7rT0cVchTPQ/0
6T7zs/z9zxv9L/vAER7mIWG5To0VmRz/us03XPjL1PdaBksxMfQifEhFY3S4p9fX
M8fg+WV3JeSrUPEtF5Y+EEsBXiuV0BUpiBrZ+ssLNQkb3VQB5nzMEHNjNHEmeoqh
IQWSQQwSHB00jHvkyfpKa/+eeaZdtl3gE1au0eBU2DFJMF/jLZ/PqhuGfbgWBfE9
vPCIlOzWGNI93J6BG988QaUl8WqOYiNmaIt8xWUo5XuwwdP38QNNWa96uLunbBRw
e8EgxB8FxyemAAprlfo6bAKc5llqJK8toRhaGDj9C8WOoFgQJgo16EltAJFN3uX3
ThzgN7U4X0LcBmo8KUDnwdejQgVtj60sPQN/b6Mz6z8jmkZxJxu4NrVWuCYrWxvf
BcR/YEWaT+hvwx5NCO+IOiooqOM65mdAmMUPunm+a5I87sXakL8sqOrwvIf0f4/C
qy7k9NYbjEJireTKE/SegrTvTcv/23QEKyJZWEQeQ+cspKbuPucBioE98YQkB2aa
URN7D2FiY710RGibeaIFYiJOz8f9LhCGYWC5oAqHpl2rVcrPhvovStjqBR93nr/n
H6qZI+JHoBfdLfPl5918k3Is3IQYF2XMyz11pPmY9/uhVa3W7IdgE5dkF9fuFVEu
35xc/Etzoi5Jv/Wy8D0fBuB08lSalDG4jpC8RY+kOlPeSAAAvcoItKS+E9Emeh68
ALEzuKx8SOYYeB4vm1ZrSHmJNHubGH/AIH38o/E8+/Ku99fjuR8TbuJjBTGiHvsU
hslXQ8RtUvWzgxwiOqaA0/nw8lJDj1W7kCpVNy1AAGvJpyBsJfzyJ1hDmQTyGeFP
m50nCXmvWr1tEw/9Ii3/D9nnf9MMPjZS1uCClYxntkzLr+8hC4Zq3ARjKOv3AZdA
DltfD7PDpNJd2WNpm1xIrNNMWr+qtDbvvc9w86s8PbSiOpH8B/n/7DoMf5pQb5IC
72KSbnKqD5EZk+dN/l2NQ7noQfUK2aKPA4q/JweKigCn6obj8S+Jtbrp+pix9KC3
MCZjMOlfwGTuPT84LPapVmsbV6TbgKdn9Ma4Q2GhMFHEflNhF9oQc2lsU9d//bhI
xx67fL8PneswPwFmi7AXoB2N2tKkgYzR3Ylo5Ci+poUcRrBlC4+qcwsA4Tz/9B34
/u4vFsuoT12JtGNWtFF4GwIOB1MHEsZ7crJqbXpYqbSe/5Wr0ato7pjDVD80A2X+
rNQ8atctwZao9JGb0LzNAWpxFQLowYuc1wWknYh+RcRXRSf1HzObXnxswi/vrUqv
jh89AArZTtWptgvpQHpOV5fCLl+D8eow1t2JUoJc1dgxYIzjQdRCMmuEyHAmJnFr
7L87HHCxuXMDZQlY31/eeeBgKBZ1xs6lnpwFAAm5bUU9vv3NfDeSNFeyuE5gXVtL
3mU8flmlpadoJWtcZH1OeizN4vn1S0IPcZp0IeZTdxmxorTx+D4M8xv+2tNi6cAS
wf8UqUuPRSLIQXiE/c8ygvP+Va+9fPw9leWrju/z0JfuxdUqviSa2vYKuVMiR+lo
olubTcUEZTlOvuP6jiWVrF/AuuLaNbAem0nMqEh/GJdfFUtSc5zr/LwifwF8MRRt
9rniC2Fc0E/tlDlxIgYAfVMF/r4EENUofhkAfscjSTcqN122jUpAmM6A3MJiJYlf
ioaweSgkHbG+JwVcjEJSOuAlM4TjpGcqSUh+lkm9OcsyJiYMUqISyKoPlTzkanz4
B/okg5sEHplGgfuN/AowECDTBFjGpCUbEu0WpOCgRv4IPaVxhzLnVE2T6GRwl4T3
ZS5n+qnQbXKWJCfTaVsg9mLC2NuK2qZAT1uyFp7zF4oNKStpYTwtLk7PJjwFpwPl
MDfppELznqMhJZVVpmlecev8Gb+yeY+8UT+QWwrrfqSWf8xAdrBUOpqLrZQj/qoi
2ZhhlG+zGXAqrfhzyeLxGHDE+l3k8AAgzBTERJNbHW2slbT550YZ+e6WIpa/SyqH
1b49NscmzeMJCbAyOCeGlEydSUUBnyEm7ukDF2pDeCIFE4x1tRaLqM5jnTWRXfCR
S/7XH6xipWSRmIFGCq5RyftvOSNMJdr0U2SbasxhT7sxY150cdRCKK+B9InWzl9M
9LN+reckKadxRL9JjE/q0x3i2mFlivCoNFX0Pa3yO3Ff784MKkJBKx3cdCKptxto
eBuI8Zz6ERt5rOPxVX4L/Xrrg3ai216LCRUllU18b6wFgzhkzZDBSukpJl4LkX7A
bWC5IJHy/wKVn+w+OTmFcvba5JMvKXm705QqPRcDlLLtxF9DOJ5K82NUlK3VXEKm
MzFexIVZuhTV6QtZiuWDwLv8L4VXz1kHtdyErHg2Te3UInM2hSc6bWByDB4BkhB/
h7O4HeQvIPJD+wuQv2xW4uU1Yl74Vpg88qXhWvfJ/O0FWmF6NYx4CICYXw3HJrP1
7Ydk+71/aNX+omJsz/CWyVrqQz6ucZKDw0d3MhMB48JQ3wyCDEiSTHWftcGnIKbs
Z1OjfUvneG4hpFNkahPgJ5RfNIp9uri0Hji7whjFPVtpuklbjnFgvbnM4oiawLdo
QtdBi+VeP3svexBUnbyn+XrxYoWSYbD1nBmpyYRr+dzAKKnsdAXHzvrIma0MPqeG
K50YghzXhxm41GWDXWBhmTjZVYA8RyawmGkJ0OHQfRv+f8K5GWQptx+16JilvvTv
Om8Fr+F4mTjMBOBwF6sMsDXZ4EHwNeGKISMBjFcSALuFAy1nGpIKwjL6MkBiJapj
3DMTqKKfCHEcIgCoq2feO0JQbJhGxIzuHXeYpBOyKxXK4BqK6lTIFVzialu2+r4u
0FiM+RmUEk7Nm0XkDqFkLj/LxANTM8K5gc3H2b5m95ID9R/JrXgCtqbojqvlaG+e
HNFi2hXT3U86lbziO9uRiLRFB/uVLlLJi220WFtDMyVjXPSeXO5v1ZjxG/2vwwkT
HgGf2ewG0W8TY/dq4CuUmV/JNwnrNLTL636pWKQVKLjCR3PySJuDnEIBVvdmcwZ2
NvbfRcBRjIIFtYfi21tKM0knhHpV7PXp7rmppu0cZd8wPt60O9v3SCa6zw0acXp7
0WbkYWyzC3WnKXwD/XpuCa7EU5MP8R+BG3R78a0O/9hLwmcjowjC3aI7n9V8+XUg
z6SvCDUoR6J/Ni2vvKXZ2FzFcMxO5UMnG8kbkK+M3+l06CnUaM2e1erlzNdE7KvK
0Kz9pF2pW0ALYZ/fje5MgQf/38KekqsvGIgcO8khKcWP4qLhKUFGyyZXD6EUfzQn
NE5yQkPO+ciwxefWLjvbmfRkQSp/vxfDXm7T5srKxZQndX8DzHLs0YHCrjqu/1Zi
tLkwWwDCDr5Yx/2O5+PqWZxizUMMI3QuqTFVt3Jy94YHcHXFrAVRORSAPiQY+QO+
jdLtOKiVa4DMrnEy4W2+2Z8XSx6Pmimo0gPzvaDB2+KhuRfzuAMiYyxCfEUEsnx7
nNwSjB+1pN/MRyKGozGYg3yEPOpWIXoAMihiLvsnfEIXwhU4lZMKCI/IWSc2WNPQ
Sbr2BYZXhbjDMsvA9LLKzMMvIkLIEolCoFKwwNw2P8M5xGLbdetGRK64Ws78s/UP
U9EikwioCCTVErTzg+Oswj5YoEg3e8LY7Yzp3UMbwQxYQYzlGOu9sHhaHLsZLDmV
Hi0dvjq8eiQ2i75elyl8MTTlgZ+znd5H5aCGeouEM1kr1xAcVIl6ZcZMCiMGaH42
eewo1hMAqFIVMumVkur31PsQSPjcdO703RMMA6R6Ad+DCQ3SaiB7YhKbfbWIXXGB
8V+coTOdwqYXoSAoUnb1E3Rzeqy4CKudz6i6isowzeGyRqK/Z/clF49+QdTQJFeS
wR1fz6D29cxPSgJXU6gl6oEcnNYFSkF5VfC8XSJhtekDhw2Ft9kC4KjFs+b1tSZJ
S0s00WZLDFccPb8vSziveYZ0ifGFATl5R5DwYeFUQddU76+5JcV5zL+656H8WoGz
B/qHSuP30VeWdPrvFPauxVoDwPtVQnRVD9szAGSHC5cajMnhAzF7IRL9iWaK31oB
cfm+BxQdublriKxgz3cJppGclI1uwKEtI5gQ+39F6YwhaSNl1STfZFqnOBp3yMNG
ndpIzPaV1xpmXOm3JjvfSAHJjz0G3sI5D7oUVDfkBsu32WegLBvhFSrhDzYqhnfz
oVoraKgD8PqQldgOqucHiaTHjd/nIQrkDvpwqUVffaFWP+TVu/dAADP/+/PJThM7
snIEwbC0N22hUTMvS5AceXXB68kRs4uRZwhQGkcdOjEIylevko0eXB66d+7IVSaL
FTAKxVCmr9zE/TQVpMIN2lQvwICVvr/dLseOVRvtPByTuWoN5TYXGW3Sc2TMEBII
jIlz/WNgIs339kkZjj/uS/SWMBmL6AViM+W6rwvs0ptU3yjtn45yuTCnfnAexGR0
RRBIEBJxiSUz58JjLRg7MNcV+M1t2cwGf4hKYYwx/Ee1b6P1iqPU3z5sXjHk1tKm
6HC3/++BV3r7B7DfJZejlMvcRBexKn3eF6NXaKnROpur9VggCBdt4Fx9O2C0B6Bw
Zz8+sILT9SJYdlDL6IG0u1Bl3fN9gv0hBr8L5ggiz8ssHJB1FzWbcIOK7559Qrrj
D6LLYaSQpcZ1PCgW16yyaUPKOkPkCWkfQhLOFZDAoCt7e38lBoX2GhCEqwVm3J7L
fXvZBhuRaLuWkgB/LyRAU1Za7oxWV2sUzIjKBEp6Z6ra7uDePBxqxAPa0358p8uj
Z/WUpm0AdzyAwl8A8A59DDtfB67Wlhwa82xz7jSQHicnmFU82gHCA5fg6kUHszaY
dMoc+PAqkHh3Nrn5SEn+Ll3U00bNI7PhT+6h66bT3KOhuqwT4kGIAD+G0i6eWFCb
4WCiptuSBg+9bUFUUDiQZM6nlL0/mH7oJpm3NOzTjgPduQANZemSAxck+PhkWWN7
ZAMG2Y0+6QD3VPcT++EpXsq39wmA518BFnrU1F+9arZdNi7ZKwehb6cn/nwk2/G/
O26qSiXfkn+hRj4iAl8fkdHcWue7tF4yRA9eTaMeyLakNpA8YNkgXSH/Dyl1M+sx
N7a2UcYkKuCF5bt/XUTsb8BszChGN8QucWKLApmfIBqaJ6bZWB+f0yMo2kTyFO63
vTzgWZsMH3TvlSWq6m6fB/HobisHBSFEmGoZAOrnWDNfXhLU911eGOUcUDXoW+Dx
cQerQyeZ0MG/fLbU/VUupr3+VpIpfwCl7Umq090vu2CaHaz10DHgyxCOg/9xsSMp
6Ui7e1QsOSD0OUcIishXu/NUlgvq0uHSbxAraeUgccerbMf+kP2+eccnovPVeu73
e4meJxXH7hysiIeUptGZqdFsgPZ8Su3v0CBEUH/ZAyG/PGoGa4CNJJimVKWLGHf4
R0hI5QyIKoelk5hWddoe24VUlNf9xWRLz6QVfwLQ1iCV0+92vvy5M1jF6lnt4OdM
YPkwPzuItKKlDA6H8gUTHI63f2/qeXf4C9MeiXXsRbg2HzXADTKWFdMZc+XjSz4X
nYJdOOLtiOlpGMayhyxGQiuYoAc9Nkqbzdlwo9EjNfuuF0JojfO7VSMRHxPpo2Q2
CkL/5ekwESxPRqx2Hls6yFBSkegw6t/pMcSt5iFtLWx86wW7+VUmEsbH7XeMUaiU
2gHZKDAsFjySz3AOj9OgfuR0Z0MNJWq8lMswZhbDf3FAtJtGCQOEGnfIyBaJJf1U
N8PoRihCGhdLueCgGMqGHN9GRFuxL2tdRoZduqX/xOHjUCmbXjL/oOLz39ARn31B
WbaO7Yo/TAR9gPFODckO/aNky5jYRYZM2ONhk+oHPdCINt2orfH/J0BSA6GktK5v
YW07qL8t6wrSbX8ck+YF51//1bYi2gYiG+rNJGnVWzod4n1u3AFbIi2A6fpl1ada
ED4714zvoxcBQraU89nKndUUZ/LsHzhgvziK6i55jKnVIMu5UWJV7TaEx9q9meJW
PPpKJgBfXKdX3zsx1PbktAXeqPPKUAMr1GoNRlmZa+di5hO+8kjT1ZaljG2eeuTZ
0pAnLn1rhKCaFsXJlH6R1MXR3TiL4OfE+5dDjYYxMVDVYaSjqHffEhFXhfypHZ3U
7JvqviW82VXTUredzF94q7GQp9P+M6hwCnKWPbQtjE7EuUsc7hrTAFff2Z5EPN+c
SJTL1woHeCzv0FX2zmAhQkHOQMv7h8ZDsl3Rcu4F/gcadbs6VUVfH8FUxrwr5FL7
8UhuI1KKGMOobPxXdDO2A88JNZpYBVHi8Twrc0pEH2eNSooDj+y71qLOrFPtcTFe
kkSfrpNtm7uDNKtLDWqPbFhPy7Y87verBRRePE7GVp7TKZPXypywj1ByDz/LJJWh
jwMPkZt+TbW4R/1ZjUi8vw5NOroo87XkU94boM0h0p0qniw3CrxcdLGp5NsuRWcz
k+4sEOgTjHhAzeHVA4Br+M8x53bGQgYcqO2Plr35Tx+x1vzV5RHeRwC9XpTaxhsT
no57/yLO149tfNzymkR5jVOTONgNfqhydqRIchG5yOhmRcqXjd88izQfU/Njmi87
y8+mUzj+ZaaX2RGKmBkg4LVJUaXpaF0Ndoj5ACiyevDdVs8fj7av+0xy2mZc+AKP
OAW/BA5/XFEkUxfJL+EDQX2sRA/q5SQTK4dRd1OY04eqrbbAvT9/17VLU3o1gMjQ
Ok4955zVLZpDZ0H4I0Z6FdeWz8VlKsmVFhnHYcpr7JsonG2whtfUZnctkAqyennx
g8L5q9gnEgAagL7eseeope8SyVQ2D7SBGABuyyZ8wF66EMakap1hfTxHOhUWTdh7
/q6JF8q5rVglwfGt0ruk4CTEE4f11xb1EM7aavSljigGF3OTsMk7YZ6taSMPQLNS
5eZhXVafpaQcWtU+yG+X4WqLRfmy03n7h/UKGBRHGOSrAn2t9y3az1oU5V8B+edE
I3LKXv2AsI/lbs3NGz1CRb0DTCKxOEUzJso1KAyWBX9YrKIywwkIGRgVMOKgKNla
QOnfQtxepw8G1CToE/YYRFYu+kjbwMIWwYbuOC5JLOm3H667sgSpU8k0iHNaQJKp
StvKRIMwHX9n5zuknsDxKUPtVdCDBpQ0WlBdWPCTNW3PwMrZUieUOjp6jRTX2d8I
tqJnN43Qyyjy7tfBRKVUt/G7bc27Pni0vxAPSQbjj6LCNiqwWZd56aIkdoYUReO2
QEHnTtTmjE8NJgl0D59232VvnDDUswz604gxCCEX+BG/DJ3kI5sX85xWyg0ICwXO
lgL6AJzogHWiMdu/fxdsAOEEO8Nsyp1+PkSXti39pEz8Wzn79Cq+d9DeMtpQ839R
PZYE+tQ4kDuOnGm3vJO62H4zQ3T4ZfuzfATQwml5kraxVoaG5PkUrPmBlpvtRNz4
dK3cQKXgXssP5w2Be5YymuUeiLoAGcjJnJdmMmgbLvZ7zDo+sITf7Wrp6MgHcv3+
uIWiducMYxTRDSVIGGFBh/k0kfWl3skb6grVAeFqGcSMoCK+DzBfSI2I9+VybXWY
F3O0ADTRkJtF6o9VBs29hdZ4H/vulaNxu8E71IxCyamJEhQkuobWRzKltGiIU8wJ
ljxD1Ap0wh9husQ2zc9UXy07FSJh8QPteEisGs4FfKQylQR7IydSI/tOnjf41ck6
qoKKjhU7b+OKth9OzQ+hJnKFexmsXWe/wGeCshRXkg/RKRPpAzgTZX4A4mD2rAS1
x1vZYTxYmC3LfDc4RZLTSBK87ua27ZxnHq4Ctnywc6aCWLiKcYoSxycQ6YRKrM8q
x7+6pyd7CfPAmhzl+SOGKbFB/lgEIFCYn9/4w2pj3rm6ThFVRY8vOm/CEeBLvTaa
DwJQMJGHdMpRWV0RjJwV8NkI1Fi8S3Mu9QAODiFMZ53xy5/1WbaSnn2JWyCV1cIR
AxDaTddPP8YrllGp+HgzVznfb7pu4X0WiffwMcjhxVvrmFRN2X41EUmqGrZp4jJ5
U6m257Spx6wdJiCrDgmUAKFzP2U88seha9rj/VX2Ed8nwh0uF9j+MAvsjKY0ymUO
kfeH7qYq6vIuF/Wn+Q7XWvV3t5zfg7QIJuckuQCGrkGtioSwDg7UZ5FLP5af959q
NuwqeNz+tnzV/wHcZxzJSAsMY4kRazrq8CluwTFKUF6DgL+MY2noSAW3bZVoAwMH
Y/rpd6tR8LhF8ecKUKoa0so/cEmwuwti6Tyq58aW6U8uOJhQuSw94/Xrli2j+IJh
btTCEUqUTvKObtILwBlEZDA3lU4ipSi04D/JosYfQhSXjTc6sL7oJ7yDYk4IF6bi
H17awSFKjLBINsTLcUhcx8ff+3DcchFGFdssaYdr2+R23WvDIlpbeqclFSJEpTJ1
zjXEcNondJxWIYHzpwZwydRPSXsX0GXQhv4J7gJGk6eriIgMN7wSh80/kRoe9eYG
w2LrdZPR1iCnWlfOuXcdXxXfe/1d9fPrU6XorUQRMo46842QSYF+EilfxR48mCX9
3JDfJBWSdGar03BFxG7FhHJUTdMWDZbfH7/cEP8lMwBBtIODnN6i9BKxnHMEltKz
jCmPsu0OgmsX7yKR2ZIbkBGMvGNK3obVlaSz98SIRLovA6QAY+Lo3vY2a2+7L9Gg
83xlm214L44KCUOttZeJF1Ml2hbKciBvmZwQBIOvBMGmOkOhb4fdxXRYv5dOEg5q
lnhp4frByHRx7qR/H/pQX7zUwrmHCmiwo2ukD3xBdhsf9eXAWqWFpS1nmquv6xYa
ZilK7TGwEqF2xqmmkUZK1BRP80PkZSPDF0pjdZ8aaTQg0HSBnIvaXypxt81FzTgQ
/94ab2nU5d6hb2iEMIkcG6lxsximhnDGcpaYM36+YiWUv1FfGgTUVBECsQ1pC225
i1rwjKDpG1O0myMb44d3xGTdhdOso4j7tpHkZx7bBa+JUcAzC3n5LsvsH3zYFkf8
IQtq9/qwYBvZSgI6+RcDCm1TNDaswyZxrffLNjTq3mndzjGoXtGJJFwDcPLsGI0e
qowKNuew2EscAoKehv2J/1i+OXFthT2qnkVkBjsSTlx4jqvdFo9Oga3uTGlUvmPH
831fgiPXkkYxO6jCsVzYPgKIXvyZm0mvsTDEfFyuLqfvhXEY5mQkFvf7bGZurTZj
K58cPzF+FKjjUdlQ0k4O8aFNwX9+JPnSq5AK+6hiNfocELqo2lrmRhDzlOeCo0H/
pzGuPCeVenyXss9MO561wnNeHCfW0QzESbLxlmJs47x6E+u1Waqtwrw71AMhovcW
7HqLzoxmg4hRHNzakRprEgmkUqu4WBR8PFSrj5tACVSDpCf1N5nJsKN9/XuyEgXb
rOZycWb/OdA9ENC6/toyHzh50u1csZX7l5G2lEwqcKrfpjSUXjbVnD2QrRGokPJ9
j7cnzbT4TCQCrdm1pGpOxDwiYAlIDC2OUJpS7M3U8eUiDSQOVVjzGv/eaCsMF+xu
H5CTYEr/7nkhGvyt7fRhxNMbLmeQLo9comFuOa3+y9WzfPQF9dw55G2deZdTY1vg
QdAUbgIzPRM1Wpc7hLJGwFiDeNedW8qk5LCQPoky3gO3piTpWPs+MMILEfS915Uc
VNbBDd4zoy02p2RD3WapA/yyG1hSTMSn6/1kwerumavW/00NkL8dJgtumZv2kKA5
tAfGEjTmD0IlLuumfGnNU1rw2joghJOsnsaeMPmQoyqogA5O8H7Pj+/x1voPoKsu
8SJtTlnY9m0tSIoYGD1SvpLEmvk+6j6edOaDkpPdNN+j+vZk4lXOzRe2su0dED7W
odi9OtoS9TYeY/vaPz1jGLoAL8omrh/d9P3VXVL+q+VUfKfNL8Ct7ge5q1f1Nptr
eohiOnlkqeZDJoVhPUpAIeCI1WBG3faWKRa8XarpG0Vkp9atrO5fxw5kfTEr2Bvt
cRjm+RUhFMJp3CtR6eOtPIAUhOmRz3rF+itk7bmDDHKahu8jv5IN8TGdvWoGNYEr
Pv54cYPnReaACaiKYRTreWc4BQwN9QkAh1qvr0P0Js3kW3XyVtr3zbZTweH2AUu2
ndjVIzL8Rz+cxPSFVl1DVUdq519R+BPa440D8RhlOjEUJvDhhsmDvPgbBwp2ETNE
csDwnNXK4G59Sz8sh/fLjU9de7qlhBFq4Sg7D1CBrSczAFGs7MSiDxyUb0+HUAH0
3JiMoB+Krw7fANdMBOcKX7wSzd+4iJgf0mnQacM4gxlChHXvQ2tFmck2DjH5ryyN
tJe4/zMynJhsvQSTY+CVmeDwPiwEPo7JELsERH1CX4JohXzxUiGICjZnaC7CScZU
q/yVwQE7TkUTKIZA5SwnmS7rnN1pRUwiEzlzlTkUa509jRXyUf1XBqgKnBaumLqw
hvud62kiWUima/QFGz5D4ZE6cdPCd6Q73f+9KJuBZYlKqRZbmPhtvXA3pYH2srVb
GvvQwsRMsylvZh2SeRjGudHYDqiLszbC17P7hPKT/tWxNtEJ4fYd9APQly3/CqYp
NP+3bzRyDDb+rFC7Npj8cvRtu+QBvr+NiJVWDiHSVzGIaLCwOR3s+g4Ra5khQiXN
ssofm5zClaflGy13qsGzGGUCrAM/Sa8j03TkSNsIUx17fIMBHsRRKEdSeNMclWpC
jN+lDk65YEEDC+tb/5nvl3lXSNU+pgUWz2+yj62+OxGPNUQjQTKwHcwjfxD4DGYQ
vwX6RWMePRLU0STAZya8oa+/8r5N/9jRkrJTNxd3wTujUK1STRH27pvPiXFYR2Fj
dHch8Sm6oEIgpLy3LDfgaM4ORcdbQwYn59+ZfOB5L7chkrOKTovWxFZacWjf2WJx
zoHjzTjpVd6Jx7vc/Rx0ii3xzsdmPtRR3TDi2qEMTwFMeL4eIjct1WpoR1j/wF/8
TrBF65d/5JiZyf5sMvi2rSPxNa/L0qqFjZbxLd8mjBxqqKGVy/X1YtpAyZ/hdOr4
vb43PkIpdGHOc+prZt3pBDEpOEcg4C4xLDq1AY+NkNm8JwyYysDSc5xWcbr01lFi
8fTT9WYfpoYKEy5s4jf/1thWqsDczz1vE5FoyABqVEh1+QossaeWfY3QfZZUMLbX
MNGBnKJB6hRzpT2Nmv3f30w1Wb/l1QKJIq+7Kf7gdMY0wlU3tGyXvOLv3wWpR8LG
iQbnhAop9JczF4lyeFJ8UFHtxov/VlEaSwOl//PgEksYrVXL4xN1MAbSG/1zlaKP
2c6QsIghwYrds7MTFB8vyG7/9ED03fjydGlg74n2kTfPM3KUYl31SpHwCwQakH0G
h9BVusmyvFYIrvTswQ6BrFsQcIUCZBkDLrqs6dyoKDD/6UvmfIevAmcWzdmR21dN
ofCKkHwJ7Dznufozapu67gv12xU9w9kOU2Ge0i0l8xKxBqZJY5nvO0iAYw+6xJje
nu4N3OqIRTfQPdIvTgRZ+Cv3aRSqz/rNxG/0AZZBXrtBySzFp5Q8Vy9iBL169y8y
gL33cQeTmTg/VOxxB+ZG/poSk6NLD5Y/3wqudL94g5MBFRHKdeMKBEG1AvmBVlS8
NsOJ3iYZFkKDmE34QkzAUDRsku7v75Ez7yqXZHrDjrarziIDVe9rjkNZNi43yaUb
UW3ogSFVyR8nzsL8r5Y4owshYkO7PfEPtivoH6ZtacgD+tZRlITEHDp0THizO7GL
jTdtx51fIHv+rcR8zrZJxuV7HTTqgru+oYyHclTanthfYHanvfba5pz/jRMjgXk4
9osUwkY1kE/cPlrmVHjYheaNk6OTf5C9MlGtAq12ky3jJYp5lKDiqkVUrgSw5SJc
w0NBBdnlkoxWSqwi2Wa3TrT2DtWtnTl25IaP1MUEQt5FZ1fFDNr0+NtkXAALwwvk
KYv6E61viTJbY5bXV0Xq7dz49jaOmmiJY/blpRpBWeKknjOPX2z3QY8+Y+lZs2jW
ziOh0Gh150OQg61LXsYEbVGlw4Z8xxbaBQxaAtODCDXrc1cRTpC7wpPOXfCd6EVz
pu/bgZPpyCmw3E8daVWdnjwzOF6vLZxGoqv6w5mh/DHhMQeJPB7+0YFi5Mz3ovLg
oKzQgIKf2t4V1UDvr6fx2BQmPdrWoruqJlDRbJsyutTPIWZz7PXYPdHqkMB8KhLd
72RkMuahPpxu2yvV3IWv/repqokkATFKNv57GJrqL6WMplZ+McLH+k0i6h3Cfag0
6KeRH3W9UGeV1Y+hLV2y8xmy5u+7JtMFBHirjuXTSUzPlqdUu1LaCHikBKetRCBO
bVq1Ks5tizeIXcbM9kcl2qN+IG+juqgx57oSb36YABz7SQc6dssRiU0l8OqK81d0
jO9MyeUqCClhe1te5y37z4u483k2ClqWoXIDGkFkqWn/+Xp4Lk9l2E4khK88bnBP
DzwJiWMu90/+Y+Kft0wH2vE+8fk+l9zWLDBbbRrT70MnmtaZUlaAVzttaTFZlnox
KC7U3zdRy1oWvQY3LIAM+/6VbISlIEA+0cIfmhy0CNlM1UrJh15XkX/aOH47iSOP
CvhsLKpyAdPznKuvCpNXeVZiKd4OoZqazO36n6E9QVU73rkMVrVGOYeFot6LQXiy
5gBN6k8vtFIhzjCNZifrOhLqIik3v4M2yL5iBdghyeM6TTHJqWXI9l6Afr1UU8mh
KQ9ej3J5eEo8PBjJ/NjASfqk5J0jts0YgF9RSEsQsRWptsmM+s4HHavRArVma1Lx
XpoLkibGSu/koPJnIhWJTOmgutqP1zBZ19YuarmmWDukCM0DyYPcNsEDnLeq6SP1
bHw5tINAxmKBlT+YcsqQpEQsFO+qMKlamL7s9405JsUztx3Onfh5T9kJEQGZpL3F
g7323GvFF+tIyD62FlFT1KdH9KtaKKl02MlZ2i8RR+qDFb5Gv+i0rDy7wYN4fWKe
dXT4m1eBosWHojnp3jhi0wadGpZVm32g8sZlqMNn/afDNAGc4iOHFpfDl5X/+1Mu
KHsffOI7bsDXXpfJIroDqQ8HnDMzco/1V/0BBtC45d6AeqIkaow+lnAWUCjqxyNi
ZYwusXuZf9O0inM41C33x4WAf0sHdYSMVGMczlc120m0QoJQ8RvFRbB6JZvyu0gh
y5Yf8QFZ6cHXVbbfsm5rLE117TxWSww/cs6QXRJlqMAaeaR9wy/qbvmx2Wh7JNWl
4thMi1NfNrGLm+Y6t/wM4khW+2tCBnQIR35EjbjPWE/REptXR3YY6U+Vv+knUXBn
0F109XK9ahI1xuSIHnvlhGRAhVkLC5AcyZoR+z5O18UjfsgvrIWD4wBKpa/ZmhSE
kXxWJ0ym2j+EdGdC+qhIK7N/SR4or8lEobAxhekHTEpH6G/VmkPmF63c5I4qDV8D
AFq15YF9Jm47yiMOv8ee+uRk9RkBomm1ik2kW72guVx/wcdOu41rOPLk1CbryUxf
khds7/zzkoeRZUkUom7JrKocquvrqrfe5V/fkCFS+khu3pojVDROYyFk6KCTpU9C
lu2nA+F8MRlFVdYR+XYdiV8j+8mxk1ZkjFlY/muswOJs9t0ueTCywU3t9g7J9o0B
QW//p0924E2SJHIZgHguWctJKYlq6nn2djdp5QocjoWuui65azm8ZuzVNmaCdL9S
9/cYMR6gIttLHeHdactuMRVZImT2ApQ2PKNEzuDyy2bpJhDBG+Cv1DiJsV+2wi2l
KFtuf4oaoU9jHotJZpwrzFGlunY00Lojv9FhosU+KJ8Qs0RbV3pswr7ea2fEGwXF
ZJHMLot6sRzcqY3c4yV9u1iFs0RG50KLSYYtnLnyDUw8JsHD8MitgNU9T60C4YWk
7RgruQZesOBp6LpwNen12/+zuDD/xNlTrFiEuJe2ljYBuQhfMm9fHx0Pak4Z3Z0O
rNW3ES8XmsDDPLpbZTsy5tC7SRw55dLV9s/V5xh94Q7sX41gIcqnI5rxosfMPbCy
mgpUSRXpHv863BX7eSTyjlDMEk/jgfzIGUg0tvlM3LsHRMCq3EgT6U46V5hNCuNR
i5heWovLuP/gTw17tJx8OK1kQcytWrf4zhiuat6UE98v4T+kFV0y7VY3srBcdjhU
hAlmhVJ56VnHLWuvH8NXIi9BgsNBeKDIcbe1KbUYXqfBvDn4gczo9HP8VT2HaETD
qwRH9NDBUwJ8bp0yzcHXXtbWHhqca3UR4P77bkOrIIDRD4E0fzs3I0hYgf+2QaPX
uxhKIlw6q1iNNUf0C/Dw0B8s+OZlGRFzLMm8UdPbZXUSSaT3vmbWOeZi7f4dmuQF
lb9i+/zJsn2ccxaOntGNjIpordrFemraK7kcp+SSHiVUdQUewOqEpmMvzeF3lA3C
3JNDanstNf7btPPMU862XKALHy3KCwc+GNlBHdnsrUVIpN7ch0CHFH+C8QqgusKp
duSAG932XPJNjNudjoXHdIsyOmyNDHf7Iy6Bu94ciPSwNqiSzIbwGglzMns86oir
4wKSnowLPz1swgb4WsXSbPBIcJh/k8fJcCpkUMidc8JtscL6+qz7AJxyoG8d4Uju
iiK1aN/2XBsU6iR9EbLRm3BMmvEDO80brgQvnvm+dcfhw0uy78YbERaXMKcNssPP
6G/fRndFRu0M8sMveca/qKdE3bwTPVxgaAKLyQn96warzxbFCSWGSPurb33/SeRL
86IPE0wScxsdmjlq+J+OQmJXQ9jw8oOYwBu9du+e/2vfMxns5rclgKXC5qafqMwQ
BR8NHRkGEIPCY4nzmmaZHqppDDtPX3hdtu3J7Y8weJKto/mK9i+32IsiwrNR+R6r
cTWl2pEvEFdXyS1nDwhA+IntgMmC3YxZDAn3GHxcQBoNB+h5xoBouY5IH9aXmuKg
6o/6TtaVYjFJacCH4DGVtqBxqJRGi/pNOYB3MipiRCsoOJWVBZEx4b78FD+U38OM
lq+DTZgSJUtoY+rpim7l+DE5Enh7bcr1H7ze4Po1mpoShDXlfvvjLnYh9HcMEdTn
Sf/IDQorsX3/2kNslVO/mFX7cYrJO/Um8QctLJaltzOtM4dra7nxvAL6gpz9jDOb
TLLka6PyEODcJFYTfGgu5xQ0RNzMw95MYZ+KXwYH687T3dkcjCWKKU3IZvIIAMYd
j3eUES65nogK+JQlmVVwaj5MWv/1TRknqp/j/doN2ukznP8pHNOWy6hmaVGg9DwC
bd/6XKqZiZ20a9mJkM26azTfIuP/TIRTbuQjdYUdqsUZMJ8KdRo1dvVmFlutf0Qv
PWQU7YC1pUxj3Nv/fpnr73Pct2KZvf1dluwCVdRDR14dVuOLEYF+/vPe7T974ITr
MjXZGns0wrCSDQJiMRpzzQ3XwNqw1u4bcZJhdOv6YEmJVLbDw9V48rgbiqJBvzO6
wyXWUJTYJX8qnauLbsPH2UkZKFK2QJtB14tAU+BZvpStxBsH6kOqYT/SKZnnB7HK
NgyguViS5b/qJ5kxB4RPBmLozKt7AyEOsM+T7lp9xMsmqOS671s7sXhOjJ7sx/zP
p85x6msJl76xf4CHxQJDyrmJaAszsGEl8MxLswDTvQ9N0N5qlGk13LuXIRfTElwQ
Yl/aDEkStIWepDXRIzBoDJzrCmiCkzSk7xnxlfGYJftADfKyjhlmjneTlPSttm8D
WLtRkvkJRPLVknJ5tFTnw2HMJxQlSRkuLmKpqEcS0BQGhUEIm00wII5WtH9XcSQF
QRAI5+BMpws7qgf1krhLMJvx+HnilRBrueySrfM6upc/CcqO2VrnAQIgE9ap1RRd
Qp09wtuEd5rFHuaUHLE1m0rwsGW5u40gKdwuh5rUkRwFw94ZfXN6gWcTmSBR5Pnr
z0NXQWu+0iEmCwakPwfj9UANbvpu9mIMeefKPfRi6r1pDU/t7RRsj1JZJUsmpygH
GAoj7BiVlKJ8dd5kXZNft4tlhLF4yQpA05uFnzomD195j7YE3QgCK8dcC07EbVPH
2FveAt8TAtTYVOyLatuMcc2PR944LjIBm3dFQktLSL6okfs9Zcuk+y1oIo7bGmID
BjJp2JV6Y5OhkEDbqQdo41eb+3f6CU9e/Ep9+nAMZ51IwWZ0XRM2r18NR20p6WEB
17j4IwyjeFuxBjDUB12CDe/xwSNzdm4JFTsrOtZRjHBmnDHoTkkBAK9KcRFXjljN
lL0bcd/BUBf/Y/bs1GafTmDWel6Ri5CVLSnivfRprYuBuNA891zuIIqzGJZXg+HW
EhzSfRqw1bgFPFthgKKGJOWL+a922ZHoBDV0bXoBxLAUe2WCZoJvODAgFYTTLH2/
efAMrkwrGcqbMWroDAvi4YcPOpFQ+lBghMcuh2IAnsqpuxaG/D/wnPYdQCR49N1X
9PkR3AQSh5hHCIaAma9eL1mwhNBOqKa4BiLCX8MO5DHV3Nm0y92biDYnnmiGTDao
jRBc62hyH+f25kJJlp0gFPHHFaoRcWn6cXhEGbCzCnbuoqeFtacIM+Sr92vtk4pp
U1g9Dga6rLvY88XgVZfKXP5BYjTCdtiDKBlj4FfpNI+RqQIb40f47rWrT++qpo5T
Yem7L931+xW65mcCKnI4DfFChl17JS2gyFWN0ilxX2YZ03rXFjdVCTivZ9GVd93p
eRjVAYQ6P6XHXjiOiFvX93qEOOwJd7ZcTQYTq1Aof0Piyn6WxCWv4MxTxfIIP2jV
9mvdO+TB6zL3jci9lfAooNVm3XACSxV127b+cj3lEb0Upu9F4I8zh/t0ojihhmEN
IkhDqls674dq4A6JgNZCYh9+WQ+z1A1WnWp71KScHiVpvNYvo80EGULqYRPIt36W
Cq1hFp9mzWmylTYEvgAvetigbCVst+v/51YzI6AuEuppoPVbQ7r/ehBJS+n0MD5R
lpOVf/wyKG4/4GINyChjz3n4w0pSnwKeQbnSkTGUiabz6TmdGhVbY4/ba9IqnpHc
k/kdYx3hP5JyfHiARWFZqk8BBTDUS5E8Mcu0IHceKI1qrBG3IxxClrBeBTrd6oFn
AJSM8K6akHp7rrFkdcYJDhmbgXx6oGuN166vAlW4VmVz5EEM8H0TWP4W/EkJOQPC
QowskHWJZ2kbPsD1LZbqXkvCqLOgLjZakCdfXJG3JakWBRwjkJwmy0AiV35xKXU4
H90LeqCR7PazpN8DL8i1Gpaad3hOkDPxn+OV1/uZJwNrrCyTGHekTwmw0oEWJkTL
SXh4KmOXtJ67Ey77pAc6twqdepdnZWMWdM+y1ejMxoRXo6i2QRTlWhgx1D3JKpZz
Igw1+xpIiN7uflcWddF9QDHuWf+KNA30wTM1vXxBL/Q21TbaiVHNS5oGimR7ZQF/
SjwpngBJlx32/KiTp1FGHbKutgu11UHian0HBON+CeQ0bZTkp1IJP98gKkcGUlYC
62H//FJqSCgpP97flJCa7YeDcr+u2xl9KJyGI4uQ7alRYwiTLtvAe2Imyx3athoD
IC9STTy7ZxQw1JvtppxUOVNwhKJupsGXuPu1LsPfVH7TZDLdNOCczuOPO4bhwlsx
vKXF//holt5Xb79drd/QKjJExCZO/QGCwzLuqXm32A9kkF1CeXlAeQQTNhNQ15t+
w+JkWx+vxncftDAdpau1OXfbvrWqJr8gnhT/Rm6TpE9N/YkCUJGiUWZq1RPrzNdF
P+lb8ggNofAGpIXijNhQ7NfR4atfZTskQ8grDfJ6DLC6yXCyik8CfPJ4myVE7TdC
O6fvORzdjS0KXdF1d0vHBFmLJo2Foh7D0rN5BDcWzMbagRBE+ClYs+qJSAQf4ESE
DoL0kTQnIP2rSGWsIu7lmFhXtO4K6vq+SdRZUMe+x0ZwxalVNfheVRJB+VPamHca
P67hM/s56RuGdzHCdwoc2yRgMglmbZJJAhRF3sZQ6807pazK+TgXXMQMRChqkoB/
o7nOOXMriq8HMvPRdbG1icsDQtJi3dC8s9yH0adar2Ht6T2QqAQhnO2sI9N1NfK2
8o+h1nodvdGMRxTOWRw31H2LR39O6drqUEGiyBsF+lDlXEOYM7+6HlbRLASLTYEy
ouZjE4yugstpxKwp1gDKrTLMakhijkeA2URHx2HaZKvmepCH16MXU6VRcuFzfV2+
HKYYN+TeHpHF41RcCPC1ldspNX3rHXmwDzfRiGixLFnxSVfzqixoGwVve+4SClwp
JUTId2D+cThRkKmev5u4+tmcVUWeVuUjTLbNiKCxs3JuEn1B9SB+i//PcjpQTB+n
YueG05dfi9nBYW4g/orfELv+vGkS/5cn0QM5biknRHxIYBbDGAOg30FiggNZmF2Q
GmMYhNYSwet1vsI5sAWtpfuv1sb1z/M1+6tk2nMqanwvMst63hOSQ6CQychKP8Ab
Pi2CTHTETz1QDZhSPokaeE1qylhBHSxth3QqDVJm1gFnsXgbN8i/Z/EzJmlUSmz5
63FJMmkwSMv2K42HyPJXAlsCmxd+SlA2/Ztr7DRGzk0H1Ho4Q4ORJ1oz9WO/t/CJ
8MCwGgH6NJUJymEkeJUeGyNu56ehd4AGumcM0u3RYCnSE664mo8IiqUd9NNkm+eB
5Te4Eo74p+UgpczXyaPyPsIIXXdd3r/opo6T/kPDbjdKyPOO17trLT391wuDSxks
7HHkdcEDWa5M1iu3Z3hMkr/8+JRHWV/tUQu3SS7whgJYOO9k1OdIQ9V3+6LUtBYP
1J1ybrJyKpOW1kaIvGQno0VQQ8fUGwrpQIUL4OIXt/HxA+AXyJbni6uZXYpJCV5u
m6ItvUKfLjfVsj+/BMpjthmceGi9ku/XlpC1qTsZBpJpSsZTQZib98i56kN+g5mL
Ws7MGo/Yep0Nh4XFx8E5KDp+f8EZllLw7yz1aN0zzoETSpJtqPv+R/t+A2+OBGMo
39x/alj7pi5+2crQYl15tVNrOa/r62bXqEQU5xWOBEHcWYEvVv94c9JcDDYtY/hx
9R2gCT1mwNAy5L/g8vvPNx4HZuWGX5m5NhID/IdU9UWg5czr4Xq4r1mIcq+zmIJn
YPv+eXhQlrCC0ZGUax1Q6XNRVMX3jKQ/ECfmqik0gaJDBv0GC8IHYqrTBoEp9CfJ
Tnnn2s3jz21tNs3XQZo35Dy9hdEI10+oT99KjWjRn6qxMerbKk8jkxxd9S7Yrzzl
odH4VZlBhE7z0+eFdxbD+tobZhDS4M8VxbljZXUxjT0mDz31314PJgCo/C9Bx1oi
yTOH76PyE7c3rW4IlrJ3S1wYBB/6Nxg6uuM7Kqjr4qmDB5R06EX66B399NpsmJOW
rFGSbBfKRkWWmK0T9Ou0J1i1C6tJdhs1xkf6HhauAZM1vJkk5SDsDp/6FImQvgOX
A+3XKDaaYRXtELad1B8vhuokv1M8mHwT9Rp6BruOQWKGckemzZV+tjpPcmc2RsgC
755Xz1R8uSRt5j466PJ56z2JrvlrOhze4yt+PHxKLPXLtVXH5X1r8aZAn8Z7aAF8
6wniedz+9DAMH2O+RqJO5cY73R51aWmeUDMQhiMaE8A3pviOPcDiOb6HQbvnVrAD
KHPBZOT9rmp7CblAG5LxVhT0G6QxnBWswYifBYVABf/aKhL6wysiity33y0YowAr
701DaLu085CLGtN4WnoHAvTgJQI1hSRGwm4a9zLiHf6nQrzBeu8ryK2ttL0H0FDq
f0Ti65aMRcutfYUqyfJ4fgny8s8AskIR2+puSMHVm2HmJNh/5cPZDtaWkn3uIRZF
sWFSwYbi9Oqv7RK6JjGpf5ePFe8BmzV1OS40+jReCsAATYdNn8x2OLFELDhsLzPO
/xJ0bd2cJ3XF3PR2lFeMHOljJEsFNXyKED2s0ZX8+p/bTwIZZOkApX7Okc8XbE3q
rE8Ab4rxcz8RMO5RgDxdVIkFzNFgVG3IoQrVtN0vJiFh/LWWmkTPsiRFgN5YP3Is
gnUObRMnzYxtxr7COBck8D2w9fpgA0gJFW1B4B65lFjpambp4WoQukAQBeZXC684
3H+9CJZGLkd/0RwdoHfOtV6aygmv87e3jdqoPSzvonpC8SeEdl6gR0XXdFZapo8I
TeyHQLZe0clerwJIJGG5ZDuFAkmt1BON8KiHx5BqUMTG9WKWQfBYqOvl8CEuGrmD
K87buqehdjZ8Jk/X2BZqfvSCaQwXzAUwUqYCbUX4/9PgkycQ67zrE9gofq5XNC1x
r0Aw0RX0oH0PDVO0JnFR5GTUUvQzw3y1QVfH6AJtNjSOLqZ4mh1gqUD8WA7Wo2LO
EUmM8Tg8YNz9LDL1r3dmVKRnl12c2sBdIzrvnKgZhJ2XEPY8OwyceC98aHwJ/Rib
2522N7TTr+9TB6r0ONqiUqpponQhFXTMHUx7xBFZEV11A1Z2Fm91Gw59WNFiyKPq
D+/2XTN8K1bJcyRFOO5r7E+bPw13j8F27L6AczhFdF60t0fSg0VNXEfomXqf2j6j
WIF8cUU0rnz1i/nCHhnswBgY5PCuDhl/D/OBXpBaJPE+cPZpwaPKnITFgMtx1Hlv
3FFYwL/43ouT0ewNjRuotqzgCr9SCeXGX0NbEu+xy2k4iW9yf5z3lgtCdNnk9q4Q
YujPiCW3NX7umpH1vDI8Js7YPg3jclX9Vx+DW2u4klQdq4JR84qCczXmZa/r2/y4
W46ko5b9cqYBLCmC61KTTPn84vYgHUj6bg7QNgVZal6flHYlF6mriMFUbmq3oiT+
k+pSwlhkIsSrAcYUdj7MQ/tTFhgU3LKHFp2FCcQIlqUW4VHESrvHYyvHfris87f5
GDMKP2IYsZ81UXbxuFpUCpkAJwWchoSZfyhy1vqIzyDaj35sLO/DEu2jaae7M84T
kNM08EW+w2y23VJiGQhjPR7P1e5+jssU0IfxN/R7/AYjGTrgQ8NZxS5Jrakb1SL7
V5zQm/DvimkaN9md4Ku/rhDb2xF/sph9xd8lwuC5vfbypJfoclCUCiLfUmU3o6gj
CFH39tdxSr0JN5kw1vrB1HhOIugmsursSCC3TFjN6q1G64jkdjU+f8OEXPxwv+5M
I4PNG1JnjzdXmloedD9iqWXy+lV6bfCCkY+MrejGB4zBbnrrlrcbjpi91YJHmT2d
kPWoPYtESn4V7OsBfKShqZUFo28SZ8vw8vc4f3Fl420s8dM3aWOh+eegVjdmFfzS
4rE0CdFmsKdmpeAXJ2vg9xMQTGraIeuB4ANlAQA9tgCM7aoUxhy4tpV1KPQWSZza
m76WPMFfOVBd7+Cojpjy38MYyzcZwkY0XZ7/pb3Wo8uWdLWw8A+DzAObDgJ4lh3r
WUUzirQ5FEsuzWA+Vevk4wMd9WTHmgHS6Mq//TmrvAiG1Us86/PrA7/FCIZaSdxi
iZZh6PJJtC3CV/RSoBQAejJAwL4p3xefRbPVHBHqaPsL7JYCqMHNyR79CMrpjfCL
3u5cm221RDRKNrnpE86QlOGfKP3CERkkdThWK7U2D6wzGwJuHWUsiW08Ir/8Ezv4
2uxqWtuFqgB528TPuxk0NFG14LpF/hu0ue4+lgVjxfbhW6ReRFuTQXpsVOcS5QbW
A9AD+0piqHm1IXwTMjhXvzgxOjVt1+kCqG0CRO4bEw8jbPseJ71f5HTktQ+fbIeZ
WKqp9cC/CSchHMSS/6duegikU2WdRNpg/SmXGb1SQ1aeRQtUhTnhnJ+uAlYzsa5H
E7y7b+QDNzPN82Nb/1VeHKkEKWG1+xF7WMZNs+a5uN9A9U8Cc2GBabsSjXz/KOs/
9advfB2g4t0tSdnfK3/+TILeOEajIcD/8u41IAVcIutAfu+jgBK/9tuscs1ZQaQt
QsUXTofAKmbKvyCk5UhgH4u8yyXNO7RieSBUwhXZqEWxd55cDUSrq0i1+FVz8ZNY
aodHGRzBsussA0UILjsHzSTZ08ZqrC2fs8Of/hVRxpgrmysYUkrd77FLQe3xXZeC
eRJzKZIWXVBeFLw2YVXUTKMC8uvahfi5x7ueml1ZYJpWArJcTQlxg5DMUCqQUzmi
VeklRU3SCUT02trTxtQiU0My8LdpUba2ihO6Psd4Ijco/vWkP5379pACS6cjWMVi
sSFaWS4Yg+fXLfu2KCGmnvwpR7hzQnaCw9c+dfHzrzl6eHm2vzAxfzv9kbSEZu7t
w0xRhC8TI8BGhsaRt6iWe31oELMIoKdHB4eGRLKhuBaod6IyGSPNpWcS/Y8Ua5Bk
OMKq7RIAM+Yj2izxBbM6i/lA+/hEA8KhpkLCy1PmY2bh1tqNE222Uo7s7PiYjSer
9CP5TY/MbIDDbIHl0jwRkgMLNQfN1uPpnYUjEtPWGTqf6//xzlmR6C73h2bDqPHt
enHMPBJst0Ml2mOOWTFT571sR0gweY3uhWTrKVMCm6dyaUMxaWcn0/lgBKXp5Jqk
qf6CVCGTHmbbvPQKkoxFJ5j8dFgt9yjIZbZ2Oloz/TqPiIbpDAfcliijtT3tvM+F
O4LlCWadDEAQ5EgKA1z88yrYaqD7vGwsi6SwHfVZX5a5Is8IFO8pFLQJqKioIHt+
NeBa9JoJU8BiWahCuIAtYteEzj6Cwjvkt5hP7ozQh0Wtr7tIOXuXsy9+6T0+Iwq7
yMa50CazpZdlbAKOdVlogZSmrAYeez4GyTlLkpC7YJA0LrIDrGMPFI2iybsLP6xC
43s/y8l83m68YNgCW2OKbFLofcNkM0L1ZDELfGTCUvhy6ivFmcdquuWqBhRJw7k5
r9NmugwIEHirKMcW8NEMcFencBc0EAE71AArcrow5CyGDXYC2AsZoWsQYSYreCu7
b2dA++8NKOg015KpEH2t5PT7Z/OYcxTBlUYJig9FRmLZbxQjq3w3E9u83jGo3aXO
5Px3REAzsCZgbzJCVbisXk+zo2o59LHjyHmKaHd+FQaUcC1PUwaqt4SHU7wL7FFl
cdMQBb33recXjqdAn3S7pnCpyrqlTDd6L7bpZpMFBwqMdzagsLaffavKMOifwHaS
+icfHDrCOJzelIRXG7LJr16z9JOugRhXOhI0Jfh3Py5XO3fBTucY2EOfd3wu1C80
IJwMChnXK5T9no82VYZ/NBeW0FEMfU4BCK+wEwuI0pkeEsak+9BvwvBkIIgRGiSJ
2uPRmhuFiCI0/gxi/x36LVvircX5qSuh95zgu2fijMRSD2iV6QTzA4mNPgKwEPLQ
X8K+VTDX2IMsjOGcFS8rH+IlmhOFjy+675IPryZHiqMqq1MIwbuUjYdqZw8jgDL6
kqHRJRwhMlroolQJwLbAvvsabkpFav0kL7VE1VQbKcvzm+P/V+6Q03KXGJ54fAfV
O/JRg1TQ/75VhkA9dkDtF5IcJxun18ls6wEDujm5NDydxx9LNqv2BkFsIT3G7pmf
IJK5tpl+nuIz4SEABdAVL1foluVstpuw1aOZO8EWgN3ortFRni+zhcSP7+SIQwVn
lin5/6h07gUVF7lURBU9XzbWLsiJjYsOg0Fu7sORGWmPDLafT5qoZjB7jMj049pQ
q8cQoxh0QaywqOVxn/93V0DA/PoXqu8KTNgD77FJc55I5n+Bs3Mg6gspr0EjYpHr
rfYK6t1SKc8aEq9SAfta3gGa678sZD9KMMp5lkXtnJMU3Edp76FbkMDWHTrZASUX
YAzvGY/XG/iJmlO8cBFrk6V8cF/kLsT80uHD0R5Yp630V8sOOkbvDHivhncD4GHE
hTNscJbyIS7AAMpBG8rV8hdqJK/HCWT0ohghJ5948XSHy7UqlH+5yGSp8DwthQcf
G5gfW62cHJHr12f9/9gqzhj+YLLSv6DZRkyfdiYErbjc5h0q+BlYyMhlEx6b9iz5
sd8sQidguXHjPH5C5Z/tjwblx96gBjFvKuYq7EYig5vhzlQbSnk5ACsGjmKm/XJw
G4I8PC5/gY/Z/fcijg/yW8BuZesCiN229lJ2XcsIeaNnEXrZaSYcNiX6sdzgLDsR
2GcjsNr7HQ6G6zRXnbSvw9XT/CBgh03sEHEy5vjbGCV1MiHcZx8FrWTWY8jhuWRK
Tbl/qT971wLXCBf89cKHGDlYUBsYPqCCAxjtJLHyrI2r8CI1D0JjoCR82cluzo8s
eVhgbovMIEKE/VxwMHcxBIXYaKOEh/IjapZEQDwUD2djCmI7i16PbxOeLtx8IQBi
VjEAGhtLB01GedllbotrJlj8pDKVC5lrXLUL7gbiMoLEN0A+I6SZqLms3BwVVf1C
l6DQdjzif6L4iWPSs+VbIK1ZOytntzjbg17GIRsm5d3AOfdvxeJd9r1GMSTeyRlt
zgTM38q5I69u/crdntZBQN6E6anZRvvOZzIe4MXHaaushvSO7McI/6Bp3FAaq2kD
qX1SiE6LWtXouH8pqeisCDTcucz2/4Hcz3ewEw+GiSMMeT1qQy2gsPkxw5zpKWjE
+f5cwN+JBnhSgYyaQqByCrONON/2+KV8LCknYMf4jVOa6dEKHJ2gsw74YGsJxAFm
IJtNlWdfl3Z8YNWH1wtfrcGe6P1TbontbKyP3knkPpRwJiSTWqT5JJB2c7WEHy/f
UQxuMhswQ/MBXsg2q2P9LDwOqin3I4kk9tjkXFv6bZke2BLcsOV/VuTvBCx+MATw
BS8VjIb0ZsCx9Ihe4h0ANQSs9XWUDPyu+RofT1weIAKKenM5Sq85XO4BM1zWFJwk
DrcUg8mwWKKVUcUd+fKu0bq2/jbIw6LLsKlz2cjQWE+4zOyW0kxnuB2vIMhlIJFY
JTSX3RcCHTQR9U+A8ZOOeYfdBwT6GcuXX3YUjR7ydAwkQVnRUWk4wo15QCpV2uS4
DLA9QjaILqPFUW+jcnLBhhemMAYpc5Jw2rzD+sVvI6kMOvP9c9LMS9FcuKJgGMvH
eoJJbNzPQ1lbu3u2XMUM62kiA+orAzON+iJjZnf4/Z8CTrT2mdaQQFwA4NHmV6NA
7tOl1gYpL33x/2oh2c3rT+jcFpIuz2qfCZF/3z4yB61E7TBkTxEip8Yi6ktsKyMh
sNpINL/gOUjOb/Ew3ZZ8y4BAjC2TuGhp2viF/ENl25TW6p5HS1BdcnyiqSUtMHNR
zlsYluoWCIHpmORrDAosMfRiKBixK/FCzO4jlwz1fAuY2C9LMgBSNi7CLKi8Q9Q+
CcjV7wByDKP28f7rh/PPE2ouX79855AnQo3dfzOnBfHw27VQ3R3eFUNeYAOmt05o
ydB74s88iUPDY1SPv8jHhpWgOEzT32G2JYYRpGvKsUk+ngMwOxZy7eWcR+UNrr9T
SB2LXEQU9CkcS6iWDLmk79vHq/cltWltlOl4y62EoYSGIua6vq9/WG/bs8nuObcU
T/B0mQCw5AlOGeKoTUDhaFGMxAhyqVr8s0p48EqarUeYkfVxsojC/q3k9Wb5bZhs
ojjIxAbDtVjdGVqeTvWwjVYv8XNkhNnDeQKpkbnUA9zC5NtbyviyE7VR/GfYf/3u
5dMIk+JiIucD59EE6VTt1v+u35BVe2eRa8nVPpYfbFykOwNmq1dLULsX63Y64b8p
WIlZY4j/FYRzTDO401Urml9eK5u6L7NI+xsSZ2SmKU4CyPoFATTRvef0Z4Rw+BzB
7r/ssKJlwxPWX7D//h34i+0mVJ+vJTBbikUSyklq4ScY6g0U7e+VOxpzXisc8f0u
j29P8f/2YJRnlOQlbqvOv6N/MUwEOHN/D4TjhjuoMtxEISeH8B8Zbz7DKEzlDu9U
XvJfhpM6Egw5NjehcTz0Gsh2OE533lMNOZ6z5bsvwME17JRUZbMYyAppRbhxoO1F
GXPWGzskosjwknTcHlzw7puZkv3xK3zwaVkVN26yItMy/0ZhwTPT8/zegPnoxsT3
/8FKChvu15cZoJQPrWPAfwCjjbHATBVJnJqRMB3jWUw8b04E6kFGg8DClO3/IBIl
YenAzf+dxkiI4k0VXanFx6udGtiQI0Dm7kQgdMdBhoihVkrlfXpPuGnW8evsgyYR
hy6wtDfAUZ0USqp41FBlk5iasZRttD9x/3doGypABmCq3HjqJUWVhGkxgjVgrHcO
yKHpTCpuAbe3MHH/qvxln7ABccUPpaDPtOebt2DKo/NjkmMxxgKz7/mkoY8XpOsk
U/wXIh0yRe66ht6RluPcYuY8S6HEhethyraikx0Nn93CorIQ5APhEb54J8bY2NVq
czS+1r9z7ys2f6gO36IlfLGE8wyhWU61Gt3VeJa4qCVDD7N67AFD7LeRV96FIdt/
UDSseceQVXolpfsOuKAmnsjLQWcPZLDR/5IXKQCYb++3b74zgFcg3gqq+LsMF5ca
NRCeBfqiH3+HJ7T62l9aCsUhPe4FVbwmKfeHwfd6ZLEJ3t7YuE7s2RqRVSctA5g9
MYzBa0R4arIn3HpnJySlDbbXDifwPIgNmskxAfNXq8kShhl0j3xk4AhSscZvwLth
1+UpU131SRr8bcyyLwTp9eVh3LK6MTg0IG1knsyAXd8CaYz/LSAdAUseio6jMGSt
XuwVyZu1S4ptAkoc56InTS9g5x+JGekRNGtDdTyqftDOlJOsPR4h9GFlOQpg41LK
saLca0aFYB9rzO1SIFMMpiC3n20wipGpGyQ10GI05YnlHVpB2NhLAVtOWbS1lWUf
QmM9Db1xZ+cuOcgxDGJhFo2IJdhkvMCrD8xbkKR2OM4zt9tYhLV447MSRi+H7ptY
0sEhzTI3xRmnrYvceRYFZn59QZ7spYwrgI9TsjV6/Mu4kM/Wm1zyvCYZ0McySIOJ
cBLXfqwlrNkBkG4CvdV+Pz4TOFv42L3wr/Ipv+Gv8dp9oAvW/PYPskp4UAqc9lXL
I1K7V0FfFZfGkJUG3JSYdTAt115hfVC7zDnHVBgg3QGWl+gV5ni1SxpEjolbtAeM
UwrJBFT/zsqW35SrKHRBhQ8PgPisP8TiUfhb5NvhC3Z1KGIzuGWSHFSqqEsPv8aX
NHqveqqCWtsoYUdXX6V33OrqQwPGJ/ip4CjZhv9Xo9JtMsDU9nptSV4p/vy4zye/
/9orWwENl0RkTAln0hLOAoe8V/Fxidp7vKfS/Ilt1AGmRbcaHgrGukRBtu9pjIFZ
7AOfjPwaNU3JB4yFmGpj+ZOuxLWvZ3flQi/DGHGfGNbk0K8SBrb6GVu8Sbt40l1F
nSX3qPJwswsXsCFOWD7jLXMKSvIHQ1u0z1349rDtNxc46tbG636q4wEhYULA/eoV
20Ww0+ZV2pdTFIPSmdlvbkPfDm/mZQyZU4oc63dmPC7WFUvDGc4luHYMw/KKOjzz
ksqeFjytk9wYrL3rJB5qVUlpNi8Y4Iyv2WuRwmUJGMvF5A8AfeAIOSRZWga65IvK
eFQgzsqEH92allTXdUQfGThPAM6gz8M/ABzdKjDcichWyrbJsv5tuhN2nkMrOo8i
6B+Us+lm+4R5u0J3wy5J1Im+DYpuLvh2jcwchsA8QG62sSh6039izkmYTeckRE4a
QbZ8IqPmW+AwG2Ntm9S0YBmUYEnu/4R12nnYAUhXcjIJ8szFMMuk/9UdH2EDcjym
pjsGFtEWlTglPcNrfCA8I0mOPZGx+qUHRUDDj5mBf0GTQOG2DbrdA4/XMVPhP9Um
va1ZzYnx13DhxDdicLKDoSpi/a/JEoLjXYdP+qTN7unzMcEPjlZdpEX8MhE8LuUd
q07K0m3iddLt5wdKM507SyJuWBtgq6ZP7ugWIxsoZUoB+n9on5clSO3Uc1Z23xyN
DgBRWm6Wy4JTFKdioPATiUnc8gduOGRDG3/iTTpPXiGZlCh3Hekz41DipVqHFqEf
cjAz29Fyn2FW38weOLV4sKNSL8xVYG2fdABlP/5gwFS8MHoTUnQBsKfIRDJ5Wb5O
FZZQImTX+fCOCHDMWKocAH/dk23oB7MdUK9S+42q8aC/UJOgZnm7/DpfvjjkUjNg
I/e2y9IcoLdg5lthCJEf/oVCKSyo9oIcd8SFOfvY+6hbXB0Ey41fDsfeVaZDhHEE
4VX/2gjn7RxDr77jXJ4aubue10K0/4oWR5ggYoZlakeUD48/BUPtOa8mBYcDRu0B
X2/dpKiLi5Uz/Fv8AsR2x/5n4C5+4wRewr+49zKgNAKNAD01HY5FSirUjEQCrI7C
gipZmaPKgJvHXjfK/xDaqHMbzGAnEn/tn8NOjL7Yq0ZxCJs2hif11FS1mB8wghTG
aXsRzLArFoUyfMfw9VjWi4sjtI855I8XkXCXhJSw2rsN764TeBbQoTZ5aL+aGueB
cwcaC/GSZuq7dZi5ywy7BQD0vZChx+IqwB7DUYhR7nsEBYvwP3RwYUinjY5ABPaV
dmQIyV5LDZlk0GwMT/09lEBhUIJFyNnZ7VpJ20rSmuBawHxQxaR4Y4jQZmnxa+gD
D7JV7VFNQZN1OVuMabhLVVrofs0R1ps5qZt7OCsde1cqde/37WX7z+65UmUreicQ
NltAKvAMw2L5gpLQTQq8L90JS9adMUtfcH0GtD4UCVrvoHloewKWO7BicUEBe4LF
SB+7ICoqKgTc4J0nSR6Lyl57RaX4x4izKGNr/RD7nRhJ3skzDldAMXrCE0dAaIBs
DytldFJYulaGHboNqfBuRh18wJ7p7u3WWdrZeUgJZyko7KdQz2pNZEM1pzxXmn5r
SXgAKT1K917WY4I4xy5NcVpIzo5oK3gKRqEZ2YSG77VPU7qDBU/DegZjTL2BkxeK
Ee2oGzHvwZQiH3PTzMoJ1+W4lETJ8dlSVPgOICNazvIow6TuvYuEkI4lIh3c25G9
RmAwtjMDN8pQKspr97+ybfPy/lzD6uX7BRqNkY6GixU36ps1IYDxlinXWDw+kkUI
f6kZV8MtGdGFGjbFKUaMA8p3bXrXcwa7Czr0N7Q2JyziKEsMTN3RM08UBoR3WNvv
1kU5V31oLdCDuA0rhXz74qOxkxBzd0ZfM7L0mAuCC9N72lx2V7QvQLP8LTJ25Fod
fh0f1+XcOikdOT+RcKKcm3k+V6jhvX42+A9M6tzIApMU0/5O0EkapUBtlnVGnxch
XGZheIKF/GOzdL5p6WErtClJhJcQory4ppAw+A+RkppfGhbcAY6nYL9dnhaNRstE
5lb5Uy8VHSpB/+7gsaRO67qCyaMrU/pSzGXSVS0iGKqyakdtXBdwM1fbcXERDNIv
cTfLj0if1LExHnNTMV2OiFgRhPXZgCqzGV4IUfUnk+lVmVPWyshHYMS+/0U25e3i
9XgELZEDLNv9y6lH315u+4gOvpPnaIJf4XAuRe7j2LaPjSsfvnmk83LAMO+RLs5Y
XNhMFBqJJ5GQNrCvicmXAXuQ1V6/kgrFhmF37mdeUAmQEJf+0JAFq1xYuBCYiVxi
Fy9AfhhMcM7Cdh2gUJpvrv2ZPfeWg9tZ0SZXC67285j1Kty2fYefS2gqBcpi5Ypx
eo5A4rdPhCpEG7l9xC6MvCPbhZsqH0clLmtdsqton38VhE/X/zBRI6FVzHE5XJ3O
LRKorXlnQUtiA3rX+GoF0+l5NgLsNyDXuJfSvXjiu8t5xspL7I7eow68HtPJOSo9
+wSYqtUqgyFcvjO9dv591roQ2QsiTuX8rISaZazgH9dLPI48SdwvA0NPXkCdrsL8
sAUtzJ1MaE3kmqwiqPhog5zUxFf4IpBEYGoKh8DejPvrvqvGNXpNzo6tRkgkCsrD
9asW/6RQOjOziSDV2W1j5droFqOUzNeWitaeT5AaVeisOWm5lS5x9dmTl/u2L941
82RsreZQ+1SfeupsyTYpTp3eOoth1RX607WCbPlB0mIhnjbf6cnu1nMPyupic5xN
mjwfYBcyJ+lf3vEbdXMhYjoXoUWqqgjmTtShguJN19Vjk0doOKrAzQsPGd1M/Mlk
95ZqT7qrd31RoGzOfPuSrmwufHTqa/EfbHGFg5vFFyySzJhgvVgzCoBv7GlWYiNI
8axqLlYyPxQARvujmB+duVdXvVBXJju+fXMCegGD03iFQJ1/B4RY/SdNVyAAtB4U
leMRUvsrB1bGoFVjntNx81XmAIvCqVxJCQKSOsxLRNdeLSqQx48wTH7tFlN0j55j
1Vwza2SeZRcO4iKB2uHsj8Rdcsfr/WW466fFTUx1K6qQwRlbHjf9fidAfh8J+Jb7
j8/5ztKTwrGBPadnZX21pV0Ek+TjCPyS3zD44RLDpZweQXyay4YPonzeHag7cp63
8stv3rBeWzye1Rfe8xwZeMo/kug9vjmKieo2KFng9ddr8c1980feAvi4BAV9r1fR
5VcaqA1xFRYtKycJfphPlzAGJp+3NgabyzKOlcYCnajuRltjTvGJeeoYneAQqyxk
AfFE/Wi/ZKWtd6v3StOuBJw5J7PTXhB41N7RbEjy57hadcYHdfJoa3IyaeinBd9l
H8+Mie1QVKOUFVZ3QXRFH0XvMGoEep1IUUlXuc/hjI+FQNR+oXRanTqaFyT3817t
u5sP7IFUICrr207laN1EkVCvcRhL9h42GysBCNpW1gyN8S4gFquKXloZ++H4/BDL
DBsihUccPkC7urCJaIKhVlEcPSB6bkzs3+gc3+8h+TKHqjPMBxOByyqnz7gyZnqV
wPTH7DB5Lc/WpHWpm5GQVjtiSSuEGvHdak862b/OmfMARiaiPmv5xO3nc3+2FEL+
7e0YspxCr57f3TJa+4S/QAiAwyt1FU7hbd0to2XGIEbGWx9d044gM1GltZIivJIX
oyKc0cxgEH1e7EJlJt1zLfH2ir7QiLipwYi7sgSAnCgxHRfQSq4T3R6oesGoq72A
hKY8ATH/refOD2zSDIiYw8ONSemuhvB0wWT/M+eim+O04Q2ixbMtHceQKO4LyEVb
8IJ3r8wiIvnerLXD2SBh1kNQaQXQ33hWy83W4LTzf111lo7Lx983vsRGHrU5fQoe
rDolKZlaXJTOWtrIYuZhye6AvXi6cbXFlS0Q/w+wbnLY3yEMfQSrqcziMibGd4uv
mBeYJvecGcjpTJmvWt7XOBOuU4TG3DtuiM1FV5ZGdD/BWUGpFiPs0CeqK5JNqzi5
u0MJLggRx0yDJaXMaU9e60WAu/fPIEu5lA222alr29azbEq27UKtGT7EIfCQc4hs
PbQn1hu7NCs25JaNu/6lWh9iLj0+vE1w6ktVQ0y3zSD8MbyX2MvjyA6+CGDaLr3v
dhEy1EdUvUzirR+R1KdYxGbiZp3MlUbyvr17DP0CQNfIWy4JTQGCIcTtDZM8aGKO
EsAoMW87Yh3/9hFy8V15Qs32EMPvEaK1duqdtK6grReWBTnuMbH0GnGerPS/zCVB
Etb/ugsROL1w48wORnpJdqW2csgCuwu79VK9SzPOKhAFm0WzWBfXM4/Lzuzgfzma
exkWVVP1KGDlIN/YwqkBBVq8Gf0hyzIvnsL/wroURm0YW3iOdMi1DwhthofZ3QVv
YObZW+7TxZwOo/ngiPSHv8vS9WPGIOtJEEiNt3E7D+H6WoHLeRNG8xQI4GLkSn4q
Uyp9jF0/OkZxeVd6ueVPLo1lWS8NMJ3GvEgHpq0qpYfYGQb9ztE2IIGmjQqThR1V
HFHTFMs49JHDA3bygmGfY2AnZ60p8Ul2mgSUigvT6qRw3tJxQVpNJjJoykWSUcqO
Uekoz8kidk/K/xNuUBCDMWYXclEXMIpxT3A4Ou1U+6OpqEggkfKUng/1zgI4Hz/6
NtWb8FVP8kdaa+hT0gjp2i5f+MV2neyWHEpkPE3NflsKlZLcT++eJPrUGCoLr4Ao
1pRlJrItWto2xQ9XtFTzpJ++JWKDSiQuQQduJ/CmiCkOhjGcB/S2V3HSae2BWuFm
pkoXnQxRo1AQJSsOQFOoYkp7PgRq7Z8fiagdqP18dpZRAVAKf+n4DfpONO0D2tDc
5Z+PqV9b+PvLxQshum5VjPC61VThInbP9K5D5F0o718rhSNQKMMVFHkCmWRDNYFl
Egar0S6134xTz/KkEWGxEYaiXzeQdO1nkoBtxfp/Pj5QAVKPse+lrEbR+Nn/jLAy
BvdJ7dqPH18eHJ+ohberQjl6MYAZep8rdf9XJgFxJfAjoKKmvqYqqGbsWClzpzgv
Y4CaRMOdFJvr2w2EdrrcyN1orD6j3rHLHYYsj+YP4ctk1kUwMDrOuP4mvBSRWrai
NS+hbP9eGXJQYRGFCvvbSkmt6AA2xRce3nduh90KhrvOV6Ne5rcrh/iQc7Mxln7a
qOBYosEP3eW4LoAO8P0w2NDNb7WP5deTAXMo/Pi1A8pGFQC5+RKt/ngQ9AyBWU0L
R7nAG3wBpriz9bh33dCnryK/+4g+4vJlMYD2EpZMeJJgn/mIC1H9u2tWP7PQcORL
2B8G3kBQufOiIROA7TigLPY7o36UBuoK948ZAbzeHkOp8GTl7Hs56v09JJxg+BN5
covkipyoIKEgHj7kYQYv+5uIqxsNgwOeIbl7Y7l88/opoe6Zc/ZZINt/SOwoYtBm
stnTJrnGJzOoCeYYYx+y4+2ooQf39RXhf7REUD4ETqzmgAprjh2TxaNPCYbXcOKA
y6k+ERXhMJqPdzF/6b0AOZNd61lkRB52L+GAw2MQoG40yztR8nhQKTPFI4zqY9iL
YiOVWIQFAQMN5j7dcYBXqJ245cKdzNWmjD5ZgyU6MQNkoiYfMZZFIG6Y4B3P0GOT
y0WrL4Ip8DabNAXQo5xWpqx3DbgltS939jIqk56ji4dROMh1gcB60FiR56E3cGf6
NPsynmO162SDdPY8fanqYRmFQlyTSUZg4fq/FeMUPcWaRthdm0NeSshfTjr/GiIY
Na9GUVrtYJL3kcARsPY0tx2rcObiNRiLXzvglRiFvZHJi/KW3ObKZ8P3isnNHWg6
T/XwS9PcXYz04D1zb+scwzPufC6Czz7GZkGuBhG6ob8X5sup6f5LbP6yW0uMVXVx
UQZKQdiPxPkUdOp7lNGtg38fZdZYylqsfztx36ofSXQT4UHhIv2fKeq7RaKr599g
a7iikyN3xj92yxNVspMpexyDHuAyG/LGFPHgjVVjHajr5MiasiSfTjIUedN5y8eV
+g8zWluKMTzQ/GFORA3Qch0+XopCNP1Rg6RzQLQV5fppKFOuOndttSWajO44PJrw
td35MO6uQRCGBglQxR/Qjc0axzpHDBmNsvTmFiOf30jiHQ4pHj78SXRm3bHQij+Q
QCBkl28RpksXtAEjydn/B8ld1QsZ5Ng0P40P7CLwtLPaQwt9mStuuk53ylxxNU7s
3pq20nWuSIr9w39Ht4ilZ2WyVxVt/HR7IBPIAAkIvtfAAjexUswj8P3vlXrdiFho
TZ3JPXqXFFzNgbZ78hydjzabYaXmkQWpi2nnYetyuA3dzWyMAb0bJjusdn/1Q2qC
eegWf+5kb41/Qem4chSBHqylU6LIuadB2UMY0DhWHB6qAeYJjEIvexcT8KQkFzL6
0cFnvM14Y6r/WiF5IZ3LzJ3++OrfpsRv+Rk7DeXsmo0Y9KMLvaVJXkC6yeqf3mQ9
e8+h1h+R4WXqjmQzo1UVwrwWGjZ+F3e5KZa26aloxjOlxwhVphA7b2uygi/ZKk/3
omgp2XuAvqiaecS3VTvmJ+TUOXknA68iMd40rQKsdBfrNFZ5RrhWtrnv6sG8qrBr
vROTiFdcq7XZuz5pRk5aEd+9zE6HoVuJeYfStRWDwa/c7x/mLKPLQlUsVzF7PZKO
KoCdFHCDPNU74XrsfChFR4WXS5xqpNimf+e/TZi/2xNvcU2gToktQ7XgcaQYIRxa
e+XCokt1qEQc+Mrh+JJJeY+T1YYVzEGqg6Jo+jdTnFNTHNv5g2f84QHanZBAX8u/
src+IOqhbsiuTp8/17kZ70F0hxWmN9VIsMb+SyWMaMo4zCGfJ7AfdHlSEkNZBVcx
Y4SB7FrTYsoeL/emJHMten3UoKweuuAiWlMjqXQo1z9+IuTi8AN+bkieOyE7nVEp
bV2aqmPIIyiuLeOWA0M7vLiekUtHjDcr0vhGjxqfBCpg1AU0QqpKMjR48pTpQGdL
SVqJZJfMoJlvfKzrFzCiKFH2/Ei9YwLEHKh0ehCvkisDGDx21TUHR9UPnNEWyavw
zrvkmkGHMcoj+iSVhCwemr8hm8aeV76LwzUMQlj89QAfBDrYka1nYxmeOH6yiVAF
ZbpFRx5pB5+dYBBKmvKlBqFVc8IIdM6Jqw7dSjhySADwnpv8utTvabxE5QXaTo2D
9PtvvzaI04H88ZYEvPAb+cHyCf4OFdZ2Wsq4y9txTAqUCxTWE7GsxAs8aC54GKgB
vGyb/GZ6K5qylM+ufAqLKUPpqCoXeuy2cNh04Q+vYjshmGgn6GUtJlhGDPwesRMn
syZ3eeMyVOEpndzCtsa29aSeLhsOj4MQKt0tmywDcdnOENUVE9MlvMCIaZT9IvZL
essmoMhD13PSW+p+R3kdTHtv/S7DXoIqLKQJ3saYkA4lphn1rLcy3iCx9+o3zE9j
b7SGLmjeR0HXBx/vpw1JQq23aiJjccP/0764O2S0rvYqeTgVhZW1RguEW7hq0EC7
yTXX5Gc7ENXYVCrNe5LENmeUb4OqD2ddNnApDQQ5fgaN2fxVahyEQjbl5Vaiq7bW
H9+w9gnSdCE1M7wBAl5Q3IBba2VgdO7F31EwdYpmUHySB82OAylnWO3BDQfyKd1Z
J5na6Wbn8kmFbZRIWdnRwU2YDFMpShxbM15fkUqaNdTUVHMc3Q58rhyNtOMhffuy
wHWQ9cThoYKPpM+0Ao8vTPWMtv76ILwNbXo2yuKZaqJjAahMCF7svfLsNMPUtR95
BSyH4A5+U6mEQBXcBDVx3Rt8wBJXjLBNBMXdIQEewUcna64S1w4NX2u4NURRFXMf
3iYNJ26/ioEj0tFTQY3jNYT8z4NXa4t82iOmHMpu76E72nPE3qHExJlxstA0kM4n
DaojhaA0GTosh6gctrMxlSsjl/vn0+kaYpFiLTcj516n7W66zMKNQ/Q7ox97IlS3
335pMpFA5PMq6CIuVBqNL88jJyx++9aiPiRS8ZdowFB8Wd9xiWe7n2iEEUQwzKym
QB7C9Ems37u02Oe5ePFhOCZYy1XkeDd+5nnBSPNsv6OkTXnvNFW1Mztckw50kOQz
dxlOTcgW07+qbAMWmYqgQXXT9yZlqyXTQEFblAXvJie5UJ3Mb5JjTPE3Ow/ZLQCH
/eF7eed/3SrWh/0m3M5i1d8SvCsccGgkrCYnXBzN+yP/8G+WPVAjbscY5F5j4jGF
jrSkizidO8p7KFlWUjAtmmKIDy21vgJjLLO2reFUtSL+U2NLylrTOYu6tb/OhnEc
E8yOiCCcRCZX54lmnPdcPr95+BhKwd6P7wI0pFVAKLWUhFFBerF2KEmKJEzjZpnQ
wPGRRXECC+X7u1YmLPcnzt/ZU0iF0EcoO+5vjYPT/y8te9DL4zFYfE2/SJuiKBmJ
l/yqCtyk7VwNn0pvPrKr9BwIWRbQd0UBx30XUFH/auV4nwDDaYK8iVLiZCr1eBIF
ljmk65zjeiaAa5WL4tvkKk75Vy1P4ULMJPJhybuy8bkoxbfH6mKltJgbjEdD3osy
lysUHaED7J+U0iKDBHfE1NKc7QJ8AC7tVzoS7NEAwZrAldCgkC3WRQHwTxo3cONn
nuxzdXbbx70j46zCndjsiWrPEp7iXcpI48wgEQIs1TPGXenf9qYT+3MoWdVjKZsE
fsJLyJ88S4ZCpkmUHf2G3RoXXXy/TJHItBcmAjSmGW4E2+aVuX5ys8EykXNx4YBH
MuKYZvwr2LN+UV3mJTKu7V34n57b3z7mxvUWOFm45oHgZfioluu15Hn9RjBy+Fud
6NSQTmtBD1XWDE91fPqC9Luc2TAL8oaHQH79smnz2PQQYxXSx35b2DmGN7N3xpDn
MB43kk5dabXkTW2DY2kw2+6WnJT1NkMB/m+ODSXliwE/YM1rFE5hwgKBwIuXwS1Y
lxSlwFiE1QJV9/nZmHCDostBkT10+iiwratwFjwlCHZUU95K5mHg19891VAt8g+S
VChSMvsiSbi6ndg8PlmQlWu3e+NywLsTTR5U+/sOQ9YuHZJHf5V38HGBIhtYaxjb
8403UVuSYPBS3WzcqTeZYEtLFeziiklN5ucDd9JL/YumD0abhdIDYXeKybz2jjOS
oShwmo7Ydh9t4JIVfDQOsWauGt7AjtiW62+PANunWsmx53EWPs7GG49b7VwyiUvA
hXIeiTs+xmsKsbfMi5jDfujpUKOGoptnC4+6Y91WQoceHwV4qPNP6QWgOliqVpPC
Sukb+1iLjzKQmgw+BOKOHEgvKQ8xTxRuzVmE6ZYGH7nmjzFRn0g5e2ePSzf95RhT
rskMDMcxDjW4oVFE1O0QamNhV+Cf/Onu13yj0EtJz/bSbQx8Un7GG2M+Qm407o2s
LtlRUb4TVwdsMBULL95vVVLr8NqJ9FJvXEs0AmVzzl2pNklbNupJVwE+IOrVYu9x
eGlYpLamhdl4LBrjFPouoOlhFhWxOsuTZYBkmbzQtWnF7jmKBi/66FQcis8Aoiqg
skOqlOQYswqGIhGqpDWSwHjbCZykB8KMQBuh/q+sJTwhr1AEDFuO5VyZgz2LsAdD
2+7MjUdvnCs7oggSzE5iRPyG175IuV9AZvAmQkFGATJC9ZMo07ZhPay8AV8Q+SBT
KLxNEYQYHxiGNtHgA3/ZhNrcQl2X936PLx+Iwo55Na0avlyshVcMhHbEpOaUmSQP
CetabVDPQBO9HX2DtCLWBI88gRjTmIVjHL5pcJkLt1IrU3IstmRQVIr0UcfIs+/1
Ux+B4PclfudxXuXM9K8DXCjKKHAh9QOHNHcXmQZBF3ojBUWHPnftpPxConZRO4qw
VpBDwfkXaJpi4quDrHDOv1HUEwtOzD+1sgFt/88H92Uo2NW0sFE/O0RoTlFWPm7Y
u4yOhqj3w4FE3xHbDQhLcLvDKzxjWdNlEGBJCLI2W+O0+CGRTxiRqADguTAsIdOV
uccEWI/5+XwSk1+KB00rpMcETI1hSzUTj5pAf1Yf458R9tgBpNk2zUCQgpnHDe4D
VwxyNLEr+jfnqL6jJBhURYFrslJ96azsKpYk5WbsQFOMqUBA+zRE4L8CSzXCauF/
GCTdGpiqiHvOsfdZmehcvwSA6Zsoeovulmqyq19B0MHI2dFScM465HlRSKW2NoYd
TcsPsatiHlkEtY00g0mmbSkqkyKYaumP5lo+3a7vjaFbPkfN+lfudQT0AcJVoKkD
oAaKlMzImU+Pn6AuQ6XM5CO2cJwANiLOCnrR29zLD24tNwTM0TMAiVQYNPYZuTB/
eAkzPegkmoD5GVtCTN0oj6KHAOvGZssRYwB+juFjTA7J0AYOPOCNX5IObwiCx5yh
RzIAqcZcLhVdmMU4N6LZud7nVyVyq68+VT2YO3K6NhUrc+wk8JVHUY/RDWbTgK81
tvgI/yRF+75YYnoeXw2hyAdT/Ya4/yK///0rqxZpg9yxqJc2DAeehvDBjTDCBYrS
5CBRmK/m9f1ILsvayGTSsJom7s47bFebBASR1QNHh3Aj4cZ5EUsAUZVSsysywD/C
fH+ZE2qZC7YnYj0smMvjcXfA2H7sZezTvIVU1XXKqLu5JbfEw91WLB+iYkdwijvu
3GRHm+lELWNQiEztNeviUK8A9KOWcf5TljmSp+FpY/Vl+5r7ppG75R2b5iXOJtOJ
YTbZB0txkSz1Dzdzp3viGpp5FQMKq/BNWx25pHc20ILkszamrUKII1Yekj4nmaj8
70kkUj1FRsU16rMQzhS4Es1DLAKwU08W/C8HJRkHy9JEcE+39GUnGw96H9vJdv2g
QDSSt+XLJ4dK5Xi5UL6w4lrAv+sfW5JLvHOUZLuWevvjkrQgMopEgdWEnLkP25Qx
ARzisdw06lu4Ovj4DtzYQpyT/6AZIcY/1ioiVfaAGrRIrOGYa8ZOQ/c6oWSz9t5T
NhF/pd2+sx37Xi5/p2oYvE4NRIgoC3B60b3qHCGbJrOFQvaTBsgyPqRa53QHH4vA
qkBfLUXL4AGb00EkKCF3WGBnxTBIRnf8Jie8FImmipXq2LKRlRls6gRJ7g9EvQq2
nUIx0SzU4OPUA4SCQlo6y3FuOkrRMZCcsW/HXnSpgjNcTcxlkH4aKDwQb+H54MAe
h3LKBxGfuIbs3Kv2atCElNWBtOPGluBJMRfGfMiLa7MFf7M6abd1tFHlvNmYAOr0
OarKkBfrjApzdOJC6LRAV25IUsP9iFjw+U0H1ScDDUz/g+mOdymOS8vDbvYt0aAH
14pSlkkKHHH9ETi4ZC9TC425ixg4DYOUXe5rNQsH3kzQ+E1nSFjckQUUspt8A3W/
3Jml5Ni3F03n8krzPdEYc17VNOjh+ynnsmNFQx3PVu7bQKAlFnbxZ4HgDbs4JpAg
kj0fFLlnK4wjTQdQdAhfoTF51pe4JGGpcSSe3xQDS2Td4RQ0j/zwr8wDUHx6d6fk
koi5ZP7AHXfIm2xtt8nXrmA9ilDQfehQr9QrCFkSy9n3cLFDALPUoCjTvqp0TGf9
dCM2VOmBUqhnUdE1VzHpboRDW0xTIp0l0WIMcQ68LgFfSSXU8D8MMzusxLFDd4gC
Ox4fiOrnjjDpipwiWdQuhOeSYgMohHGqcSd6BVWJhdoJihAWfxd7cu9e/W17hMRi
2jlKqIqh5OaQ21vqk89cpFFp9S20ytk32FiPAuq/GL7UeDmFeacaI07nTC/i5J1N
oDwBL/g25E80/ph/nzIn099tHd8qbOowk/Mx4+RcUiI5jkvxzAKMkfvS2jPOgt7t
qI4CZJ7daEplfJQ8WEy+qSUj4EGuoVPvefxdDlhRT8qOpRt9Ce1z9413MBi0HbqB
tCSN2V2Z9Mh6zPX3w65EH/u/e/EWnfxxI83BPbkZf/SVZQxxqHU6yi+q9fqaVYGU
Db34XvFrrhmEVqVnaRK4KrbSMHyLwL72fYE7hpmcdA8BuLyE0cUazItgA0lJjLa5
Jzam8nW7tzXt5iAl4e9pYHOBqEsY7v8jwprzB101OusXFzn2MrsYTwFyjPAZmlrR
xb2aPpmtAfcwGGavWdBnqI2/cu6+iNukPYTLjrX0VxO/g5HTS3UkOZJujE/zUQYK
0yTriXyhw9TM68OVerCftr5waUJiQMwjHIIPptetmk7dy8H68XiL55DDOSefBDuS
XLx7NgxVdZKqf7fgEWwoVmOULIXfks3sgK5g8FcKzLVAeLW4JBk3lQdsCFUm4F81
76y3aP4zFytwMyfrr4ZuebgQs2cx/OlCSik1RCpUsztoLRALskEOlXKO92J9zzdG
hY+bnZZRXZfOogSiopZniasazoKNE4+YZbizx/2g/qf5uFm5to/UY8gic0PAREjh
7jgFCr41hv4ozNxwh7mc/Pnj5OECDF0cwo8wV3YNkNd6HhlPv30hNbLihcy2VkWB
Hz8yNl8Nl9EZ8cHwI1zjyqhB2xicHJvZNkeQmlYiDp1k/nUX6vu+9mL5DHYh5NH3
n1nZmT/kAC7oeoGOnnMNHH8oxb+bZTMVYmWeGtmk/tDL+nqZ+L/ifJw6FhinURcG
zgTrH7v1wSMChpdl52yyyvEnvNuDtOHA1lh/y/rQfXVLCv/m/nZgJ1cF0NPwoTzf
WIdo1zkoSLglvB1vFbghxxbf1wqbMCXc53zumUela+faQuRXwrLgEhfYwY0Dd06O
Pfaxrz/jh/7X/F+IdINckFQGxp7RRc40GmMwIbRfpZdFwWNNOEW6UXodtIzqPXn/
ym+j5cuEHKmmfxx69jP6mBU5iEHhNJi0Guhw79drUQPNz/GRPg9Pb4RElDB0F9fF
FbbHxXT9ODDB+gsbSLfUW1PSWH/SdyoM80v2FkEd6twdWoLoZNbCv5747jzbLkmd
MShbsgkyyP/jo3Zl/07nUnBE9GHqvYqn40LBkHRPiPRDSvcayHkbGtodquX6AP7K
iWYwWzRzUp1obIA5lfLA22UrDKIPTDoexfSJdhzUTAlR62GD1HtpFXGRoziGBOnK
jy6dyxtXa3aSlk1UY6sUOKNh8Qzr+ETP8/2AXRn/zD7T/nZQdnh1Hoxt8UHF+r+K
pXGyh5HEYveh7jy36BMFQXeuT0/QonzaubGO3hXxxCt/yVrHhowXpPUi7fMj3tgP
yZdg+DAOiJHKCdVeojtQXY0EDWwmJYXJWfKQRFWTWoViQ66hs+Lr27mFtIRtQ9Dd
yXthtUFLhxerGN6WxScttgu3ZQLpEq2YQrRWIIAOuEVlAG+J6OpWHiCkP6F1iNoo
wO3oBmh83yBaD9kPfGz+jKflCTFQDISSE3goTBYhJabtMRSHK6c9TGRtXZYLUw55
OWq2e2e8X3p8bWcKeKfm6I1lwofLIThQL+Pf0zYMCp0+f4xJA2/MVWPwItM5IZ8/
t7Aech14BQxsx9JR9f2sH1CRvHQKGMrw/FQ9UvFfAgIjC8haUr52BQFNfIjMrobl
vUnkD4AVjYnsV6wCQfU7Q2gYrAY4NTRTF5YiNXm46X43CmqJ65oxao0Dvq79S2F0
mE6WiqAS0FaLuV+3fum+AzpoQnnaKPwlns/s2ohyUz8LKQhWmXP95iK33lFajOw/
ZMxY22L9nvngKa4vMfjUBz7ObhvpOr7cG03Zmvn9X1qMA6xESa49QsCfgivoVePL
lWValDXsUPvuklDw/nXBx3W/7w61iVBYt5d5RqKsMCZZ/V+koqiHe38FfPEOQzs6
8mgFrimiMXYE3cPRVVTy6gllEU91pHwZwHp1lGMQHs0/guPebqrKI/B6WxWLAnqN
aUvF3qzT/Dz6MRKLkpRXONaG/2X+aTdr+NQVFbWB34rAU5cSqv6SqChk9DaYjJn0
JVUvuslLeGJCsRu2O3/PnMowzn52MZoZysU5sVkj5jjkxKU4SY5fb92OUJB18WKb
20cQGxO8BFIrq1g0fNLEyX7SFtayv7hVFsNx7m+9qP+fRVOKEsQzt+WhH0wgjSeV
ijIcGc+2t59WRdk3mwsJDPAc7o/hlC0w6GCWnQTH7QXU31RpBKdDQJIatVNpYA6w
gsQOlSnpaMFlFyRkPtiw1afJ19KqpLJJVAYONwE6BandTXauAw8/eeIgCtt0NHNn
VCm1xoTV30nZsMXXDZDCfqPop/MaTFT0XRAKbh+DCe6wce+FRUoZJIOSsV2h/6mB
P7fchDx2z243IckHURCBw2q8R8D4Xz8+J/qFHAIVbT8HrsC/NAK70FhU/3CVCUoc
9t6JfpZqNw9Dycu58XOzjOlDvsJGoaNdGfniRi+9sZPzv+J0lTU9+vUrMkYNmXA1
EGWGhjMnUwlbiV/wTI31Lgb+KX3nTEtWK21kNhq6Net018XbocWRTSmahmIVtVJT
yIGTKWVVsUs6fhBcTmSuwnCN1+uvn6YGmPIoDX+2PXL3XbSRk71fHQEYM1m2wScy
6bGj9V7Lnlh0/Q0KU3JohgphpFAGXckkcpod/I2FSJKPrySw45MfWIIVXnNhqls/
o3sKcIEoksEfKvZ9J+g3vLtz/1TA/XUCX81GwtQ8Kma7WEfFzG3Rh6WAYfbc5OrX
41O2PTO6Dl/YjdQMCwHgzD5rSftLq28WroUAKljmq6GubFIUtdQRcPYntQlJ69u9
IRghxnXDN+n63JJQqY+I477UcMHDB71FZswwzy1f8u7BfDXwk/T7dpEe0NKGdgmi
NdN164useJvY8IJ1io7eVmqpdidtMJsb/swtyPBb5Slx3HCFmJmZMUnaN1OiwMHN
1LjlJLab3wLf0GJAy+/WGSb7hP9oWHhDUjZj8Fu2dV8fGtkbkkxjNCsLrLkFSKyU
Mu4Xwb84YSnyYKY83hBquwAW6IvR6Z+mg5lachNwe2PZPbsjQDvJMqx/rXmNsCtu
pEwzvs7BB+KdIfvFsXTAB4oAZeEnsRR22qoHFNfWsi07ayUUTiK9/CFjhBUKpSj8
USdvFSX7dEOH0l5jW+P5x/zUoKnRW/JhIk5yV9bMbbE6Bojr7uTfgB+J0Jw49DEF
PR6hCOvCoMhB30xy+t9byiCZK+CMWPOzGskpG3XzsMToZ9MMZ8UiN43rWm2fXrKo
tK5oBU86QvnXbeiRu+5jCaLJomPdeOwdSuInNpVfCEmiADqaGiM6WkE4j/z7Pbv7
UroFRk6PYblHl8APyKie5bao2eiaTY5HnfN9LV+ZJ003wK6VU3QEwvD+gQIy/1Ru
YeBO7fEaTreIBe5kgm3DILqjXbNw7lCejARyd5CUputTRKQVclOvjPE5w7cCXiEG
SxQChBUdGEia/HaRzIukKeWxHnIADTD6/A2CIOkcdtrC3LmqUEDBUI3PDyGwUkEP
n3d3UHycGVB6rCbVlAd8+ZZFFgA8Qo3MNXJYhMtB+A0bEFJOUY4xae/bKpiqqKNU
ZOFJdqjkw+1IRBDI0Fk2nQJybzlm/8CteBytMGXKMWcT+Pcgz7w3AstPBRUQoaxk
sv1NFNYAstwt2y5kjX/EQS2mveWt+ufYEVv9HU1hr6fTcRN1je2oIbXHT6dKJjVO
vumMKhJlcl5dStu6QKm2oZ6qfrpLZejtRg++UDxbsKNVnNjZ9sa7L8b+7jDo8Tvb
VTDQGpvwaBUK1O9TuYMewoM/82MRbx4Gmpp/gVfCFMJsIm6RI2N6UZbkWF16ktr4
aX8cr+HAhIGt3VNpZgXGT4iAapd1E8LwWOoRwsRtV5ofN2bzB+uiLjRpCfyL5Y70
rofEekAw1ulx9Xv2u9SOaRCoBjBTQ9R4hu7XdmYcSCyPXq8eo2OdbCX6fYewmDGv
guY38f+nPIYu08aL/eQ2UCHg6Q5tTY2CVcY0aO084qdW8Yn0V7JBGWsVqxSpX+X7
2KFTA9Vw9SQMpjZWDVDrYHEs9a6w1r4GtF4IBRAPt3vnxCQzakf4vARxLU/u6CN5
gQUjHAqh0fSYr9bmnawcpEO/x4T/vcpUKQa3YBQB/iwo6wO9MCRofqUddSrB57gG
7PgnytSMVUkmdpByEwXUSed2Qx6LCFWHs6TcL7mbtzOzPGZkAVsy+kgd/YgSg+xA
9WKvMb/C5bmNkaiHbE/5Wnszoa4GPvUEKHffEzNV9hbhWnnUKLC0Mzgx//iWEbkC
PQHpUrGPex1D3Q77qtms4GzQqL7pYx8DiA2dChNYyPhxgsxsUaoIwuY1pX/tfyin
7PybVxeKZnco0qC9LKxt74P8XsjdTAX1nMVCosWQd+SUVL7/kAtjw0RfqWVckTVk
t1Tigjace8CD3B86xzQqWlz4KqWeg1oxU+Ev/qEVdGJW7iSM5Wm7YKE+llkHj+Oo
RFUhOxaWRAPaxYxBttIj6Y/w6CgR/FeeqwGf/DFk9GVOcZuJNDLSgJ5YQ+haHNR3
koZGl1rC5d3hor2lMb29J3DseO1wX04kyt5gwag2EPpMJyZOTV1xBuhqjKEhIRjz
1XCvDw4Vwf4tKu4wNAB+KVlNGTSftH3EAoyOXzhqVJKMjv8cadB1wTW1uMHDDe5G
KoJE3ifZgiR1zrsExFVf2Ovhn7bdajIMHE3yRo9bhwMKa1Gcgm2S6Udhxjur1NJo
qTTRM7Y0b8kp4u5HMFyO4pITjVUYIP7crUswA5jMCNE5Xh5LYDfgq7PyNDYaT5b8
23zNSyMEnn2pnjPKs1w51yP0qXXNxnicdVxvd0y0zY39sOOnt5kPpBJm7G4CuorX
2xun9yoJfU/FDgY430nPQPDGu+yZLnaerR4XtWKGI71fNGJp7kkGSU8Vv3Iczn/q
UPZlBEEwYHF4Sc5FjBizGlj4TPu9uowRK2ekLXFEZCxwmBNw9f26u9OwSKeVlXfZ
PkLhKaNjF1EfpqFbxekoqY01oIXCIIKeZ5SPdbr6tWLHImrtWy4gChzV2nxCIyEm
RHBH+qn+ta4aGJt3l9uWdnMBF/lYDl9AWJbD835i0t68xnLbWTL4xVIB1VL86GY6
/8i3QSXDyWJXOpZZzkpGhHI5Tws0wz6LjKsIJjoLBRYzTzQLa6EmEnAxZQgaKrDz
fLJn2JZbB1whZErEsg2MsJuYXWNm6spNAtYdJShIihm4jMssUaojMGa1mUazPVF9
qhR5Sab4PWyf0inSZ05L+cOJ6J/ld1mUV/qKKApnVtvpR8fByBtrvmNf+fP8vUSg
X9KyBakcxFP2kFhj/wezDoy8k7pAYoav7yfz0WcMFHzQxa3ao0y/A5+mFewpu8N7
+CzqxYglez1Wp8AybZGXTXuygvPJTouDX3r59i0PgkrP1LYET1XZb7IslzDPAPEW
WoYejeBDXs9eQ/Y6HQkifAT4FhoLXF+ouHznY1g3Fiz05HCk7xm1HWJWNG1ar9CA
pW0eWlznuc84vwkykkc2kvUnMgEFQLgJZwnq2ChvtlYK4P/ocvJEqVBtiPxd0Epu
t2L6Ss1P0EBBM3Tz4+fnvrjRpDiHTcWDX+xiM54kyixBeTrRszKrCrqQVlyjgYy5
x5uvvtVjkjuB+XGgt7nzudgDtd8uc0kelpAzvV3LMHwwp8mtT5YHM5rQnJJHm2dw
sORUzXmw35Bo4/S0ui9DRIfSuP5jguYhBB6JEamUExNvoJDP1EqPg0XDcGwavt6t
BZrZRTQCbGVy8myFfe/tiVmwgoci5vtimDWTmAPiu18DoCjqP+3UzBJ/VGJnE7KE
LAcyqjubwXd4zkj6umTZtk7DEYrPfMXrK65iy03M4/UoaXFam9y4ERYs9jpr4gSb
20x7vMIGX8wg69Kw2f8abrMm8AiR/GCWaNsyzp+qpwG80QxsQIa2/MUgrZctil3F
p+Y6t3k0qLO+7bVghSynop1+KHgDSYli1ByyibQPv4QgKyQ3kBpHThG2FW1mp+HN
ieebHZ1qCqoZjQT8O2I8+Y7s0Jd0ciEx5c5NKeMnGZJLjdqMj1Qe+5sLShnUP3FT
fLKnv1ZZAm5WMC86xUFhoTuLGjmrb0lXuSAiNEMaQyyHJ0ItUvSrFVLgObAwEI8z
1+FLKrzQ5ouA14Ju37SVVV45uOHfeBLAvX+/Lji4Ao9V5qHlsN6NIzMjNfxePTMW
yW47tWUqms/xp4fooLTM+4mgaIeMvlGObgFVgH77/56/tKjdM20bA3ShFCyHUBOI
OEh4LZlz4460tlYZRVMjcDKRvkK+Y/ct+I0A5X9dUE4vb12cGF/cywtZgCWWi3qE
yeDGFvmbQUtDF769xMpOxm21UC3AJ9yl6kzue8MNlKRaUWvS+SDPgqAnkpvZ31qD
s/goXrrgrQe3pZ+zaaVGvQJ4dWHg6DrtWMm0V+J4Nj0ja8YY/QNsRml4QAXRvkdh
eG/VzSrw4/NxgcKtJNZVZ50zYLYf2dhCvDKxgSzRbroQ7b3y6D98tyQ/JA89wTmh
cdCDl7Ll4llrbAaXyn985+YhAt+EzHu+pJ0xyeYGwmcaT9xwNnvEVxYFNufwkwYl
raa5pSSjL12K5ZbVPkwixRYbQ0Sz35mKvh5zqXuGX8//TQjhNv7tmY8LT0dCXWS3
dBh/WPXOysDAFEymlulvAH7L3EN6KL88lG3BtUSqnjfIBlJ3d//t4n6syXynkbgj
Fzo14jE2yMxlYB39krGOMVrnyuk1grFFTHLgoUC+yAjCViu51nqOPqIIbQI3w9ru
SbFYzUV8tsozmWBPcqY7n0IDjrgvlEY1qdjRTQc2osHFDFIOq6eWJOiAwK/Sb4KU
GUR8Lo/JqL+wbFqktxuhAah0HnQ4p6NlwJ+W12in7ObjFwZxFwurIhrYblOPJq3/
JJANoU5MviPHn9ClAWh0BRupEXYl/KykiKdN6l+jkJeeUl38ldvwo9/WCVHXyOO+
yLL7LyjqvGDlYja1Yl42cd/WvM4JB2Xo36XFTGPBOChChLzivAubiz1my0RV1q9Q
sEe5Y+/zk/qNfQXLPh239xaCC6oU48Wh+Bm0+HRf66yH2sCkZvWTB0mX6urXSS3S
I0OkYxmtcPxV0VHooJeLHKMs1B4dTQUkW/ASA+sDJuxyYhlGYVBL8qAC8Gxdf6tV
xvhd4RAQecHx6r57+4uY5gk/w1hHHu/alB+8hE6LsZu+bdun3Nk3Q02icS+V7oid
NaydSu+Fwxlr5HJpXPgphV/FKndyaS/Ki6WW8zoT/SCVdBt3dfC4EbWrsGRHIiw4
+mxGaNg0e2JXHwNGeYtGSmI/T/QN8J6OzlbqHUG4nXtAmLuWvrj88kWaccwMcu0h
xZ5y/yaCHmu6F65Rppdl7fHSDyh9g+m9Iz/yRd8E3CLKUaYWCqXLa7mWcY/7bSds
C3XKpQqrJUJnvOwSN+deVXqJuzDeiBRXeLwXk4EPk+4h3pnjfMmeK7/hF2Ob1WeW
KNFL4k+0Z+LaTAPhX93ajd+7wGSim0eEkGKYyEju7F+bKYA6+GO1k1KlGoGKB8QE
MvvpK3c4Y1pcsomgIGTda4ULOyeqGy+7D4GdAls67CBdv20jrHoi77YCsF12c5CK
F/IvZrXbxvoC6Pja1wrxidBKCY4Rig77209LkzXFPBRZbvUdLY+jPLB7ro4bYRXo
tunxpdPkPjCNUMpEaEOOSvgn5dhJ6hT3mxm5RtSiG4MR+4F3qKoV3++XEoADCpfw
B+0FuPMTnJg5vsve7sN2bAYHELBxcffxT40YPnKrv/ehdHVwTMQeDEUIpaWUtv53
iaE+/A0bNXCEnrZCRtfZKWTL+GWhlpi2IMKtcrGOcVczc4NAgBysC+Mw20TP1c0+
/UpHgdstO5cQ/JjhICE1NnzBmYhHDDTXP2SMHkIpaGqluK/4dNVDactvw3X8L9m3
Nm6QccReX6Y2Ur/C5Ih/lzXWYPOYfTQbjche/vib3RGQsmst0/FLNRAAdntewRc0
g5ruNNBpJnUwoNqemRObwmqrfRUTWUX18IVuiIU+5KMObq1/O9Rhx/xAyrJV5ACy
reGl+tWAn/qqGq241QedOqCm8c7udhIQOcLvHuQsncA4wPoxbS0y2+iv+Dbj5MA1
WWETUz8Pm4MusneioTFjtE2eJ6Bz6OuhPyhEhHk2uVE4pkA5xa7gvGfY0IfglnES
0DWDXTDBB1GpuV7YBcmGwa8a9+QtmjnGryQA7BeEqU+MnJPYIYGoBDrYA0/B+cUb
g7O3ALtRiUjbL9FyzJnVqGzUCY3Q94jAM7F9QAk4FfrrmzgSRtgjNUypOfcKIA5s
HuZq6Z0GxbnJBFXWlrnT6B4/hI6gcJrlBkLGRIv+plr423vrnO02C/catu20TcL5
16GccMop60Nkp2KovEPYmUhLSHg5J3syovhXDxA4fSJIhU+Xjat9On6RMIYYIuXK
qENN09Vvjfx8+mQiYyZ10GNHZEBQ7DEcs+qfOrvgWuR+dkJp+9shOMXUydoV73yE
AMaEfXju9K35WZ6RN10dG2/yX6FtrMlb2oSbu+VWmfZBnwiUbSYaefY2dbJaCYab
tTSl47XM6y4xcr0+9vEQFIZRSJMkagoQ8q2Lo7NQ3+ZS9gJDmthdBXDcrBw7g28U
nbqWBBEjCgB0fTQfOOfu1T2QnO/caoBYc6zISngrD93gPk8dUNxotHHh+4HeVbIM
MDeIYxcGiMWUBImbKWlJjBKWQSnEh6LIu9LlbGECN8GhOpRB8MYEa8Wsq4q3kUb5
UxNuM5L3LIcSddwkE2cgBFIJ4d6iW2lQ759xYTv7OSrc9lu0fqqNYkGgKSX+dZyl
9JD7G7dbnsEbppivwdmpb41yJB7SxWWGyck1sXWy5r4j9B4A56o/bRcluTjSorRd
njY31Mju8f4jl+2Yh8Pg2YGT5shc7OtS4lGUTUnm3eMw4//N08+2PlADVOKGwlui
EbBqITXbX1T/Zq6VQUfjNIXBRCzY3u0FYCiFh/o/94O8iRhvQ4s62vxtuftmf9dy
EtY8aMYlam52aNL1a9bw5FGCUzw+N4WMveW0DQovajvz3EOqFlKrxI5fUm4UUasL
2Xw0Lorj1PfMH2st1qaqwCKZiT7SE0Eu7lREtm/vxaLKLlK3c85Ziuf6vvniFeX5
m+8n1QqTEDQXpnx4URaySDz7OxQ/Nu55NQGZ2wbBJz9kEwEoCxzq+fNxGUg0P+ZO
KGVu+7iGRP0bzt+BZKk2s++K/xW1sAiEsJuvZTVmwDpuMOg7M7qk/ZV/Ko6pWHyO
jVtlHawKf2QrhPgspoqTk1TrLxHprya9dpluMdK2oIMeZ3K2CU3Tse3MJzH3xFJK
9sZUE4c7gxl9BcQOxbPaaLzr4V3cArym5LT74YMTzHFE6Yuc/OBBsceFxm0QsBZs
OD0CAXC4G/LVvVp7zhu+fykkI94nNi/OGhM/fM7XgvEJ5z9FwUzmH/JzqTXH+wDl
ltaLP8jAvIm9XQCEsHPAlCsKkFufJDE3chzhkxi/T3VJJt5TdrmhjYQmg1H3gXBu
puHrQvItbVFOLE/plME1kCzsn3NztR9FXeqjHE54lsHZ88NZGGInkD3ZVWQAvW/0
E7zGl1cqZ9SytmYtoxIJvRrF2Ogv8BXMF7NSL+MpHRfmtsdUEPDqyRFDlMBRiozI
6DE7yGdq8DBSkFpFfwZwKfBR/mx6N1AL9OnGe23xTw+2Lq9OAOTDDQL/tSNgd+pK
plgFkimSuvo6irHQQ97xmiOEe41/WBee2/SIn6JLciA/FYtJzcygxputeu4ZOvXk
/5uWH91DzwKGIYa1+3/c+rMVmHlA3+w7KYn6oImlcxexf9YIV1epyPEjR2G/ztLP
NJD8F8oLKw+YiqR73Bt+4xY1CNOBfReCQnSaW+2EFx6lBqTmZ6PGBqI34uIUB0p6
037LF5GrAMgq/c5DK48uqTw7qyKOy4rc95nBa0M3v8tINnDdeHPPkDddh2eQw6Ms
BE6uv5yIVBqGDU2JlHSfPcSyBHXuEmMgjumf60JieahTtsrWIVhB11SSqzoULPCT
9H8Q+k1w8v885nN4tBjlKVXkWRnZUdH3TK8VZ9tTjAP0f6eYsTYj/j8xgPOoLe9G
PQ18SsKa7A5uW0V0F4T8/B7NEFNLYhhpACVbKIiGEzKvqJXW819UPYaLG0pzhRkG
4ZPeeWZIZYFrHM6lbKu+dymKUjPBkdYVVDbs9pr4fKJq46evSUro9rEO+G4s0e2W
/cYMM+kjFvvcygnVGj7PQj59OAOz3T3GoAsHu3thpMqPZ8Sn/QgIgTx9Hw2hoEre
AYqGC7YyhHFolMN+Qjx6x+uwnFVNiaH7UufB5QteKJHtBqQyvFWOyHK1GbUk3Huq
t4mE0Mtz+ziGeEog6lUIv+gSzuM0+CbIr390TL/gsJSLYfOaiotyKSqvivwRGB40
b5GOVnEK7fKmvlwxs0lbUHXKtcF49pzyjqV3SQp4zINpB5xqO3ZII3p+VlklTS6w
ssyJ63XCMyppMNbnhc8uLcCspjlMGZLvALV6G6F/DA8JzCLmOF5xu6KBJkwBo36M
uKg4hqJGaOWF+EGc2l8Uj1Gee9+gNSFFID3dpOiEBvKmyCde5MkaXNQ5EXsOKUA2
NxZbPpPrgHZQS/doIRIsUpCuaY4B61kO5olI3IEiv/VrKKgreA8WDCD386cxQI2b
504lIPQbiE/mKyZGpT+1oOxDHAXlQrIZufgLxpa1iTBEMwlFJTJz0HHS0W0OSZYu
lYPLJQ5SIJ5ksSKM+5z/G35YGRnhTCAwdcU3yQtxJl9R+URWK8FzC/yhdRhujTIu
7NEce8J0G/cRJ+gX4u4DUYhfzzb83NLWLdRGgcmi8pd07lJ0FH7zXMt/lu2PuzYp
1fNcSP6JLB5JrR6NJkMXkLXG1LnPa5iA9EMeIhH+yDf3BSAJsP+C+0/zfg37iYHv
1M9luGZ6oSy7lJjSmvhaIvuxlYnQPtUqC+Vzx12lQfijp8Y4XIFTiOyskGKhmW/H
lGrL2aRTF2wuTpGK6BPHtX3QeiC5FZZgvI1LLA61PpWpCpnnqPxA9INLqlhsIZFF
pVMNxmf3H/v2kdZHb/4n+TfvGiio+vEdl7pAddGv1UhWigBWDfM988ZB8EAfQrHk
Pt0OaNhoO8Hiia4lhHWVOb6aA3aYYs9YhcGyOoFAzZkobnVVH5CIxeeDUXVBEXvO
k+bueLXmHWe9JBPDyTLY9b7wqTlvTfNgMKg19Bc4dcdDLbsAe04Z6ugZcmyosKw8
4uzc91SVlK68X/cQAPVjU30lN7Bg8rT5u/Y946msnYhQfBIK2XCWuWF1KY4uIuM9
pxJ7z1BPUenHpjIbc8PjsDgd7SYbj8ECW9NViyZUD61/uLyC3PWoJp/m8L9Oxy/n
28a4Jr+FQGEbnv/Haie/hS2KYk61EUbcEwW4i2NLmWM8m7wSMvT5hl5Qb7dOwqZB
3dubSRkz6QhJxdrwG0WFS8WoP+nulxhEi9HxXS3E9Z8b2CN9VFj6AGaDLOiaPpaQ
qRZpOORILwPyNz6IMgliNSSt3jQBNwanqRUH9f9+9yxznCDyLrX8Se8arHPBqPV6
b/iPYE+TXFTFda4n7fsyr+zKgkqB64ytpXpoua3rI8+uFnERqBMCOYnlrdEzseQB
CFbLKPwWmGTonwWkbPsdGiPl9CiULFXRZjjkVBFVjLYSDv2pbf639twpliKepYxV
+Qv6HHSN9LtZSP1HgT1o0ah0ihr2urfJDZLo/BJqqX0Z+IQGBQMIGsk7NjEDT7/j
N5qgoRJxMxm5oGBkVdUVWsIn0sOYnwSdS4+CpA7DbTIWpimyURVb5v1fOLOM85ev
fE21+5wSiYOWmaSwDH0RXcrkY/E9Az26tCW1HfjVi8lbettftICH6fy6vOAQUqYR
hqXrbxTCu9w1mamC971qF1ft7HhaPY/2mTNSrNmqFy3ToZ+5FFEkfT5ojq9hbBOE
PgnCEAchcIADmjDWG8jgwnwQPMsMYN0q0bWsKFNkqkw2fYZL5wbfNuH+BsN6JK9d
emY8XvdPf4QQQrC8ZxLf4pYLSnQ5PA1i5Wim4ChItGWRdckWB8A8OxFDuraiiGr1
q5zGAlmU0/SDi1Y2+vQMDV0BXRQaeHGFMRAz7FyyZYA25l+BsQKTBqXAWj8YyOVF
QmJGgGN2TQTxnWQBhUGB1TVXxtmuIqBHOnuDXJrcrKiqHTECBCjICKFxTytChwlf
3Ba0x31R87TdfvncMg8+TetP9VVFdc86nCd3DM6fJ6pHSi498MXDcasTwvHymmX1
5s35Nmb8w600MqfxhTog2QAbeQytz0XplG90pfpZDGsT0tUq1gYu87jaMYyvREmM
gqFe0qPmvDV2XNrA5yWcQAc520b60EDHyfN7ygStiQUl7fySdjSh/0PrYxJlCmV4
zwaYcDroGBq77jqERKINyLymvLRLS8B0UfGtmlDuZPK0+ODvmkwi5ERWqVZbYY+b
VfG01ybPWbob3GWrhtG3nmgmuD8YMp5lDz6lV673TYwtyQFsUYsf7mG3FvUD9mv3
vPeIcZsFwWcW8XDu0q3kcuS7VJ3R5WPocCgCWjuJBmnOt5Rqh/+TS6WJgomV7wA4
GNYBl3A47APuLrVLLdIMHFhnweIzakMWTHvmTIzldMwk3P+syHUxi9bKG0X/uFPg
OqlSLfZ/qWDK+TNObXjoZP2XAve2MQ8VHw9qalLiSOk7vHjjKtOWaytDhBvkBV4u
ZgTzRvk0C9cx0O5cEWbbCXob/QTBINEC24afizU6dgZJnYlCVPMXJbjm7Cc2n+Dw
W6rI2TiPdWksmtLUenjpCQa59VQNMLm+j/m6YBhwBf5spzXctJXiyQGQMJv04mAM
7qmpKfvYIPRb4xugchvq5nk6zfJMQbMOT6UtUcJkWw1h0e8OXuTRofz9Gu+7cjyo
yC3zVnhgo07ZOn4NTdZMHjHvAyowGFsMgbfbRCOPD3VHZtC96pX2BjaVXSw2aBhy
8+ZrwnqUuMHlFnb59go0fFDuF6OXdVRUtJ+UgfuZ0VQ2IBYEefWoNPy9WFDKl6hS
ER5rf7IEOZ3RIWFfEA7jRNmrDP07yapWdDmm799Bq9VWSmjrIj/WfQ1rKMT3Aptn
ubM+jDh2kkyhh3GfmX70x11LOaU552zrlYluubYwnwzFzxmc/YJlESnJtNx2hPXc
Zhqb+TnU0EhftzY1Hi0MhyIEmeb4lzBshYuE1Q6HSHg/UT1kX1+ylQhZ7sGpNGC0
uyNTyWOTVhqjg9XlGe12NvUZ/Yb/czSvu6eN5kUx02ULqBrxXIRaaurdYsosOOZw
pzhY12okd48pmvdWIu8I0Fa9iCkfoxE+/C4C+O6AIKFROoaHaz0KCjU3JHhGFRe7
u8i0BPoazJBC1EVNB3SFIBFeomwqC7Khl7rnOMJqowMeOKzNO3wyVAiTJ3Nb16un
PJvwmzH3nDU5CfV5JODC9ftpA77MraQ7JoAQsa0JW011JISFU7LtEywMp2gEjXkF
Rp8FRZE8yJzb2LOi65v64o7p5/2tGqBGhlIusnyk5JlJsVlXzWTLN37KDMI5amOD
bKfxuEfkclOfBSH8/ptAg3W1MCLHplcizIeHfLjPyZrhE9xaJrkYcaFVYHjzNA3Y
HJQczvHCZojho6SEUanFkcBmh/O4EGn+s8bnbUmaD0mi/lN56s29SkkMinuw6M4f
ZIifCHqCQK0kcLUG/ATguh1ahQXEAEtwZpk+Ps99xlg02FY+KHrEtMRI5M55FrRt
MIceymxmCg8ffqM0tkzVu4VIp9UqoAm8CZ14ey0SWPIz57lPtwn3VhKnJuft4GP4
cRS660JoN11b9bFcvmkV3neehkL++AvAttSHkF3pWZrm7Bd2Ajansk6HmGjzYdwZ
EmjfbxWHguCtOKSsVRl0s8336fobwOw/0/Enr+ZX2hc83ry4b1DtiUBR2jaWK8lI
dXD3cmpNOwnGoEb1uijrvsumA33s/Ip2d0jUWHFxZNjSO3vpmjTrc1QGNwjvAl1j
AQY1uFaEcDbhqd6cz8qmIuuEjYug9EZ3e1K9yt2/BUfVK3BztKh8NWTgmLnIFY25
qoa0wosvlBMoK5SdST1sj2UXFVqJinhp9paQNw8AVPSwqwh+IZ5RstLCSyA3yXWN
nGhTxBtv5V0sqrztdD+6lq+tuitEXPnY2mtqN/Qnlme2rwV2iaPb3bUHpW28hpyD
7vorwULG7uRbOQGx2azbXMZsynnNash5WswIVNnXxtIaicQvFcYJkiZFdDZ9BCwB
zrq7a5iEEoUl5jcGGPk61ejAMC59boiZWClXXyxWJL7fTlCM7bDfXyTjM4n5SNCj
CrnfIa8ug5uYYF0zcpBiOOxcTVzhflTYuRnFS3Xa20YzNdVhR17VZ5tIEdeHBrU+
6Gz8D1smPISnNq/3CEnsQats4Ucsz2b6mrSvV+QRTHJmW+6rDSW3GZu93rioO3F9
Qs0wKQQe6BNdoIqtzJQC/64oppIldZ/RTZyZb8urYrZW2iie+NJmvEYRz0gSnthc
HFV/ia1UknPNZExRZFvq3y3i+hwuRvheIqyBndnB4KnvIR5gd9TvIFX5OaRwcxUM
cZfu3ZlSiv2uADAjygYo+sXK6LBGwxMDkOfCKYy1hjKdhGygW3BGPLKx3Ag6gt9p
mTnSaC2/PrdCnOiI7o7Nbfl6FJiSB09EQ10NijJ1PyQnymJGz1cMxoiVxXoEZ1a1
28FEXBfcLguKmw4HVJUGq415KmFCgWWpR21XQ7+XXOn8tmc/exKOq8mZQJnW/YVJ
A6C5N/ok10Zjl5oI74yQ0eEcSIPJJTI0HpcEtmy1CiEHACHdP10G122WRZrCybPM
to8lgvw4uprbCSnlsZ3+CEJOJG/rC0mf3RXYc3RqWMEzUiNEls2YSz43aLiGTg1Y
KccYrW3pn7Z+FdTi929JZ9Tr2OvJq4d5BUtoEQThAO4SI7iH3xvbaY4pxPglARdl
eBPgxzFudV9rtLcbmeIdRNsVf+4zkMW4TvjUS/XMOFqOtdYcnRRDCI5zv/kDJiUf
Uoh93It9U3aIk8Rl8d4W5xxuzR6HCJP/CoFn1JGKw4wkcOidqBlGqmKKppILBH5v
7UZUava9Ffv41ACWhQrC4cyhe1zI5VxAnfZgaljXqExFK/dISLHzaT6mjBMgofsZ
GdvRy4peHu+rmy2RubnJBTyJFbLsJgVJZZ6JMcrrMSZ41++rrafcgQkm6sL/rWjt
KP4I4LDkwA8+C54DaUQrcBFlpi6Ur9+YoYyxnkNL1cLamVwnPtyQj5O3E4AGtXR2
PqmB55cqAx1HULLx2shEbZ/2e8s95FVQ37YFdbIVyq1FdZ5NT6euvac+6S4Blzls
hhj8tijvThxJF0mYdRHPAu9+MQORq1RmZZHFEeRWWiZ3YIQYQTqKRzHHlboO34WN
YGxehLhO9YURosHERiMbzuG0jUGV3wO8a1/sn2y1fPXDq7qQce1QLboB07XAPCdK
DiSwinhLKP2kgE5V0aSSpV4/c5498oOvAXDYrK8YlaxY5VWHkIxuaiybfD21E8LI
giwWfK+adE1vt0zuv2sRhs42El/BzFkMCuAClQVxBiM7POpcESkaFCjnjDL4nedN
8xO4q1It6E3yknCPqZjFvhs5LlVvDGcb5bCAzy4LzS2p78pD06NQlPgGtjEhoZLN
6PHmO8dqDGIljFCiWavjkqRet67tJcy7reF8Vnm2VDcoMHKiXgWoS6ruOa3iz1vJ
g1azpKdm5mbk36kor1d8tP25y1L/1icTXOtYf1AIBUBWmuKJWUAY1U68lhZyWpWs
6ff6q+3AtJNaDFKAAbB2ZYD3NCi8drSbfKz3137iAPScflMTGws6FHq4NoOVYirQ
7bruitwmOsRW7SRx4piXt/lKM5hb9fUYQ2JDmJCTpIw+oD2Gm2CXDdRIKduuwdnk
mokGEvzTzEO6D5B3eG82B851HgvmzW8JdfaGk5o5y82awLhs8K/mlINqWBSbRU9x
NUGqIxhzRbjQHeYKfLgfk1+L4opIkYG/iVVABx4rV8cnKD4FiLa914RrTq+Uz3oN
rWBVpqUkteheNhN0TuSlImo6LQRpXcHg9kz802ToodpPKjvARTCEbCwOtzOD8u1+
1MAvH7hTLn1fo/bzcj9lAjnscAR/FTFtsg8m8kd+2PgLSYFa/NDJf8DwF8p2xT1i
4NtjWE6ZJJoCJhqdVHlMAA3Lh/VYO4cWtDWW7+I7mH4iLqCL7j5SK/L+EbsBUS/b
8odX+qU9TdvuFQvi7d4UBC4dBO82T1uit9PFaRW2jYsC1fV4n/w+PiDtH4hGDidu
J676mlADT/+p2niRAwVD61tGYYafeLtQvMxal2J7X3vQNHi1hK/lp/nXwtgJ89Tr
u/z5FC2cGRlG5s//94NlIwg8avphhSdGEc/o/IK0ZC/miGcUF8vnb4BIE8B0gcYX
CCeqcuevcBQ0uuZBJMPqamet27NgpvI6XBTAG899op0OuS9DTU3JTut573t+QdsP
n170Hw6tJS85NFVNKdrZXd0Qbz/0Pb332Bm7K9jpNWRLf9NSFxUuyzH+7JPKu4K7
1X/WBV0CuB1ZEF9Mmute4a8GBKgfPCQPhCUfIEPwoZ2987UvlcQptktC7rvEmmvW
O/8nyDN5DwCh7zt/VQRIC/W+6csMAVXIZ34TfX1Vgn1TyMBNgdMFvDle+2mzkdd6
sDUeP0XynpPOOqA1iWO6qtJrUelNyPkNtYB9YV+8ztSPWxNb2JfxFg3Us54t20Ei
UOdTsGwB98+y4LLB7LEPWWmnFLyF/rnctrhLklPgzFo0s78gCOyE+L2P/sjYZHqs
3vq/NZRLwuC+0rcS2/ke19OdqSGPeg3mRxAaPdAtIIasHWag9jx4BEmBQDutelPl
LES5QkxZSrXUxBtdq1pjIfWf93CRXkYhIBFdSXi6HtGEHF+m9AHoXjkOzyt+gWhi
8V14z0kCJL1eMR9M5SD7isEAqjaShSMVPwAN6hp4io6XPQhzZaIqHaYh7LY1udIU
A/0Tun8HzGybeaE9AkZb5LHchFhFFJ6/IVo8Z/mgi8Jfk44E5j5j/1U/c7mB+Bt9
/zmEMPatwNUaFj2F03ndI4EulK5ui2Xhm1dS/qxEiXRdUWXNTxV6JZfjiW790dkF
IOyB1dZ4ANbRFxkwLJ9VnwJ3JqVkqP7z4Jv49yF0kBicSBVea/uuDF7Z08F9gZrL
Wmm9PjHJz9ySozkAhAZkaCwKKzeh/N0H6PPga4GfSym59TYbTT2O03tMk/ryPdQs
w0yJetML1IEN7Nl2w5Sh6/64wBIDzIeJieTOTHv93bGgirB8ATWEYIUiZkPiDKBk
yvij5F/eautqyDoIFX441e9zDw5UhWDjRiKOEWHVbV0/bVO49a1snqqnEXYumtmh
pJVhfaYnQWitdH2JuwTK2yeP2wInNRQoSlyvGzhIXa7/cW3yBSuliYBLkWodiBEP
evEunWZC0h8kawCwYE6mkDirfcQkglkVzj8LG1RUgFHdIlOnw46UwPG62Oc2o6UJ
HRQTg/xlxwL6wpi7G+weBLELyNSgRu/invnLctVcSVTqrGKgM6uBMVKlH9pXeufT
U7G27PhZZTAdnfi8AcwWBS384LozhahcIT5xcdPsACg40qMzJmDCvPD8IG9K+vKi
D2t1HE6TOApv9laJ2pxlNB+GSJ0AECloaGlxoJZpK9q5/pmZv4bjftOXOhgNfTD4
9iM+d90BknshgwrBHm+a2Xju8qH7wZA3rkHn/WjqLsdWEeiaU6i0rviaCleF5qXb
2ht+IGgi0u/Ojqe1gpiYF0OIUY5Iuy9XZD4BJCVDYazUJPTqqHEapbxrm20KcJSk
1sheNjd3e+KJSppzn2njuBAfQOUunbGYxaRES+pbbBIg1E4TQpicLQJNvCPqIB5N
pSztQpAy/O2WeF6UWSJP8TpJo8fNAUaHHZs6HSwOhakq0m0ocTlhJgPWOGhd8ZXE
uavIIduYVT9n+dCVIaTD5vD0mbrjfOQn5mS8WAldLpxUwd03ZqrU2rQy517gEaBb
Z5R5cqQSeAc/61Hohr1rdJwf78tKk/2nVW4yjFXMvCAnEvcjKcLN1xqLBcPTECvE
4dyUuRTJr26Ummhpx7SzHC3HZVRyJ+hmnWvkgxMk+c5jNAcLOu4F12jcYvBTw7AK
4P1zR9Dweoj95WnspsmTMDyPajc3SrEYVhPMJR+40wg02VpUQnHxHVohtGdDYxbh
eUUMaEJQXhyM469FI8AIZBCkPtxFEBOuAB5L2I0BrvJlElsLzZ1IjgV0GR3cGVO+
bZjaMOSdc3iB6NSa3OUCLgibvnKRAyz9iRYJ2P60+u0MUtNIKHussfLE0bqjYWWy
OcezIWbWh0v/W9PJ5nrjrSp92ydcYbli2eHXQEri6Ik6hAWzdWo84xgQobRlaw2v
+HEv8oUN/orDCmw7T9QiS3KgpZyxf+O6A4YDyjk3JcMHsZNOFrON0JR4XxnoL2rl
JioEibCRgXk8shBXbNUDsATQVhI0M5KY8a80j5ZFozo7AB4YzBedgAg7NOEWBlQz
vAO+mvwhKgggQpWaqBtKi0iPriY0rf4WdygDpB/ycp2Ivgiqs2b/GmWsUfPn5AgR
gDB8Z8gO3+DkMiKfcwykgd5k6QF4jnhVdYvjWixG2wge9ovVpw5j/vH9z0sQZP+/
zUdU+bRcgoGGreSz6fRW6l3TeDns0b0eHAAxlbz9ZTHl+JqFP0Ii1O2wDebO/TcX
+SSyDQa951Oq7zp0sGI/MXWZQp1i90rbosEsl/WH5PMxE/W/HR4+2LmKJ6yWCFjz
Q+f4aABw8+VHFHT/KEAIq94IEVeMlM88qUBxJLgfM029o/QDyljky5o3iIr/8vK4
NnBJAsm4zvjKDvuvcJ0zwLPpvVdZnIOLu05+7xISkB8xxzjEF7Fc/lrpzrZ74KAY
A2r0E08OsGLkJ12aYpBnDSQgnDv7stTD5l0Pe93QqOKIh/LyZjj/fTKxknZ8TRdR
o6c70IpMzKra+WxBKEvKbn+bR0vBzftPM5Q2yajC3m/u+IuX5QNGrNQQiPz6/wRW
v7qlH6TWSGA0rCgzMnnsDy8RuFxkHAjBhbiGfJrDwWM+9XQ033upbRHig7GaYgs9
fc+bJQUS6M5hpljYZjGEKF60EmiAJP9LbOoisrc1Gj1aKCAsDio/dnhJAUgehExw
tQrMeT/jzLZzhvddZIFrSzVuUKmi98DKA/YPuJNW+SRug3A568J7NLF3AxVjDJSm
M1W40R+5KOQDvPUEJn0UPci6z7q07Q0QXCu7m1s/uTwff8iCeBRwiIOhWy7vhc8l
U+dZpUhnFUtaymzYPY1K+U+1WGK0ovrkdMLfAOSGOxwsPCT86LcwdKhnMkn8OyBt
54moIhJfmiyHjedRqT4dgdQUwO3aL6BKcD2ljb+0YK8DAOaBRFs1oJrL2ZN4AkBe
mW5D7QHBKBsYvX7Hm6WYxfDpCl/iFI2fdizwpCAG93x59QE0/LkeVuH/YrI+b5L9
tyt4rdXimbuS4w0E2f33xtNY8s1O0nGapfqa4qTHMv4cWFZQytW6GZspEf7SsTve
GTGu0WaOGgIbTCv8PlBwU855GDfPtBictq4WnBxMWrbTkDhSq4/JDZlpDpVN0SYX
ifYod9/nx98atPGaNItMpR54LvClEObDxQEKQrbbCrrHk2Xl24a3xVYJpuZoI67v
JJ4FinjTyG1jTdf1p9afZWF0t1ljnWIzlUTPr4MSIKSXRIO7X/7r9gI7NEYtNN3s
xfWCZjbH1KKKeJaUQ8UaK2GUy9BmdB81N0JeXG96cDpyEBF4iTFvLCP4Cns8Ksbw
m4jHAoKBTusoBi92A7epyze2CmdfCmH9ELlEfUV5A7BDdaHiqsehDwFjirydQXZq
+aSa1lgedOv65QW4h0XS+utduniJTMIStoDOQxoT6VOKlsYIuPfhrgsAAmsSshpi
3tOmXBaRNcRXHUb52zzRWs1rsd6vRmlp+E2YD1DZ7s9jVo0Kjte+4cFhqCzcxfOV
hYmq/p9gP+7Rm1zxrDISq52u7a+FAvSgqXVJ4BgAUQ5D3qZItfAR5rp+OxWEH/nC
emMK+QwjyabwRHHCxR9UqEP4KlOUGiKAEkYAMWEPucrlJ/1LEsR5RGq1GkC02hsv
KjeM6YVZZT+MZWj+yCuOmdaGIcKVmaBFV7dpefmDkc5+JHxAPkzGjVEPmq/75XZ5
AVGHtVU6gbETDVvtxK+4eX6bH5sqhXBcOmT8p205vrzLi8hneGCLDcdK3xyPmtUg
31rDgshbY1Lckogp1psYrgUpqbpGoXLglsVXq+8k/klH4jgoOC5HjKNmpLIH7Jsz
76I7tmzKNMzzlKqIqIXEXpVTOWhPYOLRZNDmCmFaQB+WEJiYCJw6buLX2yjQqK02
O79JxG6Aa67U3FqNL5AdO9L7dB3nbW0RJDqCmdr+x6Zy8mZbpNsOW/cfhjKznldm
eikBBzzsZHl52uO42QiE/zMTIPFYzgEy8HQQpKCuexMI749jhWBsn7W9JrKQum8e
u5izRa7gjqmNY2hcfXgmzfPx45d3ltCwBMOtZdsiZ62nHzHEWFPEZuSZZe9sZl09
Z7UipcXa9GQtgjoMZLPBQIBqjCjKzshBBJz/Z1uo0wV2/od4q9cugqWofdgDc/pl
oxOPCMkboVe/skChlPV7Qqx4rDaDamYQvJmGn6hwldwGcfuSOtlolayhqKmE6OVs
FA7CFPEUCdZsEPdCjDFS0Ai6cRUYTXiFs9KMYUbnpaXh7sSMSjQQrwzY21G3Y2SV
vLZiwWAOV5QpzWL/NKLyH4oNEN2XAx96WklekVCNZB9gPhb8VDSm7pcCrp22Ukr7
iBX6us0ZlJWgXsNOrPVN7SPP7Scy9kr6/jaaaq3Yd6vhfo9l8Z6jFPL+slvjVqvd
cjHP9j3BwUYzD92ZWW2nIJl2XEGvzUhPDWzVTv9+0As7n75p5jJHGIMoGPpf0zBZ
/f85SxfjyTGJcHj24PHhA15EUAypKk1Fc6a851uUNCreBlTss/NKLxSL5PiYoWc8
lw560jOGklGhBHbZrc3Wt0tgqA00z4k+PCieA3C6VotvyFA0QUO3y2s8t+BOalwc
82nGwyY6nRqeyZR9SlvgGq6Z8ga4dQDMv7oOAyRL7yTqyC42vkCJEO5T8SIbTfVC
vY3Fr5IWk85IkeZPBapf/JDnHyqdDw+xIMosJXnLHGuAbQFPfCy+r1ChwOOTk/UU
PSb1H97Nbrjz6bvAa9uODvuKNarl+7qG+Uen6tdmgcW7v1IqjsNva9C256P/QKX/
71FvcqMqsHxKw6vxP6yWLBLh/lYHONy4O3CTFaTSJCrSf88UuwquIQDHqEPK4bEY
dfZgGERoQzFo+2ozzh0BcWa7mZ8Mt94/ARwKZC7JwplUFJlxm/4Qx6YzSE5Nqtpj
9fWnCd7abxk/lLZ9eOGQgz6yv/3ItphYGU9dDJYcCtX0AGwKLeHyIGaOwZF3hU1o
0PKVzX5vcajKJGSN8Z5/ef62EubeWaKMX7ob1Fd98INK8ncmgxr4eSN2du9+a8Oc
URetq8Ycf/gqspzFnhtpAWM9mDHO/45+ajU4wm8IwDv9ZZFztnl4fBfKcUG6cxuk
iCYfoxwFNWOdMiE7hvIOZuHb8Il+pr71D3eJ2PQ5ZjVhNgCv3GaJ2/8rqsydpx3K
0qrt/xM50v/0TYaRRByRTwMCBMWQiVUlYMQEJ0C2QDoOlcGxI1tU5XTsRKbVtbHu
uZiLa7AwqusU+PStEI/V+iV3me+hQQqXkuCyK1ER9BzIKIbuH3cxmMYH+o4OEUeH
FbTUSMpNMIr8EbgeUX34np3cbr7D14LUNj1+UZ0elvDNxxmHJHxL0rLgkQFfOdxo
kl0SXeNhuTqzIsjkZrU0NXoPWXZqxUto5jMPeJTSciwzieNekxBEpMDHCf/s0yn5
gbKDqTkrzq6o9Fb0VTFEKfdE6Bh1Cnccbip13LmmfcFVtUc57nzw7RHQZP0tI0qd
VnuBldvYXUK2qww7/wP25joU15o4FczzWwhea815XwzmO4eGYiwb/8sZKve+e80p
yFaGZOhNhj6hmY55ro0Tq0y3A8g5fokOSnA7eYVT/j0US6KaezRcp8mjh//d6Hw6
E3bVCNvfVDEcD3Wc+ZgiCwbRmuLMGQVUgeYi0IJsgVRioZ4fi7QTsFh9lDyvu45m
Ezl3owUIcUwBU3RDC5w//iZJoCspMfI8nD2ayKAfdaMIo92VGHVL1WaQ2Md8w09h
/xpbwCsupdpXbfXlGJQKLUn8wzRJ4Df/HVfl/rOOl/f0RSDJ/nTRmhn1KJe2VO6Z
/e8b8tWt3Iin3L822L/T27vCnEIp7krJnolqdTFKA7tKi4Ts5FSGqOhCaRDrsgZm
TriIFzg8aK4RQLcpghIXuTaW5lH7eCCFn1m7wX7dwVDtqvTFu5XOzMIRhs93dQBr
qqj8YCLBcgjq7f3D3WkBEFZ7GSctyPXjIxUlIXvvET1u/2j0hLR76sDgmZib+z3a
n2FXL6N0jjrTdiYNgeUMNHAOQ/cn9TQejUsH8i5Y3wJVsi0rU8cBTNiGycmbvfCl
cFzYXs43BaQHEaSemGzFPNBnLFHBkVsc0SqzXTd5DcdmmVAr0N2HOZ0jn9hnmyA1
Pk0QY508iQzb+34wZ3/cacc4usOb+q1nEtPU03ryetJbuJXDr1jyNU6UtUHp+bgg
W4FEVmVZWlRQrm+mU1YoHnpNE0Qdk6pwxt6PDnYCU0R8FRaCLwLZA9KCwTX8x4gm
QlHLQTFM6JTAVHmvXWtHf6cUQ19jReS/KcW6jv/ItJGoSC3eab1FwV/3KSFPllyi
5jo4VVqGllXmeqT/zo7dUS+c2zQh+1ebPuuE03833eUrOT2PKWmRSvkl+GpD6jwc
cJ3peTTLDjPq1NVYGE4ZRGu7GMXOVSmH1JpIOUA91W8QybcOGDZvwj6glGfUp+hW
KlnOYTprg2mJ/cFCcfKzB89OU/9o3mMA5EyTT1LWKR61YkjTKWrgR1GZGx5xS4oD
m+/yvzXrQ+ETsX5soPlOgpumdXpWknXaMNX7uePNSlPRfGyvUQ5pAUX3wXoUQiOR
DRIYOdfcwRoCOpxnZ4lnSn2N+62gevFJsBs/r/BjQDEkxepcwDqyDaxvdqGjF+0a
xCO/inS9tEXojrocSVr6s/Evft1HWcIKOEqUV3FcpME0xveDFIA+yzVQR5jTCHEL
7ptsrUm2rDnTzuHaCAHDvZE80mtm5XymfcOvSmmx8mdZHRaqTJrGlnz5JPRVsIz+
ucSciZ9Rlsh1p17Oh5NTR/aLLxtJwPABenFEgXbJ1PLCa875tHWIIb3PzZG2B/sc
heHRZyPo3DuQbe+8IFiyocqe1xbalcfmu7qtX7m9PJygilk0j9YtJ37sk0fyeKHH
xP+c39v+86nCaz+IXMTQJFVlQ2MsgQ95U078VUhNbd2OtwMAeVgRQuhrmVJ3ufrS
NrUamhIuYiPmu9zsJKYT4928Sjwwq+0R1lmgsTRm84/cISnKmYpg5Wp51WIG72H/
nQV4p/mRgk+Vt9vVJnBmcc7Me7U3F7eLjFXFOIbzEuYbHx1ulkxeA+JuS0ni2SGg
tWlfH/0t01e06h3fsk20YLOjTSIbVM8+hSb7OBOqiOp3OAXuFfVki2k4AzdwFUyH
LEz/lhzcrbAvLfjd6jeJAW6XBs6SZA229lbgmFDi4ex0Tc8lJBeU6T+zZLVjMpyN
AzVmfX93iTqBc+JXjleV6T5e/gdQYUb9jVpvK3K2bFbCDZsvbBSJ4D6k+Zq50wVC
O7refKjivoDvUrZi8vCumbeq/pTUSQfGNFe1oGVIxyVHehvWT4gTY4e/F0uR4mEN
kpGnt1l5MCgw77I0CJmHKeNLmEFGMSqPQhq0BKmrNSWsBcGCSlFo6sEXgM4dk64F
/xTUx/EPlzLujgMzgos6vaFuupCe2Fl3rIbtbdtbbjRCdOHEmdP1JmGeaRvRytc7
QriXa5rETba3CNwy4U7sm49UqjAt8EleBHruy3CrmQa6futN3nM3RavulV/jVt8s
CvDsQH9Ox2+T/rOU5L3dD+9VEr8yIUx+JQUIgRMKcLJ4CRN6UvxWvfrLp2OXFa9P
4MdznQenM3EsIH+ztxpGIwhY8I9RJYbgL2xFWczEGxcYIOdGL0nG9xawVX2q9Ynl
3GNV/T74hiPuZ3yY0ORz4DgthbhoMtwaIKVy2nk8P9B03tUcwHvUHR16c0pgb/j9
ZTSFNVY+6TO0F8e3R/aPz4mI5eVpGqiULhRMXD+rnDq27zY78vNEO4KewQDRjAHA
DUENso+qya1j8JGabWOvUvTKFPjagvaQaDFl/i6FWXkqiaEO4VXGNQ6QcxzUJ67u
Fh7RlLj7k5T1OI6HBNYI90zFzeh59moy0qxlVdanW+8dgakrx+4PGktaFktyBbjx
CUgyEmLJtj1FOdDK7Z97iK9oN1W+4DL+vFegXSNukX1Vfvwat6bvtpMnsTnUPIzB
cljI14hxw8G2lsCwug/rSqv0GVy6skraQUIlTSTvD6Q9tckl1nHpaynsHd754BVD
SPsdTdBuJtowblhpaUt96DEQGDHuq1kHuk7+WR2QZ0hQS8Nm7oGoubUIqXfZ2eBt
gdLsVU6JXWiqGa+qlbv0G5Gu/w0nZwB2qlvOsAMNMyh83IzYkIUKeJksRkFPZnZn
bq1c4Urr37pdSvgSiWEQMAFsOmM2/PuamnWVfCiBtGiT3Cpkjx/QxqtBumFrAS/2
emEhUjcU8t/vD6BZcfDe6dUU6tXA31I+Y6WkdayLk4cdlsFcMEBvaVw8ErlcY0LO
KObFJgLnAGjzOmc0IY4KJvLHldqnyTlBjk3Yye4DRCAjvKe2JpR1ZB6YnIGndO3H
0CgIPiQrLfHMIZG60mWG9HkGfIbfnbITq60625tXbDBTF65fLvHNfwUocGRlFmvs
sGH2biZ/r5LyK9+EHzx8BlLbaC3zn0RXtgAvnIRv2rBNv0npZYz5ZNDZ4pgJXFoP
aDqB9q2HbDPorFTtWzWE404cipbn3C0zFqzIEVtQJLSDYZkuT3oq1KWpYJEKN0rN
fGYBzJE6WzbAYEznR5CKVut+uMhtHEkSbQS4dn92qosets2Nr1QlK072DPPWDtxG
q02VnG2b9SId6k8C6soC6uWzt6G5RuCWs69udKWwgKbrx3E/PQgoXXuvQssJK2ZM
1zJcn8XLLVDo4NTeLT6G8i3CpZCM8M5NeKNIlPYx/pXFa/8/z1azCSAt5+Pyb38C
xrkEL9mt3+dGc3agWJYYHUYAzoFkOUE+2qOPU35xXztkzyDj5SyOkDG2XJtFCEdB
LGizOYooNe7wAD0Yl89MmpBHisG0iyRDKAZ4PJi9POlnnzYUVX6NLKEsfg0DeZg5
stQGs2fN2KPf0krI2/Pv6zqBwv44YNbYQKEyxHr2965NDCIsjcUqz4eZXnX+rIQl
6ESa6teTBK40yY/Hqfj8Af92lJG1/oFdpUEK+k/cqmLkxGF1lyRcfQ0spXIT044D
qy4cMPD/WyBDB6lvo+XB/MKlRsSlfuWcLjw0Fu5TqyBpJgS2RCIsz/B6wGiKFaCh
5Hk7DsCOKK5S1P7N1BU97/9Ngsg/I2E5UfmEmy7ktwaTQeh5BnlqmYVHsaMktUjF
cKKx2QQFkiFi3ndxdjMNmO4kXaK6QpvZI7iMK4gV7QWXhKhkl6/mNySvaE/wimCm
yc4WG5jNTfPa5u/LnO+eELbILt/0i2PdYRyphY1Jf5wlULkmdOFd2dzuyoBt856b
dQysjUg+iCotISyhFv7zhzoV9hEB/MR0OuxzWCNUjJ7Einl1wcricdraBS6r/Tuk
A97i99uPq1rwTHJ+zzwd2d6LXATECcay7+5TweMWmyRg50pBuanlREkHeMacC1Xv
sWzUMgIIWbRN6ai5HwSS+HDiegglIpPq1cWcYhdnUx7IrKMTAPLdPtSTjtQjVPmR
yqDJ6DOJlBawV2vbnEA/pCfhSC69UIKxSFCvCMsSI8qgndYKAMJRuMK+tPhjKBtn
zEIn2XECWYxcNPQ/Jt1LizdG/PwaOGoWjiPbW6dw7BhaCVdSi+rv/EN0lPgMKyNS
Ua5NLG1J3zFV7ANlTk7Uuw/QS1n6HFFzzq+pa1bqGZZgklQG8/hCr6X09zcLlKT9
z9YVm1f+yDu2jcMZyah5GJ5hwTogfaXtDriOPvGR+krBUUoJLGyDWOsiNbFCtnDX
IJSU+445dQKtzPAVm/I5Y/JSTqeCLIO1slQlvRjthlDB0Ej6EB1jT7DqHFRL4Lnk
kwqWI+3htbnxZA2lRuUbI/utdF6c0eYo+gmfUUln/eTvDv+AmQGU+YLmyEHzkNg+
UMZ6NsynFc5o/BL9JOKRpqZ+PYDtbyPhgm87LageBWZs08HRzIwl3k2VC0ookxza
6nkGm20TXxjSXg5G/CpdiXDzxX+kK0/dIpTyXj+GwhUBL9xKhqnSUo245TRN62pi
yENo4Eb51UxKD8SXjgz6nxrZA7FFSco5zCMfwMODnvYgE2QXY7co1POcI21L3mug
gbDLmy4jvIo1mI0ewshNq36RbMAhpQQy0DQ22M+uR8AKPZ4xj3PqPkcmr7obmZet
xDdSoNhoNXqXLb/ZpVRGtu4ZZm7AGjqIsFuMTh+f5jn4JBLEyVKK1Z/TMekbvJq4
zF6MhhdK0UuE+UxtJVFdTTHrsRDFbLbAhumdhrMPTpwKAXT+kDypr2IYX5F3MhRf
NTsr3V4QsPPna7cgYqGFO/s2jvS5HMmrv0Ib4wWnK82TfW5aUNgareEPdFQappfS
xlRp6lZc3/HPt6jQSG7RMSdgXlL2TVGk4QV0sSvYta4PfxZj4aXKIZzO/bUIpzn5
yvUfbHQhczcY5n3529Gps2A9oHnzZyIIf+kRkFX1wfKm7+t2kFzGswvXMQkiRnnL
SRocRZrqjZAV2u968XpwwAKh4HpD6L5/kWoL25ny1AVX2eFNTOqlkEa2koCnaaPw
qwNk7i07buHf5y3goS8f/qotXP8z71htck0VsRukjIqlmrVvycdP672IF62bNx+y
8apfh3FI/wN03hm7n9dsge43oWe1ZMn4XLhpdK764hA7W4PNqaDQfmqlGGx+P4ki
Hp85AesWEd4RYSFBsQEQImU0VwqCSaME+6S1nmxPth00ZNZBp09HdP3vYLMifb1c
QuV3Zbao8YQjyVPOuR2zrvUkv36zavcmuQzrvVRiQ+ao9oWdQ6XmhYaaX0OSW2i2
B8c68zQMZNWZSywK3O4dxYywbNMHumKhQgYY5gSnm22KEBtcWBkq+bFkgDTeHn9w
r5d7CcWYULY1PyiQjVV+ExwCdsUTPV8Dm3TPviqGCO+J/OBFeNQhrKeBW6/8Wq7q
0CGRwpvwrHRKQxfndDJRFEWytLuKEn++bC4u4yjfJiT8QG31z/jB2S730RDwAYul
bQcPizhf3J6i/mWR+nE6GtKSKDutrHTmDD1zoezIwhqTt7Tza7nig9JgpznJveW2
foN7EMU6PiVPeEjN0O1Ay5aGKF8WTzdSU4LEZ4Hleo54bCIXPfiCM4r/urYT5t4D
hMO2LhQIeac2XCDHSQzCKp5tvdxYDAvWQdBTjiCE8za0wO37v/9xccwD2+9nJWwK
ZHqf5xkiNrTLU0R3FkT4pUmMlk3U2a+I9B5ysfPddjQ/aVNBtLk728Qoj+tnT+Np
daJAMc/mTXhi0Hcv9ep7vuk4W4FaTcaoq/ntctCy81Mh355XNY7gObAHBFBhnxvp
UoDeu8/WzEKSowEPcdKmfmHu9r4e3uNzHRviLCIUy4qD6vW3im2qU+WswJWAlNwN
NplCYgiD7w27dSTx47LU4nXHy1cRO5Np1cnswq2kNd0RSoVqwV/UprKrMAUT3IoT
hzbgEzUVSrcd72jwwO5HM0U7dcYa0OX8vKPNeXzm6FYvjbAqzlFX/NLsGfPlvLbs
H8HvNf9Vip2t2M9sUc2/+olPfpt+rUCRUxob92Q1+3Hcw8A8cJD4kglaxCSyMDh8
CN/TUhTqljYjWwEpg1QhVumRT3ia2VTqDgVYtiBG7sYaFVaoSUyMAIaYcgL1wf85
0uDrPdZaPK3KrvRTQkaCuMHD5War0RqBTs/m4on2LZN9gR6dWD0n+T+IcBTqKOHV
sM8dibLT3J/OIYrfDeE78OFKsmkLDXfkwINFRMy2OHX+Pdjj6UEqOiMEwJ0akM7o
A1ikamDK82uy1eEAoy56BduqWIztTRBospK9bodXbt3SOmnlc80v89TGwXKy2QiO
zCSG+gyf2QrQr4noB/OfHwxPfPtUTwPtQMUfloKMQRkjjAMBzAzLyn7v54DWDcJO
yCnMCIZKqZNH9akwADihbaMOmLp/DshMlfISErv847hh8ESUL2ZGGvaah47uBLTq
Rse2xPQ6NN/5B6f3BegCHYkAdbbk5kNgIxSrXfttuxxMMhTDwEExwFOM8hbcYExy
fuITd4LyaHkd9DUc4ftsdGCq1S3xR4+5rOz0GdDsOKpo9AJAwp2tkogJOkzB1aT2
GES4LQFjgoI9AqYxFDBpRvHWmYFnzKNYkAFIWKwJEhQWfeKD0E3qI4u5ipuvVZrA
QemlR6hL2yp3i/xaj8Igqz1ER6CVWK5nsC8NU+McjpZyx4Bj4/50G7J8cTEtJJMx
N44lqU7TK9GGUANuBkBBmwEZF0lb3DvqyBHkLGUe/paG0cEvUVJT39REtjksPyxM
RCUzOEWP0Ah2n2oNhegB/d010n5R8yEN+CSG+WQv80buShIMyRHTTGCq5dc2SyxE
w+52NJDTioat58oles7k6o9CZoR1vtN8uoez5r5w079A8sQMQxaYLbAGCAeuTA6E
mYn0ri7yGg6vA/rDT839xj9XOdSNIw2sBGrUZPA3oeRQbdsaFolmO/mWsg19CsBK
A5aTpuOtvDTKOs6ioi7P3aC2UUIATrBMsOdoeR1utIqbe/3luDEUoSCafBxThUeB
qSZ7yJh54JbrWPZQbWhJSUQeLxAACQhCmrxI1lrw0uKyvhsr0HPfRTshLs7IeiPL
02aTpNBfi9Z6NBRwkJ0D0NHOFSdgcuABGY3M0gHOvydbuPJr5eyUfrLNW1jxAlJm
P2D0r3dFcA8PpiWjqEgDBqpID9sv0Wq8aMNXe6sIeh+Nf3ih0a7OaAo3dMFvblox
hh9LS9ymj70sZ8z/oQfSJlkUsjmSy8N+GlABDWvJK38iBftbh63iMt0d9IIp/bkv
U7P0ACWXjwwaITVDKl7V831hrK1j9MmnLfD273ACNohOGNMLNu8A5Dad50I4yjA6
tSBL0W8UwL6JE2fuHMU5z+M6deVzTU8csjz+h/1TKk9woi7KLtxFri5f49BNbh6L
8CQ1HskU25hKSmGUmpt8lI7neZ5EXLMaptzzJwXIu8NHDRuldU9D5szvV5zmfg3l
CC+K9q7J8aCvbL8DtRuAyohtvAf+m+QFOFiAHrU268toFV/emp9VMmW/gDGmglvv
AosFhshfWryqR0jFUunSf+S/YpHrEUBBSd8o0xQXqGDN6jEx1WCTAn9vJP5bL1Lh
2cNglGnwIXUAWDYT3YvpvjLA6t5klxR1jdkB9Sg7VkawOp00TtuWrruZ8LE7GJO8
3H5V5Km8CgTGPttC3cUv7BOVSD5O86oo2M5QE81QUyVNefCgRxfooNvziqT1dQrH
4Aalq+ZztjM8/5e2Lr+/bE73TNbS85hkCuDlmDyg5Y8+w2ncTMQZ/Or6CWAYs5cP
PsP0Qwm9+QICEbQqvjJM6Sja8cbPYEdfrQUW+F3yQ1a4ebrGPNjodebTlwwNyVSD
0PM5OGIq5F0BdysuYw8pgkBirbp1GWdUJcHrKItwO0AsyBllCQpPXQR5eIg3QmMU
2V9fJZUtDqrd1jE9wDukpSMTSY5795W7POt7/l/+jo5bRpXt8OFK4t2NpKIlSEhS
M3Xai4p8CjSMtBqcHbftDcUQ/K8Uf25TPy1y7ZVj6uUXzpruQ2t3y2w0FOU5Vshh
83xB4hqDsMRbWVKirHcz7faQXgC2J65pTJ3KuLo/4c6OxboNA+agVg24pFmXsAe1
C3m0E3HfexrbTPsEVFwh3x7fPR3ZlVQouBNLmLyA0LpQ8pjPJpEZuEyB7SzWKg1F
6iHVHHlrQmW9Cnti3sfCZLTk1h5iPBhxjky0rvjSaPhy3vogwCge0cDZxmhB7dGM
gOQvmSFo++oxKpSOXXiyQYer12PduETBWvhoNmeBmIyTrAeVpPC5/BlGSsGkI5vX
Rux8SAedIVfFg1jEwK/6N3SIpZJifXqrtz29+7tfAd8tBITGmGxdzr1s9rcPkeZf
eZ9r/HlPeNUGWc31wWClGl+aMwLGOgEv1aPPx6KbnZoi2YfxvcBpcQTvSQgjn3r0
oHAKRZvExlcsHDStdW0iei+wE3HwP6a6CRRu5EaTLXnq+cgIJiNjoNseuONdeGG9
ndNCslR1vZLk5udPSayPONLgiEsvvTKVRmxZBjJQoopN/XrEoAqtOLOkUKtG5fiI
Iw4gMywrm0M1qFx/ZYUplhbCAFzK2z4lmTVwV2qp6eQlh7U78tftXs9uD9tLhIrW
CswvKheADVhi2xag9ROzCcs20mu71WQOj6I9O39LFrKmtPmVrxUwQTdbxxlfy2DJ
DS25jIXaWn/A/QzPgUdRryIQjH3do4E/Opi0HwuEyapqYxzfEm2Q7cMHE8jh8YxW
jmhf2MTKhOwYTGeARfDcN5+CUsECUo5GtWd1ZfCzUoYCLZZADtQwAQq1G0/F+BtT
bw/QA8PHnFhQeOHftx12bpmaD5QNMXw/YrFUuUkEWLC4+Rqq2+3I5b14dJE4aheP
A26EB+c23QTN15qAJCeFvlrQT8FtWFf7FONXG9FTjvBAoejAT5Hrpu7pCuP+mXiw
oW15tFQ0qklPSsZL2RaVoW4wfPMssfpxI6+IgH3fApXLCQvPerD0uU/NeOF7OaMA
B+9ecnU+IaCWvPJI7K2+vx9bVKrc/3vL7FVbF41qdztgF8hzazeSh8/Sn8YlDoyJ
aSYhO7ksGXIEQnLCbEmVPzpi9Q9fgIwsUO6Wh1I0BUnsZq+oLJsNW7nqwzGWs1Bx
jPHnNBw29VNf7H57inpcA/jgy8GZO9zcbM3OTKkXLpq9FvCmxWQWwZyFcGgU7P0f
GCSyRNyIDjxCmbqhdQdP534Gs7UYTJG8bIIAI23Ec3vKWKXwfjBrzIjSaS7v5K3G
4Y2y8luzowkKe/mdvcvQzQeCQpj+AWY3mcwXY+dzlrXz6TfVfmzkp3B5E/do229G
GAZ+r/vTAG3KrH6JJVAsV+WgGP4MbUIiAcHBR07HjIXlxcBLIaIJdpH5g+S94x4f
wds8KU+e7rof39wSKF6397dzuP9HLUXWsoBAqBUsluh+R1HndT8WgAqcDdV5HYsm
8Xp3YcYu2zAKVMiunMNhvCM01pc43J+zzUd8q73znbOLmAdIH1NbMzUX6k68dvEj
vAo9BnlihdKr/Xuv2igbVjPACpol9ufGk5w3YetE/rn5Tz9yqzQGvN+hlT9K/TV3
M94Z34lngEc2VZtwYsCGym7NYMLM7XJ32gwQZyIP6P20r4Bw7IXzodmEzABNV8jL
gROr0ml00xQrVilgzUENAKM85KDeXfRbM649dgKPTxbr+fKxRsnrOwLrf9THauie
U//BApvSHQI8cEUCMhsxOL5eIzdFUbWKAlhjqRZ0MfvvPsTDPjEwljuSH+9uifIN
Eiomg89kSPYA21VDpMSnTRR9Mj+xQSP3Jqrac8Yx8imATtgr6vzHnfLdJ6Zt+XZz
K+iZ5FhsA10CJ9hPhOHqVN7zjwS9AK4LnMEYuxqUC54ahxY0p0O8sdD1FM7oOMii
glr71BKHMdNRDQzWtVyvyyoA1EhNPJwNkJ63b24fRmkYLusZeCrtlojgiGYGap1x
iAQuHYPgH3MPYBQU1NioZb0v0/zNcrUMH+vUX9l1bt4Va9fNUb+NQkSdFUtPV9yP
oAxLa6JmuswSjkNf4OF3gCubPCifmWF8+i0lF/kwbDr5gzVSD0IOYJBt7F7FjkFf
UYP4HYkgtD1vVH/OHvdtG+aBcO1SJ1xIKBhOpLoK7+AW3M+mplSHhVAT79zqNHZ6
5mYVBP4klMiuYwJPV+BDDS43P6L/mbkYHNRIQu4okBvPLiCMmc1o1ZsfX3GPyuCi
ueT4ZKIW48+jZD2GrYtZMX1wuSvd+mFjj6m3WotVxU5g8MgwKDIJqBIklDsqO2O5
AQMlSIno5+4nxez1IXqegaJoylT1XTSE2VAxzCQZ41IJhUIrNuuss83ojvqeMd+c
E2YGFM07U9wT87lswaOUmpgZtHRrZblZl5i6H/HuspgIVp2B8M6jw1PMiqr/YXMs
0ODN4Et0odKTGAEFMgYPUQoGSMt6iw//tPynM+DXRNSXXNh6ciNgTHUJdMJb4IoL
/eXSMtAfMoSJZsnAgaNAkUxtcNCzwwjU/4nixu9Im171aaTr4qaFpZcDAPTEpmC9
qPEdNNQtJlklHcMeXM8ml9dQ2NOTdf3Ur0BeoWkEBCZ5qjcpMOzdYG16IBU1bcOS
AjOIY2WnR4XiTxFx9wfIn5JHaeVz5ZGzAiAljSzcCLz80hQAmPRSab/m83rDT0On
JpuVntkklcwea2IxngSTRm25jltI7SsSnO7yqm0hDmNwLvPBZybDm7wG8Bf/SZDz
DZhjnEjlfzrJYZ482tD3++NnBZPP/Q/8lqA+tvpVyRpbxit+qiqgbuxWMImC4FNa
haxbQL+qvFv3tKzm0VIlDMh3xr/ywgomumFIVwkK2RUUala7gqwhRDcfIvnyVGbk
KlyoeFOAn01Pi0iX54vmO+uiVN2lF4BZojC8rHpnKQhtMMOsebth4zD1iAVXbX/O
FQ6K6YqRe3OuOfiIAG32VZvbMI8URQNRXRC3/taSvvw0CIsu6/63BCfuE0fjuIqD
mJN9a2ORd/Ln9LD4S/I0HJ4iuCxM3ZBEozomEPQsJhtCAXsEQy95ZKMVDYKfWwwV
vWm5VsY+e87P12IbcikR2VMFpawietlHPH92H1TBA7i0qIbd/7uMtvPi6CijKzbx
yq6ELqfoC1sLRiQn1P8nxGslUTiQ5BdJb7tIs7EIVk1McewdpOzgChSnYtE5nSJo
QIlfyYULraqAn4EuCJwaF8zAuwUeG3ieMZP855yWEeqiiTdJ+UNARKhjaYfSD4eY
PaK1MLoLQ8vTs82GNLyl0lTs4Ik+WMaCxfN1IQ3k0L1ZUqXZFskOcZCbKIghIOtU
qA5pMEGmhDyJUbM/6z/6IjBZ9i+Giytmx7SYcp1cLgU043k3id1PH5yJtSv+3B6a
Klx+PemyZPnKM6zwcuB+7e25unGG1vu8ApneKqCtg0P3SKBpTUhYgHlRo4ZLDFCZ
+0qOIjl0+JdTXEg9NiJrNImlhlWrhEH0P49Mw5IXyyXvic3TkCluVFJWci8Cwzhg
M8PSX/l+UY0yQubztveQaz3Vu9F3WtiqRMpT8dcv5stDk74r1CoMDQb+jnF5V+rP
TU8+pR3/aV8FvWF+soiy4Qk0V9Ky0W/UwGPq58PHZo/XYTEFQn5SPXWSzRmmGF0Y
DmvO+iUE8RylB2lrvbqAr8xzNwH3b3//k8hQqTNHDNuaD1TpYLL5DHl7w96WOu+P
uBS7sT1tnuDcgo/peWvwel350XhMSOvhesaMFrk4v4yvPqw/KoM6JyqznApK2BzM
IdDhvlo39rXDHmSp2bdnPWZbOjdaj0axvEg0rwnW02hhEEt0us8exjglEe1Uw8Og
wa1oWW1x0Zyn2s/P1K9UT1lNIIE/GlBC5w5jQKIHxRfjtD3WSSVIngWKDwpp3Eln
lF3dO8SNw2H7VgDsQ1JIpfoZZqJ/YhpzsYlj+UgpD+1qbqqckbdJ4wsMHbIU1NnJ
eBM1IgfseWj9/lsDfQ+KIJepCiIU1NTU7sHTWMYQEcJTgDoPptP68ZD/wbCnlYb4
HMDn/D6S5Y+x+MMzwhEpGgQ06OIhRaI221A+0a4OyaGDuFMIvsGNwLp2EUDRVm4l
BtefEouD9VvJBIQOFc3RpLSlqpfxwKtfFkGMOhie2EiU2XAAigsRJLwoLaA4RCOZ
IHkdCwNMk2c240eTadA9IkT9K1FqEtic7jNen4Ld+iOoRYzL4SK1evW30dzdODv6
g+jUlpBznTak2vXjJK8vL1vGV96AOvNO60Kj/r9hJ6+3nDFbjXOEdCIksKzhPDnM
MFYI3XjO8KieW8dXt7j/CIuxInToCoa03tw7wNNDGDJ1ow7mcZ/OqexHj3mMPtJv
GPtsAz7RIUbthng0tywMtnnSV03GCqsFlTN+LxF34m+gf8Fhm52khnO+XCL5y3W9
MaE8U+sys0mfjtAQr2k8TqniAIRxbwpHdnsV2XGik0kLyY6VIE8QdvlboYRjrJnM
V+YuoDilDcpzTTxPPRD+vIH5wJO9qpah4ecPZ3MrbKq4RaPM10k83wYltCIOW7fS
P+B4EPj3ueyeLEchqtYlV5v21EqE+3Jo40evCPb/N2KZhu0rtnkvWmfGqdKlQZX8
BtajToMZzQwBfgeNtqbWf+u+N/T6LYvcYP6TI9OwOPaAOuKTQbsR8JKwJ0yOxP8m
Axa5D5dhpDoUTL8M8rrB2eJQvYoON4mtIJMrxhAcaBrxf2UJ5z1C3ElM8L7L5obo
1zB9NxfDWXszlchOaCrEo7N8mdpm4drP/YKZLkzi+/4oCbX8hAgcKsujcj5EMpV/
arNwR9pEQENNn2fB+uy/oNxHL1rTB2htMXK849Jy46n9xJmxdX5ZsxP0JDGhBQao
lyTTZZZ6wvMomvfcFZVAhGQ3alCKxsc0Eaqal0vTJE9x3+7TvRYY5dRyni+PDS9a
bjvHxOdUtaWTU7mMynlM+SGGKSdUxsS+4yApryapre2LLC5EvMvZAxCGFlWO2nQx
zOo8QAvuuhqz/hMuXwDmrq0jINdvjH631OE45qc4h76x3nqnUUVwmx4HahkwezdX
EBEOIFmcdiME497Qd0bvoqHPMPmKmjwO8F2zNMaE3ydl+5C19RKyd9bNBGqJb1LD
JXpowMFL7urcLxMzy20mLk06P7lXp/OeFQKmPuMQKNeeNaE9RkII1jqcNeKyDJ87
RfhcMgCk6jeArGlJjiv2DqL/turaxMv+TPTXraApv2ph5OS/eYyNtxqcqDyPD8wn
UOT86/ASIKft4X7/8icTPPhK/TVJ4a0ayIQlihp9Q4u7SAna5eCBoxcBKa0npvK7
MvCWkAeWM5gzHRpnccDovihqxbyHUx42aRjOGnWXaBCn6VGKu7zpAwG7lbSexmM7
4LVtg9jAUIDga9KmCXBKtwam++GKVBeVtW5BlwI7cF3lndSQfV0lLDet2UchTC1f
C6Uxqs908kjGV+eaiPXkri7PoKa5+/SMppzaRBXvsSM+CWkdKjC8Ha5e7pZ2X1yu
NOCQhmwCHhV7K3DARVJ8InhNLNipQvcgXbETmp+5dgGSgAtDFYtkdDOWoVi6W96W
qOwBa2QSTYlki9l+8+/I8jHHgYLqgkCi5XCcA5rtJVOi8E8UMp4sh6UBwExLQuH7
tXMNylP2uw4ROd6VpNOdfa+DWPjBFXn3O4ePA5bDSWWgA9f19PsylwUhCj0lrhuG
IUbsoz2H74Na9Y1jO3zEmC1zEhxrm8Q7I2YWdmV2mSdOTCb0CDhlTz1SDKVOKtKD
tNLMBDGyxTvPlxcQF/k7JmaWUH9TsWUWRdqeR96UqNf7hViyItrZ4ZHP7SEUkyku
IxBL2Bzf9RiBgLvCstK0CjRYLCoMfK7H9C8U/+/G1fb69SDiDNhxYFv0UYOTG0oR
sVQ1chpAwUc0TOPE6CthIsCJWV57j0Q6Pt2t/PWmgf5Mcwcpr8z9fzK/eFIxF6hD
GDwGtaR8J0jru58p7Jp3s3Va4s/T5bCCgt4V+3k3OVazreE7PgEjd1yNOsJvG39C
ft6MYbCEJn0b798i3G8fmV0NjY48EfDdXGKPzUmymQNzavwhbhPhkVLxXjtWJpJQ
rgH3xmwgTcDbk/gi0crFadOFPKIGOXPTOCq/BmXAu5Ce21dk9X6zwPxWGHUSpwUP
Xsvj22bkIiekodkHdsQjGIzfyAtXOJJn+5TZiItdJ2f0eLnFgKqqI466gWgoNpz1
QSeOFk2bMxwEROvyQjsS1V10aXrQ8dbTISQPXAbZgXdm69OxyIzAB0plM12FUmWC
C3t20/DaVWevrjGJGf1PzLO/7vl1mV2L7XtryAWTE7QRa3Z6VyydrVSaAoD7KAUF
TVwQOCJjMYXyFf1+4WD0KJj1Pd3gRVzgbrYyt6P2Sx/YBFUDEZm6tcS8nSijUhnX
l+ba2gdzuD6+43Qq75U68htJL1CX2wBxBZFXn+eKOdGlK61ZN4O4AyXYhgmvNdsT
dhd8bPFe45a7CWEB/hoz9ZEidjC3WMa4OFyDLC+EXikSJTNBjW1WzhlnNkXmmijp
Jc6ROY9U9PWQlXFi1hylH/V1vv5aEFRP9I43MjM0t2zRhFHFL24mLtfR0h3WxQ8n
6j5R8KVEQPChT4G9HJhUDS2L0MasnweHOxT+nyT/7mi6K3s9oV5jACKzWARMDFnR
+k8EI6N8EN8pPkjjXByTMxOWBFNGLoXcNyDzxHJ5c4jA6Co2x4uQgXPDflGRM+kT
z3edqToSdM9qCwe7HLgsYotF/Ivb2rY98nl5gVNIX3AUkaqnA3mp8BXSPkP1H00z
3shUygDOiQAqhu0w2DM2LXS3QAUyXJbAYbTbXCPyKLc1r3BIwYvehbuNWTFVzVAW
q+W6+mE4q7bU9UjmtUAIvDQuAU1zYulHifKJZ4frH2L6fqJmxD+aSi9FtnL43icb
wTVDcRi9ZLCkEnxW6lMLXPT39eLD8ls0vIVCeI0FGaptSPhH/olgTSKgIXfdIodn
ALNZgjxQoRi3/PPuQqdhc90n+aVskVcTdrE8pafR09Etpcfv/rY8PMlKRvChJJ4L
Cwjuap7TCjg3RKY7YNKf7kJ7MikBrNTgQ+VUGR09fwInZWggt7vEV8wWh15CyQn6
BhMugH/72lIKA9qf7EcpL7nVBjDhbGoBS/BxF5RqpdJYt7TZXv7gw+sMQmws+eDg
rnpfOPLSL3fWthWwdOdQguAV3uX1wNN7GOkTLvMGdSmVyM2ytbgBGm2xYKFo7bbm
P/ZBg0ehfM/cCzPH0vig+w63aH+CMHITos8r1s9LdH/7nuGHKrRP7+NyjzBU6CvQ
5t4LdsDLcQSaP+i9rOzk9+E7paiQod8b4AOmUugW/AiqGtZ55bWcjnMkqkChXf/n
9g8EfOq8bDdd/V2+Kgg6C6ZNDcOJkuF4ooZQm1E2dkkvcOJ0epoN0fayOtwd0V3K
NQtzftRBwUTXYYpjFAC69SK4boZDwhG2DDsaKB9CVEWCTc2I6hCALxcUHuAIhs+e
nqYxMQEdaUZLmR+24E6AZZZrad5vuN3wGubz2ZXJ68xMCkt1miYmIpSbqlA1ZjIV
Nvwq8cdq9BS9fERLPDCKW9i+AUF/b4ik16wYnRu8K81cEVU+ZLRXMzVZNARqIpHI
5YqLwUfSUE/VMtr/x2HoAX0zMaj9rYENEFR1YmlsqWJMJi55KtZONpTUpyQqzppF
F8Z7aap/HtTFtyyoh+Bx5X1lHcUVzS0NgQFgRXrzRSJTNmSdZgAnMDczT1E3e1Kd
Gal8TWTd5VNq6eq16jjPwkeTSvbt3Xa03uZNiP/DajhVo6Tz2EHT0hWbkvmPX690
B82I0irummUpVypBZChCdMghmG2ZMJScr06A32ob3Ax5OI6dKFom9KUk6yMJu1k9
sztuTWU6H6uviBKOmYPIlzXD0Z1GZWa2txwDNS2zLuPIdFiF+1Qb/aAkYrAbSnDs
MCj2ud7bddROmNztdH2moOYDuk8ES5oAe6iArxMtDpjIbfQnYBIvOyV7aSR6mbpt
jq4Q73L/HQQEX59aKIzzdEhG+dv1VWLfUjac0bMCFNQILIR9O7rTR/p8J4qaxvNP
a6G581Nv1kOSLfL1jnHuifaAJwfTyiR7xR8e7D3XrCfoUbq3HgZBuiUxK1bYOAHp
SeMgNzj5V0fn28dVYeEa/+2mTQqdMY2kM4YXlRsJw81G/Wqjs/ms13qKlqNzgbX6
Ss0enjTMZYV161qZIY5eIkVR8UnfohM7YMuJyEXlPc+mVu6cfkdH7wrZpSlwnqg/
ubFdrXk3LxwexNrMLhrGUSMXJtJMG+PaB3IEy4LaQFdNkNYjWLCfjNO6tn8uwrV0
vObvedopOAtnLE5PKI8kwsMHlsfYKklYQhnewRKhVSpOdZ6wLgPQVWUP31wSi23I
3zc8rlCjf1DgY9jtjUqOzwQWctvwygTYpsZzUO95Ur6HHzugqgNCk9EnyhAJmheO
rXe6BGb8anxpJUM4C2Nrakuurjg0O8jLZQSXWuAYweYBYbdNawVN/MhctMLDijSg
8shx+dbVF91SU0LsBO3rUVFpjZjN6ppgETblBGfUncivR5hab7mXYGLWHa0Nk5ZH
91qsP5NhjRDU14vKEiEHvk6LyAOtOY+YPDwjfC6k3SPQtn+ERYqI+hLdJONQsa9C
RPb0Vn2fHxzmICtroNte/u9wsxO5ShKJKCDd63SVPthzxKbrGcYF8po1seOfP6IC
T+CtX+dwjMZPRntRlLI6nrWiBDXNPkOylGoLllndyOeOlfNjUTwDHlTsS5Ecr7wn
EUVXMlgPqUBErzDfiV1BCr4uEnLdajCtxZ8sJrA8MI3OoiBF9C4VcxbCg47mh9mE
mUFMmszbqdV8Qniy4kmyT9HpTQA/zLbMFPqQM4QMgBFy/+1pPDl0Iq+o53O6NloU
PDkDzVR8jtp3shURmRN6Bq1TWFEgBRNyGnbVyBGr8QYAIxPe+G92KtNt+oVnsfdY
vcSmxO2lId1hmJJLx6W0rcFx44vyzXoCocKHfTEyxZ40QiwghL8QK+ihWEAelvT5
ezeIDaXouoIQ6QZ6pF2aqQeXDbij9n0waP1aOl3FpxUrWJJtYf39G8RJCHrnJJRO
OJZxlukblOA7BcEV2YME9txOUR05qquFbhRsG1E6JTdNb8TP3l4OwcxJvIySKNJ8
9AqkY2Wj2BxOAR0JpZD+VEOQZ6IuAdFvP5d8UXZXcb5lVI45Mbd8z6vsl24sbctN
3quVBHRdVLmlP/P5q6ix+XIJkRB8WOFiwKSnCFl0j45YvTiur/OBv9rAIPjTEQFu
IWEcGLgwN3K1+ZEP/5AArjdzjZ+mXhhshpUfIr1HEj7PjzEM4Nl2a42FTEnEA0Us
+VAXpQAnU8gSdiAYPWa19eoQS2Dc3KGBGaG7c2EA4eZQA8Zn13XcQdU6R0ZpK7Yw
+XFHwv7w21blcdQTJy1xMUiVwckM3DhGQOXRBQUIM54IjVuioduMKswLLIiY8pWL
nkmSe1sq1sKs6a7H/EAk0gj1CZFEkEYDGO8B4UvFNd6DzEAjNmt4O9pPKClXzGI6
Hv1RlWfRiYqfZ7N4S1YjVwAVkCX4MEBQcV35SYQyYp5lB8N+kBk8uyIhwcjbqGmS
6N5HMt4MrLJpIG+ey3knDak/8rXI9Zanbt4WzyaAdKUBNjh2ftjnue9ARvH002LW
/RsDmq+Yx4DvPK8/wyp2bPjaMAMK91OI3gbRJmIX8syboxqh3rRR/9xsSZOTJxYN
X16W8vADdLjIwXRT2/QQ5aLs9sxgpSg3eSHOa9JTMzlXn1fgdo0ERJ04t0LUQPuX
z8K6polw4Oo9kBYC5/n7KK/ExCQXM8ckxXqZp81DrgfAg0BJRHeLNyh2tycXznj+
bgWuJvAeRXLLQrRTUGjrVh8WW9v8zC8y+pK5trByPjlAy191YyfmFfsM55a8jmik
WiEU5Sl2t8za68ozc0n4gFCpmc5vkPhsdLVV5qzpfIZiQ+6g/FHYpaSlgLESb6nl
WBIrtkbYXD63rkYS5DHcsjAnXOIJBXXQGnCA1psu1zrwcG5wL30bHLWFZbLZHNG3
rL4Yi4dnwnes0e8NWiNDQosfjrW1B6VVVzFvi8hwgpuS+aO6O2Q4w8Z+SiZEiJZD
27iykQP/fPK6qUEDu0viV34fSTuu6L+B9BdGPgdRbmJjKw1LwdufvbsR79aO449x
mjAxOKq3257enH3ngZ+7h6b/GRSdj5Q03jO+8KsivTpFs5teBbRUUTNiG+ziQd9J
JDKpkmXRbUASpJa7lqNupIfkTWFFDL6eq7ThHX8iEVgGN0kQ51KV6Mh15UTkInbj
y5x0NQuJX00h8XP6QCYeHkkUb0+F0IZqZCedQAMxcAfQRCHvea7sEV8eEd4OqTdc
4MDt7UxqoXf4pjL7ifKpCoEhkKfmZtNNqHiq+lby2B2jeRUwgBoNl/oXkKY0/IbY
JDOW5ZDvsOz0t6tlSnnIeNPPrpM/aEVgVQ0x/9p6PwzukfcYLxfd4msIULpxB3m/
mZE6oUjV/fhK0ro0Qa//UOUQi6JoHrtiHAPbBCWfLUq0R69myX0iPWilQv2x5j9J
TYgtPUVuxPqz3mpGAxPgcvEeNABYIc/6AKukwedoDKZ9c2Piuh/+p6ggJZFgUmhq
p5R1Dc5cQ9x3HkCpJQSOYjRgEWblO5NYv8O19w+l3Gtz+Eg6+DDibvPQcxWCLFGr
75BlYD1P4cgAQsZlzS7eIpgku8fvOEgPRYKUmNlZcSJfRfhhPHrnqRt78FDCWu5r
2jHeoQaVWV9y1HbzrVgOMHkj+nwlSxpL+Wr/d37QnvvoxHCCFShRcyPvPLMuZlpI
9bqCC7rPt14S9HU26fj9rvD0FNtcpZGWQDGpTB1OfVzyPnBrMv94eGmLpSR4Yq02
ZGpLddR5LyNZc5hu+qon3FTwmh00vS8+qyI47XfPsum5UBZZ3jG7FuIam/isaV1c
PcAzPEcONzPqyZp3dV/+b/wRCIf0THFvmuvgkGM92dGBK8nVP6epma3fN+sdKkaV
2bv1Beev/s2XAm91o6v7M+OaSeNflXHwAnSXkQ8P2GOb01IEgd8OYhLjDt7KK1j1
thsQrUOHFWAnHKY4oWSmvkELHLrf3HwIKDkZ66by5mUQgcDpt0fyNdPsBIm6yvld
vJBG1sgahn2GlGnH8+8o0kq9sN+GpKfgf30s3ebQQcGocn5TjGuch7ptEIT4q9ao
IMcFp6Syh4/82hnlM/jnxpVqe2UUFeosQtTphVDEuSS4fO3ZfPwHWiICWrffLcqB
0RkU1+lY8KeiYo8dHXqc2/9emX11jeOHJAwjKuB5LDP+y5BJFUEwZaKgE2PC14MX
tg0JqDwIJK3awCzjz4hyFvO/KObOEDqdIUpypGZNA7xo5AQsack2WT6DaJuxz2Nv
uhmwLvy/wncpU7qp5V5Y+kDPYDXzp8nCCf3ueQF8U1UAdyug1TTueJq1dqzAM8oO
UsasBYd5tbM13I0MrbSN+bhh5/xPVbXB28UgFgWkf0L8OJaiccCjTSgXyZ7mXqqz
TwUKKPzympexphoZZCvThFKzuVyNTIvZS2uDGafCLgiOviHkf1yeXir7/Ozyfbq4
McJf19KDxt41ewy/9HkEG9f8iAMHwOB5iQJPcRgH16hJtWMZlSliXY5PyAjsMqk0
svDxhHgtE1oTtF1V8AWOgh6VWJUwcmuFQCwbqBfm2ApUTScXrxnQG3cUG7D8YF9O
wYfX5wQI96YhWedrAcY5MYCFw0VH/Gp7Si2qkWhhkvw7TodgsZNtqsaNpcdEyTUx
EZkIlfZnPfjcoeD0M++aJKPk0sT8aHFsJuP2wsBCHNJYppiA+IudZJZ91hqQVbV6
xB4bV5WBL5qQEBNSrQuI0tHKrL2oFU0W2lYjTPx5R1Td6/pSHp2+ADKS3HiGVQne
qbIlJxOIN9YqlXiUrE+/jhDp99Idhw6NoDpYd5a4/kRMlBA2VVzXfj/+bxPAErvt
Vyx/OtWt9i2HX7Z7Upa3T2BdIWT1qz7TJ5NQQgMp4nFN8xV2n+DYkYIpePiw2o6p
nLaxJwoLiEeRfQjXgrP/VSItU3dqSCmQ3zIYYPq8hWB3EcBWf/n4MXADW2ZvxrmR
xgYxaZmiSdDiGngnt9wur16hhAHKoSY9m5dwQ3JoDAWbSHVkK8dBPy9aLMjolOT5
XGF6/2r5mxVaRQBegEAHSCSxrUlwxwxNxvHM2lTSmmmjbfvV5pvNno+iPcYJvrQu
YIpqVOqpo0D83DXyo9lItSONo+Irf4f2NrTQ5Q5HkrdXQb7EZVZ9hUoI6rYDn0S/
TRfhSvjWCb2ppWAKN3KEErRlXx5jlaIX9qwL0jc4yZNZGY5WPHlWv1d7/ucSEl9T
EmEMds/4P6ihDRTgr0VMKSXHdGgkuIcmbl/+kimRXYNi4EmuWy1Lc6V+XsVZfJAg
ZAr1Dm/YLCHZEis3f1c+lz2LvGJtlQwn1Gv/CH7z5jdTMgQgC3s/7/MuYVoymlOd
/QqHDq4m0Has5lREZVsyTRyYMK7M9RpRdN4FzWJvH+TVr1fBo9NqwV/Ad6r8A4qc
skwK1G6qCs9J3nYAOtYRLu6QDb0192DUba5+0lyLZil070S/N7puNF5rUpAhKSG3
vc45LpLn5XfNponkp9DPMjb5o+OtMqN7RkHWFeb/TquA5Yfz6+4Yl2dIuoh1+E88
Mn4dn0DFaLI19zouUZoBNpAPEe5nCqNVV3UID2fJQ/m+st1jR+oooZ+JZu25fVJQ
c5VoaMcTLZRnH98zg05WgkGMvqt7xpnAugaU6tBq+UAIfWZ9UIEfWR68Dj6KbA5H
MBemsm9PXtMXd/sQoBHV4huB+kbWOf+F8/T7kJjdJCBimZvchdeQ+yLHgMAyNLLW
i8JObDQN/SU6mQBRzQ7Mz5QgMYERSb/gwJ1+6LoGbbh72VcSvioMPAM/KsVTrWGM
mf66B6sd2i3+33SXzSjP7orfM/uNUL30Ja0JEQ+2Hw4uQmH7PtatSHjRQh3JmHY1
CJWdGPUedsFYV/npiQIreZh58vNJM+OdDzbwlM/MDE+HnoZRI3WJPcikygQovnLu
jDeowi5Pp8ZJ/O6GiPRdFOrL4/4y5ZZM+GgX037ZwqK4WR5U60fb2Dvtn2wBLqBY
zSIR7oaGvyQZd6fiLZ6kXOZ0jovvSWCRPHO9w3UMczesiB8xpIiv6hdWb5XEwUu3
vlhTewVb76vgtGZKd2EkYMMzQJEoTKMJixqMcSDhqkxkjGiDBoxGr/Y87LuFgDHs
7MjC+64Mm1Foh/eT2vzlGP+zcYfRGh1WneHXUkyxBPwikrfBdMA345T9vJ1QGv3X
kwKEMH3j1Gegc+d4e0vPa262d4LZKIDYyEkkFhxv5CmGAA5yPYKmK72zhapjcICF
geojahhgvN0oVARku9VM6fooFjsazSQEecPPNaId9jW8/cn7QMEyZgrr1y5hI26L
gHJc9+2LT6uMzdT5n/rC3tpWleB6W1fk5AP4Mt3IRrySAU254lx8ZE+dp403+PKu
8y7YKAVxlUwyYzdhlcjoQfxA3z1w3rvXzSo31BznfQwoG7U1qmj/JMufBmEBv1Eh
EM5baobWRuGlI5CD/HbryrWuL/oceKY8DR1X82kWN3Jp543cOWm8iWVwnp+YkWqv
2WoNPnKXJNuXcjN5/h24YT9Lt8OvcyCQ//43VlOE7jrLpC9eJsOdFaMyLH+7JzWD
IvcTNPdKCCgDckU6ONsGvpZMdGu/9eSmO/CMZrxlLlv/j7AmZp3G4x7GabKC8KbA
+47XEEW/Uta/ZVNNvLu5foOQoOGmRGM/3wORAKb3U24ARNsRbJLbGnvWCQHOhP09
PG5NezDjv4Z2CGyynUSQAkg9cPgGkr511gb3bfml7N1Zken1XMK8sNKJ8V4/xo+K
NnDDcB32B6ILepW9FBhAM564iIYUPDo+rNBfrLJiza5oSZmmZSyOfpZejguc1QDg
R4GLjSb80o5IiW9VcPE6Pgt1vhla+uedvXvBNbqt1OxfqrS1yZt2JJX5CzEr5wB/
7gTZQkRT/KtZETh3OvVNxFuSZSmZ+WO2UxOP3jy8G2ZONTFjAGtdVVppqJQGkHZ0
0DbWvidfB9zrHy1yNDW6RJ9UKzO/9Ru54UTfsWDKQnvCxtQQJxn/srpP0bN6wquQ
myWawK7U0r6ZM1wz0iHWtR/x0hv2vHxLV7yxuMfD5UinEcRKFblc2MBA4/3WlAZx
e1vTOZLUkmVJQNsK+pz7SVO70gZHVzrHL5tETPeB9wN74hAph3aevvDK0Md3L7bK
Nh3fcRFQPNZMMvzmUn5TuDHQRiO2lCeM21Kw24guVfXmnRpR/lyRfN+N4dip244i
1opmYC/wLcNe2/REBYLcXkHBKXtvqmykQLqKPSQyyA5QktfyWOe1C41AeWI7VeJt
0KNSfqvxKYlSOmAJDshl0si7/X4Z4aEHeI2fsr20dO9rpec0+NVFfxO6r/+1gSkB
kq2m1dmp2SA7n2PHL0wQsGAsU/Mq97XrnM+/qE8hlZ1VOtzL80KXFQ8P0hkerUgR
Me74TZC2CUx98wPUxuvmzW6JkEksE/ao9t8CZAISOzvoT+axI+xMKuEkTtfTmBOK
rnXkeRRDt45c6WPky1W2vK58uxV+aDMtwDYF+JibWZAFUD44MGPT58v4nnowqPoB
Wt79oV/rJth/fxy86+ViQ6yqTArWL7hK9n7fM0NJe5ddN78lUW5Eps/i+HYmQoJo
Q9g7k0HhegXeG/66J7DOUzQhdGml4U7iz0jCqWjCxsbWyv0APdptYs7vx5SGcEep
2cQaRqbTsB7IhJhLretXkKbcmiWMe9WplCluHTHVC3e1N6VWaDxxHRvIeFc/AiB2
CgETAPewHOefKD8ltBCFdZ2rctswr6A6CRDzpRfKmIVRmWM/HQ/Cra0JCbXZyfB2
N5+sfKVJGrT/+XY3BYUX9jE66FOJyMxCPDzhYjlxC1uq3BQ2lE+nxdE6AnlMyTyf
upErooOOjiDDaiizZSQXMrpL2zRl2LqS3LFqfpxU0yJIJiOUbJyXIEVDiEPAY67J
j6jfZU5H9ZcPfe2EEYij9yQMM0cIGsCGWaGmEgMvLW0vOH2vEtGqHKtnjQr5Rt+C
CVFhF7sDyJVDXFN6YlrTf/zihksi99jdG11SB5sHHGLBi4O8Ob9nHlMI6zKgNZgU
P9PX5poDpjaDc/3QK2fgp7jVVKvDW86Vo/ZuxAnnsZ+/qWEQBHvYDIJfNw87IFa+
9MNPOAWRbYa5MVPT11vhfM2/oflfB4a8/GL35Bmyg0ucd8QWoCTWcsEADbB5aE9d
Nc518glnvDge9qpM8KT20L4FaSlVFHqCQ51X8MPr1CxnL61z5l8XfLzFBOiQzmSE
CVCxBXBT9kNxBOAPYuEDQHpEKPh5PSgRzImF5xQQPwauAbbRcQ2Nfh4Hx/2pGm5s
3LZq7jXReW/TgPgC1KxUj0ROGgjHNQ/ljls102qpjO3AtrjHqsXD1iMbuG+syMAQ
u5oumOfhUNYiSYnyDJTkyhvnSlWTUqTD1XNipzeDUjvXcjyB7exfJnxQh4Qeo6DD
vs7eD6WXPVNfCHcVz/1CwH1ClBeiBkyO/vtJduhLeCUCmYa357rn4GV7EWfzVCBN
b6HomChlip9iTWVQeJ/m+PLE95yjrP0sq6wG1PE+Etqz8xDA2Wn/44NTymQVvsS8
DjTINDaofuqf52bfKquUvclGT94Dt5FB2nfiT4a+hJPi0Q9/JYYrXvFwLaVN0USi
OTI4xOy71hY/WA1L9G9aptUPn8biRcGHttbWNR31BHBap+2yzqntqqzIGQ33wt8x
zVOfhRwdk1jfaHKrLrRMzuokEdG6cxLNNJirQWk2gg/spHwvG6ioSrenO/rpLz7X
XYDTVddFOQgBi4VWyP3is7kkEs02U/ERi3ZVGAGJk51P7fpe+LKepfwl44NLQCYx
OzUtLXsqPjyvMGVkyhPIepJTq7pruictmpc97i2WLHPSjurRTSyFS8YbfQD6dEKD
HWZlWY8miirJ5e0YbWWcRnnU9MvsHTi+MNK0D5ne1PMed2cOBgoLYdXd/XGgGVN3
X+eFDlkE/hfWZssRXCbBTug0A5sMoK1Hl2xXTv2qvoWBvl0ZS5XAVE1IC4D9jrXx
AHy61bhT3N+iBs+DNp8nHSkrgZkBczmFlnGTA5IvDjJRkaPNzLhoJjbpRWAmsgqI
RxPOqgVl9Dsc3SgZNq8QQbjBow+QlTnAr8FFllERWUjoBp+SgbpewEXzEzaNDfO3
QN7rxVBJoHDonC+o5EB1bwlGbASsanUfqYSgIU24JPfcN/aqwNwqAN6N2XORAW2b
0nrnYDEycOcHo27vDDIMNi5XYLU2uqQWrgN7OzfAzxpubxfnQYmRnVj2eWkRlie0
QompFHgPfwih+hNyDe5TZ1/UtzpWPOVrwyc36yEZEtO/QbHguYVohsYRZo/VRQCd
jSxxFxTB27NyV84qq93ibkKK3PUrXmcwI7RB4rQfktmgWle9miwDGu/z1F5mqGkX
accC/AcUTxj+L18H+5RUQ1xIen3kfyv9u3GtFc/7Z62sC12heaIw9J5wKSsPpcfD
qkPX1Mn9TaKc9mrGF5wRtBdaC8Wircxwjo5hzHOZz7DDD3QtalpCE/Twwo1wJL2D
daksZQ/BNxom0DG1O9PrgofhDilPHpZm/istNsBN6nzDZb1HzluP08OnbKn1uxdg
Q5c7V5Utw1KN+pYOXMRqPK+pLTRbrdT4enbIP3FOCPH8F9MoouZ4Vq8fDACEiG2w
bxiagAlRBo1bNjlDQ+XI0aVjSpy5mGw4g9tPxOxgWSB8g/Hn9RKIdiapU9DwKoqD
Vsb7ZLvRuQMyixgnGRWCIV8YFmIApkD07ET9VY+CUrDBU6kAgumWB1U1j2CasSAN
AjpgGoXlbBxlRc6rYSYCXCua5A3Nr0CUVCWzBQwaWeYQDjvty0MKv3tHof/D5Mkx
gZMtaUDcw+4nvwSU6NfIvq85+3osxmvfoLJrlCaUHhJZIO8uP8aT9iCh1jnfgSJC
a8rKJaqZKBrXn4kmDAOctgqH1J4tGDIYwxVQWTeEDGrpaAscb9ir9EPnec3+TzRJ
l0tZwfK9uuWMdsV9gPgcbdoMO3SdPi+DqxS+t6GggRpPu+uR6QGSuBewUxXLnMFZ
fYC5EQUJEUkZtM3txjXwMXpZDQzpCCLQKiTD4e5PcCjaHBtYVWRdxc/datZbjUj+
c+0ykdvU1nMpsVIZ+ilkPjYGudMSBZy1Wdrw30cCgS3Gf9pSJGD31Wxdylu3wx/n
xGAUiwZQIV1arOeeMaEa0LusHVqo9aIEMTAMoq3iP6eW5gx6G621IU2C6j5N9mc9
zWY5Nsd9JDO5jeqvv8e8MmYkp8b6kbd25pCN4kPAOqMm6s1q3yu7PRQ/Jfu68M7S
/0bgOEM49RyZNh2AoD4ZAFgmK1O9RkE947ifBWO011KOu8HwGF7Jw/hJmsowE+Dq
/Lk0/fMDVx23rRuMsj8l/b1qmHRi3C71IP7T5dgQNGFYd7K17Awrj2lFh6A6INFA
UJW5LPNwsVJPVpIHyoOMzEBVLVGH6x3fsNHAQMyBUXDmVNWFdPfCfzHtxKo9MIVc
E3Vo1BN9J929CKzULMhlgm5eW8V0sw6/TX2O6r+/fVB5ZQXaQZGHngnapvx52Dmy
MjxM+wW4ktGCYYxDXhz01hM2+RBk8Xy84bf8s7zCF2nCRZTVsxPD7sFI1j6h0vXR
eubv2ncX/dwl3bPGWKw9IhqBk/ty/lP5Z1IOSAEksBPOQcS1KzWY1zN2LxM0poOg
SvecUP3s2AbvQUnbeFzkVuCJzSGJxJe2WvDwe7Kc0xB/Lbg7A3i8G/82MJV3UOwS
/FKk2/Z3wpShTYe38j058huOoR5xk1SeBGHJdcHiejSr7k03paTRks6Y9NhaBxx7
miQRNACPDcnuIpctQGojvfGQZKsVmTrv1Pi1QV0EXa77mayOw6EQQ1ADR4cO8QVI
cQHuKOqY/3G1SZnUZh/OMfnWITB0TqoHeGYiAD8ZSp3MyUQUjucaW+Q2RR3ClZW0
x8sOHe9m7BdeWN6ZaPbm4PoyS5JwzPJjJT2cLIkt09W0ruttSUOMRpDbTEL1yAjR
RTwfqOAuplCF29NKLBmn0hzArSkImYK1o0tAUtnkNXjtBVA1EOI3Q2c0Nu2yRchD
HHVZeClTjdh9hzB7sTHOqGDhlVwh5gQIJ28oVX7CqrdEg/7aoiZ5EnP/VTf4ZKdF
sUB0+ATtq/SfUxMtfgjrzW/rLQ/vuvyKSvnYZkWEdh6fDd3PQdWXL0nKqUn5o8hE
DN6s3VYSAIS5M8SCwPSBQc+ChNa6VGeQ58XQu7ZMMOolIUw730DFAqzTWT1TAUA+
sD6zuKT4XJl3fnigNVxWmwryyXXKi4ZqZq9NkZ98ddzfHlwNFLCOfQ4dsnQ4AfTx
1YDITwDu6YoTTZd8GTQWHUkIFb14U73ME6lGAOi9ijn6z0DlsbOuyo8ZRm1mxRS+
686RWKvPQ+H25bj+Cuxv9F576rciBbrVbmM7PRNic47MBFuUvJelfuhWuZhb8XRh
3D4o1X2tRbOL69RIRE5yF0DaX848dlKcwjLbB8qQUtj2Ta8+Ud88i+6oprAMyjgf
gOFKQ6DAGkCCMsm2i0DXMODXjN7PDW/P33e4fzp1q9KONP9yXbcHx2PQT43CEBZP
iwZavkEVX1UcYrV/LrAEMIWEbBeh1r7WCVwkQERrfqo4D9mkcVE1ZQV9KSudQRlE
Lvx1lhra2h8yOtxWFC8TMO2h2EK8gwvkofdhnT/poyc8KPo/BIgjL9+km89eBKX7
doxSbwCggUzdK1R/+dnG7MQpGWTgnE7NJCglGlYaNhLJt7Q+WQO798CR9sQxuCIr
QbrCq6iKz/kixhW1+5POAW70fZdMmox8W+dY8bE/y+jLgiQOKvlNZ6/9+HFzGFjL
xB5enUoxCePkPMgWEEVXeihY8kBG/KVgR1kFrjnhCIEcErsEDerhbvAGftnJpSha
+Ln/A7RkwnS78v1vhxBj/dg2fdvEc4TwVOdBA2ij8ZkCn6TOyuFoNnbMduIljUov
uasAT5D4ejmGoplVkcEUeATCBZ5PqMjc2VzLoIX5qfox7HTY5UcPOCejMI0f/eFD
JgyKUPK/k1h6c7saNR/Jo9LJdzIeCt0nHxem4YpsE4WkPtQka+gvh+fIqaAqcw9j
NfjRvRKoXrrYp2Tk4RdD4iMmw7IMtbxoyuLjPV7/J8SCFqijImOXhij1iNt4QUiW
Mqsi3u7hBQp9QAPRogwcy5RBE0U6uxJgP9dXN+lyaZG5Z0x9nrp/Q96Nk0MBJduv
5iLZ2agrx0c4vLpTrQJm9MpRc9qxAY6i+6LD7tYS8J/nvay74w8cB198WljYN/bd
/Bmk9LZT6R3RYbwOFSJvEiVJYsPOGioMF4t2KnsJ/pfubVoMCMNOTBq1da+nBaqP
Y6qRkt4dPuJKSwwphYh4jZ0hPfTt6peTG8VeKx09VksgKjIf32ET/S6wBzPI+UTs
Bjqau+VDVOfzxuUVevhD7VyVZJ7aaFG5e2BT73bFfn2t7dfFT7Smkkxwde3ZhMKf
4LnsA97CXrxqgRdG4AmZdCQSdkHOSHXXAjzCOgW7mR2e0hHpUybkeVJq95oLe+01
r4B3/tKs9XLVsGFkPvtuiHz1nUwCltVCrKiFaWUJDLoQLltMaKnDuqC8jnoDbtav
SMriBGkJ9gOlyXecKEQuT8RwBdzd6tLiUsS5Ww8p6JOoHYq3OFw3enCSHCHeMDtg
SpGRr9AYvdpG46jJdL3BGEkkrJH37mCm32xIL49quob3U9kuMzzuES0evl2ULgFv
5TuQ76tmIqVKUb1e/q8XawlN3ABgLhlc55A7uLoIi/MVK0c9AR88RZFrvh058/Mv
u1uvXRZ+6aUneTookf3LHHS2LdNOw+wjMco6/2if/7Wzw5esJ4rzsxeFuDCb1wQV
RhighQ57UCXyqsAsD6LSrOwPyrR8X1FDmXff41eiv4j5DWcdLgCva8Qpa85uhmgA
BeGdGu6fx0rr+URcxHDlc65emZpvTUpgaLxW+RnAT7/WKg1ruVw95flW6Y5ZUmdd
zN5I9xPeKHQnxYwwhTUeeiB1ATrViU4DrQSdG4o5CLe0hXfHVuN9MAoAuLrKshHh
tZQH0hqyBFnUJGBCBjbUbbNxPuomaAJR2Yb1pfSO6PVWoHs7vrMt7emjCXGbsKAs
jH6/i/8B+1DSJMiYc6IOTSF5wuGnFln/OL69UGeVhHL52FRTd6EWib1Ag0E97qyy
XgSN9TipJYYN6eiHl3FDQnONcrjVKHstUSC5sbRfTEyUO0AT7Vtw0XWW55/x0NL3
ecEJX3i0F2yy9GUQ97+HPl5ogSqHF1CRM0kmWCrrXM5Uaq1Cnpjmengi0Z7MIF3Q
nPcAzHnt1egp5/VnZ/MCudYXwJx+uezXxTnrTPvUyo/BIHE209fG6NAqYyNeWohW
OVNYfILP+1fZex4CTnJ6xlHi3uSASUNflFe9j94OJSM/ATkeORlNwB6i3yWQxnyS
SbpFflYXW18VEZIix73rKR25e+FGRtmGgtKDc1wRHzM5Epy1tIPsvQ7WHxpen73F
L6DdHJs0HTHxyEJx0oOZK5sljOEZuk/NLLrrShKvfL95fCb1O++/2dUc7keoDCuT
/HyYGwPJIke/RFXQopyib8wUKOfRjQFL6HicFLc2ZoBjPyDPdq3AMDV7ASd/OpsF
GFPnWNK/Pu5wm5oVME8GEqN1iR8NZ+pIlSqXw480LNdadHdb2yLDz+FTNjnpa4FP
vQ553WpkWJcW9rzsLy9dn0Q0MUge6C87bDj47d17z46MhSowEV7PY3Re08dS3uRk
La+ZgOO/e4RsuU0X/mHHCM1MJXw0X7XUX42485M2aK++gf1K8cjSluz/nKuKOYb2
sMTv/ogOcfHyumYVNimMATvGn35k3UqfiHKvl1f42UErC+8yYslTuHju+fNF15nY
93xmG5ScSJxjLFAOgPgTlXoXiTPnHSm00ySvEGMeQzJtvcPQUedqdCAyHQjuyrlt
w7Zym9pX5V/VxZz3iK7bD30+4Ha9NYLWCz9NcygdZ8kjSFg/pGh9cwnzCXCkV6a0
nCKeIoHHraOtUDibe1s6fUj0fly/5Wns+X0/QiBNX7rjzYHp58OEN4bkmZxnOZR+
+InjDxkBOb2os1Y+j0Z/BcpLeARrNRrJ+17VZ4JCNzpDlVT3YPpp8QqeVAizIDHv
IQtVe86sgBmk49+mVgnTcyTJEgclsjnsB7SMx9apDjfY2c+1QcwbDV2+y6aJKyre
mKAlSUwjp59hPv8AWxWiaCgaPkBLhLSY3BZHDZ4bTlbJptUO2N8eazn4JOWva9Oj
tDM/st5cEX7u9f8hanJVMgZsmhmIVhoWWQITtebYUtCk7jH9yk2mRpP9jq0NOz3S
31urB/uorJspJJuzZm9hqH4uTVkMHmeuMdb2tkZpdc4bFtOjJkdiRVblDzsm2C41
HaW4HccruMgc4kYf5essPPWmbMjO9Yd1IL57lW0niu25ur89Q2TZtk2a94Pu40EU
3lGE0GrVZneSSJX5tQg5AdpoUnFZzx0G3wr9StC5Wl+erpaDsV0Onolf6iex2eoM
9nVDvPyUXxKPxwZSZaMbbIrEEsRxjqjPEuklNhThskwyKGQLsEYQllLniOUxP5N4
+AKBd5weGRpDnjsVnOr6k07a335ilMLPGx+zhrmMsFZyDZYWhGE1IbPbOR54xmEW
J7V2isKLMP+MzPzrTGDAGmA3j7bWJr9d6DJxlFih+jig0CAIGaOsp9OOKRNBf0KJ
d91c+9FB+GXCQX5uBAgjjRIBN2XHgseiNiQn2jqrnoJ8HQNzdYWQv/S4cKUt6bz+
g/OGOg4HhTKtylLu8xP1M/47Z8sUDFvJbc80O+yeFYG+nIu2O9ExHJzdAjBgpcwW
AqtmdBdbablaqEweCXmQVDhCbY8yeMtjqnrANgwJqWtZGWnWeqNMgj68aL/g8v/w
F8WNO0VNTT7JhkCop3BXUcor5vcQU2208isWcSuMEfKTy4vr1vJ+/8EjYIuBSWuH
UVKNJ+WcQoEcjA4zf4+kEatTJV4BoCLAO7yzDVOuj+wfWZYYlhND0i6KQ3QPbBPp
gKYYoMa5zCknmLMGNifhuodT4wI6sVnOz7yKbkECQiLBA7ycq7ePDA0qhR8T1Wxd
GWUFU5wdvGGZtZEUAuHZl6R77bn5KEBxmLfFBm6LOQkAoIDRUjv1OvZaLf8FcBdG
EOUT2kyX1Z0VPAP8g3GAXAQZiiMRxgcu1T9xHm/fghhXuxAt2bxcgQ5WgnA9D1g7
EmK0P4oRmK+acsZOk/ozc6DorODBZ+mAXusLWosXWLQ5UHDaSuejRg0SljLxC5T2
DHTBjxylzeeqJSC0YLv6GyvVTS9geWfhqJ8OkkaxiiSH20r83ZYawUeEWSYeRkNo
SkaOeRKswI4+JiGHtcb5jvSf/Z5rqEcgBjI6J0q1S3iJBF1zJX34apRhyAbXAz3I
K1mgpLeV7mSH3xDgzwbGx/qp7/F0Y8ujliFS4C/ZPNh/dRS6pu3C2LU+V8zP853Q
3EsD+JDaR0aYrSN3UGbj/RxBkBIbL84KAzh6kX4vWxSP7l1JK56yIPdBccb2kiYB
YvT0IR6N2UfjuHPOm8L1MU3ptDBdUBxWEIBwUqOL+NMgckhcz6ZIcoQwyCe5ROR2
QGyCgnsw92kQCPT7pEnyUgkKSrvx6sAOx9NLq0dzmpHLsGs9wtp989s79VP6cxl2
eD7/kw56b8ljAHkMI5k1VLn/lpidPH/9hNVNOpitRbZcKNowPoEIMoYxz68WCxxv
YrW5QJxHti2aVh9yeUQoY7Bq9+d0wYtzgUFgIZVSg+5ZaVnQOyEpk+BK9iRsbb2j
PvkcbPjcSdK94kyn5kOuO7PqTqohanIFnHQ5TIB1nZtjmDBnrg+m7Jx8kPDhqkSf
U40bl5Ixxk3pNg3R54Ufdv4SzVnVjlCq+0T/SGcN769O77cFJQ18sAnMe91PaZxK
M2h+2sHqhLbSHRLDtRax6kfdz9G2jiA7KtlaiiMwvlVMJbwCT/ke90VUvD0LYTQn
f5J60anoI7QvS/Xz4N3v4K/V003jJci0Ls/7L3oN8cN8P3eGD5DE7TsR3O6sOEvV
ehMv26bxAarwD0O4D8Q1U6dO4gEVdZ/cGGFV08QNvj/15UgOr4SHq/lT3c7eKI8O
4LBgymIepa8fmXDlsvZHqnasKhI7RQIaQc0fLXIOhuU7oOsFjj1/8PaF1g6ntenl
jKI4gUsXPsa4HD90X10DCl6ctBSnQ7wbC+RkGMqlu2IaL9nHRswH5BVaGFXe6Ujb
aRqV94v/w/E5xwhG3If0GPJltm2a98joSEX+ZWHsSl4nZvqh/FJgrxyy5YUttz/n
F4FZalLZBXjTIpR1keYj8B6NaecxDC5cOxBzoXwHsTjxn2XHzsbBefhhyr2tIrIz
z1SBjq9WsmFzVC6T3Ou+ZfoZlpYFKi5dn/gJKjI7sCKpwF682LVHihT9i8NVPUSv
xDRH1jVw/XhPgrbDZvbkgpK+iIKts4SuY0Wg0RJsi/iQvhcJgi8GoV7oTXNFWOfG
UtHLE0quRmkazScV7lLlzkYO7QntYYBnSuD8vcdppEe7V2ytnCF7K6zmMs6PWHAC
qn1/nOFPxheD4yQ/C4AZRcP922WJ5HBOTEac26m4wuCm2nOuy7FdxfszjDAbrz13
+wiO7BQUDwNlRnSXOOgIN0vzB1TpXrJAx8pBSV/Skoz4k3ZgmO0ki69j8nBqYZYh
QQoHJZtWo+oYWr9lQloLvIaVu7QoCXcWoiJu3okF9Vz1oTRuIyHNTuii+yhfIME1
wRzUOzqMozFeoAe71MfR/XdJpEzU+WAFpJuzYUZVd+aNr53CH0jZjHqQ0Q47jVGt
D3EYCD/grlLNmgZe8wH5vS3Zijn4KTWYqDDd0Ke7ytwr8bINuK27iWeomdNs1Uxe
yunl89YNxuyR8i9nVgCzPTmepl1mbEFsM8Spp6Q+3wiDCcffgOEEcBkvBaiioLSf
/uOb0UwmgB9xGtP4Zb44xmAcorLLJ+eWZxIhPqG03SOV4Wuddr82cZc2QT9ucot/
qCVNjosKQpiscjOtrwAbUURfB05Uybj1kqX0PfYD1UGSKiVK/YnuXn/MeTH+kYed
xbpjLMgDodq8YtS61/rrEfDjeoNfyuQhoiPLY3PljqTfn5ZznLmaBjjEBz4PLW9v
HYH73hWKF7Ue85Oz8IjbjbETAofz0wzaN1o5QtJyW8ul3jfC3Yq3K69NUBFgt/VT
TX6LQL9jTsZjGaWuYAxKB36HgC2F1Kwu1xI9g53iRGXdVZsWrZc+DdfN4TATOnPd
+rg+4r/fJNfntDOa92eN761NXujAGujQT1mB8DksaghkVxhcfFWJ50FwllIHWAtl
vVZPprJF2Vy3duT/suFSbV8C9iin/hgxdu0tzlUGCQGFWPtJBuseww8jE2pQOn+p
Ik0GIH4n2LqSPiipmaD21TJHx+zgSp/gWSUToujoH2X3AR9HG5c0BvJaMiH1mJVm
cbmmNfnOxXbNNKs7O4g1IDESXvyBpeau+QgJ54fNnpK3+rS1+ED6WCs5OH/qkU+2
1iZZUWDoq1+J5wPUCmhzyvu4GFPZoljBcYWMX6i1J1SCQ73k6xjN1YRtEJr2ZIm/
+ZraFpQ+uI3z61Z9uOQLaQULIlwzaI58sgLrC4xN7TzZE5p0PURQ2+UhgAsAT+wx
eYTnd5rQsQ+k1opBvUL+T5vE2cEiAzAYaOkgRrS740INfdeVOtmQjJutg8B0OJVm
9rzGJR90cERmLl4nblGxe1oqbxdFqCGsAmLYHp1m5j6BSMrKpORUm7X2UW7r5qGP
IB4JbadFYcQLMk8RLGpBX++BdtIs/TMHPMc42tws72c9rXvIJzsuBlzhw/Ft76tm
0OuU0sMUkEbiIDGTfS6+xGqfrHz8uVqeW461nKj7/GvQpb0hWotgzdA71CeMZKxW
FbmN5o8B7jIGC3tKaEto/DSm9IrlWm9MPXggA8zGzWdPKuMXDQmRLSWNwNrQk7lB
mXPGYuRqLuajF0e1qjNCjTaSkADxSty4zeZmG7o/7mLTzvxxa1EcSKkLnG2CONF4
S95RzKH0tZrbfuOKrI9iFBxXJM9DkZdrTfffqCwMeZv/qBSY3AnCyYPVP0YHZKWE
wj1obeqU1zlVZKaceC1iCZ02UoZ4VfWNJAw8GwIuA2OP2NzmNKo6u7AIoi/DaOvy
lE3aJJb09igIC2lTf7EpW0FnvmlHpm8hUtxXjrAw7+f2HS0KVAcvN65CMV8Qtie7
6DsbRa+pyz0LGseq0ZEiFhDLn9RZ/CafvcwmIYx7v40Y+WLr4wBbBpBmBwpsZFFv
poTAKWAFJfn6zW7nTCIzR7PTEhy2BOkuV/rw0tghclEWl7ZINp8S+goG89ynrwRO
w1vGkWhN825YnNu+R3CWlAL82jJdBOiObKX3w2S4UYwvFGr6LNi3Tyd2517NGA/N
m2OGR1YOhMva0BQgpdeU/bebTf8C1uNPqqcdoxWzyf1gwKsUWjqQZqnjh/g/uvxI
UoDdNdAsxxL+Ss2CNuxtZmc528yMOgOaKHuifqfi5jWuvxIF54XPveMzMQDT0jSK
2Z/eQABWeHIIC0W96zvjbVgWwoO5D3GY1TpQrH7GoMOVCiAzvg6RSa6yUQzJwMmY
lMNueIpJkzC9CnSwcP8+lu1gk5C+LEnt9YDdiKpZ/LN92WztVPCsSH4/bq+GLupn
FDsMbr6dgBeMppAi698tbuuS2K032WiOr4Ak1SrPPS/sLMw1QfVqQV1GuC6xPy35
fO1NF22a0/OZEYBMtJCt/prphYxgWnoRPpPwkCK+MZnMvVX4/bKopSVtl4+WXjT8
0cjwwq8ra2JTNfk3sucUX3LtObB1rfhumq7aLOJvEQKvrp7MZxYy6EukrcPSnF5n
Un/hszRPqQzQ0MeSEf0dXv6IFoQwqT20zojbmxZy4ODaeTCOpQ90XPN2jvpfH/Eq
S4igDnlFJCg9xhgGAsgB7E95UUXoO/oBqqFEwd+Yj0J0zRBpnHvALrEaAIblKgdY
KUJYIG+pFVgO6uXTTOv71yHlAVih0T1pHQamch9VdKIvTkxQRZ7r6bTYOTTh2g4n
HHAcRMh++yLfhH5NVU3ampHV1ATo2A8RGDR34YEPK4q8+kVjVMfv9Wh+/Ma719Jb
XMUxj9k2BEjMKubJL9TQFli+mk/yxpwG8wix4ViZ6EcmEUMZmwfVqxWqDZrWdO5k
8yaTt5DDtLFPtS1xnADqaPl4VVG6EFD1OgbMrLj+I+RkaFLXgOf2Q3htIPiF+qha
VC3fQ2zlQROWjNPXP2QlIQNHb4kByyb9k7SOnztAyM07hG98QFXdYYHFKaNDg8U4
XleESfPfuwYzMtz/KZS9/NfGaCkeftrTILi2jtqmc9GI8jlghapiI2POdox/+Mu4
rllJeZPNR/Qz6DrAHEyOQhXbFsb3Fnqh9rUcRJqqZz7nN3dZo5Vj75AXEcbRURUX
lpaQ3hI3ziFinVEgV9ingg4w0e5kqE/h+3QG/aFS8ObmLKx4+0R7i6RZHzvxFEpg
fQqha6igc5iiJQQY2GDgsi/bdJG/jazd+qhY7v/UzPtI1E3h4VFERCNejfVrD2n/
UGcSrkPClNG0hAZ2XGP8J/qgdnovIUZ7bx1FvSm20MVuUrbly5W/y1OE9t7LKXUX
kU/i5nKoS6L/gvJmA9dFplXBbSafgSY+jTQLls3wWrFXCgBB9XNyNX5zbpdegeWG
JwOAX5e61Gvo2j8GXHW2RbKj+Tn8ehSmnJuXczF4GnGB+sWOHwp94TeVdwWmWkJG
8W9JXo6oZ/SiBs84fRy+ln8cvzACYdsx8bf103vWVMSbDJEzXRFhenNf4npT/nU6
4yYGFuS1TRfBKzyZJRgcVovCrKidbnCfKtY20DO6lOHewFs/oPfBoKYw4bI6sB4n
/yTrh1MxJRmTRdusX4Ij9H+KJkVo2J66GOjmPkiIcYFtaYp23IwVixvD/O9wftDG
JTIScxKy0DwjFkJiHsKRx8Z+7h6wWwPzhNGKbdin6sbXXIAiiqY0J/btp89qJwY1
8GN1GbktQt9SyZm+Pc7K+65aHbCgomrLRUwHbvJ8xqdVJ2ER9nj1c78BkcQkEmwI
vltxYDTbMkFAsFXT5/0m5qjGc4SB5BzihXmXZAW6HFGLOJILQhbZzzCteV0xYkzi
Cyq6qeqMTZ0QLm2wME0oTYRB9xF3r2iW/z2E/lDiY9U+okzNdtaOh54Q551Q/7iN
hE4aFPOHlld0aKWucakVHSU5dU5B5D3Y8MPU098sG9unlp41hvRCm2xaEzUwuliH
Z57czYOJUDhfSYnqvTVxNChrPoBu9T8e8dPpar6pCccjkWlqiaO6xMgT4eD2VlOd
T+YBV6yOaZNj1p5rBsRhrkj1Fkql5BJNiZofZ1jWpfz22K7Ekrtrh589n6pPN40q
ynmAXVYxEj059PNTKncw1FNMW2E69s6YXmsJTmCI0AhUJCU5WhXnX/kvaYrmHmUO
6QhrMuISlci2zLG9slKM4LaX5bMv0F4pLWBlzOo76/YmSMNyhBggfR+BC0KT/IP+
jNaMl5/86mODXNIiFLDnK9jdm1p8fLD3HsZygIblteadKCLyfuUchqYLz7Ohiuqo
JPahzqIQmjCfXW9S98hN3AS4XyV1oWX66/6um2WkBsX5bGzbw0pTZ0DMbKlopsty
xbkAD0+ryrALne/kDdjVqkvoMwTbWkEA1dQB3JKkVJY/j3dZPHQYN2nA2cW7jQvY
8AhU204Z4LvZkx2oMQYdZkHRI9hMU4dJCaYMoXbTQ6B8F8YkvvJwMPiGwZsgPRtS
RDgZBke+4HSd4tdAMmJLKYLMZYIJuXeHV/ChvoaVbAqTOPvSCqtpTqeZ/u5Oyry8
i6k8kIiMkjZisaXe3kBpQtdwggk7kZhfOtV/aryQ9OYNvMkBSnpw4LSgqRLmB6xu
8mrMhQefyn6nknbhHWvwrAimN4Mk0Lb/8PQ8nBFAxPDUvDn0tYaAEcx9WkNqFJZX
cr+TjWB7CC+SQxiCARQSkXkJx+bzj/6tpvBUiyWvwDNucdQ7MOU5J7EL46T+4zI3
W4bdXVfOlguKTd5FEeB44hhXd25LW/RI2FvDeGATmvHPTTYUPkgMv1Esk95pUtGE
6NMkWvDI5fcIQWaaNwUEdOHZPabVu08spxcliNwcgmn/lgkGwYApIZXNxis7vPb+
wTmkDPuN+GNsXhvG7XdMdysfBruzaQlRdT/enab8lYSxM1FKFMKNGKPyaMbPiIa4
jMzn8wqVfXbtFsEo5HYovP+BOWp6ICpm4pwU6ZNyQ87dP7b4cZpVP7CIzcPGTUTN
sWNo6FrTV76DOztHUvDFiLixTfxdRlnojlvmr02egePhrzkwqd+5MRZt+k77hG0E
ED8g/P/wBLjqsX7DQoVBd0gFhERzjTbBbFwD8fUjNHzbqB4/8kcMmLocmC9NqVJZ
dupHaxQ3rRoJszDhq74gGm3GOqZ+Is25cjj6vzD3qUnwqRDcVlvOp8wnRPVu4TpI
/2eRWTS7joQYemLC+LJkelAYytcwAuJAc3A6CgXkdFPc8HsoW/7tkx6Vl8deOJoh
zCjRa/v0w53DONcmqWmTmYt4v8n0AwGk9xN758/RTQ/n2s+R0JQdBSemoi8sLKGn
BnMO4LrXf9rIrTP3fAoSgJXoC9H/K09fAKEY1jyTdKMVrp5E414/byh/4TmI0bdE
6frdUkgGK2jpYX2iIPdp7MwcYeyITvLXNCwXRKC8/hsS5tHeHourhnR2nhlMJ1S2
OIBqV2A29oPK+walNzP0ej7WGKGlKbzACgrAtqBX5hOv2NkIe7Ep3/TGtNDVe1je
cCkAnhRkPKsVQYewcwkHRepBYJlUrG15Fgy10arE7HI3K4vvUTflrlfP+JU/O/Y9
P0sI1EkPsgcDjSgEa5fqoDr7Gd4NA/MVEcN2QrzL3Wypc1EglqrPIa3OAEp88+/C
Skjw8tpe9/D8YrXaH57RA2QWR0fU569SEyqiwePhufRADukNyObw9gGfsyLJRLSd
8LW0AUq54uFRDCgpzNlxXI9nFwDCdtNPIfaKfZjNXLXQvmvVdCWMql+3Idvmztkf
RGmdLdEAywugIwaktGOZDAKCCk8h1oqADTCMeDcHE8n3JsosubNx0L670/CZ5akH
m5vTIyz+5J5YivSh/nu0IwLGVNNmNl8RTlqlBeymQk2+/l1bzQsSQY0/Zf2fHY7i
8ZLOB+yG+sbvrtpVtcMUhrJTOERvH2v1ZOGy84T0MK0TY0rw326VwPLokYYsV6Ig
8s8MKKlo1RvzHzLOJXxDwf7T9x9h4H+VCPCypbbEiEnZTGXTZH650TsSxf4YCW6l
1RTLRWRK95LHMy1QVpiGsVYokChnO2F7S7rWzzFUDLCwNka+SVPk53pmjFlwPyd7
iBvRfu3MWkVuJ9dJVGtWcwmKqC1eJKPHw/lICAZACH/NM+8jjZuLde+bxplaUBfm
n2UxHpQ6HX8MQ9JaRnQxcnAsEJXkbvvYnafQnHXWCdJYvI4GcgEC9x5JoijIsHWG
qauuA2DG96F2H7xwipEtKh8/25k4mQ+Tj+nCjAralEC9lD4Y0+fsGn55FGXa5ewT
ZFoCMLTh2H00kZGHrOErtyocH6XiroDViHTq//RAFbBiB/eTBF+YFFJ6z8C3JzPm
SNFlEu98L6swiF+7kUjvlrXWwUZyVN+wAr0SINzsCACbjYFPcdDC4efY1eo3KI+z
M/olYoOHur82gQxQMmORUIYMvTJIExZQhiGLVwZbr76Fn1k5O7jT6CSUIXlp/C6v
76ZBYZPVw5+Wpp2RkW9MryP3ZvWqqKZo2/AdP0QYVB4DeNIUD9eYg37/0gMN4SoF
cl8sjoRJjLxGpiwGCLNfMxjDLqjFaGUAZ3kVm/s1CIgVyepiqyOCRTfNXxIn8KVl
qHvlgMTx8DQCeU/gkRZeYX3nl+PzFHyMYjLKK9a7nu/bB9A6vUlEXgJb/VjAQD43
ivT2QGUfxSDA4v0yxnLFdnzEpHJyIN/B6F7P4ulnYKR5PULkwke7En8OOdk9PEuy
G+5OJbHvJPBuzw6mp0kFKu1dXvBwGp+gvhdD2TnHGMMpj5Ynq6eGxtvK605/uIfc
MryMf8U0rq3lkytFetkmCOfyF3wOihtC/dC+xIlzcgvYC5pNE3x0LsqgshDRluhm
FXJdV3Y5PhoP3dZNHPBim7YDS4RM79LnSaU7ChgMvrm84VxUeVVxLWRsQWnF3i1b
HQ3pvXbs8UI9hjxaf5p1P2+q7JJn2JIr/ZnfEgJ6dwJKLUMuaEc9xUXkQ9NEtTOK
QhApqesvBF9ToJR2KPiOAjlSnXBl4TmNQ1AN6qu5N4qzW+mzR6RjJ/e1RIwM+Onm
qQH7KaGGAK58eePv8Rmdkp9H2H8a7eIQnV5g81LvA+sLYqMWEsg2a9icyin2vafE
7cMjrX3sPeI6nuvG2bdNVaeFTpR3gFgl1UXTGhBJMwB/WOol49DDVogpPl8tAtjg
5I0l/2FnoiizImB5iGSqKI80rXY2R9VKGF4/xHl5yVtXIxE5XKX9k+sne2mRl1kA
XKc8wVehBfwdCxA8fVrPRJnLcMn3d8DWLMdsyFQpg+22QjfizxoWHAz65u79iyOj
BYr53lKO7IE47I44pSFG5TkK3HukvTfsb6UTD8P9A5AHwZvD9uH13/sMrTlzVONy
CrOrBNk2gC1eacHGGkGQdpk2FLmIBhhb5DFSKKrly9wn524nfrDQCzBqw+93Huob
9TRxI0nTifRcONf3lRg8l5cNxtkhaF5DEeoi1tXe8tt8n+OFDkTvZ8H+1eNgRqFB
z77RuOMzlem0+7KjDWbRHyQ86JOFI4gb8q9zg71vwMAaVDt3/nExBpA10FAB0cOc
ay/sVUlik5crkNKN9pJmkShVeassiTgSCf4kId/LfTKvnw+ips7xqc4Z9UoMwLPM
h835CMSxhQi7vYR+gfvBOAR/aIu+7C60FkZT33QwqlpoZ8oGs4hT8sgkIq7IFfU+
zINUioTZ5v0Woj+oeztrTx/JL8rpLm9+7/MqbCIKv+ktPHmcbnm/Eq7RO1Asq5Gy
LUR2gjC1uLyo02GWiiiOHXwx/cMI/pAVywD5VtuZocrXYac4UfcNuJzEgVo6ODkq
R0o/RebouIeIucHgYmEBj2IfvskufUMvd2OWYO4w9L7E63NsH7CXVIyx5xeanrzM
zS5kx2zlGrYonW7Hu1EY2oLpnus+6gfRroGv5a6+CI6E7XrVE8A76FQx0C960Kw6
i1gXFGrFAEJf0UXZGHG0+htHLuosqt8ANcxYUnHvmV9mGVyhK3YQNr781/PGwOMO
NaKRU+328Psm0H45xH0WIxyQ56f5Pmn8UxqrzFNVa/evToj08ONGGsQpkBIeDTp/
mYzhmcbVoSpNAUdHJb0B5wOqnzWMOCHlRpatpRwt95ux7ZEfm1YmnyqXV0RR0c5Z
FoXAhwpkrFWGbmP6rGoe88LyBh4TpoSHABGv8aQzGetFST8cjaNTea/phuPZEXa4
Qd83vzSf1GfdIW29MlGxX8zqO6UP8kZhR8y/Gkcgo/7m+Sp6Xt5FkDdKUk1tfmLk
QfDLoeDHGTz5bNtw9IBBOnjeYYEmCuvZJ6NWM6asqJ5wIEuAGoh0aiNP05rYd5hy
PUp1ZI7SoTYArxbibgLmiSPOX0iicT6bHS55mdtMhp8b8QkgnuPeVurAUN6iZNIS
5cdkXWMlBYNkyGZAU4EeFfdnp9WkqZH0rUcjF9mOBnWIdKlsfMTsVGqHfRwhiJ7B
C702oaZ0yImg5GCfWzq+6EXb67mxaPyhVvhkaUXFHh6XyonHZNczk1kKSl91kqtt
kLV5R9+AQ2HJdPafAABOPiOjM7YQq9BYhRXJIbnsLXcBh/hZ0iUedIFWH6kqHN6n
RrMXD6XEohKqOZOlkvuJsBFayLlNHkcPwekAqjJMRDrtHWzTuhfudca9UWqlF1P1
IOg95qnZRELGzgMJo6sf4/VBuMhgpDmkFIVlve1oPYKMzCiI2AiGc9Y7BDEjoLUR
/QaDXdv+sJxvCvRURfs54xxkO37U9Mo9QMwl0mGI2jBBvLVf4NhrLAJ6MRb5Oe8g
WsANKMDfsteM3AjvCTcGn7bHZW1qSiSVDOgcYv1SFDFBlLONrJuugXb55iE4/B5Z
4nHW3QSnJV8wSL+X/OT8gbOcypXzu+coIllnm36W2b1hB6KtTBh0Jz7WOhZ64XgG
b3viYdhUiKhBNn3fkc/JDQTbXArFgc4T2Jevl2tDoDuIn/Zoa6836DOx90MdRjw2
M37h0kQpY67+JTUnzI+i+i7Gghu4Gpw2IdGos4+fQTxdFRzY685v8by+V00aR16M
EWB3qwQmrEwdifqj8xUSXpOCaMcwMNr1LWAKIrcK82GxMrFIL2TLpbTWG/5bJi1g
UwPMN6gImtpcnvDsq7xD2BGKIg9Pct4uNaAgG6rNMfnZ/z7yqbNLlHNuLCfv14or
84qqdrIr98TYVbXfE3x3uqlMIcTtbxpZSQHa/d0gKoo5nn+qlA9u/vZOYd9HD5iQ
M7OChTw4wQm9iA6V9bQ6+k10kztEilLmxaqdpwKclp2dBn3C0SxAgiq6+KM9MNaf
4C4ZjyX+SPWamqcJ1BkrFjLwDz9M1BslV8nka29pJUsl5Je3pCerDMPC5l9Ew8J+
pKnWCzV64iLQr0G28liIh9bW1181X4G1dMkaqWbcUVBC2TYdTfErPHRsLnWtKiO8
VvgUz3s4611tft487GX7iEECV/6oi314zWH55bARnDXrRU3KJ3cwrEcHM5mGu1VD
X66ERvivtzkrSvcL4SYLXgD6riXDNnZZ3M6mhOQis9UVqsjsT6JsNQ+w9j9WUZqG
smvjLKWKA5A+m+7EG9AFQ0fRn3YqCpHmT19VVQrg/I8aFnPReER1MXHYeVhaR2/c
/+jXb2Qus6ayDS3+XKfG2lWsxRl5wjyrGs7Q7hFPOIxKn3KfdwwLAM1fwkNeI6Pj
Q2JY/WWQ1GJW34ijYdOawJf6AahhIIXtuWInh1usJo05ECA6M/iGQcvo8Tp+Z77g
9YthlJxg6A0dH8Qhqs/x8EDVyCOZlZHEBJGGtD4F8O1fNTScV/ukko9cruJJeNES
OydGvgtjkIZjzhUnHKKwXJ8H6uwUSFr3H9ljneqvq7VgJvizQtxOSVGmzDS7AqK0
OTn4l+/tmwVvEkkCM7stemhBVJZQOf9RPLig3LpUT2eawFeHZiDWa+38BWDjbBlv
iqgL4/jJ8WbWOV9e4+KuH7M/+xM7OzgvBcdDkRx4sR8cwisiHkCBPBFPRXgPI6Mg
LbmoGplzjp7GQOgn8Oq0kQ6MWrL9NQPfDdDD3lh8pa//BkBPjouJTwUpVCDlAMHo
Ku/ZjFuk2t/afpovOKFpatMtkG96uFYh7DOuXZlpRAA5i+jkBugP/7UI8qRhQye4
xN2/t0A5SUZf8jtDlfP1fVj+t+yapi10eOeldJjf56PNhiq1aB2T+soHWe3DcLWk
7Wl3dJbBLxi4Z/HgUb7uizZ9wUE6NqW5AyQgVu24ixXVvvd48Ccez1hUx9pojBOD
wM1q8qMCzoJM/tkxN1LP4eWagRkRlLvHhadojGRB+gW4vNzrQaVoLbKz3pwnwAZ2
ZfrO4dkMcE8tDs8lE64JodKAyA0derc/egAhQuMu+mYHDOcJ+HYR9AnBHvBQGZUu
O83KJVVLCVu0026f/SBKX2Jc/k53qxhJZzLjy51l7gli8OW15+xWgi/w+7VbES/U
m6pXuX1+lHIldxRdGV54OrTs0yj0XJSx7ufAAhUlSUnuONkadKuGdLGHxQFkxcar
R7tDzvRampTG4ESLlLC182OeZFYTuBA99McDV07GR781rPVefKkPJ+sFHzdl3nvs
+c4DAYUaKaH16p5iqEhK5do6NFbmwHghehGaz0/4fJVhSh7ImH+5T/KJZletn9zK
x7vOlE9A5Z2sgz6b74H3fjXnTJ7/0fGn9Qc5Dy9jQsHqjKI7K8gDk/zWHY6rSxo/
6l3xKbmOUbkzvXlPHr1xaSrtCfL8B0ohs/Yw6pzb/pspErHwi6fcxdQpmO+mH9lJ
E479ZsRo2cSgO5TdQcc3WUAaU2lFB3wJ4G1KYC++ynjD4tapuVota2tppqTieCEA
bGv+RWeQpk7VjgJVSypqu6yX5MJ6iCPw0tM85cffXvdVwQKsEGQklbRo3WVSxbHB
e9DSlbRfgUM1mCaylu+icDolLxN7ODlN3MXb2Rx/NWbYthFm+XiAbFMwxlK1V9bX
7NRapogobzID3YkNTD4H7uRTiqXHhYLDoTFPDvlGZBTOLr4FpOdP/u/ecylt+dNC
pLuVQVNHwHzYBVtQW/BIEx+zCyNiwDchi2321CXWN8lAunmPEqVWzBjGfhCePMoE
o/q9/hHfCEd9rIM/BZBSLDof6/onUEZi/P/Ih/EKKbpB+WZdAkEPMOwFieUMjkEl
GtoVVfiUisiunMUL+P1ZSFQwk2Oq/Wz8M+8XFYc3H7Yg+vJaw8PIomy478TYPH/m
9A/2LEPFbyV5RXGltHhIIKDUNi9TWbp6y7MH0mR/GjuKVQwuZKMfWxyLa6BR5Fnl
7ExoGXawKKY9QDujuMav/jA+jf/Uy4+Zpbd8VCrmGNLrNi7oTFXZK3V18/Mj9tO0
yWuMxEP74erZC7y/NP9/Mq9Ek3TTMEfQ1qr4/LoCOrLx5oVumu2oWBWnGju/j8qy
gQ1LxUM1WysuqCM0YCWLZVJKq3+ReSL5N/4Zf6iPsfh5Jtx74lT7+dGrcwhjgX2Q
LvXqjGTk7le/mXFhFjACnoOVqUsOEFnhgr4UKVxBhXqAl56pLogXtxxx5Lp6uuZf
wfQRmaLJNW0VPKQcdD5nIvCzpehRmwGxXAX8ejGTm8shMFRAzWnHW4S7ZTzhq4vs
nX6TLAWy61Gh2a3xBdvtUamozWz4Av9f4Vh+ATERPAsgSwD6kcNjDZqd9HfuZUg/
hsbMWmxmXQilAR5mBrtHRxqa/DVkYEr+Oa+gozRvgB5DWL+WYkeKQ1ZCRZm5stLf
ouC733nRPoFI7U17T/vLGUlLLAeS5WlNmpOXHfzRsfrfmRH2uuyKjM+JA2o2SW6m
CkYnKZHvpWgOUANlHNWdQcDfz+gfrIC5IvYqOUVdBPN1/LeeITfTMAsJff/ILjzJ
A8n/GqIVo0qeI3iccylOJlIefqwFo/GWV6d6y0WG1YvBIj5BLdkpOfokU+TS0yPV
dp4FJtjxTkScsdMtxdrYpTnDyLamA7hUds08uc+4puACFY4nJrfAjiCmwp7f8IuA
d1QMB022Av7iRsWOA/+Cn7D624EWwl5x64uUZxXO0qLPSGJ7qyWLnXDl8P5o3L0w
2tYao7yic8OpF5FoVSpjxWMU1JnFB+qQaUnbj8b/3rnY0Znb14pXrkPBoZgt5hed
mlzP1lhqAaYU5co5OgDi6w6DKVkJu8u+vla/CvCuKkzh4uguOVzi1E5cAgkGFYdI
T/sLKRDO2mFQzyzgSZVH5lRQWWJpgLZkEpDflcI5BjUEGA/fCbPBa2HMrNVYQMJq
VJrsNmT2T5sNd0/Lfp2tIoNF94sMM1wPWXhEd2qNrXJarIH0psZoOsEhD/jjm/xi
v7Kr7svzNarYMizuv7YJC1JHWV8jrIq56+7rmHjMA1ihPhmlhXXgcAodKjL1BpOb
kP7/RxT0zQ2J9oySAnhL/gRpY7tIi2fjUUPfVLc1tmlK7PaHDJY88+S3BTyRF+aL
5QciWxTgODFYzAb1jxIH8BCQOACGsOKnWWmKcMkFeNK8lIwv31uyTH4hyLBftoXv
NinTDL1xt/V/Bh+VlO9XP6W2GjysNSnzmekqxxiTG6Rx0lUNiq8Gllp0dxA4upjR
J7O6HsSy/HaZZJPxKy592wxjQxaCPsrEyA2wNkvHjz6YbWc/lIarKF8VJYLRs/YV
nJeUXQ3biBNvrvxfa2FaLQS1rxQbKdIQR8bWS2KLJY55ChM6YY00Og+lV3uae2SQ
jSLhBIVJfqJmMtOBi0NGR8FGORz9KRJs4ZetjaMTOuVYvaYuVKYLyZMQM9lLe//4
On4kFt8BMCUU2P2cEYPNzWc2J5xCK7DWCOcG4VKK++G7K+f4woAP92g4XAEMeJMk
jy24SfzvcXTNPrHdVEgpQe30Ybdta2Zh3thECnFpFngC16RneSmigQpkzN+609X2
5yD2/MqpkEyoZbCnBg6/ZJXw4wcYDADFa8MyziiSkNN6givsZcwqYehkWg54w/WB
80b6sXmsn0OH5sK1aVFrxrVAlqv6xwZL/v20bFOMQP8E1Cg8AQUdrWahdDtPGF9u
UqoTtHMYCL3B2psMUTRqFTqGSnKFTdiFFllqFFsBMkWANl1EJALjCXFd6phBlX6n
fosgewOF+qISxwORiCGCGbggIc0963+NQMZGitpVM/YWitF5hoXPZ2K88N26WhhL
o0D9d8/YntNXdltDfC383W15Kcu4wrH7q6a4COUdEndaQv+GBV/xaQ1LUiwgdty8
O51gMH9xKXB5rggiKpgHuNR1ys7yQNJRfkVV14y2ofU2U8JObw+75ROWie3oRwZm
qE+zrqjgRTQEPAKurgCuWzIHsDvXr2tJTfw5aK6lXTcht3jDAseJiSqQTRpG5O4G
H98TWfRZ7FCKDJV7uFHN+JP0zXUhywX0Nlr/A9fI+lEJ5KEh2s6VltJGuqL0Agmm
VkQRCVxz9m0kmS3p0q+9LbO2KS/Du8TW0go7kX9CC2Jy2HKbQROiaUt8w8GJ9vUb
a5Vy/5iZuDjbG26/jEGHhwWOVauSBcOJapKJvHNiOshXC0tLSFttDRqww2cT5YL8
FYLI+uCT4rOfUbJ7sBW0j4PrYaQ45DWqzsgdgqC93hDbUq42RQ1GF2RyC9+x0lZI
s48mEKaeMGgLy4TpemV5WOKK99z+MB2Wy3TgbfHMFWG4Wy8C/QSAzRhuEP8WKmeu
WqsFqsq8O+A0z7JtDnvoPplqeoxGN+Spn3uV7kYoPQ/Ij2cXRgL3mlr9hAMXQSkl
EX6KUl5MDv+kiGvYF02N34SarZxOKv+wCmypoam3aIgYFbuRyabcDOCbZYYGId8l
EqsrhZekvtwyZeny3UcVmpqcNkiBnjcmVC6wdsR0lclTTxdhD3hPizXp1gqW8+HM
ST7RQpvLe7x4Tm930HP7anqOSwG+dd5817n3v+cJclKTFDwesiccIRt50wSVHCqU
4U1KAcrGvxqgfsXj4ypw7fZcoAYlqBWtxV52qSx2bQazJ+zDoa6t/w+1pd1JiiFP
Erhh7io8zfd6RaHkkFXCCXwX2/qKfike9/TvXnyrw0E+5tdhbHAwKudJKM2xj20P
JnPV2+ymTHuWYZWdbUgtQLlsJIqDj4+6XnLGKqoo2rPSzXIM4XB0AVLw6Yl8XRsl
o+UEA6qH237iQcVsDdNZN69N+auBV5D3anI3/+KfqzlIVRpL5kI4Kcc6HytI6dDh
WOtSuC0Fq42hhUAK/epaUFrBeVp22Heq2khF/IqWCpI8mjLT69tZ3L9C+vhnQtLp
zXM/yVvksTwfwJ+Py3C78AhIqLh/kYi620ZMQYqbSR6UuW3wcpjbxMAduTR2edB7
Y/YYyZXNDGDX/kT5gVKcD1ZAoNX6YVBg/u7uMxwfWZv+w5Elb3LlYgixSViwfPjp
uOK8LOaoO5+qHaUUvcaLCSVhSOkBYEbqw8LFh43NfilkyWQh0hDjSOdf0pOYKAcC
xSb1zePkeDhJQR2/VoeN+B8ZfVoWSTvV92PZqwC4tz8T+weOTbuJSQpNubDIJTUZ
qtVBOXjdVRaEMWmO4XFOgI0ZT73BPvmOJLUapN3+yLWBlEeemLIEMEVzxhBr5Rt1
cAmLkhG1RzLXtiJMD1jRYjYr60hwDg1VlovznlCQGPTRyoR5scBBLqdERGXSmk4L
evpwls5sdRj+dGFoRJQPH2QY4zZ4xsWdBkXLTIhoqIubeSBrSAWly3kAHgy31Wc4
qMH5hnM9yEd6c6kJ/kD2oPdVQ2QgIhd7Yq2mDMvmnwRVMLzgeAP9mmkvxVL0XKgu
2PtceLu3Uv7YnNktQsmBmoCFR5b1QjshEPTXqUU16NwBaSOxKp5GhuF2WVZR8A+W
WWEwHqvKI86/y4UkefnjdazfnrYApGOi3QZSh+7X5WmIxw/DYbOMv2C3DV7zlHWX
dbsywfG9pi/3FiKdIxc+kl+c0/irSRPbJRvWG6/7WHzFMLVY2c5V29wjtJCNKWCt
Y0JtHopIxljcdU63H30Z+aaQ8UoGf9aVsh9zsgXM9CvoMilhaaWaTiaifxW/R5QB
RMrSdf0JrXD+PabqdsBvLkJYwdxHNyUVp5ukXQIXASu/UU0yTgD58E+t9e7gdPQc
OShIvDGn5ZAIYBs9ntNLMhncP5CMeRMWbxR3nol/KlBrUnZkt/xyHZOEH55zTR4l
hhRoTzR0jH/vixugDP7hX++4d6mMygteonbrsH30CUOL7V7ZadXTuEACZJk1Elk8
B/l8X+sfqd3GIl0GjGpRabXka57WtvDB2kYqV4Do8f0Z/hLbxa3Up3pEG30atdVF
+ioLAHjpb7W0j3bMYwgsdRcE5yUuxYnGvYUM53mNSohjFmIlUiQegkjNYPrqjrt0
DHzjngdpnhjv6hXUcH5fwyt7w8KfrSmpq8j4fXYdkpDJQWLMVt+IS+sFwL6YZ757
25y+vbTFZu+OzYNaJk5XY5xwxAuLpCpDDDWj1vYwH/ZUb0EIeXVr9r3eT99f5nte
bfmYe/SZpYInRIUQPAaP2RqRWWhLBRpJBCnkkT+g5EAW7xqEebOhW8sYBtrW8yHf
Rdsc9rk+VqGrj+muQvhz+oN82tgDybXVCV7SZzIOWhUuiXXTc9/3bYqzPcDfuEo+
zpnCE52kaidOoxf/J7h6D0OGtSqf1bVULW3XihUoui5uMTTHa0qURzP2AapSVWPf
S1uh9ovtxehHg8GhmZAtEg/UPMHGpogBcWkYCz7lFKF5UiPjzpHLAB+AlkmR6IHF
A2z8DjDcF+pSyx4xJcA5dMV/dFib+BCdxuLonUt1lW5DkYXOWAuhooRvatj+rnBq
LkxMp4w21xWnHTp2u4q9PG9K8xKmDHHxyk3bSbufJZUl6qovcSk8eZSy1Qt0I7DI
KKrP+VxwY5Fd2HhzjTaqOCvtJjX+RzoRQyXHqcr02wVttMGZ5RNiS06mZwWylXY4
DwNfP18V6i0irHuhvVSG19ZGEHWLr6Fwg3qbgGTbse1QzihDY/1BMCvjNrl2VEAh
3XqM2437YBmkIvtdndjUZHHbT7CNxF7yeO5s5/xZkowJrkKDwdJ4tQs+dXHt4fks
7sbk+Oj81rnOh7GO8s46HB8msZB8t54aoGj0aKTH+woFItijM4ZRT7ONsjggEUjq
VhGdxZS4Fa9spFvyVCWKlXZbh4fOKoIcBuVeNOkY/QdA20mFn3NQsPXJ3mYymzq+
BGIP0xwmLNUtCjLKebuqKghV8JEJnPyzq8rhMLzyEwYeKR4NoSeftSIy8xp8JeHX
g/g7Q/xfPq2PZ31g31dHslPBR45r5b2Q6aVavWEuPsM5s+9u0lDQSLB2Ejkh3VvN
3qA0uv8Nd7NLGViNKCTjcUrLQVl1am6/Vl70US5jH7vspS+7hLBdFz4iQurSaGcJ
aBCi/0/BW2tG71aHm5ua1oUWlApW9GpYIOKnLzwcIyY9yxvq83Me+BxOtSUSDIem
0xb7FvP+/WpIqIpzPuUdWevu80WDjmj1LnxTQjXGDFr6y2HVlmTbCliCldwcwJz5
+IU1R9ks26Ggu6Pk/xaxCH7/igWyw5PhdBV7dELI29/4ar4pdL1ZjJ943uvsvF1e
spPDTeRj8k1YuJAB0TyiKguAQ4fJOOCuTkjSiPm7J6AxBYGRYC57Ns6AKc3sFnPT
w/hNTZbG5cFuloVcILbALv6nFx2NFQTm+YzxeO9QeEMNmvnvkP+giatm1lh3yCPs
uENmlE0AFrOA2jnVpkSD0HRg+e8FeeNacKVEK6+txpMJ2vYIbHd5XYvSir0SOjda
SJK7pnP7oEX7GNmc8BMhArrZgBQ9Ve3Dm/p5V3ZK4s0l32CHaeuFItfxwP7Qz8RM
y406eSif5g1mHxWQ4IjI2k/qLwXIM1BMEEwXAPCEA4iEaxD2m/J8kRcX2qzqyxgT
s5XRyjmmtrPinlZX3UtPkGvKvIrTdLilcGHP2ugLRxjmHkmHHG5WtKRr49L8ihsz
aZlW/mdRN8HOBHG61r9S8KzvKOHWIO7dS3h5/DcJBV9waHGYzTnEFccxHIUzLPmK
Fs4lq9MWXKTNIjkAZR+mlPqUXcpiMZAV5TX5/ZZqT/XT3Yj50cKeXvrVgCA/WjqK
JlLLca8BTrmAqhumW0LGLAKwsaxxwvjI3gbhefwfox05LefDxg08dc8k/U6GO44/
uek+1IvHclKR8399kbJdudJ/2aSIwT3+Z0uwIkaSaNO3/q31jyvF/AeQmkIOLPs5
L+g9w7qxJNqvtJ6Xp2i32mfpEVNZHucJnSFgEiNDgBLjvsYNvPtHGk+hbCT7DIn9
xQYbuC+XgKbh/a3HvY3qe8TxU3FWR8Q8IU5Eeg1R/UapIopWnSLySe0C8CYEntow
bBEc3HaDFHkvlIvq1VcgJPxqfo3li8fbeSIoEKBWhxfyBiwip3jQpXLYs5aQ5UNP
Y0hm43+gz8zLjyvcUCGNO8e6T42gaSnylorFT3s+N/m55ibcQ0MjE0NcG1qIWxv/
NVVczy6geOJcFebBO6dR5OEqIIeiNHOLYIFprgC1F6JXms1tTIQPnfo0acjDiz6g
1/j2e73pCV4ynIvHj/KywNpUEh0bak6PR6cHRRjAH+OtQmXF8PT0qHfXm8R5HkLv
C85QoDRE4rL3gpOEnPGuw1V+a5yZoQTmOHXyiZ17JveBuR2ZHHmp8aofExYAeLHn
5v7qSJ61a35mowvfWR8ZJr96CS08+pvNvkP7JuGucX5lBMqmF9bjf1MR6T0bjdeO
988ikUYIlLzhVPl7z6eZo19J3bFAuDBidmNbuFIWx6kBUz/ZnidJFIsNqKNujV9U
y5TB4B5FBy1DWSO8lIG8mMt7VWKnnU/nyX2jUcB+2dOy5ivdpPgCdEdNYDv2tkbp
vK/2KW0RIFGK6umgisBXqjkALYkzHF4TcBn0m+7WogYWmUnVnemkwLJNLxY/7GQY
O0kI1jC6rg7Hx8/BB/zKrYPWRVgjCUZ/duiWsQbgXEQxDHCtKnqV1uMVqq0Ux33Q
oPPjMUnVeMiWrtyTQwKEpjVjK1lcu2A0knblOKAj7nE5pUstrsU2Df3n4FD6X6pe
H+kwrvPqVJgIv0dqVtzrlwL5ggNw6sUu3fplLOD6VEhd7eG5WN8TpGl1qJqjK8gr
F8+0TnDkTlEW49CHWSFPSw2H+BZZzaO9IoD3ubMhoYTeXtYVcwDmBGig3jspy0ui
h45bzTRdfd94ACAyvD83xmAM/abEapH2+uC8+aJkvqGGNzhhRoJrvXHUtUBP3mq6
UAeZchP/VY6RTCpUL/fHZQS+fiiy2zqE8ZCW8FvW5JLdxcy39t/8S2q2O61xfpLQ
Oy61nFB/bsTwc2BcsDA+XKtGTdh7BE9hmEO1tnHIJnRzLIJMgcJO/2hjgV8D3Od0
6B7cqWNl8ucDZBLLUPDeaEge9XzYWsypIALMNg0H387pN0sAloHUe+1ONLWCLGK8
YutwkTJGzjqN14hPzHnXOwfq9tohuTLl+bMvLJU0MmVmm3c3Hr9RLuOdiLN6zJaz
r+8Pnb9MZmAByyasjXqWvHGeUaEKi5b+y+GPUVRnh0Ci7o1Ng+Cv1CgLG3TzcsAp
NvqI6s+YYti8i5238h33WlVGCtcUEEePlPoJIYRU09RU0hopMfnMqRl9qwD0BJsb
Dtspxnz80MfNetNY4/jUs2dJqvEc5KCGMkqa/l0zta/DII/hKwMYdGNAQHJA2xVe
ZjBNT8bZnk7vtEUZ74YIKXNXa6xHeXogCr2Q7EDayXeGUKTNnh3O0Lb6SUUoUvVX
bYfjuXuNaZP6ZU+TK1HwLzUO0KHFLhr9PnD3G6bG/Y/Xhenx533lC1C33eOwqUw7
YHlf67IzAj87k4vbUVG1IibILgArLAAa7sD+asC8NA1MksB+LNDKroNJMJd1/eVU
cZxIcbSFrbffpfXLHAptw2oZDN8MsNLnhyP26rZYcCp+FU5/qJ8Pcb3hTFhm27Bp
lVZwSOUbElByM/HXRbDifMAlTSDyzOmFksLaGcc9inAyqiRjwLrDs9Noi5AhZg4g
g4Hu8O2xcj2wTdHtIAX8aEU54MqvY5o8zT5XsRNJfngiwSZTDnhtBHWtumhXVjZd
oeBqenQM+4ODPn+5V5iQnx76y/5Pt0Evxrs7z2pSh7l1HKPLdBD11N76IGSSoJQf
WoV28vMeT+8O51cL6HwLh7Kyrj92fz8meLUAkGm+qhnl/Kok0N04OQT3poIZBUvg
phtNP0+ZNxdsVmkqRhHa7Z+G+OtPcQoEO4S12yvTxwlMfRVBw6i8/TV6eIHingfz
2CROZzcmImPzAe86wrleKpIYQ2HBiDCvsr9uAod0RIcClJv9oAEjOGVlsBpuOkLw
QhVApxdAlcHodbxGGNSx4hhy0O3qXFRkvXSZKywr5z2sdgukaFzmLBu6XqLIQPJP
+f8xHikWtvejS3HshayL/uw9vZaTFSSB+qQ6nBwstLueAcpN9qtgiPv4XSbfDd8x
2CjsiM9T6lsPHek+dPH4/rbIwio8+wzu2C02xVhO8fuvzdm+5YZkbX0qhNp2UaYo
NAeD79GIwIUNPtYRfTCoE+5r4NWCbocKiwZaTeeB79XcsnYrmP6MlmWlhzaeVoyg
QpBTIetoFwA3ohfg9WQjf5Oz56h6oj+RQcCJc6Kiw+cTFe5i7q0zzfouipKhIIS5
FxQ3AqApQZn4ejBtxs5eofMKqHplX62TOL1i9601SEFxOZ07ymX8eDy4ebexatGV
O4xOFUIBWTlcDjrvn+YxumtFGs4eJQGd+oz8dLZqfa8TIMeK/0Sio8RDgm+3CYaA
LxW3A4IpbgBzbU2p+Os7DlE+GYO6GnFsnvWHs54jS7IM4FWYry/N5ERbdKj7oukU
Qbgpy02pbGDa/erlH1adCv2+Xy+ppbPRImvURSvqsiJJB3cHbCtx0TNwdn9Ak1BP
NdUxSYvoZiuNmWSNWSvq+C9Z4PqX8Lov/XNxxDNUvuTVQphecv6Haf1o9VNLPopy
Y6LX0zZECw6NaJgoNMQ6OPnd8SxXEkbH+R0JAc8aqlVLjvtUSLY7xloKMke+rQOa
PWFtmkXH1cU/8kkjMeHM5yt4tDtd3s2BCM6MmwxAITNpXASKthLjhnBjQiEHLlea
ccLuMyLs8XjdJ8LmR4P1oJFzDjS6ZF2cV3NI5yrbcUCUi8s//IA2GiuN/zSN1h+l
d9BcNtHZR7ljt/0ipsrT5bCh6FQDTykQnJ2Fw4jCa9oG2BeGZ44qDoew9oGLk2/u
WOSGB2gLdFxJc7sXnC7vpXfhSRLV+iVb8168EFFLZks+sS1ZVFSruZ4BTQ2tDYvb
cL69r4PXSp2O7AQq1hMUexhWHaCkA9qU44rFCPdVIH2NJ0tUG1JQ5E0uxNE/3gwB
fL5iC/vKprxb8p312hGQaOMYYGeee7eYkguz/eo/Jcya+IE3lK27z/+1k6LTddd5
G26gMkZsVboCQQexL/4s6Rd2TWbFSQukytmTBMw51Z5tPxR8CjjEdAI9gEb5TAdC
CpZttpHG3Z1Uop3Kvko281JDYPHRmCVi9G8IKJTd/1IXuj3Gk3fx52Dmi0/CvkHK
7WBlX19S1jTxwgVTvKqgLSiA90pR38vSfL/94pr14vfxtKf/pqv381B9Yrln8YNj
goocbnai+lJp+5ZWfiGWqzxEqjXVwLU5ISRi2rW3dt85Q9tj4AdvIPDH7QL9kUYu
3n890zUSZ32Kk8hy2bvgDN2yYVu6RPQKjP+e4r5vLbfMYKwVXtIYtmn63GM1GUu/
qtKkZJ7/SfX8aqSDn1/yMfSR8knxI0SyK3nsZmCQujvnZkTPe3vqb1stehdqlIyf
X1QiwAeRHQIQOXS4iO4vSq/kvwCrUdGyVbYYVOgnTC288HJNXWiwi5sGI3/wYmCG
3V5AKJ2v+7QaQIl45fqpbvYShd8OXN5HiYCelHjKDBNhMHBknu+ONJEvu3IgSCTL
C859QjSOKWg7SHcpY3m+y4xpgBJpI88rxGfmcS/2nOAguPM0XV9QBSMPn/9YY+VF
LBM4FqEDuSUtEWdRR2R3SdaB5rMDvQj8DQH5xMh2ZovIpZ91oOy3jAxxJq0/c5qf
go4xsCpsRi8o8gKxoA3L8kENBuwi+XE77iu/Jns3jki1VXdFprribLfAJimUxnVv
gn9MOIFpYpfiiIox/7CmrURF6zHvKFuyInZF50e6Uy/K213isr/pFDNedc8k2+Jy
mLOqABhza1qKj8ule5tMs2O8Qzes1xDR1pU6fuICx6gJVC42fb2JEQTxwAmb8JKn
lRPF2wxt2tAURGtJAvPa52aoaG1xEp/UGDSO70WzSEAdrLoH3TmjVwRT0AeSnrzR
mUqM/Qs0aBT2Er37Ld2N5UJGOuYuwt1Kk/8c3oUTTWhJuAe3NNHF4mjTFeg9Kja+
X/I1wf8k2ptm3DX1l+K187AHFFNQz0PKWteQ7mv3+cLqiOKzUgwNjENJVlE5arhx
D/xHi8jsHGLshKs+QgWhzfNGxnxMvkgSH5cMEufJQtDEwWZi+w57IUi2Qfgno3Vz
qHjPZdV011FSkjEMsPyzKXOihlYQR8GqSNeznwi5uTE/iNfxkcy7VwYOV52s35bp
k7WB2i7FoHwPzS9POn/2rIiOXur/MKr1EAay6REF3cCk5t2xst8XmAlHc6d+eaQZ
phovSRINj1BpG+9ck1N3VBuCkY1FqL0xmop7JeN2ez9tvBKS/KITHOnCkP8LwKh/
6eBy8EuBndMcnp6P1oQw51b8r2nXvb//7uSlvK/7nipzB7oi+sQ3JR9v4wpQQtAi
9rj7zuwEnNCMfKtg0vFURkRoUsUxCYOK5axSMueb3iFAQRDAUfDbH9G7pDX4VZWM
11vpHkzp331FreIeykz9TVkCWfSz7o+I2O595T8UQo5pD2Arf3CixjsDey5EkZG3
x6XrD+s0xBO1Lv7XSt/G/59TW110Lh+IOhjDBI3cUfM/Jz6UBZL5vOqBexRs+Nco
TlRhPNb/LSKKVXVhc6vqGYegtekjYxXCgTW8KOaA7sUuEgQsc2w7sTJ+Tx13fg0R
BmdERgC71A7+AcO7lJOb0L2WJ5uAxT1H3uiBODeR/MHa31PWfz5HvQ2AS3NQbZZ9
zLoYW7fIKPioH+fDc9MNPmDAvlNi4KFnBkPSgDeW0HuK3ELMutV6CdsnOWCiSOSF
wyJO89xqfVN/XmCmcleziJKmZbQGLqhw04tENR6fHzipkY73EpPOMuWKugNOUpAL
TmR4Y1vrwzrj4kMWKzSVbnTrON4colgfGWtcJM6Nd4hIWUnXKTjTJl6iOXBaasq1
k1FdWcEr+gsDJ0LW8aD9r/8m94ipsrgCiaLIFGJ+JKlxS1IaBr+ah/uZK5UKilcn
Hzyjw7xQ88p+xuEjx3yaQ7+J/cS4Z7sdcLA65ml1YUb5URHabW99IK11boLYcOCn
TckgYP6GldUnXBiKdpKYtKMu4FDjFBHS8alhfJvcgL0NUZGYAQW8Q4ttrOnhfQql
sq3d0iKRoGFvatlf/hY0nbf6xPE2pCXxeAvBBlvcNsLB8IeIzv1pCUKRj75FSc8A
NVU+54DmTM32gLbwE+FF0BA4fRjBWc8C5amiT0Nrgyr0/mjZA3aQJ9fjQWziUPV4
VJzzSn2xI+BQoQUmThac4KY+GXxK9PtVAXPspISUYsEa6Lo1tkAZWCLAVc1gYJ7U
XtI7fxdMaoSRx0XZBPZMUY0o4hMdqk5pO7BD2Sx+H1ScAOJQm790cjzsnJelbcOc
hj5oS8Kh4tffZbY5VYu4DWvKtZsRWnCgBZNjGhArGi0ho2X2LxYPLxhD0wJhzF55
0cdIf5qiBjNYiuh0E3Vto5e+5uKwcLz3Ly9DUqkfri/12HFXAeK/1Z5MD1o+2VHP
JnUdUTrg32lY7hjMGROhcpDUFyOX+Xs7bo90DHOvWOeyovZy6tfowlmVKZgzWqi0
ONBf8sobMD2AO3QlCV9eVUanRgt3K2vPOMhC22wJK8zL5/XIEbMwgyWjHSE1/tIj
9fEjH09blI/70AVC7BRH2tq/rc25DlXh2siw2OeP+PVTcfXTEetP8zhqnUtqn6se
8uoH8xefP866Fx3rh2Y4Ba29Vvw1UyhdJhGWa8MHdh+ElwbqeVAa6Gez3wPMJiNt
mvibe2QY0PPJVFtzB3stwsnCv3+mD7qLpfx1EdLsivyYA+DNe56l7bzZ6//wjeKe
a0yoeL2Iwuo5JjTtbA+GiWT/xlZMViprQnt6KcPk4EEBuP9G/Pid+3K5cYItdHNN
Dct7t631+w5WrmO6K7ky0M8BgS4Phl7+FJ4xGMWd91VmPehCEtHFg1RZiFNEHLGS
1ip62EdhjgQ8Pxyujzr3bNX+8R3+BTsxsSOYX/MF06j+UYVUzZn61rLzq0MpSVCs
jJiCmMW16zVZJn8LZqchQZvflgLf6/ZVyHZmOrv7XzkeItBieuxq3dlJ+/GTgJ0T
Em4PNTzTe8v8ZeoSdaDJaw7HJ5jXyQ/ksEc0zbzSwgMudPI3Ap8gwfXR8YADZnj8
552SZieE820+/1GHx+gFBsso6Q1kzON6evIMLhDFSfR0ieyQ+2C0PwpnXyv1TdHi
6aKrugVEzeqgdzka5A5egOkL4XYootXgXTi3MqEqDHZ/fC+DoYx1k2ptAMCFG1T7
f5KsunrcEhl0RxWQchzsV782ChzbbXyKm5mzCNYKzt96r9uMtr8/alKY5+i350p/
4X3I7jw71QF4Sk9Qndc0E/+RR8O3Hcx/efeb9CMgxR2s99ewIgfjjwUUq7p7HSyl
JdCmgQKM1QU3h4XzJcn0/KASJNUwXQn6a23vsryMl8cAy3Zw+JsYdCYP1ESbPzUi
Gg9F5hSDVcvvL4kl5iP6ydH6mLSXluwDV9M76Lr3bgn5i4xRJdblxSt1/t/eUGGG
IjR8UXXenNsJTPZGYq1dp7FRn8IL2GqZMv6ORdFSKeGAgHzsHLN0jSbXfyxUkH6I
rRAqb7WdiO7Q8E4OS958I6vvgFQXHuKhFCzAJFMfKGkejlkgOo/K0qVWZfDBTlhF
4gNgsoP56Q/Tz6m1JLdwcVX2VA2JxZg2LS2NBQtbjzq0fU/Jh+uQwNMKke2bMOmQ
4K4qSiGDts0NmDGa1XvVztxDb3GWwA3U/a263gFUyeJS1Ipv5buQ354PK16XKqgm
wjT/cNNQ1Rssw1kikY1N9QvtlJyAlaGD2DxQeKjqoyc9kYx9G99x87pJZ1fC4exW
TABIarcwihiIutw1o8PP6csgFYm5Zp7Eg/KulJyKJUqdx44aEC3CVBrVHKhnhLHJ
baHs/1c8h7oOKvC/cTgLXpsRm/Duqa8did1/RneskDxk1QDTRC/pQc2KOTdlP/Av
8y8sqzMuyieBnM4uNb2yC1xVhCojtCZb3P+0QBRYCIxwEQHa+egSuXc8SatAPAls
HJvca4RYJeAU6wMd2g3J8hoJVESPbb5mbyD5On1Y5Rf4bJsAem/TaRzThEZ7h/Db
/5w3yKM02E1V7VSFNZPcktybXCyeRu1ctpXfJB+yub7QjVqFpKWYNli7BCcqtUXJ
kcOwia5LqhJZrUCk0368jBak8Mdidg4oTei8QFPzxqytSLq946xwAf8bvNjrSMJ5
q0Det+I8UaNCdd3N6pmvJoZ+2DAqVHcRhgcYkDl5DpgTHiAOLyVRkEJDZIju3tA3
6Joh/yJEuUgfYp7Rnl5QoADH2sP9BIXfy2Fh1mdPnEoyDc4FNGAmU7yXbNwkZI1Q
IB0sycDDODHgZB7iF7hOA3i3r8jfLVEepUURglwA3O7v90AJvMf6XpnSyTC8zC1l
X4XF1zQZ1y/RJyametWxs7fVTm4qxXMrMwc/vaiH/afeDD55AqqppIrTZvRu/LOa
my6d4eL745G4+xtotV0knvuTCZha46wusX1PkxRdKLZSeqy5HqpIALKiT0YAk4FX
jANUOITg54HZNlJM3miycGxnrRj6NQhGU1x3YjajffJ+H7HB+CoZ8C3EI6vaCS8+
zfxlMT52gZxqzJ1RiMcy/JkITAj0cfQhMt+AZIJirJpa6PuVTQT9DO+zlDeH+K9X
IWsrI5kAl36VgaNbXl7pXPVHxgMGuKawklyzVp/BSHLA9SQR4410wNAO2li0+PT6
DNRWB3X71/Fvp2HxybiiO+8xf0EcRGwNWRfiUnYL+fz8zyEeO/rgwphFJ6DM6GvM
Z27lVxPnb27os2jAkWU/ePXvxTIOAZcxja17G6eF/VpPlSP5V7pmguLuwEjPxSwP
e/Y8cf+fd4M9zDphEmuyL9JNnu5bi+sbeeVJGj2/WMTW+FzP5byxNBNtmZsKm/SL
sIOLtSb8UJFf/OmCoxzkupD065FR2a5Mj9Llrg3BW1O/yYmcCVnFZDcb9FgGlfxp
JqdUuLBuji7N25JokQ0aSsTz8sjFJM32VtEuMJfO/CLAL63NwXBq7FTYdVjOYNMn
Fiv+maP9sfkmEpGZ0tIlT+8Wl1UmjbTE+XSHmWBy3HBD1rR1iAB+RdaTsoAlOwXB
b7D8HG4GhI2ozNCo549hIRvhT9M1MKZWSujXC+RSzJ0FzV+RWCGApmVWdkJyhkdY
U0IGloWIcw+5mK79/7Z6akcoxk8l7HfHO2ZRE4yrn3+avE1i7whC1emZu3JtGCTE
y9OkYW4x1wDS149GUh45TTp9tX2LZa9zGyeRaXKsJS/Xmse1scNir9RViY2zmXb/
diVFoI5XRLSKgZDv4m1wmV8jpSTQxyrULcjOHYcOa4wTKa445TAPc1940xAXHncN
aDNt/iRJvRdXiTVzcCO+d/gD32RgNsgSk00HwL1f5BqnoPEufRpQFRD9Z1N9G55u
GWbHyupBw21emn6mVuWKnWzfRRTJ1PrReRX+0U/ENEO7VqjEctVw305TLgGJs28s
Ki8lcmbjpkHnCwMMM074PyWd1Z3sAwf2fz/NGwz7kVo90Nsjbi2UToFr1ACNsYDf
n2WrJsa9o501qc+cXGZdwKdZDsTOH1vSceBXBqdAzl0wa2FSDYS+yqb9RPuysnmn
u4XJlsoKi0C7h+lZz2jM6PBfV5UEuE+MhaAdxRb/lJZwDo2biwRtIP/bSakT6N0L
3ZtJUHm7sd2BGafk3U2aJsAgZdfARaOhjymaCNqAXd7vaIZtxTE8rBF2NcVRf7gi
AP5pRb2ehboRoZ2jw7S6t7klrQkJhcmHhn/3IpaQFokcQld3DZnz2SZPmqvsMhtn
0Kk8V2g0ZkIKJb7nZz+mGhd9xHQQaBlwRXFKyhHTN7IjXQ6wOEmuVBNH3YVeAsbQ
3YX09ILcL59AlWskDU1IAN/wWm1MPyuRy7MHJ8iwPIn17ntMH/LAL/lAvf5PVCNw
KQbuMSK2wnTaIMUktjnnG2aKLQXkFP1lBEUWnA7KymijbPUCJuFSPOfyl4NcRGxQ
lEjHwKkxkAErQIVLCNivwvFeVn4+DNbdxkDZzecfdreKWBPOALWj03+nng4WLAOI
cg4RtbYn/C0+/71+PYrWjzKKCPbbe+FVsq60TPQ/FsKzZmp5Hq88Y/+6mnaxKNdb
RkR96j+/1PhLp4KtGudUglh5ZFD0olQA7cmq9Tk/XrQzjgPyTfH+gHdb3HrKQzU2
Qa2cZp6Jw9LFz3W+8zZAheQxfc4/7l0wimikN7hxQSyL0UPs39mDR6WkMPil5jWM
TFBSKpFEvBTiFcJIKkL9JiP8B01H/Rp4EGGxL4Klg0Mb4U5g6vscL9fVc0spPp2P
UO3sTjBD/Tckv+2e6E1osq/lCtrE7bkA9yOSBVp8I8iye8xrsaVGARsYL31jHogT
tHJOCnrdvysqj/IzfqQpO/a7gRc9WyBfMbmQPPxO2ZZvAq5CBSYNTXOYbQosX3oW
+9ft51YBOovmfL81L6tMzglV/FjVilnivHZUSVd8VquzwmD9uda0vlqfeD6EuOV8
MSGl3xijZLJrmCTBtUtQi4Dnxdyln2tI37OUoU7NQWMLOV7Lv8+YMoESnMm5T0yc
pIFzV37RauT8Qn4gtXU9SquK3+sxEqrjOZHoI47KJyDD22kKKfjMOfgGvY+T2tTh
/KPI8iHt0dDIjaCr06ZqHMcyUblJszBHXPeutHhgSmEG+6o4VeP76w8IKZB7QGvE
Jr0VXLA1xLSYDNXwK9+SiXU8Qh/dVO7/QtVHQCu0nSmls7MTxfajI9ULC/0l+u3o
yybmc4fbptqQDPgksGoONLyq1J3K0qXCW+NZFSF3sMtoxf4lfHz2kSCYSO/nHyos
sY3xJl3m4YPrKWTnIhTXE7GvOaiThJnGwfZOkIquCmzNUWDBobb5xJr/gGLBknOh
49gsU8GAV8wsO9vpaFmTUgRz2rqtsyyi2g+bVTVdqI6oHq3czygdNW8aBzbsxAZB
YM7V1aOtzrC5BwBsEnsN7J7Q6ZTU2V1y8YNxXBEkobyTCYcXUWq8JYWwglDwJW2i
4zWbSzwilSXMXAHeZTx0RE/1L8LWqknq63gxknf36GTd4YzHgLFQDe1nSCpmp62Y
rFdK5lK1TqdE0hfirXMoEYmS+BN1+vSAiwrBeIiBLx9N4BBrsLefAyPs9el4J/fK
Nr8+ndiXKVvOXKYYPgcVwlOl6lM+nbNDj/SgBtGDCMf8Qw9PqmqBxcKk0jS3qUt4
69T7Xjf94dnrhV6xi2O82ursnt5t5P13GtSBU/6xOhYeMeSYwlBLa0kAGw745c+Q
tDGLZQKQTU7SN0bmvLAaTfEklVIvYFZ0ZW8zxVHgPvBqtxUwuytKCcuMXzC3hEse
uh6s9vKjZW4/qyoRLT9wRnyyQRfMmbnck7mo+Zer0HWVFP0h8eMAYaTPu+5fvQJP
C7DoucNPjnX2frLuQz7g+vU0t6Dhltn7FSVNAQcBD0gasUU41qgcmNFbNHepNwiN
s38NyGOYMkx/JHVnKfAvfFlRKORP6NLUrw7Iwfqv/J+9dk+Fa9YkbfOxVoCui66Q
wui9wKucrZxUGNOSzwI1SfzVkVW3YP1/A4Qfw4BheoULPbZnJg4L/CKk/sYFHu9I
6jtUgojZxeRsSTTfnGgD7ziWZK0SnmzprWid3267ksvH8pOWJZ7eHB+6vBmQfb1N
B554QkidipWotNZCeH6okvDrvxbIOsjwL3OkwlEBLsDxI0IwosSa8XBSER2qUQSx
7lyRcrTKYVx/7NQ7UPZ1TiWA/jvMUCGkwW4pUZZyULGZ7LwdQrc9RGLJeH5LVs3R
xRw3Em4Q5l8ViE5iSD4+BJ9zqcyeq5aCOi5WklbvlOg6XS5ivP2szw1bbXljoGmF
C80XUxuxUiwgVPxlZguVV2WzulqfGY+MsJ3c8m1Nl+y4+LzbrGMAe+6d4JnruiyK
JsYnUG6OTTay+Uazw6QtgwcMB9FIOk0WJtpSaUhLeEiXvEUBsSpPDJAiVisXRq5Q
4HfQ4Ot12nlG8ZTDjuWeAl2f6COmuAoDZXOYVusgDDoElmn3WaVqHlUkkUzwwOlI
QkPz/0Pvh2JgVvftjCc/EzRY6cf1Zk1I/sjTJi9uE/diEs8b0vQbYEVPgFio7/Zn
XzpnqheG9C8rS0KpLMBzCsNiON2UPxOW7mlaQC12HIfN24qNEbxUydb5w2BA0YnP
KWtClxQ6/bgMMtgGCkMYH/+YrxAdmZhmssFujEtUhofAvr/gS1NFzeS1yevhmgQH
2OQLx4P4iBS06FaZq82Dlj2V4Hi69/Ab91GNm8YRXuLXrEJ9sSh2oubHQ9BzNypH
/OTZz/hLxeWIJlZ/BgpFZgn1TsF2ZXGqAiIBk5TWJ2touKwHfIE5QYMoIJB9MwJs
6XruVcZiLw4T5A9Ad7aAxJ22MTZRsLC9YcmXxKp629zWWvUAMUfxgdI3HmbEhRi3
OYkRUQm1bPE651jOG7dqf0jVtjI+K0yeATpEBupABX5FpThtptG4g8gZxSYcWbmb
Y4QGoSaRjuFAFNTEGacdY7q7Cj/vVFHhWS2St9PbJA8INjhP/Bz76fRkGsyP8UNZ
cACxSmndA81GakRJd+kIi5kNVFKK/+TXbhjP1K7cs6RLT+su2u8gJZliXt7vEyJz
/2fNEuZXz8MKJvJN2WSgXrAUjH1f7RsWj4t8/OHEqscFjPz/lUztP7o/qvD5KNnL
EJkbnQivJNtQvt2fo0BO2/4R7KZx5iwlwC/2MVRiB+P0apUJyAv+ZZDZ2i5B52I/
49spzxGy5Ze9sx/m+7LmxIjBXUkOH8rxjMoRypG6cktmChDkcW7DljCzeef6Aash
crvjxtwUQFpuiSFrhKjrf21GoI5ONVXmFjC+DqJHz2BQG7G86Lbqh5fvLK/NQWyn
jBrX9a2dEsso4E0Qw8pv1oykUq1WvrCxaCoOiAtNhYeteuQ+mLuXyz+pxJc+IsZc
hNmgMnRrYSGlzo2/bhH9sPbs88Chkgcibxd539wi21y+sf51twP8PulOXsWxjVdN
+XMChk8r6mv1OnZiKy0/VemTswk42aPvl2HT9M/AFwB0CH0xBRCwCgCXeZ6SJv0K
5B3jbIXaGJcyVMLClcvdUysRkX+m2xDLXz1Cjt/4UCavDRolu2io12thDTJAFG+j
q2ZecWyVE68JMzX2CKvmnNlaOAc9dOyNqJzya3TMxhXnUz6YZUpiBrcb125UcPPt
op2C1cqP9mdcCfMXyMlSTOC1VMhcLCpDDF56NGocQxrftnm1BQSBiqyEJ7Y/v0Mt
qX4bE6PfpumzKk1ZEf7Fnq4AvbZJShtkZcJW6g8sfWEU/5/jYIPjYspHHu2EjwNa
tAtEo914NpVeWxCRw7DcsuHzLzlZLpNyDr8ydtoDlajt3gCx1NWOz4lhVOiYYyaj
0x8/gQNjaJEwtwghteHSVBhfWlk645l0U8Hf9RVkS9B98AfFobbzDSGueZTr345K
7zTm1yTlHKL4oDH/nGV5KJx6pqgLYI6Tg8Z5PsH6gkbmA/I0srJaDpqgQnPSs+ZV
cgJqiLNIroCfu7Rrww0H5+l6V6Fo1/x9D7oXbhoeYmt37SNSEor+FxUS6AADcZcV
BVyscLij+I/t2uuW0njqSdvBT7pJfeztBPwca7lRFBUn0IHbDkR3NoT8vL/hE0QR
rorEV3JWkLwnTDX2+dGQYJWc3ZwoOetQCardsN0kLOaWgDTrUsOeFjaetQJhq+pn
5DSkVJbBuq8cE2qqkKePBQHRnkZ1/joBuammow/aqvMSp21z6XJAowpkf8+RsZAv
rxzNGi5KX7lq00ECdhDLrhBLDkfCh01BMnXNez1a46CL3qjAXy3EIFtzlw5HBvaR
sBtTEeCfLvFjengUG3tJeNnhNdm2DQUN4Fk5rV8RVdtN3uShIjENzyMzAxX5VWZT
yECN+FmJwU98Zyn1UMW3V8tq8hUJh4GcyynTiEFCuafPHbmQ/JBh6L3SeA9iEaa0
z04GEg6Xly5vKsZP/jqNxR7YdvXGElGere49/tWI6NLtc1Ny+H7Tm3KFHsv7UKRz
XKIbonotDq/p2PFLf0Ri6HWrVZm8BKrYDr9hbfR7f6o03/Ici17QxzpNPTkYigFL
ECh3Jcp/g4D0r4slCj9wFyoeITd4lbSyOyXSB5jfxQxw4I8AqI5BRTsKAd74Cthh
u1QDAYbBrxfNroLK3FWuPu/HejNe0ebpJNjbKTsJDob6jZAXV1kabDP+m1zWvjF6
CqCzK3v/nO0sQaUuVmt5HZpwgsMukZrf+p6SdDhxQhuUOKP9wZeDcfplGbeHDF8F
CVGo/9t3yPI1N4l0HvJRhst4k+eGZMz9GdrSZIR2JgTkXe2Kw5tNu8IdLdA0jC1Z
3H910OncdOBGDV03bpuqaKHRbctB/nUXS32CcPOFjQX+dBjvHvdZbvvf9erWwZY3
GGF5PvyBLEYck1rlKvlNR6TB82JN31Q5texCrxuegyzjXcZVfYlHX7TOeJvPprEW
iKS0oT599FHkHqubgldqGm6M4UmysokiMP5N4acFEgX1d0P7nBfaK+s7ZYQpkTYt
FQtUUN5vUgqW6SM4eHpCFLe6q+gm6r3HUiTHaU//Q9h9KxQOs9yMCb9Lxs5ATLxS
3SKoisyZKyRJiWQS0mV7+MDNDNvTx1w57bddsCqvPisqM8cRE9ffzogwMNAY5gGe
Tq+e3xl3m+dyMm87PMnMg6FDvi39iODIvvWqe8R/1op91SSO8Wgzu0uUCYEyBHiY
LKUkjvmO0sQfQC5bTWeDOjqRlKTxL1Hf/yW6hdtO4pKOwGY+fyKbOL0YRNI0cmiR
H0emCA5Z/25vc30cHBcrJNFiSgl9Stg1GjtDM6skG4WmuqWQpQN8AH840gy7/rsS
qLejicrU5N9pvFZLSHS58xXSEKKx5sDSLkR14o1IKaxs7w3vcKM9WeGDtoNN3awG
+8UAnzEewLIQ3StJnBZZwpvVfm6ycznNE10Loszk91BK54WMPfWgXsBh62Kv2V88
SZs49/qELJL7m7+LD6KSkZn2mMFeN8l2U/i5cMiUPWcRPLmH0ZpWBOK8bc0Mfl0N
Tf86am8oyxaI9L+bPq6tNoyM682TTLVdN1P38vsNxjCIGEhrUT+NaEBWbW7tmF4p
JEo3QazHYfUfdW10uNLRvp3zghLODoTgL28FGhgGMvhHJSDZ/QdJto1dyeteaMOi
bKEpULM9Ps6ph0Y7F0aRYW3nLAJL22BFRqqJUbG+fnDgCanThwEbUHVB0XMTtabS
UWxyBtoXWWPEQ7f0SOs9OUOvtYjFqizr6JcQSQK/+zZffM0KteudqpdEZ46PXr2L
kSRCqAqVJw4p9l03T0zGpbfBxsI7RxXAInsXcsfvyY18qavHwGu/7CMts1nPwR+7
zn/zxsUUw9IsdmqMa1jSqu3TiofoCGIK1aPuvZIfIzy/spnD7DXEjJ76aHxkZcau
KUI3ojA7yu2TbMXIZcc5E6W2IFYN9tNeINgaCkwuHT3tzPNimILk/GRld8F70FS8
UL+VDVLENI9N+n6I6C+I7m195bzvfuD/uTt/8P3JRIrLo5jF2sjMKVPaU6VtsKuL
E5COJ318dbtTM3nMfe+75tgUtTIsh2819lI4ETNGG4jifp6inE2paA7AS5fN774A
NRhsYTss+GMtwmykFmr7GT9bHwX0swO9EONOGOMGQRayH1wNqCpSHgndBs2Fj++w
zyYv+MMwEMwVL80oEuQCv6u/EUJ8dKbrMQniC6Gej/Imv2YRBnCUkdgpw+Uh0eQK
K+t7pG3ksspVv8rAqIJMfgzXtXXEsXU6q88pDUmRcRgQ4XYI7eLdsrOUlWfHfQPO
DaTM6cfoYoM5fWWl3IiBU7FSTQ+GvgxVMXhXAlDO+6ezIj99F/o1GZYpseB7AG4E
ZvBK+k98EhjIdIWrESjmu3S9YQyN8cVTD5+1vdMciWxCpTWykMpnumzniClkmSCR
wrHBm+RQGf8q4EZgmOxuK0q0VE5+vEbwGQzFQnLBc9uUpx3noMDoiay3DWQmoqc8
Yd0PSMmzR7E1zzrkO7Knu5VQEsyBHqA7pOhR+CQuvSby77Be68cZQRtvBtQOsvgi
kbZVVfmvFkZXuvCrQih0XLV1zKCuUr+Q6Jgp82cTk2n0Iv6/+5PvfaQX4sB3f20b
nX8N04DUXz79ZmPoQ7OTABaUxCGEcRIZq+wDmOnx6gX1nUVQ3eidLfDYEDbBkYjm
M62qGrtYutJot/LfT/aE/tSHbS+k0hbX61wVAgfbNHRdScsDRwxGXvwjX/gEV+yW
6b3B1/5iI+f/TPDzfnrz8QYKZc53SwLikdCXNYmfYj+wh167MeW4xdbWx4XjCzKV
M8rRHL/5Jw3/NAf68uubo0iN14rSXQVbmbmkyKb1BM9Q8k00tvRFZYgPk/HgHl5x
b2nqzUBdvbrKtHj9I5PsEGruj+hP5xwltrQZlfGF3fWCWpucXhuwqymOdY6C0Zn5
vwVxE26LSeQVSssS75avLymSzaK7wUIcZEUty8AdpJnz/iDtzHatRVfK8lxuLXhG
CZS4adyehcVE6VfLzVRARPKm6cF79ldLpdaEznhmsEb05fvbQyCudgdaY5moD9R0
oujByO4PmvK30mGTaAAJET2Bgu5Qi3X7XdK4/df484iI1cTiS3KlblJNH6xYfurr
A8aP0tJDAnWP4p0qhQ6Lu/E0XXsCy7rWDFuyofZEnvXO63s03QXV6uNWN+XUAwVJ
3H1kdsA8N+17IRmn11XDcuCCcpzDKSVilLNcPoBqJT/ktyyFswaBY3g2Qok6Xm/6
XrNLAPun13mKuLOMAQVLNZnJqi+oUwlLM1XHkjiUE5uhUFZoklMnEvdNOYLRnGlq
WJWFCiw4QAiNXneQ2vbgP9j6QxURn9g3ZO7zrSumfHzTwRqDAsK9pFq/Dsxhzxln
fFUuOOCa3LGZzF9pHsvvJH/zOhhQ+Ot76gy6JWFVYUXbLlEYQjNpkUFHz8FPHqhz
p39GaoIBy8TAktPS/JDkF39U1c4E1jpKDZnXVeCfhZdkomuSSlEQRtzl4B+3q2r7
UEo03wqdGV59Usf3wOt9eiycdzCWyo57Rg3wHwG6AFiP8mldqg8Qat/XWRANp/R9
0oNu6rxjIC/odXfK5/XmWtQ6LNWvrD2IfprVm9/BYZ9F1hYoceWvUytrjUEn3Q+s
BcsjD7MmHWqKHgUbcIEw24AGohrzELrCeT22aGeCtGmi+rGfWAT6Ug4WT5SPwqAa
A0xGWiQ01xXN+HMrwC7y+AHT3miRcXIgHrI71rr94uQqNHe86OtTdgvUjXPmK5u3
ZYAD+ButrkGEH5tiizD7PrDIv4juEnPahRJAAmaQnCMxiMVJVUIBNu9I/NGOTKlM
U38oH+oVlvXml25pi4nFJO25Wh2F/0mT/W10EPUAylsAOksptMnIBlnMuAQmlvyr
oQoxE3iZ2BLbI0WHjGrg0rJG+lMA3FAlXym4Rw4JurHj157GdPXCe64TKlSNlSzD
pXy1F25Cfb0R5i0WGsZLy+Yx+lK5GIPuTxAVmdW2+PiFQvV8GWisIRyWf519Fmd+
ztpTLMEpst4QYuh+9ncG1h4feHfaDmgAowCju+e30IybnDwFRKtBLP2NARUNeJJB
YeGaz9SdDI/D2OWoNGDzsPFmBCU7/wHXkoughwqXzBkBazNJmRUvlgHdUncQt/mR
1/1RmEXA+dxEADmmz2HxmfyE9RLFh6pWnRHfEBy4ndubPZ9qnnhNyxwlnQIqXtV4
pswy08mMzGBgMifYDcsXYPoP9iNVRfcEr8CgI3ZGs5rlqMOxbKeig9DoOa/UNqyz
9SboSxLnlQJLIiE7OvUlMffbvjmsww4Byxhb/wDjIpbL0PIPX2xV6ZZts+Ac6/FF
LnUdfgmxtocqll/yK1z03pvZQxivsTh7tFJJtetqRvZ+hmhLu9T9xODDKrB546rE
HTyj1zwP/K10DujE1gkGnZXmRyzUG/Bv/ezHXedCN7mAO4gZfJqxCCiTmhb31kAj
UOVlCiGBI/XhOVMd77Vj2b5gujmXiayg+erm36Bj5Y+Kt2E+40ro8YIowv9RjUsj
ZiTMB01qNblD762vbsFAYfB4uNDHmoPcga07YP/zBkcHy8wAeiLFtEtDDKfizPNz
/GxDT9FOpVdKQOpFEMzyCckrERZ8Y44HAEfapsnG5cdb6yr+1yQ7Bc67p7I01IHp
3KdK44lEnmQfYBcEXgflgRsm92i9ABHBzEjnA/lLDpgtOJBwOLpsgMxiEPMfckpq
OXuaF23qcoEAlLKyxKDiFNzm7W0IN+0GoCM3uKUdhsiEJF0/Dx6ZK6SEoJrjwjtQ
9IraY3GEu2FGeBn2DibWzNdCIXbpk7pHU3zofTK6v4frZbQG5n/NSZnuKhtXCdXm
Ok/fGd5TdPBVnQL03+mNswI3+wivKQKlI5kNBZvr5LtlJILxCdUpkyV08+R7nuGR
eMv6PCXnoc/0Vl06vQ6ac1HkIVTw4pxpFW574zZbVJqE18e5RbrosrJ34Axr1rRQ
mLsfSh6aw58gPNbfbn7MIY+Mg1HyC5RXEA8taqVVp9xVxuPhjf8nFQnrrGhDEoVJ
1h/U230zWqGgHFVbCv9B1wv+0gcMTy56GQrUgUFBBlBVkzPyIDNqnCRQk6yhz8x4
jirt6OC7OJhsPgPocRcUEyvg3swprjkZVAae80WzsHjeTCZmpBT9aq78Rs66rgM8
RYkfwoBjT3QQnUkDLegTFXkDZHQcE3GFAcCAm16Z38u7NWS1neSgrLuP1/gfABsx
9qwjKtvpX+rBhwdyZ2mIG3+upiyvpDjmrZxApyiU1iMx6+KHFt2/jxBBvYbQGYPn
kgpLWIqEsB0+fQiStWttsgyV1Pmh95ecPGRlfDHcejfHjqkSltT6Srqz/JsLkP4W
sCI84essqCR+IN3ena3fiw0DKUC+ie+TjA4t/LBW0yWDZxJIrOaGvaYkku9/s0Yq
dP4tgT0BVtBlf7YkcYeCb0xsQHigB3fdYx1ycvLzJNjHSrLm14LDt6vYEB6dbRZJ
9kxVehCih86JTmskvhi1M2kupSU5By4IsiGtJEAI2gilx6R6EjgaJQSCbfkXtfBS
dnN2NE1relYoCumeY0p509hJB1ByO5fKsXGzasbFfL4OAuRmEWpOUI1gs7miZSv3
okXpEfT0S6B43cZpcp/3v9wHTc3svs+7fQE2pIhjYKecpigN8u9uuaeJljQ4EfUk
GyhS8Tz4Oy/BkYpYsEeeLXO3Lgi89qQsg5YGN4k5vflQO4kiP3Kkufu8HLlUKI5q
tAfljY12P7mAMSTG6P9LeiDG8ucWxYcRK/Bh/mVN0J+XHmNFYgF5RhBU8t7pM3jD
KxcT6+Jlqd4hIbidqx1RCgEjIBo00Ji7MdlyewiBhfp1FgGV/rf3ye4wpfaoGPpJ
ZNhNqg95b8KYSAhKP0xI3HAdVYK8VHHidfIwcYQ9rSWJUL8c8CKpUAmF7U2Z79+d
w2P1cI8SN5d655x6vxQ35tsB/hbM1pdYR0Y2Sk77hVdWp+9ey1eYq4bbDPYZna5F
inrOdbwR5Yp9gWInbxk9oZ2Saqol8f+KBDbsjmezhAo8r14PZs2UhRfCJ/zi0CNy
RK3b2iB6t6qXjEJkQ23aQ0Yqx5z6rC0mMD2oAFC+mLJhjrV8UUeV148gJdm9xxXf
pK2U2VttnXrjBCpOqqVcC/5QkIzZ8HOK7d3fo7bm7JCI3p7AbhJFnXAVmkVWBrJH
XOFDAlY8C18Gpj7X6KX4CKZmaCs9SrwTWjzatij9vvMlhloq7N9BhhIPGCDIpk2P
q/e63dupHDPu1eDd11rWQQjyGkEIuQnt3p3FzmSog+1SA6bmUXDwFPTAnxlG8Fxj
MFCsbJRTMwC376Ap1wMwryb2iJZsHTrLFX53zMw1Uv+4bLacpeMKjITGyjmCXUA5
h/k78BzSb2iIP0N6uTn4JZYPlAzjrP9DoA38IsBoM6IgbfKDbjOH6Q8TuLFNe6wi
OOK8kKcMMkPkELsW3ddUErV/hDLeYs8oDt77aoFi3QLQEdTHW5XFbpZhcMlJ9W6v
DBK/gdTXw4yhqB+RVzjbsTs+Y2GijqLn81zZMCn0RELQKew89FR64cQ8+wcmA6gq
GKYgZYjxE5JRqbSw4I/JgswRevWik2IDoXhL7Ksbo7k2JUuaJ/X1l8ikxKkvHXQB
eTOMnzVj6RGHafkqjPFcIukO+4adTZ6YSCyV+k91eDfYgH91zlILuulgeWHMcN/U
gnRTmb+PzzmJnYQcSU9NLBnL5Hm8uNIsuZ9Wy/NsxXjdCwgqN6hhp/umXiIRH5TM
Maanx7aEY6epyPr2zY7WkCN2YxBTQ4vLWLr1xc91sC9dDGScSKIo5KlGnKdrKTCu
kEH54Ccx0z3RFZ/8ekQ2hdxSVNCrIfO5N5GtUh6cGFpYTY06NYpWrgblvtLK4bTR
1YeyQrkuWR8IiqptRFimQTsKygaPfmwi9FK0FLLZ9HrcNtxf3bE+jsRL1JP4aow/
8+DJWljagWsjYmUPVlR8zDCSnJS7TMPtF2mdXxI3Ky9eiiKj3KVl9B2WNvevzp9T
ao1FwNJMKnblMoTdXuSNOBAQqx5wJE+PvYczdiFxaWEogjL8/f5Z8UvzFd9cBcub
ABxndTcZn8/JLTYv9k1dDE3pN7TEidMi/Ho2Zujr0n8OoHiBq3A4xLCevhrEr148
OiLPoyzB0JGvQ8dyQV79aeP09IAnIzFznLHbpXFKXdqpgd5CZIpm/AeNYXFuOccg
vspPswc109oE+JSHl/+kxtxT7s904tZsGogn8Pf8+2GxT1Q4jC5MFVEh8lyl5h5N
qGaK8d6uWitHDlqu+bX4Km4FO63jZ8wujFd9qxGLNqbc2PTPhl+lNKSg9LJNWRty
0sha7v2hV4gP/TvJ/2k3q3BUbRfe5MKk7nwlKgP/ZcX3fdt4PtgUFlymeXx4MlCG
6ynApq5p3ddfHnQ9WuZjPCEF7BqM6QFZE1zpsOYWunp8Crg4N1/0MQQLTlne7C6b
gEc+bkPG6lp6xW9Sn/rAHBjp2iRf7/hMpmHamJhoheMnJGU4Korr1FBO8Svaan8+
xRz/AFnpI20//PPsy/lf5MJtPelXYZ7OTAneIQ5F8R3jGdo1HfRhlWW8Rh7LxwP5
7MhawqTm4dRQkeqNNHJuhNSqpypr9nkiprKlBjd/8+UdhXPd6cxtNUC07VlSRIHn
Lh7J0natez86sy322IsehZyBo6NrBBtCNvalr13xnaB8zLs/DI+EMxmuq3mH7nYi
hLbN/qiZmRmyWXz5LLjSUhGfGiD7uqDMcYUFeXBqdZNo9XBddP3fmSFwihhkdRvx
a/5rPW14et1bYaEmnk3gcuNneCNd4JIEvbGHrDwb0oo3T9Znp8OijX1S+HbwdIt7
+9qBAb/uj9Lp0Bu/SmQl8Lkm4+HZSRm5yWfGHHU2HQtOt0uRw3JwwguCjESQZ4kZ
F1VwpfDBjnHF+U+n0LJRA0mxXsEuaArxJStwb1k8uWOYPUfi0mAJe7yIoisOAtGc
/Wkb0kepdcnlZtYV2/411iA81qauvjM4cVz1a/y7z6JCFzgRcLLfKaRzJ016aGYc
VTTJ7EnX2LutZq8cnWWcFo77eCijWLB+pOxtD+zMxQtuDdyx4e9eMkfjv2cNrFvG
+US8YK1t9vzkd2uK+TB6FtKzmxEKs1L0ueQaR234x5d/VDdOe+DFQxdQSllPOg7J
Xk/SavnBWildR5+AkuXTc2/gWKNex0zOg1dLN8hDpf7NrEM8z2IhgUdt5Y9PPBkV
IjOs1RHIZAkE7eTZ+dmGliZ6FLaEKDdwkYUSlNES+bJpncos7fbLxzt6KeZ3DHnu
s2IzYlZiuKxmKE33Dj7Xl+ddUzPd3IFQ/FLbb3sBzWil6B0JzE6NUlbKtKb5+VgU
dw8Ok4KMW73opbzCC/4ax6ZNvAJwaADjsK9cUmEwRU3WQk/uePa+y6XyHUF2wVnX
KuaLkF35wZvhCSZUMD5ZtLyOJ4Ko0xGQZSANIJ0mkif8Lj+drnabE75/ywmpsLiy
7JX7U1JvBOckrMWhXwgq56KWzSLLwl+W2OsLhOj3hpNNsxb7QfmmfrJqrDmUSx2o
ZFlh2mXQIs61oNRFryhlr+CCYnGQnKPcYSvrw+MiAzdkv0hXrOcAJR3NxVV8oz8m
xvoufvqiveGs98nXAHtO45LqjTklGGvlCVosYnG6mJi/WZrF/E1W2GQ1h3c3j7bI
S/bZGmFKkAsJr3KpPpGCWU56fIQQCr7bcAb7//LMTJ48TZHUTeAm0lpjL3mX3nAT
1ob1JVhranTUkdfIRjpErdIVWDxRGZbdhet5KgSCXKGnHVeb4lWcdSPPkEToJzX+
vqy0YsL07Rv+4yrvGdLHnqezunXg7hDScC5r1YH5c92AleHQ3FvNg8zgIuuP5jg/
gQwUt1Cu3CBRhXzg1H/SvflqqTO+ctpewDo99YnKOTyi+Cq6oS8mPiRtQhbvTbWb
zBclxAevFDYzXfJavNkBtJFhKXCwK2brZBOSoe+UhegdYFgeKzJNUqTCRTbUq+MO
+crcBLdG4wdx+sANhNTOF91OfbbGXd/aR0XKDy5vz4FTDCjUZ0dJuJfGsKtJ/ZCC
Htb4ZLV6YRiy7TFBcBBtgp9tGQhzEtnC8G0KWkbQGuncNlVRXhe/leadOjelG/NZ
mb7njSv/pBRl9fZiG+M4GdoqNpygRT3kLfyB+1tfLwLitKnNwHlpos+6hWfNzHuL
2v3BOFvQPaYH0Qwl53HbhKjtSGOt8/WzDbmtYhDZSst4GBLcR50dQMXkrn9d3o09
UK17y4lqBaKmNHSLtLQJZK5wUf7xgXoGwvpp67ob8ydNPaCO3N90I8vjT79JJb9x
FgOJnzqDV7/j5tuoeCngMszNcxIMhH3YXV2divLlAbXxkaZmwDKsH4qTccotx8LA
K2Hnwxq7oh5bpEm2Sgo7t8Xzih4uZ7s4xbkeeCmFM74AA8jc7gyBtLXSsubzXjRI
+Xtr5Rk5PwJRpi58CAfAhoprRQg42+NNmsHTFUv91wFmhntdcSLm+8Kq8EdXOC+J
ElD7jM23cySwkoo+dhdYo1cYJwnk9w4hqVMT1FdopVI1rceQqYfmbQg+gEVi9xN+
03TnTCLzd7B7QYjL/OnfjhqYL2BHl6mcosm0QpIVoTE13WZFVSI+N9KmQJjIlMpT
YVgRQ9ZBstgTyGh+LXsV4COgm1Ybt1YqM5HkEOZ0Wdb/st9xdvVhzL+r48Me7UUb
yea7EwAngt8tEymgWiqg5jvbio/O1skUaQeQBDCD/v/TzCb8b4sCSvSWkPfqmU8P
S5go5EcjSNw0piyb3HI/oHteYiH6DDyWO5nvp5IZP/itAxN/yjKUDxeQ+JsNKJMG
U7mP1cn9jTVGmqOfNQMEG7ePbM7QKTITpv36y1zWB332kBMOD4AHvzn9mDgZ3PgW
RnI90kWNFGfq25CPeu3MRuYJjFmAyDRn4bWaoUYCsQCR9E20O+RydG0kqTao6XSW
pfa9Ou1G2qOygaZepE9ZUqlsGCZwl2CE4yIn6wqyCfxJWrGMeZ6+ULfribTH3bHe
StvO8jU5gc43h0qQf+Fxqx3kFO1b5U+drbz3c29DDxmZ4OPVRffdfVBSgWty+fr8
JdUU9JDc5L9rGAeJjufsQUoxLqWcwemW3PbdLzSzEK+yq7PuW6Kz7a3BX3FHa2wC
qu4xHM9ZnRlz5DT/y+5bXyqMdGBeV4bQog79XSobKANQKzzEFx+LW+mlXMDIp5+t
jC1A8yeIeRVderC20JNQ4t0HSyRZmrpmummMGajvC2AvxAp8wJNdn8zpW28xT529
xjuC5jvlgSEALbVIvKct2fQRtfA1ycCtY+IeLbOOj+gEWhhwTY2wwLKWPJFuIWIi
cgPSDRq7qbta81lg1zkMumj1DWP6Kl8LGN+GZdv1LCMvhSNUcS/5HyAMMCl0iUY6
Uk7crL2KQxbqyC49MTPR5yU3ohC6yLPVhmr7wi+VJN9Dmv7Eh9Yd7FrEGx4FVJwG
ADTRNjdZrwmnKm+RVI+Oc9mQ4bbhhhkNb1DRSKUuL/jDsIoFgMpWCfdT0jo5K6JY
xpONB+fah77H+6EXF1YdfhiRhJqiZHXyBH27c7NPewyrRqUyx/CgnlKxaYULadLv
X0xr1x+4NVt+wXGjdvF95ZWJbMmY+pWb0/AfUub46X0xYHzcJ/LeZ1HX69+L6Ev6
YYYHvZsK+6qYo5KfEyJIZW4YPaY0VhAWUYv5wTcNXYPonio4ffic5WEpmsuy+efg
CjwIwzl/p+NsYscmsWv26xe5XOQdZ0dFvhP2CFGDWbn2HRUq6oYkTkvePrumUzkm
fO5UEWFXEC54wS3Cb6sBrpcQCW4lae3iEmSyeQRulQH15wrpvCkt1tkRFLSEFHxS
sE645uoYV2J36MesFioSZoIxlsKvP6i2RbmOzI9mf8r9DYr5aO83aSEAn5QQjZ6j
PXdfLT/GaMAduxwYkQvYtrB1cpSMeUJaUYnAtbbKk08xt1F5xjpk/c9tYdbOgdfn
8p822E66nAJpYQQE/cmFhiJWbGrtSWutY3aKwOzkC4PSj5lD04vX87UvPYnHvS3j
blADAb2zlWuKkHc8wzakiJ3dxdzBl+jGvvQEaLNnpZ1iEq9GRTK5/ka5KZxt/nr2
i9QJautSgCbhA2q9FftCOVLirRrSf5h0uzhtyhe3fbpv3swhlPpp0BnbMb2YkIFW
OiYWNzlv6x4mP9oRki5gohWOi25LLqxxg5b9Eb/DGp4tKGOGRL5f+Ds6JE3yqAMB
7dl7dO37qz04z/a3MfDn1AGR/5EJEXhq1EUZeD2cB+L7EqnKrAp/cjzaEa18dXf8
qtnESM0eK3f/uDyD88T3yshrhVm+YQEzAvj2Dy/FeVGq2Jkk7RpBiwZZBAdJxJrp
5u1a2MnPDKdQHwZ6NXdczgrXDCXAT2p2U8fMJq6Udm20R+Z7bEtFqQCKaRDw8IRV
l8eSlxZ5UI856oC9yfqokudjlIfNIu2Jg46rnodh5SjhT976+cj8JDmxSHw5370H
pMD0hIKv5tg+IwAiiwO4X4jNzdOpQrjuXuM8qsA6JIdS3x3ds1YROBb+QXnf28Q9
vtBi458+eBQOcLA8Agusv0KerFUfyYHwdAFCfb2OVJ/Stu5552LIQqzpKk3kPOUn
w8nmSclE6mLnTPiNQqd9OxBYrQxBF9kXI7aqTE+cg9joEbK5I6wenSI30+gAbHjm
tb3tB4b0tYNL8oTidY3vV7CgAdRI8fMBBxm56prxRrj/BsGJkkR/usvQpHd6HmB8
bbTR9WDGjuSZgYw8oj7x2SP+I/lVU9Q/363jEYRA+O6AhnYxs3t9aw7Oa0bQgOJd
5yySrcD3m5BTy26iSZ3hVbIr2W8e4sVjANP7K+c+kDiw1zFadJZTiqd73zCtZpue
nFCY6UIS65SByQWb7/jVpZ3F13y1vi95mc+HkoJNUwbKOVVmEm/1NPYzyrUahUOS
yQP6Z/NcKPyZQ7qebbhWA2dxHEMDGNDqTCa4y/VKHTIAqH7589XCKSc70H4y7I4v
WQmgVhvgFd+ZKAB4awCwisG+Y0ipFfGB2yv0b/mV0xDhvqYq8BoHFSABTOy7hBKi
aBLtmubCs0ByQA3suej7APubK3mwRMw0vfrmm8Np+OnKMU7hgFPukESdFHWxhKPz
ijGhJL1CwCPWRTEBGAG3Dg0dJE5wEvRdTq+obY/1b/KMio6iZqmPLCnwIu2DuwYy
FNxp/gIm/DmVRrZ9hChEi5CwbfNeRe5s2NegNFulNt3TH0VJ6ZtsshkN9ZtZYs9P
P+0oKGTtC9rz2wN60V/vEu6aFfh9i96k/2QlHxC1A+F1Kh9zQUj6hI50D+F8UOnQ
KeJfIVgdUrwbzWHpwr/2hkEdLw/pWn++wB9DtayjjLZPCOG8YA1Gg6bPC375+4Pa
HpDIIiwp9rbDz4N976h32UOgNXavfbV72BTNhGtiyM3VsCacdfaHqoTR+LLayTdr
kWIB3WD1yJr43Jd8hqTYLApGCU/HKYIHzgaJQUFGLU0hOHJCBbQHpMUAyKVSyby3
db2OF9zAXKre8BwIHgKOw6M/cu+GIqF/OzGeVp/lOSIO8g2WI69zKqE9OwedYJ9a
kSsGr4/szxsJgKCIGxPaTOC10sC7fUk7HPEsLIebUI6kzF8EH1b0X64/MMDR958R
Utm6E8WWcSp5HOmP6CmHRgkPAI4FS6sDWdg2TN6pva0eDwPpUV5AGG33pb4/M7YO
VM0ARHor1iE5pLAp2BB9c2Gxmm6IyefvQGG5bxAjmJf7tjFYWuVMo27Cw5S1p91B
dFvAGOunf1tJf0F6tn/8CKnKutYS52ShuxXkXDN1xZb5nAwc6F8v+HAV1erGlPhm
Fs4FNJd8KiMTUuK4NyTq0TCjfBCsqHfD5JmpItTZDnv2zRHUSi/WaqpdUnhEMpx8
QqTBYro4DUykNWxw2xO1vieQeoyZ7ffFmdHYaRFnnZng2Bko3yurHGAgw3R+jtcH
OWEIEFOjJPMz2W8mjPGBSxAg3YLaocPezmrBPJynOmHMYgZWsE8PEquakEsuxp7V
e1ED0MNCB5J0YbZlhSS1g1qWaU7suxkbgZMuwmnctnCfmmiqy5KWArs5BXgEdj1d
+pZVBTeBDxBwDkmcEgv1ZCpm0ddo7/2jomw9GKdla+GnHIOeHwW0v5eTQNpi97Q7
JVIyzw7sN1KcZ5z4Y/7R5pmtOpUlJN6ZP/9vDyXBzqb72Lqvj+K0+zdzG5srZUcC
VRAogeQpWk90Nn+RX0v3JyR8M8ygL7rHSBCtukB48eBdbCmqHB9hzQ6MXw4fHzKY
O3Tzwfa8fBuYpHkncVTMbPMwwposOr0G9mDG2hZGCPS2Ro1K4zphDIm45FgMIE0C
UiYPH2xGDPWokFNfKiYLh7nPjut5mzNg/6oM6JJTXxOvbL+7T2Ze/R/VGKP28MNq
Sg5k6nnQ8xEPwY0+NLNihT3xPJe9LAoJ1ZPsixJI63zALp1BsQthxQpt4PQD9nro
ECIsVSesKSSdAf9fZrcGexyL80Mara94QWFMb/j5zKpVLCsgf+K2RGf0mIQKkVad
3os/at4V6aoFJ/Sr8gsI/oIydMF+hG9LN/L9INmLWQhpmp5wS+II2IOM3uivqaeJ
TTMkGLIP/kS5w+6hkZ8MTx+acM+MZQiA2GwNNAwDV9NvVRfi6gQdXh7UdgAkTM4U
RD5dwuIsZu5hbA3joJQfl32g99w+bdRfRmEr1TLqMTH88F1YpXa5B21aRHVzl9Cc
4EiiQybmEtaR+BZ6OB4OVL1d+X6akjL3dAw0KV5/xVaga16HSH1xVMXMYxii5R9Z
ufRORiUZizn1qoABy2l/qkUhpavGlu3g2SyqFn73msqqTYfx0Q1+KdpFRFK5fLRw
jI3Ie49qaHuGfXKmM8cooWsry/5El9fFJX5vFP89+989WtpnBhJqdx8kzO/SmeJP
ZB4sz/sEo8noH2V7kk2ptFYUWIaJ0zWVYV0w5kDQMAbSq6p3yF4csCaZoeVFUzPm
jt2BPpKospliJ1hEbFFENfdXZ2pRzGBqCZ1FmCGgJumzbpgMbB0my2UVKPildd6S
TDU0lSJPdqkj/V6amw3dXAyWxpK2ZWhGZ5G4HEAmHig6/IHrq6dXmi55ZCLb42Ja
MC4cjUO5SBcWfFKNVZUaxkzYKUxsFr/UKVPhLxmW7kOUvsqCionQmiecmimfaW/l
HiBlIlEu12XnC4H0im70JhTR/zOj0oLnbxeNacZHfXI2UT82/0I23/0JziEGF6lB
PzMSNR8mMwjuc6/BEt80uijgY5UbTBDr+1/Xn+5D685vxvDj8BgjsogHWhuZErKm
h1Dn/8PYCmLEFhOnJlp/XfVUJELdaXQ/32l/b5Z361O8sDh3ecI1LaWelfa85PNy
WjLTEiero8wPHfEHCmwiKGuKfyR1BHqcvi+SK4/4WK+SKrnHbtWATTX0DTLHx/4d
NSKPlZvp+Q14h8qWeOSgI3/zoDTnIWMPFA0TS400ZfjuXDSGhg5TSu8NETlEfOx/
Wi2uWlieEY94wtch9JsHh2s0+QSI+d/PZV8Q8Hjv3ntF0NvulULsTtC3JFXgos03
94xxvJZeGImO/Gr3ixSUcEorq0TtFoqqONFRWwpWJ3lFBTJ7p28R1FKmJODqmkbQ
aoiplz0Hha6ZoY9hqEMbaYcVRIn6g5nDejnBgbrusiiQodL1jhbB3XLxBYZhW+M5
quYoN1Np4I9VSbw73DD7xyWbIl38eMShl/GLyx/LyT5c7PKBWSXRauVTPe1itTYX
1es93NwA6Z4cMSPfgCpaj6k2RZNepoo0wgd1DqNyWXm3VDWdsf+KYSX04OWq8z2M
5gleqdOTPdP+6uXG/UDzdmyl8qfE/hstBcYSOel8zgyqtgBgb8otFN2nyd7noEH/
ln9G/Wll1+Pyroyld4MHBwj2wgBTuN9bX0OSjctO+DQoTYOshXUw8srMWpcOf0zK
7SfjSdRTnbtoQdTk3aKIXaDehtHNARNvU0SzMmNfQYQsqEDgNXvSDZ6dbgDAfoTD
6GR/4/qjfRFgXXO5928TgyxKfyktU5+lvYdVaKx9snYP8TFMLm36KYcrhySgkvEP
s8tHtZ4MygJJaAI0HHTE4AKC0qmbE9DlffigzUsyzftMfJ5z79NGqpzvrLM6wyzr
O3R43XeyX627oOtluuTQbRIP2Y097POqYqKjfZnfEPRk1gO/MCW8sMEgnHbjBMFg
tyJXgdXrlMJqYRj4caNJBMvDPlIPvT62/eaLm7ps2a+v0T6PYXwXPoafohAus/kc
fAHznl7CDtfhXv5h+KoeT2Y2K9f+vV810fy84cqAR3p88ICHnAQqh3w2iFS+wB8z
LY75af5W+xx579/dghvAwHTlWNxxQHoMMcqKtp9TIWiL9wOUZsrxQ1aBlRsGeP6e
BscJJ7aKgqDalbnvmrPkd5fu3+4wGahX0dQ1djYkMQeiRHaWjUuAFLDUYkByzHkK
4m5YkfEjeImxue/CPxVedfUQVuJNiCIojBtBuMY1PFk9OhGS5F4l1tCZaDXQhXxQ
H4lcfkrKW1EianLGdJxysqFirW4AweExKE/HSp1gfGvVcvqWoBPfSncebc6SkYyW
jPjTuGkwtlLMx4z9VI6mlu7s9oUe9gxouDELLIsFX+laBDrZ/mSJtcPNP9gfaj1h
0syIfkj6flp7XydF7ZsLPZD90NRkJKJvrx6cmLkaD5fzBGdpV4K5XKyN5BEeUses
5RgWJ8Jggar4ZcqGnb6QStZZDgKI75N4kKf1nT0TxnZeV2dhFh6i+IfMVQ0dbqm0
D5koNBVJ4iu7kWVgwBRN2TwJgPdKMeo/qjMjMI+pounK62XZ69m+5fcJRyYzBlks
6iT016z2SOo8LdLZpt93PsonLTZ2vgi6pbZxjz6aKLjAr2w7WfKKXtRrp3+2qqJM
+DdfQUtZMtnX4sDEL1gzws7QoTHYcoxraDXFt5S7GsiihSF6ioPUvvNFCBogj+gX
xeQ+LTXHcAaankdv6WxuOXOnIniWQbVu71moRrKoObLeScskMalB+iKqWKdtGAG0
YnU5ff84Q18cGvGUjaNfof6RYGyNd+O8M99FiGsOOM36voT/zZpokbpYjI9ydRJj
j4RZr+HtGz04OHufrNybfvUjqIRpJ85W8UIwH+MQxGwNiJesSdvKiLJb0Vo9xqGo
sm1dUaOf0oK7/ZFEoLnGTlf7xLe8jZZuOMNslKiWo/7bykYX3eVwlHIHvS1C+kLO
rsgpvRMzHj9kEBprOiH5kBbC2KyG7gMD6bJ50MaqaHwpF9hx6N1c+a5weAGVJQVc
RxOe+oxYuyi1Ihq8O46r2IA6YsqdfIs+8JYUe7XG2MS9lGyitAE7NTxQB4TPaxcY
5ONlsXIlfPVJ96zyaBbErNJHWSqGcqt4HyZpyKcFnZkh86yxc4AZMYrCJvXpjLdK
lhXpi0pJNKenCi7NvGmO2OTa54H77Y+k9OvPr7AfuBE5Rck5S/f/BJdWEyiAEFOx
nZgNABLvmSF2mPuP5jQqDUP7PKnYkgbIQankJVAcTkQzWK3lZu5NrPnR0GpMVz7A
LQf3vWLt6re1ihZbJgdQW3nnkO4AkMmHgytOSKyWMXDOANWxLxsNHK5tbSukFUJB
14Qn1IsYtKGO8FfW0p6JtneaYo9QNTqrpgzFajd8Dqmqnhi3TgHjBiUUqw78pwV8
dNRTJYBJbWsMchq6xd0mqAehfpIVlQFMMOQm8M87Wf0N8isntevhhm4wcOA0vka0
89+4pwB2cW7w7rTB6Adxf9/AKvorVfUHRn3tFdcutuqbG9736TY4v803nFHguXcw
6hcpY13DHsaZLXc85XzoDGA/4YW5LHltK8uknX5sxwN6xaMWjkQ+7QVze5nemi8a
85Tl7OAbP5p6jMKigA1BLx5tjSOk9vN6DV+hyqzXdBik3EgF+/ZocWGZQTaoidjF
cQu6eEoYdVteXF5KGvjZgAPWeVYS0ltUyFRag/daDpIdGKo43ggMH+jMQjqGJpfp
ytjpyA0kRuv9AvIQD1SlPGaDtP/KvS78x9tmAk43r1kPN8B7EflnQLULSRfRiPla
iBXV52ET2YysDzsjhrsi+UhtQ0jMJ3xQVNf4cg8HNOejM+JlU2nM9wzd1yryidIh
3RylT7a3wF7PZ/BWqbfemNP9/ZH/oOS2gEjShjSZl4pNlB8QKaIqRyLMwuGlHcOL
D3XZKTUMoLblgY2EopkxlZu2WISialR/nGv9vF3zCv86zAZsaihPf7UnxG5QGNar
dzzGHfUUE6FO7zVWKlw2zu7ZUau7TIZ9jE+/3ZMlnuX1MCi9j5hsl/lknROhehie
uJr5Fs2pa1AJ3g5z8Q29BMzUqC+YMJA4EvlhQv+mTyLPRf1UYhuNN7pMIhtYXM11
lEgh0Fd8Pfi7+wmsI3iOIUheJ5UzRF5x4ICkw91SXJskI/djFr0HuSQQejrTolPA
5gbmbcE/hTkDSIJF6kd6jTwmQ85wVk/6Mdlei2fI8tZ+QMthf8SAnJSDK8Mvw0jo
/BzqV70OPA6VfqqAe4xhI0rJrjHsGY3eNpONIaFqSRCwYzNgGeUji/3VYacfY55K
YPKomz6TPTOfESYydBlH2pklqNhG9Sem8+TtY9wM4ofjc7O36SIwprXnwZtDfSTK
YLKYwX4UmLoGvBWGBikQ34ls5Fip2epUApeBdhgKI0WZITs/Ev2KW1KXLnRZ/TRZ
e3j+k/+AhRviWm7Duyj75WdPHZ6DwvDGrmBLy6MHCG0fOF0IHFBvhsxit2GbXouN
6rG0CLHxVLRgzTmypSdD218Ab0aYNixc1yTxEAkXLHUNJGBwOPaTcqPUIdK1si7+
d6V0PKttntu9mFnL/kBB8WNxGtzJE+PKyeNEAtYjf7UuuTx4AmNPWTI4Zy/5gisr
qp6uzEFZXfnRdemP33vH32FW9gWf3/eb/4NiWxwHv9e5vtzJ6I4TSzP+yXtuz/hl
/SvlLEhDwfGB7kXtcHphGF6rgR/O5938BD1Z4PrhsKAdP7bVqw2lZVM2jZVeAdHP
6U1QdHrEZ2w1nLGEgbaPgFnxgy/cytWKXaElUlI28j9kmHr363oxpnx0TktwA4dR
3CS6NJ0SZZ2Pg7/NsCY5eWVa9+mIrodfcaGQHzjUx8LLIqefoqiOqIMeQ8fZPtXL
rYLsFS6KJlU9P/VMzQvFqZYSqAB1EUBfsGo6P0xL7IPnhLcySn4kyKyOvHNpG4WW
YUCBqDeMiSMGsTPzK5sZ6zM/VabiuMLFCHQ5uamjVarbN9BmDpyhQDxQhxoddeG5
JisOKmPCp5vO6OaQF+j+TLB2JT9ejt/jSj+msSkXMqZjoOPvmTlz1+ITpCI0fmWa
W2E6YEKhidZLrI2hcrAiKcZmTXPbBpuvXgdjb6leF7yZjLq6L2/I9u0q0V08U4bs
gOkaMqwwiG/aPXvqwpQZ2zGNm7GoCwL/ZgKakOMXQjo8HDlUH+ZdGIgngTk2+vrJ
W1Zv4TRXNLuswRh8mrT4qiUbMKZFpZ4JwSa0UN5jMJ9OXM5Pcxb1wY3jG0eJXyXU
7qfCwadfNP6YW+CF2n9hn3cANbhF1Nu+a0YMSYjdE/AutX2WJ/XwFU7KpHc1/gDE
f1wbIllF6E5h01JNs7+25yGDbHbIMHwvcBhKU95+3Nl1QfubR+42B5dH3BNcA0fi
nHCp4+DkaKKUBWtp8y8s7t0/cYnyx2fQpxiQeOgTgM3SXxPIRViKMpAJ8r2vnNiE
UbRkRJajYzRGdxd2rH8HlsmXvRQdK/qrmcfqpDB8GxkJ4pD5hRWuf7AlpN1EiD78
nxvgTvshv2NE0i8JuXSn+UDcWbzmiK5yEu5BdkOC7pqvDBfLPXVNH04Lciyx5tz3
7TAPEF9eIWvdqv6kf5W8KK5ywl4Z+uO+wHqT0gDU2hIeDlKUHeItKWAhH0fA5nCH
+rswofivkgkyC8ji9dTlrLyuyp5eAYtW1nspNo7dJZIi9s6XzFKh2oGbhuhCr6h4
8TdIt3t9agHgeBVYSwG9UF91+6/tvP25geq15diUYnN9zag8kaK5UNF5dC3uYSGv
7eVKLtRhsZc2Pk0qrKDdsMu8PcwNH9kXyq7F9OF+c9mAu5KjLXMYrSYmMZ7UA7W2
hHdCZaUcS+5AMpS55AUy6Ol1vuYR9ehWW7rUCubQde9Gx1+e9heIjCXtYg6HuYPU
UvJBnIRm0Ey9IOjIfn7HjcwHKA7+lynDYf6yelOM9iOlgMvfOrL4a4jq10sH86g7
4q77kLRjqkk5K9KxQh8jkBV3fsTh01Ofm3YZAqqtPD5c8ksPNLVzzvadbQCideZN
f8SrN6wgpdEbVtWGkdSjCwFI0e8c4Q/J7ykqlbhTUqAWqzwgNhdjaowlxbhllMvl
jdLFPUfhn+SmnvH4ErJCsodv5WvPN/WKU7BbkO+W9dqJnh/DmxBSns9l/S2AaMja
xubx2bqugHs+AlC99kGWonUWnkCdTpJE8SL4oZsJfIyAzpS2Jk++wX+ODIqbW/dn
pHM9sjQ7udJXEi5pjcjGtEfFD2AD48SrXZY2UnU6tMgQMskdldCyFrmgOk+cVeeR
9tKTAWhayTpexeSB5VpEhn6lKM5TcDOgCry6/DgpF9iTbZqkITrUATbuLls+GenX
32NGa0SNGmzkS5PpPJQ8ZE6dJUcEH49JG4zXNXS36xAmJWWS/KNfxWkgZ48YXQKT
/DHhw7bRSPlk6wURGYRsHouvkn+igl+R2JvyJ17y2Y1d9VZkHp5Xg3gFnjcn7oT+
mmbIdhhj5WThHWI7SPUAS/ShgkhdI6F51DQLgCkSBepytH/jUdrKFkaTCZQMm5J9
UyKDzbxNTeS81UJTTriZzahWuJdaW4zbvYwwb983s41/d6jxzIh0Renfly+huHQF
SY56yt5ufn7LdzFqHIavUXDYm/4GGpIHX5PIg6WDXuYO8O/RX8Z/rfG5ITb111iv
rdWOLEgFk+4imxEv7htrdgmuJje5LgH1tvr8qkELnJmNc4sQlw0vPpeKYr3A5Qpd
tlXjrwXFxaap5cu0gqKrDwvgN4l8um/FqSBBjbm4uhO7Zv78d4uyfwSea/qtyuch
x4UJKihD4AJ3NCdgwpdkC+0v3bgecDWmBsiQ8wPZJG53khx09oyruScyvK446sIc
+pJywI1yS9zsXdUsOR9x1mKf4NmqJur7GTfzz2zpco1Dvm2VLnOfebsQSzBMlbjk
B5hAZowNaAGAZFWmLDN33V+Vgvyx9mSJ+rHps59IcP+NCc7MNjgOdBl9hxPm4tig
fm1/a7YHjmoA0zGNHv1dg6cm6xqbl959wk6V19fs8Y+ZSXBBJ7WByWsrJxIv0cYZ
+U/OjIcxEKr09ufCRXgioNBWOoQ14sdQcMWJM+1ImK4lxhX42D5kJ3HaD1KWoHZX
BTI/fu9LTQj9+F9emLy54FsKPqQwZrqzV1An1171iGfmtSTtx2q0kdWS8rQdr2si
aETB+Gi4hvzpuesMiQsSqpKmAyRFoYXiouaQEJp0GbB5RDfz5hURsQZQ4sruX1r1
WK3thFbgWsdkoyYErP0kty1ITQ/83vKWMSBAPh08NtpTqKxe/cPzSYLRcfcxMfxS
OYwH0MtaijGo987m2NMBvshCXmws0FK9PvHH1SiWvEgIbQYum6573C5m7s4eJFFU
CcjLJls+h9NPdFad3qXX1KcRRM+sfU4PfeuHTZxRVu0BW+UXh0baebMsxsEGad8d
ftxdxO0stZBh2ZEroNA0lGi8VhpMV64/SDRS8SpPrtX5Uls44e4ZpO24iae5G/7x
y+l06MYjuSpWH7D0MclTNevLTVj402nEpov2QjYD5XVpg2vJhodlsPXqVneSUSzi
+cw4J1DVgf5AwuQjgyKPFOARZNcHXAkjjWMrMrqYqryCCzpzy4MHyyyVIAJlDB1Y
CqWXXTLkOfAALCT0yF1CEfv3hpEp1E/KNgi9ECFd+IdIhVhzY75Y6wzbbGlaHO18
WKIwSdqb8x7yfLATWlbjo7wQ7qoya+Zk0NLQqYSbtOVFRbZbETqRr8liS6LBbwLv
PD0ljTwn4mXjiRYqddES7e/mDRGZacyVXgTw6r9UWSSxeLRaNOiFezB8VcHr/DBr
XfkVhE2cvsadu6e0h0SV3HSnhzRoYsq2TgTVJpV7M89ZIGcaeEMc77Pz4wZO1nUf
pYt/nXSuJ5r63D1P+QIryqXODf8J7lWbTHH3fv/NiDHq8nX9LjJ+tCsXKG2N9lnM
iS7BxGz2M8ZFPA14SmHAlKAZmnPL/PI9kZOW1pb7wyJCyyHQsk05dd9GxnDoav6s
HwBAERRHoCZF2S+hg9ngoOcFRF+e1hsi6Eb3AaNe1DPo2u+zkfIwElJGqOMeudLh
jeDlq1Qi3z9Jaq9wcTdDezwY9RGs5zLhKYMmRF/yBEJNWw4EXTsYOiythokx+814
0GIAmArXzbtlH5p95ENkFUiOrz0UM2ZxnA7CrTewzms6PH+J2SuB+CcOO+5VMYii
Kx2j1htguZLaLZoDUa6BkJIL5XssDqpng60PrJFAXwnPtTBTUuUU+G8jtFUxz3BY
7TTWcXE0UxBzmpIKw1aflZSf6HPCrZCV+kRsb0/B8YipRPiTKV8p6fcbpD1naiFC
JT1R+swR5WNtX5eb6VXEwOobUBQSf8/+FMduuuaWXZde9snzx+Mgb8LSf6jnoiLI
j+ZGYWVvaQwMwMCJf7QhMFhT42bhsVOa83oMxbb/G0I1aV9aMgA62gi1cUjDaX1I
ZYWr8U+/35m55pNN5DkDzt44yzXQb/3sjVS9Jwids7qSebUFS/amiGh85xYpW5wZ
VvFJr9YeCAHiN9OnYUgfufW5vjFdekZHdnO9LKw11ivuFEogce11zYUGMf59KctV
xPbOThHZMLmOkLGlWRuiJxb/YICcAyvFM3NzU3IIVlZdrAAXt71fiaSIRHoLjHn8
vHSM/sCWiTBYNtn8UF+atKkJZBp8vgNFTTaeDhrK1OUswSZmkUQb5Ydd6Ka9Tqxf
f+kBTzVt10pVrXkoyDB5KokTifarMSqKrgKHzsynz8EXTKWqxDa/ahLC4GcyonkR
ewU2t0VCJGeT4NcdtqukfaLlX7CHhFOJoEZytykNNx36Tw6fWljxNwcyGWiO4KrJ
7F6e1+vIJyEsTZoymWJ83PzRVnWHb8AHBGqRAPrKSYEBqoiYHcNhiyIvP+574kVm
9l0RXDIjL/dMd5enJp259UGquNaXPjzKMGMgCJpANGmFeHsnv+gx/1GrdvJlwj2/
trs0gAQsILCfKkVPCAeVXEaBs58YSiVksYeRu14GUMGjcGjkDXjlS9dUS3f5I1Is
HZC0ejhkfcYm2Xd6WdOPHU4vzjPRLEDyP/IwP2CcN9BboYoPBYSJurb9KKCznJOM
BNNK+b1PB9rcGO7jLFTnpSlOrLTZc8EqUzSeFkd3LxZ3cP2ipZYaJwOm+rpTq85O
xQE129W9ornKMfGpo1W95JK/Kz3boKlxaENsRB5Orb7LaWpVmFXyfkGzLo6lmIxE
BoUYsKrXf6nCLyf2zWdx5I+A0iTx/f29XRZH4ey85wxhWImzI83D8yC3kUL9NdU/
e1iQRdcnZ4fjoa9/S87hEYEMh5pIc7BC5rKDZbR+weKV/fUAKIfxs2RPVY50ZK4s
RRS+g1veysPIgMwedsZs05hFew97vxvYb85K2fd6cQ/+3R4pT4zKRER/ZIAzJpkY
tv8Ae49383Vs0oz67j/B7q4joBXKwOj6wfCnbGyovY6WbWSJzx42DdJE1qHxae4P
xrOeOFj0s4mH34JNYAf3uAH+IMrMNkPrukkzJRR6rKLVEeV/Z6CLUZsAZweHfiiD
0cDxOtwnheHA4zBQt8ND63XhkPe7GaaC6rIjeMCDvt07vbB+FaLZsANEwpJ3Zc/c
G6Dp2DJHAdY04xoQ0j7ZQ2k3MX0RIJ4jGJ+J4aH/YnTCDerBzNMAB4qrRiiKYe2w
c/Qn6QeZZkAbZLpN1mw4C3A19xnMsNSadCpIPVsHPQimHDhNxPKnrsXrnjHrEsgZ
GDk8myXR3D1keCGlrG0qywwWz4f6DkLzVVs3Jbm+vJiSICTNk4Ph4djxKxvaePfb
lmeUClg9vyiLdHesrv8jbSa3uY9+hNtOzW/d5QT6tebXQD1J5lbMXQ3isOOAyFEi
HoC1+W9dkFeX4s7SgYMgWCLVMK84Rcuqgpy8Km739vmIDYZziEVbm8TSR2HWCCfu
P66zL17ZzhuhkdeKvTZDhnR+3xHknjs//c92VdOW8MsLLbzTMMTEc26btr8moK5S
Gbof7Nif4xTncq5lN4cAsS/1ShTd7y+Gmvbp2HAHFWPTZD9Bqire0zJf+xB7XjLH
d+R2fgqtwzynNKNZNIU3SyELmqWhUMw0Ym86nluuEyE1u24PF39NbLnzCdl994JR
obP89AlFem58filckQIOooK1X1V2iRttb2LxU+1qiXfSVdh+NDYBtMEvivRQWSPc
vcp8wNruaPSDBa+rB2F6KB1SEJI27F6zIFjlHSuEoHaDF9LE+Cl4zRbVREM/WRNg
TS+0yOJv0G929FawB/+pGo5TmLoEGL+BQkDVmfmulM8DJqv8ONtcRcklQHQJO2YJ
NDR5GZ9UpsVxar1D5ZmDcQNzCwDrr6BEFoAtFQRf9c1bDw3yytcHjynAhH3QFiPT
tgXI920FlGQUarWomo9zNdOspeXZE7MUqlpwvSZuo9e+w6HbsanPItrvc2zclTly
sJ06JhzVg6B4Jx/5c3DWyn3LwKQmuOWUgoizZuEodAEFi62JQBGzAzGy5BeleJff
SDCDinkKayjr9/9b5bHwM5Dd8J1Oirpox4RMiEjYSfsEZMCqDP7nawmlcHhJ0tus
koXE3o0P/lMLbD0gpKISuKfq2PvhA+wi6Ub1iMcV8iCGY8XbJqd30v+2WDK+cjvt
YYgHxeqBQlij/tIpmgfaLSGYEQFJQ1XcuNpCkGtEx3+dke/LEAxr6BhDgJBtKDr4
Pkcg60niZDzb5tJ+gHdtcWWTJivNVSlKCBr+FryZqA8IipQHOm6vIinhO342NrSS
qRBTrnLW8pr+yt5TWgKdWkUgjhu54m/6SugJUqGHu9aJleNqyxnMi/ZMfrhQX0jP
Kvu112I6aVEKWp2SgwB5jqt3zoDpFRaCSnQ70qS0BAWKkQVpOKsNOuhfnEwh3+Lj
HswUpC2hc3JEtL7+nX3Poi3JfJ93OnNSTILazOf/fr95zx8YVhUTrAZw9A4+4Z1o
5vVp5jbpyFfEzFbqH1paMh3BbH2aBu03ZsbRnFwzI/bwdv6Q63GDDIEjQDg6CKcS
GB+iHn21g5TMRRkChwNe7ly2d+WaXH2F/2o6a3gfAi7/XbGUT8cTKLfUBChq+OwY
E5nZ6IMDgJYiXWCtKm/WnVaUB4di9jgkQHuX7hD5h3xprzQoRDyv6PVsHTnUEmiO
d/qkc0jebqDnqH4/OKIw9H5W7n5YjSnnVlEFeM9rAXZbphRNtTul2lcQo0aZZjPR
JypXz+SQ5ean+PBtyxzzSbdlrA2nXMtGly26xLuKo0OWYDdzlReThw0ErCGX3cmB
6ToZVakIFPwzVjGinoLTRe/Ioo6rKa1sL7zFKopTdGxQAtLOb0tzZlPmDCCrWRow
sBfMw8uyHXOq/p92nqJ2OW7F8OV4LDucykw+vSJDK6CFAsb/t/+o9k6uU5PtmnUU
cjOOvvq+JLoZfOTfgeyD73mnxx/xd46RiBFEkkxe9RuFeIWRiEeHU9xcZlbRkAjc
Oy5XLXjXgl1dlvZMJiXN3v8ng3EgeHpNQ8VYT3VjJQ0xFhSMIVY+IGMOjxcLD8Lz
ArzFDtvgHM12xGhzcj81zq46GUWY60ftr1GQ4CnIB9OKkGwuWEqPjn+x16keCXiY
OiHiHslH95bhOg0wEQclo/jwkYmu+hC/2r4tUEEBwR/WjWHg3sCnNFjHVamEIVwA
/n+ppoiyQOifujngE1AW0PHgvw9EhrzV14LJ52ZlWSIcaqpPr+khxdL9f6Ze4fFL
GDE957ZkasVQASxKnYVBIzhkPLsNqvxGGbxVnRK/fl9li7JaALnik3aMkwtg7kN8
0lXkASxLUNLP5XA1CLh84s21Zfh1SoSXS3zlEf5UbzPWj/uur1v723JFMjxVNslh
Lt85ojGxqialBV1zSR1GKuLaUEfnFTI3igW84AJ4vU+Ono34PLxEtTegE5AeG45B
M07nUzqAdiu10dtmBZFNpk4ZVMFi5U+mjY8JXTPNAlk9YFaXoNwnNtYuAd2zgXwk
6oRgYjJy3U16Mvuo8k7/aEoTXIfH9kftP2Le8mpjvYMsZfcfc/CV5d54wnR8cZnw
g0OtwGPV/JEIoxdvQRdTDEJCqtInEarGqq+TBzWZoWSzhz7DK2nBGG6Q6p+2a6SU
Esilafq2eyDttVPrC9svpxwYuLELfuUxVLs3k/3udO2xPzrkoROhzDfX/1/JPjtp
HfMTFykQDmJAdfdNT18zL5Q8zdxQS7YBjLbVImma+Mo5JwvHH6a1Hn6ZMgRPgp4w
GC7myATZGH4cFQBc6q/7Tqp2Pt4xdT6WtW2+ThlqTp08O2nQ3XBq/+hRP4lY1oBA
4u5FY4ZzKBtYd0gCikQ8FJjQMTkq7TCoCb4OF9cExWPDVZ0jFJzZwTBSQczwNlqz
ufwp6NkfAcoSNZyowe06rkIMdR8+MzTcnYyqdrddqt8kmV1UV/v2O28YEMqGiKmm
Sczh+MbfaqZCM4N3JbdoyBGlZbOuYmRoZuzhkyTuN70r3lO+YEHRN47XdVs3d2T4
asbTtu/KhyDSyMb03VqeeEWLaSJaKqMN3urBm8SYa6GK20oyDtj0CJT8tIXTAhqx
UDjrnJ/gU/mfMMLJSvlcdN74uSEWGMZ4Dbn41J728ecd60uwhEsKub72UJ6ILxn4
+q+86BOGW3xMuMpFGOBCT2gVMuSYfEdtt9tG8cfrwVfEdXBKrFkxGwTN62EN915i
RLJaEjBWCjxu8L5PdNIlNlu73LczikAAhTmzZ6jNDpri/g1aawV0AIgyni22tLJ0
OnI83VwWxMpi0/55baRA/4af7zGCJCvpIapmsRxNVy8hpxKaGMaSn6KSlJxnlBJb
CXW4quV3qWQ3YPMtA8ODQ9EA84WIFetRLDeXV0LLJcKu7k0Lvowusmbx/wdNlXDD
zFPSpK1/+dm0TiGRE3+EdGYrq0mgYT3SuUtjuDNrYo3ME7yf4jAl8hRLwQ4ek1hG
KnCPKoo7IcGZRu7PI397UrEBptBlAhn6z2X6VUneI/dKtzmwKFliLGC+WQnsYab7
kF/r/Twh/PTBeop7g1IOepruq8f9EEX4uucy4BAz31RdMBnCa0FdLVrpb1fiL5te
jUd/ACHwt8ww9Pxf98vAiDxXhWEVKjHwEIBujaQHUI4pj6ddxrTjFjDycng/BdGO
Kca7NgQwSkO/NAbm+SnRJB0lMuz2Q+/GdpC6q/sYZy9cy9wYvfyqCCBlbhFP/4mT
kqFv23sTgWYKjw7p7Ux7p5r9yYp0bYXPTkmJYJbNMI4+xmB8zdX6q5zlLAOEIWKB
++adSV00kia9AcWNGgA2FlzL+2Ep+Mg1UM4akrxevV9sC3LYsna09cRyEXVvgRjB
KpiIGW9Fy+lMcpBBfVf2IipO/uYZEcoE4YmgXQoH6Xvl862mB4L67xCFIBW5Qscq
VDM0n6qMUaiSR8/1iLfMW9DMqkgUfAPzK5WA4GT32r4tB09cJesVeTE6dQaU6mkJ
SAS26U3Io758JzdvaEjsZYOaP8hTGnPdYprWDt9oIOvx5DCEoppwC5GYtFoz853+
91D3z+qjA2+kTKcyrzOmRoN7z5tknDjn2xgYyRwjdgMcjTRhZa1NKzCJCcLMWYXP
o5ItYOWctRNpTMCWrX6U3s/4SKI/eJCfq6hzoT/Kfk7xXcCrsb2xJSFy7U24yZlT
3cD8HryQ8Vf0OjSNGRbv76kHB0dwgeCdds0OIMv5QCE9Su9rB872FdeNhEPXJYD+
40zA5FMlpWLt/p5+s4/uOK3jKlMOdzKkCdNtff6uyqhPIg6N314he/OkeUEUOwVJ
7Xja6Wknne+h5EAnaCafO0H6mcfN9Ol9Yfd2PqeOS3QZvHCM2AQlu3PypqtiurkM
f2fT01fz/9WEMxNfS63ac6vOQ8lvsBDNI+TXYCmaftAvd5CS2a2lluB5Rx/cCmpL
Ha1VNr5ICL1Q5PzBg+VShzD8TqQvX3P4++qfbF5ZYbWeetMXOdrsXZyZzBLrkuti
vuYwYmjKgEVxIxZ2nqAD/nEKrLtCE7uVzYKSG2S8+3M4kjQ0HBGTRqZ+DsR7C1CK
nh+tk0omTv3osjBpwdTY+3DZ4IVqrE/UMR17uKU9WGLT6vx03JrGHUK7+vlD9zg3
+e03i5fjDoBBhRojg3IXoMw3GAEMhPMDtuz3uNb9JfYEDosKb73nJAYgo+iGddYJ
nl6qjkq8xwRxgHrCfqzUznx4326Ne/pON71XJshHi7rbFuJSMjk2C5HXWaSNNDV2
wBdy7zhGddgOwCAnwjhV+5TbOydImSalwB01UfiqSDQB7JsTJS2HHtLdHiRvaXsy
MTux4Lzx/kG/+O0jG0d6irxCISZsShIripyg5CqWxGp/PmNRrkxB0wF/NNyicaGB
wlmwnaLELPYkpqUpUul4n8v2XqDdMsgLEtGIEi04FpzR/QEHOMS9YRD/V1b9oOMy
/tV6vgr//AWBGF/2V9LMpkpEcznsq0WdLQ2i1ROPcanJFMl17DuCSxJEIYjvkcgB
k6PPAyenBarYTdYMnCth+9SYIdmugzMNZSOsn/tMzoAC6DZ1fyTzqdqTQ38kJg3Z
10wIYPilZo4+gwezpU7EZLbS2XRplFhaatJ7wZhZSpYClZJF/oc3ohnmZWGLOjQ9
pboWrAv8U/C6mbLMWOGs9TdxV78hlUOpWHdAz1lvQV6EP7Rte35LReAdgFyZuoQf
NT/zdfzTfkJzV2IVvhc24lvtjp1y+Nnz+pd9OyudlWyQUfeqr7Sbve7dDmkVUSmO
fqiFqUsquK6TqxdTuR7BQtkiXFepW1C78Xd2omWupFBWFZP/oXcWBqPS7p9omokC
y1lQYvgKQmT5D02F0LHkIiUAhSFKdRN/D/OWTafXhbhgADyLcIcngzxvjXWmFShF
prchEmSr1lqYveLHi94xTbdNQb5QSiS6JKS0X3HR93ijHG+OmZe56WlexGWdfSOG
H+4LCfvallgbfWbFtRCAPZhBetd5Bvc+NcEqnQPC+mdbNhgLf65UXHcvdiwonN/B
t3KKFC9+oVCFPvGtD+RouZKOI/eqzDQIfQUDuShNBWtk4ntpypzb15LgLTLHBRRU
/OV+GgUWWZNFi9XXcPhpscY10ug/J6YbL72DS/aqkdKZslxb+gFW/33y/+iSnHEq
zrPWiKjpqX457Rz4DpNx1beaFf5qGM5ONH8hGgF4RSjCH1xdXqAAZPEkPx3OhR2O
JdnEU8JqpwmStXVOwCFfMtxr0IETxFEmvWFFnif1Hzk1mGEzH43hAWn2zjX3cUii
E/f2/ZjgYgpgdE9w+V9qs9Hml4JlZWH+PnJ1MfX/oKVExxlR25/giknQJ/OZ8LtI
mcwbUw9IeVayFVaZS1lBcJGg2cFsoXhvZz0Vtw4paEy8ka5YibO9tbg5P1K7LXBG
kxI3U2BYTGlcqxxtBwdgwtBL7p/W1+t1ykRBIiOilCxVaACaOwOVLxi67+CAjTLn
r1BOQXnG2W64hucbZF0iVe+i0tT13nrUZBtchG1jjhw3C2GeyI4qjFdudYw6qTFr
9mVmfB12n2x/XT9GBtXdgTyRyTit9WYQb24Ah2ByqtpdEGSxRId14f+haAm8Lp2y
zlAj0j+O2v3w8KXVyWsZdwAiZI9rprmtHJ/tTCgIgo7VYKsaYTW906EIRjYG2IhG
NjHWfB79Ae1CATa2nHKkhxXc5vGfL6MUwH6vaVnCZbsqQzMm3ndR3FzXpOtjcuYm
BIAyw2VtJbzE5DYqQBbt5kG/J6E39JuTWpzqkAOwgE/28NRQt/U128s81ZrWuZwB
Cd8XCn4oAi9+orWAb8DSJb87iP9PkVod5ZUflwiSnOuqO5yrzC3HGI5RCZ7LRGsj
uZtXCEYuLIGzhy0f7rNGG7o5vcl6ReBFmKru9RR/yryLx2QRvmRptITLPWosALJM
GhhmIz/Et1EjRhvlr++ym7sASd6GQlldlfUB/tym+4JHWyvWslYlzRn5exmyoz8C
Got1+0Gu7TETzuI7xKgF4euwWeLk7udZoZuwpJYAA2lTJFXKa+X+X9Vz5CKCRu5r
+asIQjtzEq3IUgC8Hqy9n8Oj9uRqNVCaCeSM6xCMtWUt8qkkevW6MqKqDrAcbKp0
KvctSbMJSAOE2KOVFLCqdU6OEO2zhBVgN0ePSakLfbubhC6ux6PRVzKklV615RPa
MHZFE8ELy+/Oon7UCEuePV3JSIGm/ef4sqS8kwFViokdFbiN6G3uGu7rr+xqG3tL
IOORsIVeGJmHHm4BChJWM5jA2nfyj/srIz77i7Zb1ET+AUg1gIptlOcLdlil2624
wVzL7ctUO/mzCm0iVNGXAlwS75llHxpPikaPnf4BOJYcq+KdKj3oXscgJpjx7TyE
x+tjb1d6mxSoxUvUM3Jp+WvwYmtWtKypjEHkJIRrYH4VQZhDzUf+VUAs5eT6Ck0s
eCoq28/wlGmHEEba59EMoOcoCl/KKPlfJzFqzCq0CwD2wTPcgQ7yR2jPc4pwLi66
oaLXWTKyVdejavkKZN93cJQsjXLM8OMjOBhPX1o0L2gEcqNTTbEAonmqTWAfwSst
dnLbtCMuTmSnmwQR27p2Noe1hQjjAH2PieIn+ZDxNrlysK1DK40kJZon8598/CRi
APShnUn4Hcc/XNFKWVyPvJo0Jk+MhKiqvQw83m8yzWcCyGLzRi7ke8sTv+SzNyqq
KBSPc7xkU8PnkOT9i2LgwYpwKHSy5F2er4PiMOFsOxv3Xr8TdLjFyOR2vfI7Jj9H
eU9HmnmOLSv3u7W9HTW9DB5enNIE4SDwUDvBrPO4zIo40oHyIGgKC7OS08tiBJxC
fMmqgnEye0VZqECVskDTXUpa7+6ktGv5Ih/iVs6lAPrLMzYzTBbt7CJTsE1DCnPa
EduTR+U1niI2/WvrRsiwwcEB1XMI0sP64QtmXp3r4aW4zwWmR5Ll88m5sxqv0Fkt
K9Ui5vGXh3/CyHnCImUKc+3kJCI/Mp7ZAgq8WYTircLT01NSILrFgDd/ufpKVKwv
9cRMm4rlk+qmGPl69xp+8GQx/REqfB0NyyMJ4UGvsdxqOiY73CiIbajyYkib2W3t
vab/LLSmxRT4Wfc25rlTWRqthyJLx70GojLQCxZ8J9YMylxVytA/mFtPJYt4SlqA
14pzZUU8NJl1Rsdv2TNmmB8yMCgc+ha+pMFGZg6/jwkvZF5G0fNSq+3D7LRCvhyr
JlmM7LEA2c/SPAIjB3ptaQwZRGjgKZTW9YRrxtJWNKv86Lv+tlYVGHWaCswRZfbU
zZ3ENlBbUEJ8j3ts6AkSJ1uDHI+302FR6FRUi2DGV0i3DET1CCZH85J0ZNF6FJxn
ZlmTXkWdjy5gumdTtwl5tEpRsELLA7nO8b1KWtc9wIGQMZHu9tL9C703n8aKD8dB
RZJDW4i+EaBM6+GPZHLBxQIT7ZWUX9zDH5sY4VPRlvUORy/zsOroI5WG6nNY3k/w
7KTB3RA6sKLiFZCybf9ovzzJa3CVqPoPV4iS7jv/Jxm7fzfJ2QsXCMRrFpofNAtc
3BR6uKEjMnJcO/h2GfLkCB0wuKSVMEVFd92csnkvj/noR74aGG5W/nO0fx+krXXS
lQr0pceUwBX2yh0hNjqv8UCWLNGSha3oVa2+uJYLXIg2z+pe4KPZb9ZP2XnqO2aY
4pgANxy+tY5qekUoE/T5wv/QChgiYAU8yP3i5cm1hp57tTXeeSrvufeV0iwgErIc
3Jg4Hmh/xxs8u+ywgCkNfLZcXvH6XXT3Mh2cWM5YdL6wxQClrx/9ZMQXo6v7H1dF
rT0cYb2vNZ5tQG14EVjKVa27Ho3d6+edVo0ZgWjNExPZ+U/0vkvxyFIS0wDOk2mQ
EB6pbb/JlVCuii3/F7u6WUYRgRFMb+JcrxtzSbACCDGOrtUzZ58EgC893nSbAbuJ
yx5SL6m0bCaE9Ab1D9EVx/mNjMSQS+Pl+3rQAzkQatnipe58XAAsnbWJKHCOsJX/
6GdW+dNd8vbuN+7Q5k5lt8yX7ZIxpALJeHgNa6hJocpT6JOguVIcpf2gn5Yz5NSx
Jtmem29ehjqGHxezvuKUC/VPx9heowkvUDuLHs34MG4lihbgCcv0ZPSx/DiQCRh8
AASEfHFhSCheXwHbrJxlCQxXiguQ96BncafSnSzk1mRmZ42DGCVHYYRmrJ/fzGYy
2URJOj0iOvNjLa6pgJFlbdqeP/LrbipcG8hQG+0vdRYoHl82HzblcYJeN6fVk65b
xek9tO/+4UnYeroFEIZfIQ0Sk9LPyauXt3ygmf8Ir7yvQ5zaIjHRjOvgd++5S39Z
cdErf6mxkPAvVynhYhBeYU1bz64HBU5RILMNf4PbVeMvvfo3jWjLkvEdidX+SahD
d79tbTndEPciYzKp0x2JLWqO/c4gfkvCdnj1/kjcAwhqdBWMmwB8dT2jC0wUEXf6
1Z3NwDGzR2iKybherwkbH3D6C0oIw1xr5bioXvklUwdjpGgNDasIPRVadE19T9jT
iB4ZNJPQ85IishrBruZpSzZU49UlXg7ti+Q6s+6Rft0uXstWUJkqHSNrbcHobj+y
f9fTMoNJCoW7fSd3OoNRM8m6XaJr8l9mN9PAYuttQUCi/G6J0ZRGQB6Ah+48nNWw
Ue/yug6ZPDk3esS40Ly3q+TQS8wQWZbNEMSNNmMsCDGFEb3g49wIPDtxgaDM2Ahf
ANc79hjJE8esPnHhF1qszhbXfXMICIAYEN//VkbsrAaGhlE3bwlVI23mI2tQsdBt
QpOK5rrJr/8VKq98O/o3wVJVFbAQXVcefTgiHcfMGCx0VFOn5N0HGojCFFkpkAXG
yGxeemno8kL6Jgl2UpiGyeRGl9zQR15iSDVKzjTP9aSM6Jb2JHoOdXp2jKrtIizf
lzbTFsx7jO0IajDkVn0qT+uBH4yN5OwlCc584iiImkJ+Z11kbCPfMtrub7qZmzYX
WbuQzn66B/dVLdlzjJNVtw8YkCc2TyNnOuApSDtydO1rofjflP6vcJV6OMyFyY5D
WGsCRIGDbfdhsVTvnX4yvnBWla+4sZQikqXkj13iHnWXOynxPgO+VIcIzqq55QbB
ah6HGBFrKg3JLuEWQ5gCKkLsh32pRZ31ePqsgDEPmIBiwick5uZlttzqPjv5+QCL
IIHG8iEKrLHWWiVNqMDibwLO0SHREP3Zp7qnqihh6fqcKH1Om7QFRn9hzhhYxXrz
w3MShA/P6AvnQ4FsOKyLzlM2MwwLYW85IGD3MzFk/wy8m7ev7lNDUirU4PNKehwu
Nc3VkQo9uyyJgh5uC+Z4iIug+4ixAsNYDnj7lOHvmRvXl374dbU/MMNGeI0fzl/c
2WQCa0x4RLklPR8qA4GyHyQfYTRalE5lX42YcuE9fSqGqAnyCvr4AQKtSEcU6aNm
TwNkSjdp2A08+jApBLIkrqD1yLVQBrC0BG+e68WkOQxDr+HiTPyrjpkQrTlIcVMQ
g2k41InMIkxnQ+hI5ZMtfvN5IAcWLjsmDj2rJEKwv50y6uWySvOSodxUXnT/OtHY
ocVVdsWYPcysJkvZWkS5MEjzkFlAq7GZp2tjT7pBbi7PBATFd2y0fivnpkFit28b
sZgZs/LK22NkgvS6ErJPmrbVt6hvcE8WfCLArHE/D+kREUw21GIcOHBuq+Rw6sFz
AnNSGdZtO+hpTQl7IrrZWHzKczpxZqS9TexeavPZ2vyubcisUt9bbC5RB3kl1+KV
+nxFI8FdoksjnKNoKpZdrl0rJTNilF1B//TmyQ9T50tWArKSAm/AKKAEvScFuvtD
qpjGP9akJXgW6kS8ZDdEHJ2DJ0bJlxyAv6mISHRD+WNC/HZXSfzQQ+st6ST2VmSN
vFEaqPi8T4mes1IPGujBzj3tgtItzFH6KXuevAM36xWScPzU9e6hknfyU/EckH7q
c1/v1KNErMwf2og9UllJnwzJxBXsIOKU+VZP9SseG970ANML0wBsq9nJQW2Qaiw4
LEA50oH4joG13REhELEAh5Sdivdg1y81+0XnyOWo8agqwQLCDBcF03cGv2kjbec/
In9Q3AMOLO+Z0TTIaCzudwdp2MkSrZIRcCZ2YO+OVziW9JEnZWzaHH0VpVTMj1Us
GroFiNJMKFkd7o7YHaRxuN0OC+2dFUyXB7GUrZdKVYSrT3glkwncOnEWOVgmj1C1
2TXR5r6fFgs/iv96HkWW7SRSu1ODTCmXzoUNV1yXlC8KdPl7KCCD5Fw8WwrRiuHb
ybZPU6wzMAfnF21D/AKX23bHZeGQXCGCgy93i4oH3EmiCiKQb8QrdM6WXOtBeAn2
w+Zf2Lf/MbIIDPBKDivgaa/fL64yJvxfJPWWvV7JHNeu5nJDoZgcmte8h/lnZvh+
yqUoFZtICKaoOj6kwES4k/jNIyPLY2V0g8/fL9Y1MHQYfBhoXeRxTtTXxbgwTkEE
aEu9ZS9VipaFaZpOV+S8eMX4HGn4MYo/u8nyN1yGxIatemKrwkojuWivqIBWdumM
ovuXa0szr7Ux4FoONw/SUOEYqun6YqE/sB0tNl6ucj9z9JoSOdg2FwrERekTEBpH
7bwV3s/kD9TpalGAlef11/YCActh/M0U9mCyCVcDvSi3nAuQj/octoMaz0Mfa2ca
spRqiAcve9rqMa+DN0+1X+k4NQtqh9URJDxmaetTgs+L/RcxJ2wmy61FR0/aecUG
RtJ20WIntBT4lyb35vBCXSMnDQHqizlkq0I9B2/7CJ/6DCDMSAEFGTfZATmO1e24
nC8iGWOtUuiYn+HZDiqQogLfHZ4W84BvzQ1KqN9OKyENiGwU2xfSauY0Z8/dQy90
go9zU9vm1X/yNyZS7cb7AswRnrW2v3PEnMfl2VECu+v9R3Wsk0ZfcSpxBiSAPtHr
8YaIyQnt7HTqxFhgmnENzfKi50qT8VEkuxM0scm+/562ZHQqKud2Iuiqlcmbysig
UnB8EhC3Kn6k8abo1L/U/+JguQuGQXD0MXUgyshCxcr/i/mNlL2y926/M3L4Df7r
ggYJpkJSoj8TeNTT+Om3RA6xxAVjl5XktgJW92hb4tdfOGnB6QD2i2Phr/mLJNjo
MPQOvULgCdoyBF4y/UPy1a4TFTOLkXn39m8dgctHHlV4sE6+2nIRnpfkW1gSH5Or
Fe803//r9gn3OjnWOPvHefK384aHGdwFYthIVNf389eoNdZUAbvIgmCkJldoh6D9
vDwk8I4bmk11P2GmJgS9W9ReUpwXIM94/2xWl2YC7sym3O/a4VK3J+1sFPJQoH6A
vrjoilTcKqdnrthdXSSguQzOTMy2Es/9NpyG9FPihDH+WJbc3T+K/c2MoweKnBRM
EcmqXVF61LdU12HenWXhm/dneHCTQAPdsmwdDw2F2KwpwZmKQXKX1HPUU/91wZ36
8ZAPV0/qK9VH9q4NePd0nnxp5l70ls9MIHQf1i/qjuzkiXaMcoQtz1QUOwTmmEO2
03zq92j2DXbe0bJdaTva8znFunKeG+pJXKjmH2swZg3r70LxZIgGJ2XmHsahEhCB
M5//mjmF17DYZxDNS+gzqZIjNjDOjyfmofzGKIYZbrUifutvAwljeOBu/H7fm7xr
bAr5vnLIZPC5Js6QuZOF/X2hXCReWY3qAhpk8xOYUEDfY2STjf/hvnnRDZZmwm0o
zxVn4vwzhjKcjhNuan0qxCbXd3ATPguNlSRNbb6Wk5Zv28jd6Vs6eXmqCMYdgkQf
hTAflZLJIYyV7r7v+mCo1JSj6BYslFVymh+hKXJaBRhVB8+Jq5sHD70V2vuEkBYB
cv9Z9QNZ690R+5Zs9/pOWAsy1ho1pWJrkW/WM0YlPgxNtY6eijGLn7FYOpECwIjW
GQQgI+sPA/sENccPmih46GxWoujnaBn+w2jyxUiY5EBmy9Ypn79Ci/QiBkwRNjCO
IuUgxuvxCkSDYkdUgGE46QsZnZUNTB22d/KgywCPUx+ZcpRwmYIXqc2RzUSueIFG
yWb9fvuyigNwxXREEFOsDXVY5gHetasikfgyqlCwY+SmNxw96xG2IJPyM9nklCMG
Vszm4PfJ45RcNhqIy/YIYXfdTs8B5UIVm6h8/ln0SJ1QfnSf6b3WAgZ7Us/WEZ7m
xdkgEAWDgEgvs8ZAuDk+yT7X7+0j1D/b8dCrL+uNp3yeeeHF2wdghI9SgNXUdeUF
C9hYAhht4r8Ul3o4XNty5/dVsZ0oPOaPj4dzdg6ZnMRtLKOb7EWJYeaeABJMoR7b
IObpN+JARaGAYcv+TIT2ZcULJ1gjKv+ErBmj0XW6W/rBj4XBFDLB7BRQxpsqQDmH
WZq3dDyXqDnARCwgL9PbRyRZ+Ukr0Tzs/mMiTZXja4GLaaWkX0iRGA+lbwY8MDrf
H85LsfPaok/0a6TMx/axAC0CWkIpwvaEAdKeozMAOxWhFFZRfevzydHOZ+HKeMRo
nQlzFgUMRWIvJQiDf7fO7dLPNbu2ePsCJYEm7kzW5xwgZO+mtff1X0P2drse5OrA
OVyMDrqkafiwr3u26//NkXJP0P+VaWPkuGbc3vO/oKZiC+FfvZWGBdROuBLPaaA9
gQxm2ENlMVxxtEFZJvg6FxNpA4Yt0Wl2T5aY7rVywmVxLJQSMWYhG1XEa0e66Vpl
fhxNB0GhDlsrtUBBLr+ydFHL7YeaWcrPmCXFrUXBEJ+vfnzavmiB9CmWjWvb074D
rEQzJmrhFVv/i1bDf2LobOvG6fHu71vHwwbHwcd7XJ9P4/5XKol9idsTmorPAkE9
17Y2TRozGEp6Rhiwydqqvk+eJz5yBEnCn7OhonDcwFGRPPPC+fhV84Xx+Y+XItlN
Fq1dQOTB38Rd6qhaiKJSb/PGk2sxMr4UcAcjPATsRa6mHZMF8w6Rzz8DTprpup3y
lvNLKNqMBCCIPyV3OcxmK61UY7dxfYIaKHIv5j3XtxtXlCwWKXd+buaaIrG3+tHz
Vf5dSvf4DE3RMgA2lIM0hQEVnA2lPJO0rbwzK1KwopxA1bBD0xsHr24quWZFiufK
iSJM1mQKrnvGHj0pHlVGsxHiTBhnjKDLVCvd83KewCvRclbwFC2MnjpggiZNVxNX
4WBnJFB+9C7c2dPHCSKVLzdYwx6jnr4Ff1oJUMFMRXpw+/Wk9R0Ranh7f3QlTnCG
kTJxpk3P1tBQk3nmLz8f1JExqC2nWVZUETBKCQhVKZ0+O97dir2Sob10pNuZkjhO
k4xM5HyNFZC2uanR7jM/VXudyHvIBAYTxLAjNz8a/JjDHBN6JyXTnGLMvBvvkfHe
U7Qkt05RkDho5GzY/aEFHKpuUuSyl6zF9aMmEUpE0Tkk5FU+VjeszMMsDtHMMsB+
SMjrAMsC4B8BhcZNJqOx+xawxZeW9/v+L4wM7ra5O1qwOaANxg2VEOMUNk8oPpv+
Q7BHCfqvjd7u44FjXLGpxeJ0K3XgnHZPWR3Y+gm8zXchgxoR/eOLgJgj+dqaig1S
Cq6Dkn6/Rs9e+rny4Iv5tAZ2uImEP27NVX+XyJFNPMuPxsT57yDHX29UWMbqoepj
UXBuU7KGhPIfU/T+ePn/iysiiyBvFVtgFGQSgdefKu1VLO5RBLB7wTPeFZ03DsHL
invhDIJKqQGHulBdqnPBNqcTQCtcZ+EwFIvf44RM06jWxjsFJvsD8FeW0DPejXWR
/FD04EDK1uxJtPp3/QVvyYhL/anFHBbz3abHnOmaCQ/wHn249OlQo7xxxCX7a4kT
o7H/SugrD5p4q7wtGyK0V3Gcr8Fd4oE7azRn0vf2OwiUQ/Diwg2+Ec6FhivZl993
OGYBThAXIFF2dvG3HAMRGbpnWZGzBDlt+Cfv4/ra/rkhf+BdsFHz6UvTSdBdx3jp
C/Rtmta6BPuYA76KGZjAUPpeIdpDnz7N9SLA1sccOcyi/m4+ij4/HAx6BCH5fVfc
b5WuJ+ESe4Yta4KuE1leCb7JQnIdJpX2Hhkq5DTjtX4ue/ZMhMpZ/Sm0N8MUUQXO
RqCmWFceAkhHF9xAsRrBafwRh5ZyiBY4sRegQOhrNaaO4i+K4dwTgIq/1uML1spF
IryTDYqKwpTUJZaDK4PhypVIiGiZmYZd8pTn/866dnq0Vc35r+j+6kbzAgwCG0r9
i8pQOXe1l3+yDOWmy9nNwTjxyzm8/NGuinoJku9VuwKfCjnxXoSMmSLnL27MwGm5
zSYJLvygL88X1u3QCgsS67yK7YgK6f3nocmnR8f5aFjMDl5xNfa2H6z87Z0pjCSK
xb/Xb8NzKu9tg2QNUg7R8/9pB61hkwb1aCt/1z+YCaQZ+y5TIqglLw3deb7Dc8Kg
+b9PtkCA5jp7+U1Fr0dGmHfLzh33joZ3OnqtuS3NkgJ2huID3HSZTTvXCyf6n2qU
cebkcVVV2D10iE4Fb11c2Ixs2C6yNV5IJ/UvZUlMZczGUxlpQSYoD3fKoRE6qYqq
UPa7CoGi6PpQhWnr/b1/JZDttDftFYi0kCJLUN4MXO+GNiMua/wUg0DSM5gZTGA8
lRU173XrOGA8nf00rk+znOG6H1kcVhFh6EWEUzPkGAiyVdzPM4SojObXMJv+W8N7
OVhOmXWfXsQovCyI63KPvLvHY31VOIK3i6KpDFsUVe7iCMUjdfnETcdUPS25s/WM
YnL5irmd2WzJgB7lgiJ/sOHodB/t062O0Afv6xQEuqEW1NW3xugtWC6ylbjhQwPx
0wA3in3uJE8FoF53zU4oYbUDRAy90QKlxP4V2gmZo+TGM0NrQ6cVP1xmedd675uU
2mLtxiwK1wHsBvShz8qKS4yMRFewNQbOIslP7HzW06ShQO3N3HMVqQE7mux1knWk
YkPw9BacSc5lHH4BY7zTX3imW3tzE+0AXqoVK6ulGt1hFrVzBooJ+qDW05/CjiM7
GI8pRCUwKT/ZQinPjE7Kp3wP9HMIHrjRks0JiGR7MZgKLPuI4QNFiJT1ptJmTsIx
gcIPk+RS4ZCeN0EQsJSsqXD3KuLn+PXlzUkn9gKAjHzDPjM+pUyZ4vRk/pIKLYwM
hQyrMIHWZpnaemZZtza8xL3CabIUuxF+6ihHBBGSyq7rwIoEMg5LgLMmjbmVsf1l
2vtELpXNPH75pgraXmwf07bZHty692KhOUwga7IDf48mPE2ikacMKmrmpITmkDIc
tyZueJHYLaM6J/WTYmX3qnQnlRpj0adevWZ4wQNRptNC/0y0zlqsPdkpt6AvJ46G
Gc8Tl0K9pSxc2m0Rz69mhG0eNUpPqX7AFZpL5m4jpJ5ORCRyk50dudFzWTy8Fuqk
XQj+aV+PapLTrbJtN3iq6s1/ZOawHq1MN2npd29JxFS5qs+qCgZuGd2NVpPJ4M68
4Tto8OnXfRqanZT0vvkYS4qYAaif9HdunNaanwAeQpcaT+uGLEKTKfYO624B18NH
yieI/ErghGeB2CYqONSmVcDMz7AgAtTxMTenuvMfnLcLfOri5lBRTKwF40Imf2Ay
V+frD7xeeWpPwRQStgwvTTb+PxJOg0pu9QghDmJFcZox03+ZETTV3xorty7z7iaN
x7JY7ZbV25isJIFrGcd2eIO3Bq4dCoiJV4bJhaR9eo9fJZRNuHMhK/a1atw9k2tL
+APohP9t4i/4lEcKINQ8VUIqOmtdC04rL82rVkXEoGSYDjGzACK0dnfL+f2VUaRg
o/tNaE4ilURkz3tIB3YUeE5cY4myu1h+scdBnA53PrVpG/eq030WhbS9KnllA+o4
6520q3DvMIFL/SgnvkZ9U1Hq9/DRaiDxbm8qHHFrRGwcfaVU6qZRLi2drWMxCnvj
K7zm8yYdV0Xka6eg4mg71kUHdw1GccvzlwW0ABs9+MzX05KtbD9WwZqmUGuzYnoi
TfLrdEODoPpVmAeKEbewnlew3fbU4mUAQpjLzPa0UfFKIzwtZ+mgOC9PHAdnFTmB
PZLSM9Ix7rAN6AjBzNHZQ851xlam8pr7xSue0HJgOCz8vegYCo9gweXfXsdXNtAO
8CPuXliMNPGSxwORbCJIUlyecCa/Vd6n7Tc0pXEmwKD3cY3MriwbOda4YhBnx043
hK2Rb3O7TDy9zvA7FZWH+Cis24dJg06hxv1Xikq2fYYDdGF/VQTXzd2qcsDORbK/
ykWSvmmj2TY90S5cL3S80yyN7MhFV1kxG1zR7SpqCiDlAzpfAfvh8vvqSoIpIxKl
UXqir+qPhjLMQ0rg6RhieJZYVw4+E8Z86IWW0k2dgfTxNYkKbwW91+oYU4JI3of+
SefD3i9N2gcrEOU9nHpCg3OKZsvotdF0nJd9zKNQVSA5HAEP0EcVKnP2p7YFVhqk
K3tj05oGo0Clsyo9lPjH9ZoYT+mrLyzz8UfZ9asG3YCXpiGXJwbv1OJwtkPvpIUD
1Hw+M8CHO/7XdimERn+4epSjUnDz1GyktpS8um7gMORDJ9oTjORHEe7fwjZ5iWPN
Cc6zJsvloMiD+F3aMuOqm6RLF/z77oAYC3gNUKRlYDtmB1jsysUkHu92xE80ayR6
23W2kF/koQQfncSsDLphavGOw1LTDRxr0ZD+E4Kwx6OvhiHntQYp11qMbF5IS+Ao
KxYJgQrQ7bNGG3fibZmYwCWlN7S+CQqUcvGdrPTaxmsew8oxbiMS+8AM+JVv3PQM
mVGyHPoFQ5K8+cSNhQIj8y6kEw2v3AiLIp2xensQ8eu7B4PByeRlUrFqs+VmB6KC
Im9blEcxoA80KwQEHClmdAuOmlAxHtdd5RzXNVQ1G8SUfRgba0DH2ZSIhTkXPjRn
i+2V4g7sCnWXQSjJdrlshTT7f+X7tYcFAUFhOymOUlLXpgxzoIyR9dZuoolBoO7n
KzuVlrEYA05gjCZOzL40+eiBnWNVdF6iLgwoAU4tQwirkgvWWxotpGGJeGGIg8eI
7AopAWZmB9pIP0JTmch9HHSAver6tqE51XY1wNLvxmrC4Ue5D7/GIpMvsYaOCEwo
4RO3km3iGsmyd7dzN+yaswhbwIqVxQxyfHWhiOnbmZBbuonNkPk//9aCKOXbIGUT
9o2L7n9CdOLaltIubTWy1TErf9yhDzzs6Ug1y2mv//o9Dejckl2+iwQKNHv6Y7xA
iaaUXHOM9YFYRVqVxWN4Ht8xzzobVFFkDmWPdvD4MK2oGtEZzOBDHUSlOruUpdLW
2WD91eTh1wRZS/DhKkc2xSLvwQXD6wdXc6hfpvJlggmk9Mtj7IJIbK3dev9p+Ga/
likxk9xmo2NB6uhaeYUXrYcPqoJ9m5Vzfg7rSMiTLK0jlwiNrw3tj301K5MYIlfd
x5QZcBJGcYZ/H9L88MtL3c6VfHaM2aQJSzZ7cQ4qnTyUTOSF9ckUWClZwx8KT/bZ
zk2QNiPiJG7lLU4Y1gpeLxJqlomgDTjsWSgOKU+TP11bNRUzRGnmh9Wv/lpvbqoh
hGTT5CNQEgX7TQL2/RbzRMwAYaj4pVrEbnr41GtAoEqXZQRnma6Sx5Sg5G8uebtk
DoQYKeVsIHSDdvf7HQouZCbOpTYe6e+OzPsJ2XkaJHEtR/wah/XV5IHMxt9V+tJZ
IkURH+uyni8BRX1YH9xcx3jGuP8aJ1F8XVWOaHkKz+juPi4OyD/Zc4C72j3uLr1q
G0S/P8yTbtQos8UqbEV0HMJoTJedABphsd0TxKwEr5Pi/BAhBrV04ZVwtrEehcBC
p6hSr5i/wPu0AxJxKcZZ2vj35z0qZtXnB66w7JgazXAN1LB0wU3HFXROwI2v3sxW
W4nCZSI8JtIyJoMbqWjyWwEkx5QP3BtOckZQexBKgW7B+M7baDyURRCLVIJhcF60
ssofPLiIRGITQ8FDZZWphl3wsBkgUh2FHLX0WfEjrWqopOS77d4FT+KAc3Ts4D+T
V67rpBT9JjqHawL933OPOiUainmrN9mx9jAZbGef6HW0qDz+AWB5XnrT42HJ6CRK
3LFs3MxEjJHZS1nqzaGYewCSnLpW+Q9f5XZYw8hK+amdlVTCARdrw6zLOfj4dTxg
zGEf/WLuybvfTFaJuYGniVohj77IP+KvWgenFJoCkzrDB5LHNYusDB1DsIciP16b
9UxCRj6Ye2IrSaMPcrsV0DgKKxjspTo9xTrv3kiqNbSJQppQlSjYFP4FSTXsCpDH
zvFhc54aTLGC5CFubzLQAAI3TbR9mxdRFZWIp+C+ZIg6h4qddwOJzzaD+fzEn/+z
rSAl60mPcuZyqgWrtqTCa6ad5hiO49ELMUrvyWnzlZKfXdRI5fWj0L9eN3YtjzCJ
tQDb4GedChfuHmbkrVlXtfQE2a/gf+En+d2ys3XE1YaABheriUPpeLFFWxybhFiv
oHjLYmYQ3ywSndMgWHNICfM+lT1pgIi3ol2zCbxbeUgU+LpVpcBljye+Cpw8q+Cv
3sCz6HqxV18d9/C0sav4oFNAh8mN1APr2Wiu96Qm4FyDzHHgF24q0+cdNYzeZw4s
kx+e4AVhd5G+ER/s+5Go2Z3GIOe4IUCRda173vaXc9cYPubakWJWIQx8nrMwLrL2
1EpHMbt1080feAA9B/YpBKWOFxEeplKujiZBD9lM8GsrSU7tND6RDK9ysRYIDU+A
Wy69Nwxr7BtZrwD/bRTky5aFw5/9x+hi3z8Q+/Kdx7Nl8zTO+d7Y4WXdvyA/zLgQ
ye4a6XkjLmStlOr3uKBHw6wlbrENU7UIcKMd69pUvB3JhI/SzXSRDA9Nm2s0Jzf0
wE3H6tL4sud/lDDkeVUs/ZRWyxTQWjKZl6GZcOnHv/+fshpxj5VH3uqD/siEF7nJ
BhM8OLsjxiVKgEtmfPROpbkT8xZ+28PDPiLiLoQJpQQEE33oAjSAQymGnTfIJDIc
QieONojn8VrPmOt+M25mWaxZ/Vm97p7CJo8R+ZMa4DbZbx4PQBfx6l40wBu1+let
bSEmpjU9vAxzLtdUeCOcCX5i2RxIqvIeMI40HFbgYo20clrxD7y0pjYPki72H2kk
PPdRsQ84H69kVhPYRAwhKPiKP+zz3lgzYESBuPPbPQJ/ZX956SB257IjTlxHKq7c
z2V4yekZH0a1+DmEC8AuJBIwhFykHCkdXYJXjYTCSTV5hHf8pMWiQ8W0zfg2zdKr
Cs3iHUPio/WWVvuE7EAY9cVrd1K9PuWz7PTUKGn/yoOQCQMxYf2XQb4ht6ZOUo7Y
AjZ/ongtBaZlgHRsbw0ikNdmKlQ38A68evX3E7SVhn/tVVxl2BwbnRRtgetfmhFl
7BdiKY1PkHGu0sJX3ot0KkbZvcGtLlPAOQrwcORNOlHBGpMHrxIftnSJ18x0GYnK
llz5qcvrDZHeknZv2kStv81PFFJpb41eX7SHxY2q4wFBt2esO3AALQf+t+QpRyct
+teKBVIgRYRVMKBauJgekdxsd81JbpWgjzU3DGcPqQxrqWTDcI1xbSbJ5kGYuA4k
UsdkWn4ckr1fLBpH+/VuTlojBVxWm1/hYKTn3PDWI16MTL9R+bUVOtDHXxo9n0iV
4ZFaSuCF2NTBrPNoVCdZ+bnhaoLq97Y2V7ayqg5tDRSjItmIsUMgeEMFIQgvvm61
ZXSj6iJKKIT58Rv1ge2q1WUQERK0q1CkYtcPIR3AzoFtri/nHhd3vLb143YSAK4y
2iVPgcLa8HXJgqBlqVbnhSuPengT+EmgZHHzedqUDl4tZGnUu6oEKgRMbtdwKk08
EU+zevp3Nj9k+ICD4nXOx9BKyNAN1dRul8Ves6Ze+6VfTEwUacTUOMEwsfmm/SW2
dclaa4aNpgzhiMjxoYOz2nFn+rLd3qb+O7TJjYufEpeO7ihM8snylMu7OhJLJY1j
aRsHty+5j23E7Zo9ImIrHkuv0zlO0IQEKBnP0BLXjYAA4LVuBSSAkZBHT4/1RKcr
eKIqwFnOs2dr6uIhoJ9j16akmkti21BMrG5lOSd3++0vKmKbro1uj2SX+BVEpdhM
Pdfk6o1/8HwNK5haKFBq8LHSDBnTI7Qtm9QeimB1k2/ISrVff9piE0aj4oHFLzQH
yalyVG6r7bk9n71EQ0cTa/Jo+9DBW9gscj6HzQRkKDpwG83WpvrhyOT3yTGVqoxe
DcXVVrZiGzUJNix66iCmbjvXo+sKdnByliH00FfuujlP3uh8eUozsZTbsxq66+jX
qbDOeztYVTOWM34w3ay/eqYHtct3oHvbhzK0tEbrZqTYtlHI7+NfFRITvCfgiqHv
yKSHckEZvPsFiOktZXK3TXC97t7MLLmf1K6W+aVnagtBfAVcnjzQAiBP1fW8QbiM
wKwQSjam1Aj/3CssO/o/soR3xZO/40UHqzuelErn7+xNG4qa5n4Ci6VlM6fXDfro
u+5Ksoh7hTrw1D2OemxO5r5vBpSKzQWq1jUF7i5FD7GdVE+TKVotqO/papcyrIvR
dDfobH7VEQk+dikG8YwdKDm59N8TSu+C3Od3o1TRK/vOxHac2u/4cw4eeHxK3Cu/
H4XFfInk8YHJjhhpu6rL6LVOwWQbhZgPGTKcaPXuYtrxwcNfd29xr7PXRC3jNHh3
k14owbp1qT7ij3Sh8vqWesm1/SQPzy2bGIXPDGbpdSEdosabTi1kCrQM3GU2RTy0
XnUMsOZK1JdX3zLzxI5RMqdhq1hjvnHcj/lK/WGux2piXs2dPkCzi1v6VB91G+Pm
ze1ONI7GhxgufR8LwBG2BUCsxsrkxRd7vbimUoR2S6mpE0tW2YOuHmQl/CX7Sif7
+4vYKt6u7AWIqEdfSewn28LLrCehgpmcqrG4XeHHGVXaZExjWdFumGfVdOrWsjQ7
0w7m9EVk1kiedVImIFG17bC26+lCBDM818ZhvV0m080qJ9xtTx4+PN2noDQt4cir
DinHLyVCx/FgJ93J9ZUu/ta0AnQtBp0hfp/QjlS9WJNU7bVX/C4PARsP/dr6PvBO
3LLs+fzJwqkEZzhGfiyVeC2MDUkHQTTY9cep6osFXUQoTtwwQ+ZO/3lFs7p+ztok
dBGaEv6Pvv/pWpEOBW/SFCCXzD5JWQ1NavmlzpyiGCpb2UhdxoS56Zy/AkV1VvKm
i7II6C6acSpWVvCgQIXaoyoOMPR1i1SAdZ3kUPeYYfqYidiW+0otiaYAueOcHFVi
BVAr3qIeIcbXXEWeGkJ0X+D1a2XdwjMd4qBHEvxRpcOvaatd4CAZO1+9LfqykJO/
9obO38QAZB8/+N+VeTb/k0WOdDV1ADHve/SCcD0vcnPU0XkWLVOQuhjEjpqCMAzw
BV3PWO1m6EeNsdo6wWSvhdtUiTGYELpPvElFfpyFpxJOJMo46T35JgnpDlXsjtks
ttaVjDrLJZJUT4yhSRcNCWU5AQWQ6HUdKOxSI2cFReeKCFJcyx3Nq9mtg/AH0PZg
MU96OaVUt6mc0yWOn6sKXPGWh3Bh+ZcgrXQJa3aVAc+PqATe1D/2tTspJDANGkK/
j+4pDtipVSk3Mq7rBegbk26zr2eKfLaj3lOv4O6EOQ3fws9iVAGB1KNYujXQWE4y
szBEZW29NZV21GRmR94n5jx4wVuPmGNtL0IrmmeiIEOZLj6/UZNOas5129VaF+g+
CnvqDX3nLLB/vjC/f7PQDTdVSJGdonSSDY0oFgIf+YENqQtUKkH971MKc4XMg+Ye
EddJ9nTNT/XcbyKrfOzgr2yHxEjyrig4FBwuRv+dS0jL1RR1ilb3TeLqIinuG3Cf
3v1h1UsYDGrZTKnqCRUv9TS7EWwPOSEQCIfVbrEbyOPv5zRosxaVBv17yR0X8H6b
EFKyJgS9F2BBYKlnskuCqcBlKQxrg0dMt/HQOhBNdM6PF43ikd75jkr0DMS+37+E
8W1W2BgEHTs2hpZSPJnqZ1bpyShLHhzcwgXNnLA+L+QktXcfzXdppYeW0rj5e+n8
J6mcH/F+RMoT3jwYZhKn4PFe5TPBSXl7p84a/CajEwul77wtva2y7fz80ev0wv8u
4wJmzoJrvtQIJoPTKvbfPnloItL23q/D6xuEb4Ft9jTiPMIKMjKuboMNFy/5Jza3
AVOXif3eRtkWedFkxjxwBLqgcjqmt5duoSshWVumGcxIauLBheiSfBqhfdNQs9av
5W/EhspkvZGBTTVnuD2yLGBa00N0WTlLhoI4oaJfKqJpzUm/v3IoV+p5O7wZ/ZXU
AfObqR8DuTrFRmN65Bj4jzrcKwJ6p32SeQYfR1w60LYTpOvWJP7BrVh19P6t7qYb
Y1vAQFbv8FzqNiUxyXVcsXaqBwSSPqS7gIvUT1lhjJvhilRGZHWH+Tj0s/9LTXp5
IkAUOpTptwyB5Y0QAPwiwRDqg+8ofsvuQX61bWB9txb55KLYpcy042iGbXiqsxYX
rEBhsAGfjlVj7U8TbBTP6+35PoNCXDCTxy18Za92eyMqAjMsG7BH0xvesj6yhpb6
IuU3p296fkYnye87K9Jn7M7FaAcuKxJ3IRufAKH+ooHQxi1eaPiIl9KEImRouqHR
g87HWzXiB0ordUJCf/3+jDDQWVSAl8s9tKf/mUhO/xkV1pF5M6p6J8tgA7A1tQZo
x9k0LfDBmgTxknJoBLkJtijH7VnhtXqBdb2T6HvdWVF+lU9+dW8PvHaRuQvj5xGr
DNF8R0z5Deb7FHCvo9Te7wgq2kSz6lIsNndjp6BlegoBsMWuq0IyOqcn2jnYCe7Y
3p8micgQ3W0Tml6b9gtkRHH5GfbvZK9ni8mzF5bl4azJikiZc5lGDkkT3FwnwgEt
S3WSng7HrGZwscZAj/7X3DrqOtR8S2fZH5bZgHdEcf6UlXyH/A64y8UDl//H+IsA
AJ6tmmvFzCUP2YPFB+0pUxjsfiChIJj/iqbeN835VW/07JtMONx29XHNADhviabG
UYo2Uf5ulGDEe/TbZHZgWHozgEY+YUcES3L8vwjwkZ9OoYCd2v948qjd6QogN6ru
XznVUu4dINDLrVZB26ZIu8VH4C4GrW038APF7jAagUqH21o9H4Vs/y03E+xysM4R
0j6oDJ+iVPRlLxicD9KabFipjhV8gxwrQNM+bMUgS+oSIm+QHtgvuXRn7jFbvfMQ
3zQ0f1sm/IBRp+QBup4O04sVRjkc+iw2bX88djuofLYAOb46jxsCdaueXkmGMTrH
xs+4+seylBNHUo5tup2Xp0vdE/x3vjp0nS4zY+FSFNtReSIJdPT7pl+yE8zDXsBL
OVZUcWaPpneOpH6pU9R7ReFNtMbwd4lI1D1zDCEBxZYc1VXPfYyzwi7kX4lNJnu8
qnOVjbxDmryvlzhHaMEUx0Y4KnFu7Vb8KMS/7uob2Ukmqi0ROm5+b7rYnl94l/x3
jNf61SJWptvpmCXA9fafXa0CeibUTFa28JQNJEE/ZJ+9834LSdfJIOZps5VrfDcd
x8n238japImdQL53pmYnbWcZi2owABgkReqyUcr334GE1OnSJFnKK9sVr9vs56rL
nOqdSDX8LPRaXwqMdaayzN01ATSiAFsBu96rrR3gKU2r4ijze2QST6vIkusUayEZ
ZwZULnP+ztX28rjZBZezlEbNahQkSIaCKLq2mLI4vOMIYWU8F4ZbJoGaJhR0AWyB
mDArgJLTO4s1PZvATLi9y5pB5AVaET8/sKYnoyHecRvdRvV4BYemNUrOmeB1FAvL
zqyHcJkDGjCPDcbd+DXa8Bh1u/hcT2piTMk4OL7OFWln/c4KEOjfbL9zIWyMQ8y3
8sC89IhaC858XeIyRwq73Iln2L+iAEGjxdnfHftHJIRubO5zQ1k/9GmzuklTslRN
jWyaOBzcCW6h4dRiI8CkoeZjXM+nRIe76RZbro8P4RCVfE79fU0VbtmEonJortbV
TY/Y8q0unMN41Wg0cbMAR5CeG858f7uXq3CU3LIT7I64F1DSIYxfK2tEpeKdNUP3
aZRD6fB7IlYXaW0I7ti7eRlN3mIy3lgATYj7NT1/8vKM904GzlIgZbQ3zRuMC4y9
ZbihCSbK4F/ukrZ1jeQZNmRKxdiOAUzeLeJyg7xuh6Xy5Z/vechpjvobndEzHH2Z
yZ6Gy73hT23iWnUczeTcVyQPcV4uesGpTJCEShR8bJfCp/F5H6/g4VM56YzmmOlt
KL15+arAL6EjWOy2pWnMTtmblKMvQp55bboEKnzfYU6etBFdJYoYuedwlJyIoYzE
8conxkH6/+GiUmb2S/hvn9WxKYM2H+C84ImzbZ3Z0dls6ClFX2AKwp5nJxGxhF6D
rItBLZpK815ZoNe6msC6vZeYepRlEUyUTvpKrdV1A4FoO5EeSfBtz5siC+bKhKa1
iZl2IGsqHodMKRroASFvV16dlp4iKTRiyXhAP2UgZhxuL4n5+6zB2ESj8wLXav/v
Bx348zQoQT9NmiD3pGOMbEWcLLKpi4Yky3x8AvruEIKQKiOL1dYSgUQtxv2S4wgm
y4roDiHMfR5adDPwi3VWF30swr2FSGhgW6epEXihXew6tGy5QO0J15jPtX0HNWpq
fbp2UNVE/DM+vsqXFDaOy9SmGIVtCsGq5IxZ//C2ICbNeiWnSUbgdwIJW1Qqn4We
ZLKgUMGF2tb88d0jpscvNUh6uQczA/bY21fGANkPfHVdDjww+3kLoWEiVjRlwa1c
IRZQag7ZnjltzDoGR02dNS76v9cwDYgKHu2HQHKPYb4F6do75LoqyEy/qPPBZ9iP
dBXuzjV9TXBSoUXeGZy3ensToRSSoeY3xVT9AnO6By3QGavXchYoUYnr1yF4J5Dv
b/h/UOqDBBnOk7rcw2d7cZmYR8xNzhIclx+EhQiYuAFGVD02qm0Padnd06E4FQ3q
TgywywEnfEBULKix3fDIWeg1jvy3zzMd/xzGru+tjV0wD8b6y6d37S8KsE7u3kR8
0yTgNXNWxNgHtCdrkzfjMc1mrgsCzf/jYUjoFPTkab8MBH8KwT5wXLVNu1aIGFWF
B4+Wbch3thsYv+7gqW3vTDrrz3c1P8xqJfgmUiG/IqCU218NtM7Z7llJ5myRTowB
59pnCJA3jF675nsdcL8GZEFrLXflh1rN42bRcne44vGKkdckKxe4UrtPDrw2c5tF
tEYwkrksfS+dZBPGY7GdcfNAZ/lfDg6PqJrecmLHEQ9Xp8pQ2aAa0A0wo6W4Ogvf
2B1vCZbFsYlOpSxiDSdjKKVj2mG0YUXTRzBKgVnj7J70DGUiBkk4210vuUGwDLxF
meyPhz6JEgDbNKiWaUiDD5BlMDpDDtnaEpFLqz61KXBkCvlNk5ASeJbIJ6e+Mhc9
GPHQ6aQGrXsQOhyrSfk7TJbXYruGd6M5RtaL0W5U/EnveTVH3ZIocSycXrlOcxBw
2fiPhL8y8IHQi/Sg98R8SA0jTuqgMSkXWZrMZOfiPSahPUFLpkpOqWbvBZm+U79p
a3xw5TEz1klXD2kIiim/j5gTxmMHSu+mRmLv+xUgMm9EdNl/Lu40kmGXK4TSJrP/
htbm3HoUWYlQgAJ2GqXDdKC5GqOK2+bmU3cHhPjEIUX7RiP4QYPPOTwkWOwwPWbo
OXa36cbUBK67Mut3mAopm5pod+LaIYfomKaEJra39ApsbM6UXi2cT9/P1+f7Xc64
TIkGxY/XBMj4sPYTrUdrfzsYaENKmuroeXeANwCEbPBXDyiXj/3wVKTYaEjIRr1X
w4JAqwE09AXBVMC2PZ3z0upU9HSwZQRTmvcJCpNExdVY6WZfUrzR4ocVnVDRGDMO
xJFwCbfW6di7AqBUoa+O/DYRtrtWrZBvNLKJYZg4Ay34ywJ51ZND/tqmgHduYrof
R8P7EdYneU++2kvwpD9jLucfUd25C+ScV5dLyMVxamAc8D+3mx1Z+p+JyjXlQu5W
37XI2OmiMYS9xlCawCvyEepw49LUHRHeLyefRAOPnpTFbD+CWWa72XR7TGnoez8B
wUxLavpzMSbUqISLcgko8ltcPxrO6q5NNrLGX2BCkAqn8Dxj3sIed+wty3MGDErI
PqrLwqQYfk0LcdByIGDIQoqgHTWBXyR6+SZdDsjxxKlmQXrHLh6FGHH15PZ0XZY4
C+PuL9YH67YW/5DA3iyO32/F35Hh6HTe6ymVUWdjnPwHHOip+TiiL7u8a8oFg9h2
Fp3AAzqhOuyhOyoBU4j62nsfFDrD2tvHS22M6uZD9+UlVf7Q1qaRrwsDvW/5a4J5
fwfsvBhdFLOktGmVL1ceuyRy/dwLKkRRJdEZyfQzNoyw4TCfZFZ5+O+Tl9ReuWrP
Rwi7y3Sb+KiyrQ5EvWaUFfFH68NMKSH3JMSDmNdcJs8R1dYm1/DRTfR8bX+S0+pm
gFTo+6/hnvRCVntUp5tJ03IjWT25116YWNteKVrYYDgzQVelFLVuUd8WECIwGzXg
k5Bgi/rUdHouhcrh0yA6fvQL4H985S9M/ZkMjZ2Yv73pW3BnEr5VcM/NrbzloDo+
R0foYmfmpm1ewbSEbBL62xCqPWdKOQlVQWKJFB0WVJRVWwLvQvGN+8Pa5PR5wlwL
gv0lIXPYWSZaJjRl3nPf1IqwZfeRZ/7zZ7liPRlNdzatWHutH3bFlBWsShxXbVyX
mAUt7CrjG3zksFhY+aBQWbvMbl3G+M+bFXpguuzvtl4QymqaEXhJvIGDewGsQrlN
/K6ODAb4PrULNhnvvwzUxO4rwUKYMWoYh/IyUSKvYQYJqZLIUBAlfW93LfPE0QN8
hKZ88N7/llt6aVdYHZ3gDuKdI///HDF7k5GGajyr4c5bAkvpjKfOSVmVnJ03UX4Z
yYMEmosWZUeC8zhGj6y01hwYY8MTLyl5ohot4tFb/2r1EiYY2X78E3i4slhnHdXh
WXmWb1Mhwimm28RuIZba1fNFvOMgaN1dBR7yhuO9dreZ9gBEhhu0fLa5Kxv3J0ut
9jxGOtvSfND5K6uiwd49AMk/hR72W3943J5Ko7gRy5LbVjavPIvmXTR6oUGz0UaR
UQsVhGEOLv4zYGzPAgqQbGv5iwOST3yAsxg1dTZ/NOrElGUK36nsYQeWNeYVFjh5
Eg8bjJ7SzBmzG7dGh+556CJzPgTx/JcysTch+AZYGI2A0yBbMEoPWF3LHWdy0cj7
qZa4dhDihaXLOqSPAiniB4vpV+sqlWTys/hBPoReF22lFdaywonUM/g2nU2Nr61W
d/+V6D2qK8DtJJrqQnwu838pitYUeZZ+TI8pWOoj3jxiH0v4t9ztiOVzS6XlAQx7
o/+GAV8BuKKOaFTkLt7pfnPnTZylmMI+/NkE4rZuZwQCJzniFjxJeeTQo8WOM2Bh
tUlgHWbVZGKeBsksVdx3DEawz3kMJherCRGfBr0T5uHuek1tGWlbHgfxw+iHyIvS
8/3HrTgHzmUBRURSINOa/Ec/+uCJU75CSjy/DpC8iaRnYq3Fjru44xVUcYaAMIqm
B70TkyWyVM+aVmtbpNsVvf/t5S5DdObnwkFnRmzfIALqRRdxbzxgC5jPXT+0y59u
CY4O04pHzXGyCLWVH8ZGsNzZoHTk4aun9+Ll9zsC64NpaxUKiNnRNa7cSdYhh9MC
X59lWVT7lFo5GC2VsFuorSMl1QiUM2mIe+N/sYhWHcVQP/JxBj9URdmXjONtUx5O
+CGv60DZm9d8LfKhMwS3T+o+Zskiazg3sKDZkH6t9vzesw3SqJx1k7sLNGCgYYz+
Og0LlLfiWgAK4Q//Yw5RRmWMPUw0qUSw7oh9OnMaQ800+HID6+6HBjmS1JAZyoWb
51iXe7U9qSDuw6M1j/FS5HWcwPCqyTeLXEKdkLHTGTJXKAr2zJAbSF+7E/7p5YjZ
k7ZFJL71BoicjOxR8H1JI6KGrlsBMtg/zkn6FJtGGsGaDPTIbjsKUisGirIzVxMY
vkyQf608w6772mpPGwRHJs7z1BIe7WYd3i7QSCKidxHzmcxMsKztu6HO+d1EH4cL
WZZnX4MhRd1RbNtuklncYIyqRCu1Dq07mgoe//TGfe5t/o/ZUEtnan4hCe6RbEXi
3b+/EJXsp0X+rRKTwz4H0IDgidIKRDFq4bX2umIatbcH2YsVyjVOEO021jPz2IEQ
GD5ZCr3k7opLScZlMTmrRb8GY4Gxmd9mQWYGJPlYox6/iXJe3ajk/IOjYbTeXxC9
mFWyIfxBU03HApQwR/4wz8otIcp/eik+LhYSDIcUT8NikLhgyLPXchn+tAIH0l/J
WThnLlj4kdwO8i7r/pv540j51jGCNfKPPf+a+F/GhzCsCl7T1wxnJz0McMn42fE7
XKa+/5HN0/7beOdv9Gv57ZE5SdwW596IqPsZKZ8189xHZA+nKpgJVY2EDuosdl7l
Fdvh/k98pZKk2igKZw6KPef+LyuFdtPZNa43ATy8uwLBIL4vKKTOeSyMDppvwpl0
MK1Ud49YtymPZ/VDscDfSVr99NtvyiMwwaCgUKyGIMXUumHehFniiEKlZDv0V3cj
/V/QlkQg7PYgl4Su7O3gVUhtEkDeWija5kux2gZVkVWe4NEXl6uAUQR2QLZeZ0Ov
CHOTvFMrwfLkTL3K79qHOdhy22P8kvQ94S+Qw/s9zwBjmgIad1lTRnMz2DzlIoGy
/I+GtE0eXE62rio8zkjDoQY/aldg+sFod6E3wS+zdXH8OH0N+CYmGb2x/c01Klv8
+L6yPdDwHMwwOLnKM8BSYQuEfqUr6CFhFy+CpKa20pIGrB+TKzA41Lm3J7NOKPa3
ySm4se2do9mYwP4/ww+GHS0DkoAMJBHrdYN+eFcoC2d7ZNr1VOgZf6CTfInwBDHu
fpCHDGugiUUDOKg6+mVr1mkRfUHWDX0qo8MZPJWloT4Wq18GxLAYXKscYDvCn+If
ztVpFrDub9+bbsri2soL84Lu7w7zd6OA4qVskgF4r/5Xcld0sdZ3bGcwOxi6Ga7r
nVyU6nTAxmuyXjj9lgqiZF2gsGdqplrcEYDHZvNt7G2FjAAdLv5tVufHwDLVXTch
azE64RyhKY52CEm8vR7m79QroGS28e91tdh2fdRYhoviRkejN3kmi83S4BIT7cZR
DtPlVkeY1jHWoTOjzmt4yDVJQr48gT0g048LW8W6fk6R2tNKLhs050dbRYLXhIro
W7VJcjztqUveDxqFJaQ0/hxMcnQ7SFWObABiYnJUVh8sUL0iQlL4eg5H4BkrTtbq
684aElu3DYAsI7NPvNrRFuZXlGgxtZ2pvRBazTZRWZjXSxSWxCyLGdDdfLvGJUc9
L8C99kzqak5ohrA+TxPoKWdiUvuyBR9D88BSl1lzRKno7vTEC+wwZUQEbazsmOtB
ZaR8i+ptC8S22krVi70LuhSO6s+mXcTeGu15PzFngyuOwTrQfYUez2nm5YXlanll
wvkfMbJ3dXPxASD4/2ILpuoQpo9QOXUd46YnhBLW25m6z9d/cDL7f6+MfEezIrvv
ENulYQKikGFxBa0pwZzOFUW8QliuGjy0RAnzcI90cw8dZ7VHACP2UtPG5Syv9mT9
y3esi9bI3KN93CMbBTNVTseRgWTQQEnpdZetPhuojTqEZoWr4Ar+5bmYn+T18+bF
pJnZko19VEO4bP+7OreoalgW+PmwNv3rI9/FH29yWIt1OPU1aegt4PZh35FQgffa
/4g7pyjOblnpxBhLf3PEyrTkFqe91ZuqjJLoKGSeKqzZTNroeZFrXi39fPbkWSeF
Y17lhjsuyn8E/mfDy23zuNtX891ohFos/ET1WHs48O5/jsSqBQTnQSb6djsms6Vd
uXTl1JC5hjYv/HpSMLgtuHV2B3tKjm/psNOwDYMg8HdIoky5ASjT41ACPJoz78As
MUdbOibGFbB9psFVkVKiIXsnXCyxSEAeRZbdcPV85nTjflZNY6h8T1ZRd/GYLSuu
4Pe3kHjxrcisrNvaeLuA2WzDyxIVaLlcE/Ad+GNHvv77IwffhDwvvDMe7Gk8Y+7q
KQmgGE4elKsNT8GFXRp9TnWzxbWp5/JAkwd83tD2mcyH9PnmtPN94hiVNNyuVXVd
x8wNYz5S94gFPjZx5hjRB2L45XRn+uvSmWYa/ytBnZXCETXREEB4Wtx8FcQhISW2
qZj5idMqC+PpIXT6CbxhaLa756LB41tiDlsiGgU6eUNnm3zESHAmpLLVMizGtyGv
sJ9/mRNcQWQyDiRcAUCTNEy9k80+D2LMmTsQu15UREchLkDTFot/oQiWrEI5fuJI
ZqjSRyQI4JcOKCIx6LkSMl9OcCp5lSBPN5uPcdKU0XlIYTqqR2YvrxtQCUdBWY0V
o+/+9paGcfDb6NfhxxTvudIEY7KR+LbZO4mYdupUzCC1BM6xEN2whg7XyxN4WxS9
N/zKFHCkmJhA4tgYWZMaGDj/2UWZa1OPZgYQ/6nLOcU1BWEplLG9E65ncWhXUPgl
e+x9AaJMpSTQamqfH6Zp3bF9VH8A7Q5PcD+PeDHSzD1XdJ7PUJBkcfMeR8fLd004
mhWM+60v98sb3QSAJfEv4Et7q2uaZNJbwDN4rGx88FUcwHZCBRPyHW4jTRjHWZGc
EJcqOtG80Xwc66kblDFparYChR8uSjlxIfM0rWRBo15QVRL2mLZJjq9EmF/8Y9mR
Z+9WVQONfFgzS1/xsmQ9KZD+bX7cA1Q7Wo3JIj7WzrHAegJV7Pya6NJm0J0nLdv7
/ZOG1/1/5aTJyDxrlBtM21n/tWBnvLiLwWsbDOp81gPXDvWhepfPeuSNcThaNsE3
9X+TbpGvSlQHOk9JqrDGA2eJtqGRslUDhzIu4iIJPfo5wR7p3Q+/bclVTFlzfc/t
AD9dj8VWBPKz95d2X/4sIiD/ddpVXR6l72p8q9uM233coqNv+tnwSKWlmku4G0wr
hQNvFuA7QY0hiu8iHHAA6NTcJRgcnslIV0rEiiu/hk1XzxjBNDzEpC1r+zT3EYy6
xs9jeAEBsTjU7RtkVQXXp1eUoeWPtUdpdHeagRYSHlSO1KW8aYk1WIWcUd1YK+yP
k6A8N5PNNjbHTOW9rwaAg9beYbj78Vv0OlksXOFnhBfu0k6QY9xmb6fdsUMLy/GM
AtjBcjFVWDOjMlkOX2OCRpoivKP/2gokOsAFr0gYlpqSWwFnG5DZjwJkxKe4SRM6
vZaJohYFGBEYM+7sn30OXShq00p7ylGKcdrE0ebndqQ4Q21SX9yCdZqOQ+MGXIkX
iHP7kA5W+3shRhSL7/rxbiVijofR64PDh2dtBp1iDUdxciEK94Iycf0OkpZFKoO2
Ar52/yMQGU9koKO64ia8zEZXG61D2rS8LVFM3LZhpTZAPKlX2vQiOn8ma7Zfw6vj
bSrxFjmJJs8L5nuQ3+oZ+BRXnpRWVSqNjF5qXTnXgdgv3L3DtOZzxTwCS+zY03Y2
792M75iPd5bm+wztIG5dIus3eGaBpHGuMPt+5OYNezeLhV1wlW+td7NereTGkJDJ
39MpmydlTj1XrsoGwy7hVL56u3sn06GO+MuFKWH2gscoyLWQorrCsAyhoZfnNglI
2fDKdO2P3cDAAMFwgjtENkpphEf2g00zFgneV856xpVi3Q9DkyfePFhk/zlDrwS9
njgSTqV/z8SaMGZYt8z2r+bRgL4fyN7xdWCbP4eaxYO96lavzcYwWPrwDCVrN0yl
qKHBsT1wOTRiOVKVkNeZaG/g+s0FocpevgZLLCxjku07CTZ1no8rIasK72Y+COsW
6mlzMPe25oEkXzHX6qCfcgkVoGTWvKRfAzYB5ki1T6WFt46jS4mTXIh7qFUdMjDe
2XSS80k0u5AEPJfQpVWoAl6w+nCTXUZPjQgwYr55QjPWIK9AwiM44AVTup55AQP/
T4jNNUpqxi7d9BRcFWmRZLr+bZ+X1MtBonzamCr/PD2NtNtNmX+Taanam3Z0JR7c
flsbFQ4ACiBIcVhwCddaKgnpsnjnCECuDsUYS/brg3M0Vw+g+ALX9m1JfWpLghSh
G3IEhxJvaZ6Jb1Y9tMXNj7QKDQcwy0hc07MP8PD2wIKxxxX5Ogdl2AY6KoO9O8+K
ptCpizaTY5sqWhsIXZvbzQ0Q2VpZJ+Fl6tJrzhUJ038zKfb6FAy3Ke5YF0yFkJIY
OzwLdHWXD0WscokOLs0yZux+gPL4zEQoY5Zw7Dvv/J4h9pz/DDNZPU9WAR1bet4N
o0m7VIa/aTT5Ltqy5ELPhJ7gcKvsTIUQOLzaqw3xBnl++Pas51G0kPi+O8NYZcpo
O0GvsRzEm4XwLlsHUhJkKOdRd+QyCIwDhHLyxctxLMT0OqOUlh1Iz/B3LiHfp7ji
BV5zDhGegTKw2IdwRT9I6Mp9PJlPW8G0JG81fTYL2eH79HHIQvwZkIPSWLQ/6v0u
ZwOnKKRGBp10CR8cL4u8pP/M10DeIax0Erz3gJURF2dVusaMYSd0FYEyUUalvR0q
1SZXfBKhNdNPWSbq/fiwTb6jyAsjEJuBfMlrPtiAZJnEKG4Sbssp6b3bkOx1u3Sd
KqBck5xQEY8ileD4Y44+efsKSjR1hFXozesZROPdQONrtpZESHjUxepWezuiRWH1
mnim7a64apX+mUNpZu0PymcRiOi7oEctdLMTnOE7P3NiUgKmLNsOGbpQdwYiPRKm
/XhSODnNdgC8MbpLdN7UYnOOc+WPW/LdILIAzNyZtNEgSW0WlMP4BWpYCTjg8Hdp
cQZq93xMkRORB2eYEkRqdUaiyEGykYv5Pd/LgocjnXLoMz6kIkRP7CBfm8f27b+h
M6PInrvuW5xw10m1ksaKcb9a+9XuLPFY2bMyKAdqDF4X8maeDFFgBRAocbMVDljZ
zDbj/VyyESKp0aRgqgi6SXpGdU9pLfq+mKHAR+3gWxJmc7b/Bh+U++/2aJ541fwB
9EY11ln3c2CKOkSXkCSeJtDqTHtztRfuL9AlWrarwTqsI5PbgmwREMWm3O+pv4e6
DJpQsnH5aspeyxCAVeH3AebFRwh3DYu5cttBwJMJKNyv9w8HZV/TFuFaUmZwEMFL
xUkeSnMbErxaV7NQOjDiVMa2TpGkQ/lwqsTXH82sj50w8CGf5+pR64xEcarjROrx
nuBRxljqK1LhcFTf6yzb+ls15h5vAPc6gmAlIGDH9UT9EI2u/tqm05VQwGNUagka
lQkRVZUyIxJDYa2066lQgMyoXy/FJoKhxOGcWzuBTAQi6jXxwbMIAvNehqaET2Uc
d78K7vLxltCQoV6yQqdxuMYqTG878N14ZAOxpw9bQagEkkYerkVIbyWjF6kbc/Zu
YAGOVZLXKSA/d77GuEvWXazTChcpVIbcthLjFRRaYjFkVy/JhqbYUTy+AOXnLpwQ
71VEfU+LDYc+XM/I4wpe2DoEFMg2S/40wKHX2qGZ9V6mlmU6WTxS7ONVQMtOakAZ
jwKKLz7+cspDdjz6K4IKnR6DwFP/RY7CrmSIrTPdVq1VOYqwVvVCcqOA9U6Wochd
5qDanmbnIgpta7pDsL9uVvil5AnOpNCPcrmDE+gH3kjo762AHeba0uYFf2fBy1uh
+WCrjBuo4328FkLpEh6gDFhzjk3JTl7P2i4dKvphkXfAasLGxt5G8ZUIdC0cMA1y
H/O952nabWaEnckI5EWpPsb0wCmk/639X8kzSKDG0NQcs2VkFvvab1NqatwEHk21
aTsmTrJDUM/ffSYu333wqUJmtSgz1Mm9REH16T4tQw61E/jUWKtGBMv31I1ZvaS8
Iw5Lieu09R2OXniOHd3lwaKkSPCNZ7xgN4AbqYyvBRgf0enP6SycLsdSYrtRU2kd
TU9oe+RtjaL8cXBT1GMTzf4zOmSRrROcNP2HmhOvGtTqYEWOgL+lTWs7ycZ3DKeg
N5Cs5IzHbHMxPnEw0xPLfU8zPkogBoj08AyiKF/Y5g6jhWw/hfmxUwTk7Ext9k1r
kyGE8wBbK4R//cWg8UM6G0ZmHzH5oV65/OBvWv7WjcgNSFskFHyJ+i2oIy/PO2PH
F8GXB5HA/BRSbOZqHtB/0nRPS8KLQlTy4GGqFbcFPPy+fuy+HiNrtFzCMkNPE2eU
XswW70yIuldq0/EAHONerP92GwYuJRAYHtzWylu2nkcSSgGHoILMVWg5DSwILnxh
541iF/j+w0I8UM8zVuIrMwLyHU/3bLE9YX1h4j9s9R5lVt4+EZ4xIHpRw9/2tpBs
/76e/qY0uyQSAq5xCNcGNsynzgP+2cejyembwtxXsbC5mLW/OFS5CccecLbEL+n9
QuTWNORPZ4eEPy0XVqYhzm2wxCPfRsEejcVdYVoiQIRcrqBSqzcUo2IChKrZfNXD
Za7HZ3iVuYBzS9O7xlhiK6wKlVnWYC/Xj39H+dtSwi+YSQz8wVlrgXeXX5hgyhTK
IsHIbfLjVwr0OnrlpxVu3Zdj1XU8pIiiG+aJODhwMI46YCx4JBKLh8q+ytsKCpYd
GYVm81vICYonj7IH0Z9FINJmJfJ2riEQpyp0LpGB37SGwSsplVm1IWBamQrPbN6G
8aGHUTn73h/xFYUfFOteATtTc7RJM84gLGj2ihwQgma6ldyQ6tC/7T2FhxBYR5YN
rdO3s8tPmfxIi24kBJ472JFy/4uTsUZB+Byb1c8vU24LjFjWP7w1HAV2RAg3mv1R
2krpUZNH+CeAQYJnddUvoOK6Hes8OwfizOuSQ8ctnqAFMmSaG8f8M15OWBq5z4LS
0gHzmafskHCUVnIufMqp+El+H9QOnaBwy7W2zFJ0nzYw0tLfFGgWE8TcPwLGVoOe
Ime/PymBZ+pfEjfi6GuimWsBXnxYmWeUOKCXlgGHVLJWstysVTSac6BxhvJdYqBE
4eRLqjJ4+tUg6TVmV/kU3YYNXXEowLojbV+renWSLD8Q8NwisrVkSRpbCWB7TKC4
+ATOuxcesyokVoS6dTLOgQFO5A9JXx4eZN5HjxrJUz0WG2qwY7IbptXjLYa+NJRY
w9zB1UYDYSPPbVJztnkn3UZgLH2t0FqgWewqfZ1H2+0XxTpBnMMsJxhCl62ayip5
dEuMBDPm8bm8C86TvX3egkQWWA79D1VbN3yHhWXx4VRLECUwOtSJqAH8JcR/R80p
tdqBoDG8i9xH4RoAZL3NO/0+roWsYa/vJHBm+Q4f/zIwjUAdge0z0qs1qrHu+/vs
j7rguI1AOwX/ShP3GmS8Eck6StcuUEWEET1hc89yx/SYnW5TBWQ9XXP+ugwqnxN0
lfk+7/Vsutf8lHVhkcI2hOCmqMAxjQ1nJuHbKPh6X3CW/bG6iOHzQJ8GpPEJ25va
Z3nHrdF2bxemTWbHfWiWl74bIaATlYSL/u6XuM79XxYKvtZmM75N9HVs5Cf6v0wS
HFhSuHAoc1SvVDuLGMNNY2CPZsB86vO9OF5akWVh6v8jd2ZQACO8KSwYm7yhpNg8
eo+8HBjMB1YVSWcj9vCRPg4ZJVvJkOeQzModEpWYFXBTbhJkKDtjlZ/529ig4XjR
h+LpYpT+N3FfKaA97OPhL3aBzcxz1DoDnFav9zvN38t3JV4+2mDvCD7WLYK97Tuy
zVQYbuVYsOrth9SgFIHe3f6sxcHxT1j7XZXN2Qi17pCWYzj9ojXSPesEA/csQN+z
Tsx/KaIddPouVH7TUkps9fxC39vpsFdTSygZO0YcQxfChOD7aPdX4vTBMTaUf/oG
37M/diEFXKmZ8Mva8KeK5LNWr7wVXOR1m7HsCJ2BkG+b65dKYYmfsYfU1BSLE2kO
v5kGHNT/z27UVbGa7tfZhnUej5AOdIHk+GihaKmNZh1Dvi7ysBqnkIBTp5tqFB99
qcoOaTJ8GXXCgr79hRQVI18Q9MAoH5K0Ak0z+SbphflWIBNeLF26BZqDeVnsYAjc
EobLdgmWHl/Pos3k5js7lzypfMcMmUSEH26k/lOaz/xfV2fgTEjFXBzVIXsAVtQ4
abd+++K0cQ2QUXWzVr4MrdJpJ8RT63Kuzq1hRJu5wuVaTbumm+yBPJZ3IReUpGOQ
IA0DGu4oQcDsLMvUEJWrs0eg4G2aZIS037RAOTgAkbViAwOb4tx8WhDebCNXpeV0
R8ZUnHClOzDtUCMeRSvtKpXY4DBplr5P/F9SjZxL/zbwJtBf54DiMdz7YeNUaXo7
mvyPt0HwKjoxZg98sXdSTLN++0JX2Rtj7ZTIqIE2bOn7aiUzgEPlc/5lOc4NAqct
LTA2CVM5ZMQxpBUU4sPEDDYd70O5J/sY1U/ytrA+Sy0LqP5H43MNVrqiTmjwDHcf
VxOci9LEVSXcteqTKjewjZE6GB99HJVgISQMK72YuMKPthXWBqXaLjH3La8d7Y96
yrk1fK9AoLktCGfPPDc3+ML12zQsVKrUexlF2RiGq1AKm6Ccx13qgibAUxhDspSn
giq9obgLzxteZZUJCyQr5SMm86MX/bRHnfSNvXZmkC/Y2+M9fszyUQREL/d6/23O
fq0d8NmxN0XXMEZ0+0ocr9q66ic0JJVCfBckFEsE1a6CqhwypFDjvHG86NlSRZ/7
0CJwKy/wUjHSAM2GYx2ox2aIWFPeoNRyIEyT1akTZP8ZqLHRtfxf/PG6Ccpxkt5R
aXACnunso9Vb+waH974d3BzBr+HNT5jaRCVHrbiGo+jtUjfkbRU1xFK9HFWrsg1Y
dis4YGOcMMct+jD3ZUKmDUaqWSV+HPTYs4U7t4c1QAkCjU51PrAy5SJMvDfPD3uP
DRlJKbsE+aoCKOjGFNtKUnXDqz7JiPSP8ZUWn14dURWwJPyafhMUi0IpUInBCziy
2bgkCUo4oYh+TGQcRha29pcWlZfDZtk+7SK033VUWBYGPbbwOH5EuJso8iPlHh46
SN9VMkjxeQTCuXYhu6cDU/4TXJAFWY6SboSasdlJwkQJmEJqQTDTdzd7GWXPrW3h
8Dgxd3+AvWXcysukJVH7bz960bP0IDf0gjW7yWtPTAVJ6I2wEM1OrxJj/PHLnuxt
AC6vkoTQXG1zqg2TquyzWTT4yb8HKiOoJiFNxB9amUtvdsN3aTZFq0tSaB8OwIS5
QeCrLTkGfA2EC1dCjdd3yiS8jjQl97aanPROeSvBsXwjicvgFUQAJypHi4lC/tYc
L3RITGveHUtjMPvTTceBQfWMQbsIowiJZtsN6EAIAO5DmCqWqDn7R/1OfqRUzl3o
xawEW2RFGlCU0XyGDygsJ1wh6mU9IcXTyZui71iF/IBpgpTNU7Cexg8e/ZyBdLqK
Lh3pIVC0n2Ey4L8OdE/0td7XEuQRJaoPmSjY5lf94ABd++Sa2YmsPUa/EU7h7UjL
HpL1WzDVK/HPti6VFVonTr46dEx0qXu0e1KehDmat/pNZwkN7q42oVMpWXjcN0bv
m/C8qVWoKVd/ENN4PVgAZJH0GNxBUpDtSYPudAxKYmkSNnyvaYp15kpJRpvk0ok5
uB/Yg7S3Z2BAB4+LKcisf0SzFxkV5NtZ7qQX8tsJL8O+bw2TgkAJae7rz8I/5r7U
T8NBKCCnGjHvbKksNZLZLpUFxtWl23liYK4U9loAPFzvcgzLjceYi4PDd88nWAZE
Hop4lgU5SdawNMW24IP1gFbhaylyPeBHWSiLFRLxV4y0PTjhQF2YED1ziJ1bKdtq
ogsg9mKSE7GJ4o20ARHO8yXR0bgIDlfYGNoRwREChREdo5r7S/eu8VOW+k2i3ww2
wl4fNALWoNZyD/dJfka9I/hKYqwdn0y+ime9+Jn/VFXrnaTmEY6jAO+a4BEsitMG
NYIC43jEVaIhTdgYMGJIKaKdjgI4aiPHxLPEfevl5CFu+SgWh6L0gTPlg6w7bkK+
BlSV0NryNH2EKKbKzdV0FnCzqj6bVhTykRAWFZAq5JpzTgt52CTy0Hh+cCIvab/8
9+gkxA5Fh633JlPuwC2pllp83pL52LFj2f9yGUVNWlhM/iwL7TUILMCx0hYXn1wp
5YHBiiYJJeLl58nDNZZyeDDrAnxyURuQMXInXQDq8QotfnjXqT7fOVbQPJMjm6qt
Fe58nCFJeBS0o4fGhmpIftNftziHWIO7wtb4tExZZigPeL+/K+5AB6XaWvrzitTk
xSFY+Wi1Qq/+6hR+bQ3CAU4ooQ516IbL8OVZpw+1VzlQfT6nvedsTJVDnTp2x5+n
UhExsQ0kZcQgq9aFOQMUQj8ItOLykimvNpAfMrgE+f/mkiSG93mGgdye2Fn2NHSj
GJYqeOvFyYsZ1p5sUX22Jm4yTCpwQ4UVNDmg21GS4rdK0J99bQjZzUVkUYZliTwi
PCKKCIiPW7B/E1vS7c4um2lPIH/2D3TDbmOwSXAJnM80VpvyMjGTrQbrzF1oAn5X
z8hkxDWZrQXv4DnvT6DkNj11XnT6NbcBMhjoSbnIN1j9ufVPmmqyX8IV5H8pwzWy
wXD9OkOpxnZxX9Unkhe6JXeztiQtBIAMUhJWJlt5Omds/u8jZecHUogP90k4Gqu5
dQ652QBrzVwovyJ3AtOISwBbgfEKetqrsj8ffEqKLOrJQ50aTCs5APS1Krxqiy8X
nLnuVjEUQuB5JxNQsmzSyk4EftrX81mnKqYl2KlISfimCAWu24dA+fITBpXavMaa
rQUXEM/hU+1K3mcdf918RER0bao3w2M/VmQpzNNjrM1fbFKG8ewg997/nMNigYy2
v8cmWm6Vv6xXZqnpj2Abl6tm2ZXOta/yEF7M79oe6zpBGwpjozs9/bY8uInW03+Q
jcbAzTVJPgRWP2erRSW+mn8jqL0RhfwJZ4Y9sMKO7lFrvRbugtn5SKnoc+5XlBb+
BFjOqg8JVkWTjnXw++OUXQ3eX5b9/IReGdtfn4VgYVNJxafAq96E4/HZyR13ZDKA
YLGGodMo0dw+ta7eYh22o8AvJ1SAXlnHUGxuEW4FxiwqvfMiGuok0eLod6IQZbcg
qWsLbNPk91a2xet3mZgl3Ltr/8MaPlikhzVBL2S8+yFiJaLXGHkWL6KJHkDC+VeG
S4PBFoR0USwKGhAlbNQTxm4tqziUvfO16KUm26Cgz1b0nOh7Z9l9hLCjyIFk3NfV
RTCNbez/Gzh70ef1vAuWzmX1tfSNdMGNVzG5KSj52efMVs4sLKl8CP7za1YGec4a
NSVpLt42zOBegsrYjHbSOAeGdmYnwHdPE++yPKnSeo6BYap62daRX6PwhUS0DVU1
CmVyJZ2pX1BMsuQHc8zQwxZQbpJG7PDALDdxvbQPS/DADISAybCTtXk8uPZYVKKu
oVmW2HO9GXrYbtiNh4QOMoMLsCyUYRFYZFD+dO3BBmkd6kp2p2k2SR3vuaIIQt5Z
j940B8fuqSfQ3G7vgwOwF7UDbS9goXQLDANc7j1DkxpoBGtofyUvkckHRoa6iJOE
Q/5S1LSB2fowDgzor5HpkyL00zykL37V1GFcJ0D8anyAABXK4VfrQD0/8M6VWgMR
iV90VTGqQr4iDyZaXf+fTLotml8o5CSVXYPS2p8PhcQbg8g5t/EVcNb7ONawnDY3
2JvLCtZwvoVbbWS6e+4eCuXPrkvSM1vXa0b5+aACvfUuWcWG4n/uK3d+JYhcxK9j
pP+AC4Ha1UZGyhNLB2D9rniJTM7DHMQ5RdSJugW9l7wdzvxjlTEPfw/UGuw1c7RS
gmAPCZmAbnSIPm11/RscFX16YQwOg8HkASRFjj/JThP2PMte8/5J/kd9BWAAOUSt
RXfE2BV4FOeluGG6Smpm7C2F4mmMl4wM4RU3+bYht7SMh82T5nrRnl7Thyx3KuTr
LM8CwkOYeWWXw/b+HviovibKZumxGzc103AMUyrYp1ZkO/ffRvA5PivN344qwrrG
83Fq1iodl+BfUGCdQhpxR7fMDZt6qpeS23vGSa5xLyY7CRePKYTa0GK78pKvxd+Y
oB0zgjycqquqox5yd5grS23q1vfcwS4VqnHR+nLIx26fU8DFfoGCGvmDh+VeHri0
c1p1fG9ARhDkJwx42bIsqJ9GjvY4ci7/MbNmk8TfqmxqW6qyL2IdUy81HeUkNIJ2
a2ZB09YHnzZqTk1iRLGTvUyOspN4/agxHADERcLMVBZaDz90VVGW27lRjdFilqyz
X3ETT0FSVTXcoXHX0pT5IZFj9sN7HZqUlhE59z6jS89qMXsVMvAmtvR6gZiCfyOE
t37gvLGWexPEWCY2eFwQE4259QotAhhX4RtZju1hm5Q/IulZDyC1sMbJs9OBr6dF
z1QLYCsvaAHgaquQ7buC8d+BR6MgxsDrs4oHePxGm5rs5wDYr2ekTsFfPf/UVQaj
61gFgFf/nZqbXU5oJXK/oSt5w/003G99rzfAHWS8TP9yRtEvybI0oNItnoI+R8E6
g7t90P02idOkyQ6UFYWCNjfaTZLw0DF+aKIeWDetM4FXnpTpwRcuJHB7KGZnrqB0
jWXdGrf0ThRx/ofy6/tpQNqdLtDsnsIR7zWXLqZVWw/T5R84TkhEfEK/Ou5o3cnS
Hi//iAntbYkWcOkTf/HzbizAtMdRuPBF7xmzmlC4aBeYUTezLIQAO7m8GOvyG40m
q/fTQzdqZdr0tQ2wy+xgtaw2YcdKq314oYJNpE601nHD96j8vfm1zrFWSmZUX7xY
+r6slmX5EuWoVsfmS8ZAry18f6uIlXD4PrzRI31jm2Vp1pk8zrpJJEDQvpzAwi59
mSZXA5JxnJTBaQMVi8rB3M57Bh7p949lmHitbNAzBIVagb4aleo0ktFw2CUsM5rR
prsstd6b+uv/St/SzrZAt8MgqaoXI0P201OCQVuF6EsYnZW4+D9g26hcQLznEVIm
pxts6J/7WwKYLm1Afpbm1o5KO4XPh0aOcTf1EPByaUq/jbsr7Q6qWBgbpNgL0j3I
LrNr7G8C8uSAAumDFkifh2iUQ4HeUYHtTzvkDqnnsYFR+TIUDLqgmtPgng9Y+r5Z
GFcshIiGodID3meB1STJnKGbkva/STJZrO0TzFhmU8XBjcnLFNgIp0C2Snqc/Nvv
V3BxMvz1fqZwgTzSMDz3lVtDhni10twIBzzsXG4g+zhp+GX+R5PZTFGZlHKGwc5h
ND0/IBOf1vmzgpZJvu/ydKqpzHi6x9AC7SEAWjmhbwHM2LXpZXaHZiE74Kj2Zwjr
aRXNRBRdj7mqlH1bJr8OEqcqTOY0hR/TE+OMSncHM+Zr8CFt22Cvq2n47+wTijA1
v37bzuQbBSek5LjLwRIzl5DyS4/01yVTUZvT57f5ktRK7d5eCGfMNfWb05k4TSLQ
tIA0qnSi1umtEr1DVmKwqf1lk3RlTkIZa8uxLAD+AoPz6cmDwRZ95wcpPsXwQgjJ
+MDjO2iwGQzIdGncu8sOIlZSk6Oz4BmDmn/OETEyiRAAC1A0OABqK0FcbrUdMjZW
RPS051ylL1L9Pjv3QwxnZm4aR65F6M1qKnc+a38d72JFJdMrjz4wUakeyQ5+q6cf
/eESlYp1IEH8BXKJ/KTYi0tKq6p9LlAYSu3vbNNJZ/4427+LuQsLEvBPsFRR0U//
LoO4jY9aTBLjZrQ/RTEswwCGGUbi+n1AD+Wt2PBVZKtClucvQNa6Uqh4Cw+lOu8U
BbLs4XtODVvMbFrZdcs6UWXTdy9Kx6Qk85rpCeZv7b/+coMvOsK0cgKNsWCk2BHu
rTVxOkLzp9Iu5pVTzdsoMT41MRZLDyqa7lgSGxb/RhXBVYzNMcRViscLztlEfn+m
tM7r13HYvc0U32bG/h5g4CpLZyXtsPFAy020ij2c+2YsvWvbojWJoMloxJcZOMT1
xBl9053vy1zMoMraIRzRn0vZJosoywL4q9auPFD97Z/+LhlJjjBWHuGbym0/QuRz
IxIzaptYucGjKJ0EUlaiGYnciEbOiytxjCtPFPzbsbW7+dZefABA4w6e9MpQcD61
eX32YTOj0CVdbkiHP8UDrm1JbpOGWfzQFU6qcuvzVTqapumOOsWF7g8g91ZQWUGp
fLJ9EaOQJzzsU7iWW/xZCQdADE9eOWBRoC1GACOd1sI8R7kgZtJq82eCK2WEc4mj
NiXRTEIEYBayL/akENyY/yBwH6gIsxo09gnYE0h3cByjieNJGtKiDWKWst35QeR1
oCfJPRAaJCDdaRmvFw39jmtd8njvW0oHZDuID6pWKukyMBci/4e7kB/MlaMhMaKn
KYBOkUx7IB9KUU2gJIRjbC4JoxxDefEMrI26ub57OJK62aUzytSLru33dFf+Pwe0
jL4Ty/z3xRL+Af4MqFw7x0KLxlCXlN64K0PBKsrFbDvifjc3OyEM/uE7u+DLJPTE
pc23kRrkOoggn1/+Ool00uVng4OeUBPydcrMrBw50z8D3PobQq9qqsZ/L2Hjj246
23MX/2cJGe2ilkkXo7NpGgSddshHPfixDxtprPLCESiKnASokRw6fimP8RGn/1FR
15MIo9WXNGIIjfDgy5fCPHEXD9r35ZsFn3Fyxcs9JXO8hxcAuq4FWVWriyoXYRZo
ajfde+FtigguPYR3zlT4nPG4v/D2i1NGGHPnH4ocyaB3Thodp3aatJ9lhRZld2xy
wHUpFRPwHjaQKlYznPHOkwY16etpyU4mhdaX9wmulYwuM5wPoYYIBbgBth2iPThI
cqBQRmwhqzzDW/m+XtIMMRGgx+EJdT8y94NQBfGiHpvZ+6zWYnemHtNwqfxxIZUe
7E3FqPVWGpuVoC5AvACCtIuqA/DuxSDcKOfomvlJdIi2U9mukka7jhfioiE3Qbka
hz57eHP3tgU3qaDbuuTr+ktjcmPZnwVIDbxmRkNgpIcpmt+16VeAT/KUhgsnqzIb
KlAQ+nJStTC1KBjt7LRV0t6jleXavnN3755TpYWIhkQqQUlAylW8rFf5T9uXP/mU
kHBU2U+s1ll56+NzRZ+6UxfzTXG7rv9tzM2uv+NJDvQvLrX6N2nzSVKdKLt6YTMx
NwLHe8+3s/gOz3t4rZsrfdIbK9d4Jsj2qSArNuFkYATpYtLM+/BbrfHnb7LLZXFR
+BMyeHd5D+gNOBjUDq+xxyMFs6fQIAO2Elm9NnHGuZMNPEccBXpdVvCi00Bnpi66
ejNeTksTMBwV+EvnJSLTb0jIBKAGPagrE/TIWY5n7fWmEr2Z73ETQbNMQNJGGE7M
KiHtjYoIRI5x/Tt4tz/QEHPnV1U0DoZBqHNTL8X0ongiX0ilDK79IheiPKYOdxNo
hazIU+QDZAMddccJRhamfdVUtRSf+aoSN69Oto0d5GCluOUHdogtFgiXmIFDmycd
UrSgyDyauU5hvrioDw1M3lkioK4+N1RfEbubTmiuOaKHM0F/fcOi5KnQg/UQWVE0
fOHOdoEUR977BOiVEepQmk1H98i0KFxpwMRgthnb1bmgaKGuwAXfMUEkXvx9uY+Y
hd9rsGgHUraBlCTwI7kEGxI+YjvYgksOrj26P8fUrsNY0lt0FQ+z5C40LkHNSCCf
EoWpQdxRGjxLh70XhWP1miATeumKdtW36RaFDHRdcvpYBuJlkicMFrO5fHXz19Y1
OCV7q5aVJ2fwN0QNETTPD5xQAMVtEEwQc5NaSWjTI99RtpzyoKdL25K+SBusS/66
nHzv4HBk+meJ5OReAIvYaXO8x3mOV7goSs+OoGmobYjpZhNtF47YwEA/azh9/cw7
ipgzGim/5TUjcqKkIuVirzusvMau3u6E0AYb0mh2JWKEAySvEKb/ZJqNbUAMkzqa
OCQP6RUugrxGn5eewkx3Rh0qwi94UYHszMj3qtmunYY5tOjEhvRRaaWv1FP9CJbB
VQBwBgwZGIEsg5qHk3OUc41YYKB8QqTpCDDifZSf8C9RLpkZvAJ90jz9hiUTToaa
N7YhlPdtZPswzq7DpoyyIVpu3yxYddZHsOBDWYh5j9uQKsqZvErEGH2Ptj6iqDzA
FpKdCGXYw8i2bZ3X5FqgFCTmy/W7TzKfOfOV+maS+CRlAZL7ztULxQxRWRuOARLY
/WiRc7YL+jvIpGroEscMrGo8kli2Wyb+TyinK7aYTvuPQBV4tIMC0QXWyrlarWxp
5r5DhyuJR88LiDNSHIZUbK+83cKOe/w7XzkGV5tMJNQdI9v9NLdz7+PpJ+biRk2r
Zp8SWQSDxeHEcaogCkogv7P9y0FeYd0aMs2JygHZ1wWc+p/X4eJRvS2LJqbHO6Mu
1YiK676GYzeyy3oAMWJMYDn2Jh+5MVMZG62HwWFQHjK8THWTYkiuJNIc272/ymCL
aKHjLBUilYAUqNixZ1wjE8l9VsSDD1f5TwdzyOsjwfmk2eOOuYHmiPfbz9NH3YGW
oaqHONdaNt4UJeUine5Eez6KGlu3V4dQUj3dH3z34cS578r4bSIGShnagILI1a4F
0L6LuKkC860KHXz6o39l1saEdARt6RFcwa3yzav6DtQ+gZnmljRY2hE443Pwjd/I
MTeQ33lX8/of4uwcX5C/mELbQ5rsKQKjmu2LkIgja1N/8cvlz+HrRORmYBE7EPot
f4QweNAbHeHqSYs+kXao4bN+T/g2mjM5A4uKPaPLnIcIzekGlxj7Qio2eTzOlnjr
+ZBYin0IfuDbgWLBLlG/CfeoWXWD+Cj/CgzHAEKk8TbrZo3pF1RIiTXlmoM9foI7
R4+R9u3EfVhHP/VnsCXb//R/ud8QbTLYVxcC4wFVmkR7noKt2aKopBgJ924xPUQp
rExDCceP9BatfutLvSIzzDFlXQ9bkyOoUKT1HYIdvPxx/WtHKvydXs+BbZuw4JCi
V12wrOhm73kEZuM5rIzrzByMqZcdDBP+QE35BfLU6SofwyL4zznKtyDyuG+oHnML
2MJYslSI/RZoTmg4yFDVo81YaxuvsLH+kGx53Uofdn/cfZN+JijtmSAOD410b4QI
uewgqk2CoG2DIvoVMSeHUHbBusNE+Xoeo51DNnyN7hyTVdQGiVrn2Hn/iqiwg5ib
nA8coTRwL2YxJv3cn9eJk5Vm9p9Gi/bwxYakmvNXZjeo/WbV1bnUK+5xkgDx2/xa
OWLjF446fxP4e6jMh9DwWRUrWYHox8rP7b/LR4OKMITMpTof4C9skYednyb2FSY0
/OP1NcK7fDZm40aaKrwB+AznQvgpGgsPxjXnTp4faig3Mct0Tg408miW4/KlTEuB
oLA7XD0D+/pKHdXWHcQv5cflXDZN1NR8yejuISNZbJYOE8+t387ITui8knTuDGzE
IgoiueUDd0snJDOFPheTio4zAHEWCdyZ8i+8UasM2QLZTGm1SA0ypo/R14gcincE
l5Wt5+Rkrm0HvNLlJfBUDVafg+JFbTYcodtxzaPNySnyDDlrAP3DenlM9V8kREOM
6rXpcJyigDZPYertp19faD52KHNTXsBhaWXdPXIgzKhMMx29cGDZF6G2dmUGVcxw
Nso41AV83Urn6ShV9ICT2xWtpRmLMqvfl8AmLpFyHnqEo6laQTqWadkBNiv00beF
rH3Xpep67PS8QLJD90xqNSnlMlfcuEgJgXQSG/dLU5Rf/6mnZNsRrld50QfLGzTV
G3eM5HFECX3WWK44mRcHx+zXxBkKghWnwYjnYIS+LPH0Zfs+zuaXwQecTRRLveUV
NqsWMhZFd2MpGkUJhIWW9BKe0z1XjBL1hFMxmlrSj5mLGl7C0TJUXvnZeVMpNJuv
oqEievaPlujSurhlmiolpVkHFZ9/fo7Gs0dXUEn8l+qMGEeIxXdkEfZ97gc4NoBb
ESP5mgFvYckSpDxluQkghgszlVg6PQnnZSc+on/PUnTI7mLV3NWoZ3cg6Mregke2
mnhlw/PYwXlmOa1rbF5jKIz0v77ea3hTOG1DeKH5DTxFK0kYFahjnXhNoiPWOF7M
LBRBKlrphNBsyetlct5UT5sA/rqDDfltgBJraJbJQ10y4J386eeqZuS5I/ybMkKC
GgYCE+aFC4dF7Jn+50tAf72UQsNf7EjIrC/s17vJ2OzieEBV9EoYrK4Bfv8c0EsQ
9PSoAKe2wBLNMUFeHhxEHhL3c7ZThywcufeRh76lIRGyCoSbKoZ0UO1zVbue24zY
UStpes6fEQfr4e3loKper9nzYP7dGnQvskvCtaVVX8yzymObc+BZLsOAHf0cNzMI
AfwJAlV+o1Ex5Az0jx3PobBZ5zZQcfxjLtk7f8AIolHsy154sGQMkCpaISb87B91
wF9GcL1he7xcCnHs++rKRsCJ1aU6s8QllQ6/ChNriK6QhtqXXzuHFcP8uBQusQ+v
pu2h9jUfCsMnIzwG7i+ot7lWBnbb9NzrCs9nPFEmSKubR3FLLThFw3n5bo2FEafo
iOhE53UxXRT3YRnp0S7nAD9jHhF0Y/qbF4goNwjNsuC6KK2PhRJAOMeUfu0Vp/Dq
Od4syG4/BuAtezH5+g5OndhmpGqrAGxtcv16oeYe6uDpJc1Hxp4EooAYBNRVN0RU
C1aF8oKuspzvhCC5T1zSmp6Ob4uWxOLJU9CjahMPjHwnrKQOZUMpHxVke8adFbtn
Er/qutv96eERRblJkeu6qhWiLTVQvG2AMITofzTVim/13YD3ujjpOuQrLz9SWoMT
jhkS3C/3yBgQTTFdQBxiuHR85GU15nrmxzEaurbEEHfKlt/9nBp/mqXl7vxac5xl
Q/Tcw6FgVit1DOvK6xAo6N8JeomKgqNq46nM567PXYzrtqQLK/UhvSJWUdx4ZSvK
CBChJbTHobJ0SL468js30oSCnJbizmXrOJPBqjuHFDxLC9OXIDXcXjrFgo3JK/Qf
A8d7xC6zdk95GKdO2x+vrGWvmwPjfktP64GyzwVBgPtY5X6CKiKJlq8MK2eQgjRH
ob9/Cp/9w3Z0XwLvt7JTAlrahioF1yMd0IngjwzEbKRLopMlmb7APueCaZE0DGf7
ZSAlpjo8wJGqkS9iJQFVcc4/22stXDr9ckiILoqNRucHj0dkJwNVFsZK/XG9/t4u
jbd0Vqf4XzninxIiah002gXdOZa3bO4og3vN0EJ9wDn17qGz3BcPO0xLHCZOjGWx
s+3CnUN9OueaQ9W2+oZxvHOomDw0EugFeywfqVFFq/fufb18vvmjqU7mEhLyUXEF
eRP0JEfdr8bU3SNvohrtDGM7mwpVMU63g1TeMWMmMh6p4y35NRdjPQwKZVSDSESO
F/+HZnR/RKiFteQBAc7BNtXGWWz2Y9PyMSAOOdfv0VRtz+vBhseI98faNieVf2o3
XYFeHqwNq8lk9DpMoLJe7egoyalc9OcbTGeCKnLnQzuLgtip9EIJ5fngjIgG9hw1
+CcRGULaqzdRujq4mK6zmkD782S9+hPOVLidUVe19435ABq6CMpi98VQPAwWuKsn
mQaxTGDaF5Mi/jnJOBJZMTIb802Hd6YsklMJPY2vpYbTMzMlibcELNhVq2/hJ7Li
UOcmtnrS8epqCDJQZqOI8QcWMOzeUVhixrW5Q1W2d4Tu9n9gASNL+/tZLox0qs6w
zGdCUkor2/Jio4sR59ZKXpfMqDPU0DyOP7clgH5Y33UDexAyxQxwSw8syq75jyBx
vZavo4zPEfBk9tauZu9SOLry6YOpBl+V3ign2aSkNMq/7pZvFyI4JGaTtyz8UWpP
TIFlf9hd1wbkkfdSWV7riFrLErS2ZUhxFIwO1dLg7tBmdKYlF2Bg69+nuvTPfeDE
9kdot9GedRDmk7aIayT9R9SmX0BvwpvNVlQlG87G8EDSUA42bRg+4N4gzD4vVrSD
pYC9qevYblnv/dno4mrWtxR6iLUXce5Kx8tizUtYQ6Qi70ZW5HF1wpzgkIBebXiV
jQ2wEfCDPTzkRiuE4Zh5R6JqlStUYbB+zSbvRA/EUnbt/kwuXWTuJ0FlyeCOn0wF
uMua3vS0vMwd0FTbdr/oKlFslL4p8FnINrsTiAHeTEicrdwlUOh8pPprf5nG9CGm
R4clciYTzTqT0wk3Mk2OZrudRzgNz8Eoj8wdQTILvzpZSYC3x5QTlvDiyanI/Eza
vRMZxR9XX+2tuIfFJW4LUrwy40CqsXPYal4vnmFvcuJ8+yABZvczIk3GBXv/VuDn
n5g928KVMwDoBYRkag3nB97Rg9XY3+GQlc5rF3Ygm7hv0I+fCDw0BWWKA/MroagL
1GD+UHkF2FdWEVyOMdUSt8pmFURle8Z5vC00PQdn2QxIjvO6ab+pVPfU0I7O8VaC
qzCQrYGfYtuMQhe96W33O30txd49rri8fftFVkTL7dbktM5vs+XuIoOd8Ifr4XNx
25viRdCZscpGA2tzRqfASc5OkSlckc3aeSkeJHOiOPzYaQm+A+LMAj3YidWJDtfd
She4t0zylfQYdsbn7YqgaPc00GVF4xTbOYnLBUuuuZEoyLzrS2vTDLzhgeAucRRr
OtauO/6DbfbPMrAfrWMq7O70y3E3BhnQ0tir3iktAh6nkVr0NeolhPA1raa2wlps
tDWlNAN2Ao4+3EKDyA+1tIHHP2Iqa1AHc+nvxEMH5cD5u3HF0SLDg5h2qZ02Ub7M
bFv+8oTNlDZIZzkbx7jHfBQr16WGipxkXXoMTukk2RTSImz8u8zk7DCBaQxnZwzB
EJg3RzJFVXkXBrvujaGfsukcnEEbHqv41QRQOQYPbvIe1KKYYrBzNAWQdkWSsFMb
bGmuzutExSF84YvJUR/rdOuSnjIhNkRRXLZqyugOyvQDcXKDJaQA1OQPnpyepAJX
iPF92XvLm7t+Z9GxRPgPSbmoelrd2FFighciD4DjqO7H+K1sGzsfUDlrWdNThyIp
Wacp3D5WPo994w7ccx+g+zao41uIq45ewxRmdrsXSivv8FYV4tBjxuqn1bRc1GM0
N2oCDu9rM3UAxinJ5qu2cvwXaE9adBL0TpW0B/KSMfF1Q5shcSYJ+Y2nRov69UIA
8aYytyDd3JnTTnj4oHxBKsRbAV0V/Tr7rYO2h8CEuWFryAd+NRxWyUf4/elPwqWE
NrAgp7pfrT7ZJcfZZTXLN9JtWo3YWQOUvBh50ppZcmr9ShCgmzAt+1KWhNl/1q/e
41dBWxM7mFMg7ktQXiKsXqgtMcxAG9bWM6+zhU3Niw2QrordN/udtJ1nT6Bf8pBf
0WdVCZ2MIRw1T7kZho79Oo4x6rcRpL84wAxuWIXdvP2sDN1ZQoQHw/xzTWXZ72z5
P1reQDKi4vm19l4GM9SPclosjlV2paUUdFrTf7yFFGE4fATfVi+8aouQE5X/yCdJ
yLQ9cdLGlqjPjTtLCltDhKip/N0gpNZ7lGv5mJktQqqOl5Zt1tlh5zI0J8jm4S9T
IEk/v/+FRGgYHVGFxat+/v1edbhAz6pPgGVHjnaASwn9JTBsz0HW8lHiIDhfBkk1
glFSnu66XIFcRq9MPw/qbZT1r5b1whmeGpKxIvSnklZz6jaa7fVgUprySpvyv1zO
2u5NizzOMoRENPgi4ObqrVEC0G2WxqIP/KGHFpy/Y5kRKLqjsw33vpqT9OE36GtW
/TMDz5XZyO2LtaQywJkVXirZrbJaWc25wWbxpnWvDc9jSZzSOSRx43hJtC55N8qO
xJllAAE6RTZhuFrOj8J7LfpOI5O2kepjzgtToURIZoSxyHpIwOm/MEmgis5JIxpT
SmoTmIU41oG4Zdba7zwRolriGCb+DIRZFDWJeo9jTDVGwVpdhEr6V7ikGgqphgXG
OpqfLJO5NXW9sbu1551O2rHvq6L0Ukdf0Z4cVf2JZJ6ZnbYkdpElzCfUFXEqPWsO
Rg+H5NDpr+YPutOViBnIgsHO0wHlFkxOLd05SWXXeplnmwN4fzgHe+2S/W9zWgx1
6vgfVAtZDoz9pmSjYDnRPUwyfGBtUvFks7e+aQaCroOVIf3NauMQp82dmf7EbByA
FZyHFj2t08jQmQgWZOX2cXGOZA4mT3cHjoOECQMPE1pgkfCqEG2TNpSzG/bezRAi
gwJOzo40ziHR/dwuQjj4cxs95ogVBQsJ/n3hWdLSUHCne9QUjmHBvC/QWQE/5JdQ
woMfA4Ls+GlGxq941a+bhDtlrohTGKrtBF9En4VeCdXdQdbRj5QR6tSsIpc6ztH8
VsUdrATaESjcVVHlvPKYj34RRHOEOK3+sz6Ee568+JOdnFvxWb36yoCnpvlAv2pp
U9ScDh+M7cBNbIFLtNL7qU7AbtZ6Xej/EAtw86rDES0xL26ECxRRycw1cB9mr1y1
J0zW7Oedj8cvCS23z/IQlVqVPUnT1QV3XlCORJwmpTVnex4K7ga4C2AsO54dL5i3
ce0hIGY0nGom6bIH+K1/RcIFxfMS/s9tcBlVSOrd9fNGCXfcntRBwxvVh0B5JAfs
eLeIY6eg4E6drFY8icQ7JQnawCDuOypuAGVsnxW42ig8c3gOUeZzRHbBPpm/V/1+
6l+6kAKbXxJ1j5gz9l1B0AH2KftGbohDGLHEgVP+EZ3F8wEYxrZR8pJ4V22x2lsv
tEMa+ShOLkru82eKfC2sFCEeJyCT6Hp9YlV0icunw4QdhqOrsYWHG0XV2FXKKhWk
JjnOLjzJFYgv0ysgY5EPfDMu7JKdMkDmvS8HNlaer55PhREmKtXXtn6EG9/6UiVi
IweFUi67NqZMS8XeH2Jjn2uxq5S9yi63patQ/KY1c5Y1sEO+iOqafHo+ADk7AatP
DJYuZhC6QCpxMdzgNgxN/tU3swIPUysJsOW6q53KIvl5igXHkCiQb2tEIYWI3IcM
PME2O/3LkZq+h3t+Kq/jzWDmT60io+ExhBTjcT6k8JfTK5a4l9F5CgDdKtk9IJP2
0yi/4RKAHnH2XU+b2ZqNWk9LXFegc6nF33MfzUWu3kxTAxZwHQwyoqBwVCSBq42n
SdYPDnG5k/124uJWkDnDh7pXImvfLWhDZkcdAJNM4PqKZgO69eHN83hMAkgVfFn4
aQGISVFxhukBDmDcmraCZILB35bAAWdMeXXkuiuuOWnTM/5bgQIrALrMwperONCu
SHw+h0RryFtgcbXVBFlNrPgals+6eJjPzB4vK0VVHdIvvBkXLAhxkh3O5ZkTdCuE
E1TNiCFtVWi3DDZBO8VAIBZ8TDzYpRaUgNwPpeLVPlYVuFdQinOpHAK10P7B2aWA
KBSbVb02or1mQUhJVJu5KMDVBml9Z/PdBL4+UfKHqkROFRpgXyKbSo+ekW5s8KY6
jV4mUZWtX7q4+G6tpvn0LSlgKql2+zCYDzzNBbu4z7G4FjmlLvPNLrYarMmqFJdI
o/2emBBobfEpeLLskxx5iXLJKhOiloxi0prNz/P/rF4H1vfZmgcGpl4bf65bPeMb
bh/W/7fBue/lgctdxlriK9mmKpQv2fXeBHZsAU6FE2+x07vFZK5PhLIc2TX4J/J5
7DYYyvOqpAn6eTd4AtwCyByHOD0wUvwP7MG0CbY69b9bVnlIbY/CIrAWNewRrjDN
czU195618rRwuxaBxT0Ad4s7PZUQbtC9W1CMr5WAp2qI7qdcrzzxMNW9juhoJDJ7
F3G25dYUEpdWxx+aCb+txAfS6K8Y7EpJSU+bftNazxPwo1+xsqJxNV5rHU9rpdSL
oXasvW7H9YWHW8oGZlEbGoVW0ankn+aAR501PWiV+PnOZXfMW6ZHy19SmRC9Oofk
Ze3ZewhMrndz3kgZBUAZg8JBCG1UFiMLGPIP8fTisgBykuxulpfFCy4SDLt3rPro
2G3COe9FXgR+OymJjeXZUeP43CVq60hZQLRXZj4qBIumgPuWvXdrr+59uTz7EoYh
1cq0sEsr9XoXNiann3WT0XAjA/TdswjqqcMwt2NkeYmZoTPdwz16e08prjNcd3Sf
5MEitwEDBB/P4/BUhKVBYmijWcTOwSvxKLjnut20CYuKXdkGaBYMK9CT9GIkkYLp
F5MKfJX+jcRXdcDeCCcnXWrH+DssJXtgLWOQSUnqQKerwRxfS920KrrwVSXofxrl
6qnrjNW9byjw7RU77vkPWE6TSVDGP0Nf/NvJGiqgLsThI1KH/Jq913mhtU2yn2ES
WNl4dg/CQjo6ktmd0xyAQSa01caikUUv6VprTMlLwTOtIv3f8kmmui/ZN8PIl+dd
71RHjDWb8WbVfoXUuzZAOH9L9o72pbytIlAD8AS1KZbBk4xygUjurRM3YfcQdTu+
JxjaflICJuzuNmGQmyazoBywTJYMYP3RUgsTY7EBGp3heXcqfDWnWZtSJjCc5neA
KXGyA+lNyqPHg0mohaiWrd4LqmzqCg7kihkt8J9XiqJNCuIiF8EiyEaOFDYS0IKf
GXSGZJMyKel39WbVRXQ5mSnZlaGaT0ixzob9XgEV0GO0v6hWsWhD00UUrZlIA8n0
y6g+CWxmo1TmEQmNwiWXl+1dgV0HnXVJ13Tm9E7jFK/WOt7ivCIT8+pQinF316zx
ffRFI01zrRDvIgNQgUIEvFMa8l8ToQQGRRGLL6zphysBFdfMQ5xfPYFguIvCamXf
XKlaDGo2I/fxeNpFBKp0sIFwgrTXYvEQwZTy0x1cv8jVvaSiO4Yf5YiamM5CCwtD
ZgmCiJZFAmSvc2pLuP+hieMmkZawzmzYLwC2Biuj2i74lyCLdPnACh9g6SKEKaeY
+YXCHTFxzi5wZZfFW19tC7dEA+8KJNsLfslWv50gJHaW6yoPKitqJtWh1Yr2Enx8
Nx24ZD2YWfUnHlR3hcYq6gZzi0AuSIUUecoOiTBcEgdJeOEGoG9fE6GuCQWRLnZF
7aifmKkQfMVqVv+PClHZOSHggK6ZBaRe2jfONZ5BbtOpAsq5hWMrcLvJmAnPMlWE
lxkooran44XqIPrD16bTaUd/xcrzcSfUxggz5fp1JBQH23cuIEMm70S2XTL5yACZ
dLqeFqzAQDZ7+GJ/aE1SfQ8Nm9LUgOzzjcBvFXOD4xIRIDz0lH745fnImG1mQ7jr
JaLubt5PkWmS/wF/zD+G65aoeeJmLAiHnXR5cS+hLQIiUToWFceol3A6MxMfATNg
HY9WP0g2XgrrSM3LYmtTw1BY9u6KVrIdgKULV6PWN6yEmVacW6nSJ9BgtRmAHkvC
Gz9jpuKO9dXep3JJluC1dptEJPeLGiXBbm7T3uiu05Qh2kmhsUTFKYvMUeeRfmsY
2G0Q/aTMJQ6N4P37ZNGNUfywBPdWRZCu5AgT1CnziL9eSm+NV+th6z/GSodTDMNt
OpQ+SHNcR1mdGp2rrtHPZDXas3Ui6VB7RPfzTipA5uWNWZrPZI7G2txsvs9Le58E
EWSqa0oPFNgveW58FX/LBwNJK/tveDc5qX7OWTuVM9P1exYT5KNjpPIR2NN/g9Mk
dF0oWgr9ViXfdk4mVXOQjId7wrKxvFHDUopNevuBPlxAQCXdvigeIACiOZm4oULY
mbeVRsGts6aE/OPynAxf5kIScOPLnxeW60ojAmKhSwu0hbJdLXxg02S/mHK9lnPl
eRsoU/JMT48d8Y92nih7AcoJVKVDGSFo3bT3Jpc6v6MzjJ3lMTrRe3DmSll2G5Wj
5MsrVBQW/9xmB/GR4guarKSPz+U1zTO9Jp/HfU5OT/yVVKKZ0TYHcAAMgPTc6uIR
l9v4bJHrddrX/tnM9AOxYk6owqYvOD0BJrszy/0xYrbRcObmFry0zxq8VcmYK/ct
w966nhEBw91OnIHu4it7G3dVPNRdAR4c2ZMCVaBwuIxBz11k6IqsMtXpvzt1tuM8
01RWncMHBJ0NfiM2/NvQnynIhqAF7tWewGQwkC55CzM6JOnJ6My2SasPC4WfI1c3
46WR0jIrRSkhnkACILGrDbBB1Or/VXADVkBsqz9AS7tmpE7SkhKTqB2gm3gi4puy
5JZnr7Eo6bz83fXuZIl+0Pt2GMBNR6OPVkbmi25z49U7+5mEtf7fSbE00c3YVqme
XI2BeE88e45IJqXXNxdWxyafpi6HksMlClQxomY/h6yqW5DKGMW+UbYngsf/V+MK
0YxpGMn1b5JTUtA0VQGfsbJLq3/oqZ6J5+LFmZfSMBFWumCajcbolN7SwDGwXmPE
pNDKi7mAY5X5NIbluFLpb7r7ay7JoJKclWp8XmDebSILxdW/TkFI9ISvH2wgLpEC
0L+xzppw1bkDcTtCBkxBzVqhDf0xdu4SqCGE1O1qUPbTv4hVjaDdAB13pHAyDNHl
nqgGKW7LURbN2JX3kmbwE89dv0kE0w4zJ/dOyiCIHiWFusS7HLkcllb/DgdEl1ax
QuqfZbqFOwUcot3MxahQypWenQB3XF0w6hRkf6MbULiwxE12+8xP9dJJOM1TIfU8
yxjNEK/QT4SHLnAtxutVQFpPpOS6efecjGQXr8stLu+SGePpkIOPkF12N3V2oh23
NJcef0VSg8+jzKqmE3agUirQLFHLPLI6ZyqodWiqFoX80yUx/B1wK9Anel7FlGzb
c96EN8pbXaVmImzqgsDt3qM3Tc/l0gyd2sVh6FQximYM8C4ASdO6LARU21QmD7N9
vSdVew3rZLSYSIZYQETswTo+c5cYFYDbBvh5B4/5mChGKgLKMjgXWxuqdn5Uja6D
r5Je1y7EdAovFUaqdo3IQyrK3tv5ijeeKcOHQGPEIVJqUS/Rlho7ppnhOmiXmqil
zjjdM4mY99ofmmOfBUqLr0dmRTv6cNc3zbJyS6dZsJASfx+BIKnmxNTZ1Rq0ONDI
urk7N9t1Gb2jgdppini5bdbbQ6zz4FZB6uiNLG8vfnE7AMiilXlv3gxPB/tQ4jLw
d1DsNLlbQnDhO+z0DVTTx0IczOCu8m2oYI0pisRfmIhoIrffnHhyvvP6xD25EAvt
NQGTxgxAJC9/qTZ4xF2DW0AZX8kEVD68eWgnAhGE8iB2pUq2X+F5NlKRyd01LtO+
HnKlLojFByOOMNT0mcxhH3Fy4hkYmgvk/gMsNfwBnYt5JfZCFlS+1+aeieuvW/7U
d9PuVD6mf0JVWtfBmBhpBLscGCg4v8qnyb2IGj7yUnai77cG+MYayoITKXTH5Krj
ubpKwsTMipB5C3M+ncP2EkLEnSIooCOObqZ9P1Fs7fiv+5WuUK96exdiPRXVaPcp
tnqJmL3MAHkD4KOT2+rOuCXENrZqcyfK8X5SmZiv83XPdeDHWtHBcK5VMFMA2qCp
uptpd6Ry02vUOUJJFo/IvZOmYAfs9NuXtNhDiBmvfA7SKQOUDgEa+1gyp+tBn4X2
/EJ8NhCdJ5Tnl3o7yGjv2jnSXQwxHa2LB0Mv9zRyMBa9u9RuqVnjdbEbLc1zXkXa
U8oz5oBemkE97Z8z4eEnAPawumM6BXW/0L2ytYE9gKtmHeUIgD/raxwsKq5+vkNS
KGNZ1AkUo9q/E1G5coekQxNOjYYkjpAGmVqdZYzVshO+UaE6scvREPneFIdV5vjj
H4Ox+xV6qv/q6ZuWjo2e0H/7IebrLzIwvryM4NIcfuue8WOOxLDmOBkgE+7o4NVr
zf6qoiBNn8uk8LkYMoPNITwsVkpEQEdhFW5NpEhyj78QOZ8PuL3n73nq1jU0FLYC
gh7UYqgemhefFEuLsmt2Y0BzNQYczcPntJPOE1RJJxuJ1zrfxgcklXJX9FcDNRYP
2ZOTRpA/Rsc9MlCDaaMsWoEPxVdCteYvOysr2LRbKEBBaoXtA+88QSEXKAYrTDq4
K9ecFVV6FixvLiOyFfUm3GkSL4jOSUBdcpTzsT5YXWL4M29CUnuoRzjwpSUzhUUk
fLEMrUqah/FgFMLLZWd8vh6+s80UHzNuFu7UzukL1HkaapthTM+7pjWV7Nfkkm0o
Tqvucd9sWUyfAhpc1opVnL4KGddbUSEJqXkRTtyurzyJCGNbE2BZP+B+CO/ygd5/
F+nV4C6M66nzGC1KyRoMF3j0XhBuS4v+RMYxmJguD2V8FJcjquxyCsCVB10z1UHM
olIskrqdQialsjaxAZRFbMVvTQhHHO1h1lGCKgU0as+mU70DFILLFnLpUiOP7RGS
oVL74rbfYb5ssFkcaaPvoD0JAW9LV1voELcQlhVRRu9Zt/KQAiUFl4c5SP3Htdxu
G+OBMOULnHT2u/WEwLmWcqE2Iyee6N6TsIwCGh+XRNe4jCi6jSWA5a4d6pBxb5mB
roqakuEIMDV6yKEwDpWET0h4vLdMkjpxrGQPNE0N1hI7RJ4RYfnUppn6vO8fXP9H
FmYPU59X0VvRjdIasdii8BaYk/cgjo7GScgqCGLLJMcBVwCJim92BSbmyvu4+BL2
TdaPG2SJs/J5hGUekqENBry3gPyG+pOVtBh1SrKvp+4+/c09yKMwDfqj6phXQfSu
/AwtC3TmdsXlMLd4hgexkI4mucr2q6Olp2VlD2l968y0r4cOMbo/OPw2SVaGfYII
t7XToAlZLT3CY9RgnBxW+afWDArmFyLtqcDjZDx1FFvCDrG+0uHnuCBsxDZQ5nRZ
t7tsTY6q+Dzmic80QBQOEGOFwohYOm2QSiu+KuBbFU7NvHsa75blMJLHppMS7A1O
BTwj/VTAxbYc5kUh80sxynudCWcX1nyO864mH0fyvd+P9ZoX+Dz9G+WrAvCg5zQ4
jHlqJMJkANM6BS3TOrskdpQ95pvgftKsq+sz7pcXeYoMfSvRhrq2AN/a+KKfta6N
u4Bt5MhprvjC4CdjPL1Fms5RtvLpWqhEpbCDKpNyJDUrIjqNs8whAhJKCGknrj/S
gflmknydpXf+d9HDbaRMS7tKnTeVW/hoKfr7SzGafi7I6NES6EcoKcM54+WgVcD9
VVbi5WQRgTH4kCl4V6K1hiZArwIiFL2WYGKxSk2RbnrZJFhJPcZt+vDL8cohXpXm
IQnjyZsov3sHpGijqV/I94h6wr+4MMI46hoBKkP7IlgpFynrubQWuqNJycuz4uoB
aXxONYjSkLQkjK3nN4S7cuu8s7XOfbJAoUcum076ohFAFu7kJYOZ8hhAxqDjtHx/
9xKs6xorq8FzKnF4/JzLkk6fe1CnUymGjg0Ll2ZUQoY7S1smstY7OqeOd8y5z3hb
RCt+ixS61+l2Jwtru7XmfJh5KaHCEkPywWd8Oj8Eet7yDGfTdOR+FseIzVEMm94a
Jelu5jJJHaD917nDvxP4P/pi6CmQyrgxmloAR5MaZexxA6tSRXuFiCE+Qer9RaB1
lJrLWEnxcYAjt3+uUx991XmvSG/zrozjfZs45T9kUY8Trq7P7zPuLp0D0jqVyDbS
1B7YLBiGBN0LjS5aWhnpGTsyJ0By6thNh4N8TMo8pvX/Q4rOpm4arcm0fbdRxWMK
5YP60RBQYG5tAfRLA2FDt6aEQwuCFR7yY7OASa692j40Eq3UQAQhT4e+F1NCDaVG
0YkOuonOFwr92Xv5LO84GhGBzthPQFWx6mc+g6CC8GSKOEsryuhk8KSyqJjuK2hr
d02YBApdjgc+bav4cU4VmZPjJ9yX/ZwpC9CW9cnpPwySU9fOWnZNjhRai0GVpddi
glm7SrfZnlpN/CfFFldxqxYXTjrb2tFL6TChGO7ym6MbH28hqls91MrlEupYCwYL
/sWcgOFTk6HIqUTB78hyMjsw3HnYa6fMfXjAIwv5asGd8yjIPig6GtrhgJs1l7fJ
VzIoQ4cnU3T7VMfVodcEo671+jKDUj9Kg83ehYS+b9Mbs24gNkS5HAqg+P+O96nG
r/kTyDG2k4Yi9amolyu+i3VRRBo5W88oCwwlwhRp578Ylr6Laim92TO0mbzhGq6U
M9EhqME8LxdM4Je/q7FKgsy1RKLcYTqXUbj2RX/Xj1vgN0gkIEA9F3iWCESCWtuR
AIfkB8dHE9xkQWhyZwy0xn+t/QnDGws/lswI9sBzAoRCJznLW242m2r/LprQ9B6f
utdXJ5YMXEW6AbLcE6cXQL9NpovgFAmsATqPMvfdnZWPoxz5dXQtaJZs500Q3UX4
1GOCPvcFR7DkrTg/MPCS1Sbbl4jb6SucvTLomrs9y20V69aRq6luqO4JQVfeWMFu
oT9Z/L8sJpl5oMMma5iB5M2ORVcEG69dLDWM8F6ZUuLSSz+VZ1XlS2cZOA/3pVO8
SlGlpDO8uWYNRYY7ZOTdD8d9k+ew82APAixbaj03Sr3fOKklig2WObUgf4Bv3Zma
yPApHrh1WnV6HYdAnmB/EAdKVbiGIBTrAPBiFRkSjxSMDjKp/3DAvl/CNnnVS1E0
1ReQ8J6kTzCdtt8kHPTjGcBeJC9V/b0xQLretSX+SubjU6SKGONZE1tu2+lQJCtA
wU+6JrxdiaTwfMvbNbyxhCNQs3PbXs5U+6mprUseqq+I+NcYSHWvoDcr2U7fc7i8
dxOiS35/QiTlMmfpZ9ubf+w0mPCmr30wbjIlylECCENSY30VPlwjWtf8jndwqB1O
J/DRvmTxQdSi0cFuVvbqhIHKvj3y7j7zGM3X90SPBc9/pWfv+LUE4/LMmSouWwke
C35r4pS6WvuXaAKrvx2ffZ/b2SwMwsl2hcz0N4p8hURnzN8PaqKF98POB9oxnzOT
IRj1+tWQKKcGJt8z98Hgu4Nm8m15aOXV6uy6lE6ZPoTp0uS5QPu5n0t2A6hQZc/0
CsGFg/zxa1V5OhZ2NjMccWPFNKLUlojpG/MBIgcB7IGi3jaErIwoZ0DAhS/gEhi8
FwO2Xw5a64ieZARnsm2QoLMGGn5th0o8UUMcfVpA7XlyPhqYWfGIOId8dPtyrmlO
uqiztU9wGrBmQejKIWsdanuWaL4RWTPFLjoTLurG5LE9mIUO4Zimu046nijXbqC3
pvw3HcGBk++j3VPCwsHPbQZQ/SFla6Wgy2XRQs46RR5EzXLsvy6e3BDnimy9QeXo
URiw1LQSrxWzKmD7Gh6cnuLjdkEaZTff3e9xAqEgZ+qmgTQaDIM2VOGd0HmRVcUa
p5XBrmCrs5xYcrUgQZHYfEZBV7jcnRRJPX+yQiHi1Cq/BBywKVLoG2Ismul88C0a
Sw6cDUupB+DPwtxF1FlYf+cJSpoPoix+yl9hGn7jCP18GU6l4zmxepzkLhZm0h5G
e7O2YUf57dkJMGcWIw07fIk9SuQeaH/G3L0jea/eBNCIOjkXVqEMphPryLIX5hsX
aNpSFrdNR+Hgx1UyczZP/Cj9LVBNYBxfCspeb05/SwC9zZQ4mr+hxkru+XGkYS8T
tyqrWCwcgdQE0bEF50puEv8dfEo3y85n+r2y4xpO+S8NPcIccLlhctphda7qyUA+
h09F2pgx8TvXCUZqXVO6Njx0wNd2LcGqOpYOatVNKGm84bg8zDqmOaoLCUhamMEj
gvw4XNTHM0SWPSeiaC2sQXRrp4Mxk6r3JRuydHv9HO9F8J68n4aeTORJMSkKtR8c
4LUXqwy5lAk+uacvJJz6h2iF/bljwIiK/eicU0MekoEHvQzfSM4lMQBqRsywaDHr
cf/mlIUKZtgPh2QZrtKG5uEVA+gnn/P9ony9qEhq5jRo/JHz6OJTy0EGpMS15H/M
cfR6sJbfiUbAQxxUfso2ectGEXmghIYc8CCh+1tqOfp7p07MMg1tHyt/SvJUATCB
iB5ogp6ZlZHpiRV650UhV3588yk/WMCdVfiVAweGS529ypJhqArDKoEnRWFjzAC2
FiHTQFLIKkXNC9nz0P7r8wQd0ZcunDfc529OoZuBG4rol2HcFGfSQER1+MFfiYzU
Grzyd0r7bJsAIGNUUpTPCs0c3lKlYvBUAhkce1C/G4HXTGBsJKXk4Ot/rLmqzCNy
4OaSRc6ZGTAs2YE8dVBt/9mhIQsxva2WzIfk8M2EkiR12ZwE98Lh8P4INu5qG5Wk
q5hHpg6L9DYOraCC8nlCnMeGzVj9INGXCFO1csrhOFoz+GBelavRFnTCtXMf1F5w
NlMvDMbsf0fCQRe7fKIpNZij7rpL3ySRSd2OyCt5z4d2La7suO82AffodxWmeljm
3KMObd+xSNf3AD4ZaxSaBy1h65cbgZ3L54z/6EMBJyV2R+6Oes7phBY+9ebjroYw
h8GcDkKKwLIffHgR2mW+t0PsRxiGCfWjdq3U21dqHq4uQgOMgcHXQxbZglsSZ6DO
G6zNeDUZ9eNzalwTCUdZZaFZeezWf/GWgPLSpv4AJyfEY1x/4IxH+FfbIvk0Q98h
7xO/XpQU1d9ay5bK3tW67poswL6YHbJzhvC33YO13Zcph+QffW2w/YFhhFcZRHSh
X/t7xkfgASoWgtpf4cscfR5o4O4hUHqn59F9Bg3UvBqc7aZHT8sssUJORXFqL2RS
yqP1TFA3Gb0lugseOjMjXSyrpB2aBaB8Djb3Xk2uhQV26pxyiAFSUKfnzNP3rjph
IrB5moMHGdMJYbsvVSS6IbMVXSj8AmuDfbrxG5k2LtJfKY0lLlLPuMVLkPznXsk0
RTOdhfW7TwxjTAcM8HnZ6hRuLic0bqPB+Ekn10r7/18pw/iuzKZNrosUIZ/XutJ2
mv+gPXIPP/iBom6y1ds/eK/Pz7yiVr+CV1JaiQriczjxyvxEUlNc+o37MUomHWIv
5bjC4xbbIFS3XFQSKBZyaywY6VsmstehMPfilkySYQaxsoJJ+G9epkBenArt5kgv
dBIrBwNXsp4+Su8npryU1v43KH+gndCA4wunz0kyES6hyfX+PWeWngM2aY+Yo4zD
Hb/0YQGYfUzNQYch2ZuTQ/k4SwJStfBoWaChtLafNs0WZZEiCKOpzowZ64cywyIm
NlSwYd5dIp6jA/Cvxt0tPM+DAYTRcyZVH+3kGmVjHiM2kwaIUuzFGE/TP58wZ4Rc
6G2DmQiZ8pon3ESOLRLc8RI+g+zuShcq2cZJqotyqUCIGo4oQV8y6zTrwBrkxIiw
j/AFwS/rMGJKqKtiuIXFKP6wn5obyv71cgrVhTqLOcPJAEvHOxALwnZ94J14MYLw
k/WMkdeagOZBjtTl6hB8ZS69CCeydH6zmLYb3OT/Yt7/gU7plLOs08R1HIuVniQI
bZNfMp+vJPSTTxlajdsjctmnCZGWLUmhpzz485Ko3cXdN/Fihy6fC7QSOKWDkgBe
KDM7euR0axVNpb4v1rUCoQVtzyXbnDD/Aa8YqpTpxFEBAjyyPxM/31LZLLiWVo4h
YcXLd2gypeSzYQjdXPP64ILMMzr4RLzLf+AF8U5BhqazTLaiBCrUAWBjJjcYV0Uk
9/c4iOC+1l0l+UVhNe0E/m6SANb+WYq048RRwKXedd6c73U39a7zoqbvRa3eIQgs
3OkGOpT02qffhrYVHjEAsH22zxBy5cI2bIcgkfduEAW50f2xIlwbWuXqMFrZOqbM
6GH+sWwAxznNjvLJl7n6CuhmabU6bvT+3fI6wHDeTetk1jqe5J84A5kmCnRy3JhD
fDiYqvtJB8oy5x8aY0XWyglvyuMqTaydluMwqBzFMKLsLtWwKE7E3oLkWrGjsiKS
JnvLAn+ooc6T8gL0aeFHXvkIlRwm6E/YULYrPY1wY8caRXFzfrOpWLF0aY2eb6j2
QRKlcYBAQ87qopOnBGFDJ/m5PmD+pRLprI1aGdyx27/QjYQsAi6nZPrh7SOF3Plu
sJT4v0O5NL7flJ7fWXmaBXTqbw6mJihncFFRz14C3kh+u1CY2wDcI9Y0XJtITuRe
cwSzF/KYulYiDhC6izQyVALnBbMZYaU0MC5oGKwx3NAvLqTDeMZ+T9KAiHt5AwcQ
HSydl8Tv2HJu4FlFcPbhZgeWg3/K+gf4z1vs8aEb2xAV6e2noCbW+gXCmnyR0LsA
CgIZ/Y4DKzV01RbRqwalX/QHtVZkjxAiniH2HOyQUFufmjds+0fESg0v7GiqKD7S
/J9AektE3R0FUwjdGSTlQDc6AHZz/PMapVh1h+g1oIjrSY4s7jzfxcxpmyGo3lyk
ywViS5FnNgjLhWFGprN64pwHyftPDXT3bNIYrdic0xnwXvzs3kYTLG+7z0J5Sh8g
ehDaXZzhr90K+AymHEZYyf0qIXKO7TJKVKq7LFIwBevMs4O9B9TLE3ui7vVDO4de
sFaqpXmgJ7mGAlaciiC6DC7C0lqWoOFGGTTrEMPS7mC0HeDiCR0x6V0tyeK5+ITA
KqhM+Bgz84ppCvLoQKEviZ5rUlYZWHN1eyQk7ho4a3oipnCjIuyEhEFbHAQXuDQO
l2/C1gYRF7Hjn5kvc+uP/MjAjzU8NqqMt/Es+uOTdF8+44Pdabc5wbD9+3zn265S
4IONEvZfduLCAYDZmIqOQKHxwlPkwc3OnIljPqsA3HqT2v6oSj8WQIoDSv7sbNma
9GqFhj4YdWPQNYINt3axdwPtfG0RZIz8yf8SuPjExM38LYabITs8QdCYs8zv/wwu
o4zzqalkKk9aiWDYf62tV/5aoOwES6YgRLuEZ/1cnMhNCFTynJuU3cGUR4EP+DW9
S2kOobnPtkChaPVjqgjIKF06RZHbGguP9WyrUob6gOd8QCMck1ggTAC/4WGPZG8S
xhlD9RA6cZquIAqFYf7H+3YuxwGPZX2M0xYxyxphcoaAkvtraQwm7Rjf1AdYORKQ
YugrNRzZWdM5Kon67NH45NbBPtwXxrob00O/wXZUUaGNvkOsQxE/HNRMQMxZTs8+
Ty3SSkGCPQQB9L+yp0/+H3PAnUCTrptV4o+WFkaX+4VZEHUkpcOQO4VNgzvA0n8G
kgL/W+puavA5J4gx3jQDDxFaJhjBhbAAEwyYfYzwZzDlKFMM3PBsplOse3JyPgop
e/iF18HYgctAPJ9LCPORwphc4RcFA+qpka0W0PAvbqidjFGcmaTieOoIezxx7JpN
0gsqBhNid65nua8yl8Biot6Ne94Js64v6Rg2Zq86NcMs2IvseVwdvpjUxN3Hc/j8
yBb9QKE66PBzPAbTMh8JuCJD2PaVyR/03vAdpj8rDXUfZM7i8RoUu1m2Yqm3QHu/
EtA0qpkgx2Ez/e01swkJTCl9j8yCNeri3k+YEF9uPXnZOo/I/VZqZ51GW3RHfJHF
UEBnzrKWmitrvxUAST0+sh2pZ0eBedhf6haL9sgaulo5ICEB2ebKYwEs45Ma0mzE
uOX4bRcwnw1zt9ZChoviiSjdB3Ra+A8TCh3QbCDWs/nExMJTJkU4pqjfdg0wO65D
/4/QKlkpD6KbG/sULAXaXqyrEmj6vBhzj5kAOvRMAA7XinNHkkLATN84xHj3ahm1
vMkaJyKU5ptCtTtTZEmhTYxjJudp1Oy+gaVZSWXe2BJD70YXnyIpSlNLzTePu/oE
BRjnFew4ezAHDBbOsmxYg8/K8wcX4ztl19RCMo7A0stVKolrkOrV7hvLLIb2xoyN
un3Qh7KZ2aqrYC2TkPGteKG1+0UytVJzCAlCFW7u9w0Bg1kOlq/cO21LJKmh7BOS
k1ESkOm8dYCI1B5ck9MR4wo/qiXszXcdoy5olQwR/4rwrrVuZC58KJo8ch4xiHXu
zUp4ZnQGjn8jF9faNMpjva7zjzIWDPlyUIRKaMUblPnWS285+Isvq+HrNHJhcwWq
dxAnWN70Nu2h/O2MqPTSpRxeGD7RBaDnfAwySEX5nTbySJT6Q9yRryP7vLwcbQ3F
mYuV+4qPIyOwecF5mbJdt8gzHZCxsszIo83QPVUcGiV4hjUa1Uj3beVsOdRjVCVy
8wOBa0B4JjsAKIMHWxHOCipAKGRh4K1uA5hMlZV3luFmMTQhcEriRRoUjXyN/4LD
vCWG6kWBpaK3PliV3JatnjSsryzaVp84COSuoIX8ydtEIRQvsVC/7ozyaguIdyTR
NV96iamAmB8+T8KMHQMZqkYNBZyumeaeLbAberWvRf4S1UtfT/ne0kDKmEkNJiFV
EBklYVbKZ/1NCR7FaZzQ7NdQKyjRDnHy5xEKqEDBcsHPSwwHDc99Oz+9etGWTNbo
g2GQq+YqOL0c6QAJxIqtRom2QIHak95dm5JlMkIGJHYXCZhSDc8xjTzblMcQUBXv
6AO+z9ocE23m5tjhbtT6yFhGmABxrUiP/BdFvCcjaAf/od5OmEzDiyEugqAI/x/o
M0v1Ld1QyvmIq2MurRKjIDrmy2XjSxgm0F85iz06X30hlVj/aVX04OlmATe8Stp8
i2LMkdqPAI0XPjFMGknwPeVDgxluxSQ7/7s8QpW9PUt+SDtCvIF5fJ/4Q5RR9LFg
Pusg/aShdrcoWHuRSCcy7tsdzczSDuCh6yA4BD8HhpMrkDvf2OE8G+56iTVlgA6u
3hlxoddou5hkW8V5EPfwo07gXmbhM0RZas0IrJMUsUSm84LAbbJvOK2OmDUzfiol
bE1fMxNAg86D5BQc2MKTv5asILxXrxBEMmn4ayH0Ce4fcGuuYlIRTNyxM64Wk657
M8mfz1H3b9abJSYNfmWtEwwF4ygI4dkVnLeYlNZ0F8xh3i1MthyiSkPvj9zttqXx
b8y4FIDJqoskrY/xvx5YuycN1KN5K0mAUemaaEoF8JB64+0rngu/V1aVyVuj8kte
w5NMrWqcpW0CMccP9RIKbgU9JwgxxOUm2AD1OiYHIqBmDUvysG7ICsYPDiflhJnz
Nx5n1bWFSjLl59Fquo2AbLTighU3ULl72Rpwhm9FyPQCbOzo27jJYFqmI90yQ4Mx
sebgbRe1tMWjsA7/TEB0revLrZaJifyOnoU02fOVDLy+SPsktMbbmG7LqATNBQK/
p7Qjhld8MgXpiW8OKH6ALe/pB1Oxk56Im2oGiGYsLDtG1F3yvb5r+3qLvSshK84L
AlgbY+f2kzdtcNGlUPfuroHZ8p6dZAlrIGp4roMdY/MShQSKwWz3iX4nWSJqJpQJ
s3Och08CKuxVdG+C3ntdPg89q59z91ckmKlNkgo0yBzKSC9heH/Mm+g9ldTYg9W2
LJnpHwZBNqguVxxHKKEQ+7GguDAGO4cDfZjizDGxX0balFM+kIUD+JCISsdZY0bp
ax/qJzyvGRdeDcZslJ9DRMif456uVYjLUnnYXZbcXtzKcfwZKSaCyMs+TnYYDTqO
0XVqwhPzgsIqBUmFZq2zNtaR2Q5JV6wzKuaDa4dQhq9zITCxMUouKD6oLR7ijCK+
mEW5QF+JQy8HmGQhDcfa21cYRvtZr1LKXQq+kOqeGNrIIbmW+GUsoSLlh6v9gUqh
y3JwqHkTYh7SENFTl9VYnaCuOClh99pMH+FN879I1UGOS+Jvoup4qenpYkzODtGc
o/Fo15DlEFHAj2v+kG+o0JBcz0fv2SLyreKvjwZ34n+XwnBzZIWSFYcZdPMX+2VK
dz6e4SYqz/jaPapdp0biGLn7joyCrZVNKrS6sW4TKKoAJxpieqs7T2o4ZH3tXAnd
KVG5+A6HJ71ubu4FRVz87T/o2+d0q5h7KNWNiTjPX2WvlvEnPWwoFkxi8DK1kRsa
jJoG+6dlqTx3GuM4AecURZhc51tJkgjZAjDPYe850A9HM5IgwsaQTYW/uV9rhw5v
DFZzLRZUFUU4afl9zK7T4MppZrpofQkelLScal+2MF1gCHMXXF2MzJGSMByODaHI
SRSMj3yoq+/u/1y3k8BNwP/Zmdgh/XMd7u3RK2Xrd+oPth77CUeeL12IxNX/shUr
4Pyq8pnjspPUPLjM3+oqSahsPA28KdMA58ZbMD6cKncukXYZWtDp1J2f9SjCuNDK
cM/KwglXzN6ZceIWEFBz1EzR7QdrT2Aolf06TnguuidANLCUFYjObnPi0Pu0JSj/
pFVt5BCodxBJiKxT2+d1T6Rcq4MdPqPJRO04Fhm3PD/tIwAHph68UQkxk9pu4fno
DaVHk40pda5Tb+yYVRW01FlmS8UO1rc9/Tbapobyzsi2cPAj+hhMQf1kv0CIKEZu
oF5OT15etDZivLcmL3hRskWuvfbyvAb+Gg9lBCkE0zyge/Z56iFTy/cxgPpXjWf+
dMZeO+NWFOcm4jv0ozNq+GinWWHUv0T8t9HopHK57OjLiiLWSA71Ypv2I1HMVhuc
o65NhKLJu/xoMmSYa6clYZNVEpF1qpnlzuJD/tce5DJ3MCp8QBEHMQvslOKz6+5+
UYCiYTuwOm7PEygT17hUP0Q/9Y/TLgTtBn5Ml8QSwSphcXeQ6TNr4TVcsPhw/hxf
iVBmoR7g+HuCgDCmqzk++DjwyaFMdE2YJSxFa3EBWg8v+uChFCg58rTqMzs/NVh1
ZxrU42i9FUahTnw/3WhEmfhqiW/uQu+94bYfH+mu2RWRe76CN3fvpoMPYquiUHzs
0ndwZJZYtNTO8QVBBdJknDOs+Zq0jTnV1TXB6QW6WPwJmCIj3urTwqWBhm9flKV6
ymcJDkQAkrhWrdZkvvqUpYpex3A797VV8a0bogQwkV0rHWiWvVvg1cdIS0HNbeUT
4KoRRF6DuPLOKlXQo6gNiD2XAwL1f+sAk5k06hgg5Sv34UFZMJ/yXn2I14/v7XS9
rtFRDrl6vZV84zpMk5nB8j3PwuYmPKMbSHhqzLqHNjfweuGc5rmb50wVwAW8e4kh
QeOQSiBdFwQiF2X2ID1fdm/f0Z4s3UdJL8LklhOB+qy2cfxtBNGMEdtPPV7ubhId
UbDL07D3AUSqh3z6D4DLTAvXjTbdq3AvJ6f5pZlCdotFgJAp1ENUDtafb4lR6R6/
5ijGP9bPzvBeIMHmPOwz9eLYpjRUvbMZgI7VKqb/mXFA1de/7AT3Uyv0T4mO3SL1
ejMHoT2KMhlSiGRpF59H4bAdWEex5pMJqucKIhsKmfiamrS1IuNq84mmYW2cYQUT
KjuJ/f6CxapFIco5zLNhxBNusRzZyZIg+clJHIdKbuiLBw82IEP0AuszEfg9UTbo
puJZsHeO5k8hwAhHJNn/1i8yLizm5AkT+GuoX6IUOt+ge67IrGEoDoLeyJNzaFqd
ujGUdSL1s15GAA/GEAy3Ab4hMnd+mdOlorjFPnGiWgeYbYxpYDwhLik6NH8oikL6
oWavmcyv6J9woi3zffaNv7glup0+i1pIhhh/lOlqvxwzCBCsZxU1lYBEQwIR5j5m
hIH4yYtsInJco0g14F6cv7wwGdH0QL60YK8qL6AELO12xXXGbplou7BFzXCpggWu
Xmxstp+0N6Q/or4X0t25OyAgpbH/flCDAFjcAegM+Kd6TFwoO+T80BlorFTcLt/h
cTyBIaygNtJ7YtchME5hdc5+vik0Z3tkfFneFdK/tUA03CoVgFoMJWvN6357PnoL
hXZdeCqZp/JPc4ppSgJmPMCWEwlvwjhMnF0K9jMIZgOTntEpJZTKrksxXN7cOmcY
pxCSeazIUjiY2dOiumHfYL5YxPKUPKFl5fvZkPa1WYq6ghpOBM6UgSCeZQUKfEGK
ZulcgS8IHPwa7JQ7BZJYYuChB17sN7t7mRmIrR8QTdbCTp6FtYHESjwrpzZaXCAy
/Dc2XB/BjAKgIskQs3YH/egRAkwBjKvTaLvYN6SLmDfrTduYQgHokg/Bc+bcftvX
+2AXzveOwwf5gdNUXqqnfckjhWKpZspTvUdpk1P533wRjH/y+oC4DSOL6vph2uB2
k7YRjQRFqcpwh/3KuyrH1BT/fcMZT7nKb9xhQPMnobkuF/qRj3Z6PRIX1lAvt/Tu
u2CRz42qHPETCy9yV22DMa/Ue1at1aEUOet7i/3CHOMZVPm0ZHt48woYS462zaay
BdGCT58V+DBJZO02+OCfgcO854zUgcB8DaTL985MPB0MmDsT7HJSqOhMvl9xT/a1
B2sAPZuP13X6BziM5Yk0Ex+R1Gq1h0dBm59gjMQDDcjesXwAfHO45ouQGDVT1qPX
LeP6oNR9iaRFEXCO+ockQG+YqtBemMBwV/q2zf3KvCs9qGUnllPU/sP/JDiFHNNx
TcuKoW6318sczMLDqFsfDsLGbbSOSOw9v37O/fK/fBY71Y6SsX6vUhlAfX7V+IQc
m4Y3QkeUcK0HZQGygq2JwAPtQbilLUBFQoOD0+bhiQ8lGNaL2R69kN8JeVeJqhOv
giaE+SOFIGtFgLdFiBA6ENuIEMmQ0E7weRq7Ha21oDTEkIZAKOSSUvxKYVAE0//w
2qKihRdLn5U7+Oewzs5H8t/ItZ22M5RjMb7tP65eGgrtQTjKmowO/dfgYvNI2Bk3
PvO/Y84HFAt4nEKpLh3zQFfeirxOC2nhlT/7gBln1MHjY2sSGJtjcviyvtNavff0
Th586t7W7cEVSotYCyh79eM/SwIatX5+f9wOuhgsB4P5uJXIYciTfXlqRElBdhCv
JZQJGV7GQodLUmj+cl46jgWSf+i60m5dM7yO2GszGQlGS0XqC5YaPMSOtpMhPbaw
IJjgrUUBVCsoR2CWM8X64kQ9kbjAipyryaNDXIImdcTL74adDXrt/5jWg5QBb3G6
gBRzdFccUTSrfnmJ8oJ2rZrMTxOz/jA3u9OZc4GiYkNc7EcUUgXyIWlxCWLgpQxN
uGJvBgcHmG/1TRbEvRepjHcojyXo+FIQlHQkj8Efq7fan0XiMvasVh3JEish7cWQ
jZz1EmrCruOLoFvT6cFTyJyPGmRQu+ldvonCoubbyJ4dtf+rk4vcuRJlk0CIFDwi
Vevkn1PfnSw/g8KJ/ipAEHDXbLYHLq0AA8uu1RTa3b2oHU2Nyy2KkzopaXGsKUgy
dcGhhS7EIApjXtLlROx9Jyuull7DWkibbaiD/ZnFFHw1au/aJ+0+w5OqeIdTj5X1
ie+mJRJFoggOqmMAJvCjxr+2tiXJDjiTtPkErowsZ4OUeuPO9QvK9DE/N+txCe4L
U22DzTwU53pV9DF/SfoJ1DAOCWc+fZwTEwnHCKDxUbkF9imoOWRU+1Z813q25rXl
ywNUhzOTNlEgaoPNUvDr9ksnowoiJWm46iKEwlcFV78sff9lF8/+KCleFmpZezXO
jZZLZVkRVNH6vLKx12YDZpg8hwiON0gkqzuFSEgHfKzRjJcMlbNJc40bHAA79lJI
x/CcUNP4RJjYKH5+X36GLv9LyWbQIMhvjQaVzVnm/psopPQesTKbVvGikF0uGVa3
8zsffjcE3apvgwDMOf9FK23y/4/LXikfIX+CAVINs/8XJUKO91NI7xV3zbU50WIV
6BI4JAhKix6ozHNGBQIh4pHLaJVvGD5CJ7RmQr4nuVSn+wMt1ygJIob8GgDCZJ2b
C3dajAq9QLZMUWNdFefinCkov8n7etFNQ+FG8cp/xcgSdv6PSshBSCeUafDDEkyS
IdbiJehTdZIz8aCcbMBUxyD2YGEomlX0rswCoPNLiOuvGCDP6GWbLAYKVIyk4x0b
wPNYtEoSLgwOd2Went/F5p5PGW51K7hn+/+0qBAav9Z76CYJ+qB+MNfWsrxVnKu1
GQYHUD9hfJjG/PcqsIgzSyC9sodRDNb4ZwtA71xPoeUG4MRBEnhBrQfPMZOQ1FZB
IPZilvISyaeKT54ViBe96N9n/+FPXigvsf+jnLbHoopR+HKBazMQy7Dq5zc3fW4d
si9Ew4IQEdsX5mKKiMgTQw67nWQc7KcDACgvY6eR65F/RKnW/dB4qAwD6QfBvaCz
Uaq6BrU3J7em/wY0rItN6ufs6fCCDNIT9sqrKnDw1NDwe4PAxkIREJYYToqNV9OC
Pyc0/kyadgrpmtIjQpRoJub+M0ZIC+cl/5XpIPrDDAXSeF8APamDkd9zNTwW+x4P
jQaYvl5M4Lo4zKKEg+FTZRXgl5TbCVj/tcNakL+sxhwpcEfbLc4JuP1n0WG7cWIu
QSX3awadERbdoM36gNeOwQgeOW0pHpZA9MXWfGp3tDLjN1Fzx3LOdZxLHlo1X44m
psYtBckMGuRdTJvHCc3BVr5GU3spKV6JWnPav6Pq0kv5VlrOWF/Marzx9GwHXdIG
tGzXVWQDUjAL5EePPX+XKqKquWlkMvC8BoNQtLtDN8ANgdlcwMGx9atQxFG4FPNn
yfOQpqFQDQT8P/6tN2hE/5IU9IyGbckKvyhI8sDuyzvLfon//C0XuDLrZWsg+TZx
K0mdsxyEJpiQfk2TTNBKyHRNL3RajveiCSAmYNpRLoSVfZ3ShbSIYSdByry9C4tg
iGj+eN2KNOk4+sGQJz+lSMX3Rg0n9/rf1sG4LSBC1WZ3RfLtWSOwmE2sGYpV978l
CY7JBYnBmAy3qpfX7YhdZe/PnTwr2xc0gfw8SzHmtc+mYb/GZCzRvqc/uGR2K8Jl
lvvMPpZEAHT++nqsu+9g9XygvJ6bYGaoxt1+ezhbmRNvuHdj6CjKHMeA6115RyjP
U37ugm9LoaXcniljbc1tpyb2HkqvFEIOBUQ4RPAPP3NWAjdN40MIpf3Bg4TvOwzA
uJ0YzMwyvsOhb3H02Z99oFlE1S9Nvueuw5BIKXFQhlriAbYGUIrFU93GafFNfVor
delKuYZDGvK/4ipmmWxovvTqIEzLoG9dSsoje/9MO5N8wkQGkggah86W9T+DT4Pj
tg7G28MORepKHf53AHLuqGDkcD4MizrotMeZtGJOoxIXljtyqqrJdhaEdyvZP3pL
bW3QO+vbVwwB9VyFKlns6GEhwAeyu6Aj7l0n6SA8yHdkya3/LShzelSoSYKWxL5x
iQZVEf52H3+oKyTeG+7mY/wfycdEKzfoCOcmONexQHhcFY1DBwKhiJSp8Kw4ZCCa
q/6hPrzhtj5vYg/nbTh1O7w101pGnQ3z3rbW72xdhdA3OWCf4NihNkPSiqgIFInT
e7DTgQWng3REIv7KoYwpAgftiem1/uFgiUNhlmZ4TIoPXIdhxzBi6tHPCbkO2suc
MUXRB+a27JAXEd5hoEcDE1wP4lwwyUvS8CfUcO8Env4BrIfD13rTgCkM9dCGnWc3
2oDc/1v1IdMtznpmT2+dBSuySXZLOCkUN792O0P5IwsdF3InnUIq1DbNUigPjn9E
Di4mgKgP9bWxDtqMdb+b3TjpDAmxra/V2lKiBCXYTWHoPKG7y4HPFoHkbUtaM6YB
mSg2+PAaqGgwpA18A/T8PRK1F62hx2egcYqzaI6ujx+2lEhU4zdgeQn6h0agtGda
uYOI8KfDpkl6CcfaMMiJvaTGtfuD2XIU16Q0wfCfPpUcWnc2VX5VzwyzGvdaAXaK
k+YU7s1xCmUsyi0NU31UJjMLW/E1yVGQnV3n/E6kYAIX0om52lI/MRi9u8vrI3xm
Yj6CVHZac3jPKegq+IRVD7qanb5GNYGk3V5qxhZAaROYo4KF/dXxHngMFuiVTg2c
WU4N9+gZOfXPO9CWX1j7+AHE0uCSzWBgdF88gDYxcFUhaLD2uGVI/S2CXBodPuG/
jrQI6/iON0wVAgTxgf+VXfJeLXA5xFYk+fv3xsqzEfnkFZ+abjHqNveQV1ZTbLJp
puf0NrSiMUOtiGUtTdaO8dB67YFtn+5BRp+LsMUyl9SiQ+0G2XXOfEycFQSBbDzf
MH9yC5CGsOJ/HKCV5LMThN6yDTz6T6h47KUpm+OBAxSPy1X1CnmqwO652yAMhFck
ecYiof43l639k/qDzY53UZgFHMGL1LsRc9A7MDo9jUlLWPa8JIpartP17TtEFXGU
ydIbtNoWcypnSP4UL7fTOMGz+qh5IoC10Q633+YYdO91VgBh1rLUbO+oh584LHe/
HUbO6MvOAPYl64QALFyLZlZu5Q2I/Mnr8OiRoN/kCoQxtVMR4x2o4uUfs4xOQZ7Z
iFNnhV8tTH65zSXF1ZHeu4rKsgaGGv0tGR1bUV0WHrZWGARKL2K8O0R6ZMprh27u
Pgz4/sFvV7zFjAL+3/8vbL/ptV6Ssj20yJKvmeHi/cah/3h3f+Reg9x+dbgj76Gk
IM9dfNolvdkFRFgJhvZ9RCPzsR/g0KRdsCYVnpTKM/yB29/gsiOS+0OpQFg1hINa
5sgQdHDXm0uMJSZjmmstckATfkVd/xPklt9R2TcrXnusu6SWGy5035hJRVOE0qpt
0uNhlP/gfdWjhR3g/g9ilgEfqu7rF1ASdB6LSRzrthIiFpzUv1/nIIUEqJDJFsfd
x1bZGzpmzYKIYOus/0kQSt/NmT50cNYBSw6l2vWDWdr8r7hEnsnx0MfxJIwWaImf
YOOCJf5ODeUno6jMT4lBP3UHlAQsENrl5BgvYdUOXNyM4pxN0IzIsc9JK086Adtk
57ZB/f571kpeJyzKp6sY1v9Mdw8Ke5XFoYvSefs2rNg7uXz4ystCfw0Wy5FXOmfx
hpqb978kgheH7w4+AcHe73ZZVux4+TAadkN44ZKnlO/1weh+BUg3Ovs7D1lrgeIj
J66oZjL76rkUynz4bhwJ77RFugWNTGMPX7h3O08AQ8YHertY5IicMqOjq05fordM
MnKv8svhcAMDYUVJq8MHoM4ySZwwQJJUldWVkEB60HQtSM9f9OrJTMACxzhTENOr
HwCCgyzk1vkfh6RbxWoynUH3jCz4tz5PRfMc008krVw6sporLLsm1E2982vUdNDW
x4Zhf63QMoNmd3vyO5iAqqFa21C+er9oUayq3r2G/ogtIXWaYCNWI3cv4y35zL+a
xsSDVzoPPcFscQGv9NnUT3ZfZdsF4fN35JDLU8E+7kLVJocT1jpsrnn2CtO+tGRi
TzcStBQ/4S7xfoTHjjSPCe8aoUNDJnRMYiGYdKiYKb4Da9dDSyhi0p8FpnSXCVHx
QGLDCT0mjbkXrC7gLolTIIWdUyIJdSJNC1OcVFqi1KZqzdWzb+xY+ep+oKVTRfvN
5KyNsFyf+TtnbZnQd4LhJdP4kKO08pji7fma6W/t3eR/7IuBO3RbtAIMBiHLmMUp
C10mdLjLynhFk6I5nrZFdXKsYKesul1P6d1RHlU8jZjbP+VWQOzk5V6WpoWlEf0E
v9OU7AxYrEXLM3gqYPZIixYsPGwl7Rx6oBdK0bj9IVf+w4p/VGVo6sNhkhZn3jjR
d3QbyyAqhYTMpsVS7zsGJfmiv67pXKxmkJX+JIc3BjrvvlNpqPEtLJ29GnBbeb3X
AoswTM4iyZq92waF7Yp4aWtu+Ytpt/Ap6I9ts6rtjcBXUImAO9VLxN8FDsWXCaJA
2zCkVeBp/E2gf+KauPeW21YrjGWSKsX4Xi9NVsDIN9DAXYGvxs0phKL2ja07Zu36
QNuQDdx5wU35gFeps5IQVEOdY5ijkDMQgFxjKFPzLapee07gsH4/CySTTfgl9ABz
Ehp82+SY8p9v7rAUhZQynz5A9q72E7EM9gr7MM4bAuxExXDtv/PFZsj2pvAWvvFL
XmiMoSJArLrdPFj7KKPrvbyD90JF0Ry6ehfY9syVosRXUUOyLNbErEeW48CxPZn3
7jM29r0qwfqdD1mbTX+VE0K1TrQGWS64D0cgHtVCVRAi9R79yr/LjR+YfNdZ6IJ8
PO5Zvz3F0+IeB0aYFM1fjlTVHA+3wK04HKQ5ytP151U21w7ZEXwJdycYrCbEJTr1
CJgpk0aR681avzk2laEj5h+Oy0Hp4GpltxQgRXp0NIwZ9FGbPOjlgmO+jkdKIOqy
y5YnNz4ww5DxnN3rPZhWcjy5XhOUR9yewzkJNSxqnU/DPaAnQ94VOfn3jcBxpQAv
RtmCXL/OpUbLDUFZ1Mu0V+e6VJ9msEpEbl0yNcIcwxEoDjMnT2iQRXhc/5CHHTsF
GzNMcLMZj76t9AGeyc++Ep94pqpsXSWVSwb1GCmulvUR98rq7gWF/kYX5HN6O2vc
bElF09C5IDugXdBhBEhwXFJePl6lj66eX5P9K5PC1p1gHAROPoFJeAXGOskQfQt9
LV/hYEV0QaIjiNWbWdzvkPKkDqDRZPDngmnsLtQZMQmsgtH4eoZuh8zU2IRMlcEo
yjZyTj+gphwI7CbIRR//6pRbxoNGupeAUlJEmFhGfhWhwWPtCwO/00E6Cf9wARP9
nZ80W+3o/1gf1ygoAJ41dgyLoWh8Zomoc9dr6sVdRY1v1rn6NRAaUJ/q3+iqpkt1
gLBShGEh/4piL1LyQqSdDXl4D16VuKmPNkKiJywv8WJr8jSM7y0SUyo4Afnxm2r5
A/MKkzYl8s4DPlz9ANUvs1wTXxFu9SSerL2wW4iRhtQLzb5RiniomOOf7qHZvux9
Tl0yAZQ+sx4FOLOQQIO8pXmYKDNa2tBy0J7ZE0aXLE/4BT+NHCLgOO8pTkgrD+hT
/k+1L1MbKqzTIVUPTecgp8RFjwUvgtYRDC5rcLhRNBSqByun5dqEgCI+joWCc+mV
/NM4gqm9EoEgphDrPhBVYeCNl8y4qHEAqctYXhEkXOstUv8qmertTn+Skbe8nbCC
UYnOeKEkOzYZvW2iNEfKmqhGhQUmj4fJUrY/or14459Fmkaxazimp/T5rKIEK59b
94GGvQWqUJHtSNVUDR/7NW/bMIOsQxUbw4o1uy1ZbLJbMoOob2+i1JGa3GtZ7ewm
ob1/2AhFsTGr5brLeHci7WKXOYPXklXO2wtxNS3RG2LrJ0Rvlz5Z5LJmplzzJiVb
/IxbB3F+trVjRCY1O9v9FZ+fZaPul7M3EkcjDewJbX4vKcaqWw7d1K7JUwy+pUtO
8jeIvxvhXcK/vID7R/Pp6SxbsGag01afO4xP5FEqd0M/HktuE2orMPabBKTZID1n
cfrH8QOo+bvNT+N0TMb30dpsNcl4cPu4A5ul6gKM9EbW0OSp5lMFKDuKCF79AaGO
GfRm7iMFJwQ76xZ4Lvb01fGQvPeRAgwnluC3jAZ03JBYlzR8ur8TS2jsdP6X5JIf
XSbvriHsPqHfOyK/LZgpcePe2bFOuApNznlRSJGYVxgmOCzIvMc+48TkYQCeUXwq
YciqdIVP1hNWvFano/LpVgnuFvw0a1VAnCKoPWstIjG+cJu5IPWdRzBMjsNRfPgU
1NpMPdmzTylLnFDJ7HXh8tuS+j44+ZWrdMZ0fd6cJ+5nhBy+NONlc572y/ThorZE
YgktH5S+06nD3+AF0GpWDQjlmHld3uqGI4HS+uXEu2QVv5e41pQi7AvoBNwXocY/
gAVi5uP0RYzd1Yb9FOaVh3ofZrxaR5nSngHaB2iKPQiaJC/1EF6DdQBUo2L1rtg1
QegH03dK+hmrrIB9nlDjHvl3jgS+aIcVkx3YEsaDRn+dYl35quJe2e1XZhEf3pgu
MaJabPO4rnxh/+zalJpst4WmDM4/YiLc2AFMxLBmuOkwDSZ7jkk3SBtDxi+wyX/9
uOeIpbpaCXbOhptoG8YDV2/FBl7UQhXdiBmd7KWs83KhZwZo7PtREO+Blv41Zpqf
QmKatuPuLFrp2xi01TwAO3s+3YnAzIQjCEgDPLxQsQPvn0NBn473Jfnso5gXTcpH
77MPYlPv8IRRyYoj4R2Fflua6/dGQzl1LOzAEFbWlJ2ALyoLYLGQKFdoNx90n5Ar
J6mLSkZIepjrEHM/8hwnA1yt5BYxxKtr+DFiytDQKh6achC12Xnla6WrqcI3Ai3e
ihG7DiuNTEmG46l7K8ifiQLtRJAiQV9c2oGBWnTZwbOREhg27nm/PXwrC//KYiXg
1TA034PzxMcdIJjKMHdO8AyfROPp7mWFLjtn1FjqxmPp+c9Ltx4w+75Kxn3npboS
Jj9seMZVz9M3p86o6+ZnQ4crOc5V+xaDOAeOXtNE8/7D6h77FiqeLKVl5IBOS5Le
aEjJNMMg7uxm0uZ+6f69MHmoz4bOsZmYp0QCSISIg5TduuJYK4YSUsqj8zyaR2LJ
oXnTcKg2gB0/ek1o9IhHOThg7u0/g5MVYLcDlGl6Ai53K3OKE2/JegOa+WzjTssP
FZmi28iiiJeunAf5qY+AzxstiFlF38cUTzgKxXjVD71rZDrtkjnw+smm9ZKSSglm
DN89JBSvOBSRlY1qArKxSPkrXoWaYsF/3y81DePdYM146ylQ9QAQbNW/7dx1yMK2
UC2u5B46dFXUfq+6oUgryxRwM/meF+L37xHwIF28YwnXaFlq8/JAOOwIZROToDaV
YsdTaNzZi6iG65aqbD96rxu6Jh+CIEdZjfOJUVkkcyRmg4+lehPUg5EeUR46yMIP
o58XnHvcLIKa2HJtMzrYb6Ig1ssfXAQP5+KH5jrfaoJEA5sSERuH3U7W7MmkhXHS
L1mZV/24jTIX2GWdAJwrXhPfiQLlQ9MziUFnhhbPsC+8npw9/t/d/mWBhqf5xdl1
3T0Erxuv1qHCL/KZq7nRb79O8St4UvT6g2SWmqleydHN3j4z3IUJHn4QRo6eZjQi
N7zGeT+6CB24s8E4wb0R5YWCcq4LcsmTuDOqhLVhE+j9fPBdsLnCHiLFTJtVtnei
6hNPbj9TayklLT53cxSKl6p90cZHfIq4IkBVn8ahyxuk1hxxhuLBhe5fRsJ3b0uZ
dW/6vzAVFNhF2PXeCCZypmvcKnLQuthtTYkRkUfWNl3jcDRUEMHHC4f6ZszxDgiM
okIDGvVUHHTCRb48AAloj9Vkkmc1Bzz/LGif4nswsHG942STlZrptr1fDZ3EuXPY
K6EZzPtrnpHiAmhxhQifFCQ4J+CNKzlGD8r6Y/3l/aWZTz2+IhSFMO+EcCDfStQ9
XWjFX0A6BSW0hhWHz2fl1cbvZ3g3J3oz9LOxWzBi/EqaETBw86bf7xK9qI2/ycpO
qatNaVnhyIUQfyBOKCuv31QmrYX6h03vTY0TPSBmGfRVK2WiVMqJXsiPlGFcRb4J
9VWVxn1AdKvLRYMOrqvjdygbatdgOtdkjoYlUlMpty/Eww14uPzcMs3JKbRmyx8F
cfR+imREx5Uhe9Mkv61kwOABxrnLzgWjqYR8qIAb84gfedSusHH1JfUeKBXFfJ4w
3d+pAM+y/QkFMveQoq3I6bZEtHNO3OlxvwOCKqhLf/KWoJngsWd33g9WBMLf9UUh
BT6bCPVGf5RJQC618IW/OV0kx2v07zKdi2kwfmiVzxYEoIzUee5xnekAfXprYmmW
EnGbJs9vbTjXMXZaFrvMzTw8S5AEvyCPDZ5goReyG+OxLhKbVLZx+TSR9ZvT5s2y
gCvIVAp4lcSNI/HQX08vujkU96wAYrFMTqKk0f/ha2FwxzjtIzyJF0CNclxWC2U8
3aLqZKkUXePVkFZOQFpL7/CkWemsc0ABQ7QMjuce61jxRWKz4u9BMLLW1mMx1rfX
tTtjgKYt/64l16WHC3LWCEDdlX00XRAdkV3H5jz/e6+tx2dMAF+P7hLblAwU5QjQ
rgbbtrarRIcLo9Fkc6QvKRhC81YRW9GqPfc8ZnWnASg1IDsvokVlMtTEIHczGgpQ
kBJbGv+yrY/OgIgWWDuc/KkNmX4gJHyOpQ5mgGFgdGkWX4mqlTkpyKsilbWU4D5k
wq/OMM0YG8pIMQ2BvUzkB5W1KoVj9LFd13NmSHFNPQ0FfE3G08Tul+sHtf9Nvs1W
34WJQTnIeAkgNJ4ulWK43aTNe/gDbS+sEcVOnHdfpsjZMFx0PRIpnPZdWrWnjfHa
t5Ki3LquhM3OtwdcMwl3J9dsIAXBoiNZADeoKTvBFHSlBpVA3iy1LVxs13PfnlQG
h3OduU62ma836+T0zWR8BG5bk3sJYDiwdf7j/L2BGUsXm21Hs8NagsWbHrvjmvrC
uvNFetmzPoQslxHyDcES6wGlLY8HE/FfPuFsagAiQWfO0QN5ESbyDVRk5/fV53SL
KjtDMo4O/Zzm+xknN6TmjYcKEWxg6TJBJ1D+qgvMwzHryI6gl83T5xsLVWcf9dsR
vGvZ27hJB8l8eocOrnRrHxaXh4fNXuQrOjw+iWMWacPbXyf/XrBA2WxBuHA4PCIw
jd1N8euuVC/ArzZyrHHGlwax1Eb7tCaVRtsFHvyFEbuC61tGPtB3wyx5hw4up8vz
BL2MGRxhKf7cyOmP9EQbZ3cIhW+8chRib7oNQoFBfIl6lSXXtk/qasHyp69OvL+a
RBVg+3WEeWY7u2K/FgLrp9k1InaiDCyybZX5A1ho9nS3ZLunxc7hIrftDXPpq21C
qFKWvbZ5wNHP9Gdoyc4ZPTGuwOIfJpDp1BH/osbNIURCPG5iHFm8IduXRbmSAFXu
Ct+IFgtULpjh+FXZb1YlY6JNw44mmn7+c6NF7vAztDV0xg7TcQccunPGNB3nIaFI
c7h8olbrfH+F5oKDmM3Ew97snT7AJSuscjAB7ArHljLdoqw3krwUBUbCTrD7QVxp
M/qECP+uEkwJRPIK3g/uZZXo3vjBGo1DwBn0f1kzGH5MXa+UXHISjRZlH7m1KC8C
VBdu8rhfzHrZx3QIlc8VmnHvTEhLrCJN4hr4vpg1GmLiCrete8BWDZuj7Q0J5vKD
Lk13WdpaR3Qfuq9FMt79NM+p426wL6Ya/TdUUrT1ztPlQkojMr83uOPPgFcTKZk6
bx6Q+zjxib3I0q6Lg68AtNSEyEj970L9FukBSmqjsayzEcScgFp/hVQ+zJdIgjhA
poBS2fWzd34eheeicsL5h2Dn12udeQHrfTmHYf5h+hQVcm4M+uXnrGPwM71NWHV3
YGpHwJu8kLX6DnmSgOp4lWLSEJ2JRZO459gnbBfuOWX8istd84Ipt3o/29ei8wUx
pA7S2hNlMZnUHhL94VqB7PqAfIQR+wfsRKN2lmYfk80R8D6OBuWWBY3nmm62ULTY
BFn/g4AJwzIMz1v5Clp9FmaiJDPr/MI4KuQbeC+jv0tWoZMkSnPEY8B2frKP3vrm
lf21/qisfMzvN1cLsg3zp5AdrJfGuZJYNYFnu1NR9NvutMIJGURuIyOzOnSyJb6k
Jh9uNWMjqxGmUzrgIgnV9WqM+FtvaYoINgKby/9Zs281tNLRBXjC7LqZ+VlIp4YT
htEGudBaPtZsxbMwYRZ8Cb7oY+4jC9F4Qvy4U0HiPpYYF550MctgggQnnpZGFf++
D6gJyTpZGpaiNeTJm2tMonrh/sB0wwbaChcHmzYroGF5MGM2avVO7JzJR9XJUyCk
LLLSExve3Qp1If45NZpV2B5l7C9ems5R4iuQJRnY7iHjhgCf0XhOdLKkZ5K2plNB
G78F3i/kP4Nm5mDd3fcySr8z5ba6WBkIIH5kMCtcJw7K8cC4dX7VKpgXggXFdu1U
bCggX9W3z0Je8ubgdrWY0HqZnIrxl5BpIVcLaq/3+S49e8OFcSWIPI7y7pbSr/+4
lYH35ItDnZ7F4wRijKJp4slqB7yIvlaWZro5+XlFGas7EROR/CVvjZsCIEoMmo5T
Gv+YiAXWtELadVdWFFpSsWZmNbYXHOV4EpqFoSMAUow3B8zuW55bjinQTuostCIf
GWh5kt2Xmff+pzCJCvgFTmh/4PNCeCTObHD8Tk5tyGkjCDI4q3Uebs57TqERZL/G
5iiNDBnUQBqknVwT4PLKlVANsiROeG8vPd6qNNCQD4r4++1z+gwfCC3F65Pt8Mzt
7coX2N9yQXYQIS/ApGOQ8BEKaaSFd61qV+k/TYrF2YHFFKEIq6AjFrhEn8CIifgM
HOSIlPjH+e/46uvANvb/WjiTTH2q/oLJ5f39n7nTUPGFoD2XncB71leXNgjQoYCN
0J8pJa9LJjLef+ODcJ+tMAatqusVtoZNG/Q9a2K8JgjPWJhI8vg3zU1NGS/rsZmV
x5mQdIBDxmIdqjVh4I7OyFdxuXDtHH4RvmdWNDc8Ga8a7J9d6qhIOFD3XdrXW7uq
z4QJd17Gj865BI3x4yd5QeHaqtAAUM3q/+wb+HBXtQxiESzjunL4vAqBqf5QveD5
sY0urtu5khuIOAdTgKYRvvKfdPnxgQo5+WyWe2Ndviu0o96JJKOjVMZcXD/kNAoD
O48MqhQzh2gO5W/oUokAhK8agO7GLQGILqMjEOJX6azQBvcTpFdR6DS+PLJkbqee
liK8EIBhQf3jsvcp9c7oHYLwbWeSZ4VhG+8U91hgL/vU8RzTYapoOo+bnppzPA4o
pzemtJwaHZBzjaL7JQSas+iO3gU/ZSnVScvij04m1uux6WeJ9Se8UaU4E0L4FEpS
okEqUnqMDoPN+di0KBE+JBvf35gWHxcld4lVKzpALLh8VT6JJznIYODMKXGnRxCk
xoilhhpLosGkLlGP1ny7SmZUsi4MMeN97KhQ8bY/y5OSw7YEO0K8fufSAnv2wjsP
aiSZ9KzES6B3wimy9BpLSKBKWxxgqSelCw/fe+NkydbqTq1TdMeYpeBrlkzT59Ai
SHaDhqb9mAiAfLAZCxA6j3IzlTBDH5S4h+LE0HaqUc/afJU/HZ7Im6ABEaQRT9Mf
7g4fhwYJd5x9jXcdDNLtYGCDeMKSUjumyt8aElVXB4abDwuf9oFSkQ0LrlKWVqYX
z3MCCIGlH3jT7n7ku1wJ/3JtDoFJMCBRc9Zl58gQFXmQ3agtm3NF+dTtHCD5tmTY
ZtU01oUPhE0EL4JLF598v8w+4QehJaBgFG3P/om5tO462/KZd9UzNVsIvmLwYnPM
YIIPMVbPXJGFVhVDo0oGRFwww47JIK4pHYD5HbwKG/Tm3SJJPmOhVUA06QeHh5GQ
UyiZADQI/ZYKTL2w6+4inM/cyDawv0v3S5ImzRZJop6eS0C00FUGY+qP2IXo1U1u
jMti+ZZt12tyAivy6sFVPNyFHAQ6yugFkBnsTNzgW8X1wdARipOWheKVt+ed1WVt
0CXGoy9d3vaTGDh3iqREPswdHcnsjnlhpELoha01/IewnN4b2t+X+xj7R5Q/bvMx
lrHrJLTBDKg66aW1P6bas5q1xBfsH/krv9HeuYl0jriLhTsP1xsf3p1LzCrrJDAi
n9r8x19Qk4gtVhKTfkNO1ENo1vSTmhtAus8ouTUOQtS++2FvMgMkxHDMwtGhyYwT
dCrpuOuyYFbn2LO3XljNmCDSs4gPpYu3+O8zxy8s3JMVk3wyAKmepcf7/3oZ7ejF
HlcyT5F2a0W0CmpFd6MQ7jJ/eh8pLCihnGOb9WCdibevX58FyglwEwZQVTf04T/L
Y2KrkiGTzkZRA7UzoGCcQ+1/fdEjU9Y5BjBfOg6BUMhJsXbl14XMpQwsyZAzSeHd
rIeRFTRyHDmKhkIaHAuEflTVUFAFgMls63qjX+AdHpBgppkPB+jO87svgF9v03YT
mlqfP/MpTOmJC46eII+F9yYMH7JmpBlZmhohdrgHUvLnGylwU4fkW6Zezt6aLSV7
3u6JrO32IgPE1cCnr0KRPbXmQiBWTSDLpMMfidQ5rKtxD1S9Hypy8qS2x3G93y4S
RSre2Jl+5uGL43NOusFoBUTAnEftetgwS5LbAaX6YJO1clkJcwian/771T3HXmNM
FP93163L/O2yYZ+eNPk6SYC9D/8nwvVYZC9BiUr+b1hdjycFOUeCijj4WcymnpCg
GS6WGGbQvVrDbf4ho48Hue17PETnhohLQ2jExdgmAqyh/o6MRVuNsK396FJv291Z
83Wjn4pWU5SY/FAa9IZ249She1+J1SFB5Ns2YAyF6dw5yhER66HPrMsv2JX/1t7V
AP8ULWpRw/E33+Oglk3F50tstAqskU0NAZHMLK3+pgBhE7JmA4uwowLK6xFbRwPA
kDUhAD37QB6M8KrN2rVkTbo8jvs3QLzR73ndOqX9siDbciZx9OQoNz7A3xa+AeWP
CddR2vw7+0cBEZUU/A3YRGXIC6xtQjpcKmsZ02qERC1Zr9FkQIWJ/vgfceBZwmPe
Yo2r5KbE71UFror+qZpoW6PG2823rON4nWvmGlzm2HGPF+nzl0eCDpTZDFOPTnlF
SOR5sRQQWAzTuC+R40h9ZmQ89Cd7vqZNGglT94VPRxQREI4tuHl9muKs7Es0mFDu
kmDAQAoVyoe/NzTjHEk8gh7lB96qdjhvKiuuS2MPSZL7JXjkQbbDfbnwNkP9hgO5
EueUY9H5r1cml8ORcfvTWCoxCpjVtEZSBwX5THBxnzVRr6a+jI/e1smUzwSCxfd1
6gJS9q93M8ids3caUEgPQpXjP9JIc6rEFdM+wby85c9dJCkwxVaGl+vx7IswwoR0
0ZGWn3Ocp0C/n+WdC3iaHXNc1zkmsqmMSDMIWEfmvtFV626M9TtQNwZSewylSBjB
aTpJqEDc4VVFTfeNG91f9NcOm8KTbCSNuwY+8PskVgl0Vx5J6/8g52biVmOoI4oa
S+Ge1sXkISjUTueD6l/Stmj55dvJdnddhzIgnPmzGWZT1jnIZ+10L/5V5zhfs4Uj
9L3mQNMt7Xr54Ocl8m2XvtWFAMO8pIF7LxMc/eWCLPK+n7JFhX1lV/DnrbesZL+n
qxdxLEdgx8FnbDWDG1JY8TjazqLm+8cR9VgIUIuxORl/k1c76CJOcHkY9jgCBcM9
TmXo3m/pnaOIZHRqUr+BOWooTvZIsECldZwAdu+gPNv1OpleeZrOB1Cm7u+To+H8
OJ0G4o2sqPi3cAwbMVmy8/OJjGPBzF1lyeTVGdyme7+sDuYYCprVdKLRNZXn5vOe
WD8rT2Wdfz7ZQDZnx1yQNHK0v6bMCMZtPWQILGi2Bpc6RFoh5vkjhhSsXM1mt940
TNfGUTo5tAmX83eS/i8KDS89JP3ATFztenveTbxyZfWeJHsqAYYBKMXmF/3BJpih
Zz0CwcPJB9FPgvXZDrqGEZWcq8YbZRP/5MSzr+jP+Rc1pF5Uw15Wrfm14+AhvVN1
MPRcItB4AqQ05VNCFtaR22yvyu5cADCo2C5geLK3csoIOY4479D9N0Wflxl6QzFU
j3A/rkNTMNDe7dngHxyAzHKcJ6yiMia7oG6k6i0I5vxpkrpsQNyATEO7/Af9r9pt
cFFIuYGFHtlVWPda76eKHJCsLXhr07cYK3AaPV/fhROGm3HaFcdKmTvecArovLCR
NbVVM1lylQ+waR9VHZAHD9Ck7m5MzvrB+VAYz1/pVIEq/zK4YNmZt9ONgGHGIWau
G+XxhXtKK2gdCdyrChV2bJz4X0iqMyH85srbd9+Z+vgobZdEIDTWk/jiBcC9LHzp
lnTO9ce1MSKKGFvlO7PimHEgBNWoCq5w9lPhEjLxmVZHQa1/2SYQ1MUitqt21wtd
wXiRqnUXgQ6TfQU6n7nWZqV6hiHohLaPQ/8QAonsVxG5efkWsckv35t/YnwUS8xa
uGU6Aj8AwyBYWqxBa0Cu6gW4Hxwh2IdUZpg7tePYuJm4tsgb+2Eg5NKscB/cGaYs
k6AJZLSgwuo1c3cakfnREFNJbWWcX6l1C84SDyMNdq5rIxcfaN7DquThuIvvuOKq
OUrsKK3xV3wo78PzFikqF3yPiyjddEJQAUkAud0jcXJsmgIAtIOVwJW6Ao5Eg2XU
G/vB9VdCCDr7pYxhzHOSk9B6gT9shNQhhhDP7i3KmosKyudHnz+eHM20fjSakw0T
+DbsJ0O7WzVoXvmfBtNPejlduKA4U+IVikuQ/eYgLygm6uqiPnuFunPFSeNFJgXf
EiMgsa+qQVk3H32GHrWeLGfBm5WomGkmKmp4ePlKwixZGDo3qsvfiPkQz7j37Crw
KEcFP8eG6wIpq8Ffm4IbaFDZQpOcM5ESsLr1lT1nzWtJHGAaRKXS9hYIkTPkWENH
2uo8frRf+UX7iAeoTUsL6KoVVPxkgsbwan1L/6w1zcvfIFEJe4bwmKkc1gQsJkHW
wdx8115n4L0VwKxDBytFzQzFk85ANhdCVyq02ZNmOCYD5Icxal80GHZVMaqtO/Av
KRKNDBx5pXBBr4tGTu+nrntgB2JI7S0dyA5hWhL1Qr1B2tAmI963H+NczoxbspnQ
ZJS0MdjTW+D1bRFAG43Rw5mA8/ltWDnhmi+RbJIya2dYUnjFcR4XduVqOjyM5pfB
A/oLl3VtjyL+lfcbQ/oy/vek/VaGPEJJDgJn2q4jDlO2zDforJ0ec1VIgPTFurFn
kqr5gYUmE4aO3cCXZBax/HAam/RYQI8Gfvt+zeNCBD/s5u/69urk+GgGFCpZG34N
EOcJPAzOEEgowTaodse9wmlTE6V4Gp30aqI1Ni+NEo7F37UJ1aetyvgIdzDzdVHM
IoFHBJZBm7P4cscHAzhTLpHhaKbiiQJjBEuLakXN3MAcwcrGKFtt7X76sn4Ht61+
j8JlrVKLgKlfSNKj3LJiUSsGaLwjyflZ8oe3+if9y2G4ixpRSluvwlxBDMmQv+sN
UfnwL1tERzgVH8XGjfIs0ExcSCSM8EsGPhHOafBkovDGhtR+KdRR8O8GWC/pjkZO
uAuw7XTFWzitEKiWaqw+I0UUEcSere5qPuz0hiASBlPv4zhDG1LrFbEcg2maXJY0
3ACTmpQW2KW+cL8+9wDcyjX6pm/T9rZ10uniErs7sCY4bpmHhXumfx2S6ylEkuO3
Ju/9NagIiXTg5RBnZQzBRFG3tBsywUn0Do7vPSQxp4geYJPI+mwYI5P8cHbhTzXX
qcWGCIefFUYisGC+EDHqAln8hYnIj76yEptbS5D6/27XaOP3OTAKY7Ggg7txVXf1
VYUju0BI0+QnE/JJPviZTE7b0WVA7k4NhtUz0qxMSOMLyf30j10HiYYMOB1Nuhn2
Yv5csGQXle7X8LYQjRtz2rb0NtBNRvIrg/Wt4a5CRXgakEhLPWGC3JRRGxKB/kqb
n6Lsrv3zT2BjiCc5YSe2NBUDYSzl3BxDM7wqt3UDYCLeG6YaUixsKZf7sFZ/JAB6
RL/fZiLnYEzl8G0a2HDGkhvRBOahaMq5dDYsiKy901jIBmXt7KoADVon0kFr+J55
Iz+La63O0Pnml3+1zcLypNAfEYGELfzK1Ms1J2xinR9MJx5nlZTvhBSEH4RWlyol
5AoHQd0Th7PL4QBeqDNN5BSmMedyrPCrA4yfyELSBinkdSxNJII5Ln8LqES62zTo
+2NZNZ3akZ9q34ORpr1KabVQOYKeFoDXDaUB/39vcoG2DsV3eZ1rzIrSC1b9ciQ0
Jsq2LfdViyVDmPSvKfReA2HfdeZ1GoU2M28goN4RJeBFCxkr+DSWSFlkeKs+1apx
lSjtV1YPPqaHGVjPTKu9mot31oxa1Bs1nio97422QLUZkbMeQQn5N9GvydmVIu46
Cs0mklU/Pj5N8EYTUwqdBouzEWQlbhStLZdpwiCQHqG3fS0w0isgXY5S4ZNQA4Dn
Fttm6pz+/6klzkOMQiS68iHX/iPtA5XJlmXF5vL/RfVI/+L4nShYjgV16vUZEEFy
8o5BkMxrjwUsUnFhE85lPUH5/3glES/Qj3r20JfgdY/pfO5qvz2h3IAguJRwH4kH
NNALI79qstZqVkRxgDwXLeIyCv8CASjYQDbpllOjbZSv0N9/UqjYMt0tPlM3GGQy
q9IULdoN+nmIajNxvfpD84Tcv92KFP4nDOyudWvbbDvC8Ibhb/cy6eygfMbmQ5WJ
CmyUb/Cb2KnudGJmpH9zkzbi5vtNyLGViDY51Vt1d7Pz5YTD6w9LxkYM8Yt6y9H8
TyCpTpNHKLQu0dDO1F/pDF5Lr/WyNHAu3YV4Ghm7YP6OpPzX4HXRBA/kzH1mmuC1
qFXq5egOvKzCpCwESFFL1SYKj6R8t0e7UL+WpZapCp+8UGEWHQL0rzpsxyVcZ+eW
cT4QRifIMne2skwbECUkP83gY9DRY6jcY91nT4SzZqn+zdX/z6rjGiJXL870svIo
yh02lJvY29wvdyVBLfG3QM7+/+IqUiMMIDlJoyp2d3Ou/yKUnrWmW5myS9XnRMw9
+D53H2T76frf3fWBUkPrV54tLKxokxfwwsGUmWFjU7kTgfNku6FlJHaeo1Uo3B5W
HwtR1PpzPwxdmSuSAdQ9A2C8smDZy3F6kBHyhSYF2MMJTPLJGyOriCZB26Jd0GOH
uiUa+ETMPpwv44DIpEwnyMKbnSiFC+A/NaxogZEG4yGXU4o9e3OSTMkRANY576Tn
VpUCDcBaO8XNCJstbAc8vFEpP/nsdtHl8+F6KcHst93b20APa/ld2K7fl1wK1SAs
MhaZewdymInX/O5E9fKO1prmg3gvLRY7AzQDMjfey4xttyegrsBEAOSbe4prJvar
5xPNPkC/nX0fz/9/ax51A2UhJxH6Mce9UVMtq1y0ud34aU5PZwbveebUMD8iqyWI
hKOSY2T2REvOdi9QFyF1XKZ/bskPQDLBpjWx7CPhuDFWU7TU+k852voOulQ0nVvP
KwcD4KpJl9+D0dBQw+Tt7tkG7jeBWJ6YUicI5UfCwbucD7kLxBSwKreb2nRJi/Fh
831x0MT8+vxbdeODn6nAfxZPaPY9lDSNh5F2oaHuiSaBj5RcifIMG2ssYnKp1NP1
eKqAUsQ1AF2QQqahsnobB73tVwHUgTab+JDN4gQz5XDdeX1p1wgg/7QsGoDQtaCW
/aGFYgUzzGTnEXZxFxWbOQcsF4Plxbf3j7jdTJaJcSVEiNwRKSzFBOweoULK0LXR
A9tgiCY0urRADo5GisGTsImXANnk7xBr//rqhResISJ5nwt4Wz0a+a+5DUfGpRhz
nvvEZdLaGG7zcJVVZMPPr1mlXzcF1mhrBX9YsuStT3cp40IfYR+PcpFLU7i9Mem5
blOB7Fo6fQKAFiq5cM2WCwUmQRRMj8gwYnDMKbumy2pNX/7TKrtFiAMLbpYk7OP/
DMSuVGT8Y2EY++twZpGCCFdtLq6iAT238OGsR+CQDR/+QIp3au0VYNOC/v4UfqEW
O7hmvPzB889ROIzqAQlao/sYDd3iewKGwwRH+pWoE1pSJbRJgUWhHjp4Oz420D9g
SZ1iQ8b+U3PXjPQafKi/+SvMhgPqAA7XdEgL8ClsLMrpyd65XCbqSvU2ElWGGSNq
QzMSulstHPO9qxMo32yujOoqf9YIAKFxHWwmD7f3nd8QeUlplvIY6S5vQF2K5fIn
B4k9VzI9NUf1UplI6q8OyzApsNCBk++nV6Kdxa/35aBHKNrmXWGXpaYW3acVBg6B
EyxyD0mKw9HhzN/0BuHfwVup1EA6ykP2rsp8v2/rmTE6q7pBPimLbTzdF5Eduqee
Js8pfdW/AmchzJgbjEZVQ4t3qgi5Rdj1QqygyyZBWfAymQn0rXsD89HUs4JEBIPa
/lPURk7iCwcXKdXnuM7QnSkepHYxlEvXCwJVjaadeGQOiYaZtHs7v1MjHB21sw8T
jVhwPAVqccXZZnPuNY8ye0i3D8P6UQVM0VUdXqy3fMqECkXd+3dhg2CAutOuHu+j
bOjhHtqEvIaz+3hcFvUm3qhFxbxkSjFBxvIVpgEgE2QprDnyodRXteCkZZVTlBna
nIrIkfL/py2NIGZhiD3EfIFw3ga6qqP8E4cPoR0bYw08uuVYc/iQ3Y6MPiSMJhVF
C/f4lZtMkfUrbFDzq9/2GfQ5fqOQwB/JlN5On35V1K6oFZUBbvzPMzuaQrLUVfMS
5KU/AouyY7Eguo6Vu9gg9Z+1QBGFJqtVS3SqMTmcvKXsc5dIoclBy6II9RCL1aQX
YAJhT3DErclMTACmGpIwXI5QwWasoS92WUUEcaLLtKYt3ZuJkOWbsaemvOls0Z3v
VYlp9ApV530CLaNkG2hFQ9IoE4PxAhxork5HZZkD6aKVqzsHUfSoyeOSGgO3nVDA
XT8hsJDKx17Fz8C6osKQ63LHr/6C9eiwIUP2GF1dSxtsdnt5O/C/OJvWDtWaterR
vz3ZIs9hCbK1SZ0tgsFqE8t7o9zJUAkyJbivY4HSddV8+4fm0Ogqvcy7p3dnJ7kh
c4W5I9ZPSeTBZorq4HPjkizyBYDL1OrlsH86xxo8XJ/08NPQ/127ro5+dJ91L0Ev
nh6fMv700B5hu2Iu6w9f1/S3gEY4HC8RH7yKTtyoQlfppikb+YiJDmRyYi0xsgPf
6go03MhSbUSxP0ebjspJRPutrN8UzkEX4AXozqjxpd/fAr4ZV9dfRCUt/TtM/Hgf
bWeoRI/zlQuZc/UsaGBqJ8sIddZ+/jXKO8yq+JiW67HpyJSXXI0M1m67BX2vHg66
BwIlM9buUlZXf/q4y/3L2n+yrzqZDrO7IfkWrNbpzQoC7nbuwlUMuNsxmH0Efch3
btIhfUvci0AaNiQditpncKElQIrdS/XtKlUc5oCp09P07KYy/fZ6Uv7lG6BDP/Sr
caeMPrL2r28B2oWYcM+E/mRC2kqqSD1lNYjMC8r3fl8FsAYv1mZkSOP+BqBn3IHA
Cugj0PFF9Pck+8eQze4lXqJz1XL6jY+LaLOHPu82esoakpZsUuApyRyaL1omxaGq
nrJqW9sIHujaXDdzO3T8shnssiCiPClrSNfyKHQhgyUCftfpIci4shujvOK01M7d
XnU/qctb4SfoOEtjJhB/ZTNamhDld3wJrtwkOB47TS6H+X3dLS57DdYciVQPrm4Z
4dLxsBwMHnsSwbWZK4gtKJjijRtsCsYLokv5ria1U5ORHH1C+V66Fim4wHj+Z5a8
RCNvA0WgZv0yFwZK/UiGKiXUUQGhDFHmDYPS2MXdntgWQo98PqzAgHBoSYKIj0W/
K/VMFIXtiKSpKwIEbgY1tzzPGPukiFjbjydBOIem7zgdF0/vZZtdU3tmB6fVbKla
gvZUJtc3nWC1H52fDJjXBO9rlqFzr8deBv3gQZZuWwYh7/KJvCgzcS5Yzm4semXB
nP7fiEs5uArIX3ZeOolIN20XQDQgNNoamtINzZ80Jx47cecbPPZHbJGKbpsvbspC
h4lmc8Pn0yitgJwGqGcL6FSCdHuyAbyFKNpUVA99C0e3E6sajGzmoNk0zRyTCbz/
KdSJ4jrDw0XnAsuyJD4OSpFOe41Mib2+QA7sdsW3EFBqlImoPN73gADbSB+8ZUD5
6DrtCG2y/rM8pP4IjQBJD2rIcRYH2Cvb20IKlvvXgzoqeJtyyIJrpfwNAEXx5fTq
0ct2IUDzNdydJ+SZQKIyDgZscIS58ePQpHcWbK+xG1mqjbcRuMdtCe2xUwGBXqr1
8DewSQx485c4Nf2POp6pvXgzRsZcXenarZsIiPeuCPUZ1NZqP2SveNCxX3yfeV41
fRVRB/FctiTQhFM+NlGUYtgjAh9Fvv+U1lg5HzoX71wAtGPdbr5QGcSdw8pDHHlv
8gCj8qZ0yF1kR97dqx0/3wuA6T/qHc4Y+d38rfHop9QL+4znbgU6KatNOdm9GIyJ
kyaP5hfCVQWzXnh9PfaqIKkf0LJRG8eJJHduQAAxEbEPuQ9ECOxPYfBxYv2FdPT0
BRiqDNi2DEPWxVvtFp5p8OQU+G9E+RqMIJZoMxgKQ94uypCj8N9tkXnBLU94M1Ep
cCrXQQBrUMX2Lm9OpeyzYOvAb9b/k/oPZo85ij4mFl1WvkzaApRR3bF0lxKZe7fR
9v9nAHSzKXo8+02hqsSf8sU9TLVEphrzdUTtAZTwdY701YiJLuyzKBN3XIlucnXl
tTRJWCg95nDV48Z/JLvap0tK/Q20o0xEZbFYayeWF7i7MqoVjm/AAqDRD36qH0kB
HadY5viUFef2AuxaWlQ4S+yCtgiYZTz2KmBCCV0euRrNCUwdgn9uUcOg7MpeEeDu
JBfjtmR+GFhxLnJfgR10PoPGPi/MYpBk2KUcQOF6J0RgcnekuFNnoA5KHWAki8az
iqONO+LUjrrXr4FZ0+ZNMpACr4DyLtAzGmj+v0Oa0SeO5ecPDAMBuXQjVomqLW00
ppJonV7hdp+F2Gxgr96EVUIDP9WUOd39pDNQ0bbNIfavmeavF6WFFe7cDUVc+h0d
HfEJgnMS7mnokRI8qB1eTSYVihIWxw4DzrgJ6x3YlD4U5/vg0BzjI/PiSVY/9s+Q
TlbI2j0/HmKTdOHEqWQtN0cVKFfZZZ0TSJdbbFT20D5hKEMiwG9/DwDXdKcUh5jr
ARCHcYBIATf7UK76eXEZdtQMFWTgSoalijddIYVSZFwPJGCMnqjk3xoaXOsW9Zbv
ZxPQYA8//dV6+WzsRbt2HItvFZWKxhffroMeKkytWnd7K0NTXaLtBJq+4mzwVVWi
tuc3lp7WRb5C0sbJlX0HhSQDuPJdRolI8LQNQ1B8SSo2/nm6z3smDi1fOyz++e4C
VHT7LkeIaBSRxw2tL0v2XttJIl8AgkUt1jn0g5NEJmsl585qI/4lTipx8h92ER4q
IhZHROZ4fyGN0ARqwiV1UyxscXO+cy0+MeN52PgA0s/OQgdqQbo/1YORwP6qXHne
kVrA/QHNSjO7pEyOcSGy1OIQWAJsl7DVFA0MPVrXpD6k2R0L0naYDMPIdCVujCar
P3cw5dLK0a6PRc1ilTTMwvPa4SdS44OSQpLdNr32wfyjHNfVWIwIv+TZ4m3Nt8Vb
Rg3kEmY6FXHMmQ12dRbc/WVZyeGMlhJWXkpG+HZC2DA0clhsBViq+qHlaRjPTZN2
WhFsCHG2t/01d0hNYd2BtEprnMemyjY+nbWp7bTA+LCDNJ9csU4uW2Un8lQsCpQp
Ts1joOqGyo9rBn7WdmGECWodK58ixPLkdfopQSZC0j6Qa13VIGe14d8boUjxFJ11
zQUTyObJ+JhaxnQ+eqD1JDhc3vgw4kRs4J1YuNvCC5sNWtg7Qod4KqYXUsY6sYeU
CZjUBmv/B/GrR/vQtw44ytQx/QEmcORlnU+BzXIxdapSkPPIly5tRWMIl3P+3plm
Z5E4hBC6ysJiUfr5WvF0oO8QBLc4OmkIBXGI3AwokJRJCSRp6R3TkLlykIYQcHn3
tluKCPjVwtvAQQ0MDwx7+/sI2NkjNdAD5ptwI/ZOzscJYC/+yISRMgQg2Ca/SPs8
AzDQ//4JJ0puVmxZC0OLshuzgds1HZcmPsOIXnDZkwUmrQ6dENqT/vNHoX6x8iEk
IpHrkfN6134VJmzT6nKbJwUfq43daedXs1loeaLf/b3J3XPJCGTaJ+IuvOyjdvgB
D0FSsusXZQpTWNNOPv1CwwhoDHlVbTyY/FiNBMwszjn+iqXRHy0vNy2zAOqQ4KEG
0pqcneV4uKlMmfals4fwzG9csKNLfQB3gU3Yy7xWk5zzE8wQu1w/2jnHfr0Mogzd
JWGlJJHmqMIUdKNaZSQn72wruFfJTfLhGq4AY+JUPRWdQdSWCxGrRDAUeNkV4rnf
5I9xAQD9ZFDmskol3D/F7bBECnLLsBflJ2MGsIaztKaotC81E/9Z21fbBWvWgwdA
SrLsyKbcx2qXgD/0V7VQK16iO0H9N6sEsvV7jeMqm2fq/qNd0RFQX4mcXT3VCm+g
HIPeVgq7e4XclyHBOwkCGnHrxSgbAo537XXAFkoOxmdy+pPtIOSBPuCCb02Sr5dQ
bjSuvVOtFC0vUAV2ygB0y/ksZfLIBHWUW0xgp4ItX1ZWWKHBeHkC/0RBMvZcJlZS
fmof+m7mEAAReMnwdp9JHpTJKDOplKVbfZLFz1k727tDmDNWg5dw69OLmclsmwyK
V+NB4oaRf8yYUAvoYhfrbN2fHLNYwxitXBrQBmjTfTSDZoikEVtaP7cEj320ppyP
HXK0guUamwHTecysrL5e14pNZ5HqqjahILL9LtCfMwlBQXfIPswPYa7Zy83Si4Li
hXLViGgPnEo8os4rHKCAcJBR1YJFbO2cUXoMvV9riVbkS7d2pGLOFrKTORAVIswe
Pn3vu2kWGlWzJzoGsuPIxfZCA8AOuKXX2y18suPiORQNm73aEOXckbNo7GJ7tYZw
OGt8ireNOkXKeMby9go/7554eLuH5ENh+94kBhocRFgFpK37/4Iu3fOKUhpIPSSI
LaQA4dQ1tATJrj0ZVQYesdhIBi0wqrYaomvItAEXZGd2/1U+hFMe5YqJyydFtEBd
uj3KWfdtdB28RHWfj/94x1EtxPVKQYAzIxrd3PKPpuMIBazzRIJyV16QgbUzL2+U
H9C90cbmtXAIi0GbMsS52CWSIQIhypgKYicl4bDc3tCFx1OBvwcyS082LavwxZ6t
GtC7fwi8W+dMaIwQAg5Vic7z5pJHDpe1It+Bmrf/EFsJKAgbUq/TMozYQ7Pj5RRM
eU+0KPHUeF7QyY3w0RBMjfUlluheQUsqdP5r5Dt0Pvy+aiT5bi5w7jDfmsoWIlhf
lGKUY45lFUUoI3LY8RbaqPs7SNX5dBVGsb51HVCHP9EH0MfBsC0SAG3vU/RdpXLW
F4wedxOqPXoRTWQHLLsEkxPsDpj6DK4G+jkJzl+f2yMw/BsyucVQPUrvmCypvA87
Pj554oBoJv0Er77+ylqBDKwGHiYVKkXVUK0YEIfDenW/BGYud8dpInpM03i+UVDV
LuF1w625/Fgg19XRlX3PXIfKXxifRzFHio0YwCBf4iE2YmU9kAgydCzoNe4Py0R2
aG6nQ3XpbIYzNzqXFKM5S39ARqJFSF1hzaNmh0mDqAq+2ix1gLSEtj9E7ChSOPBl
oi6B+I/E3hbG8326LXKJf4uqZmN/BnB3784TnmE7rlKSQ95pzu4XfzvrcLRm09Vx
YdTKa2lNSfCMcQ88K8hXhFJVzL6oj9JV4V1QlFRtakRYKVNON5AgbZLZgu/HeYID
6L7yer4GtmmZRD3fK0pS0HNJgAz/EVEn4LBfisGuXVVpcnDvATgK5B/xtrMNttLa
95U1gOusujeMkbM7/92PxQElcpCjt4dFASGiXawoOhc/vR1mOBTJ8UF+UF00L2er
Vsh2SmGY+ty8k8rRaRaCFaJURUls8nIl3vqF2UeIjf/w4s2BTRpmGhT+1NHOrJLV
tEstf/yVT9OEokqDKZSD4aeP5YD2DAgKoW3M44oVLJZzxvXnNWAofyFrfC3/NkFo
q2iLtQKx/l7ipKtq1c3YlsR+GpzoJgBY5r3x8eCAfVHBmGGqgnOnuHnd00UHOlvq
dhuAqffbc3ZTe2Ka+TiAObLpq5EB04Sr0XQ14kh0xNBj9VsQ6LyUsQ5/Ua+z3yYV
7qc+fdqVRMZqfdF6wtKGWL5j/boDR2N5h+9+uUDF/9RGtDbsUSf0hXa87+K9+ABy
VtwPj6ZGC6/74aGwRGVBY1zZ36Cs79VJrtgJwzdOVxhqgcWrZvknjgigB6qY4Twg
rECndgAKR1jDfqKhUpEKzARSrcaLE3PHiMn/Rm6Hv6Sp4UdKCuS3MSUxoL6jrf5B
/wOKS16i+qMMwchOxU6HLE+fgb0Y5dXNlZ+5ZzL4AiYDnwh26dC2LM+EK9keaOY7
UmMdtXW4enFuNjbsfs610+Dl4QUBDTl8+T3mTHPAMD032JkpLmYYimUMyGClpMKc
9eAOwg0vE3gqN4+xfi5+qjc1e177LnkH5Y70gedP5IJHVJ3PXYf6F5Oc4S3gbnY4
+QP0L8U2tKeBWrdfP1uFHmkZ4NbG3do2BRf6skun6/o3VzrtCzIxuhi5rK9FMeWB
I0O3yGEtjwthqEQwiNDPFrDeA2wFqV5yQ36r9FjMAVX7YdeBO9BhacxFqXh/AKBc
SvcOjMJfIzdPMPUakTVQsJSeLtB08nQexFxOntrg/DvztcoxTlv9S1tv14AmDO2B
XRgGbitCreaqD0eGXAjjALsizlEiajCMomTcZzAglXZWRxrYtwF3CgFNvWhZPpc2
ZOc+MOpx1mKJPcpel1YVa4/1hMQYHDlFP837pYpGCNcAvkVZ74bEZQ5Q4u14Q/gO
kObqZVPLc5Fc3wOTbXHqC30ZcJalWLFsnnHrkP7EXISziF/+4cqG2eCtTwN/vZGd
SPtC3FaEsp1ZnEhfQUXTqT+ne079uJ3miK/XDISuUpFcHpSo4cLBLWDvoAt9YtBM
w6kah1saXMz7rd73Z+hJoH9ij7GT8Vj3REa4FMxjlcRCUBX1xN8dYnV4dpUsctSl
UpjB+Y/ZVgv3+TQrIRcSGprSrCo/gKtQ5AneQR0RAOa7MMqxJeXMRs1YC1KeGdLq
d3I7VU3OFKB4r3DQqJTspsKJXbKPa2vqTyi8ZoyE7nn6ed/4ozpw38rhyJ6Py6qh
nONYoOPAFEThvqTfl8huHjvrN4wGWNBLyFGfvYT6rOeb5ekS2EXqCMulAezE3uXC
80vscv5G4JSLATwaBx2qsop4VLSocnVCGCn0FQQHw9FCpXp8udV4+28gERxmT++L
e5hbXSenpDNFAn3aOTkpTYNZzBNtCbgoq8m3kExoOdgG9uUG2JLU7ZgR21TdxlCT
ufCkQZiYyJ+qP0DBtkEkLnew1leEVToxTm8Pv65uVnuRCLJ6O2+EDBfwiMUP2h7/
PH5L1KlugVRbQpocczpJd2CMAiOtHTdvHehxltOPIxAw50v7mObgjENEELd90K/r
Bt/qslkUehF54zgRrqvlXdI5hdNBr/x/raOIVTXgqZDiYZ7zdQrMoJBGPo03FbRu
9YLaRHjh+pF2IGCJaKDzM07nVZVxXE1w8bEyAbeRbSsBaN10QN7qKB353Rj7R2mS
+4M1/cfriIYgIfH8Wx3LMG4P2SW3bqhuY9J7lYQ8GxIlQWnoe+suZV2i+KY/LFPF
XVWynsi5J7gUh2Y1d1GWVZ6Qucgf7lbUJ5Ia3fS+74ZovdEh9MTukGKX3OiIebIL
kTh30XCJMxcN3JJsyRPiEHGfKlM5NctbstrO/zkfyYyDok5da5nU4mCRIFoNhxSj
S2sRdo6qXdHDdhssAZdFPgiITJvHUgRYV0/MQRh18Ti1ceIPcltz+Wqji7Z0VpNk
ZkXNweCFMHyFHISxxt+ZQZy1vQlLTO3nXqHz1kJiya7f05Cm729YIHwtnuSPPWnW
RvuoZ136gRlpS+j0/OErAWatK3H/ikYF7DPFKpWEjnUHXxLLi/iSBSBxtDKjFnPf
51xQF6ZnWTo7NiUc+i4xUQ2OljAJlF+cntm9SN7xZ524nsp2db+fBYgGCNuhFWlr
n3fntwYPgMP1VLNQ7Njvy4/La9isA9Ac3zkTxkln4dwkPuXHUAJZTbDR+FoclfuY
wUQ+g9Wfu2w8Dq7gG2vVN4tFoJaT/pyfcyKxnAA3Ks3yPX+MP55vwdqaOmMo7gxT
I0+oVtsQeOQiXuMDCKiN64U699L4VeeGnUiGBbtLjYGieYlH3QJnyaVtwOY2I6xG
sW0GG/XoWtRBHZ7uMUcOjZbw7CUlgs1DW9IGzrt1yR5c2Rrgdfw0eMafrN7d3UCY
j4jusGb/QzALbZMHzgSqhFgRKxTlY4w+YabwkjjNAcfX1bcblD1YFkyeRfmJkITq
d0Zst1q4zb437I+ZXM0k7+7VIyjZJWeWRQm3gch0h2vh01hyy1aBGVWrgI3cfF4E
VOLd5rFNFIHfHUge352zfc9SBokw5gukE5cLcfHjYvfswMkLbpZaObt3qJOLHRxn
7X7oJy5fSKbQKCQfZ4QCliXgu9ZWaMCXa4Bv4uQZ8t5h2z7QJaLtipy/o4Vytjuh
oSlz+NkW1FIUdsCq2ceSQ5c4yQrXU4tLlq46JB0wH4f977o3q4J5OwY1f7gKNIWW
jqHE5peEVlEFsfG+QcaWUdOJwUiwGOjzbQvx1GWTTg0oYLuvTj5LQLvVRqrmvLF9
O6/+ERmlkODMPorWnXGsPC8g0hFmkPvzI6o8G/QD1ZOZj/gky285vMWE9ajT2dLD
lMGwQsuGIDTDOpzEd9Ia1vXaldy9sVCIlF8ze1eppbcNSrEUXr8OlQI5WR1at/Nr
uEur8G4R3qbi/AMrjmouqdOMODkQDfvdyUwGbl5Xz07ATCpgCe0gz/XhwqfoQXd+
uOCRTwRNIQ4DHVPn+L01lGXTbw7cICwiaC8Sw+OIEr2nNVWwZmooI0pTNygJAqkj
EDdufYwIoQtyyJ61eHYIQyTly5mk0YHtV+oESy01TYPYU4Wtmb0Fj18uV/VfmiLO
Zl4Wf8Po20a5XR4V/GZSgkqtiPviChaWB2JiQWYxwQMTkSiOzGDMbmXYvaAozPjj
IGA7H6ptnGnvPBoM3LBjKph/7v4Ra7rNbGETMEYADYW3zS+8bIpXkdB589JlJhVQ
hmF4UjvBvClErSi5cYAOtqj6ZItJEPIQ6aOEssTQ0YPfvHTMgugn/U65Px8kjVnM
aLXnYdr6CWyBaqKKLuj8594nIEDdIAZ2giipIOfX9xNozK5xnGoZSN+5y7TLPZSu
ZYyfzrGN96wLgSB0b7B9yWVs4lp/SddjJz0UcfzFT6IlWZrlgAjPnSgQccCyypHT
m8R9kgSojIpEDmuzDv1lHidwSMunoEetY8pktPTbHIxl6aqz2nH7zxnysb1yAIwn
zQCvSX82kqiu4Ke8OKEPXXckldHem+pgMblRmgCR5veRY5pjBsEWgBT9InLxYKJO
vfBpiFsb0J0nc50udV9iNUm0OA0PT+9Cc/5HfBdfsgJLEaE6Im9xCsAtuIuv0PPl
CmofP+1NVrTWqdeVxJ7v2oxcWBG1Ene4CyG7Rjel8U5TmJSpe1J644BIYpjugrfU
2W9r2QcjX2CsFsk7nphqU2WFc/WwqJLvDtVSijvY3kmdVh8u95/x8tlzab8s0g//
xRJPZMDOuPOhrUwESP0TyqQYUFx+GoDf/VuKT02fMzGkk4pWacFAkTrx1VT5NASf
xaAg7MN8SkeG9nZZ49QZ/RJ4VG+N9Dm4dgO49XPf4CNUq5xi7cD+a6335Zwb5k2o
kCWkCbR7pMDMUHN/31eTqE2JOkHPsdnLIXRFc+AooZLM37Xh66YQzE7pk3hzPP1F
rS+E12BmEH7xJkAbcBSBlpOAkwFDJ8aODNdvJ6Sp1wdTklXQDBpsuPxepH6/u6q7
APWddhEWDNrSHPhvRIedHgcQnha3KI1Fm37+GiIZNDNd+FUdmmQMz3RP5tlcAIq/
gvjIDVok7/Qj9k6VSDQrGtQbuQF8gmgvay1uMX2pH1frUxyRxz2SWaTlaofEp/5l
ODzegxCmexgIEe0ZZvW08nlUU61NGMxaCqIYfvcBxxfXx1LjcZGgkz5TvKkoq1X6
gwKlvxezdCw7inCxCqIqfXRX9aZ72od7ZrZH0mMulJihgbnJw3S/eAti/0je5qW8
rSKUhk4ZKF4xQ7lh+7ijPJMA4AnlBohPbPN7kVjVWcFg7/7gswPHduIUGPqiqVuS
i/ugMWEPtMLmtBRdlmwhTlMzPV8W1qzdz7uBWvxbXxnxwUQxmSEpb+wJbbtYNzv6
LfqdYCdT/eHZ7nz45ycdxEQFbu2xMhp4kAwOcREtXz4jzQNeuS6xQiIENqgXBmBX
NkDTXLRZgknVpmDiRn/E/ros7fPE4+AEUbB381qx/BnJOtjx/yj64TniT4W8CKps
yN2DJF3cupunwszCemsOGuVD5smTpCFI7K4ZNv9vpmG2AKxcJo42Hwzs5SZk+yMl
BVAMTjSQBmWIl+dBQNkwvpuaEZeq4E79I2twFgSvaBCCEcl6WTmoBu+D0dOohQBM
9D/gY8CCul8b0LHgOrtSyDZ9mofm5dILAf1I39q6AshBJ6sMf/evIgBjAqMGZTKL
QlmOmQoKomoEJ87zt/Q5pBmLh7NLsdVvHTxbJe8DrGX/hs81qxPV9ByT08SBHkNX
bSMbyhjytukGQOSRsiYdFACu+lV6xnPkbbqSOIcFUkxGSN6l8hc++lqGehKeV4yI
jlQTOWdagrzrlUzpGOyiJR97ZBYiDci1YDBUN3YrtXSeg3BZFNc4JNIIZ6tbKxYY
9YV3erBB+FITBoTxB4V/jJHpklbhYAjA0dn5jq3ctkzJ6U+fIXvQxKpD+OBuQubW
q1QQrooat3RNZZZ6Q//7IEsVaPYyeAKSGD9Yah8JNXLYVw8m2mdroKYHVjJ745oc
rlOyWsqsfAS6cr89c1dFfvTww1dGiOzeD95ICki7R9jJQIXfJaeQCLW0C43eB9wN
SWZlcFLVOX2vw092YWEEkLYNt7ynjjoBEOYvs/MyxMLXRpQcUZiloEqHx7l9B+Bc
aV6DZCDVYCP1/zNWnEXD3BfpYNRBPWwIK7/AWRmJklqrvXnF8OsIo3rwM/+QykWp
WBY/7lRL2er19irO1zn5Fpq4mpaEi63OSLc5J0PnV0wN3zSBg6xc3uGbh+BUA1pf
3tC0qUDImVSy6hj2tABrtllPZIzlIUSewXT//rHZdpSMDghaajylU7LIuE553vit
gPUebCGZg8BN9lL26AeYUMus/adD2CE7E012T7FicXxOeK+ErE5+wjDRhgnW5Ln7
7yqUI+Ynbt95Pn93WeS/KII+Hm2X7/WWMDxyQ/5NmyWyl0vLrs4nnySoNr0NBzMI
xMZgrLGJzdMBbEm+YeaHnk7Y8vOHYssxsNjeojGIG/CGwR2U+XGv5unXNGRZE35I
zWadQ7Q3HMPAsy6NjUqMncNMMNS/oRHWc6cBkA4hliDaNd1plQLa2iDqUmVHWksO
s4PnXOxqOUcVmrQryqe+9ON40boqxi0Lcx2xlGFTYm6SJDqso5/+vHdcWALSeh6W
7b4LG3cpLzlv1l1V1fVoEiP84FJ2beC4C5nJG6/3aLfvmhuP9yNabgBouraTDgpB
p/SxMe8bvAeeEchOID06kgq6Be3nUWvRmIfTgoSWxZCBKSOD6C0xcu8IdVSU7mpB
6yz1F7d9PeKRlYzSdQLObdI6JtwletE78RJ6CssLXwPNQ1U48g3dIkzQfUb24WSo
2WQBJp8C4GYa3vnLJnVwVR3rAv5rVHQcmYtVCK0iJ+J4iJXFeoW2X9AJgM+Doohv
Dvzd7LJ/ijUc9qLK8jb9jemtbWbFkd6AG+p6D+TYFH8+HTIX7C3F02VlymxJJd0X
o4oFvOvTSu7wW3QBto/cbaM+2RgLmUM97cKpfBIqfneh4C9YkF6hg7w7g0bvcU7d
zyUfaNl/DPzzqTOGB9akfixXlvMPeRDh9CuITDYDnbhOV/7dPlKocMq8eYFzbxNB
iSsEs/LUk5/wLbZ0A1NltAXD2biNtBJJoFpewvtSxIroJ6b2reYcQjLNZ6hvgOhS
/nSDwD0ZA/ZN5plSdqsqX47brHT7db+bA5eRExC7CKd8/LXoxr8JAIyIe6XfC4Gp
XnMaopx1aXCxcu4el6PK6IP4fNcGTijGgZSlE8kDL2S1FxzWs5yY9L+iwv1x2A+G
/J9i/0zhs8WoYBcRofuhyu88EKdWnTnfFHat4lqPHXpVY5nPvS6xQ6XHJUE/6fEQ
F6HSxT4gDeQ7sawbLdCV4GEPz9joO6XZCFrwGttd673cWX8gsOP2W9wPC3U524D5
LFfUEy3eOtJQ78xw+UflUVteh8w+3RE/NW1pFKCDEIfHkd7Rp55WTcA5v5AfXeSv
pHbUt3gwdwto2mXueiHyo1/okbcu/OFEKoXuIp560VDd4f/+uUMPj/zTBkYOa6x+
2+Y5mGBgkJB3VCJNdu977FE8zBi3Tgd0T1/6aYGG+U8f69Xn0EakhcsPXgBekiiu
kfEjbIOEDYs9H5OIzsHT70laIAAOQMeiajMxf9GhcVvY791cOn3nQ9bIZhrZtmF6
/Z3a7vFdgK0LHQTpI/kNClRUPiJk0Am6vGw5b6PYXaewHYfrLfyeoUuLOAMkMoqJ
GFYx3q++Vq+dUxFwNeTG7cFaqWKbmDQ6nLB1dST5UI6+H9Jipd1/oo848bBN3rxI
nzFV/pUpBX6sJ8W5sAjwX4hTeAPLWNjmn8xD5KTj7lFVTZo4UUDg8OHGux2wlG+H
MaCzpgs1oWEMgMXA5QTh2apeMGq6wpspxU5WoSLaRvHEsVB8qQuCrF/QD3GYz5iJ
Gr+AIFhQ1IY4TNbs1NBf0lsKK2nyhiPeNQolZ31J2gMA1MvEMSUQMzNDu/j3qcPr
hnROLEey3zUpB4yBVl/e4d8H/XMVjBtJkIG8csaZav1N74FMM7UXlTFT9fuoatGu
QS8T7eb2B53xuXJuG45goFlh0wB1ZgJfxr7k9W4d5xW3RxH/7SIRMjRmnNiXpYAg
6r3vD4RQX3TTQFtqtTX99Tkfsy1V4EQtktV3f9EqmEx1abxzMMCW+38I6VYM/UKc
TludQ1UYC7b+VQgOJ4q6rm2u0nBYXA9cEFBBdkETk7FNON/Vq3g4eNEIe36PRJUD
Filp668cFSqFq15EZyRZWH48lk6SCJz+mbS9DxsSYwnB0raizenU4QoEp7DQx2CO
r5/4/70IDz6UCPcvcmCA0KRJ2Y5qK/Dt9D+vD4H+5PqtsNT1vmfJQ7bFrUzBKTcU
3i2PbKM0swyhOaoGYQJ8gUlJDJePtA5R4XRNagA2wUhLoED9qX4IIB+oTP7b5HJ/
buX0I+sZUYmVr3ZH+wI6QRFvW1ZjksXbZud/yL8qgeyYYnxz9nVfgE+/59xU0EUU
nAUu65XWRQZbBqfyhaf2yXJ5kv0nfmdrlAKOVWNQLvOzP6Ti5ae9LvQ2f9qcB/cN
OmluZv4jhcGrVJxu4PzWKSBvrEaesa9hSjXJktQ9RKzMFMYrKfcNJRFKflETNlLi
8xYQPHP9WCJrfjxNEp5K95ns8b2Qm09tHFPVMhBpyXpx1qzidzKe2IcL+quqfbPl
MEAp7LySk3f7vIDWr37+bduO1hqCQRCIqXMlsVRAZIy5mi4jF9qr1z/Jdd2BMuf2
1Qtj8UceyGDdxslt3e71GhRX95r5N7w7/x1HJgnl+DQQcSQL+d0JQXjq7aKFqoU1
Wr8Xq9TIEy3+loLDNyHPU9JMNK1W+cgU0bh8KHMU3zax01OpGnhvlzAAhfXE3iw+
j/J1hJNxLNXK1R7T/6pc8iet0ZomoWnQdgzg0KeBeMi5VTVcunSCNrZhSUnXf8eY
YU1WKFJFpPWYNsJHdTT7ta365uJVBcSJOTcrK0LXbfbm9vj5IwDQdL/D/Vyk2gcv
zMnxUqQ1ldG5x3FDDNw5eUTWI9N58OVskqbvrvyZopjl0OjeueebU30QIjuWFoKS
K7jSGMEKuWxpAAncqTPz2XC9DbPiFqGTOuldPoB3pT1AjtpeKtDG2cbB0zi1ieWy
dshw+1+XM/nXYOerUF/9gSmEj/sM7Bbw+HmtSCsuZnYW+H7dfpJKro36fp5UHtp5
+ezk4DPE5kDNwxnmQnUP1l6crMKjr193kZKZ9IA3NBxR/QyaZ15IAs6fPWo69QKe
7PB4f1uzzuT5T56s4Yqh5R7mLJHGawnFSLSSoSqePbTnch8GSfs/sTZ+kDoQf8xA
BcOPTNAqylRZIIm6Ez1ANLMN5G+Yls0uHFHXzJKB6m8P6ONO7dLPJ0+YEPaMUFat
FhdJwLw6XtZD7GbFxAZ4I4UmlfUoQjiqfvVCT1dDZsJ8W94t4ran+RO47sfnCxf2
/z0c3HcABtUCt3r+jIE9l20xJOohNQ+AbLVi1zmkSPFCg9CwZt1ua5dCkQ9jMkSC
uB+M5SqMIa/eg8jAhNFUMW4gzghZpNy9w6lIpzJOUqFRtZ0Se/mXn6TpXJjMGzqD
H9tCag29UTcnSCYMv77zNwpC5laDB1/j9V5bjTQPESJeZgrUs5kdNXi9EOz/7Ujb
WDD7F6Zy7zU30BBsi9VmzzMftRiW/R/ZRxyQUv0gk/ZYzLgZZw7YlkVdQYd0xNWj
/zEwA5LfCvF8Um2xMoiSlsZenXP6JZQSfK/ldKjzQJ5paZnFAzBKkduQHs6o5BKB
OPU4hY5w6xDpMvzGNzmb8RyxTdls0d8gczyrNiwYufOe5zOoPn0oQ4Fv+a19ORvP
056yMQdMWbiQfBPsvE4gvh0ThVbO6EJBeiBoN9inJ0G5GcJHvjEjHLnJ2k5k98EN
YyEgmP0CdHSS6B9ohg2mPkbJ6TzGwpY3gRLezwWPhzp2S2S5CmhXWD5kTzBAy5+0
OOMOoTA0l86UnxAcCvFFd7yQLHKCFgsPmFHd562t+GSgDwFLpvB8B/efAZtja2t6
r9+vk5sd4x+ZR3uUZgXpHVEqbEu6lUmsTfVH6Td8/tUmtpBqcOrys02qcynge/AD
cOkLB2FtH5wPQ+rJhj+K6wvnf8qx6Pl1/Nn9/dIHjyaDhksXChEqfbwRe36PLUCZ
2WbttgtkuaRoo1I7RnEwN+ZrN5WsFKeRUn/x861FnPMLT84dzKtxqoRQb/u3nnZi
PYFaj6T1lWPRBDTiO3yb6CGUxTCxuHbpGNSBe8RM+OSrdQjAQYjrNRMyXxJDaavv
Q+3ugr0YgACidp6et7C3CC/08ldyOVrB7tmi/iI+muJa3HySbqtQs3nNzrWHrIMN
55N46pcjLzjCdd0NzYDdOc3+Qrrx34WMLHHNmh0cabeRsZn5aYRuukzCnznWuBZo
sUYp7dJmcJ9irTuMBhmf2mAOTxHi6L/hDnqc8D7Qqi5ydNUQxABD5nWAZlrbVz+i
Uv3e/INR6c0yAX+WQv5CseJZDTeIJ2OcQNiC2xa8h7RyC3X0QxrkggcF8zHEuMgZ
21XXD1WLAQ3xx2XKi9/REAFCdIdFMO38H61/zzCdps1dTSb/KkvdA77KS3CA+Rl/
osKq123UEqFZ1j5bSKUpIUve4MHl1rzWAfzyTh1tfwfPQorL+quBNcTRRbT5snjE
cDzS4isxHNXg0kavnHM+wDhgmYvf321xYjToH0z8A0lVrCmBPhiAgZwgn92kkX29
Uly0XiY+BiIeAxrULiYrAk9HEPR+H6QZy8M3uN0yJcJ+r0VRC/OkrV7AbIgiuwHo
wllU7V9kLhhWd2h+JlzPAClqTAUJYBlzLT1Kg5W7eC0HxLpocpAcT7bheLonCzwR
r/0hOeUVR0iJz0gF//YJ0nDjS2NlQf2r24Fzp2s7+kdNqk2yM60hz2++IN8fJkV2
97EF7O49WrZ8G7rGe7FyZsmS/GrUDXtJe8QT9WFX2YnNoyiFgc+17haRMYFutnU1
DO5PbHU+bUr90tqm5ogonMVqQ6l7NiXSIzOevNrQ7ywkdpNLjd4o2cZJ3smzEYsw
Kbvc8ZOyWxjRxDv5IWdqqFBFowmplH1ZsHXXFEI8VKe8LfiFY8NMcyWE2DQ5kE6e
YZeLdxv6dudeQJwQdXJKE99cqHahmbRvZyjpetruqOVzQoD7ZAu/D9vbGIJZJdFx
VdzlNdIv64E1qoyYRb24iEwAFdNEMb3Fg0mj4l4Es6HUDr5h2bTkhtjZl6r+GmIR
Lak+O9AuPECT7LguAkRhjEYbZT2kCvcfvKJyX/4NdTjzOJyMrlQX0uAU7Tq9Im7L
ipac1jgLoK0fkYZxrv8EKHlfCeFivjEvyrjBJtPihMlb5D3td8krIla9DUeZ6wLU
jXjEvQEk2YKO6r3lv/BUCKE7qYLNecDwc/nXWVhfUoHrVU5yFjiemwOckVvoLYgv
9OW8BjrW3GEKReIKCi2XBJzqnHoAlP2bgFhhCPYKM87XulGhTe5kfz1eASXLHfMd
ehdeU/5gFsUqG198V8o1scCvP8B6YUIe3q4jQed5UOQ/xiFdQk3DIolTLMs0cWTC
jq6jn2LffLkj/NE8M3WY6L4HJ649SBk4r+VrhwRccQby2uYOn/BCiPArki3nOJT6
LXWvWPXoi0gtoENcsqfT9dnwLW0vQhxg4LZX7rBbaPoEuwBaLGN8O4TrzHQgWGEB
AylTUnhlIzhTPQ8kCR5SkaTOLtweyVJsjRfL0YxPh0rAW49dwVb+ijPpfoAX2uLI
1GgJwJLj0sFU9nyaR1yBnL24jUlnSi9/vZNapD2D/QOFN4emWYTu11zZkwvjg4Gq
OArioIuDCGJQKnAkctlWftdoeP6ok9LZYgt2J0Gi4vKJzj2EFycj7ZHmzPynY5wZ
Sa0UTVRE7suqyKlMoiWz6HHLqwL7GjYopsqihL5qZ1ZMGhELADER8YtntVEHhUwt
UJlKRXKyH3r5dPGVyMybKn0a95OEs8y4FmTlJ5Nv+75xVPjs66LLSiteDJXzeV+k
ethZKR+w/Zx8nyBj2d4JII6G5xSv8V8LxRaWWsT+NbZCsrSrz/b3fy63xYvK0HHy
KQqF3awgVjE7d02l4m6lf6sA1l4HH7K7Gw53QtNbHaNrmWMbz9C2yo7mQAiNDCTo
Zm48iEjyc8esb7AFZ/ImryKJBma30iKr8YdcYTIIl4Bap682QCjccUYrtDIA9leh
e8Pp/4061jm42sDUPKTM8gy5c+EJbwHP9btl3U1PtS4UhQNkBgiRkD4kk/FrfO5+
6N0oEncIU9Rfny2xqsPEOA8Y7jfhrW0W9w2s/XG6ttAtMGHGVfr/LZwdJNZEhHeP
jq/j7o/tcQEIbedTh/ddUl/TtfYrpiIZqlFiEcXv4p2rJtp5FBUTojTTbGmB9rwr
eiL00luxla2AfTNjc+0wL/9aLOrXChHnYZTdEqgry2K8AZt2SbCqzG8ChTs/hT9J
wZXrWk9wup9cWNM1msNFTOO7W8Lvn/xXE58VnJotvsMo5Sla9KOjUcGGV6Qf5KuB
uyDp8vZp0ki5d5SaKnYxu8XGuzHqIjG6yflMwYZSFSfRCMu1Em1AtCPNSXqm/KqU
6E8rtNiASm+6qPLXbtT0yvoIC822f8UrLv9qYaA3bKSZ4b+ZFSVg+q4PCUL7hNYz
5lzquxZjgBVW7w/1HB7dBq4E4buKv+43c/BhBI0nRMdjylm9Vom3SqyxIlSMpGj4
wmeDTnSOoH30T1nut4l+mOoZdCr6HnSvjKEt142gfMvY4TuFk63UHS5BHWyvERTB
mCFlMnQnhw6SgjaIPJ+BIdX1MlXD0k9YJiM5IAbLyvknhTGbloss2+qqTd8k6X3t
4hPxhZhV1lLg78t3zvg0qiJvGywaZjv8rtX9U+kWA7hXUFNasnGlw0AEL0hYApL6
5E8fkb3pT88RQidnOumyk4V5bCzajMzq4HnzSE7mz8A7Zy4dnn2IaqM+OZqGuskr
kO2mgYGkDmtc0Bptz3kDbSwRHNc7FmE56bvxDCbFfwPhGTcaUTXS0fPxqM1kL0/z
liitRZvvi8mhuAiKntgfuh0io/vDWqxe/vARAFwwq/2vwe3MIou2YZcLX7xBqlcD
YEVtYwJjBp7pN+O0Eoe4LvM2of5+/l0IyAoMXC6twESJBhcHXZhh6zvheWQE85Q8
UVzy3WuGYcp75rw+sGaqfxQMx+veMj9r4/tjXUNbJK2v7KVAmx5dCV6sNmpaTHVg
IIR//3vgOwkLSbiQCpumIjCxFAFM/9K9FbThPr96gsIQsGtL0qip44Jb5Vw5UE/l
vdY+ROCj3Jhkld/SoPsDzJD7jQ4+kNUcEU9sK/sxCRDalX37zHMk8qkNxcydT0pZ
I/8CBcLjMJJuQ8fJ6ek5ysTN58++AHBMahbiRfsroqyZ019Yp0gMgjVxnQwV975E
jb+Bqa3kr7Y+M6kAhK3+OLMmVygMHx3ojd2EzK+ZeRuD9qusFuqc1pPTtUiV/Rko
FQrFyhwZKM5P+FbKEoOb4fRooQ4A7ve5DuvWsPbT2OUfLeg92B+evFuH5Uj/0Ftw
OXxcTLs98Htb/pz514nKX1GJ0ydgHt0b/mfQ4ni2DdYvYUfsoGQE5RXAiiKUMlOM
JPGD5Xch3D2zbVALveIYEdvLOC0vumYS6R/IKG5sHlFtY4VDBbNKoAg5Ji/WbYek
KHgfgnKkrzKj2cI9d0QtpW6K3EXxXsyDgXUgpRyupZ0bB4ioH6Es1YldmVBB+SrU
3kqHWKXEcwYHFQj1RW5wL6fpd9bEELH/DKMy6pZRcN8xKZVmXA6Ck4jqcj+1qISI
vsELr1D8YF9l23wYlTXe4tAIUiMJJZh/opOx9laBqmL81lDOpxpZrDCRfnMSF2MP
y/Ki79H3SmwCgC/JbMJ0Ne+ZhXYcYf1ivRhE9f2z62P7oB+SyoRlZQapJucf15il
Hlk/w/bZkbrzwarXwnotIWy/4kMsHO7OPe3UtqKmxXffWFemUUMncUuApqEYQjnv
I5/9zdVCsEmoscjrGZ2hmL1ZBaULmHLGmW1OgPPhzBbOskA1D/lWUwIyokpVt3sT
utyJUBUzkkNG7YEBb36VVbkYni2046nnKdsxVrlMXEnaUt8yYqtaELBNrVv/mdp1
M/8wiwurEQeehocpOOKriX8paFIuBoA9shS8rAZuirld0N+Du5h117VgHyaPVOV9
EFW06KgaHCqQBt4jNuwSraBilTUnHqA1kVWw9zJCJO40vdanrgeYaLLb0HsqcWrp
5KgwIyT7GfQXYPYrn6ZMhhKDPKfW4UDXK3BpxbEFtEO5mKHL+TRGWNGsclrdA3Gf
lEGGMcJ1IxM+cTyeJeySXbQ3S9p3YbYUTJdxyF8egnjppYSI1kXl4QiiLrILdQSJ
aITew5fn5i2LkEkqWwX77cl5UfLdBP42Cl2mJgcxqEki/hjJK2JRkBP2gniHFUqc
VoonvZIgIKKfb085Tv9nQJgc9j4tldyFZwphMRwHYH7O9PP2er+r2xjGm2Xo6Uiz
LlAyBQzzZHjxJTwLhpV8oLPFiwsg50Yj5K6kOtVpSh4+Du9T7nxhotb7cbuDEv6/
ai7vUmTJ8aud0NDE2/amGUPpkmvTbJEDnaWxAyJlTcVnHenC6KJNYQRX0y+BvqsK
dH0E9PQCLUdHhExflpsh+PVcTIO4BsXEqE5yJ1/fXCVYxj7tsd1NH2FVMc0OUyfu
6OHu04nUeCpErsXXoMEI/ilT6vKjk7NOYIyOS/pIksXiHJX7zn95aiFkS/D33r+r
BVYqsK5TOKCd4EPGbqcuiz/dmlROSqvcBViKFAONx/m4BPi3l9HRaW9bZIINIui4
jhGHgOi/PxD8Whdn/1P14bB3C/fT5jXm5zfdY6JqFcNoXNMF/KzHWAfDPLF+OHuV
0ca9r8hkCjFJLha4SaaMWWQQ5fHUwyyNR61D7qTRV0h6pQBep6Hldp393H2s3Owi
16ygb/MU1WwlUV9M+XBEsxJXcstrEHK2gyib2BCStMOj2sU96DKUC0/WuOXC4hBr
XDRoRRa/HxSDrPjzaKjAh7Tb46AnY5xQcM7UnVn14J23aGUoEd7tTj+Wd8mq2Uxe
WtA1nNZlxHubw9AjCPYhutJMC16q57nkRaylath4htwXqPyTZl1QYVnd6vkE/0JR
oTkDJia77i9dGBxUqmESA41/OEi+Xkn9zpr6/PisUThDOoOu5nzZBRn05ezfr0pN
7Dwy2hh6fC7cKcMMW/BDuEsgVCNve7RzLVdKyAwiIbG9ngtvzKJzn6mMJlGVoJyD
+lLZ4zRizkMhBcafdvOPcDX1cz4XAzh7OQc3oJc1lI1magMuKmHfEBLcv4BLQwuO
qA9nNUhw7roUOpbj7wRVq9S8Ggd6Wqp4yk+/c5JF+hfFNNY2TxNcKuC5OSExB8lF
am2hVfyNor+84DfBRzoKT+RODs+TP53GnLX+IyBKdz2lmocaO1vRueqmvfLyvVrZ
hkIsI4zUAy02uDHisf9QbmwU2+6iLTkqFoN09uL0/qBXcMWhMsn/xvNkzVWJnHTT
ewxRPeI1qvvfS3ex2Vjq71899GFI2dENULm8tDwToiElYSlyPNdETUzkLxK7Qa8o
s4ROq5zfRrV0IYjutyXxR9zWzxNve/gnjHeL06UzIpmtoFovvCvuUlAL8KYNKGoU
cFXaDMVFmZqn+hvozxLDJ1GaMxjjtcxHlZddqfDnh7ozTpPNt3DfGrsKqt62xt3L
gd4XJt1yb/lr5AGBZ1ytBSUuLnyAwDrWzUW5MXKXoaQpF4JJbhwC+7N+r6zWmRaM
ggv2L1V3SMaJaL31Ra6EZOhJHcKt8gHnSWtPWfcSdaZVMspBkWBbBV04alcKQTCd
XshWFQr9SVr13pMdyIJJHZ4p2jcvTcZxBbWGCpOFnPwfW0ccIGEOpzO4BUMCnAjQ
2GtM28l2aC01ZnwQqrvqdx5U92tjiijg6oKubykF7ngSzfkkXOw+xyZ6+3jn/DJ0
+53Vm+cfQEATR4BUXn60LVighyJC+7zfWiOU6YpsVEzRFHVlRPIylB5W2w0n43GO
GqvSpcR9q+cXigFVJqsQFuZ/KcOcRfegXi7GlHWB9FPWtB+xU2ipxp+CV6MPgrsP
sr2C22tGM8mg5FKA7vcAOktf6kfmRza4c11UYlWom2QkzKwSVbdO58MVAijyrqdN
SoAG1kQ1tRWxeR2zUy57hRGw60xbsC9ZpeScMr32qD6JM/9qjFmbmgjuBwpZkdRm
LvrWfTIAPB013fywMc8FfGxbvUB/ePYMx2RHW5PhfbeJgLvB1ZcMim019vt7flNA
nKs6a+Ilcj5JL4ayWk34ghCt1YZpGd0O/rnW9LzmZBlNrAh4YcQ1yy/wvBUvkJy0
zie2gS8x1oKHKvFTCzv570xpAmst3hO4Ed0MPA/UuOjbeAh/lJS0CJ8QFTGHUKlO
IP7OBfAHPYWqymFYnPGD6Rl3h6wShDt4KSWAFjeKNFqMK4jjKQVnUyP3SZoEPkNt
/YW+A3V3oNg/lshb8tfkv9wgFJw4RXVBhzjinpXcXu+AF5lVvJ2uMps4zfzxVQuE
MLUmR14F5Wawg/Fl7IeMoeT+jXWQ46tuP5S0BiqFJA7smV1IT8jgRlwVnVONvah8
D1SCMthqTSips+lDPXE/218BnCzAzqtKgN/p6MZOPFBw+Nk7bluRVE4lY4YjSN2p
DAstMyE97kQcI1w4++LfR8eqJuqKCw/Z2rt5FuKUiKRXpUPUA9wiNcQHcnnp2dRT
DbMoKzLbCGshv3xWpoTC8OncrVO59/6/T3+fueGc9gWqwDrsnfDv4Ehq2NVJ642i
Eoh8ml38ZwByU85Dagu0Qf1CVH3qeQ+LDq62gwEGF4rpu+KYH6bOyuxkHFu7R/Gg
si/cptzGEUvD4PeE6kisZCNbi2XhLIPG2v393Z56zABhuOQq78ABAZS0JhkoKpDs
Bv15og2zN6XgXxYFIclIw1o/9zvre/kIdkhxwUeOV+eefK48RdlbR9Mq50VCvuWA
6QpVmadPPfi9gxEb1RwRvJ+XcBvom47wD/cuQpCS2baeW+TrRIme05oCK9wz13K3
htqRAfvIIvwjkyoM7Cudvn4cYopVWaztibPQA3eQGoymhZxj1DvZUvrF2DI0ajyx
Vll+OQEjDZ5XVhQnUpymqdsmcM0/McH6RJTy7F5sm5h4hXpQhj8cZgfhvbI309yn
6trF/EeZlFVWkS8JCwRRIE4SCMCfH9uLTBMNknt0NjiHXXcd5L8Bo9HvEU3ZvMFU
MVVH7mMZKuEtaiIdoD80/xt948UHPtHprYxmtMFVjwJWs3//ky95GmwA8nyDzoV6
Rxj4bAM6MNyUOzR1HaYIYVzfQBmBf3qgDJMPeNpEqA2884qOWTao8pFoDU/uO9sr
xG64anKCW9baLOHQY5oZpZDMluNz8JbBExdoLvyq5sqMlC9/boFgAQH++qngVnWS
RGDh3trpwbuLPvitcOSzc+VN9Aaa2JDVCQ1lyqgCzerrOxNdX5iQSavygPm9cpHZ
6ItvpkCa8qtyf6XKw4Nh+ZCMTyvRNLAtfcxv/1Npjfo9NuLnoCx+qbNuQJlmWIqG
CDHycNT6QagzryyzJZ9Ews6wUY9wsgNbPx5wAleh/OJwlXKHvxaniII4e9jbsorj
TfKLeFH0W3I20GmUugiVgQ0A2XIsLndZPbC58oDQUJAU6cjCKw9O0TrEmAwMa1Ek
tFn4Tn44hzE+AHPHuzvJR+RFevYXreF+gEnK/Q6XFh7VfTIHhVUrjs3kRv6yRNrE
Qfp6gEtaaFd7MIjcyt8t5/8mq3nT8+vHUx8V9zpElj2iuLa7kXuN4APqxYxnkIRN
nw+ZE7/gL6jou/Gq/Fcliz7Oy95UnNlVuFBpuMGxWxu5bQe+XDzq4Swpu+Cepvbx
Ec/S+ZMZbsrp87CDAoQuDOTJZc1mxgcRZ8HXDR5+eYPxvhHEQls+kHvzEyGD7h1o
cbRBApM4Xjbm6NspmaIegFtvETYzxdxTCc8tcxyyMTaKec0wjEKLJlyVnhWU0Jax
3zFXuEHyzQnSczpep3zS6cbyqtQyROJsWmU90jyhWzXwHlrG6Iycuxh5fFjhuevb
SlgU8OL6RsyKicOum4Glk73gZptY7MbthZAIX22Fc2Q2qnGiUm/UbY6ru0DfBWdC
+Wv2/ce8QAIRYDW4USw7yuzC/B880PbQzO/dhkutkiRwev/FUf3doyQP7drSRVp7
flT9Nl0DXe5fMSIa/7Tj9L0OeuON3Twlcv11bp4mQI7hwk8WSNVCA0+iGEMeMhEd
/S5ic3ak9mJuzLfEAEHC3r7oRQTUSqxtutG3BhLdoOXmIH+n7ZaEQIZnUz2yxRp2
/D74isCcS6KIwoOSStkXnqpDgEO/6v/tIPwAhM45ujZj+IimHLUTG9InNxLHb2E5
F0Myt5Town9yKAg7/ik3Dv7EUGkgsWawNLNHQiBl1YcBqAWRi9PnMe9kTm9vAv+S
/3KrlaVWgDXixilUL5CJfox0G3MAenqMc1qr3zFgWjXY++uYHhi+BdZ+lBQadNYb
nAAnWCuTxpGb5lMrvfc0dcRKsa+Cb33J+IW4fldUqGQgbgUN9MVV4PyN2S+j4t2M
qkQNowxwFdpU0SexrAOFNcpgQt/We+E95QRdgoCFkUwN4uv3yPK3XfN0udKjIGUW
hf3cCrvY9H5yQH3lH+Zjer8KNne/hKmjX6BrT126ItHzRsBQ69lUuV3kmQlbSwnx
dzt+XVQvjQr9fKfaH96xEU/vrvhL8Ukk1iCZtA43gaX1iHVKRnoIMwp25DCqQ4Un
7rOpOeB++n+iUhFELsADb4tuEQU4ckr1M7dLdUJJw4k0t0r6K6RejDbeq8y/FfyH
FiCuAjakQ6gSGliSwtleDuhxc/z3ui5RBxeTgsdpK8Qs9PbZPVQ5w+XYUhK3g7OT
NTpYIW/GGCi70Xqwco9gsx4NXVs0eIsbkkVMR/3Mqem/0LPtWK0rQMriA/1w3jbj
ts/Si2muo8lCVcw88ciLXzUYZglwcBL5yBZXf+xdRVGsPKmPrCCrTkPAm60cp0im
FVILns2m0QSwufJK1kwTthQlRmFHFLk6Vnu13yUkbDyWM9UI85yDy8el8wNPPA6i
iq57T0KsC+739dqVfE4ly++p+FRoyNlmX/z8P2bs142sOCVZqdv3pwW2qEqd5xk2
0PzJ3ucK3zwT1XQFVVGuGlOPRCCnxZyoNRZyALpgDd3tQcgi/9X1mHlZ+kFHuqFJ
ybi9oQ6Ij76qks7EuCxDxGRyeJW+n7mK3LxIuqoBXxzExorYrX1uvosnnYwlo0QW
Npw+1U3BbN8CsTvm4Um0efK+1IMrL8wlCXw906BJIfmNykS4mvqmTPMWO2s1C3NI
elWHcIe8AVBCi36YWI8W16iOvrn6mPWqX40MVwcaU/7TDghtswWQliKJQMSdbCZQ
M7FrqkiSKJ5D9wkrCBSSF2k5NIQdYsbcP6rD6BHQwOOFfvMFyZOmOAsnErMPtq4N
VHO2a5+YAZChnvEZ1jUncgDy79wGY09EquuTa5+poPeDi6cSsrv5jCnUwasq9Ohh
mPLFfFGsRj68Dx1raDvhK7mKHC2+PhjposfG4AutykwRYwZ/jOe8T7Wc5H1FsPQu
FFZ8fMZLs/pV8ik1GmeEllAF/O4c6DlwuQOzxEB+Cl2WMue2hQ6mbTv8Sfk00cZv
mcaAuf3fobiXOR1tZyd390DKnjYgefIXo/xwWgO8HoAeLRwg/lq2xKWFIyTJPeXC
mzxOYLQ+z/8QzyByt+je4cLwgUXnobRSRn29KhkhFzgaCsmBICQ8+7rtjvuRdwPl
pTWDYD0fVyoG27svylniC1/rQURPCnbnPOXzHZ6Ns9g54xvTHiKjGzRZ5uU9Evz3
Vtb3Fmu4WHy6pF/qhMk5t9t+9AZzOS4BD2BQQd7/PhVm2Ep9rPT1EV2I5VJjTZ7j
OWvE/z1MUwO6FBntiBPuklIEJ4Sf6zSp5MdJhk8quuhJ0I8kQVL1aker34a9Ujmg
TfK87aVuFTxLs+zmEqlO4fF01vNYfNFwc3rut6XRqTtjwjPq9jugiwl/mGaP5jha
vSpdeMo7h4OE8y5KBJP4p5e2FkDYL/8UGDKloiD6oviuVgs2mAciwXYhftDFCf3s
xiWbPLw/asAJ9GUbCtPcrzNyUhesfQOCTkkv3zQoHh74a+Fp3K3t/pGIqgtgpzJo
aoB12zkkZRQcvhJ5kSwyt9B5TWgjxhOtWYizlJYpaLxW1qsCdK/5Hvp+VQtsIvZF
YfaLVHn+vK0SQftMclwx4sPpj7djxyONdAU+S38rjQkhnPlc520I42fohc1ekmwl
SJKKmQ9okZavmjBIo3ls9I9Ih4gT9dlZ+hjc95RbwU50z1OJ+hRrtNPRZt4mmjlB
3VGk4aF+LvK6blN6HB+mH4w552jeuPWCUoJVVqea8V2gv6GSMznRMUFX/Rn6RONf
OdX3yi6mwnR+bqv7y2KCCpcFS/OuvMhZKMnRl4ivcP5jrogh9AwJBVsfz+2LQ3rG
0CMTfFKY4dVjJ2vkXNtasjm9NTttK73jX57HoYU1ItNa5HnXWOSR0t9+2TgxrF/g
y3LB3fRTfLnO3pfsezlV94s6nwAEB0pVnuX76OVM6+YLMyahBeTJkbKVDY1+CIgs
YHcPj+Rc3Yub1BJYFuDwKLWhGC5/R58GCP3s89LNC9bbaf9nESBaZtj/mEClz4OY
tqh6LDPOY2rD1bzTozstfVh8h+1x6shlU2yE3BPjD6GeMX13N0gB84sAimE85gS+
zLKM3zA7BhIn+jtesfVQ9C/KVoEoKO5idP/Xz2hS5eCqpnga20QZnTbia2sXoNQw
ePjvjZIcFLyO7B/v0J66PQSKc8VDC2DQw4pcfV5OIvn6YU4I7M2mjVN+ajoUe/Ct
QV/ax9Q4VGkJzt1pBNrPllKt6qh2ugsmuUFBlkU67jbA3nenb0TQTYhSXykGRVBD
XvSa1MrsE81HzzpjzQKJsoAmgTU0e3SL5YD0Ok5zTdbLczKgetEIDtcW5JxUrG7x
fK5ZaSCGk6hNFvMOfBQUAuTRs6op5whXRa01I1egx114MUHp6Eg5q1l1bJNFkGUU
PT0lscSFC36j3tnCXfh+KrUK9ti4oqvji4TaMMjSCXnoUJHJzQe3XuVYUPTRx3rH
Aq68Zrxf3373/lXsm5Cmw1gwi65EGvwPqlF0avbmPqW6Jt6fOtSZhaQcwCpBr4zq
+z+/BF2zLlPG4BpkRfo8XQeQNSEPOLDt5Ac6JTBh5rt1WoMfo+kLvHQC9crNM7Iy
jTDXVdg73NFEFS7E1gJqjeFOmO6tD/EXwKh/uDjPEhZgpDvQQEuMpaCdnHipNJOf
pI8XbwvqJ8gkQPLao2ll6KCfyA6h4V7d3X8xNsnHhpvx+WuSl9e0nJiHGMZNIIKR
rrBAPnc65S9zEpuT2CkJ8r/YE/af31rBSsSWDDPeMrxmegMoxn8oLWhLbpukq9ZR
DtDDn26wDR5eiTcPWBt4iQsxqRMlovRHVbbtDttZSydLKT6uf9ccxPz4BeNnZF1B
TNQNjVpaHiUBh7VPDuwTkIv3xb8EzU8CnYXYgPBFGzuIZJwpx5YBKzFIWyXak6Y3
NUom26B/maOGO2azQFw2MyfA54pC3VPV1S0Yah3LGxQT7q5OX71fcUXIXVkVsCBy
9AJnYKz4zTqwyRiEKgNKwc/nEd07yeKvrrM8ojeSeHlcelmXdWMTdqgTlTibiQx6
c87F6yEnMcqNRaUQj46nD1DmWqTb5yguXK1dBGmi396qhCitl5UVr7k19g11L97Y
2AOzzXfEHvE88UKgLdjuncJ6kpPCkitIn7fcfN1TE9NsxMLiBOj1VCRy2y3BoOHj
F+4DjAoL7Sq4cIaM/iJUmAZMFxfJBlbfqoCyU1pZ/xF+XWtIvbYCuZUTFe6APpmp
O7qcqqOUCMejRZboQDx2OhV4TlpzWGFQeHUF5OjiYg836Mjn6si0zoZFy95pA/Vb
DcM+p8T3LuYmM2mkEi3yuImgWjgaepEKC762GzPeSKp+nsLaMNtWD4umTIK+Tiyv
/yI8KnZc6ok/0DYz/1BcoXKLBav8lv4aGXf4taTNuT6JbEMvy107vTEwByXGbmVs
MYfHA5uUa+PXkdqzUXpHnZE8ornIr47uRfki0xAOYMek9b3cO9XyHi7s9dAbWdho
2aP1XlO52Ga3X+/CLVx4l0MFmSyXrSKWuiqXbxxTlB3vN2mWeMilljWJm3kVrYoc
PSFAe1TukU+qZEU4bE7IORNYkLDR2+oiRW7NxAyngHZGEFM3GDu+iAPtxRStTNR/
fqYtdASdXWZK2KxZngBLWmFGMC07uQeUZikEmU+oQbxdbnEsPxoyvSNf5idANNni
fhrbkakRxaJpIppH4oIza/SWgFazr2OiFPYjjotA7IQypt1mpberqq5uRm9YQNGN
0SdfAFdQf8daL+bcXaZVbNugH+TlI2EOaPVM0TAenMU80egzK3F2LFozZspfLmwl
9zVNxff7LN25GYiX6fUC173rSgFvCXwijWCuoQurwf0WchSOrVskFbLJ1hvUHjiQ
N1bemOvarWQxvXp3nbq13sLDm7/QfjM8HbpCST/i80RNflVkSaVEO1SOsskjebVr
wBdEL9oxJ829J+tuvgSq/mCYNu83h+QbFM19NDgPlZar6wyHBJF50xqQ7puArJ24
ZJXabpvzEzNUxOlb0cqNpk8zPy1IYfGfaO2w4ElMBBUFn9psTXfKPujauJCO6fbM
9MKmOB4O1QNz9gNFB3mLt/uL8QYgYg3wQeJEUnzehNPCMZ0+FjPclkGzPwX4g95U
907jSC9nHiKyXAxYT1F0V0pDnjfYNai0jNlzlCPZTIPVrnEYXzGpoyb2cgxv/JmP
edLqzRo4PTBshdHIgf8bP5dryWNQQvW4msjjzOGUCAVyuPkUvDubXiSeJtLZhyek
yNS0y4MeAnrwDQmeOaaLlYYzX2Kf2hmZ8rLZivAJa4/IZNcfZRlM/bsrPv7b8TFh
r8rOJaA7pAzrJGPUfDrgM1hCwW1haPwiQNbLeShcvh7yGFmYT5JOl0drdmuDKRw6
fZZ8kYf4XuBD6ST4n/iYXTq0PBpqxBKCJWqIBiOiebPXWHh88soItCTNSCaJTM58
Rup3Jb+BBMQDABieZUFgfluVmWsDnjU5lCGCWr0UnaM0UarNlqOsEgU2M7ONMwNX
bvCA0tgW3jvZwa5AmOVQyXm+jeosMLxqaoQcxvhIdSmoQMYebDLNgAzs81qPXZoj
NwOs7bVIbTn6rL8V3FXVo0swGEqvbjlyY5dgx8UhwYDkEpnNrnNRsbIQIiiLD+Lr
/pz25duNwGx7jsoggsiI6VWfUjEiRkYraj5o0BSnPCKbguAreUeU5jScoqr6IXlE
feDDIn6JW4oUCHKMPnWka1DB5VaF0VEJaMFSjl9Va6ukLmufk+3/CI2b2yPr9mJT
Zex4JFjpOFWxZN3gBxdUrmT20zpjRWAtu+HBqyK9AMFprnwHdpM7oENGqaB8zeHg
qX2vueFYnyhkDbCSW3X2a/0fN2I0aGfrSPjO1OIqRuImIZfl/W5jvJ+pBqwdIrlM
kBP0DJAbsWEtyNAP/LSt623AV8lf1IDE+kEO1IcFB7P4/wNpW11t7TD2M/ooegxJ
aUQXYOtpouj6PxCtBuUWT/jqW++YFlHXkaKH4Rvb9BWDN8x/YJBg0CVOPhL+9wI8
9mNC7OsTqADhj9tRC0u7yTVVOsYLH7eGQ9WFMd0+eNsWQo9JwaxvqQwWxYmBsVGx
EvYO2YneUTnLgWKug4XPaGV8FGYeqONa22r76AKqONDdrHaNG48qa56C14wZyRCB
0d6UqUe1L9DkVDBmdFGH0WqXrcckN+DTz7/hYo5pa/w9gdBLiIewK2nW6JgF8JtO
N0MhpUch0SpJjEtiUBeLwGGk1OwcYKRuESCLC2AQRu3OLL5WL8H2Q8sB+pt5OvSl
UQ71eQ8XX7mccyYgCMAxCc6lnbLgWVjwAhsFuMUM5hZobQk9DD7YFZ4LiUr5p61c
blxxvCxENtLO0ICdpsCqDOYPdXWmJRQemLTcC6DicbcZtURPlum17w81YkZAxiWn
zWSVLrmM68jm8IUou1W4KTBRGuFklLLQNNdpIf4m/VSeI3PxFbJUCFxK+XG646ny
iVjgq0LRDTNgeaXK9/IOTBJ/GzBdO4ly87AnuRq/B/ycSIKLhDV4CNrCwru3KBTr
WnWd6wI/3mfAX5lnQvBREni6Ao0UjE3+T9ALwDLoiBLSMOEwyDQrktaCVJffewCv
r/BvVwYcz+C+MKsAvvgEK2WpwWU3mXA52s8qzzp6LEE7F58a2AK5Xnfu2l0o4ISJ
wHYI85BXdKEomWezuRXn6B6qU+7xnoge5mB/bDurfJHPp9VEG78xUfUAb6KlB3eG
sJWdZQHaTdFWAHRjMFJQmOSRf4cJyddyxFeKUPFUcF1Q0+qam8kBBnN8dtIHo+ov
a98eYqPCzqq2+0B+FaydX7isoI8OHlCYyj/zisKS6rxejnTOimclY7/su8EL+D6k
IdyRBmRqMUO74BWON0mj/ffFzur9MZMtj/cQNbQ3sylE6xubvSDRjBbQ98rAf8DM
4jMQzMPvA9Hgk9wWyVIuxWHOzw4gAoJ7L5tQt5OeQjJ6nrHcKpkUlTDxUob+FbTf
4/zx1EZoxVjMLFPGXRaMoXEnkqz2lgNZEX2UyXtD0wnxDapJma9QYS3bp5KWd3Dg
yKlv78HYvSW4QjVYtNhcttnHNMsRYgjyVnjFFVXFCpVtb+5kZXtUvaTUcWgkGW8q
a/ucfOVM5oLE44AxKR0HvxpsnLrDpEuFkEVbgDGV328O578iBU35gZEEGMZul696
rsC7bN2AZ44MmNWu9t7Ja3YbUp474p6flKWZrlai1ujrj3uwwHPo5uguizYLjM7t
TvaOqXzLAAi/mJKiC4gUPBFgimxdCbUQMDdsnhtnWDtW3+L+dAxw5NDamHFR2LvS
4otBTY2DL3Q9yuYofXGsaxDeTEl/yTu5+T8fw+Pkxjc6jhQ8vL/VUWC+99j7zegY
GFKTVu67qnYc0UpNmQVT2O5KFT00nZVWskuZag5Lfks4ut+OPBDyOOrg1nOAv1wH
9O6JvWi5dJahKj/nv/UlZrY4H2UXktCfWU2phoAWTWG3za5lo+k9LB2QeszzyhkA
V8YOxP5wubRQSZm3OurVYLb5DMlCf6DoP/VHJxAc92MrPFdW6FBlLyrsUZc4sDWe
VJO2mB62oUrZj+nr0s1vnXhqyc5qSbclRu3aDnUFwYf+Qn1oBe5wFsBsp1hl4Gar
NbS4v2L1wvewiRDBAQcwWUx2lvukOLcmcmgi4rPEf98xJyVByhCO4uHr6zs/ux4A
MQvxLNNExK8WSdnOn+mfjBkW9G5BninBbWPerznbN//k/R7t9u+FW8xhncJXCmKx
hMpiyNngA8os8lJpOktOblX3glok69zsB9mzs4rV01gPmmBZeAz9qrh8ap51Wv1C
zD9V1m+EqpNidW5Cz8E7niBp/V9hL/hy1BiBSUu5vhXoqMz7McJdmBA2LuxGLHm0
xw2/1d6y2JgBxAmRjnnEE4F2tBck2H7aOP6WuQ6IYR0vn9LwqUkZ9CWyTK+flX0G
7XLiDPJca6pWgvwg/kOAQFDo2ZqDrLWf/DP2W8p+hYUr3U+5mhtaDUYrhfbiUVki
5CiD1jTTGeBr+pRr0LN1XikHq9zSCCKJP58zKoeq7cwTSk9BVPgg9WNW95NAnFSC
AYrYimExSZMY2Ccr+WHFBjh6EfK37hR7Wgoi4FE9B0kA9Xitu4zKsyoXhzPt2kNE
0KBQgD2vHm650M3W7AKFc11+PdumLbJS0LqVyJn7xrWCIgDwqgLGGbBhMVxtbi3B
5yaWXFh0uBTDMbBUFgAvmzZH2PQLoTBagUqec05/sarZ4lD8sJnfgwKNhcPfbYUK
px/Fpkj/c/o7VuzD+OqDWPNbfyEusSWdXKIP7Rh4giBO7ARJJaDnhDDeEbApPEyy
OsweMWQwq1jIqBYyDRRtnaQfWZCNEVTdKBsMYNLh+mzZn0ypC1bJpm3ZAw+Up7QE
TQtc5Bw1Z1KGqNY0Zh8GVCdS2K2LvK7uKZc2KMGa9YpRr2zLJohikVt3xeAMp4Kw
C7Eqpu4nrJ4ueHpfGFAp/YcHQBNhabNHwGIEfS0AQ/XxY7mUVQMEgvxQWPd946FU
sAa0MM5ilqiOx5afxZQKu2YZ/wKH5Y+7HlYQcVZHV/DsQVcdqYUfjPF2q7f0z8Ck
Ocum5k8qRwsBhi/WzOMhcrlyWSR7DY+uzoiRLCgSXhIv+/MN3NTdHb0XhTfflI2I
SbTBxAdM863Barg/ij7ca6MPKB8kg72eLxEFgH0oMT2Zk5cBfAt9RzULmGU8AAW+
jj5URwrBTqVpNmbTEBja9q9TJTkOW+jD05KMbZ5WUzsIm53zZemcwiUOxu8A8lEa
nXl/mZYz4lycDli5RM/FFFJjxU2IX2SZ9sJeAAbcsi5SXjhrr+E+RTCDAD43sEmW
CDnnDslzv8FWawbPpP4Sp1LtS//EZisxB/7WOa3vuoxp81iVsdklBOg1Rwrme7wy
5A95g0pWDRUfSwGzHvkbOl3WdglJn5UWyTX/F+V4iOU3p4v0Nal3RfKm6jB6KAJd
oAKBH4MBDedyaQoXPEKask9wLzL3ni2bs7IgsSTT4QkA27w/1VvQVYsDfkvXGZmN
exZn5RWmw9eDS1HsvbNxivOG2CZ9EA9xmUQb8A+Jt1wVmysySG6abLwfnQS0EDBn
IF1NHYjt29RpTcoeq5Uz1x4Zs8DPBQa/+Gl2Vp+cI96xiNyultfx2x46r6jqTaTN
8vQdsSLnEeCvcnecgDSXTsEIRfgq0qp++Dgqkib+I6TcK3tJHGR5XzWzp5CuKRSZ
pCBW+tAldgvllNwe0l6zXUQtPO7UrKbUQKWCX+H2AtBkqfPzwiC4e7yEXmffnc5F
IgxgWrxKe2gEqvtUueeLmsk/paVMhkQyobITa9ymUPjE7otJk5jOQF1hfbsX+yxT
SSawW21lsEXgO3YvCud1yO0XNXxIWIEXxpUxzJs1Sj5jKFE2G5YS0t0PAhANjqIk
S44X+JyvRyOL8m5eCrXM7rB2FnEkiUPSdlpqPg+WE+WA3nxdSsvpTN1HTusaBSuM
XuOO0X9POQk7pTcg/ouV7G1SSmfibHohOTpXoYNAb8w9dtQxxBM1LB2NLvHR4DqR
cF5YekpAbJD7JNk/lTxSUK+0sePQPSLtBPU2IwMFHLU82ZGAV8XcIjirTEjERrQ/
dwV5aZ9G+5XVUAnOf6GqEJwyy1qZUC7lML+B+97kE1nt5hoZIMrffedZyDzfmOlo
olstyFodkD9RV6lglvnQDi39aTirCLuZcrITaj6l72w6XfkghrLJvfyzqnG3uSDS
CklSmQ6g9ceG8+Afw1Hy1sFHvRjRgnU+Nu0Mi8YNLYlj8Gu0YY7cltGPF3ululyC
UOYbqBAySkM7rVgNiXVOc0/LDFnpbmLGVX7FZjZHP+vOhaH0jyNWxenuunhaB0nc
J04rrZR+vXdBSJVm4BbncWycDAtAfB2AVNyD13jpVgLMh95uRJOoXRjvKk/c50a6
b0P8pLumXzWGUBzLg9iSHzhI2/v512zzOWvt8bffn3zU7GwaDWaPRKSOPyceS4Vl
yEZ/Y6DIa5s5tzbD9F/e/Isyosw4LClyX2WRHJg2gH2d6YvkQYMPpz3L7JwKCzSJ
ltPx8eQQaf0KQLZSOGKbHgNPVeAmRBGJ3IKtc5eBxo3MdyuKxoPvDshQV6pPf8/r
4sQY15gFdMmg4Gwditcih2A3401W6kgHrLOLlOQClQEcd5sM17A927HmLzUPBW51
peQy7TNJ80F8zt0GS45HhTMhBH8GZL/AC4AaUBkgjpvcBmYHdmC+yGQtLLRbrddZ
RZkzRYrQx7DvLVjHL4cYmT8GpMpM7740xsldEh5GehDGWk1/Fzeajo9OGPmA6XOm
OQ2TXlbqi++j6EyCoJJjgvCR8TmpFB8IPos082uQ0ouYdCfqVSm09NdRYB8LPV9t
hgGRBYrQmMHT7EU/5Zkaz/sGqbFjihTiUDur0ePlI4H408f3DpCw3JGXv3Owk7uK
scJEkoxn9H+HHemc+W1bZuSzUKSFPxzZCkDe4s5ZP13nL1/y3oxTcKrgsI9DaHZe
Riovo0H2lHOMiNoB4OgI5b5baIxFRcnZgeMgo5Ba+5xuDAJ8uG5cliEVMssJUCFV
pVpm1/97cG48DH7eTjQmGH4EcwJYLOl/f2jUQkYYC/gx2BagmKTpr7OdhMPTY0r0
WvRbciyho8sdzPvOzhns9uGckA0lnA6OB/A3UAID6K5zUxQ/Feqrj1zxpimZHlLm
Zx4QI6LE9LVvKKz7AhJrb5yyGMyUjT5eC9mTegtcgqJHDSGvtF+5s7aCxcenu45V
fl2TCUqsECpueeU1vy4iYZBwo/SXS3IDDCwkTxIkBIfqk6aLac5xNoOeshWPnfaq
/jsowrVzw6FAWdAKG3bK+ReLchtq443KTnliBAfad/6FoQ8992xAAqFZ9IE4mTPT
JgmOC9ct3Ch7x/05iL+FWcQ1eui8NH/Rbd+OkQqX6Fk0+YBqolKW+QhL2uelb5pm
MPidvq2yKCBPQCMydcCzWVBmhmiT4PrlZXvnwzCC29zVTbXVKMigo7SwjdETeGLo
DiYfUfZdGRmPTfc5A8GCcw5F47owD98iwO7uXxw0+qB2v/ws3tLPqEP8Q1XMpdMc
D8EDIT+A91oo2uGJ2/MnbM3mMIXWaqAsOmSAeqMVaHShOx4TMrRwgrnfw3kfHobe
2eF2U2pFzJEDtOj5M2A9mQjFaHvEJIzn7K7cw20ttm7zFvMGq+8HQnQjg9202tZl
ObK1uqWgOzh0WLSgZdNekDfPwWh/SeOoAI+hCItUNEZPmvvxZgnhUBvJcWZ554xC
PUVAc7kS6j5w/RcDt6/cmOCxC8cDbdZNUF/hmQKePW5M0jWMmiO/DWhL1dmtc4xk
IMsgBGGUBTDQthHVCckjiMY4L8/clVBFcIa4MdyrWagPjyjbhgwmgmYaMTKgNAPN
qPK/ZsHoJ65fP+3rVfA2uEefL1FrPSatUkANL4BH2l4NdNa5BZm3j9/vzCu6mpMZ
FttnFIhgOzuNhp69lvdOTfTgjf6ZgMgfUw4FrZXJkoQz07CSYnH6WghpETUzoSxP
4zrrDKs0jF3fJU0AWcIa/0mRWQSIOr/fgdK+LgbnARcbGMxjnVqt+nWzEB/9wSbK
D1okBvitPFvF/IflXWiN9P2OhAvrpbeb6lDPj9CY6vR/L6HavQH5dVx8HPJr90xb
jMjSqy2rkWRrxL6CDxiYYTH0UbPCAUpN++sV/4Ini1vsH05yF2WttXlZ68Iq9TCb
jUa2/yZn22Z8P18gwrDI8CnYPdnp/mj6IhJWezTeWb5ZEhBOc9fgM1mCoNn5rxQZ
yAClSEW7w8cQbzeml3LyXy+ARHUqWoKqA7dF6Jf9H3rgtCew4+mJKt3+sMtw4EQ0
Sj5Y1YOFHAew0xxTMU9iSfgtZtJTw7n+uzLF3huN3Qzv9r9y35d6NUhRRCSFjeWQ
rUOF2AEuxbx1NZMygenyhEsOVirly44J+znl6zDWNUiyvEG3xssJv7NUKnMKeIRo
Lmjv80l3/RSra2GxIzTYvUdGSZOsJ7GMP9of9IOGXB3RRy2E1Hbh8UT9Ty5HTOL7
f7uglSoqoovHODcsoNNns6XKi45+8OldoCpMBJIGG9ldAGKj7acCRAMVVjmd0WPB
g9/Pq1qnyCs6Nbv7eLveur4xMftWTCI6Lu0NQFcL5LavlLBpQLcd0nqAY8woEioz
/+8F/oSHeDdAPQOyTEBORXRF9R902mE8ZtS0LFiKbZ4zGiYUxShrDa0Nh+9RGK9L
VPsMBLM9yJIq+y2OFdaGgyOOPIDjPxjqxK4EaJHSVUqSnBWYPny6RJM1/6wkDu58
NrvXB9RpcyPxOkK2XxQMVOvE/xsSHLa1fvuc9YSTPnIYSR2s/KrimUDdlqFsPMCj
ZLS3xgMc7XA8l5MOn3RcOvSEcgJB+QEXgeo1slRrYVENTtBcYWJ49HljlQ2G6+vs
scoguGOpNGKJPelOaUMItzM5+IovhnyB2enFJqpN8sAqCs24t+qP08NLFbnWCOzl
c6UOvSPdqGTXg2f4Ph5HqgjYbTJtXXENNvJlIpyN6oCdpdqmllBLU+VC1iuCHRi3
fOEkc9imYJVhA5f/hPdifY2GXs4H8gLPf0zrS+piW4mhBhch34lqWJKQS4b9bSmB
lme/ymSM37d2EEnbK5yir9c8cjswWmrL0mMpWQrUuH5+QHtCwpCpPRyVutd2nJcz
8zqtOPizy0PJQhFs6ByhrLEuLiPLAiBUnA3g5TUhhyL29HO/2qKjBY4WE2v2npMI
3OcxzrAu3t2JXjBDBaWGHxjUk4YA90Xi1KWEOzGJq5efeGpzVYeThE1SEQIVFti0
Giv6IotRL2mAUe1U7+5ggw1Fj2yd/s+tHgAAYO6MAWfm0Zg5TS54GmEDrjU4Z40g
2vFg/U5M7Vqz1ZbD2n/x5Wqa0r+AzyiLhScBK9GD/8IGRAsy2LCLeCFpA9jJWkTA
t/DWtXkR7PxVRa2GSh6ZvyfkrYMGU75OJwsIYsIQSilkjjol16vj1IOmq3XYtgUT
TXNDsyvvUCSCgnVODAgy6HDTGdpSdLX4Z+jUHNcMvlT5X2tpiCbtPQrXLQt+iAzI
zwTzh7dqb4A+jcM4MXyi0UbScOy1EOwXOvXGAozcvubUA0jL7htBRY8CD+ReR1D2
p55cszdDNuhArmaOrKKU53U502gawSfcD2aoPTLcXS6WHq8qiV3lz5xD5aI8i412
FnyRdu1OE426Yfw0M4WQ1DXlXr6GSUQcT0PgaRavSI0VxZ21Cq0W4wbb9y1bfyc9
isqK9ufSdnpzfWxgx0O49xLyt17+bQEtPpsqqi8OcEVsVTdI5WfLGA/mbBdXDi6T
kuaccyBJiTy7hb2w4O3u3kQj4PVs7zhjPKqHC9fiCNpoby4WI7twYEd9i/NcfQnO
/cu2PLrKxN4tsufSDAPca2RP9DKxJN0ATbFkntmb6UNCaMTfmxloB3U6WubwsoPs
X+61tVwA2X6Rv2TeJ+lGYj64TginbPTqYj7NZCrmSc565Dhy693nibYFVj1Virrt
OiFrQJFhens7E2tPCMw8e3Pm0jeYi8YraE4/BAJPs4gR7tcFgjs/1Asu4nG5sgVL
2h36vnr8wxG+SopIiA27ShI0xjDUt3vSH4J6Fo5xbN+rg2cZ0CnMXPij6z4+ykX7
+AQSJbgzW5Xk9VEIUg672nqyPaoydl+lnCD6RExRRyJF78YXasEAhYswUxkDKOoA
usVmUQioHtY8dnHcskSxoFQkjLleoFy+MTTbrSTFeSbMMCNEZZpgenhO/8TBGXsQ
rIzN5d8h9LaeN80iPg3sDeTbtmNuVdqAkdndtE1EpxtxS/Xt1cetnj+hYYqAY384
+lMGIdRfje5p367dJxm943fRd1dSKgVhBp9cShr1Sx6xKCi2EyrjboN81bLX0XPy
Rm13MVZst98sIjfq037trCHw3KHW2BymStxzGYbb4jSDd18lx2SEeMrO9a6LUr1/
zXm4PnPAUt0woUs9on4tRKbRB7hqkULSUsvUKivmoDzpm/TtsD02K6CGup4YCVnJ
aZPrnxIiU71tU8ktzTu2xA46aSTZzK2MHTbFcywAuQIC24GafablZtyxQgRMgoK0
khKjfkCGxUavHJB55UmTvBoPsTqIMmmA7QvqHS3ByV3Gb2DOhDkNXR+ZZ4I9Uc2f
RTUiuI3M3uxpPkNQfXQJsbUb2BDxI1z48l9ADRksjFPpLMw8iJWxAW2Ky0oCRsxp
ZvRaWLiwf7TWNNqVxxoDyJVGO4/qYUIHD1CAJWhFO7wgt17uli+liGQgGCPFFiAg
v3/KYWaw/88B3KKAnMqyqbmX3SSeEqOoxraH4xD2Yv13KtvMEr1kqPReEz7g8Dv9
IKr5aHtunCcwyw0IVDUbz4O/bnUyN5LfY1zpwB69UUcdo42qhnR3inxQ4hzgFSdp
C04XpsCFGjOiH9sCYDBzTvroDc1HX//ExYViMJIn6EPxOR2V0RXbHhf6WLt+74F5
oZIYaDG0RISbJeYvZWez0q/3sAgpBabYHkQNLOLz3RDd8fx8Uv5Ian1YvtJ7v+Ct
/A/Q0gzFeVSx7G2Xa2nPn5F/bEvUojn7u6myFUsa7Yf4y1kmSOf6c9+p9V7yfUHX
DaZBZy2vIhQt3hjTrUqB7yK9MQ3fucj76dvvWRadV7y6PxCE7zDN4j8y99fGHxgH
mxugsdFez9//CszPu/mxsbbRN7bECcI6mB0o+Xfa00fzVbDoOBUCLLQnZtoCZs8b
CQfJHDnUP9NCs9I0AVJ/loSp/2AngHcFAd7zZhBk8UEtTbz77XFqykhNfM/JtjmT
aRnSSi2nKdNpHHcxLU3F0P0B0siTifVB3GKoMQnJUWIMdY3Lxw7+o/8noGlWnBIH
bA6SAX2MTb8pqOlkYDiqb8tvLVMpd7JQgbUBVSyBvWt23Xr/HhhsLhLTmd8LZD3T
BucXmpFvocWFvmiqwzVRKTC/wpk5aoFvlnm4I6yMXwr40sGV8CdBt+/taodQ56fV
hMFszwyc1X6ZrhAHEdofMPVSotFZM4FbrHZs/esP6+Q+A6LjcyzxYQVXRcX/rWF3
/gnQwpwA3RY8Lserl4nnG3bXVCklhpdmWlPn0qrML3A0rdcLuRafXkTApXcFPrvl
ZCf+rF0XzKq8NsjKW7PYTbsybsuLgxM2hFPjlI9xzXVXqLeTADAGln7sTEizF9a6
LuR/KOlSRW9YF37rDOMkIR/gMOM/CE4WSWoqTalG2C4vECL3B1lAu+hR6t1M7jbu
P8Rf+HN8UN2cyoT4AUmEA9+lCDp7QfjvLtgWxSfHj4L9vh1t1B3NNp+dGgeBDEux
SkOmYC753q+KjWoTye3aPlmwQgyGpTF3hViTpmefu6LPWDrQeJlOghywARedY3KY
PVvToLi0MNtaMtOtcNI9mTgvmGjl4N4st2/kOynWYyWiv7KB57G4/zS6ToXMvRKA
7YTr7Gq9LYEwqIZbIGvoUOoKOjEgNTiS28X8oxFF/uTMLEujTMMijVCwuRCg3TkK
qnSeozC1eQ3LVCd5Ml7047/K6qNvk66hwtF1GaqWRzb1A7cNllJQbwpg1F1JVlA4
TU7k7kGRivrxsV/a41n1NXLZJRM2VZ3X+GBKA/JIio8f4lTWMiwH3EOmBXG5Lddm
z3Nc3w/aerXL0TNSxTGowi0VnMnw0VHfiHqOEO0OHti42lJ3Fnu8WQDKU0FjNPIi
0+r+b3XgQ7iN7NcpdnZAfLSMeeGRpXqPZDf3p4avG0ueNEEvFwn/agra3+pvOtOm
ealg3/QPBl8OnsHPeiulUEO5C9Erb7aDvAjwPVdAaEe4EH2U/7N4ke+HiY2lwvlF
n7q3hHxoziVD1I6YBODONdvUxRZVw5Y2tJSvdwgo0r6m0JYI2c4LPxgTdvL3D20c
Y3SOUwOFjrqG+KZbOr56HtBFicIOr4HljFcl+5C7XYhAtidhG+Vy+qYh5Fb3RBHV
NvFZNA7av0N29aZ0O0Rcc0pFUbA0aLZvtrRLN/xlwAzmy2TtTv2PMA1mzL5O1ikv
qERRgG/f7pvXrHlliwHIbLWZamDOVt0A+TGLefNQeJHVtTedjgIo4vRDX5fPfNdz
K0NgWNqAC4Wpaa3GtaQTko0BOjXkxgrRArZfP2qkrscJvQAxjtt9cRy978onY39M
X/Oz6qybNLwo9sa3d32sunijgGkgxm9AsPvciTCwRYxk/h6gUMPR8VOI32fKkzSQ
JyTrcUMsoPj0ZNgNbNP/xrIF8FNd59REiUff3+b3l6fie3i29ShF7tBxpMNJd5TV
FKPPUyHjXghGQrzYwvbWXMToKxh/sY9PLqyc5jXmIkafcGtQMSng+j6B+s/WOg4I
HAf5VfbNWfiyaEm7GM+yOY08FnayfnymVC4e3RAxNuu9/zz+d8lH0s2c8qVAL1RZ
xxvM43CMON+RqtRoCyWxz3BedP1WnQqDdUUy2fpSI6lymMl78trOE6C67kLV9Ajq
EJFSKoUi06fLmv2jt7xe1r3WxjSaEU5dWkRjZSL797OqUbU1df+TqBb5VKqZ7YcM
Iqnrl3Oku4pWopwQAo+EgGHKqcEVq9m92b9NZxCE3Bk5OzQ4Xj7AMilQlN14ui3/
0uBG1a3CjulD40Pp0Q6sYCbdIghHrZGYFHbpVKbm/K3CwdyX87P05NRn2cP8QHZE
kgGZaHKulzxEh2CIPPPi3d5seskYfXxb0Vk41o5Wis0ZQAxzHSNcfX3wJ39aIwXP
ZrzqtUaXRFLnGiEWGLTyUo4KLSsrcr3h0JEMzOLwVDjkZovTPM1WQ2F1H5RyY43D
48gbk2pM12T00Mt+GtV+q+5SVV896/vE+cyhjOhczvJA5ueps2CF1PCO92fVktDN
7Cux/ZFgmRh4ZJ9YIkRogr/3wV5sqEYZwMEuXrWIDG5e0T/XYW/3Mnl8IA1wZMiH
octVj4Dbu/ASco4Rt6U6A6l7bIO8r16zzrbj81s3+ICzNAnzjYWJJKROGQ0t7fM0
EpDsf1ArhBN/JXiOlFWLarjs1xzcMPMKjnXG8NynuJx5B/80tbdegaudY8019Loc
sJ9KjOFHBn4J3sH3kEAY5hWByJI7aZQHRu4Wnvqt9BSpbY+WMpV1uMlDOSZbWVSt
3aV6ifDb07e6O/O7JPPosDvzUJvlrrOrEXv48Pc1qwxRuCXd9VkiLsJxFik5VfVf
IUIvz35DtnLX871niEsOHR1Ftk79gSUpD5z9JS3s+AezDSdhPYmze1sC+oS4tiAW
UCzbOBlU7XPjZWvYv/vzJIZl4D9psr+aIuzliXQw+AZMAQUugsK8UmDoDtg2AEpg
I6qCuocoZmYh4jWMTwNh69v54W0377ZjSmuDHlCqsEhplHyc+EmjIkz+iNdzPkJ2
nPGSdrw5XtVZFfDFsA0p+jY5M0MBh3ZCPoqsALR5fA0suvIWmXt77zojUXEP1av3
7gsStLP0bs5vURDJhgfsqTA9efwCBcOSZP23ZvlSGTuBp6sXpiySVbrHcnnH5j64
8u2J4VtEa1IJ8s6PNd0uEYhbr3e1fqG3XJCH+3IujfzuHl4GDsdDhGCT8n/K57no
+qW8xI+A9LoEfFZHGLYGUWgIAtm5IzKpg7gytQYtfcOeiTsDJTg+bmYWnhOqfWdP
9Xos2eC4aY7EiDADdMB+d2QIgqc3SIwXUeMa8+9Gy4bIeGQVa9TYramfcQVtCnY5
cLuwOLRsJUmT+uwcLPgSnx9VJ88QNwsxxeN3NM2pRzin84vk3on3q8Tj2bhr4RhL
4ArgqSKMPxz3e5rHjMUTdntS/pQ8SeCdxv+9JpEu3zef9gIHzn7Udf3sgYdeMbXE
PtlChouxcys/vHwdSJdhhxzcgcETaB8p8L9EbLs1jpbPqPikVUVOXG7DPum/+icP
q7LKDo6AoTgw0Kvt5np9jLoomxbNk+pbWWpkzo2ZFZONXn+kV4wOsnzCdqOf7mMk
3EgLg9bD2hcNETVm6jllYPNujEXmJL/NAT8TafCGO7OkUZ4n+q1KQC8FrzeN2Khh
YFF7gUwePH/g1djl8x56ElpvkjbyDvVVaccOs3cQTXvtP0dU1LYb2OQTJhGOUUEp
EmiyU1BgytsSpulblpdSHQJjFesbSwQPzY1OsBUzO6VK2vMBKq+AJc/1ChZSA0s5
LW0N6wCKK3bo+c7TFZWSnmvLHCmaACEI9R35wGgL/Tv7t5EXr5nxdIgufqtIncIS
rIHJx1kEa5wiB3i4bAFnDqI4OGMX0ScV7lNCP53h7zq22vTA8tulFwiGArFO5cC8
s3CqWLAGB0+1SVsyuQEJJ8dOqVueE7hHFQdC59RukYeA9j9w+G9Zlrxr0ED/45GY
ufNvzEamm0o8JcXWwcVSzt1DMtZfjvUknXfm9vzSXxu2nzTtZ7ecemL7DLXzMFXN
Eszz1YX3eeWSZ/3pDtCYwjnctWySoc11c8CUYIHGpBpi/p7fLZKRTO0K9kKdbGLY
N6IvY+/eqEWWJYYrqouW2Mctrlyf6+bv7oZUnYt7qfmbkpNcnQLsRdgEC32ADZAR
DgZaGHcSYr5SlR70CSCFHTcl3oHwYWWINg8N/eWxQmTPMu0Xpo+nzPfedH4HhSGI
7AeML46KpcIqmWatlzO96dWXC5y4PocmFaZpjFH8UjiQ5rRqZRwh8maFn5Is8bkR
HQbZn3jseEbg8tlXzqBbKsUdt4WZikVKdksu2oXql5tqYmKmmkath7rrLPKiGw1S
UbJhWxSZixNVHdF5bUDvyg/lk4wLxZOZtRznxe8z8UNGJxJ6otkT8wiFs1ujC8/n
qtwJT4UzHVTYsj/obY24/LH/VokYMCtSoLZVmoh/Mf/QjjL3k6hztO6aXjvOn8oR
B2nMoXgz+8lqKJV0qbIwSPr4mTzVhTIEq8s4/oSJFLkClYUNH9aKkN7F3rNPV2Mn
DilOZ68dPKAQ1hPMYTBGtujWvWP35/Lr7ksJZHJ87Y6n+ucsHwnFAh+406ZkICBV
3cD2LN1K3dPS3duBigtJsgZ6imN9KpE4q6n0eb9lgiX+Aqk0dxk7rrShOdKgKc2M
0zRpYU6aurLEkQdPIgrqF1YSrUZeIEFXk1tqatjIUqlP+CRDZu+RxcDwWpil1eVF
lVxje9LwkaycgI41oosqg836FCREm1uuNU3nhQwuEozQ5gBiLmjS9MoVdbkV89OG
UI2FUSx0HGQJYnK3BxKAZfGEDcyymk0k1CIN64vtAXDN2YUZyLrVUlGZGIcZiiQN
BPfEZWc2NtqNcFGF3wtqpJsAIJwECdYWK3mvjRN9pR7EMRc+kr4jqdeiPfhe07O+
84UQ/T3tDQoh9E9QI4GOUIGNRBw84cj/Fifg8TeYSZa+9pV13XeajgeOs9S9ra5w
vTi/zabp7r2pmobbCk5IMJcJSuHynQvVSocFH+UArRMvAqcm+fOLH6XqvTxTyCDl
oNoAri+gAKasapbxHCe+vMM0gD7KjMz9q6DhCWMcuo4aCMWE4xgytwQMAUZoMRuE
jPBPDM965BJTD9u4fY+o0lSYa7VCi4wKoYDjjg52L8pVHarTMlPC8vSweJRFMjbR
Fg49kyaYgm4kZby7x011nEzRl2cSthun+vzeW4zJEjBC2Hr+6vZd5ek3TK7hBNNc
nCiFzYrIBKhqPibjFTSHoSRmlilE02mTuaxo59CuENnANqArO1cuBwCVl+Im2NvN
tBpCDhQxt+1lmoPGZLuN1p67FMjd0Rq+OgQhBuc+PAAEOptNy21wNXit3a6bv/kT
aTOwb4VzkNj5kcrujBQsEzmOf8BFUb6WhWYE5wiA0dxzuoK/LlbVL+tuCbM2oo1m
FyEqIF/33nDtxlFBlFViYZMQIJtz/BEqdLEZTHbDXIb7rahuE8oJvia0lrrfzP5v
3DlrYgtWpm1s5T3YtC21TEChr4h2eUiyvlRAhvwkGQ7IXnZL80n1JvO1BVRL9KSK
ggH3cdJkaL7ZSeHHwAEbzPblnFLMfmx/ueNyXYiaq1fSAcsBuQ05+WJz0+9in7/a
rBcchbgxZv5fe3BR9AHwkiJYgCQWM9TPXn3djiMnrzj4o7C9RvNVq15j/eQt4bOu
TjrAS1HSfXmssuKlG8m3CCJ8wtL7b+pVWntvzchmpLNK+iO6QOTfSmoVNRGHnSda
LI0TFSyoQFFob0GTQZJxb7aWww4/vbfGAawdqtO1S9UhDecx8rk5xNygC9jaSN+j
nMXaJKPThmNE7t97W0p0IYjYXBl2gsbcilAD4adbr7CfI55aS9Z1GRCPtwqkP8iZ
0Fj+ScaFzMyXbgKCPPTwOsBqfy0cp/jVMDOhSULmxMedJpoT9VWDwNp+rBkxz5Ew
2hCCH7W2N+1tOvKELWzStYoKghENUIkLlaSLf+J5NrCtWVWcEinBbZlt8gw6Qx/Y
9Pi9/rTuXZJG8/x8W689Ts4Q0CxCwBOjI13qKWMGMOKjwm4C3gEiOOffHNCuDCcd
MZThV6ZJi/iPYJfQCo2sFjrz4A9e5JAjbFZRQIWkM+GP8p2cR4ZytqYo/56MucUq
c1CROdnc2JM4GDkRMc/g1Sk3kmBezHEh4qTX3h8o09+Xd0VwcAmESMWBZRfZ1wrH
ZFjGlM7V7d/J7UVz9eg1Wn7DFyvXYcAbVHFaCZ7TcgC+4DzDmad2b0U9Wtrq2jBK
K2wZsym0W/VW/5pJYcpBFblfoIJ2iCAnnaHrlPVM7sLBkOuT6/htMMccPMq4zAMO
xPv1PTQP4XtmYbmAjhFylgrYThnPF6lY/qShShx5n9UHnZ3A9cKv+0NnO4Trpy6R
DdGTxc6Ej9bbMvPpBh1hehk0YQ4HKAHGib8YzZ5PTDauZSJITgRGb3Q+cmy9QeSK
G61wSOJxM2aL9ODdlWmR39nhn7fcAjSb2CS55acji7Q2OQrgqaZmf6qtypNrIGKa
358s/McVxEVinz7lS+PsWpt3MPMe8ERdoJEN94OthFXq602HxnzxumVCGm/d0EN5
IU6zAjoQfkalxETf+wW0mbd+hiIGKrTX+gLS/A0B4U6jdbmr8L4ph/qf/sn7s24c
4kX7iWJmIiUZh9WzNbyk88w1ATmDNtswNrOkR3//Q3G8sZcgISORPvY1SHfNvg7p
GrYFy7MXAqz5f5WweBDqYWVxTlsw8K24yRJfrWc7hooCVO2kuF0jy9w7ZxTF+b1J
jlxWunVMMbenj1NzkB1CzCvudgSEr1vfiMhyXp0cpy8Am5Uh64YebSP40DiJMd0s
GLVGr5PUHF3AQynBnCcNkd3kURa7kOele3hlTZOfZiy+hEDUF7re4WHgOV4ENRgt
VtlbGSZqVweEP649jZGVUc/C+wpqQ84XkPpY0scw8bCgv/7Yb0U2aVCHJXLV6ZDm
4L6MKrWmTDkMupsY/JboPoFkqZ6tjSCYRd48IOXBInHHVOm07ADsSQqf5uo9zHLQ
0m4lgldyViDsVfhxYEW6yJNEtz6TJzNeGkcYw5JvmDPU40ce0dKo9GFpEPD6sKtE
f5DyP9aG1jHtotkpvt0ir+Gfc9IePyPz0v2TT3ZWW+xGk/mPUYLzB38UdLjWgBOI
GGA3JKlWT0sMwnR89eUx0ZDpv1W0bJhOUw9wba+4+3MMFvRXowjO9lDhpoX94/66
T4Glu8uvZWFw0XbRBLrUFM0r32CJnTclZ4M2IdX6JPb18+nIWJhE4HqUggKq0Cgc
e/QKJtaipqixdSDjO1Ab2mQX7+kIFSNWTN5pLaPHb/EOZn+FhYfpSzWaC2oS17qC
Jzc2srP76FmbmwRF7xz3t5tMrcka7qH88sCaSFvE6JxnMVTxYcm8Xt3F3yzI4lmv
OcEf7z58acT6McUQT0cWpZk7XfJvk+5390Mk3kBI6bgSfU2HXxtBJUXP9BZiH1Wz
PlOZs3WgcnX0PDOwp6Zq9rANyDVLMszdu7c8DbXBfZiEb5/YMq0Y5Ei8hCEQX3zB
ToZ4tzCkSxs/9ke1/yNeXSZdYZKDTJwzbsnWhkzhmMWFoDD8GLBvuPZmoQ+Vza/u
V2PWeT5wat1m6fxDzBYQW0b8uXQvA0aiTKcjjUXHbcRk+gI8H7ZlkNH+8W3sx6kt
ofJz/M3bxjpKQl/Ykuitzfy9MvTC5aSHBUWSuiHtcsZ5Li5QjrjoDeXcLJmEWvu5
6CeoTCju0Xf9N78sdgodRkjRLoGOLZghptzm8RXRxmpKTmywbBPMvr1+FNtC+deS
ocOIeZel/RofhTeJk9Sv92g/xmYE0jGet7CnxuQXnFqCWfnr/b5T7A3CPAqCfq2w
Ck9gh8nFXDL3Vx+OE1JBLRYILEVvkeioJx8JwKtSccB5pZa6t1sP7Ob1XR/52Pl0
NO1PlGgrHrHuxdjngG6rn1bUTgzr9a0cK3FGd/AeTto/i7JGBRzUfjI7sz8zs0wg
HcAOTXfvzqV0EJxYk1ZXPT+FL/iQHTOZNRWDDWBRW7kqGhqgPlKp5JJInrCqevqZ
4/nszrK5VLTXRZLsQzcArtZsETJo2TrpyO3/giqEtsVatM16bpp/dN06VHfuN98y
spCrmccL0YtcJU1AyAWXa01ouReXt63GjUUuROTuFLV84dXPlzIL8pM0AyRw02tw
cLPIRsNP2DTaJYlfdybFU0NUVN6nEA01XWwOx43aCS+4Jx+uQ4mBVKqD7eJvP0OU
gXTWqdiqCs+JMDzyt5zV5D+j+zx3AO5QBBOstL6YZFi+6xm5MId310pCnYu2c6+5
iCtrynUNw4setxllH2VgdT6+X5nqqGTEwZW9ap480a4I4lPXcxiV6wweOajmS9zy
OWr45fIzjlEsZUW3u2nx2+IPu8VSCzoTdVzJoG9R7L3uFtoovPt4R4dBcnTo0Sql
RkTCS+e00dM7L9ZKR8tBh27opYY+OMoqjaouBZr1i/eVbm9ea5o7+6OQjxm3A5w7
foQRlW44j5VA3d80qv4b4iP57oRZ80bce/rjUwUONPl4GdUP94PTKb0ItoH7VzyD
zYNbySDvzXJHz4nXzBnsPnlyGPictdG88jVUEP49ybz001ByPAJ4SisWtaXUDZH3
3QuUkgxmAwIC2odxhAXEWxacGOiCgtvLQ8q5/mvOuluZbwm1UF5VkO4F+ZvnYdkQ
r1652zWyALvGANiOhKuphG1VadKbKIYQxTNvHK9QJmnrPKmwSv8Klsu3Okz4BFo6
QowZwZGPw4TPz2GZr9DjusCqClPmz735+vpQJh5b5c3prZ/d06CqYKcrBIIox1YB
PYGT7mMomJRMOe4tlh5M8rHWGAUBg1H1DP249dwRSjMuAhbiIsiP1bwHV6sm4cFC
ZPi0cNFBKiCx84SxVUXnLXEcODIK7AEVTxoi9dLiX9EyJEhIlYd26VtwsnL+VG8e
fwSXcAGOkfKE9U2tk6lNAMo4Iy4NbgI2VoFAlZbilC69FRXXLwApL5XUjEcsI+Qb
AtQek9fzH7neu94eLHByLPZBHW8kJsG2Gz5zNBXY3KNW4CZ0NPjWF3iwSOwVT5Up
VTQFoSnCBLpYXn4ngbJ6yrCgs7X8v7NkmJwu8GqYrzTBh73SqpQSZVgTNJwppcRy
l3YufvF30+eS5M39+4Yu21kHssQWrM+CacHg7uvL9jkfmU7bcT6qzco4Yop0Cqpu
J9w8XGGQAYFU7WDyMw4lysOBICPPIiKhyr/m5vu8d+SyahJ3LsXFJ4EZe35mVsL8
Si+OjC2HBVSyj/e4tu1of3oW384/aMUWYWecXLPKdVH7vVh/HD7cKxgCCteoz+ph
9eU15OHGDkFRnIlJcu1nom/xXK5VxE4gXhnzSZgP9DZTph4S3sGRlbtKgGNN8Ep/
g7+xAywIaC0k1lZwjqDNcSR/P9+uxTFIIz+Kq522XNen9z6lfnGPYCzztSOIPr4F
j3Qu8qvzChLR2qTQqeuqevO0hPa1Bd0HpRYNvPgQ2lk+3HTRpnNXAM6uwNynCDtg
3uSwCsQQXRvoJN83+wChHTb+mg4PQeBJSjdWstqBf5d/g+AXGmWDO1v3Y26a1x6m
zCm1WsqnRfel/vYm1T0/SBxKOjhB2Hxzk58rzpUjbfh0dWtG+XGCzySdmfLPQq7I
+UFfbw7ByCxML5lsKHaFUJg6KiTAR0zLMWwD8fJxLyzBsEfyubRGtRDn6UJ5MME4
81kgxFT12W50X1F1pzDw7W03F3r+B6Y273XNI5L18LelJXeqbsFT9xxnNrJdK2te
zJOXrS2+xmAzEZctqFM+v1CZPKTXnyZxzF3yc7cDzy1nWZCcN8WIpEC4QZxLrPjD
hg8DoaArIygJZ8M2eOjunMkIOLk4JShUvIbQGI9bx1WaYp/LDOIV+6M0f9FbrVDb
d7Gu33doOefmBEi+mUBhZcaf/XIuoUm2TWJfnZEC0FV0xmQHFQsV2y2IeCrsZ+a9
557w8icx027TiBFXMY0vX+Xmwnu7f05/4YV39a3XYwQ5VCAcvoN2LEPklzVP8zKE
A0PoCL7dvUCBvTtHxkrG36ixvY9zXe/W18aA8eDpGb7mr2FMSgHDrUHxjmUtI0+k
h5b7yJYbdn5hnOGwIl//YH/wd5sGzRRKWOMl85bI0nj+2UoMDynBfQfZWNkC4Q0B
ox+ayn6HXfAEeVlnMJCnDi1mspTqULmcNItSJdTT6O4Tz9yPlN9U1fUDRJ+as4pW
n5+lUXBh7T2e+52qWakgcYYM7MqEAT7Ke8OjPZx0bAxhywqW+LpMP7dL0Amm9+f5
uo/Q/EyW/YyqIArgDYjOdtl1QFhI1HpPoMfHNTtjj8rsDcalX6IPZc1Y1DeEXOf4
c3vL6tFlOsl1GHHMBzOmNFl1GmvtUxL9IGb5R2JSnISDqAgQvov/R23TFbyhLlFs
761Bt71BJ+U6urk7MIyI0RbsURHkiAN3ZmlFUUFMa/Z4ObLuVs2e7GNN9rIZt7gw
+GnOrZ47MI3Yh+REFp/LnSyGV7GY9yqS0dwPMIvRKbYFDLPjw46rF7ys16UpDkZ2
m1eVpmS5icZImVUvO7fYFPHgZz2uo/imGvuEvGs9Bu+Qyh0Vkw0q70RY5nE8ysPG
/3aX8c3biKFpU5Wv8HN62P8HKrgpun+vQOapWBeF5+lWX5YMf/djQNQ8XbMAoELh
mXyS9XZmrT+5O7CU+jzKZ8U8k6IhlDJdyxtbfGW9by2p6tI4IiGdYBLq4wPTdWIW
dSrh1V45O20Kjx4byN0rOssPxcOIIxnrfAQNDvR8FAwjfMMHKFxXjKewpAcujgvF
Sfgqric04bvMYwdfDhBx1wjXJqk++iPEhmJQ1Tv7jsIyFAyl5c/zbHmxEyA9ISws
/m5XWRHZt3N7ho5v2mAYI8Tbepm+0OFlX7SFnP8X9k5AjX+Vi7UWg83+b936aX1l
7YXkMXtddZkpGucC/g2O0jVKIHkcW2+ZjQWkpuCFrqTUWBkBj75cTM9AllHTDWV8
9Dq3e00s559WRzwz6AJwo1xRmxoQmL9URfT2ct6z9lij1BNJcycnKCJMfP1hvJyV
cUMg/OC3quTD/S+RqShKZycDRRoYNGC2Qq4ve1cu0qdD/ALq9B9dKTWs+EFgwf3u
tnwfuvRkKXG5ii1kHxT2NgW9vBdztk3wNzMA0msHRuCWf1MY3tWZYSMdz+aN1kIg
HHZFufAnHd4kX1ShxvQ9znZEnqJu+RS9jBK51P0Kiu5zOgEQ+1wAe22lCX3PXB9Z
ap65fz6yCco/md/vgPmWV8WtHdUVLuDB3RrLamekoAnV3mTU+73EOSK5LeD9xQWY
Lf+fpzk+yqq6ZqbwRlIN0jH+lur1eUJES3JdG5r4zP+VjPeVuvu5es6AojBs892Q
smgK9w80luTcpOse61YnyZ5SdupKvL59spNa5eYXnwizkOHONW4ujdaUrOEHs9gT
GTWNlpUwF22KDWQUHwZkiXIvRn1rWkGPQcMlMQ++RE8BktRmBoxW6he7li6UJ7Jh
+j0AW9ZUmDvfJfbqa5t9MrOMJtmrBQAtPlsZ9ngaT+M+cCvx+4VoVtBf5J0+qFmn
A+EXA6zbmGlu6iaW/xbCNFyGccPQ/tE9YQrLtw0fwuJBcDo7YZieZQVAm6SW5bRe
iryiuzjhKTCrvyiaSVKNU3vl9pA1gCN5GWJaCj0+yqxOolxcYXdS+ELYpfWrxATL
QrMf1DOGJ4wSApaXTRBveVr7QbqM1AqZLfdWfEGA4JADsw3s5SvuhdO/m8/p8zWr
i7hXoMDxLdejB+fCsNwXnEnRZzeSXQr4bIc/UKq4ZOz3PnLhjLheX/OWpXN2pF+u
oUyWoNYpi8XL38mUlHNCEWoLudnxmQrIoHJAnMCavkmy4NbCXiIRQUvI67Nl5wZb
ZKkNwlyOudPH9Kcg/QqePdY22FpTN+ouSquGTRxjlbCAkQU0aUmxgTGy/atENSOy
WneUOTOyHyDgUKOJUwPj/CmbG4Ou8UrmMilhokElpiFf/koIk6eq5MwwszCg5yXJ
l2NI3fF0ptxBepVD/1iddR3q208UYX1ybo6RK3Eah1/5NYsiKYAG9cNAhgky2NqB
1/PA63CNZSPf8c3uIfKAstufEBlLUkaIb/D4pZ9gjk/VuC5DEU5MOkj9GSwkZJIz
8xF4bzmnhtB73F85Eme0t0r/zRhpSzFicDujueg/xev7Q7RduTA/nBat2PL/ffta
kgfbGENrZiY2XtS1cXQIqlkxWw4BgkYZYLqiN9+JySR5mFt1sDXRiG97yP2ZEjvZ
uv0ODSMtiKaCFqvhM+i6q4xo9d8HRMy/LGmB22u/Or9DY0WezPcYvJvL9O9VP2hh
/nDVwKuVgEQDWhSqzpY/i8bvv1LLnsRGll9KvIc0gdnfKO80t/xn1B7+cKVwxZTq
HBhVFy5wEZcMrqFUnMaAInavB3W8Wp2mbnPgh6Y+8pkg6sWxe1J8u/Tup0j3aIaM
5BMkG08v0C+lVwCX18o86hnPCHT/hkrutwnOgJosFqRfjhekLd/2HTIibn714b2l
5gDvicLZCjF5WJc/CDkfydC5O0jzLSwWIxXpKPggRug0TeTCavDJxOx7iGVYAuLU
Gg+KJH3e8aQBSe8vzAIJHjsc5BkZBjqrA6ZAD927DRsqwA3/wxHfLwElScyEO7BO
1gSJh4srGPyx7mCFee6Ar6FCCG54ykjVieAaRyttA2n/7B0cCco47RhUovDmm1aM
N80ViCaakFfzhU4enry4waAPxN3FG09MTnIQJ9IfrJqystf9WrnDanYWvpLW9UD9
QmvqBQ8iPrwOgwsnuZEbOmSU1jcLb/T5LiESisJ1VX/RMvi+oG3kF+sAjztUzzyS
YxLBX1WTKavyvkGFqMtERq7LvZo7ywJ8vXEeFMJGv2tp931uRI05/8w5ryzUte4l
RVY72ssEIzAqjBwD2PA4xyLbxtUHMY0iMit0g6QU6vYQj7jS0Tfgp/mfLSlV0ucZ
dk51yHnMGsugQE3SWFu2A4EhgkVAxxc6t842qXRIMyz3mVGqrQ/ZdmN0Krgk9m4h
qKv7Z94cfY4I5T2aRE0li8WELBGTJW5b5bZCW4ValvjtAiRbPYOUbNuTkDlVMKs4
pgLZo/fVvffiPBlHwSXeRaWxmynUjxR3ZlPQalirVaXzULvyay3nFTigI1fQCFwk
VvE336rESyQMAhnzyQDjmIJ+X5Rwldiz7ltaKG8mL+VkMggDo9UZwCMjEnGgwgQl
P79PYxccj3szZpUiRCapHuhmz+i2ujMIcXzShJ30h/vNQs6rOzo60QNfrkB3X5hg
2SJCpDJap9hA+evBtTWHT8hiReZJiinVWuzXR/rJNZNx9ISN4iwXdiR+djlAC3JB
YaU7KHWPEf3BRthONcjFBaGAUbRjEMKPqsQd/gclOUywW51AJI/tA8nfijLCb/f/
yC4sciUSSFSE1KJ4bySUNEkBNgNXZE+4HEYXSGhWakINOHfusapM3zpI1P4kTxuR
4vcjsMFDiXkkGrEItUusS/4qlGsejc5j2AP1+Rv6rDxJTFP62EPL2e91wcjpxjeH
FOOwfkrleMRNZ3T9KmoTKb0UgQ0Z4HUFQ3bOeHPAfk0qecWiadwcNHR+88/ak1rb
0pvSiEnIUBKIxGgTDJ9DXe32j/cb95iVGC6iW80n3batnRrwRQU/NRrNbX/NZ97E
OHZ80PwI9edwU/ZjV4wEMHLxGR0SpQGvO1BBBZjfXIGnWm04A0Dbe8Ps0UZtcOvr
QzxG1k40XmdLwlD1zm7fyZkqrRkMYdLXYZXt02vN3BsnwPOFoLGPqvzIulXdRpF8
REICtYHAPLjLB2F1RPvscVFuWnEXuZH/EZZA6hZ0gngB530WnUKk9FcC+1021sv9
/NlnR16CP4KrrNrDjsPqAUDOjahC1A4wnz83EZZ/IjHM5yfa7vu1Kemf7ROKL4fI
8A6IuedsMhBMog2JaJl/OT/kReklGQ1SJkiKyC+tjTkPwWuZxXIippdS+Zbep+F4
brOzIqks87sPEjlURt/iPHc2JEBjjD0w0XjGrPyNhSedLtzu7epgqjTnxWeTvuGb
yLN+cThNkM6B4oN2NdjKYcu5fTi/0C2J8IG8lgXkWnUF+oRRey5gL4tlen4t9Kp8
ztRdbEZ3a4qiZgUalPAIoKlkknBpKXY0Ws3wr0Z/w98v6PzlF8GBmjFT48OJqBxf
92aDEoG+xF3DqPTVq0yeHXbxZJuQnGyw08/jD7FSYIoZ8pISTDsPcEHQk6m68Yyp
NoQr1WexNvzOFCTDTcU/QzFLeJ9UWY0F6TjPr2aQmZIysMtbjeeaByq1S/f+tT89
uUUDlNcGnIKE2VbU3vkjRnH2pzdMijBKA+qiUExs2Gq1STJhk17tldbsG05OzKy2
u9K8A0rkgvwVfeBgyHJrZU3UVL34JIte1uM+SLgG4ha4zkjbwypftm3UFDfjUf3I
C87o97Gj9vyG3U9cmf9SBKpsoMpG4we6e2uzA48i2b0ULvN9QAkUic2DsqJQSkcQ
4qpstqP5FscqrE/kb1gE5/YezT6qTxNBBzFDtgOFv5D9TCg4x8OEvac3CVKx10k3
Ss7xrS3EpEaAOl0ZbF6ezXk/Ewtv3yup9I/jToS9uQBGUUFqv+zasmcT3Jmik1EI
NQU1M8jQ4eRT8JzPXUO/WZ5UXGJY7kQ3nNq3KXQQ1rK1l1whjidTOhqiqpynDJeF
FjSjUrmgvv1N3o0JCvBFHYGMT7+ypr1SceXDoo/HmtixE8C7qg3318jp6IVBvMEu
86uEaKFsNMhvpRzBX98IYZNMsy2u32awKfWGplJ5K43cGHfbhSqfkLtj/IXSIaHH
qHaSN++wxoZlO37fUFoGcXyeYdAgPqLrnjVwho7CvQMlqx/u0r+pVnu0rarF1N2l
FvA5sZ0mT+ePqKoIRYyocVdKCXjthf0fGQimH9UNj/fxVcqeuwqmX8kOF0QSZs5I
UyeLpG32I9YbpsNA2UQC2MaV6jMN2IqsV7eiyaLxpyAsJ/dwK/U624+E82iaFKej
z/KAQs3Wq/PglRXf1WLfUHkgj9GvifXzOpOEpbLSZx2cwl8ldP0BCW9uT1lvZ6lf
WT2khyXKGcnsVT5MQ9k6RE2/7q4wGFA77pWBZiWom6ERS78pAGCXTpw9Q6qyyoWb
Ebt8X/DwznsXK+LjVlrKA2rbXy79PitOOErqWvJs2qsSSDo5VtOXYd3p3AT9ScNe
ys2zc/NswY8d2A8JiCYUjk2rzOOLPpT5Ql8s2573YxDoN1Lt3k8U06LzZf5UbKeO
/DP2oh19Zsduo+G0BOHw7EX+zmXlAHd6ZxPDp6p5r3Zacs+OiKA0a1rrLPNn6Z5+
PQqD58feNDDQNBrfyua/x1Dbv0mJLDRZcl1AtNVqBxWyteLWSaiSjJaf2GXzGKK8
jdmKMeC7Yakwom4ix8a3H3wGQCFUJZ0n8SaNG1ZP7Rw/NrC09ICQG/GgD5sfavId
1h7JafJyl2uU8wh1Rm69DgtLUS9Swg7rfZ2E2gjDdG18HMuFVKjlfg6KCqM3ec7c
4zV5Y9xbkKm7IY7Kbs6FY+mXKxCRy312emIfhXHO0kpG9njxCgC8qxLDxZtEXl+2
rh/3lIhtXveyIy8oO1pmTtJeiZtCbGbp38I3in8FuB49yVLzX4GgWrxu/6tU/O+N
Gwy04iQqkIDEtukknlsEHtS9mmwkEwXMqeD7gs3xEjZjAFJhhqyzDGcuOQAG5i60
6GXhydSK/Lx266tufAZ3xOv9pcQNy0PB8mF0npCOvjA19C57JqDiku9idhBjyUgx
jjvULNfwALpJcRNRePOh/D8PMKSHPgMMHa38kb+rBar66VH7/92DSqTZXVDFG5/C
/Gk437b552iTb+h+Bw84xAfE9NSHjdSRkVexstiDE4G1GULF1F7JtybTP4EmXuxx
UUvxOd3b2KuRNV4RS8WodzV1sZ/xdFTdalscLFDAfjnSS26F/nHeTNsPMoaaZVPk
A5HW7asoDVlaDxIxtqrQlRAEcHtuQ77Slaim37gDDVTbhZdieYJ5gJfYOYixad75
yDfyIJ2fgNMaKMh4d0vx83aTZKm1Ctx0hIEcf1h2OG7SJYj+3znwIIyunj/uTo/O
UAlHBAmOfESbdk8VdVZlXdUB7lT1m31Vz2cbi5xFAJ7qUbb/DbX1HfF5XfjbXaew
CA497HTXw2Rka/Nr6x7UihkDbLJ+18Lq1i0+Aw2m0nFT5rHxEwmXVuhQYmH2M0Cz
LpnLbIDLYDPUtz10GfwLqhmWTIOQkAIvSdh2iPKNdABQrNBrcXKyzoB+IQQHSfVL
yScQ/pPKQ5TAXDK47/hJnVJYMVKEzmfAM7Ygjwv9DR0RYigMTeP0uXfxj3G3vRWm
6cWj379MPi3YrOax6gsWbcucSj4ECtx90EOxLlzpkPYCGv10wN3qcRTW7ViAzEgk
GD0RuYL5aV/FIyzmSIiGMalYtRAJFdzjBhfvjGlON4+B/f9njQtfoevpozifEdis
m5Lx0c5VCyijQ5dmWl1UwLQzFZwS1WLrnzhfO8azYJcUr2y2LY9YPB/eC91s2HEg
2CAbF8Kt593b7Rk+T+y4RDtEAgG/WxhtKDuPyYoCoebV/uJ8V2nUy/oICk1wfV6O
mqNXAOl9NAO5YU4r+BPCAwvO/998tW3daJM62iK3oQcQ75FT5qyFlaz44bK8vr5o
YUK/TeGK96FV6L+Wwzy8hJTg8fkEzg1ibtBld3foUQA/0XTxppKm8w+D2yK9FcOG
1uZTcZclNce2N+jgH5+Z9bD87w8lc/pIgyDF4tcPXZNrVJLaAVUn5itdg/AusQ1l
DddqIBrotGSty1ka7e15iCw5aaagb3MRsFksnw80zahyZabOT1EYgZlCN68osEWu
XKln47JLS7Ixk5+MocWq84DxaOfxcEkhRTEqq/+77Z12a8IMDpRGilqDsgU3BDDM
KC4XxactRDYgZGzJ9lkpn0BapnIH23eOESFZ8OxoUJkUPxY8TAptSq5Ro+/71F07
bGjUVSFSkaJifiPk5xYNSAGBCbf/GrlyO9NnXRBdTvAJzOXb+3s76WTIh4r3frIP
tY6IB/NGsJJVKda0h7AIxc1IWJYcoIQf/KLk0obPPcQfnmGXVjDoISwLAcqixwwC
o6GgGN15LJsksTXGllbvA7hW4Uza6T+ZTsNo/C1Am4ySdgZzHqMQkHuJQGqDS0VN
+Tcr1liog9DDCpsPBeESRwfUZUqokTEkJ+qHQgL/cMUQMtya2Nz+Lu1044A/ISej
Axai9Cit1d2TSxJXAag9dywzgbM8zHFx89sxoA+xU+x8xKgcLCDHKAHnjdgeQgNV
qnNft4hfjmo3FSrAz8M7GmqDBXCMQ9i6XFFXMGNV3MFHWomUjMNtY4FrNX+gcgj7
WRKA9dRRkjU0RiF92LZF3IXQJyWfszZlDMz37XmW26KxOjTYZlfNztYZ9Fz7hU4Y
3B+SCbkT38Fq7EdE7ZPro5ItuCoPckwQERtZZxjCCwtZP8SWJ6+H7XkWyjPLvvKT
lYtFCd94setM9vzsORfz38uFnew51Vs0LnoiKnQLSoH2Eh4ohY9ed9E3Z6PqrIcc
tQXJxzDzgxWQWZCyH8qKmCCDT+TC/YVFuxr9JU26L+KkxHuYiC1wteTuG8UfQXY3
WyOYljxfCaMOLRRbcA/Z+m90TDZYu6m5i8vuwksvcVlbhh016731jiYVhw+/73QZ
cvHO+vSVRuNs3TXcPPoXIK7NX/frx7hv8XTjCiDBl76BHTo9MNHE+p/rt8t3MRL0
piWaFtvqm3eNBDBFNGA87sYSzz2yeefYjfUEhe+3iGdZ3lzPWTBa5QKIv0y1tQY0
Lu9lqSoRTVD6oT2vCGJaiF55VwCPLtgAH4rFYGgP4qEtYGLZsj0bG4/e+H4ijcF4
cHSVnwpHToG7MKuHCnNRotP2kfKKNZ5pc9ctejmsPg2egwNM/CDUKCkIEXesPizV
tNRFT5xiSqz4e+qJ3JDokzkCWVgAu9qPYyeuAkN0LYgZsCCRWgu3UmnUKr1margC
ybkqrNVRdagiuG7d/TDB9NtxZ+LwD+o0Hn5TdeWAtSUpZiY7kTLrXeuqJFkyO39Q
XOloq3eyG8seygv19niu5mPkbgqPNwjDsmfI+dbXRXvWrbPKp2BwWT5er1oKWvFq
FeKNRdc6423rzoxDi4PaxToy5nOUtMtpcYVDe8WYTWSzc8PwJcco1mpEG1Fx0CW3
/0bZvVI4hpVq2tGLIqyrAuwl4+wuwqBI0ySsfOk3JAYZhF8SdcjyKk4L1bq2DpcL
LEWxW6mAlo4QLPrARbkC+Qc3mM3oq9LlfEJ327ftFwhiMRYGclaU33XiXwXabStT
IQYnC9BqEabcXlA7Q6iuGKevzQ6ZXBuWPvaoELfsmby+4rhDR1puUfoGbE1VVOxe
GGxLDdh3StgMhh8kr6XypbTpmbps8Ad3QUIrAqw8/DeWTcuxbtuw4yL0Z3XG2bED
iZK+OmKHcO07ZiZKVcn92S1TtGSO8Pvdywu4gY4eWUbOyn5JspWH6jWyGCeON+Cc
YyZvlSYuvXpbjVPNTr3oTWRdhL5WkOFcprDzMXosqgvmkBn7hkDKzVUW05EzD11p
+26wm3ANTuAKLT254C9PgMCrys993YHU4TNnTC2ZiYU8/WfR4kZ7/P5+sLimtzAm
bdmcbDQbtDgC+HXT64gLpgoXeT9Cx2nS6rY96AGGohXFFgCfd4z2uyHu/HkF1rZU
AvE/XaQuinNAWfQUqLVDaXcKBpWaoBRTjC2Z6OLdWSr5I88OiQacP9Jwm9IyXahO
XfOW89xRcR92qlDHM40X4oJt1PYwSH46Oymz28HA8keMP4GbyB1I1eMob9Pnp3er
/HRGXIB2xpNMQiO1Cmjdb/F2rexJb24kwAYALSwmLqNo8A6kiPZhGE4HtNAu+JM8
dfuJceRlxTL9qfT8TsDqtskBrisok5qBYVngZVc/9BH7Bu9yDzVit0n4OqKQj2PH
7eZsNu9XVjkumsojOd/sbiY7HB1rJVCkj/3JY5dmtPD7ESc5aIL/39F+nlLj10nT
XrHNfSSVwpO5jqovaFMTr3bfRosNumzTozESCA80t4OUN+5U+y3p9p447gfmqkGp
UYtyWkd3CgF5VZDwF57TQ+ivxWOWfJGzW7qKTp8SfmcIUR6awQFHEbTi1PbJOSdv
B5u3LydY4ATvKjKgEi2OoZNU58ASAJ9qcCHBujEcfp6BRb0Xd6WmeP+kz9cW/DLN
OlrLSf9Einjxp17pm0Sd0KGGVyfy6l7ZfYkhxX0SKcVuQ5kVYpdO0Turm5WSlpGO
FIknv39/GxFRR0Kvbwr/R7qS7YYNZtxGg7FGwwTvKP++oITC20COuanBZMYIAjSL
ABAE8Hdf8AffRK1PAhmg+CWcrLGcxN8MLFxHkEzGBwNry9sSyBVpZjZfmLKOmafa
iqJvCrbF1WFyKnEX0g/vVVP6CYovF+jY0aLPVCbMCenXe+1iQ7clGrEze26QkWQA
YM5aHbEVmaAJwAuvfJVqFbaR3+JHnJ4jclJw+0tJGpTqKOzIJ3djn/DWmy3J8+AM
3QkZGvROzbdGtySTovRcv3CcMAFedX57btUeyEff5/742HTsa15NwcH3RP4zwBAW
qw6jErzZh+8idowbJUnOLk05bRN24lCGVNCCkqeCB1khyV4gix/6EBmBvbOUqMbr
Fe6fvjkCUIFQUL3uf2AfFQRs+dAo7VZg16kPZ4KyMpjPcsGOwnrhX3RFK2cbBur7
ytyu7o9ncD1sZ/vDUfl53i1KJbTuz8BjQbl2Rueml5uzL3oOIQasAO+qLaW1YAHV
Q0Yb+o6bU2gXV1QZyB4GN3m2hPVAh0st59lUSsFXelhEnCAkSnCTVEJZr9OpQ5D+
NHoxdtr/NIvX1s+K79yynzaDuecyf96tDW3cWsIfJ/KT7BA228OIIWzclNADYkQa
sOYW/tIl63vtURR7wilnkDT4Xz0GNX2vLRNOxO2bDmBik0Mn+qJPFBocb49+OdNY
VNm/ZU6zTpuRUGsPcwP37qPsF5q/y1OaQCNnPBcKXiXJ7RIQXoEo7shVqnQcs70I
fpm0abeRMmT6ut6ylTDq3WU45pwCRRP/RFyf0dphGaFfqR+h+i4OKQgBO0+/qUp8
9Zh+xc4hrEy9jEQ+Rnubjg7vXs2uQbYUFk7jl4ALrO/2yGu7/bkz6gKs3x2SSRpz
Uoi/VUq9rdirQRptgt5AG51WanGlaX3pgacFKsAykgFfzq4GmeauXUg72EnR6ttu
OlUr5Ptw3rFMUI36vgzWqYFr6yBd+Q2bgFXNFfLeVPW4xlG0t2zUf7Bych+GFcBm
r+NfSFpGhc+65RMAC93vQ9vhZE8g7tegAz1oEobccK6R9kqcrrOJ9TOp8s5dZvCd
s4/cn4NK50hwsYJykNhY3DhLqVLFJKEIsgrv+8HL7Ep8r0HLVWhnYHrkh+i+Lr8v
LtXeZnAJiGa8P7gTSwFGoSKQELX0coWqZBrmOJm25Kl1HXW64+ZkR6Nqk1PgwIwS
vRd41wJLj8hj+JKaldR88neqOuQ66Gqys+UBgmWo4co0et1+Gxty1RmulTSiLx+F
0lkqJv/8ZHBTvqcLrqwYX0rvg50/YOnkP8FoHNEo61UYKUxkyUxt2Gom0Ql3dHhd
yBWDrWoL1HEdDhIggVdfyDZAupeADhXMC18PEEeTp3aNF8/7AuIzdx3mP3K5pSur
NK+Rz8D23a0OE+w6brohyhKa6yodSuW3jfShUSFXzMCkjr0etcwy7QHSpuvyNNae
ARbkmesv/IQSnovCC7hZGxPFhXIPnWMtAzr4Ly/ynotjayKURAXCx9QWD3IuesoB
Ojtpq6VpZMud9r4A8AkefQUENEcDE8Y1M/QBcsvHdZf6NoJLPy2De5Qjym55lODS
UUFFtUlcxRFi83avOWBzgvIOsqULuFRud5D+x9v3JKay/SjsfWiJmdwVsoK/SnUj
zZHoeROaz9Ekf7hlD1/4IEPutQadrUUZlE0JbL1qfFweCFIOJ6RJwNyct/LweNHj
i92MuA1A5Cp+N/CZejGws9HXpiA863rjCaJjjPe1++VcFMj+tTiACSu7LKiNX10M
5h1Md9r73gGBPVNvnBW/Md2Re7SPaXamlvXCwLKcAd0ORrAnnozAhf6K/myLFsqa
kmIqkcNP8HYQtuiWS/Vfxwh+3LqYVwnC7LWCWcRY0SZVAuVaX6c5F70YwFrqz+H+
3tuB+Q5+hH9P4+ne3j1frh/10KZTyILn5jWgKVKyRe6VCLyA91CjgeG6tXlIAoI/
Ju7GxJ98porxkysmgKXqDEWLEQMS3XNOPZWzi8oe4jLCIZB6VHSlyH8bnwQ8xtZJ
SkaUYWMFvoZ2TcLmrt7Uhj+4hrKFi0N0AGYuoC3BkMPgyk/w1luMdN5qmD0uL/WC
z+AutRgzxkC3vYQBqmUG0hhGEGfhUbxznWoRDriXalR32uiymqcg1wewEBkevgK8
jXjJxZ6gnEXQdnha0q3e9OGi0VV663zuu5QuCq7Vo9HbDmENx0gUuLHrC9Mb5xeG
b65GvSd438Cj+cBLwZn31kzk0XnzZJAgs5M3gaD/cMWC6GtcQ6rzel+xVos4CXLZ
Dx+MaG7K/goTTEz6dmkCipG/zW84RM3/Z7QS8NeXwusQPggpNy0kjGgKQm31wUdM
hRAft0542pTsZAlbS0EYnSE4ameSeuOxgUkRi11By9T9lZHJsH3sWxVAPxgUR90a
R9+VAnfP8kYkpQJ1PLteVvX3AN1JU9A36ZpZS2019kbF1t0Cp855W+jRmqk55IAa
zYqISMgI5CXwHyp+A6nFhUTbgooMLTywhfd55XvPwK5VmKuYlbP3ozqbnXXVWOjM
2K6B7bVXRcKE2nXrFeK935d2Dm0dpcuVkVPBD8ULU5esc8zYF52Y1UWWPf1jTu76
4lTEs2aJYo+VcHRwDKB2yTCwORUckjfZERiL0H52rtHhoDvOpG5oTwkqjtI8Rje4
p41WHjkkSw8j1K12Chqy/IyFzyrolGPV8hfQNGtwNgiADUq9qMMVx8+Y1bHe77lz
q6yhFqqZSZGvGDJ+z9yOhMAL/umjVUzuQYUZcodIj2ryIoXHk3LR3IMBC+8FelS0
UciDavMJ0Jeqd/8NVqQUj2B8fjgUosqSoNsNk+eIf/Y9NNDFfltgM3V+9cfEvIeT
o4b8YJcHaDSjbJHlyxqCEJQDZV/WA2lGAy6/Dop+j943jh7ABTi+WhiyX4lM2/6Z
Tv/H6N86y8tXzSHcHPZR3mtOOq/z3IR3w5HrpZbxgsvSTDLLMQmg2SdFySNkvRg3
OGfXK+4koBs9omI+aEj0cdAMlxsGgywOhTcH+NUSof0Z0mk8FW3wSkl4OV0BFLOe
pT0CPF5T7bjoKzofsuN35Qisa7s4VHtcc+6RDHgiJCMVlD1asyN5goIJvRN40vNV
Uc3VNqkHjY2gOmh2FNkFIqJx+/QQOzus0YKAyvtsLS6WQNaBdxaIrQzwIYg1SgH2
+eLDchASTdizh6WcK71cnLsVMa/GBAJTbd8PCTIGKnamUpDiPlWx6x+yI/hal8AX
GDZsdT0JUaojEG/5IKDW9hmGl6QNRRoopVzfOSLbUFxTn6CGOCXWOuoslxWKPoPD
jrcTyAr4AvGkVueZxJTRNkuc1HSBpO0cHfQofDiT41js8x1YMppBzZU7PnVZKBmB
tUAmUswx+TY7Nq4gewr/o249UA5lzgg6HsxGCnDn0pqmAp19xOrK43x//UILBDHC
6MloT1DkX2kqc4kJP6dcrfXlNRSFdDM+1l5L/3sG976U7OxCve0Bd1qfdnjdINwB
WNv8uKQDfcIA9CAQQipKpOXK310oq1f3jXOvARz7FBEFyqWJCi0NZakebk+dTP5n
KkwbZErwmTTVP3P0NJ7RBUq/XbkSUrsY7S1qxV/wvcfJUHB0+brjZjHMnlAnNgxz
uX4zuqbJGqDHd3o/yYk8j52M6ZWBrZipfTIof7GVwkOzekNaeaiOa0mPAOyXUHEx
Wwm4NJwDxFQcepZo3CNOZ/e6KG6ba3NIGwyYZuG1dSid5UO9QqhtajvoHD+ivFk/
+ZVixn45V0KHaQNT/TmIW0K0fSwb1MtEV1xANN+c12lbt0YYFoQV5Gt40lFn4r5w
Z3MlWa52Zy3643Jt3/NA4GbFR2ayhCJgRiL96V/3QIRbroLberp8kC7zJgJNakWR
C3z/iIzFiOMV7XAKHWqkXgFgzlBva377kR5+7skSiwA82Vs+yCzof0w6pN9lSLwp
vk4JxaiuKjhWvV1gp8bMSBN8vYi/oy7koO/ogvGysLpSM9NXtE7ELrpcrGd3p70d
QQhRlu5CW85y1m+skY/6KJibpBhuFnXCGV9P6kHxpJwUic3CYpuF4FDDiIySRpe3
bhALfQUoiQ4yBa6mibOY2+zkQ2uFFb2q/e11vKWufM8pqiDhNErB/+P/3OtrBw7z
z1WtADABYCCFPipzeTBEe0nAAE2R2F135/e3b9/Px8ss5jURR2sqPjHo0OQKesus
UnYrbeTQQdOgS+iujZ38fPukxcaNRel9nVhZZahCERDdH/UmyMPNCfI7M5oYod+r
doqnornINGH/c7Dsacbg1ERAyOfu+6sah7RfCKj1frLA7LdSk5sesivLmu4gBg2U
Hld+yXtW2RfuPxwL/XL1eio8hDv4vaMlWJuszrwBtOLPb79SUL2EewRgD9ts1idW
dAEzcwjneTDFLYpwu8YIAqqiHacXLIC5BY2BTFjX87uoTHniJMpoXJWtw5OFk7Jc
R/8ELl+4lGcIcg2wFOi73GjKJRbH2hEcZ5shrski9YOB2iG4RUZ2FHdAlPKj2yUP
bsj07NfM8bbTL1yA8Fohi0cW/rYQYcXykK6gExSQgwD9shGXUVTAMQBbkR9B/p3r
lFA2qctf67qk2PYq6TVpvfWRcbbIiQEiOuH15iG5pnXaQosSjJJ/0BVi7O8rHhB/
uJCDbpguVKUOqFSl7SEOickb9aQMGwDZ2q8lGC23aunxwGMuhnPqku12wGaASYul
x5G6vqrZLk+sPxs1YSysvhVrvob7ROXR/xZvQ3xvu4Iq2G1a+5T4HFIeeV4ccMpM
7WQG5R3sG0ImStfB2bJJFGRRswww4TA67MfqwriE4e0+/NEu8Srr1M5d/Jaa0e29
cbn478OPdl0LbvFqSzwaykdKriUDlg8FUnUC9tfxBlvIGd6K4s/+GtpuJ5vsY4nO
h6RhG0Tg/dy3fWilF9ql/mUuVJ1NGJ3dVBC86ivB7c4L98YxF14ES5sSgcDriDbP
1VS5OkquwRNuqF2h0mSafcprM5yr4FIgYgAxbe+vzM4/FgyrAu07YTttYmKmz3ka
RVacj8ZrEcNQnJB7Y+Hy+qoaMzqHjQgQu2gah/vk8+HEd2jmlM9qmZbMAvPEc+Oj
RZ6RM/Cjql/a6YWchenhsx4w+Pu5gsbnkKWeCv/YVle6kfhB9f+A1kZNFpIVcoQ3
JRkgGY9+kTkbqnCFkSxJsrPcXLJHVEUKTZl91tMJpMM0u9cv3ldWi0NkurCJs/Mf
u8SwTmP577B0bgs1QCHbLBSD0aI35VFrBBhgxKRM3W5clQh7T5nlU0lF/Q/uFTYF
0bN4dt0MU0HMVDWtZ3+uxhZbNmLtkSj4BYS4g3QelwsiFVYiSFeXM6K4CM4KAvzd
z8c/5BSqcbhBxRjN4H+mnvvvCW5KEQdKWLWLms8HAYjuPIwvCb5oYv2PIuw4BeDZ
LMnztO9Bk/xQTy90tnHZsWW0mwy03x88K+1xuyF92MZy+0228yvLe0Cb7iVKHeUZ
hLsEqz6LRCQECh5IxUwbMriRJIXLT7PWyIvl4kdzeSAWYXdiKJiVrt9m+60Wzqxp
hxMZ7k0SDRltUSu5HBTaDCt0063zhfoaygwcLncNYtr3rtniiVOLJk8o53gnzaiT
AyS9Eb0n1IJjWsyvCmgiyPIztA9uJIBaX6cPIDY9lucBPzSyE0IllF+PoirXIgc8
nb9snZE+7CCPRuJ4agtXAPY75RPKquWKCciOJutbH2ZjkK1LzblthU8zwLAuL4tB
0elfvwKCoESOZps6r/fpYSeNcpb8xzNxtnS/j4zw/LHd7iens+WKTaygz8S7Snz/
9arY+WS1PYifw89LjdkR8XCAcVgSS0KOY8zdTW+Izel5MorAJXc5kLlQPQ7KkV00
pdSMrZbr2foFWTJUsBi3eYdHZPMXHlsDxODxeV7zPtI2OYpPAnJWobxKjvlP9dZR
nVBehd8grrmxv7jOY2RzLE5mza7W6fpxg+0xbXgdAYMmfnZyP26qMBZBnp/Nb0R2
8dv5GJ/PY0Awzr9/hZX+4d5sHupCw2Pf/ktELVs0/NK5DMUOwIlQOym6LRG+cH/2
kTK7vUnyJvYo3jNuh+lDSQGy5la3o+qFQWwoRBtn/U2eHu/8CJxZJ/4GO56EHe/6
dkEK9Ify7mmf1n799HRhTBll18XRUlDJZj6zgZxmFXhQDme60heqMzkIBQ9d+DPU
oTIroupzmiNjv7OgRdILiD+kwv0JKz3SFnPCYHp7P0Drjmna+iJQz8O0w7wkL0WY
HTczBmW2/Xmmi271Y97omlAHd+Z46UZUepcEtqpDDz6LFUM+ysImNKDp83lxdqT2
hYkVVXFjqWbQuhb2jYT0GDZzamNbX1UdywBc5KFsctq+V1ydaPTWheHPCFh71wYh
0XOLzKuWuQO3uq0Ip0iYhEe9iRtt8avo4F7goSi+rkmXun2LdRrk1P0CzMGZw01v
PDtSyqUiPJdQam25CU0DiNsURuXE/2DaScv4ali+I3mi8CUIWpTMWvcSPxTmP7CC
8H3CCXRxU+y7IpB0zRL5xMjsm5CSrq3B10JIF+58EPa2T4UfdrZMVUiyQZM1ffxR
pREAsEkRzFCwLLVw8q4CI2rJ6f0Enat6rgZyxLFByorzW3DTxCJipHqyL7z4Iqly
CuU7lQE86keUIISlzufVwDisjvLMGD8oCJhRGQOixkroSFzcTgY9u9KHlXT8D7r9
2gsDmb3kYF0E3/FqnSh1h6eEzKX86DUNQKZ13mpXXBcNnJ7q44+ofwkbSHSFlSXH
cGEBFs0BFvP4B/vIKgGa809XMNvXgaP0d4ggZXxmg7ti6m6I3cSwIimCJXis4IOs
gdhuw3Az2WFIQj5VKrwznY/ym+Aw7w+HSIrz2Mvgs6YSQJvwpTwZsRgtbiskRDu+
UCqgpdn88Ehe01HuofGAASnVolTzzbFu4a3DQhcw8EWIgz9gpzrm0D07NTmLHdcN
Lj/JWTrRnZee79unEs9SWv3d0VPjeK7VJfK1AcplZGZP0blIHalVnNLOjGe3qrE5
n/BWS1VkZQn9u4F4GRkqWXRQMjPiG2YKbaMPMZFVri66TNjkNHQmSKBqledAksB2
hZU/RVKxoBdEmzFFiphol/rod3gD8iVuTzbMe10iBur3KLd478sjvkT3GMvqAWsW
khZ5yI36/jK5XM3Y3Sj47crebSIEMHPxcr7TBXBqfYa9HQyWbTczKObx7GAmg88B
x4L6/29jVU4oGsqDCPZayv/EJMwHInc8zeOJ2UQcWKwgRD66Yd7qp2gxLXtU23Vk
mswCs2gad3G+PAZ02qP+dka4Qo3bq/uKCv441mjIKQLRstxUZNUi/xl4OMNUzdAq
zeu6XROvheeQi2D9GvWmktP8N/QEORxOACJzoa9W5boC7XD83feHsqm6T5CYqJ7x
cFag0NdVxYq+BUC9x5E6xuQlEOBGIFtBghQzPhyIA3jVhIBTbG6vJ52/F6e9Q9N4
w76sdnZjYUn/UMBmbYea85G4yk9jUIiJH/FaBAGZLxowCf96K+dUGw/mQvW3JyfF
Oe6I/bdVhwx/jpu6ZpQVKqlFzG4e8/t+y4WK2gikoKEXOxRzkI9KU0oHC71CY1W+
ciiFRCZ1L9C4etooINP9NhKRlToWFt5dDGB3o+wiMUHSvSjfi2G1wJendWAAPoD0
APlb6AmjCjagZ+aZwrA4lMGhF0GLjcVgO9xsM9Ge1SPCXaI2UVp/rwf1QyXk8dNQ
KGAp/5I0rbrgRnyve3X6+h96FV2nSWgzMKYkQ88LDvS7lsXbIboG0MRmJUbCs5MP
o/8wyQ//8Lj0/bd3SxLy4Isx4wsWhUm5SD9RrHfK2sUpvhoPeCidmOsNMMYnAZLQ
OFAEChegWT9g5Nah688l6XCPiEivDrvyUOdBO4AYrmtVqhTUgo4K18ohBzbfKkv6
v81ZGJAC1gL+yEOsVnJsVQLYQeXL7Zzf+ziPlEkQDUhnxdL0BEBgrq12b5DfrlZB
R/yAM/iH1HVWpqyRM2Hs4YSbVoC4n9O+MGUj7oblUZzlTKN7VUvz0swUNzYSWN55
G0RDFt4bfLUddJYDNUuoj4uyD+iNcMnmMNVWE2fQ7pXUyRk3+gGWcJSAE6HYMKnS
ZlLHW76fehMrZ3F4hJuC7qHDCUt2ryAl7IEYyjRrvcIWmyEAzS4aB043aw9QB0WV
wgu8Z0kVz9473w9wBb7uXv2okkbiKsFsLoBGynqwpp+N2TDXh1D4SMzwZbt5gZki
2mjQfnzvqgNUnau1fyqI2T2i6yhBQfJtP3RPut/A8YBQJUXhXPqE4xXltSH7te4W
PFQUAsJ7+02VGcSi15OxRYHdtTfYKphiweGijX8hNr/7+8Tm6Dy5agEhMXzDkPbo
aU2cTJpZcVCHGoX7g8RqhRvbyLiMFl8Dg/A2LLX+RpsAHZ41JvRPdq9u+S7OuKfp
riRMKQA27ST+2qC+zx92f/dNr/6TUzF15OHLnY4Av/kbVWEs0R++bAOWFVlO19AU
Mv9C8vDxk6ZS2DkCWwHw37gKuQi+6oHNhN9UvfGqKF4/WePP8W4NQj9CWBOXWy6B
Ufjt6LGBMEucNcdDyPgrvRCy62mRr46npY2IHKssFdpCWhZDva2HvQAGsbB7CxHm
RPC96ExDwThXMUaEmXF1KZ25GlmXZSuzep2UYSpmgBmQz8uxjHb7TF/nudDOFJ84
qKu929r396QLyvjU9oHBJgS/MXGPnKSbvqR9jm6qLzfzvTbJAeCbuDOUt39q25o4
Bad/UcawMM8KhYbIXkdW2MLNA6H3hndFQt5j/fmjYjkyNOjEPy/pZN3iE6JsWFFu
xkvcgqESe9SHrGoOX6GKVSsfa5WsIlha7z5z3pnzdKU627QTmTsYxTMr0DWp0cVU
3YkXGfpvzZxLASb/bPxDMCdSP+CRlX2R/7aSUuuc5/+tO8b7qIapVJIrPUh/9vF1
glh6RnHqVG3ZUdrnTfLWnYx0EvLW6hFIZ2ljQ7Hbz1C1VcZZtQmQgyISYV7NCGy7
9PLvbJ5Hu2XSSZRE1y8Z/wwwl7D9DVxSJ5vaE/Ro/ojltoLSLiiqjjs6IvFlmMTH
SiaAtQTXNBjkjMj9SxMjV5E7E42LhmqeTQ9xobGQjc2HzKqGabDhEZJRoPnfk3zZ
UAHVBa6S6uu8CkPPJIPMT2+StMGMoEqWKIDgmcgcUChHRmbmkmeZNJ6+AEq0sISs
Waqsk6MEJ8kwWkwuPe/vrmA7bTy9JzrcTDLwZ6zCvJRruaYMhhdHF+YgNd9ciRFf
uREWkGw24UvOcZsyjUtXpMhknyTg6W4UXTQ1lqvaFv3M+4K6+H1KxHfe3jp+AFgw
Gnu7h6KL/tPomTKmrM5jFI9ge5kEpV0V0L6DyRjgK3UHoGlUniHwbN70Q3NaYXEL
1I4uQg75LoNLdxIjn40OXnQTUixFF0D5KcleG45mvPLOai9Y4PgChSkGMF0HbktB
nIuwnKQnwpPt5qI+CfQpYE5YwSpt+ltVf76T+Oqs8rTSP2s0oyz+dN8P52xi9Rgo
NvK7EvAhYGn6TdzBEXh6uSLxhfu7B/oo874PXPdmRwpGXE4FKf2URwQFNf4dE/Zp
SpTK1Xl4sfrXQvtJG1jat0N5+AV/Sud/NuE05HspAAz7KwPlcjIhtc8sEDg+lvRK
0YdXPow405VbYWnpfARM8laEQHV6ucyyKqnMu5G0n9p+CuTYUDRvN9gZiooMFpL6
Td7jf2oFwoEQd5MTChQLeLXijZ6cQrEMEP3fDbkmfxRnmPB539m2nlH7gd1Fab5T
rky6gQ3ktnl0GXMH+Pjmp9pki7G9tQM96EUFnZqQiNa4+X8RkhVXkCImpKfetq04
W7lqLfQPOxNSxxeUr+70HtBrA6pDAa7wCGTAOJWOnLCKCm2q03HrBZ50VxpFYgAT
rv90xeEgTftMhXbeL7wUTKHYf2Ylo7alHoiNgqITNKt0LB6k92sDZx6YGwQZeXrs
ZqB11WKB95xYOsEvW8oKbbBjj4CQM7Ejd/fJg3a9Y5ixs/QDA+faU2VA4gtbpPbV
rS7GuxHdyIRrwTdpVW6IOJmbIA0YO9ZX4JvOVABFdNVzptH6O0Ww3NnMkagJWIZd
gjmhyxj1PzU9JbVpVFocU8Z23MCrh5vsKA+RwSaae8smQ330FRLQBiSBvzxIWTk6
NS1eDZ1fiW9QWo+vshkrUoFanO+klQzNtiLBsU5vasP73vjhntT+u/ec0WUsX8DS
12HSIB5ZeYKEI81QfiqOYMfnQwUHRPlBaHt4QX3HWT1S8UihfLRxluxoSahH2RRV
C104l+xP4QR6B0HNA44ByDT5Vi7ixHFg88GYNm7l9zO1v3eUc9s2w2QN0o0E9/bY
hWfAqiNhUVUjjQfFSRL/g0pUpU0p42DZgaOsvAIaeFDafENayn03jtsbEtm7Mn2s
ZC2b4DIaruXqd3tNRXDQXQg8O3v0CCaiefckDwwCCH/XM0V3wS9gNrbZ77yJwdVR
Ho1Lk9AO8/OHftquJ3qQdrSBNhwh7t9rVe+R5JZ6X+xdVWxJzyQm/2BrBP72o/rr
JxUoo5yUKWmpP0hw29/WA72C+GQR/xsTlg4Dkm5Ap1/ENUT+uoMuHusscrT512ij
k1L5PG156wUy6ILtLPl11WMytSOztEfgHeU6mEN3xXR62EtDaWrotyh1DbCRh8Qc
YK69rv9caj5fkDu3/cSNVPE7Vgru/BmbdeAoZLD1Shxku23mDD8pTHGX9wO7PXNK
M9MhSRN3b+DU7BRhTG70pvcAi4T6rdmIxgQ2gjKZ2NJ2OmG2Mo2SWJOTO1LO9NUa
vGrDhFQbxH98dD8UWTzn/Ajah8vNzRstNV+s6hpDIqBmaRRjQalSWmmU2QsiemMm
v9fJ8yGgsxY0xIEfa80cwio4RS162wnSXeHw3mRhxWMjZil398PoG7t2Pry300L8
skz0fM3YcV8ZgFxjSxnk9Em88V0IxPhbcC8WrtWdm9xhpCF+1xmkxVMGqOvWl8iw
/Vq/KSdQCuYHCAd9pLYKGxywvtYfSWxtilbqkO+u461WTYOzdO6oPzeeUI5h6nCW
F3c4qt6Tn2/O+bsNMeXzc47l5wgiooVvBbxNnqsVuTF8L87hh7KoNRHJEI/fKzhA
erhTOMGK0L7pGF5bkAint4716tqKq44kg9jZ2ZKKIiBT25yUv788vS9ed99TmOHX
QZRi20/B227wIe8XoKQpl0sngN8KIvJ03ZHbdnWqYWvy6zGg/hfl3z5Taiu8ntOr
uLS3hy7OFgbsF5RRlhsKUQ5SMjDlPEUjXzn0wvm0xa4vSH6c2alCS1ZMn0b31zYb
hMbhBpDhL0lYLhIXBqyuh9XAAR+6rNFOdc/dndkunBh+S/7Jlbbdh42Ue5gYrYq7
VlPRpdU3DuHMt8Ttn/nq1GpP1OJ/bZo0cm9hVU4afiVF0EFt9R2omleMO8WK49rR
UmiuYVrMlayIMExkwWHsVhWVcRXM4oD7czPY6bsKp9k2y6MflGSrrVaqao0sRJ5l
bsihIldQw37ffOmw6dyrf8NVTs2AKjZJoM/0inQgRhCJRznwtk7u+3tmkErE4n17
2j8PqhrgfFCWO0fQTWuZvGw9Stj4iukd9zEAGPbxUkuRf2gaSew480fHbDrdpR4k
B3E5TOesivK3iewMnABQzWbES61CJyWcDkOi9O2rz66sgVHrXyjQwh4B8tCIP9BF
W4Z7fyh+e1mQ3zTTnHkajNKqTX4Tz1CmmY7AO0qDgX/TpTBuxdpRuZilDfEI0YwO
XA2eJ1sS0fijYHUeqiPAkvOr0lyQfxwSYZA6XxPqvvSp4/vvZbm5yWPfm/P2D0fi
HPx2Ptr880L8QM2U2UCQX2aKD/uarUcsAWD86jlCVOc2pI8vTU+Fh1DKV404O+Kc
FvBw4BUjpR+VUVQXMpcFGWCD2EKwZ7jFiLjTeMwbCXNw9Gg9abM+ntS8PUEg4qiq
szCzYyHnO3MRrwF+Fb4rNWfEL1Wclen/bqcyWxZ+rEG2q5wEEtqQxA0qkDii0J24
nanlJoiT35e7ekdkWIJ/BA0zJ0y1gXeteQbkKoq4+Jq33KYjeCxuaizro5QDMJTE
mXopkvnzW9VIS8+doO9HTQLnPNqM8EGTUZX1q2UHK+BtPE2cLTfSJBpapdesEHlv
8C2A3WZv/FsAxdAjkXgd8Qs2cHy555zZnQqHi0dShLBPcYZuw3pekPB7BHeo/9Mk
pqrm/UBIKZxahQ4h7kHWD7M7CqJmcxeKqakMx2xHyzRz36+CIhJE+7dXRNTO+EwL
Yy9bbMyYls1ylxdcY589Ez7zs2+PjHf+np/o2/OvCQSWScWCpfVyoaYCtnC7Yvdz
/zWzbxf4xQ00ou7SN8G7mwfSUG2MEiM+ROQDmjDhxyi0zKrBWna7bVBs6doSiunU
g6dXhYDV2req/ypnvCT86NesqVw3Vmy5gAWmibgmFZdRH3zNE4k2QdCX4T49J9tF
OwDABBwxYLN1uRJQxJe1p3WuKn18kMP5WFpzcArSnxmuvgAbtXWWbJ19Ij+SK5XJ
+PsccWb6biDTM51R7Jlt7BDOdlylbCmXYG/IJHyrF3fO2ManC2BryIf/uUlvjqAR
rATvZJaxJtM8rLnAViDJwI4Pdq1bRaQBGyOHrNGD/xSct4k19PUH8VaZgQ/TMUaF
NQMNU3by1/pjIb7rwFYQlQkiZwPHfV4J/Wo3RgM74WSpTR0lHB/Tu/s+lh0mnMcB
tlXaelD2qXWIYSpBVUbZOGoU6bNRhqk/K7lDOcpC3t24wbSeaJ08B64TkvhADTzz
gc7HDyTLh4AzT0boY2h7RGtl735cLXguQ9i00zTm6t95Iy/CtJJKd8lRmAvp9jbH
C6CpAWTYuTYyALePpSp7mXIM/sXf2a74LoUHGutPqxM4fKiDiT52X4K0kKx7CPCe
qtCmsX/cbmW1SNSD29+w9Oqw6OM7Vxt3nZ3U5Jp06cB/LfT2ryeZOCo4eTe0lply
CVKkwKm5D74FMCc6M6cksTGv3GfzxCaAhVDI/sx93r7oc40DFxAXJhMGhfs0Ajte
cd3uw6ceKCK1tXOgUpq0Kjdsh/nAdUWFerI5EmVPbOWl0XLG0P7UYeNxwQL7qhdQ
nMPUAiRNWXbXZuBf79tFWlFlJ7V/xHfmesIvQiWm6uomOo40U8UhkTpodVbc1Vp0
X2d9/D871qwxzMuhIKSAZ6eJ1UQXh8WFArSJ6qq/cEQvn8mKr85PR60bvyjquOXL
052x2uO6X5E27Xmb0remQxVOB8HmbnC0DCXGVxbCMP6uS9RFf0Z4alqpFInv4Fu6
4sbYACF5Cx3nFZGfrGBovCQzpk4mWASWcZUkSvMstOoz5+RHWNpTbAVsoNf8PU8A
hssqOUIp1kAnZ1VRRDWRJNM1UkS78hGNdRhnF8MNvsItsdqykUCqOTvl/cKICAwV
5Vkj112C4UHlMXxX+mJAXE9zsgsEaVQXQNwJVvI4108+IkgZZTd5ijmX4KrPU+e6
LjBNLCg0wFda73Xzom/gXIb1sV8IIFbn3PF1H7fPIBpHx9dTdXO6iEGLH2jTIkjv
PUjaNZQdVyJ8xKBCSDYwr+WwdqtgKJG2s7glq86ePkhGeLhteYuHOdxDbksl6/nl
NKbR2bfKeUfwGLEI5GTcU2u7MZnW4+W8PP6WWg7BuhI8szHirXzHpE3/oEwBoiEr
MLITO3KWfDiX0f989s0LquZhwUimXNk8hhUR6MyuyWZUNfkUut1JZzonnoLwrA9n
Fy/Wcp/QFMYimUDNWiRPWuiSJ/4hKOi3L5bL2bK/kk366mNQnp/mpBRzqgHUbKZQ
4dNhEt8KmbZaOz6qSipSujYQqcli6kd3uh+QhUo53QNK0Yc82CoqybhmoglDkQzl
D05T6B3gOxcAYu9Gc9JmIsvTDutuNt6hvRk4uKq3zc3AZedNx5EDQ6Zgi6t8qhZ6
mfD34NHQrrWrz3gEacSQ18Lg+mel4JHfr9gKJHTCUiCsun4nfOCUjwyrFRKm2qVe
VR9P1eMqVDmxGhpWwnyyP2MTav8Agw3mxAnAtmXCzYrNB3L4SwMnWPFA5/YRjEm7
uEoqGV50XvY6L0ljWMvFKtACB1MIWS1k6woS6AvP0nfcTlDiHpQD5icFnjblA0xD
UBycQoh26lB9GY0qZzcLEr+jO42ZSHAlK8g47JkrDIlAJyHLz6Qa5gpu8ORZkKP6
QRuE6QAp4lQ/W36teSV5lgduwkS6x+4a0uMuqVLfv//bejbVoLqEq8uU1QdENLE0
6v8P8FPZ6lxOoFMJ5/JfEDCfG4y39Ht0T29lfKyNXH6/qmxqM+71bla2HmYjxLMu
7OHwa+dLoAQ6YgqGw0YF0aC/CsXevrmp/HLrZ0QvGT8RFwrTn2s5xnwZDO9MkMhT
SQdXVdpGvEotBgts0fdkeDfFUWTtC8tRyu4dHIbUOI2enBVmqMbEbAH9I1WaS0ST
c5pXJq70Lm/VDxKGNLYj5ftkGHTUdhadWBRfDNyHxTveotJljMahuhkLTEyw6SRu
IvbPItuJulNFTlLFiEaHeK78IO8sC77oSJZwLwya5Mf9V8Ec/sSqIZPLpXk1NYcf
lxL8B4ZCQfjEI7+IbctPDzLhoW7zeWAHi/Rh5/RcXoJGaZSjAr715U7dd8x/2q7g
wkublSAI+CXsBdkLpj4qOtLKSYi92HjpfRin1QWCHE1VwnkHvm2MFBCC/OlMyxgg
j51fErPs7CJaLSGkoy2LRTIni2Q6HEDXBmMxGObrXKBu2VceZCtPiwT2EX3HDtxP
4KNsAIfipSx8meE1XAcz3wtW4wdi9goItE2mpzwHWPKnkzIre9OMSJ1hNToS5Y6d
hEzKbnQmKQZvaJwW0yR5gec75JyTnIfOCMGNVQvUlqZZEpAIE1MlNhgNPSS/Ol+c
OtEWQyPuj873LhuYt/PKLmKw3TmjrTwgkiPJ3svWpH0JMkWwxYlF8pYHYftmjSmU
a+ibgNJkf21U/tn1h+k7y9HhxQv72E2Gj14yUtE+04FVkNRJjoNNNklN1HpTUBg0
30wNxWz1VwHqAV2hPaBGwoK4Wq3fJr5bRfRhoQDmTrg6P5o3KW64HzHE+SZONwHL
guEyYQ9rosJEed9tFxeqG2U8ydxMo1T5J3c2VNAYDGL3zFzQYL41q/D026wwep0R
O2XixdgcnFRicZ7TsxtIXsYk0nvJO5YMRytzwJ58GK47lVCuiKk/2q84F13nkeNS
9zR3gbThXRzdAiQqwSGSyU0iaMXgl6XQxBtkHlbabwepmL7nXcL4w7o3zh+5u5kK
HxaF5ktXhkGmy3IBHAKxv5sgNoX8XnKzVWxOLZCiGzdhD9h9scPHffieig0wLoVS
xxznagTZAQYsfNX9l9YIfTkXsyomuYvD6b3UIllfwVZPJxZqKYDREAfnmbZ4+Ew0
HYxnfxsGcdad6zpa0oGZGeie0XFKnlWg+Inr2UqZKf0hbSAEKqrF8sleF30U8Kro
wZQIah66As+1rXp1muL0wu4p6z7ZQhDoMTSo0hlheVBCK+0OW1dFfNplXrYY4Oxd
09xG1MQ8cZdcuO/IZdtZXNildAdeEnnTqTPAx/WJEorLaKOoqFqe+7TEESS5pyXW
aVtzy4uf/c7d28MHF6c8n0Lj4mY8iG8oJeU9/XUTg22774tWNqOA/Ga2TU11R6IY
ndArvVYOJZty+YnGGK19AKJQMgP+OpSVwod+KcV9qXXwCN2nB6lyoTl8tYMy6T+g
X6ORcfwJkU1SORWPzk1SXO5MfyBSLgEYZlEUhLp5gwi+6nz2PTMLje/FalpONeGu
gmQOEWdY3NhA70TpnO13ldNRI1Ie/b07SY6hELABA6U6hTiJb1Ze8ceQUx7i+yrH
b+MhNK23sTRaUdDBydapbF/Moflj+N3rXxERomw2cGkvfKoA9jm36mAx4NgTWiVC
33gZEGjDhHVizKtjWB4VHDkquUp4Yz/meLLwTMl7E8y6n2fnFwCxXK79+LY6nKKQ
VI85twuIKXFKiLUfT3zOdw+zPdvZI3yEIFDdFAC8QneXi50ckQV2hFX1LjhTYVgO
8KmA6s3dq9yTsbpWXH0DEW4K+OAHwngKL+Gjkz/uPN9TcEmlkcX+hn8hLoZedSbj
Ma1evafUsJ05xPV00fkhPul5Flo9mxbKb8wfFiouIv2FRDDVQoBtThTyavD9CgR0
u+7COfK+dGRZrW5cOvIQSUrdgEntufeQu1+SZOInEK0FPVTbchdb0RkAtjC4c4nE
8NDnO2mDLOdW9Nv0Rv3A+g4mDPwd7loL6k3QM1xOiDE38cp4OlzD1UIgap2EqT1u
3gfn8aioDGnyyx1OfW5CWLT9cX6zKABrglrWe1v0tpGTZ38jGf7V1Xl/qYxLhVUW
hKT/muv6qzqWlQqywhJwLY+QrXzIRaZXnFY57fcEVsskQ5j25VvbxkTNL9M/BAA5
6LMiXwgkINh+7604OcWZIso752R8zF3woQM8WafkBe6CpszxBX83w/7fMasJlNjz
tBBM03Sjlm0QIv0cYkkPtk1FVgDTfweTk7k/KIxWBnip2/nrbY8uKJCnEa0p6Rca
GrlD0dx1bvvM3bgNbYRHofDVQQpAGWAVVMR0tXKfWIwnOm2frp/pLDLp9TqbchZ4
2oodrwFeCrQYrd5PxEDxm4vYTYWypOXLGgRugJ3Nhb/O0/1tpmf/RRcCtEwR3Ni/
kKmj8NExBDQ4skdRWyky1LB1nMdiFOS79zaC8a31/fJM8HRYhY2V7ioF4mH0rMiM
BvRjbNryH0phSSKcAgA2NwOzIGr35uitGVuxJ/EQRRL/wRxYWWcPYGT9WjL2mH4F
4aQpeGWio6QTIhHjAe1ZaQ1k5dOuFGPTa4SMSlJE4MmEFHJpKAzUeO6h7D/m7YC9
Wbf0LnKH8y5GCh5yISzR7Nd5yNYWZRaczsh6+FqcPsWmiE8HLHenZ3/K0E/HIvKn
2GjraPwfR4KNdNBZyNMCXBo5zW3D+4XJ8s+B5QRpJyrbN1J00xiXa8M3ZaTjx/hm
+Xl7iQCcB/BA56ySeEsk3weT37AscKjeu5g8GkNgkuFplNgU/38PYvd7dBWbWY+V
vLwmoKYo8Y9DmprZeQcGHSbgBaXBJh/tkS2jykPAV3W24kxMAm13mz811ANd+XQt
7+6Wkn9ghoVPTFnLtiOqfBpMLk/t0jOTWV2heqw/qHCfc5Bx8YrcT7hOtBAvDlBX
mEryRXRUI0qsw0XZ1EPxMItyhqJ4gOVYgm+pGe1uas/fp8g53eL7B1scDMvJJyGH
J76LhxeXN+Cvchu3oGvaUPcudrGnzN6WytQvPRTCO/RFYN9bFudB54NXlNG5I4ZQ
njwrf3iexxWDYc6SIoA5PpblDQ4zXy2548RE+X3xWqXjai9Ev/zQtT9NzD8+keJ9
k7760SIFt6LIAJorUSoCG+MJ3er76gX4mtxwwBCjjp1Pq5bGbBHsvVidkjtwJgTU
NNWO0e9bJwi6M0NoXF7ec/RJvaEjyPL3rOyk1XSTkliMAQh+KtXxKYbK4/md5pSh
WAUarL9KSCbDVWaJV4gNMn96c6L3h3K+bTZXaEK8UaiYCVlYZAL1sOyxmmQXkUWR
3Jx8SuNuE4Y7bZxkKL0aK+Q1n5XMksraTih+ZH30VPwTBVjxXr7r3H+IeCwvghx7
iQGRpC9fYdUbwF/GSJkhiFfBlasti1IBxmkEV+F7atGXC3MLArgn7pwQA3hXgyNb
Ykr52krAIpp021Ox+VkYzPeaNpjRl4Sd2sndM2xkYW4KfZKIwejwkfYcnt/jhdw+
e3X/h2pvqA22OqNNbGXAuptKmiMqHjLyyGaEqhO6y3mXt0BQR+iB0+jDw5AWmM4W
U68i2XNSfsBF/id5v6W4toBooqYizsNoKXpGfjNi+uTztIxkj3hTgE2NpzQWJFgU
Bl3NFv4oZWiQ0wdTs3syi3haxNIxO9ghKUsrqSv/88YaKmFg/C+sRNnpMabdaiF5
qtsq1dWwUJmcDCx+QeEBAACeD0B6l0f5DCrmljD/nIUxheKwifautHn19D0u5dMP
HI+JvejgB3l6do9q7eAr58/0xFHaOGbkq8zSDtULqhq1OmQC0jp/+TbeS61XOkML
+EXcNLdOvN7pPBT73i9xlci6IDAMZs8A8jayJKY0mQtcq5JbF9N0yLy0ie4BfgRS
goEIDkDdwpITxRRZlg7W9VGNj24m3UVtso0VNvI9RGLGQ4pZW/2iW8BH0jWT6R9V
ELoMLfIqkasJXwVOKxcDvkZTz1afFk3fA3OKQJuOxE7YpTTno7CVkhQTot6mKnhj
LBPN6kQoG19uaDwCekrG7ZGGIsKJuhd4OufV02LH0ZJZUIlJSdZfloS0S7YaixxJ
Y/rToMwqDs6AicfBH1ai2xUDgCEVMzgU7150OwO0365/wHQEZdW6ChkGBvjnzMER
Vh2x6asFoUajRWJwi/5j+Dq3IlpzFGCyZVrbYDUlXdpYSduR1aEmnRUjiBZ4y+Xq
tpPNU5555WABMH9y9CplvrXN/eRg9YC5XRvsPYFZJMQPn1uhONkW8PuzKIaOUfoX
q2rrqlPqvHnVjHtF6jxxvupHIaUWp1aKLl9MprR1KYnWuEKgJ+p6ZQu8a/1pNEqN
gJH3DA6gNUe/LTGXx3HVE4auRQE1tHJhSjR170L24FXzQ29JwN5fTEUsXIcQDj19
uY2EUnu+o31WYcD/aUi5vEPD9q6/5RESglaNNyYO2DotyzEQOBh9P1FV+HtA5Puc
EpVMxgoMtIiS5rIrwLIQZMlt9BMZluiDMeA1hUqoTopj/RxAroIclAKM96T176YH
LtwAT7+X5Ewouwqkb+5X/Xf6FmH7IdP0NVC1KZC6UdoTaVDa1ymcK+zkYD2M+Y4z
xcgDBqdNSdawMNFbg5G0rWUUQwxEGqqJm4f5TZ0wn1di7b5mv0zmataeknXH5u/I
OlGzGMcgPm9nJLkx2vYEwbo25ftrJa6Qy8M8hi2qNzfbFMeJhRle2Sfgv4I49Csu
xlsAmCw2Idx10mg8ruUrBhzS+vZqhgUhN6ki2HhX0w9//cQJNCmf5LKi2FTJqSye
MyUmtNaGwpsy2epYw0IcN7eoYl6Q/MmbpgFGQ2QEgAztMrNU1oro5KP9CCB6V7T7
mpB7B0LqAQNmBFfTsxn6RqCI4rMhAaSxkyf73kVF6j27zsGeBfAYeBgYIXfYikYS
Eaje+x6LfvExPVB2osCJBv0AMRzyD0WvXH1xh9XNi5tuD66UfAvdmZrlOKxGWWw2
w5cULvsC5ZJz5eRU0g0gBSPTqqC4KJ9ZpNKNueLFP5J44nNxM73RN3d7Uy/iYT7b
Tn8dLgMxXQC0tIy0ox4lIb8bmc89mZTdM7T+l0RKz5+1HCEdcO088Au7FhKtaq9j
OResMs4o/No5m9fSktjJlRFBbZLnxKPHOOBd1BlaeyqvFR/u57ms6SasCaVyOIGW
yFks17TMuIYosz9sTuCQf2F1ZPADe6a0iw3wjNgzPSTBvKuRVCPe2RsB6jUSceqa
geaerHtXpwo1KcIgthyD8IGTbzAPOASu4OsUGuvl2/j3heNLN3vPeOC+AWsmfQUz
pMWof8Ktb35eiJ2eW0d+JT1v6ezpUhRW8FHitVm5fd7wZ4UkfEyDkxXRZAyn63l7
L05sVbqmO6K4Z+408/5zRb8QXVjeK59FcMnG5PThZjIvp3iThnz4PipIkqdrynNu
EPMUZH0w0BmN0f+yLU5tn+2+G1Cv2biL2mcJbS7EcSAvYXYxm8/0jheNZADzmr9E
ozSwxmsXQ9RpTPlcaLtefaUAk7qbaLJuums0CjJ54QkFvrgFtySuK7I8mk68Cbou
QwCB9MVxXpwEAbBEuL9Xfk0xCQUYIzl0/pNcQSgtsPSEwC+g+q7o7txhzT50O59S
yJOefO6RCmMLcmA/IRdEUg3ztERTubArYNkaJ/zYleXZ3/9YzZPgnqvHO8MqEWji
CPNElShWrqYruGPXB/osWZ+Wwve86Tp+jvxAQSf4ayWACsP1i9I3rOewJpR5j/n8
iCwZ8sd5bTZxZ5osGcqrvzXdInceHaoFIyoKMtBlrLUEIdSwFn/ptK+M0svxdnZx
17BiYkf9jn8Zu0av+Cp2G/Leb3He43p1BI2IHj1AGJIZvpPg3ywte2D/TSGrlJfP
1+VpQm9/l55Sex9QZjtnzXVuvAn/wilPgSnpZkbCDaf/C7GqV5ycUwvRCaZMmclm
ptNekHNjulBL3q4Ajq1WnCHrPDtcqvtBCLsasddC7g5sgkkm699ZvbyhY5vqOpdL
gHi/zlZH5p96lobCUyALFvCLgeDle3EcoIWqkKkZIb69+jV6huL1N9uShE1dQK4Z
WVNj5/BXjr+aCiVVCTul+rw6Iq4pObav93kTkxriryOMBeJArDzkI4eTYSfyyxCG
aYq7sjBPtkDdrNqyE3yQ2wbBU9tlgzV+s+KvefB696gASH+6aQ5DWeSup0EXzvJj
GPIFEZinmiuzN2xRabP+TZsDxZDEzT1tkgmFktivQVL7xZbDN390EGVMsyXU+Ovk
KeBfTSBipGdZKusMA2/pE6KQGTREKWTqIQuY4s5N/8rU/di5yYZ+xrf9kaPYNyLJ
XpY61fz716XQVW1jnTnO1pg5zQNJHs424yqyNAeGuVd91Uq0cjmZiILh/5N0K7CJ
6Z5BgZEVAKM9vWb5HWreVZHFCpWUP+MIVXxmDF6bFCtN7t2kpmoVNL4kRIkouHg3
p/HDNNyhJKCgTnz9ivyNPQL6IadzFCHKuD6gpVLnm1xFP4SAMylNZ5d6UD+pDlqg
JMWvOOwvbZRLamhWhRpTyx1d36C2nImZq86jteu8TVOuG1Ia1dYDv8z0lMXXUVyS
7O1AeyQCs2EqTZ/WY6XmOE89j+DhSLs5UD0ydswMsjZP7DbJArEl/PBf+13ZUVnX
Z6UcKXezZRbMSAXgqsumZon0mhObPwn3jJqodOHBwB7skKFwiYxkuTGMorH87Xu1
s7rQ5Ga3dWSUrpQdT1xB/Hw4ZKzq9GCVhHSsel3+q+5fT8IH38LBFs17Xp08Gtiq
27P6lhQisZi62gy73gqxfpBUUvgDccxKNUmAbq6EDREwWKNZQBwhv1mrqQubRbAh
unCSERbbtrrc32coKvw8yNGR4ABmW0ONJf+ET2iybM5vOQO1AX1EYxhhskf0kE7F
DV1gwQiD44Z6wSUW7fFCmR0FIe4spp076XAAXS05HzQN42qhqaXR5LI3rzzAC3Ra
ww9sgwNMfMGt+tuGCePNtjzB46a9SQ8wCi+4r/7QmeY3p5Hbp6n3dqyAQXIrfeLs
o/ImcVjWqffSMaO8WqJYod2a+spCzTSdK2Yrlq71C6QAWjAG3/l5TxTxXv4Sz441
WMer9JfrnBFTyyWvar8EKrqilNspCkjf/4mZcP5IVzexfy2m1aFbq1bDNdz4cLYU
1BwmKydK7GEd32+bh3gCz+2X/gQ+Iy1hcy1gOkc/ia6ghsJlK+Mg1gOb6boD6fLf
O2e1dqo0sj6MKHwJtp+s2IhAWM31DmOa3j87RERg6Cid/BJEjxhGYHc2JbAMbDHS
qCkAoDatEKYnUPJIohOfKYr+nRCsmnA2h+TXlFdDXBwXK8ClGSMcsiKYKV+I34nR
FwRglDKWbBcZILphh6uUZ5CU0ENIX/puZ/3Ge+lrpmOY3JGt+TJUhUkn0PwEagLt
vBvxEqAm4FYx+Y/KiyiyHyjkuzmW1PhuADSS3DKK9usCLHaQqKbSKH2iMyVgv74C
7i4u6TN8ZNxj0siG1waxQC6h8mrqlxxqX1UW/xdz8Eklhuy8zccXhrDnP8e3oZUB
sUtSagvryn3v69vj8lzHnKwL6amycNUiZK6FkuhDHmHv8t0Tfa7QVbbyRAWO9znD
l81jUu34iU9SBj6LFSwePhZqpABPuKgavpE7+lG08DBDKxsPVXq7MEMPmUR0e763
sY1m8e/Ti/JKddQyrIAqFLrDi/4shE9ft0k+uhEZVo3szyMMUSINwRM5q40RyGnp
rW/YcuD4DpagvDu18uLoMaKAovZlF9vg81HOorlvhOaldRMdQXC76IyleHVjRQTF
T4KuQmjnlLop7vjzbfQ4JeXvtAkLhVmp+r3TwXeIuYMIx7FdvhbyZkxoCX0OZrxv
ijhZ5Tp4ASpow5ufbnDp4MtHvIfJTU60zhz60V0CysLpe1HlznvPtsS0aj+Oqan4
YCQnQIUIiJHGw87wFDLF+tn+ppalwKWqyQPCaLVrf0VuELwHLGUOE1/sRxDg88x4
d5gUG1IsVHX01cqBWSIvW2+mEmh1jNzDgm7n05/xqweLxGGTc8enXpx1A2Amoy/a
FlTf18Qc8AESuUaY8xy0LECHMCYyeXeRcHjA1dkE1sSIgRww0rp5qd2gNxLWH6R9
q0ugFt6k92OiM/1bNUORPcNCmW3zJw98euUquRog625IjpBWEh9mS83cZ2YfgT7s
LC8vNN5VNuHP5X2AEKTjB3IVx6J0SnppIRRPvbPCUxznCtWGQWKaUkA+hvi15eFG
xOhdg3qBcx8oK3XJZIh1Z7OAMGH4AMoi/LDNJrfW+rj4KMmGoQm9N5Q9lD0RyIe5
b5hOpIj1dipljlzkHFberG2djvsP2y4UAF25rLQiv17z03iDX/R1/BdVFUnEaXSg
sMPpVjuNgqvjAIsBXZjN9L3dPG7EtzHv3ILJbaWD1kiSHRdbD4xQGA4G52RDktln
45ySiijWgAk7Iv7Y6Po5YhXrPpLvrcv6y+lFkAVPCZFgX7ydqslJqFmryUsNRgiz
8yo7e3eDLoCnB3DGgdo7wUOT1P0ERRMa5RYOZbDajqb1FMBTt7+Kz3FmbDzSiypx
itKXf96e8haxAdyDvSkNWsYPWl+ojjbe2/PxW4OtU9VNac7LQNrtAEh9nJ7lOggi
fUikcGqAu5MvHrp8dRZ/FPqtqeXeaf/7ilsCPUJQ0q6KU7C6WosyAGjdfAzDKDs+
yWkooQVtldqZBK0ASnPF0Ifn/uFXJtu4aeMJWsEOukpVme91rMwVYJ/17sfB+FS8
ivmRyoronK+g0knUtUHyo1hSN5Wmo6+x2Fjc/5oANnRDVA6Bwv6VaNn2cK5vL70t
kvZwBdKH0jQevwE719l2fGEimw56chjJWPLnkEu80IzmUx6I7LyWpb8c72dRksJ9
D45CVjp/38H6OcePktZOlZ9WtwjbYutSuyaBgHWF611yH+5etRQxNsiw+JAnyZPL
m4IlttHdRAI4Z0kvrPjNmPoDdlYGd1wEBQwLeAToH1+mr0U5bTNzH3in3+FJ0tlk
AlIB4WzbO8ry9L8t+oCyhKGiKCdDX/SR4nvT/uRRTCfYup/EloMg5I8xNvZyJ/iF
Tpz4BFFxPkvpbbn+AvYWzubtKSK8yTXEIT+bIl7/9UG26nFVAxRy9eXA5mzbqT21
l/Kq3p77MRKunqRBH25Wf62QNZ3514W8ipc5EEyyUDS9FW5KNEY1DFQzKTJSQ2tE
9Oy/mzurhG/2o/bRcM+GSua0llZcuezjp8zxjRN1mFQm8cCse1sCIKSoSBBRi4h7
KmA07M+W7jFKIQvrBjg8K4pkMQ0vWZXgS/pHBUtqhiAdZWi9o2LgmQy5Zl77yiMY
vooIdyy3zQR6swsz3BbyFjpL6IbD8uyhAGPSkaFwgIxEYVxAXiL8JlESmwHQDgh1
ZCqnFAUE66Npm+o90R67oOL8ypK4i3/ZK7bGrTHBEy6jO8LqWJJ7zERlaR62ITVm
u/7rlE2g51CAXqthCQ5nlQGN49A44ARlgmotnhXEzmH1zKjU1DFLpzbffZ1T1uTT
AujXOkaKUSzMNjXoqQL7mR9RViyaS7ZLwud3Q6Pc6va/cYImsb3yk5sF/KXDqxjA
CrLKVtStQJIibQTQPPI+DCsP85XmSOEzSFWYyeVMp0Y0039CQL1LXahMYqWPhHq3
Wxdg4pFAM+2u1nLTaE3RzdHN30Tg8IcX/u62u/Iopgj8UYuqbuYhnyjECPCJjQqw
N71vMmW7l8dHM7DdteDhs/HPdFbWhPYYvqYS1UocBh3ufZHy0jdf1uUSQ2YxYghc
aYkCsu590ActjLrekImPvtIAzRx5JfikVn/Fo0SIqDgSP5PW/NKk9YiIWJitU93u
7KiRhxWvb0k0COAo9jNdOFiSmNaiRIxdoMgmUmbIoQ9lzRh89PZYvt9bgyBjhIwu
oW5GUsBsRwcjACDP8RlEwthPeD1Ffxti7pKvvJ9dTJ/YK9oWcFsYBJGo2GrA+4cH
MSuLdD3RX8oK8FqMdRP0lHGkV77Ww35ldojmcp1HciSlAtLRTqqZsVEsk88SLY6u
C7KMvn3VNOUpRmayqKxMGTygs2Kevl1Xt6EgnFeWT55dZ35EubutBZQaYRE0HD0Z
G0vpqqGv1jLCi0BtcYsNKjQ+NBDMLt9kq3NzT6KnvhmcduDXMJ4bw2kq1cy55vER
CnW37uDmbQuUE+jpWWDETd/XZ3DjaEVqKZ1D6JgctKLeauvfblYGeNd1OwccYpwz
Mqqje5ODhAXdYylYEiROee2aFNGKVBlc9DvKWVDL65iA9kHcleQK/eHMK34M5nyx
9QHgGgcDcwvTojC9nbh3c+pJfanQBE/mIER2djTJ2podVf3iLJkvGDdaMoVITpav
xey3DlIFLlDu9jlr3IYXpIXQp5KAoMGFZT8Nbn1EzgUCM1bf7hRZIUFYhgJJ1iSm
Qhaqer1n6D91C6HMBP0laa1dNUOX7hgqAiIXHyBguzJeBDujCeW6i80fxuxB6dge
jyh72tSk6gpMi4PXkxRLI7fkw/x918bLouKWEpyEDDAGa1jp1gL3VEp0W/x0n1Or
JACYsF9BvNS5WyRhBZPG4fzqnlGYSiBWEUpu1+GCtev+4RKiG3HZ+1vpN4ZrQGge
itu9GQmo5KeidAUcT/zu7EWUNhj+jeAI36iMACd67WmJrZb2NSH+hKc8vabyg1RR
53hgUxJAKPdZQ9QjP367xTS+SquGMuIEfqxDurP8FhAg1oAUrZXIpEn+bN8PYCKO
a6jrvf5N74mrmrB9vMTE3Exhz8WMUThbStoyrBFmoQum7omxdrWzm5yM5dvSdFrD
BuoKFGYwwg98RMSwu0ign3eAlyq7VwIyI7hRtb4tC3nxF1Zq/dQQyev6cJxjf0vy
+fFJGGrGDp8RhdgcBMPplUqY0rsMxFQmvhYkeno2FB4L4dAQOPHT46y6BQwHbCgv
n6eqstavfCcgLC+SfR9NtAI8iIRYSPRBwI6m9UjoqJZ6q5AAxF2qIj+SE4ZiBFmQ
5v0vTmZP5Lax/oKQWuwwASEkQlPtqgYdR5s3jiXATENhWttjAlwGhM0msoxwN3pO
hQ5MJD3YokjQL6UO0kPO9rHEmukOd1u5/gFW6UqgsDowDZrQfkwiELgLFXLZoPiM
+cpjNXkbx+RzSEMw1uYNtDd0y8G93BwJtoyUyiBc6sr1E3dZnTPf5fd78MVAShR7
rwE4oVRCY0iZhZjcgHpuivR2QIgWP1jH6tHd59SJ3+hA9r16l1joYMc/Emc3ZIxM
oYhN3oTxYSXLc5WSmJM4033WbjCZDog+OpJtpzjdtfnbzVY9ptUJAyRvNQsXNt+r
YTmMY/iUXCGcs+ereU9jAuN8Q1L2B9Lz+AvcBXNAAl0Sflig9K3tD+YTlHQWru8Y
MgzNbH+jrNNHp00SwvFHxBrP7EXAl/TG6hQ5x104itRWzK/12mOxZOSeqStPGGTK
/TPme9mOkg3Nui1zJ5U7KitMEdPLtWKqLAd2cZkapDrGzRGUFdmScEpuZI2RXA5a
Kcq+sSfkgiOW/M4YIRyOpNX8Rggf/lJSTRarOWbr9aC+6uk39k56o7t3aPdbguDL
MqAUcWsh+3XSES2uniS7KzhuNkFMk12BKSPGfWxD44PwEyztd7bz3RG2Veno+QlY
dj6ZB2JuKkAVlye18jlXNKjjebVYOT6pQ8RCA8nebPhktdJYX9Kei/VVg5xxNg6L
IMtgRQE9l4BhhEydZizxEvttlJqDrskWMFLEC87NHoVPIhV6BxMGZVhWrXmjzFR7
f9gcQS6eZ/DOMwc0AwdPANKEeW53x+YEBFd3CYN9pCuxpSV4S3NAqVyQHyh9ZDKE
DeGTqfWyW+WSo4cZHxgw1c3VNm6pCtJ5WviU7soNsHLci+KsEY294PvUvGxltwkZ
SUfv5FNoS9M1j72HIPBoAaZN66F1yDbGcbK9YiA1tF7iGArRdt1SEYpYxaX+Kn5E
lMPKSTvLX75lmiZVQiop5iDZ5s6OKBMU78pwQQzrxFC3bzbjPW6N4PXDInYZ0NBx
/O+TN//S2q89Q4IPOfPe0L+jZJlg/mx2MEALp4XKORwuQUzPWqdjGOq+qd3pt7xr
iNXfuFevcQZGd7MfbtzX72ZsVw/bxFvj4OWD2AAHND5IAS2pzjj8BcUDfAil31P3
6NsQxsCtx0aPYkI1B/q09MH06qdHdbdNzM+2Nw7rT+WR14G1ffvmIlOwfdwZMEj7
jyZ8ZWUFwFZT2T6KjVtD8qDHu8YUQiW+OXFQWVYwYR7HdMgnX2/oV6IK3aHM0RzY
mEounEEltdeF0IruwYARqkVvIG2s9WTCnQtfOWc2x4tYhNP/JeyTMdFNhJT/UeGP
mVQRzyajRux47XXKlG8onsZEYuVTV3Jm6y4g/TxkbKBZvMeuPkk4EEFqA5vwvjAG
cok82VLWtBFJaIyt4KqBzil2VkSMQWmYT8gJvgWWUU+ZDqMcPcyRJAg4jsQ+54+Q
TJ4FOzjlYsj/lfbLUZZAnm85evHbahvNYA0hNNW1Knsh+gs/Cht5G2uWvjcyCKcA
tqrZmwrd8dfjVWxyzoyNJhRmJpw0bPCEnEzr3245xPr1eaXDzQu9GLWNfso1ZC46
ptPhIBN8QW/cQ3tOT64+9wO29byY+KIcEgYJujPSPgDvbkUOlNRdMWfF8nGOJ/z8
SwjBQ/clg6thzzWbd3iFUSDAVC0kLchEUOhEaStL7xyDTId6ACPrXM5WdD5ODJ1x
NdS3LhXDDMVZywBEgX6UIBUuSCiZtbFp/yUaNkqQsv08O3H+Bwm+a84VOKhc7ERq
m1YhEBagp9QZOTc3AWQQHRuGrTwZlrzZySaX47i+QXPYemBVvCmsLmgd7/7Msiqm
Mc+duAv6n+YG/zgfqSU+KnAIeyaVF/HYjgzCNx7xJIe1VPlxJgWOUqhojTUSF9c5
jz2mdXjLJp3qIoY8Euz3zQZKFXxIvROcnu+lmK6jCM5+triKx0powpWb63/MY13O
PNVRN9NoHYs0D1PiAh41qQT37n9DwVeTJniP/uo8++zTRJby+rOcOtKHyT/9j9QW
ls2xqryqagNPjUADNREgZfrLXTOIGgJTT0c35lt75VSG5SMDb00K7Y+LsubIn5VI
RG8f3NPMxa/K/gatEP7QOffCbDc9niJwlqU4me2PpZNPlym4s8E+tmC8sMrgC6ZL
TVmN8WrEgLT4DGeU18UrRBBO/9ZU/rOP8hFIFhWfv7RoCkiycOF4aqPxRpRt4hiP
d9GhxhzK8DzH/eh/LhGHGUiFQwfnzwlYcuAallmg0HHIrSjxAhcXDyS4/UQUpYjz
9pVQT7KQGnNcFsaPizD41KZXq1B9DBDqHzcl/Qu0VjDCUdD1DWRplH66+CT3Bekt
Qw5QJ6gw5qc7VitMSk3upvtVOZhJmMAJ+Vy6EliZNpsWIPlrPe5g/EetDnIguU9z
qrRZxsajSQyAMdjB4sdmDClH4E8tC6R/K9vLoOsKgEm7eymIdV4dsBWarjIEOduG
qpypU8VMY/Ta3d5ZURaqeT0Kp5GaUs7aSV7Kns1OdDavIo4IyWmtyAXjXuQ/WOr4
exXEeRV7NrB+le/aPEaqmlhun6Cj76OJVa+gxzlIg5kfzdiQ5PFi2LY25dEJZG2M
zhcJRdpvY9cbWQFCwZI+zjnxlxMOxPFjG2MHZir0/yldQ7vComhDQDHYZu07ziJE
NDPKuZ5ofeyxFoHm9rF9qS8SLAs/lHBWKtg7DRoiDaIfGvPHhZWD0qkU5938A6t7
XmwHRxmyRmvm+VJcp1a3Ow/W6ZfvVBThsIODOZDae++TPrhfD+uYzSwu0XGknP01
cgQm5XmQSve8Xi8X2H3Ff9ka5c5SA3FRFDm6euOhT1J1rKRK0NQCKL5XPuNt70Hp
uDUcCyPJp5AD7PHC52xykQWtpCpg1h1SxoMTpv2v/b5dxcHKjSGKb8wv4znjfFLe
yROh1H3vJQEZzcEB8itJ61XZWC1kC61Kajdy4jcN2G09H1BkLg8Dv4CF+81xkIif
UKw7CdkEdawC4AAkLrzboEe3w7WOTFbYD6GMtrqjsrPvfw6FJm0MgidqB1Fiahx8
WVHVskLaqE8t0+YbHo4EfV/2cCDyWCy5/C2xuQWpQkMniBq+vnCMBOTU+kyYpzCZ
i2cALdBbzg37pRWqFx9H6k9mo9xyzlpFD2GrB9zSOryMuqK6DUgpezpZIiRB9kMx
Y5IH9MOUGOkOdqdhHWKFt5sYdYcQnWQ0tiXHeOjgT4zatRhAzHg6EB5HaRM9bune
W067bbfWn+LFIC6Z/qw9vPCm9NkLCTZcJ23eTMJeEgnvtsrwNdyeoIfVu9giVX+o
QrmyBdr26v/+m8j1RNoOUQk63H8+cm5NBuP7TTjGUsXQj9TzjsEtiPVwovApcUFa
YCwctsUbqar8MPPDfwiGJUAgriUTnI6IHoOEahpE875MFt3G8H/leACk+r/h2LT+
t3xhsohhQf4HNzIEBjIraThgBgi/rCII35dmo7MLa9Nv0W0a2I2xoj/z7MC3UOTD
9ASD5TTLilGQ/CNN6B7IZu2UW6UAEsXMx9D1TFhVlNpN3neRyYzU2zk8eEqm4it+
Dz4Z+NIqtqbS9ZDYIaQVUL1bZmsqGzLabUxi+Ml1JchcYr4lps1e0LoY3jRh0BMl
rSJy6mTtfcBr6aZ6w8GAzI8ZB08iDSFNJbq/KGttcuX8cHoIdZZbbJ+Dj+Dbzm7K
PsDWMPcD0T6EXX1s+/koz3Qwby51j3LEywcoxeBJ2ck0Pn7Dc3xF/lHBHRcCSmD7
J3CzQfhrNIZBadziK3kVGKsrrY0A59vwTOf+FONY0oc5O3nhZwtR7aHC2Q3ZFpxP
Qk9iQv7HDgT8UvDfKcaDct7M/lEeuR3LmBnD9B0JfKHOlm7jlYL0lJ0VsbGCnc7z
JQf6t87gVwqvV3lfBW5NhZN1Hh1duUO0uWZ+HHS2rbzLZVFJpUdL+iQ9mSyri2RY
mYoN9jrtFbkBhx/g2Ei3lU5aSo9BcR7OxFOlR/PP8K3936VfIvnv2e9dSmamA2y2
T+kj+d9UFxef1Ldf1q1gx8Rk5y6fyis/0YcghmLdCw5lzjT8QdZDsxrx3QBfesgF
WX3luSg3BHA2ORtG4oTFvvqxTgtxEam4meOhY9eVeqDPlFSsHfuaOo2Lr2YGIIhg
wt16MifD47olNbnuN4VstFhwKMrge294eC5QJEpw+vfZ/iGV87Qm8Cr5WKCNjGTk
GpMcBZ46zaAfOHd0SG1/yuQ4DmxLTaMKq/1T6EU4ogYmZGjqy7LnRPHsRv18/XXG
4hTJDvTYNFL2u4aU7RhpFLGD50OX3ycgj7JmOVJNjtiWlJo2/HTwzESeDz/4G4Wb
f3/x4IlBLxVVM9EUrHFrV7anF1EwazWfe15p255R/7wXzXyfZk/+2t4nBvSXZbHJ
22sRstJM9RTptBtdXNNbtuq4jOALZIb1eUUxgNwpJV9gtU4h7e4S0qUH8qxmxOGL
WKVEMPO7tM27fsW2SB9gfSxes1W+hRbyqHKmsAXF9MWQ5EZUYj/o4XN/KDOc83Uo
Rw3W+Nq5dpDc/9+htKqwxIW6a0orlAW/RtlcKfG49Qjb0UhXo0UZCwELtJgmHZl0
KS3rToqo7BHQrkUy2x7xIxtXURXRiH+lBCQ3nfW2bFUKMzM6Zr38FKPkMF0mq6NS
Z8E4Ci+VNR0lB+4Ux3p7i4TUxIOfUkUy6S567/rIhphFLMKQiafbUnadR2lIM4d3
C2qnO7OBFO3DgBniaCCTpEtSqUcDl3Z0eH6YOp9BeHrINIC8s0XN3aZSVlK6h5nO
MlWktwdo4orjyBZGRF3o/wvDOXumc2xtyLu+M826o3QJXdOxtOSOop+NRhAWutDU
OgEy/QnvnIA3J99eLPAfDH5UNTmBdxTytb3gcM1QnCF7PI57OVbGUYfiO0XLMwKr
kUxjp36Fl6+73ny2PCEOFJSRU/WCY1I3JC8/eTeD5/HD9VSUiwSS7XCeLCqs6PuA
19NT97aEtAoxF0Ijx3tflVeT2SJJFZ2/U8FvLBXdCEXesVVCE1teJih98Cp8toV6
E+VXVgP47xvIxI2L3x2hEvdv1E2tK4hptTwMIjrXoh2jsX+VHV2y1bktIPdc61+J
3Gk5Q9+obDmR7zox1Wy41QRBm4BzVdpq0hYlZ2rW9Hmtkzahl75VQ7J8Onawnzhe
BcBAG6sMk4dMKtBeUEWgG08MQjPQam8pw1EP1rNWBTFHwS883TtkZCkkJo+Gp994
7HcB7YuqapWEmFm8bGHzbXEUo1Ve/CWF1Uk0Bi2rff8CDf8xxQbzq3K/3O1M9g+s
ou9hf47I2lbOEoE3mzqV0ZqVRKfcSHnQWFj5qC1dOBhA/vGb61ztNjFO4LLcQN79
jWa3NSkLghJ7pnP79IJjPd/Bz5vuzZ8rUKw/Tw9kiZ7l9WUkNJ0Iwse2wWUeDdHb
sR22zDP40+B5QNI0cNWLafuOBnH0bz7cPA5kBZrhScNigWxrc10asgDzp/TpsjkN
7lVU+ad0sfY7mJdAQzmWx1aTNpUy36BEVh9RLjGA3YW6Le13tbzJVpWWEWclRrnN
Q3buZFBOpsJmLBgoLXIXqkejHtXp96mjfPewp6tEL5yIJFonBPDfP37u/aZfDnxf
VpBE9obmBylek0k0XseglWvpw4VHpofApidMyMIJN3a5A1hEhFGbMFeZmmJ5fLwC
TTIYZGd7NLPiLrhjNXpdS6fB9S6QMIdY/mI1Fes9oBmnTwrBtm5Vx8Djn6DslC6M
Wk90k+NQG1mOESw/RisdB/kRQ+xABR/pfNuI2LlnEFUe81vlP0vhZBePo33nCdBA
1FrgR87+QuTfGHIDnwRzvCy6Ya0rk4AMsaiNqoLzak/kn0tu6Sjc5Ct0DbXb31pu
kMqY7c6k0YZ84AkKYOb0bbr+r6ovbfutSaom9TsKtqDmqMhVu+jubiNOPeUsyHZk
HDGXJvSFA3UPvVo1q/Qi3tFRrNkuV0IC4B2RQIDWoADAH9TRmikz+NrJx/BRl60r
SJ5Ev07HFFsoEhVYKxXTGglLikGeBrszWMKrPrG4i/mTme1yhzxRdkfHqMFVH3u5
2U4T/cGDuvx/RYXioagn6EsUSddz3kANthZiq/i8JB+PBv4wsPHjE/LmDql35jpa
rELwN37naKkH7ksWuDI7afvZteWjkQEOOK/SR7wkPENla/6RzdlD3p+SHoor23Eb
QyIfQMOZFNYW9yEZh4OAu70Cu5wQqEOO9Vwc9kFT2ACL+3FHPoimjvoAFVO/K9Zy
fcq4/H94nVunVDe2ts6BH1Jx6BfLHlNZAdBD4lCABdp+dd9WViNOmrPMgdB6a0hr
RFe/fnS5dRAvIQNdXe9hyy8ncMK1ynN9qFayKNRz0fYaisIpq2kW9Z91QD181dWC
XicnlSkG1DMwc+5dMM3cRIvvKoRL/cEl0L2xx+oN3ZkDTbL7frOFNqE16qViiYW7
/eGmoNgTt4nAO8gDz0H2BW022fyk3ykqW43jitGoZ7LVieFbEXmZ9dd8whKOeafa
zWNdn8OLDgNLooNDrB+C5DSiyNqwKTi2IxVQdmsrO89kDnFyftrxRXfjtp3GSWsR
HYa/Riw2/K/LXxxmlYSH6Eah3XWyso2W74mHXJDyIYWYHj6cXGMWlEZ7oqoR0j4T
G4AC9FhjT+lG8oIHcnK3Se77M/nG8pDXQW42R6jieb9BczzK4Urr7E7Dwpf/vmG9
DLZub1FitzpdEUf4AaqMPce7t1fsZjex7UnYaHPvajRXDbvkfWHaOyIuilKY4lwG
ePhe2fMO1atY7QoZ8a2gVF+H00d8+Zwce0FWwckY6OkeN8G+iV73KbNmjEogmPTr
C1t91xOcvBFhnbZGckL1Lu6OQvC4AL3gZjZVhUWJpWNos4FlzhyY4z7nnnN/uwPx
8jxmtY5GgjGP0XfBoz55R+cJ3qo2kFIREuLGmd0epjbpf89nzLLRvTMhCKt8omwN
TVZOkihY0SkA1VWG6nHFW55vehrKEyhSONfuX+ZvXKgHctAXqZztaASp2FIg6Go3
wCbFPRVw5WOhw/3CjE7/4XPZJ0CKMgHNjR4FC/TvV+VnpzhnUoANoZ+7G1iu82S5
R13O2z9q2HU9d7Bixg0M/QrkZQG2LjVXXXcI4GfNi/ItfJNknZcToY0T1d34RPKI
8WMMwrFNCXcpRYiwHeT16jOojXJNSJxgyfaQe9cuZFv8sHpu7Tm54XtunMM6HkDz
dbzwAGwYqnOpyGGTErhfJTjruCqzdFZeOVyzQj9uZW7tcF5ueSsQOJEryoxhinWq
hkmKsrQ7cw0/lXtL0ami1nVOEG+b9XZnJKKr4g0a1ZSBnjB77ZhqDJAfwyQBGinW
2JXStfzC4Mv/QfxrqA20DetVwvhEYlVXQE0McotiSvzTSZoZrrfLhj6Pii54rxA+
zlRKb0hwqWCrdEkXPrCF41GNNc2wHO7JL8LDjpAyNoumMqIWhEQi3XnCTluwj7Bg
Ui6//3Rm8wzwyvgctHTNqnJ+xpzu/HtopjJLulHMUJUwItoEin+TzLfXcmFwm1Nr
uR2vDiCoWPAXfu9EZWuRzYWvLGSfnCTbE/NnAKx+9nW/M5A5qEx5XEIx0sev0fol
HWa6DARFPnmiKe5QFI9VuXMg/fUYHA2gE7DMI75qvC5RPRh34BUG39Aod850pUvc
Xb5VrrmzSeUXWSCsKseotD/g2QVswInr0lnscmWQ3AXbm8QUt1O/S+6RJgns16Dh
6U8IYtbvQ/4ZFnEebJ7LjjsXRzwmv4UjfUTTg4UZjU3xUVSGwJndOdz1jdtB626N
U/WISDt5syPvObWv6a/aUS8uAnJjVIMWAjU84bUQmt/OIhakOzyJ0qNHeKFf001e
3YR02Z+8K2FgLX6yKWDBSCTNV8AB79qsMBIdNwE6gAx85/vx1ywa/Wl//9zMRLFu
EuM/9gN9ruv7h72ihsnqPrUd9w/HzQZHCrCCsTG6xbtYJJspZpNLJrRMVBdsjWoT
nUuvSOZaezACtjhxIJ9qqp6z0YomZlz7m1L6z9fDS04OtMe/lcVsbitvd/ooYl0a
MswsD/qrp7E0INgg7udUO5HPHnNDD6oBWi0UElEh/JbCQpqTY/hjTma/O5w7lDAt
MD3UQOqM+9luQ5gtmuyyguoNnrD0Tqtzzq9uuQglV1LBRReg47MDG5ethe3fIhQd
wUG8WSAyb7I44NDRQWmJBj98WynwDQvhsx0goxweKrIIEELmrWXMUUb0o5FDr1tq
qumlbJDKWWtRWTNp+e4WOpTs4bfm5h8xQogwzKHMLuA4/zTkXmJZZ7Plq0zBj1SU
Pez4/DLw2b3KPJbq8H0NFykf3L+jSssPzQR3Rl12vpsOS5lnXWYIoPK9iWKHN5ug
ZlBTeeKEM3izCJEGn0euV8Ag1ZWT5zaVLkfSNOoRKe9TMypY//eWyWzT9ltlB5/m
j4MFhqi1z6v/0tFcfatCcxww+t7daFZjpSrIlf2h7JC2I5ad3bqVWF1GiHcTV7Sn
nSwsZ4NWSHLVgTroM10T50zSwL1+fPz4OTvAUQtaZg0yuBl43LjTroC8U4HISwaa
/A1c/V9ll48Lg3+FwIyGsKHNYEVddJH+O8ZcDzkr/bl9esvE3Hh2gq21DW9IjQTV
ONd1CTvm3Euq7YySROKf0oNeXd86Ie1XcUvADNjC/pPxlUerkjEIy/h3YDVYfEao
upH0+bAPYdJlnT25hrzDIomXnJVRapyHpw4hVoP1da9wIvZ6pNDJgLSx6TwU0AZC
n5U5H0cYNmvygwuWrM4gUdpUzVcOb+ELHFE2Qo9mS+Th8LjOIkexMgoSKfJARYlE
F2xlXfend3A+1TeIgJNJPuZUrdg+wKJ51huM5SKyDiZte1UfwiG/IjgUIxMr4cz3
8RIL4wbS4XBfR0EtJL5dLrEzdJSlLWS/D2qDFyChW1VUHW9DW5ahcxXpHuMf7wBN
47gyJuo0dwxMqjLY4n76wjuEGywm/hdfuvKCSi0I/E3KdqMuC+wIheCU0JVIdnKf
oudOAqgfIm4NVyD3kXVQvDAj0EBNskhLFVm7A6U7RIi7jWajlGvJ9xVhe5Akze//
d/4cIdxrPBnCc/+BlpbPrBpuRgz5c5hz3bpl0cQDpsC6F/XWyoGP0wXuD2xtdgFR
xqUBqa5ua420fhCEpL/NAqi+jdRGesSoTK5JXxltm874Q1Ey+qNbVbg20y/ZQgMp
KANKR53yRYW4cpPTZwa96S15jHAdPik76CqrXK5PKlWNFOV7CuSDEO9dtOT+if0c
lXbwZMxkd0OCuSWLIO40azyiXG2HFmUWVG5ZfiT/NATdo/MRPq1j0xpxoStQ/DQ9
YCnh+6GAJ2oFZg1jtriTPRoe59WCJ3EAN16fHGUKKDXofTyVD+EDFHzPFhXfg/Fb
uBwQ3CDG3eCK9tFE2x2mHUFwgCIowMXAZr9Z5pUV4XxVi9yEVC0SCCWbUgH4nyNI
GG73HmRfW0WVDoFruNBjhCp1kuW589PyMFVLK4VFmv0WmmeDXiqJ+CVRoS/UEFGx
hsKuZlqZkCoWA33YhW2qaaXN734Cd02+sVy9KXAsWE9KeCEIWpYr8fd/1ulejtoL
DuRs9cwQnSF9pUwehvdcVPZsoLOyI2od4Z7EiJ+vSG4q5eUjlrov2Hf9rCtBYdFs
ZKDJAn7JPeBu7xufzuDhdRyCGvru43Yb+ldvAgB32xgS3Ro4uHO4otDwf8T/QBgx
gkdCDNoYp7AMG61SaDxjHDidMgafAyIKG0OsZZqkbZ11HBYZWe1+wju9FwAHW6B2
9qqccI7W1O5QSPS6RR0gEQ6Ill/OWlH5ZYIx9Tn15/x79gUpX8aDGJEFdLDMiw1F
YNVepTkhADEK5Brc+XJYT6CAHrS5AdvFbuMpCnl2NWlxLaqHN/k+j6+hfRK8+Vxi
O6MvU2gkQ9FOH1hWHOE/l2suy13iv14EyIdnwRTL1jR9ldsdmo6if7lstBnw2MLw
W4uwZ23e5qsB2mW5u+xmPUXWyuC9Wslc/k21MfsX0v8LDVgNe+ZBlmjHjEZvR2Mr
46YP+a/diVCUzQbcjeMwt+GhiCCGjPEt/miZUdOGBPDtSRnHovNBL6RoMP09YSy9
QrqiX3LZI5JwwEm3MQ6RahvJ9q7ydLlaIuueLc9ELVEO5KwtdMZa9nK7/CTAocdy
3ox6b4/xF2lM41jUiDSByh5hDmgg1zvdVa5/Jpmpxd2/Zy7DUbhs7W6YIqafwBvA
uB1bRhpBD2SKic31Je7tp3QqGGPQaRrr6k5IJH3uexoZNZjDiT54Dh24VEXwrbZa
ax27zf51yqjt4fqzcwnZHiNtU/eQoahVAVdEZsrgCbaX3ExvH/1jPZW0dNAslq4L
WjAIg9osEvQpuVAf7tZ99rUbTNmMjCVGtW37EGKxQc7Dsd8SrjwGZs2dX9hejPa4
xgnRy3X9tfn7UkJsCQ9ZXyV5NMhWwMBKMYjQGkbGEhEGAjA1L6UNosSRBIpBa7Q5
OqjUGvFlUbjCQeHa97InlxrelzEG3mP61NPaH4+s4mtaU4LQ42DhWB8O16DgyDoK
qsFo1jpcyHQHvYEIoznXPX4Y8c77zCtUNBs9bDHqGVFFeoq8PiHsqadsH8gnxPiu
yxbiQ8Er45mOarodO/8iMd3pFOz9IsIn/buJFXYVROZLM+Il+kk39ZiCk6vNwSeY
tGus+on+t+1XWA2+b9mducXg9J1wdfw9X/GtBAsW2cEcv8lHC8w6iG9dLB4u5LR1
s5HVr+48/5cM+fcSpekDxmgGhrxWc5mPsW4K9iwiVCnt4zptEPU+rvKUDEYBt9pP
Nx7F4bummOgX2UJG6wf6RoUsVkG6srwVD+mZQu0gnjqjRLCE4g0aAhMfRk2H0qxM
dVz8pj9+zx0UOmZEBY8zNsoTlReiMAx6WPjkMfSHziNfSu6X4Zqadusvnm5Hc6Kf
IWCyVqnisEEWZuqk+4fIXYfIGlZVrFNjs0FjntMNh925//T7HYJVT0B4j+iQnN+7
D1QrPfKugn/uewOTISqGTDG660c+Zc3zWB/IxxJUCnM9xzfM0io/S9rSBc6vKi1s
8/aZKBp8jslKSIX8djTuZG2EoHCLgl0DdZeIBoeZf7nsXITEpDTg5/WhOQge9Ldr
2rClhwmw+CduhE2+fMmZYvTY0qzDuzrIG8UEe0A5zQHs8cdUeh7JR01H7Fwf0xvR
z7FJAYU8ba+tpx1Y4ysJFIFGXIG34tLwiCQgXqlOnUWsXJRqJ0TXpNY+gpHpV4u5
G2hTgrEKiGVLUrU83oRlcrIGC4nxOx7DLifLGrH+5RCOtvdsucgwpUKY2jiCVU4N
37Hmi39as2Zh0rdm0VBi8jDy4RZVUMXWAey5aFXHSrgSTUWdMyq9CoYnBAuRJ0qg
dps68J5vU0fAOJ3CL7KPd/PKqlu+SVZnSxbbFBulCpQ4vzlQf5pfX4PWxx8AhS9Z
X7ZxaNpOXIqfiI9fymyQ1OzvyCHlca6h1RXaUMaZDQPQJXG/K0uLDx9s+tRWQIy0
AyYRhP2EVn6g8cADwTJsytJX5vXli0i6+gVUk3V71kSJBvPuNRpIdqDk1ye8uPR1
MxBlmWKoi5Q+NhUZT0lyTS046H2js5mUOB1Avrx4ciVWUQG9LF3YAmGc4jTMi015
7K5BYpC81Vp6IhLqdvD04O/ymqLFmMXsS7f9swcDoE65c+lWXKowuX3oReSoD50b
30vA6glvQrh3LRkXfjrKCVz/TWY22ZukVXC19Vh+b0OKTAIawrOQhD7hyP2b/WMf
4ae7r4EJXrJfAePAwIK1v7H4L+NEX4F5OrU8vcCfww3y1VpQV+PCrg3dilCJCiWj
Dy3sqcnLDpiUji88MzmsV+Cb9hK2XgxRpJOpzm3+cwDehzak8cpjffV9ZmpWQOf9
2O6f1ZiIwhM33clXkrW0bmy9wz2ba2A/tUjv8m8OUbJAQsUXauq8aDsDQ57s9YiL
6GIHnw3ouQ62NeG1HA26xuy2Yv+ag16VC3zjgbe1PVpiU3vQWfY5OIBQ8zqLc3el
m0l5/W8f+sdqm6ldHii6T0mIaWo4Q9G/7u2HCgMttHu2j/xk90TItjzjcvMOdKMs
hyA3HIG7K0wAHJYiRUjR5z1/gaGerNUbtSoXHYdduM9jDnAE8opMl4yv1UpOBpX2
66nwXXePfII25ou6ldCeQWb1/Y57WiNQb2GPM1sV/A9j7hANkNQB6kvXgML7hgu5
8rdOYx5n8clTHUcVZqkzILpT2BsuQwscraK4VbvUV4pryTg6ufmc1aXre3Xb13Uz
y6NVyc8XJYuxwf8kUi2L3LYV8P1EKNJNBafNQD9r29RSbqg0Sj5iMGmQ3MILXWlj
BtmDsaZwdJRCM2Vvki9NS648kTw92p+8CdY/gAI9SbriVqAHkrwk/hNtO9dH3l27
V5F0jUVEWMnd9CkNL7DVoPTwimYO93fche2FnyOEEy+xNFaHnHAl5ZMlxVxaDj29
ONpJ0wsGKxJYKTtFQWodHZfL96It+JUVpU3yiIEUBQRC1+cY97LO6lqjvX+q12B7
EJGpz+vSlZIefNJep+gy2INvAdzhZQUZ+D/zfqfg/ZGI2h1m+LuEIkZZdeHY2uRK
zjuJOcrbXsIcSmPXBab8YqSTGD24k/VGeVfEgM3robQfYYVSnuqn0/v4gzUSVHhJ
cfvfNcvCdpn3OO/JuT5TivRzS4dTW1pf9zP4z/5BjXpwI0QBoVnLMcUT9hVPgpYC
kNFIY89kUSEM6ivq8xHZg9V35otp/EkGitOu5XRIDFlPfsLosM1+GgqHhGDUZA9X
rsiMkS5/jpyG6PnaP2/r3cvtN5Eo8nzzPp9DUvdY/Wt8VUQA1cMBxhnpw1Y8Rb0+
yWKpQY6a69Ze2LYRXJRPyJw/VA/dP7RgrkejTFRrRphXyOE2v9bK0lApg2FVphMu
LV6XSLHXWmhdFqic515VeWfj1mkgF/2FMincu1njdYADCYOBBpC3xS02lVDvydp2
S9aGLgua+03PRbcVL4MPNBC/ZfsOKUZDoe78Gle+Pu3tpWjKpd8zXGRwo1nMokE8
+UkCQE/aYDtaSoWF7VziFvvHv1mIqPG4OcRnUnc28Nz/To9cU3bqmyMa6fqkW+nA
cmShh3UCipau7nHlax2ASAV+Deg744Dd3rFWg37WRcHVNM3cUlofs0Amdu4t5LIv
OQEU/l4z3qXpgg6fK1Bp6k+qJJrZxqa9HaHiyhckrE+nY+K8nCGfHHgAIm417fIc
j0wC5xVDqW652zTx0/nURjwU3W5G4CAM7m1bYW8GtM1Qdwu//86Vfsg0am17i2oI
TCQLSN10bRKm6YembzLGCeA/DZaYqXV7jYvW970RbnPS//famu7lWu0VtxvyPBFt
jFGD+1DAHOBPYRfNigToWMr7w85BYpZGqEmY5QSxTyqtV5LZgyY4Sds6FESPlwE3
/MoEmXKdUiror8eNSHb3wCqpatUqq8rNwUCLroW6KrKas0ieSjjbdiWGefhFMWkf
XUrhOlAFlWMK6soD3Ryt44PJDBS6OL0GtTOxpFky8W84+9AIWxuHhyl2iC0SksVW
FeBzEzd6+snJqRqMjM4usCNKnTB5Q5JstMasIEVW1UwY9byFvBEm1dSmry+vmzkN
+Rzze5Fw3ViRbZxMsOx/NTX+FylkyBmhsQmnqVNn+DHTlkitEAZ1CV66lcfFDTV9
xSn2L2jDPnU9JnmO3Mk7vgPVxLdSDCMOVCD3E4x2K+wQ2Nu44/fp6Igh4Zev91GK
CHxFL4qhBnTBoNnw0V6pYSYFtkVh7OfCLdj83eBT/Sw5NPMlc76wbhPWZLw8xE/F
NwhwpGKW8OG+6IzA6W9m45rVU8xwlamEqC2otvLnNl6hYnnxktdL4m8Uwdi9jmWB
yE2L4WQ2U70truXT9psqmcy9deC7zNRUfpvL/6iqiy8DlyM4S8atlOmgfOGoFoR6
Uor6fukzQ+2l9vw93o4JzA1YtrHtRPBb0RIlllcvakCXXyUfIp3C4qkz4iCp5pde
oZO+JQ88M9aY86xRxEOPn/zH2OCLulePNyKB23SIbr6XfU8RVONi3pWVsRASIUGt
MXBniX22yrbZs7q1IIMa1/rqw24zOEHyYyQwjaNP5v+89RYgR16dOAAK6gH95tDr
zVj7eZhjvhNNMQ46yhJ6TnUtkuWC6AmT2nboNgfkLulecOb1QSxyYZjrQlBsBn7N
zmdpcu+I19jt8eb0AnbLRpZtND42OCy67QwuzCf0TqxUcAh8BC1Nak3VTP/cZGWA
PzC+BdLOUuVZ9zZHpSH2EoRhDxTjkwx4tKYPdudwnVE9tTLRACEhqt3JQsKnQ9hz
A6kp7rls16hPZ6QZowWVu3d8WOs9J7FWsXSCmZJNf6uuXY+RncDyvbakUvrqC2nV
4VuwIbzQ4eW6nVbEK7DDuFJdqgnZ4YCHUpocoTknr9JzK9mNAIBFW8p7eIX6TemZ
zWQGxBWzAf9j0lji1Ut5GhmKrk/PIcz18ZEkuL/nYek0lwDu2tzV91GaFEZeSlxK
G4spob7deNmLMB02T+ckSK4qsl8ztKCjsx4pMkKyF+rWReLceiHYTW0YdmPPi5u6
bfRQb5YRPLMi9nFivqvOhoglNLI4IrNjnbH1AeSw/g2e+krN8tEHajzJ5LNm7G6t
HQSugqZwfD95w6bxLT92h+JH2xa219LUscMY+KzYDCxoKnpVocvQlKdnZhEEE3bm
UBbn0Jr2rNztyfd7sMYsfjKhPiqmIaKvleVJaYDQ5a096ZAJj4NNf+5ez7l3L6Qg
79CWkInVv9/9z+5W/CuVDGdQK03b/vpcWv2HTaFaJbzd3KqPZuHWmtTaUienVmuL
oZLn8y0vwO+1TXmpzmDn6IMHboSakoO8iIPQZ7iTxkqHOlh1DfSizeQQvTYBLave
giBVQiKDouZr7dvpG2nmwCT6tTP/2D7spude4Z4uPkoAh7VRxAOnQYu1oYYJYYi8
bysG2itxU2QJOaC0vMhEYiaA7qDjDDxIZjJTEKpXEuVZC0+YSb6+qC5SE2OhlttF
xrE026e7bLg3BvgWyTJVyhg2eVO8pLxCQMXl8/B1WRQgYvg0takT3R/Eapti4gTX
NK3TFikvJpRSL5MkM/cCdx3FTY2jsa3l/bZ54yNZJjWgPDpLOo8t9zktLlkOlgBE
u7dGEOt6D64vcEcjnBJY6ZkEn+Hx/kyKIt9jjqlCezOL44XXBz6Sis61nzKcp+0H
IJ8KMJ7etLWx8IWAK6g5vnZymLTdQpsxK1zLrzBQBMgfBmKzglYoJx6GZRdHkceI
aRaT8X+tYF7xR/WBuxgOMaxNFIZCPHYhPsfBt/cxJnB62Y40m9aiUvyUnJ4dvj7w
mzQQILoW3Vo/rJ9faKjd2Vk93yTT3ufulX0yPEBiYGqnoWPpHJZg9O2pH9IJB6ir
JPJwDH4JkuuLrEhXkqckFoLAbsujxgujed3s+pbH/GSi2t6tblVNTyIh95iVNPwM
Zkbg0aIgckN9+eQWpstSRYzb8gVEzVxYcSsMenJxPnG1z2L888Ix6UlZmhOiw8ss
SSh+ezpspSAJGJ6//cL5gRhA1dtmvkUQaIlQrfhmFn1ApsqkFsIz8Q7Q1YyXOzED
ktJdQglPjMn7F+cCVLF5bGY1ctOce4S8gKR9V2nnPWjFVFfpsNlRw4YDB7C8NYxy
ramRoZEktb/YrCfKdYeK7SLqpYednLRnoZEPHCNA9QhMapDzLvdNLdyfSBVJE1wV
21jqQ0X8VYQUIKPhQJCYIdwtnkR+SW/IYtovTJteZNvB5mJGFT9lG9whs1xR0nK2
ifaKaD3maSQRt+d8Ifu57Htvh4AGiEzeDntZzGmaVJ73DD8FyZksvNzoQKaKYqud
k1yKBoS/SMT8SdVba3pS0Z2JgBJ9PKHuuCEjWHXueoLMo1mH2QOhB8F9QiWN9y+P
3LlhTOI377clZEng7YdJkJ7u+1uqoIFgBcuBpptRb33sUUYnqgE9YWxlPeta5JRS
Y/zk93cw0VR+t2GYl8gIiyuybp/Nu7SjmA9kVglb8xoPQXFvDq5BHJtLR7YxW5XI
rkuCSMeOyye7AL7woeDpD4J18eJWdV7EYxdv0JlQm6iSlERfO4WEtrYkfSPtQDvG
6yx8d6mGSxf9Lw0FXjEkgGMNpv6SWjdn3f1yi7CxeWQsD+pto+q9TRA/oiHyK9Ll
Va1kv0iGjd+uLaGGmCp7iUOT2BbAbMNQ+u2dCsXEwvKjBg7lgndCfUZ0/rbq3BFs
sCY/pTEeC25hIaslSLk4ZbqFPuxM2LYph0Yv9e1+TzLfarU849AOX0CLUAxHotzE
pkujiGMfCKlsbKtZcu+xWxURvkhylSmi4Yot/hRc1IPRoRaDCf7KyHdIZpMbWrXl
tDiUOgxh+1ehdrXAKgyLH/evx/hwtqiSyVH3ZEwvYOStzOpELEfEOZFDeQq7bAKg
dHbNk0qLDL++Te7o2b+qNJtvfAbLbFO4PAmJFIyzdRAQsFJwWTyl5CvcFSVUoqBH
NUNSp6IzP5d75i4zdDOAly9TyNEdSyeTQpFasnXi9pdqKevvT4YPOCYWpWNagqZU
lumm+vjmbtzhplWTFNuwGQOlW/osTJ2Spjb2bp6nAY1wFJR/SH5MlzFaJpFa8z3C
hdH/1xyoYTU8QLu1kgSpHnC2CXtzJQVc+CuqWFjR8/jhRS/W1Lc5Aib9ETrZe1VY
nZLiuPb5l/g39mZ0cMJNtZcBvIzef3YvFBfajNNplbyTfAZw8Kw4I+7t3/1QIWlQ
c4VfdOz8U5p+exwEPRZM37K2oobwnfnRRNyY3xJVNpVOdJeZ41As/MI1p+P3fIBS
WC3XnGQz04VxB7fg76SLBbTiah09rSdF0bkNeeBf/AWxQ4NdIxAap3vYGMFHtJU0
DRriYfLhx3/ON3SYOsaZJxA8p0z/pNE/SmqfN6S+B6iLQ+rRAfr+9Os01F98cdBq
LKAuvIwCwJpA7HzWPk9EQvEDSNHns0jDPOe2h5zx/GNuBGD5QxtVs0yVYw/Sm9mF
ZGzm82qF68kic23EbjKlbPF3Hjb6FcYJdP2ga7+RYAHrZzkq2saY0bnFDgf85Af8
SEE1y9hB+p8S1lrE8w+ltz2ommGf+74XnRT2Q7Bwzi1NF02gqmTGoNiejDkVCoEC
66j6WJvtv6qtwcW00sVgmFbY+ig04kg6v2vEBGspKHB8bTo0UgxXa2lKsI4O08yG
NxGHiQ+D9Bs8Vn0X+lkIDRpq4BBTrRpAJIKaKYcmXMJY1mzLQZfgc9NpJEj0Aa0i
6TBcImwwaNrNJ4PyEo9yAw5GezTY+BCvrr1jkqkU9JHGlyaHW14UrZ2xO3OXVkXd
w5HodJCcmq5A/5Vg4xl/1ogx3MZINAvWrhCKke1ysmkc8p3Jux023aMtt1KTGUZS
yOjkm3G5rWHK8YyTocCCuMdM/8neCHKdP97chpTBaMpFfwq85HlsPzjK8ytmao+c
lA9xq6Sit4N4UdJdfUTdn0sHvIE5WHNOG5CBhqReevg+OXYgW1n4ozJGyH2X8SvI
m6CyGg9kNUWIZ+U1TaY6V2oaoxXCmTCxVmQ4HeOvCSdOz/Gg3sZSfpk2pkAeyrK7
w3xMmeCgTKX5BiIL8G0P79a1BqF21KwxeLozepa4TxNN8qrvXZ3H0n5MXpb2eK+n
jVM3m/qdNHpQslo8S1gkCIRilgtU7rQzFK/96wERUuWV4ki/jXRymufXc+66LlHn
AMdotBXIWCzVsyRBcmA9cTO1F6UmrUAeeM7+eN/6oUUJQAUKPmw4FFLyI1sB9ruF
C48ebmwnePvDbLQmTZSlwNVqT0uWc9ZnFIRECOhj9YbOtuzMkYjuVTFLcTalIVpb
XA4PIPYM1HEFEcGj0DjKAKaDcXsM8eU4em8Ssw9LxDlE1TE6nzZIXlnXK3i2nFr8
t+tmuAjwoQ84dNMZu2KP0e5jm0ADMos+93CuMWfu1VrCXkSUuLOKdt9TaLhM14OC
Sk2PrRD4NnAYXBBxAXp/fD88ySueyQhzoYVHoZhyp0Dh0j4DWJx21/OSij+xFPho
PTLfRznQ8QFAGUAHPkW4QguTYT2NRMnTca97B+QU5pLvKyLMlrmaW2ESnf76QxMK
Cd9YxxOVeERyoQpNMcg92iyrM5OuyCyGkisVKnxViucRGgUWvv5JpVKTYEzaU/jY
EJcN38G6fZsaDkJeYXgXzJ9hYM7PISQAf/kcegM8x1t5OjEkENZIe8TX2YXS9PRf
kPZhWFLrdDF+IcTlfGx3M6aUfrErNRgyljVJgfusJg7w0BtojhVOyhz0kfb4MXok
DZwWKI+jDS3Vf8+izzn1ydbIhzVL8eN2g808h/HgQYdQvSYt6psuVteCEkJjASXg
8TnM6hWdnkGhEITdSjhkOkzRn+Dq/ZCHWN/GJF7hY0/xvbPgqeAZNDtz2ubuTb+P
Bl1WDjl8FadCoY7ewgpM8lNNPNwTZhIOSq4ZMYACaqoNXwlXTU6Q+xXc0TnMiH+N
RVpFWfLcSrzEcgZ9FE3MUSX5qlFpM/K7TR2ceBKlUYcfO48++1nZCoStkHqLnItJ
m9OtUvhQbUCe0iqn87FrePnCKZbtNAP5DPS/B1ZnJ5fUYi8QYBMnRNzfnzODbsXX
rxDL4bHW+rmjup8aBgQCoQQDAidhqzt2EgIvAw2E7Op/CY+UbSZ4EZuDDCdu8TKX
LLpXnmdgWOjBIBg8ubPnywzcsZzeuEnyK5ZX1IOc97JuGD2TMFB3GgW3weRlioDE
cuu+3fuW7w/8JxzFhohn0jwmnGwYmYfoXrACyDiSpqYqENAGCUAmJLE2BSpO2neK
p8OoBjePjM4mMJPIOcSL+w0yZG1GbM3pIKmRm/drFGjEoQx0kdwFrWDv10CoJGan
oM8k/Ua8dGuolFT9WWMwFA/MnbYGq36lm2Q0tAUOzh+DztTBAxpH/LItBCfHp4kP
GFLdcoJXxVd5VA83WIcxRlJYtMQQIRjDlgcKfoEzZhNnxvVSiqYV9UiCjW4oR7Y4
CuQ9RFiM4WojuzAXtvNchpKYsIf73KDlft0wEeKdpvG/5nMjMjB6FRUBI9GHGdEi
3hNFlG6wgd0HgC7C5YG0bMU7FiKZ82qiFNPGPi1iJkfDsEkpxxpDehcaoHMddxIk
l+A8r2S4B/NddAV3FQDecDwcHTl2HHgq0Yvgq8EeBFixJvW3275e3Lq3KmG/LwYd
mrH9JYq+39UExZJX00+GT6WWSNTHitc6DXZPjpUM50Mioy9wR/OB23fMvCenYdjH
E879v1shLaNjyahywIuZIASaFn98XEvSBHiBifYSum35jPbOgqgkc9FMIh1En1F+
ROfpcQVBCxevLnYs5K8ecConKYoBeavcDmfqFx3bLQkhuLfmzh1w2PfHu7I/7Pbh
v4tV/tEZ3wwFT4fDlGWXQHHW1AZldNquFj+d+UeHPZHV2DmCy10UctPVztqeQWiv
/Fu+vJfIFLP4gjpVvep9QixrToYWlISz7SbzuLBrJ3UJNF2s3VkGTCzbj130r2/6
zmXH9tjY8pPPveEAEvHC/Bu/AZGD+ifbMMkgwMMb2PM1w0XgOEbSE1jcf93PZLQm
u9DqDTB+2t4ktsrlGr5SFN5KqpjH3QYb/z3qVHpia1V/KFOHKXakIqkdVRiuK7U9
Jvxd4tcfOkK25hQ2jT/zGV0xYEi2ZzOsfLKe6IedFRFi8B6kVaum7Ga7xGIy0fFL
tP47CnmA0J12ofw/F7Ek4H3M42PdwM27GqQsxBNJzByDlol/S5AoAli1qBNsrqk6
icUsD6Dq54n3CgAObT0tSaqFnO7r0YXmuJJ9xC4nmG1yyCkEQl/rt61gH0vmLJlr
C5Blef38qGAPGByLqcrLhSR1QR4+XkmQE49GztUDmyJvAHhLK3km1Qc7RZkW6QLa
8zYvDFBGZSk6k0CNXsfssbGcmo/Qntiec16frWvRj2rTKZ6c840LMg3N+O0TcDgS
pAcowWTz+h0QoM/Q/klzwoe9ZEkT51ur2ScgNWBKvs293SYsrnMsFlpN/zPKB17u
pKrElH/W32qNFuGMG/ZaudrjN/Aeaw6fIFVk1SEgiDTvfkaL/WDXTSpdPQ6a+X6h
r9DENUwT8YglGBYytKOxAZWnJPlyJwtC+fGQBDJqpfSkbZyRNDDTYklH97t7uT+c
79O7ZSCi0FBeriQyYTBt74OizMDIdHAoZy3p0FEdZa/pTKiYCm5cXa8+SvC9NIak
3+P9XDdBveNOfjv2+x4GB505KhblOFf3F6D4me0lcwoZc9aW/+8fxnzZqM9oKG1W
jrDnjf7BjwQCRy5xRhgr3PsJyw+bzzoMbGhx5M3ASjRf+rQ6c1IqilybulNZrd+I
/+9sWiUSoQvhZyyG83lUw41nM1oioHVo7yVBSe2p0Fh4AUFNJgoLS58L0uhzWeU1
mQ7wS7ATfGjmRCOrQgz0VCqnM52CpSMV0xiYi3+RT4atXZwTctMgm9Q6gPhGmIeT
NCPCdzuBRgkb5QNY+krOus0B4FuaUNTlnNEHRO1ZDQDevcy3o416qs2ShUmIK9+3
IVykj3bLJBPC/BSrHxHu6oWart+90qZO2yR8lwni2kghu1gkJeUytLIvyODr5/ZN
vAhMaxWu5OjtxS8SaO4uqiaWiUcibJMflaHGWGayOMj2QdUyqNMEfQ6/31v8roe5
6l6pextxf6rY+GPvK9w4yoZZVYcvUBvsU+lBUOIFl1KRRjwM045uezJKq6e5KV+Q
VIt2EcUByvPvkmt0Ji0li/LIxjuojCTUE/qNMalmzvm/HMIcBYzv/a/Ux/2PYnB9
BR9JZYVhihluhjMDOVNKzOL7iusxCR0TSeyUvAqP94c9WD2x3O6sk97PoybhAaMp
vEMSrTAsnAPuYNwKSZ6Q3GZbmHURdbSYfKG0iVrBfG4kCD063NrXPTUXd7kBnOos
aMj+nuKTfzHKSJPrJFcjT1x8FWY2D8ynhpPs/7Wozn/hZZn1UU0b+JhBVVj/c7FZ
B+GjmHcfdVmZCiXtcJz709Sad28KKfQ0pyHKhhO6B2nuUYchEzemf/alzHgRp9by
ER5uMP2if28yyau1fgA1N1XG9eHAHG1e6rySAFZ4fcLtw7V03zLJ8leB90WSz/Vv
qprQva4KD0NrD61AwNZXFVVh9NLHz1gvD5h4omweA35VAa/acn/4xOcp4cClqJG/
16rBgFO4QsMz2RdpxnaZ9v6cX9GrcauGKDsYlwnYoNrEFRS2grBrFnnHlIusZ8cy
skv3ksIa2IooApo7pliqTUhBdFdaBBvYHUd4EnDFvUAiJP/iL/ISftgAIK9iQeme
Dxl9Vn9iPloS5PaHxPjYRyekrVKXHc/PflzMoZMKPt4e1acRHzr1jNTOqlQzXbIo
Gsl1/Z/U3z4d5fcFhHzelpJU5msWCXf8MnICDgQws+8zcYFUhBFkuFvovyrHUVDZ
QTh2YGsKw0KpbqFuagTRE0qQIP1pBqDqjNKGxTCPXfeUusPf550Mu+gh+Zi372x2
UsxAQ9+VKKH/dFlJKMcOo5bJLgK456CaDmIWCgPpeOL0PWDdSvZwYLSq9Q7INT7N
7teNLuEvOrPA1FPD3jyNJ+9SPnKlp1eqpJhMi5d29QX2lIvP9wgVO6RJFjAD8tBf
v65guDLKaDYsMrnQti5XVC7CFngmpJF9oZxxwoF7wWxFXPSAFt+8axaEdbJb4TOp
uh/M2FcBIMbBrUZdQClwwGxKWl0LZ4iHCmf3H6pRnq3HxRdKCuowt2onlwUdYDI0
edfwV75esasconbLsalHTbYSdXUoOIH68a44QUzKm9rMUJlrKBweeG/0RIv/6h4l
9KiI6gbzN+We/TvuxOf6/mxMPbLpHBmDiRyl9UkKiUHFuNZVuDjL8yU2eWOL0+FR
YGNaCp1rWLgTuQzG8TmPEkbnVeld/EoHbMyMpd329NRh1OJEBQwdz2udrvjzsOG1
Ljfgmm3H6/qhy5LmcMO47y2i+wepWcfrij+Es+PS3OcbEfwW9oVfZdEVvWViKP6Z
t1J5Fs3oMHwq/lmhbesxusNDOYH5aEWRTzoDoXGtDOtJiQEckPsLhL1HuO34ZcbT
f3uSfs34oVW5a5QdfqtwANdUGw/r10uKGcXNO2ZeWNZnzLPLhVJBlBoznebL8imY
J+YIBEekFGuDXfwLLqhc04AssQlkKtF4JTdOR7OT2e7bnJdGZHucLc7Kzdq1/Qzo
EG5kT+xbNAK5gwGSUorQp6mVYL4Wyuy00T+ZWjK8IX2EG4NI5SCI+j15H3zdbYdn
LbySORTdo/ctGCot7K9IBAxMFBEQk/JJfT8+P3OShdWBwoRtru4iwPOKG8K0Hx5/
sPnkqFX+8xUKVGDhafVG/Qg5s8dlmsnYO3PXQjBJDDKRt9deRyMDmupjqz7X1gmK
48ys9r1vv9eADiJo0SFdCwvA8rIZOZ8eAXDk+l3ZH9n0nuwZXAyw6IGxvP//A10U
SNh4/95WRPosGT53v5qyDQKVJC1PkpMJaxdHJV386SMc1rO6k6Uzw9dN79T71q5S
cl+MbDxB1mzHpXvoEokQtrcfrFuLOFX17hfvxwHjeB6197wHEBDrDQikhhgBsZsj
nVeDKKJ7PvMj9JZK4y6YDw+yd+2yJvZCusRRfR3XLwN5DYEqjdvKI3n+ePmEK+rK
EFACKhhm8lz0cOChb7FVQ8pqGaIgsDrxpA8hTFyNo8c/vxwXyuGhEIMaqzh4JWm5
OgV8Usyhy3lJ1/7VxXh0MpESiq1VlL1WUSOwmnD5BWkGgnq+G7zPS+v5ewMbITjo
/1rkDcsJ19ALpaje4EtyGvQgaU03bKGxsVvGbiV5Wd5TXe9o3ubkDVEbs5X3X9fa
oVOWK1af/pF6Qp+c8EmK8UgML8nG6xULSX/umHtinmJFa4o+iq5/rbAfkmuloS9a
vSMk1Sq18tttcs+4wMWMKsnNsAGT+IRuDSV1r7jn8Jfi8MGPaUKSdNvaAez1+JSj
inicGXyD2X7KycBmpDVBKJUZt00cAu5xdTEsQ4k4qkHocFaT+BLT/sBbrteeS2On
JsqgbrbKqi5iBkYfOgljiX1ilxrsITj87wXUbiwulejHWhixOYMVnQu6n4XJbx/x
XWulZmeyPOqt3OymrTKjIoEhB5m4xw8UbDmnLEJGdS+KXsevqEwglXNCKEoIguDT
99tS1oGTqDwXiRGQqWuRs53vFgq4VU88b2+ijUwpkLC9JxbwmqgL2C1gDA0i7rfA
vzoZ4LT8twyNB2XYeAywl8iG2fzoZJmAiu2hXEpgU+p8EkaMa0xCgl2EpI6seEdN
+B1oJKmxLpGtwBShkcJtcowftv5Dz/gfCGGlUuTvl9GwxVmjXsdgKG85nYgTzcgY
J5ZuSNzdWO/W9zvUfjGBsx68nVwMkB34aKgtaTTRmtwpPutmVIcrpsbZBgyigxkc
4m/lPt6nu/7wOsyvap4t+BFZiWYxtVmjlkmbLqDEcJABnBIbSnzj/06JmAT/hbQl
RhBHBzgS6oaEkSB/OfaIlQobcEM4AFEB45vLikXPXD8B/C9iOOU1+PU/YyesP7jU
53ESZVfCJr87+Sb3SRVhXkM3iFsbiglyxUh3zRT5oHaURXDJEtwjNq45otxu+yeK
TTCdbELlfTrWY2kK+Wns8RzqwjJgSoLOH0UPMaWmfIXHGzY2XD0fZVFxxJjQIvlp
I5vDXYi8APhrGAv+PI/PH0eN9hosQ87E0EKxCsCbr/vZr3VHVJioHw+4dwTyjeLG
2Ug63mg5RLU31aCSVv2JN4UXuQwLINc0OVDVg+qTIPZSr9GIaJ6tmXD7IPCITUHl
eDa6Y9ORS37R6719NKqd/IAixn6dGA65e7kHAXc3/3h1E+1X/2yiO4SBJkmFJnLk
EwwGx+zVjVSs5oJHsYTO0aZ65Ldrh/8/DKnF7joM+iPqzY84abqjk631OTHLIGyH
HpumPN2ubIoetzDZ5PUqKVfmP8p8mdy+f/T+m28PhAgJTwFkujW0cJtC/OCKSs79
8DuJpJ0uBA0s5gykiP07AqSrB5A1jyB84uqkcxRyEHA7DQqdp1V0vEVdgMW1qfnN
ko60CtFMk+Q+YVnYuKdDPCaIvwfYHT8Ze4O0eQACTzSrx5cZOagl1YPObHD0r+xr
WM6VpVrpec49rDlsGPnTNCS98nE1m+xdcTMhAwVMRPXVKlaLsnzMyzJF8Jul1XPu
/s4ByNCM6A0itFVNG5YfnEDUIN6bIxSObp4NYd14j+eApMFAxut42IH4QWr7cedA
wF8/mwfWvUq/IhyIx0nDgGo6RBSOKuAVW2aWhUr4tFVPbzQWAgJY8yYRnq2Dpppv
p/Ih/S7CP4zJugMDaSf7viAcP/frhWCJWJR8gkY1j0x+B6ApbtAYAFXzoX/vCHKi
KKgH9HjCnqXBFn6HndKZ8mAf9zCmfEonSGfMqCsrcPa3K48C/1Toogi7sd4jZhAJ
URaCCp+Zr+jgI/Z9qeDEPXJxq5RpEyHGfx8FolEvD8g9K9XiOJDPkHW+n8RUdahX
4A5eqiEq3QHbWrs9/x9fRY/TYktopCfh1ATb0IyQmstIc5Vg34Urd6NtiN68LOUV
ej+6162Ar5VvFLMk8jwEuuup2b6I8p3ahIz+qauIp66d0D/VoO0PYmLF68HAXT0q
wkOQfE6VC0OajAoTm4lLWgryiDm94jgZwq5c1oMeKYmMi7uFPNYdTNT1eaL5eHnX
f/viclrTUtlNXeUu+eziwDJb62iTvVjmbZPe2lpiXc2Mez3p0zMW92VFACG4AHON
3tQ3CiW/spr63tZUNeFfzbAZinOckQvT9DlQ7GjuoskHaUImjK2UzVUMSPHXmQFJ
96TppUixEUvtGM4rh1kQ0MRGHQsAASGtXkjpP8lJ/yt2/K5WLxT5tXxm+lsqspBR
Obdv77nmUDmSBFs/SgpJETQPBssGV6beUDveaBft+AX6shsHzfLFefjACHTbwu2l
HVRxiXs66JCHG2fy5R69Fd0v+LUq+JIl1vwRLwsRLAPbyXnGiRuPl1F6xVRYsbJd
tN80PDOK+5mVaF1fEEjWd4jAE6SFokgdqNvaCWM9H58dzJJrW/Qg4/a8hGEvqGdT
xiB37jbR4yGDEc0llL/96aUAzbyAseRP8F8efX3p1J8dXhdpe3OgaDZVNEtodGwa
BPWwTDVdl2NMlQu9oZorawbnMpCt+c24Q/y5it77ol22Rf3Rrg7wPBYjjNS938xK
f+snOfTmsvAPjwX8vZZ41d+x4DtvXubnq3GIykhF01NFMVcrO/M3sP2aEXs1ew8L
SrrbBJap9g0KBB4Zwtv/HycfiqpmzcLpCbhU5Xkpuvib3s0Ep9sk10Dkl9HN56yx
awVdDeB3hxKtU01a+X9IK06qwKGO8TGC3SgcvDcETjP3auKA4zG9LGFwHjYdYzea
K/wpf+wNAwOY7fA9Ubfi8PcN6pV9Qiea2a1UaoxiGGmYDsT/KsrkKiCyuYizuGxr
vD1fsnMMD1ZhmjV5w7cjN5U5eVEcMRu+YGEQHF0z/WAepqjooIxaolKaZWtZb4bR
dlQRX+BfLysud4bzjt4Dnrtt9VR+lC3OnrqMObwpewDBg8VBeC6Ye3Ujd4Y0dD4y
Nl79STBlq8zb/eSzBvJesh538Csn6j5zmWhx59wu4C0IgS0Q2puRWaxlGqO6ffkA
QR1h7gW+pPeR1u4FsFZmw1ducv8NxVRsBYsPe13IFRaPZhcsHhtd33d3dJf9RqNx
vOMzVOy6In17hNkH73lWrQvcnT+kDWKcEaZPl0okzL1R1/HVXXK+WoutMfet4oNV
w+7YlQ4hATbTOk9XRXpagRsASoqid6hUwoi8HfYiIlkbp8++3V+A8OTJtcfEalDf
g/7k2ZPiB9RYcgfQAVbXmuxP/082B9wtHy+ZhiWwsSD08+dKsMNtPJSHJ/RVY533
oChM+9jA2rRXcczlqIuoQS6dmP46LOfm1XLg/v3dOqYtgqJU+vB87IZ4QnbC8KG+
vLWB7040a9dVWPHveRM2nu3bd35dkYfKSi5dC5075ZqbJC9MHtuqyTYpiS2+2CHw
wa0yNgvna4Ohjkr7kOwAOvTLzDIJerIim+dXDktTkQokPBSI4YuZT3l2RkdlUOxm
UmJ4ZVkZ+Ie98zCO/edbetX9aSjLK9e/6QttyfCGw1lgyskDWDUVy/f/4/noBQQk
GxgcYX7QXuHqEQFDH3kxzm129I9mq52hylqaY+mT11j1fK0AOt20LHPkaM9mHFkS
UnSG13ROUTQq83p3QI6Z/n9/51hdFQYjmNblLU8bl3L2yIplfDgaAQo28rqnih2j
KomAlWa4i0W0YgyXkOEW9pUSNbVIKd0EeSeGLedEn7OXlP/itQ18LcSul40R0p36
ztstduuBZ9CtiVWmMYiSJzfqEDssoBfmOHFa2/RSSB6wms9rWN0M5UCiu93X7yp2
Z0OmA+Pm371zFQp+UWzImRjs3I98b8fPEytJD5ds5m6wlcpO+EUKNwrlRkw7/bqD
S9LduF3RksWqipOrf+g/a459tTVyblAi32LdFta9R3B0ZbUrPvgR4dS7Fbvj0+2H
m161IMT0xC9xMWs8lKDRkwHdDXxGjJL5YxzdHB5PuqOoRte9gQiijKgm791s+yKS
Xg2aE77iqzwnwXO/itsWTY10meonciG9mXtZ0LEjXXivCdnsezRoOnmJJUk+RCYS
v7uZNBDLf+xJe2AkeyKluGdUUPtDJ9OYUVYXhMXCGraGIQklmcKKILO7OuMyqhHo
Gahhwnq5IUbFmVUOCRICqNI7N+Qe9fTmnLy74/Fy/A4UR9Cj5HUAuA5akhPJhtY5
fu9VU085IJKf39+dseUDsa5Yyig1ATl+ZjnNOokvo6eUqyaIq8alfkyrGdpbhLUG
7x3uQR4egX3YQATwFPNMPi9gL8gqXT4N7CDINyh4YzVEWQ+qCo57hRvKKfH/GY3U
UFKodEqt26WnGwNb4hcDSSDwARoF9V9vOeGD3ostUUIuY1809hhnXebbBzNx2FTy
tHF/uTzWW2zc5XnqlY900zqmh7ihe0o88+aao4Ao7ZFBfeLvMtmbfUdlqOek59WX
08iUSJ5sJ9IYPcCInVoy0tn44XudWcU7lt9nr9cpLrMN8aTyNIFBxHhV05Lzfhve
ejGjhLiBGfoZ40V+Dy0f6CK/Wvs8PSsbq3X/5rFBXD/kPSKyXPl2aocMhZmKEzzl
xbN79suGwGZmmiTFqIh3EeMYvHDFG9bonvI8UeUCk6Zhc47qS8mGyWdCvw0WnK+y
cnmY2MSlrMLKi2h+jcQMM7FSc+lhIU2LmCx0gHpohbfFeGuboqp+1x30QEGCWr4P
0AxqZG02gCJcZuCSgzEJRp+M/Q+rNWDf3+gxHNuMaj88aiSCJqvTN3lyAk4hv28t
tN7VvZhsU2yZv+VAPxMIw6P6NsAJFu3GX78NoHHL8e0Fh1qagNwKVL3+lw/NaAaP
ooyWR9rHrpLJDTCRdyzy68DqDMphcOF5JaJXdsj9cw3aWL0lDgq5Mtidkh5l29wV
/3iqptGPv5oy5OY0Y7/+WugXTGfq0Uaft+rDVWpfhlPvri1Xt8KN9bKU4lqIU9D3
31vEcPOJSn6lR3E5U3LPNSIoRAlkQdkFOZXZEcIVIZYFe00F5NPdFZ+x9+8Gg3DB
mhXKXLPJO6g0USux/SzPY2OHHZKSlIGCk1hKTz44dt01ZmcW6DLrTubDjAxSiFiE
Jvt9xa6qE0HbicHnePdp37Dk4dFeO0EGUORcLdcaVd3tsCehqJP8IM6M9ktzJtqY
QvClyDh9D6TfcoyPhcjGiJ/x8BT+hGco1/pPpPZCuEGT9RJs7BXP3F+GxMdfZWYR
gEXcES+0UChijNxRSClhysHFS9SDueCuHassTLCr/bpTNJRlYqg00nAhHAW1XuGe
q15xTI6v+mLCqS2ad3YHolAkR2hqL7UshPSiTKMqbODdY0wmRzKp+h9KSHRoSiWu
p6i0FFKVdeA9xujo+OJtwjHqSO34Wkf/5xejAMoC5jmdwjvQe0IkFV5JosFVmY/Y
sPAI/eckZVwNz4iv9P3TvlGdfbSOj1HnRnYv4un6trx6SxFZSXHvO1AV8QVgzQgD
91S48LGceczC2q1PEnjsgvBA6kxvEDO7IDfKNsxjkl3WHjsK2hQdM+syAnKhGEAS
1h5+moaRkCkW6ffy0cb/0ajCUJ4uKabCg42B9qDwzi7WuCXJSOEd5YyebccgMCGD
w0qYLuZWMpTpQas+otvLv+KG0GwMcoEDLLREgijccB9FLAMYfNYHi/AdP969f3b0
3G7xdLGFehOWMoX0ATlXxDuC/G7HN8o5XFTeE60hGZVIaxjwX5lIhtiUMet5XA7D
vS7sijGQ9qWaNUVNqsA3bBOH69b75g1txDjqOlCobMglS5TJHiti4levC5YSxV1u
bRwoI9U3TCKVUVdG8/MVmy7lO6IMBxTSRFuEFUmtfAhrqStDTUJ3oherUA4IotUY
nv6F0O6fnER9i4Q7RHRw6VJ80xMt6D/KofQY87TNkcfIUJE4LqxlEftfbxtS8/NE
PHxazxkj/iRSJW5R933Ff6CQalQXNi71iO4+wpoh3uhqAyDy36t5uiAtYc5PE9I+
hTbYEWw4cMnK134+EVA4qieO/ZWrBw4uvEyyWAsoDT66A9d5FnlKb9tGE8xZnJTS
68rPt6Js9O6baZJPrtLHWCuC99RLk86SUNKU1XskM66LyX99vcd1wnzkO7YGSpgS
lICM0f3bLuPWOzCWNglKJIYqx96hv8RMqIMorhPfvoCy2XrMq7ga7PMvTIArlqwX
p6xAtLyJg+9So6iqFfsQ/xzLX+LCGFs5VlU+XGq7nWmulNRwbYQ+SmJWuiVV4jWV
izdY1r9yTX/Rq6ozfRNW/HAQKy8M6OtPphmdMtB3QS6j32dupELI2Gixdb3bDslS
NhX7obrOuEMlOoB+OvhTWeK62yQAqli2H/AqHIzQlYL8ndHppwgTN1w9pDnQJuZF
UHWrl3zG/YtTvhWlwatUmj87U31w/CPgbIQfX9x09nmEMddhDszNxDdTqBiPH+He
JebcxfcwAIpBGIhPcZ9wiJj/9UmKjNeE7jBmNcpwTFlyiv6sD59yB6sgQ6oNKjx3
DgjgefEdRNuz+aJ5KUC2A6zMWa/g7vGeTcIOO9i4KuB1etTqgNj27XO3U/rfbbJo
UYk4AckkAXdIPLBf6CbMrykDmwhklsWR/Rlsecj9vLM94bLdCG+eqIpq654CgNCs
kp57i3vJDEyVj5VPF6DsC0rZMHOMJ9tncrX/4O3MDSGz6mc1LWLiwqbKTH1HOhgG
ERgf4VhCk1xD17meQL28BiIsVRe9Goqlmct2OGa4tIXVSvjYPeDAqwsZFmYwPbYi
FALdWxYFTFDGsS1pt0KxKCervmMuq5uCnTmgJRvZvrAFX2jFrEUYo3kxhqA19l87
J3h0kr4OIfGIz2eyJjBrnvBYP9jgBOKPsblgQzvMSGwlC+8pSE04LSNXO1pg4I74
wwhiq7XHwElkSpTuf0Yov9+AZq8zVZ3BVOreJ04VQpyWFRoqDWywvoiGSFmjrFpP
9Sdoe1UY5e63epE4nZporh8H+VxZkGq+/LjsYS3vCNKWnjy9WvNm7839+aV/LNsP
Plk8tH+2NppIs4P7k6TaELkt0eObV42siVSa8wkSJirA2DVWXZf1J4Hl8LKpwbT/
AXqccQLQrCpomLu7I4QfdG3+Eb1BOpzcflFssuD5Usued0YHvp5Uurt7R6a0sGYO
Lr3QCUS3KfxCPHKnLf4Am46g+ERjL3Thhpyd95eIuJ/C5LdB/pNk/NdQMUIHLUNP
M7OaSDVX2yGgknfWBAHJ7dcuWxwiCTW6B/N4NtGEKlDm9cx27GyUJUAoj0iH1uX7
Nm/bUltvlNcbhGc42fn8FlDXkm/bwPUYly/UqKNRT1AeFxu1aAjS+s0w8U/LfpFi
Bg3PC20ikdNEpDwMY98PBoJXM6d7mHQdu2tu04WA7H9bdiuEzEwXMYPZEYK5mICO
5Fv2vr753Ljq7re9Kt2EYrlzRnNcZEAsqwTVLLCAZYLs5CHUVO7cCahCE77brLY/
mDr2c5AElgqeXj/Xa52OA12ZUqelT59IasvuMCf73ygyZEPpvTZX344NhmRt5hJx
z5u3kL+6PfseaqL14O4bgEcj+6lC4IUG6ZXAvyD/VuaSPA2DDtMBmQNGklvWjrz4
S6QFFM1w2YNwRHlO06vu0dQcezXCM7dlMn1Q0UYJW23Bu7n0exWtid34CfmBw69l
7P5hS3JYsVgFcZGlribZRvGERnUnOIu1nsscM2v2X9BS8j4dzRwaHQRtmGGG+VPp
q4TZwwEYasjpZYbkJ8P2qodc/n8YfiJCJ2ydE+2Ta9p4kvY5X5EwdBXqf11XYgj1
q1ftucB+1LwuKPGPVe6Wk3Nb0d0Z9j/ilVbtUQmH4yV2ifv/75f1cITWSCC+YFCQ
UXEbkCuAAzFargokVqNdZVdPaxusC9KjbMv60hW2LIbA6p8prnRF9I8R1ecX6bfV
lWqIEwVNOwiZgQgMsHM5STZZY0rv1cHapPXHK8okEc2NDmhcP2QddlNuvUbihIUR
9MgE/kOTglaZ+N+dy2xGxUbYk5M2cTCm2zCng1SXQB+aIVubPanMGD/zsTHAopEV
Ihe1ogVIk1JGYjcFaGn/YCY3cV36/jo2S6ayL2ZQTT+e2Ex1C5fik+c0nTmch1xM
Bqg/ItFe+53IflX4ZEIlCUE9CGSg00rF70kTE5qKMiS/rMxTMNNZ0zI/GKRlAXf+
SSu9JrRni8dISdGu8M5UUXZEkgSrjuheQKtwf+Brxq+pumzoP5NJsDXq4tOqBL6m
kbjg2WjWBmMtCF2k5AbzY+0G8Pgy2Bjm1v3L3mogU8Zh26rXDisKdESLDgP6q5lx
Q41igqV1pavKZinlSw1CJENH4Gp8146KFSPopSpJ5uLYkK09zgJ4byo/OU6aPgY4
Emog3Vqu3rvzN4Rmd0QM5y93IQivcGUEkzkg5FMo8hK9BoWvUi3PXq0ZEoH3Qmdg
OgVAfWImL9qMM3vUkFxkYvHfZDBXi2DwLe5C9JYyRK/th1pWj3Ldhxnk7HXvnmAh
Zm0Tjvp0I9wylTdwxLCEjTDKX0pqY9fG2Z3HLCxtpqjay8lHKImuRnNU7rqE0BnR
gxfW0oO37xRYGdmNhlz++vw/tI4Vph4WeHpyYPfcVvuJGuGlD5FG4nFAN0Ra3W+3
mFlCWHTg3PGqn2JS4X4aZTAcXpydJG6nbZmSChqJds8tDgaiUv8Nkg1n1tF6IrtP
xB+hNZiItMRyRbip1CzIueCaf9NZqqyXcdToi4rQyQGcR6nj2rjb+WpWgXrvTIe0
mKk0irUtJ2sVtJToCBXQqKYcthgVOZUdxynPFjZzIsBmCHjZ04H+rsIuwhEGEGXI
hSN2o7/XSG0RaHP2O0fXyU5wf8vqHBYzPWSaYqXIdRwJSHToMHFmQ0k7z7HWvrE3
xnlFw9gqK0BZwq3XRvH3BpsXmjfmgKBTMWF8Gb2M9nOiQreE0M/HHOIMd+W6R431
EZUbjajCVN9+OqZb11OYUzDIv8vGsko1JELL9UC9PdRdjRtFgJ9DZMVhUJHFWifP
/cXyxZRhRfRa+CXROeNRHNZ+DdTn+YOEtUD7MNfxV4ImVS8jpiCrBtauV/Hpw9G/
e6/r7TgCxhtnpnygdfaArKZl+PaJSOuKZ5rNkK9AaxFN0Xh5qU3MNzb72zDXffML
57CPluSC4U2BaW9sFV7rADHPDPq+zQnRPY35pIsiTDvVWxS+NYBShr4NXfiVf/m9
WyxcyB/mKVta7MSmAJPmEE+haTus4liqf3k7szTZ35c/x+rsD41Rb2lzKOKFuaB6
7DSjzggZCe563hVOKVHMNSxvS4CRLEPhxSTk3zRc0HB7JJg9jvKWGCmr6L0cPIYO
8nFKsfrgsDfdV5lb/Ebx9EEI9XFfe3lqlS/hQZ63tbcZyIzwO2TgFkM5x3Mc1Oxc
GJlZyI3338guffc1YG7K82lMFOq+qauWYdUN1i+VPHuAeLHnMNYVO/2mJseKSk+V
JcjU12OYlwtk3fF3eG/mLXeZWjxYZY4AFk7NzUNJk578wh8JO27J5e6on+BXK9Zc
i0NaUiTB8MP1EVXzklusbrAeFI3jXfPzZeXx3pp1iSBs/ZkNZrNkEvMAsSoMDD8V
jdSLvGHcxvqXCsmfnRMOxWmhYleitbz348p3HDUoIj7U44ye7FW24jSaiOE3Ifz+
BffyTiju61xMD3yZQX5euynqkugAr+NKOJqwcJTL1h63/ppXfi1+bpNgYkWBpmpG
nvJCXooWQTxwnICfMGWO+4JBkV4/ZUuFMPT8rhHc8gJ+96DONgl/x5KKCXWle0d2
w6m1VCareV6TnfqJbWX0Ke0u9jORvZPnXfgGNds7uzXF93arkF674ZdkGBxANVce
Ea8CmTCTFEHnn2ZBMV70I1RYOSbHDQo64YsoqnTioWUs/miZDxTZ9ey0bM5cpxtV
QOb3Ix5Pz5QmfiRAKWd3H8DCii8VRcCmApvKkUkBjCJaZsMyCawAXor/A/5Fqwbc
Q0eJ6FG7m+VL5N9iYNicRQSFyENfwLdTgn3DW8WRj0dfnFNWOGQDxxmH9qPzt5rQ
FpMnclAIrcetJ2oA2dNDql/27UtDI8k72/w4Ivz8FP3MYvGSbEt7ONh7faXQH8jw
lOSw0vHUOAKK3XNVf05H3QdbOFGJbdn1CK37AWfiFXr3LYzpt9eLmj+8438Q2P0g
EV7rsc8yG/xAI5jeJfQWPwYgVsk6dqUrPZF6aPIpoVFPiaFQzP9OOTm1/1gmzBWn
mo1oiQFNjMNRsoMygup3XJ3moq77A1nMoEvJgknX2fzqvKXb+sYjYJ0ZDDcLhneD
R1zE8zGpS5g3if9M+34oaGG1T5C3y2QO4HZnyr8w01rpa9CmX2bONtAaq3d5v/RQ
yHR5EOHYfMa2WoqKkd++Tz3P2c5D/q++aPUZw+t38ky5RtUZ2hniE5ub0MbKvRYv
Qv3C2MPKy30HXoEGrFuzXFUElPX/S5/uuydsBIpfwt25yoBu8XiuDDc/ny7mHu+C
tVExLkMbVqu2UgY4/SmGtKVoyQqirrrORJQNwZfyyEnGFOAADNsSvnrv2EmPk3ji
wPaZ+aqe8NSH12cBRyXMMtY2aV6pH2HxrAzJL0o8ko//NLB2jpiPvifysEJCZrz7
efmIWC4l1tvsMCvqiV7do7p+GxjCHVhNaTtX769foy27HxLfUr4TF+NdaviCelj2
lbqcJ2E8eLvi2Fi2FOuT0tnpe6LcJodlGdcf69LL03XwybsqMi2Gr+GOAMIjwiWO
HvmKxMNuTk/h+iOgZb92z19TJFP1CCXXh9nhW6yO94dsGmapOxRabL+PSAh647Ud
DF4bEZ9Jz+rziibcvj9nCnPhjc/6wXHjmL8GSh8jHzGOYN2HTTSvkhDfj+aP+fMG
nrbRVELW9Niz2vSLbyoQGJbkaQpToS6dnPVaCUMkNjOErTFqd9eWurGtcQ82axft
nDpw1e8r0IY0yp9GNodnO66Oviu0s/BHmvwB4w4hBzFfLDsipffe/6bd9kMAv1NK
e9rczz4Sza1vZasFd5P9gojby5jncJFI53iEhaDCWqTr2EGUIUw7cHKMlSkmL9A2
QbX7bAc8k06gvB9ZuI8tFmjs/WCf4vPmDZnBtDMkxIvPmhIwkWyIGyEQLlG668LE
1n+l9xxI7ZRNyjxqfMVtPb1y7M7gtK1fu7lvtB0HUZgk1Jeioj0Do+oZraICuYEF
6McJ1JY1RUCP66pC7yAsMeuLU6VhZKRguAFuYzosUxe7vJK+LYhZn+319x2jkwR8
S4ugFq6Da3I5/DLLr4MvWwloeV0xUfrTtkIf3iEF/pqNMj8fmx9eFmWiAWR3KSF7
cy/ZW5csTE+zjYIIStqmpi+HbBF92BKMtYiS8SGNQKzsMkzr1WQjNcXY3F9vdn7z
PQ0gxqzvFHFE0+eYNCMcvluciswNy8Ao4oqm3H1KMNQUUD5/ArUabocGvzwrz78G
YD9mHRl+10iDD34NKi14T6aPk+oiAQ5F9cXU9+vBpyuTtdbKXwFF7tE7d7t0Dk3t
t1ktOCcXjlBYwcoX+ngzWF75h4MI7poU41OUzL3HnvNV4c8vO2FMMXJyHVjVMwMH
XSzsvhU0M2V/cU3BM6SYmfLMOb4mmQbB0alYWVy6MmYWAGbS9xJ8R84laDvkj6j5
8Bgdeq3rt/fnqSr8w4pDKzBIQMXLHqX3gtXr2Ari+YjwNA+wYORPECyCyFE2d3vg
0M9NpY8Uhyekbus3/nHvrP8v0y1TUm3096kVsn//2EelcxQchYB9v/OpzuhGOZpr
K0fVbgf4EbdrM78Us4NCYPeCEEpN+5q02yULM2CJQSXWC2csTclPbAU6MFUTdDWM
pwxa5p4Lc9RSSnbd9vWVWRGxVq7ureyHV5D5QTJUY3uY7V3A60Xsz55WmsgnP364
rcL6JJdTdx3pIXkW3QeSDP4y0hdMXo6McqOovmgEregvDiALHA8DZDr+pdPmaIIA
JO3KCSmdgYQcGqNdOlLgeSr8CRvgtRaQkcoi3rNFaBZTihBiJPDBSWfZJlMRvYG6
coOPLhNu5YH5SoarjDaEVXpqeQTd62nwgApHWitLU3SFsGhKx8YsJ7eILva1iEeA
BHoL5cHCDRlJ9qVw2sRVTFNO6dV6/xXvURHINmet2AtFtqIg5i+tTI0lrbxwGeXG
ap3MSyzrp2a1102EKEGS/eUE6W6KUekYnuGjguwdaySAXVh3wfCpu99MAdQUDBOC
hY+ddAPloEA4l+ZspqeoYw0xjhtn8efWMaNNcbvPOGFd91KPWBL5BVgZkDuLYZ60
LwYCcNIDfiY+ogB79kz6ahunK2NOLZqq4bCDlEBDFz25JJj3C6SkxYccFoAEXopa
W5Mnv3BXGyXd2Aa8KNy7CJS4WlyxOE6vepWRQOX0Fu4lNQY939r4Hr8JOFI0KZVZ
H50dbixMqOgNj+pULx0CiJn5VL4aRvglJOS9J3EtUYvDcpB/lFzAsagXTbvi3X66
zi2mlTUc6vwA8/ELiMHAHmOzsI+MZ/E4VfCSzTWDcFPI7+biMsP5dKPbveffI1Af
fU0yv2iIp4uZD6+XZXWCKvv/EKnzXluu/uVq5TL5tDvojjaVA7QLD6KLCe6+fi6q
KglFkH3E9CdbdrDi2uOLJ3V+hAt+7O2KaqP2F1w6ADq1qjV2RBf451pVpdnEGVEY
GMJgpcNYdA9i069QVEh6UDk4y1rKwvd9ARP2RqOgOBOnI4msXxaz2g9EO+5YsqPh
RfxnGo/0G5vB3nnBQZKHtz2yu0cMdjkT6ftc561ljAghrzyNs4empqqLacxjwa7k
cbqv9+vVHnU90CfmQK/w3ijvppZZqgDa8e0tb1TmeiDNlJvvqrXoBResS7rJxJfn
sEf4hlm1xfpYxiA4n1zH9IcWSqe7OMaHnULrv8ZyQ6BWtGH4w1WXIov5RUKmHADm
/5Iy/qgOFCX6tMO8ZcEJCpAK86iQWUTf4zEmmomOp3rmNeyKgvMjOGCyulI5wL9n
uJKjn7X+6HB0FdKP6JYz7OFBLlo0YMhtI893U1snuzDae84EQeqW0fl4rtZhj98i
xB3DbDwGBZgR/7VZn9TFu/4dEIADSRoDI5HQJCm+7QVVZWI56altHMFRzHxR0lqH
yCzonVN9PTScz5ksdzgp+waS18hE7JHsDIkqGbg0OfE+GbqslEve6vbg4WiEDyV6
Yyv2kQucLZZNFphzqIgow8U/EMNSubetXKmSyA5JKtGS4OZ8DVGG4j5oU7FsS9W0
mMhw5GSqSpwBxp72QM2DiLVuNoA4ifuaB0hzxPK4dGeY29mh4QtlkLHsf/Gsoh9P
/Czc73c7V7Q0uQ9XDNvQrrLZONJv+prTuYN5R/IGTniNBW31MEo7+3NAJRluCf9Y
5wIYQmROAoBax09CGRjeQF6Hcgd5qNKnilUQFh6tEDXI1XeiZohOCzu8N0iDvLBS
rZeCj8ECO2efInVO0+6JR5QDGT3I9bLBuh51dGmstnRF/683OuMfQn4CMmN5Zbr1
HoMqGvzW4sMguyxvO0KH4wRv5AXg9nzf7DitUSbZt0oSfos4K5SkciGMGRx2Phdb
wTcKqTRBS+LmBt6lZrwnOk1wlWn9ZiLDGgAkzWO3fqH/5k8vYqloR5eejdraEeCs
L67i8vbOjM79xhD6FTO/Paw2AMU8SEs2bxYHo7kqbecDIx0GH+/gU4Rj1ZVZKtzL
j36c3TRQKbX+WFKHFC4txOk8WLrjaG5p+guKvRflIqkR2b6cXKXF8kM9xVg5+0Sz
n2xlyps3/JxfJYMG47jpSLVrOvKNFUAcKMu9jlxrWLNHsmHiRcoq9FTND14gastJ
2bEQ17XQhGGhyszXFro/91S6WoFBSIhz8sd64SUgS3hoi8ZCJp+0rW0oD4MaMIAr
kqa5YUn6Q1PCrkDQaAaO1IBj9cOia6HD/1k4s9LWR5GlAfoCuVG4oXH+fMmh1xGX
Qad0zvA0/m84lf7ZGWy/O1eiQBRnUZUVJJESWHlcqupZoawqnSyYZoiLNbs1gCU/
t+jJUzSBC1u8MEcwzwMCa60q8xLsIVFblBYsBg/QoOqAdrgPIqFsPatVbnBYVjo7
7Hv3TwP1/Xe4I4me29GVt7pvGAXQ54Jj2ia5Q9kEJNAvZJX4pMghzMa2kvf7dl4n
4DGq0J56lrwCh2vd/JqbCfcoH2Iw46rWCw6Df6b+FonTtrypHNwPDW8wdgMKrLKB
ql1ILj5IFoOalGYwmMeZNrWruMKg77LVn+luqGCXwFj7G5ienXTHIPsbJj2Xq5Lq
BAUwKcC+zB4/soljH8I2/FVH4ZHOZLA8OhZ4uQD5Qc6et9muwWM+Kl0NDT7NqkQ1
HVhhNNC+ZHHLTcQ9KR5LxcuTkUKRDwbOrMD4TeyXFXiesmuw++873wDthTWhK+ny
awR8G82vKvCfZafL9t3ylz7e8SST2DEdWTmShS6CEKYcasIUw1GZnyieb4K4Xa+j
HkRCL3uxDYfagbjIveWMJgJRFl8dyLFsN4gIedmmqJiMZ4ybFNwmbvVf3dVSaIL5
FGfwmD8iobcp+4SZADBA9wfv7r1uM6O6HJewmmq6yeTvTH9/pvgB81VhWD9s6Jax
jupWJBoGrQG6Mk5qruYy0627zMnNJnNdkLFXyI9TayCe8vxYiNjK8BRMnu3oGRpb
GGel6JP5iIGrkSDRCieQPjUxXwX/y0GjUyUBvCMeQprtEoSS+Q9p8AacqTC6+M3I
6lGSGZeqjbIaGOMFm1vnHkJl62VGo/X4v4KPpGQGlJSmlJ4a3FKFCPlKWwMhFR6B
muGtUB5gLHv7E7NTZbseSDIf4EH5wOxNlf1HoZx0QejUCZfVOMNisWvQaYlnk82k
O+hNR0wHbyNJjTuFY+di1z96mMLbBpROUqKIIJvOUvDmvTkmXlwxcoKDnSIkrdTn
FfE+4EqGTdi1MDN9P7IejqO6gFGhKLAMQqJix1QKF4BRCvDepgyWhE4yWhH9g6wh
eagf4vcvN1VGCyXMyTuSsMd6HiGDyVheRRbVIGeub4vcAS6tuykT1M8QeLo2nmJ9
5AXazjGom8p1VX3e7vy8GC2qTdEBAF+ouoc1ok3eisuAUEBjAKoOVX9d3E0q1H2n
z4olrgVCzeoo5ZrADox1921I09jx91c+R5MWIeUnKPI2h3ZjJqm3CPDAf2Ao2wE4
/Szo06BSJKJWGzBB+wWHQoktE7OXtXeIqXvl3+0pIVev9s6hUHhsutINBwK/diN8
0Sc6TTLYwzSCNpI0b1D5WdK9ZA7CFk5dGB0xpnr91lBVBhYJNmf6NZybbOEeIDut
8NJxg4kYuut7s3m0pGyP7op7D13N/0ZnzaO6j8ZUdmwah4F378e/w1IWTO8JL3x2
W+dzctq3NFj40YFDt48qJtTNlqu12OPxrnzvXmdQ/7RqPqSkaNFiMbsWTvSdpovq
YqduKxA38TjtVYOsdywRs1DveborauD4uKV8zIQXs3bLlJZiC0h/QAuQUntYifDq
o9jFXXKumb4wV9xn2daQS5Plp5jO83OWH0ALI9jZ3Ae9ps7n/kQR5/e9xz4uKe6g
4B7fzyRXA6WynEAeMmTmYXMDtkICVix5VAKbMOK060G21KYKz9w6kwYQGpP6UviO
XRE6g1L40rUfC1OeVSmqQutMMeDgvQZVOC2OizxiHqYlHYitHSQCC5JSn+04DmzI
EMmRXCmOUay12nkkAD6i8G9NZQpiUnHZW8zf4HQUtcnWq+5ws/NBDWDBbburAf4p
IRV1m80SJxd3EZOmBJy18VvBHgfwTRTdrmWHymMD9+Se85a8yz+4gAHYK7LyIQQT
xzqUu9UZBkzKnLYW3VXZ7DDHAMV2gNNce5DJOxN8NFoxhvadqxNaxdaz31blsgm+
1/Qdhzz5hmdcTWEQsBn9cwe7RU0IRl1DBMroJnahZ+bEt+iVHmAcpDO3n2PWhhkx
yco0S44O0alaBeIzUfPIXGavU7OaOM4wvFp/A3+2IO7im2Q9ZLW2mII+Q6nTgWDo
3HPlaFWdcC9GnX3+aQUa1s3xhAnvrUyIwVD9teg8ifKUMudUmApaKH/ficH0eFQy
IdCgRHve+IgI3cUFNykHuhbM5c5GSQW7+tc3/ClNkYEydm0R/bqv0LiszzQ7HQle
Po19z9aYO/budSfjPCiW7MwuqlFLFjGGPgymga5u/98Ow9tEViWObcH/KUz57LI6
mWHoz5hwpmk8/fH1p85HGwnwG93f4TzL+MfvknDqfg4PApf/3uDjj7H6dGTecDyY
gc9tihW7jekd001kGfk1rTl1g2tgVSAI2myHHGJXZElztnri0RRRkiXZmBYFw/MP
JGEeQfRvnljWex4urMoMPDb9cuD0/GEBlcZMLeGkNXp1PXcWRF8fm+1vLMNotWet
Di8wZliWXWbWTW6zQxbArv4Nlcffc2az8ifWc770ktMe3QRg9YHOLYqHzkQ1xRKf
y1By0zTQEgyvPYHaA6DxwPzBU3ub/aVzeAfg+5BHM6FphhFTXNGt4jd7rfOdEh46
W0dkwKtLLHzIQPyMkifGKq3oLQ7Y7Yk2azvuES9HMatC35V383t5gKw1qp40GOuy
kT54hrpAAECZpaEs5NfHnFvvwe/BAqTqsAK+Zg39lYGlsHWEZZmTMVAYy/6fq8+C
VHmMOGewHc1hFUMDSFKyWAudZHjLh+75RLJ2hjgen+OSwuLjAS36gp9lHOEs8ZEm
UE8KZlPgB7pYeTn9OL0kI9NK3rS0W6JLNP/ouOWWQII00rcyBjgpOEt0GrCWQQmt
gSJ/Wm6Dj1G9+9HBKIzpUklfJMtraG0YgyPIjYfz0SZbbK2QqIWkCYckJW+zRAJj
vWv72SEA87mlXG14noD8deVbDaJvaZ/jZEKuT4LhMhXyvshmmWu00uQvkrwCroCM
l5jXdDVRTjvAhZ0EJVtdU3mR00WN83gb9K1TcfkRmu5V4jUCDtd+PAfDqdLHyavw
En2RgyJnj7zrbdmTXuHiFMTr5YjNMK8ICjOw0G6x6Zh35aDahEd2z10+JWxkSgZU
Nh2Yi6+c+nAPLHJEN3qDKAwN1A4wEoD1sEgro60ebHawCQtxEEuxXgYakAdee1z1
hfsImDqhXtcxsUkwghZ94ivS5o/mpiYm+hqCJhQTOjcj5mut0y2KARRiOOtfKhIQ
C7lpoLit7nE0CQ73c1Cb1W3DF5qmbBKx6fJms8lXvJ25xneVfdQVNsgAgPkLRaqz
PeUt6oQ5POguTysqSBP1TryP7WmKr41kvy6gZdl2MNP1LVUJm0v5eZfYJCoSv9+q
G7Sm2W3X/NIPvq62jsMJEjZsdDJvGD81tENqLOkjQRUIqFHR54DR7vKPfEOLarQ0
bM70KY+tuC4diF2ECfJf8kdECY3S+NnRAvke8kG4u/oQsvhm/nJ3gJBr9tMC7SYg
wGbyEZDJUZjVzJcy7t9PRHWX41hi+YdovR6C2A3dFLu/9dCx7cSi9gzJ21NxtjE0
P2EsSuB8RQzdgf+rvIwwof4kNIEgm5OVuhyDnWIwN0RsQWL4jqFI0K/A8j9Yy7wX
CQZesaxzGahdpc2wPFRWOy+CSfFNPfI12frgsQqv3cLz4vCAeeJ+SuwhOmoKUc/A
6BmniHbyWb/OrdP9H5R93kz9sqNCTw7rapjRCZ5hU2ZmMJXPutSPnDdWCYzVzNvw
eu3DccqPtqAOU5ysoDkimzajr5L9UEVJ1PyO/pIHi5Re4ZgIu6VjOMD1X4IagKyV
FSpVFGJRFMGifp6ipubOBRttqH1k/DZYZJHCdId4bHJbqxP8W49CgWxzkr8cHRMw
ULtFwfj1eqUveEA1ijLphpC48xP9SJfF7Ay+VOS4a4fx75Aji/DOLB3UKZpsV2Da
nvKF21jj4Ov482ICq/oOsgt0YxKwTTceM05pjoVMOonDBB5zIOQttungX1PjV3cS
ACYOv3nMh8A0cOCXdf5xpTUgCKgUSv3MhYsCrdhtMeQqG6utTBSqdGCrC1xjW3H7
bUGVcVeSkTkvYf0dw+Vi/V6yn4lNIpgXYzJy03G2j4vocpQ6cvMxUEacfSDv81n3
Gom1PQL3rOrln1t7nsAcdp+2CvPug4Dc4pgh426sFRIoVLIte/ce0B7g6g/OP91g
JblGAjgP+XaPLZZuiNZQZtaEc8xjjz23D1dxVJiElbIr9yt+YvZ9wz8gbInrEGOY
S9oapCAWmpZTUhLaf88PerCLbXdEf97X7QUyP50fcRV4GT2q6VvlKo14dzmFASq6
NIUBb3O9+7l5RJFJ6heZpCllUsR4tN0MrYoVhP1DesvKB/pgH8W6HDKtzRVIK8Ke
Qeyyv365Y0sBELQ4fanAL75/i2zxScee0MXmELdx+anaKuNayclvL/sLmvFvNGXv
FhCaL4CUv5Dd6DXmgWi2u+So2dUYxhFSaNnefLp5ABVRqcQu6QzlRKNO7cVhYrPK
b96O3Y7eLUldDql3A3DPknoZozfA6Wljqj6AfmqNUJYZ1h/7+OYgLuukwm6SA13X
ATS1CQhoJy/Lmbe+jjseHEMDWPOltvhTDwyOKMpFd6GEK7Vp+DjiDY7ROA2Fg6vj
etSkuMid9X9Mnxf1kibFz2NwOARnwi2VSMcanNCja3rJkQGHuVfU9DpcDF38yUtv
KeIKu1u4gEhZGH+ZS9nfItk9kyvlavyGFBXvrR7L1aBEUAIUl9LEVN8rZTonrpDO
ZEVPliLHz86j0dkz9/S0I5BGcJc+G/uhvCY2ALCqnbzC2sMae2RyLlqjJQ1XZTWP
H8oIxAeL90SGLegzIyYeh2L1yPleqYgT8H5qozJTzryCKPWeaX8NYiImUUVEl+E8
GrzsfaCjq1FOQ3PNdkdgGcMjrN8mxVBmVGwyapCMOQMz5IpUysFE3utaGW2exBCy
Cnecqne2fb72sDkBZZW92QaFDotthtFpXUXmkkjhEQTyYoDM4X92bpdoIlWwkwbH
h3zAv0GB3bZ6CnLAz1ryTROxl0GIvPNyiBWk8e6T7htIdzfwvp9AK5DwrZxDd9Jn
DgUfIb67K0h/2U0rn0AE/XjkW2aOVjbBB7daGkKcdbWxDcDoC+dqiUUBcdTxd4Ip
V7WHxZOZ00ddubKBVBjIx3MK6DRMHb8GDj3o8JK7iLmSfxa3DKED+IyONaM70DfH
piPonL124lQAP+YCLu1KkVRkXxXo8eGM59VeL5cn+Dr+PYZvdy6OsiXiPiU/y3O0
VJ8SWGk3EUbYYqzAcdTbEueyMP3hL04OM+F0XO3NNzufGsqRCMLnLxbk8peHP/I8
PKtxxIo5oF/Mre9wYSrqj7Am7jTzeguiaJoGxjqWnQyEDS1N7Q2b5uvep9f3F/ZL
cK2qmeRubf84dKa1YgkAgieuXRuRP5K3aBgYjq+a+yvVTpANqnwbkfRFmQzrH+bE
tVHsE4ylQceKT68OkjXnVirEBFKQBkFfF9shrM6pOMCG7bkMgdgj5Uztie13Om4Q
iek2azIhwmiE5qR2Lb9ToAkPviROnt14pE7au4lVazsH8o5uuFcxJTh7t7YOgW9d
DUAt6blqoS5DSfVOwwPvy3QVH3hbvvE7qRRjqBwLX9B/xbvcXG/vUfTzA8/+PGG4
xoQ1RXYMNTaBcTJvyJIAEMsWRyJG7az4Fw4ej+xAUl4zh/ZJ/05tx255jdUarplT
SeQSx+EawxNPHBQDyQ48kdSgvyo44pnbC3XOydG3/pmDrDVBcICie7XQs+bzgIcv
nMRgDGX46MKHYerfQh/nkcSKLL4aNXV6h3L4zN1evGof8POHiINKC8vu+q/cVmcC
KGW1HKMOt7zbtH5ei/FVvX5SGu9wyjzsszGNvGF39Z8zVX8YNXDBN8Q8tgKXiZKn
09pEbzRduyP2FoX+EJ6I31hnS4lsdBo7EwUTGO5oE+RmrovGlXHnIhT2F/H+ZNcT
fCxh8fls5EH9juDknQawZ9sOyDfMzVYWFJYfRtg+L8UG9fi2H1KCbj9xi+IRcrvp
LhvpX0MBlPV+CG2rk00MVx/57apjMpdQgQ2u6i+3GWKKpzeevvoczJJUKSkmifOn
NMnVP6PVPwTP6M78rnIm3oWCbqXeraMGHS5Re6uM5WLuWOg2hjjRqnir0N7U/IvN
k/DqZyT1PbJ6/KAUNPprc0mMW8IfJt2ufnv5JmMSfNiflBUuRtMRS4Aojl/d7DBO
OXDaOW/kVT1h7Bo/pciUS+oC6hEx6m3I9pXf7ekz/8gFodjHTjCQSjbLTDrXR9Hi
6vEATZesVW7Rm/rRXZBayEAS3EQ2CVweHUgZZY+5+0B7Kjl8MpX2O8wcKnRTsZTC
mrveDDWY5nkGI9ltd0R2J08R8Q20xkUqn13aQBRiZfFAR/K0B92AnrwxZF8X6azv
RgWrL3CSsAhuqjJMwz8GSIWav+gbSGwZg7sKqp9g1r764odYY2Q6GOn08clsD+os
mfYeS1sJg2H78tET1F96dg1qdeiHA1j6kMAr7h628TdHSlzcFXBr0/m+wlvhBXVI
/dQB7POBC+HNMbG6tkul0SHyDMZSWl4dSg26WGN59x3W+aewMZNam83QKV3Zur1X
5c8KUplxDOdyj6LxAeoFeXcJSveRxFwczKjhSwC7d3ygP3NckrrsL0kGJvij4hZI
RtZulXXPUzLwMNxNRTj3EfCnP6c2VJSj0gBgLA0zHjz1kW9b/+xYl39U05V9vKWN
nq9BucRjNa2ep7hfYQUzDZnC8y7J7LIAQ5yN77+qHoJt8wF3kqDos1iz/PVjwBZY
NshVNQPTsfdZU8dXNM0lZebeSf8fan2CUXZ1BKYIDMVRVKua4Tl3YLvHPS3u9ifo
xW8W6AzqqUpQxFXWpnyTeat8xQOBPxIYjekKX6ErgfvElXS4v7Mc5SPd4C4bos3+
U6hHnfN4Ych+Uw3q8V+ekXJFA8iu2Gd9lVsPrSuWuKXFVT6XrOIv5ziF8aWv9+cC
MnmoXnf1nPQjDePrni3YLLTcpHc6PHmr1N/kzRPUZlPlGtl+IZMZp7aunt8ifJuR
pO4r3e6OO+gzB2rbiXIHmzmnO52IQM1GqLBgQLzoRTq7R289GiPlzTiKO0Oxwogp
0qOMYON/G4+67lqToXCXuBr6jusmnD/EJ659PqGM8tXx93QnVqcX6QhK1WvmxNFj
e3eSl9L89nnG9gqM7QWmFzQPNXz530KwuwCOlp8Rx6NFGJZu7NT99yS5zwmS5JLl
yHLc+hVuK5t9S4bDBdoFsYruZMbj86CkRjtdotSd/jWtMqxwAyN5vTHdSzFOrgJ9
xcC4cUgGu6fFbpQ1GDbNi1N8Xj50y85OY8xOOJ+Zhu8ZoSMZiurvCcBompk3rSkB
zGU2nAcduPwWafX3Bfy7aOgCPB1gHrxHGHXRPK0hFhdHKvoXBeoYIGD5vw0kPk0e
VjPFgGE/4WyVwLptCu7SyaG10ZFDnEWdlCEtRHu7JKRdmSB+lkVHbopDpBzl6dq8
cJZdODQgs+nK9BcHHG8iJR8z9xjYFCrrphWUzZgaJuNJRw58pCTSMB8OqwzMYy5q
9usx2z/g67R71vwmjoPiG2LD+aadqPzlO1ESJGSHGTmbW/Dh/j5BD3u19IxeKXIh
aBeo5GZM2Jd2WuYGGxe8jUX0tPG5/XrqGiJLg3YTv/VvmOZARekggyqXfWq8HBpc
jlA882aKfWTktZGSSU4rxU9HyKf2JTnaMQ3nWWM/56zs4ob9Gkf6+rySXHWWXXMw
8R3EZbcqj2H3kNBgRvzMvp5f9dCvo1180LXqUAPtdLPlNrb0XxtQZD0oxUwjPaAN
Xgfktsw/K+Wp2VrGZjFmlJNwvwy/c6mERM58msravcsi4eVh9kotq+wHpUkC86Bk
HuB7uSR5KneiYpZZj17DlURs0GWsYrIKfkvSuZC6Dm6ikKjoM+lPywWB/9WrFYvf
MBwtIG9r6CBaA/vyrLoZebL3JCvgHks91BLfIG/S2T+6T9JqZZpR1UKslGFhScYH
1jLEPZD8hrvpfYRAbIIBdaHwlsV4n5tEIFpL6nhLAKfDuI2hL6QkNBdJewNu3ulN
wLK7jSvv3jQ9G9DOhmyOwPYGQgXU5h5AtTtuol754pNKSSFFc2nPlQjRK/E26kj/
epenaCwwvckSlWTc+e7+Z/ZFO8UZw50Abwof7UcPZsxxu5i665DcI3C/4DAk3MDy
fSykPn7w3IndKtF0d7dI6Viyraqa5YZbhlXswIxiYOkq3MB7RJRPw5l+RXqOySss
0UWNRk+eohQE0M2DiqhZ7Iw8y9VE5s1h+R99ITGnl2PBF8vtSIjA3UK3uQGve089
JLM4befSiigpeTRaaK7rl8b7LuDayL9Q+dzC8TuRqbGbqSS/Ilz5uv+qKqcDFWxc
RgtUewY6XrykO0eXTjJ+wMqnOZfVvwKmpCgYV3BaeDDnT0dmaPfd9dTZivLvwlIZ
uCLfxvOegGwoXpLWRpYHsMm/2gphAXUIFD5iK8s2maXkoVN1yxIZsMhYCvNVpHNj
2BykrkK7w6O6HelLSQoKE7XvvkRRZn5wZrW+HS3jMARrRevc+91bxP+OcbslLKQf
Qa94qncyWcQXPe8iFe2h8eWEH/z+vWaMVpYYEeLMMxCd3oUw6xUSHTUhnoXiirPk
GBIc42QXCA6CS0JZFEEQwnATgjWxarAUy7NGf1COCMbrZRwYQLZ4FiCthocratw6
PF+QuGAEe8zqMgahUyRWK/C5nzbyOEgcMqww6Z8htuk45Li9OZ4RmPmjVvJj5Vqu
98OVjqPkOm8JPqZlHSRJh2zUQ2w2qe0DUFOyuMtmUDHc8+5tTPvmEsF8lA1cuOio
sLi7aRQcBGngGJo719/13ZPXFvi9+qA20wDi3M/Jk5OkeQC/phVaqHbsvKY5us3g
MW5RW8BL34bsTIuCR5lLGofr7oI4lWhdgaZbiG5ajANYyBjYGtlP00s5NHHehSmo
TSB7ktnboaBbetOKctegEb8WZxkdZxYpGUynDx7WymE2hVSJhU2XPj959BuRdcAf
YCLUDSk6wLkMP6iFDcyikCx/HdrbwOk+hsRsvj2flmSVvAGq1qg4zjA18Df5Xhds
bevgnXcJ6Ajz5/3L8QlyMVMbJrIUibA5OZkfP9YrTq7Fbt4y9PZS2uYBRb+pMFx3
tBqaAgu4T6r1zDOUU6Nn26Aa8Aa45p2kP0d58Oz6ZnFKGlv3LM7FcSTHA1VQLXKk
bz+k6o/AboU0VPdTNOQLPKQsVZ3R9Ng4GzU20eQryYbMKk05DXbgJX2a01fXPsFL
AkLEV8Z4Bb+ZKPJNORjdMOZx3qOEYrJKSveohX4FVAaMpwJX1fHxyTsdlZzeRF7o
QolBPLkcHRHUJ7jOg81gcdacC2fN+jMBmF8UYotxYTS9uNQwtL+XkXDKMF7eNx4Y
xxeq81HT1fgVkVQ+8qg2jC8AxYeepTEFjewTzcPb0NI4dhp2EU4jNxKPFVEQ2Fdn
5HG+u2cics6zNiI4gDi02mFOSX/DUZXwVFkAxhuvFbc6/yMylCFLxiCxFuWE26i9
SUxwcH6CRKqzQxhKl+FwKtGX4hsDfOPElKkI2OuHxvxHM+3plxndVE3Fbrr+6kJu
ReE7zu9GWAV9VYbWZP40wo/Cb+SKQAjzVBWg94TMhkDCvqKCYoPgXTQ5hejqwa8X
TGYcmWKPrux3kZ/s8qCXrraCivMKMIqCCduhaSSIgLVPXP8Si4+C0v1PA8gelPv2
Pl/4S5lHDevozyiGucTgLrU6i8TWTTJ75q41tdDXeRRE9nWYKZkFKCFlBlpY9fQ5
8R+pmlDTaL2ajMbEjiUW/jqDguUzOb6fCl7nKpl7PVP4ymLa7DX5QdhHPY1G4/M8
RQ876PfTtPSLrg/bgzemJpzNkmPoPXI7XakrPdqloU3XjIA+eRHap4z1QFW7mmlp
l4Pkn3kPdkzNjVRM/p0QIc5chSvrt+PJDF8swoMzmx2lrIb6UXNAlfD1yjQ2z2G3
pNBBvwa16njfkQYsL/jp/wEuyuukeesluv/0HDltJLtf883JCC5Y/jpDz6XYMdsh
ZjG1OXO1H3VcZbNJzTT29x0zftqwBTd4sdUCtlchYxDzhRJv4numEcBwu/wymf3t
U9X/hzrHKNmSWoisUtcHoJwn8LJb994inpppEIymH8ZCOvdjl1Gvx8SK5oj0/4cF
LzVT6BPodjX9FalZPmNgKcOPpcxlizFg59ctCkCdK43cZ16psXaHv33T5kGzX9ob
i19q2bb0/5uDRlFnN6QWr82uNcrmQWO24PP0a+eQcOMDHrVZdjyMF8dBFId464U6
UpasVWQwtIUASdQ1BQJDSQvJ8du9LW2mD836Bc+q8hBjHF9k7Dx4nAqqvXWzsQ+c
D/8K7x2Aod7tR3sefXtUz5maALjeouh05MGwazdPmvpGACbsjtcQkJQAtIPDJmG0
mzOL9Xabm0WG/qevLnGSLmYHmjDGE4vqT90t/6ywik7GZEm64UYW6d+yatvVtbGN
q6R+gH5pz6sq/nJ0YCtzZrv5fdHAha5gxdEBDVCf/G86l7EyOgSXheITMNGBQbJC
9bpy/9l+4Rzyo7ZaXMCO6MkWldmcJE9iTAUc68ixX+mEsZmx/IWi2v7v4X1cgb/j
m22k4Ms+JIARLsp8aWF5Han2w364AcMjaS6gy/QdiOZRZqLJCsp7x1ygzGio3i+4
2GAJIy+CYXs5OSmte44iMgp0VV89miHDe2bgI6Tbo9Yw+Cw6d2dynsJA0dFnXill
PdTzyeBiQ0LvjACMhWImT4ol2of0fciziiYkcM/FgJd7EWgS54tq5a2eLuikOkPm
FhlycHIIrhtiRfDFpKbj3myVYBt/MBfMm6dpukTP1jhRzb/3E3PK1lEUv4DJC6gj
Y0aV+zzLZK3tImxN9tGGGxj16htPosQNBcCV29TsWAx9NAWtR53/kO8g75crZ2Js
CbhGJ11m+oWHTht4+Uitq4/68gkVJIwQMdBbSc7MPhGJEI4xGd/xqCRBwRNedTh4
jCvUuqj8FRfgR6yhNsAUlDYRByWjpCvhOzAAd10IfFFvbxV7S+ioFC+F9jWaM/kJ
b/FOkbRBUtF8NYDMUGjlzuldy5+VzfVlDgvIhee48P0/Iw7safcbUdoRQ+w+kzta
o/wlB9uyOLkZnb09eqL8645qyrh3OMT9WxX7jOmiZ7rXKjkhkRLA4fH4heBXEYHv
FB+6LvyT3mopvPPeJIfxFSeIsLOwTmlIzHP0DtI5Q1QqnVqYCJmv9lotqKYxKqjS
H2kN4SrUaNtQDCplMQnRo97p/c2yVsQLuMCYlgd5ambcoSk7+XEE/x9talGolMi7
bPfM8lxVduDokQ3QPM2toHqfLWLjtKqg2WvPO0nuGvHjxvbmWtvD2B2u4jvjg85l
sQ1eByE63Uf+8diju0WkOqbWDjLdYby26/tohuOceg9YUs4hcIHuL4Xm7ar5Bb9q
ZcOToSThmUzke0KTgE9Kb73YIJyq2oGdFXbJ7pYoNuuaObhOLR8etE3yFTFUABgQ
NBX39jrUeGpAM0q9jt8zXpAnzORECznKSZTEhxjcnNNPZtUfjGBRahDYpU8cEoaq
0oMtjfMoOVfvzKL07k8eeI9EDkEJubYEWiloHaBAPckPbhtELaoHhs49Z4UkK7zD
HOO7Gh/B4BmYuOFFkHvuOQm7zqcrdAIReR9LEbpgnmyC4iqvDwEOMUdztJ3uShMH
rSSnfssyOg94R4pojgxD+42ND9E4hh0kzg/CNigkchDnKebdAeiF8gsA3Tcx5bZ8
wmYCwL3EH6Zelxm5MgPLzQhZ9O8b1ZfnK4xnoJjig55NOpqhg+VE73LMpkZWrM7k
EasfEetIqp7WEjCbfOlnPziCe/erKGzmXaYAiKopkvw+yIKXZHoPXy2Hz1XobIUS
LCL8KQ6/3DdYv6IGUNwtP2N0rkm0TBJ4wuslghyxtYB+DruUrFH0RXi7cz92DfKc
Cc6+fclu6XJ+QUMUgiGQBSZ9j9QRXRy1IvD2hGg1X6DeCBE9prx/rGuHwp09jSHk
4jMzK5Cbvh+YLq4maT/3epv8LKo5DB/6PGqS2fhRJ8dE0/7uK8k424s9oOiG+eR/
EZNJvS0H/a59PBulWoZCCQbI30nzuHGwWRBvgUvxH/2TY+D2KD4Np2OEDhiWRx9X
Y0q6vpxFJqHN2ap0TCao9ltWkCq0lRPCSbDd0Yt1qLcNBszcnbHom1vRVDjSwd+P
OWd2MgkSJJ1PQ09sGLrA9LRNXvtUi5my4IlMDrQX0OZ0zyAAIzZsuY/faQyzSRte
c4XLjiHcPgKtUGBrqjeZlLFEt5dou+uPiYvjdwYNagD3hAhRLEXfX98m56bzJ4Ys
AoGGUfHJ9PKFrli/jXwbSTSOfab1DAkKL13sk0Dne+sp/6Nfn1tCnqyFFGxnuaJt
PF5OjyrhbnmLJZ98naBaRK9k8CKmZaQodxsvtOQ2C5+V4ywliSHkNtqMlTX0wMAg
5DzyQrSDjHcY4GfE2BF0RF6se7zcW0JztUM3tln3djT6zZPMzktwdRMmKNiEqu60
AU228P5Ah/oFmPntA9YdAZ4T6GZx8rJWu3J/RipCDJhk+BKtDNVckIHnG/f22arS
X7xvr8dA7LSlD+lQIb9HfIwnQN5VaLuUnBOyYiRvuPWAkmNPfCXwGlWHX20rRi/r
PvOMSV2eREDF2vqmisptZYP/QLRp9unn4quTG7Xo3rgXY3RwG8YEFWAZBmRM3pgj
J0OQ2W67qtPTN1M+aIuAJrkfEAmNKu/zc/ILrcZQEE904sxXv4rixiXTkodBLtTT
BNlwCEAOxZRzxAj1f0OFNA3B9RW3Bsb04tX0W/BUALRUbae/73lBLyyKZkXUaQSw
ZEjr4uuzDr7+zhlssbHAqK7KGWK+PgOfGPAqh/QbkXITii6UpuGnprqQNupgIdw+
w3aEnnqGwCSgtB/QjwyiekmXMgoCvD8US38y82wJQMkYkOnCvDDNcyncUhG1Y4us
fNLGdB8YTGmBDZSQihL709qbJOAue2ki8NgMJLmo34+2ijWfTgpd5FJgo+ap+RiR
is/WKNcixqxfFVnrd+88mQmBgfQPk0d0fx8Q6bNMdzN69zQMMuA5Kw61xDIESInV
gkmlLAq+iNPW7eRnVMcP1p0IFJ8559HhsFT1LXBtohpOViZtuRUqWr+Lvzb/MSbF
nab963GrEs3NNA+p3y6eguWRoNoPKbkdpJAHjCbp/ybO21MDvEAqzpyUIeRBU2k6
v+ABsReicQ51Tdr/5RoFtE82rS17bUFSO+dlZx4ApgLfdq8t6xZmZOzY4n/MR/2C
EhkPYralhs7egXmKRLJ6czEvj4xeUT7JK0SD9DLMMGlOaStV9/ESo22WFEtAEPka
9M71FGJs4+5TAHRw95kDTbAROqWU40uBNxZmSxGuW2F/JUKWum3K8un1LF0ijubc
QWnj6FJ/huYnu5AX9nzXWWV1Q9JU+U0+Ee03NwKXwEr5xBV9XaoyDRhJEWe+RYfc
2Pn1bMrtlJVk78aBLIB0XC0S2OYlGjBo73ARuN+JKOwno9WR/7yHuORRTL9Esd1o
fDxSQ/E9KJ7b89IZ7/ugB/o11eebRQaZa61dOkcsSzAKCPAAuoDeycvKU1LYqkDo
7b9ubw1QA0FB0nYNcPIpougodDLpzStH4rftUiyFaiwC+gdbJmOHbzgPFu549G9T
CVgk81CxER8NdbrY80LpZAGafzGZMuQvJMAWhdoqlaoDZobvy1w4YFtMbGeA4yPj
tFVLTBBVGc1QD6xR3W178aofUE/DC1Lvw+ffSgb9O7Y9h7fiBQEbNngIZ2sfqEWc
xIEcnywvkc01924opYWh/61tE3pLCHO81F16ouRmcFjyk9vCHFRgqkgqS8S1H3iX
h32VapB6nJR2cxGeR5JW0WhvtAVXunA0tVgBWd6mRJZNZOskF9bcIYqMGpTEXSF1
KE+x3TSTZ7skle/OfMKNwoDIRYAkWnXd3cD2qmg+c2+PsWgMAU+8Xq0qyL4ObQeE
AXQhAQjKKK9VFBWm2H0PfDeiygpH8USfPQ3KyrZJkPjRRkDOZWjnvsS5/xUg6FmL
uZxMArW7EgRyDWWZIPFLJnRjaivMCPG4d99cU8Vwvr4HClBMlKDRPuWRKtXayhn7
0KQiJCw6PkuMbFL3EvIv2/hrc3f3TO8TAGBdBaVMFe3hGDhMv3eBqWu7jlasFigc
Oq9Az4Vu8nkF+0UbLLNuR6Q3qsZcPtS19YOokzs+l+/FAFeUMKbI+sKHH1c1+Few
b+uV6sFv8U8lpMsIDE+aAUJR6t2GWYRB5opI5H3Qnxf6Ijb47OGoOGsiNsGq99nm
qQp+8QcF0W8asU1aI4UOhFJoYxd0BE6m+linrVx+W726khzSCcOsGXsNmWutdT4W
MRDoXJ2ZSlinWCLmdfO6VcH7mIw0o4C3N7r34Jp47FuOeXBpgirPhUgAERxLBzcO
v3jRxC0rzYiFTga2WCf+yKJSPd7reTCySTCpouKNqGDS7vN4LqJsejSYgHl+Y+FS
KLnAIteWIFpgtGPGUjgCXjVjAjtk/L3Ng3reeYnvIp271u3ls2uozrwp+nB4uEkz
gwZu5XquXvAYWZZajb6UtO9Cy4bN6naueAN6crHltA+nzQe+8XRtRFxHPOUqt44c
64S41zqMw9Wr8IBKQ3uZepA+C5VnCPcc9K3cTjBaq/PvBZX/cCHp7QwG210h2J7f
AQv1fY8Hf22xMyEHHcWp4rCRavUnWly1/frYJyj/gb5Wax3EDQspk+lBaG7IvdoH
t0thz06ghGATEAJjikZvSQB5hyt8dsjmCrzia8k9OIV6zwx6hfwO5tYkjs73yzH1
bzNeteKrnBYusSxYDKV9kH3p6mNt1DZsCJEqRFxn5Iw8PHSsiUZlGq4R8TDIEs0V
t9v1euTpXl6cLTw1uv4Gpzq9Hh/XSuA63uWLnRK5t/9hOYebnop0qDrXgB4lnrUr
p1lPNdT/sJT8zhO/mGCHZxp+3vxcntf1QJgJn7dbdJxXha8x66/LlqHOt4o4smku
4Qdra+K65xPeguGLc3nN5ZQpXIMe6K9jq/hOh6B4x/wkm51z4H6VErDEDnPq0YO6
jYAAIrayqEDZnM2r2XWe4IffpXFLWE1qBhAoqJvYHLkdSBvKuDaZs/oxNXs/Fkft
7192b0TOdbGsJzDvIuDnmz2PVnTFeHse7xm1nyPtEfHKpoSuyrlLHF/dMSkHqVSK
EpCpYCMnRiQDGH7Osr0p7bXilFrYHKqxJr+EXncB35gGaZNmojUwRJIOrERr534Q
bwYKPOGAuDIrtZYqBd4nuRqSte1PxKUd4b9w9CmqegbO8WZDTtAEiifCLizqvMGW
5gEsrFXIfvwoees450ubIYxMFtpbdOMzQE7de9Sy4d6M1vJgEjIJvNAvDB2I9KjF
hXKIIbiJpM76QihivsAkYfCS8Ast0KWJH7U2UId04JB7ogTPjXTA4rdEslNhwFXn
36L26ulzmDKbKf9nPOlEW2gcUxKiVE43s0ChBjG0sSfPRd2E+JnKTSoFFO7GNmYZ
hfMnlbjkrYvIa3k4NeJz+Yj/zVskbS+vMUS2rKu6qe7tKgFkDM/LhsL/xvZM1S0R
A8EvzIfkJBx08M7+VO8FaK4f9S2sEGcF0VaA8L4OJcJZILKdtiGLP+73ljdweke8
WvBcZ18L611xdO9Hals+sX0V8uZBDrWX+fpjcDShj5U+bvCNLQ0I8ca2EHttFQyB
gWNgzJlq66h54z7yKjEMf3PYU52Kl/AoRQEJ+DroRdIxVtfWT+rtwIwUh6w8ZR6/
rJjka3cTQ7MCRUbdM/ILCcjoj/nJnoBozsEFRt76genV1DMKGC9Qu5MGu+2Tb6c7
/7Ms+D7MsaUA+u4kkpYF3WJZqR5mZP7p277hy+iJMjjFHUfwEYFztYUZ+RbRdQef
h6I0HuIg17Hlu9VFyN2s/b5hmJLbm61PZ0Qxl6SBBkkO0BkWnFC1H6hBtPdHD+YR
u7h+ayBVAAie/aOSE1ubvRB4fMKYRT5E1rwiVajfZPHfC35rH06xqIbcPo3XQob4
NcCeTGKqjI0vsnXUIu9c3cfkLK8oiB8Bv0O0bAPw0g+zWJ2w8V7vQn6v3SEAIJk+
nwqZ2rPZ9J0hb/5l0ObOHoCt5Ym3BmMQMveDqnFym2eBO4gli1rZ/E95zaT/jIOP
NW9qF7YxBpGTPbtv7w8ok21S03ui5lIzRfRGJji9oEC5aQZOtIl58hlygywzFxj3
bMS5l4XiO7N33S0MTeJ1WyHvWo035bKj4jJPKHXWg6hBnyIpSGleuq8AUcd57Bzx
tn2tT8IWJfMTXmd3oZqowFjSXfi2hvBDxtgS1ns7lDtmVykGnv7wLJTGP9kZQ87M
kmFIrfrMOdVgesbAWj9BUVfP4F981G30AwAuUmjLcQscE+UK2m4m6y9XiHMkq6yY
cnMJFKrAaIxmXhLGadZQyeUCJ13mKIi3444B8JqTkEKtjKltOxQ+koJh5q11DTla
go1qtMDoTyL4qgK5xG4fT9ZyHnKyS6EvwxhcHSB+QCmnvvLHtw7ogWZAJnk4i5ND
6ehi21Jb2u8fhn1H6sUsn3tvjRyjpa9SsuRHor5kFG/1BudnOxDlXpFeDEE1j5M1
drpS4Mjgz0VSVTbArdNMYLI4u74ottRZiYCMa0Luy4+jSzP9V223k7lFtFfmBVi0
/LmZbVZlNpa3x+2mOs4SNi665HszLb/P+uZ9esPT8JIdbHjx2OBmkOAjvUQIQdlQ
rZzmiKnKMDSMfHk9sLYCsHenzJQ8TVMOrBe0dw1DwucHgdL75OSYPyOz69NwkdRe
Sb6hxp4ps9pio4vI92Jnq8SV2azy1CjXFPJMYxmoXjsCcaIzg786LlxAbsLH9JxU
2urn7KbKSid9Ki+iJ0zuSHbrOKSh2770Bao0hlzvmkmF1LYSaSKFOKtYXDvAq1Qb
o9hwIM/tlmlCqcVPZXrQFN0DfAeCzLduUYmsoUoffNvH5YuxzadC+XiUz2KdbtzD
LNLF19wstCT93I6SscUGywVEpp3Omre6hewu1LL/x6CpjMAAMWFWV1KZh6X2wFQ1
Q5hBCWNQn8V9m5T/NKgV3Uw9D+19MHjlTtUMis/bQm5+b5hXF/0VXaCUg9+W2meS
6c97JK7yUFHhQiQEh7TnN8WB4mK4q0k+2dmid0SBi/u4EWQ2v9XKtI/SW8iD8NIQ
fTmhK+gFIlpeJBl/vHLem8+xMk6oRNvMgD47HZNewHFRrPTBN3moWpH6zGvlq0nq
JBfyyGf5jKCjddOx6zdlkqO4lYov3RGPzj51/w/Pq2AZSM1CAaKZoXT7KGFWQno9
v+Ii2AhjdkQWZcSXmHPzEPvgkSxVnEKVT18cQGGeUMHDrGQDA8LWASWcCBLXMxl/
pndf7EfYss3lcb372azKEEx543lKgDmahHvoV8z3O8qXQa9C0iOcp9izlRy/xPnf
/8lt4ySZtTXmsdoXv8q7jVanX6okqQoDXQXcnxChX46UWr+OICepkZrQAno1ge+f
9rIYo3yBbD0LjKVPnXcwshvy2CcOYU6J3q4f/W7zwrABINeL9y4NPbwZANMDwEy2
1DLRBIHoKnYs0NZMqtIWivaBgCDR5Etpy+ma3mSYvIKFZiRS06w2HkeUjLjhlRMJ
WZCI3XB8BOY1GNgcmrrASaAaq0nN/tqB0opPkL//IgErAx4HJ3bsVGOJ5nQSs/Hd
1oIbSE3nivvltAboTWsN12rGonGGeLPBULCGImduehEWTFcMDAw0/HFZvuPx74q0
azUsRmyR4CIhkzsbqzy5/0x6qaOq4jSPLLYhY/+1NER+rizfylTi6yvRqqCxCaBh
EP5/heTXju2mW9Soi5gIIewNgE5uJxYGUHHFn+T/GoiHa7GzeqvPwFF+mLBO0NWy
zQGk8Ux9KMBFOHNOdRb1Rj7vAlQyDXocSslh+LUHq7c0pxVXsfEUO8Qkk9j5QfbP
dRsXPVAMEYUVljnHdq7Q4FcbPwed1NPestuWhi8g6U/NNXujr1mEyTZktHBHQ7G3
F7de3zz2sUUjEMv1GKvfn6BDfso01MgeYqSV2aZkNi3+mgrb3VgZvgKsm5T1uXIl
P1dqmRwWfmjOz6T/FRRslD3HuFs1c+KcBNEKvJLiKSAHjfEHhWJkdgC4zZajR5jR
gLmopKHPlfsYV2GRX0Geieh8ZVDNeiz4j/1ijhb1wdanhPdKP0MTz4EDt+pqh81f
P6MFrgeV1wp1/aK3d2LIvyIVNRW7wSie5wPYK/yFg1Ytptr+2dRsZzdUav88yTvE
sX9YxdUt0dVOgW639sEHmgWOxDWoMVxaPsB/e/8Zzic87UwmYwLDS1lWn+mt2uGv
u4F2Dg/TIc3mmX9/NHAfsZDIEFN/iTCgBL1bnuV/RXy3clsZFRexcYe4sAu5ca31
UMuNJpQFyOBJpHf8zvOT/y9EAsNa2SJSR5IDZooPPMzCxfh/CJ7cNvypl8BW98v5
JU9eRzP5+dYfZgYQuyz1XPYNRFiiuvIePpx7n1adVbtgAWrlroLi1+ZxHHsfebtv
4JjSmzGJiH1x+xbAxu8oqCWP9PtaAkGVlCdMoBd3DcgPBH9gZJ2uUcINUcNEkyin
Hcg/7zqf81RyLitswtj04TO0ILoQ9x1nC1mwv9F0Zj2d5TWNjoAAE0Npzlg+KWC/
c1iNYD+OcjxQbaoYRNiOzMx9jUH8Lm0eVoeA0NY7kRRYsr7Tvt2VqqRXVEhr/WAp
/SZ/S19+f10+DbJTcQsP5S9sAUHgfVznIOgpeWE2/cjaLYYlB/BH9OnjrTlcPFb+
maqmpa56JsArFf/tEpRHa35OR8CzIOrugStb09VfG1IlSBOjUia2nKQa0i/weCAD
iPPmfKbrA8wXhoA1PhI1RxsPAcAR/aPurADu04hn4ckZFqRzKXaLRkKfmoJ1m06v
qWXj9IwP3lhNlsJOBNVeV2bnVhcP6hIPZM4RshWgEpXpF6bkcgzM7RSk05sKLbOH
qMsu7nX2iqut4ILpM6+e2jGSFHXKWOP1Are443wsg9+izu/cuu149sG3Bwtwq/mR
vZ6YisDIQ3Hazc/fc+QXcL3rjB2CHCYjhWZ0j+K3WubxnH88UzjoVtw6Y3brFq6h
xLf60IpaXOkLp2TMnTryiHEUUMotnHaEHUode4t5+4L4lyXxt0jLc1DS97gvvPJv
Mfy6Y5KHgID9SsmSNoi580HBr+QPMv7AGa1qOySPD2LYriG5OyuajHTbFQWBMBxE
ZMypLSetMIk+caELSTk1XBg4OcF8wfexFN0mt58iwPVbbtY6fYvqTzLMKtypGPlt
Im2yBlFCq/+B9Y7GnvQ8J+xe0o3i4mB/qTUGXbMs/RD1Q6JfzgqfimUS+R1nXTdk
H439axVh/nLPcxor2qd/HRjgSSA8jtevwRCvTWFrIQUcFXVI9ABOrWUCaCcfhI9o
EpglY7AYF8gz4dER7I30CC/aNQzzGPNRA7vKhLdjLhvIKTY2KjyUVosuEc6Jdu6c
MZ/ObjT2TIBqtI+IENiwOEAf1kkWEEzD1RGbhp5r9RLPEzzmRz5b1K2W5blRKB1g
7i9cYSJSw2Fi8tAN73bhVDNK2kj7F/k32Z5+YIEz/jaNNJcw5BhZHKhvqJBOUOm8
c9Vsn5cHb46nDQS99xN5lfzuL/nXMHtKrSIVtgiTK/OUk45ereI+Pq79OGG1fxyb
8waf3DkAzj1OQOROa9k4Jst62uU5NtRLQc98SSsL3UTWdUdxx+e70sOcMyvxjFBq
Vzp3gyf/Y9ZIEiCna38BMd3RfFRkkRustgolPOUiUgGol3AGR+DS8JrTH0OQBiBS
AHCiQeyzJxg2kBMj3LKvbtc03JGjdNSPJkT297cOoU1R3KSHYiwEmlwD0yakHnqs
AZGimpnxuRH+YzAy6DluTVBG8dImamLIUcmOOl4iS+mHhNy+mrsd2FWCx5w6ymei
zXYM3gh1iu81VBuahlPQKFReNIbbdlFowzwf8+XzvdEndOeMu2OorOqzC34PXfCC
CFqBkvAqdWcHq+Dzm1xzTSczXl/nQ/kbH9dlIXYazjBEDdqXCIATId2A36+qQ/Iv
gLz2fjAo1Kn9tBoA9BcpmSMbLR9Oe5LYR8YiEeoiQQeSx5u8HW5/V1kUglogRqG1
uuW29lM0d8hbBrU2h6WaUGTWkJ0kOdcysfiUv843eHSF9Oz1QgY9/1QjZflk+Ta4
KdINL8huugy44zDZo+D1X3ILUVB0Lr53GIO1OqwRrmgIvcVU4Mn3KIUTTCHhWxe8
Pxva64LD2T/h5RpZhBWmnEEytu/aroncdt9EXbvKZMVkxuapduvwR32dk+VTu7z1
1Er4bg9if5F/Z9P8/qj4dqvswyLm7IxSju7IOWGwYsxvjnL6lF78FdJg91ZBq096
jTfI0sAwYIMc6Uto+gC4MuW/th4kRMuxBnZKBwpxakF4WTJKjhOgDQTJ3MUobi4u
DHlAOrSFvFU+Q5Qm0LpwmlHv0SzoSIe5lZc5hWamWZzRbH53pTlex2J1omYvzx28
LEcxDmiDu9Jy7M4q2e2J/0cTbC6I2fz0zMNx+eTIbDsDx6zAjMsQRxr5X/OAanNy
Mxr4U40IC6kKzfk/ExoeQwd1bMOKLHv0v1Bvt8kZ1IPCz9Qc7dwO8yTQm6Ine+Y2
DGG4ihZGK4UMZEPXNrts1dryoddKnTGWVVoS9zNJYP+rVcXvYBVH1jOmrGotEYYv
m8Q9RyR8LB+bS5SM76/YLAyma9Icz1VqUjeK229JQ1POJXTFx4AVy9yGMNQWIL9U
4Y+fRG9wkX174eRKVIDMxMLi87gEkXiiiv/4S0yazgNPcx6QUZtcn0wtqfPivz4r
AnshlIB1ra4SwaGW4IqI2qk1frbcmusDF+gYNJppTW11xKlHecsrqrxe7odNwHQR
rBY78eLYTqtcKam0q2kjzWEPOAK6WWNcwVZNZ3h86kRxpYSoXhfDxowOg53RPO0r
FhAj+g5d5JQ1gQQT1HqmDujiGx3Mt+zliWbaqFtBrSKH+aXbnTq8xjyF/fZmAc6S
y2iz8jFEYGJgi8pE+1wr4G1RVGCiYCQQp5/DcuebPip3UCMMNpuVj6vU3dGfvokk
Iz+ZhCS3pvwRXILzzjOjcdHHVWJYJ4GmzpLnOE66/3ZMoUgnxZHLOnjbyho6tQ/b
goENMyXsAoqXtnpj8FxH9c9yD+STrrKgwcGOGG5OYervvzNYsZFbSNqgndfHMuwF
8xBUjuckv3AJpNhXdtVwaVH6G7hRcN/Uq8dwpLLNtYpWNQAjyIwkIRuUCDDib4dB
6gaMT/TUNRMzcLfmWp5mg/xDi9BwoOW79A1l7x9TXowqe85GBr5ZEvDNG/8ensf+
HyEmfDbu1vWTSXgZAhby/rky2w9y644QMXc0JhEAIu1foVdoe4SgzApmwOMgtBFb
5ASFZiVW1x/p7gDLWgGjH8vwlJ+M3IlYdRwzEeMk7KfV7wEeWjjKb6qjCUS1Q3r9
Bu7vqLcBvGFID4HdH9cq7FY4Wgboov3Lhnp0UY7oNW0nMtXXy62dEGknyUL3+7Gi
odP3e+DwMl8EqR8HnfJKjLr7ePB4DVDc8b6UD0XwQ5epYaqZpzahvMGFXyZo50WC
OL8INAL1izXqQwvW6sbn+gxfwAHkWDYvWmDATmfXgzY5L7vnc7VyHj43KJhsvWO1
tAhYRYaVsk3MVQFD1DHu1oTafdZimLkHltboDbbSG8xR13cG4JRTJC8Tp1vUySGL
kuT4f5PA6Si5LACtiDWJtppAm9HFVj3Sjuyy+vQgNXkCfP3rC/LIs2b5PmetD7ix
HrBdXq7jPLaXfskhYZqg8VnfCleRGuxv8iSUobIl3Mf12/CBr+Ku4JYt7rFI04GA
3wct9NzaMXPqjXdbIsfCGOTk/KQBkOX4LzgLWA6vkK7vXAOY0SAcncVky1hMZ517
f0jXdM44n4xwEezdrudTHVh29WLAflbxYzC25noRL5UjND4uOAwzB7W5cx7kK9dA
y6FpwGeXhJc6qeyNu0KjnRrYbFteVjCy4ydA2rcTQp13d4lhXfl7aVxH7LAiWU1c
vR1XIyA8j01XL4/odes/asFB4pK3MQeCr/nRX6XcuE8PHeELulY+6Wm9nnz5aqBD
Wza1+K1TNgJ3EemVBLYf3BikfaKz/QVwpTPlWE9m5mwCiGHDbGQ1zkoHQdBH4/Az
3+7vbnkQpbHG3qioptVd4a+y4cXWqDGNQHqvo+dW9SlrgHc04nhN6VPR0mkY0jKS
Hdf55THPiE/pJLAUThI5QSMscyXHt43zCD0IUhSQsxyIzQmOL0efFyJGOaN95bHB
Nsj5HhSUsFA11sd78vQQg6VbA2wJXmd9Xi99Cygh/HMa/RfMkZTEs+V8cq/WmB0k
TcA0yeufuH+nH8kLYn+k6VENgJ1ZcIeB8wk8E2YTgZk0GRJgP9LNpmWtzdWds1j4
knV85YIvED1Ls5Z0cvCbFhY0WZsQ07ABK/iIRJUeoSsTHqSnjr8qVUkcOCAQ3bVD
QujDwJ/Ezd+oDCCDd8ZI0xDSgTG9CVyy3MoHo/Nm5wHIptZQ37zvL9J0voc+Tn3t
jv1I5mYdvncLqNULCuJBvqkeLi7Wx/dZo8cAg6FXJSkdsxXv0ZJS0DFkl1WHOYa0
d0ZpAMvPRNF1hlIbe8licaR0KBjLtT31TfJjmaofx5kbekAGsD/b94YB/8e9n8ui
heReRAzOofrT3t7gZnEPG9yTmoI2tOQWcjEiWkCezpqzzQPqxjtMd5hgNRreMCTJ
656yFiHb5JGxrvOKDYFD3BcYA4Gw1ub+j/3E/V0OPC9eY/M+2p8wgG1m2SPTCS+z
rmo/0OxKmOlbnii+3hnK4+BD1r7F+vAUDTGPbg/urWGB/NYf/TWBR5Wiuj6P5fMi
1btnBHzLOWqsOd6oSgbLII/8DgOTObqQea6+bG2V0kHezmDDY78tflyB5diXo9N+
j8DGuynDi8YTZGfJ2thR7EbUmHYpWi/tTNYk3S+XIeKAh8tTGa+3Rmx8KS7ZmUq/
hedWubu7fhdwd2GREuKU8Rd+zsfSHM4EFnRbYdehZGgRitCsIFHzVjUdJLusaWFW
uzDamiRimQEddjY2hMKCMCUN4CExAeCo7M1tMG1aj7QKRxYPO1MUZXtkwdpIHkO/
bE768zKK90Vixo4u7OYVPAQ3m5pbYSiKoY04ZncPLxNKgjwQS5vN/jMg2kLpe/vS
ZIkQUIw+go2MVVpLG4C0PNwksXlbf204DMqwgmRYVUvSExtifU1VZ1OysEi4QbDE
ioCiT1ikoWpaCcOIFkNlwvEh5Ome6gObc86gqpaeiqCMCcm+oGdeR1c0aKcLfUJ6
xLje1M0GJyClPLCj0AaxPG24cU61hoe/fn0LiNhpKqZTrd3ND1BPw/YeZdm7WoX5
/n8PW8HvvQOtXGkswVyIReRozRaIp26kiIglqU+YzTyvP+gNpYVa4EQoMQjCShXo
K6fZfprIF8yGaCQU4jkUPwgDNlWrH4wHEmv69GH9tpqewkGk6ILLVc/XSlh8No1D
ztQWEmCRNFp/HOdCPjSbST21UHOwLlieIFhUzUnx9SogSom48en5xfNlMKSQ/0VD
QBHaSMB3eS3U48xb93nVNNE90tn0x2HWTlEFYBv6p3dJHxc/tTXZ7tgvHHs+9Kgd
36Jz5hPKcJZj8xnt56EX+DqZnnfwlB9hYVapWx3XsIysv83oTpLGacku3oW/zlM9
pIdXOBEwQTqkQOeEPXbzftZwc1WAd90KWBdtNuBCWUNMeObe2a4MJjHRiwSnn6R8
mrkzL7QHtqWHvWizv+laQMVxQGt+V0txID1CZpHRjm+yEGCvGxUv932M+oFlLxv+
k6BpaWQC++CZ6axWaikK3H/yzOWkPaPtyn8xcaz+8vpmM1anxtJCn2T0xmp37/QA
V6oLAjL7aT4Erb005T770S5uN/JQQ9cHz/bT0iSSU7ijntkc+MdipJD2UDOHa2Dg
Gzmuz0rUDcFvnKlp08CzMgSPgRMwF6v4xQjP8Fa3cwaT6wXgTA8PiAX4Ajg2MxDI
698ZVywuXSVRe2x355bccU0P//qljJ1H8DRpyMe/WdDV2hGpHDgt5kjkHoxvHnxq
8AaJ4VeesEl2WU+AxHRvPR8qu31hpmzfgacAo/hHmgo5TEivV32nqU7EWfqtFqTR
/p+9yPWdRoHt4D+CXP5P+9fXcHMvyG3HGbE7hJrY3ef5TS4t/t2igEguoZ+TTzmo
cz/E/6NiSkK+VcInZNkJHtT3U+YlF4hHG5adWsGZsnfsShZN8+pBNNcwnpm2fCQX
dM8LEyTXd6fwubP2Lf+R88VfXgFy8GprKHP25NQtPb7rqAzxFHTPtlzbtlESr7il
gWd6HxrofTuiR0X6Xa+/vjlluWkyepCZSN/wkFcQrznC0Ajnk1ML5/vNYJYMWjHc
JqwYbQiyEImhP4/A2/N6oKst6BN5q/lJsoFjd7FDCamIAw+zCMHjVEYxEuJpJBxN
a3plcVNEtG6OP+tBpLDl9lenG34U1FusFG40YeE8t7NcE0ulUR4VhUJDRG74lkLV
G9cFb36sA4HLC5MTEIoUrr3SA1GttJJ6sPkdPuX50EYhZGIXnzfUXm1TTqGJILOJ
WYDC8EnZQc0aDDNN0oBCfTB0DeY6UyljovkshyY6oARzHAqB80dtt+cV24W2AhPl
aYfKjyBXE76poZYB+lQxOKK9YSuNi3qsErlzvKBDVa6ez67VuLBGhJKtrjPmpXC7
i19xhHO6edlDaBlLURvO7MGmMpU48uODlmsey6N0KPNBbHfa6nj1IMOinHqqTm5N
MJAbJNisoOFtgF/Wecg9maKrr1nQkObiwcWuIzP++p/Per5nUx9LYapJtigz46Aw
Th1BM42IpFRhAGQ5Vq3AdM0ofeqTQuCCO7CbJ4SelBoEoVDtFJYiNpgp0LPvPbq4
Ap/nUA6JRP/ap6rq2rqOcDsVQeMO5pun+/sVIHurouRBWO1CY8VNEdyHsUf2jB24
QTVnbpbapQyewjgJthk0jWESSWioe90kL9aBCSHBQc/hI9h5oE7l1gXzjEcy7fr7
FGY1EBBKWb0r4BEhdef8kpgCxIhNqZbDDFwzwhBQL20Z51mTBLKKeWVc9DdeRpyX
NNeTQX7WQfvxbtBYSrZByby4avLGdBJeV0fAizANoyr/N/k+SgOwdxk4y/5vl7S9
WpJ4FySJph+nZhNEcNl1FU4jPsx9lTpSbmVgF4sSvvdolYg9z/I8BoGST62NyJv/
IVkVN2MHTCMlfyrP/K37goKQx3NmyqeTQFRqIH8xSjkorAoGgur6Lh4LfeKaovX1
0hso9jF/tz3ZdLL7CnnHXZlu+K6wgZFAKqdxAKbSllj0fkH6I6+OOnTm9bDHbWxf
GJiyEoOJQ5HnqJ6emk90A6EzAG92gKDyEtiLxfdM93NJplCj+fRYuTIdmpVYHQRg
nlNYL/p9T3DjLoJZ4TKksaMitqHZ6JiBvKR9MGFjHawHEA4unLYk+bexlouYCLek
V3t9LlYd0Mc1YJa3df3CC8nTU1tE0zp+yduz5OznoE9BknUGH8rrCA0JukAeDx4J
XyKlwgl/TXACRxGruIH2Qhx1TZBCA+uZqyE18jd4LNR/uZhpm3HNDtG7NUpZcN4X
081Zz5YYjnJ8x13QaUIgcOANC0tgP2GzqficLhaVOVQClUdB3mMAGRbqiLQTlPL4
8vkaKUvKXKL9guAg1Oj3NdSQ2A2kxoCp2OL817yBmtK0WcOFcCSeoh+jv90etI/8
jL56WAQ8sS+dcNer1wdjUDMFqG4YGHVLrhGI7/IP+Lfwc/+jFruxnJEAMNZ+Z7/N
cO9XlofzmaW78VbQLwc+lAjIRWDAIHP5kDqqHJK8RI/KPSYdShEqkc1n4ze6sRz3
VB8ZZngXVQN/FoIJTa0CdQe32gYRIkzevZ/rOXi7EDzNZ6gcrwEVcWkMwCtlM61b
La18K7Ci587pHyiTSUetcm1ClSi45FEyIvLo2ZArpc8kD7Ef99ZqzjAjesUYbQfb
mevl6M/NTmjpQh9wGcdURTkhanyqMzp6Nu+TQNB1TrMvzfBakuMeNAgDt8leMfCP
9LDqcrTfV8xY1LoqIA/uwxssySUVvX5MWtMNjyMlzbi+M+TZPCKdI/XYBiQME6n6
dNuMEuTU9+3Xeq1iFFwWmxDcUJabVfnSKBdySueVh4FsSvin/rsuUpy+WNDoZP/5
4YJB7VBSKdYLgipR0LcftQzGl2JmxthmAOJvs1CLejd6S/yjeU0EYLRAXGBPXvwI
m+kHOqyfR2xiVY1nF3tny76eo6TqRguRYjS35ZICN2TL8F5ExBthEOmZDQmgzSU0
csja48A80ggXQbwKIUDHBhRaN76uZVG5ZMsWbQfFBcc7brZN+IQ1eRNL5jBbZmsG
qsqeJM8iR2o4TnuRX9Xyv9BVMBUCdB8RmK3/9d3tkk5TTGoAji1jCP9V/MA5EIJt
rmBwGlsKyjl2TE8tULyEx/ufJQ6ANoI3t9RWJBV/y+3o2n4bpyOZ4ZBDT+FeSNxg
gULKunSVVBu2DKjXngz7F9s3tt0f5MBA/iA/G9Ejq/hs6NUVskuxrdtxLHqFbKAB
XtCyJnCnafZmqW71yySAwnjUK0WHob+vFoeUuTZ63sArhtp8DQaj/2QYfZ1mxJZU
5jQ5gTVzhqcXCTwf849Zy77IoG6MR/HvU+DGuSdoMiAdRFwJftu2odAw22Apmtnk
KHnux9NFH2aGriQN6lDoGNmrUb1zxuFlgpb6GX1m0BSMI7BfMNZ79MQFtTzdBCp6
FR3+3XPbT9J8hIMsFHyldFCkVZN2rQd5aymbIN632O2sjLKmTKYqgoU+xW9HiyEh
8v4LsNqp4aZM3UMB3nNYaVZlhcNBGMz/Z7dcX0E82J7vM4OfYd5tvPtqj5aceJZu
sZ9CJZRFy7NSaLUTcuwIscfLEdAbFagxqebZ9QIXtluHcdeyy9KUzUY4Ho1uGd3Z
z1ii3b/UUr6P1KuHwlPNtu787RcdxMr18jpfJHsY2F5ZnP3TraJkrURQKyj7KrpQ
D3+eCVtK6KRx19oykagD7Lj5pPEOV8c/Epmgrd3TBGvB3pfXcCBc0FvwLSAuCOeg
iGJZEdtKuLRu8957oIihVjrvZl9ICGanTYjIAaaGGEKNvgrIlVV4gISC5cmDR6MG
TgrkZpw0HXwS1WLpzQ83dZfZd7EP/6RGrS+vyBefX5D7dAxis+mi2mrTCvuDw8A9
+VzAfYoKfri7fT/fPu9A/tKrHSTkP9TLlixpTjGIAhU7XDpMgu1QXd2iCVojkBfe
zT7F3IG0b34saaIg6ZnzA21vWEP9dIcoMSlde4ID/PlTfTVNVg78FULEWOf1sMO8
eK8aC1TuewUOKVY1MCOfQ9Bxq9Oq6TQQ4JLk0hV0GmmMuX5yOQxQYzirFte4EV3q
IZ7ZC0iNwCp+yIghfAMrl0sVY/9oskVm8jZonuKv9OVe5KrfR1RNCysquSIFR1AX
rj2wx7ILpL2kTUAahBHVUlGlnL7Dr9EujM6L95sFD32szpdf9SSvXWtjLCSSiqV0
s9rSqJvIh/hke0smxTMKVaV9COTXt852kam42rP1Oe5bACY9H0+1Ww1fGl9Y79mu
M8MvpuFhiGuNTueRPxo3DrYrywsXK4TNfgVydt3s2LPpBoVvXZlgeIKf0gvtYFnH
I3L/hd/x/ueKfjUFq1PIUznLGBxQH73G1KklzNYvj6v3manVvOckJdnIp3RK/JyW
luSb36Yuf/qUX+m71q8xFRUu1fCMXWUjkrO2ZPZAgcMEN2LY87wItHUeKv/qajSC
ZDOZGGD3L8qe01NVjstSwKHBBg/gF4unaVeW9LT1wvczl7NNFOFDEbfiGnw/xgUC
ZzPEhxOotVCrP3iZnnYjXa09+eXrTazKCHpTlOuQ9eLmper5OeI+0UhAQHvu6rQk
rd0DVxF5utHw8mS3ASlRdJuarsiKibtlw7BqPwHpyQ3FYqjjfEsFto49S4X4fwho
eteT1dDuNOv7xy7IslHVmLon+idXIkzXPe3ehx3+y5j0W9hVx+2ri75n/o6OX5zB
OMI9qPakwiuFeuTopaWo7sghwc1N0DAwc/w3Tc3j0lvhC/eQ57HZLmv+6MVWQAkw
neAT8/QQ37gzerbQnuReKOMT9CilPLbXF1JmkxNWxdAyabkKB4yg7w3VNg5+ju+7
I/Cad0A5YjhWJg0BjxKZBKOqiMGzoi32d9KUH2BuGPnRYvCRZjI8PvlVU59KiIrk
Pv7wuXROTuEZoTH+dzb47aYNM5zakTvozmfC8Gf81c/7elFWqxuQth7AejjtsuOx
aQ9PFfK7hdNYFMFOOQ+5qKeB855esW131d1tpgKq7txRAL/bIpnrGLpc7mzKUJNp
z+5DLZSwb1NUaH2mc2abFoT2CmMS5unvkCjOmhWxLB+4eBYk2tFnGFfUnNYTZKeP
wj88txkS4iSJHC6Os5lGNKzXRmrUjY8MUF0V3Cbsx0Ica5ioKyyeT4Yrktv7eB8J
hynamyitSStVkVJKxeJF/z2Ktg0rKj8uN3byyAk7L6R66aiMuzzhdSYJj+qxIlxF
5YBR2WF3XQjnEp4ha+bjACrCORS6igAhF3tFDM/StB9En+9ZG2WUq2d/NjmZUj8U
/i8vizXAawqA9aR1f3eeofsULIr6oJ8uviswT6y2UGu7Z3d7UTV8EF97zbbmI1uc
+zgQ3EVKATHlJzhteRYmJjRsGDOzDZcnt/9I0baqxd+wdzmZ6nM0k18Rvqttt0JK
hYZKS+OCa3hrRM6ZJHV49M2HzM2w1sP2hOJhcBhO5fiilOBtTD/pOoZDtHXT3uBt
RE1fpdXp571IV5DD/0RMUXTw4A2y4F+OrAtPqbdkROALmic+BiFBpzZ2Zs8rnYEu
qFc5pmAleVne7qGTwO7x8L5rcVSlobTzYnV/L7hZunelmeV2gP1uH1kZkAreoYgy
ME6LbiyCjoZNF9UCOTUgzDvxP76L7N+z1Fvyea1b4MdWORsnCMVWJK6O80QBGQVS
omyqbiWAiWi0fKq78UPkGqdZE8ygPh3kULe3/NkkLerAjTi6OFelV0Yz4ofDXcqk
XDtwBPwSTc7bv2KwYoza7/F01ubXF8l3bbDFJNcy6HUqRb6ehzksd4FnC3PUTTzo
JBlCo92zpsqNfH2s7ahtrETnuMXZWhx4Iwd7st573EAZBbjkWrbDPBiFrJ7CrLbA
nUfSMfhgWysrT+Nxf5ITsRQuwOBn29y+dJomZBoBlVX+zK4UhXzqYi66yAQZkXwy
Yx5iR10xAcEw+mt9gSpfSrPFiNjLLfIYDXHEdI3ef7xZ7gYuGj3Kps3SvBjn4B7R
l2nU0XBU7JKy3OfWMIexKo3lhdNV6apw+u9maFQjieTdtQ/4h3qj1i+TAWfGemK3
jo0RzdF7IhPOXiqqluy6H8HbH1YMLKBrdYa/U/66dgAqPmMdr2ou+ZK0mNfpmsip
3tfwe+GfPzOitLQtQ1zAeDqqETxj8baf2EFHYZhE3K+oUiikX8Kcd/TMnwxbLHEP
4e/7f7MjS6BNOIiClrjwFrDz1ThjYZcRdk0J/7a/dthyARU6zWc4iJdj8NDNVQs3
eBNgtVS9uJffETVa25LlNlz/bCXxid2FS/ilzay0zcafnj+aPOvcqGLl0eHntsie
74uIeLJY2/gnTSSwoPsQik7c9JXNcWxvt7UIpxyyGsQooOB8m3OKvhIvfgTR35re
3M6fx5ZRadqVFFdFmHl1l41+wqNArYxrzp7Q8OFizfHIiBjfeQHxbgl4rEDwF1s+
GT/X6M7hates6vW7aRpehTCtAVIuHdCzf5qP9uibp87JlM5MSN1n7OM3gwkUxMrp
VDx76wNGQW0i4YcDM9sD8urAdIkqVQ4+DuEl0GwDLPqRwzu8nFybQS0eKnnszp2n
xkZJwX4C1Di948J+rKND1bspZJ0ElibSUYbqgupyclyQ9nvgGCjfX5GkGAuHu9x2
AtAcfC2XGmWpeuNikmT83Kfktedr1Ube1Oq/3z0LhW5WAanjBWRiqoGnq14Yhbrk
Suna9+ZrVg8U4W91YfsUMCwxOt8SApG7fNfonrIN3Fo1U7TVZRzw7D7yhHFKOcLE
LO7nohLkxUJDaXyQ2dq2qVMrnRV0kKf0qXcva/Bzejx6xGQegKxPLmFkuf5pam6V
BwyYdZBRZHwXkWfiLAy0hb6cEGPBKmKN3pn2b81IRh1MIZf9/TG6mgjZmkAtsIfV
WinaSu2IpLFFCPdSGItxkK9x+Vsvlil32r/ksqAwy+vnDbW18e7X3ugYrppIPSCj
1n+U0eSPwGvKa+9+65RTl+lbPAvMjb/i7ibxqnNXxUdJtLtG2tIxSTxPIqaF65iV
+IdJI3dZoIAaEAWz72cyx/++NxaXlKRZXZkXv3La7scowVWXg9bNrC4HU1/C4lwz
m3lxNGOSQzYisqeGsTcXek9dfq01ekaVWUVH3lOtcw6p24NptWN6IzqU1m3OjTLk
piBbiAnLKK3ZPSlf7njAFh897xT2FQXSDK80e/dz8BXEn2/14eO09GXTAwqjsaUQ
nkEYjAJYWDcoaAZTgzEyjf//XmpowAc2jOhaQ4ugrv1B86/yIw28S+6ntsg8ZHnJ
f8RiIMtLxp9aDsM05fyM+X/wIoyAyO7jPGAcGIq/gdW3Qsjj3/R64VStvLVAVFy4
Q3F8n0vFNdNY69WxUfe2Ri1PuhuJ3aYQgIt2kAb1BlXf0G6vMC3An79gPcC5bhGP
s3BYHA7XxH6rbUZFrojujknjqMzWYSqBNPVU0l5byi0OhQp+E0ei2wZ4pCBdnIwO
RzFjkZDHQwA63aq1uZ+j0sHdoz1kr8+4IDEGOBhjF5sCyVL7/2xU7zIObD/0IBbz
OpsZrrej4zw3JRjEfwvg85H9+bqI9DgG02fSkVLmesbf0iyNfn0AYCzt+HUOxm+q
qg6ZF5j9TqQ4zMmiUPjxt+2E4B8ZP8be3eBUfMGRmRCear2ivaebL3x6OATbFt0G
W9FjViJNrOt4n7d6lzNvB7IFKPjXMQzCvbCW7zQF64bWJ48s0PuqVW4Ftnp9gSiI
BW92EqrwPJWHrDX6KAWNWZ+DvBKrsrRsZw4J1GNg4fPD/jpErXbj/2DCCVQ67lLp
Ut5SFQdmAatcP4vzlZzaRFycDGCd+YonOP2toa6JgBa50NQw73FKNQ62WrpP9YsW
mHxjn+mxTlTgYRFsDDk7c2y1tocVGw4rOiSntMsln7hlxtwXTMD4+u1XMbIuAdNK
bEix1tRqn0En5J9I68iigsoxOmWLaPOqYPpti2yXuay3OVxe4BhMcm6mhpemQacQ
lgwxBkteoeM89F3WcB5DoXLBaC/rdYCl50Q4yIWCVsgq1AN05jvl/g2lhWciagzA
xCzZVD+qM+r7gqNlZ1k9/Al6fSLGI67zRM99xdipqoA8Cy5f2Z7OboBv3yQIs2hL
B5gNfRscwG5FTRo/5C1AmhsOx+CX7KS/crFOL9FWaeiyxzwwOFdGWdW2uFlPT8Fe
R/HV6WhRF/5ivCheSLr7r4MdyQsjpen87ghjxyw+HQdfSbRCKM/k0KmbQL71v789
6/tosAT7rZyPohYyDHLcbWQfGnl9YKloUrwZoTGdY2Wca7tMjCH65SBwkGudiuFb
NRo2XB74MDib3v82TNADJOsZgKF3paXfXV5HsjYvJxMkZ3noTxo7LsKbPUTQppPF
VRYcFLt59JlTXvtZILvWIFku+0vhEjy71UYJhVAsO03a2PsaHGxuf96OeiNyAmjE
UUdup/My5vDlJu5Z6ilXTdE8st/hBs9dvmEb2Pg/meLE1vHOJGcU7+3orjxUsmgv
vnHAKj2hJCvc5veU2fFfVzueinl4LZ/QT3Nj5cqoI4wH3EEy3EH20JZCiX4Cruek
FEXU1EqdbrTkwjYOMwSY3HO23t6wmAiWNUa0VgkeCyDe5b+6ZEn5t39JPgT7ofIq
KdxQbVQNDWMhHex3ymSi1CkLEcVcvXoqB2r0bMFJ4TtCWqOJ0dyq4dyKBoCXkWLs
6QCLlDY8VZcmAKCGn/3aWT3xR2gu0Z+RrY6+icPKWmlv1U8p5mP1mK/RZcKeeVRo
aO21nvMmsyNxWBg/AabPjbDmysylIIvoahoVpQj9YCaNeD7QZweCRmMdtClNYdIC
Er89JCf77OP6+ga4GgLb6qaXGw9SzKq0YRLUG8gnAoVTCgEVSOH0zI+4QurIU6NF
Ti7DF9KpKe+yB1YzDFTWqXIbNIlWyr8FYLkvU/UWJUtg5j0LRHLBMmyHehohmhU5
+E+4IBKTa2N62ck/98wWgg9cyWP9XovGhUNklmwPZF6XBaZE6xCtT0LAlhU6kJkN
CGyMCSKkdFuBxLvuJ0j2xKB1PqHjA0ogB0cb4PLC6uN0dVDb5C6XQ4YvMfHV3mU2
hYIzrItFe+6mkht91FqiYZ5DyiayGzw5oh8ZWZFBN3ZK1uLWKAyGFkwo+Mr50zJ7
8Ze5QSosUybi2gzrSLBvy/dzdPdgtr0EvL2nnIuN10Tj1eu6iYEw/bddMOC5p7tc
89pJur+BMuRRLW6nh5GnKKsF54BGfsAk4bfGziLMxHMP09uEZYdHtNr24qPfccB7
AgmSunpUUaSovJwmts2F3f1HLLhtySSHag4fP/HF954Lh7I3dVGbG0xCSwOWE891
MEtiUvF3W/Jd97HZCwjrWLxNgye+vLm828Lsi5ye2gZvN0FSuCNtSsS+XiUBmirO
cmMApDmoKR4qIv8q5Om3QgA3e9iVSLmzQhXi42Mmzyw8FIRRJdVAbU6csxKiATNU
WWKMw+waGaeyvnF+1O1U4v+nPI7GMyb0WVkTP4MiY/9dfraVxE+f6MxSS9WSJSBx
E6CMWYPCpTKRBDqmbD/szWETX08/lg+ytkKtTovnFQr5nwD3XMcWHrjdEQhucc5C
tnRK3DwfkFhC1pfTjGbnUujouT5mlqIg1Mn4R9rs+jL+6jxWXwIbZfFMsm9x9gDW
WksALY0yvAizHB/Yz156lutnoK7OZPwyPTxkCopeEd+aCIwyu1Q1w3aza8xon+g2
10mPno5eybicjUJIaKLgZhhYEY4Xq7fdVRypYVS6njFcf97+53M2igFEFgBCtH8l
kK9fQvLNknjnDthx/W5y11WPCZE9OcHoLBa0MslED1ue7s6D3lRO3Dl5ThHBKvau
VLMskflR+KAlw/h+Vo4u9xcSJ4yyQN5Q6p08RZZa1n3dvhHjeMFeGjwQPudTm21x
6X0vgDNIZ+UVTVR2G2uAzSs8tW5j2D34C/Kc+CjwOpQAqVEHDlkFmgWYJNdq/mMc
Rqp2fnu1Cu4UWYLXA6NLqwV8/84xHDr5SL6fqLSFHkFNabVLcI3IRWV5bpbecy23
VqIma5a9TxMpDkcXaD4bcLBt/zq5oO/2GpcBqgWn8DUEZLUSC0hpSFwgHFk43jIy
FV1VGVZeRlQrMT/5PqMwRkMpP2P6Kk4d89iqT+J3t2OQNjEWkXdnIbmfaQv/UePM
fi5ZcNg2YAnoAYGvb4EngvMkXs8OkWwSX49n3w+Wx8Y2xsnnBihAYosLEdXKApmZ
47Xxry1xW0Ct5mUC0qg+rts1lsyTg65QjW6uFPnSuJPT8Ma21vbNbO4pClewlsM6
qxAoIBHJd2b/bB3RXKZuaG6SjU4k+9EfbOtgmJTofDR0C/P6OsotF/HwUs6IIhzx
4Sh503R2D3t8e2+fQ3qDW9dtYREUHvjZ3uuLvMjI2PGFDAl5xbSuM7W4C353O8GP
fKUvMvJEw/i0PmyG6+oklW5ElIaWC30ZC8axpl6ltHwanaOI5jwGofeihfgGG75q
yyaKjLdaUmGhL2vEFQceIKnjpoFF6QeMSiC6LM0zagVvEcXg7w4pRsIsw5/61Wyy
oz2nRZM1Cg5AFY3R4TFcs1piEbecwKK6iuNuQrtjPYzM5CQJwjMaipjwYXICz8Ap
0nw55TcxWtHcZNHBFC+WZ/ilU6OIc5qILhpJ0yVY8oawugR8h00MSRce6nbDVnyP
UW4/8Dxv6Y3wBStix09j3EP2MWREwkoiBF09UtKnRd8dv94/sFelZmDzg+Z9Eg/5
g/Vo84NpiW4nylX1caqCwpWeGeqji8zbeuesY4CTx2czOAEpbD4N2hyvOjmUaI7E
BjMWviMSLKgrKLBZ0Xk3FtPOU+lIqBx4xreXPaIK/JHzXediZhMNwekx7FhkW8km
jO8yn0tz9qVZTNGloMCOJTH9WE1udb5BPdy44ujF/wHzCSa0kGG+eC3yNDm4k3Ss
l+Vip4Ro4A0jce+dKPAzvvwVmaxTJleWm0q9GW7UxA3OFreEWQcZKJusnIwj4dv5
sjCldnKKX518yJoxDHuuGo+mir6gTPIfTm6QIa08Md221EnpEaiT8deMQkXgnRul
eCN8IIo4PjR9/0r3KpEYAYsH+0WYET0DmG4i4APY3OYeNl8S3Ag9QCespXLtFDVK
in36nPBAA7ufzRaxL9/4mnrBpWbrPsJcepTCCG98WZesFF7RhTuUNYcrcNaSgrPl
QUxQKuJhLjwRvUysEPhzWievk/u2TbryhPxsSeZKtW1F33XOtx72Ke8/Dl9Y3TKi
HhxQtSOWI4XTwJw/Sw+c3RbpJUAnWYGoJ3r563PaH8I2B9lsU3y1K4eBlL1MxK83
XZcKRgkobluJTf8gzcBlMJ7hLAf6fK9gXh3huxKSj/wfsaUkidcPSrDAzdsycdYV
0NoOourZWz9/8qEmQnSMHSDduzcNrh3M9QMlK0cuM0p3ZdMTtUXe9paV+pb3jlZB
XxhvODhHK1J2TQibsjHcB2zpd0hv8JVXZ5GhPcVeOa1dHoiAsyxZPVwY+SSIJZTk
rW6eRHnnDfJ/ywJewHTxS1Ldh0VU49uQ22dZVfuk3qleRhQtBDsp/PaZKmm97t9p
gb4xSoTaAwX1Ww06h+A1HYuBT5IqpBXpb8rHGq5MZU+uDAi3J3o2EJw0isLkWTgK
dfXlrE+38EVUJtBLQaJ4bLEC3Js9Wk5vsvOcamqvcqoTN/evKYmkEssdTiDW8cHX
SmP9o+I52zdy3ZlMqHs4bnjYfhn92VSuVGJDg0HQW4qqzTwCy/VOWy5eHCvzdvtv
VPXEnMIjhA3nMz87A7g2bzFWaBRTcKJFnpKGOdFc8U1KFoNzs2PGSXrrFf+Qh22x
zBQTVjMpDgL37fniTUUY9ohnfl21daBpS/m2m/MMaljmZ5D7n+snHAWAG9nX96j6
qfL+DawnPMwjGw5fmDiIcJK5iykEpD/Hh5e+bgg0Tt7+vsWV2dYfRpb6s+kbDV+u
G/9pi1h0G5RD1zrCdQQUsQWLMpVqfjfehY74ToohMXGfSMl+givzqSHFz+zCJn4L
dfR5/tLOZZ/kHEd38UPeo8UqvfCC9aBMQGpujbYfLUKWCCzZq4MN7lYxmP4ICPaE
F7rK2LCtE9YYd08ONaFkfEFHY3JLwP3yN8zM2t7lbpYwzwEexTAymu8XQeuN+l7v
DLBxf0lGayTBiTpEZuXHtxzYgHQRff2DN1toDkVFiRtqe7WvxWp29aCNQ141P6Uy
1x9EZrM4JV7UN8NxsLsQvR1lpyLZRNASazN2fmp9tsYJJKT8agVP7FC/Qv84T0y/
nLws82KkiVrGkJMqYaHH+jxEdrW/8K2D+abPpdRQedbCkv07eUqvsPCxfcMSLi68
wNve5hZ/LisbyoT5Dm1wurqiYlvjtlRKztveTEOOFSvifK2XbLwyP77Bob1HbEVv
7DKozW/MI4XDJXKVAVI4IawIHKd8k1NLekOOYDrl7Bzaj5uTyeVpHZghnE+iaEU1
A7CuPPcZy9I60SncqxDlWtN8AtNDPaWQ6pj9zNzUm9TV8g3ybWbBJ/FCD/fMyiYr
SZuIGx92jLfwwynSh4NCXU/sWl5z15pVtfMRTaWrbf6b7jqehHDEJ0IVC9t9CADA
EEjKB3XG4FI1hN7sK05tRTQUP/yYNfjnGe+lCEdjmzAEBwhSU6pL4p7IRH34ag/h
tmkUzL/R3S0sqLLFVkf08Bz+qQSDhd10CcJPTtXGa/EfHiL/qheNFdMiYl4tImbv
NSZE3kAyxXTWF4e4+XgAmCwU6at0djXUnEkGg6dDhZCvAQGoK5S/s42tkyIXDrd4
sc1oNlPhQbbqsTYj47VB+1Q6NxxxG8U0URhL+ozmRNNQXJW8TN4+9cN3yfWvZW7o
PBMMcwcY1xM+T99/xqttrK47vu6GOG6RhkifX+fqOvoY7ZZzDIyzyyflBNx18a0N
oRc8HXSnvEoPO2xC92PVSAdxZLoO2/Jl0rZ2DAtjU7+ZtuXfxtS+fxA1+0Q17fgr
aCMPc50GXqNyL/CDSEshYHCSKITWDfrVpqQKmpjdHhJSefjZGfdLbaaIJltlLwJH
LeQx2XXP5VDpc7341JShVczVjceqoUBxEGWl9DIuIIj8l8TFpmJGEK1NoKs7qje0
Xo0M/WAgdF6MF6+t60G5uyeGcydJlcH5y9umBl+gNfTp2hUKwGXOG9pLva2pc+3K
G75HLQv9CFnnmJiWTd5ZwmysSvP8sR98w5mJuBTjo9ZaGGEJkr/UuJuu92ZUeWpH
xl/b/EA55fNDS5S9KXjg5ZTcQ56vfVoJnOv/DkkwYV9koIQkyoQUGlwhSBNPtky7
/GJcDA7Emo+sXOkGGfzzYDVyV8/dZJksphHiz8kcXdAhuNspaB1UGaCmbCDLoPUj
SP7630MTfmxQWwt3erHjG9X9g+5QF8GBtBju5oYMH2ledEt6WQB2W5as71zV2RSJ
P44kAAYzzNYTwoK8vx8eHNSXS8lajiXHXE8lw3UOQNAuSZJphcuFEOL5uQNSZzIU
2yUIKwYnJXDdk03n1gczFgeoBVFMK9ffUdgfUYPoDfNVLYCEerSfwxrfmRlfuqPm
zHsK8+Oy75/nSVqRU/+Vk31Bpo2/7pcc3716qnmmYJvDIWqDKNNMJ4wAw5ivyCLw
0JlmcRLfgxvy+fGseBVeCH4ec4gqZvZnbYGttuezhNIwvtCJjEQBUP9wCNW9EWgi
FWJp71GN3k8CEeDfQBVPt4OYlf0MdlyT6gMXnZEh5onerftNG829s3hg9C8S7mX0
WyP5Njebi7JWkJa+XViYZX9t5c8jBmbpxCJGW4N+N6iRB+HReTpUyvAOekTKrwaW
MekEP9NyQYKH1mHmun8CXCpj0pnxN8BHgJhJRfOrsE8nNA269W9T9kwufiUTQ92T
nNeYawzQS2NTR3yd9GHlnL1RchMEoaIbGYH6GyiyR0vEmB7SbbSR98N8S28ettOk
nyX6GevCSn/gtpanH2aRKcp4ETHtBKdemf+jqyTNUzQPQqStbErmIHXiglO+IZ82
2/hPrEmGq9YWohU8hPrTu+F1vXS7Hh705l6pMMXb2psfKovGu5S9FBA4TPg6+U9K
dCPFafLV7EEL9a+R9+LjcquX3sbu0temhl5CPVjkyEbhgepoErcrPzSm7sRlMTQF
fZgWhnub0fHXlmPxZKWPBPjpGeNbAK3kkSKW2M7KVPi3yeK1O6SK7q7COyAmBiH7
E8ePuMBXz2eSI11/CDx3INAv6Y+mqtxUlmXcfhYyRQuXifMHPVAiZuMBveUl4iTP
UeNL3aKycaQLKV2++2uSc5RIP87a1sZZTXnUC2E3fkGcVdfnPPlkRH5Bh5kNAuTE
F/NyFDp/BMGXiUUAknNLO+z5RG+ybNr9K2tJP8RuIlCj7ibLj/ZnBZkgY+ALEzRv
06eBM5kfm/QmbGaDBkvv/fNFv/8RRqF0A12TrDITwembUV8UV7ihnCHWmqP9Xaqk
277TxHPRfABc4gp4vdlh4ZRSlI4wXNgwTEE6b647LYl3+FPdI0S4Q2fBW7golNzh
gkYthdQ5AGwXm+/uRj9f7Tq+rLYOgx1aTh9TsP+ZIXcE5QBQIPtnq2IhY7qQC4N6
imRU3uFhZ8SNGQ9wvB2GtKdMPvTVXAAMbg6QrTHyvn8zoQp5ZlJXVMyDbOyohsSm
BLBw6ivIMhIbdtVhg9BXG4+vPvGEml0elavu7ZJM/8YnA3fb+Kmq/tVnQB4ALyDI
cYGXHC4qqNgEFpgah4ffU0Rwn4AtUfdheNWdcX9jye6FWVU+0Wiw44Wi8aKZpkD3
jnQR4mdXN0D2zDxZfZ0g3o3z0c0PgkaHm6XNlrp5+6g5y1TXKxWjcinMqdenf1Ek
G4EQAY4D+PaQUWjS1ZlTsATOoiExWAf+xqVWWThd0js0G9hNebOBf4A3HvCZyusX
55Ak7SZdTotv8hTFguS8opPl24YeE2Q1y3woa+6luPpjqSOC8JUhqB644B9wl0TS
LWZd3pTN1GzS0vqaj5FQpKs8YorUuzQBqXnkIypB116gNpHHAIveM2uuHQKTGE/3
mI/8NFZCw5yr8E30nLBQtdsaD5DZoRxwBtwVxn8DCwzPdhIwy0kVkAgjIX5BHbSU
9d0rNM9R0Uiy6hPtJRNHpcKrR6y4nEzWgYvcDaQgZiiZqBqqeb0Zg1Fkff1UNco/
TWHEDPDeOh5nIEytzWmfpDL8drYxe+Cd+i8MTKHpiX9CT5N6Bmv9ecdrzBkfikoE
dVsQTUq/PLHTOO4SdUwO2WkxdL+6Fno4CR4RrHpFeGC75xR5EFX4IviTHY+BTezy
sl9YfOBD2NYF67SjeRM1bbsmRiKd3u5rFSvF/dbSp7C5W8qdOnthNMTM1IHyf0nn
G5XX0HFcYQIlxF67ljrcJk6E3augf4VF1ZMRUj9+tse3esZoqnvCKi90cE/5mhvM
KNNMXRCXiM2xKr6TV2sM/OZoTa722ZBLR9lKNEcETKelGpCmfM0EWjrD8hVBMgDt
pP/MTMYjjCBMVZ32hTuOjg1W5bQGeLyDRMVBr+liix9SiAUMHcVh0OK5ZZOQXbtD
raA0ZlJ9Ve2donJQmrDjPzvDz/qOw7j4F6FsN8IH8GJ+yHp3eSvFRbD3RCYIqfRi
60UP9Lj84uv8wyIlMK0mQmxpCCthrHIZ3+x6jNmDsQnO7DCLY97w0hW6XieqkBLp
ZGu2blGRcRa4PKId6dw5fPaKUczNxzUMuy4MLJe7MpzLybMJa/baAWAJBgf26AWJ
oAklYwZ7lYxw87ZjDziacPVeXXR89LabFBi+dygZY+yGXNBy8Cxcx/nr+K3ym8of
hql4Mip6KICcEhrCNm4+MjUbQsVtPTRr1qoQ3cQX/mnJoDJODqwNQiIyuEqq9CFl
D2o0eD2/1vQPQbXDxYuURla77+GJJbzstNKaquJ6tkjWhGLNt3XPstgPWTyGbKG0
PX6pzJKH/DVUDqiYj50Z1fqQYNh7VbDGR/T6jqB07urBhmv2vOEcY/pPYzZET5AM
8rwbU4nGhwF7MIyPlxEJGMnV8fTBDsEegXkdnVr05M2TR558ZV9bOGfmjyf6cn8B
/9yW7aQJbaZqdf4UB769zGWWkF6wYJ4+ABzUGf2aO+tEcMaPwe/KhHs7yqg6anBB
Z4xNEMqk8dryGXBluPTXlf0YWt1OM7qQOv9Jqn1xpJs/75e2eG1vGupocjcImoRB
d6I6qdz02hJpgJX8aISL1swoG06a/HYOyrFitB1McbHGXwvMJFLYcts2V6yzYpxX
TwYAZRd0STD43Z/PADkxjJSEHamL+C8WFrE7OOwozeUHpg1qnAJYSkRniweIIvhl
/av2jzInfQaJwlh4AckbehAI1e3LoC1EEQIcT6J+FMDqt0EFNQhhjlcF2qeRSfeu
Y2q0kILs920piM0qbf2gUDzof127WteRup9SLVJ9gGRu5mEQznzu4Ivw+CDxDwO+
9nwhWks8q6N6460Rjzd1J+g6VUUD54HZM24N9WGbXpa6Nfp5Omh+E1ZIro5rTa3S
5MKNR7QwfmlEjuoMkcBvL/jkbaGnDK+4Bm8VMRkPqOBVTOdDpx3gkimdt078a4p7
HizTSRHRktLJJokwpafcVVKtEAWU/IdGTHtkMTjXIsSERtO5lpIYvJwyyjkCyRaA
LFawNzvFaCW8Zv1qhWByeZgk/2swXAYa8S6gpclrgLhNxBd9Qrj6hlharT/eooKf
yVa4hFMrPITFmu6ZU1In7c+choboOtRrvUFl+tYL9BcT7EgXslFToN3u/d+zEgry
+Vxx8QHGO20bSNuXGTfncSKUdjiFbrZYQxwQ4tBLYRILFzD9Qj8HEi3CjdAGZkXk
LY6p11eQvgza9gBFxxP5j0s6XlVQMIRI83vfgTK9zNL4Ayvv5WYFW1mcHDPOOQ6a
FrNgf8bAUaKXs1nQkxAIdHvK98dtK+Dpfc+5kkA5vBiMboHdVDrY/+UUaP5Vh4X1
RY2O9MenRGk7df6gMEoScVk5i9xeIPNPlnn1sZfUgQJ4jiP4fkq0sUrVWbY8IKuU
RRuGQrPeLNW1uagcJ0qgIp6adOYaC07mHLZjdka8vQX+wg4atApjncUHuufGe7h2
KEH5PnAdAgIHbPLIMqtiUuZPxeiht6wkio2+RzFc0tspdF8sudpOogSA2mC8fM4k
nHX5WNh4+g/tKlPr0eJlz8US3Mjli146UW9Z5z7h6k+pR+nJK1owPHaoKrl+bI/p
PbOROcUNltjpd/M2F53a+KwRlFHVhNaBsZRU8TOOkgVo5wA/mVDzaZWA7SCfv6IB
NfT0ekY19OgT8x7F4MxoZ9UX4iezgcS2won6K+WWe3uhveQ1MWzE7/9ATAgMvsT7
WvIKi+TUb0J9ZFjYNIbg20yvgA1D2KXFm64PnRWZGhIzh+2FFAoLQx+7qAs/GjMe
FEbWCaw0C1o5XIHYOTQ9aYOo7DeAYD8PN2PV7LRnzuAD2vD/7JiJWQheHGLq2PgX
9VdKR5ab+zo1T600cYGxddDzdx8vBkixCOyYbvr1fW6HIr9O0XzmX9r3bM2Ml3Qc
cdrfWB1DsmJOvnuW26GkS//jg/hXJszxm0Mxcb0+ZxTbDBHt1IojIVJaeUYVgjpG
NDK4G/Rpymixul9mrGEXAFIe4jRGJefz0jlUyEt/bJPyanjEF2MzdjQJmM9L1cFK
t6QMhbLekTCLsEx/USb0VHNnN2TfQnSctHCNr8sybcA3/FTZLJ2+aIoSiNWdBJtD
k4LueFyI/Kho8zXvOmV5i0pcstfiNEaitUxk3ZMMBU1xWOrKXKUR8DKykkhm2W/G
wuCq4EOxru4xldb6T07TiTFJatIY/gI4Ln6O9xRQFa17dwbgGSmZvLQxOvIsACoZ
pOefuaD30oRdkoJtGrcD80i4LAJfQ4/VSDXSDFF3yor+DUywRsbvJerV3CDohi0J
RFueJWwSir6yzFajugwCNAuXCuTVV9HX+90lKXY6VolMCgWyXUfTqqZR+pvzXl1Q
96F/TwZdaS7XdgbxrKAS6tSXKwTOJcCFWyut5D3I9Joxn7U1jodwmFghIDyFvoR2
NumIRp4qEQ5XZcHopePLIzzIcqkw+9VfD6Gxspz9AqynnKaPoq0hrb8JipV6zuBh
gDBrLUkEtfKnwBGBG9SdtiqooOhtQDrQs/SNiHcyza7AFFqWf66SAxXhJQdju+z5
KMyDF0ufVcUxlNIcKLwnrWKURwcJe+dnz8qYFkPiS6peCgx+9UIdZ/Lu7SKoX+L5
ji8G+COqKvTbXu8EtHF1pFFFCvti46Win1l5kQOt2ajkbTc45me/FvbVp7UVs0//
vOE6gslecerOtbrk2fyQ0Qv2ZAXKrrnzYYmqoDrYmiprOrCd6DhiylqTM9n2xQvQ
a40cduy/5GwqpNyx1n95H8UO1bmFjM86Zv3itrL/wbYlg2V3lq1eJb5ZQ5IPOcGu
UqCXxJ9R8ROcPJl/vNPBb9gYwgrnRaNeRbWuGKI1JXINjRlKxZNxh/itpvaSCrQt
qykw+JBVvGDTVJzme1jq/+TdAWJ5r0dIzgKNALkOfI+D6WO6sRNTLSspmt4dFb+l
8RnMq04BTKeGNIBK/VBbCjXcms0ib8RZE0d9Ad6L1HeNhEBx98G3Gj5xI6qzOkNn
VwAfNduX1SV2qvSZFZbvivHYTxpQr9S4vHadH4aBLs3bt6gtEcACx+tEc3G9HlZZ
HssXEg3i960UrQCsVXOrB1xOILVXDoIZqdyzcnyLilRi8GYWLDt9BLYWPATIQvp7
VwUU1rSvG3upcA9ezhpHRsoKFj/jmM0xGcbxDcpzBsIE0a8eSUQ4YSjVS9hyJCsL
hbnkaRKjnEZ6nMZrm0WS2NtjPBKhrwxtxhSrn/e5xVEcv33NcJnRfGs4qF8oPKPf
I22VUExbnNNVSWSsjFpJPhgDt9lt3gp4Ra6mdPlLMYNyOHDUUB4ceWhCA98bBIhS
narbhL0wml23P4uYewPbwrVKNuSalE4i/IOnX7rk6qJnbpVN/0vrzAuhxn/zvTwE
VvnGuB2694g0L2QvuqO7KWCy55Q36VuBZUOYeabGNrkjn63zyA7kXuadR/Naa88N
Q1u4NaQdcva9OBHMMJWqKPfLwE9ogZ2KS9QrYrW9dM1hgztVHYPlqlNMFGBdKJkf
U/FApcWL12x2atV4ExNoqWT0cEX4/8HuRQQ6ZiIX9HJBcdsM+UurbHSxvatvDbk8
Uu/oAdYJClPZ3fpsIapPR0ZW+KDBiq5L188QHWzOZj5nwo5nrYcC1xpRZJqcA8yU
npZQO7SwtN2Pb1TSX0akiXKBsqGedL5VHlkgx86g1I8opuNxOeuJ8nhjI2f6abG+
r6HycdAHPJp5hXHxDRtZiDhEjOojBgSOQRpPsEC/d1H4pnksXoCjDqsBdN9UU8Tn
YsqsYR+L7JKcmNECyabGqlzUyS6dk8IZd37mQI7LRfi94A5FHGoEBioSc4JACa/v
Cm2UjUGJrrSnALWWSGE0rC2mU9T+5+NH78jSufOG++inF/2UwkBUYRZUqHrZFKds
VzAJusqwYHqKEPwrs/7JXWmguGiOMDB5qJTkYdlcsLJoJ5m0pXRAyToYbAJhr7va
0jpvehq8S4w908eirye7u76Xho7NcCKjJ1VPmb0pT9pgJMHC9x7MqIcmwGWAyRJU
SGUahqEIAieqDvdoV2GIddZp5FAPfcbmFnNbk8Ujn1WtU5O3xi7j9uIyWTVAcQHe
Tbpzp6SzJbg5K0SBOPqcM3hDaSFZae/IIh+P9dT1D5xaem5HtG2prFHCuA6+v21b
Rn9Y+mH4L0KrGA55U2T84VGJK3qAg9iKMSqmJHdi7mIJo3J9l3Mkd4jfJYO0wkvc
IIvLBSw2XtjVMdh/t6MXIpDsq6Fa7OJWpWnUkFILORa4nkZRDqS0xTwnc5V+mia8
bZ6Tf3IsYDMhgmQBHqKkf1Dt2xne2sI45jEC2/OX3j3ixlWeSnCly4A7xtP3B8VK
01yBYZteBUy5PLhbtXbA8sJEw2eA/UzRCRih8nfj3v6t56oEs24M48whse+zBa7A
UY7supokGr0m2lM+VakvtpKgzk4MipokjyJwrK1NkUv4BYNtaiA3dWY66KilQv7x
uRbVZhSZ4K9G7+PjjWwxndApZXfCO48rYwq8RhFsERolEIiyQiEm5klfxoUlB13Q
hrd0L5KGqGi0koQy+HDIJiDj/fFhdSqvwHOjxjLfjDBiN9mPFrJLtck+yT+suQTT
VruUJ/9TaMtQiKE6hzfwXQ4wG12kNGXNwwMYHuvb3VoqkQjSreWpq4h/DGmdKfy+
8NL6P0hZVMmuzEO0pzx9KhFm+PWKhh98qyCWkt7WnVJtvWu180CjOeea9BTDda9i
5X3vtN/OelOmGG+9J0rOUEjaQo8/VNU0BHR0E/B4PMtMy0ub7d2FYmB0rPnmdyrI
gZrbJi0oRKnXt5Vc04UmuG7ceN0RFe3d1ho2jo0OQVZRVIj1Ecd+sjXWCEqizdlc
slI1Dd3ZJ0vat6csQv11J49BUcVgfIPzUkxfLp7Jq8MI0mGQBZZ2KW9C4aTQvQ7C
0Mv0sSvrQbyrn3mVmVmdfRNXqFq14DSxcXmYRMdcpQ7L00QNFcvD77LGz+ZAbVgN
6XZ44n45CTB3r7E2yED0JCWdZN5b5fNvM4OCOLRKhBnRtqNsEcYJ0g8OddGSEOnK
xqNpNbY+1vt4+V5fpBFzqeiSIodT8JB/ih02dl6uNWeM/ahMr3FxiTlH16vBt8TU
CDXpURBrqFMP4R99bizv81SsqugQUl6gHnQctVxA7dtuS2KTEOZxjHTwV3SsQ1re
AuNih5y5exkbFdm6h3Ijp5I5rM/CVGxVKeFDkJKhHv6b72v7iSWfArouKHiVDh1f
qAgfvQ0k3e7aNt0s59xlzEFLoRcAr2l0eJfYUEseghiHZcYAbtn22x5zhHb9YHbv
YTrLe65xeUMfyEbEUOkEKxyNRJGsHPKiLps8C6guhis0xyv7GaH2svVukB1RlU6d
QCDvESnkLW62DLa3GSGN9Bi1Hu4+UMCkw7DzgeLxtlp7pRBporrrIbxcmQAVoppf
fFnnztXlJhU6NHkuxCjXB87F6VN2J0blq8eu1RGcTn9MwSY5loVFWvEldT/DHkl+
vt6tFajcbi+TO/mv6umlDeXjbw1Dh6isx/16Yac898a61ZCOlA4zL+P0yaTt6jIc
XdBwbF8jsKsQP1L43t4xCanb6tafadfCUD5O5AbkIBOf72dwaE3MVE5YQjGaN1mf
yBB5Kp2mCn7l6LcbNNPf3OdkhUjYZJk2H7oOkJQOxu/UKRbU+4fn7D2Zl17/naia
JWIMAAwGBXu5ta7GNDzLcrUbsEHGhycQ9SCZtxDSoXQydz3P8qpw7sZAo9JxuzHN
xHM8ioSE2emvJfhOl1CUibs6nRGzhaCdgNhcu48Ea36QR6GJYwzFyFjHyGDDErGn
iJxIugnP2wR2QdFh6M7eIuZ+OoKvo4QVLAQdi60Z4OfHn27DOUKZZWH5ffFxfMTy
RbXocHQPhFpV/IOZdvh/YXpGYHquGOIhd7AA5XdDNbcg0RgDuIAw9J082R2n/qNQ
0qcxFK80UmhbZJjdUQ/5Bu4BYm08MNvMmpcm2cdeh6G+cPVRDV/dBxAV1aiO7g0r
vK1DUXtAwviQg+S2FR5Fps32eZfBRfsL9uBD+euEbbf++thvPnnjgm1Rheep735Y
dO4m1bu/nNOJIIY91edt+UfTbqq2TXewIknB1aE4uR86l9AQ1TDlAMrSoC7TSO6w
wEwotaVCsvLi6It3NuoSOjCGQRhhkpy6R1WuZc/Xtytxh0htMFNtcBfs1QEZw4Ad
/cRg6PnCsOPOk1XrGpy2Sdo4nbkkwjatoXCMo8/fZAez+w8H3YmJwOe7m+a7a+us
/Wmx9VnoywF5qFYpa5ksJFulSDyLAqK73CmDlUDu3vE1RsvE9cnCUs7bgTbin0GP
O/HsxEB5uRGg8cgi+mOBfk0iX2xfIT6+t2a6zM1mzmij/sdNLIXSuQDKB+7el2CY
RwPE8IpCDOepUYj5HR+emhnlayFH1f2N0qBWxBD2N+X9Sr2J9r+ZvTyDunPlWq4W
jG0/qi5kdxb2C0zen2dJMyd6I+cIg03WxbDoB6RzLsGON5ItuxoOkRaBwjFa4+7g
4FLy5w60KCx8bMI6lQc40jLip4ucclPSQvWiEc96QCzJ3wuIjxHrf9UieUwmaMcb
2v15YKcYdpsDHFVL3XL3wZXeKZ8aeyIrBsacmFfYNTsl2yIH2/EZD5v7ATYLEfCz
mkVkcrzmnLV3KC6vQTy5LP7ROQRzYIJPOR7N+f+KNHMnJvjiQ3Xhmr4l+WP2tFPw
Y+Dh70O538kks+lM2B2gfMB4yBAUDSlLVZhhFkQ1JnjF6eQn1tIvjtMYothIwNSy
u8VUDijUwmSNUrWtoLWJE+usaGs/N7gyY0xuUhubRzcbHnFaAkFteGspAismf8V6
EmTnpozSUzGkxXwUTm92OWXUkqgxPFONhAk5W+Od9h7g/LyvWVk0A8YUS2F86m9e
km+WwDym/vc+lEbInQgaRmvbGgMoHJec56wI5IduVIj+kDiQ5/P4tDjUl+VV/PpS
jllK2r88N2XQE7SOB3lSUC1IXDjznvGHOVKzkWUQq2N8EeG0yYcdgVCyNEGam/AX
CHAXYo3jjJ+n54KLEC2k7W/0I8odAFXOtmLwI87WugZybm1fT7wmUuVqPjDWQQqZ
KcrOrlf/D9jjbAxx+TAYthIhuE+0kZDJBVLdyIOtzDj1pawo1C0FxU3KNSLMFmDu
/7RD4I/8DUoakS8icsbc9vigsHrypm4+pBmSU+qGCMfygwmAjPUJlx7XaQFUC7yV
LEkDVeix5GNGg6ZnbDdOOhYgmjPFsLDoVrzAGOgpyPyfxNOyFfNjw+neGV/TN0in
niy4Sk/6+mnDlF5VL23rYDkd3UmFbrWogF+ZFvC7C3LA+y8zSlv5cmwVnsW2g4zm
3Rq/gEzyAzRmtM5oNDafpnmax8RZ2vctkvsYTE649xPFYgqHondJYfPEm2X/Eaxu
hx65h0WwXlZ4jopDS/LqNGDxp/+PtrFu4y/BEr2t6xtFUzhFaZLSHxPsZq2zUU+a
Ku65WvtA9lPb7d7aNKjxsTg3BMbEiZcddQcnYLiwQJZJKlMNVVsYxy3TLJEA4v0m
3Uo04k9q6cmu4+7BSrMGVvvBhjdVL44P5PykysmmaSdOzYwMtvQ5P+qed7QqBR8r
3F1ypZgidnULEWJZl+BVfJUpi4fRFz9sIhR7NRGT/FaWrnKrlbiKeUeHzOJ0ArtB
p0UAOE5FIIZ9d74ttZhnqDsLmtb6TlgTHUVQiAEdZQznjbnhrU2/Y4F8PETM4evw
0fbXgSxmO5MUV0SjOqBFkSqk2Hv9RtOjzp6NyoxrQkdVmPOFPC9P5chZdYsKZf17
Xxbcxb+NhzLPElKcf/JE86h6HhWjb7JCwVhvvZJLaIG7DUqrpkKB3jsYXp3U6xBc
6pxT495WxjaRKtyxngFio0jStvcZ0Y06gpbQZeEg6P9bSbWZhVCl/m8CTBNR+LU/
7BLUw4Rn1h1qQ/hVQ+dsGbzl1jRY/kk5cPpjnV5byZQc8Dz3Tnf2/Pr3RGS3QRqq
SXdCLqz0OV7+a2xBhxXNjn6oNX8tTcG7cx0tRzQ+LHHCKIuOh09RxJ4vArvByLEt
5C8EwQZTKeH6Lwy011e+hYRVv+lstDuoZ4FbqPnoEKW+MPyTKlHoKNgkPQyJFOiZ
PCwCQWLqpNphSk0e3CRTnwA8A4lUQN2jc2k++Riuk7tQJLqzVfly6rFF4d7LpSYi
xW6mWRznE0Fa8QS1q9/lKmd+59pj/3TQdlBKLSfIZ4pYrNOei2yYGteDrlMNsOaX
ToKq7xcJ01ohlsvLeeUoQZkLamT0tmhJ+kqCwhPJQbg2n+LywAGAcLyip0xLznIV
CZwk2540cVZTn9feX1t/1ghi8eN4eCL/mVR44Z10oTd6xOEWRQ7oJwfvmt4cpnaf
3jaBoOKsrHgpmr9oYI8RQorbSUpezk6e0TKw06fOPX4hTePWA05yyXUqpIMMjvvG
T2/o9see82irA/4rK9A1hjuNUFLUur3XLL3dLwi6DwjwzJiMIZnBD2V2VcXTE2dL
gecJHWfAg/nI8T3RNJNETupH2zGJDfxXP/MWTFR+jLn+wp20IDMPgPrfMkvMb0m1
Z+1lIQlFEuPqWZwlXy8XSp3N5tFsfVfh2QlWvCd85YnQUWnabdsaXEtSq7pQmf0R
cPYOSglOZI7mONLULcAAvWxRlmO/1Fct4mubcmpPeathm1XAVTZ/wakAulFPy+ov
UZu2htGCd1wlZH1OODrwKTBB6Z9UntPZ4+ZmXG9Cu/+rr41oaJejQq4egB129quy
GGGTQYvBY5A3HP4ZSCyQE4dqNO2KiEDEt425yBy3MiFBYKO43CJpf8WsTzVITHTf
zrh/NRqQc8no3soO6Mii6vLSi9JOn7cN/Y/Fe/z2Y7boT6eamJhgY/sBZTdUBNDB
pxqPvHnkgTEiNmtyq5A3VfArhnSbq8rCvOoagesfks1tqXJVHI37h/3rtYgtJ2fp
VhmTnosep9VPVdJglje8ge7Rw1J/h9m4cJR0njGJ1+wwnBI5ReZXvwagzFAfUrM5
TApupzJ5+kwyIA+FWNWX1NLR+AJLu/+x06i4zQOCbNLco1K45Vzp4hPx3HbA1w3K
+qu645xPuvM/kHXtVXkZFQAUW4LrE+5VBW0hC5BAGuHOlLKaqklZ7yFKm/dV0rxV
1Ow2EFCxAu6BPEwNX3loc/APhSW6IN/72jDzFCCFwJJ0gI5WZCSVvMO9v7/Ib/Pl
sqszXgFNJs3gcUe5JBx9Pc+ih1P3zESM7Jz9MWS7SIpfa3HaPrrzVy4q6Yu2eqmw
rledJLQTnRq1xEda7G2yEB93rdsZv4PsSl8fMrpKioV3q/OK5N+l47ZZ/cUAPrmu
shB6XdUITrQ7zHHQhEdGDzy0fSpgaRozeCHTN8nIJ23yuQS7nMRyLHVa+yb9Ukl+
40GsuB+M47AUrupZplENPwxF6NhdD/BDLy5aErdUSH3rP4CKR7hjgYqjEoEfNRfy
EcKQUKe0+kiO/bAGFfJ1NxHMJmFoQknz9yCwcdLfya1pdUiyJAF2bzuwtdYXf4Z1
efSIcUZaWGopFXQDz9dJE4xFCZNy6BxbOcM7QTgBlg1x3YQ8mHdIROxNPOllaN9B
HYhOujGcnqmncMJbrE9oofk2kg517YH7oqncKY5LpYTJ5V8CZuxgC/RsV6j5zxq9
cVwKOJdOQ2qNK3tPi5WtfkALT/V75HUD/1br3PisNN3KlYbvTZ3XGTxbhVLN2hxP
Xvf6zN01I+Fyt7JRij5jcTTMVVoRBgxFI1T8+n8aP4c4QJygpy8e3SijyykwDWGU
tOA/fvRdrCEZ/m7SRwt/FwzaRgDDUZmBGsj3Y9aSCp1d9W+qp5LQepISfROTMciN
6XT6BoU/4GrKjugnUN2dtHU04kjl0OdrXgjF2UBSopJJWasm31H3ijY1usYuP9jC
TCt3g/TyF12F229WiV1WEGcGaEgwTH3Q+mnrS+x6cueUrXhi5W0UKOIH0F7WvliK
3O0kbpGMxlx6rBFczOvFxkG+O06WkoLHh/fXYvyMIhnxdSA9z6TgTdJiCWJ4M3Sq
i1WJGFIace52EDqdSIESI5s2EqfAxpiBSD8N3fQ5xmJnm6SUJt0Uqxt07J5bVMLB
JAIvXEtNteMio9c0BEwQkmknES7yEL4IPSOp6kPEdSmTOQhVbtIbsLwfTqnda6tM
jb8cu09r5SXHFTLuMUWG3zpW2cX4oZ8hTALwXH4gR5YooZhiyolhmfmBF4eitvWP
xHMsQVUEt+UA7J+R2BK9MZYrIDXrpjaxy5tuImuFvUHr8yY/Juge6Rkz8QGCw6jk
t99toQkXSDLmRLeW8HOvZrO6wj5pCgx/Cl7gmudNXeVymqugDIGPnZGJxRx439I+
GmJMrAvRa9kXgin3Vvqx13k9dibhxK2DOhfXjcz+G4A/r3tWAXY1Zh4Oq2YPTH0a
lB2Sw82X7gn4jLo6jOaRbsxcg3ykL35JcBDVBa3wM3qeuTE7xb6VyWPmA5JsYVlp
s49Y/lN1IqlC0ah1x4NxzjRgduTxw5v1R/vD1p1NSaGHczjZxk3aQ9z/Q+epjkTr
Ktz9O7TdLTCod3IoMn6W2Yqb+ovTdpR+GX3WUPkm9pN092CUE6IT1yLojAxJ+Bhn
ZCns3+MWLHC1bK0PG53MBEKwptc4yR2FXREADzXiVH9WLY59ghBWKW+4jZL17Gzo
qPKVl0QqxrD55XalMXR3mjUcllNUkIjAyq81pzWuNyDvzUay3zn7mLURCqRJqLru
lOXhabYKKFA70qQTvONVSSXckidsMJ31LVfg6npNEn14u7zK5+YXIGsEjZzx5Oh/
X7CHROJiHYOe08Xhcq9EpOCxpA0YIrTgi6U6GcT4C40bzS2weHYX/dNckPR5qV7W
gboavGvhEtI9q69IYTCHS5+uIa9/U7HIZ5LDnVmeMDHd52EIVkTmnfbDsw91tGbA
8o8tVhEES7yk/cUKkmZ1SFPlh/5A6Hwa05BZH+/lKoORtM2vSUde2BoRgfbZRIGF
UFvVV6zEjOniSfX/7e+sYt2/+fgxEEM9I0s6sKBKXWwuP/H+DUiIWbiJaeWrNDky
rs+S6nisIz7gVFzThqKwMGEIfD31j0wPsx5hYOlFG/vGbTZwK9wgNcQ9IjXxOzHU
kryQb4eCPlHrWW+OONMX5ArsrZfpDF8QR1/leqwUJoDLLx83QieXSMpJ7xnag1Ih
4RC6Y1z4CHs+4nftF002UsXJYYLu/ewPOVk+zfusMD8+8WCaxkyikU+j4oqi33xj
y9jcFYzLtDBhaJ+EksivIXtGxWNchF7EgETo0Yf+3jdoxOTWmquvth51G+wqHF5E
d/LvQ+aw6LQgRCUNKvTrIVIYWIKY3CX6384O3izS7YiUwtRH+xDJp24bKgv/3cjY
mEG8pGHMdq7sgWDptX17jAz8NCGTO/JIMki8eDTIV4URfRzL1rC6XBJ8zFzlAZ9a
MWvLKvaJ19xVqbFvM7cd1XMRXIsKvr6GDaZOjOwVGK6F1wJ8Ba5W76dcPlazOOHv
vqjFVnRM2V+Ni2kZQ5k7/tH5qG31taJQwLfW3VxtYfwmKKiEULO60mnTwNMtrzl6
JEpYziQjS+82iYqZq6hEIFB3SPy4Ld9tjFRikfTOw+XVwC68vW0bB8eR+ZwQKAuG
htnhQ5hhk8fpvSYaPtyB8FM1fTqyI/IeaRzav7aEeWpv1qEdpxqasx0L/WNET7/q
j17akXCZgJPzbSZoGH0vkcAiNp+kVyNUYjgcmTaQHfA7PojbZsSAmssCy64iiMkZ
j7il+/yduU4BWIjNjIUF8LjNPo9e614X2zaqFq0O+RVJu7fMWs5dy3myrGvd8x1F
n/X7wyv4wpBgioKh276GiWZCNrmG8G1MtVuWkS3aChT4v00ta0i9Dw6vnPpJtzeP
PhAbRFhpA0AsqN8kIOUdkp7c0uzglEz2UAfEevfbXQ4B/gTxHBg3C8fQqCNOX4de
hDj08SuGP3phjbNsP4iNIiW1JXlRv1LRivU3e/2qNRG99pEksDpMEkIx2X+fJvIe
GSVeTgPpNz5AvP3/tY4i9QJ7tYExGS/ap0V9XZcaY5cc/Coi5Lb1zZJCWVejatrM
Jbc+OPMIzNWJjIEV8Ks6ngRWRI8FN3NNx/xR6FxrVYZ4GJP55O+2nZ317PiAoPg1
ttEh9ga1e1iiqtB0TMCyB6xt124ZyA+8LOYih/rSDiDEXEphQq1RHIznFfloyodz
n+DLqyZLgiD8H/ARWXyb1yGucz2L6eokCPM07doC866DgzHypDh8EnaHmjAkslBa
aO/NvJ8x7tClXGWXYYpLqdey3bd2RG+nyjuxYpUCaWK3WebC6xzVNvAPY847d5xu
rPSvccpM4gd44nwDz7LTYLMwMe6WQA07BX9JgQ8ZfYZynLebEx9lzn0Y+DTPusAs
d3nZWlX9ge+nHTfIVJgEgcyK6pLM56CDi3nsnUBKKrTYjDaUGT7iH0QoFWiShKBr
ev+StFQtgx/CoHM4NTNXMm2YHGE4UQLyUWitPj7tp21EY9HM4gEJehdfJAGwNrd+
9ZFBcpopHjulJ8aOax7/JT8CFy3Bg9k3/LG/UbXn4IMbNVs+Foxtk5nRn+0zmNHU
+n572jRLBqJmNUnj8E7i756SF9BbPz9MElFamfoYd4mj86Vz+OuCzIKj3iM3cSRa
Rd6qzAvo3z/M0w4m5aycNSsZm6KbM5xPqExR7dTSwy4WJezg2xsju1DxdqhS70CN
ctxPr02liJ3FoweA7Mf776iDjVqKlUDtCnyNnMT1cBuiYegJj/yfYbmNEkIlpqyL
d9sxeQFrDwXUKZMFp+zcZtI2uLOwyBrz0G9wcv+2Cz2PYcQlbnm2csvAZxQuIZC4
gMP1eNzxvOxR/LCO8b/+2dmN8pxn4ST2blAi2Wuk6fFPv2pwE2Mw/RY7H2/UB5bb
2uOn+YezcuFZx10IgU4Zv0ChptpiLU0jtgUXTjBUzvZaCvAnKcZ1gXzmsbQhWyvX
SGuqH7AdODDqYpdqYFQwT/Gcc5KG4oFVyr7ePxmARj86j/XjqvXJKcHifNdDlIFt
Muz8RbTvuecmCsV4xi3IrBpE3QLvbrFqXmhZAmzFqNXMiFLL9NNhH6mWbZFOE8we
D6cQsVlWTrLnlwO5tBiXexuIM0b8+tp9Uk10h4KfBZQaTcysrLOjzBtnn/RRXfvI
u4plRyFsp0/8OZpEZWtdbTDfHeRPXlkazaSgtpsMAQ58p2PGiCWUI0JSYJqnOqaT
SDC8E0kVKNJE0xwi9iKESFcZtBXJekC1ifSDfhErF0SWKlpySkz7ht5a2d8o5ZYh
VA7PEYDkLe18onfA+7Cqjr8fIg1WcQBAT9eRCqeBCs6WO7PD7v0tIpwAQ/7/FhoD
JxwmehKTDroAGewUZQTjTpF/lnIx9odN6kn0iAUP3CFyUGxupMQzdUp77YeBTaWo
sPNo3m0eT4eHwKfx7vmqUUFUEryCfiFpKXSwMg2bvuXUFBiYKRMdzYN6AuOrLIOh
gvVjTyYVbwPzw0JONyzSsd5GPTpkI0I+8GfNgjOXjyuSiA+J/0XKj0+b45zL+38D
3rFp8aDinYuIHiY46rsbIevyqzUmUkGFCvKreg+Ro0al5hDIGsgJsn53m2RPvA6i
90kjTs+aehWJn1tVxgMvoY3e++4jgmXKYP1h3YgBnstyktItwf8AUhC/KKwTEpzH
WK8QhTB3fLAK5pDUnJUpAoWoTOAOYgHOqpcKToq9p0Cwp5rccocnFCDnRInr+yKo
038QDQhN5fnTxSZuT/+sRpzIl5QROZDBye8p6H12Jlz4cAxU5HPz1t9iY+ErF6zT
SW5xiaPL/Z9CQnKA4tNtM5+8G9oiLz9RrEk8UE154JvMWqMOvoa3adWts62Pv+ig
INZcnRoFYK43HPsrsyzlDL4gGQFsPNN7EhUDB2X9VB//ZouEcdeEusr/dXOkrUOe
UdEprNU35OoZYKkCcxD5zHI/pNoSn8rRURtnOTkIAyNoSLrlbBpsQtv3BlxCeA/h
vl3NIgxbT+KYZq7gMv/jlEeERqbwiaLwNuU3z6DKXyKRa/GWDxe6qeo+2xjocbGH
GWjepYp69MF1beZ46sOde4rUJ9jwcLS7DEcbQMp2tonMSR46jOLPlBQJswtlNHLQ
ZFusI/84qBgfRg484rmHSCwFDq3JUQ+UupNKUa2TcEK2cXTousGzQDzhqjKzRx0Q
aioA5+/GFj7t/OI/AvJF/GmaEW+TIYcCuKByrMRbIHcdZUqPlGopzFkMoww7LKzy
7rCz/Oa/m2EiiKxBUhNY7lJcpKdDjUsTAYrw13/iRRF6Pu8M/SC4aKqU9YXTrons
+evVuThibOnen8GuidfDNi2VqBPOB+slWjscgDLCW4zXojnf2VrwyQOuc+/AHV6X
t6GvThZ1XgX8ESAvapJc+jGBoKTd4rTiLguL8ABFUvz8gTJArSQrMPMyGr56ZaCR
aEkOZKwLux3AVRD/Z97iKltAWJaFTm3Pt/r///gv5z17LSnowjcBw5Tz0Ikl+Z8K
ErXjvOuF+shv+PeOoAttJ+5xAs7DWoIpxaI/V6hlUZd+GGMc1ySJls6YsPHFudio
tsZ1P1v3Kkl/ko7kZ56bv95UpYa7WbXHfh2OkVPAiQBKCKC7qgZt/Q1W6QsQ+Mra
u+PlGz9kVqRcTp2XNt1L2eJzRQtXSXZj05KwfnP3EDu0yRvDUYIuGXZ5+Df9mjgp
UoWmrBg4fiIYSXBgSXdCSZ6Y597MQrVs5zDzad5KN8zA9qMvvw3MY2hPMASmfZff
dqNpLKf+Fhnq+zLkuTNwGI0ouGn5NlWUIIJfwAcQsgHRqgPVordLoKoZWuMtotWY
6pxV66ssOaHrtkBU6e2+5xKLvy3f+u8eEVLr+8XfnMQoIwfkmoFHD0NdYB3r6DP2
TxVSk8qVpaFgWGIKCw9oRJ21r7OLzuZsjhebJWkCmVPpuFdBvtAHwxbX8qCxKWi5
HHjhiC69IqqQbtAfu9PHk+DuEBeJXSu4oDZIrlSa7Xjs3+1b1dzyxjGYXPgPUkBB
alrfEqMlvpnUh7JNfg7WBeJU/56yFklZBJ10ukqx0GeJ0//AfVHyCC1eTmLEq+Ux
ynmi9HHMp+W2lunSaORb4wISBzcabR8wI/g5tNsv8LZqlzShe9/VND8eVIM/VvxY
ZoroJCJrWpRRTreYMH0yv+vZcenruR1IzTTxkN32v+iaFGKL/tGg4flQKEzlcx4n
6AlQwg9MDsnLqgbkgm8oSXMIYLEL53HjbTbbaTMMeD51T0K2WdwnbpfwzfzS2Jdo
apnD77uQ/cSprfbyAEqWxng85oLsaCZ7l2v8cVwvpqOuY3pD3ukURmo6IqqC/JtQ
aiaYxXofzz8Y8IdqDTvWE3cP2TIrNP1vXcCyViAFrrNHUyZmOpJswqdVT9bK5YFg
aRO+4EETGiRP2O3jqZXYShkVNaIP90Owb28zW75hS660Qvz2swsdL/xwekLz2Yoh
E+gzyHIJFesSWmHY8v+LUOTAmU8aP0p73QaT/l3KK0bekNpP/yI5WxJ9viErrWii
M8DVtk1umekBAwRWM3U7W50cdswzVEEorz9wVtqW9Ehl9Psd/14WRUDlqH3LW/gY
NwuBbQ2QBhDsa+FtCp9fWNnqXGBxC1D9o/aRyw6CB/S2UkDrJfFSyWy4qRLzFOWK
5T873bE+3AL82Bhzwf58Mzo/U0vBDvmwWicqfVJO4uVF6P6x8kbSHwg2VQZp3ZkN
AiW40MKaZ2tnARyRM1mWwbWDRuGIbwgSA6KFLI7kNQVq0JVm1qcJfpSt0Vm3qk/x
qyWKqIGhEYFFnBmoYuO2a0uw8LCjBQdsPr/d6gLvD20/JBm/PPtJ8GuxJm7H3LqY
IYxmnAHyUqlxk6+ddOznAH52D4LM7SA0Ec7ckkVenSmO6a+2vJM3xwqYtrLrylEY
4d6xChUTAHe0u9YbOKyH7DBrmk4eU7tiQ//VjEljwkdSg2rFaArw18KNd7AidXor
IYqUtZWmxWYwDCX/9aMD5r9dPU1so1gU48AmoMKbnKzm+SfpgIYhUio1mWmhBlcS
UekrsgEyHY2Uq0NSMN2PgVdqJFzNOBStyhh8vTBgF2f82DtZrkq83KlxOGUplwj5
9n+ZeO6DfJjDDZx53AotNYyIgcfs37VeWKzuFJ8VT/V58qKyW3cLIoERAaEdU0d0
P1q43DwvO03wYR79wj0JLW/aYIAMoyu8F20a5UkqqCPPEEfBBt77+sk8hfwVoFoC
dYa4pYVBFHf8uEcV5vwsEU5pBKBLaI5cyIonVl6cEJXjMLAKYPalLTP5bnkf3dgG
9hgo/nZqwwl+bAjkHg0TKivU3EzZjLxf+ai4I0KG16T+k1oos6XRTzZOJ5y5oDi8
3VRo+/0RsNlVGhPKKfvqXZJlueLX2IZXyN7pWGwORDJLboT/yp3vShyXpdD7P0Pq
2VykFp2Vr2IZv0hx/ESlW0vmdgwoA2zwIim/eBhduNBwS98+kjM9N6TA4qHnj6y+
dAFbJM8J8jD0Qh2dwAGiCji4lqVx0vMPmd+bzXmhyQpPTu3tSI6OHUWiaYJhH58w
zhfTwEVau6iqxFKOSuURf80Vxl5SyAgaUXBV7oBN4byGfTncIbvhc09Gz3uEhLZ3
lKGwA31uius2va0EDmEsXF7kELDMS+FYBMWgiXo4MwYQkYU9ZnYIfTNAhUtGEAXx
8jNHJsQ1r1+kAGuGDKPyuwljnBuho19HrQtNf9Q5bjd8/6NvhpnzUgwJmwVuptkr
+0Sm7MIK8TXDeh+FvzEQK4Vh4SJMU/ZNtBs39ZSp6OBH1jbsv3nXnyEhtWb1W0g2
fbxEGX9lohz+dViu4ZfVYC5mrOM7hmF9zd9CG3jr2F21WfFP6qYsG4m7ylVbzzRp
0ZTi96pEQYI8FLf4utgLJx9VOG3UlJ9UH3jNk1chYb2qXCR38jLXjk37GOB/NZnK
pQGoCEwFXn825jIVokt9cCqbMvKEc0RGsDbHR939KcVDlhJ1S/m1mIajd/LwTIt+
mwspqGW2HQG4XsBF2oXGwiQwHr/5YTU9Hz1ywM4sLIe4fFnKtmiciT2z0BAj4Fjr
8Vt/GWJtrgzlxs2+UiWbikVk1IXkig7mbZOH/mWCdGjoq9RPYiqISYp8oOoyaf5U
wNpvTKt8blCKrgDZ/x0JWroklmXaomLMRMIa84zwHjfOzEc8zcgJis0oZSps1qyX
aUh2Vj/3Epydhr5T1BNduMfm7YhgB5wnTAcN01AleKOluXkNciC0poQ5qqMbYGoB
RyP/441uovP23hGsSaKuoevgd80y8CeEHSdLSmP33X3FC3xxJ+kO6CScu4quLFyB
4k/tANCXb80JXFfdZs5HgwUnOsS3WvnXCBte6gEA0Mvmgmrve4pHZNWvBF2sJkOD
MisL/WTyTr3QskKkmiEk8JIJdtyp3EDlj+5hpy4NDVe2pJLJQZAwzRhEd7azXrzU
ioDWZPsEYKCduCPAgXhkahi7qMx7vQwxln4gxDBOK9+y6QmiuTx7NDNUxsU/10sb
BnYLTxV3/HdsI/tjyjLW61VYYlUK7WhvtULGKqnQh4M7ta9uk5QWe2d382LmQFkl
C8PO5WPwjvofnZvyTnuudxcw/HMfca00W5sw6Jsvzkk/bxvHsLR+9LEQ2UCJyqnZ
kYBaJCQVCM+d65GoDuOpkqQrzTvasOvL92gsYnGw1qabsRTrga/Wr41itJkV5DyA
7E5FCQpMvm0rXn3EJsfcySVKhBm6EJ6tipbJ28fmipp3TY9SWPJ5bMbmF9xRAB88
ihMOtTChAzIEOqm15oY7uOK3Mt6Ux085wmrGXndfrRdpKmjeNMZBXdxIpGc/0uUc
SRDjaS+3VfWxEYxSXB3dtv36aP3DqIGYLvU7KpHB4HicTCqpn86YvX7K5l8YJeJP
qcKXIhK5i+ynfyZRslfzz3pD3aEnY8J3Di8rOWrIpTSoINVELowbgdxxA7Ay8IkU
b6b79rUzZvvQhyvwnEk4eGi2AoeDM+d/DHDH2RCjIiaARJLMiCpnu+TiXpXdQpKY
gkr0TNYkD3a8tIUq97l2wzj+nfyRGhWmRroxX0CnHwDQg4XONv87SgFWFhInwiIK
1RJR8yXiw3HjdYr6LsfRp7QXiM6d2e2PYwV02W7XhPmhOH5gWYwJrpHVLojeERGA
MqGK0kPB2+5S11k8aW3CrknJZn0eergg+f3J6ag3+k82fNhBaZ27zGySlmzc5ATw
0IK3mFwQyI4MB6uIRiljqOFqC9c4J9UdmjiGYulIgRpVzpkcZw2IrKgkBTNA7WW9
A9eTrj+zvRAXIw5pphMEpjIUy6DDhmWQ7k8BUdcY9DiZMDlgoMYIdnF4sse/iD1a
ME6XWmRpJtyfwfG9zWTrXnm07i6F1zeplYZWYllpaT2//LluFIoQ2Jk5gi2hDPio
BVhmPkcCGpYo+N0R/LMgg42C7SGPbMmouBaNfSznyXymCJsPpoaABq2imBFNdqUo
fJ6oqB8lla09ZRR6acdaUg5zlMfxOCkcL+BEGMx0sLAvRoa/ZLnKydshQy0UpOpV
hhS9WbDgv6Vbz623kUv9kCrM9u9BX9frLFEZ9o9RJq2FS3XM1NnL5Gi8/321mHNG
oxY0OE0q4lRPSvSxYKUT9LjFe8Kz4cjqXM8pboZUFY0Fw8m49m07aEjoOlG1Caz/
i2szTAoQaCn3tkQImJk6a/aV9PcFmui6ErIGYuS4QY5qcjikl+AlQqT/uCUFkoBY
oDYUurT2+0hh9hdUvavRkAwZRRpLDBIKB7mx7/+OmHSNBbkAsy6HJ53jvFk+7Xr3
4CqptanhNcK+dM9c+JREmMVuPvhQpfTn592wA79IVO700iMYwr0rPwHqo9Y/A4QJ
OcciA7PVtDtmxFiM0ZXAASw6CPyhmfQyCKZV5DPZ/5VhAMMNgMON/DMClUBTw4K7
68/wNDjSKxI+Prh8Gx7gSN1aDQMb9MQp774H09neVjYBSsZ3jDYfjjRBifpH2FQY
B0ZwIoUozilkMO3e2idkddWT+PH5l5q6k0gfs2BWQ17sQydqICxi3C1STHsAxCr5
OCoP9javuKHCN+4YMW9XpVpOTXsc+p4QI+xQNWbbgKWaTFiq3fp45p5/kMoGQ1Z/
I+vBqBDvpEqRK7aNWO2SkC1JT+eIpe/f4CfaqA6FwRJ1CjE8NZHcYC3dzDNpVIwR
Bqt6xkVPbsbZQ8UeMI3YaeLWrzxmtUxaKlnP4ClvuLw36ZpFXetv2qKcnWS2zA28
AkSuXQYfGR1xuVtB2rrqCQQTedjJEUroTqyZWSC1aZRG3I0su+BP69ClwaIWz+h5
teiSXb20q7/B5HItnkIjLzQV/hYLcz5ZloIyXYAyGD9VgSPABdKx3H3zMH3yNCa1
82rNR3E6jOuKeXd3Ntlwo4w1wR/J2OKB5WfkKzpPTKxyvmOq60GTxX1y3oFJruSU
WW63lFAtgv4ALKzieKEftvatZtBXAAa2UDslkKuUITl3BEGl7/jSNwAt+5nAUYkG
5+02n3VdZOMSXvOgmx6T509b2LwZm2MpKHfkUYD5CX+aYOeFrM9/TXaN6wAgjX2H
NU6aCQKPVCY0pYurRwPys8Ovow38B3EXdeutLQNN5xuJHdp4idIR8syZl5QBA1dw
iQcOTKa1zt0pTk0HPx+Vq/jaZiZw4V4BqiQdw6Ws8RP51tAB40vQH/7nr0Jwjzc4
LT8/2roz84/2271vuUVZshNy8Dnd0uE2DCnMCN9ZiuvcLymY0kzms+/qahRNkKps
7LvMJnblxlP1rhyQuu7Eo7A+XXLUwPF3n8kj2CAaeUsVCjc/hDtpuAAQt16J8QAx
OfhJTi8zevwpstjWn4RxDvGYfn095wrxynitTbSP/LQvN04k3vgixql2hctmCti2
pMBjKFfnXdviXTE51HrhC09jCSGhZj6RNd5ItjKKSEd33jzy+s6amW8jQ8W7HPzR
HCKRZrPpGgKsa5JYxuA6YjyuMdp/zFmsKgmy0/PPrW/vVD722q2FSBLSq7WLCHTU
sqUsf6Bca1bPyCuLkxcH+tkz0JA3MPVWMmZSgLJIJYkd6HS0LwuonhZsjIXmC5L1
G/E0Ne6kn7RtC33GLuhun5eCCAWjHU6OoyX3ue+A1FHy+W4WF4iHwPLS4Fg1Obkm
fsX2qE9AEh63VM8kdcWW96iMsnM+MlfRRwRrH09QELD4L52LCrmBAwFu5W+z4aR4
qZ3+otEWUo7jjlB8durMMwOfaOAKjSdIlFBQJCQKVVhKpw7pFHHijeOc5C1UyUxt
ckCZH4ST+vEDg1I2RcI9vK4SRwEWkG2VkYIPLGO40uZB14XfwdJk42nQVvjb2oHV
+O7rD0ZM6ouAJ8IrbfgMyS+vOkzVMOHmG+Ns/oLm5zXRAeNxtyHkgolvpN4aPne3
dZtI04M3+l+wcvG21aQlbPEXS00co1CELp+dplFpUE9qe6R4PT5zBZqBKXYzmjmt
wedn/Ts2pBH0bdmWZKxIuWYSVFaEqokh3quYFP6Se/6eqTNY7i52dFWUTpB61hWL
bpqGbm5B9GIbSslKf5wPyy7ZGSYN8J6K8F6/RObr6R4/g93rqn+rsXA5ogU6Sc1y
zrQjg1FDd0Grv/93fzwCD7B8uEUT2VezqTdA53GoBEJuqEq3rki9g0Ul9LTJfijv
nFOdx70ftNtn/q18/KAT213OB6h3kcuL72/5NZ9/g8JpEIHvW9SFJQDFR59Igp/5
O6lQUo5qb4KI9mZ+Je0S3vnJjL+0v9CYl4a+xka96S8fgekSCD+h7TDuh039Fr0W
kNYrG/nKO/lEPlQL0JGn2eqT5piS163It0vb04ITxSZe+1dsLFaDBmBblYEdrRXK
bpQIaL2J409yWj+tlsD3VSZ5E3FqqXYaKc/08zgv6X3JEIW/ROuyR7zeO6yZ3akR
EwR++tt5mvpOsH+2PArGrhbh8ga63WCRa3gHBMIdg9H4GS9IOaEZjqxqFe25hjU7
skIUZMI52yeOiEOht3uC5BcnTIQTPe9UNVtMaKADbU5mwB00f5x5t5WBAmfzziJ0
PTSEiU8ezEtcMLlSibEfk/9omsrw+L/8EcYMVm0XuoXtkdRlzy2rctV+L8k81oV1
FP1SxFY7omHC9dho8z5Rm+VjNOPJnMQpwr8nCTEHUyEhfTFF5I19E4jAhY5IRe1q
VpS9rMBWP2eA1xo/yFuWY9WDl97OO5YRtBEmuF/06FIQlGjNMd/klbAiBgpk0s7k
RWJ8CZVOt634U2ZPZhLLI6KzYo/7BkJP0PkRG13GpWyUMrniRpkF5omnFid+HAdN
xZ4eM146OT0NEq4YxZwnStnEU4G5+rYTT/oK/XpjRM7rvmXP8iN5oE6ojnrp2/do
Kc8qJgHTTip6PKSydkTg8HUm8CrtCO1I7ixVQnrpWxmFUsM+eVlIKFZujisjkZSj
B2DzJlZlFdGV5DBxT+07QuOizdAGD6+M5KTocX4Y4XngbNUn/5oT3WrDX4iEwTxJ
DcTklnV+6V8Ns2AmFmfbe5FgpqlJgQwvPMFrubwHmAnce2lfeZ4nNgXqEh1oB53Y
iL+oxIl4Hle/2wkkdXbnYgdUDkrzTjmZaOzpZkf5c+cnLb4fcR3hMez4+XWAX1/m
yLhtUXzOwm29ONGcGKim8mNk8GMwRgFP2ZP3t2JTXIzLTtkNiSBJYj9Ls1FUSE7G
GMz9XJDqQtiImSwUsDn0rFiE4ohteEKrlatwo5EGSLOFkI9VxbJxo4eo8fs9/aYr
c8USn3Svi6Kca/JbEK9AbFWfhCkIVrzf7ANI0rFTwbKj5+27jB3RsOAUe93S6Fvz
MKNLQIKlqsluieUgFJtDLzKFjIYlK6dfqLGS108lItt0FbEruiNyfJ76K2+KXUxK
TNuD+evMI8ffBqGLNNiboyjVevfh+BpSq9JmwKKSAaK2lT9cJME/rIpiMbj+ni1v
xub/cvhRrotokXeLizPQPu1CRmg3BSwauI1LHkmCm5JwetMLW1eJdAc6oXK2GSJZ
U78AkoVaU5gXY7z2BMw2yfBxRaT6UIEzjbTeOYLx9pqv9Kc8tLYVBzdvTUDgrS/h
bBTSwoHwohj5QG6l3dDwrhQgvYYGiP4a3D0K97/L9yZFQ7QHV2K5UbET7vJntCX8
4DkxESJjke8CybENMIjk2OwL/LLRPIUAIlIf24By22Cau7uCkAZ/lFmM3fCWQNKv
7wNuMNy4A0KNnzx0oVgH7XiRvLSxpLlq5WIp6yGsPjqG1SPA1eIuKTzAfkdsXxCo
PUFXXdDXiSJR8qFCeVVV+X/6jvV9BfTJH60YbGKpY4aAWIyk7UdArGu73x7KfZSf
KOUXByXChvfUJ572Hup6mWY8wBWcCT1VdFOCkFNj8dCSg63Wym9hMyoQckTrVUNb
+uuGnKcHI3+oP6rEvCi1lqmjtqB80QHOVlUSrgU8zah9Yq+Fdb0QKz3BJIcZDBId
azeN6eiBmW6rkKoDZHNzbaLR5UKXb1lPxDWStWp8k72ts3a3HsOJiMvyIFuBvsEe
kv97iwkY7tTJq93Nl4dVNN8PoRBH8xfQWLqxINd7pxM6BL2K9ykiQaxvszZ55JVf
S0B0XuLLDgRF5ykDorsqgB1AmXeEZRsPfrhAjaFcuUaMBH891+MkcTrBU1ptEBjv
VJQ9XDvrViu3RSVezvPzi4/k7zvEWKzVuqoTx4QMK+D4gPU6tk+3Do1opyaCuy20
oasSA9rdxhUHUNsc2/0gZWvn8N+s3DbJUHUMyBhcdKXbwmiPmsaHp+PWsAl7lHbq
aUjkaz0Iqo9OyzPc7kcrsB+iUveY5USUjeVbqkAd4VVH4s3ClaeehoD+Ur+bdErY
HWyxVoHqAPywlHtxqvTE+Q2Oe3IjIHGscHxbPzcPkI8vNxJJdqpFGsRIFMiRI8G3
xh0sAVEr4lO72PPM8huuXV87/TgqsY2JBEobxm855tpWlH/mifh3RguDSnfVj0KU
nnVBA5ZBM97ShoYx/KlyRSD7pp87zkXru+gC4hudKQgTmLB1uKoDPPRLZ8QqjsUR
xBEvq5C26bVnU06BfZEliUQBS854uV9vQMXc2JHuwGLf+mPbpy4uOXLVj18TO7k+
auS4HoMnl55MNvGubIk0usi+jf8yLN5/9rEGQNSjBc6JlKl3nBnPgWqx5HROFKby
hzvvw8yPEEUjlE+K9ECYV+IvUWCEiXFPiosecEl8yMcjdDpf2eaRhIl/2EG8XE0w
7kn6g1IdKSolhzGoGiWLzx3qZMMmTCsvhQ+WS3dMQvAMZ17lwx49C7adhJk+ybzf
I3xXcYlYZUj/uEhIFV7JZWkirCcdsmBkgW5JRJDyWidKcQ1hqzwmtFNyGiNOTkuQ
Jmz+UdEPLm0mBdHBJFNy3+6Pk6w0ehrynfjZkjOLlMCYzTa7mrtxpAjxOXtCOC/x
uDS7PhgupgBBohikAOukw2KmZ+doo0f8PCWGfIMk13vGBZcrhNlyDvr00But4jLD
8E+ehFBPy5+l9AGtDeCdOQQWVoaOKRQatdm/nPaEUhtir+5cgYWeIebrLqpSz7vE
eb2YvcGGtOYA5+OnQdOSbQD2gM8x1TvxrbBGgZ6UpQ3tTwa3zNj4tz41hgDg0gdQ
inlbEgxk2AZcxMHcVO3Aag0g2fAHiCHHtQaNsQUisdylYOvQ1SavzKiQsU0yFJjm
cF9mX/YiqUNRG/1qM9uwB36eM+Ren2q45R+Gu39ijpu01gY2jhW45PQpYtFmqfJX
eyv4EZ46EHwl/Xd2pGnbOzNOHMIsPCfR+/Eqd1a6rxycpb0nP+9AQ/mpHZfzfi4t
yzx3iV1Q95uG2zhibLT2ta5M+Qv0K/F85DnHoTsXLyCiq47rg/LP5QscphLtZXAe
YCRIs/Rff1yKgfq22wYtRFlu3T3D1lQ96ASxZiAkHPCusNpGjqalZw+aud5wnK2X
dhtQ0W4j07tgB4T/qHHxzcJs0bY34Ekc7hptYG1zBxaF10cTVD9Xw6CXP9ZutC4U
DRKl1zNmgjKOjRFQLoVXrpndvm+tr/KCqSn5Z5HQ4O1VRebpUrWkX+SXjFPewkkj
Iqjg8WTNHxZqZuiV5vtTKfRHaVAZVYlYXzGi8SkrZkKQ12gULYS5V1rVg8ys3P+X
8syO2+jl4n+0tKZTIqpd/exi/YDTUmTHTDu58H3BvYRiOz+HExtPQKBTdHjIhJi0
Etf/4c5iTkYXEexNbdLv5EZ/T7qma5qIIdqzk859UQKIP4iroSV2ECkhmZxXD2bu
z4rIqLb658CaEanOzDMetFKw3VAB/7deu7SE0Lt4b6ydP81I+LvE8AF5AIX+kDJ6
p/IUxn3rop+yUHaGKB/+H2GDCxjdRSx999e5zE54PVwEcidy5ewavgWJxlW0DHzk
iK3ZW9I9kITLfQRT15uYyr2Yc/b94OcsLIevS3zp4MXoaaIgbhd9RL4iz65gnUef
nJ/sVuoEqdxdJuFvlCnF+mxVZo+vYoZEJyggMXPiotv/UURlaL+rZLChNE7PgGrz
2cwS5S53hePgFIqwUWU+BlaMTPe1VJu+2wizi5OH7y/7gJqdRL05TiQ6gZY8i9hA
zFx7G1GOlssLeflk8glQVvKRGE45BRArXN3mbQHEQkl/9R5KJUCj9aXiDK9vDHzA
Q1hkFuAGYr5YQy2kArBB7XdkoQVbBPrxrm4kyjiWqFTebVlZ9zoJ0GXvJDbfM+T9
DJpksJBTqZu8H63Va63L/A7aLehuGY2k3usWZUDELGZRkP29hAbQPPO5BuLunkBX
wVH9L9J8Qb3qL8tT7Xvm/dOqkJWdGYGRFMkeIdv5cf8AyhwbAIDQxsFCNLmyvuLe
l6HLL+DTADF5yfj51qVE4l7eoMO1tBTYuNMNsyYzvl9mT/M3j0pmzwZql7dFpKv4
kBEwAT/vIrV/eFoOQk9nHQxqnOQaPKl40JQmmZcXzNt3GAfYoJq2Y9kgcPjdMzXt
aTl8VxO1dBQRBbHQT9Pte2hGlmRlmjI/NsVoxUp09UfAsCSviAHwVMZSvkoBOxol
MdJnjMPXu8VQgKNKhrRslGGFACcZev+EqO+SrwqoV6KcU1lfEVdJmDrkWTV/jbmP
y2XmclWLfqOeSChENZdRKrN6sXGxgIwXjKP1mqT6LejoesLS0OUNK4m0sc8X9aF/
Va3WKf1aeGsjnvZhRdP/jr2z6zPDc/NmK6FmVEqF+LWT9KEY/2i7K1tyFuEk2cL6
Ib7Il7oKKZvuq5i+ys9+6rwZMog+whoodtkCMjaOJb7Cj7jLL/sJ0QhSEGwbI6Gf
txBXN1m0FkDNLXYTbONAiY1ee3C0oQyxRkZQY3Kw/3LGJN0cbJcaLlFoyN7SdjEH
UQiGvkWVgiyKr+mN4qchFG6k1FytHpgDw7JKtkO9HJ7x2fVkzMMjEbbRH+fIHwxQ
6qaTlxen+PK9xuyjtXa5ZarHQA9uSRW3dzVLmXDJsKytUNMvRsncar8l+PXv5qIz
OJjwmg9k8Zn63P1UboE4d/Um7VVn7gBdqf5pKF0IOMv2lMY1Nkog9F+EiqRzpip7
r6rbk5qkx+gVyzsBnL9tXZceShsmICnNpaj+vdFBPiFXFVWkCSjWVZzZSV7kzv8h
o5qTT83FlAUVCYsB1v0RsWuZeuvjCRWBa/6J3DvxPli8NPE+TfeuCiokCkWApTPG
V0ipM8cpBGjeeve/OVcOz0ScPsZZX/7/ipiNN2FZLx194T/hwGErnpcrpIhp40Sg
m4mPf3y2DcU5VuZcL13XbD5EKPbcsGxzB1iUiT0Tpvns9ZKYSG6e3Rr0omJxHhPy
DcWjKD5QvZHOSBNhYCYdbjAh0ROpaLq+57xVENgFor01FiVWNuC9Yepy4T5FUB2z
KuFXoP0ky22VsBGn9aovnxvv3eAqHQJ6Cv82+8iWD6CBMsMRnf3H4BgQaW4kNNJn
vran1IyGJ1m3IzTtu5kfBeHZiN/i1oNEQrYCcqSIEbXc6c/LwImwQolbb6As9nBE
7cvpG6muK0k8j0x1WxbrclMeZmdER9S7ZVQbtLdtkaThn+SwjDVBVsjNziSY+GNH
KhNVBkGC9QS9hWUvcT5VHaF3dF9pQBswxLy/PiYNgOeFingEjdTurWrepSorQkOR
9Ua9+P2FqS7Gv9UgNt3a0emvotSnHCKFQPFU4ySr3YB0u6t2BwQ+CcPcs6LsBtuC
qWdcmeNZl9KWXrpcndm+exOeZZ0WL74RMrGYQONntyPw71PHLmnIqO3EXvJpn3oE
GYH0IV3FrpDXV1uFQUg/W6FNE6Rz5iPFXYhAMSAN/6L7Zbith7WCzPg4rEe8mnni
j27bmtBUiT6XZZkKXNQ2Faul8DrKg5vjO9NiynGo2hlEQBGSz1xTe5thFmjtXmQa
zOXe5lX/zsd9sj5kqLudjyvsYId0JNLrS+hBBDcSJuENiDoGB0NV4iSUrekiY1zt
eWh8oGEEEgE7djLRHt0zpQwR48ENga9L1K/h79Fa0WuxxlZxXLR4DjeWZr1PAd6t
eSMTIjuE8JiUD0BmQphx2GFcOQeQF4GiRyA7cTk4WTtLEUh0Nx3+P40T6UZtszn5
KsT7eWcAbLons509Tfhcg0U0CBRK6fdSRSvKCILbgny2F7i8ArTXswTg6/FYRt6u
FAe7SRkxbG7czAbUOhRSuys/UjdzGoVPy+lO4IlUFTNJfTZvURSxdFgf941DQNOy
mK2wxHr44HM06WYaHEHQbMRGCQRPLhHv7TJKSmoVywNlRrNAG3gCTsw1ZWcN2WSU
bh9e4ZEle/cfISUO8haKwmxzNL4ubPOq0cCXAE7t5mE/i2iWm1MAPQz80aSshrgr
vWsD/IqLMXXfsqaobwoLgOpEPPE0Sv5pt3P1yPZpM5MN7Fk0nygfK1X7s7xPvb8c
z7yajpZ2MQdA1kjsbB97L0Iq1a1BMrSGzqXE1WXUAtc9Qr2JfuQhcTVVu5533g1S
s52L7YZVSCWM7vOPe55Xg2yVbsrXSLzAOLhKAJESlHS4DHdvSx+zJhzatMiEWATN
g/SNdKF+QA5DpUY/xUx7NN/1TaAnb1sSR6VYVWJdKvvWwhXZz52ZAvatUONC1ZyL
i3H990UDc8eZPQ7ulwDuiKU6IGzsUh7MYWNdi7sQhmL7Cp10Y8OchwRnaNzYOoyz
DoCU1rKpGy8/7sarb3YG9mISW+TtetkXb1HxWpLy+Z2EDPLRKmLWfvx2kpTOK1r0
DUcdJTY6ngoVEVS8ec0+EiUS2k0hUIDmbjnGvuM29aDqNXDoXscPOezMGD9tc7Q9
ZeOnaMn3IWdSF1JP9fsdftQchBrKCTr721fRzqw1mQPIJh9Re3Yiw6g9cUB0T9xC
rwyYabpniv1hhC7NcJ7mkhgbLX5Aaugwbfl8ygtZAqe6PZ0WVRpNtvOkr8XCTWfU
ujILsjuNTX960MeWn9LpJDgltR8E/iK9Po/dXJVfB82XRAGQcNxSjwQkUpsBbGXk
n7Xg1R9aQ1HAqVXXc/SZ1xEd0q0p8zi+cokRhU+wvoiV35I3CDd7PJUL8SatT9NR
IKKSJB7yMjscRUsum5xYpQLYRLKFOD6gK9yx2YHowRN4sRDudGInG8XiyJqCwmvG
TQ806C5JNy9TTq0X44h5tH9HwNwPszHXVSjSZNY3u6+alO9eCWvMimlgZyXTo7zm
LIt5gOwE2yJHyD+6x4D921NylUpfhYN8WYHU7CaKf3WvB4BxXtOTWGRdOaa9+akZ
m9gXeXQRjAUOsB+aLk8AHp8AOzUazmSCGbnv9W74KAriNhvwhhaMh/8ddfFqHBDW
7y4B/z+HK7i9Cd+D9pcdzP/VuPgeLQCuPo/ZXEqTL95zSGECaJKNAzjjkWoKUQBd
y2x1k7C/tOMWl7xjys5Ur4No8qsp7aoDlmHQXua6+4Df8zAQqj+6fXtKaxKYXAWF
TpMpofNUwQu3e+qqwLaeI9wtuHN0RvHDjlEvk1tG21/fNDsc6SnutbSumlD6Wiq+
FiiityYzVbAkLjqxYAVhyNsN9uioiqt0gfdu5OhKCS3we060ili4caD/+aDXCNkh
IwXI5w/rnLYxEll5QtkMwNckI5mrr/mTkoSy7PYKFbZpHioUpclPmLGDDaZHzNxn
ANxxjQi+Ck5f6h4QiCz82YrCTNctt7u+2Y6lUGbB6q8t9JQIA07vEZ8xGm9SRzDE
9mfL2q8HPBr5noGQ6cxT25s5ANaNp9tD0qt7IqUKNsSzRchpwBAueioXvBhGhL1a
1TgACkYWJkrijIg2OzFs4SKAvbDa+zaYfJV10WkF/lTlHJC6rGaCUNXn4d8DBeHG
DeJ2sgFq01+Tq7mfVNq97YkOGlmO0LLl4mdScf3las0GVDzxGFb5VnaNA9Yb0A42
8bsqdCEksGkkS02tslvTamXCaW8YNktAtHxjO2E85KHuIEIBNRBHAM4Xl3sooWz7
m1N269EjsMcyxxIhXRPkQ+r3ccoESgOODKik3Glgy/cWhY1Z/YeXolDIGRM3Ion4
aVedEC35AGIQSfth1FPO3didnPlKhtwwVdqs+VWvD0AGHesVsp3BNJY3YWIhRVZh
uFMQWSeXGphE7kUnpDcdlb60EER8b64UXvKdubVPt3fThkhdpPqn2lx0sTlki0S9
VpkPAwpg8nc7Bz7ud48nJ59/DYg9O6UkRtYIuPwTBU+ZMMZc41TGULAQ0xeSGr3D
6SHU2m8z4gEitodHyHzAl19bOgDs86mw0g8k5b7iHHm4TXRpqIMIZkBPhDATWWBC
MiSxghKYfLf5lH17Fp934Vm9jvojda7vQ1YzkSMEFEsvpO2fYe5JNIUbolwvVsYS
i7QB0UHp7cbnewqvQEVnUoiZ+YoJtMTnpkTPOU+ntCgY2GdAaI+rnl2/pa1sxFIi
GI+xMubDc1czMczHI3Pm3sKnOOw6UetWeq+b75tJdRGAg/OcI301Q1DAYSwn//l4
wjrsuCS8v9g6iW+KArSRGG7QgidzH9n4MyTexrxU5EoqxqLUmikP9qrru9KHsL93
Uf4PjZCsTuG8tNgkTktl/77kssf2EHyMYB4yBwMF2R7nXJoTFTmfzS2S7FnGozbb
JQUXKhmY7vSfDbGPmGrJ5FgY3OZM3EHWDPKHxzdntJa97958M/JTswLS4U9km58P
LyAmwArJgj4RwvkGBka4w/CM0tk1qmPEXfFwvfWASRe/v0SIjgJB9bm0aRhIbxWN
Bs1YjiTlUUJWlKODsycKPYb1EA0H7h7MaWcYk/kIq3y5fvRHH1wgtKnmchAx/vid
ZfzTrX2NWbpSHjo/CLkvdLGspoCtaJS4WxbXwhqtjpSS5vj9z9WmDaNxvU9AmO2C
Rx6XeFvfejcr1jZJ1eXnJVwsjI2vH67eTkr1ZxZUXLbh2Dkz8Q8HrdJcfL/HNP3R
t7fjPDr2Kb950VIaZxNGQ3NWH1JjbJoewCLgLd51t8fAherR5jFOQvII6vnFjU5w
m6TL2YVaCUPfaFZCsv5YMETwMzXFAyFyG+rEGgvdZ2esBbyvTMO+C+qoZ9iW3ZUD
kS3J/jwWzX1YFr4p38tWSW9KPENUvjo3PqWXhejw9wlraDm+UYFgiOSlhQ0KuSKn
gGFNeMmBWt+FI2wmg6kdR5TsS+SgGIWhdaQpU9j93V8eUBa05VMdEVz3vWGuUQxl
+uyX1id5lblCiGqhYiuD14M9JCSrpNHNmJ4vUQ6eSX6uK4yTHy5G3MWvpUXxd7Ct
G01iJaW7od9NVLvOQCGcRoZkzbif/0jf8q2aJJYq/RA0gpA8Fzwof9VVK7l7HCuX
z4bn+IJa8l4gC8XtOZwD/pwcyj9uMEdbhv0VxTKW+4jowLqfQfldTrCAh1OBpMe+
U/6FLklOO4AbCnLYc9FTBbUk5yfmu5NQurb5o/5j1MChafUQVATnBwDvbtTW/kqn
yr/NHVIM8W62oXtQERJcBpr0jBnxRPLdsWVoT6pZLoFtTgIhubuZXWGigxs4iQJ9
OZwC0ckxqtpn1JiVkcUHLfZqomF8NJo3CK5lOLXDYCCjFEe0vEOKIGJU7Q6LyUGJ
tW7Ch8kT1R56rWTdKWd2fhSMlurx2fRvP5h5jgY9h2E4PKetDbne8Jvt2wESqryO
RuwjiZXDqkO6WkyO8/eFtKONvcU+o5W6u9tEvOq1QLfqosTBELnOAzCR4Plk7Kxb
rO+9E/d+6EeTSIUs6JX3yx7rPKUNvqmKmchXfkf0BvfSFCOHTeuStr4T/8a9i4tg
9VUSj+hXwe/4zkvyDTUvyExd0D/CLxDAXt+/GVnKMABPB8IrM8VhQCM+8/pJ5fdn
wkQ2wl71ka3opNWnkEA4eST3SbZXVb810BVIpevwg+mIN2zmLU+hv8BYKIFZHfv/
nZHpebUv861Zhho1v9CferhFtB+OhKUZvjEzCMpBLXLsxQgSmbgjiPbRwQvxA+2S
MLDs+NydM3YlcNGSnwIBP/FMrJn7r6u5h1Tjg1FPYkYKZKy4j4xz29QBNlPnHwAa
1to85JSOnLXDJc0Q42qWZaLZqBK+0Rgegl9ssj4mpkAJ7bYdKG53Jbo4BLS8wH7P
ciinaCafMzYrnfYxtRPORxwGjIV/ajKGtVf1ptkUy8OAsANJ5a6FqvsCQ5cLp+/I
rtvlple1JrR4Iopc3iWchgO3uRupDnyLiIYDjcx+QzPgNrISnalxG+olD/nnfap+
l5MWsKYZ/nmNAI9EfEzS6Fq0SF76v8/WAg1Dqh8f1huvCYO5iXpnx/+6c54GSh6/
glO4+ENW45hs0NPp3QX02AshkCIrads33fpWYPpNUBwOZSrPlg0WvjDKjoxMFtFz
QUulmUbBMsJYqmimJbxkJYzMGwk3zjq9sUvjV0FrJctFtp7zWa85tg7Omdi0JX3F
B+WK0PA36dvJFz8K7+DNDE2JJlNsZtA5ZAEPPHWyJJhVtmpaA2XfafnxlH0Aj9Y0
JkW6MsX2qhoVyuk9O3Yk2+BWMHoL8VqfkmYi83zYa+Hl1s2AjQMQI0rsargY4rgF
RWQONqJcfAA+4NvrXDQ2oF2f8erybD5pvo10bjOdlhywooIfGjkoJcbbe4B7Mhqf
xXOqaRbma1miItR6BVy6lHNRqOrcrgnIRfD7gvymjYKUJc1LqM+KRyDACcJsgxZo
++CryfuyqqqwbldMPSS4IVxTOXkKocPgheuFBo50QoaK8jG62olJZxPsch3oGqrE
ujgW26CLRoL9+Eqx9Mq8791rRyZ8t3lSqktoZHzRYEpLQgGr1bGu+hQSpexww15j
7u+ie+Xfuhv/N/k8XnbCqZU9XgR5q1FN/4v7DPglU22jlS3RxHMhpmv1V3m7tlk1
6POQMohPpXRZfLU0DtP590SDVEnlAIIjlvMzu6x5/U58Xzf9h5/e6VndPBIBZlGZ
dLeSEHld9FQyf+07wJzL8Mc0HgtE9sUjv8D7U6SI7f6l5KfOGs8NNnLUZHgRaPfg
9UqBQHc0VvFN2aFIYQFl/o0RG6cBTUT5L5evaD8toSaq96ZdKzO2xHDvlG3vMBxr
WWj+j42C+y6MJ40i1v4a7SiumCtNOMGJeH9Gh0Y1X45U03Q10UL7iBrdIDz23Xq9
yUUZ0ZdlaQN9J81tPG/jqaMeoWuhwgnQHGxcEjj5oroUPSew+QUjhlwZvTK6CMAV
PAcPeBLvviiPrPwMehWfTBPPZVw6qRP4AGpyOXU+15X75VyHpQamrsSu3sAHpmop
ULNyprdUunkHfL07O/095L6eWKn13bobQpoycT3iSKke3ca25hx49OmXZUDk/V9u
TNl1wSVf8/BW1VeUgxQFHtoEhZG1e8U/Lj2ZxKZemw3j//zjmcDEnkF/ZGceqYfa
SDFGSOpc6xCf/HjVb493V0xQ5oFOLqQVfRvOLN/VxpOtRae9Y7LMhp6YE+RDZAL/
ojGY/fMqk3/+ypHlnuEHYtmTRH3s9JTbYN2Y0tgSE9IdEQX/8kIw4cQwVD5cJFO0
OHvXrvOpKSaYHfNJYGOArFGRbY5jcnoEjv+muE/ZVbfwuFL/nn5vhfaat8OBz+5a
pvPq2bKVgxJZezbTccGymOMHhG/fE+SAbyo7L6wIgEV+UmwlyEAO17TEsVzBYknD
k5R/JGnI1jT77O6KhJEwsolzVFRiSEebz4mWuYDxx77EkpBCG0vvHT6L1QyYCrDy
Eq3TRVsi8lAWhA+dqmn3TlTI+Q+bdsc8N6AHO7SGmI8aXqKQ1C7ynL+8EVxL26Ki
4omA3XCITu/el5PngR686ZfxxQYTCOi1YW2/InkmQgqCHSQEBLHHbyg1yalvgPun
8uUJ5NkrmXyWsr1hYDotW3dM4XdtFF7/p0yX5NwXl4r4vr71D42j69cvBV3pO3/5
6W90U90bKMTCBe6LIcPf4EttIdv5QYCkaFqmcOUFhL66ZZfkJaYlqPndBvSNlk6L
346atRE0FFjy8wAk6bqfc5lI5vuIhMSQL5N/iQGVu3tFYiCnvnD8NOtlyJH88ou3
3pmCQMxpFEq/l+Bo4N09Msmi2A+EUoPxt/vZ8eM2DuZI87pJqLC8FUWH1BiR45c8
NtOYZgNs8HJeFPoM6K42bKlSMo8euv4VsPLL0Vlrepq4yHfWBeQt7MSv1u9yCM6K
aD7JM33Pe4EdtsNppAlDWu5oPUNmEsMrxrZiPvjtGxQMN+stDU8fnCl75yXdxgYY
anjtIJXMIJt7YnyQ0MaSGieXK5aE75rhMqy16NSDFrdhLhvKMqhrATW07ObOo3SD
p2F1vdMTtM2gkKD1mRi4I1nDbQA2UgmiKsrfJDUpCSeGCXICbPZb5oa9Y0/w5P3P
TWyZZWR33qvpNA86hFU3/cnMXxMbbr6hwMRGnyxg1nud+JBzQ0ApOCAt9jf1Vuiv
w8cjyhWAF1xH2sipoHe2zD8U+B/FoKFYHKrjg4XZ2ueDofbF0sJgznLiCO8KdyVZ
Q8KUaxGCgJAOlbRRiHpvHytrY9uB8tYMEJ0Bb2WrrraSUOOEMqnxknCRWAcT0bxi
LOPTAIiGPsnau+hhij/7YQu3xt62Ckj7f56qCpGKzDSsoOaTePW3yyrLDWzQdaqC
OcZIWs8QIWFWRUJAwQPRobtbsX8oKcEpbdVFDjjcTNq3GqAf0dVa5a4c8ekLnMYg
vfvJ3RH8c6inDAcaYQt9+MY2fYQizsl9f/h9IH2kXm4Nc8TLwptRf8zePougEVLR
6EDY4DTxvC6gbeV1GQXxDVNGM/f2r5XChuVwq7VN2+nUTGt7ktHou3mGWuu1OD3R
malNi/oq5Fd1n5sbV7EwCOTdw5DNbbpUP8vlhTYtgK+O3PV08HIJL0SL5Oi2ahOo
O8dQkA2jjSlGdKt0Y7bmB95FdTiitkSkpcx65hw1JjKSUX79Oo+kAGGQcbO4q/JX
SJySR9r77qnaykTLNtwtL/lnN+MtUkIFnQdogFU1pfGbBMtk+zpirefcXtGVkt9y
NWF3pc5RsipeqndebQjQ2mujp+aU9B+C3NpYbc/QevUhr7DOQMhV+p2NzdUIUGpC
4Xg8cWgGZvTN9h6rnUggxalp6I+Zuqukns7tj+RGSjKzs8lwTvSMxXyyVcAzKsAf
ugKKsIv+MVbaSAJ/MTHEbVDMpGClZzz3blC8Rrg9slm7Kv7uOOZ9UFkaA0pwxEKo
gHHJtcAG9vd+3fJE00Fb5ZRxRGk+GfnwJFqabQmOkRJ3vDH4axIYI1gDCR7wGNZs
iCEF06IRVJpef2zQAFYw2DyWqiVTPSrfYdkKoEuSk5eRNtnl0SW0lc9aaVrxE2IU
ppqEqVOWbNOrDH5EeHQeAepVAP3kIl9GZWU2JcaitkhudB9niH/MSfQZmlOwpE51
VU9G2CSxq5KyzmJegJtsfzEYrSMOghUTPyFBPhKfe+DeTN2SBIU9GOBUS5TEq/sV
tlxl5bnbyqCFx+LvOKBehgk3GtC945hBSEcKDgSH4nz/gzPfdYgbnIs1MVdzm7J3
EH/R+e6BeUNi1CCGll3Rax8N+DCtt4kwfQezJmLX5eQHkYjcbN48cTxcS375sEHh
U5u+yzlPD2XfGNO/2Lgp8VjdEWFEpkytZ3ANvKAY6PWrmipZpiiR3J5jfx2pxdyW
N614xd22dY9R30Z5mi5rstDqw2BqkdggVChP0iHUV/cFRBQiv6mEYMCAYZXeh/st
RNPVP5tqOTzMK3bwMZJXwSTYXC9psPCW8z6jReL8+JCu6Y/etHTlsnTbGVl7T4kt
2oPltHpC6VhBDqE7XNJSZ6jCUc7bvs6bjdEOsZOt/F3/zPynf4c+ir+QamNj7ajI
5JNFMbjji7fFomhmmuf3HqzNSVl0A0TgfIXWeCmFnUAp0SadQGHcC+prgQfszdnp
9CB/2BlBebfnQzwjEZvp2AzTeCMwV27ZxRGm9wQGpfYHXigzS40Ej9jGMx+zaudH
Gu6mSdJJ0YiEnctgz5tIojwScu56EF6nKky5qVEqIVH/acxVFqh4WqecwSutF3G9
VSshx6STThFsUhY4EUYm7AYjyf7ucz5++5B9v0YhzhcdjEzH/1nwhs089LXNrwL0
zVnSv+hCOt76PNTs7GDczx8sTDVr2Gld9E16RgU/snKTfJGZp6pTvcIbl2M46p3O
2ir8JKmT0FlbUWcXbVT5sY9A26YII2iXiJ7Y3zlaGq28aVNRykbERnH+wfS8Dc3h
IVjQTUJDIvNxnVNJC9aYG5hVrGbxzMXLfDyp18dX9rYo+QSi0GufInQFGeL/HZwn
gAcAXZ/KZX/5/rFdIntDVEp31L+OJwhruZV+Ho+eTgTAVM1FnTWu5vkIypZgF5/O
KRi6svu6v7WjzOKjHwX/jjK+Lr4U1IaOhtumuYdygttLMu4Wv8j5y9WfclCNBGNR
zccIc8GyYgC6WUZYZVt8uJONYeFnXw5TwXS57y92NBTmn3ht2pebXn8evn9HWpnC
5PwM4xQGpCM49AKRuXeVh8hoEyZ3lukqpK/aKC6f+lz/IjIthykDLcqZyVnV4fqm
xhlAmVf9RiHjOYD3Ky8Kn6lee5OAWJ/iwpXc/llXCWEh01sQvivhTQi5n9Z12cA3
CYNqShUtLQc56T8+boSWhuRieDlXyf5j85aCn3aeVbvDH/GVOtjd2KyfP8TPKAZx
fVjntS9Fo6PGpbKSDJfM9pZXaFecaxtGJ9YhB35OROoYnHrC98rVGJ/anjUmy+EV
v9rchS4dHZiL93LzHhUGIS4cEIt/LdG6IEkBMdM3c9acOQV48bWV6UEIHQg5RE4C
QATnnulbGYAzNW7Hgj2P8DnuhaFiD4KDLEMMNIeGRXCh2gLFzSM3eD5/JCR8fLJV
+fA+dokYAdHVd3OoMdnbu1FwY5ZaJDYLJc88rK6HOprUp7ZKNk4V+Ql0mLYS2nbj
syPEkJjtc4zhf5nfeAr7ehvTc0XCPS6l8B662UmNs7V1ZyjqruPmlH4SNHJE2n3K
3QnwXscKbCSSDPBcGQJcQk+lavq81L9j0o0rfpO0llDkIXnKBIE/Khck7+1c6qRT
yNCjqB5hNxHS5uVV5NbK5DwhqdIxFWQ7fmxN2QlcHgg1hkapB0vN2dU9OnFvBLs/
Q+tTu7Jo4nIcxB8hA9tuZ0S4g8m/vN/yBrQoI+I4vfFMcOFFdbA32c9hf0dPQMHo
8GGgsh8j3+iIMeBmdAg9Pbac7f46hpqRUMA1vteIPVolRa+YiL5dLIz5gs4PbCQr
m4fCe8fpuZK4HNPB6xjG8I/uWAJct0hpBmLOzWjOilBYi39Sv1cKJ1VQxNuXMXF5
NfQZJRRi1psuP66tEioJIRbn8W8BnVProhWAoLutjYsEXOeASLnvxuwdZAgcFph/
VrH1KNTmZnmJ+jOMaRXIiU2+5Te0K9qtzs0IanG/ZhxcfJWQEmd3anU4fV/1Ynng
xzwQCO3x8mzI7GzwayIZM+jrGq/b3GJid810VLXkLkWjiXw9NsDutApFa60naSfz
g7VRmMM8jVX6rYlOkpBNvooyCmwhEOOOpKFlKjrZa7lG9nn/sRzznH8/cVeTPHY6
uQ3nvaCdAgdf6NDArH7bLMFlcMy2L3Vdm6S5v5+DLOKrkMhpNazVQNx9C7vXdkC3
LyFblYi97i5bwTV2CZVgct/nb0a1YxTT9VEYc6/gVBis5s0kJoqCeBQYO6ucU4l6
tGoE5T0FTILXbztnuWd8PEaWgyrfGVqqvAuLOcs6i1FILPdLQ9nGMC+rW2neQ/ml
a/vWZgIeyukJ89TakkWyrkb4e6e8EI6YmXi+pL7vyDEMZ5WWPT6ZbreV09EDG6Q6
hwzlz3nCMwE6zZLroBWweZirwKj0/RftoA6Ylbf5q6eNdZduQoLopsgeqoWj8xj8
j8ukGUXx216aJBuGKbbdJ2gM5/eKp0S+6Y7Do68mCIwe0q2bQJ9wdDgf1ckKPBr5
qRrYbHIUsgBTQKWLiuB7jMB//7ScreWlubZRtRZOnrIbwrAz45z2YGMyCMdJUHaB
PGG6/FgMnzvVAbRbxHUwQ56i2s6wQ2hC5/vCAb1O0xMufw/rS8bzlr9DFibp2Bi9
ZpmRbueQyC0OeiHos/ATqqQRN0qGEQE8OtYY3kqh6F27F8VSXfOUYjCSFbDxzx6m
s1uRqL5XO6z7XyZh2t5c4xdJWFayx2roqX5xp6+4lxvUuI4kTXFcVnEluJpb/Yxn
GyvwjtbGkefjFlKelz1O4ka8d3QR75+NgMO55BLHyAUOz3IDq4G3Lgdu9Ge4VRtf
wICkbvz9xNyqbuA4tnEyheg9JuX3+fbzNqqLozLZu+i+MuOxu7b/zZ6Ew+sMuK35
7Yo9gjO+QS6podCd5qg807rJJq59yYvBmMK7xvOVfyRsb7QYnp7SUCOpY/hvFI5+
ksD0wgAaLgMKKYqX5tZ4FyBoLiJswN4eNNKB5sI6VuF8L886sUJIlgu9sItw5I2z
zoVWUJuq6vja6Et3X+SeqQTFHwl3XmKxXA9ffeEW7yM9cZ9HvVvXUUcExtrNJuP+
jgY5PJRNepzsmHKrPwgbOIRxpuUlJGqKgKq77uTFSnjPLCyu0UOL/hZanp9n+jyP
BtXteN6ixggECGG7n9ZB/wFLRAqGQ8KfpsD4bAyUcuRODZi3eKNiC/fjqmfALHbH
zoZXrwqCmzqRtDzOj5PkIiSysH4PAYG+XGOtOYwYA/0v2yRCSXfL1p4JXgHQQjzR
xiOdy6HDdGXNPuV7UkxLit746akLdqD3tDwVa/PZlMNZ8SAm06H4PZbY97dZa3CU
HV+f+Ys0kuyfzbnvIBsk7czazme/FYHD+bxVsaxv+RkTd5QK7NGAQgUpZpWYeTN4
7hQjHZMzyDys5ANFvkWeAQw0oX0FrpvpQBKHKXZEa76qNHPsCgKwdZmiHgPKxh6D
dyLkBogdLwwKCK6zpyXRrjLCzzQTVVVrHS6aqx07aFw0GzmWfVoLlgaLAGkTFjV/
oqfyLE50Ozx2etuJ4RGjmsXZadAdXpuna7/s6kl2x7Y4o9/KyEEFUxYIkR8/UZ3X
QwYWtUCY5IdwwqZZp6Oua5jPdGgSYrmpACiIvGEuRU1D6IbjvZy9gHbzidTet4hP
FEU00x6jROP/YZkA7n9uWYh81XNxww3aWQ1mAtGcvAEHRJCyFAjf5/PGM64oi3qa
KKuXNPLjx+pFe2ik1oNpll8l9asUg1CUKHnir86l0P3rtNu3XBhOJOXkTGnT2UwO
J30XAUYEiENX4XwXYq5loRGBetV7cddwEXrqHP68+5BCxTsBTauhDFt+mJL3HSXW
lMuIu+ck72JB5aEn4BOQg/Uy+wAlTWEzCTLIM5jZNlJyibxbJ61Dv5d1z9UgRE0w
SLLWu+5QEB7GHbvKmZBZjDkA2UoM6okfCuRUCIrSMd5DNbAJMgQlTwZ6J/SKIXf1
4bsYV3n1pPPO87bohJ93AUUAT/6TOagJWNVeVjS4TlRU3LA6QMoDaJGmA32OeG8O
lkCxj7TRfuu0GtdQVVvS/zqU8sodetdfXp+Am3VJTNO6Zr68rJ8lPqHRiy4O75wR
oxw/ae5atKaG7Nex+X2+XraVX4Oi55AXSFqP8woOEOmqjx9GrUUYt4Ayc9UPfAOm
R+W7Lh8lA2lLY6GY+t1B3Rg9qjVlzO8+y6JJBYbaP5JakflOWv9z1G7mJn6I9QND
A18s6ikWIHKGEtZNfQZvqW5oF1hyiniHyk1XFIW9WW5z2mTzSYKanYj7eINZmfwl
jovJZVxTxaFZ5MZIDM38iuMVXRqDCQKt5WQA7xCWP5WVZ6OlS39lPzLNgkcdnu7v
MV/nSn2X7Z/DLTLwTpnJbV/II8PcuKfdpm9OGJtlSr2frMwg4cZvujAj44v+UhVT
OcAxeycEWRstRerrpGDws12tAwY7BQd0ahxt+Dm7f/STxBz/QxybG65i8xP0Cs4Z
CwBcmuDoOE/upTPkGpWifmd42mEShBMvOtRe3CBgJGDI1Ds0qu3XDpyK5ii7YAeb
ilq3To3Mg4lpS0VU86/ZU59iKehPRxVmY6mQsBtGBteNC1j5wmTyMgEm+cVsZY+r
cNkwg6VkKax6PPXD9/Vu6AT00Xb/2Ioa2gtsWXPREiCPC02CluXnYfH1vO3ZciA9
ca39WAeYuUlTuS8kUMVZfulyIaPzOoRpyBOMEFYAcOEAePFbAl7UFuLgAbesUIny
VTzQ/7mhytdVBVA2dk388/6ocLISA3ULUPHEmQzrZb5Qfji0WFfUb3vAQmSxH9B9
sH/wEUY/nQtJj6NBbiw7VgRPMtIF28gJ9Rq8si+Iry3f2HBhl3J3FlPhwvhaQcuj
8vH121isYIF2VnV99FlAtxN976q8S4y+GUyxDLB0+/t4DK0uctP0a1Vzzp6cFlVZ
vltqSQHvBMXuxU55DOKE6nUIPucwgCpbFF9cBhOOOt1incdHh5pwl+7VV36/QhER
ERo2w6S/knsA0+A0sMmAASx9EGsNaajx05xEXAu3NgdcUBcsQwXG92AcNj6yPHOc
P8G1lJYxNAHEwskk7NcG0RJoT3UvdCZzcxredmd5NDKhR1hfj5slATAyfX/qZXB1
NBFQB2T0M4rL0CqD1WeKh8Bsi8CZ2EdKrYWwY3Or4Pq7GqPKjQ/mASkv4k0FRnBS
PvZsVS/+dsanMKWonMAziZZSQayYZwgcGIW2FFG3dBZTQpfNCRx4B6+z66swgGSB
JuJRhb/1UkQfyUZateP+hPjLmDWNQcnfKZ8Hd5wCTNNHW1i+TddDBIJq7qHsWwQU
EGn+PdZxdhXkrHuj6ZApP9f2StA1JxEMoY+HonRqYp1Da/8FP6pteBMgh9DwwlA8
EsQYkElMhfjg+kBdd7sf5GUNtB54ceA2G/8BqrTQwGTnXZUL/Io7wNAIdbRqHmOq
j10ndQwzvyGwBxlqI8Z5mgJNcb2nutna9DdukfDmM+Om29UMKbE1VQrwqBfvBxVI
1fj7Hqbgk7FNSr8hcvq61xuhVYOO/vPF3H+aqnFmxDAqv647wO18uaD0YeSnqYre
AqMj8LTbitR+EVscGOQmVY+kv54QiLp6BnNeXl93zGmw2J9HbI0QyWeAymJws27T
LvZhEaX30/By7u6IKoTDjYOjCNM/r8WYqrjFMUVIbkzPFMI747pr7aOh7nAMt8Iw
CewGkdKYtQWp4Mws8IbpU6XIZqx2dDHkttgpP5JLDOcoWqK9c2Y8sJoLkpc8qFf2
PLnluvuNNuKnNfWYMR2asGapUO7+5eHa3yFJFBBCcmHlCzJo0CEzIfLwpgvw18nY
rLhhksxRCa18hY4/Xf+3D+tm067xfB898/MjQ37tYaPMlXga1W3g52mKtnDZQEaX
W/j8nxcgvZlAler5XdBQIiha5oPjpEuOZo2rSA9w8UlhNdWX9KaM9wZ/JfNFsNmR
xVdngO+jw+7Rv+HmLAtu1feuFOPBNi8lYz7lC/l7v97/r21o7rNVU3flsXlK2wwa
UZZ9bNTdRq+f9Ctt1Zmxit/VXQ5b9XgJMsEudRFcdL7/bCAE+haDpRPeNosAYAqe
UAAQjnVrGHebQxp0xOdOoPI9kgZas+dT/VUxj1KQ1SOcg5fkA3RDeN2T5b1ZMx1X
3iBSVDBu5xKu2e/1vgY9frVIe2ljQ5zf4fO6kTxEJSaMNZWO+nIfgIBPYVN0iIsX
g5u7T+h7vhFuYTscZin0UIwScVq8KgdEESLgE6WAAyg/MMjfrXv/MJUIxpbdWr5s
EMDCkamHCa+FRCZDKp5mmqr/WfnC8ZlBUOSD7C5YuBMZbpPSkV+11ivRXAChs4uP
Gkqv3vQqdECfn5lA5kNV7Xu2w40GOEt3JNkQQc/YAG2k9XIzNpGoikZIzdAhlwpL
/HhtnREnbJp6W7xY31JUI/pZiFdrTDzGymzqDUVwJSuriqfgYIZcuxEMX/+xwYHG
i0X60B9NtAADGONbBqhdzvE0HcnzZ3F97SW2NuHNSlQzB0XdP+mgupJhvK/Ajmli
kDUe0Hn1eVnJjTCd9/9GXYaHB4CQj/Rf4W55mTmgm05gXBTZadkWXE0RaOlRTjUt
+nGfj0A/n2via//TQ5lOGFvJV2s8veKHOULcAhB6aVs7ScK3lFSQoiAliwEGCOHX
at75EiLRDxgm3O+62UEJSBzUG4EwZCHFpubqec8SDIn0DHMHvevOuUSg0fdjQbqV
JDHmW/dHHOn0A6P4DU8r2xd2q6yPpZsv+YpEgp/WAmNXk3metLKVP7nbMNannJvV
8k1AoXdOGwY7eu4MvuYD4ou//dY6/H1pm0AYfP2Bv/SmcVA2bLlbJykEJC6xjbv+
4s7UzzzLLAzg/GQlJxKhH0G4b0EnKY861Fh4T9TWXPsQ0XRVRBSDB+7LnPTKGKxw
aXajIchTe4ZGkSh20rj7iklLkV/Mm9WspUlPGlIfICSh+XfRmcOGYFGCRm1IvXZf
vofj3zQKWRkJhmmc/yEuobyJFSVcEv12U4np6m9icrc7npcjrvnub4CS8qlrJdtK
Mi/LJYhEu9phBBOtpzAMg3eaT1cJBkgVK3daExYXLLF4MmA2DLTEClP3MJT1SVvB
yAAlsGAJ3jkH5pJ5Zg1Hs8nE2gRjTM/Nw+vHCok/21N1KWVkRPJ6timv/FudSys+
ChlCWVgghr93dwGMhbgiNDvbI6fVmmTaH4gBtPIqoq3uRenVJmx4B8LTvXHJ8XKx
VXNj1/30RSKYPMrwRk1ZF2FCRD7OQgQMpN3pELSV/kG4gSBNBPm6VmAvySzSjWtE
CqRt4Ijb9lQrcqtpG4VTchSyBx8XwupbNVQ2lg7dHUc8rjU9IqVQE0UHDuZhA/dk
hTgEujt2UAZ0LGPFblkZXj85BZGi4u9spfHYj46vIfsE2ZgGlAnhRjxHEAJPqqLQ
tdJCkjBNDVVuqhwgTpmn7nUNousICVU3segyED+uaQ4ioPpFB9miAZ5vq0BQ0AmI
ZMMk06M2FWRcZqKTy31mcEOslxN1Hru2nJ2NnUZSxDLJQ98G80ijJyoR+g1m1P7J
rscU3s4UIEmH9clABNzIRyMITkdhcPo9bUvLgVFNAH6DHrCBh0nwQuziBCd6CLCx
sWAxgBjs2T04vfiIBUkNptkwrQ6syyMCN6me1L5ll0lCJ6Tai75Piru5EgoMBOYi
2BGpwJ46T1+sjJrCSoztsEFNFydeanAUBEAkk22EoLtuA5DIRk3sAg4DpdEmYrav
SFR9W/Ybrw8P8ag4rKI6/+SmaYRKM9T1arkTzkUONWeDeY7jlsHGR7WGf/lN2S/A
8m0Dy/A4p17lAuzx5V3rAEp30NdX7yqmlTquc+NtzjgVrkaaXZgAcNH5yuP/EGMq
Vsl8X8K/ndwIIY3kjwlNvPI9Yy4x9QK69dkc2NpXf9lxOHvVNsLGM2iKWrsf1jSV
yaNqCI2vY0r67HSI1den2Sg0J8j+BW7ZD4JdhHI2Y9LtZXIYDHeEG8Zy1bHiCEht
xPMEq9IykYfCaFV1cbA6AdTfDt7l9UrfYck3A1q8H/OOGxzwa56MbK0w+8FHFuth
iXfxwscaqInRzt5ExLBTP5tmDH8cwMhKfePWkpW5tPDBASFOiW99qCPRg7bwez7f
ldwGzmnFpBAqXkNJjYXJ15fi1oo9G40wD9JhUA/C3sJbQPwNvMMuBTZyBNovs+SV
//qhim4IiYpZ6hi2ipDVJyiZmrevmAofIQ6msLuOqpmMMJCY3LS9nE95m7EG+0JB
qw+kIUDk+XUULOsdlQmnY4+cDWu2xR4rNZJgJ8/b0wOfLD66Db4i9fSTnPudX8sg
j9g0Zdj549/68BofmyFQnjWkkj8cRXetJtEzeTMZe0qX5RbUmKf0TMmd9SZmk/1W
1g0WxsIZ66qYz29uhmFBb+ZtYCY8nAf+XDltxqRAFnIpV2JEitgt7x9c6LIfGQ+K
2bK++p8maA1BhZnJbwGCDcdMEbXnr++k9KBL8oT/ilhDgp8Sm8ox9hvpYc7LK7JK
XiytCuUBZuY2F1VTvXumW2dpeybxm1nZasqbQo+ji+3Qn4YECQmB6ekqGJu57g3U
neKhSEvmueBupv9z3C3lxJh0AFSkX4JnaLCPHczNu4Pl+ELQ12QaFFz+5ujwx0nP
K45ILhx1tRRXyLAxPdv6mA7j2MwFI1e7ZplEhUinMxEWNl9I/BaYADrCIAjjhb4G
14wE4GxkoEEfTc+EJaqSYRcbc7pgxsJtvu+EurZrS7TNj46uvj3N78AW+gbLiS91
wp3ofvH7S5rLbLboxOA0k9O6GEAoRM6gmR/bOK5hK6582dRXwsSg/HJegecIZggr
9SA4eAqFmFJw5rETrGAAPapIZkk0AaHUq33NGZjha2utNy09x+TjaEQnX7jlYSd3
ah+ivqdWfHNrHeJ+Huwmvf7fEJ6nwv5nxXs79o4mKbvYxD93cyO3fapV28uhsp4P
55PaCIwPMxvWrpvM6GfxAbTnPIxTl97VXGdcDsDECyb5gt2r56oWVSX0twdJlEOd
+4nftq6UC224iQP9Zn66W90/mh/3upfiEVcOKtnJjZX5eRRj1/2ijKBaAWbFzu/p
m3P9c0VPpvzVvS29kAYoNBQQ2lQZ4qlanJg8cE+UXnQJrq7ZxzTfUxNBav20wOSS
CRCysV3rqVIF+uIpbxl3+aTQK0qgHGZUHOSAitbqSF49z7VtbpUDPG4koPSh/uFQ
4f+p4j1DNr8fy+99bkr9DtmAu225YD5vbXbawfFC1GCGMjdavZy0Qkp/vcCsxFnc
oceRjYdDubxwZ7P5RtTBPE55yFliN1N4F/0JCW8sfcJZEBEnanLpmXz9F97/IhXP
IDkx9C7yXT9GM6+SHr99Cd3lXqAtPO17NkQMYb6I/Sewon2XFTbJCxi/iscaFqVu
NYso1eB6NdnJp/JKsw0XUUL+SQwjD45iD6Im2HFAcPLvflZAIgstsUVGvkpym477
BXl46q6SbpJsMIoI4oK+29xhL3fQJlmwinvSeV9cQ7ztOSGonB+Z2GkfN1NLjxVR
f9VGTAQv5PMnfVEDTgsBLqWE1v3k8plgXDvfz+IhrC+wUNPprCZdiTpCHc60CEJf
j57u2zxLV+eWITWaJBlZzI0L5rSpFhYOUHgFpCVAcueGxh5jtMey4lH/qde7d+cp
i3yE+F3OtKPfjubNMnAO+dTbJQ/lAhMjgEDdMsgVCY/oYl5l2QYUxfaOGC4JFOIB
erhU3DTqh5xiTALSaY+UKsHK/Weqs/jasQv24e1GH6zaLqADuSFNq2s7wKw1DfoH
XtJL61lhZ+XFJ572HOQpfNe9fOsmOQeUnzQIujse/bLVgDJQ9VDM55wem5ke160F
5ZM6C4bg7+lV3ia8lUl6/3DNkn4fdEJmW20DKf1tbWyv2wnS9uDCzYIl9cLDcUmZ
/cgZ5nKeTorR3Wh8IqGybvSTGgCv652N6agoJzqg4+EqSdaQiUuv0ibCqZ5aY4tn
K1VWCH2BpZ+lxiS9Y6j2lMijVvoE8WymLXM6zCylmZtm1FWy/hEavKGEgDysPHT0
aOjtg7Kj1U0fdkUZqK9WwblmK0kP48HQlnxaqpPUjEQhiHYnTYW2RUDbcPNRLcYY
sApMraXiSiLahPE0i+LUkhNturchkJcsJuc5XGK3A4JE8fwbm14YAlnYZMjLtQfO
Htxu72Ny2KIXQzsvstVzd8PqHpkNVgQcRUDt8mU6F/PgU3tr4+2Uh5wr1KwyGWpf
lKK7q7aCSL+494ZcLDpTsBU7isXysooN2j1TwmI7W/RZ8ht9t0s5bYZ7g+IovLPO
cN9dWSbiWn9dpiQPXvox/P3kpf/fbYtUUlpH39yiLQPTZUfd5SCuFiEypuH6FyEn
sMNktOAiPEjRls2dhjNyoPQi4hHeqLbOtzC+55/vG83cAc4dytr8oExb7/SXa50p
QfsNBWAfyFqBPf307zZO3saistjIWz5SD4WUFmxEFmApAO16JZGmiem/Rhg4bZtp
/xweLhusboO5IueuS4tOD/LqApFvvNMt5OCcBQD/LccEd7F5OS8CzT9P3E9Z2f0N
Ns5bC8+bWRtFmRXeA4RLx72XQ/zlo0GKEjqzftqihx/xzoPuIbPn5SWCWiIAIf7Z
v+b0lTJMT2114EfXIThyTAh9H8J+G/Pj00uWcyJzSuBFRJxi3LnxX7gNkuOBEMjV
zVumy5vupch+1+6U2MDlghnsSHQ3W5qvIwQRgx+wNlaFezcljDJEIJXQRIjIyn3m
SBIFle6FUdZ250s/N0xydk6vITHFShChXt72aS1+0l2QWYCkrCcPgsWPMotqBoJZ
NC2iuyw1uPlugyB15FtyZHNiy2UkqFpIt5E8TI6Uax9Hb2Vyy7cHMQSGnjxtwy8N
oKoAjgVs/DVuQcz8RvnKOlC9PZWbWNbodPgH9qe9tI94NYdyLPkD5Kx34vX+IrcB
t+zv/8Y6P1cp1XaIIHh6aQ9kueGHVHpvyoy8kqoE1pzeVvWOwBq3t9/aupTRssn1
6VZRHrzQvxWJ3foXqFzrvLSA5yyOCRW2zLwUgQpPVW/7Ux3D2UlX5/zIDWW5xgm1
9LqvtHVMm20JCxqpHKkoBhVNirs57uE0wzWyv7FrNh4hgtRpXmQXpeEske48wruc
KjpeTQG8VWEdHzihkDGtzyR0rpw56KXUEnaC0r0X5PUpC5CrG5T5R/XTY8utlI87
uoXoVR8BwTbM82pQKolTpC1OdupqlgLfNVfV1MjJvE9vdH4cRau3Kdmvt5Y83XUC
nk0QRLgEdjcIPpgpXhEN5wbKFSfJ6pWJ9RHNMHuamGAFgtv/yGpT5YAA3/1QshbH
QB3KX0ybc3TUx32mHVHTFe/lvbx8nKFCShKvrP+L9pXQ3LKNi8C95PqECa/sNmrX
TXY337EIdpl+l6+ICJXC7Nj6hH5W4askTmSIXBgji0w3dmjfTGlW2Y1Ak7Gd0fYd
VS+yTK9/R54kAA5zLlU/HmrQ6/u/sMIoNjmnMWAucgB87Rvq9xvHD1jeb+pTwi99
qZ6bOFHkO8ho3amTpdgo04zzTB4qZU8UcCpfsKLyqhas7j/jZh0Dg8P4c8DDXAXD
mKVoA+921+Ph7xh5LrbQbhsY4+syVPjrTxtJM6m4P+XLlCTq+hpcUyzl5mGZJx7V
4+8W75QFcdy8TGGpxJM2CIwvVsjgd1BSWPxUjGEvAa8CzBk3EnzL0YOe4B/SRlWO
fnuN8Kwi74i12DelHUYH/U7K79PM2I39CvLKaSxKUq96MezyOkLSPn71lTXCZRIc
CoeABg41NNKSB5h+waRyjBrnTw1KCDUnuTnxXap4zDkY6i6nw2AIsHiM2zeTMo1u
cNAkeji3Ioyw5DP246kKPGE4p59BdV8jbBWgHC8rjjIslOr07yczxTMPmdvveGyJ
UHlof+dzg/gaz0RoUJzUEnKn+GzqaDniRAbjVHM95E8yazdUH1GIwQ5UZdNOyOFR
nNjzmuNbjvIPlYbmL6JAlZLY4VD1Ir8VsAkeINLxmIrb9D4//D2OHW5EW4Vykorg
ETDC7PHQ4TBTrbU71BaAsn7YuzRwvVqdg8jS11aZun2ETa/nEtU5NmUL4fvrKNpn
DpbZIZnirljaetInrK67EchhW9ux2XjIHBwJ7aXdxmeER361gtyOzwytY3gIMe4d
loVdPRkGEMrinT0ej7AtDcBLBV7QSjuo3yNcYi0BQHmHdxiEHxsAt98i77Bah/rD
kOd2CmjOwuRcPq1UZZ6PeOn55FJst7T93YpnxfglTlmZcgdTmElg8nS93VeO00SD
Qtymq5oPY5ffZMZ5DmR2iAAGr0JTLHNmHvldfpALyVdbjgl5IAPDrnUh8v5QKElS
KmtlzOjztE6kTp/TjHG5T/++XFmnYh9JWYy1Xw9hCHI/iANLRINuBjZZH0d4hYAe
iWd25FJgFF6m0auuDaSAVDJ/GsWZsOL5hn2ztt1IDBET9K5UkIzE2l69FyrPFrbW
hEVOiPi1xa7jCIwCbQyavGYlXSPjPtLXy5sxgqPx+Vs/PZVdI5n0FsBPN/edxX4c
T7pFWiqehTKBDbi9ZS0L9H/NTXEEeusf5j+T8FT0frx0Y6e6QO/NclcMqvSxSPZE
Eh3TAnIWldo36W9Tkxq65MQj3Ba4ndTAvXhOO4HQ1KlVbboiDX3j59umYUc89OTc
YzeXlkDWK7wDmX4m9+RJW0y90uV6e8mUrdSXH7ygM0fSRYF6GgouiVNhWCKnyNMw
ZUIP+HPpmDJvm1+v5scbYHfWDqUsNGQQPOuWkuBvlt1RAC689UhQP9XIUNVRs8Is
bR2+XlldBwNYtO5OR411yyfyfQGYS4vkOUC0Htk8ikhqAuVVCs6HCsSmiKexn/6s
Xs99d5cOYpDbFHzMGYGeA8GQIm10T+4jo6od37NVz1AkIFtLrSCP+kR8YVVHG8PM
DpNeaMDbRvQMyPM/Cv3ljCPkVxtDvFIGAHpHMcp9B3KkoJyyMTOocgzbNgJd792Z
ESjfio58d+SWFPdcQesTPZTMBQk2ncUGUHYTlrsUhKJNuolEgOwl/PdW6BK0DEvq
O3EBuuM89FGbeVijqLriGJVPFvEHC9Odtz94SLcfw4ThizCGVyuV/towq8RuxhoL
jFlTLsWf89VPOr1f45PINhcjUvq5I4RDp96UnHMmoyBhS9ksisR+qmppfUOBIeSE
sxQadOufig+WWRRTGOSl8oFx4xRq/3u/6aixyR2yS7Kk7dWwZgh7DDVSjAc89q8R
ouPFEFwj0jxQv2jPwxHum7sece13lddxUV91l5IJMkI0brf/e69O84B/RqUSKr+H
kZPOcfGOEUCp9U1taKDEr+3haHFKybSYUfN60h0S1l7hknbS5bU5IaliHn3cyyoS
gFzPEflQy7QLmRYZsLBQfM7e27pOCnnINx50c1PKl9IuJnAMpcNzNe2lf56d6NQR
BfYlL19RmeSSOrSt95xRyG233ZpoZHP6B5sn1iHjL/edBE2qzBtR2OGdM1YknTZZ
Wzi9K5sfWg6C2kyyosUVVKbS9aBzWvdh1E+sZSp2m4U2MmffMGc80yYGrPVaSuCv
diKcQ/cUZzMJMQ6I7rMd68Qh6cLW+COlD8Do3i57fKmeozUF2GwGg1HN9r2ARSFy
d3ve0RHHPvgYONk02Sg6hVap3n28HVTE4F+BTWZRvUrdFo5UXSMjKoY+mnYleg8o
wbzn2cx1FnLiMWdm7Df3PWo+0zA1i1IKjcEoMojBM6Y2BTtE1LjXKaoTxtp+8T2f
p2n8j3mgb/YG+URja/Lfi23sJMDBDBoP3tovGrfluMb5/GNqarSnLqom3bnaDwNp
auVVuoWpunBEBtLRyGlaTwZtUHtf1OSk0sPG8MOVqkGq1LPvTnDorLN4L33UXLV2
HgtavlfFrAuNRvmR6csYy79G0p6AXPdmtva8sAqS1ZhBPOfw2/2mVhchiPD/lTqS
xQjnj0gx4EH7wuoTQS4KO/6UKkranMOID1BEXVNyt47IpvEyzdL+zSD72VYL5lcL
NZyzaepUDqfazWy22a1ln5xG/BQGP3JvRtgMBWj5oY1AK88cGa0gl1XUbP/28Wdb
wE/US++wLRX7hYUqO82Nx95ueUEtdkWQKqvohIqmSi/6JjOAjaOKy3QZwOVOUuEn
7A1QsCktUvr9WWwKmKGQ9XKLBsGN9Af8azXD1dthEHgVkuBynIXFW9n1zXcqwIQb
xdwwlnbDbYqeOz5ozAoFCZSYOLGjPqm2GLCaUJTLHvtFwzq2zGVskl+sD2x/mBiL
VOI1CwuSAIYDtXttbRlh3teq3pnbESV9ysioWp78XK6F47gvkfrViQwJCIw0+3fE
kFYxC2cYhTjIZLHfhaLaDTIhSwYzGaS+T05DtpzFIdlB1yYXEKxV3HtpiqoquIAw
fYLCVTosmOu5oUD3BVyRWPYv96GhPzv45hvAtCT1Rzl5KrbgNgXSe8DBQM/gXEBN
Szc3vz/9cr87WjXb1boP+CJGpCIq7OxhDQFTVRYxw3TrANwMqadt48DMmMvWBq6j
R1wpu8Tcux93Y5Py1AlEF77mVzsNjIGRYSD30msd8QzS8oDrYNElhK7O8p3B5LZm
Xb1GQAep2DOKUfkCHxKuzco0WUBOfCsZYjUOZImhVBDAsCvgfBB6v/73/AfoWxDv
1Qsxx7IMFf0J0wviAdq0NNw+P7Dt25lxeZhEPpZht1wTFxYS50u4JxizTWlOt/Nm
zKalEXn0POC2wA4rhtWcBaX/0DPpvuPsYapZ3ktrmCjjSs++hdOP679QMWmrlWQg
eUTxqoV65aeCtLDPKqG4rnR6f+L1MCKsKURsvcexs0CjlxV2E9M4YwcUoOl+h+tz
jsZZkeV/Yy8jJr6pVz3OxlZs/vKaVqz1g2eglA+j7wIjY/tDYyV1HrvaEvuOQqEr
0cEnD2rzekzLQdgMQkIwXkYWAz2H9W8sWnomIf0jTHZZ/yQbNqIZe7BjzDEPlm7/
Tq8vzyAhMGHhzaadDZFRQDL9CEp6CmebA6OxrlhE1LvEz4YPIsWCCTP1v7S6T5gq
s4PDqiwE24j05i38EmYXmNgX3Zh02d0HA8apkStuzhrROgM0ylMhh6mBWDBbXYlc
9tJGhJRlGoy2/qZcz2FLWP5JRmNcale045649mQPFyBAR2uPLeehvWPmBlEFKs8z
ptorCJDWqp2ZBv8LLzncYfWX8OHtkdXNP3qcTGCsAztK+8akybbDgCacCVpLnu4n
R3zjt1R/gD7gOukzaDRI/D+po5mnOOtmSRGVsE1CsZdMo1jzDogbBtM9+dKQaTni
zwnJkkxoZuAg40O2dfQeiE4AB85C118/vWdkuq20U/dpeoNjF7VKhnrqGI2tM/5P
93scqHN8T97NvQ8wf61FOhxlXjMvZz/aIr9zwcZIWsUjufYmTy/855ilrYasC5l1
rq15Ke0lBDJ3re3klfDMscBn1t3IOwfE2GaTqR9MzRtWZU3Shw5c9FoKibS3eIO5
ELLSFlTV5s5PC9GYttbZ8bE7DARi595V572OlbwLnHrdTP21eoAJZLuPdq0omq2g
NiqCK7gnDxOQatSgj+9ykDXnETn1st8sCDLyibINWE3s5GVVlY0zKNDbK1c4+HVL
uLTIHUMapwFgusChbngsry8WFKw3q4MdIk2dpo7v1Md+g7UacIeIDOgvX5aMZUne
r/TkOQ9ZhuUcJbzV8RwgVY3VHmJgiPoX0ik/hKePoNct3F5CKR9oHJLFk6F/l4qT
704GTKUdXXdPHTa3xLIrLD5HS0LV+yWuqjS/WUBuPO2hjt1rx1iCpkClNKf1WDyE
JAc6n6kZQFxbaujp83IC3G/djWLMQNNKtOPa4BDpi6sAPdMTGmjZ2WbVR8RlbYVl
FjzPP1cqdiUuuyjYAcma8BYm6wVOjNK4sKvrAJDuLTubf+o2Vg+yUOV226NFKeG5
YoFv2oVHDu1ohUh2XPrPzwWoIkDcD7H/0mdWsgv2A6tlVvayWNemU4Pa776kogb2
C3pHJkOSfs7MtHXa+kHAowayWIVv96DbdUjyB+Vqu5d99xZHmEQolYuurGJ9V3C8
fFMlnUpIEXcMI0DmGHuU5PxQpDQo9nN70T13kTQetx0wB+wk/NPV4uzCFf5ueY/+
Xw8emxqUUiZLYaj01YQoNCMNu7yVdugrQrTbW06bf0j9yHqx+iAaaTmc2M3AbyE0
FvDI6tnrCoUOZr6WtEoXzOPH1V/iSgEuGu5Uc7/WMXSeduaDcO/RPvk9hS0UYKfk
zze3yZwFJbmjYMin6yFF9zoqXvJ2E3qPlZwwUin1grYIX/G5LXsyy4LagUI7VOxr
yGdnUIWSk583A/fonPoAHLuBdeDi5Ttd7i/bq12RxHdo1iLoMuAwEm7FhSKIlzos
Ir/iyF3cT/qDWnnL3J10UWznLlr3p4yUTQWKglLB8v0Ynf6CrGyCk2P8zmLSr7mo
yjg65fPXgYmIhwLhG2TfJX1mfHHygOjVNkUnUDYxvRh+X92gIwcVIk1TtFKJ9n0/
2AFdmj8BoT3+kVnnLBiqWqK/XGVqGDODghFVSqnP94/VGanPjcvCpBsotRUPsS/o
yR95kYtVYlRpsN0go1WCflpD7Bdgz5pz40il1yRr/WS+QSGkTtu6Yq8PpTb2PlDi
urD0NtbtMSCJfWFuRtj6TL9R1yGFliHeHQRhGCKhSFl7rjeX/ZCP3NQ0xFWukC0T
d9UGDblQo816vQYm+37olMD5c9yRfGjokV7xIWjBgO8OLg8y4cpS+ICOqyWpx5ja
Z7KKP9mTZP2KHJombWhnoAllvBgvanbWLPDKo5WCryo1e4S48XpZ7Qo9VH0DfESt
LCrSsBPYVhvN1Xg31zhArCGoGAbf3ww7/13oN9nnSYnSlcByX29JYrBfcPqOK0Nl
/ifaXTYgnJCl2QJYGZLLixY8+c/Yk31RfK1C4aWGotowPEiGFajO/2Ag/eEEqn/e
QGmt2H7PBiVkPdxfcoL5sbhYwMeG2lxQJGd9+wXQuBD+V40dgztUSeoyChBk/5tq
9JXLecJ03yPmCkljwAoBQ31AD2MvWfYI6xfG50Qjrwkup3KqEH/DIw7qwekZmGKB
ZYu+kIfQML8yxSl1l2yyLg9h/UuV5ULAGWGlC4h2uFBWZQtVW8lzFkzeWzbTzfse
9XEbf+WU8Mc/N/gC2f4T09TTv6Rk0SrDQlNab5YfdK0oQ+4VTZKWRjVXBK6SpUwj
tI9G2opFIlHq08M6JzPsXfYMcrKGUlgGE8GRghp9wdaN36dl7fPAD0rkuo+vp2el
VCPMwTjcmmJjfC5SsxF5FDXPLZFGVUlUifej8THRuxzly8wJBQjLkTFlCDPmXS1V
y07nDMGIlX/bdoMX5waMzkzvhRgTtP1cPSby3jquqIk+JmKjDy4MrsOr3IBqFCC8
WjRcOXBOaUubXxfeV0CS3kzjovyBga+znHwWVKUHghCZycFwuLfwFkoh06hKZSPw
aAV3b4orQUUhU2yZRsanmrBTnZXT09x/oq3asDTJZpl6BcgMB0ssOVtD6A5Pa4UQ
3KQSRPKpvYHBtYNJu0jGdNmUekoL6GZeyb4ffHbWkuTuFOXx/BgV6vevUng5qXfZ
MNOZ8f0JVy50OsIYsm1mEKLcY7X7duQoPXH3C/StsGQEtNHeu2rLyIYI6n0t8ush
bAwPvKt7JLW81Z5YigyMNfXQnlvd+WyV3EsxX20b66u3LbxGWqw0m6Ee3AEsnA5U
yUFDDGvRU5+x5Z8aPRTsDLLYUUUI2OLY06IpEFtVE/P9G9pcSvksVtIkpMhDO180
FSHLwIOwN5BqyQuYjQDmHMD4gOCe00HuyKBOZttYYwfw7ZwxDX0M9kOyX9XY3tkf
bubGV1xc2NIO8xV3VFFNSuAny0nz+4NENBtl3PcLO2IzLg1L7Su1dazcsAIzo8YJ
tF1yg0FKxhEH8JUwURqrAMiwaFjUL2I6RN1mx4fsuE9vxoh18XZk4Zjvn2e/yTcn
ebbVrCif+AXEUalAunfZtz5TssfWc88xXKtx2nLWWWsgEzLLcrYrlyC2E4FqtX/U
+dfhSZ3mv/NOdBL8fIBT/1JIcrRO3ejAnG/Nw8wTTUacGvHEqN0yYCG1a89s545g
p53z9x8j4NECFBMk2wrZEX6i4XyPjfv3eGH7jNskGSERIRcDTnH8RhziR1QNclu3
MpV7gASJDq7Hsh5smS6z9GrBUdB8u8QNcGl16+JNuOE/w7KloX7LBZJQ+NKBG71d
0CGk3gtEJ+0rBvVQakfZTNJ9+PP1vedBH7AkOIhDgaeaYLFck8ySgIcr6ckmvqfZ
xTmpW+LKXlMJGyrVB7smJt5ppgcf+tLraJEY7SZZ5TTpxmp9sqlTNazpnP+c/PZb
XHwWo1CUZnZa0P683S6oXxpBEYV/IA2AqvObHfbELbUneO7gtLO1nCeXPPI4hu5y
lpxVCa9qqr4myXZnqWRkGGAmALilzmNy0zkHbFw7LBMUfF7KFotZxSj/Z5pGvVmf
MutKTt3rLoHXcmwwlWweBaM5+awmoqEerLTnqVUQFcdiWM+wRlp7m1EG19aOxsVO
aGlC0+L7wyh5+VwTn3EscwBg6OYhYdVIGWOk2xcPuRWSKFekth3g2R6pLCL5UtIX
PQNjWOcRJKy/iX3kukadLPfEb/f/6Ieyc5fh0n1KYNVGbin3RaF5gJwxZqQPtqxw
ITh48yebccGnKDDMlUMuFBocbnMgJakl1oCuEiAIlEscXX1fX8aNBUomCB9xTDjj
Hm5oZOqCFV+aB+7azT0EydefrDqi8987wxJmk2XEejNq46vKDI1hW8KXhvcI6zzr
AbdfrfZFZ7L8HG4TXpdDhACsbOIB8Q43GRJ1/JZnNyGpK3Tkab7jBm9Ftx3eNCkP
OT5iOu2xR0grRNmDrNymScDrkHkmwVBRsyA/nQL+PFm6m/vq2C9foKVZiua0dgkq
VHTC9yoViEmTS4wstFH/JxqD5DDk4OvbGrzVH40neneVpfNytCIhj9TSX+PkhGpB
Vz1gXOP5CZmz+rOXWI+CSAERA6nrNgWEmWqaT3t3zKOJ4A6ktAeUXIzSXlu0tgqe
r/deEJNe5E9JEbr8Y3NtQrBXqZw31j1ALjyp4A414P3Cn2rVB43YYAbmhy7DAoZM
AXPnqTPKOXzLkSwinsoBGdJZniBMVelKv5307OtcbNNOqJbfi1ZiXkT/WTmWwL+g
P/zFU9NK1YxZdUAfURgDCxmgMubm2yXKCTBw2cqqsu9zYj8b7Paw224CWqybkL5V
OqfQ7hEZ1n2Ea1Evvusej7wH2R6epwQ0V+fopO6phBwuo99dc33SdvVl/kmGbBgJ
rgZefCjJ3f9t+cVNSb+Z3GuWgbc0BI7DVMzi1pA/Hwpz54Szwix3RUU64JALG3e/
jH1AZGYowaDD75q5zq0ALDT4EBbwKSYg1RmDhtfwqVjPMNeNwJxX3SLjlvOdZHSD
sQ1tYzJ+8ZG+LXsXQQTjD+E9agHa6bAva6CMGXCHEgFqEFele97wvZFFrk1gDTgd
f7SxYQF/2CFxpzMu9lsD3fG6+iL1TxB/3RMnZqLl2iQ2nKdEkaV5mOBc90XD7L0R
JVne2E/0WS2SqflPjXPk1EWn9QkCIoFM/ry7ptkMblbs1xZU41dXaRJUSHUpw2Ez
WqUvwjdDFzAs78zWWFot2jhQ19W6ZiPHIDKi92CfwpATtQoKuqFOHsokd64fAJc9
upB7UGlq8+MZOhJvT+53vKqcJ0QSoBsAUK+DrI2V5TT1xMb1RGGWlRa6TCd3H9jp
t339sTNcL4DncE25ruN47htAEfLWznY5V6C2+RgN7Tgqji/bT2SLmC9dmOaoGaIC
g1R5j6tNvGwnu0evbBPLWn9tddRJ//dxlhfxo9zMVKqVDNwx+a+hPfnj68Gnswex
vWSUYxBChRchjpdnhZ5fy09OBg2J3D6CtOLvKtkC/fsZ2Jxc0AwMBd2zClhr1NAc
lw1GgWr+8qlb09GLWWAjxVXcE30rFFXa3MwcbF41IbwYaV+rXQNxLCRI1g5Rr43A
be1Un3Za65t2m0HRgAJDMjVdgR4rt+6Od74lyc8lBLhqmGY673bcKsRaaSXI5eq3
wUoHowq8dvSLVThdesERf+vnkOFd31hMb9eTqCmcbysUGOHCKXLuQG43VS/2S6kB
tKUDaJFuyjCV8CWrCUr6a0TH58yan0lylflR/9o4m+OKyWbm2BVZZTn18rOG+bfO
0xK6Fe/td+0pFgLZFlCN1go7tC7zKhWhWRA1cFn5E83r1jVsExxE2zcBqXeGiZVz
aTCxyNqoTaOvRA3Lrx0KONqcxrL9r6TJTCMkm3Ov3YkOTfZvIu1ZkID9Izk7TGM9
/orFxogVsU28U9TiS5UqzBTHNN6hcrb2XCvWw9B9Seey4v69IrOmzqASu57xrTjh
FaflmF55H3St7n/dof9mnWWnbaSXh5ove/1LZzxT7L0JXjXAakP4vLniJdS+bmyQ
4l3ML6canoENj4UPwXoasbZ5AXB43FaiyCL/+rSwLyTH3VE23VPn0ZHCU6gtUxT4
mp9szKltqpmaKAP7SYappWkN0AWqahZMV4EUasqVbHSiKLxiSbJiMET5ld6292b9
i1o86HjdRKjZq+PFtsADTkA6p+kDXlMzTbVDfW7wubpGxwDHNZv8hAtb+2aT6IVZ
5Q0anakCH832j2/abrLIA68G6b8HtBmq/rRQ6C7CVqiHaAn/p8QxYcTA2Qgv6CK5
6PxjNDw++p3DKeB2ox8bfTGbcQzMbicM3Xzc7JRvHSG0TIi9JUBcxr1/66bhxiBs
oG3KFqzhrEwL9rt+7fRqjqc2z1FkV5pAacGJsHy/swIumdasQ3uHqdkqkatmGD+V
hQoIKbV73J3RV2vM5MN+ZueMvZOrHroYrxn8ekCcs8qBxogHjx5K2NqEEsFwebaQ
Z1wpSfXtm72bSONWddwcomVuiu8dyvvHNj/YSk85Gnwn86/TJTO2mtNVQ/sqYU0w
j0Cyw2R9vTOQ0mUOFFksT0mKFI5E5aMoflLgR2ge41tVNYdURgp2x0i0z0AnJsOp
bapv3Aa6L4A66C8j4LoRMaM6jZ4xQy14Bm0DxVSr/+dr/eaI1W7PZmVfZsQO+Kfx
P3t2COnS8DwD/+nfvfz67HGywEVezuV0cbo96CRsTnlCm0zq5vj2mJI/u+09TUEs
JLIdNs1WCdKfhgxfGeJaXgVbSP+Uy2+hMN7lClY/k1/aLqiQlX/rXEd7Ch7vePGf
cAbs6S52fiuaMaHYrzGAtd142mq9jYBr2XNA7eTm9LQKgA2db7HoHXK4FeO7lKdo
TYHvVK8cgrsYyIacoV+rLdorpqVqomOh9MBbKfXbB3ClB+4UTa+3bODfjyBdoBp7
ckeeimT4cwptelk2OLdY2Cfxfz5V6/RazpsvHPBFBfyTHI8x3zF7szcRwS+aR7WK
EBii9N3JJIPeNHESK2UpjHPjnASiI9E4DuLjSvuiWrYQ0Dr7cwssQocqe6caHPus
J1GCjzKqd/LVKyodZHJh6tuovmopTiqvXKNzspQInrOqYVDQumAFSdslzWI7jBzg
BXZzseE/6hExBGJ/yKL69pb/PKYjxpO6JzzMpZwZ6C3iWQx/YSFuPxai2SIgwS15
SKmYr/MLNlNODevibc28dnUYbVeSfjiAJj+oPQeBcnChcjXDU4Yd1vj+n6JwDWRV
gAKRfJM6lxHaVWIV60SCvhjZ+sAypPes+F2+vwTtXlFap1YlGspCB6G9oZCvG32J
wzHtYvkwQfyXKOJQXuBlQMyaIFp4ZuyrZ7UPRNne3g8a8x1DrAbA+eGNTpP6yAI+
NymBEfG6vwyWw/lpHuwvt+GRiwaBfdBKPPeFvKHoU9/WRk7Nq+fPIxUjXjpOYR4J
YBrzCM/en4fanyZ/FZxNNkq2topsy1pap47l+NfozyYQD4V+Mlh1jYUpPffDBfek
eO2L9zqjAWdCm3SEYe5TKIFydsebrty6+Au4mEa5dLByGDPyw0zGTbLfNYNyMaG4
ayKy34vAOK7uUaexOgv+3ufIA8WXT8laBTUgMe8XPzETvmrXu+Ue3j/+JZOxM/Dg
N6UlAEaOQ220oYwfvBMheNna5RstrkgPlekrbqUBUL4FXexM2F4m3kzQ3mFE7BCd
J/GYbhLdjrAa+a/35Xf2mR0UYTG3y5CqCWczm8z7oLkn4Je1Jq2VpLlvj7neFlVv
2UR1w+rcQUrgLJOow2AhPUcIiBy/3G5qHeQZ2Jhs76vV/GLP0s+tkl5y6HpjFJi4
IrdOzofqv2WhGKMJAedP1MtjN0kSywjtNP4qh29x6WF1DOEEjQsPYf/eFM70L7eR
w9+ozQueM8mh6YcRjLc44bs+t38LHFKc2FPJ3pIjWSnPbfrG6extEh+N4NIchrsf
eHVsKUvWjGuy0iZFvpR/tiBePVnuFvmu3Py/oc55K53jDezuYYeH635nYqGGBddo
otEWClPCSpS+dey4JxY7jDPTL2BaxuDgUhee9hgihgVVbOkH1vT6bEARwB1LNlRI
eDVE5ql++i/M8zZnyNxI7pBgC2bv6vFoChoJ2KoezmfrJ3DabjiL3KiWOZ/Dl+Aw
lWkoVkiQnh1Q8cUERuxvt0MUSELxUV/P3XE7ZBZRSjkQA8pZJ3O+SDwNG1/QR9bR
8kB7mT7zppcgVQsb/X5k1+uSyYKxxEloN2fZGtRMaYt9eV6JSBAQRnK93hMvlItN
4t8W4/N8+mu7hmDqXVxRk38VHZXACIeu7Kt4j6jD8ZEVgjNP4wMf74zs3f86+zXu
P7JapCuZFs6QZfLNok7OHBweuvMMPqjBQ+M7nMfRVtm5qP7hf6IC4Ope7PcntrMJ
SZWO85nKlvwcYhyjHTk7AZjXihEBfZK5kxjqj/Ewr/NvczTPIN6Vq0s1Z4xm+NQ1
4xqaocseOb80SMHgMQR1+YQ8M4isZHvhIjUs+PzvNLjoX9HE9T+t9/F1r9g9/pRf
hMHtILnryQf7xRpxiaZWqhiZ65i3lPhRnzTRWkTbycTnLX4d2mZpc5kTBHTqThI1
lNYJRfmIi771wj+hZWj/ldXxEQahkfJTTetLEd7uSeMwJyOzcKyz1pwMWpZdw/mn
BqFU4xYJxcGifsLH+TytpLnYf/8QrNNMP/q6mdqF5Q6F5UKo/SDmReZibd6qA+IF
E4hR3H5PX0EhF3EBD8NBc2EDa8Tj5usxlIgKZurb7AzyCmLDW5LLwfpSMqcWP+gZ
4X4MgTBoKLKsaFtOVHC2JbwfLXJNbOiosCpjwMNzZ+/MKpl6K4hpfxw32TRHCcxc
SdXy/CN+YTnhUwrEK4ZnFYYD6G3S+DDTdvG0BtW0jBdMPfRrXNkGTIE4xcmNbIx7
EOR7gl3XRPdkQPoeeiHV2Nptyi2gKy0a9faVZlBYG8BEdyLFt4AzCctTSilgUrk7
tLxh0+OFboiDHIycs6/L5FiYtuzKLfLX9tMfr03g8V+NIs7nSLL9LtVYSXc8vFzF
Gd3+Rxt6c0pZMiDJ55r3jGYVK9bDIKwTx36tZuEiKIihQbWAXqQX2wKgvLYbaFVL
ixBDn6w+MD2eDMVGiMYNG8bPSdFXpFtp7BUQAE6P/O3RClh7Z8U6IunFulyd52VS
Cvi9fRCI2pwcTi3Ci72D4qR4OnkNcglYdD+I91aPtHnxXQzFdORlqA060fD0x2/b
PJRyLDzio8JGe5dtw15VFHDc2Xb3fdiMUZjSqQ/UQnzIXXnPzdbwlIBvpDbzK9BH
FBEQXE+AGm+Kj99Uh3XIspBOHpROS/X5adO7Q0QdMuLM+LZw4KwDFbMH74YwgX96
PoCLaDUm0sck1I5sQzt0A15aziiOLhXtxpLmWOCgIJ5N1/lE5Tg8juhot0peeEiK
8lyR3urG5CTJw+Ad4l0PIn0HHsAuCTL79UIUweQ6rY/Pdin5dGKb7DM9kInAUpcS
idpu1rmDYeLkJLV2M56tJL2oAM0YNPj/qRyIZuaZ4LtzLAigLSo8SYbJKQNGXR7w
67+tWXiFooLW5Q7Z9saxzD6e8EGfdyO2sJREwyaC4PLA+TLoWMR1NardebxhoTve
Y4uUq0pmLOfLw8TzjT2/w05Hl8LR2VJnDGFchGWyQ3G46DiZGg8rKhnI1mvttEmD
+s+5l1hVFXkKf1oE7YHwvNwsXCE5zBB9J392oQW9TPl3UqbdqZcebarAq11BZhmW
WlXkDa2chZsBZJryj2uJXqOMUTX+Wb3HOP9cgErqx9oLYz2wDfB7LSfMzgg39Zq+
KgJtHi3RWZW4lmZ/B36zkq0Ybw3tZC7760w6UbYM5XKf5Rtr3VZIurQ00KZfzq6J
Jz9VnWutZDhG6qiDMHuNSimyDSAuJ05fKysAMiDxJb0V6xo9JPbx0UP/fU3u2M3C
+X7t0UO/ELYzjPmm74fHn538bixCWKW1vXvuhE4DZndJkLC3jbWRE+UtpDL7qQpM
4lq40uwLs1B9bH47bxdUfZYnG/c2Z/1lVbod/SlCxtu/Em+FQ2kraPjXsEVT2iJ7
LjugQWNa7riHtSBen45WzodckxjcfENpL5BgfXWxb96tBvYj/aoeLLpq0//J3L7g
Pna83GXX+hOcjqd/Tr2emD4G627Dj4qguGVEDf3NpqE7EgrOXdlEdEFERBj/ThA/
KFf8h73bBC6kyoTORWDu52wN1LcPjvacBfOa2JV7+C/kmqmuazoCaBZW0bWCUd7/
8mh90M/728l0LMafjfTR8WA2ggWPvjFP7HqiRgTSH9+UNSb05JWaOwn8pOfwYuAD
0lA66c0iDPHgNQggb1KkDmLdY9rT1oRMZz/BaVjflK66YOns/LRQ+Ic4fDLCl/3q
vKKKlRUEEH+pLHSyjcfey7GA2YKEDFlk6Xz/s1BpTxnYQbWZm8OMg+GI37pbxFsQ
JPPh/qLkjkrbAF4qz7Il5vm47MiJzjN+/Jt70mxEoaBOcy6jUNbSvD1gnv3J6c9a
PuuiTXT8JS7V81IlOOPjkcmP1KfIaEyGlmBNzlERRy0NDiJJ2tPQhLposmd06sUn
AREPjkyvc3NV9DW9uLLMsVmBKCR97zcAt5ZAYR5q0upy/Z3Li5SIh4On+jfwKS5Y
S4c0hdN8cbSmEzau6JEl7APbtZT7ihYI+1wf1eNbiqSdEYkj31xW7MHa9vyxlxBU
IfNNLOWjnA0zqUU8wXrJcuDTtIXi/u2i25ibljUMlMBo/MZZwJX3ukAsSqKktLxY
/8iY9r82dns3z8aOu4XsC4BlV+zFTfCuL42aloLvY6USX9Ur/5ulCrdkHyQGsWHx
EODJacgJRcu80WlwadHquKkOQf7f2w7rtDP2DRFKk6xIRhDygUmiJDiIYxk8h6io
bjbunK5UbtdiReLGC1U04nCD6Q84cVnEGl6go17AoV4MvqLs47GnNSV++D8JiEVl
4wUOw4njLyAGK1mPgGUlq3y0qXMxAbH4N7pXNgAOcoZm9CeFcFHuVQD78jmY3WWK
uwnUk/X0oHvhjWGZ23JiHwxcjF2/QWTm7bfZLNFe/gO2JTpSV0fUCtssxM6gglnR
9PlAcraoV1tgkVh6bxLO+fqjVKaiQYm+r0pdF1d5wH/7zrAqzwu4nou+MQz+F9nu
REVxuBky02z81b9PmrGH5caQk0UBCoLo1ho6D9cGE37WXKVfSm9zEIQJqraXdK3V
gQGC6cSDc9s88OMC81K+lMZFYwvcWB8SQQqY7WAQyVC/LshqWxUpDhr0ONUdlm4f
fYmuxqt8iG2/+4iRP4Aw1ggZ4PG7Mrw1Q64yqpINEktUqgKiUPvL6kvxgxfth7U0
mAgylIFHbacE/CZd9WoVc7nco1DyNSCrI07QZFMoGBh3bKYYI8q6O5YPNncNanPF
J08/gIt32kWmssbXqdlR8dHzGriOz3tS9ebZkkmHrLiMCS6AR7sKuYgF3ji1wFtm
tdQS/69IESD+Jv1t0fPOs/aOwDRlmRZWzd0BEtloUx2OrE981C/01busCGO+eQ//
4n1nD/Avh6jLS+Oj6pdePSI3Bbh7ShikFEA9EBgQ48YTMkghT3ZPmOIahUaqG2jy
Lnqj6iaD8QgqzgvdbbQOr9eMCipY5ti5a7om5XiJI+hm0Gp5Kov88dpemfWfqylg
c/PtqbdK6tufAnWT5p2bytYWuS4i4koTJHrMVZ7kVDeKjRejzp5kfkYZeHAdsA4z
HwHrp0d/nXgeoKc4gTh4sE/aC16KH+1MILrE8ONXUo47gxNFWXt2d0N/LNIycBco
XMkuqyDE+5DApYVEtNretTY4iKITAEBeO+MleqhuNL+gUKE9ZHvS9AVw6drooZn6
6vVYlH7Y7busA92wVmGopLnALewsLZKAyvj3/jPqrL4YUdzdaeilE1PFFAHgbIzh
afm0B/a5qC/og3uhxmi5zWFty/6zIQSORs97uS4Wq7sSrsTCdxAYLebUd3bq5C07
Q+kMyW6JCWU2vy3ThfdhLZy0bdeboM2w4diFwSO94UY5lPps7h+fKDrFEhyI7fXo
DNzTqyLPe5d06FSocmY/yqsh8ZGlUc3QtXIgc2juxFZXio9vcavmksN4bmn86We5
qhGvUHRQkMc/ilJvsrOP+3JhIefpc7r+JcJLURoud/7ZHvc0tvrCUYCZZFxvTOpM
/azQZY0286n5W4/U1MbaqRwubtVEp6Pt/ezfX+Rl4ukic2+p/adLKreHpGTxWauo
Azlt7YtMHduT60G9iorzhxWlZB9XpNBRaKMjYizlu53cvcOZTuPkvHiOJzZ8+dC+
YuAezLBDjEbNs0w0eB13M1luJDrb4HyuoCaBEzPpFX9Ss03r3dY55qRAyP3f5Flc
hwwqFy4gtkxE/KM42NHOzA9QsaLVyUT2rwzt5Zrd/YGLFXKnHeLDwtboSJkXYjZD
ZRbBpXoALAc21ce3iOfgCK13O3/eHnk2s6IO4GIOmrFgbycuuJmYCUk0WnB5KLGS
0AcGQu82txgzapgRiDm2WJ+XSC/dsNv5q9yojQUIxlENJjPSTS1eqEP3lsNL0WpR
6V1NGNmFjy0uRZ9sT9fVKhkIXrw1BG3BIqdABx6eIKCo95hUZIuClmtnwj+14I1n
mnGZdweV5H+xj8HaWWaYd7N165F53CDfRQG2aiVECNHuo5wGlnOLNM4fKdsWrCLK
Yw6z+5tvyVInkRMHk090OJRxetK/GrDJiMOB5Df3tpWlFjWVv2BPKLH2s4O8WKMA
DKsPn2hZ08SZyFMqDW8a6nQ3qgYFkwMNbbUSSs6KzgHCyKWxcJVuv4LwDdoDAbSy
DURXZYf+n2y2vXEcMDuahTYSybFudbcfsoIxGoeLXRy5MY9RMF7kEDRN3GcLBkgJ
f6k8xLFLpcZNwbOaN2hoLxyrCFwzsf10cZLcTW/uGOOMvmSYA+a5YS1S4vS6N2U8
oZPSrKWxO6+wCuC6r8qVqsHuiR6buQFMJNWUoLgtwwLukyyOMT2i0N894PKKxJ61
F+e+ID8qsn58Y7jcjD7cSZGWv2Z7wpzB+yOx0XnixCJ2F7AP/JjStvhhmfbZCe2Z
qlYH1nMxGWNZRCVmloKuWGYmmo9JudPk5N6QYXZiaQoYZvuKPYEs1ScXLrVDKhbk
KQfWc/KLer/Bm0A1OmLQn1PJFT8d8pDR45JXxEvoI2ni7Uvh37ayqrdnWHMh/HIR
Wmzpl63QoVrCOlf80gA7JwxdUwJ2Na+v94qzT4DAIausMYOk/iRhItgrhhHsGK17
0t2EZGHCFmvaI/hLcxpvo6drwpYjL5dZk6c7N7SPXtN4IoaYIi9nuRO7hhVpzNgd
/3/PTAkjE0FXYyjrem6ikWHFx8/K+3hQIIHZNQydnK1Bn58f6mcbjfuyFB6h+WvP
wfUGnszBwDN56kR0JAkZu7+rhT+4svIskJ9Q64ElboprdU4gUrHe3tuhxig9cGBR
qEleic6OwkVS3qnahQ05F+LFdjAQvOzBW2Das1joOAs5Cv/Ev6Rc5oWA9S9rrUmM
tpSKxXOf0bmF5SO2zneGQ5+qKuoenElSNGTlBEuSzszJMnpJaY40+kbr8mzeAzAW
SKeOmXSdUNdLF2ELksdUdAglm6wzOwx/madD4yCgBF2bs0MZvg0Ovk1By6kTVLBq
ZQphCgTynXGB5EiZlja1pkUzUE3SaP9y6XB1Dvr6nkfXOO22KQn7YJJAsaAA47Sv
RosPBq9OAZeviV7DVWKfkf0gwesardIgPy7IwokP/zba8xxdkYGwWDJ4hOzOIOmn
k7boTcBLHjwPsBK2ow6ePhYGIm/kedSTKxmtUB7+CWarMd4G+Gd8W1lQ3e3rZnvt
9NQn66yO/Fss/aleF6tpQqM/tFf45Yg7Q0n3r2+oogGd/DRj5fpPIJwbV2OBYt0s
1WIi02pxcKMaTSGcjkST2DdYzgkgf0Lv5/SZgwlwq1clEf95MRcRyz/U6QZ2hSQv
dtnnBNgE/2Qkl4JLj1dsqx+IM93Cx79aVdnF/gws1ehsu61UspbYVnEGhtKQrSxb
5DNu3bBt+I/pg4ZvcHvSYbqpdzg9dMP94HJ2Zt1dVYFCJ/qMen8c5Lhig8WvWhhL
A/2PTWWm9sDcEyoevxIfT8qjG0nCYf7HvXKgGq9LqI967XiumJVktAlvI3ymiFrS
GwcAAHJGnzywXg4Cl1lp+76mWLmVLCRxFlC/H6lgqTHcjh77cl1whaV/s7FXZ4+1
/yzdf3TdZY5aI4/NltUxu1o2on1GSPjahL8OGwd36FOg9Z4VAjwEoB65Pz2bSz7T
ZTk6Wj6LyNQ+0YwiSbgznakbC9sBRRzOnlpQ1ge6w1O4mB2zS64DlZDNsBs7IExo
zVfsNMMxHiSBZ9Z83Z7z1HhNEuqrTBFaO4ErpGIG61+JDOFqFE3ZE8pAtNqsXIDh
phHzujYGxpMzMstQwoBb9KqUA2xxu+WL9uu2hDDPo74+o77QzCUl6aobdKw9ltgR
vdAwwuZ29y16MZfSKgckEu5gsqj7mprpKEnGKHKFhvTMsHjfd855R1kPi91Bz+Sw
MxJLJM8FqKrdcIS02DQGDUzU7RCrdtq6+V0Z/+DlgL2OpyXtw9lOVHrW8i+m/Fih
y1XO84zmLY5rVSiShA/4ArrvQSM0GypEPyDG+/Gijy7sb6Qd+13YjM91EbCP+Hy1
fDYN0K7fRG/8oNfZKUP3g1qWzjJecwL5Z00RLOXM1kAmgaBGhtNsbyHBHtbljZo4
IcuOEAJ3TN4JD7R6vF0CHZzDc/10pjO9mJvShZj4KK2tCgSu4ChOlBHDzirHQnES
QHVvnTw2Fn4ex+IPbo3zis+wuXOmpHDzPII1LZUkaHughIm90OWHRxH9ZP5DKhhr
JBIa9p1ExtxTQEHt/BoVsCSIaz/ivTAGPREctQiH2FHZLx7uxFv3AO1x0aILObQ7
0bg9uYAcTuKjUl9xxYLhwB19UstblJUMO15XEnVHujat1xz2zFNY67zav/7958Jq
IfoXEnWelS2xKkMibQMggtvZO7/FbZA9Cxcb9MbF2/xN2OIVeqlaKsNDvyWSuocE
SdOZ8SOFBR217D0nSfDLKuR8/8CL8e8Ppie61TfToAusFBxxsMz+e8E8jyocuhLz
J/PsYmxQ6CCYHM8Qmqe7mtuvKM5LzdgMBERV7rZGSHrivnD95qlCRp5ThNknDIiB
/woSzd3upQR1BPlxGtnSvH4Wyr81Q0fh0Fl7yb90KejnBwz8xVtwA8PSHAun/I0a
8IqUWQumuGetMK5ci3ClG6TyjM5+gWw0o9nuf0tRpqydODnshM+MM0AhG1o85Et7
oqJV/CL3gFSRQuzHNeTL52HNNKBeDcwWZaoSIHPantzKnozDP2UwIClc6PABQbj/
4wLRP4sCpTFp3rpzJ111LeclH+b+tWJXtIRhZn3gm/BM0k0jXf1pApDBKX1V732A
m3hX3ngaqS9OFlakcvyor06n/MFKCST5W35QerCkYd/qxXSTvMC0cYtidDgxHkth
N38LMTrbfPUrTzpLm7sWvUV3PIJg2seYKqQoQa08WfuvA7MShAHyjMCRcC+Ill+6
fL3D/Dw/LEG2YD282mkW2pxsPFVRvQepVjWwhkn9EPC1vudZx4qOO17f4BF+bp/2
/c2N6U5kJ5lVMWkOvmqCU4zPg44LJg/GgYv4z/EZ/I4bhx5LH2zl4io0hkRxHo7z
zErvBQg6Xf8WXfLFNvbGi4s0oKOp9nCH2U7+sMmzvCAKXSeP9k4Z1Y2CdBqDpYC9
bVpL8+TLbqXCiUUd4GT9B8x5UWtZV6jKAnvTBmyRw11x5iqdCg68g9H8n296tFGv
z+446jdrJmeQy6igpSVphjHb5HGO9UqxbPteI6XTclHhZcKk/xB1hvUHkdpCBdys
hJj9OhCvNMedwN/gKXLeoo5G78iBLT1qXvGnooHNol0u/wFyETk2g6bVrBTYQfC2
i/Fx8foZeqcVHF1S6gV9lcSoC9TR5f5ccVmzLbI7+0NIAJCbBG0DGLe/nDSV56qp
r+uUiwe2cVn/yh4F74eq+AA4ioKY6P/j9BEOb543EJCa5Cf7DuRfkmKyDqoBV4rt
f5xElrjfXwATk3IOhCsiDzYlkjccuuYbAvmy4tDkhMoKkQRzVFOxtlm67KesPTgn
wj5D8Ra3HvfU6u2mcbPLwhx8V4Jp/Gtfa8TyocEk3kLVKNuk6C+Mp4eYKtUjAZ8/
xRM1t8f/Ub16TtTu9qHA6yA77mxREHcoENgWYqIWhKUoZZyM1iu4XaO+zTn5u7ru
xFnrzwCwRT87D1DH4erfLxkxGGo8t3PKC5tQRg6zr5v/YTHeVktod0kmsVPt00xG
y7v/D8mVS8Cbdqmi8pIn4fNU9eax5eeAbsyS057u08zyk1LjgV8VjZ9NDhLf7dRg
1kgZx5A/g4g0/wIeLa5uQFQw+o9/M+YSRyybwRyMnByt3lQy8Wm8PROIFY8Evo5n
GmykddQV1I2wyeDsA8bf9pPckpN1hKafHm2mtC9nT5Cjr5JdgWC5cXhyvQm3xC/H
aQlCfkNVK6PLGhAHvHTIY8ejQOBYbyT5AYcN01IHOHzKDkpAkRLY6tsdxL9Bl5Pf
vHa8ny1boijlJ5zpexhQuDfXXMOcHcHB9zgcLfZUW7AU/ykePP6mbVtVZYyP0iBY
CASPQAOR91vG2Odc/K4kc8dgb0BKrktcsCA6u1JoE6L6P5stWiJqgjufz4fCM+6v
BwDYT/38M4hAGIJQoMe8CNSBXMK5iUKPwVYY8d0j4ARGiNYj8HdIwg4W34k9Zc5Z
mJf/SU0eJEVUaKncedYOuDiJJKoZvGzsaI1I/mDK7BY9FfRJ/RGBiPrIweBpVizq
mtjxGoT1XsJEGHN2WfkAuo7ywfo05AEJafmDK2wgXJZK2aB/NdRPXdixBlzs/st9
kd+nDHrIoLm7CZU+AZVHlRLEpnoNFn+rQGUYIHIDhksl5zBGnzfD/lMr7iBtF7yd
AP9XKaQLiMpj1RFx7YMRYB3SldjGkf2nzpoSs1Wn4H6WgwQ4TVCiVTqGk19cX2Oi
c7xbluy/OoK5GQUJoCEPAx3TkpSx94UeFXBIYFfklUr6ACCe3ptUmrVTw1AoaeCw
7qktX/cz12gdQ+CG2QUTj7pTv6VngADIyQLZXfa0p2Hh/FI/UnrPKfybxSCGe9iE
szZNLclYfZ9JgPaL64kA5MSCoeNHcgjpM5EttzXlBzOmIZhf58uU1AoAarpUE2Te
wW5bsmFYySS7Jb3Yx6erbAGNTOvkPlAUFjIi8Oo5/Z2pJidGnUK+np7c3GT3bTGf
Avv08d+h0d1ahpXr/K+XRuiV6r2adl0dLL14qWWrcx9YOkWQNcIHhm6aPG+lALSF
dKqo7qW0GITrLa4HkKPfLwXwjE+8P8Gmnvv3EdjhJAfvEInsIqLoVD0eweH3nMwb
RPn8emDDVW0nysWNg8LbgVpyurFnZH7qC2zzxsa56DjJX+7qDcn1g3x5wawkJ5sl
8jvJ7kSDYg205m4oQC6E1p0bQG1Cc3zkqPefNp7+TALXLA3i40R+oQNVLuNvsbnx
Y3ckBjocxHNRRIC5nVY6IoS2fwJ/63PfV0m/LAzTMjBrytBQ5gu1WUOoGr917oed
KB+D4/QA1H7kNEu3JzzyGMUfVRaTHlnutLTqVSbIvzIjK0JClOgisQujQH/4Y5jt
YYKZKhAmEP5z+vrYvris11ka5+JAryLZ5Bk2CpDXFkRKMSpCLHWgBV4+uFyovYqk
+guBqy3l8fQ6dNhEaNa6EFia5JgcViacBN8J1Z1Tgt8aFUb05L3QSR0kilhQ7zdH
ORuQ4YwXpmHr48fc9WPOGATt49eKI/DyNBwk7Gc/RLfMi6OZwgqgij2TIjDK4vD2
BV697fMYCEHWJ/HuUqO843LGdiKrhSvtZyeUISm1PjueBHkoTokSjoQTQJYEM/y0
UVlVQ7GLsJ+8cStd68TpjZyLU9dclsuQ76sFDq+ER+GqxGGVH3iXnOxqXFiW7sNw
zf/G9pCwFUex8Z/U8NZBaQUtIpmFX81PAgumG+ujxRVIgyF7rL+Y3ENrBmEW1ii4
7H0YEcrlHwfDAJStduXXKym7jnaUm1CSO2c4NDxNH0V2YW+rb1/PScdm958gTg8b
pCnpH77iodHvEBmqaKQfSE9/VZCLdG+Zxb9BaDV7B6oIB1VK3IsP1mkSx2tV9hWk
t59zlwzJmqZWdst3BJiRfWX0g0Mh3+W7BomabHAD35vST4ZvQ8Q/kA4hCOCG4DfG
0Bx33AM4KcEZmXxQljmCAc7UExXk3lePXbbnfK7EFeOkVhYqm0pQSyU1MOBYTZVf
rZvQs/Fj5RWJDT6Z5c/hGyftZ0haDIZasCtqAagRndqpPswE6GwxJg43dLXmIUU9
xVkGtp5QmsUiUEbYG1nnn/f8EC/79ChH2TMjN0+jwJk3Pj+TrYaRxo8BdUzyVhIG
YH8Lw1H2erklQ0Ok/6UZgbmFQfzKRclZ9cle/HBoK1YNf2j8bLJoZ495NDrbA5MV
D4ghIkb1OrV86qc4lxi7H0WfwcE/Euxv2wrrRuv7gPaxtOVsE0tlVUOSRLxjk6+g
P6pJb+i4EFGcXwVu4tPSNDxpHlVLJaVtyk0pJZRI1s4pJSOvzV9BmvYcRvwpaA93
fYWYeYlcKmtZOI1cFnhibUwN2FNWrYpHZoH0lpBv7MOc0Okj2/6aHJ0qR4rvO44t
HeqEqEl8L0PyC9o80OO0cDz0eggH1YejE6GdU81ByDmL7P8SYqJZHqaaEvYRI61R
8ezyk5MDpR2LU1I9Tp0O0Nxb560kgl71xgLevG+yOu3ipyPEyZVlXWOCQo+n7Vp0
Vi576XDQQVu4IYl9SQRbCvvOzDvxBjOCP0jSoRHmHvDOXAF9rF0L0Dmyf6L8IJHk
915D50XNojNmJCJsZeKvXWLSnVCWcIKkyAVyYUzMVSXkdjvTJkNVU2hUe2VjHG/F
CVZMyleXqqPc0D0ajvrNLN0zt/C47y68xze1DMdhelU8B/V9070FuQfUResOmuDA
la6XCOUcAWqEukn477fgP4wmlSQl0Fd6/UK80HMwLtWqyIj6LPf9z1al9IsnlD5f
HNwSR3QXfz4nhzZUTk3kYvF5ryvgEHMrDGKoFCoDMPFRpqpxpqZq+VRU7WfjPrcJ
lnk4SYYH50G2/AALNpYETAT3/18Yz8yEzj/TGRY4dnQL45GyiB/xKgYAap28ocdD
MiLX2qLLaClPKOZtWu56q9XSayYIvZ/vBrGKxtBdKVljQNrSiEuUAQkOIg0r+WpK
2zHy603+EjFA4qAguo6bSuz1IUJQsE7iUJuagilnAsILF/QGkR8of9RZJjhZvNnI
gaPdj+nVqMs6q4Ov72jA0DW9sgAbCDiDkmvUG1/cPIeaqi2VqExcAqCrtK6ONO1x
JXnZGUsCaLT79y0EriXo44oFqL0vutyYEbb++ONqdMBYHzIN+VFDgqNT+kXyvBcX
UFKN1wexpV7X+jJdVVSbDod7THS5wisvXSvGyKNa5MSmkIBE7fErs8ufKnycKi5p
lyqSgEw8H8cWxD511umuqeoMq47070q/1YQq7zM0ptoSgVU8mVUC/9ZkP+sJUvpY
3XhSNdvI7F1BLvDnFY7pPWfA8rr7b3oituTvvN7ueM//k6qfqV3xO3MIe5LducpP
sCfLPkXpK+bqcMSnDdnlTujhzkNzIMn2OMX4CS0AAlyoPM7tFY7k0aRazE7g3FuH
d+qJW9RSxPdQjJjeix4aiO7Q0RSb9OOTS48FUHTcKb8OmtGUVo1TFaylCs7wwteY
WzV2BKwKsFHA9ddQFUdyF6veLQkvHivIpSFteS+YACCTuTuTUT+dL4Lv9uTUfTGn
uIj7zeypuArQQOIPb4piztSFJq7t/DKNtNSqTWrvmoeJAT+lcsMrWWMfHwQpqLk2
zGQB/boxPdFQbIpdjS1sW2QCq+X0CVdMBTvhkuXteTjsqgZtBste86VHFEWuwIOB
JlK3YAeEebWDAqk8gLaYuGCEGEEvY5BUbzmX6rI1QCAyEujY+xgDxyk72j6TCg72
mqhV6T5IegujmYIEgBrGi9QoJMfSbT6MKhQlzlovhOBSph8k3u2hc+yPPiG6OFa3
5r65c9e5s01WYYofiygdSeWuoEknnuqW+IyGzsmWmeqzpC+0KWAoWRpKXorAI4Wd
7MDq2WRS6RYntY13J2W4EWn637DPe04bAX7CTMtDfkkKrcYIQanolhtppKvEkpBH
HpzJXUHO8PfzzWBMaWGISaSUyo1uCTQmgB9oF4m1dXemNLvb5+iMd9jxZOnjjV8C
BpCoiD7yhc/R5O8OFIZ8HVTwI8bxkXeJDKtu2JjbmAga/FUh8Kha0WQumYPkTNCf
FV2jCWfJvsQSG7BZ6uJfly3uB1HDGyQ6Hb/B7VJnv10gPufdUvAHKr/HAxs5IFQn
RCX5klh7SdAWiYgwaI3xOVydWcS5ZrcdXLEZrkId6E0xX40CQe0aMSF1aBWixsuS
tMgUjw6gEh0qIqOo2AzaJgbAVqN1z4bUphUSS/cUZbQV+M2NXBxBEAc5by+TzKq0
4jK5V6uDg36kh1amjglflMXoKpXToOrUG6ZDqpkzko5mUKQaR1QaExgU5c6dBwIU
UmgL+tveWKCSsZQNxfJtxs96CcFkDi+L85hZWFJ8Q7FUAx0ebPV4BNYi6Bvpo2JR
/BEV23sTUZfV6lQLXO9wmHFdxCGWcgCGDJSFn9aR+qrGXvJiLNENvPS2pO8dIjEe
Wsn76CI8PaqocbUnPdkFriykcase2PrdbLCalztIxnLyzRhKY2jTGzIq70EtgTxu
L7PtI6rxd3wYX8/mKhGBpuT1YdhXmw7Zq8mly0+AAkXuuTQixc794z66libHBg0m
UL1TXSTuWjVTC02t1axMr6b6QPuUClCepB5xnbK2p/e8H6AXTpL0NC/4/HcXo0oi
EWW5eLhbdVK3t5v0nW0quH3v8PCGrL7zXlPKuezJNl65GB+8Gna6jKHor8D1RJVU
iquGMGCkI4nORQyeaGxpc3OojMebqZ4T3/zhPSwy4ylx3ldy1a0aclavLY/0NEVx
23tgrD9kB86r65ErdeJHDzn1M2TPPoVSLoHkLBo7K6xKjwX3iE6aYy1gM6QJT4j1
T33EkfUWnLYaXtImxe0IVWr4fM/734FlYnjtfTSMqqMwddadOggod20owuM5yNRI
6e95S7Hxrhc2rhoL4fdlcIw39/wFD8OI6xk228H9AMUAjmfuwyZkCRn59s1S4aED
dfkv5QigQDApt74Vu8qSrfQccj0G3sO8OFtU+MUurdk5wnIcJH8H5md+SZUV2b4/
dF4yzMzJZgSlEXlNNZV4Wnt+9acKOTVQHYh+34gIxzKH8MeDxU9cqQ1buAlZp3dj
nfbFbH+Lal12VFKXx1KS+N8TzPppD9e4Bbv2SpxvZh4QROLUK6li6wRRvJMLcnkp
pUuPts7QhMx2kk13WE+6i1v3xoH1t+np+K7pDqjqlIQ4QRLfsDQSGw03d67fdc4D
co+2vDCrAsPfuBPhmqcfzRgJQpUK+M7wmh+mY92Toed+dB2MxknFE8zXr2ZugsOc
QKe7yNx9kkA+mKWEBpyGS1AVChwV1wzk/QAzSjg3v3hSy20Z2Y2OVffWqCm64u/O
YJs4/6K7578Rhve4U88jp22YcmpSMN/PHYr0mSMrTBQ0Sq2jyLzYl9wK7gP3zDnt
4VaEKOFq1VXBji6LlQAnMWNgPymajoyJqHuEOlQRbAlfLjPPt6pRjN8KwTF2HDPb
N5ZE8H4kgMqLbBdvhEOUjYfjXLxdr0azqL6i/J/GWF5OgVfhkxemNtTUXHf+1/Ug
jOP3rM7uHLZkHHC+2yLwhmHNzbowSYe668/EHWCANwHb774alwygM6XyAH3aebCD
GimkO9h4OuvotXXbrRJbZ7/EWkCi/4eGQR+z6lLmMQJN3uYuEcySi4eES1VSXkwm
Um9+ZRms9O45vBXwhQQczF82851XtJ6rklSkIjMmvUCYLIWeF2JUVC1U1gzpu6YY
fsnTBqmNhOP24oMJWbvJ9L1RbdPfRoXcGWkInPBD4wbAfEFXgg/unuRzRMbzQQ+6
rDIDUJefE/pbIQVZkdpyuEcqefXEEcxTyR01+ylqWa7Zks7lpheN3YmKfCX3Z9hE
9dw0xAi3CGAADWwcsE0QoFRpcOxR8UR1bxEwKAD4z8Vbd2O0uQozFUHx7JaDbiyO
CIF16XUwpufJc4qDZCVBpdDOIA5MkLiqH/RaWrLErxYjTt/Ta5oswbbmlTCtR9dm
FzEv3sUYzhCoHa/SEU+k34drbMLIE266oyK1evUqUAqArDsfg7XWGJW0RKmnCzB7
mJdPJTTSpOilQ8KJca6H2X4zV78w2QSX0r5t1IRqi/sMm1P98t/G8XGJIYx4Hc9T
xAVMMeEl0UqJSZg7udvXfcuyXq4W0pMtZ5Chxl6aHtv5lizIqsDtxQup2u5ns/WD
ZI+mxz7BjASXdF9Cwxu0muiRmOlaKE3cCUGCAQ0jiBBUhZOLuHJ1It8GKVHhhipZ
M6GLoIF0xK8JIm+wHvDGbaYEJmfOBbLrDYrQYV2REXFEiyWkQyhuBlkPhJZIjfCU
ahV3pe7zrs7rVingSOEYsF1tTr7eWjFVGaf1yiGKqM7YhugFjiucvwdIr6sJGK50
fkGMJDLYI+LB4ikOq23/kSENgp4w3QrlPg8Ze8577JxAEbbRiChgPsfRKgoHny8L
CjWnIOAzacDd5S3HeQ32hHnaKYc7Bo7xcT64HKgKZge+4FQP9lVV8mdhco3E1QFA
4tfI5bVK+4shNsfpT2NCK/XLhURelSXNo8ME90B+4N6uT/s2KmIwp237xig5Sub7
ymFKPVaBeu8ovHtj61DUkGcmlFpho/a+Hgbea5TBz7PVsgTbO3NaVufWH8eFVXhZ
bzu+MGYg9x0Yulb6jaM7pbgoRByx2HWJXMqkhj6cxzfOGQeeS02C3vmTxLUdsafA
Cl1iNkZ7S+AuKe25n3IWzIGzsIDaGM7rmZ8QWiPneUvMz2zlWurcZKCmoWvEvMjP
hD31hahX+TD+oQrPVeeds2yp/FfkRebtVCBsaz4Yrqq5GtFLZOh0CYdAh2hpRyhM
CTlg/XWVwrX4JKNx1zRzAObHjR2VlQSLGYeEue5zmqQ1GkFCAqWVeCUP34C358q1
G7a4AeKux1Bsf7LS0/f9l3+2q1htocDjm+Y2rv69MCf3YpZe0COttTbohPe8POuQ
ycH8Pxu8VkpngVZLUsggMHgqdGdY3/9MX3YtT6xNfAQaHbN7nV4OoJQoTkKzne3g
YLKUIpenMZ9f3mwHvpbwhXtDDi66Bqf7b7XGxastEiBJOTDiJA7wjrKzm/muKEjX
rQRSW9tEM4hy8DWMzlsnMxjWKtKEGe9eDTZvAVjX1XQRhrWQFiCYvncCrYFYq5Qr
WSIOnRo2LoecyLz3InYzjs1WAx1SifcE75ZPmUBCATPngD1DNUrj7hOU3QFHYlqV
7ZKvt8nuzConSwK30ld6SQRDbc+cMnTlV7KzoGuDdQeJEWmYCuOcDkDF8gA3uct9
Vf5uE35HipiWTUhIzp2dx3SnOuAMTLM/ARqVr7jLNs5/LHwD4Jk91Peyt/qibsAZ
zYaz8Rpsg6siY1uhF2LWINY0wa5nKXNqeux+LoCi9jp2caAh7Od6C6FbzOTn4z/m
cfR5YQGo7susr0aDlt1RMUR5J9FX2k3K6PxNMUuISIUdt2PLd+W9nk+tzfILVHa/
i6vuDPimKe+hbLEvQsdiy5UTx80j2d4kJUFOfhEHvkYLD/b5YQb2I3Il+WBc3XFS
Ef4/yyoNT93nt6LYw1HLP/GCNzG50jPYVUJqY4E9St76u42F4a1Nv0HVEoSytB/a
qdn0x67Y8BLEL4tbPYFjhDnHFLb6cU6qFFePYYXjilWdhfrF8o6v1q6tvdKwZF4B
3AH5UPm9QzioePr/Cm8QqM+vMpAso0HZI+Vwy0UaqKBm/AUhr6BENwaziwkUbzk+
Ka0S9xkWcpIUCyPb5ZdaSd+R+rpBU5tvEvQNZsCeF0mBjfE+jQ4mCDVVFb33xLLu
XCC6O9vw2HrbcMBIsmZTigjMuL4j9M627hLsd0fv4cw73SCCaE+40iTzZhA2CJBE
yfSNvmhnYbTccZn6cRRjV8HzJvN8laemxPk2cZQmlSbAijPKRZwIDuI8DLbhYA76
WRck5tflaCw0OfMqhIL4XN39+RVRWHltaG4sb0EpVP5u1ypI6C/NBuCl1JxkgM+t
7ekqxDULPDADx7eLkrZuPkxhtWVDMvBQIAVp1tlkllAKaYujd7G4KpLSp0Kh18AH
1shnodWVnt3QbpQOjhNFrAxXjQBFZT8gtTnYioSNfIYZJP6hOlQqmjNWn5VBLcHP
nSUhKa7w5GDy9xrXMJb/ISf74SIXFYY4RvhmEboc4uMUYMpBG5BFkaRwCaFflR61
zQ9lxV8cCKa+5KxNsH7Zr6BS5P3Zqwh6JCBLtPlr68WTtGDJ3y6NirxZcYdxCOkg
QiHicmB25TmcRohWHrHM4BqmlJr1oh/+djSNNhutotmkVtcCcsnzSh7Kg7adOxZP
xr1tOMymwGfso+NWtmTceL4JyfaI+KKe3fuS6nNxxjYp+mYIycRCwtb+793k3JBl
l0LV4hshCCcjRviJhvROtyULx/1h5UKn/77HZqu3o4cZ8S9rUyxjqKGy8A1aEf63
AlqsCHW7MrYqsiQQKzyQBul+kX/yZPtECatNBJ/nEysUAoxaz6K7Xj0tKbEZKibQ
v7mehscinzq9FJvfeg8erocbh3XOpEchYEntKV0Hof+AlMZD2StteO4RuB5hzidN
7jTkFgcgVc2R3wGxX9R0Jk0XEUzNkDunKTAqvaq6a17RFRmMdLfi30wC+lGXIZMk
Rt2HDfiNtOYqXchiApkFJVCqHir/CbdnW2je/Mp1wTdoXzRsnGh1Nfrml1A/aKCE
dTPQIAnXeRGAO81IiD8Ene5CAr+T0MiKOllVp0tU6bH3Z13POx/UTQKWhoiGqYd6
XlulIaw43wWzO9lxwD53DAHp+Rsnitd3UPCslzVfkrzxbMM4ZdDsPBIuysvUf1cp
a9cbg+yImvhYwf/mSY1BI03SBg9pr7lQjvZf9JJEXhjjHj7NunuPg0DI1Bj2fNhv
cDiHy2BlYuPoW+vAKwzssFq02quAZQMdvkW7sh12mlN33h/F3EaK/ZIvVxM1MKXU
lB/cqaVYXsIbt2CoXcMIAGId01E6v3RU90CjgOMWn1ThMHqOLC7eTqOk2GwuB9/m
XzSN8u5xEsUWMM8WCwRaKYYS0W5LWQJcDJdw0/5/SywU+4b7XKot+bMGhd9Hmxzt
VJmENlvB7Kq/0n351ftYxKsKDT3eCMm0C4pGWwCrgdvMg+bdwG5K6EVcDGPBmhaG
4vddnKfS8ZEPqaKAaCN1FlBUtS++cb2/577pClO2mPQEYac/Fou64gVgU6gA/GbY
vfp6gzaMkgxxEXL7bMTlH3Du4EAkPmBo49OPpcT+f7EbRqghSkJQaK8Sw8CDlWo7
505OPCdrzsJJsBziGMT/idQ7xINauglDbk3U30esqTs48UxNrQMupWVYehmHJQ1/
orLaTUlwysqpdmMqTQLa92yKWCQ9fg1YwP2FkPvQA6N8dg4CZX27GDl7zVRrNQLu
L2WMRKfVM0RSbzLALtQVQNUejOTj6tlXkd4LIq9jGO+8gQrvAnHaenkWxC9UwqU/
OI+ttPTwx6KVJwzT5bNNQFmNPgrYi8u37DSxp1uQXezvberZe9bqkO8j64/mCzsB
JIOk5PxrtGDoTNJbTh2KYbg7IjzFjcZWTcn/E9JbqVCMZDkgLq5fHtJONYPdJXO8
QEW646LAEzFoZIfLvD58o/QzmVHYAYNAKpVfoK46NfTS1aRr95poC7Biqk+qXiG0
rTdBWa121xgj7mkD04mxc42PnV/I5pobNHJpkUOod7DQrGQz9hFEptyS9r1SjkJc
17efGepC3To6BGYucmFwyb7gASqRmKoGrU/v0OFeVHzvKHqQgsGVEGWXv14PS8W8
U8q77YENP1EM4OtaYlfa1+eXKTuU46Q8Tp17CLbp1cDA2sW2g7OkfIyteiKGoL13
F1PUEZjljCY2rlFVR3RJUHvNxG4BpJ7OKLE0ZMRTiReuMmhBcIIkICiGfhZ01Pmf
CoIvAaEeB5eMQfI8yNAK60tH1Odhgt/Dot8PS+2VLZLpG6kWX1QA7gXgM8mRgore
AaZDvbT+q+ebASz4Wbls1mGOfABWaFD0LhIzXuGUc5//VCLi9emzfYxoISph43IE
vTmUHl6OVYBmIcpHJtEcY1hUu4ci/wuAq4OMLZhm+WpT0W/Dd8nFhQzWvtL7D5wJ
QtvRQakM1VDyG/7jBN7/cW2YjmR03HJHqgV93PkloXS6XCS5k5gnr15F1O8Et0b3
0VdxnXhn9g1m1p7hD9+T9BCQyoZ7+Rnh+T6mWTElBHCgILKmImjbCeihtQURcohm
ipsGoQrTF3zXp5IeIT5tJFtKl+Kp1IfSi/gw/ft0vBnDOdIec3Dj4aNonNoO4ziL
nxLA9MXO3gBd3Nh1FJLR+0ORefzyX2ZZt23TTeR3YJvdh4Lyu85v+Akf3yrrJs9q
Cs9lZkENLEGTL94aurcoNJRB3Nq2UUsrJD5prg/jKpoD931QDTvXWCRwqO09LtmR
2A2cQh/z3ssZBQvfxMjhPdJEiVUSHNsR2e1XztdIPahQgp+tJ0bMYEZrQ/fy0s1O
3pTi9M78E60baCKTWHnSvSrufPzgGj2T+waK/ovjA339olHKFZpjPS4xz0Zf8fsB
EmMayY1RwnmHyvu1hfGVmCUgiVgNUaHpxUT4zYEsIsMhrICARSCW0vzFk0CVuIkG
x1+/pbUtsGbKcPikViWpbwMe33SytqdrYdl5+udRFdqH1qaEbXTlanv4WP4LFf6D
IE0Akc53oGhGLgM/fdN4whlpmJ2YHYR/fZo1oowiziPrMf97+u1zCCPgZbqNBhtN
GDKvRBznE7+pwDDjcQ0b2fveaGJ2IGCobrISRD15MeDG+ZD0/Qc14iXyqHsaS5LC
qApPawwPHGa0aPWQmROvBiMbTWWcHPhH0pbRBIqvSIcFAt4G603PMy9ZQtSyFkmG
jb7GcvyCoNslWi9f2ACkzyGzrUjeQ69dQ4tzYLUBDM8AoRSu2hXGXGOppd4alZ0o
34N/XXWYySMZfJRjQtmZW9MM9LsblnifP/0tDO8YBVzukAiJmzizm7U+O+ZtTV1T
xdoOjL40caN5JO4WHyU3d84HfuN4CSsmX8BHfMjldY0tLrQPF532f4u8VLiYjSW5
4wCV4T+zL/PMV/EyEKuw1RmIDv7hC+npyhv1m5UkHp3+3bz/i63VcpLT9m5ZYgDE
Vx2JH5oSKVfmQ/7BkKzXRkzvILjPNOzG/YuCOaqyhDM+lhZ6xMa56vxupgZO/kYK
9+8FzvfR5Yrs9DjW6DFwv+CAApxbo6c+YKzfs9xjz/b7vuchZ3RPCcA6Pu/2w/X6
3/j132u5yKjQNCMvb+bvSA8iRJAF6gVO+2p79rrfx1PNPSU/sVJaVtIQu7AuBIJc
XBJ0G32dNzAgohqPbS8CwAsavTrtNKuITU1FNf9WFEqoVqL67Qtsj714Ystg2tng
i4i/+ulSnjQCSwZV5NqkXEn9QS0tQX978TLY0IeSP0AIUOmZSZyM4gtg4tqZmYCb
6Ha/dvK9KiH6sxZK63W9tQcU1wcROiCRnhrCaKUuYq8PSwS7UlBrP92tdWIuL4MG
GI++HaAVV2GRvLSKVJSUyWGMIyq9NDeAv1xCTL/D2l18MJnb2oN0nNh5ozXJPcmF
cR+XGrvYDhuUheaMGtSfx/ok81PkBKMR3kuGHneUEArdjkcGeUFWhdVHwfjoF/j9
1552IqnJ4A45GluhkcOJHhP/G1EwGTsXueK8P+KzS2neDoSr5MKxHCviWblIgdXl
Rlwexlm+/n0F31IFbaKgbmgdwZal8iMkjS7R7F4lLdoVW6HqoVW5rOSfjGi1Xd6m
7O6Cg2Lz8/5lxhr2vHVOXTBwe+kCFLAUTLINgS/nOioT+Data+s3/u6N/EC/qaV3
Yfdw2xTRHJWTPfGlqLhgVg3EFj0ObcAGexxg38wchpGdj9AaQv8PT2npt39Hh++t
uo8iEyaLaNOfFinNpLFehdMSctYVMRkpm0mMjkvrrojdB3dVahGHUyIaC5K5koNc
kh/Zlhwxh0iO/O9t/xUuD/ebER4cSarQjV4tHYcjw4LXRJ2OXFGNOKAiQ1wMrd1c
9wvLVPoATfMo6bPG44lP2CsNcwIqzN2ITHa2jyuyAJEPLt4UxbTUP+wQNdr+ohVl
snvbNTZS4QnZLAz+Gun4+uEDRwJjk8E10izAV35CoUYT5fNPwU692GmuUj0xIZtn
+4asDsJSrcjsO6v5JVxiqb5bm96t7cr3S7thWyDb+x3lVBoPlhHc8OzePz6bn6o1
4gI7sFaJYrik1jFb9eYng4VAr2r2NSzBodwriL53MOYE5E9yFHk2H2J1EI9I/H1d
u3K/k6CfvkSe9nY9OrChpJET7OgUcgsfFj/G34JrcQPfFOTZo/Ta/Igq8RSeEBUH
0ysobE7CzcpqcbBNoLxFilAwFCoDnMFsGyD4DBOVM6UkHWvRyhK24ll53OqjtG8A
4SmBD1P4KmY3m7SZ621DuAu4joS112UXlkZT8FkG69NfW6Mq9kH+g/GBuPDt3gch
+XiNL+LdtyqMsRMA3KcbF3NnizW8/IQI5ETjI2bEtNq8xf/3nhAZnY21QdhGzf9d
4TNkcOmWA1lXzTsRZafBAbkZ6vBloezEp8dxCNYK+j9/ftgaARGRuIFeFIUGJ4NG
EKH8/lRhwAQ8LuP+t2Xp0iKRQYghNzqACoBa+h6Skzf7IPDjYCa0VfpuluqDE26P
PJMpKOiybs9BRMf6lvQvO85YCeFLNysJW6hiGAHv0VsDUbD3AFdPsW0ZSH8eZAhu
4M8R5hBUhQn7GJaf6jGTw4Gd/VBiH+3xkp/+AQgx8Mdo6eU7YgAJ2tRe8WZoFFGf
aB5rJMLyAivTT1Zn2WTnW2vywyXHeRsJdVEPx0nSxwx2zMeanUndzOSDVBT3Afey
EDNf6ODXx6dgVQmgu/dNNhVjYq6S93Y4imhLxt8e1Jb3es4JYE9kUrUju+S+Lll1
+1ELCqDfVI34gDAylisgQsrTsQOFCPWzEPujE+bnm0RlhBnEQh+n+0r8mxeQ/2mQ
w1nd/RQOaFpCstU2sXCtmEtKX6hue4dkSqZ7/FcK5VY57gnkGtabh/EmksIqEEml
u3v9yVKX4ELf7t3B5+N8cJQmVK77EM/FN2YLS3lK3Z5OIUUAtyuCT19ExkU+e17a
IWufz8TcpbXSQ005/uH1cIFiE5n2Xdw5e9VwK40nZKINU21tabYKj3rZj22qymgg
Yn78cLJsEBDCIqpBgVyYDeKelKX25IXSfsFfZK8WtbJskRAF2ZSJfsf9jO4iGKDe
7OEjNqU/2mEL/amhkBtOMZ4vUfT9PMcwjYQuUq+qjBCXIYLcd6yMg/wekLhvYze9
9ykUdGfuvHz4p7DYVk7Tr6XyDKk7zEc1zunsA/dqZGD098K87Q5MtXAnh09mSRa7
NF9WvQHuuzg22/WY6gfVpQD89HJTxHhxPKFiJkZKkq+96fNCIbMds2LTV/Ehv4Qr
7Kx3TRkgcpc3hUCYXHc5qlm/t9PY9+I6e1+FwTTXwnB8+rcLit3S2nDWVhm/qmw7
qpK76JIFdmikO0vEOGaWZRN0AXh10CbBrf41umBzu2K+0VSF8Qr0ZUDH1yAKCIJv
L3qfqvX6mMSbvSv1249cS/+IBC1URGkLiVI1gi2COqbUMt5LgKGKi2v53wi8iGlV
mMVIdHgQ01adxhceRy3t/FVYn0m9pPzqXWE0aGdrSGbWQaCeDDnnD6DlImhK+fdm
bPkol3LcmKXelsiOrryN5Q5CA86A/h/kzprIcJ10VzmA9fT7H6nOcliB2eSJ2Xq3
0PVlR1oF/GRIabMWZ9Jdqdkal/aFkChzQx4cWtWYEUydGDn1M2g8SapAEi0tukH5
LUYY5AJTUOne2IaHaitmLVEWg5EEF5GukGTvnEQoAGZ0SBc1ogCoJ9eP1rIWxR2O
5O5G1mv0B1uGTeNUdT7Y/CU+qkyLzqJFwRuOadLlKG5+vYQfx93mkOXcAh1QzavV
JMwxiwEAKHInyYiA3fOS+f27wBiLr5GohpPGuGDlg3WycYwc51jr09jJgq6PUWbg
Dkd6CUGMe4wD+LTOVXkBbWlGP9l0086r9EVrGhkN+cw4nIF67Qmda1unXQUOXKOr
Gqiin+6XW8dwinXoXDtjk+4pE0afoNDDPHZ8wKqA5eVZVYHwFuXYSrNSKo8XdA3v
U9/IcKfJlGA8g87PoyZsMpd95WY4wHOO6iKEFaTsZzbSKxOh2gGw1K+kNCEAqr5z
1SSlNUTG7BDBb4PTyoS62Gb7dcClpuHnej0VfOx3NYgwrj+aVHHD0heOrmxn/K95
QywyGc9T1jENoi05TxwJ9I2o+N+Z6rig1rK41bsczW5kM8y+HH/1m5HLkEKhaCMH
GURmol3ZaS+XlmAnMe2GOPdbmx2ZU/SrcpSZqo2f+u+t+G7ksmTAwvnk7xDNlbiG
GD1gYA+wcg98UboC7SPhZPrNMZGFgH8md0k9tWp+MjL1MvIY1LJDom9o+6ytUeLL
ueTMBKmzvHb8cy1gwZj7/StrghPQDXI+GaT+65P5IOntoBKssIw7YleuaQRhsbEr
HLp3fGKsC0CzUK0mV9CMxpVg4AzP9C8xfMH2JVdNncHEnMe9mvvwk5iheFpYZNQo
BJXlapR50Cfs43skZAAHlEpDst9L3wsubKJog5w0r12+uhrHcMkH6XQqzC6BtVrt
+zJFkVs7+n7DGu7ejL/NOqEd+WLDNv+06tHtPBMBI+/wftHfityXS3dHgf6XF18s
yNxys0ROGHc/j4dyoLQ2ZEOfSriGBmU+PIv2R/pfPWAxgPuEnE9tfVqp6nED+f9R
eDruYUrTzpTTqln2rVBSrq5V8ObMeH2GC4+s0Akd243Um7JsLngaSdAqLTzElHd4
0Pj1d4vqaAUBr7yfxgprh6JDS+TCEvnag3PsSKEYsaMbPl+CCXJQ/ltgyS8FB414
eyGfjsAurYzyUwK9pmKBPy91h0WEajETJD8PFxA0bmCiqXbk5blMLMP34Q166ojd
sunF3dH6lJP889nuV+6LqygggXH97zmLrBs9FgmnZc0I17S/ngsbmM9WMRBoUIDE
wNuGCG48lzT5Ru5C6cSLVz9PVz0caXNcy2MIPCg+UWaxi5pbPHNE8jmSxLw+/gSq
yja0nDGp/nf3rUesP7PL5DNifyh3d2efMMGWbKPaYc7d1HvBmqXq2mSAjQ2hKF4m
Zf6rpdTVAZaOWfaPZ5WlEo5q4BXbUwIJDqT2xQsGruFazxB2xAVuLqvfHdVGoPjv
1KW4mWciUxqn5zaC6LZVlPgG0sIolSoeJjkvePr3nvn2vtJsCfxdfIG5uqo5FUTN
xVL/aIl6vX8DMKo4VMmxPMat1QygMJz0iKoRtCuFtCnBkMKpcM4T4UpR//SSmU2R
t3SgQ4eGZd8PGl7VH7gHRz3PbHxijf5/Gnhn3IM1P1cgXgXD2JUMzJXOtBA34Mcw
BPZr2TgErf/DAZSrS1ccg6jtDUhjcjYXT4lRtqJZdMEyocu62BUnJ1rbw/fVzk2U
mcoeQZFeCmpfJeuSatV3TBgYpgNe7nm0jy09MfgLioO7LeJxUYLjjvTWCTVCLfAl
Zl3rO/y4mkbyhIyG1hcthEy2co9vCC5S8Xf4TtSQWLAtc0fa5hdypmnO2cmF85Bn
ZAZNE+rtmfpR1n6ihIeSU9l85I/ODR7iQZXUCAEEs5T20i59bv0dDEM7vTF7aSD+
VG5ZWUZlkcvhDEuvnnx04EzA1ukW/VbqAgTYEO1D2RyGoAJyMBtvDP2H3atJU0KC
QGo5J06d4o0xI5pg4pWpt9BwD4RgC2XAsTJNa3ElUGOc2PfKj+SZzfpHNRJ5nXM7
SqTopAxhJihZ7sTFuh0lXYcV08dLlu1y+SJ7u6jc5+nuaC4myze1JAZCe7Hs+3qH
OWrzgIjXe6xSN0LQQE7hyPj5BeHxaNkuZP4WN8Qx4rUaCVAOqK9QQw/HnYSsUmFE
7SZ/C7BAjvoqIo+Pu+I7HNeyev0/bNNl5gAxq5+1eX4XSZYsQRirhBwon0IbB/Wh
lK+O6s/P53X9Q2ySaXX8FYoK29xGj81QuRoxcLN1B2XiOMzMLB/jl8NeF6TS9Uoi
Ck0Hh9QGqJKZ0AY/bWcl+SD1/t7NBnVWgu0xBpOtdS83eo+Rxci7EP/gbfByozMa
pihoU4lZQxIDnidBeT+CB/YLKtDLr5uXKRx/qtQFlkOSvaiOr2R6/5n1fTyVwJ0w
gJl8n0PMXIk74NXoQ+H9SuEqh2Axu03i7cOz7tWwYmfq0Dt8Tw6z7mBk5vPe5FjL
ET9UK2FCf5XDxT5KJXYXzWLciKKn0YzR+CvJeHOaREoskgBwNzxfEvrVkhvyNVwz
40GW0TAKQ7jYSUkQnlfSeAIwVm2rOUVKmgO2bILdbDDchcI4pg3T9+i/oMxuX41w
PTEOyxvCYXWSKFcY4pjmgGyhyV0iUoi6dn1YCGbW280grOFo0D1PTnNlw9iC/DmI
D2Zp/HKrV/tRzb6ViiLlR4TA1o7ilGHMOi7GYBULTenslUS5rxjT7gtLo3qs0ZwP
mGbbBgIEApNKCZMlSZTconhnuw+FCeLkQXYuj0YIp6Cz8bx7WZtL7svnxxpZH9ux
+72i52etpqFmVsoF8tZP0djl77d5FItvUmqjp4UbozY7zSsR7UsdZrAMRhuNAzbn
EJjZUCxciTBF0czMI3+zeajpDB973wbUPVLYCsrrrVgY1NTfUHIpJ+XyA0qh+cJd
yWFhZ/z0f/MsK7XpKkfbiqD3UsmypaVGgKAmzIZnNlvOjlGDg3dMXI3fni6ER8oc
4m/zYTDoQOh2ddR02fnjS50iXBOhY8Zi8LTEuV8H81LVJnnLAPX3JesUK4tkM3Qx
wNngPHTJrQtpV5AjXltOAYRGRizXCu31qpLiu8VFJkUeL0xrQ4OZMOzPnSGoXkzd
jvL6ukTN4EHcV+SBMG92EOqV74HBu2h2e9HpZE49hl76Vbu2uC+e1W7zzTtAleHs
lCdeQDZu37w1lB+TOoiraaKJqEl+lqI37sBWBCb7WmolADdsya5G9BDc7sva/bWP
J3x1mq0mrtXsobsE1sHRJ445pf3Jl8XUi5ujnvYI6QPoDUaZ9hbdt3kst7Emu1Am
BgXdQYq1r7o1/g/7Bm9ETzfuBkNbVAjVWr4xlaYYLUWCFugCIVquATpRPIO35WbB
mQsXSeiAfKE3ITJXo5XwQaVewZe62XfYWPjDGyYJqZ0PoxiUUlBv5tb7UNVshXcO
QXKZQT90CrulYM1XHyIjkK+ycmG4JRGNPwii/3nHEqMwfuyP0WP9tcyqDsOxsDJh
T2BMmsAArr2Hm3YErlySfulTbgiX+Wfrpv4moK+NkMfUJZwIVj9Jx69raH1CwVzg
b1MJQZfyv+AQuWysWqYJcJMV0o2yYjn8M2VBwvSW8LlCeyQIMfOkoTzmn0M89cwO
CApf/IqcFSezRiBa3iNr1/EMKsM3O1HHqHQeGfld2UyUGXofZcdL5vBswumSAkdq
UCE3k/XwLW9jZ+EJNdG68uOmEU2n/Y2rZOMI8e7ec9zwlQLlZ0cwtsbDXQ027H8C
RysINT8BGClMmpKyEDT2bOL2W+ftp0KLmJFIOKkF6qpoUSSoRzAz/l5mVsx+5z7o
YB/ikOvImW69gLtNo9PU++22nzl5uP8HYN5sREGTFWaznLMOtS9u5ApTW15WuDN/
dvFSINk/4s8hFdf+sFEJDQS1w4KzI61rTD8l7VxFVw4CDotgqQQcIg2NdhVcJkRz
kLZh8y926M9mNiX5c0HbmzSMKg+EuP30NUEi1yqCyo+da0qgLasJXPvmUe2OXgv9
jrheD/vBokiC1FlRz+HkMeTkLAiKKBM+o84YKiCcF78oHSaRLgOYYhZ7D+P+tl9m
rx8aqihJ8bJnLcRLspU5/lbwxbRYObHMoKD8RhCIEd91h4AHa9RFcscizqIfMUeb
Dpw5q3yXqLNaZnCxafKlExibp+3JcIa14Xw1o8pmIjf60UBYc+p/h7GcpCsbh0Ki
onKh+qNwlbsPK7D51qrHDamRtLCZWT4pXheXoAYTsZrizzWBYCrj8WowHqFdy3pN
Fo2VcmVMsY0CM9o93oX4Tb3Fth685XqGSMeZQqaTouQn6AA0OtUHFklIwV6Jkbog
CDJiRFYL0D6EnkEBtNY8hRpE+tG+/eHI6KqLWU/BZFhhhJcwYhOi3wvhfa7N5lCu
bv9IaumB4aw/VJqKHFVbT/BrGYNPo97rs1kJ6vAGIwbyYI3kiokNAy6TcF5Y6bTi
1Pzjrwh5bI832bbcA8Cz2mIa9Lt8nAb8QEoq9rnPRsIus1gXw45E9MgDQGrXleDE
8R9pxPQQnC6iWsjHS7NbeG+xMnYNTjU/7Xcv1uXakTrVVcNzXwbpV192Cw7UVS9C
fEvdWhvT3WANcK8TV/MhvegJkCHwi7E2ArnK3zydm6qWPo1ON2WOW/Jgf7PhQN1q
NHeeLMthswBwVTqZhIeUdjxJIuiSIoLeh2+l6jef3f45IS+He5JfZvG/BsdAB2Po
QjJH5IXxwKoVV/SaTJDGvbCJuUqBMC6biJsXQMxmEnUlE8DZvtdqCNc7Ux7VeGyc
uYqp+ehkNRxpEmPFhaY1YugHlwyn8p6eVXp/B8pOfSJ1e6HPpLPaD7FMqhHZU2/f
RzNdfULFWA/WcVFLAvpjFvAid0tYWN+g2FI2Tm+IyPXoNa6uLUaREPIxsPWCpYSW
AXhhLi2U6dmFs4hum3sdUbuGFZevWkbKVLUr+4U1j4NwqOE6Aa32tdgIgOAQtA4F
KlwRLIPZvwJdEsYnMD1nWkQpA2ruZzrHOAwLQCcf981wIi9D97Taq2KQOWsRdnKv
Y/qKucJAqI93rfIApgB7SfwAz2I06El+jcZQt2rL4lR+Te7eoFBHWlYVyv4RSKBp
pQ8RnjSCXUVUT5V8mAad4g6nnBxYyS2zc7x0fQZFJIcIKE/P9EDvvOaxxWDOEV+c
Y0YB/3eFFtGaaoM+8AbBW9l8LqGXk7xn8Yz6CeBAgC12/cs1yuMkCyLnPHSiT2ff
V82qc/2G5SOPsL9fd0ulsBy+tbxjwepLdoYayG+/etyNYw8LN9yzJo3rEHRrMlai
5c8tVTNeWvqz07jPDIVoa18gqLFy3auRr+Cdaiw3aDeNEW0xHGD0+1F0X24D72/N
kTI33wo7FGShKCF1wHu/h5mY1HJ+acJGDgCYAfZoMY/2X10wy5mhltfoXQjYQWeO
vS74uulsekO7WwaWLfZOMFgBYRqKKreKRufU9a8r5Ow4ybsDULhs0xq8GuB1TzfB
bNJB6a3BafPCCzEDslL5Cw+1QObG8OWjigYjC4jxsroJBcXakncsXsQH9cxR/Rud
EsRnRrOhsmVX48Wx9JnKDaB7Zacac+/rC47YkW9SqJL60iTjy3YcuiNqMaBMi23g
UzIbM9nYihYV0p4Mw5O4YeKyD18w/UJmZhQe2p2C6dk45DhRcX7BNMmT/7I0Y0DG
LPxmOjuyRKDmSdmoAvx2v1oFDjVYBDcy55GuETjaphJPMeN/1K1msRXwXJ97nYpi
w4WUpT0Vuv9C8pYfWijYQE/eGfqJj4oClAeqPTeeuRAJRNP2HuU7avOcKCuQZKZU
LN/t13ddbg+r6EZFLGKsTj35bkgYgRZhfIw57Lm5PxdRfvHE7+MyPddutI95j/wz
8Px9083ri08byAFXmO5w833c1+r+uhyOaYvQ19dqObHK6xaXFDIz/ICHnqVmlBFo
wKbqbczmLalXIb0MywW071ltMOI3SoNYpDmhay5K9218fCf9oRned1ORNRdVJ6Ff
7O7K9+0eFIP6VciIu83NZfFKFLcQXG4+JBxEjbKmknwxDudK28udfLKze7waVGI9
HNBRkGYEg2bv/65EP8MzwsIXk4ny1khGX+PUsLbnRZ4cdbRjLCCZMr55oJihH7aO
jbB6DWPO4KR1v5ZMOG1t5rZXMm45QZZSWoNsYqAkHgahqNfZe+bT895i9wvGs5bn
3sYvTMGKjL8x1zcpWCYwZFOPi2+n1Vcp7hLkUnBPKO4+hOIwE7MpOQHk6/NDnk03
UwuJRXJz7W8lyuVSizfFIOya5EnzFjssNaQcqnguQNErO1bpQxN93YX+TJ94f0XO
D+Fy3R1iBKM806od2BEghLVAVDVLDGoR3CbS0J1bsKsv8nIaY21Lx2bCkaZJnNnB
I7dY5Qon0bUT7mJIiOhHuktc2fKhoGNYF/VFTMoYtjhU/6/2ULC7aXU6C3csw1sF
8VTZV8TRqrbcUaK0nhblV+clyNhJwqhkp0sXW9G+md6aMVZkyaXgGVhoiugyo9wO
UV9h/6iMetV+XyAHpJVb7Hv+N4ZT2eBddwBfApRkaUxyxqMAe7nr4j7WVtGzSVPg
ine/+DCBlEy9i8+3JTqitBZGGulyJNM1vMEXgV7rVw41Kf31+wZWSCoI51Fcwmxl
S+dn4RhNp/pPc3/s7XyoWFT1db0L8nQ1C0DqlQQcBZC+zGOBhJUqt2eH+1kKFLqn
M/QeUZT1MOdmcJt5QrJp255GtxQEMJyR8Yf5X8y6A1fTgPsiqmoLVsqnHvKoIyop
PRYof25h2AMEFAsT1xKV98Ks+kUDVCo6UU8lng+1yHXSVlnpZEjctrW8UJgOztky
Ca1VmJuf1Yi2nyR6bQIew49iBhL0Y7BfGuAuRZlk5fWnBuhFZH7cLFFAu1EvL3b9
X9OCl+Rj6I94ytBpJJJwx2OevZq+DMUKr2beEivFytmpLoGbhB0++jLFYlgrRup5
ksiBmCnG9JqyLGYDAt/u1rK9o4PkF0lNlFaqpj/0QWdQfhh9LARU4zdl6rifN1te
ry9im0MNvCJMGUBIiv0QRgsBYuUMojVSNSjVftusIaIngmbimlCO5Dg3vllz+erG
6kqG9uuemguVp33Gzn/MmlT2q4Ua8c7yRMUcYSIdJvdzL/HSNxuhwn1+IO4B6qH8
8b+ab2WPA3Q/FwOUL4ugKc5Q4yZHyh04MvsFa5Z16Rn3RfQcq/VAHJC0uV1LHMPI
6doURuwKPj+gf0MzKp7j1N8iuerf7x4f6SUgxI9D4W1ypf3J115ZZnOD3t7IP7Lb
/D+5av+OSdqvEAqdwmz3wlg2+9UX0EU2eM0cUNFVvxc7nmWbKn0cx4EMPDJVxtlj
cTMzWKIs03WysjN1z8uDbLRuexAguI4seIkdPygQd4ZnT3hD2qGY0+j6JH+Q55fy
LHhAUR38MecAI/kp3614r+gKYrdj/72OSFAXzRgMcJI1ESnPfID/cSxRNgs5puPm
dlDroM4hSiCi7eS9RL3X4d91cqXht2dHAI/W6F8/prGTg4W5NFKyehF6DkS6v8ld
qptFeXvKb5FPMROuvaIMv/9zlDBf7Up4Jj8kFDO0v677FcAZeIEn92qa0EORFqnx
xujqE+4WzTkHKQzzPG6LZHojA5kQen1tcZX7zUQiEl+BxDSAeXOi/TgFe2zay5Ib
Ppy5WMbCx649OvrXkGwpOuhaQCwNu5C44IRQ7TTx984OeSHqtqwC/U1Y0FKvdGgH
zbtaTYhWoeLRRq1J/lx1P44VHv8l07xsHmBcBi0qr6rgky0PWyOHOsaVBJmgynmL
ZBWN15CBr6tyv0/rHhPdqwkpH7iLsUFvxeZaQ/PYbz5pCUcoC09vPEfwnNOqh6Ed
yDK4USPJXqT53N189jchrYeHbcoZ1ALtcv9863hqcz+eIWcxMH+e5Lpqd0J8o/e0
Z/CumBX8dioAND113A28TRXKk+029+VW+iHl+yspJznyLx7AbMoW3ykCK1es5WdT
uzPVmPLbp49IySzBSDrw6NcmdyRiSi1FFQjsVTwjAjml550jxNFqAQA+mc1UPva0
hzAqn5yjl0iY5VQNmI+0CGYDKMMBQccToV15tv/+wXFu8iD4vUohQOsE112gTWjE
v6JZxN40O0YHya00b+2bytO+byS3GYrFG5HfGkHucmgj/MJuYnQr8qA78RHSA8on
z8BORS+h5vpbwC/7EzaC6cvzgfMgWXN7YmzWbghmNU9K1S9XGjE2Tz2SEJsAaFtE
zyYhEB5MGSjy9XqID58C9FJK02E5IBxX06WSd5uAAkULWM6Iysk05aTYwd41giPc
9fowuNXmV3A3PU48tg59l7iyAiCLyMxGs3IfbM9aazVV+P+QlxV3gGvuxkiNrYwn
WdI/ybXs93nU3+zBrZH6h8lviItsFXq2ZvFvQliSzhFmEYBlGN3MOoWl+phDaxRa
9Pn6pVmdg/+itlT+swkoAZdW3MAvkl6lF13VJ3wUPOtQnU/lwMu0P6yha+d5WsmN
TRd9mo1CjgeT4bihO26Tv8b+ILrFJSdKibZ33PgMzMaltc9knhnDkx2PRQBA7LnW
RZCX5Ymi5RdCjSrZhuJJDJhT5bak66kgkbyrWZGO+4LRirXlZ+XOmWGcogS1t4nF
xf/u7uG8sHrWZqM2RXq0iGAHjvfoP80vvlyoL4CK/6gghbLkSUtm0IXvJWXSgBIE
lnjy8ZLleqyf9xviC22TnFbIGuA+l58f4v/DeflBCLQXaZNm/fbJL7tL4PFYRh50
kfX3uKOpHm1Ok24npCh1LgBi17aZ/WH+XEtPflARMK/oG2u+4KLdsk6fOssDwcHu
PrAeRtU31Np8u0jkXTpf0Uammo7vimMZ3Si4b8vV1RLlK9d4d+67SSvcQnA4RtRp
Ge4jvMQ9cxdsWJ3zAQcJiBW0+chP4eN3GD6KrAtOr3E+OfaDBjvO59ELHeYYJs1s
W5xPMFjlTNzAo8Y6fng0mualnoub/ygHHAzqGEVT8qpWUwjMYsR98Tk4Ti2rFkDC
xz1Ngj73LNKmC+oNMoHgZZzV+z5kH1zAXGFJj2Kw53fLLFE+QDTd8BVWv8dLUsre
0jagY6/5Lx1J3zAdcmDVfnp1LDCHuUzLlybQjzeYhc5JhfFIyQJgpfsRrEXnxAl7
WtCh79OZM59ilZpglk2oJNA3UwcmC6CQyeZyXAmzs/wOvERAyQhRDiOqaxppwxyG
IRpqgeV712EqiruTlPjLMvK4jO/bqV7JdPeAW5XZpazgVhMQBtdhDTMvT3cHlu3Z
7UaXWtciDYbCPfecsnii0zUYRc0U/BL21IXW9JCaags+/1rioomrnnu+ViZBAJd1
KyWnYHeJc7kWATLgXeiE4IP0kIypuyGT2YgCPSo8l+KriBBU7Xy2YrXoaAB3lGqe
F8O+loAdfUzfVcgDRd8WU3zrYSIPvVuOLH8Arr1Bnj418dI6gvV/zMD3/MjhxTfp
E1KlApNb8U4mZ8SUCj1qTIJAjnWt7ztMZ7s/Q24V3fqWRPXfQWFlsScx8OJ4kRBV
NLqFiBVblfo1K923S5p9cfVtTBkavaqJvmKvXamrrrpBhu5laluIbdSHsn6h0rqY
VA+UTbdhicI1scPqolX4Kc1CV0tWaBrwBF7Dob+P7jExbvFEudCUGNHRFJKwxBCU
JGV4RczHu/s71OLQi3ixFYed7PixSonk0B5KRW75O27j3vRWA9tVEGK2ViRcGM3M
ztdQFJZKyyDrcAIyVnrFbZWPGsGa9j3nyPTjRRDze3dEY5nsGGLEV8KMWx596hoA
lC3NO8dnZbloVtdBbDenkaJcp5haFCyygtRaWdyf3y6GHMotMPvpW5lZ4BAOwqwC
L/1jG2EMLfg/nnN6+RUeISJzxdHjPP0bX6ph1cxZ0tmsisYy41XfBjk1PNvIB0b/
gUHgEro5VDYSIZdGKe0qNLOvXb+pakGmK5yObfY79pgDr9Q5JlRx3/D+wUE1LzFT
0wfxfYdxH3BKDREQQAMb9D4plAWhZoBRkb55IHS67hL3aHZLWhcVX0vjFvT+wTcM
1JRePi3Uhz1N6azOdOBa8u4LgLw91f9tC7WLPRpl8omNGmjNMHPtvi4Kd7bAUc3V
BK4Oj4kFcIZ8vl3UawEzf93vDnzTieNvmiPTGqsMNftfEZwrrwK5pPrVx8/GmQX9
C4/AY8dpI3ZrZfczrJvKYtb1lS90NS/VAeUjI3ZezUzRMVNhJ27cl1LhJVr/oQ3Y
2tTQHgsHUVl7w/QLmiUOTlwvZuFOOnHMW/KzV5Csc1zdQ2A3yQsIiadcOysdE3Ye
pRkwl0bhdk6Voh8skbR9grlf2u31RO9spmXnt1TiSmTARnRXiPQiZCMK5E6GQvHf
Ak7OKg5uqmpaiidY4T0EwLKftt9Ji8AvNBfjzuQnyRuq7YCLgg7bose+N/U4odlc
mKo1sGpKSZG9Dm7so6cZdAtNOs2sH2lsj3Fn4foIaDRRqNRG50q8iquIVy/kO9pH
RjfNlINkr7kOjlt460k1ZTpWInd/npnTl9Eqx44SKS91umFrr/fnNhvMRn4Wbkej
8cyNJvuFWINkpkV/F0uUQ37ZrLICpAY+MW5GcQgmKA3FbJaW5pueXM+usizzmWMk
NT4gZzzPNKXBA4HIWR7Uj+UOyQC0PSHvvv3WIcbgYIkbjKtm05GmxYvApFt2s/WV
nh+Q7fAoEJPbcwzHAOrJxCWjHQ/zclQGvXTpVgJcP7xmhiDSwNna7n+w0CsyLI9e
Bt75bO42DTt9zrlwek/hqisNExuAvZuuholLRN3uxA+7qmnbsq5+4hPn24nYogtP
cYdlCyZrkwxw/lDDYkYrjkB3uJFijDx2zhouA7gfi3dpVCm3CcWUH9x96WEYtQti
KCpwza5PHEpX2/d1qjfTSCdUS7x5iiEYk39d6gz28XZhgXOCCuutz4lWqzY1HhEJ
Yif3X7bxqgFsWOd6f3AKJQ7vadeIxHNLMMqoz0IDNzCyUPMsn0Lh4OHys8PUu7mw
KR1ZwsvZRbRk0gZok0+Si32RzlLzCX/umRnda4Leg+dGCXHETE/2LwNQ2osVFdz8
XffMcDT3CZ/qPIhGtfVSfczBWWaMe2kUQ/MH10hb00Zghr518KL64izb8RhcwE0g
N5P7y8MyuB5K8LMlXiQS1lThimvd7oIXfJPZNTNzdj2tC9/73/Gigoh+RDlmpsO7
JfiiqJ0FItiHpGHbEElUJV9XWYVwoNcnUeY0aq3fxxrIArpOLTLtzufleF6Nz08e
lALekCOss9zFsPfiYSljjyyXkXj68nMBU/JLq4n7Y/g6PKCE7OUiUMZC/JF6qxfk
601Ew3Uv7JDG9GaRd0awvm606L+/i3cGCHDWEzNGAU+lZ+07TUp1ZBDCRBiNGb5p
65lCfkndNWSUgomsKrEHuUAGe4t4B2OAVA97oJvGkB0LV2X+wx7lnZ/atGlbvoLr
jGO9Yo2WkNrfMVp/5gWySJlQZc1ze0F4VAPl31KBWIToB0mqyvPo80WuKpw4pqVV
vrhDEpZm8yMJAU6qTW+e5q2V1U3zdA9QFUxAKJRQTeZI9beWxbaQ2Ma3xuhsvKq3
92gxO6qw12ivPz4YH9OXU+xJ19VSzb23WY0Gtgds/YAIghRbdy8jUS6SMHkwdtaB
fRWb4nV4PKL+xw0Tu9DyBPY+ggEn7nYDqVhWne212OrwTaw9CMAq+JR0qyS1Lwdc
skHQBKl+/BQokTBlVyMgbzyM8gKc0ocbIZS2YuXMt6OsxdZErIslZMLn1g9AHXP4
9ngIqz24mWuI5AHFYqRDrxikiKC+npH9hIW6Z/e/5B8U9MfM5tq7Ld9rQKH4RHKn
rkPE8b0/Sho4ApUxWdJIDE7y5r7ePeBnNANcew9LXcDdSv3IL4XVb5jnx++N22dN
2Vjb8y35uGSgtkXYKVNwJVNfOAUJkvxxrCkv4g8rSkNOtrcXVKmfGHwFuerdGpEA
/oyVMHnZsmrt4BhgrxYLcEGcXOlaqVKJs5ksXtZMD+69kUdK7ilrxZxnpUPyPoAS
mFpi83f6W1C3RB33/CUneus9n3WS2q61RR5eD0wmGr9euajK50zYwbUoXk0Ccxjf
Gz4GMCSWPeN1y8U+A21k6xAs+x5tjveRvFdUFCUwAQEcLmC+aZTdYJDK+6ybiD5y
uVeO22RuTR/c1ygFWQ+WNskvlSio+xzLQ493xNPgmSaSghgJaje/0+O/t5/U6lUF
eq4WHX41xg5m2we9IQQkRjEyoTryxVh8l8AQTVn/ZHPXyBQyZT3v4HqkY86wjiVI
tfJUUX8CNvF4o5fIVSMdPafxP/Y+rreqlSee9IfPGfl+uhPghpFu2v1uEMjn+kXe
qDceTi5wE2NNktgjWckTf9dWhQvaHZuFkqtTDpWqoiWm95JMiO8p1zxY0eDLgLbE
lwZJi4v7V1LdPR/VwNC534EdjbKluUvuk7rTWx7zttO053EUYO3uDz5OWJYvDEVH
8vMDiyce8sP6C+aDGNlbpezbr+57TtHYXtVmwHsBt7yVeRSbarnm65gZIFoI4BYP
JD5NZl/gWLYYEPlz0KhgHyXsRAnNWW13fl5vY4hg+ECoiMLFuhDDhT3/P8FjdNPf
MBN6DPrBCDWXo6jSYa3QnU3OF8M4i41qgnKC+gJYflQPlBfRqpgGqZbRXeCy1+Mn
OiAvIu5haLrtyolB78nH1qtd4XDqqdMGxAFr8M9oHBdaG5daCGYIghqL5W+45ygR
3QoY3XoHBO2HBS9fuuQO4DmyS1qpb9WpJetgWVX5gmPuIF3RcSiW/keYhv3yBlHI
FvYFuLsKqJ48vQBaUVtHHFkNgBCPrqs51ACv4RxgpvV0K9CS7VxT48UOttcHYbiS
0XyX3IjASdXwE0Uj+AzfRHV0MOH6FtQi/55UlMxNXYyYpEcTE1c09W3sXqsfMXi9
A6jV53vepCM3g3pRYCVA83CnNvBgxBvK/dG7L8NN8e3+0rox2W1+Hi64+eC6BPMO
nhgMLU+uapkh/QyNu23662pApc1X0TpNQ3RCzvbIQAsMZHgbZWrFNHajSAy3cKxR
UThmPT8/KkOCvWg2/dwzoMqxMCP9PPWQY/7hGLxdwx6VKj3YcKlOkj+Fmi4ZKGRQ
iyuo874CIDa57wSvm0LniUJuK9IQ9mtuN1xYQr7li1H8WVsFHe+cNJD2UMeOtEIy
3ek8FtKtQYENB1KiCGwFhgAW/299tuv0kZ6dYFirueWWAIAUuTF9TIj8RFv3PCX0
Y9Vm2aLcE2OPcazNaDyXT8IktIEkLPO3foGRvjN3fpbTTIsD3OZDGYAnLt7R+Wa3
lI8UbUlo/LOiuhXjIJnPf9zm4aBsUVQE2UvrPzxxX9ZkA3kFyWxuGkANAV3aH/ov
C8nJEKdBypGSdiW4eU9PeS1IxeE36XupFK0N0ENvWUnoJV8qJ1cigwWFGaURS8My
IVxeZwR3b0MdfMyJgLt+0qC8gqr0dYg7vgBziac7xJMKTBAhoh0tsglZBFoDXrlv
+szxM1Z1ETVLHVtWhtK6snEijH3ZubqCUHTx2WcB55PzXi/Dqo6NQlXse24jUMQ8
Mx45czK3SqfQatjaLxTxT7fEnzSzGBjFpL8njckUFRLqq/NIjAYLo7nDXyYlh+Fe
ywg2dwq4jWLMOrIkspfcs1cwRZD8TOK0OJigJYKekQO1ZlWjMcJ6Z2kZmyYlpA2K
WrtyI4F7dPB25p/l3TedT5406J0vstVG633l7ENvuJkNiUAIp+vle/Z6NtqJDPB2
CHmaG7AFAJRO12v1WPlVcwgbgHg+SQ3NTo1upcWomBvSCG2SBD4wbjfEU2GN9ts4
iQgVI7UWlbnpDnKSUvqg8wq0NJTFJXHTrGiRtvb8Jt1FziOxXFFfel6vLy/2eLio
V2wD47e2W8pjscphMaYDjtU0Hffj51YgxkPa3Ayan4DHzHZhBbDouMI9VewJ0R5r
OBlPpJw1TmDA6Swqma59Yf4/wXzNApsjwf90X7pO2A5Yo9IOQIyklhKU+A5Qn8GO
xotQU6Jv7WjM96pyP7nV7Y+crpaXifY2EB71jE2wTq9jmoKprmmosCECYdEoXver
nPR81ZxS7vqXoPSw7IS5DZXoOyjXEPXkzHg1hWSKTRsPCYs8NQ25fx/F/79YKW8G
pB4OeeAW1ux8h98jCNao2erViYnGwitK9aUwUz42Gch0LhmYDToMB45lPg7ZTN0B
3+lcNvntEJdA9WCqJ12b7GnaNL5u0aibuEsvGE2wn/tS2K65FCOKU0vFZSzqlvnx
ts6QqunXZWUXIW3KSUozljVW+cadgAd0UQOuNn1KtH7vH3acBiye9h2HnfnbtehV
bgFgpZRmkmOjy4UGrf2Z9ZMYmWo2MzsASYbuzVh3YOMflAelBrDmsJxj9E15ZMo1
xbYBOq9jGE8UkvcokvVKy8jSoo5DhoJzGmaXSw+7foIFPLgsHFGhIz4gr4fnKg0p
6ub2a+303eMV/RLXonVcZhjY+0zhyVF8ronMgpAzPsza4GoP8a5wnPLR2IxF/FcU
bu0cM6OnOTgw4iyuL9UNfHwSwxqdnn2hEN/8qkRgI78oMSxTAZ3hR+PLl73gj9rs
+JjJJiNznI45oatrABFdLbRfxIqpSs/kPX/URNBami0Zkzshmsvqm62ADwqhQYnF
UTmakBZ2n4IQcVXHXE6nU6XnXEhu21p9H1CgBDGVzD/04VhjWbsVQXs9jew3IwiP
oxnAXmp2SwCFg7bL6LZ2QGmT5RcSvblODGGbFEFamHbi9zYAMb/LycNbSdUtvXMs
jj+0PbEUmJ1i7OQ8d97/jDNBLYi+PKa/0pkKQg2OmS3w6RoQUnuXPux55S1WzbKt
cG+LuioKlqf/uCrzWQf94gBpkYzNIBgDmUAmoXcuZargjW9/cSjfa0M+6RXHkExO
l0LIGAQKfsho5CWzoBgIu631DszmFx9GDE42zHh8LSh2AcacfOKW6/C5FmTwy7/9
tGwbYR1wVZELdPHhY0mR+L6FgX3/lIrbBwcSuhAoMhrg8wcYufu7kfU5z2VjoXt+
EYtANPHxZH3wZaGzZN7/0jhsKhCIJ3tff8qX7gdEfefL3NFxzX8BYAu9R3n5S+sN
Gv1f/ERW97063aoFhMhjvjdcgb02iSsuz026rLkqKzRjPfVF7WGgtRE7xbcZzhci
GVMfUG9U7922MQyd+dtmFuasgPlFzppearp/KhH8ydvCI+4AOxz8xGSG+CJ+EhvY
2qAMYJnoaJq6B6eDYIWe3FE87l2Xlv1acYdKccAPFAvfmaHI8826BegSJM5w24z7
U+fhzf5vmMXTA1aLEw8kABrn5C2Cz+yU7xVwYcgYPHqz33/QuBJRUaH/7yGBRkQt
QNLgDt4aiF/cWAtwdDAqcwctlWOtcXng1QeTRQyoyJ5nZIOXp+8Keho3VZs/lm3v
4fzhPF7P3oMpQhGjMIoYPz6OjvTZoeBBa5tsoxzEo3tURiuCUuXwOoKpOVepWV2b
D1qUDdVpOZVsrjeB/PDcs2vBO8nVZ4pgMJDwcOKm2PGsmbrByQNp+vIk88fLJp9c
tezK5PV2HChuu92l18Y0exzZvFncLJPgovCcsjh9ZAql/29KmgaXthIKzrXWbDwL
SEB2Q3/724kAoKwxXixzLm+qS0YHV4ugObuSfI2KvjZqLQdBx8+0DrN+EP99ugoL
voj04Dh1Ns68saNsN7fUcz0GLsRLEL98j+TgPggCgqkkK1hDQKN0YYEfcP0jkclv
Tyhw0QpL6G8sVw3ONkftLRLqaviMXiPlTlWjJH8oWpzReJfc0u3VmL9gELsb9lpt
V0ZnnmEdsSLeieIckdcmKhPJhcCctLbtacZcnuqHLwOkZ7hG8o0yBiZ6GLoFShie
a7GN88drTQvJdP0Yhzj4k/M1XHVfJK8RruhN+V/Mz5yP3Aujjfoz+X4GDjIsiiG2
hsS59woyk45oOPmY6kqMMsRXkrrxtTe2Ud7Fnp3u7nAClD7zmixxYiQGshMEJBFF
cYyrYTErW5QjZ8rcHRDdPsct16cIMRxl0j/lVsku91kupT6/gDrzezLcwYOd0+W6
sq1o+FAvEsxODYiqmXT/o1yJcBfZfai5GaBzI/j1rBLbbMnk3dQpyQqIq1MH/aSm
rkv0S2xTDyp8zMLHXa2yo69SY28lrf2E+cyumnZcmk0ERb4QrEISRmrvz+RXprLG
ID53yRRE7wvyGq/vg5Z7slUtdI+MI9EW2HmsJq6DdwLA64Of7TsRn+g1+/DFB6wS
KxVFq4PmagTFVal4PVvbjFf7F8WsLFYggLq5lXOhl886Ung66LGJPyZjwelhYvJh
yf/5E0vYtFx7PD65+nJC3yuV+l5OdGGMgbtIu3jZ/YEyTgm2xvoJHb+0p+CVeQOX
L10Z3wUzrbuyF+bHEHEMMcRLtzpvryhnw12upt1ERZHDlouK/9p5lOF+UguzlqlR
Pz1v0UWs4bLsY0UH/oOQZwvusnlN/XEMkI/CVBlL9gcwS9va7G0JYIxmARu8VwFm
RX8ico3SjbK9dxjJ+7u5VHQxUKa8HrgSTOUFLVzhKmT64FTvjtey2FCWGkbavQ17
BhMQSZPa+crYneX9QzlDeD9koDCufUM66X6lNkyvZQ3G3XxBN+HYNS65bgIhAQQu
GEQJOvgjGQbbpb4reOmnXdZoNkM2MyLhq7Jwc3RUYWaRW1HkMibL7/r76k9VpaaO
gg0nf5GeG0BESDs4KlrBzrKnBGEyJvRmf/gY8PYr9+V4hhqxtp68k2XvcHo5qbQD
qRM0s/KY7Im2mBO47+qItv8JhyAap4FVYQcNRaWDbHMbZfMlGykjGQpQfDODLW+m
a9J5TMOIp7oNbs2nWWk0Pba5q1mdqIohj29XKCUg1huglprVnqChJCI4AGibT0l8
Ar+fVTMtNT42rSCcvahI58cDeXWkrAYbVRhyRYGeUYopARVB8rMVnvFYgNf/Z7gg
opAciRodxmoJXfiB/WNCGZTYZFSHuFfmYePaO3mqwLv0qczwoLykBavab5En9wSp
aCUS0w2XWOvX9Ep2Hq4jLHpUD6/gQN0T/gdPAzErZl9tv7pbWTKJ+D3AJSs+xEfh
0o/mmLR2OVYH/52eVlU+aOck4LjIb0204oUVI/W8DBgkHn9Bm2MQi1mpdO7X0mWW
fzHYjAPUP89CzcdywKO45mqwNSMAycW0p6T+GlNxSJNPQMPRuNdcFbZfODB+XUvb
y6137EJWVXK4+MxJK33lGG1qoC4ooRqWegftfoTpI3HDa4LGeItEfssbwvP4wWy5
ALPeDrvL3YdCtpEjIopcnItYTcecvSWjm4/oma3WPPnO4jKahx0QaZU1BMR2yRPD
rgiBTaVVzmQUUSBoU+HANEFrvsGM45ggeSwQiywrYBXFvjicePNys0p3djtEAIcA
au0x31eBHHLJw2wTwTXndw4trgQiZy/cPij8fyB+yUicZ03uv6S4w2g0WCAgCkxW
0As0GvOnFFjGGIub8i06zIjCuuF6fcqhSKR3xDhA0pGuN4JDC+kSAFIblQpni3/F
g9JDx9MT+MWw6/cL8Z0KO3Jxr6UkeBwXXLXEnd9jhIcgX0tzPZ7VDrAhXtVqgVqn
WmfsUUkg1REpG87M+uH3yCMtaY/1nfMBiV2jdrDh6CcnM8XNEN1bY0LED6j/kxO1
7A6fPntcC8mgK/JyPzzyJGntHvznOxxC/yi6fdO2RCW1k49c7+L6RkkFKjF8imoF
UfveMMnLyHigJuTljq90txu9mcJF7Xc/HhSP5ZBpWaR/sUYRw8op7HKen42thJ2N
hkF2NqlwzLry8h1CldNOSQPGd1TZ2+c4qlr80pflvMgkPPPUELgHtpBJbVOJswxb
tQxm6VDnAyb2a4eGhPMPBgbWSuJZ6U5PmPssYSVfDt+jObj32VEFcwQ54LdI+LrG
ZDU+L3NQd7xnYQPFnG2aB1RhBIKYM2gRqckF/Ce8xP873oKJ+SmcCcu8poUDNIdy
ejV43QVbMEIVorqVpTcMffuV2pdvCsFlJK93V6kWX7E3QZGDnBT43uvPKOKecN7O
Re0YOegva45/WYqTzqrRZoJaLwcBKatfLZq1r7tUZBczI34WVsJ6N4cfO5k8+WQC
Mr5uEEpuu7o0zwSN1RCOc1RaiBPirWVUu6RSbZi/AMXeSftA/rBGkrO8EwDf9de1
27PFo4Q13MdF7jxfHH6IFg/hnd5x/lyokX2R0ml4wugIJmJn8PLqz+ojZgkDTs8I
IGRbJB2LBOes07VU1JCO7yvCcy0GfzBhuN9l8KEwle5ZQMu/LUpyl//eZ4ZeAi4a
sqItPrxNUYZliKnADUUH9GvCHA1MlDFNtYozn4IZ6bG7e6gui2C+DUF5eiL8ZXmY
tN3J9l3+l6Yxcd87ZcdVQGb+A669Rod/Il/MvdpkI9QgWSdjaqjU5MRZl7nplGfD
7y4rXoFPh3gi/ROktECKyMTPz07TEAohAVnAHbgtDDm0VGsdJGUdCp2EsGmWJ6bn
QzPsi9wlGnJ/N9fNgmtHHS+ggsnXyaBdDFFrqfxhARgPqflg6E5bzn8Bjm8Vm48s
ga4/fM5pfEZ4Z8vADh2bI5suso+EqVwZJKxUrN1McLHbd1r/I57+/4CsDq36PjhY
q1vytegghAy178lU2rkv55VzoxQQ4EJ/silOU5nsvPlKJ0atyXk1t5qi1c79yBJe
/VumfUuGiXdBL6QO1cMvTaW3wBGPmk/GgCPbjEodFbnr2d2PjbkqSZttN8cwRU1D
MHrOqD30sBnOhbzx+Ya1pY8u5mXgjkYdaSPSRg2DpcXrxeHO8azKud4yh6BvPmeb
aWvYBb+iUwhQDl194+aYCw5KtGaPlRifrQBZ/b2UB5G2LtTgBHx/TQkcluu2JP8v
Oa6HO3/bjA8TMgrOpo6V+YY+5f68q9Oq7liss4aOODJSGdy9hV3nKapzEiGqkuk8
kA3N5t79gGcO8EnOLeYgWOHHsNp1LBjigM8T6cltm/PHvEy//ApYzXGdMMGCbgNi
rbGRi5CDJaETmBm9/BrG9Sc19YFF2Fm+UhAFJXYiESHlZVgxD1tum4VKltWWt6n2
zz45GFhBcvt+zuu2kTrVahjqIIFJLVT8k5I7HcHfNFgYDbctSFyeFeMGsbwmQwF1
MKq6L5M7dmS1TXuQWg+0OTYV+kFIJnhSUM054n9os78zqHdfxyxUSTTYqpLcVUZB
/0KvfIVsbZSqB8UrEMW+hMM30Oyv//kHZ6zHIKrczLQeWK1pFIoLyjAJ4pbTukIB
LxL4JQva+/DurWi0JPhuqpyuqYhxpYQrrtwgq4ZrK/frUF2ueAtvhvnnvk7iRd7J
1X3ZQX9P01F/M3lDjhH7u8eobzoswwOOLKpo+FSd7KPfSJyatrLMawVgdTq5BdNt
QorxrSX90tQCDa8LmysxisGp+3AU3n7Era2yBybTyoI4ykd7UvzETDQTUVEPEUwW
LinBAP3xi87LIVd5Gpx8nVdoAmQH9v6TcY2RxIQFh+drlKu3TzAodJZ72nhLIAGM
Lt3wM7E/MJXheD1gGsbQZ4UMtJxZSVVDe1sZTeEDsq6z4mur/5a3PkT/ZEisRA/P
KgboGFgpZeZEvbN8DUQn51WY7cf7sEKxtW5ZRChfo1cepFmjmL4fuhgg/QNMIFe0
bNi7pI56X+WFLYMJKPbsHejwl57AOa528YHPBaVLo/BBpxkgsP+Aw08VQE6XtvPV
Za1KbOYcQ1EDp85t0/T83b3I3a5BbBXzMBaDrgemzFZyQipMCTUFIAD5ZsY9Vf/1
W6xkeRDLPELe9m6dr142iuXiv5aAYF/DvTiDnscu/AIk3kcbPj4ZCAzX2nXL/2bS
SOK78ZnvtExYWlJe/U1D7pW78T3NJ3wmK4ADqA/6ZRRGJD98AcIt4mtCUgk27Peu
Cue+yaMli/CAZxBv2mYMekKz5NO36arCQ9Yk/OqBikuwmuZPkp0NRUyEBSBdRE5d
v+RicMEbEycS73kmvrZlVYSwuFcyYQrrw5eErZ6RNkwFfADtErMFL+w/za9QxESP
3dhUwxB7eYB6/9HguRouTR7qvZVbJ4nYyDDD8cG6F5vHHapAoSVlvZFgLtm0EN6E
DuHWlq6hZvJUp6zg6Wgoo3ZCxlRMP7EoVYIp5svFMjrAtHivnDoCSY5otOuFWJGi
BiziiwAoM5IxSKKeYEUATFTEGdk+OFsrQbbxT3Qj2A1m72feYHjXgcUKhBAAEMSQ
u4efyByBuZgeDdU5GZTG1HEHe9lHPfiNSiT+W6yv8HWsx+fFDvGrBfNEamd3p6l0
SSAPig7MDwRhe4Ib+92ZuOZw8SWF8u+4+pOoUSxepWxlkqTLvVX2ZxE46VTDwffZ
cFSl+JDlUX/zBG/Q+ZF8ftHGuAeiC6Rq6F52fG4RAZBDePenE+39mLEnsQEJHVX1
U5exdPF4K0f7o6VA9Zu9VqwbaUM7U6B/sEnz0h3ImCNM47eGdhuAgZ2e8AMJ8PVi
QCMiTavJiVkN6Mp/bLRCR9RvqmprwkrbiQifL6Z4JSZxqGHMvqWGGhkIEkl9HIyz
qRii/+A9yxYcix2hrGbV+vJR/272GSpm8H2k345ntCm3crhEgG4Wlv0hPreqxoDu
n8hFUcys4TQ3+66W0O5YKEA4JwfVtbUNoQEJDxZNedx8kltQuN9a0X1CJ78e6lOb
nEMtpUdIPD9NDwm1gwFWph7DHRDMH5aMeLn3SZo8cqqaVTaX+dv1WoD+bumZPkU8
kvvt/LGow/5ifQAiOaENQbuTnClV4GTQCCFTCRGGGrYqFnZq64UgxkJYeBjsSv3c
Iasi3OAsKXU+DgXTtM+vFHqT4PXQTrHXNmEfkE8oKF+YdIv9vDKPkEVJrLMzqpWP
vJ1JrwRuB82x7aDO4CBpjlUDd3DKAlIQJ1Mu3cCRKSeGc+Wymy6H76LKWB6KJo0X
Ofw/HLd8M5bbKnDcS3yUCSzMpbX2z1NCYeEEQY/dOjo5ODG0ZXKomxwEyPt43i7Q
sOIlkkUUd+55FOgdnri5Kf2Nvk6Y6Orp0grJUn8RwzEFs2obnZp7oKDjGWqIHi6G
roV3nXqGOyTBRxeQcIPqjd67DudafprbTweuTc0bTmQ0Ca8xgB4Tw5uikOeF6T/S
fRPGh12WJZAzxp5HTIaiDuvlsJFJfdjt8KG5vXbbKc5UmVmlZDrz8s3ZlWQE2h32
HfhYS8LSChb5cLnD1CA5+4MLGQH2k0ePqdmsojoD52EswcWwDTcJcu0pHLLzc6nE
x3eqDPRmytt9el5Oc54KGS9EvehiidrNk/C3byONSCxMNBU8x6Zk6SpgIff4cjYQ
jzN8TGUAjk4ce9JQQMGsFYtPyZWLXP7HgO2oX0r3fBIVj47K/ngaMBA6uNgaFNwJ
8LLYB67Va685vL6ainDURUm23BSi1Qi2Wfan7zvDU54fq9FNvhVqRSjJD0SM0R6N
lbljstSVQnaZwBZEc56pACjM56Ux5bJrlustKwqguCCIyTIhBCby5hsx8PM6yxyY
x4Vkn29JhaXhidw6c2VclbkLXlzmxE6vEj8HFLZNYAobH4i4V9ESZdBiFw4Y3qVf
KRsgXAcuqRrGVIEyT2XzEIKjHDNcQzeP/UBtA49z0eBJ1es87gye1/micLnN77Lw
e+aB7YKENtZBaeklRSSX101GrmWnB1ZLet5/H7e3DyTLgdUuPcOLrWoCwzARTYgO
+0KB9jtJfgWBKJevKJ1nckHpc8ZNgLXYc2/vpuhRRle6jrew3Xt8b9wZzPkvFDwH
oUarNpW0ggn+a4wKOU0Z0pqhMw1S9Dcu7kJgF7PhFDLm+K5DiL/k6rC0Fj2ke7Zi
OfaQ9yvoo2bMC/5ztG8Dh6ENbjCKVSsrcBDQHTWIqK1UgiYpX1mENfp/rotzIkED
R4VP03yE8HnU78gJdI8FeZTBA2RdqklYz5yLhXhNTlxH8EJsP7pxUpv5VCcO7ZVZ
6/K+jz/HdoYrl/P/iz3BzcDy4HZSiK2FHtbeS1DO3sJ6CT1kfCE8hQ8T3l6NwohB
aTRJGY0nD8dhUlIDvmeAa+yzW7seXse28OZbepdDz9Cb3ZxOJMe94tsmCDMGwcGJ
kBKsLrzR4wPpvMx/6lopQ4Qb8zejlVYJ+fkYF7lIli0Kerm/104ohluJxygKfQgc
4+LThoTiKENxrsbmDT/XmHRuG7HFqlgDwxOIdF14wwN9wm57I9aLKC382PHaPRhB
AJ/wjb9Z+r57wMDLNA1FfNPS0MSTE4WlWtcnAcTBMm8/LiBhsDvwqGaNB3mTLsFE
WDz7hwk+qMJCV9cRH+DVfl5F32HrmCjK96q1BZUVQ+lL60tHbfCch6fM1L+VdmRj
KM34l3ScbvCPwdsvMsXbcAcRHu/vP3j8Alp7zZGxdfHuzqZWFDK7HeSwC1BygO4k
8vw+8DSCAm7ZK2Ly0j8ZGdDcA/s9rShXfedwMgkgF3ETOqfFFtaqrz3GyLSU34x4
PMYSI8Fpl5iKgGj5nzzPgUgITMf42qCVyuwd6L1+ZwXd/Tck8Yf2j9b+8b2xG2O6
OXhrAH80KA0BrWSU9RNvHW8slYlIMDI1f0zf0GL7awqhM2dsYZoLTXHUjwITgLqI
qbyIdcNiJolK02Y2wPHlPn5FS4ceXXvlbribk2bibMY4sHKO2TWEqLUeiTNEqJtF
RQ+uSWuAkUsMbiCJu4/4L2m7FXrNlVvnEWH4iut9uKxTiVLjyLp7t6oSDMB+sxDx
g279PpPSiS5doJQI9zfoFzauacP6QmVrBRdLv22EoK00uIRZgcbzY8c0QpGWwmZN
k9BTQ7NbpdfYUEOFwzdBfZbZWF5rin3RH3HfkNkGpxmts7AUG9dQTkRgU9Rbxka2
7J/eGZ7k0D/KDY0rKxBhgg1gVrembLIB3DrPwn8M6bGmhK5k7M22rCXaGjGpirrU
1mRA5njGbuAAeRxoccaXJ8078PsF+RNx5Gq96HbyyaPQB5ucf/7KnyAc4L8XTPB0
ARFQZejnrVuFpODVG4qPpadaHwDYGjjTmcHiVfgMoDIA4AUXpSZFqSGA228A2K2x
VXTjA4lsyQEmkP06tG9SnJjM0YNnnJcvaFWvQZlWFmfnd0hyQW372MlVqImi4xGl
yFLh4bWga+KsFHO/eu/iDoBmc9142aGKXNVd/eEfgDeSdgxv/SjYoAwrIOF+Ywan
R4r9TS0syIDU/5QWuC2xi5EAJ04HUUbsES5jNgnOvvMBaLdxzLw0mhCUEmyHex5G
cWmhWZdD9VqmR9obr9LeW/wm0jxS8nJt6UmUjLosfArg1/8BLiDx94hZlHAShsmc
gVPIv4+2diwmY977VT8Dzbljw5PIMz7JREhhjpXhMXHOxNlxdejQ8PsXBijUVEJh
ived1huqkjUwhooDJ4imWiFWLqz5Cz/1rtZb9iS6qme1HzG5yhcMireDYsrBweff
w+DZcehH5Bk+YVQm4wfZ4+Gj/zEfkDqF1PXQIwI842K1cwNoxe/pXs/kvqAHM0pX
emXvQc0tMjKAmlQ/J8fVOO01VWKU5yH3aewO/PiXwWMq7yO6jqxnkYl0lgBCZH8h
qQgwo5yg9PRB1nr6tp8scfe9GifnzyNUM7U+fJG/WEVwDx4d6H1pi1aJjcK00vGn
ldzpvBu0+8ifzqgFK8AneF4dVg8Oivzsf6QokgLgEX+zruRI7mCwHX+BWNVZkhTT
JqOUFjnbFlrZ305r066LVAJLIiISb6q2FzA8CerNdFuzvekFxWpIPWwpaCtRafuR
wNwfiDsuAXAIz2pu0BuxCry0PK5COvWj/gmqz0P+QO/qnnu7RkxeoD3X2FL6s//A
BFzb6lBei2EpzeoWPAOoqiJhBophAsCNiRNZ//2ss6W27gH2CgTPgHnaj+wdHUka
Q7P5t/R9wX5ww/uqT5UxgLDy1vrDfPq3oaD2dvL/fNBCzSmxShfauKtfG+DFDhgW
hzZM7RZS1sWMFwBP1OUU96NwrTZTWSOtLJruwHy1pYgFnFSAi5CfBgT4vWui9Cki
6/Fuj49Pah4IIMK2cy6TJ2S6plGQ8W9KiaREgjltQSuEvrDyq9AOxF4cSjpILtNx
59rEfPpTUgKN+7YZKtYHVuQiPql0decHEWhuOaJ9hVRz+SyLs0j837WGwLJ5x/MN
ymcwzJeTWf+4kgmSTBnlYlVhOnAKc9TnwD/KkkqGAk27x5XXm/VTUW/LC6rHSuMi
MCajOVyriQSNKWA7vJ0EFyhhAUZVAq7Ne/OQtW4VNSGFCg3Y0B6JRfvmgKbQ23M+
TdRphPZfKSbhsCdg/dXYcGtHZdLBker8TbmyYf+e+zoZ+JOyiCK1jb77H9YdqDUL
5bXwKFRXUCZveV57aFS3BVpv30VBA3EEl1iWyW0/kIWn2SQTVEYGOgZl67Pb4LX5
NYCfGcgcughX5C2F3gqT7SnAB18a+DXf1clcDAKZIvzRgVjzxJthBnCghfVMjA6c
iSQf3anACofNOo/XyuAxZGwEItK/EdRgvvVIOAuldaxGdc0v97CK9L2srq29LD2H
F159/JwIDmcxqI/Kc2/mL8Fu389dCxGeHCkVKeIYw6VQQkAn3Q905Uljj49DHP3B
eT5QFmeGdglTOnCX9tZSFiGbDMCn/x2oa7X84ujDP6+48jyFkdb6zigu1gvK5Nd7
f7JQS3uPNilYevAg2Ygm9sGCnhUxt5dxwmnU3ZTNvW7hmZ7pJHZ4U/SUp/mgNRV0
1TOSUIWYsIlbNsyqao9/bJamCZFIGtqfxLYnv676TaFbLFRmGshrI/zCBcuJN5gO
jHfLC4KrTmTF2SDOzwB3Hrt1SJp+yw8SeXaNUj997rkbkxiPuVUgCEa3LyT/hU0S
c4FbEWzhQ02WRGWiq89iD6HN3XqKxQMRZ1KWRA3zNtyiVJQV9qAu5S/Wy6BwGYiV
XNea/lnutTQ7Fuw+P5iVTHE5vgExes3aAlqqPv6+xuFRCNwyYYyib38LW/jNUv/V
c5jX6x2larPx+YzW7fUbWGjFRfMO05TJzN5P3nL2VNm30s/Y6kqDEjIBjzCHKlis
m8PSR3AdECP1iZaG41kUt88kN3SY0FV90/v/OMJfGPM44IPxfoNZvwUBIDafyttk
Yr3r6wd8gYG6kqUHKbHM9EmKUD8lfsc8p3BSS81EPwueD5+4rAEMPSsFaNLkI2gv
14ddjwPNbCpEOt/4yL9GNOmKM4/SXpewBiuV8gF3kEHM2csgdyWrzWXPjn3X3YX/
wBtsmnC5H6Ni1a7hrSqaAyjkWq64hUpS1xGs9Vz7WC+HaFNPtfIm/KbBj7YuSWav
4NTvH3dbQqfpKcQwZPZTRwHzBLrVqkvb0Wrwh7P2ElEd924gGj7UIApUpbgu2QPq
pQrCCYII5HWq5DBfRAY8rNMrqbGZIYltbF/2vMSXvZEY5isiQSdqQDQPhY4h/+Rf
D4b7iqIw7uEuMoo9EMcsPBD7v02KtytOFGiWD8CWNx61x0t3m9dPEO0TggqibpZX
CK+slg0OngAJ65PCe1c1UF/r2+1cNclN9E7LreJZ58A0sIuu0tVkLCPj2UxV7eDm
SXhOHBTHd5oHQv+btI4iFHc88vINwgPH6g2dFyw0TlD6bmyCLkyY5ZSLldL6hsW3
IA1Lrr6Hyx+WgeNWBBHFsHGhy27A9cVFwWEfNYNG/gcma3nBOYiDYCAwzevCndYj
E5qyDE+8Tkwl+RvGFEoE+y+/ehZEzCH8/xUC3hyOiS8u/Q1wCWKuh3NGCkwD2a6/
S4XrweE6yFbrrZDajSg/hZL2Rpzkeu5a+aPeHVNonLQYLOaV5gUrEWMkKmSeFayK
ZWkezeD3jk3JI1Lvl7+E8XPrrAbf8RHvHbbP7X7KEf4ZVLzdOkHfm40nFuLOXHvc
VWBDxyEG3UlD3/apQO+OSmfqds5dITYH4kDysxWLwGHXjjlP9FiNqikB8460C5v+
Fw3DSki4A2eLjK8a/QWgBdN8rfCfgMq6m+tAggTlwyeArp+L0lupQg0FN/JsSprP
nHs52bE8xBSEtjjtld0rxhgaLJuJteqcN5L0VpD0M/eRYZTCPaLiHD6KsvQcRZdb
HHtnFpcOAkULViErecDa1llivpQfchfmmY9bQu2wPT7Iz4JVQeEfCGcyav6tcw0m
pyEPMtlW2kQguQCdPjIy1hsKpCXldy/mPMl0kRkf/M//S8cBjSZqgJIGj1TQnf5y
dgH8xG/eIZnKEt9c9+6pulQ+tc29qC0+DRJJc7lB4Z0PB7bjoKlrMO06q8mxIp24
H0Kwq2kJ4LlSv5/STvkKcoHU/bzGf20EQUEtVeEjRFtUx2ryLX3IJ8WKkqOjThd9
casbEYbm6bWqFaBr+7RrlRUxNMlQN3skU6l3EXS5zHuRyklb2s5Vn9/Tv62DzyfJ
ExMScDR/B0yclCRS/XUerXSvRKsS/mMuYGKKvgCJ4nRM1jPnDolvweeintEGK2HX
vasb27t8WBk2FLwpoOlXfFTCSdA/9+GqQRcDx5JwXdqay4MzGOH9IDTLgKuCietE
abhAp6rxwplckGv4/zxD0ifVNIIKRd5OI2KDgCHz6fzVeLw6CI65mlVOiF/jLJ8g
GmgqH4ms3JPhH3NM+GiRxwGIlpOg5TWg5HniDfeDptuUvy74ejMYa4FHro1WzweY
wvoqYQQoayr0Zw03b8nLRMbAlwqmgGgH1I4x9SzAH9TnAll2TnkXGw9+U6aquZaW
2QxheX7bcWel44h7a8LBNLL2IFTozFQGhaM11LVk7sI4DuVowNn23q0tWrwpBN24
wRzyfjD67Qs0YDC5nvKxeea4/HigSeIJ0MY7AAriOnlU7H8ehi13FUHNyZMB+GRe
Kr8FriIonBkq0xErWRVoDy/xvs0yZOgPON10un6/+no989w858jbcmouzr/ZHO3Y
R8AzPM16uF8yfSd1hpDDnhnrsfBrqEDTYFjZxa7Z5EI7zmauD+id9W7pztVnYIr7
LMNfgaYIHNuciKNKG7eAa1IeeztBTSvWbzS/oqxBV2CHWLl0WIChN8/14YaXpAFJ
lAxEVJ0nyiEmpmNI3b2TGCTqczIhugraeI0kouuAWAsyRZRjhGivhd8Lm/rxDXr2
R1JsoZ4COwUoveRw53VokqGDDCFrbc8wh1+XhzM2hkMmaL3n92BsKkclqd0VaH3h
kW5aaFlttjLuSorr2wAOkrzsl8RWjWCc7QYFpWzMQjCHKUYNQKzrzpDodfFFzKcN
i6WG4R9KhBZNTK3RCzK+8AE6jvpSkvUJGpvlrQmuF2/vImtw8c9Edcs95IuqOgk2
s2gVj80wHxxCuFFuCAhyfgS4xvfeCbVTe0kyk9699kXJKbNdOELxfpiEibBAj8Ty
s5BqMVhTW8ng9NIH9NrvTg/J52Nbz2Z+AQkMlzKlITrZHjrUrSYJJAIkbl026mG/
cyT9yxy/oUpA1t4EAJf+XZ102pn/jOZUjruniV3oa3VFuq0RUsrZCFqqdz+5Lj5c
b7CgQwgvQVjl6myi3fDO7OZFiwIXfloqpvjcrTriJFiXC7bqNCfri89+Wud+GOAi
IcFYAi5dj096LIDf1AMcefLt/WufkmYQQ9op9lhRhgd96IzzvcEgNlCegEvxVJLA
uWJJHQHiS/DwyhbDesK4pj/bnDqpAIluyy6zycbGemmp84fGINTYj6MIPeHUtWAf
BvuJYXJ3PGp7iq1IgKFGwL60oCmQqM4N5YEvOPcDL9SkvNNAACrM8ObKs0UzDAHf
CerPWUsiVGgteycSPgZZaPvgALUF4HxPOfy5pZ6yuwi/ZM6OkSYtixvEFRrezFKS
yvNz8O3+ud+IXCDde8qIuYtY93YHayyPvqAf/BhI8CHwVuCFyjKU3cx/yevpuzVT
fVARM+YJZhHHkrWWArThnum6rsEaVRr12WCvXmPL3XvqQwbmgwi5F1Vt8iGJ+war
+PXw6GnmGpi1Cr1Fly9B+oHU6UrwK8Jmf6FuDvIk/oxUIU+b99wiZObJj7LZBK2z
OVLSJG5Df9nDmJXtRYG0n0Da9uvoUhhIwUd8hX+hlsrK318uu63Cxmk7v645tWt9
/PHWa8XyQcSEHC14Vi8os30yXrpu/XkrSjBWxQFDV/1wl/RbB2x3kxlCjKSe4aPt
0K767UT77oU3CCWMUwAbClo255v7qjdoFoSHyMljttLpdSQxzReImHAPzbB0Gr5S
cof7uHhVzhp9g54dizoXeq/Q0YuXNpKPEZaec4cpzJZvmx6XIMmqlJTz7nX1Op+H
IstxYfHMT398J8Ll2WQZgTp1xGr7IhqPlTuA7tu5eThmc+DM509eZXgBTezNr136
kPJN/mqB454W0sEJgIZgrUPnAmKs8XphPF6lYUENcs4o2AXmSyHRCEyZTRl/b6WE
Hctkpb/86Ixw9S/VfHkNFU/mUFMKieCO+bvwqfMk6J09Z4e1sLdFRgANv2LbC83S
sj8opkh89LNpWqZo2E/gcRBV0m1shgyWLiGZ+iFNRm+7luY181Fwn7uwgJVuyunb
VC18PBeU4L6q/TiHTnVii854vFGXjexKaVrEggcQPAZ5Gs1KlpSzVIRG5O5l2ZV4
RLhEJHjUOiLSvjS4wEdMvY3i13vQSfoh2qNFHAEp+SdWbJCwO+2HGXSaP+Ducl7i
tgqqAUrvvRTRpCHKUWyq2JANgRrqavwlyat2rE6vHv5lIUFeFvbr3vZfAq2mjDZV
x3DSH1dC3ihVFoGrjpo6cHrNHXNgNa2gpmT4YtJTKcbNzstQTMucMclPIygOwoM7
Q/K6WzwVV3IVzdSe16MuTezfTiYoERYbZOe0w1zlZhnH6sCgBPYXbcRDbedrmMKY
Oesq7EBB3DEeNrEJvI3Rtpzdw63orB7LCHz/A0PSXZJUY24RYuQldl4rQXzg+bm2
HqQxT4mN+RK6MVp5RF1yVK9k3aESR9J4qJS3w3wiD1NK8kLa4ZkWxutkitQlChLe
GaVBZSj7d7SV5u7uCXYno5E4zvCk8dUzGy890b+crxkPdCniY71ElqHQ6u2xwhkY
hiV3fSjVfWBLKw/4zlm/KMQ0lvbYX3OCjXPOPNH4rCH3w5RZV4FChF8+Fw+z58zm
pXpAGtGdMxgSUqyTUWPZyb0xWrpvKNTPEbP7J3oLuifaqqu3o2yZ4dnW+b3XuNK3
pDqJCB8kAV+HQAeiIiFTlpPpVEmn9kYcfQqDNYkiYQo5ARR7P7YbU9BPpmXNrKHV
KgMr3MMd8zZW21LIhlwiaCPMXLQ1gAVVk1CQ9w+4M3T8Y8SbxZBVQw8O1XA5mFd1
3zbiuWzIQ1m4+XosO0r687zQxRAz28/bk7AjD9A+PAt7Q1X321ovWH2AjzBKYDW2
+hnOLnMgtR4sp1DZ7qyRJPtFa60P+M1KubqYZKODpTVl2qzBmAEDOuxoOEcioIfx
SL/zydVMDGgOuRUwcE9xdIR4CZXHJGGhluVU/hJEAKJYA1DLqtxYYb9P706aDN/C
YnmGi/M0aFResmJDcF/pVNr1bcKVh8XAF8e6sBsu2lK/LITF6FEdJvYTcbO9LKCY
VgstL4QT26vsQzSYmxTUg8qzovvGZtDCzt1qahQkWBK1gm2AM7UR7AaCzZROi29A
GdxG8yND2FJjNSbysgXir5q3Ctxa/BPFDvFWeCNaufuGwuYzHd8DG2Z7sqhISOCX
1M5Ytpk6k0XUB8cfpzKBjNVRB4InIobfWvU7Dpe01xYD4vrCfb/8TjuBn2qPH2t1
fyp0sNm98eZXZWnI0XWo3CJ5RprLoCiGGeYaxkuVLQ746JBE8zMg7+9BJ0UDYSUX
oWCfH0ntN24y8bU13uJgqVjDO88q5bjewlXO1EiMJTq+NZwlp9mbHQkKGNdJBwmr
eTWLzvvPDYEnDISKWFKiJwY5RsrsPF5xvHJ44RWmU/+r61BUq+LKkjq5Kn0ccUgh
eZ56H2FcPvwyU8y3CTcIWagovXpvEqFzTR5gqtD3cnw2yBCyXe9nJjH0324IC7/v
YJjAHYUsfqCELMGv6XvGyrGPiArGcaFLb6D7BYoabxPLGJPRx27gkNyjvi5OnjgO
UHlzWxaxa8pCY6V6IWTZRM28JGMIag/IiuAWa2JsAc7suS80DiRYbvPIhHMS48iz
GXUKrynDcLP4mwBGBjtunR9hhg9i06Tx3YnWuYjNhhcAVNo4URYk22E2rIR8NbSh
rspzhpwQqqjCCv4751/hcKUib6HSzXWz6oh4FuKN/MqPtb2fFToE1HT83MdmSLPD
PvBx5jHWVJWfJyGneCZ7m6jwLw9OgJyGthNjvvLG72qLuL2J1hL4K6U+w6LmD5HA
gDO8/oxRYft4DxBxmh4ebmA80QvBbW2INnFy4TH3Ja7uU01wCvjAfIDrEpCePKg1
+Z2Y8kc2Y27DFz3MyZXqFxwsIJfFsQQsjcFmzyksI4QWV5WS50r3wl5nARo/pRI7
wTxeFbWzaN5ZOj6juZ3Pw3/01JdwYh6lv9LxKT9eMTo4MptAQVA4KK02y2Kssm95
Sl1CBjLt3vH2I+YA1dJi5yF1zMJcx9yti571tMq8BCsMd8/RCWPrKfWsgdpcukO8
ER4IV2fHaLQBe/eYk9ntscL/zqQ0Or094+SFhRVRcqKRDe4pb7/tls4qg7LM9yeP
P6nzjDz+PU6i/NEzOnA+dozoUOGm6yj/MbLkRYMS60aq3kz1I8Wk61vAzGM9S58G
8fNSj0OgH2AOyr4OyU3MDrCcw+HwN6yaP5YIwt4iGSXbgH8EnBltazSJuV2thVGB
yU1emVMlo367MpYZNohn4MiYTRhfGKnb/FEuojDZWzpLUjyxPqRWt71tBmgobG8j
zhBSNknUsB0P0dOGkFAn5z65ti5ccCbFeOEOBFOR/H6VJhVltsppJHphzFmGpZtS
ff7RX48V+hbeny7WHV3/cskOqMSkCEtzb+QLRVNCUJAlUYSz42EOr86/48IYfrBZ
XTnMNqBboGhQ5WaJDA9l/jooe5qXNwOTqeLK4GjP/c9ve7kSrHBgCM848GwoPkt5
yMMVgHcaTx14T8zw1xYgLUDi1nDFJTRTe2j+bq19Gq0ufA4Dnz7GxD6yBKxugxi4
C3IskdeQYB1PikyB0lU/MGFuIIAvhScueGesjuEJ+n1qs7+LpIqZus4iiJ80tsz1
+uiFp35Pm0i2JRCq4aNkLfnEouv2PElpl4hmAb01yISsYbsBnSh3klGGL4FayM7k
I8C9VFSSn48LRX+UBOKWUuaIqMSHL++4hWoEXoJb8NStTzlMxIkLMY1wzWU5xrNC
IdygAuhW83C1ZmNv+SjF4RnmKQ1rjgQqdw4eL8dkFlzXIdT8A2zLs3YPq8euR6ju
F1pHZIsky6NDxVEcP4SJISpUpYGt5GLyo7PjR+j8alb/l5ARsVVR06ZXRM6ZX9lF
lxZqqGBx7L2EhOacdWohyh+uXbL0tZKCtASG84wFHQM0ow0dW2kTRoTUYcKgaJqR
1WXVO2nG9ADqjeIkgugU8EdoZ+JlUEl1IDWXJkE1FmR1GCg1dx21FxRqv73a+KeU
9w1sRvdbaoOLM1LyN30MlHHVAPsBzXinueX8Dk4BszDhBQPQsV2IoS+/jCtX/lk8
sicILsKBFqO+fa2xPmIMhcS3OYeTexC7HD+Z4fCi9dU01DQDVHDjr4tl+zBptrU2
RFRXCzjgjxD7UzR9Jw/LZgsZyQ3pvleipSZdzMB+VCgeCOURgh/7mLEevFu1V4mv
H23BkR4B3u/rTBc4+ooRIs72YHngMOVwdkMJW4QSNwLQg66Pq87FHZXEc83ZGkl8
O7jFtkyQDatomFnM0B4YGl5fKFls3aOzw2NhOyqLMH73T6kN601vQHsKr0tPxGhG
GIdsbnhqSsuBFBMWpUKRu8ShEvJA1nKF04jGPe+BGf1kFUUUK/f+fqOUhUT6//qa
qF94LfpRHlii1ClFCTIJSwlWEJkJHEpBit23w16ePx/4zkyHCyx4NqdZ27m1vVmr
2fGOLwGQ4mcmEWLONT/4rAkcKDLJ+lPH3JPz5YAxpQ7GCGVqO/pGDiLdIbJZPt4k
lY0e52j7WzP4kw+nHiiLs/fYhR7tJfWzuv5U13mZFj7Kmb62O1lPRE0vPKyLHpba
hsbLSlecH93yeRCra2RerojhKHt2vd2bMNZ0lgr1WJLGuESEv2bCbWrJVc42sYah
WVRE2oTMH19krd3nLF4OyV+bJmtmSl0o2pkZgVnJ1kKLea+dhx3wkGaJk4PzNu4G
pWvuS4Su5zUycEyzv4pgMV5kzcisPzR+MBYDi5GAyKrValOrteRftN7st50o3T+N
XDXGcEpi9mx0cYL+rHwQTifc8YuDKd/bW3lizHvEg0Qvu+ihioEvGqYPG5ADDaQm
SpFoctFK7KefMdy2J7HWq6EQl5MLG/d3qpXYCh8XEDgl+uvagVhK+uFDmXzWhpTJ
ljb65DFu+rOJERxef/gLW2e8x7gz2Y/2CcEFEg7yg+JXhajZZiuCvrtsKKNw8XZ4
vfwJ+4kRHKZ8/cz5uBr3P4cz3E+S6cPTiFKTmKCCg+zIEVgk7i8lUmGt+1lVVRTN
zrPDxMEHKqFaIbMiF/2nJdIDZeT90+Z10SaHcBk9JrcmMcnZTBuk0WOdhwo6MVKP
4Y3kJgG+5odjcqgeVeiKWBGhL3Q/EKKT2aOuR1wuHfezYUStN/jBF/6J2mvyqOCe
Gx/eieLAxp2l7kD4gO0gOB4+ytY+A9I0xLmD1tCicdz/q6bjlOTwud1SLnio+02q
4aPkBcFhH7vcuUV4ujvl+bl9Id3dt/P5w6jJCS0vUx6J2BCDzYTvimgYmZ0x1Og9
+KlfWzFZM/U2+kxTp9zBtOXiPOVo6NeeznU8OW288JGURn21SbG1pEOI9TmRJfB8
HO5TeNdeFbQ+2XaYxvHtgUTYFuS1uxv+vS0IImKA4aXuPWzCn2oUu3zXVdhoNUUB
qJJgAxlXfkshIA8ue8XhWGA/7rK6BSHYUH8jEGD+P05JKRgYRa6meLbVAQyYDX7G
ba7BAlWu2zL9ErIPbaxUiytrzwEQj58xQQUZxJpV+C4iQrIegYp8swcSkb1ZHkhE
eqA0FbmtfNUBR9yQfkk91s1a2ZgB4SfbiJcgCCTCdTjVM51HkYLSdk26rRrgRVLd
pWov00KhPf7DXUBEKGx8MYoigD7g+T+7ycmD2gWqgdS/uJ9VbdXRjOrlHUAMUXGy
CgO72vId+I2abwRt403PhRfOWJs7wXcJPdt4Nhp1dvB4kWJ7F4ALy3YYs1mNeU04
Xls8/V8CZJ43tSsQeYSNU+lhxrNHTAdXnTjU5qjDyVj5Tau/b1bLMrnIDv+GpZ1H
bRUNyqwSRS4jw4MDMRk6YDqVZ3AgjRU/pX53aZQMRBYHJ8020jfJb7AvGcrlkDpT
4JsjAtsUhF7jYEBAKAh23WxDe+j+Jx0toCvKlfIeBNqBJ4yXqVNAcAPNr85zJ31+
8y4YES3/vCyWM2U5UKTIQzhTU4/3J40WyIClDRZ+JTQbG6cfUTZ5qEyQLGVMsGmO
zjsoO68H4qwbfd8tIZZUraE2Rs8owY+0a/TAG2wB8onGbdt3pNrvvO9nxPj1znDX
Ebutfz0yR9Rnmuo5LOYoe/zVYgjzdD04VTG7Tv0iV6l743i2/X2cZalVt8VvnDRp
sG4TN5/saJIh7jKRrGwKItBDER/CDjxExZ2VDmbsOR9Fue974iaYzlOFbCot/zVW
D52ddsZaJwysjujzq6OTTPuCqHMpGRId3Oru3Yh0kCs8YgrWO608gFM4tuaGPMst
NyYaz0qzLiPXWIb30ncU2FWew63cLoX27MoMUGy4AR9VXQ9j1P0y71LoKHR/ugeb
8+MeBUmOL+qevL98aKLaK/YKtYcfzZMHJKkLCH+yuI2GIHQEFyYaMDxygyjraRuy
KFcpLoMxJt5yYuCG5GwjFY9Ba2LDsmy5cWkMx7voPGPGN/nBirbAMooihTDdX2F3
Mb2OzrWW4a5PJ3WbVmuVQKQbbP/3YnWy9w60L+vnavCR7FDK2dnwLcFfOEncuoNg
FwtpVdTV/f9rkW9uTtsufa06Zbn1PulYuWCZCTT6nLvpz4M6TOnAMLDKhrFzAEde
m8WD6bhqiVQYmrMHWhwnposEcloROV09qv8qAAkK+2OkmL5txTo8CUfImaJ/uUNq
NobDnPk3CkcZJ5BNq6Kt3+rqHsFzAhKNVrapyd/pzFeJ2/LIg3kDp9/4UmQhkg7t
J04Oc/rUDwe36+kzCrzmQAzWgDLepZor2C+s7gvUXXFmZpyuTSv2ragpIgwfVkHS
SOztSJbuSUVOC5jvrdU/sELThYfTEffB2fcTQy9vlD61q7/TcLMEeOEAfmqi2m+7
TckkyWEPH8duXeCcwtwMYIJiz8p3YCX9xwClpLNB8SdWRv7OLyoaBN94u4boOlBE
Q/8FRWGcTRGWH27IZ5PiJ0M84mFkuZyosjIHfg1tZb1rYr54H09l4yPEmEHxA8m/
1T87dZRPBc5WBVbykmEnvuJudOe2yp0UQE+SKf6xPLkyNNl0AhOmLbvymyiSUrIN
oMHVSgfTY7SVOBzhGmQz/XxhtZsqkesQtAMnKFAgg0gRSbNesK7gr/KaWwcseuUG
EGZtmYk76bCodWCE7qim2/Qtp8TkT22NLMMtaPdneipTPOlfItmLw8erEoLI9Fw5
mnMmWq4XndSokG8Sbl1pXWLebfJmvmMoZiVp8eT5IV3J23Ytm+KZUin29H/j+zlB
zrreGjmh/llZvGbVnXmW9G/P94l4sbj2qOv6VMPRpxKch3OaXM8VO994o/vI/eET
a/S0RKKrTrV5RX/vz574Gihxi/91lvrE1WO4F+ES6QUwRJ/iG0UJNhX2bW7jue7q
PCx90PiNe9Cg0K+rGWxZPibCbdln9l6e359TvaidJ8/RD+GunQywmfNn3KJzIfdJ
RCue7Z5E5nYI52nBobcepH9Pr4SL0L+vQdQ+E3A18F5JlbRRARWIGCsKJFmjgsjO
49Fp/Zht4Ra5tp1mVDPHM9f+sJuoU9bli4OCoG5bXQyvwF1aaeZqa/DIq0AXifxV
OK+CqDlRU87t+gW67AabQw8QXWHmMXrfp+/6l77kMpRtCIbutgYQ/Zjkfcfqnzwx
pIcHUnEgfbV+DtxrVIB83uxuC3nafQCF5KsdjAmj/dCBszIGNlzOTrK8TvRQTPSU
ZIWyj4bde/fnA5zClWC/i3lGu8DpQaieSb001Sk4pJ0o6MCIuN60frVxFWaYaS+C
kn7kRheDldbmfHx20hA45xwU2S0o9DYG1KtDZL99+JHkVw4ovZ/AWbV3SVH5fgpY
RNDX2yWIhrw2aCmlbwvLZG+BSt4u+93vS+BuMz2HErqbjBXaORE9zc4ZoRhKRDQ1
exfO/bNdQUXsSEM0Q6Bo58+COGeiLhrscaJlv3PglNhQJPuvnNi1/K/eVlbpBctC
xBOCglhyLhXwHqu+LcPpXNa4cnBw+a+zS5NJJ9dLAF4W6I7VCOZviKhqBaIefjws
yn+vBOhlJPoLwVn18wgNRmOcq3I2uGPXooYfQkf+pQzcbSHKJOE7rzKwrKn3zbp5
XPWwGrKX2rE3jN+nGPu/qsfJo11aKXMZXNoge2dDbFCdQ8XvunCAb0LDBxQbITL9
OFje+pWzoaVBPo/hyguJJEXf5A+gETy4/fxYhFow8IXZ+xc1AcLUzWeAiYZuLRYR
5JM+w+vrWCWk36rsVzv3xWzBQfpW0IucNw5GSiaB4NsySknMoX8gB41LqEUsGpsm
ouzDZ3wYMoVkU+Yl5U/ibMsSkpJb784TvIRPoSVbZxfes+cgQPckuyV9kk0Jf7+G
O5TFphQPto0mc7iWVXloMvPwut97gWaa9LA+UH7SJwqm78kj9y0m5Bn/06vzh7TE
I+yZnBG6D9hfUVgQshF0I3pWeA71hfMywAVXSQ1Xy9pZtlEROSPQGw0iVAmt5afi
fqsbYwy7Xqp2jQvEeeu5cVxdvLZsBxOieAU3R7uLcYWoXoWhtlpysgxb7D+I4A7q
drDKwEF9EY1zR05evzUaZ39AHUV4V5rfUREl/n+FZcwF6Ctu5zV8h3kELs9yInXr
Qb+pmuw2+ZI8ze2L42ADKnC5BY+zLh0XcHe/Rc2o5y0/+l13QE+XvkP0cGe3ny9v
JIA7RSqaSCiLgWN7gLCilt13w5DJLsFR/tAEl1ME8GVHB6tJj5QM+vQLvlO7vNq9
NSGy7fb5c5m++cSGOA0B+IaeAEYJ8uYgHp7MeJsq20oU+kYDtovT/AwFh+gFGF9y
64uzqHI/ILTK0Cz7+A0rg/GgeKcDcWTwznoAH3uU5+0MvB/mb8Hk+dhqhMNBRs2o
BafwT4jna6+jotJig7xr0e6R8TxHwp971OjuHyelsic968+XNDsz4P54DNs5HT0i
xAiJ3Lgl7mgpElt00Mmyyvut/ojYkp+ysWJ16zeNSlEOWk7IE0n6Vzw5rfR5RYXK
ThMbUE/fml7vBPpELdnKNlsEJxEnHi5oasrK1UMkw/8EUPiYUd9iz6ZhgvJ19yqX
q+A7sgHB6pdFGCA6bZCCJLdP6ogxa/K1752e9LFmlkYqmdSWXnY/vVtHOMgX0Lbc
htFnlsk4P89bVq64JPRUUtZqPWZWk4WBCKaZE5Y6Sh8sCfidpiAKgKduOrZeSkuq
hBMb7YyGi93XEAJGOigErMTePB0tmbA5j9w6RBQUUZVEpuL5b4WPoPF3gjpARLBy
MDIMbVz/o+akcC6b5HZQVVIhWU3IbIjKE7Vx+JnPSFpK0WpbowT6qeHvzVx+GXo5
VROgblBp36sfQBv5Ksrt6uVRLt4C5JECxef10Ky9u26H7qRfO57C1UoKbFWsHVzA
uakCB7D2OnbbbHRdXQ+niMFnwt8lBygeYfTI9lCumEJXXoT8aQm/VVhHINzSWVe5
blLj/bcTByKFfoNa/T3V/+qFfrCcDGdoZM5hJMb3kZXhSOpbz1F/1pQH3FbAIBbW
mUuZdOwW5siS5evDSeU9gfTX+8Y0yQH6/76C3YLnDv2lnm1FGXKe0+tcnU+N2vZj
/sO1C5PiPTQKh3ITCZ4hLDgt+X6hTZkVgk7yCwO7h6h8y0l88joD0IAb5IPZVENt
vcuLgX7IN8ByioWcfz4PRnIC+jlPtFr1C+KdwIvX+dTdRiO/fulq2zLkh9qhCxls
9SMUjXMnXPuuVu1IzPZBKMOSyfpkS7piwXUJn8B9mcMRs3mhK4I8jOZX9I4I9F/u
V3ZWTsl+fpNs6iZ9fUUN6o9iV2vrBBVXwNBOpkQ1JL62WONKlabklRgurPo6yVw/
LCvt/1z4QRljd49ChqcwjWA73WiPu0bcBBzaM1Ew13pfJfVpfxjiVxl3H7PWv+kN
oB7094LDcgZ0m8//skDMJ0jFzh+PdqEAbVvyezmmQxhfSfAQOc26jrMBfoIHMNHM
jBbi6R99YjH+486u0r+eaIgrPZ0alEixJPTdJQgjhEaIUdnA2L0l522Mz2wjh3V/
k+DhcN1nYHqgHfX+l+xqwrYmNTymfwG9woMyAVig88eJg2XvNl6T6xfCgIOea2Wg
XCnj4eUXm4qgkXh+xtuhZmQ4g9gB1sQnjUYf8eOseRqpXhBWPrLpinsgTySzlE5G
QuffcCy/crFQGbBOEr3Smia7VRyupTysC5w5xc7QNpcIHyJ8c9rcxBZbaBMxrGd3
s03d8r/6gNJjhMJEOgOIgBF2MxDD9/rcQkSjeOgcpPPAMcU4Od+WgnD1BmlpUddD
u60NU4lv9f7I+nOS64OEe0HPOaeyQ38vq7pBJV2xaJ8mgIV8znbi1KGSW3NzWytp
F43lNcxp6zRy1EjOVp7ZB+PNO3aEvLTQQ30fCoRpKm3cQO8bFDLvTIQbMXegAhyA
yNF1v9pCtmK1vjZLc8CuM7KH24EPoR/ZYj9ndBWUnmr1BpqH+3shvV9+kSQjWEea
5X7LC2yqAzbIvbBtXxSURe1NcXDjNiTRq1x0XIzOfnVqPCkWm7zsrRfQhjeu1Mab
+As53szB+RCAvKlYDDbyu67p++azOXEN6G/uViwwoeZT9ifll7avvfFrfh/Y4lh2
r5AvzHE33KhAi5LecIi02lxX92E+yAEW3q2DcvR884bdMAa5Wv5RaunjUtwE9/og
luRPFudtgyro7fFSZ9YeaIffxUitVGdEY/S5J7hP0fscz0CfDF/hyEKVO6m5CJMz
OG/dHlhzUNIxc4MVDexwkkgm5xg36EwAf7U8kYewImm2rCppAUn+XBMLZaP/nVou
hnMjvT9Q1saPAHdq4rVbNYe/mSvOPWGP7VWkw5OXCfmhARC0pkGxxZ8pd2J/QoWp
9N1l/kt1AkpRThKZ48sXX8hvIDqict1BMTiNxx6jUmtgUtVXxawlfuzNI4Zk7ssR
CabUqrSrRuftB5lVu2o5+4ukJPF2sXa0+31GuRgtDPvzMsBzie9nNZgYEA+dkder
tenPIAsXnnA/be+r5hoaO6mIwSDeIyMI4cZX/nae8Ri9eXh3I/KETTG45mX9ao6K
JNbn1WBnWq4nKsaDgW1CyjtXwL5LT+ZjXeNcZ+depWbDkzdA2xbsO9e9jUCs7tui
Xj/RURnUYjo2dPjIEUcoMplSXelyfOmzhwyMUEAkOevB4sDbGNeyA9M3TIHmQrKU
h5EcXWQwnfceSDg/z5lvawvuaYaSE2npoKG9hNBptKxJv6EzHVaM8+XLYtZHSJHf
gfedaApMaH58JDWuzS5ReaFcZmZ8Mc+D6i2HgaJPmiSR6TFHJt3iCR2DwumijDTT
oNp6kW3bkMLvhh76TEoSUAH6Iqcgqdu1slNZDRq/E7h2KLLrZoVjDgQnxVQMHwv2
DRj+CPL1t0wa86zxNf9tydjdaHqLx0+J9W2bxKRarflTejJ2dhH3+NI83tZ+Fck8
ECzhJ8BQeQh0+r2ntpT+yaEuKcSJUrV6yut2fiGwmktyOBX5HDOG1MtX9MQNYaAE
3upTFYlcgPGVQuLwWLNrFO/p8DzmoKsZ6oiMdE69thDqNzmlq1T6xL/ZstT+qjjv
PfTfrpmUvCf2swwTAOJecQlnjYjV9SYrrnPHV9R3pWtrRqeIUiOQWHy3tRf48hrR
BWN5I6br6JnZ9Sv2adlqL2Ooe32VqAYjn56guSpIADbFR+VxZlloCojqF/zvAdTN
pAj54Y11Z6g2qcd0wcSwjtnNj/21dOMFiFOrXVZqu07mlw1WAczDgJV8xVx6RXSi
3jwOoV7ulBDUD2BrSOzwz4HwM6OgBwycfo2not5Y1yuNpIFAVcL2pQTJblb+/s4F
t+6lTJd+rlOpRTgIeW4iXit2BhXl/6yr26R5U7yhlYPl6WkgLMw2w4FDI2wc3bVN
AQWvOzBwz6CT00a2y+6hEl7amFLa5PhbL4K4zUIn7ON27DjQD/70PrUUezz76FZN
NWlNC1YEhn/esXPXYz7Wf+qqch1Kgbcp+thX9Wm2o1LsWkfUZoCFYaG4rJSWHDyA
JsKjywu0yLy4sf0/9MNi9WP1mHlj8wtO6Zmhz7r0Zwvvzf6rtxxX0W95ERczUwzW
G7M9c6tjgr9tTGfHsovXYWdOyF9dik92ItNhdvEmLNCyEl7wJ+gf3SmYw0kri2Oe
IVk+WBWmx4ooWElOXAppXLBHA666t+5bD/Q+QYe7OOFkhTC+zDquKiBIUfQrU4uu
haIf6lFyCuOocf/Lp4R1+9VrhWi2PfMTr4Vs7LyGB/HQyJKGe1mLET6vbAjM4sGc
09uEsrJnrJ9hujm5a5LKjcHVsHx+koxeFYRsaSTmgeEFiyJDm4OYjUZIPN4tYzdK
33i2G5qCJ1z4+0RsKzqCVwh0Br0m8Wuwkee2Ea09QFyTKyrmbq5lSR3CCM1YNxUQ
517kqEYZ3vyvQ4ke+MhRKFlX0I19uTRIxLA8RhpEm4aAA6QKiMajw4zhIkNZBBv1
u6lOvugNOlgerEmJzA37uddP83WoX7H2jzNzzEDU+/xjLWVX4T1gUyKBwnoaOLWw
N64z6/mLGQuVmnc11beVQr5Xk7wFTjc48eVrRIkpdiR30D/oZPJdPu9sN8NMta3x
DCe+zdcEVht5wb9V618r2LI4KOdFsi9yGX6kw4fBnX+NDVUMzFbJio4rBTeI03oY
QRcJXqTUgjVwQIwADHSJFLYGClQqIj1DpWprM59HbhrcT1FHnz7KBkgWWP9ZmkR+
zJDPnTbRdURFmO6EQePuTIG8G4xuJsJR4/ymQzvc9iaYCInLnuv8zIhjN6yIrzhe
/IvG5IzdqNjqrpp9Qe+rp3WBvJswc5ZX3cZdLUsaVKxnoN+E/jxx70/hhsg5pXh5
3eAwZ85EqGI+GwqMiwghPN7Hx/fYqu330+uGp1mF2MtHjNo82GU7iG75yLt0QZvr
+4op4xY/BElgzpxEwnjPckX0rFMKDXd7rX1bwr4KUBJfE+x17gY05s4Udc7aTJXX
OHJv6rs3eNiaiUBStoed3xtJY6/O3jgblIBqC1eMoITH+cMlCbuay4N2zAmlvm+D
Ym9/Cj8Zf+lw5xAXCjn/2XQwN5wCV50D1rSwPBNvq83cmYiblwdQH1f2lppBDGla
QlDd3+zezoDVk2A6qgdQVvIoxdsQBT1/kPUKvtTmGoorplxjLRIjDPsWrZL7rwQz
r+C/+iRESftJO0XRDJNcxDZxGp3W2tycJZDOSV6gFTAEcMxDiCzwB/Q7THRCjqHm
QPRzilRdczcg8YizNKRdYlF79deSgS7wUe85NsOr9gT2dtK4jaKdlDKIRybKn0/x
TjUVX1vUHx30HL5ggcbU2pL1UsQU+XouoUyGkEjFffQEl9VEwxW9juoSMPCsEH1x
il+Zt82LDLIxTh0fUiVTUBYlFIl9lVbo2swiUwO8IBlcxpbQ5l41F7ISSpetefbr
nQC+l2pT9ADM2EG5RHCwqMApDpub1L5LFYtXJoN6Ph0WjBybGtcuu0u09LTY84oI
genu2O2aZKrJh/RDZPBqpDwtw0ShLmBGWQblNMO85hdmTTDcrruUNnPK8vQErTMm
CjAKq4dyClobpnKSEu9SbDVZtDyLJMq/c8irhAdrBH2qKdUeaBDqViXxktHoG+9K
UKzcZCYQYfk0WFZHYAphXR1D+bRbTQXpCnQSuFd/dsfQd+zh02yg+228JzOsdCTW
Q7ITM24/SNOMmP35dh/+hF6rULBPTR7PvnvNb7j0S5/I2fqAhlCQZfZD01G1T/Q+
Cd/7KR+P2JHo5r1f8Csf7FC2057wa26l+QNiN+KLPQQIIepttagLQiDaSmMl+exy
/ERoZnH1J+nqWVrWRch3CIlJzLmBWePzFAHDwMDOuOEtz3XPUVu0lrnxZWcsByFg
N+W67G9fobxzhdH9pvbX2LCnGGvBEkk1QSXjp+38GOasWQ9OCH7DQd7aSR4H25nb
xIGPLb2/1C68iFSRa3IuBpU7ByT7/tbubDW5xJFJFXAq3j2dkJvSvlwh0CizFnao
QJL+lvxfU40UxvsR52CTAT3NNgpIlhrhs+j8bOAZ9fq+vLSVGT93GwqsK9SL3O61
6tgeSnBKkYx4SuCZSfyFWxBqYdsDubfSatZEx1tEedshR9Dm9MNMk2tG8+doUGkC
bvBZjuowonPAllemimtL7j8Mkl6pmGVzlXPLoXbsqVElXrnc6niziecfvFQzi9TE
KG3PCyPlLPHp4BibgE3UFtqFvfYL1xmv6Zr1sIebbCS27IR2e4dLbCoFu9lorsON
CtFQ4bRtu2qo7lnDcMh/CfO6EGiDFhKbJPmsAr3hSMAELNDH931aTbCzyJeessYj
UwdscgkhCWwQCcHw2WUV2zfRY8CNf88dSQsU9YA/IpK2/zCwO6H5NAq3jx9CUPkX
KvR5lQZfVmFdOcGwQBaZnQNUI+Wg4qFmGK4LpeulgudyTDSw26b6cy+TUXHWz6yd
yVYoobu+b7ytNhjMnVW0KwYCJriR9Ymu5hDLgjpjgPF0TEhUZ3d+7GrUcba+EExH
sOyjiHoBR/fZKERTtdtkj/E68HfeGqXj+aaBnLtr4VmtH8tOFfC8vd3bLdRGwHcS
rcwvB9EF95Hpg5dd7yfz1HGNBmUXiMgdnowG7igD84BRLb/Bnria7y4wlcxt4bj6
2W4K9WQg2fOerPjxqMhAR5evdHoTF9gIzC2h2xIozzqp9uN6mcr5bjNcQGn9s+8Z
jjZNomR3uBnsEfQgiBZvnu5aotZz6NUJn+ZeTOCvuXY6H3Zwc9sBl5ixsoT3hno6
WMTe/WFyT8RlgJTjdVOaxilfQ7X/v3AmcK4g1zR2x0ETD4kSfjVvSZgqO8M+mCNx
WVt17xzBZqg6kRvb0OzRzz9ulqpJG0HV+qyHz9uxAH5iHKgww7B8tyCsOvja8Xvh
R2ApxJvQDwzuWlJi/Ww2/z0AQDzx4mIJZNpv7+afSePQeSnLpZQugsVJcbK6PkMX
trf+6TOW2VDxYOvWekCMXLXYoUYe7kyEF4L9hhpYQpqKUBEuDytp5ODjJEtYqLK0
NPSR05ZLzDybtaMV8NtDRgRthariCuguiSx7HHoyJWJQVC7WvhIiVXczS426KfdT
KgtfB/HzEf9ZTuQdAVWCfbiiPgvATHHZOQ09OjhcHKKvj+l8uAocByu2zaKrBZ2T
YxXHTRhrKBrZGOpRAy8/L7v2c6NtfiXvZgCaBkPHBUXijHDb/eRbStPvhTV6CoP1
I5BShwG0jaJsy4OBR1OhdzGT3XUGdXlVYab3sNsHpsIJbHDdkPIshyuRCOCkxBae
6/F2ws7JuDNr3dyUl/jBA5FAysvaTDRSwxuJm/kGuY4GR8sbTJZiWHeuoqZ2Glwr
k9DjsrBrIvYJ/KVp/Kupz50h7Olb+eqmd3PH5vvG+uoKwIgTb1/wj7eaLXb0vx7B
hk75QjvPXqlAgOOKaqiyRDOsFN4Gx9O4Dk92/Lq26KmcwhhztI9gDTmx6Zi0bXlC
m7s1Lty4n9xUrgzqvJpuG0+ejWAY3oMGSBAx/HzQiAnyzqiytzULmPQHoooGqmDp
kCR5Xmh+LKTJbpWNEuU8gO2uaOtOwfv3zSpfcim+75HbhtTKztz+9mMLBiXguJe/
KPFW10WzXW4E/0T7sk/owDg7LxxZiJj0E6iODDH2fi4ST987SDDwBQ9kXQRq0Blh
JEsa86xvgiqHL9eSZaqk/VXgxcOa6AUwjyJ5IxwBfpXKC+X/Vd8PIbGR+yAqBGy2
UJnrsXT1dG9+izYboQq45hmv6cwheyP9G1ffFL4RQgwKuS4tQJvpvkJxzTysS0Yl
kmvX4cr+qcv5xbE+azkNlLvbc1ghtXwjO5wGyc+R0RgAJZP0y9XTyGjmFLIi+nDQ
5sDDIexX601m4crCvswd6paYVJJmU0oXMd8Nh3npIeZCufP+3zod7hM75bM1n4UZ
fPjmXAbRjI5bf28aWDftHmc5n1x7HQbmpfBvyGvp1oHE0D4iCdz+n/ktrV5seooV
i98KuhsQCsG/JUgrdCHuyatJP3iyFEYuhdrKAlzjbTo/PsZiaWxVHzCE7YNMNweL
GugfKIBiekoOHQer6UwgHhtM6mER7fMeXVl/lwISluQRQ/vz0fmJ4P9hn5lm0vMx
L5StKtN3Y7zq8LMxFYXTT7VuXv59LjjexvPOB3IfsTfmculAM96dOJnb3CkNnJ4E
5ZDQRnpvch3VE/QaKqeQQyFCGSUIXtiL9baQs1Jz5hQ7G3ir/8mBq+piDZyuD1JV
0gYGiFFLZz8ojd8b8zuhN9+DxrhigBMPe+6kAVKp+9N1wNiNDukPuwFb3E93uhPL
76IUv36NfFgiQikHKGDdtzEFCED8eaBW5eopUrHcPtq5xQE2KTEsAqeehYry+lUd
bdZz4Erkmja6tw9+xUza2fBopu8RFqPp0Zq8NLk6iWZB4XJQemDYhJEbh3t5lJgJ
rO7yIa/UKBxrHvuXDBTKB3SIhuTpcmKPQwkZLkF/oUaotiBMVxg1axNULX6qWTpN
GNdmV1eOBa5i+UZfXurXzXyuoRfqQP9s4i7WbMn8ybA8+EahbSxjeBvf+pJPDpTQ
iGXo6zho/3118XsTqTLcNdJTzACXYk+CkeiLiuhkn4cy0HU0CHwn55Cr3FMc2XmI
eeU9LGBhTzVWHgZ7r/nwrlIS3FaTObJe8ov39E4/ANcUAuoyHBa2+EvHCMJmdQO+
WvP/WxdHetWEkBI8ohWLfCrNay0DSJo9jKmN6CFWPiaeIPd3bEC/oZ22nM5JAMoi
jh0OMeQ0pgyGvj07sX5GPzj2w2B3WXvjPuIjhv1qPmEJXpfSeJK8zqdZQSUp72Qd
F1GKx138cZAWMLuI/5KE8XrgjQXkqU/BGGBLxpDDeIzzyvkUsWikpahL8dfd7j09
RyX61cd3gMaiy33NjcQRGTY4580aej9cxtgTWAJy1RuGywCxD5AOd1cAwF3M5Iyh
m9almArpvUAlM3DsPra0FJeYQ1rPbMqGLbP6AMqd/CjhUBZR7uOVLNk9DgEiPLhZ
fHzZmK8w9ReuvouKwjajMWEzJvoZRTWyXR1QiX3R45a3wCFOh0hG7WoL9obq1OYW
oFKOz3qWnnbUEptgYvS1lpiipOHNVWeTsM0+Sf8NzQG0pLbXnyFnwEjHaBeF2aYR
v9YguG9TYUCy6pOePpTzKFQtwCUveYbweT0MYFhbKryVn9zjse3RTdAFh3GTSZQ6
i5KXGDex3x+wco8Ak4bwSENSUOcj/kX8VpWz8kNs2rqmcSqe5rlTFC4meS97eAdb
SMdbw6gKZbE2lItwzLnq4vkO9ogOhw3VyAwlL0VRtphIQ8wLj2JHz/9aDlWCSoFF
7TnWCLpeguNz8Z0z5Ae+yVUUaee/VYZh/a7iTrRXdy6nlXK5KO0Q6HIFNat1x4fz
8fb547t5ApqAxPqVWS4A0Qt5HCa/8b1STxPRHgXunk48Bj2QyRz3hShvy5ofGLwk
F9lmBQJ4lKHczlZWYyfCc0JCyGDXTSfAe/76BE42uY0f3L2jJoeOVshiSKUzPGtY
fdVu2iNrhdt4m+4fFqdMeZi6uldRXx/5rR+wMxpCGXVn0x/foafz/soBDpnupHIE
G1kohl14lQWV2BZw+N8IUaCVXgpFarbw0r0E+acdrUSnH04inlkYRmvJjimvY3Ct
z+rM3NIq9uum3fHKJ3bOpkZXIVq0YVDbAonpXzRl8p1x0E3kHmLWeYCzYSBo+IQ+
8I574NgAdo9fXJV/7nh3nARKboL5tVLggr6x+cdv2xhH4a8N/NHLdp48BDLX+vns
StG78W/sAFwIesnUMRr9XPPHimow6XP8p3hMe3ZVsTpU3L9Y8w51fPXypH4U9Bap
U4XocncZ04sNT/6Fj12ubx767KxCZPQOY9UFheMxYxQam9kPOFt/k42AU8BCx2mS
iAF+TfxU48K6FwfF2E+A0lG1xAC9NNIKt5PxOFT0lNdk4GB8Ld0CkdGSF9H9Ny/d
l8C/IgafVHCprDO6F8I2D7d+wOcucu2kNM3iYANhLpnQhaAR5zxHNQP/8xlgkJ6B
/ohBPBqkAz9X1tqEfLUPvza8Rg72gz/D9+04ZmlZxhjk478MBEVmzRteXVjR6K4k
+wtKAYnq6Qji/u3dvB6Y4F2JODV3qw4uNCrd1kSqB5Wbd05wCM+yafCgD7Vc1TeB
xRLpmqJqOJlQ3AbMLr6rgWYKBEZ9dlTOu+Bn8zObuF2d1QRk3ZaYrxJq1BQX2X+p
J2srQEGnfqbi32A0GO0O5GfL5A/SunpwEu+E35gnwAn14uaXWLBI5TpsIjzEl7uk
m2g62sTb+Wsonm5eDXq2kHyPYLd1qjjMULoq1yah+qnqnifzglNElEQ+1AUYxyKK
+v6I2XBKiw1rHM+/gkhFmDZtNrizEPJgRYmI8QukzSNMqAmEk/qgvfVyzgeNs3CY
6ffXYY0+69zmT/GMGInVaopJ6jl6QHvMVBgN/HsljEuME7SQREwzj4f714EyUndM
9jWA5YbpBD+YUBFivjJV+j5/usW/C+GEg+iGgtUskiT50MaxvAO7/qVHx9aRvz/7
BCyWEcP8pGQ7189BJq+2Lq0pWFdaz5Jh+d/FQ27mhjSciE4Y//1HrUZDfJsEc/du
Ifrbw+oS3CYrqI+KGMqeaXQLjmK0VfZhQGDif3rizfXglmvkDge5FGt91z3JobzM
aiLB0AS/GKbUB5J+LvqdLSJDUfV500T7nYIcQnysFKGIGw0LoUfjEACeWUrdYcCY
KcmmqKL7afqp834haXIAKUpOcJ0dGdPCJkqSg16lcB3rIx5elWWFEPAJM8+a+11+
53h6SWVgPnceaBkHFNT56FsrNlK1ex0XH9lSREmO2sDQnrgIOcyGDpmFjnoX+v/5
E2ltItj+6O8+osS6WKSkddGzAk0ls/NR3ZYXKj0VYwa6deXu99fsDuGnEtu0AEPg
+qVSsD7xPjg4P9uNm8uIZuRPcSACkaeBi7H/pmJ4KTgDcRpNZS2s/QUjr6iIGTRX
Re/aVkBpBmOCZbEOeY1Gj3HEF10KdBArqwxwgbfeSiiOwH+TSzH1RrQBT0CHuQBO
wuNpxLIN35F89+Z1CTxZAGxPmOGPs5Nuj9QBUGs0s5gqZErcKztNYN12sChCu7uT
05skZqR1YTRB0ECbwfNh51m2mhv4GRbF8aOXJXfjbApV5njruC2jdgGsswuC1cPI
CNpiZDtM5KCf8ydOPkmB0EHKi0j3DzOcE+xEBzpHh3zsgTBKTb8mwR6uj9ON5TPe
9En+UiNSlXc47Nm4cvmbhO8c4fi/oBQQ287Y7Mrq+hwtQUTrmqRdKSzQ4eWYv0Jo
W8dk4RTRQuBgTmHqBGo4FvEaCQStCI1/cWqF3NHH1isqGO/y7RyS2aaCl3zXQ3vm
Po4ntmsg4e3jdC/td+oN+tkGLF2lAs3V1PGNrjZXq5A541C+4pTfKvWWVDJjfkmm
GJMJ6qkf3mPsr8ODoY+va57QXNlusHfJhhgv0gghwFhrEunoWd6D/3QNJBL+j3zl
Lgn5wxs5JuSQ8rsoDv7ozsUFl7Ps3cLCC//jgVhQuEsewQuUN+A8O3DTK79S07NL
24pnEJTZmxrwClD9HGmxMEjVHhpui8njcs3qeCOpLXOKgOY+xPpBXDFziiAvKfmB
vCu+Hz4KwsAfRrUb62s+0xc5LO4NIxY+wWtO0SFYPmmAnmWfqknGOnXxiPmyOD3T
F493gu+YNbSOvZOlfXyjK04ovTLMwW5gtcvOVoboDaDSyErunnkNWlNJJ6aTxAhk
8L3vlDylbsPh9Q/K1Wmm4Oddl/28Drs3Y2LMkaSVlYUhihZpPuVsSRnytpRCP5qf
VOaLHh1IoCnDv8MFf3WK4NnbTR7n0ZpWhGqbKt0ooAoah91sX4Ze6qopg6gZBKS8
Jkic/rvko9EOTIrc1LTiNOHAdJe6+gXPyLbt5lNV/PsPE9FPN99zMXPAET4HU99b
5TMXkt+EFAr1l2R/85sHzOfSxsaTRVxCLEhsJ6Nd7nyGKxqPp2U2p0KfhL/pFlwk
PQpXNJAnOT50aoO1TTqITaiTt+lnTX5pqWBdGukDS+f837rSoVvaYPDLThgnetDZ
bfDQ0xku8nvMyMSPCR+ofBHbjmZL14xjImydh0VW8+KwRdskDx3ZL8Jx1b3N/VQs
b7jcTUWjI543lsXevvIOq44854h9HWerI4ktodlYyjlAv4UzBMJstatSBUXOLV3p
9lLZIFjzwb8RtZXCvWjVWhJ4veg/G0y22CGVfyuQn/ZiAMHR/q7cA3vwQswvC2C6
xID5xMTUHlRG5jKzazw0r76UEsbAVJr4cda8M0hx2Jst9fdS76a/sCzdWGfddqrL
PxbmvuIEB/mgL6qF2Iwy51iupguYYjFFCcMch4HqXwppl4jDU/WXqMzrDlKh3OCr
Bmxn4qXNLGVa0x1Qj2Oqz8/wEZ9U1ZayBNl5/20CERqatGvFVbLjZ6vp3hxcq33X
DId6/IklEF3kHfHBQhea+eIjrAEX/qhWmRUwPApc8tqrH8aTp53gQrcRFx0BtGAd
ymRqyvOcEcMi8PWTwEXP+565jw3vdhgQ13HeN3jpOnXJazmZ+rzb/2xjd6zPhgIg
7QRFP4mU51UgvEFSM4K6lp323AFaxaEOE/8EM5tNRbqq/Ja8E+D3UG3HqmTJJpuJ
Pl7AaOLNJZyaPMLVGDQNQ/keMIw+uZr5r91mNKHc0X3FSRugqv+snBZssYzkc0jU
iTIGLtI0CluIdPrwX0fghxF8TEGyOTKQWcWx9tJbW9AQO5AoFAKDkn2eFcGUqnPM
1kgqXGtGhqPEB5tMW8ocCS7h33a5PWtf/VkZnwdAs+n27D23eSHqyB69PFZfzvHT
d6fRElchw/d7hEwWR2c/TDLpBOmHMcTtluc+H2nanheGg6at+0JCXYCJCa6NlWBh
ANDu7YshEM6ao0pLRjyevpSivTqf6WW7KzyqBHa1BIFMsO5eI6ad+S2ZWjqvAjvQ
FP99B2lkTX15wizH4eDYY2cSrV0LLMGqzsjntTG4UN9v2gGx3hHOrB+iXUooYwpQ
sxYxZPnJwlu9kwKH0ZcZzvGwWgrbPUyt/vlaHIvkjfSrRyceFFBqC2ohrUpZq8xl
9udExUkQDr9b2Pl0rzLjnUCByrBBSfonI0VN1mQk4dhPYCgflmkyaDIk5V0qE6fk
ZzIcEqE0svatcmIbVBvaXtKby/JW135vpfpLEkZ8dImQ7i20Qh3WHp4waFdi2tW4
AL/18IefAoQnM1mhZYWeyN2ZUZDFVGV+NO3qfk9+Zymhgm5jV4kRftmnsraKVn+S
glOcgZMhnHIdbRor+50eRp8byFQquF53+q3MB1UbA2M6+ZdGCd0Z5S9Ttw4p86fs
3AKCY8SvAgYzdnNfSyzF5MDRoHXZYPBAOn4ZPHqCA48N4LUdUxtgfHwEbC9xBYTB
RTFlFF94//pQNNjFoMkenT0D6Oa5lBmFkqEKvH+1u2DNZitnZUIegbdSduRISiLu
4BzuuOuluk9THf2bfJjnib8bIXAcDhBJrAceVg+jPi0AWjgwmyGZdVYebGjU0iHY
IZhelRH/BLCFDCNvRh7I/834JHere8MvPKjdTn3aX1K20r0PNxp3Xz5kPmASQbz6
wmkejIuovwEYIzSzneDjs8qaq5ndfBHV+7JnHu6+hoUM5UTeqr20Yd4pZVoFXtRT
OzxaJwS/awvk/UCg4ZuxVaF8mFoNq5neDbkCm9+Ucu4ZcGyHimUiMTOfdiKae1nQ
svIMIIcVGpm5Qi5yEAFNiR8ENdZ+Aevi1BhK9ebTmRlvIikk/f+ucjMz1YVWK6pM
SCdAD2Q3HL0YKi7m9iZlYDrkdL3TrivHe5RIpC7kA/nVyCAKGR9skaLXMM+qyXJW
ioqfelLGglMF92NPUO+6Z8rQBDhkTpkAiONprm+ZJ1aFf50aYPkQnGVc0BCiClh2
k7oim7+uHGN5BYP32mUlOfRmsSg729wMjIgz5HCgY/ZW6M/D+Ha5sYLsxVMJuX7H
ZycLCTAXso09vbg0V9IaxPDBofszF+nK+NJ4hJvRFALlVep68nM03UERCtmG/l6/
Bzy+1B6qAi/JUk3NgMqvwbpHt4Gnw2olhqYkXwc724O6BqBs94OGhk0+Guh2f70q
Y86A+KSe/s0MnoihIdmq3lX/9OfgFzhU/PccusdDjY43wQu3GiLgxaebEbiMOkab
94KQtb1NNGnlCTG4THX+SYMYjEBLV6Nf8+TBbTLPS8jdu4f3/ivb3u3uJFjcmLiN
47zHjGt9RgPorZ6iziWgChahtTcMPImkHVXRG5QxOEW5Gt+4PEIupG0k690uc9Je
tz7SoDMLHmWI3jE7PUONbDZ3qDJDr6ixxVzlWyMU5DpX2Livbk8VzpqdcbOX2Q7Z
8+GlpU73Ly9oV55cvvZun+VuRRRm0tdaFdPeVqVUmsdODOWv5yUEwFvewvH3ubM1
dTfWPgBJPVgf3si92rP6MpOpReEGtyx1U4WVanusLSLCip2LoNf2OZZn7WSdBDLR
a3Aft/7V3/sKTtKTah58Xze99jYvOslIhD/wukgM6vjN0qKhipGVNVckNU7qW9cX
KfZoh9LgN8Z/XnA6mPcfthFsu9NL5t+dEnGNEZ1fKXbO3jYnUeVwvjI4E12WEQt0
OoOF0Ih0OfmhXZ3h6oYym7IexvPHnfofYrwM8gDNtilcrb9RZVfFeehere8i38xa
47KtE/dDrIbOYn9StEGQmzUg0GO0FSB/RDCa5wdO5/f2RvDyG+v48+Pg+jHwaCDu
6xHomEPq9PptE1ze/QT6mZrxLmgTlsctTsdJF5T19B9FkffaZR5YvZnsi0YAxj4n
q8iNDt7w5yH71TrRX0TZbvBUFojzb8ep9lpuqNIslGndbPbRpkhouh5cvwUP8GzS
ez1qGsYQpDVf5cApt8bXY1+ijrSbYB9s9qRT/uIdZd85e6GauxXzG+UP94L0UX2e
CKTn4rTPgncG/5ga283YfxFMTeRywm0rmK7lky2S2W41phuvF843sT7XiA+Y9FUK
WsFjIcABC1JLcaaGvoDji+ZowiPQ7cckW4WPAfPIZb4LYfrmCCedMaL9mcMENviv
DWy8farr3dES9QORqt8tmL85fHpZG5u8zOsi4SdeN58CGQblameOUwsiYNf31zB1
6gjmzL7SPr6GNAEheDGHGo7o+MNLE7+mk5zp8+lCAB2u5PcF43GmnKUIyXNU7VgY
/Y9ylneMrGmOBNTvmeB32kLYIuQ3g8zHfGGEPemd47v+ySX4Hg1wjwJKZ5u5TmmE
8RpKafG9SxI31L9RWrzn6wzSHz+/QIbyh9p4lbC7apAxt8qXq4MdF5zCpDatmx26
G3J2KdWL8VqGFqFn1C8wUgH1KBiLVUNJLjnspLQ9FOKxUY6XHJdUSuZphgpSl7ai
wgoZKT4WXIQQrtXQZwoN+lM0cnnsR7vpvRWyo8qwQcaKHNfPYZQ1tQSnCR4aJLXA
p4p2Mm+s7r171vTrndM5hPVEgD7iTUFf1aue6a1XgcMSRmhYh3A4QF923st2FsxD
KVBPwrqdEOdri47HS923hvNF1CqV3iV19C99Dx3meVUcn5jqQHXZT/ARLRrjc/CC
mUMWvK5xpbMV6OACfudYGQYGRyB4D2RPwViiy3SgdjbCrIAfVtKZ5J3cit/9F74f
XckY46MMPiYmPznCFYNFDCh++zlu/mfxcnY1ydYTe9668/N6VCOKBrqWjr/Xksw4
CWCAb49L6Fum1Q5FNrh1ochpJu0izvsjpXVodqkjuB0mU0SxweQqsP6roLKoPXPL
CPv10wLtIn9dt93Pp4VYa5YwxtvpWRMqudm6H38qq3nzmUSAdjAG83r5dnVKgZgI
L+cLrepj170zIzLgMhPMIqRo4jPwCIl5EBDW8tN37HkfPv06buBu3MzdTQGGo68H
LHzCwTawPa3r/afwi55tV9jvyHJ1GpcA088j4X9LnBtlFqzYcfYF/wyCTMudDDJW
Pu84A7FgYsh3+6K+SKVOvwIgFBt/3WDpFgJ7JqSCk/MTLkmE6qhI2ATd2Ye/ZRxX
GZT6gBFNShwtC35sUz6Nm4TQpBx/aHcjOoZKraG5kPNEdEReWyFQXLMTjvRWsL17
UOizHx9v7PqHdSsNxZR1PVEQ7yjAQ90EOF2oIlm9TrKMhzeAcUxKoFf6RjitP++0
5Bsy/can19+PQQRsS7AADap7dviPK7Zv/tmHFwDH2AP1zVApNOYd32zV2U/4ouwS
GcKaushyQNf8XUzytmUTGx1Jt0goB2L//+DO6fydTP4fPTTDDJUYTKEn8r3wbckT
OwwsQehTx6rQ1iNOX0vemj81/XwPDFWi2FlYAyhpghaaGraqOiBF3DvjMDmvBeIN
4PL779Sr2F4j5EuBrY7e6JcYv196R3HfZp47bFhW2mLA2ZvLfB2PBsc2f2xKM/FL
oju4y8DdUxJRAYmPo8+ZsPrlDhK6AokFZJzT7oymWZXEhoI4wWq0txOE2taCxjYy
L+aQHS2DNH8HJ/vGR34MiLt0tDQtiYkOLxg6pnG7yGZA9GNTwLho/HVCZ1vP5FQ8
heQt76BFLaDXDnF67TGbqnjYPCAeiLV3MQYtIepJuiby8Z1wbB9/UDZ8WVy+c3Jy
JOEZSACJiSeKL4AL8fJ4uYuqivNBMkNTC22mPziT3ch7q4iKdMp77Q8VGKmVWtjI
dQL4AtCKJMN/uoKqJUS4f/ISpX5ma2RBJ2GZ3edY7y2UjPNfaywFfYys2shRcxFG
XXHxuEhXcxmuW1hMHmI6ixJNdPCaxalgflXvEq8W4ELcHSB+YmJtlNnFEUToIoEN
/LqVrjDKehpX+05stsD3tWQ4WfdqgpA4IX32LLhzyhuFY7kYC/Tq/TfRAmPyP1ST
5pyYIw4jm0Iuu04x2RQeAF+7xyKkdesueSrFImEpidluZG6VlBnavXh9Ln5gx68s
QTfsIb9UM674EE1l2kidqfGwamPEiWEP+OqYr7dzhlacDn7jc5hw7oeSvSZQAft0
lPPirNIGEptrMWBhHjmuLEyIm+Mq4rmt/8c9cOxE52H09NdcXmjukfRM038VON7Q
2Yff3uSfs0zVbtMrqsp+nQWFSnGL08Ylk9OdRTMB8ySIj4shNInLvASITxOxVUoh
omCpdwnFSiaA5zBdpcyPXOs90gdHyiriCohZ4BgBRDr1U0zqFg5a2AZVlJw6nEGm
FqkzGi3a4XEt7IBlydDqfFydXeyPt6qwJZJ/XgRtZf7cyXtCVVWDcUiTxoS3CjXi
cwjd4ClIhegyssZCGbk73eUrCCC0fm+X4zm2rg6lGkSRF/NHVYco8nbbB+hZ5jBi
AqEkoMWpFXwGofGwYLybP+OzdkoVb7UzDQFXt4ja02a1ZKd77nvUvBXFpJv6Y8jL
XXfZR2YYSo8FOXvGxLB9Jf/eDJOGc15hgWmmyOZRFp/cczy8ZSGMkp0jFyMfFLsx
iVpKWhhDuCzGfs7OMzu/F89iESQrt2hzaiF7YlowQCCuSXI3qV8KNiGEyOvTcYCA
kScORMoPEAKYxUD7jPGroWI8JK/EckzhxOvXBdd1k8wgepS4XhepfG2m24ZUU7Ms
eiTcof2VVJWLJwp4khcoUjB38XbRDHnYujsP6pL/Eh5P5UOO1/nsa2Vsm4UJHFRk
lafoKU2r5c/wNmnINlGkRuD6McdWPZDosvnkjlP+0/FPGyKQplCyNjY9BtCrhnG8
6mY+ltOitpctwqOfRB3eOmdGbk9xwYLcI8dgjrotCO4hyjEvEWDmFZO9S99wuxty
ODSnLeMyi4Xagnu/+1V+9WLytb1JOC1Dm+McTFUY0Mtu+v+DzCfAxQtS2xFc8vjU
001AVW7mQfQNx67imYyMKTN2tZeT8XfGoYBrkEhHW8GNl/DFXn8Wlm1IF6jJeWUD
XLVAa89vCqna5POQ8iVgU/HFwm35gldcfb1WS3gWLAig7QDe5kPN1QnDByRPwssD
CcLzDtmwYKWwdteOdSPCSWr/m0NeL/DVCAm3FyFIG/+jAulCQ6Sr+TMrFKLI8ykd
CAza9ZXSNf/iJyZBWwF8ajiDwE5p9bArYYBl0r+9K82HulDRyjV1NjSbyhea+Prk
iSN33zDit9rB23AAbKHC9oIq24xQImpqYESxuGiwtmP/K7lLZZM2jSMajykbO/rH
6SplMmDwHXt7TEvsE9BVcA7tlb8Ot31SI+W2AxpemVcvPPIuvjiDW0i8VRur2jXf
7DrehMwV4qfYEVZmOOIT1B/e9y/KwpdvO0Zadu7blqRl1szclJAVE5FPIabHsiHn
j+Ie41d4z4w8FqgtZVc/TtfkCE2BwtDR2Bi91T/ei+YJVL1NusdZiHx0/JqkHFIb
ShzoGesgnxBXQPfvdHixZgRs4Eo14v91V0kSi5G7T0cqJgq1L/IILfyyuCoujF5c
lq5i+zwZMKdlPRMnl7Pg78cmZFuk0bTkEvwX0Cw0Cwpb3cpp38x2FzYf1pii/Hg9
r1MOYCzFyppgX/XeLl5aO0i0jHWp2FibjdOlPhL2YOQXT/zMUvC8Zn6rRDO5eF0j
y0SPNLr7nfjYTIguvP2a14WNwdLxL38UD+6Olh4LxMGoE7n7zKZFPonrxDAUs+/m
oS1oV3EZCt+sbmDW5vBkSRv/oMgw5NEPrSyMfW4QJnp5em7d9biSZiV/OhyeAROr
wBlGf/++tdbBKrsq61JoaO17qtZMScBDbR0EKjk8obNtY3Q/jhNaUyCPvCvfzZqP
3/xU04/S/7XZOc8UI7UCh0evSdsjlZR1fAFQNEGxJvq1WT8KeCNaXGxIZbE9Si+T
AMwkqb8LMRZEc1Rl+6KPlM0U20NexXFBd74ppxOMRvUwi8jKDAjDbIU+uWgsUV6/
oc8qQrG2Lp+OwtYP1Cl/ildT8UPHhccLA/t8NEUmW9JMZ0+fuRqR6Sfg0W3yEwBQ
K+/5k09pRuXXUhb97QhOTQuR3/FBBAK1TcO9mIphx3woMnWCJ4RQV8qqzFaMJPzh
ijZTUp9HEQfPvHYml5GefAtTkTBTpzGk6q9R+i8hVRdSozVe1Mpjqu4F5heREECD
myiaZzUtbYdGgIy/lrbKUbkN11Z02wEfYGkHkLUaGzJwugyz1YFyw/d3k6UqyvfR
l8IDy1ywQ+94tBJ882AP+G4gdR8XKvJ76tfAs37+FxQAPMnr9w5z9e00iMcPmPO2
h0COsb+4yiVd2d9TWor7McH6l9xrmiEfzX7k5bpXjlSOEFScflayxe2C2XXrURSE
1OtCJUiLGT7DXcjEiZypXxv/UIfbuBPcQ/26Og8IeT56mYEqjce7SLF4NOOKqhos
9iLuSWBcFgWxrwRrib4SQ56vq4U1BCQkuvZLCschgYHrClVBjfSNnRhu3+/GTf6O
9GxdjVXggwJ53Kid6r8UvBK+05o/Pz1ZN/Ec4/QRhPv3wKiuy9zen5PB+2k+oiTs
HAFwbUOLm9lpNNC7lUaKf1gSTTZYe3KULLofL2phOtr7FoGoDKpViXKa3dai/OZg
BFvWSqmyeiLoM+Wgnq0/Fc4GFa63s3p5UtMpnOx/cZGjn7GkVSW9+Gk3VtADs9hr
3zCNA+7DUUck/GjmXwPX0p9sYula97FowapWop6nOFOL0OT8Edgq2xT0n8fIlWHG
MOnEA5BkeTQteEF9v/KcCGZO7jylVSkxdJN6k8bZorc07vFq1zvgqKYbiQUj+gih
jn6MaPBMkTtFO+pDkVkCukiayeZ+gmIlOZQkal1K7T+gsHMEU2Uw2CwnfUKXUxvY
TYwFhaqST9VioS7GzmtBjucbytS7yB3Tcw77ccBLxK1/ljfX44rxCTowRwAV3ieI
+ZkbbqDSLGrI7PpCml+7cDD7QABB+AmOdBZT3DKeOW9qK90OgdZCkeTiE2qavzAp
t5FdFs0iT4WdNVXMnNoB6HyWG9XAmnXqlhUYk8suX8+FxvnuC3TKBX/R+d3YAKye
DCYUeB9OZ/qC+Wy+A7MMlF2oD4ZpDxuW1pETAtomkSWPLybybyYoNcNpy2V+9teb
S8ediBjv1B09T5IsapezoqqPq9o3F3GU+91f+j2oqNVSanVUbzEMUne2mPBJSaC9
EJboL13/hlc1+tgv7j7TBGh+FOjXVgPDJnUAd9mHLEZTkBqaYeItdotoew/ul306
6A5i3Ah1PmuBgjdfsCfMXrdgbV46QjWIjQ/6fvAn2n0EdNeF0mLNcDzOB/lOblb9
bXnSPJInfTrTt8mXedhz7fCo486rfYDMHJAygP+hg5Tvxj55o7/p08CBsEe/dREk
MCYI4l6PTbNh7XxR561YzHxUUzn0m2ZjbLibapuIhn3JPJowafHt9P1esSvYfFDH
uSPKF0/MalCnafEGcIzwx1EVvHINo4GLnDU5XgvnFKDGqQQg7ERnIdW8ioeqP78m
fhy6muDbtCfbIyityvFuYf3HaoHcrjCGOUts9lr/m+tV7d1dgEb6c79dH1hGMiBa
owcv7kZ9vcyVzqOs5XJDCFrTUb1m7G9ObnPBwVLoL49GQDl80Iofo+Kq/mig4jpj
GF8AqH8W0qOOgti1hEVECSXOoIotDj+yyUdCGRpiobxRuz7sVeNZRmcpUFgah6oc
U7cqDIS2+J63YAYftYtXbo04i4t5cTUzL/WLVP/MVwE0n3SoFCBDQJw6ilAPZkYO
6lQ8exEeUfBLTZMY6b4PF09e/9P7Nxcj5umsbK34/ekpTw/88KTTmXMCwb0ENMhZ
8C15u6tAizZzRS9U94Rda/PbaBa0EwwU4j5R4HKPJrE5I57x2YR7JoMAVmLY4aNv
u0/cetet5v4p3J/zM+UW3L6EcR33BBqjLJOp9uqRwtNxGS9Oetlz7R0r0g27T7ZU
T7xb9sARYgD1YXxZaJX4X/+bra85dWTPRQQATWKs70YYTEIbzZ6nJLLRI3eTsA0r
EjrcazvXKK5zyAO7YVTsYPBZouhUNxcgUhNeSbzBUEGzYCz+Ox5xrd+OGz3TbxuH
n8eBC3dkwxv6C4oLtPZQsSLThjjqctNPw3riiUsKO23Nrl+neKO5RCcVF9Jmzwh5
vk8MKMU/ZNZCLJ7CGOL/fVZWmhcW2TrWdXiJcslAn6I6e/XnTXAJ3AVjtSGipXHW
m5jkbjplsBHIBvrPqGXqMjqT1g12esT9cnhss8NQWGihGoNoYXxnV3hAs3YeEMER
fia1e62G9Iso/0VEU6YxlZAMSBKT1FS4MB7t+b9gF6+cDCgyvawtxbjsGWUlIQj0
IddfAloUW2njevUgdRP/56tJ6lq/mwaNFPoa6kmkWxhHKcKlavKMY4hoeMPVGmTN
ILrwmvp+4N6GoEN4UyM/Ua0fJc9lllRyMFHriCXRtQrro4jKDWxw5IHDLo+91ecv
mtJxrA5BJZWkbje0wp0yL95hjs+fjXdXDFUpiW2sPCH29SX4Oab9GMbs4FTKdkvU
wodxCkDeiiqhfxiInY2FCFL3lmpfQXzQgr/rHzSXdZYgh0sKzNeeHk5bYn0ogWhi
0+Yhr+3CUPRvab/gyNTK/n1+9X85JfT/u5q5pkuy9stW+u9N0SxwvoPXFqdTF8Sb
kPsZEEfyl0B/1unnfGi0vUoWhGMgIzb5rSxceoTNrhGXDrx3s7PjlAtzalQpXLee
V4VKZfcnkDTIFAOcpxsbUtG5VLdh8ldcIQlLAMGyce8ZsqkjyFFhZVldOQOnAG/U
g7tSuJ5pAuUnyqZfoNCBU7Hx9gxtpNG1ykv6cyitLerGBFMhaRNezDODq+Y8caqH
6AOLeZRp1UEwvd09BGlZHF8FdaDF2KXVA3nYvqvPNfWfG5mHCkAQHAISuTPPKGhX
j14KcI9qR6nKUaYRr2MAPOB/jbik+2HZ/UddtVHK+1t4zqIfQiq9YB6SsQe7nO7T
zhizy7glw9c7RNgiN7+SC1mJz8YVA7GYfDhiS5Hwcj8E1TZEzGu9e8wL1SQzv4Ep
4OjngNlUvDwT3ybsPzZqHkd2tAYIJLgIEJ2OM29aXITW8c9rYwjPhZfBjXFB57oD
MkX/dsaHd3uhKfB/B6diVeCb3FHJCdkD9ZDltuel+1ETkD0nc5atisFzSJRmxuOw
RdwLzouwa7McUGc7QHFMXcE6j6n7vakYjdf96aSu9R0JGtYWMAMcptuJGpK3M6uU
RB5mluqjB/5VxkgrpVdaeJFailtYjcC5QTQuE1b6xLUfyuH76uoaLi+c8nrqwxti
h3C8hfLyUxBDutygPM9qmJugYVtLd3QvHZRsHBS1VgUSZimF99TVyf4YOOgzFHSr
yEuWa4zGGUwc9jtRdYB54WDsMzfbWjdyrTQrvZT7mYQ3+64imRb9/Mae+C8H1axC
ZirPhQzfQLpsmc2ZkImE+1NjVbTngA8ekvSSdzSl2O9yiHv6wntW+Tu2mwUN3UR6
Dy0cvLzBEolNBf9nobCUMH4t2cUnCsat5v6bz1zK8koWPK1XDbbuLdNYFnaJfqw6
5GPqnx4wf0ifFjQqv/+dqTee0u3RA80TpIAeOsEeGgYALVLSoF23BIFaQ2z4rtUr
qbBANmiHzZa5GSm3xmJZvyHy1hfyoDbn0yBMbmyIkPK3swV+pJ1Lay48Tf2fOMzh
HOFVgfM+Y2vLZ3d+J5SG0WhOxV3ADJ9V3c6+lnlPrA8Vsui/hwp+eorJWyWdm3qr
cUPAcZl7a6og/uhjUBnh/bTj9gQMcyzEKCFZf3sA2jL33Otmt6SAPNBrbZztXP22
nw38PZELrWftVtxKPP5t52/kH8z66+nXFRHDFwqiAEoiwoQLLEY/BqCKPYFn5fk/
lleii4nmyvd4N2sqvnTmpHO3sVcIP/6wXJ1PNdlEQUHlO7JNkzGeEf4PoPLUA0K1
w7eGrN2LGOKPVLvE5lrFemfXNqaFLBhqO77GLZcPOxO150VaSKSCWu7wBCvtz8Nf
HwXs6DBnSLeUZsAoyIux1VTJXROhU2BS3C8JUULlclR9krod1i0SwVnLpbENIZXV
/l3U7lm5ZrRqDFkY3BwS1qLwDdwK9V3+7N2k3/Kq53efa0/OgWKMPA2q5bQhKPSt
v8kpMbIvgc+1xGC7C7BWN7+nIia360+jhIE8/gezEFLFhLEHqGpAVkfeXRaU//9t
lm3YjNL5RVemc6PDGuR6DFMgWwn/i1ESe5ccqlJSlyl4O3Gnnh0eH98C/CCZihzm
GBVon5fHuSFG98XY72QmwxOsNPFXoGmx2hp8kRTd1aBt2QKjV3hst8BiRjtltcX2
dimrPwyYRtpsspSflWZ2gUYDil5jkw2WrteeKqZYlPBGWiw6wGHptV0IJekADyEN
kCMWjMtNkLSt2KmqV2U2OOtAW+gh0oNj1pOl9HnmiU/K2F/MAGUHQdVqdxigxbb3
a8TyOVbwcRzDYU+WRiftQFjYrBaSKNynbG4SWtl07gEOqgBHRE9+j84+ZEf5Y7yD
y9bE41FOf0fQQnbIzEwA6QDX/dR2unBAya7FcON5r1z50obk17vaQpI8lPOjqzmh
1BLRA+q34FGO+KkOoj4tXG11nEseAoaMDxU9Lzrb0wWDWzKC+Gza5pd4FhBhKAPn
2pT4Iy3L+aDFgrCGwQf2qVBsrSFAmzivRltoHGZmErvlPHQuf3y6qH/zUyITQAoS
5tmeX8Uka83QRVJUjVaWvzyGZa1md7/5UclNHHeL9h86PSlxDiTBLscOQ0JFpYNT
/SBkddVYZEgNp71tP2MtdxWxCGbA69xQRwSBbESAHeMZU+4pC4meO67wklhbqTFU
KHBEIjc8SagJxu+49W/wcmYXkCnX+p7wqtWROeCmAXoSSITnxn/Zr38BNasi2S/P
RNplCToRbzxQUt6RBsV9fy4EexnwTJV7DDKFgxXDAAZ1Iq0cxRGJRHcIVqtWRYxo
AhvkGsTY1ZB/8mKNPLJpWjedAOkc7T82QtosPJG3O4SVR8EN7yER1fSyfyCTNWc8
5zg9UhQhOc6UYs00PgHZzHAzDBRYSNpM6FQU6obo7M4O9hsh2hW3hHskCaM55fBg
wuS85gB5E+ppW4sDCrsw7I7i9W0Gpb6lIq2bjAdwamFCnMM3aUjhuM8m/vnW9y6M
+rXPBqXBH0+fRBXp4evp87BN0eKNC2INH5CKqj2edJaRxj+0HeCMR4bMvj0cFB4b
ZK3pub7ncTBLKdmjmFMHIufBbNRtiwfgrVV4owqRz1pTNGbUCtjXd1moCtjkc4VS
3Vzrh6qGqFIQY6NRWtx6rK6YhvOtFVx+MTDvu0glCx0PpWGkgcvCx+nO5HEMGKjo
K3T+ZeHaXNF2un3xVytu5VJTANi9Ec54xtdiVIFas7Z6xBMBH+MzdFO6ZzGYldW9
Mr3qCczpYeQssYZcZ23YW9wIc55AdV/d2x6oFi8UY1q/kvDjLsba0TkF79q+ZTkd
Eux970oT2GKft4/yxbbzNthzAO+ErnGe5bpySFeXpkgVZEZUu2roldAXjc59oWHy
c1fBnmj83kggorqQeJaOwr1E8efaa1ZO0qY7DJC8IEFkB6ttlith96jepfpwogMN
BjJYph+SafAbjcSta364Uox98YmUscqT3T88R3TGfDp2hQaGAkGZH4fbygoY1rWw
Kcc+wHFi/lYEeln2L4wJwyorU3I4vdStdFdOxxccuZ0zAa6NhPOyoNVE9lhh9SNw
Dm2Xv3bW7fL+IiYdfmqp82rextmS6aof9FYSvs+PuftXQcxlOytSWqpXVMl/sz/A
0n+mWd+iyT/9llftn9z96CxaTBM0eBifL7rq4TFrsyiUnv/4nm1jvBJxW7qdg2ua
au2mbX6zD/Dqrl0ZNUSupXsJEs5Rrpx9D4YLBRjuRRETmFL1dx/TFb8N4Npb22m8
OydazJLpgraTuGFfN4NLVlZt16WO/15Svm3tYwK1Vku0d0ZIdeUisYMKoXZR79OW
paH/0IvBEcitjeIwY/NSMsULwNJYOWVURYxrmT43ir3dRYQ5/3KXtHaeDZVXorC4
JUuYN2OPFTVQVGC5mj3V6o8ogcVqZsbbhyu57gavOD+PuLy/jrM1r7i1pV68cyUc
5igH1ZzcG3nvIWGYJnE6UdF58acrYx3rEH93II5tAWaYP8XCo1MDElE2/HUP8Rq5
xQ9j5GGKFC0qLbmqkHMTMFTCQVSHsB0P5/RfqCKrbsUG1DsNa5tEKNjw9bp9hE5e
6kPpyTjUVVPTUlySr+8MQcZpGTiTAbuj0VNRNkBLRvzfh8jsWyjBERZlKIC9CeMm
QdjQQiFVOFblSPf1n+1e1Ga8IdTtn1nKKahm5apSa/XLagZpbY+0rU/j8g182CoQ
qh+em1WR5cjQyj7OwVk7lVIUlvCYyCVUQyyEyxoTbekHez+j7RRoAjxWPF2FEd7D
YU+MxseIdulYk9LOUvroWppALub/jJBJJoyDd/MJr+CSw15NGvNDgHQIry0zFbtv
HyZ1WN5uvEGY28yHoDpyy9S7mi9xMS7WJD47mgvSzo4fK6Pu8A7Aob4PSgxRBvRA
HNUzzRo27MJq0MVoAxFwFd0ABm56Fh6tQpyoo4CXjn8geSWfflhKO006TKBfWPVD
J4+JLpua69DAM1lUANh/VlyhY63CsTimYZwJ5x46gN7YW9CR70aKFRdHtwg4VZNM
ccS8ycsQpIx3zRexqIlesgUwLwZbG9E8Vrsh2+8WntVrT6lNEcsxAIfhriKtilVs
O2VelidxqAak0hmnkmPH9FyDDNMpb+fwcB5i88l1ogAbEylBkfEaM546sFgNMnoP
AztjVGjNzC7wsOKiX/lQ/G86Ka+UlLI0lInLpV1090FKhDuWLb0F8u0nmSTrS7BQ
kpc4c/EQAlabJhMGo70yE9S7RJ/vDJwHR0EBLPqaIUNzEafKVgYiHdV95SoJ9f3T
y7vySFOPPyC3JAG4BuOVxueGerGHQnv5jKaHYqoaXkPHyX0u/641GB92um6J7uTe
Jm7Tb/FwPEzARwYV6dc2P2ugGyXLoSGkIZcYYlctUjFxfe/0EmtdULJQkQViN8Ph
4OnBjW2Vu59WY5+WFLaKjHZSFc456n2LRTT5N+12jjbxMxb/Qr8H095GXSuFWRi4
Q1x2qTulhII6bUIJCKAfViR2X5lUR471XcmaF5CPnnAdTwMrIpDgINSwVaZsP4SA
lVBXlflcJHHscD1kk7Ntg42yctiubbHeCwT2c98BtOd+zkEVs/k9Y1dWnZSY297g
TEAqGtwduf42StBjAnpda2M7pSsRJZ5wHkD/DKysEXvuY+c2FKfU9/D4RAkbe0xd
JyOkc3QX7xEg7/783ST8JHd/i/XSKDqTrQhHDWYQbILqdxVg3DOGkc36xjqPqJib
xYeMx+PVu2vHB99Qbbt1Ykta52qodk76mH8in4ieuO8oXfm3huakYz8jX5p4e/j6
yI0Q83P082fBCC/20O0WL60siShOTJubKK4F0BpWqnGVlINwYJgg4LFeMHIrH9Yb
mfFVRdjjg2Dbin4ggjG66Q22m8KJ60d9oO2HuAmOd4wa3GHGXxOwjei+TwL1f4DH
Og66s/OoA3PrbCpdBlSn1s/+0gtChKjzBvoUZIuxpqXTxLbqfKAT3Fk/jT+Q39zF
JFFALXFiViubj14u/FJyj4EterUwJ7o+XyjraiOKCE7+fhKPx3/6mdd3PC22LHF0
5eXgD0aCF5EDAeANcg6CpZpveFo8PwMp2pQTMcGi21IJD4Ek7TiFZO/N9kHT4Jf4
8a6A/XUTGIsTKwDliQ0zHV3sL1AmvICHs99pdiFJ467fDVkLxaahlTnkFHKWwS5q
NvHG/bL9pB3qzz28MqomVB3QFh7xrXFGUptmbogpgKtH6GN70YrWqKLWyi6NDdOB
jtdjGb7EyB+qVobC25n3Y7WnX5AOwIijh9FYqpHVg/g2OiCwsNSmo2x4xopsssiD
5MU1vH4RZqbAH3Xo1P5kDfBfnzGA+NzG4trHkjwMyUrKxYiSQ80qOaoMxZXXBA96
JfA9U4CvCHI3edo5LIlngZNpnH6ZKUGMxSkVHv8/zFjxEqjMV5NgFSIn/M76HOdN
SX0ESNkGFx0U5YOy0WD8XsWTqBPIJ1GoDImzrb2WUuklbzzuVZRns4aJ4xJqmQyN
Kl8bE9Be4LD/3WeMf0AvIWUf/gen8lOkmEeXBGMGYC/AO5ccwizXTtMKP3qOleUM
7NR7/WFTFV4OiBbNvUrwL3pMqGU7ziNg+L6HfY2fnXJvw44xGRAEyw6TuudUEHEf
to6tOLAjmEN87mslMEDJUsXjTo2SOKCYfWCBnaEbCnpqLHIJBx7pJ5lRPCMZHPOP
vN2I9PG6Jw+L+60pK3mAZQflUbApL5Lg2E8NExerSbYhwqTLV5OIPzMivuMRxUO7
0q66Pw8by2w6A/ibZArr+CDejqTrVKQQDcqpOrLmIfOwETQQeY6ZaOeEDzys6NQB
DisJQPyM83rbRgYv+XFBcZQ2JzT7ImpgdZdu+6Y1HzpVlfzSTdfxT0DwOER7Z1H2
I3ZL2BCEH6CEk3mAVF8tjqJ9BCyXurK3vulujL7ZZCPrbribdO+haxg8VSvmRL6P
S/guGFcPZu1pOGrMwlKMANJKwLvDs10WPiJpw2DY6Hu1W84npte9iVb0P6fEESaE
I9+KEa01PuC7st081Qltw1PEI8VGJsZEJsynyw3aP/Gdf+XFKiApaJcgsR0a+Uuv
CFRLK4aC4Ubcb0nIUkrpWu2q75Gn0CyXwBWUqlIxfFR/8EJ8JBF3Yg/oB+hMUQOK
4DR/ZXbkME85idEHjH9y7TuS20xdUriKIiweHU0UywBFDPs/Qsfo3fCy+14+NO2T
c3/FXq1vjbiQi2OFHiJxPzKFOZf2ouBA+YIg6tEgvphiYiKrcDahwrX+ggR/qdEi
u7d3JK5Y9jOYrbVstssOYsOk216DUTzNzc5FQth4nlEN3wLjmthI2fUDUpwWQo/y
0AUzlGJMeACb7XtD7/h29jFLwxJSy4pXVv0987bd/rTqkPntwvZORxLz6Y3TgJAh
yn7sKWnl9jjU5w5F9jhlxjjqKyr4lS4Wtpr+qUDwpVGO11ZXexjZWk4iBtTDC/zv
IKfWDsI/TRVA+NOxGBumsgzbomEr5X505YFHgvSrvSrnwKS2vKWr2LbFZ8C31F6z
ewhWDfrJUjpWwe8YKIhzf5euqk9kbHn13UaPns5IbRjBkjhQ2bWdz42eRBerXmT+
4gm7uvcvchn6Fs5ub06rXyAjOY9QUsBS/fX79nL2T6rODJyngySpCLKv7wsEYOUe
0BbJ2Ih/06N6UN60ao9UDUv4XY16Av76urphSgMP4exFxfla+6TiVVWuq6Lg+Fx2
mjC+ZMsDolcXiPErinpkHaYIuWfp+Ef8QHHtmvzpmMl4PsnDba5c9vnNf9GWMwFZ
E0TDcfdgXGjmmTMbTUJcQklh+93RSA5b0RsNrZVa2helzU1aDguKK19gLr2WLUNp
HYOvfXq+kAHcVYGtmp28EAJA7WU9IBfTzj2QT/NPNsi91fIshWWmsyl8K/ExU7E9
lmfb8iH9ZMoH/sFjB7b2yCKSiAldwsj/soAxWRhw50ZYqDMW02pyxWGGLxv0Viwu
pyJOFgu9aTHiOVFgpyiZswJ4+P8u1auKtZMJ+z0kxD8N+Au130qpI03bOjoqWZXL
Hh2ZY5hL9z/HOlIhmxFd5kyi31h9tAqDWfeL3tYcChaNe/akOa5iGe0PoEzXV71s
4y8qE7132k4zIjDjnrb3avdM95cjnm0D6cd+b8CeHfxekLV5Op66kGPHuiwoitn7
vTRDRnZgIe3T6sp12hKEZyNfwvlTOVCepSw3ypM7tOrlEF+JS7bHVdpMgeuO02Lt
lQDHLErokc772/hwXsoa0gaBpgTwHBCTzqRLFXlFhaZS4JMKBn5Maa0nfarLj4Bz
Z7q45KiVcGOEXKEQIAQ1g5Q7fbp9teiGal3cQwJYTAiW00ZWAnDDmmXxRJe5bpRQ
4xf4ajblGohSOQENQK6sCj6tjONLWrkjn7Rj5gg4HrJy9baftCsffpGQEvtk/JF3
9sQByMVQTKALHHLf14YNeCgDdEDLVtaPfgFm6QBlesh6m9ttlY8eM7/NkLjuWivT
FH+uKIvfsNib09o8jiI1eJyVPW1uu5wr1U2ViwtHT+YwrrXjEgwUqOGFCQ71Vm3d
2U8ERgSXaj7MEaT4UydQpHoUuVOcE7oigpqWOKqMHtEuSDr0+xV/xk8IR/BS9vCv
gePdCWNH8byeS5aR63Xp/GTuMl8SInJoZ0nqZk5JGm35BUVdiikUar+zPOLNMHXd
92jha7q0iC7cab/AisAu8y0hlGHWAF1otamSR8lzfdQhfxCX3oaw3T8J672A96E8
2w1OYGtJeyY3YRZPc5hK4xI8kH2lOrRpSA3Kchv2kcftG+TxyDtpbLOYvCb8nU4A
wSNYbeZqtE0YmN5eKghnaKAvKcnWzQXsv163asiiYn+u2fxuxbtOBJSAaytSU/WB
QkRYMM/pAZi0Zgefd4OED3ZcMmauQRtaxvvZSy1+dSe5xZSuofuY7kKO1z9AHdmF
s24Kb3/YypYdAFY3pOUGNxUMEkVHpEJTrbbxcjWvqWSNpQ1segAsZ/DXW89BumAB
yJgIzvTIE0PcBQg+Eh/JxPvvDkoigWr5DfMbq+Z8yd4pWO9OhAu8/0TbOBfjdIxh
pJu2g0SEJ6er5pxefwNjSVaZkpqAKEu4rfuWs37gnkKIFnqu0cABZ6WKDqTpNmsA
lU++sGGIt+Z3tV1E6gbkPSPJAr5djoQ14Bi37GGYiCL7hDMYVdngzMw83NNNy+xr
deljhqbxPVX3Ty6na2qFu00kj0/XtdB34n38eDGvNE9CVFF7aeOx8jh1U+3GCF7A
+8L+OdBKk1znp80e386XKE4HBiF3TXtPv2lC2gKB1xch5RXqG7a5lcQlSW4FmGzD
errAlOq8dFWveeBLv5LMK74Mre7vqBwfUxSSnc5xMVsjmrkvqr7q/Rmx2NApqZcq
LcL4KxxfWI58rcsijASygPlWv87h/vpSsfwcyPiy2785/70zCwgjs6ZEffd9K8l3
ydQZgCM78janA2UkR9N1eiXmSWmMVxTuWpDgt1Dun9Chd4gA5qqafm+B2/pHKHDk
4ClC6v5FHoSmxFIfo1tNNeMDhjw5Mclwt7KOg+VfHcUj9WbTlFe2CXy5tY/7Kcvy
1xNGir81bWA5MjPtoEfzIChimBlOmPUT45DBMN35rmwxWvM3GfL4Ml8+l43dLhbh
EZhuKtJCxY/cH6yKwGynl7IbXMlV94N+JxvF3/RHn7OGyzj3KpJ7cDKgREWaEpFJ
xQP+lkIvd1/e3/TY9JrnTEPRwIU7T0TEPVRE9ykNI35+y8JUIpLn5RLDcvsURyRg
WIGdNw3VxPpUHaC3FwBQ8cs8BIT2Bh67ZUmnHBvWBrSuD1mF3Ghb45I3moStFiqR
7lKmutil4h0cBUIYFokQMNvF0rNaF91Vy1EQ7LvM/XOy/JGckeFQAl3nd2U6ho7U
UJK47owcokTqHtFapteyZx8w3nIeSl/b3FVFP34FmLOVZ0Ql6EyzDpPOG7hYZln4
vzA3MbqKLe3KqtLVIfiEmowE92Ag8l4+EUcd0oGirFiilAD+LVXc1ZnBGtCTF9ZU
3wT2RWxTNiDZeCoXBPxUA4T9D8qvY+8uNIkvzjibLuuYcs+nc+BSW1vr7N8A28WG
ZwtJRmUz5qeqLXf77KDKLlOwnj3HejaJgz+z/Qc3uaoIEl+YA8tYFCTJ8nPUKbbT
QV055PoqMjzTFInQL8/FroxEK+nu1T2NetJwmeZoBDckdn+O9R4XKBV6D4WF5ZBU
/LvhOqwzMLvUAEy141GLqbSpySOB1cXeV8Tw7/1wMgCmPHei+GiIIJBb2OGU1/NS
pmZ+j4y1olTFqv4qwz2cEQwSAWDVcPgyPujuzbWpGbttLhAyv83YHzL6jVJbvzRS
3SRoUIxaag3win9SK38P151nSZr8MIL+an7xBgQebQ+2Janhr/yM3sMqrKxMIwxP
VUjr1JvWxbcRNfcfGykYnJMKmEaCftTDiLjTjR6xTDM6ovRbYoFWKprYjzn/XHSC
mhs8y3p/T1e/b/1WJnTBq6NO6BVKQokRCq2UW4/seVxQBJpHzIISTMpvxzse5imr
aKNmwIzSWUrTUgR6eHhzuTVRBmqaQD7hliOxCArBljNN0Pg9DVlWmVIbVcYRXnhP
pEpFN8HbLmTrdqldWRzKLkYpPLS05EsUgPDfhyQdo0TE19exWX7kpRfIOmcftgRU
PEny2Y6tCWfdoaWHiYq7RF1rffmlUjVCpfI7kL9TbJfudQHCEl8SCZGRnWQrIAHW
d2GBOHT86rv+TcjLaIGfXjmqWDmBBOzMNugWp0xjtbyiv2lxrNNZ5DfzZFut6pH8
BBIARCG1Hx7P34x1V4J0RQTtADfkkOLQB5TDP3j+bBu2gdHF4ARDv3X1gKhDMobv
33FJ5PRUY3/fdSGYOS4zK0DEL4JVUCatm31tXna7IQ1qeKb238D2H3jt1qVSd0yI
C2yLLl/frnpd4dx1Exx4pbTrr9pKoGZnGXk5VKaLkl4XLS1gkLx3zspClkZef7L7
YmR5+POsSvSbvNYRLb2HKw1GnG8uwPQ433xR4J1XxHwtCemCB0sU0MFWL/0oqNON
iH+J1HEGbMQ5/f4yu0kBNaiIHIoU72q1IQ2zl7u1SZNDWH+5MUMb/m63nGREFkNA
9gf5YcRS0xl4xjYDFKF7M6Y5iGJJfgTcBWJqEwn45trrboKasV+IDGK5dOFE4RHZ
piFwe3DTwDj8RahUta0fdtaoX41dY2Qjb4cPtbvTzryj0s9SdlYJb8H46QlBWtaR
fzAyGJenaORSFolDN1hZ24Er5t9ZBX5FeDQKN+laO8Az6ChvgqVEpRuKBSz9EDNF
vyNdI1FmKWka75W3Tc+mVt3PmAGA82eQF/t0hwTzN3KVodxq+Rx/DX3zXSWcsIuj
taUqDSS2oZqEQ679FAM34vBhnoDfh/bTnR2inEH+i/UKptZRHSNr6PHmrefX+QQw
aagDaQkSaUFihDxvEHduaXo+hcxSbyAKoBPJqEevYCbNcs2cIDLJMoAJCxEsQPtd
sISs9YWPSG28dZuvVZ8EA6VwZ9CPMn2kkzI/R9rvCEyrYllX5+yE1Dulg/ejJssj
i/BP+U2NlUZF61BbA4Xiz9TnV2bJbXdSzDmC0KiuRKin4OxCEegAHpxkGOyKEha5
jdQPIQ80UVdGtiBU2g3/XSxOxV/dPdRDuhenLfw+4AyImgCa1gRQI1mlHPmIAdA4
kt/hPHrx4IEWwslfq7im4f/GKMsAFFpDkzeTdrkAmrTSIAjvF0FdTyhaEiql2D+D
Ft4owQfQO3WSGouijGJGK/LwCX6YQVFcbYgrjGWTind3H4o5PDituL+S01nJD8xY
Mkn4NWkuTb8npqQ79Sxwl6Cmpynw51fSnDTQJkC0oPwMLxUe+n5CFrOSMLqlaOLq
02McEK2NHVuEDdeluaf2XBYJtVHJHzrUyvGaLSnRwhITixmvze9N7opfbr9U2UDX
BgsHpEi5IshfYMVIyx3axNE+3DAoxGWYQF8reEjo868A01ofIQRQJSjjPw6+ZJsK
3BUL7W89/iUayMz4RoCCfuv1nZbUXrknF5j+JZE/ch2cufr32Rvz4yyoWXUMhrbj
3QK7DmNKGJP8nJSVl/QKXeGDl5hgnaZK3FvZvxSTqFhuJWfzp+DlpdgZO0EKW00l
pJra8GpjsQCPGlnYLQvbWxdbeFukWXJXCO7c3zwY69y5u8NYG6u46b+TNWPzPTmz
DFx0xOatpDM+k6Pd/JApMgMeQPvAdCTSwayQDD+rd71Vi+IOiknmYB+Qppi3Nako
H/v4nPUYn0qqLAMwNgPBzhvuBfJvZMnCDsXIoRyHQ2LIA0oPSXV9EAzahr8btJh8
mnRcdh1vEy60wA4c9htOo/Rz+9wK77Admq5UxbGjt7kMMR7LcJ07SUTVVMebmAE9
01ira6DqDyERwpxHgZqyLmURvKy73IKHRtHQutEKm3rT7g6FhKUyrhVWt8gcASaN
4UHPQlkLbVE3qHv1Qrt8ppL5Udhs9jswC9048JHmDiu4HXZkVFNmGX1TkOe5iLO4
39zMJ4oW73+UWMG4OxvCEV0gqx32J3Kja5R+PrW4llHwldYonEKs/WYLnpD+q8/K
bitLVMbNHRMl+q5PNl804dF6kz+7juxKCpWL9uMwU8prWq6nAK05ZMkBixzvzpFc
iMP/E0+XbpKshDP4GTNzKzJmd2uh7sGmPjWRywbpyh+TWIT0D9uNcQI4UvtIz1Vn
xtUgjWP0+J6nE7llgzb5G/rylcoum3d4fMRI33XZFmoA1Vfl7jP7W2Qn5P24TlUZ
k1b5+U984R3KuB6Ol3K2ANCq4bnR0e52YaD3OvjHJWuxtgnhEMfAp5AFv909sLWb
ZUMaXQdbCg66UP+XGJzZFoP9jFM/gfq5Yk8F1JfwmQrpMe4tz4QyBkv0rwyEwUg6
5fN6R2VHYwjNry9a4XK3DFAiZakokrGnuPh6PNi8RH4v8vBTTJ1BTCGK/Rq7m3vr
FoFCE6ipHe7V1bSn00e7pvM1N1sMjOE8pRm0Spny0DHl9Ie7xQISF1HUgVwBofw7
hG/LqflpMYBmPbebFZ4YS8nX72QDeXKRoGolWL+gICgobK6Y1kr0LWb0lYUBiMwH
klaKPdkpFuPGRL3i81HrlKbs760og5gjP20L+NW+o50N7NFPN1LbOkNFYbLNBRwn
QujFUZOjhXRw1MLcMWF1EeTnJ7bQoBj8KKxafLa3alwbluJwbZ7p0AtU9kcqRRxp
oHw36B0sTA5qgYL2GglabVlaDpNYZTZiivbbcm7vSb9VnmlShbvM+xTeCKI5B81E
GS9TKduNXGxuwbYOHFkP30uJa7VU3zZDg+cZUoQkVgfL605GLPgq76bU3pxkUkRb
jsT/oKNYhHgWv5vQiwFp206VTIwwa18RIdJBuQ+HthuODwvV/n190c78Nm5JTgGE
FezTBYvaHeSXxKx14Wkx8sqG/qzDrikCuU4cgUY3KSWeyaBysUc5fZ8QR2uKY7W8
m8OjNBTDL2hyY+EHkAD2IT+SGWQb3py3Wz664RWyIP4WuIVu+7Efcf6OeRRS3gMn
5FDOWjaENZd8y0od/aRrD2Lf5+r2ieuXCY/Dq6Yo+lmWnHcKRDdGV8pjE7Am3HX8
BLAYVFQHnlHa/qWVqRsN7jvgmULq34HJ2T5jn7RCCiVjIEUd3QiSnrA8T0yQ+l/j
KWajOFgL1c9TDxveSkT0JpgSsVN7/cdJPQvAsmZVcnmUnD3iUARUIgiMqsiIs2ac
SwF+nnq7aEeBNEo01aO4rZyOMBI9yclVLsW6aezxQhxCPXrdEajN/yEdGgbse96C
D2ydY1AyBva50fT1gUCTSdSk71GrRKxoRNZihxO7Elc/jNTsNuWE5HRQw1ZQr4UY
2SDXc5gXniHl7KasisxR3DnF4udUvkC0awd2NJhIQxP6ee9DiGbRwIMWqJRQRXMd
LHjm9qmZlg7r5d2xFRqJOAoV41u/ZnLpYbHgpdH77Bde8872aO6qqhSr5p+eijQh
GTnqCjoA6ccqiPu2g5tUHJyeIrQauKmzqGMWvz2B2/qB22ffctxLkH69CBY0JZxX
tUxCcP+PnThJURALZoVyM6/lqk7NysUylZLbeErYNGxkwAeQ/EprEMfXdXDIcHqc
Ju5EZidqWaZpqelpYt4ZspbpZwiB8XhQbzf5ctZyjDY44WKczB8SI44WGgdGIksM
MBCa85QgE0pUGjBsLmK56pcKRV52NcXZLF7lBOv3j9Yj/2LBUcvvPiT2AVRnVPxq
r8HnHZuGXVZNSA/DSre+6hc93+uJXdTxPGgWML2hJzZKbQ+TiQTdu6t/5Tz6cG5h
5QYBGW6EesV7HH4AWnhOsQWrAfM1u0L5ZnU1OJRneO29pJZOvF3xuosgK5spfukI
CQn6+0kjx83w4bFA8djpgc3hTSKfyvHmnHhBwUpy9YoeetzhGo/1uUTA5MBMOeWt
89mZQdsbPF+9G/gAURSQu7zOt46yxSIbM9laClC7phiiI6GNiaqAxoeFzvB74Yz8
OhGBRtLw0WhvF/EZWF4S6y2v9xqeJTStZ+MDHWNbMdyXpRzMtgRLAnKxjNvvpJ13
PawMlOrKgyk0KXrH+oNqUV5+0t/2C5rjrpiBGGjbMTiXGwiDmsWVkKr0BSYsMJWX
Sq5/0P2mmRBUPZ0cNH48DeWS4WAnD77OSwCy3B9m0LnYOPECGzveGarTnpGIWtXx
pw1c34vmVdiQ7F+AyFwxdHwqNarb+e6/94hvqFO/zSNAqFSV4UciigFlARv1oEF6
JRc8+T3fJWlJEJOiqt0wmcJBgkJh2If3fIVhcd+ab3YAVWEWQVOf7Dt0t75ilVD4
lMim8UZrJ6JfpU31U6Plcluq+6f0hzKR1pUr4ScdsQbtQdyBxdqMI4OIYJuAqWzU
Z2JDKNEW3L7m2nPfxaHh7W+hCiq9kvIqRleEjjEwhrtT9B9Zuu6AmAMkCQsbgA6H
hAxmHvfn/FRVgfM6ld50Wkc/KRy2t4K0ZkN6ivFYmnO6NM0oyouZIXJ36VDLgmEp
PCoOy3ttQEeY8iJeiRqngEWU12V0anGE4YHmaDprRas8qxx8DtZyIFEzoBiLxm/8
s6pl9cEcO2WfNto2RztShQ8YW76y3nYExbC/lx6PbAUzwQC1wBPYU9asmRZEjz0r
LOngtWBAgtip22IotEW87ooahH0eu+cqr3xtyudFwz4/u3blGPI5nMjEvXeZVIU2
EGtsqM2mRp5aslTZxjKSdXrUgv2V1vhHoE+aOKyK3An3Dl0pom76rQzqCbA1Eu5x
zw9gosSxvWKceNx5sCG8X2DwAJUsOYZxCllOP9Rn4FaJN0RwPU2Qj1MR1JGwWBub
7DHBJ+cbdSvQVrZ2egI29mwaDlkmNqgvyLvMBeUyCq7wruKphKiOM/ku7xBc7X3h
P5GxGqllEQLVNjiRkcLwG7bCb/1boa5QhisuGWXX3+WQK6kJtshIskPqfjOdKh0K
5x2eQzc1lw+sFkGCho4iu0BvYlTdDnT6vMexqdkkoiZyKQ3fdvkOv0IGIptLVbea
THEzfilRY4GptQC3P28OzeVDEgU/S92nZbQfQBZ8vIm8tYKwGhqXE17QaZo2322I
9JOHtwX2RaEbpTAZXC5pfo0Tg1dMVVu79wr7Sm4eYAaC5iLB5lLvz8R1/tQK2H72
hSOcOeebqkrQSHpmx4km6qa5OcIIqFatW6z4lO/OUPucqyHchgdHS7suYHfAE2pJ
DSNu4W24TpTwJm7ZuQiQIhf5lgEsb9FCZxQlPamlgujnfwuVn2oEhFIXa9BgmkdP
1L90k758obwBveE2EHmsXlO0QzZF0E6dvqI7CqKsjgelOzfKF043ywUQAcfgUfso
Nfx5mgKanoKwWjUwJT+kqWjw1vEn+umatV+dnTdYQxK0/xj16SJmn7R42wkaKReX
HsrA3wvQuYdOZOWMSEF3JDJMFA/FxvxD5xO6P2uwnuCMNB4gyg1bD0MbJnKS61NR
sNHvOTirtXKkhBueaEa7JNE2X03MUlfC79YwAGMiKReRKnHTQM2HNFDYTeH/ApbV
/C+r01GwEdqCyD/IrYd78xnSQdu2aQ1x63SJy+KPTBkoMWcjmFNOjy2/MniedeJ4
MKsEAS0uBJoRv+g0o6TVXf2IuZ2rbehPqhZqxvk1IMhZzuq1+ZCzNOvU3hS1G0nK
qR5iWVmetrpcUgTrSn5XifBDge+k4Ys5xqjIdExZBtxaM/heZOundPMR8oC67/UA
6i7eLe9hKYSVtndozihzQ20wVecw92XzscAoHKVSaYdw2z3NGUuS3b8cS1q4r76R
Z6TTwNxUfAibwLnEv+5QAs1PFXyK0IiIBEQLTw0RIgZeDfiUw0Uqc/vC2A1+buuM
GM/nSWHmbugMwKtCU3scP4wAwP4Bvgo4H/297GlyTDon9W9VesRWEhfGJqiFxp7E
cCKbU/wGhwdHiHL5zSvQl+mEJBZ6ewu7q5ZJ9LFQpiynO0cRG5yIf8TlR/zMB53+
gyXJY5SLRjhNjPXbQO3TqmSv91uhmeN3d+9japERcWDeQ/Po1jjZWBrp91sZp+Qt
8Og8RabJdSKsqO1kjLCrpCv+V3kgQY97L45DtBuBtlNcFwwonw7Q5lwKSOYnvWge
s/x8LGlbERWqmdek9WZ5P3MNsCULroh31O/ADV4mS46N/IJ4L0XfA/PH551S4dTP
ubFHE5NSMuNb3c6KYHgGqN5ftS74uQ7se4SpCvt2rSk046i7+/6kO6K6ZWr/6dBJ
OvI7al9fTRp43ivXQv2QuZ1iKCYlnXxUkRVsb8Xdwhp+ax/vIJkuPtYkTmGug1rY
oNp84gGk7uzBBPUehJt0MwW4PvuZvov53CatTVJeX5/3y96JIby6jFC2JMzX5fGC
cbdgD9TjvQkMIAcYfYA2hZY+xS2kgdgugqM+YzOkwi7agwbnZuzbmR+Jep0bjLSZ
9sen1zC0Oxe2S3i+N7u0IZxjuBoJRG9f2Nfcy1uKe0nQtNpBk3DjBi7iSM1eMdtO
Z8Z36ZlT+83XFmf5sptmU38loeZoiKk0T3htR2E0/Vw9wmbpkLGKwRD30AdoVBGR
kJ/9F2yyocu+o4dute/sczPikmGSm7MAJHEjxpkAPvvMOEgiEZl+XrkTlFlseUXN
/8wQi0SJRNTDBPt7ot933qLxnTezhd2V+3xD/Mc38bdF/ECn9yu9I/lq/nZNY7kv
ix++95WS6k20O71GW8KcK5D7cE5ggsSBgskd7g50GoLNhqPJYeJYo3qIqN3mKDH8
2Wspzv2Z2c8pwIpP+XYmS40HYjWlJLu5QbX6tDEWnVlJ/6DC0C6u5mvdzhDepL8F
/gKrfx6Kb3wcPlki6m6G2pOGN8mVRRrJ4ZWKYDFcGZ60jjIozQOqOrXYNsXjRe22
F+oIbLzM3UnPJCIRi9HydbiYFUkDjTrxpprzyKBxXHBPAL43F2+6PbU+aPI2pbAU
yV6MRkwcDxkSkgQ50Q54nryDUuA7GbncCJS63qVb5FYwjMqLAcxjEBRkVOg2wGUs
gFhHJWQt4sphJexAiEPRTGKudF523GlxSJJ5ln7MICJV8zdI6x1yATDEILzO2SHi
Tq8rOoAtKFUYvEW4d36mKwNr9xBXcEXTxoqMC+lK7PwXuPaks25cXfqS78XvFUyA
NbaFykeMXmx06vGrdbQFHyxz/Iftd5sFy/R8DzdRzF0F7Y2ybLcJUWQSH17Rr9NJ
fkZ0KqowmAXe2gL54LdCBtnTAOQ7lL81M3vsB/iP9odZy2cnhaCkg76QdT63VD87
gfnag7va9w+P7EAKUi2owPKwW7g+2x2BnUktX7jy/JYLL+gigD6uSRIVS2Qu0bjU
prAJV6MQDJiJXamuqTHRAb4sHKsJhK1Vm1nBC58mOZJoDDB/kmBTq7skDwg2WYIN
iKmvft5L9E1D3y02EgG7e2FZ7p7yOwgrn2nL8VqdDNYDc1LNDvA4NGR6JJs7I0Zs
/XynyYEJpzc82V65VEx/8YVCmQ1a3wUJL19Gr9V9RhOFX09QpIqDWdfDWW8DRjyH
f9XeNqx256FTPhfrq36qRh79fnQMi9X8AN/OaBkGpCz81g2m5NSk6R+cFPRQRiLW
U3pXvNX86/KHJ55KgC6YcKU87VNBrcXmrQXP0/J6n29PeNewq3Ym7a+QG32SNMei
vWynVuXkW2wrClE2oeuO+GSI7+82sQtXB+KJe9uy9uawEdd3M9CjvKNRPmCGe4+c
2+P9/rZEpgbqM5GtkJ5xxNDoa1qLhH0YeJPmXO9C8eOPXKokFe1OUkIuGjgrVBxP
+Jm+YQwVKmZG8u+WPfvJrrkU24T5Wr5n9txD+l6gh2inxBAdCzmc+t4k8LyiEUUl
cVjQf2ieVAJFeL9cVQSF+L1bL6HKMkIE3COe4IQ4DGmCkYUP77XcJnDonw4l842i
lSgVilBYbriuDeYssE8ph1wl6V2t48qZxkTzcMAOek9T07beTRelE59Y6PvW57XQ
aAjO34nLQqzRT2mCWq9mOa2zJmbbqbJCWUtC5JWZiIb82JnWs4yqyxGOsiJ7sDKZ
puilMjwSLuYdipipwncM00T3nzAuG7xyjPfElbR2LJSXnuZXzPt5fOzOnjwNYXaH
kpUEkPPxkr7fGgE7I1E5MAirN9jnzz32i4M+jzHYI732Hg/TiZtLeVg1ZsEDjtkp
y4y7ddhhVtz1KZOXJveA4mn40kw7VE8dzukWgXbSs8+/T3FrHm214MRQPe3xuS5G
GA1I/PqOojYLgiG0o1Go0ASijv668v+rRvdnbqBgQhfKQdRoyIi8GfVZS7F3vNYy
OYdy43l7xS6S4n1Npe5RSbrf+hCx1r7QNEVFoczUBqdd4DVFkLnT6krpD1QuNyv5
Z88FciqQ6Falwia5ZQrLiyVAjTWMzDLbcBfo4IYhUyRyJeA9vrrrxhAZ49773HZc
VHWGh9odAW/GL8HqZqcUBOu4LSW3aBunPFV03sWbQ1TL6XAnRbLFwabhndH/J0K0
Y+noNp7tO+y0PG6G04BoYhDuKHSWPGQFshiievcHiLbesr+3hRELF4EHOnDX9Fw5
EPLMnF12oFP+L/8ZZabeY7VmLdtwSVV7A3DizBElSv+vKlTEoJD49NG3LSHlMkbS
SzkLF89p6i0C+GqDM7aGiE44tPcrb7+9oUYKedhkr12MQGXGe3X2sFuEyuTgUY4R
6iwZgyj8ESOMufQMi22kJDMB188rhPMPCmBiR3zrk+we5t+VnLAoAOAEpfoSJFZj
jtmeH5hO9Nlw/QNUv1Mg+IRjc6HEVhVZXiXV+ZabkfxboAKtoIvM0LpMAJGzbMlE
LvAz9EQi9LbmXRgRzXjgh0D4lALNHT5/N7udj7/ZgxeSS8JqjQYbZ7q459jvodYy
hR7wZ6MFUIdhElkX38s7XYE9B4apaDi/KoaL/vTo2qQVf6R/pJvb9nymeU5De/Sn
rggfDoiVHnbB1Rw9pF1JcUX6bFZPH4lifsikPpXAWWCFc+J8vuBx6l0ZvnlwQZQd
q21FK2JNx3C9mVJ+VpT9kpxf04bFWM/TpmFJRjarxSILZxk9o81pXNEdcsez1Z+e
nWMfKAHRI5MqPt7zARZ92we+1FRPT9AZbCTPg7YH7PMWHVMCziYVQpnDYIhMRD3g
TJ/qyrahf+t6G8TqRs9qIWTnsBPjmxI1sCIibHjqRi4S13pyu3uCGRpYqey/FNMi
jqPL2ZaIstrBA72n6wrfdIdwqmybtJtK8JumlcPafxXXYWMIambhiMvuAfYrEqZ/
9+RNvs1KbJRrrCfU9pFDAkht4vgWPg2gQuHk63pDl8LhUwldFe5pdR2MCD50C+Zj
v3gERZq60dhb7BmJc1DottJ/XhFDifavlsNZCvXJHHsXWmy6DRoI63BfIDIPY3Ns
ZYS6lP4qSLjaJjRNBzwluJni/rYVYXl6yvPoG5T7cjhQQu1pKjb0lES6P0yrj2Ic
lHyr60/8cud0hen5gzpYXBj6Wz1Cj/P4S6ozAMM6gkgkxZKCqsBIPv7YtW0Tf2Xk
0Fm2Ji4jQDZcz9Vz2b3YimfGm7jSNqhaS12kUBnqWu9w+y+b7zvRA9fyKUztTODx
NCo2wk9imR67rkSgyMpXcn2RkZs3dpWVAUdGQIiAQmL7IaoR1zbJeBna9SBjSii0
IefjLqLxioe7+Y3H8dSYxUl5tQx9B9Zzl4/176ntQlCPf69uxkSTOsM+WlTgpsuv
WNXe2C5qcR0k0pRQFs/fWDxj9LuPplmhCxTjDcDaxKlz7PXCugVSFGKX9k/oOFMS
Y251yy0a4EbCyUT0wmCu5uFdDVKyLk9NDLBMMzQj0y/t1IPPcIuHdG3em2ZErff4
RL4BQfNjOV+z7h6V0iQ7WMA0xNnZPuKv0KKNakdkcpHgB/JpV00AAAIj4kNI3K0e
9kHSwo/QWVW1p3buiwNAl6qaRH3UYchE6a+VrPwuC5Lch7hP6RI0SZ0+VFEww/gw
jK90+g3M43hoHVXdbbE3r0KjJx+xsrS/s9t9wUUT0bKZbsIQuFw8hiZqxhGBOvW+
0g2j5sJh6uL4q+50aCZYJxEZx38kLZnu1NhwE4F4/Lpv8rQEZcOTNZflQjySGBcT
k8DK4H2yKN/OFM0Ec6wMdCT9Xt5L/4FcGt+VW04EMGxkkxrhl/M5M2PhX0WMYIIR
MVdIRDOfPtLNZjWtZk0bFLcG7255B/Bv+7TifDRd0uwKNpOlkTUHmn8WK0nszlLx
h3zlFyZg5zdnvd5gr1oG6wJVv35yeckMTxhaQZ4VWg08E16gARc4DR/n6nZQNX9z
TTXU/FUIcwCZgityEHh3i2jueqGIXG9Ejn50fhX/NmQy4quOI7M1bMigHXSnwWcE
zyRX081bKnM61YdgDuytp0tBacAe/68ND742AcHmTCMoBimds3p35Z02eyx/PKr7
w/GaTlmdojoOtAgUmGIKhoeEoe/rXJy3tJVSdIqDjHcfSaAd1vxOFy+L4/FA5mVk
uXwr1USvDRrNSt41+K0WSwCacgRrcIJY1ciDlO30kOxb5YzRD8hSD8YEfeRoaG1b
4FYourO9Q9hMm9OF8RfJqxpjLJv/mOAuLU7Ztvo8nPUwMOZCp6XYBfce08HJFtFH
L4uIt+1uwRX1O2mvMrG+IkmLV+97wNEH7m76ACuBGmbgjl9RaZCE3m1gFkQQ/VXT
CHjormxsDaqBJCJS37Hkc/EcxcjY+8IaYDmR7M3V3QuWaAkO5xvdWLv87gqaNblw
i3WtprOoHRL1WQ347LJaIt5ECIP3P3wTaoOhyE+eebpfDuNVYCsCbWdm3V6adMqA
uYz4y3C+7pFH6zhvR2v8VwpL8rlU/ljiBcP9Bb9wOXSiA7qwkPLZUyXMn5q4ukig
vMgce4PiBwe+jB1jJNSGL2eNYKI2+tDH9hXVfLdB/daFlSYYhrO9BxEWU5EQtM1P
PaQr1NfYMl7WVHIVYyQXq27Tb3RTUOafg0bLblKewc8sFtvqaK+RaEm4XiVqr96r
iAOEUuqTK1SAlTuPQSwF3FzpVc0UfkUZqXyDFOiKgzhqoc2/mPbgU1RJFKiD2duB
0t0ny8dm0KOlyQxA+6s8vW9Fc83K4UcuDopowKvJz3CJesQCSnoZq6TjBznSxojJ
5Yt85bH+PGCOGifDBVANR+EIXWSlroFdajUNjcj+xvkCLjI5TlVnYvpgxCacKdaE
Fst9JrMOHlaRmMXvOhwKDrzOetNs2IbBqw9hdnRdSau+o/rGnA8PfhFeC54hsJso
y27SQMrVqupBzCeYCOknHQPvzyzpLDwnRIh83Geut2SzyagIyabsNuzIfJTD/WMF
XWlliU0oFAyFdF6fi1xG/Ipr7wIOkqsGXltO9qbVZM3TApt7KuIs8ZjxOgAEffpL
dGS6PzJDpplYQcsY0r3mNAUS9uudTWQJ1BNAqC1IHhvRxkdjhac0OVu8DH6dzQmL
IhrGI0ZZ0CTBpIB98f091ycGMhgY3rO7MnOPLvXS63+so3KwBzBfDB4jd++auaOs
0yChuN0OWvnx+GYBbUKP2lOX4gZrtd7519+U7QJKJWtAuKNyhp6xNELrYP7L3GhP
gaZVQjQhlRNiiYHMTjNq7TuzVsGF8ojGoeXljvRLSZ3pPZh9GSole/v2Qvl/zRdV
tClX8yeeZUfoBNTEd0CWVbY7EEKl3g7ZrtG2YZWSHkOAJOTL4L7LdQ86pIMo2jfJ
/Od/AheHLvI023dgmiUshHZ4VGBWUV1K/TB8GymmfWPWlvNcYlhkflFSI0+SpG4O
0abLyYChNp+2XUYMbVPNornzZOnP6ZxqHd7jUGqL7imjoeFwMV2Uqxt/ycdw9mco
oMJLp9BFviwGheMd9LhevBJyHkFDdb01nzNWvbFt1sM8Kfa9awGb01JOPncBowXR
l1NXRKmvN2X7zkPdiPIW0fDfvPZgWQveAV8Xpf/8Lls5HrrkXebrBxTrm20v/34D
gjycA9SZ0zznbKFgPRKFnyr/CIjT6j1fmXX4qMwZW1eIawZQkkkFWOlCLBGsATC/
ly6m73Apz/KDdeJ90sbOfbCaivSLScku1IXW4fStuyYC8AkKip4Ua/sshcKQrbid
pTpkgUIQ3f5DUAQryC9gqXoeplm0MLwdTabEmMcArmPKpxwGdYGYmG6FUzInXVGH
A4VrhmWicsUkNA8ZMmwP35ZkrRN/ejZt92h0C6Da/8Vb4dTqYay5OudK1cq9+TTl
4x3qYAfAKmSskSiyOZQx4oFr/WJJaW3tXbeIK5zsdjz5K87KGsue8QyA7HK7dbvF
qEcg5yBzNpt+ewuc3+0qoj1X7M/WrVLQBMOi1lWNmPgS4Mt2vAJN/f0b/obFHfT+
owGDVpWJcdFTnZXQRBT/ylwi0DS9LZ5S5VMKz4rX5VsWJbIBlIGFevc4anwyoAbE
efS6C2m5V9kCyIbceb3kM2MXc8Pjoi7lP8ZBFZpsU/XS5pQn+sCNZnDJF4m5bdiM
ukQb5sNopebk8Eb01d0LJsX6trRa90UApFyloQ22h8Y07FrAhIRoWI0wdSNtzyQc
hs1OPmrqH3UGfXvYYvq2MoQNzg0+r4Qyjqt97WNPhLH8NGbn3f9PKiVf4ty5daDB
o25ZOQlyeIMf4kFxVbwVCEcvT8huRnycx60cfTstCDveI6gqdkZelvg/JHZkS/hw
Zvg8mFGicqgvQhcW8chdJvtXvma0Khcd/RhrB0GQTy0PIWf3S5C+UgVdy5gF9TDN
6KDjrGe6MJwgPnvaAtHsVTj5t062hy+5UV0sPpXvIO/mmEFkXd0xRaz4WkKZzAq2
ee4+PA76uZZYISBZ5/WTnSjwX+pFSiRtpOOtceFI8m8aQ1N5OM5a+idpeq5ZUFVb
yW8VHmfyJL1TYkzKGaKMHgeOC5rFExHnK0FIhagsiCmkX1FltUjnLH71jCMOLPtb
tsqXBngBW3f/PmO5fPMAsoZU9tP+xA+RtHiVzYZunlSfh97U/nv8KpF3a5ZSC9j3
q8f3JGgPH3P5p4X3vQTcOb5aCzcgaeOfOXu32MSHIYGMECIRdzDGdEGIOSZptzxP
wOpdWnbh7s0vh5EkTnR7ZEXSGx+ZW3TehVcMLUrxe4TqPByl6mswXgbSpLSdB2FB
UbRQ6c7Y4IsLX4NaRHXIyOPgZbAatoimFzpXXmmRGz9AFhXMg13PH6dRMAvXUnvC
8L8aQ0m+ri9R3x0l4kZM0GlIFsM11GzzG9QO9CpQvVlTUSP7epQsM9dPIQ0WR8I4
udJjIq2GrjnypGQi1EHsQD+CWBhBhDVkUR1DfmSXfhYh2sH/8HZo0R/l2yZ+X30D
mar8yjrgNYVb701GV8LWHo/119MyPkr1ZGNasAvjF38jgWxAHPbbksaqezLkFnlY
Ef+QzLXljRvTKefqy3juMDdrTp1zcNopMeqIxbVqELBrhxh+8pWclX/CsrUqbkzc
dP9I5PVxtv/SzLC6GOlQBXC7qPrS/x9fYDvEtsSJ5SdirT/ndbbfTufH9D2XZjWH
5a8pv7ZSx5YYzcmlpERBEtEVAM23TXrSlN7b11iOh6fV8+mgP14M7hOfD8pB+APb
8MByA6a6BSpMGnHb7/THFw3GixKofz5PxPfY2/lSEBCDHb84la9OFdkdKZ5JuzBj
tthWHUN1lp0g6m4g0r3zWlUrk+406ATHbdtKjRe+CT65gMr8j7Fp4kiCU3uZynJr
k0dMz+pUiDPztwRYOklyBDKG63UG6CT35U780yVvaKjfRyI5q1zIpJFZe5Qy50MK
ixJzo8L5omGcsIGMGZtp9KEgCWs8PIbEliTF3H8XRcbwRNfqg8Y90psty/fHihAx
whlnNSy/aPhftCAHA3ty7gVExBTpkMGZAb1nDTlGjP52iLWwMJl/fmgwvKKhXQcO
XIOcGE+UjtI8jdYBZRiuyxxGnCEAuJ3MWl6Re8HFailXXDhhFGWmViCpxWu1OtD/
gSa68gJZsdQXZ2McKys8z4WPZreI3xAmF5rkAUSaE1GEoFQeQoz5oxl0Mlarr9Jx
+ogYQER0/bw/IdNstlkZKEm2THU5sYxBzx/xaMo+KbCG4Ow46DxSyKYILTZgIki+
kLa98EiGGv/9GVpvz5lRbcQ4qNKQoB7y1lzQTv/SGVkhzClgVnJtPVVFx0IL8ePi
GjgCTs6Y5q99w10VZhbXxe3i4PmLsYgdjTPdTY6lDOaEj7Os8CmBBnPkEE09vHlv
+o+MjnXe9FFN+pSzrNHlJd8opNlyB6crpKK8J1S6KobCyywY08LQd8L8LfEJ8NqG
iPEVxC/vPbxSGHMY/czO/LNozEkluSQh3zMCsWDN2vIwQ7sovb/CxzSn+PujrAjb
mEdx+Ivj/NctMla/CPDR15B02OJFsSt899YhWHPrHkqdYpM+RiPHiuc8eP7RIq/z
12lyQEPaNrOqYf59RoLDMuftQQRRlPcWjMVmtWmWpKE+sFwS/ct0EPpWbMe+nTPM
2BROcQM2o9y7JHyB6MjQ7hTPLrGwz/xX0lXTf5MW6HNJLaojRxdiw59kMSi6pMw6
XiWAUb7XT99eRqSg0K+cK27jsxJxN5Ak1+dg6aF3QSpjfoJWSAHvn+vRB2P1D8Bu
kavlvbWhir/3BIvHuQK7tVge6bWElz4IcdeXJ0Z7N2uEBYlg3Yx3sVTZi05zuV5J
+iUAIUyszQCVKpUhP4900FPbosXdQfXiDtkoGuljXj8XOso1IChcdp9sJER1RQm5
416pTY0XPYH/lEDH9QI/e2iuSn0GowwYf9fJuqWga4Q+eNLYdyV05OhK0j0xbbcB
+splMBfKyJUL2vYyFRZGdYwjzUJBRKatiWH+o2F0cXAUPQuiAzTh4Zc3Vgpw+s7a
WL92S4TuOXOv18fPepA43CVTswfW+TAmXJETEayXiQ28lqut6pLMs5JQbAjaaTFQ
aP/zMUBhe6YBTgrkzZjSfLLXMKr4p9CQC85bvdauywHTugxFvexlYPrT9Ktt8JPX
Co1W2I+5MoZROY1pABOCXqwKXfr0H9LYbMihy8Ct4sSCfc5OV931L8OCoOmM4/ym
5k9AuR7NpfywHUxTqP+5Yf45p4UnGHkrs/sLY4JMlY5C6yhMqbJfm0zUOp5/wNgI
uYKjmKoZSPdauPhobA1M5MSUEpUjIk5LJtfk1k77IfZOdLGNU2TyiwnzCTSZM7iT
z3Zn2A7VrWozmqdRWX43IhDGp77Nzs0d7LgWWl2GvvCf3EUFOb+/POPP/8keNFM+
A9h10vzKnHkVXzYWgJ8T6gl6wMe1eVRP40z6lPmuJzPBdljX+dPb3Aou/4VY/FXC
V2IVCl94vh+dhKzw64BRPaS//Gp6dth0jQWo7rxcI+KSydgNNfh56DcURtafHMrv
aR1eo3wxs0snQz/4eJJVbl5sds48gcEaTKxIuIqT02moFSLrKM6xjCg/z69FZ8WK
SPiORIw6TqZLvB22bJ3S92uoLa0rfjP2K2UVCSMpMf9ACTXa92On7OY3GOfq1iY2
b0hS9MrUKRG6PMw9ZXd7198PMUs/y48BK9tBfzlzrsNx1YeSMPQVxqm6gkLLCFnY
ESkz8JF4HTurf4dUpx/dA/BXnyBjSOVutmlP0QvszdsZzOj5f/r+7gZmnDVjGmns
XVt9rhdjzsxiTtb5mWzswKyDvutXHmPYuauMAYrHhwrYIaj4yYZHyQa48U+EPGBA
mj37yWQZRZEDo+pRDEaEk1tqvsZ4kGD8XMGhNwX2OuRIB7UEwA9GnAImaPVDrOUE
yhUMMdykHJ8oINouZ7DhiwDP+OQoRFRFx/to8tx3iSZcsuADBx9NSMlsH+ROPkzQ
WiSn89YYQqpi7ZDa7PBIlazHtPOa+1ex8eem3hmWfsFDQNEqBxGhHqEbkXRc5y34
j6CgKf+ewmFY/D58uR7OWOhlLAVUr17v6bDUbJYnZz2vGbi9VMQP9G1L4CkTr4p8
ZO3joRz9h9877rhD9aiD/q4LZNRph7ExlrsTQNZvvkSbBnWBrTd4rgbfZB1CYEf1
MuJQILF/tCu0pq1L/chqBenoBn6cwWFwYhdOwdNDf4qWc8uryNw7W77lPTQuoHIB
HPBWpl3KUjA5AGf+BldEnyhr7vK7yDUgMbI0sE8kEGCRPQYeDmVygUCWM14nVxmD
SNiWeJOQjSn2vmUE47SSaVF5DvkCrQIC4FfbMO8rlWiKN+48aHubTa9FyNMUg5GL
kunhWd+laWsPmgPkZUcJVf+KGfIgizllskF+kQIhjxaEvDxfx4wejxnJBf+swLf1
L0dl7Z8vireK5ZF0a4S+Yfi8DTb7ZC9odBqEMJO+FZknv/S7k5WgPQJyM/U7xaOe
fZcrtYu6CMb2XF7RgI5bGIrj6sxho4Eg+AgzwcJ36Dq9rX57Ca8QMb0OirDQ3Znf
q8KJIa3DhcGqzKrsOn1J+X7tP6rd1ecrWaoDR2Y/5+l0PkkwgljVdHeiQG5Ay0e+
pbJF9XiIp7Cq7KaGKp+cV7rzuvbU4eixrP7muKLgx5SroizLWkCwt2nfKEIwTcM8
JWuvxOxoW9cWuaCnMy7pDXkn0HP8wW/LNWgBgjhd7+Kv5xYHaX7oEgescx7ob0UN
cYbbdTsIsBzHGtVm+umP7eDhjhbIB40X7k2TWlKqDuZXwHD0sB2oqaJZxaTNeLe1
SuXJ864ZocmIV3jxlJysQpJit+2KKlevQKPY7CyEeCR/v7ePKN/6jft9KYsDV+t7
hQoMAs4afdgE+b+m0EAqohVXSjpBaa+8Ctv+409cAXBQ0V1rlZiKzB7R0tkiAFdv
f3wKNL4+1fjD+R5Kxvieu9L3sVGUjlwmLPtuE1Rt8cWp00GdQjDhzr8L4f+aAWhq
8lAsGFlsoUMFDKTU/+mapmebDltgo/lH+KAgL52wpdNSij7gMcxaW8/2AYiKbuBq
kp5+KJdy45hUfGVbHOu+ff53yYiA4i9tKGO7BRoMxhIasrKBt7VnmbZ1W+0MQU5W
rRsJUkD0u8XKnw7LUa6pau5SrVA5QjtbeyRGQzlcgBGQHmOUezCS7/VWH0TkXCU4
tTUBtIUrGw4snJgB8ETPBLoQiHADJGCUamg0b9lKle1OFmEv4K7gzd4kI4sS/4ko
NS0pTZ79oFPMvD52/tJCLF9nhe3+VVoJ/1BLDCASJVUMi2ZACml96GrCRX29UUJE
QQlhV8t2XKL7EckKAlDh/FxYAxNAkgXtSBVzwdH5NaFAQ4ak8GXNG6Cgwx9yPQcq
cFqicKyrDRH7LJkUHA1THTBvJPgIxHRm1WFh2xG2GL1pKer3HonzD7d4xq7IezWQ
wvdmWvOfNXKBpOVz5ml6UiTneI2/12ClWxYcHvWGBp47uiyADtiR65QbnNMQR9Tb
Sv4TbVazKzCsReJ+4TSOiW5vOUyW5A/SRTpSmAKgizTVjkUYPPmA11EewQ7cCKis
fT37dYJb18wIbA/T24XOKo5tommSD5/fQKVIl+FZzH2PggRSGGfz1vS25PKJmbzE
FM+v4S4FAUhFa5unoOEx8nw6yHuyiIyvF2Yw3WKoIx5258689uz7/0OQJgarSUcb
Aw7scxp1K6NssYwv8ndlnGg3YHnhyLI5tGMmDlfbQfNtpH44w9GqTOZb5wEBTtNr
ACjV3LXCChoPJgGLA+86LlPWAeCddn8Zg0h51xMVki4EpxhxfrdQ7GqoOLLcBcYZ
/9u6QV0lOFQyxgAXUG0LrhRlo2IaMEBDi5AmniOVRaG3b9SMcG2EwR+yJt/VOiUb
XQ4n9lUY7m6qOYOVQHUTpAEex4K1JFwAAbCcRK3fEgJdqS0gJPnZcnuC0FYiqUwJ
RReYpMyrdgqkDA+3jFkEjl2U8oJVZOk23Y3EF1yZ2w7FbnxChQdqLgnqzV5Y95JP
6uOrHLMqKatTuGUaLiDneS7grAS2BfsVZYc/MQmI+Worr+uYp5Bk1NK+6kZIJu3E
lCDYJvwvWtv4SLcQAOxz58IUEWFt4tw5zyUjl0zLEZG9te8P39MmR4BMX/rTFIw7
mdb/f/M4KjvcpmdQGPZrqPfvAh5LzAdNAa79xBGJyJpWbj0rCrUJ6o3Cm2QOlJ7W
ut1P0yumdvS1rfTH6c+FJtEBm2YkPN4o7e/KuLSogeGiDYt5bwZ0nz177roJBEtH
UD9kxoUMkMn7Dp+83BDbASe36Z1NqSdbkTME01tGd5l2kSJ8xw5vo4mrOc0sQ06v
4PEc3FKsG5tTuDC5QPRxShGHR3QuIik/uNozRpuCuCD0sV+1RN5ZYHCvnEGopMfT
1q+0CHHkSgJSfjPcS4Y2sIvU+WBScnAflIhYcjitP4qxKw43BeBEgE5yowutSXMK
lncBsmYmJi8dcEW0FlYIxq25OS0PBCfODftgTYV4ETubIqAT1bLQ4kyahnaN2nCJ
B7Q+xdIpQd3v/GFm45RuLstVgKHmtVywdE71dB2qxOgDBnhsWczdbYIntlHyvTZm
1botqJlB46+MQEgCExQlllM9+N8zEgCSuz+HG0uNVan+k3H/B6Ts59OwDfj1uFLE
YhSY/DkDV+ByuRMRRLEV67mySRBZpFtdYpe6VHw5ZOJ20Ta5pJkWamcIlGNK3Elc
kHo7ppoeUrewv14KduJFkTH4ANm6AVobrOOSreFqX70EG5vQGjh4kAuudm23w5/7
QbRwfu3fXQYJyu63CRX0KzIclewYphBiLkCHpGYNZwb41giZSqJL/n3YYgA2WimO
zcytrhaATz31kXG48xsEYvl2iVx0Ckw4w9BokJyQ7qvs9TjywQzcbex0LCUrmizg
gTmdxxc3PHBQwZ0p/AlHzb8bPAca+dpWCgYduk5rrVmdDjlur5JkYbmG3+oovBHz
4O8Jwmt2x0jOQ4z+OkndetmwjCJrobaP/6rVMaSApbM+RZrOts0SH4R2lXek+f2c
qd1OFR7ZUrWFQq1a8EefOL1aDaOxfW/sAoK5K6dmiybWB4vVpBMpP5KN9QUI+Udy
nwXZMWwZXYJHioHh8WeR8tKy3Aj4I+1VvrvED4+6QEFP6nlc4jDOwSiAaXBiRTI6
tN+wzpgy5E0FswDrOYpc5UHe69g1xCCuZBJk1ajk4LOJhTiDhaIeJiM7Flirkv8i
KhIZmvG4JQxKa/D3VBWsDJ8vc5387N2ROsOAjDC/+945QWVQoWwTRU7NmIjDBCvt
cHQQau/YjD32ScWRILg3MVBYF8Rw959lNP8P2Ojn8vF6h/5RsqO3E/qySoRHlqdC
rGXvdQELv+FNgJJrf7F8/SCwz0kFHbN1GBz+FU4I6SIyBrqmIs0mJjMkTWAPGufk
gQogvbcEgrNdMderonLS2Y/k+gN91PGehLlVjIZFUGZ+VTVLfYCAKKvMTolEoMM2
uLGyLItTXUMgdL5K1e6q8f3TokFR/oos/RQjBJnc/2ZoViU9inXJAh0lng9lZBU3
OobshcNgXcIAwGHB3PEFkYEkJiqCLGodFTuhrCT/mAhKy+ShFIISrmqd5wqej/vB
KGXjVKCiOe9NlXSddFliQzpV9KSjxPzFf7NS8F8V5g7bA8fEvjcLv+bygr5xmWVW
ZjJYBBDGQdgV64ieLdgWu7rhgLCq+187pjjPJjIC3dTY4eguCRmL70bajA+DXZW9
ilSNJFmGGQmbCZC0vfi9XSYdB7A8NM0SRrJ/u3uuADCaUMKYQ//akk/f4Bdq+0cf
MKbcBX+DTtbPVu+hvVoiLuszkD8wOlTSnKP5+e9GUtdupEmqdH+kbDUG4zbidKXi
aPaaqvt8M2dUha1cLrHc9UHyfJiVxHVR24tyVokhzGTYFsXm3KBzUHVQ70juBYFR
qxR0vtNerm16ofWfioKKlGYkwJFs5LmJIrcMasbRqc6sC/JtcOydpNhLM9KtIZnT
VRjqFiUq4XqlnB7PJ4801AKncDGK8TsSsiQfg9tJYOfuwdiImaQeN7NgOcTQ6y5K
CF1zHOk6+0K/W4ho7Z5huSs3fu6XtfZ5w05c8PHZ84L/Se36qw05gW8SKnWspsqF
gVAP05Ky5tJNfZCN39PpWv2a14vs/8nEG+Q4xMGbs4FTDCWYboqL9hOFFo3f/uVk
O64kumnXphVCAGYD2U/6sFAH1/Su2/jqYmH/CGRIP0uv3ZF+Xl7vBIg822EbqQ+3
WKj/LrpWcxe/otXLzWmSb9V2QsGer9+4OO7wh+5KT+HUC8WP/NVw51Ql69y2GDv4
y+hjJmOYN/4emmOb4D5rktaANMv9ATv/QBgrtV4bwayYBUfhaVylZ/Y4RE4GB18u
zADNDnhctSIvRmrODKMADppSNyq+AGQd6ImTdu/FWhR/5cSdq2VAys62u4qIIKMt
0L4BlBtwjETpq9FgJ1yw5TrW0Z9nnlWcFLNsthW23PSGJeQuyakHFe7byVtlXVbX
rDAdGS+Nfne9GTkvdNOROy8kO8zJH+6A+l5nLKov2JxOD/L6wKcJHRgwrzA3o6W5
+B+RO2ul4eIuACA0yT9Ks+FQ3Pi3Jy7i8nomTo6/oZq/AChB3WBituyiQxqDZC37
BeeMXF7aoGqmnWLnVCYlyrOAppinuZb5cLvew6JPReJNLJ9Db3a8BEvBQHa3/Eia
tddj+2viILRVN3BG4bozr06150tCcc0jJwgp3zvfi5aErSUDkzvi839f3DIttFKd
S3p92JSZJ2n3R1Tmzxy8NZ2wCv/T9RH5DaWlxFNV2lmoafQD4EJFcC8dZgTFhAFt
jLow4gI1yc443++NoKOuoj161U2v/Nfmhq2+bq7A8sRQXyH0mi8onduxsrVWy4F3
A67bsiqxnG7RixB/7D+3nS7BvIRX0oTmLubEwzxWh4JUxIWXdvtJ/HWFXGbJEYGv
Zwj3zL1jQqMBxYTsAxMWV1cv6D0tvI5+hMa58XpHQTeLE4Xr8KUPpv3D8/ml8vVx
Cmxx68EoRjvH5Yg4lpqztSspZ4/kuIfOoqAzsSXbyIUvDheyzR/BtOPMiNTk/XK8
ea4U6IMx4+j67lHoi1IOGjGPhDbYX8Qixnqz5ubQOntC4CGLXM3ntI/g3dqZoHfN
SqWT5dNXxGpXKFoVgudSu4sodzXtmVkeZGio3Pm+MbGSdkIEYGKccIYUSvj8QWUI
oaxEohs1P0n2KX7V5ZP9o2R2936ITyntcK3JdjtW5j7MEbegHXo5FFIJN41tNy9i
0At0XzJtnj/ycU5F4SuyS7pqOZJMWnG94JKmCilSkYMN971IZWiFxChSN6aDOyRq
5tAkmqdIRJsdlIXHmbjoVlf+NPY93U+Ms5DPLCpwY7YtB1ai7EgX5HMnYSIW9NPC
LofLj8pzPYiic2e9zPSoYteGRgDjtkzh52olY8PeUgWf5S6/d9WGeVVUtS57F59e
8Punl8jcyfNf+SLnlnrjyDYDzJvHmgq6lWNSm+bI8sBn2a8FFHuGxM2ccx0ESpcC
9xh5yMUnQOQsptDYJ7dmZx+l5SA2N9ahm3TAAhJiQTHpJLkOQhv1ac3pT8msTJU6
/tQAOY5tDV//myVOG93Sb7hDIUxsY2yqIO7x+F061QyFDAxLt+hvo0vs4m/OhPWx
yO69DDdalVowHI5XelIAyHLdYmpW4ITcrF7P/Mc0d4S0ArhOCKP6/7MBedGu+PNP
ok4NlQEaBcZIb5tNePmvh1ERdBgx4S3WD4cgTuHOs2nA9Arn0m7b1je4ULtToQR8
q2v5I+4GH65tGZVmlaHBHodgRzW8Klni+IRs3wolrqAzxyIVl14xx6rvdJLOWKRG
oi1U8OPo911S8GJPeoIePbogNgxbOug9lILRA2tOiwc7S9NrBdsht4bQzQ0B+Kp7
pOr1re9ME/dxHiwrpPQ8GFt78vj74lR3xZBv86X7STcAe9gyqdtgm2hJtTG8SVqz
Yc7elczj/pnQDkZX/xwQSdRlNPWSjZjL2hAK7C6tWN3H0OfX+mC6NsvI9nhvrAYn
dRnCUym4hAKPfkJZKxgKoz7xyMQUszR+VX0Sggf+EIsWPGKqbVuza5virPx+kHsG
sqltZS9gks0+IEueL1/Am2L3NU20KOruTbWjO0jIbg0e2ANenbQfT2SUC5fRci0r
hjF7gvnkDyynSRgO0jVJ2R6/dX8lnCSg/r/cVnYt2lhM02qG70YwIPCHzR1lkvox
wNA9lqO/WoDqQhlqoFjBflichTtqAtL08SCGVDBlxQ0R9d8DMzBwims1JZfWNKkj
eIojxlA0NaqOLYULu5/KuSaDr7kIAukAcyNTJRLyiBLpJJOS+rt7wq1V2YaajpeY
EjxEZ1Kf6xymG1aCdvYt3HB0Knhjmi7KhR46tNfvDTC0q+l5gonPeHmBXJypFgYN
kNU07jGUpuLVFzuNHo0KoUiHcUSNN1erGYvRG8o8M5LMktKZv9Pm1f3yMiOpNhNo
cBjYCh0ZB8M1cBffIgfbL1UEsryS1axtbN+2rUca3i3O+gNLQZLdX+QJwwpWuNIF
FGswIccDFh4lmUafd5xmcS71v+VHjchzCwhqeIOe2L2kVWbTKyo8sof3ufZMQ9OQ
4QxDFWRQ6zukavCbd9d5Fr39qNtz3SykR8K9l58GQpYqWUDnJZbmGIyqHn3wls5U
hIR0kfA5f+AEFHuFcbUtjSjTi2/uOzHA2ptV56Zo3OHfO3pRW3tPMdkKhM2n+EOA
0SgG+5a3wn4qrI/E65LlkNiz6yUWth0iBl70UN0GE0K/25A/BdkkeA7gICaSC8oL
p1DMdtjUh6NN91CF9yH+3AHBpsnEJuH+Oi5RlM0NeJfKD1jXtrplBcpo8C1byuEe
po4o86Uv623h4XJfStcBPeW3EMng7kSZXvGgrERLZGCOMIZocZPrZPkRyS68eQ8I
KZkKI0OKwFcPzIXam/ioXlH7u+GyDqEjqV9YbkDMdbH77KRvpqtoaHLKGsmq5F87
2vAkpqEe+Y1w7Gt4vTOJghIIvZc9Yia2iQdDlYGhUsHoEp0+XX8KaDvv2zhSMdF2
MEL9aC3mEvq4bEecO/ZnxeMJlUrDuQvyaRDcd8L1mS1y6VepykBZx1Wfib6nbWtT
IpCYqYr0x33fahVrguNj8LvK11J3EyfchpIGsrU6CV4SB0IiGymQkNAZLMomhN6Q
ohHrzT+Fm6Tx5N9pjlAZT7/qQAlR3i3X3bE1j33H29ZD0fwHLfsesNY8DVn23Yn4
vY5FS0jChv9GsqrvVeSMcEQ+ciayke+kSVVhTDivnIkcRd/BOI5QEbsRglltbCxV
8UsIXcIL+V6pmrVmn6UFnz5o9qHp/hetdOp/v9qh1K40otzobpRYT+/bincnLIoT
xgG8R1eLenU+N91LnPLbeED7MDwEXLWrc5OUMZ9HtZJDOy7HbRo3byTthJ8W3gGP
Dl2w99T6+YQ8IO6yR9DThtUb23wbXlxI8MJa7H6Z8+IHypOq1d03Vr93kty13DQf
XkfoQAt3Xo99AcoLIPeycn8sbaJRzl/VvNtVg9aSPaJ8G57An+/atYAOniVFZML7
P8URR7ZeZj5NEOESiXKagxc/wtqQUcnfYLF+Q9n+IBb9HZ4salBRrVaEO1nisgs9
K5gBS4bhYknihlVh3yqkxcFDTRGxEF+JzRLfAaK5RBb9vmvJwEoqwMLX5fkAvHkA
hrKlmJtH46G2c++nwiJmk9eMJ2qHRWRnoPT3P1H7TpWtFuS2CIdmkqLV1ek93wtN
xpy0orzNXbC3KkHBXHds4RLQN0HO4YOdLP5uHLWV0GX7tmoJnnIQSHGKmDcUSY6m
nqvON442o9xCCzggdCXNHzeEoYmMoBbAy9Ywd85bX8DIOjXyI5adtcALY6f0Sqwk
y8c7Wz3j/H44iknxbFtF8mRWGeAFsikTjHFt8U1MWXtnlvanA6cCHpC1ohn0/aM1
l2cFyKsYmdi3wUa5ClmqOfbWrX6cFo9aRntljsHR23j0RY6Yi5ld2egMbN9HnY4w
EtvcnXz8ktrpsA/EOxp7aLSK9uMtP7nI3GfqDT23O0WfLM/QqvyEkJ55x7sjQJY4
jVB+VZJ97FxwI+XwY44iIY3QgjtJMCrmzk5MHYe1L1qDZyNXh4rmDssE9RH9cIbe
XAIM7hfXSm/IJm4HwQ/akO+9YwSISwtJdRBP4LjnsKaOcTNHBDVEofMHkrEJdpxz
XSTG1+8JvR+ZYtKbGhgJH4gAZDUGw8jU4kZco/3kprjMWiauZY9a+VPIC4KbVe7K
D4Idus5OXbwvOzk1QUG8oy3onIQqn8VgZzrk4uUcjzjF0X/PL3iKRxy5EEx3MQmN
c4Kwl8bCeDVKamPjneKEErPnFs+QBf0+BqfFqh1I8NqnrqUKEDmcto14hM7giC4R
7J97hI0cU+JiegzcXkoKzrSJSBPa+ptNro6giuDvZEp0KdOa3weYVZFgXOy+h/kr
R+TdRIhmpQVpXWysIlJsdVDEdC0C3XV4cXbTQQEu76oGwJ7MlGWP39aq3227ffad
lPzo4ZpYnfVdZzMfdbb0SULxbr3Igh1f2/A6scnsXJDiJyRYBsretF6l4ggOSHRx
dY2S3tlz8uO3JGgDEKLIBQ+xi/IKcPnaje6UW++Gf5iBnQ3cRJM+HRJsCB/eX/U+
CHexQZFvZpTAi0PAXe/Gq9A9kiwLGEFXbUexykhj3wsAbWZwDbILm2J+MlH8cjzi
z6vpMRem3LqLYVpIlLcc6eUnZEutNuBGwPLYV1vRgwjdEELVmlXDir3ziuLn6p3j
WEsECHoK8P8JOYfrMEglHfIw3/stQDy/Py2NRnnrqV1/406V1J/cckXkQBtAQpq+
dJ93mBtnQTcecVj4dzIMv+FEravKLQY34XBZBkp6JTSYnbeDwd0d2dAk+YdrDC79
85QRybNOI3lonB5pMCwYoA8d8ml6F86zP5jBkg1hf1g3ceI2vNBbyCa0u6XEaweZ
q7pBnBD8YsGRjy6LQVL75EifSOzaED2ZKaK+NiLr+1wV2PtewlmClDVGddSDw0AM
sbFO6xh4oHfIzR9YU6vPSoY7m92aieYxDrBhyZZ9MRSdnDC1/vjbFSdfSbupzgRl
fu88pcTmJ1/J9RVuiEUiYofhZtEj9xIRZK6rojiGDSbbb0zL240vmK1pp0PHswjp
6L7alD51+aHUfXhF1HpaeHCM/8LF1BVXIn6FG6Yg1wZfFj8Fq7ncduo8u9CqMqVA
/mHUxl0qZC9w3ZEobFzepKAd5YTTrRNI/D+0isEJ+Va8E2KDMETy80j1uxds63oz
4pX150dizKuyM914yI1027vXMhvTg0KxD0k7mlCZrDvJewmOnIHDtyeel90CII+U
OkuS8oa5bEVOHBd1Cp8lVpzoHnaGAqfWbfQEbKiSUL3EKcGfBk9wwfjogDNFHWP2
DmjiGnlV1vXT2vIML0VmYcFFJ9BfXIzx9sCywT4MLuQhGxdu0ujVrubXw3hHUeDA
/8+wpgpdG/eJuJ1rEyT7D9ohXQHpGv+25g9gpiTvkpXoxLE8x430BW0Zm2oD+Pfb
r8sd0G2zjWwCHKRMF+UYFTFkKndE9XM6ERbz20mT3I/3N+Zs88vH00h++t1VNThE
E7JRaKnMcyZPY4Zw1w/D5Mnji+d0ovjAXRzZP/8PuJpb+nr6ALlKbaXTQtfbUGUP
9+z+CzGoCa6TwOhRVAkeaR5ST5tiLGU4rEwK3xEAcdyHM1rKWm79drOcF3XOhPmU
AnOf2FuIXEB2LIRRJ3Xn/KuqGMiLHrvFcUJ58MFoT0jgnXzr7YcsWb92xMTcGWpZ
ouKQLVbJZFD+7vj8xhYw3U7Akedep1kMUkKIGv0ozOiDmX5TByOCAOWbMcD/PyfG
NaKuvMAWut9VkBpXhSSrkCs9oecmIvycSckogmAms/Eg+t4kP4ReAFfZ+eohRvUj
BFQcsUS/c151MQhh2yTfmYRiS02boYd+LF+NxYextYozrp52ZnOIAgLv3v+pTHAI
ktmAwIWJmWZvIfZHORf1RXBlPolmc1ASrOX1ZiJITtnJrwabiJNSjG+DvleVuZhs
94137Bxw3/nWzUks0dHgjg6i+9GsQDH53JHILenqbXcAABTiFtLA9yRDfeO+CZZV
KQhK5NSTG5rA2ifodc7p28d4qqmtAVq4R8oVQgWassbBO9EzfKs+kpwm5xC2/QTB
pPtFq9msclKIvz5d0tO7TfYygviCbX3VgqK3Y/Nvc/Tx1BRl1+tFk/d/yb6tqKso
pBI1c0E2lWS0JKq2rxJ8IJ0JcCAf6vo57U1YemM64AvdQcYRznBPul/GQmIkZ+UL
VuXL9MV2Gnx23YetjbG/00NDTYNqtwaItABUIXsMcfMsJFe8V0wrZeQxfW7OJTix
fgjxDZcmBdskFSjH6Vn1VZD9SvYu+0g3c+emj2DFWoizsNDhjt9U4jkgcA5DFHcY
JEcXVo8reVB8kuXXq7Bh1huKNa6J4hGrR0TbeFAkgilKJfaJkfpZFTdvNNyNdda5
PGTWrP3GpGgiKOelgmzo6TSCngoFvugrtTaLVpHwEzQqSzbS042klwUCcEz8V0f5
o1hHo/biYv6qDrr1UsRZY+09qIIchV/K2G67FVKOXqYDmwGRCtUfwsfXsIRGuAIm
W9E/zVGqYYfGSMSauH5wGLPO4dd8Mj9QYc/K+koEzqijLN+xP1ZB2ZHWcgxivrXd
1R4TLuVjC4E87j4j9HeMnw3lPopa7Vv1ZsizessJvRO8MQv9rrPnx0pGwhF0GH9u
4cygkwqn7VKGbwgYF0yeMzZvR6YqHfDmfnJN5tyRY27VuhiOwx3aSAffCQSfr6D8
UGI9h/QgrC1k1FEPjbrTFahJhmFrN63aHUkE/abOR/CRAugbW1oN6OpMuu1H83+6
J+Ofz4YFebp24JlcK4Xzv+3bRj6kGwp85i4eSVKoSqIrOl7SJbJlpj27kB+BwD+U
dzNth0ygVjPNyql/8C7OsI6iZFrZzyNzV7hGk4uC5JJ8acw1iO6MDhL/YDfoA1Ie
sUDftKpbzoKdz1KnFi4zYY7A1S5Mkbb3L3sRLbDbgbYpyNo72S94uPPsq6KGs/SM
pcbIAZyxPsGFbGeBmZV5khKCatZGvs2CBcCsY3ugLT8UzCB+kYdAGkoBV5Xyope+
obEsayTwuCZZlkV34MKE+hHA/GNYvqg/ZXP3s/EG95JX6aZWQnDXBpXEYyJX77LX
l9OxP84cMmwDz+k7hpBSN8G55wTOPqhhVn0YBvDcmmh+wgnGehJaJ+0GYuPNrq8m
4bqllLW9DXn1fkqOlXPCIEm6zWNYm8OCAuG1kTpWhOFTDLQlIjAZqt8N4Gp24nZd
GUg2D2XjlO2qZtacruRQ1peumFvW6+4Q8eXfNn+rzE5bhwV4tAefRoZTTeihXox6
CsRDplJmnYjd7rEDXT2dysjar6G4hni7EgrpJwQDsTPb3/rAranlfDisoCBqOU0U
y5zuj7lQA1t+r3n1gWh+rbvvCUYEJFVKljXua1Ez295y0t8DDoe/fATSaKZoZNqS
YOFJ+U5snYZrmqs5+xwcNFLvarskU6BZUs9wlXXp1BdnsuRDE9tKZSnnYT0t8RKS
ZMkVtr5skVCZTvoFlkHkRifZr+lAvtQ6dBCrp/tIO9yh5BQyfqsLfQc1sXG+xqEk
o3dHB+DLX4Hpv1U5Mk4ssg5iCNpgyivjxeWaofjsOw7pcUa8ZEERcucvt1lqO4KP
KXlotZ12HsXMSyulYnoL4hE2WuL87+POu8ulQ1YJhQJxVAKtOKyTsFcC9uSHxlaP
OeZ7mjqBB+qcsmUdFAGc2dmHLXdKK4cHxbt3IUEzuzTY5k5ObOo99Cb2b+54x9Sh
ais+YOVzKAgbs92brJK5XSZQjO0u7YHkubhsds4QxfNdJe96vMHG/EgdP+xcnc+7
eZsm0uYLL19jtpJOVyTU0K2uJjbB06lhGAGebZT3Hag3aVppVlUFFruo5KLj0esg
xMOtU96HWwhPolEo2BuptiodfN7OxjhPk1df9Bv3WjU34/5bz4ONnRVFXgoXNg2A
R0WC7R1okKfUQ0YIiy6sJt+Fhv+Hw5AwleHiN8CN5ZKS7pMV/jbkM5QWYzXEBCMx
ZBXSCEf4EoB0MdgSDo/1VT2F6MxyHwNp3dEkPR5quuhHwNCTaNohE5DeHEQtNbEc
9lpPrUGy+uGsXz8mFsDVVtkWxcAwGukdmUE0rzTxOnhfmHnCuQo7zfXfMCaHUG4d
pCf7+pYb/C2ieSxbjMX5LjSrOyS3S9CTfriFml15yi3s3U3L0VWVcRLXpIGn69Ct
Q3owjJLlmy0/jmN0D4xA37lGF9DjIX0ZK6JKDuGdrS2g7d003LHCgkEm6CBWy3dQ
tKbmKs0LeMKB5d9K7L6i5uQKiSXmA/LHWB4HBK6Hmy5AUA9YkQ3AlZR646qeuHWa
tnPyPWN6tTg9IdZXFcIqqe8lreGzD7XXXLO49diSNNsZQIiJb5PJRg4F+u1O+pZg
Qsv6B6jL8zDx+UtMOaAfvbad6ommzxF0VP2ic7523k9eKOBF1YVhdVmaFxMLx3Km
SES3R+WJ9yiqpJn/c4LsLF5pvOLPi+jnQrFr0jF+6bdmwpBbU+rueox32omOe8j/
dzIlGOSTmozkT36QwnnYRzCrMUOofUBDv6wLrywWluBTlfEx+KUcQq3dKFf/d8/R
cwpM2f5nE36ZUfzQprIq1XxXnAYTBGFXv5IXH3EEHFfiAOrF8+3pQ1XwPQTdXykV
LQHcNM0UoED5D1g+jW8Hw8gtaz5UJ9NEW1hiFp+leKKLnWFqy1/d/CASw0aHIvQi
RY61Gk4klyzgf3badNaxU48oML+RLbxbiQxUDjI9Yc8ZE45iBs0E1Gz0PJxzYPrt
iyWd+owjZnybLb9RwD98hf5CguXsubzoyyZrcFSZuXgCOAH/b48+AT3IeoBWfI10
473nZy/kHFvHdEAZxHTTPIDXQ9AQhLoqCFY9vq8bAKuF1h9FNj6FhskHr6Cl21CQ
sOBQlG0+23i1AiY+k1ogdDO6w+qwtfTIyrgxi4isCMmZkaQ5Ld8yOLXAx8ur4vZ2
pHNDkbXw8ecAK4C8hzuH08Iea3O+bqCQeQPgThnO+w2UqBQTWeVn7w3cxyD/xc+H
dD6d+sPfZWTeMWeOEK8FlVbnCzZ4Xf6btIClYuBHTb7sH0Qf5Msc5CLg7qumf6TJ
l9S9YU1RPEd0wFtTWtWgfPdR/sgKtVB4q++qZuxvjhwz9vjOpjO1M84J770PvVmB
IcD0VEuQzYmku+YwgMaOfRFaRmZZXpe/3BGj7+btNT/G2nIA1+r5B15xMW9o/GZZ
baw8jLuRqxLU3GGN0xdtkVVow0FwAfqzMMLB8+gd1gkTN36B+AaolAKg1KgI8Mc9
XEEQYQq2uaMgwcxFOmTaidaA63sGpIn2kwQLcjC17UkEk5giE8Vi1UKpTFsqNMuP
yuljPSctlrQ7oddSCfQRtidEi2DwDzTTNgLWy0SA0T/jO3vhXzKnK8mQPh6Goj41
m0p5gpl2Dr1OCXR76+bA5h6CZHCB0l+twuU/Gx1b2HqIujSwIJ/ZrHRQ8roYmpYp
FUvQG0Kk0RCxijJMWagho4I0/MHlPJUm1sG4/gc5S5+n7YAHkY07No9FYqxp7+js
aNITIUBCwDHVZZPR3Z4/WoIrBOPrSDiEIc9DwuuZZfom+lcT+/KIPr4PrgGXIRUl
MpMlNShUZ6LELv9xCgyKXcDZxREuoYtw5aVaAH3qMTclTIQi0yTeDsex+nI6EFov
QyYPv7xszkyWQsWHAI43W5TaT1WAkV+A83BSHhGOP6kEOJXEWU2yUBWPJujWgmv9
FQ+o+yVCodwnUDNVIZ/dI6XPk//jzyCdQmgYOOQ1O3s92z6zFclyVeGQgX7cQosY
/IMTIAhODO1ThWUV4sI6iJVbkCyAF0LseeFqWmuoqwTHVJFqz5/elr2WobnG3jVX
1x+JlzqN/ugywse/WAbY07LoasW/dYUPS04Hwc+seRJRigynsczgQgEJsPfymaI8
KTRt/BGZNMSV4VaghBK9XjwwsMkWaZErGd0PQjjOZpnzes3SZQ67EK+TWdJlET9G
nGBkBO4jfmjejVAIFil6ilLBj2D0i/zrtWTWhEUNlAO48MykSv9/ctTqYzIt9ZcX
OgFK/GV3yUohCBtVW+CMKTrS11n2stFXn+hE4+/keHnAuC0q781tLMeFYbOxPXlr
s+dXe+kRq3BlVs6wPRdX9fBXy12q+SuEgqpIRumSMHxPQKGzv73/bRHWQKd5/NNs
uCNh7SW04GHjUmKHJ8BE340DmyMP2js6E9FYo3lugK/uEPpLbxyQMjAVtqHPVopI
lt8PfttDM6bn9XtfqyXEmVce0du+WeT+OmEYFd9v+dpPOpGeU//z77AoQ313JKFX
G/33IJq9nvtEH0O/z3M/xiq+acNT/ynSvnoGDnXBUmOWHwUrRCLhHen7nbXBpcls
Avr3G5hbbvSHweHxNovSedCYbdKlJB6qyuryVK5SKaB7fr8B1G6HzQZYBfCXBFGT
1Mo8rpRr5dkxDQSz5qeR7ZONtL9MSyfQsTIBeL7Q6V6ozG+KNe1zNKd5tnGlGPh1
O0DgVIktepB7t4RoOtdhL9lfKGVCC36ZqFIw5vdvQ5ODYgJfULbj/9PBZMdGuMU/
hnVe83krjycJ9Y4yhSCBw62+WAOGUa5Ct6OUwBEWcVF0hvekcd6AFAFanGgpZ/WK
ZrM4ifpRbqWhXR2W3sNZt0RH03+a6UnpMnyLSkCwG5maU722XMVH+44NNjqhNf0m
YRWoCY741W+JNQF01Q6TLZBbNbw3N0eIVuKFjUtLJvoGoiaOUSXogFi+9nKHe8JH
hXp7kIjVaFIKs+tgvZzbJv2fxqH+uxaDSlvgP3t5pV34Qv9ixFvXA7uv4erRZI1W
gfiRl7jclJsZDNpkaRHqse97V4p2etbe4I5cjK8IwxxSAtcha+/21kCvaewj9xQD
4WL0bt4xT7hOKfCU/KsMYJaj2w4CH+uHyd8Xsnhrr3BQJ389WbZIJNSOccYbBfwx
0XiI09mL0izr8d4keB+PLFhZsBO5cGZQuzqEyix4uqgJYPC+Yor7ANUaHIMbWD9j
c/BiddZ1N4Iz1gZyd43VfR+3JoCMGm8e+s4zlwH350mYDc8O6EChmiawZtwcsnwz
o9ZQhrubyOUUQugteW1/Di2wBCj/RGGNf9fDnxDRBs8WZSbPFT/1C+KtaZDCVWcD
OO3FEqOCP3LzKpLqhP7uvUF9uSwJ8FpBWDJokRcrmBmXr3ZQunu40VnrZ/WpDmUl
ypf0Z+JF6Y1+dxo8RLHJu8VSYJZCf/TQv1zSACQ75idOZ1TrrEKRm1UwV3adg2gt
k4Ant6E7d2nmdq9OwiBVJHuQNp1r6hT1q0pFYff2L/g8/fCWmmPHdMlKon8H7jmo
O3izfT+4uSJwP318YTG2HK5SBcwzTornJxhbTUvzVzE+tPOkSjH6QSoe6KpKEtVS
TP20XY5/OVmEQ9bBv4lfoQNpAbGf/IL52lbraPsfXz9DsMDYLQ+MZ9B5Wkrc6sI1
9KXrt+IyiL1+CH7HNh4S/SlCN/46sqtUwUwDP7IWYCVlAl93TCBp70IsTwWEQUv6
wCDGK4uMfXGGB/XJ5DC2HnkAwPx+kRoMr1voSFZtLkyE3JqsyRzurMe1cthCpMTP
G51oUCCtYQ//bfngGT07thKn72eOOcHAd1rrhXniL378eOt3s2Wg0Jacigdq4P+F
wSLBj/9VdbKv+KUH7NTRGNd1lGAnSEgkaM670jp1Hsydj8E3540BnefMcSLnGIGq
zrHF/HNknNZZiJt2uHg54lb6kwokTDdfppsQaQ4AnQ38OzjjZi1yQNpw8GmfJgVL
KJsKBJmSGisGjBGQupNK6xCC67ddMMlGnakQ0dKucB31nlrQ/aVX+Jn+qJZmmn0+
Pq0sB1S3frAUDu8hws89p9JTv+SFuYJwGT9pNrHzQX2c39k61i18KHx8q1HOAxsL
DnbRQ7GhKx81+pEez3CwwCakBI0OUVKn09vOY0xCF259Edfc7uqa6E/FaxvznJl0
5ncr2bRP107rdKyBp6MAiUXoaPf+E5wigSF6Saj6nqD+8NqIDUw2DTj7wihaOXtT
WM8OtilYYS3cbz6/7iFQznF5WVZVcrQ6r3prw/NFf8LpsVzgru6Yn9zSA4RmZuJ1
n/NjWZELMXMHjJ/xMdykgU7GdD4fZ7rdfsJ7uhRQUCsNu9YQeWmaPLop3RP/RoOx
NrVddLt4HFF3Lj2TKMQv83YbHvKbrQwNI9RLroEqUUkePl5nTAJGA/iMpc/f1tF4
ch0NpRtYLF/X3Ltc0HW++jA9+J3YKmBJD9O91rVWX/4C9+jwD299DRFROdwlb8yV
61ADUcbqtejpZxZt85plT3mqBDMJ971/Dl7BGUUG8UCUndM62Ov86lAD7fHk3Hu3
MjhgaYqNFUkpV0SUf0aDEaEBqVSkNsVm0abB62e9J48f3vfRNOEsx/tcqw2gwGyp
Q3qfoBPYOxr3sbR8tCfDqeOVMJvVYOIGY6Y0+proiNrEcGG9xwNVfdDwJ7QSKIUJ
A8GZAMx0lAnjYI4lfEfYaDurq5wy+2oYBPA4OviMhsy2l9EJFeqmifIIvGoTLsxw
WiD6ohD/fuo3HFQrG2aBGfu1DoNYTMUxqiyN/AFE4wZ09tHzrMP7+q6/RM0kE5gT
wSPw0WC8nmRX6ZGL/hYOPPeFCDOvN1Tb1nMAbqZwUFakq+NP1tALDnwQJzShZ7ED
2UrviezpEU1jYIV/EhaP0UNzuvcOiVGFcIQZtC8lvQ/n8IFdFvmG+jNcNZS1Mv8q
nnCOTrSHJ/Y1RLXtr92l62j8kEq20y8xOKbp+SpL8qkPgkunr0GdggWJEvOl535/
c+xnjBom5UHixKgH5wMWtQeh8eE97E5e4MzY5OZeAq2XxLlNhOUnmp5srkL4zl01
LjKHl4rY+2GgSBXzRhReAYsudHok1lDHJH1BCo4JezrP1+cbz4l2vYpTJRz1x5j5
iK8XekUPkpHgKEM03Ri8nVefvPCkcmbTsjYtSwkvhYWhqBQQkXVZVjKggswzWa1K
p02UxQ9t1NE0w2fWNo/IzgUenDDsMmai9moIeD0qTFhQwX2amOs4ewqv4rfoM9BR
Yh/xuYV33NLl3/llDDcryDVX65OVtfXr3MADXnxD6OBFMmvxLrPXJ+1w9OR2mUoa
GZRzHV3REEd8wEbISMGxEdNSOz4dSaA5eGwz5L8ziRkKrV26SWSMm2rIFS03hqNr
/+TZHC2K2L0Eg66p75OmKG3p7jIC/rIc9FGeQlrOxmLdfpyqS4GjKj5s+zezT40a
oNWV7HDcztz7XhWga4bWhuUPLGo9NH2MpYS651B8sHt6SLTxbRlYBe+vRleCrBCj
+8B6p2DickUeEJi9M20XD1rHzfC6MuNrjT7d8LEzSjra7AsPRkKysAC1dln6dn11
vbZHpyCfNYt++e+qF6PymaL1f1GlTRdslV1V1p230dgeMUxP8xW3ascvp7d2YOxm
rR19XmtTzVqE6JcBUVY16+xZ6mdPrpFJUHsj2ysiqPtc2zClaZHKgpymkLPlbcNP
eiSPW0qe1/SVuc8DG3tyIYO65kmSkb7YYEq4CJE+OcyfgBwZtUMFxbRiKEX3ThHS
93RO+795oEFcx3ruj4KCs2q/PI0YYwoigW5rIMmU0SX2ykYX99rZv4Xq1QJy6l16
v8TYFyXoCKiqlALJ5rjNMORjV/Ihs/yxnKhJIIULyF1dIUIosxii2WYNEGdA6d23
9Wk3hAz4ZWgdmIcbeqJ5vjcuGEpY4P5W1Mex58NplgSHR/6EGb9vX3U8Mrh4+biq
ZquF6Jf3cSjmPAQEe2s+6uRe+iLu/9sveRQMwS+9Tgw1OwzQ5mT+g8YB5E0vTPFr
202/sHrJR15DX+7G5zeT3E11FvhWwbZWK489s1aTA+ih08zCGkTSsJyeGrQB3Moj
H0kQjF9XsITQmVFi2fB5ARYNpXEKq305jUgRBG/MwwU9jwq/WwGnaYfzFiWiR4Aj
/2q/dsj1pDlQVe5RLU+scU6N7Sq1Ah/j7FP9sJfSLvU6oKqFdh4yfA4EhBfrcQW1
cxln9kJBQkoZj9KWkHAtCsfTeVf1GT97ZNQZC7KIAwq8q1rJm0KAZdds/AtU8Boo
tD1MdgJZjzO+02roBuPOajuk2A9FZMn+7qboEA9mEIpyH5lVEsURfoUsFoXrvAx6
hBlp4zjlP6XI1ca1tpJqoBJy1b46erqXzPT9MnFa/tAOuK8DBKo8MUZOyF/3L4JL
BA4HxfmyrtZKyIeglrIVt/8ldu7VQ3Iaur7ElfBqmEiFfn1TYMWVTMkKiy/I7Qk3
NVKp+Iuk97n7JHXtukweDpBZ5fg5hX0HyeEVfvmPKbkuUsqQMZAcAZcsbZp2QMEm
SIrU7aAeHbRGQthC2sEgFfNhR2oJQ3bv47DnNyzJ6FWAtMyeVjMkEMFcNA27ZyBu
BpkQiTZQ+Zc3krjaVyyOiTICVIid288Yy2vm8/Ezc05SAGR5f/8b03+DiO1sSTYW
ZswZmq90BlOehK9UWhxPJ+GhcIvrTzoRIhvNep4nGfN6eefH48IBrCvXr2+4gOoh
0qTQOMRTmM65MbU1iWITRNX866fz3+yMofsojrwrqDOR/Nd+6aw3F5ymw4YVcyPQ
3kIvQTU7kCBoBA/H2YGmZXXhy2CJQtz8/ZObdzwAfDjkLAE3lpI1T2dRt0z+naAu
Q4/raiNCbuT+y5KRe/aWqaFQak02J8bmcOq5ya/SWnSzOC+IjGBd19g1pBcrxvNG
L+rf9/nnXm2Hpqx4hHJvl4YhFYePMq9X7DWkHfzSuuI69ie9plP7mRak3msZRGDp
r4P3TVhvacueq1Ff7PmcL2Q0CDT+DPhqEuMoyXI1lMWYiOl5KStdgXqglvQu5dx0
rqQfm2wDJLICbEctyKeM0UJAFOQBzwESQTH0s91wkZI3HNfWOsE/UyqdvnuxXwdJ
bu2BpvcHBiWuMOBRYHhnz1sv0vimlPbUp6FRn5WjMCE5j9X3b1k+aAU6UZ5lXlnW
nj1nZv3J+Sr+HZ4rSM2Yzf2Opiaswfrg3l7xRkGX+o3X0ikgVVaG8zqcOiiHIGMv
eLfZ89qYFJwZWbYF/y2owPlOriwmde+7ZpU/aqjPih7V7Kuw8XmL1+vg+QzJtHcF
r3n3RVvjnOw+wPpyEC/dvF5Z2WeSmUL4SoH4s2uA/NfKQEjWelE6NBTKwkVR+856
cy80jG7ge5zXRHgS89pyhQe526RQ8qjd05plDEkomoRXcJljk77JxpbDjZkOl2rk
0fN0Fy4LhP/K5MLmGPn9SEOiM/y14diR+Lp0M8HQTJzjOtdtZPlvSibPzJagnYHn
G4NJZKyuIEvpMJwQ4pydWFPewXYxnFYXacJEb0FkO+XDkciQM1/8UJCfmvIvmAjw
K9ynl+M9aE5IhrqzQ0N1QwyNviw1Fvmdno12zGSTt3JxildyN4TJ8nH/dvWtCXB/
U3fpN8ruhKYDf1vT7CKJdUaMA1lNfmbRFZCkRiFtrS9URmyb3SbmFvn/4PWY9Rz8
uOYV0Hj+/upv9rt5GwEdomvm1P94L8wOLHmNBgWSmEDHsB96REXLxrv71NGL9gV5
PIgvfJrzoRQCXBOS+s7ylNZ2+EOBSm9rVBiAg2LJZBnBdpfJPw77amKXa5g7XxFX
k8s0/XpraMWuzW8WAhynI6rq0AIxJZS3h5VogVKbc/2ArzkGA7P8cXIf4c5itbZB
jcWU45lLPnc8N8dUu74qCEOcwgkcgOxCygS0zZst91+KjJkDjfvFc67fxS/dMGak
hD6ge7TMhGL4qLNaJZolTuJ2BUowwa8Z855DWvefyLQ6J/WNxmTL6dSz6H9zi55a
wx6Jlr9eFphvQ+5QCehRP4jvCoeU41t5LUz7tldYsXkll1hlgVJSuXJ6PPGp1CBq
SHl/2fZPfBTeE3HxAzoYAU99v1TDDMBDSDhgTHjGzw1nwh8aInrndFLl6jTLo2rN
8s02A/qy7attaOrXN+S4UgjF/oG4+UVm/j5T2QzdEeXQyHrdF3fBvUa1wEkXqXab
DtlhE+D0pAD9ov8aqESkJLkL+BbXm7fVVt8iPc10gX3YZXEg+05U3mE86xQYuR2g
9zU0TBig7hEERhxd+5J5xTMLkXTMMxSMHeHLXisarCHcvv5ujDpRCShKQwVt8y/C
WxEI939amX7qYwSlj7sbwvmlR70BqzS4I5WNfNoZ84Lkhf/wHu+cCSD7lMYBIczO
/aN36WPbCNJW0iziCg7PuZksvfFk7CQrOFsmOCmFeNAW9pKwYpk9gTuikFK9nFyC
aLVZkgDxKyeO3yQmhnpBH7IF2iCagbVTvCZZCQJi7sOk4c0/9ReM5BwxEV53c6dV
BHZOjw9GAAdCpmQz9o1/17IUk9h82vmqS8DUkWOAaSOA8P5GBjyVPyviG/X40G/D
73TF9sPe6Qp6TQttlf51A6g/FDVddLfC+BvqEbf5hs1ws1p8phUSlz47K/7gpxeZ
i/BOs+zcNtx9VMlUw1ZPr21RFUTiOxRbZlQ5gjbWlxAnCHZsxqZBOiwQSSnwojR9
48EhSW9xlyPJDcBDy4S4EJBR9wH5PLLvyRZqOlrMqOwkeVWonzG67s0wHIxk8Zfa
Jgam2VWcdTY1vP2Zctf16n1Sx/fQohmVtwDlx8cOr1lcYF/UL78MTFkg59Xjx24b
TGUObKTLpioTTcBGxbhja6WlkgLzZwJjegxl5ppGfQMTaFouOY+O68e5zC+U+ToP
1SkWqWJQbcJnfxeA+RiWjem4vMMRIgwscdJ1r1vFo1bQ4dbMCGhqVetITTqtWwvr
6sZCgAdzLYAyNkyYcPXGlVHXHI4ZnTjXGSxK2YImQw4vi8UghRY78wQE1UcOo+8I
wTnc4B4qwM3JDLIu8rJfAkdnjgIX9foKA0SPoeLWG8Gp6iDR7nOwwo26mAOOE2Vr
hMm1WlEGGKWexwJjv/rgKEVaMkYQM/3vYDefm5TvAIL3wTB8Zn4X883T75yuUSIh
+4eUm3TE+0/JipSqiDpMKEjFhmz8NRFaSyuZR+nRjR05HlKNLYAari+CF1FLF1/d
Tm5l07p9ll1ijQ107y1Y6OmhKAhHmmXpaL5MV2px/7EU42typMmyPaQ1N+iDxVap
PdAEz11WT50l6d96kZJmbYVuqtBwaQFgnwfzUuIaZDpMJmd9E2B3sGT49U9bM88T
bjj+swLNSI0vlcRYtYcfMo9eONBnLWLtS89yJ6jyKSIdHcSpbk4vJ+zax6PEn8fa
ZsPoq4jaXUbhhzumsmxSUZAz6AqMqRABLeXKw92J/BeZqI/RsCVWBIZicQb8cHuS
asuTuNRqOFD0nL3BRMmB2T1FwB5qJYybPtal/W1eAPRyuQ8TNwxMfQ9fDxSuJ4DY
q3QP9GHkGB+ms3VhoRlBBIFeQDrlJMBQcRJsB9cMBWmN/Yvy3OvHHTtOBymMDZ+D
zcsSuIl8ruJ5i0UkBvGIBv5SNr5uBEDM5YM27VMxqG4Fve7ikkfM1OFH6Z1VLbYN
PPV2c/HKxzq5idveGkpAwWJB2kZ5w5cmI0WLtIe3+iy1mhWk2OfKDgje0QTfUTj7
xFDUqQe+bpruua/dtDh5/TCJgRUBM0SK33PKwP58DJDrYXADsQbDaEOutkko1jYg
H7SIgRnMFuOBHShudxZuJUjtAM+kyXbniz4Nr5ys9UVIoBWW2Azczc6iJkAElwQ9
7cOmyJejlGcDymirntajU1Zyf/jHBqVGhQzD4vOF+d5OpJAMtyzRwIQUGlHd3so2
bkcTR/uH4DNkimsVE/ZObSZGVtG3cW+iRvimXpUvUkj2RIdnej/I22fiuDraag/G
P9xPz+jwTvchrRCBE4EiVL/GjRXniUPSJmD8uLy6MlzY1Of7RhX/LZ/X/mbV7hZF
zKNUcbZoor0DYqSijxzRzKDSiqol5qBfpN9538JU/5J6ym/yA0xOgeyrplelyulN
cz+uFMGhBaWRZnUOdGY5dnsM2Wld0iCY8BhGrEIHd2LMm1Zl8gA8ORTw2UZSu8dr
kHASQVgg8gnJJMz4fo9Wc3c2Z4c3F0hmLQ25bT60UFWonkHzNLWpt2HFu8bHXg7+
x9coEmXxVUMs5MfKXhhPOqAx32+8sc+0pSIa8DZW4c4HyFuL+bjnXJNuwZ5tUxg6
qiQsGKmgfZHmZ7r0v9BtNcr+FoHXH8ArRr8+7uZK7auxXJ+SVgDtbTQJaRB/Ea6/
1OKyjLwYeTn3LfyciCQZvWKqoYBNxKBFWTIvL3APfP1XR1oV7PvTzU09VBE1lg8J
xJL5ZWuf32+kXXZ1fklKNkjfDARvpWMV6DDmZ+gdD9lAeqIG2UIRWG+VMRTm4QVe
LsWd4nucleIxDJmvxCylol7TcIkqSNEbcBzNV7jGoADEfZxUnu6VfsZNbJC4wM7q
zo+aRHUJxw+stDzTG132qAGQT5TxJ1XFTCPD6jREbTMwcJngVyWpLF/j5Ss8amRC
4/WnXIbIuebyYwl3u+1qWONlE9JFEXhRBvBGwB0RpqsLRnitAGh2rZWBT3aUDwRi
ZiVpXkUiw5zEczPcEQOzbt41bb+dLHrO8OMdGw8P/27B7xhdHXwKg58unyZib4RE
3fibpBl8Q7hJOhf1IXGwALU6R2qdm4O1vDpNIuNflgbmmqojt2Tr7KOdoCf/4d1C
tPjkMV/ikxinLc6PSq3GpvDNesqP7xGonaxg4NSvBbyVsUXqlKMyBAavq5tx4kmp
egcZnqNb16vfFcaQ2YjhKTnJYOK7BhAfvG8Ln45u0axArdqbP09Rm0sFrOa75xsT
6mXbswb2oqFSfLeMmh+e6faL7ACoOW6ZKA8q/PplaUVEi0RRdF6TSdgNm6ueq4YV
89cUsf3n/OSTOKK1vbw+wLd0YuVAPVircT02csp2v1181rDibLB05NVmlkmcFaWo
LU1nMAdTdvysNJmBh40l7uxbvuVOZcrpJfxPQS794XH5M1rptUBFvNqRL3uAUxlE
LaRssT/XBbtsMYbzHWVgMHSenWWdYcYe23VDHEQJ+8BeLMar7oz2t7plDB21VX2S
kgeYoCZtKqFeBb7r+IycziGqv1B+YWn99PtXsgnJ6VCskkD6SwC+UnvloT8RKQ6h
SvL1r+0aTsg/jG/IkhLa6ezvVdoiBLQvg56mXDwgRpRx6rvv5S5LaAOzGfgi6LDP
TpvWkjO746pbd37mGTeM596fUYkE2yQRyXbqQAWSnylKXQwo3BMdfFaldG2WX+oC
Gd0KRbPrG+U1/tKrejofQjNE4LO+2YwWbncC1zTmCLRy99b6HY6Q2EH2Sg8ooHeS
nRG3lKhEGD1fc4j8qzMa9X5Iry+P/Mk3FdBDhdqqctqwst4dJCqjFXDZ/53ikVhN
763IJRFCj+keHGwBR6t+KKpXRSDP678/UgI3BtIzMjq1zUiP9SSRO2vE9z0W87Tq
+DTAS018fYz4Aj3Z7Bot8/gVHj0+EWpTuXehIDxEUY/9IV8qXywGqJUPFICCNs+d
ZNic+QDtL7tni8GuBNWkurr+gnsfP3jBc8DNrXAUQ5eToPa48oONKlDaAhvyhBta
KLGtcLcNigpbwtY7239EtFhVz8atupTpdbvvvFTNHCOPp8NXk8fGb2G2L9BfafRy
AFTb4buewpqdh0kWufq/H+LGAPRkMfHhZu+/sQ6ak0gl6AMbabAUBIWnDp0c9NWu
tyDKBUrp8ATBdoRpm1c/0jD3SKNMt3O54AgcO99Oo6ox8yolS4LlFoh7NoseKJKc
z65W1u4KnF6OF7RAVZD/2z39OMFEbqKClO3nTXlCL6otCxIF7W9yeC/HVlX/+qMd
rndtldHG+iKUKqEhDhG3P7vy49BpvWH4FBsjY38qF4mNRbEsyFTmZROY5nfm3QYm
37iD4pZ0VUvLmmKnXr6ZFqvjutCXB/7fXjZXGYUOGBH/YSzbu/+oce+/xXd3b0IK
GVlv13kRWwl/o5OoPF6lWHEYRIMRRbac/yF3GcztJ0GcAlOCR+GPsDWjcbBSTEF/
TWKEBmpEb/UKXXW4eaK3t+5V03KNIRmG55u1gGzsyvXUw45YOhIix0KjfWzzJXEH
zib7Dz2TYTD6aL8pdo8VK+snCBIgYdeM66TWKqblpje9drE3E0Azn0LfaaBdUcZm
z6J36blClwSnjfIN5oZtzy3mQYo7YsIH3PW7YGTJEKKFT8ZUEO3Y6Ys+LB70/ct5
ba9aZnARtcawJzTsc0R7PgHgNBj+gbngrcVdHPkLp507Ep3xsCrYJlpYAgZc3zRn
l2v8L+8qxiPsWb9d3j1zivk0bz1TM/pMlEovd/wqckP0PrmkWk6x/I82DlFR7L79
/v+Yl0oE8A3xy5UidKIK7MPmp8IhXC68C1I3INKbh3dLPsaVggvW12YH/hEactNu
p5+/76kmcL8SI9/i+danycYeXa2m/BcjPSw3gOJ2QyXb1OcpD34zXkMk4bsd/Amg
IwVPnaSo4GTT9C34xpC1S0lFpsKqaJth4I/uaV0pbiGRPLMRn2PAeyaR2cuTdtNt
aOrk6pPOxrS1TxCZP6MJEPrcQr4u6oV2LiLbLbqKhh4DfatQrpxhTJmosteXe0TP
2JcY4yvRBhO1scJVYIAtu+3Vzaj70Jfb6A+4uZfqJoDvErOD4db9mWU9MIu7GOOR
lGKxZdcRrQEfkxMYy2lWYxxDnm1vU9ntSBDfiHWbFXka+mOS0Pt8ueQpkV4rXb7r
WMkcCARBkScVl3qXVH/gfJLUfUAikvwZsSszNvSMjdSCwjPt3rL5zeL0dqwJYkI2
muQiy943PKTO1EY9iK+0hGKKnV+/6XMHarD6mZ9Bw4EDFZwfbezqT9QzZwOnjRkm
MAVY5mDLGNdC69H1Y9qelPR5PGobEj3dnDvYchHrmwO0gdYJacTevTpZGHarFNo9
sUYJ6sia9P7WqCpzawvyj8e6QswITxCbzcVPlDmUfd7Kd7RbUi9KmuFQqIjrbTQf
lFmJgy5TfKVkTzfQgjw/lYEtLjkBtz2SKRw6/vKkpG6BXj65KIKPVwOJV/JheGUw
2AjkFisKF06n7Rvq0zagaQ0ijzCJliwDolNk0vWKDAwALSJPTC2oA1dzkPPQcyo5
u7o5vkL2/87F5uPS9rCS5lnfGkro03dUBmJXdT3omW9y09iKnrPrg+ikm4TTC+ok
15ubeLs0FjTza6vc7HXfD69Xzzv33VJIiZ9ud+YSmsOPCNrmz36K8QMqdOyjfyPx
pyKpj7y7A6dFUCpY9udIYJ1WsMryT84qQn1efBxkMygpmNr2JVHqBnrpCCE7qdzD
lwAq5xnJJVA4KbUZsD0u4Q9DF2UYun60lXazQpw+oaWmuvDM2qab0Oh/74M60J1A
/NebF2DGRr3+HH1NxGUSFTgpi+rTUeAVAyK+1qnKzu1a6EJNBFOzq0nCo38I2i9z
CSWpotnkBKx3fBfUrwrJz47X6DrJyMJ3TP99bo1nbNV26jPM/18QrOZr6p4ZwgDP
w7mua/oc3dn9ezS95kxESwJlZqkkpFhvgd6bQScs/TwMOQcsKKfTKFVZz1/iR5Hr
hkM0SaWSMX1oLGbsTI0G9kwAQG9rnWR0+CHtsOyBCYu5D3WeKQo0dSbChZfQVrhk
t1Ded8zKcWEC0EX2EFNPHKJ/9NzeV4zsN5CpjX1QPA01QL23azHx5vSS6SxOuCCY
C0LtFznWVr0bajklHfPrMfvh3RUeqJVYYVA/EKBlRHBGCUUnCZkaonoB6rW28UUG
H/Tl4k1JlQvoityIa3xouU1DcZPwval6mW1vl+sEFjAmVvcApNFzjylgBJVTPCTV
FT9O5or8PYl4qFvdgBe4gSubpgu5PsmJXjKKL0HZ2xJDRO5jjE529YmoVc1Cj2cM
lkS9pwv/nP1+DUed+bsSKkHiaLl9v6qc81bLRxaNIIn5HBvKrt1+pn5DsIzLOW4q
QDaW8/1vwI7GcN5DRJPKq65Xy7CWMlb1bQA6rnzeVMufz94u4aUvYsHpm21bf2Ui
e0zWhNxlavyeec1IuRJyz7ZkqxR+JLRHu0lsoS+d6KjqyXEoEp3jWGaM808WFv9T
H7ua/gRKhGW9R1sa4OJBE+inUZMCWdRPOvTUhujw8JaQ0+PZQEGhzvaS8dJv5i7S
hw6W3ZioLA4PjnVCRvLNHxWeyQ+JnxMN4gaAF8ryms8SAnALrGIOpe4+TY9RjtXJ
RoQI7F69BO8P0R/DaQ3+y9laOzgcz4NdhSUsIWfFPlJWf2XtNGL/d1lpIiDKmn1+
DLEU1yiOAsVMUZw2IdyHKV/dbfQyQcY14IRdy6Te1/t60Wk2dAOKJ9maJCi9+uVL
3CFCBX3K3SIYPyD+FE4FTGNXX8EW3xO4VzTi4b2ot8WTpF11/wacihLcSrXGym6T
DoVGkr2/NHS6XeBhdC1jLT+uOeLCM6ejGahTEXmitXsxSr37OBzCaS32SqMo2X52
a9gJGMjhqL7cn8c9v3SGwePN4Hv86twm7XjOO9mrF5HEvBIUr7yo4Et2s9SlcVgg
hNXfswrrw72MOrq8p5inbh/IfNHoZVFOpCkGNoNFYSbKP/HUa2jeGGfAOBScsbP0
CcKg4+JaaStRdv/ez8ry5CABsIXxPzn4G+ufwunn0DtnEBdvd8sanNks79ofxbL7
IpuTlOKwJUS+p2TALnafV9pkw8V9an75xWcNL/qnOoY8Q8Ai7dyrj5hIu4gn9ls8
B2iL//rudWm7nWoanPsHTFTDPf7ObHB6QM2OoAVbhGVkEWWYMH4C3BcBpJ45+tKt
SvWBCQkBnUgBcorFO0xYqtJ5FVdKwl9dL/TsOQya/zoWAJt3KYLz5pRiL5s0yjNp
+3+wKt/DZG7MKI4mTpH90j6jYiFFHGbRN6Si/PwAWK8DWeiUcL8DaTQXWgvwfsep
4tT5+vEg1UweB/rBKEyZD8BAEw6xM7mAFf307Fv9Y3sHEWVr1E46zwCPPuY1IZCz
f0U58kUaM/k0MODJEYipM57YvnNEHmzEvZ2AnNq7JRGZ+jAD7jfJWDyTOe8XGjc4
ffSSTCF8R8CCB/IwYcLVD+1jL/8snGE1s6JI1ONLaRGkPb6FoJEbPR4GEARXKUT7
Gp+3kG3P9cOPmOBEYX/lN6lym3S0iQ9EbzuyZhKaKrl1Nr/KY5BGXIakHMepszgd
vsbsDH9PSXTnKTjR6jaQGKCETw2VNAg8J8lEUIiXdhMcxkKIlLDC2+/hgnB1qSlt
rSIsuq4Lijxn8XIravLhklBFL6mWADbJABpHlL6KbMONXZ/vSJ5RGR+cVzZnfG4z
4Or+zqn5j+uGC/SbvgeaJO3phKcv051L3Bywzi4/zAMugZHBt7lFq9gy7j3B9Pdg
I5h7anZLqgbp4YRhFcsjPgZy0ggDBobY7uMQ068hp4mvXwAhqjqUnVn4UyiMgdAf
uwslpnZMoJNv5X6juUnlaytI69JiFVCtanCIM6SZzPOrmLDQ8+T7Iq/01N0X8xZj
0v2j5pGLBfbmDxdwORH3Cs6tilyi6w1M3pwhmrz53REMt8enU7JEXsDIGQYJn3h4
IrGqZLlyNKEibID+umraIh/0neIUhXaMmBWsx9im+4Qit0NoeWC6RFeletxB349A
Pby0xABRKl1jrqnFHup9lbcjZ/3MYpkS9wvLqmu3IrqIJf852nxP3c+EpCHI/5W6
Rz4LsTmBPGMatINKafhIjROvYk8PRGSlzPIn4nAfj++JZ+zBWNfAJdikyLqwPXAh
83eLOrJXqe36sf8BEXZrjUgrExKxcU73/7vvNIgzsd38PaYYgNUbfRJHFG7sbyop
sNH8u3WkoNPlTTd8cjBrnAIJINcaZJzHPz/Hrk3nNpuRqsKM2muHch9xOyA830wp
t/4XhkIyP7qbhGlkpnR+Yu5vQaAkXUJkAPbraohXm55waQJXInNvU4tNrba1mnIz
5Ta+4Klbt9O8PhYCQVgw+evVPAY7UNj+701h2DYSCPBWjVP10wfdEkTDV3ZAEFuO
GPI6n4gYP2tLlPZlmMv270AG1pdjwNpctG8e63eGhyCGRQtTcwYdSHN+rmT4o0oB
iUmUxV7r0fqb+JXmUASUF77xjJvTVlEPDJbSmgXFAm1gX2rH3A9AxPey0ENT8+lS
FaI6knGH3Mf6B6gQyA5V+R+PfaAGNrwbGc5tnyEWZwS0ka42gob0h27GWfxwVEJU
DBp8PGAbkQZaXL6Xva6rbL2N8JxHwE8XWGHLVNNmn0d7Fg7F0DIvqMSuVPRnGr7V
3UyzaxDXojYmGkRSY2BdtEiUUZyn2kabUyFfwvublSaRlTdV6I3dM08vQ9Tdu/0z
kuHqaX9ohL8Cn23W3R7n/u8oUHKn1jaJwrebldCtEXWE2wCvs3AWXiOajaHLe7T9
FxoTJRPtp7gmry24CUuwAPbM/+AyWG48R3VO9YrW4HwImmrKexIl64eKsoKKmv+x
MOrsOy1Zws4ZrtzOLa596jgkLWxq9G+QqttO4i3A73FXoPSNBmX4meKDHgynH4E3
+xpeyALBu1N+E5Shz3KgR1ShxjsIniGDE3cHFdEbrAxUZ8CTj6gFWnmkzcqv97Ll
mnH4sAumt20W2cxIiDA4oBfUk/qMBmKV+cZkSqX5DP6tJTVAgoXYubJZwSenEHtp
xEaEMc3XQEPaz5p8zLi5d9z1a65dRpLs+GnGipQQ3etjKhVkKUpDr5BBDTxvxRiX
UP/iYv1H6O61K9U0mQ4k8hKzuxSF6+iQXRHxOhxJ8XN7zabYWcZmjfLdI8aEhPmD
FTzGoAkH2INHLuOos96qYKEWmw5mhILBNczT4sEo9dLdqmNwmpWVGrKpddLLyNFx
wtmZaNoq71rMjInlSWkzHzRz034psNL8c9uUYzk79jzcWl8ua+9ChU3gtAAswvCV
iciUWCoc+Li0W8v8LVYBQZa9dDSvuo+MY0tjtrkbsQEg/MAt0LXPv3Yw/cC74eDj
3hwNmasTuKo0UGXj9ZJg+9wrLFfjsF85F0+WghGxNx3H3HGtQ6ZOLiCGUU6tF4Bk
AS3ghFgjHuDGzqEA2K9M4ykFfRlrcqQpcD4xRBQFY+WOa+8D1KYS8uqhTxMk4Fdf
tY+I5jTe0bdNQNOfg2OQn56XYUeO//VwE2mncGoNQPUAIphPvjJe0ngOpcZe1vQr
+8RQZ1ndp/cQsxcoiBKAKLMgNX/largHswtDJFhSakq3Ys1dg9Odu3ZAMitBEqln
tr5kleNmxqKQG37lif682hSnLKj29ezlktRfLsHPi1se/4LicLnxh9nyBwKV0mGa
9riSpwbKDwJxWFZEcL2ZoRjySnaRdm0dlIaqO6qwMsOyjUafcZXv/S2zg4Y21nLn
UXXHR8KOl5YxNAd5aMIuAaDIRs4oKomdkoL69SYiwNX59UXc1ZUh7FFWIS1mHVKL
bN8EYP9yAfOQJw/BDHmfZhtTWlmuCHG9XrCsZSbypJDxPA9ICiK3F0DpI1zjtIdF
x5IwRm+qwbqukUejTVAogd5n2z6uzi/P1mw1oEK3KtgOIEJmi2/Oa1xV4YD1qfT5
eZ3vTmK2eXsD4S9sePhmORSToPfdbkZsVPe8VrHirRmnelsLgQIautXAf+yVpyyl
ACAJKjYgg3h8eWwXs0sqRRChvoVPq1xoLq2pDXWVdOeOQwpQgd/K0AsVSFA8XAvI
X/pTLZS5eOCtO5gATdbuzcYxI374ziQAPmHnrF+rZLtIClF4TIQmyB35yJG5dRfH
Orz7E60xlIqVFHzZvgAU67/3S2WDifULKU8lPzDhtOBp3j2mP20d5RM+YoCgb4d/
ZyvmNeFaMn084YfnDcxqFWgeI64o/h2Sdx1QT/nvor7CSAFAvt7DN9gzxbmX39Ar
TfgQWzNct6DJc9w+NZJbQcPXT+CqXfv/QPzTE6whrw8/XN99b1acq68TedjH5vo1
F2TRAuduQ3Q58HgzWZKw2uMSuU9kq9XgPv8R+99d190sbcVnBygot1LVTEO35lu7
YRBgBLSUACDRvCAeCIdmxgGENud9Vu/TgklY7YlOdCOGZsNC2CiUtVjZhGELhMYy
+HBAnbHAIfO9zN45T5orGuP0u6YVU/MQuqY3r926LLiA+n+XQO7EitVM8ql+UGIz
piVSrIzn2P4UAHOA0nBfdL2OzwjppLdQrfyVKZJ5cm7Dft9qex0/Y+IdiQNY3BU1
YZskU7OKcTVDVBQQrIfn2dn6Brv4NMJtOpcFMq8g3iJ8PKM23tX2Jhbth7i03KMi
jAQzWFEZ/Sb7PO+zNDLqatQkMjumfFG/0LaiqHJvkOSbC+LiWbaWvS0FnpuDaofx
ZystxmmNhcdezUeo2mZtcyL6kKQGXwUqx2rj4jIBAtH0yi4y8piy97+FqsernmT5
YTdDFVTmF8D4D7PiJdpStC/65qSeVtsapDv7UiHXUvszmh9bbBWAaVG1lJh1rgqk
u7a8QEsvIMI+9cIEFyOm/l7KnkHncRTgQ5PsPyR1tNfj0K7XNBkoxp7nz/GV/QPm
PXQLimfNQWpgU2x/N1nEdHNUEUkOluaqKT3QWDOi12Br017rgTSBr8W9yAH6aUfN
HHVC4DcAOqbRjYTLrotLHkroY+96E3iJt0rSlNA70VRyIHN7lEloY82RlzN6NBlp
5djyAjjPYAKqee2VUdISNJIPKtpZ/Ha6juu4BZxD2qFRCwlMO9egCWEH/rz0CmWG
SZmNv4TCWLxAwEkVMO6ZTxMkOP/0Tjzw2xIrhko0ouH0SC317HsVGQwvulzI+5AR
SLSyvydgIwYfBkCUFMP5CY8Rqu96dAZcQadjL3resBukmT6hoiq+4Ng1EwzKAlxX
aBqtT61tQff5w8/HBOm4gj+DFbdxZ+UP0c7jt0R/8Om8mGWHWh3hMZKpqwc2FnYd
ZgZK1qRGx1pQj42Z8bVbc2YPR533RaRrqG5HhZ4EZuRZM6unrbJbzPHV3bW+oqP9
K7oZ4btcTcknwgjSyfgRXx+YlGccEl8LctBlKBpg5YWx64ezAZJN13bwPBopwJxX
4QDczvyur9XkMhwMKedUxBKydPgBFLyLzpQmj8yiTbr6MuHH9Tc5Ug1CARbKgOYG
KclPcZF1Y0Tnk23POs0/tVUicflCTWtPekmWTyinS1lPett3Qti5BsCAEy27S+ig
zS2q4AOvXoHwi+s/B5XSc4wmpN/qjg+0Yg04PX22240Ny7wWPM8ntxPODcIxPLdx
drp5qdQWA5x6PeswHurdtou+1BIOjupaC8E6EixKPuzVbdhhcsKYr6rXvKgkKTnV
F5ndb8eLY+nZUaDIT4/1dWM3XYyouUG73sDE7Vi8b5YYz6tFSz8ky1o2wVV+MpwU
bZk8z0aDCqj3NNdfZ2/mnNRzlZLs6u9/Sfea0IXIbcaGGfiFFPO52stc9gvNgrpY
OK+qEZ4/rdeYmuwxjYd4/ue6nVOh09g898ppJ+8M7l5AO4lHK4gw+9Yj03DqVjzN
O1lQMvAEdK0IrrDVEQWUBW2tO8tF948G+McQYWO7BNsCUyr3EiKzqHQPVhilTHrk
dGS3GKs6T5wcvuCskC+0vZUL//d7NsoIocZmbDfBB140z1VHJbRZgXXSYSb9ZgOC
GJoGXGrjL0efDvbdbiBytlvsMY08HbaVPLAfTenIKu7ehDszvT9WqoQDER2ifhvQ
J/vA/6KTtytuSYU42FWChJppk/mSp0fKb68Us6KF5ubDQRJgLKH6lYWCP/euIzXc
GtiwD3nVMiMMVpRbMtpviKS0e1K7ySMRn23HL1ClZzx+Y5jMqfLd3KTXZ8tMLh6w
KnHk3imp/4litf+OY6evpwdp+Eo4Yj+DuAeQhOzMclxp2G4mpMXAG2lnFYNk4DAB
iyBdYGGon1UaH3iICeb9mG6GnT/FjJgo9jR6UyRqmQvXmNNIIgOd7EEml8tfkI3+
5r99NpvND43o+VUAGLVuWN/tfoorZwCMSTTDiPCHAzlncqRSkGwNfzOdh30gBdVy
uKTOmygJKhIn3GPym63Hrh1eMMUpaE8l6ya+MnKERBO9ySZCcycRqPeYWlzDkl2n
vkQ6MEh90ro2Y7YFOu86jhGbdG3ap75EW6McGNZq7vGWJQYBgMr0HrCeVs+x2Bb0
iEUPqjWmJDAkXJagdFLJGGyzhe33hWHa+Q8yEPWS+HNcm4/uTJeEFrH+nSv9G0hA
l7XqQhWK7FNokatUtfsQS7QO4h1iK5GL2dSwqZp4hvWC9Epu0UQpK18E7C0mfpcC
NdWWGgGV6kvhPQD10uiDYM0XQRrzqxwYCq6n1/wdGNEGCMYtUshv4+UD6Vmph9zv
Txhw8lbK/TmFRbBzCCXLzbv1jIH0r//hV13PiXcBg+Rbqe3pefZpcNt39/ONo2Wn
a1UYWPWbtMeQgsyuRsGrCLSHLzw2qg4+619yzYzVklOEyIlQPn90kZicoYAak0xx
TlSnGRHu17u16Z7cniAQg+Cj7cpF1GhTOI2crW3TYpv4DBp/jjvVkv84ERWZK9YJ
flxaxJd4bB3LjPxYKWoWjNZxp4PeVC4IufgLwZ2lcbMtQ39SIjiOpvoQ8YoqQ+oX
ghOTGGzXWpt7sFdk1al8zQpU1zSYnVJYlQyMVQe5qAvZeD3pv3/o/VHg7UdtRj2u
gRpUAAD94zVkouOw/xKj2xOpu7A3CI1EPcSVvKSZLHZWp0TA2GTExswEmGiFcHH0
cKIGgk5OfFjq2EdQkpA7y9wHYom/5Ik/REXEEYwwExrXNMO8lXY+Rs0b6XjJjzQs
6WH7Vtt6oe/2fBh0IwqodtihjjQ3FqmwE7phezcZVMS16NNuRX4+gzDWxL4bOXJR
mmooSgqhqT00OmnNoYntFF3i0R7QW+PVQWhTC0IlaNJ6mz2YCUPhzd0o6dX9SMkZ
km7QMV8qJTiekxGGX9GJLgZtJKaS4TKYDkmcaippwYtzeVyD6TqUGi/rhQhMT8YG
8bEUvyAwWGk07Dh00BJDA5EkjlaRoo5ukji/5YWnqEc3/NKYkhPKbiyoRIr35B4R
TmYMG8muHjoJ5EZ5TO0pnb5kq+SV9PO6Ub+m807nWFTPFWfpQeYOxCyNI9buJIZe
3hDqD6vrX5vHmn0tQ1mewYsJ9v1OOZehlinJv6yX8qkfUKp/NMt6bVdRfBnWI4He
QejSG7PJkLcU0Wg4Uo6hrSbAtzSGhuIMvE/+H8xmQBXoOXzUKMIda0H7guGIBGUZ
7g+zKrhuQ3e/2RWCZcHkdCxqWP/Xm0PutIcxd42PwNgMANi5HsxVyt2Dg9rtNgKQ
97gqUw3LrnSn6WFURwfjljo6DzlcZS8sICqf0XQ3n7jK8koOIfliYY4/rtPQBTQs
pJnymiem7fl5OwkXS67AxcD6sDXgJQEaBhMPp+kWi+o/YmjRShm1xZ2DebWkdNdf
AFWGCMumaYvtk4y0sqR2M4UH65Xt0ZD6xwOjUK57HwdApkrnJ0hDGUosopnJDnPG
gazehar9gxAxz8Mjm5dUxRGR1NJtVeu7nZX1pWU5FJKitixI1sQMLmV+gFbZ9ob4
Cnnl1HOraeSjc/2nV9G3Ht//zM3uBlNgWvrGD0BFgWfFgqz0uheFFsQLWSL3GIz1
IfGaaxfGAGt4q9Mb3FyJQl0J+KCAqvAbThDglRZ72r0ZOyUSVBgZ0V5OmctjCN6d
GBFo0bH6lBfTU3aiQEml7AUL9MlG2KN+Q4sU99WE7TW1lDNQ1lPaCABWH0ADmDBe
kF1UdnPGWQtniwF8mJXAxW9znW8/WOivajbmUMjPGfQHZ1lvFj3ebp25P0G5qpCE
PGSnY6T2ql2Q2hYOIPfnlvUwsgD+Oh9epG3JQ2djkjWx40itUqnm6gU5PlefsNwj
/EgFW/Oic6AGExJGdM0Ftm+A/9DuOr5kXseFxFPz5F6iXobpMdoPHv4Cjqw1pnbJ
u3BaHDMPbbpMm9Uz7Xc8PGa668k38tUfSfPXmZjPoyTSX6oEaibgLdMvCEM/RZWU
Ccrde7qLvJWZ50lsJrWoVHqMKAqg6wHkbIwUmg9q6OIJAsjaRuquPozctJEqHSB7
RamHtl1MGwmMvrROinhGkp8rmIkKBEXsbkgUnMuQcuk4h5gMT/Jp17bwB5H+G4jY
8TfCZqgvnhL5+9GYejPOnpBiDlQjhB6b4tEtuR6H0v/kUinLg97ywuINBsjC/mm2
27KPbPTs2UJSCoUMeyvHBHOWLMAJ4TsIpjGDGpIMgo0+AonIcLBkYH8k42dZEmdE
9/0ry0/T7zkmrxqzqw6R/UKl9aaFhGGWo4+xn1J/CPrI9BzM5dEy6nBSYZQVVeIM
LJ4j+bsvd7TxMV7Yb4EndgFMJFdKOkfiRizh/tJ3/6dvdPCWJKhu+mlSE5zyOQSJ
aALxGhYBNMsaePRIlvkYFb6jylQuR210CxLckoz0d5VoXJkBAueFgHJzBfpY3nQm
La4NL4Os8D8Igz00AseMUV/zSeSw689bkDmlO+QtVxGYvVTn4Z/5EU+gV1ahFCsI
6ZfZsV0Il1L/f6KydtvrjofoSCcJ9ni+kb04zRlCmUYQmtLCPljViULShcjpvYej
OpNJlm0gakR3nDWnR5/9GsGXa7dUb2BghXgqG6SxRhnF77ouk4UM5IizXJ7vi8p8
39xEcg5sX5uuQqDuzitOBA5cvKMKkrCa5xZp8HFsGi9HOvVY4FaLFwi7bRI6XEFJ
PCTXU59CKmttSr+FB7RXsW//lGU6Y+QcApEDhEk1nqxSrhjoggIhTBRSnni1MF0Z
61G0hBEteRxEd2/p+R2+EmhNViSivKtdpAWrU+2cflu7+7Lr+CEYAtr/tn8FMhCY
F6/epMby5r2WFVp9hPBpTjD0bplYJ6XFtmuFSVBQh8rWCr4wW5d1c/yipgzbcQ4C
1uRweMsPo4+hs8Nkp1pCkOACDXRkmLlLoAAh0n8MM4lngudwiRRca/LTQNCdG5kC
MXgFJrPud8BVEsGx6kFfIHfCWEGsZCg0ZdpUqA/KDYaW1SmJqUbvcOoabWUHDtji
uKvgpSWqUu/Ue72V6PcrjUC52XaCgKQ7f/tIJWYxoTr2aVode9NaDc11iY2eYHlO
SnyUFMpNdrTlZH4ra/rlx8xayMVRSxq6Nfe/8HGQbs+UF+tgolZrxhnZT8AaJTaM
Ceg9eyNaB2GkefYJq4yAl52Z8QicaTQEcBQryx8zdfXDyBnGExulafIuGJy3Hyzy
j7oO4U2e8I31ftwNZDxFsBPDjt9jgk8pdhwAQ8z8x5/zE2B7gGWOaX7E72HpH9pc
VQDwV1hAKDZH2Mbv+vjJBe7HHt8UgrACSUtQXWhXFH59HBgf6MIni/2ECz2PK5Xh
3wKWRs4AeQGTWZ6YsHeSwMO3acliCoqxe63WZUcCCWeu8G/Nc9ukbWqJ5HL4pGCg
2J7JRz5Xvul3L/fctuzTXmolRKOTUIqShdEAuOglCvIKifXHpbPrvk+aagmI4hiP
V2MySejgBh9akdqUY/dFGIJkKb21Co+03Rw8yPaI5m50fL39e4PlD63adxU3oFtT
QbhSoVHQZLJ7roiMoNY/6mBuAo3UWl1CkpQyF/EpSpwZogW25b7JupF5Q+s+YN/7
jRIzZWbe2i7xoS672yKLzMM8AJYctePsaJhOMv/GrNdv+ql16PEfUwP0RtLZaIpm
m43OwkTBrNbmoz3+C3jtJOcxxV/yTNF9MEeYog4pFo0czqVoxHrB35D/IaBa4Fjz
A80YkNQViYjL+8XOH3aSX4MtzHbaemfMXY+D7xktKRmwwKGP/wnBh+jYW+dvkBTr
EQNMVgWgZ2THs5JO7EdLexmFXjqSKPzrJ97/c9PtK975Sq6KcMmu5iZhMXumcioU
wARsQ5UOfEdInGc0lJskkTDLZp08l3HEosjV7eCnrzgxMaRMPl1LkwJsVgqw0vrq
NeODOjolyrGh9J2/mL3KOwOTSYqnOtA5EgtlkMdlHvuC5X3ua0FYIHdHz/8kVBbz
UdVrdUzKPDmQV2CfDFVMCtBIXpea8Op/9KcHcRUX7UpT66cwZnwAwNtBcTrhyWhd
U3PNuI2FEyNpiuIsaX3SzlnCON5E8yzKpRIqP36eGpx4Xx6sWztgQ9+qpIG50tOL
vnQFYgewO3NL8iJuhiNOxdI9fHl6XmRGsF0dNsIRD1zEow7RIP5Dh0pqhYu1t3ho
Z7k6HqQGKONrhUWz3vsv+R7BV2tTkQ9qClgnq4usY0xi0HMp72vFMU5zK4Fwks7L
RxhS8mi03lDvWUZYh4b/vIG+a1uIm1iQF9UWqlsoUf0umpHqeaPuGp3WscK0g/vF
UU408OaW5Y9tJVJ8WsahfIeLxsVWSiD3rjYovDVSkynDV7aYlxDlq1yHs/VfmDZq
S+PlK9NHif7eiySDLmF75bEEff1QtyyJNO46ZaAbDt0ZUKIIB1Nyk+fyw5nGLKxA
HrNsBC82iSadnIepFMhFuur0hcN/BriX1UZFMM5R5iL/WOO5NmJbrpPsp8F+J+vh
GkX10pjhs/dWEXuC/uQEFDxkCS0cZOq7gPQikbWSjLsGdjlPCpm4uDaa+Jx1vB9d
UHoCi7RvM+16+pTDwHdHgEGXl3HA3WaKZhNgX98rY3Ht+3X3a0PKva1C7uNbrU5G
kgbGM+ChdiSng3zUUZqUH8A8LJce5DIK7mTDUh95j4blAFfU10IHfWatg6lzfj65
vaQsOeJ4a7wAibw0rbVmaoJx42+u2fpfT25Y9jAmtSN11EVmhpAlh4B+pVT3qEhY
eBGDsetE1jdru1ubN3MCa49LMHafnOc1YS3Z2fyCN4z23ccAgClLd9T5PEsGj8+D
CVIMRAnzjrDZKxHIJMJ4rMij756kzXXyUVyAoeeS3glfF0G/rgApNoq85zX+uG/L
MbhLRV/Cc+sr7yrvMp1sIf7cUwmJlN9VfxDybq9+PdU1WAj4jolXRtWxRDCdqaqh
M+Vb3KWbB/PVL6aOiAqkkg+wgk7VnOaiEAEGSIjxtxvgIh0TwsHOtNB5VCv/LrCc
0f0qhnyTu9TRE2MGW9ySPQ1VFarjdi2cy0EhIivmnRLq0otl1T7i+c4SGn5J+HE4
WPXcv0SLiVmiEJByjpxmxrD+MAPBKmulc/d97iogu/0hVPbm0WOFca8PS6oYTzUo
F1Nuxx+iIPaqzdip82LC/3M3SNHasNAPQ834n1x5WV2szt8pK9V5wbbm6OwfFA3B
UrPbdeItew1LQf/v3mBLfxlEldrVQH3DvBFNJNpszhYelOyuiMw4IO939GbTTyF7
l0hM7bEVMAH82DMCtJeA9bA6YYx6Ofw3OoH/cVyC3COa+0p/m3hs96kifTPzINTQ
6ti20ynCF1Sk/Pq/Ctrxi8pya+6QOB1frYWbtQyhGHHMf3Bsyceb5R894KMYzvzX
nFqqWL439mKCs9fFhP1ar/mvMCYdR9NJWi/6niZpokHtgLSjZulmicJJCL52AkDz
s/Acs5KqHe8h4a+raSC0uRGwjqn6I7waF0oWpheRJAIPSY3pFuo24BZUHQoKTlkT
EuRDjHKn/aVSmhipMixliliDbgLr4UF5hK9zhHmEgZ4L+BMCae5kWbz7kfj496cJ
yfiGnkVWqVr+WS5FlX6AYoR1PksQUysvRWmGIU/Mm0asciRk1WYgDOJZQohKjzlX
LnE9nR63c2eqYMpCzh3hggVldeRx20ECm6MTEvncEzkYReKu03HinbzEZrtXxbZi
uR1LotTVfT63esv2BZchnPGmWIJ+j/TR8koQCqpQOL6M7EOycb3xuQt9PkvL0wz3
S8c2B+Y7qSQMl08xQjOSUSpizh5JzvpnKl49iLbZ3957PN7ZfkUgLZV8V51BFUoT
h8UBOAG0rr2p3Uc6ZO/lqCBjAOPkULuTBY+t5KHJ6/AzDRi5E+orAlt4yBzrnbzO
19cNLQBEszWm8AcdgPPVRaN0ka4zpfPqsnlZFrIIxb5q3JPFv7EZElwWyvx7/Oht
w8XPvwg0w5Qrd1av/ecNcg99uy6Y5KCFze9qgRggqoqwqDKvpiOuWilzRq4SPNCT
vktajZmrKW/2QjtGQ8N9DK9sx8qSND6Tx0R3gvy5L+0xmlPSSxwd/4ul8nDSr4Hx
Hd4/7w3+bW6+USxpPy44GvG65EbfCXOg0yebOkgEefvE4F1/fjxfcGEJnxJDz2ti
7/+b2c0xwzRi/3Hnabb11Tn8XWpvGReVuW5a9EBv2fDwpRoqlyYd8DlZ5fGpnD7X
QO3PdD0Ff9U4O8hYgVJaYDrqUDNB5TnetE9uU7OeA91+lndvwreaf7i0pJAv2M8+
IdGgMdVmLuCJic0tNwHfZcEpKglyMmJwLhiboH4nQOR1G/RXrOjUPTUk3+kgyaOj
UAopChDSn3x2PFUJ4mIrCHIp7wy51mVYjWi0MNuFsfalJO0k7qLrZQO8wASWIwmg
Z4/sKSADo5mfNIOSZB7dukQzZq0vmWWdT+Cin2pPu8cm9OzI2TLkQnjpPrw2Vfvx
Cv2gAgiNPBYrYJiRF5BJnRhPd+uP9SGxqA1alg3U7RGZg/iNhGEb0xc2eycQ0nD5
+Glv7l48Lh1CoPv149czizLsF34K7nqLmTgCN7lJwCHQt/xpEyYPdVbqc2SDP0Cg
LfvusGQi5gZ+BKk4xkPJsr5nbGNe3QsNS+PbQ5NyK0iPWriNDq/EqcESalwCs4ED
2PEz62nHwH8jjQCyCq5tiRajak1pbXJL7HjvFVBBwGc4/Z8qpnqSN8784eyVwoEw
erMcyOvUxADMjb2yALi2EtjZfEScAgwDSMbfvAQkEurwWAcWzzKkjpK8pKbBMeKF
dDkMhCRzcvT1I8g0qRxATyFOWuzScGiZ+ctTJiUosmVk7x6/1m/YLP/TNZAJIonU
dzTNVYzBeU63YjTWYVGeV6xT5SoDC9hYXmjFZXbqNKwFVyr7MUjfygfipyTXhGmh
hBPkvEnqU4Q9IMMT8TotOYAzZFJN0KEOgoCdlzpeq+qKkkBtuVLzMUpYf+EJRmAN
MVAYD58xxVMq+pQwVfq53ZGaHuY7CfbtJfWBr2rFoZYOVhXkwGgaWALnQaRMuCIM
IzBgujEBKFEZfupYu8n82PjqvQf1piTgih3ZmqSHJPLi3+ZMNl74x93yjkndOFd4
dOSXqyb7rTjHAltV1lph6BYrPeaYdA5gtGu7GyIBm+wPB50lkkcbhHmXM9xhfjtC
5GEstqiRlZIZGxVyIwq1rRdZ9wPztwosg6MPrA8z0mx/bpZ+0ThU36C/Ci6UZhJU
X+BP6C8GNSAO2bNcWWPBl19O0fuWAmQqZpkNOmgO7OJYlqhwxcG+8LJTYlg8C6pe
SFE++hDypXa7Ej9SZemqDDz53mOhc12YO0LSTZZ6KmWeQ/d2TMT/GqxIutTmBWKL
AM8i5s2Ddh/oobcbBVqeclw2O+n2g8Y4rWcWKnvvtFQcoTZgJgfAzGKsDxKfsKij
kFGFTB8HSm6LyG4oE6txElajFSdKsTpLvSp4jXepwWp/Hn1CfcA5/UK/DrdqhcEg
b8cTMsW6BDTpFBgXZv8qcI7yQTyJzJCosFXjPzR+cWamwNbcfR2MgT9LSlJHi0YE
2G0J67Lk6OTmrimVzuw0J+kS4SGj50mxon3BbnVPePU69x5XYO4eXZKA0qbGtFTm
H/IeqAR3HGvtC1OCKDa2oFrrOjt1SNw8My4bwPuMmkYNOF4c/z6OD8IQvNiHzIco
Nfm0ev2KspipW1oWM2z+aY05aLmzR/tR71fJAaEtmtY4M2gwBR7gmDLEbuC6TWTh
DvKB+ESfJi8nkrKcZdPY3rCtYm6zQKOFcL6enUSKCR/WS3r3p5AMxqvqd5P7NPhi
SUtbb1YVUY00M2GEZeTRQzQOJOlT/qy6TSkTMQnU+M1z9ObWg3w36iVBHvxmJaah
ygSO9O+4nH5l1opHI34NiYJS6DZSfqxWYgLKW/M/6yOsgYkX+JCue4WZXtQK12mU
zHnFnHsvNKbY8lulMiuU+Eg2sYLQXr4XL+gx3/8+7VrLnYMEyjwSJ0QMMv1nw8vS
pHbQiYhYm6O+1N9lBceTWS4JNGpkBtiXKuJUKLqNvPI+44mlZd9nbs39V6o6qPLy
wd7u4LW8zO6OaXkqZ2VAYlco1l8Acjbo+T7CIG5pecwHdMOGQhkia6SQDkMdLk4J
Z48UsrpS9ejaXdp9vF2B04UVF0lkfQUExK/gCi+T5GTpkG1l2YnEQfSNlcvZDWwx
lgVGS8aQyz6i1al/NAXqQMsCq32+bxhBGi3+qvhUccg7vwAV02jT1biX6GhgDpd4
9vqBCGEIwxd08w9Mn0I2sE1WzYw3Sx4l970DS8LEj0fdeMKql8PkR3AUiquqXej3
7MkEZQ5EMJ7VHnl6c7duGjSs9lp+GqWyjIU/eJQaZHKlVW8ZzF+cGr724oCT+Z/l
VAgCTtoVoTkUGk7XXJewkKxMpi2jbAA6c7a6aXE/7d3mLheF2+IyOoCLyQHXipcU
3jjGWe0Yd3f4OpeCEjgebrBrozQqJoKYX/1mYMx2MdVFAUGxe4c2aoX4PEaXugu+
5lgLf/h4yZqqRwMxi9vhk0h058IoMI3x67pWCi2ocakp0kDGxpVGqkIl/9jJyk5E
nf9pY5ex9byaEBU+9ET4F3ueKTik5XEAvd4OMSfw/+guvCXZsEODmOzSrcFmArR0
jXrHVYT8qXt6qHHtxLio+Ngav3FfrhbV/oDlCbvmS8xdctlZaKD/TMfX9LwzbikT
cYy6q0g4/w9rAzI4HLhhX/PB8SIRbfK0/rvNl1b5lif16sKe0b2lsjY8eB+XRkd3
Yd68ewi9Rn5Ejqn/6zjVbrptyiMhQ1GBLVX3u63Hgyt9KzT1ZHQAzmYKA0KQj8dr
/7l0MaDnR7korT5eLB1aqi7niEtEsfh/2lhVilD9y9MX/IE5SeJi3F1w6YBBzfGx
mxl6rAmV3QAm//iCEDJjjWdGOrQqllilGnuLe99xiibaaHRmrQ+/G1//M/BRJN9F
aFMC/K1GETG3YJxi8RHEuhdJ2ZkJjy1Aomk4ihTRXfJSbuWVYxAe2eA7r9IMzSI7
suHFo5CoB8DFCpRGwUho1BFYhbH+8allKxxgAeV1CqUfW+lC6z+tjSqgeUiuae4W
AF50/IGA8wA5bbcRXaDyb0227nMp9I59ABTlkcyCtdF7uWF7XX8srOKCvBOlEtyN
NoKgbAcV62KuB03eDpdQ2zt0+wqxAhOZeqmZbnv0cVuQqO54szMPqEj+R1HarKNb
HRV4FMuvKBVhEkWJmgkLoSA7qaWKjwzPvu6BmkFN9rxhIxb5O7zbRbsPBNudHh5i
w0Ar9GQnx283+s4dn8vYG+doqEogkL78I6/p06Bf2Uafej82m+E81kl5PfUQwnZx
QlmUlTGZxc2IBZvQ8QKIcAusdbkE1B1uwwklV9DSdfBQocsCejTTVXfyrIvIE4Fa
Zgw0ftxVFOYBbSBn4EijohkPa1FLgn/xQwGWakaALHeE6Fsmd7GBjmZPj6fFfUZW
2BiyThPKgBGdDneBRKWAIQ5d8A5MrOpwaC+rnJrSrxu6DEyCGBKLfhoLuksy3Lio
dvQGzIHVK6w4SxOqIYvFDFHWELBVSMfc75bTuuI+KKXSxF65y99+pMaL8yAdA8la
d/zRzD1B7ZcKulfqT9yYFqW0fSaCjBmanRswRFDoviYXL/KO4eNJIK28aL25v8PL
TDxfgjv1oq9mIgGmQ/eBpxagWHehJYDrAGIbHqiLIIvi/kQeYILCxG+hYPfeD46x
iC1vyP2dTBy2YsEJLzHMa6s77oggGvlA96xEu3tozkUHCvYHUodCIzhHKMy73XBR
Eu5GQmOurmMXCklyltQBzLTm/LJ1CCzAEM+hsb6qN6w5rDG1hwT8sdcn8AmMAQCP
E2KPlrg5q1DfaaiSPmyYA2zGsU6faldeHi9AqvHVgfPillWr63awzL6RcNhsdETN
TcNmFgGz3+9MQIjyy5vTMWHGbbiYboQ+KOW8PhOSGBow2myRv1xwjna7loh0sY2G
VnNWIpuICGjozH6BFGi69MifyhI4ABrqbrRlM9MXpTWXd0snIADKxpY2aOHTW8ho
oHnZwIR4uVyJUSmkx6y4+ZZQmhU3oyq9lrGEGQ+YCozUFvcGVWu8wY/OQ30Bna1x
9gKjkE/3iKF9lZ21uzEnSrFGGauuylzg1VcAAAHxpZgRJHp23WDNmj4m6j9X+1eN
QP1KIZ4jwWuwgzbKqwwX6HvO95oWzY5i4Ppmo31uWVORuWdR1dNhweYxaDU5pRDy
yf2yoYdmPbGjEXsOFEFzZpUOCd1/t+Rps7FayaisTiAYT3Tg5vbPxgb6Pdk6IKjF
dflkQ+k3hY768r8a23GjlL+6zwOJCa/xiD/AmeDMTQMAvdduwP8+FzzanDuStvLA
VIhYd6A3C6Rnea+xgsk5bMWS/37O6sheCVn5Jla7wPfSf1cy0GqbO6HWhgOXR0pd
YXo8AGOYa1ISPgBToFDPQ1WvSf80cylWk+Ap+3s6ook7EuXF31WIV+f2a9fuHssj
fTptA5sNvhvxGAh8ddPH8iTglSvGiU4dpT6E280Du1FlBGRZuwb7q557gzCLqfEL
RfmsqbQF2XavrLNi/0EzdYe30UIu8kIUu22PtS/nlQPmosQy4aYHu7vWOxSft33L
0eeDcZc9WBGH8B6ZhuxIzccanVII3Lnl+FGZCy4uHz/ecp1U+xhKvq9kKo5HwjV7
WxNj7nO7Qh8KaXLqOoIKRK5bSxCGo/ramoCvynCDpAwvVgzvfSZRz1XixPrx3z8m
KdtwIpXvfcvxCJ67+p6Ugrtxd2E2GQd5CDY8rXxA9h2ktDO3DgT8rJmby8vZ/cJV
chxDQunX5R5mdwA2BVf1KgzL13ib/c7RXh5Qk3FrUuCb+GaWGxxlQLuo339f9Ofi
WHgarwQQ1wNaNIrRT/GKRGLCBuxdMsYEeq0JH7SO647aCPFlrkJBbTHGx28P7YeH
wLSOXDMg5+U7+EADdxfdcDd1KoulJaqPJgJDuYLCKTprdu05PvtQGjGa34bSp2q5
17V8iRmhHE+lkvFgmp4lgIHSdtsEPKW8P9ROEjQhfxLzI1c2Q6Q5RrHT8BbbV5LY
gdNpBzMs8F8tj/2H79ng9SLlXLUw76IDM7zGFAhAw9EEsqNPHR3A0LUbCspLPuUx
Sl3TFxNb8uOqsAG1nAuN0o8hXybAivTUY/Dmhi+rgHjg/nGTTWTAyFIqThegzbx5
XFQzzaD58N+CKTMCmx95RnuqbvVN7eG2Gu/UkNjE573rZ4BYsDzEiwTqPU2n+meh
C94ksr2+jGBvAxWANNBP8dbGs71JSrDsc2gbbwSP59EcYHuvOwnioSyysSrFDdPx
k6Nk4RdXUj8p4WwkWG6J7fZZICq6WoOBQjCSXdSvgJoN4QJuDxNJIeGf8TZBivEC
BmANMoXeFKaFWZeBS/n2/bLwIimhdWOvM1RHldctPOU3j3Ljw2x+J8TvoqzbTtsl
SK91qxXk+ovTWLcSAfKMDD1G+tFlmmQrGvYiaGDzG1MUG3tia6d2tBIb0GxyX9zU
p74UiCJs6LQ0mYIT8Z7GpUz1gHyaR6a2c++4A5NdrPlgM5m6yGyO/uEZCGH5QmuJ
/Wkss3gtUC2oDMR4J7+sM1Csx1Af0NFjbEcrPyln5sVlIqUt3RKgvXb/JYbn8rtF
+iZg43CltKWbwQiiLAsTq8JGqWqLIfNXPSZaGwj+PlEpr9OxBEvLiDiZ5aft+gyJ
Kwkq7Dh3a12A4U4trH2p6mM10+FubT602Opw0TK1xGw4xBq/bisdXrSAxGZtkFMY
kGa9oB77aXZogz7JwcCJQKhPULQeBOaVx39ZilFpWNrX2t+a+Y6rZrdmyo/v6fwo
pi8rSDh8MVxdDxcSZxGPQh7fr2+pbXFBqiaHwZo+YpEQSr/nD+nQ/ibmu9+5la6D
0ShKszEdxnqystV0+vCow2s1dXvAI8ScDPj5Os59CZMIrh0HBeOlx/pG0BpjO/lw
z6TNqE85yJHlnoL0bqTKKQIjOos2ntEHoEwb0ZavGrwAtxBf130fx/d9thbiwVO+
Gk++bWnzrys2tpap1UoUkSNIvC2E9UEBnHeJL8Xp65/Ew5Z0H5Gte4bDiDtfwa44
2zm6VLLKpkGescnndCt1j41QtioFo+7/gXXjxVlBCy7gg5+U1X4cduZtjFu9GcP6
nhncFcTeOuP8W0836pkckK+2B9+iutG5ADopRfkAotU8fRd4zW8al9M8oUpoheTu
JQ5qu8Pi99EArIELl+c8fCWtWL1rJbqpAKSsanNoYForKFjE6Df5/gU1qn4vHN3N
3uWfbTJLvmE4AWJIvhzi+y2Fer1/1fL6KdcWH6l1WZzJKamA4llhY3MRE09+IxK0
/DRECiGAo7agJ6ivUgSYzB5RYZ8EOfA74DgINIE3s40iOofhQ+vV7mPMBGj+3ela
Ej2cU79EFmIDs1nUypGKwez+RcX9XovCdj5ww2+RxFyPCbpfDGueouHSjbw3LC27
6RSfVBi3cNMkAUivRvISy6LEgj2emgfEF/H1NZIGK3RRAEjrMUQtGO915Nc9sWot
dRyasSEe/m9ECWiP4q9gr9sZZzXcJ0i17jgsJmKpxELYTmR30k27Nh4SmcYrptBg
vCDXrjn6r9rCZmMyJF2cWXBQNLWqE78k7uHcCTXKmXdK7HjitPZA/M7vmDP6lo+9
knHhB9oNU2i4RvBD95rgxvdNgHshI7zr1/Ey2AQAbH0wNvBGAEuqb6K/FITdseU7
fW9/MBc6DlqO/TFqHO9rj2F++V6FHOxftcBrKim8lTFdmn7rMmfwzxZ1854STlGF
9clemAo+Hd2yKHdMWZqvdBwXqVG6lYv9UFVupBcFHdVXr6lW3HsaiR3KJ8gq+495
l28huDRu4Gt15jBiRJYf4KakJo5IY9mnRRnQOv2J+XA3BvFDLzTaG3/eCVkwGS+D
Ae+m9bjwugmDiPBRfW+L1IgleANGLibS+4/EvNb3Dejfu8pyYQrIO9QFpc4OjSfq
ZY0UmvnPfT/x+DJH7CkCXToJ+JemN842fkJqQhwjvQ9kwpgk5C2PCbW9sVwDNhKA
10EjqW3YiqjzZdrYAIc3zUq5SV3TUmMw2jyVJy4T2eUu/7TdK9f81MYrTgwGKhfa
GB49iJWmBppokkMjq6hiMgdiaNI7f+tNzWFGoFUeoi5kHpAUucSGP17h4Sh15ki3
1uTZlGXcMen8CkGRoRItOn4o7nUinXsZqWjOss+yltAImc61ZsX/A/3PEU2II5+S
gt6ts2UFdNBU0NyO4ZbwoAg7/eEVFqBh+8ya2kR96O2xSyccxEiKiS0agxHWCn9G
a1AEDPdhMpZKqQHHdUGg5y3Ignb8ehVnGIz3rlUIkDzKKE9K/dZ91biLGgs2ATQN
dAfNrfQGdtCxTI+flzMv5DfGa/qFSypBo77FbtIeLA1Y8Z77/PvtZiovnawuMkXf
HyF+27zQCLOu35Q9breRXfBQwqbVimlZNqrBjgLcc0tFNXlPwFCNQaVi/fB2bA96
gVJmWS7efhM3nQhlwoanQLjMSKGdNPUx1Nn0cozdHucJh320nOi/p1qhGAoRnItn
bNvijJXUkiafCLT5x21/fWRbnX4Dcc5mMXzbMwClGC/hQSsxWR2Oegz1au2GwYd/
NwTRBhB38kmjWLG334SeJ6KEWHIv8p72a1TdyCIWfhmCGn+upj/su8I3hcInqDTs
KEzHi0wquRVbrU6Fp64LH0ii7vhABVUf6z8Uhd46HQ3xn7AOuinHeYexkbyvJPhx
KASqYcVnhSAQqsPC37oZCoZ+iQX/wdeLkPHFXO3tOIng/1/F06CRS84RRRJ1oeGw
kr3YuZ1Vmx5O8r0zeHcGNvzpvpxgx07070VhFaAch3zpLcMGkg5fvlo3tyMPo9od
ARRr8V/YtVOQI2N7u42mS2dM/chFPxn+gS6rQ1YfNmegrnSiTKifZEvv8vNGBsNa
T9EX10+DuO3eKQaQnGV5hOs50JQfhopRbwUutEior59s0791RLPovVrKqtkFeaso
Gek0eO89xazU7M2Vx4WWkpVrnm8Sak3ZgIN1fnuxsnOeWGI47TR2Uo9RJd/JlL8R
gc2nhLB+jMMpBVdlqokJxILydqD1QdXwEUAh6JHDil9JeiGSh0OJlqj4JraTv0Nw
uLNqvhRH5Izhkgua2A2BcsvatPzWfRSAiZ2DFQKPucjmttcvSbXwN0OZZNxFHCWe
g/7ZDAiPmdFgLChkYfG0zJpx/LsYVm594rVAIOqG7RZR1KZvnM0GkXcWEdhacqXj
FdUvVxIskryjf15vDalhggizQ95s3BxfDsTpQdI0Ft5JSy7cfmaXN1qaVm2t66oo
7qgG2vKXHBnSaHofqXpPV3iOVNo6zl8zbM6US+1PDmVelm+4qS3bQIokbi49gKjm
VJz30S7g0fHH2roDUMXAQNzklAFWfDNeetwFQOI1iBmeScj3QUrVvI6OffGvWI3T
R7quYHK93wwUMVoSUnCR/Y8KN4/n63IY8V5tg8iD/7Zu+I8AqUaBzI9zXEVzcwyO
CNVBf5yCeD49YeJ/Ag1bb6lecP2a5ThkwvjHWxMyrSc8Y1CULofIDK9GqhMsZzsX
JHVEpXn2jPAMGTw2/aDQE4unC2lcPthneVpKicRhosXBdlcF7jr4R0XefiZ+Q8VJ
4C/czg69/UmU45ytTOwUKqr610CmnOKzeqNZWQNz0gl4rREDO0DD4Skii+Qe/EZ0
42Yh4GMANj1dZa5f+bkv6e0FHVT5auZ3Kj0QkefQPelY6SNtoNkDBesUzaRg0YLq
uuNGZ6xTFg3uHlu4l5bl72u5XbUZoY2tlghmNOPYTuxHxjiX0SA2WCOICJ+XC5Fn
9ThjzX08+csvtSRWJ3SsRh6YFa7kHra/mzjVAVfhp8GdTJmpUWQD+WF0ZQ6RqOyM
AhTGQvGXr1Q57MEmbDa0kVrk8kt3Yroo9lPaGSRBiEJCiz/zQVmiv17bC1LRrKSe
+VTUrPGZCRPQOPS1zumCv46OB5JW0Zh3C6xva3r31Re8UPlyCpRwxfE046gkAGWo
SHQLIbMRH0cat+eEm9SKxeTdRWp00rbUPvJDaiFuK1BwH6+maQr4kzKdY3FtJk2M
tHknR1b/VyRoasdN89iqK5TuBlAS/WUdP7xyRa+/cph63Su8+/7WO1l+bkENnEBM
yyunqD2djjNPMTetDDc3oN7SC8Ozkc9jPim9f9+SAbUZl3tzRr68gPvTVVvMON1C
t7Bbg7IEkmUdkaC+9KbM1yYxkh5HMVFvCjrYQ2qE/7x93znZQ0W6ctcKLVsalfxw
ndtvcgy1/bnpJlLq1Raoj99Nqcsylglerh88v++h9hJvz3g++iWiVs+bCld72o8R
ydQZ4f9xNpF5qkZCZsMk64jK6pGBpVtXV9bgTvWZebTyKwQXAe3CcSSxRsuxvXRc
S/GhnJqm669jkugvSuTid+GQXthE9YjKIuj8GIxtB0F+lhE4c1GHKVlEztQjfhH5
QV8FCDKLaznktT1JPtXP5FkKyVdH0rUAC9mYR3Tt7+08CstRfX0ohxut0uA+V2+p
ThZvK3aiFPVZCusIhc7MjCpIa+rIA+ibyPbzBUsd4H7cpTbV1MtNd824FUJzfhkY
XZ/zArp7nm6maOlKja2ZoeDB6fCn3weWkTIkfAmYbia5rpdMsXdQv10b7+Gwofdi
jRQ77n0wQ74tSZzD3jR40n1QKnvC9PWQOO8ET9Dqk27iMrEuXyC+R79GVHKCrf9V
yqpXmmXqz4eEDCBINyVEbIcBKvDoCBULfVYGvxmApbGRUwDNrG3Uff77Ww04JqWP
pkgUVg6gaHwUhR9BsX7Q9QH4pVWqxqW8C4wtehov/bfXcDYm1M+nHyX/UnBB2b4V
3ORotk/b3IxMHDehtNBisG072OCr5VGRJbY10/ArW42Y30TfKZswRVW5cRr5NPpd
znmE4gLp/fNMYiwMixX52NXsusOUnXCgiyNEk3b/eSV7RVuReua8pDy9bTnpIT+/
YoTcij57AnV58SmkTgB+VQGtIK36U9wNJ5IvP+pQHEVsDrZEj9kXTH1wW+H89mY9
2QC9VK/BX6FzkPBvM1f03fta2NDrB3jJ89Ko0DNRApnqMjTMGCFJ6cNtKJpEyvAq
xSe+gkF+uGfiqgdjuGgKsvDkK7hvRrGnoVWEIb4vI/5jKr2VsYoz/7lp4TTbCkxS
RfIyoYpIl4RQi8Teg6oH+6p0Xk84pI3P9+rnjEDM4ah3S/lgCYJHLQndoi/c8c6V
NyjIf90ITmGBOVfZDROZDDZvhFGDs6h0/moGyidbntHV1MCBipoUskV+rOzJ1NPI
SXfG6erl0ipWL86Ma6NHHj3Os/IxHcdTYHeHOa7DWupYTxNYc4/XYvOT3OvFr2Oy
vSXnDlM32dkVoshYF/KLgApQ+XOwNZO8TvoepRnjTJrKSuEs+CU6HrrVX2TGvYEg
v22sGavMlW9mSZbQXcUoZuHdJep3GLJpZQ0BLk3MGAxEm+pnzEGfY8kTOm5LlsvN
j604XvQrAilvZHpgTWoE7aX4Wm/ljPU/D0dGaezrx/2OkVeHJCIkoakc4WV+6ncc
tV9CxEs3vBJJdhvjt0s+UNYYfmhnSrdDC95XhEP7G8rwXYbm8TXMeAkjvSfRBkxY
mOOGGSqatR1Ujb8gvmmk/o3dOoFMJGvVRp1BNgh8loZU9ECi30BxHLdwEl8+cl65
3sfMxgX8giSMJ59s5c9luHXMdlLjp5RxsvV7nY9RmzWdabOW2L7o/intdhsK0knK
8dQBeG77kHgK9m8+ae0xv/DRirWC6Qajjs1DMsIS5Hi/RgRGJnjp6fD+A9Zl1iTO
yCp4gOlsi+kYX7MzqcidiHmJmgQTsiTPDMF1FVBrTd35gmV8PbgxSkiMtoMMPOGG
+B0y2QPZK4P+qjg13g7SiTDcoKqsPrUFD79CtEtU6/z5eNYiuxCH+VVsShnZUcYo
7pYG3e4tjIYBPa9MRRwit4xhHnDWFaZnvkMzTH2VyQDlLZJXGId6xlBpuq3QtAs2
BzX7kjanxgQWLjcKnd8T8OPx2VSVItfZdLrrVCveeEqNfhBY4ukXzPG9K+OZHhEQ
Q4YZpE3zcZGiMwVczOdlPEpnILoCSYFM9fDEagrH3ARKYTQWl4OPlaVWGFyLpZxy
kiQ79Ir8ibCpDrz5nWLBj3nWW8uUAGdPT7S2290/lIjsZI23DSqasLhb4bAkybeI
tPNxgv47g1LgP+5jGBtmgFfb2m5oCSgRYkTwvYtTaoSiYQ4Zfw7bJTqTfApXon18
zVOkgs//9cfiVwEWsNgg44yLhxa0camEN976NhQXJZLt8M4fzWgNQ7yDtzHfhZWk
/DFkgdgn4GHq93BLw1EJDnvjrzgfFXqBuVuSxKpMo3iUT9Ns2UxHeLiF0W6tEkTa
kC/kQ8e3odFpwZVkGZRMybbwnB9ElxVE2SWKoVV28LaMdIZqYRlNS6YPAIU7YhM7
w4uYgRzB6LoZFt1JplqnwqNgSI34xQsFqqmhUGzFBwEsW/YxJJv8eVCI/M4zQsK1
ulTEjLh6luSwzHk30J0HKvUVcomrk1Koo8AqO9nrE4+eSFQj5S6ACH4QeipQ39OU
kUYlSHQRYzMrCYmglJsKDAlealhlu0S3GWyavCqJClgUBzZOQdhbvoNTmYoPuXHn
HJnVUI34+Yi/pwAHzQ45lYtZTsRTJcIz2hC0xN44MmHpoIbXbqqaxmlZpGuzghbi
AqETQW/j+QwOvS6en9utDofePPFklk84McrODJ0Pl9MuYE42IwI0ypU7SM3dlLub
qmL++ghNrCPB++3P7yi/ex24GpnuKncQlb7tV6pPWtKmMRDgZZ4WBLGz9k6Dl8BV
wkox4jZJBQdDmUe8oATfY8Bi/ayp5WLjXMBVCqDRYsHIPcXaSP1TfN0nHY62A6QM
mBGbjD6bG8SDkjn/QtX5+YTANPTfs2cDRB2AVFakyNveADzCD6tpUCZXnWWQlpzT
B5aZkqeQAHVGI1rJqUkErOJTuMtw8mNV3IP5ozc8IxtDforzGM0/P54hWaMYl8p9
/uu6qigsvdk8I0RKBF3AX1ko3cltls5Logjrah1FrrpFJ9BmirCkqm59W7GT+FiA
VBWYD9IVK1la/hXOnlY0atO9y7tTwzebK9Qm/VZFYgmLl+mciDuF9KxaG4SU0XDQ
WfzeHEb6nAeBg+hAC7e1C7cfQ/2H3AUc8+vA0OTkmMXgxKIloLrIcgLuYmB2KgB/
3cVlXNV4sSgWsE/ATklQA0uXSUQrBJ7VyD/lSlOA5os5TT0Z25tW0llARYldlPb3
O9cBrrwZ4TZ6673yE8licd6+X97YaOEGwLeQ+Q/0+YXxi5taOhBAkOK6qOmbokdz
K4ZbJOv5owxXnCfEP95MK0/ctcBOLC06ttIEIU4s7x4ZHSVtwfvwaHgAB5iIw9Tl
kY9XGjeRxo2vG0FxKf8yWvxGoHhnyI++oflJJrAU1n6Mjl/gqDIkd+ZNFige3NMx
2SRU1qjSJM2uKAnQf00ERKCiGXRTXsqz8XItvfZAseb16hzSXLjZmgXH1pwRp0SR
vKF6y6Q5k94CNpM7zKz9o8B+3NrFcE77yPhEv61lS9EswB8uJZo5LEIXtvK/xWpt
E3Fzxem4MkbEkEqJYAOtiy1hgHrGz5rTDZoCyLqj7hveOZ9BlIQSdFH6emOGz8wj
2nbs2lh6w2AkJpcrVsHmmVHt/Ajk5jU/uvyaQjxZIqjCNidOTZJ2UI1fLhl/Fk4y
A99YL8mkWxLw6C6eLsT/yHyKq6KercOKMKw3HtAC5/XBRGtNz74OQrdl1bGRvQOQ
iqQ1kZsUiBQpQCTEsxi8zPNa4fHOaS3SnZDVf86z2v0r5LcxgDafSNB7cXVCHUGy
BhFyEIw7SGEvLb84dI4gSGBf6XHPA/OJ90bJ9CWogLq678fFMDuxnzREJ9eWoJKe
GcLmvoCunEy0rXkSO3/xnKdmT7BPH8r+spQTXAfKiRo54Y+kCWPAlrFk5PHfKN2a
kT2WYqEawbuYCFTXmhnlRP3qG6j8P/5mLidT8A4YhBviKH83WboD8TqUUtrHD4jt
IQydzmFH7zPtXxCCvwzFX8GYxXWHGLein97/qhd3qgRFrQe2gWnI/ZOkjUJiuDQJ
BOsSnt2MlojTTMAAQDt794Vat3Lv+XwL6G1UveDtolV2R4qFLs+7I77jx7zfyPuG
aTWoIfwkeByfNn74TjYkcGzxexEsp/TOlKQs+PF9kgTnA5UdngskU4P6QsT85II/
Uxu6ZGSfYQHNbpNc2O/k54AjYSPMJ1m6RCE0ETrQ0nm0Q162PiUEwPMFMajhxih1
X3LfAmg99EZU9u6HbGhjK+epTfxZXmJMFVcwRgq+gJYMcPG9iIVgXIxcbc9bK+Dd
St5UALnNXIncrWPHVHt3R8NipV/ZJI8g3w/TOBRH20Zm+7vPhv9ua3ILL0z+My8o
puX2a9357kyGn0d2gBom963cJ0+hzcbPNZPCiC7aexFV4DX9DxBuOyC5MVHLirq9
Fy/XT+MstBa5ZQiXoqTMht263BO4bb+MlWdR9hYbO3yK2ZgNRZif2ycKTV71wE28
/1FJu0+o6+O3KJWF1sp3bpk5OIIMpELFFR+56p8+cgK+jcvX+kZ8/eSfc3TH2Q49
siiNYXuG092fo0rFzfzqGYzxwqjt6xIj5hj9RkfjolvC8o1l3q8UF787SoMRu6x2
zdkSIcUZuiCyAfaJLRdyTDA1evBCGoK6HAmUgHJJpeEr2prC5AVDBDUUuRumV4J+
SneKggJT4Phuc7l6yyDFkTegDHXEJCUiLxiasRzPnhPR5+Pka0o1sXojO2aeWALl
Am6qTjOOnePdoBnXbVi6+B88v05m7Um5m+QJRvHn6KfGpG2+y91lKkLAyc1oq1kw
ff++3GslYpWuvsOX0O5gLfyjz6LLxz6fUzHt0D91/Iw6oOQ/V/BB9sB814/zmqr1
Wf20bj7kcu5ElJMw6+Zlv5rwvl5AzA4JcHG60PLuR6zroffEO4aOHtnHoVJRN5AH
1Nz0vuOvgo4H7kt0spodC/Fpsz4OQe8Xisw7Qfx90TvA9BfSL2frriShgCE/NqTn
OzCzp6uelAgIcUOzwAdZ+4iGx/9eKcrI4IkUv4hHcFXciRLj1lMWbVSrDvEtEGkv
VDAL/n61YJ7cTDk4+gg8V4zQ+11xlxhtb+7cIy3pwS6mJyJ/ldo97MyhkmgBkU/c
oK50FPZSiyCgZrIXM0QO7bhYsLkAzNujWdwRMT0oN7/AOgITBr33U9s/oJfGnH8F
f6uNe+QIZGV3sMrbnZzSp9rQom57hWSGikngNrjqmEgJEgn+3GwF+Ri9dHiQ+x8F
iqz6MuzgZ+qFo5JhPL+z1x+hHhP/5bypl2JQL5AE9+VdHOJdomMhnCuHPG+WsMGI
sWW1pKFQP/Ajwgx8BQJxjdQkhAfmTLuFN6JwFj0Tkks2I3xUYLA3EGTy+1qL7V/y
oYo0MH1W8s/LZvqfsrz4npC/43rMCfFu1jnaFz1UpGRMDgOK+8Nue9zoSW1Ccn01
NlyKyJyRmbh7W+5QWQs4C8JMN4xB+RnWzHO+Hba71F/BqBpaW6mQMsf2THqxS5s7
SD0pE1/bxfuoTtGidewKvLyn6RJi9FJjd9BCmRWGMFH/dstqX5QxJwpDG2T+S5NC
0E4EJBmZKLSTVxNi3ylM9HlpliVy03BF2+25vXAndLp1kQ/hyna2CpiR25bT0+4+
LxulPw3nloAFik0fBUCZC43pufCRM22KZA/KZDbdI0uInhSvQBsXkcZ2RQBksggC
z7lB4PaVG0sXmureDia9hhdvB4bQol/N++ln1jVRnAk4lFnssTmkSDTzTNDbZeqq
KHH0c5++0eXfrtOMQW+nYkuBomj8I3w5O7TUEEz7PQkqshQaXIaK8dfcBf4Po828
bN9xbq+DFmwKLlHpgXFIxpAN1LNicUBZuPrWAurYqfKvtC073Cd/N77vDVz2Nvk/
hAphuJi8IFMVPcqOmqC/A4Fd84kTOo101AiHiP7hIQ7Ap4XKZEQoCFSb2WadkSAE
zi+daf+xMrvOhJy5SfTestgmcTnk/Y2bBHltZr7nNF5/Xs1Xhcjb3RWiDGHxF+67
ZPFdqZCiAVV1fUvURLK3ustrVeJnV2xhV/wxu5l3+g+m1LNph/GSmggIw/ft9PWn
AFsEBGPVCWm5BMcFhtxbnXJclYvVw0SV0NJ329DIo3b2AVDbF/DA//MF34+UdbhE
n6Vjh+g1x1lY0MPMr7E34VXb0mzs89oCRRaNL1kxje/e4Lo9v1hoRulcKawyvASW
ALPeB+k0ecjk+TlaKEzL7BPzFPwtDy9h+hI2+TZMRffcQ5WY2V5Owk+1HSSShjpn
w9W2llY5bEhs8ilBm1NRtbnGrRpnxjLAmF1DM48iG0M6F0nCq0UfsgJmiTlDudYB
LfYNhervWOshOzYG7VuxxjAkjnENMtakKwgGgKoqgCbgfFqLWOR/DcjbmUWEc18e
dnIBXDeZqw7LlCynZUkdTp6ZGQk+39udw4qDutVvMcCsPDfYys2vvpHBwL/GNY03
5eOHRnZJOA9UGbb4SvQWti0L3//jrk6MRMqINxxdzWybyQTt9b75VGTc88tjJMSW
1IBpg+VUVCotwQSnPtZY4yVDeQVx6f4fr07TFWGF9hXIHokmjCp6Chibtb+9yyc6
tmogyvgbmJejAZBqPbC1f/I6I11NlaVnqv9DP2hbfdtCCBN67iliv99KtRDTDQ/A
QfTaFVes0bfVhCMnO2veAitPX8yzDe/JLt5AJL80BGo5xlKMelIZV4mDgAuXNTJU
tzg3CxTB8+Eg89xU0d0XkWMLdKudz2aQqN5s6ceA79gobVmRVTnCg2E/4mfl1jBS
MOGPOdUJGfTx8ntqyluabqqBFVaHIvfXyaEzyNnuRqJWL3kelrWr+lVeZC2D8q/4
l1TrsWrcGYT5/wdVNoJ8I/IiNPrA2f6OAn0YPyvYUit/j8PS+4j6pQMBCzf3+dMA
ZDUelj8bt7fcBVY2DXgoAvfKp5fasS9Ngp5Caq5vTdSeS3oeyRxRti8q9KgAQnno
6yflSFKHIed25tiu/26PEiVGXqRsIMXW3qg+pQgaJZvHTkaqJKQE8+kPYtk4dviI
n5a6iWyqq+NLiZPKxcqGyv6a9srWYheWPaRnc7s6yGCW3FjatCjvj8oD6Cs4yb+B
iHa2sS3rn3+zlSm+iTmQ0P1PjWLhxQOpM3Zvimo10h+OL0snbgg7ZjRJmiErNr6n
G+7oN39psYWx63dIHEwy1lSfdRLZMhavx1Mk6fQD7G3q8mqrRHxNPbICZXO83OEl
hFTriRGEmrYFmX9w5+f9L2YYqit1cO6jbLDtaXIZvpYFK1SPeWkGOwKwFb/yXT2b
nwGXtcjhZxwz+EA7k/cr44ifiRaWvJNk3c+flmULazeSjhjvFwCOwGNwkB0ta4Hh
5ewDXi9VLAYay6+q1actVQeiGkbAmuathsc5R/Xxrw2p8uwamohUJEutvYqr5Evx
+AJHrDgs6eV0SBohMTGnQogXENSWEfrrsD6E347tSg0Qji0hNe3U0dekhDfMSDmz
5VIM4qdrsX1aiCfmMVuyYtbs5pdxlfN2vBbagBSmVB415qeT+wAsV9BV3AIzCLFA
Soo7j5vRp2h2e4hVsUR+O4mV4mDbgkWvivW92GofBPx8NAZ5y/SagKEvSqMeF0ST
ztk3bRpw/TApt6knHAfBi1zmMVV92Ht23chcelIA7QG+5pDSYj2NoyrkHsAZkFol
oOaOxdznWAclTIZjom5GuMDFuPu06r5LtGtpsLpILsCq3YzBY4vhebqAxHnrbgTL
1gEDtaahteyrwmKjqx1APhZadaW4b9wNEVyZLNYHppJBty4cjPIcDvtlS8dQwKGA
yxUQ5jiVuUkrtliUtyvthbsxCnw3oY7syMtWveS7oHfSfJf8AcC3SKJX0LFI0vh5
5ohm3Nx4lqq9vtFn3flsKXRrROu4+6lrZVc7ogRT4AoCpa3yg8Szsh1FEfgUqsDF
YYekYTBVjHynGD/BLyDf+4t/kRk6qPZb1R5cYwKJIsS2RqBMlMcwwzV+lCU7JNiH
HnBaeGdFnhDdq6sv8eljxgkYZUjhF+bhTrkHbEepruS2iBiRHDdfxk7zmuhkcWAH
asSbJdyyPLeO1yYMMysxUeAFB5UihRXYVatkvsODTCBFWr+B3nbfBgP5Ei5NFifJ
7n5Fvxg4KV0oF7VEjSh4XxawRtpXSHDscbW/srWoGy7bmQtuMuKCGt6+koQHK0eg
aGlgOpIvWdPFfNNZyQiXkznXidu1Vs3xmOuOFcDkELHU/rMR/sXU8hk/ot1fjPQh
aZ7AwehjCHqUUS8Yim5uHKKFCjO+j3dLneflIzIsZYa59UE0smmuxtuos97ALYjx
yijA/M7PrNuiXT6BcsJO3BXRh0BhJlUCqk9lKuPGL1t8H2z2Z8OMiyIIkWcWWwXb
axHiMIVcPiCRAnSopQtGK4yODQgh6jAx1DX+D/QZtGg5yY+kCw/nk46RxJOE1lfG
3/EXGAmEJDUf1vjqKRJEdGjKKAjBHZDmUDLzxR28iIXGQLWgkBKqWbNNhMwqplva
KiyKDO/oFYTiTlBe5cfD8KyDj57QibgaNPgPpcc2T5mqnLeRXoALLx/3agmRQ57e
Z4FiWliPP7es07kMSuwhackilOV2WeX0+ItFqdLOejgziFZEUXeiVSYe3Dt+A8p/
TxW8AWt7p7d1U9lX2oAThdEjDXFrxzwsyIUloduyH8+qYCWxF/YJQL7jHfThePvQ
7fvOhNSGmu7T1ljTcG3hfB0s1tmMw8WE2YxN0DG6G4zeg5dx7hWDTwEkYIouvuj2
+MmzQEbJTsqvhNXpZh9Ff9Iw3KWCgb88xsM2bmL/88L0WdlZO2LCGa+PH8CFGvF6
EWf5O/4Xt3CjJnI0zhYmlbeljkZ9TH86ePRTcc/9wQx72OjLLzmZkAw7e3BIyITW
qp8AarO6qJP4A7ldrHCRyoXVtvzwde00mPNcbcHwJL1tGsgoZiFoJ6WRlEJ2uP+x
RiqrS/+l1oN1+q11+0QoiTl8gX5cNj5g3vTQMO2lq0orQqVH4+s831Oh+jqfX1EI
lpqYaDJQ6Wl3tNDuWlkok/FcjqHFnL2OznKrdcX9U/W3/G7x9jeARzVol0Uvuk4h
uZ7g5T2YtCf+dP9ekrGx+POTZbc/3vhtON831kF+VuWM5Ki5E84WIzsWMzGZjCYb
n39qADXdE+6vjJ58Z6oBN8yLYe2atDoF7Hsuma8Z3W8x6cyu/rMNDrzOkKc7H1ba
isBlW/tWi3Euiqzja26XYoPnfBh0/1uhroxB64zrgmqJsbFxj13LM2u+efWTg3kJ
ECB5PGOaaQcZ1V9wGIR+rOyiqHyXspvIJKdxKy0Nj8tpLdbwq3+PvGJQH71tpf1M
3FWOdMlPYUwptNcQc4ByM8vzteIisW4bIJOliXKcCWiyg7YfGWGY9O2NDMV+c+n0
xy5vpsWNFXcmpldiSK4Rlv+XpjmdMjr5wVugvUV6UxnJax9Rsq2IxqelZGvQU1J3
3sMVYLki/EK0/2r8pCWY6PUb+pLIrqkMr3Bb8ZQa74YBO1wL7aWV1EE0BH6uQ31X
eLvhaxMX9nNPsRgNGSEHUvS2jfqVcF8/YIbwB5ZHQJhAX++LozP45P1QjRPfnKT7
Sv7h8cAW62CQffiPR1+P4/3shKUelEJvvRXsKhdH3K8YjgAmCuElwUD19nqyvXee
gMpqwUTw6N/fsCxJATXjJFYxGxGW5yi0vjyn1zN1GB17WETgJNKsylpXy903DIDh
UrRPwNJ/vFrc4BNyJ9EFR86iYkVZ0LX0oyS0dkKnM44AGVcavgqyxib3pzH58DM9
Z9BmNZhySuZZj8rJ05wuAksZYGZoydgPLHJuPsHHZ+NZPCO5gipYr84uAjEmURps
pc2z26O1rrWr8XH1dPE3Gj10VNzZ2KrhOTi6+z1VZ6hwcWwzdDLiXtmjuWvUQKTa
QXzkFTFFOe4Se9lKRkXEnvmwaEMifNhPA0ydejsUPZcaL5KZZfYfySM+bLbPaJFw
4fFjdoqn0TY9SK/xVRl53Iqwrjji00EU1vcChAjntKfrgfHRo4Ulfxr/dgNrHq9v
cWDBEmX6OS3y+7b5+pD8gDlJPx3lbLu9QednZ7KJvYHXqBR2YgUhlSeF33Qu2dIQ
NbqnqbuhCTSxZBlYbIb+0AOM37CpHtornEEp5wc4gXly9QnD064WN/rdOomC648A
NdY2ocuDPC6FzF8dYXMK0VG8s+LAH5dveE739R6A9L+pgALr/my2fGc2lmOwx2h6
DNMAhZ3GiaeGMscVmMeVZa4j9WvvX45v6nN3GRamVn6iRioYVe987+//qNQ0dH7H
X7/swAQXs9a/LLiaXephrlJy+D20SiB9JEPNKFAXh8FNe7rGbjB4hW7tbv7m993U
xc46YBtNUjUDRtxpWDiWAX9xW5d+Kwt8vHWIjDt8/qzI1ibpMuBPSmEVtHDfJRCs
/CxLs8Pu0xVJINhzyRn7dCIP8NYhjxM3RWKzRGPEKvPnGfbkKzoy6rwJbjoKg3Vt
tLI6L5QsL/bebX/p4oEtBIP1ef9pLl+qqpf/0RcbAm8bAY2cIipB9VQD98bFUyev
N1Lzm+cxLKcumWmFHP/S/N+ogiiuQg2Tn0BxPo9tZIvm/ROSKEgvDWJf5jRBF1uq
fICOq+CaKV8YjpnGuD6PUs14lHt3rXIKi2EGUOX7BU3bM81BDHNaHCx1VEdxoE99
MRX4qymcNgUzvif/JWpDBOErxnFyaGJokNmKDt4iwfhKSGBGx2u0Tmb9viPVvzNq
SFtS5Njd3n6WlZoW3m9M6dlLokpmDtVbIVqXqc6heZpQoCmU+OD/u3j4BCEXyv6C
zWwFaV+mt5Y194yRE3RdTUeC0I2xceUmvrm/Hd5BFv+yN44ZQfNyzdH+KYC+b/oK
NLNouoYjXj64zdjJ8uQ4j21HVDKo2dugU7KDBfcHvRMa7dyIptjg1FInoDMk/cJZ
3lvoGQUIn0XTsKTss/22VoR0UbqJq0McV2l5sZnyfqMiy2C0TDmb3esxZVwlbuB7
mgA5p3zomBysvrHznhlUDtdxnu+hn2lEo8GD97WzYZICflhW6O1QU0teHlwp3Fw7
VaSHQEWNSDD23E3mfPC2bqLCVW4yyLswZFUJ4sS0wowzwWhVvnw9TGi2cGl5RsMV
sZXLRFvEzDphlITEJK5JtyRfhI2tF5A8J6GprgnTE0QLpSJkIDqcjmncddCabwpy
LdR0gi1Hw+MSqQrtnSNPeFwRa3k3l2XjDWrP+mzeltYKEs32LxCbCZS3IZ4fH2IN
kbDBBpUHfC8OQKRsR/CY9afe8YvIr+uDw0T1XYNdDJaTLDLEu2FA3ewlBOtjkAfe
vqZhYQM6ViNqoNMmTgX64V14zGg7ZwvwuA52h3u0SKzl3RAmBmZaWPF1PTPyzedX
Z/fRgqIbcs4x8+jl4o9unn01ijactJT2udyh3tMTnSHfVWR19hRAEf1rhQ/NY9KP
IcfV0DBmztkEYWubMfi/KWKrXQmzVfAjT+GhWt+faAu9E5fi2wfbynv7nDiXFdMI
u8suSqYjdyi10kJCFxDE69lDFMuLjjrrLutO7Di//xlEDqa4yncyUldG/Pr7AnSA
xOUDd23QhphaT8u5jMbtRhNgymuCSHP10OfJ0t2wM5+H4wpJdZm+SXPfxpEXWf/g
bo/yLqyI9b1ng/DUEaC6mOqaR3F8iwQPr2dR5FKZRvhHEPWj9G4Zyg304LQTIG/a
BHSUWI9x/mPoSS5STzOBK3xgFGdt+EENOS/6P8XClEa7Tpq+0h92tbJT6vw0atIM
gH6u5Q1q0cknxORicXZyS2Cge/OjPK1cwGeaGcSP5id7HWqjbRhHlPUwQoPcB6NL
2rRfbv/v7mO2PG4fWdRomDpalpiqy+prG+igsZUi3mt98InVrbTQlYsN1NApAsiE
WPiZQFiqMXiRgQ7mTFqLw5A7hxegyaG97btw3vFidFyGlDjycyp7QHU1TLx44yg4
FERzBivucLu4aU/WQTp/BKxTEbuKRCtMidNjOGisfXSFZOiCzT++re1K81wdiS2Y
rqE0a1OSjR0Mjt7BLaKT6KvXa2B8wHaHQ0n77LTikyhuJ/AZPQXeYkiSCbHHYEaj
pdH5Pm37wlUmd5vrU1yWHz16NyzEYmudWEGbUulwU5otPu/BKR7UD0+cVMEbf5ud
N0HsCr33pPan21ybeXt6wziSJW19U1zTEtBsbLhSQfrweFg6E8DLwHFPtR+qdCSd
fJi3ZY2NjmNd8Cj5AgBDC12wlN/lO2d/QknxycFPG85Qpj0P2eSrfEz4CPFbAaCD
BlNJtvAgTw4W/OP6JthclagJGpcE2m3KZw96xDh9FJP7kWC8OK74ryZJutd6DHaP
YUCNb1uAXXU+Sd4hiX6kjkGIED4xaRf5A0wJMU789BBKYVrTwMq0f6w+C0vxyjv/
wuOuJ+e3CeuxIGiIkcXtKQepyrHCcIx/PJ3CF0cjs1WQCEdw5QpDLAaL7u+Sh1Dz
Rv3a5nJtT1t1RBLHJV0ACc6Uzt9mIzG9qYg6XLwZTnciVT4Vk567sNGXoEO1tX1k
HUwl2bq5H3qt4pHEKuqqwzKzLy5Ecxea3OMl5dWxq2pmfUdIdF/o6ChyfITGi92E
3s3fOeOiPUaUZv5qwkvlmCRnuEPUxAPRAYAaWrRBFTN40UQkYS7EwH6xPLr6lDvz
R/nrexore6Ju8Le5xlPR/+gUg+K+T+SPO+ul3VSrZQAfHHWPBKzHEGFpgF3h94nE
eO59jmQBNfDBVDPUAmQJG4PPhnalXLnPQdQJtTmNN+bYyHm8LdVAGQ6iQ6Sdj6R3
6yiieVzdMxchwsgQ32e/olhKfeJvE+idwar6dNP0GkrEhV3MEpJKTUwmFfXMfOUd
GJo3JOQ8Ywti7w+rt9Jdlv/iyt9XP4WH620pOLXhdPhAaEuG68p+EnlC/FaEBRyu
KPAOYyShAwqa/1J5tWLEe0Hw9byo1zZIlEMvhsrvs8UU+Zw8qwAHzfND/TOGdCRn
4pP6VD+tf3nq7GdiwbxJcGakMcEe1Rqpxa+EEPpo3YeJ0SJJk87QDIwkT9IpxrJc
eQiht/NULJ0A1xbbzFLldMZ+jh0f4Ux2D6TGVcXcWAfKn3i6fUdR8/N/K3+k4or/
h5XY2O9bvocjwkR9AhmeQSwJScPQZMP3yFLC1gUED8H6GkJMMj0DcrBfdCfFqNM0
HJ25SI31hPAj0gqrHIyPopxLDjd6UOqPEkBFVAmW0aHfCxc9f6cLu64LKYQyee2M
naYiD02wVNg8x3Cv/HrzhU6G8e/IySE2EiMTsx+LZ3lCnblkegVBs5A1K0OMYrZ/
WiuRyXlFb+l1rSIA5yp35yAoJMbD0BjpjRRKISfVf80MkFbICo+gcHaOItNk7qMf
YY64kp3CyBE4G2TDqA904x0zB8rf5w2uJ3WuDvAMXCS8+4Rnt5IIOAQ/b2frN5te
GtNHY6CvzxWYpP8cc5Y06gO9ehhNQIAWLPlA1W+mEkbCZGg6TY+o4TYvmE2yhVXT
ZlnMk0+gBBEcIHzzDKIICReLwP+/Cc/3NaHFUE4Z/z1Z73Aevs5AJzcuYFygoxVZ
KpEbWipxu80VWrBAH2Cp3wQoT+jn0ZBT+Dz4DDXimkGMplILcvsS9fjPQVblwzhP
jUvTna+F8NVMlLomN7H36fvgIiC2avmuR9mgKO9AjA/wZIKS0O5Zwnv5oe3Q83Vm
DywewKZMuOyweEuGY18y1tXwchpOGz2xkJldqXe8vaxA8IPEBRaZ1IGxRrW/gLv2
7C/8T8WsQQ5PmQpaAmvmjWc+AenpMbhWShsbePKwinreOrjdoP5EYJFGrx7kS6/A
PRj60vxjkk9jObdB+pg67nEr3KnIpnuGBa16+dkjyOB1Lbuty9AQdsE2WmNGHgGM
5cswmdBS2Gom9UY1Pjev0iEC+PtujxoJsfXDE1CZeaYi/+glxdov9kChoSJoCWjm
QbLD+fkNH9pIckpKwwyDchNoo3azu8Vf/jeWK8y+VhXxUJ8DUuLo1vA/9XnkvTJC
4HAxL49DPKd/ajBYZB/oYNHLex1aRYDXdhWZkeG5qgTmBkq/847WsgRmM3YEsTFA
O08+5SnSfhSjS5bNh2zObZ/i2+gfIC5N+HkvK/fi8iOtlOxhqdCevCc3r+j2KlBW
gbJ4B2T+zVyYW8ZFvqv4NIkDCjk24ngKy2SzgUE/D2bEoewCuGHnf38bJZw+K0CK
2lBmWjaUwL4Lk5/GOB8sQD3FdrqN4GTr2ZlgdPIw7JcXlRQOoAbyVtyIToQLxIb4
9CNcR5kNqgdWheHOmLWVLg9J7jOaXtSl5yUFKEhIvBD7rNvs4i16oIZlLZ8XIF03
sC8hZwmE84SeIqvLpEO+td5acQCXiF4lseupyZ6LJoUElrQHoE3y8kjlMnBLdtTV
Y748IrBXc2xTLEv2DWXUz1At9oj24dzuadGO34yL6DOSXDHOoG0giHhGsYmLXqQB
sKTUDuPbguBKOpTWXzI1jPbnz1Tu6KRvBccf/mGUaFK7V2x+cbOrJVpfFbfYK20o
VzPU8QYMgc/mjcLFrOCgKE+FN3r8ZzmzZiJdkmyqO7QN4f69pWnJ1LZTUl86mKkX
gf9QpinziZYv1xzjoOU/XbmnlUdPga5cOR2g8WMMossS53au/kTJpTpnGL0lUmTH
gF4m1feygWxC5k/VRT34kwm0x218g58A0DsaGyPDEBu+IfMkJPO4xLxSQzbXXPJl
560/zR3cUnwV0RgwFjX0CIwjDBNXWDi8yW4bgWlgoB2C+SsE6uWQfM6I4cA+FhGJ
Kk9JYzDTom/0X8q/xcz41CEr+PK4oo219O/JqadbNtWvIIYRfK23ByY2B4fTFGj7
iS0wIXy+o+L4TP6HL6qY+VJNvm1FF1Kq8hEAfTs+IfYn358hkvBmjwHSM7a1IWYZ
9o5DOdzaZnJsae2EcYqFQYA9Tg7hclZTdEBtsAjhUSgE9yGRFVC7o3FPLR9Jr2Sl
1uWPQ8GPrc/bUDKeoRX2zKz1Gaahf3QoDJGFFvqqnuHzBgRn97oCCBQ6gC+e4wiX
IJXk9Etk1A1Sq9yjSSZ9VoRlUl1+2BBYjgi8gYyEtSYcuAOS5J/ypuO7pgKYawam
QLWmg3BwLW7rdvqXk0ZE1hqQa1AL4TDYo0U6lZw8nVUmkxvwlcvnK8iVeUgp65Ri
4ywRxCP76S0SIov812BEj8rt38yRJ0r6y2sCbg2/dsR/Of6EMDWuq30Kbc0lu1PX
2S+Az8Hrg7xikCvIl19sdvKc9RV76EbMtWoOMt+gc6RN9CYIbGo43vJDISMIQvti
HAQ2jUsRP89KNWmyC4oTfEvqf9TAGo6xbCmmGvqsdv096jn69ENWea+1mZRtm5NI
a5D3lS0B8XAk3SLrleNoIXXMTBE2bWdt/0sisvuiFjwy6ImgDEI+HmNcg3Q4SUpW
mMcu1LebK3DlQRoKYyZuGGFGuyt4ZolG+gKBtJNBoEUYeuJcpbF7k/QqvU5SDCzc
uQ0iic11qstn9wqyh+EJTSv6J6W/MLDZ7jsp63EDEvMAyH/Nslo395DXRT0lhBp3
J8r0kYqrc3/L+l+0fiE0CyiRLr2C8E1mPUzFyobH1YHZns1sUzlI1NSuEog2NzRO
4gU1a4XnBe9zXBPVnliCm888RtVnFS8IQ6HWAQCgQY0BzY6SuHrmiQRqzOkOnYq+
A0dJOnIxv9Rfbd8G1gDw+l1dbgv8CAfJVt38CcwKUijAaSZzZ07oR1ni4L46PpHV
0ykPb6uKEqNon4I1KFrJjV9obJ3g1vQuBBU+jo89MTgLt1Vuzcw74+9cD4xM7VLb
4MWkHhomsWVYzVr/oAkPao4azTRCpq7I83i05vzDMZwfKXAo0Q5rm/yBSMbQey2n
l1yx4xgfQz7fQAYXISnUKpOyXV468gp6J4ZOBl/ACIPX7R7LVTrhhgiOTEzGMPhX
K56U77EQFOuF2YNIcC2xaM0K6ZFfbPIcEQZIstRzEvqM8hQy+82gxNuw2Ehr9g+G
sJ7QPuG785Cul6rDqfRTMnqK3kSDcGVZauxQVOchtYIi53KgB6kM4bMlGKmRS39E
bsF5grL7W+zLw+K7qdJ/YHmG6Bop50BI3FRyDWG0wMmmxX/VtqE15sBCu+6cj6nr
P1HymU8+iBQdpUAv5B+S3SzmAjNTnczYolMMhmwqK1nF3dOebRjOpqmMDGls+ero
+8JPuIXKKgJmtgI2lTSOhJwyqrfXay0pO9IRgfWH5Zh7uhspKeoZ0ZMaI/PdFJJk
QkvWOyAyj1+/mzXiLunsstc+ZPs+tgyPxjYpNj80AP8X89ptSNaCmD/mx089Ph0b
0rvrEvV+Nb7IT9mircUjdEhzM8vHKXOOTl7k3WTHyX6ImF16kdjim4Osa6ql/8zF
3eOA30ay7YtqjSKoF/u8UYLCf8grM4oYcRlWXaCJcj87cXVSwjcgYp7ALhIsk6eU
i4ql10+KWtX7I8rNMjHxKBKtbsjntEepDPtsmGf10oGPEIhwBNJZxk6yD/TuJz0G
Gh20n5/j9rYui3FnjQ56WNjsl4Eo48YWPQMlJ7w3ovuEbuMe3N2xLc0E8BbqQloc
W7/zKuFeVgvFT2NQUcF9t78fuidaiB6nG9Ggn8fd1gOUniAbf+jjvAEa16Slk1x5
d1CBD8CO0f7z318BHtrWa0Lm1lEnnlgASUklnSdGhTvvZScSxA5oljKjAfhydeq2
7sCEceKmG8f7/MGoCajRnznxJjoxCtN0XQyrWVYBxswWNkFh4VTZU2qw5QiYxPuK
aN0/g5DKj6OzC5m6/n2lFwX/9XFFk5Fk+4+PpoybKntFxEWuHbZpLGAUV0IgfLlZ
x+aiPwIRmFMNtFepciiFRWol1OWNJi4+t5IClh3k1UrhK1zLx1uSqabWJmOluDl3
Eqi/LQJCC97ilNV8vA1x+CkHUaMgCgg85WaIKyQ2ycnu00Ph3sCJ8D7Aws3nXqPC
VD/SvshPC0r1hunyJYbah2jQdw8nsCxbmZ16H6iTSAJVgx4Me+N58/2zSQ1Gwoza
RAA5F3/ErPHqBoaUTE10DjRhbreMe85F8CQm8dZSHpOJVJsa+CMX0QjE1C3XreWt
oKPvX1vkB0ULlF67IRn2QZRr0dAuQZwELQLHbtDLFEZT1s4iWXXFYZMwLlHfqOo4
mOAgnQYj0ramVVSEVUvBoAyDxnpqJYoBKDFo0CN4gpgCcfi5ZVXHQJb/3NMF7kZp
30VzZo9g5ZJZI8HqUVHfd5KNuy5QXrT1CHB8xCx51X+gPT2bVQAYng8km8dF1zdw
DokDULqEPNuwjYxxhmQa731eX9N0Iu7VdswksxKMP9f2qUksd90DD8yzbL+isE8K
Sisma0gxbbCMx1ZKHFn79dPfVudTm54yaind86qcXqsPw9t8dTZZEzKJ/HasZ1Nb
tSYhstyItdvx3k6/EvyPYoZMwEgKoiIfzEMkhZOKGmcm1e1qRP5ps1yPflp4ocy0
ZnKslEl1VHk5MTO6WoUQk0mFjbbYMWai6r/2OPnW11OLdn4MU8gJJtyXA+L7srUd
uQGJVG/CjQq3tzrdzZ8XWsFXjzhbYOxnCQObj8fA2GeM+raI01Qr80gNMqzsLEoW
3yW2DgPTtm8A3EhTAJ0u7G7gWafXxiifSTKxHaqUBDEx1arjeeW8XmBpREXylJSF
oAGR6x2EeCNj0JYJI0HZqgCphhSgC4gIVDdkAqTMYeZQyevbhICZYolnKXuVAWTb
W7fLABGAFU55FpqHS4U1mDPPG6p2RNP/JNMaESms7Krv77B1sYvMiZasev0oppY9
DMk+uc/kU1KJaOk1IiShpgiaV6TKdTRh567Nymg+kQ56qwVr7d4idehJ0OnQaryX
z3l3dcvKCf8uSWJmrWILrwrRgUqV/pRpj8QboPpg/m9ZEy53iNakznePrbmR66GY
cZlJUXecdeVZLE6uhk6Te+h+xOzdtYQj+qkd+9m28li/m21x7bXhciJKix9m6nij
dYkwJrugLISHmRuUKyBJWSkowM5xPhWoMe6u7HIsjcj84rvGaqJyylaFc1HYm5bz
7wEa+u2bL+p5lNX1nutbUcFrGfjT0PWH373dBbTdZw3aX0mJZ/m/rXU0h2Ek//dd
NE6KY5ZdHKIHpWtupYEwdhPzBW/hzC1vMNhwo6JqyKLFFD1V+cSTdUnz6Bhgq/UU
Z0MdVDUNGqRMlUhvn+wvyEGWNr1bvVkojNi7simtHuD2nSo+yPIpyYzSfSqEOCHB
P0h9Nu6N9SW6A7ZY5FuzPZY9KUChNiQQQrDpSSRdColA4aC7+7GbO/DKvSf6VvKA
iYdNdfTPPdcc9b0SYwpyd7Ti/hNaAqGPhWTIqkByqvA3urSG+/JqOXAgQW5ChzGM
MRt8LfJyLMuP1FN4Q7gIscnn/4kyfFpL1cRuHahLXlnSTtbYFpWUWRwZQjDQNTkl
of+RhBzkbrB+7+5iBxbWDO2Ako8W84gZRQue1MhPkrMebaNNLS1QKFaEjE2hE3Cu
ls3p7jborGvf+YegSlEKoXFb4pd3poxUut28WVS44ZOb5UGSwOuKpOqTlobTZh0C
vERtXj8r9dNxmkdkE3JHXWMP/pdpQFv32SvR1frWql5lXt1AQNFhW3kQov9PIRtO
wxQIX2GHOPlC8wofcL04/F7VM7uB9BVjEdN4VvrawKkKX3n7Jxmd9vf09ia4Ngw2
YOznEcaJSEbVbSXxVttloAu2/xbO5/svC9tUcLP3sGUXgodWYj7mrP/hrYnDcxL9
eCJPhaYICZrf/afcDVSP7eEh1VBSL6z5ejWEX0B/NWryCEk8TKYZsr96uHv/v1Xh
lb9F5T0xsA+SyzuRaZW9mMRLqyd4I+icMkCpkAprU4wWmPix3uwN0ZqkKfNXsMhW
hQ/6V6AB6goHCrMoHkbf4KMLf5221JmQ7YQVaBK/6KBFnFniV0PiBYFwN7KbTzGs
qkQCUB/H+93Uga6hs3yCoQBvFB2voMWZ8ZU9n8tJ/rbM7EJa3BcC98SUyhD2RbWY
9GDEEjI9LfL8FdQf+Ss+12BTwiURRprQWb6Zj3Pxu+sosFtCMIcAg9JLq+rDkPpa
I+Zot+r0B2DR56PO/5/EIr1OvYX49EFcltVqS0rdmC2Bwyh1zUBcdyH1AZnQaRx4
T9Eg47GMOT5kmsQGU+tt7FcHCEYb5HKEqLy6dGylAA2QXA43JfGKK0Vw++R9Q5yR
JM2YcMoLxDkyu6U7uFq3wHQlHVo3zTqsJcyBnM6eOnd/qoHjdHn9sImqtX+Xbkjk
qSsUbacBngGTrKhNj3kDKze+e9z6cIWHB1Kq1uPQQ/gQasfNEe1M/EAWL//I5QQF
CO4bCk4jLwbXDB8HEeB75viTol/rPS7epI4+bLXtPDERKMm/QXRQKGDdPLGNuEGW
JSdtZPo0/vDgXiU64Lz+9uQaEJhN1wucOFcTghu+lmST4EjAXDlG3+7O4OVGW0f1
ky4920NaHeoP4Yt5s4UfZlnVD1dRm9rMKW9KMQ08qqiMJDx8iJXwe5pCesnjnJeR
7V4MYNmAZDrH09ZCN7mcO81/rop46ktLmvc0KS+i+gW0vPEKZAC5gJl3PtQIcU/X
euBx8/gPQ5KEzNYyPOnmJvKtf98YbCouUsx7nanqEKK3027YifIWDqJO9wgS5BGa
l0Qp9L2/TApPuGkO2seK557GB1C8IktvWLpFFrtBVkgAbxlVjQ870DjGcynEWhq6
rAQJBUZ+ss6DE/gslrQxWgfO3t+QloHBZ8Q89v6qWwpVLLI/CqUbOYRnM6SwBX5p
VNiuiiqFuhEtAZs2mJyZUcFmoYyNPYCOPXJIEfNVEw6g1KJUnF0dktmt+EZttzzd
St7ZzUGwHeQqZBYVyQaHow6TrgPpk5p3tBHTJVP5Kq5v2m8fOpp6z/nLzkjmB7Kn
vYC5lnrlWi1kJI8Nby61IH98haLFGREBnAxqvphJwvOpa6PGJ/OwHYq2//2dob0j
Z2XqlfS1c3vvHAOe2Z7jKqZ4g4EhQ1VXg+MfFoS7Yk93so8FjPuJEn9Njj3DjAZn
YBW6NbinObaWPI6qn+qMZvxY2agdGjJTKIU/i9Ij74/8hqDadkGh8r+KA8hiGVbs
ElbycqbK0bEjqulfXcC6/RxRa5rxIZxKQFU4yjDTRP8lu/iiCnDonqDTDg0CggAy
G/cDaK8hvjsHTO+pFG/OeDmGvNryAyUDGBf8lw4NAWNMfr/pCl/CpjuH6cvSZy0x
+xqVJ5foumLht1vDLau6j8f0gRFp35pReLZwove1w34+5I2EJihg6Ahf1W+8ihPq
54DUfJIqFyfYfhx94hGB6eHVAdenmaOEoQhMOZ6kBk7uWHlCqFnRBb3r2W7Ee/FR
OfJ52Egck1PaR3zwkOoDRlRoi9YrHvlx5SfqWkyCnTmPHuMwwWd5xMeoBGJFg1vg
zES2+hZzfdjEPbB3Ib/Luh0c/fnJ07sjnMDYPP5UeAXDpd655VD33Im3huZ6nWDK
iwg+2lRSjgsoz3kA9qqtnpKe2aNDuBzUj/dq74ir1Dj5caOCtJPQlCz79R3n6VhE
j3O6IAk/BymhFVowLdkDzHBcDXmGigKXAb8UJl0NzIZurm5kvaNnCtn8JwwKQKQv
3ACio3rhB/P/rKflsdCNlaVYtFbeV17KNPH/hbtQZZVW2WXkhsE+xhmL9osm7RSS
Xs/ltU+SStBRyPjcximQgP1nn1zElBzRxK0kfuPVxHuBs2R9x25mjBZRMenroz2J
6veHx6GLA1mir8FgEnqRwhH0wrdhDXLeTVcnx7XYbAuxHfnj6Vjc9WNjqvdNs2Cz
D40mh9Ggb4WKiW6aRR2T5Pe2DtX3HrFUcTlMJAlxTfBzAKV2GXfoJlb5Yu6QnJW8
LIdMmXW+fcV45gl0aAerAhBaH3bdoOBK9yNLVeIvQjxnDWDIxdvB1XhbOf+Wvlij
JbmPUUZVQWV41DCMDG0Kbiaav4PrVq8jejKNrBAndLVR7AEgi3I8TjIGkpl7Jtia
cbf2U6khso4/GsPjAld4R7rab7maIvUDrDRJ5KC0DDP71Isb8iqm5kN7mh/+DJJJ
Iy5Ymu+cfBtmBOsMuc2EqxQg7lXL5laOunD9P8osF1Nn4cugRMmeDYXXtHkOgKPV
GEJSoBOqzTNUg3W8FAUZKan4weMmQ6iUf4bCOkEE79dZCdNN6eI93o5D8sl6dJkI
b2+QReTYcA/Qdch4nhCO3RAz7GQEGeaeVhu8MlGNNqN+fC68CmV8KzDweZjCrl/P
EdYsrwCAZtP7VU+C21CnsbslBrFxhc0/0jIyJYzn/2Y7qt+sxe6p0GKgpGnfB8lQ
YiFOqokE+kZkRw5t/C/FXnkP/JlZHAlI7hvlGAgYWdUVLe30KtHI3KqchoiC8Dcf
U3H0wEQ+AgSrcvIHKRlXSYTGIm5bjeVKeWt7IEOTRKuYbcdcn/2lE2gV4ohjVp6m
EvCd/aN4PxGf6lsiuDvxMHjBqPDzS2FvILXigjfzx8N5XnbbzJrqmTaxqwcsPNOW
LuWh9aEEw+n+skhvkwCQBHdkEdrmovJa+uJaXdXpMozDYfciC/d/4cH20E+/5VCc
sWi85Jhys70bnyM7HuyHbPvKcOgIx1+xLTL570Gu134ooOZe9J/kN+SJiEiwmyfG
OY4Ghmj2OhuVb6l9BVC9xUsPLxJGbtf6uSEd1FAjHWqrLRYYipyUnWZ7EVmNWxrr
/CFtH56WxwzlU+IsBmNF/kuTFoZ8EdPOoHU5DPGU8fR8xR4oWkWFAejYqlyVKbuk
dWbH6Xk9jfLF2ZQTTQaZ5TqAmsBXR0kHPv1R3zOYAdleaxbciQ/8rLOvAGTatdh5
UZw8obRww9urcWym/C6/yKb0Tbq1qHxCjWnHsJ1UEsqiUFR2x3GkBBlI+JmvTn9X
1UjzjnvY2x1TO8aIHHqIbL9HFKV87N74dwWWR4QNL2d4K4gr7/+tN1azlWb3vkUQ
MEOQNngEzF3SAhw63IhzLpslWIN5NbOD5YceKigb1AInnrKjhY2GY4Kmyxud3C0v
CU94tIE1QE8GFNO+lD4bbkRLeLDO6CK3j3uPD4OiIZUtHcDSfxYd3B9jWE0waJ3r
551N6pDir4qwzRJvW3wQLRsQ45J65/GJpOlnqB/offoOSmMzAWK/xDa47TOyOOGI
zoZ8dz6g4SqBIAyuNQJJnSIi54EGZTfBq0URDCf0O8PM5hc4GPZSebKDkBVHkKmM
WsDL91Oz8It/aFK/iYkMWP8zqhHVbk/yWeqEW6uX2/V/5Dm+9aOMeNrgULrpiZMp
3kzSUnr6aTj02fRWn7RvO/V7E+KZ8CVljRUka78aPn4jfpP6rrWW1hc9QBbgxMkq
mEG7ldaz1kO0ae3J0UoptVXQrlDSCOo4xL9TDzrFZSOaybvs1aNeAdsWX2ad6UxA
aru4f4aSiv19PFfeYFO8xOhr3HQGnUXEkk4no9X06T79E3hkRxXUaLCCQF+N9T7T
ODB+OZcJx588RBinEZ7gMve9btNnthEZFaMD6iFPfBLQ/7KgXua1cTKYPuEAGVz6
ya+1sgM53CBFf68sXeakytbvFsKHONzrEDcgOMkltMzcJe7fkwwbJZ+5J5AqXK2A
h20KndEQc2fYNsPT+4toslBEYIDsLmTyGmrZv41O52CoD4/PUVhq/YPvAgXBddBX
p/BGS8iPzQPa8UYJo+iSHK5wR/FvmniJi/xTnOtdjInyR3G+CRkGRMZJvVnKKbm/
9KZQ71hgsOiBk1z/ud9KWi4ryObPGrzQhX0ZObT3x5lGnZ4rtBWHj4ImOx4w/phh
8ymZwT8myj+NllEhVnff7XWFhPrt4CVzy2YF7TMLyDSIwxgo2Mh/9I7DeL28UQPe
dWBkPn9xydggvPtF+Gh1fY1c34eIRCdUrVoDNaSmqQIBOGl8Aol5sV+oZCzpZj8q
m2o2mTCVoZLZjM+AkRVwtVlT9EzOTv60o+eCSV/n8cNJfg+VFoK55taPOuVgtVXQ
8LsYM7Tu7oMngwGWfTma3pcL8Gp2GOYiW/idjRsl9I2UUNDN72vLsFl7HROu7UXm
Kdv74gSoB/F4rURqJXmdTUtKiddDEPnSgcPcUm9/ffj6b1NXvifji75sBRR30ntN
15jN0ERrk3a6moyocOM5oPs1M9/9dGJMCCStOTFd7p2GIdhx1kunBO42pvTsFepW
EPoOh76yFqRjaIxgjMuXv9gZDRKoBoNpgB4C0wbILCIm6XcJkfvJ5HmW60/nGH0B
okDMbLZHrisoEDjDiAUr9rEfVtUOT7j7zjGTJLIJmjRp7+Hlw/KNhu9ZsdPKOXmQ
LXBYHJ2zvEMqtLnvJ2dbD+kffE+Y6gKGgZjukLNDwqwwieELgTaedjvYycfaqKTN
2VgYi9KBJhCLPqGRDUyyjFy8tjq4L7Ii0wK/eXbF2XX30BRC7zloGxYasO0o+E+3
kghPRR3pniyWFk/Hy9gczjWw8z0WuItddU4dEivSQlOAiR7czIKI0z1nzXCmgE5B
SM485sqcl28MOXVJRAkMRJDzs0LaG6E/SEJxRCQDFU2gB+T3l+y/z3Aes2ZMrTfU
ueNVJAFk2yUNRihN8Px6nZ0p9mVpLognPf4KM6lxYZH/dX6VZQhBCEgKWLVf1Jz9
DqLHcUQoe6t7aJKPmggBzeQ84w6jMRD/C2eiOFI7oOqgrhgZdBJSBywhO9oRYeAK
NoqWhITaPZA7eqhgASLOWR8lO7Pn6lDU/Rbx4Y1++UqYI+TmTOvNJ3r+ORJEq8LM
FyZG0VUcYmkN4sWXTYu3w4FH9Msylg3tXQYQFenOAfeqpGi+h8pyXOfcSvjh+q19
BYD8dkCxMmecQPhYEXl0f8e+UY8I3Gbo07GEr9V27aJPOovjPVSphRxwC7ZiFTCV
gtiXGNK+QOMhS8ZsCcbQGbSo3hGJht0GSeybPwuduXHyZ2F53DSeHmOUoNOCFZX6
F/xXWKvrnaJmGT4B93qJG0pyIwTsx4WQJmnMAbw/oS8p3Xt71rqzi9W1UxjYboLI
Z0vVm5J1BS9AXglZqmrcajsxJa1qhMsLGpj2fL/SKzu3LOdZ8tssw5L8LNLpjCv5
X3ovD+kBlA5qykYpFCxFuQe5/ZqxRf/91JnlXNlRbY1DDuVMb8LoM7fhXmCVGYp1
hswtoEDXHd10HNHZQeP97lmKYWS2tF1GGRs2HPqtXnGtJAof6MhCn0JHLwOHQ+SR
dYQ7fUcKWJr51L703EWz59nETfhrhTb+wZSF+85QmPZd2vbm6CB7NMOjihPGSINe
SA9jqzhhHl8OcWjZBZcBA8D5JMFIIaRYZn76DiU9+SjAT6ApdpzQg0CMucWSSaK3
kdGOrCO2nq72jYO83pp/igRhvzRr/tahsdKBo0WqtIuMHZLlDktFAfPnYn9VP5hf
a9mBek9ooTl6b4/LFZQXY6kNXuTuj8vrWYKMIizLvhnhPnfo5gaHBxIplIk3fJmo
Ghy4cvtmk2Wf4LArT42pcoB4WxnNpgxWZz7YsLZGKnWl2xeMs5kC9U1j94ZMglQf
5sKAkaD/O0ymqRTTHT5hmWdpRTWop18M7Clo+hTlrQEph7byFS0TftCjhkm1YM4L
Sow/Y0mbT7ngBKlNubgFuRkQiJLVlQ89tc+AXZOCfgwrNpDV/vJk5NFY9969N47o
WCY5SCj8FEv1RpqDsH7y57l1BAdDSeumJ6Xr1fu+hvG4M3jF4FQ6+u/wrwGC0M6i
j06C3Lqx1YEvDQbamC1FAcwoE+bZeBKLOGEC/WVk088JAc45m9xr9wQDCDdn2iF7
KUT7pbgZ0+/9HCTVLEdD6CuT4GMQumLfNQtuzzoc5mkBltEpyODhhLS1RXQu8DBl
VbXBikSe0kA4BFC4VYO5leq1sycJyupXnPYPqNsnO5zPefRz6OyuC/0HQU8ZFACd
VK9bDhn4sF4aeojIrykJqumBztR7dFjqvwESslXt4Lmx1l3dDkk9jtvtTS0UFEXS
2Si+OLZ3kBkyqZbT/v0/WX9ZQ20esEhbKKTQeIbFEx1az7joimT/NgnoS7xykgHH
XxmQVegemnygwLWNqN3xidO+8sGgInDfv/4ahORj86gFKyLNvfzKhCLMBb1B0Ism
Nu/63RiRthGYBnen3vdklBxLbAxsybop6DLGUwIHbKI5hDcVOZqTNmQDx3S6hzKe
AL1HxZDxQ/4XLc846QO/k1j+o9P0UrRfivrHAAeapvhJuUw9O4KkM1lAVq82SZ08
OkbQat/VNvE7Bkm48e9bWkg43n9o/1NIGoJhu4ljoEcFt8WEHY/NZUu9Vw0EHBjC
lSV0aL8X6yO1gePg/i47lR+wOzJNRG28EGldKxyGhvjyFTSODhLBV9pbQfk1sEIi
RjFdCVJnSZnLOpG6+5dkvIQv7yv/w1S1IU6BXH1Z4lMkZrqLJFYp/l6JsH2RErhB
NT4em562Bad/22qDyPILQFtUqnMz/2SZpU7nnSobB3WeGpfvO/fTxXbaeAm9N+WS
r2/Cg1Hbosfr/b79yQCjejk+KUj0k4TKaBr2j3rdG4DaApujc1dfCw7ujI73koot
lHQJcpytkNvfACptYmdVZcQ+SktCxDye+87H6KNl5EcvM0523TOP4xcyX6m1wfpF
gSDwRB58enNOc8bl6egNy0WjyNYko5jn2S8Jz9n4ZCfEBpj9hGavKux0vGCz25Lc
5B9gryqpjJnctJFzJEovMrv6mXdr7ZFv56qCvi2N10KlqmI+FvWXHUFkOVizNPEP
VpoItruJfXW3P5ttypaupt57cascLFs4oqsmBuiqTGFfGxKwgCwQoH2BYYivl1qN
KkRi8U6wCpCaK2ZQp9usH87jQAbYCGtgFMbgu174jfBxTD6XOcP1ntorFSXrRnsh
+tdiu3sLRDrijMQVJeVTm82lt/RiYWwY0MrxmRutL/cUNO2NCkKTOHafmxGWLJik
i1UDFdxH3QdhTHXf2ceb1QdqfKjscWEWvZV+AJ1UBO3Ltg5Xvu6eap/loalHl0Zh
bfYxUylX56osDwitfUooPEpiymyy4ThvVIaTIVc7S4JZ6tbQprjVtqVlIfijB5IB
O3OAEjuvdddvnwVLNAzkrPt2t5D1yixncrI8ravLn6NFUk3j2DeHnJdm+9umADn6
SLDmIqiINlLvYXy3KE+BClQN6gcC0DQmaGoQzYp0uKTPnF6BfIEJPPYmuib524jJ
omlmSzK+gl36SS6Y0F18UAokoUIhhGzyQCjihp1jyRi3H7xwiyN8Q2m5eeYhiyPI
Yj0Un55ZXE2JywPXZQ07BwiBDilcKvnZcdsZJgqiGb+p0yRmLOZ2nt/gNVyUHqA9
y3x8+o+GkIjexBNQfT+JJE6IJjPpjy9ZO80+zUUxWbya+/BjGNOQRGsvKG/JIhG7
meA0azrKewfQjhMzzjtUEX1kx3fW7/cJFwEMJgrdSPzm5l4n0gzaCC8u1gmoUrju
R7qSQrpjT41fbuCCJAQMVJIA8qpEkcVa6HZNmRmnqXdX/brO4Da4T1FZpzO/4GEr
P2PPa5f2SEznV7UVOP9thQANFvN7lKQdDtJ6X8/5SongszOEIbbhqLXoZCcsR6Dv
waXrbCxa9r5pZBd/Aw80OrZSFbs5f8FF5M9R4WSoq2f2S01M4w8knHNBv+QZQLQo
WM8WUh9EnCP1Kn/LeKG9G3uxajFvZEgECd6iKeQRpXAKv1hiQth/1rH9VsGRZ4w0
6dwndE9l4h6FHQ7EcZdvsLuWu1jG5Mhu5d8iOXey07qgtPO6xH7HA/LG+aqn/u8f
uiuCyFcYAJVxtaWvfcKNOW5jRu6fzyQ+zCtK8gOb4VGh/tm417mBVgD40xCe199B
WRJWdoeRg2zXhBqN748j9hDgKKEoAhZ4G2Qn9LYDeKs7Znb9+lJXAFMCRGNg7i8U
bBmBonlxfq8JJ1u3fjYISiHSlHq8mI0AtK5qi3CIThIFQowrtMgz+gimzARUUWZq
hfPkorcCg4pD+udnPlmvNKqql01X0igVvjeLNI6LjiqmrGSn5IDEcMKHgeKfpVdU
q/zHF24gibDxVpGg6g7j/J21ejsLBSLXJXS28hlMZqAJCTbDbBxLLvLAzaqzRq8N
dpVqA9a/M4Zdt4DcOR/t49N4pexWDqUvJHGGgVU8j/xSd0oKtEbiLE17NDqSUpzS
bAQbq43egJAHykhWCnEGv9irVNd+4t9LQ2snS8v9AdRtyiXknUeJx62GYgFKwI5e
sPNCXwnDJ3U+6+TcvBmZnk7lmoI+Wyyf2RkIXRoC1DHWo4jx9agmScifhWA20wOG
v0QGd8trwSpfdE3H/VJHlacbSiqAMIwPogpiKsYFpZcbNzIZGM6aZttJ8XX9+mUW
o6ZxU0xYZHSKCouUTohuk0XSU28kSB7w8JSC0NywQPQhrovyZQzUMbh1FFHXW1Pz
MshrosswCaSCq1af5i33FyMV8/DTEwkr7LJ5glgDDSlxL1k35D5SMkY7Q1p1jCE4
5nx/u3q65Q1mph3MzWL7l7eOm+v3ysZBoSo+Pb9ADw1Seoh8rgCKyt8EQpIoUy7u
zQqRiC9gCzuSX4rEeUeP5tD/buLzJuz0h2PiJNIfARYUlUMnPCGn8mFtLb8uqA3j
/2VD4J/EGO6PA5ShaXvcGng54L3JhzAIigVolQnO715b2USH6ytwoWZEduS44VeK
DkFr3WKR/LFj+005EAT3IHdVOEwzyf35G0kICLuEezghewGlJpBRvS1izof8wx1i
muP1dZltejZxw+MbHnH1HuJ7r/R2RZMpDCyFzVtfuo7ZB2YnJ34OyP1QXO4cN4SK
g/cwYmla4TVmOXvuy3wgYw7TD9EXFZOFl2n3NLyu30iT1Uz8S3DpqoCly/zcw4za
Zurj6DE3EjlMO+3jWCd3CLWtpCanV2GcudDFHdU+VJcCruwpV+Uk8tXnxYSr2QGY
f3pg3hTQeUDA+dMwm4n+9iNe8KiqNi0klKm8YeUN+StRHwBrwMmUQOKjFhJ5nviN
TAFq6xbJgHSJQn24ou6r3EdZR00xRLo6rxZylEM+1S3TOzcxYGnOlZz9RHeKLhEQ
TELS2NkZXwVl5Moa4sYoYqBaQevAVy9hulh9nqhx3v3GxKMeXvbFbbuBIpBlHN5z
9SCA8iatajVGqUfRyyCEzkmQwuK/nR+FxWQifvFlvAYZgSJNQ6wFxV6j3bOyyvaK
y9C4tK5/WhtDX2wb+M9urMQQbYXhE2FgnZ67RM44TQpVBUy50xyqvv4wgiZaJyZt
0EokstsVpz0F9XTc9m6DmcVR/6czIcJobQP0LJSDIQmgnZtaIV7yF9UYIeE7IaYC
/BNHoPGDqeGrO2RLGrq4F6Q8PzGWyhHL2m32Zm2vp7lUB6Jm6YM/tuyoC4gwBGIX
3qikRCHDKaDPphwW+3WCWhdZWZwmpKMx+82EeqgVN0VxVzpPn/2X1oyJ7i5aJ/St
eLLk89/cWLwAw2crxhDyY+18Q0ZwMgdd0NO9I/KVKsTTfg9xlNSjmvG2PntM6f5u
pW0Op2xvhmIj81PkPpL9btuvWHl0PBaPRFstrthBe3BvKiktmMUJrFnPGt24n3NM
TlyVHrN+/lFlfnO/EepiWz6le6Zdt5pSTN0ia0uuzmR5s9kzKt5Vvpu0Y2smHKOq
HF3D3sZvlfFtO0HtfjyioHezegHEjxjHr9hMqNIDcBe8naaM8lZWUSE6xhzyfWMC
jbZs7rbO7n3i89I+fBKahc2hqGv4nXWKKAJRMSOopumx8+SWzTOmWwr/ptCTARTx
8MGxSDTpqfP+XUGI9UNCqA0MgUWMxWILWWBw7FXDzZ1A0+4AHUom0SlqLmE8m29E
THdrtwsMu4UHXFVnDXWWSkcItixaz2S5VsLilyDULj/9iKJQP6lPk/KMd/JSiL0L
yT/6Jqe8nIrW3WGYZoZ/4ngcBA7qQbtvt6tnwyLwDoauF3libjymTCIKUkQ8IkFi
U/oeJ6f8JDHFQmjEB/QuAiikmZO0Eb0+yvJux28j5W2hlf0dvIghOPi5CoZw2nn6
iqLbbLxRa6L2+0fl5jv3j/fgB46gbEuWuJFtT7+O40UUVw9KnsJMlPecIY7XRAtT
fTqNNAVaq54rpsVaojeR+XQ60YCA0rerRSGO1XWv3nSsFgC4Hfmv9V2DbQqh+f1k
NTDrpJUJi4Tt+IgeKQUflGBQtIWA2a/mkDRBa6DSpoMCCdE5x/NJkQNtfx/TOpXm
xFmMwEjhY6VytsCjstGNppqUt7aFwBF3XqJ+9EFJZRLha0YZJeNC6vMBdeQitjfF
CUFEgAzamYSegps+nto6UvbYx5mu6VH0H49fpZXePxaYWGwPyJWg5gbT3ojrpfKZ
RcuD/K4uOGdTDdaJ1Iry1FU978jf9q9lb7cQ24jabYZqLX2Hi/OKbuviWkobN0+L
0QdE7nmutq1ArCpAB+NeJCr/rq5Rh6CRw9WO6ilDVVIma3ECpaso/bsLLMtOFGiA
I0h69LArdJYlTf20MTk1IgceQBDuvehBxeXdK0NUEb47hW6/mDmqFIUA9F8K4Sjm
agZFkkDwXVQwfmsATPxanXNxq0myMWuxo/kxdoh0mtpSfOvCrdxxxajU6O20aSUw
Kdc4pI7LgI5PUtqzfF1m8v1iNWCb9JTVgyoTP6ZD3CYadVJlcTXtInNaYlzaqpok
TCxIqtXyPM9FJ8mytzqb9PFzhMl8WMR+0xYWrQDDc8Gp0P5hXoAMVy6x3Q2uMswO
uhGOkj+Z0oqRNvaMHnoQ8zsvkZqJxISSUtG+MtoSlRzYK+YpUBH8gsl+8GACQaJJ
VLgazEjG3bhB9PVCBaLLTLtNx42t4vluj7ffjZfcgEt97Y5G8T3NBBTEKpYQ1VyR
H2I2MxzhsD20q/Z8/MvAQwI+e+zhOJTCYjpL3OOUxfd6agSX2pADdOPtKo1moYRQ
dqS1XhG5DjWBgMdb31YHxMrkrbi1Iu78TnQ+k83cbW/UtkVc4GPMTXr/H7EGMjSe
AxWp94Z30SguJLFI9O1lVHGRzuVwffJeeAiDhRzfoIEjxyg/T/iP4mpIu6U+yCRo
VFlHP1/g8pxT+sYUU2o+UU4GUxEgdp8ySrE8fL8hPGBF7KtZN7rcJ+p32OeYPdL+
KZQWl4cIti3yvbX5KH6HNdJolp8NRuNWXe0vvBA9ss/skA5+QjhWz5twVyWkkGWY
GJOzjgksms2OWL4cN3T4En1rmrvW5oM/YHfY+FoNGmJ/eVEBRTYVRx7fPZr19l2/
cJA57M9HasD2WqlsSNrZs2U98BgZ6FeTSuxh9mpJ4f3rm+b3SNkerZuGSGFsf6ND
OyFe3vaXZGsqmWfE8ItKTebh2ISHQvPHuppP1isfwdczfRZvT4NtLS+WDgBE4wi3
qnKkjKBM0MZOlaZR4S5Y2Rwo0JxMH/xsla+hJ3j+IoVyL19YxZSBDp4zmvd4H+KP
2gLd7i80QQPqs/iIeeNPOONiMCzq7tylFXJyNnDfwzawB6479cZl4SoN4SMAf9gU
RGNJDrZ8GlMPJLKYYfLZdv1XMooJOCGPvO/n+iNiS1AykGUjUTOF7bcEryvAUfUG
IJG/nyufdnjYjU8xASS+E4noO/7GBgEGvGXTYNvU1ObYXKtOLiBhLn8AJFHm3uLH
HOMRNCh9N9sy+a+HJmg1SlZcY/9195h9X60MyzUlrgmFvcmScfH2LxdgaEbQdkWt
cCOkO5j2igc8w1CsO9EyqprX/iXDYCWX40klR7QRu1USTG37kaz5ZAw5yCLxN4WW
XxTdbz06jSzQSSzh9OYnA0UhbleKosWRA3XzDY9tujmLZvB0N4x2Gw/uXZ9qdmyA
kEZxZf+PXb97BCKYFL/nLdiGdm1P6YImIgkXF9v1Oi+FbsmJAwYjiS9bVVEd3HP8
5wn0Ahtp9Pjy3FRb3OYdZsmNhuIye6r6DzU6e2ksP8emsddeuaMeLRGKjPq1I3V3
HqdTD9k0B/30ZDDeRJ4idcXiSHpuENVoEyySbr/9UCd9Mh5vk/CvDh5aTNYsox1w
YlVJbvTL0ejY5iYfsYwAQ2Ij66Wn3nef77h0f9W/8gaeotrSHAUMaPnZQYJkC+Ke
UtoNOC4gP5p+JpPGN4OttJLt+GvpR26/g7xkt/wBAGznLE63nPRatq/csLVX0sZx
6vjtbYs1EPgwZUJmCBRb5MnIAOGrE+iZHA9CxbFnqTSTIy1EL+/XAYcfRYxXjzh0
542vLuiPHFeF3mxRzDmP2YU2apvafVJAsxRvXrUKI/sgiG7wLJyd1nlYNd/keiGo
Gxo8LnglQdCA3M7Dbo7t778/yeJE6qpTQJtO/TavEMCWcI/FHUx2YCbMz0eS8waR
2Iqeb/ov+n15uKW2IvlQ5x9+uPRf8pk9DJRg1bYD/9oWIG0N2rmYBOvxTqp6K98F
VZ7i0uREyKvhEd7FYSxeM0WL22AJLGV2EOOdzHSgvN1I/kpsqo6asHi2Dfqd8+F3
SpdpmklijZZEg0lPn3b0MKSrfl76ILNdBaFFaprJABboowiSYGMdveLtgzFxtt7q
qxA3ZQQ/uA9DoA1KSxklub01D1FEpnwgJgMDF4+opN1wmvn2szXPki2zxgR2db45
+d2v521DG1qfebFVNDnh6pFVt/tMX+4EhPqBVdwl5tz/wa0v/dLuIOcT2CstudrA
Suh8TI7EA2Lmfvt8zgUKIZUFYvpT/vCIFhYrLJib1FYP6jLDklB+yQyZsiznZpe7
78M7ODKg8POHQ2tCOE6lCJvK+hza2z1+XuSI1V+oTGL6ghwDQcrs/ReeQSlfR3/b
FuoAOyY3Q5t+Zwk4bT29swxmMLTfTxhYmBZ+etsZPD7B6DafP7gnPju7chIQsFdl
UucF5GvDrjc6xOJWJT3mkOs6un00KYi95n14tDC0he+PzwHXaFOcmxeAnfFrmNYr
G9hOgzNw2azccUvHngK8oQ2GbhI3GPe9rL0GE9wZrVLlBjZKHzFtdngvFfK2gyDj
Htoi9gER1CTn4oVxi3u9HcJd7LTPopA3dxCaIpjVTjT8amedvsnFwqCehhXHUmOM
rQgXRvX26ohxWqzQvbdAIr23DtDfkiuyrOHL2OR9cmEiUunK/kZFIIru6YufTAK1
jit+J/1JRmkwTAnenLVIQmcMoIYot2pOLutWS2SWLLlwyDBcNFkj6H5+h5yvCnPp
e0uUm/cQAX+lpDBwV/bnHBZvFr5AQWBd99S2LpnSxJpXEUzumSyNc/LOjaAcU85Q
H2/rCU0JxorV6VjY+coPDCGFr93Srh20RHs/uxv6rbfieAcKvzUzdoJRtijCqUO4
kCN6YvCzPvh+2/Y0wewpVjf1axllW2+OZLJBRIEY/db/nJmy0CYq+AlmydNy3g6y
sBOpDlmYqihFuO0s511KwDJRy4MQUPwSeoA5V4V7mScs/gtAwS09M/gXiYly2V5y
Kuqy4IkVu47N8Mk3Cwn8Bq/5pOw63vqpDo5xn49j/R/V7PU9sip14U65pU+lkqZS
WPhEHY7Jhzq34xmg+HDUHpPBO3e9++IS0JR8hN1DHv0qGg623XLCQt6KdDiwpGAh
ZYAvDU0nO+7n5SVehQv/iVpPu8GIhqx6nPlbWwoqWAxE4PeDksWa/Tv7Kzq+KTRk
EpddkOp8Az6cpge//0xTw8BC0pmSqjJAiclywPv8rZbj3GVUeB/+erOv2euYG43H
GRKGVJds2RItSRYzjbpMn6moThdmewBI2Xv68w/A9DfUeH5xxYEx+HnC34ZnYvM9
fs8z4/uGpu6IGb59UMzN6Z3PxbdnKRoJ2myvE3AQMgv3+B+Bu76vSzyYy2bC4XHR
FKvwcwa7VEqOrSYjtlgGJBBvuuWxhLX5rD3is0Xs5FkGVizlp60xoEIOLnljvr8A
zO7/gKMB6UCVzay2CQbJpddzwfg5h/kO3bAxLpNFxeg/M8W9+fB1lEPrDe4MTtZC
DgRFS63urY59p1w8diU0ZH/doVHsIb9/HqUz4YEA1AJp8O5B019FzEAZv0CnI9dU
UQp1mstBnplHRamTGINSwNHUgMVLS8jVdJeEObRBTkiN4WMrneENt6u6VT4lyiYG
FY55S6O162O7R6WfgpDNRDKSaluSUwZHZPq1Rkv97sUUeby42fGraRc28gTXVsRK
g86Dgw0g0yRyxQk2HMfNKtNuPmjiudLuumY+4yFctgg8ejXRkbuL1pRWeq0+KuOU
FYOU9mLia5Pxo6o95TLxzPbyODVOVhkY0NqlK08aSGSbVTzL+bfC8g/EP74ELFq3
4cS8KLwnqKBmxspzmdRwfXusX00gKxt0jxrW7gVTg7FklJOpTGsRUpAE2rbnqqKm
0YoF5uL5iLoj5tGQ0A76mMxY3tY6+unfb8ug+p1Ks3xkHH+TZ/Fd4Sbn4Wd2caJT
p4Q9ve4yut5eAjYfAENiRkuqNKUAyL+4y8dL1wsvMo4c1YC+tRg9T1LBaG0fE6sm
Al5k7a/Z5p7BIXdAJUcKtff9hxphPZua2sjVezL679vH3skKdjA8s8AT6i7WS+s+
4Rj4dgh/moWephPeMvEReoxCxPOijwixrwZhOK8ezICs/pCyi+oD8nnnphvx0ivs
zxbUpzsWQYwk3xruBaj2o1hk0xrf4X7I3EBY/d33xQUcCA0BJMM7mpVm7VRee+Ji
eFM9sxgxpyK2R5LZwSPghc/usPN3g7lU/q3IMMwTIZhBQXAE9soDfyCUTY4ocQpC
IGGAqKzMMcjEkpNvZLeGeteRjvhed15vPO9aFsl/BLWUJ8xTCS6zavuABjA1kEKu
WHD4ADTNr1OhUAWOgCAU9vBxq46Gnsg85yOrhJ9MuBgCUXIBNXHBpS/YHCxKyCdl
bcndmq1b9RScBfkYYHtFasWPT3HN0B3Ye6o9+rQxmw6vBwRDahkt88CoBFWApfwA
nKGv628Yp7LcRIj6y6h1eoX3NkXB+4qeYyDC5uXR3WzI8t3Jsa49i/7AlgICPJCu
frFfG2Kndj8PutPom2khUfOUsMKlRXsshB3Vo9ApdvySVRklyBHzTCYgObwq1mg8
tVXO4FTifw8Tw55XvhVUVnAAPIlwDBKCRG3C0saLVm7ZvTlQUOJJQAK/5HI3uwAj
/i11kg6k9A2ISYIgQ7HkqlEG9UwngwlQeFD0Re0iH9sWv280ChMTke01sCrVmHPu
o6wrDXKmxyD2tuZjz5KVzDaW8wjETObIjHpAtr/1k4ymAivMDy8x+KoeXgp4a5hu
EudXoQgkv7eqHoGCZDJCckLWj70npvmEcMpzuJ8yN31fUVKXEzolk+YQQWwx80hi
9gIBl4gR/Tcd8MXwGrKoQ30qNiIjrewgeTv34LCibG3JpaDWZ3nkutXMeYFVQEeS
8QnnU7bbwCy0bra+PH2j6xk0SaV2vkkhqlvqP4XZfdnKopiCSO+yQYM6MOFd9zDY
EuBmy9kpQ2Tf7YNPlYq0pP/Mly41nN54ggXyF/djRzXs4xj6UAQwctNZO8vmhuJK
z3Us5JBJpZZUIzuQjHH7gpQPzA+kj7eZE6HEyyV5AyF23+DomdhRiZcAldG3RI4f
fot8VBWW3sACDfisVqY8BNuIH4NaowDEJ/yHrFD8f2sIiKuJ2AaPR/LBUqDrGA7J
6/HiYNY5P3mnzh5bcjeLkHtjDZbd7cq9GIRxIErPqFMjlYStpI43lv5+RhsB/F3w
hUQyijAmkLhZcXionXGQ7y631RLZfACkMejxNI3UXKuVmYeVa4tCwXLEpywoKEoN
+gsQRlCfS4bpggV/+VI9CBxm4MIOuqPKUaVLoz1cK11/0zwVZPb2dPDBD/hXzG4L
gNYkpHh8MamJ13Dea9cZXaXXHm8cpjVjMzep5QALW2FiNBqWvAaLbCK5lpaEV2g+
WUC6npPbZn2Z8OgIR5cKT6zMrPRfnExOMknvmhgo4pcWl1okVbzo+4nHMMPPbH3q
Hc1zEBoTQqYbr2XPlawGyKR12CZnQ/28IxsGBG6xpuaIQcLFIDuKYc+DyT2Nyqp1
RpVrFVHevj7KXZlbMyKXAxfPDJ/A/keJCMV5VdgV0SlNI8guJuqzUlizGmGjhYIo
vI5s42FwoI87AVy0TRcKUe2KK+fM2WJL8htVA2GJRWeHDhR/mzaxzFI7VmQzSDaD
cOAXIWYcgNpnGFli74MBf0u7vqupXrnTDmnEQ7Dcuf+JNxRu5HQMFvKfeGdu32QU
LcIgqwXsy+AViFegCW5zcGkSLGzvpzi64oIIOL3m3EgFj8Sy8+TG6MmK4Eqk2GdI
S8S2114s+0/vTIh9vF4r6Hax/XwLI8+RNMvxqA+78YFLxDT9qfwfoXk1cJ+3rwCB
Cqdo3IsWEVciNlJx9hldnqWAiZaB28ZK1x4WPYpRuH2HLoqjOO03eTVM9FxwujlW
qvSCmitkkaHGEdDvWdNF6vdiTS8jgEo9sJWhUIDWv/PQwKNx7wX+BCoWFq3h/bEB
IYrmiMhO/4AaHe2w422J0vxYhBWsFTE4p0cB5mHnUyX+hYrYgGc8yxLnOh37kOwq
qN0Or8KAkc+wg6Dry3jLf210bGEELo9hh2xy1YpZhXvhIMJZlR1dkOq0MkGWMHi0
RcRhvEo1FLVkUDzy53slxlhB5dp/sTRNR5f9f4TO6iCrECYpn2VtUo2NcfWvNwDB
4jAbKIXgTvfdUdrJsXoA8LkBEB8P8h4GtpCzpDzJwrXtriopHuvcxF+nLHshnxU4
tYBMgybLE0yBDElMD00uuWd0A212XzYOINddiVR6AsYT+1ezRC4edNHvBW/VSoDX
UJGoYUw4wU9YifgR19DGRPZyvLOmDOobGAmHT9opgeK1pysVMxysNd3zujkPfvLK
FwvYTpcHQeaN/WW8xQ+Sqyxrdw+/SrVHd7J8/Rr3++Gq5RvAjnP11LXAm9UAtdwM
Gr1hSOlyhuXNna8sEsJz4yC7CWhDway0t5n8qyRFa/sH8bF1/o813sRaQA3PRiTk
ZV8erg1kKPgUXpGeKD8Mkk03p+nwdHhXTxfQEXTCHbbsYW3K6r6ZMpfifX8WNMY/
VRgGWPup0o8hoEcjOZTyxToG+kLoRe6FD/xhi6/wEuWfi1qwr3RYqRw9i4uTHC/t
/+RPUD/P9Mf3AAOArjNldk1qo1VmZ2LxsJH2Ohq1fUxoS+0C5ISkxtI7Yu/26RA6
HNa8X9QVaCQcwip/6Dti9LljjAPSfEFxddOgZjSqNOOfi94/bX5cDP1dUV5Feobv
J3iiGQwzIqBNFMqsIFrnyqiHV7iZ9MJFBk5shEqStFAnx4XnkI/xRXFpwdUuK8wG
2hv2GcHH8v4rejPwsM6s6Z7JnNlfuE1tG+eES7j6rksg0JsFVJ0qdBGDwueoodSA
Dh7iltZ8GanJzfGiS3pJNdNDKaCF8F0jLoXR1aPH+hsedvDwlAOtXzCUkFF9G+F8
QmJhZALmn15td0SpjRwzZd85OmJjSJn/8slbYTsgCDvgjKJePtF9zvs5wtEbeC4y
J39JUGYcpQUyhMV7iawCtnIJpOmhIC/Ld5bq/hiFnCivk5N6G6box5vNU6kyOqap
X63GtA73qil/49oYpG0QO52HB/O/Hay9AfiBoYIftsEqA7raVitt1994055+uMBK
cksib6YZtTezYullQyb9V0P55QEqz868qUbOFnUO25SZRwepvUWh7JBPc37VME8D
iUoDflLOnsv5F/R/rZ5mY5H3vaAoCZ4gk3nXjDxQ14A0UbybBo0YVs4qYOBfzWbW
VF46DhcDO6GiNHp20ySmLWg1YJeo9hIzpZw5PNMfB385fCSum6SdMr6+/GHjtdLB
V2hLxNONp2CeU+eixepaqhJkCqAnn48ZaQb9W+7Tsr9xo6EMFeE7s16HUGI50GA4
0UvbDLxQ7NhgZkieK4IoWKwm7mtasD0xLw9jshwQYt4pShNzjSKT89rWKdtaNOdb
lmUtpUZd3LTAwX0wR5mhrKqEJ7KSdYs4EUiiRByGtxiJYkJi3PJRlvNBdBUKidaY
T+oR4eldTOTvYiVEy1lIgGuOiJDftRNqYbt0SZmxvrrGjj5wemuklbSvqzFLnMJJ
RQfEr3LrG4h9NZhuetk6GxzXBZxs7Aceegcf7icnCw8lT5V+pOtkjYULJLTsj1j3
IqzmUQBk1cFXcSEpiG1wsY293JLhDWcIIbEUVATw9eclrdLgz/5j4VDJNRfE3IPu
gdAlCePhOoX72y7+Z7GSPHMql9DUz0kkmEDtGVOlr6TaCFfRPJRk6ckHAvsoQtmQ
Kwz+DlXnoraKYvFs07YFmMTYYgr6UVb2OJTKV3FoDg3/dh6YAXd8TfahMklA37gd
z2VxsutU/lWEvy9GaAJAsPhbiBewWh1uZL3EuPy6Xe4Dq5WrzbWNYvreycU8GvIa
VagQ3jmDGuH7ou56aN2DlGQpFDkIyOnsBnqb/ZXzTN2remqTka3POigBj53tuM5I
Qvb+qLOzeg67nb7lRnoLPFVkhOPZDO8pzqplZA//0xftQvCI5MXQY3PQ1KlLmDDE
v7UyjyWFFvRzi348aAP4V0XKOW4+E7Wh4chhow+lqWjEF/xsrtIxbtplTBgchPkr
dg5JqLM1LQmRN6qLDsK7rGzv+miIwZPLGk1g5OOwqYoyYDIdKSZbwwrrpRHWsp6g
rdLfGejRU6YtZlXHvNqdeTF4K/A9mCsWYkUDTby3juvhNxTDLCsyVSqmRirNSzGz
dvqvaXy6BCrfpazdH/Accvp3ViZ2HvHwPB1zIBSzJ3dbHEg2fIhpkHpx4VKZP0FS
jO2kClmlxC4Ip5rT4mT2xlaKtLNQw2pMQWwu3jEUl+0OYSjIjBo1QKvzfRL3j01s
JNKWXkddiF4+dWczEqs/v/uaoy4KL8MEPGES8QBLX67KwaGn7DXi9eTp7H1J/x5x
C2fQllTsc8SIK9QIQD9Dtgp+u30kMjnkqN+GJ4wYlsl2M1uhWx19MWEdVOl1iuWU
zRxqdYWMwOQWlj7z/OuUwLnIGfOsTwG92lFaCguVaT59pUvcWXYuu8HJCv1+gpzU
cBUjhnrXZAcHIBP1G0uWEqY1X3+IpazOetxIhH7Tdqobj3cOS0Cgngzym5NEvHoP
Y6gw0yUc92UPa9czPpI+nab32vZUeK5x4/L+ItAkFBVDFC1MNMsrx3gSkewzV1l2
ysNjIjHC0ucqP+9ypIb8baPeE/0hUhs6ZyD2+eUcxKFd/y8QldPS7BFR5vy1P96A
SmeA7+dhlbPkIGZnEuqvjIjyhpsA8nZRO7CQhyw/RthNWjyVP54/b0RX5tJV6hsC
YSpM4HBPrM3uG19LOFFsAGmDDvG5cLfYtbkNOhFngqWEHnBc3R0lyDXV6obIYjw9
oBgYEA9YXzykePPh1HYSOHeJklJ67BGUDp1Bt5wgVfLodW+KyXHoC4rft9NH2HMy
5aQlqUsuuK5AN5Ws+gHua2vWAbrfr9c+ms6j4Ki0wLEBy7GkjEsCWT6/UN53vQ7D
hviM2+Vjm0oVGkwlSMpdZ+IPtltmlvPBJtzQhcEth2r0gAUzyZaCHiDMGe5eMKz/
7uVyCamynz+XkkiWL1XAJAAxQYQzEIZut3w5sLgy9F7qT80vnkc7bwmA4M8BWvpe
aSb3AvUDh5IfXm+hDGKaFDACAiVh1G/6waYS1zbO7DEmB8YzYBd3l3phRgXEJUTA
0bCiIVsVH5kzomh923zI3tLkon1OL8Cb/8eKkzvZqDk9qd9/rKg6Dton01+Zh3b6
ehWZb6oKDjKDuktv/eVlTHcZjgkdQOy1XeuEYopukSFGkLN4kGhFYTMptgpd9Oyh
ZNvIuOno+5lhrHVMfbzwDKSQZ5ttSYzXazCIHFVJ5xozGqJ/JBItDGM1JnfFlC0C
N0Ax70yWJuP88EXD1FDMOUM9UcPPLZa2yMSx3sESQJNZ35q8jKVKmM4oGewz1aBR
Lnq859a2iQiDyDMH9BWO1HbT+fsVK1qmjD+Irg24GoQYR19mdrysBFh5Trm6c+Ku
OndWA7HMMOgQwWKDuY13g4pSZNJjz9NSspg+AQuVCIe9alISKPgZ9qtGZuGaqsYF
a9osIKbb5/eb/Sdn1sObdPgzpwxN8kFD1c0+8NSXZL3vyS/lsljpgI5Hri7kEKaa
BrpFJmkXAtVSOxdTWTSbjh+zTcKMn7lQAlSgiNllhWluslptuQAJY+Q6kwPT8NHn
M0dgyM1xMG6Hh/jb8jp3A6AdgZi+ARCXJVLS0EA/SPyMjMgeSI5vsPWVyTsi+vr4
241FSgn0TILqaMS0fHbFff9dNOD10i+e8hqMU1wSVhUArthyVqTUsPdIc7MoxJWi
LgVSXfJaNaPzkoBk0Wp63PwBsNaqwLWzjH3ePkxHDdR0/GZJtdcfzkLRrJ9jlpfz
1Md8BASdI6fw9tfkpCecA/SNIC73vHonDxO3ke8QNTlWg6iivNebLOwn98qsguIG
r+OF/SCC3ZIcAOL9TAcj87+orRhQXinGWj8CB9c2zHeM7CeQaPLqnYQqhZhZDBHs
2UKVcyz8mtQDZaGnN6PtcQDs9GwWZVV3WBGTslgXfiA1gX9y5xAeJeG9ItVEecH3
hLsvJEzlrvOsbybMOA4FmNOp4cpOYPAjCzcWZZry502T7poWPK8g9yVl/bXoRYep
vUU2NWDSRDl6WxoSrZGyevgaxmnWPP6Qcxi5Smrht3TFEiUzLlWHYhQhEtwr4m32
qLR4TaLt2yyjNUHNMhnnKIU4/idMNiBrwwmbAPsOBKdobY6Ljee/kxDRi1slwnhJ
GEerGIk5o1m4+G+eU26M1JCfz08Q6debEDEfsSDk3ECHGLPp7InxM5m7VdrTe4cz
MaUlPxhd/TdyeMTt0Lg+hHLb+jGV3HktT8f2n0YU4moy1KaFYxKzsdanHtCB/eh+
/cRWp32SjKzoFbNpewvWgOCiBimxIyx7EUzPZoKcbEXd/TVxt8BOlpmxFIU52g4D
Desm3Vput44xeasAuFkSPFtflHUT8cQrR0bqsGnv+P1Sw2xkmWC3nLGJfnEqgi6h
Bdv6kHAz18vPpbe9GL8SFZXxRhuDCjGPzVqMaA+b8VC3T82gxnnSUPFh61qR9tWm
WtasVnKixGsGc48hwqgMXQ/hsf+P/SxfHp662GlaIJoVKo3leU9x0Qipj1ogzPMD
ZG++eSglhORVKWmXUitkBG5fK2pSze0N9jq6dfZLBrhRbHeJCRFITI8rWE6pmktJ
gKEdSYugCppwQ1YD+cDqDFcjkzhTd+bUloa1UthS5anyQD/XawXCX/qXQMgI3yWy
cODU8Tpls6OC1pB0NosZ4fPJqIeTnnI8ZQ/gEc5MdJQ8bkd9c3sBpr1gVLIV+0yF
Ik5D2uT5tuERMv+sKrl9QQwA1cfuyKO9F605/j/A4ru7EDaTsrqL162ryUwOS6Ma
QOx5yh9Zr0eJ1A3m/Iw3I2NWd0m6XiXmqMOUx83jmsGQM7UE9kSDGeOtkVfcH0oL
SK57OdUl/XyGL4jKlPuSzJA/oE2ShqzP3dr2XaxwluGIefmk3KsHixqnVH7BusuY
jsDCeOndd7uv/eH3/Pc7DuTiwFh2DqeewTzm1NiFeYQheN8d0NATanvoW8mhQNmy
zBh71SoIe8srqha5YqCjNz6PX3s4YrxTnOGOEF7hK2PKCqVAEeYBE35OjkQl06vZ
Y7GDxt/aQHojfYFoyRuXZfRfzNkDHd0Lxdk1hgCwAApXZBBcdY6SoUot2UvOeHH0
SY6JllJUDPwd9485uw1fiEDMI87zIIF1xWxoumTmmD8RowRU6QwTjY1Y2kM/CehD
KDxtvaymP5gUtAz+0do5iwp55/YNVjWjT7MneCF70poH/p/jED+N5T8uiLiKzatA
pGZUFTyjLSL52cY/XV2n9dOjJqAlTrfP4jE7tM2O22Qqm0VMMxs5S27/CxV1Hc3v
H72Eip3eeKLF5fHahhmrkgu/+BmV21korYx5Ok7jdDYx9tXlQ17W6dxmQn1w+rSj
pi7jgxRrq6QGJvKi4w3g9I1j8vtNM1FdhY+trrMbtZeBaEgSKR/uVon1f+w8Ho3H
xEF+T/+8bilvphggRsZr45Hs0Iwi3qtk620Toc859l8g4QXheDpyxIArRF1+6YOw
jQUQgFFgbpe/GrtpZOZ1o76O495SvS2KokFXNZ70BdVRGZ6Z7spCkE8+ZPjtCObv
GH/jDiwfw5GZpuj1bjgKnyAF+BWeahVle7WmGh+BNC52XSR20T+LYdOKw5QKRc8m
jq8ka7xcyrI00VzTW4qM3FFkDpvwrwpy+soCeYoSdjFfpdP6E7bDINcNvQDJnNH+
E5DVCy5IRr+0O3yWCxbSTEnUb1+DTpLb2nTx86bul3HDnIBnZNCNvlRECeou/53f
f1fxx6VvasSSiK5eTD5u8wwH5p30zK3Ftm3A7rJn8umsR9NW+8BjVpAEAY6VmNd/
RxD5a3TQM9cfxWi3duUrZSv5Rz1syQZ8NWfAmn2q7v9tp6f4swVzyGtJNxC0pXPr
cvIv4TNRn57cyYadUQEj2jtzqF7ctq2kBrTG91ovpwNon4h1Au96AXiYjj+NfgOF
K7WOLQRQt4GuIa47lokVbjmbQk2AZ3MJ21azVhsYk5qT3vd7VS8VN3UjLwMlnI+8
CHcd/U03vBoL3wVTVzFGZJs7pDOjOFJXVQV1yEr9PhsSYzwWYwN/7ni9M9iV/32J
36pgJk5g13Obp5/cJvLpTtkKkxvw0b/toAL65j80RQeAYhyOk/v95mvNqcXcxAK/
H0NE+i+rMQx60JChmOfBUiNytkFs4Y8o7KrI1UFXlTHJ+mYIyl3oyptfdWlhDfIK
ZckrMut7IEsZTgWzst255EZnzY2pOS95vi+YZOrE2loRmqhKOCfL67ED+FEqsh9e
0iE5RaBsi3EegJfaAnc6k3IHS9z+7FCQmo0emYwqQaXtK6ZyIJQ9+XaZXm35PpmV
/EkzN+zBNwS5A39b8827otIkPVWTONK4H3jQ9B6FopL6sdEbB4eUHmCFynRtHYP6
iKotqGU+ZRhiqXLvBb+NifRfr8sMzX3//8/KNsdYDPj81nQLrkd/PHsvntwqxd+h
6MyHL0eT/DUv95wa/0LQKxK1bNGzod0lT2f+CEptkPI3kNyAVdHbMFopm5Sj6f7a
+568TDMY6Fo6Wr9/xiVFfEG52QF6FklPFmLIwTcNbx6R+gJcAJNcvlgLMpI7MonR
XCsxVp42LjTYJDRWjUktqTNz0ojm1zyekDteXZVJrGD27r8LK0lAMq/06/+k5vgK
SX7tEh0+M9oUjFwropTpKpFtET0XIiPLKuGsD6Bf7vG+rcuXbfpebf/b7BVh3j/L
0Ibf30C1dUNKIC0XgkrCW/FtPJK3FB6M7VIoHWCSGy/KYr28WyAxOn4LkfgNVzQE
9aetPcwbQy+A+5NoCgS+h4WiI6EoO9/b6qh06eDiYGFbp7MQCSBXOI+6aZK5/uhc
KdFZg16ZPu2sNqaQubW6sR2oHvLYFRiJKw78MmJVTmwYslNd3joWIVqClJnavDS0
Iva0B+FD4yMSz5o+w5b5EDHaW7pEXpDjJR4M9JljmoFfNQqjoHRno1hbWXsg1VtL
l2eLvyOqnecdWBdr9i1tdgKS3TUgK44ukfPJYtXMYEva6cawcihdfqSxmSZetvHf
3X51pJNhY2u9JkgANAUjYWCNAvy/84T8AN7/NyTWUH8nVyrTC7CZ/qZ1XSxSaGY8
LebH7LCW3tqqfZjevBGjkHDXuSYcxnPPIsep29m+iat1nSTlGH+XAxwVIgcF0V8m
Lnbtby6rMJP+QLjwiSSkQn7GTa8FmMi9lnXLHN/MmSX5XkVCPnpQ13Z7pB5ZdBvL
zX+19BnjhrWWpVG7yr8UYkwmRMe/iY/+vWqXieOAab5c+CNhh90mpCZRAzs/BX8b
lq0VzmUIuV1eQid8Vl95f21S7aDjINah4aJ51A0yzPDkw0lMFzQjW7iAQH8Cmbq8
F4DXa78xI+p3j5rQBh2RzREDx59tGoZ/cbnbFJeZrs0Sw9ZYO2gu7gGijN8gtC4i
uIIWbwgH2PmteseCl/KyXljtZ0yVyOLNxorG5CAGOWhI3FHGUiChg9zULQrWfFSN
jyuJDRQqqpkGA9XStE6/WFaQdmn2lxqvAqElpVpXCLla1v1XNc0FoEiYCNogR4a8
vihE+9CVDfaHgj0WHfMUAXCYZcp/AFOgfJVrDDEyss0ap9GwHaZQ59tjozylAlEV
dSCNp6p20HBCofvACppa6gVoq7kXvpPmstNv3eEXPSCqx9CZnLlf5zP4Z0ObJXDP
Iz+FpfqM/oLBn4ZNYKc9tg1Hqigycbp6u5E0wY2M2XXEGC00kU+rFywTJ8gdV+c1
o6liO6ayEjV1vvvyN0d4jMPI+X8MHL31C+JLvJYr5I8zGZYxryjh2CPus3cjAXcb
zQywno/Ef7w1LcS8FyZ2gE7hgYSyhg3fs8LiDW4Qy9kJ97I5QlyDx2V1QGlsWpp7
fyJKsekV43MSGXfhgAAH4KO/9xRY7aa0qd2ssqqfKEEtbIvMJheh+AS0UNYGanRa
gnYv2+B/Ys35tYMGrcPJfuRry9GGQmipmWNpBfdclczeR50V8BWnO4RSXXY5NeBz
kn1xWiY8IPSFdzlybMhA1nAhyIg1EJBcQAlYi4VlwBMUbNTYDBazMbBwrg2XA8kc
RkTAvMTjYHQWB6HhWF8wtbxS6APS6L1HGg3RNesEhIC61MHtOVSZUP0YN70exeBp
ySO1Z+zUl+ambAcNgJxsM2kaXWEIBPBQHk+gv6RIT+KF7gUSxxcAe5Ran24ekONL
+HCLmJHo5viYSWAowbN9SPBtjQnIQuO0cLySjRerUYEDIWtzM+J4j2SCbX4HYuiH
woc7vSqzHJFom0EyVEOtOf+tGUfM5RSqiwrLryHIKDlifmcBrBsU1mAqzI+qF04c
pXGz6jzxlIqyhCGcEnS4daepd2DfsH1GGC1Sr29JhgSaBASgRr84BdolgvC1kaac
/wSmiJbym4QwJU1EJwxXNmQFqZu7hRfqq0Q0B3dz4lOREfxFySYuD3WZavaXPMb1
RmD6eMG9aSU2IwGP2CT0xcWwgQtPYNZz54QUDAKwGPSxJ3ngW/ZSO1uE7mbA6mPR
2jYoVI4gG65a3jnaGc7KjhuBpNosPVdUIODeDP86vNzsCvWtsVeG/NfXzvPaJ3Qb
W7Pr4v33gvn1ujJPjENGxuM1IP3o7TY2YPqUUXVraQJF/5x4HaqT9FGsCqOtx/r4
9Nb6BT0jM8t9fAjP9i6EK41ZlWX54W02GjT/kvb+t5XZLcC6y1ZMQsoGxJ5WhlXu
d1BJtw4eZohv8grmi0Dg9jCwDhqRiMg8BDMYv9ZwhqG1outA28sy/TFDnC90Pu5t
a5cb88v3YZwRd7Df6RxKINupg+yOzEMgSMeQvCTsHBZhUnEik2aXZfJtN+FwQI1A
DbOaWQSwTH2GO6rmJsQun53o7sYPRhEW255suRkLbgi5h2UNfAI3/7a6Jm6OWney
s8jSzsXNj2SaXa7+35psrttNu7fYjfCp9rvAV0CUlmIwkf/vgVXWcE/GyOXYRySk
EbjT43MqNVX1qbbiiLKfdyIOaXUrBg07rj3JI/foXcd6mbtprX3YHDX2dJEnusEu
RQUt9lNssqEWhIMSyDTBAHKkrLdZj7vEdElPOTJeeKObCIdZFVCh093yrRXpIgCU
Bxfx3/Caeu+DxdVKLHoeHtK43FbkF9EuWE/SsGspXnylzEAGKXGrPwnXAxtfdy89
KEWNzUk2P++FCDqGIc6zIVMYGJjCDuVtPZaDKXRLVsZ0wilHgpdkvIeQkSeOksYk
h5E41NmYRXFT+7Pi1STPRVawekomhwMPktUwy6bYDB47dGKW7obNVX8FHxgByaUf
Tlli5u7Hy+n9hDEOp+bolsh5CZUq+eza8b/IKw2ozxm/xMZ4wGp2kKbWqVu1XeLK
mCzjp3H40M5Ynoaw4y161UJ1v01ih2A7VE8BwjkvADqANIhX3Sx7kc1OjlNSFbdq
HLysLErYSRiQJAIV9MVkyLXoUQC8APFr9Qrj3qnIweASlWO22Bb4lm7TTwvrw4qo
asPjrVpRgMsb0f5IaAfmNSkP3QtDslyIKeTd5lJCqG972IdMsVHfRMoRJP1VF9K/
Ul9BYZJPhV2OjREcYXAADtR9l6ZY7fFRojDxhlu1v2jkbT4LSiGza6HAe6C1IW3k
eYPOJUJrCUv+EBQY6VTm7Ozn+XQPFu9wkXoiPMY/nz4Ex9f8cgnoEtV7EkdL5QHc
CVQgF9gXs0gDnrjctVPAtovT+wTCjjoqCSwH1C3Ora5N+QjXCbMtWaimcag+EqWw
kyg5sG6pSKaSj2qMfVGW6to2xZgk5/8wm9he8Y+YpgGyYdbgzRv69ZAjzzSVzHHF
aWFs5sGfOUvuSJHlAOcnRDWcB1rd6qg7BPTCQSeNWdQ0K27N1C8d4BJdMA8I0nTJ
cwTXHAj790Iybi4rgvRGT+dZTk8T3Zm2l0N/FMCUXBX9NGTRIw+MYfE4W0gf5rI3
eZ/RGSGEGEZxhxEGoerbPdYUITLAieX0ZNL2MExH+EwXwCd6SOlmhCDRJr8tLUgY
X6DLbV38E4rXycNML4LnwW8pbAfS5ANJ4zxBQwq3gsUnpFlNEFfYKGGG/o2cCq02
0V6VH3ZWIPpMJr+UZdmPB4qj5tpPhsylBc2Ko4NJHXzdPk/0x0tjK8had1q6zRgj
K+ZqIg3bRzrOzDgcP1uF9zdO/Sj0vTO15SbIfsnBtPV8Mwb2Ef58ZjkF91I1Bn15
v6XX6++btTQi2tltwYWqQ4Lcmn8t0B029Oh5RvvgrCAX2keLcmFzanthHK/GB8vD
OZWbvEGbhwq864+649NV8Vht8/2oOrELxr3aXlUC0f9cAx77gjlt1MvPu6oB2B1v
/ANNE1j1YbR/fP6YBpK94sGoBL4MBBSByaN8D7GyjHwaA18eZoSEMI9o+FdZenT0
80ikFxoUdV9GLe5NtIv6RRCwWmLT/UScIt/TwkgKfPL9afE1zDXAiyXyIPxFp1t8
GaDg2qvC5e41a759er6EpMsk5ONKHSambIu6So7m+k1XOet0DKO3XUNs0uXW9oTn
B77q0IoOsdkS/h+SSnOZnuvZU33koaePOMXTj5ciOjPS9tIWEh7r/wH7LH/tDoGt
6dTl4beLx5rpLxeCBGKXZjSlEbQnKaflVkIy0L8qKFuNiKoTQKJE7bxbZ1xFvErQ
45ZqizOYRBbeNNeKtrpbE+mQeTi9vD3CpUWGn2c8/gMHspUPJIl34K46xwm3fBSJ
zcUF9W4R+tUujhIhV3hJmjX9MTepj7WyG4nIeiqD3rnbvUSs3raKTV6Ym5GbOPdh
1Kbc40CEiNxgXP7kGOY2KAf5AX21BWvZUuSJzjnjU9yW1m+saFMu0HHk9X+Wcq/I
gUL7agdZhPbJUEqD5LMzdwAn4IBXS5eXok7FMK/sHQAnVoOtFR6jfXIz3cHQStv9
XEIz7QrbONs5gFVoP58xGvk+w/ijfr4RQogDYAVU22MASMuvYsZvVcUVSQGhhpTa
Tl8mYE4pXEUwZsCuInaU2EeNU3UQPSDoFkZjc9kTM6bkdmffFGKbuOKx2ngODX+x
qjToxoX2dtnxaJ/+WKmFnzcRjDzpbzaqhvXcKGW73lqOZZdC3PrlLwB2KK3juz75
BNAUKb4zAMlJgWT2fgYs21idNTc6qtOrO6euttBEHTgPF2KuvIWiaBrr2lgqElKm
2xs+bjk3px9mBZD9o+mCx4hZtMURs3a7yT+9/WPQtG7Bm/KQx9Lw3tEXo8F4qA5z
Y9Wd1gK2lenJZQDtmk9pT7CgclWeERrFdmuGNdu305qOYzxrtItYxFWNnkME/fiL
xW8h+YbTCU+ja5mweSBZ9ehShIfOeiT4NEqvnKHTdwpC/tJ8INokaPJUhuqXm03G
ZmWRxsYaaXvErRo56FqlktPVcHXtOdoOK5Kr7C5mNjjzKFIuEyCNkLZoimDlK1Ck
YBGwjBCq0QcM5ZiDjmo+5UqWoAXgcVv2+bTO6z1xMncRsoxUCwVF7/omdIAbbtBA
Qd+A0Qchny0+4c+UXLPj65fjiu5FO62i3G70eLO0f1bxkmYFWeQi04pz5cM/wHZy
grAJtt8aquGGa2sqTWyO9HebkUl9a+vDFzsptgjFcWBMt+s2BqYPMl9G1gVr9jWt
Verj2U+3nty5IjA30VfEhIF98wfGQd693wlUHnU9SkknmlPceB3VLh+rMO7fpEGG
jNhGAZDCOa6ecK3QX2hnPmfcT36VI/dC7PWvqtl5mDdjpmAuDt6q8X1TT7sb6Yam
2FOws3ym57LPd37Zql2TigqNLoFmxHrHwzsGB+bgswKfwQbnEABP+2AaHB0DfWBJ
U6ecBOG7omzPVrVJUmg4WqThbbhjo+6tboIp3k+TrQQM2RN3+qEilhu5jZNDoxUs
Kf7+iRnuN61SAXjNtznTpLR2/ikASJVUzCJXhj1HLZ01WpG6datkKpO4r8Iu3rAn
a8Y4FlmloI2Lv3DaJCg7KXpjBjdFXmh4yAjYHFClACKiejOP4dhp8wEn5gwplIeD
LhDam8AZm1R4I+9a9t5Hzb/FD1V4PoGvSrp1Qkad0GoDInXOvX0KraNzwuj+zTNs
9pwn0FeBf1si+wwu1hjozas1gqv6MVK0KIbheiLyJQyiYAbKTGHYtP1Gmr0CT4h7
pNXDMbj69flt00iut19/JEPjoj3p8fkj27KeukWxG6peObrS+zJJQzEUAbEEc92C
skUNwtT/wj8OQRQBQ0ujMQGLdUri24DP7v9gjS5Hs1f/RDum4I8QaM5Mm+RImVVC
oAErfCowk0Vt8p7SgtIKIsghEwcDWRGT+wuXpdBad8OibpzAW1Q4Djjlch46hWcu
kc+eTkKXwN9S0M1FPZ0an6lkzruVFJrn4tTEwiwk4TU32SGrEtJIp8QOgo39FJwD
lyy57+aCy4Z2CFpsVoBdWssUVZUX4jZKoAQqHxq8AUKcUleSjLKPLLMKoPU4ao8R
p6hsZ9U+0KYU3yoLImCoY311D3p1hzQyMf21mRa89xAuDgMbbnPX3RxEKbfgAcfq
4PKfkREVC2N/HIh+R56eHXM8v0kryO+/DIyyVt4GYBWNpra8D0pill1z5XiVFhqu
h0FiNKiELT/atQ2JQyqp/iL7ySDZDGQh8OhbFOz+tqB4bGM53gzFYSrhBEcsq/DM
dTCZENfK2wBkEIGL/VYyunaqu1Q9CLtPxgdoc/P+sYZEg1GvC7qLsVnAStZe5VFQ
JRtz5cKWbIsgpUuVKcmmvbOf7Li/HHk9Aucst7y8pfKvJsmgXhlrh1/oWSB7txp5
x35IDuFL7GskX2CcYdq/yXqG9E9EXZgC9GiQr+3/KeypQFjj+btN0hckFVfQqpjS
pnDmp3Ztf652PPW9iOR0OkQdZoxNnm5ylfvK9GDnByVfVsjHoTnsqSWBCJhlbDoH
jpAuw1rOETuUCViYapAMCRWuloNhRaWHynUY66SrsOno2TFT3ZptFit8+TAZeaTj
KC6rvNwKssSbtuA/4q5RTAb3QY7Op8rgW0Py52mCqpQoGqzeNmEoxvSWIU3JR5t6
vCeFixIHwsS/7951QbyPgcn3We+3QgFOUgvx7SFl8Q+BdzJYaetBB80XX4bna69I
rXV1sc8R1DdQHy9ifzI/28ZJVkffkR5lPNg5nEfZEJjIM50kFzU5HmciBgSmlDjt
r7z+vrG5CDfZCTXEMECioq8M+kbBH/FwEJ5dScSnlhicl6ehZ/1qaoieMhKhmULP
pbB6lXVcu3zoeIPPnykcH70kR+HtTg9Y/i3oW0wpkbY68DhisRGYnmVfi0UfNSGm
6Jvkg3UnUmVQL8vLPh8w1uTB84dVsB17Xc+h18h+Kh5v27IM481V1vkkSTAhlbB4
ZMlnauQOVcasjtMlROGnt+p+1aYG2JNOajQ5JbTRf7UVhZ6zWLnDwtU4oXhUz59b
qbBeIfBX26pkNlmbtLo8ftFr8eukwUahFJ0/r1vRkuV84B/0RbwifX+SZiwFiiP8
QEuqCa7EbAtiHb8FT6I/ASvjYqLGxzEUHIX2RsIj93MxSN1DuDlVwZaT6KSpBDwi
kea/4B41h8iUJicwtoR4IaB/JJJl5CkOz7TWJ6FCfRBibsuCzEAhvXgB5nZuYR8R
c61diadMRlKgOBvV3bpRoP5wgD8UB+dEC+lQFFZXoYw47pK86jqkI4+n0itHYm4t
dWpT7NByR8RERZ9NHvrcePBv1SBBZITyfD3MQ/+Vf0Qy+i9VFtqIyrkX6x9oKSct
Eyv3MqdIYLoRbBCurE9CfLbXqjVs5uPIA0R7kHwP9Cs2H3+bOUL7Vng6y1Vk/MVy
2SutOQ9vkDcPz1LlVnicS2HGVTUGWmvFocSSKu4r899Xt8MynzcJFRhySIHt9osN
L/cqbZTeOuZFsPa5DHcV8G1sWP14QHUudtZRBjXHmnYsTuZPnXDAsesy1qRL4rft
RW3wQeVV92NcK2TBJ5KFCAOdePMRnlbsq6xOoc73tVVPLQ5NNMuECSolGlr/BVcE
tdT/SvxVbdbLSNkZ/vXLmhqaSW2952ejc11k/8+WAuCZ8dgqWL0iS7yqZWDGV0W7
4OtVtx9ALb8bkbPMWGQSkz2buoc6WSwfkrbCnvkaNKBqDI2eiGs0g14pm7OvrLCJ
npVtONNwb5XgquModWPHgO1OfdbDYo727MP2DyQrU6zhV12ZitwsZldYo6rfUIsq
4liwTFW23rLd/W56nJm+eX+zmQg8h33jnfELRpFBsi9hSyLnyvXuVvfXwEn+fy5q
SwFFZ1HZeb4Bwj8Q+0oOmnBj10PXoYChKRJ9A9W2FRMH1v9rx3HQ6abVvX/suf20
/asPx7zNfy3ahBfAigZFJ2A+cc1+63aMnv9ZAjjSuiWA9NN06CJ+Vukavhgsj8Z3
qhk/kFJbV7yXXofHRIKQZ/m80afPiZHcIiM8ichAsJppJzzy+lY+5zYIlAwUEuxQ
0j5dmA/UYndpp3aZugS/3ZS6JtrkIcbtW62yUbt/I81oqiaGplFQTgXJz5dPeR1R
e17Ia4vHrPasueE16Gzi/0S7dRUeOlerauk+wat0Wce/hwnZghN8qE0UhM+hZrVm
xfz7QsB29jo2bbu4bLdW64qF2RiymKjCYqRJ7d4PMTfuj4WW0538lFWsncqg+ktQ
ADxnRilqalh7s3a6IvEJfaxF33r0nh2NATR00kfPOHi4ePTJhEAAEiT+qXzFVW/+
shDkw2yYDA/NbskDPQW71IOeH05zwY86c/4U4VHr3w1QylA1q/UU9bqGg1vUpRus
3vtBAlm6D4+P9FgzK5Z51l7cx0KtH6ui6Q69SD/kTNDHEhMJcpUA4zOc9t96AE3u
0tRUDtwwmlKWcVohWgiTy4CGR9h1fbsyGgmK1KhMvN6z9S8+Kei7ERZ9Dic8KR+B
Mm0+HvfrdVseo5N3DoUUCQlvsg+z5SssxtEQcOG6joSxC/kkz0jZdJUP30sIRu19
x6MoPnE2+qEy8X0Iwr8dKFCNmhply//O3DHjPlywdIlCnDfKmnyTnmxjLYEVUakH
90h1CdfFjlXbfIIovtD8LSg1acQEych5yWXcg+VlQvn+Y0bHbb9s5CZ7kH0jbI7R
LlN1MSkZ+XZ4Zjwp5ndXWEWClvGRP1NkqW+73erRNGgrAUScQg++94wfausATMKK
9EMG2/TscM+qahjPB1fAN7d00SdeN5oAB+8tM4yZasdLTI4wqfFr4zGTSh8zczjN
W+K+bmDOquplmdzlLawLNU1Z1+RI80ESKMi7zVmBHiJlvIGdGvBrXTX/byukSzp2
j92u4yG5w2Y/0OzmIsnvmHbHDuy/NHbw6vcPaBHlUBvyHgN7Y9nF8y5oD4QYzYVa
n75jQ9io7AolPyZfcfokjYw8Ll45vlsxhYusgiIl3DjtwfQwVJA//tzvQVfAC3wd
4ApqbsFFQ0JCOVdNvp0wHxubA4CLffmlqI3HwwdcFhwVY8QvNjpGvY+DaX14ymu7
Qhoz0J4Yz6KuYfd+ZUKcthtKfCXrQzwOT7XUx1x8mwM6W8diykL/JLtbAMBCHe2/
ABLk+nXGfOHCeC85DzsEx7RfvZuNROOF78Av2GHEa+FN4+I+gvyxDd9ZK2nfilS1
Os4KswvF5e9eFbxnHQ5mtKXGvMGyxowsdJPR/vd8bm8e+iGexhk2TZEJa0A8Q24e
GhfQsMjxGM1If1wPRcpNl46tMqC7SB7wbLAgm3bjL8Az95+DbhRQKG26qypv1pUS
U7qydD9MHKZSTjXykzuLBf7bqK6msR9qoG8oXkiOvr2MgHA42Pwy5/xQaLcfDohQ
71eTsaJVYEhYGWH81uYpn34k9WLVizDIPjNKHFPXkIh4q5lX5Q1uQAs7vrJ8O85i
K7Tt1Sp0zSid2cwawMICIEKA9lbDoDwd/NVV198J087mVataG3aq/kYxgL5RFSoJ
w/e+CcSaboPBfwJWfplXh14pMosyrjANupAfVVktM55CDb+D06Ug3FRnTCMLh+LY
c4LChWhNA28Xe8WPnbIKOXEuqRuVbUp+/D8t5A06opsPOPbkpHvs4zqS/lAmU+nE
YS9ORBQIgn70SX1B6xVF8nWNlEY5xInULmE2GVuUO3F1Zj9b7jfNOL8j1HALKQKQ
JsqsY7lgEoTQTRpqhiOVogeaRO9g/uiUBWo6rEW0ZG5LQEbiAXlT3BWMRfDtgGAB
JxKXy4NufhA3gAEPVNRRXfbALOtZ4GblIXGF8oyLj4CFNTYZtCtwONC+RpW2gDcm
17l/YoH2VcCGzCFgW6dEtxHM5awYA0eY+sxsddD1HDAk8BM+d9nILnhege5IJZr8
ChhQvND3p3KMCkHZSjRweVNqFcqtsDGmE73CoML7iaZsqHDTTnRNSZkoMQof7I8I
u2+iotlyvWTQPPUh+Sk/7FponkE2emP1Idrj0Dw8gy9OjQ81GZfHjY1iGpj5Sbx3
yC8d607GhwQK5PSaZRaLikxmc6ecUnfFKFZ0BIW3FelZAy2jYZqk0idGltZjytlH
6m7QTX3VXJUsin/mtJxuBKP+D+Fun/PDNzRWVsw6y2ilYfap35D2lSoHhm3hBu09
Be+bHrHeWbkaTbTyRwbIoNca6LxAVIif1F1UVSiMjH/joFnkNZpAp3xbSh7ULffi
yFQy8c54jd09cmqyLYjKAq4bHYSaSJksXbHquKYphKqX+rHmT6xK98WAH+hRsUfv
7Qxv6UFidz0ireT8ScNWPm+xrmUNKIXhFwhbzR8IsirNh2lNsKvGfrKKFiKm+x45
Z8b65tBADtnGW2WmXiAvFCasQPbSqp4KESJ9E7dGPtEQqGkLdr7kNX87Sv4BVR3B
AKapw2fBiWABdUP5zXh8lnPbZ+QUToym07I04pxGYG6ENJWdN3Ba0If6LFLzrDKB
w+O0UBFmRIEeJhlL4aozIDYn3i04fLSeFjI9wbPVL58bdPe7JNfbVrmrzHzryCOI
8WG8SoUxWlpAi30k2aPCDfXVq9LqfiJZfSoGa8Z8KegA1rcE/wcCt4tzOnf1AQnV
Mm8Mi4U9HQDPyqa+twD2xhACAngQiEeY37ckidtQrjOCuK+FMs7xoLgCHIdJY8sE
PA2hun6xZyKSUmovXjnMXyZwUoTH2DLZJdEaCL3IdOmg7yH7Bm160qWuWGRqQjSN
lpU1KY5uPfFNpHpIa5GWJ/y1QAw92AarYsyEMueF/r7+21GMkAdn3UEFVH7dqwFW
QOFP8AFUMDTIc4O4e+lyyTKeB+h2teLM+779eZzGYJZ/NPdFaJPELDnGAgYM84DZ
du9oQFGsy0ju2urPUDq8D3VVCAHLo3ZlVVu44rj9fFsHT6AA5/KoEpFw4HlfFUoB
9vz5qdCpFiHX8TdH/Z1PPsmnw+LPzr2ejFkDiQry5nI+vLoR3qmD/uxKvp/roxW6
X1Z7Lhx83iV39ERQe4zyyPU607INuvqFt5RAygIR2Yn+OZ3e2A9Spf4JJGkd6jIi
/mKDiO9Z1X0139nuHVyImEtqh3GJVlIm4zFfXnnZBHBZJJMZSGbrd6qFRk0hhFZV
V5QGoCDCAoLqxR1qjfFAWYHyyDGC7JAbroBslGC/wSTuU3p9KlwQFfk4V1GgsLbW
blm58yiZwCio7Ll2PB4gMJI7WyVVhSqZmlFlLCibpjsIM08u0OjvHeBD2pVCWBYQ
Sfw4Rt6Uk/2CKVCfWU1FNiKyNpiRfPc6XTAhsqgyoljsZza++wbedNOQ5gF4Rv1W
+BdIdQ6IQ+nK7LtyaiZTCMNH1z7ZAoTUGT41+Rh/rFVAzgbxuoBp1JuWnU1+DGvp
2RC0jz1UNa32XBFk/BRpEGqjIQsKbiUIgMGM/vXtIP2suLHxnrgNQFiF1sFN13OA
UW2cJF7vDyGxPUFfbOV7PnpU0Cv9qKIogFPY7iyo9lN8b5KZX6IOJmNad1u089pg
jz0Q8L4bczOuzQb0sAqaYAUkKg4I9W5+06rXKsx4YK3MT9VUNvvnqqNeyVkQkDwo
lmLqz5alqZ+fJEd9l1xp0BWIRodJna3gSJC+YQBsWUcH/FFMHLNlDrvG0dYCjzlY
hqCUxP3rFyrSuj/hm/PzHvTmsfKnTAlYxqZ73+Utq93jgizOfjefLlRxqrNMNc2O
ItzJBjrrvG26pcSuh49bgTv3yUDS7Rei2tG5S3eHhRJlnUKjhCgzh2fLKI/W5vM6
1OCuzQ2EYWy/kZe2kl1tYy+OAKJqWh05kB0G/Wj6BMO1hPO8ggyMb3lEj/lUtIMs
p7pg+wcEwftZDR8gv5bPcqutmcAg443QVCviip/wdImMcplxnwumwZl9P9+c6Q4n
TtN+PmzdS0zyMjnmfqMVa5EEbciLLSIyrE7/CS+Ol5HSpo8PzXXcpB7r2/FjyIZY
xN1KhY0bZUcAeAj9Gk/788G/jyHSt7wJOkEV3N7pJeT983cgP2NUhkO3kq1mBI6V
fT2uqWJrxRoxjj0UFtDm2G6gKFmR+XVaQwGOamej9stmeir3j9LsMu8ZDPKIp8bO
UdL5G57X4owA4PTVTdzzV1cGXhXlKa5zDfHEzLFjvitJmF/2stvvV6bWMw2aOXjM
6CXEvFQI4yb2/i05LPhFonyIeR2c3VMPVUmaUNAeY9vMpmdLMrJi+x99pDoa2as7
VD5xlP4Xrwu9oUt/BF2x9lw7VICgFwcMbVQ547ZGIvUQFSqv7Ip7bV7keXWLVTgf
xwFCVY90dW5vBxbs1IhmNDxawP1yDHe3t5IYjE8bm/QrKDRV0iDpD88dIxca2MdH
orw3lrCjxg1nNNwGdyBuzbdmiLLNE3KkJQmXltiqRw5UIqkSYhxGtVqjSZ4PcSwD
Q9fHAR5h4b7pEPanMOR+QU0lIkUDqDJZ7R5napeDf3U1ndWLUUY41U7mjjKsV2TE
rv4s9BuEJer7pG8oo3mgchcV9ogFApup/STptaf6fGCP2CzJPF+xpLTi9Z2Pa7xk
QI3VudS3oV1j0NDVqyb5/Jc2JtljeXcPZI6+hddOCf91MZNlTnAQc6OBNQyJbUBy
FGG+kzj5mpXCe3yVkz2QHVnX/f6Q9MMK5Y7IF8jCPKZZiR/EKgmcxcJEUdgYw/0v
RaeSvlxY20iVfupEu251eFVk2kAHyKO1Q2mXenXzMFmG6QxGe3lB3jZrJBSS+3g7
3rGslesJBLr/APxOb8T0AM95FzYY4H7juLm74JCD4hadkwW9WY68kFOc7OyzUC62
iQPQarlzghOLyo0bhtI4epmpPyR5ri46i1dTm6bLbEBHcz6NTWSjQiR2KyvW/XyW
EO4JUTxIE6ntS2anRq8xxOYXOq39PHv8qn1mx17RRhLld9WKxjN3L6qOe/H7Sgu3
n7oP3I3HYtCH6o9E2V92CZX1NBSouHXpwM6WeXaXPWxhQsPci+kiCtdyNCNWPq0E
PXMeh7D7G0fFArcaeGuvDUI26tSEAAqoMogiFuTSrQk0RebYyrdO/BSZTbrVLl91
bb5GnkEQHoRa6xOKs1n+7/FjdscmORwpXuriTFQ7mC58QdlX9UGvyGHI5Hfpt/CS
WW2ld06RZVjvvZl3dluzWL16mV7QOP/tcrZwQpGvm9Bg9RstL6tcdw/OiC62UGOR
nZQe7SUOCSm2TRHWVrM9+asA5zwV9b2SCDN06g8uWTcWqCbU+7WFmcSP+rj4a4tP
cydy81NAwQ0w6GaJpC8q5YtRxU/BM7z+6cVoWf3gI8dN5fMvtsVGW9IcuKn5li7i
/5LCDtAAIGhIwo7r1/g1Kk7TEy7pbWL6kqoN4f23FKPYG77bdyAKv3RFRRjZtt/g
srxqTJLjiMKdS3NdtfUYhFl+Vq7GmesVQAZjesB7/gma+xQqHZcdditNEjkWiIBG
UBP0VkK35HwD0pL9IlitrzbzBb+COkfU72+bNyucBVmeGg/o1klSBXb26FUNbfa0
oRbvsDHx/robYQ2m5TtXnF9nEYaY15X/WFHVHLsLtApS+qedHyflGCjqqIIp0pDL
Ic5nbnJLvJpU+hZFkIfpk7BjoIMC29yCb3vyF1DvedPLnDGlNEdqXRYC+SqM1fPv
B9esMX/NJjKUK2/F2QCo47MsOm+c7o8Zsuj29xGEK7XcP/kNC2hdQE8tnVI4HhF2
pJcv5MhM2QCK3ytgT9IPM4XAkHCPebZNJ/ND+eNiMv2LSpLU0KdJ63JXgJsQiqFO
KKPVdjziNWC+2S3gTep0GkOBKdorfyOmjFiiU/AbXEq0RvF1+IveH1Ri8T5enkG/
UJabJfIrpSUxh8QRCjY2kqcgi757gcS7D+hkdAsu24H6i9FQw1i2DTAGS3DQ4unj
rEMmQGDrI8w7CK6gdiWE9KIzgz0AJK7X/2onZLMGaP6R7l3GaFYYJQSnDrcVGZ6U
5B9c1gbQ3gjISgRJXTt5BTQ+1e3EtGegXDZtMGSYPTMaGnyzfoCz+5JR0RXgI3SF
kEmDNmxQF8jK8ImymyhWPTdLgBQ+NLwES99WT4DbCvk2YiFkBg+zdAnSwPz7prkh
edMOiN+xLGj/qeXvhLKGf7Ve/20rPmw5fKaSzLx12EFmjYnHPwj9sDi/pTU3plS1
S75En6v5f+lgS2/oND9HMtnP/879pZ90iG9OAP/nSSW9jUcgMoJefPCiPF+DnzOF
66iUM/T16lYEGIF1uwDXkuosarfhRTOFTlzei9V4BGF8t1sEjJV3uVvoi7MOpwB/
Y9GkaNUMeQ8Gzo8F71Ekk8hIEq1BMgD3E0m3LGfeSe6KRenSY6PdeHXXkZSpxRWi
VRMnq6XPCoOK0Rk3Cin52w+8RWyKA9EjrSq/gZTtljhp1F854M9ITOno8lgRZVG5
hDR/Pz9nS4AUBq2T5AvPyB7BemgBHNpTPm4DG+hVFNBk1xhvjio9mNox5KLk/mcE
tvEXNIH4nlOLoD4o3CSECYNelwMDn2UNHM8XQAbK1/gcJokasGVjWFuJkoCOAj3T
Rq/si7w/KbBDwJKu5WCT6jSPllnYx6SvMCuLBpLM9aZtcnJtmOz67qyJ791gMXoB
dNQoXYXJe9niIgKt67xroY3OhkLPvhptGG8QiGTkJDn1icvXcbDmc3lknPNgpSGE
z9MCx8LP7k+yMAFc8rMntrFRq55HvfeDugUNr0q4wLeOK/eOMmhPIUsPgaaLdidO
36H2ffnfD2kqoXOdRLXl/TWjxaTFlxbA/+IYPy0jUOZYUQrsIYWjj15nF2aWV4ON
Yf1swqF0sompPaeGWffeUf94K6akJs+/p+8o/bemnR78r1QbMArD0ghY5i4pbaln
v/vq1VvKg31d8Od92l39Tq+OoN6ktYsO4fjo8cV4DD29aqZTUoCiV9Rz7c2D7RWe
hFYu4D6TTOgT0PiTR+US/G81lDEO/kSadQ4yIT5ZF68NM/NiQCi+ayltApRQANGL
HPZdsCd3pGSP1bhI9d1KCs5UI9sjWK025U1uYdbRF+UBsmouTZQ5JVpbKGVkZAyc
ufW8S/VwSvmucOE7EzVaGc0a5TvL38sCV/sWWb1KR/0v2yWV8rogqhOR36JSOHrR
s0ar1QO5FF+JOJFh+N2oLzY4h82Lb7P9JlqGWFrUrCGtHGpoubE8TsBp1Y6QUAar
3o85nhOmJqM4QTjHOtjf4Rk1TC/1fzx6pfmq5S+NNStEcgsFfgMzYVu9BUo6kc9u
fUKhpcbEfUafoVjGKpZiB09QhsEK0f1IaybxYjJzza0IhefcVXXTyaweea5itLrg
J645tjhP2trFPHeZnhmSGFfEPjB0Yx3x0S3LidCFclOb6Ld8Kp+p+XII0opO+rrP
Nrin9vcQwovRciHVdLW1WGyXGEmqiaeAobae+G0loug+/2VeKFeZs3jx8lwDzO5L
e6hD4viuLhHtZSrAa5rMEuA2pynFYxhvC0SyfGOUX/F0Bw5rsHW7vVnkrno6EJRb
2m7vLydZiqshwwPC3vVG4Yvo6V4M6+w9QkwlnhFxtsAyrgRvTOPsQrUUiTQsn+LR
UITkYYiHmmjvS70Q8GXpa4efoHfMvq5NbOKxzC+EToxwf16Fotq4RAr4KOvMJIVk
n61ah8hFc40TFPXBNItqjAT8mFO7Zn0E6TXnB+NPBoeRgMRHhEKlcnkBKXJMrdRn
5GZhWmkRxOY97fVERuhS+1f1sZAltvkoyeg15XzkK8I40R7Qdfz9TYrXPHwjTOjW
Zc0JiUtuV2mpaLtVvzQBgW7VBDGWEQYHIJO6BWDbjhrIg1h4PA9uKM8QOHLMQXy8
BcfwLgdPCY+fkF4jqRYwZcIPo/yJQkMBFpbxsHRoyNgDO7Sr3+aTKgZB2rKfN8cv
2AOSYhm5Sp5uoWlfgE1F6Fq8vr3B6MtuRqeadSToBq1bM4ZtPsZVu9M1Hl/Nytp7
9zvfQeAQg0BbPkfvxLP5M63zS8TxQtrsBCG5NIQHbF22XhMPusQgYiwNrISyNfin
kbwiIUCJu7FT3Ymos2blpLBO1RSRUDHufCWwNW253ruJP6EEdkppCusiIKkygwIe
kgc86kC8DLjUEyIEuTfxVrJI5bKubduJO8J1e/0+Jh4sjotQZ4WivW2SD+ObdHDK
ecwsiRCyf9ED8aU/1tNgNJcov20mDCk23W7PVMFtamTl9vk8eOhlTgOghn3jznCg
L3+QLe3PamPean605p7WBb6ugshOA39vI+3Zmo5pKzr/xYLbjQkJSFCvArxGx8Fs
2gmr50zT/hk4OsvrXuLkoTwMaqZp2U/Ijw0IwtjdFR6kUwrY/9h4FTSn28MD6R+Q
rZkweKNkJzj6bG8NSJg2GaDRE7nB447I+iEWBKThvexZbJ3gJhpWDDo/ZcUKhErA
fSS52HRPcMgnRvO57FjAkJ6wDbl4WoyFnOaU4TdwgtULFacvoTHUSc4gkFDd8IOL
k0C+8Xvyfpc26bgUQUn//RPn5OG6cSq1/p0MYFJlo3qrXQpzLIs3Z8IKxQnSX342
BT+PZS/3bhn2ADphOA6m6KmCqDlXOLSOABl8JBJQ80abk4xAmcuFmy7baxO0SSyo
PJqjZB7T9rLIzYVL2vANYxVei1ZZWbjzpfCsHnEN7Ra30j5y8kFUyilD8wGnKxH0
Sx8pAuKDORhYatEtx4UvDJ5rctVUPUrlB3LOP+sk5QQTPeNqG5wxkBr2UHcoiPqI
9ft4P4HOtbApDUgfefoPb+LLDLgJZVkr1RKklwN855soXG8YVqf63cZhl0c884gR
eCEfCueH3sJ3Iaw/ne+fgo14Slvx/oF1v1KiENyVr7N9gOU4iaTXiV5Wy8femj+I
qCLvtNb0L25Ejiyjr6uwz/w477i2PRbUKm3p9VpTcZlhkqyAMsFUoiWKkfln+04G
ttTgfpoIOVisWLbaVRQp78v1zNCGwrOCyLiQhkDUePfhZUYuCFOriouwmMeJ0yb8
Si6T3NvRFI5rU/+NMZaEePUgbBUq8OU2NWAR4bT/rnNfMxGl1soD4d6Tiuoe2UZw
E+Bfg6wWIK8ixs/Qp5iDJatV5yX5oPJW0UMjlxA9uQX6JiI1kDIEK7pVOi7eOHT/
S5mjyZP3F2urz+0fjrvCmIbZ7+Zv00ccHGdJzNAua5ghNphvmdbIpzv1K2y1GaqN
bSMf14QzBifquSnVzg4B+0JmtujK0VVEFkSO5O/OP7j8j+/PjY/sdZAzE8GUOCn2
STp1Ii0jCHRhnb2h5I3ET8BGdfRLGwCFinVPrlZBGJYU6OauRQ+PcHfixq1Mi/Jv
xs1mwUVSSV3Pfe4ZKUXOgc39KMCbcqrHZOEYub+ZY/1B5EKKPBTzeZ7f8BZSw/dQ
9iGJi5a3xEfMTC6pfOzMxVztLGl1rd7RHIkQOjpJ9K4EfnCdpvt+xyWidrqyR6i+
HH1yQI/rbJmm5eEbbt+ZECDtn9KQpRfachCwMLxoExYq+dbkbM3h7mB2KA37gJvo
qgJpH+JONSB/z+qx7ph5gIUMV8njKx9ERW1PELHMkBKHFichwtFHSQAuUjP1eOfU
r6NF/eNV3zezxBUu7yQYX+Q24Ot079OYh19rYMAHezu5maPET5R3Gnt+HO3BflHR
PVWfopKcZimjHnscBv3IrGb8UWnfsFVr6RYnIvLZ2uJOapiMVlGVkfA3GvyRAubL
hQyyzEeYTt1eXMtJ837+G4JnlWHlkyzTAnUXF0gXLnGn5Is9Ow1PROiERq52O9fg
lRtYBLppVGMANOtL+Oz5/hP8+dT60ibF583JpxdwvR2z1gbLAZF8x1qPNCOLo8Ic
DhOWq5qEepCyH8PFK8xZ4ykQ1qyBR+wxDlPsXlzXmvZg3/iCAABrYjHs97nmhb1z
zINvSVqcxvWtQW+pLfZe03KLmdMYIkInd8V0VIEsfKudW+jNAqH/uLcyA4QpG0OK
/Bqx0HwPm5tMk7rcG7b96zy/xRhb2SrQxgOGufWXNaNlhz74RL+SUN5nU7OuvDP2
uca7nlsiHVCE4H6VA7KBUaA8JZ0WpvAGHnYTD8owclm+3mY3FbqGSrFpg7xjXZ57
xWeZgDpdftBDsd1P7GKl2JLK8xp5ApKXthq+rxoa0+0X2IK0AsXt9SIYrOmNIxvO
CFyvRSzgWGwapOvCgDqlozkKVrshF4DyataW+HTEYHvGIG23jmIzsfI3XqlkuXJg
MB5a5rd9JCXSjCJoS86bDFP9XDZgQqV5K1BwxMePheD/ghXq2hAwxGf1hu9GjN1Y
b7DbQduYTpYQyJQu98FJ7FkTRa/vCrnU4ir5CqeiGIQRdZGDEFCZoCeJX0lcvYuU
UEmiVHUw3ixPBCScgAUxtdXPSZo1jOm7S0kcFariFw0E5oY1Sx1XjKZpsM7vAnB2
1IgifAHZWK0NKwAte4bLG3ebAYaAzS4loHwk2dmBxceo20a04RU6Tld++hgPHi8O
7hM9tbBc85Hc4CuXRtWqp+3Uqdjfmfo/cSEtrwaOpZEsvUMS4OBs5sr61BMwL08N
AW9qYAXHPYj6NuFnlB1kZLr0y4KnPK52S9YfB0WCXZc7UyH0LwKXbnDSVRkWBf5u
H4ZG9yOGPma8FXhL84QzZlSzgw8fbTGFM0QZnzA0UasNu83AUXz6qQYmSDHGVBUV
FYQ99GwvWx51kuINWyb2c66UCHTKitJ7zR6AOWTO8jZ2FHZLc8nxXraF6OTbza9X
2+15bFoevC1S12S8HtHuf324q7oYhIoyOfFCv/w+s4UpUf4QTHVa3mnc4f8XRJKz
OA8iMJY+TI7oUocEuV4/A9uJTqALWghS4UVHy/d1j2EvUq+i9FHwbbQu8ELUYLoa
U6pS4jx2GemWBrcunwZjRE+fAEYGQ36y8yGPKmRm+3pndDaMVZU3ovcSGCsuoI/X
KAHaCRjPHkkPn8fEDXj/VlQYo4/lWWeFUAsymq9bM4n2VxfTF4jL3+J/cfd7d4xK
qJhSNuKJfOLNdLl+IJfpLtK05yRCqIwIBIKv1W01E4P7VxGvJyBBSAkpo1bVOdWg
i9TQ9cXF+w4zb9/Sn6pgS7tyZSyAtWpgMxEO5xddrL5I5r2nvJJqfUspjwbS9qr6
GzkekMYeVLjAaVKdIRVSYRP1FB8RjlitexGw+guFB62oxJbIDEYsKNCl/8SLIPpp
djw8biABE0lxaFH6P/EGKACRydU21OMNgtQ37QuJEITSGxmcizi5Dr6Q9AM2DYrA
Pj8KOtrd6kymBmEg9Jrset/oEZ0jADd/U5yg0xGnwbGOzkWNgK/w6ffDP1qNU7gP
Jl6jX128kPYzvd/phCn9+4USQwtXFU+9glw4vBIDgKYB9SMaOssz8Ipb8VdTVhvS
fHUkH9Jq9EYnX/7C8v1EbtdyMXi5CSpCMjDeJG0g63Km89xkCrDBC4yzc/EdH64h
gY0rnXnp60V3A3ILwBNG5Nyte1jcXBV30HqrCVcfr8LjZF0zY42P+uALl08shcyK
8sItlZut7uw48agb3Q7sQ/ofi57VwIvWOnrinjWZmCX1bwasnx6NrtBhlOwcSYza
zXAtCe4Et8tFvmoawU4hcT4js1QzhIivFnC67T/COrROEmCDGVj/Aly/bYK/m+Qa
HFAaUeWPT6K2AcVE1x0KTm/OjuWaZxlBXvn0jzD2FVk6c1RE5NKkDjlOSM+yqpIr
2JzL0F6q7LG+bftNT6SQx25VgOPZqV+9jmADsekNbzid9UpfLs2z0Un6dnTLY8x7
BOATrpywA1I4ir/lzRRBbSVyC5I+O7VcsmVwUrjcXpMzbth0kcFki7oACufxnFII
vZJvpKSdONuTATg2SjcECGKksvZJotUzMtllf919UbXgD3y781iZmkmC/Nh6b0em
cjlayKvdhJt1YV3sYYt1NhfFfspKJYduP83wCamDE+rj1chXEoSZ6N2APh/otZWP
NmyUZV0Jxwrv6GFRJgjG16OUxq28seQPRlsjiMNv1bHTG9EFG2zv1XTgY9kQZh3I
yuWBtFWLAHv22r0bUV0Uuf0100Y27/yY0DqQ5OhUdNLU33EZA1koYuUhgpb4Zmlj
z/eECnw05PG0OJD8Xu9omgBUdtIGOQU6m1kvcrWfKQEQCc/ztxPNa6fe8wMPczb6
Vq5qLTJ6//Q/2QzjwQpLI+6gbHlS0qor7TK7OiTc1Y+q3QcyCAhVK1FMKTNuLjS8
hBCJsFvvJsMsTqc4OeNTv0AMyYr4NWsJu4FyXJhTvBeba85GXsLqbJyOQBqQbA1Y
yhj9bsgsgyYQ7vAHtLwVmYdCufnasKtY67hxnDGIEx3sDL4UKthTDJpX7Q5wx662
kSEkhlgBYpc+K1IwmUj6AVgCvFTUjXcrBVwDcW7Tiv4w6K7bdovwNGrNTXgIDxpc
r2z7j3bWpKEk7EHymlN2gL9NAwroqBKBP/kTGk2YDmk8z2EhYopU9lCMjQjluCBO
h+1wtMy5FOs0DfF6Z2Bg1+JbWXA/lsHL+PmyAo2ctBXJj377UtW7YJmLQWrSGJlM
Mf0pVh5QpGa9Bei8KaPqmgXwEvPewV86JEvFyluIIOgCh0QaUVu+KHy/QscyKf3B
Z/+WtD2jJoxamZpd9PE9SHCndr3UqIffdC0Fug+ybAsTYs6ZWZaBf3bP8OK0U0i4
E8cIPWLAkLfm0BirNVNzhZevoMhrtnmgq1ireN+MiEUKoezs6jz96OE7+4N8pDYH
n5y8MiqcTGgqjDIqBfS+WAkn6PoVqizsOgz3oNU5/iEppBGxBwF9Eg3QT0r4/vmd
JFeWKdV9sOlC+pB6Bcpp1RivgBdbtQJbnuHO/I0svvT54EMwIEkR2mI/qmej9HUs
v0ASS+5xH22uywhnsBBVkash4nz1BLB5mCVveWxQyAomUZ6BCXCNNTzPOePpx6vH
83xKQyOTarvs3xfYwDklT5FHevGk4o6MxGaDaLTgkiC6GAIwMZ5/bfJ7WWAqdxgt
Jw6gbrOB5O1yX2VTadt66wfSj+HY+zXDSqn1XhXgD2qd8qz1Uuin+X+KM7wzeXkn
cUckShs1zk2wDxaB/uETuzpJ3r3nL3vYC+d2Ln2DMSXgEIBf7T083cLPHiXuPna7
zOfeRVZIdUW6WIOpuTbnLTfNPEmrOf53Sj3zb0epXa9MAt0yqtI28LcyWDiwRY/l
oAgPy9DF1Fy3zoS56fg/5Y6MBRqQK3SOSp2yAhsGDR0PZCo4LlKh0vXuSrmIC/JH
F9ZVj8Nqrap1janyla5mMyM7MYO5rBoOIz5ajaDWmZfT/E+faGxycFzBFIhbtBgP
AfQh9s/aEHx7GjB6rs5aKaCFSJz+YkSHfz2bAO1ROYWAvZzAB7K37tyNkdEmp+s1
W9K5Shm1eP1cx81TGqeB6TZhARs7IZHOTnJ3pYYYD/Cl5JmDtrDMt6FqRn1U4fN9
n90VKssnSPhIsXzTM5a6rPCxC6MMKli6Tkz/sHHLYQAmV00sun2NeU9AbBh2zvlf
CxHcnwjHYxd7huk2lBWRXDnRTgjoTI4eD7SsgfJDhZSc5oWNYl88EZlf3nu838H7
QfNJ7dltYPXksQ9cSJnUkYV2AogOk0eoBUWOJse2qWmycxFB4LcWW8AMSnAtU+PK
JXN2YRQj7vRimLEbi9DvYxtyvQntGhUdoubGbXfWZvfRHINBbKmjeKqWmXRz+Sqd
12BBQ+fc4ZpE65soc/76weT1y3wUV3cqrtxTe1R3n4qe8D5Wh9Q4YcDl5ibOC/go
wLrx8DZYpFjhFMT/EzqJg2NZ23YDpjyRgupnS/Q/3AScQZMjTgAARFBJy/Ym3aVO
ukKn2Zc83o5mYpxTkKrBaknzjKDSnjgX3Aj4DcygjrJVwfQq0MbYzNT4TjR0tlYQ
uKhjpdT22NRHgCEsFYolRcZ+heFOdMItZjPdjA0IGiMA9u3zuhnsPt0TTkOXZeSe
e4wdlE6BSKtRwhCa1NNk0OYGMnfUqVnUSFVOCa8sUw9GkEGHNTJrrZR4mhkP5KBl
mh1H9ZlfPLHf2uohEHqh1Pmes2KMChAAlJMcEfMissofX7zfcICxUHAxpMaWYR7y
8dpxsCsPehwJsCvCHfEoBfxmgN3n9PcqONpnlFSl8lPrlsHIAsyv/7XjYjfr8PTh
fVLy5DZqlbRsgBWmq0lnlAYqwynTx8vAJv93nD7aKbZN2hZS65EIVEGPUFkIlUtJ
XBPYo4KBJoHA1jgVO4yTHbE4lWuLiCESJwwS4VVRguqAUqPXNz+HPYKC1VJe0ql3
waTabs/yg9yAiXlyWsqfMy62ml5s/uWtMYw5a66BaMIDUvD/+1vJGOHe8gIW6kKW
uVeeGFmEIxsy20CevWVPspa2W07Su4V4KrlmcSMCTkh7G8f7FB1/2ZkN6Hv0wDyn
ydJFbjdUQgGs/AOz9cZ+/JDsNSstiN4458PA9dLI9lmVLfUW6T3GCSj28gNrEO+m
mrZkYDwAGDKOagOK8+MrZwzq6O0y+NGmalxggO16nPFmO0uzOhT9ivso/3WvG7J2
5dURT+ifqPGCLpVpV1N2BOrJw3ITon/iR7amnfxCquDJMQ+wCgPyjdXhy0b1Ya3+
GTpr+4ZXDroJhxdChyUZrV3M1i3hBqF7PzXcGTb6E0iwtycbDAUWRcEyTJpo0D4+
XRzVu88w8c1t40i/fl+aP1Dm9rI+HunVkKj/tt/tUeCxijdNQLqKbmS0UrHI0lcC
ZKAHZQwykIG6PBwhIAbUGsaLv0EsChJ7Xi1lEY1Idfi+C9HQ03Iw1CkF0mRUjdPZ
vLx1aiJaB83HciX2OpDb8tTilfDVddWq9twRnk2fCzMSDhOEXAyv02z8KjJSsiWF
4EiDwLns3DR5VqnQD+pL3UzzFXdshoscZK1PG1YKKHmGw+SIbm8pwAm2vpeGz+rF
lOIn2D/4zfcyAK34D412xp9nPOBm7pX6hFfY6wmAvr80R1cCf00J/O6WrKePolwx
Qvw5bks/BHUQXdAylSkLDKVzWZ7zTzSCsBjdizG5f/4I3buuGGwrQLkrV4r6NnK6
Wa/LFv6WvAGqz88xMmflnmQrLSgeDnhFX3SBgQlu3WwwWjoas64Rd87OeKwelcQ4
gCCT18wPX9vgAtrq9pXJSUKbQpUy7WhaJZWaRR9wkUWU7QhDD23t/18XXklyypj0
cyhNiwETFI4IP6ShpBIdw+9X9h+PbVXrWVdMfghNGQwQw68NtIM6wgRpjYFFxOl9
VJmH5qNPoLwY9DsGr7GX+PMS4RXNi8XCyEolU9Ps0Q+6hKqNzAPIYpPBBcNFHFTU
82ZQAFMJ73jFdxoubZ9yN/WXpoJS+3JtGpRmyrDNm5ag9+uGmXA5L5H7jtDrx2S8
E2JE9I7wQRG0QxwqK6XeNnfXy4fDsTn4NdR4MP+25iMVA2UdfSJQEr3l0uJRqPhs
0Qn5Xap7/0zhyC7wz7m15TkeqaJUrPG2flJG834KoJHxlH2/18pWsRT2HtCuFXJv
ePZ9AN4cy2OS6xnaj4B8MquWbx7Vr8OElJRSp+6Xp6FBup3YEVB79NQvQfJIhUy+
pOyJc1CwpeVEoI9OUS2oUkhpPXjVDH3uZbr4B7Rn0re+pionuS6XdfPHeHwuY8Yo
dkPY+ZZYZpyLVW3488cRT4Tsz2FWIp+eB5520rViOSymKFYSp3o2NeBDgvUFfjZo
FaHDOC3upsYzV0PS+CGmBIWJ8Ef/aeCiXlK94PU8wf+TgItEdO8cpIrED70IqshT
/hQGuMK0QB+Lp/HPLlDcuuEuFY+TF+bhKcs2l1K6HJrVgmMAxSSJRLbHFJpGPVop
1gSC4WgmjTh++nhbMFyACr3fQ9F495UegQ/Wpme1bqGbdyFL0s8S/i51dEm4DnV4
hUgs+5Zgm/3QoAALyoHq9ELnjdvGgJ3q4G2mKZJyuNykiCP8PMjSdTn8C324S0Qx
5BE/OdLIXWTEZUYD8sqsOmam11caSBfgiqwm0mRtwwSFe5fwl+PLm0jymbIwURXS
M+Wy4YSu3UB0JCgGC9h769UiCwWVdgcwKipUhMn/GwlBmBJ6vfiUS2DkYDWcoiK0
is43nzGFc7czyglDRSmq6dFLTUJFhTuJKWAXTB1Yz6V94UUqRUSG+onOW1Jj7oDZ
TU6uPNf4KkqaX5t+LyIpFd93rkd+l1k+XMnEaHlRdkcC5f0+L8oM6sZiM8p1lJg3
azgZqB+/avtqMyCofHT/+qtBx6orgUPCvoC0S9tqJ/yJ0gDKH0GVkYR3sJONKEgR
+gME46JSfAcfzciLpGC6waZGPZm4GeAAXcaaGKLZMD250nE51hWm3Gdk14sy1vWC
7PWlBDhgverwIemb92oFdZHrac7Mxk6v2R3J7ajDTmEFQ9kt2rvY/0IZatYQ4yTM
ipAqg4R809TMO3mCL5LCI3D4PZvSTPIr6xSQBaB9mEV3JB4PRTFCJ5cG6efUE2pG
Wjp92vb/jV0Yoj70itoiSMeYAoIBdVurT+WWSalE9iVGdTTpj6mprDHy/oNBmUzT
R8ZlZjm5d8D1asiWC6q2itPryVEdZcmYar/mQwXsGVRhSbQaKthVxbKaR0Mk+z8x
x0zOwUDwxrANMiQxve2ZT0zWfpUwhdOxqMvv4p59sRxrv5rxNFP3DnGWz1bFc5wn
9aoMmz1Avi8UeZkBD6owua7YpASYThOvuVEN3iPt3xIgRxTVG99tIuFbB45phVQo
pv9TF5Lq179zV7wZy6mhbRHQIU8N1aY8tlCUfyYw7zIcb+/MI7l9w3tCw/DO9sEq
o4OVFisVLMbgVeHZUIprG5D/DWKLS1SmxVfpl6iXBdRb4xKAiLCIb+PoWC2+hL7N
r82XWDW0AeQNAAQZqaR02gsYXY9VMlO5DonQxoYFNkhzkR6wQV6XT1X3dgmathEk
1yzgN66LYmGYUiXfm+eodxiXzNvpJjwNeajEKLqdYQqud6HchPzIgvMSqCbV5s61
zgBUYnqjsrVwr7GrD/lpBXR0DfKspFPz6d8vlWnksGErH7joeljO0Gi0KqRbfDVp
FX0B58Iv7Hk+UjJkHw3cOGRbsfJ1fLenW3LqDrlJna55G+0tJm84BQ1DwMcfi0j+
sRuj2kCOo/xK1h/dGJhFQ3HyQzXu1MPsWXIhaCfWWDx6ZFfStO6ffcPNKaHK+XRf
EjUOJFrtknBjsd6ww61BwKckRVdKSRS26xHr/NwesVnE5wNdMT8sLGcxPpF6EJS3
97DRWqyyB9bmHW+U/is3GcmT9Yda9wwN117u7DHp73Zf08Vswom7VxDrGehVkRy/
r7f7keqF8RH9sxxc3UDU7WST8IhKWwyhWo9F3WEXCdOfT3ohXopN8MHDq0f0u0Zv
Jk/X3zD6IionwljWpFwEcWzCTxL5Lmf7NuhUB7KMLq6SvgILVa769DVXHm+NkOUC
UtsNIyooHUiZSERT1OMX78fuMeEMxtQAzn8iaxFD+TyAH1xZ300X8xuUBbRZngQ/
kw7ZW9pf9fPGvGjdCr8TYurBbdB20f++Kl+s93MVkLe82BCXHTZd5tfx0W3mU6xY
NLbuEWj0IdjSiJVTK9sU+w6AzcLc9kPDorC+RjNY0JfDbyZcTEl5Z7I8+bedBezT
Ep6IqGVNMSAqeK8U6FDFrPb/QDQ27HCepeCYR3eeZtP9IEISU1SaVNdT0c0RlyRO
vQI4sJXnZSmtu1JRpEepQRblHWTo077f1EKO9fLFCDgqS6sIA486zPQeCu660fsX
8Zl6xUcLUQdS8elPWUgOto/1TYpg7Gr+ikiLrTzQzdFfNmrSbjdr+yOaSCej5J01
nzDcRj4jq+AM58uXcVzdkCk0lM3qLWjboT5xmfL6c/1CbFI6pqAtAlp5D3uNqlg/
gYxGz+7tmJp3sl4snJKaSG298DGdzXCOJGoOLjvG9CxrN973KgZmniXS8sKn920e
K0uqgZUWLNmMq8O9UGWBVaS5Ab+xlTdnhxovb0shJ5X4cjPCYumxESTsX2rRREly
fFq0Dp5YRCMyd8xOpenID+3yqo/Bv2f+i3KtarbKxQXVOyVEa7bCHxQUW60Uu7vP
HUb3Mp2jLcbo5Y6/QzQSicmIRmuswJaUuK2TEZgGatAz53cOt9Xd3QJJHTJs/+5M
dQqYnVW7zvqsrdOxGaeccnF2uWii7JWNBb4NjIOeo74WSVlJypL2Ez8Fl6lt66E0
gq6fsJJnLy2QJk/EWJLLRX3NAehWdgYS8zruGacy/KNoF5QthqxJ+glIs4hO6cSW
sNYlax1kMc7gSslaAeLzOyGBwu0zkbRqm0EGytkv3ewQfd/oBtVFWbdno80YV151
aw4F56XkbUEV1t2vXsFfYVCXdofJTKzCCAQJ4lx/xHQ5GSJv0SEYcrMiTOrZo+X5
50T+K1V3AVE+hGdyWxqJYKSf0/zh28sAJ90qkpfN0drxjr9PuHDe7HRyu5Ktp+bO
EtYcs9h4remZHpWP/JBWZKja+5hgEDXg6jfHcOulUazxUimuAOCLi0cTYy2uY5WP
VKuattpPihOKpqCn/Z1RZDmUV9GUEwRc3a87znelsEZG1zsJQJpK+mC/Yypmh2GD
Li2sLLQ8J9z9zyWJ8yqhgdxlw49ay39fGcKZXgAioDN881zhO8SfbbKQ+xYQl2H3
KWdIoXyv2YACyApBR/5HPbnelwxuAkgDIAW0gdQli8jLZyheVM/rcQ9nycA1YG7i
wFwhggmCl7kwWulUFmcWPFOqrfmycjs+ihlNZkvkAxAJLbQcbBCwDvowVg1o7b4H
Ad4/bacwrFdMoxyX2bxGvD2YSzcipfOYoPi43AZmJEPFVKFo2hF+TlXyvazbVDwc
pNSpwHEz6npHUYGqADB9qw3NAvzf7YduyEbUvOqiIdjLju1xhstsdXxCVz9hIZev
HANBeiCYTjHRRsvTTmCiF/VHlJbFPDOSxHeubvbnADPBQ/368ERTWQZetaUMyqIk
MvL/PqlemYq3zLz+iaTNRYzE/x0QyZQ89iJHvTWgcSiGro+5+90Co1pj52sI34ca
4/ZMC0gkX4Exqf2cSpZdLXS1FBpb/3vJR6baLD1FY7V15qYNi8z+4joKm80M/5Le
Ig0NwgG3Ve1vWm8vzcRW2DbYXDrD6UN+PUINnIGyT/2kpZ0vdF2pVcbgucCXko3h
C/QQ2t7Cre1qKji9CSKoEiM1UtLkgzv5stUlKxzQ+nlFb06nwBZFMGrUotTiO7xD
N1pg8ZUZWPJeiniOZVJu4Vm3LrmvHS69teOeoxevNQKIf4FAgQwILWFpWWA/FIT1
uJkvTStUDmCBb8a59OA3ZjV/Kpq7xGgn9NN+sKkaa3joMKV48dfdKrgKqygNSf3Q
J3vtMB2yNg+X3q7VqAt40CkmZLtpCFhV8gRa+++eGzbK09A2FokTD8PKpx+rADlf
BwmcbRFPIun2uLYt+EVgfN2oQGaymrqfjP9mLOJtJFt2xjFn2odGSBvFSTrR0q70
e/B704TP3P+NhTy/TZ8Hyz4kcxxGqEpTcgL9VF8+Br67qG3fvtlSoUvMiaDkTK7r
ISgKXUG7a/96qLEfHMy/p3MwQqBwS8TKWJWi+281YlSu2isheEh9vuKqzTL022/o
OBdaNUL4XhUBbVWR1VsvXNQG3xrXkdHwZgEQ7wbjNBsBm2+hg7nPQJHOzzvbYZMW
DcrI2oYUvevzHmTL++vyX7ENAcEQs4V1ZfSsGZxPkF1KCCQL0YCwZAjimg3+VzZc
me4fLtq4M/B4a5LduYdNgmt5YbWcBhy24k4nas0zSVuOEcyUxSKwO6CmP15cQCO5
ooe+RqOIyo9ZojKSOLUIYm9wWx+PSQR7WTYGbhdCxAKNsP5Y2CpcNqACHJr2L57C
QfntKo80mK2LkrMZe9PqHxM4KNt8A6rJDe5zoMkIvEor3Ka5AbfVxS2Wt4FyUFXL
gFExkTYyQQew+Ar+i9kfHUDulEIdJACdojbfxkOfgQlgGOCRUNA/vpcAVkGWW0Ir
8vGQCbFjL8CsSGeiZwiUtPjMYNa/V0t5Fc0SMUTufecKkQ4ctLkz3mBsWPPOpEFb
Vz75W/3x8aosffpSmMROAIwjV1WlN3FFFglNd/sCOdBVkWDL+AGSo95Cv9uZXxNR
8IZpGXM8hTQt5lEUmBp+otx7szitxgR3XzwhAZukKbfE4uNa4yL8Ds/Gqy21/nQ1
w9wacGTGOoyoaQhBHO9QHkQlpjMiamlHg7OfGKKJ6b6R7INnZjYSN8ykL26KVG8F
oEiP9xb0s5XgrolvaCdcXJkhyJkgDtfJkE1eRiDHexdEoQLw1jfK5E98UG8X7R+9
dei5BqKBrKOteRGc7xE2AwcGDXyH975AvOr528Sr4TG1NZn+8qywjKW6saTwlK97
vRUSe2WNCk44At+rOGHrT1jCL5YsSCp9pymzc01fBo+1+sczvs4ouyhpTwtBE5F+
rV3OldYSZ93UAFCiLMlqNZe8NLvRZofcS0LLsYY2ug9OT7N5GN8syNkD3rlJbxL7
apponQ4Dip7DHGKCqmVjiDAK/Mz+RoHOKYA78sZx2sbvltrfKI8U9iWo4PztGc8m
mhCQiPCRM0cgSMt2XYBkskyVjGG39EjUMEO/YozByZSbiZ5LeEdKaZTm/1pI/C1a
fDCouYhrsbrtGNJ0m4hEOT2KHSm5gvgyjnCbmlnze5xGbXPzyFA2PNQl1YYkauPd
vydTfCIuSFdHDrrkpWxGqHqeH0Y9D1ECwn6HOJ+Qhpu0O5XquRvvbJMch+FUBeYq
8bOC+ruJ/qCjMWselSNntKBzNWv/gmqcGhwdc4M23984Zw4yrwRKgn3Ih8M4Tqx4
dBDIPg615nHkzVVih/km5F/wiv2rA86z2BKi7IgvPj8OpsFXx2F6kDvxm3n9TJKL
8KTQyq9iPNFkYceMQX1/AJOyWFl3vLa6d4R6DPFF7oTgWPSjg3UhO1WmG5VLY/sV
k5PwmdjzgIeJulkT91/B3rwd+QKZ81GVb+H6zCWtZa4DnfiAllSh5/NrL3fqBIr0
wkuUPqkJEGTjv4RRcjv8wzBAylFEtInvsKdYPSOOCBmOrjn9KQlwZ8bBTiF58783
QkOR7y+TZZxbOWLxq9cTs5LSU18l71VeIXB+YM+zQz91XeKqfUunCmG+lbNuM8Xe
NwifezAc6eBplzmDzuUA8CfCOakmKbsoaaleISJcccfimhVXgce5b5Zi0kWKEE2Y
QBShgyf5e7lx8MtgXAf/JnZ9Tp8tIFXwi7vVa3Ca15pjA9C4xQt6dBm7xjQq7AQ7
9P/+ujUw2YgW0F8VMuHdcMwpsrUYO8+4UPQ96uxWDvDbZrZmHblO/1jZ4RcduK5I
aem/RlITdt6bX6QptzY+1Cy5C04klO8In64cNIUkQcPLkRGUlGfpHmKTCNfaFG/R
K16W/yTxUipcjP7xu6Lp9zJowMR+DyKoOS6gX9JLjNlRPOArd0XzlwPxMvLHkIWn
hr6MWw2+x5rhWJj43Xx4RF+qApze3OUhji+c29r5hktupj4d/29Srf2tcLs+8vJF
0EO38FRFCL5MIBK0Fpguh/Dcv3V4NXpgijfiCrwit/H2wa/cHlR/1vehVEH/efuo
CP2vYW+bYOUq7cCrqSkB4EDTXtt/rTkI1CIRlcsHKDBO/EbV+lbqEZSExurXCWkX
HeBnXeVjJiS3QC7KIVHSwzUxWXbMmmRdd3P7yyWTS1CP6nsYOes7YKaWqZ9bGl8J
FLXXVV99bKPq3ltesVYGDRDrXkifau1Jo1xeZiQUaUcA995VT8BP3brYEj2/cQki
fvc9TIQgHLfuB2p8pKFzsHOLkJ6aZqFvAn2VEyTy4MYKSl80QPByN2RSnm0aqrmn
CyqJKbW77y+g9qK+akXhISwg2g6oZbODtk9IKsFlu4NuuyDOkaoH88QLYZXyJQxG
2V+E5sVTWA+5QOLcP5P206tZ7TltjTqsqV2FyN/xaNwZ4lC1aWihhO2eOm5NhZ/A
dimwlmkdvh5pjdO640YTNEN6Z41AiwnKPz7zPrWqiga2Gto3rrYnG17hib898eto
d6xRalDJlxmvYOiLmyXKzkk5x5cy+Vb0Lo/ZTFKeokxZtOiChwJ7BYDV+8LepQAS
1vTsMbsGVs1OORJDuciLOGvVl4+BRBC5ISR+gffhiCT4ppZdxjTgGdpi8fYl1H8n
uBNllDSBUypmGST7RNoxCmoCj/himnc/b4dxSkl8sNf3kwxwM+Rx2xMrUmtuEJro
0Xp2zI5I+gPmrfA/kNIVIq5vkZcDL++mySW0tFBgTeVjTTbjth2WDzjVYqyUsCSf
fjOmCO7qQvXvSMc3kiD9vMm/y9IqcxIo+EE1JnQQvHJgCLHAt6bxXBna3t3o4XVI
Mwh25p9tj1rf4+R5U8bAFauW/SwXpYsyEgq3cqxNcmd0j6dNl2meksEYzpf4CzS2
V9MX8GdXd7l5KLipE5v/TcxY5TBlMIizaG48qR6jN9cTOs1WFWtCMxO+rWGxQ5py
o8c0cDOL36kJdreaz+kNzB6vzMU3nfGxm3ZFD1vYhvUcT/Q6qzGZRv6vElz/616H
+jToG883Bw/fZYf9ACtDpf27qnVzGs69wB+T8hcqGTISq+jtR1Mz9Nf3S9BKCYbX
Io/NRzSPD3uxHVNkh7eov3wgIN34ZBXxzyi3K4+cCIf6qIvSGQ2U5LQqxgAmsiHk
ihPlnA52L2oMN39PF9E0WWkoEnUq2ElEx2SyjVyRpa8XZFfP61t5bj5qIPpIWaFR
wH3oYQlH7hjk9sHMnlTMg+KvpWhTjOq196/XDD2cEyvWBtN1Ls69Ldo6LD0eZzWN
ZxyoRgoIYp2GA8FFPe99697gDDNx41O5A2fMIvQ66wJG6HwiXnUC12IJFpFnSr5H
Nl9HJm5q8nvgx2zU6pIVUM0NOiW/+cZdrVy9OYSTJI8ClVL7e4HDL+AYTjUWLtb/
7+Uq39CG7CcTjl81ZdTlkxpZJAOPQLIAaq2OQde92Iv04l9EXr9c/jm9tfQmp4si
dZBiK7lWxZ2p/xyj0/hGSfyHVHGwkaSCOwYZmc8cFyl0+bkec3LQWKXigPKaKbON
MMlH8VKCQnBUO2YraszotO8BQsmO5Zr0NxKvIFOvqZomIbe7sAXIIAqim60X5B1W
jRGUJPC9mtutvjo0RdzxQczbHmkzlTzI6DL1g4Bkr56lgqfPS88VtwXIYc3qjqpF
F/4kqIXuyLrdxqO/Nlx8d51D1wHLwqGZaOqx+H5FAi2l/mqAbKTq4M+xTYOhc/Ym
cF4BRNmVbymrFYJ1SuSSp6yfBzCIQXR+ddCrdWqE7ks05wOHN9auk1YesUN2P8OS
LGnSiOvy9Vv4getMZwNHecxxVmtblBU16qLilSGRY2zWrjnmYvU/FXsVsK8CSEBp
9OzdniZiWgwazKJH+Qmf7cHMiphDEeurNKPH3W8NxzZPjgl0xZy9QIZYLPCzQrk9
Nzjla5QjezGDHojDJmAuI1kuM91Bl/+EOFTJK3B8pLxMcwZLHSf8fJp3B1F72ItG
b9+kFONj9V2hFBudhCcU3EHfPfxltKvMYpUtgmebbzCf7gp+A0uD6YNKoZbZPwR6
c6m6q1dNYKtYMe5hEk5Y0blm/nac2j3G4OCyNAltljMnOE1//rToLsv/Qpfm5ZFr
jKij8lU5wCIM3Z1RCH9M4H66L2+nA8+qwjyHML0lyGY9h/qRJjBozbl6nZe8rBwM
FNF3IWpX7mRz+CiORPoZWgGzL3vPNt1Jfv+m1Hl/La+9HUJ0PRLJPCb0y4IQ6H4S
D2W/QaBggJsqlad5YjE0Nxu6qg6KcPi+vO7F01gxj657ogEPmnnBBf4PPRuUaZmG
YwtM7L8dDhXK1BuV158bC6vNW7ZEm3ibWuTKHUBc/cMXc5TEEsSUL5TI5zrrRxbM
CtpUY+TE8pZr8HtD4gaCB0iH4nQI04iaR1Xioz/GmbSLeeRob7wSLvFeADLlqx/2
9kJr1/HPkP4epV5ARRccgM8NL0CajB8iVlMeTfo23X3+2G0wZfINcwGM59oHZLXU
CJDdroQUHOZKWJpOi4i1YLN4Yr6iBa22SRwKag4atM7DKpv7BgIE2Mjoy3GogvHg
nQ8b9+ImcfcTEY9gE/k6hMm5t7HFYiscg154WDw7mE0H9Aur6IxPPajV3kzbibms
AucyEHkYnSZQYWExl3r2qrbLl9AW/rkHP5rMswBDCibvspZ9IqeMHdFaK7rDiAoh
7PUkddY9dA9cnCSGlYlaBBaAR4benSkBa+H91f/mWltUOfrNEvkrR+hsvUMJxklp
zZ86EYWNIMLdOfioA2LOk6OG4tO//nn6RJS1z/zA9IhH4blCJ7D74N9arjANllIT
InimN0QDNHyTwC+IEOpcGxkWTFCUFstYIJ3iXz6mkvvuKU21O+WHWqOdJ0O1kgZE
LeFdw4JnEFb05ldOT7f1W8CNw7o+4K035xM82ASFJ6a5WGo95490b9FxLp7B1kQn
Sg/XrIKglJPF7hDGWIQD5qJqiiyo2jM+Pm7CvWrAGwNNNcuwg0J6HtS+0FUOpJBE
9t/wMr3HDfBgSQQkFb01ogqjltV/kT/GY6cxe0uOgmQAlmJGaZ24k4T0HWr2n5wa
N5U+HotlYK2Qnbbd+f1wZi0JZAjAAZmTQxx8YK5vos8Tph97rgxB+e1JB/BiiuTp
9cO1SYy5YzacncRYTN5le/hWT4359eyUOLG1XJ0BqOePCsy88AkZXPcDtaEkpdHF
HNoOxleWa/tAwz8+mXPWye1+WGcWbrZwNIvowzJ4gDwcXjZcqPL9cr9CtkXA9U6H
3wDSQVoxie3Qy5N2401kFErtJRzDhO1G+xn9W+Y/T7u7dhb2OqXhLnYKLklH/1di
O8UkbYF2fXMTLxBPBaRiEnBuMQmhl7qyGyz7KuGWlsVm1aGe/U+tavI5B+oneXkz
a/Pts7RH2e4Ua5IZrTDDtPETOxLA72Nlmy9csCX5F0Rv7e2kcLWt0+rPjmlpb/TY
jNhqZPGajjXtVZjIO+7Nrq8iwPSHnZ8nhUuDvJYJt1J3clPea7Yzp/+AseUMY/rq
Nz4+QsQ5lRHj51Xl9n5wU4jRUaJeIUuT9Ia+r9h4DiZhMX9AgtK0SCiFywjeKbWQ
swY00u3WDVI53LGs3UVeQBBMZU7ayzYcR/WWM6g/GmBxGMoiGgjZDRejMfez3jt5
ezPUb2FpKtAbI55o8Cl54RioWE5CPAuR1aPTsdsP/LMIdkcvHs0LFArArOyOVR4E
cAloy2mJY/aNiL1xtO4qsXnVlCWqM+SP6mlrB3EjLRy3BCvdY/RpqixH3MSAyXDm
TZkIp7pA+InCloeScLOJLLQCYWKDwg0nDf2NCPYXILYMhbrrd03nAKbxg8vitT0B
aAfFVs78ntXrCcrKdQ5tp6Jeaj99BF6bVWJQg7W6YaTIQSHvx30lfauRH9YjJ6Ph
hXHGA8yfRq9Hpl6duFVgccvle4dV6mGMekgmTVWsKvqiNN0m5FVM67zSoP6CEgL4
GisbS6VxoDziMMf2wksMAYNj+m4kI4CdURIfzc5s58o3qS2shsf6ufNDesfnVnup
NDYFpiw31GBBEzcZNnG/+IjZkzp6Kcsm5n2QVKmcIMNX6qTMxK8AgMEMfWLXBAFk
ywTREBZ6BQbnAuco1s6JVkgvTKjmqsJOhc1dn2g8O35sd7kJcw1gnyYKmlNleTKk
JEyHWka97IY1tG2V2atzBKd3MyYF2VC4cgFtdbyntt5vzyXI4LTeHJanfkRh7LEw
egCthe2JzokswatlPzPhxU/FtK/Dy7yxtG8vs/elRfnmRlmX/z0HTJZxvYP8k/SP
DBpCa1tcSG9Tpdxv1a1Bi3nDwKtw1i7BTiwg7WYz+x8Yeex1ldyWdLBYWlUT7xzc
eXKv5InMJhF5wSM6h/CgRFRSE2XwFlg+cshgqRlGJi/mG6YkyrN3V1fXMxA8yPJC
oD7LxqyNPDnD9T2FHzOnjm6WhASxl2+J5XbTnKEmHyI4aaYXmgRbLR6LxvfinDIY
Fs8mfH7uxFFv3NRIeajn61n7TbFjQrkAICX9BeUJkIwvJhwnG3E/IdiygjZPk8aa
qS8AqiiN+bttQWX1OIn1b5gKUiFQ1e+QT01EoHB4BBPLEe5f1CR9MlRymEGA4X9f
eK+2KJ1OqAQthC+yONkkgBSuNxHxXmj3zYGxYJn+a2Lr8ldYo0xSVdFt2PyfcsXt
Z6GfMRBrOurfG5WQ61IXsxvJiEGdYkHSEt0Zc09hnDEZgi0QiXnzUXY8zVa8ZLby
0WR80AXXIpBe8M8OHxpsJoxMQ93JmHkrkuR3JCoGzUpWRLozcOtTPP0QReX8NpPi
+R56lg0fBPF/HmJb0YXY2IhR32B+0xPiDq4Jj9Fpt7Uabcbv25dIxjI/l4WuCdGA
zP4QheR8nPstVBA/mG+IqEpcXcb6BfXOuqXHY0L7+ZJGl3HgC3sBaPTyMOML9ubU
9o5ZCnrU2uzlrXam6tvwQYdnW0eOpZNm+L2JIoN6RzDUgBvidzxTmerAVNKyUqS1
jcB9jL0MksC98HWO0P3GrPyaYfBpuf3LqAirxTfqym9pgJijWVeybEnE+uaDVz27
FwkfjDk6NX3IphMLpQe8rwBGTp0r3R0XwKkbqVp6Lbx73LGNvw4TQ6q0gpteclRr
0UMBtOdeafkTd1LgHoX0Q38yOLEq9KTljGjuXTeVTUrnhbmrOpdv9E6X8PwqGJ9o
2K+LeklD4KQV9jYqfksLdQI1BuEiAC09OCiNHoCYTV/fMYLtYw+rJVXhgF1vwbjC
ziWWx5c+/zXNf0A4CIpo/w6IWUbuP71qgh8DfSkU4UFklXIeLg398WhsfrtYkBd/
YvJLsHjEQnvWht9EF5+w3wnz0qZrTFa4/VzNWZxHWepxohIDoqYh0cdKSnT/r6HR
heIKTd30f11iy5I61m0as2BjV5pEwqomecBKsYchxSZWk+o5ZpZCUguErnZi7JOe
ZgWqk1PEAkHijnQ0QtmmqhwTFcLdB87/795CBA+9ib8HgaR4CVThxieP9jPW15a5
dZmWd6pRh2tqZUnyN5tAVNf09Ttql0MkV9jemmLEpjo3PqU+9IRfOTaMPJxMDRl6
l1b5LqwU7HF7yOTvNw31sLGCUsDJONuIH3/F1XGsrUWEwhZSX2F7XoMEpi8uoXix
+Mij2UBlAcTCj0WUw0PvdOGDq6x8bPmSpZ3LkzooSVw3+dvllRluEuNHkdPXkmBR
Zqh1rpT16tyvyhig8OnL6Yfsow60BxrHjzKL9DyXOEDwZ6ig+tlJtMh+FbP3IBgF
UkJHBEMhNcRBIVudCsjIo4h1WkFaecAiQ+ezwrOLSpEn+f3IPTiJhRwd+R/PWED2
z8thSBk+v7T6A6mjZX506NUsN55/hQokd4eQNrzLOdN2mAuzuwnQE41VHmGhWjit
LkSL2WhomBSSr087+3fWb5KpiLIBWc2U7WW08XH2qC4jABMb4oBXVQBlSoMUZamn
d0MSzaRYekyKxVUTK3GTJQwphhDnM9X/hDmRxAWREjp9GjnbC5bKgr2FL8LeZfo9
k/r9/ZnzXY01Wu0QjVQ3CJPrwHoW/CwSBNPSSvh5/Zod8bnRidkD0neYsPWz/dzQ
TrsRnT3AVDPreFvFINHcvOLUvt7FoqakkUGlw2GR7v8K9WiMC5RH9S/E192bWvv2
/p3VGnPEguGCviEUJI5dTGtPPGcVzkaEWDWblO0/E0dW30gU1XtaAG2k+23ohLG2
QbbWbS1grjXY9cPAJgNe22Oadie2ja5JYFa99o64Bn4upPW6MFtEVGfzfgf9odNy
B8Qh0DBK4PZXZySIM8OI9Oc5yjVJOWl4MBicjpIIgCsXX3ikHTDIpfVvF07Zn9v4
EWUYtwQJP7X0Wk+rGtQMjQysErx8/Mdt9GeU18FXU8HUtLpEgKNBeOOUOLPzS6Wf
um9YMq4HEuy8J5AuKx5DVlbTRmxE5/J/A5DDIeCpryT7Z105xRvJNOJ12SStgmf0
SHsDQtyzVVu6h8Y/o6nTGpG1cyr9twDhbAXpanDx5aUFwNLGpeebxaAyQSQD2OS4
avNNat4s57aR2nFYVkilCvWgu+8x2wCcP8LnAOsA9JChSTkHKnVB6iQulDcVUXl/
LZve+VbUlcbgeL7PHtCIwyOT4+eDjo1dcXnI1MHYbZkZ5Fpb+IdSo0ui8XPBY24/
it4nhN9SBE743jiV4sVuG2yhfQuJUajZW0Ip/QAW31nQ8fHa7MwCOYto50gbMjpm
ps+XBSKbXMCEeQtJC7LCQR2NRVecEf/HLd9wke5wbn8KRtos+q1jkmjPxHRuD03o
xlzX8MdsRcqswjIf1iyFUpn/es7RSwzUH4dpcpa69fycXsJ2qFqGn6LzZmrPM5nd
G2P2eLS+r9q2oxyR8L3FrGE4du8ja/rJf+xl127Jj7FWGZapJ0su1dsQQMi4wbAH
nlJJwgHVQVxWPryTvw4oiPEu8QRk4cgIOLwIyKSfq7YfPcIV5CY76gWmGSqZt0a1
eRCqe6cPzCsOsguTzS/OKangctRXrtqWTIBw+l+qcZTsqkjMskKz6Ennwj2VqKsT
ugjU04a+x2ZfceLpPHASQwYj6dBF1uWTV8dJnksHBCA5jba6Fby7PpCN2X3OJEcu
CcMOTbqWOf5eIjuvgQLv2EY937UURAVeHKri4XVi5LL5biHoPlwJ9LnV5Unu3sn0
/2urJ2/OvPoa1T3EOefcBfZeIhuZakDS6rRfm62bC022udNaGs+SDU7aEQftGoe+
08G7RE/oxlTn/3o1VUay9rkI6l3bhuJEyfs+kD8RX7dLEET9hxsC3goPUma2WAPU
aUox8VL6vowQrPs4TXxRW5IZZtxD/HZSHp23WanWO7/5LVYtvuDpx95y0W10mh3t
sqYCiQjsxHV6hBHYEjlIXi582Y2QUnyF/53dVEql8CYRO4CsGBa0P8MhEy3qqoXQ
AYOmjm/nLhlJ7kZjQiP1wdF7bnZdHw3DLEBglzie7VC1O0TqVWYdjUA7Ouhjl5SJ
D3ORwXgbuDElW0oyz/naWe4rgwgbsZ+lK7PUGko4crqvSEQnmhKZOxMLZEDPegtR
YyNZurkBnWbcfyLfH85+Noiuip1GLQuBhg7EOMU9g0wb8JZx1i0JQYKpZLgNr7Q2
kGmaumCR6YjoqTbBosQA5jGCZTXWjQ/P6NVxbRWEkz8CIQ3eBsq0GbhsFQO0cCjZ
PYuWmalr3rphNt4fDeXL2nHXSgkyhSWBUx2RCkMl97ymNn2lHtR9TYj6KwEl9d1c
KY2aXFi3z8wy9ziS2oyY1yYc0otvjoWmEid7Zy/0DB8wAYQkVMZKXsalBzqfapRq
fSxZu9e7fJzaPzMxOVuL7oTNyay4SkhjL1w/Bmww89RKLk1JQv5dS7iGwenqWFcC
oB18pKoLVaYEJI54b3+VtgxD3rREGd/dTmzxR/1qQfHC7GY+7WE0aDlIzIyVRiPE
9eQ+GYYvKSXcTIdbcIUuhLgMVD5GHmYqEVWCnKbO9kppCQEmh5WZPZP/rnzUbwoy
yG7pU4ic117s9F11tcVvj/lzlmsMpF2Nu+bLCZL4fbMTrsEziX6B9cvVaocFAta/
/zb60GK3fG65Cz/sSlIV3GogR/ouUZbpMgW14LCOcKzqsc0juWiz+yAWUkWlWxOs
E0orZftsZAM1ovge3CKtTepX2xr1aRmSkniMqW+yVpuJmJFCkiPt7yo6jh++nOU0
KjOmmRkE7ajuAewGE8B0zFfV/4bZN/yVsc6VMU1tW9yNzhWwEPCvGyrzMzo1kEUf
MkHaJ9qGJYiFJzd+E85WPyE+Fd0Grey3lRYEkbw3jBUJakm+NPN1/c4OjAwU2QqE
pJIO7UsO16Wnjg5DcKKNGt/OZg4h1xjRnHuS0J/lUv+aALjojRnSud8z2OLKJN6q
2klleqjcaiLGHhtfkhfwp6mqdBN9qmoB0JdJqisqs+QQokLFqdqtfuAoVjritWzW
PJwgDP/C5564uY/pSBQSCUBPd8SOokAQsVaGWlyL/XaXQI/Ddb4b4bz1BQ4Q/wMj
QwcJReDBQr+j04xxxBks8zwWh/kcuBvDegF9g5PGjRSHJBylNmkT2Sgz5JptqoSU
dvuwFHY7pIVEz4f6ZvRGCjC3PAYnxwhfNxEHj8GnzmyQokDJMIu7Ftnxpf9GRw5l
155iVTOzHzGEkrk8X2uX8wWO634PbrjmwYKOG4WSeKQ38Fll4p1m1z0KFMaavIzj
Wr9juHa6YJU3qItZtJzMo1bbSpbx0dqAWTMNi8oAxTjJ4ouol47MBCylMPZ1tKDf
+MCq7RqjMWCX/KgTHJID2UfJrJ3ezz0mV7h1zcoYL9X52NeLSy2TopMETyIF8Grl
ID1sLadq293GBvFTNjrjgklizLncyVgJzaxoShYyllZnkDJvfhxV0Xf+ziuCmS4V
sjmsmPL5rUom8IWLv/vtuSCTZ5ERpG+Y0uBtkeZNJca4d7J7v5Y+iSVdXeZZoHu6
dswk/qUdkC+zfMRPcmg6tUdxiEN7oG9wPVHM/idOcjVABa5/Ojnc/yF9ML2oqPTR
BdPzlsPUjJUGr/HqRo12w8ijSZtkmhqbFyLjd9RvJNQ+sost4av5yFqkz2QKI9TA
8kry6q9p0C2LymRBTIUmu0j1QF/rPeRQBZo2eTW/B5ofWQ1J+99s9bwZ9AVmc70p
UpEQNxhGD9dFUGfjOkrpletie+kb95Ymu9XvY6JGB2vVuxC2hqQQ05BiR9WOnprk
dVOVFX6WwVHxOlKcB6Ya9WoWtMVBcvTOwAp21jWHgCqN/efRhJ1luw5TEOiLGDK/
aeyzGwaNdYn4A8WTDbMb/bq41dJAqHvK3EKgiulwPaH4swbOCPbMyoPeI6CVFvHV
7EZtejf/jS1djku2DJHPpxPubfMXawYanVaDZeCVgOAZBnAsioemLdoQbQYDNwag
X6XbxF27Odnp8ElyehQdgbIF9atNvTnL2DNk6DwwQoof8jFv1ymfCZo7jevL3+/j
6gE9kyMBQ4WwlMFiq9oE/s00IFcPgQLhBvgYpBK7SEZPamJFqAXbB90qCetLVHuI
6vA45LEEhUjQdBBNcIpSOd/4nssfqhV7iT7GruoHNMewU6hwVFNHScWw2+vrtevp
WpjRIIn92pqCW3UnoTVH0/L/d6yyN3oPnL0KFz86Sqn7uCEUuUjaCnxvbi2ghU/f
Qa42lSfQRcICUsY16p6kPo/AYiSHbYQLm/K5ZOHXioAc97CPR16M5UchCWNPk2QE
mZ0z+1GvBbmOajNb10idJvIwDNruaNnUNwFy5OCNwG42qmNpV/sDjRipAIezISmG
jwZgAoM13LUABJW309FA1W3GthFwu1AaypS3lHsd4tuCiyfm9Yu7lCbsyhynIZgZ
7RHbQTca45d8P094OPzUVZpG5MygTJZUsiG3pjJOZN4DQ8b6ywO5HitOdKL73m3Z
/ngsdlv9IvXc2OhrEU7rRn5BSlA+m+rmLwrdGFwDZ+4zRLox8lx9MlSj6apF0tjs
ONv41cogKd0RqJJtjn8Yog9FO3a5D8NBO2XKQs0bmS7UbX3KbQjvRGK4HlF1Nri9
lb6Uf7W1TBWkrIcF8Bx3pMMumCZ+XP2CD5o0EIwbEhj0809C9sOQtMYSFrhoFSJg
/sa2qw77r8KG4Fs6UxE9p5OClUT6QwYUaAgi2O8rAwz+TjWnyZ7NseZHfXWrnWC7
SxXgbSgESMSydZFl9QoYbQnDM6YDctBGQ4fxHg0kseM4upByWsdD3pfsfuiBHUZO
0UqOUqB9khNbsdipjqFfXluIg90I+fKsqu6KwFZSQzJl3S+u4HQtI7+YN5modwxI
yaQIwNn7npUk1qp2WGCDM6pzk+jdJRrDEcTrsjyzuCTk9N78Tx8xpAirZa8/FLzn
3eJIAOPfDqJSor3g8aGJ5qroVYnndL8gwhiZppSr/YVSjEs4r2eqt2FTCMKd39Eb
rQzgwcpmGesdaCXTlCDCtGyXLmpuwoftExdzE4eWzs7D6LuuqczNtXZHC3LS2Yqo
4ZMBUx40tV9R9IZoiIV54YmZliZY8TZWqLsQUz2O/iCZIIVthKTxglkq/wofhTd5
W+7te32qi9lgDk6HOX/2BAN2b5pKgbUAsAzQWF+ZeZTvL+Xqkl79LC3Kz90cm3+s
paGpVlcCYhJIATeqr8u4a6qPqDK2xvUyRIsLg4KOPEXFXOeFLx01bDl3E8yztvzu
JRXVjKKLdVGkhSVyh2QpPKCIk9XiQvMVHi1d6EkWraPSa8rQeCOoXSpHdBrJ3MB0
5EklRedfFSEVV+7xGR73Z2sV91gV4zFRcbQ7cFK7BxYYtO2ZLKwdcy7s/JlXwoCG
hrcbiGW9x1fNHN9I0j80DyGpmFfnVuqzF+Rb2BmpjcfsRKL22IXUbPdV8/8BQASg
2WzimdXevYxmj/xBrQaWGmxEU+J4Wyb1eLXnUTu5F3AHrRYN+KxHvd5wCSwgItwa
3dJ7dg0brgnlGHp+8Vb5DuYAMUTeOBWHJe/zX56pEICXRWDCllD+c0ThaYb9lgGx
lOhpOaNYNl0SeGz5TTObOeSn7yASr81VtzoV20gFwjCKgA7XDcQwBqcd2u4LROQ+
VffkuS57DoWHpW+BHeh/hkWW4/JyBEMm38H8XGJCX+AXyFaRxtY6F2Ktv47n+Vr+
zdjrtmJ+Y10P4fqJjjr6rf6YJvPgIxNYjfqhqzBpKCDf/e0DpBIbiPHFEZLzYn6z
S2GXIxtOVb+BJOj+EaJUiNnPgE5Q1plqGPFLr5G65ja+yWNRVt4obUiEwR699++V
mUczl5HBHio5xmwj6CeXc0At8Py5ZWI7VNL9HQQxcc59W7X+is/Hhg0lckh29Q4P
/L2UMJgSTdK/IUoSUsFZ0ibWEcZjkmYp57GvKU+Dzhaw+t3zBFolfmBARvW7M4zf
iNlxgeq2RQVErYgcwKBTAFj9/kjcZrWGYSDjNub0j2pHGhpKVa2WjGT56LNW2RXB
AIBvQQUINxw9yzGC3yoo4rn51OtIhs647Gz7HqMUt8QsisafEx2nVv1U0FQTkOV8
xDb0NXJrYBVykOohBnjbPTvWO5q/5z9hMK/EbmQw7eYDi97ESPnq1NDXBVUVSX0k
KLPQOgqtAdZ+BElx8KmH7BIadRL3MdDyotOtXuhyWjzDP7y3UKDW7YSFv85hrHEK
YSiDG1HLGb0EhKXslZoFLwstCMe/0YlrQ6hrBKB9nPpVYc2mEeQ+IO8l5ij5+dhK
0Jy94gZ2o7T0QK1xkXpJ2PE+zxb0D6Uj0aAW0VSbuMvt7ItYJ7/drKzk0pPC8ktU
5rCX59xtit7T6FCz+CxQaW2fY0ckXcWjHqZNLn7+3PVa8Wgi6n3nbTRMnXo4IUBs
lNfc1a0tQxKQcQ7CQzOCsufe29Gz2YGUWQDDYX/1rR5Pyun19r6tGNy2K2oxjeMt
0e71Y/qv6VosFZjQFU4f5IRgqPJWcMiKys92vby5z0UOdQffDHNOso0rqSzPnjV0
zxnPhlvE8gyST9nD1FWgZFCfJB3MAb+76olmmwNlRytCcZI9FZ7dqgheglhHbgwn
TlQ9kG7+sLCJ/tnoTE4K0ApsOJQeG9EZXCXhksrlb7VfkJ7ww3uLw7vq1SZwEKsD
4Ze9uqZ9CdNRcJ2w1pLRqaKqRBJKxAthUDtac/ZeDIjDRMC+6/Ki5i+REQrU5Jpu
y2pEA6W2RJR6ijWjsPzTSL/iir9xQsEug35kKD4TGf11p0tzW2cM8Xh0jDX3Odiv
P87E60pU+dsbenu+Ejj48rXj+PcHA7j8aSDOcWTz54LKetB3A9y1/A9NlKYlRv37
CZiVorL8PWquP508AslaD9tkvjmRTxmWDhr8xlkWjTNUiTzZ8xMcbRL712Js4jTo
4E8oSVqL/V2oen+y7Sc+N7uf40v5Icw8lXbKb5gxWX4Dj0g9dRoZADCiChzwKo7z
pRcs6LSg9n9f1GHPzgSSmXGAKw4bkuZVHy8GPKOQr0N/goVyIUKBF/RlJ0VHYn/D
0fQr9FkxSnzYTm29ygKxVed8VTVEFaLISO+Fa3ac2mUc2bx10uJS+VyBVbVXO7tI
SZYDqZei6dskrp+g2yk7+aXM76YU9Cf19ylgYZBcNqdBK0D+pyFrhiZL+YcqXfYA
TO2MMBY3H7ft4zaYwGplLaD5v4VFrdXSyxwWi1Fk/kTqLorxl5REdeSOhMuxIWJx
kO0zPd4cuKduGKJGSTJJgLj3T/EUzsEtxiUYRRxcHCMyj9vOVZRfn89IZrUhI6F0
zos9s64VJ/nf8QGXzXJ1+ZKVOCoWfJQi2M7XO/lJFStwN6rF5H0Dkqegznxz/QD+
OBSraIlQsBvJs9LmN00IJokKOxoh2+rdqocvgkxU0yvzzkWTzNPS6zMOyyiGL78w
d2brtCHADbfhwj4xUiUTvCDrh5tDZxV9UrdeFJSilWDouEycSbRUq5/73p0WpJ9c
O0txgqVjDFpZK71DxPI2Rp3saVLNGJInpH/9c3A2xkuQI6swBprbLk3tvZ5ejnOY
pBQPcuai4+Mlrut4eKobVDNSXeZOfJiwzmCT735xQOGcPJMONw8a/H4IzbWfvQSf
61V70fMlJvKd3iaEHKDxXP6m1lywEePhcro1wwrxYPI95+gpzNIZYZN2Uh/um7ly
Tqj+/GgcXDkHNVPaMEKYF6PuowtSwz14885zaK1edLjYQELHsX+7i1GjKAAGQMXb
jGZ19OTLZIFETzQiS/WCTvwQerru86Dl+Ecf7IMHLu9OMk0ymNVJbsgyPSfMmx3I
L3drMk6tKOhAOLWBrrWkGAMaRZuDCDykVE00LcYJmPnTgUnVBzkD+japWo6x+pY9
KmK1O+dcRkap7NZt7ak9gKiST4msZh8ZrNsv0IpDzyIVDZ1U4lU08hkT2MU7j+qD
oi5cozsd2JMaHXmwUnbr0KFKL2RfNI0h0CyNnQcrEyE696DZsnvl/yzW20T/M88Z
Ee8MCq+KYzXubmxmbnln6v+bfGXEEectSuIbryA8feg7v2mhJ8MuPBTJhJawEaHR
PS+qGQK2iFFoOvm6EzSdqmHlu1TTYPkJU40t1NYkGXikME3zbyILzo9epZ0Q9pYA
D2uVfi09yMkj+8aAsh+vOvhUN2rIFJDkZNbtSMiqFH3/HHIt8RdstlVG+SC7awUK
5hqcELHUl8lCS2d3k2GYHNq7qeBOuAgtLkFb9n598gVSfF/2EXFEzVlgsbVgbe84
VDdRSM191PZN6pM6KTiqGqmE9FrVLbivgQS+/6lzDkxRbWVvVOaCuPkzbumX2pur
aWYz7YBdQ9aGcWtciAVJH7FrdjvgVoFU+yNeIq1Z5g2DAZBYS0gPeigmsC9z6k20
aXEe4pDmyu+6rzc58zRuF23X/nOz2D8zCfgX2ncWxuw52KPKKscHqDFib746/lSl
qCiIY/sFFHi6kN1OYzzvCztnqVJ94hNz4HpoZn3HE3bpDcaCyixe50l2H38hKkub
HTX8TIUnyvbQd1wyaJUsByHqP7vQcJRYufZh3nit7semnuV3fFqkAQ1CoZaVxs53
RnqdgkY+yKNQ5ONPhcyp1+ab3h5PM63z9lxF2VqU0q/xA4rbLL2DTT90gmcpRTFF
6+9z4hCdpKb5qEcZmjwuNdakBei0XFS0E4PrPyB026axmEJ0ceaUAXH5O26+b+Rc
eH96Ew+RcguYULNBIuXNDuHj4HxetkgTAXGIHdsO91QuHjJtNK/HpR4eXucq2lh3
E4gTSI9zNd+DAhCUDIknC0Aa7e4X8uMTeuKCMe2VOnoUfynLY4qZZZGrx56qpoUF
iAHxssdmpOO6wy0IKiz8tO7wO7uOkBLCEWuw2CoRQoSbRQTKAhlbV3PBOlECMGCQ
ItuGXU0SLmuSFkdyQ6lCXRsefGw3A1ZCbwbfaR9TVI7fGSdnvnyINhgbkRsQpYHx
yxCfdeACHKbAlK2GHImLljNEuad3FQRBflxBaTaPM+PQKwppGKTClofDCDXhNvPi
6AZK2WhzdcBZdGYTDl6SkUUjZg9w9655veTF2qvAfpgHWelJ0OHWwT0Fnt/kUoXo
rxAJOq/04mB6FXI1S/pF4m8Pm6nmVWNekJZjSGhggc09YB+g6HOOl9gEhjE4XV7N
/4DXnu18CLjZN/PCTsq6HaQnunHzULDmErJwssjEIZn22pYU2IHQWw4FcECSjkLk
QZ8Z0cx4eSlDfe58FGcrU0BHt4+N5eG1V4pQb2PhSv7UiwseCDfSYxnlW1g9V9vP
CayJlzDEevHH7sr/wNyd5X3OR2g7sLNcYVGZr+NZpJORNWsxe0/eLKHbVGO7edIB
GfYAqZsWmFKHlHS6yBJ+6pUw6du00SMCmhwKaNlaG43rf7ZF7XX3GmcdtK9xHoQu
fMJjo5+0cmSRr+3AM1nhgkzEWbvFbc+cIbSXCaQvhqWeTyKFl5cbbVXVyrocC6ro
xkW8WHZ/hBh/wCncoyhBS6/QLfGGzleL1f2vHiZ0f5BSrowyVbGYxzmcLh5/wZ/Y
8g69cNkYWbtVABlcU7co4rj7uKpyLwQOW/TTasIarCdczpH7+MzycR+7zBOzkh0C
BlxVI7BosyJWohDLE7g8Rt7F980j9jiug4tzFzI+5TKie0f7xkcZQWzpxK0sWzBp
2dsavdQUI8cpJ5ukHMjagerX5mccpdj8VnunhCxI+YKc4lpF9droz/3I1eqRvWAr
t5Irw8w+ou6lgxVnbbggeqBK+/b8zrgyeFCcFJVzaKKD5r/9lyfRsNfdpywp2Bvf
LHCJ20w961vRHjfGWKE6JlI8BnMv7Ylb3adNoEGss8gCzGVosebWuvepBNu9HvaE
qckvKWoNUKpQLHRM17QqzdJ6eJiA1ROptszfO0pX7aQ/2MOqJAJrL1tpU+VKqMHj
K4AryE5cUxF4E7IiPa9PtCznXEuTBBj9SVTBkLCfIfpaOgPdIOLlCZGMIZdXTA40
hPpJ5Rvn9m1L/ljboBP3JhhzREo5iew6fh5gSDMebUPjakHnpzZD9CCI3RIj6eFC
PLl6ef/53kN96rQwrsuR3at6BZc910ruUMaNkZ0SY2crzZQGvqgF5S/jr52Qvp2Q
/P4jHVPZvggtSn0kh510IKq4JAzafff0Na0Zgd9pvjttLPOmXHl92MJ5u19CT1xG
pWR4VWnAm/XlaQZZAhebPrupbgsPJTTG8SMActlmCqxy5grKnnwUc6yHjKFRl+ET
UlFaMBMuctKCAJfsZ5GUE3tmUbzcn4+mR0PZpiCREt6tbKIVYUtgmEXps6YKMQls
sKO8d6RHCqdBUjkqCm5QgWliO/3Sxl+AjZZD+QLfkJk4dw0Ra9YWkBillY3DnKKu
H2DEUVDmiALDGJYp8I6t3wk6zTjvW/9MpZ08jCc+9wmPBpN/WSDXgKqVQWxQhqjJ
X/KbNZxMltqG9viSb6joCuD3w2zQuHq8DvXjg6tgzFrESskxFPsMMHPun+bzA6nS
PFexqguFAylyihQIgU4z9crLXezbJSyWO3+XQby5WHYWouEbyn91CPBfI7i9WW9s
t1vgB+4TZzwqTXf7c9S1SVgSsGw9bvt8v78Lcxan6LsWeTWvLlG2S2buJP7efn45
+q4lnevVMRjyNIB+o75xzhb4M2GsLabtSXOArEhPirpY/63Sv/K6shwZDDQE+Dfi
1l8DLZichCsVcCjj1L3tg29MFEMPAWUFIY57YSMpz0i4fX65P0BTqQB4POK1Y7Rw
PXUb7BTiIUIQnYYSIUPgLbVK/2io9ssW0beRB3l8XMR2ubxoUYVU0RDtkKbqgjxT
zP7wcbwpDJCLI7yNC2biwk/gM6y9PoMplLrrBFU8aJV55obE1SbPELYoQaxjMj1r
AOwhPWBHGwIs36OG0awz1vQcutLzv3uBpq57imv6RZUBCBpMr/tRnQBuxZmOBAgX
R10r1A4xtUVDsk6nwB14gVQTo+jQTcOGu5bjmovAhrCWUe6Zblu8DRdmoBvWA+we
P5ojEkskJl/cft9Fe6Bx55Nui8C6ht9HHSKE7LsnUhzC+SXZ3MTCnC+GqctSQwx2
efpxGu8+X/ivrCbEsOlCD+2QARigUeil41y/aKnIpoGDVWs/aqfFyXj49b0VXoBP
FALzo2WR8/t1G983ekBWzvaGWqlg3BCEMoU1rGAJETfXNPf8Qidb5R3pi2GLsiAT
GCwrrchHB4qrnekyGfsPSBx6uzjuT9jjU/zvBZBphpCdy48OCEA65jRe/AeStpUZ
kZmEflHxuUr7t2lA0q8tJ3wHlEQDxBtt1wICThvQRWfE629TTjnKW9IImSU6g79U
tq4rKfM09Szx1xhV0CuTgLy4jbYljpF/IzqhcpfT2Kft+zkZGTNrE6JBff4fnfIx
gF20XC7ZpdbeNE7n86CYpmwcllK3p1uulaspN252FYnko6SFHvyU0/ZkFzu7llfQ
o2bKUfkZ2qPTYefJOYlHUvhEryaWbiK8B7miL8GbU8BybTLc7M9rQJA7W53ElFoF
JOf1/IBU/ykXoAEpXiu4hfny+uxwbAhapvpf0G5xQUsgNneZcmPIfn4G4KQ5Lmhz
32u+8IwmEmTp1CGA9pB62zFmMZdjjcq8aQyublEPAPjAydhmgDrxXkB5m5IYlm+X
VNt0hFtiamnFogvHSiSJ8yD7d2dnAW5uHNqE6asrY/MvXe5Hwe1cwhlJi3vbcilJ
QDztj13S40kLRXNO1ItlpQ2wKND6mcKZJvDL9049hO6x1TiMioKJJkAnkZNnCLBq
CC4ZLqA/vwM/K93j2XibNUIyanQD0XABeLvtRmCElw/xGDS9SH44+UuRrSpfzZGr
Q+0xuLONJuxmnLmVobS75pgggzcNy1JE3Mw13pEsI1fHQ7D3d/Qm1zw7tWIUYeTR
nt8y3TMjaNmdcq1HSJl6e6+73hyPGEp6adfy+/Pj+dLeD8SpdJoFldpuQulh+K5e
8yYUZ0Pah43q3F5K1p3Vg/dss+WLR9H2OK36sUZJ4uFs614B3CFAIVpFZfgYJvzb
BVPvMZjWVH1WWGjR2QBA2MslMx1ZM+lG+aadwVmLHzKA4AQPkLnMyX+OoG3w2YAd
Qdr34z5ZG4Kg+5sDCuSWBlMBX3Uzv/4dM3M83nY6rU2FlyxpKWsm7+pzPJWAlYRI
EybkG//pkM6I2wkFsbNzJba7TN99C6Fir4DOFxzHInaFY15JcuxZccRn4zWYlGkC
2GfgGyGsf3CThUmTkhKg7DWjoBCJM+aVunm5B5/BAuQ44DthGx/1sloztjsk8i3u
nzrUSM9L6j5CFVpWL3XuRoKHKvNRc6qzZfN/W/NIhyM6IyEr1WtZDoJ1ysOpbJl9
CfFO+VkqwPQBJiR61pj+ZtIoAlI6K+zndIcn+j80UT9mrQB6mBEfHIPH7npCkOIk
Y3ooFchHSVTDIORBn59+JJw+U/n8f5GYvV/venyzdhJ/kKU5SEsY3ZeRhoOKxnmX
KXN8/3Fhp6fpgFwfHsNjghtov4mvnHYEEvRTDXQHt8MyxIQnjrYpCdx9iyaYO81t
Aa9hl1dyLHSv84AWbOpyCHH7Zczt6EXPifXWX3UbQAyEEgRLCAFToGNTv0iQnQOS
ujf3DR0zm6JnCYPciwGJk6clGXuob1K/dStFvt2KoH4ItxHPo+p3C8EYw5W/nvZn
AGctLzxE+MGCQ4e1PtOc5JsV6ZLjzFr1fPun31d/U+RVSCeG4/ldPjBNxJAxkDur
YWKYkRkhO4CDhZj7EhqnVp9uuqOwdcJAoYezWfPzIeOrvmbUcH8gpai4tlvGDdBW
RclGnrEqHLMqW7Q970/8VBQXxjOu4p3hPpM/bMYH7URax2SC6YBfJWP//Qu9lUSh
xIqY8SbyrR2islZ+TsRuMKL5qpiQ1lWwAwEDhHw9LTNtzhup64kmFix/xnI021pV
9lB8d7aUJJwdqRGv42N++c5VqbC4XSmTAac82rVNN+3PlqhIdO/tiwpCLgS5AQfV
CG3ZVWzZTzWBL3oEBgFal8Yd1l/t9lTf0uF/W0UR2/xjGPHgpg7XUtnxb3h44Eg6
zQNCVHeSfTRZHWzOeZr7oFHU1RYswVDwsQeCy0MB/f6tjPoyLzgTTzqfSoPNuM27
5h1ciR8JseOB4eKPF2W3dPCB921usHth2kWQGVH/6ZuP4I5p6i3IPXcTUtg3kk8W
/t932DKlA/s32s0hhPI0icYkTL+Pa+UnmvctQjx+1eX4CN7W40FsizkArY0v5pSp
VupxJjyMl6/Fq/1r1moF5nRxKCovFi4ctGQrJaSb8gHuX8M/20xdj2vGhPA0kANt
VajMl97AdgRd3jewY6y8fJPMjuF4tSK9ozfNKiqwyt72Zaq1tBOklPMMyruqyOAC
OOHXjbby+lHKK+X3p3lSnxBrxV2w/A3VVCMtqtGGU1CL/9BfJfff+gGRQIvughFW
cYTmAE4OTpIik4aiykHBMH01EBqPHV/+q/44DEl1wwdhsp0B3MfAg3J82DVuY4lE
s8Oh8KzoqtCzDt47ZR7YPZiRwFDeRMkwlxOAqhSU1iU78LPySZRUD9cOuTB1WLAB
DsJxfKGVSdvsLX2+xzlk61uuLe/OYgkY6X1yRkvtq5z0/cxo9Vrjy84dzG5l52cx
s3Ky7/bOdHHH4iAM867vsCBPlcST6uVm/obFkBU7FBtQyZOERdyURGuMuDF6mpmw
4CV2fXqoK2yhwZs90Tcq8qALbz+DuKIpwMngISE6znAMYIjBzkeediq0VgeE3byB
ghUUU1UdDOXMk1EdZWlGAWu/lbr/fWTZ8v+j+RiUVv6JcbltSmd3+DRzuZ1GSA7y
6NNKRslgmcPCLxU/t6UMQGcoW0JaZoAXScdfDhYDlfYCxPSr4BtMT5W88J79LuKH
deSM1d3/sP+1Nm4gRJktHLo8CBWV62PIRY5w9MeIbLSpnBPnhcgsynP7Yq4rrKCy
do7cgRzHsXQ81NfA9gqOZtmmZHLYexM5M/GbnCqeSrnsl0Gts3iOLXvzCKij2TNF
DYGxgzXsj93xs2ynV3uby/VtQhupYXUVSrlgDe4GKBXZnT4DaCpK7F05tEoKU+BT
isN7QFBcz4LCfXXBkkOG1WWOUeuVvr1LGe+WpvDQskDQkVLzAG6UtMry7ThgFtdn
9RjmzhSWi2NTK+ROMW+8bjsYK7u3vy9Kz+Bu5a5cJvKwnJQbd+36tigEMBMZq5YT
uE1TJrwI2Gi5UVfaf3MlstNygN8BCjlWIvkdkzhaoUUkkH+XHgszP0wLkRLXL+v9
jcqvEEfBVDmN4afx9T27c+SFz9rhpjKqfyCN/dGTk22nAArzZIh2hf2z2d+HJwtB
4M9JOAuvjRYmBJPr9OhkgnrJ5f6P16TA3/GvlIJIGPAU+YyoA46hfQS+q0wdTNHJ
/cb56RLRSVhQNMBspvr+gmCUB4V8p+p2Vj7wYYg2xX6ed1/LtX/KKrRB7uiwGKuB
SG8I3/w7BjcSkud1QSmDI94sMCwQ1ORE1syz5UcACd3VkrTXn9DqHc5+u46rsCNp
T4RrWxc+KpT+kVluJy1JhF5Rp0g5hMjL7MUjdrM1oz+jui36aAFMwEgi1qP0AKAI
PlZ5Wfa1c+UvLS2S1Qhy3IdGE/LG84v0SHpJK2oH+ZnyuXGUdvGYMK3sUWIEf1b5
HmOwrF/+moAbj5JhRPnXsYAE4pyxF26R9DW1aPO/VsCtCppv6EPHWe7s3PXAorqN
x3rV1CBx6igRvIUxZTzryqfBALPxxNGAM5EqIUrtUEJlab1No2/3A1K5RODgFAV2
+2HcpEHw3kbZA9HpoaaDUeUZB+WrAk0qTef9TP2AZb+UlZMYMWDRh0RmX5q7YESc
CTcYEkzn9K/YtbAiLcRtQTr8BNHkrYYM8rDxTtxse4l9ItUy4VYhi18L/u/Qo6aK
RXwfKAvSeBvwIBRH195g7iZs3F2pgtE6TmJAzTcl1roAVho4DqIEGXp1Tl3jaJln
kX1r4MQzopa9nln/hxFT9rPTzrNpd52Uj/WVrBS52ABn60r8miDfdwovvZcDQfPv
9NUeGaKnNFVAhho2oogdqB7wW+yMjzLSkz4lvoAGcguq7p8GQOrYwfoLU0Frgn4I
0Q6Dhi12Sof4hDgW10HoJKexX5jzm+IQ5BvrfJj9sIrhyrbcjrsIu4ODO/MpSbnP
WGGUX6l3o+nsgQNUqa8KcJ5Fi3zymqV68JGIoQJJuwpEG1kHqWGe5T9r8Kpnc+/d
kBNwa4u4wJjulOWVAUSWQ4/sD75RYmvg0FACKKmZIW2V/wbupCLplmNcRZgkc3M5
XW/0r1qjk6k059sWzug1YIBuwXMFh+ohSeA7sls+8LeOfpG3JlaOeqibqBIMo/pa
A0VZYh3wRYjofWs3DFuC1RFzGzOAlusUA4MjF/8YpOuF7xUbT78Fc66U1UXu5oKK
2/77LIl72AUBmlueSbm6hnJuh9Tu+7WH4kzTGtTjpQSuohmwDEJjnAfSsDYJ46Kl
a4LcMhs9SETghIHaHKwvW7AVrCpsQNYNJinahtZDTBSXeZqNqj/xwowp7ei7JIqM
aBWeDAOBue5O0MYV8BLvjbBTLy/VTAl/L679s5xpHyGswg38ThsuSnZmM+EkezJp
NatHdRjUQqLhlD85L28frDm/bYjEsYw1tEyEmOULIC13qpqzbJLrVgZlojbzquOd
wNNhVW971XJz0O0oQNGuaRDhEPQjFmXj2EXN6TosylkeH4xM/ZJnEeOt7HjIkxAO
YtOqMIHqOaEIEOkVioSzyP2UvNw/HZMKlgjFXJv4WciF6nhySjJSf+8dxrf5EOyI
oucyAQditD6UlzF5DXW7o5Qh66+Uj7QxXabqOC9tujLKqs6TKq4Lp1OQe2qDMVQg
VhUXDJwxrC2ZWP5IekwUXtg4q4lAid3HpNIMU0FD0+H5EZpT2prnr3xk/e9tVYA/
fH6iqKZYbkjUDWRWMlhpvvDZIXvq42Pn4DvHmrZeK5JBvn0jC2b9LoXwx19giA6v
J5VPFteaNeI1tz2H1lRxWXoz03IkdowvI2/hBBRQw+Uzn7hty8FT8EQHj529uICG
ptHu3b4ByjU/U4aU1vaJP9VAZihPtblJfVWnTa9S5gPDqgmC7Sixsjc5lQbQFPC4
IupDPqpnt636/ZCozp/7KtdmtADj6CC5nRs+lIlceSvsYTuz+DOz40vftOsew+7g
+yDpUHEiDFAd4AkUeHLzllCQLfBG5cZsL0yDywgOdnd+TkdggVok+332Frfpp6KO
qIui+62X/CPxWA4aV/AY+JjTLySoGiRQABygEm04gdRKpNdm1nUmzNYfuIdli8jH
st9YOgL5H5Sg3yQ54YTKQ+r60Ly46SwKdpNzwRFJqnAz7d3tiK8OrZD8ZLQe1piN
5VqURmWb7FSMAi9zuaVBUQktNO2ukPBeop34WV0NN00MbV6M77aV+dqxAVWeI0uw
x8baemfWUjag96P3psEYxMTfPl4DpC8UwaYZwiUWxn7TP2JnHTrux/Q8zmgjJPx9
DWM35OZ+wlz4OHelPtefLR3eTeiekqe5YSENAoblOvDmWadhVQguaTatSI1YjK+s
AAXJFctJWgB7WQMjVEbEjy5SYzjwuSR02ZSJj05lHYJT8g6xFOXTkw6WKUoxFtcB
2vQKmKTC2Ki3NswtZA3XCK58M7QicnvGeh9s72tGC3s4K8ErWMcOlgL6Na/4007e
ihJO4JJb6MyMsIhfMzO6XRHKAONvzyjUCxJcZ3ul1j2jLw7YP66rzoP7JKfcj3b/
XDIh9wLtpYmlJpOnE3TVTgMiFeZqmH3CdAxgikY2fdWRNdgR6abRK0ajLxDoPXl3
onqSwhnWGYleTHyi8H8+09nX8/1oqCK9CQCMAIJUpoMOdhGDyylovqB4UceYtKfe
gDdD0Qy4XR7ovVJ8DULkRBMMDdiFJ+STKxRydg6qkBEMeMrha84XomiD4IWUOutq
UYFyvVyVgpauJY5rAYq1+lX93T2535OX2UkGIA+itW3HhbfJtIyvOxz1Wl4QFkbC
6K9fB4YXKk8vQXAqyZElG/pJHewL2Z+ia+hgpPNgHkQ1cLnYOFk1JWL1nNzGpd6H
iy7PgwWO2fkKQwJRLoHXbbvGO1WuiLtDqXPzVVXnGIGQ7RzA0WFMbkia2gU4VCW+
ZMSVW4TaaAVlKqQTxFwKiGaBaspNkLxpmQKWNtl7UZThAK+kvGSI4E33TnP6hMIv
IJGkTVAPt6Hg4OFr3deQeL3uZOmVgnEgXvPy9y36nX4Ypv6idq4a7wLvziKgxRT7
Ueq9Gbnu4DeBgVDxZFDX01UUPIUubMiJ4rwgklCOj8tioxbtc4ITI8VJeRUNs4TK
UaELRsFTtV+rYb4eToYa2GxVZGzSO9dE2GYGw/ILlu1x1sP7a74kFEtaocX2e6aJ
2gV7KAvnh+jZrfb4OfaqwzZvEP0L/7Yt2/tA8p+1i/lVc35PqSti1HArK1XSsh7Y
vHMrzTjQAHqb/5lYfwz+YyezlcycZLAZ+BJIoKG3fQ9aHgJB28jzmuDZ6GEfWT9Z
ufupkc+vYoJLhkY74+bHlc4cLcMx5tVamGdcNuNKYbVLOip4RW0K13ITc3XEqtHA
SsEfvTohAjudyv2LxlwDGanLjsoAjiByd0DylXS2fpnq1vAwCxTcA2fgQmNkP3NA
RwE8k1tGMqMW3od0uie+Ye4OQfv4YZyCL96oVC3gTXWmHrGDGXSBsOgUuqK9ZexT
O9QQ+doI/+YvhO/R8EHRBIDZrZAycFRVkZNdpMwCeUZotBLUPbOP8lw8s1b8CPJY
sj+/aKefa1cLraovhm9UWpn/hEB4557/e1Q3PT79I7EGJoxRS+N6cukB7UeKxOoX
sWrxWd5bdv9jmHoN/gvHLwPT0fkPw4FRHL3rRzHxGUjYgf9ADygQMP0/dImnj6lS
05httGilmtdihm4bPeU05TQE7X4zAqMHpdYYWn5PxAus1dktF2lAExYo/iFb1XFj
H1eXFfCHd5oNjN+jqesTLDMzh46fkR2NgELUqvGdk+SiZ1VjMnbT3rdayuDDraJJ
cNBJxHATEX8RI+OiCVUj0zGYsCKmKxAsPUX//4KDeSxKfsMj57OHGaMslXuKY4xZ
afCBjOibuHgawYQL1yH2S9j7el/Bj3KxHJWrvXpV36qrxqiMrZEcb4V0jNqDXzHt
2Ln4a0a+W+MnOOSZT6DSDr2AFGZHUsanROL0ZT/36qCAtUHOCXAeSOeBurhWI/Q7
GOZNqXWpqDtN1osi8fcVk87TtEwZuJJvU1GgJHaQ9vQu0TgtHQZ57bMKP1gP9Pxe
863H07nRr05nHOTceUNDO6fdA/FZI/kA8SKvjKLT+LwsRlEbjyVgzcT1PbkJS7Jt
whBr8RoFyH6626ReY08/PrfNySm8uzkF5Ub9HzcSxj2AFZwZrdpSg8XcqdwJSuW7
aNYJ45uSIMVmyOz9xWC3H+DmJVj1yLnv7G+pcNDzindlMMA4KKycyzxckNRqoN0v
y5MbSYXBcS6cbdUSTVeJDF8V+sByn7Bkul2suMjC1neuz8AN4+06dh6b/9HImfWe
jj8IKQw/36DWuM8D2hJptfWxSSkCcaNmaEMz1/E++KNVfVsFZ6UMIzzTotShow9k
+zl7cxEw+i8uv4sR5bgstFPxVLOa8YIB4vmFddyEHZEo9nKgs2RatyWqj7jlH/8b
WPWw2y3DAqEfDd/4e8PTI7RzKt4KLn1e4dfaCVSWhIHf6/H4dImscJfmlwXWU/ak
X32M5HWIyt4gMXeI2C4mJt+toPKDuJkZo2LRvexyDwkU5fOXjXSm4pQoVq0qzoXm
Da6vFZWel3GfRkJUdCI+jzudoww/VVnR1nPcktdaxoAMTXKawYrxVKuR2s48MpTU
EZt4YoDjP4CZVmyLoNnFZJR+cDJCrxbJtkD2G03kcxpd5ATMn5BkyIJrZJjo5XGh
5v7fjnZzeos7xVJQnEp1b7UQIAVmpO1TbRN6kWgaN2nrg0FUUnyuRR4rqylxeJef
u5YlJeehq+ji6UUrZpMzY99HogvvowydYcSGiUWNBQMwS89fdYlI9/HQIqsosQ5T
MopSLsA3IlvzSSDX5l/yPynbNrjUtJhYdKy7htoZeQSJKlgkBQ/tYSlkopTRWdRK
PVeGSMsJuW0D0fKW5PStB4B+lBR3jACVcucImoeM/IZOKBlYssBrh4roBmQA1oc/
nq3q1MVMcumo8ye6P3GVeWS26pI6ujd6zRk75PVRcjP4lZWO2WN3TBWncyw0uNvl
4LJwuhuEqqEVkKJv1hiSDYsqBqIZ+K57pGYlftz8r+sdYsm/ZWO/D9oGaLB51zI3
rbbDiysYniQnjpvJl4pzU87ui9y59xtx3/FxLundZaJoV4MwHr/eIaMfe4KC775m
bEdZ5sy4rIAnhrDaEIuu0q2uKtAOg3rRU0nj4ktcip//zE9b1xLbtJrKAbMUKN4H
HwjzGiDozepfrHP9UugJCtWNJARvx3rTgcOKwtfc3NwRWtK6A7+jOGCxaBApFaqE
KN8sAOv6bHPtntgKOcYjbA7EsAkvfN64UuAXVyDlTytrtlbOdmNgiHHAmLKN8atN
q2C5Rbe0kkIdF5UYeR2a87NwWXDcbYg8zfwG5xL0Po8Y8vMQC+4oxZ+0seFACovX
PfU91brJojorPYCmRwlgVV46QRU5IgR8v2lGvyLbq+Q7733O8yh+cj8+D6gH5NvN
JTIIqsGKQhAw2Q4FgyLnzr9doBbeSdX7BNq9r0K08/ZNNIso8VykZ1wfjsYELz8B
p9neVFwk4DcbG5xZAlva51vxnYf6QNu8tOxyiiE91rbQa+vIQDFaUmL4hDJuyhdj
4cZJ1tKsyHPdNT9fB7OszUtCSc6/BQAl1XCvgNu5+VbN79ckRxS3GDdRPgMQGfc6
EM5rlyW31G58Fi6Eeo9gBN14esfkqnsnqHnKjGKHXJ7zrSDEGGS0j5xDKWwXZKkk
W1R6uul7CYm8IKPv2AYcPJCmoHtyqldvzOMZyonMYBSpQxv88bW7BCsFObSJK7Cd
05EhD4LleukhJYylO07VL20Uop+wPaahy5FYfW+Pf+qGSjicZqcXXwfkwkU/wwYX
+bqE+HFWu9wbn7uMNy2ufXOmZnjF+LNfv06gciRflGSQ/2BmERJDy3MAqSl/8L8o
ly1rLurEbZNXePrCaDtRV7VJX3wgFzUKFQTGS6TVstA/10pDxFgi0khqrZs/3LxY
ArNyb5veFf4v2G4kkSZOtwERtEi5mwEidSg0GnuYMm2sVv64qqMcd6VuxyFuuZgX
MhdIWpbXQcea55vmyJI3PXF+/XpRh+5146gsLDz8x/i1Vg5s81uV/Uqjbusadnc7
NJ49NZnSSt1aJ52O5Ze6w1V7d4vm4Nr2R/7nZUzMUamRacHHek1SraoqVZ1s0rsH
GWCQ3NAfbmaPNbL6tO9UgJxBDTpg0vW0jGooJHiAIHGYCMKRv++1Xklblf1/wY4r
v5mF1/OuqQkCujnZSWMrG1XUa1i0O3Lk2yTIshO6jxnNidxK/dp4QlzqkQUogjbf
8TebrjneCQmTPTLZ3bd16duy2ij3gWLNhNg6J9Wcy+0KwziBRLqp2CutqkbUeoTW
tJv3Cne6geiEY58mFNjnQ9P5ZsniIPkLJpB07pJEYTGZe6Kzh2jxVKxj4LQzuA/T
RkqZY/NfcBHsfHqnSvNvEBLEOagq6Vc2gaH15MtoG78mI/eZ1YO+4cqIs+kPupvl
xun5Q/RCC0qBLK4LVspmcCIq/d5xYtX7UQ5nngAraegGvlvsx1oGRAR36ZwldERa
gz8xYqXDPSbKnm1UvqYSaXOYbVpscfnZhlfVytTCD1AqCfvsDRZN1FzWvlDt8Vhu
X8fl2V/eeswkZXmXOtOKZfMeSR8GwNxyGLgSRSt6L9Tk9WlFyac7LIbIwwqqieyl
yLVVwG1VRvYdwEWVTp+2qGgmgnl5uHNbK68dmW7B0hCplhaMfvhVQhi4YCItPQtM
yu/UQEGAsCg0aEc3faURvxv9BZ2Cv90HrWukFiIZjwvhRysfrMoxgxqSNwu0QXSo
cjlMzGHpLN/IGctd8vJtjscT1wnoLzFMhwgXvQaD1RBCyY8Nf/dbv5l745LhefFA
JoJONMsJGYHbfT3tZah8fHzsqQ6hFLd3Q+e2+C7nZaTJ40GjvLlasbP7SjyQWBao
TJ8jN+NuC78EfZx9KDygsxcNQpujxJaiCnJcbkMOY9pgwy6Hc78pr69hnUCx9fLq
BInJ/G4z2T6qjjFGGfut0Rt4f5FCp5xSFmZLuDCoH6xw4MBuDkFPbRX8rmktzuTY
QXPZafQ8O1w6hxyimn/xoNuPARFv9rv9clVsbXKbtpEK2bxt8EFL0FAXln2Wj1Ue
dOnMWM915uI/07Bjq3t09D4kCHWtHExVjGgQGn9UH/V4Vw4TkKUjkPbl3xIz6mGS
cOOvsV8JAOyHgfOxBPXMNwgl5nHj8pImi9Z0mQ2K5HSf0w2THFQnUa/zhm0qBJSe
m+7p82SFWCljrFrgMyonoQBlqd/9D1ERGZiR6JqXGdGwKo+xB+1vJmGjPvBvi7Sq
/ASVXMzu5vF2XEkN1dT2yhxYhAyz3+uKwr1lHr/KXOThWux/6iujuqrsNlaJmHQw
O7IJM2ERy+77ZlElgHqz7K4i1qMYQx7pizD+dpjG/KwiXmU4q9XAdbaudyF0ZAU7
w2BGIragoBvIFER8FVX3qaNo+Vs/naIZ8KUz+eZNB8Ei5U5y/eIRoNvHQQ3EZQhp
o3FFUei4h5bp79IAuBIWK5hZpkhypl5YSzEUdL92WrGY55TbutUbSfGd4QwZ++/N
cF6NNXhmDzpGFJVuh73fLznsuvnI9t3L8E2A47QWWYF8wGm4YYHHbw9uywKt1zwc
L8DQMQZWf1guhFnRykxR4tlnlpnNEDBH6gjlYJk11arc0twP5ryG52TsjMMpHyfR
itSGJDW6ZSiJiEiS5tDCPlZwZouPfZ/Lkb587eIBHk9byE9H5XALJKbpgI9S85LM
iMi3FLr+NIoWYj2+JBr3RuMPtt7QHgF6aKy05ZIcBTa3oSoP7ghc814OEkcBJk0e
H622RGm/ttDHLM00omWwQBOXPRP7zwMle1IL2lhrGhnAeM+VqrMPYk+cwGGh500K
rVgme4gjOii+gP5LuLfpYiDYcpU1Nn434fnKWun8tFZAYTYPWm2jPMw2feMUjFtx
5ujpbQXVYUeJ/ZxyhEpCrPXCPBW8GbKP+02etFhQfg0linFpGzQG2bArVhQ4kQUV
s8ebRhnqmD/lkvJjhBXYXHjYV12Bi/x2I+3nc4tTUUZEaoQ9m89T5rcLSiYVtABO
ouGi1Y958goi48grp1W6js6VNY7sxZoLhRbOjT5VMgdxjDi+8DHM0hs5uG5bksom
PN1+WofQLfve/UH6li/IR5zQyP7KvQrnA2tm/A5+RBAAL0Itf107Yve4hr6Bd8Wz
QLdV/Dw5mz2v0VEX1PSPJDRWbK5KjdPVhhp1TGvOWYNEksSSop6WfjcvfdyWxEYs
H+frhkA10FwHSfBYewyy7alSZnuUxYB1+GwcwEdzKHkKGvZNcuggnSqd+qDf8QKj
9ZqNK8Ue9mD99POpEm5CuvGoU+ngQDXWvTTdP211rNtgaOu7J5vPKp8TWZDnv+eK
qBsRghVptdvjGSvBBeheOY0E/al9fqtWKKadhlCxqrpmv33GD+34vHv30t0FIErv
Re3BHZ23GYN+VD5oJEZAdNdFroTXC3BpEGhGUN9Q1qRuCTTr4EOD9YPKeLa0kh2R
rC4Sd747jIbAaWxK3BLFrjoITbZhLbXEA+NBKpFD3nPf7SO00oIYR4wbKzes7ye3
R/dnfse0bVg2rilnl/9Btt3MvEEDNGgdwjsElUhuP7ikdapNDEvNzjSL/FMaJk6j
/dkRlxZVGKN701IMhOC8CS06nfy/Xi8NnBAi44xFiWD7ikhzMMIGHZYHHaeVsFQB
mMPlI1AjrmeLocKJBVy/bYCM9erGlDfoOja9gYfCW/o9jb9P0LSbTXt7saCgqLt4
20Unv7CTLrLbJUyJwa5xlu5UaAO3qChqu+bDEqPEAi9gX2NEDHTybKBCua647XBM
pz3OpJYE1vt/qYM2iCi3USiaelDn/HheLlVkyJI/6vAWPdYh6/YbTcAZpP5h5c/z
G0euqA/a1QbVVLmW/6a7XdTwI3nUKD2bDw+qwUc4dtV+iFgH86HjZGVlv6otUAUw
NeH70k4hywhvl099vM8pHROLfeEJESgrYootLMATWTB8bFDl7tw9TAAg6lqUzUdg
9qbFiKC3D9mMujxy78eRBVcClLtk9E/hj+T0Cr6G4No0lYsBhk6OeAcXAp9P4xpO
kfvWkkjXf02kx/F51MksGSr5YYbXyn93RLG4LxM3fpFbgO3le9itbrpC7R0fVFti
kEy4Z7bcEdcm9Z70VSoT+V5nzitySnDuS+X607GNR4XDXnL6XqzMZ+x710+Yuy8k
28ONKMr5MRBz8tGNh1v1lwu24D6tQp2QP3HZZcIgYNYfxTbih3R3dsLYz7sEekK9
gukOBZUYbvmMP+myuuL99CYTlMrFaKcBBIKRDjal3AjctX13StzErJ0VY/uNhg97
S+APjHWKm3B/0l46vkF8lVsTpBu7LglrVaYbjCQnvfhfrbHzY1Sz8YxvNJOSMSqL
VM9uq8JlzCOD0Br8ILSCoKIGXERpaGE360bzaWym3rjBTgiOBxPZ3mi5F8hhrtTw
jPwO3WyNsy+0AbGXGcMqdLWZbGjIenbYxv2vGKpN/w6aLwtClpDQOflEPeIKTz9s
niwydiSxNK3aZ3cA/jup5+D38yHYzHHABBKY3m2Qsu7N4PMYmOk3rFUSyiYMxOt2
aN4RlSUbt3rIhLVU6VRbIoE2N7tQGIN7fCbcse1kduYCsUNSj+Kz7+Ji/Dpu2g+U
sJVNih7Njf9lUi/3agpNW8ORsaNKnMjWN9GFBYqbgTea8tfRTJuvAHY11MEVfg5h
aD3EGLr/5/AAjMgmPSG6VWhdzPGn2xAKoIyYKJA98ye/PhKPb4pIQ/B+JooBIMgL
OV09MxbAKQOWzmaLdlBB1PH46LoSyhkG47OpxPq/gQSc4kVDm7Cxitx975q7Otrd
IrEKq2H6EK4pDyV2KhLD+0Ys4x9Z8qfB7aLr5A7N1xkNOvr3g9YWO3fSP3jRANZL
GDXz1NKPa3NQUUqlBWTt5VUTMRBIIkLgGZ4SSo3J67xPm7c/uqO32tQQL+kJb+7F
UCcLGtCDSjOQLzZBfDsNl4vNMVP7jHF5Zo/9hqf7I6t3uH0q+YjBITo+6DWZBT1h
BMxiNx4p379QpkDQmwRxWp2PluKJhKoiH+0Jbr3La1Ukm6Tt0NSLJKtrX0alpZFx
ZCTvi+3QdJAJCaDthHiU1t3oxEGwv6KAv0fCTPCzo2JIVnjdF30g5sLKucVBf1Lj
iwEGF0LmwRKsfihiptzCW5RIdsWt93mk6ftJGYJfDGU7BAX4esM/F5k1Ia5M6s7m
QjhSC9vVyFs3Z8SdVhVkpBEgQpnLd/+upO0EHXW2hxpH7eIm34IJ+GvL2jySb4ch
z0l/fIOh2pL2TjBTp40941ffcTVR6r5cH5mkzEWI3GWXag2zMEfvH5aTtzJP6wOj
k2DVPtIrsPqW/IDaBHO5Hbe1Xt6B54uqYoIJSM5W+CNhU77RNIMn8pFqD0F0UESU
TwV3a4B/zXy60u8dP4KyretGNAMTgvYWku53lyCY952m4PrcuoHgRJ7ZgW7alr6P
AIoU4s0yihRLKXPZeHmu/NgBikPpPYc+c9BYicR7usbnEoNFZBNPI/CXqjbBpNqR
IUAAdGgRLTi285IAG2KTRFoR8vo7Rr/nD6zJijKfAoIITTubePagwTxrOt433a2K
q49ibtKa//dw6xV1rdzYzMsSMlMZ8Wj9tooLoBREI5xz1PW+ZdbwHces8PsiRxTi
+AOiouLwVv+2nV8Pp8UNP3wMJmB4o83kWl2s+VK08gEJt6m/bZYjWcs3BkcxGx6j
iWtkSJwANNKoyEpzhU1Blmt+N+cvfjc4LccfPCKSZ0SOg/41S2Np9jWOvTEhV8nG
mdEf/GsfasA/zl0T5/eH3HdHH9HQ2I7L8Y8O4lDpcX0qXilFXt5DUxYuUggyZslT
f+wE7uONRycOt7K7v5J1zGHpFzD1ibrDAEEXMSAdM40OjYs0QHI0NSXbwcKGDk0g
PmcdeNJC2Lv5YgewTwgNwAlaJg5j6UR4Bcp3uL9jis45zfauHtC7e4MXBQFlgFnn
gDYj5yjc00y3ms+m2shE2h76rSMDs17Y+HCQ4v+qoFTBWClRdI5zbOVBrGwSiVYT
2Ag4TquUGwDIEyQyWL/5HJS/ArwPN3/i7262JWZjabEa//9VebcRbeN6nzKn7D+P
8tNzs+fRcWAjgOsdPP7vJ3k3bCJxKPQRs5tC0ZZmkuwJSG5Y4aLC7gNi8RDcahlc
7+OLmITe8udgY9EPwRCmVlhnhmok3e2/URsqo83RM3t3Iu9OHRxYR7glwhfgiw96
EoQaXftqY4e8KMOgzY5ASDJ0FjHHgH17aiR66OszRsrzRBDN4TaghL60do1aqsC+
V5/b63R74L9OO/eUjdcMd/Q44xAchIA9tKKP8iMW+19YQzhPpU49kYk9ds6hSN3U
VZuWGJSOSDHTrn9KXS/r5ig8xYX8uClcyLK91tCbUn2z3zygyNXAc4rF4oN5xzGp
9++5K/iUrtaMQETB1kLW2eD1eJztJCyon2KNpKbHPT9gEWmnan9UacHgIumxPK2p
luNGlqX+98BG7e8cMP40Wir2ShavKjUOw2Dn1WYPrwhG7QjPEGGGshmPWDtwj+cj
IkOaX80dei+016kkgyrx/ktZRhN50n+vm9GwAo9qM3EnYwV68ybbthjXXQjG+pNg
C57hpX5eilxMK+Bvu+jL1DNoUcrls607jN3haLSZDuOYfct3sXQqIuSbL25qmiKx
LMkDm17zDDZUIqvfUs6JkWWqpxUc0EHaNE03j0YVJWTNLPrluocI8/qj6PKcKWZ6
Gjl2qY6CFjDIK7LOm5ATi1DFgyGaRNk1eDMeUxGIizVVXrW3eXKQYMiDkwoFi8HZ
pbmyRC8LsSpiaE9ArAwbNw+pZSuxDNsDy/fwi6XcbuRUpAwEKlLTY3AXWkzvtKxy
L8tuzzklXLj6wrcuNPFmwtvah7rX5XsaEjsxcVEHP5FhCaeuhVss7YK1JuFeUKSb
6vymli3+tU32UeTQIqAD0u3Sj2xsC1ouB4C/KpK7EN2L9oX00WpqUQmlw0/67Euu
rVFqagB3ilVaPelXL/v4fbyS2KNwHDDBj4g+mWuahsN3lADIKcvuLOcJjD0x1y01
moZJSRicetA7G/CFzF4TJpmM6rVl1Gvr6a9bf3STg9apuYNdptAeEd4B1+lJZ5UY
sPkaEg13jYZQcfe0sASaGiy6qhAArQMZ+v8x4S+bJAc4+IavKFpy+3PVKKzGiHr2
BtY+l7ZMrKi8lXmLIXMU9VBnYq3OLBplAzCqVAN5wsaf2S05v50/1MYkTyt67l0s
3rb0BuqfNjyusm1dU3khDMdxWyI+DW6UAMv2t7AMeg6hmsPoJSHGxmlRwF5So0LA
yhcWwhzMTwt8ECMLF2HeHQa/Vcl/88ZoIni3aXkJsWtYaRDTCSCj3ev5AFqzmWSu
q7WqxILnI34OXPE4SQfDyv1G5//eHliRx+iq2JLKhBTGKUI1xyAgWdITNxlCNxq3
7C7I/76iw4P8q+vlEpjuCpzOqFUxa4IVldncG3/yp4MnlH8VuxAb7Q6JSdpavKMT
cWqJvhG1ugzYrWo5f8grcXsRkkyBPpOaTNr67qDEpKfTTOMNbh69wGwu4lDknZGA
E2oFtKrsrZEKiw+5IgOgpUrgiqQF1nT/hqY8yCQse8alEzAcWY1Zz06gdaLaC0Mv
YtMSfhdr7YvekUXLWlUo/A/I+mNuAOyUfk3IrMtr2urQK4YZ2Yu552Xl3wVp1lmr
wMpuXWOAA2h0YXj7SUknfRwRyxFp4EvbDT4+hQYG570bNFt78Xisc5en8QVc9w8L
5h/ulGnKMj1YEVP+9YFXflj5/gprRJat9aIfwkslMBciUuIo+UzXA8pU70jHF/a2
eIENwO8Nq0wVGDBihuqikuzqPKZEfoW4B4/ovWVg8+4xce4YyqhT4omCl9E7fApg
Hfqqgy2Vjs8OKuPE3bs7lIMwJwyEJtaJCzDgiZ26HS95P1mvoqsnwEgBL/VaYG+v
Fca+WCD6ELOgFF85sGRgJJYhGHP+EWNG0UFG3tkvlb5ZbWu7QxcuMXJAKHrdP7oq
E/M1fyZLyBKz2RkKdGH0LsJD2UdY2m0M/AXuLl/2ofxmhVCLYVNeVym9MICe4Y8i
t4xKymRGfDrMD7YLz/epdbrFpn4CWVBMA6+rvPbO274MQwqojneoPmxHBnYHa4K4
XllotUxRMl/x5i0YQRt6WSEjkApIeFYcKv8rCmFMeCK3MMnRV4SVG6S6U5Snr8Pd
wHAN671JT5Dslzjtxr9CnwyvHzi7vhUYo6pZWZV0gPd+iGkogKtDvkehBq2GlnTx
51iFJPuDp1iiAfT4bhr9Tnd+mrEslDeTHfUO9w3acTSU64o4Q668Pyeb7bZkLAZd
MruVUPH6wJT11V8+ySgviXZd0SyvtrRd2RyyHls/Y0Q6ufug1yO2Ev4i2yRHLWmk
Ao5bl+rCuWg+jb3gvZklwgDVEPmxeSDQpi0TI3UkG6D44c+lzrWh3NAzyu7+BtCv
BLpevrSQJC6YAm9xC0DNSRJatds9roQUnWbF6oylOHsDiB2o0Zoee/0AuXGqZWVH
cha7gtn/XwDQ9CTPEGfUNPJtXHZriIuhKNeX13Eli9NRAp5ywKmWe3hGxGrGR1A6
jRlcSb7CMyqotf3pZ9d0k44P8D7ofMdsGLPONmIHzHeZL4VTx2o8G++DAwUZmuA1
NEbqxfcEolDfm6W5+qO3uk8v1xVHd5Hlm9c2iysW0RKMvRn/Z7FN4upfr9DP+om/
6v5geNZMzpjaE+gschZuUOMaxgNcLdAgah45PiXVvolqKTothFHH3UBPW8Fqg5vE
1ECAlseqt50VFpiQrkKSx9eBQyztXer4DKfJ+sgaEvIMb+PZrAtrY6K97iJO/q/j
HCBrfq9eWM4Yp7dWToL4nUCYDyCDrMcjQRd9EZnEOSlbmvoUKSV0y53WmaALX/4E
DoNfuSzmCYmFmdH2lb2Lc92usBlDXcItGxOfOO5EONdJd7N1bC6FWyhX7ASUpdCv
Xu93P14r12wynoUmo83XN5dAELcAB1SfgHIkSbz2Gkzh9t4tJTEkAno1U2A87sKb
4CZpATI2dcpG7M2BTWA/aR1ELPnuaJRNGUzhCVG2/b5THlJ0uL6sI0vQn8QUPSiZ
ayiruZay3XpIMhNPqFhmku5FeWpiVzEQQHkphKbvsrSVW1Cqrf1rrB4v/uK9X10N
XYVA9ckUHTi4O+t0rD8OOHqRBMWAFC8tr+EEwliYaJIFBmO3l+QB4GtMarxYd9ML
vEtxTfoKNMAyJyMfjTAiAHFXqawQYwo3fAyhcDA1S9a423qRgMfpjZBl/34ifp/y
CwroTu9LfDlIi6wys9fa1D+PON/0um8XE6VcYBlwOoxrjCZGw3UUIQzCGiDoUg13
1jZQjC1bBYdIequEvO9edTFyXHoaAfQw6fl3wPWNwT2ziQ9XFbJ1XY9yVFZdegdU
csJZcXTZMg5iz8XhmzAw6gDLQBPaJTbZm7ZOOnIR4o3uW0svCFOs8DhteWz6lT0q
00yEIjuzeYJdZPjEw+zYzMhekojZnw+nfLpOW6iEma4RalzIVVWYD/BacZp2n0dd
VR/n7SUOr+NCUYHo4wskZh6r3lJob+do3RaaubnPgXKwCMNU2GowO0EGJ0VvY4ny
KEPjPh7za2jKTlBMFKPBo7t86ICxl+8G8WCCf2PjnvGXPXxRaStox6/+ezh11bzL
8jJNRMuRYCqu3Wb6B8QfIcYLD4I5rbNUtnvgKyACNj8ZTkxXocdrav/mH0Eegn0J
thEllWx+/sHq7oVmUgaXbV5WTuELmyRac7xygY1W8cT/Axya9ddv/+ckhnpuzS35
0HM3EfdTl2eahYPWOpIapYqbofS0w0uT9qhP9i8E+DiUpSrIZcmeXHxWRgwky7+s
/qW7lAneq1d/nfoSImrNhfzMJSqUrGzg4VFe1EsOLpiouU0jVJHc4H4I+PkCQcyG
F0sF5JHBgFxtm+320VmXDH/pVdxEDo5gdIwKmxpGfGhmSTVrEURCANSNJp5Srowf
cLRz5WOk5DHCQ6nQs/Sh0fyhBc8NGnCj8xl8DnldMNTDkUcf/MpAgwwNdylQ+xpS
Epr7qoi+cbHiYbgafOUvqy2wD/WP4zFYic3BPHv2Jio9VWtCo8R+b6SC9V3mBjwn
OwKFXp0u32Uxak3WCNAkaVGKF+2E4+LdUhn2SlpKrJcPWrrBJ8u8UOaJqNOhuYBc
IBK9nduI4pl8cvASf3vGmbZVgjj4Uz/D3jjh6fmCVSPtzMaWmHgRdq1Xv7fijePI
xbOny3yGqXznc8VfRjWI9QLYbXx8Rj6r8Ne3MWmvWjWaUlJ30ZlyWx99g+PlIov2
JiovHVB91667e+MB+VxwUBKDyBLJ2jAondFF2FzDwuCt+nXhFjT2JMN21+7wEy0K
UgZfP9Ftxv1bmczlW0VUU6Z6B2N6GNoiinD6SIM1HEphR4l7pLPlfEPfqvpVjlX2
vfA9hFXxdDtX1VhyZzFrhlFlRJ2ebDbOHlpqdtbXKYAB6+FKB+g7BdBA1DS/ROOl
MyCnakYDveFBjpG6bH8tUvvr/Jj+PGLh6yYxWaMqdchdoemJHqdf3OdGeIoS9YlG
blBaOj31cx68tDw3f96zTdRydfbBh2p6OSgmrRevZhpE40mhkitAukBXzQHUJowc
tzoBPZUCU1f90gKOJ6n1kHLERIVzfOglOn3I8oSpehVmIwc17GF4VrppJImZ0+W9
aXUMI25vAwadyII88W6pN156F3zBvCTL8DIyVAkt9tX9yxdNGH1auAYUEBPkjbfS
S4zrji5gUAvbXdNiSP3fOAX0m7YC6bdfW3VkrBRaxVVNIDh039pR2PDhp2ue4hm/
Htv6anGipcqlkHCB7kxlNvMCeG5gLpnsRYS223oCUH7kR7hcvOZXDy/i15Eo836p
pmOlbOmD2bX9F5wuazmIHs+Ldm06KGIhl8onaIyQ9JjJQXZsdC19/YufWMQgVEi2
cfi2I19Axef0tvHWQ0a59csxvu4WOxc1lPi5tYjaFsVMtXsgsqCGRCvLsqNABGR9
KbcckBejz98XvYyOC9jVaPutiEA+rXAsRLdz8XWo9enye2MaqyDy+91Jcn2KJ3h8
SPweF5v/4kZhUYu0nz6lfpVxNfxkQ/75Uctxnu0juBlBIinBNYmjfqh2UGauBoQv
ZSCW7zMTpVYAXkOPVF/8pXd878Iijwa/9qaxkSHC9msrLDm0mRV6m/BXnzMSgmr8
WRW02Z+kBVOUPCGz92G5XJNCYjp5OoqkkyYfeP9w5fXPtzC49jKgb5k75uTDk9LN
6/UwJs7niBPMsr4xFFAEP/j6x5YrpIUXTY4JlJrs1IsMOBczg2WXj90ufWaoZg67
dOB1H+kSAVAYglNfTwLTGomAP78e6aeQY2jxlkkeVShmLKjN+O/c61GoesOk7GUT
YWupC4Nfgsy/FTchi5MmDT6T1OcraLxNfCwzfxiuKg5zu9DseWVxVEVsC7pRvT4C
jSqvSvJ5Z9r4KGkyQKE6D6ZI54w7bSh5Hd/tBeWEfhbcDqHzrwS6nAdHh7gp+ixg
b8J/5NXkjXKzxCL3L2FYuRb/VEdgAeshSMfgm5b5e5KRnLDmRn9Q/knhr3gGcCv0
SbKFmzwwu3MrTZm5c/ZiEVEdYsWADq/1b5357VBQ7oo1TuXHjiJik0RAyK3xHjU4
Re1hCTipLIODJFMgq7qyUKXAw2fVPOarxSiRpTUT9P7JScnv4FdNTvZodq230OUj
2EdBEVwk/HXGaCYlUcOHU4N3ML9Dv6qvn0/d2Se49jozhoBRuspLqdJ4FgSV0FFg
YHrEDuN1uZJXZBLimdKZULVDpMp5mSRZqfGUvSFiy4eC+uPmzCg1rKcaeI4Aisrq
IlRWmr1qpCWjh5gQKOqZu7Mvz8NLh0/r0n6H2MPN2hctzAgQuJTxmSeF2XtIO/ap
0lrfeITNtwAtVxCbvrGOdoGWjvB8rM3kLABsOOcfnmKeLlsMeQ2/flfoaGc9djzH
fFLlDSIwphkKhJnP3cM09m/UbY2EabNICTB85kJd3YZ/B9Ik/COJsRVCK+7EedUR
M+lfuykWRNg82ENAsgwlkm/AUgedd03xtV6rQuqplosg/hCqYywvBOny2x0Pj8V+
oLHQclXzBMWDqofZXsME84Uu56rC9HeJlsPqa7jxU+aTzqkb7k6dyZdPA73j5o9n
dSt+YWk8AjYBn9T+6HJX4ByqlTS4ZF99QgE0UV4M8vnQ/ZMJeuzaDLQe+rCWM650
CUWvNsGCG7umRAuA3WFtbs5sGRZ4xtJ6rmacKfOi/dcj6ZyGCemwFd2jdn4kGFYy
ZVxikhqkObq8bJpJ0Jlc8nxtmcgwQx+kZonVdR8KUSraCqdO3/GPglPBaDTTKc6t
cT/mdPmJLmWrknjGZr0YXxho8jIsKM0lpQWI1XGL/JOsvP008pKZEwsBYqR+ibvU
DIUP4PpsxFuZtbK9N2A2DLAmov4wO3zU7sCfUe2Dac9Km0b6p1ScEW8qD+s54rhM
VZa+SEozZJTuQpPdOdu+4yqPBdmUDAx7oZUpaMkHsuEDSi7boTaVIIIpX1fbvYQG
7x2ed8A82SQ6amwNxijVqXArj+xPo/vcGnruNGJBYnC2EetxgVW6k/Lb/a39/Ua5
vvcFsHEFrTFJUGA/wOmyXqZFg8BbqiWODdXBJLBBdEzAMoU/8T8ueWCQ2kVHLrH3
EjzE1dxeWXEGoFg1hFsPEIIEzDoSdV/grVhbeg4UL+oBD01RbFu/EmzjwEUM5FXD
622hGDR4xeL6xO6wNTSya4QPOLIkxr+HMJX05MPjoqjCliiYL5gfv9lGV233XfmG
qQ3V2TR9fhIN0C5QlJvHcIhQtr/Qyhm6AxzRTqOog25qwdAiTfElYkEzI+SKnwmO
TRzTwxrVAKmoUazCp0axKSr3jLItvwsScwnH5kOKG0T6He1s2nlAWSMSN+0guC+0
v8L8XVwD+pTQGJKEzkgx6xzDl6Pkc5CA8eyiQBn0T4kgUan5qL5EPfGiq4k+pY34
wNehxife9Nxj2ISOK6OZHYl/wrfnE8kAfn/P+VOUvyCOWkRalqaziaRl1dyoiDHp
KWrSKMq+3/shRuoJwQLY7fNiCBqhnpFNjwSbeViKKJ6g7LTnbn1do6lGbO0SIHtP
OFHQhfAgm6OiSzhjZgltmG/mzawbwyj0OKkHdS1qoJMks68rNYm7SzqnJ2pVg5pv
/3ysPP4tqNvFGBUeCx5mb+oZImRxyHiDeXUQwH4A4jnZGAOKyOchmFCQ0//S0eyi
lDMphtqIx9NqZ/XRl/l6yLdw+WkzPQLJ2oFk7Ryha5YQnbxjT+Zg0tGztPheLHD1
b6WaxB5KixdatNojWkI7U5t82eF5d+tRKAyN27Mqz4j1PSYNrSpKYIBgezPSF470
8LsM9OdINE/3ok8re3veeEmA/E+N/a2Yaw30txbpzElPhAFycYnfvmF5ePj5uCz8
N9Jok9v64BJjszBVSGyyMd1UMPMr1h4XsbHznqxaOQyXfpRlhbl2Ms4tgTqgfTWh
dTJap+pZVJY7Hsn8zY0B/4VUgkc9SHc7XmgBHVrq5c3h6iCYuobNpB0dLZ9UuK6k
BuZNPp8PhoDycupCFGpbHD0JNSBTZcVnMVHemSsxJjN81eE+NAYxhEfn1pKVGCTM
HceVIavI6UhVskq/nridYQb5J9pUzRgrZFhPitWtc/SAGbOQuq0eOci95xUfez0Q
WY3TSflmcxNR5fzzLEwHDm5/fTlpHrnG5IgjmoAaTdp4X5NEgoVpgL5uKNWMK5MS
C9yIn038LYq+EwgEYQD6U8O2hzEuoRaI4a4ONtYuwD45BPi7eYGrmXwX2QaNx8MZ
zxu6YxYtsTqWnFBN9eHDB+fYM4XeKxKRXvV9sRgASzIu+mZbFwcnU7LzFiOtIIRG
dG1Jf8/ELrLZBxfZnHHoc+4wll2d0Xc3zOKuLSIzWMShPG5rJQBjagVHc5fEzrMP
Cbw6vM9Bprf0NZU/4rSbnBSpz0yhjJuVKnFx54okaH7IqOzQiZ6kEUSDNnAewvkk
P5Oo3TK5YFC8u3MqI1wzq8FoHaGLDxqUVPQCvq1Bkgat3gRZd5sXVLc7Sc7qlufo
q0tHRhm6u1OjegVQ0xUsuHNriiNQ8N5G4rjI0EqhLsTSMqRxG//eRdKC4k5aktto
ZQ5Iefa/OHLjce1JhPg7ZBIIMCvO1vkbTWGWuIUV85DzWjP5U+9YccTYLe4zm4ip
vCgIxSudNB02XlXr1NkYNg2/3q3pqgtczQFplYbN9v+TU9N+kJeFPArIF9AHTp94
PH/UKpeZzRc1jNDgwp4fNBHCnYw8P7vNOGlvajV0+5NlYmeOVc+KLq9i1HlWn0XV
gJl23QabMDWYO1EsG2NOSg9vuUWGyRqBkCsMcSv88MvJilkigLIe0yg6d6WsArkc
v8vQLKFMmFIUN57yjafjcm4r4QiL2hDs/ZFbEmLiA0GCIy7S7pUAMcr3ImDhpf0H
YC87K0zu4xXS4YP7GAtBme1rKIVviUSvNsMNKKhOy5/hlpK9ZiWpsWpvO9qucnUW
znNMjrOalGSjR+JK5cjDmBAadkDSlRycVPR+1wW53eaxRR9w0T3T1P2RuBhCf4Kw
64fOOuX2dQtrQYXCvIvBQH/2WcdcWP6a3no7PLVtb/uWFoxn8HY0sGYW/SH3HDbT
6GGubkchkMF16E6XA2FqrL2Ey8mg7F4vMe1YbSENFAZTlEKfW7YRqEeJNPXBhXY1
fEQIDtGPjvK7/w8hp81Qr9UT5syYz4pEEHykZ8LONHkb2xGVW2vhYb3Sy+ibCq0t
vFp8/34mP9Jju8Yt+4jUH7oPhFywb52rKVFzis5ipEgHBJ4tikS4ELZO7k4+z50P
dZK0G64jKvzoLTDqaILZEQmPsyg1u9QIIu3ppn5n8i3A+Aj2bkzgWQrrIyVuuHw7
fgRpm3XKAIRD/wwt0QpUWr7ZOHUKwRd+3MD9l5JLuK816bmzziKZuRG55+deXri1
Jb3+jeR1Ch7s8fRqbeszJoHUxLPBqAmvb76d6u7+7eJlKB2Jhpia8PvIZG2XZaNh
KZuwKNsr8votgkizvFlplNk0KJXzPxIFrYPH2dnszbHYA+rHXoK2wtQsdBuu+MNr
zYvXDpDzIVtt1mRLFVMyu8QZKH9uu7vXaJO/pnPtIq2y8Ipz3N/2cRB/QI2QB++J
vq8zduAqNsGoBIqdzkdBS/+4lcs9EcqYO+Ce7YSZ+Z1eQbQ0T3DH/axH1i7lbsYF
lDy3ZPeRXHbQotcw4s33TSLBKcK/LyypXd2X+KRbLpV0e7OSisWhb3jKHN0PFhvw
OFosLYkB2d5xomk/QuWg1sA3WXtIPsqtIpewNSm1xY/PQc8ar9XRsTwsf5GM+SSN
7zDcHhl5+BJHa6/0BF92j6MiaXMy/OwnnodSLEIW0ofcvpur45C/rQu1267kd2OI
4z2FoKZC7PsoW2fUSPxXSDeOvKhOwyuYXhvxIYSGDgyBVUIRHbCrQiRkTgrObtZr
wdnfGCepEnHAYV0arHXTIMWzYAqE4etEq1RtIS32tBx5AOMuENnm9GVxAJEgXfDl
lwCMCj+PgQqR8W8C9tLfhM3H7+cG4amxGoZAp1s+0SQBEpehwcB6+JNpSntJ7sOi
TQ7wrEoslxzSJyMGqZdtXV8lbAgxCf01LceiVo3wvdv0X/i1zTTPH4P74fummc/w
4GIpD6r8w2ncmQp+AE9VLOnRJpdlhf2QyTymYM0EEb5vpon6PHTKi3QjQYxGOu7Y
oNYv83mWh2w7bzjxxEnF2K5K6dJGnRXEAbGMGLH7W0PPO2uHHazuicfBw2Mmd4Jx
BrAeDV2X8OFEu0/6RwHP241akSR4QrG1xXvcJHaEPi8IV2TcuU3LMk6wi3pt+c6I
uzaXvMKreZ9GNjge2QR33kl8XMaEznNSwYMeq7zmsg+/y0yWsxRCGSWcGpbn0cHP
psiuAlTEIKcbkgJxQKkomdvOfWTMk9vJmbEufxR4If44j8vlkRplZNdH8qWsc/6m
UnHiU2odkMhXnut/QT2gAGJO6l/WNz9/yMbV5EB3USUHZVtd9VO5ROHTTkPw48iF
Kpg4WFKoklqxxdj5/f1GeWmXJrriESwNYY1F2FCJEC37eXNnCFhG7+KL49hQSwm2
cME9+7wWrzaa1lMktF05HSHqLpGMfg3mZK8HQOzuLTGJLQ0RStoJxlVgT19hYXCQ
L8N9iEyihJOtPIHmbSfc1B1xgF6vKmOMwZx1vWaNE274npsW7SfuWeME3cnkTq6p
/icJwE5DHu4jZ9sgASaDxydTkNAQCZM8Hz8+QnrqxTVX00MvdIUjLQjSR9lZfkZG
aCGEEbXJm18FLC1PAK8OSJIe9ZpQm3SBPHI0+W5LPIi2zLj9svtY7550zYpBksYf
MR0q7mgutf9pKKRKXWTgM0fCiohH16SDs3WuAuO0j2c8zLg5o/oZ3tIqPzoZf4tT
4rXSl9J4Wal2yHh2Zq4Vn+b2bBm5GKxSvDIBW90KuCDanLd794IHwoGXFLvt4tQJ
uoFzltTPCRpW4DiqoOHsspjo5CwNTy6Ptuwpttfqo5rnUpB/lwEVgszyYFmmQ7yV
dCLV4IIzoz92d9IeiVP4tdF1t7i8QCy7Q03Q4Ad/cmH0+8XIGTQhP0qm2bme1IRZ
eG+koFEz/XZdoHV5fhZcjLyBC8l2WfqlIOz32VzjVTQd9/U2Meyhu5eIhLAa0s6K
QrchrKxhR5wVaarXAdU+Q5xycwEhuIjfP6+Jhzc4wnyKlR3giAQspMmf42heUfWQ
WgJ+WjssirWUk2bbPASZmvf3LrwR6h5MDf0oCSJEhHBvYGWmRp7/UPtBpRDwxIDq
ijW5CSrqXZAOqkhA3JXckG+DA+OLsTYUyozcVTIRfxuBSdsPDs+CkNJ11NLdbO81
SmN6qwPk4I2h64txtD5Fn8+A9rPCmBkBqPNxj6KjVo9toOmbObyvFxUNIldKVNfb
8ocDl4RoA/rreq0DLZABJ1yYhmV8CQKq1embWgjK5TA9ItViAIox5pRKTw/V/20Q
P6hDQv08VUWX5QTMCTgfwbI/lZTSSwP5Z2ROwIv6JSSIOyVEWImRrjqxVXjq8Z7B
Yvn9rS0OwD3q1lRr6dqDuGve+wC/ks4RevdJBW4l1iZEHsm2uPsWxuPc5jZeFiV5
4MpOVBXpSDPCCG8lbgU/QEGa0spTNfL80KaEUijmdEzF496yIfXwQ6um+IrzfnRB
HZ8K+E2vJtpiKbqLJ1E2CWDSeQWiKMEGPdc+uiL4TFRPZdDklKsZIcSZbpUV6JgN
tIks/deOue5rRk52xF5HpY5erUfLVO5Z8E58K/WWN6OSw6s1QpNvaEu6iV4EySGS
BYAZKedKG5SNsJNWVwmje6PpArIjVMAdNI/pGKH1p1uwL17xLKIzyumk09ddQKt0
Yhh2NMbeudwQFFq6hY8nK/Jr4EljIQlE/EBTHbVTdt3IxQlvgVTKyod66zZXj1ry
tkC2vaoAmDUjXBNQxjEeJNUkQ1dTFOo25PLh4hj+MM6om+/MmAbc36F617UyWdce
xO0FspBOuOYa0dOp/Jx3UmSyytpcjo4EkTAfO9MHOQ3Ra1Vd6Au8qk5rAl+CbYMm
y5F76hFEX1ohCNr98l1fkh3pyBxQSxVn6fV36J5zrYI3eacbw+2mgrrMoWEiI6E7
Or4HXsSRHHQ/sPCGtY6PDUJSkpDTLWvQs9Sp9698P/YHDhsLs+txIKL3v3V3vyJK
ztyUfSi0rjQTMLrAPsisL8vYB0wEkYJl39dUQkXNMCz4v9GL171/CFx0VHS6WZsX
1mCRuljySMMoMxd+qnaYJRXn/O7ft84AqK0BshliYgmaygrJROE9avJLZnN1zezB
Tfe2aekRujTMz8LL6fijZmTiqCbUoiEL9j/CnF3/jI4YE/nT+dJGdl9iYh4k4KO1
BxUQ+8W2Y48aBH4SIY2VbzPRIGTAKOWsLM5QBbkt/OEB3kQZIdn7gJ76JFkcIm6R
I/qPrIY6k3He6U8E7+FCs/8g5pq5kUKmvZlPk87JneBvhTtXltqhJMhabDziRama
gPvL1UD8DY6iNUqQUq9th0hauD1fShAMoLrgYapNqSVFGDDQA6APMStx8G54505m
QJEOPnsEjKh2kUTQtRAIADyyOsf/baZOcxPTP0A1Xiw9ImzLzd3EQszRtwGTBs+l
FY7+aYipmguy4Dpw4MKBGKEMjrYmb25TB3V9Pqb/HZ3Oykm037J/2wQWD2+fgs6C
/4wePc8z038+x+wq7ZpL0yfiT6V2ffwJblgGApnm2Ce8efxxuGzMlpNB31BTuzEJ
npztROeFfrJzXEVA0Ldl30QruyCbeuNByfcSOh0SioOtFo1np2qy1uMbsNES06Lg
UMdftuQNYVuLl9kBXIQ7H12V5LLnahlaTiWGSD7fOplsgNYg/ScM9IzEoXkmS4zV
Sd1sMcMLKBOG8APM6ulMKqbSRHzNn1YS3lIQP8UJuXRHAARuc9Ng4cxHjGixNp7h
/9PYzeyoek/QP73MIf+39jQuewea+iNC4VQ+0X0ycdvuzojgGFw6oG+dfja8/CTg
vFKr4p45Z2V6ERmjkfaGE/I4PSAzobYhi/r06moJ6gGubfgA69IwNQ6fvq8VeFcv
y/Z5+uOtyDWt2ea4COfXaE2FKzu7PQnm+yX41qSyj/qoV+F++3H6xoiLcAaI15KN
IPsqSaji/epXnKqt5t20z0l8dvlobIxgNrqJV+17Xdj/5MY+Qq0BHZYorJ0f9R7B
Gd1X5W6cQfQ/7aAPkxlkB5ysruL/BKtAs2fe9zwa7WBM4JnL2/SPUsuGCyNkUfMp
AAqvNMd1gyWIGShGZllEU41icv0VFzRDpBjK8I+PnKHFxES/KGjGKCQBIz9MZEzj
KfHEuLP5+QHWpGPyTYonGEDeWfRiludo3w2W5S2mkblZTI6/wZ4aCLOhNNuYhkmi
1XXgJ10I6CMpBZjxe92DR+a5W7MISxRPlQOLH5+RQK35aLXE16uvmRn2q2nkQZ/I
hTKW404hm/xgPYf2XmpTB3CxNdaOPSTvyj/U+OKAj+tj4UlFLS1yfc/jFV+zxD2p
L0SGU5qtnWgOH3TU76SGuOLaAwAi2AvymNX8bEVIZCuRj1LZrnUx9vCYo4EaX5AX
1BGSgUwwH/pqa+y/jP5oePTfXRkgTDOIEGrKz2QhLhynDumAXxORm+rMT9Img2Dj
rOOuauOS87dHVQR4vVwq17G4smYAqRrevCBc+aZ5TectNCmVYmpfWo8ZVmhozFC4
WbxAIuFzitZmMCvX+wwREHJoWWjFdNc/Uwnoc7L8vHAD+rhdnAoSYVvxVRwgKBea
y5cVUGhnTE4SRk7BNU3HVHLsX/gk/d4PM0dBuCSrfvAl/Vf5EzZHSA5lOGux6KMf
dHLvrSMFpyfKsA28n6kcvCCOkfwJ4Z1pUtKANxkIKFcN3TIsXHvlFItxdHqQBZcz
MzoqjPezsEyfWLRHbkfiRkdv8KkPo8F1MUcvn75pUi7OoDCIa3cHnzlyTZMw1Y9O
BbcqRiYMVvE+AJRZgr3xL6Dz/ZUf3oouLpq/dYzb7HqmNRShXh7R+7tKXtxFbzaH
xblEjDMAOXk9fFnqHFx8uYnvJqfrK5JlvutfHzfIogrdAAPRExIzkcWXgWav8mmK
Cfct77XUYeI5oMcriDEjEsClf1f+cZioSjxu/OoQkcmg0+0ihNPmWrMBjbz7Ky4q
3yN9vJzfaX1xJbdCv5lBDARrSEzT5nmeIxINO0mjHMDQAxLqLuDmBPi1SmzI6OqD
aciYyf/AIRkwBRUb90usJ8FEiErQ0LArTJa10kJFu6ehLNQbdYlsTxHOgGieeK06
/Y28dzm8Qlc7cLDA40VImfCkPcDpAkkxa9hfe46K48pm2Y/lNtFVsL+KNE/jRuUl
RWN6bheljO9kcqbOK0yOuDyCsqDHy8E6IOHCCGy8u+QmdpuFCOKnr9FxOwJIBwem
jBamsWYajuVR5edw8jTpgi9VcFtNsGWRIplQLFJGcgFyc6M8FdaJDZqdxrOXX0GH
zcnn3RU2IVyzT358MRQLfSBFFSyoEBlKf/N65brSG6VWOSTDyt7SqS7BYw7jyVr9
BSfsd04t9fFaxbZzyHh4Ahqbx6W/CTOB9NtsZx2tl/j886DrRQSb1qV1CEvPyvtj
TMNUQj7Dv6sBGVSPhbMByUIbZYjD8M+sgpgFs0/KlWetf/kmH1y/rejoNl5xw2gF
IpkxoBP2S1KjnCrqkDrj+8R//jNm5+TZESppapFMeQb68O1PfDZJEnAQg7Nr6gVk
j2MRYuFWV4eLqWfgKJmojDSWspxkjHn8s0bdKbPlXWMZXejyNvIYfRsZxv6Lg0Im
6NKigWgjiO6eQaeR3TWrr1IWM4iAEXcDiSwiZchhGtisoZGuKpym2Z40A5pGep0o
4WKboKE9VILmBsWW5kZMkKnam2+WvvGt+evCHm1x7pSh/0V8ZqhBo9pQ0BZPyK1Q
ZLjYLkybg832YnEqdiuufsvb6HzQ2bULzugPgqQoguisGDk5lylu8RMDXRObIZnK
3tIcsyTrbCydWAFjXtx6jAHeDkCD0RgSN9FRUyzjdBzt7XzwfwDqs1YZz1yvIg8X
VIfuiirIThfDpnQnpv2+hhSBOy/vjva7J/stLkZvK+JCmCflCYSf6wJaeUoJSg7r
UcmlWb5/xTvQUCiWeT1RGxrVxt7lBqG0xLRkgBLenQSTcTOJv3fTlwoVYpx4SFop
551fIztSi9QfsThYJJAXKOR6LoSVouqdHLINtRezImKzd2nBVf5FcaDQNfrPReRq
KillDmmkRVgB4sGIs2Hr2NigZpq089FDbfdzMWOGat6yEg1wy69hy4bpA3pTYawV
AFWhMRypjppPC4rKbgK81lMNHBuP8VqmXfbWpM4Pxbd2QI7UbZC4Z1uKthEq4jxb
xojJBYVSNACiYQFL/6BvEfBC3wPqgN/us0fek9u1Rdpx3OVtGU62fL2tOLt/9JsV
ETjR6LIy+6q14Sp6z2gs51Xr92u8l22xo3rVijk+dAZAtddL3dprgAvRIxUeY+K8
jygwQ9+6wCX8qR3BFOTEYMPJfNxX8cwgAP9fOxlCY2bHO3/lMGHfit+nHBjCqqFD
SnG9e0OiwdGeb2SSSWXEcNK4/zkSoQYjjEMKgK080UYc3mhtTGjs3V3YIAQ7nCNC
6MjmNJzeds+iTR7kZHIrV5uTrE3qthW8t4wa742VEpFlKVYW3yL15JhCjkMHx6YX
Y3eYFkvb28Z+ofsBUokvC+OEbCVxHDljQolvXgOajg+eAQpYjZ5GgJNcJPSxtj0O
ZGwB7PWp9i7jZQhQ6qTEgg6hfS2h6dpfs6D1U75UeOlO1URlyb8HVYLqPde6gUfI
BucWP60XJrJ4jfYSjB/KYh7fMLvng1wfM780TCqpkim9yCv9mBtl6/xQDTKj4dhX
oULfgpihYJPenDNWz8XJxkpsDwVd6VFhPc5lPGTlw4BwHCDHrTzsbClBKcrPAt3e
03O8IpP/clRCMsoQvtQJFN/qMWKDasCDoB31NoHPQaQPZaJUhZC7Wy3bS4rm4kVY
IcL3kYm2/xVNblMgqfRfWL81/HiWY9tYRNyVDaHQ4se6qgmRP/sxgAWQ1JsWXMuB
GPh+fFFO3irGV68Uz45Ip0OC8g2g1MoxQIVc30+ON/4/S7Kxk1aEpkU+ZUtgC7rN
jbCDFratyulfkJKUBPwlakmM+JzQM8NmdOsrAtRL9Ep5GtoQ78PucavyRw6BIGPU
fYhq80YEhqIpXhSwHY3Ljt4RXipC02n0rkqmZW17QHTRMkHbDLovyNbC7+7iMWzu
Yl4N2X9V8HeP+8HiV9kFMZcmLVZRj7SFrvKzlCJTunAE59WLTIwoqgyYJpzu0XMa
o6UOiqly9ycXn07sAsaJ8spNk+nyXZTVVacQ9XBmqtDExUAKoCWd8x5feUOxTSzg
rxohMLKfJT/vWBxqWA1O8cN6XkROLbb84u02HTHCLURxE8fHb3hJwQIDHX+1uH78
BQm2kQ1Vst2CcdaDKkE4de0jIADp0pDQP3rqqlhYB4eOw5/SBPH53coA8sc0jXx0
RUNHIn5jCu7NAO5ZM+FF/Uo9Vfi4dtShZv2ZtZkpLSsH+6YmqmHU9zZldT3aSkUN
lipVu4z2yaOEgelY1vUqub0Wq6T6zqlU7DmoZ84W+1kg4fyh2ngLgvpUU8vrpH2B
jk6FrVB0AWVMBOwfPfckMX3WbgR6AIvZoymzNy/RZZ32ntQD+b5zU0Z3WpD4AD6Z
GXFetZmXpAqWGLe3Q1WkzKKd2NVzZpI7Pp55eYHMsm9GOeYoazBuYcn1oFJm/AZP
CloCkHlXq7Aba16cKnJZsLVmXwdz/esO1mlw8dA2umCp66fr/T19AvQdeHwD25sM
auAm9XJyU/LroQcv1YBLDwDxT2rfluNT/WMOXDfx/PUVz79cwW4TRS80BySGyNI/
tdvMgFFDU/JLJD+NI7y6hiCxVPEbdNAb04bUR9F9pjH3megb5W6TdUxxbOVvtUS4
8HaPFyaDdtHWkZj+Rg4yZ00X+v9eQ6HP9Pm9CXQOT6FxV22JkdY8eAaUALGrj3gL
AzZWneiokJrZpjhqjpbm+0sx4lZS7hnAhFzDmT8pCJZZ59T6hAqD4rW9wetUR7fe
dyVQCrwUMuXlmeKNP95pIXAMrXBG72vTCADU6mPv4ItJ4UiAObemqMBljKxNbEHf
8Kj4ZszrTkVuOWdI8HMWneq+ZjutinW6Kq+AC+x37SYI83hclnC7P5czn6SXhSyE
zscM13+f12+YJykZmaLuME15qJQwL/E2SFudFa/IDzYfre0ff8EHdHYBCJiW7V2A
BOmsTpRKDQs7YLzSYFKRFvCihncvj5DOGQGjmtLYZhA2tIOqF+fF8D/lbCBLmpro
Z5YJwQ4GtvaQWYDDz1BBkmH6j4jbAX0pdDI5DZZVn5TClUpP8P/9qPJhPR74H6G7
MPlzHNSza77dJKuoZhagT3KzNEo1E9fqkk3GPgd4Uo9aWja4iBZYExPsIlHQEvqh
hFkpo8igN51gllWASfc5LN2GotfvfgKk7rzEtP1e1IqpNEskIrWa1MrpFagNYL0P
h72ZNQrqm/4CWJmCb5AuoIFWXDYPHQJZ9cr/5vOBrhq1y0Wkwl5vU2P1hIK8+mK6
Ghv4P1XrVo+TBPZGpO0HPaEqOA40YEBXfkYTcxFrcZfVpN49Dy5bVUOyoudQTQmk
X309iAS8xi72PAddTsLKtQC8qvrtbdKwIJ3YzLdZ3lIvNCwu8qanvC7Iy5HyDZNj
6Rbao91tI3a3PV3yhBpqSs0dE/YbnJyduurV0a1ZnU7lWHZC84aO3JXfWe51aLL4
WMAbDxoPqiIhHIhds06ZHjCmS5lmWMfeP1ZYm2kyj6zEVh47V/Zm2kKfCEj8tc+f
vqdf4X4K2G/LLz05ytVyBoee5wNlZfwp3xTlAHKyfSG4jSaD/ePIramI3p4agNqp
MtFCQeBMXOSuiJh67NtPx6HjewW7n/hOtGrCt9C9j982JD1Wv9PS2y+OkmpmRGMs
4w/zRSdDBSnAaA1ay4U82D1CBeBV6yKPCZA2faUelSYGVQFgBTRK05GDERa72XpW
EM/mCy2ziGxac2jFgPreqGC/MwYy99Z+KGlMTkf7Y50HjBcyI2gAz+GU0yRa3n2m
9JBBZCa4r3o/K2BUPZ77i6CbtvUS3dhOwNtRxEL6dmQSuneenTTcPDCBP59L0fQx
xCQD2egf5w7d8ZXwiM24eLC2BI5vzHj9dOMNqriXzAOEfUc3f6mitwOAHrm7C/RH
ccng+tFesi+MMkMiFgOYnLkQpw48Rf5YsSJanFHYXDRRDFzReJyR7wEXyRmoICfV
XiblPCcgx859KipI0aNHXVM4tbtX2EswdP7xdGHWooittKKNOe0Va/9gdsXthkx/
p7CYh6iPLtXYq5byMXEjX7Ray1qGEk5f1Sx4UBZJI101xQSXhEpd+RPQxAx5N69I
z2KPghvy9b1n9vFctMpYDCmY+ZhcwblSqLyonHoeYpMm4VH3Ve9R1eTm1OFJW86t
uIprhaIut37wmLpphEzniRYmbMY4SN/+nJx7t5ybrLUoegTmPV503V/d9nWnCkf7
UCeG+7a2jdhJIk+hcZOvwAId4wlsXAZ0Kvb7qsvodp8w1tuNTqgV7Z/QYSPFjADl
BYlT2GfiOHF+Qw/aFKNnAgjlJhNqj6kbcW9eSw6ebm2dF2rUQ5c9ynaI6mwQJd+I
GBiHRZrORDbbabuCB77HUaMWF1oJiymmvrZIiYLoicI0Cwv61rB8ld2zmfNLczsA
OaLne1fpsRi56R/iFFV0QB8RU3yY6Uqw+TvN1F/LfZyAOpafFf+S9cRbBTanVZyF
fCGWQVs8xPNOLdVts/Nhbj85+lK9uXLK1c/HNrlwcITA4kvxJfA1x6wnswmZ9iLi
X1llxjfGMWKwJT1krjvctYHwgnSwT1nlkS9ehB+e1vPYVzUqIqPOkRxWWjyyo7U6
/guSXyroYOCVpnQBvWxM2OjVGak27nc5SwoaUHQceMGP785QeYIuJ4A7TderzdsJ
NqkCwTbbpEUUynDJC973dAbAaFVeh5PL9py02Lgv0ZG06CFUhVqSwXP9M1rxH5vK
e8/n4kqm7gYhyu4E/GmGZSYj/8erzPhMBimOU7o7u21T8OP4F6Lon8S0HF+xHm66
2OjRxYKK5ATJr50HIWv2WS9B88G8+3tmLX/RYRAaIGpqJCDwN9uksVyOVGSpmX0W
IKPwd8xdxqIEHq/HazEnwbhZwKVrif0ZjBP9ny3pQjgeNXOghPzk9u7gMlMOXkkL
Htyel04pEXBpea9BsnG5o0ijBWKN2bT/dMiR7zYpW1C/CPaQn99ZMFdrz/YDbPBv
xyA04ncwURGml79wl9KfhDz0rpkkydR4CCH0bJHxBHUq/g5mnSskmIQ3pSo2PipU
sACTV/S3VEJpkkkmZXvUkaZPDrqFuhQUs6eztC/y3PSM6iSEt0/CJo5YT3ABNUhY
jifOv5cLhUZItA7YdvnONDMoSR5ziVYsPgaCUTqmbPALSya/9jpQVyGxSZTdO5/3
P6xorOHD2VAaX6R3boeSjQDmwJnZFzwULs6hRIu7VFj+UL57aQWZxQ2wobqLUd5q
ZYGbTPU3mnzRSd+7Hl8IaLpHmhgkSd4FhkzIwMRWtnb22Yharz4nbuJa8xgY82Qs
iZN6O9RJkXUsrS08ZKj77aJVWZCejnMrGGS5bTRzKB42HDm8ePUnRek4q5Xe+MOT
RWPot0KgQssOWgnuiXD2DgJ719vfVX34MXOIxOujSwscKzdbOVX21+9evY0mdWWg
PE7MxUJds9Km1gb1a99+y8s1EuhXUzU3PZhX4MlvtMUPKU98dvS8xlvW4KNykzqj
AMAAGoZXEz5De9pzk0uwXBke5Ge2fGYr0BgPiCIsZ6qA7qa2mWt+d9DACSuBAq7O
nh2eVGgGYJE77OGGMXbt0GWtEYSh2fIdsBtESzlNVH3kL6e5YxGmd0uFVIGgZ3/C
OAkfq7sUVvM8i+PIEBTPmTlf1/9HniVdDKK7xbEfRG274z32N4ng8egayPYI5l58
+zldUbKBbF/W8uKu+Y2Z6pJHv/+C6FtE9noJpIE+lAS0tnzlhN9ZPeGTrT9Cy+sQ
xJ1WwkruvUuAXMJWhshVdEN1rsHEHEIv+QsS3ZQI8SjsuceM1RFWuxwKQ+3hxU0U
qfHGNg3/KzBJORIMQz5xduXIX+J/gfeu5oIKiiJ1Z9kAwThMhX2twIChxjxwJwvE
BZtotMDyVFvRMASWZYGAgZm3j80aeodDYr2fz/SWLq5oENbPWzfUgltFZX5BSH4b
jePWzxBaZfiB3H7oNBeB06jP9gz5dq5yp3q1Wj+W71r23EtxiKO34dLLGqB9qsm9
AQ89fUdE61sC+jf8dvtkDjshk93pZkPB5HNJQkob+npc7r5C9CN6RTjSCE7lkZwm
/CARD4M8LVNqWHCEerkShuDSmsfx1nx3MGGVHACoycIaYaKYj+5lZUiJUF0LenRS
92NVL8fR6C3OaQTTd05YDPPASy01BS3vYIHGRb+2/oq2YoYaSI3WuZy7i1kJIMvM
wp27eqMhVYuUhZVKNgZK5Bcs9YBKgRnBk5toDFiW+Y5tTJQh8o0dtP6YC+iciw0Z
fnwjxhGJAjadL8D22fuenoDmCEgaAIOGbXwi8shH+ylia+KGeFz3fKzhdI2n4I+q
ZYmv6cUIRSvLE6BOjY0H5WZJ9ofhXIogModJdY1jJxoS025TPnSclrhcTu0f4oGg
YUDEXmjsAcBGBYuQW0ePGLVczlCsV61HmXOhG7xZXWH/8ALWo9bHJjIJ2SYQXpy6
37h8eDHeicAkpPaE/ihEA8v5ISGTAev8drHpt0MHOqgBHjB0UemEwAYywMHZyNXh
nz0yaLUSaS+YaQoZlpfJyUgOyoAAi5qKstOoRn4YxMPV/1Kvj7RcTADVfV9wqZNo
UtirCCaK+bjTjafVZYrQ5Qy1sUg15VeS5d5FakCL95UHTF4Pu46LElK6ljm6/AzJ
mniiLUvhSqXNG+dN/OSJvRwL7inEovDYrqd9FmLUApB91kTXE779Hg0HBv35z7re
6mK0gSKcBxQyqdto5JECLzXLitTXp9TJpH5dMG4bLc8E3NlYKZw2YkIStOCBGbpC
4bWYhPOWGxSs5iQLSYob+/Ne8X41OUsr1Kb8raq1BRzWuIC2jnWecxCqCvwmm9Ea
xAn1iUNYnUgl74MRpcUNa38z2UDu8zWkzs8ALG2jx5W1x0py3Vf8aEx+W1MlKiIM
bgCsYIBvlgSgwwHB/9g3xFWSiB3mA6EoGFfMvffqIuK6Dl6ChLnM2THfrPMnfRv8
VSU/2I7WzO3yiCH0nc3ivmO5wi9gsRqzgedlwC58AFa+r026NAyoNGtMeDKGMbBx
2ZWGycjqAKx+zwRLos6bOdxLVoEQL4frHBNXZRmGBXTGQRCA/fYgS1+vVRPSjilK
iMPGlL3NvjIuZJyT+kKYhw2sl20YeqcjtgbEglteZqqN6ICqYNvEW0k76IvTlv/D
i25ezHXjAG7FKKTiP2B30NOuVhsmLbCK9C26UhEZ086+v7XzH9W/CdA2k3IGR9eu
wgM9dthki69c6ngKC0wloiQL3AlyReFypFHfKmgZhQPjElPOS0rTkoxenVyLhuiV
UYp0FyVX8qyWRJgqd2w3MdyPxe+ETM1DghixIjGFNYSeSXvZnclhCKPD7GpVJ/hh
YxzQn2XqbdzD0hICt/M3ODN33ZuudoBoX+aXJmcr/6+ltPycyvjp9WQvnIcIEIgi
84aYyL1zJCiSFTHvwwHpFWOhybSzgSEXCEvLFGWrI2GOUvie83ZMm6H12751zgVx
+0lQu+ccda47jvvuLd252afyjuBo9FYVpjTX0TB7TLEoQtL4J3W/kt4httTu5CN/
2NW9dfn8NrBGIWnrzpfzf2vJqlbvvFCKbR5aRhg7LtgPQkuLblkiZSgqL+Ony5Vv
RDqM700lV8recinJsfUIt8md+N9U2BhrQv9hCXHvVCTioyfKEfVnFobXkNEyReeN
g3Ph0peyltWHrwm+6qEjwAplLm/koAObQ3R76212/DbmQ2iQMhyKFcy0nqPnWTqD
q9DKQtEzOgVts+jydASS0P6dR35pIxqghrF+s2aZbhZBXbwIy2V6SFMLw6nsGKkr
ySjo89QzZf6kzDV0vi+c8hUXht6E6aiTmCf6fYrxnX/gieY2RgtlTNwvpeBAbtdL
Nu+4fj4fiL7VfhzXxnsklRzDkP7KBWAGLLY08kEE+AhFVvRDGgJ/BsYfHGLiDDTO
6cI5qEDRsau8XhGPgwr+kzbkX448LcR+fR552m6rElRMctEzgORkKyWecdJA9w1t
Mm22IL/SMas3rX9p7cRFDyslzfmF000qOPhew3ZpwQ4iIXfwxDTAi9K85X6Vr2Ia
mpv2Zt8RJwqSE5mtFX+jZUezLPXKuCYpEAo05f8SCGC1qw85GM3YMQfjYgR8Z/CX
RjETflHIdWKi3CayY4fQBDQevhRm7M41Tyxb81uQ8B+geGCD+54L9wiRkNlax/O5
bZRo8wiw7hXFnZmQcpdYfzF2s6vExLqTX4B0VUmsUKnx8E2O0cMpHe/LJZRD3SFA
0JoVnyKm89ODBRJbF99c0Xz9OHHviCutaaDzhW7wEAwjv1ULkAAKDGehVXtWvDRM
HZICZ4BpUgNzOAB4NaQuf6ajsBv31EcB9s+cOS7X1/d4NvJu/JvgVMZoCdWNeC1/
2Jw3755+ivsXNS0ysxRT4EUCk3WqmvsvPgVMDTi0ZDHTO5XEFEAdTCcbdvi+x4zW
gpspw1NVo7IYUyHbiN4zP2W7ROC+hoibbUQmRozj3/dONYkIDNqKktpbi0Lm4sQO
9D7QhM93FwIa2Lw/Fkrlw2EPMjgKvLDP2mEf99HHKDm04E/kdL7EhP8SAN5Fpxjf
c/F9pSDzREywNiWZpDWuw5i1AAdAEdAT4XeFznVcNvcY8sW0J1p34iLmtDDLMbur
l1s/+YueplJ4nAwJJCcBQPLdWtIEZg8mQzIcGdB11x4HoiAcyMDQWp7Gw+7wAnUa
2jsMcJBeOUiTcI/kdHsJz905yYMrh+CzF7m+FJQj3nyEbZPgPFnXp8EjHaq4+YWN
+YYo4WZhdH6jAtJzW7Wm0p1RMkOYOgBYt+8vC+Ho/af5W29BfLo+mC5fAyVMZ2+W
SekrGtmxcXUXGlErRs5EL0M7ER0+fb+8O14UoHZQvWbElapUXmFi/LkP1auqKyEY
t8nbQ781X6EaMgljJYR1/zLTIeVYK6ovZiwg+SUsfAJXx0vWgNQppgXFlZakMr6e
+sYujVvzR3ODYJzAQx634yTjcZO5P9r5ro/JIDn6vdyv9Gohsl01Bbt9RhCFCne+
UOsqTuG3/51Tkq2l/bNfxs5jeIKjcOSUspUQ0Y398rCs6aRw9NI/5p0YLdOyvU8u
EBl8+KWWMRXfCFDZGCogJtAfQBU2ckLKdUGaNRvYw7TNS9t96LSF9QS34bkqxn6/
dOYOV+soKaqNxQXSpcxROHVBExtn3EXRXbZrsaOR9hb/iu/3lCNA7uBfrwsCzX5V
3GlZY6im1Dpqtm4GGz2LIm639m6lJRCpI/OyHj2pWLsxozhxYxvAelVP3/2NmNmN
oYawGGvsBgm1tYt0QMqfyMFJOLMqahb68zwZuH+31ren9CcUWGEoBIeOKjrLLpGt
7ZDFhYIFY9aOhBM9LKpNdFzBn1qAykRDwXlVHbdoz2EC60MSd7SnOQ5QAk4mYmD4
quNh6NI4/o8IOjNOWt3FZg7I/KeuyH7SzjQi+qmPHBLVtpuC7JhoStlfBk9yHOYO
B+10TOGy5Z3zkB42SRgf6aNz2rhXSiSZlQ1B3Jbg1oZb+ba65icMBYPKOPbBMy34
TdTnfvm9m2lzmenFFyhI0hFrxeMd8hSHjjEmDYyUtTQH0oniWNSc3HNtjwdt0X9P
u0evgvTKhqtSQpWulhcPHWppkx/4ONcXWXdLk7YjD44GN8zhQwIYEuGdGJBRbmO9
3fdin1BjddClgTK18ZfOA+ddhWPL2C6BHXuSHlU1e8JoUECIjIG7siIhT0rz8wCN
gRMWdRfuNQgOZ8yQiWpF3m1fFk6E7voBVV7B4lHKLqlssJv7Es5xAwHM4ELrUBgf
wLJyVKKU9/6+MvWozqeU/RV3HgqYIoesenIrTjFTxP1mvkxqMGROYVDJogEom/VV
b4+fGZBWHgBUgYkr8O2riA0Hw3DxyUA+FdV/zAHEXO1bxPGTdoalNpvBsflXSjvD
V2eBVQoc5t4dn/eUyU/JiFyJVTGWMR7Js5oKC6t+3fjvJQxLyFg2ViP1VUdXObO4
5AuSghHfB+RItwXkhkojD+mckHWFJ/9Yxct2gKdPQDvC+TWvGSFGWZ1piYOJgKQP
42atV0uu50p+G/2HMkxKKU7HCxi9qQTE+DP7d8O20uopZHxFpPFtHOP88vqhNMEx
EP3DDeMsLGOUxIYb7ny1gbxuiqmFesKVGh2DhnVhE/eY5FzdjsyIeQ9ePjh9FDxU
zGJPsaDQq2wL+xRerauGgXZUI778K8mFGvUbUtSA3lBv8XTT5VDl6rVRlh2ebPf6
4MOriybC/6bzYPwzskq43ONxvCytzBv1qIjPW5Og2vxtF1Uk1cUjvH9AQ0cQkNd5
Ik9o4b7AK4TA9MMUS93wu4HD4T0Qx1XzWJ5p8nTbw9iamcGVjNaSqYVZJkdiErPs
aR6Fb8TmUMB30QhRityChpiE6djtpiaVG290GEpFunC0M3clthzjU11RNrnrKzL4
8fcDjxhnhkDJefaKkXvBg6h9UFdSKaC1Rg630/2MdS/GT2HvB8RDq4tPVIew83Ew
oLamIqHVtCxkNAJLRqM6BwNdbDm9UYDzoZbEdVuxTarzLcMsTHrmP+lEzoitm5kA
mLsS3PtANLnfhKRID2k8zZ5lJYXabpSwVY03h6G+XmUgO/lreAnLuWRnEevAbxVI
bU/xJzVZs1BDG6CBU0ToySfwTCu3V3PSfJX4MS475dqRNLn+dD0vrkjme/WrPjhg
fn+CWMk84LZ0TVJIc3z06iDyvaS2w6nlPEWDvQ/Z6UR71C9haNIHb2roKkiJJEKn
L60j/wb1qfRdPbcK48Cv1Ro9E+WigfuoEjDDcKttXihAX4+OUEiwyrBSDTDyDnTv
85jDszykdfA5qAgNX/8R9zf5foNbeuFFACULqlv7t0Z48IF1UUzQeMDPoHmMblo6
2sTo0yw5HZBMnTwKM47YCIPE0Dpku3bcNAYpD55uxvMd48Uj/1Hr7K6ly2X6yDJc
FKnyzKpdsz0tNXzN+jORvluP9vJ1J/sCj0UIFx5G2XGxZLywsZCUaP0CnnzbkvJE
7VrPrK3WK75lctQCoZX0i7fxpfxPdp9kxYjpLYKcd1zCdi1isZqI3Shh8Qtjp2+b
vJkEbypZ4q7X2M5sU5QOahTS8FKSvIk0TCSWq0sP/DEIHjGigS8dZ8t3VLyN8mQn
xQP5mwNmMXO4YakEytDTNGYC0qdogue53Ld6YSRP5yfZqFLSSJQMN0yHLnCyR6Yl
tnlpjW0sXziXs8OuxI3j4gtegmJQzaxvRuaHtGq68jsjjQnJ2gA4kfbiVj9UGXys
1Os/a6SKPDV/lRgjni8fCUVFoSeUiFvwTOiCmlxJ8Lbf02IM8oEdT9cfKxSHa9Hy
GFCsQfeyrdF74Se0jEtjEMCiso7z78ylS2QHAQbUng1M0py6V7XEXCbxwJ7ug0oj
1uI3WMuVNerhx6zdB/M7cI00RGMfGBUQ2A4KHPEjkl53ltiw2bkJ5OEtzaPnCgIX
Tps7xiwWaPYAUNr65vDwdE12z5DpDglC+zS8Ak/+baiLPgKH2zUzXGHuAG2k6q4f
MZf4WV6uIJTCKojbXlZCbO8j0oq9aKp7y9gm1Vx+xRMoMvP+CMATaquwMHeCUuG0
WOtjn3IeSiJirJWfkwirpIBkjn30tFXvb+T6cojbsfkDLcSMi/QtDgCszipiu8Cd
6eI2e3yKa1qDgmZM+WQL62hwY/CIIS0+pIhNErNeM1QDyenwN8bgancDjQqSzbBO
kaaTj2sUycmZj9DJBnpLaYpN6nj3GH71mPXPPTakv/SZdJc5JVkyXdEtrD6l8cO0
Ri2XSDsDM00FzvQ0i/OghTBB4gSyiD3dwdcEaxNprBIUJjAk604CgoE2IgX6yh+D
UuG4GsksmPihdzitORZWBjAkCRoKQwcB15yGgoWuWuqowh5im4sv6EvoHIeJldmU
5wmQVeU0lnIkBm56u7qVwaTV/F6lHsYoVXNMmQ+Qn7nyBd5Bd4S6EWjL3vfsJRkP
U3LOnqKiRBvgppmSJVDZIixcc4GYbM4VCRoIjpGYazrvUywoQiiCUFI4DWXpTtgQ
Te1ve8CaVZUNj13XQfjVZwCDanX72nbCe/eLHNJmFTXCzHxInYyFrIqx44ps5VNm
q0MTpNhRYpcGOSoGibhnBDdQUh+6YKIUTUOGpaAZMGVsr5Ane420+8udKR58rYIi
ulg2HMk5aJp0lblGkVso9klC/UvPsyR3tCm29E2+x6fD3QwMQsF6e6gQswsIPI7E
0S7gwAKvDinpMqefsFJ6nyjlo8E4vYen6py8KKzqQtRIXBDprzL7F0SNqd4SwZlN
kEuhmqRsR188565YbN3Br+GX3NMbqF18dqr4NG226FQfxm45pDL+xOFUNI9cJDdg
Zk1Nv0aY/7/rhI8Fx5qV7NsxKeyBGNHDmhdOCrnomQjvZ9XBu9EnT6zezxGZ4Tz1
0lFk4uue3A6QKdelcjVCUxoL59zZT3aCHlgHlgk0OJvBU0m5Yc5ObcFD6SFHkmgg
wkFzeOHL8YCjw1DHIk7G4z43aGSIDKoYf1fretSpvlOwgOJO2oS+XlygjJZ4X1pi
ecX/YS1lolnQJDBlQdS8bq24kpL3FIXTwmkfBP/Shm46Y9w0JL/gbCnOFj3qN8N+
2o0yMaDueum99PHtwA6J3qElujuHXIOs64fRDLDBHjTvEvtxnQ0Y7bFhBxivGGT9
PovvQ+LfSGMVZGO+PQ+YvSc8AMnm+cvdQUhAEweDLbckpmOVnRPoZc+v/ussk+sk
8b//sIMqx+0R1WTkWP2AzZnfFOCyKbgn8JRLI7uSNlCvWHWunp0k7ZMnXUfNbLB8
N+b+xAxuD3T75jSnQNILHdKIlwnIoaHRctSlpmK+MBaSsLx9FwW0vwnIilgxBeTG
lAmMj92Owvb5RfEYb9Wlre+EMUaUcC4OE4Znxqk8tPXoqPoc5c6QN/f448LLcvjO
wh2H/DegMT7hqSCJWwU7hsaazMDHVvOC9GY/a+gguX1bQD8bRVOFibboJc8JGakZ
KoaNyXh38k6l8fa5fgjJTyYkInJT5u6N/VBr8r/2Jr0OckoheZxbJR2iZnalx3LC
Zd8z09lLv4XLEBx6/tyW4/0nC4y/Zuay1GctsIGU1220uG6RN/q+0hwWbBmMYFoS
mpZYG7h8qfMjGUTnOUjNPSoyO/fLVr3Z3ttSG4BS3vWbYrKwcCDrHVhbxoFoUTXG
CbC67SCMNgEojVcFBlWLwukVzavY3i0laMAOqXO27wZRF2GKxurinB8/Jpook300
//zUsfxOfvKfS82b/7nyhD6qIDBQA1z0NQSyZkjFSCBSldnXM0dcqFhv7+2IUGIA
s0fpGQMRIJp6/RXRsFUaGuZRq74WX3FTRgU/UptfpeC2cUJ+s6o/crBiWKerzZUB
mC/WvgC5X1/4ca8zq0beq7gBS7MxdsaMEEI4YKgs7jTexQeZVudPYIBqQXwLUqo5
51UoCuBY2ZVOqg4SMG17wIndiBco46mKyrnHnsgKEz3FSo26qdjG02PWy5tWGqPN
JfxgTWymO4cS1AHpNBKcGp4kvvyVC2BgidAfG77ni10NK6C7iKMGh/h0T5g0I+KP
JZ5MQmLTydlbqEs+lnsNJX5FBBfoSPUI8cGrKIe5ztIWE/FSWgYww4ENQsOw8shZ
dgpGODTZUaBh3v7B5biw190tmDHCRVN1gy11I+uRUwmTcc5NS/Nlno2pOqdIqwu2
dB1H02EI3JTkpOyEKxbeOJaUiENn3FUopysdUhZK0T65XZMDVtZ4CAM2cCPTDOKh
RTk6W0Oqwj5GdwWhvMM5dgmFU/hsXXHcihvhm5L0kHKSSYRgkW5F5TJ1TIGTyyM0
DFovURimCcmHUvKg/FXnK+wfF8imGhTZPQrjxCTv0RybfVYFFHrDve9oqkLklvZD
LKDDA6fKVLbW3CKKRPnGi1Kd1KdBKZQwHYm1bM+epaWt/2T8n5ArgUF3LE25EYPo
6bsPU3FsxI2xrGv1Oie9R86IYbQuHspi9UQK8UoNTjGlM5bSplMgHLIzMaeEOBJq
FO5dmBkyR1BRu8Arfhz0EVf+3kDszVjfodQHbFXNNMtQ0zw2yyyMlzutnHlR76LL
qRjH6FzjXMXi4sd81hYxs6uliY2lq16IKzKhwsw39TdJtpkSJ5O7qqyKpH6RAksd
va99fIC/FJYmjdU5ihmga33veKw9Xtkz29pM0+jfAtDctEL9TP7twAO2hMNt5p8K
jwL2qNrbtoT/CWpN0ISy7F6m8ORzDZRCDGI3Al2sCYvddAY/5AHciIG/VQNE0/+C
aPTsSwN3xI0USu2qvXOEm/gsBwjffKRUa0FOiJ24HDQznPStupBU1j1XjFzsAq2b
3ukU/x9+sDEzICD1ihBJVdW7YIkhOp7X3mkAf3kzMipXKwqAQBtsZ3m2mgzmkjQo
VALDMu7I7OGttF56YTsBOW0LtwUKDATMv4LcNSalhFoM//EIEjjkxXZqTOGO3DFY
pmBLm9HrB8AdyiX9QA0E8XBLmC34qv5DXrz6L1PLSU/CpFIe+HohkXRf2lGtOS/s
2eGflMjOGWQTurSyNeQIDggVKP9b8LD8bXUkYXAfRTIq++F4um1REf3L9oQdzFg7
QcJS/8vRV9DXCMlxxyUCn7h6NFL8na8UK/a3P8FzQifJEVMQeKkHh+j452bEZr31
0EeX23rmqPTLq6XgIF8965Q/W7hZEzcg9dfkNbuV9egO3EplA6IK4jCkcF89lhcW
tY9IaeNZnDUKLU4Sy/yvUfcKcy3cAJiFqLSX4qxGe1/FgVx8326KDHAFHE4rduRJ
9pJq9g1iNd3hUnBLN4CB56LCyFSuvQycHV4+e1bmSzJhDd11qHYeQouRv4kTJU8D
eaorHNMFTErQTrOQYeWCNBiF7rmnV4qeO5GsJi4VQz5dk70EucvJSkb2N18l463j
l2DJtV9ZRM7bQZ3y47dfLH5gh0tWhhX939WJR/WHGUPku1nDnEv/4LC4sI0efw7X
6tC2O7xIW579SwrJddRGDa8PhkXx2+be5pbQh9Vbc0uc8VatO00bukTwSUcguTay
Nm6eI2J+6sXKcbv+my1jqRF+VKwBBYjEupkSWwmvbeeG7xRQniR0BZb7zAhlbtGz
V+/LEj3q42u1YicZQ/fw/zO7ASBAnWuxa2J9oOhPuqf1T6T69SYzV4dEBBH3o3sV
yIUaN8Vi8N/rgpb/sFTs7/113C2I3L6fDP2ji/Np1JqG9exN470GRiXbxYlPitAj
C+0ME+z0hJVIGYB8X82rhyMy1JQMmOKSqW0Pjv9qdsywrn7nBa7bcrZfDj1WzGup
1+OrYiYeaF6i/JSmFou3vrHtx1E/T3mQ/qY+8AegGRvaBUSm0xWINxQZYPTR3EX0
s95RYS/L5vC18Bk3/dRMvdTyr+q3gapGbQ55sRqzXWi3GCMCj5zoyEDmw/UPWs0W
yB9I7u3UkytSoV7+GZ1l/n5uPNn9abpyAjwb6tgFXiwRrYYJit0PrL7BqxpUIkKj
5CTAwYfiRHPMJCC3heKSnqb81VdcNZJaDdNadgo4TIDZJaa2FGNKVDmJaJRSCC8N
iGOxQ0idy292fq0t/bv6tYLQ5JnAx3t/zn2BLcLNcenRIqWPNKXjMS6RleG8nikH
c5VxTIcY0WPlwp2COnRo22h2Q3CukN52r8rE65hZG8SMeqU09ePQQ+NklOC8IwcI
/axUpsERVMSLriAOZmvQyPwW3zSINOdUo+V6Vb7ibtPI6VTOzKdJcoU8HX7VDk9D
E/3hdHu0x5iBcNuSGlWSkbTkMMcDD0qXm5wNfTKNcpZvp+iLuGzWPm8gqKjbEoRe
9pCVufDPDT/cwV8D1DPeSCX7hU4pHZb5ijX+283fAIRSGGVDWwQuBGD3qMeZTg5b
vwho4KHo9ga6BYixBSEj8dQzCdMgwwZbYCwPwwC1kcnkPIwRN0Bbs9vf8cu9kTW2
ah0JxFHT4R7bKvOUXqn0p+X5FSBQnv9S0mAUAR1Wu+FH6hdBWc3hDuca/yQVYluJ
Et8OKEUWrGFHeIdLPkgCauclPx9ZmWz44ijHt5bCa6fM0ttLsgkTrU4W7zthaJqr
HQCLBaGPO4nmuOwJ0QBj+2Nnuml2GTesI2L+JC/rqV9uuBFJ/xZ0TBKc4FqYtvHe
SgW46y0q9c5IKBjm/ZKTUJSBn4bB1ED3/yx19P0QUOjkJpaRa/W0HyifgoHjbag2
adwrpASKD06IiqoQgq7fLHGKMteu+KSJs33xipmufqb/haQUxh2+ww56631HKiVO
cdPYvut79VFWUpgghhYlXH/LESZkVO9dj2fzKqci0hUBoS95Hmi/Osj7ih5pGBHS
X1IbgUgaUthEuNg/8lYdNHBVq1qmW3EFMQfUG174OIiqFnR4dFnXaVEOf4SD1QKm
ZTcK8vh6duwPF+I/rc6MppIXSOUbz+whPxCWZWaPE4QgFJWePg3q1Mczo+bTK3Dd
lp6zm5rjmj6hnhiQr1BNEOnXJy+V1ATROmiFesEOjx603lccNzUBya9QrjLtndJZ
EjW/bRMbtGnDPbVAZRlO2v6Sm9lBTXLN7S6Rx2iHbMMRRQQKR3nAHTCGnsrCt3LE
+zN5Decj7VVDqNEJd81WyUuhbJbC9cx1tvO0kD9RazOig3Vwez2rf1dfgjh4250m
B0H+RGs8DYewDZy+AasypIvf79LS3s9ylYWuxHZrYkgWUHGsN//FicS6AbljW21V
3+Xx5S8+k+Q/RukKevQpfmrJXztM8nDZaGRKYkFNhr6Hj6o+ksIIxz4DTZAFL3Kt
Cf/5g5j8cKWGpNPWgF51Yng0GOXZ0hCYnbZiZWOObNYUBWs4Nq27EKXYN4uFP/gr
cS2FE++xHTkXj4zH8yNIPxcG+pC/Id1bC60quVeXRARZmsRNcjA5jMe1miuIVfIH
eVjDPTRUhXzsvWhj98orwUZFzTzxfVzZv4w4SeWbaqalkKI4Fo/cfVrKPqLzYshf
S8XFaPcM8dUztbOl2wm8/a/dqEB+lSv/HV/OPRbnDEsONKs0LVsfJH/dQ6zo0weV
2b1lVXJoJGpHfRL3L6atcnSdvoYjeT8BrjfWZkzW2uan47zDD0ij7s5WPK2zjQnY
2oNuHc1Q5bGJN58TlVCUTOsdF1zqYgkBw6SAS5HckyYbe/uIj4smGCt40fFepb8i
x+TAtN1dzJHzVROZ7K5ggMOZCNuYrLHt+PA3N8EqBoQKEVHDk5dR10hJw6W/6Fdi
5j3wV3In+DLa4DeHfLL5EvLj4MFWV2t79h+fnItl6h/mIPGQ+igyAAIt9Of+mopM
yvKY/+MCOTUH9rSLUwnM4FpRMtVquKOTK9n/BbxYtPmySoZgiKE9U0RSY9xRwJ+x
ROGsHIYcD5DxXyDdHWxl1iyMfReRgDcsYwGpagyKQhqiTk5YTCy1h4vk+cQWvKE6
EJDlzDaiZbtZ0jl/eG+S9Mtx+mWFHgu1Y8hu7onQkhL/xgygtk7SGPLWtaaxGZAN
8thu1oyG/tzAPl6xMD6Bn7vcnoFrMz5uTXLMe6dq2YWlro2ZNSXGr2DJZ5s4I5rt
saL0B9l5UICT93RoMs+tvY3Et5/czVykmPGRT46i+HsyUlWphNQysh9G6sVHJ9tg
IkyLxVJxsu6mT16Gb+udr/+JGhZzv/sK7h3+ahv4GGFoH7v95UeFXzBNVqOTfKP6
xbAxQ+jHWBI6sdRBzI5ncSGtdJgZwlj7XajGPUjNR8LkjLRMv+VBiFnAp1qC7Gba
Bs19NGlxUvMKIgmg17WFrgQL2hmDMM4pxDTwVsK7rBu4P8u/okvUyv53UmNpij5r
+N0SCs74qaVlCj9ieOAcfHQ4kRuYjVUiC+8Yu6CZuy5U7ivl/7PpvzY+BEVIgzjW
nQrKqpxXaGMlrd8gNFxEFldz5wbkE7IdlsXLXP+gb8QyIif1h9vfQvQkPNRJidNQ
TCXCoEbLpaFDjXld+NY6m+ECjpyKAf6/tNlV14YJB3NUFAs0fO/NXJxZ2+vd0Mlw
FH4kRDjav/a4K10sQaBSsDX3fNwH2vMD4pZ0xyhx11DL0zf6vhpFXsiAZD1b7A9U
C6cU11tq/QKdq49NvzxxfoDb3pi1cr8OpIFyTmaXCLF3jjjEyrXfBuAE0BjW1kyG
Zyb8tPiOPquUM6B9vGCOgBmixgtxgIqjJUNsPL7HKNVVP9AYNgBiEk9b6d/2iHcy
FC1/xH8I/aSO8J0iOfWQ2uzLzFEmbU4sr8c0KQlScqkMvPDtktBcmjbEyjgUs3P3
aGfRhdvZmW1SVgvckVRb5w6hIvzIwGnwysH40CutJAEa+mM1Qz8yYu5Oc3PeaVTz
ffKFkU/Iza3WBJtZePKMzYzRlRTLXaSp7jlPDjOBS4t6gCjfR4eor6FB2jDE4oUt
xquD3jod2U09idJaMiFxG+3CNJnBLq6mhJwOypJNpqQnGzr+I1/sKiOVZs0hoZZz
sh+hs7LYKFaGryJI45Y54YWfIa2fTzCYCh0UsPRvo8NrTPMnLmRQTndW2FKP+xez
Ts2loQqxeSlRj5picIR8mo/G9+LwaUl0A8/gt9uEE7d/aooTvEb+EebFzKF+4+8c
IbaMDd4pM/OOdPogzCnvfDic7TiuCqweszer+3KjHm3tO0irziC6R8M3dLAmn1Zu
Bf4V9NGf6UoNHdKadykSiIJJq0XEs4YOlnkUJ2Jt8SK8Fw8LHrhMTnk047NDzK5Q
HEYIhfzomnxn/EviXlhS4/xWe4+VpBfuV2X/FNuIemxpF+x229DMY0o9MK8EsGs/
26PmsCI5WbCeeRCGjwP48Z0ULNgurtdnUnFYTen3ONUnIfrhyEMFpiL30/V/uVqf
WNpLepiYQLp9C/IiSYTtCw+sI+6B/L4xBa1CraRUbsqtd7Yz9ve8Pm2t+dFt3IQc
Nh8rR4/DbWu54PI9ao9XHgYGr2wPw2WFkhFuqgu8WBMfZIs9l/+8SNvNJLl+3JMg
UnH6gKZ8lVZpBVTc0i85a6S+bmi6LqVFCbgzg8/5v3a7kAFhWQwpNyR3dNpYBMZ7
lx4xo8MTxRP0FLYJYGeyIo0ON5KhgldsS6/YraZz4qlMSaigNQBo+JoRRDPVHOOU
1haaL5VQ+MQxoj58yob9ECWgIRVJKIHmkwVozFkgzvWK5ALf4PAZVFOyaSoQfFTE
WAEVpkwMDV6kTeGlJK8KsKeOXgEMbMuhaIcTUFLwO3Ifi29VDEWyHtNaL+p1pgCE
R4XGiLK0ApQWdQvOXzAQ+Jq8pvBBAQ1jWdLEuhkY5pfR4ah+jMhr3w3EXxNYo4kg
5RKZ+kJ8AcMYKcu5gco9YYF1tBY8NlPPdasNxo19lbyAPZuX/KxOSp4LB/rdLuCh
S63vKEgD/axdh19I2OS8Msc6YJ01ZRXLgZltOZcusgVGs11bmp8YxWGf+8PREXxk
O/8SZfvkVzmLPPOoFWdRSescz5vV9ikv4v/Hi1VRxWBknkDPZnBaTEl1aY9FMQUa
HiO1KB1ehbBpNiAfK5UQV9EnKWhglCgOUmzQtryZxF5bwv3X9NeoHvTTeGZ6lWzy
Gm1Ysl+6t4m0/8dOf4w5HbLSo2bh88QhSUhJNxw6UI0l7LaJyoxXmTaJKd3LzPTz
Ztfpx7NWek26oqqAMNq7UDQ80kfk+lAYyBqYO3x/U7Elqf4nayU+zilDnqOlT970
Nn1Zv+rTL/XUwVmONKvX75WtCcrMtPRBjBdaETpYOs/tMzCYtxlPcyY5fULcUyWe
taQDIFpiFpAAsfhHe6/5viKW5K7RlD3/V8JWpcBxcYg27jLKOtJc8TYoGhUjFsjG
s37Lb+3dVbww8dafUTeuzjALPe5baxRcp9MgWkK2m3DqN/aAcswjYx+9VwInplqU
aDwAmsrs/Apkmc5UoliyVczvorvORAvWoWlQCo/inXRVjdcw6T3aQ7IvSKMRFV0Q
z96xth9BTvGreiXC8GXDPUcu3nMKQ0cSTrWn0hPedLSkDmVT5zpfvSqWmWgLus6Q
SEhBpDxX04TezSl1tziPpiFuoIEDeKHfreDRxzg2dgGc0QS6EBGZM51t8h/HDUqj
BDLX4VAe8UQCXpG2M8opbWMX0CUoelax8I1u0XTPqBhssfeKi8qTQ6EtX59txN+b
/mbxNMsNsVErRvNq8ESPBvsclDuTL7+T9YtoLlPNv9IoYmVHjOTpkqQOcAAhS4r8
6a7KMrijqpaAgiFtd4cBeV9XPnsMCoFhZO7v3U4/PEuxOv0Q97fGKekPDu5IbteN
8MLnsP34QZjZca+LAFkf1lxU5eLp/qKCQVIQJ4BHeEo4GEZquEjV8xt/Hq2okMCc
6JkkRN7HIEWh+muxHEiWc+Z9wHofufqZ6U2SGqG4u5hTVeezo43MYMTfYoFxnMND
AVsEhtw2ACqlgJVamkIp8KnzZy9/qFZxzT/jYoDtWsFsfBIskCrIp9YaZEitzK1j
y1EaNvEN1pzlRzjl4sYirP84HXb4+XTKelGLVu6yaqNaiBSpJv+apqheGXjm0/Rq
WCH99pxHYzxZayRG3rM53HJxfYf7qgHD2DBQwzwb9p4NJm2/8V+sg/sM9JvHNypV
HBNLZ2h0389u79CQ+VFEtUUIggVZg17t1jrt9VfzMJGmtUGTv3zHh2/mlXNOsvls
wVzuJY1y4HHLkrHSc62vRe31qXXvDoiWaMUjPPtCAQsyU0vEYDbchbP9qrrSjLV3
m6cE6/rtgCyoa87JsnA7wZbK5jK4yzTlupZh5hQDYnRDJeeui6pN68FbRzxLruEW
1gHHI574T5HeVAxhCrVkT34RGRdlI48O1M7G6G+CD72zXQC9dgk+oZDPHzW02svz
S+C/pGmijoZNWMGngTYMsO/X7o/qcjHO2U2T69RFaSI94b+SFJ06lsxOhZy5S9RM
K1YN1nKXaHZSU8L3tgsgbX2CI1W8yBUUi4VNxLaBZo/3CDLMPPGWTsPQXk/5BZBn
ENeLEvG5375gNGH6u/t/fOplzjtrpBAa8HRL0EaCmzSir8+K95FE6gJVe00mTKTv
VVcV9OHSCtSN94R1qPaF4GLTyM+sUIOXBwuYVf38PGWBeTvMPU666qw8UNTx+rq2
rVOvi6urmhJWdxsctpicHDFLOMKqnuf+acr41iOkpHC8qb5sHH2Zq5JouS645t4m
/TakZIcZTdSNlQLEj1pYljbeOnaIZURx1/57mbYXNhoF4ZkWAHdSQMVqD0ynlfpd
e7h43oYJOsFkQhoc03yw9dJmKiDr+5wuZfVGfxYP/4S+974RveGu+cfon/PcTVf8
t9Qjy/BXs3ya/IDcMqnoH6V8X3bgIbd4/lMuhCsBJwvm6dhQk7R/rSfxH5vKrM6A
6+cMnBKSXcqwoBEmow3WL67Gb+GJOf7jXan9rtumfkTiE5kSKmRa0dCjEJsYSHvD
G4VJBfCYIIxHacbZ7gTCJl7A4CIlekDxzixmWrYYxGl//Ok5OWPKC6J4qSA43TnC
IZ3srO8j1R3uQJohnD5Za2BjwuFMsJ+TQEJWrYCeFqHXxi1sFOU7SwPLrjA2Qlyk
ramDVuIm53PcI5eUzQHDQ8GCzFcHUjnMeciNb7qhmUuVoxBmc99B4GZDV+dDv+Ed
bq/RuAVmWxQkyMFBpXnty3kMAf64moYQzdjynQaCENougEvPXXLcA2dsxCM6MN6R
j0/4PO1GbExvVdh0EtM4IzqhcVC3X0jF/3PsdpcpFQqamhrLhrFdi/jUhiU9kq8k
HcV3HA7gg9Hk3hrvu97Cjjyel1kV4kn1HElpnTLa4FcGAF+H/X8KJGe8IkbIK/wg
xmFVUK7EUb4fM1eiFLK7Ktmy9TgNzaAikqu6UHSpiDs6ez4XoEoLL5GVnv7FSbXE
/M/c9c7QXypi4Y6WbHV9pbr1Bddfw8upArl3bHTKrZCx/5uM4hq/kVbBu+Pj25ek
f2CJBtYflYVDnl0fWv3gtIkVdpzBlG6okTd4XOoDkZlebqF+JhJ/A9d9t7HYXSfI
pVkANZz8Yu3wGkFHZLUEKYyzu9W+ltqOpj7iUGrc6b/Qm+nPm4evvXt8oI2240ew
ToSpvm9MMEiy50S9fVVILNkpINbPEpcvq9rfGjgW28hogaao5ClEV79v0qHM3EKt
STzZ24GCan3FDnUIOGSRpuxF2cBnssUJReKma8Hb7XnIYq/5/B2cH31BockGy/qU
YT+XlfHB2pBNk7GbAmFDrP3vKHVimNIst4jF2OJ2duo+MtsDI7ejaXskYQ9yeMSK
SElUrDToMj6x0d1vObIbg98z5cSKDeoQxnjwQ1fAJY0wRsLkBeSglmaJygk6hYdu
rfW+D2ovR/R0VOlwyG7YS6aTxwI9Hw2c0/SsQqDL0XJhFrNjaU9L6Kdb7i12qFNc
EhmHHh/Jf2ZCTZwZQt/BZjEgD1Wf02jc7y5OsRCW9So+1MUIcuZgAZiPYA4+/pTB
DzCxj+P04/hmvG9+OQBjlzfmZuIkCf2uZBluWV1v0DX/HE72xZZ98PZwmzpro1/C
eBXDglT3RsrcQqIyD4YBibet1+FUwq1FshOitg6VoX58dvzlm8mziL6hEGLUukMa
WqJcxt1xI2L+p0hUTSpvu/b/BE+GUPX+tEEpaL9fnuirWHnGmq8UXUFeGDyZBYpV
DBPSyacg2V5m+RwyX0J5NS6fUCfNCn2ZiZ/Q90wDjh0ewj8SE8sn1QQpVnwupEyY
bMs9Pbfihn7kW5y9/AwIPB6yJPZc7nLJOFS2+tyCaOKSHcuApqapS9la5y6OYYGM
Wmy2faRwKrA4M0jZ3zd58okkUK3EGaYMV9MfctF/nT5di+z6cuqwIfzmsOIiixP0
WWfHo1HhDrOlnDVoWTMu7XFGMRY36WFQWrD85bYWJdV13tJPQVV9M9SNYObX1TTc
aPrDx2DkJa0352qnFwzxFcDrp477AXY0gg2Dm6lRnSIFUjXpuIOJoYmE+cb/qJ+F
rKN0n0YckRnH32jMeWCscg0MU3rCuq9QHUpT6TDKs5OCwdBcLo04SJ9SiK6gXuuE
s6sXrQ/3SXIB6dKEHxqE3WSqh8EL86Jp2TUflHDIjCs5FzyDQK9l9339CAGtHdmg
HaN5U13wrbltgfnzIHiZ2dS53t9YXHtMXyEuqZm9VFpo6PSNoYO0iI4yN1XZSyuL
aZ02O0ji+J24TWHBovABlEfevAiaW65cahlE8PkGK0wV0gEf4dRU9ZR17fXHjMVP
Vi1+okZZWoONaVjcZaj/i1Nr8bhaqNcCVj4UYmvhRetWiyrvDViqE748116hlJ47
wnC3aFPirwCUJSCDzjbDyXN4dZrfGGbnXkNtEU37mcKFlQ1mG0YwjLHTbiEblIHK
nTev3Tfsw1z178/A3o8VkWUS2+qDaWoTdeENhzY9/JGXXRcpaFK8m1oX/l4EZsYo
SsWw0o4LutYXbSVmvY16bOcnzNB+wtwOaXM4Yiy2gX5ZDMCHw3sRPXVm1wcBhQN4
YU3x3E+ktJ21keDHyWZXwK8j5pNRP3Vuessh5w6WO8/tFFDN0sO+ZDoe8smkOuY4
wcREqMX0idAAj7ShDGtbD6g/jEXLlM4sDw6/4qhhX9ExtBd9Jkm6GcKJrbDGN/ly
1mS7Jk8uTu2nq3EgDngOJO0YjmLIrqpUHiKrlQZK0xorq2YotKSPS1IDIGYrwUdj
l0U4Op71UeDVXxk+5YS/OMW1QLtHa3ScBhh/lmikbYC+yDlWXRkBMev+oWTXCHgh
g4AcYOzjsNzRmYS+VNIJmMle1eCDNKs5aIbtv59+Y4VckqxKwTjVkIWs53bNeGRo
BjM+11uF+Y4tRmJzNp+qBHqgC/FTYfYI6W+hyCM0T1T+saJb0Bm81Vwu9YaWljyR
cYHzg2PgbPM9oDkM5UCnZ/LViufpF+5VcYb0nVF5fNyUP/z5ziQJA/SorNDZPWXM
I4UnT6/oNkULbt2hXpzhGz17z2QgZG37QBNUeajtw4XRhIg3GLC96bYB7hmy0gWx
blhpIPI5NW6vg+NWVHCY+Bfctd1Qxbyl9yEZMcjEFsG/+ca82EZ6zwlTT9WvYB/J
NE9p2zw5G3hRBpuDE+bqHDN3G8Cs/m7GyUeBfdZKuwk21CBeVjU+FVLwVzLNno3u
BUQEenSIktGPdRakFTEOTPfEs/EfOZETzUDqD6hq7yk+SziJLRiS0iqTi6AG6kGJ
FVHhTJWakkjTf67dVAKyfknRypUPbVdy6As7eQQxP/tPvuM8WjBh5jn1eQfB6Xod
aIzVCwK+WAEJrAUnDBNCnT+eXsH6vX9Sq1oFsQ5j1ppFWk4gRUXwI2rntDZzRTqB
P5oRZT77p7SWAyRhPUzI0V2LIXDlN73pc0+UM6pzpl3JugAtxHTKaG3BvRsZNOBQ
kmJGgIaa0Q73GcyGBHsbTqtN1fiRUXxheU/afJnmvF5lSczVu+RKEOOePJi5azVv
FZYtA72gKB8tLkEFSDToKxpbZkU2uePLOgohysb960+x7LNKfGarnmPhAayFDvJs
J3TluzExzEMEVNc03ouA0tTmi7ssl9eQqcLgFsvN6w0qCdOdHYN8OMftcBOuUbbl
3vaCyFtzn4yKyZUh2GzJaSXmNTH4SSwfI5WA95IiZZ61I280xkoQ0DMyctoiXwC8
Ck46KWregpeIHhAthGlq7mX0RayTYAq6g+BWr3iKQ36NTcqti/nsrNof/RqH2EsK
LdHIVHhf0lzXTzsU/xnHV2N5V1OlR3A6K9A9EoMw5CZU5hyx31X21KmH4ljd31+f
+DrEOd+Cb8Iv5jNj+ekRKzNyPj9+jyEs12mNjg4nH5Q6/pIo/wsc/YKFY+6Cgf9O
TvfsodOOmXeeUyDEQwBdjDvg+j3GiWTsTHZdT3wISRwAbcPloq/s+WlZ/htgGMOX
mi3ftlEUvFH+3AejMtteBeQivrozbp59KeoaVqC0YazBcVKBdJApwhSdTAkUKu6u
MEHZTObtpphSxU0/I/RekaKnbdJaoyqSATHyd3NVrqvulDGNqmOIicjPVs63nfeM
kN4bCAlGyTQwloCakgZtZYmoR2GLsHL621bw7dvtlUSm9M+5L6xG4JyVnwCHu2zp
ohaiG78wcG9/fyLKSlpQahno99Z4Zr97vW53vXTER3RFCqZFfdZmwx/bpUXSAxpp
DCs6MaCEeKVKfq8N/rRtYgwJNYS3IvMptnGTcA28opv20wQdI1Umo4tY2y/LYqai
6jkWNaDtSxuZvBeAWmMBMrVY1bEHzFOakNiXeIwrwE5PI3i10KsdSxv9IZapEIdK
XAAlmy0tnOSj5NH8G+BUw3SaaAKXziTILoVOkyyd7Z/EXhAL54WmNzlgFBkPcEFX
cdt+rQifRtg+CP+NAisWks2NI0AfUKtK9XdLgexpVyjeSB2L/lCWTiNYuvUWNkqR
YqYqH2prElpwYugjwkRbDZhnDb8F7ikycZKmi64AnUedxUBEKRluL2h9NxdKOh25
jy+yZIqpOYul7WCBd9DIr+h0l+/FDici5TXQikwNommOYVIR0+Rr98EbZRcUYCZj
lKPTgtsQQE4ybZ/fc/YT5eBbbz6lRtLFZoaoE9UTeUdvN6+cwCJovWFmBViHF81O
jjWaILIo2GQ7U3izpP9d2KhNoHDF3pXxow1EW9QreunKaQKd4AVPNT/xUYZpz5AT
BuDPUE6HIzk2Q4BEeobwjl9bo5kIJWuqDCnWgRnMoUrxPKGUl3iVIt3qiIIcIlGj
4kOsNJHvm/2tupOkeMqpUy0nIzSOJy78BGdriWtZdzGsRRpmuo0WnKxfIgP+qNHO
zy4a83ANW7v+e7+/zdFxNncTJye+Lo6maeVE9C5O7cRljYW4LMdcPqqzIZShf7wd
VJsAwk2asU6hn60ufrKK21gcinQFumykuxXCM6eC0oap3c8898J4fwsvu52FZKpX
K6cN4JigRhZqtb6xU4vVcv5ZJyFnkmUIKf/+myzf7LogEWhCJFfiJGAuA78skg4q
FcYIPa8beGjiY42ARyS5TCgp1JdeN/umTRpAyFhnDUeruVsDKtQ5RKWtrBaPoNtR
sXxsBAsqj1FVwTbeLsJ2Dv7Z7w8jfyKQ4YhbBwDgy/SNH7o6lhWZ/ShDCFqETAoK
aSW5hk+uAw9V6M7deBZJKmSUes9LaDDolMdl9++DQ7drmB7fyMProjpcjFkqIuC+
CT1EUK27ewrfDJskMAfQmaEjuswJ2ogoI5HP9Qh8GNM/skYxbq8U56IXTZdQ1HmC
GjNBrLg2IUa0OXpRGvHeURyeEVCtFOdzocr8IbmPX1GxCiuvpdJdy1hFivDpfPIc
MbyPzJatdD/bFvl3ttQU3k+luvmgqzkyXaC5CzUveyiSJiXDrhchzjNUQldQSg3d
1iRtDAS8jc9SYTfGWx9eTBcmjmRYmki2U9KOXkjZTlGT8QVc0RkRII5ArDsL9IBQ
PoA36wdJHphkDbY0FGnHQm4zz8lq2HUzw/qM5Kta5c7cKt9YsuOhjH8Z1fqO0Vpu
0W9cSeaAy52BNWYhICiPf5h/zdM21OyFs5u9z18OlNOp4U3IGaSBr7Akq3USRFCn
2PFzjnPIGAU61EygPOhdmuJMdC65/xwN+mJdx3Zw766wBGzYYc33OXvgR1ogvNmQ
v3s+qqRoPWpUY157zMBwtlrXRwlyeeQiBJkVHQcUHcT70b7gvHrrU2fiDi/6HKT3
JbITg/KSCr3Fc3N+JyjOKR7M/SzrO6P11kwM/1NG9O0pDT4OkSyuDWnbE6+QSf3f
5n7XfNTC+wcxfhsLxe/ze+0wtbpu4mdH/ZUo+iW5zk40mMy3nstxVc07Yv3Qh6rr
tWeSclH6pGQBYOX2S8ffT7/UeIDbL0HIrBdikaDg4Y0Ko1UUFuUbLjxsNQcWtkf+
hQw4796RDYwQl+Z7LhFQzBfRa4xGLxDxN74HEuYPo/9K/jnLyPvkvxeyEbqKLh+Z
2/qIiRYMPBhY907GDG/7o4KwcOmjOyW3E+iYoNW2jztxY+AwSaThwBpe/PUcQ8HB
9yVv+6fvqcqSC7EdaFfW6rlX9RFpH8B1oV3QITCB9kh6B39+CbgQ0hU32KQAkbPi
3XIkNVVBHvilX8tjte7KoONc7f80krMOJTmqV4gt//VcLQ8OO+E4jbcIAZO4ephc
7azsWKefzOV1K0ZqG1yhSVROkUxTudgx9Irr5vP+bGo9P71Q+94VLlmk3XgxT+hU
10Q4QFKdZyeHfcNb3g12oft1+Lcbz8Cd2KwMCh7PP7PYZXdwiDimAH322+Dcm5XC
dSVJDskjiDGu6f+pEa8ZFgPCPSdWMxEnpivn3DyM6zrCoLCi6rpdFwxxGPblmugl
okVeZOsPMWjvlxF0lJSozankcknQ2qfxf9RPwGtJM5p3ZoRUPu8Nd30dRCtQlzFO
MIdVIk+IDCxqQvjropSPlTZta1+ek1aF1lQql2vujUwvBV7VoM7OrkGXplMDzp6Z
zT5Hgcygp6CLhR0clBCq77auUBTBrAebopq+R0Q9FCUTcXkxDqTMC4U9wEPZYflV
fERXnHYcO1EbM74DLQbzZvmSM8teq9oVD2z27g72T38LW8rxd/rJYtitpSQzCw7Q
pUN2I4HW4rtcdUeeS+w4Hy/DcwbuBiIvLH2nNsUm3ZWlmgvghJ6xeVCFBVeL6W85
jI0X6W03dmeOSrEmL73Q0NQBA2n/HzvdBZ3IhzOGPLGP8QUijEhH3Oh0PIKGBvux
Neqr2B+BbXygciFYrPPJiMrUz5ekkcaLMci1wFvsb30+GSxNO9sPS0+PRHKDIKHQ
Q31JdVoCfB1RuW/Ax98wlRnMJiDb5VB9Gaxbyx56CZjktbNalrpgQE8jcoG/BjAO
lojvgY+HlXBT5Cv3UYZooBUL1qg8QWkgsw9EzpTNw5iYPkkp3Ujb42EGjuas8qGj
QigUMq3pGZsNxHvCCj1R+UQnwbI0IaEdxWDs7w1A8g37WUnFw/QkPa5ECqYpXJoF
PFV1z0QA4qqkBGIoSlOVc1VrAUeC4QryaRrR0b3adFsstIRYBvVlJCn1cHQLI5dm
l/4P29vOUhMlb1+fZ3Mfd4z7yPSgK/wflLQ0G7JHzlbwvkxx6dBIq7ILnE6ofybd
HmfdsL2wiCQA1BMhHKo4LFlzrGNc7UBSHO4g5gmR6Y1PeN6EGfgs4hJq9i+iitXo
3Ze62CH8cxRiaVsoZv9NM5m4qy9GDjj16rXXNlRGUyVlynumKaJcMkRLNPHS3dgs
jHmGgHFNcqpYV48TEQUoVI+veM3h2vBSnzQdjNlSg+qvUoosLx3iMpBHAa2YyHhj
c9iSVso60nXk2qfpTij7+HG0sMUfGzUKPdSTuW5zC9HuM0ga5ItC3YDC+Ft0q331
vKgo4fFM2H2QhtbbyaEvyszayg3TujJNp7yxxRduLxOebjY+kS9nRCcvR/yY3gSm
dpTgNTNl9SBYjg63bho5jE7Ttuo/WiOlXThY85xpFI+WgfAMPxl/mObJaFqUUhCN
yTTRLSx0UB9iT/YvH8dnGZHw2Kq7xxQF62LFnqdmU0rOkJ67ztkph6CYYDJwmJBO
KU2JwGs8ncyerK1fJn4eJdFIPf8mWXQ0VdIy25ueq9S9mUoYext9YKilu5EjrXWj
H18H5imTl9NWMUWrRbN9CCLzNaxoZj0rWF0Z8jIXZlNZH028YLV3mXakI775pkVE
mQ/jhdrOqXOL0umVC67TNqUzgj31ue//rg12IFHHN8Jy/rf/F2UYlI3JirR5+59K
Jwk/C6qQPVtgsNoV1ixH9ULNMSHVtDKtPE8YcquriziuKKwNGqWCjJ2gEheNfuox
RbmplqQ99NkXGHl6lvPWQr+GBm5RbZ1m3N+ckXS+POWC26NaFebd+Q3mjBS/7/xr
ILVZEwqa+9DKwdnXfhuCr23ZI8qOnU15Ocu7zdqPfUbo7i+75/+okRXntU5Fa8Os
gum+oStDFDmiB/eYt78Or1koL5oK9TvAea30euraSZ3Tn7i3O/4FqLUdqtzAubnT
w6wPcNxW5lY9/VduK/pasxdCKJHIZ91kfs9L3mmc8nuV1LR6wyBjWqW4+6UtAN8R
9EU9sLIvT5aer4EY42Xup87LdoQjjmASRO1tB89Zya2qJI7PiZIxNZZHNqAHeeer
3HqhVCo8Xq7CtyJ2NkSGdQaMGmJKQLUtzL1Sqo2etYufpftwvkVfEXUlE+9v6hx0
TPLW9wETxu5Fq51rHlobmT+EFlgiquOHRF+Xogq3avQd/5ULiAhJtKFnbSPKcSRI
Tbv5Q7az7jSqw6Mw1E08zdHMzlCP/9PQ/pdeojpwUbSZgHAh43oY0zXxZg/HogPD
O7NScX5PWfI5m9zdVhClfi8RUZDkVRRPHOOhpTXkoFxgSWVNu0WQHdlqXgwElhBV
wL9yITCGZFivLbyOG9Cb5x+I6ONMGQ93+7CgC9ToMrhopPw0heShUM1LtpFoVT2M
nVZcB85IYcsXSIy5c0Ub1PP4PyAd5qUgeMX4Roxps8EHDOgzPvIi9f+uOK85n8rZ
RcJgmbkroShKj63a0eSANpH94davDtdS5a5RqUbUc/jXt9L7kW70QLEC7Z0Oulkl
XzJQMXosX1xcxaU6srC6I+fhAog5GmlPbOnR8gO5KKr2vN7DY0Mqp9vQppcKGnj5
CR1051eB8u6O837JnnA+W5wqzeKXvX1WktaBqlTZTSCAfwW2EIFtKjxZ/0V/qGkS
laUZM57t+HuMS5r4LPXEs3jUz/LrVzvz7rnTo2qHc2Te4touQZ4BmXNnOwhkLvIv
9VY2SFd+CGIS/xOKy4y6s2SOj/5y+/GO7xsv1isSQ9+ctxZHiJ9vgipQKurPNhsh
A+Eh0CHAV79tGf6R1LJNmUnYLWCKS8fvDFwnDSG/DLyO8kJU70W0Q1YECt/qC5H7
0/c+qLIcib1bruvoevgibsGIYFHF8MVhKKxTbfcjmZRC9Khk81nH4TjQrGhykz/A
/7JOAVfJwlOUkTnRcUOvx+eYMQE5v1nMrkXOvau71GQF2ol1HUC8sDPu0K2kVG19
rgEPHXKz3yxdzQly0NY0AAKhoh5Z+AtywTy3MTfUQsnQoV3bqtMWKwWYdbIOiOgq
HMlytFJXZviYW4yLuPULf86dKrvYSQX6BsMgUMSOhavViiGy/rgswgRWf1A8tR0C
u0awq+JnTeM/sXIGZOuKUa22tJJ74VliS4Mp36Xw/hP8bMBGmISZeHtx9Y/betMb
mljC0gjB4jJpEBwhAQUJJr0GQg1mjaOIvWB99iEtK4DNeTzILJb5Em1pP7D4qmnD
Y4T89AEy6l1VKhDsAzPtszw1jMDiU19Qczi2rT3bTpvNPjzbUq+H0UDxZAnTTzK4
VhVWYTP5Fx0sjkgfVH+kTqBy08boHNkWRcavftKSaGzRnA073A/HiATP6h2VWneN
369q9zhnvkPeazsVtLM9W2/0vJuJCLtIJp1UtvpDiQgRb8CsVqGviruLVujEmCVq
aBKXlnSv6a52XQ04lrI4F0MD4JwF6/HVSifEXmiDHFt1+Psbq7vcjNjqsBQ844ml
RBNmzRxPcRAVwEodLfhlbXrFeojJDpEaZ8xccVH60Je8G5paT5+SuEabwljxAB6V
cKs/Rnc0KrVX0zaN3M560qM8QTjzyKJFQnQxIPh6xWKAtx/9Y4W/XfQrmz4iXES9
CfJKdpG2zV+Dxl3yRaOQsMMqje0MGnc65Cu2x0ShMTN9qQY/77s9Ye53hkZy1Bp9
crWKB7RInkfJ/cj24LoL24mdtH1LhnpDhaaBIiyptYuqlWC8hRVjwFNAdIrAyezC
VJgtpF96wputEp3ptLktX7MrDUuTUbDJXqO4EVojQyCLMkFke6vc7tJWvH0YuGiz
aNJLAZimcsh8NJwGeGsh1YGUKgVOea5VpBYT4xBiZKqb8kmOYizX1ZBwa5ahhBbT
64u1LhhJuACPTStTm2mIk1gGfPFbpcPa/SOzEW+uBNZlfU4NEIFufbufVBzfzO6U
+tl/adAhXbt4qOG4XriUfDzA7Z6rSJSJz1PkaBS6ZSdbZFjmLupuyxcPY9jtMafD
2gs70tsN2SsER7pmleUbyALTWcL8TRmUodFMb9mo9GHoY8lo07WfFcSkDoSrbCeb
Bg+F4zeFcuNSzgFsHFzraHfEXO2u2HJ9dmZkEM0fqP3gMwOWKrHK77Rznc3QN1cF
6eEF764bASfh0nL5b7lo6fMNa3wFdPVIw7+HwPAbMj1ikWT859IFVb2jxjaGoAof
qEwO2aWGUARVBwedUdM1SKcttedcoQbi92rzTUwGXfdNF4/uegcBMAg3QVmHA9e0
SaTOGg7meERjb3/o7NPji9xx3uWCLdbJ7/agaIIDZNE4V1ra0yTG/hYQOcLhdRLe
r62jdxyY7sBVpS64JMWp033BdUPDpB8J1vIoCkpDyfbS29r+JztLVb64M5TIdoQJ
yh6Hux/CwUZiO7V/R4LY3TDjnxMS7+vdO/9GxbTEt9YY9O16DzfHCMrpqj5hxtxX
Gts7XB5gz0AUszicsciePb+jzTiwS0OjFsxiu9e1Karf3n+f7nvfpfRcBGT55EkI
j7DrI4zFxvmqqWsytvIQpy+Kut2v/OhoGS9k7VOG0dDOxAdG/3U0hidECTAGZyM2
AFOgJJjodYoIIHk8JP2ogZRPMU00zggghNIKHBH001LFxRrY0N+ZYP6y01yE6J+p
cnOiuHeDdiFc8Uu8rdnojpf/YYTojmGBQmBErz5oq8v5wMulEdUWE3GiRhAv2hf0
CBaMUGEeDjINcJJ3jvcDpQrgG96XjpvXG7CdUBCoMqKM+2cvFbs3zDeix+U03Owe
eNFVBMTYlXrcVt75YIUfF9pPxuOuqsgafDU/z0duaD8fsJe1/V20F7yNHmF/XXS3
pTkT+nCjG9oDf38nt6j0m1RvKM2uJ8oOl7P3LXYyBbhLfIxWySv22Ibml00akUbu
wpLA4do9EBNRFRbDYu2M0fXal6x8rbrfhN13or6Hgn1UaDCTckhDPQDgPwCDSWco
JjvTGn7GN03gC8p1Op2Q2caYdVKBrndVl/+hjitKaI7DtUKZ1WopL9p34XOOYQtT
Kdrv14EY2t3VLQrelaGcfDDY+Ce73bY4XgI2hSeEOQvqyzd0pZzQsP6aDVsrSKXs
/DwPJugRZnhZm4lO8pAg6SKZvdCvjHMR76/p/kwLZ+SWV0en6ruUlxbQF8iNJigB
v1xiPCEm+eo97rNAP2vVryStAqSRR+7v70EiamS4FORYAsMQHK9p/qPTcidD2UkW
k/fgwkR0SL2qrZ/RbeEazndcHInXxS0JyonlOQSGtj+Rd8Ydaufvr9fwxjHHB9gu
AAx5YZgI8Dp6lOzycua8RRlj++Ev0SpJ8pjyavY1n3bMPvQifmRIlSexFq5JpgaL
AgIHbg+4ca17NPJwY+2+9+eoGzzavtThZNVN8NxCIZEqVuTV4LQsCieebyjPz+W0
xoGtsU0W8mKxsaqEr1gMbOMgDWAtcC3D/1G3FDerQWcKdauUWeLq9VMHjYM7/g6b
frWFSFYoH2dF/KYTyqSDDhVTbwPImlb/m9Q7kUyY9ajIR4X0QY1JHTQW++S3zXhc
a6828vkZY8cYeaUf4tg0T5qmNK3FV1gIowYXMNw9HHGgz9YNdxApB3/lgsE5enGS
dAMNxp/HrcpzXFfnMv0n3FwY04xpaGRAttnjQTq7wee+Dau9JD8hBOB0DBrIUKYC
ED8eM6uKESGSV/LFjvWwGQPAaRqzZsFbaDahrMGiDjOi1CieAZigZNFShcZtB+rx
DYd0QjwyIiVRbHSgxhV0B96/AhwKcoQKIWNSXqNNQw0gd5f5gGDju4IGaoiYPNJU
BdvkynhsnFecX6xweMM3jGYm5eMY7UEHPncNPYkkE1xBLRmycqpmfzXL4bgD6ZSN
ysFieP7BQ9O+QdP5RPqmEF7V4GuTv6rfmnL6be7GUGI+J4GROPydlsnrfV91u5hE
itjF9NFWmp38NZd7NnDWm7RR8diSB09NqnLEWdNZQ/h5jjDO9xa0eVfXG3IMlsHV
n2kz9yOIylQRR+0wanzkcdUGqDv4tLltIfhpEAyP/hlHpgcT5321hY9FUXEvivYJ
ck3gxARCdG5JaXXdoNjFoSb+BPytR1ZvJOI9YWpZGLk0x8VwoJRCaFs3hfnZLwpx
54XxmH+EU39/n4OFz7nVUga2cRCk37ZRRAjw3IgYAB4SzjLowJRuBWUFBYvxlu4O
tsjJyKvoG+zEQSCk9J//hUI/ddaILPO4Dj9o96sVry6NcISAYWS86YzLkRyVYKdH
BYAbPuOB1A5CvfkoNZOLQKl4dsqoaCecrUY1jejc8PckzPZX8AeCvlA0Q31Wp50w
mzikzXEl0qXUl3mpQ2CI2zfC7VFz1NOApQYwxGwar9yWlLyyDL2YQfTORTmGcyol
T7Y10LWkQKAc7QdKMDzH8S8R3HHCv73gyPfZhxDao0aYC4VNwjgZM75UDqSBC7YQ
SU2btNpMRsAE8oJaGd9neyxLvx3bCS3zLMOFaEeoKji1uB7IWRMBMKpg1XVPCjV2
Mhter0Ep7nZVax13Y+3MGGtSOdmuOMbO6wqSWUfOXbqTegtsuQbRQucDJMs8kWVl
csTwWVdA05RPNKk7AxCWjGBtiCqqOkMBb2AbkyCqmOEtLeOSR7PaqI9hEQRXDFfs
SIuK+vA6MfYNDARzsm6kDXzg3ba871UeHMFsjAiGcI1BM4jhd6s9icGYYxjillYl
hLzjD9eLYVBqCKDTlo7nhKRjXmKlybkNotrlhvm+q/yST2WXjfSLNsiA+ceCnaPv
1y5su4T61pKYn2MmFip8TlnWtIkHCGx65s3ErqdZTGSlG/xGQvBvVpVUHxPaYJ6u
E/l4QOYft3vlZ8D189F8C/JJBOhSZp1SgReTjs6V4+FKDi0+tHScjYpFtlBdHPFT
E3POfEkfEge/fIXrpV88VKnGYR+VBazzaMrZUWXzD/jqk5p28k2C9ad7pvkrsFpU
MMaIX2Uhq55YSlm2VFcFngZywT9UpHuFgjZf/lIYBOJUYCtHxA21vRWAouvCnN+f
HzcORP/KsNbWpoQSUKIeebOIg/WLiy5bCMcyZoA7ngRwUSgqeNOw1DQAsO/cOiuj
YyM6KfEljTnqw5PO2aUoX3dATqGdMhkw+WmoSBRl3ObdAODypv6wzWQq+r6+XmFM
MSdR0P6+n8JFTr41XJaoyEJrXb4YhU2rC+voNg18NTnq2L6YNqvu3/KAIGK/3vvY
dzKRsdvvkjVbzZUU5DtYBaDrUAVboGuINhXyZkHPgp2+ZmfxfMWVcr47vE95UxEP
XTencthOuXyueWQoKc8gc4jjbr+P5M2jpMMX34LKyb0Vf0BbrNcapJK0EFXN4KV7
K+78xbi434k7ZWVfY0zJjLQs8vZ5RlycZIxdn0EmoJU84c1pg2kSA/bl7avVVB4d
vKrGgcV04jTkbSlz+W2aoe7saUvokor8vRTm46QTNcg8CTiaueUOxa5aN5YeHVXw
XcOVbguCLkNm8wkZvwPvH0nyc81QuHIvvNUfbyj2m2kechc/Wp9Sg5Jh6XggVXMD
wqSX/yrn2iZV2Z05pgpczrVF2Z06IqjKUAE91UueSX4cm8Des1aJ/5Y1eqD6uObx
53OnbjsUWvCfiYgOTlffn3nyiW9NXCvmbneYJ0AZ0DY6AHIiTOUyY/HMr2GwVzKD
eXvxDIrbRZL9lmbx+c+bbV0MWcisz5sfAdrHKX/CPYl4EK+tbynFHN52ytNucSX/
hHtVXjj75c2sid6/limjOEXonKVx/aQq+W6GRH5yVZIFPshibkgBdDvZTbp7rK/q
IbGWrbFQichWtU9wVaoCkEshUP8G2DwbauXRtdbd5x/eaCOzFncLTaf2b3OhgIgH
aN2/BdXawIIDuXFwAHo4IVnrJDaHbj5qzDdUVN2M9BsGT4PjvyFuRT8Tnxmz6Qji
o0Jsja0mABTnpC4tcjwkHPVQ7U7XluvfvgS4rdy/A/bVfNKXgsFnZSsfi2olau9F
pABqsKYvhkclU5UiETA7rRA52leGdHjmu5JVIjMghleqcjviCRxnQGs34Sa9Ftnq
l0yDKAlczNeKdy4mzXNflF9ChIrjN+R3mM/wEfj3Y1jFJn/7Pck0/5HKDP/j3lag
k2SFsPZT2Uyg3rcysE/lAynKC8RU1pQupFWhf4sAJqeM//nAw3jndz2JG5gDHoJs
lBsceYauYiQQsfeJXVtir0KLC3q2OOLykGwW6DG4GOSSDuOuX2iFy4e3392JqizA
NqbM+IwR/a5VDlvcnJczGuByYdxuTTjVZzkmcZt4kNoxSKu4Ynwd8bPrHocTGNjQ
ZJ8tw8NpCeoIDXBMUN8zKGmEcpg5rlBYbMDdD7Byn3YQgkksrOE9hFjyH/MsZCuM
HmyXy7TFrWTUG5sbQDJfiD8iLM1qJHz3AwjIhitOh/trdR7adyT6WNRhyvnYZwP4
Cn4X/dCyifpRnkk20qCVltM6+j7edbMTee0591x0R5xdrs+IWLGWFwqdrm1MnLGF
dapDH/NJCOqmkq7luNnEsJmMzdFvYte5fj57hvMP1WzM22RdM9x9QjDdEt2cm+4v
05/QdnDacqdAtLAfHxviPSbFTEx8N6yBPUzl9Kl4SICLZLW58FJ2kVyYKeZewhe1
R8ug/GYX4xXyilx5OnsZ6hQLloV74lFnBD+9hL31sM/AqkTVa/qfpdLY5dmgaeHt
UEGMgCSGZmxvRQ4m8HnU+XAKjanKTQ5cU3ylRU+Z+Y0e8UxNJcvMGOTRyMHHLBbf
FbfnQAxxPX9j03Jd1vBYt05t0CzI1sS1gCMWPXt3XpunadituwwUF2yQnxnFKZzX
StsYvK7Kb6lx8VJNrZShgqP4teO4qUDGRs/y2z729ytng4Us0CGg5nosm572TzF+
4rNzxU6rkeJFzPuFk4sYo93AVSy0x2mj1AbmkybAJtK1i4HIV7KUIkIiYMhOAiT2
7i65ZyLEO1kylS38EJ+aQbFswzJlAFcfWuYHGu1aqDo9Atm8AggI5yUdSSyLMttC
TB5sFqzayWMlCLFt/F++IH/ifKr0qZMjMKrc2+0pNlPGuhZG0BzPZRZ80uvrQ6gI
W9fJDjVf7/TjN1P9BpQMWhz+0CsAjY99PFHmN5qYCkDgCFr9Hz5lDm/fKHuVr922
/r+gxdLgINGcHGYrnk5ZAwm1cbDTBuWXgeusBFhuXX/ElnE674TIG4ZV08mvntjp
ObBFGVqn2+swQeHSxYooMcgJ+PawYxHLD6FjMopSjeBMwUcWsYFmGuiEMW0n/nbY
sn5X7lbMOr+kaI8h79jn0nzZ2gGiA3mYMMJUncIVOqj7HiVi4HykkYtX8klQ7GFJ
LoPe2EzcwrlFtX/GUm8zAJlOqdz7dFKa+YQ619rEhzYSZeWQumEAtw+nvt3m2XV+
w20epKuOj9wlX7JrK1zPyt/ZPx7GkLPEQ2HKJNZ9uPCp/1qaK4y0i9khLxmAcrUM
y558hG4EduBvte+nCwrKt47kkhcMLEOx+jJ7Rnqak2IQSAKHYSoYEn6SGTwKt6xd
LVTy6hUG+1E7GdnXVtRIvltit1nzwd4wDIbUztnYcIV6P3j3n0uQbNICumbU90kX
HG5b7UK0w1SuRatzgGjX6OiSWovf3sqjt95Dy57SuAB+rbdOCM7cVJffpDjRHrs3
ezc56WbPUHbCrlXzAck5p2RvNjUNjL5y/AByXouc4Rli2EwmvwclkVSkOxYjYWyK
Lk0xfLc4yFVX78XMd5gNhAsIBYlw5IHaN4a6kkIJWOOk27HcLhN0p4E3rciKzgVc
pMS2g2na/Q0xDV6PAu2iPWoHufhP8lZjTjZLBhhfBssghKUXS3ULzfH4MiOeTTuT
ftkDwHw+4Uetw1yJLqA+NDNlhUwvRFWrBd3y4dlHdEQqm7vSRYAjILWLiVJu0Ktd
Ov0lr7vlyAEX9RzGM05Clqccx+xBhuID/DLCNbz09MAQGKF49ooTBmDUNrHLTb4M
tHsv0PZv2W/skF3n0I48wwSmIIM7iZw4my1DqVBbAvfgtGFD9Alm+4WNDwKSVg5b
1Baj8NjKz6qquCgvhbpjONaVnGWX+UZnOI4Zjim+jaEPXtj3H71GJBhIiE3FLu0C
wj9uMNTnFs3HC/hVugmBVYhhhciItPm86BSjp1y3z6Ts6HTXOUYkKrCiDtZATy3q
hT4FkP9Ira9VGEjpYsrpLg5oKZ8/CRyQ6rCfKgbX1kT9OVg9KMH6gudOt2vAMD1i
WIroLOU4i3WNajqk9J4EEpUGtnCJdNIT1U+mkajO3PyQb6FMf0UEfMjpqTuac+CK
ny4Z8kHOKWDFFsNMTE7yDcOS8tKP65pRhlFUPa1Tlp16EEHGFc7UJfKXXr5YRKlK
0G2p0XD8ruObHbvA6jADz/y1SYlaZ+QfaNxijalMUhkimGnr3hCT5TnpWM7Z0hcz
5reqXGk8+r3ffiKjbNBMuReys/6v79HCj+rW1ypr881TM8TvSu9BUEmXEE/V17Sq
lKFKIygyewYNQrfupC6/wbsTfMXiNn5fDwojDgmZAw5Q7I+CjT0kcQ/s3uSTeSxB
TlfTlgFxwowFi5TVPurr6e7bobc115EuHFimeRwbqoKPhm+UDd1vFb/dFSxF55RA
IkbTsjmFd8Z8lYRX4tv/UzUZhGs+88OVftssmyUe/a2mLlZoC3JGqI9yk0k2njya
pFrAhCz/cl8rDOdXktowaQG4w2xzPT+z09w4VNGf0Nb7fjVkueg4ApyspSrpEom1
jEH6/uvpFAladg1mdtQbjV+WtHCP5LDuMmIPvgRBoakq7dxSBTjUcxirvTquQkmM
Km2BCX6HXVvPy58vCdasTYQBYx73QSa+JkNla7fmtEmqMrdDMDh2DQ4wAmndjUWj
urjjXPAatv6Pspy/B/dCsLkXJNJarHNO8ovK19Nfc+g+nTQ28CgjYG5YDtdDdaob
c7mM9EvOc2Mogsyeag6EbrePLZ16di/rBAwcgIFyBuBm/ZMAd3TRAWHpjauXl3IX
0zAiNKMuHR7tcak75ZgDPop7pJye59mfVTr1Q9LdJY6TaumwdJfXg2otKSQSv3Xw
y6hBbpIZnHV0w9ummkoN8AViKvUuN+q4zA/DJk2W1ld0nCadMhBjTWKg3MzINp02
lrML5eNlf3w3BfuS1MxX5+emYnWpf/fAFk4YkrZpch0axapMTsu2tlr4IbLYRvCk
LqnHeqGRNM/VZZT4pEL/C/X8g3IM0BDlxnA+Otma+VtcibMJERikuxXb9IoLH41I
QhTBoN4aGm4j9HY2lB8Zc2xXFcNu+p/D+7/hyJk2cuA3LpULcE/iUTBbF6PbPRRM
aOyBfFSmh6+t0KXGEkWh2t1wS5Vvg3IaJd+FcdsPTmPGY/9PXLJ4K302eFV+28+1
PceQ0KV7ihODaPBBtgMLLOU2FbAahoXNgtUme73Qfto058859+YTZbMi4d235Vmp
2+ftln6iyqO7CTSx5ZqBSj3Kilnv6t6iNKzv8G+rcL4onMIiXFSHBa/hYQxJukQX
LnkRK8RNnaqHzBs1oDGUp4I5P7IEyMSFH7gA/sMeI/YA8KeIFiKBIn4cfrtyAY/m
aNX9ekri/nxVjrOUsXXsrJ1cklUAyKPgSW30kDIVr7NdWSXDR0pKF9xRryE8cG5h
vmNARAuDydPghHHCrsp+WQtnCHzdiNxF5+HSLRbSIfnqcPtwqpE+RZno5LGM35lD
qS7yRNwb6wPYMpvy5y9jZDCX6+0hom1UxP/i6lZx9ppHftH0ubG929NnF9qypitk
aW5oB/cptJRXQlDy1nEWrqdd1Md41+QRm1aiPcYsAZ+MVU/6JMHjwpECXC/2b+17
957qemQFylLJB63EtH/pEqZZKAnVOKkf7EZulzlqAZzbITIGiUS5ngguEceuSjfm
pyaCOoLn5Cm4bUnjwSSSg8sQaAk3LvmKbzFyknIx18IgVRNjuKvzSr37Ap4pJThi
GkC4OIMb4I3LY5vnydwelCes47Q5XqK2BVHky0YMjr3O18ZEZkljaVmgz1c1IIkk
IPN9ZtNK4bFgmiXKlNkhwl7QGITQ2p4nurEQjJuWaqk3INUjVd/I2MzGj3tfIDvI
mjCVsdA86jxcy5enG9Qzu86e3vAM0zBXzRKWRsFx0f1c6WFikQQN8x1/68wxueul
nlGtSVG7wl2lWanOtETJZ9+WT7UQf67N0cimuHF6U1bkCHF7gl8IM4rhW2n1yenN
GrWq+Ca4QGx8OLJ6bCYk2fDrBRm5T0v+cKt7zWQNp72tvo3wxZzlVgqgLYOPVDl5
sbleTkWOxI2DQQ+lTpH+zyISL8suLHiVgZa0cWwvgvHFb7fACStlPU47Z6wZB4X1
5XmWlW4iO5PbrtT7RDqjM1Ht8qevcs0nDU1BduuO4mKawYn4I5PUupBCvSyG4Sq0
HK0M0bp6rDwFm9JeXcv6H+xBz+IISzibQiprygLcS15m1y1d7M3I0nQ070C/ATqN
NGywGndOAsuq1sUtuJFo6sE1rxv3wCJyUJprnFd/oPlSwakofeIWB+SmqZqa2UeM
rIvVgpNvNuRGaJjLzuZZ590ykqUKwE9OP9NyqRl/pYyG6F6sbZ6/D1HQkSItQdNW
6gsng1c+MUBSNNXJZ70IQraxZXZyGUGpuSc2NBWjirNxsz0PPV9jMI/FnHT3x28P
3kiaoFEt1Jql8jcXjdQKs9oHoQAERa7DeJ3qXSbBTUY0Xl9P8R9PH/lY6HNwknmi
6pRrujpHf2j8a5W4NUWM5UslzFKV0WVgwPzAx6TGRlvo8wYbQciUFSuHoYq6I9Xj
X3OWMWdz6bnXG7i0Rx2J7+lMydd99cf4I5RDXQbSIm6CFl/z6QuBSu6g5RCgGBmc
Pb0OLMW6ZlwRNj/q97YFPIqih1+gPWQmCkx6MM5Sofb43QWVHN78hPSvSXfTWQ17
VZDlupIALQ/yiKhmCzF3oyln46u6wa6SHz0cOQ8ep4tqeHMsuTqZg6ws+eveyqrl
Q7Q7QPmkm5Y5NVO48s5n0pOBHvoVoXQcA9VsFqDxGKUO6tVbQH/5TZoJWdzfc8CR
zOefNDwfjUxRrxhv6ZxazEFHBpu/V50ngwhDmobbVhdmen/staVoEj4ay251+j3J
0cQz+wkgPI2qbAy+DkL2vmocdB5USdQk9w+aNHdQWoi68d8ItiMWfgMAhVd1hK/V
lPRBWw5smPUELXE13K82AvXhJTG85+DfbSLysBoS7mQ+DQXLiMZhOzeyIVDutg/i
HZkEus/68XmhGqLt3KzowYreFOe5w1WthebelSql9W3G5KOJ/16oYtvV9hnE54No
/L6XEX4ubHhgpqUbupE2+nERBvdmTpqiLGJ6pZN5EublDbngSWY32+35a7a7xDex
qi0aquZZAKTK8SXpWzbfZxLN2vevxCKnXzw/2oXvHWBLlBpyZx8HsRn/pHS+RkaL
75PcIdbnhJ+o7DVkyroFrbHVtqETIjVclynk50jUTPDqKEiaZ+KtJQJb1ThnLDmI
CjzZ9HdNI5C8n++Jl+9KyN5K8GuJi1l9P0cAsi8Y+n0MiSxuy4kE3IVqR0ZIl1eG
SB/lluuxAbGUvsGUWRw98M0iTk/wWx37vv2XqTmbFooGiVt6loUzRuRTqxsyBUns
F5kUTvPGMOZ4S91v9WA8v6kfs1tNTnYPLBdAdNwVaQO5uhkE2GeAjb0e2CPWHOVE
VBWpf+UzOTMDCC+s2phKG0MoCwCB8ms4lUqzV/cmlv1aOw2/EEPX1yhOseSePM+Z
JRBmWhx3BWJYnrkctt7OmWi9NgUz3EyYdEqUPWKoX/Q0AJVekpHb1NcRhqH/4MyU
FA4unnLJNoRC++PE+xbcX0Vw00JaJIHmat8jNGcxtkZpI0MyLifsvRodNPaUtRxr
tsdI3U8+60aHD15URS92UgiD6K0IsW7D1/HEc6OF3X4xJOoSj4ar1XCy0//5xuS0
A75QZI0UiJS6sbM9hPQCgY/r2pr450F3gY0rqqjsYlSvusNu+1Hm06ZBYemlB1vI
wLMXdSj3oqtsDoOeesHqUc2Zhe0ld5bnHJGL0qj8D3iAU9WIH0ry4D4rC50uPv+k
0ZfHTiR7jvLuY1QmdRQJDCInPfEEiYhAInnSyfSvM6MLVe8mY6ev2BWEQV/iBATG
7GqxgZWwvab8AVlIDOQ88ZW1ENUuRH37hIvlMtciI8hcqB5ZtDrTiltj1lNVbXBS
u0UiBc5Oo30B3JxiP8n9rc5stD9GAb6i30uL/VIdb0li2qen2ipOBuq9FeHTjR5P
euzyJIEdo8g5urRQ9lMh/s2uZNRIB5ymA54H9jfnWdwpc/INO7ekU8GQ7oblVwFN
+LkP8jhHOZASzEPSWtIECu0sK9o9N1gXTel6s2a3dPChmPolIyVfMncZy6s4Nfan
4SmIr6whDGvIy75jIJOrIRfYTlaTIFeN5/n2TagJeb1gLOwtTpxZTV5bqowVgFz5
W7GSJw31WlOFfVmxrVmCyP+5v3bdxGq6Zp/zDNLvgDhx+Fwkxi9R3RC0iIIOWp4l
8dsreAryggHKbbNgaF1RPI1ZfT3GUXVHb6TzgtxDjeXiovW6kkTdDXAsbjcnO7hv
ID/fZvEpBYSeJJ3BzV7tNiHPORl+84oGjWFBFTFvFR3kz6wzv17WHEsWEsW7K3Id
eOOihPmh15852i6LhFhzpsxr6McbDU7DKKJLTcBFZUUuCGo0j9VgRPYwDzlY629E
g479A3THFUJhKa9+E0Wx8745NKaJPgp2gr2DxO279mjdJioI8WCgJKpKfFKz9/2c
aHil8Ck+UEPCIEdYbFWh6Hw/URwhYExBtsh6TUk/zeF2V2vP8XY6DqGdsjMXx7Fx
oqO27wVvd4c83OPp9uh62o8LlC3tnu7xB1bwllU8vLl7tuPnP3wEO6KxY0V98IE4
U0BZipjrciTq8PTidZTXeucojMEhKR7EvV7eo5ypcsqoh41ZhXIuyGT7MVF6hIcb
Inf6Y/XDxYh/rEv0INBO5CAE5brUzR/zwJnZly5ASj/HpYq+EtfH1nVQ+WdpUoqb
bqkeqAherB6+CVCy4GUs86Ee7A8X9Ef9OEodpybkPbtN31xuze2zKjFp67WxFMPg
rcpXKmGQJjP8UA4t0UWSihpocXXeq7UX0UaPOojQh/uMiv33lwvGpnvvnN21DW7Z
YYvQgITq0UpjDyBVFUbsUqFFdirmU9Lq6Zjel1CNBaAsf5D1dSVGhRvwJTzcjYx6
V+rdpnyxE16aBsZ5GBddQmvgqDHK1lBRoHjfwnGpo7X9W/4DzaM5AVmruUg4Z3x9
mZRT0lK6jx84uXsIo++698hodLH/3aM/l3m1jHaHmmeLcV1MweW2u6CvVx2lg+X4
IyO/RA3hK+V8qFMYh9NEDqnTZzSH1lT6wUa14FexCPVDNhKe48LUJ1TQ+3mDLDCr
XEQ+rC4F8CG8tbvFq2uHOkTh/njxOi2H08guh23x1KZCAAkCylNGmDxk769WfTXv
jA/oB/ls//3ARhhnYXobPljuqazvAtMALZGE/0GCwUoeSVRBOgNacUup2IlVS5/i
yiYyBpfibqp+Ys3RwMrLXNibPr1L3Hh12dI/vEFzQs3zBROHq7OvJpgvRJ1dZtGC
PbkCdOwpSSojuasMItIB5PEDw9vApsRn+F204TtEXQT3sYQ2s9gaG/XDc9wwosF6
tpzZ016lvZg9a3SLCOPze1Xgf5zyEzQ69/4SvT9/AZG3ngweGFpaPOKtE2gG/9Bx
uQL7oja28bWqrPMRyrtHgbwDPtJetQqOy0PmDKQYzN/jOGPY9nXV1QqnXVGhEidI
teoG8JAf2Esfj4pCHJpeOm7OMewv3w1848Fqo5DZQmuzhFA2Of9BqTsFC40whzE5
LCQ9MaX9O3iQYJEWr7f+89vKZls2VvrNqGFKGgBR/jiZ06PpGmEd2bQDPdAfcp/s
ucwkQvBgZOmhWWJ5npdr/6IW8BWg15j9nyoU+TqUyhuvVBYgb5ZIMnQFJ+AHlVDX
ljPyvO+bYrzHX9WN+CvNYVrTndiUmUQPWAW+KWZwwY5TvdL0KpXV3kiOlLn71FdC
M5YA2Sm4joGnEH4FNZpjJk/E12hUk6lMtvZrBcbywcDUEvVLxBioZO5d7XE7SZtV
/YO330IFGl7oiYQiLIbU6glYXDQfGpHNmarvtcah/OnkSf6vFHucZw9rKH2CrwR5
uXcKQzLEl7l8Q1m5KVb9v97qs643Pmzs6htz9Liu+AHY70r9LMJC6Jama3tAP9e2
A+05TDKx9hbFWk61k6nfQrURCKCBt1fuetieF0HZ7HNPiv4tC7TYE2qnKkeqVDqP
2zhPrWie4PAFWB7Z3hSrv+7T1heo33RYsy7WffeNOwPCIOgEvOXZn/tse4lSXmai
CVSmC/GVaswDruDEEL/66WCwCbyiEpo4XMDUvP5LnysC3K1DfwTh7ctzLEYLYGrE
ndtiTkLmQc7DfdIVKieYbeybtkRukbpQYjpKmjAZubLONL1Lk036A1HJ1V/OYlyw
5FBd6IVGnJIZRGkAdKYYkMDZbK5l+Hb2KE09zUxrrE9kMPdkyKkk5Lg5iGkmwB9F
plYiI583vN2luTeO4YNHOZkydWkk+jzRQiCOdpy+0sGseMPpuelZg6kDu/Fa6AKr
ZczahFRUwPXKXeT7z7UAdPrPJ5Dfv7Nmvm9aVSfhYNjp2FlalfCjg6oFVRJHhb7S
lTFwVrFFoAD85WH/otLwWMOFepwM3DPe5OoWNTnCoSEwTYeUVgip8TOHzMFSOisM
irX+5kibJJJHhrlrOzbJ9BJtKna9HXUUyPGJ89GO9T84W1j7W25moC5m5rq+GpC4
mZjNSN5YLUU5HEv0mQfWuRyZ9QZ81N6Og4XGTaT2C8flXzRhc447e0R++Tc3W+Z7
JBEePTtZy5B0JFMTUDG8VqgcxYK6hs2YhCBjEGGRibHQpHWjET3VhMyme7wWWfwI
vZyS2J4kuzCvP7jFuXkVL7JZZ3/UaA//QXwWxrFST4gufXxpWo/VPD2XLLaMTz3J
glzPStbc9cPZMY/7dDar4rziJNw8nZw5Ji0nZnTVS+tDGdQ3tha1cTJ11O7TV7sN
UxljByuVvMbhfaaioHUAKYT329ZP+YpZTjgtEoG2w/6k0aKXBVbCUoKTFEeBlD0Y
HXX2Dclg+TVdtL2ihVQqmVhAhaG2wU0n/mvRpVjfQqfAqZc1x9O13g63B5d3Xg2p
rm6a3fstdSoFCPPuLHNhcGldnAw5RLF1DyUDkYcq73uSINYDiddVRMvJdvwGNOkU
Av5/cIyMFLNlKDA9aRrNf2wqbO3vdTcIvMVSp8u5TllunRlt2I+ump2KqvBeO+2H
IRc7jMth1bBITObG3rsC7xMhxHvbQTzLoGmXBRS1wbZUgA9SoWhC+zHOAoNm5jrA
PV97Jj+133ngAZBW+/vlzAJhtysunsS6sxS5lwW3+u5y0josgdeB+tnv4vCHk5Dy
DajBvhcMOMfu91PNAvgHR2EEKLkyB2mLiAvYFeFHR4g9ykXQeBL1nIJta43s00Q7
vpbcyryRKfFmxbNNIXeTh6GP50Hbakx1znqUz3rITkHjwiEjXJgKRzGunuPsgWFo
CodAktRsT/qonwk++PHgzhUW7cD2mHyiWJjsmcrl3LxpXAnM8PonMo5VPubQLMxw
kMTZRU7JLNcX26JRmpO8HfpdVy6/EE1t2J2168ays8yHwxB9ws8g/Qa4qLAykBNw
zJ/ulxlN1IStZ1wMupn3SCD5wh9xgFiE0fEJuOUuZiLgu7n/Ioho1VVcWZoziISi
AgRRXYoLM24+M6Dku3tboG1Ix1jYI/C2QSsW0tfysvmEPKOXlYHRrg63q/HAyyJT
lcBXsaAiA2FBpA6yCyvqxm/EowQ5fG0g58YzrfVt8rtMRsLlgF20Cnm0vsyeQ6XA
Q+Xa5Cg2VToOmhq1+6288t8EJG8FJu7hhAW+JssX7zi0AWsiXFITya3L+ynSQ90q
NykFRREfbVH7OI45/M8+PzBMSl7Nv/k84l5WVKdLKqsGE/c9Yhy5VRz5A0bllleZ
YTaToNig5oov/V4V61chvo+qWpfr0+aRi7JHvjZ2qqqNYsR4ljC6D080vhUIQvP5
NMmDVnR093PyvSzexzWJIMM5Yra0Mv/CMS9NXGNFE4bbOh5OBlv6tMl7jIetyRLT
3DXN08dR48Oq9a+61PQUt76lmBgiYN8ytZzwlHnuBXeax0Yn0WqRCFcfaIRS81nS
UTxQaWnTQZ9DjqO8fnB+gq20LTJZMVCKfF+3P46nzQVmU9Pg6Ye6J1SKjeUtpEKc
TmY2F/jTLTelLxrjejRd932xfst3T6EqtI4HRRQm2aDyJecol63PATJR34t5sdHM
gt4KuFZIRYo3LSM0NLAiUB+E/DEtpV/b+e2XgcmBeifsMc0PNKEzjEhnjMOaS5Cl
tKIm3hvPhK3b5sLl8ZBLDVLgVWpAK5empdRKZuBVJkRUk7QsJqq1eUQKkJr2E1/y
4oUrH9RrWhcJTqCNvG+NeGVdHI7Wkip3/SS0dn+Q8mWAJ/hcG+rlKid+97lc+g2X
+3SFmT6BPbjRke6UC8qRlb7wYr4/eD5wph2S3tznU/F90iCj+uBftj8FCMgNgCkZ
Z4xGPrjBlDkutu0rgpuSZCc2OeOcHY+qFB2LdQQu7tgSJbTcAZ3Q8IKkGsgsOSZw
iyDLyQ826SoQaGP1oWSwlwSc6Ylz3T5+F6n4xe/3Cs6hAFrjJPDwlWqtGFtbGVn0
8i70coLb2TrqPoqjH3I9HME236bDVFHl//u/35i3rzNs3Grru+q0v3MSjxnyNF3Q
nyNB09A/tIyqlA9OcR7J+sm78jquFMnjTdmid85XGxx8JXRN7naUS3hBcWAeIwc4
sbeW2e5EVM2BE/qtdAbi4u3oZA0WNvA7Ipo1hQve7FiVywBLl4E+kKo0DdXOyeUd
vmTl1UCfWKArddiGpl0Pb8B6y85JLdORGgqvM4YOMzRuBBM2WnipS2iKCrxSC09a
xTmEsiM6Hx+okPd+IB8vNaKGNmXcHUYNd3PAOi1PTBxunLC0dKiZfDJGr7XLdZj0
tRSQMMBoOBx0qJSdIy03iynJukci0qCQhaTGQhPAfZ4AaSxyYiHIfnvKBj0JhjNt
nwfnQA+cA8KARXmJpJ3NWOY91FeUjy11XQFwXe1s0twYnCpCHBVgq7Od9DXIxnuk
hL1TU72Ecj5k0bqViSCnEvN7oCSPVV68weWBXUFiu2Et+YRDGcn3Q0KRoLaSTFIl
oodjOSqNpnCi51Ay4nRAZ9rJDtEs2i5Ww9ZrchK4R/AghqFAA2dLvRnl6mGS9kol
5866j4Nyn8VowmVwBZj0ZaiOQiECQ8mb6Q6NmEyWYw9pPdizRZZVCi72+5NdKjbo
bzYo07ft0bvsHHhwrvoPPMe+ltWyJ+OitYOQ/5HvzuzVGd6x6mqvMC3Mv5fVQq7e
emkCS68hM9cE7Wk2Goc8XA+I90SeCIy6qLXk+udSbW7+eX6jwKs6hZTyza7v/c1a
ql8H7NoM5btU01AEXCok7P1IVWA4KXNTd7Iapo0bWJtu/KGWFpo/rsuijraJK4HZ
Cr6L9gslogp2ENk6NglThfnNGlInWuhJo3db89ncC4U0YBD2ZlWq/ie2kT89PFpL
DSE3DyBwHFgTesABX4h/Uu3CMxYK3h7z4CpZVHTzBzFpNkC76lMOUHkKtrrlK+oq
nljpwrgzAqWnHiUJjv3BhnmiTQbBOci+cbqwkF7hWg3N0aMzk14X+V0JEtw7HWCy
HVS4Flt4h31cL+DiLdMv7KF4mZw1vucz2AP+lop5Wedsrr6hGk3BuRVNyXScLBy1
bzSK/m/Et+KFVfoiRT/jn9TzxKd9V5KtFX/o/kgr39PaFa5Uf2uylAple930WGUw
CjtJpJP/v+TExGj1kUy+8OD0fqVh2x8ugxvsmVyF7iIDzXthvPI/zLTiJWLYGs2P
W25tiCcM7fa5Jq3GVcDCoSdurBSmVWifmkxNMo1/HzP8H1ufEM+Oyy+yiKLuZjQA
x8O2WyO2Kf5trI3/VRz9aAnsA0Vow1BFKmqVozqdiDJS863cokBPi1EGY0n2saUG
VL062IbLZLjh4bgggvt3c1U7pCALNFM9cDIJqaKivavJFL6q/UnnuJr5qNTmr4z9
eT8NxmbLQ801B754Gv5dHwlaI75ZTZ/Je362P9iattmiP6CGiSfnh4I20RWvk4HK
FkYgZ66KT2F/7glO2yt3TwTf0w6iaNkOuyoRQkzvXTtrgGbeYNPvuiCU9W82w06I
541WgeCOuZr3gyUwMD/vgXBaH8p9QPfOPlAGpO60krm28We+ihqCkELCvrYvEW3n
NArIWA2on1xDiaAFsArfE+tlkboR1EsgcISIF8+QZHK6amTcuvMutpE/doTbMSS0
YGCef93Yff/6Gb0vmrU2WlOPpUdc8lBiXB3exaQw5PqV9ofmXRnZ58dWe+z20E/V
+LP4A9g6DbBEeye3jRQIs21yTjgDq6KBtS0lX445Y5k8S4rzfyxpFUMGCF+Itr/g
M1i6MB4wkRoPzDE5inio5eQUiOh1ei+IOC01KDtphO0U2SQjf6qq2dRHp0zJJXt5
xAoSst35v/W8LF+QWAZ1eRn0O4YCSxjeYPDBZT8ED5cEEjkEg9aZ3GMEjSTkJbId
w/jK6yyMLxpq8wbXdEyWZ28QOn7WiL5XnsY/q+7UrltsFasIrH22iJVi4wM8Qeg/
McJU7jsgoAuqHyIQ7FaPCip5EdfDUT4qA5twIzU5zO+r8E+Ual9i5u0FfCzbz1FJ
d96GrF5QqgjDcIafiJlFYCM/IEtMEVRXE67jutsyMAHhSDnD4UMThR14X1AOstSZ
eLPIOgCO4meeMHc7nnE9b93pWdSu+K+46ZoL+NROsZ+xZac73eapCDXXcOGSGpkL
rGSXg1LUWl6yzg03KEfrYXqEoZfzMPnyDa0XTnL0OWoe1LGM1yPD+jnEZ9ff3NCw
iIo1YlSVezJwKcdf04m1PK5UblPJWs+aIFdfDM11MW+O10L0tXVgxm9ckLcUkHHQ
FjMZBP6j+6Mt1E16VIcbq2z8Nmq7RQNtw4DdMkM57P18YKBeT9QWHyn2xnLeY8CI
M1U59hrWwLvXgTeuXYhg3SgLbO6oNEtJvwuCFPzaS5/1dLkMHaMFt5MbTJ9GsOsB
FvJNN2caXRGVpJDCy9506kiCsO6ZoeOpMdmS4GJBYR9ue0MsEbzAEVHV5Yl8thNz
Yo7dqmJxWfWdDsH0aM3e/rLgZMDyHvxFGkBKMWJXJn8R7LIuemWvCcpYR4G+oNlR
kov9583xTwwa4ICdiqm0JmKCkCksJUEbLCCsHWbDi0eSLuKraKyZe4zJP/KGpXmT
j//0h4XmnQwjK6NN3oNif4MDen2wZKt9Jl49Lrfqmlrr0cci42EF9O900WwxsRlB
CLyp5WJpKdd21cix2oWKa0ETl0s0lkETxd89flyz6zJizB8z9z+t9h6M/XD7TMlB
gAqef49sXnMp2L1tTPlSenZebbJGyhMtGqix4bNoZeudugRxI4PN44C0R9r8FE5N
CBwbqTNgaWZo949lKepFWRHXGrasCYnUSHWCQCeRTqSNLtaVqLEL9iAKKpnaeDs3
1qqMhSXi1sjDc6F8y7wzUHfGj0osrL3XI5VhkIkDpSsOcebcfAUx5H3hxEIHgMB8
liJiqrv6M+nrhsfSYuXwssmQxi85IgdyLJmZCAuaQ3pyDotor32i7aiNQgd/exRm
zCHfPqLyzLayoKTjWxxXp40V2L2nk0gtsP4jVDTixgwE+/phiISV6pwH4uO0+qHx
inA8lr1ZYAM0A9/N1LLvHI5XJZw/VBtwbVcA5u4LPXXFFohMZ3/bR6Quj8EpV8bE
cxGA82Wdig1UXZEu0NtNFhWyaaVOo/9xdOVXnnwPoUR3EqCosSiV8aBemPOpNbHW
ur6llmOCz6QFabubdVwxHebgyuHcemKBdyx3ZGOdmUAk2GI4a9U6c9GW8e09BZCu
l/g31QKhn6yF+cU91OAU3mlqnzIBQSMvz8brMK+9NYLR3I8L1byEuxmWWdL1AsYl
+eh515hf+lZWPxLD+NM24O5JIvssV9iA5usVUGojA4furzWgwtPlHGkX5O+SvRM+
+g5caoM1bwTYqsr6LsZm+xF7aXLu1uBDSLje26EU/ygPN4TIiD135Jl+yMAuob72
BQqCamuBQ7KowAKWSuSMZTzFOzF9MNhkiJa4daylq2tgmqMgegob0v6x6vhPvUNw
dYEz2zdzsfwupa2TUYIexdwuGGmlqmzGvxNFyqHzUR7G5II6On34OVdHK2yEtK/5
zrZpx1aEvZQUs6TdpJMo08yw0ag3b7rfA+mYmUTB1kMCGb7/IJ735p72VDzk+zh9
Rs+lBdrvNP5ptsxLZSYwW2mx48i37blF4I4OjFpUG4aJcFAZVKZRSQcv5lhU1OC/
q0kOU6v7X/Zj9EvtenSFVinTmup3juLwy129BG4yR6F53KM/nqgZlFLuH6nDzS+G
FTBCNvWjznN1rfJIPVlP1HqW7qiigz1eLPAgVnDlVsjNhf2qDu/ukaSG6R5h0836
XRms3nXx5Ji7urKzenDiSAkQa8b6fgsjKijFbgEBEKrWBo6RMns+e1wL7zYaw2Ve
gaMdzv9HRzU5Xo4hV06lStENtuDco0pH2x3GxWHOoMs+NbxBwhisi//V+6fc3C1/
RjC+/xMPxCrpwteg8ARQWvPiei8tEdDyBmV+r7xQ+p6PC2OyRVTPxJx/OENh7VOa
drZ4o/ANjAeBu9Gh9LsG3KnMXLkYQw9cGiYhQhUFryBpIT5FuWeSGQABfcc6bhIr
8zueRZbp8LZdX0osL8omZg4e9yL9e5ceVx87Q5wmV0cYqHxsyfjxNWDF9nFDbAOD
lUIZD8XMSTlEL28vxBx/dKvxVd9p9HGhbNA+74m5H3hSsgBqvepL8YpX30GiRT+U
u0cdaqHcBw0zi5C8bkUfObhARH0hmLZMKroA5YrF8lmDNIBQpVsKm6n45BEsUbB6
sX1fn71NR+Za0Z536yvpZ4TbKk/qS/bw94A7j9PZIeboueCc+3bAF8R+INMFgQ/z
XUyLx7GNkmCfcCAMA+4eemd90fr/PyVhTGp96ZE3BPcs0DrVWakZo/BuDLVHkB/T
Xg6ww9mamskp47rkakaJF4SBNfEo9sZWTXU3PJ9biJ9Yz6jpO/tj3M4YAVr0oiid
oeGYXVI8pWnJ2c0pYM2WfKcH55ZGCDRzBr6tTxoe7hJs8RuV1Dqn1Ct8pQ7MnPmV
2QWyxTiHjCL5yBjo10m5wePpP1A9feFxVuiONvqbbzmfXVf4WrT5/dLtFKLx9iWl
a2P1ZWEkhrgLz6gyKqJnl9QlbD5lHwBGUvQAOKBiD21fFStIGvQPV8L+HM1x/rhy
GnHGUkNafEwNXRk0hvOb7QFfl8hCL8T6BIBYk63vpu8YfiM91l3+kJzRS2rnkVTz
WCVdbbXVUIygdualDvFyVFGznV/ZSuVey2KXiPC8lONtmdfl0tUGe307zpi4Mq70
SElZfhxx7GYwS5oOi1LIJsCaCEAoJXrJdXQowW7uvKQFQ7dbXJRe0DZSNNFNAb8V
5qMgVcuE2cqpTxVvHpNYXwb8MznrrZa3DWKxE2A80OsK6mbsSDtkQCoRx+4oXy/U
F3bAnZ2IGB9XLJ9Hfabdhjhh++LyeeNXsamYK1pu4LtE3szISzTHFbx7WexHFsr6
iWbVrEfLcnT11SO4raCcNbZAnrwgwlaTiZQ1bg8iY7lmiilRb1eh7udjoiZQgRuG
xsOcnr6rC1PCeZAe5p0Wam1GVcpQF8OFhIDH8sgWnnsN7j0HbXnbxMXoDrycwBxf
BEHRjbWjEYPNBSKnC8RVK46HQskIFHixwoEvyn7DHSeIa9EX5LrL8beJd9d5ddqW
bafYwlk8n0Cu62eYAM0gguFEN1YhrhRH6PKzpKRoXdXWWIWgNNPphAWR4WUyiauG
ScbEZFSR2bRn0WazNYjWAmk4sA+gZsSdxXhGJhJFoAXnw2LADHlYagC4Nf2ZHXym
Bl+cfjE7PPpxrHCTXe1h05kH7mFUqYSSNUJvPYxZnVf93CsQdrkykprFvUNQ6Gki
NXbRC9xGq/pq6n/ZOtYhLHdPwIE9ahW07jHH5orfKEnRqg+v9bmII01Otrxh9bdd
UqPjbs5su3f5sSMG0B3hPVelvn3wyONm/uFxvXy3M1+arNkhJYKkJAZ/lTQL80o+
JlzreRO1odNmQSVI/Z6wQronDM8QTSCaRmgjfF0SduAV27NwW9CEOkRXrW1k33Wa
1/B5phKpflDfVaGWRNBa3zcYsOAepVCmjC840ocHusJwdvig5U94s6DtEaAoT8IE
3RaaVs8ny446iziJ/FbqYD4NGrQEb6boghS+88++u0cQP9K3vMOM6WaKYBtDMbGX
4ibjpz3j2fjrRnMBYkiToqJC+nGRgSAnTafQiI0R3FcOOQ2hBnkX/aX1+gydGtub
lf2sbUYW2I6yGYNfg6AHSspSUWU/M/dP9MlWRgb2kmMAO4NyTP3k+l5sMNLyBb2o
Nyucb4eli3JokcuzmRLBvNfbZNCkA9wLfuyv+di+BC/Cak9KFAoaTryhi03rkBni
tAYf36Dsyy9Wmz5Tw0YJ8pHalQR/q2k0/jjfrvPKAn13ecON5cA6zJcK057N2Jdt
sDRlDEtKjDZ9wpBHP+lCqs18QcsVqS4wcxo0W9ANg8nAB42u+oWFmbJtrlxGvJIO
EzJg9eDWMl0LwFYGocSqvfwunQXxX09oqRhF2UDoPdWnxbz9EjsdCbkiGdSpxKU7
Ukz2Sp2Fl+fUENGKPTnWbBUbcjtpd6oioN7x0JJZd1tf6uUp+49AIPzEARzTE24E
xLt43DhNYn6AiOAYjPrx+Mec3hXQgdqsLUqp6iPp+fkiOxNGiKIYBZ5RtBV/b2ch
5l1z1K1xVjHXC7HlpjNnMocA2Usbp3cZN6JyCv2ASDeELo/tRmQcSgRcgmIwfwUX
tmCWYfihJoNx2CVWAR/fxjUWSBr7vR6WAtwwp/GA/SYQriM8VezIoDIgAu2RVboo
4iLnHg8Qso18XuajlmuOivja9tjXKMHwZziZYhvxrbjqczxzCtET4zzARxNP9bkD
KCIdFnoSzUPvHzpKGkgfhfowkcPPeGSwQhUZh/39Yke9qMZl5Q6Hgaya4dIbV1S1
7wuQYIYOYf5El+w8EYo2854/bDXXadctUACHOVpV0klnxVpJlHg62/zqrHruWiY/
I42v33XVnFN8imuYFnzGERt5Dq8JO3GPJcsiiYnzUpQ4SIT61U7845sMpVo0ay60
Cjcdc/UIncgsTmJSa9YybtQWo/Tg9+iwSzkrhG/cvIPFrvM22taZl5qd1/00iGce
4NuPSWvx4PO+ABwEv/NJhCgw3KIhUJ7lcbXRV03zKKFRMFerEtf+bpLnLur3Zm3D
UOPTr8YK98Udln+5CChkcozCPazklEiV/FsZN5hKW5PYlLxdM5ALh8RyaNlbJsI3
sPpfi2lWPX8/0YMxsgBRZQTpiSjkLZKqvaMF96JNA/HTwTqj54I0DLkughkPaOup
v7CjqKBQ+V8iNzWmmwmo24P5AwsYflnZ7ZRXKF94GkHQX92yepJBP6jBkfDE4o5w
FL7+cp612yoXITIQInt+FMpKyt7wm3GPnBQDFd1aNcQYdbzderGn/9Ce6WcIcPtk
gNew7XsYzoHmKToSBOCg9DylFzcCuOcLbFWNztvTmf74pP00HPiVhUWxy4nZEK1w
U5iCJgi30Kwirt0kjax2eXQibQgAUkMLUY/AniSTjaMecL9cA2OTRnii+pxQTWtK
utVhMTedwUNWCj02YAHKdLiGDQjqS1/1hmuK7q3seBR9/Wdzk6qejnuutmjPc3WE
u3jDKMeuvpLedN6oE7N1iD1MP8J52AduFf+qnM0ThhA5C7EGQOZu6XT7JPrQOmuX
uZeJiK8N0WmvioHsQq9CM7cMsLYU0UKtZIsYc6PG02F4iDZghSK0Eyhgj+rW8ZLB
f89q1GCPO3ksEXRWPmaFMYFXM2odjPGPjVYEjH3tVDY/I4CAToS6bIg/zHVI/nET
Lo0u0OTOcKdgFMH18jX7Lb4YcSKMLWrcxLj8GEb7MN2sS06yOy2+J9gVqgpia8qI
Pi8dntIKxD4WVEgi/Z5Plq5q8ot48kTCbj3FXUjC1CjjKzLk6pMGzHxNNKpHYEUA
U1RQlAsHpZssOjKCmIDyVjxjhvqSPg6G5cBw0tTiFyGfdjrzEQ2B0njyK8vC3DND
xu3Lo7HFBWWNSXqGFGGlaFhlmu0UooGAJ22Uqb+EoLI6rxHxSbEFW3EYgjAhuCgf
kDBVPEnvIXLVYypto4+mwEEx/APWigUqK1EoE+oaoRn9GOcadv0glJ3y42n7F5SA
Q97kpeqP4b8JB5cxwU8/hNCMNtLsU6EBcNX+G1up+ewni9gH/V+G2yzaiBVjGYAA
em98/7wiY+WBV6ksguD+/+A/VqYZZ21PmVn1z93TDUXqHogSSryMnbvFR2s/+PU8
RquNPyH/7k8W4fkUPdwWnJTuN1Iulijh/F8OSU+5hmIDcypeNS/YkJ4bmQiG3ODd
dIwR4GysLzdP+iCozCAfQsfpLAgdiyEICPemj5kOB0ex+zqtrpDFi1OH8AiRHDB4
JtUYUEzKux5eFc8SpRbJtqjPOCMUZoObaVTLUvTmHiWkMj2ZH/s8Kdz1FlhXS3ny
HLy+NKNCJMa+7Qy9jiuSoA1+J3HkP1xF7T8+vZx/dm5SZtErbPu0yJF84+QtLi/f
QolUGC4axlhnSTBH9pEbHVkEq5avX+g7ynnm7hitKtGuU8nDEokyqMIla59HRqCq
IRR3GRlhANg94h6o1DBRQQ5JSW6Z3bRIGh5HfvGrAR4mMwnITDHoj4GMWAsuMCNo
puxnPw8qSn9Ehd8sPgnXvBpstBkp4iTv/A7kc9JP9Rii4Hvo2elrlX5OZeB+GAeF
Jg1Ng45CIG38YkDm9rKpLBv4NhW+lRSBNIWYBVJzGVG7PXSHcEss7FTfAb9oyCZP
eeExTytY3l625YB4vC8lmsZ3OvRsowsxZG8ZyvEyCbuYaftOecQ4Fd6RzqrECEMn
y8JyNz/pVPehW7imRKt+DeqwL9mVJEGGSjJ5pyWCm07CLUNPx+Y1AgM3TvpWQfua
uP/tgabiMI/Jy6tMRTIlw/fAJ36Q/qyqAvlaq+g0mqFwJpkoldITuzACwB67lo/H
aZ0YFEQi4yw3Kt8SFt/T3mD4lucehXZVHhPHA5+TzgDSrdnGnTn6F18JsNBbDrWV
o5OVGmYKGKEa3WuB2W4MUqPlOdp8k2D/osUNjoW7RiNB1yvZqCQrSvH533lqCOyx
G4MZGqCV3x5SPJly2gIA69kshRemmv/NM/nNaeE+5EeXpTmCyK0pYVsIspInjEgM
PQDZbPq9Lfc1GCS+OsFzmDhbhoWzz7iQN7DpPWE+n1ZaN3aFs0UygY45/YJxTmh1
TjhGtqETWA4pr9TvZEDHFvqU+EfhlZAF2u6BUaP1+60g6nIyoLfQznHwoRN93g32
CcteUxN3OWWqrVoTDMU5Fw6zLJ7JbkyqGcXc7Wach8S+JAtpKG/7CGO6QJswVR/M
9r6lyPYu8ROvwoTwIzIy3CqtACaw4WD+MKzq82ZDmUm8pXhx9IvRJOR6+YXW/DSN
Qgs+OBRYAcRqhhMFK6CNDCdadDTWgepOlwJTRA99No3oiqk8aDXffu2M/MRotKTD
/w8xEhMFQbo0MFgaQa4oVCA6u4MKKPMQdckBuvnLYk32oAVFqj5ZmbIz1JGuwYkN
QuyMu2D8D/6VBvYi4Rd8cTOUbXX889FQx8SvZLHaEK9K/qW+m9sBgiwhp/zSEFQb
bZbnrIFUJNGWQ2cu+S52Gz7oKnT74cH6zjru2KGigIIiESlyt3s/jR3g9AyTvwgn
h1KZfhCi0ZfG+9vVnzhZ8LZ9Kt82QHB7dEGBCzTJcyc993njOnAL1Xbc4+8NFzRJ
w4FQ869SxiXeOqNnaDPCZplRwutv5OT/MZ2lfxrNFpt7nWZTH0P4uvRfJacBuU1m
R7hQRx/Co/upta0ApXobi45k22GdY/23QuYxGZfr+kwpGpgQBKlY9Jh3mbnXaFKG
SCeMV3g6WUYUtQqpH93FjS5sJ38vov1yRIKpXbeE7gRW2qR6PKJLmySCRN5THPMM
lnUmUBsOaDpwQ1WqDxFSt2KPv+CFd4D1dqL7O+HCDXPfA3L4rxm+jEwBptW4OcpT
sUnAR+Mn+R2z0AvWrv6GNRP36MHxnfcR4S6akV2zO+hL2NroX2fdc9EUwwLeKQHN
7rumnzzxlfBzkjyhhJpNX2Mlq12pRggzOku6NH5VUjxxf0lg+2cOGPS7lIACykSh
oa30q5EA/k1aRTr7/AiX+rlsk7xtM8ol3D8vzb95cMo/NAR6Bn8h6ncT5sGp0E7A
2iGWw57szWfE7oefYs4Hq8VePyfBruYeXhhhSAuvlWAW6UDMsPA4Kx0H3ER43Fwr
QfsK2BVinTZgTuHKKEk0MGUO/B5VGkvS12VG0K1aL5/PQ4sS3WsAlY2YRStPfIsK
hqniRsDXT75kDCZvJIPGsjE4mqmhBmOp/iYRS12YL1NPfY2II4CdIMittUzjZ1xQ
B7p90fE3XJlt0vlF1Hr3GBEjDgZV1N7TQWAeCfuV2paIVXUm2Dn802TMqEvd8tS3
fnl4RvJysJY7wWzGrrfgG0M85xzc+4u5Y6ppZwxM1KMAdzoCekSvB6vBHIakI/D+
elZowbzPhMxQBu7Vy0i1SRAgRkbi5Z9ZoFMqG6FLBTG89aS0uYUWPLvZbbrpIOzn
1B3jf7HhRf+QVxmKf5BI65Lv4tey0UBWetXNQuMjdQ43ucB4IZrd79e7xo94B6s5
0XOhODrPxFxSLHpf6U+o0ZxCW6nElNYqqeD6GZAO1m4kx+/jPhyyLYRzRvbXWwpC
Zl14kfjorcHDhAB4y432YnM5Oae0yaFiGS0DNM3/XsjgUTCexnjsNDxYSXI21mDg
knEmaocjD2p0l8aN6dteAO8YtIvhN6ZJ1M/WQwKr9bwT5Q2jEc8Ryb6A1OxFJSNY
w/f1ZVy5/uh3M7K2vslSFbjR+a/ilNyaz6hSx72vqXCktk5Y328PbTnApTIhoE1A
vYKuU1zlK7Ohjr2m0t0b/rXtNnj8cT17lRMeqzoV+b9p1SLycHLPVlmeDu9tGjNy
YiMS6gA5KbrBjxkYpQYk0ZMtBeQuCiJmeY8Eyu8ciioOJP9sgGHH7vPwiy5UgKo2
87/kmoJaoph4wCk1Y7gCLIM4kI1tZZaccfi+P0YFkqJIWLwGTVP/sAuY1LPCnony
MXZQsfYN+QoR+L0qWNAM9A8e2z4cNYgXxouMRg0mmOqDksYiGx98tEAVelis4RLX
ZfuhSk7B23EAKPWRPKQC0BD/HjavW4Qm6F+x7ncJeQ8Xk6GxRiWootnAaCH0xqnX
C30+SznSIZvZYdBdBOcyIAXBXb1jI6eamDHBmGHPdQwqAYtTPFdfn1xVnN3WN/+d
3eIcVB0OPVk+oqxnRjSagbXx1ehF8WAdqKj38flVi/mPwLUJHfmEQAHO5gqLAc6J
aOUoSbTOBlWpvTI+PnxRgMlMCyaMRX9GKO15DVYrdtmeV0AxxnUDsLmHyWRqrzVL
EqaNmryJbPzk5RIQ+r7Kij6kvSEFsLPFs+x6q9bvnXhJ/hjFgrEOSQMJI7V817Mx
/5lTyo371ZIKm+F4JZqNYOG620y2M41MMBkvd+nyqROdBo3pYZwLSLI4lc2uQYZp
jEeeJilq/MPkj0XTobvgXiLAeVJi0b+fs/akkEP99oPyU7ePuPGr9/iJMIJJWbfY
cqWDs1AN/rMAtVQuhOeNCTEoRtG5sN0WIGIYh4Ury6duZlxbhCCAlHLo6dymVToA
RG7j+a074wZxfjXHzaWT/rtXdhZW/UbhdOMkLLGo7VUign5abeAXtq8ROHaYHoQS
+Dre5c05AJ5forkns9acbn3w0G9SqVnZymtrR2bQ+agcPyqXj9T9pW+jUXsyNWrT
Uoc+KNu1jG+JyMVQ7wiE1a6kotVE8g+Pson1MbWEAWAglSfRD1SfhgjHfSumGeRv
j6YkarZQEtgAsd9m2a+uefgieuCjZSolgZ4WmSZOAzCba2y3ZGcj4OZ1EqVm3+tK
A0yMBM8YygLIcFTJBR2rqquf6y4c/8L8gNnVHl+8UHmTlnjC3o3fDMgKMpHzZrRi
Suwex2uAfz4zycyQkhfuD1DDMo1AREllkv3i/w2ni6mLW5LIEF550/Txw6xUSc4y
Nz5LfFUUK2SZFGmgTUX8PLTS7v4CLW63/Udj0OlEXds1PCs5qhljsyZg1NyBjrQx
EG+P724KYi6OH/Vh19Hnhb8m7CuPITeWwG/408EN3Wl70749EXUud/EKb2IULGpf
tFHJqkvvTsv5ixASpq3iWVvCMA4VCAo8FFbOQ1XhJ9ucfsZYoDx0xh99/nBJyxZR
UmlQtMRf2NYltLa4j874ATrA1EiaJIiPfAmU9oqXVRXJMrSYP2n8+1bzj4o05r18
oKr1i5Jd59FleR0eO76v7ygXboBatmyWR04LktzzyJEmXKBDFJJGhdpJkAfEaVrf
fNFvd48c38xouWxadTtrxaIB2a3gdEziKe3sdo1Jal/uVXL0g4nxjmjgnZFjkPG5
nTK8VoabwF48bdLLeTWzalOQUyVC+aPkE6ZE0G9oXYVWUi0vyzdg7kHGbgtaKiWe
J90AAhCgq7C0Lm2WG+2jUvciBxIffY1xpcEoAz8qmaFsYoA8u/KQR5LzIwWT3c8P
wW8RZPi1j351jm+If473Kt27mpvncmLKrb7QeWObDVaYbcf9dN4V2174V2ilxV4B
g1bKfeD9xPCsuPLWdcqOcEdRjiXzM82m+PqZKMygumpiPiqaryVd0k+dqqXo8OmG
waXxQfKWIdtttuHfasTknCMMRiYMl6aey//yK36SzqWTOGwfzv59XI9Nys7tmsdu
kuxpUoPqwNZPuQ+zG17S2SzjCeyq79dtXjOQhslJ7V1DaYqDD09ALlKt5PSJoIIA
nw5ee88cxDYy/bnmUZswbpct4idawM5uJXPBwzsiFoswTbm2EdWqfbFAGn4zEdXa
1JRfW7pcRjHOMQCAoHscjcDEMiZ1YCC/vNQjZznP6qtINmt/rEQUpoxUPAncoViV
ENp+0s8ojF56Vf3mlx2rajpjPhxFmRAPMH2trNjunvMWDJxhP58J2MmEFFZMqmuQ
jV6L9jX1HeB+H7OGitoiozxhv91ZyaWB+XL8f5j89j//mojdyOARsauhPeChtj+9
TXM0UH48mlOehNjfPych1eTWL91EEh+NDaPqHBuVuYXixDtGy2sfKZgoBnX7pAUQ
bkyT4oLQL7Ql4YpLhJVkL+CpL7+s+9nVlCSXSzl8NZCfcuTOM92pX1Vvi7UCpcWF
iMNG071kIafKli9rzq8NOY/nucsenHUvJVp52l5xrSgxWT/Zv27O5NoKqn4JmNNB
5iv/Y+rX4rEU44lwi0nJMucTlXcV0LqyoS6bJIXtqU2G/VIS7xb8EfSAui0AAIXD
Izc5u7NzpP3E3TwKTqQkBvgVx2KCe2wfbSVZ+8uaidzb/J3/VAqmEgOSwFt3DA4E
TGRE6ik4+wayhfaTI1B7YdRnblTGbw3VZCuR4BPQa+FpUve6xaz8XOnn4Nn7tYQ0
wuu7rjtOK8/hgHsfXSZrBmWQp0uOT/Sm5Al4Fbshtvc2EEBh1ZvaiYUhJ0z2zBL7
yRBUUAImoS7CzW167cUGe7VPH17zEGWgBYTRrVPwXPQg4jmjoOh3pUV4JXm4ttxS
yttRLccGK3ETcpEPTKrMUY6uz6aZ1n3gjf55udZDSwY3MQ7jJL8MsBUr+vODyQxC
aA3H3nM5pH3BMsfGdWOfk43W5He3Qc3Y1oyr036N4A3xn70KAnjVcsFj6oDYu5NW
rW/iVuSjIJMyHt3Rt4Lr5Yfr6yE6Xjrd2zlBkPZqf18Zy9JcGKsVz8Hx6VH2OUav
oaFl7pwZYqO+vR+vQCpD5xCJX759T19hCTwjNbkF+XYl2PtcQLkIIT45AlJa32t0
C9mjRoGMzXt6++3UI3nla8Ie++fkXYMG1ng+waSOFZ1KmuTABLBnDa+6xzahbSCY
HVP2lKhO7bt74TTnlG58SWfAHCtIteFIfeaTaLZp2bsjhpkt5hr+6JBJNmIiXvHT
DQ2j/8REYAL6inn0M6FLhsFP8BVO8BVrr6C1POMAVNpcrQL7rllQiCzB8tPKLlRg
Nw+ozc96K5fvMyKRDuXzp8c6gQWR0oVToEBBHF5rUJgVUOyrX4/Z1zE8tzHM+40Q
TuR4vlavFPwXh7DA4ci2ZdNTJq/uGPUTpQIrkw25RjqdbKctaJ3xGa+UR73VdRUw
drHj4KJ7JzenQy3VP+7H1vNZK1fWWA45lQKm4bSZNEow/olIzdfr6UQ9TsL4vhB8
YEYNA2zZa6Wy/xBICvSiVjR3NiaN1X2KNxHye+6dWZ3frZy1fCVDhrj2tD5HG7C+
YBpT+GPoxzC8YhslzmcLlj5OLlA74dJ2rPt5+vNI9CQxZp9117jY4ysxdje6M49S
Vz7/Tx8eb3cQpb4K32QSHrAMPt+FI01d82upbwnhARYRdqd1n6qiTf4YSi1+1dSF
Xcsze9wm2qxZ+TcYOguMowX/n1SlmhQ4wy/uJSadsoAavjHEtkYPN90M2f1y1MKV
qNKPKU/fr9URTsxfqc5QuE4fXNzc9o4B2m5nxBHtEjonnd4etdqH2RsyViU+Mm8D
z+0nS+XWntRhydbhAxFY3cNSf2zlVB8H6iFfsBU7jqOfQRkLWyDWpaF6AM4uz1He
PBmrPAtRsOg00+mqtxBOy6GS50oFmKCIqdQZOYuofU+/w6emkFfKigHcJzrKILje
kEy/+7m5UZ1tSulJJp53NRlLZP0gv8APZya9IQirELxgE2S9PpsjW0yoRjtZjk3/
PfKTbeaBy6po67N5sSdyz8QIoP80mmzPhRJoL4a4Nwupi8QvE0/e5ki64VaYMqdx
Zz4Gm08FE3WXLJcK9+JjPz6YTTrgDv+stv4Ct0zfDHLnDyCJy64zacerI+RqscHI
Zm17+EdNBMi1c4FFlSruxR8wcEM49ORRYtGsaJkwVIjVHB+Lyh2kz7hmrrpjdpiM
FXUjxCD2eRqIGCoY3Xbsi6J5asoUMKwyQyWYKhnUCveevMe6vGAGVXFoBIB0yLST
cS0QjYm9jIvtF681Vi1u9WyaG+69EX5JBodjUsr/Xk+QMnG5c6rXubOt9fMZ80So
dKqTtif7DOzsxScLQyfdjWkmAQHwpulmK6U+eRVrEVflMDAyQLA+iXEu1A8LAA5W
BLxgGjUKoBhRpRbzYu7idigGrw0am4Ih7jDAc2iy28nOru7O+04gJzF2e+AV0nyy
VdKneV/TY1iwErFjIblnx+3V3TO6rrS22w8TNkOsT5qL5kJj5vOVlcMBUHD4rHcf
1Uc1ot86nWVSQG9rH8KYMIhScB9RRBuQ47KII3/xSRquSVi1gIOw4vRIpMNtlXh4
OTazrNOrug78+8VCNL7Sf8gZeCtmPdXBJCCMmvVOhrrTNcmkGYRQMyAgbmxn7vC5
ovOk6TfdfYwx6fqpuzGqmqzX+o0AZNTBtZKUqkIy13UoPh41+vdNzr8PIYbDpDUW
vyu0DAxEUUD1ktaLFWOadDrMK1FFc0era4YMo5yDAm/A1lFGbjI0y/KKZ8VWDyv6
4YSS5jzw2NWnmSS/fbHHj73i6gwkyZ4wRdS28Q6S/lZYC9KQEzghsrAovvIDImmk
K4rzxOrp2mnrM5DfIMrCRAUR2mTMRsdX2m085QquxrSDb3tcVKM41cPayD8956pY
v2N4g1xnxdBFr7FYXMCSGI+AHa0Ctqcv7REQrSg/J9zFM+/2pf6im+77SbMIgAPG
OQrlzZu0/BgKwHo28wC2jU3AY0lqLtL9Q30+bCcTb3vSngLBo5ZXhoCf/FzcNp6H
tqEWOfJs3KlHRqzETizUT2GzGflyZCjyKqNjbZOw1ONuwrC+BzeFwmE92cwWaMSI
mOWaq8VxUH6mY2EyMFVXxyl7IzvKO343t8lBgSiN2QFkMJ1Rc/eCayHgpc9oLWs8
5rqPKpVmCJyyEWiUq0/v04OV8r9wXeWDPrKWSjc1ulicy8OATH3Ly/9DcvdegoDz
iK+yHEa3vm4qTlFTOoX57mj7x0TSPxBl4R6AJmRePMLFSv6XFN+CPa74/OlvVXCE
VTORKSdyYl0LEpAR9biqPQXRdc2ejw9rx4ckfQb4a9OO+x6tq1mVFwmXMhPq5owu
SwE8AGrDIadf5Y//+9OXR5C2PubQvb3ut/aNleVf0E5dwaER07GOR6TnUDOUC2/8
pg/Td0TqwBdWvr56zr/ZRhuu/ce4oDJLWxiKuBhdju4yUpoHF4enoZEpi7g+bAeh
KbCJlxPcGRU/0zHM6rMHiXqUnskYPwWw6+tLvqaYZnJw5Z6Z4rCsRQ2goAQ9bXBz
bdw4NEm06WnwdnuKKYePshHiisQZNTX673/rySm4JJG46MP8stFxw3EByw6V+VXC
siSlZIU/NAB2sCJU3zjoZuoLiRJ7rx3DF/NwwViyDFQhwHM8+trbGrNQtww4Etyf
TwOH/JsjZQ3QhRPEQ95H0Tn69TdU7l8bfLMpzlbVtgGff2WnO8fipeFJ+Hd6tgew
qOWDBftksLrFT6AMfUD080sdCuRMnkGxV/ucXZN2G9waefo9j1MeyJC0uJHCmnBe
raVgAjV+XP1dktv3NG77YliGJz6PcaU60ygGk92eNfOvRGsZjktkAD2lAHCK0Vuw
V1x3L9CD5GEyXjXZ07eFTyjElZRSXVREUzExedPcKqRtXaIATecH81BjjXZdQsy9
hWOtwl/FPVi/bW1jbicedZ0+xw7VZKk44jrIFNLBPXPPEnZlYnboyyCsA32x1j8C
zkjFjm9g6HJ0BNqhcVptopQXuzk7b7aR2G6mhkzIxrMMeT/TqPcsRVBKpfMRsV8i
jBuJ3lvC1MZVE+h5AGYQX9fxZXKR9VAhmNvKg0dpx0y99fyMpQiV7W9UhUjDqAWM
NroeynRCzXWdIHuO5rAvbNdKEtkq4lKX8dV1KbrTCxMbitHvx0NlfWr5sFilPyoL
6irGYrzkKwMzQqxHboi1GDNv20vgDHl/X+byBLhYmDP1alofEYRaP3/dpeWxJMws
SlfIMq61kDVFFBS4OtpnsNs8puajFRWBPkN4cTNBA7yZaphlIrJFiAvRugpMZ+0c
huy0vaSqoyRyTDXe85Y+BSlbpJ1qHhONwVU5Zd8WZwqIgfLuLmzlAPKhYr+oeJVv
J8+/Z3zBfVuJkg/2se31n2HsphZxpzp+zQhRBXtJPTJ6ys8eyJkvaioUWF1O3eJJ
ueA+c0NBrltiUzsl0kOitPeFH98anGiTpugxjWgf+kxeyzcmlWImhoLoOox3z8CO
ZabvTsFFBFozbhFrgfonpzAz9eMtS0dKFXC2+7Wt8AE3CjGKRGOUkbnwi0ArUFHo
3ER+BMfhDAAmJ8CRFlewaPWxyPlwDPWfafMynWuhNAX8pa6i2RE5Aq/F0SCopBQk
kCqNrUJwF9wSX3gXJ1qMO5c8eN7ftdijyfPdUMcKVFXa3MvJAlTzIL46fbjSuTJC
3vNZf8KoVMy/YdooBU01BumDH28oN0WoRFmDYBCYX+HZBAG6T0gae7pU07Ojhagb
kFI1t+FgxwqyMoPyuGWUY6NK3lq8N208XjYcCVSXcPU365QIGRjgEmUgwTf1Stwf
QQTlhMH4yDZ7qsrHmxTd2GIIrLf7PWYrrdJwssiLHkvJBb+2iCoyKtx3Z+IVGJB0
ep50cy0dpPwkCAQ4GRQJFsGK04qkS3WtTyO6mzgBHh0DGaOm/sxkS96DdUzD9N5G
aV+y5O5/9wxMbLbOepMdg1MFIqbHwAgEFgGOdnHuIye9pKANx88c8SSiQFnYJeiK
vpI1r5wpeda+OtSF5ItTQvZKbHqQutAWSFfhh3QG1P/Xudj83KfDJA/DmRSfTmma
a+C+MPEWbGVBKVMps1yowg9eXhGvcHShvxLPz619nqOXOtiQ/CLcGyzq7D2z7ECt
PMKaPkyEaI6SqODprFt34/r09aHOkK6WAofyzTUwXfPwfbedtHPCtLsKXxoooFAr
E7nQBgxuLinMmj5W+vm2x+FsNCZkhZKC/L/a3lZ02m3+a3B7TS3NSlfonXQf8nb9
Aq42hto6EEqbTmWrefmfia64kGnPQX8MHgLqHaW8YyIwofmaxtgGJBfwCEa30vMi
vYejhYYYSz+RRDMYFG8D/i72jUXZBfRbpq2WnTN8l32gFhe4rqQw/Jz9mGJL1gna
7PdHvT95/SOZzf8Illbw35hctS78bYJTdw7/geQPQnBgj0EE+E7vyRpPbDBL9EvP
2kUZa2Q7vxn1Hh7j/9bKf+z2GWdqNL+YtZtmx3jPvIsMx0H1s/bDU8FHYEsmJvD1
RhwMl8zWzx51WQbhttkeExHZekPYUxYzdqLi3vNxNUe6ej+ouAnMbPZEahVP3eka
t48xi/1HUO9/C/t9ab2ZxwCkYnVnh8T7Cmks+VwwVC+dyalXlSCekmBhbCorTzzm
i0Bb59bAHEEZNb7jBosnp1OAVPP8wNia2Fci2fZtMEnta5A5TiCJGCZhRkYVr4dj
jEhFtvCpPnExPI8dAdUU0ZWur45H2Qb02jrncJYQobn5nxpErhEjIDm6vzmcsjcX
I4n2GikgaKHfuQ1VwTiTlnf/3bbMMU00ip/rMDOMPrSzSC+8CymIZALHti3h6W4A
TnqtbFouEzt2ug/vUVTneGqaiPSC0kJyMD2xIbDZIa3+Mxv+Nn0R2NgXrA0wHmvS
t0AkxPqxnHqVcPxvYmSV6+WSGyOeRMBn9Sf3jjFwumBZlsJzPpXzYqwzvsM5ELx8
o5QWkWn0DgvKoNwnckMzELw75+CW3NPcFmaDI6D6+er9ng/H0iJauj3Otylk5ogo
7MvhpUC1HN+ik+wixPdpiORIzy9BNCHGG3CFamJfkXySE2PJNXsGqPW6dtZmv6yc
5Jt0erJYhaYkmMzkY6zdQYSV4LD27JxMWYdYkwnNBrnGFWWey5vn7BgyX2tNGnMw
VsKCLOknDKWmURiKabAnDsR4hwCVJHSVgIj/BB9NmvJHlgr49M5tCvqI7ciFCL4N
okTqbsvVvFixvSQ0Vq2BRG5RsKV0mM+pEppgLgCk2lREdyRAxx05S6qWGT4y7BCC
2mEH5B2apdbfZFCb5g5Iy1GtzJXvHT5EjF6FmFsd1MYtoqZwDatGbiLbP+RL2SGx
BTkafflO6z/Hg/nON0ETknHv1FLmeHOanQrIg6VyNoN40BO7etJECfPxsrcKh1cw
+oylh3996fCZd4rkBJNq6S6f2el1y+8fFEHQhrk+xrkuunv9G23LKkazd4SY1oq/
pG32TGaGwxs2TKUFW3ZGCejSEfT78RPLP7RMPJ2g1jj6LKmCcjnZC58/t8C+QO4a
TJIoLuedA9YSyvCX8raRXYpNbseElpczzAVAHtP7giy0e0sNtLuJI5VdGVIqnPKw
fcKOLbGBeMSVQHAC3/RYWVvb2dos4/wJhFaOQnyyiK9GRipUGlw9lfWb+YLItDOZ
LIHiW71l++NtFMAMyirOJ0Y/0uyBhhidP/Epn3s8tV3kmLmar/UpGxu/5FiFvepR
idnwzfuU763EVJFqzg2HjDHhLZvOiis8NP9LU/UreCnHQoUYX339IbIcFp/qQWcg
UCojxMQocRdPAoFoSvWZYohXli7Dz/SMNZzBGHDyGl//DPvmcspEmFyLEdJLMLaW
wJs2zyXPUTMSWIDlyvGMLwgwwXCH17o9HZG0QZf9cTQL0bY4gbg0kA5rK9Q87ngl
ihHDZpR8SNhgX1WvEThRO7psY9m3XGGbCJn6ho5HjgfnusdlLANFLPWjUkpV5va8
H0PjJu8aW07MnI5A7n3/hwJAC/RkDGoQhlQguwF1kMWmaVJ+PlIpsQUXal0XCHH7
lhkeMedje/gXVFBmYmihBPGVqwfK3TeF9ZC4Ps2pepNQr7s8ybRuevHazH2lyY+p
BjpZBPCPNles2dpFf+JluK0xH8/VeV/IZ6+DHsuSgEYRMOfw4OCnWL4nSayv6l5f
1x1ZqkkIl9SzgjShlyUSHE+Ntf2vrkWeWZtxYrBdQpfmWW1zQxKuOesoNYElw13y
WS0flXQmrzpPvu7MTZJvDFNw7CjLsra+1q8IwQCsoq1G6on1LkJnWvLsJgKO0eni
rYtDjS2z2BiXXWQBagr3cYrYRGdQGKnZPyX+gwbKs8mKMB4WaiAtW+I3+WYjYyvm
ejRUZZ0GtXxmPGcWinLFzsn+uaheGhHNdKDF3sbBrOx7nxwP46GAnwyFiKPKxRhZ
dSIaXAy/G/em9O7KzAcJ6KhcAZGcn00xsyat4+JS6mEDqaPSqyX7ie+zkYaAj+YK
FR9auXtpbTulafYgaHOSynuCle3zduyfTMxfz7S+dI4y9HR+riaUeY8fwY+RxKaq
jbtnpxqpakZsHS4AlXgyK21piuprRzUZDSn0txEvvroGfe+Tilw+bwaUxHTWrqw6
x/kp4NzjX6V2t+cfo/EGCdKukEBTvAIOjdbpmmOJOAmrepGFluUsXMfzxYBJY6si
qJ5MRXoEVbPabZ8iv5X8MvoKlJuZeh7FTwIzMnHTrDD1jIE+XewESYJmGkTpKAFs
iSKmYdiKyMsU+PQWxadH6eN3MGcyvGzOJdHERSkxbW3jUP8KPql0LOTxVjxzvc6I
5fKXwveiFNwj43er5i3voqSaXJROxhEmMBNmWzg2RQbdktlAv8M0v5suAWdCL25J
0Xb/aU9BF+Q0Hcv1qZ9WzGeTKlM9zHFwNWBGBmH0f6cudi+YkCrB52jRUuQHdJLA
wArcGgoMBdzUkByyRpra6AH27niiWX7ZYuiRW990TlJgQ7JxunU/xWB5x4W+24pu
vJ0oF6Gf704tYoD5STTeSHWR7uyAF9Z0uHaxh1+CSt0V8zqPU5xtyn5KE3StCwyz
zqZXqRHUWV7ULjLfin5YII3sIU3gDHDnEo0SWZg2ZwGID2K9zrXBytIuSeCDB6cE
GtmrFHq7xzlzPgVe5DKuBnrNqHp4nXRNMuQ4LLU68P6OFnH89w1Saz4DDXq5a4GT
viHUX+2RC3XDj2QMlV9p+cxtQtPDHnjzXMwiKiDWT8ZUXVzwmdPAdNo+i8dovD7Z
LLxeg+JBT//Ham7HUblSxcqopDEUL8l7k3B93fMAqGFEz+i/8fvt2zNL1YaZIBZS
EFGKRla3aBKj8aHTW6hA1rzPTl58tqAx8WsPSodRhk1clH9p4XnZRpJ6odCwkf5G
emNbKv6PB1eRVRwXPrWuHXgIFnnWdEsW80/cS5LoLby2KJujoCc/VI2u2sjHYdun
1hY/p95tqsBh1CXHuIiHnD7jKvcx1Y0urMdBs8zBga6kTbxrByCymJE20VYLT/oX
ERiLVIdxf2TM+Ae8UkqWVbvx2jHZkO1hsVsLPnNYtColewNvvOtIjtYEs+BYTYnz
Ypk3aXZB0/Fm6RmfSEVvivUQsGfecGIMARPeMckbA335i6evxaNcJEPuANvQzKbi
sITsOUX3c6XqI5CJmGb8WfYo3vpCMLdvqGx+i3KDfKsC88wMCV8u0Q+PZBfnKtFe
gPWw+ObGan8Nzzzzg6rhLYwQ4IKb4RT0mQjBa4j8eJdAhh/C6172fErt1agkvxa/
Lab79b8qqr5H8tOV6hvNsRXsxNDkJgQ4pf7F2NMaxOKLOJaJiEQf/hqxMzbTYkAD
mvnrpTrDkrY9I0Ho50Ozk+pO+o8H2Plai4LhrVn9kmhlOxz6lAGsY1iVLt0xtLYv
+PZHiCdwv5jftpdgBQDRb4A7AWrUq0AI+p8e2a6MY3Z1FfGRRUWC+1K/inJ3u5EO
QI6SpTJ35WjbffBJQBepeXn0RiKlqJHZiuj6zuZoerOcZJhrHzHBAbtXg7dQbQPH
be28XWPNtlOaOJOpZfJQHtlpPcq77H4ReyP/suQVdkZbV9nVMzVe2CeoK65CQSHg
t2f4t86alZzkjbrHNhFiPq5+fhBBfrcnpvbCts8GjU4Oe5UsFoooH3ZiLz9S6vAR
DmNXKq8RedVFMr5zXIvCngP/sEMmVlBTKN19frOMmYYQptUxD2OTPEslQFhcW1oJ
i/kP4zTR1fCYae3Ru5k+0jbdtVIqZW4YKPNKBiKtV/N+DMdx/ScU4B9M1YgvNIW2
TeNNccCBficuwjVEx8jKh7fqwRfirV5dfLjQIGtWoOykSn4JH86UwO17nTDSQwYL
8LbUAyBjRoJFE8jY68IzMRFJUSI6CjKsz7Y4lm+aP1rlwQh9kV17ZNYZSi7Q3UeE
SDS4qb4nxNqu/fw5sF1M15Li3PHrtl8kpPhzWWbY/em3zBiX37SckuOz9ildpoHN
bp9TEshCms2Tf517XX5qXe/52T3jc2JNnOCYolrwSft7iwyPy4N9imbHIiWEIsW8
SyiqY9r3yug3x+3foBhqL1sVFdYIvAay0GuwKsj5EpzufTFNvPU2Bc7ytt1KLR5q
g19mBaFYY5tROxkTyOlMqyYgdwsCmvOHjGYevoBiQSiv3v0hFb5VGjEEPbYemMHP
7eCUtznf4N6pQ1xSFwjFss4YkST51yUSyo0fG6FCX5HnAemcAJkKImM7kwkPTBrU
SkFoI9TUUuG0HQ1BgOvAJFXgvPiOhuk+IrD14KFWgVeJGmEvC+Nu2Zwb8O8e6k6U
+VP3weEltkQAbcIN61RLhMxmJwNhNI8WTzZvtnm1mLIta5Cv4AtQW8LtCmLAx2MR
46dhXDygwcAb0tNE2ppaG0WrrtpfIdzeC6Zr0JNe40uUNoPU2glmW7OO6gPbFljd
NnlUvEUYc91NHH+geKni5lgbdSNiYqgJUHvtvUeowAPIvN5LG3aa6FJFZ0S0XBqD
WJFuIZyto5RAACIRkRsLleQ3I90r0MOa6yRp7dLXcRdmAqj7sAO9U8uF8rEMPQXD
Sa2e8oFj0Mgpm0fTfFlzp/iWhxZdXY33nA2iVm0Dyy1Le+JOOITBJTmxVn8vl0CE
banCGgjAHLAYNOWM5BolClAuzpC4ucVPVfrWtFx0yPDXXeQOfXcGKZ/jvbXiwqFN
invMk9/FCTo/PV5HejRnYigS5Y9cRnsYix+LwvEX7eCul5Riyrhj0IMXOlMA8d9Y
7ARBKhfD5St+tQRNfh4A7PJNPffWwEcqarRk9v6S4t20o0bHSk7NB09Vxw1WyeaQ
+ICclzTUA+h44KhI/bQsjr9vx9V3ATmhSOcpzmh1m4+PT/sjYCq6ZiRt9ZVkkJ6Z
4FoCuWOw0+6JyeAQAziXGD9dO3z8Q81jgSYJcoXHAPBv+rYvZQJSXWu4U8L5wpoU
vAPuLjm2nmMQCYMMhG4PBof5tZ2pxYPXybhWFMvDJmNi0Ucaunj9ZDUvsaaDRLp7
GRgcue0ZsKbQjIA+UiuVsUinG5UCIL7oZtd0Rzdc6WM9n9PSNuyA5QgR8/2goreU
Gl3PmvGQvMvYosZK6wOseikdmdEdHYiUcG2Bvwoqw6fs6XYCMMwwrCi3GGyeeeRm
HjCr26LRerp1Ua1jbFDpgVRvvpYzrxOk77freRWdJEvv5708KzHFCjX70bmvptoE
24FAY+SAuDcD5sfidsl8ImpVhGLUsPb1jeQp9aZSyiW/NW8tIt44ZBxCJZQmWsBt
tZEXFhdSalRxdn2Omq9x6BClQUvitsL+gjU2Mj5Ph8JOyFfP9+OrQVBFKZjOCdhA
N2+f+Zmh1BGXKPx6ziAZqQ3EtctWbLw9d3ai4Va50IJ1G2Weh9rOX5E5WSA44Nd3
+2Fy40jGrrMY/D9jY/EOnnTFIkRwV3U2HwEk/yPASxH33zm8/aWJNZIhi4Gyg18E
1fU9oW9hQyuQgSo21XAcv4TzsZnMqW+OwU4TBhBMYJ59EteaVs+T6N1OxzkG5p1h
sBJmo9F0OD5YXQFGhmrfVYQf8fQbqGnJIdrryjVXarh7IV7MbAAcDXEruwcBTyRV
SeBCfaZlflA+eKMWJm88pKZ0PQtaBouVLKdaUpa+ZXNRZuhV1AUe8FiDh2QcS8aV
66RaHZVbTCMvX1arilQBWBj1kWHT2Yufe7A7r3bmHNVz8L499OG06GkADJgUBub9
WV/FasqExrj5eNNlSArPBX3dZC4pnrekm4BZaMgcqDFtGENbcQHs4m7+xsvVlswQ
ZurxPOJod6nQpgmv7eNwh1+fx5Ga/up8WT0WVC1srDQyAxcN1AsQX/ydEnXggrJb
U9qdR8NJtQSQlRfvkU4+sKDg3YikNZLV0s7u8wVW0dH1CQQw1Hq4fox19LNpgzap
Xch4On/i1lKpAs7gnIY4EMMIHMlUBee6Rh3KUff59VM7cpI0M7RdSGxYOZV6/lZE
F/bRDjB+Xu1ZFCkkB5HCURroHTUABitzvlthhXRbJFj8rQxMloe6qWsUEbag/Okz
wJ+cIH1S20k9LwXD46SQR0Dxr1Nos98o0eNXoLaVZ4zYEwU4gNOUdiRZ+L4RATta
YvIqnC3fB86yAatC2/kt+TO/AHY4CPP/kZgwm2F/aN5FfdE67Q83vmGBDvFAjIav
jNI0YPLJrelbIkq7hgzFwmZ7e/yS87/FFqbIMWyieuBJwJBqybBepPzBwT3uP6y2
3uHiRzYpJKX3cLpuRLuRJJXw1SbkcrK+OmVYt9jvdW5ahcVOGAfy3/8otsOmj8QV
oR8mUi/fqRfkPMJEASg+/wVwV4j2b+AqIL3qb00RM/O/Fv8ZmvlreG2MS9W8Wac9
JbMfGqO/ysIyIe97P/LKA2BxgH+4VmsEgrl9y4iOjFTViXdSVmSPofQV0zuijpX0
5T/WMXK2xo7gNC/99/Kv4ROakehzWeboFaR7ftypxInRMbxFJmgdhKcEPPsx5273
o9TqCn/FprSJ9MrJTCezsA8UkGHUsz+pVosAjVh1bg01h7JXi5G4oKoGNGTdml2Y
v38UDReVzucGP9iJBM80Idt3hr+qXIH4C3m5StvP9zwJO2sPNjNs5rEhWJgPBs88
ZSb2bDYeiq3ZxAMu8Ncj+lIOx8eDSpehxjE6dSyV22X1tB7/VtrMXWJL7go0DsLQ
hS8wtoc2xD+gJ9fp7Q3/7t2reK6nOhyT1/pHjrGsM8E/iE7D3ncel4XqQ2ULAonB
WmeHeEzJObfrkS+2CP9a+g7Pyoj6C69pbXt0rNz4qiB/Vvg0YRBHN6CTcnWZf0fM
ZL6R+Cjwl9h3WIuQKv/0qaup9L1HMzc+QmmP5cA2KERKMEk9CLFIUsCwlusUEy65
HK28MvyFkG373ra3dd7lBIiwzLaMZwNEeJZBdnwotOZ3LpzDzm/2VDyKa6+MhyN8
+759EufiMnlvtOYiFsQZzqwFQfa3kUyRh3efJAYiznsX9TcipU3kosGnVAy27+vX
jDf9GD5BmUjekFCVTpMU17vIxwshkTNqMLRjvpVvu74jrtJevC/xjVDjiJBQNfUJ
3NhMRwSnywkFF3pM/kIFFzl7k9NDScCxNKvd2aCwRT0PE+o6bBWX04VzZxT68xOS
JOQg1Di8oTU3mpYOrJ4JPrZJwZFGRv0VGhtGianjdhGmCWkj+8c5uR6dRcULWn2S
4cynjXu93SoPd88u8HseNUoSXCSbn9cvt/d+ydziq7DvSHDiyjBGAP4vbm9yNGnA
jT4EvIMj24cjrH34tmjLH+DLt8QmiWVLcp2xC2h8hqeKoqhuP3bvLcKSaPaQ+7x1
nAjGgD0n5OfUhYo12OnjuMt70BkEBkErog8jue8myf9xYezMCkmYbVbpKzWRA2WM
06G4b90VwHaVedNZ34V7YE/b+VnRYt/D0geNujRAHLPXBSwzi/fSu+LxROfAsAgX
Btf4yVWcCAa34WTOiqHhMKve+ARXH33ziHeRWrBBQuiTWgGVAsU9ANAuTFOEcKUJ
izktAnWLMVqc1F18HDd7dLIGroGykRV52+bmLfvVw/8y3kHwO8714O6ixbLLylqF
fk+erkTN5wT/SLZUQyTnNozIwL+2B+fCOPS2sn1NYVpvbV7d2MM0WJFmCX0BjmMP
nvBOJ/jb7Kx3UbBZWmrc6g9wVnQ8jRorLef8NDXGLnl/p7wRSe2Ot5+UDJS2iezW
wZaTVPCXuWld5cGPeHzZc1XFnIYgeBr4WfkfbwBoyJGKjklp73Zhlx/hPuk5UNmE
6BA3CV+Gp7Ui8qRNF3rxiUJYd0VCJj9JIwMiLq58T3Hon97rWsx7HlP5ZRKHnzBH
8sw813xy0YkKrN3orpcbghu6RDzx/8K76fJW64Rd64ZiIKBSMzNm8rNKIOjQajMs
yY+oszliXLFG6ByduxvvJvg8vOU7VkVXZ6AVv87pfihmYk5qzctJwGTUEt5FsX+Y
5Qzo9BlDitrfYKVr4bJ1XAEBji2XFI5DAUUbGpY1+o6y1O+XEfKbLKDiDHM/n3C8
O1tdvr4CTEKYJirUFkVwg9594FPCQye8Ph5buc5RIqoANeyqAglYJj1diND34cDk
AVmyDPYNbsq+DsNQqbXtXMSz5W5+KyR3PeJqLoVJyoQT63d289HmR7EPgmFWClbO
jl+EopwgwMAtTuqoxq9MoeNxKzyHYAZxmxIBwAHegISVu7awrxwZhgd03jJtLd5N
Toy0taOC0RZn7dxItt7kvr7X6odXoY4GXvMGa4qD0tFHpkIZDLXOwqB6YInbSEHb
S7iDaGxDxC5Syu4n8zJwTUoxjoukBFoZgQI2wTC7ds8IfjgfuF9n0oYCRtJSJld3
/DhR8uuii/4IMYghms0XUUtc/P77vYjOWIU/hHVnnY8Sai1j9B9T2zw7/uzKF/xs
b8r6sYfRDnQ75IMxPl7NbaiKlgTJ2IVqdGwgCDHvtEvzbXxxYAkY9zatLfsUUmwy
svxq6HQ0aWVwmf8xIEtMPZPS4FcyJTsG5pzg1bnf+j4bFV3wR+xYI5TCpB6/JIze
aqAhDT26CN5vgQbyz7SVFGjnzlYqBhvYimsfaCAJHzQO8La+x4x460YnsRLYEqIw
koiNYFLnJSyOFdxTTnA086nx2RcA33ShrEjuWyubww9gZLEJpuqijUM+j+4WP/Fj
h/DyDDtrHtuWzSr/8xyPR33kSJsGvLp5OF0uEI1tQRPuRnVV5asxiBtcEiknSE3Z
sYKTU7a0kCyayyD6afywnT3Ip1jG8p6Rx0B5dliQ6+ziv+e+7Wc0h0S3qTgdeO54
cuN/Q+LCFROdQ49iBOLN7lHliVOCXz2MW9hVge9Q2pUK3ZrCs6JUDTFw4NDZibKi
xuUpobsXQ9EiGB/koCbKFVun55vq+dsDCt5NMpaZoGDdLB9pjHMvFTAZfzCdL3gv
I/sHjtmLWnAtgGz9BrYtEYDb6p/lPzsMgwWZQGBoyMVs127qQ6fMZoAfFhVrbeZH
QEXAd4AccA0IS/Tyt2mZe6RqmGFBRM59poGmWQQ/GyTJKgEgXBTFJ0vI7e9n4A4P
RIC90Tt44ucNG+B2bM5S1xURpHE9ZaGVgPSGqRE8WTvS5YciVb+17I5plT3RcAmo
NnSnz67MBT2aT9WiQn/hnVq71Ndi2RBeVtCFcNIjRLQM6ANe9DAvN8D9MiNXS/lD
BFoQf033ZN6A3KLlsyBUQ9HsodUL0XobifcMGd1OYWnoz+3KRbsugMDNnhrsF5jD
C2tlUSByVj49mOpVzlRUh+uRGvasWy6ey5edfX/cx9JIPSLSsKnvBE4lg+C6b7sr
AvNLx4Vam8sN2P7TI+D+lWIZ8Ltn5BVPqMies+8JAX3noX5FJLudVlL3wJE1eelv
7qmuV/exGQCJNl7jJ8K1CSP4v8XVwLoqLprmLgWtvkg4sfsBxqHKpfD4cuj4gfin
fPL5764LZpUzVb4ral7GwEVPSJYJPuspOijH+4v+4/2sNNeJAWoqkfRvjEeJP9OG
IvfkmWjF7UgyVj/bhIaS72jiFW4YFcl/djm2sQjJsJtkMmTwvEcaC9HSjwlYLJxJ
Z6259wiQcm+bsYZdHJnDgNCXezRBq4822qlHshXTdSPMlnfi4l6cj/7gFMONJDXR
6SSgiXtrJm3FItyPulYV6bmuIS2vuKANET2+JZiP6ohBrA+1LNJysUMThq0yMNTP
mH3pUZm8enKANxa2F74VgLXZO0tFicjecNCdFBBdVlSMxBkkhG8X3w9y/TVVlwuc
1656y1VWGdR2JAROVne6lmH/C6BvOCQa323gEycgGfRyBOrEjvTQSS+qlS4bE6s+
7k81qpL7Vir6n6Csp7xSmvO2ADwxZ2DSR3oCNqRbY5FwDfe/cJxzvtlvnk8swZ9B
7E+mNgDmXEHjQAFQkOxRLSGmxZK4zfHMdSUqaaiAV3L1A650FzYhZRqJp7IHC6Uk
82YZY1kV6l3PSvV/ndUIxbA8S3H76tGGlxmPglbrue4cgNDVTLeirdX5MIQFyNV4
+D72I4IhHgaFggnmRoI/Y49yoNzBoYuKYv1l9Y1shNPbBcXtNH1/YpPy4qAn4oYl
jNAa2H0YeSwPUR63oXvxrcuguaUTxpdlIdf387WM5d1BAlsb7Nvtf68Sgqc9xoRg
UyWOLeH2qxG2bCbntKKJv5taflxUgiOgP03yBULcR/+IcYzawsig6zcXdkp3A957
OnLsr8ts1jRGI21RUMpvr94HObbGt+WfFL1TaxoilaxuF95vw6YWZZGXUWh6Hhmt
x/lTIYtEw3vBWV++aQdXJBDaoXabGVOKsNa2/wOcFp1i+dNCCHAxpjQn614M0Th5
Gp6D3PfTZfncbU4Y4KlSGB8Y1XTYyV3V62EYEJMAWDp2ZhH0k2WwCNisUsRsnUaU
7ch4nhObG2vqSYmCvnuBq7wEHmxypBQr+Z21AZ2g7sTtXEnclGd60yWQEGM6gGkI
oTnQM+QU7DJLNdTnlPTXww4uLmNgkl1nd36LDe4ST8mEcmedYsBCAtzEptRtNTqs
brmjsrk1QVrDnifU+dV7uMsmViMCnQWYGMper7RzSLF9fBQ5x+vMiQi0JQLt+vb3
qOVl/qEdUn8lekZfJ+y+AIftAFQEwKdtWN2eI6DF42BpWyfjItUp7QPidCdAdDe7
gDOFsS7LPcKtBZY1kzKUGTuGNCp/TE+sMidqjiAKAD62QEf6v1Dj6Pl7gZ0LavTL
PiP7L4AY20wvPUq3vPgyd1eR2d9srFIG9is5d0cLXdZ7pxcc0uFiBtHZNkl7E7mz
j8GJAdPeaw+Lxu2jWvAplIXtSflveBPFIuAsgq0CPfNgV7SlkvDFzGvkMa6geD55
U1yhmVQEGfIcbEuFVQMe674BhQb51/Xfqa56xoigGW3SK4DDkGuzc07wHQ2CDZzO
QYqvaYnxJ7E7FqeVTijlf5pb4bibo8YYI0bR0Lprj4HBcgMj827+jBeqHGOAG6Xk
JxL4UYNsuIljlKaqAp+E07H4J0lE9tB+pgibClY0GLThwuu85bSpHPnarkOABlUd
Rh/jGY9VxCVEQJCaYrEyznIe/qtehJkULYFULIC1dXkrnz9s9FB5rO2H8sIz4+RT
CzRynEqjKC7ff71xK/1acc4GZvJh3OvMwRiXaw2lBtdjvg4Pq9tprwNGu4/TPRIc
3uEgOtWmM5a6RpqZg4SMRjpFeb3uN11yPq1yNWn42EgDWdyxBOgFmwN++elQvF9e
RhyGrI9s4JsWsnUPhMcny1/WdLx9OPag5KvMIxeRpa0O51dqImv3lnwsL/G+1YXc
zc4Yj5OopwUuyHoYXN4AwJoCCBx4NJJSt+QRn7c/mr6QGzl6edgEocn0o+iD/Qnk
bbFKtjzbmE18xl/OqKbypW/+px674U1gQKOOAUi1p3TtTjDqJiIll3tv8GWEVA+y
F8xF7TWCzxSeIzpLglaOVj4H8ta7pTgX57Tl2cpGpzairSdcnwVDP5UZNXExEjXc
VFGJTDX1sGYlkqH7xRLlYVm1hS8/AKvPU+q0N+uvvpI5dQdCBIxMDrv3K2MIHz2T
j1kUVKE8Lh99BPiXb5/4D/F1YZUR2OnM5St2ZA80lD3MGdZpTgDfkrJXvPLG3Kon
bJTeNyDOjgwPQwXmt9VpOL3Pr7Z2ZZXm7WFjFTspH/sBsGvh8Z+rDKFxmYzePVx+
DMoEGellFHXD9gvdXSJ4/eTmYUOYaByxA73b4RPT0MQHCe0IQ4SBHaMqqHba8Ceh
HZ/u32d83tg47p/92r9PSIzKwYwwcucvVRs18CG17SLBxxIxHjE1iajxjkxlE/xf
7VSej4mwzDxmM+mCuuR57vgtVI0DYKpPPZb2Hk54vWIzrGMwEBQPXfcpt87DURvZ
vVMaxD3rSNAlnhB4TA6egRLB4XK3Lz5ZE+gSE+cvC5qIgCirIfORvwhuglaD9E/U
uKpwFmzX3Ycnb2acPh9UBvMzg2XvvpWMROmud9G2fEHetiGLHyEBgflCpDIsQfwZ
hVjGXtGoBuBgaYxw/eKOMHeVagAELlGMc9X2w4QhAoyHBdsfZEW+GeXxxkl8f263
Sbtdp66Lh7l1LYEsflSMfJaWw0AazQwWMGd/w9Qy8PZ6yllRZP4XzIGKdQI5lWUR
wnh+7oo1+1ac1ema7Xjy4Iu+otAAFUSiWUhfKezXj9/f2pSpGp8wnLISQqyI6//t
DemnF10uudvnGMOV9VgZffbY7DcPioU6/vCVZxHqHTsPcu1EdX1/HQnUaoO+Ms00
kckMAx9h9gy+DCqw3QEtCyryzNP/0kSfwYWsV9GZEFJ/Qe4G6Cc5MX0angZawVPd
ZWziB+7bA8hwSYrqgKGGuQvvMRjQk7i2sIohxHcW6hdHh95cMMjfbeATa7ZxB6dY
B+ertLl2YuEPExpu8B7fDexYTF+w+i4Jv+40ZnW2Y95EzkxVeWlX+xYY06UhmGFT
ZJknGHTOea8SqXLH+bEK5JGXZy/aLepddnJbvE/5dpNEQPNeIa/n7/eVzpr0Mf5d
BYll2gKuboQrT4MS6I91ubwwMvxK/TlaP3pn8gPf2+ezlG31DL8jczFD7Z3tqxoz
9W3FFFhWxAiiMf3276xmo2k0J42vHdw+f3jtmQXYc1wCtswz1+xqEO0r4YZn7A2q
xK6YhPM6jyL5DA72eB/7HdSw3xIS5xK6Zkq8v3WcRP074Zk3L8aMx9w+VR3N8DOa
zahqYVCGNmEj1Cj54lFjGd/yIW9GYjHBlZ8obX7lkpkdMq9pl5FPuLD9A+ac3jNn
G7JrBgAy1LXa2VFDvyypwvR9MZ6OlyAYg6X2fCe+Gae+kYc0CcL5y5lQs70Ife/8
2axPBNQpBAhcWDJIN4hH4HqZDdPwgUKpMpSinK+UBxaAu58BZJr+NeFQx5gZ5PrY
Kwbc4h4OZrwxNOYp/TOQ0q9NCG/8+TXYqofTo0pI5o+aEfdSNrj9tTTBzn/9bTPw
vI9gQmifHnDbjwdOpin1Jqx2XSYmwvzVfaFLf75kl10r9rcd33wpVI96orbcKuRC
EWHBoofD2ypbI1k9NSmDr3siCi7eFxNLi5nQPMgbBt1jBtZsxPfiDudiW7I/Tek7
GukZJpn0m9cgjGbhlhn1rM5bN4JBxMKxnVYNP70RrWLacoEAWCc8Lto/yVdfxwBF
nW/cxo8f6XR4Zmh0hmDEjoHr5Y4JDkrXJ3qShb9qPzDVG7bNI1X+/qNwzLn9kFpu
l3oFFkKWcPaxpPANXQIqfzIQ1urbbWA8kL5OaPBNugfvuMn3un347O388F3hSvj4
2OYnzS2NNZul07sjD0sUXq2YzBtanmXYC5fOMm3W3A24YorfuFnji12ILu0Wcyfo
GN42F70GeUcwkC6t2HMJFy8/xUjS5XhnQ09HRiuXtAid3JUXtr2qv1yEFotMgiHM
5oJa46adScmr6GDWnPjMdD0PWP8pZV+Kh0jvxxedPcNlE22+gdOEHb669AwzfitZ
DWty52puGJ49wZU7mAaNc/RrpBtfnWMU4KjWcMI6aNIv/x+zs2k8pE/Lfw83jCXW
eTZYSw6HZMq8IQ9aR9SgKKd8PKxlBaSI3i6JvM8VxDMYG0/sJLc88FQIQdZ9ETqP
vmd3FJ6L36IK4eDL19oGiSRqCEJrX74d2jt8wLVpH7hiN/rTimjV+57Wk+4nDicL
gcNc7NmnwTPcX2bbogLnBOcx+JpC5DzDmc0bGyBb0DBL6TfCUElxCpCF4QXOT6c7
31PgQt6J9F6D3p4h8qkaBegWN5lL5CX8+MOX+bIxkI93z20xx8JgPocVX67O/1f8
H/sZJ28sNlgQb8prgs2D5/QtyOOX1utSv+XBEzdVdX81top5jnWwUVPhs3augHaZ
um9N8n8c43NByBKfwrS8pOqw0WaWdEGE0Xy5WttNaRhAKdbJZMMA1NxvppZlTPjj
IHgtlNT6PgXEti79o9htrL3QWZLMoeq1stUPtDiWz+hCslTH6+8BNHNZWtr7gjCT
XhBlpkASJMAch5QW0/Ibb4bh75oLeOy/ive933xz6n+RNh8sMhCZ1Pw0EXGjq1JJ
4LRlq1xOpJtYjttdSpo60zqit4/5O6huilaZLMSxVVN1yogOW+Z2vwOQy/oPt09y
P+UYZuT7fE0Zvq2nIJRUGK64WiIxIddAVCdGHIuJEj8ECGQ+GMLoNaMO8O4EaN2K
q2LM2mXwKHMxr2PSIeHckbGHSGYuYV5Mz+igl41PqPl5S+QxrFlMJbOo10YxyQw6
mamPJLIePwqdZQqzuqqRcBLUI7TNDxKK7p6BXMXHxog4hs+8hjjX4tNEMxv9xa6v
Wr7+E5dH+RzwpnPLki1Llj9Yi6wT8xkDAuAjQpOQKjvSJuQEImKTacnHB4nQQgmr
d+IKbx+VruJq6BiQHWG3KrLR9Jl4LzFJkKn1hZvqW63NsB4iwQnEYuMLCFGKduxI
7mP3OKtCGjFhFQNspd4jCKGbMTsSq5NZxcnfN89hnD+AXp7oSCWLh+EkQ+gsr8D8
qZpQfnCTstDoSiMnPFbwyLAWTruJ71KhX70jWTDKyW6SR34HYWjJl56Tlz1kFJC5
0y4gMao0c+MOnlcwnNaCyr3Pfz68c5WQXH1I4gakJmOyv2LET6RbznhsGz1SEa4n
KfO3a1HzzzvLeCz8PxYgIDx4XpfrSokIfvk1xmJwxfspBpNeK9vjN1u8ZDAp/+9P
Fy7KHzb4FkARnHkuXpHzV6nPFBMXxP59+XNS+0HYLTQkye4WRYstIcO/OsoAx+H2
nl4NlzjQKyEi/wNawMENywFqkXrb2NGi0dVmrI7iB5QdggOCZwPkiA9AIbXdQsRv
tvZHEdNeTjJUcNgBq1ljTxdeR2XCbERvTWrJXLIZkDzktE0rorfjAfqD8aLGWXTa
hidkXsKH8kPzlDMNW3o5N8AfR3Rj3RBIgB4ylHWoeAYFmGjDLjW2u1knZwnbgUgH
Vzv+tHp/LFvD0HrbcqGeLn5ChF9eRNJ8+aYl4kZI14oe9HpOdY1TFUnX6ppECUiM
seI5Xu4dZtFZalH4V+/trRWljLRnypGQK1mwyrqLc6evCwfrIswt+f/1HWB936m+
ulT17f/GxIkhqNmnGAAtQCc8Bo6cTAk6SX84qB/mwn/OL8zs40lZucmOwktkx/5c
1sOpMXIpuVgqqMaO00LL3jqzFKJf1RpMPJhddPs8D0243l22t962ckv+UHcMJstf
66243e3nqU1XEvCB6+vkqoJH5J0l7Ee2IJd7a6Q8l1LdsFvWn9g0kWZEWWZUS+bO
JvLDuboQ3EI3hqdshaRN6fu/by0qVIICVgH8oeN4gHXssB+oojRhsxOIyRsk3B9M
SMsCCFbSsojhz/z+WL2LZFvq+G1EezkOYf8PidjuoyAAHhcZSrbb0sDRGa9rfM9j
g4x9zA2oeagebWLsWpesaoCoDKgMS2REEpKEl57IfyZpgWMX4Ok7SVgpcqgNXmCl
jjR9XP0RFb8tOmPFLCX7dJ5DKrNFO+eqN7pGnFZhkoscHTA6gas6dXiCqicpRuV5
tR6rGrm2S7IP0WqDqFPTb+a1HPC+xD/DQRvhVZd9kalI/C5JZgREt6W566s8g8LQ
miR3YiEJMANKeSxkc79LM5DfobZRaNja9/kBW0q9/bIQeexIJvImeSrZKSSusChw
bJgtopPEs+RqrWuXgEQiE+Ga3P8Asg2VgHOMbWqbUWCXg399IKNzTkLeQlvYpfdL
f+hnrdiltspfD6ptKVHNQ/RsniwrtjdQuYCetxq+L7Qjzuxs9UBKWOEzMYx0FCgB
3kktyyS+PgCcGur6ZJP5n1lKsxYuBUp4aPlzyFEle1w0NeFzX1v4oykdTg9x4GvX
rglo2UhHFdIWbZymqS5uf4HX+i/5dJT1/PdqBVynnpIKTE3XLqrzJxTKOwDbaejm
9KqqVDQBaJQPVV9+HiyDYo31zbzNZ50/Pt13xhbvl1UM/71rg/qRdEDf7xdit/Za
xJ+zsncsXsU9PAseIWA7fsBYK3yIjATuEyka0CgZYA5tycFLmVy+Itq5EurHb2iS
k0e/fOPbWetIt39NgdjG/Sj0n1nw1Yowu/cGEwBtPCfdDZ5jeUoXPzkMVE226x1Z
waBbQ5c/QcJMWLaYoRcdNzeSIKH06/HKx40yguwUd6MPsK3C3TN0fI7Tzo7VPSI3
SF9lifN1WIXfI1rdKWXQ18dQjF+TvFMxmzkTiWcK/dTu0CRGRgWlXjdz87NB+sif
QLeX5f+kZZJfpy2rJH1XRsqEDgdjGp74UnMvzBqGAdZWqncdeFxTokobCc2M8Nb1
hWmmUyzcC7nOciAVUXV/2w7Htg0tJ0mrqN+2UevK3FfYHda1pXlFPHB9iZEXuJsU
Xe5ioWKkJ+zwLV4s7XjL1nZBPXZm4KuvyIHtaBjmuxedHnOHmSdgHGq3vzI81CPp
adKYJzYTqqnV+Q0a0Ln5zV+rO5PeqwhiIjwMaeoYCbaFWgmM++N6iJw0CvlhNBCt
RRZ7gSXIZ9XNauEfEHHQZUSCdbv//kFBl9auHXDX0z7X3PaXysoH8NQdjQdaRISi
LUngOmPw8YJTI7rukt7WWAoSARfimuE4BYJJt9EoZVo3mbCqCd2Om5NnLOPX0Fav
CZpE59LbLDB7xaGfOTYg94z5VcBCw7w/xQ3HOq7sZVmLDUVKLI5P/SQExX/O9nV4
SYXZXSS8fB0/n2TxE1F+Q9hPAZZAQYvqrYxty6g6MLrpY9sniGda5q7emxSkZ+Sg
T/paxbcJFuL6mRVyhK4p+2AoZtJsQm/oMLTlZJQktoF2mrG551BI/JuiuZ0PtQ3q
w01gBuEw8MaPfo0BLCjbGWxtwBW0O80VGkkfZD7G8B73/jupaSRSfqcnticDRXo7
HayTJbJjrZWtELLHJ/du35VwoCjHr9NIzoxT1WJ5mxDdzoJCpVbSVkvSMYuAy/KB
klrCf6DgpzSdvhXS3ZKTNyz2CJI4TuEaATBF0jpvZkF8QuwBAA0LPcn1SqdDbNvR
x4QnKtTvwDCDc1PScu/C+7jeriQwEpC1SrZKNXaQdLDTvskUKPlmIst+CkdSl785
K3owljCTGECph6q+3bbsSG6FVSLWNXas8FFOKYXkMHs33fYlhMy8nwNJ+Iru120m
/QO1NOkqzKyRn5V4MmWtrCM0MGhw/VBA0ksvhrRnSzpKs5VpbcD4hN01rVeJAQTX
KP0NvWonGS1kSHvj0ktC7aEU/QpvakdyzFjP/PJwkePfff3aBeGRgikNDotIOzhp
n7koVfuF/yUwoZgJhKwDRbEab5rnCYpst/rVuzM2R7sxuuPkgqOSCswR0+NJ+2HI
OkjjwilNqXvOCPTiMgH/p74e5uvvqc8a/mYhSsY6bKOeipiW54qtYN9c8VNbR7Ug
GiEFtU9Ijhbq6TRY1ZUzGhknIL0duKYTFlYIGA15s1MSD8dXplX3EZsdB9veXVI/
M6kJQ9MwOeZjOz2jJEjemp0NEp9TRWUwcY2678OYge76tsNpJTGHQqCy50w/HpZq
8l5AGQI/ZFb1dpF10GQgfEjaqxrYJyUZ3ufsYGVsz4zBQNXq6sp0PT+sP5JfovX9
/H95sGXawWTNpnlNT+NiGOIgWeACclsBpXOfmXhkWx2b849LOhzS5rAj4Gh736nR
9ViCch5+6u5ktUErnoiiu2dw/ZBO1SQndUgI5Etwb6DaVd+qBEfFBqjw1w8WKxO/
/7TXXSTg8EqfEdYfMq9932j07TSw0KfwoOYqpNFh1cjf6rBMkG5k6UAtkBK1Yc0q
XHUJg/E97/gYSDePt+IuCASRtnB5HnzSOF+NhM5PPA27lkCiAYJMDNlmid9j69hj
UAVn9WCQ8mc+vV1jbGTezn3pGTszeUh5p3S8iOt80J9U6hBbYjXKbMvwlqBBrJAK
0RBpqGHHiSAYecmRjO6N05KnFis07hVIZ0lZEjv1EqLh16D8gCcasFmw6WNFnsHQ
ApJhoxQbsNGSeJYN2PVydYze4aNA9spn26PxxQjKkwxXf4b1hhrHz5Bdn6NrVpto
7uZP8DyPnGoZ5FLLRAAFwd3eVU6V0pKiVokEwZgVFN6UZ0Nuh99ON6TQnlQF5vNB
xNLTmC2dMkwisDmmzvzlwcZrt848mw5iswuryyaEmqvLaDvULpjapIRukU8IMpIq
8u45l9rVJNHI4FjXlxdqdu9BLw0nsbNAmldchAhr8wM1dO2y/8rsXzZ+8XZ3YA6I
W0bHJoiora4UH27TDNCGIi2+1fPcHPODBYp5N6BIxcXQnRJQ9hdJxjcupRtwembG
5NPR05WNothLmcJY51X7in61Z01V9NBRHZAFSenoadoOhk5gt0d7uDMvM+KnL6NZ
1kZUyk/V1AnBNU9kxVJvhhsd4NcuMpi20Z1gjp665nkOa16lSfzR2LI+3B2OV+a6
+6KK8dNRw8Dv6VnXSLziVn19vQJ3YCcqxb2Slty6dHKTgpuT9skOx43TcQnW/2yK
2DYHJfh1RrGIP/fWxaV0MD5L02Ssz9VaKoKCMN+RfrnTG1oxcnWnooowXxC9g3FJ
aZKn+fctzV+4jm9E1iXaDxKMQ7tQWcb5BgQ81XL8lyLdp54/mOP3VwOAXcJAV4W/
8m3qiOv/zwrwoO6U2EjAV2fkgCZKFXLeO6gnoPO8utiMp+lCZpWx6iNPDXlmUXeb
8YJcpG1QGVR0ElmLz+oAUl1wyDnnf9yopx5wRuzzx+lzoxnk9yv/U+ZQaspaZ62x
egepgH4huYilKDnTn3WaFz206sorSEvC2mF8yBAgZojirYo/GJBbMmv05rRgkJEh
j3ADeJv34nMDJ8i+Z4Labv7/c4R1Sv4sRQKHx4izd26vhWToHRTC1ptNRxlar+zr
0jwdR7bUVQBuw25qhtqQPP0l9MmTD0uDO44nh8ebseTnCK0rL7i0B01fyyrbsx3d
R8DzJxCcdbhld9ugn6BcR7FvMJOLtHhyEpVTEmKO1L0xWbIk6EPJcozBLFc+EL6N
UUdvnGtavnzPWh2Wrgn5jkbfzlLNSbfdi5OtEyCtf91HP9zMQZa+xM5Tj8EwRzBl
5uinDi4x7nqx2wePm9o0cTKdyRybbcAxGaGKozlA1ZErFg/brTPxryi/jm55Mwc0
PFzSXdbc3A+Oy8YW+7fkgphNu22s0O2T1WmSgzByPKK0aGZgox6ig/ftu84hGAo8
5JIJsZTLjo8U+UvmCYnM97RGBj9iQWxK437Xw2hiHaKZuMccabmaA9AoMZdmdQ57
psy1YVGUDCAuqUgae8NBV3yjCGYlcTj1ApNS1fOQ2TAMzfZmVO/fTPN+Fscp+FxP
05lBwr1tkVmtj6pKGFX1YRM3TPgjPp3aDs2VPnVhaslivZEoZ9M8iymm/ayY4WE5
RPCS8cxUpeQDhFVbi5BkD/EXzlpSObxA2wiwNv9tNvXSFbR7sBtaWfEXEETmnanw
qqh81q0AZmdEyH7Olya80JvlNFUNDg4l//A0aAe4RzbmxjUoP+tAavlU+QhKD45P
xkOBrVTZeH+jnfKxHb10VVF3dVPem5Mh66sIsVCe4knDXHmOyu9VWh4ewYJLNMSd
hKQxjDoklnph7BxL+qVc5Gv1q3iQMQzZy7TSUHG/zh7UgdsGonymLhSecvTd0c38
nl+UHBvP5FqWhYfbbV96lgA/U7gTRnpTY5k91ofyFOpoCcQpOAWuklQNkhBPlCFf
3pIDvCD6F/iRMwLN9yR7txudnC6gau8U1fbPQR3L8W1d86Uc8TswcRWUoBTYgm1I
qmAqdNFnl6pL6bFkrjgpl/vYIBzwIXuKm5btyUeIO6TerdMm18MODupVHVfvrng0
U+TlZwuxtVh+cDbrXIWh8JHUz0afQYqxstdL3hFXQezmH87CKN4azF2gblOyWL4O
oJtb3PiGROoTddjT4LV6at+4tbcjzCBPXMpYtqZm1mF026bR3JEpVr2YktCVf5Mp
MdwKjmqgi96zfxXlM3DbenXFnZLKzGdrnpyCLYKieIxlXW/yFyHdpn9/Fad3uGXO
B+1uvT/HMfkccyR/hilhEvKX2b83wPK3V1evri6ZoJIArbsmsSF04iLABiasPRO4
QnCekxweNXxCQW6lqHnXzXw3J9M3/901B9fifnBSnYRGgPXptqYm0MI1ThfDSzus
hTGNMlh9rGb6plbEr+57OeInKXIb7q9qFqEePgwENt6IUT94VaKEpqWHhlylnyWk
P5odJAPprRztPg9fCkwzXs40F6TNhIueyYcJeojKNjdghwnWhnkhY+BS8RHb7Z/l
KebHMEOYxS+rr1A+ggjhU6vWCGRf/RioKYmRK5fOP8jeWUa+FeA/fwQFzDGnp1kV
db+jfFRIu2iIC0u7njkGNQjrZAaKlJ8qtQHQ2l08YiKkfMaCGd6NEG1YuThHRIeG
Y0KHLSt5KwFrFJlhAdos8jcdVR96ddoVRU4Z1/zsLiaxagN4YygpdrMx+ARw61qs
fPYhMQLsvXFsdoyiy11fH5ecgaSP+gFZgNTvGb4tlI3bGBLJDWzxfzk3t2Bxv6iC
IpayPeK36kb+S5xguha7DT6ZJW9PHBgx6ew9bNjKT7O7q/oviIpIpIFCPkT2FsdO
HU0rcRUxtF6powDXXAfMjylnC4TLp2STcF9yvO9+p2/b9L2U4EkPeXdzCHdH3pQF
w95L1as9sZ9xZrN313MP2r144qXgZtFZ6TNY1ZReewwF62Zr36CZiKNQk//LvGR7
RWGARS2qDTX728Bmy3VZsuws0O1bHUqVbuzvwiH1c6G9E21cMdcfHYfrT4g68VXs
QrOPljQF/AQZQYJXZeAXSH4c3vJOGdJM2zJiUeFUOLduZvHSPEQ3fnYmwPxi7ho5
raDVrB6nOe5pNYeOb39GaWdOw9Sg6hAlY09MCSJx5KTls1ovyIy/8EzD5DIZgUAG
Q9U9QwDaAJ5l2pnJa41/BcMS2PwWnC/LX47TqPakTLFT+TKvzYjBdA4Loi5BSvhV
99cc+CjkBhs55nt8Kqm/VYlTXxdBAlcOZlwwFqRAGo4IQJXpw13nupRNdPizDQD6
8tQRIShyT9t3fcXiMLuhOUKPPDCj90cvTb+Vi9ahPwWI56oG1wqNWQmYfofCM2Dc
3psz2mBOQeNTTBFeOKX33y+I1FJOtlsy3coUp68dpWsXi80VTnp03fQRj8fQqj3v
Q4l4/tevPOwJpGoeatIwct9EzXWfgYiT3ss/E7OaMHs57r+6a0kmvwO2WL35zk9a
bk+dPSEgsT4OOEgq203X713rTH/Os+b7NJVHMgae+9Zw+KSO8dHG0W5LKNz3TLYf
GTTsX5FFSKq7cPb+yX3P9b0/mq/AWO7PJZMiwauoOycOEUgyLIVM/d4XGArzXe/R
KAr+Cgr8AawuMOL9KjqKJwMi0nkiz8FU0JsoR9Nl3sQ9LS+7377pcpi6ulnqdHZV
t849+lXJTpH3mYf7S2Z7mEFIF8aIden+3VVoXvxBq+7wCOqHhcHOK44sSAfyqRi0
g8gv5NC5OtPJu4etDYX6WP8DgeP7WjnHXPhLY9NdgoW4ozmndT7aQKECevxaNvxz
HlKBxJzmOLYKtbwsiq9YYbq4pzXqjIQ28+PRFlAGTr6fl0MeB1aqCrnjcT/qFjrI
9zYEe/hSWjTkh3d2s+V2ETMwmgB9ZV3dI//pbj632Od/62icp1aXI+c96XAXrXdy
QTYUtx3HUrnaVwTkdLeJAmJZTfNHOry6CMTeJgRyGvHhP0F2XJbwV5TgE3ffKxiS
woau1lPZbgRC3gNqaX7Un++XebDMMV9Eg/AGzNqE7a9DsjnEhvQZ9la23QkSE4cF
bRhIq7q9LXrrLMF7rXBUZgUbogMvrCZfcoCANFfyXZ6FmAlZu5Nc/U4oEmPiuTBM
G69ckgbD6NMZzzPSeK9mOH565p2R2ta86QrdjPdwGROlYKWZrUIQFLtiMewUXeKd
mAMP5zKN1WXeD9SQ2QIuhvGX8Al3cAZOqSgGHn3O8gIIxsnlM+l3PJj3jnlXcZcQ
CghcL85AWZ1PSTNVHZWP5R2QK7lbDTQ4nQMCV/N52uGmiUPd7ly8/JwwbgBcjEea
UdUsmoBiXN5s8i1lqls6xViQq0gYDjOlkaMOSLGiDYiWPal9rN6wWZcawdMNerp2
TFCmVludt1TacaqAVGANllXltzwQWSmYtuFjJq2O1n3k4i+xoatHkqPP1d7GgbR7
AnBLaI0qQYlgESnghsAXeXBGHylSmqwIq0WovlC7UYvDDMFO0KscAOf2Ye2mRj2y
gJy4cygAc0e9ETZKyWdX7mloiau+s2/62yWZtvchX+yzqenn16LoIVYnvGvDmZYv
Wp+6JNlUh2ucSJckP79lzp1vUDWHpZlUvuNmq1epGhSGzsKLABTjeg0SwJG8APJe
IarZjvRt01FjpY3upVqEtQjLUA+uLVt6U6dqCbtl99YtmAk0JlsF+UOV3/BkXw6K
hwMoW6gJYnV8bn6lfpV4QfkAeWYxUEeUQA4UYTkCGpTAyeryku1SdI6PIYKS1LsT
Coo6UhFS5GEr2aCHlPc7WgFy9meR4wcspHXEr/8+kOpDFuGGNgByVTYu/uivod36
2VEOV7YVrxkhWh/uHkC76F+K9AncLpe/KY0XtYULS7PtQFk7nIRY4HedIDxcQAzK
sQfbAWqyVufj6b2FnwHuJO4Bc/MEuYsiM7HqIOcJoWyL3YLESuL3hOp2knVJr/ul
d/kHTFeqokvWwhssmqEz3QeXz+FnQSI7lcUm3rtbQtAyflnjXjy462ta+4WXSLIH
iSZ5HbaiAj94h7gLo2GC4iqC6ByXy6S502aJRerWvazkz4cl2EPMHyV7phFAlMlY
MCLDJnpVhhmPcHLqn8JzERRdz1C6Z1EptSOnc8hTM9j1xY1lQWm9K8P5HU/3Pzqa
vZfi5WOrvHvnzaIPnxM5/GYJ+GjZCb+IfO+7jAD26HY9qiGd3vt8rXsQJCdApRDY
TgsFOy9lwUr6AHt4PEZV8alA95ei/BqATD+mXc364heLwe9gl0rdsSuPhVQkj/xR
xxcIBp0zngn9f8R6XHF9T14CsZXslch8VhHy4k1EaPWh+djxVuh6lL/FiaSvl2LN
4skHnMIr2SKvQHZWVa9AssB2XP3g0la2IlMcEo6/2CafMekljAbq9C6rN7v4Z7g1
+6SueZ3PWjMZLDmY569kd3s7jgyjFdh92UTw3NKvlTFXGeLu2E/IDzXUxGl84CyY
xxuugP7lDKqg8HU4nZhiEdXqHCdjS7GOu3lyWi+dr2JEISh07vTVu8dZ2nv7Ei6m
gCWw7c9u5tRdmej6re3MkCspw/b6z1k/xdkQxSla2UZ6GGhqPXtvOFebZTYcA9io
BTaRE1BpEg6CoQXnaXp/C6CrdP8kE05K21f41O5BMybZ0U7xC3mX6O7K++aQH+RZ
GwS9ySWFUBzF5aMt+ZUri/hmL/3h+ql1/HWJFDn+9xkwFGrndxVSaDVqa0UVx/OZ
nWD+g+8Yf/cpKKhA4X7fBNCztghgxlLvgqEfPeeIbvzK+7rWZIu0zfUJ5JmbMz5L
38QuNp4jThzc8GsP+oNkax1xZe8O0eQQ7o0Fe7KwGkQkH9OmmnXASm6WVpVJmiql
CJkg1W+whHWk+jsgv6RwecmX4BNbbeWvTl9ZECinKg/thZzuTx8Gkp9DeWc1qwJl
rj6aB4O5jfAcxA1tCFk/evwkfdlcWdHqMJwieCRT23aI24Ln8imN+/jOiVIuSeGd
o2uuYKaBRjjGigM0SzuR4A+ifolXC45LI+QRrEYgkkQ6UxjZnEo4CLFTYa3jdBHm
JixxyjXiVi0zri8MmNmQaIyqqP9qGWjouOv+S0t4A+V6txO9JCOQDollwuqtMFJw
JD0AszbHKZOfMydPLudxFu2ENCwm+SDOYlwmaZS8wvKwxk9Ww3cM/bOY2JsXrlQU
1wJxofd16F60B2LJz1p6twOcgh962octXB3fek4Yqphg4LRKb4JrK5ep/Bm5cGJK
gSrCEjhKWK6pIYP7vFq+jDoNqbZ+PsmVdhRq7P0xt0Z9ByZkgY3TZca9t/HJ2AA6
fS9b1aGoVSfqXWiBQ7lR1ZtLVN8hNgX9iVo9jYb54xvxmD0bevzbxrrsKUQUiaNO
54HH9H2XClHpDbEbFCFGmXJbssq0FJcFoT36LFXx99vFhw1eCiOtL9Qb/iamBnaH
VHY6sZgg3FpAROXkPvvguIv0Q8NHonI8ckBqmiljDCOoV7jY3dGTH0Mlt/hKwuJn
mehteEqYAtQf9xJxgZ2g4we7B+EmIjmLTeHo1Qbbsd/iNlYo4UElkiBQW7mgV+UP
qqQHLHMbjGcSjKgQlA1KHx2ADYzMGffmBHHoloR8pW1c+VP/chmvwqI/U0udNgJs
KE9YKA7Hi2aibcMg8MJ9fZeyw2M2LNlktAD+p23/Vq3SPXL5a5n8Il6hv5lR6To5
xaXE9VY589G1tJQhk+tAQh17gsWsEWRtP7bm5zEcfz0wu0Fadzk9PWJIfmA4qMxW
mjvLoXwVwBBUO5aLN7PH6TYwVVo4f1YYlcTxlWByMAARgLjM+oYwiPmWjOcgosaQ
8TeNxyWwi5K9c6w/sGfkWJznM907PcgvUWmaiHeszdQMasybTyGs8E4s5RqQmS3T
KAfHffdqsNckYXxeWMUVYU5uodRViATr0JbS09pEP8oQnSs3EPN+KG8RrywNtMGZ
VLhP6zqgp82dJPofXo7hmonKNxk1nb8r3GQqaRB9sF4/3HDOvpCuuzE+QEiqH6yu
zKmEEQcvAMOEZEZke2kN42vr5WK3Zu/5/nnOJTN83k4S5BJuISDNzNmRdwWyL6Mr
6w5zYOtVvv1NaLE8ZtgjenwiO2Ew4lBJtmkt2kStQq4i1eHFriNFRPWuHrcvsasm
e6XdgsyrNrhcMi7RTvDi7nwjmOaOPOxcMHqYlyCH1vzXSDiGtnd4UXjCuE3pEWCW
F/qAMaTRYgJl/TrwNJIqDYm27CLhA8HmLSMTbI71XncscRLjzNKvgJfDE3pRFElv
Q0bZyia62+d5BNrocHUr2EvG3okJDxJ2mKRsidSI79iyrBxsUq7XOJHVE75qDmuS
XqHhrPzr/xHhE8/9Z8TSOszTUPw3HvhBv1v1YCDDxxKotb1q+y8mE/SbYaUY2cNd
prc00lGMomML64RWi+sG5TuwOpiYdR8GuxMwU4IUnVXuyRaI0GOp3zND8VBL9YfI
X32Qn3B85ZPmP3YHB7LBaTuEkgDHF+vM6UwR1FCwJF6kmI2MrV35v+YMC0uZb78d
5jGGXyI5xrfPCycR9kkKfbmiqPxVdM1Cn3YTBtoM4ADFM33ZEAyWoZrRvnuBGzpj
ZR73nnjoVlxZ5mkjZ/MYeU78hKWaVK1tVKBWiaGOAFCEFGPQAcBCr14jn9eZLhTw
wBIuLhqADCU/c3yVV+s7l4ZnqHY8lljU9PP806DJr3e+vSuYWc19RjGJHfbldsjX
LlzNidxSlpJuY9LUMx7biyLTPoQeMVUg8Tfi+J1o3Be7It9rZz9B2WrGLxXObqyS
uofAm4f1PkZkwwP+qj2OHj78yevkpMALAcYRBfQ3AdPKYn33vgwtwpKTRyp/hZZa
ZAChEireMIt1L8DbJiVuMtGy5gGtDtBeDdDBnGVwoR/n31LKXPENtAZhcRIvsUnG
7uPJaCTxR8k+pPIjrgXGBTsTzg+bZ7HzE/rHfnmWMtNppnNQa2qMUE6dwTUqQw2D
Q8AlF4nMTudkzr5jrKyNdJSJBrciDUbd7y67Yi1FdK4TfZJpr5cBKZYTNKn49nHi
KLlYcEntAQuPPupTOmFOzJeKFyO5G6Arpj3DHmtA6+a4z6NmUrJrt/Ly78kUXFME
meuNiUPD7x1+H49N1GDRepw6VQqK8OnTjVuQvv63KgXZi1hKn5SUMbL5b6v0SG14
8pqRadrN2sHvNsJflTDEJZSu9ejWRLz0AYLQzaDTTawP7M7Bkwkt5n+rIVW58zvw
6G8zevQiUXMYlqM0crnA3P/fRnd5HK34P6B4kvRhE3PZNa0nW2fk1pXGx8JJeEL6
Y9o6mk3JF/vGTrhVnPDp3dyzvMvedcAKyLQOo2ZWbyn1eSoKZy37aohJxPMoJR3b
J4eyn3zZDXraHMzHD0hIJiH57sgcMXHxtT1jIhBYiIMpofoaacwytCaQ22zjDuy1
Ql69QUg23wvhfKA5V1iw5W44R4TI7i36gDoFC7mhXtH0L3+VLmY5kqNTCIzpdFA5
aGAWuT1Qf1+40aq3gaEhp/ZkKtUe+ieR/LGy996qhNqXcEMIOFvPPVDT4XoCaQj3
yJbuCUhS9yRbfE7TylNfjaYkuZmjWXMB70lxaQM2lXPl2kxCwkov0UfhJ2V/DOFU
7CDbNNYxxiaIzoQG6Krq+OgAGQiVDaufN3/R2gRcBmSrfAMWQ4NcioaiGpb9vyt3
jQqu5TPmEo2gNj+gcYhbfnFrpLh/0mUkCYVAb46RMyqbeUi3kn7Tuf2LpW4Qqltc
udNqH7jaMyiZT5NM2TOhT9OGyTaWFybfGHoVfuKEjSJJqK8RTpe7IwB6bnLZr8hu
96PsRSdFa5W93LyKXzJJGXhumDx7Bf/QXklQxklX/R8wsrFkccwaJoXPoK7Q9Ird
iaTai5DtmJ642jpOMwUlrcnR0fP6FhCAbUo52caAMNeuuhbfEMxwOr52KeXEa5Iw
zHBrd5nNffQ9xG8vhQIAqEtqnu1AyXfqRWIRFZJLHKaayvKwVvX4u3TF8nsZiRVo
gRB99Z1mV1NMjzmiF8GOiOd6NVBvKRuzvuCS+fFIEc01imVwKMrn5k1G7KG67oCs
ls3QLAR62SFEL0c1/pUunV83E/rZ3ZANikB9FScukftEgbQCXxYD+qADveSBS1+v
Zydwco89gvaBT5cZfmM1Hf1W0SIuadKZSilr429ooncETkSGi3ArbGJGq1kGGAh8
ucsQeRQGVtGowhfED7rYMrFFLzyeJgVkn5NJrX+dG1hYEKtBosAtLHSVvBINBNr4
B7dhc2Uz9bcIhrt6fAMRYj6Va+2OoMKgEYNzMRrzpgRH4Q6d0BRXkFCKTQnqvN6x
FuCsjuTGVYno2CzFtehqxpvMh5S07fWXotAaDKfNjHr26+qrXjjT+bMMD1VpGabv
6v8rMKQPMNgZENv1RX+s1EVcv1kcA1bICm8gsCW/eLJTyVK0dyawefnuq/MhRfj7
bIsgOg6Gg0fDr2mBMtZdoqfTljB6SqTA76PWPw/wp7Zut4wzGLV8iTwXKzupKoeg
kMRACZ/eeCWnwhp2H7p8zLmGfCVhk5Co6dYseAJzMhxPWtIabMHL3DaDzNwHjZYb
M0s24sXOLiR4ksSWNAu6kkQC3sUbhfQCdg9EO/M+IKa4mc6HZUjgi3pkeycSa1bW
QwrTBNcCDmdN7BtpJaP0UyneV6wmhe82ORN7r/RTfGWCD71Q+LWzQ4AJEbxy62Ie
ZkeSOwuHqHDiFKT807cwsGDP20aZZ7lokPY+lHTSwYuR8lY97oMmubiSkYKqRK/m
mosweeore8wUYI5Ld2aLtabuTIxaSLBCex/E3/rtlhYhja2RbBAsrGrsuvtetR4+
VObhJS8/L4TSHQ0UJ9Y/7m8/V/7/csYIpx0NUMh8erGB3mxu6DchmX/fOdFLDKBy
q1ruNV4fdCdw4reFsnc5kGyZegtz1D6huPNSxSd49n52cGBtxg95GKo1LsECtk+l
TcqFW64Jo1Y7FQPleWWGONvNQea7ferppBi/UzD6+l028eZSED5fpBwz3xs59LVH
o6QKPa9FLHriQ+wm+YiM6aYS6NNGOdj0cygKAAu8vMkqSYGHsMNIGquRMsS/fFPb
DqyFvhIslFwhOgt6erqKh5aUbZiCBkuHVtnZnlCQmMRnZFeinPiuzGNoF57VkBQ6
w3hzLpqcTHmkLsUg6KSKz6h2k4Hp4mJE4j9M8/wbouscM5BbEuuNJxu6ti9+8V5N
yX1XW9URiFb8uwIAuDoGYsizt8EfulYXLu1/8hh9ev+NJ0Ab5A3u0S08oBVeieQN
D8EsrvUEtvYha39QkFKqvRcMzCEUZyfEa8ZeejPmS/s+noxe7fo8uqhFRjjVlevK
r1FLsXdYYfXUZUsEAcmItwg8eJNXB756vx+LEt93ANu2XYwJVKF8Bh7DhRrgtp3O
uri/r74PP38mPcrjnPRg2HlZUbUFyrIV2A6pgwSZPiXpfEtvkB/ljIDmueU4M+BA
GVFhVuNIpALfHGj3Aq6EJhY1i3tzpNZJNpUwTD43Srw+E0ZCfhiEVLsiXu0I18fj
5N0AfjhpI0fXwFD2N9Hnmi5xcxTdgtIn0Sf9LdYTHsMbdHaK3xm0io7b40G1WdLJ
ttVtxKRqOinyNDAl+0UlaWfle+5ZTBvX4JgISBvDOFoeKDoCVM7dNLiYozhcagKM
I5DLA/NWw78cVavwqOXnDytGAh8gzb2JFha3yg5nDKeLx1YTg86L3XHSOzgwiejO
cs+j/hPkV++OrzOnfdVQjfnQgS3AIXhyKxehZuHwruYBqFMxc62XSSItib6gCTAt
rsQX7BHYJdijnZm0/kGK8C1go7ODKHPdRsWaRAS6ZVMOEM+vVtE0AktMTTto0YKt
VfqaibEnRtPV3Mv8pOF8Y1HI/GneKqtQ7RsFM/kavl6hpwHapzrmX1kUeA9pTkX2
3gnVLgILzyZ0jgZelonF3IQEdyupMfVQ+8FK9Tk6BIFr5OdSbbPnOr6cgGxX41Fw
hkdemOP+MqzEu0CP+alLqBbUNXibENNPgefyfC3gTYzCV5PtGf2qN1WzxEfezAox
G4navjzAQBfsnYYRHMflDMMXvt8xNZt4k6gUcEUdg6wz+qce6rBcjJ0qXs4EVbiu
MPrjNG95EjIbp4lAkoL/RrPrtGCPbC/05ImeJvH1SGJM61bzF4d6R81arZal3Zq7
rE/wI9BAd41mktqq8xTQJvo2FHQRJE6Ducd71RYvhmf+MpimiQhswCJpg+J3aKFw
kfsLlr8saCcew99z5KYkhzfvesEQYk/t3QgHg7XYfFwzUMqXfZp2PZMg5pamHLNp
KwETiaRCX7/ozNF+vGJ3ONF/aU6M93u2iOCiQ5szmTueCnojRiTWz9BHJLaIVERW
9+BTGnvTzWcBd7O2hFnbPmL/kDMmjzeigB79qXUxBdoVAclPWMyZtS9+xyW1s6a3
qQt9PxOeiq/LvpVENThS/CnV75mi9rYuz1WDDP7ZMAQaUoOpA3wcKPqTqz2XkaA5
xtoPu7rImst51OMi2yLCbgizAF8+IFpLpVgwwkpgA0OG0NdWLF559JGUdT260o0D
bt5Uaf4c4Dl7lOFGttbh+5XBLsT9dpzXCe9R54EqaXGA/c2ufsuJnHIt/s0/kzTT
fQnRDodvLIVV8bNN+7ItK/LJorhmLjBwJ6IPRV0Q9PDrULSooqqfq5TZlNDSHy6/
IETkQGP5WauZTW0TxA/C0jXv1jmYYUpTB9LSvVFuFTOsEGg0LImOvQzjTeDjgFF4
gKRZI0Bti+715BGl/qmD+bFgP8Yuhvr+mKKdOkKU9S8FyhhlvMEHpZNo2EZRXZCM
t5+Wl4hlqyJ3hh4OFZ+jlGSWOhEqfZQMbxIjvAmHEOYyQJ54c96dBHKTAQq/SNcy
LxYT7uq4mzbvvfCHyfeh89l8FrPbk9OgU6RAzBrvz9Kzc/HuFr1YdnTp7dWDRV4m
VWUedCrPqQ/fDu0w+5zL2JVwWbWPZZAbTO+vQkN2Oef+oCr1F9/6KopmnfJd3F71
cuQoLQ5rKLfwVBtYftSJ2vVeSUFGmNzrqdtiYPU3yogopHQQfWnTQszS2mDzbIBh
ZGgwKAqIGLlz0BDk52/w2vhxbNdj7h6fAVjtZckQeLpfZruaOe956Wv2T0ad7Tpn
38fOPK+wNyynD520PCEs0NiuWZ9yDoNYqE+gHQkTsdEXGxZBs7sdJSLyLFZRWnNe
puQJ77qxD9ngFulIuHkfVSZhzXh2Dr8k4uJFLIgRKgfVEnsNiOSjuYe/S1PiU0T5
5/oR918J0Eqs1/JbuXB3J8ZlhuBgtXdu7E0fM1jbV5EML2OiNlV3MxeJbowRwfal
Oec0WoSkKC1O4GbsoS1m90bCtRrG1XFhwkgLwWXL6Pulb63Y40z8w5UQu2h5Jc2X
/fRTpdgcH2uIIfuHMwgPwH+4sbsRCA7dG+adbSw/gYztMOBCqGcND8HooqdTdaGU
c+zECaEaXl2Y5g3P/hhpnakM5+fG0di3lSCzEUSUxeLw5bLm5biOi5TLYg+PN3GF
ZloeRpS8Zs8dEh7CI7weM2hSZ130SiouqcwCc8wakecFvqDuy9vSzEPpyLcn/OgO
x6K/5jP7QKAhGDUDbcUOK4622E8EWDaxUJWtYnTkUximkzkzqmgeKlombebJsGMk
IdkLp3Qf5XBJhUI359/0S1kq9JsKDLBjFnp9I5Ue06mAA90b2vQ1fxul9N1aJ9t2
ISJQxqlyBlsmCKi9W6brC13fNHyJUVcshtd3mEq2MkiEL0f8uyUDYDjXQ+IhyCbj
mAws++VPoFpoojv6IqEAcMVLk2h2oqCmjuzx3HBXm/XMLn3eg88B6n0Yr+9ompXS
Zhp3vuUOfvWZt2xi0IFLGYL2B4ELcZhNoGuupDFzxXST1AjVF43fx6BqnPaZQ7Ge
IiOQRafSAHc1vXARXZdo8EBtxJEPR1ohlvkRIFsd+O4f1XBLgeGNRLiPNLyWFI4O
c0Sjuakdr/jJQuVK7x5ims8ZNaAICg4WmUt/at6kj0pv4vdhG0BHAXBMMU/FDdGU
U9Dmkb2DNurHMWNXyV4YWK7lqKmwByqpDPji4zjZRMDLQfDYvhhI04Cub05QOJNF
CNHKDbnwOUb3J02NWI2YgAUY3+oW5Pe9/k90LxtkxUBbtQvi/cAAC4rED5fQuuBW
G4Gbug/d5F5EV8U551nCefU6KDuU+ZyeSyCDnfNKJ/c0oYuoU4sN2P+RkxUTk12u
oNr53oraGuK9agr5JD2S5nBbXpzN5rpnDGZ7DW27lhxnLIcVuVI1Npf0lhZo+Tbo
pNIGy5965+1/92sxW67n0ll1H9MhoARBM5NlGmVkL8aHDhn+/52TaLys3CGiCgMh
Uz45KMvHVo7wZSBJCA4H6RltYA+IQmOwqsbI66/tfqQ8Htkk0YrLVsnn1Xhz5Msx
vxr8NwBkgpv+wPPzqS2hVu0GidRz1TFuA1YbaH9Y3QDlC1WIwNYWE//z2v1UXXLN
CjlfuqlJ0VAbLEpEOoFwYIF/96XDygc2zAMaFoaWBl8ctBelGY7CiZvwE92d6iUi
ivYkk34vZObcL3+xO9C73hIHblsn3V4rMjwmB1gGa6GCsxHKQSNWodyIVicxP0j8
KmYVey8NOonyE3XZd4R0AoBC+9Pz4hAiqTDMh1fDa7xOcHRD930BHLCUsg77ktBr
sxeFpb1i0a+X5GezcfwXhgHph4s3XpvM0ICneQduKRFUKd20jH981jDiOUcd+/4P
ZcBSec8v0I4QV3Ha3mMHxbCrz1aK0PKEpn2BznHBCYv8WgYJEYkAvuvkT7k/tROK
6LgMbhaIpLMYo4HvDOLIg6Md6O90j1SeQO607DYW/wk0DmbEkKduSQp07sHv3dyt
LxIYsQlUmHl0IsAJijZmOkCfSbGkOu1buoCSpywiJzdVrqNqqfLGY7G/CqIhZy2v
cjNB3KnG3iHnctc0RRwqF+047j1tgBen5PHHBcoMKe6DrgfIVxji16wPoBJzpUeJ
9Zc6o9ObpNbxwM1WJQxAu6NwBMXoEcLzwYBHJN4HUypGCVHyeNC/psHcg9fOBrPN
qk1FeFpfp9UXQ9qCKZ/9rh2WC1lrYCVfIAcaWCnGpqPj4dOQknuKoyinUgqTzcWN
2qcpdjhHcYb6rMZWqDjI3htqC7PWU2def3Fz/9KCElsMcfMMwqtMOkNCIAtGg4HR
LaFIyVq6HvStK71JLmJwnywE4mA3ecyeKDUQ+rdQ3Urh4fgVy7XHVvzhxKNGqkeB
Ce57cGljR+Hrr6iZr7O+TzRsER0ZK1GFyG0agokdeUw+zjczR7QrVwiS/6bryCBM
qfI/wmk1rvTMs2kQYQJrR2OCfv7wbgAWCb2RHPkuf8fsZ/2334ADujqeCN8b83tz
eM97DrzJMfTOgtdVS+MOoAiOM4fo/+Ok7pUKXptNLgyS+3JlPC8XPLFCWKa06sIp
Mrn4LAxrF04igL9GoDEKJe1aJNdX5Smj7qITYhkjhZPv7EriXztTDXInXntBMSKy
7oqBzgZ1UXSfFG3MInnf8W8sbpOXm9ytUKVIh/5rErgvQq+kRTLWvh5s2jem50Bi
58/td9Y8algjuUSzMNUberx9idMOVs1RifFxcLpJYHlyqVFuhzCJNaVYBzTUbzeC
jIdnHyINvgIR/URxvUTM+NFVm9bS2FXQuQN4O4Iuc1N1y/BYNCPDVzGUDYBNRpxw
DorKKYRORR8ugWqQX6WsoqwaCL27KviRhkLhM1dpO3zlOOEiMsZvkfOOcqq1SuaO
K4MMHVdk4rN+OcSUXl3Mm7v7/L6toIFvJgMiu1So0+qYAqCr3JOtcO4TOhmFX3n+
bdIA+Bne6BEYeMevkUgw1Nld+XpZBSBLgmMmWFeAjoKgRQeqylJTCY/5VqgRaoOq
Vj9jAUELsBDxsmI40OsvCLFV3bj/7q87wU6qB3gZufEl+0DvKzC/q7qmjCS0XGi3
PkeUiehr56Bp9Z1GV9LjtKSEN8cel8RFligT+ZzVgJlbEYgDdS9JALhdffTL7GR7
/mno3uHdW2NGu5l/fUUqiUF5hpC7rU3z1Xo3KE1vt1b7y9Wec+/gAgu1vvwSFDHh
DneneKE5vpNhgXVmYUKJLJfe8Y1g+UFNKrGYatiOVI6Tr6ttRr2o0Au6e/JIVk7t
7qJEa62itpyJnUNiB/RdoUMgj2MbtCrrcBicFG4OPFqFWXMxfrMHpdHz84/cgfEB
50cRpWbMfAiqSa+UMxh3eCY/HoAHZ2xbiGFeG7AOW9EAgcyAJ8nSXpCQwbg/A4+T
cD+EQSimZKR1DpkUzI+SpWaeftJYo+i1Aubnr8qz2+Nj+O13woZpDe9q1WnHukRk
5W76hgpU8XBQUUsHiMhbsuno6IY6tKUG1QQn+ETaHz8PK65KfKn5tsi9rojMDHxS
ZFiehuiCqjOonXdqmEWAsKhV1Z9mYTHyPa7j5X2LFXQrQFy2zMTafA6Twli4EjKY
9vUf1K0E7MU8Fi4Mn9ziRpDOjG8E65BCbX7MnywEMgxKhqUI7FQZuWLPKT6hJ/gc
KzlVj0sto1DX2WB/pXSgL7Yy3n8dPkHuJD1hzM2bAftqN1Dg/0saz/KMlsqUEMR7
WBkKu55WOp5gUDWvUbZEP8Xi7pVkSrGVbtGohgreWn7TCDPUhK56LpL0YNySQebk
bpdkuwkTSDjJeJUTeGCXNMmZtgAVyGYL00MIICJHsYz6d5GbJ+vQel1jkOL945h8
aLCgUUd3JFAt/811ANvqUdYnwtKvyuLKza2JegWoBDXcbXU8eexjsNmVeb1TqsRF
5Lkj1E6f16Or+WPtTjcuL4EMT8mXrwIthEeVPZtaTKlHrU2Vy2ss+m7zIDhBF4/j
NpjRh4tCa8r4ry3ICqiBVRpuF2KIEz7EX5kSN9oRwEX++ZI8blARHMl32ytnCIuK
ejpge/JfRlobEJLcHmazf84lS3lvIjVos1pAGWFPSC0uox+TBfWrmSTsk7YzWoLg
zFOJsSwcGXrs0AY4zg7UFs967TM1q+K6rL3DfdbpI7sUNTdcsSsUCEb7IkTKwBBy
1lHlAElq+dOrbJThHdsQQ6Dmb6LKJl+SMIiybXF9zSZ65X6CtitmfzdlG7iNDLoP
tt5JegA/dTq1EuGV4hosmkM+vWv+R945SqCONwo3u153WAQCYjWnKBkeu/De5ZkI
tMdHWSiYhyMCFl/ALp3sJ5X66lZKpxRfAjvcZZC6Rk+S1KOjK8auHaGVZifQoX+b
gjhy0E7rnXFWnrBN/yS6+e+Eb4R+a8ZfdS1s2oyt+pBzwFRpLXCzWFOSttftHIsG
tNEs5pzZUBBvl9U3Ump7oE09nmUQFLBFKgQcLWCfL9v8Ob9eLmeSV7i5ypL68BUg
RFT1FnO9l6a76yFANa7BbKR39hBFaXe5rTWRMRHcIYFTov/oLktfalxHLzACL0Jx
NGwvKJSapHUuCydlGIyBMufBXSqNeS8HQ3zo+xRgFvsR1PkIEEtqsTYw8OGKmwzx
0N2LAbBiOYmB/ky/u9Ly9kCYPh55oSiVLTEvF1V6u/4VyJJgp/yV96EjrKTjD7P0
st5ZW6o69GoPnxcW2z2RCXvWfsWX69JDISncIi/CI4SF0P6EO0jXntLMeyXgrIEp
6ZIOYIaRw2Nkqal1w2PJ3neDbynCMumkKAAMimeS+n+uSGzgYciMI5YQfbPYkF1Y
R9hVV5FPo5bBfhS1HhMme8k+YZBoLEitX4AXAeNanFkskxnbky71rb5Y1Bdj3NBs
zdJLF2D+yUbkhJzCiTRb7MakDRFjQIjm8YNqYhzSIqAlbUyCKSRgWyJzlIHDfVp4
wyJaYWc2CGVOzHszwlY1k1wEQisYEVBgjYnR6pKQdh3AkS2Wzj3bX0LlnYHgifUI
hk3AcqayCZ47fWkTCsGPNsw45OHU3n8ZBkeCBdGjcLTrYABVinebtdeQtiKZnYqA
gTi6yf2e3RcSXIcUTegLFvK3ABPc3hNQFPH9bVyzJ5HQoEX8TSHwtcuMb1KNI0b3
8MLccWrlLZ3Im7KWHJ9dz1U219dXUrtK532aSr0dj9+p6Hz7qtEWB8k/LeXTNy+s
RWQeVNa5mqF5hq3zSf1y3VKlwQ4lOoni+hB7QfUZ3XlWywY+5DKostbfMdCwNDGa
uzSKmSOp6hy8E+qTtuF+cei11tzBmrpPr9ePKjyoITam8gO2wgIztsEQKeyGI1sq
jRx84iG2lUMBWwxPhiUCl2tO/cMuUFI+YErYjf2ra7m7p9H1PXWJaA8lPXEHjwBC
/1kRDj06zaFkZzPnPmdy4rkJ1jQW9NqUnNR54c8Lt4THAYtx4D01pbSDjs1+19t7
+b2iBs++trBpVCMd9t1kgdb/sz6ZggBn5nsPheMkibSeenPHh/v4quL2lyiYkUEw
Athh/ThYV8Z9CTlKPQ1Fa27rIwILtY9vmSHdgsinC2wccnaZXz6XuKLv/W0YUNGL
HHpfLbAY3SN2KiohTOPDZnA96moiUZ0NTpHX/a0LXPz4qe81vBqrmYJX6Xu3ulVD
vdKUlueatymrrj8aejKd146gU1hWp5ht0AGNjQuG0twQPwAK88a0krfXFLguCpMT
SxPDsTfHYXt4XFN+jFLNxzBrAxjygEg903+g0HdhvYzPLoFpsV3ZzPqcp/PLSMdv
7oNefvFlnMx5TBn0ZneFbuzi16VtqKYBOs3T5O2BBEsn6Z+xkGcNH9RafujzbFog
5hFfP7pcfOWxXn/WLQ337bCx/rGbgpCs88mPtzVIsnwruBMP++sK4MF3pF6sycc3
K2z8JHEfne427fwovonNOMN1HpQxW71TaDLwrW2ZkLJdTCyz3XSydpsLieTELOBK
qBoYbLkWdeWhVXQFoaVYlCdp5a0Xm0bxICCdYT/oYqh95S5ahtW/JzsKU/Qg56xf
rtcvwVabEh8LFDsiWClnpPzJ+1FlqPLs9Pv/LCC1at49Dvf2lIKbE1VPNqIyU/MO
Kr/RUGpgLsnUgqrVqsG+HBeBZfdF2i3Y2AntbDltrLPtmAtq+W/RW3Zp0hjpqCve
wz/RhA3KU+DvgD1aPsZNppQo+oBr+wRleKr1JkbYzpu5aFE6yxZXz3RQjnv35tcD
qK2QnpVAvkMRoWKpw+6VYLjFS+HJ0/9FaV5uyYiR8OPqzEYh2/KBJqrBr3aSHh0Z
LhTk9q9cYAerWXDRnp28Dj6ICt/tgGN95FTHyQE5lvsaoER+6BfiQ5QWZI0LTIsj
G1LvMjjJkzP/+r8rVuVivn4inv0+VXp8EVuJNlypgcEdWMeHQwVvdHFRjLQGR9OG
5SriGEEqnn1MErHQ0cC8z5kRokBtMbXimkqMmY2XgH4UKZ+JxumKl84RUMKWbwUB
eK9Q0RRkJKj2ai/wu+tYRKqx5pN/s1OCp/rQhoSFrA4Zlg0UpAkswG15eRIZ/wXa
Lb4eMpC94uR/T2n3OfR4g+1+uNDdVaUUubxGUiTePsM0H7ANLzYRDtRXHDR7dDxM
rquQS7bxhh5SWXMtPRkdAcZYufVYwYWlGDh8bYzd2PN5ggvlENMCfUJRAov4lI2i
GHjv0LC01v2dQkJyxwm+dhdkQO7RUSWC00LPs/598mQJFgFKk+nEBwKJXRiy5Chl
Svwu97PSiz+b0aq/tjYs5f4gJ1p6XHrClvxYQ2aOkmLbISth1/SjltxB/yBJ3z6S
kTRMBL7vtOGOR71/F4lWp/maaOl5JR4H51Xcp861jENnJ+jhkHgKOHZBRxV6aCUS
T2Y5OEIcErT9754Q48sN8BZxB/Bkd1tWnhdH05TKhWZOUh5kPVJDLQ7KP3X+pAgR
CmEs6w1n7V9ZrBhPA3hedDMC4Q5ILHmcHPQIvT+sSfQU25bS7uRVTEdkhrO8xbbT
SHAW2IzncKI3IOWgWHSsbaVglmFvRBFnssT0y/2Ce1j9KlGhXyzAoZS7FAjTXaG6
R2WvN8UmHLBKI0IF4xd2JI9n8F4ykv0FS5idq5o7TQfKOtQnSpUlMt+bdQb+r1Jl
+7kfZQiHZ0+5UvJEuDEtqW2lGs66L4RSzRGgpaJblkeqiIuCTsG34opTfjCmEXCQ
myGssCZCSe/5qwnGtVG2LjOFRTgAQzRpxnwZYnemGYeZZmltGFMdjHm1SLs11WQo
I6Fe9fxH5yGZ4KzKtwtgm0i/YK09SXx63xg1jnceMyELLoItjKz9bTOdfLkP06og
RE7Yjx/LnzUQU7d35PEY4rtkA2OOPdmGbM8l+KXke2uEV/Ik90Uv7HjjfoCWYLW2
UVQrE7AXZC74SaScBWZdfFqw4hVUAnnprudeabYXS0fsVDRh10wYqBpidR0TeJbG
PUXhcKY9VANRx8uIl4EjIUP5EzGecg6T9Qc1Y5xADSBcg6hwb7vxzmEqgJ6fM/yE
VzZiZQGjBKA1OjruvWRgbKFKjE1e6v6xyxHDLQ0TWyf8Sf3ZXW7W2G09VQNPoJkj
PdOdIgUnEhPCu6ysSOSFTpO5eK0BFGt8MQaNnXTF9ZMUxovZNCabDpKB5NiNrs6y
bEbsrNv+yY6MkyNqoE8EYHpQyxlcvXttLZjOxss8X1f6ahdyjK+Ci9qQG2xspfWJ
mTQomkMq9omUAx83FLVjzAT2zGozVzf5MUKjzuZu/NJ1a3nhmJVToNZT5dzmwWFH
gcbF7TqRIHrmHz3KLZHkJrGnf7m8a7uuJw90C2L975W6pK3B84zczGoVez3Pn4jo
QQs0ThdcOyo8I61Sg1bmN+O1TAohjwYiEk8JSSqcbqqvyRbBIS1F5jUTZieWfnbs
CNCQZmvUFo6Fx4NvW+H9p3gMnAn1Lm1tcskaep99uUZ8RTlBpgMxhw30Z02agj6M
lyVQgCatwxNxCLi0a0/rZrvsXEoPYhaEHb6AuJLXxgeE0Rhr7uqrA0Z7xml9sQ11
MmUmLqyGmOOW/9SRTiB64GQ519fF9OMoysL+JQR1mcTXsC7MIs4PKSPsQoJgVMIP
AxdWdnysWokswXsKKmP658qbHJNuARfntufDMVPYZtf1BmGIVOslImrIhsBczZPj
myvyBdqMc06x0XUsZrqcW9jRLEj9r10cVXdVMJWPrFlYnDzO1uRcRXS8ZCulbgph
T18yz5lZrYqHxEbgsnw8KPETpGOYE0SAi0QZzkvGpmy4jjUKGJWJ4IDFj5BoHFFR
mqdmH+lS9s6S1jZxlX3qvGQvU43MLZcAMAemv6eJfJOPAr1bCalt7t0QT+94AeMR
UNJPY4LtBO2AEe9AsiUPvt0RWP37SRNkJ1zvEqLqsOE75dY2Qoy9dBPKXcI6mpCN
a9xnQ5Tn74/yvy/woN9id6MhU5jAd/RQyfvBDJ6OhoZDagOoMboLvGwjtddircYV
ACjKrB5DhxiFsWST3iX/XOHZCsbQ0GiBhCkP6p3PELHbxZFHZxTH5RvlfWmBSiUS
iAPFm4oqLHIpRcHHMZg8KICRR9uXxcTO8K57KZVJa/ocm7RaJ9/e6L4jXxEyceJ9
6aZxlJY+jpTALAu4kvDQOvMZbCvD85whz3g8KM9gNd38abTiVkVUIS4mydWOl7OT
qxvToy+tmNhUyQELe+AKpsiwaidrpLm+eLylht44SSeYmJeJLVNX4bj97ygSzA6i
UqOIcjQI/aF8T3zv8Nfa0t49UyBSJKr/7OT/FFiQa2ZTZOC2VPte1EmFyvASHSHx
Gm636wUUUvn66kJhkxyzShnVRVTiZLy5UVjVp0IU4fpmyzUUxaPWuToVOl6Xv9o6
EVN8q9xybFBarBTBYPWNwsITS9D0k+iihzu98e68ZnIs205sNZg3+OSs0arzn6Kc
aPzFNmBDcy6U+UDquMPhG2Tf0gUeI3gZ8KP3dfd/fg6z1kPuhs45wmBgspLbyJrk
Iop1ScRjJTbYn7V3fsCqyJoQYP1MOgKvmi36J8nby05eON34F9bnpKdnvuyEqqCk
s1SL7JB6tPPZtUvU+I70AgF3dqz0W9VszmDJZCxsoJTj7yiy64LFwt24n+40afCr
44TQzF25n+BEoDgEDeu5Mm6BnhjRmnnIyeMNahCFJbBFm2qkFW4JIbpZZN2d5iTC
xFD2eTr4zjQWZjMbinXWa1QqwThFIDspcZGhG0xZIf5aDm9zOpAoBPEjrpBqHEVZ
m4nFkV1czxYyNMR35w7RwN82epsJC+Z5Qtpph/te2E2pIHORS95pNtmYvARi9rTw
ca8xlXUJ/4sXjwRMFHMNFQI41KfNAi0HvqRz5YbAEv03bcRceUsXqOmfmsQZ+y1L
1IPRh7z8g2qeGi/mdH03atVYmifDwn27DJEZOK24nIqYeRT/btz6JUj2RjeXTr4a
eduaP7DahUSiQfJX0ybX6RwlctogxXPGX7QcORRhfqg9HTpc9dhOQT/khf6v7icg
DFaO8vx/f2u+kx1U+PefArlPyHagrMJhxF2xcqK0Z7a+OBovKOcXKbsGnrWSAl+f
lB39SDq2yHJ+NRLIZJxVwydFeCG/uqcIEd0SY1HWR/V5Mxbhzjhf0jIcHSEOO5p6
ig7SShAyRIY/celcqbBm2pT+dwIJIrZQ9vM0g8ieFN7gzjGeQGzbEZV058KPznX8
lzu2cC4CtKNg/+eLe/cHR4QaEYTy6PJEDvCq89Ml67LMr+WULj8p89Xz/kee85nr
Z4w0tCs5Vz4LE0kBS304WN0BGx+aZyNHrGzJESg64BpFX99pv4CM3s8FyQivjmFa
n/Rw+uZ0mvAVu+BbyRDb7w1WvGu/1zGDXdzZRxCFB2Y60OT3VLjK5OtUFcRBQdmK
jl+VwiV+po0fqQoEQ6j3FGIzAMMWxZ+9u+CLQkcFMIA5YmXiCEPosXkqtxDrPaPQ
Mda+b2rVJfXUAtlJ6JThHZx2+4e17sZu/4Kc62HkNkL3WNG4ouuUe71MFtsBOvE0
L1DaazX6oQDqhz/rCAoTQk9DPOtpPHY4Mz+FztYxOF5bD98XwjVjXXUWctzyXD+I
VQLSdRYd3sg/yDjXx/Vz3xr1U0MQJRTWejrDiz3HtE+Y07bE3NXUv1o+QjtRDTCG
Pk0tFCBzAaHGoTJUUW+QBeTEkgjQNQkj8IfTwbpUrtWsSVgA6cTp8WAwBIQ0jicC
MYjUnUskvsLWqK0gauHz6dW/YTMUT4Wt155Bv/kFC1EA7gpkXNuHQCatOqGjoCDf
lIuu7zSbAcDXJpEjxkQWbEq1kybMiZqUWtKke4jiRcPunNEsgVUrJr0YGYQt5lhC
xW99jtpjgkDTPyRBQ8qgten7eZJYP0+Kgb81JsxQF7L+5E7BtI73QWo8pUCr5tsc
xcgS+UQKuSSNN7xWuEGjfS3nCRIvdqSSLAAm//P7ApwsMCWrfW9x2h5N/VEd343B
33Xzfih6Vu6DosidnPRy+ETJdRwolkEyUrxGi4YtWqxIjXsOtYcxzjoRr162V1i+
0YmSf4GGTuhA3wrZceCCty1r5Q3YoGHT127RRu7I9XELQnAQGGs/ambeZ8wYMYz8
8HbxiSZzI9RVduo0MWXmq/kTMrNxNGgO/nWNDnK7rL/da+GlNujFfakV2Q+xvLkv
W0l/gLWLiSQHZqZoR8MJLRAqNzFPvtWJkIPmCxtsd5CvOhK4+x1miy0OD6MLexNu
YCKoGH50dX4IL9HDP8FbAPP6M36GmESZOyBslqJhMPDY23jzY7hn2sWQmOAqkx7d
tJwiwkEMet9hnbIq34FqclHuABNyKO7T1aAAdieJkJYzQMo1EMdKg0mfGsl9LQZe
TkqjNDF5+grG8ZwmDiuTMZ8XNCZz9G46RilP3/dxEfcsGwbKLPlYj6zvuVxqvAip
idqvIMl8IAlXHfBS90fAfuwbICyRGyvAvtOFnGmBPSa+tAE/PSYD1skk821wryL5
+lfG0CkO24tkY1C1Y6y19zeVmI+GHgqQ+yjb8ZdH2Lf2GyYfRT2yJvvLkg19Llix
+rraFthUzOwcUQryVp0n+DKu4kOwpKBEAGLGHVha2hkIwJzvXlQmmCRY+aP9xVFa
hH1nNid9MWYqMtnDzpj3TIx+/nwxvGONz6LawQpxroJgvJkkYaU9j/zVU0gR23tL
Y7/AHqXJHWAfoOOVvnfwx5mm0wzoukaVTD/wwp0b9ob4cDJASbQIc1aYM2N/p6y8
ldFYd/a+aJRoVs4aKDYQxiazVZ6nPBuLMh7gxFrRjoTEwGUK/pL1U7UTvnxHe41p
SLoyipOdrPldsr7wBJNCY+hIqlZRv/tRZvF6Ee4co8QKtdiIkLniru+JN60rAIMy
ilJtTunizF1jCM7I4BvgDDmvjQBN/X6peEPcIeZGv35Eu5TZe70I0O4DlD3hbc2/
NzZzT7iJEmHJYYQ3zzDLivBuhlNyNpnEvaQLdSiCgTtnDDDUsNfABXdWX+ffr7t+
DhGN+dMUrTdYzGJeBSZIwrKqRQ9JgAHwHrgS23i1oJHj53NX9uAAR2bVWdBi328b
l+XYELj6g2k4D4glHDKKuoO09QFbMvLDHOq/6q7wXvVQ4BREXN3uLmamP21IHZIX
SjVCJ9qDvypDziAvWKmX3DLUbl9ufFvD7see6NUQJMxjwm5rLfRpWEA8MQYtrABj
SNQHhIR/gsIRixhlJvy6vkl2RXgn3pR8wREo2SvEhOat7AAlbzibHgfFX3faybos
jj85Wgo13SGJ+ki3yPkv4dpw15yvdzQO2li5VOEbu2CFymdh/g84AQrI9AwsiOZi
2va6ObiWt+1+e3duQY/EoM49KbJo5fN3jsDLkcTW89YVyR+L3/Mv8KVmHuqcSl9q
jocsP5y1Iikvqfe1EPvuanWJzCDf3hhFcRfpW3Z9fnGDO32crmFtI2i0xAVvXJ6U
po8Vh6QaitRAXXy3oUOalhPfRDg4LhLvU7npXjCDNkHnVhCuwhynQYJ07CfqxiIJ
XeZMtjm/cP6kdBHHaoO8lGs6FgZf5mtPzR+a8/RSz38plaUY5AkB+FHjzoLH51Mw
3tLVzZUv76cVPhHHxiLyPKuapVOU2B8kZk9DAAt6te7Az2XAkK1LDjoo74SOa1Bu
gmGEuTot3W74lZopS77FHS+TQ0YpjNl7Q2PC/qYaTqF1Pb0bNlSDTSH+iQFm6Syb
4RmXsn7SjzUVQwOOL+aouGGh/WPOsWjz/RdW8LB0w7rrX0NgmAcigpnEuLfrWya5
dofaDlqZxLz4O9N7pzRvUQXnn7eXXAoGMaqLYJaOA8lWrBMj3xPZDScvYqHzVvQr
kwLIQtbpdvBBnytKbBSFblfFK+r4ejJkZY8TrgAxWsA4LJc4FJ5mqat05NM5KDAX
lPHHinPKQqlndq5FEoCblvuHoB2ymGwcPRwv62ty1cjTSqWhlYRecAaILgoKn985
s2FKzAKaDyY7MPut0/P+ol+H1iM3GWl4ftg/cUv0qxLnCcBcoYz2yW8N06N/gEuf
OLE5cBfncRXgPsw3Xfx0LucczqCDxGDTpO3hIDJYawwHgOdRngjvAmvY6sA8GKqv
EjHFDAOYhckNSHXwqFoWySikjlA57oYMG8GOBpVODnHQeXh/5sxRZQfPa2X04Yq9
M4Eq6hoUXYXaQ0pK1AoE5yyfIIrWQXnzA0JxhHiiQ3LynKD2MGhO1EQi4qRnrDis
zqyKJH7TuYaiwDXr+uxcKnhgSIpE04y5VhhsLQ0dAeeOPg2xat+2HKqggx3zioQP
3I3lFrDnO/Cm1Jipl4FXzgc2ewkPeD2e3ImlgCYDTxchyCPLs5ZEtWw244N6Sjf7
lB7L8CJ9jmnd+3Vg+u++RiYrqCVqhXOlfU6Cs5XC4ux7FKDPpe1YhfAD40InlwGi
MJPpRTZWrSYSw1r3ZQn/jH0qBfn/KKqFbII5S8kFVSCKLEdlxhu+g4M/cnZluToR
8q8ryohvfD9aiQtL68N5hcl5/Mrbt6tUh3FTTr8AqGOgth1NQwy8kUj4fDVo0Td9
KEf4okpKfdwV4OuNsj7x2t9rsn8WK+fOf3g+/A+HyVHK6eyRr7EYhytau7x+Qs5i
FO6gfy0rl8WUxcqj2Kq7iFXUKPki2kh54JaKBi0zdfDP3KG26nYq64pcypiN5Ghp
/U1fmPiXGSNotDNjBB7kUEPH1uceio5IFDsz5/+Hd4AvnHbH1R/wmTAtUKXPF2UW
D6ssJjy8NgC5tKQsyuCrHRXvVSYNCD3A9XsOZR6HpSmpylb0CoOEB55YT2V36lC0
M3+156UMJGehs13xHY4/0O6NvrPE26N9nEEN61yzVoPuKEEvZCeuFYZbPVh/WSgo
1PCH0mSSN/3IzQjMk58QyQgsjK/d5pjqcmr1ToFJOSrzCxXxm9kkFHUxLMCyVNDU
2/IdWzquKYaIJNDvBz8BD070nXEzl+HWt6WRjRqrJVbnDrHHiNFt/Uz2bOwjrw+F
7SRNXkwqPQidA1Zp9q/hGvL5XM4tCR2YC1OB9clQeDMkg3ASkgpo+tXYLji4gFjr
pE5Tg5Vy3JK39iAm2lDZi+D7klRulTSktatWJE8urI/uSuEblTHRM9D9w6ipO5Sj
tltOowy7rlaDU7/Exkb02q0IFk/MCmu1HPUcFSoUjjtb/S7EezQ50ASpVKIA6b8S
cAvjVEbdlKONtexN3Hs2dBUFISZA+jVHRnc1G24QFrsRXRjXUJ/dCrAkdc4RZibL
+ak1YlH9X0Y7LDLSGVXPvwIqGfcFCEmcHlBS1rMqSqa6HvFAR3yglJVwAMNTsCjZ
so0JvEQcNBMDFv+hwhqkAs4lcu3n4VU+SGlN00YpUv3iXKVAPBusWgtfajF+O2u8
dK6BjA7Q6phkmR6SzQXumaWWQMkglVXkj0Q7xEBdp7c1lOxXe/jfftB7DXAjUrKu
iWiV0vEwfOyymyicwT+Xa0Zr2BqQ7wUUMyXkvmsDNHHY4b+PPMxE8a/ZKUryKBWM
HqhnoGvphwmTb9Qksyzx37OEFUhhqWNACLgTKaZbRfe/LDYnkfdtrpsvhePI58nU
J54saSD3eJMiLZdwf9FDiLhJdBGJ0/7t2j2aGHmelO3yxEcf3Qwb9DSGwvweU4jJ
SzRYXD0mVQ9JuAK6ELJphZIt30KnzVVI5TVMXZuC/4uzuwWDAqbpBkEV/NRcYUmF
bbD1YdM/jWNscCeN8T5BrnWKwgIx3DJm2Zvf0E+g+MeoSZ0svCBoIR+tdYc6Nwno
ZU+9s1ccDIEdT1AthHfLHGGraiSFAqNRhcsH1PAbNnogMVCiZ1DVvupck56+nEo/
4T7UihjXkPRpN7f32reWjQS+xH2aphzmcHytrreEtCfyWvwkNiXzmkGTdi26M/m5
R9DTiAzATCunV+AZ3cBAvK3eC1eLudl3id/chgisBfKRRu4PLtuIgCwxt3YD1rC5
GOEsuIFH6IcCpHufzJJ3QrQ5cxtxIPym9Yc5eZG5ZkoGO81UTfC80LVG6aEqm0SJ
OeMHooKMMBYx4Oyhg3gyS3jECmhSmLZsM9IyY4lfZJZ9iqz1KNcFXD0zZJzbdpDr
oCnGAKQcCqtB5Mqi/IKUrlcWSABzPtvBo0bQJlFh65oMUUfutS/dzWGpuAJ0tt/M
BEh3s3n5uvLryT/1Zo0hpWPtBsMKQvXlg11sY5DjwMP5le7lkik7rg40z24hf9K4
UMfB7gPJdc4rcVjBjTiwUD3f9Sr+akbUJyPX+8aiUfycu2NG3KV3uopAeWRv3ezZ
NzJfZ6SNVWhaYNpYGg1oy63CwgUwuWLi+DqfuDnDvg8azy+OANDij8Bx4dEDiXOZ
YMp0wzE7WfXz82EYJFQaRl9TxOJxJZPQ8KVzCT07+iCsFbwOclw9MLrkqAqWK7qF
Tj956HP3mY0L0+/aqUqyDtCnBArmqso7bKggBkCknU9/5yCIB/UwrnfoDOWeC+Ib
J/1vZ5nnR9wQDTJ2MJB0qbhq8JBHtIaa0qVqJtDtqu2WfYdlxHluDlVKqV5idOWb
k2Vbdpq1XPz/+9hcjxGCoaAPFrvq6pht09rVlJi1dx/0ZBN868XrlyW/erx5YteV
zhhdlujJMuRmLLuE0qevXXPZQCsK7PjJ+eXz0G3VuhfNoylrEq1JSAQKdX2UXnwT
+4EKPWYTMT/pVtACAc+6dL8NWpCcIB1RYphdzUkXzEcPBiPt6oAcNJRlgPYYE3AB
S6LsrGvkX2f7t9zL2fUWK2muoRgAuyK58aMUWb15JXZzSF0Aq1gGjuhPnjnLbhzG
todzCEnosf7yHwahYmHEFZoxdVZmTQIPGtl6xVZyG6Zy8bu6MuGnd1CEKYLcxFg0
9SOQatelNLY6SLaHDMdFsPcQTHp1VUf7GHQGSYaDvTiQ+fvMuE8dHguMS067Pud/
QOOZ8E2PZk2g6rh1rQkQ1PfbeKObyGP9pteR5+eL8ALFhT0IAfLpyQn6WnsI5JKR
s8EmBIwtNGZy09eBK9xmfkiFBG4QOPneFrbpGWvu/PdnuEs4wiSHW2ZjknLTtpHC
aDsGBm73esUOzRbufWqY9wtPuJ+c56R8bYvw2/hogntMhYJACuvaoK5wyhVutrz7
KcfbXVTZ+GKahQnxqHReEqoQk8grUMjFKj3vkoZBRMNB6TQjZEMLqj/3dxblX7an
542e5/AQl42l8ZLIul583dIBJ2ot0TDLaXm2r/LzmVrJCpUrk9IV7b8vY9dF1m4O
6SJm+U5aSDstjnJU4f31JCXWIBE8bXo/iVlRE7/VamqU9VSg2Y2U76qbSPp7j1cI
bC8sKXYsj4jbxPaJJn3XUo3Pnf/34HupIaYD8lE3T9rlB7BiFefD1WaZpJ4uahzj
L/fBVdGUN/9pZlHCd79c89MQchtlk1vvM7CecX3ngZKM7zGUN0qe1w7mfhRLE9W5
aoJy0VDObiQORfF91TnJ4ujSsBW+WMLRuwuvv3FuePLWeCq+qedMa0/YyN4xcNWa
uD9Bd4OLOEVXQXWQt5YEnUvk0Fo55mRU6hFmBpJUHhXhPmU5SVDtsDEogcH3cTuk
fYAxdAbUT7Xaxo4TLjTNKL6qAt2ydUR9sgfBD1v/OBG3U9DfjFHiiBq1eJZ++y6z
C8xW9wkei9EJhFOXwg1GJKS3jbV7c90y8ZGXV+5F/6wXPViIUfWNHhg+i0hgGD6b
FNw7yEjZAf8qLq14Sk2HodYfzHEUvsU1MpverFbCxPjoJL37/2ue1K3e0V87jcPp
zOjRzmMkgXIzXPMzmrQl83YqIUWeomlZjmD5ffTcfTmLnhHS3LB+otGWNV7FET8L
fIFQoXNBGuTpKjc7JchrceaM2l1WcDnWGANuMjnb+56s4CnL660PcL4g/ioabjUf
Fl0g2LcZCpvDRTvcwXbIk5jJrfbFDnPb5PVFt022Amt+opgPfH2Jv59Eiz8ovRsk
kE//2Y/fjkpwNEBrO1DcI7snyKrcO2WQUjjbczwPpatU4a5uhCmfy8Rs7Y2/RC5E
Aqlrput37WVPVkEW6nOZYIbP7OKab0x4Hgd7fvDii+KASBZLN3BUUoLKOGOpttf8
jV9MK1k6CybiJnEDKZp9RANMdHBbb6rBKCuGOHLhOfZ+VkDgXS0Wb/y7EUpXfvJu
sosUbqhKbLb9e7ifz6r6c2WH1Z5CpVsb9Ws6hJtStFMMHWfjTDzF7UjBCodUC5w2
eLD6UANT46MBCuSBvTVVDhn2FbnsPD5aHaLGES4ytp0K1YIbIG8EQDuYXxfK3yLJ
guA5nhay8rLTIvQoH1dfVo9D5N2d3CiHgm/wvPzTk2Ibw8dy7wDaEID4tcAYpVKg
MzBqagEWG7D4/gUxxoLFCppfNA1XcMpRCb229H4H9PnQAir7poWvOwY3yAAGGAqh
8yU7cRKEPmBMH7v+wMQ+apfgzYS4WRBEPbNJpeEc7Irkl+B3l1na4iNTEPpvmTcQ
3XcG0OJvFRKjKJu+gixOGEJz5nSGADbIIE45EzlLygbKNgEGoojgwnZkrz5blV3h
syfD+pt7AY7cubuFkCOKyXgGRCty6Z5bBxf6othiJJm4o6wd9ygoLAE1LRdn8tF4
+Hr8gQ1h/7Yt8WA1lnCpAsdfh2gpbPNH/lFPWKzA0sQCDqvP8po1pCXR0kHIYHqV
bxG5OPBErJ8eb/x+c/+zJMjw8UGU76qG2yDfpiwjP/qvcN8daqS/8oCUBvwk0AT9
13PRUpkAWFdwiCATikXHT7EJqjWSxNytVjWDU0QEXw2zNkXzaRMXDvrejPmPLVsj
ZPR32nfLhjyv9eofMKjsJ9BVyO4ESBmn/m37+oxUoEugtuFqFJO9KdZLsQlc0YtE
S4MXSLIIKdcGopg8zy+zQOi9v0JDGTi5l+iXfkp9vBA8M3+DTzKtocULX/WP0ble
Cu9FcD2H1IpZrzTfe+49k19oKsZOl2zQV1fViSJdSbBzuE7BjV81ugHb8H7oksiS
lji7z6veTiv1uZLDLU8fBr4/G84m6zfTBz7CNOjZmOxUrNwClI/NaY0yIhRJ28re
RqrBHUdp4Bo4g/gnBQNJakwzZZe7xt6uOuFyOROjup7nlK1G1oFH8WlTM8bx2Whl
W2s0M/b2oTcmE/+jxWuZLK8jfh1qvPzug46ANWIURYZA9evY7/5zEmISWbgt+5o3
t/ldGxGwtYg59RaWD59FTdaB/FrMJu7YGNwSDAG8HLLDLAnbTyg8ByNwlZNgTxu/
ZJvL97NjidbdJMt5MuE2NJkoVjIwVqsQbf8FML+m8v+OaiG5JW5BaeD3hs+fvyPG
cYhS/enthNtS6jfMnEh+FUaI2Ewit2e8ma6NZuQ+Jwpsvdf9uoENKNIt2M2dp4wF
p/hqRynZYFxcibTLv5g/lGbeVXGa7rF/vOdirv5FB4g9oZqgV1dcHm/7UBfAYM/N
8Dcbwa3dz7gQwnEXaV5t8qkh7PqhQk+j7x7Q0rW73G6R4TdMKTC7evEr3CsEasLS
TRAQ53MqKVHNCyz70TAh8m4jYXnBBxyJfgJPfkQxHBn7jbk9y9pGg/6pQH7ciEdL
H7Nnzg3gLPWnbxrhY6EKo1H+lKBvLdWjgg26eZZRg2QeX/rtxclKZFR7V28/as2F
0p0AAgfKu0NxmWFjcZs/2g/8/OSup3NF8KNcvLAOC5EXZG9QcLDtxYSL5I+sh29d
ozzTe+n7M2eRjuzDLvMtcA0DgAFitS3mlWmJKLWtTxPwiBiLGRbrDTezoLu+rqy/
fz8ikgIV6e3hRwiQtkwsKnKp4AMibbDhKqp8e/rg0RvMw31xNLsAISq9j2o6Tu4Q
/kUiTIxWG2Mgt/05k6mPFC5DSFgNVMM73k3znuxhmA/hL6wD2oEQYXusFLvEuY5D
J898VzHlIv+yOe9ht9lJ9o6o6IuzAHZnPLMu3xtuzFBsXqk2udYQ6Q4i2fDVjQEG
Zyn8SMCE+L57eBAZTZN+Uf7u7WouKSIfjKYZ5KqyRAy9i9Mb52NzYfs1qNZWDjLW
2qVWRwRAEnliETMlFUAznV4LZ0/lV0H7owGeGsp3rHM3tLxfQY4VYwb2f/megdo/
YrVfffqINmF1eW9YuvIfDj9OC76Uojg+wdvMOSUaDPoXZz/5B4Z61I0k/+1hea21
Li3xSIc6fNchwM1i+DGOkT3fgA+D8OyF2PSZ9lcaLsZoTfsHNQ92pxDEXf5/E1KJ
0QQE7vxvH1V1xIKJUJlaX2Q6NkoURqMDRTNTWZEsTPaWYFP7ku8Mrxth0BAABs0A
5j/p7NN/38xcX16PzNlZ0F9mj9PPB6eLZ/NnT5hqtwFetnN3Z+6wb9BR1FvrGaVq
t/x92tMMS75aZzUaHDhzQsMKHN3zC9Nx7u/2EZCzN5d1KNJPp+RP9gZz/a2XwVy4
+B+pybBg3JMWmfyWWyMg0p2C9AjAwj7mej4L3qjX/USzL3SxZIesluEKqpjCyj05
4StGFFKfYxE8+0VCaHeZyj3/Je+or21P5rkUjpmPmBGIW5xtUQW4F3oBBksNMjVk
Zc51LyaIoIqHEWJ5VedVvQPwNte49e2O5D75Mve/uWsjarIpVEZDh3WC4XECblxE
vpDfRjFWlwp1BTBhDVBBoD+tVIQDXzK2HX9wmfrF5ueMi1dMepBaXfPUz2+/HjM5
C8x5snypcaX1Ah2G7kivQ7B5eT08YjA4UnmY4kMD0EpeZyvtAOUGiMzykc6qbEio
JAyJfH2Rt8I0vm5AwodFJ4HwAE0zA+ZFpEG4mypt2ZO0keXw6f/jzy5kSEIbCNRp
91hhfO7Iwr2GyTZXeY2/KTbdml7FAfEHyYCyWZQdlvA+BN7fbTLqkoYwNaRpaCY6
g0MO9/t7Wr+cuSQAKR8o0/Ta88A7DjGT0RX+y1RMe1ys+/LsZFwabgDr3V8D9EOf
FS/rMmHRIC3saIedxIcVq3hw8E3NgzW8cmDsjvmmHGos1Kfwxgqh10IRhXPNksfz
GutjC2AC+k0FZHF6WVvMdndeWuid6vt/ab4g8ZhurbeoxrqyRnb3qxcDXnxrbyoG
hVYYYASxCamd+F3KMXPPDiLi6zGR+TfXc3/Q1WjvB8m3AFKYKxQKiKqf8xsgY4t8
so7RLB6T1OWmhskiZzPy8XzRKyPXLS60a9CHUvSYoyDOjJt5LrPcDrYm/3a8N4bV
nwVXIOC9Am/hOafBMmAQobojfekwXZXvJ7MYayYcuHxXWn/Z6I9QVTP4W0o0rNL4
IRp1fr1hl0GAJP7OSu4wdMJ/Eq5tF8kvddNvREiGue5UyOU7STjzD5851GS8ideR
CJldn6lUi78aYukySVt/EGVv8WeiyWn/wTOyA4XKmZO3pXkW8cRzp01AjYAN5NfE
TvNArAn/ZyFnnb/+26I8Sddl/GvGUAjCrMDGkBUAYjQCa3xUiWRtVWxIIIO3zHqV
QZ4HQv5+oY7C9Zot5cFU/MKWMfKPZUxsl/BdMcmf1xb8+2jfYamPjmzwECGhkwUz
0evchQfe+XQCPC6+89ryYNPF2wvpSam05mWYAdUGH1oWHyxmwKU6SAmXx9rru9My
yPKl8drEmkxERrM4xZE6nd3irZyA6ZeZ/h+IogMdNDr+0qmxP+XYMDKq3Tqehws6
mbz8W6Jhwd2iVnTZBJ+l4Q1Ql9Pp7HnzLK+xhUB1S4RwwI0G3QAJS64oZ6maGUlE
Cc3lUj//wdVFg/Esr8fJVowNXF+OLCavpYtm1tPq/X7vL5Jv+O6ZLV5dDA2+tdwJ
xb9Wb098RWE170ykyN4Qy+h7pl82w5PIqYUPn2rJb5peNmlGigYBCADIpV5CiKUk
7K0PuRvH21N4atIClMJT4zr4KctiMZm9S0DlEuLuayEysD0M2aR6R8EGBJEB7d55
SYFh3DyWDXnjPAmFxZS5E2yIcVAfx0QiqZh9dXU94Zjbpic4D64/YwzgfIuSFo8y
JymjL1LNwq2WBkvGifXrAmICqtJde7UlPihJYyjXFSWcf4QBnRtsOcprbwjO2mAZ
UAXmgwnb0u9uBWEWs0kLuryygvV3oGnJMmMwITioklTZRffJaM9OzaxMAPPxan65
piPg/8gGTKMtRGFpcRBV/56rKnFDwsWjNzQSTTdQtfKYnd0XglRBbmtrrVf5Punj
SqTiHSiC8F3xnTTd4dGXYJF5oBTelWCTVgKrs/v2JZDU3I0lO5fMgdE2/LRnwGU7
9Shc3lwsm7IhJsZrhqptNGCi186KvfVdJGvfO0ENu8VU4iGdxyXgzi3NdqT8OhNj
teiMIHQJT5h0vdRbRAfouMolhpuH7LyNpxumVGbBqdUoBG8K5+icHBEfqKqPfgke
SuG/AXbKjAtymTLjqYfyzems6G2qsMfMygU/jOieLSwDihw02Re7zBGZUCD5ONRn
rDVdvnhNLGKUvbeghn50gyOztrP9qqsN20o+bvRCK88x3svbAuphSGPMR7c/tGmQ
U0sM7Xu3JN3jNo60z4dzoJmOoF3ZV59BVlqthpbph8rr6+c66nOHyFd9ikD0KVqV
EqVqPHneddYVJT4UgjkJ6838G5RTtmkHDbwMV2feT1FguZO0vmrbVV6Ckai98ZMW
cxN/6FpUQrA61nI6nqC0d+yu2qE9KMD+INf1i8qOzDoGIp8WfAkQorbNPR6URQlb
ok9KI8T9AZbZNiUXmT1WWsBVciZ6Gd1g9GAt8k6HUSaJet+gVY2pNUilyr9xUpeM
FuSuqOL96C+RnLP6vuyxyH0TFOoyoJYDHP2Zq1+5gynA4cCF2IP/CHreJcYxzjzD
+jWcY7StGO+ZSdmG7x0vSgERizN4itGeiVHUtFtlQ3YEbys79j4zyHaiu64e2/1i
eFr+VqQvZZHiiqcuvQbDComUdp0IejFPm9Xh34Jx2W14d/G89mn9cbxB59rBRlKn
j72AGi3JBHEsZ9Ept0vfUv6fo/zs2uil6DoQFshBEKDfgOIg/qe/v/wrcF9ZL80B
S4HQq4TTexD5JRZhyUJP9s+3dZD6nmSsKKssm14XuHu195zPW1f8YI/yS/Rqh4/f
sahBZ+hbej4XgKm4cJXPj/YMaYwrKFqCry2Zrcdnlu8okuQVY8t3rvggzbTwTdV5
BWbj1p+EwtbtKBgL4woPSKp2PXzqtDTW0+LyzLaZZOOJAxFetu/XP8ohYZ2OJSFA
brYraodXAIenp8BP8ibXs4mj4A9siovQx3WAKd7U8A9/PKpNz73sC4ZNMtozYkRP
A7d5TvoGofDLYuLyInNTWLF4lZAHH44laC7IxIDCyx8nrRQgFB2gG0s8MjrgiPKN
hL/YJKzC+0JUHO0/qPTn4lV9cbnGpqt6xAQrqv1QnEcNFe1EbX5AhksxlB8s3seM
+KN0dL4NgOFWoU+CDNOGNPDurUP7jn/pSUKujEDTZq782XH1tVY00V5dn5pS9Q5v
mob6HBREDkG0ZcpykGBhW2/snI0ln9RMuleTpTwjWTFfCg00Tjm6zGIBweosSNnV
MiKWgxTegHF8sUjFdwXb2KcomV+jW/nEJUzmu1udB41d0DZL325qCAS3WTHuk2jf
ZbbO/BA2eyK1eWsIzCbJk0iNRhNx0AbgUXIq1Vw49gLY7Kc/PU7dsSJIAxlSborQ
YnV+s92+FtYCCrwJ9DWL92VZMlAORuiyQIJXJZ5TDqc04DIvcLF1oXcWlbxk0jx6
9qWRlTw8wNe4BlXGNfvLzST+aTeiU3lU8x2byroCYCHoMtQ3E50vZR7QKNJBIqG5
AWqgWAX+kpGbQ5jARs3S3IlVenH+J7rc857LDRBQ2VKFECrm+lK52CEl8yXoQ5ib
njN/IzsWKlxAzpQMvdez7EnnMMh2307IOx3nOMvlUf/3AN6ODMKIB++AB/nsJaGd
Hpd5vjL8CwgsIORecTplYqlh3QbGR2IVzaW/Rt/IQT0b0SdczUIgBp+p9H4A5G4o
gSAD4h+k3JtApmWgG78W7FUJnaut6uPtnHLNJSwgU17yTojqzf27VNrbwcXwNz+l
nhdJJTSAoX8ZEZSxMKlzVWxXpIJXuEyTdW/Ltp9qPslO7jU4mpuv+M/N5eFMGkyu
Okpada/ZapxZ+sc9KiHwUAwA8zuo8IJy1hxuGrMoyY/f9ofO2lsFNqrivIcTOqv/
OtwHUSLMlVGYPOylx2DSFF68v37a/LISZ08N4utdd5uOMmS+cLTpGikl1/DTGDya
r/0bO15qjJNyFl1pY3HUBJGLadmrOrBg0+JrKml7LvX1D7xoLgiS4CQFdTgH4zIi
/V+RJHmzYKiv5mfaYG3UFM4jKHA8voZdgRBLuQTdPR6xXJzdRtz7LB4nUfDXEj7s
aUodlV+XtbUcJM+KGx85HitWnHT91zl9adljJdO0NZ7yIkvqu0Lc26nrt5fuVRGB
E+ousFUqtC60Y/+ZmPHi7FkGEZ+avsnJJDSVj84oUvBMeTKFuSjVZYeoPWBlFq3r
NUiJ5m0P+Cv6TYi+JuXz53ByyHXzqO0B6825OUBeVTbeDrts+GbJ17dC73DOB+cy
RQoQEeG88tuVuYdNsVpm6SsxOWz94kGfGdbrHZ0Fbvy5Q41kqcI0YLi5uMxlYfj3
vOFOYbOp76B8+i4tf2ycQK7mOTx+WbeJEB+VH66OhYn3tLJjtTw9ckOh/fDt/hv8
Cj4Y7KqWRKhRRXjIeYJI4/dh7ZxsjqHX1+AE4JkPoxApb4hIpxrTqU/MRC8k4VVT
o0QhXXfVpA6pgHy6N/H5Njbo57ww9QAKG3b8mSV+kQhSUhway1tIqCIccnuvLV/I
qCePq7ZUhpde/nO/zJP1tyn9uHtQeietNZrnJ6IChKZPFeD+DB//6Mazvdp/49EZ
UDillMZzqpNnFLDOf4bUFtKUImiHYBL8Boi/gaq1bff7LDOrJz2hC2bfyUq1Pvbt
XAl4xhKdikVecFRGnaUBK7PBDO1tLxzzEH4lzPuaPAUOEfzu1oSOfi+znqGzW+wz
PPC0PD+wsxDy4jJ+h9ipAMu3VglhlP9fN/hi5pDa/U0CzH0wHQOkxc/3jNltmBQx
g1UEsyXqYnDf+ptJCz34JWcsesjKmsQLuG2t64DorjJawmMFV5omQT4WwxMmtzPn
SPKmNRr9vnNf2QYNDkaPDE63wBXNReGPxzx8toxdKbCPFDjAv8MQF6L5q6eHrfz4
vq7Utl3PAJy14ku1rEgAfywquKgAYJFPMPKIgEq5cffuv2ICvp0l92vv5cVgLLre
IA4eXZVaWjGvb+11IySApaTX+hv/Te8zMiEeNrpRcdJxefrxq/mlB+v1if1DA9xo
6TqmeyhLxVbOUPQWsUI/tFoxGPhp/RNyPQyrjI07iqQF5g3swQXMroxkwu38JjeJ
sCB963R0GU9Pj6lVaGl5/ZJTQZ8uY+lOjfIr1bFAsUIHUqLPpxRkwHy8vKcp7yW1
wcwUBcHA5Q6Hio9jFnmxZ6b9LtqZBi1VbLU1vWXfPWu+Em9znITkF2ht0xsSsohm
ikt4Ef6e//gBNMAfcSkEm+dC7HyJbpc9RffZ8XfajlgDdtuhjSBI6bX9wiiY/5gA
7qBtKYiEfB68HsZcgcwtm/jth22NZ7bdsfCxPGX2Tm5/Bzv+onsL8x2ulI8GGAst
YkjhYnIwgdf04X6S0LmOt8zBlLosmUp2WSyjGbRr/Mn53wy+yJJSCMJ72oZul0xo
PIyOXXvh2zt+OZhrtlPVoYnTXVDuV9G9HON0AQadUEUuxEwgho2Kg1QJEtMNaESF
PMeX7pEgv4qInO3lNn4x3h3ys03YENrvU2WSbPcKvlM8zxh3q6XeGWISXdeUIRE0
sFdPYizKni5plJDsU9nCIKNnIwrw6lGpZQH3oodocG4LL3xsaJbPYCQYsfuSVM24
gIufKHgtqg3FLk65pUSAaYzQbd0GdKLLn0X6/ngMsVSDWUFTTXVsBXsUmp/T/XVK
UR5yNsnf5cR8YTAc2JuGkSxvMZGBYJAN0+Kv6Z1SwWOeXEgXdwlb/rahcf5yPmLk
JQXCN2dGQtKhx3AmhpQ1s/OMtSYSNQyK3MXdK9deqdPfhROOp//CnbvJo4Nxkpev
4XWfclyEJDbxk9oxE5U5y4kEqU07D0rLtaTIlwOB+WldqMaY1cEaB6gwhvDdg/ZS
UJy6fiaVQ+GZTTKvJMB2IA/V5cD1f0pRZ9xkcVtu5R0BdzTB60R5VMaC2RrpmAvw
j6VIezChlFzeRBxe8lZkIb54LWNUl3hz9i+BEoUoRurUmOQWZlzU1bFyCu2/Qijy
Qay9gC0nqFyPhZ3+XK6zaDwmGO3zXnil6fGleJMigMpzN/M5zRIHCq8gjZfzii+k
VivCSa2RD39Jg+xZTDlgIZmLAlWm4/6TRz4f3hRDyTvh2Tf/BTeAdSDHLc3KyW1X
VU8h0QWZ6X1+Gy0nockJ4Qzq7KYq3Dm1fjQjiNOaDTOFkpKJWRVnV6+VUk1zynd+
kw+yUgPeXlcTwZCOfsDJUT7iBGckqogbHj8hU+2ySq4epx0KEC3I1i2vGvdMyc5l
cSdpjHZWbHQOXDO2GNOzIAus4hk2bPA4KYjmZvZVmeoU56qg54+VxWOshB9rTktL
tIrfLcH53yo/afyPjO5e8H8NbDGitoOmkO8z1zF7Mrrlt8G5Jmvd/AJ5kjX1tblX
wwYCK5aYQYJln0HyDw/YGr/kdehayzGbjH/vXFxcrphDzKCghBA4IRXa3Zo6nlOp
1OGzLPkO7Zj7FOrOH9p1VNghaAGATZ+zlw/XG7/yimIwfZ639sJVQbErjXuqL4qW
uamMnV/NsbuxUYaKj7guXxpdVmzCP+uh9poQnwNwzfMGSgtVf2RYBmc3KZXAqPHf
BZAv/G29YKnqYbh8THtZQIUAquSMMwp7i8+GyL0JaM9Z/UNN6/heu/sp6gVCs9A1
l2U5VcpiFiuDob1TGuaaQOPBTA7LTeRyQ/wkffSDnkDnrtOFPW818CPhPSXMja+Q
I/GOJD/9Ag4r2A0sLNvoFGFbk9o5vWrQLkJuGsNi1ySHncbosN6dFxx+b4wLHjvf
mbUI4DoHIo4HYpEKGpUn27A2YLQz5TEENW0YgNjcHe4Lyf5lVLFP9UX1iY0hPc4b
9LT0XOa4TBOQG7tfNp8F3nlq4ggGcnersqwC9Xba3dj7x5Z3MrDz174llSdntJ9T
4lfyw7GRk2MI0ELzcvfPcNFywITQU6GsQB/PigntRkJZEGYxYU3/zhxWQZR88Jy3
UzK5D3wpC5nwkrimSabXrpzrpEGHjKmdODNYK0YYwzd2nx9X+GUsDZLk+UhbiE4/
tUc/rHxQsfu09gkWnkJDwBU3fmD0fYCCPuOM6XdR24UXOF/XEnMwQ03qQjADFUqm
RvPD1Qmt5+stV/TCf4yrdu550caloSWhxE/3WWZGW3iYLSxBmORj6uF3I3UxVyDg
MWUJC4albyHRs7PBK2KcrE5IU9bdHekJsQGeCHNV+XSzX1SXSsahV1U4mAjMQlvK
fm5OrN4oSXyrb3Lw5cgqMiZHpuUsSzugSKRb+yeQvktDxy9AqrdLOryO0ungFIKj
W4aVdb6yyI2uWqLXq2Tk2eCcdsi+XgtEZ9S0+mJJtFIVHXfiH35DG7n1NnnIFcIH
rolMc5jlPdE+hdxqA6arOvru+p0A83nU+6zFY6cC3TWkE1Z09NvJgKcXhpmR59zT
35pV+XmdPThiAx9rg62I6KoQagCrNv6bdPqPqrMOr0MgkBy6B9w7xOpU6F8O9PHC
abag5DnZ8GqtkqODqAkF4cqPMKaWc6FGpQOMKe0d6nIWwBi/z5VK1G3FkTvJslvR
jKnFkgdqtbPvSznhnX71jXaNxZazxYTEcwNQGc3tflrwIpZNbtOKorVnjaywgmPK
0/71XSyiSezW8HjXNF0qdVHOgSNvBD8JjzXB+MQBYunjHnzO8C5iWvmdC+gbKkgl
HOT9nwCArHY6PtmknSnnKDvlUTXmiKJsyClcPirOKyHS+rOSK/4PJ6zs7zHcVYsO
HgTEdFKlYbU6N5LcZ4jARV8hUrRJmogqF4LqiyblE0CXwf8NBc+yLUcgboIDh8r5
xccEMNmHyayVEncl/qE5w5wTAMlJSUpeQ9JgVqbtKgMCrPpuPbhdSt5ZZSU/UlSm
gYaDJby+CiaYA4WNda3iiVkWi1OgXyO4QeJEV5cPEHKqLkAwTy9fZBn42ZZWNVLl
/lLapWFn1O8h421Mss+rAzGoV9tMFBY3VlaSfAwWnqA75unn4dI5pshE3fbQUxxH
nVcOaAbW/SWRGtBpw5PTRjatEeZmDhpV5dQ0KyfHl/B6ghTvj930BGYizxPJm9G8
u2iNG2UmyzB8K1TERCK/TeMPmwoMJde6mzkIzIcrGJBYyUcVEn5Kw+i7hUBag+br
wYsWFI08oGSntmrU1+PkDZZc/+Mzh77zpN4ZLzrnwdyJfgeiteGVWtncT56OG+gl
ye6zxTtYmMMgDIg/JsE43YDW4wg85iIqWgYRvGvWxhJP6uPDMjPGOXC/6Ixf1gCL
kYG/5q1L31Jge7rgiXksBbqUx2p4hcutvwkwEdH4xlqhEMkou2U3lRwWQkMVj/Yp
PAzYnSO5hv9U77Y50ZU+5voMR6bTGmzQNv4+wQuBVxWzjbJTK4QgI0BZZP07kJQ7
VXmtINqeDvhLdE4oi6pkgeOvZvjWEUvrtw6BFSbTEFqDiZX4ECoJ6zPhNWX3113X
8G6kTmkcICaktnoGKD9zSqMVGWsWySdmlgoGliuiXjDH/xr1bs2S4LdZ53GXi3BU
TDOUGjV9pH+aG88QIZ+5nrbEGKIGortLfxj2ljwQcJMuHXXRLq8N62asu3dJd0V1
Np4ycC3wpX91ItqsQlKof16Q5u7Ft3zcwvdY6L7JCBB8zLkgd30u6Rxj23xXbHDt
eAod83jBZT1V4d7ILp0KfznFBGp0DlYb4VPYCzrmCJvXTNoreDbeeOD2hoZS0eVH
y0mGRk/xSPBkgkhhYRUSpmjOiZx/hz5uk7D12gFPeDMSpteY5sSVt34mJum2ijCU
SwE2X4l5WPFGpq52Z2iUPBV7o+TRDg5G//oSNDTuk3ygHWwrA1dZTmiweIFytYHO
68g4BwATS2rc6BIMKpmyJxPvqMrntRDdXRzYg/Z+yxz7zHEEQmS/f6QiyYVv2QiQ
YM2qlT89K2C8vDC1blLQe8lnYDoj1nr4RDIA5W8imKoDOfxU3EK7kchDnzQknK/I
tAunYGFqdYtOhh1NDMDcxjPr74jqqc38/gCxasofIf2WjEd8fE5OXJ3fzMBBIAHm
fTuHwLsQ01CZewFHsyg+iZrafqQ86z+r28o/4Ncj6XDitxkiVZ+RZw9D9meO8xGr
GMVNIapIx5sgxoHxAdMQYBZDxEURYXB0fh3ya9WeKGP0/bw0iXGJbdZShNLGsZb5
2INQTEHM7PnnqYBVvQBjXFgKJv4o8jNe5UDFhv9SultRMuE550srtLs8TzvlEccV
exm9u/kgufpkR6OnoAfOoT9gi5BK93XZciw3q9OytOGFN1mNESl39xa/0YKe3i0U
rjdFV4C8mxhc08kmD5FzNiGYbROX/k+VRGWFgPzqy8s4ASQu4ccuJH757XhFc2kc
MrwfWCzDIVeMZoI+IS6Z/8B7xyO2SFEQqlhtPrwCZspxPiNfd+Z2pczLtgZxRJKh
V7hKMYb6SoY8bGYMt1WCiMre8LooOFtKXF1MIQ2gbxMnRo2hPG17U8rss0GM833Y
JNJNy1h2ZI6339b//0nl8gVDdzr8MVowXPYrdSkodpWGeyOcItZgLBEjYoay4qnb
IyviSLuQSp33C8AfaXk52suMFTOf/bCctb24qNrqbtKPte8QJxCZJ7SGZe9Lvh5a
53HkSP6OiQLLyOuaVPbsCD9Nf6Zlt7aXg58L3QMJjmpWe4/H2Hf3OgbR1f+GR912
Nt85krGds4RXlBu8aQNfaFNcDQiautpjGvEUEKw5AE9y35XDz5JomlTzWbaF1eZd
1F6EwimHYIWjh7FI4x2VTQN+xgYZAM5WziiUYSC3jMZhk0L+OX7dL+X0Ws1S4YtQ
ise7Plspii/bn78cVJHRN6YnXBYbt3K3CIZ7Ic3meS9EHxVFbcNjDkD+MOeDFk1O
efHLvhVDMOAx9x85PCpW9keG1iM80t82ukUOckL7wl8Bfxq61XW/Xx7yJLmuKIWw
LoKcT0jpMlx+KaHrUC2IcX1ye5se++8y7+HBu4z4eER09luVNksvMOTBwXJrM6vu
sfve9Cl4o4Ve8eft3162sI91GNiOtiFyat9TqeVvmBdxdN9zHK+vjBk7xXFIH9c+
1dWMt5NeF3iCZn9yPGTBI1m3WBk/2jYuCCB50JWY6KFPinOqANnrJybLv6YSL4T2
gB2aKYp2mT/YK0QuuESeKw6I46j5smv/HNtVZ7pMA5g3iMkkxLG24bBYK2FT3uiQ
CTtIwD9RuqCPilv1T6M1ZEHmucsqKvEiVk3EF4AiiGZm7y3HQHu4rp2RIGsu6BD0
hApuVu52A5nzuqPoaExLqfqBPI0EYiLWXQ2wTWN6zg6XFFh/N0f8uYij+HWW/GYO
7vgA7wIG1B5M4JI/Bk3zm8xKl6bQqdYktveO5/Ws8QoG6yzY1P/tpwxnKKKdmdiR
ITVyVO+ukxAxXmTHYmf08ZyNZdzn4Aw6Nm7KUBBJBDpm2s4HG2B6JYDyaJvQwAmo
uUTzq7H5t2szVPI/4j66vx53FcciUpIbd2CV0d3u5N3veqxAmW+a5UfKj9lnmA9B
H4I4t2d0ZIWRhMjl9m57vLKiKmbJEXuNOycndw4QhJ2A9YmETikXjtLMC85odIi8
2iuiOvN3cHSUy7oaVwTS9e1rsYWPbjunus1kluWQM0ES9BpFOuYofMOQx08PLjdu
BulI9iAEiSw0cU5Csfb5p/1gOj+6rU6T0/D0RuZMumlAMfeV8InkLcH7D1WLh/SK
hueWwlfQTcunoUCnut5deqWqu5HUOanUi953z1/2OsalTSNMUoB1BDhXEdv00o39
M8+rjQueC3rrVv8pelWLY37isE/8lfa5BbC3VwWKAV5lA1o4DyxNdaaV653hr93z
gZXV5xw4Dj8zFc+TTOldAab08gBHiJNeb33g8a8VFavaDmOfZWiOPz7dHPg8clRV
gKgjImvrJxXPPmhYa6i85+1cjTcpnBJn7U1rbKKWZGdVr2H9KluCTAGr1ZPRMAyc
O1haPKN/TdXvbaiIwmejL2Nfy2VshZvzu3MuyF4XjSKWOKPpkA3Ii1HmLk+eJfDH
3OGa3cIhXY80y//DNZlifz7FdySfqTaJG9hjU8ofS38TtzKXMRUrkaCwBFAmXHpD
4zYnKlhb3VB25b/5p3VewpQGH8CZnzSTXfJznAB0Ca4Y5ljsraBFu025nnMSYFZs
KL30ovuEidtbedfCY7OA/V5FTZPAMMtcjiIxvhBAvS3XWgvc/3GAe0EOtFcdauMp
ykLidCg7FBMAppxOuMwrLlYghAX5RyhropnipLY+K9RS0/57JKNF6e8Lznoj/JTR
oKVkZcIVOpSpwlHz1lLUbqyZ6UudkwmD2ZfdoiEYLHDN/ukQTfswhJvYpRDEF6xf
6PZ8R/HxCqO0yvAhZYjfyPTF6PhdE8NMD1TpxCXP+Orq4ZvLdHM3cdPG4RuR4E2J
NXFydRZjF9njtFzsh20CKAA5qL4lX7FZO6YoPon6Y7FMhZaNMtnoEHPIla6ax5Ik
tCLx4s7SdWYAthlSRW+ZZOdUgGCP9W16fH+qB4rXwSqODhx3BUel82kp2FmKNTtd
uttInZM0FToumWKUqLVZxbFqRvH4qO3+2diHRrIy2Q6exgEFNpeva9cD2ze1K0zU
xnLgK4ahO9Ekyn3McOoH/EVnvvv0vSfPaysn5PulsZTL9UCxQHnFT8K6wCjRbs+y
HtRxEiz94zsjFgdLh4gtTVtoeGbkZQ8Iv1WTe7+jKZYRb92qDU8OFjPmxY25g3Ay
4LLnBq3V+RUPGVMMfGbmNeQDQTa2U40mjirQgOGBNzFoFD7WWVXygHNxd64tCuqK
rMgOhLOtLUlbpefuGnmZBRzK8499R/1+LWFY9t55dcmncPTLPiQcB7EBAToknwkd
53xTGfIaNEEyCLDu8/o3ipxkvT9uIj5TWWaYJEZi9PnWzdao8iFC+X0+54quX/LZ
fsJOHyp5frW3mYJzgOEiMmBVMfkC2YPTzOeF0mmVvv+Tg1gHTIVq0Cgha3t1xRmG
Y1XoOxF48C8zVWJBhuZNYBn6lG5p/0AYA2EUvN//4iaNSrOMVbV+6eW8yeZIKGIE
2lCw8A+J8csjez3yt3Pjc9NBAlHJ145LBCwucZzvyEnLjE5hGSOlCsmHR5AOmP0z
UAf1n32WfMMU28hRIXfxRk4dpgRKyg8TjGhirEelvpd8HBHYtAUIeEk7l2/RjUsp
51/76yfIuRi0C/XwtxJ0hPP18UlMDM5kkAaWxsWs/3mPAUm2dNmPlvxwzW8y382D
EM4GuudBsvz7hSgF29TVzruIuFKuUV47qgxS533qLXRvEANfwH5YwJD+VOctT0EU
V/Z1VpkqBNZS9E9CYdGmASsVr1wd+4DNL6CeCsaR1oVMMOJf3WWfrqk+fhV7KutM
/+C9Yrj16pAaReRijYb1PBHz0A+IfHIuVWDbMluk1u2oUzjPd2OvKYcqimcMwXyf
JySFX6vkH5A0u+XbIaXRsW82xmUUz0QxnsqRZzaK3EZYyE/BtBWKkwDZPe1puurT
GSkt54BYoXapMrkV2OCLcr+LUJi6OmrHamNol0EP0xB3gXT5F4ND4kkbE2t0tkTW
W1GlPnpq25S/dnTL26bnxv6kEwZ24NUh8g+3lOETOXu8r968K6PezpWjibLiBWv/
tHsVp3mcQmRQyhFYMDozMBy4vX2UP6Q2DcfQRhG8RNU/ppXJWCskZBPbLGLw7zKj
/qqH9os/bjwfAOBpduAR+hmkmFZGTc6R4k5kX7dEEzE9EGpea2MJG3yFzHWzNg90
ba6LMl3yBZqF6TmHC3V67/RImz/PiOUweD7ZY/IcfSqo84moYW1A7Yqi5Buey3uR
E4d6Bko5vxEn9DwuzGDcZlZpuUpaVuKCoVrkiYGiWvlvQ9W7r/HSnY7L2YXsvigT
Q/5q5CYNMjMwliXnBgVvKReMCvSPCvTB0nzvD2t1MrNULowvyZadyfXv5NX4rqTG
XDdS3WPnZzwDln0bm018pOXjWYOOvAqn7D0dTcujjv82wpFpZlUdtE3IyChLh4Fp
QZjxVodnIKNs/l8ENcxIUmqjU9m+LwRQ+VeknSDz/gRwfJqpNXxlPAtekZQJJdPb
z1t/kOv7aMHCrvEJhgJu53rckNSJPZl2ePp3dSeHaG2X+NIiNlmYs+a/GlNqj1xi
ZBieGD5aHRl9bxCFgxj0O7vZ/J/44hCy1NdVJaqk8pyOxlqP+851NQi3STu+dYqX
QrecZ3flpHM8PzSuMnQg4+MeOwZtwbfNRhXb0T1yJskNhxDEKS0mq9uwhosCDbKb
3FUBehLT+qSDLblT1qYIMusqidITR+zBeqi1/CG5TllFgZuPV57r8gAW/hog+WM5
eTRjeirUYbTmEvELuVBSR1vcxa0asDpQ0MQiA5D5avpT6ybHBCp3DM5VhIsKPVFI
Isx9cayQ75vYEN2QQqSFUXdNE4uTu3y+9dHB4NlzTeDmHEWpjJFI18X4UyTnejeS
QDXw8TUY51xHUVbanJTLFTIVG5VJXfvRHg08L1v52Q9+VETGAcHd/IzNZmUwKvEl
mzRWEC8/3AaUfItZrlNFqScysbpVj64IBqEABfGDppiNX6JTPsZVG/r5KwljnddS
bWRgoWzfJzBo/6idrnXmdgXhnQQaYt3ekSwUBp+PN6r01BG7lzvsj1YZUoxLI2cv
T+C4Kwo8CqaRTjs8clRY56/Cx4k4nXQ0ziqUlFLHJLaIaDeus/TyinGdK78mkLPs
s4tLYsUxYiHWyLxqbPzjxstop4567U+eHNs5A5OICtN8Y9RDP3p7Gd6KGzeIDq0T
WRIV43eIwKPfg59MLUg8ITp0EMXkJvWSo9FsDku4e8Ut3TzCvst+NWEyJJAS4cg3
Z3doYYyzxKG7WLTph9JTYsIBTUxj1pLE8AgCeVyVttTzfKj5vAlKvUyDMxxcAEzP
dDR9zQ4vhkAxn58kORVQqqq/c9mlIHpCnpPmb8in82JvpygZXM3ZoqZYxG5Zcb5k
ViqyJMsQKULAyDixVcVP2K3ctymiEVjwzOozfNAqAG37SllkwkWUJgmEYTvF2xKU
hZuuYwXpu9FmeuEPxYj8Y2aGJ/xkImIf97mVjtHrQ6wgFD34vg7O48lP53CGuARQ
C4NyTMNQEHcqKSPLk4aRPfrVF0Nrez35ItGxq3nAEHwezPqd6GgxL2UQyretwbp/
8/A4tZ6w+xjXOXC19YyIurOlGJf6T7KcBE2Ouv1jtBTzVaIJ7lLgyQmESZVi0yM7
KtVOXUXIYJr7AVNEPC6AWvXI79ljldyU78VldI3xCvZtgyfypk3/r6L4mxIzRKJk
gghFViLDfO+DezZVaG7aPp5ebNpbX41A6gvceqfzZH+IprMZmdqUHlvnX/4uF9aQ
qNxORZRsf3B4eaLC7guki2eemD+DPpRmeixkX6bI+XwXWPLaBi2Loh6tMJg8gKjp
ntC6q3K3IqS9SX5AT2mPwDV/lK1RAiBFGQofccZgWZfKZNG5h+XuEmB+/qpdJFLu
q6Vg1yb6YsvO9LObN2eIPRqVuzusZWpa9heRkvbSn2Rn4V3duc78vhLnlCIy5wFb
nAex3PK7LvQRAQtP2cJ+WdD2sy/yraWl3CMJgPiBcxHFoN364mwbAe4HX18lAuGd
mRyiUGw4aYCTuAGK6eY9SbN9FXKg7ZxFMMxT9iZSUX6JFruKGIdpW21qL4G31xXh
S08dsBOewK5bcmPMZOC6QqskhcnGXbEYxLxKnHwAkk3lh1wOEP4AtneZ0QNyA/01
a4fIxhlDL5tPRY3QnZv/drNM+UqltMyZAKS8ejb619CTrFmlKLhrQLP4GWKbZ6zb
vlPA0+Wbt16iDDu192hGtkCFzSSlV+Kza0BY7VDPqU0+mm/BQ+ms+YXQJ5QSzlGt
AThvwCP6b7hAMK9AXRLLiBA8m8TSwbxXvwSpfTowHe2euQTib30r+oQpc52VUrAm
YmoqTK9+fYbikuPtae406T+OcOXs2UurCyj9UQXfARqekLXIq3bt6YZf3RmW3leS
iMPeVhmYI3QtCpmS7vemS3gWnQ+ftkZiYMnGhNZ2BPygfZX/UvjX/q/gfbKnBNWi
OkLP81uA9DOTDhEXzhKiCSuGEznT51aD/VCE1hlqcKUB/ObMYJ23reAqZ8nF7D1r
XXJgd3s8/ajpvikdPAXvs7iXm3maYw/3XUfmQofb17aOvPR1Em8ZeI1G6bq4taKe
j8NPbdeQ2NyQzv6T+oERN6CpKmGl3YEZGTbvLVjld7Nx4wPWOKp5ZqFgEihbXzYJ
7qOUp9/T0jh0hoWby3+ooBnR4/pfjX6GhejZbkTcC0YexStaGY/pvKJ+wMFaJs/t
zmIT6JF4KjKfRwLASVf/CiexY7XvBjBnTuFja+yhhgx1oGSCCQ1oko9BNJwvluXG
uXSAFruFcd/f3arqRU2MLxzwg8UVRaIJnQsPldQh0aMfwdeYgsXQZYjt1t7LbVRV
8Y8ZhL+Lq4ATL1dd4hCFvgRS+4SYwWt4NPtFXgsqnBBSobDDcpUmvdAZyQR55UJk
jFGAy1C6OCqGAdS1d9dxQYI73SX8eLsTLR2yjD2aH8CiX2CoV851ZgxGofvsvoEA
lv9/dTMVDVj/5iTcoJMnM3ztKWPJgewBtb/ioSuj9r6GCb/IPm3t8RAhluYJdyRV
/Er06mYa+poy1Wk6VWb5J/dDxMeZ0eukFLk/NYzFXeqiqrdHcNovP34ofB4L9y0K
vc41Pn28LswM0yF9m2WxN4QK9BCKM6Sa7B51zEe/wr4HQbmcUUUeTCefZ5nlkxVH
X1SeIDLfHrFsW7mYCiuFRbBlki7KgB1EuOfzzuW4ibuFzvXPptMigAwVlrYJN8S1
5hzYrBM0onqLrYNHiZ+aKflEwp89wqugdOx0eGOcXpKVAucY8kNMFz/vKxCS194n
OyZQZj8OXNYadgZuBRGF2qy/CQ0HQCPIszmgOtnh7phOu2ykMQoQNhposKVO4+dY
V2+IBrbz2oRxMfxqJ9nX9Z5gUtcOCgtdAoT3Yf9LV0TlQg+ns7Aep6i4x6vP3/5y
Zkvx5kgaKFtNQyottaGH6qjDttQ1uD5oMYXm4olRgUwN0V2yvJrekELIelfprzrR
kRnrs/Cdkoiub4d3oYgD1BaK5lKc4LI7eAcmUCNxiMQQQ0AiuWKQEzlB8G1RHJ0w
L52y5bL9NPMYwJXeLaev9iJAtUA5j0dYEp6w8n+IzJy9sWnpAu1uQXIbIYmkfNdH
TQ7MyoyRR37jkkgA0341F5X8qBW5B/BouZcbzMJe1NIomirMvF21SQ8DBe+79N0q
RZNqloH9v3F98G24LAhVrkxDiL10pYPRApyLsfhrjPdwu1Hb+jwMhfnmPWu7GfOr
djDrim1lCyMWnE9+OLyEA7YWRZrK89ZZUhCCEsH7HAoQi+bBOf8uwAi4Cl8RFs6d
wWrr7cz9mlsK6c+His7qUNBENEll2miXHwnan7RKFsQJZuzFtnK2o6DaMzFFjPbv
KPcj0uxHuaZJRCjorYOMq8O20njJ+Y3o7N5pfveUADZMFfzu8mY/jvqpgEDch4F5
mVhOh3SwuRReY3NdCr5X4OzWwkLv+l1iHViapJVee1k8IzAyNLPkCSE3vKM6uXkE
izd7eHNTKT+EBuC6f7mOcxqQH0sT9YuCnVlvZuKZh/v+1rDhxZBG6HLC/6Y4bBN9
zO7bHTbq1c8gR5jPgMVCNMHHJylR/gkc7JkL6eRnFDSJNNoRgDjd3gplMPTu9ZCw
FnOTekzoyYNiTGB1o37ysOdPSPgpgxy0Ks2/mxEM4zWoGv/9c5HAwx11hMWcvWrZ
IJ1EO4z8Vd5m1bqRaCjnZdrYgQ2Yv7mqD0Lr/7wM2VGt2zYIbA5Txx0d8soRDUKd
mg3vEmcm4g/9dGO4WEjWTSzrx4nVS/MvYsH9zVvVjcIhBoKU2V1dCTMeVEfAfb/y
JjbxlJvyO5/j5pXJ1S/dEwqI4HzVTYAMd+MuDBY1qRiHR5vfHzLW5SWmQjBz31Ue
naWX6G45hhQLARrniKy32PmSbZDgB1ZQscDPWL5vMYnVRbPPaNzJQSgmWqs5QDAV
gFl+9M/OpvQFfIxqZelDGx5/JwOLr0HnL6AgF9D55IRisFYyoazpkqeWxsXuFEzR
TJ/qbeyTbpICs8OwZ2m2Ml8QJPifVLXbMlBiC67NZ7YDPvt2OJ1rLS0yeu+dkmkd
bflXV+60iGPng+Ia/Q8zgGcndkS26T5oEMi3MDOYHt21LNsovVE9I38gZgc0lIVj
F10kSi7dqGWkyqNc67AchZJUm74G8LxOExPnU7geLChQ6mES0uSY7pckrCwHy8Ed
pzcG52rVYlJ5O/7u+8LzBTj/AJQPjD+sao8RxZe5MEAGzXJvH1sbFHLmvzx9K4+G
lLeFCsB2ke+DgJwEvsnNnVCpSRzljlBmAWq7+uPvxB8V1GHqpZZOZ0v5/h9fbZX8
u3BAqQGnOVgEInMF5xDCc4E9DLTQiWGByu+A5jg6hVmB0SaLQOnYHYrPp/HMWb/U
73iMoSeEnlmVuJBKczhfTP4ZYn3kIpFWuCa4gs5q1Iq+DBSaM2TvXvIqV1WaCyo6
ys1BpPfeT4yo2ERJ6+fwsYKjkznv2XyQ7sDMcOGObzlgie7jKv8o/REiZ/9W0tSH
qP/WwGZCr8bPKQBDBXSr8l37/fpkaz9sJ9NrD0GGXYG+zQ7K90lHStWD+p9jdsPW
KDtcXAmwNBpic4rIZgQQYcQ3uhCJveQESzn166lvAns9bauhkrwvnfu/k8DTlsyq
2uwGGEq5ylSR0ix8Y0+q/pKUKWBjJ1BD3F5wMLtd7VTKmPywjifEXxz02E3SGUMS
LOS+5GvJTzG+lSJ9oJvRiaGVIYBXhIfxanUl2l9ZrrqOMyfSZ1TbRiteF0/3lqkq
vR8LK/9oLJgOB/W2P7m41XJ49XAuyPubKXL3wazAJNbNyCL4gneqHfDivAOFowct
yzDoEqXApbZ5xpCyCD6XoBIZU9nVH0jcruR93+kjFZDJhsvYySUPcSd+M6vT69yf
xhnFlsbquvLLNVweXJg/oANdCnN5NOYMCs+OKJo19GmZgpRs1LzkJzhsJSGtPOVr
/bUGvR4K5T6t1Z+vt4fnosw/bPiYmTFTe3W5oS0RKYDxCmZ4ECKO6L/ymKH4Bk7M
jMko6D04Y1MyMv8V/+hSnRQjFJD98//Mwzp0vvKBQfK5/2UHvD98bCMhPatNzev9
4XHdKFGubGE7QnMCT6AR/Zzgb+MHvOX1rCkoNWTHMID2nVTscdeOT4aj4ppGwsnD
hFof9yBziCc+UjiWEiN8QWEGE1+Ima/AqGLbZbsnzVY7oZ1ScKof5Gtr67QcF8Tz
QTzif4Dc7j+ksoEMQ3e1blTh8pv1xZ2bB43min7XGFAZhR8ydvK/Etq8frTzztP3
mgbL9E44hdfaAqBdbDI60ioViVSFaf7I66Fu9m6mEPlyacoPbiDmFbyWCUS91sXr
EArzbB+YTo2ZQVWsEb2oa/3p0Rqly4eeU/7o4U3m2uGT9CPWCxWRUvj1KQui8aZf
vhnf8fr/RbyTm8kOaKFZeRH29ELizMe6YfJyMEMi4ds8ZXwK7HvTQJXHVpRlm7wT
Vzyz2DneJpNQqt1wKmrCB8kth9C7rjynGdTLsuVa2OHNbBY6/GH3DjhcT6P6O+eO
o3pGQCSVLwIZDOXBm52UY3It8uYGoUup5TikrgVNMRi3KEDV2a6dlsVJDBoraQ4x
LqKcH4rVwgVAHZXB+GBH1w5vwaVhjz5RcfBTpg4CNwVCse6j/sDhs5OKnKPk0FEK
NXi154zewRzuGTz9u0GoU9nrFxvDwgS/vkQqPTzmEVxS3ePjBfZOfwoV/DrdFMmK
oBusfY6Mz6H7oQPQeskNn4GTgTZAKUEj5enwbesv8kUXXgEOHsK/eZa0Gbpc33PE
1T6hT3Em+u2MCPOupyzPqTqHYVAR4v0jQNnqQ5Q2e/jyuN4d4nl7YBCIbZQJKRKo
9RAfRVdohWObRVDFhxa3TfRI+KEzbQnmG+//1aixhT94c3tvc4fPt8qv0bmwHEHq
65RNa9B1mvK+7od7HHJbPRvbHyai53l2Hxwei2EiPT0RoPlROqBDpWdzOHKG0hBm
ok3ffkj5RHrcFmQ3sH7pCYkjz6o6aln0ED9Fh8V1eM2RHeYlirpbnVXvtqmeI579
w87bI40DJAkn0z29bBeLnIphyZqRNxT7AsiGygVJ+ooS7J0hheZhXcCXy/7+DfCP
HJhvqe82wbEkqckylg8wdSfFjHhm7GkX6XsuM2GJhdu1woJzgJF6mh9LQ9hKXyY6
aab7Shq1MSmQSyqauSNeUp+btWG/58E/S+XfNCrXa68wlVEC9eGFBOo38Z9D/Ca8
QeG3+53CeMJUL1QPBCwmEr1yvV96NigG3Uv6KaJYkttuVTD0HPcBGoctoPF2pa/b
zUna1jXpIJY3zsMwyvFLgoNGQsS/4JP0DDvtC29oyeKjINhwGmhd65RLXfZrzGSh
KwJVvfQWk7I9phd8i6Ez1hd71sEdyhC3lrmGQM7U8u1XumCTMzN5d72TQ/S5VwLr
SbzhNENOeoutbToNVzegUuRGGNwUkO7Jt6RLLnxzBOwg7xwvwXJ/N2NkzVUXb7zM
Gf6nWkSgkAm21BO+FUvgVQmIKF2nAb1baMNlQ5Ed0K0IyVeRXVB6w593GFai69SV
SyWgJfYfAzrMv5GtRbG3Fjyks9tpw3YSHsMN4zONyN/XhdpPeGVWzTa3UnwQfsYv
qjwKHHIT32UHoSGow1Bo1N+AVjNCXL/q32ef/1xtY7zEZ6JXHKYMLnFfSHYP1CCT
qEgQA6HjezUpjH3eZOMAdih/LMGbM0YCtJo6vmYHJ+G/Wv+aRIWk7wPSHyXcl7Mp
jBH6ICJFN/DUZFqgYVaxsWGcqtCPA9agSzZQiirp0zQaKkmMhPXhcuI5kYZsp/Rf
54NnoMGQkRr/tKlAgClGb10/jOEaBF+wVYLiCgrMLrweGuKsZOHm+rJWkUs8QOU6
SfbHmjZk7bp/IWbazpNni2Ua/BgneG9t44lC+a8X1ObGM17TJWuBqYTnVsYoRW/P
uc/bYru6Lvf+4sIwf0qZf5QhyYTCcpX2J3+eh/gxW3EcS2ALvQZRKQlnXVjoWgDK
uDaepmQR1HW0pj7beGHK5m2c5q/xi+UEg/kolfnAUTvBzQ+Gm45i5OdSDOjuT3dJ
NCboBKpo6D09XH2F82uwHdeKWN5eeFg/q/UpCseZoDQsJ+PmrgTNPZ94uKHqCw0j
BJAU47Tz/m/mYZAP5d8To9VpseHZ0FSnGBSHr39qdDCqE0fgsxV+H4lBGiK3HsJC
1Hy196sV9G0lJFB5kN9Zzs8rKaCC03WbyRrQmqo9Rc33YtULbUFtk4xHf/hKEHqm
hJF8WCDIInfIzt/geIOaf4US2hiUpXRZqjfjJlZ8sQ/n3ybdw6M7scfAeficORvW
pkIAwIsYrhmK1mk9EK6RmVX2Cnwrv/jAY00+paCsjOhsO2AEL+g8efgVEQGR+JlA
HN+u5Svj86SMHMnHcz5ijLpzVmwt8IZduvBNIbPfwiyEb5xXCTtOZFQ9S66G/Xqa
h+TmTlxAuyjq9bhkRcjTpwH5CSUshzB1khxZJxVihtvE6jBUWTs7n3/j8rKJ1+TZ
mhQM3WN2JbMRvK0JXu/3LhFNY+6IcRzVFzyyJfyD5Ac8JRTKKWMyqpiqXPdwzwQs
6y2pHI1tAeRMK7JxmKgw6tToNICvOvzxYWvgDYnK6f7hbsYsli+kc0oxhXRp4Ks4
hNC3gcl8HcwKl/ZlyW1Rz9uT4Dgvr+kuzrfEbARdL0ig2kGWUAyU2y6s07dp1NWI
20Ax8Ok7V7/Sa0hr0B7hT2f74yQxUpX4yR1SWMOA+9+i06poi7IE+yRPyB9d1zD4
bx8UEhhEZ48BF/x+aPqyCsXfBEHtQRax29iuk2WdcDRvQSlZNYlivTA0zkQlrwdN
arIq/Qr6XFAtxLY9S0cFvEea7cNK3RGuzsuJWNbuaNj+jtGpIYaNdy8upqw0obTr
3AojcnVZVtQIgHyloQxRjjPwnO65q/wOr9La6tHws77NWU5KVy/1Fe9mGGOZXXJJ
IeuY3Wk/JZrKjaosKwrknkOvxbbB00qfyVzulavgYESjy/a35C/PsiHOOlpYaKsU
9vj0a7nBNs6uz2HXgxdBL92/9r8w4tIYDsjk73jvTfuwcgvjiGjzCs3QNJ/fSwcZ
5Q3o7VtEhh/KJYGovHao+brIxWaRcGb6t21tERXxZ71yaPJZoPSDyXJa3ee1knz1
X6A2FuRVydb4Op++8R+Meq9lAbqMIgHfk/sHYcVIADoJ8qVo5O711ZkgM3nn/Ded
RaAGgAe0ARYEjFFwAMXG6IupI0kJu5XScsaL6iKKcf+cpSf6T3QLKwccXFefExkF
OZ0YWiLjwjimOHPK711WilBAKITVlyNdxvf2QKJ9lNLxJjyn2deyGU5T7oSOYpqF
OD3gSowLLU99VavNX5WWFgbvKu9KG6bZMEEDIyDyqtjl+oim6dQRAwvxXFcyCgFf
iyYpOeULgwgBsu0rd20OF/mIYcndv0AEPNwFK7ZykjS8EFexPNIk19iEw2HfTjtT
Q4ObMauGlPNeoy62lNw+i4Nrj31WJXuThXCJXZLRMWY7+Kbn8D/eRp/nO+Ml7wVr
txAgiSTAXZIJ9F7KYae4e5pq3WuLyRWSE8hSGhX+tqDHooCGJonhxSc9yuloZacb
P+vKB6DOOFRhMvbiRp5GR3iwKj3qmc3p+WGQZAzp6mZiZKYVscedg2nkuvye5Fyj
hsjLAGAFRgwVwAGZ94PyO/PZ46H4s/xhIJa+M7EcuUDKPKvien2YcPbc5SyVDw8j
sEYUU6VY4yui6+cYmWWe1bAnBfHKQGyQDQeXuY4jb72MPGKUyOgoX9oWre/h2/1v
1mZW9FC0/iWLWsuBLChZVkGmvlof5oYdKZq0LKjNtipvHckL3hM+oxbrbhrVsbpi
AjiNMm/G56LNkEN5ynjn8fG5ADgaOpSqZrhMVT4WsOWLjeV4OXiCR2L3mHIZKJxC
dfqxXDGf0dkWyDHMsMdKJIzXbJEf+yu4CkJsvSxlmkh+43Es5J3R/CluC+XoYoPL
VFotF9zwvmAj187mTeJAGSvAWt/YYfCiQSZF+oiWy7R3n4ohubDLaiFEEU2X1tBr
drfuhMd3YUsfhs376GvKwOvsAKiYC52GYA+StQY9jz4z1PfwE8x1+qCYqkvvn6HD
U58Bxmx7CAWbDD7SEEwxTu2pWr0JuVXJhuGcgNeHzMovYElgcnfqsKPrawoeir6n
ko2IAUm3HgRz3cLGQeqULatK8UddOmSx3JQuHyr6ziNvudTONJEgkI3VkiR2wC45
lAnTcrQ+O2MdMH2oy3VtPJKnZvEret5GPcOxmTGDds/qr8ignpoQ7wd9h1eRDnGZ
vILiog6uvt6JRP7cMMr0G/stzzJpo0YQrIjhooZvf87pQOfXtznDwGXbLHNufZPI
aTvoKBGHql9EMu8rjihJaPDTqQpYWmpCeHIpyhE6udK4Ygc1aDARdF1Ff1xBTFaL
UoXypwE8H0rbHk0uoLzlkZVn1VxqCpMT6pfSJtjwFr0R8h1jDgoh0ekDn9Srtikq
uq3pxPcjQQAW5aJMmr0mrx0t/COuVf0IFAhbQ40lUSrhG3z7mulOmZT3BAoQoTDt
JEx7R+qualuHPxdmJORynxWT4FpZBlfTAn7o6RlrAnyxSsTNTSxewAl/wnNu6O2s
//o//+LR2xralPBfodmhbr1vvIDWvWp833ye24sYH1/Hzl3T9GhqWPUAjjQwP8uJ
HDBn89++PWfn9M883IX4MQ1G/a2P0KK9pumSwScOHKqgByga4QuTs2QBxJExwstM
whNPuTiqEHwDUAx/qSdvSMNo9XnX90NbT4shqDRBCxkXkrNH4UxVHCFU4B3dCjzv
NyYZAd1/MHg/z49Na8uewJVPZuPefjGEtbEj6jf9eH/DQ7h60TQzqgkhV2PTad2V
z5HuyaEeARJ0Xa9skz9giMNFr+kwU5oS4dSau/q0Vcsi1UtK5WJGvYnl6P3e1DNf
Ho4cxOYAR2SuBlrCwmqdmjC8BMddSTZ1NQz0KrTmQSb59kRHSeQW66Yl96eYuHvg
c5wjDKs28nWNt5atiRA9S2cu9zI3oga6rEFOOnbpfchsp7kMz1PpWXC7PvxlBvqd
aDt5on51kVtyKotrNFjtMHSX0Z4DxYK4hqOR9fl+cRhjTjORkNoMwiFfIurA41O/
pzKhMPnQVqopA54JMzBkM8Yvp2i+L5vHKEG1/Q/AkMnxF2f7IbysnkEeq+jg323i
5kLUsle5SUGl9Pwthx5nA3XBxVsFSJfe49TN+fYnm027sEGFHM/VsPBJ+UnYceqY
VDX7TVUnya1Wxq4LtTmWGNE48492We9XjPNLTzMjdDPFhVDEanOE9YehwcmNlr0y
Hvbt/qWkKpcFiMkYSpYRandS0tL5AbKADxEb1pTmL1uzBQSMSMxagur7LmFLXvUI
f77P+2Ep0tcxbdbZ6Nl+gpkhIG9JmdV4KWQ7++OEfXSCTmbqBvCGMj3440LAyPD6
yiQRjq3WdzYpcUk0XtukK+fFjcajixnQQD7lcggRHar+1ZZi6HkekUoUG+6r2jz5
zkAl5JNmj5ZN3ol9hf2PVIdK4we3WkC+opubXMlDTu1yqD+VdCVh4R1uhRK7fsXd
yrTQ0SLixorgSxUZX03Wx7RaTbFiy3AQE/kYgwLW13wha2nNnXRvoHeJoWWwstz3
vlTFQFDCMdoKqtPs4W9Nav2lk3+qhC7b/VX0WZutE4j2FfP2MDW/XvHeViU6AR6L
fEXikYI2Or1dhH0Pyi29x/d9KN4N5MO4fxGZLuyP2GKw1ot46j6lhrsWO3/96WaE
axDaxYEZ3pK9KjGeiljCRVTrsFpmw0/tqv+IYuNQ6aklDYSPCGpyNduOXlDG3+1D
KTcPTnrdmei2DSxD0kxBf0sExwcUsH6ix5Kqe2QszkBL1VfmvAsXxAaIqscs3fBz
ORQ0w6wBlMrqlyfJSCCKWwv9lA+qf+UHcITduaxnwR9wJZfLJNnIvvAYx97r5NjT
glN90og1dzohOOEWsyX+P92qchyMl9utUJeMT3sQ0kthq52YVNaHk8p12fgRKHl6
IgNtasAJy8SbjjIlH4jcJYVmRy0eAw+uqfK0+gEa+xgKQixp0LjQPDBdPc8M6nMG
ytOad15i8bPYgfCHshIu7GR51jtviNIfCbnSLKRlloaHyahxHjOf5RquEzm/yrCF
INhrOX/7nPoP3iHib7L6ti5O5W0u47alr0pQV+nl7hOAm0+x+Si2M+hY4oyoSETJ
YYFedYEzfnWiXVniBQsmXED4MM8bACJjbdiojGmBu9QVQ3Jyq4nzOM78qKqPTgHY
hZIdvAVVM84pkn1U8xdwGo00JIqrmFi9OwSgrxFg7O6hWmMTFFrSZxHxSU13yk1p
cD2mGM9PObA1A30lXwU6SWBfgh6xLSW3NcY+cQ5caI4iRb09uPGLBfmOTvI4OXc6
rGDZi5SQ9Tp1k2HrIhVMgXdJc8Jz0resaw15tb0B84FeOPLSao8evtUxE+dtUcps
MG0z8ENhx0xk+UVzzee5IaKRS7FmbEAnEQXRQaohgiisfl3Dd3cqEPWibLu0Iisv
6Rz9iG66T08Jr6WKMfJP87e86bU9gZ17VJXPKyXMMFmjKT9LSCrjD6k7gJoMq8OF
m1GiyHi5KkZ3U6hpFwV0/IrUMJ+ueylvKXDpHEz9mPW1duLLG66JVT7+TFpHd2iK
qv83ZmTsjAuPlaqThZlHL1i06Jz0QduNGZfXWG5SoQnX0//9DtrbQEC10Alprdl6
zz5ivFpLjxiU3O5PcVjpELPtU3Rej9rOohJx8SdGUNdvK62IVknQ/X6JPu0nUE/8
TM9ORqLF3rVFNwHZTP7pxTjk+gqAodU1Bzj/mg12TxhgcT2DGwI0f158AhV3F8qG
AvtaMcuA+ubu6NfGr1XTlG573ccV6Xh1LnWZwnVz5UyQNakLKrAi90njhJMJLOiD
ricUU6R1LpWIqhTmn6jqRUfW6Uwz/Kn4+VfKLyVF7QRLn66hsMphQ8a0wu145M75
jh2Wq0hK8xW8aptFFMaokH6l5tkfi9mdJRs8SuZYmynbKrnbMy7xKBMUrgSF670q
aO6PIvF96EaLOWb76RAJuApEoGIA5rilEkHE4Tn9bBewaNnYcVPHf8GoFr8lybeB
2n4TUJeuK4JhjZgQdtz1e3IPi1aHnl5lMsyMXDsMh/iwo9ko5ZVY9WRYH4Elo6pA
6bav+PCbn9B9Dk1sPkg3a4XougfXwmHouGVs0OTxh7rTTcHFgBtjo7x/GAMy9h5t
wUWsRVI9HNHTegqig44ZhxuYTTCvORXtWHp60BpByZdbdK2d+gp6OUG+Fk4THIos
jTfmxTVtNYq+IgG4IGg3GuvskVbDR748X8pcNCXe1R/qSsSy8bCzmF6zud2mVDHx
hcg+eqgP6VokJYMQQ07ylkqJ2Flz54ISoE3f/kkNUdneajXAf0OIOkX+PoaErB/g
1hWhS5DMKmx/POEV5UH5s/X+EC6ZbG3KssLtUvP5LnmtDmCPTxjE2iPrxRiu94VL
XkCa1Dy4b1KW0cjjUrQX2XbKTHG4wb/ML6ginDrg7YUZSXefiv+rSJ1/wQNySn0J
NzvWhZ+8vcTRKnAKeIOH+FTZ23eG+UtDbnsAyxW2v/AKgNtWv58fcWLscKFYeUli
PjzIQ1NB3HN2I+B49nq6QHmvuFCo4CzIpxw7Pgsc+d/M83obmoPY9BI+LXaw5fW5
1EWvlDglG5KLL4pgNz1d++uIGL7UfGpL1jHPB36U/X1cYhrPogMd2qkxuttRv2Hn
U89pY8BEydc5NgFUfFn7EB4ZKE67Nc8N1QVOaf8+Crg9GdGOTqidm+p9EM5Y6tPb
sHegv+JlbCb2SKGXxM+d+rzriMSa5YcghKj15mwK/+1LQbPqGrZId+Hc1t84ecft
DW5aotS+XNbj4PSDgLvkKQaOPHYlC8nEDYuLdXU98/n8E4DcVo2Q7GkX0LnplIpf
+oTUuqlc/Frakvl/Y93K5dJxEKz0czU09GkqJSrXR3kArFG4PajY6hFyVloBuVUY
/WGkZWf/99ncLPCZsF5pXxSz9UgJQDmaTGgXYeFFc0i1RJeKPvXNyqW8XovBLYBg
DXGU6Y+f5xBuI1dyoou+ss1Wntx+VWzDPvl/9+WAllUBwqXjIrCF6vxW0cyYmdVn
DDF4O9NBGNdC7nsd5ESTrHDgLL58Zh3/XZe5lI4lhddQvEbSPQTFV3751hb/B3H3
bNmep/5H17xG1TnsAEuaLmKGWN/aBpWDmpEdX/lL7ixnfV2pbjV5pbHCsIjuiKKa
f9pxCTiiY19cweEAdBNLJMaQ2R0rGCk2q2G4JGfI52qQMBeXo3B8jP1rD/Sxi8sF
vFendoklluYsgF0neTYpeBFhhNDdfCrGiDv8Z9/FHQ7BTH6BfsTZwSsoB2Y5f0LK
/0fQqiz3mi+G2SCb71YiX5XCd5+f5Cq/u4mjN1eypL/ZflMYImXEkSZNnpVY/+wK
gR6naV1xpAyLd3Luv83f18d/u0qL11jKqvjVflb9x5Tz32xlBcL1sv8qPOQwQtBk
NXOwD7uTBrhCSOJmYostvr3Vo5b5bMWD3akdAQSF4zm9dyuQ6+QF/O43fQ+hW6TF
neHLZQwGBPkvhA++55/FEQDalZYq9a70zzc5+ZypCMLhQxGncNMB/9NuijMS+UiI
mgJI/LH2IcHIIFO6jYX6Squ1CKu3yna569JU3ljyK85PisXZrYai6FKIsPnE01os
q/3XPtdBZ0KkSP6FM3Zo9kOzQ+q1ZekasFAZH2Zm/ienzF9oMy2Uy/462sCAggYo
mBZN5GZ6/zv1xML8FBcRjtkrXzJyH+wK8hQ0q0zMmXeZFnz8hvBWRAfUUU4SX7TN
wIEPhPRE8u5YqoN9F04sg6O1ebnRH8CNdhlr4qTtMYD5J7bLhTJtTfwAPGTdn98J
bJVHvfdKOYRWXx8FehioBCOBdBmtTQYbft+rDauEzeVZJyVhTlpQ4slu6SrZEGHe
Bo2W0QmtWV/8/YdvYqpTNVnrC21rvUm98F4UPGGYxWTGX/i4dqDpkXSf87yJytHZ
bxVvDrm+zLc1XWH1QAMICBkZdPOk3EBWKyQYK3cWgYnlyhQhRAJCUso23fdNSJBB
kyKzsG8h4ZPHnKbOD11nIk4E7jmMD9hCCX7cr4Wj4TZVq1y/C8zEca9iXFsSPrmi
JlrvdBwih+HDUtxOqL2l2PVfj40mfNjG3tkzDR0QZGCxZxy1oGAhtUGr/2/sfeuY
J4BaT+xC7S+E4yZYmbDwCteeiQINT0YBZD37QiTyI9OZ6gbjdrKGa7buZNLgfakD
zACX3CT8E4a9MjW7pQibHPy7Hj4SrVC5jl+hdmgHYqNV00IP17qtTSms49Tb5WCU
nICSzE1ZPsO3fMgGAc1XArNINFEZfsJ/2kBqJLIk+tGrx5prgR0bII9mu0CNR+8E
mFRV51BBcwv1qkjwD7KdLCOFvVuMYMn11kor0lHjrIg0zke7aD8++goNA3vHCnVi
7jQDXiv/GVVaZfseLp4pJU6NIwo9X10zSkGWGj4enoS3wYASlpJSUu9Z3vNqLOok
TgdQa1vp4FKd+2vpKb/zZ+NRChXlFnC8UE04PM3s90Z4xv5/CPCk8JlPzC2fx9uS
RXAI7rF542rsQ8n9+VwuX5OML0JBZR8ARWv8qFn0VOFdNURsKv1rYwu5frL1PUsr
wE5D2nGlI1TCYlmUM3F5gdH+tT9KeBxoRrCq9CFvAuQxoKuS3lMrk0ufCSWjfDFl
d/BbFNOXOtpyzzHRD1ScpcmpOXreUJRCLYlYVgYn7yOgW1NzA0Q2dcvWbwUslbDm
LJzi4GWIcGE5tcCeFqZeYeCEoa5v8do9FEyvLi1cFKK6FkLYfE86H5rQ6e2K0drX
axzCqG0RY46NJIOp3nVnEGsfzieL5Hp2uD9zdIVhb99u+0omkQZIdUdQ/31ZxHEK
WWqsEJhhFUssZ1124+J83tpuLYOtjTKuBaV/8wDge5aFkzGXZf3B965NmUiKmpH8
anj3GoZ5ev1SbUv/+1uaYT0wqBe4hoJG7z8LZk4TN2KMJnBaoFmTQY8yz6J++gJe
A3HjGUw0xgSsFtihDOTOARKj34bLQ/OI3btRbR95sy/40/ZVcImGNEDwgfD3Cz7g
MpWI9Df82+xtggc29fq7JtEhOrKFMJqCjLRJWWjz1PXFTQiJes6fAR+3c/WEmv2C
S8plp8dPTVxn218g2VSiyzEzD/Ct/S1xAujEUWQdhbrOmZ15TOHRIWhsO6ib839D
JZXrdSmlO0eTWHooeS1kRJ/3iS/QMPLNPltIez/ijzDYOs755J5gYzHYPBALibZl
G43XzMBDuEJkJ78WdGfCSxnEc4iiThZKnBlkilP3kzN/XujrsL2uZhZMLZb359QI
JrpRJyS7MtRXSaf6mRWWhjNzn+Ufg+Tvn0yfmM9ZOEeDb79hgjxZGHUMGk5mRm/H
4ck0FzR/rqrHNLiOF/2Bf69UHn3iPcU5bhHVsKoL4cXF5aoiAaz5lTZtCOJS0PNQ
X5h/Uqn2YO91jaWBib2kzn/Lkq55v/rlP5gSKovMneVOaeph0eFE+TfWD9fXCLoT
xgl9la43SjVpGGMTKjmE4iCbMRm8zc3V2Mt6ZlZqVz1cGvZyKtsOUEGmG7zH/mzk
v79VoBHAPOn8Dk+u+7w8/mscHZnp2ktnmpCsqOKgzyKeBgyC4bzJ/FVAvH+96lRe
2YBMQslEWNKPurQrBD4/yBsPMXSUQMpiReuZsWCpPWk8QfTLNw23hCIkpoToQZYk
O1JD5QsCXEOZZ24oqvCzgb+qMpaDMfI0KdL5FSnQISKD4ptednDzPsXnf8UQI/BY
4fYepIumPHE1eUqwhaqqXOXpsc2umOM4bDSsmn6WBNrxOvfzgP9YQdS+E6hjot1d
3c0FDBSVQ3tR7eCgfZLdghRVzE9SCEWND6ovloy+0yH6qQBdGKzhYn07Nu1HvlKJ
DhiRKzFV4ztKdyBUZxoZOUempbmMk6WCSncl6533LggOh1LXdRgH9P3IWnQ8Y4Rf
MYKyshvdj/npS+Hzrt45UfifPSUQJUsrz2SdCr1ug/Qe56nBB9ywY7XsdlHXreVw
TabM2i2ANYbLaDR73Kn2RQBXmSTV6Ty76H4Te8NVT1WyPHlFicJhDa9VonehvWT8
jvdkGhJZnzwoV0hUHpunx3Qi8mM5fmOPwBPV0BTfSiqsf00YRBONjLCyK6lAgmxt
x+Mnt65vAAMAAP2fj0Es2T2KrcP2J8Y5XoKGbdaJLEtPmoLISeiuKXeJni8CjmwG
jYLN/5jJvWXZTXVc/fwk5JSb6p9GHLIqQc5WTQ9/yRntzIPnPqloIUXGEQn0lj3/
1h6EDxpNpCRBAXuLwz/P84bq2vqJktrQ/A1UVUxhIQPQeMMyUhvc+B7wsybDsP+Q
qILOlw5AVUKPj+JTRa1kFTgjHtyzgQXb3+EUCT03gLqt8PDhV3DFrnfX9Zgo8J8E
ocDkt23QUWAZ6cRqi8yX4E5aBfCQSDu2hU2hWZRTcL8tDP4hXyZdvwBDqJGgW/lN
PrxpHtLLK6Nd8t/7zPseyjnc7i9rcf9n79WsgXhkwGQI7ruLnCJ8MUZHojnzKQl0
sSA2eA0tQsyL8baFVkfCUqTABIoovRVeCb2oSVPgC2mR0IGGiao2MnxO8I4h1cRs
6MeCvbFgrhnJGuUnujE2CU5SQXUhkoaWXLSHWBCAPKChze0dparAH7eyIGm1ddeY
ffLo65Q3lL7prjV7gmkMMDfsda1IRyEfvdOCa/j3a7/4xrCzhbtlEGiJKrDCrvqv
Q+XS+ahWcreiOt1Gfk8XH8bSl96JpnT0thle0GMIwWmAE0MOXwR5aqM8jiaX6tmt
O1QSW5RaTznGL4cp1FoEa4Owp9rMl/jNRAo9B4gqT1UZmAvFlrhoRHLPwdcc/0ZH
G5auZqj2R1y2UA4s8W50SSIzwTszfn78DaJilCWiX6dMtcwtFibbHrAfLIzt0Zel
b8UVWCja/qq/wF41L0NiClsDkrAt9c7HvctGiiglyB5/eXu91EoAD8nOHkOJbS7S
pCnDySjXFDYbJdh8eKZHGrk9Ee1zw/g/v/ZcRex9NKhv6RgxubgQvdh4u10gPZT0
4/LOXiKyUspvyRW24q8Hq4n7CncEuF2aByPNenHMRnlYmU2HpSDdlkIP8B4x/n+h
FekJ7MB8loGg1SEFEFMZXcqMTmFWgOZgdNx3yl9455HxeX2asprFlUZYYkI6Htda
ectIWWno6e5tWz1/9MA6cxd0g4F5vHnPUvLirTlsR1WcFeUYmdQIMHLM7gOqaCTk
9ruxbz/FTeWxdbD7vt7OpXDgVOE7pJYwR7Y/50mKBAGARU+Gr8ER51QIXJDGcSet
4lA1YGzDmTOfEJSmsaAnr5YJcOGSKmYUjUmSWCk40W0pAJYi4xVWuqYp5a/hHt+N
UN0lDkC4DsbZ5VoKLd0PR9eNu6Hzm/sH58e1psD0DxnUR1J5R+RZkWJz+a8E8Nko
eJvqaZYvvN0aMyUpzqYEhbCw/74EIovkRSC4rpUBBemBDMI+vyqLUSWaro9wsLn6
GEP64luJcrh/6KTK/5icK9b8VXqTFHOJ+FK43+4mAh/tiTcjLcaG+vZCxM42D6mb
5tlEg29F3nz8oqlo3BgK92NtfqjT8rPfVpqz3cfidHER4a32bW4Xjk187QZ0NAyT
TbZhOc86dZByn87qf2E6/wvQqZT2/BoZWwOOndEeFiChfirfFGyZpT6R0VBwwTJt
PV05AOwkNva7eu9ukNKjXzLyVfRmNm+TLsUbHiglqTLG5puealpreUvbRBgl18r9
ZaO5l1SYkz6riIQeRipjtBYT4d15bTqi6rBNTs8L1Za/wKnSxmOTU3Hev3k752BJ
FxyB30DbyvxiDVUv5oYG5y2FlA+h27vgh7mILEz3/ZofVfcWi3gcR/D5TD7U+8Hv
f/EWBYh7qBipOLuCBMkj5+e1ox36MKH+3EH267ReokJAnI8Sdxo9zJ978S36ntcI
n5THPbaQ8gV797oc4dR45jSuE5V1or7z26bUwImOuqiy/RPjcWWb6KPq2rrZ/yib
GH+4/2pJC19ntZSy/KEutxackrT6bP2ZfFbVCsXRnXUZmJlNaFfnh7jOJUsMMkeq
vb7DqdUgA9mQHhUojowLSvh8/zzDD49kf7BjQg6zos3OWfp9P9oaCD8dzrP1rS+q
SYGvrxD3Y7gM0sPj8ABJq54cLyWaKQuZNIeKhlZBEFtpZAsT/gf8WwdJ4KNoETVt
wVcW1fETscX3LwOj1sAbzqzwwIpUqe9WIwH0j1g7KrbKfbpSRIZv2yeLl0KWIYDF
9AYr7xHri8oOehpLSzYmYdmTcWlzNa19RY/uoParpfyBGbOtMOqGAFH36ObDzdVY
xTKCKH4ZlrHvdJihfZ8kgA2qRSOCcESGqabuu5gzqrCXU+eGZwMOPXiC3i3CVjZQ
OSgcODR368olvPlBoqCAhKCk5GYyCy8XK+t1PROaZPcdRQnRC2xbbJ8vNCekY+1m
NxRbTxHi03ZmbLqpgU/cABZC1f46A+J9m0hPqW3PeJnn7cxoeb43pYsYVoG5Fdl2
lTtpWUQr4cuRvJiKvgmDhwJHnstDw/7wMIITYY88/jR0UMYBoSDhbqmtGESloqzY
oB85Segp8C8UIsE8ZAZeIVWWzvCmIBOXdOyMKupYPARO0lvu3ZYVl64Uetw9JeY1
ApMJLR09PQkEIOo1PsTGTv5X8opubS1TiPuYmhbSsUbThYUmlCyDKKAJv7VnFCXs
cEUHJrjhlg3N+oJOIWzv8ftRUXZusHjCyCxaehTLpakVrY025qX4Kerf4/YI8YQ4
DdnhHDOwdpWhn1536pFem43JPG85sBntuwdUzTOul7G+L77fK4FNO4sysXAgOG82
k+r1kMcGL3NVqUOfvvFuzxPtzaHaNJqXS7vF8cfhBOY6xVQiQUoyA9q10wy58N9U
5gULSz6EFz9WBi2Ca6p4U1lwpPw5qjI/TIua42Ci9gFZhMs4ouuCqj1IyRw9tEOn
aGGysXZ1Ud+LMrR+DEUqVX3z737bEMNZOLe208RZEXJvMPXAK6lGQtiDv7YePTmW
Ih4sYNnpS3eYVI+rrVKh28gDX5ZDnGyNgSMau5p0KhR/81ywM0q2V/f21dblck40
3x7EnwAo8WeJRqjTc1HGHgUNvBzDU28htoX7RtFNfXjSWUd0a5/z5oWhQBPmcc6p
wbCcFQDizWss/cyQ8Yz10hPfNSbJufYVuV5H+tyBrqeu4duewUBxZ/0FMKocNGYh
qA/uGpzuc8zA1hzO0CeJb9nDaqJux21lZK7KRHc93IwAjv2twPW/J8X3IQE8mfzz
M8rTEYWRJfIougS3O2jJtWf8bXJcYzk/5cDF5n6Y5K32V+wMKvgFG6rvqr/r064A
0Z+eza5Z7Nf4FHn26kh9xDPStIrdKWbAvN6BCkQ7f2i/NEwqWU8aMWzAmE4DBJJS
HTeHl6+LT0XWwVevKIIRxDk50gs833DD7hD7/WEZplxwbvEebUEA7ctHuFSrn/lq
B9trgmWeBAKyxBT5yhTcMLMnJtWAciC7Z2gjpPZS4Bnb3l9Dxyn1XrEX++SNrR87
0iyUihGB7ln8lnE7nUX8CWzj+s4tIAq6ULGoi++n7p7LWPggIRXdPocDdm/7OAaP
lOGbjTm3eluns4TeGcfx5UdlF88r+e11ClQA6qgjkbSh7Z5V6+C9Oi0yhD8hEDjN
on9iQUL9O7eRK78rxolU9H17rdQ/QiPvT8mq4R2F14PP1/H4fDZh1ZxtCuF6Umj1
2ei2/MnpetWsL169P8H1Wcu5PLgEHFbdgjwMZo6DMHQNpmnpCDIOf7/USZkJA9S/
k8l+AamHO/BakJJcR20bUox5ryJ7szD00araBZAMVKvQzXf2UEml8ZQwN4Iy/Ean
msKGCkwop3/xLSR8xOiJghruSBt/8oqnl4Acy2dK4U8A+J08HbXKlKYDy4XCh0bg
se6XLmwAquug2FylxUQkteEW/FsGjPcpF0DTSnWWEnF5Pne77FJp/qL6OhKr5ktn
xR+7o4r6jUx2o0CZYU13mb3r1J2QEbs5iz/BaQErRwnzuRvQj6MExhEdw1qxY0x1
J6XqQuQkOrYsxnVHVQMm755xfp1HzSaNrPR5QBA30I5Z66MK0mysxsbT6XGi9qCZ
4CiWasPwvoZjIBtyru10TZVm3r5ZXGTQdV4NbP//32MOG0e69WWMmaiczKNpD7aJ
wJVnwVSifNaR+vFG6Q+3Euwkk2WdYsTBeta1Lcskab2XgymiE8ckjEq/sW5KEWPY
S2bUFmOLRk46oP7SojJE/h7GgksPfCcX1fJt3BtLt5j+PSoPqAu8nyefxzNgvWqQ
jj1JYjdG87nL9cQ+mWqw1Gi1mR3Qr2m111B0HRwH2GWs5K/75yyTtO7fnIlxFfkC
uVzkrQlrnDaQpOOhNtPjOyz0s7F9DczOOy7UYx0CFvR9jLyPzreoME6dbBbbUMcU
M4PZbXX0jatqCzoV88nwwwJWMV5fuK5fCcZgXRtXSMSrhHLdfcgEEjocTiTV8dz3
q8ynoYykLFkX3hlCJ2Cui/ew8JeoYlnUDapT/+ziqVnoszHbv3nVbNqrEKNoPYb8
YrW2vbnXFehAva2COQFOELuor+wL3n6cNu9CGa3dD6cBVNrDjRaXig19KUXMkPve
G2Ia8wYKk/NzP6IbacijxkJ7T0jJRMwRln6R0ZUsFNLhjoK+4Gp2Fw678loRk90k
FayJYvWgfiRqMwH8awjnH23rGdBBFsQahfaW5JHQWEipYVSiIRJJ12C4cd8Ox40o
RBGEIl16cvj/wUoEwwmWoXSUtWFHpLujRkSpIukH8pbF7m7CPrng02V9Z2giN2ke
jSgZGD8dPzJmSOEXQCZs7xdYNMmIMr63rOTP535+ZsfvztpZulalVv3da5LHBUEb
yLXwoc4e14I5LgzoKCfiXg6OCwcbTlMZrRbnITNa1i3P3fTeDG8gSp+1qZElyWVr
jSf0eTQfjXNf2HShxpT2b1uCO9SK1QwgDXUAdWNJXZZJ/w9+WKPFQdj92pnyedXf
92cC5Y/csrbXPOSv9K0auEQXOmQ6mcoZBXESVZrKDgc9o8wqQwrqLg4XEGikNmAI
6w+48l8SISX1Is3rtLqWflV9ThRiNpe7U45oxybnmppFZMBD3B3OTRNjjbOa5nwo
9OMrm64CQUSlSwqSos14EvP6DaX1LpgVC6bQZOBwmOJNvUE1F9nGN3m+Kj4OHuHn
S3oO2VVLSFJQ+5/vFJ9fk7kFjptljyp7evzasQH83GRm4Ri0hVd8R86S7nGij3Re
HtXNDSbIELOLRfLrxePZRwvnDqLy7zJiDOs9kzJL72pqnU5nEoqAgBXyKnQaas1o
OBv5mwvmnACHVmbrOuJNAfQp2cB/k3cyW/G4egrmmRjiWqCGI8rrzByKVPJ2kQCZ
aPui/VNFloLg4CbnLyL14s/dsifW09YpCZgZTJHoDuxZdyatvkaxiBdoeGbSPEq5
CXa/PJh2jbrgyYZgxV9OCyO//CdQ9R3x+kw2/xz48qPKQd3QdlQVvSYte5wV3OyS
crHqESbCJnhc2vVxiKqgAS/6bE2dO8ONnYS0XD/hJHQb8wSs1ZKHAn7HeNRJu2Kx
eKsxNDekJTnIkkkpcRbUxDSNA95c5E1BPDQT867GnUJHB6lzBrXe37hhzskc4f8T
E5EDzk8YWL84FvzpD/rgdWDj5rELHIhLyIvpWCrehoeXU8pmXPW3ZWWcBoCFUMCK
ukgyUlJSR06KaWVBH8jxgNaZgmWyYOSUftNX8VMyiAbaPm2uCI9EiLPeBae5FGUY
jfnhMQ0//M9ZtTYJTJWBOBJI1wnfUJjl3WEiDOi2SRaxYNAvvBcsmqEIl7m4pLqN
S89z7GYPD1idMnH0zBz2wmov42lXTQStM3Xn/DmHANyK4Zsvado+AJdL3cVJy5G3
jEmYDm4Sf+L7Q30/4F49ywxnOJJEPjQOoggAK8Kvu9csYScMgG0HvKN2qmoD+l9I
ZnPTL6KIORGEFMMSXM7EqmoFXBjTWBxDHh1ad/cAEA6E+J3Iah1ROVPywZbQXwDW
/5FY95PYWqc0sqP7jPqwjQwQSG7rr8JwmAO6fgWOBL/lkzsHEP3l5X9IYI5So/Ii
Peknw0mHm2WdvWJQGWkMGIK1+pC2FjMckvv7vGhyFkL7NRS7lwuwXNzGvGm9iWGA
TMHFlgGlrpENOlCu4YqkMB36IN5c0mOSLmuioosWpwnzpN5URoPCeo1vNJsLXfa6
yZeNgLqcO0rmgI/Dx5BGZwA1v82zhlMyMeslWfR06EItFMhTcstMsuplUXDXHuKF
5ngrToQHUtpX6CuwPWBnPzTUupjweNp87htKw4LXXacaAwKB/zggFrFrGk1RQUdI
wTLSvioDgK9Ke4K5tKXWsZE/OQAKBKaJtq0ohVVa6L5LcekGc8WiUWaV0gYtDyeg
hiUbxt6p/HfwnaZ3SbsxDBuwVNce1uG4JKObHAcRtnz4GGZGBs69ZIVCWZcqa4sq
oGmBK8Se+3Is2tTE0Zd61kfFnLVC2YeJHbKqABO22b/Ys4T2I4qLEF59r3RwrVQ7
35JUkJcxRF1PvMKk2zAfeqCJMk148sPDBexdW3zkjEyNkkvauK6TMGKfBcjNXS7B
w30o3yV8hsCy4wqJoF+A5M/docfPmrP4DwsoFeiU+Id0vHr8l7iwrVIejvTqpvl8
GIWvOG+JYFxGEbBR+FJRFpUeliclWURuGwSt1/jQCKSxeSh4Bm0kbkTPR6JfzL1e
o62k/3ZKADXFLh8jkgHVL8X13KI7eGi0SOdR1uQti39mD1GzT4C3CX7oPEuWU9EE
6DH/Nv2jW9iM5ZjEXDe6UtrbZ541uyCDF0FgGmdOucom0VqIyVrcG/jTCyz85h+q
tLaWXciY1ZjpUJyfTbG1f3bv2qeK4E6/1iHZdMJMyNWW0UhMsquIihsX5wXMfn3A
+Uj0CQGgglihI865U9rdKwL6ZwHDBDWUB5SINLgs9QY9wwviDLqJRb6b2ngtlV8y
9nNJE9ZBEAn5NmR87K+wtDFyZTUUgLE/lqg6BvgugwfuEh/Zo3hnkFOud3Rfbq3E
MyhWqXIqAQVp4Xp/6QhKF07lS4oF1oi0L+wlrItA/VUTN1lsMLff1d/M2BWaqZwS
2MD/VOUM2Ok6IMVYbpYJHWFDJFn/1dA7JnVJwOlXbp+/jJs2TCpGbjmw8Vzyz62t
nWnLa9oYZ0wU7vJEnfUq//kOIbafz7QeTvBS2fFfUtHZzDtmA9FiTwoiWkPqd5i1
qQjIlIcYUMhRyhAnGpgnvIGrI4eF13gtCMni35Jpmh0PhDH0osLddvhO+9l1Mb64
V0ODjBWLJWSln1d0AWRJZP9jpcHhkUqKILtGqSy9LO6g060MwAEnIDtLSrMBul80
eh62KcpCrEmGjbhOBPKGzS30vITYoBsO6btFu361e7Ay/+p2IrxNu2oaT9mimhgm
L+UdhV1AqbJRUwAJAMZlSsnzWPSnMy+zbitLkU1RYtVcuZWYFBKDqzeAi0uybn34
ZER4tiVh3Ydn560Aqq7alltWqV3kKwKjlIv0M4kRvI6/CnKExIdkUgfTGPDeKvAv
flgpLirnirAemfmVSaUHckiqCNOvRhrtr9ehRrgZMsUIaInBmdBU65D/vlbFnm7H
Cky7yk+JF/iv5q9d+ysB4fIrH9M6N3wQPTrUpXdcE6Nymtd4Rbkf3ofS740UmDF/
JPXkvZR1UNJhKG7mN1KO4hJhP+x8S4QTdtDNkToekk1Lx99IKMsYLuuURnIbAQzG
pF6krTdHxZZwoIyh1XPBF9OWVYOPG5MZDzo+gdOc1j1hh+aT0jFWdGLCbEffwm8D
h4fxI4X9q61LNLSKHGTgMDwQgpzRMchmIWTZZ+I+RUoarfwenYA6xbHaWOacXosc
KFakZEeIvZFEAeKfo1kzsmKihom98TM2YwTRe9q5qoZxMre0avDVj9Y0GaVkB+pc
R+afrXWeawUIq40EHKT8Hw/SLLhDShtfijdSQ0qRf+e14fl/ilbM5LqztYWosWNn
X+YoGSEHTH08N+8y5xz+aSOCOfPwM32bc6MM3f+qQzkGZn2W1RiQG+Z00xCHZ3S9
noaxIQd7v8GQK10EsVDJ9fMEwyVJt9nHpFAGH/ahEMGYnu9QS3qTAzKAey/+Sl6Y
ZQWM18MBLgFkz0CSkJ21AXJ9BqN86RahESZD4qmAAYDGg5RGnaZ7F6LPNtGWgi7S
UXcu5GuOM50vSrhWbfu0JKdRFJzQ2KyIFXUopYyyMDFEuWj6raF4xFVlJ1MuICK5
Pbsld7fUCwSR20pIDpZ6boHIzYPYB7r59Y3Zx7RF5BCQx3cGtwVyjpG7TxISXoWB
cNS1JJvycifCGVDzsQ1gVmmaOO1IgKtzV3TBQRQmnf/SoJ4cGFgsB8Z3akHDbcGO
7yeXUxQeAmQ0yjqi6jQKy7cxLPs/TB6hIhYgiRE+0SAlosJraIFOH8G/MvSrXWNz
LTGEZQFlskccN53RJ8ieAr+FkyHEE/PbCgIPQ895+2aDAdJsLaGkJDkvpYReumRI
XWiBt3QOMNBjmtv7hcj8GPUJITfRweIZSK4Tef2F3ijxGLZ3ge7JRJc1/bWWFo/G
2YO2E06SMkGU47BiDRnvZi06D66pNurKgwquDioMBLVzIxHBBWrJdk530Ii6JaqX
7zKtywdZQ0tyJl90xlvyJjhbA/RqWSY1OqNtshEjHByrdCtGc2VIFPQzKbfvocTV
tNOVSaDJg0JURrkzk9QcOE75sijaOuLhYnYaNohCyK9MP2dxjBNJ41wStOJKA6Js
12sFOaXcDErWEHgOxlFEQfKco8meMaWeTsHBrIZCpqhUO9DqVy+Z5i9Zcv4j3/l+
BJR2uy6jCYS+EZiNwRo5umQkKZ0RYahL4pWqbQB26Rjy9jFopDWhpisQenor6xnU
kypeJPq8Fm1K83g5m2d/+rFLt6PTFZnpeEifFd1FTSmxbjPRc4WLiSBA1CFsuPIb
ZohJ+VotohTO26yJdoRc7HGay0VWoctEdcKXETy2iX5GNgV1I1ngHD++aNV5AkfP
nCQDCDMpXWbBgOtj6DRDYHPqUUL8OSsApwW2CLzXLmjRB650t2FoedFtPbFWtZ4S
Zgqvo+okqXCu6Ftvo9OLsnN/R9KLDPJP2KSj1ydsm3TxvHJAcftrTNho74EpIpkK
hEB+qzmRYXkj0PgHZPOBUtCthnkDuxIx09wonrWdx5q4tQQrR4fwKbvRMPg5idoD
/rTV2LiL7kfKacc463W4UW9vXOKR6FGxiNMQZcTqC+Nz4YjkGcqZjRlejI+rrW7M
dQy7iVktH2orKLnzJ0Gpr3PTWtZKnJc8xhr7ergwjMx0rM/a6qVS49qkbL2eVo4e
T5bQEGnjLNAEwvV4uEyFLjLJj558Rwk0mc6FfkwYUXQvx+xCV0Hi22OI6iA/UtU2
XHgvDQ4uxE9NvTFemY48DX93mRmwScBBhxAW0JRofzi9yU9owey5RDHhDzTQPcf+
ySOyDB+8WlZFXtRwIt2xltWfGkKFn/DEO17aEu+miHAUJAV5W/g79diSbBv5s4cn
LHVCJbNh4ZJgrotiAaHDTNXJ/LYtLUg61LM91Jacuyt7u/hTitSSv4Wz/thdO5Kk
E2wpKbUf0vbu0LaBKIlZBCMUxWh93AXSXdUhXKkut2fHgD5g3pDGpolmZBeRO7sX
w9rCmeoINfQEwimq4DqWSVaznxY0E5kipYQDQZMb4Z8qQPPpwkE5wk6RIghI0huO
vWS5+aKo0TflmBQCwozYaGgOoUgQ2iPYcG9HtitvERYxIa35ui2IGBk+40Ta2Z/w
rduQJrKkT/isckIsgRMAl1reQyWYuGG8E+AqG+F15kJe33QFTUH4FM6YanUPsNeN
sWvbBtTN8vfdaa5gyyh5bELpD83Rb1kuksDDtQGS2/5fAFZzfux1VS88YpRNKjau
1p++wl0v1B67aKKHHB0Rk1DgBzhJ0Dgi95soUD3RpVEsFgKFz5JFM8tAkGzD/PGL
L1tM3FRbSZ7t3j5oGc4HMRpA7Yaj2WfKZ3uKm/jZl7lGkDUU9tOjVBLofaR6aPut
qoJbhv+WX2p1scRMTiL2/NoJ/5fQKAPF4Dh940cWCJjrrnzsukUrdDCuJYjcIRWU
XHAhiLaZ0A9syA2aUlknPFedX/30cR50mp0H2e86Y6kWeWDXEHo0+hOXsqvvK4T8
/EYyc/hDKDoZ/wHXVjgnlSIwL4d13NjZH7r4gkWDzVXcxPAIstKc5u8KOzovVN7P
pNlpZ9FWd37RDn6jbG0k3ELSHGWR2C3HEkZ/vCcGFISBY5vieGZHDrcvnr9DsBYw
jSk1Q9z+ggWfX6ORYHjDRej764iP4CHQfF+Y+AfS4ZlYUb2nT3NlKNJ8z97HjHlJ
r17r4T117yjfOY8L1Ek/d6y6zXvOB85Cjojq6rrduSoV5XmXFGt7iJLm1ZP9s/9e
t3/e5SUc000qrVAeE+bAswX+aSf1f3EGBMzj6VOx0VD7bgo9DGvp46svGvsAWf7v
3H2r0c1Go6G6xkD9e4ty1VeK5/QF/NSUjqklWZpj8mirNxX/RE71b4iBKsiyCuLd
KnYxhaTj/Sjulr3XXDHxWTmGHnT7zYVXMn2C6jsizybEWTE1IesRiAJBgagJXEhg
k1pwjc49vIYcSa13NCvcU+Ylxv4BqTpLGxapErs6fCI/YN7Itjk/NDkM1bjR0ZWq
7Rm4pCQHEo1jtLNK6RL3BRBVlAvY9Kx6d9RvVNTTjqAnljamxzbNek42G1x21ktf
TjSDi2McUhW1Dr1cKB+F15HQPWnE9BEn87HW7m/WXbtrtoOjCIw5BqbnmAMrAvQH
uiKEhIalM+HU9R43g9v2kjZE4ekwzqpU7JfKwimjNM8gLWH1qyBJySJt8omEWOEk
seTTrlrReg6UvY0SW7+Se1jB9HdvYj71EEGcGE/OBj8RrWYC0RNNdJIJeJqu4LUk
jOUCdhNn2XEVLR5WUDa14MIMl7x7L/e5bTmGxHNciyk2vxdNrMQ7BcY29QRHiEKW
QbbbbeD6jpDNlBARU3L/TKu9m3VCmgA5ZY7yUNpC6deJjFWFjrWfLRdcFGPXExvC
m1Vgv4lgG5d3MpGOjfwdAbyQqRYrFMGZUjsA1TM0DeHXu8H76CNLjXwP8j04ay3Q
Y8K8ECS74lhKDqPXfVmwDfaY9xBOCTcXu/JYUvg08UFD00XLMD9o1YzFfY8g0Gl0
3UbTn4YhuHgk1+9OqLZEYsyEwDPJebX/RRpmC3xC4nJXW9FLWWgq0a1caIXv1iK/
gJFDcZakp52k1H/eNTGDds8uwPHrbBcH1ByiWG+Q3lTGZaN8Vg3qhrFspcp4V32U
PcyxScuiRxdoWSdMnT6SiSw28Va9OgYGsFfSop7AnbJIvM3vKCWhsF2vlC7xeScq
HwCiwSpQa6eBbRiLBFiqIEo7whjWbrpUKgAN/DlMGu1SItgnl2AA/cpPPJwXIIrC
ngi9AF2lDk3PEgLU3C0047e2CBsg7Yx+YhcZKZplKWdIBKptnhQTzmPbVYUzqgFc
0r6NQuriQtw8Y74K/8I5WUBLAlhRCYaHCb6+Da09DW9/seuO8B3yzMOp7XLDN7uY
r9mfVXqMHNb1X8FRZBNA5Qhhi1AWH0CqLuh971hVEtuJ9Ed/cdazOq7AdR3N157L
XW5aomGnESUl8Q5jAiv8MKsBO3LTqk+0pKHDKldJq8AYlyJT8gFPw7icbWadWl7G
3UyeEf4/dcJHMHydlO5jIkH3vbwqFex3tS/4X/rCh7FXqFNoTkRerfyFnN7JTyF+
/ic5Jwz0Uzxuw2zygEieQ5veOsw1JHkM7BF+FnqdaJtIgLxneOp8CU3AZ2LQ+Yta
3ogXkOay012rfuJnmegYd/x9T9icmQhagncWaM0u+PVEbVaDLUhGQWEhVT9CAJwo
YVYKoxR+o2ToFormhRHE7kkiERqpEXyL/KD0+OFzh84qQCkJkiIBDyM0bbhlLGzQ
s7H5rk39Y/0B2HK3U+4DlJL/Bmg/VgkGMRnHh+NVlJux5HoqOqfQujvNqKevDc8A
V3FGlFqc+VRmPtUyPIM5ooQ02PUAnAEAmINcm5MNdBAh67+js/GzY7qdQbgYmyAc
V7e8v4tbc+vf/0pM3SIrXW42m5nGMGtodxGAKO+uyVSe5vA/PSOrzufyfAWRMmaJ
NnGywT0ocHEAZmyWZIiVAjJp5kaSmLmXcnw+9tsnkERdrKTz5aBKfK0oZFzn9PUO
uBuDA8+x5qM/HpSkxIgA4UJ2ocQSVnXCAZF7p/4U6RrrC8G9NFDK8SjfTiyYJw7K
/IZiIiOe9lK5TNCSLQb2m7fU6aSA4yq+r78+QSm+Lu95RobYW4+aQTJC6GL8REI/
CZOvtv8gQc/GCq/zvFut3yg6XX1ZsoySb7aPd/cfms07l5C1bjUMAZ8zvySPJhY8
KGs5jpHXijPYw1thvkxpKA35DAKnyKdXhYvCydUC+pub3DSrIjK0fzta4ND5R7XB
T/CdzHZcmiKlXPBmfHpZ2PqRPQKDU7CnmNAaJt1kjIBtWqXrtnKFE7+Rr+xJ054O
TEMwrs/dzmRAmIZ49U/SQlDVEgiDsYCBbDPt9yDlBaEqSPQwNFJLPVg5WmeHJKTq
mtNkXJCjZL/gSgVsEcZ57Qj8cFkvE8aIhoKpTnoL3O8y04vxjFX4fwI2pcuJ4duG
3GOe7ZvRl3JRp1oROqz1+X0tlXqf/h3uUN8wKqnNFHAWt+3zFur+Q8Gh5g8zEv6t
Hf8QoWkkqGsam7/fYBKsg+2EA+/Mz28l3tdy2LwsytxpUpQl6lfX/kH4NYOGFQnj
mrwtyypEEGgRRhbOpns7QvREvCM7eIxmtd/EscF5yvRTIa/1Arm7bI3Q3MKGAdUB
VObX0+f06tiuAYXKzEUn/MwVWbZ0+57sZTRlxSUwpqe0xvtXa4++/SewHGQxynlp
NACHjSnirfs6zHsz3dvnndi74BbT+vqU8XcZsTgij3rvkaDRz5wrHDklZGPm86XR
ve2DXxon7YwGO5ihjylhMXMkcVeHyjltZMvON4wiPOTXqGpipAjpNcCLGKkaG3CS
N5/I0l94d5e/ltGsfULYcpTS5h8oxPEuen5hPtg3Vw0M8kaSpbLA7un5TSDXqay9
bXaehvvhmiKIfUdh0R7vHpw0Q/L9TP7iVPtwqkRKRFBNqfZgJe4Axlni8UPyRi11
LE1F++8ZPc/rDcbmmS1TRFBCzq461c4QZhgUpxHuk2SNibL8V0j/McbZR9HXLyDA
6iqJB5FSYYZOLMtUEPoQDVgzVnmz55LL/i3bbFMTjxk4/VNS5sSW359GZNZe3h9T
guCT/kwJy2DOGIS645M9We1yFWqN5uIfjIxf/0AwprgidF+XQsr7T9JQ+TD5iqkS
sQrWN844/1+CTk3ceUjJORFBepWeNBCUmYSxAwWA6n7C6GC2APxRSHm1jPF4zOwz
IboCUFSWbAVbmV0PhystiL5U02aGN2DyENvzhtHbPPFbtoHUyqQQdbFeeDA1mLfN
3xDwU2ah9DkY1bbkFm5g8ECCZmcL3zBR1AGfnQeev5EIJkudygNQKG5knPMeO6Wr
Vgy2X5LdoXbAGHZMYVhBvsMyHcgREymj2QGXK8Vf7me99eq+DbrJrwWJgc8OPUIx
f3R2CmxVhKIrEy1YVbaSg8xhQ5wEbvSII6XZbbIYAjhgfUToinevS8iEhHIoF+RT
PVm1+2s2vgMIp9RmD8KNyGDoa/ZTuWixP89WQIDqRHKlzyu1sO8bSfJm7bDJIokm
ie8kJntXJA/pKeoty1o/ZKjZLvvnTCCdLXuouCtKw25/gEuUXIWanUHll33VHfC5
ZfXfoXDC6s5WndEkrEmiljP4jB3DLqlUyPFqdbq8Tn+11bSc2SwUELGZZ5W4UvFc
PUOxkYTWvMTu/pKs18Jhn7Ju4L+ZribD79P/sd6UBzSRNxnkDEug+VoblhqT9FBQ
PwxHAQBRIbiMtYUEnDBVVhaKET1Q31zg8a6Au35SWGockvOMPdi1EbL4AW0vDS4p
bC+FDKnLX+NUfL/kUU0LHyNu66FJB9nKBiIEoKS4m/V1Q4ISo1fqgk1giTibl5lP
S/FJTqsylIb15i4lYqsyQTvsoyeLRtW2G7orM6+ReOGfqwss29s6FmLPwjha5+vl
WROShL18DCwb0U9zg8dOppXjnjwyz7uLSpy9RQo6ZV++OZcXnpCcW9CRMVsyIobF
a0BXmB6SD0IeBonQ55bl92J9OuHpFwPoqtO8lWG3jRN0We/VQOZYFRGfObKjgGAH
PcSDKNFIq/HFXsvVqd/LYLNip7q09Zh0NG173xSzlT8q/ZrfmqxQByXr2s6YBOCl
7gJKAMWhzyNC7dIIIUXt/w/fL2m13ubB8HLj23242YRpT608A8/cxynq/mQ3P8Py
G3RlkRPMX/X0a8gT9ybbXkgnNTqN90mTKKM0EzZgZoTmAlHlFTZ+1Hk9MgFHIzzC
rgbaLplTybciPNcamhUW7R/a4Vvvm44tpvxT4hb3ZeD5SirFkhMZaJAWAUmv/VBo
5TGSGNonP5qAs5w04Nx25eML1PfbDOd/FrvD1iGlQEuOg9jrD5QGf4XirJV2WrJ5
zNxDDqMiWcEHayktKaOjNnZ9oNKnTXSmYQE1odh70tDThLqqoxyhFe93cVSxIsHy
sMz1BWBzVsY5+PUnPi1FUr2h8a8m2yJIaCJek6GLSZGlqTXiKW3R0SikF6rck/yb
GZNef1Z+xjxvGohF69tP4ERW++rEtzZAnoXW/dtvUgfIwC+dhcMpk+hsdDdhg/Yb
5qD5Bb4ZLVfoqWLg2KCVFOBp0AwTiNX73q0g3a3DbKxzDvfwSZzq4v4TmxBOWjJr
840rKZN8SkMoVULa9DB03W+9s3AE0ASWMQQoCyckcIPbyjQyQ2B1PEUyQgxVFrqX
QG7h4iQcdoxdCHjFTpqHksKbV0PcV9UaoaJKrUY0oC3v4q8VxNlWLiabcKMH3yCB
m8SMI9T1Pzq0mNuRxW2MD67AA+uQWlfnMRD0TtXuI4GOUyOx7gy7C+bQTTq8p7vS
3VWSB8DyEYgX56NjDYp4MuJUZY0CSmbCPeqORBPAzx5PLECSzv599z83KR7bwyGq
5EV8xP5C+pPJJMZIk7zZ1ugPtG7LqvOdsEGZESy00Dd9bU3FlJ5vUQCE8fjyr9ss
zb3bvQnS4X6ncHVT5PBqjfojr1CiT2lFgQUbutnCh3DqtRmrAuH3p3ynol5U/q10
sFG6AMFPP1GjcUyzqbbwtvmcDZrcADSmgDr/ySEtSLfWOJY264mww656VdwPsM6L
zHjFJj3FJPMIe9DoKpLvTQvyCLmW4rcxcGW0iJwed/MeVj95Z45TyhYiBfVK9X3L
aKQE5XN7uka6YcfvliEgN9vY6kfIegd3upg4CHvp6HU7P92iEMA0Qblzprc9lZ9E
r3kmBiw4g0OYudoa4cWw14qMaTdJmRP7HyBVK/49wJLQL0RjM0M4wo8v0VvPEo9o
SvF/XkHug1xCWSoUXhyaOmMjVPY6opdbJIIU7IVK/k2KnL2Z4istMw6VVWF6gxMu
0/vvoSvM9aU9LlkwmpMow9KnSuVlPcYIyR6INtxJTbID32EOi6DqPmGsEFTv1Tma
eHBA9dFbuoJG3KBxfDWcOz4ksfWFQSKrkKaLgx/5NQRffoJ74d7Zn0+NcA4FWUPx
szfy4ZxVaCmq+iHIAIbKaOh1wvrXD0NurvbtjlIbFX9Zd/bx2WhSahXnBIKTG51Y
hd40DS5Q3JjEDpfFYX0gd8+KVeD1DXOpQPareQovtPTtCz5BsP2r+urBqgjyy3OJ
2pZ34H85CEwz2KgF8DEw0ibxHl/n51lBOqHp4xjdoB9equp5+UnC+XHRQZUOzJh6
KoiDZDoKt3JQ7hEGogIj7rLWC0jedvtYAE507FaZKch5mZplGwOuwvOznT9a8AM9
pDNvq+e0fZM/CvgzqdBZHgqwGrHOOyL8LZETg85+8CMRLF8qS55wN2bFCddIq6le
9cQXSiv/NUaKB4WM7qhCQ4okvEvDQTwjFPYF42ZuWq6fRW2rSZ1VIvS3kTzqSGR8
/Y/014I/kO8J1hkL7N0oI+zSwoAcQP05O4AVl/ZaofPFRRoPgoYkB9+vkdJVZ1dH
UFY+arDNAjZqyUtNdx6mXvquYzCw5RzfHhOrjSwPjbZ9wUYWnRB6hirnh469AGHy
v9PFQ4+DY4tq0UqViEQCAdkYWocy0PdpEmVsvgu3+ipLUnELwATg8Y1j2O7hbb44
JA8/VC+Cot3IAG1H0a0tEu/9lLM3kMgKbfzXWXejXuB+UbbN3saZH0PM82F9Y43J
YYoFk32fUxc+9/hvWiTZHog0IRAuhy4w2Ld+r8A/yVvVLmsh3t3IoKu6SK/3Ss3e
ZmL+1fTYCWPWJnrmaP3bIXGZhN0xGkTU3rdatCx59dU8JFFn0AhWejxm6i4ExVrF
DF3wynOc2slSff6dMjbObcKjEQ7uXk5ZQcV7t4eGZJ+Wv+bwa24IqiINMTaJTUlg
54WlSbAV29eCd2P1PUVDYlYTtANeYBvTFE/YEtVTw/QhCho2IG17/H5XtVhc4qpS
CAHbLSzzHDU2sABBbvzDIgwx6gvwwmcnNpr22EXxci0QRVZppQM9cUkJF78lGGv5
rBqK1hoe7kfEALa6k2/Bk3eEwLsD1FmH+64KSkl3OUoSQnvaKtYlkDxhTALsICtp
eT7USfcRQPqBReYdn8+rDu+HE9gJqLeG324CWdHNvgD3SC0Ak7vjfHpu5QFPrvU8
/ZeiuqERW9itzSBhLm7tkrKtWlE2pyTBkMGRiAPtGPsgmtIZQAbzgOOtGu644ubG
YmRz4+UJaWvuGQMJAmnLro4e5EF+c6FV7iuu28uP8kptj6jnKgOUn+AhxsaPozWq
QZ/SG/+T67f1c6ul9JD/igXu7K28RXxjHi0acavZiqurJFeyfOnnqw3FcitKqtVz
N4nIkrQEHa97g7jZjr0Q0ZuLzPgFb9T4Tmi06Yw4vQoc+Gy4DaGnte4szfL2fWfV
BNKCLqQcTy5BQH/gYQlaIfNqoPVmng8a+FE7WRTrPF7hsFIXpPpv6pz8Iy5mJng/
WnGgiUBN1aEhfq+wI8+Xw3wVxcMVHaZQuj/VoqWU9H2Ft9fehSHjjYC6pJYy8LIv
FR+iwyHiR8f1GqmUwdNuEFNTT16rpW3EcBkU7NYmgxmaNOEaHhxt1CqSqk61kmDa
BYeyJ8sVXvc2kfI9MLejH3XWruAxBA7fKk+PeblUS0Q61VOfKl6AldoOTVdCW+59
othqhEcaWppz3i3/buzNcxkoYWhbuFQuVv6Blr6t6/Rrg0NDLItKbL7LKI4DWG3Y
SwO/s65DsVPn6ESHAEqFnqcHtbxYMqULQR/QnFSoEYk3WjkTidfqysm+Rw7ggSJp
GjYljY9vQSlgwcVzYKUMbPfPShUIOO7Y3E5S7izoDexmZvepr3wQn/ftXPBJmjq9
Yf7axQw45XFs5iXaNKm6jFSMJmY5cqt9liJ90YxLkV0GGqhQdZcKS/GqaUXaQY9c
Encwx51pC40CvJx8nC7ozyCvHbI54VEEbLaosMZBXBWz6pw0Gq2pD/zkM+SlTKJf
Co7kIwbAe3pulsSsAr3MnL3bkZmVVcv6T8YPKj5d2SzB6FPnOFHulJg5h/3TLbJ0
GmtmslcS0gXoqLd5Skw9oxfAVe5Bj9T1kjsOo2NrofkrhQlCxWAMOIYzcxagwHv3
Zmx2K2CxoHxVrOKYsfRzyLuH5dQ2NNx7XsqqYhlBnIP+E/OUB9NL6Zf8bRia/rq0
X8wR6eh6ML3HyHo90MNJIx1Nkmz7IXYbX6PA8cnp/uNyd7/nIG8RkuXXO6fiazTg
YuV8TBqNBEgxm5hLNgziZGXrLviZh0GMAJGG53Aw5IRJHfJLa21dRTuPnBLStFUQ
LOImoTlwV5agJgoQoN2sRUQSr3PKr7jS17yH0o1MxrlzdQ/PqkX/i0hjfwE2JIW1
GVwIPnjvZGh2Efi/buttvXghbKcQq06xBPHVokIr8+psWd+0jjRUrQFo/Z110qkZ
Z5o0Zsf8WZAc+OvTqxmGi7H1U/HVTbswl26ay0JROGs/gvkCTzgVhB5SuB1HeHzK
Dc7N69zdjK8N9jom1gc3QC8Qa/Rsh2U+Aogo+PwZ6h0M0nBgtAKffBdiPG2l+uhF
q0FQ37/qPuyoI9CBF7OzFoXiT0l5UhBYDCMKkgiHZxVlYKhpmjTPlhXhr4RnKszl
cRyVgbabzH4LZHPugLdApay26Lz/qYau32AdpC5g94r3kBSunDV+Zglh+07ic8K0
yl2ggQXGQODgDR4sT7o+B4d32POVsI7NDFgBjNQnBqO7z189nzICx3iFej/qQbiR
cyhOVZDSMHRQ8/H4FnFQ/ntCvxGVqSRQd51HzL3zRzY2bJIIg+40c6/Z2y+eEq8K
486iFrzvEck2xff5M5tYFrJyX+FjBil/a04cQHoavQWh9pog+ZsJxjNMY65izxm9
GNHK6Qcs32OS6dDLv/qZ371sSljDaUOTmsJ3ASnCsbQ5ERGpPsM3G41rM7ABCKE2
NZ6LGFHRfrajxhwDwOisbpkr5GhR/M5uuqTymgVV5zzRGug4km12dQyGC4eW6PTt
CtO7vu9NcJsTqhpuee57zd7SlZHEPz6z7SDO1//DbTPuTiysuyRrOnGuZrpPyGgE
+OR+1q6KwC5SXyzzSmEswP2TWpU4akceZ8siWL9o5zfoZedmxMTyFSV+OT2zQuSY
LcbC5LN0no4m2jUSWsxwrBvATIv95CHY0wJ98xsoiBas+syN1vOvBtuuGwtHUERW
+KAjtFEHOHfZvUlRP+4FwHkyS1zwj/deXVGQIVGcbP98yzU3faNEcZNtNt5yJ7kB
0kkDenY0YbPuqqVec3gYn2Vh8Z6bZJP0mbhXeyx5GSNlfYgNo24FCN5ofrYxVttL
envlUwWlcoidUGvj2nClE3YEH9eNhDGFk+HMTZsbVwVugjFqb0cg9esyZWuMlXtw
c7S3k3qNlOVbpJRexY4BwlF1/hwmFOM9tbXCqqoa83MuI5r5XFd7kW9+zDg5vHww
Jg5d7rgCM/Vktl2p5Apx5YtKd+TI0P001wryeAImnJ9A8fTE2m87XscyOBOJ2rh7
+2G1H31kTlfYzny/lrOOFMbFpgSkkaSI2DSiNEG2vpj/ikTky7Lj0mLaHED+2a4R
HTNO6bXUOBag0ruLEJa6mVDaAJjmDppb0CulbEzb2FpR4LVJTftT6EU9mGS/vwMH
8Ox3Axmsbe3hsErqKy0ctjH659ksIE/5hwNs1G0NYnbEwwRB/SjJRDt/xbs3BmiK
/PnyJ7nPWV2ugKfHP7D9HkXP80XCRNviVW/VIV3geCbxxVwZzyfmn6Djpbc8h9d5
zS9HNr13yCOVLIiHJofJps0TW04o8rasSpBqcJggEhHPlD54wqDUd4e0V4xyh2J3
Lsf0hLlZwfmbP3JSBQxrZLfTKmHOxqKZNbXrperRYG2IYFn4e++0RzXKGBex+Jui
mDiler0k2PMfjtMNdDTVUU2gTbslqVG6rxXUwTj2pKhD/32l2h8h+sUw39QqhOE7
mtI+2j7EAAMKJ20eCQM7mHDgp0PwcCJi258V2WE1G4hlp2xh3E4rjQpioL85K+PM
9hkHgF4XFuzV52yKMFxBzINNh7ZFb1rzetLuhmv9dZ61dUmo5TBK5tP+3xlDHtZT
qPusatDDVuYnIqQ3NqOAYX9V1DSHVPQAsulvOoa2oLXfskRmF2baYLyZasIEURhV
qd3+Y2nJq8jANuNdv+i8Aqh3isavf0gMVCp6a2f61SuKfKhYSjQq0sQZiWoiADlF
g1w5ZFx6KJXYZ2YRpRdkOEL6/hMyFb5zMPZ7PeaoGfRI418RCjp597V8h/WSanGv
SMkb1Q84iP/8MWQIGtohtIYcNvNCruhT+/1QePuy2paBnhOek0lMBHpDn4mY0HnN
PCoWJ1qSHsf1wJwlPmJyob3dk1k9xwAtOXZBka0h/aFFvwST7Jb6HC/K4/HoW0A3
KFX/dIbOYjmyuCJrsaKF/9/W7pJs1sMA6LJB6nJ2oRgrgQaTxNyfa7Y6YzcxPZAN
jchjjUOLbdRNtEOEvXT+NKRJ3gwcIWtnM3RxNOU18eIK1SgoOAbtN4UI+MgEGod8
/UnOHbK/kZFR7Dtw5wscE024/GzL47RSbJRoek1+XkgHWYv4KQ+KGOZqSl2zRYwh
VTvKGfG8tIign5sRQgEBia+jLISJm6i2cOos0DyUgQ+M0QXsNWAk7pNlkXfP9cvR
+zGXaLlJXrbhoPy6o87cMgqCDLtD+1QKi4JUWUYiDrd1NnJl3CcDTgVieOgqTR4q
7Y2iJeMKXA5dUZDNrXMguUF3zVvUKkfsKWJfEkkiL5BmAdkPNNzmySdEf81ZniK3
dVXAYVD10EcNxOuR+Pa5/k55odfS+wt9V9c8eWoqvxXMdQ12WKd+noHKJQEvc56a
JUWTCh8pz1nAf4roUa1Xke0a4TtUVBptNqNe8XGwisCpeZex+oq9LC/WPJxdVSGY
b8vDGX47D//0YDXCoDR3VW6/tePu0CJC3ulgye0hkcHKrDiJ/g9JJj0IdLJZxM4E
4kSuY3XRTHdOsNcuBfyL6bxxFRraCC4/NA1C1qUu4Q2XlnBuGiXCNKGeBG8UIXjJ
SrDZJow4NBOb2dZDrNrglt1tmJaHp+n/xuLNRzv8a5cp8XkyYWLeykJ9hN9NAI9T
gEG4I8iTXB0YwU56Z5Mua4NkBgIPUfOqWwsbUl1nSyq+3hO1ZhkW2MjPjT+Pipex
cOCVW58f0tKPNcMVqwe6GjDbijsbSRzSAWqKIThK2GuYdwQI3qENndu136dfmJij
DPPuXceIgB8VSaEGBKZ/OUZ/d504OM48yBPaXQOgAt6U1HakHr1DlFfBB4VCGgmS
0BiDHW0r53KJx1HOvT//NHapuVJbGL6VKLz4p2D3KCTNHrtz/B9z7PngWfQZFkjP
n+dveUDO5Lkz6MU+Xt/Swjbw8DhgE13A+/oP2pW72lv2c8oGzqYJNxZ44DQleNFj
0oMMFXst/gB1xMFEhidQPoMc03tjmm/cdwwMstHqJkeG7nfNUUE2JNk5FxvgcGuj
CCjs+GM1DbwHuBFM3TRxdeOVkkxZqKun+poKFRqI7fi+q79P5l5Ne1iij98u7KWO
AAQUPSfBYSVFb0na5mdI9lUTN8kYah73iaOV6O5nKfDZiveqtvSqbZtFGY3OozFX
8Z7GeZ7iJRC6H9MXYOzswt6UNzNoV7GV5AcGU+xevggZFfMwIJJW8py+luI/5xCe
IqsNKHH+a32+dEnh7bMaj/JO0m/YYKNm8e46y1r49a/Ugm9b9BszRa31/K4Im27u
SYDCnXsXgqD1xJn4xc5y2uYfOu6cR/l7NM1wADL66vxvWx3vCjiTzw0mfNhY0XgR
2aSiqE5JeJBf+6wRmBPqLhTzVoHfsgr+BhcCn2mLK02AHPA5uuZFhAPcefFCtjhr
Y4j+0WPzoUfQ8e4W771MVrvdQ+PAqdwIUnsU0tI+MiMWRNfumg0nQYrTsLKDaIPU
Wu9jnZ+ix+qWZ88IFJ4EzOa3us91mcnc0rMP1jeUMys9aI27v+v1L5fzj8Q4VOf0
8yNXMjaHA2Ea2Y7xUr36puTcPbGyelVZZMBAL2jrdqDpWPmeEXNbDg7vu03kqKTC
UHxdOePQUPVRE5lpwwR9RQ9LUEijK+MqYf4dIt1BVKTVaOJjwun85v9zA1N3NvJh
Jp1Es0fFFH/eK6Dh0tlrYuERNorwX/+zQQgVXUHLcxqNZzUjfQgG5pCZCGQTyUJA
3NZOGZ0TiHYy62Xighrlyrh08p25a4Cfnbk92v/o6QLhA2sr8nqdIXAgMGts7oi9
dxXVpDTiS6UMxcn12WkaYOKaLKcomA6f1N8KKkzsqe2bomaT+xJ05FcoQju6Ayrs
VPghP2wAJQhyexilF2opACUgfG82gcmjhFAFQGCzMKppHhhOZjFDn3kLXFQaGd7N
JZBcfagnXfhiU5GSDbloro5F4ZmBCWhMadZakE/QBSby+7e2UZVIW+lNe656sR/V
LvA9qUdpZIEDcBmpTrs01hilV/X8COd0kvnzWuJRNvtrPZLLGU9P0xTAZFLltR0E
JCamxXXkUoz6eYsRyxS9cMxXY7m95YEDppKilCCXnWdscj/U6X0Xr9KwHU78jsvc
pTTUfsezfMjY+q1DCpWuAnXoB94cP9jklUXHHifSk165BfP7dRhOCL0h4MViBlCt
ijK+eStgTu4eSzspv4jk+lU2P3LlwA/aI9y2zrMJmzekAoL1x+i96hDvbMwooZ51
AMt1ocOwf0R/L5wIkQTtksNrhLpBP40EiIt+2E1/qzYyzWQmfNGXVDUhDDIHvdmv
4gcW3Z7aIeXrgU/xB5cgwvrnCJSZKpwZacnqGIJbEa/h5XMa+DP6VBdz4rcWmudY
L8Pmi+a+7pcwCZvSkDM4OVbWsO/lyFm/f1/VfiCUCFql7jZnOMgFNydmA1oI4C9M
d+aKrggQyOdiIfhx7mrJXzyK49trNPYZGGJUAUw1mccNPiMCAqi5BmT5DYQQVcMd
y0jVGbiELYLf8oIiDEgDg0M+VFKrpc78GZ9S//NfIdr+xzfnGBCR/xEV9thus22o
IOdeEyFyVGQxuTR+Bxa2Ct2uGvEf9IPIqwy53FXApuFzvprHBO6eSw1JksP1Nm3S
i8SeuEtbuGi+tPlz/Ya/MuJ9Cf4qzG/ANuontIAMm9Hwfg6y9f8rY3lotPC4Z3Xy
xv4SSrvHsJ+n5j1P/oe4o9cWjKyOT/aG46dyRx2Hdkip5IWCXJciC0d2wS5uqCPV
nTgA0yGOMb+JxjgTaIK8wBgEsLXpY+yvEYvya/GfG/laA/LuJSFINVMT3PokO79u
H6Ok6sD6bPWZH6YGXihd1i3XAm79jl0mV6EyVxsab3CRpbaDZBW7Gs9Y8xz0BYdr
LTeQt9lqV1uuEz2VoK89rrIBaP7PnBZ4EzeAsG7iqpxUvm9TqrElLpgLZbeMzH6T
xN0xLBwIUXFQT/Mdw928z+JM98On0eBJgL3Q4lsQJh+Av8Xmkg/VDdvgkWeRhjSf
sIVlPIEDTI17xRUz8Ere2wx9b6OrQj2vmsL5uJJlDytvLS+ZUmHQmlrM7gbw9wul
7pkUYKZfN/LLzLHBrv+PAF7JJtdFSuqiamJJE0P5QYFSJdzpgJ9+eqHKWoJSqeLz
tR7GU73tkcle0wWw1I7Y0TDoHJoKcvn8iRuEzRqx5Lok9VSkEmkfvwoKs5j8t37r
ChNhNT4E+FpV5BSF+fqWFk2LFzAkNtvoF20bHDFlG6wAbnYD0T+RgAnXuwYFL1Qq
a5FxooAKW30Jlk/GBQ5NwFR5Rf+a3W27wFPlKlMELnIha7qLeaX2htexsnLt1HdE
bjfIOsBep5MpGEjQmCPUAOhEaBs5IFCpJSOi9hWXH5LJhEtIDNwwAvKik3CTd+Rr
ZSo/+x+O7MF54WqqFKGX6NsGAjMOwr+zMCveAbDdZ3w3HpotBfUUogetuqPQA4Gd
qC1e4wGiwamwRLFKUbrlWehk3QRFsUEhYZDGP8BevEZX3O9pPAkJmsBrEyA2K7a0
kdBF9ghiaZqWswHbiwnZAuAeRu/BZy1v5t7P5tg1pkf+t4ehtqX3OxBtWRuW8Zul
pOlXbPZUOEhm9+PFgEpfTj97B78QUUQESZtzZ2BvIf2kXuA08YP56IG6xe5K+oKY
h+87dVqgWyXpnPRYw0/J/WhhJVTejtefhFE/IxliH7oTWzDIuDq2FoDb6mJhAQwu
P8b+ZV3SAPJ+TTZNgKCFNBhr9Pr2T0eO+ng/bBK8liTXSJ6nI1iiWty6Hg9X+0P6
v7Zgxaa7FMXiiZeNrJSLfE4vh2MLlgQIp1ySukDQgIiKPIo8DNbImU70tdBeI9F1
pt62s+RAgzklGf9oKjZAa0wCbmnLVFbFck8P0TB0Q2kQuzqSKSwqow9f23eeaKYu
iC+tPKDJqCFDf2VLs+FtC5bQzPShtENe/MwEi/Pz9dgbRlldL0n1ow+3I6/Zhgjt
nsozzujAz7CYVMVQLn4Dhai12XZfEKIFztKuQqBUG5p26/ULoJQdLVe4xKHr8kA3
dXxi8iUlczzIQTj5GWeSZgC8aHKuTO8kezXSDxb1MwOmtETe8x3fcY8Rm7YxMJfa
EHkityNoTPJ6OwcUr110AGL7MdDue47bExvzpuyXlGlhX+jLr/JcwPUWBfKw2mBr
qrWFRVigHLZIkjR/eO43JwD7D4DNR1ntdHIEsPq9VccH7r1HR4oFQaTRi9DazQAE
hYbS28QxLAsOB6bI0XGO3CxkcRz2f9RcZCs6+htSPJXCxO/aoo7RQNavdim5ENfX
Vm6n2raxS30f+GIgsHrJKO7TaCID4Z4JPv6IdrkfxEUCVgs1i5eOOS46rttbbkQ6
6vrQ6MFMNtG9frJfMbs53y9kMVlKgNT4VspnEvzePKWpn11QGK2v54tBg/eadHmV
r7PQdmnNnp9Xsrfw1NpbaZwDAjkyDjM5JiDCFEnuaO8HOucYNlRXcMSb9gLMwoQ4
HUrqczJvz6Nd05PJKQvrV5ILTlYqcFnxGNK2sg4lSNtFhX6s9fMFY9Z4aEaJSLZF
dBDA9Re7MQ4dT8qf6r4D3KTp0VwDsRHx1zXKMJVWUAuntAP6PqSWfYZXC7JphYet
oxjc+g/m/m7sQxP8uTXfFRAVBNQoGX4kV0k8I/FgKhS1lPd8nHuo6v3ZZnM8XVHB
UZt4WXP999PTN3Yz56MzLRz6ckyuat2AGIwhx5K/tNcSjoRGVfZ2dSMfLuDxj73d
+N/QzL+vvsu0EpW9RCkbu8hf4OxomFNvudWxu0wp+wBbx6LVdnYx/TE8lWt+ysQf
1XF7UlGqZcol65tTX+C/mZ0z9jCze8L6zuhLrRv4tE9PaBjwEyb/uAxwsKcnSLEs
zQWYQtBLNOsLXJpbgK5HaIbGHrpr70z0OYaDEIhMvhz1ZkIkrRYPMKG2F7ho8bpj
cK5spSdz+Yk60s7srb4KMCej5UX1FqR2ca3WswRO3WdFK62TAmxi4TPZg05TCMEF
2x0ESQSDJ0fVSYfTCAmqG/w+sgT2AeeLJaZSSQIUpWRiGBShulWQlBTNwYi2Ucbi
EHZqJvLK1J18n3ppQJ89yjq2vlg6k5wGpqmwHHhyGeXj1CjE3qMk2spv0kxPIv5s
TeKqK/Z5CoWGNL38oYllRydS1oUPrE9v4OX2ONzeFoS3WVv4h3uvWH+hziSTKlIm
TvCezj2E8jptykckO1Fzs0JqdZAXf0MDyM/DkpRX52urd8ETx5k2Rxw9XpR1CiMC
Rcow2eVVbzY2UJ5lC6p5wLnsCOwQaH8oebRwaymNgV+Uq0USNq0AyuQ64UInou+i
KSIyexgH9HwXkd4usyk303jCKZ0o5rJzqYaeFkBb3tmxL17Xa6FSEwzVYU4NarGh
gZQ/gF4t2jaFusJe6faR5rhxDPyVZWMojAK6AV/48bmf/JmWRrP8eDMfgZ7QTnme
ymhbvBGThbDfdf0nAMz49rp3dtJUV7+tLzPidJAgZc4wVQJnp9H+FuM40AFOaQxt
Hx1B8T+d5iMwC65MLVKzQKrSbiRPiYREHjCw5T9bv1apSGupS6xVLxdSEOKMmIro
oVBzOcZ99YpjeLqFdqiBFuG/vCBwmTFDI224dPU+j2u7TnD6qCjSDpgnkQj84til
Waufq2syk7hMih++i8a8UcDtit86L6JZiktafFUIyxlGX095wuAJXnGwjTG7G4YU
ROAe4vXFzPYS72MfojJoCIN7KkRHBTRNxzsA6gOkFC12v0nb3rVLLgUY4mCVtJab
vFzed1Qlv/6sY/gFIYOODRrNhf1eGf0mQC+F8N/Rha0LVEqHYhYrZbt1lslexwqc
sh7rd+a5rknu730ffxLSjL7spd04xutNOvictgRRPelkwQdkRmGg0JRwUtL40jjD
AWj+cvEyxg/rzArwucqhQVOgLjV5P1VNvJgu2Edp1+7kAykfAc6WThhOwBecS42L
XOYssG2yuLL0hVplelnQUo3oqygJg4mdGrO8q1L0t/XmKecEpikitR/i6TV8gB22
F+Yt3SYiw0x/WuGmh4BMELBLvvOuFYvDqUYfZ6qE6K0QNlkeo81KT8kOdcKgNF/R
+M+s9TkAyMK990B+noYvuZBwEv2+9vu6j2lB2jX+m0jnZX4fHzxd1Nqev3tgYl01
LlKBtgWhL8LUMtQE4titiaZGQ9TpKowNjARb4/LX5bwT/Cl5+q9nw0REcYTQhtW4
NqcnyN9l9kU8yV+TLllpZWB7sw9LpyYwhcvkltolUufYBExfBM4h8/qik7Slw45D
OTDfM/CXcl/hVeOBYAeD1b/KTwkQyjTM09TH36nFbZk6em3lnMT/mvrRUflPWhZw
On1Dj+5j+5nt/2+qxLNDn9DXixySKjWAr253F+4McldFbiHAkLn09yena4Q9vJ0n
UcWAQxZXz2KYfrYtCWxOgplxysMSGOmvHOBlCJy+v4HKb5X3XgM9s5iVQOCLpDwB
6Vxi1PaophR9QN1Zq+JlJUMSj96dnzUA9fyWyumckQNQz5Z1Ow6pV2N6TnLZmrfC
uowTX0YnJu5x235zd51uNZrQj6+iLS2yblc+D0THvZ++/2ERXHseQpL6ttV1iVj1
bP/6vxsz2ISxlK9mY0OHaH8nEGxqFr87h5gdnJdm7cWkCRHuz5sCmpCw0SI5/5Ja
+xuw9Rv7sInEXOlrD5ToMiJpRg6H2TSRB/fPZrwfHH4UxvboYnZjDabdbDWMF2bh
Ee3g23A8GXOAgfbivSES5enpuG8iw4HDHEV1yLZlFOa/g6l5dthWvB/rj/bnKgsu
Yhi99K+bYLCEZVCTU/so6TXxVYqfiQ2JNqStDZp/5plpeLZFL+Bu/kcvJRJ9Zemx
fFSP8W9DLw2ubWA2HndE4i7y1DrOJ4Ug+H75uNV3l5KK2+zRMNQcNPtVqLHdwoiy
ogplujl9oPJZg+sxTFh9mDwdv9DtxOZSCZuuBkTx4hCk03NM7G+Iter0LpCaqeDZ
TyybyH5uHFB/0s0s8ADwCxzrwkulMkS8thOxHBB77vT11ODf5Ygjoar/4u0FjqLC
7uNLWaNqllj2Lz9056Pxr1LRvIRug28Bwi26rZ8El0TQwWknhMw9BFBLF9cOMUak
bcTcOgRNdJSzu5ObmHcUu/qqEN98/cveGuWWITfGRXyqfKm1y8V3ZFNPhC9UX1mg
orR/GoklKz6iOOfmpZ1MXqy13EDG0ENEKlZRQfv8OO4UIasTprBqPFP9PUJFU/lv
UsxfO5KEnNcDjo8DLeaLvlCv5YCbEkAJEVKAH9bLvF2xaisRXPdWnOVAJ0E1WjJg
j1JtmvVevjmuYpIfQHpo8SxvWaKzAqeXwrqooNL80ytfydmEz4vlvLCBlRB1WjCB
vNR0e004k0zHc4b8w9WeKopx14+1r8wVRvuVP0aq3tTf1XvHS8jzukZwYfCyKcrz
TTeca9M3tPgdQlztrNPGw31idP+Vty6IopI6P1WW9vPKycz8qdXcxcA1wnCDEE2g
DqcA0m7wu95Hx86rZ9ERbGUpEKMs0RPHIGXzH8UEgAE9fu5tAYw/BuQelpGNte/Y
YDBEu7yYJbCtaYsQoMn1LXjgjytkAEAg/p7D/JgGzo6JJEGYTBS6xEO9aTftpJAk
LMRphuMGN9summ2LTNT9OsNHgZ49mhzYG/8yQykch8LxSVsYgzczCkBz51XOu8WB
RJwv8Fudh4hYCzYpJu77m7d5Lkyh00JbpfMRmj+pp6s0TiD93mvCkIt8qzRCWxHa
hRCe/QUndVXxcDhyUDerzHnv6FWAUsd+G4DMyFZs0OIlh0zA+cdA63N8XMAfU+7C
rOuDu5nVdS2V5RfFhLvJd8+LAkR5LkN6M7DidHaHPvqFboaEubw1mL6CS9W1TIEy
IeHQlW3dUguWUHfMFpP8CH9o44rJ1HpJc+eM1RyXHOCdXOLRfhTQi69l1PNVAwIO
ro7TSIjDlHMrqXUkISDznO5cptvR3tPJGqmkW07EQt5nCZXEkniU56TONwqCQQTN
kmCRg1kCAMoHCDPzMJovGTltzDy7tsiFXFt4rQcOUQc/pGHO47zp3pqlVBYlt2Ej
HKnfSG3lphyKVLx+CnOgpDoe9LMXjsPbe58DqVNUF/CVtufqfCwbClmCaQwjo7F5
cg2x81qQPgCS3wi0u2LT/Z+jOj0Up4rZoiODYUDxe6uPMEoK5AvLtCQfXVMVumIQ
pVGnNABWGA0Ph74j9F/liUYEpF+Dh5IE3kgUPytuSxj0hpaG9P5U4mxEjXWnZ002
AUoeW0qT4gsT0t+ktBN4erwBOdMt1FS1FX4ycOhP1IEJZz4v/uSZqPuhvStv5c/B
joqc/9e0v49Ks0ZVaFoky4UycG4QhC8nkylTKByF288mCu82LoAQGzNmu2ujJd+J
2hYFGoiDZSEeRoMkGmNC0xLcKc8cB9+C+JsW5Btulb4HDdMCgwLUGXQoHfTHH6kD
YrL7khVGJVasqLfZS2pJCLG1+l3ihzUtsATo4msErCiMrwbKOMtXLN66vFeylmRk
ZM3gFhPgybhC8WP8GxMvmk4tAkQqzXVgmO+eWiHKFRzKVs+GFh2JjmGA0K3SulJB
1kNg35OoHgEkPoxwNOI5EmhmQ+FB8auShrXLBOlDItKjjBaJTLYL76cOSo/hJrv4
hTbYkyxWxHYBXdCIu5uzUpe1D/NZ2GdzB/RWg+JzScWxQamfwtxrbEYUtfw8F3p/
SOgld6xSNbGSAebM1Cc2lG1oJ32Qn2yn7ebOUQVZJwkFT1XbqZnWxku3AsW84vVn
NCFRGhEPj6SsEyvy7J0jVl05vrjtDBsGdC5HXj9hiTsYpusoHOaU/D0dyrONg8A3
vuekAgVZOAZ7TxvMT1Qd4Dt4b62oTRCs16PfLkbxntI2hNwwrd7R4xLDqeZkQVOy
uaG5IygTIOLAsfmEMuQgentNBc8WhmeBd71bWyQPbXRZS/orFzHZjPKAAVBaH1D4
k1jE83MYymUuSXZ2E1nVfGhZoP4IJuYGR110RQwTfpj6M+6A+6Ir5H14ToeB1wrY
4SdHXAzhrR1BxXzAPT1yOLrr7ooTJjloq2r/zu8e/BEDOpRns0ry5b5XdSYvGzwG
VM8LxhLmqQ3AXYG43NYMij9aOssikpp4oFqhR51usXs+CC6u4gv8N8de5hNp+5ld
sUE9+Eyeq0gBexERSQjBJBHegPDc5Tp2nYodzGlPoliOTABcenzy2zpGq/fTsZM/
uFeCbf53BbZsBCLhDDTOAekTMm8OX3Qp/MdN0DE4cp2DGM+wrTt83TsXG5jdJ145
vsQHjtjjiTNMjt0uU7tr4sPSLcD5CM6PWBCGiLZFCMIjo8gWJW0FugZT/E4ToL0c
Aoqt/IWt7FhMmOOAZalzdWRR7ElhgqS3wAD6J20W6Nz8rbhB8613myo9IRgHbiMQ
N9ZUi6NXa97txrXMKcDQFd+3eV6GPaQfIDZFsQ6pmH/VXbGD04fjBdrwcqCvEoft
HNuZfM3QqywUp9sTTfkkFmGb+PO3EsXQdDt/J28k5pnzdgZaKSSLJbe1KT+rsWcN
hyT6h1Em75wad91iZIc7pwRqwttXGc3nZbxT5hGlTHbb279/ukaFiHZsANLvjqPs
bkeE6f4Y0OL9OqlxmOwbpXUoyGSKB/gwV3ybe3wVa+mRx3zZ9I4TS/TZpy3ofP1O
6OPdFwVRZpSQcecg10OoEuNNfVEoz8mVKdx1gZ2H5aj8nHG4fgq4udDAG9gDvCh5
WlLfSlD/K0P0qzP0ioM46iBFrPFhS0NmRnQUk+wX5FkbeQDRz8OmkVbzpdJ1XGWw
mz/Dwf6CeTHlzOov3bWplXFIdMMwg8uP/xeKTqJPxcStdBU0OpiAwkksPBAoTdhI
jDiO086FqTZ+YJQRiAPZQCXH9ixdxZErL1OAf5LtTM4yLMxO5aEv6l1pViPYufxY
T9sbzw1yPy9SQPxDgr6A7ycyCTmyMNBTiAoeROm58qtXN3jg0FutCmuD59rglzog
nsyy4EQDaT3m8H22e3X4Vd8/uF0JvqHBIlk61HOEfB8eCoo9nFihFI4IpzlHnugV
R9UxV6akpgKtQR9daSsyE5M+i0lu+tS90L8q7XLJpLlC//JnapIdaWeTJcAcwL+E
Nb5Gkj+xwYeN/66IiGWDp6SXEElJm2XWe94aBiuridcL7uTsDV0xybJLxaSR1/On
D33lX7id7i5liEwkcBEf8SAAfARqpbW6+9s5FLYY00Pg0S204N9IZ2M8GsErttuW
wIzr8CaKdyfmAV4cm4SW3EbfGBm6Y0sEN+gYX12m9eTU9hZNaF2Eoy5iuQT8cVAB
uAQrodgpe/fZm1gP4tfStvR7/AQcnObdYa5rQ0KtQBL9YI/wYAZ1J5AQm2FixOaI
wwDcEg6MqPxTETeRLsexyMi+SLheYOlPHkQrceqkEHvF9Cy3KWfXidjrALPH5C4Y
Sl9VRc0/4lMQ7oMSQUNeXYOerYqgx6jXeWP0A4j4/jYDALuOGq1F+fp+/eBiLMAz
KZUd5D8DuMFE/cii95lq3hHZ2/bkmMfPYHSb9PkhkAfxYVQAr+zwN8WrV7ewYAw9
rxq0jWjz0K8/VH0zuoG55/lHdKuId4/S2UPY2lLZvq8t+OabH/uuoko7ntF1atDX
2gZvbYju9IHE5+Tmc5iVuCvCjNlZIx3GfQwxLjgf0mkSS15gzCJhX8ZeTW6l4ObP
tC05fAoV2hQ6mo+t4Z3rVcMADg6s5OI3NhvbyywJmXwPpELIb8yTsoHsm4QaYo+e
5BlCSqCznHvEUC4ZKTkyAtmdRv3/+xcuDR0CdWhyw7vb2/06yNiN+toJMNyN1iMO
y8Iq0tB3ZE/ZCH/VzdXF0tLmxJztEymdLegJt8yULSOTa29A5SgkUdlWiuOxKpFd
XtHZ0XA2iOsIG0/pUmlRpephFoLMYbjwBo2aKvalKLzPunA1/4Q6FBBkpSEOstRL
Z6YPUmn3318/kLmbHvGDaxUm3NL+1YFFnQL6vHlKpVMpUW4V1DcYavvrUHY3eAwu
0QUCX6HgrnysUNWSnLoceKJcDS0NxwSxfHUX1DJCqmOLzAkjiAyDuDWhwe0wgpLK
M9aCDg1Nl9PZCYyMHlgsbD1F3mnRx6eoFX8VPQNzjLDyG91j2UI9q03HKfjsoOEn
VuyajXEG3j+lGDDlAgdeWd7fRFC6je1JrJrlaqHnNiCaIzAPYwNA8UYg+bcYS47h
Ot373VEXOFz1fQtIHj7FNZiwY35U879LlhO+yWIBQ7buPVxZdc56zc7pEsB0nvjL
wfrmGynxuMka+lFZp2IY6X6JipdOC2GYWvIaUpGesKwF/39Or8HSAbrgaCF48VkT
6Jd9BZcF8DxJ/Ajj1VFlainiegcPfZZqqUuBOYOp1f7R9hCH1NhoEzHXeGmZdVg0
CYp4CWjxFXxj4pKev39eCWxzBHUTmf78XJ+VsyKBzvBzPYq3M3uTqDt9ZazyGoiU
6QPmwtEjrOGQ9QPIV0eMidc9Sos/62hfIJo3kaJmpk5KoebBS0BzwIDI7tQC4fNQ
ThPz2a3uJM+xX40jCnBzkoJdmW6nRPPqgrpr1AgikeFdmqTyC2T+1EHN77eU5scI
9hvGFHj3CjqgmxAlqFJwH3hsoo+Alhm/Now4Cc0+zV1cDojzTnyq/E4KrAiDuFkc
2FPEBDzFYpp7V9XXL124ADxuhLIsQODT49JoBLGyfK0VS5VFha0RVVNY4+YKnmhs
Zd0Vq9+VRgzgs368RiMBOQ199aViv7LPoCTv68lPlgrIIrfl51/e/TtalEMih6RX
Djj16qQzfWpySRqs6R+89TIl1LKXGmbON12HFa/V7Il3U40F+p3x7h0Fw8Q/agyF
u9Kz0tuTdHu/M+bJAyEkAl5mYGDw7nLiGS0veatgeGINMMioI4fRdY9d0U542cuq
7HzNoeB1xUx5KkGf+IBT8U7MtoBMdMh8OvHbkofJWnTdLZwHllIP3Ao9fHd1nVMu
oHO3lj/pFMmzN5p/lZs393strP2iRKw3qQf3wMY1N4h2JwND/F4M9+PFaZCIjNyz
bfr7BRTZ0cqrwgV490yEQo5e3watIjeVFfru3iJWJaeWxoOTXzhO1MV0PF1t9JnA
RdkJYFM02Wx9dXJn3AkT51ORHSSOk4Wwj/MwdomhCaeQ4fXlnTPn9YbD+gR6Tfxy
jQ0UMMnRidy3rsOJN02vlWVOCEa6EFi8S+xKuJ6v/BRFb94upfInnQlC9m1tWXzC
kaN8x4/0Zul67S5N4LBwZ+HhOCikMdBr02r4dR34izjtgEiXB57FvxeWYULPCqBL
P0ICWIQHWIsNLhK7iFkCTrThsSk8nWx1Wr3o77OED4vZf00D9WvfhmTcmZHrDx4M
vyEC6YKKnOGFNPrrzm9AP5yEAUH0JApAVEXRwg1ySh1BCQagjg4okDBIm1Mnw0MH
GHsMCmq5clMwuc02LDLSz8Ki8WKhNLHOQo3/m5l1igzvn3df/88j09rNe6uFc7ib
uzM7Ptu2IFrUNVQK3tQue7hCwBrSZJz5yapPCGLHiPaos91+VVxlAOgioXsOxTNb
E/HQDYezw/xHiHomST9QZR4+ovw5OkkdV+q2upFKHanz41MnaWvTTcX4VbCNpCMc
cvIVA3mQG0P0cPhX/lep4i6KNHM57WoG1ELwJ2uHKAHTP4m8KVJskUg3PA4ypQef
RKHn0AWcekSXjypy2T5LdUsG79XY5RY5J5F/q8Df9qSPckdDIa5+Zt6XOtpQ4/iz
nCFqkBTSbvpzObuCspUXbkHAI7igrt3cNJSUKR0mH+uSj3NNACftHz4D0h8ctMxm
VLUIUIRWRuw/TQcnNQlg+FYtpip2+vB+A2ZOpW/1PYVXiZG+IVw8iyg6sHWcHMNX
0QLcqjtcb+mWP7L1jXIFAWfWY7kZJagWv7V75hzIslNObGwzfmH0Xph4kwHrBeXA
dmqMcpJKd5sG2FH7b327ncXsvODseaJS80UdzkBdMV6VGWMY3mr7m2qDZDI2wxbi
2PRSvjzgj1E0NK6pF3fdvS3xs4Dr1LjZmrVeSoSICv2ZCo3x8v4/mRSCvFP2ymd7
Jl6F7I0mxviEBKO6fo8QV6CVUQMTO0fvdFmnuXAYS6+Z9K/zC29G68NoPtVTB3eA
BVGZ8uye4iWCAZeJmtbNQcQaGpKMGGtWSeNbhQY3LagGEwr8nMCh3UT+05Ezl9xW
Bh5VnP6lepFi/orD8mgtb60hpwN3a3QyRCwXDqCHB9nuFqqs3HILYGn8wcMbJh/8
EVDCU9F6qFWyuFjGDhTNAYoiaFAJWXwn8fNNlXqtxrGivPM4Vhez+5uV0h/6QgY1
/cqa5QVdT0SDU+04vi6bnG4jqA3uuoqSkcG/vF5HwGVYyiky4Owqjy17P8PXYE9Y
nPffGamT7SyQBJpkVObOQMnqu7duRzEN9YZqilIowgGgfcEXpOSIul1ojHqqODN4
ce2OcJiv/dm+jK0U8MwMeA0ifom9X34DQk8M5bFVdgIfam/UGMS+aE2Hw/tKE0v1
RIxIci/CYwT8Nf8f0lEx70DxJpAdcaiCX/bLzSP/ul6Bn0N2pd9eDyar6yd90e5+
h/WwwYi9FU/wmdwohUaCrQT0KBFMyCgZfxl4wrqi9RMC15p5F9CVKAbXoSVRqu0G
ckR0C9VIRQNQuuBiPvvc4pmLyriKYqlOM+GnX04nOnN5CGmVdhM8qWH9lIijT+lT
1q8z9aZ8SY3Vd7JSe5XuDxfUZeTZHnC71tSudYzDmlCn9qoqq0bhLELCuqMxQhpP
qQl9Lee6bPLmxFoLnMwmkOYv6bFELptCTWKiroQmcOROTeTtVyXJNSf4dRokwMyE
wuH9IpbkQYCjf1q03B1rl7lyY6sFainEouBCMyYhWTcvLnauL7Fdo81JR2PDig4m
NGJiHvD2RqXUq3xZ0EZhboAvKQxZqqeJ0kq8+q1k3vg6VRt+y/ZKEGiSp0FjxWRA
8xZdBWh64QuSaBqWLN/9aKj3jRum8vKr1tJcyPk/+juGgaUhKNzdRD6MWIzLgtoO
IzPBQukN+C9rL2gkbuArtMRHJgz8tsDrA7bBuxHGwgRWCsBRl6ouncI01mFr6qyX
lXijcx22v0xIaR/QTGDAutrh799THpgIcIaYle3y2QCN2PcPR9y2Y7WN315LJ6pW
/6F+C4s1gw1D3uxawMpGKaLzD5eAtmQAbD6nbUpIYyqwwwXyy4ALIFEcTbKTFpJp
pI6MuD+mhQN754LxIVTqMcpyEpGjlUAk3MBOwuHM75Gh8RilaqUGTjBWw5IG0Mja
nv9eb3RpUpGjJdzRAEvLQyKVQE6RGMWj1STXo/8CTlWSGQIbALFZUshJKXZjwF12
QgidttyHrAx+OaYnz/q/7PVDunhrRzKO/U8ae9nKUstJV9B5Tl460os+GVAEuAOI
esYgfYGJqgQNLRRAdWjfoBEvCz2aRd5t94nxUtvHnUtTFh24rU6YF8cXpwE8pFKe
Utv0E7rZuxor9C09E8L5eKJEF8veXSguRaqFRqvOqEyXDbGyUjvcRha5sxo5HCxr
dcIwQexCVCw01pf4/JJu8k1lNe5Fzdrcf8TImTW573XFbyJohuH4JhVp1Ptzke4+
da5mqXAdpKEzVg14fY6M9Qoc1wVlCetKnMmnmxKc7iy58aqyuG8ovt18fC5KZ4sc
GvagZEHxQUb058yBpES8t6zhj4VYNDx6/ANhd2HFs/rOyT30LG5CMGmTG3/A+PSl
vbSW5uzk26oY+9a56kQoiJyz5LSMBEK6xOZpNnI+SBZU/NX+Xp1qG/Q42siT8i0O
QRnIKlepS1kBukkta16yFzNgnTOCqYua4XaXvXQlM2GWFAuFlWxI86CLKQVT3m7/
PjfMxMaefX28c7sty6+fwACbhiEJbNsBCxQQgnGvpNhexHcRGFGFKY+pEXNu+nn1
50vDdCoLg5EdIgS1KMg+4DVLbsUM1G5A5im6i7Unp8fGwMRS9Y+sUloJfX9Km2Hb
ht1mHDKI2X9aXL3anEBJio4RMXN1nVQFhpibRylW+UpFhFuYcVNZqgeB5IIt5ZpX
5CLkQ/1q4Bo40yw2lgJkqic48/2TwO/bZRPKFsZ0VeBbh/31S6amLHUIdNDhHTAT
EWUjbE4tsPoERvZTTxNR2fkaCo140mT2OkikuIv7powDUnOnegy74oex9D6+rsu1
kjT/fiesEtgDb2UUhfwYwwcPffWIf7KgIce7TTBsMd5cRbg1PqGn+tZ3jBkFEOwM
3xtkJI8idPlZF87Peqt9BcltVtIMVbs+QsmUpq6utbnrnESKyKsEVJT7cA3l6av+
2gnQ5h0y+Sr/yroepqvEFo/Sravqv9VmE2XyDSE5YncBsEGpufjWG3Jsw+3FfZyP
t2/9jkvdf4vB/9E+jorWW2THdcsCOI0sAPK0b8sRoTy6OZiCvYLNm5w0pERcUdFn
tbyMvQoML9uwWA/yRAvYjavvvNwG+ZJ6kgLrJA0eD/JZkidp5USmoK3vUThyRIxI
SOvKlM3k0h51eia8bBYNBN+DYpU9CUxrDB9LPaA76jDmyezSo7MrY+uY2QJk/gsk
y/Ha2vXL06VpMiYBTyz7l0FZODQgnTHLvIQ+MFlfZANNxYhnzdNYjhfNiWpJQnKy
LBTZZOWBw7b3BAX27le4f968ZbNvrSvvxQZ/13TDJ40fH1ui1hH73Iqqc7oC44Vm
gVdEcV8DLnMYKOg71nnRCcPz8x0ApOOCoXLEy5CI/MUkdlZI5DPu8Vf97hgpowNe
adKOh4LnRidi4HQHo86ZfUOllArpoPTdtRHrRCsO5LyW0Tx0I8ITGEZqKlMQjXId
YEZ+kET183Q1HcPOasIVu7IYKUk/XQDarHM2SMNMKQwDKm42XW0z1VfKaz0GK1fx
WHxu6ghU0nlcShGoJaQRUKwQ7hLSZ33NrGvGN+IdXGuavTf9r3HZl+eqBRe30qP2
z0Jb8L65WKVYVqieU1FRitsA8oRzX6StxUKRxb2eucWm6AlQh/tqCfVIBvciSsS0
tnmYtuohsV7VVLFMVxZ0veg95mCl1JxSuLwa0Oo43hfyN23X/2iLdglgLmtDX2Fm
W9xlJhArJ0sTzrcT36N9gt8/5t+Rk+Q7EJ0yH16n4UWcPZ+ioZ4WzgQeAmmQhYaP
3gozQUIcr9FlxFwDaRMkzVdZI6H6UzWdcl3OfPB90I24zayug/qp0zjTMxIk99kk
+vVsgdA2JZ1XG/ubw/6ZvEXB86zlSHHrb6ZUodbBql7tKbTPGPqQ4990XA9VQIQ+
N3tZBNzkh/slqzQ7srpK6GOhNrD6rjAY/WW/CAW7JFMafUb/i4xmtOhmxnCTdzsD
DHtFSV7tExu2rQ0/13NgDII8IoyRBFA7Pxix2TfKfnH/dgooCpu6LVFg5wTbE9OX
wPTBhECeU8qXpAIDT4pl8DmeQB2WSidhLkwH8cr16NpfrOnYudhs1/LJ8fUN/E99
t/Kb6NqjSTbY0KqJ6uXiwJRY7fEptUmktmvMktYHAe2nBTkHMpOyvgzdgXX/2BYY
tV8q/I/NUCTeEuTWvPPbXGZWkGBokeikBZ4FK4OW1ReRFLikXX0bwpOceNwRzOFl
sPp+veABp8T5th8sPQaXh9vRkxbXjehbhEdS7dINH3wsDL3omfmQrcYgT4HIxmDy
RWFtTNUmwhLMRFltyXdbZmblLoeWSLt59s9ar6d/O1yDALUlsHKlCzQvULSxaBT2
HvJpaQ7Jz/UGZ6s9WQc3nkRsETqOBHLi1CidnHfHEHgMuADTx7SejrnIMDSlwAme
yM7sqvmVH5Kk81Fwknw5KMhxk/2KqkCXjxGfBucVFs5Cd1DWQ4OMf6uyYwqWvdCs
g6EIHuX9a+oA0u/nD6j/AMCXYoi77CeGop61UfGmZEB6HnGiuoC3sbT7FoSBWeDr
6UXEgvDOH7Q5ijzVNRNJ7KKGSGaqBQ92VgL7l5hR/DWRfMaV8t2Vc9uJfNKchz23
hIbcIDSKnpv0gIsTokTJLvwnP5kq/aMladobN2ID+QQYU49Cs84eJd6CvM6Pg6+F
rRDohv6yTKxwtACHjAwrBYejfYBqlgTKU2RS1qoYDvMW3QE4/8J4ts4xqJiTX0m1
8BBh13vL/2S1nGrd/kXhbKnQADyVhMQZ6FE5Zp5z9LX7G42WtZh0ZHvNcuoi/hfZ
NFzTIGEGooVwSdnwm3SmkY+gvM955WTGGkj/sxUp3AhKLvDORmkK/Gofp/jPaCld
MlL30VawXRpQ+ksaOolFhSCPLNdmHKaU9QI8LKEyYQepci3y2JBYbnZYZnjMsfPU
0KmGmbuwGhF0dSuviYMHPJS6yBfFho6dqjaC4LX0R0DC/lVd5D8yln2BcxJZVxEY
sivTA/zyqRmOaS6uyTxF/woaw/PByKYIdwUXL+3GNv/z7iB8XtyU2NKM1ag32mWz
t7qPUcwWQbtyA6U+l1EcftFJ2hl9HCyZH4hyrtK65fUl18krUFBfxZEm3SwiusjY
NzrjJnVgXSXfVeRkmC5ZIknsHivcJH6+ZpufxcYNBkYUVlbeUNonhLPzY2zWAR4H
0vhQ2Vst+VBXv8gKqpk8/C20xfUFySRFYyatWRQKi2mYwyckonXmrqFLR1t6DB1k
26yJVGHs3j7Ir5F8yV4HLQp+KWOssR2zS/AUmGAAIdRfZRD8ixF1eKp0yPrFdIS7
Wrw1qphkzM832gZGtvKT93btYEUqeR92cAhs/aBmyVTv7j1nGejdx/zuDLagPgA6
SWQjfYFO+Psj5p0RdWpsLOMIzEXt0RaDvnXLL/q7SQEakqcn4Kuu/eByPRcdgTWv
sDX50XOFiQMbBvfd/xD+GV167ompEyBagqsdRxLl0vme6FlOGe7OagBMifJX7exB
T2jfIyS5h6DqJJSca3qTylrAuQ9G+dXh1yYI4ZjS7UTtXSf0gvmw+h+l2N3eENC3
q01CDzvMarV0V6p7WT8NTEyxYnuOqxeJ0qsqVQkNLqwiJYEfknjJ0BPLYOlt2tNw
nSJzZKQlv7qHW7R406uwmfcF+kVzS0ujCl4VKidh/AbguSsm/mbzbsgMMLgQqFnO
hLgKIAOIcNEjo4JELdSK0YiROJwm1HJjdpxxxEAIJkNpoawz2iGFJU84t7zKgyIP
SsllkH2x8dF2g2hUeKLr2d30zvNxVGFwwEgm/hsLSL87TpeD9yuDWD3nRcM0oHC6
ISzsdZaU+rZGaqCp4Peg7F0UoOSnDA6p7MfFMEZXx1LK+gcZXJYfms2Mol8OWy3M
2dZA9Zt4c/SWyQxpJ2dS8UyRmjRfgxLfoUtY2142eWFFR7VGQqMYxdL0OiN3CtQD
30kKHNNIfIYT8noizLCsVkQS28f+FAi3jvo7svKJgVg/nX6oDAcKUGoH0FzTfcG8
fntUr6jiPRJnF5e6/d7tiwdxgfMg94zJ+tJX7B9DFxYnnjTzgUS45f8xYCHfhXMt
QapyNm7rArTHESebB5NhCG+vMgzpCn7X32qCDY2pNzpSs0hoNq4mJ4jOyf5g8Ppu
AJct3bML52ss2Y0L43iXXLT0EvqKvOxWShHC6af9iEoSClBl5Lqy3xz3nScSu4RM
oOMhjuLcg+eDoc+a6RC4c2XsEvWtK3x+BoBoJ5PBCnFX+cF6leFQ9yjx2ePAAxmS
8dRSIDgYBlwlEpaJrXZa4GnCkWjoY5qqLYAB9iCkUlvqDKKhvRxXgZvPOMOJSJEQ
Iy9lZ0P2Iq5X1+0t8dfJfY+dUULXgXa/HKkm0aATNX9mVCusZI8+zTCeRjk6MujE
TpcWZt8hvC81tO/jeKzoIYMh8PYhfU0S6dOPkA5lvDQs1k2aRQF3nlEQxRjYn600
rCoaqRsALHbasqc1j/ZjZ1jbNjXv4x66YPDNwUjOPKKcNza9N1zSr1K5TfhZJb9U
hFWdQKTJEY+KK+zVReb++lWB2yFNrwUEtCHaTP4JrOftk7kI+rGfyS/wwBWbchZu
lnJsoblHPziVbpY/nwfSkjgqNUTMQjBVqgkpXACzBbTrrvsxXLOQW8BhxVyfkngN
A8z0j4HcZi6A0APAeZYV0IcjM2STje8iZwtp+V9m61WkjEKrilfDJWwQu3CoeiDZ
7F+cyZ+xc353jv0VpBUUKq7c9Sk0zGDTYrTVwtBsHoC9QrF3ouJhFK+s6qHoga/A
lZSTIekxlmgW+xhJkEOXhPXJqJS6N54CEEcEiCkfbIGJbn4Vev2HDKCOpcr9l5ox
wbdS3A5nlpoclo1Ppngs/PBkIkW7Xx6igiEd6V+tDC6ch2CwZGyTYER5xBhlj8Wz
zyR8FcMw9hShbV+XRA0D2G98+d6Zq6+85JsLBD3DVW62kExRaYHWKk+P82117udU
zqw5hrWaba5tYEmzBF5WNaUkL6T0NsBqRlEGdz+k3kb2BjIQY49JyCQ/wYa8dCJg
1Pevj4o0xmmMv2iOxUgnCDWH8JxxE8Mu8ATZC+/p9HRWCN3w9rgVuiQXyPd8divt
lhbZObS1frosYQoqfpwAmt0iHLEXIXPxwxZobpWm6W+yJo6FWv3edHeZnENj/Cea
Ty9ODy56YwowgJWJvUtejmgoKpxdi1Rtv+u+ORMMHRPooDG5w42b7qGnIMyWSmAJ
kYEIhBarSdhvKb6NTUH/sraav2s4cuDKvCm3nWwjcOy4jn4PzOFr2WiFjby0ICIo
903RcBPUnGHwpGrqEP5hI9dZrtZNb9RH632DsymZktEV137bpkYR/KncOs2cHpaI
B+Ik7vdk4PsyS+SMRoGbwNjQ15YqynRIGc7fGJapKLk4UU9zJeojtTrpXmi5028i
Jtrjgq5jhk730SqESuZC8mNfPWvnJx3Z5V8HGqIDpgoLWY4OA7jTH/EMyamS3uf0
YRZB9+HMyGsHR5tK7iJML9/qG2atUUOap+TnkRYJHUughYRT9ig/xdZMOwoiiAxv
y2uqIJiKZlQjyewASnoUNObcKnFqJaflVoUP2lL+nrNvx9+10upK6QGgvQvub19J
cQ8wpj8xm5wxcqxK0f3DE97TiuB1C/xMm5/FjQE5YVqCg61gnIh5A1PBmg8fDznk
Oni3BSQFXaIgk3ShixJfkDSf48NgHJkrYFZsXZrnAZTWDMTErxcV8fGkETWV2k0s
IZM7J6p5pPvBvfILaOVj11md8RNAs1Z1uO5NrT/O2a7gkxz4m3PSprPcOgkOAEeQ
1Iu4u0+yT5+PgkXG/YpSwse8UxMKX3kLb6xGlwtNyIDUR+lrdlnZdeSRA3fkmmZj
4ZPTPAsJtqPFn+cr30bNpbhaesN2tiVrifw8wUFNbzNmI2wvECYlZun5JZ1EGNFZ
wC0RNQs/+hRgtogg0TG9u31UwmtCD6rEpxP5XuRAji8eGo5/enMpXH8MzBBshS/2
gP9q6Xqs+tn9rWLZLHZowPEvjU+CzB8GeM3AlkO20YKHy65ON2az7HRg3FdrufWn
vIxlb7CZ3jC1YRX6BA91603UltjzaVvhdwbT5L8UiwmwHjmcOEanJN7EPCHOkA0F
JeVZvHRkgSmqO0uC1gmXRewWoUjKqq5Qw8Lkp3SZtclKGZKLY60JcgrQFOWVM+tC
rmoLACcwyqtPGaHFmKQiM6A6twVNx2nIUOrJB6JroAF2xH02AHqvJqZDkrhxWMRU
Km76fOyNGfYvtp/yCCNcd70TRieqmcvwkqdtWINXg6OJu7e0XSexHMib9kjH69gO
wu/qjrX12FiEW1P3y5SBoNDOsd/6f0DfxAhtlZvMDnvSHnQEjJGGkdopFA/kO3jJ
HVMdLyHdhdwgL7/64Zejo+8pOCFzhdeyNWRECWOkicCOeVf3lj5lHpiMzwL7KRKC
jbKRvChbj+1MjOkz1uQeEIREvOTIwiZVLrXl9a9Dfxu516NzH6tHJHWxNmRLubD5
mImGRwh9BJKhgfzdjFbuUHR3ARkckgdkv3IgZXHFNlU/fOShbnHvevKGin9/bDWM
pOWPwW2FH+NL2mRP+GVmZ3RWRGwxxHoK3XtiZBDBidp9PgWx46GwbqBisHhj4aRZ
hFvOxy6wrdPKxUWX6QfkeP4QqR9+GYkWx1jCvnDufEy9t6IY85VECeQzw4JlARny
CGk9j7rINZTOWpp6WY5RapJ1bUmCj40f4G4WZ9mPdPPzRkCOh+Gn+C/m5GiNXyGY
GIVoLQBmL4I3daFlDchiG43V/vA0xLA1UwU+q8o2GDkBnAdLmnpAPRCBojhbvU5X
R/BsZ966gAM9rpqE+RrzHNePWQL83+y++CgdDhJFwgr/HdB6ZkWvlLohHMDpI0fp
w2+GS3d19zIsdGZUPByPTppxj00s8YlhUZYgsXPVl2njwn6OC9bSo7+/IijQkujy
KTEjBNAG7LUS/5vXMiyyeCvUPYB6MUGn1G/FsmCBTIEyG++38EvuPlCbIZqg90Yv
MO4ARNIx6Om3HUPVfwX+PyLEkCzCCBF6MgC8aeHSGvu77Uwe3xKJSImfIvLLB6XU
oBPRRdI2GFfSwDl+VQePB9vNr8Wkjom7S/3Tb9yrsbp3a6QVVo9yqGikLf9fWjhZ
khgwoG7UmJyT2C2bVJ+9HJaeYIszCssuvpgH5QMShIui71KAWduP6Nx/m1rUEgaw
ihrpcVOe6CtFhH9PV2Pttpeu7vQoM0cv6msGInFWflZwzq9lBFIK1oTSEE/IQrR5
9+/hEicUZil7PFAOdCRjZFPDYBm1CrQseoBA0qgHiGvnXNv//oSSdqKHN8sMnQS0
MCe59rKY5eFu175c7GU/4byN7dGQ1F4IZ5nW1D/5BfoVwNJPl9P2FTuHFWHJXXFz
Sn/AWXy0zf8b/Cjnhx67FN4BAXhMFWYOvZQbkzymPzfrVPW06r6Fzgu7MRbjVhj2
g0bGckLqUr7/c2L6B7WZko5FwAcMFd9zRzo4KSdxhD/L9a3/g64tbZZfjBbeIjCD
1yuBTHRxWJLgh52dw89916K0tue4KzqWtz5WIcZmugkvj3RcLZUmGWi3dZSigo1z
8izT3towynP2w7w66pCm/jAf4vdqlxkhhYvAtfAPYdoSr9MNxVf2SiYMjjGBPOzW
wJeu32jZrfeL+TXwMk3UcN6Sjp2/ofxEVVE8MsyQLK9EYau5X0Ctf0smd65bO4NC
WWaJ8InIcEhWpWyw/iCTpFmR1Pw/hWufTbjFrouVJ9SA7oIu1h2KK+U95O2c3Yrb
MfcRas40HiS604Sri4Xk/xNnUxXiJ+nokHF33F/U3ac17Ifox9jtcDt7yg0dQa5c
O0JlFdnc/I4KwI1afq3EjtWTT2XvSeHo8uVi0efCcjJG342yUULjTH6MtH+5bIal
CKtml8ikmKnztNDAaR4evcyE/oYEpfz/8XYFAYeYYUBuD2QBcVWXFiwjJx/AZiCE
71kGkGK7VdQ1qOhH478M6Yhkkzt67cMn78X4uQBW/rBv15uPyaGJd+fv1WFBDOV/
c21EHaaEHpq/2qWDObIZ5CnkYlyd62tBw5sQrPLDR9RwyJYLZGGnY5i/We1lr+Cu
cL0O2LvT7I/ZgkGkHf5ddWv0widOzzBSB4irraNIbOJ0f29aoNDXI79B+HTyJOes
UQqLIndrjOYo7dHz3MNHWWFKve5z4u/H4/fNTxtp63QCTBtPa8RM5zrsF0sxvOdF
/f9QJWnTTqM3i1Y3Y4RYDUdFPaSA515TX41EfItN6q8oGgKdXE/Y7WuHFbq8gBsT
aKweLAl7cM+1WJpzNP9eEm4vTVYkP2hVgD8RxeDuc0b7XyHnJ81HkgpwUWd4HRqX
hXzzzkqiKQqNuIWH3G7QC+gkYhNivfVgMr2jqFESWHdeH//jS783g59uyGQG2OZy
rbCgs5zZiQW0p4kIfSgCovRL6n4miHVoaaw3Uv+YJrR1m781/xSb8yyHWQ/J65Fp
gI3xFz9U+OjDsXvvPsOUaGzgZsLD6DzxwBy+6okeL6Fb9pkGerAgLPVZhd/3+lXE
tEZhFCGJJVY1ob/IqDtg7re5O8nRlMUSuXfxLXneWWYT00GXkdwya9pEv+RpTxYS
1Qac4eeWY0wHPGm7IfufCTwyQVw8nRGgAfBS2IAbLQ1irpmWM3Ra9/zvHGPowzFX
ZuY/ASc6+fu7fNTx55PSUQyyCnbX3TA+SCofAPpDnGHRnN+utftHUYWayuTq8Cl/
8SebEwrYLFqBPxBx4LOarV1oy/Dfcmsl5aqgbTD+tkoDY+wbZxRPN2MqD/WZicdX
thoV5i9sE3HTsQDgfK1quMXeIIg8rpiTg/Gw0pcGPxFtFBOdH6emXwd5Pra+MEJZ
5Kum+p/z6DB1aA4tYced8dZ6SVfPkXE4jehxAZAvmgBlKm4cxO4QlweIjqVKzosz
0jSfNaCR0QO0xfKsooYIEZ8/xhUtV+bVIy+sJqQP9ed2KJITmvadJ1yIwWDaqDwz
aAw2vSH4dfzA++Dn4PQmre60FHHtJBLfyGFpq9u45wnh0s6ukb2ly9SOLuKRobD/
/nQUTPsJP+VItBGXHiQLFXqEZjI7QFyoc6c4Cb0qaVzcm73jGgv5VM5ExZjCzp6c
5byUDvEEWny1ClOHFtmVmG3LkS6ZN30P001dk2eMf+R7RP/u6ULn6CY89mlwd+T/
rsJLZIrOh20lkT5BlVlP7g+q/8FNR15BqVPwb2b5IgVFK4chhyZ523QxqJChSyNT
811NUUqCBaglKPVOitChMskKkJ6qHz986JfKK4o+ashsBsSfP9ro0QFhBiMq6KkX
u7NUjb8D9+fRnbNihy7QdI5JQX/6QFHzlyRCFhsnYHSy47jcC9zyL9avVvecX3ZQ
OBAndTZAktmEscKEAPSuNX04uGuPe8RP2D471rNYfFgj8+KR1eLSqQQHR7vDBjTR
TPXzUUhxnaI8duFzs2Oknkw9PeJGqjFW+7irr39btPfP0jKMrLYVyn973uBp226r
flsoYuWGgkQE630vLWO9ruIBWT0GqGZq2Hy9EpaDq2aFrmCvpqdfiFkohqWhpXRk
B25VGAmJxYnuFCiWi9olBJHK8Bg16IuS9Cd1cC/xuvrjeX9BLAJps7k9cSU1+/GX
pUUirH5YSKqL5TBHVrMnciAJc+/enMEagwyHtbgYUxtS5F+bMrIBV90DiqOefvdt
00QneVYYieJFyTAKC48oL1iMRNlq+90XLa/yfFnlIMC/sjoX/fBHrReU84FEQgYG
NpHYOhyx3U4S/ORQxYLNs6SyMEDr1X9bnFy17fHdtKk4AOcGykfWowZIlMv8EZZE
0LOmO84Jsb5GiFNL7S5anuB1CPvQK2usQEHroIZBShzpTdyg7tjToojY2+90SNQL
xv/YWTMBg6cMYgYvZGArnWnuYE5kObeGcKRA9fytsgkMbGJ47Kb/ljmLwzVGoBOd
7C6QEw8gEY8DdpVMuaWAhKt9zqCItbcxqzafiZ8vZc/KlWXQib9Kfx+VUxGEqkUH
y7SZFg5DhXDYUtyrU23jGsyMVjvpPgd7Dgymc5zsAjhsBnBDTeKXqUgAHAtoncqb
OuvBJQju6ryB+LGtSffMjptuxMKXE3pOuw6TUlJlJUSjqXNKlWxM+rH/NLlR5tyc
mo9rljjuUlq80mZhBL0kPon8hKkEaUrfOaOrfyL7YqfYul7zgU1MDRf1WpDOKMHX
wTRLPjSlu0DX8Mtr+AcnMfTjGgWQF9h4b45JcIOzRZSXc6yr18nCA0xc8B3vqJTu
nV4Ey3l5beOIVtdqN0jm5zHeFlZax1+JmDl9C3G6SmhUXaWwVC/a+mgEUDWJ9SGp
Y7pAsCvXLd9yFjv2Dn2Cfm4RRI+bpo7ER5hw1Y9cnBOP9wFeZb+3N08RgeIiod/t
acZWCCrQx+BvKArKKI+KxSZq9jvN91jTOcU5rfpwvK9ccyLs9IGBfen4Lgxfa/x1
baU/NBqZ8o/5OlZNJww4+cbtYkYEPGTgeDbUffCIZ6JzDfPxaJEUApAN31P5pchD
R0/bucfV0UBxOOTQOH8Y9zj/vuqmyzabsuplyh9tXFG3k0KeunaL9U6aa171Ahce
MESOrOL9zKxKDUvo1pkV1Vnpz8gO//jgKgkOd/8Um8TaViIuCxHfr3G63nSv9iLG
aOc0sWa1asPKyTDrjOnb6wPQ6c2qAked3Q9YqzJ+GVCRDPEFFZg4upDyHUPxckac
Z7Fm5LKObsDVCY4aWsE8URGBhmSpFUD95vv0c48M5m9Lz8MHRZeM+mInBB0O8F2K
szLYINzdTRb8z3jQ6SbhXOlu1asRFmmsQIEsaxhBfr/sJYwMVL/CpXp16ScvKkek
ul8AbxsNw0ZwjGSYIEJaBGxIEAgMQnNINQB3CWnXq3ihYoi+YgAaTs5ZUgMbv0PB
sVyoHB+hsl0FGmVGnxAu1CLnAGC3keEp23eiZAZweVjDuXh7qMdaVxk9XTElAaUo
Iv9nzwIPtAqdbCSzYCOznhpAMtVf3a07p0HGbyiTQecM7UKVgfMk+1/YR02wmADN
XBquyGfr/X8lSOy96OulhroytNcSSx8CbpVN4FkpKyLMRxC8pP8GAuIuniAe0822
A3IgFcthGVjoHKCEcMzbqUTvhcCoSAIMBd23ljCz9IaDyM6kABkX0cHw5hSF674n
tg1t80Hpx6dzb76y5H01ve9+SMtmwgSNRX7+ekMTVAAO3egYgdu2v3IRAlVwkkC2
xu5AZkgsm2HQIM7ZdOL38fSOigRCUQxu3+tvvqDrMTTx2QL+d2//xOiKOFIV1jtG
3QlxS0h/cs7S0s1J2kaw5VX2BvC2M/Zh3v4a3wRVhE5+lesfD/LrpNVWCYdAfjAD
unk6YWQ79+IBPU9qEjndDxYnWKh4U+7881AlJ2KrK08uVY2qM2Qs7jdHrUC3TNbe
Y/zkIdr+J+bSEGVEtRejl+LSa8acVQ+cFP2bVseQDfgq2HStRELNsDpXhz9pqB9P
cWluQ7a2gR9+aa6YSm01un+rSNeEyc9YuJDdm5UnTvkxQEUuQy5Qxoqptrk+QrQE
PUCFt7yos4dFUCiCRvhJBoAkNWeAa0cFqNxj7R47XGr8proibYPEmoUVANmB5vh6
I2tYxbaQ0K8wBsqKu0347IObzD4gJOkwoUEFBTeFh+Xbd8AXoapV4CKJasze9nx5
ZehfeF5yKV+7/mJuqaQj3P2SoLG7dnrFVCUo6NAye8xug2aakXjHRsMheI68QqB6
BhCyQ5mJOKN6viF4b50039D+IGti4cfp6O+pmGxb/Oq5yzBjqxTJ6pglJ5y5NGZ7
RDbsBINlyqUj84hKCFFOxm78JlbLLb/LoKcGDWjfcYn3+1/RkZnQdRmBuHNIqfXP
kFgG/50pDPrSZAuluUaXlVWp6P6dMF1UpdIr1i2K3KdJubWr3/L9aEzugiXzeJSg
W0bl4H919KQCzdj4e3CRQ0p043NKIdQptVXnIzXp/D+PvUX3Z2IJeyFQQ2p91OjY
e9f4pyzxN+XvhGFoyl9upi/CiLAdgnIDu0tKE+wh7tbo0hvgksED6N6LrgvakxQU
0e+GAUfP9VzwmMXjAh08R0jqVEaQL95O8xMYOnLu89wES6OdS51oO2qeQLCVhiX4
JltwhNJonGg5XT76FgMIMM6pgPItcZ2PrgotNnEwdaVRDrw/nPI6EvXAwa6aSrxf
Ko3W5cmXi+P3y8XaqGFTphbML/xKO0VkNMOZtcsA1hu/OzwfIoAggJbgr/pC7vh1
LvX5LcndvbUiJj60JcE0bhU2dnog2ENzn1VleYaD+MdNOAMonq2QvqOAYoTgWndd
PgLSHOQPquk5dIYHeEB86+lgo/f0wR2jLDgbAyxHZasQtsKL7zqPDzurjaXhmzwd
xBJJL4qa4Ys2CtnTAUXDTpG+RWO72orGZAZCILTdYNgBaEkzy2f6aIRZf9woWwO+
x0kRIGlSIQ6uDP3ktwLo/UHOl7iGGm0LShd27NacgAv6I0F+glFgzppWJijMI0RX
vvBRFvTvTaz6oH8ZEdnJgpYaIOWWeX2MfrxukQQf1U5juYB2ALRJTAqEHt75vYTd
brcp6XcqSMtFErn1lTTkAzEIsZvs+3p0cTvI8u7FyG8uQS/Dc1cveRzYN/i3YPFS
KPeS8xxUmohsAwV9O6SG+9sKhhrF1yZraj/VXFRV8hhgAx2GU0YjKP3nXt1afhQP
sEBPypEGq2/SA08HgwqhhEx7EPGZFH3lRQ4DvoZbwOBbWU14BQneWcTxv/rCAFAx
YB8gek8YkSbZTboj9OsCmttwTyxfxOeejz/QLBGO2nIiSxxqF+ONxFQhV4rnn/M7
YI/uTjDvJxHnItIIbN8PpeUzco7apoX8FGe9mb+6x20kmwQ8qnnHpq98TpVLAPcb
rowCF8bEwWTke4YeZDXULqxpsgv5xzcm8klh01uj9OBTQIXd8lGPHEkkAKWqpqM2
vSdu9zK3ynUTx4EDAKiyVQvndCOEtoj5dD2adbuYi9Jia2qV1nApLH/eZy3h4h7G
G4Eo6+KXqCcIP/fciz1yV65Vekr86xb/shtz/eQ69WMigYRoPFcFcXFO3/ulbyFr
c+lC7FaOcSgeytHv1NF5UtFeUQUnyzyoEbBnqcWiZfkIOFwyw2NHjW8BpfAT3oQn
0pWrYrnEWGR9EL3Qup2CTZyGWT0jM7a1gTBbP1lvPbq75sucX4nxyk78wDBG7a2j
BtGr8PubiSJmavJbLCyctRxiR28OyjjlhgrPu3NV2rVKLPEgCiuhjLiG+rBzxPpl
67doiGnc/IwN+LEEVvwOMxpHt9ktIr6OWaOzuM+EQpmFMc0v1gi4P9PA1ofXWh79
w3wd6KC7GvNk01jkNuHULj3Zc0P86JmbGmUdJ6fsA0wCPVVzSUR3zPgW8GBr0fre
EW/brvPTArnsfm5xciwpYv9DNoQOmBW6FvR2skKAH6sZEEeFU/Cwf9SUkTBgBKg2
D/xbmt5OqnFQhHz4DZ6wizRs1LZQfFl5H011bsXv1wTbnR4eR1vQDN0jTDy27AnU
dD3JwpD/P4WAiVyBxJlsy7iz/pPAnMtzD3ET2108EAlmn6PSSRsV8sMo8s5ZimP5
ucm3//fHVFwX46XxgrBDMbAsFNlNxLIp5RQdmRbcSB2yzRmG7d42k2h/B8ORVkJi
0ctfqTvPRJR4dro4b1LCus+6oNBRLSqnJ6nNKqjj3EdwW5E9x8pz5CJh2kEdLTKt
QhWt6EqAvfMOxPiuaw28f8mRsOlCyJ4RG6uSJygi4P+4+90AJ/fum/E3BEh9/jzd
LR856LPn7EEdrB66fHqZaAEpKJ9VRpnbtz1jROjVzgL/AeUqa2p4r/UiaWDX5FBK
129BGyfYU7c3VMRrDAt1zn7l1eANjwrt63kqPLChTlwb+lQupKj3Wfx39/MnIL3B
QH91A+yIsFVIeDieIOuh34+WzPErXPYpmGbnLWUfbwz4Wb6s0twZxUe64p1i2mRm
DfZ0jiIV/YQXMYq7uLCbnTR1SacYLK1jrma8aKXVymmJRJeJOH9gPEdOPwSqUXgp
Ogrh/GSFzRCyG8W6zkfMBTtNL2VNRs1qdndjn4v5pml66K+7dDAWhNIJdC5eDI3s
mVdNpThSp8mdqNLxouKq9oa1y2rJjrATruDRTn/4hs3Ckg14osT2XHSGgGlN7Sw0
dz9I4bNwKdMNoIK2z4ryM+83OYex2oCwA1IGW/G3lgGacw+Wg7K7QiK2zPTWZT5Y
RGwq74IDguHAJe+KHVGpZyPK/k/XQotAFcL52K1wHlxfXDhBsWNm6E9wMO+tAZWT
tjk9FqX0aMC12GYZOZm77BQsLzjgrVVc5WCRbgK01gxyc97SHlnBUS45Phski4GK
O7WpRjKir5Eeq7SN8Cm49pE/7VBGRffWUGJuLhcsi6erzok/V7LeQnEq19x9wtCH
XrU7zs6XLRIdoGEEJ+j+ue4/xy83yap9bVze037MONn5ZkDCw1cW8umyNzsjENQ1
qG6kXIKqjqgAhf5PxfwzK4ausneu7CN2AXjVdwc194jXEEH+4iZCdYc7NLnt5foL
oFGh4IIKWUG+zeiJDWG+/V+gxfx2wbm7OxUsyq34N4v42P1TvCM1lG4gzVPt5sw+
7qxp2pvRrcO7UCA21J4Ss9+lP+4Pfwf9Cws8OPtR/llKdlY3MyVY3uRF/tE9dYMY
NYaOhQ55qw6KX7l/PSxkMckzCEn22VOc0r5tbp05IlQXYSv7513WvmHPm1gVGYV0
UJ/p53K0zzqxlT0In/ZrFe0YxQBXGjftmpGwMVSU3C7BKZltX0hdH6SoZF0KrsQG
lyQGjuWuyYqdPad2FtzCgKigmwCW+4ltYuRZ2BhM98gxp68d9ZOqt/vg483n+n/R
kDF/eGTciwlIuHlPwjp5ehxW9gTuDaV28xz8hThNQJ1vU8r2YrAsyKYsfuB+rwc1
tP/1CfUD6qSOPi1TYluncMur9R2PHp1XKH0dcsNhWJyniNacuufiq9PcWO2hug1o
zhcmAG9ei5WosT5w5mUxVGx3LIDfW4nTc0DtOOETma7yn4JSFyfYROsPCd3Q3loR
FIsCw4+Pl7qI/je/cRGWIpzpQgTzmbNPa5dofjCrCKff4VL9+kfTQDSIUOjRkxEP
AxzwfY0o24yOiSsyFiZrUx4SXTjVoFQ9honw+H2JbyGKK0g2wJJSidam5KRakRJa
kWxPC8AnHpillarhLQZAhiOIOEzOsKC8ADZEYtJk0ngrn8UVZt7/8ByyEWSLL51b
AmzxAB8lq+cC8S2baDWnjny2Atb3brw5zFTQpehrGOry/3Y1FLXXEBj1cYx2WPAA
9qc34dXsuH/jNgAR6AVKRHlop8aepNqfa4ONe0cAvRP0+6k8UzMFg87UKIYGtWIu
WsTcmlnBKQjXFSOci5ufiar0z34ZztaRLorb3nS2cSyH6k4DjYOE/yJW7LqmV6LB
WKwKD3zCTMmieJXog0QhNDCEU5ChofuBWAuACE5TURtIg0LjxHHVSWRokN+0hgF5
d7uWrWSHeV/JImnxtkMCVSldCaKOsiMjlQXLP8L6fFjOJgQEPpQCc0ufB5tyJPrU
cbXchAR6mqg63sPAZSWUjcMtltE2JuLMltxkp6ubm/lP8EHpf1Xu5kRta4+Ce7OE
6Y+7kq0k3OdniTEGgP/kxT684qKBInIQ/xKpurNYgll3QcDittlMD1L99ZMlBerJ
vx58jB356fBxQrQKDUi/8Ssd7SkH/0hoJMp9wvwiYo8Zuja7mXjyRWruchFp9ncU
Fhzeb2NGCS5QY8HDL8HN4GUikET9U5sMSeycc7KljhombKq6U//mkxqaREdU4nP4
/v1RXE+xnGwNtUSPgWQRAKsDVmO774pg1ycycsED9rVWCHMdefQDuN0VJyC2Ds6K
hBeEUd41+ZqiECSVcDgpfD4wAnbEuLNsfuXddmBeCokX6cU9l4m5vHYus44MNa/S
V5eKF1Js1aaiCGSiR6o+QczAbtfACrHFmHvw8esb9+XIsVJkYwdl4mBhaCgLggLh
UZ7WFeyXz2blZHzE41HW8kZKnt2JDLyStIHWeo+hyvcmZ/LGs8LDCdf9O0leP6gg
7MNjJoJaEPaMl9jmVPWanu8LCr2zoQCq0pcuW3B1i3mBQJjQ6p3TLmRV/s5Gpua1
1hjh79eJPIPKVOUIrXsAGZ8KI03MeXHium804C1CoatT7GjAv7cEY7SsLxHj3473
7yiD6P3Uz1I/Noa4bqhGpK6hRHu0NnDHlfnhvdGmgTHZe/K4WS4oI0JXW+me4qIU
3vg2NlTgcqihS9KrUw8I/Jgh9+r3hn1j+FMFVcE1YMD/0AFfynqxF6CAz5tHd/5g
lQ6HaxgCdQzZrkwqncfSTz9x7qyev5TH/TME5XOOyCIJoOQuKKUb7CJ1PmQe27zE
gcUE3gXG69IBGsjgTs1G8+vP/BUlaDd6ISI5wWt+dOOmdLNGyK+JBjS6EBVAhBfz
EhCfYkC4Dq3Dn1iRPp1R0d87GXluHEhi5FF7V2Ko5Hci51opmgJCy5FvbUFGRR8I
/HrU0L8HgZjA1rKdnOJxXS2x8YkJZrAX8q92uZqQ3LqGY9/O4ZtjbgEXR9qOCNpF
1pMjEBw8r9BEQq+nV9U1oEUfu4G6gDpSJhYUP7IL+td/mcaHuVtJVYz73sHOo4mS
O5GOP98RCOwM5DTRYYm+wgirs2o1YgbUniGc4RgN1gy3CKK+07WywU2yGu1ZyWhj
WSyZbcJXqhpJjRprJufu9CsmicbFXC3QP2XHkBDcN40rY4hgii+0EHSGiJA3/XJX
5AtlnzjXDRBMMut1Kt/vqJf6hQGepDZKgG4yjJfHtv99xWC44488bRss722T7H2H
A/JL8Lznx+5DtxLmzS0JXYDVzUklUqIrX9YyP0UzzuEVU/nyvPv6X/Aph+dvd2Qc
PXdT2X9YDCPI6kapRhP2cF77BMKCuWVjyFmxnW5nwRaPric8mbdkKNz3u6CHODgH
k+LLVrCrwNQziEKTWpFtvKZAve6x3suI+WvlDHxYOC773h+IsXKDZqCEaG0hQ1c6
5DeTpf3unGDgM+10xDfQiOxJBEoCrJVxrLVsyDf8Bx5NLjOZ36Mbt/kjRHjv1U/9
D1Hcc3gwyCCrwabyrNjcr07eRnOy4eAlZGIBpay4J5NTgOh3gdd8UBbpmjhZwXZL
CfzyEjsiCkZsJugpGbr3Pj+0+rMdpA9nZwwwyhPRC7KEMcnTRnVYYuwA0Y7KxVBK
tQbyz4RjxLNVLGG5jZ7/8wPp8qaGWzscdSdmhSs3rctIAqmqmNaHznbf2sOh2Lfb
3JLlgVFeLHfTPEVZqY59BzX42zCwv19hoKZIfauQWqlBNF3GifcOZwfuaFCJSu8d
ZSTr8kNMXvJNKJah121dEUM572V3pEbvgt0h0WrwxQWG34rDJvkVPeeGgKN1LBxg
FO8UYzEDwecx+UXbsGEJGhTkgPogDhx65K5YVL9CIx8+yaHrjLRUBtQthgUWIHVf
ei5uGyZZFsYkGwhVORQJxGV/YerF9EgATazdxH0+Kavo29q817N2Tju0Hbj3huFy
U2wUWxi4UrHBjKw9Jw0XX3dd5G8V074sVzxeBOEaR3GRPWQIMU9I+BAxCVDJl7Y1
CfTFFpDQCGqyyqJ6rE5325XptwCwJcvCBXyy4ercdtLgcSlX+TVjoLQsbERLlamy
Eq2ZGbF8/dIxtIhiegt7bx6ks6yjht8Y9RJ918Zs+zPnCdLi/BcVVuvsSmi3pBnG
9tZOWCqhGKMrIuwWGEkTZuF0vmiIGM3EBWi4TXuEma0bOkJFSF6+q8rhwVB4x/RR
wEasEb6L6euk5vad6G93czji5d2zV/xnbKu3KNtaCXQXkfWKO7PHF1cXNm8b9oGU
gTn8XKLorN7ul64QVII3ZeTrYUjPH3N0KDIIMXTjUbtGAzbn5wCLjEBZqRawG2mI
dL8uClkp6Gs/yP5VTLE/+uZCmUXVoVlGapcPZX+dQq/c/G75UlOLfPlv2wFVX8bR
UwiNNtpo5tLpt4rULGUTN8HG5LrXVh2K7+dmNWoCvjA1eYaex7OOZmoffc4KXrs2
nkiuuyRly0ucH3gJm2dhHGFRrkh7A0c7B82Rqw27ctiiVXN9KmakLWfQV7LWZNay
taYRCCr+V4UaS8PGVzHcT8Mp7c2JCEe1tKwhbgytkqz8pdRePeLpifDraY/8rI+S
KUcuKb9lTtY5M2D3X+QMzUQ0Jey1bJwuWVVUVf2hA9siZP6a/7zIGCsmBpJM7smp
WbvzpKQs6qOGJIJNWM7KsCKswN1vjL/ndN2Px0PeQHIp+QFqZV5wFUeB+F+2pDPZ
/fTDvUkoEqQb7GnmQnQmNpaA343LwdE8ES4uPu4PAnAn4/yTISHIyE1YO9Xs8Q5y
Sq7FG5JK9tmw7uhUwPG44uRT5J5mqb6BlX2OKRpSb6DVfWzRZ9wCMjVmW0eHuuD3
bWedKnLz4IJ2dyC1hNSdLK9gM24LexUpgVp5LXLIlU8ZHbkGnygTK55IF++Ukna9
c0cRZIIofxZMwpfAOBzIg2KTAaE+QJwcLOOJoy7d+XPMCuRrZcp/rU52JUUROWjt
7HFw6VhUAQns3rY1vy2ogw8Kc7QT0G3vmb6PSHPnjD4GFD48ScvXyHZnflu7v2/G
sHtDk33fC+kGH9fa+7JgYGGQ99on23t388hGcqvTHWYksgSShtF15+Ocl3TToicF
rRlKcDS5CRx5Nlj5S31NDdW0O/9krgnmeWmbsYeM4WyeXjsvII1lr+DwUE0gr2NW
lZyCOWBIcnmLGHfsFKAQ4k4yJTn7LDBLlO5K50nCIaCaaJ/RFcNFUi7bKSCiOqXq
7mkQKAsWd5gVB7YrgSmTa11UBNf1QwfWeav9L/0EaAJB80boCsV2rk2yeR2iRFbc
o5N7PKRLw8D5lgae9sJjeislIe26AfsG1HILTQCq4R/qqbFFrlaOKqd9zol/36sr
Nl1n6Vvw7uv5z8z9uSE5ffGImzpo2cu/Zt2Ue3r2c6UFND5AOaIPadyVGLqW4aLc
G0x0oyrSFhaIP6kxjFXtNESZcOsBMTJyH5jf+VSvoYlq/McDC5imWpaseMK0DaHA
79PWmF1Gfbw920i3ncLr4L4lKpa7HnAgz/kl/mRP2zv7XCTRiYmriqP90D++HH/+
CYiVt7keRqvmzYhgM+pLizVppCCwGjdPmd+C6cJJSYTlftWbkhEWoYg+avF/Sx2K
N/5xz2CKpsZxO/JUillusulAtPpeIhTj995p6s6aZ2txMJN6TeISz6bDK5D094Fn
siFonW/IoxIvNDMUKWm81MhNIdTEZevXdlyDlwwuEMfV3DqghxTf2sENkjQLjtIq
yIaTstwVtvhIK+w8GNvd49O9ZuOmUaKE3J/7rzgJuWIOO4kDvKG4e6Qg8OvWzF2Y
pXh/nfmgcCYrh49JPpj9S9S5ah6O1qmHCzZUP22kMvPtZs4lLuIawAvsolPYrFhy
gz/WyAWPM5/apiwvdcfikxqOpTDoBD3vf4rWaLzB+EA0NF/nrhawAFDjBpYiqxAH
UcIjoTj/po2BRnJsqcFGxDulSJPFRL/D56l4Ud/Ss3r2IIiHaQxBweIkZjKmdWqC
7g7jv9FRsIvhjykZwSsetQaiL3sOT/QO9KijjEnDkxJSZQdWJUGVaCJKpp5X7dK2
F9/kUmfqO9qf+lViWKcy91t+eGc7I1i/hWiWScGEnMPTZhlD6rqVXMoBL4HkCka/
Lg9Z2uSS2UVetuk8F2PLFyct+N+9dT3wAQXXa3R+lGhBbFm3ol8jPZGKeiTJ+eJe
Q7B5MOn3oGccewL2AW9sLGg8I7Ci3KGLZVYqHLMfHk7BPX9U7oGQdJAdhBHG39KY
Wi8QZZWPJNnenJZiZfkToS9pyTG6tL7Htl1HwC62PuLiIL8uX/jrqQuXpvKdmPOJ
ZnitG/okkXt4CNJquBRjCZWkbYqdbA2fjVZmNJgJvq6C0B0DPhNa68X6X+6xYYdB
2Rj6p+uzRPtmzc3BnAJm+dQ7AhcZ8pxTjwZENqsw8Dhg6M4EpvcGjA/A9pWYOECF
lBO8iEsTr8ni6zIambZSpCWXnyFcvQkoqX/bcpewcwUoPg4QglmAUw+yVh1thGv1
bqy5gDM8tKdhOQ9AUqhoyWgnORc2vAjhDNVYc2Gd4Qzt8/wek16fEPzGmuobaVmO
cUSmRbUt83TDBqhQo5o9lEDsZGe5xktgcLxpL2PCtkI6LTlZ/Ibc8BAY4zZvWjOK
cVwt3lgb4T0x9pcxnVGsxoRzVPGpkbvN5UklPOHkrbX62tg0LHg1KWCies/5wr1Z
7+9DlXKrv2cU1FFlNuff2xUcMQpAaZGtQwjGdZutq471Y26f2dyLKFwQWY7IjsgY
4IMR0eoPzyuD51kzWafkiRNY1OBBoqy7VWhP5I29uV+dkZRit0K1Zz9ajljsk37f
2Y9g5Ptqh+U3Yv52a1l9osDTIj0Q31xe5rZQurUwYDxoVtWj4ZiKzWXy7TlzX5zl
kPxL4/2a/Tyh1Gs8QqOuiyeSgqlXvYB0bZNI/5WpoYhJFED5c7coWb1NM/pMuxk7
ka990oyuyJEDLKOm7uRcq1evP1PLVBllOVqEd2rGh4Jn8WkAjhtzpDQaEXdpQC4o
lTfbhqdo/MrWZh6CohiYogT8y2z+xpVLc/u2tPhfPAPhGCwZ/JIHpydOzzHOXAZT
+x0G9ghxhqHPZPvUCEgaGVeQ59B4IBNlNaqp+0S7WfqqYaJwc54ufLqrTctslSHk
ksxqaEmdPzLMCs3oALOA8iFOvA/KF7+ovX3jSSAdMCGxaZLE62O/KCQOwsylXcXp
AfFXS3g9QWdM2ouphBzyTI5vJIa0MOSULeA2uzhEKamnIAebnPrCIrhFGuHDZUcG
kcJqJM4ozrT88fMY1KGE3bHZaEYM32e2q+ak3ermApOi9sgGYIhrn3GD3IyQGKlG
zU4s3eQzuTD9J17izOsI80MGgbT+AHNxQBhGg3FMHYnz3GUCEBPY1PL2x0QUc/WI
RNoH17uXba4RigU8bZpul4Z4temO9IRGR75MmNyBhzIA5oAbvo59ScYK5D7YzJuo
56weiqpnEI1FjIb15rf8qd1Lq+Vu6fJk+3QjTJkf/+0Kbh+ZtPIwshmpMnzEggK6
iDDUjNW5nbQqfQH5q9lN3tR0LI+OEnElPG/OnjfwM4WZyFs9haPQoslqNWFURI3J
jp4BvrqbZ9dhSo3fNaJ9+WXrcsslPub60R+0MAwzrPdfmufOao9c+5ap+J/VUoNR
i8GlH4rXZVkVRGG0Dn3l2lK1Om8FrBg0aN6/es1FxPRXKHF/qWwGxa6BAJU4bVre
AIw7j95BaVAAeb/qq3MoLCBF5KS16AMMYkCKCLKZyWnbMaZYZgpnWzkX+wMQu1Qq
9m3YCH2VgFolcpAYw7bdlXfGGGthKawSW+l5LOQ2F8i37U7MamYdqMmEUX/UHZTH
1V+l49bLnlg/fFkI1IDYYXzKL+j3olyUcsxvup0fdebsECfpZA1V+E0C0dIYebIC
NsknJjYFO9+pBsZ5e/78z8Nr1hOjyxFG8oIvy5tSbPjiXCwFDvUSmi0oC4iz57tX
8OlMLBCtUHTZtULDe8w6uK1Hf2onDxr6GQqe1VD1KK29IezuA4uUk38uwmQqPOlN
DnVXVdJQe6SQARClnnhHyAUsJOMfTFUP4HrI5L7HK+nhxOgKciCF3uOhKqICVITo
mdByDg/Q6Su+EwtsyrKjX5xlkno0/yo66rJ+KYsrxUYX901jsRn8AjQirwv90zP+
wiuMhj/XGlbZqkUgvlwJX22z88ODdAKjH3WQDkaETR0OyHvs6wtMyV5JpSsmtnJC
K0FE8ZPzg19nN+I5TR7d2zbg7ywgW8Hui7gvUP/b92rntpdQO5nJAe7JIRpE9lFl
/8X+IWPnJjk7G4Hr7f6DCWOj8MNDZWofnTiY//1pMsz492cMxIcYbhFB62JRKUu4
jn2Vmrg0srFytZBxxp8TRiOpHwoQNN0hqQr1SjY+/uLWKlzp+1oImI/c9jempPYH
A7QPgc4Wph9bhldq9thbil/vq81Xw2QLTokLXLfu64RP0L5e5rxpjjxmdOLH0qYH
54xHbQ+fNtc5U9iU/Qwg7WgabF1cSkJ5lTsKJsqZeBdaQQur7FOQTNVEmV3H/1Ex
vCnWKyRB6DQxmHl8xFattTPT3pw5aiVg/NYLV9/kSFniEf4i5knaDYxOp2XDnKLf
CUvdIf8ztuE7F56mqPJ4i9FyA4tUbbNux6hAOdgBX+An+Qi3Zme4BbdzywsO6tOR
CmcLYfrB9yo65bcEi9336dq8Q+zkJPUiPc8JWte1+3/cYCKOCBwlgCL9JEuoWDwl
JiQ11uTwqpj5ksUHCn2DFrvYKipNnfhgqOZeRsQN+j9IlP6tag9lj52edtlFHVf0
qga7fyRq/osa3DdqSeO6Ff4tVpK9bEjEwJVdySwFdWCuU6md3GosZSI3iNaFGPI3
u+15odQUZQx23gUkzfeePULpM+RyDcy/zeibH5zIRe12wjr+9sbwAXelCQPyDyzz
RSvYQ7HuuoBJz+g8LdH7YIr2BMaNjVImhv3hhV2WPDMmUecL5SNbsxVttZuaBZV6
/SamBBLrCNBjfLwQ/t/p3hCCRMC24l5iQ1LxeqsxEmhHFC8zdvk/m0clVdb/mpqt
RuUTKHA6cM/hMm1uoiHCUs9lUab1SPgRqrnSXEEI7tScaFDo313bm3B+yHxL78+f
dngjLtdbPon/EQlhGoq9NzIBzq32mL/ColCQx3sJmUG/O15xubpbZTCQ4xrBA66a
UMicBehFWC/drTt3L2MPOJ1w8kB8aogie/B+81SWSIhe9+nrio68/G2qqT8R1fzU
xeKuGLt9HWw0O7Cp0AYTK8NhjDVzgnBs5EDWQJ2TsbJwn1NfPQHK5gpfmKSw7ps3
HRQd5L7i0fVTtWI011JIFPfB2igNCtEynWDevJ6I/krm09vZWUOw5NldBSSUTMpp
gXPepHvp0vYtKbmn0RF5GV/zKfOukv0YpKXCg/iQdrWdwH0SiW31jlWUt1npfvm8
7Z7lkMzMpdCxthZlrmKRIE69HyFARkbZVU/eFMSozsOA5JJ3XjR/HemAskeaB8vp
o8gK2pwCqEjR3JlBohG/dgOJ5TINRbAbWViWiv93dS4YmWthNkaNbxTVNRpafv1o
Es8Oflg0bdoJbFuGuQ70Auqv5iuhApObIWAO1gHBjAQfoZ15twLD3IWpnXYpVNso
msCd/KGQGCixjEq4MioWZpbZatgm+7jzMDLn37wdS5REnV+WmAiiuWT3Md6y7MRE
VKTFYzY1Mr9YqKfmKa6F1K69k3VBuNB/cp0petCCfyum+W360GBn4vro6qKorEpr
rU2/hDuBWoLp6C+HCmDezbu6qDQROhmoq+M2UcCoV179iE4+I2dI99xQpKLnz5Jg
kEuWht8yWArQJHsxHGsKcenRZ+ujA386DJR3yYVtPHjCFhgJTasHuNzDmBhxoNKW
5aCerZvNICHEP70MmCBnCIqaMY2gJpPkaYqEtgSJyF3pDo15Q9FIeGOg/B0/6NnR
pT5vZVFUBmRZJmlhCYLYQVrgSQJ5xSV1P8SyuXf+azf8u8cXI7/NilS+urNrbwCl
DIolBmb6KgxzLkKC72MgpwAmtUMFVbUkho+weg7l1uJgX7SDqrE2n2FBqwtz6vJz
gibms8el+/uXiiFNlMTtrmA/l/c3GgJEJv+Az55LQrm1qqutRBfFesSSzuuJg0as
6MhX5KnqnrFis1XzzqvGobntADjWgKlUwnjQr3dCh/t7TfNtjvRKq/E7cBRAILRH
Sk50K2MkRHXYy/mllNk5mC470hjDXfgvUznKSRHrQN2wD4LzX0vWP9XTaW1eV0DG
Djcm1hmx0HtJShcsVjjQFPJnkHbgcuHs9uT9q6V0AzhTawxcPZn1WjK2SgXQkviV
2hrVeRVQ0mOcTQ0aT/3a74o0NfZ5TscBvydrF+2hd4T1dsD9AmVtsEbLMVQNzGYK
ryuyEh+vEQYqi1fdyapHQFXo6YZRmT3u3LiXux7mKtPT5mfDNFCzyEwU3sKzGimy
fL6CGBomSiuxXYa17dWVrrFn+Fx9X4laPekflU49ad9tBSz8xV/ARFD0BTp+m4Lo
16IuS3YYMhv2yI47g8Wf5Kkj0kHEAdXJTv6WuKrE5hrrd8bvj/SprlU1Y6YA/ht5
LGVg30n+bcXfSbX53zqCmHtYsNQIvcISQspM+2dFNCBn6CHCVQmDGbxOFGVeoGHz
ZcAzXdQj8TL5q9C2teYkmOmta+zTDqWzrUp6Fz3bNY8UITDSP/SdKivJmFpC+f01
+jEOSpLAafxg7WLtNnQtWPec1dPpTof+zVngqX65o4Jj+xWtnLTOk4zT7uAFXRZg
hKTkzS0KVtyHahtSv0CkbDycaB41BJW1lNts1++tVBfBegWdY+wzQs1tWQ5ekAi3
fIkhikffYlJd0TC3FOWo2HQ1lDUaRFtzY43snpDDnbhQF49h8Igt/pIgvn3eOPAB
nrivz8yMSAOBERO9GpXCeoZT1X/W1sTIQi48wd8rLtoP8FWTIS0mNbBrb0yt9MYK
5TxhRhgy1VmDmsd/lFNVL1OnGOnIwhTvOsO0eQzjPjo0K/hNCXm2Ms43yJMMo/FI
90f2P2kESQ1Rf+rbbDoKPe6ANRyHloNb6Tj+WYavQ56yfsQnienCMuG78iMZ+jS+
wFGXEAeRu4plDl18yLK+MV1DzNbU5dk+jOxAyR0SUldCAWGbr8nEBPFqdIaJhVXk
pAujrmT1ya51vNG5eSrkJW38pA80N66gJZVIwjSxjYdshxfX8mU8nDh8zkTDeFvC
7slXpfzNRxsRh36Tg2k4fhyeCbuRxRE6mzasvDYFUKShpiqtxq8bvVajPf6TcpDX
qHdYwS+QmmsQ6fifn8m8AS5fbKGzinsqlBfyQIRYVLbK9h2hfxi/fefhd11ObDP1
KxzNXxur6BjubQdnOSAgGD0Nx+yRQCP5tOhBZe1NVafpzzKEEyXNz31SvkY7xALl
aJOb9HNjvSeeh9MVohS0MCvlfBbPG+mWXnhSuY6vDXjk9/WL9wd81xOSZ8Bdol47
vdAecMECXqE9BvTWDJzxDSNwUgdY8g8IlO43ievBJ6Iuv39Z5gJjq9wleQ+Wc7HQ
GPhxPH2QlFPZBOiMhOEhFaegw1hdILdsGnelyfbH3iXZ/wcN/4sB1myxGKw7bNKd
nNVsciwpMAr3RJkBg8Ndc9tnSMexNpVEp/PolfQa+ldAAow8+fZ0e2B124WXVJwg
re/1O2xXPOkerh+w82ncxJaP8MgrOlgfF3mcWZNlV4LKuur0vBOmxwqHebHSSxcH
NWn1kUuEPcc+Lwrqwksd7W34QrvsQTmIq7+GTPCLuneAdnRxIGnpnN3GQFNeX69z
+Wi6BDdXspXQvKeqB2g/8+irEKPZbH3ajjZF6zJSTASzSBZKL+RWzI/GqfgneDVC
1wmD7U4UhkQSt+0rEIxFhoE20qb6HHcRNw9srFo3oJiX/gYm2bE20le0+OFCUN20
7CLb4YrbNHO7QAB7pT2+bGY967JoTg6q/JtfnEtZeCetmLRta7m0Mq6TTSWTw2YA
6HA5n5UlZvv96PYyHHPOi7biEaDxpOrKc+cYhOb8wT03oprJRLC4OBRytiBcN1TC
IFG1aS427s2ZopoNo9oKMuu3OTYUAi69gZZlglcPUs9DKcrXS1SVmBSECTFu5YQG
dyUyx8Fz/vyBQhxA69XjYJq1QqH6BJCBEoHU6AwR0cAhDEOyrrSEwGOmPo/pifzt
+mzi578KaYeYHEcVURZxbGtzsdOIoOsVVBG7vUDs88IBOjDJ1Hv8RPun2+6olN0t
jRpoMfSxjRBTRSwEkMvmcDPcnSskoRDcfFzOulx62hBWGwqWHHXvkGpuTdYCIdOn
XpWTS4WsCRTBAryMl7TGSbyY1uCTSxPqb68msmfTw6U/7J75VUP88D/EUCkPg1Js
XPGkWOT8KBm4YUXs8ff6m0u7pCRP1niHvweVg/muCxufRxmkzA4GBV+EAWBGySoQ
00PEMSBRiuRcK1tqhVgWQ3K97Ioq2iZ/kYzmlTsySGLY+8LJwT+IN5gX7GCQbud3
98kQ8jYoO1KT71o6flTrah49HLbZop8/VBhFBhB8+/R9mkw2rAZAxb7Z5bqAzosJ
iZ+o1HQ6fIqbw3H/M56yNmsmXrt6azEgGjmlRTpIQGDP7+tALT05uwHIs4C5tFLw
vAfEmTtxrJ/nAKWMoXzv0Ua6d9/OckUZHuj7KlsmHnnJMAxF96sTRpUptx1/k/p2
ompSOZoEFzB4VhNm5G9q4h9vj6vjisVjYFU8n3j2YW02ck0qGhbkZMnaZ9nQ9uQG
OIoUmDuCdSFJJc3oK+jwcbkKweONV9gwrJKpGgkNicqU0VskL2x1eeBRaB0erp2k
7Rt6GXTjIEbSYl9iCsvk1Tp0/UA3vXxo+zmcU/HksHUjZ3E6DR9ajBhVhXBDxoxn
+dB+aPiysgN8YK5O2B7Nh/wHyj1OqKHjz/5G8ag8aOVQ2jlwSEivYzK9T16gen3r
KziI5gzyvMWNV4HiX+g8s9/h+mb4jTj1ZR1K0znRbP9ehNDle6oKB1Kz9FPP3bgK
HEyHL1CUKfgzQWp14U/kuBiBQmlLu2NF+uKuMhAPS+d1x34U0Nvh3+oHxSI56XKz
irsKE1DDiO53VVcLkev8+gCOPYgv929uCJ2RaIX15W3SokswgQpFpz1LydYwb+nm
bgOuR4QZA69F8gsKNyd02fzqJ+vRUwgqjgGz90hCWOTjJWCQ8Z3BNAzWwI5N5ndN
tZss/5XL2bjRehNrZFlrvrQT3mEYtj+SFtCVqO47klm9f9c1RDRBLMxfpkYzijUJ
spFuSes3+ViNYE7g148Ko1SyVnu5/PPly1Qc065xZXZLoW/pudTwEzJOKqmhkqlZ
uRGBFW4Kk6vaBJP2FdzcOJmS4Kq5kjluPhk9hQSzFsz2dh2nbQ1wYCNtHY9S1loz
/rowCzGUpUj5+l2VRfc2lXHFwSbWWDPl/E8sKQpFS7vbwmVJvbP7vWc+R8lRixUs
X2uodtPGLBbs7mN/qOZGRsREg7aZoiVk0fKDxLkEOXVY+DWdRib4c9MN68M9tSpm
xgKav0yOnPBzsldRgCtBfQj4Fx5SVzknSNZmUWfc0Odc/pXeN3+gl3vmOqsOm0kN
Zx71r/IYKVH4j/f28F8W8pxFkaiNffDx+MGt+gxqh7MTwyctm3H/MTzRHRuo/vj/
mCevpPlDC0n6DR/de1THo9BCsBL15HgJyrK8wIpJCmHlzsEIclk/qwYKkxbpKlWg
53Y6II6lw3YDJm/+VIL5o6QbNn//R9VVJ7All1bJX/DPvsyxMZbRW41dQYYrFRmU
iCSv4/M5uzxu4uesKLfOUFwgYNIDR5KGYVVe/cCAO5URsco+NTtY6cwrJmKhDrG4
RAesby7U4aOPsZGokUQ7+uDzvCBpvM+TIFLLo9G4hI8s2ofiaYshJNYaAu7EYlJr
8zIL8hJ78hwIitkhBmayjFKtsIj7c32DV9NCvzl+hH2gTsTa4cex1MPsfWoF6//M
GWit3+NBqkTk1u2HRYLRGxhjscCy5s8w93ZfeJpiGSmlblOV4sWfiXRwj06BBIuF
9xGze1aYwh4iM91fE9hlgthr0AX5g3qYBf0n4oxfVRNTrRHov+l0/VkOZCCPzVVu
nmM0mlNfr0CphJiTq0p9vd3fAuctaeHlGbcosdVwxxdQk5X2U+ZGKQF5MNqHBgtL
YvGgW5TgbEPokFVKg9f5bpDwa+RzhadWCMQiMxAjMaP70ydJBRLz1cthqP4F8z4/
TcsXT+IYZMC3FQcsLUWzfy8GVRg6PMyODgkrTWXSrx1icIf33Ka3DwPVZoCFfRIN
/Hp2xeDzyLd21X8gYGNa4WZOrlcpXWlI2CFVi2GkuK3O/5n6yoYunKYftywhR+/0
o48IwUjKuByb3SXcMPKjn2vj/iSw51gxK+l4HHWurlNIwrM6+ataJ/EJ2KEuxDaR
Aye4vjjl9AbJ88jvdZMnPmlixJP0wEzuTWxDukb8U6lmdPyAfI/JvvCF9m7fYWFF
wvTYWZFMPw/qMHbjIEo+bj/guzvMiOfF4wngbGe1LabKj/8RR3mGw5k3BThTxiMx
VDBsGLzrZaXW5m4lqi3DJ2cofgyeuDog4aA3j65tmNjlQGMQ1alwVnO5YgYlOpYN
zyLqtkGMp79tQzSotuoKWBy46+ra5aFnruBKrb0EyeQInakqCsOHynAe3WiJpKi5
lG4m0L5+2SN5VxnEV4Aeeh4bL7IstzIMRKfoxWBoPV608HwNCWrNkmYltjYpDyVl
i/pxlyo8LSFkt8CPW2J5MAddugbXc/IB0KjuYv4utrBuHx2f9Od5ma967DBvhWWH
1AgI7mqS2T9oKIYwA+Hkca8h9GUmoHHvz2lSSAT4HGsuczc4qXmJ2c2ln1v06drV
RgKe5LuQd//0LARZ81WFo9zf+ffVBD3UWglN5IEhs3OCJCchbrJrjEZOdzhkLoA8
+inu9Hz/EDtwfkgY1CqOkhDnkPF7Z4WiT7MUc46ygxLoM5PTzoTzzAWIhGB7u+Mc
3natZtx7qEqK2cE1QFYvR/ASQSwaioIRu6Q7Zd+3Xe+A74YivfIqsRAPYajSCpy/
qCbq5TPOCx49Eyt5M/pkCsr0Su1pBpueFOq6YAIvmnm8fcljKhkdiSWWLGjWb/Xv
PnPNEvvaBK3T6fhHDJFgbYl4EsGpSCHzwc1sakqyM/t05/ndDCPi6X9XZ101nIUP
sTYbOYaqGNjIDQbRJyZnZFDetwPh+UfFHKslNcoyC7SsnluHzVulg0mf/vdzem/Z
IhGam0GXiSfhFFHmrl9c26MncQarMeS8z+pvaoqancaYwXPq2qFE7jhkbYmVBDVV
+AU5YesgbbLUZQoYeXK/f5uNo/mdvZcJVY6mttSb6vtJoO5PcBUFegUdzgVFL4q5
WdI+eiAAHhP4ZL7qk04GunkQZyyXHjZcFDdlS1jhsZMGDUoo2C1T6uWU3II+HmsS
gRDR7O7rYoQdEW/BwGuucmtRUA4g+5WXuHjcLE2SPuixtRXdiNyQKcrViJyt5+vb
dGT2+fA6BYbiEHhXYmDMeGa4t6GqLhRYkH4G7gG1fCTlLCAGHO0C1TnDHwnAQa1L
S5GtAJjJTNq3Ys430LDYMA3fAJ2suSAtZ3DBZb88bbUpvAEdamje1doEDnFyJIU1
Eos9Nqcuh1CfVv5FGEWqgznOh0wt01dy0K4a6qgJSygB6zUWgnNPF/+RKW9w7Nqg
68zADRDaj6+Ypo5LTlJIHzQ6gHvSei3/3MQjh3GD0RsGHrUkq2p6W9bhd+qov9Z3
tOCeaqxXKVVpDc0k1x+oFflZovwwkG+7Hf4b1QvyFbgxjbWJ3s4PFj3MFaLuaac/
7wnOZn1Oaq2rKEbfkx+aV6zUWAhUKqZmAQD9u0sSKQfHmg9iiKliedzwKM79sXtc
i+zleAv6sDhFTTKKJ/JyziGOushNGO+e6BMwBDgjGPDJ1pm/887ZaU8RBgLjf2uc
g+IlARqWJ0wHKzM5KF4+WgDREl1wFjHBIbAmlFTw60wEaPHARa8urRJd96j6m28Y
hXqKoUTeHOWA5Tv5815tlXJ2skoe61+vIw9SwUuaJzDIeO98CXbVutFFzu4L8rn+
visehQvZ5x+SsEyyfgnbDBiV7pThiXgJIbwr11H+uTcOdRhQuCUl/NDpL0dTPxbC
b4aHvPvL2zh3Hj1VQFzaMbjisR5CHodmheiyPIV+S/QKws0szAh/rsAl1eTHeHvE
/Aiey5QQpuZTYqHwsAwY2Wb5ITCvhDuR8qbMDl9vRUdKRSdnu9XcAna1yPlNco85
6B6/j7+ssf/ig7Fkfj00Va+ImWOUCBDMVAEzH9oWPMn9Z1D11+4acT1BW5jbqrGH
xfLu+cuxf/H5mSgWmZE6QsPVKG+HdrpEb/5XgrwktVeA0+WmgjXDLiPudnk/obo0
XTv4i8bX9yGeHODkdwSUnaXXPNPXaxvl9uoIBU3y9L7VhmFIloY4Kug2/5MP/VIM
sYMtSlArROv2VY2+uupM1LybQzg950y9G+/Ju2Zw3gOuXJ8MyRMp0Bsyf68/I+t6
ZCBIhiZCuqg/Xbb162dCl3SWYuexMjUojZCNsoGTAHGQQuxZ+mDrg1os8tyYEIKM
BRk8vsoq+b6AO+lEdeCi/Brab33JgnVDZWo+58TtrUVVUo8YUWlj8imkDbalhtbC
rKKLpmSePfrRNscK37ofbqyVrcRS5bkJTMhhNYa6MbbJIwnSbdqsvB/yClTiEn/N
MkdVp+fQswyZlHHUhN09nnMlZ6uX4h5W8FjjfP9YFsrxLRK0jqEgRuy6hjiX+Yk8
fLFrayY4MbIgm1GWgHSDi4IzxPuE1YjdWVwzPkA3KIDZCaQmU2B8E8X9RpSxrXTL
SguHVET9TyIXChkvUBhrRFFLqXq2HK2/v/F4oCTYoTS+LR4h2ijRtu2ai/aujJPl
DDQI4IZvo6QBNWck0A0EoW+eecuyB1GFMDMLfZSo4jwFSgYy7LFZ8qG0s9KScsDQ
Y77C9NEyaAcbDInjk4l9uR6koQINRtdYevNy/RRjxu0Y8JRpr4dxvJ/OrRil6ohZ
aJzjRnz+maCDKeyC+ORIMysLpeIwVjnYLF4ond34qcX83enjcTc7KIgrW6VM4/g2
DmtemrDaI+A/i8xKZMN6/O+BQZBkUmje9D53jong7yAAfZxIYuVS6OU4BcPOcVgI
URBFtsm2O2Nd/x8Pvuq3nc5Z6qW2VJltX6G5po3lHL9l2w7yKG0XFNv6zMDpYjfG
W+u1dfxrv8xgscx6Nvxu6esUA8v3DxZUPl8qpBf+A+dQmN3S7OtslPrV8CJpRQhm
jxQmZzKewmdWOZSpJTOjVbAbdztUcODZv8KtrE2OFr/VxBEAHnrIyJyXwvWVDd2s
yim7EMFZXBjlPFicQG7Me0afK26UDxgjnWV59W25avBv6MEr6+9Tabd5KysZJpt0
hauDPU4gnYSnTRuZWsBk3tzQh91dg1/i9/kZ+14Wg/eDf3NIrkZhpTW4MaWgkT4R
EXYOOf6F+8rG2oznhHLSXKOGdgfPxdhXFAeJUXe6DKKew/VQ4T4ZvTFHKrXm5ZL/
GMKT0ZKqfDRZgU2O0rFVzCV7fEFo2A5kag/oKgBaq/DyFJ4Spd8kH2+pleXqslt1
MjdBzsOU6mdrqzv2PUYx4DW2JDNKGDQpq6B8vHAovMEEtvNGfTuaUy74/viFwVoo
49erPUp/pOPLrtIFmzJHnfuHNUFtK2tG4iXSS4mEzo4gDS/F7aQIWBakOzmP8GFT
PxRfwhLTtk6U4ai1ceuwX5pKVV+3M/3mzqGDx66Q4qBrxbQPwAohWQ95ZpvHKxlI
VZ03yO4I5TcLxM1MkaOIvPyVhBYxcCMm24565kJeY5JCb47yjxx6Eug/rqh89iKT
qIEbVTaCJFjbUGyg9KAPN4s3FmuS4UU1kSHItFF8HN3BczM8KrFLoRw5LLgYSBWR
k8ul6RsCymOb5CEXmGisQKW1qSt/FkwgsAwYnHNxtEQmvlDpNxysoKDszPI1IMl7
Dq42MjtUg2xWC3HyeDvj0K+NfeoVZUrN++/nLu19lp5CxeZxzdk2xaRysisJr/YU
ayxWK11ocL5zCJWt3lYAerHbf0FwXH8p1/yJeHSp4+bM6bE6fGq0DW766FTBh+e5
4QCaH3tAnC6ffFkcdugjJoRWFLCO+cqak6/5gHst5bOciYr1p5Sus9bZfErGCQv0
SXiEWG/QrkV3CJOeVJaPziyIT6ch0Bmj36TInr3Z/cHwOkGIXlmCtdKr6290jFjN
dcCGGka8LeTYDwbqzI9MOPzHZTfA24eFbH17XlmJ2qKuwrS9ohEeP3EtNiSdnVwh
P86Si1VUIwO7zCOV8eb4KtQ63HeT1Q9DkcqMdlVrtNHFa1J780tRq4HzYhYPdxJM
UhFD17/lbUK+4KsTqhErQ+PZr+QhDRVhbxfvXGDUiLF8ycS9e/WZib9fb57n6GtL
EOBwhUW/Ho0teee7NV/tCmcp4RaGn5Q0ZQuqIYH8uWzdz7Pbk+Zfm12ScNcV9UuW
1DQ+qEYSLXKAdsfj8jRBeM2jSp8/HQ8M/9UUEvS3ZdOUe9c045hBe/q8MmZQlT3y
QkSJWGmKN9Xmi77X9xg9qb3HM3cxqr2Zfcb8wMJhZXXUCCkQVAYnM6ED293Ly6xb
iNeN4PcqjLQN3H2gZgEAMPsXpRk6E8n9NeLay2yXanU/1WM/yCIfDimZuwagB+yg
flwe/UFie/HpumIQ3HQJBOlMx502Fmh8esUjoSx0lvgrGKyDFMQQ0VzmOwLE9Mj7
ewO1vufhxAy5sHFKyhYWblrEN3+/9uCAzyB41p5xSKP0xdvff8jMFhReCQ4zZuif
D9KWXG9F23Q2imjfNqWjsjlzOBAhAmEWTQ9NdkQ/No77AHFmBvodIcHowKJh+tG0
dk+tqKakGgBp0N17On5c5nzGopGBFLm9Sq7AMBlKUzhoZ7MYHwG570GBJtpahcfF
j/dHjqP7b1C3MtXuaQWWLYrfHMNNI2WAEq+YMXoAgPodueYciNJUDItT+YByelAP
UTt152v5PI1mT0w2Noqs/L5vL/LdEO8xCY/s/8rSIMR11YTMYbFMjHIVZaXT+qah
LRR2PWYefIXWe/+/DbpYLJeW9I5SPSBymyr6gJkIrFULbLM7TJYjP9Lr18v3ww6l
lTkZrv8Kch5bu5hO8ZfkQ3Cp9iOGGKZfvjI8Jcl2uPaJDFGOGKvnjPgDO0O1s9zF
T4QxZtypEDLrYJ7WRdGmkYRkxM8K4OWZnWGCeL76dyAnu/sCaaeUjUjRljshx6Fi
uWURYXCbxz6vupA1Ux4Dah2oLkOkJqdbGZgovyJlyOsYIKpPpTTcyOu98hKhvYd1
GAxa9XBPkNkItp5MTcNBk3oXm/EgBKM4r5zDi8aNTbdQTqc9fCldGhuH12COhMQa
gxVNk+AtRh79djKgNH/MMrVZCeZhP0Kivhq8RYDpoaqvvdfUpiYHTUe0GxRQ9Xqe
PG7WETNd0N/+Nixi38ljF6HIgDEiRgp9v9CA7q7jjXUeJc7Er6Jf1u+gqqJVlC3i
AJ//T6weGZMnvteWFKVysVmAtjOO5qdT0/JS+LCaGThJ+0X2aR9FHeUZXHMONeJp
MQwMSyO0U4kQimg/BqsakNAZYF357AcfV6vEHXF0fynWhdfJ2VUeN7y6R+rLJAZd
HaRNYZ5mIc2pBiXODlOTXejn8UvC+R9n3qPMKsykiErVWK2rbiWSH1SWA91Blxg0
+ujY8t4tfhjQOyFCbBXrDnFU7GPCPtxae0+6b6nvfQTTA900PKriE5fD2AyHp7pB
Y2E7zt27iLM2BWtYIFvcJzZ6eVvJhu+oZFsbzePu2Sx9vN6Y+bDNnvNFbh45acx1
8gv2glQkAEqmCeVcZ+co/xZLgNw3Tx0RgKjaEfkQOHJAeOmHKAkGAfMmR1THvFwo
cUB6Ku7IbKbZHTNElaBYRVQgei2LEMlOPocPzV73dZd1p5nYJm4zORmje5h6PLD8
YVycnLfGwWfYuJ8zJ/BfDwGy0PNMiNfiYheVHeV0B/rKjnZpCVZl8xvJJBiMiQta
99AQcfXqIaMUKR1aK7sTxOeYY8u5NMLzBFL04kuqZuEbSTGizd+MvxXq80Aq6D0S
oSeAmRUrIBMKkL+Sl4J8rZ4Kk9m0CPo490AhHpyxzgckYrmFNal0N5b/US6zlGX2
kcd/BDYNypjJA2kmXZTJ0KBLRqNObQZ5kNN9iCTbes7T/osZfoNR2z4TyaO+QLCx
+qd9+IqNbaQph9/QpnjUHzIQePNV0L9r3O/zttBd8+G//Clmtkiw5JOAWs2uaZAJ
jgPmjvzo7sdnn7W53BmF6VOZXwFA2MYiTUgKLIIjHSHE0i7mvEjtNEFKUH7bFVEd
py1ZSLlJ4Qsz8czJX4G0oaQyYzMoVeEyUat0JKI5kZetonh1yOTEBW+3K6FG/M1P
VtQcFYt6Apux1XeAj0+wvmKeYVNUxEAiXD90aAPg32f4dL+oGfJtsZDvXv0GzKEI
DMEE225yf8F19/3MpPpOP4jHUoJ6oRpaT00ElUS8VG8x6WBzIcaxlz1XhDsHfZJq
Vl6QckGetyJLxWfOnTcIb0iXHQa//c6TGqnYJzhfxm43d+hK4US5aV4wK+woWOiM
l64EvEx9O3ldycFPa8VDz0rKIQt8S+VYiWMIRJJJYe1dsPWBATkUjvVfLDrOUrev
0qjPC4ZaZFDnYRS0zYZlKbIe39YZ3J4uZYDie9IywWPR9cFcDmQCIIaZVAeQDFDL
jYqFY+jnMoKKmA22TjEjPKtOh8PSLJMZTACyKo6EfBDZUTELBururqDUIj3qY9yS
P0WVKu0VNCS2DQv7amb4lE9AClko9b91gzGeYm+nkJtFzitbxT9aiXOuBIe6Nxyd
wd9pcVxfb7cYugzY7po7PJ0Sf8+L6+1j//wg+Hj/MAfTiozE7OcynHsVev4xS8o6
A1Wz96UpwsMoDV8hdb9UxWOmHGqaFXNmtr82i7OUsK0xOxZZZd09Yuo/Hd4Z+8nC
l9TigpDsx3+tbazIPAmT4x0zapUNj3ygeAFCIuVlgmwofXk8qX41W49ln8Kcef2q
S3e+znQ9826yWol6OrMTVk+Rycga0wWMAvYtbaeRnC1o6AayXZ72jxuy8qBQL6eM
+VFmHSprpG9EHKk5bipGfZJDLBlB9nVJFdJRTTD4GtmX89oV5w+CTqqYIA8mDbu2
+mf7xdbipP12O+PFYHsqzArBmBWzRP6USGsuKBRcsvhGR01rnhbYlGzHGYQRzoaq
npJ/NSxfpT9DD0Ml4+Tctgt8Mb57zmBJ+5miTZ7BVox/f2RMbLh81BD0oEOKf70j
pwSKXyQE+WEbHHzJ9fFj+UY46uvXT37Hypr4eAZggGVchcHs8lzjnjisOCWsJ4Be
WxyzqoOpKZ6OH6FE5/ArO6esh3YnTk39ZDzFioAsTfvnJGXVx0BHjOMMXiWORZJN
zx8lINeamJHx5cpZE73aFxE3DgypbKgT5dli6LBjL537kpn+UJQ/ManuofS79JKX
WKffIW0A63xHzvDIvAm6v57X4dBPrQzVijJHdOngnhJlRbbLtzd+xweDh+Q7Sguv
9iutzMEsoFoaT8k2ffGZ0kVxDoz6blzqT8x3AqRpB3Cv4bzWqPKtVfVOblJYng99
HlOLcWXqeasF8au8zpNweEl2YQ/F0MFKZ/a/Zr36DiPmCvw90CYo9lcQCqc+yoOE
7sqMrnX+OOPG30ewHBQjVFJhL55sV9DEI/SLkpHef/qMvgxYMRYFOjJ28FMlXP67
u/ynrTtgWwPgCvkBq4XQluTrxns6zHxX2YHBECXzrW7QYVxR04r2GyBYY1Dzx30l
m3YHpdu5pwsBJCqQCvFTlL34Wfg+f4ulmDbj0yeIfnYvEgoISPHWx1IWYsD1CjAM
LXQdwRV8L1q/AnLsGyAh0042npeYn7V0Up+/tzQVHqWX0/vtYPCT2eJD4d9jFOSx
BfY2HcMskcjqCUIzA7jG32Blrg55uSkcblAQ620ml3OOb8IbFvBgHFtEY+yzD71n
prlLlKeYJAdXSr2wZYMccIjUp9WE8sHdFzPu/UB3DkwWmnDviiO4CCBTs48AdRfU
mUO9jZT6scLL47SPx5fKvJuvy6Pa+BI2UcDOf5kaKm66OPGmKf9nHxlzplNMctfj
5DD0kb9AfjpMiMX4HD/kM2gifJsI50st1yhHW50UOR7hz+CE3pVsr13u7QfBBWac
JUYqN5xqCWwwV9jSJcUQ8cWS1Xd7ReekCdBzHi9UgEiU0WyAv9n19dvTuxvqnjyJ
h1FWxQ9p+hIS++wZQdH88QwI3V7ntTUbeVzsfdFhAAoPaeErwu8kuOXs8BIRR90Y
wpm4788NyvfvGfLJRYIsXjp2phoxbYXtU8OcACgvA0fDdbrA8FJyLTCkTQV8oTiB
r0p12Jjn5yiQFqFynaYcjc06td2wPRtJ6TGEjuXI+mWaW6XrMZecxC2CFNbwTa72
hhxpLSA2vhliq9TkcualYkkHAsj8AY/nqBZV/golUEGLrOoaXsWAS2nqjTckViX7
Efw40UbUWEni+RQVHwTKXXcGVeffbaVNc1MTHunuIatNPbS0yIK7fBJlpt/y2M5Z
uXep5t/Phy4wmT7gjQby1AQKJbq4QVZvZ4+Kv6gafxahoNinGrlGJOQkv8rVNyTo
a1C2nN2hieJwGpQBXzIUdhxUDUkZb50jhe+oDos/HIWaKtOtkU1FMRwSXI/MG3mH
dMxdkaVYkD3HtcgcLNvPzZlbT3n/oR4ZbQ8vtr9O3GEvaA+y3Kp1EeLwYxgz81rT
nOsQIZFDrHrjkmWqPtQRX4oExjIeawBNO3P/7k/CFB7C5qYyJgwFziLaA1dCn94b
5tolySl5yPv+LV4XJkcKwG5R5pVb98RgigpKx4eyRrPYSRtWXtUosO8JIFu/5dk9
Ff8XLxEWZwih756kik2/VjA7SXozHKVA0ZN8K2Zzi+vMSmah+zoOgH4NTdHDw+X/
lnxsVTR/Ci4UdVrjrFVt/jgkMwiup0YQdyuhm6PZNXGcaEkTgi14Sum1a5Q8+hRl
8WRYvG8OmUcoozuGUkVwwMLUuyP8wQaCpnamgmj14FYAizlksIUNr0lhWuVh2Pyn
8I2yp89xwp5mRafAI6DMQAno9Zd3v0BHqDyEAsDfODPPli+7+JJdlYvS4j6Qxtkv
CU24ezfHDm9qzqhQPF/PoOjsGMU+t0IGGyRNxex5HYPrunjTDpuC8o9MSigPPqXf
asFfXD3HLeHjQ8zHBsUbN6OF+wZfTs+FpRTlwWeStwdwuQsTN2SzlBauk1HX+EgH
7a5f2gmcC5bAU9UAlEV3OC1/xOORei2AYWMxXYCcfmqLPi4VAruB6ZEMBW1hSkwb
vQ84weMGXrvDP0lWiJqE68bNV1c5Kmy95c9GbN1CUXfKUaqFlROUOPNWxsLquz1L
eakp9dq0M2UmQo2gf5r3rBjKLixoa+iG/ACF0hccpSL+aYb7KcqD9RiZrgFSEYBR
LolWxBME935FickvsPYc9Hih0SL1ZaaWzawOC77/2oUQQo0QJzZgLhfg8D78tip9
6eeektIiDmxC9VFtpXa7ZnW3lPodAyAgoLRw3mXgnPJ0631l/OAFP3Rp5woYvDFH
dP1XIkjC6QcH1A/qIPGSTnBy4ylXwsU4MFqpmlf026ZC+/bsVkqNOPnF+8p412Pb
cGki2zQv1Yl/LTf/j6TiGiXvw5SkBzL9YAYwjvZZGVBLCoYoH932pNeIQAuTsxv1
uJodHicq94+cPTjfg/U2nutfO0mDAMn2VXSBXbQUhCtCNUtGJIR3HzUipGtk4Pix
L6gV3kes1MtwkVcSKFr3sKhVf+Pf3a+cpwSgXpriLFVkzsQqqMneOUqlMVyYbFjV
/fgrOWktHS/PzlzT0gz9elt2UDGj7iuwmltJ4wIE5m5OjtgxXhR5i9LYcq5PjucZ
MwERJ9LUYW/BVzC3SDyGMIZXcssx7q1pw2cAR3J3C1v66s1lr8O/jzd74i0Eubim
apMHjCOsC7/l+VHD2rX6+A5Yul2im3bNJAkaD5Ww88LhJ1H+PQYH30CK7tb6XnfK
LVf1nM/JF+J1yzJJVbE2X6uI+daUUSNb3vs2MtVA/5/xuf+GZBHFYzMFJ47M9UYy
gjn32P2UQ7Tn0CA0Xfg/NSrHvQYbtZl11KIC4dSMeo2b9nFQMP12dRMjQ5bD2BSm
UvYwEzKkRoVqfUUEGZQQnjdr13r07uwqWw7kpapoM99DhUdaO5FJS9OEiQG0jucd
cVZP/fO1BX31NUircoERJmNFc+PcM1g1auLLtMahA1lpc79li9+hyZYiFE7MTQ88
8jwHXgMbuxBk31U1v+xiIFCyltra4bQiNPX8QlvFH4I1qV3fUdOBKibAGnmnfgnL
PIij8DF5NuOfKCeGVb5GFjCASyKM5PMrt+DpW+Vrq5WhlI1GC3UfUPW/R4XT6vSK
sv7wL1QzsFPFolwIoXjJjxku/T2f8fl4IUX691zOPvGUFmPzg7xE3lLJMzHWYZfJ
mH8S+qcjCWXDiLa/bWeHWEwQf8pHFkslHa7vgEOjOmKBcqG0/fqP2oLfYKRHIrG9
g3p8AXM9IE03NRsJ7dmaaUNqwjzeDcj59qRs9hP8TksDla5YMF8acnuxggkweiPD
TcYtCWHpl3dNVgYgnNPZQRpn8bpXtL0wCGW3cLEqf/DDWaZUcnTrlRXyD0ZMjFGK
XlDEV4j/D7LsviAcejWHuBxqmRkUxR1TyWmFabAzehhHMO00WfO11DwBGMg6HrFz
Oddprsl3bpETeUonZVrom2ltmn26Bw1L6Ngk9S2t+7/3zxEx8GEtlOGoyZAFSs02
etjRa/a85Mz55ZZcknbP7pDmBlZ7rAtYhEoQJkpoDdVvoN2WOy3NhDXQ0jbMfHJi
GqR18qSw+zGB2y2DZrF2NDoKnlMU1DoZPttauZ1Ftllm6s/PpuBrY7/69Op0zD6k
cVdlYKIo3wZHI0hMcmHTcP/4GicN5CKbc2FWqG0L44PFZ+wbokN3G16Y2kaE86oR
K4jRj3UwpZFfc20zd2MpIGqEcgaGuc1vb693uYC9xV3LygECsAm85aDNhIWsFvWE
jndPA0tidcq26l+l3Vkge+HTuVswEDuou5b3N3OdyDZTSdT0cHMRtMHrQ8bhG/Cr
0LOzB64cYFCDMVkNn+dUte4Spgn0Ug6Tfdi6B7HLtQn4yCEONFx/oDbm/BN7+DfP
TH3EkxdT324zFuNAya3J/EaZ465fPV+BjqYe0cTe42jfB3f7rsDvx3vJ78GrpEIV
azRZyjZhmu16A7CmLEGk0ADvszpAv29k5GE8NGG+RHKc9A1fEM8r5lF0I2hMlw1h
rrwgT63GVz+LMwX9NP5WpO+3mynaa9GEzasv1AzwvDP+KOlZ/snfAgvAD4ptJB6K
+Zd3ksN6H3+FTMsyc8XNgFhW7jIJNGzqIDffS2FcVhNPGJuS67Oysm0eS+Hoqjwm
jH/8OJiFUujZM6loQlUBep3WxQz0NTal3c45zEEEdJ3EiDS8QjvFxBAvLG7PuT2U
X//rg0gAupehZAKJdlSrd5bCRbPPpDMX6qoFrxyU+FQuoztmPjY2M4twb8V0QzyS
+I/rRMDQrohwBEkNc+Dgknsr4NmBDSNNbmKSKY785031L6v65lyn1/QqnBYOyBCN
X+KVtyqlYjU3mFmFy1UkQx1Ceh/gYjZGftBbbLqgBw7jzlNvI7CdTvrzQCrSJ5qu
GxscOy/eCHMhLaZ0+7ORAptGOdyNLlm1z6XdVp9Em9TQ79Qxre2ij4qVOP+aTcqw
utl3mH+T7AjDj08JTqi74fPjU8dte7EbYp6xS7pfQJgJou3Q0lShB+4NoAerFo7r
AbXLeBi34fKRvHijFtlt5Ygw00n4ndz6ACNCjo8D+vvPtGhbfLDPu3PwppxVTfo2
+Pr2wsyuZ4+dcelM6EQxYEexVnLz3V3F/WwP2TUlrQGKRD8QAi9hqRdaHJieAbqY
9Wt/HH+0lcRCVbVq8A+J97ayAewhyPgPCFW1aagXX88lk22xgJ1uzJ/p5zkwtH/T
nFVzrc/U3m+4pyVTXsZanvHOMuqTcco9yuSsZgznsNx+9tieLht9OdYyeEHuzIpr
3JxOm0LziFeNpLh8KyH/t4WNH2EpcHZL+LkrnGZBdudrf9/L5FJwfitfuC6ERnwW
7MFkNz2xFAIeN9j7CHbmToFol5iZHGw14M5gCiTx6maYy35c791iKjMeWB8q4r8T
+1zeslVf3AwSx2NUo0azOQpcraajQsA2r4QsLVj3RYQ4aMBoeZC2Y+Yt9JolvuIJ
eRc1V+4qOhZl78JobWD0qNe0jZNJObsZJfThEDzN7jqslF/ZTwqHSySei7E1XP60
LHFUMbRLbVVyjYZw0nS1yCatl31T3QpksrPweo8VUW3am6f+PcjT/qUS8OMezkgO
uRnEZjnNo4Kve7iexIKXCrRfgqHHvr56eJ3Zc4WF6ME6oxc/uMUSVrMQiJ2hlv2H
GFu1PVZiLRoS5veJoshEJmEnpe8BTDlnIweQzWnyoSgthBcEzcgBMpNdqgC2ltJz
xueM4jPdpu4mOOsfi4vT54KGy6UBrgckbkXfattgP346UX2jEB23GK6t4RpcntDW
CfxKU9qj0HaMBXq+ceKU4S+Mi05deld+5b5A+bEozAIDWiN8VNNcOZB7BGHAkDFj
P39h5RoUpTlIDN/7Y9g/Vi6jiStkjNGVzcvSZ0dDQ2J+IdH1EztxnFQQDqtsk6ii
R85rNyxAXdTcuZEOT9XI3+WYHSII5oIZTOTrOgaAuZfGpWDCgn/gC5cxbWkaN5IN
iec0rnL45i8U0H1QjL1/a1OGIgefOPjK15ztWbqACjOE+qvcQKBITUzWwI02IPlP
23MRmfUBX9uBupagcCUZmeOv1uyfj6mXyP3fca3EfDTyvRG/G88MIGJICNbW/2G1
1ZiFcvb6aJVfRcmnXZiB0r1OS/M3dcmJr9htxU5YwFrEVtlluxxbrCvqordF1HjW
XYbdaiMBUnq3Q0E8s5v38ulifJKAbwecL+EgqXfx91y+h8ajMzAC3f+n+6G76fpR
P6Kny4SZjNRna9ivkZADHnoF42/xKiIAYoEgh4880jYI0D4A+6wBVRYNpCaQE/po
+QGdCugis7kLFTEZQ1EzK/7RNqmRSvsKG6wu1YNFEcWw1dOrLbZCuaOlMPvR09LR
u5SRWeaxcDnf88eN8bMLSw03sGUB3FcIIt4dU6I4HofGwkZ0T18dMC5EQEkaORlk
kSN7L7CPGAC3gtOm5wz9iL46Hf9fHcRxxKytCV0QxWKj3CReeIozb/HYDjmqdwkv
ChANv7gN49vsc5DCj18RxZCYZv7UHBO6ClLDVQCm/Yrd/TP68bMGp6KtEGWmpUps
A8yjYQ3pTtAOUQxmInUHUAIFtyG6BHhCKmJeRK3dyD5mCepomOvc1mhnXMgSqqI/
tGnb3ZkiK4U/4sMi7XYo6LdBqrm0lOIZdM3LQlsfsX0n45/inL9cK1WjlmSHagOV
owOy2sAUsmwtdzS+O7MOaZifIWpjEhUyqVC6MmRkf1CwaIUwvGN1IudI/iRgBrgx
5yta5ECPwc0mmTp7gGaiA+kMeWYTeiprkwPew/pfGttX6hczrHx+7/sjXishNJDz
Mjo+LTI3bM6tgR+y/SnLvuDe56+6JRJnUlwMJRL+Js6amjVSN/lxZZ0ED4y1gimS
EDI7H16FRFfqpO67lwyFfpX/1F4gFo8eRsoqRuH8xbzHKhOM7U5R5mvNZaWgBape
PLmpwf4CMBuiNb4DAz1uUi1gInsYpFa3PjV8UtHOwlVt6bqaVpys60thNZv7xc3b
8y2xwu8J6hEbzjoGvuHNH3/53kA+Yam85MGILNLDgO3l2dsnm193hg+bAnvWe9MX
hEOAADcc/0rr9nVf4iwsiGI3R2zwCJgT9RsX2pc3NbmmKI/Jmrn6/PEcAncjOCVU
hStLe9SFqSb/MkpXFc8jSBi6+jumhChnjUlvcjyBxz97gF+x8VBR4bQEHCYMdxPW
PmTY0rpbW9n0c3K5moUQv/V7KXblL/pj8lrvt+xBV7WxM59n2LgAPBtygcn0UuXx
gLX8bgzBrTgRW3VOSMO5N+LXrocLUHuq8rADC/jTzyhUdyqsBgJBiDJPExmMXVIQ
ukxNXrK8SBt4OtMymqLvxncS5nPYTV/Uk2yVgOTSWGaB9BuaaoSv9yR1YZhw14Zf
8uwyMtop+ZOOCNVDY+9Wkg0t0le6OyllD+kjqLKsQ0ngESUWzPw2N/d82Vzz3XsQ
SKoqIO9ogmwrl6IjUBL6/ZfU3334QibqdEalaktkZkXoLO5EVMA5vgEODx+0Oos+
4ujujhYGB36QHP8DbwggCpLIQkg9fyWAS6nh5MydBRdkp6CK6EeI0H6abLfFDbhO
0SnS/cfy7ZjaQb9Z+NcLnhIjhCkYEbm9BExKVxqFzr9hGMhyJ0mGdMebqd31A1Yp
AIvWisQtLZuMRq7YkUBQnxuQ/hRCB/8EsjWYug/4qT78AHU4MNYoaKs2kxCO+zr7
F1h8rs0uaTrT4h3AZMVnBe/8OKSLJeHLFFDQOYgItIUSwh6Yi2+OPC3RkCamuvnS
9lTDeMz1b7/w/YUoXtf1sh8v/dufuhFfwEy7Ipn+dWFLQ2CA0eWfKCem9hg79r4b
6Qmi2jMYGiYm/6dqeNFw55SspU5Lc6nPme4TrSA2zUl5cBNYEmog5e+LG/2IFMqN
RDjBy/+TA7RBxWv6mDQkYw47WQDZVpcv3JRNR32dbm6Hy/a1NwIyxJgz1toWFqob
UDsGfitlqn+7gUV9VMZTy1N7oTv/IFVv4mUuSoWV2dYRLY6A6WOkaiY47vQZuiyz
Cx3S7lRhNqUpfQ0TXF2lK/SAHoYmwcTNDticBn1UxApNyjJ8nlp5ooJwFQd4AxDi
KL3fO3C+Z2r7TpLGYto2NBe2nwp0KeaIvGvxZ3n4qEwCjWWX29WbH4ogNTC2PLeK
wlZQgiJT0vjIGgBLMt8RzHtaxN+2Sfpq1Jn6OojMG0wTpcx9QPkg5BKNSOgZTMll
y+TVTW/wYh9V4RkhyhjMawBLZrzI3cVuiTIE6b1kFvVmE2AUgXT2aNeZ29C12PPc
VvZeI/03r9hiZ0Jnm0Id7HRrPoUpf3EgxcyArUDkhBT8/86OnovaZ9Mb+bn2ffXq
coUbCrinZS2HISq7uWlLyjEdl+274jaVjB+exyWufANpL44xYC6kNJbtTRG6dZ0C
/DEZJp27jetoJwRUZjwgEp4VYpZCqoGCGQ8W7gThQrUITG7P+jlxqSqGSdN+ICc0
MI4yyCD1udHsdF7PBUGJFOPyykwc4PmODK77Q4KW8mhANaDvgeYwacJTMfL9hV4D
RmNKgRo80soI5bmQVOeOtUSzpBDgbHukm1K1hQrCPX5lLuilj/ng3ejoIkLzP8qx
uxa0alPiEIfYHuc15oqBS8163eTRvxQI3TQR+wd9tgPJknoFYY42MpjsnC5YJiVH
pAI7VtpntgfYnQwnMpvkB4RvXS4j4oMY5YXp8opRSNZ+CDSwKbuUQNovDrDx/r3W
2DcuZiyaLp8uYdeTNurULejjg8AvupeRCOegmlh8nN0x/Nr4Y6sJpkTwevWEB+XK
WobGZWMOXPkOGtMMt9DUbLVA+nXJCSyMpWlfkmkfzdrAVcaIfrZlCafZz4JwY96V
RDsnFN9lGXUC8JueQS7/WF3iCyVReAqZ2a3GnnrbT8dHyoV2t98YAdPAZcS/GnQQ
gcmHkeWb+cvIUZPqJLN32OHhgVZ4+n5FMb7JZPrXc3gkykPukbLE0/DBaS4r/Ozj
xnoYYWDWM8xKFE9aSq3siEUQENB0EF/jLW2JRZdMU0n6P86m4e0MpppxQXSvria4
v100icYgLW4IjPVlk3jJiJhOgXzGWHAU08mCxkcAGl2xLh1wmBxnF2I0UXk7s7Fa
P1ujCtta6CQsB+VWIqGNfZOsduIRcO1+57eZtAXb39Hm0L2XCEb+ABZjql/cSsi9
Qh6siLrkaRBZzZF9/CwvyPFjoKyKfXqeMj1hdtDRwvfaM1+I6q8AkuQIHJnlCa5V
CzjtNZyeL0aFDVDsGF7li+kjaIZh5qjTRcVNBpNCcGG0SXAStX7ZExmn+JYeAPNg
h1e9NhFgIjI3FfTewxm4z1HjtFIFFxEdtjwICESzY5UTBAH8HG7aQ89wP/SiVgv0
bhVP/eFlOvMmwmirekfoijxG15G0M7CSV63mIJUlHe9J1kYmE67pd3JW/gJ0TKnF
YE0/D/4pdQVB75nTWaVFn8i+1Kfd4gYWdedgu1L3kJwbBUNUWhkvUaS/R0NMW8NY
V44L6SS/r7xaXQ+CauLgj6IIgCCPzd+86Xtn/9ysklgqPdGhaKvbuktR4IvKNUYS
4WgLd2cPw3ZDwkyuEA7AJpWF35Ao45iPpXYmndG/1HjX0vnYh22KhxOZz8Gby+87
LeviOCrwtzeA6H2N8Y50oulpjzaI5CpHHO5XQdsSFceJ75JDDYWvThLPeVlq+3Pg
treSSlaAXcr/16Xc47Z30dEuzDn6d48PLfH5J9jeAe7wHZaWKNdRRaQj/00YZyZX
ue1/eTdD98R68KaHwHSdY314IvKdjGtnFpe4B/bd/CfqaWcCU7iFeI6487FWq+Jm
NuzCC/snS53X/6le7x7J99A+KYilCsrMVILuUcE6xVLftTH7vbYRtFio2k0R8QY+
gaO6K4UzfqQoqh4Hf2B3ERAlDuKW/unaZDihiOL8FL0h23imOKP9s6Ij9Ah9tqN2
rpZF5ENMlTfOeAqSdGjC9T2eXbR9BL3MHsJKa1QpAgII31g961ZVjXCLB8OZqPx3
TsKEryiEXnxNCvUol78gfF/Dompf31i34Hnt6SwmgnAyRYQZUAhhsTMiyoMGsk/t
45BPLQJJfQHs2LrL7hHMR2xBjVxHGTh+x+Cl9KJeY9AITL64jvHI4ChQoj7HoWe2
g5Nv7LycM7kkmbrMhy5OzR0/HxuLLEfqgs9kunlZ3y0i239JnmDesffTeDN1MPKR
AcfrfWEYOYOE7S6d+Cu7pxw7nr2X3kZiJEzluB748mp4FQ5fCo0oYi1xg3CDqJDY
TuRKU/E99LSyEqv1EJLUIVvcQN5h9CscBSZmVwu9/xjdivlY9bIoTkZjOtPttNxI
HjQ1Wgn0a5TbBK2ihigU6PnxXaeRyIXCxkjyJNsmcHu+eJ7SRFwIpFj4p23z2a4m
mvxPK+LANlj3xtuWwP3lf0NBrnsf1N1xLiX14uhUi8TRracYM6bBXvtlo5RObv22
RRIsHu6FnoAGybreDIQtu6x2z1j5Nj4D0AwAI0QWAFdrBye20uK7i6aW6AOQ9tx8
GiVuxnVeFD3A+VUkbM4eoOpIeP8M9411hfYeUYz6AOQZVqJc0kZUCbo5WG7PVbAX
NrfSv58a0d/T9ol3nv1g1wcL0BnU/YlDzsdS3yeO8uFpbXVzrkRqS551By4WDWlP
qW4c33jp0mZoPNYHGN3jfFAMPU3MGPyk1I/TEIVr2HjENtbs3r/H46PhTvfoSplk
K3fgvRsxQPGADnDQnd7+m3ReMbH/n5zoZ9yDzQhWcYcE006ExNHhtb1eR3z3/7t0
F2lt42XRhBG61UAoUJdTACrgA4B7T6wtAYoAtz8TcCA7yGLUjohF4FMZCFipsANA
WhdTnvYuuPlMtmtmgJjF/gouRRtHBy9m8Y3P4uaXtKvoou4Rgm2WgQ8EBeB99ja7
2i3q5SsWTX7UaBCRJjAMcLcvbG6yi3pPPZp+1oYtpu+3trhLT6Y989Gc9WnCxZHW
Iffqy6am2U0SRF1Wo+kaIg/w1DyrLg3kmA7zIsIdeUasmmtAJUkwRKX20hmA18Ig
eYvi3IRP2UsIniJ6yQdf3KzTF3yEvDY4GoNOJZEDjZ+sswXxb6MgQ5E2+ZXchaR+
eIRb9WvhB4KZGkIKqvjuRHfgVFQTjO3KZjOtCDj1M4uU9JMQ1j42J081NsDq3GYE
QXeuqHbgdmiISgDndNqVty//JRNhcR+Ai/aHYhIq5zyQt9SEf56pg8GceEPZjjmS
nWjDEGpeyuuv6/SvSRdjRewcgTGf4zEXyjoF0fkkLfqgRcnYn/y98y5GRSxuMszT
Ny1FJX+y0g0A7awS8bLS0I4/recUiIPE3j7R6PNC7mpUCBJyHL05njL/9tN25jyW
0QD4ojPiOz1vcFnSKETF6KrVt49Jvox1qg9GfHnGOEDFmIbCqv2Bx5j/aLLuJ7Sp
lvH50DlsRUtfE6jxpKSkddTi7aLz3cuo+ABESDPbMPM6yjYAcuMy+BDsPBhZYbPV
S/6GCYyuZ5cIQoqCxigEvCpOl9QgWrKPjex+94yUtueObI9SAV3APi3w8YyanLpS
Jz/x3Cryzw6UGCpWV7Syag0aPyZNiFk8ho0F3CjaVEilKBGt+dn8wilZEU8G5BAO
3zCTFIqDsqgD+DX3jl3lTXGC5FUTyMQbHBFSQMTGKBzQIq+M+aNw6gTXTs0KIcmG
quVhufwiiG1Ito9Q98yKyStjYhqV9jpjDZIiJMRnBbHQwKEdcNdFEiV8+BH1Q26L
c59DHMKV7X34m35ywEYKw24jO83+bJzbGEE86ayUQg0SyeVhifK2M8N/RkBPQAFx
THtVyuk0s3iGD18qcchpxyPVGkLhQkOP4SwLOLzAv14SoeJ+gAb7txs7Sod3y8/x
MW0w4D2C1K6cTZWLjDqGVT4HI4ZFLj7pjOOieExAXWi2JJiu0FshWfgW7IjqCeFb
6poTWWMIfLTkp+Wjf1Ea4uZ+gmaMhr7D8XqG+gNpeCzd/XzuBW7S5BuikmUxzSng
1YwbG2Bq1PLfIpOkpb6kiOkIrVWRQvgmusqX3jOSjJ9bUgxZmP7oCyL8+UlFu4v5
wZi/374EJDSHPNWVC9pu66xpa2VLUQcP0nrtbhHirwIQdpUxgxvH2S9Uv0wT5Cxo
LD+W8EeSxwVZLnozgA+FZ7J+Ri1pJx0rg3jgbhh8lzZyFjsMQQpkIHJAGeKuAU2H
shlpbmPUgdjLgoR/5wqF+KvLkVvyRzECMLymxSHlNrLIJfeWz/+9rK4wYq0s+p98
M11J9hdv2Bn54iRihJ5mtQtDx9I8cwPLJsjCOSCEBtUqypElysSbnDK07j4dGyaj
495v55m1fLsPYO10dRnodswTXR9y2VJqopRVmWfEVW6LyQozytp3F0zkrHY4k5gw
2LVLtL04eu7veJG/w6988N0pM7d54FODG2/6rbTi/qOmojlT/rjIALNBhY0nuZky
vkZgC6LWIT8Qg0OGFz0Go7KfZDdeVEbrWrjP15QQgyD3NVuMdjc+GmrVLGRJUaVC
yL0lBo7otHEWUsQOCcyL2qZaFxwWJe6umWpGtu8gkBYkYzaob5EDWO5ZO/Mby6hz
CT9sl/y9w47YDpKmokDjYpLvQ3z7GXFvVFY+65HncjklnkT7i/jO2LnrUBui85wq
/J4llNkvojWDr0xyrdJ4a8tAW+owxmku+IlY2r6tF5tXsPhsm1kYPxsRC/Mba74u
+69cnhgJxRjgok+cqddf/kXwtNZ/Rtmx4hChEsiAVQjgEMV6DzRkC1xgx2tD98Ld
RmGGeZ7x4GvZAvP/j7yGifUxz/4PhmgCYEv+ikR6PAIr+EdRpIFhf7p4pJ3m1+Te
wma8sWFAwpa8WqeOTOFy4EOPQML2iUxRXg5oEqomRRR3jhYtJ8WMkYZ+Eqpg5X3c
T4rKbfDkMcD5P23aYBLuGaPidsrxCkBTyMtr8gLcfLYSOFPApWTBdyY6WGuMVjr6
NbxWpMr10ZO4WIFVNaM9jj/1bptZvVfkg4e8FS+J78LxxVoeMd+XwqEGPszhjxD/
wLSeYj+1PwsTyLEtW9jVVqwDDjjr0MkBHsnIm6Sh3tzZkecj4BuutjQr3tQSRjCd
6/YrmhodMSc+PJRco7X5oC+CrIPrR1ZTLST/nnZGYQnp6sqbp+G0yqYx0ey9U65n
QmHylRyBYlhPtqdWM2QbJiRz+Wab3GgzARhIreoC12bNL61wTTJ6PLVRlRGEgjzY
SgEMCSnYhGiiFOthwW/I8ZVSIuFrs1BSOQy7JAbrgrAneNyYmEZ8u1NnNo8Zso8y
6liELb7ZrQ9c82ogiSUo9P6RHToT1VPYD99EkSZaRUC9t4EaNxDL8L/0MtbYtRn/
P8ibFg2IcfkBDzHQpRdB3nThxghv4dGMozqwxbZm1zhCxlrlIIFcHm0ixRqQxXrt
7mF2pzHYOzPwaSw8+tS/P4m8F1tx/xnAFemJxQHSOFbV0nngo/bIgw7rhWUgQ/jC
OCpMV9/MDHbNLlcOsq6OA8fQPtYK87rOyC1B83cBFcftpSDrPJ9sWG/KTltx8/0r
qxTcsvZRw2/WgkaVZTSARFaWfGR8mY8DT5mZuo7MrbAB/jnXCX5tdXAjPYGPEL7b
0/GVEYK0yevDxHzDGv2yKMAatJEVFn0Hd1YgmL6gtrRPBRAt8E8EYSoOMb5HlYvt
qtKrVTPjn5VnCnu3rGsJTguMUce0PuST+4KDqtKc9v8Wn4XeSimWDpG0U9iht4lv
MCCb1xcg9rTD059IG8bDoDZaC//q4KuEK/sja+xPpIERiA5JmfyrmiEixMOLuvTk
mSyIxRfgZPwiWyqiR4pP3JC4g1dOQjpFAz2MwqSM6P75rfSzQo73Pd8hzjbuIM7k
qOFX1VES8SW368GWXtH1bqagJR1GUnW1ql6RZM5qekQt5opOcTY41/2+KZ2Prx+Z
q7Dg+mjbuNloyh4toruejL1kaDXIs0tBfqMD6PdFGbw/jn2AmjusetQ+EtGRmBiH
AilECGWuKXDW92hv3WPdP511bvpfT89K69OsXgBgPVgnBrUVauxiqLerGytvNibD
8iQAAs7bjWsh2+WToGD8jJ1QNdjil7Qcoe85LH1/QRNurIODF3iArIkq0DyIXb1O
3nL2AKhAqCNI6vn422rN7lI2aMprGUja8AGsaVzUZTQsVA4gXhmajpSDSCuhsMOw
WcFw75OLRnvSmfDTYRsnXktHlOzHSLHo3pNktGJ575ExEXnRfxuyhLpY6NgitKeX
TIONuhKpDLGerLivEsAFIIB8HotKoRcIhzkTPUzLtw3jxBEJQzQxWwyib5dUZCd7
eGIgme/6LcOiZkiNqJs2GQifjH0GD1TbQH2Uu67SNXWaQ4cKP10vr96+dK/52F48
asiYoR+90jX86cIcxhUtzTUBpSX083XsvrZJcd1jkDkuVc8rd7dOKEK/c6rhrh8s
4WyZLaVRfiwqG/7cumAGNvjqMJu+nDy3TdQy7VTC6haozNchhfObazv2oklpChb4
Ptik7IArP8bfvb0ZFkXugV/ZIeJgBDN33rGRP6obc8opDg2rbKrDnVxJD7Wo/mHZ
Loy/cRi7CPKUlOGtvbQp1wVJgzRm8QqDiYYF0hF6DPzwKCcwXUeL4rJ2Txkjc7XG
DM2c40/cVo8VzAT9zqGCEHW5oTzF9DERoh4vd6XLth8808ZPgyhSKkgOIsBc05bw
9Ntshoja27y8rcr/HUIFI6MmFkWL5gWVTdH8cZgA6b6sVODXPPp+ooo16DbIkPFS
AmUfmZL4uEwMZsJxvm5b9yaQYdf/i0M3KyHv+WW9lIYzhymF7r8VeZm1KurNCmXZ
e5+unsxFEhMmZwuTEu6p6YzewL8ntz5Gj+BTThMD0sYdc+oiDkX3Ojd6nN8eeq92
ZBtjIOqBqHeBJ/zD1tS41h62exLDRcXAC13H2LMClm307TL/o5SNhkG2+gso/Lwy
5DMaH2Tx9b/Vm3Wy8QI28T7uz9L9GoDnAfI9YQeRLrR2BA33UD1E65tmtHHAcGt8
mEvXtAqJtYe3K7VTASuCIdr+NvRiDhqsWJ4GBig8kSvioycir0ciAOX/cPiYTdu/
no83Z4KCzkvknkt4m4I6a2xVx1Uv6qaytL+t/MFTXJVAmn5WElxpVz9g1ZjD+Qzf
/qAAB4A5z/g+2l8hNfFWKLAOPhmupKURYXeGNZee0DUFCDmLD7twdnk9C9Lq5o+p
WhcIFUFqj0oVTYPRHyOjZy/sEO/pBcCI8MIbbVI3HcvKeHtqwvzlaOILYyIrxzjP
jNcIBjz7SaFDnLNVZGtii3z12k/gHZon3ech7AbsPIggKj6HPyMMSqvwn76lvuG/
YI6z2SHtemyb2oKkM5n+clwjC2exNclmdMc4wOT5cwg17y3zYJ3ozKYjTb7EvPkC
u6M0HYni+F6bqfmgoG8HLyfdYR9KHRf2KfREjofbv2MOExU7LhhTgVF0t8CHrmZe
sQCl8BQ9KVsTo4ViMoMH1aODyE51HD/S3gQo7Jcc6uLA+dSbn+FcFZ2qdzDg85aW
k/we1LmXWnF0DlQ8A/VxyXJgjpyJ0YKNboQ3cdco+nO6OE/k8UjVNAHj7DSjM8BF
5/kH/gs0cuEk3EE53mVryuUzYeTRtid25l5ijaiickWLxqR9sJ4Qi++vmlIF+640
lCdFwIfaXYSmGI79+8wTkLxA68GmCYDU70Oo9dzcv2Ip+8znpLpQeyGr4P4sR9Lk
OJBXj4zlSgQ/PGgBeR99p+Lq9L8U9hBNSDCrgaP9j7R5P7WYIOx7wpQPwOc6pbbL
10kzRNeKvrgfRYdMiHJe3bgQIHDI7GeiKouFU1dQUXRMgqaCwWcWdz9KUwrYiOKj
NnkVTSRpK7mtIM6KY4TG9IDMRm17o7WJi9tB7oAza2ghjZ4Oa+vjLP0c7N5xt8lV
ZA+k7Nx+P2sanm7gxF2u1YrLL530hJuKH0euspmlih6kDzgQDxv4EQmgtYUCJ6FA
ZRIOPzjmsJaGqSYl0J0873GB7foemvSz/HG5i0GsxA/XEGHMUbm6HW04l0b0p9Wf
UspmJ8MS86txYvkxEuLWJTOOcxrgDnEyTntuRFgzHdwudvrQd8Eqrknbi6rt/cPA
ifWBQ+2meQcV5MKylSOCwQvd300FzXhR5ztJPsFUNuB37rfQpFvJCDwR669qU0cP
Xp7IK5z7cWSE639c/x6P6bVB3mUuj1kfumIJg7btRY48/HXYr8XD2vIe18f7yKNX
9Jzg599bX+SvV6/MkghphOdWj58wZwkJ+gDS1jxBzYlm0c8tTW2j8gHdZ5JQDXch
yi9dnlSw51OyLpCjyc3Gtulks+AhdXNmEc1dDjF2hEiqyBK3v89iPq6lI0oySBIR
P8FPVBMZ9hc4DgAQokNmFkKryREkkAs4Nqg9ldvyNhDOo4btsLoGF7zljW9qq5aP
DW5GpIKIw4lXmHqNobGrC81Znxa7KpbJnr0sxUtnBDzX4cscbKcyc47DZ6yWFbpa
nB8NXja8GwjZd6bQ5eLJY0NMwoniDbQrCJvXkOZa4US+sft+QiAizCRbKV9AXlFY
oz9iykAgOS/PIkMzyRdPlWkY4SIy+9QlBpCvEr4RgKNJb1mJ+Yw6GaTQh4KQn6qe
zmWmfX1sD/n32W28iK7p10GjMZ/XO5yLoFVd4PNHTST486fjlnwD6a5ztXMmNkZz
yVqfTcDNjBvYZKBC1KoN7IAwgjEx7aTMgAtL0GHqBRzh2f3+IHvB9hPXm+HQIg+D
QEdECnaDbi3pdM2mSyy/sPrk/sPKdC771MpQmI+x8+Cu8UN1ZCqxXa6suQJO2nRT
1UZNLF7ogegTo10upVwgvGprNn/X6anMs7u/hrQxpCt5Jx6Pc7mat1CkuMOHvKEA
MxUmLlnqz717xM9uGUbM+X72ZHr9BEQR2RCim1aDG99X0AN7jmGUoYa0owkA0H0l
IT26oF2HQE/2SPdt9l9ZW9RT2zPkeZJGx/bKR2mHZj63WQF89/X12MP516WPdoZk
9eO4etWPFH4su/jN43SkE3/KaoZltGk5q3vBsx1viC8rzgwokZ3DcEEdjCut7ZEG
tAysZK21EjkUaRwT/0u544kEvb8Zf8Nm+3ttuV2cRmAGnV7Bmza2aR1BiRK2rWl6
45nKvk80GS9gAMcS42nIqoRu5n4n+v6N8LNc8XbCaiQ90ObxaqcjsISVyQKRkq9I
6O1p1chg3nWPUJrNbvc9sL/N4/XcmRaLRO3+50RtqXYZxz3bO9/kQ0GF3uZTdnyN
ZDqQvECZhN1a1EOY63KF2NjlOx0Nzrd+xzLR0MxL4mKmp9/+AhG/sfMguFM3IHVB
5ZezudqFWTkgADbG2YDOWIj0vnlKNXCqdepbRhdzpKmSVRkihvtm6rX1R1P3OuEL
+etlZFyBPBU/1aYa8xejdavXrzd0QDDTa4wWJao+z34Zuce/R0bpfYCwnxncbHSB
iNMhHFSTHkNWxxopg43sr2uWJlWjRSf2YvwklqCpG/WnvSfw1taf1tPwOQTAn4Eh
g6oHAVun6ChKTWkVrOc2gdFuCSVT7UWq+KFKWB5al/9Z+CPJk2hKzOGICHxqdws+
gAKUnh95De0LSTBWC58Hs4FHniLYX4woX2AXdvOzMZQwphcSk/J4J13gy5++WUPC
wDjzFNZzEyWJzuRe4F/5rkLUiuQBk9fcUTQdksWfhUYr7XG2VUgN10vmPN9QsVYu
K5CXmbbzdy2LQshPfdJUatn+L7xmFni5RHp9waLTJX6c4JZby1gJBh0vvj5IYVzJ
WVymdKZYLzqBbbqgCZuWGZ3tVDNVLWr5pvzwwfizg1LDlIfvD0S7uA/kU4rCHrPZ
UCYe0i2Zy9J27cbLYal+0s5ANiBI4uJn5CUC1dBxmegUtVV2HdWJwxQ71ITom9Xy
VVI/Or10Q7O2AfrD7kisvswKF2Z60/nyObMHz/9F0ALmfhQEqyBBiTmjfPKaddhO
d0ZEy3Do5geYyLvvDNt52CRqXDb5K7LctmrvqXSWNP5Gh7egFWBPets3Lh3VWW6K
t34lpBCWdenEf2Er76TQhD8WGIVxJcvxzAz6Tm6wuhpTkNqFTQB9K3o0IiTWRWaN
6wL89iqWum9Otytytj6OlQ33SnD9HBsCnjxzocyH8EqhtFuT1NzgsalHEka0EEjI
/z8XP1Ang/M41UE8ox3BvXqbARvfb0MjeFsKsxyViN3kMM7O3RjP+gWz+4BnlM8s
Lf1O9gR/sAuQIdWBeOCM22abRBGTmkb+01evtvr83thf4jSlNFe4ED7CiirbmgKL
ubte8WvZvfUvuIQGmY4HYN+Klrhp7lib6I+PHx8GdoXzZj5jMqMXfDp3J7Ht08PW
2TeDC84mJhEBWqSBrLxPlFI0kyIDkpsK2OAfwWO3ojCdijTY4hK8YdmAM1vSdXuq
e9Bd3obq0yYH6xpd1vt2UsQ/wEPYTIaIW6n9kE+e/D2ZRLFuuhEjiyCKUHxdsjj9
S8QXb8A8FMHB50CihidDtzh/KdrvIklMqq8uknq15vfaT6V7CCCHRLqMfVzV4NGR
HNJC+FGvPjyPOKCA34xWcWbUearJTbePRojhUysZlWjUD+2bEsVjLUuirvIXPU3V
gBN3dZsr5xB6vXOlP8P/ZHfdoAZUw0sqQTeOPYLuln+57QYXp/JaA+BxbnFz+OBb
tFW0DlDcvc3ZmKMnwp/v3gEAMTEBFRogxlenMKXbgY2eqIBoJWeisOr4Q24sYMQI
O0Le1AnuoD/T/nWAxqDFGZfoVK6UgItAyqbHJcPIWVnJIPiHSjWq/SL/zB7QSQ4W
taX+y/UiZU3iUcPg6Ksl+TophX176aObtjDWcyLLWB45x8fCA5NZSIhqmLa19gSB
iTwtJZFrK6+R2nScD4lXoLxisDdV5hrS1Xu5IdzpcbAl8sxf2BZiaORHPt4WcYot
1Yf7NQDGF7yLtrzXsFOg686LpzktuWc68VbAUk3tYsNw0qK7lnJFN1rgLZFpKFis
fInJ7AzuqkXOh3MgrF60+N7Zw4r5m7p6UxVqck/YT3VJ+cEgJUqfcGxG6pM9aqt7
1Y93AbXHpt9TA3YIkP5QErbZDSa56XY3I26cZyM++VaLa2W+j3QyG2osg7Yg0ht4
1mIN8PEBa2QiGofMCArsgS3L4hYVAMLM5k/3pLRjQl6ACvSUKfXrIHCzLln9dao3
yXwi08F5gIulJzbEpZOkJWWmIMNc+P3kBninJeZsXZ2OtjgBneKlPW8Cd9o9J6Pl
JOEjyGD8JDMifHpD9gPhyHPJFEhizeff20PZNaOvAtV0Uie7l19lIH3ntWQ11Erm
LCfiA496SmAwashYjKWnlt2Dknv/9kak8CTxxzfJrHYw2jTFFp/JS0UJjZXwBm3V
JVyn/+d9enBcj7VkWYxcg710k564Gzj0Qk8fzPaweIuRBoSabo0CQh95Xf/zKDQ/
p3ncnMJBk+Z7H5lC/EcFRkSMTngRt912wTJRHCofEnn6wcYq2Ee11jgoOSU4S0Pw
fLxkyvoa+ymniaRVmrK3Ec84oyqvR5/QW9H+/6DvEN7U3EpBNeDz4KWOb35OCyua
+WKDZz2UyGRy2Wl6LWHYrRdb5UOPS/TJVQ/nJ4lW8dTdZhNEJmnj0IxfNAbf2mar
Ecl/jS2ZfdK2j1d/b+UOAdT9v8OjU+pbX5ShKbTQ1OgdP3z+Iv6EuFNfZ95V0+FZ
NQYYOz94VwSPI6s1QLkVD4ShXh4E9wqR+TsgLUD7cWX4KoErz77HC2fsPYgAkyQs
5IHpgyu0LfXM9+Eh0asMm09R6CdVOScAnBonhYNthtns4fC3TRgR4UgIkZBeW6r+
HgD8hZd8ijNQW2kIdYR0oXbg4bnSrl1Kp1R8LOpahhUmZbDMUIq8npMAQ6hrbP1R
ophyIlT1JNv6nF54LdvFXpMqNcUxvKBnaPhzJaj3hZ4uB7eOTGZxndWBkYnCVBLO
zWDQ9MbOGrTNkfQaR29Q/0rDA3K//W2MjMbYCAeSy4d5YFVl09ddwcUKIMUBSOlv
PEgLT6UrSks8kvKw+ynlBI2PmaKdrVjD94DPLbgm2UDOvXKLoEys05kYuIBc3OsK
+qDHRFMrF39Gx9xtVRAR9v0LlRClc8I4yKlWV1TqvLf+zRIBPES2NYlk2dfNE2oD
GhSjedx2EyLFbDfrt8MdMwc3UMiTHxD1j6VBSiH7p6iX5qVYDhV36bGxALolUQ0d
+kAYGydW0HXMzKMrpQFjsabm5y/DKFK8fXK/lLBtPAlgtkeb0s4YVruY5luxZD9c
gvH2peJADMfpaLxfd7fkQE+Fo2fo6hlCaIZQzeoRHe3aOU42FAzLpTellIRQmx+/
qtYaqHbzFPo6pTPdPAD1guzA1PBt6GNfyV3XWyWe2tS3YyeufRw3q+ol3TpK6wJY
oJX0hFFhMdhHZ7H82qa5G1+bRlecia8Jado/Ni35fhWkO/3rEakB2bPBTwMXbohq
EPv3Sxk0RuTXGnvcD4XPQEmkGm6EfHC+qETE5/zUaX1RVZEa+FWWB6yv6DDl8Itm
sgqBeiWvHbOsOX3Pwor1AeNC2qwfGCLOUZvPfDQJURju3+JK8Qt06x7Ljwm6oGHa
CcOhtyXGYdy4niATd7SQqnWmbHyVpvnsVKwT5ZFstaGt4G7vhsLhj+8TXe9MpSYY
+KWwyQEVJole4n1tdFs9BEhn+CbyARr0nJp8NpyofEdacCMCt8DbsUWL3//heyXt
iX1uxzYizyaZJOCFiBpd7YdfUT/5WQiRc0z0XY8FxFfuDoMOv5l1oSy4yQsD0ybu
UilEZn5btzXSVYfv/wtSKMgvOe4zfLnK6Vgrr7PREZEHZ7mhpM2DRAI5lJ6H5awP
ohoi1mfB7UHW6z1TpJrnD/Qhumctu/uCBOgQ3oEFBF6VG7mzgo6bDzq/bpveHf6n
rclyqZ4KHYTdbNz/YJBhVnpUJv00bc8aY9eswwTJO6q+KIiSoAlHui1hPOmURrWP
qt0Ltn7ZvoSgpszDcehzOmreehdNJ8M2T00swUafvkZGgFK1Y/55UNF2l03lYkzU
QQ/Jgq+lOtvgVRI9WmsWJu9JnCeYn1WGnXicNGvFINUF2jzkv0qcfN2dY0tcfbFj
xfZe5oFqveyC7x+HAa4zGpgNnMpHFd++Ph6D53d6xep+34hnW9bdBBkFmMdDIEh8
jwqbcHGerEKnHqmzR6eyWUJArUZuFfyMJhZ0SoBKp3W+tH5FG6xhnxvEO/YVLf8s
MntCkKgCaqO5kzExuKsmkvJODOK3N3EEPjCWK7Z7tIrhzRTygKXHYnl8piRC/reh
rMfT4Rqv5VJqeAJ+iJV16TJwBUuju07GaD0xLJ3SUMexL6+pw+oj9+XY6J6apXAJ
sfkBYNpDs0gZqK+C2M9RmKoizB18l+pm8KxUCq0C9iVMmThvDFGuC9cmJojoNumS
C7Nc/kTfCFMxzxD8V1gKaLrukD4CjoF5JkkAxWooebvd+fTmtKW2OQ5nuB2rkh2a
jTJwFe7Bh6KfLs3h/q0g+T1oVvGfQDKggf7UEVmRIRv1f14t4Q/sUF3BcDh1P+F9
qFeoozrkJzFQFUyLxPNSppaGgpbo+1kqr0Qn0g2Jkrz3Dd81qpBAugbxNHY1Im/A
DZZY6GNfzTBKLJDapM339utD6ibc0JRRLvTexfYzQd+Yt+aiauvnaFohITFsoxBH
CWJvv45RNLsQnTvqS9iiWo6dZTTQP49TCXEFhj6g7xasKKTFKEK4S3+NdtFLkkmH
rZuJMNCaOYeohdp26enfDcdKaXRHBlZGoC65+aTCrDqTdi+gxrUOEQ0cY8xNsaTH
L6wP5Vi8cz4y15i7h1/6BugK+F4xeAb0jVh2o4fwwtjY4nQTcPunQAX1G3sv04wj
KhcgjIh9d8uWpdQpjfMVw/GkcJRgIu1OjZPgAMXP1urjODZl7mtWJ4FR/WXCClNN
Z9DwJ81TkiWCC+4mOz6UsueqWIsX4ePzfeKl1UjG0L4Aylipmo/WyG3kD96J0CgK
TzlW+DB1hfgS5+Q1XA+bItolq1w2Ebw3HgAUxJHY96VFyPsygIPZG+sPnIBKw555
EIJcM0haFzJAEJEhYzV4laveMULZqOwrguDaDvWxy1PUXfJlZnhjgHxVUZwMBqg8
2eo0GADzql08e76O7tXphEG3GgfaAWWD27KIy8pL9XRBzlHDzWRAi1B4SS0tF8eF
MoT+BGiSs9X0MgkHkx4nKEHmEuKoupg1N4Ji83ZkbrJ8QRZb586DDJUsUhpDoSEj
JrodehGddMRv5mMlYoZz7Fnk3dQzWjQVQJxNfHHpSjdBXEDHsYvNm1c8CxQl4bA6
oXWflygquuhec8XgUbQxEvWJHFg4zTrBbBZ7fdZfkNmsCdLGqJuaC99uxTDbhRTI
meBAhsqFS0p7yoLymU83HF/0zS39jxj/4Kgo8RxVFgTPTUMx3VdXux7p63wDZx7R
C85ATKxrY3DEmqhg0WyLMblYjsxDBDUusZOj/vL9uRomnxPw+XLB1wx2F5kFvOsa
4yIoBOzclCm9hsQ1GcGqPpajbGp67pOHrwUhoIZYMOqP+Je4sIgIgQE99RoNvn8s
RsDI7HVSj0l5qHV7IOdPTKxyOZyw2SCPPX4gnqjJVI6tOABLAlTHzBlS6TQgCP9C
W1vrGLSGnL/YMTD1Z4AruMNxu2R6XFzYhyYw0+eE1Rsl7SGhZGQYLMXwEl2SVNFj
xSDIPB0R2WRF5KwmHv4U4vhNhrpslL6HvxAy2h6l4dL7OiWKO92IQkD6IldJ0H4Q
hVMKKljvcXCy+wD5x6naeW7/OGS3kITexXZgVpwT6MAZcFP+Tle/8lSBhjenCh1A
2+TwOHCJCzle782Bki2e1e6FvgdwimwOc6vP9yplHVPQoy6LRjwEoMzm/K11Pdnj
IaKIyMkF3MDlY9EPBl5PMHNh8ZJ3Fiv6bPDkJHXVZeDIkunS+gocdW8aeI8UWtiy
d3HOzs3hf10Oa/udcVjEQtuG4A8vkGL4kbncd+7HOJkA7vBZE4aeqiT3ycJ8VF1m
CJo5KhI4gfm6iryoGHJ9O/H28a+4E8JDQ1PPgq9EvE3/URLr22IAMrHCHW+Hbxng
bGiXrsLupZp6i1fULCrJV+5f3xLEYCLfAVThPch9WCxgSVC99bdtrZQG/0E7qGn1
xOl5i5QvDlqg2Xmi7febm3dI1LPgOeWbDwrgQPDsyFsQAPZYQYlfDZuwv9Dt4PAC
fEFuJn/8xJoCuaqZERx40S32YTjHhReuxDrblXylTHdGi/BuVmLkv3ba0n5X9PaP
QVzra5GvgFkOv6GX6WQ0KK4Y9hcJgY4qjAfhnzN67s0K7/OBJEHwrNbs2rMlwjKs
LyVQCHC7V+HyL61lHtjzT3QVXsyeDokWNaT07u+V72b74nSitroAkfFnQcrcpa2f
kXqn8doKy/FCVtuGtJa2ySzuGEnCQEkHPaNkpyMep8/IOlbHZuQINg7lVsFWW/Nv
u74aniBA3opXMqpriQ9E3SrFr+A7XQP7/cwpAWkl4hKdYVyZTodH1CP1Oj363AL+
yeL1x8+4peGNRvyXIIaJUTjLqEb7+D4mrmUp02lcOKq+66lo9gx0bgm6gA/bQCDl
pe9h7+ALBxnudXjVIg34yQeRoPCJbbY2EI7kNmi4Se3lS/Fuzmfi9nkf2Y4x0DQG
3Ke678gOeIXYdmZvPsTV2NIStI2mwblMVjSMirqTqmRlHEvWJLhsGdZkxgv/FY90
2LA7ByhAjjQ4gEcgqO2EP5CB8mUW1WsNVhI2ncMn2qeyIHHD4VFqEszrreS/le4L
Gd7KJ3cg8eGwaYgUck52ozzDpYvrh7o7SbUsnfGs4p42VlwpBKwoidirjRnqmTRK
CUPS0+AznfEyw5pUvMBAlqYBf4N7DSV56YebSpd5OZ5nxvipE8hMwpEe9iyvb4Tv
m/NoNBEE0NevXNjBZPOFd0qBCyegqQj48KfONhR7nWwZ6o9ii4mq51ZSBjTbVWuH
igAkC7u2TlEza+1sviVa13M8Lojy3DYgs8p2/2Nskr8kmLAFZZ+ESuyujNmhzVTt
5D/bvbu4kqguXdZAMYUO3+jHR2prU+STTST0K90mX89d+qiwo4r0EYJ+7MbLYPm/
bGL2Y3kuYg6OktTfHrrFfSE0UQl9LvBO+83jHWliao37KPPzxAF8QYtNRUCJyRrl
MZwFiYTu5AOdinFJPyGcrNZHBj22YHUdW9EA+jVE/zdZx3QFSkn7urjkNenzJd8r
3BObjhzxA7J+ZVIpfMI5CELzsXdLXz8gVUBqpHaPt+VjVXrzwSS1HTSwqOHK2xkQ
zFdC4HASz1R+eCi/NDVMHD+Y8MOJiCpeqiVTsKQ/XYVKe2QKv3mwrMMEJvpsaQQt
Zyvca0GB5eaCcQONC4HzwTYaIpoF4Paq7S6P/uWO3YAIsFfxUMaBw3Kgwx0KkcgH
sc+VGHihyKa2KhUq/tUDRskLfrRXaDjbmA0OmJjjdliLaQecZQ7zTp6DTLB/wvwx
qYr3t53vtYigptej9TqsKBI6HvSYkZ33ezoE1uz8zJpNatwZ2ZLsBbfsTPbJlda9
a/itM+yISW7XJShV5kIEeKjnzQKfjCNfJVlabhiG4nxnzSNyOHaKPoCPI8rs21uK
iZlr/OxSUa+0dSwKmoZfwuvVozXs02fcOsRFTtQGZCWElL/i0zGH0JXdgB5A9fZK
wn5gwTYemfdgl7CKabeaqV72C+q6xgKZm2KNW3PnqepDqsTgdaiFcDM8JMgtP914
VUCZjYP5HwcYGHJ+JnLc0uLBm9kXIyEMs4AxaN9iUiQTZ8nXzD2uD3WO77nHfRx+
ZpTwHkqjjiU6AayL/0iLASOgYanHsmP7iuEaqRBmFBmPMyuo9UWBpMl8NHZ3nIhx
q8gDWC9yqwnVswSvtSFPQUUzZBIOnvGzEETDTZXI2feWV59EN0kE7YXvS2JXi7g1
H7EMsg8Yo9C+KOVUO4sHC/FI2slhqP8exK9/R5tqU0kD43cKtjN6jTIupkV5dO9R
NHPicM6V+XbcIqTSaDhLo2RmNQa8hjY0pDbtdKz/WtysFgJ6rRbCr74SmsdTDclE
gpY8R57gIVMea91lkHLqIufXYfkEv2MbB7qLPjbFeRoLf/x4HB6rUdivCdueWflD
szZkDtaXvvWqRpZf0+LLX2CU30mmKctmaxn+yCSd/6RjkpAerWdmDVyYiODrCvPU
SDEhczPT+0SDwFsK+oEWbBzrilCfP+ECqGIzy9OvCLl2JVjNps9IunUnn3sY+ty4
4oLUqH8tH2ycm7Aif0/29g99llFglbmRqTwJ8rGaEcmU4a7E5ywKooJtLmoF9YT6
iufYza+3PXsnEZinOb6J4/dIl5bxazdsNII8Mc/jMKFVX71vdS1wrPYTPkjcI/9f
4Rm4U31j5/fxh0TiBLxWi8ZHHQhQco4jKS8T6jeZzZwYHsZW0p3SVAVNHO+75Dc+
7oZQ8wqayj7n38KL1g/yJmbYZbkzA0+Yw4NR45hTbk863Fams+AMZ8eN4dKuMcoY
O128NBkiwmtelOxYtqtunqrGP13gad5aC3Ou13Mu91f9ypvQ7PuffKRwDA7P18Dw
6fn5xb8FSj/mwc41oB4OAVNAKSHji8/ZdT+X1C1gFIHJ+oBYeSysxi+rPaCy84xl
/vJOnyW3THqshpP4SeTVdZfCtMjI+6JEblpIniLHrdXSZSdt2yqnneRGW3tozzil
CDMlwWyysilG5PrTbrAOBePubveByV26+0dYF5Fr6A3DxU36IuJA4eLrTlSqH/6M
tH00mCuVDTnwQELIKXpWhF24ldYyP2Urx6GD4BbL0siLlKWzWXpi2YOsFxmtShsb
BPj6C9LKz1AvxEWwSOiK5Lo+eby8z6xPNT7WFUR6O+DPOO37IBzIavpuYNagc46M
06R4CFQvBZ+zEeOl551BsVIjXvAROU30UaLsjwNsmh0hHj8A6XQxN6qCc9RwRt7l
3fRF7kvwxvFDN2MUblS8qTcD6z5yueSXDJi/prGt0IvTvV2SONgf1ioC0iipH3CZ
wZJmVBhek+BD2ft6zfLqa/9UQ7rrAKk/vMBv/RPXAP2WqwhXcEaFK41rN19HNc3x
mZNO9GtwLtb9QnQS+Fo8AzUCk9hC43jC+lsvJaflben/BVgpIb+1mGIAuETCccYy
1OWZDIF+6ulefZD/qRwQO3UGKjJ4H3Uk2dHdBPFXRX6T2QuFuB11DwsIfzq6WIGY
4VDBJCZ+gYbvfO/lGmv1C5uNgGF3rxLNY5N1l6xi1s2lqlQXObDOunnrYbDQGLBv
+/iyWHGeBESxbeKRlNc93L5zE3tZ9HzgdooH3S6BlhquHioLrFWOjWvlLI2YAGCL
8ZV8AdqUqaYiKz4DAudv4uLkQqNUcT9FC/igQeFGYNGGC3/X9JJcKUA8L9yw83+/
2xJZFdsRCb9aQ2YDgkFoqz3xP2g/FrJ7HSIh7Xp+sCw5ctY1aNxqEE4He3iG3PUw
f7IapPyXM+uA1+IjVRdfDonamjJvo85UBudDmlqMJMlLZIilsj/ne7dXQSLKefmb
0gMdA+biBevuE8BzEORAKZWxnPPnZtIdYSNb5RAjOghnIlSFAPBYMFVwjdp2wvM5
vzYsJ2pimrcsUl6wazK8cjnw9ilBn1r85r+1O/f+R9qy4OkGWbJM1WTH7yTw9kZE
0LLuC/ku295KSSl8mPeNmvvpC5iCPZm/SSjpaIABS2f4p8ofrCtLQfSo5xa+f/Au
nUk9hciuTNLw7KZNoWNclct8+BpZUe6NB28NPkXccp1SBJ1ZZ9QHQrR0GlIRzhq4
NQ2JjFBuI5ROqeGR3q9ZkASwXz8Gv6jXThSUNIlY5yuwjtooJiX99oCJECBw2p4V
f2cM/CMrl4SA/F8Pm9hNioFfL5WcottPd4RNDJm85nxQjduuJSysfdkKFcWSL6Wu
TueLyjGx+4f4TfnirTdlLlcFL/50E3e02IhdfzZyFL67Lupt32cbdGROk2iSQDA+
jY8XU8MfHbMMsPtvbd6LCuF5k6s2IvBgTWB7WlGl81acKIIM48ZL6DUYZ52IE/Up
Wtl/p2NOGP2UtDXbjxMupzE2+qrvXJZQMRmRUfWE93z9iouupL55YN/iqiGmObo6
k6latnte1JO+yIwhrxQbH6XioKQzWWFU36ETiazMkYbNe+aAWEG/bgW9uTMh1F8M
DofnQd7cA1SLsNvqlsnjppPQKSspcYl//IhPuhhe16aTN8hVLiBu3K4GA0RB0y2X
d+mdkxe8FhcIe5/3SYqexiRaSw+GKY5GfXk8k3oNBKUFVJMjf28Q8L+OCZkdJn+5
fCort/kJVNhuF5f/KfBze/666Xdhc84d4pKPld7z3QZwL1xCKvBzq4vJysKSZxdW
++yQEI5QdZHR3Fo+dLtpem/GSNboy4DPeQndzKwZKF1ZIL1FCZSKGDNBX3Y/aI0Y
Oy75674Qp3BZYukooUpY42xJ3PvWKpljqzngVNFe5nWiOjPCRqscJ/m5kEeMFCu1
FaOMRjXXj6U7ByGorvFzsyTR6e/g60a61KZgqFuLDrQ8bD9mNMo/8ZDzLuo1oFwT
mNbZdKD9/iF9KY8t2tDaN7TCRKPEYoDWFQYbFHBymTiVxe32bJV35aouOhrNmOBn
J4a7R6HRlagzAPupamXCRhHYb1Rf1P/fmIkQw/SAmoy2Q1bCsTNTKg1f7ok3f42g
vs2k29g3JqGT2O6GE3utq0j8FTokmWpgdDPYMC87VQreXyK/pFYEE9D7ktjCyceS
HWJCgdBh9eFd1z1RhEEkYjMX0ngZ2UAyADZSlHpePE0hapN/96p9znK5T7lv5lyX
6fcB3GDTNziVbEBROc0LdgucInGf6X8dj2OdoMw7vuQgXOgsNUPYlh74Z4h9Oh3T
99czk+LoHtnOkYHpWWWg+fXudKV8/isV7jbnx0RpzG5gkOzzOp9Tidk8AwP6G+LJ
X2WTmCF62YGjd4WtWIhYxyHLbQfJwXfmG1zpwXhVVck44WlYc+BtJRRqBC6A/b/0
MCOIfshZKr6NiG3zZnls970CvXXbLGAxFcWzXTzTmKlFYwaNSQbYAEtVaRSXbs1L
6cpj2St1Du7pLMnzrZmfaEUMxRm0nWJ/hlxwEvk6WlsABFX/dFpMjXlHu8OVuVYF
THhg3gr2FaZhI9YIiPgo/qNuhN06yeWf/r5HpB8PToXRv+I2uqkUtA67kpe1UC33
YHAPx5mKGli/FDEyJZiJMH88udBMz17EOZoMSzMlIHrb5Q4Cjb0Puuwt0OK7Vu9R
zpSvHKGMIKdBuxd2LpOcslVN3NgaZNT7KP2kfLTshsTNGajZw0aU/4EKV88zVHxv
jdI8LAnR0ZuJrRuLNnrMMEaixTCV7xs6b1DbljUQn4oC2ku3AaG5ejP1rS4/ulGu
Z907e45NlmBUTjd19YYXzRtraefYPjlA3K8r4i7daXlbz03t9a0IvP+9cOjvQv32
EZIGu1uBGbTR2ZORJ8fDdTI3F8NYqd9l1OER4hjWb+/wspEPnmlzx4TTkhUSPJ4E
DQsygSCXdflrtPkOHoka0OqW77jeqJCsvvRchIcOYPox5IaP1HAUsPunFGoSjXXj
glYPdiKzxIhdwLNbwKi45fDJm4mqdwJBDRmZYKbkASZIPqK+bOpNzBxD3SK/MOm3
JstT4R2XC4wB2TlFv7/YmLMhgGZaxVfmXM1ecrjjCZmYcRMtD/6l42V9uQnG9C9A
6wYdl1FV0FKhc/xPMvYGSvlcrLPaIcmvODHC+WGL77bERPgl1C/+r1kmuptqVM7T
ceSPN/wS3qvBTbYNy56wNcTQ1Ui4O2AAX4Ne9enpDOX3wz73lrI1SIHq7AAtHS+X
ud9D8GSBl7ug2Nc+Uqt91AJ9z+fU7jh8h+xmatMmhUvL7/ha7HEo0nwo5s8MaeiW
6ZxaceMXO4vONbRezHkrImQJ/uUt74kV8zVA/yzimeDDd8KcicE1Cg+xizHsmZuw
MDdpcMDMc6rtwEtRLfmrahEAEP+GmAyraPb/hzrR6wnuU1DvOcu38trNUlzZRuFN
FkxN/uI9fuUex/rHqiVs+7Jgsc3at+qrneD3Khg/VLrcKVpCDhxejxj0wg2efGEF
2f4TKDTI52Tufb01sSsl+29DsT9lmv7HYbvEMq+ImoI3yTckyQt5LkOKYZ/VxMbo
2+zEFEUHj8VCb9vOl05Wmrr3TRAaY/xzRW9bxR4NpNCBERpwIge5VM1IphYB+KTk
b+dKeZtLrmN21B7+q+r/qtO/EFCeWBW318FnG02TZ9PQfRLBbRlsOnsKYG5Kp7A6
wr5fFMaaUZQL224R2lxOkwxr3U5zIuMti62jeHIONJ3RKeq52lDvBezUIHmloeEn
lVAGPMcn80FFTrFZnbv0d9SO+MxmhkcT+G1sBsVgej7oMMGZZHJVZVn3IhSN2mPP
geIsgMo+iQgDPi6RXo6UE4Ky2UM1WEQWC6JS7TrQEo9R0Kf2Cov/VqkDG5eMfvZr
MuDMJb8w+tdA7Qvm6RcmTjuIV47sAqkKv32iqYW2xKIEEWwkEUGZdSQoEnou1jZn
tjBWr7IXB+WcQyn7ocOFN1cQhwzW7dixgf97UMTyeh96Qu9AMOXBrPlVvkOkfPDe
BhqSIKoghYxL44+c9VjdO676s7wF8gPsnwFi5S+JCyIkJRiB/oGX7emhmVan/UZF
I5Qld4cxEgAT8eYSPx/8XOsrz4q0j3PGgSs/gLKp1b8rOBdbELEDUfTBzvdwjhW3
e3Vskc7XvyrzFwJ+PdW3KZYjHe2vY9Zmk6BFfGJOztj3dabLyt24nK2D5RupbfGj
BvUyOOVrfcsYv3hlpuvqowA64pOHUiA4dkYEWRIHk8x6nWjR/jOhoBciW4EeCgpv
pAXYhgWP2cD1gEM3b3HvgEEJav3Fljc0YzxQlth+LpX9EClGwOaLP3WoDQSFLRfJ
xG1e2U4u1BQnUMQxahap1U9lmLEfX4OZ+rQ1OMCe8SAcAfKAoT/SscBRQWR4gSll
/NoHnU9OlwThWDH/MMkOqHhp5OESvXLIPvVxupFfedVPbjGS8N2dV/93gtbiH+MS
HHz9snefT5emZdImG9sal4ccGgFnSYEdDoUkU0t4r4Ir6+d1g2qcQy4tS0zdiFMt
Cgj9QqkHccsKHi0EYxuM9F96PE3+UefyER7A9HBPYkV39z1z3/q0Z+weaxPp/vnm
4I5PgyFtqTvIeIpQ7WTtm7piQBSBvYCfwcwiagY3xd6GS74ciG5KDLNnl3NTYI4M
WNQF8497ysrhcQy3sp+O5BV5MEhPr3GWUDRVuHvekK5mXZNF+NmwEdQ4AOZ17PEJ
4JlPJrbGjv9xj4CH6pTczDKsvu3ePnOdv2iQEJvbAWndsIDO6cWEkz6y0nclx5o2
CK7ML7WAsJrOPKaqib7lOMHvb+0pnC03ryumblLC396GNEWfRhZc0k71YmtTvChT
VjyEPRAyrz+PSE2tUkDBLBbosaeXDtBRpmuhrdi1iZKNf1LQpxZIvQrTYJiA0Okw
yLbOMVyN/0Or8BZvqiMrVlw1OFw1Tzy8JPJ+L6y353AXnUjo8jsYYyaiP6xx0chV
WctqpP5QrOKjvQajO8zkqvwKGlqabfOkh1WF2NdUBbUDp261AkTgzLJrvkg+UzXJ
Pt4kL5Ugd11ShFdWTChnB/DRsr8F9tFgw7MAL2XzxLlxXVLxJT7WGs+2znT24GXQ
NYgi+M+amENBaVGfVIsqOmhjOIsvqFokjepJG2J2L1iFG6BWIE/gq7QfB9jnwXCH
zfiIeS4gU467IYMmYhv+T08Y27TGuPubESeuaqX3XRIe98p8zo7ee7d81hNWRppe
WnM5jidSCZBGgO5fFpkvkaWDSFm2EDtBLI2xO9YGSFAojSDUPGf/Dymws11txOc9
IMP9r3jUSO4lU3a/0TAMfM4TwP/CMLRAEnrz51FMzuyc0rfgD1cNGYCzmPCFxdWz
uuU9GkaulN0V4W6XXQr2ftw65UgL36zlPTw+ErerNmKETnJxSBUom33snMt3wW2s
WzKRU9JMNbDjgRAt3rGMCsB9+WE3xQfMK1ETlh5ZvYkWEBdhQ/NY2Tx7ljgdkJ3m
kyuIfWCxazqMFlLqvDWkbPWcgjwE1WODVRoSeQKZIW9z4W6x9lgR6AzfPKYVvwtf
xXX4jpI3Z2EH243vAxqmhHxm0nuqW0O7pKzF0grmv+tVvHKLp07wvXfZc1/hXQsy
FaxoebVpp9XBobKz903UhhC6A43cFNsRbpG/eRKCqGapy9jcR0/bAbjF1peg946N
LizKjW+p3YKPVmH8t/ylClnHN2FNeovUL49PJC2takEfSMP+OGr5GQSGxjxIfT3D
STTcgYKDlXyxwVnQsyoowXZwDwtt/vnEbTjyJZ3UWwlaIr78RemX9llwu2Nxn98j
RHtgv8nnR4i9DfHS8/UhQjm/b5EV/A1wVMeZXoyOS1pO5hXTTTvjDs0i3E2bKAO5
T788LvoRT9h4Ds8rvtnTEER+TvblBdwA1tyeWZmufUbqjNCeEQVp9rcY+gDhEwAC
FVak9o/wuJdzv7NLGkT8XMj15N5kb0YBgwoPj7RbYQDZEWlIPDwfxlDCKdp/UnxJ
piqxPv7H/g+3JNsIRyQI6Aikd2cp4Cro4+TcL49AVIFX2cpKcQkEu5yhmqnI4FQ1
TkhEagl8BVHps+BAANL13guw+rEz1wLjndaPb+R7AQ2Q8tgtldDpa4Gw/hqJ0uux
OFAloDE/JoUbgSgrCjjHZP59jKBO+xDtmtz/AQcbUsU3TAE/cqdlbzi+2wMDj4qZ
OXDUM+XxuMzJChH97CbMXHeQTpcpugaogSP977nVZ/8OV+56kKZ5WH6ydfnrysIR
57WcfBwXGdOaHEXtSPjjzo9TKwwIYy/Fv33Qf7lsj2Jgi4pEmNiXM1miVbqdzGgi
v1z9bZvB3y5P3AonrEq7taJf/TTlbP9kRH2OyLXqJA/t2PDwd1+ZbG6meDQ/G01b
nEuuUfk879SXyF2WX9vcbOECzWKjFosyodEpVItMykU1umtp+nHdMyS+7/tDmh3q
60Uuo6Rod02/f7W+KlgwMNstOlhavHoFLbvtZTWS9iW28C7J++/2baZzUG5qP7nW
CZsyPWGZbjjoxVRAokqpdlbX7XE3tfWq/78OD7MZicsOPEEWDnOe7QTwpk5kppor
eUWCGS7SXHmi9GOCjygx0t2W3RtVyjrNKMJJkslSQ29Y6sfftne2wD2Y1RTANZKS
FkuS0/VFAK+9zX3RzUEVnZ0ugx0NPmpuGI3JDqihWtSzrURpK6lfrhuxbA5bX2az
flhGkzaG4FWzXjv4JoJd9umdOMdnrKzeVTqL9VuWJArt+MgSy1B999lK+YHBdHr0
L2l+sARxFnOJ0I+dhxR6yOXvFMxEgxPfSMKZtoKZC8IvsZJMo8o7XWMcYhdip762
Rh5sYQzvVgHKOitC5zAKb6R5tsz+DNygZaeWpOf7jz9dPb3l946+pZ5wdYQQG6+S
IjpQ9oMStwMWDIAW7J2KripgBV1uKK7RBGkTgffqt5rDIn3ix7ZiS2tmMMzMREiv
4hd4H7qRmk61TvmA1Bn84HMcYw1JI3JDhA1z2TCDAoB6wLgGIK6wacymQnrGbrxw
9+94niMJhqT6563e7Rhy53HU6oQi48YzxCRWCHDny7PEdR5yPslt1R5JzwzkTWgh
6DBW3+Uzh9nDw7d1qk9mZujV4MtExLK1ClkQwTxRlmYLgP99WHZj7nSxo0vnM9yX
dTnG1OTKPOySVyd859wHLuMpiPoZFWkg3IJV2bRKRyRlDvR4P/4dwXaAny73DQeg
u3m3jsOszzw7IOdduZFmGKTx7kzOjBfR1Z1k2veDOOzTPgLhedmIDPliurW815YH
1d5it5JQGG08o3laqCR6SDMqui3KrzJKbrIc1PuNSr0N4Sh85Vwohsj3I8hhJyNp
sNJc5r5GU1e6eQPjRfBjfkXUpi0ZR7GaxdhisOs4LCN9XtEBWEP+TFOgy7CJxnRz
k/Mn5j4VFCgIkgn8gnc+hnR6hAve3zaI6e1/FZHzQ6Y8co6tt2xiLdqNE9g/r6ms
cT2CmDGGuKFa+VbYJ8nhsOUzSZ37ojdmy9HTtZutXzi+L26H/uY+xU6iR0mUvc3J
uUxzyxaiP/1J19i/w5vV6j8n2nZgGzPAHxT/uIS24PxMAM8idiifXqhqjnaJDRNH
V3sFVe8lD1BeZ5hBufFIJJTMrLp9rL0Bbqg7ifbUG48YDQw7BJULVS+8eERyvHs9
uSrZj0tvmEzWGSYM2trfABLzROvZovlXywMYv0w5633H/MTDizbiymqq+uEzsIKo
KofyGy/ppbADiO9P3cmuXwLt/LoTSaM/+hQI1pl0b8i6+AdlnzrFCcJ5kn7palhj
OhJhOHoUcLfB0p528braNMT7iVAQyHJ86MiILMQzDgnjSWpNE9ZDXdLK1K2neKDr
F/9d0EaYOBf3E/jufD1c3pbO0BjxNO8T0M/x4bWARAIjlyMWv7n9GPDTJDmS/xTR
Y951vEVofN7zutga4ijccvs65MUTaX8TtZUaHAes6HD4LAU/WY1mk4Ktirv6EgGn
o5j6O1Q4PDLOMSes9oIfkR4xT3x9G9tqJswjw/2Bw9lsbYUmB0+arTSSiqo7/OBK
MhAkXHHnZqdq5P4624W+mTRWMWoaKNq2rJIURRT0PZXq809VM90WA4jUHijr4Mru
P8lxP7mCTs4n9w6YcVZkGYSNJANnsTZ9yTDj6nAhAMOOv+YQCaAPvvS4ZTMV9KzD
Nhp3cqj0rkQUiWd8+SPDf/F6ATf+XpfP6kxfKpF4S4+IviEeH0GUzFmBy4j1phry
7NwtzAoJwRw7XKajnyf7TCB0FVqKm2+svb791feMDgfiVF2ry7SLCYNf6WgPzbWG
nq0+8Z/AdTQVFsYuzeyte4kApuZqNxF8j7Jc9prIcwGVLX1k7Tmnhhxq8mEat8j+
dIY6lc3wLY7U9iYiENq0mmnT65oWcQcIOjF3blRWCgnGlrKNB4V8pnYcm06BwkCe
A9SLu5agSpD1MTL26LtS0hZ+ZhxkiTBmj0ugj0b5C79kUb3KKRBkypTT3GVSntMN
0d8Vdy99DAKzurNrbV2ua9XSLsAGovcF0rw+b+bXKIVK3tQ4DOoUvU/NVwta/+3V
dIFdX2iV2Kpf/EzFGjmHPPP81UYfqYYfeXvBd/12+qUNgqSebeMhFDOvcVMXl2ND
puq3F3RlWbNTn/+kMEvlDKhDRMJCb7KMAI+L+Gq7BK180DSWS5KVGhf8/FOt8RFw
SKLBT5wRZR79tOIrApsUvxNCYpzhX8jkGvlPMdLboLaD12Ls5NvkBoH6NLCo/oRw
LFBz1j2Cr4HfrjA7lLrCiy+Rd0fW2ewrgS+oPjzaoDpGdBOkGJ8ECccs2Ro5ERvS
JYaXnlXUU4iIr7qcxhrufzsy9U0FUdYeqCbULRXu/tNyVZqQ4nAcMU6e1COH2iBO
9j9ROsucOOYVgl20pJ9ogZr4mE/g1GPSpNwmgBPUwBQtURq49jZpuL4zpdDA3Upj
JXWSoK5dGNKppIai1bSt0fiFgaNlOqwCLZi6Bn7608N4g7rJTR7pIHguViRp5pJV
GaVyiFoYtAeQTaJSfIW7LYI4Iuc+piJzQNrJbbJbnYI7WPdoC/YeaKX3x/OgRxJJ
BeIbtJOxrtsz+xMaMYXj1mIdj2KFNzI/gdbjxDASX1j8LvSmFhoFs4aRiFEEeVqv
F1TZkwZxUTkSNhQtx3YyDPX8khrb8T4XRzut7IkCKjuLtya/Lmyp4V7NeFu9S0iS
wFGmy0GsU8hfaZNpxkfy7cYz7OWGFRsPtwyZ92o3dxYoCQdCqmJCVfBuk+DmldDf
7IPKVxuX/IU5hObXt/ae+ojAiOLXOFCUKFQtWfwpleOS+M2S7x0bTbAWwUCkvzIZ
zcMf92WHQbgO/f+9lGMszDdZosIO2K8EjWnDSJJ9DvhWjo/E97S9vdokwN2xKHNb
+VlS5gZ+Q6E+h9+R4R7Rk1XesLemTvhPcAW21BbtvAwl7e8A5R5b8l1vPA0eV9f+
DwXoggHfQah1f1+TwlUJwQq4ipIEHAm5y6YGGKzz0BVHYWBD3TS2Q8q5Viu7Tse1
mqyw2o9kGg6JkBu1ql1S4Zp8FoUoMmE8O/a7+qAZpSyTLYXwciwmAkqX1/BfI+Vh
TkLR/6IhVg8AmVfZi8XxCS+ArLaepiCs8NWI6ncXmXzj2v7yQDhuWa/5PMueXdap
C4oAc6bwKKzUJHaP2zcgCw7jlLI7DHjVlkWOtUCtdv8sVsmW1pVONnxFh7pmJn1S
78adiAdDr3QqKW6MbPYlzjuq1/S+v+gQXi29oRILn93LlCl1+eu8fLMpNQhhQ4Oh
jyutQ0c7jMkmPVeoP6PP9zP+PNW24oo9oI5wNtqUL10jkJw4vv7N7sT0JXYon3Bf
SjsZ/yuSAeG152nLtbTp9qWzw+aEi09o0bCiAnxjz+N43MqZ3mzueHJjjnWiRmEb
lPY3WVJStR387fk82Pwqa8sOFf34Fxmg5KkzZdkyKfsRc7NEGlgZ/RZNoJuIt//A
tPMZAq5LGMzhmAgT81Z1oWm/V+oSEEUr7mVDEGc5K5EGhJa5VuYDvjGxzZuIcnty
mUw3/V/gWE+3B4bJIT3hJvdZb73w7/7kyNftFNTxkOap7L8wA8jl42Om6YtTTr5C
EX20pB6/zUSCmetcG+T5KHUe6tyUzjkxUFEwRxsSPqwwvs8JVSSQVhpEONljX7n1
CwZO2yl0t9krBMjXC1t729MJl0QVYGKALp+/n1k3A87GoIs6h+bmgMD7jwCDyK+x
DFAsDk0pPm+7DZQdUtFgAQS1sDslFjcZheilawI5mRm0vH3DGFK4kv4sAkjVnGek
1Z01nzLmCQB6cv5ihq+L+ZHj33ES56/ql2nNnbTPrly6Hu0EifOFRgG1j6JfG5TR
3mhAyEOIyu6qnx6Ml8PznQEZ7312PclbrvnQVEfdkA1cBCCb1C1Zh8T0a4XUoCHA
EyWnpRrLusw5p1+z54oQFusU5qKPUH6caKuEuQDbVy7QrwQFoyXZ9KLe54tNgW9k
IOdHH5MAQo2bi/06nIjS9KQjhzo1YdOoKqYhFQErPV31NQmAoMmHFNHw70A8kifc
lmm9M6q9tHUg3QCYQuh9cCdQZSOZpXeLqAB1JU/00tej3Nzkh5rXNEpQnfdOlJR0
J5/qzN33ICuAJT6/L7tF5BNVN9Z6tftWVtW7vupNQsWay6TjdhZt/dP87GLleLqx
7xf9RwOWRdJoHB1w2AQYYZHOml6zbMgn7mRknztde5hT1AWheUQvdYUQlNrqfa4M
yLUdGci9iF3K+Z2nck39Wx5882GrpQ4rE2Bjra9Xoxw68/tA433YOi9JtsaqO5uP
e5RqkMPXJaSGRjCCfXPy/dTzFNo88KPIXGp9MG5ftOhFEKsZ2VskBO5akdKosTSH
U1LceaicxrLOr1x0aTvzPH+dr6xo4MVZFj11Xye56o7qcG1yAZh005tL5EqfHgDQ
XJoBbAk9rkl4V1j0fYE2CqS/MGcAzfNiI6RGvNzbnG47B5cKReGRIjICC9W03StG
NRTF0AByRF5L7cHAImTYvPdfyMjoyQ3p26S0Mbuj+wDUUBXBkLyGhdrSsjBdUIkm
NRA7tr+exPQv7ir92h0UVqGf9klEhFewYLN6AraFKwRNKaVIoJZwGk1giQmxvZ3+
Eib7CFoTzS2VKbsuhHTdxl1ADd35VEC3pb9yE+dlOE3HtUDr14FefoorhS0R69GQ
VheQqesWjzCTX6BzjlkZ4q68q0phLaM1U9n25My1/CJFBEPOIxUs/cC7xx7q8Sy8
+fJWfwIqXnDh/7Kw1NEyLwMBzpUZOQd6K1yt/GdNMJpK2V9U91AUk3N+L1HILYfE
0o4cBbYEovqT7SqtEiqxTb5/oiGmAAFXbogAYCgcntj/9II3E2dwOgxzF3xwqQRy
fEp/I/zr0NkrWN2q2OjaVHVooeV33VHb27JZBZqjeTJqA6IAfWzPiBnbkQ2hxiLD
gXYAbV/vNAA6nt+VguEdYtrRccBgZ4SV3Mi6zNdkQJyD5IOJ06fsgjnrBFZwrT1K
zIc65FYNlYSalDdp7XsJVWBuWeArGiClpujgwNrlnhUWNiV7sZk0+1+639fMRXdb
d/6Mx/vZldkmrSbLLQed1rQWI6x5S9kdVDzJRG5O1QW4FnSPrqobgaDezmklGQ45
dVoWNOVdDjm+bQO18tJh7UydGeqI4B6JsfcFh+9eINU7tOJ4RB6jAxePiUcSxcbc
irJrnvKqMlLo+cRl3m6xJSMSy9N4I3oXEt948g/vN8hIPm1g7kUb3R/cWeFyMNXn
q8Cjq8kXx4hfXuTgrsbJ6QedsxeS9pQ/Q5dbDCuKmRzwcT0YK/P4HWtm2HcvtLvQ
60AYsgBlSmtKsJfcZ1Uq/5DoSqwPIIiAO+q/rUOWxG/CdGIQ7psBMbl6cVDo32KL
ZuatDsBMEV3HaaGg9HMcyL534OMcBiOt46DsDGsrd4U5cDktt1JFkPW7WPCQKd8V
n908K2x4Z9c4BGtNU8TNmutLAIq2VCC6lztol/XKoYvbhL9o1mryltcdM1txlcnv
M0Zpba+zVYljP8abPizYSoDBe8mzMitgSeOuhEwDcqVA0j4Q2vvgA7URWJm4wqrJ
K2I/mP56+G5teXdJHzKsplUFj9NVqg82HxrcTZsq7Rzu0woHiyXNW/cnc1/jlDvU
ufWgG/+UMyRPAWG+0xSt+N9fpv1Qv0qW5YXXXErEl5DOmDujGoQyerVyi6H84F/g
i/Q3LuzelrrkgjfllHVSKzsIDCNKy1ADlJeaei7fV0G6c17RPDenC9EZdpvbHekC
1f80+OU+5W7rxcAe5oSIosZyaNNHXRKD/u6pDagjB14OA9s2lAEuZ1PFlOWXFzTC
rPJ2gnv/pJ35uN16+KTL6Acd0mDZMtNsrzyXbFP8l6CL4rSo5bN1wsSz0Vcahz/L
K/GwMLAE+uFkoTEHKXlU3lReIbgiM4d68gSQGSyX6CD3Xb85UbdqrzZDdXMECYnd
UrThx4fbuvG5VPXQZf1656j7AiYCpcVcmU3YEZZJgI56uAHlKj23JC7/jq7e+ycy
NsuKhm8Zfhl8QinApI7mfJ6Gi4iAU9a9LGBrrMvCBT5weKKxEy5o2qSUoqHAlvEk
1Q/mf6gecaRAg4Jr4NBMx+nCf0KM0BsOFgzPsRuwY/28aIFvgjDc0vSzYoY4REOg
BFGT6as1HoeMJQJ6iPKoaY0nByvhmio7Q7xkVglXRzYgxy5M296Pg5rhyixEHp78
o3T1m+mi6nxRpq/ZmhMtlNepMvwEqJLnu4SSzyY6LFUUfk46/RpYvkn9hz0wJqFH
V83WG4znyMQu1mhJOYSC40y8CO7Jyv3/7OPnXA9lcAMQGisDhHM3NkPD/+Qz044d
uEOZsamxuzAEP7CkMJ56LQtag46FpdfYgVfjIHD/gcFz0qZKr1GooJ+D2gu2rHsv
ZMAnjFz/uW2fnDYGxyiKVK46fHow8Y9LOv8ps8vGnXYTBjxUEyryN2ObyxONMoVE
lypP+DSYTogiMTDjqVjML3ODIFNkjUtyb9GBJOwCKz1EUM1D9tb6mq+b7w1Xba8C
NRh3C5iDVfmRT5TAiBRt5PcDR9H8LLAsKRxUUIWg/a5TYP3GmYjooRWxpiJ9P3Uo
XGlu3PjILNe2C5rRIykJWg0rRJB1jxTp8dXPfn9eA4WhyEU1PKhe+P0TlgH9iBk/
98L5IfUefnh539qqMHenuzi3KNUtVzk+8YvUb7RqhsEaAW/IsERbPq26m8dvhHbf
bj9J5XBZfGxAdJxM6SxwnmI2Fe5VPO7NCwBS3+BrAwgw+w0XCGuWhh8CRcFKCY9t
6yombmMKBPV8vEhLswrTgR9L2eTC2X8WJ4NrCxm6R2yVMd8dgjznmB6pmwNdECNK
s7PhQ99gR6+0odDLsKSUv19sCC60ovzvvD3YebZEjxbbbmoUOtiUOPgUW1AKb+3R
xqL8B1dqIHZAaGNQFJqoXJNoRk54Acgh+VHemR0ONgiU+b1vxkBSiVP01xRLVwfA
vI/hD7cLHTDkl6AOxMrg529c2dyH09K4s1ChPUoT8OYNYLgSS5e7wqHYI8AQ79oD
mBMTt6IJdblBBTpxtxTVOWkpvhUwNtDylMMe0nMBeUx3sVZaEHMC3yn3sDj6QsdT
1eQGPtblH+17lDff20Hu2pa3zL4LYVSR/nsrxbrMYd0Vjn67KVGi1Ms5Yk0T91WH
/Cc7CN7wAwm4dYEuYA6tcGrFZxUSlcq7+AmpmZdibltJ2YLE3BkJbl5K8cUQe8m6
f2tzKU2V6wVJAcYjZG1ZGz7/PQ6AZb5uXr07YVaBsHkZKKd6khtETSxBCBYm9xB/
4i7KRMd1z9wSbEdWdYlivwpB+1oGpj57m4oS1chfs9z9JDv+XIJRqpNw1ERd5pN1
QxLTESqwvXJqBSxreDzEJl0tH+eB7akwj3ss+h1fKllbVluUBGXNPgcgXg9waOtV
hYuEVnJtKOVjRA9/ir9/7eBhHG7Y8wQ0JErHc0VmIsWtdqR94WnwkHOrEIzSR1UJ
3AqMGg0Xt/+JSroX0VFZbBfZ0Z9Ac3/wdyUh/RRasnimPAGOHEYoweDOSt2Xi+jk
iwVV5OeIj0H03afEYxGHKMtz8nVdUSRNzdKr57GB2rY1zK4ykyLYkczFB+fAH+Hc
+RauXNYLa/yRJVkwi5xk6J71JnLcWNcK2qrZINDw0PsKb1BlztuKIb9p/UFnCSY3
C4AVIS/sorvwXZa+fGVRjOtruEpmaj4vl4HE0akFy9MFDTNPv35ll6L13PxJ3UVg
6DCiJqsNky5ZQIWapuCFWWaj/J0ICJKS/ehV6YIdT9G1+7YeJ2g8OntWO2uZBEHx
MVPZP6Rra6WiuadXd48eHXCCHeEqhOHJlEU3xucdlhvOVErrKl6QEmXgA2YdjhsL
EWB00eSw+GiHM6KLFgYAShucriBvE3cmAoa7ZJmBVLdglMTJJvEpYg/TpCcQEsyl
PmB2mvn2GfyGZWLwrs031x2G322yxuTc3X/iQswt4iIwxga2LGyHv5DZFOOrv69n
M43EsrpA/nTVCSiXc0Ob8WLz7QbHPhwomsNihMHaDKLkv86uIt8tA0meKnjq2JHS
VWeFyn8e48TqDfbxtsCGfyQRqq8jSeli1f7vba1bklOqmARkE3aDfOXgicgb3PvB
OyhpVQ8M6An/wZjLD8/qC4LSHNkVmXcHVwYlGxYmdR5x3mrRferUJop1nV5BRuRb
nRqZVd1qHLolu4rYwoKbhhFOIAXAT2eIIa/brihEr3huDctOCvMzNrhTQGdHBnk4
QbFbh2gfCF7F6cKDf2R0YcyipHT3vg8UqjJ3++KEJYeMERKzu3vL8o4AELeNNz9o
Y9qD9NZB1vEfn0Y+tn6ilx7w92DCyaU9CIogPPwewIXmZ9d1PViPOdvW9i0tsAaK
v0/YmY7c/meg+MSD2LoLHLTN8RFtt8JfoYXp61MQyba3pY5cNCPKobRncZ1bug6V
PH4CdLxb8S4K/Fk5AvSPNLAubjmyBRvpJXsadRFWcwm+kKntur7yvitW32YY1EKl
y9U6jCXBoN3pvuRlhsJvQl9PzriVDhUi2ssCc2tz4LYH0iZ2cWWH5m9HwoR+0S0k
liidbiWkNaOjkGgWA9UhBlUZDUC62F2x/gHhkU3q3tBBrXm/tQajM1I6XfsjNBcj
EIPxknL8y3uqmqjyXOG6A4tppHzaKE5QACsLnS8DpdgibpBhMiyTHZdwHEh7ZerP
aQRIMP348OVtWdPXyyP3wcqbIBsYo3T5cv/8rPZeKYS3YzN7HG301SLpaqiqmNwl
q6pvBfb6H0szpdyLAra2iJgRPUwhuf1y2kDeV3RhKu0UyOd1+tAB/+b3QlmMMyPz
8AtXAA967dfSEEl7y5idnnRJ/a9G0jS9DZFqKylnOylE4JnuLjvYGO2souhcDxhQ
gNXP9vKa3DV5LX+mbEnfiPKEQYjR56w5IeMsRuawzZPjAoram59HVQwBL+tphwFL
ywrqIQZb7OooaWBxLsBLPmThJQrlgZzZt0lwn3Esc9zbzJGZKKZBSpiPIelpyOaw
sZg8ayf5GcUB/8L5B+OyCM/hPvduX6WLhulm4syPmIGyXmALAmcp2jk4uYG5D338
v/2+LlyOY1h9WT84aytxOTCxQVmia4bAdELDSPzCeDh+2B7hsN0Pf4YwwTCeHAv5
LT1Duq1sKF9JG5ILPYMOj2x3jgzIcUz9uyOpXfUEuuBjF4cipBV9iFkvg4YElnGR
mEpBKmlSLwwfy/V6xrzFJfB9cNzRr08zc7Rr16T3kOXZjv+KHBVqZ3VGb1Qa19E7
cmN9Use6JqrK/0voHrLuTzGjyTKzGBE6ju6fPO1dj7X1nvldo6HVvte0dJQDhUZy
cO8bcbHjm2PQnT/DsSXx9T7NMiMvquVza4PUVuC+qIi90Kcs7zu+l0jq5Q93Dxh2
ztWSNtZZ1G92XgKXue+oxESi2uXEKEcWCGiemZhB8UEgPq/Bq47qydbOtQegfKMU
vtJEsFGve7r+UYGi2WdF388dFnVtGq4nV1IGYkz287oY2G2EMdhnYnWz70rfrZnb
siDDK/9XAEjRyokSIktvQtS7zmiEl1vwVStQGHdYzcNLrbPaCOeCoNGMm6imVVxv
/0Ddm/bbkbIs7fuMii6eNmDhvL07mCFDE5Vt+MS4fwskRVlXs8iDG13htQTHzqO8
ybmnbAFX+tPm16ZK6vSKmIcqPCDT5cOcEt1DGQQNRSieC1/MuoZZFkAJI6HXX+vb
HF1h/wHDdK+iJ0RP2vH9XN93WEHFGV0lhcDffGTHER+FZS9ViStK487okx0/9U/u
COJ7fVrbLmWRakCOMe76bc7xmi1WyGVkXNAU/Um/2LFpNzuAVmXkpb0sizmYhmEs
mZBSjGHBu4EaqnqB7GIc4iEpn5KA1LyWcvY7lciS5PV3iN0RIQKHqgGP6Y2CDEOb
9Fkn6+C7yS/F4XwxUy4ub/41VtewHganqI/HPgQuyvJTrzmfoQiUs6bjUgzIpaS4
8lwQUbr4s22Ujvn67aKdnVU8eJCeCCurLOW67dmJFVj0BTts95GRkfkC4GzOKB3D
jrGLf4Q8oAYjo97/Afe+t78A9EYDCq/EgZEoG9Gjq9AYFwxHzFMVdXzODNWtrZh2
GCFAkPNcTdVFCIH6koes9UVqPB7KIBvxwdkCLWkEygLtrLnHVDTI/VdGVMwvwhiN
ZFSJWyVCKcpiL4CNyV417lNOW8rfy1Gg2rJByde2rbvgWBMhN6Vc5XdITQbRw5jn
m5cNyRZ+2K7TzM3rEb8XwwJCLs+8gM6IutlnLkwlpjHXK8Nsux59a+P2zpXXk6oy
/qGjzU3zXXsQ8EO7mi3o8RNpODPCUx42xdD/Z4VHXg48eyJRxtFl3sScAkbSH+nj
qZzPh4lXX+EIeQU3dU87Btpt6L6UZ9819kmsrnmCv+nq77M51v+T2ubuJoIeomEI
MSL8onQG7nosI8N3OLOKYOLaUCmJna0fPINwkq/Q4U27ssjuxR10y9CaHrSwCBsn
TNy2UFpGqQe8bNjxoj6VLOx44a1HkPb0Df+cRgc1tFFw3rNd+SvFe3oGS//PC7QJ
M1bXwKa9xsKKSrN1rnAHZM1N6MPaPhyndvt4RrmY9G8zWj9VEZWc9pbbM/hInz78
nQ6Oojau1Xb6ONFmYsy+eB42pIr5QugATub/0rx1z2uE0mXzPTsFi9WknvShABLK
BVkrN6Rm0aFJEzHWXQnoIT3jNKIwjneQipwRIpQZlV7MV4h1oLzA44Gm/KI46H+C
+lxTTXNoADm4OO7wZ+rd6qRZAkUnEydadKg4BpRLl+J2RwowtL7FOF7mi3NJO+2G
COzXm9K9NgtZVNrU2AhmKQQVaKeoSWOk+cLximQBwn5npBPejpy21cK2CJDpkoR9
Spe0MxrNCWEUL0d+g+n+cqmM0P4O1sAlitex4rRBh0jr6fY0pwlL2X2FKSQvemRF
Fdoa+Zlpi4lih1jy0sRLrB+OuWrgaXDWLnZK6I1VS2RbrS9CajYJCmekGJTRB8cc
XfBGqbIHWhwLF30XN0gqlhX3yAPBDIbOLF5q6F8HNXK6I4aqBIKgCikuoI8+Cous
FeqBwHkyKUSb6/XftGjvjlJ4S83q36YxtD6sc0T5OaqxNR0N9XVXvuDWA3Hlehln
hvltNwwe+1u66Ns0Uiky1YcCCb8+UCWeYP4v+k3kJl2Vs2TRQHhYznIZpCndb4yX
C0MAULWfGmNpCPxq2X+N6H8grhaCxSgmwoVx9q4gNTSz1MV0qX8AiR12/IbwGivU
p8Xy75AUWTdPr28g07Z4753AgoWzvvLtz8JIlzLMT9LiptMt9jeXWxynN6pBjtdK
TihGOdHve7x2G33xmbqOovres/0n27930trAd2hqDyimPzazjCKgTUNyBTJzerWV
A6PJOS5I95a39K3xcfIcepsQPpOM6VOxfgwi5VvtTzKBMRW31XMqe64EQJfamfDQ
sdtCgu78TvJpXp9GHg4zgpLPgVK+6DY+U+0FOvDhRuV123+u5cum0WPev8OW6clz
dCy/FIFUVh+qkgjle1iQzoc27vkor0VlFfEjNVaWhphYt4arbLkGEkauz65w3WMs
jPArjeCGXL7089WEEh43pFyP3Mnm6SU36CKaigrhqW34mthECJ4NFN+qj7ksJU+n
6REZyH5Od/C1uwPaKPiGeOPmN+1L6sLHr4+piRcQcPBeRKQ2eAM6lMO0WpP3djch
t3Ai22CMNJffZCbJWyRcnR4/LaKZZumDWk3NP2dkqIB4dYKjgs5aakBxI2jwqJZJ
RFkRjkg5MtsH9gMR4JxVAvY0QxTrmwZM5n0ENTnXcfDfv6xGvYHaAGbe3OwTnk4x
Y3CN2V+fefNbBoFG3sm5tLcftIruR+w8oMg1IuIASXBZlfQK2Mwg7cm8Pjc9sGEx
MjxAzDagAsniacDxKcwiq8gyGSWv4y2rS7nztPATzK29jDczVyk2//Qs2lV2WsBo
9NkvdcBJAmzXLxGowZ0Iu3+kzwGQi9Hxnfsto6N40E8Qi5x/qjJeaBs4lBQkqdVi
r8RHsTGKYPG2a+jI94UAkn0dOaHv6gWszjr4PF+o8EC8O5m2lzugzEx7OlqgtdiO
StgTNLvhzeYb+XOEhR/iCiun+JkWrTgHEOTudobIdkWq8S4oWnklP15qg2PDXhWs
dy01TN3UQRu6F9uY50YJUOGWbSjTQyv05oLV40PvalHtbD+dD0Jf9Etopr28qotu
yhIiTKmKmIimMy1xG9bgOjQUAvno70xF/3DCAnP9tTXbnB7AyGcngX1P+XicG/Dh
8JlyRuoRzM3xBniL2jj9dldMD4tz97F+dFwfGXbLeqjoLOFiCeNbXAub2x6M24ju
gjVH7YqO7CPdAJjdorb4WZxbKrhoqImRwtbNFJYRLoE/f5Mp46Q7OyYNyWsviXyf
67C6GhfKsvKmuVBrXHqCgohrI0GGryxg4cGq/2Lux06thKFV6uMDxyKQLLiFF8EV
1yQJ6HPdZ0Sp3s0sEAc4rYEtlnqFKlta4igZgTpRM/Om9YYwR412rh49T2l34Z/m
P+5YQVMth7gIJdqngI4ma5XfoyTFXp43yrECDa3q0k8ATIgYJCIabpVstLr2YV0w
MZov89kjoQ3QCC7BRJO2D1kztO+Z2k2SeEOLiLfRfOlt8FOv5CmECUfEoThhJnVE
CMUAj9/kvzQyCs0kbQFo6EWrLqhMUr/GN1udSWetEjTYW/t5vkxKtdWlpjwouOgO
2BDE0smTP+EQcXsj/1hJWSpatXJDtrTsj6SjMPVTJyMFFjh8uSNzZD6F3lTTH/K5
x8xJmd/tYPO8OfPEHTRB/YcveughPaHR0JIvMou4fvzTqoKa/8yZ5UfbGadxd186
G2dK0Qn/+QoBMjaFNCW6j52Si0fUS0sfgNpvtVY0R+KodcbTMsrVevMoGVvGnHZD
ywlHtOx0sAj7mD98aQek6SeLV4K11IxGN2wZHfNrIUqJTBeWOZg9ij107HyOyVU0
CT9X0/8TUdxIOrMLKsFkVjKNWH3JnD65onKzTFOV2Zu9fJl8Q5QcnajeQBSmx9Xi
HTbqh2m2KX6O2xPDHWgOmK+xd5M/00GwduslI0gtqIizB1GHxq/SBGiuCydSRU/y
3rR3N4H5oDsHBV/0xQPIdrsWw02HNIMCkUycRmxz3mfpYxZ6tLdOgyJoMGH7/Gfh
ks9zuifof4KCwt/9Kfs0funpJ7q1m1vRVStcoiO38MQ/Fo1R2AmAgCqTfoBmGhXa
eEk45LgAK7B4jcYcJ/LKhywZiOMmNsGTjXCVqqo4iY73yWzdXpvBJrUpuicHmAIc
FLi4u6uIjVC3+RkBwvdH9VH8oBnOStUZfdD1D4nEk902twhtPQwF5rLY3ubUD63e
f8qH4MHPXYNeoG9WbTQjdtjVpMHMoRHOZIbtuyvmKobL/ut4g4AILn9ReBZVIxqW
04CxdhAdpe8JxG/lRrGTaYLBIJt9rBqAwbGTDp3qNdCVlWgtmUetopEW0qS/8OGK
/aCYCJGkb5r27mIqlLsNaC9J8FaO4pCdZYSExoYlvlv9W//0g6n/o0ZnnZlRorWw
b3b6i3IoilPKb1fTAgIO03StnjTG1jGMvwbqR95Sw1sYoG5eObKYb6gqO/3CkMyp
H0fxuszfqhnYNFS12KOLT7f0UuwPAxAujIeu213a6F2ZHAJ0ZNiZNMEpHY0+RMbz
DPJ00ACl5ArbYs2fbefItM3KBIRzTwErCdt5OZwYHWHazY9ovI1VV2PJbTb+QgXZ
auH0h39Mkxnc9UGXs+N79r5T7TZrwG42FeVsBLR3GtuhwNrEWec8O6SdPrDuflJr
APVYULiCfm1hX2wJNpq1CQnruDk/7oSrtfxb+tMR6RqIcAKP1FF3Ei+Nldua+AxN
lKvD0GptFGRrHFWrh69hs6nMTFwuNYfLlxkATPnzU/HZXxsCi+NTGRh+3ZRWxr3N
zO+QFLjWIwgPd8MQZNhlAWWskw8DiAMCB61SYCXu/l0C/A59NNmwUhhmSF//CEmg
5e7Fk4phU/yH+KFqtqh2oKIkhgP0O+1pE4SLr2VFxMGes3mSM9g4VKDlEJRqCtMx
RRhezonPF6vDOCffnOSz+Qv1McFCpx9ZVrax4sa6CuuPKjgD4r3lTG67qVduz6ev
FXmpJeswwND4icWFFjuuVUJAiliKV95xxa6LXkmQeH3j7AHyUzomwFb4KV0Pn9QD
Kd7WYKPvdTTWE9iQ9rOFbvZZpP5gl7IRPsMx8bkeaG4B82T7GuZPk2cfUD9DgP68
0tnwLPsVdxBXJyh+iLP7eIA3JxC+U+IedICDtX55HripfYzQftCJUd35Ka/597Sy
LeC66cJIQh8a7QR2iR4XprDlWYuQhdPgpZv/q5ade4lBwjfOSmiyGghDlaMavYoe
L7rwLfxqIhjaAaxhTMRH8+QzhPIPV2CVGTwUJOJ0+5g8OGU5Onh870apWaz5lb3m
xcP3/84LUAUIwiUzH3wwGiH7cpHf3V0Oa4WEA/Omf9JIsjtwsVJeTu+k3V5pBtVo
GoBSfk4aYun5KlQcKK2+tRmYLwK9ZNnbxBrDoZcJ6fAkGVNXytQF2LC9nPQGVzKY
lrlByA9B+U/Uv80cvHzT7nMQSFVliS4sB6b6M/pcjUrSCdh7PCFqJ2ao9qd41JTQ
oJkdUimRYiYd26TWaK+R2BejTHGmQxTHgCQJvf7S3bYo0hQOHr/9pXbl/oaW+HZp
eAxXZZk6L2cw4dMGp9d9vkjNHjtHIc/Sy1oBJtTIajd2UIp2GoP1RV+sv9mTSGSc
0YbpKnCObpGUKiu78LKUd1nsYgvf8N8wIEyO218iwJ5U2tWi8R8Ox7YHj8xbYXqz
Z4v5TArv4vSrWSNBJHHDd8BDdenD+lB/9jXy0o8M5DlbEW90231uoYF4KA1OK7UO
4XQ6C6Yj9+kP4Wu8W0mEX9Y23a9KTD7ZJtRQX5fMjhAkVXjhwOxTP3yWDhZLjG0R
eK+qG+mFFyMkEN8jvgT7xFsX9BGBYGHY2Q6Y0gCYSYU7Dxzumo0ADxEXJbfGP3Gr
SPR8ipEWSId0sjsjLN+xjLPYR+VNifklev9BcGq1sHLy1c3jyC3XYOLL6dpEamAF
Y3Hs1wZNG/NE/WCkbggDuEGI7JJ5GH6vOzyqiCvjwjiO5COrRdtoGAtzvrcvMjLi
AolvjJtgf6kpX/SxpfP2/w+jJUglmfaJuvGDV+G4fpqMPQvyeBfnNRXwPjQbITIb
dkk53ci4cKNUovc3tRjVPmc1Zf64fehlrizkphnMcO7C4NZDoxViA43otk/L3HuH
cNR2fFYQQTCEntg+aWi0N6xV3lNw/JYpXnen8/Fw3h4R7GwMscW5CItzZEkoJye4
rrul+hIPRkNkvDWAcPEd2z+wfDh7zkdosoWblfv2DjAcQ7rox4D/4/7zP7ju1yvd
7zKQyThu9yFcIbge2otWt1UJamJqKlKPBNg6eMGb3PzgiRjaFygwNZ6SHloacRRZ
JAjI/kBO3YvbkGCgtvfKS+SYcYcLKxH/DTcC+tphkcJtobY/V341KHYZM24H2Ief
77u0myBxs1BXjLlP+3CH+rNEelNvk/hTN9mEPGxZ5Qh9V7O/CfMjzx2Qh9iYMWus
GnR/d6Jn26vfbKPvP+3laEzp+CrlCPZ1iSzm4kMyZzGobbmfAgnZ3jfkHlMXQ9Bv
IU0lXNEVUL9Y6TULBiX5pjnvl8Aap96UMjKtiCDagETk+sQuuap/YrdOTCNRh+/M
0wpodJb7xb8HLiekT5kpNPugW7kKWtvnwE/uQzFqbSyGYcUkSNUvQ1BQVdRo5L2s
b2Zz6SBewZZndgG43sHQVb1J2R6oyAZBdyei4pJ+PLFUj7jzvv+SMKFcv+pdqdLy
/4sRRYA3rJNid4Trjufs7TEvjzzXQJuFlAElajLMkeTJwXf0vmR7H+fG6iwbko7e
r6PEQVsUpWgHqoAw2feJyYlm93lMWFYdgBtU62f0x+T1kUzYKKCgpw+W8UBILe8F
k86a9N4H+RMUlVHISv10FMA37qTY5kNBOcu32CrZA/CiYiT5eRvgCE2Nl4L4gvGJ
kmRbC/LdFpuY81VLhPY8m4x4jw4K+AQElQh0Bq31Zc+kz1q2+GA7yiS5efJJ7n0A
PQRwiD+Z65z0m5wrDxCpRzpunLcA21y6hXZZ12IKQIEzgMBponKvZfuj36okC7m9
FLuBbS2UhZ4JsOOh17EnNcS661GQcNgWFIBGRfbpY9NkNJrARG0l5eqS91a/c0UY
LC2Y8/Ni49RREdbLm0YQSEGaR2nRyvQVZkuycQbHL18CxrJR8igaeeJ9isEXGXAH
c+jv7F49ZZ4oYv2hM+m2lWA6Z7zrq9ObyKpwo9HztoNxBftFRZC6/TNCWE2sZJV2
8Ryra758BDxb2jypMU9MRcuw5VDjJ+20XLKE0uPAAxnRMUmEFcGaNXbw4vBIwVv2
3NUV33XEoWT+IaitbXyBjhQt6jD28G9KxKYS1Saz2d2vdigLq6B7IizOzY4Yw3f4
JDltPGLuHprTEfb4LV0I/zGFoxcCxn0fo1eEpZobxovQgqdv+gscwQ7mogzV5uao
8Yp7eQzeW5HliNrDNBrBUme3Rkxe9n4ouo1mWj8deZu4xEqCrilGmtqJAbuCuJ0L
Zi0RS+MQul4neR+De0+t7kWUXF74boAtJHN3FEIpTJ00BdZ7nGH9S2gpE9RfoAQO
7zGhClkbHoQVWI788S4/UtAh30wzqS9brPoIELLgPwi70L0necNvfTsjP2zFJtg8
SHbslXgO7DQ5RQV/hwdJg4xmte84ayLf1gWMHyo0/7fVVr9bCtXLcoaDCU6YxVLQ
Np5bHTNSmbOM+W+BsdboZz+CnlbUOgOmZB99LcUOAhGfMIXgVhXL7gpj9+yMXNzS
FWLttWxJPyEuG4+f5bDVLYR2hEdzKJNC2KzKmgFn9k8knb83a8C6gHkwC20rzR+f
nXeClsJ+pHse8bAykpYRvs4KqD/UA9H/f9Fn4qv8LWRpk9y/xDZoN+dbR2BEKoOb
sGrAUJUR65ontF4el5XEWvOwOC8d2N2v2FZP1oH6/NrwBB8Ud5DXwnZ+Jw3sirg1
DhdfgsuI8BjOwtWWvRB8WGJrcpoHAOQtjRdm+467vc8190lmB5F+ojzqWFJOc4yY
G5XdSJdjJeYF0yj4nVyGsYJTIRf6I9sDYoVT2P+cxTpS4k6mYhuJTpvVx9V15lCV
ReW94/3al8TWtVK2w+mwyDGP+mRsLc+Oj7v9YImiJDVNnAs9lxxUzaSU4SJvIfHe
vpCNd/azO6j4pXKPtFEK1b66XPoLq4VM2xStqaKck49EbNULNCstWNNN59eOw+zT
cOm7i6uce+tCtlULXod7GIEe7rvnR63v4RYPiPLKHaaZp1ScLBAcpIM9hilGOKKP
zrbOnRLn2idbpPIG2Y4/xJgkiQGRF57568mWeb4TqQ77roEhXwgZRXPpO1M2qwtE
ZI+GSjkWD095tonBltymQ40odK4Lk1jpZCeg3OmU9C7DKKxSPxDGM/y5R9z8aq4M
DDEfkuMKN6xc/9I1op1rI+Lzf0/NZZS/W2D58/L0EZ3mldS5vxuOo4dc+7cD/b1v
7Q1s0dbYYfhMebnYxwwqdoBpErTRM3dZV9iKQuEr5QqL02ovTSnS6Pr+9Ng2LE5L
myj9lW0sIKT0KQGz/fGw9RvU4owrM3TzGe6I0b7JwcaypHWhk4omYOBl8AJ/2EGi
LYaEowVFeidoDicCH1yz3fkarj0D5QFOJQabHoi4xdkfhEieqKiNRz7PlKVr+mMZ
uXbIm0H78L4ypQOgwXo+Kbr0YppRzZVPMoDh8uqGflz1yZ6PRThUnD51luAW++QQ
5vmlZaJd8xDiEVLNukmzVt/X1Q0g0TUvftPoHkQzT1dAAOltt/jsrbapzh2WnhqE
DPZHDWIrkc/MgUPzm7TSrLkIixrPQnVx/Ladw7MdYQaEEmJIr2b/G6bQ3JuI1iVZ
xOcjn0tzQeUtUjG/bRYdVwmaEBttYbnnM2AHB7J7ajjv7BRbNBREdzBN/V1ipBjJ
VK8nwLdqWlQW/cm1yejlpsxKT5SF3oJEbnqB2qeiY18RpDKpyPOldWvsyFL9gnvG
9HuNrWpyWmbd5T2bh5HPDcSarcKhMgn9JMIvDOyx9Ro5z7fUSpEOcIyfi4HZeq+R
o5kb0NLTiSzHmsOF238lXmkl6i6R7mnlonCXUAG7ULhfO7sLyNqCEM42Ph9l7sUC
92UAhUDeLQPGHYTKltHksOcwg/w1hynKjkM2jWYxTq6YYRS0WuqxCAQYpIdMIz7A
AfgjgasHKyL3KBfG0xRoUcHZYMom2WMtK30aG38vOXByn4MXEF6DwwVoTjg40pzP
LoYnEF2NCMiN+VkTOZyjC5r88ZKRLyP5fiZgqpufboeJ8Dxl+sObo5iiO6/FjV1k
79yoZbJnQoOqqkULSn2ANaHeICgZtDuoDEllva/uHcr450YXYl7imfWoNQKBCvh1
SymZ03tOXMw1x/H9FZeBYhokaZPw7DLOXZEDXgjAviat62ScoXm7prwGp3XkOTkI
0YLc4TGkpZyNa3yDaJo9xPMi7s1SWYVgfxq/Ooa6towr83WdTrlnNV0rgSyqoZI+
a0U5o4S5w4SdTflssXo0FcC9hXxph5fWEF0+gMorQuZUyV7oCCDvT6oJ1ePO2tsj
q3Hqj/dpx8+DXFjcm43N+AooEagMZ2ivzqx0RMCDIMvRPv4LUUpWx83+W1BdM6Td
dxBmnGCE+V12Yei3JbErQhCSqfDEx6BFrREU2NyU+jJ7InmImqAdPfm3NKxZXvly
WkFKRrQEvnHsBQMZMG0btkFvuYu6C3PP3QRBE0HlfFcNQb+H9flXJc8d6sw1iYjo
NdkxSNX9+u9nfgidnclGCJmQkWRbWCKrajqHL0kz6eNM17pJQCeW7S/ymJ9dWjPH
7mszArYSRTQOw+ygtvJ03cwLnRmIh1sRZREKVTZZoSmYaFHiEEBP6gpZCRqnPxYw
gC/kIuKk6dT6vl+PMNNeh4/gTpms7Qd2WiZ/7HP8aSwIuFQF79z1JAIWJcZ3x7R8
/JIqkjPuHKlIsD0QUt5VjNy7ioKGA+KjRrS55jSEpxMfnFz+OZ4QVjLRQG6LPMVz
GYypmwJj83q1HSPZaeMdJTh9zaPN0QmfiZtRPumcPuX01H2v2KHbkjEXojExWm8F
ubgYXg4VSz0m/bB7L4KKMCn0ASZcY4zUqa4+fm2uN2kh6016bsVgkh8kwpZpjEEd
TeJtNfmHgLJijvlA5qgqsFuK70TheQqbEaXx3Madg83Hcl/bm9pgJMaNdtXOmgH9
vR/lCyzTL9yNFjQMHJCc8VnD2/UEDaHzz81u3Nw+iINyPVEsKEaNanoY13vxAlrx
GUWrgcZXzEigfC40IgrsT7Vm7xgJsBgoSbOu6+wwp5Q2RSwzRHUu3Z6QC4uxgnzP
OCoKuGuhWwhuG29kGhqSG9R5dNS/FW8DoEsaN6acNGUqbWIi7D5G2DnnVPE8jZ1Z
opLOJaenYiXmBjaws5f8xDA5Dya6rvxVjB7jffylXzNtnKkcUHZE7GmBH0E5cteN
COhxvK5lp1ctA/NvO+jwzdOJQDfRdfw0VJydLmlHe3XLZUyuIA/iJyTi+6/Y4tZW
vzVq/Ox6qtvrSwR2L/awemL4ZHz6IFA+d3dbpgKdep6Up8rwzYwKly9IiMKOzH2H
/f7Lv5Y/+hHZOjqP6OpdJAKoT1zo9ueEWJYYpm52AwxmR0UkJSwp8ZwIXBC4EuBL
bCChrl3u2nFFHr1Pv5gEAS6FzgrtRXOz4jpPwJ8FWz/+Y2VKIpr4S61dKyMkSWQx
02UGX6vxAMF2KRvZ2R3QBj5qVRGd6a9RYsIumLsDo8EtEe/Fb5zbeNGRGgpKMX+z
qCGUdQuUM4YkqeJeAU6SXbmyaD8H+plG6gAtEFJr9CeIGAP74kyOV2wSIWrG/tx4
DBMko1oMlpOZiGzO7ziATrvSM92cVMsOCIcLOZi1auxWjiWj2ZDlHuAWBtWcpIOU
hlnjrIeLD9cIRiCwi3SRsA+UjhOYjlISnK20hpvZmxl8GjeBgKWa+YepaB6nCzcr
kLYioYQ7IoMH1bqLKXMfkPId27onPZHlZiHPuqShORc8RablzjiiqPV/LFGraPv1
547/LIgDHH0laKCawRMCLCMvthQ36F97pNStZPd/7kFQM9VaLQENK+ndW3m+Sgrp
2sEyJl4zi1GIjlbeu5wD/tc6sAn7tTzD7ytBNKXm9+hzeZ7r+yatlhhZelTYn6ea
JSwpp64yujvtvd7undKTefMS3BxkaqXpYKpR2VgqXvFnkLVy4Yp4ChRdAuDLR4lA
V6fWt4o7DGLqIwe2/xH3EANJkiAmKIVD9eu5o7r6gnIYO9hEpOtJnGkRQtSiZ8bs
g1LpSaaNdDyQzwK4txxUeE2BWEdffhAmTRZAtqrF8YdvSNiPneS7eOa+RsUNY2m7
8w2I6DTxlfnpVHuCGEYEwT/8HjGxoUWoZ6p6f0wSxURXQj2QBUE/XwWd63oWCwP5
QaQzFHJXR26NzGilb74Xm2W8qEBY+Xz2/3Y4uhybSyMVykLeOBb2QPVmFt3dWkZG
UYzqvDeIWjDi4ic8jMySZPzKy22dTb52wOfOlIwMW2s2vkNXTdYcYGsoR/+7P1j0
gyk4PsSo73hKJ3y7PJhkshKyAYZssdOBXyYCGfPtBIjyAftlaGDrYPSlKyqJ9l8o
bAi4Po3HXioD8VOwxBnU3hlVx4ifsARMm2iuSTOiL97GGZVCLQmpYfa+EfYX/aMQ
0gV9nAf7BSHVmLFWxHBaQZFZp33hBQHWLXg+gc7PyGExqazn/Oq/A8ToN+QARgxw
R/SbM+vNS9i/89OtBIsMSZy5EobKvXeeO6hbWOSJT5ZwqDoXtoQk96ySVF0HSA55
bNnis3kw4ADuzBpHILitaZDk/uhevt82qjbZb5Pivh6/bewp32x3d92MmOzpg0i9
MSVdv5/5KjUhY2GUI1jqH0BtK+WG9v9pyI36tRMXPkChdh10enNnAxzs4p89LCKo
hXLJkmqi6kts9CNrvrCNF6IpM2iJzdQ6ESSh4f1TRe7LbSPZLuMjt8L8amdSQSvE
PaySsxYyw+ZIT4kry7qPnP9Q5Os8dUQOPMu/WHz+oeFtV9PTjiJfuOt30ZqTeXtA
wYvdsyPs4lqcSadkQJrw5cn9qg+O7mAExAGo3s+bm539cgAcEX2iYeZP4N71xOyO
mP/EK/4lAd/UTmJM2qJfUl1w7LOl7EQkUDYEsnCZHpMHV+U4P/PK4HcuaM5fQFAa
0c2aSqYJaOkCN5C1TcQE69qPPkuS8mMUY6EoUFsq/MxLjZKWLg05toty6ikGw9aF
nu2Yv4GloF15T9qQ70jS77Kscow9x/6qYHcZ1F+UqGpvnwJDOjFRww/IHX061MaC
EhcoKwkQudPSshrWlDJJ2vW9h5CwPIUWPY4622mUcyXJcSWLAIZLRkQ1+nxevLVj
Juuv4wM/64Jfk5udOMfsRPJ+OnY0nAi3+bROhSN9SaxpcqqFGzSbKEoUAL8Ds0xD
yO7gIEkt4NFEV5VGfCXmEui3Cxilx683pmaOjjvzOoF/oSBEZZr8duStGuDEusn4
je3dOyoQRuPzpTygdYvxGHZ7r4D++knMCXRYkxu7uN1hktwVxVXYFfkudxNxSIDl
MNppOcKb7uZ8P82Py7LqKyByoYT8ipdYAfRcGlAtUfT0dTJcuIgEJuyxhbTkoQ4a
b4oXWgULs9iRu/yUkO+rGcJ/e23NSPUEKVPckR7uTY0jiDSJ90YBk67W7wNbfDVY
flMQNbYfLilYM8cGETlxK3X8Bga7UBMOd2G2FlvAF001AWl9/T38ZHU3csGG3KZM
gZX+ChgE1CKChA/yPM/Xf7YHP84MHRmxtStgWhDSK610Q6Qv66Qg/16rF/up321q
5qNfaqRtljKk+xozz58ZfM3IfC0knnXNf+qwPA/S2xBxFnA+XqstnGY++R2GnMtI
rNapCFee4EhEvmdDP4X7y/7kMSHw+kns8BxNKb4TYLghmcZpRaDkZsVhyYSeaNNb
9LXEl6II3i9d7ELIrBSNiDtr+aokawMHWcBBkj+NL0JdAR223MniqaSUSLs6d67o
5dXHLtfzS2kufTxBX2okCJjRebiXpetD9sTzk7DNCLm5oCkDp8cL9FzNh2sO9Jrv
LgGgH5b0CgKfHDzspXh2tGUBlrSvHuItX5GZwuD3ywgm0liFAexaT/8n+6uOUdOg
gu3modLAc9WQHay8o3Ktp5SQbm0gkxBqtYgtWTmgnX/gKuqqJit6bpimLCG9vtxN
8gMhbUN586Texr46X2PgwbEquvJx/wIo9R1lMZqIZMC4jMmSz33L5O5RGTMKdwQx
/yvaP4p1K/70AQPEm4SkBq5deuXhsWxqI/YhueWZl0jb3X2B52CUI2Q9XJivbphG
thVAf6szuGBhGXFcXuotNs+u30rgkr6bYUtBjg/FbXJ4VJob+6YNyehRnM6YwSzf
fV0YkyRCpAAWOI2KzEI6Xev6E/hkh52itY1b9SODGPikEW9kWlyIa7BsQ3H4WClH
/u0PIzIg2RIJlFQDiQC2bPFJLnt9xvNXASjFQGn8/QVyMxWdPuqQVDyC9ysdU6AR
3KxsBKYnVGZB9/yxKtJv6ld6KtOZiTlAAvRFO2ZvPQg4UVoP1aGP1CTUCN3N3P48
ZPww+tjqo6d+EDA/lrX3H4CicNLjrUvrzTPzbOameR42gjcly8ew22Ef1JriaGyq
tXMDcOZ2IVjrm30NKWQc67hoGYmBgUnrQ/P7vaQ/0WVOWwV2pJvqB3CH5zU6XcpS
BRipSE1Q95n5qEeSoiCcaKmutivRKwlELnwb1bTZA7en0h8KQuVzzagxxauvFywO
s/TreHoXzJtth7ptoe/vu4r1lfNE7ZZu0JBEE48IMlkkSIAhhgBjqpnPaUzGBu/q
9InjtowTb7OO5lEtwZP0Csy8V+JCUbz4xvM48X+dwJpHS34COdrAhxQBOBFTv9zI
8HeLEEJCzjfqnKl/NCAshJSr3JQSUMsdxpF3Qu0f115IZmBuGsZ/AO/wdw34m09f
C4vbaMMjHzDK/Y903RxKCZqHEpajz3dPvfnSkogvGyAz51RRHAvM7HrsTSGMFJ+x
C1wHTIkzUadiq5E39W96oAzJ4n2G1ZjDCtRsbKiP7k7Ol0svEZRvy/n84/0MZ9Ti
PPgjayzBMlPc0klSvB5GFWRalOpGYdbLXgNfC7eX+/063yKs8KrK9Kz8yLf8GLmG
vgBY4dEhEVqDxyWomdLqzZA17D2HqpIut6fObYi9DvVgiTcXdMcoPQUJqi970j4D
+rI41kMi4w1V1H8x1Kpsf0ZASJJCM9Rjqt690WWFbzFEsv495ATftU0uS8Vez1Ht
2PsXeP6gQGl9m/psu4zbODuKPaGGmTejC4FXTkd0tBURanM/gMISLdxscXvpGyCz
fzzqragE4fkOopRUrq9k6BnNmAT9F5jsYYJ/EVzMpBex8Czf1+e29ewEP7vQHPcA
wzedIIEeHjQPkwBJvIG1LyMhncArd4p9x06TzseVfmVFaTRoFrfdAzAJT9SM/3mv
voVy49jCu66Lx5Uuv5EA9eWJc5mtzLmKxlkBzDv4MjqoMy21ncXD2irC5hBz+3b/
KhB1PctD1aVyUCpDSvZxMIQrs7yFPOWpYjvDW/s33lf/EJu7sQ67QdzMJrbsQYh5
Mdg1LlovTiwksDV3wPF7XPKaWAB2qsfLP4hub61uqR0FwbY2gTvLqm5x2CJYfHxl
bR3ZaYlMu87cIPe/ZjKWsF4Qj8S9OkMU7a7ykPY0lH51nWKu15sheDfBYC4lPFmE
TL7vFrwGNJqF+nnsP2gOJTTvZBYbNefW+MnLV1P34G3SowT5F2odIqeIYixcJTbe
umLVsDyPnLvDw9ps324GSo8EDIS+Y8JSRQvR2lhIuh9o9lX2Qy6IVWwPO2CCaNAK
FWDrqpKk3HZAZ7T8/caeV2vg/owgfOBRAdogMyykG2vl8vDp+gnuxs01d1w0g90W
lRRwux9zB4Pgbr7Mw2m5wq0zBvhEryIdoP6CJv3QNvriYcr98FA3XJM9eZ4plIW6
pCusJknubczpYsd46bT7Rj7UxvzQKc0AS5ijOZBrrcN83PJaUcRALeZWJYvDn5XZ
3en2z106QpvUncBs8FdQj/ZBBPvb+bDFb7rdEBaWaen3x1uONaXAeZAlrCElovl9
nJhzSL1wLGWgcbMp13x+SEbJA7cXx7HLCiyQXsRmAPiveETx2bAJ5TgAhTUELjjT
ax2xk7238Ev12N/zXP3CnefQtxXKT9ij8qH0qGsnLVgtRtlEi2uxr+VH+m0of0ce
jCsyptqIrVaP2UCbOJPeOaf/E3IVYOGtYlHKjYsJJWuDFS0+wx1yrFQQZUG+ysXV
j8YdLtzw3Trz++aN9Q1mRHYKBznoVZTcskoJP9VEEpUSvG4oplOLYsJ1zwPpbKGi
kD40NP5l307z2PPSpWDEFi8aby/Un+cfZXs7W8lo6U4Mxf3O9hAi1HySaLe2JD7B
P2rI0iOiQ94a0FKPMtHZ3GF97cWdhaq7X2UbnY1WCIQbyYFDPE2mMOq1z+xl+5e1
WWcmceiCanAK0xsMf3zlwa1QHR6bFAOeum6gy72lCDW4LorlbdHKWLA7uW3TBB/6
mDJafyfx8CnduApxYgxeOcop8McmsCZlf0WBIxI4fxRtWIzLQhLTgejimWDMk4yv
PtTjzhzXd/S1t5jLr2/4U6hdM+uSwbG+2AD0REvypx+PN9xtVoWcL2Y1cWcOrbyN
aHWIKWJUs9LYVzUG5oswT5p1FX1AyueSSdpCOPa0R5BlLnNMomJi7N9WbNiBBMAF
BkZdJIWVoHrQNit2KuO2L7BID9krpWM/7faWQDn/QsjaK0OftGwuetXvzOSbzwlO
nVEUlMn9GoMi92JgXgeBwWWsoH9i6m+n3FwyH/+1fcT2FeZpt4M5ekijIUrnkVS+
HBwgqK854uFBW5v5O/mQBUHuSqpwAzzTA5ZqgUx7KHJcvgweVmgIm5AgeyMYUvXG
AsD3fEqmkFOVeIhqrcdQymdOhq3O3C+Q09tQEdnQxifMIIEpjhyveouoj1La/nrJ
3k0hQX9gkV6IhSJyEnarTctSs5pMExFKU2/AWaibwhNhgNIhBokPcKcZ3EruYVBW
8Wwa4JDGQTxC3ZdAedDU5ybxBB5Wh6GbdLWGI93MeQ5e+3ErpgjqaU7kEGGs16Zp
LLkMijtH4XG1Nw2RpCd8vZUEu2nxnTRSoyIk3i3W6Uji2hz8ejfDZSTzbHLxuLnV
Q6UXifxu/tZBnMmhyPYqtQJ0sBGiV7aQwZQH/CMsfJHMI0H2lOrtcwji8v/LNYHF
hi1H/BpJC25ILGIk65lFaMYhspsUPYUW9F/rLf0A0igV3FxevZtcZfpihWrOUdIv
1ea5mhqHtZdIvLD7MN8dtjrwpbs1fX/opecucpGVxysC1uC8D3wTsboRBDYG5QNf
rCjTlZphEvCPw6DLWIPY5FleP6jp5HpDSMmU06WmL/IWQFyaEpMHanfYinqahh6j
PzZuH4HIv3eDfOM72J1X3ZtH2kvVJgQkPMol2QKQoRlzDfAqwdAWf4gt6c8aWKvH
HUGdL1T6SzRR+0z2UDz/HVYjEDK2UVlUZLGKLixOAJQnpODutV6IRvyIoeY8jNws
Ams+faGx2MrAhOIoxaXt+CDCI0Yk4rRGR27vnsysU+N5YYvzhPhDPA4XXdWPhuX/
kyjE80A6lEGD2zJBqUvhyTVLL1TXG0OoJzzhBBRprdQ6lVxPGJK2OJmVbfq1qNL6
XOMFbEs51KtUPqfMaT9F0GsHtfOlZcAh3YuUfkgdGLzGZsjy8PdoYkUZdIc4m3pU
phHAnHIa9VKhUSbK25AhB3VJ9GmZD8bcFcHcWUj47YBi0wr+CI0VoqWElsrWnVUZ
JnLungU1qTCKWO6xWZeZMDiwYZg1tpOoSgJJynwDgZdeldD0am4HjBfAcMPw1fNS
qGoE8K98gm1UPfuhB6+IEUwLOtBZl2sjD6utmRfT1K7YueS5OR9x3d0cKI0sg8KG
CPC8o7bQG+vL/QXGBvykGWnKIirZjft6nFE3L9xoGoLoJarIMA8zpDuc4jkt9IGU
GV2wN37gUy/JmZliHx1H4hAuEidqm1l8mFGEZ/QCmLSfvbGdtjV0zxDbxX+Zd+pb
ZGwnO9jZdw4HWz3T/WsP9J4n5B7/wwVyHER2Wkreru/dGcSSW5kM5K0rAg96FrLG
bAUYepgSYATWyGOYNfKYg21kf616jhNaV2f8vkph5d6uApNWhqxzv//kHcW4+Ree
BlnCA6u7Mpaa02TBAuhuT8xTrdwBGqLPQ7B4KEBscBBIWyQEUm983XMTeYp/LxKn
PnGECdyHS2Bn7E3d1QaG8VFmguVQ5zATVDj/1ud5FBcdS4hiw6LWqGIfI03Q7vrt
3xeza6dwmcXZagrRQhKm+B64QISIN6jHDK6VVkvHHxY93p3WoFv9KgSV2t4pyYYL
zem7j3DJTa8dppEm5aCLlwZDR2zhN2aR0iFk908v1e7F4AAzQbnIzUvUpkl+pw2T
vu4zYMYNZJLDmhFwOZk4KVCMKAIkfr8xpugN9yOuAHUXR8LzxoaY/Bi4E+kmDLrR
/HVg0Rg/wsZBtkCGu+6DpjRg3LCHts5NdjauSDzonCqKMBuik5dh6XepAWtYqX1e
tvzAbouq1el3/B6Sozb8PuepowxIuxglTO75i8nKyWm5Qbh7irUDTB1+PvRHYiZo
//fMBI/lXmxeEcC1cdBmqqDuzzvGxo+vbrbZe6oNzv2GDdCD8d+f/UduPSCesHCd
+18bDPT3Skst9mQ5pkbN8qrrmlQhwQy6p7IJf7xZkJr8leriJ2tP+azsTiei/f8Q
ytItvmKMcnpj5bAAvgpr2mZybx3/bqcZDADkI6yKS08IwXsrkRBsNKS/O5SImNZM
9td6Nih/8ZPc8FGJdh1uf1+DwFlnts4mHlgrvgqaNd2EbfXF4tfiLuRII3l0axle
NThQVAzbTfz6Sto+srj/mH2E1xb9aByeJqMYAw2D41M014IQjqXmj9dwxGdyIQbD
goXfYNSYuK1JUbMJMZtM9pN0AAuif5T9Dq8WoiypK78cASahKT7/KjSobx+4SwCg
tgo0GXwtuVKw7862MVJbx6kUwoIuBnTNufKjocC29W4MXZBlMn1qiLhGJtpDNBnd
JOdd279CP+V9bYfaD6VBCGqVoCipmzCTf3HhfJCHdC+vSw5vASvtczLa3+MHUIxE
QfmOXkomG4tSVT0Fi4DA9KO9u6CGhsHM5KFa0q25M7v+e3uWqkgOLMtxuPjISjv3
6Xgpmlj0kEezMG0axX66OZhGppaLGYE0vX0m/wCkMaZuLz8IkWNKfA6bZVFx34Gj
MTJ4ghpnbI0cbM4BHFlAfnEu7s8uxuxAyblzcV2gKOPxwP/zOf7ZoM3t7NAGLrWi
93G/iaKBvNr2X2oiZo+yt/Vz63iimRRIlVI24C0Q9ezJU5dbz6na9iyd4fPJeE5a
zIwrnh/AfWnNgwZRq6g1HuKrGmbJtYMQAoiCp2Ws5AN9tKUAxctz9ub7o65eC0Nl
T7Va5rNLEemZlo5Y4pHv5fhAJp52VCIrNBU+p9nNoFI8OSEc732naon7J/bvki7Q
GZDzXoJMliH6rI/g7zmGkrmyTCd3erENGd/vz/KJnqL4239W3MTWGbqLeNjo5KVs
AVN99MDjGlVJFKD7W6RxMrGvRB2BOedwsKxcv/yfWtaXik4nQNfalTuhKJhWP+eT
hfFXM/0lX9pgPDnoIVWc9PbqvD7Pldowr4aB6a4ZJwHZIqgufu+vSqShJlAytXn7
0T01UkspucsWPRedZitt+i+faJxCvIUqeg4RNXUz+nmgdQiD0IxQM1sUEF0mowDh
OcyUqunvl50SWYVUoIHkVBxffKpQU72vwH/s9zfSUssxWyT5w2xCJvMYqIwySHdT
JgKBZA06/9+vpPdD8tCQ1k6TIuweVd/L4vuz5PUR0laFTXq6dU8ZizrxJy0P89Sg
mQfULkpYT+JBjek1b7z6oQoaRyam/ArLIKST5fKeiCXyFsDUuEuVuFaOCR1QNl5S
B9roQzV/fK5uPzYPbprUd8ArIg+hdYSfPRH8TId0h9N+DPL7oTGWCfZJrcJMoMV/
076qFY67POvt5pvknoCDSElMzUCAUESmA4VOGT7Wk5j5pHNaOc2pixW3n6Xhb9gl
6zadhgHV8/ticWm+sUoJdhj5RryGgq7c+aW08G2wIywgNXrXtzP7FQwUyIADPblE
pnoPjaPu1L8acevQHNzx0C2ph+/72k2FUKGj/D7fDhT06R59llxs7FZKz0P86qEW
sTwe83LvrJDGl1hU07SlxsuyjRHXt2XAS8NdjLyGOH6raNWiCLzCTR162MISw6vP
0w+PvnEPmqGicG+ZkYiAnaEK6IpqYa9lsHPPryWBmeR2IVjAM4o3XOTPVy2LqFHU
9FGv5wgfxpA6kJcNNOEyjM16AL+s1QItTy9tdaXREokmc8QU0d5uuUS9v+ywaTKY
spdZ5StnSVbvqXz5rEk68Ky3RFaJQdTYn+Kv/Aj3+L44lUSPC0ypJ6jIA51TDMkP
xS5jG4NQ+85+pmTydjpoBacOiJtatsMJDcvt95SuaodeQyL1D3TwhuzW0H6wnG2L
Jiil5pB7M0rTFmdgXwnbMxPQKZhpefGHEE4ZMx+rrMXVJTyBLmE01kRkFd8BrvVy
Sk36UqxLsXFAP3kh+zzC5vlVVIkls8kGVkwsS+BW0cr3JGbB7koELShhmWquLUwR
9ncLHQi2qsy1QVBrhUz7fFxGTDIFuJcRgS9CYalqDEHbPbITBngjjINgvqFnBXhs
AL68tqH/fKKhbiJUNruP3U/B4+S7kui/HtVzcMYR9Cwh3Ti9T67bKb82u5oLf8kI
MAT1iiR9RhDaqXtfbbEKwPyd0BCIobTZi/1Dk3H0ugzVhW2mW1QI9Q5019lz22r6
QsaYn6ViG1rYWcDMnZbbpbyD9ua105ws0JOUA8kNz1hyDHdnY5BH9ZafAHbOxf80
+lOvrzGOFEb5YGRGiMD6v2zzNYslVrkxW3vWRATo2G5SC6skbWHDoBliQvBBy8Vv
i1F3PFIgTT1xNyT7otRR9rsGSwwSgh1qGHd1fExFX0XO5FkQHnjX9Ld3DwBe1ol3
NFhv8yZGfTgXJmcUsXw5GszQXFPoDhKk1E7drq4rSJtCnnaSj33dELiPvzqDsBuD
yM4FU6KVvRz26a9TmU+5qcr6yJ+mmp3c2DJ+cfmNiIDcjpSziZSMUJ2yoAEp1Trc
Vy4iMEIpjDzl8U49y/nJiFBnNuXiABzfjOKNIE9GK3KcWi027wjSAFbfpsjFo2RM
c+I+h9/NFeiGyqI0SzjqceHPvjyagA136HGV4PpZVnXFBKnTJL8jO1WU6Yrch/fn
U/mME0O84zSsr+Ent7AXOKZdxY++ueZ4kzSFOKwFaiRwFJLoLEFOJBkQWtxMI3pG
gYeFjhmoky4MSQT2lVAXM6sVGwWI3+0ESNdovKKi3q/HAtxSKGx/FrHeXQW5qjDP
viH8vpu4f/4KuigDLVWfROHW7Y8tIK4RhD4jkJ/bVTQyep2HI7zCaS8leJdAroOu
aWX/kIQVynulaP370E054QGR+VCjLaMLTjTyBFfoKOFyBhQn8vCEhDcMQCYj7T4a
G2CvBaMKiCWvEsKAbiWe0OhHlZWeg6FvAkFACmnsMGQkv0U+xeeYmMlkTIwU/m6O
alSHog4KBTYJ64dIXP6ET3ox9eZredExByKMBNpd7041MiWLj8FM+kf9q76RcUHw
+3u/P9fAVn6uQwxC9b8CSjZA/v+hNRs7BW/U1l7N2njYUidfYyy3yip706HDQtpK
yr9LvZXvB0W3JUFegks3eyIAOo+XK0JDoSjQgeHe+Bb2TThon8teHCi6h7E6QUNi
d8A0vjpJNiYr/KH5krfMOvCAjfEI/gK0kRV9CntOGfXxBDFej09dOnyhqM3A7DPN
MCqe86NHNPQa9iFI19o+Dwr+u2rrfZw+zYJhpD4XFxYyILe2kyjbTuPhUCyhP1sq
0DrCSlbrQ6LbBVxkwB6fnTWMZuxRVETis8WprRTDX/t0ke1hClPKExISkVxuKhDZ
RoA2wJm6tDEKR55XcdpL0q0/ZG7G0e237zoCwpnBVdczQlwN/Qde+hiESsqasDrq
8lCMXYtMZBINjNZ18yBl0FXeam7My6rWJwj/Mu2gG3oxqfr7LCBffxEyPzVR7Mgc
6ojmSZNcA1eKnp4ZnP9T1fm75JNccnLGYG2CyJXtO4k1f0SdZBYGi6MSKyeR93M5
N3mQWSSj8ZOSZXgwcKz9Y4yunnMWLOhFfgsPWMRws5wnyblMX2v7VAmHFzjmWMqe
6l2JiyCCHlK0AxvStj1dUC5EyyMD+aMN1VgJ6SsG6y+wyWSi83x54aADK7fEAbM/
EcAnBbC+2EBQZStMjS1iB8g25u8cHM/Z/D3JgYtn/3hgKit9PKCRANmV/LAaHg/E
W56lgdB2cqRXKqfyL7X14StVTg8UCXVP0HIxAGLw1dBLaZNV/QzTwq+5ls/h+wXL
i3v6h+6EkA+sSJXxgCyvFuksRrYaJvhVya4jGCTPyJecZuqjrfJXs5EBjFpDDKlP
cSs/cLUx+5113841UNlnpv7ZHz0Je3vCejtVqO87lv2jj4lyZrw9CiF04XJ7/GhL
/DgZnCRh8YuuBwUq8Na5f3BogpJNbylkIZ/VGWPjSI1dHTekVizsLxY3fGxywTI9
iZqsfJ3L0IHHFD5Ds3Hr0sjOcX0eRIM6mumOqGQCW7lQaMwZMM8wgzD1soROKhZH
VlGL3YAEMJPN9P41fK+Ak0U5NLsLb3tAS9DpLpSjTiS/rX7BJzcZ3/XuZc+uWnSv
6+aK6qzS1bJw0MuQ9c7osWrSLYwGwladi5ep3F2eYuDwJalVgvE46s1vSEROJH3M
yKBgon2SFcH5KUWBjckd/36DKkfhogFonOL3wlEnJVgb/mNCxuRTawc99BZDJiRb
fYFBucgnFfMQNDTez5rJYqwMsRj1JFmconN8cpjOQpIos0ipP8skLNy8ZHFr6yhL
AL+SodpSLVNUab0zbk4bzvIzRuS8FVmZma2Jmin/kDGvDP9BhGvfz+Pa/5JLDBKD
3/Lov9j2hiZ9OjQuttNTE9lXSdt4fXq8RXXiBAYgEZ9rW16aDoThIBpdswneb/Rn
fMWdm9jHmwO6dOhZ4fY0xheSNkFjN/D0tjRnNjpWyXeBHG2O2W2NcFW/ZS27MfDk
9f7SCKDYt6SqwYeVwJ5bsA6X+NctJYyUHpmi3N6V2MkPMCiehHgMzqmF0aEHvt0L
egV8L04mR6/MkiJDRc2+eyo+fqSeSp6LBahnAyVimM26MR5ysLlsx17sguy48TTu
uKiSzZKqesJNuaY9OXuQamo3O5cq/wBUUfSo7FCR4lSyKRE6qkQr/IpkYh/+mV1l
jx8YnIwXV6FiSShhGCC6/Q3Opg4+cKTGMdrpvUqvqOWzA3+G29KATbsKkpDjAKxS
PTOUU1hCBZwgDCtCsyP9NhiV0tvaVbBC96KR5Uio4P8f3jQQPxngvkpUgHEOy2yT
txitil1nPj1SAutSwTigEgfH1vYCWVLD1klk76EgGXvqpj23R7XbDJaEYFxJ5qv9
6ts9TstxMKqPbrQybkyyuNLEetxaKCgjkTMf6vb2EiSNalPG5fRj3qyYZmNcGVAG
gPL8NqNE86cgNQHbvvCNFpMG9CtJq4QnfMF3NiA2TI2vPvSFLELBSDtP7Js3jpx+
+3kSgIJ4ZAcUxD+Apkv6qmOz8WnQ4w2W5nOvqUt5KD0g0sF1/j6Hj8Ak1MKXPNf9
oEylgeyftVMuyDvnoR5QFaTDLeryT6ZzqvmTMM8+Ep8z7pI5NkX8V6KYJGhiPgei
IXrnccD9f0r1gbg7QxuJeuP7KnNMjtXw3NhppKfkt1Ef2Tzbk2TNKKmnSBsoFG3D
Do9hcPZQD3wgoQDY6dF98QJ04sCVmtZ5+APj9SOnvycEMzmxB4qltJjtxud4bBq+
wwLhv9oSSkqeOY3p3EMg77BwJxIUJpl4Ft0FYWa7rRpWxoxOBwYuriu5NOuBGFtL
bmFEXPQ4l3VFb36Pf5FJC5Tp/RZFY9LEmEdzZOcZHInAszmU9Quls5Yc1hI1RfDW
UcLUzL1dPBR8IVc/ccTqsWPw/WPlgxUl1YBv3HirPuiBZyMvNu9R0mg3QWM0sfVD
IU36H0jcP6W4Eb9K7F62UcPQPfiYLOYTBo6906rKuPOea137Fr+gjXFtKoqCShKC
FXKi+kTk0EzPpZEhA7/feMUI5SezOIKYxfQBwCdoYjaAHZXNEjTun5h/BWkhf15q
5wXSQn/7N+euqM7E7AARIErLRwuPuXvnIdCOM61TgV/c42KKCBYm7sewu1K+uaC6
8XcNMYiAR/eXWZc778RkhgU9CfV+bybKJzT5Xoxj7jZfG0Fu7FQHybDVF0830Ng3
DMzJszz8XuujEHhyW9SVviaTGzJcAYRAMfWmV0iLpewklsjBOVkgpp31oGrCiPVy
7o2P2e3Gdv6B3fv74GecQCMbStDCrlnPnmUUL5URYPigE8n7kIxNKK745LDILMeG
mJ8eBpyBwuaNB+X3qCC6riLuFyp/6IX8wqCEJz4ujeguVM4b7BLp+36BT0sUqxxJ
IqfIKAvjtLgWienL38Cr1tZzk5fGKKdb35iZZm2SbYnAeWYOwkwb4rMWiGMQuUmi
mmGpg9uFBO4sJx3M40HaZkFOCgLfw5oRaOBgw2C9fb18PxxdyjxdnGjD/cadVuQB
ECckk2KhvYOyKhpzef9mfnQfrpj9RQqHkRGx/5esSsJkr2lUoYzkHfaPaUokTyCq
yAwC4yc38VhaU72xZteGOFPaxRxZp492HfS1NJmyDsu5bKXTXYAH9jd23mJTJsvX
gtpk4HG10snkzwFYygAG5cda1hNUg1jX+U07oduZaASaWGBPeHULcpdvO1r0OEVX
sTje/admgXz4pX7WFukWGBc1M/JKhUdAW0D/LPkNx0kmDaac8FBkSfdrTkeC1sEt
CnMp4MBTy3GbdpNAVFNPqxsHr+DY4KZdhYkwaH0sNv/o5q+xnqXVZzFNIE43Kd2l
P4bl5aCRDLjd1el7TA6Pakd67O+LPHQ8iuNTkNUtebHZDuNDZP7bPM9dZyE0mF2E
ZHETGyBqHsxYaRAeXPOREDAXTjgeYgwaSV7bgDzt5GwIiUqNKv6dCwhpgxS4Dyyo
JwUOa6/uY5auzKMZPwlY5Nl5ElBAiXCiS3zNcjWSScCIr9jKSsKOecogOjd7vuQM
qX/Xnb6/K/dInTF6/Hm/tl/J56a45KEtr20kUUN+dzD3iPtCIX3ZuvbKf6lznq3o
aeg52X2cFFLohnEu6L6azVOI6m8GRvmBs1Ik2OnqqgUoZSPMXair+nApYz8GeduC
eE31mVfFo8vFhPChsfQEBmKtvmaXJchnHYwgZ6h0a1bnz9Os+HgLpprrc73nky5W
4eJjJIebR0CzTXbKjkahom+OW6pXFfQjb3vBJOkKsm/ebPdiQXhBOfzV4J6a7xuv
IZEImEqJYFhi+w7bkle3jm049N/ry2hHqXjpPGdzmzyXAGOnwCXK2Pku7CEC1uUV
NJbvUi2DHuBJdwVFeW/5/AtIfz1fNLNYVCr4SytQc23T/6GE9QtHG7xE/6BuEXAv
28Zxj4wysetJGE5RU5//yRsdWyhKFhhU56mcGlq+EgF190+FgZ1I5e/4oqrpXzDv
NfVWS+hLr7qtJtS4UMY8PCsfLOs2yhSifTXOGnlGG54Y+7sHnHPkdGsNb/luH4+L
hIda+GjZ4OtKbZIZo25ho7/QXOPVxC97mkpIV6Z0q24BkGoCEN2MiZe0SSg+8GjX
K4NzFmd9T8BF6hv4qNwsSvofHeU8PCLAlLGlHFzve+Bk/lKMrcSf1pp6Q1Ec4Muv
J1LL1HNVrLROZs0dFBBgHrybD3X6gkZyZ4UqouXZJZT5Mtj7wBpf0qKHrbCyGFF7
DXN+g3lgbvWw+XANOreu5hVLxQ9vPXfVzaeGqjhTQjO/tfq5fSr2RlQTdbtQ+7x+
0mbsQHOJkgKNMHQTBax4IdYqge1UfLq50ccor7Q7Axbr/2gvoJkUYn7Dnhz8qZgd
2c95NDU4WvhKVUDRccSTyWk9aeW+/CTsH+M1MmjobuX+Aryvjfw+70PusW5tQ5dE
Z3B1pcsL25Jj3eQbdyB+SxwELL5pp8S/uN/aqFbZ06oBT9/odHEHzG+9Q039OTEj
1DggMFFnhyfLnGli/oyc1cDkft3vhLVKPNZT5LdIMUioky/cqFBTys7XW8ih7ffF
MCoFPGg9O+wFR0VZ+U9L+snmvF/BDwrG+y4c6yhfQASaQrhnPiCcQj4ejTXW0JvF
USz/NyMvZWCucS1z2U6H4G351SVvBK23SNYfgTYvpxclNn0HYLKI9nuBDLNCoHz6
J3nocqDTgnHdslHP4pLI2nUl5HkAhYxfgdWizinI71J79d+ANYROWg5z6oIkKANw
7+jOvKQCLurDXcRxHJ7BOVCsz57vJSSkiIDR0g+mloov7ay+f0RaNfTeDdpJl71e
YaJ9lr5wrsxJWMLYmJ8nPbqu19Xmp+ZKBv3UrYMrosKNBW2PuLlKTVmMED91UcbR
euwXGwgLHmMZMlfEERkjO6rbcFcVkPGpnXYFbxlBRf1pqRkos17CF3zTFsutpXsV
ieRy4V2qzocJF9cFWZBQT3ZbmbffpVP/nHBzcgdPtw+PY6LcMcKfgd2QoWdTuQRh
ceKuk+Mvo+i7N3c58mX0FLXULepmcHDa7sJ70xrwBicUfTT9xE/NEace2Xoniibq
Rzy73v1/bLDQ95nAo/AkkO6uIJh29aC5GoG38POU6eweQEBVd5HNsaxHISsyHIBA
NOG+FmqMdpCVfaU+mXNhaUaKDU/zIUgUnOIyIdY5ImPv6u/1B6xA/EhFpu1ETU8c
+sl0uzy+bkrfXY5wQ5eR3cspWZWkfss5PhVwCkSRYbWx99xQoCHjU1KpC2YSKu6V
DOhE7w932Akqu5HdHKTUmesrF3ALzUmAQ0eVqF4iMYAhzLqmFRai+NhrU5eMyGy7
aJmK+sPRtfG3lBYgyA6nH27JswjgcvwUlxxLADAjzK+AQ5LBaYBK7dmUsWUH3ZTt
PTmwE7k9AxzMNt7OP+w3TRGhtFpEMfaRgNbrnWU8TJlgWpZbSEDw/f7jfqsNQiya
QF937DWqou6wL6D0RCGzultD3WdJf2UQdspL2cy2gTmkwhephGuQedL0vBMVsmH/
L/1I/QeSDpXBK2aJ5uju17+drO2Vdu1kPwtG7uIgCc7H4W/47RtZjoP1tPJlUtFN
I6dBV0RecH30/smR3NxsEJUbogztmIcXIM2cgDY6KcaZ5wTG14RD/npsfGDK5Jk4
NxHd/glSvCG06uKGFBJdZzktg2fE1ARj7NZYk/JdxQsfwwJ273mEHEYGh6vtl9IZ
B01cPyynxP8aLxutyJBBXz1ft/MrxPKeqE0JYEasAxu0u7kvWc684IeGv+n690YS
JcXRi1T74xyH6HhpPwSoUwMbhnMG5c/4bGi+tEQPV3VH4dY3QFUszBxF/0mFrISf
l3Lg8G2o1fF1gOWHQUu6kyF1EyQJQfPrHDI9XuqoHhfRqr36bp86hs1AMLf5MYHo
CwAgBAbifhmv/FUfLK82qPKfnTHXbsqWtzbYH526rSIU8WEHYGLdXBIP9GXDqHCl
7zAkzLS8XvYcno1728QiB8a8f/GUokxKeAiBOdrCgkH7xT7TA3JxYHUk9b6t/ftj
ZS84uXFcF7Osq2wNqPZXax4YRpHXYQEWIWBFE3nvbs1PBaYyTc1KvIuc3k7PFVFs
snsSCuuv3aNxYnD0UYhddYyqYSZUK9Z4lzoPCpjhE7/r18n6DE/Znuizva4V/2Wx
ZSk2zcZ9sskvtyElMyzNh3eC5hH/7T9rikbvXMhwRajnwk2VE6/Tj1GQKEYKnWjl
wCXwFpVXRpD/S/dHdiD435g2dOGNeWOOb99LGi3a/qoORmtQE+p3knSBG7SvMAxB
5150WltF97P/xhvf5r/fat4CVjjggHdCA8HbiA7D4+JQ00VR/rtRGEyz27G3eXeu
jU68jfmU2GNqdBLGn9anKkgE/96Cw5wCUhvpAeqEwDlu+Q/KH1nGpsZIigCBnrAU
iyXjbIX9UTMVmtH2q+3xyngYpwPgqMinJOuhhgqaEhC6vZLUVrmVT+bPkhD3znLt
/+4kSK00MsXF+mlaAIuqnmU8De+rmrR/y5Rrnw1fGkreFtjwbOVy7hin233DkHfn
IigU+1x99zu82rgkhXBHpbGku4iNxsjTkeqp/hAKuT0Eq52WjJEPYFXzJ2BSoEu2
FitK0E/z+A4cwZEykHMvdeDpUqHEHS6TsuN+XSgCtX7fY/x6a/ZCalxFH6iyCzTY
pP3XrzhedQDImzR5OLRibXhok4zwToRhMhKEj3T3qeAyMKXOjf/BA83jY2zQImBp
L/fRGtsB+pQ5H0LVIEBlblLW7TkNlMDlW5RGg6hoUe8tk5r31//1llHEHmv1vYtb
VNl32iNxvLKjq2fwO0LyZPLC9cdkFfZMeJ4ptn0weTaPcQJ+iTNGySLiywM8mtjj
awAXh2OxVAmu4+86tp9qwt7SOcQvMSUjGawKW53xagxXgj8uSlBc1SjoWuBNdirJ
lOQgRo+dnxt8ghUQ/48H6rCR+UtB34Fb1/wFvDPwp3NcnNNYKd/QeAD1+VDt5R8P
7LXFQCfIietJ2Yacz/zmylqlrGgd3pzFGCBFhbcJGcv9swAYI5D+q4eNqD/MYu1L
vyeKltErEWE55Ga+VZGHKtVlh6lNNerRKF7Jz6xoUuh3vPmdV5PK0ZzUuJxsWnkS
06WCd+OzS9eSD96zxbnXyZjizJwfZiGDtoAHrLCP39Ak/BZ86poq00UKY9Be4WBO
h/PUkzt0hFOay/aki8WKrfR4OkraSHuEIGv6Y5tjDnI8gEZOKeHbk6BNFMsiV9Zr
tSSTwgPXhINl2T8YEGWfUXFBQgez0045OcSE34p+N9a/EOlPNOtek5ZBFwTXyRXS
W7CfMI9x/5YqEqywRIZZS+JFvIkDcKBlmazBaiUvFbcqeL6gozJGJ+RcrpgOhP7+
VDKDug8UFbPJfphwplKTSAMvzxjgkhGXMiyTPFhJJuRm2Lhmy4e9k7vz5qDMIglE
exss/ItCmGGu3tBhGDo6p7U0GB64H3ahnankEs7ceQVdjdJAVZRebAk5bKCroPM3
nSneHCnPnxQLS8HUHpeuIelzQC4suYseBPILe6KdqD1MSvODuNkryEQ1oxac8c9K
XZSO4stFqBL/QbscF/7Qw1Zsi65xOMKBYDese5d6ljz64vcu0eGQdNIZsTsNkMUQ
jtN7jpS4E63oBW0UMIYQB+IwNjUiVODxU1V3AMaeTtYdLbt6hvOVXglt1kvmzL5z
ktETC/bWcI+sEpJ4bYc9AwtJLzAQRsTmhRTUu3/6IY9zJN7QLqSArJYA7I30YKHR
LlCfrpgnnA3YnYsCXemyXZ6iCBVf4c268Ti+2beWerilqV5A5BRhqLj3+eCos3gW
xddG1VKjkh7N/a7gnuLihr+iMB3LpqP2rFRsTK7QRE2FtNvYgRPKF9WfGBAAlg00
g8iMFsJD58J8m9uwHy05vj7m0hPlg9RfOkhlKI0NQhlNz6Jo1kYf5+FPXGTqG6JY
isN6nS6p4gvL2fmZ+eCn08ExXVYiZxlfw3A8znD6tEiuN0s9uSxB4+n6wtbmzvnk
JTVpT74Ff7Gudg6pi4Zb11Phf52m9FW3oQzybOhVknpHBnCAQKT8fv7VJaXEn2qj
dpGxXchrZ7IeFZZ5Cr6CUFN/iwOXR7jSwv2DurCC94p9aaHP0ILj09+4AAtjmWAP
3XOU6bbOOxOkOo6v9FBQRo5fmQ7g7J785AMY2GPh0a6iAn0cYzACUV186ckhlFcX
Da39s6Eeap/OtwpD2dsttw3+Ty5lcrpFEm0SxX0OVrvebx9orBR2a7zOPcRFmzaQ
jbWoMtFw5GQs+da/SCfTzedkVTDK6LbzMtTCjMGIezhl2mQlm64pT0nFJP1+ZdQq
M2013T+MKj69j6muHTrXd83lm3jGFjv04PFOk7G7K0pWFvWymPqvghP3mrQCy64E
sKPsw4Qm2L/VsH24ihZ4eCrgdhXFeJwgpO9L+HRz/NXcAQ03kC/x2ySY5Dfr15s5
EDDWNLoLwqA4BMRIGVoQUrIyvStILM5kJX61wxbA5cS8cnoVpGBrHfqj5umbDLoc
zEh3YT4JSF2YHZVrT8UJFeWPJw3zZQXBbndutPOuuwPqnwBtZujRoVcSBy9gx3Fz
BT1ou2KOUjq7Sso/AMXurqPnNQ2cQzRqhdg59MVvlgIvWNr+/KZsZpiSM9DAWU4g
33AXkFOZkHGy4389JoZIGVEZLhFsc0h/v9WlyTUMAuby35hs07Z2VcAeYc9NvPR1
q4az53Xjgmhw2iv2l4QqW1jUoQFeDODMcZv5d4kKMOyQqboorHc1VpEdkQne4DYB
spmpa6yQZWoKgLYLRwDsmvRKn3tfwPsHjJLaoS9/mC1L87buvs4vkQsk3fZS1jkm
KNW+WQqp9o37HnQJxO6Gauaktr3LOrC0DRiG+pj692E26DYJnVXA9oZQQtKMbJw9
80/Gg+QZK8lOd4wu/uEwVGbl05dIApa1uxejoQt038z0eIT7jHh9A4Oyc5KpMTgH
jC6eoE9vR6ToJJcx+wuR+s6hIAUGnO1mHIqVbc7/+VpbbqDpLw4eqHKUkcu/y7px
wadgYN377bPQRLgqhraio+z8o4Tjxd/rDitbgy3VMWUfimf1+cHajLE161S7P64M
4lFKHaU+HC6hl2fXqt5WtVsQSUYqbfKgZUpToDX8b2soVJjDjE0ngQLIZUk8hP6q
xAJlrS3q3+bT+fwVV53fZZ5/Jzmoc2dhU2OHDNfkYFtabe9yB9ampAoAdnmBbTM9
LPs7R7feEzXZjGha8CPwTuSA0v602Y5UCDLyGZeOPgH6MV8gl7TLgOnnBI7IcZue
I/m4+Rkflr+l223ViIz/4HxXefY83vqYLBPRMcyqYLrqaWPuP3Zy1bjTvgLPdTU3
fgjSr/Pd0tiAsWw59klwb9/NBElrsoEnHBqcaCHO1VKt4BWMb5trjgaqRPlF+B/Q
tXLvOl4rlyG9+4t79gyzh8Yo+VU4wf1D22Vk39Uwv8lIyU4I8ulpZXlQhtYBLFSZ
qfgx+G2lrVP5TM4oOoqYVbFGDfjk+f3O25zwEjI/7r8ywE4SkXGuqb/S2Z7REInS
1qfAZPGDPayn4BckNMhcJH+4a8Qhxb8TmqFP7DAygxUUEtGYFOK4X3ZAc5OQqu4Y
+QYqNf//pm0COca21HtpSXqcmhjJqa+XRv4m9j7rWrY6Xs8l7x2tTE90wH0+q9mb
bxpqMGZHdseg/JLKX6JQ+kCkJh+hoTRzDPGXBo/YN748/Y55RmYTZ9n0d8RQJukO
FlOb7vt0COd67P8MO5nfHWI0PMNdYK9N37c7QZsZx3X6CljfqqZWpqk6uu1QA6xv
uLRVEGR17BDPYO9iu/VvNl+blhOTTbOiMtiEgvBBLJMoDUF3gpHDvjd0v30Zbi4a
AAwX9LLdvIV1oDhDVCNepOQphtW1Aj/FhNeUwrHuRHUq22tt4hw0deQLpic8Zev6
73s/zC5kaR+4/q7SGC9WmO4du2w+nrGJcROD5NjFceAWDXJUrAXBeJiGjw0jml1d
7v0psvwByo/qirJPbOek9Fxf4zmaonLcohpl9G9juR32fyZXjtvw83w3KAxk4IIa
N77lEOCULRU1XcOXLTEtAVAFJf4BrTvaVDjd+yE74yRo/EM+KS5Lmfwv46DmZF3m
ArDFDrrZ7JWvWvPlVFtAPb3C9gpE5oJibKMUsb7xQh6Vi60DVD8rPksXzVZWKSRQ
vKbLqo5phlcMMMZz8AVo8BBGJqDrYjprP7BZ/QC+bf/kzYY0QReJ9a27UQAedARp
KEzaC83MQk8JPzWwa6Vas31sjDBb7AUujVox8K5kSUwGkeUQBwjp40hqCbdUVtoh
FSJOWQktitjdN1bilHk/47POj4KrIZ2FyJjOpg7kXAgE5TACMOWakFdgachSfaT4
gRAXUG2nP86oiZRDrGw7N8MHdQsIPHS64Z75qnOdbJeDqgr/A6sgN/WzoTI8ZWC+
vGdXCbhrIFpquHlSfHYhCEdXfRZnz5gim4xKRMdd/fBxFQsHaYjCPJWyEs2Cb1j4
OijejPV9YcpMNlj+LIbefGh6XjVyxkL+eY11Qoj4FaCxez413qkTU9kx7tJ7mZ10
Pt13aixf9FecTGE5t7EDt9L4J8fyUxnKoVWbHRZekHvb7uCBU5AUBsFo6E9+S9Id
UHCXwKZUk9iSiati2+arug4pPTOUBpDCQ25aN85zX0BOVH/vUODKY5VewADrKkWx
NpvmvitxysPTaEzMK5/wY7XcOCsrgPHRsssR8Byn32kLegXEjOa8Bg8V1RJKp1ft
AFTtOQa3AedyTeiNi8rBKrwRdwyKB/XPsmo/USttlO08PIUwCjaWaittlpA0JA8k
OKsCYxQT8Q6MTFT72WDzumLSxdJ1ugAPEemktLpOV/nXnKFhQyLBkRihUUgrol6I
1dbCryal0sM3uYgheqOTvnjEEwZBEUBOBhyGVqnTFOhY7kb8tWPHTo4p9VIjtKij
5IbE8Gl2T1UGOCw6du37xC+J/Hw4LrqxV1+fBdIyNO/jWm4BUU7kcRI0E6zHMsDZ
IA7K8d0TyP+wAo+9BpRPAq70aprtNSay00IWy4LvZQujnkoCJWZvTmTw2qXo8L+0
mlMtLkC8UlUuQ0y+y9vy4scJMWiXvWQXd9xoEopZUASMth8Ni8qtC+OfOyTudjGs
CQqTm8BjrQYGW/j49yeiyfafOpIsLBsbiQkO3cDHo3MSsDLeV4HZZSJ3kjFyjMkP
O+ddFl4pqPfw8FL/Wfw+O1ELYQWdDLL1zDIo/2h79OQII6ijVQF3FH+Wx6f+8ZFB
biDk74ypYGhSOaMXPaO5WLAt8LNpztBhN4IpOCimauPgIFkwRW3pYsesLI6GHbGe
l3+VmSfBuZsT2mEPlTumHLfKY4kpgUCZTDs/Fp7L8Jknmn5MZj737gZTkbb+pI6L
St0HQrp93b0FBadTq5NZGcyv19IXWtvtgW9gTK6BonKnjdGPI6qEAQmHaAVd5ScV
BvRIlSgYa+xpvEl9h8YmCftQjs6C3Ai8bawct+EOPd7db0ayGksyxto18K8QI6ty
yn3FbiY05kvN+y2c0xN1ZZNlOOYeir7cGfxvDpQl1TNym7r/Riye+FUWqLSYZQi3
fLy3qj2LrrqID72HxnLHDt+mpswAMPQYow5lqrEFllb801ilnD0Zrott6/kPtFW4
8fFOP4iBGT11Bl1v/y20yl9RaqEgIw+aIxx4tldG5rPBiUtU5ADkYsO/wkvqia3X
SEOGI/ppeJEgy081yX1p2uPugL785b+FnQiXQws/6hGmxIIBWsrfM2YrtTVmoFao
vBev1BzVq6WjYMuQynvXTnSD32a1LLkLWB6fDjX+L/jDToVz5b8Kdz8t6RYWKgzN
NAp4y/8Tmm4EKpOTodtWu1QOozXPVAkPo4M4rkrTILH3zG0EOyI54DhDOzjOURbn
iWj39OX1rugDoblF0jN5HeD0OgOENi890z3yHXMBcBWyBq/NL5xfmOxAzutQtL5y
K2oSlkjUUqwakjtXIlnUgh2ITuqIV6Bzc54yko1Au8LYTxwbqnbOFGEAe3nBQF5W
0VGi1pJ+5MHRfHlu/E0oKNY7ecVINlmjpJqSvZSnRSRljuSBL0TmYGoakvIpmiey
+oK1anwXqnOWYwlANohBVeLWFH45PrUHY7UXeXb+j7LkVAVusggGk5QvRIaZNAeL
gj8nldT9A16IyuS0BmYzD+4LieR7PptTMVMFPC/0EHqxpZ/qcru8BwYriRnElTKP
3/rZ3pReachXI2nhwWtumjpsOo/t9uDpLXY4nQI9BssLZ6ftV4ZHJ5zV0+gHA2ie
fm74y17C+yFlkGkrU9Nt39yRwXYYaLyB1i16+gMww4ROHV81ePmzKCAHCaIGZ8uX
8BhNTudg3MBxzzKNU001O6ZiZGiJ1tgAhi2mBejLCyzSmeBeJSS8/K1qa8NR5wdt
Z6TCiJAr5Qad2P/QHW7NETUddUMhCOV2rAuBxuCMLWWyLEOQXNDVyf3ahFq54Agi
ak6IPgR3rP7JoYu4sETgyBvAQ/E15EgILPgQOh0I8d/b60PtZT6MOvc+gVoLREkV
DoaiqGX/fS8sgBAlvS7k6dEQlsJoWpltMyE9baBZPq5lcS1EGsRT9bwY9lILueDN
2dZHAJbt+F54z8ke8LwamTHOnx4oF3mvwwvvpYw9aQVeBLcObMhj6prEC0dpy2Qq
UFGBrXVVwbgnsLsYFnMIL421mc27sDIvzT/Vt5nZiuhYLADYnW/Tp6pa7vhdT0m2
BBIPrfelZvDdTw/HgmKKSD4unBGLpo0+4TUDFRcsVpQ6poUJlTQ1J9XMy3qQU37N
TyYhYWHdJBMmxqM8WP7NulNDYRGlhzdoICrWY0B1/UlWUI8K7wBsZ3mAr2ayU1II
2yoRXWfcw4mF3enGo9S5Dq4nfJFcz4U3rxDcdWLomT8n0s/hXtP3u0/UZMNvvoqs
vKnAFIbXhumFUopMm+aK80LIUpJtLwl8qVnsvOWE4nHpR4b0zRO2nVw4DbufrvIF
akugz/s3r2ircvSSw7t+kAMgDwGjCn/eXM7XuWuIJe97hUv5IUtjSkwpiyYCqXeG
52bsQbjHQxOxKMHDYXIhwA3b4b0BL8uS0x34qiw8jG6LbIkaEd0OHTrqy8qjaRkm
klczdv91yE/5dA7QeV7uWis+56QRuLlLdSyAHSb6RtAsqpjq3MT1m0HptukaATXl
m6wu6+WBj6A+8zJ468SUKtPfaUQh80oYV3E+t8/L+133cyxpdo0U+3sdaNmcJqOA
o29fURnLjxAT1y/jpPZFZP6ZZTZby325nmj5hutLfUab0FBURbXUORsTlRFVyMbr
vHAU9b2O8tdrOO0/73IO6NxFxsJf3+9lCWevQfaYcfVUc2dTjpcUMc1PItjXPc88
y+1eSOxTiwlK8UsUnQRR+CSZfkAmg//5xQodLc2EmRUiPKPGB8rJkGJ/dGddf2la
P9LRh4tUQ3YxkvxKRTSJnxfknYN0EWgU07JGr3D6hzfLt+InCjDKT8aDs0LlJ27X
9Qi2jRhZImhrLh69/paDFIPHK3Fx85aof9WvE9dSiXTWb+oCp4+6jv9Svu/yhvFA
kD3kkiN4JJsXcC12yTAc8WL1NzpPeV0rsKIs2IjVLr7SoprcnsFIUVW528hQUaL+
xXuGGXU8FdCZGz6elj9C65AtK2nt3GXdMcYBR9OW0jDcwXvccTOr7OBTMnD3tLfK
yq7NQ/vc/QEGlokjnl9HyI0D0xjQGVdLIjtwgWjq8rbukZdh8JkENAKBwkMHBObW
+uzTaoEbXwjbqsYmlgeVuleju4ZwXogE2EjCRRREjTnLtypmv5T9WJdQ8rNXxjzz
gFIXiUUnQKSS+UXI3v79G+RitbFkUIAaeexfHXgqxUsY6JZwKRtSIGu1/3e5V5gR
TAubfTSzvUTrwIO03oaaE7eanjehQQxXuiQvU4qX22iOPyGexcUQxMP78czHBL0r
LIpzrY+lyh2lrAK0sDGytACt9T0Rhr5sjMDY97hPqDS1oAzxAODkgycDuJ3mdbYg
jqPBsGsKymT0LAx8i1dHXj2AWa64JlrRO3zazLqJybNpIKh5aHTFKM5yzjoCMGmA
WUPGWjQFxnlxr8aZsaO8cHdbT3n3iFtRWvtFR/tMgMfse9fsRYESInFUsT6ezVJL
YBQstOXxol626KguS+TlBXJzjKgP5MJNpS/34XdcAtU2Y6PRdPZDW+/FBKhRcoLQ
u+zolejvOmv0LIFOhPQoOC6wY2/tZpp6UrcKoFMvdZIwLzRQ5YqKHJUCwla1t+c1
D+h9S3bXpI6gqk5tuWVock5JIsu9JDKO0x7h5OZ9cq/XbX0PCepFwlTG41tcPvRX
+DOYfwxfX1lTa6/g+Z4SW2qmDh3Bq91MoPFyQetzKDDkSh68wd/2AZxYwdyvkGV/
Hm9hYMJd/O0uGFUrQuFyESMQx+xEYaZwjvxwBrBf+VqQyY4igxKuOMFuR/uea0gs
XSMMleAgNW6bJQGBFYOGtWivAEA8eSKkEtruUlg6Y9yh4irT20D70NHRzXHppIqB
s9YS4gLIG7CYI+Z6Db6cX26EYHlRfHgl6AYC00TJpIdzXyDVLkhzPZZoX3t9POoe
edNSEiVUVl2qVj2i4b76VfKGVLz2UTJM7XsFd3hnkI9ZF0gnakeTvNn/MdVXZFTJ
cv7wHYF5wzvjtUZRknz4M2NxmPCF2faSh6AFWECo0tHku+z/JxrZik4q7pJcAuyQ
ogAz+xlPHOt0rv4UZ9GI+szxVasSUpEwdyRHylPJPNp5AqEwaFrUxFduCMe68X1y
dSsfuT8jxOCb6rl+8WG91MQBrTaHmvUH1YJN/9NRH+gXnqI4V4jx6R2bFiIrMwRv
dRCpusYwTceNCXuInJdM3OWzJtraicaIZ2W78eVR10ZqpkzWjkWmHGmZMAHGx83K
QgCzWxBW/pjKN3UtokrZDvlxGR7PGQWmj/BNZ9yS1i8YUTecYD3v1QANP3ahIfp7
3/HnbbfSvFduT5bmjkHb1yVCpVUJm7PzKraqeRZhdJQfbcOYV31L0Z8CynsVWMX0
i2hfYVdoQHNQEv3eDFGH7C+K7T5kFKeTTlqaXu+oa0z5SoFCKJDEMl8Ppt3RNPlm
ei/B+mPxsyKOUz3v9+CoDDJ9aKkNSRkemEZf09aDAaRoQrrLRMHIaaIN0mp9GwM6
t75To1NyB0D5ewQWpdA82sRXETUMdTCSaLszOYzJwDYMeuit1Id9uJYilbBTyxRD
utRFINRXagDqfREshJozXNCjvx8RxHUwlukFd3XrO58bGAgYL3Yo+qc6I6Q6Hxdn
GRSLm/brH6h725P/jGF4oEVo6V6xoQcMs5sKVNETZ1FL8TnDfZt2E91cDMVGoPtJ
WVPwKkkLyKobgjbrt7cmbylW7QpqGhT1mkAA4lT2FsHBEYP99q86GVev6G3wbr6+
ltUzLao+bV7sHgu0TXuPEq9lR7kHMr4SHl0f1yxorRulwzaEEPlUVi6soSE+D7ym
3MNds7hBhUOoRMbQevH06ciO0kQotR+ZWNuX3Rc1AUdMU8CHpI72DVzE1vdmAPHp
N6eX3/du38f/uHNRvGnmlvpNij/ygpVsrzWKElZcpCS5dR46Kyx6D2dPkwZwpz+O
jTnq8QFODsvePcDwdmeuOBCa90671UIztN1Y2U/4xX1COQSeIC9Rj3EB9mdypZ75
r15UXJVnmFh3s0cN0zrSh4T8JCN3p+rrjb/f4xoOO+Trnk8NiGvyu185qx7DEPAP
f3c3Cm/AJIMruWG5HBWcHZZCgu1U2PhymqAXyi5NPOZK5BZrD0eB6kY3fjkcNIL3
MNba86BaYi4CJD+Uy2n9mqYUZJWOqGbLapoyUJ89XOR552DHYDeXOjQGd5K7Wtwm
8vRZph0/C0L+8WLF9bs8KqPeLRZnw0NGR1w1woIH3VOzfaq8Dqj0Y/lCgcdhmRTI
cm1LOMIVNDpr7LDQhp2ediDV/qKylMT6L/0lbcXcXmnZ15ANsp6Fj8Ro3gAxjewu
fjVN0VdX8e9jq8cdy8F9dIVGuEhb05uki+Nslin6ww+Y5mbJjtAXs5RQ1AO2mZ5Q
tt76qmT9uAMHs3HUcDQLRP4ySTJDyEjrUlaauCwTTJ4FZK1LBAJpsHXR5x9/szTF
2s/WV91i0VoIRdnSBTYU1TihrmdmZkMerUn4Cyku+ThU0iuuMrDQRRftCfEfwTFh
VWHAQGfaA0HlUbyaMF+xPLeoSNHs82cpz4v9N/M4bJQkMAE7nPlQ4qW5E9Ijn3oS
o/+mtRnnG0+HsbsbU+VzUvok5is+NNwaMolv4gA5KYgMOg+zyZCzwXAm3XGzx12N
r5HvyQIlLROw6NyYfoJ+vbomiccBKrf0GWiXIpbwHovVKgFU+9Oi/QgqHoAxlYcc
xtobZvfAWk+R1cm2AdqyrTa7NyKYqAvyJZsQ5mx6bQjvwvoouM6guJn5Z/BSIgnS
5CqzrYXEqUyQM9NV0hOy1E4+kzUKpsq28MHEICM7Q5xiQ1v3VfwN37WxMOUgX8p6
YqX24FLhammp3iEkm5xaCoo7UDEaSk5W19hcbp9JX7NMB9FG/bejhIFnbranYjV7
0cBWIIJHtAbRp2C9P8/V4Bb1kjNgEwIp+i8gXnQfS0U53z3s3gor/FOcaBzoy9lK
Nso+NnVWjBM2JG3zTzvvStT998HKjrkBDbMF0UHlw1EwVNUbdCPysdxm5PkFOCvj
7+bjkCCoSwoya4wtqOFXgBnG3Cu+FwWpdEwFSVA303dwdPd1v5gvOOgWFlGYI+ij
M2Q4AiXMdLZzT5WFvQpUYrkPCLtrNjH1NxHsP5v55rbqDlfv1jOk8JHfCXiQugaN
sXaPYXmQTka1NG3gE1rfTEZ9O2kFZ/lCq1p5gxoch1+Oft+UqyYtWs0M2P09CduY
1w9vdQIeWzv53NMcrEHSuSv292d17dKtHFkUhGD3UmtVqHzhBDzSs/73MyaDUc2L
FKyxoTfDsrmJxn3YhvpvVj7kAlGGsP1nnf/gxL92JE7Yg9uP3Eo7toeFTwMsRDmb
fJOAWDpZdZwq85QwCZscXpWMWzYL9GkAqVxGpjUXpB66rit0W5WcUaYXjNXnvz8v
2DriJXDVSdvBbSr3qoZXy8T4bFlxjyPDeqJC+1F03B/etOQdCLxQxVm0stXLjuin
nuQqF1wyUItCdr9cVo9XYyqZMdjVntEB6BVtJ9yJ5lhhH972UL2RO8hvtVv2JdOw
UZwPdm5U807joDzQDcDr7w+bc5tBZ9IGwm1f997otIRRZlEAZMVsdY7ibQftxkU+
2E+vwmUeBmQ/JJuozGdJ3zaXunaeggLQKNX9xNiu2R+bpbDSgGUtGP+k4ujjcNwS
OxPzixm5vtM7qisJHpi9kWwzZO079p9ZtbYERcjquoR9f3oSZtqwZ0CEFEcKeQA8
FeyshBCrMbnMdFfow6APjo2ybDevPkEaGeBFpZ2IBRUbEmkuavd7mpuQSn5R9Tf3
j/ncRV4/R6Cc4C105gKAuPW9/PJdPyl5c+vaKlaLqFFMDaJMMei4Mdx6vRI61Eme
wYP4KvL0vs+rMNFwW4OHvuomKchuU6ab74o4sXPVT6uQRS2ITk8nxrNKVAUZ37Ei
Sn6x30tYJnTnJigpRVcG8WJ+bGoP16M2jmFvTPaLdzvf+WGlc1XKoyhA64UEIkNu
3UuCRtwnkRtDICyAHNxawBSPMtDrObsuhOUUYpPnZL9/9fqvWfES/NelhLFQFHlk
5oW0nMs7hyS4jyr+gDcaSejpguNRU0qvFqPCCFU0tQbRxC5vY+u892EtKA1212Tm
gYA81WS0X2Qpi+uL5+exccNoUvw89P/I0d4d2PqIqh+joFYa6pGQSZAXg/s/ZrLN
+54i5BxnZpaTTiuUP1Pf6eXTVeDJ5KmLQE00RQ8JutWxLEGJkJHg15TB8FDeqBEI
HOQqU+LABoNLkXS+PNMbtLo89K6PLCXhDuQbXjRi8ylXLzgDKB6Ha0qTnv4ZGIsU
qTwIa73qahal9r3wsJazIfwIjCiB9wBzEicvy3ualUGoZiPGIgQlgKdq2Oh3LQw0
aeat9i3/kE96Y85qchOawOXr6wm8/Qrhxs+e9P2D5xGNjTBUNK7K7tv+jS4NxVoh
24/hrAMupAyqpusYDZtBQuJHBJmGKyPOqse8RHF/X70HH5ot7+jCN4z7jHeQ5R4a
3GIQwNC2hxW3jxwqSXgQb6K/Bi8zZl9CA0v5xt2szdeQIWUVD8VvYUYutR0K7nDI
hHyKBfF8llyNSsBfZHPKsN2I4x59kYX0NkvL1iVB9FILmUKeAh1ThUXHn72B6sYB
4qAFpIiX1EPNIGib9TeXBN7ZrNQmEDZyCW02INWkHf9HrsgoJYYL5m0YlvGev4bj
mtFkbXf8UtK+oArCv3yZPPtSae7qgoOKkdgYodXOgmJhx4huhFotOVduHyZ05w2H
F3fIvXQy+1wzd5ds+Apm7330x5mdXZSZJOoSojA+FKD49g85B28oLoUCSTJKRIWu
JfgeVltjw2oTtLjlwm8juzyeT07rm7eXhvv0GD6TRcbbDgYjDJkPSYPsLWlqIFm/
JVRfMJhH/S1Oe7wL18ctelEPs5o4S8i10CdW+lQ6wOAjcupYDICUzUJdXQeT4KOZ
tT4Tid9Potv5+Lzu9Zo+iKXrLQkdxPnCz/1wECTZKV7B6ZfUhzQcPLXK0yvHxmBT
zxMKEysOYGjTUfjO/Q0jGUyTerkF5qxQfefydKLbubmVr/1WfdETu64xgqKlj5LT
YkfMVwpec8FIGjVvKu1tHhiVHy+cKnSh6rA36foXQPIg1oMH74vUF1Q78Itv5Chs
Ki5fdjORZReBCn5eCG4/WeRCZYYGByBrkZlAxEseBdaYRv/STFY9T9gWkfZNYihR
BHtW0RX4cGIREKkoXBSzVwB2wPGw8U0ee3tXiW8gjGla/ghwY04Mw6IjLmEnfKgx
HhEw935urkHWy93Ft1acMQOOP9HIUWwEiZKfej4CgYWZcskc11DoJXiMiAIv0Tk1
QDWfj6S/2c5rYrf+4bxcXde0nEZSFAx0OLb2F5QqH66nquDZpqICE6vibBoGtMNV
prYkXVZMp1qr0CnlAVOARw3fESJQvquRnkHx+Kd35MLnk13xTiDB/8lsoCJSWYUj
y7Rdac3RaPzWbrOVynWWUKnrxVUKZcE41/gQ0QRW7nlqTIiuFC7wWUIBeYJpeOb5
h5MxaXT4HdBQJSbke4BC9Xb0HutWl7IeN4y4S74wFdu+m/TfsH8DPEKGbuYBzDEB
V8gsGE6QzvpRktcwQ5FtpkAgz6rN808b9Sile5KUz32G+cCibpOpd78iAAm4GQ7A
yszXYIUsVm2iZardxLG5e7ablPJ2tgaUNqdlUvUjOdYn/dzJTPtr2SpWwaGleBFZ
KQ9fINMv9vFT7drGPy4ANJFLZgZTRdDJOeejJMppBXMaILhTtGovsq1rwuv+tz0u
1SPynRjhX8odiC+Mi50vXq85zUAl96+8ZICffB33K5Ortv9itkBQXBZuYM3WpsPy
2LUrsiHm2+Pl+sjB1e/VjfWPb0rZKWhmu4mS7/g2BSCVI411+gtq31MQCh1k0zWN
ObjYo1FY6GpX+O/YdM8t113aaWMjDNzB4kzMDZOuuc8942sN+B4nrQnfkYa1X7Q5
LwShLSqz2wi5RFdL+yqtH4u+Qf8xfjG6SBMRMJoCtZq8k3qmbF8po63AkUqX2kf1
wLaTxkpmWdI/o82HAn4O9QyP/eq+udJVMt1+A0wQWNdmNVqy/XPu7bfWFooIbxs2
+2OeOrUxqEwHM+ciD5fNvrNauquyfdNrRnHbhkjyWZUmuVIAdPdAFKgT+9eZsEgf
yvfBqfS4C8+ESwe9edbD0vELXKTnolv6lyUAUMYyI7YU3SFApSt95yV7GwHkQpL7
I+wMBeAdltKb+wBXh+P4qxZiZ8LBi8jO5rz5vhE4WVdDSOR1dc3I8pfo7jARGLvv
QSPYwXNktDzcIC8uNPOUhoIAtmsl0eNKZV458RxDrmFySM8tTs6kCE8I2OQ364dQ
LwJtXYHojlqTjFoLDJAcn3o0DnEQq2Bi226jOekS7GHk2viXIk6DWtyu/y9It1fl
Qe1Xh2OF8DBcXGj1FpD+5d9sQetBiZ6OYC5t5Cr47+h1japzLmQqEpiupb5ofWxw
5rDdwFjv+X8sSuuAYSKXcJ4GfSfLAi5tt88KKShGWOO1jHUMfoAC4DQu5cL5Y5kc
EuBEnIN2MDrwu/xi4IvnAsoacKRjOfXNAkAwAm1MAQiHCS0eJ1ycQTF0gh3TTiRK
NqG2O1hfl/ZXoegAswTCOt805lD24M3P+B+TTQHb+/t7XVilyBaXmOX+Yx1rtBNY
OowM2o0oIdmW5Rnld2mf31jH+YhbsyUo4szP0Gi0x266DYs+aSNhmgsqMe16x3Kk
ngTJ0lGk/rRhNKbakUquWbzsdt0gmH8eJ8x5Oli2M2mgkqzaJ0Rql/PhczojctYW
2nzpT0AyG+jEe9yo7fZQaahobjfnelqHamWV+UtWI/+nplf61JFqs6FlVNLLexZQ
mty8FaqVwm9Nu4J++P4104AAaTppAoOSOe4McVjqGctTiK/x0ScnhZScZZzc/kTh
qpj6q40P4SOHTZQusX+inyEAiTK3Kfma/tE2aQ1QHHGFf0vRNHMvoBdnzadmvtvo
GGnV/5kiKdBnA3cYkx2dypy/H3R8BFo7C03YpRpaGpcSZ6n6DwbLaniHS1tRyJTx
QsCGaAooGEypY4oyi8ABNRtA/PJujETAoTN+J19/27PrwL/0ukXn4+zAYXs3tQos
LiJX57iAaqIZevN5co/i5ddxrcVgprxkuiMdLwkFUvHs3HDI4HfE+uxrkLwvVRcc
Bcqw07l/9dE8fpBqKKbpMjs23AjG6zS2S7NmiNUWIiftO5B8SPgBZEWKqbheoX0f
RHBLG3ICJNYZ7E/PVISmyUWbxsi6V4TgZIQVQ0eUHMn0Of4nnjGu4afU8/PMPcIw
R3hlVRiqKGtye7ko3XRKsukflNhZmrI7a6M7cveKrNJabbbv5Hwp4OZ23lU+DicH
rn7zQhVsArSIXqUGopcJaP6PY8bFN7v6rPJ3eJRox0biS24cc6r/q+jmwBRWEcNz
b1lcUeA+AP98vcBalS1WE8nUt+NRQLbbT60odoBRWBiJEebGU1efJggGxgd2gunq
s1PAw3vTXiO9TwBQ9s9jJrJgiLxVvMg42YdH/pgvhI6GsdRNQu1Z5G0y9EeurUbJ
Q0DXue/XSIqm/jOgjna5CD42o/0hKU34YHMxHy0ZuROYCnwiVrJd4dlyL4nZKar6
FPTMfMhV3A9epz7LwtB+v14iRIdqSYjiEoiQWQpSYJU9bKxXc7QDLh3E8myaR8Ao
IsqfOfNZSukOo4TUuY1ldPfhHuQzAc6kaGk0fgj+DMaF0wtgxDlL6Pn5NwCFkO4z
T/MqnIuPqoKWPoutYGSp14l8xf/XnCeE818UWaaVKD7e1n5sjksKZ1kN/mwqJrxF
/S5galeQFgQ0c7sl5NmxRM+RvwoA0K/rNoPTFwfma5lRe/+cu+6q3TvqaN49Z+v0
PVlDVrASKoHM9AuSiL5pNpndC2Gquc0/uKG7Ma9d1nc2JBL5igbE+pbTeNJhb3T1
HbzJKiBFBVys6GdcPaNsoaG6Gp9NrzVoV4IXM8l9Mh0thtVNbX6ytqybHKrsJ0tC
S04G64v7i7dEGD1MdArXH3DMEyCbknFOL2Fr46lcffnKRDdIwlvEewqnqN92X+70
EDjqjrZYernB6pd3nJnPhBKnW2tzkhkJqD5dnU95SybkQ5dOsuVhFm9sz0ftGSOS
xpGbRoHTne8bpzC2c0TCadrj6rvc4a43x9IPNFx8ZXwZJETw+7BzaLDHwt6Gr1+G
MWM2tEchii1ccxRTvykLR6yxpbAxBhoE3w9Uvb1FL/QF4Obz8LzlaxypY1DWE3F4
irrFsEH906i5TGmzXf09ljrB3KyGJW8IuenKPb2SYpVmwYMehIx+y59yF86MMPjV
LlfrjiqWm5jJDs3KNmSRGSJ98Hhsv0rEXQC9hJBKybQ/XFzwrMV/XHPkEv85bWc7
1cXwL+JTdtOET9Luw4WYw9E9p9VVkk4hvVwsvyuU23MFpzLQuhVIsf7KDxRLBlaN
KDepb+8GiM3vLU7hLUNc7KoHVI0wR//zd4NLfudzH0TdTBzfI98bqgUyDwes68Yl
T8w3ctJx3jQFwceZD2gzdvulcN6o2/tbBsyiISmPtU/CGvzJ2lMRMcPk8FIyFPht
GgR1hmBGGg/leaW+NuuycVaMrl1pElp64MKXQegdmQcDNl84o1TumH+w+LwO5JuD
lFiDXU5cVlF8OM+fZNeyP6AbIzTIGvKwrlAzStoWzF05wtHRJf8DAudW6ah4KGRL
pO0k6JC5wsF0ykLAWacBg+Q4DPmgWQyJ7byHNpput5LnfVup5cyaoNX1in3Imlb8
SeNxRm9gkjeeBl0Lsofv8jMR46SGNxJvpbV1o77cxr0R9CeyY2Ph861vJ1Fp3Mov
WduBxn0UPZQEaDYU88jFf/Q6lNPD15UPmt0jQbFzgkvGHL8RW9Kn4dGM9OpySwTi
ldUwEmOzSTtFCSfN2qZ44WZypJXI0R96qYtWtBT7OHjI/nxM6F/osjZJnA5cRPla
WZx6EluofgjvNRzBoiBNHsPx+mFDe0n2yCOkvEYquI1tzL2QdNtlpvQ4jTLc21sq
rCwUpq0yfIByLMnUe4cR8/O2iM2nwRHzquobE+m9z73IymBba2WuzS/eGxZVjQBa
kCXNC1QezQDKWXtyJd8VLSUCvXNa7aHl5oKBC1IhkwX3b9scbJ3Y/l0qwc47TSv3
Yu+YIuNUqU61QN2ALpvSu9nIyz267s+7hT5u+or3aWqEtCMIHzNzV8DGi8m+9we4
T4dzzpmoljJ1P3cIGcP40HwD1R3/3SfwCn0Vmzjf0nFQnb8E5pojTXX2o2QymSCy
e0mG7z7pSakURVJRXLCVUF6ACqPopuy9NWDwOqsn/gDHnXMmZ3w3H0PIGjgDI1Ku
o3Ex2iHPG1iX8MeoucHi0pRsqZq17/MTbWmcu8qaojbg5YTOZMYRJDow1A2kxEjN
E2U+5m84nnZdpxgqsVeP10YBZ7PCrlVAcGSo0+I0APp2WdjT6X+m3gNtk+PCHa+4
e6gaWlxMyKHliPdXDSpz3BUjVRcIkq5ARRrf03pN0x25knm7w7UIQdI+/DS6vN+u
RtkNJw0JN9WIKkFtgw7nSc7S2oU0kstPY/xdZjbjj+MVgBmraH4SsSeS2pflj5ef
ERUPwrOqnt2gs9dw4cBwUD64KtoMx0NWMRrQdrZ13ihJ542wAe7NJ7uLuwqHMrA7
oulRQRO+gftPCZDCuQaK4QPbxC5uqTt5tUVFPOjbjdoLOTcpkCBJsVMMC932NdBh
xljWZWqqa+SmGP7gKx0/zgX6W/yJ5lxHBv3SakVPZRY3JaBoxrvLImK4n2cTv/Bu
k2yiuR6c/CsJR5DWE58gdJijWFjrKzS/+3AF5Aeah4nopcsecz8o2LudDvhvZjeO
yK5hx4eREk/IUDNjxqIjZXyrupXsrkHQNGFs8oEWh4rofBZW69nWQ+LGxgN7mNGA
CsMg3jHUkdG/nSp/m+/u7RYSlVe9IKoCg8ik/wNujJiPXizDRxjXEHzGta76MOMX
ph8EV54dTmQGacGAR5Ib/Sa4dVIoslNg4rhXMExLjP6QkP0AecoSmihOH16h46CI
BbQqUcMX4UhiSlMOGmaRNbv0enz4c4Yk0mpceFOsLm69g9Bd359/KNytfN2yuap0
nbhRI4ul/0TVrvhbNCYbdG5tkpLtjSfpzeOzLrBVF7q9xXiP9Tw5IfvVlBU1V09Q
PZbyCgzMjV3CgdGRDPT8b8+7SmQpljmaOTYh+2/x7kSoaoZfY04GFqIzJ0PQp00x
W5lMqIcTjAgUnzRa/Vt0ElE4GsbDneKx/QYsonqt6xgJYPfz+x1UJXZpPDw0xU94
0o/ZAWe5TpWxwAmYJ7+ALbIjEGmDnanBpA7SmadcZNqLzK6a8S941Gw3uUodLGsU
ZMGmAgq0ZR9DETdDrTd6wAAopXhv2SoUsz2ZVgxuHCy6IWBV+Upd4QJ+qrgKFhCE
I+xlU8N8rg0bUiFBv3K+xNcWEuYaB3ThFzWXwxLIXD2J+MHtpwm2g3cr7JMkeD5E
/ocqz7P9Cv1zX4+/WaZVLoYY/uIEndKUysM0u0ZVBF8VHRkDBEzdYwK/xRrPpZKb
jxtE9NOtxKOhASEDTA81Nu/PgJiPPO5PyF7T2n3XLWMVmqfHw07R7rIqxOO7RoYC
V2dQtjZIBkF5ed7Shx8X8lV6Z2J0gK4TDvnmNpBCPkWotFODMekhsOSHjMDwpAqU
dx0hjGKbX1mf6xPoM7tpYS+w5WNjOBnt5+SVN5sOSOEnzqogRCANtfvZm6Tt+5e1
b6LFFwedNSc+FrD+p5wlxuPgKygjz4cBo9Cwc6ENfJ+3IecvijoX2qRXG5xjS/7r
N7j/Fppb0jEwos81Jfo2wNF+xJxygvbmuvSrSdlE3+jgL2yYn8rSldaxyZHl7Pd2
SiaYM7Iluc1l61cDptqxXFgdxnzGD++jvKSAgaU4L/lVODoOsxsabb6jXvYta35q
F2uiXJzXE4oHn0BrYmqW9G4zOAWNr63Q3M8s6fIbpVG7Js6x+CEGZ99s0bTYfSu2
kQFH86uxJjNi/nFsv+pfC698ucbosQhElG+SEJrqkcFBNq5fvlhQgvT/P+P+B1Za
vl1/SydvjLOdeuBNTQlS7EOK83fDwjjk395zCKl94v+IP6MYlEp7+LD98asdOfDd
2FUduwcV+AxEnAu00AD8ffA+l/+Qe6ZjWtWMFAMRf4EKN4tNNkkKIYITy+E/LUtT
ZIhlXafyCTCQnStjL2jkfojnV0SpxtIcuOlk5ubR/r/AwPRfTKQWe9jeCP3ssbb7
cr+y9jfc/ZUDptE41T3tbTn9fgzugxFZM1uI+woudTdjywe6546ZYgAsqNemPHg6
GBVY8itvApePh674KmP050rSNYdZm8QHjzJBwKrhY7iX2fh17o5ThnB0OGf2VeK2
Jmn9k3qRaix+cUPbYQZC8y94lth6cb0OsYxdSVJcft4LNhQ8bcQ4Azyxi/z2AAuC
em0eqxMN+ufAt7hqq9yD0PtyXdxMg1mcDMashcyanR2Ie9FqvTxlfrEhOgTy06J7
WNqH0FQO2lpQmG0hD23k7SxrsQNHd4S09TqObqpQvptdirYwlH4TH2pvowMMJLWB
elDI6QJFQZ4sP57dEznSD4H0ed464UZpeXV48GD2OO4gQkmj/lWSF7+W22j9CCnY
2I3W0pf/qTZoHAHSx/e6ZqOohBJZc/ys4QrVt4V/1qDzaHqq3HYdTnqmQDQxEarR
2VZxwghZDkJPX9EfHeg33E7JGT3/ImmCovvt8pBaMAVioBgNMk51AGat/RLhR3Fe
bl/h9LYpLfJ+84OnDAyPb7R488qTAjgDWtWb1/J3adLpeNj5Q3ZAzEHXX9KtJY+B
o1bXHeD+QQKvl5Qd2d+Ai4GRn40n3153ppCAN2WqJuuF9x6XAE30bN9dIoGozf05
gei1l7F3XSO59VKFERnmiSHk092UmraMWyeu5p7xxSAvAWQi/JU6ibbc77sFW8mL
JW4vImYetNhJt+6bL3su9w5nLxp1gFlGgjdRpgZ4ppwfwoyFtYnYQXhIG/T48rRu
WzdLP0284B41GzIYvZdyOJIYlnqA5HhCaaffXlQqW3oirzQouwuoi9zErooMHOYi
1p/tgkh/DGz4y77VQDDG6a6072Pe0/ji7wx4Gj6AJq2ACW4LdYl2w+Fv32NvaS2G
+MI9qnWPM8uZlD8udafVA8WXYRr5icXDODBiyTOauhAbUqPleJfjRnu0hw4LL0kh
gpuVpGPch+/fV+E71NWtKrzmMzSP8HYgePq1lrAryskWtGSoMngw1hJJghVT0BmP
4TEOsYqqOnBA6sIRRHVIdR0xyAVlQlZO5p07vMX/EYazr40KKN0vGhn1XBqlXjmx
h77iyH41oeikUSfxqNJLIpZIQgC9fVkkA7HuxKD8fxIUFarbJoN6Il9BopuQbxVx
yUTgnbwzNIbstFG/Af1pqnfAIroAMctp6sGxv2yO7XfYfqRCWb1Xh5nLfauA0tOt
jhxSwDhgyhQIW9Dx1uXHnBgSd+QMWMfD0PUYNsojQpKTsmLWZiH+YGIlS8GoPQq6
p+vfQG1DN2X0oHSyp/iW8J1ME770BjrX6yRHmt1DsNbbP+4aoQtnilGVqBWBKs9w
KI1rSi1nGjEto5IpUjuSw8+Cy+pnz8lTS9GuX5n2QaaGkAiar/0CZ5wNVLdnjVxs
bt5YudSzZmz+OASomQRrrNXf8+LgQUBbc9zJvRHCJETIBcEMlMr1zQUT//pRCosg
sAyzDfhu6vnyVtRLFV6AjsjWHU2RN/of03q3ZVV9NcXefEdJYB2v5kvfr3kFfq8R
Pufxq8XEo5z8iRJN4Jcd7nO4PG4WRaH+WDvm1RuTGePq2058BPOwNS2W+PY6ZOFx
S/zzw0NJ9Y1R1tZsF8KZjcvbu4eB0g3Z/0ZYrHJAyxENl3zcmAsBmuxEwiErrC8O
HmSxrrybqrjKDFIuyuWaf+aFtIKUZghnQdqQoakJQxgOkCfADoTAIvqY343fUElb
lcr16Jsnp/O0Lx5m140Tqvb6dzFTU5AOmjRAhqtakcPVg+LnA7HG0bJZe5iGtJnt
oXbYfLujdPbDggxx4L99aS0KQXHvXpsAEjSsEDYdX8fCaUnZj0ivR9TX92VSruHB
z1DfhecmihFTzCEVVinniTp5yJry6WZDYKSOyzue8TzXZ6RjgP6o8l6NDCPyT23f
yzk95+3J/Qu/LnkfwycCaB3pNY7DxjE4s2zcCTzRi/pTr8JH5MSrm3Uj/Cf2v0tO
S+qWhdvyj8CbAu8Uf+EgcRsi6EuPAMjVhxltSBzMFJo5Fwt/Plyz4TAt9XO7MaLB
7rIs3kwvyKBoagvwi7GHouHszOK2If24WanK9ND359hMAE85HdHICSobyCgCKv76
2J3Md9KgYlJ3km+Ff6mdLOzRRXvSQyKxU7vlgufwdYn3EyngUBxN1SGjRpyWcOmg
0RDJ2u4/dR04PVgxw3xWJxbh0alMPMrWoFDG+sbEscFrBX4cMrjh2q3ToNELNOzq
oTvMzIdHQePrve9ftzQsJeu8EUrc72VJlkNC5XT1I1DzwfJV+jPwq+B2B+MG1SxT
fLvYaE93v0Yl/su8Z4lppa0qyqKqgdjL6QvZZREbt9G8NZYCsqu96+kXp4kr6exM
cNdpyzRRo4NFdLJ+NbCwahidT4gL903keXRaX61npfms8No2Hf5aTv6V7lJfv+h4
yuJnttKFHredA7XLo11bCCDy5GKIgBhkKuAS3Wln2WmbsZGMp9ZXpMmKTPXUQkNp
Ii0V6ZTnQA/Wx5s8S1kt+lY+dy6dv71DOC3XZfyroMWwrkN7d8kbzqn7xlata10n
pfctTED90YOEgQbVf9bg5NxvkP0FLEZdwXIhCoeC6dNw9eSBfnnH0sHPyt101WZx
Ct63JQbyolVj14qZsstrHLZWcXGa+l56x7+rcnPsuh6X1t2XDvfkkXNq7vwOQt45
UJ8G6sfUtybyB14BiNUii/W9rtWkedrwFxKLCx9NUQDDNRSefwYPKsBOPcAejtZS
+WxAfYaWI2svx2K81ayAooDG3raaBACWsTkH6Mj28hZKTjjiuNkcLXmhus3v61A/
GJKmvSPhvf5z7qaj/0YIdnK4a4yb7hHdxE8ZeLEtn0jdeCLeooKtMjP1iO1sabQF
pr/OR/7r+7kmuxSI/pdVJYjR85siuSnV2cNlCrd2Ad13txH1yLSMq2iN6SByLK00
D7J01LNfgKjRVE0/LqoKxgo2uyE0UiQmTDf8n04S9Q5wn579TTZErCBZZv9GDcM1
kdEaZaIwbjCzVDfwsJCBFBCoiUVwAmFMLWKNhqcJaiXQtyYwg9crILC9pDzn9dmq
hozuBsVAz3I2Sgf8MggyOAmoq21Wky5XNHNBpmNUonSxJHL+KTyjE+6Eeb3JXhQ8
wv/quxEJzDOUR57OnhPCsZAKBHh4zD7UZl8v3jf9a+v3kHdoIw8JXhQIzRUzutbf
n3PJ1xIRr7LpcHpMqPQ9UG/d3eSgO4V4pG7QOxdezyXVcqyEVpHm7iA3WRfAnV9y
anjRzOkFiRlgoe3y5VjPn+9xX22WPqmOiofV9kUHvrvo2q1tqXBzYBoyLw3eSXFD
dTV7WDKTxeJnFRNY+mgllnK5ZnMOFmdCiL7FY/Jj5yUMAW9jZzx7wQxMd/VBKSnX
L6CCuOceV5fNPATS0xuSX90vhuWqQ/CuuMME20tr1bUbU7LuAdNBTskmbpDKNUbW
PscojVmOez5Dl+u+5+Kd3+eUTAgOsJTLkqcGOtYnT6ggN2XZsubcQ/o2D6i/x4Qi
10b/mDoIiLF9rBsp2y89ufRUZTFB1a59VkLES/4NjoMnxfUO9YsWf7oYhHdu1WA4
5nQvUZMSexes/hDFJhTYYqA8wrfbMAVD5Af9zk2sB3mj0l9a/iVNZqrIkWjCKay8
uNcast3OR3E2YBKHWgFakPCAZMcxl4WX+3jsA+iIn87jeMfj4HT2WfivZWtSI6JG
DqC3LkWsAX244zDIuPxRlheJUEtV/Ta9yrgVWiOSgjukv/+7BxSgXKyvqrk9Yzx+
qC1m6LJAZccSf99uSZayqoItONtPqjg3xuNnL9WPUJoROMEPrEQCP61yDvZJbdDQ
g+Yz+rsvPHP684hTcDyYDG4yt2i393rjT5MIOMnjPclq9IGOH94kKIPqrKhBT5RJ
rvhQ/BBMivISkOwuwVNwfg/0/iNOBfMsJsTwlm25z5DTqdd4AkOsTlLMtu1Tw7P1
8oUO8y0Pn+sCfQ3cWO0QsOI5BwGPdycRdY3UDtzkS5gyBsbSBJgpio31mGoJ0XRP
+CKhahJRXK8YrX79WffbCKG3pMCOHMcyki84eNe9vqG8oQf5JQHdzP2AogFPDATY
ZrYoSrarZnnSDV+XpAwGlJJBMbbN0RN6auLoLgH74/tF++Yrky95IXbkRJubGXtY
ZiAQs4Gt65+nRLzytdI1IEoRlqKAqJEWLfAM9vhZBhr8G36q+mDLSjFIg3sQtvok
bJJD//TQJ5TcLJvAr9K0vy2rfnAdgDb5Mfc6/KDzB49o1T0yCZBoOrAhluoaAyPU
q/YxussTFv15yziIoa9Bur6uacGorefG25UfdoVU/alyZ1rOpLcf0O7yX5K+lLew
FGELx/HhrS11/8Ih+bLJDZxr9T00OEp/wUQtwBV+ahj3ADwqZFOzAMm+yY+5Ty2b
SXdpTml7METrlgLgsOOeiZZF19a2V6qzVn8kbNpMYVHnog5bEmNJ4HwGpYEQ4fIg
Yi/nRCsJUtzRzPFLb/akOaT7R79M2FPS64IZnaKHBAXGzZ2bn8iwk2+pBKhsW2TU
UAPgmDmTffr2GlQwrNDLmx1nzoR3TmV9L0vNXcck6psQ0UhySZYevS9OuXO/yrsQ
L0Ud44DvtRQV0zA3Wqm5yjSOpsrpSkUXj5/lviAwnhOyxfyTv9S/3DDigTuy+rEt
G98X5kevU6rUOMBqmTXzRaHZsNmOTMDjLhH4mOKJ8Y1N2jVmEmAfp+tbytroDIbY
7Bmnre5jZUJIvtGt0YmUOHp14qP3FHq8Pok1CuGk5LI1NJGlqI0RnMRNrFvpKbau
QTOw49KvLixvykEqaccNUd0WU5c0Hbg9Ai4IKRuyNnYB1896SUXH9TAVvJLC2DKd
mJpf4vO4zk8hepDYR5mFHeZKI2DUxmQWPP5H7uVxo+/g3vYdeCBuqMzsn9WvQ1d3
8GjzdjUPuF13bYcrajjctIBzAJVrzwLuin56/1PmKPYhlLG11gDN2w34UoerAlrD
mAgP7RHqs0w64GBHAeMTeSciMkfvAA3fLI/uIZTttjibOeZUocUQnoc9LMuTeEEx
pgzqQQAMs9buvBJM5iNVMM6bAHzHF1BLrBf5KUvKgSClRmNG5JZDaFE73K+fPkZp
nnLhXlWWdF5GdUwBWa9vsZlXX7JMzzsuBWemT8EeBJA/QL95KHjyWJz+SHfvDXzt
S13vZiXQ88nFMfe+1Ysn5r7dy4VC1n3ejivYWp32o+NnT4mu+kBJFu5iauuzOih9
5XhCZ6zRNeiv8tBjYZkoVWlo8nrJVSS3Gg7lZ+PL9IqUQZvmrIFoGYNUW6v3CKyf
ChwKhGdOPdUsW+DiXIX2q/zY4mVkNyV8Fx6MObriCQHu6yfUX/a0F8Ai4vf1Wkr/
SvrdqK8ZcZGXRpf5o/fM7AIuLAzYxz3rm0/401puPco1YQ4CKtII0DOVUKzoCuXG
GW6HkdPTYdYh0sgtagTLDUkuQNi/FpTsMBfmB+DCF46fn5dY7/GOhwds5r1558Ke
c7vcXUViXkiiG8DF1Kir57bhnFmVgVa4iRIQAv0t1Tv7k5vQO1I5jdsV2UIjWic2
5XrQIeleIx4vJj/BRKz2t+WWPzP3mNN77qVVxRWR7f3cOVHNkAybtqtrGp8ZDolB
JIVJnqX1ehJtoKg1BNRnho2OZPkr2UTbGU2i1vZ0P8imZmKm+OD01m21Vt+QoQUj
LYxDwXUWki3xPrTPhdZC/8fwOllsQv9/9EYds5oF/+XsdXEhN8kPfYBqdKOHi+z9
FuUUO68G5NubcUO1v7GbzAJcz5yXMZpVVucf9OAI4Yrgmi+25NbHvCCrvUy5SUq1
eQShb3cvARZyQ0za8n3Bb6P0NRCKKY+AMg0v28u+BVBUtSfJZ9MNz7ivzabLrDha
TY3bD0wc/E8McumyzTVRUcL1EW1G+pqnPXi2mFL9nWOi2gr2+7/Hwn+eYebgRSDI
3O1sJp4b25xSj8hlMas9k/1mycm//LDjXLN5gon+/l+3UEewGWwOqv/9tK1C+jQX
5eZJODC8y2uMqR3XUTeYjYsvyYqpTlVqml/euTJLwDzOvrf3F5jO9x3eD2FsQkXy
6diAYKHd+/M0wXOTlJhmFJrqQxAvDu76kvcrLMRU8R0LG3aFIytNMTjFyOzwUhNq
9K+dhxEyLnGcRFpl6W60JvA8Wv6iwiWuqP9jPICXWvtxedZTeRGGfknSOXnImgSC
MswpaAGIZrnE3sbdcet2BtbWNisOi7Uxls+5cos84XHjDrMgJjF/rODZptaMKAO2
xlymSvF0vAPBXgtmVH3UkNtbq4ELEHshAX15Ocg8Lr4WC0JhM8LOS11HV7hD1hjP
Kby2fJscTdKCyrX46NQlibxYQhVJOyw5T9d1QhYg8oHt67Yeu4btBEa0BKlQdE/j
sHBd1ltK5HDVRoVJhIpJ7oRCuGwN27j/q18MLfBb2ZlNU1vg7n8bVFSMpZbjxBTc
2sxV8fr99SsCdUC4Wk71DfzFmPQbfPivzJFlGLqQRIHnoMQjK/69px+S5DDG4m5S
mZaLO/VIjGXgiORf2deQ18T99LpGR2+zg1kwMSDU9OP5Op2ufDpMvGHdCIkLqGiC
BKPKqrPjFchc286MDrqv9YE/JfjzoaCZzuVkv/Nm1j5FmMtB/mBkUWkVhARuVfjW
3V3d+lWoV9a3I7lnogiMtLesLl/F996bTTugXp30AJ2utDrDTMinGCTqckxcJMWS
P5Cmjmn9EbWfOTWoFEBv/NRylMYsu1l6diGPy0Nq6KXO9UMCSDTdrKVPhmGVQD0E
KNQwgIeIByBf21CzbA3D6w49u40dJaEiYiv2HGlVhkYwse6mo2HM1B6Jr7+9H6O/
l+EYYn1KEo56wrEmPs5dbvEbgWBKlWLP3nRrZUY1JUL8t6Yb7Qo2Mcrxu2tMhtIN
MQ5+g7TzSACiTUM3rYPhZUvsKYD+X9MZu3PWWIdi2HsnO+0fC3Sh6jU+qDkUZH4G
KQiBJ9TVGX6pks0mODusFhzpIDG8kyvPEga9tyrWvufGtqtTCOtEGOzHBPln5Ijn
FzOeCZqGThzOmCNYSoMpJA9SnBYMSpYTmd9n8Db4d+uorOrlIFny+zp3ubD4s+qd
DRDbkiHWCRGxsbKBLXAdIwU8rlg6wgIrGKu8+6TYsvqFrFphmTuhkB8MMjSyPqCO
Z7agMcgWmOi0odT4kdIaenQUlbT/xAMgy6P3nBRUFuba5qyLip0tWmyUmJ7na+wq
YmOHfERG3QdvzbARoNfzLd5YYEQjXVrLtrhrBqdz2yOKkECxOw/Y3I+Gth+Cv14t
XtttoT9oUHcg9yt5avCws10vzU6ZDspQGOGV5QebAXXqq89LC/41WJfdlJPjumE9
qP0mFHTrQ6zKVmZVHUehKEGvkK6PGA4SGp6ZoYSe8g8uPyKG7eFfMbjNRNu4+JG8
ktTQLFHPKQmX+NPyirjKUtWRjs7AVFxVY/fOSAXkdtGSUyvGm3AuF7sRVDW25ejC
5DwlaYXwWOUV1Eva5ke5jpLZg/k/Abdd4xHv8zX82a7QwLQhJk9XOm5zZUq4vllC
Dkb8dAnA1EMl61O/Ce+ibC5IZH9yT1hmFKoC62g/u0ACCX7ZisxHfL2Wn1DUJip8
lBhs1uomOcunlNfcym4vGfQxqJ1epxpJE//13IT1Z1T343n74wTmLLVIDyZGaaRP
Lfn3dZCJpvOjblkMf4DpygHYufiskquR1Qu1j2djmZVax9AMoncHyo5FyiDX9Qfr
OThOPoFgA+OhW3Ju8GtsXCB6dijzaJQup/RTyCSLLOw5lxebPVHqXRMH+EKNUToF
JXLDBfgpSyylVrwJ7ptqjEO6lXE2xMLVeeychQBlpF4MptGaw7Wx47fuvfDyDQk1
vFwsF2/pCqCYipUkcITKYG0ubKF1fFYKkDAj0bDnL1hUcenoXJAeZUHziDZXGPqJ
78mPtkG7j2B9r7ppQl9kcldmDOT/IK7I2aVCW0qjiqWoOxMfg68ppsHQKdhKDDkQ
eTPqZssN/fJxiQdQZ3Hds5fWP1hO4pZEl5tV3w83wxq/ztyYRse7AaARfMKihKgG
c/J2Ing/FTZBEniNRqS6nYd9eClMPFgbHLDHF4oSoKxAE/Gfg/JOg90n1Vp4VhG2
IFP02WlexnzpwTi/2suxSlo7F/qUlNStTzj9V4yR7yKTypb5FWNdt0WEj36NlLm3
W0Pg+7iKxBO2TEQKPvrERgJsCD607tICV4P7tbaIn1kRHYS7Kz5gtgTZJjMuWetX
Xkxpf1h4OoqnU5FWyBB6DeAPJIvEb0BYku23I0mEld21p1XSnuVOaSP2FCQRC5f1
hDPp6K55btJ4g1Ya5o28SVf538D83+AvigYZeqwFGy7gS4RXPATqLek8pJmSenWS
Pi7JnmK7W63z0aoVGKu6pEXO/NXFJXVWcU3nDMb3Pwull+wMnZ4DlWozyMNbxrie
kFSU7xQfC7TjxL33bBxrZaarcsAthaYBIar+rdCtRJIVvnLVlbdeCpviJLfH0ucX
N9tiC1mpFzh4uFOyT60Akg2ne+Wg7Cxsz6P+pa1gbWQDOz2oXh68l0IOBWvmLupj
TfThzcDQ510sETuq8YhERRKxafJ4ZP05HFSJyXhBq/EVJLAS/XVBEjgx3O2O/2Zi
5SJYJNEAhzmypE6f2YNkNZ9CBcWc06ilfFWnzdRcMGAJJNQz35QqMnobR8LMve7u
fhgaDqnoN202ByB45zogrKTJ0RW4ZTMWIdk6GKWFFVwqzrGh1pNYwkRYofSKDOHc
kuOWr+lN9Hpwbb1NOIUIDRwqprw6w1Vhd/s9Y81m3X5/zNpHe7o6b0tzs8b5NkET
s0OIBwd9Nmk/OJK8J5vtnjf4l+2sO7BBe5D0azQjgc1yDbbT/qAk9XSQoxYTGC0s
LxCFmh6UgXaQMR3cJZkystyTRMdpZTxAW7EfdC4wJ9LvNfd8peUbQhs0G2Z4DL7V
ztURA7JyLVLNocrNPu32vzMz0aTfJw4xWtIBQogrc10aFr5SK5BeG0pWNbVW/x9L
vActl8B+bYb7WCJeHZn9tGlRI9pH9Mh/4Jm5bb7oPvK3MIPTUULKq6mcBord1kzH
kpKR2eBOjKOUrEXgwLVnFIu8AxhuutGUzZY/9s5obX31LiUZ6/OE+/Nm4cngra9O
Vsv3hox9fw9m26wjZlCZWn62JSryA3uMHRSuz0G2OceWQDRZKan2OuCw+wpnjtqc
DfFEdWT62YPaTtfblb+C+cIGYIU8+3RtpfSi7E1R1wG11x4X64vtgszVImtd3Q22
OPN/KllkaVJZPO/QQsws2vqPggge5Vw5C1xNfEtPPTEAOcU8ZlX6Q1ld8PbYrGI6
U+no0/2FV4hK6jWWKbxmXJ+8AYpDKNgcKo73AR426mUdaWDgS/NK2Iw/obM7Vbea
8ciZC2X3Rc/hmsfTkirFxVQptragj0RftBrjbDNjE3jIh4hlSUTWXAoBvorIJI2a
QIt5uFPwmT0WM2PbyGnWuh8rOcpFP1awOkzhgnpjOMrPID2s98dp4fbT1cg3ejjP
UI4JFL9h/Plhs8dIo/I1ApihbT8IYu8sCpM6n1Fscket0YqV9wXGUCbfOb9g47iG
wJ8nMMPIji7nb8eHtsi+7GXbQRFLaMCseToCd8ji3budHSQgQRWznFIlghmBkHRP
0o0zYBcyWezLQkKSj+bwdhAOxw1JeRwSIKcthj41+VQ9xU93WIFp0z4M5Pq87K92
JF/UMyqgeI+kHfj79GAh7OLv13JzerD3X7DbYxwNmFAlnY0uyMY4le0dnjIweFfN
XrAvB1zUgJSXOIXcjyaWmoQgl8loMgMiNqzM0p6j4doSgyF90w4YN8WJ8E4hu7BX
e3fZmd5sqTC72ZwnTP+G5YGhHoVa3o1bKjkjP5hqe9EEOhW5hzQtxeQkkncUJJkc
gRGHI61KSBjLh/TeQkyNRs8LAdWUCytz8DoIBGsmTy/Z7CAKEPhlVrnIdjrrQuIE
Gr/SwEXUNFzuK8A5PQJc6c/81JQ5qiAdeC2CVUowkZmYEbxFjEcdrqtewhagZhTF
X6PHb7u1r79ENQRYD4fq4a5R4JnxrktGDXZrfuF40/rloTk2FLWxUrVbWwsU+tVR
M5/tCaCN+Q1wOTmUhUK/K29eQt7Owr9LFf3mg1D7SitqS8CKvn02MMDKa2ja+vCR
/AJ26wKH7s5o9GQklEjJkzAhzfov4o1bIseyGrUZFGh8jwWGnLK37jpxB4GmTCwq
xff1J2fLLTIoIMAXB7IASJsPuAhLPtwm4W8IStGmEDxMXlnS+WggB2nztV/IA9wx
UcJHKSHX1pUPXdqZSAazMDOiwQwyZ4grfbqHZXRtEWL9UThv94ss9tkkpmT4yEko
tmgquSUs/GfSufsbTppI2Hd3ynHwqzunUVMIzjv/M2W+MYsTI5tQZ9MTlWlzGrEg
7lABZOhgfXXeV2fwLDJP0hyYFt1g8IFoQ5KWsmA/LOo8vTZYfN5H9F7zn3GOXjOw
x65s5h+rnz4DXQbpQB0aH1hb3V9jqt7pz2abcHUaW3AFs+SbnT0LYUUtOpKEttUJ
AE/VXBHRzGpfeMqJ5q3d9j4eLasK9/h+MTdGDyggGDw6uJcW4GRMcVe7stf92JFe
ZkhLFiS8RKmQFENLfPmFX7Jvy7Q2Zdj3Ra4IEwK8rIp4+gEoJcODUwhdD2cUrbvt
wTTPynif+k4pYBLbwHFrlOA74qbSTQRLWtZOZFpnKTxaOq30kvYTDQMLoW7AfWqQ
Q7DPV9jVgakkz/ZZF4CBtH6jr5UL5bLl+SCL/mOZyxbj823raLqC93w+z5xftgX7
P8AYK/aYZDh+KV3g4ndCOIHVMCT/wFaMdtg176WLK3ORgfCUklEJdvxYuPQ+ThCW
RlcQ32Pu7bulLHEBEZ9OdysbtfaSd1vFrxsNWwJ56DsQCefqv0iTgb7iDOt8f0Ys
XNLhq6fStfGfsf32bviUpuMOyP9KWZ2d1kAfRVnGMtirpRw1wpFTvN89TBDIQYjO
OcjumU6u020cw0VrZJbcVxs26Rd3WDoD6GkbIkbxL76fBkFsycZN4lE8NLeipCPQ
OSXAx6kVIDMZyBeVZIW0tN0LUDcVBx8Dq2aWNNeV1YJGr2Wkt6TkAx42tXC08ndB
fwefZefog6Cx5tnX8ydLurUfgONbG0goD75dS1qfX7BYCaw9+Ks3OT0K0Xn0zyz0
YmIDiccXfNm9qQGACPDyAM3ULYFo/wv4Zclkw8i0xtESrO+j8/j6MHf7bANbvVfy
YMCFEZ1xD3ohBAQg7dVrDvXzNwYWwKhW2v3varRD/gPFbdUTIkSAnL0DHJo8JZJ7
7xVTXZeNOhJhPNHb/RTQILuNThaEMPMs9bdHAt2vZUxOuvMBTDYYYZlCZy223m01
Cch1iM152dB0JbSxF7NYnKkYu0vMlmK8HtumY8CfjGJRG3swHJ3hGuL3icN3QYvD
7aKbN17VnzX1s03v1JaLDBsDoq+5XZ7zFPT2oKTotxtPYeMavtPUDiFcHMalL6jT
Hup5HzP+Ey5ypNQz1jytaBGwdw/V2Tqol/hJWSbn47dzZvBoX+5O8PzKC6rg41M7
1PxeweqIG2PDJbDyEBwfyOnu792yhqI20hp92ZjnMXC7gHPZa1L9BNv6LGxD72t9
hB28Rq/ISeXff1d1eUQBOdxAoufHikU4zIUGvp8epETI40VDq5DebM9M8ZVzAX24
FW/jFg8UIWWzr7jKPigrTjPXsLodFZ6RQb7has/qIJTp2NnJqa+h5tQt96j9sOal
KoeesSVvE96gJJOYpTgptbsF7OEfMQWQr1QL7uKcX9twiVWUA53DhRxlJRuMQv5W
SwIvcW5bCL4K49WTPJE5Sun5IuL73C1vk5wViuslEmEAPOBQBFTBzj58ohJaerKX
3HCnMpoXQmeYfVkwTF5V/f4avNLjDNBlLQKUx5ko9gJKU1JhE+7nidJyicUWQPc8
L1T897w8BRq32zmDvvH1xNdHeLi9v3vzXzYuZR8+0z6ngRrrmSycQ8NQ7SY6P0Yj
U4hMrh5t0kk6JXWL39Za9n2GCOIjRfpvtzvo+VgzzoHEBJkn2ZUga4hj7PvKxSUt
xnirvDrlWCZ8MG4KNvzpS23SpK/A5gn6PWD2+D+bcQnSEXY0v1/6xxZYwzg0QVu5
rNnag8WTPndKkBy9CClFGnF0E2w4TnpPRQPq1PkY9P7xWGga9zfiYR54K+eWMcOv
4rqX5UDsg439BOe1h8U0gDWUe/M8nDs1VJatXHpVvzhK8TCmuquqk2TJXDSBPu4d
JqSt8xvc/NWfZNLlmj0HlJsvZ0THyT4Z/QkuW4oeVzwJzaHW+nZHLSllLi8Ofk/R
/un09JzHWk9efWQE/n/kJe+ouOJ4+PUHL7eJ+TeaWOcA4vX3NWAy9q8UlXaTzvbp
QkLwv2XxApmZ2zcPda63FKo4enPNiDqn5PHpMBuia55OHuNv3oVjs47HXQkR3WXe
9mGUbFoj3mshgtK0bijDU9D/wy0fdgJQkEa8yeMxnu/WXpwCPss6xG5ZZPhrnNuE
L67YhnRO05mn6SbGs7X6mxjV0gwQ5SQu3MOKo1eizan4Af6ZYb31JA7BItxbXWIZ
NauKoLEwOS5wDGCruwHIGGb9AWkb7Ptj4ZY/hcM5Cv9qrkQROBs4MCjhcGsET/wT
n4/AcOJ6OfUlspbm6Nv9L+q4FVskEtt3fWSXhaaNsdo1636cT+TO9qnDCSST26zh
Yj/JrxV/7A61owyWjHWMuAB/LlXc4OqPMdlwQTR1TlBncZ/FcQfKegvHvTFQ2Sjv
J+IuXgOTg4FZyHEoq7kkhZlyadcL+arj041pLn0LN9tg8psB31pEk64lkIZ76uo1
ZsyFVSHoh/J6d5zeNUH9C5USZVv/pJSIk0q8JSTVVpAPJBRss/Y2eKYs45D1t/gm
7pF0op1gzKML0ozthaE+vo665mep/tPKamH4pg+aS9HCnaxZJ2itK3vjdI1DEn6u
T1IAs8yQChDTgorc3lPaysGCLB3ggexY769tVe3wz3MPQicpqb8kBEHZBCtUw+Nl
Xoe1H8SE+znB0ki2faUwPhHDAdtoWsI8l0JxnUZAAQhFC//duWjNkZnwh5+6oiLT
egka08VcY1ja4Y+TdOYD3tVrenmyyaFQVPWZdvjsDjfxp4IXC0USQi9tsoq10u0U
/ktPDs68cRLGFClAH5AJHKaYkeZA83Ax3o5NSCsnT/bED8kPMqosPFzm/9zYmMQX
pU8MUfn/S53JAMyhCHHnktAUfbED6JOvS4ZpEDJCzmbsLRw5ug6zhlT5SI7CC8Ud
m9mvh1fa7uy1y7b4CtJ81boGPRdJjNu7LH2TlKZAghZiQUGkc/1QsxZgL3mj+f83
kmZoUKHEtPp6csyfq5YlxvbetUXrQYEKTYuLR9UR8t8jx9Rx3JGjBH11NKoNJ41u
5/TXDkF+01asCGWF+sE2k13FDvG+O84hTGum7+xhocfWhgFw14a6ZbYEgETbQVxO
3dBHWx84OO0aYLxkvc+jR8xQYYxjwzDRzVMjHCP00IIW3tfzcvBcd3c1r6dUPtEf
wp2juxbNaQryPGUGtqAtCtd41mhE12bYto7L0UhgmHufRU6qgk9FR4lGJvwN7bTh
lgHsDU2H47KoPUWOBh7/xwcHDCpcyNv/ZGWJWpjYcKF/C5gY7s2zPcZiu1SVWdck
/qNnToilofvk1csevsbwVfLsvOv4Atd9BbN13mB3cqQoNEC/Eplp8hKoGMgGi30s
alL7R5mVX956qQ386zonT2FwzUp0jxjEuvEvEx2S0Ik7UqgJtx9+3hfeL5j0IgT/
95Gj/KfcdipTT5j0FyeYudg1avaveEm2quCEmTYFkwzaHvRvAZvZH9IhCCL/nLl5
3dJbKH5HDpPJ7A1OYhMSy/dptjejsDowZIev5sJrVaMdHmvTIFQkZwNDdKOYXq/N
zk54ropjSMuTqi1x4eCKQEL/qsGGV3NVTHFoz+z3SO/HAEILc72kYR5RTpEBuwLQ
D2oSDtGIaVM4fQJVP3HLWWARwFb9acAGLhT1uKerNOCFsDlZidoKrTlP/EN90dJo
PFVvCTIY45KMTxhPlCqI/IXMGdVBIRzLyevCbb0osQF2kkg8QEgaM29tQmpux5iR
hi8V/7/hkltCUGo9aMDJfFRJ1zI4LuCFtTBH8dsYNDALfVItnXg2B9tw2TZI7Cc/
EF3kGOOUxHwHyHL2VaqjbpEccBjs0Z26da09tcV+07l/AfktPH28e4WJbypcXoUv
n4zcH3RzzWXZcCBl2zSSgq3Nf7GU1mjZh62h2hMe/fZrFcbE/lQr0KFoyGBDzQbh
oq2Ec7lc/AXG8MNhwEnzUV2rt1wuKVHnJbh0LZ0tiFLK6pIZoON64shHFMaEHC8O
FfvAIffeHvjVBqruKQ0LO/zN72mU1h0KVzuEzx1GM/pws536SWAUdZV2rYQUS5dy
pPrdUltUyRL906ZUO8z+kbwA8B55BwvnLK94Xc6MgZrpUHM8xWIq1HAj8cm5v7mF
i7tcAabWPVIP9H2pVsgy/1p4S9hYWpwLY79Hh3lGSjYI1LPL8QLsfGUYrPAkDiuN
1cdWaA40Axi+8o4HQLM98elXB+RbzzO7huCozJ/Kp9bC7ut1DKr9Z9UPMD8j55ig
WTNvdT+uuvmdFb8CVg07OrkTQBP48inbPCdE9LnKzLKBru0p1qKtZvLsV5f5z0hm
jNIqbjoSyIPIS6WcteUAlwtx/nBdm8ccsO25SxvI++n3c8JHFnUdNYu8HUavLax/
0pEBlwSNYzctH1+yT+83Yn/DtCHTniiruYmUU3jVltirTrMtsmksBCOOWZg8gzlf
16hIkXahOZlU/7CeXI9LanhkniJF0T5VSYaGaokrnwKUGGzItLc2Oaiok/revTYY
swBpLm/dRSPAE7lL0Eoc7KCmsIJ4V0vpurDcDCHW3dn0FfqLd/kIYIKmG2tE+aXt
ZTPj30sio5HaqBO54JVj0cE7ZVLKlDv5wlowG80ZNIqzbm3QFF+/u8FeSxJO4rz8
NsM5AOvofWBdrv1fU6FGF6bf++sLfrYn182zIjwLjVX7OL2lR0KFsFIxWyLRc1mn
6oIy0QosNcw+vnLz/ZjIJM+P14g3KnuABJRM22gKbK7SG8eBYEpByuAgwbXAlc0k
juToBo81njrjbCiZAG9RCyhkIH5D8zZ4hY2vAiuNXT3DenAmF3Lo2/hvqfPEFuc+
KvSkMrNJNmulhpTvQdF6eA7zDCPDYv8YCXL+zQQi1EjkkzlhemoATWSTEtx6a0d5
nE+gV+tZ0K5JabEyKFEynD6geDgRbuV5mOdwI4XM43VLhViuk/zL/wPYkcXfIja5
zYVXpXcTv5ACnA8181gv9G3ghvhcCVrCD4WLTiilcDSuGn1NVzMPWfFxMRQfAnIr
j8M0YoayC+87afZa5Suqz69A80ui0JLxugX5TBlWL8zEhyl4cG2knXiPaz78N3c7
dWAqUcmLt92x76HSHK2Hkx9e9ckHIYQKS5acrMpvTEMVBdkBRI5jLPvPMJ9x6V+T
ZqeWu/JuLEewUSC/jHNhTs8UnOr4TAWKqkaHe1WY2n28fBO3ZB8tsr7zzfbgyDMB
ferTI3U3A3Ens+Uy7teEn24aJUOfAou6+DfdE/a9nW8N48UVmSrqxOmuRbgjRbzL
e/wlgi7ZV2NCrcWbzyQh+OY9xmGwbv0xuDeetoQXOFGlP2e7KJTAdsBIE9Cp61BH
SQEPbWM2dBhSZaeuuJdm++jegVyZ2K+IIrqQRcJejDe5NGVVggzLl4aoX7n+VKPE
Wxoi41v8O2H/d5+3u9U9vqtpmUH3JePy8yRpT8mmmSLF6yZ046rBcNS+QGWBVzmP
ftWzmogQMCblNoRCzW8f+Y0x5xUv92A9w5ShfkAPjfB2v+vD0mIMXrXwkDoWHKm+
Bbi9b1weKe1qSLDPREhiBCXFsHq3KJwHBc/DKP32s8V3TeeoK2U2oInhsAabyJ6p
fRZrcetOU2oZ/YvUdCyjbuWO4fZ2X6JCZPXjPYDZ8/YGkZk2QovvU9o3CIWold48
ZueZqHx6rexwwIDEsxlkcfk41r1rD8cTTMh46NH3bpop+zM6epJP3JIJ87yMgykB
6tbqVPM389b+7TtdAIMlwAJiBjQgSuj0qjDq/JX0ZPPtOKbp+dzHycmCf8HdxdXp
v19k/7npXM52I9uTXrIb4eWQ4OSiXN+1uaWPeVM7LmxjY+yjyz5dfKrZ6tKyqGqr
/D6BdmnyHo1TY2W3UNeHJkySYTRiKh7N5f/QdputN5N9IcWNqRTMAorqUZTrL7xO
Oy3+bIvq3Vv6885fl1m13Szk8CZEg2H4a3VLuYoRbXKbFVW2N2tj1hrKrfzCVFkw
dZzgS4/aF9JvxXmTI7pecMtyeAetHs/UQfcU2To1ptBSol58rNynu7weCPhRAwra
KU5YxFjpP3vulzI2p7YW+erecGHCf9YcxH3lByr0iUfl60lZfqeVTyFN6UB9iAKY
+9c/CrLH4HtSVgtYA7DMshjarDP/gI1xt4Z/BVcul996HHXNY90ROtSSJ+8WpbR2
FS2PtTTGAmCCRCc8e67NhavLvx3Hb6BMknFw4/Ew9HyhOE+ztrdIu/5oU5v/2cdR
sj6fSAffgUXkzEEXq2gip9DzsxYh/51FehvnAAfRaJvt7CFCDz5oG++CaJhgsyjj
9LOXoZ/uFDsi7QjmIdf4fpTSl8jd5tK1PYn7qND6QDhh/JOm4xFZ5HxKIGhV6zxc
72Lao9IGXFlBg5s4aKgnb7qQ7O0TN2Mc3yduF+yrdjri7/ODbOtPZDy5XKzOM3Qt
1dhDpoEyabCIkgWs8jNN/vXnRkeG1vUwvTpyLFKzQFhN8uHmT9XnLcpOMdl+5qY2
eri9c0SOOGoGeNCc4vzJPRj5i0s7LDuamKC98gauqTbV4qnXPm+FR6StWD5WTRM2
olbUNxY3EeJuyVx5O4PytyvP90LHsggIZRIC0IWgBqWKkGZf4CKyx++5+VsNbuFv
xYosJEw/owo1Gf35PmxgX8aa4ENoJhrF/BMuOl3NHt0w//4ZQGL+bS0zxuoWrKYV
umrXIyh2UXQhRTmoFmhADKEiYve5GdYvE/w3ADxybYuxN9z/B45eCgjvMihZerOU
M3Zzo8oGa23bonglnW7+mK6TiaX9qnltz6jzJEMNUTjBTMSnfAIkAid1tfYpcXJ5
Fbud9fu7Fr4LKPv3kUBiPHwsJ7y47im46DlyjquIw9euZYPGoKqUa8tFnEqxn3iM
7QMBY5iqHtJtSFM2wDnD/EzpI2DgvRnnuaHKkeKgjQm3GzngG/92evlOaK1Qu6QU
HxE1tqW0Di2KdoEIqodC7D0Ou+kyW0QLoHl779+rwU4ehPbfrTtPFuxSK8c/8HdQ
G2h6Kk4llyoRwzkvYgBmVsM4EwDpitYl/DU7aBz8tNblbzVXWHfg7OK6X/hDfVWB
JVXjbkxLVTk3gXPGYgTPS4p6qaAfxwU2ATQVq2lOlCs+KcGTBXTAue+VJj2zsUQF
9W45OhsafeOZW5/+VhUVLU9ZjqfNvEv/6rzBqbowZXVrsAK9St7D/Dil17OaujWu
TK6my9A/cXK119ExdGd3rsrLjcdoYHmjlV9vXSJwq6SF/NfwWstolxsByQ4RCgsP
IsVowiAiz1Ifuhu4jF90riZAaoRLj0sDmGXz/CPS28S6xCxDyVJLLKiG3i68TKx/
my4nEVQhYJCVFWKm52MjaAxD0DzNU3pYEcXAa/10D0oLYv9HcbhfefGPm3BoC2Y4
QrAQVVY9B0pb3/QKzLnEa/LuRkZvC2B9H+z1hYY/lBxC/q1p+lyM5G32BvVbWBz1
pLtKgr0doo7WI0Ue9wQP1XgSx0jbyT2tWgqP3SRZWy/sCoklS8Wth1gs9XCfbUf8
g+Lc21qz+c6q7ybju4IQLps+7Q7Hx/SRgWF+9b/O3PJ01b0/zToYEXO3Y05Wx+Q0
Y7iV/rL3iqqUbCB1IIrTdQSZFhFWzcykDrofgAW69yUoudlXx1xl+ESF5nQVgZwR
gNj4b12R2v/rqdKIm7Y5e7vsAe+aZdVytEvYaZpX89oCm1PzEDBwEQ8NpF/nwEmT
wIaPMH7Z+QHCvdqfr+Iy/yO+wFKymZ7tuLl6bwsgvhHS//JKeBj8zfQnl8KjuSz7
WrxbVHMC3Qr3+S6ISohK7xw4UCIq7vqA29SKt31HgX6HQxGdN1TIcS3Sa9PpdRCc
VM0VIE9joW+bsux41IX1TLV/1A/E9enGjxrrz7VXTFWvX7l+0VHdW6cCIbryTQmI
e4KH86dEVg+R7oALrkQkP/MTVTfhJ7ubu9ozdIRQZcghmdS4h3Z3zTJAUC9i4hQo
pJy9jEAHBg6k7+1vnLcTmPNpUFIQDdXXtZLOOb+JsIWV2uDlnPdOC/raHmL2y+uK
d62pC7Z9tkt6H5VpPXR7bEd0lk43kJGZ/FQhSlgMK0R5WAlYgjyKnGgG0h45m3cy
js1e1LjKeCyRnNCSja2dgNHeYIK1QTy832IOG1pYEhL5ASR4eTnjDtV9ok9dWpAZ
2j2jCQUTDm/wAYgnh4bmvcB3mOzwTa1AsC6Wz3ZsXGOIQ+lMaly5CF97lb+2yv9V
tBlRlOEcbHWNDWs6EFTiuBOru6jSLgPjJ/FRq5RQ/69t3vk2N5P4UC+lpxF6zaXP
Gf1CJMR+wa4ijudtEx+pIhiqqKhVQp0WuM6tvAz9FW4ufgyfx+BhJleHDe6tEtjJ
i5ELbwxRoaCQV54fklI5glMQ0yJjF8TO3Jq6bN0MXaf2LJmjUrnUZ5dY/dUO5bcK
A7omsu5o1x+TDVyo5VtHqkBiXfrG+cD0JVnli9grRSzKazjyAn2ylqT/I1fXtoLi
E0r3Tmgt7U9FaiIKJ8rR9KugBElXyGNnZa0kdXrbq8fITeTVQ5bBel4rAAh1jLjp
KHFFzO/N4+S4uMdjxtUz6Oc7g3kzirGUULrl0E/IifVstv1utHwY9Bf+nHBBRWhr
es/hD59ywDoqY19uPmCurNrnz6eQm3qZv3qbEGoxFg3F2G9v80gnqQJTJuBNKwxp
kRPJZ3Ta/VKEc8vg3pZAwbe/CvuNcH4rN8SyWR3ihGtnPysEJXt15ssZQIoOc90/
+Qe/i83S8JEmhHlvlbsAayv+rVgQvFW1jxYj4ebrroEx35rXJq0oOaOiVdarS+GN
xkbsykncxhIwIdQPu/MQ0ff/KUfmMBewRDM9FNDkHLkc8P3BFSYmFEvLs2Nmvxzq
LpX2O0GFB6gRLMJvPiKjNRYP+AAxYEDUVJ71JVm4VEbRhBa1mQCfVIVt2UKAHGH2
iYLpm3E3G7EI7831ysyC2DNFdgYTsuXqQe13OxDOfHVMNgfi7b10fVsTSJf5p6FW
IckvT8I6q1QVfeh+gqf3EkxhZpim/t55DHU4sq59oBMG6WumbvooGy1B2mb5cWhp
jQI/sf1Zey0foYxNoGIAYT5YmxyK6YBDohjqXSkBDUCvD+j19sxaS8MprH0u/9zd
1Dx9iJO3WVjXdgNVINabrgK7cLSSHOQVFmVTWGmon15GEkryTDENct8qqul5pwSW
RSJ8tFhXsSWbcq7lrm2NLBgNzx0XQ9T8SjFh9sF/gq/SyGk+HuBBqmJVmDKCzBo+
SHgmicjZdNelQThSrU17jBp+mqUvr+2i+SLMS9N5O40UekKy85FJqdi/ayaQyKAV
0GwGl4PQ2Xgqi/Ag3JyV4qKxYI3WWTLvW1v83wkIiSqATuXH7g7OnVuZurMjVTYS
/rymcdGoK4rXm21Wtd9lIG9f5Q95fnZU2Q4DrWy5V7UvThKDuGq/dInzXL4NnwBJ
xQ8T/AUyL3KyDwwSaThnf8/+ruXyzYVwp4kkUAPGF7sBoA4JhZ+t3G+e9iH/dZqU
jgsKEW4m4kZ+JM4o5loCDh8yLfzUkjdjqLcLqvPtFDcGUQWRFEDW7cWtlyi9cFdW
QbP6z3qK+u6FNFC70hKMiNoaueTzEy+ub2O343O4/eLdWVkLP7npzwyyGJnbyiPa
EI2f6gMLxZt3/M2F8WqLOZbbuZQ1e8MlWjCQlOOnlVHTs2bS5rH6mCRmZqIYrJGd
d76pMzcmQKdwcy4YbJnhhI6mvc3OJM0nXlZx6MrGNqq/gQdNWXlH0v4Fhc+ZLLhE
08Y+ngbArfLYBqBATtLHthYSw7BCx8ai4+1cTsA6K8zW2zHs79X+RmF4j5DVhT9V
MdUNoh+nvE5UfXeijzvHaueDQ7HupkwTSg10Ccxnq+kT4jk3MHrgOSR7l10vV03i
b/lxFONvZxLXwCUYYclDGVP03Wdis7ndlpFMElzZDZyS+xi4NITbWeanc/suZv0i
Y06wmu+ssOleAK5NtOeCGYX3NrmB2sbK94pWKNu4brnhyHzuHxd7vkq9pHYxDZWL
Jw1LE78vVM8U50dIKOqrLPAzk3cGsqzCgxXDyoaSf5/gZItxgIAynQkXHEb8RIQf
ZzS4Pq3NJG2g5hasNMRoi1QpVOgK3f89VkR573w/dU/y+aXSBf1hAQ9uuwabxbUi
d9rcMbLiCO32rMrfuovbrV5ea6eb6sL7VYFHRtoukgCEpREvrO05fDkDbUg3v9pc
tgM4+u1VSRsfWuTEc7ypPkG8cpJuBseKv6qhZQVKCNVUIxO+cA58GISNwpFuU05B
sB0ct331QbVLdfSy2cmn1zFUbmDiT6cnzi523ZaE/uUmN3RbHLsVWHL8im0FPUKA
PRoE0MXFrHvPkdYBUtDJ+xoT2AmNmcbFAc+ynOvzkCzHwaSxNcy/XVA7hsUBH3AA
Q3OCoDbVjjQ2i06zY64QR4/qLnYW2RJBDjQVbtARG6DTgfYT9KNuBBITrU1xhob7
0NmmQXk+uthtUyEBvDt7Zi7NXusq1qaM6L2qizZMdfUnPVSIbxzgPGLEZozxjmwW
sbsGeg39FrwGjp1XDGl07NceNa238e+R7WfAQKaWt/bLLl9KG7LKZc+QU6s5l4NV
+Wp3fyzyS6gontPoadC5pZlx/xsez72IXf3o+Y99fIz0Gu5MBkfsJMiT6xJlIeGv
HU9Ujvdl8x2vFQYRcz9NLHzTmv9i8bgD/tN4PyCGRA5PskvqnoTDiUeW1jJ8lXJC
ZitH1jQyTyQNzzA+YQ9vTkT0bAQ3DOVcDxc6XNI3zZA7/2KOkWtdoBq52xTmh8Pr
hnxU+0hAQmYMVPsE9JUyYpL4/r+iFCIOV0XCwHp/kOInWKy36Px2alW/Rr7GABhQ
XqHtDzvj/eAXt7RaZ21y/giIXYmDSZ5dwNKJlikgVTe43lxcmM5tyhr1WqOV2LN8
9KS6jP3HgegLZxheMOeVbzMQejmV8goYFcJKUYDN7jFlYplkeWu2v+ZCfMICdocT
WRw2Zh8gY2AdqkXFtRxArAevQCNIAcTmd+aF/XqICxW+zQoPuVKJzEz+KrbBTxC4
XftTbIdmkyXzgTG8t4fYUjF3c5EMRCqDeu/dEeciSIbfpiNuBEirZLpoIs3bERev
Sj1uONUBwsk8e/bwSDJhiJ6Dz57bSHWqFevtcnYzLN60BPBDZ+5mNVhKtlkgKTND
ZdG7Oon++R3Vtp+zeHSm/GeH/TDbBv5hN3Q2X7HGHgeNu3V3t78x5CVWcaoom4T4
GQkhHuhjnOBWOEfVpRnb4qGi/fc9q7f6CDXclnNqc6/+T4768XI4Ct3UQFDqmjKQ
jZwquO/ehFYlNkaBflSle3nupxBHpKcaw2PB+wb76DCsyboS8D0FA42DkIGUpQM8
fDNxJH6w7bbTd+RtjNpUd80EvqhzYFGTd9CUOoT9aQPSBLJzVroieWeuOwCaN8PW
yG5rdHEp2bDLgWV2suGClhQoz3EfxwbW32mnRJ1ePX5rl7YXSGxTtmY87gr0DlgP
43M64aGGE6ZNpn4NR9Z6aerR8q/tFZfVwB3Oi8fYcwAFhfCjyDEQukKOkRqoY5Qe
HJ4zFLDxv9VFfNKSsPxD9P9F2wo4BX3TC9OPd5q7ruo4PKjvdA6YsVwHCKmBX3uw
PD7myoVFpHqrYiDzheYYECRpjDCJzNPLQI46M1K8lsgGXG1YcW6o2sMWbUK49ct4
QJ6b/k9TVBc/RHBn6e5utoEylqu1W+tms07YYMLjJlo+Fs+WmO+7tBs1gcKYOpqI
uBYYkFGfzrtvHu1Dk5YacoQ1GRgDRDPCAba75epdmVtmVG2iHS3hA0p85bOAa+f7
PdN7gh9KRcFYKPxBbIlIQnqQ4pXaEKbtEfCT2FE8ieCJfNiBmvptdh//PU6T97yr
XMv0diCyOWugUfwp65k3ZHOZ966EYf5wmBml5zXo27afnK/DTvC+BZj8YB66xdqN
9UAJLvETs0v+n8uPUY9xLdSOTjYWFPHbd36KvUUzp/WQeFKl2ueu8jai/tp6upqE
Ee3htOdhwAb1H6TSXiAgvM21D5bmuqAPYPhfFyrJRE5krbTW5Yydok1ejYRfaaQU
ep0UanAiQ5tPFuvknrQQjf4NClbiw4FvabrwHx5+GxmqCw3rzxcEtXgZ5izloOsw
UDtfKB6bAjvA2/fO+pLAkDOwPXRGR5sjCx971iuGNSH2p/jYrj/NarqZk+q6iiBm
r7xtrnQMUY+bHOmAi4b6PjU1ZrOnc9GUTbSTTovLU3OtfMk0BFrXzY2xyupewe66
zjgT39RCuCQ/fThm3zLx0Uf+4L6n8tO1lvxlrrMX/uAlW4VWLGgaDjQP7TkFoGO1
dd3N9o20DkiehA8CveQgsJ6ZaFBT04tJOQhGsLRhK67HRjjpSk7ArxrICflbtUX4
/wMHGOHzqTA3logbZQrxqyW7+NKOls4dhCWH8tKo18GFYamd1kR9tFlpm3uSmeIk
2S9tH4qL51O7xxxJHMWnwX3ZI8O7qMv/uQBJHZGYRUtXTwkpt41aTr0odCqkQ673
5ikpRJTCmUa6b5g0Hm5ShaD/zDtMVemH0WHwKCkduOfdUoF+550Mb1e5iPTtdrDi
1SR8DF4AeMuzZ7YeLblPz6/izYEWZbe+g0bru8P3TIGRWJDpdV4+vLX4PySzptDv
SUjP8f8NXfaWX+mcVQHfwc3Y1AUE6hED1k9w/4i3QtsTt8j4P4C2Aj5gt3HVD9gp
LHtIyv9zw/09Imkv/4owqWCV3i4TY6Fq4J0XrOI0sCI3Nl2Qi+ybogpJqym457BJ
+rqYH8n1CB9H2MLZKEQXNH1unZUcM0nhRuABgU0+hbeElaiPISI8p2QkTwst+nkq
vW8WsExhsC+FUnYpO91hYhBPbExsMiQ9Cpkz6lariW7BULSWrqm1//BvfJCsjxJO
PvKLXVmsw5q7AApnLsjdxkWWu+78yq1NO1PPgeJHwUe7DacAVE2rgM5ra61b5fuy
RMJBQcG7yM696u551dGeNRMYxjKLdr1lMzcZXWXw79eiTMwYX7nkVxYbS8k8YcU+
XuK9jq3Ehht22FXvqKaBIpIG9H99HxFe/USVMuDEAGxGDK/qsZT8yjY/lfkpHZq5
dqso8y2AwF9Jvh20xbUOX/2crx430CA7+A7f1XswsXzvU8RStP/54ee5CQLHRsCn
+We5JH2zV1IIllaaUaL9Q5e1RfKkh+lbKNzWjqYu3ncPBZeqFIvDDXrElOotyWVv
uI14+qFaMbnMdL1snDPo50ncXN3bpaYmEkws7nIUr9drBFLFfPYKMPYoOxiEAorc
2jIqvT30Zq2TNGuWEeyQH6oExg3nIPtisV3WpDLFtiAP/zZnIdY8vxYK1Oa1fcBf
tewMUcwGEFGm5r0RCKjFlSfWG7hzOJ6pgVJkyWh1fOqDJIssYpazlVXjLspUA6r8
ueLxwLrfEL+nzOOW8HqmPrRWgWVPt/HgMy9x8aGx5+It+Qj1oBNo2B97UjllIAK8
VU9wXNTwMn/K48rCuIpJLu+O4QDG6I7TuIDxq+X3h9Ci2dz8Sn+ZmTafhHic2Isa
EGJk/0AcVCZfK2KDWx4/5EpWy32ntinPA79+QA6BawfhUGWzaSm4Wez8//TLoUJK
nx0Dorkvf6nOAvgh9K0MvIKNJMwa3cAH1WK+4Nm+T/m7T7sSLWPdPC9q1OkPD5u6
tRukT50Oq0TVF3WC5+jIAm2gZPqUZPrdLF1dVb5YQ7LcDvBRGwfaFwQids0K9FFN
+or0ftI1LE2dfKJg4WX5twNJeZac4pMjs0RO/RcLDuhYVfwXrAKUBwf4r8KWB0SJ
GsKug++EZnv9WU1tvuF+lSXBMZ7LTr1O2n8jwWlXh0Gaa8J9rMjqYdKDnzIsa5tZ
e+p7a+oscr6HvRu0oTfMkVfAIl+H5Bl80FHgMCxGDmIMgBzb9kihz+Z6xOtjWQMy
y+E7sGb2VtUDhZOV9OPaV9gF+vhyY//Y3cXhNWcY4ZK/H1uccpmeTLfYDyWT2UiN
Eb6P9ivRZIEnikwx1ECJmLFDJGJTugMusvFoRq7F1kqW0UM/hsYQlma26/lLgpxT
WHyGFtYKQiZv8ZRiaubYRXZND3ru+UL6+1FrcU7iGggDnQGXCrqWNsPtmu6Jfs7F
/9DuURgN+tyNg4NtQ019xS8SHVlte68F+l68RpGdFf8uPHpKy/q3D08jE7R+eYFT
AvNDqqNmXDEZOocV65V/ijxvxJPdn67MhEselk7YgTQ6aai7HMTENnX+QjAGJ+lY
AWDr96L6txscR0bnKOhFEMdXofNkiFM2bwZjABpPTxt+nVZLG5ueOi8uGPb5hDS7
IcZdjOIWTQOgmYgjWHz+NuMnHesvx+ARYmirDLvjqcfT2DKrQasGXU25HdbQX53E
f8X8GCwsCMBSdBOVAoH6K8J7tl6e5Jv7tcuKARnf0gn+D/2c0Cu24iPBhm/KdenP
lnRDXe3Kc62EwjH44hm5/0Ek9bjS0NFAmjOR6bB5FOncND4QcbYkMiuNBgRH1vd3
EDdUVBtHQ/Qf6PflzoHbm1zL4PMx4fx2hFyLkC+nFiAKSrRNsEtnRWACw+TmQ/Po
hhVMZ5q8B4ztq2aUq3ORd26LmTsv9khcpOW7QWc2VrTE9rCN9/7e/v9CCNydXdg+
hpc5wfPeI1Fw5W5twwnWV5XxCN/YMfY4HRY6oCieQAHuLZF7iEYkkxBxKU40/x3P
q1mni0+NETKwLM9yzbfTvMFNnYhZmBIbMxZjJwxY5bTvokx+mgaUUjmMD5UNpa29
EXXzxf87H52BqMRi5TY/cjGtb1+SpnwtA4yFN7a9kw2soha710FMKXXLsU5PApuf
nujh1KiHyH8VLbd8nwNO2ijWTOlTRSDr7JSlaj9U5JFLRqSNd0T2fQDQI2uWZLXI
oh8LjRLRzeT4VoCV6rbtHJJEHcr1LXkNKIjpKK5xkn3e/G/HXSUCjGLFilKFN8uj
sVkYJ2RQHTkXZo/xXgIDpVMMjVzXklFYuYOZNo5Zb5TLd5jtdsJ2IfBizP1TEzw7
fN1qJrjX/Vero7tlsV8Kj2ny2Z959u9q8Z68XtpTfbZOW9YErbNcA56Vr8bMttGw
li/AwLBmd9WHlPYvrLOoo+o6XvDh5raX5PIzZjBjwXwkvRXVz8qYa/XTh9G7tYhL
h+wn1BrGeVVvfORg8D6mnBD+IEvyXSP6/ptHlm6LQKuEsNDdEqfk277tGZ4t8SdX
21Ay64wpE4kw62LM4vyrM+m+VHCBc1yKUU4P0US50IUXbM14Wj6mIF0sa8bPc144
aFzPppluT7J4/bWqqBWpjtZp2lWDFGZcZIyxLmhEdGr1n6VTVG+p+cFSg0eBRVfl
ctGF82OuekpsEpSZqJvIO+Yp0bzww3DorA1RJ7/2bSrelbZQCn1ths3KWiJsQSIV
YNpD80EKRlfDIxcPhpox8HTZc55xh/FeePTguySIAr9YxpZ2OhDKVLqvinPTyQBJ
3f8uLMu9uYZj65CpuxeQ0gtaR2tQ5eknixqV8Ll3asegWpv/9F6sA1VOGtrTthEU
pvHUBxJh1NQ66y0MnTYwlJpqu+5TURwVFfBkyqCB08OMzBbrAYPXs6iY9rL1vxZZ
lclzpk6NmxpSUzNT//KgF+w/6AEbHzxHyVWQrrZlr1rzo2bXPTQE6qf9s9G9hDrD
FlonJ8pYnjlYQfcVFHVLNj2SVxeLEvBAJYlum4qGepddEShoUSs7iWd/RUJNNypD
Z1l1lonuws1kI/1pyxXkIQ2tPVxJyvEUpgtxi4Spa/T8TbOxceQavcC+b5VmJSS3
7kAS0nokWvV/ytfByuoF+uTeoOCT+SBe277QAHnKkcVLcsvLw2qwNCg4kNEEwowg
V4DUD4ZyhbZ6bexVRLBfTLhPetFvi9sLy5UMrJbI9BnJBMFr4CIWXFo6g6q8wstG
BnzcPZ5ioCJ2QuSW/jmR/dwepAIexvFe66Lcme65jnfVNaqC3r94Z6yA/I/B4vg7
ekxp0oonIPfB5kHqu4aZYQb0DDtox/eSXWVPBOjiZqtal+6cQDFG7jV3uFm8wR8l
g86gwFUx+gHy91ogHV/RPywOdEwe+JryZDf1gOMoEU/yVAhAbZYtCVaXiwmhywxo
qOY7T+ok1UR/3EuNICyNxX7z0smhxP7aL7lbBDAAh4Yyc4S+fwMuCefBWxHf42sZ
eT71uNfFGmCZ7LArbvMvhPVvmHybf2KONo8wLlsBNEh3tcHWLSF9mDnF0vDVzw6P
YBWRhnOEcZ8y16rF0seAEhuanURKH2HOmx5qcs9KW5BAesM5dT6d8wHQ60f0EAwK
bUz59l/7Nk+f+d0IjsUK8cgf+V5UW/Jf2h2nDt0HKg09fW9fKS/ArYTecBWUCX3J
e0s0fF6CPqH4+HInA/OOOXCcirw96Hy15nh/ToTSijIKJmQlvVQ73gSl1Gn/zBeh
h6LP+ERrm0gov8Wq04IgzgDumLsLZTTe8XDZmRiD68ietDpCJ51vQvdE0TftQAXI
h2kRa3eeIZcg/vMrXXbUujU+DsZRdKx27NHdQLP0DGDOpM8owD1yVqno9fJ1hy+F
AjzRdxbezic1RhNAGtSPGZAB1ZkzrifrKFJY6KDLegRYB2gRbcarxn5vRT9zOYPI
SY7grJwtKEjaL6oIp0g5Asl7ImtjCdR+moWnFXQDgX/roYR0IbR6RXHR/LNtuP0j
icex5a0so/iJ/tLJfeOPsojh+GrC2WMuw9rjvaf8zxa3dRstkRqNeEtBwOnnj+zz
FiQV7zzb8DMMOalUiQdHbpvFZnmCfzrWdUDmD7ki504jCHfrT+2JI18B6tPXm28o
77WX/LY0/u31PwNVaiecGzhD3miLmdDIage3dYOAUvz2rubD1BbtZBqJE29OB3SV
F3rYi8x3MV8d89isMKmlwQW+GaIpuM+yroPbixYaA/dcFFwXjU+tfI+Goku8GIbz
zYcfjPIFhnqf8ls1sBdR8/5BXOBVCjQJZ0OFBaMy7KuEw0oon+g4nrkCUUys7a1z
v1ZVZZ94gmex6BxDWCby4V+oUDCOgpa8eoCQ3/4NxCgBGprpgGcn+w6wfyTkhcdw
uKu3xgdedcSY6fz/wKgalS7oaVP0w6cNeWjhZJvcdVpHdWAOhZxvw6NMpHc9P3f3
abS3Iykid/pezWivobjiLw8cPbTIQYH35W1ucuIkgEtyqs2fj+1BNbJ+mzc2Qwqv
rlKIsl3PObobI1uI6e075OdMl4RTko6wSL5/V/VzRxQodfl7zjrYxv2A6lYEY7ug
iIbBFn0C+9GvtHXIcOWJK6B2ZH/zpa4ZjrWf0ZOi4cC9OzSLFHW2W1YlunfCrCOz
8Go1Ylcd17EvM7cOd6APAnKs3lQ2+OUHJ4go7d/Oc+ITjbc9yDFJ8BByDH+n+TGb
GRXGzEjYpJ8gJKlcOQ1lj4P5pN3hVtt5AZecKNm1AMqaT5O7SL7Ct+y0bQcWB5zH
FalvaM5g+HmLTbl6OwNFHa4Fifyf11Vtx74UUkaBX91L9TndgsXSPvFJjGfmdwKy
Uyxyv/qWXJ8I162LZPjvsMrpMlO1ueLurOS4Ooh06fvc+AgTXe1VzcV90Uxf5XDE
G3t6++PVXkSK+G7lLJONFbSHSfbL27I6NzRmPfrsEW7bhNdAN2XQE7qsw+dFTLnL
3pnN+EK6g7O3haHtHtwzZ3IKEbGvVaTudkf9Ecxz+N4Xlqz1atKE+XcDgQrZxB3l
vgSqZxx/3uNyJMXQULC87MRxFS4mHgkDBHJ9IPc/nZTAUwq0DcK/alQQA2YupyKd
15R3acR8tFCh5WT8fcrY4TemHAfchozqfpaDYTAdfjEY0b/87wbHps8bqjdWh8rW
Y4Gg39hIlsxz1pOeMWXupr+jmBPWqjOd96R9fQQGPISCAztlvIWh7G23UT6/VsjB
PeIakMZLGA3+mFDpvsb+8UtWDxLoXTaX/xA2kNURNxpxFXV4pAlw6pamDcH8dI3l
w1VTYENv6YSPel1Lu1NwTaxfCUXn7XUOBfwWTqIGVleMJ0bJ40zMK4kbXpngpv8Q
vXVyHAzkbEWbQ79GZH3e+n3g23PhWJb0m4imP/KajaOncEzwXeePMnYb6qV3N0+5
8ihBwBiCnxjKxErfpqXwotdxL8BR9fIPUdCQr7Ugoy69EL2nr3Fshx325dlOO9yC
GH1F04wvOr2uZGr/PaQaEmW4FRK2603bYJrtRAEhdpX/WJ3pHTH+5Zz+5J1KUreS
6iD/cNBG2BqnzAqNasMR4bAfffqbLxcp4+b1qzsabiRU2jkT38XO1Eqa2eMRIIUT
1eligfs6D0qsAcOf+NFP1sVdSIx3txF1/sbbZdeLJSH3ptE7gl0wLde4HjpgGYFn
hZhz7Y2ZtIdOGqNnPaeTfeRpsTCiExnwg1Ex816x1eJcQlPbYsu7ljkKQrNIauHy
O/FmFoCTm4fmDyhlmKubj0094GOC39QddrrEv89yWqF2CUmFBFJkQ2L6qXzlMLy/
riJzhF6uFw4vUoByqytVd6fvgeJgQSBRiB3Aqp7MILb7vzCtfkTHAZzGz2djNxUz
h8dWfICfN8Cyp88nUQxGqEgrZkviZc4vivx7TQaxbymPc4tfolayA+EYkthayYV1
chRlvhBeOMi9XlJeQcQtphv1yI/GsvpfYelpeBCOL0suPwDRjGtKPWT4mbBAlFjv
Me1427CZ3C213+zV9UJ1PyWAd8ajUfOWFwFF/85Xdp2PxEd4PkahAtT+vYwwiBvA
F3DvsXj43KqyB6zN9Bt/rOWMKv8oYo3GfW9sD/GQAd8U2USTyT70vDlt233t5IEI
yiykdGbFzxFE8b8oy0feV2QWt4KVACCFqzQXWtDbYLwTpo1VFE4QB4kQzRJI9daY
vlFgeu9B52/U5dg8lyGVuZk9Q2fJR/D1Lr3GwAP7nKu545zJxb9tr+EgBS4+Ak/C
SlQiJ04Pf315leDSCGT4HFfWtaIaCdVI7KLsDZmFUE6LdEgBmPOwHUBAUjPSRO0k
E2bwrFir+bRFq+G/CCHhDOSeVuOi5QI8Cn253/yUeWa93HdlnBhqU3UZjylb+Ikg
69fGdMYZHSgtjU4+23PiBYdC5iOSEI3XFY8z+A2aEfCVejm+0Uob+21cgmbBhPdI
Mlofm1xhAz7LBILmf3BeyLSx6nxSWmIJZ8IIA4Z9oGOfcA6NPMy+Eq6E8t/P0UEF
iU4iz3e2vSk6eir7oba87Bq3sARF6PRD3VA5gK+Tmv92cSoPn36Ex8Gq9ZNpbHV3
X5VnDQ9imrb3Ky36l1QVDMAi1f5GXdwQw229vHC+E0Sqr+KCHnx8BiwNcYJkQDsV
JVDSZb2hTqlv0jIKq3c8FkkFPGd/5psz8eHZ9NjfrTRW8InZXlVbNe0G8z89mby9
UqWUbiLYx5UpVoG2HjP/VxMsRzAh5k/z+rP7extJUAJvyB5k0gFRAEHWhGZ6uxnc
zBhnztYyD5CjA50Ixn4JaancRmgOLIUJZkO+uv2/d+5BGAR+IKeWUPiMBh2BpC6+
bRnOn8yyHV/bL+OPFE1J0liTm0hy3w7c1OGqjwvNkkpm+GQJwkWTLKDmh6LK7UkX
LHkVW6SLT5MiKTW65JHH9Z5+43RFCe9zjSdxua+7R0ycDcWS/Ey7IZgW6bDhQRBV
Wtj1w213m/hSjBMzVPrlXlQ8GK/hljLQMb7NejzI8jAsheuv7eTms9hx2zz2Ced4
e1S8mbC1ElSihYHjn3IjTAaGGCrOsk36a4p9GeQGl5QCBTBLUr0wS9TMOuBZJrzk
3zxn4apoY0K7trVSFM+0KuwsUrOqJ0KQEoGPYO9XmmXL7FzaSeYVnCjW4Uyo/vtw
7uaZubFHJjfmk6fjpbGKc5lmAKebCe49RnXOfL7B86pN8nd9Rq51SUdDBC4PstBN
PgnOOQXRSVY9NRj6KGZVy5uG79Z4bcZ/TtTkpHpSdU7LRISKolHtxwKq50idn9Aa
OEIV0BDtnwyQ6aMWNxn7784HbeCBZEkBnSh0Xr2JcHAvGvIrcl81ZWIRQEWX6uye
NBGcKtY9qE6sFk9XAMVOYQkRR76QvUruigiMVjpUCxtkGfhOr2c2ZoV1OIGmJY4Z
lNFpedz+GR1p5DC6kxFM4NvhxOt+3r/wyo606Cvlqkx2rZ66fPFIiGtljCleEBmB
1R1ZC1wt2a1WXdfHispCyATbQOprKVr3cO3j+m+tLrTTuwKGsAxjSRsOys3ErvH+
filgGTscYLf7cZJAIved+XTB2YUjC09QhtHyf/Q78JFSPaH12TsQxKziyKH/MS0P
UhJOIEsxcIunhzBT+6ZPvEDp/kCM2Gy7ZQUqiHLcqCvi71rFy6AEkKqr1Nc4g7sE
qiP3flC0v2pu6Op5u0CUqtWzZcYjmqe+zgQlKw/XgSQtI0vF2B8pa6uccofjRqns
um9onBjVebvhYmtqPybkJ10ylaUXCeHDOOmnVNVxL68vqqH8VS2gbcZ3NTIqY+Ke
OQuRU5WxfwnmVlHeBAOwFUmc93XBcE3LDdLpaylextCBX8kVCCefWoLo7wvubx3W
cNPLJyzJI11tQKDg7/AI0coyAaOqlApKcDVHhOIOqz1vnllkAL43GsSoD/CBFThP
1J0dBjb+9Z7wyEyHtwpSfSQuoCqLT4lhjS1j9ABSy+lUtuLQWOMjdI8mb2Ms+Exk
RtwC1tNMFBzmJo3xKbRC13mETrhwA/NFqlX6CPsGMCGTZddQWDLqQTtbgN18xa+h
PGpgX6UvAMzbeGC8F8+lQdZrX/qpAS6cE21AoZ9rKZ3OgqfFQik0rkdMZ2/n542k
voZtB8UkoQoocjDPVcNGaQhnBDJH7bMvk18u24VfMMyCV8A7RKULUaVEOjD5wXRO
9qyjZ4tVz3fESbgfXMED8ZBE52e+9dqypFbeQVJ98I+5CPlgqVyo1I4+u52Ol4l/
kh+wnzfb5eeMwIjxmo7cdtwxdbUSKurcLhrmbrVuMWQPKdTac7NSmCDHGSXbWPEc
JI/CZJX5YOaQOH0+igagTJVZDm7ts8YXHwdQ+0LiWTGMPFdh2OcL/PGOLWdP5Qw1
aMYwvy6kmR9dCsMXlYihBdEH6DS0v9iXbbrWLf82PQLqVKJ0pmXtOdvhGWvbkgVD
wAhMDJDmlbDIcrov+W+4UV0rUEDBCloeEn+i+YrUV5ZMn+gaqgG2Iqm3owOWdOB4
8BOhxQNpQdzYm6a2SB5eq9GvE54Nnj8JT7fXbd6tR/zGxg+tTzbwvP8V6OJgYeFd
EvUOZR0V8d5jX76DVurXXowOryX6DVVnF6ymrzJGAO8vm3tSjU7tGU3mik5FOgJ/
QbAD9aLBZhEO5eEYSRZBEbM6WkR2NijZBpBtb7hjdWbL18MSiacmg7dIP9fRLma2
E7Pvb5opZlxHZHk/1jf4rl6uQFjWdLIgeb6YUgsJl7jXN9PMOO6HjYqYx1JsRFpa
QudnGmYskjFhnx2aR8sbFFxw55v+5yDqjTP+8nX7FvwH9DZetYRGItyk8bmvQOeN
krlDbKpf7lMRaVvvhG9ASYVQEbOj9XSFrJ1qHpSdUi0R6dbmTigB7VtNPxlvcaME
hM1WMiVKIhvTzP3CVcH1e5Nqwf+XLPwOofdawIH2oF15jZwig88XFqixK/782m2B
T5RRSvN/gB1YrjdfONKVwcq839bsxZMVS2m/ze2Grt32IXAugRqPHvDWKNhvI3sz
a/q/ljZy8Me8YBDD29YDkDiF2CmMgFD+Qvpdb/M6HqP1FQSbeRjLPZtHFOchp5sF
yapLbS91HIi9tn4TCd6ivkcCaV/IYOzvr6fditgvl+NOoZkshlchGqmIocZCacNp
W/yb+8hcpALfz+10OeFpzedxY7p9qET8gn/KzMft9huA/6mxOTFvy+o6LZvW8nOP
vIoUMXxpnDFEfVWhKVIGb9NlbDOOUSP8oDUXiwNCzWDyF3MXhfNlLxO79dlHPHEI
FMcCJKpEZ7yMIEi35A9n+zp1PJkbFNDS1YplG94r5dW8dOY9/UXttEdF6wfnh9Bd
8kl+NbOJHMN59TLCGcE9E8bYLXXGqsGUHUYdKDOUcIJZMV3KQUk3O4U33sUnAIlj
Br09Ab/zwV3oTfaJoagT+f+Yr5R9mNCg5gagItXCk6W6lKEXSCMCIqyOa9SF7Z42
9KkUFotFRGgigJ1VyEMxCfvOHos+VkmhYrdo0NOzqs8Bbz8ULoQUCCNODk1z3FsI
V78WOUslN5jD/OIL1OQm6OevHHQdsQ2uca2NgxT9U3KHeEeZJScBhapzNRwb8oK6
ryyK96eaX6R2eD8ekTcwTodS9RF9aA7awppa5UXihs2UN9BUuRjlhRn3m5F4bjSg
e6nFWk6rQdzG//sxM1d4R9m915ExUgcOgFNTz+aEofehYXAmB7FI5LU5lHiY2qwD
7juThrlSx9ne8im+jFSa3UK+mV7vD/fz6tocCIQLhOx3AqVAOxqXbRCHlV4pdy8N
2sgqkK0688ZVYb+EPWYemGcFZvPULSFJgloNHKTDR8zc7Q66dKUI8irjgk4k+sIY
9cO8p3H5T84VVTPAw7gGxrjJnMhZPjKI4afXLA56UEjX8z3WYtCAY5B/rFTqBOic
riv79xoEbnjHdyjqKWCKowZpHbZSQLe4JlAqbKNVw9DJ1VMK9dyYzQZCLuD2XvSr
lvtIYkOyv42q94g+2/sG7GO3brEuAOmtwaPpZoidnswytom5MsO06kDJh4EUJj+Y
Ct+9OrWyI+8HrN8Ps3nrEqRKiulxrqEjV+yyIKNdmGEUMIG4pVAewTAh8QQEajb/
0RI+KcM19WFvqC36U1RIS90IwruBSZ29PqIjiQluO8L3AtD+VoHmskIP51tDDtxX
AOomDKX6hmZfpOcQxwE5SGSvipOwkhr7jBHlbuyyo5fv3Nd5LQg3Dc6GKtojkpFo
aUr7NqH6Vp5iiSpEwbl4UzcTIl0sOjm94vGTGe8LjIkkOxR4JxAvcK37/qQ6jJMb
EsWlxiCpevrhSrNY2dG7GpGEAenAx+0EJsljEtOHdZoDlyHVC/YgwX0eL0ivTqq5
LVqgL6TSUzB5eq2HV8hMohQiVAnsedKcVLJfs/9ROP9EKZGqGjVAeWIf0YK1ntZc
OKPNeC42wYaKKb87vHowQsBKedGjqHsQggevyWCeVRYZUpC30IfwD7rbMQWK1Ofl
JLDJ0BbY/Y/ZGeuEOqGclw8n+DiM3ly8Y700SSUvvjvNq+UFxtXD2LHWjeTq8Txh
Hp5H43HjA6khh5EONMiW+ad4jJ9lFs9CTuAEjfcZZzLLR+j9xwOuV+WP+6OFqd++
IOQfdF4aedN0suiQE73401acwgaxazyb1lsHqUuBHoTOusb/l89NU6Qo9QMChWLF
QNl/nXPY7kQta4S9ZfBQ5pYOiZQgHzjQoLpIpBT2hx1FKBNSeKd24/KzBFPXzJtu
TCw0P5XoUwyyPxjBTR9GU/D+tRgQHfdoHEgpw6QPjvZdSJiuar473CjmMq/furmo
t9bm+cCnRqZvmKj3xdkZG9l0ixARbrB/QFQWvTDII+GxR4BMrWsEkv+ku/q9nti1
7Ccmw6AA2ckoDGTjrspfsooQy6A128qRH6vBfqVK2tfx8HslyC46htUV7vm24JAo
RAe1R2JEf1ElHGTqmJKooxCdVyMjqgddZT90qkpztneRuZEQHQQJAgHrhNrJAD9n
KWenXW0GeiCpYc1IFry5+i4x+/zLyjK0Ja3ZRhyQoScZlnCPdS9lW7LM2qW1MDkL
5zbi4K/zcNXpIseZz7c+tqx7sKTkfdPKmfMnvkYXskzGQBFyerMWWqeQg9pTomye
hHpiKK98tsQms1SMW5taZbCynXgfxHvPRUjONdzFvLB7FWNvscNcGd9vZhphzS68
q3qZ7pg/8b2La+z9bbUFmntW8YyN5V/i4cekRTpchthZ4WkTVhvsKs6Mnlp2f4cQ
hinAZHHTZdu4Cu/smRt1A61Y4KFMba3n7i3qwPB3OL7/43ZL55ztR9jU6j8jDGyu
5gYICv+2dcJylu9ab3FkynwiJ5NQND/gL9Ta34zf1f6w1Mjq/qwi3iFIopGQu0rc
W9Sat1KzVWVe+8EuE3OimcBw7cJcilPa9n5J4xQgyoWr7VJXkXdqoEbH5KfCsj+7
mdC94852h63g9sD7Pn1oLrHVgGJbNywsgy1EgB6bjhGhsHJiuf2m0NnBOm+nfg+4
6+oyKwDhf91t40WE1Dcob55pPO+4/KElJ4a7+rKiUO1YCaXn0LV0NYo+DH0OMXLY
QpJz/RCoplsOGMOa9D6MDRlXkQpl45SE+9KBjn3qWjzrvqxBZVTAV1yQUVUNeHVz
FcMMS0N8y2EGeR8zkjsvdorHzSTF1dCuARPQj44MkKYc9HFr/ga1U8NDDL83fJhY
khQh0b1PnADKQJanGff0Z+faa7OBqua0/NlrqZQL4EE4vafbCLDopx81NReEzlw8
T+P2jF2sFBiaYX9kBP9TtCNZ+5QjGRIW6uvfgJ+amIJNa5XZ3lnNeTVnXIWuw6xM
dZ6HgeYE/6EL9OEGYoYPIH2cm5kxlH7RBkxREmNVHzT8W7ITyE3H6nr9U8nD5UmA
jGmBPRocPI+GqhsUo4CG+zPjlK16+N7qXsommVTzVdYqkJSZQ1HFGlLRcwcvajmE
48zde/psCX/umCfbHvXPxOU+D6u+gD8VTYLY7bcVJQNtILP2cpsTimGT+3m5DY9d
aFPjy+83w2kxf9CYWFq+R9kBmflu3RncJ6gjvokvMABeWuSMbg3EX0dWPHfhL5T8
/xwAdew/ekVyiPPyIvLCdrdWv52p18tlIYXHzcQcp741SL9Gcnwe2ouDIhlGdxp7
zQElFA+j7Yc6OOP0bUJjJjM+XfCr9G/7kDE1SIUFo6/pX4V5MREh6uVjx5vc8zPo
M8MUVtmBKrPw6vdmfynDV+pSaaPrvpp3Nu7GaJiEARkJtX1a6nqbk6yNGc92JD5A
6QwMwz7berQ/VhrmcQMjKcy2m8Nu9qf+L7b3OEzVaos3hR9I8k1bSkCXEoVqxi9y
R/470/BsMHGTdyGaAzHI1veP7rqq3+eJ0uCkmy8vBz2ut6xFcT188mVNkZEClKVM
iovQ1ozQoPc4QA4g8AkB6Ue5IzhZtZaUbhh8kKlT3RsaqCep5yDfZtBneOSjVdlu
PWBU5AL+Se526NWSw8JG95rRH2nbRCWLFXUnNcI16z4Dxy14b0K25naaNwaK23qZ
gd3v2g1T5xlSEuVcz+gE0992Z8jVZ1PVS7CYoLVT4krFbxOPEuxok7l8ZWUbOZv3
lSApvHfi3lHvdB0HewTfFaAw1xvGz1mSmL8vcGcocYPMOrNZ1ZrHni7TK7Fpw4JT
aISVDhQrbwP+paQ6Y3z7EPqBh1ejtV3kYQPLx15yq3FDYGOPUqZ0jlaijx+SblBD
9OEy1+jxmebYJBu75EvvpFuZP+ilH4i3jKsnMLICoH9JKNZUxYY48IbFiyRbgVaJ
esF8buk5Din5ZXyAqs2rHiM6VzNXKcx6tZ+qtUM3Pq5kLoajQHzD4qwMRTq3lEYV
Q3ArLn5xfPStF0MbIXo7l0PKh1cXS3e+wCbmBnFxTQstILLQR6kMdwctuRib7S0g
ommpU6ibHfxQ62WIHTGrX79toaZwhqRjs0YWhIO+Pe1hwTsBs4wNzSShonmv42Bj
lKCLdzl2zdixtZfNhE0+5IoI9cDMX9iPmeeh9cGtVuGkvn6heghY9is3qjAtGvaW
m5xh3t46zAvEMInp+KOGBD+T5J4A5si18Cfja0UWPSiMmzTymftFDVBN30F3tQcB
N75nctKhLY9JdkMD+Q9o4ry4BSxapetHYEXtSlO5huuEV+xRqjMyEmA1hHAtCDFd
X3o8OYxafhFu+o3mnR5KVGPBoBUDKT3IJhdIcSwQ6u7Rmp1bqlvyO9hy4FbrTQEb
M5dpTw6licKpRoU4elEXJTKenIk2n1LIEP1bMVHxVuWjUKhW6ce0/DHadYmm2Dhe
MLiKiui/JvPPB5OMUPUsmw+o8MJSluB7+BZdh13LWGPWTlnziKkCXjsahC8HzQHX
sdNehc1rrKtFbXc2A8p+gPyaf3h2FqUcNJFVkxl3BsWcoQoKIZrFU2Bp1sjGhjoi
pNnct+cjfXTkNKXic9SuLXyfq8RW8X5lnZh/f4PDSt4NfMh01kizfOKf2f/AlRa6
zduoiOw0gec/AXFnaQyIaS2yGHxH8kGEEoXLr9YA7OXqMgeYX5d5bULDcg7Ss6Fp
X2Rz4Nf/Icb9V01L4dTgelwNKgKiczx9ZFZh4o6h3EoxhNfTzNgHKnLeyP7E3f1f
HM6Z8+0vMZlQR8jHlJw8pYSvSyXYuTm3ogq5F28QC1sMJuz9kDNwHy5JCkezxrmi
VMDxrV44R7Ydz3F6Z85Ri7+DO4zQaX528p1652tyCyQtCrkk8YRHZqkDDeVB5rmv
9DG7gLA23DCDBz6jtMmO1noct6bfUxMm3l/q/wpeQvJBVE8g2fsSHHrHfTV7fLeG
WBmrCxw5OGmKgDoT5KcGTOMjr4nAz795LwkTiX/9BTQ4FCZ8adKv5YFGOU+USpNe
H96kpUnRdqOtlATnHQY4lFcnAcF8KbWdeNi3NBwFyrGyjQe8e/hl8Y9gTQS15Q69
82PItpalLO4nNOBCp5rVzVMmCEoeYluqf0vV08UnpOYQ9jjDYuFtPVX5wUa1Nct+
doqzhTgmg4CjsEbDe9jzeSpcaZOwC/zGpk7u1655trRc9TXT//kPxVlEm5bSlisP
haO9+xlf5aWKH6fjVBQKQf4QtB+5ZjFNzdbhYiH2GDfAzwXBoIepLC7hw9aeYAHA
foi4jBKy+gaGkqpqCsVrXChI2/hOlqtLEm73cvTGxSgR3O67cRQqEjpQ6nnTgznb
Z3RcZYwbcciOf1gZHn/l73J+AZpirCnY0lcDOY5/7jTJ1Z2a3PlJwHTh1B/7z7if
TnEVOm20yDgxpzpuvFaTlcZpBQKB/YvBFR97YBKvfoZ0/wTJpbISibYW+u8AN3Zl
kmiHCs2Pq0VK2WmaZ6RP0oZsLYx1DvkS9ZhiTCh3/Jrqzsy/JdMXFYIfMW7f5wrb
cZvxacgpPlK14W3k3MyNcPX2iivN228J0kNJxOhBjmapUj51GDiPA/iyX/6FsoZd
/Qgv/DHYDoKGy2xrPe/+Hte0iUYNZWwkjdE0BSKFRXeb9zNbFjHLVgtUOqVNoQPp
kwuim1FGLs9iJw5/3+UXfVvX7hVC/HM/smH/8a80oW2HkV6uxbCPR2M/KMbY6kun
orMwKX4SX3iBYq739cLpOfivDh3YXRZXNxsa4tW8aIRMILqjN3pXvaN0n4h1xy1Q
MBnAMNwMhtl1QBgMTbwo9esvW0TxZArJWdgcBGeTXoohSpLfITdbRYqsLACWUHL0
cx2UaHRqq+D+si4iBCT3bKLO0Nf0uHkSDkM6+di6VD01us1s3GWqx9LUvs5mDNt4
SYv9z+SZmK2TN5bLyzfMOYwip/HOaZe1uDBrI896xEkU69WfWABx7v6pFQV3ZQLo
mEIPFtpZZEQ5qc2553GH/tE1ikNcbGijfTRxyCG3t3tnSbhLWp+UWnuJgsOh1Y4M
RBB72mtCjFvV21rq7aHzVKT0NqA02b5d4Inm0e7FBMJs6oz2OYQo7tWdWA51pDNM
hLt6vOSRhTE/R2hdG9bgm1JscwM0dl+ZC6eWEb+EUyK7ci+AwiuFGPaItbQ1q1K0
15fZuEh81rSTG88g0XM+NgxN5n33KoTMkw7/A13gpPgiiQuLek11Zr3mLxDwU3mR
R+Fa3PJ9toW9Yjt+tOmVeW9Gs51mxkGpDPxIuR3DIeECWP4Nm6ZehL5MqyPRASe0
p8EdDcK+Jk3sz7JAaskkVIfpXUd8gDCpUVGBarOBiQcbBCdhsuwZQWHXJV3vsuSK
qm1RNKlcKn5yPPuqzkZjlO3Pr/vHYBMCZ8XuyLaw4YhA0SW71Sig/zUDNWy91Zd5
5mEWVnpCcj+wVg5REFkicFBitz22ZWjCRehlukjPlmXvTWYtRdiarEZC3VQv5N1J
MUQOL1M3ImUT0FRA/rbwIyedlQHpvR5cxkb/vZ0X5zXiPGL6+jj1QGwKwLfIP8R7
rD75uVPrBvkjJaM8hvWmD8OyG8Wr33m+GWQlpb3mjACo+yQ9wUBJXkQT/BlAkYRv
QHYsPa4dNOPnQZnMLevRSNjNGsbjGv+VMmLiww5gmGlKHZTXW9atQWouLfPXG/j5
FxwzywOe6B5EnYErfRZi7zCO+DcOqpf+V7fZwcjwSQsIR+hYOZk9UiR/znOBSL/E
KaifMAOB7cpPY8e6F2kETTCiqpNeM+mtgvg/E94dBRsRB8GbFAkIA3X8BdK4x3wk
YDJNiGhfyaO3V95tIUUNsJUL+6FxMcavG0iV+pj5Q4rxhL4is5Y0z9aXq+xqCmh7
AXxDxyL/IlZjl8fcOZMcIPSN+COdCCeos+TNdntr3cnWnLyPCi3GhpSpkKQguurh
+OL8JKT/1wbKYJR3K0498X916qFen5JTqkO3do9Y7XVcr08C5Wjz2ka1qyPJTEc7
KBfFR32iQ+zAclDZPucjfTRaMn/aLUO7nKArFC9uieIrmt1n6jCYCymLU/irqZ/V
yotDBI8VIsRmnoP254dzIExHMfXWy+Qrdb3sZzb3/lc4jszBs3HYJqoElQ6NimuE
HlMYtlZgjK4Qp/Crc00IpwSOGEVD/JTmVpbv5DLqNfIJOmYgegIrejo4NS85Me88
eBnjz9Qc0BaodZEdVm4OHD3H0XNEK5Xq3FHk3vhRRO8lzrXU7bZLBu/KxEK6i0IE
ekPHv4fEjQaW+N/5Lqq4+FdkC5yF0CoMAGAguIJENYfonBp6NU7+Mlo+0Wz0EtIi
QEb0DQS2Gtfg3wYeZFgiGuBOtcMRwQMeRECeGyPJ9apty9eXRh0IiHuua5iz/fKG
G726JiQsEWxV6KLdniZ41zjW7Ne5fmmu733dcTLM58oJPDbX9+Wld+jBDe21YJ8w
I/OAT43ji2+cPYjEL2bQFAj5zUEi+HpC/6x2iBWfVhOyQ/Mi4toAj/eV8RSDsaQa
3fdz4ghTTyJ2rihOHP+k1MCLo4Wa8c3hOPqnTTRvORGgj9GOeuzVVO4WfobrTOGE
kdSF2WBO42sjYl3cgqVEsAUkrbyGzPUApxhg7ZRzY2dAI6WC9KkJ9GVqF/AaGAHV
VaJAmWvNQZqkHOSnkbhikn760HbnPF+e/6Q3/LyOnhaJeLEf+JjXRhbtKa7Szfo4
Zlct7naBpoBzI6VaEdc31/NY0Ij/QPGJaeX9dSqkwiGPJ28SuAJ+YmRVjargvdZK
ec4Kc3JOJyfP4fA9kkh6ljfcBgfGH295CiLuaTv7uZJayqAb84zNwNVgafbsLhqr
HbFjXoYTc9b0cMPKOjhI8xbtcdhv6+DQ4MdkdnV8B5lUYRXV7E0Z7hqzfhaNaDQR
6/ljyZIPaV5OKYI6Hur2PNBRHkFWTzUDJVzU26IAP2Dicj/zr0MWxBbWtpFoHEis
Bz90rUomAgkB1Nllyf/0G8SoY1nUpM8tfZMrqe4H0u5RPoc4lb2E+f25w/+QXBy/
gf6hEW1izZ9rgeD0cyVIY1wl+ze7Pfbp+ia2+J15LejdfuMwzbdhgUNa/R3N/fxY
tJHIdXdlLKqUkMx905t7vXXjZ4GkWAiNW9bXrRVj8+mq1Rz8Zirk8EO3V7o6zVAm
8/cnIOWS9L+iLErpvNRKg3jSYL3RM76eb8zCLiHkMSY1w1D9zNfFJk+/b7G92kXQ
qf81FtkTWr/lPPR+VOmRicgx3pMgP2xgVzcOY9wj6XYkOIKqZ8LtFDGSNJUOBJSr
CySGuM0JLlaqrgXPv0JaHD5xuUfFYDTHQa3QkyY/8EowWN1TmRkmI7JHj0bu0vOq
tbhUiDQg3N0XD158AjOQZ84oplaqtSom9OfNtU80UkERbsfSXIwYAps2nC3/RStW
xW/oSH189MqDYH3+wr56BhqsWLVzG/DgBRVUry/j1CMDwV/TyuikTB3ixZQbZsnL
3u8/K/2v7qeAM3vrep6OHJ6iRS886zWlI9oUbNeTO26ZkXwK+ydGqMggAiYxZzYR
Lxx+/9ytVsbd2Mor++Mo32DtCK1bNyX/3D+hwpDCiKsOtYEeAerwVB3dB97liOIF
g7/GcQPGOX7PHMojEMYoVwoOTeW1HmSivoRnNNl5xN2F2nR6dSal8g9fN62xFRSt
zkNjoXzZyRs85Wa7iwwCT24Hgy2/rXAGm0PSVAK+wH5G2otN4ED9pS0fxU9CzkI5
8ItJY7Y6wxsHa/L6UiENAHw2RenoE6htyGS6oc39PNbyNz9f+RfTdRN5Vq7oZiSM
p9l36yiG9A6F/L1miPkTz03wqi06UKa/RrrI2aAlB0UO+odTJSsX7DVVE11pc0rI
l4SmWCUq9EXEjHdMVrd1FPJKZNYBMuyDpSj5usUB0i7JxSw6JvMT7v0nMFM3hTvx
ktM/ZevkKkAsWGniNnUdxy0ZrDOw0EY5CjMKVkTIquSENdjgwmzQc9RiIu6DjkXi
Xu5cgYYvWOQjKoib9v6CkqiCkfVZUpEWOroHVY1ovG0lRInnra+vzidujXw9GCrm
TL4cNdS6kgbAOuxobi+CSD6o8i+iBu0UxyUuOTdxFAyT6CqSiRqVUHaieOFQ0KKa
AOC+4Sb8JG9kkTayNcOZrPsWRH+ZPGjYVbhqD9viHuWzQJeVzXgaN+VOCsO8kddL
5pluk5M0MVjffLn2jEQmTW3BfqvECpi3c8LbK6PXMsZuLM20fteTNOeAu9Ha8eFM
y+pXzlx9FaU4Bdof/tLAVHmqW5r34PBeQdcn4Wv84lD42GsqDYoyt8WhPwrmwHF0
Wpj/J4MKWbo//NbmCI6pYau39ltATs5UeoywGwErvKANKmBSeHFx8C9qknxdZH8t
gJ2naeShLPR24v/Q3+bX7nAi9FbamNBKxj968s9CeGLsO2KMSv8ZWixZJ4ZhPi57
tRGTUWvf7gSg3f0w8BDRz7/8TVec1hsuhou4NYWbTXguYb+SrX+r5IZEfVUDMxLB
FQPDRzNRMJrTq+rfxMdsmSsYkRtSCbZGqHqqxI2kNZygTD7lVpXFs7aKizXsB7Lu
IlFamGSClmDfofqNsRSam0Hcdc38rNpGZgKsnvbjC7+yPjT5RdGhfdbFiSQvh/fD
n6+4A9j379gPyqGFDSvYoNqf3vjbIQgsUVjXWmJdCq0kFA4k90uoNVdUt+qebZkF
4/FPPJQtM9b5iKnoxZhFicLRypWlbzYyte9qlX2l02qtmkt3OSlCYOdsshnoeBPp
Smo0Ok4X+HcNUBEob70avZqGwgw3g6tyTp9tINo9kkZgh/Xm8QWHn8inny6B+KU1
ZixNKJFolt4/7CK8nxENZOFtRkFC7fQkRWqMgLE/lRSmGQ5HP4ulpcxxZ81rVqRK
ZX88nPY4bLfZJwhRcJjiVRldFFWHb8FIbO6+ZI0KFZfNJRF1hfVQt/NlNEBQde5B
G+n5VV1iJrZ18ZraiUzPrZgFTGASrMBKAgLAtLYTsFI490i8vM4cjYz6YUZAYwWt
ICs+eOzlfoc3r1Kk1cbqTgo4QKnmGQyoO0/xBdP2ec0jlXbzm/YtSUPovJocN5g4
R1UgOX2/8zzwL1lbv1NRmQapunNmC/yXXWm7Oz/M/YSITtkulHMV5MCMEjixUfyG
qLMDY9veD8vsUb7C75mMCAHrxHdD5AcltIni29HenScCfbrZnOtGGS2N98Gek58E
GX7z8Sp8JYnLG+OILZSZzSQjFs6oogzlgth4Kfpu3DfD3l53O7Xue7w4uqnYnWN7
AtHZjOsVui9Xco29QyZISdMUWbehEYtN/S/2zCRB2IiYDdnXQCobC+GdzzcEusnq
j0WKRxaDn2Il3aW3YRH4h36oiGYnlmN0NCMU4xVMfdkwI+wnAoqMnqNojy9uR9MX
7l8tFVMyA2bqogzPkc3bJHezB4rcah2TJt+LeWB8SvY2zA/zj0tRh2UXhGcR5TKR
TWoG3A+b1Fc70p0G8Pq5mdfCC5EW6KK+7O/maspfrZoL7IS44x2nXQsP4PtBbvjB
Ob6fXlkfjp2/bU4JYHmenNjPEBO+XcIQzsA32U1tNKnH9lR+KSvt6uLYcYf5MOWO
EUSMYfKGhV/lVPvlkbwnwIrMDAUjsEQOt5RwN5mVkUcJei+/z6GmtUbYwFRD4caA
Il++eehd3Ud7JQbJysnyPI7sM2qXWgzTlfn9JG0cFrFFeu5ZN5BD+9TcF0iLikwL
rJ6kQRocgtz3p/nsNnrt1b4/DytvFURxtfwBTu1KjJmylA/JsdzNBoQhYAq8G+5I
QNG0sZfXs0F/6V2D+yZivVCx2oiaNB2QfJaEXctglpqTRvVwqyj8cVs7U5869zun
4TTjKrOpN2edqXU2AsV5C1EKhUq5Zi9Ta5NyK1ORP8VtFhhh0Ar0HqhqPoxmzB/Y
/kGlwyuiOvTK3+a+ufYs0KJpmjmvLWrGUMBbaZiIwED0L3XbF1vKsUy9p3yyF+2U
C6dR/EUxHiMBckoqsd0TsUpG9FBm9im7PxJVJ+u/GlMZExbyzmBUkgTVbO2cjNj1
YkDh3NSE2WEsIDAXwaTpy+/NR0FQ2uRu8qrVjF+UBjKU+9nGS8Dbf0l8DQdLMYOZ
AKTlY1WNHZf+JtiIqxUv3HGIeQY5K9VXM3pjG6hfZtZMyKXPoE06gFshrx5OpG5q
ph7LGFu2hGp6U+LEv/gQFRFRBGDn+eMaamrIsk0i3s7oPiChzB9n47oKOoBJpnH2
kM8K+S0oeRPYr1WjVdUSejnLqnuBDMj2UQU0E5NitPpDgcSxGVYpULG1j6G8ufGC
jYgsBCBVgTP5QMJABKJQOAE9Dr+nS9XIt/jeexKLINEmctCRK0LQ0jxEMJsZCYXP
iiQl9b3fVXVRjanb9YZ5mLcYuB7GALW9M/Bd+M8Rh3CP/WFRK1IBYZUMlnu5PwXR
seTpBefW7iqj5OqyaM1EASK3nY2pbGrb8UwbKXf1Bbw9tYmAmr139rgfQe1TcONU
o9iVh0kQwdHpO50Brp/P8TvFRLr2OAJxjI9WT0dVn/apDvTxhpBa2+QF9KDGwOI9
Q9sn7z5MQKPYVPSIj076WBZtr+053IdqZGLjGnh6hpLUodIJyZshT33qlLvljiwZ
SCOx/G+sDaOCbloaw0cyDW5K6wGMpwSNOEO0PZrdWlY1zCNtwOcQoSTRkZkAe2sQ
2/crcIwm6UpOwxdMgiGvkXdDbCugRJNQ3jHiEYdcYrpQ6eOzSdo/FnD+sh42rQLi
y1jKSTovHQJve9GIQhuUJ/zj91YZDG29F56Ksmes79+r7m2mRGDuD19Du1FxdO3d
XZOC4XFN+xpt9WDDYah+Z267UPVXWylBGMhtiGMPe/u9h/BhH2H3QJfoE6cHuXQu
hxJ86X0JnZoMTUkgJhI1trhqROYarUsPh2JrkZJNPzDhs4005fhslAC7dQpdRe66
oK/T6jEl1IrmIA+sKw1r96jAOWfxBCRozY11GNPv4/QmLw7fgwuLRzDR5/lC2uFh
kDfTL/7rfiWBnp/0NlZYCqblurseP8vAFKSg5CwWuDJBlBon1+YbMUt3wLOmGo3a
8xwWicuWu1BxdOIq/thVV8qnujUjUlu7EeZUUa/I5u405KKwcU0W3BO8gzxdk+tR
DnPCinDd/SxL/a2FLBBqkIgdJ9xYxFcnxHu8SDtB0Gi7XcYP9r/Y/ng+Qq2vnZSU
47EIFXkHMyLDvvLF2eVReA3JNmeooapTAkSNGi/mohRsZOIJgnCLRKFJK0iAYXnG
5zFUMfVByE30asAq9n99YXysH08+s0obSQHxIRXxiU15FzQe7xV/nxYe9FBwCG87
jkXbE28K2Sr6aH4HrXyOieZO9Ckw/mc79qjcQHMSXyAb7wJsTvj4LL2KnAUoPioT
etCVemQhY2BpuvI/9Kl4ivzeQyhgqxxX/ZWSm3a+Cqqu9g7bpxwXf4sCmHhmjtls
pIfRjHHaYtCxAmBrl4adk9j8rpKLC+im95OPqhA4zP80gWI7jDbjQG/EiSMRFH1k
aDojMmHFOsReFY9QaP4gWwSOevG9+oy26lQoHsYhMt3PPDHmWrf+MRiV4J97xB7j
akh0qxq0wz7RnSkoWoSDkqMibP5Y6loVYeBKGd0GRng/E/1rFKXjdiX3EnqE/2/v
0ccI0DYP0x4WYrfWP/o4SxVkHqH/7gHCibpXRcb+Aj3isRIGaKDvhsGFeA9pgftn
7XB3zCPM+fAhJ3E4/VO4jAQL1G2HKNj3R1bNFuu8T8otX7SnAJq/9/+2/q6+t90K
wZHp150HVFbwMeAkgpuWl8BQXWhzP3h+GEk+/Y2riHPzZmlP4Pn1hUWgjJ5Z1agL
vjeL7+afGBfX+38Yn0D/maTv7VBrV4Ofn4HAk8Mfk4HZwNtppdBpltFZjF2PX71c
n8+qK/1/MMJPx+yLSdnB6KF+Q3pMdcoZtRyxTmgpiV/iRiLs/wr0AxoPDJvaE9J4
y1AlSoMjD+zqjLXBLagOYTKZfPodHiaIsSt1rMur640ZMmznJQDjHe3sVIvH9ren
K5oDPOp0l0ERiO9S6/PG83Ev6KVpLsPr14MWQJNAiKOKYNuIRDHcdwL1qTx8s802
JZblF2xTb4IrHfQBoN8IosyO7hFyyR04oKUCkEfQnZ13bpzwsJVvL28VT3pNX+Qo
FltAhlcmOrZXLN/QwO5sNxWQ3OiQF7Fz3cUS+x0Ul54vZooBK/2WECn9dD99lRZJ
/uaF6MTcnFDPX/kbkS9hLVf8oD17D3nBC6H/V5mfrHyU0BfPcGBG9khv2U8ubNdS
osYnRO0HPrbBoX0qSFmom97o5UnQCzL7xK39YLpFzqMuYtSqYOjQF43Z7KSZHOcz
kSFxoh5dJB8D9bdBOyUt3gFsJKHQdGrpdupw56kshGhiX2AmCiehNkgPTPK4dO5t
U+xV10Y69LxClsrVY3Ns3hqowalmcZ1grTJoOpt/73hxz6MrQZF681WiWYj5a7qn
EYNyshaX8MivueQEKGPh1mlN2XavSmvhZ21GgiwIy13an7UW8WWA9FkRzaXyzqLo
Zu2bi9EPakkQQviaFzeZAtWXwEsKnJIBGMnYs7ppOoLtaNHPsW8q6dnS1eN4jRCq
Hk0BYTJ4FbohO20Ej8FAVhtkQPWZniyd0DswzbhsXbEj4ANOONO5S6E6Ao7vedLk
3RPlIdLF4V2Dw8sQdCgZPGycCj1ZibQtF6tHOm8jYdkXi72rN6bRyC4tcn1v2zWU
JOpwngrhsA03xi2lkJI918HZjmMuyf7YQYtYN+F/F0lmOgTZKisX7Uy/dqAnFAvS
yXyhBJiI1DB7a1ev7SbFiWXzjNuXXuZLmuYcDg7CLO8jItO9Rz2WC7q4kBOoC0W8
OBigGLdrdPbhT1g1o08OqV4/Mm1tV6QaOXdNnZD2tiPuoEsQ4/GAhCi0iNqgsAbd
Snea9R8nVsz1Jl7vRnesLVr3TvBDvrstEeIYJKeUg5qspXxBMICLGFxRMbnykX1C
/WUCnGapj1hX8T7qk9BgYh7HOowg/lnQrKemjY1XIC9jGdOaLFWtJD50hMiWgu/I
hemAswu1J12JHkPUOExTkQMqxrGN4q30X8BWYqSUv8Pw5c9NLXia0vGrHjE01Sn9
ZckFiMWMkI0ijUTQM/wO0stom+YOebSUvZOJv4o4KTVZNfSuN1aKv5x70kdNK3JX
vWzKgv1LojQKfnwDbcKVkRWJItqMQ+Muvtn86R2o5339I+zyVm2r0W+TQXz21e32
gfRpyeG5QKaijRfo+gHQireoFl2TiYGoDXw3/ocu3T1IVNKFQwZtNR2LjwJmMp1Q
t0QjnSd3ylrLLmtEYGMPTbg9nh0Q3treJwDTsi3e92jf+EptmgP07F9xKE4KfVLr
8hG6Mlgl8H7PZEdnACb6cUPE9/+O7j5F77CioAcqpF6MK5WmCDEEDedw5mcT+9wk
h4lQykYyGOKp9XZ0kVEh8KdIHDUWDHUKaEJOMbaoSKRSeJiG6AHgeXZHTC1tffx1
BVlz30kySPIM14recFEhn2DFqZljk9tL2UJYP0ZWWGQgJhLgrIyUUkbrGwmKpqgA
AkFlbkqhmoG0QGU1Xto9HKDu1atoakTjag0+UXi7b4SFYQK1EZR9140akfz3n5fD
p4ExAsZ9VTvSW1NL2p6EghroqZWKL1W+E1nCfNla1BLn1MaRPEOcGMQECm9gJ0am
hohV6KkK0l+BEsiy/oY9swf1Fnwx/GXM8oDoJViPCjD5jLMClVYAKyjS8eZ59CK2
Q5q+4R4/bMKPNTgnIfcpPYJvKx43mwwt7ctJqnnkXQ0HAfMgisdl54JAugNy3+L9
50rgHdyY1/GMvyCRrRu0deZicbpmJuSj1UgjRs/0nz9DAbkTWBV1m2CtSLubVRPS
CA+MQwzHOLvLNnu3wRzYzU8kIzDKGEmYnat7S+2pxdy7UmG8iBKIUTAvR2KrtaW/
Opq0MbokrgyGLVVg6rvrfwYjglbWeLEL5uWu/uFt1AbC60CuI3ktaBnHYQq04bVD
DyTzdewgyttnMqs8j1a25/JLJ6FvmrZjxWRppI0PlaBGeaR5MBfkuHn+xAT1a6Kx
jCUxDIwUC3oDknuvzoagusin+XxG8XRKMPzYqwu0bkFZOW4Tm6BDL+aJiIMCXIJF
PR4BBDwHYZdVHql7Dpuo+ucje3q7PtX1WmS6P2jKcf0rCVYGTXYG+p4gAz5K+Vkc
jqEmVkVpK2iyhSLorD0PRJKVUdKfR0wt36AapoVZMDuxBr3gj+hkQOPWst+/WNHA
/Zd0IIgIECJiGkfaSlU8fhwvm+XHlf/Y2/CgKW8t8XKT3mDUmDoitCSNNlUXDt6B
+tXJQwf2cVaa6yjVj1dtDpbLWTnuugs7Ii20C+nhnQPiIL/hPcmjEcftYvr76OJE
4JzQXN5Ifa18II8UgyYUUICfBOcEeiMJtOxkHgeoSIB+9piPJfVTmC/43VYVLwjo
0Hl0f6iH3mEFovlnfgEFTvglb7GXAn4DYKAi46cG5P2rYGabysLw0/DTstjk94lc
/vrwo5V0x6xVJvDVF+0T3xDfezymoFna8MIlKtdallN+8/kl3TPqvFvMtzcsjX2s
qE9396z1ylTLOINdUVpDua1TGBQgcNpdMrS78XqgyDbLPKH71xBrD91zeunrTTHj
0kHbfBLzGNef8WoHmtJ8UgeZxgeHazacC+AncuhguRKiU8DwPuHEduvcE11gBQSK
IQLiqFM07g2L2gLlGWMW4blCJUkv+Dnjje63K9sakO600JVqnhJABHUH8/HjX6Ki
YrCUx3TxtQhR4BBAr8AwowV0KIGLsTBtyxaFDKdmYA51R9MdN4HPrQvc8i9/yblC
5Qzvsb1mRUrvMGP08bbAgO0jxdT7aFWwb6kriO38e5Vb8i0Dddi/wCcxS6cgqCnP
e5MV9FleO6JIq+p0TqMCrSwce6aFdBbHwLGjbujV9Wo6b3UskYrlBf/7QGdB8r7m
13PBh7r5mx4EZhz1vNqgEwntKvgbPNg7Ic54EQFX4oLW4BYF3jg/sSpKEtAENP8Q
IwLV62kjFOSZ3EmJeQMfy7CA9GdOeDj2RB6HvNZZDePImjttVuq9v7SzGRUjbHYP
j9x9+DkFf9VyXhtZPsGrRf4lB9rEyCVzdaDmrFj/G7dd6JkL9mRK8RINbHI5rGVV
HAKWEbeXAvPqHuIRZxu5yApAtcsux72IZvhDeq4QpL2FHCyjJehKTXTDlUoEc/Xh
cPUxrJqyqonA3tHknx35un7TPT+Ec+bq5/YyugiNJuSK3tG4trFmqIIlwLpWopDP
PhmmR3EIKTsg+083BsclfAGKt7nse6zX4ejzGm5RjHmXFZiPDpe3jfBWfCoGOASc
opsHFeQ0HGDEOi6Z4IyT8YrWI5qrIkCEtWrhf+MUOcOeGE7GjYMuQWhDZwOf5Wpg
w/CwJ+2xGIuoaB2L73h/8KPlhspyiMBPB6VCzG1nBdtWxWuFzYeX+3V72ktQ7byo
BHI8l1asrrPOPsIWZgJ6wY2Q7aOLVuCri2LO5yAc7gcD9PCAg5vmShPDpqy1VHi/
pz0hHjiihjkCI4Kfj4TFxAr0LjLWI/a4b034nqM6G1kjt3+Tc+sKrO8zDanFNxgE
+0AEUKF9qfaoxFyUMWH4DyMlBysn4zJ+twrlkGKcj6uxsPgBDiD5GB7h0PiH48zV
g7Fx3VeBZtlpPNUsIa0vsPZiOw2eIcRJQu+UOf1AqqtJBdxyjARvXQ8tc0eG/rI7
TyeAlHJmxF0fg8VsmfGLXKyNJYdo2alL7dUbGcvEI8b5dk+xskCnkbM67HB89ahb
AyPdAQcvhySQAZXHfGoaVZH9dYORg3SkhAb3vMX/1PwH5cwHd0vo9+NiARnx3gVI
I4l/PabmkjDWlqIgQxpna+6O5m7YNciyUZ7O8QYF0a3RSVfWuzafZc91C1WTtlFX
2gKLer5ZvLYG0mnFaIDNUSywv52UegOEeOB70gVB6HySLFLYSTnDMiDOa8ZzBcoZ
MgaY1eMYAGy8hfN+3fMRi3Si8DqKMjBy9xnPyny9hjhlg9pHHH7xxj7vgVZi1ugB
HrRK3QVatcT+d7BrBkBvqhZtLUaYXMHpl1YSGyvLPA3Y22/WEX0//plbuzNA9ihE
PUP9wMMe197jO8OSbqeiJNmqK2emV1O/zN0siTt+b67MnJrrUApb2Hg96AH9ylz6
g+yLnbX/seUJaYFQvBb3I8YKzmSV7OgM4DqAihcGZ5HCb2iBd4mYQ0i6kdkVgsEE
o4STmfv59jvDJfx8vFO/Df+ZPzq/P43LQYQt8Jtwa2NBLvLdUip9cf/MGEzHh13Y
gFrORfPz6bH0mLpM19auyY3tPMXyAJhXRBrYuWFqXbh8xwbsKsV5IWr6C9Lh83qR
ElyZSNMKhPgDkLDc9wcnzCL24GaU3yPfltdT4ATz9SzsgkJ5z6I9s/0EKTVb70uK
CW6KzJxxuq/d5vyjUjmEJLxPIzU7KpOfRl6lBToge8ubSmywVMyXpjnVW/bosbyj
4gz9WD1ETDuL+Kint2mXr2Yr/N2nptLmQOrK6pMa/4HxdrhuLHVW/3FV/PibTHGx
Bfuy/JAJ1dxGg5FTMIbS+9yWQ8yCAwmJyk1BpfOjkRxh4BZQpB4sxAapWnNX+XrD
v5Y7qpj2YQZL3G60ZsUmuZHmd0Quv0Ijjy8Qw8l8PNxkHjKxm77/AB4pt7/D3ZAm
9Qd4h/DVUhSqNMIOmT3pE/s2Fo0N5jlXlwW5CeIAcyJ5esVBV1zjsMg3Bc3Jf7mQ
ZHwzopjOlxpAwPqKzNtMb4hJMwyphqD+YDvXYqysMEo1NxJpg/G/8vPTfmJVBFn0
gktIKo7H+kYw0R8+WfBtdz6C+vhUCqxgvfnwGgM11gUoVF7yZ4jJ6k2Q5aHKsAhv
Tc42iNPFhc8s2nYTRwQNQA1ar/gPi4x4G+RizSEy5bhIXgoJBZgmozlWUTB/xXPA
sL2OxnFxWcxZAXNkKPPKS3RArLSArx5K9PEYWAaj6hiTSAdsvz9enaUVlpmYHMWK
VbESEoFYK3UVnI5iEh6CtqUp9dDrUNAd9nBJOaXpXK/V9YO6/T+SeGJEstTvbfne
CXqImt64KnoQEovwjxX/bDIvTlpXwlBIeVI2qTSugs3XHSnuQKczoQQa/QVa0eY0
h2JoMixwjW7ia4xNFRgDvrl6tVeE4rmxkOPc5Wl8gEBrYE9pqPLByq/BurkgAio0
o36b3rUjzGTofQpZpofXVWSx7wud2UgloBJZIcH9q88NR5dtFKFtcj2zg05pBImm
luWrYjt6Ain/qP+GpzEAojg2TrJpBbBRJENrKr7cY7cE0Cario2PJR/d8efU9hWw
RVKnhzdRDkHKXdYz6lPD6KAUoYK+7QqGX63NO7MtHK7c1GVfoiTVG1l96Ljfwodh
F8Zr02efXCZF24SGG4AZ+ySG63sgrKFIENZS4zFnRLvwnnLFwWeG7gcULWLROnyG
tKHgYXDbubJNhBlfPfgUOgmO7nvqj3lv3X+c+6l5Ykgi65ylfwJtsw4Pj/JTroB8
0qmttuB/06H4wVVPGX9jlQeUt+ta78PjqW3Uo2fatGiD5/V/J0wrDGQEMWiBx14W
tKqfscbD8M6m7hLCTiLA79TgH0q0Eoo+kWltdWPNqbUEin+84VoBryLj2KmrV8xX
fF7MxOtvFyblGIVByZwrUAQeBiDstFgaP36nP+9VtbnGkgEtmKVxZx440jKM4COJ
AYDMx86qym+shAHXkaH/RfzaH/EU8iYsrNl5k48wSPFqBF5TJISKKZP2kVLDxnSY
vHXDf7R4ADWXPkWrK8LBxKYtwtEHRHP+cVbWI2a1zq7zbU6f+rlIKHUdJyz0ZWQC
QawuIzltR+QP2YrPSlJGqKtOQdEr3v6ulDL5LmnEHK8bb00ClswTMLe6FeYAgi1L
0KP1kM5qatzqNdSWGth5xbTJ7VDNqWZRma2GpSb9E14U0bDVP1kYc6gre3LDnHtW
7Bba63ht7Jq/OXtVcCcE6FGszEyhoLr0AyWbUJT27gUTdHp7LElAH4rccOpU1ZRx
IQI39+qbkwCCG6yhAyr+WACy3giGuN7opbIKuTA5GoPTh2l08GfJc9xcExmHwTN5
TIAKnU70gdMBlBVGDhJaIfVi7B1U30c6Jv+y6wzCP9XYuBXn1dD/pKzWgSZQOJKB
siEtFp9fw0ssAoJwChMZA+mGooEsYKc2kfaTT3Yf7P32MSf2NBXAAXZ/ITM4VYRS
LPcxWHrnTjFE0GUcuzlKkTrJyakTxbvlc2l6iNtqNUeVmvDhRX2NbmQANHuBrtF0
v7OkNcKSjGo8CZm7ExCWDZik9HwL5XU772i6z0fciw62NCqBEdAxCDYw30zqByUX
9hrrAdYdjTwkMJQlMNlQzCnDOp+L+tlx3+gLXuYFJQIwScl2jZTnAyYwJdj6AUfi
Yk+An4aX+WGAskCMcip6L+fzOFxrqWwYQ4dlAzxsOhorDe/Sz9c1T39kruU9fOA8
J4WmYU3tkQ4BgTAZudePl7YDjxhHXAyppT8Mn5J0hNZ60e7C/LNGoKcn+th3+cx5
Ie0vrhrwjjVjUqhLaZjBqSsQEu/ozXczA+Bf+7KTWic4a+crjGBWhbmj5dsAKg4m
iT0xy8NzOH/1sCk/26OwohrgSvXUwuJ0uYvgVShgFco5yX8T9itHqOzXOAc3xw2H
gg91IaGyTwerbTVWMiBsS3DpyVkJUBk8YHFD/l6HIXrfEAk45Ex+kBXWdr01hiFE
vkco5GfUCW0oMfB4rL+qfSV4JyY60R56/mTQ+7QrnyUd1SrtkRdu3gPULGR7UBTG
NN2irkpA45nwM9US0lc0wyRsaAz4QlhzpbUoMxRI067IvrbXJclmudlUbZvqTMpD
fnR+VYdQwlKZA5GV2v9eEnyq9o9Is2Xy4Ura8TV//Xh+lPI/DUAE5niUrvITcHCu
rYJLVX8/cdF2epILLkF7B5qsBSQWT7V6xnT314GjyKibhNHblE/8CFIU9r0Rc0mT
OyRbcyvNuoFdITmKT9vYgmv5GQUN8XZPg0J7R2p+3hxVt5csQ/wTfsF829WdWQO7
pii99ZBhvhjrmk3Y6sJe3dUEBo1duoJi9+Gr4NMSkBHBMTIp49h1bdtk6iu/XGCF
HS/mciU9DS2a1xDJfY5aIPQsqXJRA/YKok/oofr9iVpNvjCB2pl8VTG8MHahy/FX
UMGHOD9pzPasJI0xumhPhCWtbDXSjw8HVCVY5HlQ/S7Zv+TwQNsHs1za0U9kKKh8
RZs5qgibmRa2I1FvjJuQkd+SgPi1Na/09VzLhaNydVNC8/chnK/Z/7EHWwhLFA58
wSeQbIdex42JlLfBgrfBI4RwdndKGvvwwHfCH4E86bQ/pwTnGa9s0nPY/oyOv1rJ
ouyaeUfN+vytl3+nCyWlhGHJMbzVqdBJ3i2iMP+PXitpYDnVQvNV0qEh653p3Kl1
Vq0qFsSR+FLOvd4HmijUx0jT4WlJcIUxDt0jrv/UCSYEVgwVRVB/BSAqNQER+Sgz
Ede/b8wDJx655+IK/EVFzDtyCVYt1Hhx3Q3URGTonaR+D5FFHstKbbi8bgOm/z1a
P3wXcX1YCyAiDWReiRucT1bltq/gy65X1Sd6dqf73mzlO1rSOtk0epF6FqxQ3eVL
1z8vyAaFX19gxWUUghHHYfP03WirrSqz4fa6AgrnglIJmuG930uCnbKEQr/X03Ni
sv6drnZQGJhYyVDucRveUgy4h/10Wo6roFgYQp5sbKRqf4ztx2gwYI/UXHA2YoRb
jvIZGHrjUMG4bpmozs3cTI8+9gJTxlHAf9KHDFYZi3iG7GD2xnDMJSvUc6cmjcso
4fKEz/tKEQdILRBIFCDSvjn95bUaGfAOYPQLLGZyBwWfN8wkhzK+inDrDEbujrya
OLIUfIXLqUQmb4kc+Vn7jhUnUawwv7aB6JQloY7OF6goT2kpCM2QHj7ZdGCldcbR
vQTN1Rul/doLnIMWkNbTWzWUNxLk5UbX4tpqb2Kjl91KU9YXEi9qvuQTlDKqzeUZ
aeTkIEuM/QvRmERa+kCyxSlXnoiSeOWIFEcHAeVAhz62v4vTBwRWwuoXUbUrJzzU
06pS1LXum7o0GpDvCPz8V9F2KeSZqRUHrNaQbqslJ/+ANczWZLSUU8tL2hnJhCsz
OyQfnudcY1HhXqWwcm+55Vvr/QiSFd8BMJcyYr5PQ2YAUke4QkhR12M4dT7BjmGx
HUhNSe7FVRB8nWxz+4BhV5RDfr2o0e9xHxKuXDDOsJg1kr3Lor9bmxScUSz7nteC
qugMHZb4Fc63QDQkfeAF8LIHOfVUVvRfcayxT+yGusIqdgSW5fXE2uEjRpJHQD9P
vSqBVxu+mkbT7lzDrK3jhouxGG1AwRsbIq+/ENKLFnZxbg6YBtj/SSwxM6k2KEDA
lLibmpm4FEmcqPCXeOMttFnbWAAH5qkoRfTandiXnKAaVNtP/siV8ECs2OhUz/39
+qfH52dAZbJ5ZSv9Fl30h2UmtNNGZwyADU3UEdSrSQFaHGcwFXFdouCepF3zu7bc
VEeTIGk0ZdGz5xkbraLVjJiSkPDJ5M6mM8MSdhSqH95dNhsc3kYZ5Mq8xubV0nFz
7airKgb0PWaALWz4ZekwQSYF88geZQRM2Gz0wV3Cg4ADVzBHt8Fb9oOoRxIaeR+e
XDXF5GsTlDqcLbr5Udgx7LcXGij+moO/dejdutNqrTZljAF/1fNKM6yCzon48EzV
HjM2H15ILzRSnPPASVVhC4smB9eq6rM0vHWbWWlEX+uMs0oK1TT+x4I/S+QLUzN2
NyaIeFN8FI0zSHuog53SYbJ1Tdn+dDzo55adE4iWFxifVcpULdnXI5bSUlOb1JVF
zN8gJs0RkWJiYNByq0uhN/V8+EWPRM09Zm029xdalf4DosawyDMbYBb9WjUlmyBF
F/XZsQrJu9DEdZXpC4yt9VUNOuw92a00MDjFrC/ccFGBKZBq9dKabW1DAMXUd4b3
Z7P1t1nPetro7D0u5qaCEH+zaaYeiM06rUbeA8bBhcDE9ozGTufk/zcfKaq1LZCs
CJBPCPXbfcw43GDAb2vPK6Iny+VOp85+rDgPhHWnNFi5Li2/EwI7Yl+m1Gb0J2ul
RTwfiQwcnVhFZVyuqLXHCz5m6thndrzOwkKdo1yUsPpPaFDcsx/rVd6aRMeoMmtt
2neJqM5KULzFrBeyUsMxjpnr6PzhKVP1TQ8GfAQ4YtWLgL2lhneTLsZ9dzoDACoy
8ll8VWXGWcy9YuZ8TPJhRd09qsW0Ahv3HuQeedPLTVrMrdeHzqmuJiU/mHvzaQL/
dYaB6pFo7U8TW5N2ABKv952c2eaRf27H4Pc+gYvkGo0IdX2/Xp5sFRXRCXRt5HgQ
+1mn1nkCOahsH5dWQEygUBbBTF76xo93GXYLdfc6AmfrQpNEbTtg3GIBSRtCUSGV
UgZtV6L0SmPgAzaviZhE5hNPVQsVqFpMOA16l0eArTyS7hOpY+KJJ5iFJuKBLU4K
XS9MWfSFgz4Orw1IqwvG9v84upHex8bTZ3bvel50WZV8FadjFz5MLni6NyG8bumB
00SQHSjBMPd3GGg2bw2rvfodYhdebeZxhVZBWANqkgHRv8D/r3roeNt/uWqUDWkV
ml7PYcAxQ4aN7A0erI1Q4MJIdcVV4jwwWWODtfIwmx94O8vTZ8hlR0MPHyslBaCX
6tGZwv2o9wkgegiyA6POxoCO0bZQ8K8aihHSe/lp8HfIkGwo8V1vOZz+d9yYZOKf
NKJbmQhJaPzybYIYvvpdudgl0atDKIdTgq+fbt87P0Tcd5aPkH5OMbZqD9FXhWwQ
BfUAXMQDUuqMc4iiRtoeT2ZRJqpaF6ZfOcpMVsYcq0znuxC9Q0iAyOf4Wzo8HUHJ
3grVoSDMDlSXFJrXPxyqlXmDUxRDxK/XgIq//WQfhZj6hF4qr6UcyFUVt/7SS6ux
sJtBeFuuk7liSir86AyqlzgX3OgKMqi0idMgZnp+4rgcVn12JXZF7mVSABUcTG57
7DOmv1hhmGcujMfehQb9qYyie2ixi9hfwAa8eHMSq3EJIiEMgocLcNGq4lwmq5q5
nJLKAQD4fC63GIZXQdt3HpL77C6R6wRSd5e17x8dFsTlpBhDUp12OexRpLFAmGgS
AP9Tbs477AgyXGSlFcIaQ+HXQ6We0cX/q1Axrxiw5LOq1nB0lV3FTgU09YSZrbfG
LhhrRgCPgDDkFCdeym3BaoqandWTxsZt5HL2HWU5dZZd9QgEhl7MfU/pxvOGjLoy
LjDxEXYaNeKVa+QIV48dvD7dpcoxgQY/ymrWw5UWLyF6FZLRQu9P9SFwpt53h5B9
FLa2NXQFzkeay4iekxltQYCLRjTU90xV199GrPXRa4x0RQrRabtp51FbOcrJEVQ2
KTXFtk6i4CzbwSny1xt6nANJHGgF/1mzGyOneuWV09pEQX2i++hQvIFPHJ3GE+9b
RYGdB+q5n4+zvGPKxUybW7CAyG2elTU6rHy2GxHYOI202QN8thF/vrQc/TVzSJJm
47P0+gIslaOyasAKoV2xjcFA9bCg+wb+lFwyBeflCrjKixePWWv5qtxjDvfLLD5d
iSqdmuDxp3owRJ/pERpKcAerB6916ZHf5vjYoWVPTOSmQSYEG00enWSg8+xgmrew
Ex9iJKHep6IggAqEnUSdyA6Z4flDTZo44yJIc5jsD2eIhj+NSgpA/ZhrECFoqHPg
xO9RrfSFXCejGfWS0eu5LEpHMlFRsRmUPcR1f3qsrMq4ONp1x7KzOBJcCvcdet3h
r+vq6xXx3Zs6eIMVu0J1E1cC5O61hainYmoMCuhcUlOfcSFrvbDvy1qE03DaZEbk
x0Myapcva9nKFHNDEVO39ccl3YNwOrhHhSRm1GXLiexY3m6/nh1IWrJ6mCXxSIQt
sXI3q1dMSe2fDaSkEXRS4T+e9CipPRWUzXfryh48ncfoHS9F6U3Of8RhAI7rNd57
1E8/HOoi3PGL6Ol0fdYaQ+Ibzedu1IjhsW+zpj4B0hMeA6PdRahKhgSG1ipA4s6k
kJzoSKE/Eag3zpZL8mI4MoozRoC/gjbvKkuiViIP8VfCKxBhLwrVJlx2XRSJ6ngM
EZj9V8+N/uqMJn7fMA0d7rrCPkfOSVsAau+fB+RzfbvcMrk53zYgVJ63mhEC/VLN
U08ntpmeplXaHLyCkzxTnq68ZvJhxkcelg4adcdmMLzX7t87SUlgyW4yZbFKIVls
X6sMmJ1Tjvl3dr/joStmqlKulTKeQDM0SeHsY0LXV4ECeat7DLUObF5SWmGVExA6
/CMOj90OQbmXf0VzN6wnWc4KM7ymtfCLrnlRlmqjDd+/hMrP0xgPWSX6FIRvRjk5
fWPPBFKkOU9wUdV8uE/3n4E7KLZeH8z3tjIicyRB5spZBwEbG9QfkjNJjcJ6yu74
VZfI+/nTNJoYs85sBIbX9syzjrbbw0zB/r6PaXoN5NXxkXHjC/YET0J8MDGi6POH
ptZOBuhpT4nXp2e3FCFKBYBISS4kDC7Qm/LT6od0q8D1WPx8BGBpguTZ1w+xaeGr
Pjyl27HDOOGkX5vIovQrIuevQm73q3k1ssc8nqPzi1fLT0BLvEZl8VnbG1xX6lSq
sG9r1stZroqa/D/JZe6QPIdXaohjjMynoKGQtbru7zHnCXBRgGlLgAwSoIalilVv
bIhzNepx0SdPjLVNMbUdhY2pamwU2BdbvJRXk5Z7qKFFfFZWR6cGMhpv2c6C9UXr
per7zKfvt4be/4zuMAOLzmOfioNIvseg27PvQS8zMjp332VR/uvg1f0+wQ/YNw+s
vCzCUypOo38UzODrwCjHwvaNqejr+WcCIGnvpPxv9/0g8uNtpe/PxVaB7WPOItQK
ytHnZpN+XnYWEYkdIIP0fE9LpKEr8YWyzOpFz6BmwmxvCu8eaog9el7sU0pKQ8pq
/X9SjRTEbJ174hxvaLlNKMXh1XgzLaMiGg+oPJMdQ00t4tD1lY+0onusL1Vihn6c
25kopdq90/Rw92KXQjchzzAFx9uTUtuL3KE3psFkc7sq5MkgKb1zh4Tk4T58Bhnz
44gyaVjxnRSFIXfz8yW3+E49dc9qIQupsCrem4mjOFz59m7gSlxnhrpeTOoNq6DP
u23ntsiY0uq3CCsLcDUYuSDFCUDCoTzneDFowam+OICcSqQc5GKN4sCm4HEabU7i
4IkvkTiFhzJQqQ7E6HhMpuGMDmJNvm66FaP0rq8jNbk2vj8PQo7jjyDjXLVXxb2M
90DahzTW9ke76cpVUq4dx5FIRGpSU8+abuQ7K6DU33Pehcr/BUNpAX+10U4pn0W/
yuSsgOVvOEH3qiW7vhHSpjpauPtzoTchcvsAmH24p/aVech8gikWiHmiRIZDJD8f
pSTXSaV+Kq9zoBtVi9u6QgX+225cm/JS6030e/gy1ZfFwWwv28xQlAjQa2OgDJ09
yIB4TMfx/e/J06bzLOxhXvqZ2Svc1ebEQE+Qi775jf8uJI3/YmnJNIw//wJJAYt6
XgkzVhkI4c2VsaK067UY5iXlETMBaER+7q+5DxUEhD/mTCbLmi/2Yd2nDVtWROjP
zyLZ3s0BmM5qwN+RK4AQavNjC5rHqv2X4Pwn3x/5CjuEjZY0aCOEqC8dqlLggRlK
Wuqxl5tlYX9bweGWSsAWpgoRUC00qWz9skh68u5blgNj5J9Oy1G1PWGRMav+ccQv
aJ84NBuQ4ZfU8D1/9fH2yYopz8HKegQDwL7ZKsBUD7xC6iPaxC1CD6nyjY73/eYH
UEzZc9sIAdrDbyQ5rSxHFD/SWMWtpfvrq3bDOmBWqiDC9TTwQnJbN3/lGb8FPdwT
xaaPBXNzc8sYW1ck2ioATOn/CnTFoyGpg6LtKcjdpntA6/NQ1ikLyJbqV+gzMH10
BczS9Or8k/yjAleYFNEfZvIK/RqKvF4vgv1SO3TjzVqjmZvM/inVzV9L3PgyFB3h
+k2wqL93q3FyCwnKyB1Rcrja5KGnLSfaNCTmHrdkflYxul23XYqjXR+wAhoF4IqC
UPFGsQ89rvSO1+nLC13bSck1qlZLF1RggI3VVZ8rzuAf2gpysX9si2ywSS1M3YtY
NThWI60pAsSmT0DC3+r/iR+swkyCudRuGAGaTOR4f140khWbngiAQXcqCXEq7v/i
Po9YzwdYumWq2eYxeA756tkHq7gjOSma1/RW2andBevDt6FuHoeiYor+pfK0BMuH
+fjPdNh8HAHnHk7m/ZtpPc4RbC8HfhwjBhA0rtWTX8LT9fHOHnQ/83h9yv3Lb4Ff
PZFMVocBpY2LrxzFx6+17vxBR2BHbdg6NcpSXaPV1Wq6c9bRxKdjlw10WacE9d6j
XI0a95gJbpee92QsoISxdujB7kqwmgmYQ0x1jtzkeYmNrnOf4LT+c/pGfflzTSeG
dS+H2xoImcgEWzFEkpUSVa8YczhIrAYCKw5qQENRsdqyyhR+SQzxvlQzPDP7CaxV
Hpg9mfTqmtLC5ENCFoYmuWsKn6sYTSKD3vq0+wI4Cj0gSKcLs7QJTgjn9HeVCD2l
fITCD5Jx9Jsm0FTX58P7RgsqR/3zJh4dmAtQY+KOREZULWg5kcd9WHuy/4ZxXkGQ
9wnlEmHp9d2Ke8Hlrb0i5t2AH7isDhLgiQ0o7iUAH80gTVhsFppm8vvbclf4iRoS
NvI0VSSgWoBlud//XGc2xEmZLu8vPatJuerMemmcBuztI2Z2je9fk0fIvPPFlLgC
u4Eu6bRZ/+bUafepZLEyilv/VxNCpnAceTPgWpbTS0/gbqVV/TAe//to5a3GXLpp
BBkBaQE/9T+0qunb0sQpWpTvuO7m1GgwWyqEuhOisgt4t835nHXxKUtqR7R4FNTm
t4kXCF3uFx8Dya8/MFooGXD/2J6Ph1vTaYLDGAtVSUXHl6e0lxwe0c76aNeBAOs0
ZPR3U+eXKKXY/xWzXoDWspU1otah25BZbqvXROYLwfIhbHT/xGc24jZnheNGnbDv
im+5tBlGiD90MLrKvHdV58ieJfAtA2VZO4W9T+l6fWkt2MDOtIQ3XQuxn3sJri7a
gZ50NWgrl34wOjR5Qc9G21MZsqC2BDgaPW2n3QafW81nMRHZvykp09Ab39v8Qo3W
1XFH0IGtGyUEZFAlWVOTaBCGwBYXhhKW8T476QRxzcRZYMQSZvWJBabABJOx6lM+
jmE2pPeZU2wQUVkzeBiJvEgk+jz1cGo+cHicHDKt3q0eI6ZSK3I1YSovdkYbHYD0
6mhx/5SaZPH/7KfSqGqWRvJYiLKQtmC3y4VFPEos3Bmm8Phw+QQsmKqQyRSNvHsI
5qlHF4gqiBJnY/lRjcPbb83inAnJSseOwtdiySAVZkvbbves8Z3IS+E07vnRVOX6
oyjmQxSMWeArsw7cPLWlb1DrvoViLhvwjLkmmygDOwlw02oVqxmFELUhGffwu3ud
xjd/xV+eWJ9KO2e/Db20rM73KeZglumGPUQeTJ0m1MSQSSBo0ez68iQRhXWBCdlb
OKqqtLXuIKZ30BXHx9kk6eMJ/YIJ8Ey8gdDFiF+e982vwVeuIb8GS6W/y4obnpHz
kjBV303EbLm8az02bwYj+YU6F4lyTlv7/ODSerO/1renyXHZr1TRSMjxiu2BHEtw
5BvvqfwoL5V675YMmpCMWfZhxTx6TM6RhB2vcm31kQQ84kMakKGhr25K1HEv3UIy
8sxf/Eq57QAHQMUPeWUUmmYAHYqw39oHxshXVDli3gODzQmOW3DfbZ00Q2cDsK2s
TG0CrLQ4Po7MYXpN5kowTOcQTMRKc2VPjGPNovyk4Z7vlLB/oUw66mwn0EJMoedn
bjGjqWHp0QZxxaE31I55FKkhJunnHx1vbD45mfv2Ksey5OC1yNWxKGASfSu0stw8
EHb7/8DkYwru/09Y6JstRJ90ABdeiHuyN/ebFgYNDerT5yxE0tQ9M5m8ldx8Sm6r
xxsWgcHYNBhQ3knGt3ao16O9/E5GAaNYqPdGRJH3Byb7xNwMI+2NP5c+u6uxDXqB
SIs+ycwSk5OSwcZcEiHJmMVUa+Bm/uFLntuZMqOBSNMsd99qcanWBHhQcTxwsew5
YxxO4XHEKqRDkiBvyoD0bAQgCHRC9vx59vA6ecxAVBxOuZRLfC1bcSPprP5jPQwx
XUOvR+dnGbEOKWpadsv4KKaFMXVzO+sHnMG63YSr/aXTp0bMqxCpkje2NLq0WKcE
GtQ8tpN3cfopuIS4+FTS2jXvdXT24AKZIaFs/hUv7EyG+ZDM585zrjJTy2zLoraE
ihdeSbKj7V7/2U16e7A0DiFtkIuBwlejG3ArJI27O3fDg1HKUQ4MOjpSoR9cUMIn
wwZHpj/Z03NtX1Cv/7VNQyJawdMk17O/a5NnYnVJSh6291zsMYdcanYum3JtBxjN
BZJwpa2IjTiHxdZPZ81qWQoMAuFLP99ANntBo/tRVIjd48JnFSNCJg0WdgarzXtF
rcq9VOv667ioYz/qBD5mZ+CzCZt0f18Udat65bVLxCnKPi/zcqZ3G0iHW2hfnAYs
LHZYrts490/48qVYApqQLoJFrdmgotIPPqZtv+EWPqbyU/QHLPgbFheHwgVc4pGB
j2LLLhRL40XWXmgR7qm5n9D7c+AGxGB14FerkaStAW7F+y6h8xX2pgsaJHkdJJ6y
ArWSIkibZ/cMTR/j958T2QhRIufs7ndh3Ln+F3kWQotiI6udlFmVYsrHVSqRc8jC
LsEbv3UzdVYzs/qz+/F+12F7RsyTEccSC5p0mf0ZIOR0cM/AHs5y9LSDoaT8DK0H
XBBN56V/ACPV392Wn60Zti4MZdqpmuvoS84J15HEP1dGLmr8zzccFhLKF1ALGqs0
FFd8SQev7w5/UIBWjQCGmFjvOKQCAL7/IYTilgscdG7K8Azgde6zVOrNaiaBTqRE
7K1x9XO4YcYy0dJxISMjOoWLwpRdEq6wlH55sYvWhrRyMdo94BYVf74+d2jaZdML
HppJ6btXZcDO7a1siL1OXahMEheDzgcNsERL2ZyJ2i+UTeJoETkl5g7tdO7Zzt02
7QBKK/bsCnQiJgG6uFMaUY7Rikgv+3prk/yUESxgTQrxiecEkHRFlQfjbEJP9nTw
CzRMnRdelDAHs54K7wZAujES7WPSvaHTIfvkgHOA08ADAMeSKvfNXFmyfkHS7EOv
eqf+ItOKIOWEO/pdvrrl5tfK6n1lCtwWFbWoFdBLG8TjGOsdgg9xaHrzDgjkGhVJ
PFrCyRYxt8BKKb4PLXrhHERZ2O4pD/qFKkr6D4IWqoG5l156pJGeAh4HTASGuqmg
adknsTgiVILlAPPrnv/9k6WznXh+fncjVIt9YCiN99pRdwRM3pbUWz0t3eVC0jl/
7st3dqjONrETgl6okyMs8/gmmGEP7eNRJRjQTcuXuREQkiG8YmF70hVKKLPI0tlx
nYvi3ql/X9kSFPmWVJl2Y+vavavJCKXEttPhLiPiBuxMJhrH/24WAKmsorU7AhNR
Nz/tZ/GdBQKekxt84Gx0oY1dd4XvBoJ+5QOxYSjF7q2d6Z9PJ/jhg7alLOmIQjV4
AZqydu7C7WQXIlnHtmYlV0WiT+X9bIiztNzR3EO587sQt5bySNfhAJjoqolJPiFj
vSTrXGc1qWPjsQBM0EqiQ4nE89IxrKsaaNIM31N94cqNMffVGQVKKTMeA4NH/9yX
JD22RkJhNq++V9i+jyfwtxz7bcdsRmpfaXQBSqbDH+eHktN2ZmX2oV7BtD3kA53T
06qr6jRoMHjOEyZQOJQcwfzZx3nhWei+r70hmiIMiKMtTTrFlOBcATubGqkhUh8h
5C3FAWzFfN7urlLIo+llli3nKP5hgnH/4ErsP4w2KXcgDYlMvUlRL/mo/suETEqo
tHdO6RKp58bLfjlnTN8UBU4Qrvlaf/i1w5lIyPo4bcp0lVHptOg2iTWXMZ32Bdbz
M2pd1aQo11fIsH6eMisE+WjWa9+0gk1LFgHRF9Fas8uTRfxBPyOB2XpNatfbB26R
yAJiLmDkdigempALoIetQOdKnMx3r1pQ8oKDDAFgvgDXI89klV3d8U1KwMeP5Zzw
MYmCFXL2NGEGdlpxRup8JoIwzusEih6RqpKt5vR//Cd269dTIZ/IVW2NrGU7x5Px
YyCjT59suJhHkLJBcSbNoQAn+eGncXVCXxpOsh0ON9KGbFK8yhYHccUUu2KGhidj
WgIWi9eJVITsjvl0bxy4/ccgaMM5wtwVthFK+eKyTdoB2o2YShFUYS/E0UkzN6ga
6t1u0n6DmBIVAQUDsM6OwvrX+JECwrHjr97Cs01ymy58sAt4t3aLSdGm6Bcvg33I
XQD5dwR+YRf8dwdhgkrZbXoU4I077d+IbEvTH+eX98LCRdwCZLBrL7vYIXY/c1ug
U9aq6ww1ZzV+KoJsgEW29J6jQhSRlEEl/CWW48eu/KXFVpqWCJ0WEMy8mvAVgVql
aJ2cG1GzTdvuA0NwLgSaW610Yyr/BnjlVAlyhqFgvOIaIKayUNiC59h4aC8aWlcD
Q88s7SRnc+M9H7pUYv7ljZ35wgu5T25mx04iqNxFyYEzihyowMQtCRtGbqgmVQVF
AIjePlOn8xxv6hBOO12GyewjYyjI4v66H0dUX21N1i6qJCTdzqVXkRKuHYdckoUk
mN4vxhCPYAJWgZAopb41f8krpPWE5v9VZ8vfe7Fcltw7X49LMSvhPBt6c9VscGSu
qknM7F7CpF6wPcdEIm2m/Pu8jc64kifm51D66MWdWqk9ccF2QmVyg2hA6TmxP8Pd
wmYGh+NzI0Cb5OYhyjpSAEiu7to3Cc59K5OROB2rwmUn4i+XYJie4FqCxE3nyE7i
a5r0uQBgrVxi6X8GLi9s3ry63tyvZqXNo5RrHGYQYvP+zexAY9w5TnGgKxtmSR/v
Ws+YNd8Og+HPYTxPZSzo3QU+bPKu3p/cAKvpZpmkYZmDr26t30Me+utUBeDH6+Dm
277Y1MnGP6S47DXfSwYIFlzf5oLAujOSbnxdHBW73fG0b2zpqnB569ActM8LIWkZ
1pj/e0v+lhQpqQvxC/jhHvRT9WyS20tA4EPTBdDV6FQ3ys0JNazuXXPDgeO+2me9
xU9DD6FBfFOT97waSDX94HkxTOHflj4Kyf0kaBbY96l9Wy0vte2OjNco63RmQp67
hhCYA6oZvDV9K9AkWZzt0lU6aTz5/LhPR5FQv20TBtWJIncA6HW6Ox2BPZBrvNla
gCZBBtZODcxaxnVtf3RpJdCTQ46wfk68FSM6Nj4TGLOTIHJnOQlObhGVAiLIH6r/
G0I8rL4HWvrmiyV2Zmu9cFIBjxFQt2qSkyRp14TzvReYnoThmGtjNtAt72s9nzQn
0dHw+sDnG3cDJYrmljze39CS9aSVemLUEo6swUwvRtjAuIsHrHoAxtJjkcSNdcak
vrA69S/7Nkn+z4qu0op56SXe/++G+H7ZKK34fMGMKQYrhGumldyjPvtWDHPLmWfg
7iStFIB5Y2yJ3LZjiDwqC4ZFVbIIDjFzoSSXEvJ8xif2iD4Smf1KF8FxmRhwaqzF
2jsgd/iUDK9ihUcovbEaKnl46Px971rMPhywHx57cM/dEH31uSlX77S0n5Q4oMFm
P2O0QxoISf2vlKY1jFZIaqF1tAMlGrvYzcmc+b5whsewutfniAMcJ60plwVB9frf
2/rkX//RUQYvoVw9m3cDD8Z4wNaHrOUuKv9hTqUTMVsuFHrSKuXCPoxUzwIKB8Xs
oKPDP4VOko8jeQE792YSZebeK42DitzNoBiHzgK1XdW+PUz42Gh7+l6ELqQpj6+Q
96jIkCIkTdC/z7yX+bTn7Wp7BMQEgDkzHh0jkpTV+JW7XzkyKvCu8HQR1YPMeiXL
xIU2eiKNhBNOZY4JtuxKEN80Uryn/A+BawwBV9U+rW3mLNJp+iXfFqcH/+gXc++A
E/8m612WrnJGjmo/EJklY0yzA8XoNRgfTHXjkpivtiteD5TDMNBcrLLWcasm6E96
MRocnM8gykXx0TZhN9wItCigcLMnPsPfy9F/6OrSBwveilHdhDkFFu+uEcFEdTl0
0VUANPOEB24Qi+dyUi4hwsCnFuqgtAif1UpTEmgNKgpid5EXkjBIaogLktoHft9u
9bHbBgpFy+WYFPPGOrhc1eU15lfvw5zvzaQ1YTxO+PSwaLpnv2E/G+zRTD1x1eLN
3rdNwT2ITtfEyJGnCkRA27AvYjIUwhjl5fV69QIUMMZFts+TZJCddft5q3K4JRlg
rmuQFNxC2fe4vMMGCcq42fFnqIElosLCe6ovOlEzmd6XL9hQlnDhKZ4pTBSIRboD
LDQ4JV6ExMS1cFJTpUgiYpqBwsv9ThN2Q4f+gTk9rgg9vvy2lnbQEvDkqp7usTIu
0iRmqnTcmRzoYmMTA4ZAAGQtiUvjerDVB6hvsXgg0+otwZ5mY1FoHLA6Lluxqup+
J4caRKEgpoBWR2T4+GQRcAU3D6okIqwPyOSOcoNq/lH9hMTIVUs1ehHN3CMfKX7/
lxv6KX5NJi6/ZcRsb9sK8jqHJ4TrFtGl9OFwPf0OUjpCRXQTLVU6d/+IMR2vECzZ
/tLLyctHQYFXXyiWgnwbFCkfFVKPBmc/YeMMJ1pICW+ha/MOYSA1FeNIpYHR0STK
NNQfcs7hyYwEiDvPXoYdgQITAoyg/GSBHUQyvQ6OR4seb0ezvm93VugoQBs7kwQy
ste/Q5Vhymj9P3W3vMNPRNWpLl2jEE7uuknvViW31DtkmnNU2L/8bhE7Ei7a3C04
PsbN3J8rdiKYnp90Sdgx2dlpcK3fsN4+yTnUpTx0RAKdgNHn2gL2m46ppxG9LXMZ
bmrBqxALbhgT9vZOI/4vT4qTk8kW0FkfknikExafTnfAttvdyBvsXdIWZm1hc662
WeQhjtqtvU+rFbE9Zi/aOHHK69JaQKF28YxwsxK1nl8eVC/ID/BeufWBz4GQQzaw
x4F/CKUc3Niw0cbOHngPPbhWvFCja7zRNUOkmwQCBNzjIsbll15nkf1pk5kdQJCx
R4R1R3WW0FWcTvLBLJ031WQ5W35Hu7osaCbz51xN/C0Cz0Q07V9NAyp2zjuNghy4
t/ws3X1UFyfe2bJ1/DG70hR0MEsZAv45g5r5H49ZAzg+Kh1qPy9vxZl+mo/cN+wW
6SHEyVJieYGIhxsnjpYlBcP2LstTV231HrgU4F4binpL0GihaJkAVo83HVZT5rg8
ttN4KlISj3JvdTyLOX3C89yNvcFKOwco9RKZS7ZfJbn5ckvdOYQc5RZx0UXg4xnL
zj1PeEifRJTiIi/7Hq1l9qtkRRel4Z/z1UW8lQ82il3o+f4DCBSPAZN6AurPROZy
dxxK2yIY1OvBR7pcksTzHyXKblbZ0o2+2Bh+Is5iaNLza06jkeLaPNIYN3Zc+fd2
Xw4s1lwcGiWHsAfEeYol/UuJ9XPVmq+LIjgrDVf+Qof/JJwSeQdbPGvMAA+aEphp
ACgBNcAoJDTf0oNIdKGtrQhOaG4NM+BDxfGtHD/xQTJFHElbReXDLkJI1rkjEL5P
0emK8VOF+bw8r5LZPeDCqVRh/Z+1qLdNCcLlNVfjwJFqgoj1eJ0vjdyV5tskLPDW
m2Jsvpp9wLMfVvONYkgnRkiKh+7twPDZKcTX0wOFbp8MEqPFlOiDxiDCUn/ITC24
aqCvP12J036f+/1FP3B/4CLbyepZrujUr82HExCLwAHO0rVPAvcZRKheMqXnESla
nQUlCwVkAdOZHIt+p6XCqqKwGNbxzLO7ECQl1JmOdKibpnMCY0TNhauBxOBrmhqJ
rLm3m9c9d/iED+g5EcfXRRljyaLPasNT4u/c3yaSythvBqrmjgoGfdgmF9ZsP7YB
X0+TGf6VjJHrr+P8XDd1aTXQbyHLr9V66AOosJVROonKXr+m7f/MCkg5F3bYT5m9
FnBfHUldGIYddE68EVBq3AOv20mLe7t7G66mgzkOSuNzmi+uCTHNfUDpvhafWeWt
DapHgoXPFF6H+ITxVDpcFWDytzvTAsMvMHrKoSvzyXwhcYFD4DBznWCrby0bVbJ0
I6zMyfo3NzE3pTNQg59Hu42FTdr3/c1RCjBm3tMN9ZF/NsSmm+Sg4MQ8zPZKbdA1
2IEwQbATMqsDTR/cjeABCUgrf2IJRlxPA8DmpH4F9uuZkt0HACugVGZg3j/Y65Iz
VsHU1WjtWpiEivhcEgsBoTIY9AiWcRKYNuboNDkgA664um0Oa+pefaZE4YTiNaJc
vhWjNNnoTzwZmH63FtnK+aytcWoZyzdYqbJPRlavFpLFyTemNgBGRJK/IB6oe+2b
kUmFsL9PsoPpxbNxYIRuq6J9damzTwVRZZqAVxEjifpsLmWXiZDHfmKRsdZsM7+s
LRpxyq5uCld88FFhVHbFc3gWy4BAL0rjvPXO/AW/nw+sOT3MtMpiwNfmrJC0Y4yX
SrkiMssimhb61aSJw6KzZmqqzcaKysYMTfsEMqFmpY9lYXNUjmvCcJDR+kQyYmaG
NRS0G78hZBfb15NxWRXLfvH+IANqQdB8guH65jcz2szPG29bH+dF1W+thpJMFSwI
UePwxWXDJX2O/h32JjFta199bpf9qG+Cp6Lurmkyphk6LIAGSUnLPAphLXwRHYTw
URE5rg9i77pLztUIxyTToxJbSXajbUmHRTWsuhlzVnGNCVOCLp10G3Iop6VHAFCv
TWS8gXL2V9alIgi4Tewq0+N9IJmh+pYmM5cGssjxkWhKCNISlMXUrAhtOVa7/GGP
0D5WoiYCBxXM9DBUYZFlq1ul+yaswZHsAXMUiDZYm5uNJI9eEQW95JKIjWweWbgG
6jH7izu2/NEN04fcOf6OubTLOJs2ZtOdoKKV3AYRhYRD6wz2RxXBN9VaW2DwU0DD
q/r80v7RMSgRgcAxC8Usewp5kvG/ZIt6oCFSCns6DXGqbXDOfy0Lty+MuLkHtpf3
8griwiB2BqturAhhHvZ4u+/nies1olJ1MTu3wnyRjOfxIqY5Sx7ORsWInvoJog01
iX71jkrkYxSEYEykgoertD6/TFvmpiNwFiaUlG/+GXqdr8mE1RCnmMdMOwUzM/oH
RxKoFW45GZQ/HQr90RR+bWaDD6mjxV6itv/sBBhKCv8ImCxMuJxA7n3k5+WHv6ZQ
tHFUsJy6fModk8lcxLu892D3EHroLWrt9NlR1iAukmjuKSyrN/+iJWtPop/I5Z0a
jcXFjW5JJtyQFLs+MlbIVXvoMfCyOG7noPcmsuPOjmSA6w9S7uruSZIBzokuyBKO
ymLoKTeH7COgxNI3Bly2FbWt/wiJvkcJ4oqkw7ScAUodReNHhqyuKRPTpDra/yUI
fXAmqRyrO/YXA+E6aHr1X2r+EaZU3RykuHMM0G3poO31zAlLUdieEBFeFMpOl6dH
j6WkfgdvghM3heZOXQZMS6xyWJk7apjHdt1uyqaEH/mky48+0JpNnl/crZSFzY/B
KrAovxCX+WgIG9/1Xi6MZIDidJBu1qENH/k1mzhwJXwvOEkaX4L60aSrZAoDo81V
FI+NXjwygh5303iEVu7rd/+l1VMbmcWtM80ZU7yZzCCgqCp9+4Z5y0qCJgkuUTXV
LG0VnOR3axpv1DIcE/4BOW+iG0KCyWNDBZAdfDUmb+qJy6V9kvWPuwRJDDk6kO6c
YAVU9ia7XN6DmLVbBDU2QyhYKkyQTwBbC3oWl9gVxCNT/foTj7AKqk9KyvOJUIg3
ANBMPOyMgbDrNdH9lsUhslZThKTzpoXY2qsN4a88ELp910HrK48VrAw43BGaDNCH
cYs+oyj0bvYCCf89sKx/Hv86155DpQeGU4WrXoOKmZ5Yu9F1QvqQG5ODHXke+cHp
EkP0QBR+6I5NzFrxnFygZz+rlcrR9HzeZN7w9nNJb1noOYjy4qslCx/S3EDsEFeh
dUFIn7wGPubNJ+Z65bqV3AxqVKGRx6Fs4AjDXX5MD/gTKq6QP6k3PXDDPpm6EYhU
4H36W+braA1O39gvVWfaapAwUXovZLO3nFia88P8ZTPbhVuAGPIfgZKmjQnTudN8
J8/5TLLZMrAL793x4FfFkUyG0x4TBi2ltLyg00m5KPem4rhJ2opNLylycEP/fMUq
BzSqvcDcip4egJ8EAmKYn4ZqkP2xz9Fq87oegYHHGLAdlQGn1kOmTwnnaPIG45oB
rKyMZis2UZD8I1V16qXcJ4RFQhFmzyZyEpkz3j+8ZWa+FpGU+r3//5fIYwngBUgJ
C6eM3DJiJM1sSqTqpS5iosmFQ6d8NqCS6Rfy6pj6ANALCZUJBSWS2KkU2nI0W5O8
Ks68h/0YlfbTKxf7ItGZO4q1wlLQ7YJXcxicIlD4lViuljI06yOiqYcjbQITxsnD
jAgvL3JbpiI7alw9Slfu6NS4DGFO6n8z/WI2UIMd6q0Y4pEVish3FpfVz12JJaq1
KsZmv3oLMoGlAWA8qXQBOI7hhRnfXkTjuZSpOGSTG/rwN6xln2hPWiLfJTrZ478b
6G24m58J5KEDSp2EsKclRI+/fQiTBe3e+tiBb+sct9cE84wcdHLajlAO05IDzb4i
RvjLbPdOxJwnlhrm2zUds1sNDfug9WT/OXrWwIJtpBP+91bgnmO8p4GkPjFwwptD
wZpb6kpk7wKyRkYJXzaR7vuJRbZ328frwpX5czfiM5AOuN2cU9Lpd3g0nXVgwLjl
o71pdepUgh0Suy00f4gbUg7Z1mio6N25XZKLMnW04Cyd1ic+vrdpFY7dJAl9be+9
GIl40/r+LniNjc64mN+kolsSsmWDm9bywRVZH2WqBBsRH9wHMjumhek6xrLXC1xx
xeQr7UYIhkMEYZEyk0L+7QUenRKugPseFrbPKGPKQhoB3/FAAomYNjBRgnT2QmNM
9Ea8o/Q02lX/os53Lq1wyyZnxc/JcbdwVx1lJbImtHjdjuuPNC+2oyQn3V4xBG8d
7k1f7Vsty1b+Bd74yhiDMfw5idnMr7rTpsEW/AzMR3E0En1omr4o0knXJHqBR31/
BDUAuy5q4X/5fAkiQ2ncxBk5oi2WmA0MyUZXSBfuQu5oqV/M4Oc8FXhJ/xJ8Usrq
iMxvkjJQDBFD0ZunEwFzZNydQFGbwATHobb0i8uSjsAIc4cjpXwln4j6GvLHwKf3
yQxuhEUvIEeRIi1Fnrv9b0RwSA1aS9N/i4VkdaeD9dAM2I6rXJ8WWetJn35GoVSS
cmTqP7Tvk5eW/C3phU6BwcFwYqc9OJEalpY9tFSov442/IPXB+xlTSoZa7jFgoAR
X0t/k9Nvwn+uZO0a1UnmyiaSBFQt1FOj9VzTQAEk+a2r7o6u3V8ryC+4lU8j0r1w
InDxZZX7Z9MisfP68dSNHPJe6WRyLw5FJkqsTjeUbBL+YCmQwFIv+YcOhq2fq+qz
pAHmawnlXRm3I6+PSAzzKczrPE/+sXVmQ9Z2W4l9ZhbOMDJ1lBFarOPU27X8Kn9d
LeHcHSgWlUmFW0rX3EyQYoJLr12/GxX8aqZ38mplRO0CAePOsFOWNS0cFvQCLVnq
lHIFMaEzP4uyEYvpHSoesuTHBBVbr/CHLaNtcDv+TW/mHY8GFmk1BbwhIFN7kBmq
fpeWfhDAbMzkt4LUCiHMqo871XNBqQEi5qO6w7vjlzUwHmfHsJMlESTFqbzc9PqE
wU0sPzVc5Hw0dl3V0pPa0SGrCRxkggyapgatandhDjDYFdTIFPG5RKRUvFOli7tf
A8+U2+ieGtJDgd/u4TKShdf9dGsuIk600UJQkM5vvvcFXSVi63TYVwgSAIvYB4Cc
qAJluf/QggU0NA69tUhaIO7mEwY+CK1UVmpOyuQK650Jd/cqlD7DvCubWDxklxN/
CtCoG9Ts+FH+H2M2Sz76fZWRv0/fV/Tpbaic28Cz0yHFVYRRrLU0xfTs+wPILi2/
l9/bvWUG1csFcn6mN4JQJqAWzjJlGVv7IBgkrCdERbzvFxZ85h62MBVZ2eHNW/wp
7Oip69as5RnV1W0afPPEQwJj01zsymAYUWRvvH9N6D30DcRQD24yEHx8Tp5tHZ/6
lBDLcKDY8G5B5GCFMzs0FugB95Bp+YheT0uekctUCcbg+tPzfwhrI71yZ5VfDFlo
/otbCxVhvd9nY3TYwF3lqolaiXrgU6IKoxpx7ZwXD28QOmUMF03za1swFJ7tg4Si
xPogU8/vzLjNXeSZNZmC9Hlc9wvOFK63Gz0WcL2LAWdKjKsxidvKQmL+TKbLH0+W
71GUbaQcSbtpZ5geSTA1o1H4s95g2/cimHgyz5ODSB3TU63nUR1gz1tw8O48+y+P
MVPVywhnpt6aKDLDq9iL3G/h8VVAFiNFa4L02FB/FJ7qgRxT3K3odld2UQxqawSE
m/2KEACedezlJ7b40zTwOTEpLtz4z9Tm4tzUETn7LpeDBYom6hT5+D8akkoH5Tym
3smJ8kqg8jhmRhOwgHbBO9A+lZGzwMTmHp4LD7dohZkvJXik/mek90d5Ue33hVSG
oh5r3+0NGBlfvX7H9QxpUsYgAG6J9AN6PtacHPtc1cMuYUWfke+w9eUdHsrxkyqP
qwJGYWGoIpXSx9b7X9/TwrbFJJO8OOL9EHNU9Ft7NVZhSdxsx4KYLU8DauMz49ob
5GAniDrJOvwZteHAt09SW4la9yPVp74FTA0wEpra+NWSatdJqZ0yzTe7ElJy6AOY
69TW6N2GSa+/xngG6sHT1S0UD6takfRoEm7wemCi8gbSY3I8SLhXDHcK+fM9efrl
1ShcnePc1DbmkuOhAyopPiOOxFjqAGscL9uxlKB5o8pU9NTgXSawrWvn4DfXN9H5
xLgcQYAqKP6eMVreOZ/FkV8JkuuFmpSbn+nVyIt0gwyuYONv3fmOrUZcK+mqXVNy
lGP0t5lcUF8HL2Un/8PfSiUtHG3NEFpUUvUzOXgWiFeQ4MbjkoVCy8wH7CR9geXh
WVlLzZzcbRVkQ34/zx9VGJ/JjoSw06kglvJHqcHMQ2GdW4tzoRba892MFzMTjd7W
YdQJQJR2Rk5a8BbEVyWkqbt7aAZtz130XXJ5NlYj/45C63dfKv0FifPd3hOGIrIS
0lXMnUffcx8T/XACOVFyWy9pq0pSh8Gz/OcPiOpL3CL/Fin1zknAYKp/RRiBERT7
hSDMXpz5wTNmQSYII2z9796EXDFnYMrUjPrNCXnShxSUoa2s0memUhveJEWGfSg+
0Mr82+uthtcX7clGzhSiZKzAiKg774Xe0d90UAMoRjsFZev5yA4XC3rxYbkfIFqR
uJVfcXFp2pSt7nM3Js5czrQ/bGBVc7S7fRH3VaydSlANadm4LAr1RSdGlcO0+ugy
PtNt8sqLRD2wq8WRwf/DMDcJrVMBEuEcMpOvx98JJVOAJAAU2oSe2bm6Y6YiwNOv
xZT3SHXQ6kfJo8Of9klGC+/jO37y8r9L/e3wKEr/eyi1x1HZiVz90ediyaVJs6/y
lgdbBFCALIm1P4SJyqtlbm0JFNRKWkMu8lTHWFkKncyYudN+s8yKoPsZaPnhKNJm
O3Gi6yNuga+9xnu2MjMjBhIKvbA5AMhgdjr1k2QYj9ZYF5fdqa4L6gotkowoEisa
xNAib7LDv/TYDrehXuM3O3EKxbwVtNLLOz3iTOCjpQDRTBeuKT/AR7Dbubye0iD/
A0fmhKNLjpDhCxaD8Kdnnd/JdNk10TR1cIGA9YompUb+VIw+kk5jq7nsgUz6NpPW
wT29mRe2XeAI42ru6tYQ7mOguhrWjh+R5LBRsMtSTVbNwN70VE30ssXgDtyPLWOY
RdozHY0x0wqEe7q8Hs0LrlgGsycfJuymuy3lHPQ1NiCP5KtPhqUcP+EMVHss0K1A
i/gHYNg3WylGbVj3HRXG69nVPgoaxwc3W+QR4SZU3NJ55OJULxCR6StlOpf/7y+j
0HzGaq0JZU3HzdehnF8NzlyXza/ToOL6VetfK7tlAL53RPGGUbdEgfLLzrJUbGmS
HPsMOy0s3ycS4ROiQZRDVv/C1h9To07stejGpcyB7fOBOjI5ZEstkLdNERkcmAlv
t3lIIoFR96hSQBfea8pwLrI6bfluBzlOrmvvcqBxNCy6yFoAraHhsDbuS2UG9xDC
TWWNj4pKet31Em0GQryKRHbfsp9uyx0+AkFn0Cj2M4ABM79Sds7qEKMmNSd0eHms
w7KRf+m+H9dgdd+5vMlZByiliICsin+ee9R7+mlJ1m3hWh0lErTL+mS6zhlQGJJY
8NAdf/djiVqdwsB4G+sI3dFM5w6+fbAD2CmKnypS1ZBXdKYiG/gn4UG7ZbYUsLaZ
PiqwJwePl+ehJrrYXbqyzX7s6XWpDESXvbMng935vmXeTOb6vzT9Q0zhd9Y3kv4h
tWQARQEZE5qN7YqYkeVZJ2D43XFvF+6poSznQAw9pqCbjwqtahl4s9B1T7GC3w0T
Eb0pwyyuBkPzi1mw6588TPNG9vHnuEY1sDKuG4RT6aO2FRQAuCnpihngEO3g9wav
giq+SdwoOUcyD0ANo/BStT0n3/sbk1jw7WtEhg98aah8Zlq+ipVYE7oYWaoL7m4L
g0SbxQxrDN3VL0vV8wM7S8TK3Z12fCrajRdZ+moZY42V1vmAg+y+PfPwuNSLr1EJ
gRPvTem5qph89vXp3KF6RUSfINgOZH6NPa5tPxQ3NIyI/pvqth0ZEdF9bOe/V/Lp
su8uKE0h9KNT/XMaSxCTEdV3JTkvPPnjMXyRrB34g8Uc/jdW5yIyYRSMacs+NkIB
WE6GIzxxBmGdRyqxgpHOq2azacaN1Se+X+ULS+grx+DoNppWZan9/EN94VBDCesU
8gsn33Mma/Mc0yQsBBJ5fhBA7UGArRRXRGEPD8bztv5tpHIum+iS92QrLhNrdxB1
Uce2of75YSbJMdVEm46SIHRsGrVLtVX0yjtCk/r1pxAFGexCIAy5IXWjbj43G4oj
AhLzhuj9fqPeDn6i2DaRnmzLGHCkCsjcsYv4cC8ZVUryhPQVoBDDgUPX+w7lxCof
svH5vHptSKv8Y5Nz9kEqktjan2fg7GL5XnOJjDRaa0SdRbKJxFfx/qZoya5reYqJ
ojJGtwUGs6TF+OYvJy/tlVciHS2+/JiTOMYbOM5yZccHcfj/dLfTaarTaRN5Bb8O
0/jkYq/vhdydNLFdsFpOX/pWGNgIpWzmeTHuEJBnwrkqFC1B0R/sLIEtls6OQ190
e7ax3ttTGzgtuOhVbWmOdoSs/9toDWg8+BKd4p4d0GcAAc9RLj49LHSHJ5AAZgbZ
7SMeqUyvcrMP6R8jZB9SbGFg0uN3s7CrvKN8pUvgdQDcNBe6kcf2fB0QmgLDlNJx
0RYgUgRMFhJvAUbwOy51FJxD0DO2oc5Fsml1jWh8mwByPd8LS4z97Pc0yrBNUqre
v/IZsUTXWzFn7hyFbFY962RPfz3BJ4ats45P2XMF3Cx9PCMYkMKZCJxLeGx1VXoA
GbtYt82kI6s+0RGFhZfaxTn/7EVJQP7fRgVW6IZPK0/D4NHMlZZFsEXBhuLTnGIO
v9GQ7RVfXhTdLt3DbDIncxAydlqi4JfiTPPKiLuvxSUjuuvMTQGqHVU3pYqre2Bb
bpQlWWjvDAVaQsWrAQPkg4FfoRbE9AM4vLNJ1pXTp43d7btq8Uth8kOrFaN/m75F
b+jKZgeI/wi4UMeokr8y34o9poc5szKE9wRi+In8qBDtFhGsXYm4h0liGprpr2Nv
gi597KxggiNIb7ES+62VwbJEzmjbBByKr0Px2y019WUnu6X302y3rHHOSqAXsHzj
Mj8Q4epoX8zdUTpFlCl1RC9Z8UA3vmbab3XJIRm4onCtx2rq/rrY5HBXJABVuCmq
SCIMn6bctscBudM99Gbpb5QDluHry+NOMChn67nY6HLjpgj2kx6hGTSHL2HSFGMu
swwLofYCBykr8zyK59OpL2QGejLSqxID3BmXN6i1nufk9tjz702Agk1+6R30OS62
7Pcb1Szb/EudNtcVNsqIOPwyZxkgeZ2j464ZAbOm3bYMxnat0jbr/rn2JMAkH97D
EMm12qgZqeBe5tI886Z6tCth61BLtDbdFaxQBhKonPHsAIGDAVm9aUIdA3fLCsVg
bqUQzawY3/QlrNuWL1lC1a5p/sZbC5Nf9JUPhWEgH4xUlUVz98NMzM1vd8kvqAXn
emNlTjliwPNUcmq+RhSmUniqgwHiQSdDZg9XAqPYk3NQvy8p38ifIPpkwPqF1/xV
HEMopLo3R7ocB7GPds0H0wSJ5wh3aT46RM/F1S2EPV6bS8t7u75qGjUOl7qQLEZ2
hDdIet/D5g3F6urgEXDcM2sb+ZcLoqIaRpMUVmO7t4SUevM5VMoWyDfkTA9or1Vq
608Mhv2nxM6h6rJOi/XHwO2JNKrL4w+BFAScU6iha3KT9BEoZC0gqqcA3VQI66yb
EWUBtxNoBbrGuo0zcl7zmupDcDiyugLhFcGRH4oJ8Pr4HTdFhO9TYcg3xTImflKN
XhPgYfllpb/6j41472Obadexhc/mDmcKVvaVbEFmk/PUyXIBON93V1zXGNAmAc6k
0A9zwziVZYaycRt2VYuDP5p5FSpubWF3wPY74iPYvxSeEqRFUZb4bNrGuWyphK8P
SOlODJRHboASai+feyPmPfh5mMyLXaWRj1QzUZTYq24Vy4cIpNSds8dNS60+A9u4
3mq/0X5EM2wR1VxqzBQXdFCfhPfUHuyaKR5dJg3i+14poI8a4n+zp9+BTr5//67W
ExeTMQsojoToFqvLAN3l9aGErjpn8BPwNoCYjpMA7g0YH7uwwsuY1UG0BKjBvKfE
VSbEYZd1zkojZ15VgyvNvQUw/GCnuLnvh/XVBdcYy3olRzF2KNpSxoKtEwy8/RvC
UVMjT8DzD2tQcxY4IgMCXVK9GkAeDEhsNjU/GYi5kRspzeMNX7FMRUUhEwsSvBfG
CFjGAkXrs1y9PmqmRSsANoumFemldgU+gNbgarisTokYMoDbVO1mem3TWPTLENQD
TT6EeT+Qpk8VBXAuJi50RJTglqoGZqfI8QUE5JdMdpvPPLxXexulCq7KrGwmFstO
y+SYaebsxkZMm4X4yrJPlAr9dX9VlDcBsrKu7zvA5rRuxCUR7yn+xTH6bFrN/RLU
H37+OHqXOlRGLN7D8lqa8wxeP8EeDzDUzwEO/ybgpM3MnMgVfSWKbPcayPAiAeB5
OSBFK5FhjsRxkW+CKhWqmvDq84DGaQAFhrEN0j7p6zq52M/Lk5n8QaTzeEKS5kii
OQHoOzG/nbkLRL3XKTBBEsUTrMXCLn5exk/qOHmyPGLcYQ9I2XwBR04sw8ao/URH
Trx2P25C0X66xlHVJvSQ3s0vX89ksG7ge3aCIdceZ/zS0Pcxef+Ft7rQYBbcETuU
n42CDcmb2HjO0BkwevB3K3Jf7QtcOlHSfZ98ae2WUoiZh0UIhhzOqWnoQbl45sbk
p5co/zTxKg6p3QqhmXsXIRJh+Qvxdiok36QBcg1UxnhxHxdJpB0ryOfvCUBtANqj
2yjmzLQYsBzRr+uWk0imA5ZDVueBLpsCgmcvCpQSVHYjKg9GFdGLeMQUVMEOd+tv
zUGFhJsd3DUVu5RKEA4Rycbr5uUCdhtqVATUyHFpOgjscMu+3WlyYJ7PIrgAcm+T
1Anm1+2F9qJDHpTuoQ7dhGcOkaMr5e2gQOqBZ6jJuHFeHyDWSmW7Oj8DCj0aFare
n0DT51GPy7x5kdtDIBqmcNiZ982Ho7AUpTeF1MDu78JMxM8zmhNZoVUtheUca9OW
1pOT2QmCMkiUXa2q2v3hdt9eZ5g62rGFH1S2ikzNrSfZjZLEo25yEAExKKQ4Wfgl
WGn8YQaFDXDwkNU1YEbXqOL5dhMY2J+e+Ymv8nYEPH/kActyrKFSLJvkQii2FLyU
3ZDZSwnikREKx7Fhme/YppokVczZ6Ey/o/zZZ3hEiqz4bOKMz3QoHLZiuuSn7Ra/
qrlG3HMZnyPECkWJTj6rWXgQefL+pDdIXP+ccDzY6hL3LfYZr9Y6gdx/16DgOu4k
8STwc4QXhFSpRE9cqqep9921E8v/wvuLYqgeKZJgOuqJy1Y+oEc3B6Z5Eso2Ynq9
TDEJm9ZK7G0GlG/A7cfqjKC0JQ1Y5VhJa7zwdQYkklfipvvf1Ex6Voi9QV0QSDEA
uQJsj9PwqbxDyS2sXcvWK0YYJzgMwemcVkdLWAXXeYyy6TGR6JR+dLZ4cNuhFD3e
coo705l/Vna98bWnRbVuw4p2SIQVI06Sakd69O12GVoQObImjmwnEDbJAftoT5+M
00XX7jiAXakzeC/Do2OJKNRanmBDwLR9ByXkVnSum2IhAKtIZeBw+hwUkmZEsuRp
Lpb4fwieWOJV61jgU+QLFVJYA0Pu56BAw1p9si0wQiOVhFqj97LwszZlxQBFgMzf
oRvV5aVtMKFTMGQgDiijp86nHcZ6moLjw5Bz0pKEVT4w97SWj6AglPzdtuGyWGHy
kr9iUWg9T6RuvUO9vpVyotAe2RUI6d7wBp+12YG/z1z6HduoHb4cY8VQdrf7QzhT
JJlJLiyrl6kW2iHfaFX3jCKx5ePAP2cVLM47e8smus3ngnWdOH8AuiFVDG9fuYso
HLQBuSW/nl1wmtDHYN33KNpIMSpACpgRyURD2N3Q2B0PoWzOPJNSLSVAmqvDpJz8
ceUi7VFl01yRFufTk4NqPUG06/yLyOlDqBj/2atDVIHuRptrtpF+oNiAprdIEVTK
+VsRmHy7Toy546e+xi9vnrMue8yQ89PGd9davW7uWXuugzQrxuVuE65+LCj5k2nJ
NmgpOl7bkM7c64UDDyd9irgTrG9MhfwkjO92xw4KgGyfLhE2y051Gqdo+RDBrRpd
Q0ifkT8XHEn5N61PEVlAwkvV7+OewDgi99HbDWCFTL2hwPiIdbZo4SsrFosE+wE2
9XegSj00rzVZiDqusRyCPITLM8RjwO8P4phPuvCUKSD6cOlQ5GGdzVYbjMCzNd4O
rD6jAfVTOsrk6/cZMu4jHL8oqfzZR74nAPnshwe4VANgLkmrgVkdloy3vVo2tNVy
g5EP97MhkaJmiRLjKigS1Wlh647GVrvzSES/1WuBt+Pq1ec7em7ify3XWJWsc+1h
Z4kd2Ie0jAlpDzX6Pfd85jXWdvQ6HpMtrisLPGHHPj541IFv5xf9SU4jM5emhc/f
e+pLgjMOn/AmzZitlyKKvHLvjkUYiSFR9kKYkdbPaX3bFvYr242NXZ4Hylx6xJH8
StoGKuOwq3mi5+CH+uQMgbLGvXlDXP1lik+Y6DW5yMJdQ4ORYPQ/nnpqg/OMUHls
w0QRT8mpp+X6U895wcKht2eoLehlUF+oBlaBOC1IP23Uib7WyIdBmO7BuIP4Jclu
ChxnKeDM2eeHuRcZanPGaAlcasMezMTMr1hziTl5iKjHWa4vCx7w87haPOdlrWFe
b/KVqAR2ZZ6DWLgfpYUI/ns1XVfddfN5Hj9uFcUBvI7ep1ImJYwrQ2D2onAUrB8R
8MNfJXlRCgf1knl2tLkG/f1tcZEZj3fwtTfV4FN+oviuwd9PUwkO1Xe+SWt4kGTY
i7M2f8ZXRIyKW+wejmr5srRzhdpDQmFpGDXS8wC3iNDODm2zwk6c3jL04+MS5LI2
aE/RC1vdk7cF7LAViOuZR9yWH2x18g8jze1qDmfcB4jSC+uaq/ugux8bGSDo+3h1
ReVbnZpmf/TciJgEbftmQTqm4/8AVZHKAFCC7jFfdXds0X5lyBR48qAklBfx3c5f
Gjx5Nb2HnNiCJooy3IqUpAMoPmfTgQE2Wj/BQlSMIzUdN01cr0wsaJYT1zy+XVPO
QhnM/WbJeD7EXMaVAmAAHdbVFODJHPd71wOqH1oMDSx/U7moWtvZDERc8mXsUyus
mO4UltAIjDfBNSLzbw3DDdnooqWPJAuEcVRinIbsO2sPUwKkcJchnRB4byzZ8pc8
SJcokPz2LmRIH9KPZK5ByfjC9tlhjdY1xUnsMULOsp4qRfhgiBR6fzJv9iYMGKn6
6s9qAj/aBtcBSXxCM9lSSD9NRthsBctLa7JGSN1LPi5fVu5GYvMAy+pbtUzJl7Yb
DWPYD8U+iFkyaa2v3gf61bOb0Zl165XC9rKZcyTMoin6RSdI9t4oTOKjqg7oRLcq
2kPchKuj8LFPUx1hw/IuzRIbzTG2Wx6zTnEDWThy3lTLZ4h2wnFRMo8D2wID+yHk
UapgbF71in4eSWrD7c1VFLLZ/S11NRc8tJeX3zAnI3HkdbhxQ/nWBw5uCpjnuqre
DAiLNuHXFVhWivuXBdVuy4t8yCbNhYkwZz7xfkSIanKn3q353EIdI/z+GAtnfL8N
SwnM6oqjccLun4kGDXoUjToVGhoMRdTleVA59l/gslryueUOyABhTYUb4V3EFNdA
IxvQXJOtnh/2tsywfFLj8A+u+AMat5Tn+K8QwP0OMS9pPROZcGOQDahvfIu2iowg
srumt7uaoih88X6IUC9ziy9eCAljCx6bfMz7qLWVl2ckAdD+Xbmv6PAuYPiE74S0
815aBzSue/DwhKOXlTf4la7RdAm+wnS6YXCbWbrIDonT/sThd4rU9fUhc8wWhGHy
jKcmdtvEP2yuuhybkaPdqInBdtPGMOc2ksJdIJd24SLcd6zOYiruPXVyVQBkHr1r
Ngl2eDs2I9uyWlbRpBjNJXLNvwVcSF5XvNhQb4WSXTK9D95k+WKHWR+RveeORBY5
sNVrglXy5zFbAV6Gk2H8G3tA1+LMDOVaiecefs8Xk7vgWDakaPilspEIqqkQuXAl
4m7Dwl+IxL3s0LPMkYTvkWCF+18a2e8FkZ4Je7QuoEryEjwkwP3sMP3Os/2pF39s
cKmW6k/Nenxk1zLNKPxasOOkZkxGhTOexDY37DxiVMVc3NTmNvfkXj4KG+ek5WSK
2ToHr3U05+8ZlT+HJaAZ+9qPBT7+yrucvMTEEBuu0LKo+DdPRr6mIquOl02IJ/6M
fvpxSeaS9R272qKnt3dy8mw0IJpmF5HMZI2R10S/EPH14h0h8FAoqQZdH6hwcu5E
ukKf1v4z8rtEugmyufWgSJX6n5HzQ1BQCt/9uaKfSnB/wVjjXUgGrbiBlbV+P9yY
Ayu/ssolGpL+F/JUgYoip1FXalTSVCVOuSkaBDYoOeXzo+CX2GfJbMB6ii5kosMm
m4EvIVx4gDClZ/S6mX+Izdp1nmvq91VWUnBmeNyb2OhiVccsFemqBllMGJhb4aY0
x136TXbxdyNv6UD4LjeOxP0NFD9pv0JUodl4salXjBI0S4Cax1v+wddn73oaV14K
IpncQsWtLBAFjGHoIGJw3wvz+EL8QfjAiZBb52wiKGZRrXHyd3C326/APYNt/uAb
TF6OMKHvwCckP2IiKzcIJ+Fl9jwhYxB38Ux0oHeHeVpCtwKTQhGKL+EH6fvEcBDj
eFYy0+cycaMDfBP2IlbAF45Bug7MyTz2v3QpDtMWW6yF5uJFoklngs1kQXEHCst9
9oixdqwt1oK/wLO1zYXA1Ito1SdjpyxbK3w89NU/ZUfQuORTETY6jrmQayQ1TgFq
5lV8pGak4l1q5876eg1u/3j5ZPLBfdQh6yZnatuzSQQUOWzcdF5Knu23Vhq0r5YA
sJKC8phuH+EW3E9gHVG79LIgmHSPAl2YMNtuJKDQhBjmSl85Rd1sIuhGD/U/mv2N
DvZRWNTY1Twmhyh32CuiEvculg8LRxk/eSmqnS/V9R7zcz5sJIdBE3OEyjRLFIvz
9Gbxwza7xJU99s7pWN9kkLt4fxrEGdEaw7ULN9NvofgfXmzE6Lq260uDDa2dBbSZ
thMUUUGoxFH2eQboqKHKzIF/jdtD8RXA7e6sEcR6YHn1kVPKaOmD4Rtawvh3srVG
Ed5uJ5jSgytFEVab448UYMHPc7xsgYTSnWPsYPW3VMCmwGMyVnHJ+MdvPQDLyz97
65L+ynhRvKyhmdyQHQ5bGuGVjQLlMeY+4C+cdRoA87lXcNX3LXBbQI1qXP6jqvMd
B92rCN8fiBOiIbE9jm+jJjjz9A6l4IVVtYEeBnae3sJ3oct47E35JN0XikU7qF2o
xDuC1GGXLwUmYI2uOcRHyIs6RgoYb0tqUz6qXuUXBAqrYHkNGYtDeHwjcp3gK17p
nbc4zlrv9oSzPkUkde6+MBmA+a/MVix+9Z76Vb54PVgwBUT5Jo+DewmftQ4MRAr+
K1Ox99Q2P25vZaDzEC0/woaezRhSssOYc5P6rcS/qjRHWtco5+mYu8s1ubFadtbw
MQ0h8IKJ9f44Unv2du/W3WDdMxnqvj6v8FAG0iLYECL9ayegHI+uOGb41LU5cfod
jhPLG45VQ33E/vcPQCYqT9z1DZ67Eav23ciGzM2zSqRzYw5DbIvkrgf5vADvW/1D
Ehdp0Df/2lJXCwo1txNjHbHKS3v9b3uZ9arJORz1g0ZPZ6mFdrmmI/v9YNNoaLfj
2ofml+pE1qUO/soMTzjaU3g6LwAudLPPwSqQXJ+yDhrdjcdq2CoKOcWun224U3lU
tWzceBBf2Ci/AbPjYlWyT2ZkZR+pI3AxR0/cpB0qV98MC85G8awFMBWI2kpWA3jV
kXjHo3ZkwIccCwOI7Gpd1W2xiF6gLnqA2l+1ILU6yiEQ109ebk8TLR3TqUeZ8T8d
R5alOWID8NN6hi4g5Sd9kAf93KYXaVCJzQqL6GMbZXWAD2XhTJQEFgtN+Uv0fjbQ
+PX8nJxVBzDEgdZaoacZ8XcbnCW4PWvIUS4f7WC7O6YjABT5cyLEZr2oU0eyma6C
xJhKWaq8phFlPPMEC+blF9yqzWo4mETnm1DbAmr748id+y1asy4GxU+oVin0uQaZ
aG8hMs939cJh3s6CnDJp+tYjd4Lhx7LABMJGluY7mOOVX7FLxUhzEPZ76g3hzfS5
t6qwKMeAPyawFoESxB4WeYtODsLaJI0vMczebL2aYiriWHk4oBa6kffR158SUi2Y
bMTfdDYsbr1zNsn2f7PcLjML8CCQlWtIJpIxYH278vlIuI1gljHdrDNIaWSBPJlA
G1thSm7670zCklmUSf+S3N9tAvGA0f5srFd7IqfoEsr8L7/hQustTxkMh2Be2qG+
+GmazuTMv0PJyOZUk/IQwebDf5aD6rCniy02qGGYj0z9EeK4K7f9clx1Iszqnpnc
cBwVj/NrQ652yUjfaG2Ol1+pe9aslADQU6VzsQtVfGUxpHlBMxkzdgnDs2mqmfkY
4ZUd98YuggDN9m5anciWlftefd2kiPt2QbZcQ7/q7BBYynSqFuQXXu4T8e05dPPa
L+WD9BKt/NO/Kbw0VLyj5VtNpBbevj1pEWakdZc0mVcBRtVpFlPWD+nlIeGZT+cz
XZoLOQqQQs9tpzKjSdY/LqkpPHWImcrhy8qCjD6xcMLVUBJCM+Plre870kuizsrm
XGU7vzpJX9KGSIcFExr1bygzAhvyPfGJvf7eWg5pEaQmGCpcNoXldrkpxH0fGuVT
zxrOciiDFdFMwVKzNE6sGvJk9kzPnmcSZ0TrCW6XtepAk1lzX3budUtJ2wI1yRCc
gUi8UBdj0F5sSypDZIqVMxkq4/+pBW2UClDkNuxHwIti2D+CY95t1VJnXDmLIiDw
PKvTQ2Dbvwd9n+jPOS7lR5jPx8LvAixspcUVlDH8hk1Jlrsejz+GpOYaWDftyjDC
mBPSIxPyfztTnNSPLyO3o7KC/o2P7AzeH4IXAitDfaagneAyUSxFS5dB3pHRYPuR
Ex6Qb93yx0aPOz1AxIxrUD/wl42pkAJpWeZyZuaW89DoVL9aFK6XYVWUpk9vw711
Cy/EPMPVnnn2E7rS6+Y5TpHHRv4hq5aewljmZbFVNYszY2orx/mkgDxi474jjYPA
ACFnTSGuHhtddO1ny3cogwmiFrIwtC8l5x91AITgwyKmb7TfaG9kA14o9f23F7JA
4asvc8l/wClL4GPRpCSZ6lLofpmA0eIcrigtdMFE/JJe0Y4LymNX/YF3FLpUjgnQ
irE6BslqcP1AEeF5L/B/bWDlaTMd5VjBsP7ev9nsOi8fweoIfzCLgiEUBl04AFlB
h/nBbX8F67ggiBpJcgb+8uH9Hte2ArZaI69dq3butboYDHCmpvW3RGTVCmQfbx1e
ws1mBxm7gVNSLPfD0qGpt/yEQApDCY+nhFhyFrUkWhx0cabtuH57u4xX6mPELmft
BhaA6k43Snm15VxPo9V15oRmBvkYCUl1CHjCY71TUrXu5zNd59ISkTVusSTRzy2m
seF7HkkwrwpqT3SKpY2cZtrowmByer/RpemvT+9TenU8Cg2wQRKwrVlYoVlv6e+a
CwHJK/U5qsNNbMg1IMxFX0lESXvFvkI1P69LrsSS2JZ9gh93rXNI9MLp5SW9j/Cr
kkQHArXbxE1UEzjK/yG7iGCsS/EFqYAMu8a9C0/xT1fEGPmp98XIZv+L6xrmUqSg
stPuqP6slNo9Cm7PUkDipqZlUcZl3QtAbC5PdVcS8qeaOXOrH2GNhjBkwWdko5eA
wpJZQnl9ZQoqczwmr1C1Q8MR3tHiHT4/bo7Y0oN1+ZKq7fwPoaVPBN+yL6/z0Gh7
PkkhopK4DFQwCObjSvRgP+RSmfrrp/miyUxIOK9n2iUqNjAYrGXdvXCHmpA5TJlx
BeT8A6/Dz84nMPUGxuLe3riUCXEc0AaRFnXK4YF8HH6hoJu6X1bwqzBrbcpfOrP0
uMP223btvKrAUaUdFi+DAKbKUO2vf7nRXZ2cQHkBkfIU4XyU+kfsAODn1mlIpbny
1uNLwk4Wjar3fhIJCp3FBmYZWT16kRNjO55GKF6+mt8tbiu6t4C5PojgyAUF06Fj
QiKr7fUs0Fj7vKcGMl80Mf5WzUyBA3nFmOKtuitNG3LEsrBl3/vmjGQnw2pygylN
AdL98hXDIXYkvarvwQzDOVSgvUBN88Xp2RLBAeJFRIAOl95BRvDg7R72iTll/o32
8WLE5BPtwrY/hUuOBWaQzdTOci+2vQq8AuAKAKTCLUiUA1H0i6yKW8H1S1b9Tiur
QGHCuxOM5dPGXgwAfTtLGQccvUNAxHk6xU6fOLAwzbocv8wKC6POPiRlg0csd4by
8tmhskdB3DbPgVd9rs+wgf1oQeuxKROJxBD0d8t8XXWDMl3brW2DtJkasSxLOQyo
Z1P6rs0Mru9Po5Myz5GyGeHLSO9nCshTDpxH6dahoeRkdlZqt/dYWiZIoqy5rkfm
rI7bq7NGm8sbWTrbUEjPGSbkcY/I5yzouNgsnqU46szqPVzx0tCe8vLCUe2/E5io
xjGEgOZvFMj5N+WNLqBEyiYM3sVFuNWcwv5SiSu5nU1YTUAHktJD894tOLBsqRk+
xQtQNyIIGDLKdpaAN4xYusUpLrpQEAWRXWG7UIsCcXQLaN0YlHNtfWUVEkvx7+id
bf7lEd4GQLspNfN4aK+2Dn0fXRUi+ozD9zRxk88CYoEvusWV8PJxP9atFuPAVDCN
eMyK0oieZMUGQdDDdZ7c4pvWmPbK7XEqiaIdfU4f332STSiRm+W35C3uUce+4e8C
CpgxUAv65yKZQT0xYDGznd3+D8xjj0VKkI4rUN7nmsZv2hyDMvRRhV5m4BTsn0EY
ilxMWMdJo9P50uchfdxrVpAcxgS4uXcxOItB1JPn6SS2DVaMsvRjHYoD5NQik5WR
jNr1jQV+lQTD7bJXijBatvUu5NNnwG+qV2ESTFfxOS/A0JrBPiFDhH1Gz3vnM1ww
cZjyr845RYm3zYBso9Q1KhAbMCbFBkpy8yLctUPEhhuFCPiPteeym5CCmJQe6Fhg
AisPX79s52ZgXTTTsN+I/vhlod/4Ea0eLTNhItYhVJwv4ICe7ktKCfmtNZ8hUA+8
WyaL2geVJ0VZaftDOg7WGUbhgB5JOZrjKB6fjp7f/yxWya3EXIgwpHRlumwuu3/k
V0yAeKanlEAr0QqM04bCK7xG/rolXyhDESB67NfbDM4d8mqdjSteE5OIY2/v2r3D
QtrS1csyreH1qHmtE9T2HvzZU79XzULOFj6QH0sxqEzottI4nP6QyWBpiU19mi93
2DkmFfdy7uLSOWppw61PzFO5R3c0xO/7eYXBKw2fZymYTCeWgVigJWr309D2BDJQ
0zDmG2qTLZ4W4PBZ1NdtPRPUQ/E2Zkpun+d6NzTzeYV+qYfgl5j12FYKfi16t0xr
8faW34KseDdlKJyldbY+rgam/umAIdT/QftNyWXrGeBikqXZZ+w21CkzQ2yGeIIV
Tz5QYoLHtbaLJRiPgiUcXLPrjYo1w15TljJOTrxQGGKMJsZz4xv1GjvtimJDX5Ga
g3/3mrF9pdVkZe6CEgMroq/+/85565/AMfZd8++87hyoyTWvX2A4yc6aNh9nXFhr
ezFOb//xONaXMm6LS0EIi/xrHRKv/erGeljCjVt2CBAlc4MgeJ3sKCkuLxGM93oY
Lkio5py8sH1ojTt1BUeJyWlwULtRBHlBpfVYVFclaEAxCUoFMVypJRKS5/OmxGvx
xdpo9hHHA8kJo+/ylyPycSOJrxBkuQDIm2QNRWFe0e4INONIiHIwC1+dsxotu4+b
vYpyhmHCYTQf9uIKBVdOi8vHxPsLIv0pivuOijEuSOTw2/Ptf3YLLxX+ddAoeZCp
+uRdgvOgC5HNJszoEhB5rOVr+CltjJZGDn76mg1SWXhBCrS3Rg3Lujus2sLNOENn
SwjPDBEKyL+CBdjDTehNjVbJSSXfQLyuNNghUYaIGfdI3jCHbnIjRBw73OlGKJpS
BnVVgLcloAdUXevIcjf2LLgO/IgHW8I3pjnqgiJt1E0PUCc+p16GEdnOS5gb0ry4
p0aClH9RwZK8fl7tHiKPwvzFv7IV+j2CGyfUhGIPX9YCSvcJGs333pWA7VxRKVcu
2gSxL3kQQGzLpaxmNpwRLWcMw9A/BBb5L70DeCmjj4mzRa2Uuitxm76OUbQ3tFX8
BR9NWtUmTNClgY596r1dZG1WlPlxIR5T8KRh8LzfgNG28Pw96W7yVqFuEVKhVtGF
VqPmoh9GRrl+ZPj91TRZH0AcaUELGhnvbu/OO+v6Hptu2wYX6x9+mWhVAbbq16d/
dtwxIxbikWRCzdmu5UxeCyMKchCpbrLRK9bvl/wHBg7vARhe649slxN1P+RkpT6H
s18IPz/o1aSOPSbHTu+Y07M5bPv0HAfkd/W5MnYZOczbywzxD65TMtqnrW8rOzU0
aDa5SMHZZki2XRtCnf/2VofscmgwdcC2xabBXQ9GMh9F2kCcyRJyCc4SEpVjMSxc
C1WK56tArQEZ8ImqLxGa+cy1Si5o0591IineSfu/GhGqFl/88EXGG5MJumr6p9N8
0cF57feLBWNnmG/06z6bOYYQ6hWWzZuUuf00qbMCQHEwMuKKMq4BF/dUMatlCddh
gIFtCRPFbnlhJiB1JajLA2/hELHjyefW8YGyN8rXGU9VQ6Q3Wq/wfd2EG/Hxqa3V
kRqoxgKc71tFXQ2Qzqmzw35BukE0ka4bEBLnu1I/dNZ4CePxeyT1k50whRxILHHG
fbScwYp1FeU4Wp+GKlBh0vibNMaiv+WEDl/EO6OPGuIOuuFJt0pwOw+l0B07wfdy
BPzga6zOcoR1JOC+sTf0UmNbiLf2UdQzNVaj1Z0NRYeCQyn22JKgcvrCS8BUrF7B
v2Y5UaQ/KDHRJHk1SVe/L+g8ZIxL2cp+dOERz8cBRrtRVjPirfnWK039IZguiGpo
zj+NPwXE+nQjsSpw2H8nZ4bHSFF+gM2aNmBu+rnWcNh8uvzGN09Spl0CVPFPsT79
rblMlWNxn7hwXjxbTre+u90iBeF4vc4wskDX9FwCRr3mbsecGbXyD0cJUhQe2M/b
3lW/hPrOESrvVQwz/RiqPFQhd3C3ZU0xezjwj3xMgjc5w0ANUstMEMKCzjNrr6k/
jGZrikm4IGttr2TQyivd3HIyljgf+XMdy4MuP+8tbEwbmBpXpHVpE/SyuEG+Z7Ry
PdQCkyFlCTMu9fCULkGujYoG+RVLCeTpGfTp0wXDV/8quHj0CLYeeGjbgJLph7PV
xoJVfC1EX5R87EzPbkg52JuqNx3QqB7+XkeUmcKfQ49Uv51W08dhNO1vfeZafVBp
6rVgeRLDC4VkUTJf+tGz8G3WBga5zwB5PricD+gAcdLyfcxArInYS9VQpVNZiD+5
CKtRTFRh4cltH9wYajgAxhpyOjY0pXIqpo0LObGfIkPqcNMlJ2jtE9cmsCGykMvU
LCnoJovc4NrJvb8M+clhn4r6f/1Or5kH0aY750p5eG6fifI00gsUZdVEXtP2pM6k
Fq23Lz0YDbKrghHLqQcdai7Ypo8yxj+xDd0qMIK4uMZgoRdaqycHqGYVCVKz+dkh
sakcfLKwmSZyZ9bpge/H64DjQMRInwm6QGmw71gepyMSMhxORPu5sG7KJEOIKFdg
w4r0j+VgEfTrzbb35czAMC8aDUJHQMyi9+J6Iaxt/CPJgERdi9iWwxoEdo8WHVme
P7F+TSMfc9n75K+KmYjtuFtgG4LF8UCcDYwN4vV+meOuDIl+3MYso0hdiHpoy6SQ
0YusW0SZFlErk9UlMrMgruHupinpo/QS1wzG/Wwiav5FGL6WYES1BEwbDDjuvKOg
YFA7kd+B5nn69occ0DyEBY0jdoDgoBA95MxLAYPg/bXkAOv43yTTachFj8hRFMhf
Ve3p0RGVdjJDH7Eu7EXUMqLbOBbQgFBzn/vv8HHv5TPqwo5d2bqlJkKhyraQ9T+J
Ft0MGV8WqG388+2eIOxj2MjpqMz7DrPOz0kPq6cGib3HaluglXmSgvHHW0baGuBq
YHtLwY4grNRuarbpJR+UPNX4oEaYZxYlZdFtvrArZipjZ5M5meawOfCLVsJPgr7B
vImjCNyjEhxUps7F5E71RfkWYfVfSvXLzjQLWsMTx0fsXMkYSsZx6407bfPdcS2s
arQg5uuVj2zvZ58txnjielyYxF40j1Ehs2bKrLfmsIvo6OE2ckvXq/ltUvTQfghP
2hvVPg52lDcQGAlMjxz355FR35DRPW4ebHy7Ih3Nmtl4u0zZNGVXwk/nHEJhk0fS
3oAzky9yfZCftH9rsqsVV8nVbKf5IfuedpIdn8dsZTaj7sV9rLda4bUs3xOHOyxI
IG5vyk6yg3j1u/v0MdwrgALifi0I9oHdocevDwwhwtzc4/0KHKyChVSUw6gscb6D
TZDcl5GOzP+33UtAmXfoRPNIxFFcDC12XZa3WerZVMXeMWR0MWEhDq3I+gN2j8ml
Ga9XlzMVD7rYBlneXFA9Al0mKiXREurAdHQWcLs9WkWD1m/44gBZi+Hvu/hEtNBc
JSAcCYkyE9cQypngROqv/QzhSkRRwpRzf36j0bqEfbjJgVG3xxcNDiiPVgpDdOZN
Yz1fsv/UJCl1G3SaQEglOW4Qp8AdWJWwwiPGs10Qeo/JzNsB4l4FNZrUUVWxuzm9
CpHiTzJKVu7SExuep0hwZtit6EOtvJ2ISHlLsQH3Bqan9mHSYi2LC/GjGUURoMf2
89uqXF4oQuddyPPVlw4JHe6QyiXXdwv/h8Zq8knnj0ihf76ZpsdqQojy8qlJITdR
78ox60W0tx72fJFG4GJA3m6ihEtbIAf3+G3qhYtN8tIxELIDJfsVj//CKl1ZzGG/
YVJWNlpbfRKzsljF5FT9JGbD5hgabdPHFou5zHxpfDvp573VJTYLffXXDybFI+vy
snW4y4KD9qpSD/oE+KE0om73frJ6INOoln0t2lKCmPa4NQw0NEnXuwq7m6SkR4E3
yE4MC0jzJ9Y6eXa8nDU07klDIwwK0xn0Y4a1eyJIP6KJ9iSyKmEo7qOnQRVmlnAa
d/heqv08ATuH9P/SK+0g+uBnbeDVwIB3syTnXHRg9D59SFs5vs1zToFL+UORydlp
pg2IJ1B3z2O6+AdTBIwc4jdiBGWU2LKoWEpAPJ/eG32iPUxmNBA5pPfk2yWZqD2H
Lx8zFsk8nyDjodZe0d38OcyA6GnwGgJRnkVWc55mBIWRZ6HPN0kQqst2n7K9lL96
1+HSKQOngLpBx3rP3cqLMRmjcnFkoScE4KAA57N3GeAY3+MZfXn2N/ysjARyb70x
kGzXXCSefjEOJzrJFmFooCUYvGZ6xKLjztY8I6Wo7/DOKlRxsYqoKLn/1nFgHkhJ
D7zvvf+ujmLqiqo7LnJ4CvdnSkCCP/Xg1nZA0O8d9YEuw28Yeq+jD7BEyHLQI2vd
6K+p0/M6wBqG9ToTvWEPxBewj4DCy3xQ0SVkA/5MXkmU30JU2gyEMEVmjfNCZJqu
nHeMt52d8bIBHNbA2NozqV4sWk8sUHhWvOFCwLS7SggosLvDrEtMleeAxdKNBYBY
2L+7fhnxQcTh7I6B8FIsnnu5xmbNoZn/kDIADBuaA74MtkqnuoUU5pnpZ821/d8T
wXQLmLRJx54jPIKpE27lnmVXW/IzbErbb3ChItllz7V1hWsjXHfLxTke8oo6hnda
QTiX5mZRekXxxqQsMD0ZvVgDtrOQAvYT9WLICuop/sF4kVRW9b1qGwHQfT6Loyvd
baDAJj0kpdxwKP0TEH7FQk747nrRnFdgKaA3UxWj/0qv1+acCPWtwIBavF5+mb24
FYcwHiBwjFgbhWiPizMTsP+q4kSRgy0FrjETPUOwdsIKUOxu6yMMkKhZSoOK5uOx
Yk/UKUjXgFTU8j91Ye/0xcorRJCUKJczxld4wWptyLrctO6PNZxJOz+qJp+J5/fD
VooQqIJoDvRWI/Rx/lJpwATXJIkFcIJNbh7KLLnf1vNXVwmLBr1PX0CwDdTymT23
uuFIngCsPMjxoTwzgeO3QRvwz4fNQjBmZ6A3GkFSux0BCrbw07RGTlIwIz/TzWt4
1qbJ4y4uo30icmYlgEI6+GMCe90NFOhrEoQD8023Td8RGLMp7fBkIyJiHXJgZG9A
M+PQJbzeOOFiMn6BswQbvdiaZx8plvdnS5ZMSkZSedqbqeImNk+j7tcbrAo4R0Eg
ZPK1bLhKG/VL0aKFqqTDhJdm5AKDp9HZ0bxvHtMIZlbrV37YPws9SOhDnotgJw6w
qofgTAJcGlIGETnbGORsx31DfseHBwkTxfFPqCJ3T1T7XSd7RXQ7dYZur9NljgV5
f47BEQIlO5TdViPErVjJiPcDj4K+vbFXNX3b8fWvwXWwmzBRD7hnm9/wXFeHtWHt
YWC/iZNsNPEw+U9h4vcWDOpj2N81JtszpXNevIpofHfjYN7I7tAHXRR9aTH6Hek+
1vao1PlebVZlfx8qmapgxcHR2AToOOCN8RgiIcJpc5w4EWihe0xVVb9vBtIV/N4z
EpstQXnQ5ml1ssAZU/q4lxPDMDlZ8CgNs42lt8ViVR0e/Yw96fdTM6SWcFjV8U1p
6xmiRim69zxKdK/IspUfzsUl1mYGKrek5mObpx2/ru47N6Yg/EJGnk3LNcEgP/g4
4A7/5avCl47XantPOZ9aE6TGWjafVB+vZZ6p/icZAQZhxM55Twk6V9f6hCRet0Sf
MqCSfzM8vgvNpb5tCFS3kUNJRLlWsHYO4NXfuR33k/A4HpWkcH76SQ2I3J/MnoI3
MCROBq4Ij5EI38XhZa+J0cY58FWDPP+IywjjscF7eUf+8hDxSxSQpj+A2oADp8ML
pTjNnYL+zLgLtuDcIQfj/4dKhm5gCm4Akk8fW6aBtCBX4O8eKL/M0KYZBv66BZyp
tF0v4xbwI923aWInG5k0xY0xPjmsFuWxCwQ5kJhZFKLJ+LqEkJGbGcgrFgfQ99x8
GyEHBEcJ9mfBYf5pMMm89diT8QWym8UnmWlFDX3e7iBiFBYI5Z4dUXEljVJEKMnB
5Vr7XY3iouH+GpIVxdul4bjDVC+h49/F/q0ata/unM1+2Rt89TDE3MaFa1G4W2fe
bq4SKn0Y3rdpkAfpEvYYkJjePqNI1dEyY+nvzkgTtUoQfkrD4zGEkakgMZVQyOOr
MicSmc3qS48vMaNjD0wKxWSrnFmhz2lM2+Yh4AsAQdjtH7zbF94VG+kYdN230vbK
rX/yxBI9zbnnA9VhKGYNvvrB1z/7zy6N9VJPItBnHFGO3LdB4VNxBj0UAlEtNAry
ZOIUJnSyszVQ7li2Kjw/ikD+lGctCckKFdxbmCFJua1v1FW0gKraxTXE5CMFmF0h
A0pS4AHviSCi4gpjymiCD+mHi2mtJT57DzYyrY5gLKrIIKkxRwCX7tN84u3P2Zqd
dowbMuFS5uptIgXPqYDFKz30Vsax6A0vg45Bv5sPF5JcBP8odiqQB4PCx/q3+AIS
7ll6OH7L1CPdjlrFQhi4QrfwLKroDJB7+nr2ZNnW9oTfri4OMKckAzljtFiO2z87
5N6k+4xxp06LO4NMPlNTrT7zUWLmsXcGFzGur+f6tglf0xOMKYgqUkJ3w7vpiL07
6N/j3x1ke6fi6ML4BShCLwb0CHMd/9UwJ4qs0sQc3DjCB95mb2vLA5m6HOKaEbP6
j7bPFaPou79vmeQUgpVn5dolH79gpXB4TqfQKWJ4mu0spt8zpVTYM551dC6mlJ1e
Cs3skeHJlGEcD+hH+OIRnPe3//XRMRqS69vR6gE2tr6wYiqNinjKfK+YePvJI6lM
I9y2VQjRlFH+7uTrJZxVnyfQxlIfkfHXzO+MbozHlqb1+6cbJHK6MkM6J8fsdvIb
v+IhPsPzMir1VahixnHf3aRfggV5w0hJBRW9AGNWh8keXD6zWYeksCZpYeCMUUDG
c5ihamCN8NeRMUTwFYqjhN3razAQhpTFIS/ImtwtABFpfLbYY3nlbjz0StOh2tG5
2VCC9apseF0M/o1VFawHn4fMNqKEQSgXq4NrBiXiZacOge9Z26TZ1CIf0zuO6/H7
k4X8f6xvSvzFB6uhBMKWwyKtZQXuNlIk7jDXc0cMT6Urot6arUIXyWCCe93ePD54
97QyMcgy1RqJ/jkAdH37XOGkKvkn6nfo73rUOCbsVuIwNZysI5jpfmm/GQNBthwI
Nnz9Ni1f9PrukYO72SYwRQSgFuv+v2FAwBDyQ48P/N26aWAzleVJ87kVvI2q4eMk
2sfa4SUrHiRLHNBOXMULn65l3dAh3fvchvRB2mCr93aab0XDeMCcpolzzB3bgBVj
rniY3cKlzAHqfX405T5ZcMrBZRBIjm5xJyQZwUq98JjV+vgZyKZMzUKX5jMbJC3w
Xn4DM4sYinp88dAI1bGvbJElHJXp+Y5/az3BzHzvAwTSF2nAhRRlApbj+fKNGaFa
7947JM0jL23aqRhnaWYkJk+J4S1byvyadbSRKMuFYtDKOuGpkE9C3mJPqU3HpL3H
3x/Qy+jv9FJbA72NDev0TCC+lsjljqdrwfbNkQagybGyVsoBPYgr7Rz0KSYs8q/3
41v8tsr8U2oQCtnlrkJKEB8FCyM4jsIGax8wnNwSZ5U99X5Lfzs241fc0ATtLvbM
h5g0DmY5xgzAx24BicVDulyUsUxxjv+jAWD2LJV5fotDjkyRNSzVaiurpmdIFXXO
Et9dSj7JFcb/0PlhC8cBJ/T2KJStBW7u2DRonZRHBaGVlNv2Ew0FeUy8vsV1nh3V
VN3E5UPZjX8yvQ+w+Dw+6yr7v9paswZ7diPdbO/ZsUp6hmamc8fIV6sdu33eJI7e
CesiA9HxtjZU72wboCNqjYz4i78+pfT8NZnoTUUNOXtxc1LqTgFtE+qzodaZCPwO
/YGwKtT/V0U5IrQDji6QWJKst1BZVnumlF4GKz+S1MKde5QpcEQppR9Xi8nb+Wx1
f9PidnuJik/o4+k1fHfYyPyYrl7AImVgGGqdEafIiJCq2ecn0UOKQmPtJNHHzRH7
XuXiN2KIYIYKTByoxKfgHm/sroWE/XJVEsWQ5XsbkSOrsGLmcrw3lJ8piGrejf16
fj8pCqTUvbqtYDO0o/Huf54HKU75h/DJe9fvmPZyUVN07pj2kJa/jx33xhedxikA
nGDBl/IuOlUS8jRWrSbIP83a777yYKP100vj7YpydINahVro9KEbV47YJRKRLTld
iCPjh6BA/5bBD2C4S93m8q/NWvnFdRqyDSPyQh1Vrh3JByV4m1YfzwEoe2ZG39P2
JISGigKCKx2ZSg+QQ7BWgW+iJF/2eiEAKV4d26/KByNh8LwIk7dfSwB6S41AJ7nv
q5CU/FyzVR06Bl6Wodzd/H/rJyUGeciXFI1r11Dq/wCj11zQVD1pnNX+dBduVhqz
MXjzVDFOq/J2Bf2iYaLFV4TOtGrRLiDX4NYLs+4hXL5Fr+qVgpr8b8YdftGoWrd3
HIWqtQEt8nYTpf1MdHKCDd//0wvF5oBtRqIF9pWd71+Ic8Yn05LvpY3rpR9sal5Q
ZSlerqvwIzWszpb3XMl8HQoWB8jYwx2F6AtdNO68KLaH3y0y7f/As8u7MvmLzMmQ
k6mHUedVo8mgy/I0txsPzXKwN7PgmPj4UD/eHgHQALhXGMGumOteUQsb6tLycHVl
oerW3mRagKJZ9587g4JIpHnum43AaSIOWApI72VwSCr84vkrz0TBoTUkdCC+r+jD
/cy0Gp4Te3wsMd849SdQBu4yJfWo7TZZ0VDBT3XH8WJTlrd1EsQF5itUHJ7e37sf
Ioc3HpCY8Ur9clTX+lL9jgNvJNGD6L+i1m30+vc92OW2qyeLZDEYZRrB2BHPFvLY
UrgFjwoxI/A1gqZLhGBgcxWZZovWeeI2Tq3HHk9ZhDKXM4ggqEmzOktHLDubzyEx
xYTQnkBqA3Z02ZOntkYKHPpdq7zBJC1PjH7zF1NKqWnQiLJdB3KcOYkC+EDOO5sF
pSeAyQSFqFz3KmCKJ1PSUZYGt9KN9Uq43YWq2h3DOAgdGq+MBdCEdJt1k9VteULy
c8Pkg9SkSWUJ95LtdzlrU9/LDLrpxsTgOZSw3TL4EFkTN/g3Ugd+5rU4diRtFqWY
furzL/4r6yp4xDEmlmzZYknRMUgnMIH+qFglqOrzvhwCdmlmDFUVNIIZ52LgaPU7
7CK5pCwRGDI/g9e4+pHjMvF/uslilrskK758CBiE4uwPhAU39cDi2VAEKG/Y9hjh
flGGPyPRnS0te/TtZA3j+2wMv23IZ7npzPKxXearHUitLqsEHPSwXuyNk8gftGaX
CRDIsnuK3PnfgvD9xyHaRoggKAEa4xl/Hg9EvdmuWtvz6PhbkggcKcRVgjt0RuT5
oh0mU3iU+yRCn+AfIXlD/qPOBUn6gV99ntnYqOYrOBqHaxz3enjLL5yrey055c0I
ocXiUN1VjpQjLqISeRto0yGgHt1ktE4oMG5qVrwK7gJ+umdK/fovDsyCOg6kfKeb
sZsLUdKdhnZWlRLNobV660KHOu1GLfPxStKLVjoBj+bbnvZ2m+Zue5pNYzDrq+9s
AKrncZBiyYLTvrvvY0dfVThOWy/vQ0/SP34SWSZiu/b/0LExcouoKgk24lFX3EXC
oy+suMGAg7jFu13/MAIQJ5qhDeIxSCqDs7EH/zFAxXYu+0GO9HfCGQdEQR/KymIa
Q9uO0C1oajgjViiEdklSkMIx5ooBqnW2iM6yTf4mU91ZKsaHOHNUaRZqCXwqxu1w
pWl+kx985EVpFpnOhBv0ivmd/iw7bdDTQV8Xm6lT95CcgvEJAx7YFVtCTmV6LIIQ
aq7COEQbEC6qsy/gW1vvm4kLdCb8LP0y7LQLI4QGh/SPQjH2UiTTpoJV1Ohw+jQk
0p+ulelPo3uod6PLipKgzHACy8TCZ13OO0krz16sT3Y7aQ80XJMoHioL+EGXRheN
irr5FkbbndlN+j/szE3PEH3BtynT1DCG0eLoTritus5Xuu3MoOjGMoiiQdy6ijcA
VBhKHRY00UQK2TSzQbwVwSOhNY290u3tOcDka+fs27ZPguz0bPNHeHA0zTqCF/5b
8OMcnyLT89m5QtXWHOTqSlWMimKgGL5dz9/EbIu1eXVkQEVclpKKGFPksrlpDOOn
TSez+Zr4FVSuOtJ/yFP5QJSpwCcd1+ONlGLswENXnHN2ChWRJxj6yACVrw/6qVt7
ivR/hgaLRYfyr9HXM9Cgb6mtFGl9jwGPpsgrjkxcDFcCjiVlNaKVjBGrTl6D1QMB
2NwRPex7qWBTI028FckCZeMEIEXAHtnXJ0gSY8zCoyY3aaqGZU5TKaE1n3GTtSOC
s2jQ2MFtRupRKyAOEWpJe8VV5Jf534AXoUcfIZNYiSuU8KYYGMAnFI5FnvBL8VoO
5efYeaCVJU7yY62BlHDysl5eOa5coBi7dY1lc5VCjy8rTFpHkYk6yeKuMs7XI5/9
GhQNicFLvMJDmXLYVsNs0HLykedOgekLSIYGE36/9UYC5BtA/rA8Se+fIlsGsZZL
XAMdepylOpkT1uYIwEZdBZhMsYe7NMDkDxAUyjQv1rJdIeooQmNqtTRbX88fV6Gf
2PM1rTJLXY5kW/SQ4gM3BWKtN11R1jnbDd1zdrsBcar9YVNzdF9BQ028FAgBcoi2
+c9VwSOr1Rgp1bF5wdqXIkB+pFJG9u13EPfM9y+Tk9ExF0sPL4KGNWOtcitXllsu
9DcnS9NxDNOmocczXBk8h68LeLAw20ZgwmVIe+YATKnWOLaq2GARfYgI6r7HACw2
0BdENB0/g9K8tm88t1XFfIjzmBtCDdGRWv2Gcw97xdNezyJKBHOXb5nx8VpdqliW
2XN7jKQl5BJZhuLzVJhjMcrM0ciujKBPZX6y01sB0c7hGUThTJ/gEfV3tCS/uxw6
VVlopHT9ypB0UxAs36PcMuAjME80iNUMeDw3MXNEFNlsiuOrfQmrmz4KN2DUNSR8
v+FW7SA792+43aDGYoER2uCY8Kju0XrBoyW0VH+b5Hd4gUtouStoAAu4VM/3LX4p
zE8QexklUS0JdHdg8CQvk19OBcn5q5vKSfiBjlu79sKBBhjmd3m3WQutvz11ow4y
KM2lu9jL1RnJZsQw99gT/tcoA/u++uU7Q1JZ429A9agUWDxdqF+qHK5snSDNGMkp
PPwW2rWjSzPuEpmjxltk0pbkO01pupXYeSqCZStyQxTCceHCQ4Ud0HZCJOkeULsB
ZFTr2YO2q8ROd2tbOjsYlthPqnaKzvkNhA7SnBWnFFMJjqWW41bdcFDfvm1Ugukh
6YBG5b3LRqXWMbWY8xXTOjxKmXpRgmltw7yClNKQw8cQ+SeoyAqQSshLrrOGyQPC
Lw+yYEI5BIbpA6SI60zNSsTZP8bBcDDkdc+Jm9R7H6V/rH4bdrm1auW1WSUnLufa
CgmRhPxQ1HFkf9bXN50i9o9Vye129JspKHaLHyXNxOfGv0mYjvszPGUEGWEu10c0
uvhpuTRCSGHwAxOAR6EdI76N+sjzYHa0AvJBJbBMCnS06txC/aImopLpOFVwyRnE
xQn86sV2MXw0Ws04wtLmZDv/90rk3epDkQ5NVZwlPQYn84hBL8MATdydZO5j2V9H
BdUWnZQt3pbR3MWdDXRP5kye+6oJuBwGWvVKEt9/MqaeC/hthP8qx/7/H6pFDUiO
oMuwK5MCK1w8iE43tJYmOXaLd0EwbBWFGnuttu+bFvrtoolDLDi+u0MOqWQ6fhlM
8FzkW3NWhYRdvSpYRpu9KNTN0km4b5tLmA7plRlht+dA+7yXmgioqS/9r/FB8KO3
GLC7/q+Ce4AkjIa8xMUDCF/Df8Zt9RebKtNJ8hZJrh6jiM9fR+Os+vEIM57OOm/5
pnlpL0F5o9t/LY9snzbU681ufJ47TDYiaCJhx5xcWdST65SKshrqoZB8wz1hArVf
Jn6/tnLePNYfm5xv4oo679GrnZ6dTaZg5BOPDdh1bFngVK8aXBVZTMHVRRsEvO25
/QNaZXadDnCW82iE4iqkdo/1/PK7vplB7pMTZAZ++XWm7f/9j0a6Y69riFPvIM64
PaUAbpethOL+bk8xLun7Sznh3aHQlgWKnptizZA1oPZrLXAY5cdHltJ6b91gYarl
FK04A5k3Iwwkb0lrC6VUL0elD4dnk5NPF94Zq5nCztsezFukygQp9EyDXll9Im6E
vjs5N+zMr9aUdqeFxtzZoUxnU+zWJb7hXhy36qoa91U+lf6Cm7dma6b2o2Lx1xqQ
FXfU7SyFH2Y4VOlxwCBnOtNbu6Vpq2hfjkIWZqlFCjUJ2U4w/OLC/7EvyzWxD8D4
cMNEE1v5HelOvM03tVohWDYGD/5urA8R2NXdleHFvCJhHr89vpw3/ZGI7c1uDlFh
94DJYJIu/uVibSU2aId53xRbqEficDj1enjPshySe0Db9CJlLffiRFOxnSquCnQe
Qkn8Hx52sql58j6izIcnABiGyB5e/AgNRcp/RtlEljQoLgctAnQXzL/2fuu9wA3Z
NGPGZuY0IANh94mul7D2/1H7oL4bhFKt47XOgm/r69cfJ8+BPb94qEAPphIWkKa1
uwKezb2EOfokfHqXhrbOiAM3/bwSS31ULrlzkSnNk/9MCO7Bf3BUrE0YYOU4oRYS
JKF5jk3Os+zlBWIP17Da5ZxR2XVzo7dRQYFODRZ0YTmwWGAXbnzsJ+89rPslSVnl
93JfHO0L4EjehQ+STGR/V/SMrW1teVwSIso/HoQbFO8x1rEff7n6xWc00JL2CUWZ
j2tz5BX/NY9Ldkr/KDOElYx2id1bz+n4cAu5RUEBcGzI6aLWaTuXmRYKscEmqnkC
Vj7DlPst8665FJcUOU7Z9Ss77yqnvpxluuCWOx8XuT0zfyAw4oT/9gR7ch2GB4Pn
DXgCGvEzdy6BBM2kUZtUH7Kr5xscVVAwpuK6JFcC8hTfnJCKlqk64dpEy3k3+YX0
qUgvnPuKPnnLxdKi8xRpkm8XCyZWoKkbohVNlmuboEkxMrIk0nBosXsEYolZMJHv
jIKtxUP3F6tmgZ6TyEGwmJIJ9reqYbdOiUDtDSKcVc4eQtGi7NWuE+w3pw+5o9W3
Ke2IYmrOKYpaYp4sKbYWa4bKwIL0YSJm46gHJbKQDrCSWgWaWKeClNa62dHpUFQb
r/sMdWNi38+V2axuuTHi+SVoTg3ef3LvYPTf10OrZ3eOd0FN7ByhRllxytYWBpSn
VYGlIVDU0Ub/rd0Fq1cr/kvVs5FRTnww+02qkSxO+zprWNq0NxGD0p4a2hcbfMhl
iXAS0TkqwDTfwE04FT7NwDRO+g7VA2vD72LOEIAKXgL1N3C7EhUsR773793MU9xc
0fhSXAXVWJ8ejK5BoqxqOAFOcNif2a2o+6xHjS15vJ9YyINMBYRVCQ2oNpfud+it
qj10eHfYR8KP2kc5dMs+pz7Onyuoyf66besEYbySWoemGSYgFVDtAl8m8+aTuksN
LlOwg5XCRLKSJSQecPnzcHhu4iIvIpFXreOyNT/21JZicXDld0frgMdHfT8IfTMC
TBGwojaUtBMG6Ak7+q8xNG300S8As2/Dw0ftPbxsHTMQ9u2Xx+s9Axoi4uRNtzzD
O4kui0CMIuBElpPO9MAJSbS8rSE0NF92yslozuDLgRz+UTVqEpkMLCHXbj79MxGV
JNRhEcPOEs5LBdoAp2PXMhP92IamcIky85KePnzpjH8VA+B2RFHUDhboUk7sDH2L
x1/04sNFSWqCFCRK+pUTHTWGirBgAdcgKrSxw3J/Lc9h0Paw7RxTKXvQAaIVwlxW
LNJN/ggCrvmm8GTACBkACVbBgFCthyqEqxB+RZE113PVttT+p3naM8IBBQKxXAt1
S1bFE7iCgK+lRCjDO0ZYB8N3vgEnesafoJ1fNU06lI8KfYjxoTEjQlR6j8q9Rb5G
5uhR24Zl5jSxisy1fF0F6eiC/+Q+e+FcYuxHs+Q1r+xRwGMP2C+AS8V6KVEo/+PN
dJxlS/yDYQD2raplJEd3tVrwBcq8q+ro52CkXUuUGcN7F6LZyt1OrUegrwG7b2Hi
CANtqbeafaY5aabKD+daEdlXJLJDOKbO+bfNKRAqZ3CNyq+FE59b0MiHg8yT6Z8H
pocRMACrEXUJFnOkUy+l01/tv8dJG4s0lAB96QQaxCkdAAQnM/xzqAGPmJdC36Pp
RQKQgNcjaIEL3WnECHhusYhNlKpPuRJYz0+09mLFH4DkknZihuUgWBD7XQUGBIM8
TAWDbydg3fNutbz7LzyUdSxy2eEBjYARu2FxAgjfQJkqLZnkGV6GZ6+jq6uZv8jr
uxBcB10yPxa9N4UYN0+LxVJn4j9uP0TWTTipzmX/gE6B/bgav5o9SgOQ7hPs/Pzt
xEbpnc/h29/5Tako1eXTGs9kFzfh5f5bEWF08aT/GuJJdrYljh2Y4uIIpgwJETSF
KYRRiO+1B/GnywnlUUAUyPOk1Xn+rQl3ahKQUj8vTsKNnVh+zT/9+b/hwMI3cFDo
03CxSpl4kFnUDCNEdhWG3lfLzIgen1LEEAqU+l4aWcEZw+6Fh+SfZVDleWhmw3f4
z/Opw30wbrFIqU55lUSOlhuvYRJ1XMRm994faqo6oqLukhAhFYME8A6edt5LJ32y
SsJMup7dCOG5OY4uHJ5J55LXs/ROW21BXZNPezW+avkP/lpJmVCcr0Aw/GUvx0zM
2Fc6JW3RbciGkx/qSJ8E92Z2/fnMAQQYrKUi08nJzw7VVPAMf/zbSanwuEu/TS54
oP7ERoqqFD739JZWfarRQxE3lfC4ieH39xnal7+/o+S/Frz08Jd5ZFlKrv3PUNRD
o69p9wPYK/VeVDLrqac+cGnFZDAzxomP5bEnxYXCWaMe72jWdWHzw3/qJ0la6fyV
R17tvBvCwc3JRsGv9HNf73hG8osjW4dAwW3De4GrFnKEE5ElfU4sQ1d3QxBhAWIS
dOlQnGQj++z43Yv/SN0WZvRRZdolnnV5CMhYKp1sDMugJEQcjYVunK5IKuvA9sRh
FqEmsik0aY2XgN8W62fSmwt3Hf+d+gEDzHueCqMGD8JYbO1mzwIRobd+sqXt2tnq
twzvD+iBpVI8ocNvlA1D7TN8V+7V/uJSb26Ix4Xao8royDkJjkvt4XnnHwYzBGnd
cxmOgSKFFu7cXKZy0JxIybEtfE/AegtNMJtECuonwROBFDH2Avklg9j3fEVqkOZp
/WRrtTO6oO8PNI/Xe6prh4o3C6nd/Q89aHqTrx0VMVKahUkFqjhryfPjGGhRDkyc
CpVR+b3u+i5kPvB3aPYk81e7YR+tzHfNzhWW/YgrWaJ8FJiuwJgQqF93FSj3IECY
ReBJ7j/xXgW6w7mod+rsYGV8LPE2AIAAdVOnvEwbF0qdBOg8wAXSlVXwQEXLADWQ
CrlhpFK3gWU2wuuN0XmUG/gcc0MgKlddTQEX9mN02BeLa5w/5uORPmlyA4TBGZ62
i1gzd1mlHRjEZJpHpmkPEwTSlHUWH9YoSPxNvPvJrvfFedfCLc3HCp6XHK++av8Q
Il/7aXBcS9JRtZ/dKyMgH35yf0fAIwYo5cC471oktvZY/1uRtXVjBq5BOpuiaICm
uNzk0w4RPn7iTekrfxlsI39YjRhVH+KSHL718mFXg5jvaWHU5d9t0B370ZPmcwqv
SZ6/qMwjbVSwqdLOYFHI4ZyCc6XW1joCQKep34Mugbpoy09LHNavKzRWi/jWJ5g4
HNk22ILLSrBGaHkRkctNkDBk9En90a/8d+qY6ecyZ/uUmelzuii6EVqkk2CTzqjE
c0GREm/UK6TUpS53KPlQNJK6bDPUtrbXloCNHMJJ0WjHVUVmKqwqJuBGzNA4nXUt
0MsuajiGIrN+aiIWl7p2QxMJgu9olVE+/2v0FpaVaaYQfiGkEI3Z17CkRdJRBRxd
m0KmcxfT9TodRjDa2Z5wN6I2kzdsZbS7USLuy0+2gmbT/2ElVUQndjrv/zJltqs3
C90CL//m73uzxMQhAY3A/+U0X9iw3Hktushv7vV7X5liw3uMm4XplqldMQpebz1Z
W85ptLT2/2GSChjPcob4XdBNy7fXeqBfw8xqX39hP6GPG3LgqopvorQZ0bhNpQE3
s7hHpUc/v5IfKLYZEvJuiKG4ToXZR5uYxQHBGOCILeWShN5NMR0H2cJwc4ywVAk6
fV64e1hhd0Q9gDH6udNl4Oe6Mb3bw8zNOV2H2oLJ8uXa+FKCy4Uk1yjYQ+xMWATG
gr57o7oXWtXAVFLqQlgSqdaH/gAgqrkP5QHHQDOoPRQjZqTKFI7C+R935YnarnId
idnFfK5KxEMnbM2omkl2MWdLwQtB0XLor4PEVUPclhvuHrLrCax9ZxOTIl7ovr9v
BUubY584upboZmqu78q5ov3tvsOewpaIN2tvZYl2sNPaHdiREJrRuLU7SdXR9fFE
kBiO7XoI8tojZGWjBY2MHIVKvqB7uDzOuZ4BVTl0v6DA3R927XqLcqMTbZ2T8rqk
9/3ONi2LFGZVsQZMNToxMIRt1aoxtJiFe/Ccx8lpT1g62Bbinp5oJaWMHVe+Q/lO
zddmzXv/MJ9PY1/ItalepAw2/Zi0ORku/SjN6Np/MHYGwdcP93P6HEIarbQhBeGh
MOe49gnzt+DwLb2nC9P10O/UjdkdFMRxZi8FHEAqzNZPy5dRrMIT7RnCM6CLt36N
sCDb49ZlUtyKm0wPGNMSr0yjconNrPekCKzqeOtExiojnpdb0nE1SWKs7LrJWSQa
ikEekXu1s518zYG1wXoSediCAeQ3zoGbHoZaPScJ8sGqZrxnQPN578sOCHOzgquD
HyWuaUKx6i2AAMuXX3m6PDDhTVummkQNePqD7/KxQ0KQbL7n2wJ2jf1wA6rSbHwr
DLLIH8ZG6xZixX569QKTCbUH56thRNSxyyY7zICc7ecPyihzDwwAd0RU1M5myw3X
cUwjVH0wdtJmZVzgIOKGHjuwcou3NMzD2EqTLFi7X7tGWU8UmF43NMHvVkBO7tL1
t/u/VTHuGpkdColTcLZvPWE24FgylbD/IsqkJOQYB0wtW+A2psAYjrulFC8CKOjR
6utegPXhdkpF1FecREj8F5tZ3UMQbcqqei+bJCrNTHC5aP18ziEdfKw4z0nFPogJ
NNVEmnsWYJwbjUKD4Fj4vB6+u5VYjD/Ld+530QOYDsGpL0K+rqFEferxW9okyACM
zuaTfR1UmwJcwQEAn/2AkRDrDTlK4+1I+EHYK5iw9Puc68DBNAzWJZUvUpvw+9Ph
9ftC4X9bNtqxbiZQRDaVBYWKHA2coxe8SHk81pW/nna+ZyIFGwfN88OSLR8neCIs
Fis8ExrS0e57RV/QObOsl9EVNBUW14kYpOIiC5O6GCWSKquPraDLMeUmeP5alyAy
THFIti8PeOSS9wKw0yvnP+PESxRlOv6vaBYTof+S9Mo5EWxo8KCrmc+Jyg+Nf0rb
VARnTknx+p0txwNNIDm1+uN4yGYNefGw8WVWUPRGDQWqHycKokhi4Ivjxe/b4Jk9
rCj05raCVp3y4bwE+OWhdAYuFe8nvKW3XmdqgiN25tOIj4mOgyjba6/qLhz91OAf
IMV6k5Ym/oiCmmIHybsAKv3ed21e+C7Y1pWaATWJM87kPCrns4oubgQUGgxO3Qeh
+2WvYIoT4RN0IlfTCMIE5CJuj/70AiblIzEa/gN9GXQG/lvpXqYKPyVeee0SbTgN
yGZ8C+hAIvI/EPhzmhoHKHKyHvWjcvEbNVR4NsiLcx3PejWgyoAz/n0NAMz8C3R0
3Mqvgyh9Wdwk+Uk9mpZQD7ilKiQODGW8xBvAmhURFYPLJ09jWuasa8uu8l55tQsT
dO/yqxZwHWbrqAywZ0qrz9liW1WlwuXFwSzcQt21r2UY8o25I89lN1l2umr6SPcn
YesUf/yga9ZAuUkKP3BGrks8HJ80QhbThLv9ZKUTQYdQ84x9gCYifkKxBYLckem1
BKz6KiT2Z6XDzQ7T8lxnXguC0WHTRRrgJmJPN1Y+I6ZWbn86xoYhp8KPT4Uq/VFY
aiKOROTlTK1igTIaz0jsK7zCOuaL1Efm7tPJUNnRFyPRNpehqWav8KW9oqSOhwEG
9HLIEGqZal1pFu7GONKQJeAdwmAL/kIRja74L5zTIv0IG7zTRTQmQZoU7Eeiiz7a
sStOBj2+bnsVWaZxi1kuizbqsPJ1hJ6rbYqXeCJB8xgJzwHIn8uMjc8pABcIAXSV
2o1Fn9n//vAPe8IeWYwdKhAOoEPuPRWZdaQJvfjvcAFM2E+uVdFv+TqxbNg8zKg8
pxAEi4ZvSc11f3gTDX/VkQ7tg+W6Wa/R1OBwtGpIdsbfwrF2CW69LFzK6DYnbQC2
HNd/03aKufx/LbhuKZSh/zrkcXW2HipcwNvPt0tDHPEnJIDLwh/Ewhtunk0/Oppd
h8pQjptuF/JnwaGNRo7krGrMgmPxyqjAUnhreIjMyUIY8JSDnqJAOZoJ5TWnFhDg
871cXAsIjNzcSbJ8S18INf5ktJYS8VGejTOa9dzp4zfEjseJM3AeDjbumIeHs5/c
YlGGOVajjtPBVrTrEs0okngl8mWraAwx3X3mthejsHNK2t274oLEoBqIFfc2WwAC
/rA9LQYkTJ1lP8UcZBIRZB7frKx8L2eml3O5Z0KtJCkfcLyc9OA3HJWS3jNwl0RP
VI+TZc7StE3MrQVtu4M3zvq4c96G+44byHTFZnVbOfBbRkPSrksDpj3/wFEpQJp1
kSjJFL6RtGRDM35/6enTDhoruH3LroVR3WPVzAV+QMHWZAn0sqj8Btu+SxU/4EOK
X5S2h8wikCrrFT4mmAvHQvlI9nHLiv5Y3XAULJdwYv+28SlkHQ4bMbpEa0DCHFeC
xUiVwNh3PJr7OXBh8SqS7CRKkPsNXmo5RolFZU6KDYMa6b4KD8i7vG2MNr9tH6BG
UX5y78UZih3MtviwWnGxb/mtGzatgDH82xpvzW9f4GtC++fPTbbY6arb7qKDeHS6
DDy45nt5R3kORkfDr+GDW+lBF4H62aDEKL7e78ZGVq+6JMhRe6u0wPrushbYS64L
CtIrrHAosnK+S0x2n0/Z3aCPIOhAHN668hJH646TW5Dtq20UK6QgPEnlnyj0V4Pg
CRtpsgWxACZg953HMhvwZuHhY7XtHjePJjv48r9syyM4/5s5n8EPe4StZGDucRjM
LgFqfanl40mO5saLwStfH6qlHJFDTsqGvSLj9L+jZeGxV6R4b4Ez7pxHWX6v4KgD
td9smQnP+Ea9Pt7oKIYLPkPthsCRIxF05TuQu+6b5ldz1JhZejxUrW0pXx2rzybn
3j0vbUQJNBMbQCy8uilzLoldTYgrWF9ZE/6kEtb3k6/UdBIuuBkCJ9BCg9OKsnYq
vEf117PYd8z6waGevQNnO0FtceYY1Oa6c+GDT5bppiP+Oe+FW199OfcrTsuV85KX
KBWI99Xur1sVWZXVGobTRg8HUO+7Mir9rbdrm/BxFa2DrqySUIMNy7ftuo5XAjxu
r0Ll9baz55dNFBkmc0UOv+iQuP6o1Y4sE262Y8oerGiZAWY+fyvu563P1AZ52e+U
G1V3wOzmYKXA3Y6HiutrHmQGI4bRgvWV0AHxZzIp68IxsVzn9LriOubQcdcqrgjQ
XutyvCIo9+9qLR1mkjXN8agPz3OKPDFMClSZPT82Q7FZLTkUf4Bk9OVBRfg9t51p
2nF4/Xyi3DbWZJBef/bv2KxyMtzml94gwvUVU4VdqTpoth4ymW5R8NfhH0DN3uD1
JNQQURV6Vr4SLB/pfnBz17/s1CEhS4bmnSYJXXpTxyac3ApPwsvv9K38qLkj8JSj
TaOBgRHYhc5AQbm6M7kLrzRlY9zg7FJ4DR1xXrjakHRsDJxS/A2gMX3LA1gFh3+H
Tew4NIRVlptLeL0LVv7HPcGMcgOtNzd7Q1fPgDNiWSOLiC4c+H+QAq40OAtX3Pnz
VEVMf/NzMq4CbNo3GcfAsb7aDrJd8hzKA5ws4/NDpaL9OhJDqfHbInX6t7ewr7SP
XiwP65hLb2MSuiTNhoFa6uc7eRZ2bTMcwbqB741Y3O+pO3ulvmSPVeoRAAaeN1Cn
QhW7Ats3S19vcXhd+MXN81mE+/Sz9vFhovQcbTTMyxk81B/8UN1ZACHV81bt0wqO
VZ+yGpx7te4talO4EPvyBWl+XMOSm5hvToKvM2mSGT1o35geoDloyjOVniMr3BEE
HWGOejJk0ZY7k1IPTflQUYphb1/m5BHdQ5ia03QeiOjbrNyMRMv8ap1KC4qkqmcA
e8BVLPcts61qFIfNtdwyTsJG9JCtipRPWpICO2PshlB9LqS11Q11gRMKpDy1CJEe
X5+mgRYndskJ7YEIw4s6kVYhUSquLx6Lfq9YHVb+r1Ox452RRt8VpXQoC9LRVZDR
u+YL1vH32+ER7naxCInirxCKF5JDkaQZ25xeP85VUfDTGQUi6dvtYnLYpT1XMdV9
upvQoppUx2JLSF72xuKUt3h/vi/V/422wMZX+4zOi1Ifpu/PBsl8K+8SirYj7zkp
jvkfq7iIHE5f7tE4wvVUIgsP6a8xKrizyIN7+lGnaNrREC82rVB9gFApKoykEnfD
VNt4MK24WRrKVXde7EEgvfRAsN7tOldoyAkzKXPSlVTAQrj23i0SuQGNPT9TGTOh
0Fqcjy5Qu789zeAgLJGGViE3vgzdcB/LE8bZGghEUc03uykZfFFemnkz1HlvpUmh
1jOyKdwakht1xff84jKjoymYL5HXdHngQ3fxVShVpTUqh+pJwySDAPUjpy8xkZCv
n7SOgBr2W7l5C80jK5IklHoRk4NuzsrXylkzu6kpmBAmicKD/WHJqKUQYLQNOhlL
RJautPjBgNnbVuUFsixM7Oa1jBLde8i5PkEkCgmsSOXitnNnJqt3U6N8daw2fHht
CQ4YMZT7k+Vekxjn2g8GQGvcIJYJ6MxzKF+3w4Z8v4DvvsY8aK6ji3v9RziS8uFz
Ot+XYVm668mOXX1mw3B131mBDKqo0cytmyjR7ACVzEfjMXVNMJ1BC0hYscn7jC/m
HTVo6m7mr3Nc786s3nO8fKnod+8FTZOcEeWvSJrbXLQURxGGVyKAAdoltBcQJh/U
xRegZr1I3803eM0I5PYj019TjD6tXx12ehoyKG1+uB3RK8VgaTMH+dn2sMt3/5hX
UGKbAG/SPfSSfY+3FvBs9ZzH0J8+ISPB8cGHd0B1A/9T379vWrg0bgHmr0ipFiFQ
xpnmy4bsEJIV0ALOflB5Os9AkMM7RD6WEJaNTkXLnlPunWm5jtR/vqWiATxMt0f0
AUSOPvECTTyCWQgDDIjCWZ8sPQom0K60PyRKD9Ur5v3YKME03uoImqkFsAAITOPB
JrdzJmUsa86zfE2C45HUIkBCnB9WRFA6Bc2/TGYmS3MPkcl3Y+cvh346u6oz328m
dwSNtcjsmKo6rIkSzP+U3gxOQU8BTMJl4cy1d6AUj9RTAin57Ya5TCc+kX80uttF
qb6uD4YGqV/MZcsqvUEIK2EgNsmTOMj0SpKMshP6210dc72qCD3AuBh2yf5fCcRv
m4jbQQuluVPXKVoFUDulOaCvzRsf56cwYOZtKC540L3flwSyxv/zLaGmada8Z4yU
Vod3MeKg+/IFvatpS3h9icjmQbd3UIazVEsrRLx5L5ucEA+juMtXyR193bUGR7zP
hqadY4+vIR8uFJmzfMoqevedKLzHIvro4Mm2yPqVESpF0SHIkfD88aPtMOl7j3CO
ihDrOdzwd0NGTjyca1Ud1E04Xq+EAHCPYylhDddlHp4LnUGPb+4jZ+9+TP/LNvcj
XMXHZBJhvaYQvPOiupG2c+sVyaVzZewwe1jRdU784uuC2WVzDvYo9r/YaC0omyr7
1k+6DRD4UBuVi+ybSD9pKLWprQCacanQKzgPIxh9+XfxiVnjUrlURV5mQTaHowfl
iee6g3rBDTU8L+kxw5RUYZTFuQUbeTXFmvurIX1IWsAZ4stBIx2bDdIXMC+55opP
RGFsiNoDCzMNDENB4OjDgxMtjpuEY4cajGi4FNB5qpLnPTatXYpHXPcN2Xv1pwbQ
PF5/z1gB/Kjvr7zT+fBTwJ9CHjPLzv4UUspRivcQwgXLS2o4jCM/Opi+T300Qws5
m4Nincep5wRezrQm5vUGyFAWc6u5G/GWtdahzxv+WlK2mlx77VZhr6XajWWVYjbj
w8eO3l0tUxYB1fQD7HaMh/Q4ZjqUMipG0sersZj/A62qweIXKQ6I5VF1BEq1WvQb
tR01rRmdQdjvv3nGiJrMwU2bDlMdENpZ09RSSO9RabLQhrbiOBqjAgYfhZreKe7s
wy8AF9kB52kpoGemG9UUlZnUK9rJA4aWV5wegyfzGq/yfC2+shkJ9xLDd9V7XZFG
zeZhQekbJr7pgEkmnA0EOYR1TMfy9ejiqyJCyaS9nc5WX4gjXdvs4CJlxWBoJUX+
vTnszZejgUXr7dEnxatkL4JgGC2L1DY5P1msTLRKGthyeSa3SgJ2920a3GMBSehC
Ssr484wCWH9TL1FPjT2RJ4ChxbTWqGjWAOE1HBdrFeNIBlCPqUFpB6G70EnOTbDV
Ber0qZfMGqwNnszvlNOdkkufxmIs/718IRLPoLgdAcLtSmyHPqVfJ6fD4J2fmmts
xYz6xs5+kWSpn5JrqBLeNLd0kRV7LTyDurp2U4kupy4/W3SheMM6RXRhc8So9F7z
a1LS6OXctAOvz5qn4LWaZqBqIak+9Dkp8QfO0vhp99Ckh53uV6MtM4tyKhHLSq1W
2A+gTc/V8LczSeRLpgJoYbXIp+RNO/RGzsk95Z9Ley2lOnsIGTcMSlz1aCYcEqIS
FoJcA1XdWT3He9gTzkotwzqfMP7LeZT1ygulmHutcqrecCVAKhPVAhbwwxjkX+jL
V+S2+/6y78lhuvKdnRvSvl2FwCdHblDzQqPSKoh9pLETrtJzi6chveXM3lIcM6IA
TKjWMV1rbf+A5Oc/0yjyAMzh1S33vBaR5Ii76+Pfk6p4rNpK4xEcHzMzVmpKY0Pf
PKz0KC/qMcoshN29R0eFjnhIl2lHTk33WPYCxo6JxN3XdoWu7x6jfYsc5Cho4ie1
lCAwgPlhGQFge2Um4YnVseHZqZRm2wTU/Jm0fhwfUWlEEVavUnfB6EaUTg+11bae
yiIsfrP6i2fsDyUIILPXBnLpNNy36M5Zu/mEWmazBRsAwoeT7fbMAhLvbd0qI3Im
AASPMA+2CI7tsNDqIJhmA0Tv+H2ldwT/+o4ta0f7WiJxgbiWrWXO1bVZXZ0thz6E
2iQ9T/K9Znq9OGhPS9ylssW+dnZyH+93mCWSJCGWk7bxQwcxNh+AQfJNYhexrqwF
DYjRwegSeUwW+ERGyGM4pPFHH2EqzYmr8LUMWvXDwOiAJFXuyDdrxsI0wwOUOJZb
Idq+xAyjQkp0hsKqHhoc8NFGQFw5WRPGrswv7pimT9asbzdO33wsDy3as+KDeokr
MhIyFT4gn/Betf7JCjmsZ/La6lH50KcoGyYAFzfC0bQ3Qy6/DzPPiTj73qn5bYe5
9UqceixTZVc6rKGb1qWUL3SOr7R+qma3gLTVjcsh6kxN0u4rwrdb2I2tZt7YCRI4
7YayfEviXmMmZR0EQm8pMiqksmqPt0r186nVX+ws34ACBsq6mOAtJprsYdmpOrIT
eYuZ+hyqKKW8DdPqgaAXTBm2tLxkY7NLG9xKZHhanzLbrsjV+tHRTxGfNwMjbBXO
/f33TEXLsA8cKb/rw9cdnTmLKxJKsjFXxy6KkTPrZIsZQ4tAEv2jaTZg1qyw1IQ3
gVT0k2G5xLtB8DnRRCLL9r6GnSzXXMxe0ts3nZO9y7LOviRcCc23BESgcR1rX1SB
QM9FaGt2AqddXrMBJgWmTqVCKscYElMta+gVm3TkMyyVejkxqoMfmrYMigPbbahA
FELgmfGzfKFgXOMRufXYB0gU+izL2zpIBLK21PneIyt39WlywdvMtd8Oe52eNvU2
roRavXu7lwwCMYU8zQsyJlnJUCc2IFwkaepTIFOgKIyLy9Tv878tzpZifoM6/4gJ
dhcCYWJnsZmFCLveywtbTRfM14cBiv9KZpaQ9FKetSaji8x0SbibvtzzuVK92GPl
/HY8/wNTtW6nPgLExzMr7WhPdZQogLtq1pKuf8sw6KUeHTKfSqzIy/KgpIhv6Zf4
9+5dpMt+1xbLmBaspUrdnf72i9AAiLjYKy4xZ0iwMEgznwEqouxJeXA2Si8Y0n8k
82dDr5UZkcF6IbzdqCOWxVyj1IlnudszUGE/ySFNWVyPWRNAYIcT97exF3miY2cn
26IfjOvuigRE0oc+bSV9DAd2l1wbPsjkpEwuotmxDbKBbJKnu0WoGAjciNTgymb9
SMyfKeTwEZ9oplf3ctaFr4MPWxkPhRIIM/nDUb/KgYT2k/OKg3A3EHZUdkbwrW3B
XZP4UfUxshnfmT/2Civ8FmA+uXRZ3+yNVbdQ5TY4cp3p0Xgc7PMd6bIJlB4Mrepm
/ZqAKXBhBQ28ebmx5IbOV6d1CC61MwEQHzrkSGRT+KoCoPk6/0bn6l60eJGk17cf
qwAmcawciyfpERobpEuLewAx2cnKtmlxVZU+so5wa10ipwS4hoML5N32oi6FFMgi
rg6GN1PhagJcFjjP4lGzkQMC0X1hDPXx1R5BnNfVAgOhdmFLbTAAm95k+c5WU1ev
o++1BW/4ROU/jU3jH1cAApSIlIlPnaKx4npm2i3wo9PbJ9DP9dTw5uzbGgxQeeAI
AP4xZqwjCMoLCqiJJhGpCfpil3IgTx4UlXotfkrTSPgGbvOknvu7JxUoskF0SpwF
9BcGnILsq+E2CJTJzuzO7KS5sD/96nNJYQTCSJth7wSJELM7x9FqDiA9e6FCNQ1l
zs6LGWcI3WbmFXFGQ/WqYLlv7J74RHxjQWbDGMaAtH3bXHtPRE6+glKgMV9HsDv4
hPJu17nMqoGlJnuGgbh6XkMgmpEWk6vdoNPw8hWvxBNde1NmxxALd6JGr/NGkHRW
WS06s1UbqLkTSGJ0j5uU3CwfOAcNS9S/ontHzXHNhl+I2y1BdUH16wKxkbBSd7lk
mRzWqDEp24FnEdnJWfgvl8TkKCryY2XRtmwbI2s3SNs5sF3OH8Wuklb6PcOK+lry
UuWY49QR0SXrkpalDGK06+xiIl3m/J9cUOL32172//ggYUo38E9A0u9TPpdOw55+
/oxvEc87MmYgeVirKSDDRZQxKOHS/MOm4mn4WgV96YgsbOcHzuU/OeavfeNsjzOr
9+lFAFr0NEteLzcPJvH5nho3PHL46XE3/O/4ndJ4q3FdktjBoQxRIeGAx6X/i/SN
xDinMzYp5opifQxA0fIx1YFUV3HD3TtWDcfdyEUlI19UGUi/8frVJOAe9XfCQ06g
BbxjsF/IrcGoOsXpSBSQoLW1RFjzYmaOn4dMjvUI5FbHkj+WVT58wQbjcJmwH1w2
aHW3nvzqgWkLiRnswob9p1NpU1eVNlvWJnmGeF7TqVz8g/7JL1Xuho8M8SkQfFdD
bA2dbMScq5ds4ASqDmpknVXJeRsksZ0Ti31Xd1Q3VRn4ye44oCkpbB+5dR2Hr6Lg
yB5WZ4APm9bkIMZR70LVeytqQNASb6lAB896EI/3TVHpH75yHlQe9cRzNne9qC0n
zVi/m5GsL+DxAXgLF4o/B8RnWMvuEpQRHB7/ArVKJ4ds1B4oichON4BrMdGknApE
oE/kN2aHpRAJKU16aOpI8twdMU5PylKSurKU4DcWZ0eAS7qoMvPRgbElrHdffU/1
3rYc0JxVKB+REdnm1ajIuitZv2MsOJLrP1GlEiKnphaOUuh4AiuVXF42eudJFvP+
si3TfhxNu+k6K9g87hDJnwd4COJdtCnKM6wlgpwaKF/E815F+JQUbZ3p4ADBzNr9
cNuPYxbbMxJ/AorlPKMuOHI+K6KexBELsf6bc7UVbO1g4V7muDkF7bpRsXoc6Ze4
ygjd5mNSSYabLa6JiJuu5MBB48nC7C/ttzjhMENQHyb8Oq1zPeryEaPoFjBKqjkQ
jG+zTM2I2N21Go/OoamBbehnG77GQ5XH+mcPgcPxWFmVKki0wffR+hOAfUjULbK0
eO11r5ZC3J4pLNZt5W3FnyQ2jWqz6aOM1B8cpjun7BLMzmLHkVzHkkJ4SeyodvYA
z9lLKcoFFFrkh/21yRQB3MqSUXKj6aixUDAh2DriCIXrQi3AT/TBDoul0zoXTwAF
8MB4Wg7Uo2axhz+GZlmql7ysQ1ohgAUkzNq/dilJoDi23ERRr7cUsI5U55l1nOy1
cFv3fqdOAzOZUSop/D4VkkBZ62yw49lV2c4TaljlVzBcIDYgLfmiekmu4CWpeDTl
QTpwbyxw48oQ0tln2fOav1BJ79AN0D/iNuhAR3p5yzrH7tflMe46gen/FTC4mxIW
+pyvi1Nhkp9k53sLakgHrup0Y6c9zzQqjwgT2EvAQLpjN2A0oQ1TJYu/HnthwIlE
/z8T69PV+VprxTD6ZGmgC/HLCgUweG/+YGiSYP9C8ROlnvlcpfPz4+AJBDKKXWgt
Ye01NVpeRXOFk5BV42WMkIt43TbTzmm1I/M3RhJa4bohfsMFm8/wTnnUuuYMVcYT
EokLHgtA9dZTyQO5ZJD5EB9YtG8PwXkSc08pVRDVtmDg4bvXsKjAE47vl8k0e296
QpdB/yOVTQ7L7C7eYPabyTTJj1b1aV6ggOW/vd4SwlO9pD5pgM6NjIktR4GcKRpm
tZ1IFXACQL5f7D1Z4SczHdDg8/rx7CwcTvnMCdT/Rp63hhH1+JxjRxVrus1KuaOk
OqOUjHTRk4kMjZ2E0xJKMJgONUjUGHTYF43xT+ijsL4NkuKKXlNy7Odzt8XiCKUQ
VZMGDNu6dEv/A5NyEkwAdHl3tK8son6XDu3MG+qWtKiF4ki/Np/pkKWzBb2TjUQS
1pLHymBhAQGJqfEREpvwGOtfUbTmWbaMz5paArD3+EP0UJtYDDpChMWFIPzftQ2J
uixANSA+hSjIUnLYPs+iVJOsI+pkmheFw/2uNoGDwXdwYfF2NlGIRSh/UVzFcuf2
93fsq9EaQR9dNfql2t9ps8BzyfevwShiuuZdUioKTxM/z6labU85QtM01nELk5YT
dia/xTEyNVQZATgRObtWUG8SUjYXolj/S5eGuWuzvJT1dmbdyTKmn8t3vyum9jaZ
BWHYJcm4Tf3IMkRs6cUFvhFAvwoVVnRHMm8PJezoeeNozo6bYkKefnWcizJiOHTt
flq8aT/8GS+E2kIAIAzyGeNyJeNOrLi894oHbIEPvksA+spX5Y6EZ6AWQVRGUrrr
nnLuEKMv/VRdmPUgWZHLdC5pQfqjsTQFFD7qbfRJy0eyRhiBLedMWH3oZpwAND3z
HWPLeqDq4lc6/F0R1RxajLlef9cAdKXYu+Lyqiaiqn5UEs8nEe/x7tKkZnn+NuQ2
rlcCoFml6EvTHhrL7C/tPqHvYHADloTSzsAZj27EnHHc+OEeFR6PFQe6/j/cPEei
QUIeDDQ+ENaJJdIhvGRsdfG3WsB6ZXTyyfKOo3t/SNfYqb8Ab0eupe9KugzxHItZ
2WnMfRa30Am0T4M//9ywQ7/DTq9AvnAKX2rcSfamRh5KKwLMifqxjCXk1sy3ORiE
DV7w4Gik60+1H9e7sYyW4QJ3yP/ZqLdlmTdL48vxmNCS1wSst71sUtGwF5t7nzpv
wlIuSQtHbvRpRnsetbcq30udHtPa4ewjUTkgPhZROP+d6uEW7osrsyyj8VM7axNW
kWOYJ5pr9KJ+KSF6dyDiyTZ8R31oZ5g46sgv+FkEwqOWVSaPT1gdpahwspTxIqlZ
8IJxtjIIXNpw+ZQ+c96tq523RZFmsW9XKeLUTQnsuY1hTEYyvuUEF/th2EtAaZlZ
PNdyypkHvVdzlpuocUgZ8lauKedewdBJaHupRa+o8BnslCqwy1Hau+yl1jTK/0Gz
UQBTewC+NyPOLsxfmtCog6ipSr0dyRnIMESm+LrapXfii6kbuuXEm2kAJRraciBd
Nk+D2AkxjZ/RePyRBb83f6oqFgWvOrLgnzYnZOVY7zEQ/eAJ9RXnkYSHWW2DgunT
Ct4GxtqzVKdbnQlGP1ACg2LwHF2H9q6Uo3KKdhpTp9FwtMnNQvhJeZnPJqlrjrcz
xRfm1K118aRo1QfmGe6pXULaYSs/739H9DtLiRpuhrCERoyNgeebeb0dvYGTuame
xGhJE8JnxBPeXO9llCzcJaj92nRaC14s0fZOOzUYivqDEkMugSoqJP7VSuQyLXmk
xpMr2BRGfCvPfXFU+8evm1yLYnFytQJPRXcmdj+jS+IqdsYD9quhLaPAViszC/Ax
Tkr8N/ysCaMNtZuHtNWwlqirpmax6lOcRw/3AUOcw0P5YGyEfTbwtGOpU4swJGZx
mnPiEsa+2+XlVAeAISjLq1ePAaPm7wdCcZd9py1NZmUbQGy4nB/cQKHyYClzsse4
PwPNjM54rf297sv0A+aaYpASUWvA/+RomEZtASpibpCvUQjLGhuS/TX1sQvTICwz
oqA2+5+qDqU92hCv7F6cqsRHdRVQVp4biRwTLczW8IQQUrw0d7y12EMeyyb/65sN
XYBKInuga7Tq2SOz+Z/Kpajyvg/BAqVJjP22m0357zTd4hLfG1hntJblVGy8KiJC
i9mgweMKteQpR0HQ3pxkxsBeGL2tx8ueq4BGoZKZoQQjiH5KyBVx56sjjpkUwTye
s31qvGRBY8/NPCUoSwI0eGYkPMcXhLjyygq5es1t4cs/EOQYy6PDp+Wc6RdJsgv1
vRCc1LpxqsssMAwlX/kkP8Wvy/DQpYkk839nSsE9kOT9kDDSpWHMThd+I130PcU1
KzmuSr/8WDcqTs1p3eRzH8Yhibkk+JJwvVTK+vUhJKEwM6dsc1SXfD5YVPcd1Mpr
VOTZQo9auNh6y0GIIUPvMM1UCCFMhi3j/wtz+C4KM4X9d3/Dm1Tg+XofvfcbWdUd
Xk3OkvKFNcPeaFP1xEgnyY26xISuuyEMfwk5aUKgdPrfEqV1wx6S0X5KZ/Hpi3aI
8uv4NVQrzUzljMePjVmIusWjadj68cR7PMn087yYutdr7jF/g/inEekGkdmNfgoz
m8LinN85fF2jp8yg+wNDJX6BkCoH+UKukSwWdrriOuwq48G0gO2P2O79S6B8ib9r
Lb8UWeb0WhZq13RQNP1NYy3feaDTkJ63WxDlHr3dGZJfVVYWVN8HItDyZq+14qtj
HXB5qsDo5MlL/Rtt/yo7GayXY1i2VX6iXH0AHQaS50cNM14OALWnj/RB1iK76ABm
YINz1Lzzz0dkl8+M3rCJ9yFEErFe4Nv2EsOILEM8nlizV6G1zIF8FjlXImFzjlZF
PZYlBCKXrccBZKaUGPK7FuMBSH8mF04aTTtfeiG/D1Q6dG5QvOcT4pWLUgd1Jfga
SlA4/DpwCTb5DOm5mp+9GX+bbX4OmPHCpCOMAGp0UcVAWAyOimiumcFfG4xiw4m2
D+b/kXLJX2swrFFIbOBGCPV+RCfot+1roe77mzCN0OU9kBNVYmGdo1ZnlZ4Tm/b/
+XTzy347kebGdhd46anfXcDWAw7cZwNtdvRzppM+sTUaPDlbSVTEo4RC8cy2XmWj
C+i9LxWj7psOVDBk3y36PRAySmKfOvOz8nJs1iqmEuX1FyxYRlE40TAxoIlLEABQ
T+KIauRbPCoOli2/mSJ6dg4ENhuJRKN3pyxu7gk1Ft5GyMYKBIKct2NCULcuzUSq
5Gnc2lfo4t/+SScg1bF7TOk6cmRUBYAjDy9SGFF1NxdxQOZejUGeZiKYR9G7+Mrt
xN2f8OElsPT8IvRpsZRXJpskDQFdUwiTB3I8HmsJpVuIhmydXRruedMNKrYTkB46
hDhZjuOuG7v8lkJ48KuMKpM97/SDqZvFAPcCSn2AgWET17wv0hzny1ATJyjIymn+
M1nzMQraT+KTiaQF7EHvubARmDGpoyyyp6FsUMgYxnJK6zsk4aY1cv7/vjxBi8X5
Wv4BNIT7pGqHhh8zHzUZqgI/CLfCJIeuujaWk0z59oDOXuAVkEK3Mc2vgBD/kRA0
bMyu+uqzVaRqJ5weZHSCMMEqa0EkUFZ+6JshbJp85Jp3n3Vo7OGRFr/sLZpDiizN
OoTTErJZrZKrKdH7uz3ItTJZXGWEWYqXrVuY0P2iYfS8sAY90ImhE9iCSchqNpxL
3mHn7//reUkYP+T/VQSkyUTwU1Vc+kHtpm+qE3ATpVE0ccWiEEdRmitvJZwvQn60
98YhOuD09eRGjZMQXbDUupryFEIZoLJaeelnYookk+gfxZ/nmFSDIIwd2ROzXNgq
4ONJJ5jB1yBPDz9fPDs1qkaLsfEfQNpsjjVxx5cBHJjKtL7uLQZ+/a7qnywuIy6W
H7zvB1aETngrlCnUxWk5o5KKs73GB6IAN8iP++le/5TxsHGJymBl76qhohheRmP+
kD+Dr6UwDO4K++I2RA/ujkWykhGqyN3Jdlx0ADet+PkmD8Ol3yB/sdF7QOgZdINm
mlFptlaEbf1p963jtKcVTyIQjyXkLf38UocRjiyzc08G/BtlOl14l8XgTVd20UDg
GOIcbcG5rjenWRA2TmiuyObmCc4X4KH0tyQJeYvI7HEDZUUmdaHfN3eEBfDe2APL
jcecdb6T6Xozj4SFGivFyUH6qwzZJ5c7NQsTmxAi+BXj2fy5mq2xl3S1TX481iLI
qwmF19WNwy3D57eLbBRgVDtRuXlp/SThGPOtSFbe4hQbgBAA42WBIegNV2hoXrYQ
XAaaF47qqDn0+YXl/2kEYm0J6k5nMGc9UL/y145Wr8vo++4eJqysJJhAaki8QmQU
AeZ6xmfsWjb0nXAhAIu8iI3GmeUQijkLuOMOEHJVNDZZpnkrmi8ZSbPWH47nwlao
VO/3Y3OM+7oYFH0KTYGHAvfZZ9J1ecPgD478x2RDBrjhwhz+kbeDWpmem8JiKVMK
wgCBNV1gQMDr2n577KS2SPDKFHaN9nLuBqI23lQHXSw2RAOsiPpuFUT9ykHABraS
x4moQlollb1LYxRBaX3IW6fqsAQcpvnOaO22jhl0WP2qAFdWY9Y+uuy9u+3X7cJS
0iZo9jxrBHu1q5Sdf0Q9x64ZKL1/cbcDiHzsAxJ/2nYwsvUbEGhzpu+tNTwV/ySa
dHE58dRV/at/qMgzZPXk08gBP0DRA5ZDdXIg4wRZwM03OtSYO+nwFBS8EF21h0BL
djWsjHgBrhinwLCXI8uAyUtvR51VigtEdHLEvRHK+Zp7X5fhQO2mwUNtMHqeMQtK
WZ5tPRKdAG8ndr1Ti45ZfsWyBAtOjLhJV1g6ud8FdE3G4qY9C7ADH4G5zEW8iwca
da+2//jnx9lXYIbUHH56Zz/CGN8SAocmVPhvJNv0pLuVsJJhqc+JM0cYwPjol/jC
mUsdvxnMHvfbWnKJCTZ9LI8hbF8qsvdIEmpieT97wk6zJ+Dj8eSbXR4jV/C6wVFM
miqrR8Mnpj+FiA/P0UNnZYAidpddbjo40DulRQ35OczCvyeM7k/28xzTNLG+RcbV
prj/INV/91UAg1HPGgvZcyFxmTrGtTDBptKpjodoraR79Dt8OemiPwMfTtjcxgJZ
pPaUXixG4gasvaPefbb8qa79MjgXxzPQ0GKsQO22GQl9lwkHDlnyf4iauI9Qendg
9IVV0QPhpyYk61Kf3KrSRdfKjAl0/TkEsEFpsoqhVd8GFYPcJBrEDyDNFtmhGRqW
LyQYMZcSyqlOERhYIy5Uo/nz9XNeO3OpT9Twi/HDXkuIrHitLPrAqPGw+XRDnBM6
jVelcVecdS/OXD2S+edq71oWUfkIzLrYTaP91cMkUYl8cul5EAWH4zsIm4h3yW9H
WBwntw2YBnkMbNfa6zqyPDP1rDFDJggFm/HFhGd9az7Gb6u+7rJGtKjocRW7i9IO
ptXNu/pvznGm9bmmVuxjBcNILXGDbNd2l9XfhJUx9ZqycqXul+dHTeThy40od20A
boz8509xiFrDACw7+LDP+iUluqmkmzPKcNu3iNz+fkNHOB6FtOFzyY69SD868fzD
fcYs41zU9e1bbMNL81n8jnqhIwLWMecKpEH01U/cQIfZKrSgwgWcAEQlBa4Sm4OU
DJBlpgxw8xTofl593fRLIdjnL46Gp+expScfwFHs6LOm+GKyhWB4sOzamufpxtR2
z8cYls5m+v2jkSkqzhzFG69QBAkfLQWbox3kmm4bLcz1SdR9MevHYAucf7eZk8GE
15bBxtU1XMP56Fc1unspWYzIp8lFSxSsdoGdaGgci26BKGr7jq/OTXwO7nAx6Dl7
CF0eVBO6fxLZJPXQFAM4kIeVDUqZDEDrAvsBrVL4c9QwirXceG9px1cwQeAXCGG8
DmcadOOVSzpyJntzXugjtI49Qn64fCYB3nBZLwViYBplA7fuzwBc/ZEKI7pNKdMQ
4nT7d/+88t37Y5VLE1hQbH0ejDMh0+Xn62EzhiNbMVcIu3e2l7ShrnW6Jls13FdH
YYSPKiwfWsDOJgchSEelXdyDbP9sO8ROYVs12QsS1gWZRUXPjSxF7UAwhc6rPtwI
lhneCRDRLgdBsRezJamvrhVNSzDFrjvdv5Y40TQck/a94yKbDmtpGCjBNqrAGjF0
RIiLs8XCalncWM7V3gCwxzmsSJAEcbo3q+cxddcRW/zc/6tBwWbAePOADgZZTYTK
L9PSchZVTFoxshh/cD/txLJXuhXqQSFqh+IDrNWHHkD3U40YVBwi+gAuZoeGgbas
uw3lDwruYIPZvWIruLA/Rk5ckPidAaEv5vTSycH2auYLBpIen6eiH7fx9Q4I2PV2
o38muNO06lxNkia8ZMHAdi9CqxH/PD91Nie8vE89eucWY0/ISWAN3pEBcm/kgxAP
ZjGADCbPld5BHFRR5tdYqhPrFf2WTZCD1N+k1s8y3w9VN6+aHEDnbT+6EJdBdTCv
Jb1EfA0HQM5q2/VAxGDE/HIzFJfemVm0XlcSJvfZdGpuMWy7ExNdA0vbsy5U4vLC
YMtzZC+Og6Ed0PnxY9iWK/l4VJuXvKlo84UOf3DmHcHY+IUlo0g+LDgYfnQ8zmmb
oo+UK0Qi14g4jiBdREnRJ4wM0WQczen2hgCb9nmqAwhKfH0tnarBHegzvAuh7e4S
cVJM6eZpUdGAXGiT8vv1sW5rZTf7DPQLsiZuCfVek9tqDHjmkiYSm9ezZon1ELL9
vEP7bSv5L4KOtQZ7lyh27+yhKlVxMlg570OIngWVifjurWhpzjgFwk2Dg3hhOrio
D8iy783DRVD90QaihJJwRwiGRZxt9tEfwWJtG9RhI4uchtCDuL4sECDLvXoWITbl
Ri6jZ9YMw+/SJZlTH/L1p9JFSHrVg5AiExcFD8TOBKUnykqSjv5RB2+xw9x5QN/e
T8XHf/LAgMh0Xj9weTokIUYtateIuiCvx9aZLqQGXRVwfZ5iLL3myXf8oMFZWnuz
lB7lHoOsxpf6cuYKlmsfdteA3eb0VqEhliZJCnysiRmnePY+qa4UDRwmamMDozBZ
TXqIMd3BU5eSt5XapCBf818is6FGrgaf5r2eU/+KWXvwNEhfTiH5NZd4i4KJZmBk
BGrXYvYJu2js8TWexuB7a0qUVI0vC8/g3ZaO9EZzAl3yc9O3NX/yr7Q0DKtB2hKi
H3qmMQ+9++mAnEVahcIAqSUxmoEFVUCTS/rg+5/PIM3rP9hJ4JGJ3M5hwtk1X/br
IXG4EaFtPTcp+iJ/iW0V3b5uDmDjrzbqQs5f7URlif0ezuBHvZ2QNWRwXvfwXj95
me0BBLHpymQsh22dcpU1q4nEMgFtXfQrAyXL3JVxpam2Y1PxBuXEr38tgMLVV+jN
pLVCKOyqsdNgLfu43GHGppMtl4zIssdeIHMf9daA9TDnOl0TKFEOEiAutFZbzOiO
kHJIbkKNNkHtyJzO+PNnUkWa4Ks/TYqFvueN07Qz8GUS4t4g7BDy3kkuat8+2cqp
6YExTs6u8XkplMiq7EOcSF3p6tMPC4Kwaio2SMHssccFbZIPpiCqE0INrkkwWvJU
M72wa4e9H0Rv0oq3CT4mm+aqhkivfVHJx2AYHDQFplqODwjRabAPdmCwMCv7hOHQ
U/lJYKMcGZNfMZsVXgTQJW3pM/rVK5HpPg7Z8+w0DPGvu+m9w3ae78pDpce3BQif
AWRkfhXRp9WWxEVfaIe4/uv5zpLTNAZoGXE4F/7EPtdYvj8e7GOD03QiH7IAXmJ8
v5sUtdpSs/3u+LvfcsBnJOq99eqcbaWR0uQpiWbWgpKk2ISHtFxziApU0msd8J74
J6nZIJRn/GZm60y7VAkXLzIJgjnH9qMwuJvuPWJ1cM0Mu/PW/j/ozeJ7U9rdK5Z1
maFBaqwkHmZaJNBUXjTqAivGk1dbbKAqJQOVAZ227acbWmSNV0faIf3BxcAht2nh
fxUwhHzb4lO0GnF6s4hjbCIsySyxgarHVqWvQIBcs7dM3Sfw9g44EdMCVIwgAjlY
QjDxiRZ+GbNWYRV+u9WPr+r6UxzIgdKALphF3HxYIWSAXZaHW6EAm/XLGsKJhkfj
3a8i565OpR6ornKTFTICTIdf2JLD8+kiTadUZSpyqF5yvu3KMZb6YpPVju53eRQV
KfUz66GpcZlQHBEoP/bkNzx9b28V81Eny1yzVhI0pN/XNfzIqFiLf5WV9e/MpVxJ
WIW8r5EQVZ87J5m2HCrXuY02jtdHPX+ROzwD6mYVqTGInu0vGg/h9IKQjZsCy1go
NWxRQUyugeWGPaGb32KbwMFPtWuC4r+ElTMFZj64rfsTta3jLqI+cqnsNI9uQ6ek
eoHSMcfMODZFgfdv1NQailFCShxyNOBPS7N9apIIY0Zlime37oTBVunwrwZdRTus
NUC3V1buO4GfQ5euejKDFQGAHJ1jbUygo5g/Zh26hBgr8bturMk/VmpfNErTeQ3S
lKz02029hbW4o9jcCaILUdAqCJjAjEiyx8xRoiKfdmpfC4+enSwAiVORCXdD1kh6
OXTZCpjLQ7zLJOOaJ/DoybebN3L8Jx/GroeETNP2iTfRibc7xvSimO5quz2r+ZgQ
SXjxZD7okAvyTmPqe2wg/nkXo24AJJT6+NYlT2iJ8sUVgkj66nj7sxklCr8JtlKy
RbRieZNKZCoDom6yAaCBXd5m+oCfzfZ6sjsQuvYa9Oe/wW6JrWccENqy+OguPWug
+mKm2nzj8iu/ZJ2dnK0AHTXcq2BICUO/z945m39lSqYNNEQ3lVC7NQgr0VktJ4Nz
6AYY7erUzKUucXWJCGquqr6QKg3DANJhv3I0OBzuJZ10fBcVKYVhtivIPAfrNTpa
EIgYomPjPiAVPsNaltvnG8VeDgDGznhQtffdxG89hr6bwuct4otdBRC1Yu00tyHf
+I8ox2L0oOF4byYf7k9pJyMZrr9VaBxTX9mao1bHntG6DV3R8FxFNzSgDTREYVwp
7H2RGCUg+FNRBAT6Cjp1NPzvYQiJyjxFpLjbTDmxCiBxessmHw2EDNzwBUBKtuZS
Ih1S4nOzNVfdAMZsuTt3rQ/5iBj6nZsrYNZEg2d/xeKdlyFpyN8Z3f+Al0/VbAcm
MBj5Lt+uLX5u0wi07x5rkUW1H2JehE2ljcypIl89zFnTYkevoR0QY+v1aiKJ7620
vQuWKVSvsRnbcrM4jNZNLr2T0CbWFkmTk68trpJuckMosSBea3m+8TLpJbW+6DHk
RDT2QQau+fQdTyWNOQnrYX/4qCtK60pPKWhybRGumvj5S8Ud/xffD0OkQ//rt+KC
lta9cRBfkvue2oAKDeFcvNjU/bLfEDINDeOQ6WCoCHNMRADU0Rt8zOJnm9Lnd74N
EH3J9LlRcX+c73olnuxZLgABrPx7d9xsfJLzrZSzEPzUn+PkTHxhaf9iEuUr4J87
nF0Ht3OjR0jYwEtpx2+AGqxg4YeQTgpVzouVhoEBskhwFzS/JtTxbJXmURdvp/pN
rNW1DYlUaYZ0LS2wfJGIRxe+XxXnOhms8KkWnO4wXKfI5JzUH6rI8xqA9j1/oTk+
sPiIC+VfPptjulsXbeDNbebeWufAxaWTxBkscZao4qcUY7fKwirsxUcca9G8iWcN
A47+LIrP71eqRBIj9XgwJozKfbn7Ua4lbkV7+haBShJo2Jb6xzjnkzYJqFZEiaNI
VuADwEiTbvbdhIlLxJhMCLKNbW5iYqCqsYTsdlVMAroiu7mSjfuqD5wP8IQQO1Xj
REDYLEIgzgL+FvLrKCAuunqeDzhZ1y3Ueh4+ykkeySTyvo3k4XVjPLceiiMjW0jy
GGfuxYhJ4xe0117seXyz9P6Y/67eN7vUxQmcvr314FqEhS9cF80bSuUKYp8/ebhN
ampzH03/oZw/VbArHgYv4/VqOXFghBcyDoH/1eQOFUlnxj8Dgxjr/MCVzNZ3ewGH
r86mQtCFCchq1EbFtdguJRNqCoUnO8HGaZ5K3DNmMx4BdwJMyZdiPTsHO/TcZ1nF
Faunm2Ws6gz4bzJSwsX6nqF3MSfdB3BV9z8vARvlJYH9l77IUXRDl2qPSyRW1zfp
arSh7Dn1bIgo3n64ucmwmiOQZJko2HDxycROeKZq2f3kKb6lzZnhCgxbMloeX6mr
AS0ChgC2MhtkYzGYkLc/72vdQnh+6napWUSYJWPcDhB6X9137lM3V1Uym2ZOJXJL
8/+WRMrO+Px4SCuXzP6BLFGhNwopv/fEKlN9KwbZSQw8qwZx2HxOmPfq1OrFN5gt
rC+emnZ+1uFt9vTusFVgUqWVgXif8H5nETjV9m6TE24RcwVTz+OCFTJtY/qfsOvW
fzExLyUj8HGK+jMvoclhmXzYE0E/PHxQP72uF4h2x1Ng0bBDes2eQxf6IVb+J1NE
LJr0FAEpEbWau7lsAGclD7vO8aLQyieoktZLpCkJfTQMWG2MLT0HbWv/Vw/vliqa
DR3r2OnTlTD+DELfzloiVXVgfRkLMhFC3wnn4/gGZr9z4Uwjxld2TCsYVLjm1qgf
3DRhQA40IQgUfwUa4ZTtfREUoUVSfFejyABI0OvxXtdjKQ2XoJ9AW+JmZcM0Sq28
pfhjpB4bCmQikk4cIIxB+tzOw2yuT844N/PBLtod4HgV8Jq1vJ/4I4TDBXb6j4sI
UleSr2GH6lCRgEbaR1uRN1iZ8tZ0OkDuJZVf3PEIWicjqGEpw14e1gHdTSN+FXRX
xK7nm35SQG3ZQEHlMNJgxFyJ3bVFS8B7SdNoeL+Tw1RCRo/NtSSVA+BbG4ujl75U
yvLv9ujZ/+vHSmFm94tdxtIJV9nFOcXwK/CDThaRrVi6WDKw9Mi3gWzeg3lzzLRB
n8VbXXmg/HTBoxpyY/zy55JXYMUrrJEzlbHmlItVuno/MohLqe//OqrIJmh87Q87
0P47sbTsXgOfFXNBxNmcBqFWsIvePfgq2O8PROcK6NeCyjghVBfqdRkLcnuSpxOE
S4gxfwVWUZjoVceWSKYao3nURw7qJXNQZewqNcASvZWKL+0lArraydVUTfelZJGD
rbcbu0xw9K1vCGo+A3UwczStTKLnGS6a8rXclPmLLuo9YTyAj6SmlibfxUBG7yFV
/XWXI9OkQej8AXhtgUFjDNMzz3wHNfJpNYXz+5hN9rC4czxGoNjP4RwA+1RHMl+3
bSsWYm8hfpBRajI+tKxBFiBP8V+++lWHAo/vZ/Uk7Snz0Fh5yZqME/OOJiehRmqn
ky+Kr1H+HGLrVHTheuzM6QjmMGfcQiBxtPVYsJKkY/amyBDprvTQ+FQMUi3LGXtK
ggFI1WXrAdmTYJYHCeBNCCSNCuGczC1jbieCWfSCwmUr+CGNVlyp310PzIbkj+xZ
AGGHABo7rifDAsCFYONQg/Ei/lteK8mFZkFkbjUnAVgadRpSj25b4IWIXFpXLbCg
tOItxAIZw0C+RGYD8xZnTSZzoc5YTMTlwQn8ZmwGpfGxfXoMjUnRym1Ewvtju5It
oHm0Qdh+nO8NT51uWIEf9EySMiRp3ecQUut/1kM0ke8adsVVYGCv52zhIizCWw/M
VTTpYfSuJ5r7zsC8+5NjUaXRhqtgHTc0n+IF4qf03TS4Bn9cNHFmzDBw7G3p5fYd
Qxpbc4mjNcrRiFWvdpHIeAlY4Zga5ShrmyaVeKtKIHdXiohjTbaTTPKTdrGrCfA2
NjGpgFMuNKQe3dag1s8K56IOsY53w1PGfqKwyvXYoQEG4LrbMnnSBWx+gJIhx8HD
GjnpHh4vSQr7EkbecKT126VEHKNq68gMjI5Gv7sEjOqMGwWQJRPFl5bweHL1KR7S
SMihuUASFL//7yRkdmyPmAAdFDUwm7uPM30ixcwa9zLMyATQQz/tuQDSnubw8fyE
BImklEvGAeTk9rMEhcPYa/QZU88tR6VqC7If6rtCI3pSKSAyzdx47fapiCe1un1Z
UFiCPpncp6QKlqTX1Fqc4kqfsltm0DCpcOA/iip8Li4vKVIyBJJ4Doj+VTx9GBfw
ApJlmftw1D/g77AKID2kIz/aargtNfQO+NnYbG7J6oYyE1+1FQH/2u2fwoKCD2wS
+GMsKUu6FGA4Ca9QeLbyhAfxu9cJSRfza5lGBB88X1jEpLkV2YvfP2aHaZlXHRIa
jEdWCvfUn857i8CJNACoPBz2i6Q1wWXdqPAFiH5maYanCfAsZnvb+ZSAlx/tY/YP
riGzf7fOgd3PgB9/fPivGzaVagVMCrt1ujyvTkCxX9ZGlDn/b91TMWyJ9538I3Iu
UUynyPoZ+C7DgeSFl5ZVcdVWQ2ZdUhS6UbJ1efo3g1TiGVbBinegjjuSi7M6nBVx
DKuiFRQJxabtrSAD1aqQ1VK/Mm1uyS/MdV6XYu9TnJiDOhp03GBw/yUoCsN+E8hW
1yAlJQhl7Rp/bcILdL7IvhFcu2A8UxOjeDSHqSvv6OwNqJygbWzvPuH9KvYyigIg
cg2Ud7hLeeXmkdQn2xj7pAoLcVPMgacsP5Fyz8LmmsftpSd8JcpVOsy/L4h+brnJ
LWfD1bM6LI0mnDbKmOfh9tYsTO72zI0yx9d2bwdfKEPecFm/qqa5v/b4kKHC2WHE
EpINv7fZJvYqcsXtgzxHCZ3p0KpZ92waHqFe582qRXcxseJoLQerhMOkzWbI0+34
t9vrnV4YrFDG2NsAA1b/0kyI2mEdKZw0IzaE1e7V+oYCKgZ8Yi97Pi5Ia3GJF+vc
5BYOGKYRNJOA7Ub1nG+0xpvDJKzMXiZX2BGW9doNGUZ3qE1BtkbM0tnO9iSlqqh0
wzibhq9OgWb9rLr3vxvjXBwJO2iBWkltMyTru7EqK18OmiY8onTCn1pv/xItF8IC
fbZT3usr5jDHlm3gjJt2rzurV7X+jYu69CGfVQ2Xipsi5rHumlIUQJzHzqq8aOTf
G8DdN1Ua2YLTLGCan60NNBV0AiSRXFGsAulZAixKaMpomNgSWalWdDTDdrXYr8k3
84IutEQvjQWJDDSfVWntBegfnfdaYUk5VjFwy5xlOB6hnwpuD6eWk3Gr5rOTth/O
DUeTe777FWSqtgG7CrI8n/OKNIlRG2HOsR2SCVbh4nZbviivgOprivZ049GLqDoR
dPaNEG9Kj1OpvqKNGbZzG4KlWkgPJkB1Wg7OR3kCJ/QWHWti7jzMSd3PfLT+KyMI
rakvJ8dfCNCEOKkDnw33us3rlbMs6y0SP5N+W6i5HvzB+KZWR/BrF8wyXqxn/A1r
hpuNThqmxCM0VM5uAISHWXBgyvsO5SkMrQTxUNkw6u9+Qr4Q1F9w104UK2VoAQoO
HLUiSdyXH742bzjsAB96E6uHxI/AhRKqzvx9zuVCXYKW1zAe8KLfhpVzz6QEdjg8
Cu3jGzoucy9D1RKHHfUjQCOzv//sOXPVsiWSrWGNJlX02hf+XohFsCHUE6o5gwIb
kMjOabWmKezPqYqoyjkawewitQHUYcbT//YuXdqT5vxHfhAmTP16HNynhlMswYGM
LCQaYCCFDNSo/o9GyRJoUjISkft90I/ectBhMQtER2b0Ex24ZlUMIfEUvwDXO06P
GpCWABrUvbWfEXQncYzgqHJ1dAXWVrvE99bNJveUgRA0T202EiugNcQwcE3q9spl
oXrFO99vpQ928f32U6Uu0o44aka9eZM+wKCYqQJD2l5QNrGIbqWVCvNX0+/sG8CK
HF5zl04x3cveesOMGZoGwuX9bz5FslkIfmX/MbNH27DODuKCwUd8Pj5h5vP/8n+4
FC9cts/ffF+sgQJZ/f92SPEaHUvy8dhUApNJ1YLO9Tm4m4Il8gKxVHlD88qsfpTf
1NKYs1bQ+GomPZ5nALnbY35WBFSBQgEjpa1xdN6xwHQ/sve9rBeZPYwR3w9j/KfC
mADWH65b7MR9tvwqzYQEh9UdR1sTHeEaybg0+VA0hCWJ2OIpFDQAdUverc6ZAI0s
2RxleTAc80j/M+dmX9SHpBhYkLwWI6rKQuscMKFJFJZSOLBscQA+fVL2IzkfWybG
S//9nyoi5IyFHQr6IzDneino/a9iEnI9Ffd80B6SazdzuivKvVlHsK2cqMdZ0CAn
mbSz1ue3PJXgb/9s9AiC4atotMlAPnA11m0KtACfT4dBBVeHHQJcE6J9/n8NiIqx
B+nrI9yToh5yuwFuz4pPzDtI6XNUzYoEAehX1zc4aRe/P96MxCEVAyGFyRYlqWru
1vZJ6DkRoUZCMDl/U80mvZlzA2+xx4l2H01+vvGlLcXXBaQaao93L6qenRCPUq73
6K6rXFxJ7TH0NoghADwXK4IpuhsN7Heg4CALi+TQY+ts7y30IP5s8wsRnBt4FEFQ
dakNDKpJd+++xgA8UEnyPUmCVmtLYODiyvfjXVcsLeeuhj5Y7poYgXwxUAft+eR0
TlwSe33I2vZxAl0zGXT1WOXku3gIYDlIDZ85+2XOKKTQNuFw6vXqmUYlmGBFp+J0
2nRWFxH4Z6UNN76oxE+ORaEde/kgRRoPwzV/Gif/0NNJlA7TCPHCTjWXADL2uHmN
8K5CmvdsSQtK1iz9M5nE7SZUa5uMAV9Vpr2udslYpGq7+ykr9FSmlxm3SCNO0X3S
BGDbtqdpbJfz/9Ul7IDnHyqeuUa8vEutug4D+IeSyF49azwD5IQsJ1d4XQrPzxMt
yo1T7CW5EF6E5wY/bkVlnZeipST2bAlK2tHxRoZIO0A+1drXrQZTGaOWb+qlLy1C
LYQcITWFARw+zw5u9T5QPK67qmdT1vgPJBFziY5mETkbQQ3dc5P9UxjfqEXYKnv+
1tcehGJwa12fNbviQAkGi8ThfZPTGgrkj6AGP8XWGDcbl6SQv2Yrs2nPBmOAwYYW
qgHPSyFAJy5aiEc56FW7XioPdB/V4BM8whmGbiEpQ6286j+SickWsndh/L3EmRm5
NrynmkKpt2WI6RE18dtDQPHulQpG7QYS0qZVDuG+FIMmE75Pz0BadQuYf+G+gcxR
hxb0LBeQ7yK6DcOmn5ifXu2Aw2e2ugliNHP0cUCPrSp10XMiinwTfV5isnYZ9enM
bf/v/9SqRz1OQbW5dCx1zLhbiEvPDSKg8pkdjitr0iwJO0ErhXVPOu3QEVTz7x+A
lIxmBEczAjbGQ5RVrfmWkT9PW3iflAyKRlViMQckNhoNetyYtk2jiKihDjksIcQJ
PKsnbkCkGmF4kA3uBvgxlbbtiKseGEUxSCHZynMSo58+DjcP/+ys3FqRQFmU5XWg
HkAlGaEP5Y7QROQHM9P63yOowbHyF3EHvYbNRiq4xlXMlcvV04Owoeloug5e9quH
KqbzScIBRkPE7Rc/a0DCunpl5v5TLeygfOfqze1gVBtuZu3j6JiYPl2sAWRKLFNK
86JBbxcO82DOJY1rJhvzhpRRhHHLcClnw43DeMn0O3L1+taTXzMu3MeNhdP0UV7N
VLYT0/q7aCVJ0fIMzFmXHoDdPMQCF0UYQM0uRfwWQuzcNCIQoLgqru6ulkP83e+v
ZJUNRe1wdf8SDXVHt6xqUEScbdHu7JPQN9zJdawZ2GtfcrO7lt8PQ/TxgRxEJRYa
ufFJ7WBRlP934PAHFvQZtlffHbv0o+y5YJ4oO//f2enz2RLEVmlD+PXOlMeHN6Qz
v9BBWo9WCHNpauaD9aYrnMPGoacynwMksdWnYCLFirObGclTIkN6MoWA1u3fZWrI
I5BbFeRgTlSJjlJwK3MbgXshsjA9QLgeM5jXt4yk95cs10opdRiBsfeFw3VPHWdu
1LC0DM4/QA1QFuFL4m4Y+QUZ/2C8Sg189qqfVAtBgLl/dujcLbojqV8ijU28lfG1
J4WbqaIS+yqT/QAixnY4n9fA4S94UFfv+Iti60h1Dx+UddaUgC6xjPfUFJWoCm6g
NEqmke6j4jCWDP5/54/K88d6zneVKe+WE2yqyC85hibcS/xJck5Bn5qUtbhvJ91G
mKVTskjdljhvEJMUNuDeUG6l2lo6y1b2tm5eUnkOAGcg6GISYaxoTqArSpg6NywC
9DdCFKr+PuvNvtJ9IYCwkDFs0U7aQhf8445im2xqKHI8d5NLJlOKRGdtDosu2Nhy
LvTZDU0MRdg1apFKRFmD2N5H7u3tM0t9vmnxOAIhtxX8o5Daq44ovFiWd3hpgBgD
YO+wIUl1aBvgYJBNEP86oGHzcUTSgy7ySCaZE2nyPTfPSdKcWom3b7tfoPL/vRKC
H7/yeA+oBqFVKFEAJj3uBiDmG7jw90YFoGzgIJMG6mzMZ1W0avBOALkbNvWRGUlQ
2OiJ9R28lnap0HynH2mTAc8qpG1KNDwes2PwIB/5tDBjnL1JqBxaR9YdRjdo8JZH
AtFGmJzsP7ck7A/pwtO67SvR7xotwZDrZLgLlUQ0AhwdkxOfqxNiefXwJsV1wkHV
e4MfrcpeVZ4tgxuueZQ7MbsOan/491SqI0fZdaKBUHK4GdusP1eAxwyQMY6UebjK
/1ZVfTdZhVmhWDcLoewi4OoMDZEV+wqi1oec91NnjwNhXS7oVg2GvImrzq/XgE3d
2D+VMVHN1x+H72YC3JU/v90XnCDpvT3aJb57tBCqOPPehLS1MprjDCtxbCJY4MIN
pUlagea8566O8fI6GQ9acqKNdCU88Syk9w3L/FHVvJCwHGXqHTkuJF7IOTXQziHy
md8xUNCFBoNcSwzUNnslQmVWmuTq1yL12/KzUDTyPb4SIRXxHEZdjMSCqoxnqIMQ
B1BPegzZpR0Pruj8ypF21E9oLoT2wXHJWTUcl98R3oH+745YtEbUbwKrwZPFWKrC
2AlYpZFfujjS39fJW5NLDlkz13JC2acytIFi2YEpb9Bbj3xadx1Ja08aP9yhI2O6
EeFOz5OqOtB2LERj36bsXGBgniB8RVr8QthPZ4L65hMZHLFrrYyzf/4UJhFIImzU
xWYJN5iHBxNDcr3yEPJvcid+tm/+of2k2a2uJS9HCCDQsjGn1jBzSPQUuh5KnUY3
basI33f2mzUdhjjuHprTxdluFmSpoDCfHJg8x1m24015lSKvHC/54soJA6mzzQLi
cXPIEeCzTUhFJic3d+1WbHQWBk5TW7abeuKjDwNKVTnWZp/wMbKcodPv3MlHdz9v
qWvS7chrjtvdaRcp/QFBaoBxjchdByLew/vjkoHicHgH8WYT4NswGcAt8nCYXvu2
WEOIlHv4Z/OLNX2V+s5x7OfSMeR7uXCsktnbHbR+qpVbRCr8hzyEmSN1yGhL5ZLM
1A0PbboVHikdv68xKI21hHBKw+4SwXbkmOXf8S+Ms81164Bu0L5qJmOiiGxn5Knp
hai7dxAGXZCUjZin23xeuCpHaTISF8AvYIhQbi0dn+rURvyOXN8JvgqlaE5lNvw6
RTTuNR8k5d77m3qXR+3kRgaNVr2H5wfP37RIsQwoPRE5vx60k8CBinkK1V5PqrZL
+KhQyWgzESTWCTK7xnciD7AdWbm+Zr8eSwWHHFsLTOx3Sf7rEx5rvM55rBaqRWvP
Ulwk0v/5WGl47j35D9OF8/ZGzGmg1lor+dP7n8bPl61ckYJpUskADFWIrs8oIkDO
eIq9iwBl7IlpuFAR9Fo2LRSoEFWu1XvV/Wg3ZlD0pDT4hkyqgfL3DoT3ozDiABVZ
S5HRYRQxl/EfCJTV1f1WaG1hgsuLAuP4oCIHL03nJcC/nLpX/T7kxrEGOHGGKDZI
DWhBRcmz7/cmoC7KRbT/8QhzFU09bNQIQKj7yenKROQrbPPB5RYqzeMbpt28PKFR
7zL+WihduoXeJIG6Mk2bnbV1P/LOaRACWJMiYnYWAr0fMaWtBVVP71dqMVYGn7ey
yep8/Le5aKr2Oql36nWVPxRpTUIRR01c58co8ZktiZ8IP7smykJOPHGaLLk3cTZr
DeMrGuDIl6gZw6FxW3HQim4GeT+PfzV7AF62OqTtKcZUn52ykzdPChvMX6HtiVUD
7gVwezxxTWy3YJ2Wz6oNRNd1pCI8EP1ppGn3yeaO1K2Pvg/YzZVB+iFQle0KV8o4
cn75j6HIKtNtTQzMOXuNuoZAq2c48Er5mnFDHUPIDxbsjvzorWCuNwyZO523jTlD
n5BEP6bevkCdB9S6B1RhAR7hXNQsMaPYvpjyuS47e/uWvmGx1Y8zS3kM1GSMpar1
cfRYrsOsWAXpuWzonhTFxMh6yJeqarMW5asK/4tEFAqrIfVXEWi3v1ADyk3SuJQC
cvlvIOkg9Rviy3VXibAUmfH6kNvvciIqWKV6KDoPEqLeC7WRsbDq/P1BMOF5hK0p
6W2giEOX0XUHt/YkHj6KCuCAUafrifqH61aXE6xXCHyNdnDuHRAayDVuZDesNiV/
uw0n7P+0RTK3yhmw8TBbOopTRul2LuzgxogNWPRKyGK5RWVfkZiKv/7nmWMhYRnY
PlssCHTkgkwGsesgupGRT1IJaNHiRMEzHLEgitRIUIEKM16WgwRnE9iYzF7Mi+fr
EUkMUsrADjsEwpszRWt1qMNvxaoS2IzD7lQteKkK9kWrAMjzkFxPays10/lpQlGq
X+YChCQ7jdg62PzS/xkydtOtjYffIjgeQ0/Zt5WAlydQhb3J7h51XMYSNFfT4wg3
m46G2Idj+N4EsSeHNcmxZeKs2gqMHT/jYH0lEmdrBYkUftUfdIzVAYzbz9XtRwwC
oG+T0W9IZoweiWBcbNMxlZ4HCVPWLKf5F9G7i9UcvRpC4sPWMSFi6k16bS2jGoZa
j4tlWbMYzxbs18bxs1lZywxPaYb3IXmhhkRp/vkQj4TjgU9drGsiT5nJKdKBiVGR
kFM02S5izh32yEfP2zvICavhK02+3xvtBHyvICxmvnhyC/k32GZ9nSqhYJw3/LxK
cD8lwdGXAD+Yo53Cis6vGAjchf7qdsZ8vPZb/4dqBJD0U5+iGaVbYzd8AW6xD/J+
rMfGVR1EsmStiYbbMI5BKj5aP2Ac7NZ7b7Sg3FaBC/poKjD3xXq0sUdiRFXbzisE
o7iyQYqcpgUsDyQkAr4Km2gszVCi/pPSB2bMl/zIIacVq/NucTY/3ag7rcbAAZSv
XNUFwo9MU+nk4L5g0C3h1hYRkSg5tAUSZHHZEvWleznjINiQQwTawrDYGn4Qi+Ob
olxLi3obNss5n9T6uw0z+oWKoQFHUhgNdp9xQzUiiP2VoqZkLzpMiYmuXJuWp309
Hsm4ZzY4KjW7vomAUDh9w6MLKFez+mzXqr8TX8FVHM74OaQNGnUq0akwtucZMWX/
2Mdd7Ahx1b1XoSZ4LwfUmazSFkg4r7d6mb38L0KPyxwfCs3Wkhhe+Fd3/OpjvpF2
PYBWBKsoFXuqVnrKCGL78uxZk6YBtdaSn/vcOkbokExMADagbXfiTdLIaUWJ3xjn
hh7vu6US5AWQ5ICzI0TDkk+ffhLvohwtLeBDeZuoCCr5IrBh3VYGkC+HXSixJlsD
D4A5LyvQ3VtsFFpzTmZlCRG/PuMr1+pdKEvUYZsKdgWF+7RmpoW0tXTRzxHtIdMd
l1X/NruSVnFvNCNSjU8vikBsFzwN76WamPQGkry3ArSa25amnXrDDki2Til0NN1H
WnvPXMrapdQhhVCgA5fR9bPNLQSiywCfy40UHgYvxKyWYekx8ZUhgMfmYd0sLxVa
g8GqMX0FF9pjbBW7Cvn9jxsvnlVnQMa+BfYJeAp8MRXFailWifWz40qKVQy8A5Qa
EN2fl/41FhofcF0+LDcK7WEPQM2P//+JW1ehizs8dOZO4vMpHh2WsHjy497vVTG8
MkQOjHg9YN6GPlsAf5F/UOS78uX08fgqSvwSv9VhY8Wv6ZCS+hW3j72F0GIQIELn
CRMLzhRw1Fal6y5HHyg13QJXS4wvAa9NOngyYl14ny7EHOXkl/7qwkDYW7O9JhLO
gfXHYwxSD1k7P9ipJ1wdnC89enB7dphBmvkZ3EP5HYFN42spxqowZyhCW4NSnVZn
tpir0PSKlmrEW247VmdoZYuQoYtOdt5o/iGG7dX2AwaSxo8svZvIyYW2eXsixKmP
Wd5z3t0dRdCBVQT5n1WEeGDJYU9AexGUc/TepPsjjwKLVHPAZ4oNh9DNuQxStjRh
Gh2a4u7mNlkhLZNs6hL0IJskKKlaL/zXf6yHG/00LrsmNqa3efA51L4/DF8a8yLO
94CjZYg8pT7933guevJckqi03WstRAEWOAcOFoFngmDgx4uNmYhfoq+mYYYVg9jy
MJGNWc3MpPNW8bzqMDQKsma9JwdOkq8CapGLYNFvgyvgXMWKaomCEl3tqNZsL6mF
UqVl6XgohecnBOtjrXnUngU0VQQGRAuKbJcVkNeF4ouZwHewxi2v32xsJtL6Vg5h
dJjwVOGE+IiFEMENJLf7XRwA0IpgC8qz6v2GGV44qbTvb7N0G3V/ai1bxtWogYRM
2nZFuT90p9yQHbQ1eDHvjiBk1YgS9M16AJYSmgzEiboj6NW2a/JnAwujo6SFzUPa
Y+1vorVl8VOmRhDr715mEu8y7LWHTWaE20x9deOnuqgAYcvdBbSjXT7uiF0kASBv
RsREbUSYwj2lQzqEtEMC4jSegtG6ECGfvy9gVvw4DZlOXnyvUNQcO9A996x01cw0
K/zhlsiub4z1OJ4SgJZNz0o9YQ2gUGVowqab9yzBHYXp6bveaznvm9lDNU3mzx2i
FqwH/u5aeDjgTeLjBzXKSigV8EuNUOtjSIWaUM8XQ2L4bPNhx0nTTnfYoIA15eOU
27YToUBs9m46ECVRAkc9d+PjnJh/y3k+3r7MA0fgPudjFqVVyM5sRJmbHcVv1kOR
RjPkhwxK20L6+ZuLvZ1CD+nXbzu6YZYx7MWCD9U1XT8T6w2b4YVig1ddh0cFHGXN
/w2q/UwEzdpokNm/rQz+wA7kU3Abm6iyrc+ixEGElvEVHq+c52GGkcSeZmGzA4s8
8Vfz6ynGQHWNztRDaX69yu70GPjOIavREXfdRJLo4Qc2G0TmpkLdqlLpvQVqntJ0
+K+X6lkpMuAbK5vz2e/eM8QL1cJdmxlFibzPcolW7P2+EXZPR+VQC1/+Cj/lig6E
JSHw7UxDCWRP6C3IfwLwWQgKRYDeP902o7iCwBDoM91NZoybmQNCFT0MgHnF5Mky
v5FB/qCV5Pw0xa2FGm7l6PeN1oRcAnkff89sW380FjKMov3C35mWYp4AQTaFE/wc
PFK49hOAy+V9ID2nPbeo7qXKHLXomf5ubMy0b6kqkiJNB0tizum4ToCmWlrQ/kgO
9uQ7bO3bllWykzeoS8iXGUSeVMmu2jY4kew3B8Im5qU01WW+u7qk+XnXWog8yfj3
/hWmoR6BHmX+D5gvcxVKneuu0FCSgX3AajBRy/z0IuYTuuRRQCvbTsFB/R2pknkU
DiR/3vGdCOu7c9lH/ctkG/D59UjSf35/mK4xIRKOeN9Q/6eTJwvdbdXANDrzzWkE
Zjt9IzF85UHdavWZxEwuD9IayLxWNpYKiMifqmNuaZrsyN/OVj4cWQfgp2eXICsO
XG/LwVWhK2yso45O423adeWoki4gmuuS4KVwT2R3j+f2lUXZQ8ycGnbMnUzwjAUc
E8C4tRZfrH4Dm1QGorT93ZxqZRCHF/8z2WKt7vni/l4wQ1Fjq+t3F/v8rbuIrEkh
6L0nzMGP/5JUv9rgMAtNjaQXTwfYuufDrvFSjWr2MS17BL5UnYbcziyy5XD/M70/
R+FC7YR+s4ncFIqYUsPhWSfRKcP1xkki3rT2Y4UtKnmmqLcRYO2NZ8PnvfP/LjvX
rlDcIfUX8igEhEnkiq5sAiEhg40EB4ZYDdFJ+O/yGFuMirnT7y8/R+UMBuSQ57a4
31Mr1Q5xeZp1egvHlGQyNeUQIV2t+lpSePFlaQEsFMMIIZGgXpGdUYMLOtnWEJIX
39KUJ69scygKW/tdGTISve4iYwZqUGSJ/qzjZhfdirOa/pdNVleqHG7yIBHt73Zr
OhjDZ+WZPo1WtMk/Yq+ACrLyXXSJjGKh+vAcFElm54ky6MDEWUmoRgR31YiqNC30
Z/wPS8OJ1oOXKaFCLplgfAikxDuvBi9iqKTuJBdtRnEJUevUMZecXNdfut94e3v9
p8Ss2bFlmpSUWTY9E/uqttYIcJ/2LcpL7zGzWsXyQTwFEpZUKep3p75yWkDy9b3u
3wHfHU4Go8FJrb6t2r+yEYTHJeE+dZLTSu02WjnE1TuDomcm8gBdbTMbJHqy/syo
3EpcAEMOWnuwfO3+Ac6JCtK8cMh/0l/bVSwLygzCSyiSncjkCtyu39IQHp0Lgi5z
5FOVTNMlMPwvDEoIZFJoMbrBdysCW0FLN7oaOb6270ZuLxWDrogQsWUpCYiwfvT9
HK/RpJFkVmHwsEm7yhNw77rLCN5lxbfFyo7gZ/lMcI2uRt5eTUogq/8t3UjthC8N
YymDEoyOzgDaGilhATTiQfj6VNcob1qVv1kkbo7N+DVNjLixQkR0fLftE1zI3VqJ
PFCIFRGsNTwePVL6rfNnrsSNm7GHifL+tePsEUldXzW1nssZipYyWMG3Ly7RnZRW
PTr8m7jM9f6an/6roPHnYEJq9sfHPGRW9NQ8XEOrmhRBJ2k4ekTvReo5j36unl/m
WkeQA6SZP/8tzz7w37u4fsrpYwQ8Fcle81rme/I/6E2dNXx6kJQ60a/hlPJtH1Mw
5JIF+LBKyxfPCYAtrWFcTjcYghDFHax7f4S2hAa5bdF637CIQB0iRdZuN1UlDuL3
lclcPvjrOCyL+P78lb0qN9KwODcq3HxZVQA03r12JRpeRY4tjimOGr/k+EJu7mOk
9MJZGv5GaONgFHVxnJdfyyqfC+MlPMngEENkoUOZLaf96FDWNerjTD73pe4bLIwP
vmmZKRIfhNtDlg/ITbd0dLQ30k/Cv3tYFgDUmZWcvkipcoEXpE6w11vCczy5WiT0
RtAdYf2KrZV6wmEtqx+OFm9XUiOm/50gxcLT41cH+uqaLfwOVi64+/YucbRew2xG
yqoIQqwhxp+PlO33SG62i4BOu54/nePB/2zbiWnnmRqDzIUPYRf1uTCodUVae7yk
/n5+unzH+/+2q6QOnwS+oXSO1mlQRTGFj28rGazzJksHQtT/eKAdvNeItYR/YiNg
viVeDNj/l+vDWc8JS9hSnfeSwN5bIxwB9aXoqp+LbkJOMuYK6DfKtOdlYBrdpvow
qsa9LSutJVBtYeD+4USieL25l5OxnuEaiFt+/zXr7rty3ZO9WzXn8bJpPLLdHQxQ
METLoi84Xh/wniqfh3cLloFldNR5pcJzn8lRWIuoQ6A2y0YJgvKCfG48wlPgBxdo
NmkClq6P+g3PcWJKsgLojxTmNbm0SWckPlHUwZEqKGuyWwZIGIl5W49fbmus5bXC
Pqp2nUXefz4nmle1gN3Ssk0o9WSe2Fdl1Ia5BmUucwXpvrRJSd9qHkpbcvbZZHFR
ERzyGFbfXY+J8cZQfju5GD+vStj/fT46/TywXyzGmkPABVO594Un2FsnapqjPYW7
98soBzf/gPMhuuZVGTLF9O/qD0bpFQ07A662sRp6LaTYWCrEkZkSfrTMNXHd0j+9
3TuwmBo8DGJB2BSr1TyE87tsuDGgeRxJSJPIXLIElRalwXxWXNFOS68ycDjvQi5I
4pLoWrESbqWpBoaaLTFQfCPPCAH9KhW2JaMlz+u62Nt5aBJdmMXcptdBa7nUfrIf
Bpy9gP3OxAXTUM1DYm9XeYqhabt+sSmFCvNZ8retO3llbVPlOZH7Jas7lXDEbxGe
HTFoNzMwcCHyMnxEFjp2DomprT/YGFmTyBTmI9vL57hf6RGJr1Cj4IhVgU7s669E
Pvc5vsRvHbxNOyN3yzCHV8gz+MTn3Q8MffhFvp1ZhJ0Lm0a96LIp4JxBesid/KvQ
6EDP7jDN69QRVJX6g7Ckz19Ws5G9esWw/hm5FtKR7FiWQsSll3UQlMW/ud5q4XIN
coIuFU2J+8JwWXTM5zRrGVZ8ayVAaQV6LgTWoALvbKlNq8hLNB8r4nwmEEN1DqaF
deSDDK+IHd1qf77WntIUPLQbYi7eLdxIEXTATgsPu7xw9qD+/l6NQsIpJLm5ZeUs
apZuoeYDAO1mOhRZchVmLVBVEAPVBGs683LOl0G4UMwYfdnnIRjnyhh3HNjOXJhZ
Dn4FIh2sWhr8JbhvOLcF74HEAifsP4XcmD1KaztJoJe1roIriw6r3t/qZ7xO/QYK
DPP3Zf5cU4t7mwzdA1JN22isUKVNLfvfOyhJTTyslTifx7ogYgYBcP7qM4J/4tIW
x+5vnYiqJfPQbnHgc8HgzglZ6rGFiN1ob81Nvp7HB7KPqDbuTcym7TGSQ1A0+RrC
GTkcBYm7YuMgWC9uz+L7beWj1GZG/ZVQWhuTXuwXUGcvPtsKKj+mJOOAjO1PVCgo
ejzyspjpe60EnXq09+pkKraudu92nFsDYkcJcng2M7vo+Hu07KpNJUfDKnDV6rE2
zv19Di94o5nr9Pvd73ZmPJ3VZKKJBZDaWYZCIQosXUWgIItAMRaZndAApPgGKFwC
RFCcpXd8jY/WT2qHjWAjbIL3l0YmBWu+fJ7vW9aO9fPzGNMJaDYCJK9FcJL8HXAg
NwFgyVF6Lp70up2OEsfOi/xEcxo7y118sjwohIkWlGJ2wPf3HB+s7X1EtwvPGoCM
TO2fYfQkPIDmF7Q6xkWstNkCHSbRNxlNg1+LSTJZLtlUDgsK5sw2UakWmPNJ4/Dn
9D5l/iCl2OZuGD6Ax1wLEcuhqmK0xg/MgLadEXLYv9WNQ9NnzJ3RkLtg9smNzR1P
izNsfoMq3QqYgTyagWALafAuiN308srdV3KD3j9beTBfehKibOo/kEdrHweTxI1/
SOlUWuTsTxUjcdf1+tvkCchEDPH1+nid/U8L1g9/wckjILIdNZEaBLy7NAD6eHgM
11uSyoE+BbFrTMiOcSWQzrkPCcZfghdfwi4KlEY2QIvbdzYTbtP6St/dMUpmrUsQ
MgKNna8//nLd5FkeIIb3Xtp10ZC+zQ+Fb+gaeDue6XRuKwDpm8iE/mBJSsP7LhaX
iDo+uhslSEtnD7VUJpHzAKJCMYLGc/RH5VuVpPIiPCERnCD4BCXlkexbwkgN5GUT
u3xUkvxX9oFxlzHnnqwcoh+kiNp4K+ttRJPU3ZPkjhlo675Cc9j1HwmsSP+Nvoqw
vCuj0M6+Cy4W11VkiENv5s1uyDLmXQJvR/hWRtobpcEvNhw+zRIDWfa6UZ/Rl81t
JUNiEHC0vMjkPahpj8Go20WHQypWZXbw2SmDSXJYfY5RX3J9+OggPX+lOSua/iMe
LMh9E+3Nj6joY7VKCyrPWvCJIitQ4W11X3rrTQDUGV5q+jqDJKVt5b9uyBX1n5j5
IQ06gn17ymQmTgtHOhpn1BtHpBYyRyKx24bUnEuSsUUbsStGe+qaIGpUrljr18XD
ynQ7+fqHa+av7NZUK8leyPNnJMda09WWARBy53CscnOl3IGVAAvYk2dlDMzwUEpM
kHj4VZswVwSl+V4hEq+MwAy2CzwrC0+Bm1dEwgI0wtstfXyOVLVIifUYtV4AzXea
YcNV8GM1mQgc4SbpQ1+WsgQWGns0aLjYmPu1G5qjlmj4xp8tzRrPUHPuscLwGgw/
m7f5Tum0bBGB0T5ezwWU5nWXRgHi7lsfk4CrC9vf9xHKeXeBFCRxSOed95HhsgTy
xZHCkWx/jhDHhmyl9cZiuitICBa3vMdtcqF+tAppz3kV04Zk2MOcs6Ah455N+IFp
vMz0smZHEJANIH/z4+4a3aqdDTcl6uEPSDqcrQyHT+AYoHIjXFuaCBpnSiURTSQU
fX7N8dtGW74q8y3t5WHs/TdqZagjfPP7VRw1Nuckl2MoqeLp5aFt3BlCO1ojLatE
X+VBT6CP8xw1o2j6Z6kmSehOs5pfN+RSKiCurcugbuF+gE97fraBIQlUX4k/gp6/
0pfFHAx6jZS+dgYyMvM7eg6S4hq2XBL3JrJFdoq8LS9PQ0+DdKY5S7IiD74FDExH
bxvOKzEzMqjUSsNIFupui2GErQJ8QE/GxU84f8/reDb1lwTL+WiT66T4rEPj0bGk
k33GQXjONlN27/jzGeBTeJ9+Mr/Pd7QTiyiGSX651Ho1neUsVwWdheMLlxerduwJ
tJeX5igC/CzlmE+yGMEwtLZKwyPBtS3LIX24wnOBF5BhdufnoSgqVhWWy+qz9cVb
mJfV/NOnu/W5e/c6zZoUKP96a1MwyEV4dT0SZkaos807++9ZNQNIrflOok1KOBRV
eaaVLwV0mR+gxt6+7gCDsngcuMwszh+orv39d8zyjJbMN6nL2HXXeYCBsaeXWc/c
/34sgEBUUbjEJaWjYJL/iX+aCPpwST8/uiPfNPZ9X3y7Xu3LeTRTeyqyUqVJQcXA
M7qho5XHgHgn23XJLAThUgDH3OUHjynCi73wjBPKviml90u5khmMLOVfHVuxS6PR
Aq29Bp4BDNdSKut+Gimi951JBOQuuT7IFDHl3QP3JYcEXl6Igkdp2ys9rlF+3VJm
Zl4uuBtbBh8dccBEAKFt2kP5rajsYkSsM7C4yfzdOeYlpawpjTHfvm+H9Nx0aN7Q
qtLmLcbWCB1gbLSy+9tdpvO+/S5ce1UrM8tEgiotRJ2/cJxLKxwJWcJml6feHbKH
UilgFoaF/GMCwEnj1r6beUJ1nm8/tggMGrs6sn6uraby9JaNf76k4a8xfDGBVWQQ
z4ToKPPFWlrtPJgoOGbKfmDJOGGPJI98r539ZsUKpZgC79X1MGCZ2RJkeG7xG2mj
IWFU7dICg6vjcLy4w7HVF4Hgp+jsLpB2Y0xCKTnQXgj6HcvTXQ6/Izmx9EUhb3Y2
sFrRqWYiSEBX6rZFoymHqoMOr6/d0vuvS03mToF1m89ra5viSD4y8qhjgwQu8+iA
+WsKmGU9iz2II3KMuwE5wO7jlNVaRODQ0PK6yRFc9pNYqAB3AFi8hF/VfarU0ug3
/k8Jhy8vNGN+TK+0hR+lHS+9Mk0Ehvjaa7cYTptqq0QDWo+HBvJUhqY4OmOg2f4G
Lh8QeV0F6r0OwMOL8PYo4tm0zaPAWeMnTChlZf+ULUx6YuCCgoqHuTPtuvGbhY1/
sXeKjpBKQXb3QSl/WPIWV/KaOjnuoFyrOieJJIk4hfvXp+w/ueoOCZWqGRZ4yewj
7TRCdu7uhUYTXTNjW1TY6i5BavdV/3DzlK1/PuG9H91Y8UHFwTs2QC8vGaG1JitL
sDkR4w8gMzubRdELKjO/MIYeNrp+RSnQDryAQBcYKM8EMFXzhcg5Ug3v8XIerBX6
ijs29HwWCBH6IsW2jCfRgaLLyfqsUlXL68F/RunZ9hTk336g/PirIapSqkqpw5Ls
xVfUHHc7n1bnscQRreZrd8t4kVdcTe9zHoTjHVCABfhYQNzS4rf030quz/u8U+QC
OAmUHwurvkZGQUnu+fvGlhY9oepAPqbBhCR/NM5PdNNjRQNNph/6BCLYkGE/o5CJ
4Lykv2hCKhVasE/AjjR87rHvp0omMh6FbwbChuf5lQR25VjsYroa6Hmx06s9IXA1
sIpClozdWkcKIW8xYi/q04xF29xR9lSMT7ADLK9SUWIQ6QGJW2OZ4qBVU6OgZr5b
ezLMmIyHUHuyMUHee3bTJ6/5yDwpTs7t9HvowzHzeDlcOD/NozxpzkZgZjtaiM81
9DRuiQK7YzcI1TjPYwEw0raBeXMxgklhbD/2YN6t2oBrK/JYMVevPNqAPxe/NaL+
LT1Scf2pQMmDxRYe2qDGi+s379cXxNp6Jblgxy6YibXsNVleHq4q9DXZcM4HPLTp
kku19OxXOhSeDLbgUueM5YPMUgWXjH1U4LLUcEe9yNN659wvw7HWWUgrQWymjVEl
dse3r7T9kDm31akRdOrmkqizjB06enkYUlYEBHOhe4nw+zWoSaQ+upj2yD/InGwj
31S4RbLalDe43YkeHrDZmpD+4d2rI5T3hIP7NjtzzaBrOpTTvQCVfq7VypyUUYWn
HFsmS8EXG66bVcVd3PvuT83WgIsE7TT4LXD1nkzKnu7zsR7ioYwB915Hy63bgV6F
+utaoApE8lRd8F/gO9+jFBE1KBUWzjtQD7GnVBQrWQhDZIaFQ89BxB0xXtO/7ccv
sQbVGMnzvOiTO1wQeUQvNmXeEqK0VvxhnttvtOCLM22IhZi3yNaeLVvPoSAjNXNJ
n337ifBM3joCWxow2j9i9P4qdaZ3bMYJ2i5rjn1I78MoZ/6YQXjtOGA0tVYQ1P3/
wm/pOGXcTdhR1geEI+p31FLJaozlpjc5dfwOlPV2oH+HW/DM3OtezQrzMWYgdWDy
U8SkQvfA/j9Og8pcV0wX7pkNOVXL/hBBOMS8Xp2hGprFjuRtTbHVR+EPgGp+CBOd
h+zScCd5zqpRaGpjPs3gVBjokYuSKYpMF4qJjXL9XQ4djc/zZQW4+hyRUNNewg+J
21NUL4rqSoqXUTM3E9fKkiM5ujvpBXqV/pluQQ3x4NrTGfZytveCEfDv5tsbx1xR
Zigk1L4OxGR/3n/L8cjtkRUvdPO/ByNfkLy6yU+6bcLZ36tz1iMSteLzhAQ4MAsZ
r0D/2Jr4Ys3ZW9aGumG//BxeqMznB4J+hXngAwVuTX/k3xBCsSxPHPa6YSVd+uEi
IqpTSfdbdK9sKAuT7tVcM5KQEYq0cD/mmdt7UDleeNnv7Iu5rcKqcnjRARWAha2u
OidRIHY9Hzq1jBrqszJr0QVIxOfvltM08WI7Z3KiqD0rLQJkQkJF3XUJu+QxndU5
u1twiVI7T3swf5eHwDY5gGvgWxkFMSPhpNRApFYlALo5/Otp2Ck9Ht01/bDrzjXT
1SKpyt1r0Fzcne/yzp+kp/ho4sFEa75a/KTxQAaTzW9oA0uv+O1pllUR2iX8EEP/
IzhjwOxh2ZKeVl6gGa/rvW+k2jmarW3/AH1D98ydJgWJV2r2e0Qt1QdjqdHl1Wq2
ZPM/nNo61JNWy3i96bP/EhxWLiXtsnc9m1Q+uiUIZLb4N0nHq68k3+e95oqh5aqu
wMvKdQgPaC8hefXZT3wZDsKPDv9xNYtmT/O6lZC8n3pPFqoqK2fr/katMBfN6Wbp
c6tGKpqWixgSwv1a/lVIA9H4LLb0HPHVx5pMhedTQ0Hmzu/ydpefSPb7htzt8WOU
xTopauZlZINViAh7VE5CGJN4WzsbZANHG9Ve3u/UEF6Op1iOUBjbdbItSOwESf8J
GSUJw8Fc6GWT+qfVrNY2UD1PoNyKbdeHUF+2MP5TrAc6GvNY53puw+ezhPibmNUg
QbjEAp8fVG5fSE2l6+OFmiHqqFTgkYjKXwJcT0OcNdD1QEu5JVxAzKRonhbv7AQM
wWgIYyABb8eBGjFG03VjEoRM49MYkE4ldtfxn9QI2yLMaJ7y+EOSxVs/3xrjNGc/
ONYMs8haVKmmG5NF7bPkBUAvUVOQjgAt0zoJPoxjYN0tqkTGlf+2tTGBbzVpMLA1
+31cGQ4V2Wg09mQK8vzbGwiwSk/Om9QdivOJ0RO2J/40GpNgctmMN9yYy2n+1fyR
hwJOBo0ckXHTkYjtzU8Jb881Jq4lTEd5elH9qJ2i66sqJouwTYJBIfDgPsUy1qMY
fSYN4NVUQZouvlwI20X5XAv1wIZULHqFwewc4MIx/CjULwLRvKma1bLaIz4RK8Uk
o1OXNXytYxlXPqKhANg1T14NFOIcHwQM5mIULvqkuA0oELlmA/fbAC8i10g0XxH+
LV6VZS1SjZDKp1Voq24xeviGJWWGr1ngcmks9JtfH25O96melt1y6m0NXKp9lj9d
iDCCijpkIzgOQQBIGaI2S4XuhXl1J2MOLTGhnDneySHK+uloGSymLXzgCPTdlhh2
xDl96EnGeBp4b53DIARbs2Qlbw//E3hZDt43Yo3odBFXS9ZpnapBlMBNsk9PGdHA
x2nVF/iTWqSmNJGBeozuZAqShaptAWBYYlCqBczAhs0euldYBSyqqqMizyugjtbE
bCMBKA+OyzKGP7Mcn+XR2V0E1LRC5NiVWyBmwBk6zv4UlZPxQxPTuU21uDvdomHw
VPjtZOaAZ0QK4RJHLnd/p63JKfWj5uPaV2uLtNPq7JPraFozr876SJeFZQ6+ESbV
ClHAMpYmAx/NEPCPLyasuoC8MaGjyLRrf6r79SkI0zZvJ/zNzloC6nYUmtSQCebw
pKMwsbpe83UJIRgYXw8p71qiPwfFxqYE5dIWoahX2yae3TIRk9JnFUWncdCE690q
hEMBee9DiXZKUr7xzW3eLhIQtZBsj0UfUPNYiZVwFtu4WHeddHHSiujMFDdcgmJ5
vnKEOm8TA+dh53QRc2kYSBWYTNJRlUFiM6oTYFu72VMZAJJLKVxrF5zY966GxqDE
360nCf8tZ7YphmkTpG7CJspu8H/lpZ0boCqyiiWYox6r1tV7sReApJu5ndIY+Tc1
SJQae13ZqXR/3dZlCs7De1csVLKIwhy3dR9AG+zpj1wK8j4t4hTVBmi+eWvQr0Ux
ahLFvLaFmD4kKfqD+i5AAsvPc9VJhrhbQZdTe4HxqTNt/m7OWmWj4/UQVYURFSZL
nhFesvLmBkrvdU62c4bHDuhD8C8NIy+dxz9C6Gk0dZCzd+IYBpx/sxIcJLFmIFR/
x3Mx0T7rna2H6EySCRUz5jQK6WaKuRpvongAuCFBiTIZNNnr79JvBFNC6nJlVnBa
Ep6TiOKqliIcuqIpx/ntx+bTFP3bNxLNhGgRO0TksteAMhM3SGWgIa0InN1kxLm/
O6XXtSBzwwNCpdr7ZYQ7cagHcDlXaZ4D8vXENHX1c6twBkX2FwvLJWIUGv6LalDL
Sqm1mtMhbzntTVkEMrq1mD2d7kUr8s4hZbA4Uhu4Pw2kriivH9nnDOsjLerTy1Jp
TlkTJ4ZmkmtTcp5QQVLhZ15tkN8GoJoHNt8EYUDZ0i+naIK+GRCzQHv2vRk267wT
WmBvz8KxHx1kEUVQovxiohR4wTjRvDbiFieEru8RtrsEYCGUzr97hdJdH0JwfgXu
CULa3XFHMS9vO2S5QCASPDPWAF1BEmZ3bt9lIvg3YcdduFEfM0dDeGRxAr8mtzW4
AgcCHI21hOMa8Zgj30699LVfPySw/u9x0tlY2WzVlS1fj8kRA4ME0B9+nLbLjSHH
+gs0fsqMTpc9XY1Zbfb8VfsgTT2EpEAZ2kAJXTgd3dWzndCkZv6ZBnSPoJZkWVZX
7hWrJOmJq+qfQnQxOQdnvuIgyKXUPNG5p0W4LAG4x6GIx6dxmzZE64sIvlUm8cRq
qqycIFgTx81dxcsFTfoQ6U1JuwB2Uc/5C46jESk6VvFYrg1UQQqEBcVClk5dcGiB
66SDjNN25mARlmL9ni7XJKMgGnRU9WT+PfnaHvmYVhXA0vPDjdL9LA2j5nOSN0hm
miCcoREP7wTIG98LX+z1R58URW7eA3iHBFD+muqsvUYsuEe0rzsGvKdWnr+Q2NQF
6fpzwXh6eX20MCKnNZgu+3p7gDnR03pZhNvZPHLWgg97nBkkHn/A9zMEkfHduMp9
TkHVKUhyTaGKuNpcCct2WY+6gr1vQYH41v6zclgv4EDfTFh8y7dYPkz2j7QBqa87
is/rq1jnz2xnpmV4Fc4Ca7XhSoiXvW473UW8HZZqa0KQo7SMZ8pcebWmBokT4rbp
Ww5ptILuSRvzCsWK0DROWsz8Vn2UXgr8uG4xB6IrfMG8PzWvHuF2tTOYgaVfzYkE
s/vgS4aHvhupzReVUut4efoN8EW5j682yDGBVUVK70LtadTBowDODK7PERTsmIQa
UWCk+V+ZsMFAraQ5TUa/D5qN6zQl37Kg/YHxfgdHMd/h9y+spKGAZjAdffoqYfon
8qvvmmSFKJzkWYqa5i0FALycB3Yz8znk8E3NcdAZk7I08SdptCS+FOZMDVzBuwre
O8I2VxwP531Dtn9xEOaALTEH9LvyPrglP5qhZ1E86ojcxVR80itVJxHakcIpxYXZ
ww7gCTJaSWBPv7X718aclBHcxTzWWfuWD2zp9YV6NnLtbp1DC8Dwby5zoN0cvcIx
sTESdmsR+Yxas/GbaxPHCp0nWDm/sGYe4nhZhY/Nt+bEu5cLMQDFLAFpudyzBAF7
CvzflAiNU9RTOyg8saPAKBq9rwqWrQ0fS1aU7Ls/1mPyWBRdCYGtU94xzivrlOfH
ez0AvJ88M/XTFlkAcJtk0HhncOrU00bRmPbcXk6jqtSGWkRWso7tJZcIqRRK9Qs/
ig0DkMHpcVPSTthJguiSnJeWU7fRn4E2eZ5PMBWyKEa7+11s0KV6m4kSEyz3BYgL
tShsaApZw7CQKXNrYzVS/1ERVbuGUq7xPF/AkX43sURcTULwI96xn643h0PiX9Dg
004BLESdQcec98nXCTpHSEOtf07iD17Xkl0hYILsA09h8nHSq+U0T2wIV9xSFJ1T
p1NUqB57UXAbUT46AGVH3PVwuAlCldIr14Mh+s239ec+pgM8Jg5xG+OQXpLTI5y/
F1t7tuhKSULkgyRfjrJeuhEAi13cf23CgbWBycz7iyub8/asAY5t1uvOVU9dIZhx
s/ZR2+np0nzVXRDowVUagXmDie/JS3ujhAmEBdzfLnao8STzLz/SuvrNinDzC6eK
g51SyFZ78nBu6FNg9jNbkfV6brtZlw0+50vRSIAnCq170NaWqAlNjnG+3XyemNPW
rquKmU7zCSHSs4ROaWLLiGDpNvtBpSU2sVXecQMjT41Q+oIUjCwS+IdPoD7XSNQX
4xRrNqzMXz1NZk+0DN8BV064HGw3ACcbgpfHs/t40bviY44GNmHzjcQrevhzYCDR
UC53hSYx5792yaos9E0LFi5mSMiegBnJg/vThnOIKCnCxmm239Mai1Q29rslY9uO
PC0qiTldf8hueOWKAInaEYusBHC+pQx1EOf95WRCIptdyRdC35+2uskoohuXvvdn
xEqSUxpSDmhL39F4kvvzu0qld9vFQn81HQLztLR4Gt1/dCiuxM8fSP8d1w9lwRO6
3QhZiWFycCLPqTWe/fxIwBqkHTJC7c3h+thfh4aljZJU0KWYq4S9SjvYIzn+Q9mZ
Ry6j+q9H09ngvH6GiZXdIZ6QJshLsWTMh6rYuiLWAppUjUDsQu5SKb9CvPWzFIdY
tL1UBxMX+ipkY8YiDzc7hxmVIrBMo4MViFchOoSjeyTtzJS6nitWUcj6ff/GFQap
UdpoJS6I9dcFUNrCMK8ZvUkLVS6o0HMdQvJH1bbTTfNxzE96STutfliJMFIhE9Mt
JRGwT0YODhv9ntW3+0VwDrSK1MJ31A+4zR3Tqa1DGrq/TZtSaKnr8isO0zCxy9As
ng4im2wT57Lii/VQ3PtBr1mmzOhB3a2s8aKTUPBrV3KrWvzY68DpBx11dmVoMaVO
SKmhuFNBlJbsLSp/fZQ6kZcB9JkOh+WIzPdWXxXG5+4Kcg2NMgpzyCaXVhTxyMbK
gagd/fbkhjT5paLyytqNen2BgB97dOi3OfkuaDPrlc8aliEtVw469ZyX66uImtpd
dDRkDjYq8cGc/dAP/zGYq7vJTyGNQ/TPdz7UILUXp7jIXEOiklVcq+KWhOk0iDTB
K77FmPXXd54mp5bTa1Pcs1XFJha72iwET45zIN7ClOFAXTKpoXdRkNcGeYZzkRgF
94uKbOHrbHdnj/SfZPfCAFiujSWacuf0PSPWgbyzCZxPgISzRIn7LJdqL3zzeLnV
NKw6/IDxZ3DydzJ9lVaH1idzcyRJjINYgpQ6u2Dc411w84BL40juyWGAnZyaxXMI
Dzwma+7s5VMenY3DnQjxKzEuOwxxrnq4JvCVCtkc+xYWyqhTKYaYWc1Q3iHksMTx
W4Z6ol2XZGZkzAXdO/j4edEYvDYaGSeX/Wf+CEwcxEJc90JQ3jyO8jrJUyrhf/r7
PinD9zkldygBteRriBpZoeCG367GT5SlFCodk46XtH6o+94vzWWckpan0nlQaKL1
CG7LuVNLhZ0I3c/zF2+9qTJBiLqdplpMA6lt6eaQlK0rzMxWpjBbBokct95Dro/C
8X0Lq15SIBDQiZcCsK5Ut89k1S6dMMVfKWySJ1tBX0ubEaZmCynbZ66GMkPtSfJL
6yLGa4UWGsPYIfaNMcygAW/znR9zKL4siAwzq9PPWd3Ldl10p8KKYp/TUSJYCWFT
lF+8J/iyV8W7zF25Nsgp+FhtBwoEpSbZOwo3hwxSmXxZcOkWtX+x/l4YFP9bfYoP
QPa5WdCK61ZVc6yKPCpHUxzlSo9qWfhV4aMnrcRDBJyEyRkiTBQYHxlxAGcTIeJa
LDOJDPB2YUQ77aWbwtGWqLAyVjxcJAc4Kv/r82wqjSCJVtCnT+epAw8GPOuR5wyY
O1Kpw8PMUqDxBgUpb2X7THRgQhQe6q+gksDSpXif8M3U/48FnYgH7El9SPDFlJdg
S6zl/wzG+jz81nxac8jwjpXq6+xn+WdxybiVrdbWKsA0yhhAmPKMLTwWKTgR4XaI
ysGPJ2JQw3w+QmDLpq8OWYRDkAiWSWfchIcSWm03S65Nj4idycdLlZ2uQ8lDusVi
wDmPKe3KZmmugC9z5OF2ujYHbUvXWiWCnEdDbnetf4OW+4j1fNuJIqIBWiffG6MN
kgdynNujUChDP+L7RGWLygPw62/SPNhhMowIxJ2lHmLMk98HpQkrZcTlehBc8n+i
9kqYtRirsIAsQSFdb4BeXUZdl/Tly4Ue/ok+xxzxsUInwi4AwjQsXbY93p8Daqn5
1WVT5oRVTooVbiu4K9JumTPnod5dblvtDT4e8g9WA9WHjtpF//81pHkKwXAMwFhi
vvDmMaLYtbTSSWUpEM2gl24tdthc0vBHo/efLzTGJkOB5ow6sdOxUdoGCf1+1BgC
n+NN3a6R2ceUXvDktM/vCLLhZqLGLkqOX3JxSP4df8ksIz1i7qSxPeiO/VjfPM+b
Vgrs0Zi1/q9iFljNfJGan20lXPRokK7ojr3ha7DPqtEwtE0AOP20IxFcUtNoncNk
ChV1DG2MhuYro+FDfKUsUlV4LFavPGIZdoVF/IdTWx/3b1kknzGA1pedYq/ckJSJ
AUhnWqTEUemPlxLRrOs09vHyJ7KHtYi2ZWTkIh3Lg5BWWnf5y9uiUOu8ZWcTnswy
lgD4QQsnNhX5nO8FPNi4qxZfX/YtPva1LBRmKKnKZA+Dq/OZC9YeyahjIN7mvFyB
ocpkxdcd5Y6hWIZ9MI9+Q7bpZqETvrF7BBGAsNWCTS063IURxc9TaBZ1SXgfH0Wd
Vi8WPVsYDoY+yh8S1lwW6+V840NQJFWbkSPGFBXcwUVgzLyQFqlmd/Bkk/EibHGf
BaQR4WQIJBIso8tMWxwKcHyqUDh4yNe0upNZ2VJjh2byj7ngETmumouxgS+x1Uwq
XTT5fmrdUtjRy5g4fbb6dd131mIQr0CDlKyDFn1XCurrB4e8RC/fMr3vIG4pJWRE
O3QpLdw6ftGXQ+Ar41k8kYndB8fBWpvHMHVRUBWv2uf/idMIOmzBMgCputnqx/Qc
WwORDqeIdFej5pgq3Ju2q36S/o679d3KJt8jyFPxkcSF7uMbTWFbw97vWLD3oXAQ
Jif7I5DDtEeEqtoE/Mv7tXvbB9RATMGaShxc/h0k2lrJaDmq/k5a4BYlE/2cwbMR
gkXTDJYaqMjeLQLmVSCI2K6/TWwuhawS/3tp+KvFy70NvbkNL1H7E9sbHibb6O5e
tG4QjdIvGWCmBRrAo1K1LpFED+aajWf999cdOEPKVXPo7dcxLbt6Tuy6iKZfby9p
uLuWRdJ60Z/iInyPm6thKiHeO0tJk4NrhW83IdV1gMV4IZxhCpqRGk7g9qkCYXgW
IN6d+pxbNWx+3fXAJJBLf+qJoYAkGxWb3g+MpmD5THsgEW97O16e+CZCxKgH+PC7
9de52UKXb9NKEEObtVTvsOopHjcZBIl+KixPWGpbDZhYCJTb1Eev2ez0RkEc1K1C
JV9+NFVv4wfTOkW3f6nqItMBE3evYyQ2QuD/5YalaAbw+TAFpkSafC+WbnF5O2wG
XzQK1xVLaYr7/FcbckIQ36+oYCBoMRnUyYqpW15Zp8AYI1TUMRX+IQoPkrODK0/4
gc8ekGLKb4hUfUI+633zGpOjH2AoJGzjwQn7uoO/ELFAkMGHB5wSUat6KxyZQJOw
PdqQDcQ+ZEeTzhO0jjmfwscQYvpJtW59Mki0xL+FC8tkwr35yJk1KMUssv0RQAmI
xgJNOk6SodP1Zgf2xqCoH5yG4ZNKZ+CnEOsrNkqwoZA3btgGFo/QBI2l7KYiV32E
ifLqcaM966VcbzJ9kJ5UkW/fMkrgi8VB7XWiD7E1O3Wqqqf+a9ZkJIHvSKY6fEHm
MTcTjVJt0ldxfnOiz+wa75F3S5nyd8QN/Woyo4H0Ngmws58iyVe7IhFOVw4Jzuw5
DF6bmfi8rva2a+WEYFueLNiM3LWHtBsBCNL1DZYQbNFN1/oJVJpSFcj8GjD41Teo
WqrbiCEgXUpghEHALtkpgE1oM3H6raKu32sko387tSR5vFkr22tZ4ZA9xcVtI0uj
rv1V6gGe4zo6qlAe2Z0fOOEi/EaNUPcWXLcQ4G3GO7clA7hSE25yCDybL256okDy
QwFOrTQMiT4ClWcHjTTfVF21f3wvpsFE/N5xTHgfFDjyEyVpLWEt6Ullb5xWXXCN
4IV+BtF55F8/NIjW4bkN5AcpXo8W8Mxxdk0HZRn4QqYfobQbr9prBYv17ORd33yU
KFezPvYwI+FLjY5Xx602SXD9eFLUvvHg7V/1LCk9XkNXSKMLFoUO90EKQ9J0P+vS
puZ+pleTfJ1i4q1mAjrJEgt8883lZPbZ6MQJPkX5j9W/jMSY186zCZQxesJlNWeQ
Il+Utau2KLLd6GrMQYV5Yn/UN3aQAveSOs7HTidiH8Lxhke+LZOcjI1Wl7Qm1ezz
eqlpiTd+/QxeSu0T9Vd28Ze7q+Gsbv4v6ONDIeNRC0TSDTKnJmkpwLCNFYRUoW5y
5eYauk9LV3PHm4a9vmBnyeaVsakJqXVHTBgZlpUUXdYC7B2g4ZNn+3yy12jnrz0K
VoIteYaI8bCTAdGODCtQYcSJLFHlQNbYA3JuWOeu3kNIEFD5bgcUZJnYIzT3i9c+
BZ0MFUtw5ZnyThJcKPju6rpgSgpW9Lp4Ze/BOIhiaWNfwoidUkN4bHUM/slUC3ws
2eBePS/oInWgwytalhSBwt1TOLKN4j9AQ/Ix90byFg8nw3CbTWXKrreQaYfcl3LQ
RCQNp58Q9dzvgkNJ6VxoHUi9D2TKRDMrNXYf3DEKz80IvuAmNbRtkjxaExXI4u6C
bZFo7Z3wblhjJMgSAhMZVZpv/Wgsuobxc5W3/hD8e2q13GC7Np10/xz5TyLV0Mwd
NsMcb4zuViO2vClg1nhvLeBnacjhohjQPwFrZPF2LL6D27Mg2ZotWAABA3UA9qkm
ZVx/+MXNqMZ6cQgE2t15DrREdxXywieVrgRFJ9dmFf7yPuRH6hULgpa+JzfRBm3b
wx6cAn7xSrdm35v7Yf+KYJ3CPDg89sUNa+GE5/rsWRtT/R1kSqPbcirFq8LuZX57
XBm6q0E/NKpRvWZ1S26u/TwX/0CRAW6BSIqwf/8Vrh/Z48sXn2H0maEQe1hmW5P3
QjQhrPOfNwKicQB4nY14Ok/hNNFky/lHNVcCshPY1CfN6gW0qE4p7XXvXMXnrkgq
kHUePsX/lriokzmuhPDxA7+mL/I1ASwzBnMaPDB66gSB+y+XYyenmC5lKj7UXJY/
zW8i+8gfVvEKJlkgvpmIEnqA6up/lgiOpj9+t4HCoEHYtYCN6KZr4vIjTumEzpcH
p5Sulg62s+P5bQEYcvCu+W1JVbKEWJHIYolNRTXjtoaCla8RHCqVlZfam+2VVH4R
OE3H2weTvWXBelXcmgRFt6X2uZ7JXNM6P54gooDh5BQKFWt8KihoS+LHXJmPangq
5uDDnm/eD20YktpeJl8kl7gZHOoFw1g0ils8EaFlj4PJZJk2BONNbNSNiASzMIld
R1A4FScgr8KrJuWTmL5KQUqa0Os+VU7+iMsbcNVQojs2NzNa6WWcAZ61iPSvirVe
M6f6bwOMIEG/MDz62N15pU5lEwaZPEvjij59DTfZMAk7ipD/ygmoqQYePpAuNG4k
C5ztbOkGnZm4F6Lzan6djxACveXilEwb4xtjlcgR+cEjomztOOZdu/t2wtWpD+rm
GpAmO8bJiHWI43KyN5rzwUa2XsIewXseqG9gptNxzpElYhnDAL6yDa9tjXpaAeaJ
A+95e229u35ETVYaw4VZ0t8khgq62wy1dZKjYGbGSz6NkDgCFDUZb67ZAoJLh7oe
nVVpaoTOAS7wSh0e9rTgueII+6PR7xHqYmnpYvejh+GJpj/EJzB0q6/yzSCcVHU4
Nbuwv6M8Pok5NpOjauILjvcjJkAEqAmOiOsSqTgjB9E7KElJJ1F/h1Q1FbNhHjda
g+BHy6jUVftkAN7hq73Lh2mvMKCE0z7FYpXvr8kq3VeEA+sQxGeNW0Bt0GY6A+Kr
CMsgHo9LUom5MtwTYtaTH2u36ahI3yG/eptP66qHMbhYHInvk0qsfiOGQe+u/8EQ
rbYLCuoWjov3Jv/FxSg4EloTRZCuPbX84fwp/7oOvK1wq6oRGbNw1HKsgXSFrNUQ
deJD26qWYy2TzqFsggBCPM/oCmIC1O1q7/4Y3EDCgQCw3N6ffYAXDIkOLxZTVgZJ
MWnkyviY8mtoDteM3/9Vl3dL8KwpY/LQ6rZcQ+7Ni/X9hpWCE+76mMSKE5YIPlkL
u05fF0MVNGpcDDsKGaZteXpQrH2c5lpE1kohKQKo7wC4d5K3PrI19xbAkYkmTqay
o/MhSuTE0EDZZGaJ/rvRqQfb3hk/M3zCaG/k24P3Agr1BbZXXWKvJN8cCNQEcVaV
dWGkFNJXt/gnvqkmaLXG4RhrElWiPHXoJpCIjWmFvN9Ey4i8gCbE4r/jqLQNxw6W
9VNtJF70s3CuVRow48fBlNSrPK5loZQ/wQaSVTG9j+TU4oIRBOKpGOomFci0rw2/
vPboSlds8rudXZkgs3OQf3A9OXsyZ9XdqZWxEdJ1JfibG7Xxi/KC1ow1kP22mquN
YhOBOMa5GU2pOeLasBt72vxc7oOHaKSOxgaKcJnpKTmMN8ktiYfo+HViFad/j0Ch
yVwj2Nsf+5M0kIr7/Cp4vrcHXzoj3Qd9guQqyrZv9H4JSS/xXDORzH60w0LYp8ps
Xvcq28Qdk+1ucJAoCOo5UjbzGc0/pCsI0JdbRqrDgfuVXxUjQobWnnxyWxVy5CtN
KZzeyIrNy7fCW6RWdDzI/tp7QQ/0anZIug4hyrShhPxOE6Q2DQmIQjXVLcuCUH+Y
lSYV2waxFlslUb1WU9tuoL4ODbGQPIVhu9il5jdb8b090RAEQL6rEETQN1zcZ5Xf
nJ7R5MTaoH6W1pKsEfyMG/qekwR+fPOdJnjvWxl82eIbLrGXpW8gB+5sQjwuaUtf
vDF4+Zl8jgv9OOtXhjNKn8sH5hLUqa/ayHDi97Tv510eAprn2/RdnW9m7lwlqDPl
/I4RBJAdd54tDCcSbWI9g7iuIVIR3N3jS+yV/raO3Pb98AdChbI6dk1/BHeBNHRO
o4S1GismwBcWUWMgDkeDo1gqVm2SW5kXrdgThwS5afzrlkM56Fmep0rxnmFfCh6t
V6wypPaKRTcWzYUN1Qo1IWesDOIBF4AK7HHazhjJ0wUBEbjapwHt+lvqYMfVhn0P
N25Rxdys71DnhUdX4NVcNt2xkRiwrPSVnbZ3XRL8ffY3DzKwbxK+PTKEoRumtaRk
9uT+uLXDui6DEI66/Py4kL5py+FYhlOS59rsYirwRBlEh7WvvzPlp8KYLjo5BGSF
7pv5ivXMeWjMbVtwJ4IrAqtKawyHtVQSWUrVnrXBxlJ2dqEOPq7G5TKTeDX/vx6i
KC94scOk4Kth+0GHlcVSSZORZETo0ciI6P9Ttz7jRVmTOI58yCKG3wURMqMmxKZW
BfYpuw14tbA6dsB/UGExIilK/7WK5ET9mDWZVuyZCP48iIyOpS9DfjIgWHGi3cMW
S0WNWgNUWgW6ND2BIpLJLhOVqB4FaYRxY5snoFJNiuxjKJFQ/wD2ior6M5b4hNnr
MN7jWyBSvyqUjEyI3nd2kqQ7e+c6asuzrBs2/5vOwYv/Vm/Plz9EAOkVUzn1yLhx
7Bd3OLLskiXFe55p4jJLyY8CSoA0l1+9k8P0dxGK69caxnlyWATrXm3wcvXnq7RS
gg6ci1ArAV7uzdEH0Izh8RjN+rotdkrTiYfPJ3SnKLJowHRMMHGzB1YTSrSOB/v8
2Kq5qeBzH+QsB5PHLvs2kTo0StUrBFcfHuHu5/g1d0OHPolh5Ed3L8CP3S4oZ85/
99Wxi79zQzu8UEIp+K0RdqSUZuMJDAX2EpkNoGE3WqoSZG0Fh1d5hzeY+luXnjZI
g4W85rH0XZQnG6lPXKow9lc8CjR99wx5FLI98AVIYcm5Qskt6ZWp3590nAwK4U96
CvOBfjNy73hrb8iYm4gc5AtBkC6ebUCh0JKeWqLncKB4xJvi148UotPteZ2Leq7l
ymX3OzJDgxpCTb/X+dG8waTkd4BecHuZ+4849Pg1BWDCzrdgCp23UimuxvJdqzZh
FV3JyA3jY4y2RdpLYRqZZsY4npvK1ToZVa+9o8RaK3zfv7wEaHU0lgQzIESTj4rn
kaSjbx1X0lvpNGCfpQRBbkZvtOU312/uZthnm1aWdfJko1pDphmQI0pZuYWDvXlL
1IXgaTpPT0dfD5rrCE1ImSWAVmEHJzuVdPUS2ToUAJu/6O4DojX7yK2MculcWjy5
tMgnzJJFpwwR1YKKM8r7BuX5P75KA1NNdKMMLfQbEjR/ZxRT4mIiHvWOniGj6n3L
tXJH4GxugNT96LcJeuHwaUXb2ZuOgJ1aABplFVTqN55fWTuW7wY+e5u/dn4nrpbg
OsX4XGaWRk4LtVviXJsrcUiFJre6GOk/y6qgPPe6bKQbKJANdzlLJbrayWuBUhOr
HusqRKoA1flhWIk3jByVR114KNBXSDhv2Z5qF4UJxTnmrH5LQA1P//sRS+QVk1T4
1s14UvLe8xo9if1WjLUKz3QVhJVXG7p0NU69UPy/qOyCUI9hwkMJlzShUD2bbOUj
fDQ+aiFOh/jPyQfSmmrFfJB0jy4baJFoQEv9GZGmRp54/0wXu4HjfDIJo4br4VEg
5o6PZzgSzIqAUw2J3CSswvKx0VD93WmVfTVvzdKCScNpPOV+bW4+HoCBWJL7yoEM
gHYaYvSAfsJWnTwwFiD0rSY0HM3VwU5vUTWm6syZ55IYPT3EBXIVoLS+gZOWUMZn
Ecp2xGbQnwUDJTzhzDoLXXoCayymrTi16siIFERi31WAJLSgik5AzJ4CAgP83uxM
IriEGCS+sRgB+nIGvUWqqX1hmpI6RP3CGbKkvV7KIbXk6dPYAvNT0YZAyczISH7j
HLBCob+rz6VqZZMTHbiSp+vJgFwfis/4/0MIvq3NhiQ1RpUgxisIBq9vTu2ZPeO5
ivV6wf5wwRbL3f3Bk0cq5QrwGFtYl0PSOPs1tNialARWjsWN0Ow1/zDFGar5RwMI
ZKgJHYmxR9puOpnSsZhjl8Md3Zh8k6d1ET1kbiTztodRtA422KSxqUSrnt0WfC7L
Ibzu6pqhQBMENrWyanW2AnUp/rA/hps2TpUMfcAMO5BeDvo7pV9+1UCRkE2MxMfd
qnTnmFAO5iMPRC7rpNCX4MGbXopjAG/bnzu38eu/4YGwEqonTSytzFNZ7zMlZMhA
1gE4cac6EIWlxWBfFQXEKtvqbX6h/fOs8nLBwpaCC+mIzO4JEJu/Z2UG/tI/NG7X
f6Dzeg+VlrH/9UeYVB2/Y4fdhELOTkfkrDllYSvIm9BOp9ERokVA4C9/wK9YYtJC
tHmfM2iRf8wff2F8aPUU12Zj40Y7WSmYhJoi3BAtSp1OGFR1YqK5+Kpzo5o8MnCV
eRmpPFrYFzjTnfX1JZkTN1B/TjY5CF7HhkRKYWDZwOuLu1vyvMlB8/kK1z/C2q0T
lgSb8H44Awu+aQB5OaqqDYP3lNOL3GXvGIvtGaxIepN1vZa16lNeGcfVKcZEkS7P
4AZLfbXHgKohORLDoRJPL+rbk5ldiysOJGsyAHpGnt8fJDvRZ7OYgk5b6WyivOCj
UrEcQRTqPMVMn7WgmeBj27H3RKy0vkri0UiCjiiGOt4aGCD2qDH0K0oRSTfkn4sL
5Wp6yYlU/kO7HnpqSWeWKhBudKVlbhuH6eMHKJSNSojnPZ6KsoGHUi/RzFGMD1WR
PcvGEvKuDIGBJ9+qHWMCEBYD5UnkbiFevY2XrutPDJWYpLCzgs185U3m4yRHZAQv
QLVmx+ERQnz3JW3QLm5BJqdkQvF91XrLvPqYp0G6RCQTTrUS6l8s/8KhVmK60D5v
2ZbIETO+ZI7iu/jkig8Y4xRB6yIYZTevLV4w6WyfHh7M20apn/PUvFqA1a3PUiYZ
8Z/12C0/05cmNoMteKyjxEDcIskB0R+v+bOQNNs2tdnRhAQXVNDExHMsdMwpgcOl
v0AwRJHoNQVcSRNUI9HPe89CCKE80Ij0ZGMT488vGd+1zSFR++XJOUgv1Ee5ac48
ATwq7Tmkg4wHXOPALxXJHLRDxjDJdpXwnLF2zNVaeudtbkYQxsbWslJ987KtSo+q
geyvvGV6DFTdbAfjhNKpdEOLLnNYkF7JiD9wZiaP9Pzpxjnl/imA9P3T04tZaaYe
SsCUdoAEqDbSeEGFRtGRXTaghLfRudy3VnD3GIr3yrAlaPMawfUtNmZ3uvmgRUjI
BM8RlajcI6KUi/2VFaedp0xxc4eKtH0a2IUbNa/CAwvA9kW3mXE7KWK+cPAbupbO
sscVs8jXVvz0xjPb06MsoDihHirg8J2M82VoyufmI/2OmqVtDVcp/S+xLaWC+GQi
Vja7Bkd5Z8Mlwx8hhcDiRDMPJqY/pJ2JUkOo3PrRtwBRWMx6h8KPpqNOu980FQJ1
xV4HN30IN1A1HryB0Enwsad90jASoRL3i517r5aw8IDtO9yV3g+FyJJiypt+UODf
mdE9mub4o4f4Zr3dDdBF3XkyYarY1yqfmSSAsM1HCJjfcWW5faVJBcHIzZaams7p
ZaUXy/9OPcTWGtpvc7lCdmtHC0OjGIH2aghc0bTMnIJVE9cQnEERvQVG3ofsayBN
es+5f3GcBIzfUZegTr49qqBWfdvjxWehE2tUod2kr18qSeY1UOHUnrQ+ScR7G4fR
TXN7UWmliL12xtcfRQmgzt9ToRw+/g8yUQaKC/g88RIbTg+fG8dBowxFc57A71To
3Dpn0DiQ5J6rS9iMVpcnK/LhvWiNsXQlM6832X3+AUynVTTX0/OBcMtsFCup27aR
Y9gGk5haHm45crWz9+xqeN/kNAXFLblVRHvu4AtS9pKAVmVMSeuVRNUafJwPrOrP
FZsH/42cTXqYG/pzGe4RYNAfMf+it63A9w3V2w1+PXzynbTlnqtV8JTSGa31+34z
GKVqFms4fD4CO3t8nQuKk9DnVN3dpbKE9iIzho9toFyaQHvPlBpi0kXpZ5gYq45t
QAog4eoAevs+OC8OU41i/RQmNSEhEwxNaWC3IdzxtjZ795hc+3xWUbW+AtNJ2+qy
V03m0HGeB4vRbXpPUUzd7r/IrqyP3kfD0WUO2yc7uZrhsfKm/crYjO/IS7tj9CZd
Dore/XFAwCvaYCQSpUt2yBr1kYrgmWrNbtKO0ky/6T2K3admxQeFdSP3hMjM+LtP
v5iGIbP3qbkwkc0sbHAj6LAmM1AwwTG5ujdVLrMc6LzaaQENuotXnE0+qL2Lc4S7
QRZezpVojYGwyrxgPk1u8KJuxQdfbv0RqEgK+xCN71odEYaO2Q3ESd8iBhRUrmcW
1hiL1Zzo3mFLg7fOW1g+3jITJ//eB3gEgWNzcVnFNJrLS6vGGTyC2fmdfvUeW01n
HGWure6aQg4c2Tj5HnRmqbP8t5f01/XI56SGz1mn22ml7NoZ8FuCPuYuDqVk5Cb3
Xc3sUC9R/6+X8SHFfvPnu/R3VFGke7UY8EylqD23umSN41Rj38J5WPFTDtZIgmh3
5zucU9CCQF6ua/0mpjYHO+dTpP6CPisS5VpdzwM7VDzXdzBnqbsNOnxvzgOhno2b
G6Avz26kwvgn4FQHSlgk2Z2XXzmNEGDTp4kNrLpqd5LlpIzEIvbPgkIMTCEcg6l5
0Rh3KGm7HsExtMR66uFp29aQtFuu7cqzSIgcxAHxuWHr8v6KwF6YGKvEu6Cl99LD
K3eloWAZiNGEjF5I9eO0+9urjS1IjpuQ5esThFQ3WBqiW8g/kIEx1DXW5gR5JGmm
VAc+USJDlgSMbwKnYevaWJpx9i1KaPii1dckdDgpHAeuLbtuUd39zlUpiqLbirp7
+ucCj7OThkzlJCUz5azSnRvqLQdGmfBN/u64Ho1X/Ct7Mo904BtViq32x1rNWZK/
Zhclq+svCBa3ON6ZUvwkMABhKcrIUeJb2LYn5kw2w/gVlk22llAswSpEE7OWB7g4
LCitE2GuM41J8DySuZ5eMLabj+g1a9H4UAOS8Hh2EA0/RQmdD8S+3kYVbC0avx4q
M/Gbep3dcn4BXT6/J3q4tET5p4wV/3sSldj2fSrQskIHGGK2HafSff6dUWzgpCbe
itXPtWr4TKrJI+YGWpV8keFexxIKwiNe4e4MkBYYdHdgTwFVIhDXFBeKhxseKWtB
AQ6kt+Ndru33CVAa5ySSEwnogSq/z56fqfV4vLGDQURxmyKWUN69W2OrUnCVGnwS
XAqvaM6+2+GlJ8hD/gOKJE+cxnXc0HiPP0Q8QuhQTKr6PwMnyAVVSP0VN3fAQr91
RVVVKPOyUf6uOonMOVbaz05nctOfZGmkladcI491g/RrYYlGFGN9oBZVk/5nfe1Y
M+fNL20fUIpE4Vuc/Pp5399nE1MUj/iAhTWuOs0ULvYzx91WBcGoryBeQMIWCgV5
vHvYdLVgLCq+OOnA3AIHGUbBpVk0UFmKdZPKU/igPiVlc5zrpaHvnA/9WLmnG2+j
8Ek0fE3Cy743w6Rdtr4HU7KQ8EDHpv6vRseVUt6NElaWofkCuIPkZSseaIjbVcvC
cRBIDZltC2pOcGEIJDMtH4zN2KIqyiCJ+2bAVIVGGS7A5yAHzEwTqza/xQM60JXR
A7BDzVqNGj9TmjtxovyFqGYwKT2wB16TlYvYdPT0f65L0HC7jIHiLYDMUwbeuc/7
AQHn4deDiGT2D40fBPwE/5L/K9HIjI8HCnY4xgfYhAcdNFRRCtPj+EsBnYCeM6VZ
QoIDkvkUKUwDsOAifwua2MYE+LJnktis5i/6B+UwN3RgMp+Wx7GLmV069WSuFskP
k20GtxxgKry+8Home6kQt/O100sBHrdlIdxmpcrD7WRXFFnFlgw3pychxY5RiB7/
2CUSFf13jVj7OEmUur8rxW2FEHdN9Wfalcg9y4rUkhxOcfgUXvVrzH076Kpwagl4
39hO88pUUm2NOlqH5HOPYllOrfa2elfdkt1d6ir9fJ7+wSZaYxexd70fOSWR4vvl
pWG/IY+PYgDk1q3B8zHKRZMeyQW7CeiQfawSguK291eRWu0jwMu39dF5l8EiU3Mf
7M5gaGkmXV4DcwyUyIu+mMydlCXiOjAPZ3Utz3yEV5DNLgN/4ROkHj4KLdoZunGC
uhElstFBPbFyUeKLTmGaZHznXGYsTZy9QV28aOk1QaJtXbZzELjnePZ4R4EO+b1W
pzjcb6w6RNik3oBwKVWf+eKwowy+kT1bjzqcX6F4AZmZQKkXA50pJpmovRQz4xVk
MnQF3I61Wv8trfjSjCtHtSMdPfmJS57C/6JZ53eKdN9rQUpNNjw58pt55wFRasjC
w+CshM8B5GBMJ7zgtG2rBA2DF4NXERGN9MHHkrzPu5irzCyEN4WyN0h8CMPD2RTn
hRWmgzkoN4G7r//DRsug2mNhsjAD1PIIDR0sluSkT4UNsDGvm3zoYB7SKs7hiy1c
e/VbkmsScxfYdmz7kDN590skuocVZx3XuTuAjqCLgD9cC5PWx6N0slPzFBrzNpQX
AnPFoXpfhgkWWHlihou997lEtt5PfKJVHFT6MmAex681NXykSBm6b2xm+wbzayNM
MF8rlqfqfkCcLBnJswlv9BUKCEXj89suRb7cl6MwfApUvVZc2kLlpsBWe7fgsU2B
kF8SGLfhaMaNi5oiwal218S77M4OA2i4Hcqwt4zhzS/3JFyewIlUH5b1Im2NP/XE
+HFYlM5Di7x2GGS9Yj+KVH7sPiT/TrmcJX/8ZdmqjrGgZKq5KOCGlj09D5LnGUzh
jpCcFcJnKnjJt5u6bsGoJitxbOMR35LWapPHQlNH4OkvUvouqwp7BYgQwdDmJyT5
R3Hi8BMNXPxKPYZDkEqFnGxK6M4o7XMDMan+SYrwOTsQyAzfdQn4dQ8gTmlJdvOo
USgAJTo4A4mCATf9vkfU/6WDDJkxWAzIcS+TjbBxBj8RMN4UoQgAXui2Ja6g5+3U
CihotCGw1qSu49+g4lTBbvDBdItldxNH7OgmX+Dp65zLicPdg4yA4Ws/KFxhQI4I
a8aGvoWx/z887vNfBNI73Ubirowx2Ner4Inc/HgpEmvqBj7tSd1lBV8pD6ZhDPAo
uZmmFuHea2uRSW/WWsiSaptt/vm4DAgD4MAVZW7GeB2hmLvtfJIKNyKrDMOH7DN5
xobfLa9fJTHiKp/4vgi25Nx+E29Yquo9cAQxWrX7+ep43OUJRlGa/cMuRpqvGh6/
amSa9SOPZHu47/MYFHTpZTRTEfAwewclmBfugGuM26H/LZNdVNn9KSlgEACvKTG6
OOTfF/LEFvHpZxyJ4aQQYmtvT/PXOzeJryacOc6bu71voDV0mseqgAvW374T0aWN
aDzsh/WV6CgSpebxcEWU5EZzamGgxWymtKU5wp6woekhs8t/HLLAKABuw116Nj7q
crEgvv0MgDOtmsZjMAsxsWr8UJOohSijE6BTg2sB8+cD9agQGLN6P6w2tTw4ZQeY
jQzanPEaw/WazHuEjInjhHzZ5UJVM9aBRZ0lB4m4tUXgQuOl4aRkssPs3xS4Qcmc
ID3Y044Nlxk6EPpcgnz2GYSw206CPMTHcjfHFpNsgK+rlVGOV3FZvN+IlHuXBZra
Feo0uQoaeahWpfNfOssp9cQcalmmZUM94lXwur+1XqUZXjQ8UIdj0YhtoepsbfrB
osEcDcaITS7/WhtVloKyB1aD+F6fddLMkIkIjxP28VW5fAsoFB6M3vk6ryCfWRP9
vG2FU+EEqQsJ6dkFJBeP0xALFy2o5EnsSkLMj3Cr8r53EOQS2sr23JsJL0vKBBcC
q26TSliXvwtz8iMWS+3BvbZQOVCBR04UtjQ/BZM7vk6nIXll4YX9EBRqbgCtbluA
PAqoUs7fQWbSL85bPyBIKFpzyimftlweeW7k5Kb76M0X+HBLfYQsH4cQ0b7LPiCh
JkwjnP6r5MW7aOni8trcTQNLP51+/pgngUbyYmS8I6goVHjKurXPQSnxdQm4i6eD
UaJkkbyoqvAOz1iWosESDROMlDW9LsNAPYE10Mr8Nmdr9+AGzKnW+OVvHc0Xrbgn
jCPdTUyAm0ARPMbcVQgpbcA08WEnP/BLkHvT81gqvDy4vFUIuOB9sIdI7fpujUqU
YZiJ1BGO4AfMNX/hYgjJ/eOt5rwnbpWK8iX0o1CnavercXpDJoNA3elSy3dDvAZa
UOH9TrEG9fqIMHeDGDL0cXG3xaXKtYQt4gSRmH245Xx7i4ycH7LIPCNoDDgKWEhH
C37wp1GI7S2u632rBLJvSEIhc25zlFU6PXRbVp1TD6WjRrrxq/W21jTimrxvjVtf
eCw4nwKi9/wElBNstYu4Euzg/qc/c/F0L+TOsHboOkCNoQeRqQc4YGqZP+AC65s0
8NEJbicxwrlPVTzY3+Ifak96bFe4ACPD77/uqixts+NY8Q3fJpcHephU6FfKN+5E
tOcBb658ilLeUSPe71SVhSKPK2BRRyzHUKFJSNVQmC53NBeRS72ACev5nMRixtvX
Pq0grQEYdtZ4f4obDzxndUyU02IJ49XG3gL31CFZewFV4y82CkmYdk6LM8dbDE9e
bKUOnqeWyE/1O2335WlNo+XTkAfQ47SBnTrRFAPlj4hhPMSIH4/KxIPT1A5fpHM9
FL23BXswv8Sx8Z1KxOTEm9nJAOwOvJYG9GbGdNuNKr0lqHhKNI+AGjQyznjLejGO
0uH+0H2a6uAT7l9ISazEdLs4IpctyvGMEblS/nhUSytFDu7+qFgoqfYY7UNG1pbC
j/BnG+4QDo5cWzPzNJunYL6K6nrbSOnqZuBogbwEtO83HPFWPHAcPxSbrrE/QzJg
dt6ZNB+XRWF94LvLRAJ7UxC0IT65/1NcDV5cKp8Ic2kDbrcB/BK8HRGKUxi3abXm
UFrvO3qjxjbuM/XlshApXF5lPmjj69+iQEhBzYUhXvkvsQY1PkrjwVdpjS0HN4Cm
lZzHC/Q/eyyYcY/F7unOHzjjgYz9RJL0KyObikEl5iNLfWkSkxLwjGlpqKL6dmiy
byQL0/amBsaOuC1x00VVmcsz0iTIUrcasx93EtWkAB0eg0yNdaSrkQwZjoPG1Fej
K+RPOH7GN+IFzGhhSn5MzCzWZf2bYnr96JAg5p/OfIc6OFlSp/h3U8gpMY3wEt6B
RxZEqbgYxsxGV2AV1qz0RW5nIBg7Hj3+mQMldOKKt9nSsP+sFzaMCMbqg4MaQyT+
Q8ylFr8BjNh/MOx445Nv+urZERn9pA7uxp5zjHTSK0ABFxw/2MKztJ9p0BiCs6pb
oEr0TGYw+qlK3p6vpuah/NYsik5ls5loT85IrM2SFRl2EuPfauWmzrsHItscHL6i
qFqBp8vl5oI0Ct/lW3bQrW3/vN8ncPs/u6cAyePP8AJ0q6RWdBqEoETVLiGcqGzq
m0CsDqlZryCb+rr9UfCnRBZ//XVkg1AmYVhiBiLL5uQ4WHTMxy4Mlkv7PSmiWEXu
HOAPgb8U4n7uAjFKkX/TLRZD2OIah9WFcGwcU2y0MZTkZTuUEukAFZ1zDJ5NDeKR
mJyNCEfm2G5UUDSG2CBSZba32ExGMcXOkTf99J3TiD92FCpwpTF/hs5xZQD4es63
WT+LbOq7bzaDaOQSe3yk/lRknv/i3H4OtKZsRfckhzw+FVgNm5XDkfeIU9nvaZ+l
/qoor+SRP0zQYSAPpCf90YH75omJLxPVLCDAbw+JfmRS8MSAWg7Y5sulyfSoCKH1
V962/ksyzoCq5MRa6Gj7O60XeiN2GK6IJXoSfCIg/YsCUrvZJufgZFonSgdBuvrs
mPo3FNn12OV3FDja2ktckWDwYC5pCVVWB6VA0tD0M45YwLDVnFMbBGnNFz/p7Fp6
G5UBUSYBwJ4LgvKMiIXd8SZYjM23COCES0W2oNHzgs9SmhuH2jTH7OSwzjfGSpeN
lFfHFgy/kzjbZVe4Gkf88/nOvQAv8OsqSmc8TY4PD2IcibxanmICiVfJziArY4DL
SRm72DolAK/1WC3HjNui6zp7r9nWq7+ec426WO674cOnrd9zfBhb5D0hfKMc9tpP
PlSilvjbi4Usqwz6tucaktVcqL5zaiIX7Skew15cILop1BbAklDd2lKrR9K2YcBT
Ej2Lmd/3qR6QVRPOaIaUeP6jaoG1zOkSds7mp/Q3N35HbcoR026gu0fjwuSubgyl
eX9JqnSJTjLOhnYJcS9hVhk90Qs60nuU8EwQIETrSSs8nncfhsivBKk0D3buwzGA
eMfxRSfS8KleOtYKkzp4Vtzagbp3Av/9kLDYH9Ph7dJV1+zcF5yAFtb0qW3A8T9U
8nyR6jGqyi3XjHNr9UvFVrOPaXIkr5/Xr6Z5ai8PW7Y2Z2qA39Zkem/b8IJvTpBk
KQxSzbO8DigW92KsdbLjvOJmImwTvTnejzWUk7goVBbSN6BLp1DygRZN0qchSAkv
qeOW4jXSeZqCeFLvsEIZBsV0bXNLJOE8at5kH9T2u8yz/nANzGEI0OtdlSCd7L8N
1D8xav7zWaUq/TIr7VLvEtudSEt4XTWlPm4qkeNQC/mB0RVCfGqCeAL7M6M4+l8r
ab87FM5rHgAJJE6nJwELIqzNvhxFohTzXa/Qk69cE1kKtTMPI2pWz6jz4gXpwGZ3
Ki+8oHWaUu9REbIDpFlU27LaRuGEVlDyZbO9gYtBqvyOhBSJx9THp/IOR+Vz3LEi
FaX2rmmunRLRz7Jf4YDP7TkSqTD9+j2+0t6EY+zMUG/P7R6pORtBhCsIzmOs6eDa
LlllRgDyWLvLXVfRgooJ0Tk0qK3v3BoOXF6iSPM5ytA/I3UE0Nw5riy+oISTPDOr
Eu0kMYGWYTgKgjFLpvVkUt/TR1U1tG9EKDLcWaVmhtLOEgr4PGZ3eM8Xr6ZKcXGu
Ug99g5WEU80BlhaDJOdwPBc5DTolROPuJ0fZ711jZGCEx1n0gonn8HWADiaAttr+
cdFtqMVwOXd54oFauxgDZvKiMGiVY3D76Y1MAp5S2y8EhWt0r4ELoux7b4qbCkas
XGY1QspOuIV81DzCima9iNxpEPJCzchRufdmznUZ82n077EIDXDc2OHFxQ6lV05u
B1fZkHi/cI0iagYAzVpKjSbfNoYagvfB8L9lJ/XVefS/ounp+4H5OO8FBmBfgPxg
nf/CFNuVm52WAoj7GaiNIMHkvYe7w8GWik84mOEVF9zOElwgAyFrKAqwpoOLQnJI
GYQ3HU3jsqbPS35YjI9aWZDbw9aVte2Nxk0AyGWGfMpnhRxNapelGWo3R+a6XVK8
sRO9TnEdjxOmmxdC72em7ej7s/pYlrXn31y3b7Lfxc9hn7/6gX4rT3vIK0bi/B8X
iEoeh69QMT5fuasRfa+KdDuYakuq2M21az+o2Av28U63SjNdO2ZBZHxZkv3A+dJ0
Ou/XvfJwD1BzKIZovTp7btPM71ECkbZr5qZm+kCQTFIiwrruEHIDZbnRqreB99cW
vAokKFLD8nP6grpjVM5Xb1sF4vdN0qNQTOrEePkpCzmM5XIhsnN7crdE8s8wbAje
9Xs5S2pE/iP5Z5lFkvZS3c8rFi02atd5XN1m5RzljzWf9JQ6SQGy0dwLW0H7lLk6
aY+8/V3IE67QG1RAqrzuQ1zCUYMxBWjSsMAWisT30ryF+A2RACglHFBZ3YWKdd3Y
fCwCn15dP30PUS9apQUYchGzt4fT+oNuw6HdhSb5m+SxXzyAAHErqMaMEcRII5lP
fsiZjgkoqiOYo2ADtCLCCCsR0Y6Xtu7sjaq5+6LmcZ+ZUlaJXtUtXbIfFhxbI1rk
S4sV00JGmfINUASBfYsQtPzGx0YoypTwOZsOPYG3QjP+LcaFqQgDCnGw4ReJpk7d
ASimdY3a9oHcZDau1pEz5R78x1oFbnow8XUbeW3wiLXCg/8qfNWj53h8mDvrKeaZ
+qU88Gb+IfK4jYpoHBEFYiRVT7NyOnVHz6SLMdh8OOPbyFrkeqfCjFCQN1SWWETh
r9sMDvZP7uopogCVw60X4FFaPF+QVS6g8uWxQjAjEFfqJWRSeAU1m9pVOA5+TshJ
gyn7W7IX5XLwL9Pa+tAlSwW9kRB5nQHtxABa8/Ykz2msswLR/8CIJ1g0PwWObam6
Dl0O9VXPpiOpUPwL7ASdmiI7QWQAUpw1+KaJ59mKBjAvKwxwsjhWn07x5pIyQcFX
DLN1fmf+tC/zh25UImOYmFFhR2lW0hgOdofxgOfZCC+qV9ZIi0EA4J6gcq1YMmNQ
s7NA/LmkosMeGyVKZAFfvp8LIYJcyNO6CDtpIQDsD4TGbSEahejfXcTa/qNJaGzi
EEY7l8GqK+SDG+x+vqmEG1jWgLn4kzeT9hJCT9VePW4JyNDf0tfRvh+njXgFXlsI
8vPNzeMTtA2GD0ksu6GgPE2SWUEc/ecsQyETOxQ52bWFcnGUDCG++o5dmnQS1EeK
x9mpTgHzFmMP9x+9m337oR178gJ0whXHtGKyG357sMdyJ2pt4A//rR1/+y3+fbc0
Bv3zO9mSCaVwCFoYif1iDelEDyt6nET5wjsyDbKwfKUbn64FZ0OzVjtdSv7wxlU8
wK8FgqFcK9lv7z86qQWVB/ZkAzSffeGfkKHmOj6lIZHKhVpmimtv4WkGrNrq/uku
GYnpRYt+57uWL+4IOJU5te3ECBJXp+TcXzHAa6o2kt6r5WeEO8ea51TSn6ACcip+
BHgAdp2gkrmuWkzfmavHqdM7T6MgUzzV37G1cmRimnjE+s8ZtnQfBE894K0/m6zH
9M2b/TSotQ7jNaJuqHIVYN3HfQAA2JtlR/mtgadgWwQw3tRzpk04jLmj+FElu80M
O3uRU8hRzYjy+I2yQj+XF2xUp/bnRTDGLPUdnU3KGEJEANJFzvvkks8KJxH16+vv
X0sxYnEPdIeAUsxeOO7g/R62kBhTZA6MVppuVD1fjZflsrEWIIi+ODsVt7g5I30G
Ds023sLf/wNUMEqJXbDkeV6LwVCJ2c5DlhZBE8iYV1uU+nXEWJybWwtx/tpuMjSr
yqTk3DSrSmTzNXZ4ijuEB6235k+jeAyB84GYqnAn/11o3H9XYhgO8AV7k1IeYNVC
dcOcSi+Lwadgey8n7jKZ5ObHK7q1Nb03ZK/OTxqcsjb/8LrAfS0JMYFEFAcf+1vO
zgZFvfcATdZKnzuxqMkur3zb9R87I6/9+3fgk6FVmO7HalXg6rmjVh3hRbyxRwR0
QMf9w/6+qPIVN2uA49uPn9vzuBf7lbD9orn2THU2COCHkTLxr0Y3FczytE8UQXQV
CqMkZNM+O/3MDnI9XKmFuPseXt8koM7C8/xPHbnzUJp1wx/J29sFnwt/3psYlGtO
IaHPvYP8AUBKvt/vyx06KQg2n5/uap1WKYDiyzlL1S6bu/5FA63KNy88VCtRcgJE
/3RQsJClb23TSAnGV6C3rXHaCJl+oB2xvnWg8hy82Z8CbpYNB4xsLYBNvyVp0LS3
nCugtyBnt5Jjs8f8NyltF3Dhsaj7x25TkZb5tOaI6twCozJFKHMImRj0fugQv26C
gfGeE+7oB7EGfLe0ZY/HozMAMjxt3GzNnjdIxRbJsL1N6Q6AFPcInQSwjRDf66Fa
uXhu0fMgvmwaQ8edCxYq5GZE3OJAWaA2EFt0Q8XgFtl4X5bB+2A14Nr53LDcUzn6
yv6aH4JI3Fa1zw/TSGqrYWqsUrxe1nmxF7g2wRnUU3nS/EcwPHa5JG5YDYa6tWpS
Kw3e+Ui9Be9P86LKrwz/pQ3DTofWm+B/8vVcroBL/lulxbS3fX4SowsHvjtg3Hfp
DjgK/ZNUOY8hPZ9baSeL/8SABd9CsHKwvrDnE+NWP8oiesguRVs04abBRFsEXbY4
BiIJ/A/HWzEIEMP9yX5xCgclOxQkLgooQ+s8tO1ArjtOHxy06Uvu+PTvYNcXs2uc
ujZd1ckUMijrejHIOkRRBzk/OthqgJlIi6+j9SjoW+o8EZwg4zBZxVSBBWwLbxVu
rZVF7JxR3anDT/EwT81ULerAdByGrRvdNRONVkk0zaufYFxun1tJa8mpsaR8cnU/
YsBkHWDqQuCghdn30fBLaEc423csiukorE4wKUaxKHyPklbVa+QAeFW8ZEy+E0fW
Uiaf9TuG1FP+MPcZtY1DUBKwmT4MhUt9Nrp2dKKeworRHyA6LfSMAnwVLrdW3PhJ
cjTI0v1eU5E8jKUZ9NzsIpTSgLZRVPdq/fiHwvm5jod3lhC74AEqN0sJszqxJMar
x+hCpsxDSmual5sQGx21i+fCr/Etz2k1M2G0MAreth/NtEE9FQN8d4mj7TzMUixd
OjJdGJeLjquGXJpEUuCuQAEjqUn/YHazPnWGnU2TQp2W1OWYRqZM4B9bRQW1qNiT
gTrP+poaESVUmVGM5qqx5u5nPxYTkdXMrYBLSgX0dwYuApaufzUOwAqazBkUXQ/x
AM2d6D5uSRMfm21liuvo0YuUXmWxDGeRGjePevaDATJ7nkM6zBf1rlowy4Y46O13
EHi9n1y77UpnEFYPUnHAfVBaKLbY10r87TcZmtyyTn+S/AObSi2lUNzwSU4+60jg
05oy8Zs2ezcxCm0QddH7ys5Tan7R8VBl+BOxdDksmJlw4zKR1tG7ywm5i6SvY0b6
ij5kgcBgZ/grL2HJIY8q+3+BY7K+OWfvuly1TvucIFrda8PGCWOaYpfTRi+5Eqhv
kX3UY+Axev97BJ413lVZLvyWWSS1S+Q6wapRIfWVCxaCJnqzmF30r80Dqs/HzjGT
z01AMlHaMKXQkWvJPPbtFhgzKgVQEOjNgkc5LsFXL2Tih2drLySFmLm/FT4eJhIW
JneR0E6e6bQLVy3OEgE2FhzXfc9OHo2qS0zpeJkDj5P0FdmwQFilKP3wrqvi95PW
8jxi9pkf6r6Qe+SZAdGyGnDbG0VT/ajMgEmcn3qCtWsvDVLhcfyySuL9alOYqqVO
mn3DTuBSfoRAQOhY6jkxJVL446Iegx3ErAHOPdGMTfr39i8RH+LarQT2cr5xvcbE
yKVNfbN0opprAcHFD2Xb7qNTQhBJV65thfVR9c9GlwfPqILdeAHujxjM2gNHKmRD
MeFX5ePS3klOilGzdetuKh5pgPSlRAGt9tSQN8Oljr+wgBYZxHGaOuFCJhfwBe3s
0+PJVa22aLlcM1Wv1qYOl4zM7SFLgiRc7PxJN2c/2Cbx5OuVzsnEs0pDXW/5ZplW
AHlaWQJBKiRBUYOtSC3/QPBPn1BoATw1n5Ftdb2ZANeLu9hYlfDk0wTroF73jBuI
tXgf2IzDg0qhnNVgR166Y6zUCj76ixyE1vH0FzQMp3/WRaX2sBSjTQagYMu8cXQB
74Nng7gNGhXFwzzCTTT06zxKI3yOa9KO6Bp0xhX7eJonWqsTSafanztY4l4zy2ZS
krc3HtKfgfC23vs4OFzwkcCq6o+ozG1onjRnrVY4M7rrthOgwoCbD6XrBtdoFlZI
rYl0oO797bXAUBwEcZLb7Xepg+T7/I5bCMsfBHSYJC7vV/AzO783b8A+ytA6Ddwg
WjBlc8IDs2w310WLZU3PMlkwWfqyIYoajhBPJa19mmK1z2KxjdKHsR3Xq+1YEBfe
KCHNh6qtzMFU4m1DT3EB3ONxLQ2YHw+oEBw9sV9y7K6ukG/aIfou9cK17znG9OOi
eTL1zvbaKE9Gf1oDTlWFAO0uHzET6pDRJbuSxyrCd0ntKgeh0pACo36YJARSZtyE
QKr3Me145LNoUUH0BfJQaQP9wwrCUyib/eAAer6r5Y2nj/hTscZkWWhLseKI2bj/
zRoAgGpZ3em4agRiAURmIuYP2//WVqQSZSDEm26Ml3uMZgBda87LGaOOGnVwQPI3
4yP3Ec3KjE7pt7qn8Qu+bVW5OgOhVHJWKIj7m2z7PqLKbke3kejhgOrdK1F+jO6J
Fia6fYlW1XWzF7vy13RFRW4gd/O1ByQzelwtBvGbldwbEncwFdOyu2h7Jz62RawN
Cb1DX02Yd5HOm9RPL31XH6JSd37sBZFaZrKstt9ElkDZf7azpGD5DMLBlquIVxtQ
AoRube8zNgfOUG3Wl65yuPo6IEGxdEUa/h27EgdWyjgg/i3cbwK9fThOLUZVU6fT
RoLoDdhhoD6H+8w8WyM7px5tJxl1hw3Y6Z/zkGbIkzg91PXRI8DFuiun9mQOtLs2
p/GlrUtxv9tcKLY53eeweoY2ZTV//7lhDvCU2mX8gFTPG67ie+LJOCiD027ivxEk
pvnBA9YZvrLhaA7HQX9uqiIp6BlsU3jLL+mgFPdUL27HhVlKRlb04ANYwIRbsZss
eKiWifg2DXlv2XNp4H7zUgWF/8vAYH5JrBwmlrnfEm2zwAaGlNCvVC4XG6yxNLHd
gyr77J08W7cG1sXEFnC1c5I6/uSohnJgDBobBqDZASWY2YyEmCxppQNHSMfDOy9D
Wn7aB8uE7/BYWbTDFAQKUTXskYwTCc+ipNYYkSJmiSIdTox5qApQgz/owbGozw3U
33l2abDbm15vDyZoebaxxFG30Zut8rbskWHdOn7eugVfMFHO8H/boLVM3eEtkbeQ
XmGHTqaXFYdYL1r7olRhMCEvWei7WK/ogjvnG7tvoVxGQkAvsc82AveU5ysQzXeD
fprWylWTYGmTtV2Kn7KF762hqyIA6W+ESsvodOLMU0Ei3/TurHcCt3vUIY6S5ok+
Cl+hdRZdxH1ELy/DDcMqT4ixtEHKilpg6XY44bnvf0Bw1UCqBEBzqJjTgh7GtLpl
m5DNtxfq9gN37n7KN8I36/+5lIV8igmPwbb5cnsxMWo6WvtN3IHNcubeyMyu6zj1
A3T4lkrNa9FQ8buoMxUEy+27pN7rOo8vKQgWT9uHmXAK+gvMTTwzaHZJEhbt2+xU
t9NgzLeWTHlkt27P4oZy9i6nU6XE1GkGypnSLCiLRukvwYyGNbop5KH2Rzt2XQI4
OaXUc2ZoT1NZ8XjDg5BjD5Y7ry0sw7Cc5XRww8DqZXXvCpL2xtXsJGF20b7Cn81b
l0DZyTtoM4GaEAliT5PLPOSEN7Q8R6f3w/Hm+q+55V+III52HXQP7tAWyTPySeJ+
U2IcrmlJXfBet/pv0RpeAo8J8NF2cXhfEdpXGXKSlW4LIsTKiE6utHZGTUU+FWDS
UnYtWnhY7XbMLkg+P/RSimylPiumSRhxSdqlfbzLBdcR0zslxJlrXDYIPd5OjTvu
h0dw4KUWvpKFGT7U4c/BV7cXpH0PqD06ofKnEls3QCzPhmyTtcAEoAd2DW6yOspI
Kh7zCL6mfLXzbK7nGKvnTmQsJJnT8lo+1m2cK9c8iUdioON6lkZXEzYdKhWyGWkj
5ah9dcEopa433Wjq7fcsI9/sZq08k6IY8ArIlXu9s8cI9biwq48jWyBtbZYC9EJU
y0jSUKNwKKpZisI66XRGvL9rBMqgpKBmm6zM6YDfVaSiiOX7RAGhTA6aUUaSLPde
HQudcyBK7ra0bOgsxunVnPp8726n+iHaReuQTgM7zejFm7smxi+konESYrv4qKzk
kc4a1eweEN6uE6kN+Jgh85k3LsOjixs3psaV0wej8JsYNyJCtJlveKtmvkmktqPO
fBdVh6DMI4cHHo8K4bapR5D1Ou2q6dgpGOR2hN132mwqBRwcfrfac3TMkKauoVTU
5HkaQqqlGu7aHwOi898BbEJcQ0ovcAv+FiSZP/6eiiagS3oMy00a/6RA08u5OeCL
ziu671L0X7wU6kG0v3qvNUWRhPG3eIDzD9THl8caHjWkh753rZc6/6ncs6adwi4H
AXK2wz7a8MaWT0DQ8YRysrKoyDQdQDwSOqrJA6L68xda1dDM55QEHDrhmMXgQEpc
P1yKFmP9w5pFN5qHnQPeZMYNxY4O+9bNxprbJSlWQ3t9cL0AoCPUIpmhqIYye77z
Ub1nD4sfU+zvUfOWlwa+tf78SkdzRSpYBKP4cjQlhOvBZoPgki60jh9ff675/hee
vN6otAQcrohARrhRBd4eBODVXumSgeK5o24AzRDgxfc1bh3KedbGD4YuixEnLzp0
DNxC8DcJkuWzxEnwyEfyACiEdimJH/UtKB1Y29SD3lqbEUJbMfVhawLpQKgmo2Cb
mo4ZlN0nN9DwhKN2p/duPHzpWReOq1LAPshAqq7e4QHggop3uRpwQU823RO2eZPe
dQ+uUI5qDbS2qjHSMCiuv15BZwNg1DoLxmjCrdcjuMr04Fw7qtv/B6fxD9QzFw+Z
vaeTZdCEfKZMpY8IE6FbVb1VBDUUgI1typPS1HMPWnhBnsWe0b6lQ9EjlKJ7TI0i
VwIO9+u0186q5WDBTLlovpi9ueG/HLETda8BisiLiVT3PaKfb1qX5I724DIuhxDW
UgJAbTBvuArNLYZnJCJlLuyJLwyHsytodObpG5ZsjGvjUVPN8MoO18wiZ+m1YbZG
s6sGweijtfZU9zkwF0VrghoktpmatBLSFywd/an4M1EgI5z7ZPZB1RXwgz/Me2by
JtpRMtN1goiZembSbGRBYvqYCRw2PzSVafeC1tBIOuI/z9fckJeOvrgU+DHefGE9
HVJODOwPdY5g/UJBM3A0M+nvn3fDihqGCz1fByhTtdxKPj2B9DHmy0LpGhFcOqFJ
DYezR6ZFMBGltAod5lV5bN1ZRXOJW9rmDO2H02MB/4+icVMcozZxVVHRrc8ZbJRi
Oz/79s3qNuMIsM1xWtVSaLqNEZaxDPAGbSolzbC3MFs/aaUK3H0N+fue/zFFbZPX
ojyQ/vS8GFTrJVOia/TINxlQ+sQPsgMwDqzVfAB6vMApTshvDol932esXSqtkyVB
Ar1TvToKLc9pwiIzBDvzAxG7C/iGz29VwaTJ31Y3R2fbvUnugLvXcdayw7nhUq2Y
q06fQsLihXbEiukH878hzw+sYmoeaGwbIbVD1iwwDv0I0CvvlCtkQllaV20lnU9U
ZrX2gy4j0dSmdZtjTYiajXwP9afL/zbAbmUUGCWECQatzFvPUwrPuuAxuVUGYjjg
HPVBE9rHC7IWTr36qzA9++Ogmlpf30RwdYLERcdX8ECO6kpKB9sx4vL8snE1M+v7
JT41T2bNckWRtN2b7ieXxdsX/TWGBTSZnXRXf+mkecS+7+QXKNY1w6zYV8+pM2sb
o3+seqeDvSM0n98lSm3x8VKPxD+npmY58G9agOPWrrqtO2GSNwc2/Nmj8eSeGCnO
isuO0a14vGINgrRT1k4fu4E/Dfz1YsmFnlHeWfciua5OLBGOHEyE4RkJyx+O7XTZ
1J9XeNPjv64NwZv7h+eu/2J/x9PG/P+K893UivnGSnd4rBQu2pUZtGLd3CbiCFyo
nFkvxmmr5BturWHnTHX257zHhIxDLC5Ts8/aavKrljfx6Mrtv/hJJBHg4fKAmMiN
saPEqDy80Rf4z7TsUuVrM7FtiF2v8FN2xg4RszbIhGmXKIwQUwnnk4ikdCS9PJ4M
SVVKqw811Ol0vO5xn0xnVhTNWRQC1OqoovRKmAmD65sMEh/CJX2Hqgv43s2UnR+E
pRV5G1PL4oxfn3ay1ewY6aAMT+aM4xI1nPd90/tTHZUD1PqdW+fppYqGdOWWngCe
s/b9EgUPyVoYnSJQkfgXmyeVnNkvQ72Pr6nnIoRWUam56L3ZhafEi530jR+HgCPD
iEsyoG/EHuEqABGJmgG1q7Jw9vxnuPO+0Lc94u1ZfCYGKTreTs4qthdgeQsk8cRJ
MoJZmQRd7qJCD+YmSOyw7hlfwa5BhM6u6p+RbP5SqVb0PDI6CsoHxX4EwDTpD8CT
T7vbzx2CYdcHbCxzsP/hBLhyqe5A8i4wffdFbWaQ0J3hc5oLqf3Xh9MNrYfsiDBI
tx6LwbiETHhC/qHgyFsyCAkZQo1/HWAb+3WRR7fBc9dyRmn6KoV2d+xTFj/4NrAI
L0TjmrAZWfpEJ8xEtpl9Nf65CGYJWBdbrtLgotZgSdBEBhIWEGKO9AdZnjvLMA/5
tHwZavNiMmKdMpYzZMAivPcz9AciUDNqMceLL/miNleD4Ry5UFTa7U6RHmb9bc+X
/sqW1PFd//FcKAdvwm5/ngSvRh7sNfdrL/Xfv3jaiYrA3X3gGfQKkcDPXvJ5P8i9
CmBLqkInx8rW4Kcx9UfF6m4qLwsctBvvrTKlEtWdTsb6sCDJbm8LDVAC82OltGvY
CqzYKO/LAaIOtPpqzdDXPD89U/msA95bH+kPMJ559eexbs29PJ9JZwppOKzxyg6Q
MwAj0Mftbs1FT4sjq5Sxv1xo1c7KQx37bBZHXV4tYu8H2o6iH8dOWdKfXbz0CcsN
dlFa9A1Ku/SOm05750RrLOOMy2HsckeQXcM57l7oDWSJOmjSVCYnDpFm9oyUFZ6C
/D5TUpN94cNEuxvq5pvDQzytn1XGymYisxDQWvhL8teeIBLeOWI4c9K5kLaraTG5
iIZBEAfD6UQvyeHgmfku9H255lrZu2AP61E/Nuive9JiHCiXXG+25zCOsXRhzPVC
g3pAl13b+GPo2AZXELRSv5HjQ3hqTNUPpD3VmlmB6y2hie6dcw+Kip7nuvUeGI7A
TtGXWal96Ygm1hGLj85Gb1St30PixfYkNeifRhMcogXMF1+tkbrSs1ZZ6ZEcMdiX
H20RrOSui9XztQqtd8BNNHttHw7LDL2z+lRuKa7M7VkmMAt6sXbl0mh06W1V+k+O
FatZXYLTdejYY37l9QhjpXB1aLYaF2eLerMdrDIwxorN24PdZIo+tX4FtVhBxKj/
R/a7Gl5MBQTyjcoHBPoeZzziRgbZMuHQNhOb0rfKLw7kSrTca9HnAJXTNtFTYspx
ZSIjx1lzAm+XK4fQm6vjZ58bf3xaQOvKXsic0fWXQrCwANXWN+hOl39/19kpEJ5B
uIwJpvMdy7Vj3xB2bZ+dazm8wKgNdFjJuz9SEejCZ4yU1w3QU6H5Nu+a1Cr58gFd
T3WeAiBjUPGbXq8sxtsbV2LEvY/SgvTy1sdeVb/mEh1RHahd8luwl5VJVt4YmxiQ
bVrzUehJuTgCBTZBbwVXqD/X+M/qfd1SQ9I+JD/F3gtyZ1MvTgMH2tHh2TPAH9Hi
isvaFbuae/VsCRc1S+Xly2JUmldlUO7RYml7uOaNy3mXcHJECbAm0hUoHPtR7ui0
Akrv88dPg1hcFVxFClCDYrFDRM2VldXHbtsyDST3zChHFMdp2ksnvvlf8oO7/+V/
n95zbbUVdhE9xWmliinTHV3mXfb1v+Df4JNSqrGln4FH3lPd8jk0QkzlY5yJ++Sh
+ZFuojox8T/ny4i+caPhNTdgfgnTzmMqhqr4e+p+aiYCiyBBxsBzyAiG+ggB7sw8
rGR9u9Xvp08PCaqxsaRt/viVuYs5j5gvTH/+VM2f+nbJ4bMzviNsBtP/G72h7G8l
G8GJK88PQoOLGbI0fNFt5lqupA/fsAg1aeXwwj/3aeMD3JCYNDlaW/9nhOF4gGET
nMQKOmbvxLW2fokVl8bKIYBnYrpBVfSQbahlZRSIPhRTzNtinMUj+ijGivkTkytf
aA7vY0VQvAVZihe0TjIDsSGh5kaNcljqyOeyVOx+RbUDzQ/wTdDNc1EkWsO9jMz0
Zm1lR3ApEdLRHfMvfTiLqN3tqTxn/N5vFWqAoTfjFcM3CESziJEXVWTOiudS++JC
9nLXqv0GFmGdwaYv9NRCL/at9/L0en8UccGZQBYui9/pUpscQqEyqIvzTkwhaqBP
AZWxYbiOzuW6qu7q/DWTatlzo7O9F0P3Pl9L4SfXkyU+ECa68c4fpEKLUZH4DD8M
8dkcMVVOdi2xdbUXRibRbqG3eu9lJFeLTJd21DNpyEzVcPPDJ7cz9Bc3wotOFK/+
i+X3aLPSX8YEr38Uzq4UXdQz9/VDkGo63bBIOsqPd3oNJkz1PcBupjihoA0CGoqD
ITe8hD48CtfyP42tT4Pxvs0TF/OT16+5iLTuSmViNye4zu2NsNjDimPDjGAlXR5e
7letzNs/lQSzsREyQBfS6266FD0xce3ndXjLARjp+ERDGS13pAlkeFf3NQBOZTUO
TKsPFytQV1byld9xFnOkTF8W8CYros6zGx8VGGbe99GHSHKZJCoT7Wf/vhn5N41r
pXai20+FP6VShQrDexdwWp4y5WmhFfMpEc/83ufHhQnKPD4NyVGLZ5dJXdQvfO69
M6hZVH8BHRoCokq7SBYO8TRseHiQCnQ/Tj9eqV0Ie1pBM3Rfls3Fg0jiM+hHP+F+
ryR+rX7OOmDhfVceIhxUa78YgqVYS7QdUN7QMbn0GbI4t4WR5AZ2BwkWnXas5WZC
bBHRHXq5V6yZdMkwUPLVZYIsitLRQsztMszIyjSMGg9LMvBDarJi0J02vn/TFe0g
xqKF4DojHap45ucrMZusKA9nbWrDM0r4RyD9cSE5KOdqsXlh6XU9ls5n673Nxzia
sE7MPlob/BIJdJuXSytxumIGdSHk2HPfXuqwJC+jqy9LiPaY0+bj0efp6UPkjXWN
/cGR11WSSJi7gyreth4Ewvt4iI7bcylXuIrEGztNzhLUH8YUsv4aUrSZqf7RltEF
9VfXF81CwVqE0NsMpEG8kGfiTLqCDsM33v5lXZ9m6HRcIh0BOwolAKjJLV7v6cyF
ZwCg84SwIaoZYy5tyyTVeUW5fX3ETO5eaFdis9nuOaHXn72rjbKwTN6XRj5W5QZi
UkX9ut6+/YhaogSe/t+zeVJ9WtOw9cZxQ5jM6es6Y2i+OlSmrEB80fhmSmOD8Vd+
JO61fNsRtcpjJdP6ee/x34TkM0oOZVu6PkZFnUwg/KEGqDsQKPxgFZc2PkXK9/Li
a5r6yoOhO4K4n05LU7LkuXYEayD6i2Uu5Pnijtcmd8lpn+TFf5imp7b9TCSmEOse
PLMZRbRvBZm/1WqsvLSg8D7nffFpJ8TwEmQHW58I8raeLMjiysYUj7juNYWi+xxh
cXwVICYxkBpQEWV7nqMRRBHooQloNJhFY/EN1gzYJ4OztKT6GMvK9k37PFQTd7oa
cV9P6cBJBSFJJ+VYj02WlPOakYrtEiEKO9r3nOw+OuPD6wZLIpGUqM6u6Bz2MR4B
3P01em8DrigbahqSfALXAt3PutfGaOPOjPel487tw9mhf0NXS7AHpK3Zs4d7BXBA
P8z7usM/4BzudNP9mQx6fYoSyHvoWtBxXL2pbh8WuXVwDZnsKCmAj9F0PQEPDB8h
tICk+Ct3cCqkBd3NSfLwl4Gd73hzAhY+0IDO8L2QP2qWz3SNgTfAjXVA5hFNVThZ
IP6P7fLX6QtGo3Xaq8uOqb6/sLk7euBOUUTdV9ah34HgGN07TY0CoCA0FXn2zWcl
UU0UJxc1UckIKrST0IuV9rG0slkqIuPsy9qyHF9C8jCbntkKdo62WRzkRwS5pbFk
npg/TtAMIb2TfDXo0Z9+wuv7YWnmug1nyldjWLU/wIKykER4q4/O27//nAb9TMWw
IKLtgdZIGvUOVoSUHybYV9yrZND33lAx0tGGuxQstWmrQXVbLel5ozcrqvxvqpct
ttDUqoeCh6XDi7KBtQBZtk3q71nf8zg8SR17GNZijT64PjIV+W7fvWUKrHl9EZMS
nf7zFVbMkfgSLd2uxztda/SLhP3bjN1N3O74Awj2t4g9IA6KTAeX1cTlCPRf9a08
ZWKOSwogI5BWwwdS9/ZD2wz96qVi8XlP/MEFm2brs2wG28jCGaKy8zmNOIJVYGMu
kZXFMWofUhwGRI+vj3t1H0reYlDQHL5G+HUubi3f2dgszu+NRQrKPXBexUfI356G
jw3kQ/mVOgjc8+N/UnOsApd4hLc3B0rk746hFMXiY9EhnkZq3KZi74xOGSAUnH0K
ajDgqR2ZX8LQPMcYSXnXZUrti4rtkL+JOfcxANmXnTChhJxcFTwkExdIrDYtGl8j
ZW9/eCRq9BsWHGk9loVweOgB8QCYgVzORjfAQkadx3ECfGXO8LmIVUx1sU7XE9QQ
LFR0BAM5KltCbQ4KmcVoNkFF3a8XDKUBZOXjs4Flv/G27kKPjyxkhPyLWP/y8aNC
5Fgrw+PpEFR7NPgIHqDVRZRT5eAowZPZfMrYb5F4toWFV/A+9skDfktD394SdD0x
NanU7yVxAjesFSaK7FTN2h47exT6GuLdM3s47SaExsEprYBjA+oevPvI8sSeKp7M
7LwdZgAtEMEaQlwBoV4R0UZcIVdNvqUetyhfSs46iQCK2ptlFaHtFwcYFIxbD38k
AslLt+s/3QuB9mdgmR9Gl5FkFZJ/q2RYTYJ86XlySZUdVteh/Tc0HeY6uZy80Tfk
hvIsz8QcO6H33LAsVQPfnr0p3EgftD9FvIJ/pkNkDZ+p3ykOrkJyJynfj7cISax9
8x2j+5McXG7PMqfOACehoEi6RqgEPEj9Ym5uP5zVCy1zbKq2jLe2316OnTewifEz
sekfapQYcWMwELEK/jUdvQZAHPZFTBGvwUSIHzcH3lZsmu4RvV1Madbgw4Icvfoi
EunMgUoO/QwOVR4wgLPx1iQNryxRlzjjGKBe+IJHtGoWRvEsv+ZruhWL6GsZTNuZ
baQPInk2Q1Zmz5RCQaKT3WDTmfbtHtERdEJpEfrqAqXm699qomOZihfUjnD6/5RC
3PpfXqaLFW2YPWliGqj1e6QJrkD24/K67OyjaRC87wO622rNWWRJSMUqWehSkJv5
J+Yz8fueGJ5uh/WP8TSLXIwmBSGKtLIONWIgkjDrJhZdkWcQTfvRnXrtwZDKvsiz
KhtBQwEsGXua0H4btX+Sy7QPBjaG6tM7uS2iC/wlEZBWdeBQgOS6v2PiD/QtL/GU
a+UJzTSpHz/J/qMx2G3ex110j7n9VEyOWKMhF19TxA+LknshzkoAPLuEvV4cRmjm
cdPX9zuclHrwyEJZYjzRe1PexkoLmfMZjcWRBL+QJxhCJXKsm1VQ8cfeIJKN35KZ
d0fvrx9P4La6HUEflHmiOolJlCo6zRP2gTXznfD01282uNFBW4b+VEL3M4pSst7m
J45Um7Doem+7wXyF4ajma/VPuUcxArNGTPFGwLEjP7NYqaabhmZn567lz+04MtAi
D9suDRBdPYuwnKdLBUSVsyYhH3rZO+7K7KWWcryVpp1T/gIz7EoZP7XHKY50szd+
Z/JwOJh+FixWPUoaS1TsGQweHpOzofUhmhfL5mXNTMDhOzEDCdVSwUrgh7csc0/9
54CKqYHOtSxR1lCdPf+65nko/g50T96wul14dr+ke9eeLgE5QsGNjcpUHttzDPZS
KUxzET0NvXZGtVnl39plwH78DAY6zgmDz9p7ubdOm+WILEWVmAwX4//2OsTXAwbq
Cxpmp0qzSRbg0lLyZ7m7vtAhnLNZ9JzcRCB++egll0Rk1ye1Wz46gX26O40YqxJm
km4RGEuDZsmsipjRHxvUgwXa2rZRso9c5k0IWxQPMHl6X0DojCCJ99emMfWz8xbT
AKGzzzog2TADPducLKndC/EVg+wSdQbK3FHsc+z38xwRZE2nJBunQTt+rf9d+LTr
cb2m4N2JDISZyKX5IWhxZUJb5z+O1fEQMeJvXgnbLfKbSEt0+HNFyQ4tJ91ZvISK
yNj+7ZJRev/ydcUyuUuWyQtZ+fcLnuWbYHxnh2VQD6kPMq9fz9ijDE/wsTxGrlyl
OxzsgBcpbGZy57UcL5ALzWVzHLhuQhBJfA7j6efNMDfM36qZu3r8rHLYX4HmQVRP
PeVhKLHweyE3EF5r17PX2I1KsnkjbAp6ORDgrdL/xXgsEtxNN19Inbe+i0UQ4imf
pNHi2aSdHkgeu0hp2ATAKru/A0yQm8TpQ5HaB+YSdCwV7tOd90f6G3KFQ/NWEd1V
yZ2hKIcouPdI2xzvr0JKT1ONsf3nlWJHx1imBe0BTMxvReAhlNM1D5K+mxaZORIr
Q1A9DSZHmhGXyOnWh3rrf8pigGRKMuHeHNWRnratrr06PBoopc9Z+BfvbqDBmqP0
r0hVKo4pxhYbGrGNKve5klD4J1eZ6i2WrdVVHqaxJ/6gTiKMlSB+L8NmD8sO4cjm
aZ3C+pL8yTr6kDtHS6eYUN8SXkgkAgGwN/6WV4HMeNfxmMXbixPr9t1rBc5ywiwQ
gFMnCDEKAoAMkAN6qFMm2zwU6NtzEEdbvpfy0+/nc2BSIrEg3yPNcQ24Rx/oRduE
BsBTUDV5dWYu734u0GhD7KBqzlS9r3BaCiPyx5mDOnGb9CwSnM6fr9tWaPYPMZFC
5gHd22/HekrTMFT0sRdU9S5IctsO+wT4xH6/hOstgESiFH6zCWIfq5JH5vDliyV3
5JmWbHdPUOsJqr/ZmoEl3rObuSv0WhK5NS2+w6cYno/KHrJt/jncjMvTO7W+Migm
geb+oH3jyQjwwpMk/wqU45jzI8QpcXlJDwrka04Pz1Mwp21fGlRXE49AafkLnITx
x7MY56TcJGRtKdoq9F6xslqV0y41GbafLdAv4jsqsabCkWar7nQ/4O0hHbYl2/NE
aLBWQpinJAYwKSpJijINw6dGRcnCg/7KzbfXEwhaEHctYYn0TWkVZW2cHz0Zv1O2
00JikRi7PeYFwC7Kh3EvHe5UoRgLD8gpPnBfWG3fuL73Mt9NtB8SlsTCyYsnvkRe
H7hXvAJ7KOa7paH5FNglGnAfSEYabKMr6hMsfTzrQj6xkkx1aKKZ5RupxpCSOxrP
BW4lt4IDkoRfR9Uk6yo4ZZaoYiJRRKeZ3P4aOD8b2GmvlwWJn0EIqlHXfpyvuC2r
NhPI1HAOikdmyNbVDl5lu9yUZWD5jAOy5Mze2ovf1ycWED8mxnjal0AfTyr0ybOj
qCBp5X64dUBeGZ+Nx81NLXdB0jbwl0AIAqO6ucOh2sqAhqZ4AlmwPUgZy6OcdRdV
ueQR3A6/Kpi6aExO0bV/na0z+/5Qu0ca/RiEYzxKazYrO51wxxdNQX1/5qXOeEEl
qqp3ll7S6BwbRg3uBDixvlW7C2g66gRPXG9+D4XgxqONy32Y6c8SSfKhqVopq+cT
nMxeYEpwOAqjlKF0oe1UKajcGoU0NqK02U/duzbCJ6fHy6q/hsy9YL5rvbFnz7Kn
EjXWDhztmvlBR6JLx2bDM6njtYssPAqFQQF8aak0H2rUZESXiOOrOknrzYxye3kr
OKqdQ8UkOvc4qZ1/1mHdtIue3ai7QggU+0xb9dcuyvGIGzMQm0xnmrGADl9HHbms
tRbMBxDUwjEdodHsbsh3B2yEp4fUovv2G6oThNZAz93M35435meV5rQEbM7unxwk
NvbtlKSyLnFau+886121P24fX330/ic2GmxACF3HaqoAl7d0Xo804iVW6U82mkap
jlTLb5jkmSpijYpRQaCs5Bn0/GWYlRipJGJeFGn3yq5Nj4sG8ncWvx1x4neu2AUM
AFE+87kDNKRNzhqzclYdOW/w+wWFJLk7RZgpNXXFwkq3//Z4mzzXeE48P9fMQWsN
6n5e7WMPtSeZMoID28FGBXuj2onHU5VgWOQl5HifX+QJ5lL6vKkP6NopF5CNaRW4
WqZlsUnZjwu9RWX5XiGTgpWtgB2SdDktQbTkgGfXbBpIO4FoPwS+/txPbccoO+xS
2MnRLgHan4C3PhrMaKlvh0xFdzk+6vpK+NqvybQzdyHguZuLrzBUWYj4lzfLsQg9
ZjTNuJJiszIDGkhGfOTQHSqWSdio10l3FZekNjOE4ZWeYxACenCcqRUMKJz75uqK
HeNbJJPaGjQUVLy6DiPpKT5l2WG5CGSDCPX8UrzdUW6iKAFqqYnA86xeCwULhvSL
Y55cHnv5t/PCUS5FA3rR0dPYzyfz/fEK2dpwOainRhBGks7i9+7RAuO11CoVx8xR
FRdIaDBdSLDkWfzI1YmO3dCEmyG/6N5BNMsryWZ02zr7OkL5lJGcR9bsYnq2X0Pu
vu175RTEjD7766DmTFUcRRys68dB0awlWWBa0MkmEkkiUbyWylWj6t4wYApbahsp
1Hy8q8IWPU/vMUKxkOZ3u/kQmTDnQnyDM0QGxUCpOhxbfVuovINec7NAZMz6qdBy
7tceWKQ8sNuUh/T9q103eYZkiavCTkMQiqBIAxK6O4adyJN5TtFb8CRqlRaXQLNq
SMmZVW8Qj16rVJLoVeTIQp6xsH7nnIazsXPW0dcoqJ7CdacyOAb+MDq6iGJ0rHDG
amu80sfNCVTya4CEIbbf/PO2lMstktCeC4pdRYslEIm2UXn0fErNKWqwExZguiQS
4IyFRV3VUiAVXHViFvKu1RdVQAE6+/EfWRExFPm2oMD3E5HXRDziyYwULI8OGAZL
DCg53AvCzgvn72vTtowDfDWKRstEh15lKhLr5ha/sjrKLsHzm1Q1xsB7ke4J8qlt
3SfiVINe5FiDwLITnr7RDa4qkJ8SOFef3H3TjPUtTlv/okJ4Jn/HmO6g9La76H/w
e+9FTeo2dyhGWMsG7Hi0BHRQ80WJOhfvDMt9JngfPcgNvNoBQYWAVXVxGTOBvzmX
jqP3IKx4oQHLGOgP/7Q599hzVfgp6YMVap7Z+oRdVublPrF7uEC0N+KNNYBUCYSV
h8BvpOh2+uWe3YvRvYpVg1eXOWMPqfzW2t6XJ7JzvRK9JA0w5s81YdwR6br1Ph8x
X7llfW75gfAX6+qaripEKNdWeQyIpzxkNS5Ig6QlHKCICw2RYnUb8ezuKBXZvngx
6kuvp3NaEb+JCUpEQEktUHac3jLhE3GgaHmRcZ9Ewhgw9eshLg1TsWjtRqO53YfP
wSn7b6Kc/yr8/IfbCL1qOpL7f/RMXwPan4+iQqvZypP2buJMuZA/94kGNaos62LC
7a1uiEe7qeUx7UF6CAtgN3q3ILA0K2tlpIHJmBb+JMT1O487SpNuxYS62lWRDXCN
hMVqnjR6wRao11ZuGu/O0BZQKAfdz0lK8EALcBlxz0jZI3AOZuTQ9hPwDHk5xrd9
VCfsykwn4Mm2Ar6oSQUEWxHrbqSRE0T23Q8C05JNcegoKkt6AEfd0y+QYR+fzVzP
qNoo8HE2TdPYTOwoPJsQ7T+spkO9dTxtT8bTFpq6+hISAaG2MEdsK65ZPt24YMjJ
GN1vPZr0SCcfIXpzQkGJPLdSnQzkgwkGl1Jk8sxDhV8sEMWnwUnXNXrk0bXEyCFh
PHYGyxudNFZUi3MkDGIcXYafab4GiWSsJT1nmwdpp9tdYFTg6a8se+kPhZpfR1mD
2OtoC2umgrEpH+teOTU9ReJ94XXVORVLiuk7fGaApluCg9UhO6CJMYm2OKDLvKIR
KFkouH7+fvK/GVJs4JpPgy/AOrTmdUrEWiWEGYcQGFSxjUPLnvlnmCuAsjldzN37
ZJlKsVEmY8eHVzR2kt/7Wb4a4qGgiJUchOOh8Ccc9o8Vyl3n4vzJstrr+4XZwKy+
A3Pvkkgjn3LjA4BI6MPHN20EVpk7VyYaUeLsZNXIYfBb07Y0y22c4L5/rm9fMABr
P9QUbsQz5Ofljv6eLxRUubsFvQ31oVOVQQg1h1YxOs9exQ1uPIY7TDTW0y6uc/rb
g/5mIYIoD0nx0fCsrBqU9W4Sik9ejec9qW5sjeIOp8ebHAKEnKQNhfI3UONop35W
0UUsaa38QdRB/nfBOpb4XS79g9IbuuSsD6lIof+QjjZeLcrGN6gX9lT2qGvth4oE
yCN7a+uCtHEldCiO+byOpi4GT7THpx106mRy45tJOAX5t3sm1n2tHXj4bQc/i2ln
cmXQ3j0YdSwCTycvICEbsORq17Wv3Vi45LM4KmFegytChn4gbh7eylFB7paLPVnF
Rvmr/dbwG51CM/7YGjEpH93Z0RaZV+L+s5iueuk6fXTTe718ul8lkhZHXQCCiJKx
/g1pbLYtQs4kiiTwgLFCWVw7+zb311S7Z52Y4MTgI1Lcl+bqryiopwgZcyVKwj8E
YOs1XbHroYdGW/Pkbtkn1Dhk8/1KA1eWC/wEHnaTWCdUUpyCbZ3MQDx7FFo5kwqP
8X4vIkOL+tUm8NU674rDyTEl7abV3Lpsi+rPNoc9adHQrroK1w02bJvjHwOV9OX4
i2C8dLaEVJBJWmqs8LrtzwzltHKMFLJYmdR17WXE/1qWXM/3fSzRcQPZmNmEUj7/
IDMIfZSyvhYlD2uj9cmxHR/ir2/tE/2TeDhDwCSfNrqK6XtkXocmdhikYv5ZiFph
yPK0zdZj7LsJTaxaveV4Se9tDMGrYT3Xvd+Y0Zt5SdWjW52cM7o/Jma2Aj3Jjz/S
bKoRaSDjvAsxwqB36jiD/j1TU33ojydEJPlViMrbQE/QsHrRamWpf8tQPwULt+rE
D0RU8aYQ0qr0sxhKPyRSPZmM/igioPOMk3nrHEa5NJKnlDN1RjtGYMgD8iBFa+7c
+RHsB142UMr+vBaXcJ0KVgYEuahKBB19ixakRMAtZdaVKNDElJwVxqPEB5bc4Kc2
9/gw80t4kp+WzGrAfHnID0+Cs1rm59QnU5dIanFuXxZzTbesQKz9DZPKPVJZnRbD
TzWPzwYa54fkX8RCF9ahuxBzoQBqLXjfjU88ODHVsLbKqOrPXSqKeDOtwYTE77u7
mQw3fxHXgYBlrtF3+/BKtBoJtbTiOY3WhhtZRZThE53kuh9ab1SZhX996+Z6sMyJ
DOZwoqRrAJx0y35OpkgPx5I8oQqyexcsrj6HYYb5NW5SA1fJ+L1v1nBKBuTBCv96
6U0L8RlaozCOH2GxwJ2wytFQS+nK+FN4kQNgl+gVvK6zoTGZtcpQClEG2jTbRsI4
9FxUzXxbQMZbdNg5OYt4aFHFMV8jt/cminhw6nQvaLMo2zEadi9Vmo+omaoLp8xl
k9Sjg6Fm3FGIkkCULl3CqoBVMgwjUzVWRllFCp3VTl58EiU+7jsk05JC9wdR212b
Jc8jgQV0a27AYSFTb3x+C7ZO8GdkF1G+4ECmtgRX258MCm2ixXulUgSBgWSwMAVh
pN5YMn/QKTAIotypnvtBHKumIphtm7NNpwUeLr63sUR1hOSmMXjoSd9HteHeuGN8
QGMMii0ytztCyOhBS0usAz3GyYxJJoJW60TmCBAtvoEESawTq4eS2tlVaUOQjokY
cxlQbf9fKM2sNnOZ0yr525hVyh7sivhQrt+SAYbC9pZXvmOfYmL/1p+wi2fkltVg
2li81u2vgZt8bWX4WFj1MSOjyCn0FNNd/YBHZzXWWTQDNYYXMeRv8POMjZQpwwh8
4DnNGR4QkOt4+zFxXSFuGz+ZF6THuiPdGhHxxY+G5v52hDquCQCD+ZA6sFUoUFbg
K5nmgFD5GRSbty8Voe5mgdS8t4FakR/BaHUETPkjLhodH+i6zypdpT7WSlHgkOiA
pG8a+LgH4/Qj2hGYlsnukSe1umTHQQPTjpRjiyqBr16aLwaA/erg+oOTWUScPExB
i5XWs7p3rMyxpBmup2H6AqMjmYV1LiD/nr6h5hdYD0oZWYs7Aj8xglck+RZ/XG0N
TUqRgg1TR23sAtgIDuCgGGvjEBEWq0h68YfX6sVy7DHHQ/F3aykjNYViwAb7IPbY
DCLY+HNB9JllsJgcb+P8MNfez5Zi2jwyDoF86uLfUierbezqjeeZRDaL+labRxcH
Mwoe3P2424jBh7Pg+q8uz9bEmh9dUnsIdVjlIB2cUvkAhXAcun/3RO0KibCigUKT
kCZkcSjimYnmSvfO8NKfBb8dPnLxgVuvKP9xdLTN1WUbdCfvOAAryeRgf0rlrSGG
h66qAmoY0+NuZIbW2Kq0SeDfa1iueC3SwJL5FwTtd5ISBw1e7VxCO6Cra0/9/zmV
g1H/fiA4zr8tOwSM3OTt84VeI9KJ74ctwOLIDjRt6MXwvEfCU15o3XfzWp6zYOsN
011W+R7euFNtxkpA6wBSNKUu0QuetfrMHZS8kewNY3+xAI1nBXsqNDf6xHgRiNcT
ARLF6ZMjV6qsXHMM+mnaw1JJXNTl73evbOnSqNv+Bsk43Ccs1i7Md11Xze7a+FrY
9LxM+nUrjbMLli2JYBJW7JTraQwZfccH+42IxBJsKsGSSvaYQO4PRusycfEY+1Fl
dtFuM6FfNXsz6+RAD59htlQbMVgmLRR/AY1rG7LvSBDWjpBA+OYOK3Jdcm+IP3Nf
Zp8VCeRUu34HUgte88BJaFG+yCZ9FnCDrNcViL12rtZF2XYB4g/00mgg8sIOj1IT
aRikP3drUKTtMS133WXgvQFl0Dq+/q3YJ89rtFM1ER/ac0dNKxgI2xIHP2uKLdL6
mCBpb/ipzSN61yVpHGhjfme1Sb/4O6UukUVjOm1W2Lx/iHD6c/uZjYE4IkvDy8Sj
jxyaAmW6juWvhbTUKOZraw92ysQGHVdk/gM6oTMxvNOfw5bNaAkUhtQOagAzmqGp
kgUMt67I7VYBiW1IS3D4I3xu9tnwwDpsvkoKQrq16Oj7L5o03XrBmuPLFFBsiRXu
VrdA3hGB4+T/5e9kevOgmnW+HkE/j1607B8HfhBKT9xLfIiA3PUCdSEcmyWbTe4w
+SXdJhNB9Mn7Ktz5w/s3saF6zBA4n6Fu7hmFm819HuGnniuOoEjgJ8TIBqXy33Hv
IaV8ASWHZCx/8fwCZ+jD0mJ5eoBQxCCaKodHb08woRBrVOnzhbYG4llerJMqLRaE
g+vh8hq95F4H6dKuCQ6URMq8t0Wdw/EpkLGdo4aHkP3f+59u6cxN7LoKz0GpAH5Y
+atbHKp1L5qWWpLP06k5QxWZu2vgDdL+v3al//lSpQgZzZAj4X/aY4sgHcGJ/xBy
9TWr1Mt+BNiSZAwAXSYCQmhaEf0uraQaK5Mv3uYmIsG55cBg71YxzUCoukY1f5+2
armHj7hdqObkoPISjI1+gAoag3q5xnOhH69+n6y7ntFaFcHSyUpsGKfbBr8Ueuce
Cdr+DpkM4DgY5yNILLYD54ecijDuG7a8HAUyAoIl0gwfNcrVJnbKxU1cE3Exhe96
A7ws1QFu5uZ94texgIL3QSY8v/7mqWXTPLIysBfkHuui3oUJjBWWnF22V7QIWwfu
d7MmjavV6dhpY9WQIFRCwkztuSWFmGE01WM/QyY2ECZP9oX5wGYUQQ+RDCgJGoRw
xBuP6gYr97K0yCSHNcrl7ijqsVPe4zsCn6eGqcv3TZ1NEkfBKJnNcWG0zbRp9hrO
PesHnUgUF6HEkST85MtZj+7hAmyqtI4w/B2LCPHsOGfuBtRnz23IY7151DkXnsZa
Q+wu3STgYACKmkTtkRiLGP+FTtagMAeAb8frPdzPfXGR7SlxiZjZW+VUnEh5/Z35
Zz1PUERCZkpkbRauhZuAynrzOoLlvbwMUEyeuw4NptLjI8pt1ZLjy5YteFnfTWCt
05adTBNvTFvq7fc5XSIKxHWF5yPbYU6eEjTAsp4fpWrFPXc8NNNbk5op2u3F+zT7
sCF/WlC0TA3DgIINZ3NjmB2+YywQLydy3RBPJxxDPu3ic0nXpeHe4BxCwewqUdMM
g1lRMOH5Tyd03zJjLfAhbmGXdzKT86Wea7M4BtRISfGxO2WP9aRZFf2WMj8yO2A4
YdQ05RAX5DL10nVyxQKeCC86roy9rv1UUtRK3noQVZTqTGoTkO1pbzEGMFlWzpPg
t+SwroDA7LRfnTfD1Ervg5uv5CvpMvTxXr9R3dnAQJxrzfMwr3AFvqV3BfV7L2Lo
zR3CJmO7CFz3wBgM5VRaEUBShqVxJSGfJfRnoDBZ+fB4sIm+kRlEPUACuLTcQIfH
zx9WJeVBYGwtAZHqmRyFIlFakgweXRswFXzya7VwkSrgaDh26jN+ORMFqy6lWqhh
2aRH/sD9fyQnRu7BZkTV8xMTYfDArANXizi0V3W7XGSKT37IPB85UZSXYpBBovoD
Up7S4focqXN5mMnLWzQqFOlGIWOduflG5OuYeC1cNVlcpDp5I3gi7r5BGiJQVQH5
eBNx2PAwPd9uRJWH8N5ITWxcRXhlAbX/x5RR5oJY3vxRQGahbLJsDD/ENpK2xVHm
3qn9oqZf6RObVxcv1o+yK1vPPtbxQyreAZZ22KW7KEM6HqjvtIpLz/b5siZK3fko
RAy0Gtmf5lvke1ahkpcp4qJHrxhl1sP+2K7eJyi/3WcSuTXuJG25+7lkQ129xUHW
oWrAMi4SYsspKlUsDD2abld2HMrt7+X17tojAyhEkGzFem7Uxjbl/hB/a739e8at
HJkTrxN/VKhBQGTjBCjF5PkJ2SUfpWE5f5tAx8Oi1Dqvb3s4oHOUR63m+SruvO0l
ufoJlMKZZmI+oE7PVj6NPVz4u1VMieWf5oBvIPZBHJZmYZoVk4xYUeleaGcMe3W5
qezcc1FfEmTxWgib1JpL9wTokqmEEmc7P1HYWcHB6dYtOkVvsuLrWLSRgv5Ek0AB
7p2JLrCkU1rpsNiPEfgq5I4Wbn5HxjWBRF3uw7iu1+bpS0NQvbquLl33HKnJWdn1
JGjZBuqTrsM0XwoZZ/q6Nm98Vapxu6OSRKe4HWBHyw5JdPtaPtc4efynXi+87Y2M
Xmnu5fMi5CUcTpbiaz8T7G2uQBZP0twWVnzmWR5MQg1wKjgEPq7WFEDSRuK0xNp4
HLGXMuO3fq14Cl+AFtkBfPA2LVD86WEncTcmUUA5BruuHFpn0d+Ckkhw5BN+PMVv
CZm5Rm8xhJLzrdKHzBVQxE90N67eVeSoMP5KQDK7hilfKoZfQW9i6kt5RtvsZl4q
fMPSWajWYUXvQu8cKkvVoYQwsH+mn1zZyfajuYMyUgLY60vMFfaRLrPJ6Y28Rx0E
wMjUrk5UsraUQaa+1JT87oJwVAjbcW5o6mYker9dg4tEtWVxzT53sQeGdTUZut0t
nmD9cDTcVrC9OWzzV/WySEbQzGjTVbrsLxncYYaCcQLjd/dGQIo0jLOYAZXkLa9z
ME99fDpRSh1pEdydENddWCCrNKRcqMa1PCR6LJPlvo0kibF7Dd+w4qWGlHb41Arj
Q2YYjjYA4dWiHoQpwlxuSs9cPbKLhkQ1fbDKwlAkUYtv5Qy39sajb8wx5iFZ8eoH
YglCLLe2uVU+scKt7/Lxvh+PeYvqW94d7S+v2cowrzTx5QwxWWljyzYK4Dy653N2
aOMIj6cJbOED8dKxVgGyf/UwWThKx/+eWeFIAz5SqG9+GtdOdI8kT/m7ri5+xNez
jj5IE4oUZr0wbdtkWmOE5ShkI7jUdAijparLTeetTmocBCh4EaOvWY/RXWEi8GJt
nSn4XRA4Ois8NsAo7fjo2LQUWJdWULKIsfnRGot21QrQ+dYpcdhAtFZzNVnAACqj
lULKZn3xr1wfegTb2z8kfQNaVyZ3AdWLnQUi6eQuSj5FX48fV4bNoztX+EVUEUb1
EELgVx/scIsUp39duey71jMfzIAXAUOhDQrEZ/iBotnadKtRmDAbao5cuC1rnNJN
f4CMkKspeZ2/6e8zRxwelzRTXiGnJtej3Rj0Mx4AuoEI38YJFJnWIQKEHhghdhZC
HdnaWw5JH+R87CUx17eYRtr4+MYumjAoOtbXKQ5TqTNxF6HnZ4z1A6RSs2ThAlGF
wTmZuacHR9I45RnS+JbfJPLg+pllOt8TXA0jW9y9p99W5LbOjfTQqjd7kLm6S474
HyVEBkudc+EeAp3RhEIjt8bF1Oc00Fe3Y/bLdSaJ8iDPQMm5i5O1wiCdV56x+21d
nUEyebpm43G8IIDPjWar0k5vwi9ACfWIXnkc8Gd4uJdZDAYANY+nNrfv+WwfZFjD
db0083zsalg51o/JEM0ykcWo5Dbr7s9ZfLXw++3MVY52asW+aivbFB7jv0lrpkdk
O7PljPJyzpDnuW9nh6/m7YApm49eeugx4FIOK1aYCwBOjuGvM0iX68R5Z+dTYIpV
huS2vJzKIgX7lmPju8Yi438ITbefGVoPizjwztGaUatRnvBBvYmeJFVksk5fYTax
fR4P3mIb3o0p9ciWY3BnB0BvMN4dLhX5tpINioS9kiNA2gKlQ5/kE5aVBGKNABbM
MeOGJs6eDM/Zu69LSlHtOg13UArtXQGH/6JItAQqEvG6qtMp0pM8zoAhFvjFEkmt
jmM6NoESd9FyVq4AOGIyUpfTMWaT7rckbaphcHHS1rZOmCcsFC7TrDxyiK+MGTgG
XXi95rDIvSSGViwrbZ/82bSwsdzXBFA9WxBFJtGQOXBuyE1oGLGzPxhFHdf8h7U9
gKC9fO1qOQyuER7qByNjqAWp7Nlv6WCvOpVhbRt2wyUbpYiPu3pNb0f72cRIFmSC
mzPV4VJPS+6C3mOjd03xh0Tvu2WKyGgG5r9IGBBX38VjJX6PEwlvLcFOE0MX0PBD
/6JOynpkfx8ms/LOBtyr0qfxFd68SVzWKYIbHVxWHIpq3nVT926JVTquKtt/e4Rz
nFqjcc5LFmUQ1v4bj+01NZotXj1X4xyAEhrbt7F2lFpzpy9WpRTr+gxAObM1NZti
aey+iGaMXw+2h3SWUEzNaIWA6DPL2wgBfvLBmHKBWM/YNBXJdTajj86PRoX3cWwf
uBcszIttg/Xe+PnpkNP7w45zNu8fJPJHpCWvO4RmKaYFHxiqF6bXNxKK0FYqh/4X
p2sjT3Ypt0ke09krjzGYFbY8F9L4qgqE/PzIuBD9mSw/iRv5OVKKAViHtyf7EGsn
XWwtHRGULIoWjStjRn7WNSzwqOMSH2BL0ls0UI7++vcWy33t9hHn0QAMUKHN1tqP
HaLYPvYnuefTXD388a/HvGysqIxD4trOIgburjVp8hyW8c4PpAxPQ1+98yDMiRvU
CKh/48QdjG5hIFYjdGCIjjlYCTaPnHg4omtUONOg6s8rbwoBlBVDmrayXGMtYHH7
TEokBpnrnP4o3NKDLUcWTh43VdgLEfwmJv3Ly4f8o27LjFe0LhNRpls3T0NRPp4j
pSCUU828nhOp5I8R8oDMgnkXRJbx5SWo8Vfe4eGD7sbwVdzI2kSrgPILpdSH8t9y
cxRH3/GNft+/FDYRoi19ybR/lR/B4D8lcNb7e6J1pFBd09jx7HOUZc/I+qtRvQBN
qqBeT7eVQhBEGIntHRG+P7VrUytO366DN1qgxb/JBUClJQOyquoQnqrNkhJIwOBF
nfOoO4lbzun5zQ/YiMaIm+JDB9xGQFjaNDnffGAZLvQe3RiySahPiIF+T0iDQ0H1
Wmk8Bzw6Q98FdB/j/wBh68H4hbO71drlTFVtPtK7G/Of6vJT7FhgL4z/HHCJFwSc
JHyiWizLwwG0SYKwQLw+j9bQVIeBOWyrLzaFKoJybdCBfk/apS4Vk07WD6vajDh0
/8SwXpbeHt3+iKvDxxPE9g/FQR3NnT1QzxMBOlYboQ3LkQZkOmC3PBhF9NW1j0RD
SkNdZ8tKobncqj8lEXbmfGMwX3/iOBUbyCaNhNLDqAljh/XB2Cy/f+GmoB+YiIUX
xG5yCAZusJJbeEJMwytslKNULnSFxCMy9+zmcPBBC8wTbkMdKQwByfMorvJ5EqsE
tShkmelQcp46FBNuVKNx6TowKFBCv5SmeDxDXFac6Tx7fUSGGApT7kfgKAaGFyFF
yH5uyyO9NPKXjZQIYwLBa2ntGI+tF+jdUgU2fbI7h8dM7xlFJbBT2DItr7wb1FAb
TRPQusdLUkq8LceiwOZ8uIW6ERt3B6zev9o7evatYube/tMu0P8Rmjuiz9my7HFv
3AhkXdDpbKsEug3QsExyi8/rL37OrEHLguuxSQ04jQ8qzS2Zfb0CihWHgZZwrJRq
peQpgl/iLM90x2/5nMtqocZmLBLpTy1J41pxWSL2sBRCpHhtNcpBdKHq0LPbqHRc
uydwFyRFaNrcjAmME6wDXOAxGgsAkJ9Cr7UlSsZMiQiZMcGhk6nCrBDTvGZv1whG
YXk2KI1tjA4TutTKFvBVf/yqFTsc17gpGBaFWWAyHgmsulKCrsy+zUQVUI6dnEIg
qTNCLZXZFv9Ud1m1dVSA16LFHBnCTzRjwO4CQWYZ52D7TT99R5alvVuHG2elX0Ug
ukJurL7Vub35dPVwNo9ck535g3LtSKLT1EGUwMtDsbABigDwcwRzD7YYNyi33lTp
ah3xT8nCOf87Myn84L0sSt7SYXnF1ITL3tMXnL8NwUQBRLGW1xuMIQUcqvFwGoRJ
l++LyvqjlVy1tVwhF2njKt4qbc8pCWrChdZ4mQLgfVaUzTentl9V60OEKauv29pK
W/G7XlaVZmuPtpQxoxdPRtCYrFuez+Q7Dm1qbNwHTc9NDralSg+akzlMWPfOp4oN
koZY7uqXTrwoE08mAHdWHEvDYA66pFXBebvHaNOwFuGb2N060gVoPXkydts0NJVm
txpxCI4J8Qf2Sp4bZX6AKwE4+Srfxu/sD9Jabn5xVrL7kP7VrkrRoNPUcNmRnRFt
qmG7rITDezmPCrUDgXOUk7/svsVfcJRK07D/b4AdVAAK0qCqjlyDmv5/YAEuoptS
jf7F7HEvpj3UdQgnh7ALE/m76hiaRrcfauPX/Y0/3I07upuAn8beFT9M/fCsrQ+f
VpWGDxOckGfoQKu1BTU2xhBVuAFS9YRS0YlcdeYVtRY2Jio87EX6HdBFtty4orlC
k2mQqNKZuErhYajHsMcNH4Asc4GC98KjgUPOIjeLQrYU9h4T1YeicerUFwWMA0ki
LT+WfQ2U/KEjLOjCtBER3lCRhzrTdy6ejKkFNGBtwYvoLSOXEfSSNWI2s7RrxTqG
Yc1gmkQfjc/mA5Jp6CKMpZJA5y5reP7o+KpVdsLmhxUnBNgGBIBzWX/NIRjA3d4s
FK5HbOC7fho+D23Pc1qaS+DolMgDULBd5S3Nsnpa74Y33HQJLHGsrVkJ2Yz/tVsu
nWwPnEySklGn+qxn4Ob+TP4GUJgPZWB798+fgrosSBQ0m7GD0EkbEKv3wmu8MvDQ
Xv/Mqtp3YrjOMTyLDsX+xKD7eD/Mdr1WL5NHNvtKU64Qc5dMdV2vCynzkrEdmhYJ
lLgBzKA0HhXPpNAKX843xAUBsvSl+oHyE7w3KTU2Q+V0VKcD9HAUdO+ANXk7r39F
i5XZTx2lnIJxPPsTwq8J+CR1BuqY3XaAkkGJVQnWFDc+o450zI33fE5Fkso+HAR/
C+0BoiHvfNCyU1YA4t0UEJhbZRaN2QQ7yu9mRbprHIE295RG5l7MO6y7MbuiXT1n
i+K1mZAh2ghwplmpQ/D0CQhPpYwMTBminrI2937XBwT3zsyw+uUa1ruBt+horFdC
KxB4pHHKCkJYP9RvAwhsCuXyi3S7GduZP0mrlKZZGHmrD1bDFaPVegU4HIwIiKri
4jFwfcNyWc38bEe8lqPiJbO77omtzRJGRKemz3jTqQ239olpb2a7BdZ0liXvX596
JYLkClALV/Uot2MZsngdUFpfgIBocjEtK2kQ6DLaqqKcvvdsXZreqS/ZPt2wzks3
xvZu+zPQDlh4OguwnjPr0FKGL4f00ekgJeKgGgTa3tjhg+5vUirBTook22f3B0R9
ONNDh4mfKyjZT/l9KkMHB2qG/Klbvw68nsgEZTmtRIlRS7Vocslus/oXElE2HHUv
H8LWef93NS1x3IYIoydpaxNlK/ItVecLhbEWMQF8rkWkVL0wZDAVoS5DiYl45OW8
ahEoB7KI7R3JyCB5aQI6pSAk0fR8HNNpaMq3GKXDOPgbQsgCGensslRRhOUwG66h
S2FlwdsJ5C5dNakQtJuQY4eM+8XYw6cxK0MCbPmRXvnzMtfFfm7Qd/KkpB7rhDRu
UFRkI6e4kGt0sfFgym8WqfUbO2QbEPoBqUJXH4iwzzvVtf7k2Tu5d1MbVZ9L9Fv6
VJeGRj6pATNzQyUhZkITN0RSNMYjCuoMd17GmT/tKt1yFkbOau/ge84TkTHAeGyv
svoO+mjd9SfWjiAQjr9/GN/nV18Qbj8Vh6+WAEwD3zUHKlFip3LhN1Lj0EaVzxkC
1qEzrx5UStbf6jhMWfH1kQw29anV6AkZAojCOeH0Joz9NbPIZATT+2R/Tdj4Zqko
2QlXXXCSCHDPeYYy+CmcqFrlpsQtQRuJs8SK/HqN74NzgSomlgVRE3XRmUCmn25X
bOyKMmp6S3AbUH9u5PIC6XKjpNuAkhb+APno+DAwDNGNr88VhriGniv7ANkNlvfL
tqh5m9uvIPYE2xMWeKwOOhy8Cd7L8jJx/SfbMbJRJiK3JKFM/oHvijSOyTC2EVzs
Ue5I9CKjnJ+G7Z4g8N8t2J4ciekxY/EdRXbBBoDkK06dJhHVrqN8ax815bpEGT5s
jHS35k4KrLXVU8G2GolS4Hw6OMwRgav5T7/ZRnciAwtAUGFXpQeVSwC/zsk7/nch
eExY9Lozm23Mt3dQEhRS3TA/P49HINQ9QR6JTmvw9d/KnXx1ZSCBYTThsdE8NYii
3cRLBl4S+sIVW+yUw0fNQdQTERhWKD/kDbNrADFxvdsTbOXn+hSEFUEtq2FVLwyB
4WZG5pBXE7SRUDei3gPFYdK0lUkGtUnI8gp66tROE1IIjeaFAJCNV3gpoOwjF9Dp
u1dv2xJ8jWjGnrREPoBYtxGHkFa9pdI6ehoN0jGhbEXF0vo8YiqJqzuvYBxWvFok
ovBqZxOedRZPRfAKIWi8ZRTJ3x25Su+vnfRh+2svB07TbX5PRooYiTDnk/pEHX9l
cUNyHOvK+Kq3YXSnlzKiP6bt9VsD33w7I5M7kCnaqGsp1b0Uf13/UsGxTkyNiDsl
DVZP+AjflIch33HcW6S0rQ7j8zz12yI61eHhRvjZebNznbxqsErrNGnL5kOjZ2Uy
LlLOtdfBZSzZsn1YNLy1RkTVucOi225iQrP0r6/VeAiANSFmsZ/LtK1R3zgJHabp
+OBdJ+45G5k0zSA44cX8GuHJKEHbZCRExA98az2vQELzFT8yG64LK+FENDYZuNvS
5NLSIWkVz7LttvjNKUS5N+SGg8cFnA0y+Q4dxsfvGE+kaNgVV53Tc3LtQAshJYt/
HFz/hX8PEu6pc8XHSh3U4hrZxRCJNXZYSDKxUW/8NrPRMMDTvEu/vH054KImGsEY
dehj3BadVvQxjx6DDy6JGcWkYvxP5SZ3fHUA+dchHaeu+KK+f9RNZl09aOUzrHqC
vTFwSjDx9YPW6aOFczddZmRRenT/8SeJNJA8im2JNJdDl/KLsE2GHir24krRP/K+
nU6G7XDcdsGd6OX5V+4srhHGtkakq4zvcwWrOqQP2yUg/uWQp+rzZF/3lbFzbXHv
gv10OhPIYM0Un6lvP5LwC19/7dSt+3XH1WfxEFElv5HlJZw0FULc2+sV6H/EO8PJ
40COAP2oeFzqq2ZzwwtGZ5EEmBl50uj1+fOA3SZJCo3zOBXuHiykwk1XSyJnWmUW
ZFnrkXUxt0BMgkwBImG2YC0RbJFCZthY7mwajF065ILjZrqT55A8ggDfS+sp9HrO
XYnkJat7i7oX6Cw4JGQi64B5n4N4xjuh+GuERinob2o3t4xSu1LZqFvK/KLJV1/x
NIlHz+2yywe7TBSXUR14EJnwvkNYhJzsn7TeSTkaNT4oy0P1McnlA8cC5/nAvqnE
9QwCeK32bNdqMdanZfPFpgiND3B6WK2tI/LmuHi6qWNAur/K38rflr3+rdKD0+iY
GjJ4ng49TbHA5GbsX9Kb/DN67I4lB+0LEZwiz5QGnera0q7pVTFuneckEC9i4FPd
yoLXQeC90GbMc6tEjQwAN//Y9B6mwE6QeRvGHfkaKhZu1gwVvzv47kRA9HIKn3D6
VFfX9EjyFuDGOYqi2O3QC7YAV3sbxkD+3CNA2tOQ7qqO3Lq2Lo3UkbRIEJVCZi3m
SkxUOtlIrWKwYisQmQ25nsWbydwQuuC81+y+XZUOkBpt3/VDlSPn01xTO27tRejb
czpDHCo5Vo+u68guO0sgZDTcppKzjc+wQiTJp6Cu0bDHIb7OR9pIJJrpyze25gXA
KFCGFpz08LTa0fFZiR/Ig9J80gyWIrHQV5EL2inOZKY+1M9ggG/nDNZLxQZSXi4E
sg54q6g4/EOJ+8Ie5FuDqxrwaCwrfE1/Rk+ubi6sRfej68M7TY77DS8btBe9/DhR
Aqqg5tguKx/R/DlzcHjWNELsty9DgolJ9Ztmh/qLauRwHH91A9wUDFSPa8uE2d9t
uECjkRofSIBjhdGyOFC3EC8zmauO5dyLEMKFsx4yDOyeUNewQFftYL6/zvRlj8yb
ZZs00qr+qYanK0hnFeWSUk78hy5gu+oAGBhIh5L46UGUDgkE4/p/Iy/Itxve287s
zaZV0NUvg+Hi9GmEzqPAGIrvyHwfDUkBIrQnf6IJSYIEd/d66cgADNMQ6L+tPeN3
Gwezub74te9aaOZ+dLlvi3tPkhlZXJHfto5s6Gt1G2xJZ2UfH8JT2yh7pl11UXSx
iJOgy1pZ8ulAQshZrHPWworTmEkE8bvK15vg94h2bBPkqoMC/8ipuLxY3DwMGtYJ
9fkrCNNPalDJdThz6akgVg9c9e7ltiWRgNqUcURImXMj9ZfA10xBXJYSfSu+UwHH
LTaypEhiIBrafY9G39Azfu9WDyoZEJwVVjlmUAETt/dcH+0+pg44DlFAoYS435DH
07EvK14uCGLqAR/Re9QOX1SqHJ5yHEc1g15hEmcyVAX8CN+W1q+pKDOL5PCfuBT+
5FyrkeZJ36l/Q/LfBvUTOTEmwySBPUNNKuP3G5sCKRAcv+UnEcoI6XphqTKgk6L/
a0WH/jQ8g67uPzGpsrxoMeueJMd1LoX7M8frlUV3L+8zScGDcTzCSpTJn0cuoGpk
7w0vqs79Bl1vwyaRrAT61LKjBebImtqVfU6GicyFdE3g3OS1I7IZ9KfM6gm2tzLP
LKcZxaEPrCT+OGtIN8ywDFaedoc2PcyFGwRXbVfnV0QBy5gLLP23ZoHpNVNfMgOS
bjzJeX9VJFzeUR/9o4mDot8tVuTFPqUu3DWhAwyRFjfdGRlXSWR6nVTGDXvmBHW5
DP3e/mCN3dm/WU9pXHsbNjtHmOAFnqgYuuQFKwJklbzmg2h2vBSXGIH0pf4uAGFQ
6ThPfyg7InUakjS0NQ+XNAgE/CJzyE+7lpYlJk52fTI4mMzQIi3V/gMusAbaZ+4l
vRF/j5VV9PbruD3OFeIhAbZztY5t/+jMWXJo4UJqq375NArUpKTUS0p2Mx3560qG
CXIOYwYjX0SUYFx01BP1Pwi3AcnlBKs0DCqHmkAqxdFpUIs9TvO5LwMJy98m5Pbn
pcjArU4TEM01wKZp2Yp5xxn+L7Xbr73swCbDqBk9wSKjrONipMCja2YDWcEG03Dt
BgtwAoCU4GhoTpGGhLdSrbqNlp17udwRCKWQcAGuRj/lYkXW5Rdn47iN1w06KMF2
Q7ztDO82UI85AKOrDN0hMw2Wv4os/vqb5Hd8z4BnW9Dl7iX1npg2vF0I8nyJHYLF
1f+VcYZylmebJ4cpO54pWdIXiVOR9gSzNvZyUPME+vE+Sbepnrql8Bg0mTVpAxGP
qcRrWww9lRl/e6Bl0URqhxE+uY0mr5UkwRUXH2WL9JiRWfturtpYa9TSyEjuTHf+
lJz4ST2MXG6urkLs3rBkjJeBolu6jkBOW3vrb0LfJ6yf3MDHYMtXUN8k1dx5PDoK
fO00kFebXQEy1RCC8+B5FKeTdQnjC12au2Iacsm1skN2PZ6G74dsiZvaH2IrwUCC
ohv3nx5jfHoeR5attmnMZt2WoNuqn6GUC6ZARJouIoyPTVISsdwik8Jh0+JrTdAx
OmrtjLw4tpcQhP6PsHGM5NKMvkhZ7VvYXlTkVLg6se3ApfQ5Pyi7etQwdkNWWyvp
FGPnrYzFPwLD6H3T8K7EN/koa8E6nXeWviJsCmnkxry/Ef8oeHaKpLq72e4hEhVf
tRUwBvlprTFKn11YoU5Ukw/rnjHhHPfPoGcxfiIHRc3pfu6okMtdJ93OFsUUo5OH
mJ3hjikPX7uJWNTYEyXA7nEU7XtIlDZqMxphzwufmeb37kc3OzDvCCScWhB4ZXmh
PcSxLIudLf+JQyL+WaYZP9MGyL35KebXPNuVSe5qrdITU1/ggYLzWE1wznrSZ3I1
U6mJ8AYJYwtOL2xDatNf34nH6I9wy6q3dHkAdAachqdpE+2AeQNdT2MYzjSkZb18
Z4t+QaB6fPk+iGf18hkLZCGSjARzITzN94TaEnTGZcPGN9D+8W599x1hm35UEyjX
18ooFYa9IqTg+YiJklrozLiSGM3FrfayCzwbhb364beRPX7dcjO2Ju1B2ZRHe0lb
r3qPRTxY4D4NyrCfc1D31YvQ/oq/O1mtwndO8JED9xwaGkBjrwectFz6ZlVsxLiP
bvszW9K2otP2iKbmPRIgl7Dh4EnbOGivk1XAA04xW14odivTJAvuxecjhUsC8iG4
NtRmt+8MiarXO4DTD12qR/mAIhkUvYf9aiV2d0aHUe4OdD5q4DOnpDFq2dX7GWLP
7AXS9Qgu3En0HFNIni0hzPONx60F8AwKbBb2H69ogDvfiVqV+XKkwvDQh2essnbA
ETeDL2eQEmzJF81Q9VUgifRgPgOua+wUh+J8JX8wcRPGNuLxjna+SWs3y5tr7KQj
32B8wCXuw53QBuGgtgMIsu4GRBBUrwpQQhLribrxkt6JiwIXnJgHTfs5SgYMwoGL
HvNUCj4tUZgzFE2AIjcH/Q65FarORxqbNcEsAvWPCtAkIzgCPe0LimV0L23qArIK
xYlQLrbW7RvDoMYXrQ4DVttpPltJlkUCaAlvMYDaFo4x4e8bBxuXAwp2PLlSOqKZ
NEl8saw43IhFXa/PUYF/zLjreq6VT0n5p7lq6aXDtCE5eJQASKjHxyCDYp7Elklp
15fvvnlBPs51p85X/63/tt7cik2cNzaVz2c7cSN5h5SYou93EXNDK7jB3+l8hoUT
aFN1BTxIbyUkziQqRM6xAEkFzWPJoQLC6J36Z56BiSe/hEQm6eLhtEPHNYOAVedV
zTFY74ADOKJISmUa/8Qq3AFeruQVsnbVdXrtUAhzY3pLGXb0KP6ZCDev+BX0/FNB
CyaKbrtX73/hKy7aETf4TCkSntMl33gqSiArFL17Mm7G6CRICGxf6yqlCnD1lYcu
mM8KuAcm1COU0xsfmQxXtpDig6QhMWXEdhEP8ctUP9e/Uug2UT+qjV+gur/4VKYy
4b4MI25EoACjzhix6gLf7r+mEJmaKUB7sgXV1AT4UhA4gVQeB9B8+HrB8VUktSyy
KrqIpD2XK4CAE3ufLyKFw39yEFTvGpAHckbFZ98nHqR/LqQmv44xATwMjRK+sOzM
a+qr/kxlhUQCW8wYEhkbRzREzuyZGXBjLyVFvBJYM6xzpOOUR8ZW9s+XqIvwyYho
tfw2Dr7HiftKk2n4jsfnPaqBegdmEWXS3NPbDSSYNKlGxbKQyv+m+sXmLsfItHxs
I3FFYdRTJFyj+ASy3uFFYNXhgT9lyYM2+OS085zcJNEF7hDlYAN3X29hf/9FFtry
hcXw+oUHD00REcUMlIe3KvpHuS9nNha05DD3xykCGziGoJN78Ha6pxXOBIm5fpEc
MG4AV+5E733783/lhr78jRz2jt3iIOPlnJGyteQ3sUh+jk9TUm3LK0bM3F9dKplA
Um1m4wr/Woynr240/X5YWLY4CFh4P9pBpmhF8U1Thml/a+im9PGM1J0vqOuUbPqi
tEBR0TzzcjZqzn93kTlLQfQ8JTijsgBoEJiQhP50e7oETJHoY1QLqFIUL7sG96ig
RunxjxWkajVw6VWvb+LvaSxuPLBR3dn6cqHATtciJ8Smm9hYeNi7vdsa5ifa6WBr
PYoNcHHRFg6I3CJ1JImDGeZu3rBlnc2wvA3PNG4ihfBCqHN6TwPeNl7TzBqlTv6M
nwM1GA2lXIzA6CAUp//GmMwZY3dB76yaJgcgPz2T4/EkdINEs6WarzAcNiMBarEC
33elBcrGbojo4xIFPOZHRqpXjQFTMh3BqGJ35Y+lHZng1VFAboog2QEQ24BCXlM9
XYJU9nzf3U6UVgrSEFRNwOUpOiYUIgOeOCEHMc+boH7fV3BI5NkgoVIG+qyYB0A6
Ug6KO5C+Y6ZXNnpLSriWurmqKe4wZf+JO/MwBWK2zdVpvI1lp4VKsgBoAXkNYYDd
yJbjPQTi9s/hDCmqy/WFMdU8ywOHhs30y+dTPucTkwl26DEMuxakDDL30FnM1lVI
1u5QCOWA7EiGaOxvuK9osw4NU3zN6gyU083Fj+JLPW/rprUsBNtJ5fDX9C1TUt2s
KtlhMHZEn6MGxS9d+utPrnHL0W/AVPK/p0IHYx7DHiXtPOkPZVipUQf24Crxm0mL
LYfAOpWDuoO62zTmIXgfUxELnwjAEJSu5b61wS9FI6e+26uMQW8THuIuLhQGek1T
/UoBxiNia9TdwM1ClPo0HpORaZNyhFNr7Tm3qUQCdM0KLzyGmjtyMfq8+/Uwv+av
nJM4+ycaBXBObv5Ra8Y2yAqKdfmodGfCDA1+qlfsrnUb7PYnfdHaLQmTkNnGdYHX
zAy2EmwXVtfrS5ZWjbhlQiMRL5tgnkKef5GBsp2mLOyZLhxIf3uF7EAZVVKchQ4o
yhNRlA93rl1yTXK21WjOcPOJq0Mr5mggxjiVBo9cEGDqCiKkDTU6BYt84UJDHfho
6uf++JOMxnoNPbKsV1kjoTVfwq49kqhSshD8o4a9OlFz2b79QkTGMVQRsrH3szIi
mFvxQaE1U9/YI9dbKG9BWWX11YgP1DGZOtLhkeD9Hq4bNeVPjD/Gh2gIxgt6A1se
ssYRqcB/FGfUOuNelFHZRpT55mfSV6JWa4+Mk3D3wtfS9sAJDpk8A1TRG+OEj2jP
r2A08c+4awzACzbDPLy/pgZRQMUe9/qIaCs4zZvanjwb4V5lSYDyuL6prk7l016r
6PvzuutNlXITKIfPkvBXK+rdHpWpx3d1lqj+xDTZrj/40YbVucZPZYb4kpAFj/Ju
svE0i5Ic4clZnfxQZxaxJ8oXdPpGKGfVC7y/P0TSYfVhKjIW3GwX5Z2tA9QLY9iW
MPdtsu1i1qp9RYyO6El1mO089AvJDcPcs58pYDdbzXrojdPPr6LjeD/dt+7MlsbE
6lYBtHybbIAo6NZ6i9nlRWmK/SHk2w+Izb1pK5RQaOUtfoph0UX5oJWii7XW/LOL
xhU2tmC1Gbdl7qzv977lwkAaT3C8w7eNoBVgHkVFDKFSrkCpsZEtWG3dc1Jol+LQ
+8GnleCI95zvbEMEhuVDUMqvGIsLJ1/o7wZJ5u/OMhPSLebYXhuZzJ3RRaiHkQL7
hUOMjWUmVxkQ9CfTr9NDESIGS9jmZwjnPO5IEgBNxVQiCI4ojDpwh3+/PnyZOSn7
UqpLTS6BV0/16n9ykW+S65vbPeEV8yAf7T0CfoF3uTQlzDy87BkaS7YGzbF+C/qV
4XtQLjasKzai2VqNQwOjXw2b8qtbuMewi3xTc4jWHWwjAvF5NqQ1JnXLtP+opKza
rkt85vS4/DJxAWHBoNG1BiNiPc7XHwaes1i9RA4RG2nbc30xU7Gia9lU9X5qsXk/
GMH17Bllasikfgr0T+BcVkKi9r+XktfWMCh/86NG/sk6+CT4sAFM2h06rGwSfYgt
SmycNnSRW7NS75klOzCQ7O0WXYfYebYdIWKANNVX44v2EGy+8+I4zNIF3hMa7LuA
vRTkq+bB/2A+MeHY3Hlce2/YeL1RL9ThWtiSa7kpjQ8S1KWbPpuRdM7NBpipKVrB
rUSHPXPwNTFSFRz3sytSNi90Yx75QdonhxCSHDLfQbI6XlTLXjlXBMhfp8cWMWUM
h7JugFuQu7QK3lP+ETflrPbfNrFufu5NAXsRo7tXtZEiAv+nA529pXn03ufJ+PfI
kuflMeT8gN5zheDqZCR3L9DHqu63h3Wq5Y5Ghw/lOVqfnJA2T/gN7B32ijxYxLDZ
qDxVkBji9Rigc0C47pujSsg5X0tLKM5MOh+XcEYl3K3mJKTMDBY7Ihh/HQTFO9sM
3JrzEApAGPab38+l/n37xzb4WwlLxduVQ5NllUpFgIMtFTdYZOBIVkvD5FGjhqtr
/s1qVk9cFt98hGVMg1VmmGMre5sEtU2nivV2GcEVDR+03UYoxb974el0rf2qvMiT
6YtbVhHITvSOUc0oAroX6dOEqwD1Lfdzt0TgDMvJ6/NNVB8Y5rvl9a0T58rzluzq
0T5puDWZVCat/p8Gblo2cKTkBizirOzEsOgcZCk8zQTyrK3OvHKJya8s4kvsHcdb
tvih0nm9ed/yzp8+xS9I3HkAhBqBDLygNE9Rzn5oNWpb8rTMnIY/HtnWvZgi3YVv
oMu1tWLrood2Z7UPIsAu8Y2lZxa+9J7P15ntWdUNB2B09+fUD0T6Ux7sxopSHNv1
E5cnvFLG2hLim1AqHXdICAPgfHMg68z7X0vgwfkFyveJdaXFymZcgdhdTsso0Z4E
dvtxSsJjd0Z+HtRYHbS8S/Kp1L48ElVFMnCzzL/y0IB5RborGDFm0a5k5pz0ucrB
X3V02z/51PEf6jr8Ip8oYQpQHHsC5GCPGT77rv0CG5vRVq5v/vLCvmbaR4MI/26b
YSz3kwTMNuRbU7vTZ2E4h7/B8zxpernVe5r/qGLLT+9lY5EVQpaZVEQ8JTm0gPuM
Qlfl5Gw4HP6V4xKemKZJbUiuTqwhosqbLq+gkPmkhIRbuCh8b7M9Ih/cAjLKNp3G
qPDmcm7tb2dbA8wE6ZSSO2vHmyddKu62GUNMGmhNO/E1Pwom0oaQTYTDpClM7Va1
i+6wJRrT9y8dHPftSv7VEWO20dIheVmPu8y/AkXjkFojjRoZudhVWvae+fFeahhE
bQJyFmfeUQeJiOpxCzQ+oDQJm3Kb7WmZUP+j9lm1J7QbM0u7FT7d+4ARirW/x09Y
WpAcD/u8IaVtfwust0gA54DG1kGzUTW/ARM2J4RoznhmH51R4kP0yFSNAk5WFKOb
6ZoKv4/AyyBCZJMyP1NQt7+3TZyXabyjjZf3Gky0CB+vu1J4qgOeUSZxwABkXH18
gcM+GhFh5OrgcB1LzxAAKh+Jy6NE73TzScpIQhx4fp+1sLoQw65YwjPFWgktuIKU
qwcPhNq55mUsJuwIogWqtwdoQVd6S56lcYDA8C+9OXSdKPuNqK/v/V1XY6sZDhqC
Nj0Kd4rUMYDbly25ZXzVd999IDZhgPj+J4gaUf61sSFZpcLBJWz3DZBWOXFXhvcD
q/5zpQdFdBxiI7Z/AxGyfLYUPTh173Z5jxx8Tqx8lqUBpSqYzmJztX2q0A2GJK7Y
sx/r5CQnJd3E9zuXoX2R65Ru392HvylNVD2My/qGZS877L7UJGVskbGLj0wq2jzX
1mdUw/hlOqZZTFFpASrzcUSFp+BjYJiR0ieBsqibe5xK+IureiH5y41ZK3lmPYE4
lonY6wMf0+9qUnviEaWS+ZQDJZuFi0bd4DPt6SPgJBPK1cZUweDbNgRXwbAHboy+
Ywk0y7dhO3WNdinKmjdmRiytQVCLjmxY48zpap+lPCoACl1jfjIQqhYDAqLOhMfm
m2oPzDprMJKZl8lLoQ2HOVXSh0nErSgBWtCDH8YUVtB8bYm2pOxRUBsbhXJY5Gwz
A3ccwvQV662AUXTGlQs8SO3vwtuTT99pwuzOpfat6lpTuuSGewW6cwejweJFHKpP
299R8YTldApyMRBjeEdQj5Phn4n6rm204jpwEcB7XQAKSSqx/dXs85exBkr1TWSb
/RjQx4rQfq1b/Epx3RhfaVy5Pm6Gy4GJL4W+vtIDdgCzOzz1zjHAxtoDK2QSE9Vs
MY1h8K/OkTFaGh4dRcwuWFbq3PSvqsZ2WeQ3XdcPi/6NkTcshu/ekem2NNW09viZ
ieT9XXJEU68A3hmJe3VsaH+IhzQRVNCxYOEWWD3crKFjKLHsdAQhgv/vFwUWcsaP
o0M36WnJg7kHdrxO8vq9eMpN+D1UZkc7qqCbVUFVshqjnRuTn+U0UWFYmhr2gg3I
PjWbcJoYlytdOiaZaj2qRSDpKv+IIr4EhgXsMJ6qyJPUc55kjyBHZf9OTmLMHgem
YSIoQJw0a5LIRadMu+vsrq+n1lJiw8vOaqyRtrmOpl4FQbj4sKgyXWzSu4PSF1UP
rIoGedutIxJnVYZ0bTF7OXvvulyRuF8I+IsgelhSDJM+R3ecYLuPPjCQdvU0Nwl+
R08vk08b34M4oNbDLmz5lhZpvX2kS8I5dUxx/cocURNoFIA4tK8wnvjkEa2LAdSe
+2uhSv/ROUzgJfo9e1QXtpjPHMrs827/nI6AFc4ELHskb9x6RcewcgFmTVF+GpjO
dW643X2ldmrK5FE96j48opSn5rhQ6jmBtcf2ew92TGLuXGWna6QLjZ19tQcXfflf
+g77xDInvfRRN6rJsPN/8T7QLNY87gZKulmmHxoVVe6Y/lhuqbXHNLpuze6+i9nk
PKc6RCpZ3Jjy3lMFZyg99/uQ7EULuquY8gTbrzo8QoyK5t67ehwjrolh2gXpS0s+
EdMdKc63SEhN0PHf2W345xtB7EaSBEc/FGkGQSv1zk7rXr+y0wbjpI35W2J8Bk6y
rdQP6y8g3w949O9oeKHcVJXZh6Vytt0z/QJcAjNkQ433va73/TbpW9PBArkvBvjW
cuq34lMIPBDygKhc8gvAoyjwAyWIpvCAUUThHsoJugHI0v0ce/qpCGEhK2G0NEH+
iNVyC2IBPOP5yTDMBPns22/7NoxgSNIRK9zfeGf53r68pcG3RAYaecFFMpn/WcEE
XYdLWvcoLv2RxRtjC39kikqMaoAg0Pu8CL7mgKZBIXmAb7L6Nl6daE5gl9iGgYWV
tZMxDMhWieJm0uxRpcAAfRnn4A7XgZ0WRRzjfP22gIXD7I9SyZdhe1/uwjQpef3k
0Bl1flpwoScU+hbwVszUtYTPKN2LXPk7ufPVWn60CG3sgXSwSxFPqOEmQwZW9LeQ
fNUUKLVyn8SC0xTLinkQ0rK/ieXx9MqH2/Gi2RDhEQJXkJSPo4au/b5xI2OVevv9
9NkUcCi1LXUthaLwYbNFwyZ3HSToQMsWlv6FqJq2EB2n4IQ4hAGGKrAt4Znvbr6J
T/wn6fbI6iHbWWoxInHun2SPhMhCsX8PiyWhaWvWD9GpQWuL7+DrF0P197yXDkKU
5brtju8mnQ41nY9hDPdnrUi2oQdtXW7IDTr8Zr/2181NIg+5//rLQrGMNAh8QLwC
O0/QiKQ7gkAyJPWwx/jSc9AMK01qVt9GMePE2rdNbCRef2FMz6TN6mJtdwQzERcK
dJsTzFtLjkN91sM81Cz2JldalW5I36/gvBBCxPNR+tutIDjIAz/52yLDrGxzGGw0
/v7iA76Yfdp/7+Vz/f7mjCop0jmhsz7FXQEbYwrH3FMyY8Y/mdB+7PdhSzIxKirV
OtAAF5FHSm65vRuJCsKSnAPXcPapDJr2VLyHpOwFzzGm3Wo9ohjbZi/Atdd4ukaT
sAjuVfGJLZwb68AEqtM6zuispYbtETojVGF1wSeYu9tUZ+T1+Cm2pcUkRN8jEpxX
SVd0Wpp+fufSABmdD0j1BUMt2kOfuN2yKIpXNOgAoNohcJ1PubuuoDaz559iGXA5
hZGHMf414hVr1FvWmkw/G91VZ9QTGHlmWDkOKY4LjSYZUe1FzVuH/aXncXYzR4FQ
FZHQfPPvZsFlpxAeC/eRMW4nfEXE+ulHc3GkwrNIFNgxgihTfyHuIUEmVnGnAE0g
7Z56aaHE7FZg5+m9MsuwsUMO835dI73F3sXlE+WKouHMvm4K5C8RH9DGcbAN00V/
1ZywZg0UKy65u3g/jue6dCRigV8hOZkgbPT7DxbZvrcWntpienz1mJ9LCWq9cvFd
wR5I6VeuKSubYsdF9VZgvXb3jPLY3bxjSjm4Trr9a4PilfHyeQer1eyIJRrpGgLn
Iru4pvJzU2BX1Fx8NoIUDvSW3YLH+f48cFbQVSl6iEJN+WxLTm1y/AWuADFhO0ZZ
NfVjz5gbVhAsbWIGMBen6+FXCM0I4IEzM7dSs7HdRUKfu9QyRFdTK2wYpBQzNuM4
5Iv5OUOMctyYLeWRho3bHF17Px3ovB/DUn9dxtersug6tusiLq+RVS9Et83bIwIF
3VyErjrwbCbXTz8KJktNRVVxPuPMoJS5iLMS3EF0K8HB7RHpJBd+dD/aAD+ca6ux
YceOiszhEno6Lxn7wqEwfnNUtjMGZ6U4Dd7JbuAkcMj1A5dJ1FyEGnk6+V7oWazP
UEmD4Wv7XAyPWY/mUHe0R8YgVUnzezgd4nUzlVEM5Dvi4d5AdkK6mI8lNTTmkKQX
HLpoTOKLqoZl6WJhnUF0nTBzmuVSogPCBCKBCu12tvDLyYH29ble8CvsEXKnBiLj
xFVNCRCdmawHmQRBHsQpP2cU0kBLK83iheA/vK7w2p7M0VUud8S7Yk28AgDBVIDP
6cpAO6/kQisWPZ25rd/XZv8chknrvd9roXQy7NXKINFuec+o7rJ6RcFeqmr8Gefw
b5+3k65C7xkMZuv2dLoyUytz3xl7C1wy91lfHmQkYVLiaqEUWjzIw5ZODOPHYyB9
WAcskvOR23A2Jh4stOzBywzfqhl/qaawInryfEJwmVvk6NEUlSWAnKhBpsgRXsc/
zsblvtCq6q5Mf/wDze4ANofFl8gAeIN5h81C4ZsRwIZhTh4t/mOo47irrGYIvYVe
qBUcaml99xIjWP5GnRb3VFZ8fJalTVE1D3PZ761cgAzQYGQWhIJg4ZiTKpzy4sRp
uQgXbqSVsLQrtB8EErDPK50KwXiwZllHDEeJr/uxLbhs98CEdMcZ2dverYe0Zxx9
LClkO9mLwESQssb36dFOLJ0XteUGhnbDsFV09dLwV9g6h/xC1fxwrNIH3zvUPFNo
72+2Q0mvmFPa+AAbPFzWBWgso2j4LQY6PKT8SuDT0+fFabd+4R98dCmvmYpEm2mR
jifbG+Mq6j96LSURmMpOPQ1355ZBPfXKInesi12+1SsgjaIp39sC+1dCXsRYzo9p
U6m1MILaF1CyhvHSpOgnsS7YFqEvr2WpI5/nAe8fj52X2rwaYERSm9JWqn2h49Ut
95wbFmzL72NWxyLiMMbsun023XiR2ZXbvyECTpSwIMXMKWv9vLNVWU04GBpuOLlR
QT4U5jeUmZqjGWNgtJ/7RXgVHTxejO5sGPjNq1zjdOHBUdzx+hT379S5p2dtuYPp
ZVHMMRbSukX38KfDC8NVgRpZhqdZkoOzvBQz5ctqg+1YSqYzAL5IbcC6+gw/frev
f8v52uzi0PbePsJihftCnJYXANDd6N0rnaQ159uRrK9JZxZvSuCXeNQEyspN+2gC
qrxZiqjD6ek41yuV1ARrQrowRYCmCcV7d+gAf86tVa2NpnRYabpy5aQEpQ/VQOEN
LhzGOBapNn9HSPVLUUOlhz1Jb8sVAi/TW5n+YKl5lVggQWaT7kUA0cxhKJIfDbpB
OoPElU5v/wCQ9LOlDaVgWdii2b7zRo4DWlIC0cZq7zCtAiErfSGqYz139V2GIf/0
YhLIDhbOyTxm67AQ1QEE2ZKJVEgEPE1nZxQv2aTfQq0wTRfkx0AOUmMQsiQh0ChW
3F6HheRY2NSbunQU7exvGbXkm54jn5GW6/R1LJVNdsE58goBcoDGoBJtmlPBr7fB
gM3eGgOcDZS4JlKUUXlwZWWlQgjA8tIGGz2avj8LgfKyEFmayHwSh+BN/IFtltAp
JKDuTFTCMGyaWuGT6BfuN1wafWxIKfZzY00CfdtS8Bvrv4QvDOd3p7EDG4BKNhEJ
BObNoK8zt5Y97CwHdLSxso2tdTZNaYCP5TfB4qvLXLddgtFRM2VJSmasXqm6KisT
+Dy2Q3IEE675sXH9utTUvGw2ksl9fKpNNl5Ah9W4mx7MkSdIxGVxjIqHCkC1gXuC
5uEzzxnZN6p1Q1SUeZ7U74pYY5MROWaWf/m5XFQcB5u1ilbcNlHWB2VlMn6ukqnO
a9ODR9prY+SS1oCpgMPYKCQFiIhFmfEx8vdwsh9Yo4H0uGBs27rVJ0N96ge38rja
CqIhOEFFdoLhTFUls8dDn1WyNY589dIm9t+B823Pz8czhrIRHPmFNuk9whzuT983
fa+gw6EkjEjGxT0d/aL05w5sdG3Et0QPNiqBipCZENdMJBpTk7vfqE2CM45JOBVo
u1Qy7KsOKxwpBTK3fYngK+h8vvShX4vfBpIggdBNhXYCNBjDRXxyfX8HNlwC671F
JoERkbXwoKhreBr/N2QNLIKQB5XP7WYAB/u4NV13+Pf+seYN51vW+tN4HLUp0YD/
AZ99HaAgStVv04Nr1jAu00gAI+B17CC9tfzcDaqF1E1kC7prsKnBVeLyfbQYRgg9
10+M+h567jCJ9PIfX0nByV1oDMOGYnbgMGI4RrZgFGT/Jm7Nm5xhgcBbxtbD9c5N
IpyxMfE9bg+PfXsmVJbzFlBF3BZ62jC80nw5qrHx4cFhE6ONxKx/FHmBKtojFDab
qrtvIEs6X4unlhRu9aGMUhgRzFuRWvr+ciY4iz1lCsaNcCa41eVIpVkWqIDtp83D
7rP38L2RmwmPEE6PerTQkvjbgGCUGuJcf2A5TeGEu6+iEcpmn2LAXPaNmYtKAIJh
cnB3ROOGFwDCjKzVJQA5No47lqMA3KgJYAzfkBfDJu4E4jK6WMt0HYWXvSA90STB
b0PsmPllKf/puFIsb4jxkvFPP2eeNvuxC5lT3g75Q3YPmY44rcpZz/aBILrBKVIl
q7BqbjZXER2y2zFMIA4h6RccwKCnFs0XdGtzFgQlfVFp5iY3pnDb0NxszKCHfmWe
Byg2TLjfb30a8avaY1intRO+yC2MYTJtqTyeWfcQpyup2LLtQpDecMNaXXKARhok
NQarmB0lsU10T+mjJFVAsLlGUdwNY1iulJWGd8AcIDvIxYagxM5oHuwNCEmOHae6
kgK4rcc5k5s8hMkUuXeJoLP2viqSu3seVefIY0D8DPSWf9xVMS7nO99l6d5Pz3pe
lOFTwyoDV9DK8b5upStm7Ozkmx/Urz3Rj/GOGZA2OYMI44ngrLLMsDmy9nqrfxMb
kMF8Yul8nWBE8NbSe4jFkQ5urpuu+vcJG8vtMphcXJW8Ov657wSovLx+66C+cH6H
k4rv8mKrN+i41bEdGHRx3fDQU+dv2E2coYlNVaK8M5Nk0OtNLPA488rKZuHMF3ty
7DeeyBqCI0NKQ1lcpo7pZ6UKvsT3iQM2hfOpZK1d5Qjt/GL/STj5eiQ5XtigPfa9
jdIxE0N8nHxBA0sFjTr26ocATv6QvCNcAN+l1smsbzVz3MA7rI4lpyEwEsuXjPnw
3taaO4DrbcT8fplIv4m83Wn0FJ7TxaLUztzoUkLeLJjjGCCKZZT7r1u7SNf7mTsi
ojHWcgrEw4091Q4hi+cWoHElM0Ww0edAgzI+SZXLqa6/4U8NnlW8PhHzwAk3roR/
hk7eRpEiVp/EfARMwfgE7R9lZR11VJCAxzlpLnBFsu2nVdv35YmAHZA+5B/oPnkd
KZTZiivM4/jYBi/ixkRafgryRapPTujnC2UGs7qBb85geFArKhgD9Ie1E76IhM45
zJk9fG0fhr5A0P9ggo1AOUuM1iXWLPexf02ek7kqeP5cXRXtnC/EorzGk7p4vPgr
kcfCFiCemKQFuBAJhQnkRhaFpfPtk1pOlT1yQfcCcNBts9v+1wf5dSuwTNM8+nmE
OzccEXLy565zIbPDLp8Htrs3ex19fYV/ZTcaSKfjF1J+XriIDyo7ux1K/OjNpa6d
DKeB8bvn9j4PFpjbLw3HJ+LWNWrwWUckplYUlKFUK8lA74TXHmL/ZVr270soM1jv
zDbFH8UGKkbChA5QlZJWasOe+vEvWn9Y8GdGXkijEY8ZNfuzFJjmFPPqnUNBRQT0
ELPRvDcp15M5u+SEuYn4vpL6muPORnIcc93YObXVJoHgLY0Y/c75QOGcLmLBZ78W
E7i76M1NyU7Urdj40RsSDiRjiEOOJJglplnnTaad5OAeYdgWioB+CBUPC2R96rKl
XwrHxraZvhwQJDqy2M++r0kZNMRoBOYjPfDcsw/qy0142UkxayAHudYkqXJemsF5
26W1mtuDfMJ4VKLenhkd/pxbKy51zgQLQfvF8IvDOCY7XHgl8K0NVkxipjp7uB+c
Lo84kUGIHGZ9IQBDXNBQ76DTfwEnMgznVPhPkAyc/HCYxsv0P/bwvzR50ixzURJe
1NM6jiJe7X9445YWwQ5jjtEVQwcl6y2Q02AdERiBZ8XEsezhZGNDJvyK4lRW7FoV
dCpZ/fciwjD/IAW/77FwwusB0fxs1byd/H1kZ8WGJKEflUSWe/lbiaWH1h64DBWm
2hWi8cNAQ7YZQIm4RTZ1ug2Qr4YZ/Ydi8lgf5A2OVNxAwYJer5buuS0ZT7CzLbjC
LDZuIy5PzO0VDW7Cxo0vIwzRZNIS+iFT/aQE6ZfBDlk4ad1WG1/fgDWSkZLVk/It
dSugR9TknDKRqTfRwttBRdChKMiKpK16pPa8QxrnP3EpegPYfkHX3sRXMBsgtpCn
nwkgMB3DjHzRWM7ACGRK6T16JAR8QaV1ZDSy3kjY0Ow5mCgf5slMA7w79RDGLiD9
iQaIN2YMelkRnphv8dnO99zslVaxtjHB3TYi/h+q2ER5tkAlbL4GSDUBCk6VLfWy
EE+Od+brBxr+n7gIoWHNQ31JDpOxskxjZ3gBvDZXulQKf2THgvJ1T+roPmWyARAP
XocIhhjA0qilpFi94E6/TM+XZ83HCQD4U72Sc/+jy34AF7PXkLpDpWSeFDJINBbo
rxKSVoxBVY8LYDMQiBM9U0bAPRH3yubIhfJmBKo03VVslYXnEfy4UkPqfGbnyB+b
8mNdRQNURr+knIoWvLT8NYcP88u/MxiaFUU1OE5T1K2Bo9HkeYkscCvo+817kSAM
wJsDhkKuRDTq0qUGAYIX1EJqczjsLEoSdSnYYwsEDYVuaMmQc66aCH+e/kuSgBY6
1Llk6LwhfuUgWiqMtbOA7PPAXRXMIHG8tOp9hK1OKpb3gxKVFe8zpyxoeEWERIjc
fBMYMxcAKu99ry7W8q+1LvuRArHXppHoqNnBgcpjpz5zpmR9PkhYAWRBsTaL53mv
14qxtz9Xsi8dM9Gz7ObfEUM5M3e2+x4UTAOPb2/Q3iH1V+OBHzbzp/KUvPWYAIpM
k69zIpQmsCMRGLS8sNseLlk7HLVFJXSGO0Ot0YDc5/tunBNpCcMOWIElCT2Edkin
5mgFw80STJ47xJYXkl1eO3GMWzt/ClMk5iKWstDtfcQ5I77lf6cnztVVF0AQum5W
TS3efknJpLgdHvaWjvODi2hJ+yxZUafM7smSgJ/us8ID818XcuScZP5WRrlVJXxV
d5eQwcbicivNNMG5juqSZXFXXq+VyMzBk0jd9tArxu+shWJC0+iyM5ZwbUOXpzHG
wfA74fGMQ3Uf6dkaqt2Wv0pg6jGcJvgOpu7eXspwgCFYxzaUMocQatmMe6ZvwgqS
f5f/95DL1ymYsCjn7chWYYzuYDyDWpXdVEUGRySlRtZms78B10OvBDcoERsUzrIN
2wT923X/8rBD8jHvG/fbgTeWA9Odqryrx22j6ZgpFfgACr7j33aV8qqWYuzqzcOe
KlZKm5+VtS61UVuq2C7i1t6sUQ+2D/Z4y3IWgXOU4N/dvBCc0zHwtvAvjrY74HUc
PVf6Ztt84JMew3BuLJI/WRFNyw4IMpshFpg+fz9DxiHaW7dgq6IK/4pxwuHQCDw7
PZ5eAAFpkTBPacdA57F4mPsRhxOXB80j9YEtNUul7qfKjZxLPAg34ugNGuyz0eig
PkWgqiUPclPXmhRBwe7kOqVt7a714Qh0WpbscbilT94ryKwV4a19ArNezQYIAlpu
CWiITkauN3+bJCECCPTaHbXgv8p+BHojBUsxTosGfKMgUWGu8+QJ6FK/iKaJb1A+
7nF3WR8comT6wMwQvexGPRwmzJlL2wtfBGqXEiBRycSdauDc/nHhS3+DVmr+/wmD
3pzvlbWQh4UyN0nSo7X3CxZQaFhJPMN2aIVNj0sdRLTmFWrCBu6XAr1IWOrf++6g
nqzUI6iwmCuntyZ2ArzoXU10SKGPZcxsr5SdU3+Nbz66oSVcconATIm+Z0hQsWMg
+fjOgwC0VMBn/kcKkqMzSakjSoVEQY647cqZbMOTn/JaK+CmOB7lpZ9gLNd/fGoH
3uyDDR8lWz8T3hFP0l6ejbSrLaveWbElhkhCog5K85CxQmkjG7B0fXm/zkPnB8mh
uDz7NXQyP3sILzauOTc5CAiUQDa1ZyygvvcnUHjjmwX396jDyuov8AktCLMcOgQi
EUCtpDlr7zvZ6P7bjvkcwLlrA78yqT3R7yg2ZR7TmZZ1uyum+TQej2VyaGgFrPqB
D9Ee0WFGeMvZ/2bM+YLDTptEhfSu/BBqwxBur1/yxHXZMF/BLfHrIN5JORI+fRP7
HRofxh9FqmC1LaV0iN0Mgx35haCrortUX9HsGrRvyNF81eDvDQn4doG3fdGeU/1d
gMvxJo98yruOnwJOIa6JX7xYPuBFdIjEJnry7HfpNhBH2InDoiqnx+QGbUwnKEeI
f49K9g1oqFthLbYs3Qs1IQCKJPpw93l8BzKjbbsKLlAVKKvFAnrLilgvSTj6jWKl
QpIewSkuw203ZvHz6P9TqonOP6sw2cOK66ABPXedTMne2Y72hKU6On0wwID3TZcs
q2N3NeZg/7ccRRSs0MEclQcTAR+tcNw+aa702dqb26d1uKa+NnIHDuIN36CkRKMJ
JpvXG1Zy+hNrgDTy0Y2qyDu8QHpeoIgiYxIMI5MEXviDd8FgzErrP0A+9+b0MlM9
hReq6ZLvIVewIkf3OANMzhsdaV6ReTGX1fQe39bY8HGQCzAgW+F2pH1HhEn+GyFH
r3tziwgXfhMKBgsVj2kBYIyv/bwMRlivEgxfHiOKEqwsP7s8egblRjzqkdMaFeUd
3fNo8RXRwZdsvGw9EQQNb7Wvqaz7sOLo7Jue1dSpxinl3tCmhH+E88iru6G8q2dG
GNLLf8V1D0PrKXIMa485NWkpS8OnOavNSXcKjNwsPRRD5Sbyz6Zolm0T3QLMiQxf
pi3hoTMfHCXnLFSaXDHUlwGthSPptDPJD3HstwzBqWjKk3+YiOZ4WQEIlWACQTX8
8im0eLfrPo2AiE5CoTiBwq9e9SG0o8bGxPdJwRd5whjJzsIsrLoF8ccC65WDumN/
5O+E+PCZbkCTLjj76OpifGnIaF7B1D8V3oSdw8uD4JnUABb6jemV5XgEacQW78bh
rzg9myAsVFt0h5Fib/dXDaVqw9naVI7lTXlY+DPb1wE8OSC4f6VTUrb2ou5XhNZ3
hisXSJ/fcNBOuI1tlgCrd45CiCtjvI5hOnC5fAvuA7OP3Qn4e29MrAqkpZmnb+Ki
8wkB8tml+69kDMZc3ttpvw5n6Z/V1cynfhFi7m6IyA3l5MhvmRuezimfNsuY8B8x
BG5pzGtOXEmSx+v8JNJX8IjZKUhW6zBvlNkzuWjx91i8viv0MpwronIa5vp6kS0P
yb75+fhcF3Ulytf0bDLhbRwKjXXJTKEBNoTCv/2dqWvIDtPbC6gPV/BaTs7eUG7J
SRen/lLliR/HOjYr5uXKDtuMBjEiU/z0z2pNebA19XCWZGPHzj4Rp2uQ+V559+VD
GIeZAkMImJD0Mln82raP2V3tfixL3qhrYirBJYG361XrXHXLh9pbRB1D5rVXVo6U
ckb+5Dhy71G5yAsK1Ry6Fwbl8uVoMJiN78EWHo+i0CQ9SGyJNTPc2VgnqzOBftUQ
kT6GBSGvlZwY5L0xX1bvx1MwcXlpV2aftxYLVbtlKF5hG1pfOqMMcInxyzYR4eca
OviA2ZvAN1RbQ7mGduZaeldvCuyuQP+mZcK7ce/PHMKJiMH45NQs0dulDnqCBOjh
9nBNF8Wgj4zhXVF/vT/GeW9L3bZRpbepkrG4kh6/+Hj43Y1grDpZpahsL7N/pZei
PnpklHF0nDHwo0CBNYHi7L2vuOri+moky6bKNNVOE9FdyWapbGOD3U0Rnt0p7aDz
9s8qXOKpxGiYLpKF09l/8UlQ9Gc6wBi7NZ7Lr1va52luxrLhAooCo+W6jadXOSY3
KVbs4W9Goz1rzC/Vv0KP7k8QqbYE8XPAm11YRdGbAI4hVEyxI23PQYSZUzwgXvdB
qrK6KyybnkAgV3rfdQFrLoRwsUkuXxBUkmjRujXzhK1ngIEtsfRvskBGBMOgkm5e
iWhfQo4ucBFhPykFhoWsEuqZvBIio93lt9tYOoksjCym5YfGk4H0HlyMER8mTUhi
WDqKPKXjB5ZoBHgibssOmmqOmy7FUUZxEklp9YvS+DaTN+/Nnjv+4/DYnlgpygRF
hr4aInJTHgibK4CLx+z1PizjlJfF0ngqSC/TgypgOOvUyMA8NG45/ZRTnI2yBryG
sBDx1RtqKL8McE7ZOZ4PPUAaP77dyh/zay1Hf5M0+McucWCylBPZ1HpwYB7IJD6H
L4FHfVWs0SiHaeb65rcVE1jaGoABHADAFiLoFyiVLdIEkYF8gYDtD08DIfEuTiYk
k0NmdmyDK9UVhWH00WfLBUCA8OGxnIoVuvnTlEiEBIiwsOx067pCUUZqRrtI/JgQ
wAjLcsKJgWFn3MzHTmL2w+qMbYsncHELiXEGfaLXN42o0wBhsu6mlm/7BtKFNTI5
Su4JPdvlORXTqhQ+39IKl7PB5HMXY0qccFgab2WYOumSzudnvxc9CuwrTheGgofm
4G98WaSQoFoRcVydMWhDMUl1s6j8SUEFygyOy8rj7HMok5EEXQSjHjFhw0nZOJ+K
GG0ktANRLD/p6uShNdv3vOt43YwD1ScwzMkLHrjxPi+BsomuKna89YJQ5TvqNT2d
k5SGTp6m3rlJnXaAlO8cFM6ZnnvU+ptKEy49cWvmmdi+yry8oGz+Y0/eTVP4s6nK
sFCqlONrVsRmt+3G5uJlluPq9rmku443MIO1oPVdCyEhMwkUwZ++NkGqxdicxoon
aYcMybZcqNgEHiPVq5RDu6QxyOM7czojnwceeOVAdhK2hJl1AAnGsD2+8XssELL6
1sQ52+CnOvYyRf3Y3RaGwA9OcQzbXoMtuVbFFTk8ujGLnsmWP2h6/FstWOvF9OdQ
N5l6BZvuvdxEgSiT8GNMekPAQ5MyZJy2mdXLqxuKo54NfZg1gsv6hBeb5k4HgcrP
Un/tUAkAU/zF+5v4T7Icda6VVw+0XCAUK24oOppOInUbKD9edNG60hoOCBwWpxN/
Om5TxhwOzBNiCh7iGvVhdqOGRKXOgQKsmRuxbWQrXVC4ZG/NOJ/YNzzx70zDZj/u
I9UZtj+dXzEVP8taXzzWw8gJPkNpjwjPXV9e+FjfeKpCnVzIm7bS9oWz4iwpUwrg
ISEPswUdW4JxjKpWrxbqbg+rWjwYGpfyAeNtsGY+6PiF7F6IobuEjKreI+v8N7L9
1hleprbkCeSjcKi0ZSnAn2UowOvtLOuCKY3Nx5M7zmt0FCNwl2mu1sPpAl7jo8vZ
Bzp8vpBcitv0xgiGzDzXqXzS1DtnFimBVH7pTpWuCNYKtYJosFlCBndAF9iI3BMz
4okOKAy1oQRhUVxq+zzpNjP+Kt+fyravc1yCHLGlWxA5FDEu41ms4DZr0jRhnJOY
tNtTWvUiBy4dgnfZp+Gyzb2t+UHkr3OI0l0ursf5KNoifNPEoZaouCFWc9qC4jb8
eBNsOIs2NfLJrBTB5Z9jHqAf2sqpPzZBjTWKPOyqNC7EOdhHT9kWoGtHYWPwZ5aL
D4vrJFI1U3QhZ/unZ0VPJTGeA5xXads9YXyGYTjWOG4aNOjqYlvkRSkVaMQ98U19
4sDGe9fZ+eys7CFy21FPNEh329pupsIuZJwz6340EukC2Pvp/GA9MmQcAmuCPZA8
NDde/pRZC2F71ECkGIcDtgZHZVxCkcLXGPkMRyhfWI3Wo/5wgYfWPehQpxctOrNT
27FNUrxecaAl5jsNe1MgEUTMRFHWztZRfN5UWItKdTfXjPrTUx3ptNEqhN/w1PIO
SnPAKWrzKUef8GSPxTGVHHgiyXuTlVmUr1PxPHdyAs/fRNTWdFrypjkIDmNA7IMl
KRV5N3iJOAoM/LflYheHRtYoato7ODlsLc4YmUGq87U3xHOlcp7JIz3aFGg48hC8
o9sQ7isamin9RxYkosMQMA9cTg0CHlf6jP0LGsfq4vWlAyYD0pZgDYo3OOHnf3Fw
0lar8VPQNeeCIzR1wUtaI36y6dk8/dJum9XF8pNWjVsVPkvSIcQldVu+7hKq4TcJ
ylnhSg+Bf/TiU/H+5QH6VHg1jPBv2Gt3Q3aCvtFN+ZNgBg21O+hWSqocgM1p5THZ
VHC1ijDCCDoI4XTfZqQPL5xz9TJWtThTRB2eAcbJGHRIYNlxuU3DiPY5/967n3Ss
jA1iphitvJ3BMSlvobxijOm4P2DR9M/qICOtiEqsWP1llWsBsOiH8q3OIqWUodmb
9fjFocaklILorPpbIJ2rpMrNE3K4z+ashCm+7vQyDpmfIVpn0rOGD22MPJ9OKaf+
m1kkQyflqT7B4zEtPVajEMoiq5eWTHje/Y31rcfTnz8u2VrxQXnlzp8jfnbf8uvp
h5opUQ+RQQ9saZtmb8YDmaQP2E0nPNGlfgq+Dzuh3g596YgL2BK1DvThfing1M/Y
r/+NfInp+1c21mZ1+LN4/K6A8xxDGpqWeOBYYlcwPc9Zh5/7hchwJoIKDTsWq9JG
B8pqNtLCUx8FogXCHJferIVPUrTB7u2NaTeOniNZI+4BSlX7r0A6E90IOpJEwUaT
pmZneRDhhbU3i8MH8yZxW6jDqR/PA+sIv3DokXO3GVPAG23NDt0nh85daW2NVPoy
vTwq81Wn3Wpk5qIHSyaoNdWuP1vsk87LWK4XYA02oTfg9ZuBToa1gsiIdjR+GAhR
0eykU7i4Ynhywp0Q7J4yuN2e+V47KkXqR7sQ3SuUDGrkJ3y22Tl66PHVZNIby8rd
kNuEZ8yBLus07EvThDaRuUtIliKDPWn/BPhrX5Q2FRxEkELdgjunO0TRuDbxRnaE
xI+eYco4dKeRa2EbpczKMQlQ25jujm0pfUp4jhLxeHaKtKJIn7bC3tBatWqL6V6G
a2JJBq1bO9yzQC64rsBubHcTZXRWND0Xvn+4ptksg41ifN61P8fHz93CV755YxSr
O0pXD8uG5CeXO8BSlqzrHNa0pPQtCzx0laCzvo9wzU33eVpjN4A4BXpQWnYyFAgL
1vJ0sVhjvhcIl1jA6SqO9ySKMHm6wWWIu79Rik4ReEyYyWM0H94rHebKZ3W+jPbf
psLMGPUjt2QCohznrE4IiFxz7YLwbsGfAfZz4547giGMC9ft3csJATvxMP5mJ3WM
VA1ATNjkuOQyR0sYDSFPxl9b+c7m894efwIcPHDhWzWzPRjG87Ylu3hxrWeRIhL0
eX2vzxIpmN6Eg4wq3AjTc/juvfF0zR6eAxg6t6C50ial2Z0xPzkHqj/jBUrQmISA
cdEfeW6L43O9EAtcHGL4ELBOAjhue0ezeV7ivHWHF+Xr7J75RYXYHY/zemVYj1NF
y/T1sa20wUpkjv9MBcLCaA5vM6k8h0wxXivJQXo2Plrq5wd8VZOtDWGnfOT9ydfL
tAve24W3jgXLguWZBxyqzBfNUY+Z7nbRaf0bOjWvCda/kjeWc9HRpw89g9++gsE2
iKjIUyr/OvSwFVVIcs6QGWckSfevsQsm1/wql9KSPrKNIPhIjnPs2FVhdIltHda5
jjxeG2iiBSUrvdSjwEwNU3wBbo+VKHaTEORdMCgeZMfPwOLJd/P4kWxL6ZQE2ren
YoEYUmQk/l+DXYFJSSdmovBAitMAV8VojLVnhAA6OzA46P9bdQ8KQHkf+cDJc60O
g5JqUGaG3GB8yjwyixLUsCaoLrebrKmadEjyzS6CyF9OV6/NjY5AP/CG5X6sCQyA
e+GjPixsm8way4CPvDYzDhOWDsNisIQTpdjNgRmqICk1zNsreHaXxLWA+BGw9NDY
gM5SPcya23r9iTk+tRYvMVHAJIykK7lNG0yFwbwOmdra1bXaYNJHA3sst+sCfKdQ
mYLPTF/qRVqwHoqi9DW/k2vgEVRwaKdWyqxpBQcwstu2/aNdOYvk5h8xSENDGFOL
tfTEXjGh5+190kdACyhadJb/I0IRR4U7AtjSYLkUCDb9/g4U7BmBbUUdyT1nnOA9
b1o9ow99ZpQvQaKMHwiGFKNGebnbWVSEUw8prX384Ea02HoS86YiaLhWepFr3vSv
i5w37p5w+6trfY4Loi3RDg7lbGqoLPIt5BxGqzpr14h2qJpejBt36orrFTwjC/yA
B8AO6Xfw5pQZ5IeA5B6MJxkgJfjs7FEEIo1hhY6cnq+cuBUKM2ide3+vZ7LGlmgv
mEaozMdSF2RdHG6A5qifIDtybzzo2nAzNAMQQ18NxaklfUVx123vOlP+fRBN99k6
CX6CcNCjDfU8UaJjD5AA9DYe6RkifCsmZhNqgqEQQC96g/BfQ4IM8jt/KsvfZvQb
QrqLJU7udtM2g4FTQS2tOCiuH8q6ASNqv1zWMZ4YmMjrtgTRKQs2lshmofomj0gE
84Wy0QfPWoRy/uHQaHO3kKumbuaf0xXIUGF5Q8ehDue7/jbFMkAnvWP0/AtCWXqw
UKY7ENq8HyCWf5dQEo+ekovpcbXPyf1bBCUlzkJr0XWoq2/tOzGVqM2YjB9ZspsW
+CDpjck6SnxLiwkpL+usmgn3f7Zpy67EzABPeooyklAgsCmt8fbblqW8VHbTvigO
srWJM+e1/tOASUvnxCA2zRchduKe6RIBsiEzcJF1qOovnVVRfG08/84J85n3jASK
chPCiLVTrkHRK7qs0C+oHT3oxe+s/Oxryrt27Y2iMR4uLbQHrCL4uGfCtGooBIoA
lFt/TvsXUg1fIsN4lmny3LewE6kwdMa9FvpZ0pJX4ew+dSozq72NTJ6tZ0n+qJuB
n2/yzUP5EGBECtMbeFRbqciD1b+IlBKCLsHde/hSpwqZvh9z3G+PoJvZV6/9O5vC
B3dvmtywDocAcaqlk4Z8y3YdLeGmaGdd/okQBM/3+dei+m42N01FEsDNX16Lq/nH
c7NTEf1ot57okX63C+Nl9L76OJUwlt22MHyRZvzzTllcOpvr2ZIvPAUjEP8cHChz
WF/z9ZSURBPt9e/J9Cp+N643trE7eviNrL4ajs/2xVLTtZFs0PeglO/aPGL5STiO
l45djbe/5zMdtO1OcEVGLJSx77E0OV3d+zbwaykmpA769Fk+Y5OOYmHvNt+TKMtM
Pka3U462GDmY/3pmzzxnuCWgu1Rhd6Tg0zDbWBKsYaxDTSQP/xWOWW5o5pKEPq3b
hMNuvV4+ir2+nmefNCKgm31eDndnYOEFc+0GCGBVWpvyPjRDrAMf9Anh7VCZq52J
AYTGl7OuMOhYEMBQeYD/p70lbtCh1iK2WZBBC0GqjBtnoyQZ3c1eo4BhnJAI1RpT
/I+59r5eQkgFGULWKFb1K8Al0KaXER+Z+oyfVqgokalO4cUT84+4EMxYTLI58yPO
UxSar16ih1vs/cXS2O8sg2u185IldZZLeByY19zRH0lH3FVKYgy70h/sWdxecQvn
7qwpRvdU5hzYSy1mUVSdgthnaA9y8kv0s2Ic2C8R0Qdi8xQJ/kCPDfoawFmva5RE
mjLJs0k8zTZwu+oRwOVNPvDrZwcCHXeCd68PBqXaB9ybyYV4s57DO41pSAJz4bhW
1AX4raKvOV/Kj2gmikhsmN5iW8oDCq5nA9vSfs6+e7gPRKt9SuBsJ+FZbA9TkWDR
K8+zL4aVGaVGK6QoPOd/BOm/Y95x0WPzsMj1KH5p821vj7A1q+kEkXwotfiQCPiX
PTenCqLP9F6aSVFlMlD+6a28D+2EAlM1nRfxgHsLMC2brtu71zs/Z+INlwke3ASF
Yeo5FJ2NLlDZWN0hL/wtUqAb58s+QoykAwEFbO7Y6zFo8zZL227Jj3EJBAzR3gJ8
8o+xD6FDBuKk6OLSFLnLWmRjiwy7Rso1lnFvHg17t/TOA1LSHTMNZd44VS5ShJG1
Ra5YIKoAJ2/OfEPoIAr5jwSBjMiIBvgawfPU5UxNAhjsmwu5z+1nB3RxglN2hRxe
QPwYRqchge3nmDOkn1xbMY/L2+O0wCtsfBIPDbUT0l6r760cVWT9WKEbARPv3Jx7
4SBRv6rT8QFtrGMCpoWP/mzu3Eili3R2o1fEdWuP6a2OTl5fkQuQcK2H8fF5FDfX
BmY3BhqYzwX3+X6OwcRBU7mVBPBpzZ0+BvrEY9xjBdkjkn87KVXjEA+SbT4K9xiU
g0LqVJOPXM3PL4zsPj/9iuPae7HyfLTys96tg16Yb2GaMPDOnWAq4HAZWXD19B1d
1z4naQi2s8qaynpWe1BIMGnDntWE4UciDNaNj1fQg+zJIDwKeYsnfTySCePrlGkE
gZ4IPw8IZI6VRqCkttYMARAIqXi9IIbt2bQKiFBZrp+Ok4BTF0bgfxKRO+PlRb3E
ehxuvJY9mH9puSQugBhCFkyQxrB/DVPez7v7mCyVzvdhTq4Ry7IUj32HFrhZ863X
Dsd3EREMMKEGe1cwLbVABmzB/uGZhkkR7dBg2a5YqBvxrADoOdA2prY9O7qlX2kX
ZuUV2Q5JbzE6gfozjUWtJ0A9axsZExfZG7yg9lahtziFilknZEyCPnQ+G0UzclK6
KcWS93+QxAdFN7Swr2jddoHyc7SzaYWBjYQr63xflAaeuVoZ9Xk+rdXvAkb35MNG
Zl/pnI5pBC5WeBDe9KQ52EgiTiSKR+DhzTb4XBF9vf6WxaEJdrNlQCXJy1S05d7H
m2exmIhYWDDVkXNoxxzaimAVbPLgMunFveZrWOam+uFcc29TbfAKaCOBMJZ8bLwf
BljWbz0ZEFQOvWIZX6BdKJ9u+tVCHmd4DP8b11soDl4r2WTvYcPmBMQBi3tZAMC/
2TBKurywWxJOpS7Df/mYkZCgDc8ejwk5E066U77C9PL7zqtkmsPhEXBhzSKHgB+o
9nVc7Eu+qY+BnwyJK8toJ7pIxJxuCvzGL+vrKb2KUF/ww8RdqoRqC5bWpygPj7Wm
XMy1QU9w4qweFO8JvWnicUh3MlwQxzgS1hk+Fh/OuyDUXxiW7ytqaYiVJ5JkLv0M
x+Q+/lYc1s3d9INj+p7saB+/RTuEWR3hMbeDs8U1FD37t+/vnH0dxqJDmCy1ipSC
SKX9KC3qML6CvphEZjU/+mORTSVe7sN7HqIC8ykD3929wPbVNpZ2Wee9HKYuQecR
w4dMb+8WITqBHBOKLmyYTI5R9oVI/TdR6+wjwQoT3KkNh87pzAwethVKb2tt2f3m
15lBUq0Fj+hMZTPZB7U8M3THLt/RZ6Fs1g/+aI33E5qzNZkjwPX0SVI2QuEeA8Vk
MuOiBHoXQcovBrBER01E3S8tGT7zteGebRdTa9Nb/aG44waluoHSRBOggj5yQMHn
X5coav7QcLqNIrEYATgh009mUhSOkQQk9HgghvZb27grfDznfVe6qye7J76dG2PZ
h6eAagRXbirjWpi7Vh5x6NVmEJTlXm5/aijG01P3IkAtGmzeyMrx688A/MUXwpvV
ILcvZJmRS79k+8scss9KEzHJWWeaG3c/wDZknkR3Ng7qx/2aCxDUji14PWoedY7L
TWDURnwb6oyHN+eMuigZoCK7ePMfN/xTVWq8wrmDEN/U4c+OWPId8dT3R28pMOW0
afFVOoBT217NuZ7wnTmP9svRu31VQN9hDQY7jV5JAWl+r0rP0Zi/2TH6GEE5RSuJ
6yuB4wKORQdsgyqVT6hh7Zdu+he7Q5J/7hcPtnkEGTGle6hDLiZCdUjR3SsS74tQ
WiTCpU6s4s3xKliK5bjMU/eFlblmXKuof+lpxw/HqOJOv5MyYqvjtHtrKEyhNian
TrkSyHoUetCBHdmx4pJ3pStwF+J7RYzFpV9bKxTYSuLADasdeKhvAK0UpDoR/wWJ
l3NxUFcXfGUvOe+UrPB0GYXpjCKyXckME6NRAf8PHMaJu0YmmQAJgQT/bEiTBQ9v
OKuff7yR2liJrBx2ThBsq3t0RjQP4fkheVhzlfllyh9l7Mvq0lhFpgMvvrxe/H9i
pMCgPopB2VUOr+0016ii+S2hw8NwsuvTlQPuX34UNc5PQSBhpQdyr2bho8HPRfqI
9FwmCmxXn1Gc3LNut3bSbncXg79NuMXgFzQQMwrk6JAoecZKZMcHfg3WpZ2u+9aB
EtnmlrJiZG+YEOm9Nv+Gk0Hy2p7DhYlUbRDKzkiaCEA3xEhcV2tSodT3pWco/Mde
hbFDFxh62hJwD+Kv/87BF8ivdEHCrM7kNBhomO3Gi1GZ/uBo2ZZM7UBYuFqHiqEX
tIkIJlt5oE/VFcK7ZNw1Dj1x+2FsfzzlI8C+aDBINIeJwFYxMZKlqd4BVzCVk72r
wwFdn94FDxIJsvBT+LVHDg5JboMIFXWdRclNM/IZKwDFzUkzSvQ9bxlKjYLFsmFH
Ig8t2BXirmADpqUs2XmRJiQyVNxZnRfTxS9k0K2BoA6Y1DXE+KqJ9g5cNfp8/lFv
Neka2N3s6BPx+P39E0N0iXHBs2oMswRf9yWR2vl4M59Nwf5dQKaA0jTUNm1uuetH
8cva2j/EuGtjEAtUOGgpkJ1HAJFe+eqXcezvJOZ6fsstXq/PjOeyPlWMorUktKEn
2E+VEiYH0tsU/ArKAwbvxwCtRVBXXryHPtMMSQvJEagzSYXg0gpd92KghuAj6WNE
eJpeoaM8emdRiaKDruqrbbAl3uP8nbEDbqcfgRQX1kaZGDoJl4mBkaT/zGVbiTk3
dSoTX7q9U11JGGAGmtz13I/OWgVjhbchiQuk+ruNjy8b5L+jjdFhAvDioAJWOOBY
4ExLEWJTM0rpLEZuWPKkGwZugV5sFBovF+a4v9T4QY15ohIuj6mBTJF6v+pT0s/p
pYDa9f8mx4jk6Kq2yc2TLKPQjpcIzixX3s9u+wGgwGiatWvgM+VbW+jDRA8UDz0Q
+LbNBcvjSD85No/vtSe9IFTEij5kcFDOG9r7WCsYkFXDaqgvsersIhixw8Asdh+1
yfA8WktLcnA20HWfkLxQQNDZTR+aITHBjREsivf37gmJkL1f+d6Iv1vr82aWcyRt
b3PSkro6oh0Jd0T9kus1gs9OYtUxSE3QhZlMi4t+ePD1Hnnk54Lk2oDi1I/L6XQE
qpNGdmu+yQhh2DKvxRSzXdBafFHSXrcsgKW1t983ujltaB2BZLdN5swSQ7EF9Mjy
PHrlaFLHl214dgmvkdxTIcMe7kpjLxBCq+u0CdHSGw4ROqOPeTudJMhWx1r5s3sJ
i1oC5Nb/yAdpm37Fq9oOGVLwFbTeWL+r0sjbB0ORYAyOHcLZ4G6eyLQowAEEO6u2
xXh5x6Q96vo/Ytydy1UvcUNoqKjl/Sm4kH4KLhc6IhiGhZCojZcPMB7lP5a9vx6K
e7USVpwVu1WfCBY+h9fMY67XlstCHYiLDWmW7tIOzRUv/raE7/kNxhUYp5dgLKF3
hhXEB8ggu9MsNF4qdKROcNVQvHsGni/c5LeUALEWJlWHfh+Dmkp6jjPxIdbjyfy5
5cpDqD0+O1mCFiNH5b2wA6Wbns5MVXn98WtQ8Dg5Gma1762Nm6mkHJa9BPlF/Mx/
2dPumhXLMmQKJ5eECJqi1F9HhuSvhHSW10+76iCkvf3QuDijZXSVe0lk4MYZf0sO
gu8RkLZjAfYU8SWe6226H1h5/zGOCD5Jc64Ql4hxstYXTzwIGPcx94YO+zQhNQfi
UNffdVeupPObNQj7BI6GoG6Q045HRQurmXBhaS0jEu3KW0mOryA8woXeFDdarShb
wG0i+/Dz1Vayzb22vNTZSnjK3jf7fud7AY3kxzzo/rOQ1FIhobX+F/L1eWqdZCG1
G1Imp97R33Im0caaUaSL0D1CQDp+8F6zZO9Ek28VJn4f54JTE9HOLAqx6XCxQcW7
FO6/8DgO7dgTW8BbslhKPbYBtMEaQLEZwb+daHqtfhNR2UUZB3xU4Q9CWrvwE++l
46+X3JjCim/7Ja06fyTzS9QAPzgFW18kAzRmB6ITVGYCMQsqXq0GsuEeWAzxwo6D
FF8CqXaC767gH5mrdCNZYw+U53nbBnCWMnTjkvcoU8gUIXMi01atfcUvNZUlqjub
sEpV83CiAC40qjvNLQN3n7PYbLFje3rZhuQ0GT5+91qdnUq0xZS+0sbRMU3RgnF2
cXcnSaJDOJQ9T0A71yDBAUpxbuw9F4JoRZ8USBOFbtd4hWSwRIWe1FCIv3aw5z3+
gkibjHsokKqSNfZA7HYh6Dc9HqoU/9Ov6IBV4PaKeHJP4Z/70yoeNfzjTDpmas2R
+HqVxunlTkL/auusvWuLHFnrghXRT13jHGTGwT0tEuidkOqsqydC6BFUWiBYK8yW
usYrz29Oo/B/QQmfLcKbCWaidksk+MU4gjrSoJAhMAfCMqp4qduDygd1nwxWcvIQ
I5+IO1EeCzzq+I65d7HdEue4HujLetz5mXS3lLiRCNKULx7mNTRbfQKyT9wTS0w3
EKFoUiAPan/oLnEsJhN3OR6sXtkynvNY8C6WqrlzYr/Q/1ctqt6yR4h092kt6TVp
kVq61tYiNVVqo6I6Itf4utWZtEXHPwYpyxtDF9AOMPrfLG1mZZKUk5Gbm5uzxpOb
7kJGitE7hVIjKcsGwtvxXK5X4z+WKsdGRyLM7LKeZFMQI72QyrmOnY8k7japG9yb
yvfSzfW67EQ6V3K5oaQgjVgkmhqJNgYndhGgw7pwHRmy9wLFGo33JcFoKCh2WViU
rXimhvk1k8OyLEak86kkhSFvktfwhlE9/SFc1tn7QVWFatVPKQcCdtuALPStmAZp
YiGDTUT3Zlm8zTHNkfL63/TGYuZejc3QmpzWbU9ir+hIXcqbBWCAhjqDy5qJ7fye
rAc1nc064EaMrTahbqlGIEpAWdHQjNt6bedtz4CdcABYxOUATKzOXL75+XcJiGU/
5wUBvLIsH2XelCZVZ/AU8janj7956ItfC/hTsg5cjE/Mc+Nimswm8HkifWAVQo9s
pEttx0BCcbIvfklmGSVTPFmn0QMP6DoCNC4Hhde5e1cLb38W1YGK5CFUH/GwTyjb
QJoBzac4eC6/X7Lm3zRNxqN7vrEWFnrHGsYaZIFnyDx5ZS9iPhfM94+uFSbCoF9z
OZgr5LsffX0fFiYZgiJVdZhsfYCZUzksyPQxcoucRNB4Vt0aLVNC773zSrpkgKkT
ckrS7RSRxXKtz+7tdBluq8aUFTKXt9+DTK4Pv2l9Q1bMZLM/gaywATeGd0Xd9rr8
zMsd7mCPVxkKDltAv2fOHucXudXCgcn9MiYj0A5LFnsV2TMhzaZc8+yAwncJ+RHr
5OXvfVLUycXequTmIBLuHkZhNE7VCbBeZxWVogYB+57kBU9a2z1/QB5Af8RKT0nG
GN/ZbQP4L56UgropeD7TVLEU/UavjfF7oIaSr1du5yQZNRdzNOFcnpDpHgUXmQU0
HHvt5NZT3wgXD2Y6s+lUfT/hbhTqWg+8ectU6ewih+H/dz8UO83tMF1toVqXpg8X
otR0GBbPiLNS1bAleDqQe3+oaEG1P4OP+f37ZrdtwZkiHirtzyvXXYEBi7t7UrUV
LPL4ixdxz0i7qtyiJtE7j1uD/44iUUe4C0A+yHeAB5+IJh0pVN/CcmXrN7KIK3At
qIH1ZPdpl9ojGmHvZr9c1NnW4/vJloTe3RlOsszSrfGT2Jt4o0l+EoNLvaStazha
/oir9syb6R8X+msNmqTDPrX3GtFhGKCHHL8a9tRxOCZPDZPkNwwvWbGSRCBVxabd
8R/prPZrn84gx9ny3kmNGPv9hsCA7KTFZ+qpXhLVr92X2fLpUixpWLCTAumr40vJ
eUODCA4C9FCHaz96IcoeD6myyiqP1jSSoFKexxYZQNATOb3s1ffo9BqJbcMzG3iR
QYcSbNP4v7bAU+Pk6bnFqp3kh2WjgjhkJPF7TxDWokh/x9N012We8n0D1wCNkTwL
rmsB6ravLRJTMMmsKYb+yEqr1+g/kE6Ui7mla4prEY+fluaqghTYcp9ps9F3kkHA
0IgcN1RI5G6qZ+fTnYMXcg1771vYfoBV0kTgNH4lltq5IIyd6GGk6uhdd9iAoCWz
vfPOhPU6QIVYATtjMr8HnVaZbnSDpR1DeZ2g1TprvkJ0no2NR97F3YluAWgRq+xK
cfAdXTV0ZoIqTMFGVBKKX8yWIQ7VPWUr+qiP5nDg9ULd5i30KMXh7BmC0ioJ26U7
L1cevc1VFiZXKFXjDnhk36QNFLtLPLlPH51ATsGgOouX2k0ZNuANy1EOdaaADN/x
gS+zLVaztebWQea3GlX3HyEQWUXtvZkIzJGowghcQhNyAnaz20yauzkWgpKPBVgo
YKwFkkxtKHxMoDvGt2GuL0YigBM10bS6n1p1Eeje/QwmuxSfLMgRerkv53N47lQZ
mVQCr6PtURf+EA2cBiEyb41DWby5HR3In89UqRI7tiZKMsWm/NO7CKdQpXWnVxQp
mKbBO3nx3stJlrQElHgU2m+1XtGVxjEQzJIasIxZFSEpXXANCnnULCGDN7k2+OMH
ujRoA3YHeHeU7DHXfNiQLranY0wBG4VpBCLZWmyutZCo8DbLt1Tyfj9emLQvYlmT
VOEuSo5mTlMPbv0TJVsLTUkA0RdZGHVkht9iZfPglbrrasTU9SCQHgU65sK/xT/j
sFkFeo98P7wwdggdI6SXmIWC8BXySmLfylvwVupAxTrfLHKWknmrAZtHvoTuIHuS
/etXLcrHsHzu/Y23+cVtNRx+aqo0lb7hinSCAx+7iOrP/C3GcY0HhqsaZWpCdJ/F
jFMHHsFj1VRKGy2v0CWa5xWBiYKjsepHfXP1za7EdVoDoqQhLfxXD4JlUUN5+hCG
iCJHNQdz6qt65mrS5w0HQBtxdJCqG1FIBgEpWgnvBxVbeRS447GGNFolZpZjS+xS
9IUYqy4ac0fpHsddT40SP3J9G+vVgJg/zoG1HT54b+WQ+W63X5f9wBBWLUazgENQ
4V6USXBUHxv/bAz2/dESTphI6Fn6lXoRu1vSYG/YQ15/PKx37fse7TslhW5YABt1
k04Ybf0pMfbA2I2unY7OL5t5oeZYXxqcKSEODqbzNXj1J2jxAPeLabRe4vrBnKZj
tf9gcIMXm/FB3CM3HWCk6RnyyFDwly7qUfjaVbdMwpTNF62XijkjOjZDGLLaxquo
7ypat/3aGZVR0uRdzyhDZTrTcxNZ76rmu2wCIA/ChefmkwlS9d4v8SZk53V8p+1q
staauP2vh+WOS+KghfISk77TLgNebs5/WPggUQcCMz59CPkcAGjt34uBcxhwnoP6
SAKoWxaVdbtYbjXuYC7DcKOe8RoiteWEKI2SDbk/Vk1oLnTLcOMnbhXhCSQoAywg
ba1e7OfIt1+qja5Z/Eq37aQPHv5DF+BxsvflLFSIVu+A8OS5EU+gkd/6ds9C4CXI
vFcH7vUu1VUJ3oaN+x0nPARQKePRaIc1zCK4ps9VXJP4nsN7RFu/K3vjaul+jMwc
KsDthG88mWBfM6kQfjLInkpTQqqPZ53cshPV6xbd4UdsVIZZi5Zdv5oWciTXyjOT
/vVTZ+Za1kKkkqkELii41HD31PY55wIOPiR2E9WMgZOSQcUO7mV11L7Qe3Vgj5KD
bb3Rbu3Pr8xCiH7o8+EmnCcUWrjyLcwHl7SOk3LYC8GhXflvqT4VbKZ6OktDKVy3
mAe0Gr1WswzIproRel8kKEnr7zgfJI1Hmh/Ej7C0MDSn7p0KVdSLIFSNn0aB2i2X
jHkMOwx7LnngQHcBac+R7wkF1mLi6e2IwKlZVjGePHRLgu5/Mh2J/YLp81Whxscy
+EgyUqjMmqo8zYOr/HrnXVmCiahXSfTenHjpjHkoW4iiqd4N7MXJWepWqg2yJ4wE
hroL6vbJVSHZrgnnFrYfO9kltl9vpaPkCrr9BwdDb5r0inr5AeF/XNO4Q9CRVtVp
SxvT4GIAiDxjOITc8CIoZ13BgiexvwbntFdEmvi2Vgn8FkbCMljD2LLzUQtg8pKP
C3Kbw0KS2LVKK2S7BvygSMFjs7DJ5t6JIDiGdub/fynEMY8bGmMJp6FqN0ydgZba
YKfo/4Mx5QndjaPnrYLtKlzNynDi+uLuaUJohShcM7L1fSaEPxZoY+HnbHM/WXBg
Wzvox6EnLJIIr7A1s6WpqMWgw5uYpS8us+VpBHnhfVutQvwAhVU8n5cg5S279fFm
naZMFeUMivlJ4RrWYKWv+l51bzYO0jAdAnH/PPEjhgD8IHX+giyaMM8B6dR35cA5
1W6HcRMYTeBeK/hf3t9PjaL9Df8Ib/ZN6y7dLEKB09kvgB87eNkQlCBrYAYyAOgX
cQnqcaJjE0Q/24706c52MSIHtuNg7B/5pafmE+JvZntOP7XlOul2MtVkS2MRXhbi
EIYXxRUn3ghl/d6UvoVTIWj4rXwBTPsqS+XJRx3xiigWZC7K2Ty1ksyyBOwNyjH8
FHd3lMUCnqUWQFVL90ZDQlyWBavqRDvYoQkGAsQgkLsiKu36RpqSOyFjUSR/B8sJ
FwZct9ho2mZ3W+glwSz+hl/4wByLXFeuKLnoI8IUBaZUhcnF2+TaaZUlzyBSYuoO
KOVQ85skasrhnVjEgpiHkJNP2yA+vsCjX1uqyPpbCglnZ7J6m5jgj2/JU3G2dAKc
gNEF67X1vAgyGNrW8pt4qOn5pDUdA+rMr/UxydeyLT1yWh2bUWcG7T5Gu2a98g6t
wYjuM79GwkmYyYmtEFLH912XYVlH7Ubo7M5rbb9UoWc8+RibEA/Q7s0ut/h4lLfj
ukBc0VeGp/CDuM1bC8CqpFP/KSLSBY8l0wUcLaBApfxi2EIFWO9FOtLdC7nm/33i
ufubMnTtFSy5Wx8tq9ut3buT3/awLoawvr0NTPaedNf30goP+YO9ZTrf0tiHCT7b
t7e0r9dY/XjqM3RDn9YWcv4d+zkKQD7PG3+mmjPAO7phK9V3u591GqPHmKd2Vq0s
nrtYRmck4liVch1jhZlZOeghKwikwXQcqm5iDF3qX3pN9lmD2XdSSxkROhl59e80
OcJb/WWsa6waFKo/TwkoOleUotyksqubVJ8GQIXqRaQjdCqk8tOhUKSblZv9H8TT
1h1+DUuMchKwwQhaHO8asPH5mDBA4MO9bc0fcHfNq+be71PgmpTXM/d+qoERpnub
VhtjH5ua0RVUylDYRxmHrykPuXrg7K7SxMauDRZq1O01l6CsKRbKLxw8LSSL7ZS8
dybQt3YusqmzeF8x0ayNl2mGiwWj2hhl9+QcPtNzZmhyJfNo176O+ROPvOfTBmVu
WwsaSK5Kpp9lGUXCxe3PIWE3xZyv6MsHgK3+RBTlnu2X8fgvPdQVRG72uZnuASuC
+dhU7Trnx2oW4JmTvXdFtfq0Ppfeoq+V2IBB5W2QKChINBCBvvTd/kvHrEBeL09C
aKbOR6vFJsTjx/GicGRudR99jgsqzsqMZe0XybzLXwx0FLxRAuWJmVz4Ul9Wc+Ua
q+c/F8uUecMT1NLIiAxK0UE+qAZIX0KT1gY4R/gxA3lNsIlVk61VX9xaiarlsTZM
85KVE7FwOvQXXtaEJ5QnPnGLmnOcblwUqrOS90A2GN4KLawFgbCJrdEiSY6hAjHX
i4yT+XF4BCZ4RNcYG+XAgVt5cPLBMnjFlFdzWrrJe5FJrImrFPMCJ2W9kXHiNbM3
EGty7JUuk9oEzV6qe5OJ7MVzLfJYzNKE3C/VbrTFEA5N324/czn8v1irzJiFxF2H
rjkj+Yw2gaQUbV45knSqVSOUbt4NojhVb6KGj5OVZfPWSkxsa7bfpeMnrQuPiHfs
g1jm294MvwIEg4HmrCGdafTD5Isx9ILID0SBlb0U20l9astceHMhqrXMQiF1Fshl
twVxzXk4garH3DM7H90h6EX/qkuiH0dwRZN4KvP0YsTbM0BKyB+Cc/loL/qENoic
LRqnumbrNDEUG4nof1nLvX+1/Z0Zg3ERDBuPa6VxEgGPj/mi0128K5pOJ/zWn78b
nToH3lLj8L4kC6nfC0a8FbowBRUNI7xJ4S0IxTQfj6yG369dzc8gA3VMTl6YtfiH
9NfKLAiklmRPxplJ7C+iaa2aDlxzN4j/A1Ictz1UMzNVduA3IqGkJ6728JfIpeL9
8x3AWr3VPvkHPw9fhJc4wAuR20pq9SZ+Etm/vUI941FJ3kDq3jz8Mn+Gs48qZkGL
s9tsy9+2WjWKnUUNbpvZ1jJZz/f7Uc7EBwmFkofTTC6es1rwQllhjhxRpF2Vbz9f
1PM8Q9oZTsn6smcIQSJ6K/XFQ9TCqyZEGje9OiZjp7zYB2cUr5BTmRvpZsxUTH9Q
nbQ4l0e/Suzw1qQ77nKPpLnfnvba8S/voW6zgYltsPvy1IK3xbX9Qw8UEBCpn9qn
VQu4Z/6BEQxn7RBZ9fI2qll0iFfS2nEAlXpeBnuEStYIHpC49Ig1YR8rvGtcoaNj
Md6rKEEqcjVKinHTsGWrNzd5oVMd+5OSudV09EO1JUPs/dpIS5iC/sSb+x8x8HDF
cekn45PyTrQh43Ud7ZscOvyEz/zlGwxF8xk5JLKOzreJr3O8M0s9PKJ7Vs2ayFBC
KrYBW0bqlT6WGsPhmqOLwfE5PKwEXMVgABNhUka662Txq/0TQjUyhyblM7E06z8B
DawxgmObcfQEe5o2QJH24B/9QS8dLCAGIuDaCfMbrq4jCWWBT27YOrcZ545hRFCw
22AepweXrhZIavKtiKTPMfU24ZTJCflnxPLvW4nZ8lwoXnRktJfY8YXDE29rUs7c
EHgNi5LMbmVM4ui74F+jomnnBpG1x/cfLuFiCSOSB0akhUZ98iU7taMG3hp7N3fB
jTOPdqD3mhUeJ7BqYQm+glG3lc0pJge4lIRhHndXedkpLq+AQvFchkXNjhcExOgL
gxvry37qhr5+TSBVxvSBc2Vt6n/hB5d43hUxIGvuInEMOCqECiF/OwheeZtNHFoB
lP5Phbu5AaQ1d4bZ7M+WX7bzmZ6EScO022ouXuzNyw/lcfQ1QNYvL/+s5V+LdKHP
n1CarVY5QNjtTDO1UGPWJA90izXQpNutqSnXgUYCugmiOmQ+WesCZ6mKe36VbWPC
DNobtroUssp/sU3CDkPN4cqKkW4gdnLNTWP+AcB2KPuR7OxPwpZF5yb0VHWm/JZ3
sQguq5yklCUW/KsEjYO/38d6Niv1LRe3Fu/5tUK6BQ0/Oz24ck3jgxWvjvU2dTao
CH6MLLBG7JGQkQSYFIF4PLLtF7hhN4NGDwqjQsnLLOMyGawrg3ixM91J/FQ72jKq
VE3v+h/UHZgndOyfXFgjbWWkVWhe+82bKhkuSheWpPxGz3SO5Ct5YFfaxa2m6U+V
nB1tSnpNf1MNiuUVzTC5tJOUGzDupPwZCOAeEWoZSoH7J9IBkaGZcNCFerdDRDIO
GKYpO2UYZzf4qVDLa3rHCJdW5WcsrePO+t+hg9VLaD8D9at+RzR3PwIVWg+DKqFn
GWdTFgpSOBVTZrnyxUtcr6UCfy+LZahuwzsZMAIf7J7EGe2oIdF6j8CEtW0rE8E7
zmDDabMdxh4vspUz+i891kbt8QVMjU/8yvYsX6BSNLDGuFTQbVNUVL125UiNq81C
aKuhhwAsmrW58XHYlte+JWV/zIB++b2kjmy7MEkwMSdU476eUBBDTpAyvmHNuzfM
ApimiW0+GvJaNTy0GNdSbUxGz59OSxy5reQjePSv9OCtpGSpXACWhNlM3U2nq5Hi
ZW7/T9Q3Cw7ocwkKAfjrJBhVrct/2s2xqkwZ28/7piegigydR0OiFn+QinzagV5s
YtjlwtzlZ14iZQQzMkDCtuDkOEqZfi9DPL1tXLuZr5CK4s5pD9RPbicgH3vXXz8C
FL5ZvMGtJYJYVjzKUz5DDFi22o30GJE0wjNHiQNlr5Xp8o5CKmE9yedbSGI4u52X
+ONLZ5u7RyL5UGwzUs3bGOOf6ZC0mSAHHqiaoh9Jc5ghYRsro1lXAtq6VHpcYKVi
vF6s2IkrA7t4ULgsfHpd/Ypw271F7OAuEzQ3lnj//YFHcB3jv0D6Bm9o9+wpLoBV
RdoqIWvHCIKp3NJZuC7IvaiMAy/wz88WQ0YyFC67fLKuFicEzQ+f43dalazT5Tbh
Iw+A6myAHZO3MY0WALsRdh71YbC78sBLzTJRmG+B07obUOwjZC+WICyJ0qw13jKi
zqRe1EX5OZRzM1rxIXi9jipaPPxDAf/dsChJD1vM0nUa6SeCQu7c3dul1C7YXdBe
NOwehya/Oynttl6RavXv1YsCugZANqhN0voVjTjwTvNTsYMjJHQL1KwvvGjgEHS7
vWaZiNyJnwxeBxiGsmZB0Urs8jkOvaKcCmW3FP0TlLTXHvqRGTF6W2FpFiPolRVx
DMgxCTnCmtvF3M6qqFxGb1grNlSCPUahhVfxrUP6U2dH0a/qa9xHPCXzTQ5WEX+i
CuOG7lOpVKvnKrye434VcqV53FucBEP8QWv2bPSHkTAI564SysQlHN5Gx5G6cFLR
kaG+W+i8KexOTweR9u4LP8j4cxNHP5qx0+KCwd/Y6FY8kw1gb5x+VowUu97QwTiJ
vsO/uqSuKAIe4D/f8FEwVKGou9Kz5fMxq7ko6Sum5aI4olgCOQU8OCjanq1vqQVI
DNDj69vD0h07qikbC3YZXSYbKCkFr6F+o6oYy0d+cuDo8Tji8ut5qwCRZp62bDUF
OV5idbnPad9zVHpb0gF1AQ4zrR+GNeqaEhHO3zcsbNxggmeiGQ5TElVAQmamO7G5
tkcfb2a93kcNO/gWpF2ZWJV8svxBP54Sv9vBSDhfzoErGxW78UOGIJgVDvIvulME
2g4eWhWKeTzHrDQNfdZXEuFer8JbQspr6HcqjLdrNPbwhmEPU01tI9pJFqUmcMRS
qlNy3TLiRCHZ54avC2OePj69ibB2pb7wJLyr+TVXZTK9IpGSz08FmDDtSizhRClV
Yqkb7o94E09W1/MGX4pfnZiLHa6vqdMeVnFKP1BN72zB0ANr8MJfYBqraA0TFERf
folmCPu+TRxXdQY8BIHpjyDA/LirKa/VnzIswW5TEViNsiiwojRLPa6mniExZ2uY
J6gUnUIkXyLq4Kn5dkAaVJeM4zPf82CAMOxDIJGdrre+mtp7hWRWtDJzIj1o6lb2
wGRWYtoeZlf9vECLkJvN+rkc9U/PBV0IY2GW24O/HX10iRv03rBLWqHw2xg0CvDA
LxzBzm9vo4aSz1JKMI2uFK3iOG5nGnIp9FrZZoFt6KZm95qJCZe35e8BpQvURvQ8
QNY/gfhqxiv7UZS3WUL558uYz8HnJNWJaZoVI8xnJKg160sbg6mvXGBehItHIbQF
h9UlrbCPMmFMHJGiKMl71ysAKbSztj3ImilwBLmSoqCB2mDZ9r9tlhFVVMzBBxwA
/Tl3uTEHVJEH7GySEtzmpoCUNpO8FgYJn1WKWt+ozMEhZzW/TxLFuqQDIQqw5pye
/MRRRKCnC6bo1qB8XZ2GNf1PODcuFF70n2kLr+S+ZphjXvrmhK2Uwq7lIqugJ6uP
VtAfRqKlxRq1/abzpKbyQQ1BLkT+J7gxh/gKaVk7IAFVLmnyRahxsAanRDkBccjB
G0r9X4F8yWB2q5J/1vYzh2OgT78QbqHjmdVJGXBRVNuhtRFT/2QxtJjS57u2JaDN
p9WrRUebNiPWfZYPUacAsTDDe/yOj1iv3FxDeqB3pxjGcbXPxGg8oklsoeA4WBA7
dG4xJFG7lxzLQwqetnO7K4AGcaqJXL3hHxr0fyiR3Gd/7ft7v9atsjES50233Udz
ZptqT1+N2EmRyWcuqcgrWORa8snvo83B4Wpy9Z+dwUAE3E6uqDVpzWfO9BeToZmg
Hly0h+CG18McC9MgZs+VRaB/eiq4dGFgYyaXTba8iL034IbakyW1A0MWzRZJDAf4
TCneErESQeMc4X/6PN6Zy4zH+7/YWxk65kYqDhmDfRw53mwLKVk9+C3SyGOhly7k
PlmH+gWam76od4ENh4/Si8WR6yndnEKA55U254lBFvLCI5jRGMHKsYGTctKTO0le
gB7kgrYo7u3T67yGeXj+XsNva+Mn6pUEGpl482ds0ZUfEKYI8gTetgUl+GGst8+T
PFWx573iIDqq4/OE2pGL0XDcIJZg3m25HLpvqw1sx2sBJaoZeudX1/jbU39bRWGY
Q5zvNHQe356wI5/5RUWl8R9ZbbMgLqLiTnAJg4ImJuij/ppkJazk0LDlN5aciQF7
lMoHuGF8wXnvGJNfrACSnC7mliT9AckemUv6RF5HSnnbbwr3YA9kOrqHZOy7/G+x
q3wiDzgCFgg+o562HhRZI/Fkg4kAgnuxYfvstxWeNR1NjPMK6bLklI07TSIIkkm1
mZGCzI3STjwC0/0kT/SmFkZdOZ1f84nYVipubmxHWW7As5FgLbbu4ty6WNCDxExH
SF8Ow2bvFLf10Gb8PnQlSW1QEUOzxRMB7UwJSR3vwIAP0x5iSPn5Y6icf/6s9j8y
q1ZrSvaXGK+u7cZXigW0KO9YOUVGfgkqWG2fg8IK+qmqjRrzAzNxS6I/sBgjRNUg
ccw1CvNbRJilMPwryZuMRerm0W+TqUfdbt1Cm6M0lpwSZ3hep9/HF5gjclPNoZzc
Gxej4vmdoFPilmrHwejeI86VgfZIOP/SZLh8dvxV1djnAeDIy6CqPMC2f7Z6BPHJ
Gx/22iOnfRt9EH69lb3srF2i9r0ONroUcu781RuIPYyzp+H9dxpRJ+KdHvBIlSz+
EBIvEyIlVT+qKP8vrFUpAfP9k+d7f94RU3AncMss/3+UxyEB1Akq1WtZvkFj28wH
DgSZQ6VekvUYOM2Z0Ilem6wVJF/AaXCCdLNgZE74qmT+Bvumg0X43MMTChgLXaNn
kuJL1Zu28Uw1KSmvc0aL6wYgZOMi1QWCZ0c7d4l2c7Te8ZwUn0j/jL6dKqMz3Tk9
31FdYzpm9Y5MOzQ7rVV5oGUnQl1m29s7kWnor1FP5vnkmcIpaJN5QIU5QxN9pxSb
xUFgDKJRLQ7/Rrl1bUKwLTrx+eI0XCS01tlkWiBtYtML/4eb5P2S2lZZUBsZRJU9
oOX66blm9xkL8Orj41aA/dUNJpzL1dijUUowpDiaw8Bq91duWTHNLyXnyCPCcFtu
SeHU1YOseuIrmRG2b8PW+44EEOMdF7jLOXyClbOWLxh0LN9r9VO2gL6RQi0RCBnS
euOrDNLUliHa6fmQbnmp0agTTflGuyLfEf4aW7ERFNN5n5OFbzN8U9CA2DXU0puP
rQnQAir/txNvVologGAPGZdMTNP7D7qhyujSBjpYtsiEBMn2gWZiHM2nkyz4R84B
uDMh+tR2oqkhPjjCPow+K7Zt3p52DxmSrdS9mBJKGDe9G3/kkWaQ0GoIXkjdU7rT
MxQIDEsja4h6pMvLDCMTsRcXWVCMzNcAsbPUE+NTwpO20qBN2p6I4Dq3TaWhdi3A
4pH5Gjxm14H0f7zg6bE1OBZJbMcCwVTdGAOC/a0D7qrG42473BnwmR0Sp3RgyhDB
/xJDYCtaxOqE1TZyLy9GP9ffe4RYfFLGuOEBxMxKuMxvzIMsUVh8tJgSk++BxYzY
FMQlosVU+i6M8Z8EZmjBDJThsPDDotHYjvoWnHuurvWkmL5OjWQeiY8hUuOmNjXj
6vUVh/54DTQa+Kh1LFxoRmP3nENcf0rc2SuQTy4IuijQviAD65UgupmnSqE+z11F
NQ1FYd5ewkWwIPZy0AMM4AHpj8yQFFDrhTamH+JS1dkKTrAXHa0/tk7V98t7rAsC
TX7vKQ3wPZk5+L8Q54XwiW7a4k7RwF7rryYg77hLRvWukD4AhJ0N2k6jWlqsnZMF
9taLLtfb8Rgvg6LHH01E0ExQ2MsldPrw0BFapHWdvvi8F9bSF/zZJkGPtaJ/Twah
487ln4AFgv4jXBnQFDIVlEfoi1wfHAsbEzNdY0VUY/zn9+8dYddQbkpLeFtunZLQ
2AKomtYsLu2cKWNPS6clPsHuawfoPxkktUL2hVpta0hvBqy+MfhZzFUXuBenRFdQ
bGMuF9izVlhgntYIUTOKocznkHz9x6dIQsd++qc/IeAumpGx/3FfU3rKNC7l5Y8c
xCvuOvcsEgQRIk3OQ1OcwN1lAvAabSOJnNTApLccLRo3WrPpupGhlEh1RKhwVoLJ
GIVISt+g7I6ddvPD1iESYoPf9R84F6SDx6TX9THl2uTStn4R4R8BdANeo+znbmSk
WlJ6Jr4+LsCte96UCSdCM+4v/7piM6L7rzAJcx1WIPrzrBuE0qx5R1O4ANQqRT4D
TbLWsgGsoMQGdaMCVZ1yHhYX2s2RNL0wqSbFdJu4n1rNISjqfXcUoH7nxKBQ0YJr
ZiuO7db+852KAJXUtNXCe19gmTGuNdZTAC713omZ+bqa0I30OlwKRw9oXr6ygEe8
QdC/0lhE2cNf8I63qMa8JZwcscy8/A4ghQlbGRhf+fs3iPaNNvDUEW2rYpiXiVYu
DVHiTOKg1rr3eNAGZQRETV3hzq8sUFNRTBzRRNo2Nvj82x+OVJ6E7GXZtKlavLLc
XCypRFGj3A+DXooGf8WmcOQhECvq0Z39XnRbSUUkR8IUqN/Ce+M+3dS27alNFRlq
eD7Nsrj6FTXRdkl2rMspi1yn9H5u2HNAIipvJqbFeIx0Rum3Fe+1VT7zKC84d7XI
RHjUjPuUnEblk+/1uXgDIFvD9S9aJLIPj3iDF1YuxjIIFgyF2Hh8C9WGKi6q2ITr
0WUvS2Dh5jS+zAvUrP/ktHQGK8ClPIiKsm7uppGbzqa650hs+swoN1H5AXm9SKy0
xbMqLiCtONscWZ41oLx57pEtd9MHxXZLYilC8y1VoiQITZmC0eHvJtTwh/vqG7hT
MyYCRFyTN2myK0MuY5wih765KxgDUWHQYepXuoY+/nf6mErkNjZNH3She2Qi1UXp
HtVKaPgpKtK6P3/kMrivhvz1/8VaMfWlnpp8PWhop+8f12VcEibj7wXfMx0NlFKE
w2lRripQniUIr3+aKO402W9IlynAZIg/nAFi5nj2GtcHp4cRQMWnep+2KL8bslk3
qp7Y+z8CUDHlAB2whyFkCGObPMVUBDURptfHThdEU8Fr28UA/rWfHTf+kIkBsqLf
bY+pmj5aMlCk97u2Ro54IImejQeZuWJDHTwXUQfd3BEkjUQdSVX1lLivPSKwn2kS
qDRUMLweV4+VekZSk0JPFyswdEHRuwO8jG50GMZQjfYb1/mkbcWVgWZeD5Eh//54
HaGjMqsQOuaKCbFVaT07eg1qUVq2ACTkh88H8uQLZYqEvOoR73rRnFzl7FX5JTuO
6ah0ODjsEVWxV0f6jSSaW6VMDclr4wcVJPFzeWoFd6cbzbU2/P16V688WF0g2Udc
8gtG5rCbaScO0AOoK3OF2XLuHqau7lvY0GuRXGvhMZjFS22zM5q7JHMnwxO/4Tlb
EI9WkTQ1+fzXxZAHCdBDu354fMrP+AeplyyPQ1OKUIOUTuLUKudIxDh+U2L9Aqac
KnETVknDOD09sPyI8ZoJaomMsbkkhsKL8wBjFp0j/ZVo+ZtGXOon1StF8RfBIZfU
S2f34wCuUtDt1REpcE7p0RbtP/2/Q0Js1KR5a7aGrVoUhBxWIuznZiRoAiCBfn4o
ribv32WkKhrcB205oF2MCVYP3XJolTEhNOFohzYp+Uz8v9JJfTz76kvrpRnEj0Vi
DMxuEvqasXP9E3ouJDfk6LPnPsuA+t0H++Oim2f866AvjsLIwVAxzGMNySTk2E5s
ETLJtcKg7k/FkYip/ionXbzRtc9/9K1ulUkiYn0PGQYdA1WJaVNp5qN++YCD+mUM
ZKbeU4WZ1ip+6KEgM11nJsgA9zRks4K6okN0K8JtkNg1L7fEeDnwjhyP6KKf0Co4
JaSOs/0iqOCjB7Kgzapbu7f/90tJCJ0g1jXtwkYCdXrm5RIKY/MIN7y2ryc53Wiv
bJpQFdCQtsazAsUKqYVIc5OPB8jmKxSkAl4u4+NuSbUthV1/1dOBDl5KFdRdiLQN
EJ2XQPC1m2DzkUNhFCBH3qNpFUbQs6KYOf1duJtbtthSGEWGh+Yeljov30Nrw14G
TDUON6X3WOd6THXqPWJH05zdQh7ZELOReSorAwHBEs5kvgFivI10DGRojY+SOuGV
T3ISxef1DYxmLJuEqPVoULhACRcIbyBfTp709X0ClqkBqNeNNCQzgMFbfcHBKUPI
wcMwEZ5SfZCeV7TCn7kV/GC7KiKqch8NkiDtif5qjnEcd/rKC8vdzyzQQ1EVEdCr
Y/OOJXWzbX2XDYKvsnuXla50APtlPfSeA6rM0Fx4Uel6zJuSxgAyOxzCWVrVGtGz
lS4njy4dHZQfvaj8NjNdCqbbdzmUxPaVF9J+5Nk9X/JPf3UBvWF5oiQbYNakkqPg
wb3WjcqFhHaCWAA2MmiVr9xYQo5qxS8cXfaC2aY7/8HoPT4Ynz5LAp9qY+erJKAx
TwlB0moIdumAFIktqADsDYbusvjilLwrI6S/7b3+Ok/0+uQX0qyrt9PBal+qsrMM
+jYenHKpNnBtUcWktz4rwepWzDeYGIxugRnBt2WHXqhodpV+/Rw9L3gJOLpOUf2Y
yXPh4pxb6g+oHWOdv+jesIHIHZ5WEM1QhKQKiCT2dwtJnRdQlKFAXOjWDr09oj2Z
qPYF7hFtRYa5AVpByDsFh8OaMveCuM8oMzOCzhxdGQkxSUCV/HLIJ4KnB/JIbbjf
/6Fbu1P06EAGUSb4gTuJxCGhh9woi7mJodRYqyWGyQn0z7XYB4OdnkksSBGl8XYp
rFzUhAS+46gfrumggJNbvSVfQRDpwZVSjWUIL9aYOt40AC8Fh7l83utXOJjwwFbX
k1N+51NrQumzaYOgkkOfhk0ArTtXQMwdHFPAT2PgzEeBlt65LlXP4wowY7OOgZSR
ACGY5MojQMEVThkP/Q5tNp549uMLd2mUm2IntYMAH95pCuwWEgdSI1vVS713A0p8
H82IPOU0cJj65UWR18PA8du9g0hptPp0pBmiUPMWt2GWn0DjlJ3a6ACRU+NJYH30
t/7Yda/aMkgNEUkZmD93hTViPmMS4UucqS9E5iet4TGrkumb2oQsOEmkNwPvP4nv
ZRcixfiHE9m18VbJauRrMsJbax/SgqIPdvl3UW9UBecQ43Qajb0UQ7KQhcehGc+4
TZQ3SQPca+hgL8AiWTCV2gM/seMacukgFEiujJF02IMcTwmBXcTqBCFc7SxhtNXM
pg8uQvkrF0WXIs8AmUAQV/7nz1HyhW339Y9d9hDzQS3v7u34UTH+zqHdmkTULbY6
/E6LKMo2uAhX/7eriolw15eOr1B3ccuNHM+1+gtsVD5QLEBuhMbyfDUSSrQgycxU
TntnybVeqKwzT0VFRGqNVb0FldEd+AODo1/UPmRAgZuCBvGYySY6QSrWKUMgkUcM
SefZ5CG/3IfHxL7wOzvkC1DhYDs+nFUi02zltp8hA9QxhDo1qKvGzysEadP4TowZ
qakovMZ4RM+3v9rOPEnsZGIkqO5t8IKZidXJnKQWSGSOW5dV1WdPh8Wm8oS12OOk
nCJIbyrHc5tdFqd2KSMDfEO8q1nBkhzU2LCOzwvoquDlI87SLtqU4QGxPaNIB11j
9udRjVHPa3rJWjQPsCZ4nCbnyitF1iAyHwCTekF/RQj/XjTKXoC19WpECaPCFEha
OhGDR6JT8HykIaQ/otUKWojAR13AG9AB+cGpZS5apAEeRogrckHydLX3yr/vvtW7
0bCSV4b1X9lckW92XMe9QcGPgF8CmhPwIMY0kzypjekuxUtl6pXXo86DhMbt0H6/
mxhWyRefqSZjOTVaBbttsRS+sBK5/WnF5b+cA8/uG4z4laDK2Qvg1BcsXWnc5tpB
K4MBgrkwt3MQzT+0h4nlqLKTDFeoerXFMOpFqh1WcYTFeCDB+v2IZ65wuus39NqE
Kqf1E2/w6sHIyi6L5dV0KWzfsWM464fOomxTDDuGKAhYtzgKw5CoW6h1r74Y6heh
3ZMAg4GLpsIalDjvtYc2lTIHekfW5Qd8f8duj2mKDlUjyzCydusVxYPjjVUxAT6i
qYkxjEsd1r+5KuJTW7RpFiWkzgjf/scNnZYh9OesEm3hdpEr8JJAG/bcYPtgkxQZ
u85gApms/vkBvfxOHPKikSjxT/uowga7cKwcJ9MdRa1mcCaf9xZAGaQSqb4CuCUC
7E6K9BZxaF1c2lBEEZyngMxz5F/maQjta0GjfDc3akq9T4Jn5Xmh8SwzVOMoZan8
2y4N/fgR4b/oghzcofas9phhAq7tH5kZ0FAWwAgnrP3EGprQSjjY6zhKJclZLLGB
IAYcwEcjcGMRTDB+Sy0njW2ZeaPrIVxttSP4loSu6OiAdjRcCntPTB88xjRJg8JK
bieTXAtiQEA/lIlSDGd69G69+ZtfgHL5HOnLFE9v6qDoOBrTrZZKpLAhmQjRbhPP
0jz1tf6uBjzE29mRm7HNFc7Qyf8UemhYwN19OnUPl+YkFln2i3Uak12CrJOQD+Zx
JWKvYPlhS79sZoUetMps97KqIbabHyCX1Uai2PEd7mlwl8heDyhFTOyeQnbiT0jm
7uQl6MJ3cQ9hAPjTaNjeP46XButDwxRuAnV4QP0LL0XsSpmiw8fTNw1p4m/EJPaD
rDEdqkvZTyFru/l3HC7CCQazs+OELW2L9JIOAhmjU0AJDgDXxb6EomsnKc1JLfk/
ADSAmRBoOWl/ZELX3rv298zXxTMb5gkdAaWWKjail3sYhUVIEb9BwJ29IN+WH6Lw
VhiYPgyL7L23ZfNJ1e9xGQH5XsDpimiTHfXufeKJGWGYpwrmYGEVlthz6Rrxe3p8
KgBj2nCZCzmVh2+VhQYWnRtKIMoUp2EdLPpkjzPrAxcmgYIZmuXlOVLHLq5IwyEb
UUB3Rdo4SSLyzIN+cB5w0OiQbSyRpP3ZU84+VdNOrCkAR9bLLuPEvB89TZ3et25J
ZB2TUsfXHLup5ugfH+vP8GEmEnc3Vde41Y1ZOYN5vLae8KCp58QQM1pua9RQbCGd
O7Uap6EAqLowHnr3m7rPBzHIujf/jCmvpweIHcWYb4qBI9DB88v8p01wW4oAMH7E
WMA0fLLSUSbJRi0/lBz1gSmBXlihSr072KsuXbJ9w0vUbPmfdarnBaSl3BLFzcQq
SuzIAzv5fCCK3Wx1PVUczITwQEPozSlGvhD1mtmQvaK5qyspcbXBVBO5PHKvXTaV
8SowlE0Kmhox4B1kqhlWxkibM/b5oKjtUPg5hAy2eHyHD0dVCS/ucK/4F0jhQ9fH
vY8xMDUwyWhT6WZtZFDPhyMZBBhrOjiYEdjJF0h9HIzdt3N1IMXaVsCWilb0sIlG
m+o6moPsZxzx3mUKQLj0MPkfbwkZX8tZIjuxl+fb/EbDZ3hqyVgR6HoYHEpCHkYW
QE7rhznnRddtxVJGV1CEdOT4igxD3T4+TndrDKtu+p9z9qQW4VQmJahYtNcOKBCN
vuZNnk9LWVQWDxC97pHMWxLu+GWddIZpzV6snhNd/S0x6K4Oc7cxQZrOjr1G/k3I
+8+ht+y7nAAuLoafWqSZ3VUe7o/0eW5MLCt89pWTpZAkEw6m4dBjkwAqiqIKlZbC
RMIBTfFIbnMZSIAiqGKOd1syTVDMgGVeFO4+hDqk1hlR816eD+880qpXy/YHDkxT
4eK5T3UYda52DdNxNo0ggBT3RCZEVnDup2PihL6uirdveXSR03qGz6cOZipiRwaf
sQzRthZrjN8/HEWH3448O/v+Yeh08KNWcctVQMTtcRxxOdRUQLzZu9LJ7qXoci6A
dJQzr0HBuGaEhQVltnZhD4VJ3TOQnGHYQuOR5jK8m2Jqn0iB3fQrlRcALqemO0VD
Cjri8op3bjVjgk+yqR2HfLlH9XyrbOlrnoD+wNG0D4LbdyHQtvjs+8wGiscXLYi9
mxYfURh95JgT9kU/pzsPmDASXb03iOhOD1LfP0MJkUe+WGts6VdQCypOh+TueZL1
fyh3zQyYRHVx/0TSTvSOq8DNFZnmwkM35QPL8hXfq31iVyCDkw9ie5PaaBQ7b6Ns
O5HcvVuFgniSfhbzTJKZMTQ6AO/zy/tU3+O56Sz+LVuIbWdr8z+SarNfuOz59Jlw
YKVIABRTSwwNXaMgjFKrxsmlOAZkVmcz6uLjfRa1I32N0xIKKFWbOhWcc91+wDtu
8ywDugEmomGtBz4tu7deCyOEXM/XeioQ5GO2sdSpPFqCiWsJACc1AAUWHAwvd2Wp
VSHh3uruTET2Lp4J4qs36CbMcYmHjuiKlR0eOQzH21huH0I2XVWK11gDdxAo3DeX
b56XbQY+DIZ6FeGmiIRDjzLFDbH5f9tW2DH9kTv4OQAKd0aDVriEaBMLFj4lYUBF
yXJfOPO79s3pO6PhH6FViv4+3bHnWDrLO0i+juNnAs57m+ZJCRy8gxXGMRRXfsef
1kHd5ZSPHye5kIxKiNeyoheJ17sp6ZB8fW7XuV+zGt2JQoeJ+hjmneDw05dtHaOT
jHtLiiy/CSwA68kzBzk4NTdJfekrvViwuwr86zbQFKJT8o8FZFF0eAiV0CInR1Gg
BI+ELJjDIoAGbzMSqSBbfc5BV6Wi02h1t4XFJ4YyljUfXzhp61CIB2DqrSwhqwGA
D3Gn8UKrFJMBKhYMw4Vf3kLM4Kv6GTYCGVMKsvxlfVCna58itqvl2Vw5P7IwqS4e
Ahc1bsdbtDCVLpKtq9aMlAqYWEFyNCkDSIoQy+ZB0imi8J+1Q9G9kRSnpq3OqfwU
2wfrvmx3n4Vq8TvQphz1cPdHG7EkC4Xp+9Uvj91VoRrI6RgacL/rDQpnUqpzTX+y
rOQqWcU9mgsLO9UByUFBrQs2MGVLLDVk6Fg02KlhHUllgRLo6qpeGzpoeNCr7A6s
icwVIKr9uZV0P6zJHf2aOl2JY/jdoVbTHztjY8Y4i0oYPcpCwam9j4PB5kXIT3Yq
Ue+CuVjrn1NMeyXpw1iU0sxv+nE9HlkzgyXyQTCf0BatYngPWXPcFyuSr2lTQjkl
BZOg2OmyGHlI2WMDpCEP7WPdCAfB5kzZ6PRVPF3N/uB10bdAiDwb7aWG5nyR0CkV
LRhoJnChIHlVhzrMcrOgrZERQBEfNVqzLvcEd8fan7G9Fz19XR8Yttr7PBvq2AZu
lV+CxqG7fcRm24Y/IMK5WNiUdYSqjbsf2YvrJZ6eQySTSDg3yODpaFTJ+CeadpYn
xDYvCA4BSGIaJl5Yqpv5hgFM22nzCSqmMrrm/jy6oW2hgucC2bbpT2t3sPMHP3Ec
OCQakBf2C/zOjnvY081SQPa4LwsNHK7UjNizP3+2ZG/hzSaW3Sqqt/l0ylkD61xL
4pyc3qBg8sKjHpGEeRsX0xdFHK7A2/ImcsV0PwshiZ71uP/WsMnWuofU9O5+/3P0
XooLWHS/Cbu2XP3fRF6EAocmzRnq7r642faK41jG5UP3I6c7FLmnRhMC3lc0I2B1
FEM5Zdl3zcIibZ3zLQaWfvq4s3tnn34V+Sk/yvfjR0Us00c75QJE3s8pEyDwvkcR
virFCafI/Bdslv7yt7i5UxQb9arq396exai0X1PMvAw/zV5A04aQXI4wKwZs+LpF
EP0sEugC6e5HXtGEfgPTGaxDZvPwGMnqyrTvVqW2qNpCmlo0790H9JQYpQ60POj5
HYbSXBeexXDhoXwwVQ6I7raB99gPJUAOLhLLfZSnzgjlYa21OZre3SF2OjO7Z6q0
7z6HYtNoL3ZTvkdhsWKhx3YhptW+kvhSwdYv4yz9x+YghISLfK9W964ONn2KKOQ9
kCKTYPT8xnt9akD4fE7HiCy6P9wEs+kVZcxTspshtlhGb8XzR6Ctr2Rw9C1FrZv0
b8oRwuJ0x7PniTjrCODExqTpkmFpG9MrVh1I/znyYjI+IaUnFviF2WWDst61qtFw
wT/daLDRPQgbwxvsve+M2G2fsWbeXBnh1XHGeZpWXuK9XruXLo2+S3E1C0L5GWO/
g0oyEo/4Ps779heJOZgD+E9RKP9mlpxBDL4c4Yy2nk7DQbj94RHrpAl2JOvNLDbx
nz08fuAS+XdxHgvCjrQAlCLJZpSzU1u1cxObObQGKf7yMvgHjfIWYj6AtWrqE06Q
7vvZBcuFLb3j+PUufywdaGf6uMi6+A8uket5UkdNq4pTIi0RYX3sJgYsFgm9ADxF
g7QTpIT23HkCNDbm3tJJQQpmTAJzef5BlD0yCfItP+6N5EGT9WoguQPc0zupuaql
HNIz64/GgTrFBUpUgmhp91FUQPLzghOkcK0rQ6jKaJ3XEquZqYXkzh8jeE0ZPzIv
lq9rwPpBVKbetuM7kdBOLMN3THNphQE7ahFS/KdRjdJsemp1ZgFdQLu/s1UfThPg
5a2CvUus8AHULCkbQZztSzQN+/jSe06f0e+q+xVeovdOx4g6Ef7TxXgE7YtXPXwO
7/j44J9ZUeq7T4aVX6uZQujsph4yu59xZz09APw83KiR/x6IIbNiIcbz6Ruw5r+g
f2IuoO0x6NeOh79cMkGMcYq4/cVD0Z0wPqiSLqfCOXYECNL9Zo4B94MUKRERudBh
KeJcrCC2zgcGIvAPkWUkoqhcJ5k8gfBrj42vxyss83F+hsCX6hgtyYhyb9WJF2/i
I6jXwdYTaJIgWmg4Wi2Vijj2dRqt8/wjK/v7wCVnwZmqMOZttVh2qM+5/LD4o8Qk
tmiryS8S2iPHiTLvi3hkpDhTucJebycnccaFp5OBhbNW8adVkOGmtWVtUjGOTkxS
IgOR9YCid4tXdZNSbCqhLLWWCQyTNRP21toKQPIt5Z/OHravUbi+y5nTvBCWgId9
Y/HBjtma0doxsgOvrUMn/zDMOGCAExzFXd0R0Pahxt0qA1AjDhVWHXdc5j4zdZnB
N7QuiCPqxQOR9GN98qSTsXDMCrYUWTZj5qeKS74Hjk13NUeh70iSEjgAQRQXY9vz
OhNsz0ZOZR+tErW6v3kgdqqltpK3n7XE51GVxo+JhGpvoaPuzpHWadqLEGAhQHS1
zIIH6QVI+TC++Tz7EZ2/tS1JMAqZNTl4aZp6qnkbpbjcMmnlauTPYnZkNF9T8seJ
sZFfYqGDKXTt3PTitbK7b6FD2AL4i1vMHAaZCph4LLDFSBSAeCJBdwJ4WlpXvDhM
ka24yVp6FaKSStEOFMzPm303IyzC1ZVbp5HJ+O9YDk4+tHKMGLsbh3U1INHKCa0+
04D1J0fERpivqBd8Q0vOLSjDmYblGRujc6i1GJUmUtsKPtj+TDaFeK2FauqVcjjS
TzdkVE9Z7VfXEc6LnnyFf5lKQQlicB51m1tg7bbxmA4QDHGG+2cxxfluKIdM7ILC
W1OlRxsZd3ee+FQjs6qBD8W8JNOTeshqUCq7PEHS4jqDQQGOBkeNPwSuY8WFdkoX
1+vUWRxAniL+LpY8XuQCEhBsppAZRH5heHO9jX2KXJB0tjAeXHyt1xDnrIbT++IO
dRdReRVQbA2U1rmyc2sHqIoNOANzZC7Ae3OV+hgZ7zU1FjJJP6/sZlXsVXItDLWy
yAAL97QkZcdq2tZ+EyiwIfWt7oi0W7Ydq4NgjxLwXsNA6TEamKp8VKQmNGrUKbxj
3G1jsCJjrgiVvWH4mYz53I6R3WMyL2Cd96wNIQ0mxGN/Mwh+eJAGe+HmGmLMd6Tk
7myKvkyHuh5mjrleBCsLMKSsupD5+lYj0nPKU4hKkwzYkvk3fycjtUC+Ls0aFS9U
lbujbAxsxdaw5is+gomf4mPpqt0s37mxDZuiDgi79SAyQzgQPXNFwMDE8VENE8QC
GzHAh2mu2Dl+LpiszKs/9K3ubWeCPrpQobj2O+/nPn2fF11uxAhV44Xa25ypbYQv
fOQJ5o7XGBLPEfQdT74JZRAzU8f+sMm6kWuCWkfGxxXEyzhQYK3S6etJU1+3QbdE
sHVqqEo/RbROL3wrj0blzEFBtJJT1LKJRcy7soGCFBrJZTYO9zNSQEJH72voclWo
UQxMm5moPOAmt8GNaxRXM80gsNE4TFkDpRofi3CdOq+NintBnMBL1vdTtbulkdfP
QXmoh8OCZCx5vlS/20CqYDZLG1XAQZUypJ7v1fmR8aJI5s3ZmAYzVy5TfxrbvwAp
fRboKHdgYhXQS3McVJsh67o+iBurnOo9iCpYBNGwF3UvAb9G/Dbpgtj2CKD2Uoyw
AiF9aikmzEp2YkaUf7sZ9vYZMsOUFAE7h9HPO/CSU4vq7hVzgqI7oriMkOqAREAd
JfD3TOtnuCccdk701OGCrsGSyp7LjmW6MrogEg+K081ygIyCv2lZYxw8QXdcmdL8
GGhLYOD3OjsK5a9eMBMZ4tZPiB8YYvBdRLPIoS+OZnLhgyGfy9bxjuji4uiOgrDn
/Z62BrvTSNylqyCGSCf2HQrLGZecefw8R8KiKL8l/R6j2kWjcnshRCLRp9pkwwbY
JKJwp25sjHc4G6SNj0fy/SJL6gREFi5oSKz6qt8mjyLqYfjU5XGBmeiGfWjhwvyz
cGoTD+QqE7d2ff1S/LCoj76E2sbgOekmMnfV3Js88lndOzk8jYwX5zSI4B6eNLl6
NouQPU1pvQr1/Pr4zsZPLqSyraEPnoOfZKALB9kEWrU1VuSQwpBqIZlK6hgStNrO
tvEwad0dLujORIgKCccccWejq2pO4LKZcp9WFo9RsTp285YreF769riFC1zP6T1w
gN/nxQeTOGqWPSavjgcLd18YFVhQb2iRPz7hEr/O0yAnNkDvb1lbJ9j8QSraOOf2
cxCIaED3nYNdp3e+EnWSoGZ5fUQU4onQIaJiHA9css1kzIdrq8tvpdQCbt0G0wWC
2shGZiBRZ7QDSgTE928zjepMd4JPDHFjxgbh6rGtimatYDWE1L/KSXsxn2u1UTUG
DQVA+HJyPFLckS7FNLHbWqMuVJN1Qx2NJLBKtsnEsREreRNLiUcx5I7ss5nIJYyd
96bGDX1qGpMFzYp//P/obkJ11+NQ8oC2/+Pkzko/GC1cbmLArWvuNwpeBvOSK2w9
O0EceJdbzDvLMBxWZYd3Bx7UXVIq9C2tYpx3VYZpkvdUIC58XNItv9Kdu0mEgkhe
XrnMi5uYRZn2rRqz8+hZwjC4kRuVcMaFvB/x6CKm3osTQbVuJU+p9+PKA+4IcNyK
ytoROC2r5qtz5AhDQ1Uee59oqKKZX23CDYwrVdAbB6Rt0ZPgr4M3Lp5dkabmE6Gk
SZqF34NKLv8v41KZEyUNz67FCGjDlHeUNY7u8DcFLUWgfHaEIB4SHggx9hFW1AvV
5W9lKifUda4NB1VXkZNA4rC/T3RcO8k+qxbH4l6w1mWs98965/ld79FJ5XTeoHDu
SC8ssmgVVmMXup/5FqVVIItcjkHkqa1H3wV1yznlly/c0D35k4crpkvCXTbERO/9
bdTQ2uXkq+y2hMEM6sWKOny7w2zQqkSYoowf5pqjfaMHR524zA3suagPGw9LMk8H
Pxt8GsRrEQrhycgpZWtndhuBHFFmnlSZdtj2UBrXgWsZd6O92fIi6QsKSBb2crwl
fioWDavj7ayiVLfyEP/87eAT/E1AaekAZdeKwGD3nYp3Y5SAwDqBMlZyNjiSDvFQ
OJDqv1v+nQZgqAzw2wNtPAEz75ahiIVQnBpd7YKgNAIJhuXAan45PHNTrEwSAJVJ
pCIrzOo4MQzoI0JSeOu5t1m97mjJcQgi/CeP0Z9WUQt+zljWyMe08UxoZ5FshBZ2
3Z6w+lu2ECVwlOhhjwF5rIIkL2Si35sa8HKth66AWFF0gwGW4Y3MdrzVg6To/WdA
Qbod7Nzxz9BPNxLrUqm5Ml2III1FBxoN5YXaLO1gPJVfV8kt/1hvqfm52vKluul5
fGCxkPMWW/M2ulhSi4oQJL+GMAuihLBwSMuaR7lI/xo5rXvVmBkUUlktr0i49EBL
UjBqh+yIKuAt0Y7V/zFEQAXi55vIgitLhSufZOGG4sg4bE/9+uWXNkhYUgWuT5/X
yFcMXjCkQiEMlrnkPXwjFjdLsHJlZXn77ilBXmioZhOEZSfxuCHVCHD/R/DglVRL
Zp8jf9jnXqQATBY3HEFxTPS5nNpHyR5k7Dw8/1pEeLZVua3hogLFrryTnNxaZ3zm
Exh5S+crSyfL0yTVVM6LMekZ5KUdEZYIiRPyWlP1NzLrHWHoz9eHCwj6sVCKte2C
cH/3yQE/FEmYr0u9uDrWOGo5qOHN8yMup6jpkpcvRTjjEkzCwXg5N4JuW3mnSBlV
wL7RgsShNGJ0zc7hLsx9hBf3DsZr5107i/L6HgRMZqzpUVs4AWH9BwRbKFYsMWHG
b8shoWcW6dfZ8T4D/o6VvQduLUWRI5Ky1/lhjAzl+Bstd/No/B4ZV1fcBuxeAa0P
pdEigQ0zMrRX3xioNIyDh629Au5B6oJq1ygXY9lgWFXV9ARZfIjjYJteqDv/XJt9
SgCtxVvWP223VlfcZZ5l4EV+kKe10/gmHlQBWwuGpWBUkdE63spLFC/3EzoXmBXq
Muqgyar4v6msoTwQd35FQK71HP3nrrru80cqD+ekE4hBD3xHKRWVIKzlN8MM9oCe
qaZVj8qnd/l8AbEbITs9ImYbyrfLXayMrCe0U4jhvp9YgQJSxOfnlGlNMcxj1F8t
U1Rwoj0WrdRLi7EAxpjtuWlpz2pBrH80RCcujfPixpJrFoxxYWB4p2cthx293q4W
Ryyq+urdrLQ/fQwXcgb6QgTYhwRbrqhknURZ47wj78gYIojmd91O/0rfppH+r2ZF
ULvoONknl4s4xXErefzqp/Ay+sVOmEoauRIT0QTpKTv3pgvf/nzQJAOSZFY/6bMn
CmWqWaZzurkPSVeaFRMso+G5VQU9CfWQjz71Cc7PL95T2o073zt3bUdXClo2gpTU
7buRoDl3V80qtmRpBf+/Pb2wrfmEpipzjNfFBcVhaVSEAeOJskmEQczlu5+eGo1c
enYiIBaksX+mMatZyEqKTMX9oZWuX3xojMAOOE4iP4iM6mHksCb194LYikYy+J/N
hYfN6hMexdfMqKTRzaPUY3rEStJh0jTEt3cLmrDURbcnzcx9iEJinx4gib1huv6n
Sky4NlI94Ff1UII5UCqbCRO+8ZZjLLOgtXMeDd2mAdf9Pf8pPtzpJZ793aEvNZq4
rZcUajwqI3uHSbCOtjOc/+zECjdgvaTxV9BHhHXMz83u0jEd2MDqDk2oCwee6OlP
ZWD93iLJEO4CNlodUK1qXqxASVw47VHe6qQloy2ydQulMXiCQOl67suMzK08wBaV
OPbaH1n3Fkxb8Ic6jNuQ3XXUXA9/9ukkrr/8X6enOlz/dFkN4FvehuW8r/Qe/OND
0Zpy5OGnWPW692grEeO3lDPhx/Oyl/0oQSwRomzm1Bz2wryzV8uYpKm30OZHbyb+
/L9UXFHJb4IAMv9Xy2LJ0jpNIIEchPOTM4A1Gz/ZmJzm9ieQF3daXmOaQnO109ib
fC05qHojUniOHdl/0qSxZhO6ybKTShyF1mzGsuWYpTCNV3lp4odgSfahDH2fB8qv
SjeooV81h6BQD6XpsQMNC4DQdY0d5LZVX3ykpssjEJ/LmvzgRA1IAyweZDT30jBN
xl+KEeR9ZwuOnTCpnHOV2QUNoCjtJwJr7UnnnjHGpRAVJiCse4+uVg35OCN6haoh
rWyCvLdmiJhI7zH0Qx8K+7t3RMOjfKtawEYzUrRicAWkOE0HI9tGH0NLdvrpYRde
PadCrvTZRN1KtTg7Y8wCQamIzU2nAs0Lq+zVQ5NzTzaS3l7FOHI/su4066rOBcNo
6/wKafdtR/jkHZEfTM2pjuYoLUtifUHMq0CjDWWH/ttstPAbaakpqt5tINZPsoiP
sjOPbHmhz1gabIswFxXb1jJBGKfQap1Dn/KcoNG7dT3n9rZ6V6k8blYr1YY+/nI+
6E4vUVu3GuImZFIwqYsxp0lujQcYvcf2JgGzDp/KmQtDF0ITyl4yGR2KCNEUq9mu
dHAxJ5CHWa1KbOydTQ5jQslP4/UcH019J8VQJGi1E3H4nurQhMslJXCZ0fGZGfFO
oSYhEIC0n9vfs2JwTgQjWkC/Q39KYFRyAOYGOnAMvwiHdzdKSk0atyQFYDyXZigI
D8Q4v6dwvEWcpOGXIzbZdG165v5J8KNVZO3dpKamgfwiYO0cI2geY7tAImKXjJmX
npmkDEd3rQzaY5FHEOAMOKeMpEOuamk4euwC2C1L8qoag9MhIosdLBZV/yu0hVFO
dNzTybMx5V4zGM83ztGT7Fc9LpqQdISIRLJWmY15+v3z7Og4GgwCNAC54OoMGkon
neE5soG4no/nRPjVhIw9iYKkgTUI2n3lc61Zht0ML8pnn587OhsXCQWADXh+9eI7
PgjGql1XpYh8Pf3bZZuyjdp8d6bVnNKoo7u1fSZOgWmvA3aK9n0Ei++fQnafySkJ
niiIDWb3HSlAxudYaemyrN9bIcwUJ2ApC6hIsr8ZWJVaoha/AmNrnaAnF3sIYfz7
11jMO0rzTEqx77oWlYseTX8cCnwyeyU4CcSRghSP5gmkxyQkv/GQjr4rBqZ8wcQi
pH0TYoBMX/0wZd45glun5TFHzuKdzJVbcHNNs4GLRZ1QckkFH+oPubbThDAi3RJU
3icyQnJFlKAnetCbzw8huWjLcRnfnTgNiTLxcXPllpo9WGjCqMTZlACb5Z3zGUNZ
yRu8J+MM+5jhXGGfKQ6p+o5RUp8n4BWPZmJr0b/W0qG+9YX4CbqHyHDSWA88C3qK
Oax8ysc5vSieA88JtXanXkq2DG8HCAmGaGdcJYpiriOd1DdLblsw92Htpq7lAwqe
jSXF14zhC/cEx2mn74kRRoZtZ66UGf5eOnumXpI43VWMO//manJ/9qmVsis7phhK
J9zWWKxDORMNXpmFYTqO4xrA29/EEU3CvmIuK44Tp3cK6mfXzzqrhnTg4UEjmgyx
MQzr5pKnWO0kxawE6o07oJ6lWlHJyNZYMA5s9HWyX1zTQUxbuXTC/XrXpZobuJTx
IQvhBKN6/43R3QV44BHcZ+cv/EmOm3YgfO8PxWzAL9ucc76KLQrkXnqB76dkn1QC
mV9VqMHgO9YRRKSvgzR2aqFhFtY+aMHM6YI7ZzR/zVugs6vTxaCgYRESFFvuwnUY
EyRzCFN3O4ca00D//5IDOh2lWbEqxcwLkO3p9d5PlO12Ys9mYy/46YxLHVSjO9M5
l3byaTQUY4u8yGnoGpcNfjwAMBMB0URPfyXXzTKqT0Fgz/Ma1pYmSlTtIArClUCG
FKDyb0rZ2YOA1VLmJ0ntKOLUjr18f2vKMK/hjkkGhhAoclI5UGCezBizCCZ0lPxZ
6U0w9kqjpYMuOoiqBSBnNiO37Xw90Rg4kYzk8z9TfNKj0XwB9ZwILm7lvsRAtKVQ
R5SAy0UEIQyZRxLzLzs5gFn6yrj+BSAK5nuz17LX95UOKWFInQt68dbyHQ2xkHqm
d3lhYThJjh2wRHTTNwWLtBWbzgMSh6xHVRlUqYw9VUIxMF/5xvCNIWU4J67NqbDG
h9BInxRJdIC5LsjxUyhv3stgL+/2YELAbQ8kh5eA7H/uXXAzaAdD6w6148ZbPa91
QPCJUf8WpqvlYRvLk2jhW+KGEqdLaD8LoUh25gH1dSdhFNddLOC/87c5VkTlfyEQ
g9ak06YyxMfBhFt98ug9dwdKQ653RumG6KYMad2e8w/09sP17qX9VclmoJwse9Sg
1mVdCoY4IcfUeESpd8chRp/DOnhwn54iLgzR81YF7SJAEtU+J1h1agIQcD5S0vw9
N/SsTQcEY9WIdvvbeHZpZ4hPQZqfDL7Gt9kAQ64bagPtjEpX5/clWWp9WxxgbQzx
/BlIJ4cln00er73zvu/3YAoMiHHj8bysEZ9FTC+OUl7+ePCayAhxGFcwDX/tMLI0
OGM/X+Kyc7XxZO95FmBqGIgNttUobcxhL3Ndoja+2xmC9m3ihCNkY/IOygWroU47
L6J7EfUPc8qGdDqRutvtPjL0DqF5KZNgPgZ0aQa2cu59w0p1ndMPzlh1/b9htLQF
gIySCjF1GEXgu0yc5c1FL6xoirPvRVx56sB9tOeotL1amgA96Q8GhpgY+A+fEDiD
9KnH2MUeNqp9EqYw85rwsBpnkbf/yeapVFWIKTLzTLy+KvcQM4YgWPwdPRXEVbND
3fuB96nGFq5Dz375RiRq1YSlw9GABm8OBWoEnhLK+A1/dHfuTSOy0EN2G835/gxE
Y5ed8KjMYsoQBDkFzwwYeK/dEno/9tlK16wKTjTP/3eePTtykXbFYCrYvtFSaVae
ThLqX1dP+Y587qPiUcgmJGr2YTDQeB/R9k2pdqZxYgdChLZDVm3mOXRz/t/mnn8M
hCGw5igZHlLlnROhC2v0vmYtMaoIsmspxsHqapggeLjrabda8O6CsgSr6xegyd0b
bB4PNiWEqXBl8JGeySrVZziTAJg7fN4vtDGPImhIDg6D6dgSk+Ykcv0cuS1SOfFm
2wdnDagYoKZ1D1Gm3Bfy9KpM3Xw+dXLRJnBuZbI3Hw1I/uq7vtZ8fvHarisjAuFn
oeELQLzE7PWlD7sxLoDXisuNPUNvSzKFAGUnznEfJnjRmjmAIq5GOVN6PjfWLKpP
unRaYhQ3Mz2uZ9C8dnrfL98qPiXyvzLriKIZ82XQ27JGcu6RtARgzanc4XPXEUeR
R4JPQRk3NtDgvg9zvJWpi8o21czWT3Yyp07MB9xZJNfLC4M6x/BlP22Sy8zgUPvr
rKHoPQokS0IUs9hiRj4pA75SXr+4UFlcIy74Jfw0Te3ihNVPN4xMbUHNg6QQ+lVy
unyxkprIlXaS1xTiVRfYBl8BvwOv5L6sCnsiLwyCTO69oSo/UrIUqHI11HAzMN2h
F7f/20t9o+KHOHN6ICSqlvoHCWmLZWrqf7lGR+5FAu2jWuZqlDVSvJaq5uCpl4M2
+FeU3xpRQb7WpXmx5ThUCqyaHTZg8PNfM100aOGDvcHus8fEKnjVcT9vgguy+U5J
0QBq9qy2KUvRazIRgd8eql7GfzjNcg8qdry2QXlloDgs6XSFU9+wjsxSLT+D+I02
2PpA6x+nWGWLXeQgomlxO8Lq0cZp1eeAfaWohGaPJNGrxOnAYyFeeEtIlZkrTZl+
oD82OM69sdylChBFfV/lvW5sERTYju2wYdItgUMlgWRHyj7Bc1Toa6tjLvgA+KQ4
qctfTji4YaCKQwFZQ+piy5zJBDtoWd8bDbUXdJXj0SeMrrmlPoMv6IENYv7UsYKa
BbiNcUcSCaadd7RHc3geTGWQZKzEf0xk+BZxeHasZqTLK8SLpCe+vqN0GWc0/8ls
ZW+XiIeAroCA2+AD157cwC0Vu/CE29FDjTtbgYbqkUMiLaO4EQwhIbhupPLFNpOP
K8Vm35fNIjQUPVHwpAlkz5Rcc9YfrQZex8yLxAeGQ1sCMxkD7ZPJWQikkU4s2NRn
aW4SkYxu4RPa+FJEKu2jUr32BHh9OSDKcbF9FpWdR7R9oRPz0QLFcDJfh2TCwgJu
xHZS9xTzIiHDjGzJa94s/wmgsO2ZFNpwPoEA8TwWXxwlanQ/wMkU/0Afjf9pyZfN
b9Esl/QXQlOI4j2KOAyjrg9QZTjjH5BgBJyGF3YFREWpUJKYL3w83sWn5T7hZvpf
HgOQ2X2skF6JVsl0doFJb4EWPa/hjarLnuafh0BBHKGKuv7hJwMRLtxu5NuLkuaR
3mfe+S0wTdQQ1Q6pXTpGu5zPPWXjhqZWcJ2xAjzM1JYcV1Zk33kpDiJtm17UFYrE
t36zUdvTG+L0dskDEQz+bycKv8CqM58kKdeDRAr8TM6swn5p5rvE9jS38Xev4x+v
MMRVo9SWytOGZwrDcCOWCC6XT7cg6D70eXfPLoSHQAhdQIoiH3qPNBk/BxlZBCFX
A3dW3fBmbUy+jLrg4hgnJtQ33D0N8//liwGL4IprPBuCgvcMxmhs/uaRmlylPefU
Pc33y23yJ/l7GtjHcCrEtNcOkzSPpFsW8g/btAY4YMNFDiKOrqyXIcuGLEK26L8X
RNhMIBFIB0XFqV83isW5apELQXfzsUBG52D60cAb9pKccdQ//aDzywwBCLUMZOBv
+awLzPK9Qz9AFSajJmTOCi5DeYCxpwNxhcHHtYL9hyTMcb46x//4ozuc14eYu/YH
GDfua0e9/p7h6mVjz0xj5rV3kCTvn0gbwQPH3g8Ytl7AKnQc9mKC9R9cEEK+m2Tm
aAw63LxJweFlKzeOOIzjGlYY2E3KICEA4LGisp+havDo6OuEcaG2mlgk6BeP0uS2
ZiFNjExpxsXfeJMQxY+ugG8mNnp/u9dLL6/Ruw2okOh7/MjuKZcfAhGHiPA4Fg0j
DHlO1N1fd88hE60B/ANH8WCjPUThLwLJXmEXRMyZ3dBTETEe1dUcjJFZ9mCCKPdE
8EuHqDk4lFrfOAynr0Ibg6Vgwv/vDh64Drjx0YTZ7H9Y+yrROJBw05EKMhLsPR3Y
kQSqIb46KVYJyEg6/6/C71kyMwnQqlDyoIsHYHUK4igwikjeKdm5HcWSvzmcNEIY
hqf4Q/rdr/Vb7AUF9jq4rVhjzaBx8h0xjvTYg7H2TRfIEsplAddaM/ilU40F+4ak
fHjF94YiMSqgjndgIoYgXtJzhkTKK3YDp31KgitfkowjQmBcwH1LnoRSo5ljF/Fn
a1hzqOC/uD4Bqv0UcVZpmMhDP7Ovk0TW/v63tTsYRH4OtYncTdHBodO1QN0BTRpL
jGnyQ3qKKOoklbcPuPTNcTFpVcxTWx3U7UwBCHXnIwP+lq91FYfgkGg5zpubkM9T
/acZL3MurqgmBNROFzg2bMhUEoBqcTBRojVpn147FCIx1o0rKcQZ6itfN/ZwpEVw
6XZRfQCVPNGnok87Qpkx/wy20Lk3HMjUXdN8na9VZXlqzesgJvwJLk76g9isjBEo
bxxnSIE1I56zNgSbuWWw8sDj4bH0sCHsL+Y2ujFkiCxCeiDeNM8doKqKTca89gxI
8zvA+RshfDf8vvITZxzsoReOmJ4wxRTX6GyLqsCoOSLXJm1Lia9CovYDleuONbpb
XPYgd+EkxBJ87PMcgauROjQLAlcAEX6Yg+Hu0OjQ6cjiaAFtMKsmYMWgLZFPFHUV
0l3jcXSijxc+2foHt13yI5NEJl1yaY47eYws/a552SbgdRbEx2chAAyIVmVTfn8B
p9xRdIQKIMZJeUF8dI9CtIVEYaBw5dflHymFfSFcnlA1uSXof+B5VO/pQ6Sdbnaw
n9jNnw5WFMD9rG96d9ElhRncSTdGuQfDPzjcVvlF5GkT0W2jRNwxpA9wiFbn6YDx
ZZdKS4gLEFhWIAw2/aK5hd8cuVV9Y6Zcxh4/rlhCkKK6wX7NHo2T+4VyLN1Ci2jG
hqwLo6MVW0TqNpY2Di3fSvBMM9O0EdXwvCGQyWJY/+rIosXrjexfkbA+zqRzH6AU
hMztZ6NmkI6X2abWOitBp1x78kWtWQGPI2KWA4XDlDULaPDxd5GaLkXDU0G8zxzN
bW+wHd5h6KDGS5Ai+stnNNorztLVnj1idyJfPPNC0mtoJblL77na5RMaMilUWJ8b
rMvHedTDCcjWly7N8EReapHvE2rTrZNzFH2fB5s0/gLVzghxbIDwR32FQmqy3gk8
i8A5r63DrK0lUnNrjhI+pk2nWX6dDIw7BhNPHyoV6qKYA1hjqKMhoobeHm6qFNwD
ZTUoYO1sRY6IWoVcLeApBE01BKeOGr/cnUxaoK0k0yhVqrQELKm7xeL1R9KWFBZv
gYLs48qCZ0Y+aGjOpPXT6FckCv7eO2FemcR8t+FaeoIkwmLOlEPbpxMojzsCaGv/
Qtvnkq/qEperiIUElucID4e22Z2uGk2TxxOtWLOjh9PEdYYP8ACTP1pC2LZxRaN5
m34ayzCrDvfK8lEL1cJiO6IC4oc5KFTE3gDFBKgSTOtUWznnrJhX7xz2f/GPtM8/
rPUdxEEdWCQAk1NlTLKax0ZqJ72AzvEtzLM+85QpKgxpIMWOrcu66vCfECHX2tgr
5mriNKo9As0St7sh1jJYezF9QFx7J2dtmf3ySVOuOIKoK3JW4VWp3j/MIgHzGWr/
PK6n9RIgTaMA2QRlZ4CjdwqLgvRmbwlehB+CnupGdDjAVug4LN3cje4Q6E8qr1cJ
JL4DqNJIjBpGZrrdLaBL58dkEmtbz0mgHVfgsS3ETAqVE8+4ZLvm195oSoFoRXA5
qhlx4G84jPxQJDVMw3Nci7f5DxEZsvsJLPKrf2B+hU1XEXr2vzRqHtp6DjZHMZVI
+3vGkqnV4vHaqLB7WMtGlIsOdetLTq6rCdBSN3o0qo4ibKAFO41zlzlPGqCRmHEq
aus9OioSGQdKLIlmLs8Uy6xgQoX/4UbprEt1hDYJEsmR1BDpXcNZaDsInD8ma3HX
p0ui4rWwC56kDa6JWUTmcAZfi+4wzS9fm1GNc1VusJrM4byI6RFZ/tQCPT5kceP9
4RcI2DKf6+UvhwDn+Xv8rm4m9AEelDsv/hcc3XO/NyonejwWkVPNSigPQmKu2RDC
551FujNSuviBYo5IOM0MNa74gkHL9CRTz0iAfIW5gfnt2DGGN9OpHHo6mewzfDAb
1l8EpKv9FiWB8H2yCrMiRl3dOXwLxl9KHcSQVzJYowdR0idjVeMKBXh8G7JSVMqk
XnARVAdYu3mFf+wUxZoFsUqANJy0hHRvCEhXHHBYcdR8QO67XxShAvJ0zbFEWqWW
8pI8XsdvLk/ML5YqG5AEwc7+4AraC8x004MdF0KVEjP3HE7iVwo5t2/HEW1oTP+a
EuFKT8cCprpzvMgnqkVmfvpjDVr8iLEHXvUZS2zKUa9G6i81Y/pqwi+BSzUhG3Np
HqGZ2gPTCL/ZT9MJ3vVx5aL2iKJROF03fE34NzvTN+oBxG5RTXZiNovZ0d6SvVjK
mEEo0G++s8bdnxmdHyt0QmYaC+z9ywLCZAWqC00QkH2Ef2zVD3j3Tz5WWKvty0J4
yGEffSK00j4ZsMRAO9hxXHqk4gnP6axGdji5TevnDvrs1WAQIp/3NlvjTqU0GIGU
b/Ss99WGWw9bSz1CjgkPe2OfWeYlGdLxTKFzwJxoarcPRRt/+4xY7LzmXEsTbfPI
FfxWj8j9U/Il5z6f6qrRnVXOOACW6au7rLfJTk65sXf2rYy7l0vhZOKzed32yJbO
YesMCenTfOQp3OxGnCLSw4hPHgTUbjRxdNNStYCfLQaeqquRCUjMxErX6Nzm8DW1
kkuvzDuLY2+R5wYfihU08EwyGb8xWaAKMz19fhYIVsJ00XCxEU45z56BFkFcAfTW
ECraeyg1lUrYGGA6yeynAYxYWYFYKmfeDJzjnF0DPFo3bqU4KEYY03ctU72MeuUo
OTEuYvpwZFGWpr3DzuD9EcqGOgUw5b78zdh4pzxoqHAPISDrRySlKG/hmhQHTHge
QL9eN6BAVu9lLV2M5NURcbrQhT02m/xHIb+tZOdrtXcRpL13AYerMFojZNa+LxNE
kAVVtpd9RWFMJLH9tpAJezx+gsqU375ewCGC2nbAi+d4K9ISrE+V1oR1jfDa48sO
nNca0x0mj3dKy8N3K0TV9YLrGBpFgKVvYLNfm65EyrpHkb1Wj3HK8xAQQ531+9nD
GkQ3m2s1hPm7RpZ721LgxLYq61QajRKw/2MU359n1Zl6IA/dz1NFHX1L3jgK6X+v
FRkP2tk9TbN35OIUF1gG6I/PB8R7DNG/DFEMmnkEc8+tVO7cFQqeXQSvMTt01lAD
2TdxB/t1uAua216upCqul7k0IZ/WyIwbacovCpfb8mIM1makZEm6Y6L9+Vyk7dFO
vq1tdyVz6h5khF1Qejjq28CZyKxX/mzCaij1KacxWlOMv8vAiTM61cjZbHVXt5YV
Dl41CovvCMAfQdRUQwsObOUc0ZI5EcEYN54hZoO23nwfTMsy0mtsyFX9RVXEy01a
OmFl0OEWBVncUlgB1jJHT1wvb6MvHseJh/XNVXBEorED+v7VNI/x7ToMcqfjK+31
tUsxTKM3N8HrqJd8Jn7ko6dlSWfj1g0ZPaRGoAKwE3WYkCv4up0R5BwqbE2NtgTs
WjUMEmpi+wByvFzC+qoI3gNc3P9mxGybB7UWM6KuP+e/33fpkg2/1GTjsyoGLEVo
KwUl+oUofvpr902oUN/SK4+diKVYXkZIm4vgs7V1y32E99FKdAPS2AwVrazV1Hpd
mwgvlegkG3XZ6fCjLUWMElK0L88nLkty54AGG4aPo5WqKuHyUPO5kzvUK40cjFyU
C8xeIMA6jFjBCjYud0BLBlWd78TBvRtpR5ezdBEO/NHcMbUv27PkTQj/XQHJUCGC
k+yZUZ4FF6TQkCe4aKCcpK9q0mcG2dxcsdZSuARlH8fxPvsc9y40wexpzXMwg6qg
AQ0F2Xgvqy3PeKW62bkKvhOR+WDGlvdEc0QRxbvMs0AuQkvOffPW4WEx5v8hrj7A
x1e05at1FJaHJAGvWV6W2flq23V2Ohe+kwQFcyOO4qcUp+fO+9zlTQs8LF6PL0Y0
4iZdy/mpg8GXmfrZ1FZfgYILxG3SdHCPu61cZSkZsFlaXgC152HJBeKlAx9ZpsMn
Ii3DCuV2x1yI3n6lGBNv17E5j+W0C7ZDMOfjGByFzllv1Yk897FcChG4d8aEvr/7
IXoafEsA1prkZK016KO4vnXexZzLw8jRUem5UKJkjs8PQm4iZgmP4ZF2co8N2Adm
0HrJOmNEyqFHoh7Ej7fpDQmovBy0OwjPHeQ0XuAl7PH3qn3iHWH2Qke+kJdkwjDT
xLcH1TSdOPv7oCxj8yradfLeGH13p4fQM2rgd/YAKH1wZ64kl1wLDVcqeDIp3oE8
99N8kvs4HdHhZMKVK47itdcXxZJl76DOuerst2TNBFHRz5Dbx7mShdgSVwxktdc0
6o2hroelsvvtAFuC3O3ug4m/NZQKqvuLJIry5WSqEkYH4ndBjyf1XcWMSnGNAs+y
sPn/YaDv6AM0QVWWvwtdi/z2o9woyXVW+lKa19FE7mslsf0fsfupeETiyMoOoGF2
On+sz1DmBPESep0lvM0qmmq+FXrou0guKzYxzmpbDXFsrxsz59K1UdWxT02AjPC/
Rkh4IyiMlxmRn6LGQWSNd5aVbTGfhi38QDfbcT7QDbfM8o/1zlEzCm/cypATmKg3
sJs+sbKsgIEFfq9cOHOx9qOv2AQY0pm/5+bv6DJlMz5knMVNBpmDBws5f0O6Nhgg
+sszew8+GoyBQfTCmLFJTG3Xjo6kPU6LWjy0Ar1wxy+Q6UM9z644XKR2ONOtx9mr
t6vIC6mmrmXpLrbTrozL0hPrJ+kd6B6GXYnTOmF9Pw7SCAX/Ph3Es6KMoMlvMVQU
XL3b/s6sh/BWo+z/9zOQ+DXVcmz/SaxB8Gn0w2uQq9nHyX2bhcOtYHy5sxH3ESet
OSH17OplDS6xc6indcQ4enPxh5G3kubQDPflnVo/TdPj8a4TveuRIl0To2VGRNjp
QuG6BSG7JQUWgTcrbPSvbLTWr35dqEMcrDJYj6zfSwxGTf49h4HruTlfBmeONnzb
fU5iF1HC+jCX0CHlFLnmK/6pkd/mFZU5AbiOdyU9/YJ7J3s1REIa1doVieokRaZg
QroOvP5Fbj1gKj9fTUWP3N4lSTLz9EEMLset9ipkPnZnloIDuKZqa0wQjBMMFVK2
N1Px7b5vKxWc4VrBgtFcHSKb6Kn6IB9+cEAO/oNtP/IRRHR+98erR3utuGgEoXEn
dOdffLNeCDBSFb6J57alOqZ13Xb9ih5rMVfRclVLqNTXX7GH0lMPpEJo42xyhRNE
kV68B3ldox9EzFhQ4BC6YGf2l3yFAfxOSuJ9YlU8dk6Lovt/22yt3RXcOE5KiCzi
BOeSRcXF4k2z0m12r+17AW2RUDEq5kver1TEDU9Zgm6WVBr/cKY+diYd5BOM9Utt
ldOFAgbJ7p3PudTqu1ApDvhln3AAo8BBdnAR3LRx1b/E/tlzM3jF25mMDNASSC2z
B2JSh9N96U7u3g09BTPrr9f2C3I3krK3o7LFEDNSC6TGKnssu7p2gsCAYh0tMTKm
vOVSTEZujtdDQMvDJXEXHERqhomakgt1i0yF+cqk2VRyMv5h/mY3NJCm49bliHoc
3B1emKVJppJm5LNwJbb/QTWExrBhXgeDkGmEeBU+Jqc5QDpo5m4jcvQvSu8cHbw4
0dIXVDtsRGfbAL9sr3WR3z+X8PcKkoA/kpfqGKGJ6vYucVrAz4XdwVx5tP3d9rOE
PSRSlUHzdi+fzZU6AuYFED6qsDQUuXKgGlSGTk+oVGTpgFcWWA3uhFYhUXsaIcAg
MRJ9cX1BirslsGETTsetbF4+wLoV2oyu9TRXMUNy0XVOQdRFN0CNaoFAC3KhmSgg
EME4V0MRCv7wSP0IDz3Oop6V5kfggtwT09fTqSrKIf0AfRzULhP4Gaa1QUk9eZba
TzVZJ7xAJtoxlKa3PyVLGi5kd/yUHDmbpUNBLdyGrS1Hx2LRnUxkx3MVYSLjJweW
+EiRvNXNVUOuswN3H237aESe/b34PzX8T7PzSuB16Q385SuwbGY5fRRMSwIA2QKo
Z3QtiaJ4c3wRJDIo+lEbyylcvdmIwmyADeArYGCBNlbDUdaokes91qOvHAbntBzJ
tRQM4KWbnFx7tq3ydz6UUKEtNsn1PL8e9gjOoPB8zmPYHDzohQAhWXMT+FsuZynC
s/5Cn5PsamcjGKokidteF+bQWt/VQ3nQfLin9dMr27sy9ojIX5CfwV/iW5UQmOFf
f+PpWNr3CqmojrKjFEkyOudORo/NdCIvWXfdUm1YM9WH/qxs0Z4kb7tS0xB6osMA
NpCluq27GUZkvw4UkzPXJlv+g0/dvVJc8iFplVGE0oYxYsTTl0HPhGgtYnfAWxAe
5QHmJibaEySuPJCPFTZqy6LLh9CNwSLdP+C1N2ploIIuFf1mPmiGQNRPUV6IhrEf
yFPusa+bwsvcsS08WrgpaPzRz2lc/563Xitw2UoBJJ+PoDTnoD5VrZn9pJmsvehQ
NBV5qK6+xSfZXPu5vp3+Sv6Fuq0JlsVz/oD5dT3BhcF2iJlCVefK0bjG1YQdyAVm
jLL3Dac8cf0AiH2kCr0NpM/8KZp9btBqHp2D3wAOI7RI4hfijjZK9xZSZWi6zNVY
mmB0JzIwrYXrxIBSVIT7f72Cg/AYfl6l/vKhA3iCHWQjBHicokueb+ndVX3s9pjW
BVzWyHn6Xw40fAel+A332aQGp1QeY98YBPklZtR2qcIRCEhV8AAu2kSG+HjAMupa
wi2qgcPN9AVcSw0GGFG+ROMRp+RAfJGOquo4o+rWam6zuW8HzZx3SLCyBDrTmmrt
4NpuIf8zslkjG/SD4xRMd9srR6x4zha3VvJIp/BGtt3HVXpQQ7tXm7pOif3m0OSm
onmy6o4aJuUM7WjzbX0PZTzniKzq1zdJ8Zbb6fp9oou+bB8fzPh89iAXkzY3WbBZ
VGW2Xkathos9yvOWl1XgGf7jsi9exWIQxyQJGsE7sh2MM2euJJxa4OgZ35yKzz/z
qTeinlGKsnEyj+zPncMUt9O9Ct7vzJ06/VR6h4DrFPO55Ppy1UNu+dWyGjZNSN7r
hNdzUdW7yrhyCU50JhpNHLHTn+POcBsYl5/hwC1M8yFj7gOFWldVwVqb+7HrXG4A
tTjG/uEqvaN8g6Q4NlO2gakkoVTzVeyEnwSCDQ0J+q8o2JT0Q9mQx44zp0GObRBW
92LpugL+7yuBmYjMjNSwflQDVVa6WVaLlos9IJGoZoPC2x1HX2+Y1XdDKGs7MaY/
3M6n1BbQaBXN0A0roOsV88dv0Mpyt0M63Bl+DFvh8SeFZ/LC/LS5Xh5mDNe86QGU
M0jEn9nxENLVua7M8BVt2/x3a0jMtc/SSANoY7l6MTECfGRb4C3DQtG0eJs4lSBf
SyBMQNVn4NBIwjg9xuPIwgV1UDDC9Nx23yYSi5MnnXejq9IMGGTkueLpfRL90q+W
EHbVw/H3sMKTnVh/063OuGDR9E1b3B2Us4NiA3pNjqSh1crOSIpZ8H5FW5Z/8xA0
EIGFy04bXDV+QBNpYcSu7y+gO5CRVLnZkyqxpz1DzwL+bMBLFpI7zBS/ISSSgY1T
96XFuCy80HcJ7rBPinKGaJbWYmgH+Z/PGSSGnfaEAr2USdFnqXJZGBY+J2FugOiE
r0wfKhZKraRaUqBpM9cBc/xAWMGJXlDkGVZueOGxLYc1uJUgN3bf0J2jNl+g5g8O
NpCtIwQkgCfXKrwrYKHByuIOEPUglx3bArm/KOgPG7qCpTIndZQvafqAvm0fbwKu
B1dlZLXeIG5rfmdnty2z2Z8U6AzQEhHlQf8EOYtQZgq2ZNFjGvB9ygR8DXxoqBuE
udtPuwqx5dVxmrJjRhgeZaX4Fcl/JYhe548JxNilvLxgouTy81vQJI6brc3A2O3U
+8eKPUyWJ+QPJlXvm+0a4hZCdSfQ6/BF/hWzDRBJvH8wyJ2OGfErrl3+dSDkTyaZ
FBYMpy6nLUy1nve8EwCt23IPkCw+XOcH5brB0Rl30bOQCJgcB5iihlwsUFL6RLWd
RjnGENowFHAeyPMeADberYUdnWxfGMNWGycW9FSRdnQ6/kBaNTLsAOS+VQaJHaZS
yjdl6ipBXV79p4peYnB55iFRTGSAabyh80rWw2+IvaShFGIXn3vqovjQsEhlxsZU
8x2sWeIxOu6v1J/DkyneYdqhXVa9uXjPl+dTPb/gGEBd0x8/LBaGcdC6T9KBB1WQ
HWkreoSUHFblo3MFsyC3Ei/LIB81IX4FyNwegp5PKK9tkDIGzfXsQ0WTL3dlF69v
ch06JnX0XROWYhLJe5kDP0U1hEbEa/v4MzzsGCOWkHVrjasrCneAE/3gm9BHUt7u
rJRI43Qv2JGDc8JEyM+zuf+SxmhiT/LIKXKmi6MTdoWiAyGuUUwkGRBC5mdDQayg
RZ8h7HtufGbKrNfnoWO5FTvX/5Fomhmy/eRnxJUBPYUz6AbJk27NdRRiPbPbklug
wBNUp7pUg97HQFuk3pRztYDdoW0km9au0DR4M67+y/5XPh8+jxvPNGtkiqySqege
RWfB9UQCZrFzKMkdpF6f58qtslM6Z2bbN/pMT5lr39ApPqXtu3/QBcCobQ9NVS8e
UO5oronS7ZCUoFSmy75zH9i9Q29d7r5y97LHMynP1BFV9RE3wc0aWpxP0yaJMsj5
iKN5kt0Ckpn4wj3koISnd+D+63jIDajrMBCrv0izlqGxgeZ5HGas9RH8NHRyx7fG
JCvBVLtEDDm24F5TWcxHHcsrwrRSJ/NUr0mDDetvZfeIFoMRbTQLaTw4XluM8/UB
YRUBEZMpLrv52Lt4IKAxmJNhMpS9y7Gz9udM4JHjV+5rCtcs1PLa388lG+aYJI2W
A2YcnbChN3xAEw30yI9ZxJFkk58vs3+HWa8KgGFjUMvU/56R4Y5+/zHl6vvROi5W
m7RzWkshOjHSPxK21gPv653+JgP8xDJzNRpnLx+Ymkf+Qw6OSyA1z/A0ePkH4OAu
hLOobL7VapbbYo3WpeMsvM3o7yhxtELnRDcsE8EtULd9yR4uJDEu3y4W4/GctvHI
Rma6jsiM7Td0e/FCYkUI9+s9YZyiKNbcWOqfVfcqdSQePFWbzugxqiManeqwArsS
RUucDzqV0hMEpLZc78U1nlEl6IjGCKWlOR9ysmSRDaq1sEQhjCnH4DzfWmpylm7P
kH7nUc0+IN393LZpe+kRSjlvbfxXU3tsu1iaj7Zm1y1AXSl9s68TeM5rKVjvzjhw
jlwNN8GLRNCBHo4I+7fqkhCNmyHBhYHzkC9KistPtN9RHoyZzPwCY6yKcu6casZ4
XgFS1F9E9ZSl1oo7vomHjPHRxXcMLw+dV0PkkAsyQG16OmQAp/+vjSPMXRPThR7n
R6z4I1HneCmyuylet4O4vrpmS5kdwWU1bfil0A++1hSIeMqGn9xagLiHoKV5p6uZ
7F0q1ggS95/7YIFHIOsP/PNU+WJVc9GqdyTQUNbksWqMQLjZ64ZsFExFZaLKb1AF
2CFILiuHbiQmzSUk0s1+TIAW83ICeQQrA1mSIIBI4Btbu5gWeF2TiwnThERFsXz/
wtilpFHI0xGPt9bifT9YnITF51c+xUPIbVwbTUyL5Aw7RacXSXBg5R7xnGJFc7iV
Q1y6PfqUiOhqFl92vITskfG7vu/ScEteFdoFc96ZHF2GWraA8mFBO1GWoPrZ7CoO
bSeXQYHU/w1TlgNtOF1ko4izbV0uY0QDkJu8r92u2Y4l/At2ve67jceY0NFK+Xdk
+s8BObi1OVXaOaiR93oCTdULGLE/BnIg4qgtcuHSw9JJ30UTfoNEh87NwXhqXHLD
CrSPKwhwoIxRtTfsJheLUuV8S0mDd0Fj746iu210vDD0QwqJsIOBiD5ZDKr0hKKr
AWDHtlS5SONRQuVhteJ5PvT/fNqZ3RlEH6hR7G8YKyYfW+Sr82ztSMW7bCIcQNHN
B/6bjpk8lI6z/VDNT0HaB5zQ+dMw+JPJORXjg/IbXzz7K5zfqxOBalNsdfeN5Wad
ZbqcNv4ueXep0t4JhZ6eULAhQsQ9b+vDf2rMKc2zhMF56nMuoFNDgORk2qH/6YJZ
csX4a5P4zSs57e0gSpHqrHqVEdm97VMNEy5/p8RGB63l/BqO1LbQK37qJXYSwa4v
5fA7XmV/ZNy4E00O9+C/c9RV3kjSFsSjP2bG5VFWMBzxPJkqq12tmuRv6e0J4JRF
issdMvUPXeuAhr3yntUn4E29q5brPMHaWdPQ0YGXR/+4pZ3jDF543hOhRWKXuqui
q/j/ZL1D38S+dKB0U2EZuCqRYjmLZsBJoBgp+1XcsU7BxVj3INqsjcPUX8zz/vfp
ep+URD7FmMKCZJj/r3a/wSB31ZP9R1txxs4GkUQim9OBkRq/wUQSBoFw3DtbGQ0Y
90x37qSBAnhkDC5vRshMyK3n2j7N6KADyqsqup1VdWDfc2vA2lPLey6cZRZlkDz5
b/g5HfVq7uiuV6Y6ZYMfVbhHvF6cGHZMyXM+YYSbz+5xa7RKROZHec+Odc6zmQsT
jATXybaFdZsYC/DvSMmmzL0C8mjqoP5t1zqBgjNNP6zRHzKW2DmRFVtrQoLPH352
sYfm++jTEPLWUhQAKAM0MORArBy5cMJKSLZZtIIYYw8cJ+IUH8l9bScM/MXzPa/7
B38Nmjpe7nnWkyGAuS5n4ZXzsrZ5buUyAEfzG6x7Dbsz74fmdn+IG7QSEbWOQ4fg
BiASWZoLG2U6P9R6tsi+OfwuHEE5qxh8r0wxU2pnAt+/SMtB8DRbA6GVqsldUWly
5rmH0fd5H0F6llSzLKRKwIpvu+Lj+Hu7JyCW3UFaZzbuZQUqdvJ64/KKOhgwTbXk
iNvvK5IB0Do8LzEldwlfaBO9JtfGj7+X02H1AtkzjGh/NrOuJ3ZxiH7bdxo9+ZRB
FSqv5yJ2EkfBXy61y6oX6hUoABTzIWQ3Zv8+njyRszE1E4KfogfRkKCHWsNMz6ct
oKZZGXV+jFE2qcGG4KFulDKOcTcUzyUD3mLK/x2iwuMSQxWUS8UjHfxH492AL/rL
bl255zUoXZazIkpGq7nzlXwIuyLQ7nrf62cLq+Je0nO4KROZVYiaeUT0YdHwWlXM
qci8rxl5pNEaDkex8xGGs1RBBY0uec7i0p6KqhsykIyuCJDFkkci6b4ndoU2ycOu
mioPbALfmbR8Do8mtCNPyiTUmB4A5qqxHtSOl9q5L4cV+UWWBCSaemcto46F7u7o
4yVTkcC+BsRyVXTFh6PLX2xXbOpPQnVv/xjnOnBKZBaX8rRIGVmUu2Fde04iRR86
by0cQ5U7N2f/f2+epkvN6j+Jz7eufnZnvdvFgP4josTATV4w4Z/5UqWoortOi0kL
mykl0LdAT+E0sqGBD5htDR6qZY7Esgc+4NpAG2m+7TdVt2fUHEgvN+u1mweYrzul
SGkRvK6tpSSdGmHZPJmKGrjczOt9Lns5DIw4vD5+PIRvM0227m5Px0ttqtPqDTKC
07R0tB8IuvBqntxn7VHp5Bjlgv3G5N5FKu9BHMU8jSeL0CD0bRMNoX90YCR7gil7
tIMx+kMOqI3/kGcyOilD7gSPcWc+VQprcEHMIV2YsQ8HHpgeH9oNH6Hqw/ZkojEi
RSinQHotC43prM0FBrXEv9IW51QWPmdiAYyzJtvA3QB9AJEo8yUUpXH70me4i0JI
1LOdaLFqfZJ283JBIVc8cawHWkfwVM452yzQwdF8bfPQgzabXf8B8T722oBoLhUJ
Zr1zwdKJN4/urCE2epezpDMwQ/duMHpMksrxVxIT92Qo5mfJqxB9dwlLU67wesAf
4Qar6kE2Q8Ujawwx6oXm71yyOzdBi7mczidqisILD/5N2qI8B9ogrdCe+xIv9QJz
CqdSHpbaOirNXhEp2YK4SvCRyaBFYM3SCACb3NA5lpdkESjouN+lDqzHKAkz1bXj
lk8DuEO2o5uAf35bSbYmOuYbwfl0Uvm5HM97xsD/tjdPD8u5At+AxKX+lBqHCHdq
L31FdVB72J8WQI+Ww4NPtMKhw69OP8HlPlhmhrQPuMBJYvb6E6ST8UZEJqhtspbD
fgn9/D/XumP4qV60O9mWPa881xtpWcJdK3l2W1eXsx/7tYOGyKyyPvd2jyx/9Oh0
/otVAobfZFHYCyEG00SuTrh+oexgE/9PN3A8V1QabQkby/ceAJHnCYASqo82L9HE
7NGeNi44EwHm8uz5YiRpSh3vkrLhwHoy2J1rP4711URo4qdmDc9fVRF42JSWqJRz
KYezfCmwHH9BtGspwyEr5tR/k5mgMsFF86l2GeZQTy2onrvG1vttvwc1WaIVfXXl
BwoQHEIB14D8Ts4MeO75oURRJxlrnd+Ss0aOC+jz0oEcuy8utsxIViB63mh1PF2I
XqCYyZSRxonbOL3eR7dGoXdDDf5ftmc+T3Sd7pruUm+kn8AMAaDyS3HneFM+r7aI
QKRFAMbXiFItYhybODgcbnvI0TMZEEx1fVofnOd/vj1o7kyjp6f6Jlh3JX+FV2lz
PVXuSfrCuOFjI5oTvNA+XrtHAeiSDHTz8IkA6J39+5LEsshuaxWyk324QdsRp9Jh
I7PIi4xa6LRemnwbcK6LXbBsFk9TuJKBvN29fzuInvS02jffjhADcSpBw8Der/Ci
s0eTlBQ/TBdx7IFcpw7ZS1sUq6/MG1HulSUpP0syeJXqc93lB7poAMnbmigtxCpS
akLFOobUt5PMuf+qS0rN2HtOoiHtgwsV/lNp3uKJXWOdlB/o64PmH0EHaXbmyKOr
7SfATbcAoy99lWDRV2dxJjkyi0gbMcKetR5QO70bjRMthnKIJiJyZnP5KfWnk8jz
OzZrpjGd7Vbiw28g3LsqEtP5HIfwIYXYQUWValX7F0s23B078Aly4eZBwXCbjzj5
y9xAlYbb4zdEcT7yaaSX+4LJorU5tCSGNrLcamWFffgeRrtaN4/x8LbDvlVC8h3R
kGkAD8BrBaE3occUqXZNvY8JPVIN6bO29v8K4F4PRsQRyLOeMf293gEn/voHk3fC
Fqo5TRwIcEozH/s2jig7m6sYtN8eRiYUEw2p3roy/QizKkQo2gKLaCcKSSS4hMEY
JoZ9FtnX1GZUiouJ4da5HwitF9JUpQ08X5xmiVqVuW2uTXOkonxUH6qVpdqzDdNF
ZznOQSf6xMJWMXLXZHEfu65A+r7r/NYIYHWfnto9pyC9MWLJx3cESB6VHpIEPVEo
eswb124jIPAYGd1xL2xfxHVTe7pdwZ3WC/nzDCZ09seovUThG3ewI8It1JYxhCBW
zBXccMH9kEJFGHCBWDRhjHdfcLscYCfG3rOIUaWmxbvwltwvzckzq4GqmR/X1WJ+
7Ub6nEZZLVrp35b4lmepj5x2FOIIJtsz60y6alGl43wtlCHRoscfEeD8hDTYY1Fv
Qkq2UCDzlgNajUQhJa/DCwCm/MZ40uXMU5Dcij+Nibnx/VibggjdRsF2AWVsVblA
WUb9x+JuXBXObnyoHV94jmb18s+UwRzWVQ6TU38eNAdPisIhL6+g6SuBzpewNqwL
aVsV5a5ZZ0pdtjBvQlPC/wW6LNZH3oAvFErDI6LTb6mPxHRlS8j6T3sPJa4HNDlY
YIpZvmAUG6+tMH8Q3BOUz+E54rM28ydIGmypYDutrd2XfB5j1hRG7EAwwWUZIsDd
gEvWxjrVB0Hduh34W3SXWSDrSCHAuz+AWGRgz1yU8h5XZnR2b2uPF9yl11wSDEWS
63NH5Kvphs/FB/uSHPCekYzowd8MRTqy0UvCYD6chrlQlk3b8gwKwpJHtOfAEh0p
67ibsCH/g3FzMTx36ZotxbhV+mnUDLbqHnXrVN5ViKfVcbg+LtD9qV0r36nnPKBY
ngf3aaSZdbDB7ROMge+L2kzlxB93O8hfmd/mevGFPLUW2i7w/AzHKltYt1wpNx9P
b42ZGfGCeyUbw2y7aXCC9NlbPpKQZetn8nl2R4EeLZGHYl7I2/MwOMLQaYdCikQp
kHZqT6wSbtzylZjLUMMGC8E1qatdHJyXzLHp9h6e/w88JUkZettUicZ7eGY4bROV
NKt5xDY1tDmvfPS1ZgNuUsxxfT5wGIwY8ZnskJ+jlUy96K5mohP6mmjqmABoo9Ux
uq5fkKN5Pet98F8qb+ds5oTPf0rYrQ6Z6dz01r/S3Zvfk0pq+MFCYzoIKAqRRoh9
4z66ls4MYaVqiuQ7txaYCYQ1TclVoJ5ScAD8euldnh0A7HehpkQM3SXA8/uSFYSA
v50H0puZQ4Y85/nfB65giOpOvnrwwT3oLl35Ioq64lrSmqfAmohqLXK6MMUI/yC3
tVEoVCMsY+mrNUZqg5LMfY06KUgWcrnoOQynv/lKOnA9FCdy2MKoxmfN+98fiEqp
k2AdQviYG008PvKML18MNwFpPm/XUaNm2la6gz2A9HGHVPt+lz0le/ufmploEQLC
RMlk4/Kw9xs/S7X1XCFWsHbUdLXsf2IhBeVIVv1JYdX60PmTggV+t7w4ozHOStkn
OmKvg1ibDZoNLSR3P7UMUu/P3FSt+uA9pLQrKPND1h1D+gWX9BsWcu1iJn2ce32f
2HoN/wt+SntSigM5zZlU8cFXdRgLJTScDPHAuQZdQ3CcvAkZCuwGDKA8RbY+loj2
MUlCUeHWP9ZkAclp50HdYfHC2HmUe2pxKgLqfaZ5HcnhDWbaagqR0jUoI4niIEHk
1lAIqj+zqOOhWsYIolNWzLBRX1dinx+asP+eNuuayNGHTyjiDVJJhu/RUfiCHnTk
W1aw8qWpxPI03UsJq9x+olz1CPPwg7gBwlMwdnXK/kM/OWOY7GUcS06cIVx6edqr
0iLC6nC3kipxg7dwAlTJ62lDQ6Acvc877U+ZZ4bvOl0jQcS0h0tvMBNhlmHB7AjH
EAWxtqu5TSw6TiUDntA5gtNou/20AEcpOV1N+g+cwyrL/0z5iBUEaZGk4YwxvQs6
atLuP/bTUU/R1HaMEChjNF0nVS1FqEP88OlQbyTbiHjdf8iPsRRLv4614qtkNTGG
E++Mf3PUpkSCaxZ12P5/bbPVxlpbpOpVYteobU/4o72hIcsPZmFClkdiiTguyQsv
3bWOXzASGuS/6WwnW4GgFyAy/fdL8XBb6awGiTk6vZGGq3DFgNjn7cWyjUV9Gdsa
QX394Gpo/vHhfZ9PpNZ7NlIJdGfrbSGNR+VS6eo795Eew/iHVJqlQoVXRfb2KAYn
TIjNzFkgaRde4nrrsMsh93SLKSGX/Rx+wHUBF83yVicvK/FkU41nw101/orm7z2q
O4WbrYZcJgjLNpB638P7wk0pK7jFIYbyLfHK7WQya+F9UDVtg5nvOpolZkrye2JV
RM5xh0AP16h19sjXygC4mbVBoKML3zI53JTwX+5xqsR8ekWoaQ7w3OK5uwAVoNIk
b5OEXK5Z9w3OhXUuHIyuFnyqLeJEhADUkTJwOHXUVMuESNtqaT8S1YzsHxlsXMdB
P0JOqan23geIiJzsuNgIC46UWx1N8/eUCMo3v9d/tLO1MSRctySJApDcMF0nZmIH
NrTzW3M8heFdjkfiUAJAbm3EmKzRihnyF+GK+p1SWwbX3ykIdX5M9dO5SzbKxDBc
olR2+C6vLr9A8ufHtSECxWFkBtnLOGi8rYzfK8akPl7c+EQ7e71As+z8qv3hUmCF
wcbwQS2LPE6YuvplhMBfWKWER7WIt3tmz9GI7CqFrJQQn31E6X3FGggFdxSw+4Wi
kJErWO0aTzx6wLODRwoUUtkGvutABcnayjUiglmvlGnuEFmNZ3dqSpU7r4oudDX1
nFB2WFWoFbY/puwZKqDcnv2RvbxKLNQp/9UqTHOvU5u5JToj6Vq4JU6PslGaqyI9
iuprLXCR1R6/Xd80WAOG+CoYmqmtDABF3BQqlTLfItU+gV2IUk1dkpwafcuHNKgG
V9HeuVE9aWziyU/JqQXo0EB0PkqHgrUmtNlCfmnoxcYz5/szYsK3CZ+d5+L/iHkC
nN7LEC3VXRBJrRHzH2XM5U6GQjs+vpOJmJOZxy2ZG599SO5pJ3zEix5btADQplPm
H+Od2RdWDfsehRDI+hApd9NnNy42xDYd69iOwpYM49v+nBht70ynWNHQsikrPavo
ufnpGj0Ea/DSQqYguXYu8+xjvyffknjUXOMR5GUMRDk2zNpUfLa/rjeow0xA5vSe
T7tVd3rvwz6CVKoCbW6hFLcMTa11VJutK7EAKQhGW6AnoSR8Ts6GQY/H16ymoq47
zMpN0dQWKyrad5ugH5cARR1gMkw8OUbDLlzd7ha3KQdyngjkL0lXXJ+jwLThNACO
4I5mMS0BxLBNP3nqxwNYl0NPt74IorhSvZqZbVZrxdZSk89ddSRFK1sVin4TZ0qa
ButsYOM45NYEiwoYm9H4zUDgFR5wttJTEamTPJcBm2BAi/dK3BYGBOPN171itTeB
0srUaOAnakGqg6Wzip0ywst4x7ASL7fgIilQhaCJwMRluzlUHSY0YR6YKjPoffga
EKk6GiSizrkFRfdIGpmQRoSRH2z/WtyQHkglGQk+9SCKSWcPtRK7kxvn3k28R2dj
SLeaZO79wOGuTEzngiGrGeZIfESoiwdErSbtBOxO3ZFz/Ri+s0BAVcH1DDyTMIzv
ljY79FKdZGT3mANhod2klWhEGNppUj9mzGFFrV9rZcfBY81eh6M3GEkXqoS2CNo7
hUGhFEue3kpkTXKerB+SePkKRJMkFKiGvOFcThptqHgXYgeOApyuqbNPYWbgTm1B
mU4Z7e0kA9yX46MND9eSf2EYzh6N3S+Y1eM3OnlojeQe52Afvl405OBq8ud+azGw
xZ/Iq4syh8dtIhlGR1+R4ZKrF4Ear+rrhqsDbw4l2JVXzZETsoY4csQBlE4mvVR9
ba4kC3nDm8cY2i7m8reVhdTBYu/0lGB8Ca9Kzd36bntR+9lziovWpqFjnYSAZxxv
3ryegAhgoDexN591tyNcLQfBv1Lc35D8LDR5FrdTV/fSfnntnIE8+Dfg8l1YvnAB
wKF3tbMM3AFpfbcOROgCGeIKzvA31RmAkP0CrMbiv/wvz6uCQqJBL10+me/JzVzF
vHtQBMOAgjOubeF7GQOLUwn9PBlrICD5Us2ZL1vYjsCLOH4fkToFEzI/AzD0ODQ5
vnRtFwZFddzWg41CFngiSPuV64BFPq+NK9OOFI+A6ov1G6KPzAMfW3VbcmHaCAws
bsnJpoYLArruraqtBqCHwoIHGZvKR+MLDYiOiTzNKDXZCBsc04ZgQwJcdaBZf7ON
ejuwrO5eNjCy479LC46xAF+xISWfhi22owxDEE4l4OKCKn8wA/r02UyMHbFm0iOe
HAoA6DKlslT2CEvui9l88uXBO3K3RjGMdwC6kdQuDdfMw3BdMl4Akv4u1ZCktdZl
4yZBXlQxxJk5x3H+oZFawehHSi2CCJMV6EjR6JmzAwW2d/9g+SfBOd19Sr3bh/eC
j5SMLC9OvVwXDWT4vGVA/NmLBMPBQ7BhFG3/4+JYqT8y5VDUjWQYbTC4P4Z8gbZY
M9SqmGCYIcwWxwNV9hHJMtsUcYCQ496P1nFUYcPbuvCE5/Ch1WZJMlCIRSgZp9JW
HBgxa8uR0c0jR66xVyW7h/8jPCVQe0Ys17I8ls5Wo/2LGTHg/3ecucEXvN6AkpO5
fl4z8xxFA9UV+EiRI6EpSToQBNQU5fa4xltTesjuL2EcKr4ZleXiw7AOwl7OY1o8
qilmY8jcECRa+6NYaF9lV+YOT8QuLDVLp1DpwrZ1UxAJDFKLU1FJpugI2CHfbg3E
Zw3forgcqgWi+AtY2eH64sqlm6ISrNgFw1yq6RQiwPXDVcN4gNP1XWdhEJJqY+kL
29dwr0i6+QV78DwqWBqMtGuSrrS0iY4/E2FN+beoeox7ZhoIXcSNTq3Xp+0QXyFp
T3LaVpLpU4gBooUnJ76x1oLJZzXkqkk0buP4NPrK5uYb0RteGGnmjDnapIJEyWt6
y2CyzghTjV8P7nSWuFZlaGTG3VlqIMxbgOmv2T4Do6KK2SS2rTjJB56PdZh0R+rE
rAB5eWLdflS2QOzVNeJ+XXgdIp5oUtX4eS3sG14MhJwqkWM3uushYEss5DUgDTv0
DIMVBrjc6j30QjlIWakjKlC6/w2k85hiCsUpAYeAbcGGQki107iELpRx9tQRbHiP
NW8OeIf3RAeMuLqPT4ibtODSASmKSBi8VpUCQsoCuVY30sIyoMLaYIYLxZTsPg2K
CiMKgKohmC9bZ+1me2B9r0bcleiigWzGoWzPUHl29oB8quEnryQ4NxL+CmlKHNkK
d05iu3ixqVFrYYMZKJFij/2OaekNNcQr5E7EAEJqLlQE42LfYWlPHGdz4VdQb0OK
cjfeDq7s7epHRLTPFnm2u5/SJZ2Mb49FGC6KJ+fL5jfXOSWmOdDpjFk8bVHXusaJ
TwHm5IF74rqZ274rN5IoQ4D5IUs+7MSp69Uyq0PzytHOVpt4fMGrBfh+w7sauPXF
UkR61+y1sB7vgCdnPezZvNcPn2rUs0o20aVEh1Nc+OUBcK+hbBe1dpq1oIlJJUvH
ZvIrTQSkdRzCPGSxbQ1z7yPvgp+2Umy18KRUwI3UJ4kfaZrvYjpeVnZ5clzONha4
6Bg3F2sLO76LqNtjlioHVKGkDF+ehImRMz5/bz/T9+1M4uvH5UtdFLktW5xD/cCd
ooo8bo3XkKr61TPnZ2p2IoyqwnbLTogu8bWW0mEeuzw4ZrXW9IiGhFPMOdcOAUrp
aehnmj3k9Cototgzvty/PbGjK53NNah9sgowZUCBUw6ST0psk0NG2TMdzt3+qVgB
EVemwQyENOQ8l8sbRMmBj8cy4Sih2Ip0Z60rn9IVJ5nVRX0h2IVLIkb83qsicj/P
dE2MfxhAMLnBHEF6wrUUH+ONWne/BWPJP/RSS+B+C/nu/rwLhym8AWUghM8swHMI
6Efuve7aaRvqXX+dujH6cVe63t7rHlgIinVuWEB1IFZWm4/rSNySEl6RifXe+6Gl
M+37BdYsdSsbloFoLe66j35RK8HVQlDgMoaJN+Nee1JEwopszSDFry42ouV0vnkZ
/XVwghA9gCYo8Vaz/jPtWWeYW0Fu7fqD0fPq7Ct+ZFyhSeenip6dRmcPfP95NxaJ
LN2YlrFpv4Dc83JLNEVHorzxb3qOswPbeC8LBYNzJmHtpoOvsjYBFBsgG1mQhm9y
y00SpvzMyWN6NpS3ipHah1VR3OwHXX5gubvHht38LpBXGpv4M5BvExupGzfhWoEA
9fn01tWIpVnADsvEylYGxSUkLl3L9NLjYPY7dmJewX7quZEi5pTwlPvUM4p5zqAz
2EgVE0sV3D9FX52D08YOiucQYnt4o0grEbWhbjV19yY/MHyEadyodg8KDjjQZRwK
lucflLZZZ/BYwskKoRVZmzdYOJjcJRIMPpdWShW9eZv2/YxJAqlG9PdwDVN3a86y
DahGDkLfxORQn2ESaWyNaVeW+HXJ/gyGZeJz4mJ/nrIiLXedYV1KR6+gdBzP5G5R
eHcObaCiA7KYUG90tL9/h8TQc5+sX6QLOZN7oVTjCz9T2m8VTvGDEqMMNZkSpXop
/09rFX1dz+A4QD0H2xKDprgvzOtQphXozCVJKJrJ5W2l/SImzVqAF3TMuAOFtJnx
12ffEYBFPC6UpXIGNLzPPr4MquWPMBUfObK2YKTBuGk3+Fmps+YJHQXwf7yS05qD
Py2ch7N+eJNhpMPFwsI/OGuQ4yIeCuOVcLGuDf03SBm6ceoFrZMmRRkLInDCamsc
p6VZkgC1noJUXcKONSoKtySNrq4iwdSfezSmapkbCjJcAv+NBCFP6dbwYn904Cx0
BiQTz4wW5u1nfaWML7l1sHi+Kjs5Sz2YuD+VqQoJjBOutRQZoi6MVNKznNFWtRPb
3MeLWIQur85r5G0ugpV/gpIrgYQOh42Qr8MptfNTC9cyXREQSBpHP3Ejy7rWzsvP
C6eyk6m+CvGSH1MdPIWbxmjmmSM0VmkR4lp3Em+cWSWeMbCoLIZEqc0XZIQak4yO
YMGyllABRTkrZvGMz6+L6DS0+V3plByTdOJK5y86VN52EBVbTx4Rgp1RPq4kARbD
qAwUqZbVkDwyS1g5kwzJ2DB6dWOS3i0FEl5ARp2xk0h4pH3fCSW6oBnvZvrs0il2
Tz781wmhKpYUChW/cYpT5eXRjPbcGWbhMXP491T9aKr1MgofeKYfnDSQfLVMSW4u
hYsl0UFaG8SkLE/nrvDxB0TNtqI7tU0Z5D6AghRr+3qFcwKZnPup5CLKMxTbF9TY
vSMEqadlf31zTujj/0a4Q4q0AWo20OFlaUNWiEE44X7cUd5lnHsM0a0BtCfD30jV
NLH6tl92XsSGjyRbMeH/Nk6kvkEqPyJOO93EPUpawSMn89TOW38UCNlZNBXZwtqA
BasBah136mzLbfRifEyqj91HaBAsATB3xoY4wSE+xCGzTazr02rMgTEWptr7oqLY
ufkonpDNgAjqw3vxXeAeVv2ODQE1LKNo69jylmEdcGOi53bKx4tEeTYrFJmaln9c
5yhXYCfDgy4sVy+kF8sNPt0rLkVxlr4WC9ZrnjCz0F1p97LfZ+nlUvxeBTmxwQ1D
kqHh30CNnITTSA7bLejJcMESytxxBMgEv31kKt2CuMzLb5NP8FtF4lsyYlH/6Mnk
4jgb6SFEOgd83riGqTGuFH9QYrSa8T13WY2pgUbloKA/zLY3zu0e6cLzML1i5Cba
J3O8CX3xpnu+2b8Xhn4LBAlLl/glxIF86kDjzIjjQX19u21phYV8ZvkJ+v/3Wx+8
KtXuNyDpJTigJSLl6bdDBNGNVFtT7XsbrbAKD3c1zE1N7rGlUOmXIgHVlIbtj5Hd
78wzECkGw/lRyYzjR0iEGrjnKX89H/G8MsHq1pQbytjYyFYW02pinujGjZH//2gl
66VZDIDlrtgkDqrl5CAoALydPdpE4aqCTIEDWIeK8BIJMr04eI/r36OOP/+1xf7R
+tLOL+vK/VL+9qrRIxp7ZLvvfTCKPP3O3l3TiPtueDvzrZAL37NCQHmR/byzDodb
mVQoeJR9bFKkObTSCdQs3HCg3EC1zJUF6+y3i0/YfB3uhq3YXYbjp3Bnxj9syeKi
lI6tUJHLB49/KphMuoUmhRPS5KYHQqm2S8RAsPs5s2Zp9L0a4m/uU3dN+455rli9
+wpsGVXOfkakcn5BMcAJ5VroJ247RgQAb7Mac7BecPvnmhazK3He+PHLij6Pyd8J
GUpHPyarSEHKBxK2aQI4ZL1dg4lNFFUixFmBnPopu+Slbgfdp4K1GS440tOiBIPV
bsoBItDTY19yGOaz0ok7yHazo6gh5rBG9G7BhcoJ2z0Kb0Ra/1AdyVphn/TC0jAz
bK+Pe/1XRIfIFxcadLLFBLoR25wB/5mI2N7kGl8oFBnKtNe2EFrI23iY3E/Yi1N1
PfYFED5rSQ3g1hQxbY2zd3aygeiT2uiRjDHYqQ4c6bObD6HQPEBgU8zQu3SR70WF
RJlK17J/wlHhD7mKPeK12vAiAwkq8jKsl3w1nUrzN8l7SHxTjOStBKV5UuLoSCcX
Z5NrDIsCSW2ESHWJ/aCq/uOZF/oDUCrFXSsIRpiKzBb+V+HQhCk3x5+dGo6UYyO4
LLTh1F5CgxDZ/vU08I/TKR2aLEJWUOt352Fsgz7tfCw/Arxvxqm8ivVO8Emh89Zi
TH0+9gduq3JDoNTS2XtCZK/9cYOMxB+4W06BU75K4vdAz9Oli6jsC2sQCPCkoZ8t
FlV/oPklmk9W7jOneHmnQ2bWapoLm99zmkywG4yttJWoy8IWmiOKp9iiT7pn7OLg
//2bwac/OXLtvk0xgaeE3Xtv6H/8Yz9lzMAr5niw93AzkG3Nj1HJLq7ALcWPzwLQ
yWtIxcwPR6KzM6EgX8CcZ7UfNqR81lW7uXhYs/7lLInI5mJ6wzus4d0bpsxaB0nQ
sfPkE3gzl4YlwWwX1dGWnZ1C71rt2RFb6EEEi9TH2Q6N0OjTHIp34WUqnXmsdnXR
0nH5UTdpAGJHj2XQCC/2m+tCMi0AOgRV5gE3Kw0KFvGvsG03srRq+//g8GNKVTQ0
g+Is9AK7k6CmfRn+g3owBaTneMW1DE1nkF8gp8Hf08y4NiDEx44AB01CZQxn8wiC
kDb0L/zyYawqJZTaxnnVpz3mp8/fwveFcr8PIlfi/dEbpn+n3IVys7Djdg1hjWRZ
3iCVYeiLQRg9w2es+/2qKBDcK1DqBodp2KgumTq4ztj1e6G7UXfhqcxLMbVQ7KAh
LM1SnKgpDKewFIJSp21+1vqx+r/7k4t6KCnbeZvkVQ3Xb2lUBUYoqN2522STekHF
GIW0Dnf800qlvtfzvqny6UX1uYZDCOGUAf+u/jqGinROAMbz58OaH27vJd4taR/6
dSHo74vo5I1tTSsTR0NcPTghwLFqzCxTPy+ZG/S4v2AZkLlbqyC8XAWsqYKgbMJq
VEWUN/26NTZLOJfzm9wlLdAEzP5Tml9Chi8FG4luaB09Rqyk65gKg00wRuatsyi6
HxEAZT756V2HDYJkD/1WsJFZoxqOm2ERIR2JT2m2FJZELTFaylc8IQjGjxnBwQ1P
W4X7OlLa8Xq7pa65JfIFXi2/7Bbj57BaOCQmgWDvn518YB8eUD/fOfATEFkqwjp9
NOqI+2OgWXEU6zO8Ig+Wmv6cAJxe3eXHJ2rZqgUr5Ir4ZWN5r1uXfJpm3c6MyrQZ
lZTSzzv3HObV91cQYKpfR33oWGRiZLUX+14KcpkyTPqn9Zz6bviKCHqP+MP0EaXB
eAFbnNIdBkIcST5s+UAoAKybOuD1t3M2H9iSxbBSEb8HMKa83MMk5BLWJPym0bTH
th26vvby/7AGzKUkhPk1hUWRprS4LEd6bb1gJcZ/YU03yYfKYIj4KUHyroQy8pb5
Z9XiV962Y8TiLNpZz6cP/q5h5cmszJYys9+U8OfZecgzTqhl8f2vANIE9sieXmCj
hvYVr18vDxcawym7/o0Bivt1x46ckx6OSmQUccJHdMzPUlpILeJDgEJYG5TqKu29
QgipgkUksmmlRL/9NYPEFOoDqEpmdadLNKuMJKX9PjiWP7+v0fOe6SfBmvruxSBf
TViVNoxmtNlYXONj/hf7cXapQspK8XojP1F/pz+O87xITaSfMBAo6x/ta2k5fQ20
Dub029nzHdcI8DUIvYW1/4qI1h1cs/CmQx6JQhbB1FJcPtDOFMuNas6aHAYr/eB2
1ZSY4skokNj4b7EiDIJHBCAi0CxEg3Px+B92VvMoJmj3jt9lrlGFKAd3tvQ7+CVy
VaUlulObrK3FCAqlWOZOPSh2Ow6Xa6mbZVAD7US8GVtMe6Z54qQdb3zrDGSBD0DX
vAi8iy7o5M+zAynurvitXx0f3OOa15sQlUn8V5mxTgWsOZ/sSxV19cn92WQ8ThZF
UmoPQDhJpmkYd/4WdE4WCLTOOBkIaVd0ddib8gnUpJW+QCx9rNCKedEjmJpyq0wr
6lLpUglP+3Vt5ANs8Dt1540Mx/Nmoj+opI/r5duDrtyk4Nrrfs29WBK803GvRooZ
tG4zV1t8obwbNRK6IOaYb3frmeDUC0shKugodtMRWjRR4vk7S0ZKk5O2CLkufIUn
OljOiwIz9OwMvEZkVBYf9hGtuot2nqic5xh9zNpR4Sq0nCMJ5v53G+JsBq/OZIRw
mpz/m6yMoSFx4RgeUtbeDkI2QzEZihJcgbvof1+UEv/9RNHgVgGdgxNcFUvO8O9J
JWRdDq8VDSWDD+kM+cw3D5Cx/uj0/SgXMa1WqPE6s9c65dtJNMV67REPF2M+9M51
02BRfSwUZ8iZlwD7j/Kw+S2bVtofKhGhn80epdvdWqWyOm27LTahXYJ20fDMmdDM
efyJR2K7+446qZzzbfW3ylKy9Fkbi3+7jo31xvdHbcGroGgrBWfaCEhcUj2eCaSR
8NUOm/ydgPeyTfc/V3US/qtdBP4wIXHzoie/lKwiah326YfoHfev8uzMTbqByyHl
e/9J8FOWDgI9/sKwJgYImSPejQkgNe8HZZ1HB8YsEgDdhubMQGKCB1GOLl+WzUkD
PajlboPCzuFAuKN9+A60ecY2a1/j6+tuIGxllEimtMaLJxNlRk0kXzejE7cRRUwU
eVjSkUVJ21dhPqv69ydHf0pp+Aa5zTYvR1N6wBkYwkmG+umXsT9J3ut/XDkpPquV
wYpIl0O618ZlqQsbOYCN51fpavxN8DTFHbQc2MYxh2navy4qyjRgBmBnPdyoRvsB
M2I8/oRYV80nOep63Nw6CoXv3XU6Vj6XFx/JmDul+sJjeSg4O5kYf5FEixLx9Mse
qqzAJ89g2JIe7Bzgdv3Olpju4KjIGigc+mrq2WvZ0+SnMVkK1oit6uWNMHwEdTAE
n23T7Cx8YCSkd+hetHQpmaGFCjW3Ia5nzbcq3xIX7perNROIrWvnKsPWJ73v9xVF
LgekH71s8Db58U3TPFU5Hv/VBfvCDRLqQ7K+ksfQyvGFDy58tAv3Yws9l4+zhPyb
p/ZcsTEgxe12RuNmTg42JJFD5uN+IdSwalDGwYQc9UNHNi7d1q44q9i+8TkULQHD
oYQTXIORT+TwaVqseja83L/8v12RsUbPFFeJRj+VQJFFT8eR6LPrwxh5ZxJAB8VL
93FKD9vTd+iRSDKEZYvSudYRcRBXVImbwPYbvM9igddrW7upghI2XZuhk08sk/it
Q9DneD5AKdDs4Ls9Qh/uv7rabOyEu6Lq40DRuGXsI1gB3QECUEdYVX7AaHCXPrmU
AbG6YXzQeGzSblV2QaI4weJdxsOs2sTDjB1R627u31EdHmXDoNGHppj7ywj+Ax4c
fSO+8MvRQBO6Bt1jmPfLEEfCcTf7eLw+YtYb7cPnV+jDOWr9UKWU8IKEkjQJU6u6
HM+831W4uqCTniUaaid7E24rkDeNWO21hlVN3h6Fm2dDtxmD+bBsyZoNX2CHcCkk
BQn3/ZDBgTI/A5c1R6BTVjBNen16eUKGXbRHxT927kxFcG3vZwmI+UsABqHVIajw
y6Bge/v+ehgW0S1nmTR6epYYqP88MInLvC9fmD+Dlg34D6EIGetQnEbZMICKwB+T
PjPkpeRNTQq212pS2i33+8F0mLMG7YrVgShSY5kEmPjjzf7wMxwc6Y4ELwNAkzAS
zgFrs9HP9YgZ1bm4orhS8h3mMp7eQMu8rXTE8nP8IEZa2dh3x34AgQ3/kGNJbQyq
pUeNdSUkeBZay7bBvw+1y4rBuh9YNpCiolixoMjZOVqdMrMYuQWk/ey71ZXjnIuh
YHhZ5PLAU7n9OZLacLP42JcirkExr0WrRF1iOllcoYMZ/HpM4GJmA98/jm6iv51b
T3qBBvoN2stTYFloL8TWYYMTHfbGnt0S9aijyJnlSM2Ln8a6Sm1e/r1cbyLPmJkZ
F8Hac6S0GSStCKFiUEDMDRGAJkf6gwYmSpngPqb9jHJoeLJvklBf/d2Acyt9pt02
nmLas9ezaDy6hY1bTZH9A1nw2bTokXcNgKPuMDCeKskdn2OOhbWVS79ZBvoO8IZE
mWL/27soqldTzE8g0B7VHEkZPMTEEqkcUcgUWUbr7LhpuAlhts4O/yv8uM+/D6Vv
vFD06TQyrBqnrUAhpv/njmWkjL6ip1K+bcVm9oWW1OLqh/4C1WIg04j/it7Zkz+x
sBBGBh6lkMs1KGH5jWCfubWF115rwA8S5liVHMpKI9pz34Z2w4FsEn3d5hO37zLz
37bl18893lBfuf8ioqY7hVnEOmfsOZLqDpdX16S4os9iG3xPB+ZLMiB+DOA/Nm59
zfry0Oo9IXzoIywG674dUhwFigUoS9tOm93MPN7Z1rAMHxs+WBSkvwNL2LXFalJt
CSBMIZ+MVNd4JkQQT7hI26MsPVvzin1BgTJ0nRYIMeslI9dnU+Rqup6JN1/08ird
MmZT8lOAtDRpWXZRv3QWHDmRNKbIE9MqkCXmkeHsTjfRcPFCsHYypquSQDavftcW
EY9w9JT29kXWtXMD62iHPWojno7NXPNzdKtuS88hpxSqg2bJvS7l8bBLJFq4kTUi
DpbbXOxJMEgbxcH0Ssi/zgKT2neQ//wu4RtEXtB0Nc874pMkz6CrZgSIkFj6aUBe
CeQ2clFo14IPi4s0Gyo1SgdmhIdXCrkw3e+EiaOCzK76vzeBTq3u8PIdeGtGXkp6
J4l3i1zGxg8DJv29lYdvTUsnB440ucVR41rGNYTKwIU2oYq437Fo9S5KuB9gWhOU
qhWrJZy1jTXu2Q+49DeTi3XILzXIacgj6QMTJFaiqpA5Bd6Qf6ltE/WPCzWtkDCv
i6qvLQrQFFrXpinu3c+uvDM04E4oBFTsAFnKAKMMh30tNptz9ukDZvQdMoC5ZXrW
75IQVZkPWw7nOHQ7t/kwY/m2/c5aWCv/Z7iw8/ahU7tbquMXHELamG5Qg/2iPIws
SVERKwqS7/h9AmHhdJj3CqnQQisEJexqqE54gI4fwSeYfdJHrw8hz5H+Dp/sbOnx
9/yFF7DZH7USt3oBxg6sll0MOoTdNqC1U0LDotBHC2OZoeu+Kdm4ln3mAxNPA4RN
JBwvzGvpV64GBindIpEOBOF8031ugf60rakd7IGyzWN6UqDWIAuFJnnQTyZVpduj
wZnloukhdyUXatvF4hg+yLuHBaql1vAK2U4r31AjAH4rxSoyZYqEWqS6o7Q9dSLI
kwv0JsWYBN76LUlcyNIM8YzCGBMydTGnBxjZNIEKql9cRLFxEQxVYtneYfvr5Er5
wKnWIuUO304T8GMyxt6v5QNMTvTvIbplIRY4bN7mHtPvTleZBDOZJCz33sVWTpbO
MZSnnhhG2/BXMD+zf8uZstNcW82uITW7jJiWZUmRBtWu+bT23+kjCeoVNIxGgqF6
hKNJb4F82NrwtHU1F5m8uvqUJFHw9hvESrsXXbu6Ln9wOfX4Nm3Vr47+7EEpXM76
S2I2+riFB9GIgFlraCBPf/Qu+jkfZau7SV+qTGIHqqEeDtnC1BrnPJzoZUIeHolH
MGkGhfeJ6lLDJCF+qoLsx4blw1zVjSsmlx8ALqYUymhoeJfLvOCvjSQAvPanKKGd
zKW39kKRvqhxaiIVqs9nG+aNxta7OZCeXUoQZ/IXOa22H8Llcgs4/I66y5g5sJ0k
ms6+zZSsO0HqFmjvsTsu8NdO2tAGv07D+X4DuQgeb8k0u+Fym+a0zoMgjdvi+6jy
j30iSR9Wv4uWbJF5z2wFxGFI7Fxnat5zGePALENS69deIl9+ei/iPAupbZIx/WC5
CzLaXukKfHCX547B/ih/N3BpkhgLoGv52336reHY4HuFwghsQsL8MYKUuWUDslqO
ofEzk/ntSbOsXvAIUxtyycC4CRIoGp1z5CSkkP1V8g8yovJd4VaQ6YjEcVaGXFXF
FAzL+LUjTskExl457VLUDWgksiQmDlBJVeZ204UXQVS9KL2EyfZQNsjzeKifLQ2S
rDCl7QtR2bXW+hJq9p+QupIciJeoT/uDnDC1uIW76P8MARbxp0cLCkC+oS7HyubQ
j6Du2FdXrGj1pASNgKT2QnUELX5GAfznQOXBUZTq+2NJDSiSLhrvakHvTaXH8CYe
eNd7OgRd2XjQFmBODU2LvMh4oe6b97KnmcdKcSb1lad20RwSEbEYpwGoaHERoAka
nd0gjcphbAAWhWo3JTGt3kNLrZdcjsAFMKLKU3PnLiNclR7i/YNt+HLt4jkklj87
1eQ6M7Xq+MHDadlg9vF/BtIM1bRe5k79aZtli1PCR3UDAlw8j4b5d4Vq13jsTt7N
q4W2spKriGuwB9U9sqZqtmJ7iUtssvKnFnMtQMwL6nzU++DhF2C7iz7h+KmrVnWd
DhYSyZ4JcZzcnq2S5QdRWlXm5StWwzJsH87pWM85HiGNhDNQCU9ebJK/HBlJf0UW
Y5fcuUH6p0cSBQQ4OrNcrzMxwWNiJhNryGfjKtNV46/BZYy0th0znLqig70IWG07
9FIYl0Fa888wL+rVZtllhURXqOQMy63KjyJNOA4NxcYxdm6RTryLd4Do/carLU88
fMdjcwGgMObz+gaBk/s8S3JI9fDbAYgecSTKRoyPpCtTIo8s7qP1kKb7kbcRmp4k
MMe/1ohAvsVMQpTXCecD1c7c+p0aNGXzvhRmUGRTzHe1KZGSdE6fT961MeJhZpv/
kFcVMEEx7ltOrQ96zPth/ZIBZAZXegWbOo6u9+F3/MUOskC3XnaPgRMSOAhE0htJ
JoQLaSgdfCJ9+QE0kgzRJIrsSBnLg4nJCpkVn8kBaZetVNe8dJ0T4EGwXJy6knpA
LPf+HfUZqDfGVTyFXzveBKmQTLtuVFDaIBZ3QaddL4mkyGKkumrj0aAv1zGAkqmY
sbbnDm8C8fXea7OWxmIXJw6psKgRk4RKT+9lA0Djr0EXP0dDogc77yUeOOCbwUus
+9xzZegY3UnyZO0WG3h4NJkwtcMX0sVHDLtDzTU6NfKwx39Zne3BANaWKW7rDu96
YtNBHtgnuLYdoIn/Pu9wFD2tvlzTfXb9QRnm9RAx9yACWpHkKEnI0SDHqya3PTM9
nKT16P+bi8oqaj5mrczCQ0DIJWI6dkbi/wkNZUSXORfenHsV9PUeupIkyQdHJCTB
qyxF33GLhHKgJJe5agwilrHvGR4YIhvDY9QG0tqGDZtDrZEPzNo8mv0MeCOUh2+h
j2R5w84RiHIri0Sa1V8sO2bpvxZ5uMf8+HsPfBgDdnQFZmtuc1PdF4sTi2b+NIkl
KQ/61GrF8/bOZl+ZBwSUZbnel3U4f/LGbDkaNxtKragoLCJHciwl0A+6g82OTIqj
BMyTCOq36Izv/sSUZpXbTabXZ6/L0F6EAB6IUQOHxCXToJzwsfNaSq5UU1vFkmZC
c9bUJkDZktCoMlF23RFvj3sp4ddxdUAZ6ojt35A5ZrGJDxsqJ5FZbGMPgMQUJskk
elyMcX6kO8k5rR2afR/udCXx5qVVTHHhelJxK49D6L4oIwrJVVIylt/089zS0CtT
L3RDTfcoWbfm92AQwPe6/opSkhc6Tf+1kaWZFAbXMMFLV7F2aL9Fb6jM7kbHJ1Ql
BruJE/Iwiag0IUK/MuC82kvYCz+S0Cjv6KxcVOUEM5loFFemqOW94uV0gJDtY+rs
areAeDhpDr89k+fCiMmmQIhZMPO1kqtyGPVOTksU8t4h6BkEwyXaEAd48belbfUW
eWHZ/MFML6/uItpP/FS4P33lU2PS0u08djQV+jfBNjssOU3U2i0Pt0OiMxzl27Mc
5Dpegvh7CaXewuoL0cw8+KY4MF/rtyWhkfJbSZt/yVkcR7ZmUbUk8QSYYqMEKOw/
cNgMAsl1zU7mAhnX3q8rY74Pw7DopH2gWt0ZTuO+qzG7IMAXGn4SIWXtAed9eF3d
LznwR5XWbeQU2BarojC8h+Afn+az1CMI8knpjlFu9JiGpSosy39BbyIj3lLNeHXk
y07BMS9i6NpJbR9gHMcnOXFbZrvYyZ7i23Vi6zS/pMAoAHWHbJdxqQEjrC91gF0x
vesWAlQCGx/S+cHiBQNUuYu4BVG3lfOFTiNBeTCiDJO2oyGVWrUkY8cuNGiVqr81
CgvuV5T+PkeNcjzHRbggGKFpCzGeHPLdCDSPZ8JK63lllRkeIxNFpnBi+cGxJZkV
Gy57GrbjB+IRy/0BeqSGZcpx70MHa6Ss9i+VpNfmO08Eg2JGZsDwhk88vB1rUtKz
ifpZgc7W1grhODBhmh2UnE+R+qRNKwC0J6Hzq7jhOESGGD3FedcApZRGKAPBMJaR
+Sa3P0iZEfGgPcd49fssCScWcuGR0PNWSGDtKIU7bRfueLCJ15r+ecdRXLzPrZyq
Gbue6B9B552SoOZpgs8EIsYdpdW96UaK09twDTMZ1TL5kavBFAyFnoxEfLOMO3Eq
JKLP4EKIqWjhDlH4TRA3b0G77JpRpexXZ2xYEuKOC67mJ12i7FGkojDsZtcFZp+p
lwxX6QPggqhB+h8FkDlmLsDntnK2il9B8+hB9ifrsUGPlQvkCbquibte+k7xayN9
Lhrj77q5M/+Q1eM7nYzicvUvN8qNkYzSRLRAYAsshhczzsMpLk1ctNcUNZrgxl0J
efpWAqH1GVMej9u9m0/RIu6yjhdILGyvbntrTbcn1+LUBX9g2NBAPQLbsEloYoR/
kRdUbQWNt6oYLa+rgjCxHCz6faxBaH9D0401EqqEqgqCB26uvgF0ajopkV9/utfD
7NkEVovnoKdJWGIt54tAjQCqYS1P4BPWSw+c33+ONI8zzAofvtIFvPx68KFwm1XJ
Dl++3d0oh+td4e8bjXs/fuvzRdEnxxtb+qAViovGHlhSRVjekVeWi/8Q2LoDBl7+
+4TIuNy/hAmzXZ8SSuycalBFYxDTDUwOWRYX3dq0lP4Q3XlJ+iliAnMkO25vLPYM
qXt8XO47tnWo1zvnSHwODXfClPrHeLBuE5wmziCml/PiIFlqUiRKI/EEdHDP64Xw
yveIUVwbA8HUowmx8wm+k1iHTwvCESlOClDSBvyVtfWzTBsrEnkWWCme4FyWt0D9
Jwmc4ate23lJE59p1a/1yEz4LpZ2i2LfZ/kKbFdkjH/bBl+ATczmyYYrmBQrqi2L
j8IXz+IbaSKkR2ll13nCHfhl34z/gUSNBCRtwn5YcfIv6oqSl6bJtb2Oq8ChHwAH
9TsZwM1YXVcI+6ounKsu6ph+bsmhAyg92unJQgV+5OyjqtDWYAx6g2aygy+yEDAv
ND1dftbmojmegwCatcbAiHq+5ZPhKHNewhtebH33wtUkhoQ4wzwQw4sYRkf9tv4n
1T3PfVqgvcQEw8P62dUuQIhA/Ex9ZGlwoSdpH4HkebeaxLoENkfNpE9Myc/Aq4tC
4akMXLn8G//tfBBTV6EsE0OFPp70nE6YdrXx3VujTk3tPpfaXPtgv48w1rupzean
NrIEEErUP1I4NeBwyxTCNFlb3Pi3qc6+LbA/VWUx9G0RC43wM5RBus2J6v2nNiN1
/gs09BbXOS78KKxhbrD+J8SKaFY4YF1PVhXn/qIGX3Ug3vX2P3qeVFuDUhRXJuaj
3vbPh6yIIG9KLLCyU/67FZIN0eJCf+BKyaqGMkoprj2xA3K6P5F4gs/vGPBJFTB1
jtpiT6Zp/nKHkQ7tO4WLFQ0HPYYTcOrTbgUlBGQu7G6TutAtxbDwnRFG1jS4d27h
9EzWhM8GJ+AdQSEUvAPPMa43l0bzGIIzBBxkEmrc4ogpjRaEN+WCpGDakrRXhfkL
A17VmgOsGSqeIkMXRSi07zLyXN38BqyAFEuhPzHKsy6wyRcSsntLfsMRgh75enId
LTUjLlJDKer9Y0w5fWzxWvnmB5VEkR9hYKqoN2r8rUbXGPKfgImIVhlC18m9Dqia
gzoSLhzn/0LhLtnxZTfOQLnSiMTy7q3bv38PJ9Sqj+UIAkAvOiOeyfyeW0Gg+ftM
ByxXvb/4qFKxR0+Jyb+HbzXLRiSNdYh24g9UFFjgH9Lk07gQyv8TU/1WYK6/Qqe5
r3W8mk+R4IZ2+my4gfG/Eou98P2DMlbVQODAZPRN4fWg7iKDBHvrPIeHt4CCdLYD
veFZJaYdIS1V2PXGEKNed7R/mcla4OpOWPoDv1nhgK4/UVSUEsAhd4huCWdqaH4W
rtaWzucXStneZdhTztSPpDitQerJT1wDK/NQ4AszxDhMr64CGSjfGW7J7j08a/NB
WJJrt1+kQYGSkyicBLqJxlqdCfwOScX7dD+Qs8r7173gpGuvVEjV8DGy6Awr6kzd
UiprvWLVU6T2bre4SC4tPxJtgq5UYk+hLWXxoahQCZ2p/haNs9uhpmfGER/nDfkK
nH19/cHKwtDypn8ZAEOslAgbQAhnm3xQ3CehUpNQyGCeaaU8AtwQnHI9cCRIYODs
g0ytLw4ykVNPXc8TWB6D2mer8+NTe9dBSR+XNQ1Ns+wg3pEvuiFkWkmLPy93FaWw
u52p/7OQftJYNrNeiMtvBqrQna8r16L+Vua5eSObwxi6YsspFv0JUCL2RGvJUMLX
740htPtENHcKnbmuOkriM0z0iw1cQ+kSSokkKR3UMKtp7VVj77oegJnVXZB/prPB
BDZz+CXld5UdUGwQ2Vc6HrK9gLeGV07m/+2QZxp4P8RlWm8DKzd+mDAWTYP1FNz0
cppkgVn5GxcMM/WLqdDQD1CKG+bKi09wC2/HdphhVYkmnmdwCuLjHfUiRR4gbMTX
FfEtJsBbdFLcQqMCbEvnuN54A7PpCmJB6eadLZK1jtaMIx19QOaw8GDrkAC4DVry
1GWO8hGsV+yliUJQR8utzYsCy7DtMg7vZ+w/EFLPLe3qfIzkrwgGM8+CyXMM3z5z
YwFZQ6zJxPzT2vHTX+rmtvhoW1tU1obsWBvR6AA9qbAaHqJe0wYXO0BUTcQNoPIh
Xul4MAUoQ8jfQCCcCglWOgs7aZ7qK6/llBKpHgAdgIWjl+6ef2GMoq94AutR4nZe
fRJHjr5F5C16lddvIEyunxK2TEfBcpCQGQE2frSl+PEBADeTmr0pHHwZh55qek/4
OTZLAMZaz+7xFE3H8Lhl09yH91/jeTnzBzGopTZEJLE9/Mbbq4gD195jAjbhQQ8L
QINY2jj051Nx72Pk6fYWfzdBJL8tdcz690jIKN3lursg+PpdmKTq888e4mjtQC3n
o1UVd1eSwmnF32cFJkv6Z4oW3hzjBY/apGCshINWHpBaV/fcPwVOeA2iqQ4TARY/
zwjIuupwfLtvZnfIHpEgJ1ULUxUS0wOaRHSJWZyXCTGRvLogLC6QjSfW4jnomjAA
wvl2p8AQ7eSSn1DtGGHp15ZfoZfpZVCXUfzbtqWUbSvHrsc5P5sY5/DGK4AuKOSK
2QAYScjx3pv2ZukmmuSnRU9yrtteH8FYd8KrMfrUaoZ3Of7R93NIOkV5rqXQ3foz
lhjkPT/PbipBRA23VwNzYn29XaQ6dIsz1/bPHcKBb3ndISdrQu73L9XkBTNCasq8
stel0OCyPEGWOtbpg5TGNVO17Wb3F2RxcE5Kam5uLbcx97TZGONqm4PeNp32jGUy
QLVa9QRePtm+TwSteAH8/Tz7AcKZruaViRwfQuSaGVH5CpTy7j5vJmL9ySCZBrgU
Qq/hmoZEIinA1Zh4EjE9RtQPA3L7EM31fRT7ZMTkLxx9JApdXZvMl1h5UJkY9cKF
3K3xtboNn6gzAWUXmx5GzAtqVV4Wi3YFNvwDDwmF7e8XKZEGfJJqzSP8wFRFH+av
SobktIepm6pisI7fUg5mWyCpidSeQKXHh/leQvpzcBqFyImZhhYxLm6839MGG2Pu
tXldyg7ei+xtAdc2BXjCDFww1UbYOVNAySxqPT6HIlaZ26U66baPIkSQ1e6jW2oy
yTZskE6hX2dls91bajkS3cEStQCvPlekNR5I8Vug+CY8OwEbo02Q00g/u7t900jW
m02EUXtO2JXJtVyqqE1ty6B6JAjkmGqdcaKdiCZQ84UwGpqPY3GUU0nCIBmcZO5e
Z+5QDzBtDXvx4dJ5mQI2ryN5dsvOX3RE53JcsJA8uSWv1XQXAUXFIiCrN6EOiL5g
Di3vcZtZ0Tlidb2gpy8xh0j64iDGknramgHT1SGtpCy87pxlvEoYwj9ngAzJSVjF
adIQVDHdj54xi66In6zu3VpRwz0DYWmC+pOqZtQFCcwM4Lk7OVp2ezMW9kCJn2ux
nANAN+gfzPFykasWMaMkUGIw3l5y5XLiZ9nGowBnqEKu6ink8ADhnJ5O2GUy2PjX
nZ0oxOIB9GEubMoUN3biXkmHaijgVOERtq6EMEaPCBcEMUQvxlcbN1ya6a2oFelA
KvrVglG0zPjCnTrVUX2X03s7WGBiLE8UUMo207gm5+tnE8tPqVaeY3mGMKlBwmZO
SJ8iUQttYmq0xzvgGnSpuX8npYBDDq6Xf0L7V/Nazh7kF6tFj1AdkVQkd1xsaHQU
CUA3+4SVMXgW4YwuqpklFJY2sK4KFf0yrYLbng71RBm4tw+W3+KuLiT2VUnQAurZ
vSr3O12rUu8/VfDn6IDkOWA7cUJ3mXuAu8vQEpz45SLWrkWKfs7L7j5UJzR/ZrVy
0UFYKXA3eDX6uiHlohCQpY94iUYsvC3xZ3JQcZ6EbbGnGXy9efqKG+i3bqxQyhu9
ysYOUZO7fuJYfq7h5t+YGasIKnsF6hQIsc2JvNj3kl5/1oBakJjY6cdp37XIbtU0
zK548RnASI+aHQvEGkkNikb8gApv9a0QQTzQ9r8gbSsa0oDkEi6SPEZTaxPGEvOg
Ya9rpYy9Rudjq9NxX6KweDHSaW5XAGvMoQnnxdDlQUz6yoCLgo0Heqw4/QV5O7lQ
E8jKt4P9D9nfKybDKkiPm+orUycDL7ibDKfeP5l1b8SXzKJj12/ElMbpq3p6n+XO
VcNYMnJL7jXYaBMcFRgv7bKOgZvg/zC3zTaU48TDmBXrUrcbikBtnDIf/Bo+KIsr
lmdwXfnxRRti71HPdxDgabgPRMvqyiORV17mlH+dSSEWQFGi6BBEt/pri+/Kn4Gy
UxUBDXRpNmDYiJWLo0PxmVeHWllbKMs34y+jAIMu/uxpOffmtETXheZHZy/xvUc/
oqCQ1Pj/q1MavemzSYTMNsC93YCUZNgjhXGM3HpPcN8orDjtDOM0Y6VAa5lqlx8g
5H1QWxr1E5eH33H5WuUw+1uJWAtYxwOW/jWfm9b07FkY0+8KLskuDWnWpeFwXPes
RACE1fqICOYRQo/nseEEg1S4YLDkuR6URcjloTLuO6J0WeCS2+tcQguC+JlnImg0
h4SLneHg0Ppu2BAlls2zHlygbKkhk6JvnhY/ztez0nmTEmlrfr3dTG0Nptd8ee6w
Sy1d0oLP3Pd9BzqssCGbDUAIlY2rrKOfOfic7LscJpMMXEIjdC/jCAphfsrFa9d0
OiktTK/lmXNFlATdmx15wHnKZVif6nfQnvq7axgHl0o75+7thbGeASWEY8ywzxry
3jnKOn9CaLJxUd5lL/s9d6eF3muoVHOtryolUoZsWSndzsrU6pdHhfTvAYRzdP8e
9czBvcpoyr1myL3nWSneotBhY0brenDD8kj6Zu294i80TtEKcYrQi8KwJSiubBhX
YTjUsoORKLvPr4JKEcrJw0W+cnbfbDyhWhkyrNaoGIpbbxWxYGcl7DbIAQruNcHq
444DffVLeQkacVV+Dti8JGdSKZwW8NNhslzEzYYN6AL4dZprCglkTPkilg0EL5cR
Rx4Ma2NEuZLdiGCLrMFwHw7di+6yYG/KHJ8JBFdKrmwzizMz85wcYfhGsUezyTwe
9e1hxIhUe46wVSeuvFJCzjKwyUfhB5ccUdEDjh4thnEBrVN82ki4GK7kUtwtj2FA
FR8doz2UUE8OZodKYNvwopVJpkfquYmZAO1YHslqybtFdUSONAiw755gulIngD5F
mbKMCv8X7fV6VSaPSmHWa0bfLLUhAPuUYsU+s1GHotXaXlP3DCV0TF9P18376S1Q
v0Nvnb3H0N0jimH6E0d4XWjyfLmon776xEZQBcm9baVH1fb9Xq7Z+3nIHN99/fAs
ScDhIEEw9LaDk5uMVgLhBM+MD2k3tcn6nCipxzCYFKKednbp9LBXWcEfmK/k2Onx
c1Gr4dmJMuZwAlSQ1R+OAusqWh5ub5S+BJcBDJd1lZ+pTJGTP3RLsXuTkkfClpPV
K2utoEIeyZTLt5VOQ8WCSUB6RGgvvxmTaRAcJXE5cj9JP8MUZIY8JcMVYjYR4XbG
bv2kraCBT9OWyrJ+aLjcEybakD3imwafXOqvt+DgJDYNKbSam6DqgWe6N8aFJtCj
T2cDHeK+8L+hnWAt0o/BPgziXA+EbbQIicmxfwyAeyxUTD5x13sDttzWl1eLvabv
9x5+SpACkxKMICuuOHSLNMq5qR9PwLp1OS+NFAqZbCbU+cI9wHt7RxJIA8/IOhW+
MiOoxFnuDcUYA7D2+GoAZ94v/ktuJ4owx2s7KDCWyJzlD2ECJWUypWFdeW0zriQk
XEOog2Fj5+uer8NNwIi+koZ/Qo4lX6ng4H7uKCYK6DGeuI0ltNnLY2QcQGKf+i8Q
IHi7ZBZAU903UvwUQzJOIo8zIQWt+qYpS9RvIzMD3BRJHGgoTU/w3UEA3J3E3PyP
cPphInBxFBBlR/qcn/pvhVWa723xRsxMnYdGSsb22BT8/3v304IDyM5hlHZcipun
gdX5nfaZgRKlCTmr7kAgZxtpWgXXRoGgY37YbQFNdRABMvEOM5yiaGlQaM06Klnx
077vViLxYV/hi+f6BQIWszWby0p6RDM2TrzF0wUmxzIqOcjITRHKPOgk0i+hM4O+
cFAFH7PApDQkahM5mmrV77oKP1NNS2pTBwkiOO6YWUcoPGhDAZ/TNGfQcX2N9bsR
jsdYZpUnJq/Mw5+ybhJVAQNrJCN4VAvKqqBXfCn4aZWCbxuwvSG0gd0lNpJ8DOEx
BoPiyApWpZu4NUiaICVNOF+zl7FiRuRs3R6fbDP85pDv+kT2Qdi0bCBmjDyzfIJ3
DZKdpgAl2q/BDffFVFxSg91uNj+pPThVFOK+PZl1r+KkGTtmwMg5v47MQAGX/ebi
34/6akGy1QXLik6PbTTzTkuaCQCllFqmgwojulBn8iHhl6JPipq6wICDkzJS1FLQ
dhEHefLm58AQiNBNM0m9NUb7fXSYt4FiPt6j3FE4bxvRQiUf0SU6haM+MJuQeKCF
zqiU0ak4w3Sn1aIGOjBxhdiLrMBgsAplab4QVBzMjDmGcA5Gn8te9KZsHDMvR+5N
DdnGhHFJW8HUQhAnQ1Sb/bu7m0omlgzDFq3gotlLH1N4hg7aAnS4DFiJ6FHyD7tP
NlarbKAk0YBWgJGPUG3erykWVuCH6lazl27Yt0xT06a2duZ4rBwcGTTaocGmMNUu
Oxj0BBEzIDLYgTwotV0OJdJS024suigRYcA8VrUe5xmLl5hmq98YGr4vJtSL4W/E
jmQarj0PPGVeVJLjaRbCrh8z08sdvpiY5apDEN09VWb4SS4sy8SdSXgvYOV+7Ho+
b/sSC/yWYWAGDZAuT/u+wBMDfoX2BbdMnlo91g4Zeh6bkimd1SHNdhu59ytKKPox
atk2X0uXcJfyuFcfe/oYJyPBbvM/SqmXhYE4NT80CtEnlXVYAw9dh4MyICltf9fa
Z07qGhBB353aDp0qZTMYiH7VCHbnvyGfT+mo1FICUeXnlTSLwvTErk8lrsHE+9p/
SqPOJmkpSV6l5Fn7lwE8xJM5fkEiSc+EmrV7hICfAehRwrBTOCPyEtZPpeL5/5kD
JB9OpeBKakIA6PYFhhwGx/zxnidE2ypSv6zYfOVnR8RClsy5IUS/GF+YNv/RBCSw
yaLRO519XUvXcrfMMr7AQBvUZwuzoisYaLVTdu9bqflyB6MmHwrdKE9Vv0mU6YXw
KftrzkTYl86Cx2aU4f2aeKMBHt8CqMeeWMLcEY2RfhDznHIlLnmiAD8WtrchdHZC
nbOMnIBUq4m3KREqtzkjuYx9Org4fYmYR73Ocwzk4a6yLEpvJpV46NuSwn8ac6Ex
9+5l3rIqcqZFC9Zx4AARNqD5KME3FnmRHxhDUuWbwtQrIXSzdFH7T2ahu+xFSM16
zfmjNi6R+Wuju8zty5PWUGXGkqIcH7coTXKI5gwnGlPC01Tc8MKyCAG4jz6wgjw3
SGXddbN/657ABe+pj0T0HmJuZKcBb87P7pP4YItiAyhk9eZVBAjf4GRtPdefkTLn
Gy+KjfX59MGtLLmj4YuWINiesnmiTWUZ3F+6JXoo9yMLhKQc2itVHJkPyZkvn2/m
eecdaN3ZgntmoCMEIiID8CyiB4biPSFjJ19PwrbdhG6p6JZtfI/np9Xih25CiwvQ
0YgzTpKDrKXjpS/P6+Pq5kvtt6MvR5jaTkJYv02SQS5yVMz/2ll1C104+KWMKClN
mcR5F4X+TcgTl7XHUATxzvl9wAdsTjPIYBjdiDkKsKdDVo63i6gLFC3EjZRWtyhn
ZfH3K69M5XX1oylxFZzvj3OIy56PIKgMuITbXDL/nJt2/igvJrvVHS5GXD/FwozK
XX0+djZeuEv1RGf9iUR98SlrzBx4HOiPvRBQ+zxJ6270lHhapdcEfNu7PM8uDTel
FXZfbtr3JrpnBESvNoUNdQlFw5fpyJEs8kOEfS6fO0Kwpb99absr3LyCMp6yrtN/
pSUUujZvshjp6p7o8MMVKK1byfdKuGeJJnQiK3KK1GnyD89UmDzsPnnQLl0dOlFj
O4fF3h/VUU1aXCL/q4ilGbCOKMAzoH4HRyGkk8gc4dXDAiETVxMKlREfEdTcZR3U
VlyA1mPpfJYuaXdocrEVoGCfpXZA3xCHwzZ4YuEQsHPVw/YL1Zlg1lyE3bZ9NZ07
4eZGZSvFBNFD8otcw5zsLgyqRzyqQL2F1IKw6ezrANrWTZRYiVU4eq1nIys9SXfW
8Dn2gkTROPSYLt2ALn4nvw6WP1k+yY+u6n0i/u3qtgFVQKcBlGjnFDyL4PTF3D8a
lDSMcPUuxyOvx96S1Wq5dXcCP5sj22JtxnWTrg3cCzHFdkKRpJhlsrDwGuCNbuNW
TbTzQuHFveYKLZxHSg845dJxNs6dir05rrNdAaOT0V5cHgU+t7d9J0GpSk0US73A
GmJ8JQjRePFr1gKz8dwDecJe4NdRBFLKhksHFkWlpgdI1OhXsJGC6ig3m1QJPb21
bn68o7i21+VSLls8fwStCTSfbrM8NSozr+JqPCt/tdssEogEVFA7yjjL/Dtlgsfv
BTV3pxqQkmvoxh8g+42KXNUXhhp7TWVy7akE1g++yar/xtyhM+wqA2t3TNAonf9Y
n5UB+bMcW+3BAFdLk0HQGyFhyikHw3kKiw/TJpM+rJ5ose0FPwx/8iBWIuVPYE7p
oIbafZbNFs8yzmCNmD8FV+a2jG/W6d+PrVJMr0YubEdJQejXl672aJxv/h5Tyl5u
whXK1KsY+pgO4D/CpfqxEksUTzsMdFZZkOKb89SVL66R2XCaoFFPXJonNamErF/+
V089cSK4iXaF8GDzdWl9sqolOaMclfgn67Ccv/BEFj1gAUaWfRK/cRU4SnhJ2UUp
q/+aY00NVzcAZI+7ABB8fxyf+pT9u+rqcQqUEXaNqr0oZK1qQRb9PoLs3j2rA+rw
sFWkx6mRWCSFdjHwkosQz2IFdQ6i4+zCzZpzYlEJ4Mv0tzsjPV53rddhnaEnnLVr
KiHtgrobEph97m+zHSqFZU61bLbtWK0dF+vUh2MAqTGQeF5p6tL/GIT2enQDMSXj
Sc0G/wSylbe5rlsMnrVXYtUwfMWYbPP7lgp7EMGj22A6bESQatpMhfbAlt8y0hAq
NsbRS1GVKraF47S4RIP9Oe128eZFEsaxHF9aLUWxpL0p80oHBxheUbtUBZQ0wE6u
BbBy/UR2ZZJPodAXlA50dJqKy1riscgVa6gvAEmxBFux1RRIc5CBtfcj0DBBDvmK
AXbwmtA3090c8ZmKvGLKhZHYywAW4dA+mRkloBru8w/CTaSSLtH90a86n9XRN6vK
Y8kBtelhmAIrvb+Jx3Ej8elOjmMRY61Q/nyRHG5NAtUGGQ0+uC44BM1SkrSyBexX
1uQPHzMw9RIfbB/OnG88t0H99itY/cuUCfDAcbT9MT4KUst0i8Nqk8UHHQNcArXu
M1YPmlGEOHj42yWbAZ+hzSpepDMywBc5GTCcv4CIGCF4aeHRswW05NL213Ondfd5
OTWvH2qdrMunr+3jQFkfZUm2JKO0LttBJzvCJHJ2P8QwIK+LWlVye1B9qdYlPFOT
wDrMGBnqWP8HJCGe/Hy3/kl5ifH+l2AFRgA5aVNM+0hfn3ulD+lg6NUIaWizwXrO
gKmljWzSo8miw+LsaDef6WY1dExx3RwcXG91X2WRxS/6UlB76nWTnD7Nx4yh0SOl
HmzwtUhfZUcEIxkhzTWpRr8Uu70/YcCweamZPQfnV6uCH0cnad/F/qOMEX0OhJH9
SJAZJEsDuJuaKXDQs3s7E6fahaxlL+u0gCoTfUNH+am9ku0K2TeH5hWhSDJqnLB2
Yxw/JMp3IAbCqoxySRrGf0ELGpqBSCDAOZ8Ib59IVTOcObxFs3aXB05m+bzYCTKJ
1Va5y7DmNhzHKpwS/Oc8rujSGN7reZsLOUR0Ujg2AKO2h9+RBb1r6Nc7dKZX5xgD
UTo+UszvuEbgHKVrz5kiPuAQETxGRbl1uWPyagH5lVs6QqlZ4e7h01vCAQRwlRTc
BMLbwmppKP2dbhvPjwuBd8LHUcIluPXE8cFC3DJMPbBuH23BpwSllyDnxNYZUWIt
qapn5k5KdPg+ZVRGsRKUVGvLa0G6y2VvUmIiroVdvgKc0L3D8KKwyt/Nr17qWKh8
wb3SXw+FPFnC2Ev9mTaGgavDpqkyx0xK53Ch4DF6sXeB7BdxD7p91eXlwWWFgkqw
44LHRNQHCeaUzrB+r5RebEMgxV+Xioj3TM1nqELQSELEGc/qiyp4nDNv3bFYUuOk
Qro/uPkZwZQErmoWXyviuuWuDky9YfkrdNjYO0GCFOzvmUf5ZdbNahvycy8IH1HF
YQyw6Bh8rWeDuONcco2GtWJ9eK5LXXAGSXoIAbbPsAHsGd0OsqCgueLPYdZtqQhq
2S0alTpP1OudX2eL27vJfzA7Zm0UXJ5RbM+zJseoibD1IpJx2BHfg83XF83XazAz
a1dOJt+K5sq2mV+DYM64yv7xMohB2sHAfH6+RyYj8RVDROaEeiOwanugRXlyFe6X
FJ3/ZHsDtCtcdi8BVw8q42MRpOaugwCHwYKbMP/m4eXbiRdMu6esAIzgmULlJjPn
ESX3Oj2zmczIjg/aZnP0KyUXtWQSVzthcDD3tAQGpI/NIlA8dEhHDZF+pbyl8Iod
YoFIGrDRJnIQP85EggRvKFD/53TbMu2uBClxL8N3KimSVEJXCC8kAOZzk/XdVzQG
6oupIPsOPCu6+jI0FAzSzN0DhSHqIMjDZO3X6UYMXlesSsr5eVCJsw77+Wdj8sWK
bS7xWrWpYWGemF1uhIF+ebEGFuI/AZm4fwdRuFcJBiBuCrVzDTee7hhH4rioyqUk
l7SNto4slXbFb6lPWjqVpcf2bkODtq/9mmBz1qyKVkh/EKNKd+YnUFqkHkWki/ot
PL3BVH+9fatzNyfz0sm9dk5fOQovPg5C+e0H/6t+QvtT6Z0V1adoEqaC+N6162ju
97b3YVQa5rt2ypTrj7nE+tQS9SXGK6wmqaU/M9b8C0jvfXPIL3l+1/7bSsZ3mR/z
jiSw/7XOlsKV8Kfecm2d7GisCSU2W+B991//L687zjAGY6DypJoB/VFWMo3kmh4F
Cr8kmXoXPpPYBoUvyllok+xapQSEqM45oBX2gTirbZ/7ktLbDGJnegReWctS1i2g
bnUJb4WF5hS39zCpEUuR4By/3zNd11+iAgKCkKtKX5MSGweqDYEzEwGVoMcJ7nob
OjN2XG/vzQR/FtVcNZy0kjhG+2zethjzAAEC3BGkoqUY65IN3QEMwcBtYPU58zGu
Qus1cV4UbmqUull7fghRqKGU+oyN/kEis38uO6eWpjG1csOvF6HqUw8uz0CpJskX
IVaV6F26ifeolep+ghGYCan53/ib/cbj/RwtmxbBtFPsSNKX6QhCZhDiOd7JuK/L
ad/aWdiuxINqQ4fJiS5NPXBjGKOZX70kqyzu+SNluIjRYt9+qQe282qeATGTVUwR
zRYauBwvOLFceI6iPzWBUWisIIxJt392H8KJteBzi8smayVm5lOOIQRt5aLVlgYW
vsBccbdhRxBhFPGl2aeLZ98ETOHUbYu/6MPls7d/HpVsS9ToUc/XNEfp5biEKQ8u
Vu7IfmC73FTN6BYPbIcdW3Xvr8RajWoQ8YjwbxdVt7Qyj0vGE9B6s0YJ+goER2lf
2RpP400P1Zx7Vtivu4cUAdieA+IoUuM889BGfrDaBMHHm1356YEJl6zJFmxIfJtz
cIDYiVLc7y7XNiU7WgI98gk1Rq60YMACtWB1nHpBtvGcuK81Dd1KlMlZKXb89v3Y
Lmj7ZuRWiE0E/q9/Mo6kapkbmAgkJO7b4buRQ9ix5Ew3NlCJg7NZE/WZP8in3qNe
eqAJ6QGRulHn6OqEGveUpw9EM07GECNg/n2CqyvRPCYbdTYjY2IldYlG1rMkt6o+
3ztNps4ytqiljde36w8454OO/Sjv06AsexDtRdpUOgpC7j20R+JPqaFNgFqBKaOz
feGnVyFOlvXMJgx/1fGAkQ0VThYjq4kk2sWWRACx6CYYdIYiBDwm104OENMvoBtv
u3EmwyJx9DaVajXwjK5cJ8nfWMW5X3lkJi0dlxF8fafeiIqvzCihhmTj6gz1D+KT
yxeA93AyoI/qnEJWK2Nhw9HTotyujTO7LAl5q4/A10gFv6jmzjiEGEYOySyEuEse
Ts3AuWN9mIBLgda2X37zgKZxY+arBjb2lEAShGkzlzJSeuabIRmCAOFJVPwVdz1m
GfGGVoLlnWIiU6aUDUiBd7VRSLv70ikoblx9mCdPAtpnkZ3gMqXBwyI/a8s5vu+C
JATMQxJcxWjvMNEJJebRnV03u6t1/TWW/orlXM9kRrKoc63+ZgwTg5pAsjqAJj74
0lxcsf0DdWWoaVoxjdninpw8JklaOqS+FaPdmTM3h5IVATYo2yyn15zbtmcOd0q1
HZueVu+5pkKFuJs/Wjbvxp7HG/SJP6zxKHrzYVQUWCpt3TjAZlJPR3F2pbju1R/L
vkX/IGeqld4k2u1TvQbLXYRB7P+Lu7Hs2JyVpoROuQuopJm0lbud7whrunq1KI+u
jpuyvYfcy7O4/m0AYK/dP6E4bfq9wTn7wASrzYosC55KOQfOTntTCiLPPPUJSDjg
4mePpLepomkH1/RotIn4aT5ZLg2+KlmJ+2U/iEdJmnIgNyPPBq26aN1KT5YELif7
ZZ86PXpCSTkcqsTcRwbal7OA3eHCgJu5QYHAdYyeEmXqLjVU55d9gDA/kqNCT18g
kcAIh8i8CJP1mjsdd+SkkJyjXlMbrcF3aBlVYbL/A+Yi6U0TAx8aCJlRkAtm+BYA
VpYVPgsahOtjsyqtDIZX3yhotg8320BEo9rd6C+BYp/zV4wyeUqvmqzstDhRYvLF
hsej0tjYmmSwWvYTRlOeViGZxDZyMqA0gd+aU4ioNC8KDTP/RwivU42N9CKViXQH
YtlyAUBrY4ljkV1Y1TZ8/vkiWv69r0drAx+U7N5niCB0Ul37dQZ4Vv7rbghnXMRc
KG07Gw6MPMrfgpjsImQH+jl8gHecjo+x/xWPzYsThUKtbcekgn8YkfadFa2Z/flY
Hxg/XbDpzgWbu1u1zorSzx2LKj71TQ74hec+e0lnIPdqJtiGseKblcGyCdkH3MWA
OGcSaRuv9C8bmTAxHBriMGpWNZrwcpA/4D8V4HK7SUY7XXYKLAYB9r/24r0JkjWe
+cW8n6P6pImQnMudmyFhnx7aLo8R6Na7uqMxUNfmuVs9g4LJhJDbjblndcgdP/Sf
flT+VsIN0OGVWuudNHfjgkeZRGgrAolr0FLmNIo3fHTnpkh8t+E+xf1eqjg9ZrKM
/zWzf60a3UcfWc6diAE8fQ8tq4g/0QYHzfncgm2tK4ykzj2kPfL8lmAIIYxIelh6
67DCl/hlL7hzw3Fhw0lULPfT0ZhXKgLiQiTdXsdmVs8S7+8+BeKzbdv4jHKlEjjW
dW2j/AU5V8QNoRMaLN8TnszEdPw679Jo6WToJeyxrsf+Md3TeZq0SRRbJj++JyFg
QnfmrRc3k2+SRs6ee0OK+wQr9djaXNGTM0FjB1Z7odoK5ds9aRz7cipg/4ELN6lR
dqvhSIAgw9GWKHWJjTk60tyFk6QShBfLOCjHMfGqu8JY7ysqagOXwPy+jGyhZShs
/KB1KHVrz1fnc34WeXM/M2BwtprJJyeD035bVZ6eMRpiUTq2rYLrJEo92SLj/6qc
rNXgS7WLQgNcvDnm3O6Pp//Z8S2WLIErwfFrPH4gGSkFGnwXz3C7joQ1Onb30Zul
SlFPiDTxEQzHdW0SBEpkg7ATVwHrbLBQ+zYgK3/ZgSjIRqJvbuwqxr7l+2YA5cib
nZPMFGNqqYLCkKmjgt1BWiD/kJHUn6v0OlQy/RHXie9Ly7uoo72mn/QQJMGim8kR
CoMK6g6PoDOTXIvoeaq5/7+kASlqgW3pXlYiw6ykZqVIwxEacmxRHjUvO8yehWZZ
XVcUlJ4Qeo5/1aKodZcSGYxLbcvtOGje1vJYb9NtuOKp7P4e9bY/cnKnfr40c4N7
aTC/d4/f3Q3Ep1FlTYMF9KZ0fuzUOTDEjaa8zRaT2p7UBHg1/UCANsqa1limt8dq
nRj9gQGnQuWFrWxp6gEHae95gYVcJtViMZi+avWrydqkgpEcKaJV1OgJYYW6zl8v
POrJtCGqb4i7RWglLpBsow/15jZFcIoMtogVhQ8iSf55H1iAzJBZRDCOD07gwxTa
oYIDw3YKruw2qnOFgaeRr2EZn6nu89mdlBUrXp+l6XcNrToeDAkGA2+6THr9v4BW
IQWsgPbwEKqRtW2EKGCptFSYLE1KgjN3/4pESajETmGXYkC+4JoJ1bQdnYo42+dq
ogSoYLS+jaWxEzIO4efFmGewJ58puxaiB0fjXYJx2IKo/D0Loj9V9F6Yg5VHLZat
x7SZEe0w/IkTKFBNlJvgHGQ/k+ESn/VvWcL6jKVkNwV2tL3iEEBDYXGt4lgHTxNw
VxSDDsvgXS2f8xXGsN59MH6/jTBGRiaD6vmh1QTEVa4K/IbmrL+Tu6OSA3UgjvlE
LwNYzb3nCOJxVyQq05iYYw3iRjx4P5VL0UuCpf0D99joeiv2zUFbJEZxkQSDfujA
2tETw4G66gCNF45gO90vvi0UjH2Hl0V6Cxhzq5ziuE1Z3YhdvWU6NL0vbLGE/I/S
cNTBdegeNCb6+LAxjAk6oGhjDNnfdjz5BgCR3nlV8sKqA5t0sjFYpyXiXuQOHcEI
CDdE40CxdHIA+kp+dZSznpU6U24fsSaqupfYoJX2J+5bU2P3g+1XfnaFgrqeyIGu
/nALKdxXciHwOqmt1MNYqmFz3mch1SKDOeXTIw4fbC4tv1AN+opSxoWvqbaaQrOr
q1aDuw02qK4ooB2On67dpjR7tQKNhbJODgLOGgx5KgfmK50MHNyMg7X/19PEKs/W
3XLSI4nYoeG6ohzQ4gkM5ffcSnFQ+3tEkwq4kq+qS1BOGVTobfFtJNRvPz65pufT
LDu64CxmLHHmRDTlvWVFvOf35g8RwxxBwSs0cWAb/NtkCHdw6y/JX/lE+6e5Yvzf
luh4QHt5i17VIE4k9yXx+zn9a4QsWpFlgnaCFuStAsjFbwmAnd34J4yCBMDt3jJs
tdp6oHx9dtWX4+BQuiOL5KRfg1GGRlgLiCSJzEn0ILyfJ6BfLRcTgr/TUwF0ALP5
CBLhReBhQ2I7WtqFi2aBDpQHy7zCIg2UJyzjf4WD+W4zPSkMNqMSaP5neZoofhbC
RQtWLsgjfVTjvnpDhoQUFkFGDpHUbLnX3OAWUdp4iVbeHY2HAI30ZtFMQ269QVZ6
v57NzMYTp1+NkZH2H2gRUmy0wEivKX48zss/Oi7QpaKwBckZBDWGS+Eo4+A4ZybC
far0/6jMaFBQOPCdVtAvjTZzwN45DNMIIiN+a3Pt2kX5YD8pFn0mrrorlJGYdi6u
4y3p/CNYJgNhF43vw4ZoINK7XHCjgj5H9pBGlXglCWrx2NS1Hjz6QUTEuU5DWSKZ
W18NPH532GPeC0Y1dStCaWYnaNxBZN5GpRqsOQnxO17G9ddK2LtUqDJiis27Xukb
v6aqFdH75O7qi7nRchn32Y6mBM6MU45j1pESniZ4Vll4CAqEPMBTEC8JLoEv/e1e
tnIO3/yuhpeza9ubfzAtG29cVB1vMYhjBX5o78nYWO0gj8QQNCKG3xz68/gnmt0N
xqR3d0nuva+IKwSeNhNLJkXrz0lVvAdtmIY4lpvl7cCloDSMJ1oBNDoFrI4QaojN
mk8d6Q7ez6UCKib7jBUoxyb8hW7lMjnUF54ip507jYAhb3RkGBAbuhZTrenOcZ3b
1wvi2aONgxrdUM1VAqWvPRqi1wL+SOCb/PeVfwcNBdaMwTfXUE3MGp4RQ9THH3S8
kgzmNu4BmqvCkVz2OaRxgGEk787JfCi45vjVZ3h/pI7iaTtdst7Bh6eebdT80mDJ
BIiUWwnVz5RPNgQ7YnnRAb7C4VfFDHVXLyk925D159ghaN6AbMY+Zzwohxbqrcjv
5kGpWLXqAmJtQ3DchIH2xPsGsnJrsbKY7co6fvwL4av7l0TEmu/chnwacjyhpZOp
ro7KyaoFEbBCd5vcrAma6xBqeE3cYttXsVYEisJSClTEDCeDuDroM0rAcysq4UJV
K8OaYL7xKnWdkkXDk3BV9whfCUfq3NW6s46YFRYKb63fBTcbNikhXjt8OyZJWkZZ
fqgkRSi6mswfUleN0pwmUgjL6zIXRrKzGYO17Mm/L5FRA88cZkEwwlH13l1VuaCp
lEo4Yde0ewBiagqQrM/qlMvjGGMLLppHcqpamx+Wp+mvRKXMQHyuWa5t7NLaJ4iS
RTdMI9wXZaAs5n7CIMFCo1yx3wUwaX4VwSpAs5gtAsHSlCeYi2d4eYASYKcAc8ob
CsKjkbL2gSsJ52vqEPpM6SwJgMqcsJmV973a233F34PFqnhxaOOjAXd11LeZtEom
y/xe11XmzRXyiRcvEsjDgalg108Q9cQ1yMrdaP2Lx3iPq6XGAKlUq3e3A7wAlkNZ
Zm1vrZuYxIhf8wlKSO59M9Wot8hVNdmLz+S+4jPgWetYxHWVjcPyl1bp+yY2WVEH
nH1CwRMFTtKyUPxDPItOCoZ8Cx7sssIqWL5yqY+TDznArTLON6O9nktZcDiBEQ/n
th3n0E/iz0OfioTZTc+wtoCDRc2i/jxThmIx4nADKzd4b8trfoUbHm7ky9Pqn9Ej
EThDYBPA4ExDVk2HSbZfK0LKmvYRItUZUAdi3mNZP/9GbZxt0EsQ9cDY+VuGdT8Y
X8GdkhaTq+fmzt7mgr6uvsKuQumGMxb3yF6IDlBbCogphH8jvtrFydV5EQulclIq
cxljG6k2f69br8GgyLeBodjae3uPObx/89cfT/KyqUe7iEptxBQbGQjQ/x/9ilzt
zCD95v0VavJgVDyVv29zhpWKwdC1YOY3zo3TYRY5sl41wJRTGrS/uOVj/Xex7mix
RaiL1JTBqOBoCPpIZ1JE29Awuvmkb5dMvjMdNMj+5BkqZOtQMcswMTnVB097L8vQ
oXKbJ0mRcg97a6rOgNtBz4iBUVKqMJ9cSKjyHsxXamBNnnBoQSCXWTdi6iYQ249K
DnENzuWG3u1UL9baRyjUygwA+RmieNpruv9JhqTDBe3gi8JngJ4Mb155ndZCdNM8
5INE9ZQdIOB3zDW/vZrrfFBaFujNUF+C6gctzDc626ac2C6V5dfLCf48FQonMnAp
nXdCr/AEo8E/h6d+foOl8TWubSM+1t9yENHAY+ADcQdCs6g+dO5TX4BQYi2VUcto
1Zd24xSybDhkERWjKZF6qUlHxLAzmY3XEIbI+HyZXG4/wEOR9mYnqyj50QUCmlP4
qNCusDFXP/v+gZCTgGKcgAjDNlkD4qggYVPoiY4JEdysd4bDUBqgs24Mhg50N3Bn
soXOWm2cQ6qOZ+/j1hY4xKuYk5aoPN/dnhxQlSiY5i1I4Et7jmjIcPjZQYjIFtDW
CDFk2TKZGv/XRnY62ptueAV0m3FXyPLgKtXdsBi+QiSnV+SEUH+/FO+zcO/6rp2R
i4bis1iebjraRDBQMdMgMH4DbowIxBUBOkfl9+UxCC4UtIDEXkDgFS4G/iQdS8ur
5t+sLCfkf0IbaJE37VjBI4fzQ7yQOzAPLWQponuBfgUlhHnqvu4ED8jWfsCK3f2o
UXyjKnvyY0PkuLCALyl2gDRRkvewBodHeVj89NxH+Rw5JHcIjk6hE/tQsZZ58Fl7
mAvf64vGL5/IZyoQo/8hpCpT88DYXYMXuGmklru/CAPmgupax+uL5pGowD7AgQrf
VOmlwKpHAU8ewFiekXGwRJz9CsmUL3YhM5Njsf4s8T3xHI/PEnmx7ciaGJJPTO5Z
ZOPsbPe5lSYbcWbhDBrqpHQX+PZaAlmEJkihB0m4tqVYnJacUv+i8UPLwThjBXaX
Nxuwqn980VtrA08Bq6Dv5pVDnfVB2/+BNJcx0I4fuN9ntDScyqrKAn08fBKVwJ8+
ta6EQPDQI+je0mWeXrcoOHRv1lHxFZhnllnJNOlTP0YO2sqV8Q2+fIwQOtFxIXPk
dm/kQCnxEe8qQFIsE2vgguiMmDjcUF9aIoburQngDoqivbcw9AMdTJ+uCX/bRowf
ATZAM63rClZ6pxJyLyro+tW1lfYWIKs73FkYVavg0zntf5P/hzkHwp2GAC2G5Lk0
TT3iOdnzj9el8eSD0XFIIm5v3FQrxobTWi3z8B0LitEAAqYLxDwXJC4Xypt4OXct
2eDXrIjccp8deRKLAANKl/ywNQETtkU+q9u75+tb/W0j1ivkcoz0YhSDiaH7agma
rdzBO3G4PnCRnAd5yOpJCWli5kThebMDMqVeC4sXl6s3BWeH8dA9RVUk06kvHlXs
/I4xzKE+Wdzkv16CXwFjYUULXSKnt7+gOMn/qi15++y1Z9bVDQZmwbZD3N06Abkc
JSBnf7kUGcP3Rvz+BWXYo1J5SgrcNfeoK1ifUuDXRY6xUXQqCmz+Z7DidwBIt5t0
Yum4pkjAMqq9E1TWNaNV6LS+VrGoOpcS8SV72CucekmDgoeMBp7eI41CKsMabaB3
2RACajLiU+4P1HX7sN2lEV/TQW5DisbSN5J46gURBC4vqkthn27VLu5DDBLyd3ac
toYJcaUSpm/edVZ7dUtKTQ9mus2YblN5NW7awKuABakXh17rK0TLuu1O94yI8CNn
cjSDHoaJLKuuVZxdYeboXl/gUC3zS9KkgpxVNu1nwQx7r16pom3P5ZP4Mg8lzvi7
Ti56xv3ThT2y3J1l/NTYpHhSpULvG9GzfpTdVLpLQbCjLzAfC9pYYjucyb3yPlsg
hBXbGSXFDHLbbSVlT2kFif5RT1zqVTiEGyDG17gvSyQipZingSHkm3A+OMPMETsH
ftBIi8le7B/M+kdV/Eg2tswUnkuJpKz003145ItuktrXHVQrcFsDI/Q6TLXRSL+b
BG3WCzorcBKWwrYGGkByxk8opnZw3g22nE9FgQUm5yZXjela6pXTT/mO1uLUMBim
od0op3IbYUT7O2FrpUQqfREbJ/n0r0N1HjqDhlyE/auJhDAoQVbELEFXYnyuhPPE
oGBaimUXHXA444bafSLi/wtifev4LJ9eECDRDSQK6EwybCpXKryGFNPaysP3h0J7
z3YNe30M8A7+yIKIOih8gSzRgI6jrCdwhtPmNS9iFmyutI6DmKjnKk/CNsUn/XL2
Hv/7/WiRfQzhdyBQTAK6hr8kX9BY9E07dfNHQ7ghWZYNLdHA1OuuH3ie/HINANmj
lEweAS/8MtBGNtKkMcqgYmfvT9eYmQoaW+prbcVo7wqxPdtyy0D+kb/UbbEBrtoU
XsQDFsPAPluEaND/cED0znJkoGR/UBzSxSMvJlkNa3vff0IJa7CT5s3bYC3Qe9NE
RXhb1V6yGH1ymab2KpiyMYuY0g6Mp7PL5VBpVbFHpHIBdR07mRto4u1jjkHTea70
x8tF2mhnTS8MwvTNA5zBi1FOtgOv8rKQSMOZNRwywRfh6ASthZBrvIxzmyFHMv27
EVgCiB81wkUnf5OzRBC/NXvTFLZiaqCperKIw56OA0RVkSy3pkBiYeDrAraXx1L6
m01u5JKdLlbQypCiFLUON4lemgpshcHF13SxVwCD+62g3sbMul//b9BQZaB+AqPc
llPouL7NhK8lw2I0q8A30TM08RsILR0T4bTKhde8hHuue2Y3PVHP3AZ8Mr3y47Bx
zCXKOV6llMmFevNwE6FqK+C4ZudprtH9GKxA77yriTZ3Cjw3uzR+caVvN0Vq6r0r
vmX2/T45yECFwko6n6sfN9R7pqgKttn0iDqEs+7b92qmrDP0v3pJaTlX8A5pAAxk
bU7Wd7f2MSVOuewh2ZFsfoMaEfUh4g5EAi8+gH8OpPaznkE8xzT/kYsvr+1TaFLV
gppf0olrLLR0fU0kl/XlHJxasKC8qWTBKZxxu1Mub09jGG+jgkqXvp5M/CASp9oz
HTL2DXnkwJ6CeGOd7fFQjIpSzwnD6x4ZnaP0ZKekkSmDZq73GDp6gOXiO3/gcjTv
H9t1susEWVsu57k3z7UGYfJEairssYlmbExfqPDkBPnMPI46mV5dr4Kmy4RszoUf
UJGC1nSSSX7QQSLDxE2JjpQpfHcIbEh9guTjoRZc5JM6e5VuDnIq/aALOOpF9Dgz
AFQ5GJmerwEtZ6LY54wMAtLrwCB25frOMBa8rbDPOI1I0zzrpiOfb1MpGit+SDal
1gLfIhF4KmPOLCIq2pG0Kj40C4GU6sPkhDoyNwE2+4f20CLPOG6s6y11zwnfmxxS
TGLajiSgbPDO1tlniyt2Jq3/NNq91QFYkEdFZ2R/5h9HE6irWlGVWsWKgrJ5ggZs
6MQV8nBD2RqcJ9lI75xPMhRl4g34Jg06BeupNdOr3EKxYlzW1icoPLzDSudd4aVl
yFA0AOH+DX8fmiMA1o7dtBYX+HvS4s6MQKkq10H1HgjDPnh84DzcHqr+SHi30xXV
qk588MqxlJt8jeRwwR2HdUy0QAuM9mxFNZyQAOI0bUgruwdX8NVpfU2JLdIIvQVU
pr9/OU8I3CkuPc47jJkttLL8002Q1v8Uf9KVAgcu4Mh96xS2Wv9yatyjf3u72vkI
nWWOUcRnfV2UOu/1B2hiLOdACl62OTYCig8D9uGLkkt4wSIn08LnKRItOr5iyuGg
fjZrpZcVmAqNeyCPNgW3mXpxUbkl7v/KRmDuNYQE5uk9TTaOl6h3cwaIWqjh0FSV
Cnab36VpE65BnYKOAlylLQzFv/TTgxebDi22R4f0BSciwIlqbCxyyAtUyDPfCILq
EeTuDf4uZvDg+M8F5ZvK2Tqwb3NV7wzSsMrEYgWH8Fr0MBiB/k9hqv6TK9JVPfKB
sPOXbV9oKkZ8YkG3kXFYHmnVW7JPoiyFAf6U+i0QiI8uEg/dIalIhToQaSkH9/6l
0P7Re37EY8N1j5yhYh7mLzPKE+C/AXLqFqjZ2cBm9gvQNrE++H9uxYerHJpn5hiJ
y024/PywPvnx8oKAKlfqyoI3qtEzynKIURD1+hcOlgQtudUeyuhWTaL6fp7HTFml
d469uw+TWXuckJXZBbkCWDM/q1Kq+R6W8jWH3BhJaQgk4zFqgFfKT3EFWl0Idr6c
aqLy+zONQFBSWkP1DV9nifQKAbSeVdWpAgWkdZKZBiSq6Z6C0lX0Rsn3NfnGz2Zm
i/L8NtU7RkMwQIYENJXvXmDMo/qn6dG9gzBYx5thjeN29QYn3rT5q71ZYvofhC8W
fCdCuo3xLJfr6uuAOwMpEsd6gN4QNkSEkzD2uASoGpnbCxvUhwxSAnEBrunm2U/M
NeBanM+/vcdY80sYr32Q5KRsHYc3UaMmPyB6JCztyLKSkPFrcZJo8QIQG3HOUDTw
m/gt9223pYngyU2/TRtSB/8Ki+onWRc2NLWwPnfRsrIFN5s3VCJu8XCiOjZuzm9U
CYRU1VJnQxRnHkdo/lGyHTaCaQYYAaP7A+BEVPKxgOfmpd5HPRNmaCFsBICFPFZi
UzbV26fyEEjnItlfTLISNFMp2rbxRjNBv/ebcUVr/UMfmiXQneljjWVEoQRQb95a
nQ59kp81S9xH/KDYfjKeFHMWSdIYQ3X/FEGvak/cw4TQsLVziYj8L9ZZ1IjBrHZo
jzTJ816wRPlg2YP+n0dHSQKakSLuvu/UHVh1vjvJsH5ZB11tpoxkYYwhx2Al+T+J
S2lZ5/VAqfMTJ0QqOP9adRQ+zkM01bxIpxGhctRTYXI/PnJ89vWTSWexRZULEIat
bNeVq5Fezp1prn6/Uwm3HUf+vUca2T+ToqLRadG3zEJjYTYUHtUQRnP375atCEe4
+zO6edOFhRkRJZ74oNGUJUxs2J0d8zIyQPgYywFQv2VqbjRs5KxfSRqTtduH8xg6
P/C2Roir5GiqMPdTd/VqdHp/7z6K+VmJ3crKK/pYCOqOC0vqnNIpWUT7YXDJ9OlC
oKq8UWRiftiCwHnQfGO6mhsjuCzpuVhJu4TqLJPnZ8O2sXC6rFW/xHYcuCGww9lJ
NmzkMDzaFruB1dopEu8e5ZzLrKvPCcOB+jRASVRHBPE/Lox+gm/cYbzqewjTj6vF
VKeqm+zZ6zJtnKboJDGJftyXSaiipSJJsLppbuAapVvwU08gHo4AYlErazTX6mJd
qBvi5mriyRpBVmYqR3mxwGPu2eBGFmRRO4mnbn2LbPk8vOypqx3MtVBEhMbK5NN+
yIkWVdV5EEYgMiTJJd29xU2OTz17WH9XYm6EDjl2jzt/DQy1mshvorZZy6F34Dl8
uVJ0rlDuHRmIQD6uf7+IN90WQN8o+z1ASClV+jaohohoRX2MwMtBy71dfBZjh6IC
3Z4h/pvEQTgUqFNRASbsQ954IjCMhMdDGQM4NHRB/LztUGzZ1Ze83NNwlyNTBSDr
CwYvfEwJa+t5RpHhxwUd12MSFKRXnkCTaO4iAkBR1i6uQUWiCPiSFokWC6BCI5Ms
b7vK8BTlgHwQKB2PVLDPhdZNM+FOoutFxDD6ccsXFpfxMDS7ZM9lgbvhkDDvwH/a
aUrSgtoluLUG9bwD3Pu5K9TxRdzdiPXqRPRFnmP2PaUvUwcVOBHVmItxZ2nsID3k
ncwI1BKEI/PQDezGrxSltUY9N41CaunLV/OvfPnGakkXjH/BvdrwxGzP+Yp9p2el
9hzVjVkJGNK1ClKLXdRGr60DO1rocuOeiGx329qCXoIsi+v4CnfdLwHIHAc5e7kP
f2upUqFxELfff1b+I6JgyxtsMASjy7S5rw/lX/h/KJHd9PvisTrm+ebizwOWLLna
V38Y8jvqZ/+i5zBXHsfCgPWw20wNpbmNtZcTPTpgWE7o1S5Dog/MaAQt1Nn5foVl
T+Hm02GLWcKIKKZLCN13GwQ8j8EJKwchgKbmaIPVILLRYGKg4rP6+dDbHpwdKxnY
/DWv4PVHtX7Kb+WOnGF4SfIQ686cupngC0prU602N24bjUZ8qLAMX+4Qr9/q20Pg
WcszJfU5XF3jnlECTXi2FYhXxRBGwuhowseh2QdNKe1ZZJDxZRIH2zP1A07l+jHz
xEsn3EiyG93jfb6h2YXdQ+rSoZqLgnEpuPsiv8nG6zMm4+gr+lKt9A31H6LtE9hg
dfbNmO8PyE+aH095B86pt/udG3Hka0DrOhigA5F4iUoRhPwgKRcwQfnIoxp2azA7
fFbZHlnV8+CtNTocq/n166C0lRJ9bdYkpEhsYyYeNQ45j2tezAifhKmvjmoZ5Fvr
O8rDayvFtC4MfdByBj9ylf1Ye/NW3I/mP52FaM1MH/HK2xQj5l/OWO9HAiKS2dex
7aRtebcKKFHOK4/xU2ML3NgLJO7LnRD+GINvQam8/nKv2vx12ykaLcz5hH5pwis8
aSD7Do+doz79tuu/T2Efaw90pltCxhPiPZB/hheryxBgUqx07RB0R0Sagcg3BBwP
GBM6UaE9CUu8la34mb/4zCfBIHqpertavWO2cg5Pd4oWRh9uKKzc/ufHl5EPSslX
WJscYPQQbY05uWBN9W1UDhHvnDPmQq67oXRolR6JcNDIIQL8QAcTPayi7ve61tZv
4Uk9AvUnd2Wap3hVYw9ew1HNMzJ+jkhbO8XktCsLMFP8OqMOUphijMmCmeKogNRp
OYsOA1IL0Xj+QyoxFq6vC819xijLYXjp8XNPRNUahi8rmVwEXQNQMk9o8hIJVb2f
b3CpwUrp9L7h7cSooak2dQMP2EPFU8F4s5KjjEKZy03oK61O5j0lYLB2TZfvlKHZ
c0RnuJnymwLRxH9ZzjCqSHKLKZ45i5teRtscdGJRw74cUcHlPyi+CAsFrx4EiVli
mWztcoDau/W1lFLUuPO3Z6tg3qmD7ndDfl+opTdH3qqN5XFp1RiKB6/Wq3daTFBd
XFKIgQHVNBtUeBcqdBlGug6aHqO1p3Pu1GPMEnWfZEuA4YtMsfN6DL57Vq6yxgQf
VwLlnZPqAE0rumHCNZfpaoWIAmweTYRO+pfuGlmovyfgrdKjF9kEewrSdtAmBnCk
86fHYfdfczHu0wXw3CPbmtaFe5zvffSM3e+UA1jWLEDOQzwIKMYUm+KndgpGRfh0
UdbrzFZslj3VmJ0wuu/VJE9NOYRPHZbDa9H9KmewibJL2ZKlUyxV6lyAjc+TS1Gi
/a57fLB/euTRG2BZins+TLw7DIrWep9UEvDKy5jOCJPdnyQs7Zy1bd4zHpsDeqto
gGz7afXBuKGrzRD5JWvusefwbXFRgr3B2NAPwgU06bRrr4dRQIS5H4f2Q+HaOP0q
NyjxNcFqDCSapgE9vi/7h44k/gQMNc2gbI+ypl6x7T1FRIlpiP8CUat9taoSXaRX
CMxRov1C21LUmffrlKL/z+II6XKuFdxm/5cs4bUkmP88K664G2svEC1UsLJuhTGz
jxxqHjeGeF0FelNZRDyTuCjKFUTbZLgdLX0aRjXnIAbPWFM2z0gfzrSQgL1ExHNA
cDykZe/s6/hnOYGa9wsrrCbykXye82LYsJMQYdx3X4qwc0UcCkt/LuKo9ilVlbWQ
ClIyrhDdj7lmAZSLwLHhPfjqmZt/x7z3+i+b/gsDZQXnQW2m7TQ0ZtaiWhNrL3mH
Lzk61pZwT8q98NEPJIOb2E7ki1ZkLPLxW8NjC2DMUPWENBQgQniK7BF4qpmq3mz/
pN9SKYgaAceeu1EvrcPUQJWJXBYtdz3KHrtL47an2OkcUsVvPFf4jX/zg1fp29nb
Ax5/pJByrVE3JgklmN0Krb2WRmMU7LokEIbpjS261Mj/VsCYUWVmZbIwd7RK6ZqX
P7OC5NhzSsugRF/7bgiJ9m0AnKgdKOscZKXjvmc7olU+TNXRniOL73cly7uiU7bA
oVI647C2ZY1wxgoSfcFuRpEi34X4pbIXtp/XrOmWvYAB9jPhxg1vluj1TfpLfkPR
yOsU4E3aEASoG7wgh763HJyv8ogcXfxlwG3ysqP2nx23gA/8l+RS3XFl1lbHu8BQ
jYc8luzoFK1LfI/mfz056YklZX3Z1/Y6Lmr0B9mMn4ZJIJR+AJwUcAJ+2L8Hme2W
OFrHRKaJiQhjCTizkbFDIHODWX6hcNw/w1Vm9WN7DHTjU6OOMA3jNFzr/gg+Hxea
YM0pJ5qlg967k3QYtcvGoaePiSbTQaw2xmwwj198c28IHn+2rK4SeEeDBj5ZwFwR
RrssN8iY13A8zldcvIGznGkU6wtZbQoGVzvwjSL0azQ3tgZ6Ig8Cbyr7phTYjeuL
Fyxp8e0s66UeoHgeshJSl3ykfwiEkfgr0sJ/Uhz89lJT2Cx2PhX7JPmrQ5k9IMtx
uwmnWh/Rkh6McPG8idYx5ghGaWWt7UnXSvYDvCNeCQ2X9JwXynp5pgk3D45p5oXv
+UqJPxNHorJPwu1grlh0ZRb9JWdGxqfOinYoWiNEJS5QXxZ9mrNQaBRGAuVJFgiR
v7baR3aodTPZfHOKG1mfB5sk1NYz3WDJ2gfe/JLKqy2cMKjb7zYKYDhiyapq3Rot
idG5ZhX4UlZONF8a7VFu6rlidkRsWTqyf4t7FrXaILs1MVJ3gzWyu1cqFwLk9kKI
dwf5nbKc4dbPYVPK9TIiXyQqkf+0078wbPS1HCPbHCzVoVRBdzyJdudHzcLG44JI
d7gGe9p4kOLghr/d5SsnLvuDHEY5aHwQu/HTYEx8lPxRySPg/9AyodUxkMLWrmz/
jHaQsyCDnS62H4wZqkTMpvN5A6upDPvruq9ejUPoSK7FtiRrz2VoHcIOMiojYABc
omiylul/0Uv/CP+5MaX9Qj1JTVQyaqYrkadzpfwsijGMasgvyxtCgH1lYPVfrCOz
zIl98yspiXGDb90l0vN7XvmU9Nlz2Ls9F7QAoT9ucEIwxklUi7MC1PVmjggUJTtt
KOmHH92szKGOBHW+3ms+VVO34NUqWHx3esvic4J3CopNuJ/yulyAMwTkDW6Gz5Q4
Qh1DwPmXY4MGzpggrSBeGKI/NiHpkSIvRMTz4HY/u9/hWfx2Ab6ePDerxvyhsQu9
I2TbdfR6tKDb/HnDz2GJJ6pP3W8zAc4B/WVFXQjqrKqRIJ/gmeEsIYrX1/ACGLF1
PiA2MhNIfI/lN9QZu79L1G9smF7OoH0N60I5jUFjodDxpH37cFR009lP9J4pY+JB
ZNzXMsqOuUCyMNwP20/WjQL/ejzDgNwcPeju1KR5nIuoYcPt00WoGap+2KLFisyL
+Sh7cFbAndsfVtm82ASrS+DR+0e0bp+vgAcEWU+01ROvvksGSdYTRKF2+08i/Wqz
SWY9YjOrYJ/SHTBmTaG45OZJw/e+Tv5SKeCRtki4IVP2PboThszEwGJAaiVJtMG9
BWRFQ14rtNR/yjWsyUvVjFTk6LZTWHueRKXH1HnAR/YkCEH7+Cj5RfB6YK6pEbGS
irjXfDJ6TvMQjhIz6RKA7lrTPWmeruqR3kJ5Ns7FrlznQHzZ270fcHFU6je5YSOX
aj5WUwzl+UI48H3kSIo7A+CR6QxH9pZGor00h315vLkET+BQDvs2Ux734coBJ5xD
RDzyi22bFba1kdolQ0W33QXKyRjQ0ZamE2/bPcGBiDxcxrUlQtwMVrc7TwdSmIct
hZe6YOL40Eac9DGDQI5f7H5RWENHfI51RED3nETncl1KvtcQvr6HecCW8dYWaOR7
khXYhL6C9dqIkLYdCQeLptfjLir3AxcOLuT33RKXDV0ebQKe2u7Ez2VXNBcoFedh
HtEwGb/wuHE6b/tY0PS9DFz3dL1WpKBtIOHfwkexDoGUAX7sWQmKmD4qPglDolyV
IXOWtv614V6BBn/l/T5m62XJZqjJySH9fgHOdtQRP8deO2/kM8S5/YOjPKa3jC/R
9NQtilt6GvA76gT+2Qm+HWqVwfdrb2iz0mYQTm/GGMId3vJ/W83vLCd5u5N6S4sS
9ACUVV8jAJEkUMpeLvVy1vDvzoqCPIF9jxcRCi1a0YfpnmG8AiNbTs3ogA1cTZfJ
LQEkem2LZuC2eOJX/3S0AgvBYdVOzC+iHAq0QfUgtHBBtT30hwENj284Q2IKvvLL
0hahKpWTfm6wTYwjvIySh1vDAaS18F3S73iXZ6cfsAszt7FmnyNwz+Oiddvkx92B
Qz8I2jk5WGT91l0NuUA7EUYmPZ3liTi3cEEoLHjpsBB6KQAV5eB5l41fOCtIdHPF
NjTbuk8wyQQ6Ma6OF5g1NjgoVep/JnN3Wqp5j/AxPaZueCuFRF6ve4blbAnXlYGV
1rD/6Mb+ecTzAKCxaJxd5H8C/Xvgbzaq5HirWfWsWz80NJvi8g864Zd+rNBYB3yU
jQR2k6KQ6SERQTYH1GV6sVl2G8FGanj2M9ZoXVf/EMkCmn67k3xDX0+nvuGgXXxf
EmTUTre6LaKtPWapuxr0Y/NfVkQdWAWE2qVjCslmsJcCeK6t9cFmSXO+EG49rnZL
DYYd4IbBlQCvy9lDUhPo3J9Tddo4GTcJ/YjSBoCSO35a/mVcIbVDvdpTO2w/coDH
g9mUAN8arELyo8bHHXJsgygX8jSAVdUNVUEiNSqxwnCh5V9wgFVI4k1VUJ6S3f6t
+SctPfuPuhX8QJoHQ6XtJO+DUWqLbL1itn4aSnZM96N2N87YU8P9fzL15l8IYdyZ
fJkG3jFpsb1O1RQQnfqMGqcqpP9RjwDolZyn/paDObnUv6LBHCU6mvhgt+Lplach
XEXNwaibHqxrSUUPk3udBO49nVWJmQYLEvDgkh/FqNgvSqzMEBoYmbOP3y6Ignzb
/uJ+xMtGZxxcPnqlvfG18HSMWNbz49K+Ds5ddLEUMb5n5tsjDj/cbbuURfHuSaNX
l9ZsNIhfX+EAYVLgTlq7arUWbuFBmjSKoSbkBFPQd+CulsKLyW8FpXICAKOUW4Uv
ce3uXej93tizTWHhn/XgykcdZvpUlSdG2IaOP9X8nskHu68db7D4mJwwilX/nIX1
eKa5hbiDLZqVYHAYFi8MkL16+NNP45OWulsvtgB6RYQ2RmpckbuvGM24Q1EaaYVX
bw5rRG5MJxYoewiwazQTsx9xvmf7BZ2hXnUMILlcKhMehjqpDdhjH68o6EnZ76vB
iYFfGk7pLRl+o3M4EyO/YoWtKINSPXyzDA5nFI9qHSXmGFeKQdbZP7/PRyhQXTeD
SiZt/LYtuR76nP8w/CqtQsjzMWxta086pyYtBYz7STom4SFDsEMlWIXal6q2Cf3l
0Fp9iPOepsqIsUCtgyv5+EbebwOGpTD1XuuVtr2tu1G9lazU4Ar3iQLLQ2ugiCKd
CrsXodtqJDkurLQmOTXTBvWYEhdW/dw6j2EhytsHSgixxH5wVD/qztpZT+kEjVRj
6Yn6d8wNmYFknSbIToIzpRyFdprvp+/+y1lJCB10o46PfVv2fRMM8fGId3D92zKF
wUINFABOqyYs5vWGP4VADHlVoqn2d7JDOAoXlUoJ+0YXOtW5SVrkuAOBZVO7GlNX
w8J2peVB5MnLZZ4Ol/5EYT1EpgUbOqjJ2nuKrGYyARuDd20hwr0PI91wmGnchQPY
og4rZMiC/qJTWvDAcDuH+nGKEG5tbWmO/P+oy2Iarpcex2fadF03+ZYkyPIngTQ8
Ous4EWQkFWzAOXK7fsaDf1hecY056FF8qOlWt6Bp4WHHosbwH0mLJySDo0p2wx5i
Uh5pban+yFnoJywDrHgqPyiWYfha1VlZxJnqdEf6UtDmERe/R1WSm/G3BE8pmbLz
6iE+rrGObD6g+4YxjhwY5mm8XBclBbF/mweYNEK/cdFCOAVxhPLJTQNUAEudxWn4
rzexu+dR5kfXB6Y04ywcvhIAWghwRQgghbN3R757C5szpWTjhUJie2msp6qwSb89
/pK6TvYKwNV4sOisrdLYZmNXPGFLHi05dZ+QqtQBsvPXdXq0lbhq5Fu/Sb/+fCel
b7r2SLEUGQs9aF1+WuRWOEOdivLBr/KfWCIxFYsl2h51SIRB0oEtsORcQ2L4d/rX
pZ0LJoPK5rbFYUu0bHKNb0c3XUUK0ez+T7OHGEDmeqo53wRMJwO96SCEJiOOSnpe
29jsASVyU6YIJQtlgX8IIjxKY+Xg8qtYe5vCqgn64WLvw4/2ATP8M4aWsdGCPGkq
3KTl1ZUF3+ZWmwwp8C07jh254KdgSqvyGcthXG/6jOAspwTIzfxk2Owg/XQaKfqi
3FzwwJUF+zdN29lnUMg9c7ivWeQX2hwUgqxicoxONuqWywMNisoy05DUi+VNPc24
fmoyV652QhJ/x+2zQO0zxX8UlDmXWdqse5HTuyCUiP8jGiJIBq1BnlRtV/+Lm254
wK0SkCHO0GOdaSUp5ZVESDNAdvuTC9I0uQZ90m2ubPQgtF5x7dZbxdsZ9QEj7+MV
XNsgtggKVgCfhnG/UKmlI4YhdlIBjNX0vdQZYnDoCw1fGcPktL3CC3HApNZBjMh9
SGG086j1yVA24qMlLWpSMhPqq3hkkV/3n8AFO2R33OvjJFclBOpGT2r1PG4k4/9A
MpsJ2bwi0z+J64HsmULLvHlu1bgJNgmtE8KdPIDauxPqE/YhKBIoj9nM0qlWBMSy
8zHnmgnKSovVOHwHToCEDvpl7xF9NMihJ9X9tWWVQuUnTBPvbvde3VcNCRRgdnHm
nKoUv1VfG7xYPxT4LtKEwSGA03ay+RiuK5otlWW7BexK9RHYsfZKoZK916EjS8Cm
+qbNqBb6ZVB8NSvHHURuluDxnz2Z85lQL0G52q2EeZBcEx3wqqgeqxBzonL9TYFa
mdcziPU6Cln1fTVkn96WwsSKvvL+NIzQ+Ia+txiMU6dhX5+gI5gf5fCxIOmXg/Mt
eST9J1+8sXCp9PncAUrePCzvqYEKnnSWmS72r/tz1FBFhi37dIm7m5PJ7LweZuFA
LQu5XCgwpEhAHPPgx+RrbFXRGxgU4Ccxoz/Az8LkFjzOMWZEJ4SmM9biQTwDdF52
Ik45X8oDyvYCXO3WYQv3nJ8ujXxvW+ZjRv4PEe5Bv0Jwj3hkFd9I34G5zrBIhoMg
+8pPedVUUVKvQWZ+2W6O90cabRf/A8HSoi6eehJeMBcRuYjSfwI3TMt6nzZNp6BL
5KTP4IpFqcZhZAp/DnZuLAMpEzD7EpZiD05SO9C0IYUZiEyJw4skTvuVVqhacMhS
xIYr/fvxCcFLu/1+A4EdRCap9Dw3YRL0nKyDimjzF8eu9hm60m7LpTPmK9k/aLox
TkT2FRyP/3UGKIy0H9Wz38+zcSMr+6BMrdrDuM5BdSICW/o3cqPAQ1/mD0xR/nhQ
CELMKcrKoqzVezhAzaqBFYSMQTLSxD9wa9Aib/3xTOarKsNYchIJ3YR6ezIPb5lU
2slOy0o2BtyPGi0q1qU+LS0aRixPBd9M5TPFHQ8gXQAHuH0WV2pESY9AIigg7vUz
mr1fDwY1eAb3g73l1gh8odFKO/908Krwn9MCOtfA/otpwdXDv1mqKLIa0v/9NPeS
+N7z8EMb3+1FLLg4ENLebVroNcUjeB4lYoNEdwtK/fyhPXJ0Ekt8tSgf2EKqiiRO
tNG9KMQrqUd1783Ctf3JNdW1dCqA0uOre/AFYIwQCJaf7UAXSh6Cf3s4IT762Ebh
xm3bESpqSIz3W8C/qrz9xdX5qPZDBvVLsxlKXeROI+0O8CaJj0J1di0hUYMDpF21
he84afe2/cuWwQCD9Z/3D0x5vo9iIJ5GAv77WSfEZao0j3xp1TLZ+Sffx4dAlIYp
iIBkLZgUPlulys6FwSF4q3HOg/iGF83rF3j07/Bdw5m/e6LHN5NILAIYPX/1TSTO
1GdvrSkwfobp0BioSc22GMngZAcID9zPhzgjybwTUr6f6Y/FrIO6OzG0AaVxqJlf
+zrHebslf7Cc1nUmZdb7O6l/jslTKb7MeDzI7mJdWxQMHQSRsQahBt/bbxLdXgaA
PTqNRdeEx2B+LvQ/kLkZsIu7ez8fjNFtpf7ay7Doo9WbZZs/hqvQ55tduiA6L1WP
KkDIQJgMc08L2cp2rCZ6HlR8eOs+oT+K3KnzPTGQxICo0Z4G/84SrS4hqM6yKetu
r0T6UtOlY7+LAwlqHzZCh9j1zSCSNwtX09tDm1v4O5h8enOeuDkHrdCOUaFXe6yO
n9/jqNPPlfqIHN7rnhm3ENuMdMJ4a910vQGtvvlNaDug0rziWD6Qp3O4m/M03mFm
amwyGzcxDAiPzMb+OrVn8lCWzgYsAhl8u3km3EO6Q38P7Q65dBlk3gKKJeXqXpul
+gXj6GC7J7497GZhKDg3lL3V7eHvdPvDBAJtiTU7pCMvH6dknj+cHwDR2Qt+9Evj
xARcLgOUZjWsOM11zejT3JN9PQM+3brjvRnbf8g3jG8xCqjX4IwyVZjw/T9moyxG
WjDH3ZZHE4cEHkiAzjZxTJ36rIuGuegUqQZOHkGPs/YoVrAKONhCdwgxGxtwzfoD
KNSXW05KLJDl+Mso7sonL3udWoAK76Tr8HY1jMI6VCPBUCLBno4CzSbX936fj1Li
RBgW8JXzaz7VCpLVPsBaiIf5EzXJlpvf42OvXjgpSCIdIK9utNI232DgM/kx4h8p
bGOjl/XwUaXQi9W6z9091iK6Okwbm6j/8H2IAd8n9aeLSPyWKcGPu2M+bFtXaICY
T7/SiABxVQ6seK6OkUhmXzTEqDxCxQO4iSwQAaqK3zLy0es6VamTgWgcKVWMnANI
vzsn8jfxoJSElxI7hCA4Ds/KVGoC5BhlGCVctemZZHtSIsEZk/wBVOUjv2CzdYBZ
kwrTT2akoxohNGHqa/MbMyXN0ejPUYrEVRKOTcPhKxawNKlrYSTf/Nwo8GavnBIT
6a5PDJN5PxUFZpN+hlcXVa5i6kbjKH+9+AqDnZ3rpfeC1kCS8GXl+qOzuv3f26dR
owTLr6/2nrKrYfVfJggMY428HULLm+kE74Roxsi4w9Qia1DrD1BZwQl6FdKlF+DO
EX9C2Pvbf67MmFJgPb0Fa6NPXdSINQoCE/vvhE9bzilQwtk/Xa7GlI2Jmr41IGKS
fM6pMdt0xmGc8op7x7lsgVFFfoWge3auvGe5MNa2m3YmjgpFiJpeSmTmd90annrZ
oL5Ph6XgNFe993PMjNTTFqFb+cHzSYLARzcvmx0Czj4Ciey0Z1g7DSj1ceDs1vVx
SnTLUFtX7T7GDOtQiRARNgoVlqOTd5n38j0gHYHT0MQUH4ISkTk/dOR+TrbpRwwX
I7jgymVq159MTsXiPUwPDvCPAdnIXwCWC+DHA2NIdwEqjExvpekuuFa+51dASgP0
6jMo/EMU97H4C5/4XXDf1ceOqR0VIP7ifjTqRjVYZYR6KDRwcPEgF2H8bGPTT5AR
KTlRbLShtaKaA24I/7olw/yzAk1p4yuFUsH3hKCwvUsgz0lait7BMLZ49Eb3mQZf
TSFa0tBANrbUTQLUbfIo1fXdu+5Ib12l7/qSVraULsWjmS68DU4hdfM/33UQ+dMk
PW66ALSZPm0id8QN1unuFkv5Fs7g44rbm2s9xpzTehf8n7ZrpA0u8aAskrUBgK6S
m7WyMdaOXK286poZmFMHcFNe6IMzMfDkUQOJv9bP3zbNgf/j61w3SMFl80avYLlH
D/8Myt4sH0Mh5EemBMIdb+5kD890vuIQG0Vop2mJ5bYEBHP76GarvknHEC4yQcb4
Rb/R7prp45NTStz/bivGX8zmwUfrwTS+3q+15QikK6VwhTukXo+/jYB2TAB2yPjk
mSPGHMIUYxMGdRYbGnHlqCWMRIIXLNoOk5HVmauj7WpDWSfFamQ6Q4uzKJ108pg1
ZWhtXyV+2yN0AZkWRaVE999KPVO5GpdAsXKf8iInW+Nlp+P1pzmJqXY5WkOLPISF
Jpc264aJBvtqdvWO1PPiNvNsKcu+Q7Jl3R7cbkMQDpKMSpket/CUZ9mIB1O/wVhB
Szke5CHAQEioMlC2Y0nQOP9lotF95aoKDGxX3y15GMy/vISzdrNQuj3SSAfPYAw1
Y/PJTLjTvq2ZenPTbORIzlkkZRsH+ehY0PVzmQUpVVHwqgcI2PBq+MPIpCITjqdL
xAlu+CLF718FOtiWywn3ijgs1hlcX8NoRjpNS8NZx1lIMMPWiKpJMFDudwf8WHkg
qa0Hl99yXgo4eaa4CBYLe19I5iia+oGQisHYZtBghHVsQPTyw+uSRuBRbVJ3L4yV
Y0FCJDXhCyAdZIAABke5RZ9rQhzVibnwaLMNnyF4yblM19QwZHJju+CFnXSu9Zps
ytc4zTxbmKjPybcTarUQdK2OC2CJDeUUYHUa/01DUGCY/pU1lGpA/iiJV8oTuHMi
w/09+1OVns9tSAbStqnDzBWTPajDP0KHGRH5rBnYOpKIQivSUH0lkmDBBSss66fI
WoMSeCX6s1i6/6AnnawW3VrTQN02btwTpS000gzfYvVn9HBHqQ95odDnvD3S6pIw
BL2AX8l6jobMoavHg/7SHx9Qpafu0Tzv9SdE1EYioW1AN+6O0Q9/2MIYzOclKRjS
hgd91xLuvkb/eYJImf1srUwRpdmOUZqQqWFvwH2A8d2zSBBsF0yqpi4uy+QR3JET
/Cto6bEmMqEZg8PMx996gubY7n/Dw8BXVod8KSD4rMhjCy2cD+uXZIg+EG/nJabi
jKKG5IxtVNA6fvI4yv4kGt6ZFl/wSNEyYSKSamkXXplEceAKqv2GUxirzD2ztyNL
W2kFvOhh9DWwtXxK5KjBtnjBnhnyOM536Bli3C5anq40+IIbiJHVV6T7R2/oSLSQ
snRYzohjvb0P4xEn1IVebhBE+RimiGKrQc0hFpdiGbafVNgJNO3t3gvuDT4c7Tdk
ZuABM5RBpkaVVeuwj2qyhQqOuZPstShIkLjdQNWglOrdITZvCwoLy0Wu6pMW+qug
EPC3hNz7JusyHJKizzbKENAdFeD7EH2hqq+u0WxXLLperc5qriobzop0j8v/TUxP
HeBBzMPwW42s5LhPNvlkBj5SKNSMPT/67i1PIifKO6GW6e18A7XFWbrjXxeRVaaX
qq3XOptlXgISdTC6T88RZ7MgE2DvRsCqoY7ebTD8NbZZ+lzD8GcXYuQs2HfuLRHk
ei1ZA3XNrpxSMFbdZgYJbm+b8QBkYKZa6yQjfrP7P7H0/K+N0tXhR5LUbqmm/xjp
c418CKGL5tpqSGzJtI6Tk+LY/kfQsqmv4QjXPi0IXWNrQg5/MF1M5sYyMM4f4vUN
cvn3EiqHgcDyoQwrnQ1XDbUlJU9DBYnCe9kWqJYTl/wGYOPPFhytyIaxWMMSYluq
1qA5wFGtv4q/p2V3bWnp8Ipu4QZHHmeeNzy2bXeKc2RUSAjForhV3aH3g7MPMq4m
FC6osdP4zwdCRlqmRsphirtE9PeHD5BKdIcE9iRidVLJCjGTuava/O7E9tpptEqi
Y4KwZT1xkkJ7HvlQj3wr5tnpF0ly1otV/38Ms2PLBCSvWitX++/Kr5KVPe924yjx
DI5X6WgpuiGYFkzBSGfsggKtQhe0biSFZZVLdhj3v7PV8E2UnCw8S/9aSxRZ5Q2p
Gi6bqrPJOjqnK5eXWpdjqIYvct71rrCSHFTc+wYIvorghuxe6h2Xyru1szExXC6z
Xy3bRdmSfAwG+FwwSriJ/JvKUgPTkMFiyKKpju80PFL+5+scsZ2QzdqbpA8Ot7qT
cqYAVzB6k7zYa/mPe9nfYIsg6FdNNkqMRywVxbn+XtOcyxfJjsCiHXEvmUqTc6Yf
FRQAnNqHIltKmRm5+znpbyRtUjNoRsooGNVpK1D/F/o/yLgZHEqGMLCnGKTPIYhm
LtvRHxth3FgdRiJFROKd4wIc9tkv6k6SbOQ1Y3WFqpaMR+P9/ljVnX0s6JJdqyWF
jFHCPywIasrsX1qfIMfQKbT05v9ZsmS4TpUH32R3KkcX0b0u5LDS997Mv2471OOm
JgneYMiRPtJBvBY/nFmLR4EcbzxUzRi4ZS7pRhfTpf5UYjtXWagAsQuq5j1K5Gjh
tqzYFh5vF1rDy3jLLurPpJ4nVq5ITXPdtMqvB4+19ua6fVG627AJ9CYUGi1ZK6Fn
Dg9POCec4j7ySgfat7nXzPHIYeuBWKcyYFZHMSlmCEKQEoOmQBQuhdGSJpd/6mMN
FYqKvznXdXCyj5ez98157NXWdFCQpGX1c1PMKip6RfL1yl8jP5PorQv2qIIPEIQe
G69t5p+3I3qVGf+IBmiB6/cxtzNhq05ka77jBZN6f5/hWS4hPq6l38yH3FUShWUw
f3Rio2ADfAveaORdr0h80PpHU2c5KPvM3jPOM1MgsY2vh8uTu8TsnOrR6KS4mcqP
97tI5J0HMW0J2kLd+tAnUVcavZqV1CLHIeWkUjrY4/zL0uSxM9EFpZJGbGQjCWuT
mBDpa2BU6mSCeJM+Idl9dXccptiMA/wI08OVdYWdwMiLJy84GcKlUJbZDpnQKkgP
N2F2iGIqESd6kkt1pAtYqaoYmRgVplAKW08lyOF7dNR9L1Js91AOQlSAGGIEGN8X
pz7TW5ZBW3mOIpPh6jBaj00+kpvNRCoFypJKCgTWDOpsEyfm/ovwgiqGqtN+/hhD
u+H1AMSxrRUVlzsl8f7JNu03VHwVkwW0ZkO/tZyyJI5ilD0PXd11Oh1qvaz4G79M
fpsFVu99kqeDH8yQrN6+vntILCX1F/J/puUQfbBgB1xBYUmRsNz8tLc8mRHjuUxA
FqTIO+/E1vuiG4jctehPw48p5UMKj2TBE2m1t1/M2QsWcNwAXjM8l/qWF1QaNsNz
nsq6IaFguCUu3p5XemxS7CKt56r7loUL3UXnr+9hO7MDfChBZKmGzCk9g5K6H0X9
uJX9M8zkWfUCrjIgBCHoRjPrjkRGb3rzeX3OC6us/jFe6AUxQaVDjSBFNuMMjx/Q
IrNlTPfoRSH3ZUEyViP0Zfw7W7PXLeap7sUiFbKtxvkRweLLtqu+q0M45CAgmUl/
K2ys7Kd7gSRU6qUc3R9qxdL3Nu2ul61suQYXMAlvzCGcagcMQv9uSD5Kgt17MLQt
VX7CtDfZ5FUjrpB+5RKgfN7Wr7M/8PRu33KVfXATa38b6szoBzJD0g9RPqWij8hx
9hJUOqSAEv0Wyj15WtNa9K/zgBJGSwkuSIzxqCAgbz31Zq72EZgAZCLxXs/jmZUA
xCVVO4Zvt1lZ05ov0axIZUrmZ89ZGrB7UXHzXAu8MoI7eTGj1MmLXXtYc5elcXtH
qYQi0P7VZNefV6N6doRJFlkmxylRlCg/XX2j6nGRjtNmL1oEOzarJF2FpXswOryS
LCvXsO6Swu218VD+K52ARIhYbMd1yVKgkyqYbYilnmyDNSZjiQS3t3nUve+x4mKO
hcZHDNXZA4c/5P7hk9gOt/YNlB/MuMDU7S0PwgbX8jCKJGfKl/4bBJN4GwaOJfY2
rM6kkpN+mIl6+re7LgioOTiAF9wIlIc38e6IQ+Q3a5UxBdxk4pvuuGjwooVFFAqP
zsFQ2TvPpgg3ynj6mhq4b7guA9xuRsFqVY2c92tPoPQdAiMMBORq5RECB5hBCyyB
2+PNElCQiG3t1LOOtfZGpqkRPOLfWPtnUYar8Wdp3w9KMDwjQM7uDQaYqq6BRfUv
HqRm3nnqmZ9Whup1ZyKwwVvfu3RR+1Uqa7XrZDz0FugfaC+hhYMyXVKI/scy9PiT
wZF0okib8xfrTT1UqXCXPN9JvgLPcVCkZeNouhUFrR6oie3inyCneIFai5ALEPIF
j2o5LwvfCTLQ1a6W34s1iAQIjzTzqyHUDBlOcn1B7vlT606AfzcnCewyFRJL/CFn
JZiMQe+UmC8X/jO9mYwrSPwXbAqdN+wGStTpdzn+MbFXa33pitybKtEBRVyyuJpY
nK9Gho7314M5lPGDSAKHV1xFU7A20hFIsWCQvmP57sK5geVoYZODwv1SEtTJsPWU
gvBvS+hsaIk5gAjoYlUj7eFQFnCO+8+PWRWShm+vwfTIqb7pfK8nq1XgE6SiyEER
kMVDhFn7KEbZoAVkwAFbNDCF4OT54+agoUtir6kSfQoauohxNYUVaZD5Ag6xrjL2
GHXlfe/j0Fu+YKim8W3EU6fh5wigwsyCLOayBj90pBz48L/sHbQQaZ5gK9oc0YCQ
X+uJlxRKQ0GlDCuctYYblUiGoV02u1weNKclMDPZHvv+3oq+Nye07DCYTv/gk3GV
Lyb+ufgXo4oV9oiCJ68phuHWy7Tr8yX8osdzcIGg7QYuGrDYTKrjISZtx9lTKV6H
lHLnFjj+5SLjT52s6JvX7hJ3ktqFt5rDmSu+MaR+tB47WeWtc5r2//fVSX5JHwO6
vqB5ZpzgQCNc7j6FPVa26wLRPFtUl4Pl8m/OZ7p+dAZn2vAL6OjCoofp+OH0Kao2
px3wsCwqMZjppW3iWc7OVrEGjqVl1tUpwh2ugOD/R2v8GJgzWRcWHIcHf5nJsXiA
jDnrR7lZBbfKqZnNjqzmt3Fyeu3pf5/5lcIiNPuOCrSRRsEX7pCr4O5Sd4ulm/2+
edgfA/IFX1EBQJk4WiaJJCjgDGJwL9omAckRmOfEuwugQoa3yjx5X1iSMXXi3Ux5
YTdNPKU0G+ViAE67a4ONFELiGM8ooCo89tgJxCxQ7d25C4w1d+W2pfSBdgWrKGtz
7fIMD079vBshiMSooxubkHu6zTBWn8ky9KTKzrXmuAsEv3n0HA7GHrCgoxzc8lac
vc7QooB81gEKKZgLkWasbyEtBpmp2oelansNutIx+qWurLl5IEkhUZAm/e+FNLn7
17LLbt3ADHyZFiRzGHfHd2NeTI8xZxzwqi6hgsv7gdtZo37d/bHSSAGggFop/Vax
MMXWCP/Sgj7lRIFS4sRYEYO9TphBj4kaXOrpYpy/FFEPVwWfkAahS85oGpgZKqv6
IvLz/DLdQiAX0nWoyCig+pW1iDVWafGW3Yq1myhoIAxx16fRe0IUoWVJW27eO3Lr
1j292BykKA3NjX5sOQls8e04sk1p8Iun0vliLrTh0SiZfuN+f2gMT+Xm8vOijlj8
k1WvQyRkqTtWThszfpW6DbBOeSh0zNwDLMAW3+RG0Zyu3UfSMdLyXFCDkd26/3au
7/iiIFj53TxNbNutEMWXLwF9lzBZq1gjOZ114/PaZYA9ejYzHwEjA6VS3ZchRPv3
nyEF1x1NrqV0uZPHFFhuC6O6e6EQXKzRnh8AxV2WMYzkykQbR17IwqAgrV9o4jbw
l3aZDUzni53m8VPpkxCBIsqhZUhBGMz18enB/KDrbjX/KdHImddisqBRb6MKGLNl
Lnrbqv4yYGevp6YxPkDt61o783G3LlWzHSIHMy14INvgClG6Bx7IPu0uZ7StXVj/
NFczga2MfU9PhKCx9L9KAzi//owvMK+4OpWseqU3rdgIFFIJ65ZWUSKhTrjWfCXl
AnWqrRY0Sk/9+3MBMOJUZ1Nr91KA0WW3ZBCPnlHoAHz33OWLtcSNTYwKYyO+Kv+I
nMlWW0q+iD972349DPYfeBDhcnU+w5H4fDOfDY0mZPLfaI6I+fyWAImopMX8Uhd6
CGYpTMTuPn5t+OA6enFahIC3VuSl25AU5Ae0C2cZHfG9Tec1E0Kzha211OyIDV2o
9ntrrrXEQ+hyc+MVLGWv0VTi5Ev7MpiiDGDhDz70UhPecCueZRFaQaGeovaupBeL
0XH13PekJ+h2jNKv1/EyQFGqwbTC0LtZtpR6aPdKLDUbs4cWsyHQc3UPKX4X7jbl
xSweFzXMHDtEReE0nDDAsPnqtNRj/E9Omr/NFS6GYrSiBdDZ2RxMJx5DRfrwtRSN
FKg5KJOfFBw79z8G+fn1mxYj8ex5x+GuGu6Bb5u1mEDk7HMJs+YJVADP9x5cS0nr
16KZayHtvDDjYlYcMXz+qlaKQVNOjYM7RnRS1HyfXtpeQfDcdOU13f/mzx7DMxVb
JZMTndsDW+fZ67q9XEDVvzR1HctGg2ozaJVksSpMDPbs/ic8D7twXO47+34itcMP
xb6iXoHZArvvdb7gXQ4oP+nhkM1hvmzl1e4Ldir9kgbYL/7B6lbIyCSHr2py7qcu
BoZbNunUfkuzaMq+j1OKBCS1j8lTNjIm9yozojfZ9s0vPaVn7Obn0Emo0ZLaEycx
+9qz3NqO5S694lWE8+kR2pJM29Fh/K1oVD9hDhpoPxBw7oftsA+01d+q7HSYuHQZ
jYYTn6TojHGk3ld5Z1E6LQfv2xvzlVtAlWz6jG9nZMownY/5+22zrbCzMw25NM4h
rTl/OvqlujjhAVlKwLLQ6uGOSTt6er9+O+WyqX0T8OnaItHYzgDY3B/Y/x5qeLHJ
Do/uZUdl1RLLeyJvA/09cpgwzezpmK4+f1PGbuctHKUTfOhLJPozpocR99g1uIZJ
3NNchf6PP1NApEajVCiPW0E+gEpXNpKC+WIZad+OazAv0L3UWPpb9gaolZams+ve
u+d9C2S8yMlfcMuyQ2FPhIc3BSenNslSBphkLR5kZwTXEcVKBhx4ndIrLkzOxXKW
g8ZN+feOFZ9sBQqhcwVTBMIDyyEHBRYav+7G9nA8OpEkzEs8hvxruY3wWgGpT1Io
KjP3tmFWu2B0bMIqmYy4nVomypD2jc6Rsu0jI+K/f9KmoLW6o/iZ6yYTzGXoqGFG
5dNzhO9v8iZUjud55cnc48XoAeGpL9jc4Lp8RxpL9BzPRTPqXwwEy2bASdPUBG3Q
GXAfkNCb3OM3GYDPs+A2ZCkfDGdisOuvo2Z0jT7MWiRhqJTQyB8jIVM+lXuBUDhg
LVBNyOXyJGxXnfKTofNIoKcOkgViZ1QfJv63hR6rvNoS0/lv/Yo0bwVBqmoJdyPc
/1l2YklFTaI0L3GI9fMdwuU9KOZ5OmKWh7mmJ93jy4i3TWUMjhI471Le/D/ILXrj
x9S7/tPRdC5mIaXrpawP8ep+JkdXb402hgfP8YcTIY1cYMCvnaIc/f75SLBLWqcv
PcKQCTGLaOcTcoc9k2EQrSRRQPeJT5Z2vsJ4/dGQSp3sRZPYVFTBCw9yLB6sblho
7sRPMHYTCUXm2ifkFOdJQYchnWoCYnZ8CWqGA4E260Jo+eWp1+2qGhwgeZczyb3f
oS6xneBHJ3u3udZV24jNaVEAWp1ZHkLGFeSWv3yxhc3yOQ5VGPlbaTAVgsO+XLtn
Lk0BM4W03/TxJqy9zLmb+8lNOWZ2zolvF6/Tes95w4bskLj3xxMsxjYuVV6UV9ud
hNyn6hZbbznCV4j+PfED9iBYOwFn3HmxIp/cy5aMGD+xaUBSpoGKt9cLYRGFXB34
N1jjzh2fVyJr+UTL26be/Mx9OcVCdKP6tb0GwZlRK29NEmARdEiAuFX/9cJh2H8/
TmrMozQxnJp7nCk0bFzRseYgAIWaejPCItZQDLT0gWxKQUgi9rNSb9TRdL5muj9S
IhAPkxlFH9TvUOIKKIyOZCJa7izYBPvQ4riy/JOwiyrjkCzWjWJ9ZdQF3jbHC+/Z
7seSfW0P9UNiJ0SwKKg9sFoJc45XIPwHB9Izei2ViA9j5RTzPZG+MbXkALaubIUQ
7K7w108oqaPlVUu2oR3LkJ7xqvqz/GPPxTEpnd33OtiEM2aF1Z7sUiebtQMFKemd
gegqE2vRoge+4Bs9f8Wg5chGYAltOWsBMHO4ilcd7tTBFk++gndeqC5pMFCD6x92
vwMm3jop10n62jv/5z6xWut8c0mRe6lkQwYzuwSd/POdK8C3E5shnsbVTvxNntXT
hMRjAVrLd35lNmw0UH0UAS+LYu/3dLGNYCjmNOwzHopFjYQjBVqm1/146GYwHze/
nb/7rPlqPb/NUv/Yx6bVMYDmJCrQG04XWML8ybsrrwFiHtVbdwdoaP8f8roC5+Xt
DwgHgAi6fGckuOGee0FOrbTXOeAVs9eWTkEyxiGi7mvLWGmTPrzKj/4J+uLCk23o
9rnaBqEk8z6OL4nLvrto0nkLaTkM1o32ecPk9WA39CZmsyWC1KE6Y0qcitYVqib3
Ft9xrDzLv9P4IOy4ciKdt6S1ikR4QPImPDwhD9ZAgJ9EzHZfLUqTFH0vu5PRIu2z
e3boACetCSOX6t3Ao221MX7kKhMf2a0ED8K6e31Udnm6KPtVWTUsCLWL2+lDM/HT
cwj2BfODCsCx4U6d+ZBRdSaG53PxyonDPdzkrG45GOlLOfK1ulbCpz8H2ivYINWv
WrCzP6p0kafnclDi0eNKG97xZ1E63oQLG/jB6A2AMZWnMk0CDzrSXeP3MGF6kwNu
XqM/X4lUhGrST3LhV+EgD9GreEEroiEi7ytpx1vbHKsKK6rwy3O3wHozyaS6zeOJ
8Vt0MfjSryM/intd0vkniDf+w7KK9Sn36apl2q0Sun/4st9uTXQnlM+jJb9MQv8H
r3IXkM7yZ1XZMi4foF0i5IdHgugRQi9TwXL7tT5CRXN5tImQZ83VkE4DfgBm9pr2
CGzWH+TXifFiz7IjoBXL1/41LFI2xGSlV3P8e0G7A8gmFkUfvcggWi1VCSrULtPV
yIZedapTO6AGhnW+FjtqJVb2Yjb6QhbeSoPgLCmJ7CcdNcVwqJjW3rzbyXYVajhQ
aNv1L7R2v2jJYqcQnhO0wtkQ3/gcyC25r+mjyA47EFaHiILpm3dCclud/7wMoO6a
x+WhhJShJj21tR20EQbaaDaaaJoU9LnwfpNG1vRzmIZkKA18CeDiIFEf/Ei1svFP
Bxj++rj/W8JdSE5ekzM00IchPQv/uETDUKnCSAUnR/STHOQS9X+LkD/hSxpu9mpq
QFxWsj9USt0QTgHvCndgSI9umNtzpCE1JEoKlvlw6idlUSQV7lpO6dXAlNC1PDq+
Rq2RbP8AH7/eJsfSOLSREK745RBv+tt1XX76W8z1dLuUdUI0GtYE4d9YaWY+x3hd
K9VNqSQK6UgIQyktplZHX0lAR3PWeSWjY7xQT9zmmtxcoZepDj9hhb8g4uWIECl2
penJul9r5jgUlxmMww2QkpQA8ti6PS5j4+Clncm/n9bA/yEFj51YrhEKVby5kkGU
+370Ex4AoG3Z5Wg2DRacqpSnfE2jRZk3C0jEoA4pLkObb/qIZBa6y/vNhfb4aS5e
NtuIpauYWbZ+XNRnO9XRVyb3pTgMJZFyQ6dkQ2XVO7iWujIi1meQygRjy7AGkmL3
f8OcP3AlV7JfnY76IWYSgkNIyyj3+AyuVicL7oQfX8TSW+QpwcjaU2YyGUWIl0Lc
9yUUzIQFx2wr1qmZQXPgvuQc0R8zXE4ae4EKqs6lAmB0aN5cMQXcqzTvaC84SMVj
hKjXFVJ5UGcrIBT9Kh+xHPagCF0rAQU9Gqlgprsv+XJv6ZBL8CSst2kUkwHIPK6z
IKLmZvF7OlMV0YHliUF4QsyRmeRedUhJQ/MjHb43Hh/igvxu+iUmQnrHolLwcPYJ
6MoJELvZ+4nGRN9A/1QP66kJrhLFI6N+o6xic1LIYZ7Y9UZ4rSEuquDGxLebAlyb
ZeWj2THf5uVcYtIt3AxhFTpeGWjx8MC5frcmy1ZRLlYdyfmRTDFORF3AuqFuKMAu
WHxYZtIVXDLadC+cOcBNnweLJ1KepwbDQyF4v8bMuPBzcCnups9FTGcDnmr/Y0qe
0rd5NojExC1KNuhiaqFQlcjEH2+sh4L4/v+eUuvv9RtJACyYPMpR+KPHGmRLgZYi
s8wkx7JMrCiP0XOlXr8e0TqTF/+3r1EjLZfV2nlkp9QiD7pO7cGCDZtmvRXmtDOY
VaQ6W4mgduhCLKluFqBsmIUqVoa4pPsYMJWHoBtqNU8uCGzm1pAFKfGn0DU/q3yi
Qn5pHfL52TriLuzV0o20iP5P+cO4R8u/0pXz1zf7UuJKMfGyFh7NiTETFlzBueSH
E/1F3tY1BEwp1E2BRH0B4sIkHdim7Nn+uxr7+XcrpmFxrFJEZVhEj/wzI22EZ0K9
gG4cK+Xn3l/x2QeLzp3ZA55RSlQLbK2mpurEjO+Yge582N5+JNTS4aAAAelEwofC
Ft4JREy6Ft2H2NGfhe9PId5K9+kt8c0pou1OQIR4kgUOqFO1Uq77QtaI+1CZm8SK
hYpM6iJ4TqboriCr5DHLA4x6cwQ17C/DEAPg/5DKFXisf9T0Cx0Z0dGXixQS1KAO
Ssd2KMqJ62fZ05pOlLRYASvlq8HiQrhcUf/BCCqSkgbcBgtA+BEp4N+dcWcEUjKc
x2nAB8hDB6NeTZk0MH1vQKj2jSsXec1yJBR8nevcwKIhydA0SbKMym+D3wPsh0Bu
IkWEdc8wQHM8gKO2TVLG9M1+X6DpDhnYPSVF/PFX4sbvQ2MWyMR2bL/Nvh725rto
8s+HESHLnUelHEZO1z4Wx5732HjHhT0hLUq+4X8pWjBoONG8g6Q1K4KtfbtWwj0F
kuRZedaQ3tiqoNitxrR0MmjYqKhFNsK3BAFkmb9Ly1h1kh+jJ9Ooe5oUEIhMCqbL
01jE+H3l0CmL6HJic/o1TC7j3gpBqiCtCx7/GOycoPAX7UVPGRE3uZGCEC2u00ia
jrxhND7PDfL5yMrt9N37kRMwsYoQoaIVz9Xk3yFnGC9AKhcUGY2EHpFNXvstp2LG
7OKKzmSsG+/6IAjfPQMyR/dMbhJuKpRFnc3VoMZkxeN7M/j3zhfgpjuG5ywB8K2u
ePUNe3m3EZv9gfX4eM4zOpVRd3mPsAu1frrMSlPV2yYzmslY5NDOSJiNfXUbrnAL
a2VaF1Zs+y6nqOJmfQ9y2+u00ejpQ3QtGzLMVSCZUnw7MRALiTYhVtDAwaQY+aHJ
89whRlWHvK1wAZAPpMkCjJZjp9bQJYf+2Y4NCUxMwYqUT/6APP3hsKB6y3P9H8z2
sVmy/YzmUgUeUBMnPZ9ErbgvXLpF8gOwHa3Vi6Mc2hL7AzOdhBfmlnY4Ilhv18JS
XXp9wucrTfFA1x3xNZkOiQrgUI8MdBXi17Vp7oo9byNxJfAMNtpJJMD4neGuy6fa
NNuSoqU4XLzmtz/reHDYJexRT1J6WwWb4X0Tlw6z3fanxQ0ncU6d49jjigxx8kE4
orlT44/AQTeinFrxw/H5ePzxZNzy2UbYOUEYdJqBIUcrQiKvln9QUyl4uowus5OH
VLod3Isx52J6mI9qZ96ceo2z93YAMN1zSyUtrQuw2AQzaU1ga5PHRNlgSl+R2z+Q
0dE3B8PtU8oHrCzPteNUzEqw4BZwuXNRg2IrzWOR8wstGXn7VZSMm7LrUKxQVlAI
IVyv1fuLvTU5rMOxJShLowks/beB+DFeEqlKunctH1l14xP9pQZG3Z406hnYkGBa
K5REPYUFzEkk1BwYKxhf0Z30yeI6b2ZBS8Ae9qYGD7gtcMRbN8ai0a0eLbbbKmg4
LC3OWCT6TuhIacjZ/+kqtLk0K+2JkFRhgWM38q8I9yk8GMXiR0g3h01KvtmAMKYN
1NPe0iP4smTVM0txFPVAkpTfiHfPBjCy9szd3ulX+vd3WohdoWWoOFphkgV703jn
m2c5Hgm0nJe9zEj2RqXB+AM13CnSP6SMjBKAvrx8xRlWcwGTBS5aljnB19gE9zqo
rHAXLeKlp6+Ul5GB3a8JjUNk52UG5V10KPlDzLxYK0sHQwYN+gDseT4Y853V7mCo
eFXP971gUDWdrVtg+qcFTRYrebcbMlZEyywz+LH2ILkmg8oRCUVuHU8gmk94qVoo
biegMuXrkVMCSezzWm/XHZaf8/YWpKBI1zGgbo2EFW+vHNjmxHzfXLOyRSC88dBn
61P0xSjOXkA+Qs+gbzHb2N+mH1K5eJE0sVzUHXldfXr/vfBg15WrT9dGSykB2Atj
0us1CbFSxYo3Sx3sAP+wcuxQN5Es0UEORDqmfcq0YH3tUTaJpPXD4rAF7Ut2O3On
ed5Mu3qDV72TB3grvc6miPvPVsQeXAYKIwXYlXncGR+7exCjpnXd/w1NPaPuubwA
DHxeZR2A2+d/KyuU3P71x6XsZqixXSo5x6p7U3rVr/9kdyU2cP+OQpIB5raGmnlI
UoWHg0fk94G7udX0ECNslyDjoDZ6J46/DkeXqvQEolZKo7HWk4q4+Wac1BhK27uO
ZrOEpL60um2aPlNcGPlbVYHBqic0ixGbqYf0UHUUhFnGn51pCxE6iWv8m3inziWA
vRN8Yd+RljeblIQEKiJWU2pS3kiwxkfBbnEEE41lUhgpcO/T+tG7iLeTwwc/oE2d
Gd5A44Sbt/fDvBsoR0HXKFQvJMuCNKbKPNaIJ0TpIvdi98UpJdGJ2O0PwfgWKCaM
tWkxvGussKLw37JrWYu7kHsdu1LpV7op1HlsyhQenfq1IggXjE8AevIrjHWD0nUD
c3qKe1MUiXZF0fMw1l81vTjvSkbx3WJXEMqyGYrE5vxaGjnEU4KnXTBB+ZpKo5bb
WS2KMQ/pKPIV3b+H0qvnaUxkDK6YOPc7I9NUOROCW95HpP1NOZVKYxURQNZc1jNM
lKL06YSQa8veJKfjcwULit3k97VIvKE2ex8g7kB8rgYYXMAYvJBLwHhs6Fqznxu6
5Orot2/Mj4vDqqX3bHNWExDT8MQ8dpwTp3LuOgXQkwqZwxqtaq48SYsYelJSfJWg
JkKq5hJjG16IUM3/Hcao/21iPPEXPIPWAV8ga/NkO2ywwiOpS86D3kbvhm8ItfH8
JyFYQ54ft7Ag7DZZuWC+l4iB9VXlh9mK2prZgmqBRQ7GU225vU+q+A3cbwNrOkiy
3rcEYogBPGyVCxfer6eLVMfe/sfi0CCi0FPkr08ZHWJBED5VrYNXthCQdZZ5Yq9g
0FvtUSNHk86HCUGdHb+vQDirG5KQ+bExA5xv8l57yT6nPx2rKgRrzd66LV65Airj
FuFfbXxnCCazrSRJPfaDYRZVHWrcAwyujDf6YF5Brcz0bKqz8zL+1kzMLauGJ6KT
mUCuqIF8OCorOh26CfyWbayaepw1X+XlufWMl2TDw2GOyRMjXZrVydbQom4H6nSk
H9wdgA1KNuSmlc0LOhXMTqM3YQlQkbjq+cYnTPdyz1ZKwuzL2gPxH/INYhAlzPeN
REk+Ay3qB10RZU2QUlFfmAK4tSJk5pVPewQPjYL+gNKWts1MIv/egTcJcQSQoTBc
h75n/Y5P8xMqg/sxxEvmEMddwGPpi7aXlmMdhTPtlvhImiqXwFHB2UJLV3K9sWJS
54dQ8zuZepWWjft355w5hEgbhW/gB5xBVxjbPHJRUiim9iNYuMaYQtfaUlnmOcNN
iCZgTwxGUrqYY1h326rM7sy70+8clSX2iBJv+hsB0acdr0CoJ329v2AovS4qWjYo
9xar27Piy0whP0h13r+bOXxEiFqqvxkR8dcM+ajyffc+cJefE5mbzHwbHa9tHXkl
c7jhzCyeD6vxXjnPX5vBUT+CKptM7xClQKs7qssVEjKEWC3ZF6ZSws0qX46g+Dl5
dEogAYmTIcgN2N5CusMQiy83rWRIUwaUr1QvPoLbihMA2YZVvSREl3kMx9+Ejnda
0OdMYhayGa9nGTsMCxSJTqe0ujNKsOo31C62XV+4oaBbI25PrCk0Aihv5hY/VcKc
nHa0vrRvZ+jK3L2squ3a9PLtpqlQ3zw/mzCeFa2/hBdS2Z//bdNtmbK6t9HkF579
uXrBWzRvy9YtP9P3I9KGnfYHMMCDlckglrrh/KhjDCPbJW3HI6sMwMpSZ5hHkRhs
scqXQ1clvV+E5kQb0abpQcWp8PnaoxMbLtRbYjIOS5yLZWYRg3g9vzvVq8DeL2l9
Sc4N5e1rFlsHxXTfPbs8eH1g4av2hMnUWabNzJPBJbuxS8ckrGEqRmZtisPE1TFo
VxgtUEiOhf6mLDXyg7EzIgcOX2MI2EP2VMnC0StPKrwqELX3u/32JbvMOof/9L9I
7ZA7KaECIn+CZSxx8NaSLCnDJ9fAjtOeA8Hodl4GpqjGwWPwr5Y4MVrXgV0sKxZX
WMHC7B3lVnrj05VEYWAoBF/71sCExV65cgUIaRP790Huns5Q/t2VK3QCmFJcrs5Y
ZWyD/bkWwf8FQdSGbwhMeo05PLMuPC2clNe4DGJ7W+i02XBjW74ELt2LpDnbPejL
3RbdzHiahl1QZ7UXuXhPrkzzgSGhqZWdszmz7FTwiOd3CIrh4mi2gkTY+dj24Rb5
eTNPcr/NJcvVD0p7Ok4qTLtbiemoxDAS60zzPjiMxYmHmOontRS1n0Hq46reoSF3
6UdGyvoRHyTQOfLn8HrDqvPDsTJvTWYI00HmVcG/a/SjT2qVyuUa33tVxYYEiuz6
z6ENjJitGb3VuQNX7y4cnEM6ExRgWY+qJPpSiK6xiJ6MBfjuQzeYmsSpMV8jRIdj
yloCeiRS6lhbVYpUsdfSB0ap8AROCTOlwbnk60Z3uPgYs0vHoseMTgzAVnCuV34o
3r4UiBoQKW2M/hHmXYB5npDYMEGcWUXRTfk3J+CH3TD5otgOPV1IAC6WzEAWDrTu
qVskASfWqyEl6nGZBszLhfVeN26Z/cuRTO8fVjVCk89fFRxqPendPi7FQ5+HBISK
/Xxr2PrdG5NDLzag4u4qe6xZFTQc1RgeurqZibscOjOeDCs2XCiXVyWM40BD8OKb
8b2d1EYWiazW7+8KXJPrDU61IjKW7zWe3cB+hXp/HjnvkViX5U3qogdarlmSslUi
OlyfIV6Voe2yV5cglKViXYTdYXYW6EZkNeB/G0aaCKBEnSIYv4cPNCw2s7YAInhK
I0cdUxgmNUy5J2Iio3uGyvQ0tV4+wR4trkxZDHPfXk0Z/1F5CfuVyiEbH2KQdr4D
ys3ucp+4e0xTpNc37Bb1T1B40SwvyJVM7lfXwt9MIpigwxF8+eaQRuiK7Lk9rSR/
+L5TsgJnLuKnm+v80eDFx/Orhv7FY+Ot7EqGx6h769eyYEtLWlM6yuSB4gpiL1jZ
Qd2w91/UY66rtyLgHK3En0t+x1/EKj+XXP3oH+0uprxL4GqkRZgpGb+RFA8qV+vj
/yVm/fSUc0+Uvks9KgT0SPSbqmQtcIiRp9igGiQ+USi7fuKYHF/edkEMGvHK4pAO
zuu9oFmzLaFlwLGPda7EBPElP9V48DhzF9i24QTI94Iheu9kVqjNCtlHoh4L3I5V
youlYtx25j4+gObdfaF20cywlYBEFjMVTwnHIhDZKPFcYO51FtkX7ZrYyUTAo3/C
ggq0vS2mwmFF4NyJa/kWH80TmX62cWVooNXeGa0iIRCE8qyqmtaUdotLUdEEKq6+
IfPgvEEvXuPd4EK884RR5Ok+PdHxP55s5s89sJszbhq98+Y5+bT+6s5V9NzbexUo
Krmh/bvJ7xqPAWKEkt5hrwrhXZ4CYVPR45SbI3Fpac4twWX64hGis4schKr1Xm9t
v8BNzRrrf06CrugNXLB6/9yiILREL5zbEgBFNuk6kQJ6Swlpl0QqU1rl7DxVdfRL
7yGGxXXFFloaLAvj3V98/gFYZKuUNmO6PAzJtmIKVgZaS3II/ulAajKhfgecI1FL
5EHV9LkmsCLRBEW+RwuAMm/kY30Cimr1yMFjLAt8Vwoj1O3FfF/Aw10B3FnZAzg6
RU3VnJBOqZUgOfh/KG2+f/9uXGjj4s32uBKON5CyidPhU/nMPVTQiDN2IkDxrhIn
cdokHiAdZVcuH59xBsZAwIzo292p/5kdBT1wvUKWQ6nWuz0NN+5yKv/VikFIOqmN
mcLrDSd+QfXNC1UdcD9clO0XnodsByUx5awFKJS+QtFtwRF5IOKjB7hnObfhjinK
3Cha10cCTud0YPCFGDIIN3yniMb7Ou8oWsdrmgo5AVZmPkgIo2deiDkhZa+heu9C
+4gAydDaO0HoMX3MbRvecMxvhxHqiqO7LRwowunoQmSSAdoSetmsbglBFaMJUFxI
CZpWMrHFDE5Gx/JphZVYDsZKczdQP+YDEUq2HBzCIJcjxdowS/WWxCiejA3628Nc
7q2Qu2/gJcIglKKonHwe/9NgQGSxKasvuTJEDV0vi/X/00BV0Y+vwX6sA4plhOd1
9CYLYbZXMesbnhRHPScqGNk8D44/6gqsWw8oubg1m29pySUWpC7Y7Cyz+y6OpI9g
v/WzRDrp8rKe91JSKPB7jz+Hz+exszUrGwCeUfORgm125VWPfENZUlQi72tepN1c
x+uB3iTq+pzcmIXyhqx2CfwI0/kO0TzUwHoI8W69KhOP68/fo445ZipSugmFRu3+
fvCMtwLexU0HWM9CWmz/A3tmt2WhehvDKdR+1//1xAn7sL4FfkCBrliB/msbm2jr
J3iehCPhQdE7mSlkZ4E8xUs8OSJJIEKgFtX7yoGL6baFOl1jG+iqu30taVZacEnx
KB7LebXskLoUFkNlKk6FHT/hLoh4o5WfodmY4XvV63vIyroSeJeSv3zLimGR25JF
bURgaaqizSuqYe+Gv8beMOfERz4uPBZSrjW1VvJZOMW8MSrE56kyEBet1+IygS6U
z24L7uYjx/UgdD0QSoIQiYMwjkGVg55DXunvXI31magvtmMtLDVVQ86HWV0TUVSd
8u7jRHmeo+E4rse60OArFN3YKTHaJcUCSTHQJtlQZbkoqgjPYiTlji03yzV8/Ihe
YnjFbu1G9Civz01F9qTWA79lpjkLDLHUqJcFggV7woUbGS0ccmcrcm6crzM4vBva
X6lSkXNXtVvsCnzCGLX7oF2TD0ylVezIAV3BZSHdBJ8nMVyODUTLoPNhs7YLVlAo
rZQxNrozvTQ/6GSSJTxNRY0Kc2y/f1EUPwvS1DqtIpFvqokmstucXrhfT+IETDa9
r2+ROJ/5Z7NMazIr82F5K9ZT6pIZURn7u8MrZwowBIBvXUgor+OLjkqT/2KPL3x/
Pew/r1ojclmQGBwvi2mbs1oZsiqZK5zJZ/vTf8w4yIKDhHUKA07yuHcXUfGsNscI
ir8EPUPsp79X0bsnP2ceMPVPulpneqeX4XFUL+xfx83Zso6wdykms+Vb5lEzaje7
RgKenw1hNiCu05PkpFWCysILp7dRlXXvbNy5DO9+br6Mqhpdlg0lpb7Ju4Lbxqly
FezkQsF/H9iqQb8yjmxRMEx1Iu95Ww4Lb66GmKxju47KS6N+kE6fknc5EeRTdr5Z
3s3nkmwLuYD+gOq3QcOYo+BnYZX9dfscs1J7OGC4lZAB8fTz9T5lql1oeej97yXG
ZuFxJWVDK1nUa7FAk4+RgQVhsvMX+mFo1eSNDG3yhEHIi5JjxJgonRt9nfCUdlbt
T4GMrQxIwjyJTf8BQPZaXVLvy+Nsk8hjKdJ7w5MUAPM7iYPaOT55L2esV0DmR9hw
/1rcjLtYlI38g0F9xcpkjzRHbCgJ/mq+ijVIwCs2dOIMBU87A9ZVhScTnkFoPWWf
gB2T8kMD3UBPKS57b+gBCLpc4X8Vm9XDHjp7H0B9/A8o/qPvlCvuQXKWiWpPtJJP
eX2TwSgr1SMnO6VapvNyI0yK5Oajb2/CKs9SgQuJH9/m/sZ/xQ+J5akVYr9D2wAJ
1I8PcxrxKC9VdRVhuft9Np2zyFRkgAS6c9VLxYV6b/bECV+elHSWM/hKXp+wNdQq
8J9e7aYY6iojsXzsq7U/xY4cxY9wMFXI/VGv2iw/8QEbIQwXhLLKkG7sRHcUKnEg
PUwc46BhEfwGZCZJfbbpNW4pXG681IjNL1E0qmVG2iS9aMyjONrttCBb+iFY8VgG
nKPFpCVih3n+Xx+PW/gjSoo2Qq/7OACxKGm9l4eVg5QGkkHGibfyLipEfRpRAkOh
iLaPatEbilw7bJQQ5TESiwZHEtq2vV/UOGeV5++m7LuUCOUFdjCR/PYoraOn6VUk
/U9zqZI9pGKyDAbwYPmJqj9Uy5ne0OAfBLC32dKQ5SbPJfkss4w0ebdlorxac/jP
m4EUyybG1DKTa7hFatEEO8ylpiXUKsjcqZ0PXhoAPgLIOVqbKVXgKqFJnahwVwg/
bfDHheqNdDFw4V0KButhBcgohpS064/m2xj7MpsBTNWY0i6OUDB6gxCM/Xg2xtv5
7/As453SYwUkZIhLvsyEB4YgbCbbE13BurZINpvh+Dz/4XhbTw8oC+4P8Lny55f5
qvg37RU5zKr8Ava0AkNwxJCXYaBNWDj+brgCZr4xHs3K65zXPCyPYeIXR2rdKNxP
tmuaRGZz9/U9g7jbAeLoPVqi05mK+3bh9PnLkKpR5La8mCLP76UC5nslHijdJWvZ
J3PzDPnxWemRfeWWz2eCt4Ny+tXBsl7sLs+4K8bScVZnBVqPxn9ET8Hj6FrQvbZD
JvTOo+N47sPmeu6C9KHSfLZ44mruXQSi6QCyZYfBmrmoPp38zNobRhLsSB5xKrh+
g1tJb1XTuV+3MHEucNRnjG+eLuWqLbBRFnYhgCDJRswObjhU9OS/ZEi7ku/PO7tZ
bI9T7ZMDn6a3AcKISpqqFAF2gy9XnE5+QV1skiSkfUMqlEHotJkpXuZDPi1PuZKj
PCiArgTnCjfWGTZUVZDak/phomWuIeTUti7dYqSGKqF67SneGPf9X63uIlo8i++B
Azi0UbfKjMi1cDt6aCV4VqEZiHJf/a7dVFi0DD4W5rWDx1chOAcRcHZkpwi9T8NR
L7wVV/iEH186EXEWCQhpa5mlF8j1DQ+2Mu8GmhKiURC+LtD6/Yx4mcyAIIWYt5jJ
6nwe2AL08SVEdcDr910g1Eqt92CNWAOj10KH9EZdOs7RsdDOAVgFbbMEiK9veysG
c6PAyo0AjhhBXyP9CSRu34941Ibi1sx7+ZOl29S8H7sKiQVOeKFMhwO0THREO+mk
DMVZmNn3NtPp3ocE24DRNa4fT5t1WPz4M9LOlkSxBw1VVSE/zXuJD7cVLXXMjLrH
Oua7RvUeZR6KHHQDw2S12FFKIA5ISEFJRyBNv5HsXB9NqPRkJrpXMHdGc+EVSbF3
QPuimVwM4eWYS9uDM9ABCkCZt/hj0AfYvTm4FHq+adVBa7ch+1J8A9x8qMoGq+v0
vojzgPyx2H2+41kBTyePIc98NpnOflrjo/O64Qm7pgEnrnjLXmPrGYt1VC/R+kUy
Es7mLRGN3awXlPEDjyPxaN3L2gBqpUz9Ll+KyHGtD7rbSnStU77I5XWY86WYQcNN
Fx643nBIO88H2mhfpMYVrRPaoh5Dq1fBOSeMMcTHTa1JewVif5M1YKB7eGNqKbjf
3nk4QMXJDq2uPPgGelsxJ0F8546dVzde0OCayM27/b4RVMwL4mM+MvjYyflSZjNC
8iMRZC9v+bC3Btz4HWMH5Tl0FGnLZUWKNbenZAJWXI/mml6bVS8f+3ZOSNLBqTcn
hseLk7B+UEutIngr7lpV0yx61iXrRjGtQaSgg48UM4L5YvVfTu/48A9+XbhE7LRb
7tj2+mY2QoqopczuxmXKL8SXAlkTWnx/QV1pJH4Aq6HxMDqm6C1q1plakUF0K8do
2ZLJBaiLititE2jEOnvVf98oCaOEfQw+YLvGAF7gdmBX1aE1aN7bKZD7lSZEaYBw
x4mqN+tDCmVodKRx8a26Z9f3CXQXB5KX8jACElg3aUHdIZVOnPiOSFU3qbA8Jokd
XinovxoIJT5LgR8wGrPRtqj+NDhz7OeWq/GlCZRpY4G+RESbf3ERykDMj4vqvSdI
N0W+XvxRgyQGQ4CCqPqL8VAE+Z0U4E9kQqyg8xeMUsD9BOv//6jXoKN0kpZTX9rI
EaRrR6ByKzcf6VkK1QSM7DBvmkzbGBDyYgcKihYQpRflmcR4EJjGeiqsj9R6KN8n
dzDwQjYWkpZwD1+TJKooSK7F5r+PgruC33yUenFQyjV2/cPJnrv1IMra95szsttu
k6YJajipBAoH+VI59C/lfUj+2MSKggkpGQijwNu+E8rRah1iZqw8jbMS8xPLLjfT
70EtUJLgUlv/+hJfD7VhNVBzCdbTEjO3y91g64Lm12pd10nnPiqBrk6TqJd/61+k
fApVkka6Ad98A14BbJ0zPM3XMEjrWRfIKtKmhch97pk8Nw13DkOCzrglZthE9eLg
4fB4wXwwCmuUbpmEs0ROC3kKqli1xh5WirtcH8tmfbZyFvljnGmO0jwuOYhJUPox
t7ufL6PTRUJ/eJMbmiBK8juCjilQCYTxcZCtK28sAY09zMJaLGG+jqIzLSXbIR1T
0e+ml7eZYe1w8Asmxji3z+g4237g9cUQ6bLwoOfdxpmXtmlb7xpNvbea/K+hqP13
2qS1L1kQUa8/+z8sAoBb7E3Yi9Ne1XJ0GYEaBD8uFZUdl2SUTMlA2ie+Ipw96fm8
RHwevjmlZo2WjaAPpLacN4wH67fYbBd+aaEbhp+6/6zelWN1aKgBWHCUvzmdzyOr
AbV4xFjMpFHbiYjcyd8iZk6n4kYGVaQAXQ0apOLTr6tywyvq5nXjdQa6digOn1PM
NewylPO76TRwtTKica25oJ8cyiCH3MHjkn19zWiyjRftkvJP19jHziiphNOVou85
g/fmofw3Qz3N5d3zCZMoAl0Nl6v7FPSGO7qVXAnBXN96OrSL8jQ38n2aAjodh5p/
BuZVH0G0z0brOorieIFY4+6o1f15jZJhItIxEqSbv1teFEe4nSPIY0UhJ/GGBGzK
6r4t1CYDqTkPL5V0PYH8WNhQovjptdwcfsuP5iWiWJpz0KwR1CRoahMHrLL3GsNA
87N/FG+4gtNSHFtKGAMrhNKVbduc16Ly4AD+DerPmHkcefryVuONXILnAOY5fMmU
V9xdk3SLZnyiQq7L/11MSfQDCP7tD080rdRYSAnIN6rHS7TnNXVh6CO7QPJZredQ
7ESiYZEMnfmW52JogdM9BuihuOHaQel9Z9YeVp4kGXt7Dz7Cn4kH8qxJ+BWL3261
IsKV8UnVmsSkFIuct13VmpG0tBSRAVDUp6KhZc/kzdQ1txGJFdDPfstfZyNK0ql3
pTzfONUQQm1YWMB5agdAcmSEcoHAQ31pAO9keco0ncDMwR55UZB4cEkfu20GJmMC
WsWhF60TDjzHDd4/4vLgqONmd3vj1Xhn07tPX4cJHwH37d5VkILY90yohobrDvzt
2WdUllERlybyF7GsQqp0e41TtQ57A7IIeDEh0nfd8/h/NnW5ycAOaQDtS+jWZIw3
pyH1MoQ1kNNorgkrJLItiWR6NgCuVVKvec1XDBsb1sPgJPvZGbgorvgmrrYu7yeg
PXzQ54M9dij1LG7N87zOkcyUFm6RFXsAs739QB0s3P++a9HMgxeZhDK4aPfEpUNR
HJ3dSuk+LW7GYaIE98IJV+kRKBJ524k93L5dIL9jLrdQsvlIT/LHAHtRsOkzGIwJ
2eN57EYOwIAVHzjKGBfxrPIAyCNq7CUsf6Kx6em6iU0RclwtOwvmGNuEIfR+8N0X
NOQ3AnzOY38e4W/qWv8vRZtvg5dwyhPTcPMwxitTUCSONTM1AivuN9zoOwkTZCSR
PWKTyEUCkp+mStYrPRJxv7BTBlcC41E8TL+iOSFS/+KGcOIJLgbpOfLdpbgdVayP
Jk9ns4CwBEwaB2ruooPrpIPY2OohmdsDi8l0L+0O9hxsn6R013HHwz6E8FHYyZVd
1YtPZopEl9EMeMatQTFRDqCHcaE3Auh5IZwODTQHczkum2y15G4u27STGfQZHsy+
WJcIAXVX1r/RhmpchLJKdI5lak/yw3s9mtI7iSTEg48zmK5mN+WWeIvDIDl5HWq1
svitIMkDOOPkYbuUisFp82LtzKliysGYukI9tdg/ttwD3+hLkjPXc6mQfI4R84kT
yO2M5kxusTqsTDcJzodDZj35tLgC8BHXMv+7zSGSmGXja34QjIW/RQ0CZy3tOLsr
3aqTBhe8c8x9d+J9KPDdsdEnt8FbV3Y5bOGOCWvWv0JpA0qslblVVWYOGepHSXAU
2Y5V4jUYiRfbdo33p6nRAeRQ7y5PRcakHPpaziiGrAvq0DdRmS1rx7+DHGTbFbSK
LAc7w+yWUI0OLLmZiWjQcJ9gM8Wrb0cHDF1mtUilX083iaNO2dFYid48my1bfiC4
5YMSDlhsDgPqHkHBQo6S6eFyKzmD+0Z/fsxGY3MzL0+P5FVPTEkV7wdaORcjLk4n
007ttBMMHt8d7JPVxJ6J/3FpLn8+RX/kgJOz85Wbddde+MhM0hW5b7Q4EPZDf+7q
pBpYCmLcaURhWQFRtzJUeTC0zYSDgmz3gIWj3DqwxWBSsqrX91Hk/SjYWEfrbNrP
pEy2TBAeRA7uGWKyIZpcXP/G86bKzTb7oQTQyIMf++eDjCpL941t+2toJEkXHclX
8QPRMEkheI3Gly5qFTZIy3iFbXv09HMVaNKZ39La8n0dZPAZg1hKFsjvhYDqpueT
xs2nEEr8k9WFCqjYBqNHATlsyj0krWzih2/sOGwkKNkXQOVvmWv2v+NUYezKfff7
lTUaUmk0ybtITeF+v+iG7bOtRi0NDBYiQfWvZPO9FN2pLWupURKli5BvvoWwSbYG
nCJGdKPlON+LCfJ4MSh5TsJA0OUyhv8+tKIj6PvChzn7mDANLN0ZFceMfN3X/ITL
yoqsyjPtDg9KDL494RsZpk1vwaWW71En7T+60RqVqE/yTJ5MLtP3qdc74f6yN6Wz
Hoi+5OEfLb6sg1+aIcBQ1ZGaswhmsgklY0SmWzCJZYIdlhv4YS4cJtX+URmyI+LJ
T3crMSMtbq3ojSGUEFm4LIQv3LiPe1YVZiZP74dxijyy+F19GQvFnTK+mK5I2EM+
ykuz+QtKXO+Qo4WOie2PMchM1qRYq3i+lPOqytuaYEoNDwCoLLAUvezhLfW2cjGm
a3ygQ4LRAS3VtBZNHZKM3aNSmYJYi6fqnYGINrIj375317fwxlPU3DobEUtE+HiO
ZEnY174DNlOn1Jbh6Ty/P6jTNzSm9LnWsjUgtmjYLLEP2SvCEaZrEZ+5ANjRpF3i
Q2Q35vn5swQDoNhwJ4ubB89ijJeGHwh0yUBYG3FgFiayrIts0KfkL2XugbfZ4BhD
r3GRXuYCi0AhXLeO/8SnnXjNbbbl4VQrQfmhMrBHfOC/VErZWDZXgiQOEEoPglNG
tUCQORe1SEyHKMDXgCfXeYKealRkOe3UBZ33wrifUqWYRNogqCnOI80X64CMpe40
4zMLAEyqllYtz7hWTHC1OPSI8mt8e07tmnNGCkJvap0co4xDKPw8yHFmw22tM5+3
WZCWFsmnOVrC37rj2wxdn92DlbpTjyH2sQc9PI5aCZLagB4eXa30HZj1WYOilotV
AgbeTNH7brwTXrcp/BoGlAwccFijbK8vv69Sq4Qj0yG3k0T+jY6QO1sOWrsodsL8
w721NMzkz8jOS5P2pGchEYLkW21sFwzT7U3BWSFAWz0vlL+TXNjdbEq4F01DoFhf
i/Gi/I6gTNGmcebcHyfrCo/4RzTHDupDc6CjBF6wR71EvLJ/r6Y9EZPrys7xj4D+
76/Vr6UksfdC3tn6RH9xmpdgbPh+9m89IFak5D0TFqPbOxSQMCQCySwCgd32Jtsa
zXxaM1tDY5BRVKyDi0MCIPe/6rCdEyJWOg/umHsgFSmXrStd3jl0qHFsd8dun0AC
XWllUsKGvtoIhg2U5jUF/pWGgdSA8jXYp5r4/xA3WW19u/Uf6iSe86/ZE/lqdNEL
OGWF8fJkjoEFl18Ojxx2EmZVJ62uDSG8MVxmHTAXAQQfpHtCRo8xHMk/wHiQHvD7
+z9E9vH36+DwUsvFVQilXZx7PwfpwKDB6s2DqheK+dnQCLF8UcSKXSHQJ9LKoKs4
gatW/wxDFs0ATgekNT6tTcZvxmH8cby55WyAopr5Yk2WalktjUh8tqDrPwofxS3c
pp9b6QIR/o2zjB/2QtOhnDgPdq42sQhYOwYjDVsLWCOo39WJF1eiHQzdpjKzNK1g
/L2KwSTCeaVoHphsiTNUGO7SLlTgDA6jJucS/qQw28vXJL0OO3gLDFFGWiasO1Vm
xdiXYv+8U3r63C0FtGKNHccBjii02GZPMsagVE7OVFAPLUU56GRzUibNRSkm7V4c
TMVLeDjKKX+L2avv/3Qtvf5uNm4GHhm5fkWItEE4e5yU40Q9Zcc/Vh+G6vqRka1d
TLXkB89gZfr5kGPeaZ6Tfqlv5xRCTyA8Fh0atoyCaKGzRgx+2M2rAeA4sQuZO2vn
NwcsJG7d0df7+uY0xBEY7b1QrzOiKBpkaXV4e1JhxinCvJr1sB6EzNcHMqKxFkl4
Zo11L8tHcJbZVUnHhIJF6KYKhaZgH6dptvDvsBzNqyA6cd85b7v6AElpw37KtuJk
EMAXBTdGKHaT142gOrFrMZXd6/qmyMo/yyMnmpsyxedYIHp+IqIRh3lFe6JVi2BF
zbjEOEjWpH0dxQtcKfsc6evbRz45O7xQ74G53Ol1hkTwYLkAdsq26sVv6B8PlVxU
9MjTmrKGTGoprNh1SLamkbMBFB2HaWnNbr0YYMxfPHDvIeA0NHJuV0rftUSrqvNn
QlQxdHkF/AZfoSc4gdjJPpJY36o5BDZvij0l+clVtGGyLTGlsoZs0wUP/6e92LdD
aAXIVy1KJGiJt0zJcUC7QHgz0jeIJ78+wpobjoSjLDBAD0NY2w9M4Zfw4bIEf4MG
IlJD/sfpJi4E74ZigwpxcsOZFmdZ+KDz4OfDK5Msdc9+bm3mSrILjfCfT5ORT4a1
004K7WD1wdOw+jK/tmCSRYo2uBiipZsuUe0ge9U5zHW+VCdYthuGKDNO+Gxho5Mz
46FcHvEDe5SNE96dtsY55CeGimBAJUFNIegfKF0Rm33CKJS+FVNrNbG4lAVAb0wg
FK2ABcvEW41jGRQUdbWeq24NZqKRo8xoTz3wV5pqS0wiKKO5FMotPUAIP7rya4AJ
0ashtuypV/QlwHjmmxeoXKuOwEkgIx9B9hOyXkSNn4C76dlVytOwmMD8EDAPylCq
O4JWp2aMU/1bKDeJqca2YVmkniMz5ju9AY50cNJfOZBLbM5wzCjflnK38krqDnKD
CmZUTm6nG0/7HoXGYK5yvjOpCEujoQMgL9AojqUn+VBZeDMrrg/fd/q9jxHORkVa
fzkZi/Bnt3JnfiYyngiu4Bf6eMKPYgcPVuwwwggHtWkwP/f3YcOb7fdb0kWAI6d1
w75vwZm0aMOuX7/9tMoCmqzIQe6wacNzu9EhE6axPn92x9TisKjlzpzVH/TCLhj/
gnV5N/xD1aMzo6n5SPDPH0+xTcva5LDcPgwlpDxM3bz/6lO0sOG/+CHFXx1MVo3z
2gdtJVya2kCeP9ZTtmG5+3Jjj9zdqwmdPTsjCHr8GPiCwHmvAjbWJlpm594kb/uX
ok0HopUT16mo4Sde0T/66AhEBOSXm6RFJUdZS96pUXksb+Lvx59ml4bwNI/fLy03
CXWm/pHxU6RYlB8TBf2raw+JP8AAMhCR5zMW8dslOtXNo+w+fJr0Qv2SzCtAYYPy
BRyhsM7t2ri6+Hjo0fFNZAeQUpVxR3YOcuW3fJ1TmNF4l2YIztquqvBpms3zw6gq
yq6W+x9cxDQLpPe7DJTmdzZxZGoY0250KzOoyTDETof2TjgFFTWEpPWBq1uaRave
BlORvwYmO3wCwcep/4SP/imUzKlTUNEek3otEIU2xYyHzym6W1XxUt6ehmoaLt5E
gaKVeRDn/F/N8RwXuZygiGBaVXjTswihAq1ODDQBthgT3gIS7ROCDSP8Uiq18d/w
ZZTcDKXcraNke9QBHt7g8B0EkaqKdlm4YArCzvMZRe5ykkSka0CISiZ91WMX4X5k
+QpUaxqxW+PvPfuBNAsbd52+koW4gaFcPEn+Vl/pxdTmx0rtpAZlB0uGTstLnLP/
8m74TSIHTwWbcqCntuYJA5n+hD7AtL3qKPMoW+xs+jCoHNHTAI42ds0H1s4VtGgy
jhvjrOh7dLHQh9bFVRhaFjuaLr7sNKD4jcFBsu4Bjr8SPL5aEOguIDGeRR3dv3th
BlnI/3H40eBlWtQPX8FtfCF8L3CzhFmN8LNA1UqveU5os9XhdA8Sj60NBz1rvB7h
HSNue12ew3nQMHDbRAhbnRY+CAFtHRhxK56hhQLM/oHte2/1KttgiS1KQ2CnIDlF
h2ibCSbw+4n5XFdXen3oxh362UZ82VRfZiAuseujMgeG5P3ePI81wTg9RN+HU6WM
SyvI1u78b4MQd+Xus2AOxKOFFZOe0CeiyHImbqlsH+2aWpvVg3fpCpjfTKqK4n+c
Hq8T7v7T+IBpazG/W+LhXTgaZ2lfQTnizCGS/iDoGRboxmVFXl6AxOQR+npP4ghd
qgCtisyH1eiseIRjzdCZ1Ylip6/ijBL29gmk2SasagKpPRlZmYD3+SaBc1yWGqFq
Akj2luhOEEHrNKhocfdhvIZN5c+TGaZCIv1zuIZbHhIj44qaHXV0lb6iwqIQMo33
jNb12WCpwUpw+g66elNAee6J79UkQjqX2TAflAREZWvW8xdMzEe/nEL2LLLwj2Tr
7WL/B6zR7i5QL/BiQ2/gW997uctYXuxf1vwJ/NGbsDr/eBUA3wT2U6fjQkLdB1F8
tK4zzvD2DvaPkZmcG6I8IYS3fZ3G9qr22I1kj9ObtlaNp+a2Ggy4z//0y+MCkMZq
FFx3U4enn0a4reA3ChiUL/8SxsQ124DNyfkgloyZCx5tbSFxW8ljgc4JLpFfFIco
KxDpbFDMlKIj96eYEKMgwRFzaeq1Cc/rNJHq+/eoPpHS9/f2xav3x+H+W8lrn37h
C+GDFU8gNpGSS/1ayB39sGHCjhRSSWcAfpckA9e30YrmTBSvxo9BBt6qDlBcHpeM
CKO/JD0LyMs5hSAsvV6darOdEs7bJjFWXcwrHsvQi9vQs7PcCQbY8OgeQey2qKsK
rwFXo5qTKdia6roLhd+6GlZOxNTL2kdmKFU9wx9CBoyv1iliNnGXVuj/s0odtFl2
0uJDTWSq8BH0/SmsUFEjGPepxcx1QuTFQWq3SEE92wg4d6YyBoqBneHyctRzFMiJ
jK8qONGerdv6jBTMTZ/GpkL6NsF/0Zrw6iyXmCdNZjbCuAnIQNX9uLv0XmQrSESG
aC4kGhrCPBCN2+Zxn9rhI0lyXnSqic2M85e77cqJgFqLEQAyII/DHl0XeyxYbvhA
xvjODP5LztWM6IV3Dr0bmGI2gAbGUICUOoZlvMafFN+ZRoInaUxlQcLnDVijV471
yEZqB6NPPsGuHtVF+4CrxwNOY//N3uFJKqY+opSqJmSJ1a5lpyUCwBz0p79ix0jK
5RzjM9yhdYPub3vbbs2JNWvXJZMAgnEfKYPJvibNXvk96Y6wDNLxMP5cLHR5GYsa
3o/JNdJXE/az2eCWSBKTgSPhZjRRgJzTJLdY6BFYL0KtDidJ05YFtan8RTvYkQ2j
ew9mL6qGWii7H0kHzXoj9qjqgwxdgEJC+WgW9z4jY+yJUDPWnv/4ieV4XigJH3IV
o8DKRTQgeU7fdbgvKaOhuIHsORQEIxEWqfM3x3oMBt2DwUsu88f9QOv1mV6RKcGv
oMVfkmGGNNikkyEc+sTOkdu4oasgX4os+9nKkLK07KX6hbIi+G1ohIgaF1Aj6aOL
j1R9SBTI9EWYf89uepk1tls6sET02XAWmDlAYN8YUYIMGlhs9ggCodQt5O0Zu9Gc
+qcheXhSYO1C3ZzJ9BjuGvGwaDArh1gIE5zneLEErNmw/vsjXoLS0Oj913jJ/NM0
VEF3vyaGBWuZaGGYs0y6lSYqtb+LQ71DV1+7FfxJfQLEPsOiGdVEudk/odrEmUoq
xYJ6MmcbzmWpcSAZIyL8ZhhF5/iUKq0N8oSjug11QeMS93xSyje5zVj0/dMk0y8z
9pGbx+qUY7aIlaFO6lvfj3/heOs6mjZtzVJjhCMhtoIg+wAOMm1jy5biujCMztgs
4FiNxEvFA7+pTkffypS+tq6tEe8iu9aZvknrXE3/axkNSbK9+cGugfry8llGtUmg
khM/sPfRPtX6bsVxCwPvHc3xgTqxSZtYkn+jznyIjycn6Z8GAeMnROx9vOgfrK3a
n7YKYyfTTmrKIXnufuEt/N9mwi5kjasaxvAmqcKPy+QkHr0Jyf7lebQMfnfO/9Un
6F2treBkvnOhnIB5G+V989+N/8mclXDMmiUddm4bGr0XT1Ij54PEC8RA4qzdfj8f
IQA/X+aw7ykBXaBSf9jqzOAmjbnlGaweiwenW4iEsyzAWbZ6SEcJFkTpfwv+274V
BxhBXsA7Yf/UpL/8pnbRja9jxmue5uv0d2ac0Bc/gQy3dpTzx06Al6T8fQWJRvVM
nJlIWW1ge8VfPiBI4H8zdbVq8/Rn0l5oHI5l6cHDuMKnjD6eB3aJEa7iufj41mw7
RcBqapeh/OBvbHjM2YPp1euk+PY4Jgk5rEDP7+pcpR02ZsD1GHh/GNlYRjjxO+uB
ityTsKLsMNvgOSNU9BPTu65YLCEtunvTKzjjnj1T5qiTG77EjznnXgU1HwAG2OIb
+lOOzTpc5Gnxol+HI2Ap+SDMqntvDYrU5PUiSKEjPIKa8JT16BfXh0VW+4ztAMoV
VsL7pLIm44XA2IRYwPxLLIpFeb678UVrfQKVeJcBwbESdPKdS+osuG0VmmrwfeTx
wEgFIPOoFxkBN+O2DwNKQtLRqRTZORN6KR+QEovpmutCzRVH4N18AnZlhaAwytVJ
xd/4zleQksptV8VLBABL/o3/JRBZae1N3yYdowvXyUSW082BZZpEjalIL0k4cWKH
ucvTe2JZiB5nkN8y7gDqLd2/eNiN89YcITGp1qBt3umWoRptHevu0yasK/GR51Wp
JeJoTNXeVkOuA2YB/uE21MIX3i4sP9q6XEQhF8q712KxgfQ8uqAQWJ1x2hm7MOru
NysID4Qv5IUqHnx5jiAa+R3D8Ih7er6/R7eE5SD6ErIv+20ceOKmWIipwHGzQLqC
tnrlPKlB16vpVj0I8rJ5VBVAd4RfOPJIMTIKdVeftUiUV/ZMue7YNEkURX6cZHRF
BezINfjCXFUsZzP3TY0zOS4Z4cSOfhMVhcaQUvlfUVZPypCiUNE6GD+nsj+14W/X
g2W8u+DFDn2E/QQnIpXnRyTjBWeStNDTu1l6YtJYDWYnOtNI12FQmtb2fAsmU5yh
8jO0S4XzG0UrLPZ6JNbGr+B5Str34kikJSLKNtHOt7hwYMjz1hnW0D7PD0tR2hho
S+2/4Bw5EyFQyet4Xir3/UwV38C6T3Ow3dF/ko4sfH1FGv9uadG6ZnV9seu9PqRz
FpizRz7E9ranRsjPITWpdmMFMlOrc335ywCBSMC5W333WLNpc+q1412y9vbcMj2D
jX0ItuOnibdPWZol8ZD6FSDNNNh4HzqKxu+Dm7yRiJPsi25K0r47k3bucqt5IAOR
0cewZMncBzQrXBhOHr06VPO0GB+n+kpd73sCiQbG81bOjyVWBAk/EW1n2jfS6Nfh
vjX54d5T/xL7mPirBz+zvOz3kvz86i3lsLcOePLBPpnckmfAvFh+o92YX4EnSz0V
gMYYMFAMvUHGgfm7xsAPLWODbSSTQGfMdMug7MYQHWQqnNdEMDQ4FirqN0wLRbUx
I3+I6d6KPUSz9SiT7s1Prod6n8gdbb9ckWtNh7BeMW9tpqnFql5YIUiAQlvWyuTn
PB2PNKMaUyEDIMdL2eVdiExup7MnkEjgtrczp8x/Gz666RqrJ/bLMeTKc92YltzQ
NWQWEyC7bsI53vHQnhqSo3M+g9JvVKjriOgqrpceRcwzBwAhrI7NTkfcWj//CU6u
C+BsaRlKKPPUIAt5Njg/ldw03qniu1GkXD+bk0qUVTxnCjnCP8INEJfvAwvxWTh9
8s5sQE8xLiO3FAYu5SFnMSg26h1WSl9+3tQ3gB5PSNRs4YQoY1mL/wbrzDHkk/FP
87QBN3c8ixxSFtwI0HWi6aomP+HEsI4eEamvcpVYl2kq08/p4USYJu4nVXZf+FBz
cZuaVRvXK4UegYcKnMSBguVXRgSOqbZ/DKgcqkTo3ayOQuUpFDsozaROF9HEmGHV
4zW3LI4mTA/FDf9RnfrQxdQlmKu136fu1ym9INrS7JjH2yTVfTQaUCCTzeGgXb7G
PM13obVo3UDYZwmQJaKIMGAd41S7+s+harYGr3s1OEQdtdifDJ0gR9y8KFICqRQe
xCeSN6qjVksijmW8+QMlY9DGpJMMAsorpnHRQFbWhlmliOzSDWJdq3N5b/zCf+60
7uooYlhrdXcQnjlhio2rksdhy616AOFxidsuHnI5L/D7jq2tKxWmX7tecOw3/0C7
j1Xjo2K+8eUDPPeC72GB3Mq32pqVXVYJ63LM4vcCtGe1+hNN6Hkojb2JolKGXTpz
XTqGbBh3q44Mlw23sEL4Eh3zxtTt/tCFJT8UH1gpt+6yBNmnkb7NoL9Q9A2HltSf
R/LrjikrwmXNvy8j1QWQ/qo80NbwAgGfupc/tqW8QL6l2JDDXVEWLU8rS6nkX0aH
MW7aGA38IKxSY/O0mPZNLz6tSXOoCu6yHC9c0yRgYK8B9FkEF5Bfh/NQ2Bm4zNrr
7K/B09s2UPQt3vcrnuya9Z6Oj7Cfze5bSsIcuKv2TyvzYuWLBKbADsph7XDqyRrV
KW2PkPRLczFBckJ2HGNlBq3BepIcrnd/T1JXE+nRUEz5gaUbdpGdYAqDi13S5g0I
MhgCvXr/NxmsKSJl1OIlQMPQCq3hGwKC72LaCr2SHf7n9tsr9F2Zrs+80iAVhZA+
ce8KL5ikMxQmNqNDxGLT8Za+c1SoNK9uis9t0Xi2pbdGjsBc7KZgLCrPYEyBNwZ2
aFaJRgVBdg3v4ooTdykuBEHPl/67WKWVp+KbOo1ewNtU9JsJeXkt3zKoT4qnag2m
nk2kO2PteFsDZKgTgUaLobF9YdbJWUjrY5xtz706hJrJu77j4XEA/vb1rvhkJ+SH
fWnMCR9OGh6nV5OR2r73aHqoKH1nn1X7mTvpqB9TMwQYNhlMIGHqzb7jZvkI8U+h
aZsIugaECPXrJ8Pq758cVuVO6tNEJpJBpOYZ4NTkY+rRSnHVtwtzUmW693lqWOST
hGcL7THDK5o5aHOD88gWrrGLM1p4Yt9KFLFyMHxuXziizPghZuOVdkPkmsEY2mv3
e8ggyykU/yMrUSAJd5FR59LVnwIGezZ+ZEaOSrwiYDPwbE5k4uKGaSa9UjDYqbRq
M+vOy6fjnWisAd/XPbODaGecgPor91xy/Fknzv+tTDQhl3MFTY61Yt+jHF/pCrbV
29nAcj+b8BD81ymy99EAeU5sDb2ltgyFdaD5FElGCHh8sK6tuC3KG0tfiCMd7ueF
yV8fjIapfG2qG9AQqPU2PgUDr/67Kr45djTo0cxrY/AgC5bihXwAgIo2nJlQ1ihX
UxJ6OqsssX9pxxDOCJnyZ/8IsMBVJmQANnqwCb2a+rfzoFXVtoNoOmwdYkQjS912
tkr+iOmfXuTbT9hMYni2HQF08AF4ZG3WWLM7oyzb8Z0sXt18MJI46tI0ixgOnJcX
JZvcHVtS3FwmnHprGWIDcXHAszN0SjDskwmsoDMQf/o8rNnArr3yvPmVBQvaqUlz
AMmUvxSeM5FMGTQG8c/NvEPP4MWFQWxB2ceCXbat0Ce8vW5E1XeL0ms456J8MToA
f4rtKI6KXTN4exROPHnXuQx/KYGLrP4awc6hBwUEiCsZvJhvg2QdNas2YiId4x34
fzlvjjy/GV8xXkz0jUhk6uScLT35ACV8fZP8dCI8wA4by9/dhLkg8zbQmKolF43t
b5c8W40lG9ImH335m0xY6GwAUIK0KJCTFO2oKu7d9qmWas6F3hAG9XMFs8Qx/bXT
n2uD78RI+QJF/hFwx80sE/M9xhb3Jj9thgMrZlz42kOtePtpSJt8yCcqKYEQaPPZ
99xnpf9aAnEG0E1o3hKOlsoBO7MpdX2z5W1uNEzX/ysjvzvSyU2XKFDBoHKjpXIr
kTc/7G/RSxmhq6K5TbvufhBZMgEhW5HzCYZ8SwvfQqyOojttkCKX96HJ1kgoSNlq
7CLuQlli8sBIeOBOxZ+L9gPR4nPQyILFU9HP9I4Xik8nVWAnoPcI7kW63lTkJdT3
1CUagR6NGqtOutvDgQoLMBCAFnlz1SIYhFWxibjURMqAhG0pfWD//C0RXXtcpu5S
BOCO1ZIx4h1mqGlq5ja9oyMxXgX2RT0bSSq9KpDCXpvxOpkv5bioOABihD/p+M79
V2wUljkYfR5W4oL2UvqOe9klAHzXEMl40Tkz59lKC916DuL1JIa9lQTti70zlbxt
gBw5mt+NgyCebzLtMCdSLKRaYws4qI4imCZqVUG38F9eGYJgNDj94C97O4gQDaGX
ogYMAQvxYwMG40tFBAkGGzYSnLZTJJ/zUEkZp3s8tRMdyxIFpM7GH/52xRrICwfx
QcY2ZiT86gc0354zlsZyRCsW+atyOO05M5ddp8iiwpX09EERpSoEUep0fSSicBfB
yxFQ7gdRNIK/k69qxFFQix01yVzl83jR6SJ70pjjkQLt+h9kg5dE5zdt+dKuNuMw
PKPJR2lUnZjvnGP0GdP06gVBk5RpxK/jCf90e2sX96oL1xhgFf4TT9vZVujSSqvU
S1Nt4jZVfCCmVybyYgnNZOSzVMYL6IhCrpgaekor65NwDIHlrrdkgvIPdq4oakxK
ChANcldHJdIaiLAoWjMRneHJJEoyiAul4yM4xdWunliGkjewo5fj7tT+EalbaFkT
bEpoE9jXPiUeR8nhq2g0a+W8nypipaZEUorwFkJwyEh4dTLlc9sng2tbd2wBknLj
HbNLnJvOLlqgxYAYNQGdKrPy2ZEXlOA3L4Ema5VMlh8dzXBfdHwOK6+8TTD63Omj
th2wPvTmnJqDtdo/JIAI1XZIao7Wx5MlVmVEkVXCR5/eWJuj32L1R0F1mIDaEhgb
nmdzgjWu+aMf0T91bOojlFosIxfhEghSZE3UxwNj+/zabQQQPUIoRITR//7Lyc5w
NPJnc9tSYCW3RPJ0LZkzvSc0ltPKhJaLPzK+O5jA60QDc0ISFog8sJ7kTUB3Kqi5
LPOXO33Bh9w/V0yV+yLWgGls8dUireAqJq+FEpPU+u7aUguc7rQaXR0b8VTbaxph
05bk2QdHPMQc/VACE1Zh6I8+oz1G3ipQ4rhSAx6PfpaKQRoMZZLH+gvEAcM5nTnq
YynrH3PJG3rOkXIIT0ks3F9SpZF+UBX9w9uqRsBxsCEtRtXCZSBpLvB1Vy1lD5+n
fqVD8JtKYmtMrtxjy4eQFK1r/2bsZJhTjaI9lgx3w6rqszdfoqOrJI5ONw68xnXz
q8lEeJ/PJbbFpzc/tGfm+esX9dlAjDuMDFOsrFj2qtQo2Q0/or8BOhp79aAYg9QN
MiGyIB/eqNqv7cXo+eR8lg18FfYMl7zX/vx78CHaePe99U9Bfa66d0sVGBiuNdZc
/0ayxC4f/Gksn+ZpUShaPAxM75ixi0GauxG13YRbXWzlwJ0KVUNPP4UYJBIiACVQ
aZGfDAI11MrgEVt0KU2BiOZmzgWBci3dLE2ZxkZA09lrDC1YSwug8f6t5aCgqOK2
QtmWJ1To9UZUNJlYO3mFKUALZadeVUw1g9weUJMrKB61PLBB/0Ek1/iz3kr720Xo
XN3HnTMxkmKojWAx8aulajkgjJOXVw/TsHiZ77eleK6Fm8gZBy0NzzyBXqbyfzFt
3REulfv+pOce8sV8dEZKllpH2C8A3oCfYbvOj+awDYT/+Vme6tFvcxHL55QuK8Qq
xrdnUYU1olky9WR5UIVgTOrlC6sX0294ykT4CdrIZ9p27EbKiEO2tODbozDI1cMN
KHPvqS4PRMctUImV2wcVooZEu9nlEM2RHwE9xDGPTAdxqOARKOFwDpqS4ppjJYCU
6FT+FxzAQnipfVEp1v6jRZtXKxMKPM+IcBdd/Osv+fS1U90mcPsGAv5AEng7nzf5
fLPe9i45B6Fv2xrry8G1t4jVoCsiumjAD42Eg9ts/ttKD7YyoY0HlKEKvhIBYUgo
ruSnR/YAYcDYWwESVCy9DdBB2PbRv85FazZw+lBayLKWMPBDpiWqBroOyf+uoZ2H
zJp1lyPFDddECIYwafebtd9xQ2xM3boxAA1MuDrH0We1OJo7hL/WCU9xsCYyDUMM
cXSodmO+wj4YbPOOclGTuUCExnR3IoabwvKc8udHElNxKa3RtKO/TjiG0mKnWnFZ
+Kq6ZntmBaQtcccNengfevMwaEbp1AIv/RZSk0N8FTWfRIhAjfaqzkMlPTYCMM4h
9WhsNTM+qaj7WU/6zYDQ+uiW0LJyLSwR4TxKQWcE3/v8EU9CB+tf3+gkcn9r7tZ0
HhvrEzpbdd6leb8G31h/w2P2/mkAOxqY9eJqxYO/G+9AuFTiRTxDPPxaFzk3F1O5
LtjPEpwtu0MGfI0z0Ll13h0ljq66GJGc7W5rprqBty+G7j1JtnO2iuixqOed99vE
MHOLsXFIbC1Q90nqIL7SbCj7kG44gLKS4cNfiJwXHnRj0daEd27GjYmL5jg77qxf
h1VMby+nv7lgc017cmetXp1zM/YVu0GfvJnXW5UHLycnf+VoPY1fFLMVu+lxZpb5
Is46tgzX71RLJyH0Ht7RHagRu+ccBw1N+/JmEV+XD0HTQBa5w0uT3De1ZNDChZ1b
9QQFtLmG0DeGay9MvWKHBqswm0bWLtKHAajVq0975LsUSzrOq5Rj9rIrVEec1IpS
NgAhd0YuwipxTWnjDKzTC3qRDyqZzhMPmLxBp/HlNRtZgOKKWpLtTkJSad/qJEk5
VQfo7NR2VZcL8iUHbWWOC+uxdxGDk9GieUSB9vn5xUlbCz3f/SV5St+L7aEV01XL
GGdlWYw/FqvjW9AsHqbyBvcx/d0vmolIWaaXh4mU7N/RtRHO6eFHsqfWyzD/KkKF
Gr91g3p2e2JopSsrYSyyo8Jg5zX1rvClB2rY5O6P9z9MZqrz/oFDjnLtHjnCYTQL
TSVUMWTNLyKQ2RYn7vOXwNAAfTgBCGmkhzz4AJU2ry7j4ByKjG+xdTx8qk9vI64W
Yxc5z2M4Sh1O/QF41fQCSqXyYf7ECCPh42Ji7TRFqSHxr/CBYDBpWrldkBUWD+2O
r4UfaycMphy04VCAZTIlQC2V37ppgM9JaJmam0FtkWjYrJoZDScsF4HhQ1g184oc
bEVw/a5rRcx/i+Z+U7nEu8tQFPSyT/wVZnl3zBG8mSwm4PSOAG+p3lvaVRPs0HuU
/jzEHFHspCizodhU7QY/oDCRB0HVTSfhPcfX+C01CMJ+OLwlq2CKXKN3aivIPAn4
V5UZ+1m0UE/fORmDoT3m0H+qeYT8Mvevok3+v0edlYNnaSQq0fiokkoYu3gqR5V+
bSyyZvaL3KlSj0cpJhbizdNnZoix2xZLVJnmwfG84NKeqauCAOT5MlWD5nIZd38t
uLuTArNzGAV9/MeagOuNJjWgQ1/ie4c8AJbUY8Nao+RtcsxELRxW+SIXCUHkIy6O
kIYg6vZ1HIcRKdBroOrEdYJKsl7lekw077BibTObJuar35pKwD2NMLKvF4f/M0Jb
Y3T2QOikcbF5P8EeHlRNtj7dDBA4TFrxGt+l1CyzbGmZNaE5sQ1HQUqLQoShFA60
fdYF+u4BJPWvAKDpAo//xVt4N3oKBaOhcOveWblvMQrSXBZBv05tPMKOGO7lNVfU
DsNBPVq/gX0ICuAlQJA5LCnxipIADwZRPKuMySYp6/cS4Cs8K0idvAi0e3zesWqE
sj4LuIG2TX3HUDnSt4zkz/Vn64g1QSYOFqW/hNwDE6PzRX7+Ws1akuEtKQGX0dQu
CflX73aXSgnZlxgV1f1IBAloGJlsYBquerGBJh29ODSuEjTRyJhnMZCM0D96oPJq
m6vTCrl3BQLBTcUbFRD75Mz0/4lRPtsiGX22IzDUGiQJBuozD7dHmIpbLDZFZf5r
mvhB0TYONbD4PYvo/B8gnw3I8AvlTU99HSh+evk500BX+pu3H+8DsSj5QvsQix1E
2pYV7doItIG4Pwjp7RrFEeiyJLq1fIhdu4yj8YhAAxIy1eS6ah4xm7ArMnT95SYo
i7pRXEH1IUntj17y267OCkYLQxakRO8HnOxtBzIUlUy9ktVCE05zG4dn0sY/2dxK
CFQsZPWoYgcYDoKZ55VFRSexegfPUWOnxse8eBdTLXaESNdOF6ZHMZge95UndO0f
jOkjWqGdnYsZFGpFLuW4CBcXIt2dtUKKZsqviin0P8/exluNJBQHhsObbJQHtLeH
nOnrvrSJy+tnreRlC4RkmPReZBtOphUIXmBRDyI6/U0CBCtRkJGSYFfb+oOJNFeS
ygxI/KQhQA7biJgu6YJ2U1+tO+pSyKicVWYz4F695JYQy37vKq9jU3gC6r+yjrjb
8GdOxqrFDGbZo80xhsvWdrbRgv7INBXwFk2bJahli/zt+J6//eaxx5cbnd8C88jq
1e92Dzmtm5WG3MWlc3fd1nZ7A2ptFgDKS+9bqtSpBWxOvMNY281bnoAXGaafFrmj
jTk7l8/+e4sWu5XYNpar1Bjq2mSMzts6Iub3TLovE9V9JgvYYkpAipTNKeASH6+I
1mBVaZDV3lmjXGyjBEsPPaEIjN+r0W0qhyLqvPjHK111SZE2FtIvI64UD6riX00b
xaDET5J4YFxogLlawVJMwq0yHtGQHvA2FDAFJ2v98+YbcrYeWytbW4WlhceybTyR
y1rQqiuOD9EdF5XrwYH+5Aljr7ukiTPMG42ueq+XGKn/t52PtQJ907PxCysvFVXG
X31yYoZcMD0HKi5D3awA9fRK+5tV6GJMWhQzHZq4EQ9ixRGvkLTdKDUUqH7DFxlt
fS5AYnRK/YqeJqifAoNQj5mUNNg8Xd6DYWAZQCRYlmHHrn9DMWLUhx6kedvPJ8z3
N39q3LIMnHlmHNi8fSLz7TTd58cN/+WyPEq6eJ2SbESopAyOdF8sO7RBbXFlHnyx
4IZfxc51G819WvMEcKijwP4Hn68kKFvwVLnls+gktpNCOnGqkBw1jOmecYNL6mBO
nmm3AiIR25JWgVA13/XP+CHxiHF9aFK1aIBttXi51vhqhfWggCM4ZWH45+ZhVhbX
iDb+eEn5LMEGAH/eG376umbo0U64EcWJysiMVP3rMr1F7EQs6wOi2qmWeWPaNLYW
yfKpMnI6iT6KHFwPMfJl8jsfPJTBz1E62f9S4EYUlSA5QtMpcw/aTdacMo891gEN
vBgVmvJq/jOncsJBZogv1b0+NNEnO9JbqRmdiELyJ+U9dp5iF/gZ0lzrgSmuBqOp
PMAzgDvzUoDk5QKdYX6rQ1c1RFDvJUUnwbXhmr6PoJ/0VL2+06YKGRA1lrNg5G+K
YvxCzgBXL+c4j6tiI9GelbPjZz2b+NcYwWnchiRL333MskYG1KsnL0ZoxXMnerQq
XTXU0noeBWoGUb5t5cAZtl1UlzYRu1v2cEfUnAG2//OW+ciyrzAi8k2AdWgy7s0W
LVHbGTyXSFt+nend3Erths3Zs20BfjoXgXvekzVnM+g8luanw/nRwV7IdS887gH9
j6clpn7Gfm2affu1V5qEP09TGRxRJPMSWcvIQgN+CEUErvspS3bEmXuY9zFBa3Tl
CUADPqmTzSC1PHeSe5h9GBQF7fKApDgN/8e4ygSSjqhmF+CuG68Cci2/BI/As328
NNIlYhoOeLCxlZ49Ldsogp7VRaic/Mj0o/rsfjGDC92fG70Su/8i92+KzGxc5Cyc
+rOcOgNyIusMAO+5mPIavEL7Yynodz7zzbK7sAyU3DTDjwjR9BoTTy3c277AfuFn
YsttaRri8zDxTLDwXgEtmrZbLTL47qc7h0r28YGPDnhwnFkROOOQoc8i/60sPmrN
P5PmiNa/gsb/X5KurHa1x3swyMMCjYxABy0KZyCEs1JaLz/C7vaZDk17JFcNglQ2
+DLQgEwTY8yuLi/PNd//+GpDIFnL2LiPxKi04sNXHEKRnIzNcD5wqptnNIyj7r60
55DUC5k0CXz5goGfF9/EQecOHD+5kv1FywXLYcKRFWl7xBzPEyYrhxP6ZEagWxpK
JixKd6820vlHry3EPbPviNl4WrAoREaH134nqn9N+2AiYJCh7siTA0qjo5badBW0
RjFqADcwvQzLu1YUyXmI1OdPTEOnUxLe5gLbScCfTuczCnqn9XgjbGfibX99om7g
R7EM+gzWDnFOWZ+HvIFuyw1VL7U3p7LijZv5AOfswG6LM2j2BW1MQcDlTXm2aO+D
QiKx2A/Rcc+aSqViAPafBKXplGaW8wo1Vb6qZ2aX/mLxeMdU4UVZtvExb7lzpnlr
bZ35/YjFfIbb9Mx9GoHqbd1u/XxLhiXr1IkEyC8gaH1s0dJexz/HqiErq0z9xkFK
6cwG3uwBNMK95L3NUq38q3dW7RRnxNGe4pLqjnJ337NenYQaKrAAXTJkP4iaEMHE
Wsu+GfKQAvZ70RCthwBfmPGAi4Z/wwo9kFyo8hsJXpd3wFlMwFju1RIWFKvKvyLl
p0ttgU/I/Tles4NzQ22h20JUciZNugGmAOkG2Ce+MQAHk3XyvsyhHpHMigtYifpC
eCsDv/Q9OyEz5/3XLLYBj0eWKIL0X4LKR8L/ow9/AjroAgnQKcxpvLaNfRsgWvka
KY+DCmR5Ua/G70zFkUex6+L1HN1idW0znpgbDXhVisymvW18GEWX10kgojdYTJ+X
fike9a+biAdMM42hviJEYB4e5/gz9/nROX1DiZfZpmMSy3OPsyDdaOMiFwom1i87
PwVZvJIuvEvYrsZ8pd0U4t0yjJ9lvx0UdtIW0scwlWf8KQeAcEDeT4gdlFtBppbM
4COdfaHys+mwlZZqOEe+4IGNVr5EbLJ/7ycAbAbKchmiiTh5VRQ/G24ozM4eawF6
upVZUFkTsOgX6tk7KdsqFMAh4s4DAhMyXA/ugaiMydRSCy6AwncXR00gctps+Yem
79dwxujIC+0WTR8S1YT6apDfUa0TErB48z1AI1GnObpseFtHSGt5Qpit4EDVrZod
bMhTwg4NaGygXCmN8aYMZQAzZDNgSJF+OxluFccDkZCHSxMErJ3ZMIRzTPUbOwC1
C/69Ga467FnGrhnl+e8LxtgQsKLdLAETmLBwlbUp6ddPkWDIzprPzGQ5j+Qer77B
RW8mvqa6FdHNoEJa0TYhX11K1BWONYg58coOFRmzT9ZseclkSyOFB2tHD+z1g7z2
/pN8wiaxf88bzefWAdhCHKUumoSvWmG3PuEj+eq8I1P3gWE8UvWGpwK7M4re9sVV
yvVXA0q1ntTfXkJGmu20crHiwHnLchyUn+0AMfKqvott/esyTEE1yM8CRnrmPHRp
LYhBttUfsLhRVqJTbSAhbC2PXyLtwIz57569S5Fp1Kx4WLKbDXc7yotPHBPejfNU
J4iqIkx0uiJLRX9rHSJeBEsuhjX92v/8eTHtJJbbbGCqcqwsOK6n/xkF+fZHPGWZ
YZoh/dyyl9GAcGNF7U63RmCeNYG/FwjDv2t4EJZRLKyFaOzIa+cdaG96xB1+zC1J
nPLJL7n4F5Cm1s0Z6ti9RgKd1pskZKcFjJ+ndYiGXi+fVENga6lr64PHUKT1AdjQ
vJrZAfCfRkeiKEAB10b2TZjXKWp7fd2KtH6enlHrDzPHedxLvTCbS+sHLKzFcodQ
SwyUtf8r3ONGcNlphhfXYVbOZlVAW+N1KeDYwCod+F2g2RbjLUKYHEhZEvWFWb6B
Rieb2IZydr28l/wK5vjcKV1UC7A1S4GIfw3cmryKvTogDkbABsJtKZfmGcax2XlK
sfHFr2VIQbXnRM5CsuHThSCMoyC7+4iGaZSGV13rXcflvonrKSYnEQlnO5u6RnuY
NGjGE40T91aN+TTFqNbhB1EWy6+jd9ZgJnVQXM+JI/hxX6vnCBm+V46K7LIrsuIc
jNEa4gHLm7k8G+xvO29p0xeX2o3bmAlQxy6Bzp3tBjy6L+P8veTd1WpuKtR9l8/B
bmlxeKB35rgHQtnWzVbpam00H54+JqKXwIgJKGD5cQ16rpT1Bdces0ARC/KoST/5
LFFQo8KK1WvYFucg8ph1VQgTqzazxLXrcI+Gc2DuKb0R8+BNBMDV6oEFagUkZJFv
ojTRxQibvdXZ9TeUe0EoxqN6VDMJIbxSrq2RzHGGppk8jBVATwfT1MQA4hjnbKFq
2d3UtapLGBSDOqmywotkvuBB9dp1YE8EEAsn1exvRhCzRzygPwzTRvMZTTC+Joue
QCb2DPz3NIl5+baKvsDKeN0aU/j3TaWyfQIIWpxW2Q69/0fQgHRF9HaiKU+Y4TxW
7/D02pnx3lDHYAZrsLmmB2yZ0nFK0io8CSQ2MsuQsnitqMO8lwg97XnT9lscEL7/
HfKzf/S+OuG6KwPr3LTpOzGSO0nirO0NLk6dSFwI15DwV4a25wDq7CmcHNvEqXfq
xq4aWnIIXXvRuhmemzoSzxWibKRThhKWyRkNHhpMc2aYfm6HJ/nJv6HakkgWIruu
4BD4er27pioqwVgynDU/qKdIqvF2WwXGufqtZt8tHlk/ZwRMiMUcJco8cWbXNMRt
puDd4c7DTGy1HFfcmctl7n6ep5OaSZpBSdPLFlUmfo/WW6RfuuMuDHD4siVfQiLe
rvaWD5lxVQFnkOhgH5ytoxC0DLD64gZX3oF7fc/LDEocRh7oFCrAGKLqXxtxcZ9Y
cPOEBXx88cprN9OWonEi6T7gMLlz21Uq4ZNAcT5oan+tTQty3sAxn+AHILRdtFK5
oZofBzLzLrje6NMPWMbU7rjAF9nT1YQKR9HuSvVTZpvfi6Zn1ambYTMxnYSWnlXf
iP//wKwCAegSJJfhrHhRnwvVtazXGFKEx+iSOkUOJv9P9RYtTQU5+3XV2HcABJAC
Jnxat3aj0LgQms4JNjTMui+lYly752ZAiNcRYjH5t/nQLaHYaBzWuIu0e8GT7v4n
Ev0Sliwj48WZbcLbRgMZmVqoNzks7QOB2oixSTVvuIylTTbi4iHT7QEvE7+/AQST
VfTUNah8bnTzMDAmMPl6X4e0h7oEErRmThoPDGAlsQ1NwSzfN38YlNUC1gO3f/48
2hmLNAi3bwnF8u9117JnDL2iNSW9gd9zjPimDQHxgW9KPOUFMBZSdilJQUvocmiB
jf/6UqjAHCsQ0sdahANt1pqlFgkcG2FMwu1WKKvoQe84v5qAFkyHEj2ZHGsyLbWq
1IpJoOUZ9w3SLS8zpMvaYwrx6O4QWJtcBWPyIrLplt9syCj5XqGnlwFJJUZgHPV2
CtkjZ12NR5a0j+GmQI03tQCBXJDyL9ZLPR4OBhNwBEFfrTXU7q5Wr8lfuFzdR4M9
kIlSPlcXNT8hCYMUSLNpbbe3wWoZwyzeAhGABdCWsORf+K5kGOfPXFyICraRkVEB
ZYJnFeWG4pvdjOzu50Xwo53VYCHX7rCZbP6CPN2nxICzsjs9BvcnubESbWMHvTGD
FhqThXZqvOiYpm04MWiGXX/41tZEEsbODcaIC9hFKSrkhKDO/qXQEvIZ4kfFc5xW
cCnXTrkd6TIGAuBMYy3fvqeM/9+q7RMin43vrCQnH5dbXJF68XwCgk+vwjZTJLNH
hNolYcLKs2wEvtPlyQv5lK3z1L9kWlHHx5QOWB8Y/L6JHCeK31utGHLEO5Og43qo
262ZS3sdJ/M8d+/Cn6QaAi9Rq4Re80ncfW6NAWaO+7uRs4sX2rexnHoVYlaELaHt
5zlq2bgj7JYv+4D1nS15I1YSNHNSETTC5GrKjoCbhXuwkPG92nTa1/0iBLGlyb/Y
ReWOFxBPWeDwfc/+hMM1IN3jRSNaS81z7ypNMuYzgaavUwI978+Z0rEiAmKGqoAk
slQTx/CmSu18n9GR/4uAWiDezRe8qHFy8P5dC07I+IoDj+I+ylckrNL/y43qqWt5
TgMj1rXqXPRqXMZXpw1jnVYK/cVIiakNjubJTNVVJLHKfQCo81R6JBXzhPXJfk4+
ntVU38kf6tNyx5FRqN6HnQ8vhdiDk29O/zF1oJqW07SxTitQX5xwy+4RSwO1bbe2
ys8eDRk/KoOva8QzoXWBAVJqNjiYsQdNuhXJgDbvDKC0aYPvy2NgBkADQLn2apLj
b3PBetjQmFTY0+/XMsTF235hc5N1y1o5erqcz3oJ/fPm+uPqKb+Fcl3baU89NBRG
sGUzBqk08AWCtTer436F2KSti4GTCJsdscD4duPUsdwkI6JDGsSH9F4HnJKNLrjO
OjRbPWEGImVA4EZImExYFFO3bGwSAd3RGW54VsGaPyijZXhNOAH1XJVoIxWNsdCA
agPM1cBQlhzZiCDheaFpCxSP5ri9hFXVtLqZKpVNYI/LikBeLMLTGKuHbOjEirav
vZgq8I+MzU029LZ+vdv/N8SJlcaX5N1ot+WNKAKcjM9TEoz9UFdW5u2O3vrqaMNl
E+kTsFNRMeJD/KcOQm3EfTDpRiRLPQLVeATPWKWsCeXi2uEIr5wqkMO+oWRaJEv0
NDc+RqUqYhghEt/GduqjpfbWRp5wGU1ca4c3n4UjPfJxY14rcSdfeYejQGIUn6Eh
WisShh+vmMhF1pEkN9u9AazSSDSg0+dNQVXaiha3ibc+PyjKlThcB+9GzyfajtR3
TepiY9M8FadbUxU0bJReohHWpzttfodjUVqu7NXtf6hlrkZWZcbd5MlAdJg4UvHF
RML7BBxVOczDehnruf6iI9RDhTfFHYdrtEWdw90/ozMtRdpMgSix7HTe76+dTjAY
/ilz/d5OhAQ13blPOaNkk/UlosT9/f9vwNv4Spu7jMHlMXweIq+jydWUWCg3uvHC
e1WkJ1B/wcEvYQfgdDRY/FK32hhG8uO44lEH8n4Olc2sSfuxgF/aSsXpOr7UhhCl
H1WaGxJd94cTXvAsfflBnfVxExHrYhhCjUqdKBY+MGhsA8SWf2nljDK6sq496zco
e11nEWx3s0JNHGrSdjRpHRLQ/cV6qo/J6TaOYAdQcrqMoHSyPjUL7HsZl/TUlOPn
yi0+J+goAS8XNCImPsR7wv/UNLcT/LiwSBLMUjPWbhFnBOifrdVlDwDWsBOPYTPd
0uh7vcXPMMW3C8CEBDtlmpTu9Tk6l6MOYWKXZi1GScotDE2nLXWw2BRDKVNtWExL
5iACCSkiaJTn2ICdRDP9NQFS/I1XTclE/UNprfMJvqOep0xMxoCnu+fXqk5RmfKH
ZO+CGs6nBpQV9JHjHh2f44f0+9lSzlfcHRIeIe0CkiLj1ZEe8nnPi41Pr+IO/i7j
bqkPbqgrbfkxNmZavaEY9Xz17/l2VfyJONWX0NFSIIdACJkZzcRl7QqP/kENs6dM
bNlGbdCoUHwLeZe/PSefaB0H21M8s//cHOQmsRxQ1/JVsL6aWZO4+8q7oxBWf2aQ
2gCixxd1S+bzSl4m5Q0M5wnMsVco1OuDns7ywZhJv9X3PJPYj4n5rBVtVcqvb6W0
VrnB99mVYboGg0djG7mKqaQfMZS3EL1zfxwDAi1/hz2GdECJ7VRkfOdFbexRXh9T
5vastkB1ahelrIjCJ+09qp7Ab68sjkPm1rxA8JDEeJwiQ4C7na014ohVgMOFwt6d
LXQYSohEm7uH9mnFA3PfsdKN8i77UiOaf//PoxtMlGit+KkCoGygnU2PnQvr7Y1H
i+4zPXKQVpfxb+F7wgg9+Bb+IrsXydv+c8jUk93oYWFSVSE45vcwj736Qhz1XgT1
uuwS0+q1RmTES8gma1fPvKHydnjMuqZruRjk0gIIeX5khL+apFm7C4xEB2hZBITW
Fb5UCRO5m5VhzNXZhntcPQoWNnqI5DvYucSnJSPo4CXxYKzdnH9jWB+pBAMoHPC6
67vgPd/Ckd7Rp1ontghKUnN03TkP52G7fxV6o4XbBQnHOo3E2csqhOksEASroICI
GBQaFqmo+QRMteIiSe0mTgpeWdOJ3UL+JgUnqWK+eBp2150rxToBcPoMmpEDmhnc
CMTqVRs64OHdEHjikj4I11LpnvW1CSi1hFuzlZotZKrGzlqY+FJO7XtscdwIMfFN
RruCwxI857Gjk9ZVsB3iA9fJ/MclYSthVGT7LySWoeyIbG8H+azH/KQMAwrSXVEX
YwyZpZLq/P1sLktkkYlNWK3i9WRoLDSI6yGmROiQlmM7IjFlrCyhE8ZVsoJ83Ebk
8w1wXlzrsTY9Mbuw6PwuLvCgpfxRgznb+ojkdyjUdvlOigv07nalvSWtb6sMA+2v
P4VmFqjELix3Qf1uQO1LeU1OlBSgGTNnxPedKlNDP37zOqwnRuPtnP29yeX6RyxD
BILzLe6S1qBbEW+U8ivqGTQQV7hG8Y2B5YoqezH9l96DbJ4ThElONe5jPtiPnu+6
M4J6rVCUiWe5MY0skAQIaoFOQ+SeQKan53nqWqrOmYid6uHmXLzJ5B2KPqv1boM3
kqp489K607/tR4B3doXfLeXyrko6IAEmGBbiP/78O6IDF8TAbgXPDoe39Z9X3ihS
6SDNKmlYuRSPlRLdPdc48QmptzGoPQqTvDY2GVM1LLRIafhSX9ikJAdBUx1uWQjW
JtW/0wdGNV8GQiGpJlisF/O8ElmMNIzUhB4Q6hF0thDRlpqbkHgnM+lPk0K8zNjr
Hvs6U414IPHe/Z8ekCltZVlPHqXzUsGZnuGC/c5kQKgQDS0btisSwPyoi1ATlKIO
rHY9JijTtcUZitf0XziATOEjQvr1esQCom01juK2aWEaIu8TNtKgmvB5HmM8PAmo
MvRpvTIS6Kn8l/wiIo38wP0czeH2fDoYv3ATSo3zTNaqc31d0UvM9BHiBdnGONlf
zr7Z9CkTADuUZpJ2mfdWQhpCII42wpumAqTCzXP+nuRvs/71chWgHxge5oDViYnZ
CzBuy5P69N7z/4s5GJMZ9qPjNPXlxWnqLhjkAsHDJg3SBVymBLB28YMU3JNYYnez
mgxxtw/LEbg0/PhL3dL8C632ltsu2KVtIEgD2gEt8OfCEixIHACWlGW4eM+kDYV2
/WzwIwTncUO2YdLysPBOrdnffrNK/fVCDjR0EFcs0PsubjT0k9ZAINB9qqCSVB2l
qhXmRDz2xthUxohNnONgfviviLiBrWojOMjWQzeet+Y+IK/XDI6lQJMh5DILVex+
FbeR6sra175BIvhPRLnf3Nkiro3zucsDe2byV/WQz0JDG3mi20Jc99Hx7WqxJIKT
vE5qgJaMRSpOaFslCWVJ5CFY/W7I5v1XCF75OG7uf1qpXW//RqClKyMz1UR7qhLC
qR7NKCS/B3m+ASc24YhxP6lF2OOmliTjFDb8+Hkfkw0mvRA/F/c113Czw3A/AbDQ
N88TBFTWbTRtBT9zCl5tHdachC1pSNTa3y749X3mYl7oW5iatkn9ZlFARTcczihx
3W2UdqtiyngCFOXSl5JOvUllDR93e67pCAHFqr7Al94mA++9+Qz99tGm2wxncdct
lyvUpHgflBeUjby/x7g6fH7mgSloEzXlSpA6B5AuV290RlBdYn/Mc7GKNy8QP0Iy
z6cTR+bjhkNdpMiGw5t55TUpVBCEAlpvEjNlhbmyekRqGWyWrpUk9hmgvD33Kl8M
9fjGGeHOz6sQi5oP/HVt2OKrpZdbe8ENKSgC4vnDQnLyiBYHE8w0Z+GHfj1P+Qlp
hevleU4y3A2D8utKOUv1vIZgHTRPdgMqYlVE68lCaIsB2cEGcd1yZ2JSNZ65PVkR
aoAXnd/ydWk5fJrIPBMmdqYFTWHmJDHPTDRoNEGh1NqHl/4Y4I8NvhLdgy24ngY1
9ZkTqq5gH3vtClQYDkrDfXvXrSsJSqf59y+c8QTeTYhWEMCegVMNqVf0NQEH5QGA
udV80+jnUeiNj/Wzwd4E7FmwaukvyiFvywKnHJWkX8ZRcfVmLOYb+DcXPwXFxVlV
KXwAFVxF6s0Tke+OPKdcitrkDfnmMAIHvehp9u9sxtun5jZiGOr6WpzbIpxiiA42
21zrkPbUeoNSBoL54Fud/ZaLFbOy71ojpY5SbkpljRAn3Bh1hcSphemL/KhiVo9K
u9+uuhohP+LD8UptphwV8uFMFiNOIDVyIiHH9t9BlJ2aSmEi25ltXl+8Ojn7SkGE
KHMM50XuO6N2xpwW39Aa6zPNNoNTdCevdLcf2xAvdg4AX2DflJvRQW3xNAg9PSVQ
ptT+9WC7ckUZ8D+58YN4+loMvw4Sn3Nj1eMNOz/f9A0azV0MBHISnLUuHBaRqJns
rOKH2EiLyqlSb8TGJ5SApaAq2SKpwJA+ANV7n5s1R/i7H7pkAcBZKlFbix4mybCp
XecDpgiJ+5UJDaMjx6WG7HSg4zeOdbAVzkddd594EW/1ZfcJ4QiI6xLRkJnp9Iu0
fqZnO0L0XAubTB0NbVI/1WU3llrrk1sA1hU9RI3uLXKtnbMGtnuRWoIMWA60+u+i
1RebGYA1KxCmCEtyFqj1tLGqRK9d1QhbF/7wHHQQhaZF9QoD1emQTXQNCSq3z1Zb
6iK7lF55LHSAtMchYuw5QJP1zg2yedWEGeYRFLS/o/5yPCTVcc3hRsQ7cDDlFlc7
T0jnkQnd6+C/VCtDmFwwIXi4AmgA3htQIPXOLpwHhUMPagW4kEAvQvwUE5lJ2HAM
4tiLxACMZuZooWJQawEQmo0HKPG6wELuwLqk2ih+PzImoKbcbKsbafao7dFi1MRu
SFYT5fnMlVd4QBSMYVE7kYCEwH5wBuQwNfZz4DD2X7HKtDTPI4xoNixR9o7OdkAg
ADjy4g/4vKQBOV0u43wyUUzgpOfB00vXyGUQUmbW1KAA3SxrpKw2DLAymJvD1tJH
wvbltoCR8MZMGNDb0JG0iAbtsKrbV5tRwyhURQQ00oI3mbkBfPgkyLoGyba86ErA
itfJZZxatW/oLYwPKQKwXxZyrQY/zEcIGAu6iSSqjutTw6o3pSvAM2Rvk8t2jZY7
RDR/iQ4IjxMhEUzDxyzs9Ktb/5zEPaGyY1ZZqOW3qIpHDdTw4w/ukATWTR6MMnO/
bUfYsVgDVuMWcxor8OkuoYQVLFAnWd3XBsfhNIWAMX/3mwI6DPQRMeVwjfwsHx1g
hKddPPAYh0GUJFoYQEPUdjFoJDBOBF3fogn74eIUT2YbqVLHirDKj/PGVeA5kYGV
Ls5TadcpRaMTR65cyJyWm5LuRSFQpi4wvHnDXnbs/Ri/dFEumvZa7BqK15yM8j6k
8zy+jZywjXpf3WDh3YXOVHgnwuOO88TTvV1lFsIx8a9nTenAKROREQsw4cR6TBHb
cP1eBY/fY/rkZiuZASOrisj0Wlm+BDCar2J+6RgIrqZYvGlip2B2cVoQBH03uUO2
VIWb5a23krDkUkDAE+sldPbU9u00grcwQjs5gxAz2xWPoiTauJ2J2aevc7cafV4h
9e8dBtjyT77r8VIWnESL2LH9i3rkvQ7ipNm5Y1uwKWZT/K2ZrDlG3NXxKpcMiBJE
A5uvy7g7iQJmyATy7WK1r/Br57xe4STjsX2L4lvbk7o/LEhVgId8I8JbLg4Uottz
W+VnyjXdeMP8ZtTWWp2DDMq12FiojHM2x+0O9w+xe58K4CV2rv0x6WqRWfkCxz1L
Ti82sJQOs1mNUHd5i8r/ws0zEjZDR9KoCfsSEaKYENe1DAWnTV3OV06gAMlMyL+o
UsFZRM+Q5zGLQ1TC3YhNrW/iFRAjYnDTQzwuo+G1uA8uK9rOIkly3Fl0fY06RFth
jAgFingBEwsQWl0Y4Ym2zLvCGlnUB3f1sw/baNLkEnG/s2Rxpr7U5h/P6U+ZIaMh
FecG3fJA98jc1orM44C1yOSmY4I3L5ooeHkYwYsyOuB68gUsg1jrThy/oPA0Bpci
UWDdohD80+0QJhg7bW1qYYVGol+Vk+fYwYo8u1EglE09Y5SJzvIiIu7ZkYREML6O
y4Nl3Rr2gNOpnziXbwk+edjhytw7MAi2BGzEVQ9icUu9WDCqW7iZC2MFJZ2Hj26V
lIF7sOCqFf9QpgHtZ4w5KUIKyDrB7Qi77JdFVLAGovdImdY++6NZp/SgX5Tr1j3J
9lIM+vDn3cJTIrdWlktDt+SpRta3yBoaLDuhyNjpP8j8+p5DGdTHAaikgiVuKFwy
zu4MSGPNw4/PCv80KKzbQRdmuR5aKDlX6YQSpDSAMqnSPwA0/atPHGl30e3Qjl35
tUXiFdMkbQOCXy55QQWOEVgOsi53TVBErrs6KV2BxN8B6qUAFUIJouogygiwQ3Dz
QbjNEWGT09p3oiQwzB4bVJPNdA4dLpFRsoiDukboHnF0UjWLAAwfCjJaWIGxyz/2
GoeZxLjI1/622xQX7GY4ieIhclBJ7dFR7+R7IgP0OxoR3MUPEJWCzKO+VTwq3C6I
xjmPixF+vj5oyFrRm3kyJDNPkQ9nJwJIjJB28zOdj3fBge1pYc+wJZMbwUYlQ58Y
73IA1b1QfBRfVPXO46T68VN0RQt0HGsR9H7wmAGYX90EMDQ1dnZDIewFu21tsjSZ
vjUJdEFhHixUh6YQ2FzUtxBSONtdXKJZmTjFnlO7tgfLZTHJBphVPQkw9FuSvpyo
P2/SyFszod/8AOsX/h4NTZbAo5qhZvTxnqMP3RoliEgTiQIsAqiLgNt9BScTQj2Z
U8TC83zaSiZHlM8L/FBArsSKtUUp2wz1DxG9MttlLje+TlaqSrvMgPlOYJFfJDYa
uycJVVXtDd3mzQPv7P+sMb2n8ZVIYNsiqb0ZnwvTDOVOUtXRP9FYrlcMecHTnXvd
fSCm7osSsvsRJYnTyTCE+rUssGtl/nvWiVvalj4BZWAuHKxgzok2kVwV0MIl/uNz
a6LrzViWz8fgxxFsJXfFIFJ/pK6jQfxH/bDjwIrf/eQ4vRZx4B3AH8lGUIgMZOvD
bsMht3CWclCo1BkHwUqNQmlGitPabQyu1QzRXWAczOaeL/rqHsyyH2t1sLxYLe38
a7Jypa029+AeqPF/mM8jr01ejLJ7TP7H3SaelEv4GGZdMVsM5DHIBTo/ueL/rR1d
36QNwqreKoLwKrgnJkxzvURuXKHO9ECSDgxmDfCkSl8AEGviTs8lugGEmWXvsIQz
p6Cx7oKZ00Mq+lpvwdldICfPnOQn9FpGKPos97ap0Vh1awO7s3diP2V9U7q3gWcM
ZxG6qA6baxv4wKpJwMszLSfGIRzPxBOZXP7xGs6qHsBdt2CxLReuQv0DyptGChHm
OJMO8UbQlfUex5+aaEQFXe7O3M2XXgvnhaN0z+b6ATSXBJTjxnN9YgFfUbQVb8FO
WmcDgo0xMTIc62/8awKjtoeFFrUytCuyYOr+qFXY7wW5MPo+zbGvT6c0Y3BTfl8P
seFYL7KCggfcfzVJnMBnX7EXSVatfoFKygtfXlTdFJ8sk/ylPitxPOr5s5oTFCx9
UUIltWxO9RiKkOLAksZrHAy70A1cKJzNj7GUXC8Ieg3Z5QlSppxlqNVobpNVpxAa
zmmgrBOSN854RtP7XrOqAk1H5xBE2zPKUQnbtbdiIpUAE9Q14MhEOZtR5MbwgDo9
o5/KWP8A+h1dr3FyCRoqz6oYlB4yqe43qhcTQPSIDmFOnn6gnusO/T4MSUvGVFWR
Wh6L6s1aB34zxVy4gIuzEOIB9cIJEQ6/o8Ngolgb0FHJ0alFwVbKKMN2PJO+amLF
c6kkAPXWgZU2xfZi9q2QY/b/NFc1zBsMkbfxekaO6ddZoqmO0ZIlHxU9Jj94HIQl
J7y5Imq5iXTlv95x5REzn2HN1gEjDrB2Mf3UXMtgxmkrz+0MIRI/jfNqq69S1rsf
Mpm1bfRNoMkd7lIXngVsrEACGXFGPUsiWX5gy8iY9E5YTNoH5+KgXNTR0+XJKsfU
hfur4DOiRN50GVENGjSR2bTYnmpImI9Xwegsoaovj8LHnyldxorblUhQmGid3Tqr
U8qxBJTGlAFgO6r/yVY0EL0u1LvkCgthfb3d8A3v+RVicr98XcNufAD7mYMmmZIp
IA9Kp+MGdHqcZm8QqfPmGMwCrQcw0FoMnHRh74AzmY34kmWFV5lj5dQhYuyDf/6h
gMbh1tIV8fbQxVs2VN3R6oAcGuANdYMR/7iNfc9wReJMejSCiuTOK7d2k7QfRvJE
QISC42nCrWI4Pb/eEC6uWIswdVCdx4puQYutIQYtkrwyiJFxbbuK1DXx04CXEWWY
GsmDa+Y/wFgDohM3NNZnTlR7CQ51eOYQvoN2tZVh/rOwvzicDYkd6jjR6sghr6Oc
nuNWMKU0ompZTG3+qpNxNZp3/Ga8LqNTh+a2OLRvx6vg/pwkibNoU9A6O2FOqi5M
xSaaPLAiCcv3qiQOCaisLl9VC0vZstNPGqGZ1b5Aas5dIh5MF0Xls3Z8gDVbT5ib
1+VfKjLQORyyBIqapj52yGSnm1lrMwtHCGn0U6PUrKXIeEOg3G5eC+Bq51HGGV02
S7GbF3UTisKTS97+y6jWb2ZfzKAlaRqr29hQA2k6jTAb+X5Fzi91jr9n4MF8HcAU
vFJBT1Brpzk8FNKeu9gnxc7Mckz+FZQBpYUXgk/oyMOxTv3bYADf3ammgh1bP4pn
oM7uXlTIgNC6VKvC9Cw+LcPgON3UyxVgED+hhuHO58t00nYwXJgmDL3dZh9RVSLB
vpUNnJ21V0CZc7fjhmjFnDBA5NqzEuuWYNrQ9ISvmyFTBw4JFg56aZezl3sv1qXL
M/abRVahn2z1BW2cM7Z12aAfvDmeDJuOp4zC51EYUI5uSNmWSGURtSCPxzpZqbSu
hCHYANLpI1NxW4QTTDJVDO91THTR7zOxZrygtE8exMxilzQ9e96WNDb9hjIgHjSt
rWikFGdsiT5+/ADCClZ33IYjdgE0+8Ewr4xlezNuoboLG9sXpwvz93gptizEfXgt
bGxwoaLl+yauo+3yLJ+CIvb/7nZfOHBxM+xbKfUiHzXIS4NQND2hDNsW4saEKH/a
4iM7/Ouf+0f0QA3R02UAqjGBN8tBF4kfi07i4iEZ475E648qejbQAFgK6k7ga4KB
w19PMgvnAHy1B+vZxz4FqQCXXzWbGVu6TGf9FzvPKf9hv8hC+iZPBBk/gVU0YSS/
poBOt264JdhEXudNqmE/66hKxjw0uExLMOXJuTryD/HLTBz2sIfq382tRlwB19vN
0iR667lGw8KMjV/czyictVKawSC7c4AXGd4BhPAoEnpd6Rb+2Xsq9vYwf3puYH06
rZrdGzzbZ57utRnazK3SPNd12/CIvGkTUetBNI6AnqfHM05+ppcriugKo/+1o6RP
EOhQj3BmAexgnOJ/IeGcYB+Kr2fNMmRoCdueYpJ6sGSKMr9PMCMTFLsNer9OLSHD
gm7hZ73ugpHudxe6sXMllVnqhe1XQIVf+5pxA6wZtFGBAazc2xLWmGypLNvu9Jgp
hHWErnU2JY/xWIExl2+nPiaf+NYEkyvTL2uOC+b9uF410j3/UtomakqigedxB/gQ
RurVodBexJ9s4Ko1X5c7ZbvFXccSesCcDhA4Pi6ze2PFYd6luFH69BZCSaGOP9qu
SkV++NbKnyqTqEQd6N6/huZ5M0z0dofG1VFo+BY8hgsNUpJ50Bg83py8psvzJURW
ZU+mq80LWbf4mK3OHBjz6HwpJ7q32Lpl7oMBIjxJ9NdTfmrPY52UIfOm0bhjzG6W
zy0lSz1xuRHziyXPmoe4EKHqkzUgpqJQ855KPanEr45dAEAyOGOJPUTnNj5xv8Vk
oZaBL5ExKhdmNJ2GeTcMAM2LQydyEX8AtGxap4hp5pNzAqNfaYeWifRklFPsLX+X
8wmocW2pjRK0eYyu/ZSfH4FgrkBsJefZZt3RisL8TBRSaqf4Lnq5igfUlE3fXybZ
tfexNV/lXxknwkIly9FV4RtYwubgizuWp850f8uZRxmDVfLI0AKP9PHmy7zzfNYG
vZT0Vhvzgj6604so8IHCI1bxBYcxs4/SFs7m6NTH95xjvcrxLGO77uUvN6g0CDgb
vLusbVczVz6rCzShH1rB/t5XO6FfL8Qj+/DKQGK4Fuba2VAP1nYKIjiN118qqnpI
KcrnvXkU/wknJNF8+Wzufo6M7YLYmgVxuB1AAXMeV/Xq0DEW5O39n2PILf3g6w/Q
U6OiYgbIFTIx5HJZ4BX82OUpTl08Ckd7Sb6DPu1U3AL35MPH6sv3n0aQDJS7oUBa
U4garf2KN3omRl38S2CzknVVTr2qCREf9boD6Fmn1+ncAMdVQfD0kzxemcbbQD2E
hUpy8i58UgELgwa3QAqH0dyIdMs0C2DOOB3zr1vw7wAB2chMwOSNxvL2Y1MITjBM
7C+W9XzLgAjLCdXVbiAE5OUApC+lQ0XeDRcc6JY6/MhBIunj4HtRQrA4C8ixK50r
30o6GDfHSOHRWMCcrEMtEkgJg6jPbOjUikT9TSRlX8+OeTCKb1/rY0GVitT+5029
7X02YVkUiSGUnlQwKYQZXWoTzf+qQxr8dvtFhpYE1/Lmqm+GjP7YJLlbHGtSab8K
kUMEs8tkmkOZrez1jlzceSa+SoD+tR8qgzkcyOOhpuclK0OSNDn2mhvvTlULNBzA
9LEFR8rYU5XaX1L7gCrNIADJIOjEDPHbnyoO0PPFcYq3AadJYjv9MOjJB+L1thdi
Xwo93MNSYCd4Va+tFhsRw34F50C5g5sF1k+MKAGMJrAGPxE/q1jL/qEsMqmwm9nq
8JrZdF6KeAuWbFsBKGm2hQ1TjVLq95kFqJsBMTUsTzW34X4ZmFnG+2HXz8i4oG8y
f94QTFgib6/1rIGRimhh6hOAunbwEF1ArZ3QiW+uxbdwmsBVx7v618eedR472tg3
mrfbKzCVd+owfHZ0S0YDeL9fwEj/JN95NM0ARNIEr39Cv4bLpaVe/lSpKjs+8WVH
c5uL86VatFclJ6uNP1fXj3qROBCyyoD4sVTy3Ux2BIV4Tod56aXk86FhWa7gwNhq
0MMXdTeFE4SAQtwZxYnLAkV0U+fYv6gxVmsGWYt77JJKBdAhVJLIhU9WsFiuG9mw
ACMm7X0iuqPCAycIPo2ORu+3aJ2pzESjsSv8ALsjG9rMeE96Ib+e8QgJKUN+CVfJ
O+ODQjV3lC3YqEILDV+fKYp2NYapviI2JifJ/HqXTK+Oess40gZEwvbqPgI5LENE
oveTpAOtgTiWH0ZglqUd6z4i7myevRITOHKGKtrqBKcJidhvXDfnKz38EQOWljOX
nynhGL86cwjlKkIjtGIm+VEcPR+SoxgHNNRDiJeMNqm+PJ13LrwALjnGuo2Q/SV2
NkVhLUc7N4TF49Dxs/GbYTD7cXSPh+u7kdhYbX7HVytCl/xvyxXcoxjG0H7gpd8q
6I54iZeXMrgqlhgpdRZViHgg5KsBl857e3VdjBw2RD5wGznoZan5kViVZGLkqyg/
3u6xw8C9LUdlgEpRGy0tGaM4rdCk+VnPiHFh7GBSSOqy2KGf1ud+RL2Y4bUz3q3n
sQd8ySYcOaSQVTxhRmgFPooqEBw4kfbY3LLF98fcuERgF5FsD9M1PrKJbGTkWQva
5OAq0MCHYqcY+OO/Tb8ZD46fb5qYWHeGsMAXykwEaigqYQJScSnyhpVEQ/9mDOI8
9QNObaB1Bb6u88qaUU942rUzyj/9fp6pnw6+dGzIVZt81y6cXzTZGPt34A3vRHG9
+jrGgeFYR/DgTUmOtsgoBJo6rLV4eRNwyhtWcKfLtNSMp+aHtmhEXBsIL4E4e3E1
UQvAC4Mn8mCQdOIJBiY3cTuy5dE/uMfiAv6SsQf3SPWfr8CTdUtBzWU71Kwbx05b
oVh0SbqMK4nE2f4fN1MtKFEUrB0ckmBDGehADNZTDg9Pv0u229xU+AZ2hSnH+a5N
PHkclDpQpxElNQpTyfpAXDvlSuaDW4LzOUiAWjruUdwqksaug0TUOOsCJ6zGKqoj
Cgs4cdjeyHfePeUM4w+Mc98ytzDnKhXs4UjAxDOhgICpin5VhjlsTtgVXaNcXuj8
8wyp23w7Z1kNuT95mzqRrJZ9iM/Eooq26Rae8OnjQekXM4Ucsj49FfvpnLdFF/HK
20R+ESW/9YMGihGvheb097fJWCWHiCQiufQOwIyb0GmZay8SH0VojiSom0pkRu3D
OHK/pUgsKO77zN+RTTB7qa2/ynMgJvcgWbQD07ugL8+GP8wzCIcsNLJJ1MAN5u+H
kMcCmwr0w4553fkjTtcRAB96U8pTWJy7AgTEeSKeNSsy6PfptehJePBKQvZF3dnb
sQ4g8wKjmo7Tw5xw/y0nxO4tds1Inmy/TcWmcLzMFShdNQyyPVgEP0eF4NbmxXZS
qPwLwy1wCoCVO+KrQXfP94qb3ykp7aShIHWhz3GWT8lFcdFwL1nlV305mZxqBc5K
A8V5uGbu9qyOMBzFmXIVuhHBJk9swe4asCwZx1JnwRlTzdKBlHCeZylu9mGGlwMY
77gxJk8zSTtAKLWaVkWEp7xjEq/gghtRRZxzI65/Gtyfu23M12e6sbJLEE86zV32
g0EXysvMCseo+7Dy1GXbX9yn26ciC6dk+B7MyO6AWRqo+1lP6/FXWF62rdBndp6Q
3fK4wfU1Y9yaVY08xSRY+PX6FZd3MTtbmm4YmEAe8SEDJ0qWYPD60DC54D2GXZaU
U+B77yx3DPPCqTlPV1BdOU3ejhBWX3VCCKWt4Bf2jc8hrbSeeIokzzUMe/CQJ7hP
hLQ1seCKdff35WuU9lt0ZBCbkSnbPCU38sT1R99UTfoUQRDg2I5rhcjOKEfgprgU
cJPQpelK8zSNRN/duISV2do8bBOWq191gubUhbPOvfJ4nuTdCMARWX+oW3dKwKhf
OJjf8APCh1A52wQKsy25llOH6EOHtSB3wcG102gsOnHJuSEVwKQ/LEgCJBYimr2i
J6pWElf3vkoEPLVwCoTNUBZRpd8Y2Mh1DijKGGmJQdZ3hLXoClpmw6tOCP0mWyGK
pPw4g0WSy746VD+2kyzHHbmtI0X1ZBBjrw5wKYJvghnjI55Bg4aZBbH82MjIDs9s
qm4cMkQVsE0J3uSULPLKD/3+aMjU6ssOEwR+FOwQYBgSZFKGzjkGZhDNYK/9b/xw
1vM02oc+cTS5CPJJpiODgEetXGdXcNGJhNGU6HgINeZrahvJZ9RJfYfDHgFxfpla
yzKANWtVSzuKJU+SkNSKhOo3PG7kzAIGj1ER9pkz8ZnOuAebJwQ8Al8dk4zqg99h
3q3L8/jjKTVqFoPKu3KPQ8JbDq6E9ZVlu7GoGg1DgkLkU43gSrPw/6HB0ElTtrFU
7hwkC+FMOinfLFv/MUOE/aE5AJg8SjbMB595dLfYmwu64GSSz2vm6bQjzNuVpHtq
kS4ZszAwxqlDaLp8pmCcgZSqA5RkQBcBVQmyuL/XuwakFHMrPzHS7TQEP+K12+/h
JnCk5/TFHTM47IKxNjcZs5F8DyiuuyUN8O3SX69DnEc55XIqxWj/QLjxnX+7i9Dj
3Rm8+eWv0HoJ17ujmLKLGy0qpglY8r0PolPB62mU4lOK76ro1f6enr/NG//ZuVZ2
tDwQ07xAFoerPBWDUoZA8vI47f+OtjRjpk+lRSqCRWZb4+OsbAOqbMTJjr6gHHXv
Z0SwW5i9xnqFdIyVQPFEjOWQWnzF7Feg63X6uZ7gky6UKTKdxXjNLzp/7QueQ7jh
xshcPttjjN4U/qkHTWU/1Owv1fUh+T4i5CWbnCh38lpo9yAD5QEUGFBTnoaUQ6HM
mq5LpcvLYf4slqD2bYlQZQDlSjOZFrpGX9TLHdPvbQ5jvMEf7cxRd8ii1x+GzCL0
GsUXzLHI1ecbg0/xgeHJNN1LW8R2vsmtsbqsAOGLXuzqvSS9iaJMRAoTuoxKCLR+
C3+pnyYfJ152LbkPUZN/1gjrSsxBnNtBVIrbJfCTBUSmNCaDdIkYfrgXys/+rT5r
QKHDXSkOyV11vQ1QHx1GicYKldEldQjnT3RB4v2rQ3dGPcISHBTIb3kxhc+oc/hU
iYXCzTYUQE4OE6GoPHHroYDih1YtzAU7pLSS3cv60bNc7CYVr0NQskpYV8Fb6XfD
qYROJyGUzJXQbfvCEsSvwxGc523EewC4LZT/gllXq7kjXSvuYaT/GnoE4EsrBJFq
jy9bZ/2+Qxt4SLv+n+oKpn6hp0WwNCScxiNH13PtDdpnneCH1qyRIwLhIp7lBH/Y
HxNhOsFteByCedunRcuMCK5F+ESdRMW9LFV9hRISaDpqBzqZQGqk5eov2UQacXVH
kRzSFbdL2RrRyJs5yZL/hEk/gGuNWhDVBl47yWvUdtkayHoVKj/D4/1GoEIOrbVE
SDx39DfE9obu0v9oGfwQBZNco4/Au2u4yqDK8+ofCHaNKFWTLe9eRnGFdtIMCcQo
hemjaIIwZFju+CVXES9sSLNR4Z6AiTaQKyH2C5qk0pigdBgH3umRDb7PSwaO+d44
dnJnKoZuMlr6Uv+D/L1FTAgNfybO/LRz+qxezYi3Pg/hvXIwi/LWwuef1UizB0K/
JtVFI3Oxx8pPUNDKQhVBIUXeILMNPb/xvez2Ymy2SE64XkCX8l8L8eUSKOD7OR5m
q/KkxZbjjTog60BVxhmwDBsSL5keZtSfR/RpUiRDF3hzBfRAHxxTOY6/BPZTjsFS
2owodYcMS1tSX1/bMhd+KFjCUy4zMF+yRfBPNczcz7w9qV06YBmR6uIhXzKybrUk
qrSwdtMGgrCYGsHdv3LeQhXqi9JFKlG0L3Z//2PbirH2dl/GvO/3K6ZqwdRUs/cE
i80Lid3rfILu2KzQvV2lyrKIZ8FtC3x8yRh/8SRmyq+UM1MeZvtsv4II+wTH5jX1
8+41cKOhb76RzxKn3z/7aB2xMvdONYk1RQHjqciSNmgNr9wTm2f3DQEmYORkf6W5
3/tzVuHpKhk9QIiD+riLhX4HC1oWOTZQYxQFntrtpPQtCnWe2PiGNXl4BnEfYyFR
GWoBiA0K6b+Y52PWBuZwHcxayGjhdckVSLFcyrgWO8A10EVy87cxY8VYO7AWwFbx
C2pXbsgr+P81o1wgKfQv2XulJh0/AalOj2dhaIqdFi4qvSFF0j38j5S/k8LHTXPs
Mz4NSyMYcixMagSC61cRAOpfawL7dZ0pfoGrECBoVBiiJx1sxUtaAI9asokUA6fW
cU8JkRTgQa6/vdaslq6uS3xDdTVKWRpJiK/t+PRhhMdHKh3soaUsC40xRwNsaRZE
CPFT4PChEfnNP2H6zGcDgZkeNnxBeWPiwShfa4kjqB9NSOiLanrQyzmfAZ0u86Li
sTkP4TYh/M1hIB+BfSWUg9XK4oZtTAUB1Q6IznfAp9pCcJ5+p6Mg7lseuO6Z4y8T
y2zuvCsYo5lwTmvPXeX0ibypj1aVMmYUHuV1EPMon2dBbNgqpo9144ry2y4nyrrt
c1oPwIh+HXcow0BTsD+YNC2mjiFEOSSBgagdIsBu1Oiqpl8VEihDdlL54b0gYn4X
8ZTwv74eNE3p3hab76LOzq4YZD7eDvdfcfnxksR9iek0Og813s0LjSkz2IEBO7PV
YO8lBBz8UFcEx5mfKvntRpXFFFr/7U7fH4OhyYXOlS8yD1ilVxM9QlxzYFoUEGS5
3bEB+Dh3gJQwjoyg2sujUGFYVm4tfS45WRVBvkNb3rE+/mvs+fkSQfZmMOFPrxtp
KwgnXJ0xvVHD/ZP4JAEdHeinjvbhidnx5vkhkHggYOMAjmFCtsjcHoKmwdzRB6xQ
oy9N05o0H+VvU3qCh/guvfQLN9CL6kK6NnmDu34JhsahD54D+LmM2ItXO2ol2Wyx
3FKF8BDgw1XHxSRs3jNJmye62c2Mx654zvHT8jBEBBNYhK2xIcL3tStxl5C9GCLT
IIKljVn2xuT/EZOIMJ9p55AEZR3ha/poI9SSXzcLWLfEkqPL4dtyuwPwaGAIMHUI
sKQ2wj+HczwIfYiZn+9+LGvTaj4++wtqIH0ZBOSGxI4oaeCpSXZQPrTYSjSqyMce
3G37G8yHQ2pBhsMgp3VPrarrWM/HtE+S9hqbSgGJBxYp20op2qcjNo4kAk+ItBod
FAvKO0BE3eUZ8lRW08FxrGsagnn9SHapHFrXSIr6D5Quwh4KpLeJ4WVfd5DmIjqm
OHbJ+h2icclLNnm/84FBd8zfh6Hy7yLsvPaXb+UfNsuWR/kEp2s0DlF2taien3qo
VbXI8uOzfXgsh7JBUWM2z9lN9b2NCE2EqG6zhzqrOGnSBNwKiYtVX0dh5bKY9qnz
Mn7gMC2gqkTcPaTRw++NnpzMn8rk8SpODR3mu3p2XROWMRuOV6KF/sXXN4xS4uzR
xG4VcwTSQ2dshztENOA91BaN8WKJGXBT1VsIuC8qtEWM2Gnf3Ps1IF8vq1d1Yo4D
5zJ4cADk990waTYcSHVe660OExknVLBJRdOVsQehm6G59CY6pOS9qS+3zm/bIXyL
JUzR2i3YemANE1eJHcA0DF4W6hij5GYQEBBC4XTC51JGNrCFgt+ifh3XK8sb+6aL
89jcY4o6Qh5vsZ3cvKMS4xhFtyEdgl2FnTEBX1OjcRFZa38RLBtLab6FPE0NfeiI
IR4G/GzYdAbVlk+qbChWVs4o4JXLRdYMBZxC5LgueZ/ZbsghiwjYUNE8SGxGL4qV
I+8+YLPR950dgboff3hpB64OyxunB9igb7Yo/eqI3jbIA6cUJxu6BEwOx+VAhxFf
9bqKPhJOm0fADYG7o4RIVKujCtKfM78W21beIPkzMYAW6e9o/cUMdScv5rZrCEI2
kPfwrGjb0sV+TOOYTu/y9MWSvYcZofvJaoV2+isghcbTjYqEf2sLsOzwIhyhqk6z
HInfTRfm41Tkcie329v5LIzhTkfR+tIrRZZVsvlce2DFDvSUi51dg5yUMt/SNN40
S0duih2xDQbmbrPx5h46mpOq93d4hJP2CO8dEsx6dLETL+18/yU+eZJju6U2EAzU
CQ2YRrw7ketU8+ujmd27PAGX7NPOcrpOz350u2SSA1q1Q3ZCnEIWEjqEhh0SYL44
XWqBFp2+o/fuh1WyeHoTgQ4Me4eV10to+Xkuko6KEeOXY9JuMNWNKXm7ytLbrHu5
TeSYqf8HdrDfoDrPWpjEmNnUCpR5+VdzWZKr+XuNyxhguzYMvm7MwdQSa/Nun60d
OGYbNEJcx7KlHrVS3Q53S5gxLR5qf0VZSpAa/PWRayRskb1rDIG9Fdb9NJ8NYxmF
80R+p25lsjgHsnVs2QeSUfMpZ7uZgP7PUs50xRRH09xL0qdY50CbIg/MQW2pc2Wo
YB0mfgqQ7AqQObzl2wR4HO+vyII5nNwxL4YrjjgAqDjUgxrD3JCeXzn7YzDtsdTU
YdMQSbPi1LXh8m8DZgT3RLCcRco6ZityHbx399TcDcE1rxFZQ3HaS6p0Z6X9RHvT
7ww4VlwVc6lN/KHYG0XY0mnvyaBoCFJoY5n47u7hfndii8i9qxYY02P9Ub/onwFj
NL/q+hmV7t9Jkp2+a/oedqirvU6/UGs7+yl6fHMr9XxU+aDhCGfdpq0JH3nuZrC+
iwxaDpff3ehLUCEQxpIqQ+mc5LrAG7iuVHubgWiklTxzrpeOHo/d448bn7GsUEUk
fpU2C7Ds3e+yjZOtSUdeFlA/qrDyz6kqfrNmTh0tJmjOCyDWzXpqmT0oiYiVXiJb
Jj/71XExhtm4hz6h7pcYkHNEPHCksritZcIjf38pEJSWeswsQX1ic5upjG33BI3d
DRGwcHIzkL8I5S9Mkxyef3qaDKpEE9ZxZeNkaQRAl7w4MXIxiUavOM8JD3c5WRXP
5f5kXdJRcm+o2rsX7wEGqelaVdDvALYYQEw91xxzN3FCPct+ipHftlvKgwca+nEu
q4LW3QRTGqKF5WQOSooPz1KE8ypPYnqSQsnlSPS9Y5YmCBvQabWUgMQrL5qMPs1p
mCKackPgyyosAnvnGEeJS0RAnCuGggw+O/W4YFFCU7zw3j6U2XtWB+/BtEprBEgZ
i6PIofL7KjLEx+/7wD928v23SGExwSvNL4HsfkIdRlfxVz+RNcQltafZbaeJ7UiF
9aWQqQgV6g5v63T/iaglLSibZOEsyeyo64+od/BTiNX+tjHagK6b0cUINr5NMK/Z
AW48O9505P2H/rjzRjSH9l2b43kVYuP2QrVUyCx+DwpJaggs+4Yw8xCC2qdRf/Jc
GpL7URhdrSBajZMdExxAZDHyRu1NqG7mDoma8tyHxcb96a1tH22Okyf2DEr4UxR8
pMLrDoKJ1FruGYxgpDzLn8/Prd0ljgJ9zd6W9zlVDHIxNtMmwTAsvBEsYAUeWcc9
AsNbVlkmKTnvXXyD3nNdQlSfJNhof7URABUGccHMlUxPMCGre8rUsrCysulb0Ozc
eGpmQoAyuJwO0ZJyXRiJlu4i5YIsIcIhMy8UUKL6j0QtgOqHNVMYIn4geDexz9gv
qGtXmLwifw3VYBzsOXSK3+ASgWu5uopg50OPdWbWmjArajxoTcZLgyVt6S/yD4Ls
i6WFj8z1HPxqA1wTIeB64RL6PEmYEz1ah2gxNH930AXER3Jpqd0ep1GaZDy/u3Fx
CLiPJG97VFlJEFwSDidEcJH5tF+tC+h48cAjChlXOdM05HbjDqekVLpCXijEiDmi
bDNZeEOmjALTRvKrjwatW6gcasK88JxtoyFwvcSyvBpnmqgJ1mSjZalLiGDBxCEO
yYb/sIdNSjNmDeyNQbZbgr54NmnWGrbKUhFQFGPMAGmxQfKXAw1V3X9SlHoV5Vc2
6IunNbffNxoSOpZWnJfVfUoR9Ep+7VsjlLreeMpFeZBDxUfBVXuS6cv26uMLQMJs
O1vdGNAl9DJ5cwdY55DuR1/thvzC5WN5ns+RfD+b0rJ5o1BlS6DJp5m0TLYVIgAa
EZjER3mSugMV2rifxb0uUouTu1Cm/kmXPiR0teQU51RgAZMGdjAOhFwKssws3pLd
XPvGwNlxhyYbFyPmbskQCN0z/GGqMo778gAFIpSwGFyOIaZVNIeFgLCTG83lw2Vj
QSj4Uu6smwiy4Skx+4G1MhBmXcCODla2T1f0cndM8QOwXoeq/yV56NySyI5eW7f8
swfuRIllSoBBqkacjJ4uegry+ZuKoqW7ps/0auAX4eTtwK+Q1LG1FdkNE5sxAv2k
XfWSvbYgXL7KyWFf/NsNPKaUImjWmMNrubdimFLvaYj7EZ0fGy5jh6LxDxeblFvJ
RN52U89BawQKIT2pq2jVRPaptEz2DEZCEBfEcGmQ86vKsj6jjS9hll09tCCh8XOA
PgQdpHUES8E8ae8Tp8wDF+0s43hieRlOPjJ3qt9fbl0kQ7gTZRPLbqXFdLSP3VVW
HhC0AmmMcd5L+YWe1uI9zJ6zSXtLIgi2OYvNT88GWvs5G/YH4G7WFJgdTrtofUU9
7EZetUByWtFAAmxEwz+A2TTD/wy7yEmB4IrDQlsOjvOWaynXDdaIt1l0GzLGkAMP
A0asl2HAZXa0okP06m7T5YQRHXk7qdxmhMDGcuPsr55yKVDz38Gjvo77doWO4cnc
bLDR+/3nAdeeUSMT8sUcekK43iCQYUzf0ZNBAHf/AbqXoCiqdWpaCFFln6nCWPMo
9ycPMA1dZjZ/JdP4VsguDRFDLM4xcC2LiLpw6+dcxwMGPZnYCdXgVGsDjIPhf4t5
OLmncNaQoyqotft6V1kgEuT32XuA2faMrS96NUhR59Ohbo7PaD17fdWREVFkCCAE
Irqf+uiL0TLcP4noTeCHazO8QLw3jURQdsnbjcj/nhuNf3JiRcuG7ogeu+RckHVp
GDbIz+SZQsSeqjkGg01tBTzG6wby2mO+DcV28whtxO66Nqc7MCJvvA2rmPMd4MqM
QTjm/RGskrhSR/tJXE1LkqK0HW6i/BqgYOhTiP2La9KBUTy+n0jLWfLnNmkGXYBf
VwhB4lBavuoCGNEQYX1saJg9joEmmbYsihS0r9t598POXeyhnldrOttc/B1xeqVf
v+nFKZ2sAmTw76sGjFwJ+JMM9qcLs70CiFQqXX/GNJGcfpUWzY9rRFLztQGszrjs
/DSg3Fq1pbTeBkkZuuH9OxBjDQy609trVFHs6v4Eg3vcYEFllIXhF8uAogPEx5wf
z4WrqJtjAGHSTpMswmYA9H7JmFTgPNZS9AU1VtVevvolIdjNrbyUsIPUyno6e8qt
78AV7frfLoywmwec+i5pwPCdwbglrEWta+/J9wNLeTq3JE16Dve50iyu+5EV+iOz
mN7HY28dvPRc+6LIpu1GGYoyrMlEVy46GqMXi8CNYqIK2QL9hRIfJjf+iQc9I4Ap
ohwnNNbF5re8H+TjSJgJxMerogV1AiB5FKunvlDTCPg6QzvBreMktekzsKPdTNmB
pHoDw6EDl2uT02ZJ0SbUcTe60+ZNSAObZ384QBsNFw6yGi8cw4XiVCOuQIG+c45f
TKKIQHU4TRhdPlZ2hzGUMbarvKb0FF9hD4e3kvjpJk7wvItIf5DdD3Ki5kH0Ttg4
M7rFKNcZCssB3z5hljyT5yB4ylhwvYGoPpGUWUTwyebsT/A6zWLov9Qh3eQBMfvK
PAdFUBzsYdrYrBTZAKOYbVJe82aUIjEj17ntDJyBGmSC70szPslQ1fnvMzLAFDpm
DbK6tH9f3rlsw9a/b5kXfdbjHjSUY3zZLeFUzkxC5xA/F5dwx8zv33vdJZLnMSAh
YMyiw/yAp5MzVArttismTzghR+lm809IGznR77OfXjkWILNOf4j4hVV4CVBs9zRO
Ng9uViVVi8kuUxMtzNlWjmErUVFT2JFZR4RgNuMpVMKOoZbql53LcVk5DP+brgzQ
/5KtlBDZml2DOmLIZHEXGcTTLQHHw946oU84ca7YqgN9iDEYYPZ70haxUfMEgYkw
VcSEnrQAx7i2EkwYzjmVCi58cXn/PreZC2UNFTocI4Cy/0JxTj9H1nj02M760UAQ
IHZT1S5UF1hlhNlgkomonq7O+B3iZHETkWOjQvukj8MwIgy2ptXm1f4P0iqauLQE
Wh2HyEoi/2mBznOLscE1GLS8PQbPxBFDM72dl9dSN9lRC6vciAhSplgtKsKTccU2
N1/qEWF9subV6BuQz/EBN/cMgJdtTwhUp9xlFmRVVqyCnqGhGYQnTHKUuEjFRAD2
pU6uqdYNb/3Qr65DRsO18K3THHmFrL8xD5SOT6EHSjgsk95Bc+lRlHjFalCZ57J3
HUa9S6KNhJSRcBISg1so3V0oBMG91AiVNLkhsvAz5viC6zJ9zsY6A3973x7Cuz88
T0bPLjIL7Uy1Qw6JhFbs1HLrFKUIqKGW3t4X+4DilpOU7Tz8BmmlsPdkxhtRheUg
7s1k1lZzxu3bzLmv0adPcwO7luQv/rFnkygVuUI1NW3//RmIiqCZL0bC170xzGxc
2cA0mp4n+k27BJA+tPhilE7aMDY36TTOiSsxca8W6fMVhNm/obA9dFNHlXkDZtds
Fuur+DqwJe3N9AxDgxV0FaaiuhxjWM0Z045d2+gryxhojr+Ot9+kChWI0aec8vz0
Wjp6mVoMNQXxoDrId/8s26A8UUqMBhUHIPIetmF8LFS89fLdi6dzmcDhCQEkpoX0
U9PFN5Dfj59Ll6PtgCClQje403OA87ENlsff28y1/sql5LDSwwATqizgrZTIrVj7
xHp44ZadRQ8CvvILAt+VEXWpb5b85hsi2jZAPkNM5+pkNgI2pOiFYzuy3fivNTvo
0ncVnWLzRKFtr3SMtGI4waxv79FnmadwY96Q29VuDgLFRmfFi5WUWyb644IZU4pi
RrqmPy6e5KyIzh+RlGXbIB0DbV6tKTBlCCP+lGqpDPtWZc7k5YdGfHBJXWuualKl
rDvJwqC0+cK76eVTX9jswqT7s/myeQ/F+U0owgaUVzOUeVrS7//QKsuhl2TB+It8
KQkEdpIxqFT3cuwbns0V9d8SElJWLaFSdSawo8bSUkvNWwOUSw47TAi4IkD1hsFF
UT5ynaO7xOiC+pqpDDXt5IFFffpQLW20fSfanWdhU6DhJ0T53ZZ47kT7xdnplmf/
9qMMBrOeh1YcC8LuQRnIbz8ZbhWDBHfu41LO264qh3B164pS1eWkBaYjtqkP8TUn
v0dOH7I9Ah63p3exZKrQYZzfSVCa4vUTj0RnlNjX+jiMkKxO/+5gKu/OFwq2uDhC
n4YeYyk9QiK4p8OvuyWZqadeUM0MHTSqbECO2QjT5Nfj232ujpvY4RPyeqOUqeUF
YME9vbAE8S4JaERDrmMEbf93VQ3JAN+2CmfxuLv/06ONRCm/WVKyutQunnVSBhTm
/qx3amfEviVIZ5D6Kd1ulrRnnm25hMYAydO3+viOkynPcaJNOIYePWA/t+/X5mbM
9ZA3+DdB0V0ANIS8SVdVgoUA+HfkM01qPgJr5RtT4C3sS8Y3UHVL2ut/MHrkUP7X
vabEurgtGV/7sZzMEmNICzLCwZ0QSLkU7kRJzj+WgHUy2Ng8xU1AFfUlvk7Fl1Y2
V+QAg75+wHbdtsjq3SKiillz6adVs+zCOD2OWwi22vEgs4apCg9IG4VlQVI+KhhN
a4fUmRmD8xOONN1RVZLpA6Ih2TSoql+nkGoS7EkSLBbrAZ/MHfZDb0How/tZuiY3
XdAGSmZ7LBK/P/Mw6XETC8leU4d/OQw+Ee4mq86CxvcHBs4vXe7PCfhMaKsw7FNt
p/tP/uKsiGBYrJkjvSFts7iI8me1ngj3Xbpz3bTRL/1m0fPfj5AkstHQA5qsMWxw
aEewB1J/z2egU0RGmOlecak8BWUHAQZPtA848Eps9Nk30hheCt81SpTG8dF6VpBq
jDsbSdgm7PGm7J4AsjcVrrrzTAb3bf8oGV/Gcf2Cp1ZzlsF8d3a2Vgmy4PY85ixS
6kuG2YAxpLdR3mfLZOvXyyPsXevNSIaC3BtiYLnxthGWjQL5P15CATjqFY8UCKVh
UoDNUiIgJKSX3aZfuulF+cxMe/5Fqhmpx0g4lHcBHYk3apPCAwU2BWKRrroT/wsF
1TZmOpSgZ1F+BfhrmKhmSE8c+95N4bZXMilV45HSk7LMeNmkHNAk7CT51U5+X633
dmJ5XHUVxZm3mvBtR9CgJh9A9hRFqOsfdRmCypc6Vu+P2IVF2LC61F6ViDpmILFp
C75JOd5WZpLfEYBceZzMip4nUYffL/P+y6kpbJ6RbVlTpysZiAT9Pc4mBKK4eQFC
yNKTV0xTujuUvdWQxPrHjLoMtAJ7wwdomNURlgWCIpZljGNg92Heb2XIhcICeEG1
Do/UezkGJk9HTIWzfpuWPWlsPy6EtjHZdRFAf6Y7XLiyAhwElc/w7aYhgYSugRUZ
XwbARdQFI+j0FwmjfZWK0dakveeDhWiPobh2eev6Kb6nMTGH2Hs02OoXGZ5Cwev1
TC+9ENnvv6EDDSh2GdQRScKvmVtyQ4poZY8YPurgsvmZiO211hdUTfrJGlOXLQCq
5GtqhalLhS95cNEwMLH3wP4clWwyqvG8kwM1X7SHNqAFbGM41svjnnQE5+RQsFT9
3yIsuMhGt2hRJEhXG7dtnt/pAttgFrfC3M1Q1crKSHD5+3ioPdW1r358TeCI9tFT
n8vW2ERQFo8tmMYJqUp1bkQussP4cNBDX/xT6cYXO2RTXplD5QzXT6k9MVGt6yTh
RsjzJq8XDNgtykgPlqliFZdrce4ix6euHzovtGhp6KScuPXocmN0vjXLKdJQV6V4
cvV9ailDFApt6uhRSeqRR6PVRXYjqY6aer5KBeN6op0qA8gpA2VnrPf0UkYzqTfw
qZGTIQmiNL+/g9b3S8vkONijw0lPnEZtSCHInBg3TaUIxRGpjTSW4gNHkzEpr93t
Z37r6XtaoR+R2pHWXvj5pOhZeQYlZDEL+o9OLOrrA4i3uEbW5VgKwbYcE2vGYIqm
x/z/SeteFQ0i+iO2Hqjrboq42yVriYPELkGO4JXPkJBeOGHe3RZvM1W9BnQVroWT
BIjcEG13tdGB5uMBqmD1wL5DonopWpigBVUVvlZrGCcUVXEE3D1mYFns1vbwThFe
lM1AxhC7Ycm36INBIr8gOBLSFqWfdCYWfSzlh7O1fveOEAbDWHWw9zgpviKb0/ZM
CyaZALCfVh52UeX4DG2ucgidQK8FXXuBHBHP0BsY8yMfuJxV7F21BTVCzZoFzAJr
IjJ+xJntjyjdUvuff6NI47THllojtM5cMFmHOkLH+d8kOMHhnF3SGKyaJCP1VXyT
K/KB8VRKMwEJfJuOwbq0tEYk9iWJ4ScOnaDcZMADqHOQETVguMTY/MqhOPau9wSX
ivlsmGRId9p5NmejNHRBciQTLK3s2gN1kYZlRXe6CYgVyXGEl46nUrW5rDDyF+v0
KR69brMOfZgVKQ/2+0eKaxJtbChJpDBtWDGlubeFr0gU9dt0akNqDpqYdLeqVjF1
xhfTUhcsGB6MhzMEEK4jgywx7g/FDBE0P58Fc965D3io+Uiz0ml5ONh8ptwDMh0z
kDpM4woGLvToZ7bSQzHCXOMbfFD9o6UbXV80S5Gf/gERi+M7UPSJMvcq7UjQ3XsG
UKky/UXB9CENu9ctwY/dE83TDTrZFaVcqWHlZLxrr1/xcdhg9/XU32p0ee+gv0Cd
NLdo97mTKHXqcZ/sjDiJ6CRT6KnmaO9usHI7v3tKXvY7k6twDZBL5RbBGNZRILHl
Sut+ljjbhtABoxi1vdRZbc6yV9RjrnDDcdqFVHVReHQNHfk11iJ733ClAyN93fi7
mdPwie+dTYi6rAEh684VZNQegfh89fYf7pHptPVDCqYlSPN7BJLBhpvvDJ5FPU0W
TT1hvnTIfR67DIU6k5D9sSk0oowljsn50QoGpW+y/o1UojToS5ZbHjFiv8mzkduf
fGmB2hFJGOgabupayRyO9KjHgCuwIAQIU54aVKB6Yy34TL3enpv95iWi4k+1bJ0r
2M+Qu+2vU5QFx6kUoa02naM/Dei2rWAHls6PnPhB0yWot3EllOFDsjL0ZflgNJXQ
sKbrG9UV6Qnog0XfZMAyKV/QNXQ/tYcFBj7vHHnv9OkDg2w0SrslsGiSRWZzx73S
kbzOVh5aJzZDj+KEpc5WjoN1lNwyQ5nEu+koCcjZ4BPBT0uM5M2cbEs/dzIVK0Ff
k1XDtENSslOkBonV7ZhsZfRkiFqYkAVmrsqKV55pm5Ai0XhOYFL0Vx7PYitRTf/P
4Ij9/J+2hbIqqF3aBhWVQDMjJYhjkIF9/HOLOzjn8yfMpah315gEevxOcgpRcwFd
UF/np0niPnJf9eafbNWBQhPAadZsppTcH91Kd+UGwgO0u3+/fV6nKLtaYzezciYf
EQyxvfB/yIqrPXuSUlsatJRn3gZu7XkQG7xfMcvfP1Jxn1jzKR2CXBbocbgfoLbs
IS7GM1pL7Qsdgp/PbqEcppr3d/SjmjGPD66MNvxUvNnWlTUZibtXKKXtzvnUmDk0
Nmio2zFDx9mIwf6or1sNTVJGoRLco0yoNFMXf5rqblM3bg3qa0W7UoHj4+s9EF4Y
gPxZqAzEO97AKKPB8zXHDxYXDZHQWtQX6+eakDyA3fNodSO5w4ObpZq0pRLTEZkF
RuFPZAgAVn15T/2kCODTCBuADVH9LgTv4M2TXSwgWdoMx4e28jfVJICl7khSg4he
PTLqpFNevcMoTQWfDfSXWFqTEmOt9olfwPENbQBwwtiekESgqKiBWUR1lJqr/nxb
VWwluVWnBtHGNE4lIsjBJo4phqQ8xNIV0uzKqeBob7CxL1lkw3LBCTBMFz29Jf1K
1h+3DbEneQZSd1GiuOPdd42BdGae7cJCmvvlkW3cSkUtlDk7Dc93csVGn/7xkr+s
PYueihO263FnVQPKNAux4id0FB05J42oTXsxEVWnyC5IeT6nMgxGHWI7zhxZPfsy
kL6vBLyjF6w3ssdqbeZfItZRW7kUXSstbHINpxRaZDHghVlmB16zG4s4QmdYImk8
CckMhi+8RA2cX2B/KrNrx+IN0/uYB06zWSZio/OXEZKJ+MaEGhia2aXAgDiautVP
HI/7HUXXENnNE3PIfA2SO4NPqIyOtYXCMfgWka/v9rm6BijMvI8NOGC7o3aY0t5c
0B/2nmJHSRFNlQstfRRVks2U07WRUYLiBBjB2bQeKrcrhigO43NnveduJX3BTcmc
dtRkIZq0Bt9FPVlhoKb+VGeHaBEGFziDwStqClPxBRuj9mctbKoBBgjWPS6cuenr
aNrn/SzJ7Y+vuW/c+nPn8Xh/bva4i0M5kBZkEL4bwZkcPQlisVX6AQPQGTHNwaqK
EH2zAtHkCS/bJlni1Ikiw9c7wk66iEHJVnsGQzmGp5sePFiQlBKn0ONJCd4J/AdP
E794fZQ8Qt3zBFpJI+P+yMvf7XpvMDfatGUzfl+1df9th1f3fSMuxCla0iVMcR7D
guseYTBRKae4TkCERyj6q7zg/MVfoUBDLgEa+cSwk23NFs8tvucF2wHsj+ODWqHI
I4j1L9fbY5e5WQwz12uBCNMJpXRWm3+Nugy1Bo8w77noQ0AObZEXKIj2Ha/Xg95F
PB26mFE+WlF1KfnbL6nmOs6qWWC9FigMGI6N0cSZJEqK+0KNC90MVrtpr//TSNuQ
/CXigS0FT4sVm7S9G93pYfX5Xi+G63Qi8i/rPraFOQQ80/NVZrMSEye7UaFPCFcc
xSmN03JiYxxXQ8jY2K6lf+s+QknkY+s4aSo71Zy094g8V5n65OV9uRRgedaVaMnN
WN/1vTBxs49xElCB1vJm94G+fxpzrZKYeitFDcFD4WT6oHEAj//XGw/A8AyJvpJU
zmK+FBf5uYb5suoazhWF8/JI6pbhEL9Iey1PnL3+WiS1UBbkIfapJsOmBSZ18tqL
iIWJHTshN1kjB1ruFcClHVykNAbSR8qNWBPeON/k4VFrAQ/ePodYaFIMVqkRqO1B
RgVa/Z+2UkjmtiL0qoSMaVLfW0ckLNQ8n3PA2YOEFjoLJWww8uuHm6WlV424m8sL
wLkUwMWyzw+SWVi4Lm3LWpHQhuOsWpuDn5Rp0BIzB25gjceV6qRK2585CrVRQkkh
ee9FP7FAIz0O0LwyOaOjcrUKXeauaDijz7NSSPI+C9AVABHbbFRHbY741GZWzL9E
fdRvTIF8hchkW4wiTPB6VmAEHdP1bwLONKsKFKiCEJxSDZs1K+ULofjYxeVK1zc5
FIrS6FgPBIjW330GFSgqOWXmoF3ynusbkXW0E/70DX4xXsuhsoF01WvxdCoNCAil
+nXRJQ9oVYN6j+PvVzQOXitn5WVBcl3ltMjs4gsJDNJHxSzgYl7aklMDI0T8gmQ9
9yP4n5vQnrXFvCmeloyi2sI6wbotkUMi2tCBFpPlj03cWB2XavabIxDhksxrNtyw
edYrY3OPsdmFzbbhq/PLaxYuM78zAKJVe9mgfjHYPKydVl13BgyVHqqxNym/KmbD
3687bA+40Eav6XZii0uXWbwrDoCZAtpqfOhLHOyMvLdUTRafhT9mzZjhmYuKZQTP
Dk+5IWuoDGBAUfDjUsHpSMhcOMdryX3wSXceC5I5uFXCoVYVbclqp/9r4khNrMNR
KjFt3SJFgtTP15+uiv6MnlEWzIK+lMFB9v+x50WFXetTDSM/6xoD9wPE/KjPuvYb
auVjmzOQS8NCZO2q1HglXDPormiR/kKzIPWhSJsNijheqtCL8iNX3rlBbCkYI1AI
s8J3VCUQqME9Ij3a4LYT+YddmRl/yhLmQ93LZaMlMgOHK5Ki2YbyPH4f4ZJno1KN
KtTDGH8kPO1lMutJRs7v9oW8PxMSOfjXhGNPVNwx6VSsV+11/t0oUzCzDImaq1g9
Vew7R31Wv8VKIyMlqHyZJI5PXo5gIyV78zh5ss5qyXVqYtaPpkasuGRoVlJrLRG4
E1e4VwMTyhj5bBEwik10L+x5tkmSDm+leUs9G5bcgP3WnA40biPOcvz/rmDvym0h
Gw8VgLAsJCUYQNQH2PsL6xsfTGwd5k8Cks6IIvffIBqG2p/LwH/IyMmh4a58Gvqi
aUi+8qK4aI2p99LsGVh9Rj/WtjaO9R4O90AWQS4qZyBAOMan/nPpo0ZqwJPhisRa
VH3zWrBtIGBpC4J64UWymoQn5cezIYs5jQrZRuXk1V2Y/bX1P3OVOSYPNNdxjaZF
mqdBpFtvK81hRs/vt/RYkC5mWiXZa19FLqwRCaXPq1fsxuu3EdeUAIkbaJtlUnW8
1JnwskteQW+pmYYDAUtt95nLJLwcffpTUvD7adj5cbdANe7dxZroeXS1gc5FX3vl
DWcv1IJCL/gYbx1gTrImzETVrg20/m+vkY6tbvVOabor60+MGlT1WQOcZm2UcXrC
K7aPv6xQTAJlvAI3b/5ZZCZhGDdjB3dbj+L5IF+bNvnHz4yMDZkA74gcT7ZbVAw9
BfrDl/hYXOwGo8wyz3a7G0qXcr4sugwxzRWF8wHhyg0SCvDM+LapcOgs5AsZYOBB
bqxjR6wOZx8HjLJu8LKIV9MTs5TNEsXXF/k/EZ223j5tjZOQ6hv93rjHyLQ8L1UC
sgg9jayzkIHW0ngHzyqAIat+bzkhDCkOIcM9GGwksPybWFOscduMxH874mc7y+Uq
bt0AY+FD2tQtQAZsE5BAhKoCngw5kKi18pgp0+oPPKV4jgzT/d0akHqoaGfDW9mV
6eXv8RRnI8BVzAzCxXZCAAHvAwCYrr/T+/baVNcHiD1BpAZC4stlU04HaFHWLp2B
hl6rVE+PPwLuASxv+8eYW88yyJpAqw+7q3QU4qLplpgce2wkeevO/3tJMDHZ55QC
zsTVwiTXHBGiZ9XRJZmQOX7GHF0CVUmpQ5vRdlBs7QNpK8+jFXrvSoCVAOj8yoIA
QgHkZO1RRG59u3Ch2xCmGeFfgn6IS6YZ+v3HwPHIYushIT40Y75XUZHTPDVXP5WP
eQ/FogIfNgZYYxt/uzzA4JOhaTp7M4D2fhYUHB5sdHPDVaoTyisp0HL9Ywxc7Fnl
GY+RE5DQ/YDU3wIzewV8roojTxuPYdvvKbQsC4KpItrJxmNxDkyUUdvmFRMEDQ1d
GR0uuZ3yozompvytC68KukSfJ614TjBgmQTJcs7xgI1PzGOZWuDVnDWZOfawnaFJ
ys89SsS2XUHZ7Fas4QoCJc3McDjF8kQ6kvlklQ8ksdR6TLvuWFytluGogAfLo37T
yAMrLwvyOkVjMz1hjE4Uxdkcjz2m1+m82Shb9aNFgBJmvCv45ExEGlR5sBfXhX9k
1Zw5dx5mJJaZHW2Af5JtHzL3XwFZPrCdp6FyrhpcR2+bzPYG5UJmsiNu0zj4u+GN
YURZoN3Sd+pVzmADq35zffW4aXW7HgSpnRIl3JwFqjd0Jfe13H2LWvrNhiIaqx1V
r8CUtXIuXVl0TX8/lC6DKymcO4yScqrnuKDQHkoP87tLS2vm7BHnDwiA266LXzI+
1KAHXN4TYnHWVlwGxh37NDpOoK1R2QsEyhrrT0TvzA3TORwxA9nm1mSMZSkL2pWb
s1CFOqAWswCEJ/t/seHkV5uIv4rrKOq1vUbdRUS/NnxFwCLgq5R8fNVijtsS4rs5
RnxulYFvWmnTO64KUy42VccWQbQwWt5+ybDJ2yfmi3GOiOAFYztp8sZIZgAowo9q
XdF2Q44MfhFlAA53bTIs4M4Re+7dJ5g2P/KMyYL6KllbDT2UF4hleQIcanxgcjTW
2F0i5GyC5RG8/tGRZOxcFzPhiCwsuxZ9oZOJoGp3HPWrMwCr9f6oyB7QQS2Ai/hg
udaqLXTvlbXjGTQsSEFFW4BMBPf9z/Wg+feyIkmP/oa1sQlmzTd4IpHeNxMHWioa
24/yODrwyYYhegnmdrQfC8HfDCAK0tCNcyc9eWj1fwaF8fw3S3lET3aa5l5KFu99
V7bpSaCkYHsEUe4FCTaL+XVL3Qs/NO4tSRJdq6/e8VseUXdb2vUcDm3tI3lBJUV9
fKjYqiFQ6aZ+5n0wBmAEDaqD6Ds7AI67p5BGrX3l+ez0tV03gUpylIFIngziw6q0
QY5nsbaISWosZu++M40C0c2JSIE4IpOAtefPk187tABFnuDu0KuYx9U5aGlEdNwA
2L2Vbjz4f1yOLEgn0wjXf/ts/KB4nA3DXOWrexeedGceaN9/bB+ZxHuUYWrPPWdM
INNlkiZROAie+p/kaEFbg5Zd7QFpqaZ9WFbLDUiRddNawMsWUMPefDMo4O6EO5PT
vwQHP/risliZ9dwrY3NUhu4dnX03rINzhbtKVS/IeII9u/Ttv3zErU1nP3NmgCLc
Lh+ieDl/SmOESrJQ5ALfLnsEFLOSwIgbkoLJF/xvbS+4aW6IZKSSZgDAHJqg12pt
gx6LnhqlpT2uI+dTGiEEuEgZiVd/6G/scab6+cPsIU319IQSIwgFBVk//nTkw0JH
l6VHnABogDDs9O/DAPGfPb3UjI3g0Jt2zkGhTrcXJuthc0Oi82ZwekBPQi/UG0ty
N0qZfVNtUO9Od31i/nuxd7TTOKtApO4zxc3k90vSynzSvpCoyWQfMVOVYttbgi2H
LyYLNoi6ffS7ds1Al3pvgJR5umwsGyMJeRvIk30Dh13LDa9sNfzXU3HDhX0yTSPE
zgVpVIIOy9sle99ohYK/BKFONZpBYqRwKsp8MM8CnQC5IXIPSSSBcpeQL+DwiAzC
vkPDPC9ycm6LWqNm3+v0QIUwoEh9M4FpEAP2ckWdiBj/kWAVcbv7TJWsDKAipEjl
OY0WAw4zKADbSpCvhFF9PHv0k9sr2U5dp9oSIrMN1UMzyvycYiUFFilc7neNDqKc
KwH2oYRXDI8LY9Y3jA9JPL/wDBOyZT/ZDg7H0vPwuAiWl+qChaNbeG0hOE3igNeM
/wRwUWkMTbfGpHNZXjFgbL6KwKi28OV2qYVJu6JBewoRR9FWgyrjTKH4LpeMV6w/
TlEOC+yD96gv+uF4nJSx8oGE3UgQMrmuTOFfRn1ML1Wezi9UKejVfKMlOpb3IEWG
LREAoGoQNeQAj9BPLcs0Ceabg7ab1dVh3JwtwO+JjlfmDk2uDMBp8DkV7imhr+AK
KIqjXEoJe9gge3OY0++2rlHig4LkUCDYA0MSi/xaTndQDAxxQ6lB/kb5eDC7ZXNA
jUuVHv748cMpjX+vQax+kK2/cbVuL47AslYX8NlZNA1pdleIdu8D2TnSruM3n424
k4lGaLqEBSyaHcuLKJQQwtBNlF+uXYUtB9nNGK/6MrTjESsOibnEpsqAbnEC8rVE
Y5VONZR8FBRfQQBBNTdEgLOADcl6yO6zx1EZ3IV52/cfr/HP7yWK3qGZpxZ9oA+3
JHCY0kyJU7zaRwx8nR4KF4tQiC+p0g7wh0Bb3Bk2uGxTlA8KDpKhZ2+AKN+XXSCl
U1fQT7AHJRKRnDzrfey1ulUSn4JDfFQQlfbZvLEPF/Mnmp2M18Mqy7elhZ0/OKJw
rAKR+ktND00ctmePsC7JWDb5FzDEqH1LGTIVv+oqZdcXKyOJqSa1pZzWIaPwgF27
wn2dZZXhTPed2o5izBOKt0TOrCTJ+X5/6BjSZpw3AUMC8HnjPz+fb7sZnKOT4sxl
0hflj1OpAYuIxyk0DJsdqaJ8XuFgo/QZKZpZW+2LUuK1exmD3T8hlVw4mY00ZiHg
Uf+QhmrdepWaif3ye30a8iljFp8JN5/RVRbXZYKZhwDTCqzBpjIpvlk0/1fcQwrN
peMjQk9xkw/56AASpaLyjAJjqJ+OD7UpU3ANPTJZTLJlQClRtKgxlKdwdD+a3JEO
xVxesaqsUcvj7R8pLv1xrB20p/8Ioe9O5IeHO82WDK1LBv6OqO/9QGilMSC5MDV9
3ZIkjyIjx6aQyAgRWKjOY9Kn2cUw0eNls5evxJ2LB4jzxMf832chZl+uriYDkwko
9/ww13H/n5KkdeZoSiBZyiTBl7QHa2ptW5lUukNsBa0fAeHT2COAs2PLpMQJAvta
PwqQEwGmUE9OIi4O9DW5JUQZtNxBWnKm0zXTxyC/cbjuVyrh5WMv7qryWas/gYVy
1wxtspdWMzmDxPtR1JV/7o3uEn1NHEoaXAGhSd9wRH9/2NLg1wrjplwiJYH2ZtLp
AzgjPT6cg2BTU/Fcw3XdW2yjAcjuMcFR+zt80zu1eqgVac0XxKVJVmBdhUmYsKU1
i4Y2BokHfu96UlI/fJhYRawKI5zOOz5nI/dOROjsW+nKUe5kCMD8DGXEXxcjR7M9
yZrcxYk5de8dM6mvkA8f/tMMbsrs4eoCEUA+wy9m9TQIE2dOIwEV0ulc1xdwrHoF
9/fA8s61VEw0rJZUZQmqCxxaf7Nge8aOLeaAL69oMiaIagKooB7vyEG99kAXPXQu
pCM+mMkcCAzLBySqkPQPI6YtP3ibborRLXdLFEYFF1eI3Mqe/dOqlDFdUUaES1Rb
29QB5dNhAkwH6nrPgbNMgSnMNqyz95cljId61r0dBWHtC5yMHCrJCrl1+wT4qrww
ETYRYD1bKJjhsvjnPtsTBohpiix7GeMKJ1n++ZtahaFZT+F5AxkdansKHGHt5oAd
rLdFgqBx4V4WMzYakobRzCGuRb3UT0IARJ/htWLyyhKpISVo0gF0EZGeHAcl5fux
kqtqZZZ12Cg57NUYntf6pTB+mCFiooX1WOCp6Og24CrqeapAkiywuabq71I7ucMa
loPMnFaQY8JalMQRIosSs0P4ujngyyNujKB8ZrXwCQhHL/XeX8DJz92UWrleMqYx
m8BJSa/+Atu2MSd1B5FoDWgrbmx2l/ZaDP1SXRrlNXxYwl75aN3WUMpsUOgyDMhJ
jlbexfBEafJE81kisR5QOrNdGDN8/bYYilwfLOuWmiN4oNSAD9YM6ESllmR2JaeB
kgjkcB0EJ/PCu0xylafggAMdQFSlR6jcGwdZUTf57s6p2augyiQ3qFTs4xsoQ/6z
d47zbpr0qWAirXJG3NeXqQl3GMX91s2NwG0tAFODJey9nF1sLEmH/nVLFtP9VVG4
8JwLwM35GizKSdgLYP7QHKDza3C7q3ruj0vLfk55Eqx/vQ5vtfu883KsBk4HtkQ0
0AwfSF3yB9Q6UyqoGmOm4qwd2i7zYe7cqSERxZhP3UpB2I5oGtIKDBERHTpl1WO5
Qh4T+m9VHPb+Sunlgd+rykFsKBBuEetdFx9aMMLk5pm2Zb0OzpjC/iGLRxj6Equp
UVUXsm9l8/jw/YNmaL6Osd6LaZNu139p+Bn6niZQTNvZon1V2QqAs8152lqLqVmf
4ruzgNYv+mMSUqlIIZLHDZ0X1OIECvgPpKxfFDS3QBdlUu3YkCe6dffYtq07YGIN
x2ap5vEIzzhyxymdL8ODNRN/catcJ2nAzzEFMkHxot2eUhi48ptO++vWsapW+ah2
X7BV70ZUKDss9maj8Bgu+zlbyCMUaPLjjf6CDhKDxtcnZRNfQ3+iReLJBqK8j315
SnyMaehvLt67O/EpCa86nyc93XjtY//XsB6lwOOqIa0LbR/X1EmyVPIdAEz1kA9R
nF+7mbIrR4XUw4ASDbtzLS7dHSQK9d1gllST1UK0WC6h2lrRYH07p/5e/HLxhVyZ
VgJvU71MtI+t4HUje1ofCKllhwbKAHAzGhiyaMjD4LmLszULu8dfwbIU/mi9bIMK
BnoTbSgVqZqPSZd5qJPLPxFtHZOpQoz4UIJ1rFLKnkVuExCiBrqbrZ6UAkYtgKSL
U7SetiWgmfCqPR55vTgXBnl6+Ugd74+Q3VLJpWafH4vsaTFEiTxrbO8FFBNSJorf
QSXJ1erPR6y0vcy16YI/Ek7rONV4Q5jCMdb1nQCocOcFZhSfDgWywJfozur0w9lD
hpwOcGFwrM4jRe3euRbEM1vEwMEKELpt/4o0us7thh/d6rXBURGVFMkztVNxKYyc
qW2E0oTDiK2wskxNDNzdsMPE3jZPuZGL0Vs+tznQ+C4YxVK7zkfAyYUEszlNRaSZ
H6HVZ+36rdh9GtfrBD6CgJs5uWi/SsMYFiMkjtCRK0Zv9fn3XszvDTFR5yOlbMNm
KW01qj2pUwIjl3InQbBH8nRXMzv9Kh1osYUDAjwMxWahftaeEHZjaRlEarME1JXI
PjXKCKP1HyF6cpE4Rh8aKltTHM3cGVOjyau0qkRAVntckfVcxbJbcMUDT3125IBV
uLYencFuW1al6jlXxLhLNqb4BlhV6RmO4B5SCQAzgtDzHPmyZc6gvJCbi1p2ScRB
er3GqRcne1E5VTMQN3oRWJL9n2lVorHm+zLw0Sal2+bCvdIG3QnbRHxjvgMng9uk
MwdRf+/FZt5I0sQx5CVyHZhuF9QU9DND0l3vmjBh5Jh99jVL6/asDTYQbJrTN1OS
/3F15A/peRvEnpueLqcW9SeAsxYPKZPrf1z1Tzmhqbg8fJAgEdbe2uoE6LhTS1+K
AFm85WunPRn74mOWs7risnJKg/cGODMQBpoiyjB7nvpsdEnvitOf1iW0uLsl78Sn
OLyUQGQZO1zEhCsyTQxljxDo6QhwdmF62pnQHhnVD1IPI9k0xpch9mBtdqAb+ENA
VtjFZ+xHkO5S5Rofeie0gK+dQinIBH4OJzwcElzocXsjG0DhdBqMJ2BPkOBMtOgF
2mpPziruO4LXjNZOcdj0S1C1Ls95StlFosFyUnLAInGpTiJKlyk1xEQ+2jQnHF94
d67cqWng+OZtYnJ7k566Kx6A5cENQqOEDbGDk0SuEv7/0ResTYOWewhe0uo3ydnY
SR93HisxCIEo+3ttIWhJvAvKvHFzn9zYCmiJY/SocQyyILsLh79wG8hVVXHkr5Ek
5EEDyvI4qAgzGr/R5acU5/KGkvmai8HNEoAiTslV3SgquG5sBC8ureG0cxeGLCJG
wHwyEk1lzrHSiCUtrSLcj7WzHf6x9UPu++dJtBiSFgGWPVkFlvRqHfzUpmz2EGty
+oQ9/DKyPPL8zNNVYyfFEfp+wVRAq/CyOs2EERBlgisHpzQmyLDYBXR/dIyzzvMZ
uKcVHXr18G96bmDL0NwsEzdtN/VGKn3Ki2R82Q8zp1zUnvPWQQenHAwUDafFjHZV
Vza++d3tZ+FMvfwsRX+7hfrwnuFX0bASMxs1SsecV6Ft8pf/uWWybjL+jPkn2MKr
Qnoo5PfEUaSvu/bI6yOXq84qgPtIVJzqaJqZrbB4lovxI9DMuG7INuTJ9uJuZgVy
YRT1eR6XHCddacd7DYYDft1lhDZ6tpPci3NnoYvioDvQ4ErBvgzujJZl6QmxrYds
S9sLuAADXRYXEvmwfgBGLmof4RosrM1GapMnsx0iJ/S+bkl/BhbqKyIQ3gFngt/v
LtHVKl5VBTqXHzM85H4xi1DFtV0MNtmaoQ5mKQL5hdfbgYXGhXdqbMh5Xa+Zd52x
xQPQaQBj8HbL+QcEammz/0d2eq0RH//mPqiDgkR/J5TNzd3xbavCTWVjjOWHRYdn
dr2lxWOv/d6WxFOM9NSiFlxyQYBzTMZjxNnbjpZj2G9mbduEy+qeLO/kCCE5C1G6
77aTDiu7MGv3c9OCq5xw8QpReGPvFvmLFZze7YbQPil+0laCYGBSFLb6D6RQhV+6
VUTr1yC5DtY1lNIe2KjQ1jpmDh9jBsXyQjSKTI7kjP7pCcMg3uYw2OAxOP8Ftw+2
4jBEMNdVgSJMhO3Sq3Q0OsTFHQVtkh2zPhuFdVvscWlan4urFAi+VAxKr/TdhxQ5
4Jauf8GCQVPQ6PMHBxDhHxCHgUL6lSuFmc1mU2dN+ElZiKUw3+zeE6JQSadi00uk
p4ScolUfV4ZqjyyZj04w8rKBxQ8dogZSM3EINnL9jRFUzzpDloY7MqGqmOVaTQYP
0km3oACzoo8sncDlvmg/AHZ86aSO2zkTuIgmH8EZ0aQAKXeivlevdUo3nn7KKn5I
6PKb4aYsechrMkEfRWWa8axY2JZLcVYATA5cvhm1h+tdnM+mR5E2MIIB/rQhQqhZ
3tFqzQi7DSddIsW9m9DOBO6aSDT7K/dhuz3sG58sHJ2tlFOoMYlO3B6UAJ95NTur
vvIzUhnOOY9vcnH2utV4OBtxvjgtCKmUEk1SnBpxzHRUwRHVTjGIpv/pB1GyQ/Gk
xr3fSjqNgiD9hgfbeufx13DHWpgoqWp91HKX4qJUc30nY90DqRozAnDDT0PlfnkY
Q+LQRCYza4ofWCxTzZtHzLYPhUdNrwxkoi0n7Bif7vmitwpDoQxXs5TysjOWq8Bt
0+cdrrx2tiEtUtk1m0xV53zCQoHPHjsXJPAB76tzt83SUlPg6LAU5s4pmLIOaYhB
jfoxqDFSWrTCiBV9P6SuzObHxQyLGlxx7l5KslPGyAyUIId3C82tXscmst94XHtv
XRQtu/nPETcLQgj3ghtB/nGHNCb+YbXGtpgAZTGBPbL0xz3CCRiuGlcu+qtfksGc
iL7eAK8J/6uuBL+pIs6MHvqSscY7xB7+AZfF/dmqXxtwYurk6omCvOGHyWsugd9B
rjFX3hkS9yrVIVAiBUgqNLg+s6BRXY/PpM2MB43FiAnVx0iQBepkoyxh+AyuIyVQ
wvIXVn4zCvi8UpW6aUnzoi3ljM+d7LqcplxtSRkAlTZI4ikknDmjv0EubphNMPvL
Cz7fXS1twf+BP3noMNyP54viZU2e0HcqIBlZzP4NIgKuMqkZyreUQQjoxgnr+YUi
f3kJI8/DkvRkArFDSizv6EGGKuTAadcEDFWlh/UOFsFylCFbEvCPrVDAEo75B7EF
Z+Cb48f9gt+NgqzGY4o1y0EWMk74b8lScttcyNOmAyBn9p96PeOOvuOBfdYFWjga
TziOWW75KPR3dYoLtVmvgt0T9iG9/t8hcbuvsJwvdgHbnIOvSEMvSHeHOk3bNBKj
iTuLqFpNK2FqaAwHp+vD3Fy/KNwRqtTJEj1nqt/kVwJE/bfolzYqlwbNyWE4dqYl
KQgTU5V71+yk3BzPtJiIhqyNTzEQdCPKRLpzXtfaH7gu6nFzz9d/ou61hR8P6rl2
lOuS6IihAYQU4ItYQCbqrIlGNVhDFa8/ZJ2Qs7CMQm7CWtOVhB/Jkk80n+wmM55c
v8oIFz9QTyjcAzMPmcQ638EeXT4eFodxPGwx3ll4JOJHMU3VVuzvkukrDDHiifls
wuktcbDGfuXH4Jk4h7aeiKVEn/86M6UXmMN7b1PydKU10LyxgQjEn+gxilkRbRf+
cIz//6eSFwC+RXBBcGbDTigceFulf984+ho0Rk2j7NEstl052uab0d8NXBgzKZVK
piZio9nDMw+mxjihEqxtdgo5UYfqviWR5tJfjjH9m/nY597bW4HhyC6ssfNIDm5M
DM8qFptzNzI3h4fBd4sOKmaE+PLVS7Gh8WpBbgsOAy+zi2KMmLlZQKDZVvY3r0h2
mo17cYRn69eui3qka3X6uXtzFXdsWBbRSedgHIvqlrZmB5KWjqO2oACkB01E46Kq
FDnrHb3nsEGbLfQmoC1uB70rZ1yn2fECdVDHx9EE2KSzNv8McxL5vyrHjRouFlYq
16OOgFSxEQm6xZKFjR7D3TBuxkfa7kJCUlS30S8nWA4Ax+aRRLqyjx+X7nFUdLFW
hEGU+UtPS5Fe6nkF3wNO7tyPtAXQIClj4LxAWUPzlFM8j92BvqewwrPZeJxMa/Ir
NMq82WSvd17SUMuInuKxkLBS4+kAQoOs8j6O/ejqzLnk00fUV6C1ewf0JiFc3Fz4
S/x2un5XyRrbBmfsOdiuiOYwqw2IhqocSAZ0S/5QoGmiMEg3iubBOdDi3/e9du3n
haIKabBDjwfrFexbTTQP0SX4SDhiDiibedfm5z2QQNqGNkTXW9umUK73IGtKkqtZ
5BnX3zDLp/kFzOxOQ5I4C2jG8sp0rRX/3aF6E0hPD49lE/2mOge6II/ePlw68FVe
Rn768STIUmeB6Vi1oJ9x8dI79pFr2UHgedZN02JLYPRkt5bnOC7TnpIgbzfpmjvW
qhEjK6TXoCZZsj+UQ2ofXi2EfUPm7GHCTRkjmOuZC+21YiXEuDOBribwYBRj0YN/
fTDSKyn01n4wB7WiCpTpsGDTHypRODt5t58NYSENkWJDN76MxMlOML7qor/a3UuJ
8KwPDbFVIgu+OlWvx6vJgGfdchMC493DLzUIib7TvoTKJzE9KBOtqhvi5Tu4LPVS
cBQSyvICfgw7poU58mZqjUWzelfqNibq1rKyrrdywrB80HXLIBwEvH3X4zbxxNgQ
pOA2JFQG0pbENjH5MLIaypG6jRA3QJbJ3PKZtLoc2pPkCHoyffnlaYap4fgwxV0j
iX66x9PAFLulzxC4U3wiaMWKYlM1gbzdVUl1a7SxcljZGuM2vuKH2GFBuSrcSh/h
Y/MYrIOq5fqOTtU3c3mn3uH2x/FzxUzX0UPkuBOM9sGz/e3952XaxRuZr9stfnYf
b5pY1DsLfSyx2ucsLQrXlP/OHG6sL4KllPM4pLYP/OGlvXI8Y/YstUDOEcj/KV4g
k1X++1pXsmS5KcgG32HcPCHkAt/eZkimCTrLCUUz90AKkqTsQb0Ihj6u96d8V+zQ
F+mpAqNM8gKOuplOpZQMuun9rrX+dsudKA3caYywOMBjVDc6sk6y9jmdOLfkTBe3
noNIIKt1fwQMrb2tgUh6E17e/E+IyCwuWmocsy7mVoswbw8ZgiZZbuQyy/mEPdKQ
6Gk8K7ixbDq+pgvZMTwb8mFSVq1bPOBFcHrVhiBr8IYFkSqFSKRy0wX+PWL6XIoZ
321SaS1rVF3GfHsl6ca4sRp+/GdIAaR5RipJgm+zdVU7WI6HXU2VibOLbrH7Hjab
cOkASxoSm0xyrMtwLgIvbJD4V6gkOmwo/mnTVTYJ4DJFXb17nLh0hG2trYpTA9+k
rF/GhqcXxdmR3IJHRz4WVb63rmMIEuAJhGUnVSpc4lQp4pdvvjtwxew5lT0UC1FD
+lHTkmwBTT0ynTqPOenvk1l7g16rZjhVzaVMW7TcFQWG3RFZ0MLYhJWDYyBalfm0
G+lNpmBANwuvRNjAMMsbBK05C/YdIZRd5LTbmYESpICgwOPZUsc+nPHxqEm/egu7
dEeTp7qbF7Mes6DjDoYg4gD63Qu57jebeK+dpzgk2FlKNamtnJ6Z9vmN3mmbNpoY
CI5O5Wg9zYNI47L8RCBSH9lNrU0u2qN0EJBGlk35FJGRh2DYzSCqafJYi8+R18v2
ngao1zc2E9eVfAB00dTNYnXKVOMw6WmyVHDizNbovoGdLarO7qk3G0mOzk+P6+mM
e3aRZEE1ja+U+QhvUHm14hLCYhkMxzh+jZ3Fscy5YGor0KYIhxi9OQRBrwL8OVOh
fnIMWnR8DpEtpobIlrFsNGDsFWsJ9gppkd0QcoIp7D+W2RaCtCX1kQypn7t4mmoB
UJQkATkcZs+7SZcpOft9dljE1LsDKPyYRgxgHiQBeEJnxIJHe6pOvOsuVx6jpo9X
1JVJjVRK+EmruQXYZZlTPYII5wL2URcgNx9QMjUlfDczcjposTh8qo74g89Bpyh4
LUaupd2QLoPcMCNKs2NGDYWSH5p2pq/82evsDnd6z3wqhse43zH1xu+p0WqzxrFy
wYSQ+0Y7tq6KCUfkXJJqEEk9xHJjaIJvKSMSGQgDGJCiAqJib10FaeizePVu0av3
TTaND9A8xRLYsnszVfDeMmM9Un/dzRzgPZUkpVuuoFCuLL4G1vceu3i923rJPWFK
LZ5HQ6ICCSbsgUacMlQoCHMDDPXyOVQa7KfDfLXoK0H61MBhXFwpXudFmtp7htoa
9K3fGf4KBDUSJFwF7cpx/F6m2EApJ/JK/gjCjvR7PPM58uA4rNr2YjNpZzkSZKX+
06HycTCNlQ6e9rkvSx8fZ4aeiPVzLI3ekcCDijcQLde5n2Q2wTEB9iVn6qg1UsYY
i3mnZpNss+j9jEiSMOJlL+8wUVRa5jdj5DaxF7bCMnDK0H/sKhmVQox3oirneFep
LvbgJGFswEB3obM41xJSege3W1XP71X4RjEq4nRysZIag9k1/2NPFeDnWx+Jg7yO
VMa7SdFk+w9QUKPplpoM1vHRcyNPJIVty0FcYcWsV7k2FkzCVs7kCsknAxuDHQnC
CAlMQ3O1vEak6kiQiAHo6/qs0kv/PrBmynIsKxMHOVTaEgmEgYyIi+4axKteUnPE
BoDXDLR2BnGFEGIWzaW96zkLuzIpUBVFpTHohRGFkvaTeN3C4H4sK2aYAlWk2ryv
xnnEGsyl5R3CEFkTvk6KWHuNeJVFOPOMRZ28mA9seSH0kF6jw1C6iIvoIsIJ/yVo
8/UKQr/0azWiEr/PW8GuC2HHh7MfX5+/Thwo68TH4bpS+nSLlGUyf5xcfn6/XOlf
On4c7mskQ9FEm+PYSYvPEeonYlMJjfZOAM7UotD4KqGXhCyH8PIAQFNWQlR602qj
sgUjgfExYXWue6r2/IQ1QZ183YlzLrgChyrqHSpzde211caqSKUWcsoetLTqhcJo
+asJQP43upzN/56P10GfQh1RyuoKP5Li07016Ivud3Rmob/ocSCnMnyt06x/RVlI
KaJoebAbK3/GrhSYQu1BROEJpXdF++sTnRB4EbCiuF9jjJNbm83uH2BzZ1mpC+Fq
Eug1Ac1Etq0lsgS9OmTc5Of5TToFIbgZn5hSgMy89xqbb7QJuZbUK3O11EDYgYiH
8lSsNB/GiEOy3c/XrYjKvmhM1AvTMSNGRVeuPji9tdOg5aBnLvKyNBibLyohjnfe
Tr30fAdFO270ZNBEGl831z9cI/zs5FKVoRMebe2eCtVLi340kajr8GFc5ydAQDxK
2a+5AFrlqUrOyYqWNlCIuj8TVYPrkl5/BE42Vsd7yWnF2xDMBRb0zUIsh6CcIJ73
68GKgLddgszGucXhvQZI6sn2XDxktdR30jf64yevxg4Uxu5UJjkQHpmGeVcVA7BC
GtdfnNIAOn1bgmrs7QQH1cn4KZSvM7VtCeOcffoqD6T9Yb7B9jpiO2ckOWnxUsPb
+/ktlX3XeJaWnvRvCDoCbq6lOoHx7naJBMIA0vfrNvMHhwTatbilDARdW767XO0n
agFEeOJQHNMmtHKRxcfcz43PcR7OdlK+sX5u1Be1Ky+Eb7dxorxnhs8pYII9uwR1
hbAgg2QZUHntzyDrgxlzBLBiOp0fcRB0On9m1/Y15RNUqI7BD1fgIM4jT+kfjJX3
vRYgK3mOHaLVLrLq/OpJle/g5+Ffj6+bU/Z4aJtUtRlMjAf5u2bBX4DT6dKFR74H
KBNHqGEURHFvVVj9OsrkgtwFxenwvwM1tGSz7p2IsWzSRTGtM6CZMoj+XcQPiOZw
Lwp9OsuYLbZpYoplSbB9bMIKENVEj+kVzSLzBpEFKlDxdrWIdPk+chQ0nSD95XiN
kbhaxUpD61iHg56zgFG8gtJzw7r2F0v3d5mFARoCrIAEFupJb6dNB/qg7Vxy0/5N
kyOOBKX6gUwg7gpqrLImoNZv0qbpWenmHu1Bryln01TrwUKFzWZqfzwE74xr9QSK
VBGXuXp4fHA9fCuI45UQpx+a9NO03gzcyPDJ+Stl4GVGBWgvnBWng+qUdlArHxr/
MWOuvHvWxsfddj7ddeSNfDGhbaJ/aHlxD5dR1LSx5+YYYJEWlJDPVNKc8u7ItNMY
gTmxZoMhLD43i6Sx087m8yjiog4RvELVGCqduUiboPPxkmKIVufe1Hzt22WIRR7q
Osc/CmdyAh0mFtxJIc8iFeT0Cle05KbMc8FMPkk2CBIoCs5e8QfaB9SuO8h1f0EC
vvGD10MoSa2LAsNVnT6DdwAMvadMGwsWGyZfe8IDIxNNPq5r8N+q7g0aauNjw/8k
EWsq6jDDl6zzawobINQEBZGdl4iWn4aT7pJ5RW5R+Ojsj/tLr+JvVV8PKNl4SejT
F1FOzEcW2YuvDVGtqlidnnHfTsmILJipYZgDxBGn2VWe4t+ZtSYQL+L9Y/RzwiTM
5OJc3FQ1DyqzwuhkptsDLivMWi7hrixbg1Lw0kZL4H4Fu/AwGsBSgt7gjn9ndcfW
BxJXlP+uYJ2SqItjUr7G63BzcwKCCq5TitWYw/8roAqsetARCXdHdGqCHzW0dAsJ
wASsTC999sqs6x7QbdKr9ebG9AxpvZj90TvqSelKj34AGHoT+NNdAz8Lf9/gHmIR
oBRXdOJhx+c4IkwLCDtIIalM/9AOpMakkY/n2DqkBhzXM/CceEBk+UtQExqxFSd4
xwjQt3TSeYD1bRca5F305RT39KqstEEjErmZkLfIA5YCWjhjnq7lUvykjbSPwhDh
J3WlSHkPAaXi5UVHxmscNQ0Yys2qdVtZElDqcoj26WoPU9gwu1yFqEQLvJpdh9A9
KnjKHlP5hC6byKCEeGHjnU9K/9tk6bsQ8HZfxr9bofTvDZpzLztjf/tEPhbx7nTP
vcDuhTTuFUQzrRlDfH/sQBal6dg4xPzd5sWmkfdotn27X7zVRUGVPderPtKl+vw6
nCLRavB/tFU19mBGlzLZ7fj2nTyMyMmzBV/ZShDP/4Szv0uRsfG0qPoxHtA4XYvs
h8E2drkmZrNDow/kx+SaA8pE8gcCyMXGWtSfTTQ4xJ2bZLlDeJzfsnHPKglO3Kie
rvGJBophsjB8zhdFM19LbasV7V5mvcMjQY+zt6/1/bYqY4QJFaqNUc0oQ2PfPoVd
7YE6oWTROvbZKPdRyOQGnF397LqRuWCYOri+8wwByQ+lVRGb/PTI3Ld0pZYjU8wU
Tl00sRWVsCmtcRT08KaEPxbyM9rMTGg+UyR4JEY/SWY4k69/fGqmjK+aM2Y/nu1h
ttnrHzJ/rl6kR0SrgjqOVgCI7uxQ83gbWowSIxBbO1Fu4gb8BdaCAMlZI/HiTNz7
1Zdh/yi7txcbw5kQGo44YxoXm5XBdmCxzxbJUWGh1ZJ5+OAcyQHIm9L0JkUDTERT
3MdSZglvaza0haFyZJ0p60jjh/OQmDegL8q+eTLkWgngmz4oQgjoNE9Aus8x/7gn
IhIYBGr2xfVhFBDORSrexhPtmAXtuk2ZOOOJPjQBczom8SUmVUPbnuMZpi5l/SW0
wl7fSAOxzmELJ68CfrqMcEPALZ9Rc2IyIsJdyUwknzUDviqI+hCxD93QpQdzkSSM
lNtNqqMWzWD6Zd5GrX70Gqkfec0kNiYEn8SuA9og/a1+ecmldNekTHJsTos1tImJ
9tc9zGMNoiUCxEly+Ge10ZuKDYoqhYyX8QEsd8SZQmZXC2okNaSEXSMenfbZZtKh
dAJcQExUHtEV6REqHJpwvrunmh+keGuNXtJ6a8QJVuDczCgiVTfT4AGtEUyBg747
E9xRLCMEkCQ06ZWFOzEv3h6Q0Wc/uKjLIXZCukMn3i0Cy9NWvguaLbNY37+NnbbF
FMXFjCUBpglGCDb9RthTjhVpEnc2m44NdlEsjWyytNNqI4hWGqurGHCGip8sx10J
rkcTM0S+7KGGK4bqalG9Zoea/tW9Hg7YyrsxrjV/kEpcejM0X2s3Eivwss248DLm
1Sd3lD6rrBEeBvodXnSkwKypOOuyiQ6y3w3UMK0A4E7Eu6bcFBdSP+HtLHi0U0nv
cD/8SwgDp5umLmwfLqUnyujIjQIZbrJPu75qQlPEU6CP5lBeVpd9w8cPktW+c8Fh
E1CGud3sT/xs6tHkq3h73x2UD6ftiL5NLewd1rzHDEJfp7pFEtNC4xnrr54bHevU
57pXNnhwbsktv9mdos8IAQ38yYg/jBrDLQ6+afpc3VGZU64EU9aE9aqRWhDpmx9m
/oqQP7O7LKt2kdIEetHAOzBZw98pcPUgPbOiqCGK5AyieqYlSslNuiZ4+5GcPqhk
Q5ooaaIPsTBK5RlJLsTduLWSnVkFD3ONypXq2EU5k0XW7xFDLJ0yHk0AK5UoXzQV
a58wqplSMXAIBSAeTfrvEdE7W3bnDE56jOHWzU9TKuZjL8pUZ+vEw0cAw+rmNf1m
JTf++K1Ykuw+EKjLsbdZFvbc0+qgAb7qNrD+yBR8NY+PhRGZ+eVZWxSI8DwYn39w
hGTsOGISxtCey8KqrMIBhGPRvesGzZSSrKdFDFBI3T6HOWGB/YyUbi1lg//GkFh7
KeLbms9b5muteiLsli184vcNMLPTX5N+lDr0PAZ8dMXZdiCCFg2Iiq7bdIIa/k6J
uE1eh6Y8mhCCGV8l5Vd4PTmp/UUUPS+Me05KXUmM82m3/L2Bg4owImBs9EQrHgnr
zzKCurgbbOb2pGpaQAkdXi5+CqsB7VU9Es8KvlsqKEDLTs6twr6mO4lseH5NNOfx
X03cAn2+/0PKPPPNXcyTWspgr2VJWldg5tUp+5cBtsO7fhnTJrbGgzLkBRmOz5et
GoHuleSaAMVgAl/1YMr8Ie0DbgqRbeRamay0jVMuIqorskCQ2RX7WGOzZN/yfZkH
aw5PYZ6oo0SYOKZS9h+pmRKC/I5kSNjp/B3gxMZ7HX83je0DDWkAP2plqEc0rT53
eaPUfaRCT/7ld1FHVqtD//tQzV6H8yZCkrzwfTgyhQN6frNIU9JaXqaOrWePfTdx
8HV5tCkWa9NhCbD0WEEGQh1Ctx9rDYqjdIIAXoTbjZvGei7mq2qH5QhkeAWTQMTV
q7C4R/brUDLaYNa0+YINRmghOVfd/yvRTlvuTbLyzTfqRGH8PD/8DQcGDY9LcaLg
fXCoAPUtT1WxnwHBT947WAW9wqeZkNoVH7h/c1G1odEJwnXaDljVkuTU6DI5Bi+8
jWnsKYkW2C0HQb0siXbkMUv2Zjzv3Y5zGMAg1YnISG0Px1YYISYADYun9f5RTb3V
eL776034wDFGR7cGCJiEN6jRoGF8I3vy6KtfAh6bFxs6rUH65M8dgoVrPVDoOle4
0oV4ygHSd7wrT5PFY9dopO0dGz7xsvTvKLDJFnZS5uWJJWZ9upVvDds1JHfFjQ7F
siMS1G4+xpcEzx01fbbXcVP9SBhKwCR/X0uEjlQ3tCkPMo9dHLrXL1PcooT017eq
SKyzFX631UFCOmExlG3NdSDJyE7+X5CRVClrQsfobYveiM+mDASZg5d5Si+tcLai
dgzBwtw++IHzvUbyorWNIVVuYxGkiF6blJUXPybDPcwTejW+R+daKpxVJE1AWbpE
+TrOv5RST2Ez2R/aPnrHqNA6p10uFmThh0xxbdX9fS0a/1fBuVo3RDR/1tifWL8/
rTrMqC9ADAYv1ZTDEDEN7jnpec+gHVgcmUAd78lGp8OPwM+ybfYdLIjIJkc8Lu+h
hWO3NvZ16ohSBeniSgP3RMpXdvx62hfFAUgnDFY/FGZqOGUUkwO7D/zqwQVL/LYS
7nq5IcZQjbt3efXCH/ilOpqOe2AAnJ0gd/3lzYjB4KaMYjhpFlZCwbeluY2JjqAH
XKmDIyt1YNXf+1YFs8shVS5CN8fUwZtR3F/Xer0cHSqRkFASx6lwYye9avMRqBNU
96bbMQUwwGlcCR1fyA+ciIkwwE90PaHOyzEcYaHjgopOk0jcGOZYDs/MBeh9E2Qm
amcXf12m+U1GbVri32DmzL2Foago1xUL30QEwb8Yjilupit7pXgOGsC0ZlaQkqeE
FDeB+QO9s+D54rxv4obqK9pOhLuf4yd5mu1+zRULmia/x2+DCYD0OZpIVwHdJb6A
XVBoC5Y4nYofwArG7Rl+prTI+l9tk0PHJ/B6nHx7okJ9Q64B96e82BKydAImJroI
W/XDOuchd9gv0SJ8BtpsbUzfHR+A1pmhUPSSlnqdiluHztsSSnWCY1WqXvpGIXYe
/3fskWD6F8fPjbiUKTGaHku/fAOdnSiNtyc6uXR4LS7C3is5jTlyQ4xgmdjLUBGK
woGFC2JCiNrp8glZADuKO2GO8khAznmwspTURfqoUlsCTZUXe1F9YuEVI3ZsMxhZ
cyzkAcvtp1MoyDxh+cyiqayD3ZbgJq1GlSZtwAJ5fNATHagLXfvA3Cox7LxLxXjo
TzAlEcZixbMAlrYWCOipBZuz7CyhpqE5VrkXD0wUPxeGsAQ658/peCalNO8kaxkl
lM/xvsgGtUDv5YvO35ubCFRqSro4xa+0mZzCMNvN2paxlaCdl5MqV9TxieHoBgQL
rJM8hPUlvFVci2JFdChdGk0rMmYzrzrThHp0deINA+YhBE2eC8BZpUKBrxACfjDL
UnNv87G3DPknDiyfrhTUojoSlTrP+rrXG6n+QlQQIvjHMbreb/TXqhCGg7sh9Udl
7aiKQEO8HQaA1smv55ROCM2fMBWpU/sW8K5npiNPNIwulPQrgR9wq6TplaTuHQ8A
BwrEU30PbeFtM4vDSq9zPxgEpGHCz+GnKTgbuQZHmX1n+Ez6lpJH/wSeDbq2fZOa
PaBzpiVoF1B+pIoNa9j8U2zsR8ayt7g0oPU9Cky9opsWhj1IW3o+FerRY02T+tQq
Owlho4afLlrbBvVC/OoX6mrTcKuIS15Ov9lwVlwBuB5/+hIiAzBHhiH2hvd/7L0Z
t57HgZXUA3FgypbSPQKu8FXQWAhYj5Eyl21wlfoPy/b4Lj36bQbnklh4SxFAIGl5
HbcGUh17aA9UjzTYdt0LP5jYd7huthw3zIuY8XJFl3iT50Wsi7Wc2Wfi0uUeH67y
mtmYNOuUfGX/9Nz8vnWrSOIbpZbR7gdKdQX8MBiALDbg2cUJjUjUhHzhm2pXCy5g
Vj2umQjOR2OR6IHJ8JEAnFlRINQVXx2WE8Zegs49SSTZb1CiGnKcrg4nR3cCOn++
89T3jkpSfY1uJw0OFcV/SdEPE+QcIBzlzd/WL+dpw+q74h+qUUlxPJ/wPrzMAxhK
/VaNe/NmaoApFQdsXYNEePeg3gV96eIzxK8wuBwAy+v1c/MEvZkQx/yzZyu1h7Ta
ANwZsRs17wx6v4dxwFfk55cazk3SZEjifKO0zLNZrY3GiyJMyiOBQyZu1dGfam15
j3bUTut9l1mbl0BzB4GArhRj+CB6HKBw030Qo5aYFzMMfulEuyuuIvlyA/WD47N9
FmmAPeNzqkm12B2YLK863FydLDcImlwO/I3kqQ8SmjRNIyquDAGAUxQ/z4J3xz6x
2cc5ifxKYlTO/9mi9kdnQbrVrk65nIy28zxLzquIWY4bmG7h9/DjCKJuqXbsYP03
/wNY5H+cfUVGBASAo5w/Aa/skucFikWGmwk8P1iiyuYa0qD39Dv/Z9SYOi8+k4l9
nalC18JXyuzK2zxUQO/FiGFws1/AXmHrcX88221AIYODkEVYF8qZWIpoGBJP6DTL
HKUwHFcUUujcnY06Gd0ciCIyc7ENq6bMP8RDLpse2QvRC3/LyItuhiFuYtf3ipo+
jjru3oKyIcuqaQWr5cWCvyqT806Z6wfExei961A9OvcFqhGQBY5dJcsHIEszgtEy
m8sfiZvusXyOyXcDeIoSOdsw8Btc0NAR9de1VGCnehucR8np6AFzKvfhWFzMhDtY
wd4mh2bYlWyR1YFHyJbchZy0A4hHtrckAyDwQ7dLlMfzzQwYMfhQyBm0e1al6lve
b49smSJ8HrkocVbfjc6fjAlYfY8CJZN98DiKvHF+mDsAg0UVS6Yde3c7JW1B+3yB
D0YPEm7TvlfIBDdTgb4kCNzQt/pDNQ8HbFPyP8oo7TA4fzfpWqlVYAfx1foJ3jZP
DsjhAJB1Li+ZzV4/IQ7yX0jkgMym29BUw11MxHu7cTErU4H8pkh9B61zHgQbqERh
bIKpGutri6iT3rzEOT7dPEqgrg4VIoOGRHMjTRff20G94zjCy4P+s79J3T14PDXe
oON2a+K5ifqLCoIraTKW0XNrL7ndH1ynceuUvBoa/vkvzOWe8Ecfqxl/xWaJwJ06
HhbTZE1GGa4rUl0khQSfvyy0BW/2H8UQvekM1fEiP4LC4UwMhdCsQED9iCaoAdKt
yXYOg10ZdrVmcrnaRKa3zU0aWmnUM1fkWZJcatW6TdoPBklhDnCjBOwJmecVnQwx
9e6jQuILyLixBC2c71z+g88F943DIrh3CsKoSoqY9U6awYguFBCeGW4UsH66ecCM
scH6XMKmFFCPyGS46vNOOLVqLmTZkT4I6Wxc164xJG2zJJ/wm2aeYOsKKiRVz0kp
LH/NqpoEBjUxFRWLQj7lUbIctuxQSbWcoMYjjL/LbP9KiLbUn0cPUbChzNSPbB5A
O0f84nAeo/9ZYhLBwwXvhraYd/l4hBGo+q47+Suz2koxS1HfXKdnr4Tnd10qi1Rp
vdzXT1sY8spo9tmlIh3ctj1KqDLE0MgvkRAj1kLCmH6B4q8ZNrX1EWG/SxO3m5k4
y7/GUXEoBXu5EURlgxjhzMjt0e3qBeaNlStjFzdpXxpjeo6grtlAUXxbM/V5q7ku
9hzb7vz528MCsrE+FUQDDzLTXzODMhvgHCLfvfhBiBYo8RxJPzydmedOc/g0qRE4
6oF4SzT4t0F0kun/NWgwLxJxkKg9eDCwbATF9sMTpESojJLrfMm9vpDa1n85+4rG
BVhFTqaTzQ61B+6fHETgWjmEhZaM8AeVo3xTXpJ4cylj9tyMGgMgLCWMbLrDqm64
48SrNfzqaTTzjpIctorthnVjWo0bWbmjekO2Zw3wcc0ecdxgag2D/7j44D3jZofj
vBEuEqORZ9k7lKvhCUMvVJ8RbqwiLhufBcn3ZKx1UhOsGNX1G6bTVhsm13Ru5Fpo
h0/hTwsIWiNMCdXDFlOLUQavMWOITCH+EB1aCf8IoOFKmaltyqoMQkmSGJT7XLUz
rfCyhMonjXyJI37ShJNQLUGgwS9Pq8hQNp+KYzENSDqQTBoM0YDh61yXk8NIsoYo
jiw2IPJZpVRX3umO9px2dBK+FivdlZvb32PGlneUwcxjgocEuAmcFPpc8O4BGRIx
E4B5DS0nd7uoPumpdh8BrljiTsvCRHdKCHQKUxRRsj0sg3a/EKOpsLY2uQfjOsKJ
ws/cy6TO8/5Jct8KbjwYGodC/w5LpDSHycR5DCmMzsmCBLIPxQ5PcYSnpLH8ktv+
m4+sJocGP71K4uAnGn5MmqyNMRqI7DuYoaZyeAvj4Um/ahoHssbbgm4pMX1xvdZ2
TxdxKZucx4UFHTXR6ijGdR/Ks0Kg0nCzrpS95yCM6rdHXW+qZLKyD9YJpfqyaEXv
puZtsTJTuF9wwr+aBKkp7PflSFN7Wli6YHp2nN4/HkMNyY3wZZA+l04NBABVLTOh
+u7IGV9mbmndpt8gqH0AQzOloKdSM8Zf168FU6Eb9ufFd8SUldQWfG8uQxHdnIYx
Fr8u4BJhHmi76lVy4uofQEpoW9UnBO/Bq5OF9iUkqPyFo9wh+/5+1g+hBoTQ9aXX
v24WprivL16Is4V/8vGoWiGGoKHjTrDtLJiI4dAhMyWft8w96AI7OPrnEaA+An0r
2nljQKPS1G9b8mjO1S5DQ/QXyi/nn9lenr4bTWeZaUPBM8vkhBeMySnjI4dGQCxf
JlWsjaLtqtv0nhx75FfTmVG0mCQOVw/lfNiorQPEmQ4g6Yw8I3+v9yeFyl40xpvL
Mzv2VkOZSxyma0JnqaPKqILhSTQOabAseqchhI85Tktrm2j2odo5PS+VcLUBx6KA
rgQaPyjumVDEYgJazeB5kMMWBPRWDWLWThjDCwhrKarJFtKp0XcOnA9mL6mPCPSt
EYFQPDPuFL19Y3CWnzZbLICe1xWqP7Hqdn46XogJVVmdsucTEvq/86UQfBwBnH+u
otOycFhlfPHIbUPKfqhWSNVdYgM+rcHhzf2oEDwKjAKOtCyFn0V5Tsy/SwZmaI1e
XfU3FTwrKyC3h0S996SNVMMy9NPaEo7lxkLYTnQorK1bOG/5+/tXZEyLaqs+xtWx
kpfi252JC+aIbaNCApTYlpLUPF6k5llEMg1cZ/Ss9UnX/BCRghLYf5f78n/Cm97p
RnMY5arlivGxWCRu5qtlJltfnAWfpyEO5GNNJj0BH3WwooBUSDYYMj5xZtDZlfTZ
TxSJ2cuTRUa5aOjxFsbLsFCjijGUqlrct6SjyQFSSjhTXoRvgliUyZ/znUo9pxWX
/d0hJyMjR+WQsseJG7LR8PcWFwu7QvaVbbN25/jtdLC2kDghKPEYb8dPXYgmxVF+
Kld4d33lMNXeWz6A+eboxmhUhgJq0aNaLH8mMpqX5TTxLA05hlGwClhgOK6x34Hy
nWCNKGHCmHmbAlYuNQS873i6GUcBuXbuj0IZJV1orwXC5YNQQmdyAID4d/2a5v6g
TAikZcHybPD45QoOCPSey8yX084p0RdufiT8rUSMOBtffyeFSjxoiKImkWUYk6SA
zWNUT1SJuzI+70ZgQbcyCBhqSMX7fE04iZkD5JIMhkjeN/GWWSAKqDsUISk6OK9X
JfdZh3z2PmXeNq7cpBzpzfIgd+7Wba+UzRrYLb5rm38NEB6dbILMzDVuQGo7cM15
KDmD9IOhMQCDxY24YGcOUl3vzluMF96Y2IsXB28eehrFPdwT+6erYdZElqfE0q+g
a9elHaKtQzmBfLECaLMHyGV0pEt984kh71JWbj4tozZKx5TUL8cGZBhHlk6czZm7
bBivQ3kBzX93fIdBjFH4YR7fAbJoAU9TPmCk+opMrdrJnuB7eixHRciNaPKmir/I
tDWFyOsmo1Vc46NJ9C7I0jfPK08/Kw3l00jeUdYmrY8wxESk9g8AWdHNobewRzpq
sV1x9eE6CDlOMmTK+1j2W0q0omTdNHSPPWjEl1nQEDF8jUQSnWwkBfKAuMMMeab2
bRJxNgW4mtQwd7nPKt00b/an/Q34q5gn1RB0dvAVTOx3KmxnNF2cGIC0JAk3p2nU
2z7mxuuXEhkbkfXbKzz6Jx7VTmMUsRzVphQwx2V+/xJfOVU3Exqm3ot5pQr70pjc
W6WNpe89uW3KgFryIaquKogUBKIRKcnErpfUpGHWFPQoQHu+HUIDCDiObuU16jD1
g7QY5eNkfPid49SH0D33lVk+0MJRQ910lLHuEf5BkgToxRfUwm+BfCh2WvE383kD
Gu5yDD3UuNNovT/W4DRW+7T92MbqSE35GNCGuh9v9zzPG9SLpbg09dT5nh9oxxAv
Qd9QJFigV1+Ft2hwfhyqpnYnaKvGfFraoi/Jg6AQPDr6O2Kz8x8HnrOXHK74Essl
PWR+oVCte7zzSwp9UyfLi4IZtBK+cjO8fLqWwANi2SSPQYSNxvURSQneTARCocCW
g5hNcWO17Af99xBudMdcTdPHHIIEzPraJPAyjwn3ssPW+FevsIP2p2rOPtMlKpZ2
+kZb7Gv7aHWiWhww0VSTe9nP/mjJXdsgBew5riM2gbiCc0ierurvqwMsZq4FbUav
2WqrYI/ACKBNp1iGM9LHLGGQXWeXkDQ+q26qm+RVTPNtEGmWtFItNGRUxeIKrWtv
pXc+6w9yelG5kMPGFlii/cXZePltu0RLWbRw32vzBjDd35Ai8Q3KmesVF60II3OM
qJbX5+jit9r1CPR/UxDBuLAYvWXtrHGYDfIey5vHy33rZdWF9eBD05x5wS6XOK36
ZtMDNDjc05UZRNd1cxZ+kCVom+Q7ZQ0XModpnJigU712noED/jSYovhfD7GsSOeC
YF+IKvjIFES2WcRtQCJRVJcxvM7YmKadst+1Mtw7UtrI1DXzg0wernfsskJ4z8nA
F18L7L9L5iWsPUbPzgYSHSfkXGdFMNrpmQWKwGgMI4IhGJd1iCUWHNF7hsJpPSYm
eduPiQ9E/D6fuEzam1f3YGBFnlt/d0PDQc3EjyBVclxv1UFKL6TLHq/KWxIgd0qx
DnoLnWfce3Dn3bgEiVf1Uu6QFZWmLSC4y41rAlWB8Uik92aP2YPNSYcfebE5h5fw
b4fz986MNUQRcpBdc1fgvGS4QZPsSK/LNps1rpfikqjNUD79pZ2QcA8ulnYb8V9b
yAcXXHTXa4QZmCko9jhgqzbDlBpIImQkj1c4Ibkz3wr6Jcm+u2YJ4Sm2eM9zCwoG
MEIxKtfS+L/GdXHbB80aO0JV7tTPe/yg8sJt7vEHpvHIJczgnBiU1+tXEyXvp9fP
Q/z7/u+Qr0PREZPcoCbfMRgcVcABcYsxScPuDn2QEkv9Rv2lYQk10jjClhYTswPm
S8TtjyUgbrKFNknDd8j2hVCS3RRy/FIQaR1T4NMwZ5Wjn0Ez/aDvIHYFNDUob899
gSkhZKJyy+k7kSAt/dOgKqU9Ccwj1ZR4PDe2TT7rU2sbDhu5S4hS4kcbjY7OfgVw
A/hLiWA7YDH6c6rBfnf84UJLE2BkJGReV3xQeyLR7TH24q4LFVnY/mxe5WZNMbgW
hcOgNinNShTosxLXeTa2zyHFvufhUMPM3IVyGwxFgm+I1n7OFKn2z7IDxpoiAD0r
PnOv15liQc9rHpX0/AgLxJfNQuDxZajdV4xp1U4GSOeX+1kJMMmI/fmu0FfrLTNC
9ZxbAYAYU0EJ+kA1spjdllyMFAjxLiW7uCLSLFuG1vyLm6YNkNqpvD9RisZNEjjz
ZdfqOvSoAjTkDSmh2UR2IjpQ83ynjsSyeiUwyO3JJde7+aTg0FNRGJcYXrNfGBB9
d0YKHBc7HQ5o+L/pXFfBGg42XCHm1kRwH0kW/Q1179mbP0t34LmmhMwMye0QyKS0
yrhwfsrvROcxTQfBugbCVgSg9Fm8/fU2VF4WF5yYp114Hs3JazyVhY9lFJ+TFI43
tcHxvMLPqnUWSIbmpNC4gmFnfnxwKl0Yd0Me9FjMw6x+f2I3dNxsm07c6bYqNXru
3UuiDlB/7rsWwgLUrgFl4F/LKT8JsI9efmTYWx3t0F1SnhtngEAByNoypL636r9s
FayHVDK6RqCIvyrKAzu/Z1MgVN5SgnOuDikWJii/DuYCyzX2Wk8K87E29sILALv1
zsNxdFZfLl/WoEDVBH9s1QKY5mB3Y+UX52SclnMfhee9PTlRV24joXIdDuh2uVIY
M0/nICMv8gu1/dpkqZdM0CtLFRpQRQXy9rbDJEnJ0JXtdDHxr4Vgm9QBf/Ost0Mj
abm/anCewl/SuZK5EmISsrdGE29xgqEafs2YzvXh7KOVlQVscHklj1z1oycOBhjl
FmaXi/61fjMjMpiWMTN8FdbgVXELS9Jx399HgBxumKfV4s+tO11OnzmnyJizt56T
9qZsSwnNtkD1uue9CW2yrGxMHcSH++cvONeoBBdRm4PkTKvbJ3NnqBvUP1j0Bzri
f/xVpmF1UycFUuTF1L3D+3kF58oFJUcxtIUD8cKnFBfSbmXJOxtiJCgEEi/o1+Ux
PxiZZ7Yk/FPVUJ85Mbop7CNJTc04KHOb+nJqIeoxTF+dOo4UvchfdkqaGaABqoOw
igLJLqjSmNZIojQTHF6pxw44hOp4P1LH8YaqwmtEzfwQEgtGKVt3LBVH+P7zmqle
uAJL5W1fWecPeJC4HawwyFo1VApsJ1G5LxI8PSeiyU3oESGOGzkteBbDtfonzSOx
nmlDf3Kns+YixCrKNYCOepsGDvgPF30zdUbsIqnaPZpiWcCx4M2wodN8OBgyTqEL
dNv11e7uCatWKjTWwXAyO9Ql8UyIXbf750Lh7UXx6cohkN8Zi4Pm8ubHdDhttv/Q
sohGxh+ad0uvfsU1gUZ6TUzCSE81Yj0dXIGOOxQX8RnJamqxgjdT5Hq02CG2rLqp
xhqdWl9AEkyMHHPUiaDDAQTbZmLpzOET4HrPTiAIunrqYdNVr81Glvzd7m/U18Nf
folg28s+btQdQPqCCALe8vRfX4HSDEFUUR0XUp8KZpIUxVoUCnppvgrayKVmRFmf
8piQHohGornu6cd1YsfdCSRfRg7BwXLS7nC5pEgwrsB9Cird2tfy3qZHypFNTb0B
1bNfR13MHotOPHmN2uZbBPA2xgztiEKAcEdSqrzQ9nqCF181xbCdAB6OTABi6SVk
AI+ZVRg9aPoOc/NyhkxARjwRpNW8xpyarkag04yQzFI8fUORqCUztxle8ssa57ZP
lq5IMPy7NNMG45cCkLfbdM0VRJplfgGdNIEGI6Y2Mawq2jfaV1nAOo7clO1nXTPO
szMD+AypIuIIAAM1LtL9sKYWc7bbq3ByRHZHqXu8D5G6DfRxxRwv8Au2Wtp63yIN
PCkJyqtyl8x3Vzj25yxjSc2qkCR8hmXp8PZzkQhW+8KXaUbPEzfE21OThZ99eVGw
eXszgSJAfO8rx6dc1CRPXcSRB01QjIiAELdpCopHdZNYjcZtdF1le+UQPANnYU/U
FLg9aP56BrzaQxkedqd2uZ5OiYOK0Uoq0pLbs6jfg+GW81dnQRcmLwekGGfHvSsZ
oIFGWsKIeVaF8jRowH8q2kw/tn+l2wqTBsWbDUVwKcqSrYeGt3Bqbv56ZOG1DwFc
ZR56q4bI6qyfEE5iSh8v0chOMpB6bfhY/u0V3/0MXJg9vhzIYX5ObrLPliaXDAAZ
iS1rwmh3QGphtswpaXNSRNAbpK5aQfSfvGfi5TmlQZUQfQw0LIH7lGmAH2SrI6vl
siXCLd7JSa5lx/92joZnYGt63UAXqX0WfFZMi2l4DLZSbIt+eLLAfihpkLDD1eAK
9kWSN5Parf0nUA80NH1VUe/wY3TYHwRVkoE9ZtY5qgG+TYZ0kkmXLg6U4Ery5m8b
VC/nScSXC5/PvblX6LbZqG0mD3gbLRUj8VgwRbEWqtlHgw1JVNXm9USemIz2VB0H
NuKr8mf0FgPf1SWlu7xVavciKdNg8p7x0c9keK1YJ2yCot6L5dJc8G7ACT4r7bED
DOEpTzLZUeOBpZEc85l/6JEy0YqDMemV1duc409lgKwY7XsjvV4zQcK49shLpQSh
+QEW90UDCHbaWbfnmIgVF8xylWBIbm2WSp/GXOu2Ghe3Roe7hz8lSHHgslwIeJDk
0YGLBUFnspsGLHQCLsdInSgm8cCXMsG5Xm0f72h22kJ2cDVFeK9CXS7ZOi9pJLVC
7HO2uk6GsWEkeb7sD1U9+EU8vC7/1Zfyo7//xTw/ogpPqwuvyAbSOfxJlZr6UXiw
o91p6O+2TCVlES9BnMushp1YK7XMhZvQlW1hMwZLsP/EW0C/7FdPz0jkmgqGKvPt
cocv0PD2oc2z9K271FXAjKDDd2/29oItsTIpXqJG7XOOWo9r2obR2HP787SMffAl
OVI8uvhcyqT5XPgjvre8ZF7lPf6fBV66HREzSL9PL68FUPyI6dQPGvkA6GWhYJ1z
GFULfu6IuUMbdxjSy0jAmTcjWHIucCoT80cCtU4r0z0AdfRHv8jdTPxVewZAWGMi
jRa3aXpHYGu1zDYub/UWvoIOkDnM6br5FKMKaxcemgc74HXQrzPWzDUlQ/e6f8GL
OaCRtY8qmT2Cr3R+Y+leGx+xeh/Boe2wkMt9sToIi5Zl4bAWql45hNIumG2cOwDu
ZpVcx7Rl4WonFc/6NKyw5QYJyesll1fAGSRvNYmZMlyMtXGx3r4cYZxFzpuOlCBd
XLmyeysK5KXvKAhBlOF3CW2+CVvirbEh6wWXXU4bu4aVHFTLIrPveYU7ECTshzJw
esUd0dolKgcuuaaP+5Cb2+QEQxFBaStac+VnpynM/F656mrUxsreAoCq01Cgf4n6
3WidWkUIqcXLKjYA7pzdXida9eEfK8gnnA0GJv9Nzua7FYK/D+NNaC9A12wzcGXf
q3BzhRCrLI6XUVpd7B4/XWxcL3IFusgMfbgBGp8z9Um5LHUA/xr9WPp/kgV/XGB5
7mAmkUVoCrGEcisn+8hno7BlyJsPlSGa5YCiXSxbOb4spx5rx0dVtQsSwJaazBdm
v9T1+1FdWRaz9zGlksRFnmdJFQmOhYYxjXTFTWoxBVysnLu+74BAdD+RufH+iexp
PpFFmXqmZOWID+e/JkaO9tDroDDeyvvMiKuT28oG6PFED1E9/96auaFIvIKXJJ6Z
/D4s69MSVHM/70fryOU8fYDIFhiiRwX2E9ZoMZmfw4/SmPVsDd57AUlSfCMaeABg
urmyHT06boGylADFD4ZnGulfR3Uggbra0r/7ba5roQU4hazu4IfB0vmqsKVojygI
hEybIOrRJb8zLa4sNu2kFLFnEJbvO4Wsv4NKtQeavLKwTSmS3TPVA9IXFKCIJajq
DitK5uqwEk1CxWvIgoI/VY25wgFwu8boaXTDLV62+APC3rqQ9skfqFDMYBwU6qJK
6h9RSaM5e4Q4B0oU/Zyn7E9ioIl9okxloN5tXydHYyADN2YzeVpY7lPPV1h8o3tU
lyL8TxEoHhbPo7OX1EnMcoICPGuMwSEuGDyLi5KlL+xh02GYoB9wiZmO4nj2MrwB
OxJGOJF8V6ET72AUOt541z2A13IMuJ4L4mvX44md5ARj2g6d5KnJgzFHnLvKngcI
JnOCuc8QOrcDIduL9uGk7EtE/db5uOvPuLreFceqXkDv3p9EDfOdmBiNVY2cUnMG
pGjM3MTYrE2mZo5LIf8CvPBdIT63UYn2I6BMWzkAF8AkEOd2CLZm6uYvF3BeJ97I
TDAvnLuaRvNJ+nnoehpC6/mphdpHVNwW+hhqGy46a1WllOa+LKnzXNIgCd+gElTJ
FrpKemKm9kweWNSn/L2DwK4MQFt4Qpguh8oMm26LgSKTChDjd8K23iyL/k3qbayd
YCQNqYGXItf3O5y6P4CZTEL0r+8lyqSElwKfCEeLYdQQpBmKhj6ZWvBVTR5SepdT
BXeUP8siUE3OgcK4h49jc3yxh9DHCF+WwDaEKTWok9ekTAHjlYrUJ4RYRx3uF2Me
UnhC/k9HEeID/+DcR4/rR65TakC0x5rPtV35mGmsBwhSS58J9zOG8sspVS7c3d2P
hEQlOTTMLARwTpJH5b+hW7eFSyJmg2hV8ERaots33acCccislJpkNW5bFxio2+Ul
w/oOBYwjZSr9z+AZ2ZS5YXFQrH5B0ujz374PwsGs9rU3A4mGDJaqSH77huy8c3lh
QFP8fSnEpfyCqypP0VPRuP4oriHtZVvyYRZTdAVNA3LTCWMlmzAqVAJp+9OeNzVc
uyatOk2sXtXaTSr0KyFUvo9HWuvxn/poVvfe7p7HHyS+jUxi7cdsLvlz4tgVCzJC
GfPtYofBp0zgkYlFBRF5Yt03Uo90g6EQlpOr+ztMNZxiyIVykiglLjApGffcN8lT
y32BSxjSiPRY7KeGqDzdaxJSYe3Ja4drq957Ap37YBe8yBsKL+KU/cXmIOqu98+M
8y134k2W2jiYLx9DA5ICWSg8TkJLop3f6insAY07IaYtPqHmA7a7Ech5DluKu3Nn
ybY7CNv3REiUWJjR7YAy6ar916V8IQB/5m3zW39CK0FK7jiUCJKVrpFUJn02Dd9A
eHo0ezbuCcb6JHmtFpoYWecKIFxJ7GXojTBZMn6tqdGAOJknSKfCmPKYn1v20HXt
SXnDmKv7Z6Zvd+KklsZHLuiDaqh2IhfZVikFC9OydxVxihF3HhqRz3czsa+hhe8D
dR4TOazL3D1RmyFPHnb733k5lzF9FkwLZ9b4uAwCT/m2UJJQ11SHi2manHVfXvS0
Bs7fSYHmK7jD1kiYLh+hOELUXSGCq3N4wJjLFiBXyp5YviAoBGvXN6AcBK4aXRgN
tKNIFAaZiI1EFT0lHlpudyJsOrIqQeR3vpnileDGRAO45B9m6gUx29SWurlW4bBk
q5/Kg1Z9ATWxtvHGknCiVzf/NC+d2APuU4JWiC7lYrol0Zp+CYlsZ5idtKoDz3rp
qZ+y1Z3ZlSLV5XcvDiLg8ThmB7VS8IkHs9Lo0kmpkEmKRpUdziqdfkORDeLquIfI
LV4o6FwxNyEgaa9ZpkK2zbkNlzyn9EhUan3K75kmMZnWwSuRruOiLhW8Qd3TzRc5
pPoFWP94Yq++UwrZbk8Fv03Mnc6PuFapOdURC2RHeAv12pNd+HQ1sLL6ESSL7MKI
9KhCxQR2U6IspTReTLaAg0OKgOtzvhgE8HXct4ty9yxWo4kZ5PUjiNQFTIuaqQTk
LUm7SbMkI1NrLhU5k5Vdg+SDps16Ww4+eBrc+mDyYomM3+8sGvZp5Jkrvsnq5khQ
BLZWJr0Q1LxSAIwCw2CWOsVxrxhJxd6Ng/ojdFkyBulEUSwx1P5GaWtswCksMbGh
OVcgNhUy4R42vYsRsFrsl9nu3VyNs4Qr2zN454aeOjObw2wt+2aZw9X4KDzMbP5z
5Pg0clOI07QPMCuiKbFuPm2lFgFFWIaQlq9irgCVTpgcmfgvR//FzumDJZ7jGOaA
gDjaKIvGPIKmICT+YJHGopqZNVeBw+9/Npuo1dYoeM2oCMQfl9rkTKsEz1bPdR/N
a8BKAnDRMNlwnzp0A/LMD/lQyVM0VVPPJYaCBUnzMlOD1NjvzfWBQvHDW3osAEYM
ThglN7Hq3U+Z93W6lacITyUlQbKbNBScvfbDBgdsHyAScEpbKYU48of7A98vwE22
Y9AFdyO11mrnzZ1RAf1MspQ+2DNOXQ6q7qsam8ThqaIEVQi3q/RMjVu0WOIfoVP5
ndxa7nB0SXQr4R0ifw3bKnY+mJFZRS07dXLodTcrGnJqaLYHO51QBQW+P1dCSi//
OoMcvMwlsByzJgro2gQaSSD9tXolXr+RERwd/Pj59OADWWtXmPrjkDDGK9vTEDVy
SX5a/YUaPJjUvuAS4JL4Ga2avUm4Utbpv2mRb4u9DiM3eEI8YeoLaui26Y1XWeBf
+VRN+FOwuthY9prkw1XlDZVPYOkGQ85jDlVkWBrkGz7KEvGYW6F6/ixRhzDKH+Ih
WePsexanHcGsKfCTQGZhfkngnXMlXi9I6U6lnpaieOx6wlwKL/0h0NQCjwVyZ7l5
4vWkg6O4dfewiyJoGXYn495Ke/ggqcBT0qmVuhbC5WTKAHh00WGVvFMBRktjmt8x
DNklDlglVFSNjz2h46DpXAtxLYe3e5ZQAocn+LIGb3SanPZOKDRCpP82yR7rlVYK
q4MAxbxUbe3kIXzXjyJSelMva8TWMq9vWsWUGSFzNS1RoMUBCHZy8tf4RreNOxH0
kCkXrwVHAselv60yKAX96O61l7eNV17DgglwKGmCCtAaOrnxmPIAGByQECVWNnOY
sOSAaYoc1h5c7OCDgPd+QyK2K68+u8ozqEvtkut2rvYIS2V5Xs2MJuDGGgpBGFfa
HN7jTwa31R/UQekOrGzbVHpMsnMGx9dvlTwiGmo3ByYC1UKwm7OTRPOKA84i13Ld
9cmXf4cttJUC1S0Wht01dqqN+wCdMDgcSrbcaFvwlepzTk/18bYtt7BttDdA93Ac
loZSS6zD+9bP2d30c9oB+CPlp4uL1dB+G2yuNRE0b/n3LXeEneeleBTRzAqhEt0h
1kciEG3PmRIUSr2Ujwh+U0C4GDkx6rfaPda+kC7VRBENESbXw7sUUfe8WFS4ciV2
s4g2omV0w3YDIcwUa7vrcAzO9PrFYYZ3JB+J8WS00RX13CMny+S2v5vd+D/0O8wu
kKqk2GMUm9Vg0IcgoTDH8OrneTT1sAIVdGuOkA+TI1tyzyAlmQodhb8V1kUN93lr
/XSkKg0/F5OVzu0OJPPO9i/R8BtLLRNNk3NzCI8DsPaIJoGJTugQ3r9/o11NmMKY
xshWZzlrBcyQmM2J9FXjvGcIW7dDx0pRPIqtCVfzGQoL3AX7hdfqq5IQgMg8i/4o
Aox3S+k2zSZPVm8qbxmKH4VOjd8KvEjYhpTpmH3uB7juTI2rrU9edaBCQxL5+g2A
DUYOGAO1sKdlP3HmzrjmmFZvXVst66LdK1do0EnznUt0fldUUbYORWzRizQuK+9u
vTl7BHPvGl5Wk8QziP3Llr+QTcXjJKn4iBAnuiQkvGmsG0JG3tyFJ/jFUyQYSfbY
TPL6rzXs4gfxx20+vv7C5y9/miMNDS0x2CDKOfGVFig78yHuDzneHJXDZXTzAdis
CGwqKr5rFwOpScdwzWzoZgmgibPKxuLfHFRuZmpl/PTHAsPHJsk2JwVKblxzETxa
9uZ+wAwZf2vnC+L7cyp1jaCO1blVSErfff+oENnolR8bNsBVf0pPV4FTG3nMYzIS
wNAtoXTVRNqCFe6C0NLJ6OW39BOIRK3jcHGymHNMAnlOVY2eHfnuO77QE/OSTiK5
oh4NLIvapY/W6CY2oueJq4wGpACJONr4rTzoI2LT/4GJS7Uw34boP0tcgaBJRhc4
XgvytS/DRGXJ7K4pjlz9nALBx7mdlnFumFeIzy0ZQCpw0X/9uKagOQgcbBBmhIta
VERE01LjYuOgXn2+hc+VRDK9s5cZeiGTIcHJmCrK/1CaV2GhJCaqP1Ut7YwkSKYp
YKDQr63gzmdzOo/WZFnDj2Y9Sgs5ztcrUx2SwJuDQD+uOzq1blaEokKTt86w27qO
78TeGvAW+nS1bihtlBM8IIJ9+msnMiaa+DdgvrlE6v/aUuMzeDWeMCnuTpH4I4u7
quD01zw2rb4MAtmq1q9EJBMfCeDohZ4SMjP2ksFz1sMFeIXiddV7urEdWTh4T38x
ZS/rg0WY2+MymLe9VItT85oIsV06Ev3lunikQzEzZkMlYO61O/lmLArl+Ut2Kvu/
ikkKs7AN+G5cVNlulA4yhr3ZH2kabKfn6WhMSIdPvX187t9MFvaCfvoXsxsnyvfP
KKwyWvBXTWvEjI9gzsbRCth980n6/wRFdIiHKwrg4w2PKlyxC45Ock2K2Umlze/I
kxUpjVlEn3IHe574YhOBcE/rRyn77JBu3CK5T/eNKfbtMQA0CIUnEtkbx2pDgtf2
SOi5VBAaxEDRyRcLfgq0Lnr5wUiws08SccotkLusdqUqV8iBdFoVOtZxpvRqSDOs
FiGnWS2vi4iAhNFTnweiKrnZekPVenfU49d12pxc0dkf5JBsonL2AeAvebrOXLeF
K8KZfC9QATenyLNuZb+I8/mN4d/lHTsREZM3FA52BkWJp9fljsgWg2zH3x9rmqlG
3N+xKoZlI+MWFYp7iQbHJ9HmIa675gAXMZtO9PM1eYGlPW3RN8sz16jOgrDzk34q
Y4zQizQF4uDTE3Vu/t0Z8cHBxsG07wCD8IKNfk/v8OJjL0raOqCTtiPX0/Bld+up
OR5YPAKzNzXPcjPlg1k+OHQigK8fGrn8Y+mYtCVZhJz7KlHuQ9gPZmkTCcDanpm2
C3I2pt60yAaOQfsQix4JkKek90cpwh1lN55AFTXeYH/cn14oM07vTK8RbPsfG4xi
Bsu550aQREbPOpGakkFbC5sp6WuovcZRsJSO0jcCJWmnDmSPkJI7v2NOFBcnOtrt
Y8RrK4zZEx9R+Jb8G8AXZ3jm3W57/aDRBHa0Qr7nbAigZetFgva3MQ5OaD81Q3dp
l5OWWu7ps6nN0lpTENmkr59oB0fii8eWHX2TDoCqSgBQ2wmwGNWvZExA8E96cl1h
EfxyrghvMqbNTucJHJUVdqUDLGgTUXeueFn2HdqKPdMi3Py570Nv3pB0oBXQpfyt
Nmd+NgElOabvVLpnvipddQkd5OzvHQH75s+fGgi6pvu+sjtiv36hACg1UtNGZ3zr
B/BsHQZqbspJS+HFn2PK37WzPE+AxKYPujdhNlBkBfBU6cUsg/A7Vx0gbawWjBy1
mHQNvwrgXb55O2qlKEXKqzfqWcc2npuFfXt9154Kcq4Uqf1sK39vxdoOvaUg+QJM
qhIi/jNK/2vIf2t3Z5R8r7GT+YBalQT5VP6UR+pvgfNqXog5vIFXb/pwr+sVacsE
eZkg1wVAmg1cr6K0WIIcY7RafSrqwRkAGxCMPF+tteOEGBn3qIBxobUWrjGHkDcO
LZCV0+2z83UCq9X+29MqLTwNA4zsnsJPDL3SShBe9XK2o17DVdPuXy3Z19j9GFOA
8T65L2yx352XirF6m9YUgRCALXXPwbVkpQXTgJ0j10cgjMedhIgKbZcfsYIRk2HE
AQmHnD2IMWUFLIf4Y02r26JGNkW/DZ5ItUYBBgm5MQcbPndRP/sFBYMJu6d7k+pU
rHAthGnoCRLW1wUQss1uyyQuF8MS0jzdKXToy60siguDQTAs3NA6zW9rX0Zr2x7M
kZITECafCiY/70kTtUt+xVbEjuLYWvk0anwP25KjT86P6gsr3dx5gIo7C8WtkZ5j
h9Sp9n60WdHkVWEoEPe36II3QQ1m4h0JuZR4WvG03O183uC6ggH0v/GF4Q2UpOmb
tpfafDJD0tsm2CoLyF9w0mk77+l4sNF8K4+UfwGNSWWLBqp3A5Z3daJumx0yIye1
Su2XR9t8d1VoYpNxV7SLbQi2r7RFJcvAOIVsQ4qq5y5NCtBfbor8HnMmRUMJxcOO
lpHGZKeAUKnOZ8WdSHzovrwfPb4R4RLLvrUvawPpIjM4nnzOw7NSgxiQ9ff9VvD/
z2ypoEdTQT40OnTGp2SMpIjq8nnD3GeX5ZfKYhHQpWYBtNcW4vLvtH6kpuxl6nKw
jrmeNqLnuQp0Knipd5kkFRpk4tTij73K3x8TUy17Ct184/DQwrkJwdPiB9Cnao+K
ubUd0hc0jRnw57X5RAZYrKizgBN9RB226ggVWfhxh6RByy14dpqIz6ZYmUBRmcEg
RZfbii12ZQKbOQhpjLT1qt+Uv6ckWrr53nHeSbHbVheHzKy7O3gf/3pkmA1NFfZM
CTFr3UsqgSTBwNjFKsLgXU/baz9MzsJL9Jqo9HpdLxZaCkwwuluv8Arz4B7L5T04
8ktG0qYSA5S5bIcHOEFkI4JhgwrqN19jqrg7vuPehnOXo99UhN6SrzGGkBsbZ98f
7Udi+tN7Lp2iasnP8Ky2Rvt63kV3FFBgVjdn48vQU+sVZAT9+QZoKqcPqeFZbuz6
+h2tzwuqE6UCCEjEElqSPDihZ54DXsb04Qwd+dEg9O/+QpwM9Y/DFpJf+sOgKbCn
SySo4SZipryciUkvNrdfwPM90Nx7yxkZcJTlomQ077M1c26Y3uUXtdFw0Ve3mYhT
bVH/nQc1ZhpK/NLC3Kr/bHioEhOv1NwDuPhUqYc59kwWDJc6xtOCE0lIU6ZoJ+Bg
QX5NjtAZWpCNUOivEyjjbkYgkyYVhWdN7hCdSQfRtoPuVdNXUzq+VIYKvFNOhL5K
JPqLrLGHgDLzSsWCmQ0vY7nUztnEqcsa4xzN8NIH+xLY9+8CEZv0s/MfzmSydHVb
1qg5NfywrWTxOOhA4F1JDILCC7uyTeg6I+SnbYjYnwLRdh0kzyQGMeSiMNe6VKgB
HAeUDz55xqd6orKGNmOJ2HIzvISlBS6IkkmwzHRwT75PKG/sHgvPqmFL2nIfpKE+
Ezbl5DNYSAc0VS8IWeHltuFZD6CWHbvFDH/AlmZYj3uEeDRf+YDbCdquowd0PUlb
iHVux7geQu9Z7KPR38yxnq5ZBfLbmhXo9dEm8Le+PNKgnUd7RsyOR1w5ljfszY8h
MraYhlFfihw8sb6yQ4bhHeE9NgNVpNxZ912FaU3QVn/jeSaxM4dbL9FJ0soHBQHY
P56+4ruk8XrVsKawj4erKTRhYQDbiIM2GcwNPpMN6Z6yXl6VE3e9JbyyIK3seOFt
LDI/V68vDilMBtw2dsdfxgSHDv8/sXmLOGOpt8ZtrufVDFj4ON/EgQAJBqyxQ2ye
fdD78y9W1mmc+QzKIMTYe1o07bbZppppFIZM7LB0rWOl9/fTciObOsmQgXHwhftM
DlnTptQ8IhQ1Hl2eucSxYzDq76WaiRJEgyAycCUMh38oBcO++sGwvxjMth9bkSVn
daYeNwSFgIu5yxNVE4DuD6AIaaZLnM5yPfzKOW+AIE7E5ADQ4SA46j7wGIZwXI8I
PEsl+EtHltITWq4XXj+G1Xabl+/4BJgJCR/uGFi5t0rZPvVPUQcFCE1xWNUapjod
wujWnPJJA9y1Uw0tXv3zZHBs0lUZov6CaguZiR+sOVBLRrcHNk+Klp31iPIRQDng
gkZrP80jutuA6o9RZcXImHJSk+eTtg+A2zO6hTFnVJEwmT8bjzaPhMYPJrD2T7jA
3vA/K5wuehmELe0AHErWLgvS0x9+Q68+0Hi8AbRmyS1EZe1Cdah0zy4ZFEBcPbwI
QQ863NEp0v8gAD5/eI01/2Vw5s/3/u5a6VjR+KBOo3nZL5/lbnFRDMIU8Up0sDig
YJzgFRVU8M4o5JFS21JwM2HAQupzu6et431BKlP4oM+kGYM8xcs/KwW+G1wjRVYz
qhP8eOjP/7SHL58tWgvpps+pifIQr029fmNlu4FCpJ+l66b12GO4fYmFSdr5Qn/z
N30yc9DvTjXQq4/fAHWWqpeYdWx/4ezpQo1hbaldpPP3EMXm8Ohv+HqhqMlLfqOK
2ge6jG//h16wnbJFjfj+lPMsNNoX6YjNtr5yGuPQX4wgp8mqkz0nItMSsQeU456t
sXayrOaPAUDQlZlJf/ROb0j6p0BDb3Gpd8yszxeqamPhFn01852i+PPwNZ80c62E
I94pW8d3zahf0puukH5Q1MESMTfmANZEppJfuWHjSFPLdno1f53rPAC083dTfjRA
fN14MuUe4DPizdNwDCC3FpdP+0QfJgiLjcmS1A2R5nBcCLr+h9l/ZChXrKpnyQ75
fRExhHDwK+KbU6SlEsWVR9R5+HrFxKNQXuMB3yy03A79ghnQVA3cKf3PAUiocPEp
nEcM2aaf4+dX3nTscREzGYe5angGIT77E3nHFzOLJWFBs/2fNpHX3sto60YyrQ4h
zDCM05YvAOg2HZ7ybZtK59V8+7cIZq8EMENloKO3yLWWil1J5GmjOg+2vLjMcI2h
+twSNEau0+OGkSzBlMpz8IRVIYxt0Xb3DsIpVjApIcAuGUbrtlqJaOe4lC6UFtQ7
Su+zV0J0lpmscGxpNPyi5S55ceBEKs0lHNjWYvUG3VT18ADFW4i4jLKyCgiWBzXR
yJRIavoj6q8o6dw52yEhcu7Iof/lTytj1l47oKrMbQVUgS1/MC976PNPjvHMY0xt
pYav2CL/ON/SlujV42+V6JqPXHDBX05mbcSBxDMfqhEUMADbDS3E0I6vIP2T3zfQ
ejbarb0lZOSas/Kqxt48WoPvgUT9b4mhDroXRiN92DUkDcz5/lAoMyyYHGAOCyPz
unKruXwjT3SM6YYJAJaP6ZvgTJ19l5Edv8xBr+mpFKlKv4Or70m2QCpkutk+QRLo
YNoCtkocpHvZNzHURAq+M8OFyFNOTor6Nire+x/KwIc1eEaJbTN0niAmJBo2H3JO
0BYob2jwcNBRz57SsBTGnYRGL+FAFzf7HcxuUWAY16YaJW349bsCy78M4q7XLpC4
Sp2H0cBTnRUFXD9OO1AOXs/YIf02Dx1ryCIWc7TfSAxCUrh2xJM4jP63qRT9ckgq
iXswj37Sv01+0VeahdbNb60Dl1uQT+VW4hTRbOdyqNXL0jhYQizEv8So8RdBBL07
pfFj/g2lFSsEymLpqVn598n48tGbK8uV1XeFWCWUgGzITA5aEVxW52s0frKCt2WN
mrMEulrFfZpSJnCMWFbhFfA7oDV1ZEXOyTqm9gQWJAZPaDqpbXsgMMk5GJRIMosr
BU7VhbXxZp+JGbt7Vh4kmP6rHS/ba+uYeiAkxlm2Sjd3LQHLEyC2SXCF63bm3p2m
DT3swEjj4CmF/AZdkbWR9+F/pch9PeDJFajq1ZQ/j43BH2cctrdTRkD3ExMxXegN
MnCHgD2ZRB3i0rRZ3QPxhXj+PQsl9hFpwPt3qh0JRP9tgjR5IIsFcSb8KMvFpeTh
+5dur/Z4/fHMg9N0K5eu20vEnTh3RXDRXUzmTr9S4thLY7zfjpW417EQwHSnbdYx
xpvk81AW53jzOPDxul34ajlFXpfHwtBL8l54mvj5sZv5KsfSf1GxZOyslAuL6vT/
WxokLc+IHNdpRI3YuZg+xYtwAeZHgD2+vsuVexvwPw9+GR2z+K8Uumuzm0X8LfaG
yybDKPaBFwGKcHw+QyKnjqtwzKcNtYOKkxxyEmeIcW6K/zjQj/J9AapdQwlHNonc
vcL6r36JD9NPJYmBy1/vNdO0dXQD8dLLT9Hq+G42oAnIB0W82DTnEXbgWpfWrYwp
8WuaIHLOd5uKJGMIYhxbr06udWGB5trKscUcK4AtAT/xvbVNDNEvbAobhKhS43J8
gYImEq9pX6OUzIWmPScB7f1+YLis3phvsWb5/BgIOC1zKB1FysUOKigFzIrNPcKl
Aqp6gU7im1FXDDogHXgXzgBAIcOzWP+r5Bxs1uslfsX4mms+QtmXlaB3uYBCAKQ5
CVn1WiBjTWVwurgTlpuYuQPMTyYk+Lr7wa9Rktm1XpR0vT+cCUqR9a97YBXn1rKg
tKIawUN5PA7kNAmfWUfpAjgSv2ytdzuXgZk5+fMZI4pUmR7f8NVGBIyeSt91YG9e
ZpMi9wwSjtkJfhjr8YdHavwz7sOqSqn5feNhEuwzF/UWGi/3Er277KlkSsJavUpN
1EG+Nl1+r89MDqqLyEfvvOLEI6/XknbVWAC4S2yqf0cV7mhzJw2QgW+VzgH1tAKe
y4WYjc6GGSWQQTbcn0o5MPoLGK3HVghSOS1VWOMvcMDRL4wsdQ4bnK7dSt32poIu
1mE/I0h0/g5pKGTDdvUMvOe0/uCau0pNHSrsOokkmSpG10ugInzLyd/yjMP0Gufi
2LKs/SLpwtIhIlxOfbqxh+RVUmSXstwwXKg5STeCvQ+pads07oR8MNAG1HZzmRLB
VxYEIvRn2UdNTHnfr58FV8nKY/Ly9NaLf+vqZ+3ApxK0CnZ0f15CzsDpvl2rjpDj
iKwGLVUzuEl1iYe3BEY7kwHYEJbgU3h24snqPXoWQLsv9eERdgwVi5gDtiwvokRO
75iu5pyYn3w4BXBi9nvZRj+hstm3EDcOAKeXAtBGA/jzzyUCIbaKsZCD158wXzd8
LPFyIMgTXj41zn5WZnSyumTEJK5F8e+B3R5wB34oX47LJ6KFi20QZi/Qt117gol3
/uFuxbRm8q2vU3RCdC2/n4AaUVHW/1YX3vaJvitouDkehYAzFrxmA27H7JDmuzxy
0OJNW7dSHOGX1STlSL4opDKD1QasnqLtqCYcKC2x7FDvsPD65t4hfh795MQvMJuJ
pa7BfUIO0fujt2u6c42u+fE32P9EXeTJSViDfd7scC/lXToW6zuLBvm5Vkvshalb
/c5MjNvV+IwprV6l5PkmpWhuic1tRA61RZjKiK/ogs5uGUFqh4wEN1+v+sOt0OCM
7ZN9ID2DZw2oTPJ51fz7TJ3NZUsfKW2N7jIbWVDMIwmLz9x7VMxpcSFbe/QY4iSp
EFKK7MSXJ/5weGBGIFvWaEAGU/IVLX3HCNKmD76OzirsLos5peFYmiIERRlG0Gve
XP4nR7iBTLzA/mKhtVZLt/WYqDWxTrZcJMP8XdFhhSU2088ccKQ0F7/3aZNJVdB2
gD0pCvkPP1Syi49xHylH7lwm67aQ/iPqxQBEZS3X6t/SdDsvYI8gWJJ/qrn9D36z
m0y+RgZZV9ArKBbp/h4wLhn9IziGQIUzjDoQ+OF9MNVV4HA2tPcCAA6V+EZ9Ws/M
HbO032DBHkLsDpWIzu+xW8EKiMAwy55Omj619S0i2CFv5I1m1pDbsnkk3929PcMw
rj/IIzROXAtQ0nqZ6flLhbnznoUoLWAmJougLDNe38AivrjpahM+4KFmXYfNVyIm
+18C3ZkA8RsuO3G3zXuQ9GJIo8Pi9zCK/HokY4tAogjbUCNio81+1kyNm8jZUoDV
X72bn/v5dDcYs7RoYdPBD8oZwYSyOnOkFAQO7SkfdZ1hDr01cqoE6C53OabV+MLD
cJhqKkxabSgsoNkRx4SBrZ+pzGGI2Hbn6qeqqHwdrPGd5n+AuygIaqIIcrQatG94
FB6kI16qPrIhRSC4jP670LK0cNZDoZHDimsYebeGY1FSAVNs4onn/UkM0MWC51xz
aK9jggqFXUnMqI77ZcnFd9u7i7NeDFUMkX8IiQc9hfqDRiV9zPtBN46gjnIpTLjY
6+saKYw3qSJKJ3Jtgr6jJhZfc1Dj47WnqbfDqxOslXuiDF7Q/4Hr5fSNKAJZyzCZ
beFIsp5sJokju/pxMkNlF6mn4N3PrrxZwxYmQEbdw2ZYJqFm0FaKg91gqU9bdxd9
jOYE4w5fWjpPwKmlwO4CHj69lFzMptwpslbMPntzlCjIj3N4uj7lYnC7BbaFpDPt
3rXTcG9Lm2nyMtNmz7wd8MSC2XKkKoRfc3lmyd38DGTQaOiGBrlUaIVLaLj91W57
G3k8ieAXcfUkrox7gTy7XtxUQ+5q8GNrkpssszvY0oaKIQcEbb9N16V8LQyOhDTY
5UxCbId2L/UcKN91LORYgxszcSOxUhqcZ/mFUd7nk0LPTDg/xRFO+0abP13Wp5k5
B7vqgv2Tb1OwCKixD6kGURbaiad7PN3M9TGpCNsmvcLK4OcJk7a/r7uwbT2/6mfR
gCMVMAlK41U5wDDddvWc26aevdWc2SrX1nZ/bkWZQHJ/I1lkFHQZfJPDwJUth3wi
2QXHqyIwrpPD9HaiHkLJrk5sNmVuNEu2fLVOnkF5jS502KfIHGYxaPMAAGEsbi82
TSsjsfedyZ4JeeiOng3ztr7NLb9xnKbmh0FdwH021B41E6EReprEc1whvjfb8l91
yavDGTLOTXoCke7fqCkkHpPof8iWDAcewUILfm1gBwXNwOB9kATMjamyUxLWOkKB
pBbOU4Dpm+Ugvj4D6JtZUJ/v7L4+OAUDMC7bz6CunKQw97XlsqDzE3+VdaIuIJzs
6yWE9mRm4HnJtm2vr0ePAcEpqYYzxmrs5W3P073XF/krzV2CKHPXtkUPIhdZiyi5
WlbX55RJLoysJWbEWIDCyQt0fnw0VpGYCQv6iPWICX1ZttlXkU8mKJhzr/MuJWiB
CbjfIY9LwZi5O1gTQBKJp5f0bOYQliSD3Se7h2zZu3KoZptUsEDFr5MOr3VbnTgJ
Yg05lerY8WonP3ZUyOiynuecMq1lGecKUw119lxCbPj1CFCGnclno4v9fruXIfYX
egJErTJ5zGGzl5ZD4rx6AHzTX6ZVRcXj0GTI84fYUPbFYBqq8oW+Ado550kk4zde
QiT0iA9abiAD+K3MGZCuvuAk/DfbEqCV90qHKZQaON0YxIwi11dBXnFznboscVwK
7qVHy+64feAZ1nsqokL/24ikX+oR3ZcfJKr757RQw8lRXuA0JDGw/FI02ZW4TSGq
ux0TIoa+Xniwk6MglsxgBi9jdJph06MRZqu2sq434NXSBggUe2VvGlz7JsLXouUn
iYR9hPm7lJ6IcmWoKVoSQTxCJgpSIPf/O/7ZQX8deOzRFqweaojxYm9U9gFgQ9t5
CT99kS0E6xGlV2bqKGosqeJ2cf2GzMfrLjojO3fpSG5yR5ScGpJjJx+Rz8wrN3I0
sK/umLPCci6Yb8GKQ/GBd4fnwcoxI9SfJ6Ce8zJ77FHNiPNsJGBy1O1N11P7sNf9
DjxjZxPhLGozigIawdXM43uCQS8f4CrJN2GSyZ7mEkAi/okfTZvQ2yxPaqiG/GMA
UZ6M6PDGYlldn3bRz606Ny329A6Pk0AC9NyWmBn2WjRELxl00dingbfhgWj5MPPP
jveaL5uLVhbR/ENA+V8HPbKz8i4h6153IX6qlVjXdYAPVlDsKnfYhU2rQ6Ozf008
tcKRbel0IvD5yndhig50ODiB+yMGJwgw3RRFViHz/d+B4WmV8q18MAUK8uNZGJvz
m1znIdfwYGacryW7nx86EnWZcIYy0b1TyhspVXk+q7edznF4FHBD6gt3En/3cTEM
FdT4Wzbuj9A3pgIfqP16Q8iPVjWCEhvSpEe8OIlTz5x4U99LZ5EdA8xPeSDdM+BG
ExNmw+X6i2MrJy1wwf6QTQSC4pFe3ptnPFMe7QuwsTMpJkyYmcHKfS1d+XYZn3n1
7CDiKd7BEX27/owoSqWQNiTIaBnEdVDuTecBS2NdZi8HXdXGj5bql5ZCzGUslV9o
uMQttHOAXq/Q4J8vG0CNuMyzD0QarJBVkRdwiVYuz9xp87CnwD/sXlcTYJQ5JCT+
8Wd7AUVmoM/NAqFjQMLJW83vSdK2I3eoQH1AlVwyl4dMDzucRYJOeqMFylEB8EGS
Isp5v1cJmNl9U9ubJLQo78A6TqM3JBBWf3B5cKhAb68n9Pt+vm3A3wP7Dc+AtjnD
h0PFa1Wbn4unyHOyq7xKNpzY8vwlV/lwGSQLo2NYDlgGGt946QB74msGhOPGieBv
Ub3KmKTb3m3iBOCPtxTEGfLyDHmR3K7GV9N22AwhiDGAViysI6VKKdbtuNHJd4BS
t711E/jVQ8QTTK4gx+0Z31Q1tV7kxVLSFWXtVJKFsHiStsCf0+V1AdqAZXTfyMBz
oMbikKdJje/3e9FlH3SqQUg0fAIY241GalcoHYcM6BuOXXmlg4wPE6h20HTSNBTs
d2paUWwqheuzs1IRsx5hsPuDhjxA6wS0SWomL0j5OK4tIK80ofwnt/0wuO5PeohV
7hKpVqkfFlb/copfCh6F0DAeiwXoUd/lUa9tfDHQTaDMZHtrhBQuGdwoa7JkKIrD
EGy9R6tiwYfDZX41N4Avl1h4Vz0zw61BYuUVrCconmLin8NZr+6ndWwLXPaNqhg9
SxxoxnDtpVxhhgp7HV4F/LmqLGmNcq+kaxOzSx7D2xQsJgDLM2Fvt789pB6USw1J
S+KIGISAkzv5y2eUzLfPsnXaenLBY1tHf3hyV5rGb6YmR+ntXeihrvi5UJMwl+SD
BJsyobqMpxtsM2YbQ+19SRwMwosKwO5Ln44yVGLnWJaPa35CqkSZSIwdhRq+Ojh7
d0kc/YqrSH5TVvDg/mOE+Yz25IEGJI1SQh/uG6U6/0AUpBmIvhnee+yUs6oXbnyu
Vefc/TRl4xczXx7tZPzARSXObIqjnZJw1Ui5JFI0n3ExkkDHDaXGTsmw526zp4y7
anQ/2rIVNGt9OaZLTJ5NgB0SbRdgeasqiBgA8KObEwZQ4FpGHZjjJFwlF2zwEklT
bScMHNHO5MjzqRtvRzI5YM+dvMBFk8Rkct77EDOk67bFr7NL64IQS/rW42J+jfXt
Gur69OLOIDp5SRzYMp+bhCvDfelltqFdJ+1VDEkWy7io+1AgTAkQW6rUfP3XVDr8
X6TJ77R9ATGrxclEiyHP1jdN2bxf+6a2EBj7cMvJbUU+jWaisz0QRGCNq32XmHKV
4ulPyKqGP1SR3wAnQ0TxwlvMtkja31FBxz8b9OVIb9YrHYq6uIrR0Jotp/tRb52p
viUyQmBhC4r8s27AL9h0D8bhetrNfuPYwj+fMT/TjSS1iusdjPpnapXcHVXQkaZy
DfMrPU8AtDsJ4XKFF4j09MFNG1fLBfXfOQg0RxuLbBKBGA6IshIEtYRcaSR8RETY
B6LxiYDkbWRE78fi5DrKYBu0GqMvEao8bqPumUboJtMRcO1YkUO21Yo4Ojg4hYBR
1JEZoc9PBhogoTT660cbSZYCrs4ln29IZCsICj/3H+H9rneO+VEB6Mw1m4DhDVKG
R4psYFCfp5cBnxDIZ82PV8LJ/kgoVCQUXuq3bUMyX7D3nIi3GvIQMkTvi+p2CHdr
6EwxTuGw+BQ1vEdnLJrkk2nbllao8fsR0StGRCDPh+5iDgQpLI29vfmZUUloA/uL
DXFxRkrKayU7dhbtDZ9gEvqVcTYA2uoCnlfDKa/XL1v7n0VTaE8kNSLg8pPx5K2S
X+GIu8dFk1vQQnwzN/dtmhSEb7ayTuSrdj9Ngbgz0Vxg5j1AVrQK9qXSasFKPfVF
kDjKYiXtQ22Y8VZ/6Ep5Ik/AhnWXwIARu2TSii4VecNNbExWlXfr6CNAWDExwyDM
yYgQvG2FOGHyqniY5bP4au37+hgI1FBJMirpRmXDPI/SuS1W31PMvxFgMB2A2msM
A0m08qmUD5TzBiDZxWk9qN5WmhYDd6izXxmMN0iJ5hTvExNIlupXYlo6dgu+l2a3
WPEHHsm3MDX+7FU3RZO9iScEObHZGsiajleMIM0U4V1WmCI4lxth5sQChQoxlBjL
VspkTRWk2sL0Xs/RdkeOMx/7KUaVOYU2AOrtpTdl25EEqMsBqlaHaNrkcpgK42XB
ZAWUw5vNNqD9CfbTXpnjO4RKq1NbC2jDhTx3L7Ho2iJgfcF8Q/+eQel4QkLENigV
lH4uZl7/LFGiU/Y+Pgm6G7Ew0TYyfb3vsSn1OwApahl864Tgt2RRlFk8PCRakzx7
AAgOuK35OPYayYvlzQAUnGn3qe1L/TPiXrNei6tQ3YXOe4+bcOFcioLGRSJckQCx
QpoWI84oxVwoZebye33fofbMPkpuaBcr3TtXwF8KiZQV0DnTrwLjpfE4snrWiiOK
nbrNxYfB3CVpwD5dyzIiFINXpQDHNBzkykudDvm0IghSmZp9Wr3fLJ1j0vm41okA
BqsNQJgolRS8G8qBfy7PTUbPX4NIW+NIpLl+rEpRWbY6oonpVSnXf03u6EdKi1NZ
RrF2s4f9jNz7lnT041lKHtR9tbkhEUlniZ8JV/JJr316lKpyhpvACIGWHUAmlwoj
GK8pqjmdopFp9yorXnomEkbXaoqJzeZ0Hr0L9Ix4syfI72+i7YFvK/u+a9xkRqiW
FIWwjKQPqJTpwDmJ3FqBMIBePXQK6bplS+4NI0LU9Qd61bz5Ahyo0MxYOZFR4dHI
QVSFngKQIwmF6n9aLeRhN6Lboh4WEjAD9K/4A4oo/Er6oRsOzoxeBcOlKgDx/bmE
BQbmFbut94B618su/Rttba0YfIfr5lNWd4iUvxPiRfcSRTaDqNTJh0+vjy4aZh+T
5Z6khsOn1DRhNGBIE7mukxcH3xt/dsZruQV/mtRYhW5hygTtjqmBLID9+Tr97IBL
IWgBH837Wng93LP+mwYa0+2tsbfByXuZM6v4DWusXL95HSJksKaPNEL3Ies9791R
eNuplejn2+qGT2f3OfHg7V69+kq9euZ8DB8neFY7ypIwyy5FPB0d+9SuLazUMUgk
CeItGDyBv9GukYgybJIIdsgAWGf6j2ldroFIJ6xcVWx/sr+VKh6DwmWSYFyqIdWX
dj9TFZV9jmUlsUxq8ufzit00a9JmHWsWJw/6kM7dRzCzoywhxsJR1CBz9gv962om
MCbmh/doySG4w2PglikF6cluLpQ64+hJTL8MLfVTX0qeeFb+QOSS6QdbxaynvLKz
zIhAGt3TTEycM3YPqDdGGcz8wGiNI+PmFhA5WYbGljPRGVHJAKXF0C10bbN6/VDF
VL1gV5u2Rka+kDqxcE5Z7IMQPnIBgrX+86cogddURbuDb9diIbwB9SwKn9jiG+v3
Zb4RSOUZe2IZqRSK2jFlhTYHRf+2XznIx2+yCQ4VNrYl9pioOXPOcPnSMtLk2KwD
MODUUkTHDPn13G0yiPo+xDurN2kaJYB0rWZoqni2WXp3qqr2Ffm0GIGjGPTM3Y5P
EdGr/HDnsv/2H8oq8QzZ/RXJn3HQfUF+gs8t8sO7EKNYQZrVjJ8FQ8PA691NXvox
pF1tj7gai5A1fAmLH79idTw2pNP37QkM0Lf8cUwjwW/5aK6FR78a5ozNKUfScxq7
g/fWDZlgcGfWSNq4bzXw5vy84IgKXZV/v8FBQj7s0cB9BUxOVGfbcQRTROP2g6hg
1ytTTRI7fAK/PUP/iNQuOQUKiPU/87QzhL2GbJBjTATd9Xkqy/eBcoKM3qs6akxZ
2lRQ2Fu6CtkcIMOp9H0O6DxxpPkCneUfOES4oKDzHGBBHAavL0TISNTUcyYHQqoU
V+VuG53kTNeHTcQNts40eCrbRGgdCvHTt37yT56TNtdIEDe1Lqwq45wI3TN4V7qg
M/s1T0qan9Wmv8+ohxs4IisBx8LxBAaP/iHyDeCQLz8ipAdiBoEQ7PGrJ4qOGr7C
f2MeDaPctDnKqDZ9DCZOX5Y9ZtEIiJINhCeo5wfq+m9IUXmNI9s83RXII2V3IVme
dZVtyLyoCSrjhWUSEytn322iK5uerZLsN0sV4RCLEtIYobHBBKo3PFcvffoXTF4z
fIkDVTNxjjNLQTibu5CDRNFgnPaN68m8UNfJcnQhkb+xaoL4CmEJiaQahIZpJ4x3
z889pJXoe5ORmt4L6kUxFH1Ms+YHpWb0BKQn0fGGfb6N8wFP98WTyYyVu3UnXyyY
jnHU8+3nL+fWO95uE69WQla/Iwxiv73LoriFeJbCu/W6WI5aeFAgHnliinYbK80k
YKbUJVIGbwkq3a4qyF7T5Wc9qw1e/vxAmKZg53UrpARC1SqhyfCtkpQhdcrVvt2D
uEL1VkyKY3lufZ7lPpvWRGl3B9CdhKQ7T/Awx2MkfwlCbJWrV9gxSk0Gos+tCaLM
wmavoR7jFUzmtjpn1DEZuBGzuczIjfdWdPl8zEptAgMstv7lmjynmRWyMBuf1cfa
aHcquyWfSx0cucu80hHH+N9cpHPB2bZENnED+MkHA108rj8PQ1koiHhi92CzY0Ku
mNHfmtaWz0cRtGRah1x6ivkZEfyGJPEUL2Jzhr1vVxst3bBwM/G7CcZnxlIuGFJu
zTLj3lMLa5WcZtOHYruKCdFnw6mBnjwJJ+7z8eL8ds6nRO0knhPhaVmiV/TJQ4zI
ohdCd1xT9IeHN6GJ9I+rwt27hGa8UOX12l7wSLZHiUydjdpn9RAnA7gqYGsefUPs
mEaESzm9KdzOm14l08wrzqfBmG6mRqvgUhyXRVy58OF1ggwkT9VG69QVar9jnRZh
1T59Ew2LKpBwCG0Xoiwn7dad+VT0Qi0k8tLLCsgI6qO0XSF+jw78Z0SiwKzTcUxv
aenxqhgzfzopmBEFXDpqNQTAxRHZnex/MkPyVm6P0g9bwYgxfHlfPaBRnvDbiCS6
T7c+c8kAd72ZuhLvKLVsHXeAvDR4HTHcK33CNumSKCcwC5mLIcoUkxeyr9KJyF1L
VOORWU4gtl+IOrODNRBs9tmqBhZEbLEbzOzUaUYO4NBoWE7XgYc0Ah/l+ZplDnsZ
SAmPBeiYgNCEIMHtfQoUMe7pku6nUSuc2rzlyZGhmsVttQryZgt6I1zlt4KgLbwF
9zaCxPdjht9laPquJuA2kFU853ZRdB9bb49PI7DCH0izPh46NTouQ+nEtN8vdfxK
uZexFAg678fOlB5gtg2RxNHtognHGrmj+B9V9/SU6Wr/EgRho3phplHVrjz4ocsh
01UzBLqcmy1j25CuqF7tIKYx+hsWF6R8FobbcwpfHEA0XiZszurHKygsNqGx9vro
lOske5CS+PkZpcve9esxwF6b91xFzo7zcOxWXBYAGghpyeVyMKbkPTjxXEBp59pp
r605h3dyNb8GPsEqVYCqbTBeCYataFe6NEEdQ+dYJGo8lerSAwsiE/OUjbtH6R2Q
ng/hrhS0nBnN/nIzEm3zywgNDi5ukXFvH8YxKns4Q8xRiZk5hAC9e6gax/mZUJaj
OWdKokCse3XUJzjsDQFGVzE1ZwN3nlGIfw2S3dw7KkBMjkTndK7Ie+dICN3Yq5U9
j5r/2/HcDdtz2mAtZUC9u8Woa4Efs+UFdMjePYQOUt3Ns9WeDRIrP4zdEEPOgz/9
UNSINZvucPkDmWWs5MrpXaTkF5Q3VGVdScdfAp+T+uAjYFzl7L8kczcOZtEoF+Fe
OV90+yzy8tBVchnpwbVEsrLKeVSu9uUqZF3wrKHbBOKbi5BKINwROKFChVHPL56u
hT8sUPyyZGyEFq7NVuVgWmmZ2KgAYa2Qru30wJ1cW5OUxduezfhj6bAs5Ea5+6+p
Eh4CitgZ/oqqvXDS/HEJ8g06mNJTfYnQWeSlTPMAk/njKWl0FEgj4FuD35q+s2kE
2tqe3zT5gtx4aIIzOWU+GyTS4zwRx3AfojsSKCPkf4Dv0+7DtrZRyVQ+z8NzFFzA
EUF4lCTSi9zSIpAW30PBzTXxxl0jkUXzegDABltE+oydq3sFRDcxj0zzLnf3OK3a
08Zkkj78e7qLuNwRvvs7J8if0nhbHODoabZkqf7l8ny1+Tl0Eq8LmtOnxGOltEie
/dyMvRzonXzMv06J8JCrU4GSGkKnidG5NZy3Zk2URj7nXh9DVzk+GGcG2KI3LQec
b1rwpeGk9J4WquSxJPmQuUXmNBma1l+q98YnL9jNuiRSTQp1kvrLnusCTeNWPlPQ
OrsEUO/uHuOGDyrgeMjpx6v9H8BAQFfChFy7itltHxnfb9YnlnEkiMEO+OJVP8DM
ZxhHcgUeRnCjq0Wygxd5qtC4FxBYJw/3bOJ4bx1tuwCGwxP5dC/+hRcotl6bNaRt
4glUIcRuh2i9cZYqY9sMPqTyko7vd8u+IamRO5yLF4q7B+qcgY8air4pfjroi5Ol
4ct9c3seNGG5yfe7nu354e3cDTqa7KoPmnzHEGRPceMXD5p/xEnXMQJ1v7Vip8rk
6BMtyD1ZiCD/GiDasx5WlbbTdalbc3K8UDcHtY28R6RipvmWgb5Iqa0OC0D9b8bB
NqYYQMJI31ZUyCNbBCazvnzcs3HTG7Z/7USB9tURYv89VKo2cGvg9E1GjblJ0y6U
dtjHPGRwUMXJ/tv7yiFZpYJuBoxDVTETX160cRJ6uZcsS7Nb1wznLdArufE/NL4N
/jZajSPDVkNmuW/M+EgPn65g92HfX2OlDlOcgYRCIGpZ8xnTPGRvTxPJnsImILOr
Bm4XM2jFQBPlHn5XW0/8miccT7QWweuPtSkKr3H94af/uq3fxfPBybdZLgBAGuaW
GFtG+dJ5I8F6Ze3Ysn/ndNd6I6PzLs73U1l+obj7/lkYXrukn9h001+K65c4pdI2
AAWH5MUroT6h+Ez9DRPI/ObgzJncHvyB15heqqOWkznbF7V8QFcqcGryI4+84kSF
oC+XNNBaJR3vMn1SJQFJ5sBY8DztnVQ+EQ2nCGJy2uJ5banNyxDQVxXAaVCAyqau
Z2P3USufzWii5BzdOQArzYLoJiFqOcqyo/3jwX1Qh9hzE2L9k4R9+SsXbW/Mi2zD
r32EF4E4EsQynPCig7pIIm5eOYbT2yefKZ0O2XzzCNaqn+stCOirpNx99Yo9rDZo
kN/3g2I8AKx3JPpK9vqmWQnY+The0Z5I4Ej+kIFp0dY7WIBu+XEYiwF8BdP4XpL5
WqMz6xnTP4N3Xhbd8Lvy98Kq9aDtz/m7OvgDlRIg37meGaXHrxwrvAT/DiYI5Dpi
uoIO+6em6AL4DsSeIe3mImaNanwI7GVPTdLT8obw8trZMcjLJwLDnsWA6OI+dLL5
clERWESHS4nFCHt/iw+YVlhc1am1MUZcEbcOPmkD1an+CenqPCtzQlI5V6D3AOl4
R2UHiV4VYsN1AwVo97J7kMiMBjzKFAfqBDWZhOOhscCx53xNfo1odHQ1DeoAzUed
nH8D+c7TI+aens0etLCnD90fxD/ybDR8Y+rRDfgUkcl/owjZTDowMg33UPfs7YKh
H/Mcfo83YiPyKMLFuy1V+rvUsfsRHN7EWbKh1cfZy7V8gYk1872J7t0sMqhdNJ6x
8jcZREkm6xs9EpLrVHxDacNGLRIEeH7yJf95Bh1uz/wXSnx+zg3RmqsbXNDYc0zD
UsgjVzNxiS98rXxjrTubjN2/lxWAA6ojtIk7ZEa3mzkfrr+wuHdftYP92jpTVNBv
C8gkarQb9DdeQ0BL/xpaTWe74N/uQ9sSttGJyhYZuAcv19szBfkA5rUSmBGlyhTH
JFjrQnvnyCRIjJrJrLS9spEnXHM4CkUmOOzJAr9Fh4AnB+Wfn0qBs7QtTSAPOVkL
lnaAC7RRT5b785vg4DjAKNANpT6dVALkgevdlA4904IDHi9R2D2iGCoY6YjqT+ll
/1acI2KRRfZmYguNW3y/0z1ngRJPLIifBaPca927GUhx2TtCvaKQsYsnswHu5HmT
CHP3gYJ21huMaFKRXEC8z4pivEBlXh19HHpgJQMUv5Rm6Xq50yHXeG0MLd9W+L7Q
BvuY8vUBRSI0v/KTHr8Ylo+dUQW7KaCwKJUQBX9YszHGKWNgSXIVyKmtViE7BAQq
rmlioRUXtLu58u9lthCZScG562h6rr84VCxRqr4JZfOglVxhQAU5LSqOsN7Jo1NH
oOAZ9M67vE5SiDrtho/pxM3dZM8AsIrZC3istYT32IgnJW2ezb5YOoyxBxd0jGjO
092QRAWCh1uhB0TRC6bLNrlF5rSWMmOYUFO3xDZ96ggZ6W4QDDFLHy5qCJYusFjF
IIVGZrzz7cOKPwXrezli/4tPF0GrIVlyDoUPzNT6pGe7GCcHVFPYFLBMU3GG8KLk
0NTqZrVIjv0oISAbGpxF/WX9yteVxxnhO34fpTgfP1UuCI0mqmQFNw+SD16G1RVM
cro3aXMXC1b/sTaWhlr+jkPDDN9rwVEbbZ5TGK+QjKvPYXvIm8s6anspEtZq41yH
e7RWt+/tgMwqR0/kt3Iml2GqwJaLWdQApb+FJDYJHd7rkBAZSbfaxIxFnGuWBZKY
edlHI03cARh6Vg4Ok+dS8y1GUgXIlDm8T0lnNd+hXS1gZhXfz9CFAya3UjQWBELD
oHVZlmSy3hwYLSNJPZrfM5yJndy6lALw70eTKp3eYm5Xxdz/VdO/0pexTPz8/Yqk
9FAOuSeA7Il2BkgNVl+wJriF8b9vbAb0yAOMWLL5e1koYNtDZndXaEF+zdcw0J/8
FjGtr6o4NdZDeujTc43zz7jUb38V0MlSBz96cpje6yaXGafLRqMhSgDruul/c1/A
Lun1gGXZQ1iGSwXK9FZ6aPo2WMNmXAkcJr2fCl34RevfxOHfE8AWYTnDh6VEkaUM
QXds4u3SgbYTDBkOh1sB2JhOAr/nb4x8x9pAEWNqznnLsS/E2fIfJTP67iu2JvJZ
6irAAyOc4Do0XlDiEzVcPJXOBi2HMfd4HgDpU3EWb2lmxcEo+BgJszE6aLNTmq/G
T0GCKkWEAE6P7Tge4UXdouUPSyU9bTM60FA2syvHDtazmrQXY5bpq94eSOdMRoZ2
pcHoxX7wQRfqs2CJcZoijG8RFLvLGjevvwf2n3qTuey3LGa+AcGqh9H1qDiE1wWC
OGn1NS4RqGiRcFPhYmFVHMIztW/A1zYR/qSJJqjjm+7rx5GzNUId+uV5gMKDNDZy
ESErw6+b7X5DKXdSPBdpsGYlEdhY9JdZkqW4td1ZC5donAGzgwwK2e/bPFg25Ger
L0MtR1/nwW3r+K6g1/SSboIaewQAU/VFROeuhB+6PyPiXFBkIZkFkp0jiH076qLw
9CQ8bYz12gOOMfJrb0ecOkKrC/7p/SVY+tG9ktUW9d3lm3MMIUZUiFvSIYY1tzrA
QYmC9iQ4lVZxPd+SSjS8HuH6fYJ8oH1Esj71G2BDAAgI0W/42MQ5LyodyI9cWVpa
Ct3FsjigIxqlaeVxVpo7n+M+zj0TqDeh1gaFmr9EwyAzpOsIAzcg5NznRMBSRJmx
Iv730Y3/TT3CfUb+nTZbDoxH8h/JBAyGdUEhmCpFVvN5y4MV5jVgZpQ9uEuiRdII
pwKs7qKsy9vpQODa6goTvhovNkiJEGWDXWB8wLiegiEQY6bODE7s4DJiJ7Dy0n5Q
yyEI34Tq5SQd4Z0B8NJ/UigBtWGF/YjXBcUVRNzsTk5cIBeqhvWnBBUPo1GSUBJj
FsMsZ/OF+bsVC+mV72JXLRnigInzQXdqavATPVb5FlPhLtqE4p9wu7Z+iwb6neJE
GogxiktVtB62w2A+5cwBG793FeHpN3C3N8gmOtnm6rvCETDU/uO0i9UHFattK7gG
92onilUioAzhmEqBE72fQhh95ZZb+oh723NwQk4b1I/e+ttmcMimO3M3JL6JfLeS
rvt7nZI0cuc++6VGK3r6MflkezuF5MfofwUM556oNO1LYfu+eI2cY7Ao1sQnF36m
m+ZJCl/YOTa3SSK3BQYyPh07PpK+D9vyysqS4kQnW4WqlPiZF3dHQddDm3bmCQTh
z54/eNPS8FZf/gZVaCPNDpJc5X+xq5lxhiGcBua+J5uQZR6Q7qAsDsG/cPSYg7DC
AZiOwkDKgPfRRV6t4cUXF/mTxVMJ9/2kIkMn6cMoAYNiEjgPczbusFP5PuDHW3wX
4X79V5b9xJLLQeuLytg7tvcuXpnmUPwrg90Z1Ea2sQ03CqRlRsgKrNHzVJDyfxYF
cG4aE/uVcB9PkMn+iKaJ2bDwjMMVYoReGTAy0i/nzqb1rN3blADn4Up54hQWbx8o
EEaIKlqQjBhokL0JUgTDdkfXl6AkQTeBjn/wGntmHAgKszJ/D1Ehnvzj9pvX03Vl
UKqiMAsUad+ENVk/qVqCODPIbZ0r5+ZPZXuFLg/BSkKV+thlGgR0SCiK0TFJLCCY
XOPeeI2WFfhh0jyMu2AB42b67u+S4HbNStsESX+s8/KqNu5sLY69wCvWRi61DI+x
4Xboy+TnysN3ZDNrzPGhcDLY5Sm97KodBxJlf++UO5Ri08z3KXHYP+tbGEnMaewD
i2x+JTipi09Ucg/2WtTuQuiuDQOWIvG+Dhche4kSY3wVsXPSaytx48SjvSzQx44t
6EI0ve+Dq4BZSXB6kjWNyG8FJErDW8y97iA0B9GNySi1A+NTWHSK4OpeGpgtwWLP
W0rNqDvw6ce5t05Zr2ybhJFv5HyF19zi0XHi1/WlToHkEMlRCf9r/5NxHFcXRM7Y
T1TSOnIjfjzageGIOdgweIZuGj2h7CZ3ox5tHRRe5nYaAcRUQo38Ocmlnnj7kRjy
kjYwEJQYTpJUrGeQsqm7wkkSV+6rxEZIm0bkmf9lO9fMIdg0mCjp0g38PnEj0KHZ
qku4gc9iPyQtGoHg1fNpza8X6P4Hh1a2CzfnYGqsDN3F8VFviw7ksJcbyVIN8tI6
TI+S3tYDcg9bkI2NRSAnouj3Af/Vz0hHzhE5QjTfUb1nuioM+i4kHCtSqkfdqKlZ
LYiLqbuy2VrnuofZa1nlXdYSrliG4RKqa9qNNwnpiSqRgDXmeRPtdCJ0ZsHAiomo
JcgRHz5S2ECYyQvqPUDw7N22GrJvaZq8dS+A2aDG1j9olkFR7pYAA+pH0ENtO1qQ
UoS/LX9m5q+nbM/yzy9zlmZU3rfW9nVo4f3krS8BzFQnnUS2+lP9fwMZCIYeqDc2
7ttOOk8sNhzlQ6hpj2VHK4mDsXXwXpKYkyye2MwE6qEAEUxDVpIEbPwCDbVBeKbC
/J4g9S2/Chy6KgA7Qiz2RB7ZCMKpIKxn0Cy9HpN5QQPom/XO6EUcZzXBuEZlNv9U
l1oqRdTTMC+Qpz6OecxpE2jcNMHF2jJpb8kBsJxQqNgCXn9p5EX7sbDDhRCXw+aY
TwMxH6ORia8ykBg47hbCy9dXoAZe+bNOPhOU127gD38KSC5gswiUpRi50XhXZLQZ
vSM4juVrThl9uEReHddD9DYXst87ffm4y9dxBrIpXtmY80JXqgfRLA3Jq4VRqNsQ
cq/xBKV/Lsyd2jEFcedIEXGnvgCj50KEXy3OuKwaTqLmAGYYvqnt7/viscV3I2Tf
Owx2AdZq4Gb5Ae73Se8w3pKg2SQ+dw00NjzX0oqk6+dOmzyBeKGYJUEABhU0s3t0
PXJ80ky6bSkVm2+kTMSTGq1IFFD94hbX1Di8oMspwFZ8HX99/KzNK13VpfrZuqUJ
2JSMszG29xSk53N9cEalCJzB0TUrhzjHvKvYzK4TTZimSGrBehGBICAJvQWDLEVC
LxStI5bSxVgsA28z6hFXJDEtzHNS9/cADq1C9AKYDQhErIvWusnHwret20OAYuGw
d+7/pz3xTXXeiFYivQjuxIx3D1rPKTJWKrLOGN3/IqTzg+Phe+7SoNmhan9ooUz2
ZGzm2VTyDK6r11Pn001m1APaLzv30/hoN2asESgUyw4oj+tsCGUOj9N+0bW+6NlH
AkK06157+VDP2f9h6e9Pmd4vP7dcGufqQ8DbABw2DmvMEAiOsADxPuw8rQvjgUvU
gser9fEiCmaX6UxhtKloyM5iw6rnm7CetGs1wVjAaXDcOPPOXezTk3OjMgG8EgX+
LQdkx8RSGLw3pQtMxwNHUiwlbB9Vs2Kf6OJWaU5uWhezZfjISwiCe+P7khhwdF6j
moiUSZIQ732oNarKjYTbxFrDhn1RopYZF4q8a+d1E3oEAWUiLGm2iRHnMI2EDTA8
nxan/CGA38kWuJqiMIbATW/YR89W9ZvoLS+AxZGUzCiM/1ml+X0PzLKDwkJrmApS
zK9axLnA8ZxT+MzRH/G+3+w3ljYaQ0ybYo2IWmKlzAN1dZyurZdpXNR7Y1OV/+Sv
P+EPjRyqy/Yq+EPHBBU68BQ2d7axicB4SMRpiuA84FZ4KC1dpIo7AEDw7D6ZG95i
TX/3yU0oJ7K07U+pu1dH0mgCSaO7hdRACxuZ5qnqcoO4NxKa1sKMjqwvpBgZUrN1
KkJITV93rhtKSer6Du04tzd24cfmJ+xdnpfHZ/DllhhVb91K8Jru9FRYfozylz4T
HEWsgp3gTjXkiMf6plFolMInow7by2B+EYoKNEu20AyHxz4XnT35s9zg+8pRF1YT
47/P/F/2zIdOvDpp25sQxjExYNzrFEiBT6JjnBPk/kDSGO/Rlo98xm8nJqO82KRz
NpuaSKdDXQJl+OyqRVn81SzGOV5HrnqDbYxlffRKALfunFI5sXc7yre8EHqIAoZU
twPjIMAog7Jb7y1SE4E+eEworEV+osqi1E3nTE5UKf08A7v5bbR1Sy8PhsHe9vvM
PjkVDVau4NbXKt2lGzQc0Fp8859x2wQeYn4XTtXZQ9mI8jVvNGnU5Wlb2i0ynVDP
WBSiLh84D7HLWaO9heJH13QgJ1wUp4OkeD+YyOnFxGqDvXUNHTmmH5U7icBM4w7W
Rtqu3/G6oaAfXnJll9iqukCvkf44usSyPWm8FyklvKGcXRbKUvlJ3DwQqPOlaYpB
x2elaWjDVbcD/fKj3KFWlrtwLlVFIQNjMFVhlAI96LQFlJN2Z2z41njaq43hSDAH
m8IRYpfQUyjiDJYiySU3B1ESCdVLZCWWLDJXm+MRQyca1IHCGSb0eN8qRREKBdbz
pu8D+qYMVICU5nL1ydxlCybNTCpPiRyLX66nrW96mIJjtCtiC9QmRTxfcQJV74IJ
zYmQUVS3ZyqA9tJXcJeZFLDTg7JGs9n1ddceygBTy5llFxWYg0pCfIfiyf+/vEWN
RsvzVFowuOnIv78J24ht2HhMcELg+kELvUFOrrH7VJF0iVswu27SWKfw+RA3tW0F
kAJlmDhpcZFa5B/RMgSp/Vc6eQ90rv88NXH5TzoN/3zadeAStzqNDYSND0ikVgzd
c8MiSSbOnfBCoWDlGqJfKkuFfY4nPnJtJiNJcacNPJJi/uvW8VzPqdxF7zuJ0hHd
/YroagzU+zlrUtjV08fX/0sA5L0YOFq5LQilxtHFjJ4z6XgN+fAKvpAoVFfi25oe
fyFN+M/74obPSJqi+4uDbIu5YFbgcGc3d+L87Sf7Nzb5TcD4ZPIO05IPbGA/nvas
FhHz7d/tgdWUfzwfRau+qLLRbq5cXSUKhKOg02F7JSsH//nHm7RtUguLJMqHRheP
gt/lnpW67G3F5cM1R9vXOzEK1xRYmYVPvq8Cab9B+dj83AxwG7MhyQ14itZf1bst
AbGNlFgrgizqNnvl5CsAQpN3LvMUbcqRCB92vSCAFxBzKaAIc1P2c6fUfBga7T8l
QXUx2xYw1chKpu4i0jmmx+sMnsMCo3AzGFv/l2LLKL93/0MHlYMs51m306x8Pz55
DA+LiflDxB0BdH5mqBQ5UTvvRVb9rQvqoRvQ6vaIPYKWslecFYXcHMNhREWBxCo+
+VxsWsmQ/xNYPQa9mJ0pkR9v/ib8eaA9KaZiWrWjDTmb6nZbjkPykiNxqGcQph3q
C+kxAweA/e6Qvt2KUN/cKQO+pCaJ+IN1+NKuZPn0lXgZKk6eXKBjOLSOL0aPbdLc
fMcK1mo55dhuuHrGZ64bPIcCdTAbJSkE1ZrE/oXAkaSuQ+YHvcR40BaJrSLqeG+x
uSArKPXG3nNEB2pXWeu7DxNIXORW0pg1vqUDPxN3FIC7DwHL2ZBso0XhrfpW4o/N
R5dMwg98hZlaA8xj4I+y/JHmp2eM3JpnndWddGU0QHuEP95/kppQORSjFw2gjcDy
D/G6WBLLDn9gGeq+1a6D+/jLH0TMH4P12h2bQmZ980YSrLg1F9XOM2kYVpLjXrTr
PPy3GuVZWXNRBUadEVYb7avB4+VNARwJvxjbeioJqpSmLvyi9mAOJoPLJ4OW+FFS
ZC4buypmvWh+KQ4//rUSVsrQ3rTcAp0hTNvJrEtIE3gvspG4J3jHLU3lrcUDlvLA
s9jhQMBwG5PMFx2TBZn1JrRxryX6ZQb7pp7j7s5UdPs+hf3Lnu7cwModkYRQ5Mzf
PcAHkog3C81c/JTc5u3eNiv1CK+3Pem/LU7IXFZPyenyrU2J99ppBXGQAsCq9SyG
oVlmqJ0/Ju6s+a5FNmmLQ7yoXZlAqs3uANKwr6SDL+QghK0gFbprQU5Agp9ImJ+7
csF4xtko+NXVblJaKqJANa5rubEzkMISvX00fjk3+SLs5Jkn328rsU+fYEl9yIQr
R2B75av1WY5py44YzF7wYNY0PsTMSRVyvp7JGhpgiOdnZ8M6TQka7RZ6hkEngJ07
g4D1g15FsM/vrKd+EwK+jQT4KLI0QEYVH1WcHiYDKzcum73EAaHYO2OhGAjPV5Gp
U3GdmvcmkKpr77uFAsafieiOQybG8nQAHKBi/CQpIEsDPl/96k7fuMeNPgg2LOVP
17wzpyq8cR9Mmq2WZM6JlWVncUeBam4c20e20JMbOcTtWBNCkrewWXQAYMOrjH8o
xnnf/DW3qF5KT4LexU4M0I+Wqs69YBIZ8L3DVX3ph6uZXCKgdMcUPVX7E0yWiyd7
PpWQxBE6ttxIbbtRrlpKbgNT7kIUUwkj7RoJu2xVI0F447AgPqxtPk4BsQC9D+Ut
h+iKBd9gxLbQBBQNVXzdYJ9veOIjEwUaCub1Nl2Dl8I1nrhAxw/sItwbc62hYiJB
DobroRY0OoVBOuMDHo6gCwhn4upVjFL55OVRa5h7pHegQ0jHm4HvKc43coyWeuVT
LCQRhSHg4gBK4WevtPJos/9pkK/+OmuXcPkpmMA7eH/wi9jojBa6M1h3brvOg7o2
zWv2Oql++bTdbdJqVUUZ4vJpPTx8uheuWp5nPYShoG1Jh89mPHVtMiN52qG+li6w
yKiFmXqKS3o8oGccAQbgweE77PePRxOb/Ghma6AxE1t0FvrApuHUvR6eUtJDVBim
TEEEukPlZbO7SahimpomVznPNTHGAa9d8msAheWo5W1swjuwRIFQbVWn7QY3ijrt
QqgIqlVqAv56/SdIHKkvx1I9DXh4wLJbzOhQH9MCqXezU1ERhHHm0+vZRINXwdSg
moG6wkuPG6Xs3MLgrvtj/YLfvZR3dA2FV5fHyFChxiBd+aaDRnYhywxQ9ZMwJgcb
UtFBINOcZPSp3DeA6jx6iC/MWazv0EgI2TqbaHOKb6O5k8Lz8lNSrrzqtDe1yCWZ
dhb7Xp3D5hZDhq9HYYByEwwKBsFR7B++U+tlGmGjvfz+9s3GIbEf5bMyACuuEOfb
2O1vhhCphMj32BYoWnVhydQp+U94LFRtRPZizuN76mxZzUbnIwt2XuRMXE9zctBq
EnXus+TImrN0DBWrYYaaPG93Pm9SL8zfxTY4nQS8m2+34YDc2yPH1PgMYd526rO1
kqiwOaKXErnu9V83bb2uNr3716Lz67N6/ZhWOcRyilcduwHtVf1RZ796GMNMJdEh
eGTnpFUTBBp8QvQ41yI4LAuzGdIG0BND75iF3a6Xf+t2BhFQlkshUJJFtnMq7hGc
5ewLblzEOtD0QH28vTIsDUV3Km4YhsXIG788GJuZQVlasb9Ot0DfIFQkBPQiUfcO
HTcmyx1xjYw1hawourtA9ZFVGQ+wJ1Ya/zKMMl6lHF3So6pH564wwkGeMxnTNDrV
yPbunKCAsge7kygDTHfDGWp6vDx4B4K2K+0hEX+nRhwNVC55m6EyPC+zwOTfFPwP
qEXsVv5bgzC7WcJ888WpDRr0wyHD0pk9r8BzdjZ17idr+6VQzIb6Vk/8hKR8FtIe
g/y8g9MCtwuDLpkmJ0FHC1jQawarLwDFfNdOVVaCKsJmN7CNpkVqB1O2tizRbah9
/LanU8e0nAe1CXw1gDjjQOMZ8A6cd/Rrdg/7gPOpVYazQ+GMOWGOx8QMMEsgTZAP
xUY1iQnpRBegQWnJ87W+ct5r8l6Ve0i9AgUpMn7JMNG52w2pITNoj9wutUrKwU+h
UfPPL/tt+DJ4nhu1Rf9CmUqL+RWZvRb/GzD21DH+aAHz02/mwHVsmnAgrcb056RJ
NqgEy5vb6Mn1v+8NkfnKsGgYbtoH2Cu/pvGklNE6xO86U7BoAsyLmw/H8vDTE/+m
+60tfO4AMPoGYMwsCXZ3vvG7mIrSEe7lNIDmqvOjlniXUv63NVbAZ4p9bZCOeIbr
B9i5yH7DNDu2Bp3Z0pv35q7vHXWTRePEmUo1GPVfFmMoRqeh2KpSqChP6aMvw+7I
4As93cBMezO8ObLwPHnRpPnMmorwC0uJEaqYjUNuObZBpE18hHYyk4dbsX8po1f1
vA6hDCdbum+TuJqit0iQEiuYMGGonJoWsOsAf/YgKW3umUKo78N4WofgIVTokvcG
DHVJbt4JyXYfDlfXhcOdnvMUjGp6MjZSWGXh9wf9AVhRAt+Xpj8Iy3SOekaex3Tw
wbuXPUjadayDKXoN/BTkhfX2jtxRQYOsC046pKIyKmgsiimjTyx7thwN8z3zZV+x
Y1NdT1pe5bPOa8FboKVMF0apjWJ4mdeKp+hpfGmCWHoWANjA1DkT8y2KyIm+EPT7
KyvT3KETLUCz8i32iaoElQGSJfFljGLGd0TYYvczPiMsJEHsI3kSJnzPoKONcEFv
EVrYeX9uWE1B24G0rpuVU6uUXLGix8Of6jKWa/OHZG1BBUAGDfczW44wBrKWX2sO
M18gZEGkCtD0jyJY+nd+z8cJzM2BBajh9lRrEIKndtxK4iu4ecb4JYSM7jb2Jcbe
kXSmn8XYjGSHHqp7LDG2h7YNZJJ5hpm1ksXvQImeGuaHQ6oAczUiMD2eGqfcvQlf
9z/ULYCeBkpvWVfWy16EyfLgl24sgnsRBcuZ+Ux1Sxy93T3ZsMZipsQoWSj218mM
VQZfs+o/v98Jh6ZHviVMhRj5IsjgAkgXg5VN7anZyirvDJ0YekCLJgWERckEgYiG
gEMrrLkzwPF87mMGBB+EMeNTWXglHXyQ4FXBbnwDKc9+fAqbOY8SzahVxSg3BR+R
M9509BJDydpqJ6EP+kroDt6lAoZK98iy8hj6OEJHfxtZFjOlbHkcqx96jLMVdF0q
BqLD6AxQ67nsNy1FPg0AJob9LDkmv6UJjEeSJyar2HvrKfHdAxITig2dUgUXifJr
Sy5Rae+B2Kk5H+TMFdHA5C93mgCARn2YuJkqKO2wH4C/QShxsvJnY7X5KrE0OaF5
vXI6OahEoXjMzDL3kBrSbw5pysn6Ll6zVgkVsGrgWgvbGDG7kArYfOyIMDhZRgLp
d2sWDSFJn6RORsU5U7hiSkZxtlYR4u6igssWrxsETFlHYGhTTWQ0w5TQ98fhVGKA
KMZDqCiVv9lBccERw9kAlDlWj5KS54t2Rdok8tBCz17mu5cA0dk3IMfVISRa1c2Y
uiLIPxs9Cxwtpez95brnHwgz/K4ba0szRpp/G/PQFyG2e/5okH8SqEEidxdCuzyz
ApD7KLeuZ3XuRUTYh6sTTJqwZkLJ/r6NPKBLx1uAz67fchmrs8GPC5gE9C63NfF6
3XC/I+IxugicYPCOKMlcCnWLWx1s7dtyeGcVvPjyc+o6oTKDYvEHfTqrQL2XqbnG
+fS2GNMjdvCozre0AxHu+N/BRdJtWsHiqvvNPccDIPyJrK86i79OL84BQFK+B3il
cG0kYYTceKPSONcWT6t6ZbVLPGGMZ/yH4deLRtZGUzm9XN3PXux2phcuFBADyYAZ
oiFN1ssyfphEOCLEcaQ36bNchKI7lu1q8gL7E1bBkxouJpGz+62SYNLYwZJZYaFT
AUStGBBJ7NPcb7y5Flct34KXXAY9rTWOGQGNXWIXhQIWPFv87uelDJ7YN0gold4q
HYj/fnyW/qMpBySyQHWwTRFhOLZ7/7FkBpuhv3RN/dR93Pc/QSlw6DEsvagjNY4E
onNAh1U/jLQYoAc1exaJE6W/gOq9A8uyJ/M1dl6MxUmBcu1/ABv1qPb93fKqDD9E
J5DJGPzx4VEaNZJ/gMl1qnxXBsJh0NPV6+NkZ7yZzvuFFW4n5qyxGnsxKbiWkz7L
ktja+/Bh15351a1z7jPh2SvFd+5YDj9NbUSCcIa0+IKvJarjfzsPRwjSswko4N/W
Rb2GkuIFDCOtjIUSldaZMOc+RSua8wfXPoZ3rd/JqsT10cgqwqXhbqVighPQVG9r
dydsxJMo3dnnlbWUtxaf62KxrM7Pyj5xY4GlC2UrP/r6bDiLL07FNMXhgNn0QgpN
ChCmlX/CLuPTKzzMqJf7u9jech70Ifj1PdbQw54huNraZ4uPCCjk8dbRnT9b09Sz
bVO3BZ9DHIachMgpkMn1Ce7EKcM9DJ9PdgRdLLA88C3yK4RfiGKMSDsyFOv8JQri
BMd0ttObYW3CbPWAb54Vdrs7NrkTsJfnhKgp2heAjyDCyi64E+3asmO6o26Jj1Vi
KyYUl1esf/yr+eb+EopLlDQaK2HuhDmZIn9qnE64pK5JPGdg04I+aloor4wcjAI5
46ZPSLm2KHhDq9Eln6neGaa25hiBgz6cF2nUeL6H+46ajBxz4jOQn9hd9V4hFWYk
nHtsBXSJhO1MsnoQuBEA70fSxDbP9R65KqLQCBW7Z9fiHDDAiRLK9bC1ANZM0zme
gDgoErArePo0xRotBwLxvfM99h/Exn+sfNj4OVM16j+8U59k5SHMcNc9xJ9HDsZS
VzcBEYEBl7O38YjDWSRlahKp6ZcDRBDx/agZqQXHoSnjQC0Mub2xA8ZIaZHF0Zan
/XZO7VLY2JTej5Hfpys+WGgXe3+F/yNvJ7IDAKPj45zxeimt4iKnY3OuB2aqONcs
by6MDlPry20cet+U8dm+TtJrt0Tznkj9Gil2P8Zo3iu/2vIh6qYE0f1DUcUf4c4n
HADk7wdH5jZezECs/W58VHsU1+zQQtr46qYb72qqYBMGMKP2Gy4iEOIrjEWvp229
gKk7qNDbc7YNKALGpfkyXAWfYngBtN9xNN4zpiypQCYxIlqAn0wuqmg36Ok6nQdk
/yDtjEYbShKfSKCJFdwKvS+H0sTfpvTkizb8wb3w9OGugu9YSj11n3dP/Z3+g8eY
g/fnRiKKcWwx+qB+iNQuT9nXNx+9WCIc6io8NkNWGS2SOpf0xBrXtD+Yh2qyxjgX
edq4ePBoGhrDABSU+PyG/V3QkMUYGNWf21Xl+Lk8jIzuUdKU8FpQ7tte32GHNByp
T8NrvSpwx8BoChw5lshdXYHPPtXVCBRY3WM9lphDuSQqIcS4sRvQltnvsgzIZfon
9LoR8foWWled7kR/bp6ZqWAposfiuJArsH5CpCsyR2pXgIQfZjXw5XpNomQmTv7S
nIhpiY2Z95igF67QAdG0pGqngo9Sm7/3oYVqM0w6IMrkDcQJfNgSwp8s5xmVJXhY
6M5N/FnGu6IY+rg5/Bd5U2IglaDiOQXLwqx5aiWXD413rSooFJd3uaT+mS+vCFSB
QOgPw+GcG+sQoZe9XdEELRR78LB0Kwa3zmTN4uCZHx/tHWxaCdV7FypMfxeox0SP
T6uSbiaDqT/RTACzfT6yVEoiX+SJBQKKvsIyXRLrWimEksZMf3f594AgLboIBNRH
pmqx7x2NJjpXkT9Wr3OL4YkmUBOiqbN+pnJoc5pUn/e6RA+tZR+gZr9YktbF5JAO
vTzmN/yYmNkOmm21kCbgpdIaDzji/PApbUMz45zQavy/LpcQAOimyGY48+T0V6mx
zlEFO5txk+go9GjhpZrD3tWQQhbe3bN1EN+XPPrmB5luD+Qph42dOX52iEqLhXqo
ArcwpphMkDjbRnW0NGPkI614e3NeGdWcc/PMkmE15XjttBnb/GsflGDcHQlcIDet
GGkfwqK7PlEwse0f9md0rfccCgXFd5SJGX/Ky9m4+VBMqAZgPLmnxHJIiXGGi/+B
QtEGAUlLH8mVSOdGc6yZNaEqNyhfRj3LaZwffPc8LZBbOsqK2Ei6qFNzUa7EMMUu
MLHd2IT+OgJdks07UHNGjZd8xuJPJ1mW/5JWGK1wgte5jC8PcY4kIOdQ7tPO1BwT
QPd8+Mnt5qraOcCWqxNItTqxEd5i0FpgyXjYAUYzBGvQKCtitVsYNTzcHkezl6AF
PRLmnqOL21yLTa3o+aLWfZF3+L50LQ4FAPQYsmzrV6czGCaDn+NAHSx2ftF2tZ+O
KVcTep2SERyQoHJJuZ/QxZTIIo+FlccmXC3LZ2C2V9ypfSpfhloOKzsbcVtNeHl2
Na9sm0t6tcjGtYhjqsurlTF/JRMHeNMzq+LW8A0fUQftqNURoMRhN/Ko7z6N7f4p
UgFMveT3Y4B2UF7NLSmy7Itvu522TsOFv239XYRdnpgvOg2LRyGQvxtVWwpnzkHz
VzNeth/wR8rxrKKkbTAZV5XhoywaymMxrcj/5s+Hjs/3o9+r6q1Vj++ltZyNuukN
MFYjHy7X3z6BTfItfobMUhEnKmxjrRQGrqbVuWCjh7iL0/UQ3k6ZSeukMDIzzbA8
46R1po+ZjoyKXwkV2qtlEhHcnzsDhiL8gPPXFYVDWbN/ewQSLHrw68ZV1MuaI5aL
Hpo7kNmkNXDzJn60tczShIWji2wPZ8t88ZYLAKnnatki+y+H+AVdAzq23Noi3Buk
a8JXRzcUQwcXW6uK2vL8zI47rNwSOs27D8GhpDzz/t2V5eZm+2GIiLCv5L8AEQz+
dY3DZ5GM93ahxOCyke7dspbdUt/FrJUibeyX10CUuc4/vjJfw16DwXHGqatWOR6I
5yi/VmkZwrT6taI8wqc6UGe4QPJXWeF4uvIJN4YAfbR1jM3VFRnqcRyaSu07YBkr
v1mWWDdtfH9ty9eBNgdyFVQ5YQKtsLIjhg3imiD170Q5GojpccsyQYB4WFyGHMJe
BCxCMH0WqNbyMvoqt+AbhqrIovr3ZylYd9rP2MLrHWqocw2qtx81nWCz86f03I1C
HPh7YL+RG7OMY0m9+W1sADihcsg6bEuaDnOOMtH4SRN2sd4sXOBF9KOSVB5neSy6
A3i+bdI3NQI4Acn2kov3xaMSX2x8rUmKab2c580VABbghJNvuKNMOglG4lY/r4U9
Dr9wz6Y0dk1Jlfk9qr5udEaVjBpXhr7GUoCAs3eG3tuIPn83NDxWR2NmPZRlRhh4
z7bpCm3wgJ1TY7xqctzoTmak/9Hl7khgBi25wzGTqUH5/9Apcr+uCLhYm1nvxNw8
W9McanY/6fzEgevAD7AoioVyOdBm2lp5+oYOL7fs0N9CBHLqyTO2MDaIGM6N7iRS
oufQo2+ysnksxKe7k2MgSJ/JAz+gpatjBLIhZybmRMCuUtHm3cbjhwV3S6VSVct6
CYkrowOkc4zBqO1hs2LyVjXGcE1LSaCs59GyJuZrLbtH12gRwQVIH9Z6vHzH3yUW
ITTJ9ldcfI3gOupCku3tW7FfeHr4vcDx6lUON9uqf1cPkJYOSukxcbQHxzQ7huFY
/kzd6Q0MQByXOXPhqsfV2rYvz3GB7wK0IoIFyB8KWmQz77WNhgR6CH9aB8hSGohJ
HXj46hUM5IKnbS2gbXOXhZ9FiZyOnA/Mm7bgqS7IVH6s860COhZLp5gXlrXOG9K5
7OVBlk+Tv+7DBoBXSHKrQTfMQaIQlj8eMf512i7hdYjcQSzBcTkK5p1zBpNMfXmF
aMsm722sA28OMHTBVTXME32y/DdE9McS8OhImyAK3vubdm5+mI3DznE56hjLzc8b
VpuL62n/JQGYMeBdImpzmqCREbVkK04buruIVthFKLzcUhO0jvXXiu01e494FR+Q
mEPBfOvJObC9tdjb86YaBJaYnNEA32ao8uYNyrRtimGLA3HBCi2cmhrVpOVf8nCv
tSsXfTP04pTRJviCzUICO/jaRNL7qVyJGvRcHKTLsTHpS/tJeWXnwCCQ/bHFe07u
a68kQHu9yb+jUChUtyq/aAx8bmcPxLXx4FUDzwE0q8Ahcarp4gNs+niQhpwdncZd
facrafPooePrY16W5+NxcuZR09n3i12oAl3lQboha/eypjcxyhec+e4torwWRwq5
AuvHEWSrii9eWuWE3lIpM+AS9isj2bGDJ9UiMSW61T0/7oHsKehgyW7yvUm4YuYI
IxsA3nh0Lmi3OTkctmCO+RsPLvGDc5Ado+BQPpczTF63LE+qkOsw467wQu2WwUFE
EVEHjtZeaTneTXRHenIjRD4IXNqWSEgIVAAy5EuKnURjlGQw3HQD3LZtrmv2Tqf/
bgPrgKtlmNkPzsdJY0wAEaqcYmE4YgzISgIIOODtYW7wQC+xcZFCdb7a1EeGRJ/X
GXD4aoRW4x2TynMsL+funo/ZlQmdCV+W+CZz+7v7zKuUV6tjuZQxvzHhl/vJwcj6
mopnNM+CirGJPhasso1lDENwwD6IHzZZsW8c//GbVbv9bWtJuAgWNRzHdx+C/Nf6
6wjxVQ6pSfp0PjbAClGH8mrQ4d9dIm7x/nQVcaHfWRWHk6DOA43Q25iJjgQgRKIt
176ZNrHGOT4lSSktqAB0cSx+8rh7sJ39STzmAJ5bbqt8BMNNKotsWa3c+6Wz505Q
v8Rc2eoqN5KbAvoNJdVIud62+lXp+loHFui+bARGI79aaHX90m2dtAL/1jissAcS
rhULbaMYE410EGyoqVszrE/6w3UtJLV3qccK8bRaC2fOLX/7jf0vQyG2W9spX+Fb
XOlngW0y4ZfdOKc7cvA74fsEzOqCG0x1JXW3OVtek6w9KDZjYpoSmljaGKf08/z9
DiSVzAAwazNpikKUB3lO3zBjFst67Xcm6onRk84YCwuqM2HBHs5H2V5Toa9kCnB9
pLe9/mZzkPV0DhTGDXm3nwp/w/iY9MQFSDWmB/uxkZW9WmqM4MCkb/VjG5ws6U3r
exF9h4xtOhRBVCGoS5pwYOTtOH7BKba8AvQUo03EO+/KozXlpX5K2s3D6WNvgF8o
MZy3pITszfXn7xPuKc9tZ39gy/cQslF6LxKtGCUUkhK2HRTnmueF5AJ8wQMyjpHG
4qcEUZwtVnKbpg1ES67Ha7GGQCX8dSfU37enKXGwwS4fsxZUbD8A1R5d3D25nFK2
qsxaM0Og1x6la/DOWIrddp259muNxG9RvhgpwCUQOo+z8MwxXTtNj6+l+IWPSo1H
kPpL3iTSg72aeyEpeGLKvGkFp9+16jMRKBFMkl2Vl+CRNRdrOZeh3qOLKg/b/caX
io2zsIF1rNUEUiRvDTPJ9yrU8n3kfEt8+p8xpk6phuqcYmSsTjclFZkOQRwPZqr0
P8QAa7u2lcKUpqkm3FMCY0ioDFi2LLXyGNpoGkL60tcCtCU/qpCtF8rDmjzee07B
feiJSLJIDZg4KCddcux5CyNmcyATw2PU4F+t1IpIVW5t9TqZnQBhsckQXKuU5JYh
2EcgJ3CJEKQnxbszr58BeNI9yxDgJIPBRNGuCsETGcsv4IqNPwoovz3QeqWH+oiO
0TnH11JHGoqqFGg4lqAxm2zWyuKlfiQNNRBRvcFd9/aP17uq8+FodjLyeGzyxCc7
xtw7a523qu3qdjzCSB3PqP4mAmJGVOPYeryDgfoLJ9UlE+FGQaZYRdFizNHqT5N0
+Fvz1tfyfwZ2ANedC742JPEnf9MSL4OA4vEIcxeqODoftx/DHDUsbw6A2p9QLrAT
CSVnf8z5Po/ucs7GrEB7ATGeO90cRwXXEgzoek9zKx/4ERxgoGGBu2yuvrF33RQb
buZwNxst82x2uigloLrQM9iNp1343vPrYVOST/dpRz9ks40mw0WKLgmFwQASmqC6
qG+g8F+8xrQLhn53Nq1ZhMGxVgKMKA5Vhfkyr8++O1BY+R6LpLJV4ijK/pOl4oog
92OU+OMmmqx+/Koj/7GKrssJyYoxqogKuIDFZyA6F1ex1e6kUJQB+Ab9MEJQHB4j
NtJ6XzsP6lFpzlJk0BBz9BL4wqThncSXhiL+2qGswg/neQX79uI3vR/AR5iHrzcX
wClv6yFV220vlpkG7kOIEeB+BrS+Lsx2Dr9/p7k17aIkOyLsHpV3xCrwlb+wHJyj
nFfpuE5/dzmzzGqn+kc5O0Wpp/dAJCrRjvyFBRzCwRaUMoTsFh2zpcrahgvjcq7g
qi5kplRiY3Ixfqc6xPp+aZvpMU1BKVTlWezABn4RjqLwkutdReqLOn5etOGZwS2+
jt7UOBkGGMt9WCnVgTmuGT3hqhHB9hAfuN76JtrQUUynZTxhQaiUdC5jlocYHcN2
4IaffJ7xi0j3pABEU3zowgMDKyXpWfdJOfHpRtHSPY2knLXJ2NHiaKHhsLK4o4LW
j65z9gMHCs28Akk1lHAvX9NKqCNByG4vccseG2Fe/6WS6eKjw2widn7dKrZEiiD+
BCHEJav05DWAP2oAy465+hNkxBuuNYcFKyDJ8wkQv2Mn2hJ9GeTJosHbDjk3ZBiQ
q3s1rFkVQDp9RP2bvmohxdUEekBHTVCfH+YpqOIS9IhFBVnEMAHkIoWQPfTWDufJ
6TnSX/T3z8WXaCRA3R75tel88erjMlb3hFZ9fl/hyKC0yniB2F4twC52YFxJ45VB
U/10KLoyXXb1gJc/dq7QB1Mubgb8d8FnkkEYeJHAHnNZNbS/LRSwnFumS4Nbvldv
u/iSTe+TCkyIH6Nm3JSKk01UuFVxTSfKnWUWcdntOwvh3Yyiq+aY81YDSAVcuX5a
+yFW/P3aQRgs/u99rEK7NEvQxQzasaeD5xbVHF8uKz4y0kxY7ITzRcDuDZ9YQ72C
j6QU4+mwznaVOftmozpQbyDlV/EVdfs/ps24a8iKzHvF3AhIgM7c72tkb86p3Ajm
YhnYMHk37ws6nuEZ9uGE+DEcgmsQcjRmoJRV7gSyV96+5GhNkuYLBHSFw1+j9dvJ
3I7zRzqBdASI+/YqYLAdT/jmaH4IvRaUEpMxi3GV2PBsAZx2DIx/vCJrCu3FHXtw
/ThTEXIYGO1O1liXTVGM/uEux+Bo7cfBb1GtCaavrrtQMKfpqHczXd9iGVh6nFZK
njMw/qTy/+HITA4fy8QE+P7KiZ31UIZ34uH4NDzyVJDJpuHgFbZrjXgMEXRl28xX
sH1Jw+PXDfhHOUwgvHM/4Gon42F3WMW3M2ORQvxyueGs9zbf8BiQ3TMpopBfG5un
jlF3AS2zAWNncBdhpdzbiPi92tpi3z+aemYwpMxumZT1BFL8SAGXTrllxI2nKuoC
oblbOgfYKzi9d44FnNA7STePhnqe0aC3uGbOE4/kAzGHWTn+Z4DeNw7PJccnqsh0
Ypa5lb+fHwdnX4OfNL4LMyPgeD8oGDPlNq7G+K4ps5lf73r/Cn7j8v9cPFP6gKBy
kPCIcnVl7iyEpWrxkIZmhYAhy1/w1bX4ux0o9el2rgKKRmlpHBC6zgIAeC+mEX4a
D+d7i4o1Fzpt8KbIHwGKxtLM8iCTmVaDaKEhT9Tnpg8Kcvu+QrmqmgqYartsbIPt
XQ5wRazUkbNzGWXQ+YnseAgyAE8+2pU5oQJhu1ee/Y1F1cd+jQWSoCbAPSCIBXqx
w4k+S/Ylrkjgf1ylFlWcSF0ei3fTJgPy1iNI3j+E3ZsqsAC+e0LJttcnqJjBKtkl
kYXgYD0G6ktNotpBuqKlENCmZzyWYB20z1IKVe+scJ6uY0kKfg4hOPFBF+MsfltD
D5AQmRCo0v+U7uqjp6120mhN6bbyeHz0TIx+bNoBUMm8IhJWISUhhzhwouI0fXqn
Lc5SSpAOoE7ssT7jbhMrDe1CUXdXSoYhHbC5wbtbodOpXIylN25FVbP6jL/08div
NVW2N28NQjnGzguUF4UFOsNcV4xbCl7ccIHWDXlNMBg3bklHxq8v0yG8iJwpfVb8
JWtCzLxLcEet3M8pR+zI3YlKmNSF7LWAucbaXEG98sFGplgJWE/XjHvhHxLC1a0f
Kiu/1vo2OPKL4ldr85Lvpw+hvMaN5Fi6wdO9ANum3j+Uwg5cqHuKsMm2ixjDZPZL
rYzRJzd9/aVd8U9kr2gi9FDnvJI8lCEh99rF4LcfrEFmO0AReJkRbQLhLz7/xm/Q
N/O7NpMWHK8CDYDozlIpGtjvHOXYOdoutgzV1ozDtd6L/xKWysV44Z9KYSFUhlMi
cyhAi6SGDx3K8dNmZfoIAY2lxBZ9nmN2WSSW4UrPhW9dWxWVwYVLs0H4b91P1qi3
sJVK7dSK7SfFWt8QWHHjAhVgqmTEJLcA/CZg48Y+xwwGm3/Ogeu+ljk/Pp3xV/zf
unG7o0wiUDlpzHcx/yIm8XoNtsKNx1rdMriSu1AVBZATA3yWxooWA2M6v8DL8srI
QsTHS8CSG8WbuER6HdPqQCLUJNikVVyLAz9xvH02v0HtCkPxnr7di+uSrtwmeiUs
nOFSJv8hz5vPcUbkiMFnncZYzt5/wOVdQCDB/7SEY16oZMONRdI9ou4WYrOZZHGf
bhCHzpudMCLBAWyapBePZyDcN01G52iyusAOZOSI7RZo2mdLoZ/ek0ZvIL3EENu+
JacBA1wwUyX902yZFgMCOW2sdic9cZ6UBbP7z32hYfvWG/llHcusZakZbzQ9C0ty
rYCoO00nkDURKJ+nmadTiZN95hPCCIrp8h4ZOspI82E/OO4H7mEPRMHwygwWkqF8
jTF7yDRb0Ni/7BzVHRjO2hzT3hu+Is0DGlilMcKmJbh49i4BJtOV+/CzA19qL561
jFAue8hNSo6sfmsPUmFsJdJxdEHZnSuXnWnRbPdpofQMQ9Zv3gWG3hTVKtqu2Y8Q
I49B/dVAbueLBZCbLYUPLZP40M8gXjnAxE0w1JqsMptC8GJr/g0cqe59mU6gdAeh
Frz0pls9ylYaIQYvHtg1XaabQMd6EiVKEORNx9uEPCkZlp0IgcX5JARVfTWOwXmU
E4W9pEJkQ3ajKwY/Dgxopjn6Ocee+bjRoODVikmI9tXEZZ5d/2u5+HpR9shu9JZq
cggsWFElENnHaqGXaVu4uzMhXbVcPr5aJyYz2MZYUcWxMy0l6hDURID99zRxlHn9
ejYrNDtgrvk9ZiF4o6+Sxig+PQF26koaVkQIfPIAi+S+95C6+Y2drsDGwyAASQZQ
+Q0iJcz0ye2yd/nDBecf2FE4j2Y5w7O+VZnUADlyrG3cpF3mueteNiIL6TO7PuYk
1Uocx5vek/kW8MRK4UFPPcnRasWMhhzMNmiwSHn5/Di08cwhw5dvTuY+Te7mLaS9
JHAaxEA50HaGsV0RIMq8ERbrQHmkkVo9V0Q1LFdEiiH3fQ1x6OMbGbu1ZCqItOt2
ojWgfH2HpIjb1/HWCkUuNCmVIM1ryiXftl1ZEIY9AKkaGLDgVfS+6S9moLX2NaDd
Tb4kRmnv2FB7B25KJ+gLRiBPdyNPjLcFgZtNT/jgnfngL4gp4n6ui25m3Xdm4Gei
8aBlTJ0msliw+fNXAiHOlnaU110o3P+4uzsyPEv/4ieVzNnhg8Xiw+iqZsKIQOpZ
V1y1LY0S4livzT13G1wp7uU0raOK+SGfjDqtwCK8pDsBlHZRQQu8DqT2bp2z5Hsx
1acne8yPz86KrWS9fFXzSjEBiUCO8NgWHwVhxT4EYW0eijRXfOjz1Lpi9+P5q85M
7Wwksg2+HlXIprEYLfP/ZYacxytOmQuKHfKZOC5gPK9JD7pfBybiTWmflGVByiWv
6bRwF1Da8l7jUnU6beNotw+SWR2HIocMSJ8JY4ULxrd7PGa6Z0QaSHb2Yd2rR6d3
wuekaJJMfB3z+xKCUnCBGqp3FbgwztxBYa5tQDv8BRfRovDiZNMyT2dRUpfSFvJo
iHCKkcbXWGpVdpiaUbjRaMlq/aFAZIhgPrTUV871uCnw+HkNRDRL2ju+wXNsGVd1
+vfw95fFNa4lUViFNtGzZcVP2y6sXEZituAshrVeeJMfRxzRUbyzwCqmginpTyG7
kCjmS/HARdPWqBY8H7SwwR9JN3L10IwwZfoK4/efbSjndZ1e/MzHQhlMOZL1fvvS
Qet7U/L6vDrtI5vVq2DffNIp80LtvNtP7JBscFBQNqcHMXzLK/WZVBjC13SvWG62
4h5sE4C2zSUfpvDkd1li/WSr+bw5N/lxJRpla6SjkHNaGZj+t1WJticEktypUKLX
urZBVSZz3+S90e0UrwjuPW72BDtRXstqPqUJkP6jt6AOz0q4WlKmsc0eLnOakrSV
83ynbyZBChQtD8zOgFPmuNoeH5hJSELINF6ZR++4OVHnbURkgCB9sVuWTwiMgP9S
k/4Z+3jAM2/pNwbaS5UcpxE+Klbmw0InD3UbDroF/Ifnv/6fE/YJANuOdr7Niqhh
9ByRYokynmcG4+YUOotXLCnYvBRq5JuEuRzqz/3/vm274T0u6uxBG8U1hZF7FqlM
eOMGkeo8smzwS6iSmipPObHM6yhw2WwGak5UrT7jTEG5JfCzWVCDh7p08Ny31u5b
KRzjtraLbA6+eIfzRe24Chd1ooR80DLsdDQnGmjhbMBqvlE0Xzh7cRX6xUKmSLtq
DwYgicVe54QMXuYwu7gYvvrvos2OK3Wqz6l0pIr4SGP6K1BXvdeEXGjku3uXdW6J
kd7zGFR978QsM9pNmfIUOdtkUojYAPCsn2sLw3gI957pvks60NlUWefPyCVxnNx4
UjwtNsemnUuyEbvgkP8Els9P7u5EMH/ULzqZRZ0EzZcVuSMDkkbNHGlCs0EElIqL
kBgds6cwlJZAg08nTbtxQKSgfT1dwhMi65/f5KDKTKLbEHDYdv24k66Br5QSMc4f
ty8ozZAkcL7EtH4QGwkuMuZAfDlEqwIteNbKD7HEDsQXHDRiIImsxOgCgMee76lP
KdDYW2zLqUSB4Fvfm60pTHqsosuM7Z4yms2EIWK7PjO1k3ADatyghWifw4JKt0db
lzn6sQ0aw4a2ugJsSw/GGPEMyBQz+mzDCjS+2zb8GXwekIEyTlu7OMloeeFZxvYT
34quaKtINDadqVVUffrZEADJaEn30g1Y85PF3aTObMH9AQjXojJlNqEGs4dBg7qI
zwp6xNpCB9MQOdr8uErFnpHTrI3+VZvNCqoQx8/Llh1Mb9ggIfQEIj8XsjpgQVaP
kmdRQjr2wGuTANkn4w/dGGV+lWe1PN3Q71fGmxAn8JjITJ2KHIEAYkKyH1PwyFee
54B8h+yvXRus2qY8ofv8lMoNdeLzewJpzbjLrO3m4xfO8sZCt+3FeSo9r81t+BGj
wAier/MckKSY4w8Jos6Fs7zAkYRMaKMMKYKereraL8KLPQc2ZUt0fchoc2Gn6ufz
Xb6rdIoa6y+dAiGo4BJcg15TVWSq1tfJkdnmjnGtp6sLEM97fMEUdnAzMsVYmrW9
yUSY81274JXYEe+8BSpsNW2+H5gm5E/+V0aTqDvZKYdHF8rKHCLEp2fJHD0XI5hG
sxmuGf8Yak8WnC5PVWlW6+Kwj18sRqfvlh73hgF7pUKYPCS6gnRYpAC4t4IClm6q
guZYH5rtVOTtZjkOambO0wGiBBrox1nsBpJrs2H1g4ie8SMf6S/SFHoruKCtRtdH
o8ex/jiLLi1GBL5OlTuvOWGsQwOuKv/g8N3PB1tLlIAV7QnGkMVArUjpTtmuGZuV
RW+hyWuff7PZAm7ud2uAooR8VpNYrCJkj7kIBIQiUE6TPi0r7YGn9Yzf7viZV4s1
cM1rh3b+SOcHpiE2gNVqttoK9DgsBvejDhdsZqeGlHUJRMqHRJJxY2kwjqmmcgvB
ruiqWvnic/bSWIyfh02aM3gcoVxr9cifSSddx1uruIM5ouvzrFNIvb5RdCmWtiRI
DvS2rg8gvoFNk1MYdzXwySK85lgj38dxQeoh1qfLZXAGKPBtc94sMId4pJPL6/lM
MaJ5E1jNxZBrcLT6xjsYV3u0UJ44pWpjj33T20G+wUn6L7DbXPvxmD10Kj3ncHtH
dWq24P0XSh8cx1a++cHX72OKGvQ5YN6AjCaqenw4ZMdr90YhJ008sXDPimZClJxg
jxCspd0Vw7TISp2fwVrAg7jRsZjp3q27g3hR9Efg9xu+Jp4RjU0QdYof/ScpbfKy
ulixUk2uOrKsmPRG3vB8fTsRK/mi1yBCTu6mPlKKCh9AmExOamXt0gAIE89KGqIK
bpgmIT1ai7MFjSyOAVlo52PAuB4NIzoKPalivRDw2Qj0+K3IP9ZRk8+4uHAswtnd
fKHE6r1tEtwy4tlL7s3ijwWHpZAflKn0yH/utvyfaoG5ub9zxvL60pCCUhLR4HCK
3u6JpmNQt5e3a6iTAbdfl7zP84+VOECBNhlSvzPkjMW1Qwu9nQ4AVO8/qzmY9Qru
JDGYGPQ2TIjeGNauQqWuZuQ7oGtnHzSEgTn5SykwaLBrVEqd4cFaej6R6VOrh/N9
pffTQP20ZrUr6f6c9jmvPx6XBS0YpB+kveIlxGj+ebCkmVlJwsJEJuJlt0vqOdln
V1s06k5Oi378BtnLuw6nTtIv34lnTt+yHyi6nvl2aeOnjOsZ29vB4QIzvPYK/LQ4
xXxc1tjVMN4ObY32BTP+ENGepIyNmICxeICs8t1xAGZ205qiujA4cWdpLkdDU3ku
Bst/OHqpGObIf1CiTn/qaDF4Z3j5nTRBJHAUwlLXOSjoyjaJ2qTik5lxHx9teHc4
pK/6SRtHkHnCM60xcgp3JdsdIVEudAv68+ogZ7pE+WRp7WByIoyxwYxXImeZ26ID
RUeH1IvUAtyDzb2r4CWq8G0qngi+p7cDZ9uqcdHv4KS7A8wkwJNuLLX+ET1NlOmq
/WyyMMMPdBzkULT6coUdoD1qKHIcsjr45AoqGvemQqFqg0E96DNG4kK0QHatwwCQ
xSuLPitq+NIUSpL/z03+21FK/ikGBFeeaQh056+5Bmsd0msXlQ00QeAcZ4Sw3Uq2
k+3ctfv77EA6D4OlKFLAzaHDj1R64aRoI9dzi99ZXCFuFD6nvn3WKL7o2y3TrTJ0
wcgHTsA00NvX8gwtl3ha4rapX/syBTX5Pa4UHa2ORfzS2tkUk6yudshjzR6O5C0L
9bQIntWXzW+i8rThgIgM/JYqgOAm2GkATA6QIL5IKih8U3cY+KVThdOd7bs8o7fA
z6dvdXeSqis1dK6U+/Obt7i7MkC1wy8Pah8fyKz6ksDK3lLAt5dJdhuGucbLPAoJ
39PuA5asuwlG72JytZMjnt3vxVWHolczjHZvM8XQwnAOccnul+nByxNI/aZbdyPD
agNcIyQjBqTpi2wL7GqLMISP2XAcTnYwZavz7JVUpS+rikIgaMwxPfZYiwLqBQFE
HcXGAXnjrwrI56LMREiO/DjnD5/IBVc8Q1Sn5smtNxwnjEhWmonoYaqODFV/sxGM
GC0NkDMU49TY35aCLAwuULH9wM5yPhmW9npcbAmOQidVG0QAqGabMCQUD8APfbKI
EXwuL6uMLt2wXUwJ9UafdvNka+7Wcwa5rmUIJfgD45QI0SN8Kb7Nu4/1hFA81CPi
JlcDBPbd8ZWEpzpV7yCrjrRybfQVTTsPGZh4LUuxAhCGZfpaNwmSTusGQD9WModF
J2kpkch8MuJpN5ngjiv//lFricRrfDw6gLkSQaLIEq47YPLANcboGbSHGhHjsj+1
+zaDLciKRfawC2wN/Ny/emK5PrvFezoMvf3bnIBev8AaFE+sg8a+IjuJBkzqzdXt
8FaUZ13BLH1IQO2BtXkkDQPugONoLvojhHZnqYqDLWtk7U+7aPRGezfqQH86TEIA
se/qikU/f1EEiGzjenF6IErnH3YjzOoPeav28iuhAnP+mkucvEhWoa3XlMTcOnHd
1b74CPhuCrfa6+XkFQxhXTrYbMJgUZlfZAUZWHi0VU1k0yNs23aB0QzTCZO/s/xg
4sYzhFnSxLQ7hqp9Ud+O6wkoc9u8rPEAennCSAQQXAG66/sV27sI5ZN/92MoNYn5
nBAs61/vAQqTfXnkjdan746+291xJfIKvcRlrQIULIaaEZxiizs1YwP/yeoyqPEm
28uSO4DjkJKye2Jy035Z7bRvt0Ni1/xZBho8UxGecNk6GdN6iAt+hT32kG1DujlL
QaI1AbxYHW8QfgiPWUZuKmvbyP80xIT2ZpJ7fY7T7UyuxThMr0/2CGMEvioG14mM
ldhWcKyROMy4OsBCI3+gVNZXNj276FSOoZipp4+9u60eo+mJuwd1Js2raQlNLZeT
3eGfdLRwLY071B5ur2YDb4tH7b9siieiBQ7syLdTscUZs/hfV0zsBytQJ7rbkXPQ
ehUSqcs3YU/4Kjqk4MinWb32CJBzzhbrfGLKL06CiE94hsUvksoz59ySkXEiqnQZ
CVfbNwNw4GF1Y2pX7DvhHjFbLx4+3TeX0lXCR60zKmBK5+1jFfJWShiJSKxLxDUR
p1YMSyIsWOeAqkiaciIukd4VY/MayPtHoB4N3xAlnCzME5+cmw2rl/UriBLHW2Rq
39o7Lj4S8VZM6HYRJqBTzlHRzpA75rSaGUn8UWZrLk8F2KAihXFaCVAve83HttDH
wiq+KLatT6CpbArEDWJcIMM31IhihLOegWFuxwy/YCk90z7ilqIskihKBQSmjk3f
Bh3fVC35rSxU4pvHnekS0gJh7PY/FxC8mFBskN9misUikdyFZYCUUDhjesBw73Fy
NFePGwSuSrs51QjZs8mF8R7dCPmZbBrKwRnPcGoPZcAVJBam/H5JiDRIr5Ygc9f8
/C+3DNuNGxyEF983hXVARowJ2eyJLAfgZE0lPl6vIXgLzUsmbrLIEmWziWjWxJqc
jxNtZrFOI0uHFrHqFSInh6dCy+j9y0/BNXa9pnTtbuiDl7q2Yz9mrKGcvWnTQuA+
2YOid/23qAgmktsyAByXchBFY214v9/HPXUF7CW0SWxH4sZJcumKz49vK+ho/P4K
vVqh8tgtJGScMQOkeWWbUR282VGly7eHOEvFAmIzHT2wlV2oxhzMBglNW8RM7b3o
kD08rNUWwSFJrxcaQRVmsghr/v6d6fQmmXOhQDbLqCCfGbAkgOaPzIW0v+T0GXjl
Ne2j37WJsy6P9HZitOTamxbmaD6ah4gbPmtsRd3AC36CnlU2GVLwEBfI7CT6XIZb
L1JihCn+t+kpLbq5C8lzMNTB8zpxbg6cLNC0T1ErQoYNSy+rU6RxteEb9Ku8cv5C
CFBdowkubNKZl0To3JpCfWe5wZKMU9IgbuN7WGUT/dGmRmrRb1y8YFVPDcjnjrnP
lau0ymtpnrlpIC9S9aZAK1q6ST/Os1IAEhCStRFardvROOD8grL3erv6qKtbiHni
apIafgYYMyBUjlEcOtzrB1jVoI3fLVAtArLPvz4XdcSckiKx1GY/8Amg/h1h9OOH
0shY7YbWdhk7l0lEkl5imtpi4TM0Fj09obC69Tjj101qULLM2kevT1SRErff9r1M
mrFxphgFXG6n+qGky7HJs/p3fSh9b/ozczbW0M9qfWjyxWKxsmwLuPSJ5JnqyEF7
6MHKRgqtfNAgZKUaOnOTX/6UjRbuzIHNHrR468/IA7JHuh2Z87gPi8RhOulV+cnz
ZXaK/xPL8j7celWJtJ8/HlkMG36yNDXGVpDuQdyz3M0eKUE98A7fYCDBnG63cPUV
Rz4+k/7j+5N/GpQnDLHBi8o0s5ZH6EjJrsbQHdktihEIKNfOV/kuX051gbEEzbuM
iHN9QU7/nFQcd/IqOX3E/E7kkJ7//XfzAuZZyq/zGwO4VXWALErcM1YvcA1ttW7a
OTuEEtzTejMoha3I20cwUIAoi8k3y1M9f0XGEChK0X912HsjmGYAQVXpuRy6JqqE
Xmj6FSmcT7s+4mK/c2YuuM92deKSFGGBgjMHtJXjIUm1zR4zf9WvF5WPcmMOsGMu
4+S9p8kjl3YJq2en5aFaaucGe6IaVJqau7POAHqiWe0jq9B7OxokBUZu+Vz4ePNg
Iza1Vq5KJVB6jtHSoBDlXsRecmMukR/EhjFjKXb8C698RWn4AjoM6G0AxhqIvsW8
2Gy4Y30yGsO0PdUIwi3yRbFcLNfMsAJnpqVGEu7FlhV1Pzj2yrhvqlg3W3Gj6uMZ
+MYITk2KTo6n/O8mJA1yFbWnAzZe0cs52FIu6mcwGAEdkrY3tltmle67Tk+hxCJz
CWT5cTBGoJGm1zO31FcrCRx7gdoq/tqGLIczPg587zIF7eo66xaPC+rnKRmgoYU+
GsuP1bB7WtJ/E5YOisZ6Myk8OMKpTmRE2ccOSQkKf+ES7uNgFa3km+7jpQEacTw/
V06hSsXtVTGRRi7+VeB2n3OPs1mRS75JjR+01cXr1wmUmowa3oSr3hV31jQT8iBS
l875qJoBKEpwh/5MoiYa/v25RaUJAAqMGxcCmP3hX2JjtdVKnierqr11aSZpsBOV
QqKiHDY4xR0RauQd9M7/PB3VU7t7IcxPsV7SyzTPyt7BuIUkO74ouj8uGN2iQd96
WJR6rJJGIv88cti6pXQftJx7AaHVfzbKJ7SfVth9t6eDQDVOqHMMPbcH7YP0Il0G
3hpSKnzYtOrXnMYdQMANnDcUu5Bzi4yERrhj/BO5ZQJfUP+Jdl+Za89FokwTvjRw
C2ev4TGnntHcYNkG/sBxBuHxkFx3hy4PtHnERPLheCOX/OcrF29uXlLFBnfkhATI
n++TchmJUf9Pdh/vJ+TW2FOWVO+UrJZpx01OayKUXMnKr22HrrX9EtQ4O7WwHwn5
Xpi5pIkOjR21c2KPz25lnJ6/TxNezlKlzdlsIm4Zxgpgnl7BRbfwxSS9QavF8IVT
4c9cpZ0y9BwLZi6ez+RcGlChY82zFJVCcA0DDOHqwMlQuEENWK+S093o9FteTkME
WSb1N+Ee8iLotT16/OKQ6BQU/4xVkF52hFZhgrlk5csE3MxjglT5WMkVpqwoz9wP
hnSzU8jLFLrn7OgN2T20gYIXyN/v34VUT3kqdY5DyJCv6HeE5cbit0r3VKgDCLVQ
kpfuJQ+cBAPG6sgwKsKrc5cOF8uzvQwY5bX0rA8zzQ/tsW2n76Tfsj6zmn+eWkHt
ijSAjxGi/f7chD3k/krHVPFjqBvNKRUOZYzbzHdQQIXE64punYjkhPl/MPPpJ0Qy
Uob1oeeOZx6z8p2lqziXIMea3Mc60f2oMyf3cQF+zHmjm8IgY2Edan1eqrw6A7zb
gt1tYn6V4XF7uMVA+E4BwluMgqehayUXRPNWka0R6NGrltzlfVh7L2GI81/aQT4X
r9CMQe/rU4qad2m+KnE1KRwCuP9uwuaL8BCDgehVliBj3LQA5ztfnWoIudzfutD7
QrCOrJyNOA6fh7vfGw0FjUGRChpSwAztmrheYTlTbtPmbA1UEnHj4znFrIcV44jC
/crpcntsoi7MpTWOYD7+j+BszxVJ+rB/58pMo11TH/9jIes7ktr1xDw9+TvbqgZb
MQrCsCb/O6RWZW4jNjJs4KLoongFkFO/Wm3ErUfqQ4gGK4b4mbbEkwy/h3O7n3HF
aIccRfkWn+DhL77ITX10KCW8psauGtIk+G4Xhu0mLLYKVBZ07hj5r/7i3bXj5cAX
Q3umDa8eQ250aS/sU84mTQQQgg/Gx87KX51CcwRXWcSUp5d6gJOGf6X2b3jCXXwJ
4iRcCFozXInYuNBimqWP1N/qXu1EdDtsChcP6m/uqG6/H/Xb8zgzHIMPhiC7PaBf
YhiueMFJd0jrWfnWcWvM+HxoCvagw61R91hADZElP1IABIbpqFa4Fvn+vNmhlBmt
bDUJnd8WpkX3Ktb9sTzVEGGQ9vmIogMUtHeQ7kE/ORtBFyKAI0CGC8LsJT4AxtbD
rmdID/vkiNcPrjAjG+tFC4BhdPUaq+BgtermQp2p7ckACN3L843p4UiOUam5vBrk
BQQ4CzpyQflm4nA2Uwk2o4n38jIXUHSyrKv/F4JuRi/fRIA0gBSWFf50amjHAC6o
AUjWUIyENGIHButj73gglJMOkB4ZM64HdkNr9gsS8YT0dC3yo7GQvlr4CgQqA7fH
uf2RG8i9TBF7iniuooYsFLb2oseGJIk45u/3YFwCRnwG3G0V+0OTErIl3MxfLqqV
vLGm5evq8iooiuTmFEPrxxOrFilXNYpBduf/a+MHnxe2JH4/3YaCcmUgfBe+y2vn
n5rKzc09v9VXUNs9bF9q1IvVPUKNDHm4E8S8tWJPe4AVC6rfgdwIb204wNI0lmoG
HG1YTAmuqL0Kh7tqAulCqyGqjcA5/mPmp1SYJ1qxDLfqc2HdODSLbPhy24ZX/V6Q
22H+bPHpuq/7Nm37fxBq2V9thHLcyHOrNicGGrnwC9kstxwA8NeeCUwwOCkqcCh9
OUTF00n3kbVnjUZIiChdi+tRg+rioItvJDsHyHFYy3aqfIKFsA7BPgQb1I/keBj8
8HgqzVjairdVMWklQINoArV6Hntx0q2IXUHFmXmfqy0YDpg+TLvXb3EA8/CZLbvf
avlRZGDRmygkGSW7V0P6cpda6ZqbXhP+VcV+2XcsD5ly4xyU7tF+yx1P8h/Q34Ew
ZzFbgjTusuyv7jfuE4qDvdiHSwuMLJq2Kj+Vunc6arhJIy2BV1alRgY24Mrd/DJN
Bn/9NjccAZPipstwLBtLaQ25ufKAIviGIz2PycCKZfKQPAfa0ShkCTF3j2EUhI0l
wJ4droIXPqN0ZdBeDGeHjLq5Y+c+gtk/l8SiJ3H4LaOE3tow3WkEbExaOAC8RrVn
Rj4uLTXGANbQd+mDWAiQXAiL09+5ogtLv2npELlyjS800iBJDtKyaDU74pr6pZX+
Kr/jwPA1SsBrr9DOUwQdAttlor175P9/QjQGXhY0loVzhL74xHFlunwLsj4AIKAF
CnlkhH5I6yb4Buv4UDohAkKb8zxBnk4w7P9k6qlaSv98KH6Hun3hQcM6Vd0V0pjd
WENUvflxBsapuTFTDtCbiRDTtsnZve+WmTyLkhXvZZnMcY+0Q9bVbGgOxXaTR1fI
VN9Fe8R7k+z2Dho1vOVC6rjM9itQCnjGwijyMVSg2iCSL1gjFQ19Hy/LwT34tOMI
KlD9ofwmidCLNrezNvqi4n/v+Vg1cWwe9fkoudmA3qHJ3r6SJqIuNj3YFmX3RbEb
gHunwEjUz4VjKIY7hElpwwnZmXNhZlUbceJJRhQ4rnodoOWs9M34PjYkUCOgbgHh
B/jMf8rAIk4RhJ45p868H1UddZpfGI2o/Rg0N/qMRCv5iWZptI4J0+IJs3GqmY+2
mAD/65jPO2ZMhTvf3YBTuPvM+yUVVOkxwMZ9zmGnP/PkfX/m6AzlpdtUmLPSpfLO
pkXKZMU8p4UdvIcUUhFonQ8xVoUUlSwUtKoUSgdgZhF9peHB6dnLYoc8BzoX8GUj
RUTeshEZbJqgkvsBltEDX1cD3Dh5ck+FoClWY4me5tRuoA2iHectQ8UWdmG7jZ+I
uZE1YsLZQRNKtjlDzwdTHYYwIfs0J+zKTESqH/mQ7H2J/38b9Q6xh9bXizKPYKO1
WKt+aUSUfZJHifydOIiXMjCqIGTx6KRJNGmJj7U2BoAW6v1/Ts385lnNogAZ0pq+
+O8ZlWIwk6he6x9Mk35XceikLTgnTFi7w9qlHbiyQJ5t1/5DPV8DMIWygH8EHlgJ
uZr6b6TsCh9PNDcAevgFfgsYTihWQiXHIfCPDLXAow3dLht5CZ0TinxccgKhVI4l
IyW7vtyeRRvMm7TK8iO857htIVTTL+0VFUlZa9tcEi18lqJp+uBE+5Si+V4GVDV/
THES0j4rHdOsF2X5HY6uev8XGWHqSsarzRDuWfPtpn7/5102mbFTg2u2IgAZwXVB
9ARKvW5UEXLbIx7tH77xrNxBt6umc9EDjQJ/PD43fq3XxsaQZ73cY62FJNAJaZZE
uqVlsp2NgMkWLTDP2TkAMlsh8BnKBWZ6qfImqA/ywZIKV+pRpdTRhqbClLaTBfPK
pEAOqkhdMduZZ698f1uhBxMCzgCXT80jpmHVHOH2gHuXO2hEhkp4oH6ShPADEdcl
9ZxM3pF/cgzT63wVEIr0srNWSY2IpDDeBT9h3Pxzjy8hVz/P7k44sJOJMtZdQtaS
iqd70kqskB8kFiG5hbzP8pFhffHcUOxpendwUfQ2AeKn1J5imBlNl/5x3gTN54hQ
itIRFKr5D0qGbWDKdZkVG7L8rIFUNM2wkntAxNN31WNFshXenHNWqi4k194t7RnN
amcjVHgLCv2mqOPmEMMIIDGBdvOHdDQSP8hHw45NoK2BNzhLS3mzKOf/aHueTWSr
R0Hjlc5dX/0A9gTH8kw74fNxtnlWfDAvBAlXLDI+8MaHnFwy2ZwfGiigWfnqLFfD
i49aUh3mBOz6mSaEJwWJdONTmT3XdF+cxDpG1mHaGXaOpD5FXwbtqRog+L9dTnNk
/RoiiwaGJU49aQZ6v71slcZqCRY1TpOVhrpRX0zrIU8vbm+xTYcIVJEn3+yj1OY9
vC6wW2zLOR41DjUGDFOcbXbHp72u3xEkmtgzmbQXeGdybfZtpifvCtDn805YcDOl
6SHOyvvtPcvUBhfSFsy1XAYabllqYSyGZYgoPsVIxsM9VwrJsOEapYCG5UbmGv6J
EGSc/MHb4adQNfv5YmRS9e5t86iuNoiWw3bOy/osxaDU1ITmo6E/z/6WTVv1wcN+
OVA65vliSse8btx0ivsReRX8V0gAJ9VmscPCqJ6o9xil0TyWv3jG3zgfZrwmkDFi
msg64IYN26efhd+hstFycHz8eRRnZi68sIVMDLEraWRNdEGOkIDDUVyB6aDlWHb4
3vVHmBCToOxH9xUrQDNFRuZFSWpP2RfRlarMIpMrLRuZsAvY5i/JAWHY6FIurP91
v9wDD0OfBhe4nTm7FJmVLNqz52Td/SqUEw8IEI66lmiw8bKfkMMnMqQhvHmsLXVn
XUe5f39NePuVG9stY4NTLSJAG7ujvVAeQAeZu9sFTHSM+PaYNjNjcf7L7Undp+jo
jw/3yRqzuHT6uxSjFh/X/dRPKqGJUaUexzXo4sLbSW4DM/qu2aAU4/4yJEQR5AFS
3ZXfDW9lSdnkJwDfxgh1Rf4GTUPiaF8Cewji5yu4/rq8hwXqwGOYBd8AWszAmf3a
rUiqyP0WtNjHZpabWkGt1ekiTWnXDi2mSvbiAnXAH2c5UXf1loWAVJAasDJcan9S
oebIMs65dRWbJsK5KNvhA/tY0yHchsHcJlHWIOiWMC1E5VB1K6wXItIAssImA+eQ
z91Gze+3R53T9FgP6UoGhI8N3DJw3S/7WverCERQxF1bXBRAf3Iw9lVIjgs4bKsk
Bho+YWTEMuDc4bUk3vXVVoUYvrS9ycBYB2+wAjDQ3qVoYnZyh3tQWwXjHCsNjAW+
NeNiljUjf2iUhgAgF4FjIGyFU4XMXJBnzQukzs/mgwck3BHCpleSAQpDauCYC9dt
/o4MUkRMvlEtExAQEYcwDOOwq1afjCfAvX8ocerpgsKVZ0zgADpfPLG2Pa34P5//
goN1EImXNK2uZ2iVpNk4NByakk/Wbtcd7Hy2n4AR+T2eTPYtHYgC1BNxj4IZO2xh
k4DINc4Qw6jfvGHGWdb49s4F7PGbauczQ+skQLNVVlpuGu2DfecAjAGIHD5+TBMz
wnBGb1YEudGIIfEVCeGS3Ep1I83Ws79cpO+cN5Z8EGdpTsqE+4wMVfYYdKEt/xEN
5ewSniYDktbXbbKbx2pNJKu0UjWTsJOZQL9ubWZea3dE1cowynHwSPU3SxQ2zzKh
aRC1zTIgUJwMh1oPCV0yUaPpDV1ZObPZBoE6a2oHKzgVKndxwguLFk4kKxuMJij9
iXdi8l92Gf7ecuS626PniHrTqHeL+DjUNokzgPxDQrqFUYBuTZ3kxePA4e53HEwv
RGUCniOIB1W31WL7ghSC6+wUnszacfU+1WR4NHG6tlpaTEEnZpXp2X0JJw1t03MI
PEbdOB4RC5MwzNw6bR6/g02ce3DW3WY6GHk04dMzJME1DoSW3/bykpHMJSG8JtJX
s4n7keTiESGIw8VAFLn4f6uXE1JVKRs+Mt78fBOdcffTpqUxiY92aLvAKgdU55lr
91UdNspgsv9eb3M+zdldQGuMmUUpir29l1C/YMtlSUvzO58p7wo0nlNmUME/LC/p
nxhWpNAWGe/DlIIvjUfvXJxxuG+y/jbaRNAz20ljABn/Oo7wBmZa9MKdsjg64HEa
AkirhR52Z9dZrI5qWg5WWJIFrWk08KSjF45JtK086cJFsOdXwUQTabiVCb339sP1
P7q8u4Oo83Wt2dtcgRx52JfaBafDClN9D/XWvHm315+DXpzJTqgvjcpefrXAEWhe
aZPIMDv3L3pULVPdCZqqaiXCO8XaqH70wYR/ms6tfFeM4l/+eIEiB7yVjKSGkWTt
LR7KUDcMDraeqWVGOGQbflvh3B/FneUcyUqqlIMqTLWpvi+cQaS5jwcj7OI0xV5C
9jlfAIuM5a/tOymrdOQWv+sSU44ys87YOjYqtkC+4d+qYn3Q/lmOXU+nk0WrYpyp
GghC4KiKOBSMkzWAY65yPIQoLHkFWjT4tONRfqELG3E3SeX0NdIHOTExnL0PG/JP
fd6sq30dkkUJ3SQqTxROvMNibsX6YHNtqBcmGZ/iHhZKXwiD+dHwDuwnCbE/YZwn
1GekL9Ne2bipjgppLY/EdjQNzqV4Lzm8WDt+3pAZmK6pV5EG1gFyG7D7wt6DDq6o
zG9ztIhddw4n8zSHJupl0YW/kJTD8HoSj74FwO9nS+viJYuWvQdkp/Ouleg3SoHD
Ne8+tX3/haXk4Azcvuaq4jtn3BCMn5dWagV0tR9S/O92aDWR7GWZhSCAbzLNjGbr
GINg1j5tXJVKWGai694JEIQj+V6Jd+AI/iOSP2x0C5mRNTxyemZ3eo7L8Y/mSzcp
tSPA3uD3br/OBKW7jR0YWA+il04CUA2p7AWxWMsOiEvhZQnP6APzTOIWZXjoTQwN
YzJnS+LGWlrwFBCf4MUcEHtRwExyONp2LfutX1WTqKuFNfdHjTJOiqLBN9l2T34X
AR10KlLcZDpzHvYfhgqPAT8lkWxopARp4Ec05/TtZIuvRWBXqvxGd2OQ5YOfsK99
RHNswTelpj/DuxnngTEdlPDtXqntdKDiSwYzrq8waHl0b3smaSDl7NombP1uJ7pD
N/85ed/akdZUNLEQ+57AGqk5Q2diOlR1c8ICxs4LweCFF9azIkIymOxEO4+tviel
5J99gedraNR+p5HTXcUsexLJVC7HoUfEdKiE09sINRYSJKxQ+WBQbWITyiQDyT98
6zfjbXeIsJnH0cPZl6VXhN7CefJz92bp2GcZ94qujT4DPCPSSa1pG6AIxUe4ve3T
o4gPYNf8gAELIVaOa5ShDPl2uzjj3DqC6TPg3mXpPk+UV5Rdb9mdLI336SIVeSBv
HS9NEkmEeSuqfLR6KjJahM5GOvbxenOMk8u8OSuPg0GeP9N52Komgu6VdGPYFH3p
OKZnIYxcq20IfGdPhCaC/V/mbqk3epBsO58P3w0lClc1nBp1dKdh/EV7Wv3kq5Y3
FlOCeX1sK7ZReHhqJF+6QL4vulbxEVJyWqQhqFhjBv3oWU4w8FChqCE0Zo1lkNNA
kFf/OZQEH2ySlip9GxU5u4OEXo/t8q+SlKG2RmnNodU7dYWCbYPV3ZQ9qICpjJOr
Jw7f/1KVCTBH3r58gt8M3zzIt6AhtCotHFGvi3eH5pLX1H/EeplodzE3WX90iGee
uZ9XKRbpN/x4TTWBRGZ35dW+QaWIkAx/G5+3N7ExDmDxWVYK6gDwQp6/f0rJfOnE
4NwAgqH9TXYgl0Lol26aP0EvRv9ytpFn79D5zFq2tZ9r+x6DI+wvIdSu//dfSJ9a
pCbB7VpvmZEUtlMukZFgPITBt7kxNLpKMt3bXW/hmk90S9g7dPKJuypzMdMj4nkH
gvRTJ0BV/JxgdiEPXC3/A2h2nXdtUwSgi/vehi50CLlka8mCwzvO6Q04jjIQ7oM3
dfrEOxR8bs2SCDXBpykFmhmLda04+9IXqqDqj4Se0fweUKRa37sSc2yeun+szDjQ
DoNu11jCSUZMmV/hiGnYWMkXyj1ggAaL6PhEQFL2JEVDrFNMJC60LuEC7F0T6oCB
FJvcILAvHj21aUjAjz4IYHZ45J8w8kdL7lZDzIxMNF4/SdALbRdpiknnE+xtzxUj
ntnP6uEzbEJv95ksPHGJlzY2n7liE7ixDSr3sf+dMG/oxnLrySuqNWKhq2XRxIfI
7+fvKgXMTO4k3mq5UBOOFQPESv3mH62ZAus7GtacCma9wBw74UCppjr7EM7Pr2+G
86KHOfGce8TDCMfwTTJ1f/5UQNBld2rYpJqr79LNo7bzRBKPl1vQYFk2t8GIb1g3
CLuGHSJqVKWZ6fdfnPT8bz5zJ4SuYcHVL9mtSBx85oYK9JikUYo9/xfXZLOej9Wr
XvyUaxO415Eo2kOtuKwrN4BvKiT8ZRjze7HwiApa6UVSmHnS9jjGovlCBrUxAgrX
IZQl6bAO1QLjJZVEiq683lFdz2CUd0zTGKQIJwOjqQtmJtgI96YosQJ3nMwQTqj2
x7AzuE2NTHXvDW/zqkXRW6siBhLuJJyxk9qO552EInPNUSDCvTsLxkDbIQ44I3sU
19D2mtxvsZcN1W88loTDCxMcCPR++suRLLiZV0jx33f52juM94PJqDZx/Y4qX/J0
PWp1xhCxk9+QtNymG/n+oBzVGTaw9tn/t7ixKjg2/EfOgH8VMKO6s90iMlAyjhid
RX9v0lqUK0IV9yL9bGq018SmZcIToKvrcoeGYsFm5ydFlkbXsWR9dNLnxXj4ZYkf
y6vkxHIY6v4Bk8WnM8YsNWvvndJGGgA8v2szgtONFQpUV91kOPv1FW+g4TtawO+X
1IUjjbUkRozwa9sTDe5Az4YFxMP2TGnTjdUq5EYzDPHjU8ixTVcBocZGoo2WZ6BE
X69pwpd40c0qBFrZliqWA4a4F+/a76iY/0mJYOjq4S8FSOgGj97e0p2HYkW+Smzs
OexCHY4qy6IFOZppRi9wY0zAKatQz54ztXomgHp7WQ9PQBHQ9iirXuZEFNNH00XV
d3/A1FgGESc/CcrwewQIe0ZXEurX/xWsO0rS4PL+aQwGhqKz5fKExxuR1jcSOMG0
a4gCTsoT8EnT2stOpCncs+TVpEKX0pPwmEsjiaO1IL0o8uvWDdUGE7jp6FMbdRbH
gJMeSYjfdFrSON9jPVjNEdsHqXebz3gbLfEUh+VVKTk0Vl1mEuhQv2khjUe0j8zf
rFOrhUeGnvVAld2JhY8d3xbBFJ++dZoVYPeR9hK/rIw437Es8BRrTWWxlCf/MZtQ
OTqvp+XojBaJ9TXXKXjBJRj83LQkLRnqBl8W67L+HlaELSysopciwdzY9Y5R6549
rS5x8bP+2VVszPhXMYTwownO2IegFlsDQxA8YAmRCEw19ciE8OJguAFNMji/07Op
alaTRei/1DKqyek7rDl/3STvNoPCk6ukx3WuFaj+/lXDaHJnZNOl0dpy9yvF14nP
ZhE0ENXroMytB2UWPNMNOaS7sOkfeLQzB+C/+aanNYrlomy+xSSObOvtGnvCkDXH
ZZRzeKhRvyhijuEOA+lBjbekIZK+xbyTAgEqW4hdjIMRCQcqaa/41S7OGr+AkZmH
e5dFMQAl0JPjBIOTHJ+QWHRrEoolDosn8l7Q9g1axvWFwf4zx/qwqOg7IUoilnrx
faJqxlAMxAcQc9mwoygJ92KrqHrmd7RYw1dH0avdKfgtdXzYgMDbepgI8PtOaQQd
wsIfMOrhr2behXszpS65EDkQ6lFcGQWJwR91FkaW3JAVni9ByJ8YJlfBRAMfRcop
jc1CpDKVPkZjQ4SnXlBH6ukAijtrMb9iE3xIqYH2g+0EUJubufGCmErWNVkFEHys
bREH1xoM9GYU6v8w6DOunqfkaFOE+OigQl4EKRK8RisjFMP31PRIffZ8nEnn+JuE
ymIcyRzcCtldNFPNHPMnI6v5dS+br8QnVCD8bCKYGA0aOZ7//undQ1cRu/84F0X6
o1m+lVSRgK26d/qWu14QZI/1dA9AP4Dz9OYVHxcVTJEIaQFDPebmGCxy++YzqT3K
+x6GaAYJN1QY8XbC2t/QqNGJ4dW/tAbW2jE+rGDi4FYNr+EHaaG5K/efp7M82fvP
mKLER56w2fWova2JRQY0PInts+jV93aXd+khBOL5nTcRgUAIxWP/q2kF0frAqT8a
0xnpz0YjaPs3yFiZd0dNywJbdyvET8ClyS1zwEwy7jygOAgxsMkvOotzpD6lNN97
wDh28/YlCpsghUI/KSUNgSm6+kvKUZwBuatZQugwaeRnYahcrsXtpzAJisXThyoy
wyRv0rOakQygd52fwNct4+03sRn8HbUkUm7zbvLl2tz+NCQRze42wkR5LgZ+hKdb
ksN3ZNGBRix46WQGSM8SEMZnbQNlebevvCnME1klFEKH7xfSbMUIEk+CM9LftA8w
M1ZilyM6uUJkuZAjqHn6EW6Y1tWbAvaXpytun4ztOEOLC3UML/78Tfxr0G8T++0z
g0Fr5vPEeUy+I1XBpC5x7n7ZqQm0Kro5cMxAVcw10dF7Og3UdqSANwdJGN8U+esM
e7G473v+zRgNzLtY+y7C2euadozuD4/JUv5eeE9ut7Y8H0sExZ7z3zEQiWymToSt
wyW/153kP6X/OV68gr2OMtWrulMeOeXqjiQrPzzdPgQn1a4py5LIiQp8/iB06GIM
oF/f7XlFqh0XUnSk0uB0Pc1TbxlnGwQsGqojgLr/jpfKlWVn0YSA+ZciQSvPvAjz
BTYG1LKLw4Bek/B6mFdgr8qSa9aWzc3sZDsIfZNLG4fhSITvt3LvJG+LO61eHe7m
CzUVK37enFX873DADtBnEhdeJ7ktKNxPzLsE0XUIfMfnrQP5aSS+ILL3WAmIGavl
+6pBnNa7GkJcMsfdb4ugzrg/ryWKr7ecCtH5tgouOVHEYS7NAQlkxyh4KIuf6rBS
TZUXAqOreD3bwKdMkqvLkBgLNuHjw7KkgbfteTv1C1JyS54JUc69wRWTW8KvNnrZ
Ruzr009KSFZXx9nIIDUuT3NintbbRk6qDG9equNOku8ZQK8+64N4DeS+QHcAeYQH
dmEkBYHXpdtD/lX2Z4QsOnhqWEX7qXOO+CgykhPy4ZAI/J90yUOZIOdHJRLDPYEY
yP/qJ1RCr9DXaYDoBv177Xqft2Z1l6lgrSuYr9aOOpumFMySLYyDBxL05jmD4kP/
/8sm2c8JST4IDbG2kJolwc5zMm/ye6ulYNwZ02TcbIX0+JwIFLoFO4ynQvQ7/X+l
qf1jBaZcR1l/suqfoFErsb5EDdjNVxne1nkse8d+rJUCgnYlqz5MfD8B+AHE6W4G
1HJnxnA1enwR07p+qYCxOJx3l2/h3kSWPaxWCiDjL+lvJriig31Y10sJBn2Rk3iH
Ptz5hltCKQBlSgP6N2A2Gy7EtdFAbt7L6kkWvw91R3B5epHAW4YHkIAq21XBkpzl
w4SwIdQXOW3qpEjuBLlQCXNAPIdVtHScmp3Rnwnb/6AZTFFeKoy3/RJOTKMsjCLq
pyPXXJmwCum24Rpbc2jP+ORdhruAsGzff/l1LOZyHMleg+7fFEg08RBF9lD2vjUW
dXPZmsq7NyaRkSuDCO4PSUskrIR1tPzZ/FyFLFcXntcpDWHlniUj3T9vumJEkJFg
WAbAwiGLZ5UgN5e0dE6b3CFMH6JPsRgfQJtzcmZbN0ogodX4BYuJjrm1IPSs41fm
qxaG6iBlx+ElerWTtAsQ2/+Refwk0xvlWVgVR2FDWCoQZaB/olarJscTDr5BqKlB
GVrqmH4gn9f/XmBbgjSA68CxbGmTpMY5rPA3LZE4P6SfzhFT+QJvpQlmykWA3x6b
TXFqrBN5B2GvdwhxGRa01RGCtXGnl9flDtqUFy8UHAQ1CgBentsKwq+vzlixhaQx
4oC7Jj+dRvjNvk/Dd192aneTQ/2ogFNAFXZD4xsovIGgvMt6BZ99ES5KQ7jluPv/
aKcVQzELPX9spQDk5p2aMd4Lo5JMezYZTMSv8Y4sok/NPI4InCcSTMyeI37Ffzit
vNZzo0yNJ/beIGYUchfDjBOWLPEJp8Y8j7sE8Y454q7bg1fN08UkyfVSEEx6wu3G
0Gx3mFfEmWLr0dGmI7NSclZsOr+EPyQ2BYyRXcxaURfqNeiKkxCHz/t4WaD0m0OH
8ef2DIir7h5bcAc59Z6/CK7IcF2OkeUhkKWc5qFMRR7fFqFO6jYUKe3QrwQkAoKQ
QBQwqKmBKyblejHLgODevyhUmwUaz2z6j35cyWvExc89v0mCB//hq1kpRskXFtsj
k3dSVMg1CcJYcYE+Se43jwOTMrgqKxzIdD2SFE1ew/4jw+koXfqB86hVTWdTAfoG
XCosTz8HDX574dsn/1B/e330s21xOq55OM7xqZkY5O8RPScRhDUVTz1q+g4Fowyl
xhC3rjcjrGkXZjA/NiAI8BMWQfRimWilOS7ofEqMJAk0ftbj66WZf2R0pJVVSQdK
y56/AC8/KG4IPAEV7z4Cb2bmYIWDEHb2/k93Gf4J/T1X1C/x+ZicPGr9+YnJ57lo
Xtd321Mi8aLyhW+MkDDCLaovaSmPh+REKLWOJdFWMlSyi24lRzyKi8JTEZ6OYgHm
EWVexjpOUlBxiwSEy5nWl5VYZG/HvTee1943jOT6a8O2x+eFgt0wYgRzkXTf0jKE
cgmW4HBWFSIXreDcVJPNALXzL6v8S8ZSoAJ9QLpna5+cJqTvakSom1Zo9qI3UQn5
j+ssfvdgWMlQr1JQVFD0Rz1jNC8n/WZm/s2+8Vo2ciavUIyZCXM95a4Q5L2iaI/q
zDuxYFbAXHeCvohOJXoZcVCHLNRv5W5c6mswGLXGfIJ4oVc3jvo+eGVhMFrr8Ziv
IhEUwa6Mla1gxcH9OMaCHp/lpF48+gnlCqC7+YSjmah94bNQTFHa8zjRRKIbBj+2
FVLjsnGo+DFOj2ygHjQ4FKH693gHk89R2e01v5lCxbRc4is2Iamsz7jHXAFRTsUY
slQ3pB7ifDVjPDi3t8ptw7M+fFDp64YojjbW3SrBDExEKfrZSQDiMkV7FeS3W91R
z4W8aOFRKEyPEPLTpHYxmXyP2K3FOv0U74K+6FLdGUyz+KXbzTWI7YP5RSdMIAIE
2ccmjF5hKLP8UyKvPwVnFn7InR5Q+WhaLid3mX1zHEAPu2k5Lh3awjMXlWhGSZWq
Y2TH2Kdji7E7hMtA8i3f47zUcnd9XIE4Uwj9x128lfo8C6sfT5U+jlMFGr1OXaUc
nkc4zIyfVVyTWzlvrm9QBW7UpUdZ5tVpYkq6iN5wrhqJTeLO3nTMT6sRxwfAFNlT
+rc7ZtLTSN5m+J8+9lliCQ096XUSqbFbQ3uYrqsGnx59qOcONzsHsK5T/TXPHbr/
q9kfB5oW3V3SnkO+WSaMy6CgloixIDpIUj+qudT2wnPRx/OWgCgowMSav253BXwH
iYmbQr+NzVwnkv5Mu/+PjV9+IFV7/YdM7mytONFeHz9wzOfZqMZjFee09lfMk986
rcpyqLcPTsflDf3YpSqn76R2eIceM9w4YyeC3iMaket7cPATbOei6oQ48HWq8Kl6
6oWU4UB41vnPvzkTNkYy/8y4GHlfuSNNvsKKeJljFyWlusd2vzKW4P4l4M1szNDp
u1XtqYfUrtVLAtFQ/wlS3tDUqG/DQBymx6nNYyJhlmIPiNLQ5caRXKcbdiqtpyGi
N+8xFISI5cSMUt3FzYCQjMFda9o0Fz/R4c1h40lrOJuDA4gDS123h1vdrzWWnXlL
1iGCKQOlptrUJj5bONb1jxDEYJbafGJhgH1+stYIA6y+3g8pV9UjZ2xxVBKPx9cO
6YyXPxy4hlpAj/hMKe2aSr50kA17kRM9Ti8D4OrbFkXhazq5sywqr2Ffc6CVYjCi
bJjjEZ9tCURIg+rBL82IMhXJzaoPJ1+9v0ouJBphxmd6sbJfSYqjOcILzUaZ1DUi
4LiG+k2uzm54vx3g5Lx8MJPlB6SPXUrm8qlScbagM6MB+Tmka2UCCf4qtQHBXtiW
+H6hdMc/c+Bq1PBzXkd8kY8xBBSw3p84ZAD93aRSNqlBkkoAkeM86DjWUTDpqXjy
ADkQWptosYg8n6eR2jm8DCDVptvV+Rdj52FU4mi4z9IfmRmOie+oIH+NN4j+3TXm
ufCv8MZRgXMBgbPTD/wVRN1z+zUZwPQoX/i/XUdpGeYz1fGpdGwMHKL2HLKrj8iK
AxaGNCu/FGGtnS+ughniNpYCj5odbt/F/2M8RWCTT5H+s1daoq4RWyxhzaRkY2Fl
v9Tf4bsHxSRkRNCgz7HAm73ZyEA6lN7N+48yXwDbD6bLIOOFYIJf8lcOeQ9zUv/A
SO+PYNnCr6c02Mso4b/aB4WICiH8IGA2DsYLkJDqcc9+JjMRAnbim3E1FQziUqVZ
+b4Z0/uSbQvYMSSnZsx2t8bPkFbyLcOGsZO812KLqvLrivhBUxelodS0ejL8/KW4
eE4p1x4JqFi09U+RHdWiRDhD58g1Hu7QkPogYM3uCFaUVZ5Gvd2SVXZp018ejZ5Z
F7XMoFl6lEP8Ar3ZnG+zz6jnHg5+V4LmVrsd4c7mdGZyDUm5bywNeaq321ReOxOZ
It6cpex7urfO/goosZ0nyJ+t+qm2Y1pTbukAFxfSChSNKtxTStOeIYwgtjFrqDdW
lvSQfYWQcql4+v09/AWatbNgU84DW5Jn6qKHDQYbauKTETzFOlZCsSAOdFQiWzSZ
L5pVjxUJq1adgoUJdFmsmhYQi7k1QQY8/rB6eDZV3m1meF551S1/LkkQCQDmB+u+
06yGvieTyIMzi+9Zr5k0+Mxu1nRDpYOGOknpfeYbwStTqMdf5EbbDGnEWmzg/6av
E55EuCZcXtm4WxILYR1+1l0xNnvuR5mPUhuLOFFlUuTimthvtXctLie928Ta4Cuq
IGopP/c0BpGKPFzKG71O8cfSR9D1b3JoIJwB+ek4/kbRmNRD4xGEqVmQXboIJ+Fd
R9PFENQwkgwl0IU7DiEML5jtgqXIsSCuCDP6NuEOwHLuRe5NilRoHmoFSU7zPN1O
R5y8eHWFNYpaCmZIY8C2ncZdZeyKHDOiflBn9Q8Whc48H/YUVYKsL5ip76UhJLqD
t4vZ0JYwwaHh/Pjo4o1yMnFliMARJH188jgn47ijlhr5QdK72/1Fb60cIT1Qt5aQ
kY7gbGRN2UX74aAmd8YFqpnIlJaWsd51Bb90ICq4ZY3QfKjgh4DbrG2XqIIoQj4u
X4aMQMj4Np9TekSd8VHjlNITUvl6XCDdhx7GSOH2EFojm8Cdj9oFqdnX/T58erXv
n5PuXX4HDmVZtHOnFL3IhHG1545tAOUt0hvj5uHbxEgt6uCAjTXfi9FeQ/2gLJgy
KIHjnOxhQj+1FzcG865+ddUxeQUqp2s+rIjh33M0DpfhcosOPrX566wfLU6j/vqV
+52pBT3QXGBo+ay4WHkML94+7i74IBOF7gTQvLwQLDcrB/NvLaHtLXSyEePRe/ir
JWQP9HbuFA6rlm4J/gVqpeWaLaw2wbSpS14b6fxQOXSNmSo4xaegbMuiWi7dV2t2
ZbmBF4Pcf6i9dLJSgxSASXKs+77yjuqiYwGaSnr431m8I6rVXo64CZRyIIRvasov
B4p+hOJCKOqerEb5pES9eejzyfZ6NPxrmdgtxIqXrxGmc+GLUPtQJhwUpOcvrHbY
ypCEd5OwbtqPu84BsEEGyMhHXfhr1bUkHPyfo1OYELfvInAhB4dojCY3QHc1ZkC9
hAzL65uSHN+2gR6eZGPqpw+vx8GuwOG65tLMu5pQPBWmlZag+tPcIhQ0J59dDzCB
4WEv948hSF6WBrjqhgY2DjBMeCFQP2Odpf0Uq4cM59db/RgRNYpSJENCx3uvc6M7
AMwvNHJSbxbVrO+wvrvdGuKy3upZnhVKaUe4MoqDr8JKJ2TZg313Rm1ixWKCrUvo
PDEpcdpMT+XrJAWJ55pxXBhmwb9OgiueeDyIuKooFc2FxakGwK2l9b190gcbvFVH
ivmki+eKvlCDR11oyDc2nhQkNQ5btq7y9MsJuM1BL3wxkx0zfTuUq9DCzTFpjrBK
9M8YKPJ9azXtahw1QSZN1hsSibRWkZ+kFISqwFkiJYZzDV92CP8BP1zZZ+HN8dfn
XCj8zTg3x3tPfO0K3zOOqF097kGxvnlejJR/fh3HCTvcxdjYhHAZtsYK1UcEh63e
z39gC5RRR7XIR1wwc588a6NJpwrttPAbxflRwbKWokpONxY7vdWc/qkSxpXeMHgB
wj4rTueEbIGq+QEajd9/mV5PY+ohCJFmPg5koLeuzpz1+J2dRroQMYWY5QObXbbD
vtzT7L3yW0DDtT+Q88AieL7azgJnTg2fCRwBHlddi29awFR3cyBoz0Nn/Q0SR9RB
goDKOt6AvTyBzuN0H1kx9nRYnJEDAVtMuKs5gECB2+OvL3vEXNpW3i2qLehONPyR
dJXFPZsluJKO7ggyk84AEIT38eZ0T2GiODCRGeeNmP/43iesD8fymqk43TUjd1nE
2hNr/zkaap7Irg+iv0RJcY298NI+ujSacyzaUTVrIDydrz172hTzsHwj9A1IU0gs
DH8G2OvBSiVC2ikLwG1A0XblC8NN+y8nWbOhu63UtMfLhCU1FIDxjX/mKrmE+ilb
KTbZ9zFQZ6fbE123A70iD4TjNvmS9lKtG4HdAFf08B7XSQR3XMrLd9zGpOabua8+
91VKrtbkUAWLaQrwJIHPkJl0+5KQTVz8TtrTgnY7EW5eE+LOAHVMLUpg2enCPyXv
Sguse/e/qTYCcVgqlqG2mIi/tW3z+GGv//TEN4jKIf/mspCNhvwJJB4OFSTKL3RS
RQiXz+0VS+GzpbO0Z01wX7DBOXfqISYIsqRhV9oUY0Oj9PcG7UbTHTi3C7B766wu
aER9qOwUSLAAPuWzxHHKZcvI0q3+37/MmYAg7WfL1LUSA1bzr8VmS+ZbZ//a6Rj6
5b5jgdQmfv4ALwoBH+vo7V0snvuSgbJb1Novb66ddR+m5jUGwTXN+qNm/YJMXD2a
q7Qb7Wpmw2lArOAfsNslmCRTKCAg5o449Y0LxTDiQUtHQTGJwhmEVqbic9oYOOPw
B/40d7/PiQv4JFjchwx3hyDNxC1eZVh9S8TKW0KkdVhOTCMrDJLkShvlrmWLqvYV
8a+ZXs/5Lw3hHZ4E9Tst337jHZt/xxPifuYRO4+2TplRenWRVkCwn+3f3tAphBd3
5UaQ217/cw2pVmzCBY4vvuzVhBMRG4viLz/P8c5Bzbk4ojWNca2UH8SafF1E2fK3
lgfpJTCmZVFXV2E0Rwo1jOOk24HbwG5Od11HDHNEJIm+qJ6vX9J4vMpOOXEu5ZsZ
anK+15HZUN+0bfKcLTc4UBWnlmOG+JvglOBqMOmdfa9WR6M4OD++h1Ute4Xffjub
Jqf8t9Yu058ylPcvyf18zBS+AjDHlts13/ihvUlQFGZ0XHvEMsAvjQSS+lSSxS31
qIleVaY2u6Aj+QS/JYo4zojRhV+XZgx3Mfct+cnGvLi1j6K4+fEix5jn+jUAYYw0
sIfBow9zG9Q66jqvXDlqh8/BjR1+RTabWDHspNtzck6iWkkFR8POinpgMHmZ7Nc8
Dg1hPmVqhMkLoE7Yo7IMvgWSqz0rjP6uXppKWKnl7eHr7hfIo5/jwx0nhVDO/Sq/
vRdEyqnt0K4aRwCUaa194c1zDdS9PNwNI8Qlybi+D8jdikpI94eprP+y4+oOZFkc
0vaEB2Kly4kHdUWN0pgYTF+/QKvTxt/eDHRRyObjSBkHHqc8cX336rDS5EjtrKzQ
mZEtW+gtoWlOmOyR//x7KWdDsyhxwUIrxXsf8BT8AvMSDwMQwQaiGDfnnrMsrjCL
b7kuNvUBw6IkV3NyNyUYLB5i6kK15y1SZGXxoA3MIGBqZCSZvAC/37jT/eIwfQGE
Ih4lNMtCE9nWabr/6k3D2AFayRfnPBpKPxSBD3jRQKO6IyIsbbavE1ahUmu/Lzeo
Wo5b/eyYTYqDn5/Wa27aUd9+NdKUE4KaEAHqIoPFReX4zKswYYY5C40aP7tLyfbC
GhxkjkbEyiII6ARY4daJ/zrUcjLBll+f90pHxmwdb19yStK0SyYNt61+1FbpOFbB
VinkQ/BfF2mYwyWQ5ocm1UKph8OOM0MKNLQ8fPTVm+OFXAXAKxE8GqlW3HwMuvsF
4rZLyRaORYYTwMjetyZOXuzSYfZTXi/EHgj9xr6WTW/Fb2GCUD2FCarMOuZtWAYX
A/AeAHSlmch7GMyX50/5/kcruDvZ1TiWbakIZG6Q8t6tTIml9ifTGPTZm/hPzRFk
tcChKN+h3jlee4LkQ2zg4n30e/sfVZCYJ48pDymmxmnJsH1fgMMVL30Iw5PDms6s
2wTKrVG2hK4AnnNcNqS7y6DhFCUa2n+DuSbkesUtJhkxZONe36joa6M3K0dajosB
DgS2yeV1z6R0OkXlHzd5Tqmk+BkhBrMrxIU7x7lNsI5EjLbIkuwIFerFgI/dbb5n
nb2QHtMekkj0Lj0U3qk1UuU+Q5tox672DyhStalFp2F7Pc66o5dRnjJL0v1cWYRs
R1iFYtENFiC8O9oeGDaFScaugE1wp5ANbhiG8UdJdMWv8LSnQgolWamzQ6MEO9Uw
SZAuVQPYr8300kLBK8binP52ixNQ1AlXBG+sORrvJDnOk42DoAYDfWqUcUi3VJuv
f0ua5kvmdKvtjy0oOGE+zUqpk/t89Xi8khKamxGBd6b35VFdTKR+nVkK3nRFvG5Q
RevPt1EX3W9sHrC+KdoBOARb8C3XRJs5RjG/cpfWv3SyqUDQxl+z7Z+D/jVQmscH
nYmaAC08xNIq2/NBIW5mUw7pf/wqtE5yN6NxFBFygwX/q52y36XUiComkaWnNyrt
jYm8IXT9CIC4fHGED9P6RQuEtkC2x5WNMmXNpMNOAI1JGEfyH1z2hKXrWT6bEyYc
/V4Y7hmaDg/TBhLKzFTtsIt1cg0HMAx90wo+3NqmTHYFcuPZMAmAdK/i95zX417g
igwMKv2wlgTag6zTNpbNBc4oaSiE3VINRoKiqJOzA32tH7lmyu2SuyQ8P1NVqrSl
Ywa1TGqCxiy+Pt3xBvdVQBxi0jH8ownwqGZzxP4cs8VPGCy7Vn8KsJO/E6RfeLHs
rativ9pxhQSLhIuVcmHjekUqI5YbA2vxVW5kczrIWVdllBljwTgCi4+Bd0UrWrCC
4oH9MhbAMvcvfDCLjcxiKV9LFEX5blZR8XksPyB6GupnIeobHGFcrMMAA8Kgn+l9
kquXo5cmwKkA93HIky2K92iHpGyLJoeKx4J8j3jut1tljE9XE5Ku7k3WpZ/3oOkL
hBn5oO7UffiKIDtL3Kde72/SlkSWPh2rRshdeieyZqO3hNntgp3PThgEbCN2Nh9K
zTxQyv8qlO0LX0z8p+ibhZC3eKQiWa/yr14JeXTTfOBfOIHQLU7fsxiw9k3J+YR0
fHe1eXMijwb72ebL0rnCs0UmRrm7MYKgp1rXbpfiSN6YzSPPrq2lDYwndJY4uMA5
z2OUzS+yUrhKpT9r1WEWpDekMfzycWKhNCgQiuBYDpGz1GOTFf8P1rZJzvAGNpfo
/yYghhgTM85d0Gxph/C5gRVOmxxi7zFPMC8Oy3wn84a9sffVu53qlkVbo8//L7JM
oZPViBOBB5eE02UXDTYXk1EOPrQIogKeWt+ais5Kp+eYvULDfupivm9XWZTDECpA
SkAMwdlXvJ5H7N51ob0kOSCmYfBNCgelIxrCn0ViINjOEbBZQwuYPq0xIkxoVPlz
VWJolaaAGJVy2dvP0fk9VJYw+NdD2J0omDD76FgkKiHfILMTpnIILEWLYCV8jAez
OHvgP5+844X6trtK4VUKAbCU1azJH3pOFylnEpCGrJqrCXpO4fjgXPyQraS1DC4r
6WbUw46RygeCTc83Ee1ceKPp8qhTOaEXOD1mfYItw0pJozfCKrgr18jc57zWJ9GK
XqbSvWqfSbGCnmwCMnwwB+r3H125njXyX14Vq9+xb+zuxogPDMWBynJD9O78+7Vw
GIJorrVvobE6ig3xcoc4DbnF2y6UTfId8/QgU8mwytpbzJoKIqYYgBHPBbIhA24A
6qVEjnW7IvGnWsK/7fkAhlQybWrtyLzZdjbpf5X8Fa8M4FXJTq0P4A3HJfPeGyUz
Vk43NPjBTSxkazo9TW2LB2EJtu32xOUlD6swu7TlMbIK0GUUFmnasmEOe6pYwiwM
WOo5b6ftkKLL/dwyE/rxKDjmEhHD8z7iFG3euIEAgcti3GVofiROUu5tuP5XxIZX
gYFLplAf8kbvkEIp6LLsnT7PVWEKGTSc51vMDJsiAOw6c/iYxRSkbJHTC8hLZhJk
Ul8DtTKywQI7jMiADsqKjF/yGj2s43zy5mRRobafk/8NCf+ZWXsvuvbSXqhx0iO5
NvA82y7IGsB0UN1wYINxcSZKZS9WWh1qKRhLvtIoLWMPDiKcGUkgBH8aAABANRqp
WnPIZbEUeZoLnRhIMVJlie7Skcg1ynTdhBy4sdYYPm5wQRUsVaGc3lVtzxLBw6/Y
NuKNvMqvh+nsxU9SFEUXJS/QvLS2D39l9X7OuoOheD8VuQQV2OYAmEXB1w7mVBus
ogdQvN5lN+prEnEUzt4L7uobuPbcvy7XhOLppM2jKbkFDL8Mp5f1xJ43BGzR53wR
kmXyMSBGhElf0iuOw4Uo6F9gG8qY7S0qdTQxzRrowOgdQ96JN6mvhnLCNC+/L2eW
G0elJEJd/TRcCVMs0beMDkV9jcf5dkmbzHpufitCxEV6ryIAHEg/JtRVAUyva8yE
dwQOi4HcpOxCIeW1g+QCtgrbitMPLDuf+vrd2pzPB/YVyAIE0JIKGs8p10ilU9AS
SqF66uU2PM7YfJ/nj0uiieLt+KI3aXh66QOVpyDpPEWGzmp4QZoeN+jrvMm0uq/a
FrumP2xn3UNHQ3ZMrs73lOdBHJNPaoPYsZAU4eHH/plAUkkX0pzEyGD5T7qqx6cO
jN93qOCBpYaaeQDEgINGh4wmS5Cd5g57DpsJdGnZTKJcxNPopFK2B7mMeiupkGmp
QBFFoCoL0FsQTpXjoXwUOkqmhkT/eW9zy20oFIktBRf5luyK20cPtYoxLFVQBAlI
jQWSkITD7XdjNdmhMuPKXguEREe+xnuTSl36j4HzL7lcIn+RpbZ9Im5/Y51SlvOt
UdQz7up+rOHp4TxXqVwvuG/KtmN6wFcztXiM3i5BO/NP08lz4cocPPGG8ldfZTw6
LZFhYOI3gfwFHDcLX6ZvlY+RZJWO/7nlNcA+/MhzILw5GbOvrA78OsvCjnOZNr80
7lECrwW2081Hu08cPgKNoyXMqLCb71rEt7UqTFESmYT3VuUt3pzOmUkhaeEd8rGZ
QLpDDia2wU97r94uz/sT4+4odRJoGCaomFRl8C7v7Ffmai06cFbWrwUB7NFwckIt
W9G21gJYcSYiDLI7LaPgTmRwLHmX6/0QSQjLQ6LJDLrd1K4dhq40Chb4yYS281Fd
MHPyelzpHp/Qx+AP8VwBpEhk7OuftKtOv1OFpIJMTNWx/iIwhHqS9WDEZqeQ3ZYp
nH87HOPUJ+IvgtqvYOTQlU8oq9SkgYsZvD59mXw3A1tl7a8yt92WphoY9vQEYL2S
ottupIytaFX9WlmBc7sPCVq8eZY87u5nulWE/jIErxDzoMnybMRDsbufEtJqGi5I
Y22pzNDfReExKRFPksVoGr6NG3fcCTcBRAkIWx+jyZp6Vw693qcG19W7xEHz8cgM
SPUBDp5KIiHiSKTO6kg/u7aHa0pVe5ns8txHuGVVCDi7QIrH0f6ks1aLaGP96QdH
B2TZJGxTLuvsAA5sB/zNWHbhZYfCBbkSWvIQLjj/EPVfNCmf7K5R2NEKZWmOyYBi
p4DtKZRYwgy0umLXNj5USOxxlOmmzTkTXW/15F8L3hbwCfhJ4MbZN7x0w49K5kN3
Zeu1N3bAZ1CGwyKhdZ7EMCh9JDlit3pMoWGQQg4nSWHqyZLEMTnvxGWq5aWJLozY
jguEuEf8tROPdewBZg2sswQSdjVgS5doM1896dDHpVcLIpub72QkjmOXIRDFzOLC
oS6HicGcealTlIk2wiwb6sVjhhiCrqLEwbNCPdt8dD2vtBI9Tzz2S5Mts8ssprei
FRGTID1eaH7xEpdAe//KHUY6rBA1GvpUMIgsfomx1uImY2ykbMdQqzeDPRBI3H15
kB8igoFq61sb9CV0GibQ8yCf7oVftCD05pDHm2xwBkG6QjwhOe6MvwVjeQGd3hSC
euCONFYxTcX2VdwaeX2ur6BArbRLXOGDJlciL+z0SiZOxBQCaTzqFnpVpB9heM4r
gL3NMwXUjsRwvs34ivM17TqSxuKCCTjffh9ShWtbcTOT/yV/l6V/b8yOInfNMJ1G
6v7SaItY4AO3HqkjvbUhYaUH3q53pHbjDgG+VkZBrsJcyIHrIJF2s+ei+XSec9su
yEKli5G1Onj1a+jbOdKyKtVd891OCJLZQrL0dIxTxeYoCiN+fMNZt9j5QVKMBEvP
ETreLKJZNsA2fu+gTp2YHOw/52CZZ1rlN13KW9I5ZAhgvSNxqDTRdi9xx29xZx3J
WuJ1KEFcf+8iFzCMU/KzrAF5SNgjeq7C3r7YiZHh3D0Z3Qwjxg1E2mP4mQs/HUJR
P5H2zi9TNYnUPT71p+p936M2fHS31BHt9QMCl43wq8WUdKCgjhn7T/1lFiro2EXP
09E465T38/uICM/CDWsWajJQLiiCgRsO0H6BBxEfQbBDcUzf9kOsaQ+1D023ImGT
9ASVzv43Yzj1wsTXP44hvfT2zba/WMfNpSZjvxQwDdFB8DCBJIFFWE23ET7rlDA6
qJBpcUth74eX+mCvJ0xwNy4sWGN6LHqh7zHyWCfZ43hrk23Z6n5Hx0MZJ+U8R3A7
IG/3SuNowzxGsCGBMce/o9/JKWt/DfgKu0mD6Rltw0irAYO7v5xsdllYZd9IleCk
qjpf9tzV35CTNjLXUJiBPXFY8v4ylS0fQfsf00aom0x7JC/T5A++X3X+zCZCCPBC
FMKoo9rt2I/JycYscR5mns+EJPkA/6T/w12DdeUBUOEXzo28Qx2Y0QZ9hdP3ENI+
1JeE9D79WLWn2POEGURsY2eRs1HpLLwv6M4hTCS9Jqr4EBMMUwPBg6UAnOJdMYbW
LuKPWfR3JzioD+q0E7gljtVze2GdHvrJRvVjZWXddJfFqw/SG2iQgMjAQv2xZIQY
M7KwWNzM6rTdNAbBPOlWUxb2p4aQki+YKsKHyRudDHlqnDoKresNQClFRUdoKh7r
jEUYjADdmzkidqW0ourPvk3a1bUgZ6X0AGRGmQ+qNDwa+47maFpzhR4E1rmD3IUO
f0dPgW7JPNnM8xCwbhkk6LMbyKG6BS8w1RdY1sA/WralC/DVTCRjl5WCfXgZfnGf
xrREIYBc107/hCIobtChOOaxCzxreOMk2t1P/qyiN96UumgW+7RwXpig3s0CB/Yn
M3Za12EhKJjL/S/Gs5GhU5NwlyqrkJS2ODZ1JMEeJ3U4irOKymG3uIiqIPBkOYYr
p+pNPRcca1fKMsEMe8tw4T8mi823JK7QMQV1Wp3TTSjzHavTBgYGIoEFiw5gD3xb
+vz1Tod793edxXc08TYhCE+u2ZKQxW3nPW9/lKon5Jt2NP8/Blcul3uT8iXc+Lx8
70payirypzLbA5ENHX7ggeMf/4ma/3pInJwk8F8bfUF2UPADQTUOvX+RSuU+YMzg
GtG2t6Qo1ZfFlxHr9J3DXPNBaeLXhGpz6XF61I/v/uMejVkbtSCNTeDQsXAs8rJa
CAgQkVXb3ZWOuyn4KfoqmhZUdWKd7hcBKd/VqnM8GeWxZFspQ8tZ9zzI4LQE+l2c
LVtcsHw8rL/GIlIcwFHzuuh8OybHxfS/LEoalUU8jjz+DSJRL4k++3XQzcx88+35
aVuw0Q+9/sPQ36cV7aAI1HnNkz1FmQyVEnNt9m6Yb9jZpgQmuU4zUcw8tCBd2sK6
BJkzUiYEaKcjAGHz5yILpGsyguVGqLHjN/tcgqrv/kgKVcH2rzxijvhfTqgXP4Ch
AG59DwMe0g3DwttX73cUeW85SA+dTshz4Dhm0shJVQqa3uIPjAVaZFXCH/yaWdyF
8UC6Al48wrqtAK1/2GSWWtRLUpEfMVruKt02Fxix3OW1qoO09wtaaXg+XRTnXk6M
IUg6vg0SUMgps9U1Oba4RpwTJTYMiQcviJA2Lfbsxl3+sjxvdrrU2w/HUKxLE07u
BgokuLLXrdXSM/N/LzE+VMb+kkwiCG0+Qd2F4E4lZaQacOMkuKJhwPdIQbBau4D3
xrMaKDsCA8LGBGBoQq4hsKLY+lT4BKV9JkpeUysmyFbZXkkZ+fiDUVcuWbQd2Egz
V2BRk+PDeYouiDMfcg1QR+yP+t/xCCdahJvbGjcxGJ2yziip/HSMrMnVJtCjpGUT
ze5IfH7xAlwxUm8K9xpLTrgViUATrOAOYkUaP1fSu3TLcPXQcIyOgd6lG77tFmvO
itbJn58fWhO4vO5isbrgxRNKNIP1cetEqDhWwKl2UZpBrrEIdqvhJhzByPFkQmHs
k8xittbuJBICFeRmDFYjoAnvvFGUn2Mow1DehplAnmCroKQQrp1WtQNUKIDpNTcC
tq8hjVVsy5c7jV0eOLTzEjrgjDaMErDFPWZmMOrCZYahCzA4/zn4VZtMrkqLFnre
ohrbqWyoFxrUXApsiSyAI/E+Rvp6YTBO6PfspiOLLsy56Q3+WMpHok4DAgP4FHjH
Tiy1pdyYnn/68pj5C/hpISodlKMtxVJQ3mkV9IwoP7CXx/emtlZiFq+894JJ4IlK
wbEF53x2EXwM5F6r9jj5XC2SEnZJdM2+2lrgZfLipxqdLj3vHBmwjv+sZ/sB4ZA5
cnTBgqQ0XUVNW0qFxZrEeHw8AQJtbQeDXrhSmUZdeXtWXQCVv6lEEFaIP2Z0NvG/
tKJ0XmTucCWTiKEqvyD1StkCsE3qvCZFa+dfx8sTgu9Wj0SKweBIeq0bZzS3pt98
9w4jfZNWFnSFiymouvl3koBzxAs+w9YqX3h5GpC6HzGKAabczgtw6jjADMnl81CH
JzLwl8oJACjesjRG6Z7TVYlwqpSalxraQQpbz1V+WflaWvwFfz7qVMsbL3YyPlnv
I8NNDuGWI+gJ+tjXMZJVRFJCCAI+1Y7jJ8rttKuA6/Hjmg7z3/nnsZpzkM5k+f+k
Z/GqFzO8DQo3FGkq0vAQcdE9mEBDjR5Va/V6bro3rZ8/oD0BpHOfaUc35nQcEtry
/zQtVwPY+BrZAjMB3Q5zr1iOTdiK0fzHITrlt8OUX2X7DHyzTxWtTIzodepKvXe3
WVVGRsB28eeGSwqu/oo6tykZjydFqGI4mqOrW7oQzUHyDJv6ZzySjg3QrjhdYCVM
DDZ+1od9caVZxTFfg8+66g20123xAAv8lQLKSbDCTAaQFUvOyqQfMArkCIFICVF2
8kc4pnCqVS1T5VEYBFYI+pyo2I3ocaifsorDEeoOgo6ZLeJLdwSh4rk29eLzBnUn
XUP3TkXHLAEW2br/UIszWuU0c9dboZwpvAQCMO2vMt85WDAPEAzclYgRMlCIehab
9vOZIhwMc+/p3XacG4CgT2vkwmFMbkguEs8rQdL/yq3hxj4FIeD3/Qu9qBRs/RzC
2Xq0hYDsu7bbmZSd+UdQ3ALiNHJqAxpglH6/4ymGHPtrBZdFbl5rP99ZNqHap1CA
L1MleALMAdPAOqWDLGTHGBlOka8ilfrKwqI2XPLmm9t4UXO+XK9a6h6HyWm79Fq9
5HdpzSLSH4FNj16FL5K59paAEPNEIwmuIqYvCFGqecPAL+do2uB1gpyUVGgEMsX6
h64TlJJALVg6nrFKb/6GsUAhKQ8jJ8++3R6H8CMIJbdc4YMKgOrFDeMWyGO3t1M7
6lmmrfzbLWhHbWR827+kDuTgNKclQijSGPHFUoZd09OblIJOux3ch0N9ERBW5nlh
5YKc4wElh+frZAd2W+5rDoF3CBOQDsy8rzcKzHHymyUgObOv25I+cH/s08E6Cd7y
lIVYfG/8pd5bGdfCZA7ZXGetQKxIQTnYJfsFGj/LCHSur8t0+/Qzl10+DJ6wXd5l
aW8zGiBPFi4697OZF5WDmVhNy7GkBOZRK8M4j3TtrrYtOM0ogodw0MlI83/yKiuI
I4C4GaCeoCoaGOMkVCwkBUo+xXZh+F3xCJeTCbAJzR5LKjq4azHA5SAykerooE21
aS9TGAt+YgO4vZ92F32yqfrqMaoBlDke+zFCvGjCqVto/3nIH2RNm9eIoQsSgv4D
4p8eyBoLgb934W2hKR9O8uTgzMeu9k15jZCBnmJHpAcexPfm2nW3eYMbM+aIAUqG
SKNKWNnGzcUqDdex3jqMIdGTP02MAB+iWr2/DMtfgmsYN888uzG++Q0d3cblPhm5
61fq33JZgBGxLyI+9B+ZNk966XxiS9EYuLGWmfgNjvEONlPspPL2iBfgK3ylYpMv
ub87puj/Gj2sssNCO1mKD4J9vkRj38jHhK9LF8R8+yxjaUH/T8hdFXUDUy66u5vK
obkm6ZOLulWUV0lmzjB1xPT+yCUAOJ2mQe2esucnpvd28GoRZ6vLf0W8Es53uLNx
UWd2lj2uOZL5N8xCd3LsbjXnAR0CvwGMWa3HcrA4wE0nweQehrKm+MymuhbP83lu
Q7+RerYOSDs03lsWb/Nkfufw4M0HtU6TG5G1CvPKUulVOvgNNl8yo+7AB4qBbsZJ
+i0NpYVbRx+nmW4bw/Usl+RkKU6D+keyiqfHuGI38wIXcKRt+byFnkzgRmM9sOKp
G64w9mh4eakzuiN1Y831ZFljORz8VO4pYKnQAkAx6LOa8zwAkjEkX+ebAL/vuYOG
8l/ha4ZJ2ttfcBiGd2EtqribyqTv5+BjZxAX2rak2j4y/NE9KAiBe3E3Ab2ZXX0T
agwFio/S4U2djr2tP9mtmYhk+VLhsIrWNZE8ThSlyVVADOzGEUCIWmgkcdhR1DRd
BDeqicRcAqd9DZXlvPI8+4T00IwaPJI/8HzZsgIna82pb7EKxgsL0625kG65Ytgp
cOuMkqPVcH2oySARUZygTClFiIxCIGnVGLS6R7kRJT9PhiOHWnPmMKlnExyeLuX7
2n+ENbNzLF0dedCJTaUEJt7A7XAYOHfj8r7YuCSwE8u0DiV953jLFcQ2UAFA2R0n
DyqPfHE7tvz1N+G8ItA+NttfysYr6pAdf9Nasi0aIjG8DZhUlU0B2gK7Dw+j63Xe
jMEh5xbM3tQNWj4aJa3ZIteMGoVI4u8ImROjcpslj5ieuU5MzHcyUYuZJGDBdHW2
MlOaK/oCvAfO2bKApt8OyxKfaqddbqsYJvJU7ZJ9QaC5WNpGdqiwZR2OVAvn7sxZ
mGQqqHcLCiCs6lKisqtgRTFzBrrYLRSiCLP14xgvcNcijSVxfqub3ZDRMbNA7BRP
HFCAVjg75ULSLellplfOmhx1KXH1vGZ2xpqi4oKHsi0dyqRyuFaeaaWU6pvzjp5I
r9GU6ItQpPY3ZicSdPPsjJJRa4FEDsLWy3Lo357XfZ8yIS8WxBlMDvJHOsLNSlr5
yRi1gkpANF53W0UnrFVYegfv468C0xF1FHoIpnGviHpxFsXEiXHx19oI2lnz/a0n
YxHs07ke5MqC8lYNvzaS80LfT41tqVszUB/B7tBhzfTcpETWqO60Tq7IE06FWQno
fpP5b/n30XoW8rajk57WuKRoMpYzuHGlvlUkqpvJckL7JLfltC31frBybOUGB26o
4UqnkZ//enRAo4RGgVgKxILquEGsSDZ5ILaXR6S/ivx+GSKuFAfFS4pnI7VYx+vl
iIJb6q8inyXQZxmsIlfVYBv37/innrMUJCXc2PxEQcpgYxQOUwpQ+Mn9COoNIR0M
AVvMh8zlMadI+nNg9bD8kfkiD60xV43HBGRVhU9LcilOAMXNCBUDsoD54/1sXNW2
oJN+YvJHGAL/nUSByXY01Ny8PkRM8SFjUB6/hOzQ3i5+4NiupQC2F2O46fW1ZaTW
rhMjfoQs826ZhAzakM9/vpaXwqUhcUxGGNegQ3YlxFmce19I7yzH9wAPO/q6Y+gb
SK1cuhtINhRYgLEU4kctj1dU0v7vNBa+IpgbxdbEoUq2TUKPeAZB/OTTFhq/PvXN
D9zgdPBN/49a7/jAZ1TV4LYg+rbHGjbXeHkFxv1dvD9YgXGlPJIKsF5O1cll6ZQu
8CSuIdqbrOQ+rqmqKvrV+3+GKfmbAX9it/yr6MSe8b8cjrQw1RhvJk3u0t5CMKvc
evyVrGm2gVxWD0y2TeY8U4IedtQRIGh4E/8ABa4jhChi7+sUd3PZkab1vn1y6HYx
R74duu3uDi/BUv8oYXu70KtBhoHpRs6RpUqxj4Gon+tp2A1r1u9vMQGhwEOUtuEp
oRMQtFEb+a6ynpzmBQA/VijJvF2aFbfgazJrCfDD9nixr72cW1JCg5gDZUMi6OKq
/aR7edHLFPc3Khk2oEVjPElKfdrcvH4WJRpeaNZKhse299xY1r7dtAGfwynj1grD
Xm90wgN1/2z2iybGrXjOUpt4zgUt2vfMLkczumsf+rXEkNjpBlHb+MiEMznLTHXX
WmP1dx/nmqw0ORSAR5+EkoyuuWeKOETqJ5E5L0L0oSaaNuG5M0Mq96D12lXm0eUr
9ub53hR3iGtIxCPtNXQy8cvzLZdu8TZxZLMjhDBkr/I4BqUIK39H0JXGEOAzt8LB
jiY39rrIkbGr2JRo7WcxfXK6GfLNMw49el+S78976LagLi9wpwGu+dHocuUaKu5I
MBCUB7jlna3hpeq25uoFmhrTN6H+mwaepEe0mMryTZM/XUAnOVAtWUXoPsc3cuB2
rH68Vxsn1vD5yY8cuQKFiez9VRrq7++6Aaygej535r+EWoRPaVHM8BTMUBwo4jsV
J1nn5O0FWxgHb3t+DXPz8L579iYGxFwf3gsjNIDVXHTQQXyRqrkkZHgvUGgpizIB
zzcQesQttn7lzvhXemZS+14A5xH+BYrAr2o3lf56C4S+qpSy0tlZM6oaXHv8GTpc
2iCXLeBqdr+WmG+bdnLeZMZysqi/tdOIn/e49ufhrCRb0oB0PmscaIeG9kdo4qMu
o+iKaAzwzCnz+/yJeEWo7XkKtO2ZsMrlR84FEAOAK1QpGq+hv/mpVeQgjgFn+qCT
EpbVbeEUxM3ve+KP9GaR/Vj5FudyotQGoR/PcTEiMpS5dNjaY0DeYhIXsKIR8xVh
JcrJZPv3NQZ8glBhfE63nohEBDf6i+Z5KqeSZbv/6d82n4k640fDA7EBWsRH/Cqf
NwGxzrOlGxswRtKDrxsIhNJ7hBXGvldX8xmaWzt7uL2uqQQUiCejgFZO2omANtzK
JOYzgMkUuk8w3AJ/pO/+tg682VeuGttcS1WslT5eVMj1TS5/dXrl9AQSJ/y5Sbr/
mC41wtYU1+oRG7taZkrrfllRE2EKd4kpeyzmdP0lKecN2P6lGkxuSWiHNZOch7Jv
xW2l6sotCJbIRSVedOS5buFTaW3obD03FUqJbTGZPacr+LTyPPmvugXL6Ya1ftX4
gvUq/uRlWMobsgNnzaxe5zLcf+3S8n4XJPWiDd0Dbm/pFYyI3yCNjBrAeCZcJ9Da
FUfAjVPBEjG6rty9o2HuhwqAlDJx1No48K6MNdR0nNVq9JEH+Qa9ws1ui5yUNVs+
MVTRY5f+oOkeeQH4lZDb+4zgROMZZ8qZhDRQTNf7FYUEtYJ73/oFPit56UF/ND+l
WVBW00mj8vGoZD0DsaP/mAnQkPti4xWxfc2m7YkqJIhsJIK7eYIZis4BwjGn/38V
qfvZslckWc2sD3EiLG0KKI9cFxmjFHXb3BPBtcvTbp7xJJ3SMgyHTJ5TA3okY/fL
Vf8a9OPpcQsoBQj7lgPPVm69asx9y4T7U96AJAsJcVr1zIa9zUmJOAjB9woKMqhY
a5puQ5Paquf4dGEl1W0iN2oXqhCjJrbpuw3CwXtbuqlUWHEaHsZcvxNSgkGG82yi
yqeEy/oIh4lImZ8IiWnIALufHN/5PB+dZnw3FYOTJGvKICFlIcO1A5zJtyiKkKIg
v2d4+yn8vMoqwWNfNleCYMDgaPVi8p6Dth1blhPwm8mDZ0hcsHfFZTYT1p7LTONI
qM0B61L6CDS4gqUyWmi1hEWSN5knyMk5/sWfsRiUGkph1zNq+z54rkcCfMP+QwV5
DNKMCjTVZnVXbf4xOFoyysDWDeQalbM+4hGRurzGhEDJJwRasELwNTW9jFGYgw+n
6rw1zS70yJl2sb0fP18H31jPayQaCH6PL9ZTSQvzQkKqoTCXaCCqU1sbq+a0wIOe
qjqLuiIXeAUzhIMNuTLCnmMFh7+cFWh4H2LeDUwEs5lKoM/SW7R5bGWUgteSy4ae
GJ+chWgGUUJ9HBNVnareaPoi9kw3M+gH5Asl5miqLa5zGzQh6d0W06YzLMQRIThQ
N/D45iVjYVISSoqyX4W0AZROEjIRdyTJ8X6Gxc3z300EBtQl2Bfl6YhRoru8uRqK
kDKEYxQ2+QNZ4XzWvKIB5ktiJyBC1wQ/3eClZlyQWaF6s3tXkC/3uQyeoHXq2II3
/CqPYYebkboRokQmw5GPNbZHdjHprO9jf217aYzVnnUNNOUkucTiZBFgMyW/knB9
tgCi3h/Tt4xS2BdrymDbjf7rloFEAWosUxVCJvUeeW8JcGmWfXPblXnZDef8NGy8
pPKGs9+7+EHzo+PT20CukmMyCT5usWX868z2ukcmF5so9bk0szGwnqtYpbzX7LnJ
5FFq/3Q/A5cP5L0+5HrjhIkArcZZZ7z9faG9EmPJTkfZhCNy11c3oiIcQ6QQwvVH
qoaK65j9m0j13hYqtGQMiB/sYMy2zrU0H73DTyM5g0bPz7PsdBTR0XuP1RhQ29cT
UxZl7Chvo53SxhBCsOypoUhyBbVU/wwstzF+pXTNeKUiEPSoHN+pLINeUPjnqqyV
KRNeARzmmcVFBpP/vvWXG/Ce4k0RDEQdqWaaZwflp1wamf0Y+L8yhLU6cNRQk58G
E1yFZh/YPGs1W2V8fJ/dCDooSo8bf13iTXwD3d8Fzw+PG7HQ0m+/WyiHGSej62b/
U99gEEq9AkiNZEnesZ80iSjac30q5PolSFe6BpUvECJxz5lHRgz1ZfZCKXhhAld4
1XqrSJk70fr8dp6O8/mSSIpUtkEw4T1vVc9P/qmmF2QRjkD6dwBZguhy37bDymsA
c0mKnt7RoSTImrIKlE50pYTeqY2EUCphqUcocWckDeIPyM0WWdm6EC4woTMoY6ww
hR+AWGu1zWYkbXCnpgZgNsAigT5OKF1aZfRNT25OF2WI+xRoCPnv3QmoExWNZDC4
jBoTneOf9p9nY+nZA/F0NLcB92xIT9E728NHWI2BDBSG1i+GflnnYDqNB6rdLP6J
HWHL6GVnQEqIl4xzt0yk2UDs/VqIOvc9LtEAgFNjGLRHNhQv1Z3AN3c/G2JFVamm
hqd4xVd/3yUEPbc+Sy6T6HTYag8o8xqU7Pr118sdShytSUh3tnod5M4ipLr6kb4F
f8zZ81XxUyY5GJl4jUeccAmsk0A5Oqzf2LmonVcV7RlTDRdnbgdtnPmAF8GLX4Wo
NRBRNlDpb/bUh3/fsta0u2JCK/ZdSn7XSGpKwygzImY8Kz2iOfkaphja04fX1VUk
o6rgpcYpgOjCLbP9Taj6JWdswLym5ksbjZBo1fDq9Nl+zbu3mE3Xd3Gg50jRHuvC
f8Tqz6Dm2nmlCVSse2IGLCDy8KTEAs1OHUXk/RtI4il5r3I92SWjgWF8uSUkrHpu
9KOcz0JEvfiicafftqlvwF/ahFjRO9bPYHv7K0EUL/gPooxuePy+Y5TXYQtsAUwf
n88n/uZVJ88D/ZcLANe2DmFvdP/KljolkCfC3H2ITShqJpGE7BSt/nmg0Kk8WGO5
/pF7FGBfneAWCORCCG//kBNowibgnrtwiKaYL2oTYa9eGSD3QenAz80pl2ZIUpGF
xK841oWEN8zG4LI1gqmGFNtOKKzwmk8h0GVuA1QEjAlZccGcsOBzEi1uOTki6Mox
wFW6Ted8RUd9qbkLn/pgKU8mHneUn/rKa3JhX5+9fLc1ZDX2NIo7HPSiBt/SIxrL
Jxbe88Fv/ze9PNt21/DYM0xMhKBzwwTlRggOcH2LSFao5uBucSoX0W/as1s6rbi2
9y46mvt97N/hjF/UOX6aU8okzS7awNPlNvniB3GRkS7C3J0gRl6Q0bO3UYpFMdjR
1Oed085OdkHBPAHV3MiPPeK8CQU8yY46IiI2rB6xhM2F1AA4QTX1pFF073bV9Gw1
AKtJPf+bL6nzn+BIpQFhOEUIfTGxLgKtNMMUeMEbWiMTT2fvqf7kxhjAw3QjNz/9
1Q8TIYEulokOotv/LY5uXGKGQHSyxSLs8FwrQEpH7zMvCpvhlBQW99+5sSpPdFhb
Rzd5+0lDCOWoU8uVHMYf6MZz88KSHd0sm+lixYHI/HtKJ723m8b86tGa5SETTPMj
nwWTGKXCB3NfC/jB4XviWwDovvmiwvzjrs1lau2EJOGwi2drOgTM1JHmjTjOHxO7
rPbRAzG7Iq130E9QPSutKYQ0fZYcTpWu6ewAW6YECV+/kgVlf2c5BSh6JwPZPE5L
fNmkYRzmP0hI57Ytu8J1q+0w7kJDnfaADKTjSHx3s7Au2d8vczbGG1C6PFdTVne5
p8UtiRtnr3Q0HSNcHY2RaiclkoLUE6srLg91FFNa5CX2gyzVB6fZnepwLfDJrWZ7
Nao+Sp4HZ9sXfv/7VdYD8Mwn3wbOfnHuOjkfMxexPTiYjH15yj5gr4FpVpvYaGYy
m3Gx2dpuP/ZCd4fli7Z3JjouW+RQlTZ6guhHJEq9gP7+PYgW2KS2BwcjcO2Y+HrF
0X5X9a5Q7pbDyA+vc3qXt36IWxbYJYcNvIUNo1C8YLs/TqhvJSPArcD/jpviF9Rk
2N0hyqW4yp+aC1WUaENHJUrMxQJ3og6zpr3cuS29hbqhdha0eY3jt2CkQfXFVSjy
QoJ1wGp/F8hIksopbXJzsQx+utXyzzA5qSZP8052NXYS2cfCQv21GFmgmKYz0JTY
+XctHrw+fncxf4hz/NO0liANb3MRQu9AfLaOvz3DrCyTm+gnAu+1Zih1TWWmCBsq
/TVH9cXr1vhjXe//xjTl9FOdqn+SQW0kPStPbF74Cl/js7S0IUJwQjBBYV6IT201
+8AsEhRO+AxygOpwZrndI8a84h/luZ+tHVZD/K2KOLK0BrzJ5YZYIhk0J8tzuBHZ
DNQUs5l8YOu+rrszvtAdbPcSlvS7MbjawUBoFjvim2S0qMO7jt3Zi3QP7O/K09vO
lLFeut9Z+AeBdRCNUj+6IiQKPzSpTwZ66rb9MILDzhEKJYnutNDAsn60j4fC9DD5
T3VkaI0bGQk1dinGxAuCwjw9kt+3ET6AYKCNPwG3TPuhyc++yx/i0Z3T8POYNGAl
wW9WG2SEFkz5c1r9ceqTIgfvZNY12jBmCRCXFOZPHEAYXVYM4YR8QipicfkEUWMY
wdApmPKQ0K1fBYcPLEHGn/3NAKRpKqZQ+ZxJXivcqWfAY3mJLENe04fm/owe5c9O
0Y3PH9i15IX+blOUmUTPDqk9rKXaU2/I2X4/ZRZ7zmo6btmD6RwcWr/vAXD8911V
e7fWWep32g1U2OBAu6lMniPgjX4XK5gFKygtElUq2Tip3HCXyTHvc4i72aedrK3f
osRotXm7QvxMd3773FEC2IrHx/sNO4GSOI0CJXQ3G4LHKdTueOKipzz/S456CbcL
rAr3HbzgIIQ1K2tom0EiNL0gUKFtLnB6iMuNLfb4/hHMCFA/eJCRqmxxK1U+uU5N
6PooGhEcrvaIfzxXQHoRGw11EWWu7qsIHAZjJ9xbWIppRGqTu6iuGi83vBmzD1ib
EaJivC9KqQrOzc90BBYQrmqiKC+N3XRothI38+QryJsPHcuqv6QKi717Vsp81NDw
nlg4DjkYIhjoGsqDvQhfNrBdcsXt4USuDmIopkLJUK50cNC1+6ZfO7W+VNj/XOJw
RsnQvfBog90CMYdUYzcOoxkOHXCfGq5TwGVcOfOBioxYDAS22B0S9rnDTcOAceUS
oLwHutr20J4fTagK4GhSWTtfw8zJ9G7Kr3j7F6hCPe5V2LVQJbNRC9bI9a5l+dy3
+5KNUWl8Z0F9d3CaEUCpAb+ety2vTpUdAnTDPZg22CICBexvF4lbrPB7OHO5Opso
YnyJ5oFy+MfseNEkJ0mxkeRqtaYAFt5kr5Rmv7SuiLT6/KhfA9kYVjj725JLT4vX
vb9G8YP+0ZrW/sO/h4aTk3qqkQXgFmmcuDnIMiMROlKuhPhjwqHAC5wFmbq77uSl
V1KYZ/qwCTHlwQBK9W+rYj8zFn1y2UmkftDCYHzH0ikiGorhfS1YiJFSeklOLoPj
C8xZjy3yr5RRtxwiUOeBD5PLLdSoCEWx4wdHnvzuzhxDidS/F99NAWUhQz/zasOE
aRee5EfixRh9IL69lbfh9/DyUaOc7ARk3lAAzw9ffi+q6o6NvRqzNN2jn6kMUG0l
l1+0Z65AFuqqyEJSQXxSO6rui6DtPr5BJSti/MV0Omj2pnTINlxk+M3DcV/D2sbK
YaLbglEiGhtG5o8OeypsqXqE/yHkOu1nx3ozaSskfyeS3aPPcdfvmJoOd+v2ucRP
3zZAkMcRWxleznjxhuc4ppq5PhMiAu7P6nz7D2CO2uDiOtKMhoqI0wF6RJYEeRKo
0O1kEXZZM9+EU8ZoYnhmfVo2io4+VJGEPJ3zAWApf/4xym9qqu7Kdi0bHowFxa74
xTU0zbf34UmIaoRF3nQzBxgc7nKsIave+DIXSZyf61SM99i0B4OCs98/IzUoc/p8
3EY1I61XyNhahEW/82Ca1k64/YptVLSNqrYea/CIKQp9xBA63baZ/sNGTtfX7Fkl
boYFPiPa04X3SY8zmA+RmFo0geS1UvbGT7VWhfTDWlMpEMozcKDUGPgLYY6gr/yn
RnPRrgOnapu66IEvy7U2Zrc1uS2z8sQlrmp9260jVzaONztfUSa/KkrYT8B8PBDZ
pl4jkPCIICbJ77mnBsvWK6WKHyZZGMKb8k/K5FdeY/wgmTS3BahJi1Dx52+q9JPA
nJRQjw2Z8ywYMcvnn2TkFiMLe0Rp9sfp1j69pgDLr3MUXYUs4eCz/Eb7jhvKEvIe
DgD1v1FAQls4ukmRa4BEzcP/2IZ+hhNmwfXbrBZ5hdKPi6KdpeaBbRN7qDEPpZm4
pPzpDrpk7K6ARNt1jipG3IvtDURuS0Pqr2Hq1TwHRlC4imNGagZuA+seBGvs7rJ1
vRZ8wLe3+irADWzv3WchlM31dMn6CKq2iACvtilOUTcyacjkL0OulP2mYAZCPWug
RCuTeqwdudJQqTi2mn/TceYWRuhh0hzLmCvlu+SH/MFPiZ+W2yGcxEHrn6tVGXlo
fJQeS1DBZ8qaJbtBUDSfpG/L6C1F0PESXZffR/mCaa4T+tqAQ03+7uDTXXONHUv5
AoGFBIlZDv7eQ8aQ/YV3e/+4u+4rE+ML/1C66pHlz/YUFN23b57aX+I+pCLzu3vH
y5Od+01YH6cT/nPMHroJA8CF0tifZJ5C1uSS90W2AAxaA1oWIdgCNIWTAINNsR7L
DefLEIh65HZATPY6/nLGtHAXtfLPEq9TumjGV3C0V19SoZNA/1eQM+6rGccxMZQo
fN6EkvtT7cnFKUHErLwmZwVyuBVHQSF0QKz+Lqku3qBoL4MhSL/17o7ztKUzE0oH
BjBi/GarE7/B3refeR4MWoUvrrZxncz55lLrn4bCLdvsufEIxp3cHdbdI0oD0uva
g4ATyW9GFF4YYaj/4G2fV8eL+zLtPCzHhNEdyZWdAciud7anCj9/ZGfO8WDhi0J+
SuLVf0ITgB/plgLHHOJvEZMUJMAvGnCYuocbzhOJB0lt/M5ZvUToIEMZJp/CwB4G
g/Oox+QrGWt+w+WUHaaMf8DYYPt0fShfH3TtCrAkogDx6jp4vez62802EEHaidDo
nYtneNyLMWl3Y1Gr0386HaxaopNpnzU0ejAPKPVyChMQSA7/eYXJ2eBfxFporQyQ
zFJpE4OqVYI5nSp4j+xDjo0EhbkfHMHi0Mz3iKrrRwPyItB5rCGhoLG0DpCscc5Q
hFAppdvjmO9G/fMWd/n3gOQVVid6RThStLRZjIO56RLuH6Z+aj1pwGwlP3GW3Xnx
Oa/Mqj4J+LGnMPZY9iK456hfBLCpdt4CxVByqkPtVFJp5l+TOBdsKiSIoo3e+jbf
HsMP27RtJecsnYlEiOP5hquOtAuQIVtLipR9EXA9xft214ENn1fpEoL+2sYOcB1i
T6QjrIUukALx3Bkf8u64dG8WZOGmjUekckw0VaVqfZAdpr0aOtUcdSrh/ZKh+Fsi
DZWsN1ZjB/F7RxiO30BDoJgZDJ6N7ePwCBpTaxQbNbNQj8ODvNDMjWzuqsKt1ya2
Y6U27Km38wi+ZhWoHJrk0XU/1Mz3ugxiuEyD7QnVjMHgjCVx37tRJUcZ6HoBg632
KgG4HM77ddwqGT3i8d5/yooB5X0W1HCCM1nLlnle1XinVeX1j+ry1TGQMvo5CYr5
XYxu4CyDVCCVubYf9+EMLvYgubmN3/mZ/BDGzM5rNOaNzyhrJA0JFa4ecnjbqOwn
lr95lzFNwCjVjkS/L0kMZ5DvP8RL4cug+o2tGT9pzT+sy5BTbEjoMf3Gmeq02EAs
qitKNXU8HJnUrnqPMz0K1KXg6TwP3++2ysvtG594xLthrXdobcpb3mpfrOT/3iVb
M4+BjWdUAXH71wk5wrfqitdalA0hSEDWpZZF7BovtnZPx2ZQRRCE0nn6VvPfYD4n
iCMGU3lBAuX5z1Y10GI9vW3VO66a/QY5j9bxt4TajAq7r+PtbuAZU2nxQikMmTWh
M7MKBv0iTU+dKiV8FAhuEF1i7Q9wU35kX6c0AFZKBrNwCvVkklmBjyUlqIJh2Ycl
cRXYN7A5H3JKp3rXCb5y/dR/7RjVa6VioAN403ELgW0v79goXjpjALQr9MBYrA6w
qdfYF/JTq4g48QwzKYDFJqsmJAqBq3rAt3W4O64mOeXSoPqLW143sstpSSSKh0cM
4eop6R10DSJziSrg3vgABshpXy3fpUVChJRMS5yxBjESeNDBwwr63UOLYyXduchL
HBYlk2eIdVUB9YfFRgof4f7xrz+B9WBmEWKEbCAfVsMWLrQkKOBBn2O0gCtDNBJI
1d32w47oPTnLF68oOePOV3DoBiiMLAa6kz3h50dGuSsFg+bKWtTHriTwGWnu0lw5
e5DMrXqPH3n9CTb2uG9K4e6+o4eevmrCBSmMLKg/wgr9jv+Pb6+JmyxGGDjN8zdE
MDRMDJUw+1HRN0mso5yb8zfrvQX+L82FTOOw37LF7LFGvaP32KG5S02XxHyqVEjG
PGJyz5vxOznmxb+9Zao24n6IIWmeRKA7tUIBA9tJNGMkeAZWCa3zAYT0HXZHGdsj
Xve/dKjcUdBgkiEN3vMNZHVFdpCrPj5c3eAht/wAdhd8FaTZ0YMv4GPgQ6xIftiP
yuWGcX8qCFXCWZe6mXRzvfEF1F5dkrL4Krmi6LT4ZcGaKSlnaPw0o2EOvjx1plaR
w6hd0Y2C+QqGQXWBhfHcAiJ5OWBBjoOMqeNf4Ijey+MNL06VNkfo9p1qzXTgKyH/
ajxHGwmswBIF2/eS8y7c7tUiZUe3ooH4/nokUWuvrJmY2qtfG9X5YTdXU9ucfGr1
azzXo3lIFPMBqLDTNFvD8vpi8IbX8KWm6JJy8b8m3TYKZOXTfvQ//kIbHc/yY4f5
9FjHoIzZzvMYRVhIm95upl801x4UlPaWJP8dc+8kYwveakApMNq79h63tPiXosmw
Ch9PRi3xlNPyp+WpcWaqFkfk2LzXzikpXhAg/PE+mtELDBFil8nUnZzO/OqVQGi7
buUYHpaWG4TLlugub5h2LblCx7pqTI1VmhYc5dSZaP54xIlV3iCBDjCrjW/eNV/p
b8I8XmP9tv1X/JyS2aOcf5WxxpCvWYsN/ce6Uc8axtHgrg/WtuafyAjWrNgXKfZN
XGqHfq0sE+66Hqyu3Mq2x/aKNHHZKcip9bSnbV2NcCVTpik5Erynte6pW6FicaYY
rMYmfLEJJLIxvzkrPeyikSAivzmE19oOBFLC1/N3YAECF2WLMmKB2WK8Fu+L3wCT
3RNIJG2245BXXcRY8VGail/DayKIQmBHoTgORPnceJYkQB2I9mO+SmqcmqLsteoR
gE9t2V7LfyEZdj0uWIw4Sl5lOK5GACOVsijGRxckOCUmmO2Z4iTOdd3kuZoudCWW
xjjLf+VbLHsFGGy/O4S/aXAckRSI2QdHSsq699mMzEt2iMUI/ZK9xuEQxR+/oKnX
AZRbS6dqz8WYQoCL3fQXFAFB0dgGAwr1UihXEeBTzUyrtZh+fiY6kBKz5q/yyMGV
wfqxJ0+7FWz2FfRD2w5wyjWI8hOUN72USObWRNpTg2MMzBf7gsaBDk91xywzxAPo
sEM6P+6HDrFDZYtSRpzmErdR1O+nlb01kO8Zj0Dh8DyNtPw7zQhj9sQrrD93+fOq
tu+UV2FOyDhkLjsqk6q+F2oUXSQuzaVMNtraKCq8Q0oCRoHwEsKUIfd96nPQ+yOP
eOC37klc/V6QwozkbBt7n/QbpfzsG9BCLsdpzG1Zrr3nDpPSP/u/wtvdpotNY+Yi
o/K/XSOVbE9JwveSMIBVb+gYf+9BmhTmeZOeqvYqsa6h+7rlikRUiaucP1y3OO8J
WkWgU/LVc5mxnisZpj/KOjXdbNy+FYYO/sOwo4j9hddUmgYnCmwJ7QccsPb+/O0v
lM0AhbD+PUfJWzrSC9C43vVnDYXWAjAYBzGnGUku1wx7lVyRDjDmbMwyRROgpj/e
9bDhMGg7TmvW0bGtyL0HbckS0L9ExuGZeX4W53n7mkQ1+6TJaUM1y97E3p7Hk35g
s++bhS5cmRagCKopfOOvSBz25X4KNqBOKCUnkeE7/ndvECDAbKb3+5LhJ9h6TXeQ
r+KWKg8C5XgeF0ZsRp82hBKJsD+yIuDJ9fn1nSe4jDD/2KYyyMsO7EaTf/84opKy
JGYV9a/hjbHRtAOKkBgchhimLvhG2hpiZ7+ThkX/Vz7vtMblXQMSjfAjOoN2zECQ
qJOcUcskRWk5XTSfJEf2gmT1A2CampUoK2l+yNGT/mGekL14o3lQbMlWPmS7wwZL
l1W8W4rkqywCE2S/JV29cyJKs+asb/2LgcKxGT9uQCiyE4RRYE0CTTOWIWA5iDPi
B1jokBD0MfHcZvoHa0dbmXPzYuOw3AQ1HluWvOMWWWwv83a4DIe/oZqdmNoWBSUX
3yaAydgk/IA8P5eLO6v+DBKMIBwaIw0YuTS53TTNqKFvvv/CFe9hygTzSDy2rf4E
JeunzUBPEXzQfpwiKwM+u2R5pgL4qe74kG0ykoMP1tLplN+WV/kLjFHxsi4YX6kS
eCLRhzDbsJhK58Ygz9pbTJmLvhY/hPb8J8CcK07si2uHA1jTLz1Ou0VlKoBZWSqT
SxQla6MN8gB1DcBtcUb8VW0yseF6h6niGMmIhWat9QoBfsNf00qXLITD/FgaMmqE
u9jwu8qbmQHL61KmZq2eMR7cGuXaN34dnNkAf6OGxAJ7wbmErlZ5X2sQuS/pSr4C
FDm6hQJnpUy1tkNHcS+tkDOS5tGYvbniAZEydTuzDOQLULN6YhFL8kDaqVhTwnRe
0ERfbd42CbdTgW2LaF2YPE3WaHwiH4TGQ4c203SElDaMj3+MP2p0xdCNVKT3kRLA
Mu4kmJHASq4RTcjAKAMUtuUoLwM5yskAg3eOT33z2H1qVte7xFNQAk2UWvr0sAph
HYlmdB9UFs7lpgM4HRllZTw21/LGzPIWiq5HfUtMAYR62MdJ/1C9Cv8A6s6qyDdu
RqaADSqw7psmvU0v9EJL9/As85GslfnR9Ci1fPNb/iQhQjEMt/Hyp0yUWtVG1MoX
NM6LoZJR9P+s95HmsLmqDM4q1VlpOxhWosgmfsfg8AlCxiGUcOJzdbcIJ38U7/4z
VbryhYuyxwVeV6/NvlJ/axyPTGg/4T8uvdOMja6+nvWoAGPHWZMy6LjT7HyJYyVk
Z0ryE4p033oC+4deniRKAhRs8b/sRna3jZBkmFeF1S4TeP0ORI/PloIM5VeTr8CX
RHQwWHrOZe8fXkVbXdIAPJeDsUCdzq87nkANnSCGrWa94LaI6DCsN2xY+KegaM/x
91KhyBP+NCZvd6LU6Du21Tkj/NM+Tu1MpDk35XiORusD/w/EzDm2b8jx4b/OoNW8
RG3TbbQ+qVVjFFe9PtVlzGhbQroolPLKuLBqX9t50w5pSuceL2BsByKsIVKqSj+D
hvMaz4/2SLzKZqFO0iwilVi4L+VJT+5hKm33FczEz0Oli7Fr4isb+fZF/2K+Y6KX
0H5R5rGcoTuJ0wEEiQaGydHsxLXCoUd45uDytw8VzkPqtx/HkxN1+dDUF+LUpTGS
ENeZry5LZKWO3BYrvlyHf37o2B+n+XyzafTFy/4WKGZJX1TTF8XontayG7GzeVoS
dKonT8pco0DpLHLlz09HX53fjxNgAak6NBHjYFqsJOQ22188/VAII90yg27iAeXn
muBCogEdEkw8l5gfoL8Qi7/fhZK6MZUkxbJzCSkidzpzb1Tk78F5MzXrNUQSLMwI
oaV8XLYMrYrQnYxRe/3gqMvfc6dsZ38elYh97jrrlX52BzM4ECvRM6cYolYyt7K9
bTrwrFJQX14CH38ZDPq05w2lGwGx78ONX782gIqr/Y+T9mhUjBkFMKsko47PtLrL
anfFZMIZbuARhcQwCKpECWBeMHsS0wK2eLGuqjBG8NOv89BpvwAJDzUMx7Q+QKXX
sk7+QWk/ESduNPXklByDkoayfReodZHCtJWydKxZUli9F7Nm/GLMb60NWuV3fbwT
Ahw6SrMGa7DfxjxN1Nnz1bRciQO67qCsgoOR1aiHTFjJwMwkRmt+T8twpyTpZL6Y
bfrFeY5ZPHWi+rId9UlbKO8xCnB2NblSR22d2+u7Tc44wrxJRXDUMqg++3lVBBJw
vXVdZMuCjwEBRvbbDdyuWTgyx5cdtNmqJGFnw7Wx7OvML9U4TTRe/YdYBzSuo6SO
3U8BWrRmYdhJkaXNMgjntDXU7TlbKNx1Y7Aa1aj6y+kPVE24TlaSEBL4yz3Vymf9
jtufT7az+MrFkApyWYLK1sz3sc7Had5gzxU3Qpaic+rNkXThraVGCDKA2GXwTquI
jOCYz01cNqDYweP+/Pcfnb7He+ijkdsxmG8/a0XS36uvmK7IwWCh2oFpPPMMeGEJ
YlGbFYOHawpE1VLEN8Cb88SvXjmw7jV00+j6lmktTTqXBb6ZhtHP6Idnp3lWzwOM
zYtmxQvIewS+DAqusPndMJWrJL0LSjPDOhJ0h0kNyF1Lyfd2mEhQ78qntvHYtMqO
RDLKvLRvTWc2ZAkV8TC//cWBs5HJMjtFHKQnNN6p+qotwLXtXku6T7eIralPHjqN
OQ68M10mX9Lu6qKCMBdEV1A72L9lhXqFBNe2ZFxYkDt+Op/75fqjh+FdZWqK+FbQ
S+UygaJNmisaOlBScdb5fwp5puS6OACIiqbayNL6Ny7sIjqnT+19/kZZcLnVkxIP
r03OZQHyoaGgM+Mf2l8lkGMnloeeb/jldvfqUb8Qehfy9i5gbxq/dGZvpT79nb60
RjRnMKtSWxqQ8SAX/OEQqtNVUp4lxmbChPs2wdiGAAuSvHd7+PvIW4RTKwFumyBy
tTblgSuSu9EVGkVHdUFPpmx6ZZR2MhlnhYVz1MKrOH2Xxdf3W7iRcVuNZWdo3uSd
2J2JvO6SifLcYarzxjHJ6rGuF0zc48IcUkkedO77B4UHGZeOGzno1oUajekHriAc
7MUnod4YO0YeVsXX491xMxTDArXtTNGqMyBKUBp6HdHrOeziTlV5O4odwFgCpeiy
PVlyx69nuPo3l2sns/qnPeTwC8MljOoKxDFioSQm6C86tHChhYlvBnXp2dHYD24L
nZAIwNqnGuO09ervDDLuxqPqAPpYdB0Z6H17o8eQBQlH1fsYH20mN7Y5LJWsVgYZ
ssSq3hMYYOMt+WdkmOXaUMqFNTQ+ljNPpb2Kj9CRCGptq3n3yE/gekNZyRZqsdtB
HpOKmwx7t9bb2aimfTL/Si/2g1nUbERAAf2SwfnuwU9gUedkyDHX72vrVsQW+0bY
S1T6XFEP5Sh7LLV5IBjmnfSUWhhqwdTQ1dzCBht9kZm2uVpe2KP6IivSEI2ybWOH
B5qrLUlPyBCQrRz7ppnnhoxPwi+7385h6aEYF0NmaCE0Suloq0ZQIdCvgmIpXpCT
YfRb/Rli+8/2axglKIVMqRe+fOx0AoIL19MPQ7HTVmwXR6Rw2N1pBmiw7NfbjCr+
NGhF69PClj4Bos4PX9oiY1HejIwv005P9WCm42q6ISbGpPg4R5erJ8FeioT0Yytf
8ttKQ2sSnj1uFJUwJWKoieoOIfIoAQWxDKoLLDme5bSHQbaULJ8UdIhDVyRhVlPY
iKJnMNp3VQvNuaK9vKWzeQlZHKUs2gEjqNjilehJarP6uMWCzSN17iM/HSo+dECL
8CI6bJK7fJQ8sgO3eR7to0sjzEa88xdmbWFBP6Ms8UWe+Q8PkLvMGTSd+njhieW6
1qQZYMCOB0ptIVQOJri+M72g2Cz05ynIsekatX+1YTubFYX4jTH95V0U4k+YsBcy
ZwDf7dPs1egYTtr9ocSaA+5OR60dcRJ26WW/BkK+2/NwLlDWQL+IvlXPCsJb6THv
L22ovhMDuiiEEVRSl3aOYRXBz4jAR8346SLhxNrdd/bFQm5T+OLnfj0Z4F7awSsv
K24tOE/qH8CD8/eA/J/OfsV9N20Ho7ENp0XgXdp8aZ84QVVYwP+BQ7lz76jP4buy
nQE2GfC9w+O6kzT2aXRIh3mbao/zGZsYA6yDfeUZv0wOLA5OVpzDn9+MIW5NmxuK
SFlsyeJMjCgbzHZgNG3O/n/Zf2jikRg6H0f1jvXiiTvk48Bu0oS+x9TKirVnttsQ
EyLjV2X6GY7KSv3Hpbx/ulJ5xpxSVEv0gGHpUV1Emr6UW6gXorfl0xI4xkMobieJ
75fVk8oo4w/6qv/vvwO87OGokS8QTJM5e0hWpFnPdcD2DSMjfuK/rUqq1aICa/Tf
4dt2UE/jM5yzSUIv702PR+yyCphXEbqbMZTskuWbR1kBqYykxHCigY2W1toT5/s9
QafxXnQ4BepAWyFep2d94JwAE8zedMiCrVR8KYUYAH8PiO5fMrfvy+GfdOEf3luI
zbHapsRrrtraIfqvkT5L+wRhSiOHHl5WQcdujoxDfQv2YzsNB5D4n0tqCjb2m62J
iZjQwJ6o0v/M8XvcidkxAEpkK9xHGSu2NcVVUjN/5l9G3/lTJFol0NhEKkhJDpfk
iaO10EaC3fwN2VFuZnubajDrRBJ5Tup86SqbWSFZtKXQ6dlZ8JqPRi0JVZW8gldk
7W3xRtT3SiVsGOD0AGhcKosI/m3fOi3DEy4iSFaJqXpSg+r3RSh1nRe5MTIRur+I
91fBYL8Usd8085RgPr1Z36Vq0BFmeqHD6qWM94uJGhK+Hr2Um7cB6rNE5ogkKX6b
+fGrgud0S1Tu51xng5Ge+vX3HnR9esEcJHF7ciVi8dfFmBbODT/DSs9bSeMDEo9+
MxdWPUmEb1K4tkoOPtD3W8BhlF6RGsadeJO1ujQr0zkNB4nN3cZScz7Y56p8jf4S
x4a8mg+UPyrEAMZMVXNOHZWAVWRy8BnzvMPhdxGiaP55KN4RU/2Ez86ygltlh087
ozUF7q8HHTPw8HjaInaQzjHsa1Fdn1vihY7+HJVKJLJSqhYsMERwompKgtsCwx4f
kPQ0oQufb1jQmxhUV2Hkw/nKS7mJATG+LyuNT4WbB1V5XL5zg1ZR3tpB5VIPINkE
Kcbjf6gqrYSoBBDNlg74YwI/bQt5BjeK+dBey7THmuIq3yJLpOgFTRjPtWAnwr7F
rGNy3thfm8vjPkZfQ5X0ocuLAUez9HBe/1Km+lzkAIYfM4mrYeZfxExyLv4rkz2e
qVbjfrkwIQhVzfuP4XW2aJn/Ya11hUxUVXl/jDmQYsy0qhU2w6n+/xBvO3CJCgkA
Jro+d8JmhGGFfSzVrTYf6ficY3KHWNnN5yP6YugJRT5JmMc1+uGpvbgZUOHGkw66
jUXUAIzATO2L7hE+nY2MoDaUzEtgdrS75XRWLZz4Z1ck2PkZoShVqKSsJZ7Lp8Xx
kz7dMgwiOKL6+vlCFx2MRgOM0UglBdTIFlm8Rv8dF0qbEx832Dj4MNg34Y84SAYP
si1T3NIRC+gq0RyL+SK/uRWsELt4CWeWpr0Wi6x+BAdV2uhi1W68X/yUy/CpO/rU
HkPS3MAixQ6rg02ddI17G7ZpbVVd4kcBSSLVVZJWzVol2bjAvJc4+5cWgsfiES9i
fhAnQvfxQ63veodHmXZIneQF1zkDNovdJnkyVdYHqzizJKmGg9LHjgaf5G7O2oS6
LNaHVcNE4EEIu8QVcJBWaih/dpEzTfNnCc+/0CLIardZZTFmiQGvzis/4oIHvCSU
XepskUa9BgTTjBmgztQ1aKT14+pbgrfK+ys1XZ0h3AfSuZBOkaSPVDLcEGjDx7fW
MF4GCMg0DqLgrTuXq+9ET/BJsmyhrVgBkn2zLKqaepZuow6KtoBnWwV+RT/MPRc8
lJnVb1lpS65D4oRWOFiHreoCx2BrezXwZ+tMuzL2WphMpbDcruG6pemoQgYCIoR+
GSQfmCscDTbU8zDcOkXQ7s9bO5C0d/ErITencMrXOukO5Dx+G91tLXATNJ5Yzt0m
I0hsfRUJV8UnBoLQEL9h9bn64N0Y4CPIUXa2tyvOnO+Rm7wbWR4nf5ciVwP5LW46
C7pMk1cKQ1BVoY43BEZHZc+c/iOGegYm+OgRlspqg4FPO5QBWMA7sxVoPUNMR0Y7
v6YhARiEl9b4gm93yRUZ9HXgdMFN+ShuBf4tHOkxMEr4Qm9vWWdJYDZiDThtN02I
KmYVoXPeSuEiWzuUmi/KNo7E4IQ7MWRb1dTvfT0yIerXIdoGt/avj/YyhH1kgClU
PokFQ6sYF7OwkXQRV8055aeGUJoxLujM/CbbEvs0b8lz2oW+iom7KwLweK+jNcif
AQaifhxPqivPr0s9edTN7Fh/saBxRJaWrmKZ8Z/uz/hwv+H5THaZDni4XjqRzEsm
OPH8j7z/9uz8E2dJCSvwiRAqKsXkrtOasrDOvVhvUoOmVBJdUitcBTqsD8wrXIae
F1mkJSQTwHtoLTjVAoKbinG769hzb2e/Ynd7IvY0DgbJCH7H7Xop4oVSCdywdzjB
GUwC3Pcj7ydp30VUtpYoE43QLzffxffKVXaImE6Fb94UxdJz1aekpFqZGyr3Dfrx
qesjXcnWJrRuJ31j1h6Zy9UvZRdEOCZ/0MYbLqDZ4cOmOS5XAIqqSP0ORrYuwgdZ
a9bJSiXyosIA1EAOUUjUpeRZDDy5jjdeKvHvihnT8IJ2cxxiojQRtI5tby+efIo0
Q/mSy53oPXvyOT/hm65ZKyRenMPcnjBk41jDHnipQQYQkp7X2qR2h5ZucbZzH7Gi
0zzp9PrHpBNWqNlmdkxd3jCTv8uixspYd2T/tVCS7rRt2VtlShr2Ae0XavvKTRAL
6PosHclTfnjNgCYRm/7RVk0sXkoLbTfQIY9RBUrd67eL2jorE94MPqSgB9sAClLf
Enb7l8xXjwZzX6Pzx7dsKFlZBlvA4tyvKeSYnZXarlPTXBM9dIbmcL1Vw3eSbWgw
XI7dCumTddR1fnqcbOLdeQe7SX9lVAlbXKAzp792/XTsnzUSmck/N7tCL0gfwXj4
0cTS7cSeQgDhdtL1KonMWSGF32/8nsb3ByIWKcyFET3TULyqVUXngDkhGpCiL2PC
2xcTGz+7rceC9YZLPxfTMunJQBVlmS2IZvcHnvq8N5xAzwDKE9tNJvFyyrmGCzUS
lS1ExG/RiFZ4N7S3egvFZuWF0P5Twh2BcdFdTOLEyRn9O2/m36f5nY7PmWxU8x5J
QDMIZVIV+4K87UG2eU8nN9rhx6yp8C3ZoBYEWO0PTBl/Y0pnXkYl5jpRpkx3uyb2
ucvNQ0epn4zfucHlI+Zwk42b/NY0vAoLWrB/raUXsAo74qwcNeQzV7Wfh1bBn7gq
vlCEvwU/kB7xIMN24zV1fxMRuFBcZDT8BI+fLa14HQl6vUhZ0iGTmbh+kGRvSxXZ
tV6Y1BSc3SXPRpof0xzqKZMUvQ/14R6lZZRgGRwk0HOaeCMZtxeBxCgv83rP6qts
v9bWoK+5I3JgFR7E+Q87uGpLvUCsuqIMpWvwgbrgUllwLhaxmwMBCs9KE6sp7BD5
97fS9e2XOIdJ40xnItQrEzUDGmVh6luz/je3VsnaRGtl1Lh7LDObSDFWOhcXw24x
jtO9Ie5vq79F7cN1bR4SLitNJRtl8thaw6bQy3NFFjMG60607Eg4K5evCbecNB2+
LUxEYCkSNBZkc1edUIww+eveH2KWglnl0qo5BdtGg3Qy5Yd+oftkte28s+L7E//s
bSljIdAYDn+mJrfGbEfIRc1r8LnJblByCfpaueUAeDezv96xiibNXWej3A0XyIoT
RRfilUlPcPsR/zKG9uVakaB600b5r3ab95yKUlE2uWx94DI2S200O+52H0jdhlGO
j/hU4RcZM72u+QMdafRXHyf7KZaHeKCif7nsum86TXnbNyxRgyFRFgLRS4pNCXcF
CJJ2mDnUicxQ1TGhzlfO2ZnAy1CeeUxbwQllmEurecIlWfHu6OalMGJGXP2xXPsh
iBWTvMDAraA7RmItpwXi649xpmwk45cMHN06DFUYjNlMZzkE5ZGvhWmAVI2IsnaE
oN0h1Osnsn44ohEyDLjO+kelO+Ji+61WKecHy767NtnDnojpvysL7IOuF5qdZiKA
nRylxp5RF3cClUDHMMiXonNOVFKOtAqCMCJC/GRvLN0P/2qqpFv/ca+mNLHvFv9o
TRm3SGQKO4P6CI2eyCxhPo+737EjyhcLPzT5Jkf5kypQohBqPp3uk+j5HHUNtWG9
8RMJXAhvXOJcyNOrI5uM/RNll/b1DVaVJgUp+iATGchxnbuMJbNGXgEOh2Tul2YL
CQAtfEqFFtnEpjvb5JQL4ciNB+QhwMA0sdR/8C/Zx3N+J5W9EAjT7PdSG5/xm+iC
kjeZsSWNS/XSXTIFFZJWcqkluvtvfB8NIyRsxugIg+sE8XM8vidhsHfoS4GkHxoC
QSqJ+nxblDLmBPjpnMA78s0CwEtejo8Bpe8WMDvRxumx/X8xRFmYmzC0o2dY5+2F
YpAQeSpjnMSEpoN+OIfuWV3RlALy4WrYOnHcCzBtbV4F1k7qnp7787zWCbODiM47
D30IpGaoEvJVIJqIkOWrSE8o1X9uKRvqbiA+bwzlGbIAq02+6V2d9eqFPNRgwEXc
kUss5q2IDjuqnZCGpCgglG4QhcDKis8Fx4dqlvEImdV8fv7kzGyHVa13MLARBD46
IGQA+eW8tedmG/UIARGNsZpvuDX9+r8uAxrJs4O409eeSw11dm+HWUaoNGbbBy+v
rS7s6pVVde9h/w3K1z4kB04BhBJWV+kbYLEm1u1GIPiQkkKFvjSrfKgh74+jbZG4
qIE0Dli/cvO5z75hTFfLIhgbKRyueNx18rqmUFVShsniOUMcX/mpml5RoBnJ/ADI
rNgpSwCVDCQVgJm62q172rsd09BvQ2/9s1WITFYqGGnOoxjBErFrm5RQalNwyO+w
mNWg3Ko3JqSZwSHu/bLiAEPMb7xDajFCs65Kv361tO+HGVp3j/kJS41EfAzRuyQu
kSy6laMb99S0/Sn1dnLaNSQHPIjksK6j7etvwNUdvKcBTVNqyTOx5meAsXlUQ60I
HI1CXI8ElbvPPpNN/7yNK2oFLX9iVKb1rQlp3VcYn5VsyktlFMGPNhbTAbDjQtH/
00vlE04bNqJLb6zHaMj497K4U73ES5mC9UnETUVM6MHjP0pLAe+YbjJIi41kiVem
Q/FlxHZIPNtcSaVS1ZKfN0/VGj8ihslaQyPTwFmnKMufRD6DDJ116PrV0+vx1atO
pVl49ELQ9T/uQEJyVvCr9C7Qzt4cgk1dy5Uz3ZNscTAOhIno9q/NaivlKwKlQjR5
FYJiNeCdaxyaSGpSAXtwv5RfWtxYDyDtISLJxHe+fDnSsk/YqEpGjcJYKdxG7IyV
9aclJgc9LwSiZ5fFSZG2WaOTX6/TJ7mPjXQEbI2T0RjRdSkGgbymijNouRGMZv23
yAbMWnesmFDxITQqJWcVmoplpv9pm998elKNR/DiMyotR0rbmgqVcql8+gEgUVcU
O1H/g6ukyL9GymkMoG8aPiTWoar/Vm1glMwE5Q57dVGmZGza/szJ3XZyq5AgxMmr
9V3MUM9vlUDdlEEsFy2CNGTg2vJL7cLXiC85EUh1LwHfPlmsL9i8TdwtPKN+oXgm
lfFD1wbPEr79TjFJEQbmtEN872BE7jbkjk0YSuf4GofvY/Iw+8owpePHIYsL85R8
EP3R78ZV0kTzoctNyjyxTrHO5eydhhIPpwSy4JNPRNVWsCy8rwnrDjEwvgzq3+hc
zRZaK5ejrUm2aZDSCpR+NtQcPROzZXWVxofweYgsjBNx2SMiEhvkQDkLYENHWEFa
2XiMGO5P+rDj5et01tRL2plEAJzGw+t1oo855JoIKD43Tq6NqIAbfqAzZmUehiti
zhWiODdiFk0YF2g6QxbtUtfYVTi0uEM/xsc+5y1TYFTUIJaqSzbsXeN0Z+1VbVrj
ATrQYef2wby22yo5wJbGWADwwhFI5wg4WFBCN7zJ5NN3IJ6K77Br9FQjV/2EEX6E
GmKerWLpMNHvKz+3hhdwv3dfFTifUqvFcLXH2DBTKLkcChYSz5+Yau8E4fRiLiJ6
NT9jzP4GXkyKfpoX/By6mJEcZgCfn9VbJwU0Tuh/0rcU8mhXTmmZQj46xzWYSpeN
t2uOJk2/WleMVfa4yaN+QRtSdBkcNDjYaKE0aR9FVuU9KFbZNskgPKwpUxONCwti
ZEtopHxVyz9jacfeOY/WCcelkXGZ9RCN270Xp32OLwP7SUa0RZ03YMcUujUVu0kE
7rrH+e6e9n2Zk0PUdkdYjElQgxxviKPEKtOLcm2kUXhvt5uakYlNN5uFgl/09pJc
XJl3fJIF/26Q82+6Aowwb+DjAUZ2aulosF5Gb5O4Ukgy64Szn19a3IA/D035jUYo
MkgDAbcYhI6vAgtBDU04gZVsYRzhYBW0odA8dXsp5ec4YC4weH4YnT4+udOEySfy
itmUK8MstYktNERTOq8jCP5h0aB06/JdKM9FaRlx0F5D59eum03tHDsVq/dQm6eI
2XKpTyr+t/Cpdf1Kfp729+X+/x5Yoyx23ks1Ul76N8lqQYEEAOpdVBerHGT4WyjF
ud0/i5u14GmecxRLP9IKxMgPCBCz2rlA6zeuSf273P4RJm0eTJvEgyzI1uJdB/mg
YizXZiUEi2Re0Fpiz2bKEmIkPuimlI7VT/zyZ+kQd1Xz81vnR3X3TsW4Z6VjXus6
3Y6jdkjIDJtbGDMDJ8ENX265/GoXLoLdeJxAQn9Y6etj/csK87Px/OVKdkQcEZu/
u08RF1lRSsmOiXDRWpvCuHFcb4DEThNTXmw5dMaYQEOa1zjr0kFyMIzXoHJRgj4T
2EI0zI2TCZhGIwCrnYTOzeNnUbxiOlFa3BEXJ0ZT2jpaQ2BMMlipfYD3Q9F6PUZa
aP/w5HNiIbKrREgIjyIH9/G75FoC+tSdzMPjKnF4+qOaQRnMSv8ePxYtrrW321fL
Tn3FkNd9RT+7Tvsagu7NAhv6Chijmxcb+WJyZ5jRa8SBEBLFt8/YI3fR3S3+9OjZ
sc0cet5MmsBZ3XMcPH4PLGY1FYDP9PjffpPaImauBUem978xeg7fx9rNlPfZl5Ye
Zo0qtlhVNVQJyRa+pqHMh6MRay8/jy0/FoikuqPGHz5JU2xA5oAVOhMdkEQoBgiK
SCzgn2q7KZL6mcOHI5rFRsBred3E91lS/OarphiN3QZXwgRrswhLttrnPsdxzry0
or5jTotShyVV7i2wpE9PSnig5lG7QDAduVHs6AqfwU61pVgwU8mZ1qmgiiVHgCtP
AVkLVQFx0G+3yn18Yki4jJ/jsF4sI9Fkslb1OygV5x0Xz04/D207pcSdh8Sd9P/1
ZR4H82Rw3oTUNE9eSMaIHpv0FArEyDlzyx/c5eICZTuSHPmE6/yaDw/CtYd4SaOw
8iDe5D4etCxQuHfV+Oz7RV4J5J4CAl3OTgp/BReGxThAp/RJ2ikAOE7lHv6aRxJt
oCjGDuYnwhHrZlVu8B2856F+r64fzgw55seWrwVqSyaoGY5SXu1mC17daDqe/MoK
rH+Ds1SoSVQAy0USQue//GGY5GwhfHlIe7PIypot6a+Nt5pzE5SmzwHkqxc+V/Gl
oFscogA5MeIVxq9R+DKGnh6y1zOLaAjUBtGTU3Wd8MkSphWFl0BK8LJ54oHaAmBZ
gH5x4gKvli3JW32C63RyEk40O9BaK64WKZih3RopvaNXrcotldYw2jy5jrP4b41J
t8PE5qOkmtaWSbIAWG1VAT5gjl/cZRTlopOtUWkEoFfSkMFxxYpOj9EFmJVNp84d
4EzbelvL5/pbWCfr4dGif3nWY/nRVvLdaQx0UBl+d9tz44PxXYpsSI7t2/bmIVfi
N1T/iZiUdX5a00jDeulVcBMh3P1CYYp1A2vABzM+pU30Kq2xuFb2Rj9FxoldoTP0
l0rBY6mHFb1tFZu54vN2mZlbXDorGyeu6VydxGy3Z1/O41l+2sut1UgabPW7lwja
96UUpIXuTF6kyiPlXpi8O5dhWzgEPNnQ2At/CGMyFqMxyICuQuPAKRCbloc9S3r/
dFmCqpz3P/rODzgHP8NtstIpqJM8i55PjvjAaZpDaI8FYeaIpcUsE7G0HC3SISP2
hWw5t3Ci9I32dqgyWcGFrfzS5sqBYlqf2DPhbHOLjFGRjBsuwl6Gd83GWYYDwXC4
czDPVyosT0gzYT2jlrA/8+NIzFZ8M+dQmtQNZEk43q0juAQ1vtDmfbldMiv//0bw
cSDT9ujKF/XJNksU3kAC3WMNBDUR8jwboj9dZjRLRWdRFKkzVL7pYcovbA3OWG+u
aMsnopBKvz517QoyBdqcNBqWmwU9sTjaK/c76TABfNHLFmH6SvA8ZZgWxYUpssbl
9rmsYin2FY2Gszt1nrA3CDdocMP0q4KvQSy4txU1xfFxdjyFMXxdrzEObjvNRxmJ
gHzXLULIlV9P8pCvAMlMHFaXzHEO4M5kzqrok+1xZDcVF6pczNkBWzUu89u2bvWf
OhCagA4JujSXlcI6iAtdd7CFT2AOfhQBdqHw28FkSVsmblKe101/pClD89J65v5P
RMmRKQsEc/sKmppthirQ19bVImW7UAq0oqaUVci8hhllnBzISugNo2GyyN18Anbk
lEmstNsdBUfoMX/j06jb42WR/eLgK/uiWRxECzWse9Kl/aSd02eSFW4snrqk5uuX
MEdlcO8H8Fy2cNlPoLgZYbPDyzNhrpXjuzH1MjrUJCIqKvmpG43ioiTdFSPtjoxk
AZQ8IhtMrVNY5wA5YTNOXX05zS99A4kpvxP8BDF8vd1DZKyricbyuqjGqA5n3s9s
5cT1hU0N+mszDXzf1paJ/0BSvXmO6sedK9UzFFggewu1y6qI/dN6JHDAs/fyu1oU
9JKTcj9T1nWFKD9QLLXBcDyGI/pjE/nzgj+Yza2cuAZ1QEG/v9tUQ+GVOL5EdUwV
D7NuBWPq2yiEBd8khp77sDWLKCrDMabMSP19KCvbDO0kqrsRPhB8yTRwezIVeFVb
teBMxkykVmq3mmi8yD4wiUo4qhFwLtPUnBVdxO8bUgNLGPXJwUMOiAa9uFfu5cE4
vJb2W9R6GIVJminJc5xMioHUs+NfcM/5UTPQGpfNA+YPyF8BdUKoP1EAyho0iSWP
w0N3GYZaCAKXbrishew9gGvyLkMUYnfbwwKVhd8Rq1NCSck89PN7g0LS7ED36jz7
ZKcs9RRJC9+N6NUW4a4jVvvkPeDRfVa+PQCSQLc1DpkL/byiKVIgHcoeJKKiLxfq
vqNiiArH6ynMSEkEu17T1w5IO42PNccCLe5TnVJXQ4rRbz5kpHx1iS9B05AiFEgs
NJ30ViiHP4GiNGMRL7jwINaMLHpUQ3hPFsylEJxS1zPwLqZduAo0B8SQ6cnM98/8
/4jLHFXpX9+abevSOpHfQ7RTmt/uC1i6Ug3Y0j0aMFUj4HLZqAWoZm7KWxvJltYP
bQmQJkvqeurH3lQzZvGJQ9mSHZsu+ZRNz4UF4UePibsLrD719aD5vJqRfAn04IXD
Gc4/aft/xUd81V+vKMBcoJDCKU+nXZy+pg/CtDjorMb4X/cKrRK/0GgJE8jnw5oU
UrVkI68xAvqwLJn2p7dbnvls3mXnB5suB0rqpcZYKId7Dgl7/OMvLrNFkFixxZuW
iRHBDeUaDSaoQHROaD5GqY9toOgRMHKWpU2PhGfPTQHn3W2XY0oaG4LlmjrzRNHL
kjojbxL2cfceOZe3Muap8d6dkJjJ9XExcb+rrzOXdIadNJmDVWr9hf8YB/x3FMcH
1s7al0+z4wfeekog3pLqDW4pRjavQJ9QiqQr7qk5UYyF9hnZIf+UVhi5ooZgDFo+
Tnkjzp9U1T9t2vPwLwQBsFJ5wmj/nbOm+Ol2CJG/IBmXRCuf2nOl3hhCqeVEvu4u
x+grpVBoaxjZDMnycw5VWEL289iZrMAQm8lOivuEm+8LHfd1xG98FJ2i70uA4ikU
bcEJ1489pMobWQeQrbG8QND+8P3Qfq4O90hTCNFukQ81aKvobiBgHKbvG1HjU1O5
KUJB7CfhiaVmarrDSNjQUUgzfiFQ2B2ZgLnut7DRBgoeLDOfL+Icg37JTF3pOMVU
25EcUDkg/v879iOL3fQUd/LzMgkgO4u3b8TJiLhZ7k3cnB71ZDzINvBxhXcgWhnz
Y/ahRzyjWQsH5uA3AaMlNUysfIOZr2++rgZDzj8ftje0Ubgvq/zfUodqWXZBKltv
wPiFSS1cuP5IgV3wkbNEASxrq/cA+X26vSLmnp5T+9OI487nIrh1iT4hGUFbkO8h
0+wVrnWUinT0X1VycwbBTebtFAvlNNWY1SlNBUlQCOHqZkrqQCpVX45yWR5k0zVK
sc2AmPJ0081g9IsTZvo7OF5Cm/Ji/6Z2LrMIeW7wCt6aSvqbCXLnu4k09S4mWd7I
nzTQ5D/BO2oBNZs7a9lTroch/D2vMS6IRKDFuhZ+hU7qtTSu6mQpucZ8BKBNkpdl
xtYoqVVtOvpcmq51KaTkZlai7zdBY017tqm2sjTtdD8yUgGbAd8JVALqoHZ3GBmx
ga8PJhbu1KCHlD0y8VUSA9PFTs8nPfhvRIzegRfvtAu5b9Pf2MLPnoQmYRMY3Dp2
LLCkYtInsC8En3sPT5DqNSqe905dJMwOvF5Aq8l8y3QiBnE7Yb7e6PL3NOcyap2z
hGYF2EgR/qbv3vG+CqUcZmb6NWlC5ugcYs/4miQSI3elq7lkpaJXsffnmuPI0y62
1xYKQ4M0HozUasuppc3V//O23qVyZJF0paQRqxYN7P4ZFKoEyzZcFUe+66FM3fAF
7kUINsI+t5DUeaLOYK5FKIA+DimNXH8QMrjMwqyLkPlpsw05HE/FCIUT/TqXCupz
rnwVmuUg3Yquqs0g8eL06K14wkF99EyAoRLm+Bwcolh2I7L09dPWnq7hek9Ea5qv
dxjtEK0qnmkFxXSCvp5eletimIaIJGBlkNpcxav3+603vbTP8lxE4+f2DFYMhHJC
QgpfmDJLyv0AH90/Un4F0Du7c0KEVIhbbc2T25xqwvXeHzp4M2eemyRuH4U8AWTe
dTRlsTrA4VGSQ22xiorecVCrir86WnjjdZ/jY14OVL0QdwfniyNYAiy1hEvY4JWg
6ch1VNybWPRD+956TABkhAVGx26X3EifehTqnWkAiNLmHD+nV16abLgZOzlIyH/u
yIFzR9NxwvjsNXysQnZoXQOWy+DkzS/2SbP1lFnEZe1vmcZ2wpUamSrQSX9P9p1n
le9gpDCpnoyOE4sZHDjdKhG5QxrIw2bsmVWEzFL2do7Ms2fzM5hd4ZSXQ8nkDtcm
Obrni5JA1iDCrpQELDg6isH6+uYaUueLpuIpDJtq1U879uMEe9FPVJsLvMILarHH
byYVhUm854YiwuJ00uVm5qGjWuD+BisN0CrT3T01Aicu3B7fUrhddGj0e3vKwrv3
vK/pFOsQbrLLb4A5V95OaNteciachFYlgbxMXcdYmsDiiJysvUmca/nEzEwm746/
HGiSae4hwDdoOs62vk0xfoWF3oMLQRDL8axzsqlLJmWpqFraQhQSPYv2umJ6+bm4
vf9KjezuKVYiu3sNC/2d5JO5eeMlrQB2yP/CA56fnSv650NeT+Zqq30T103dydpa
VKa8mKsAB8RHG3wT7Jvgf3mFG/YYY7ctgHN8xS/RcX5/9w/hRZofPq0k5VKpRBro
3hLcA/uWiqmUf6bI1ZdAgZif7W5/am9tPuBN/flQ5IR/O1kbtmM+YzZCnCuNMv/R
/KznbUJfNO7Alxchd1ECFOnE7xlGSpW8ZWg0aJEPyQLdvch7K+4Y9+hfJWRxrgDI
YHnC650wC3GVTnWjz7u4DpSx06uGfIWBbqQQoD26+BJBrH2Kk/SjwJqqIdJ+YriT
fpKFBQmzp+MjCn2J9vCTtcmY1TChMdtz1s/ut9Pw0wLaqZriYq4ElgHev8GrYhyn
crgrw2DGsW1leEXrLdlEcm+DG3n2c47a6ZCagP4aSuu1MObkwsNqHILP9gpxkVLZ
dS8uBAk/axi8Fr3IW4VVmo7RyQjMZo6Buj0pdNxo8JHEzzBbLzeW3yknV9kltHkz
wzMG7jaDx9PzPcoSNz2VXzGGgskC2mTysVzsiJUig+4/6x2htFv/qZBBEeM6jJ0z
/NNx6LZEktUgSvKXxHe8+UdrdbET3qPrkB/AZRGrz9qcOxYoWB+kKGkV6uN+UU1K
ckHKRO2e6wPcYhR2WagyAydpzdJeehZ6kFUQlRWAwE+QKgyc/jdTmMYubigPK2gX
ky373N4tNE7Ay3gER0MerfgQPdiIeqTwpRkyJbih0xpX1LUvujpuUCTXBoXXTTmD
xREZjTke0pi/4YSbjYH31UisokeewelsuOMPu2s3zyhrGvTCD+VWXrOA66+9mwWJ
YdX1iCNYxNd2vm9Pu4fBqDBOV75NuO93vo2nPI0Rh4x3dCzIO2W7d07SDO6FS8Wz
sqBU6Vho0m36l+d5IeNYeT9svZ25ZPkFba8JNsgrFCo9fLmVNpjbT+AjkXeV2fbW
Iged3ZTHmZyS34oEUaQ7aIE21h2QIqHYyWY5VgZDi1o846IGc/sOn/fa4dnbQagF
ffWPxr9l86R2q7sooBalAHOsSoeWyso776IR0v4NWSh2ty9gRSAR9/Zp+/WnZMy3
Ko5oTY7gDxDBj84oPI1D7FRw+Oaeogojy1udzz9TgivOFtOSkaYi2nD6jsa2i9K+
0MjgG4c2txk7oUxWIVdCDpfG0oE8nXi51QTrRj9++7vJ1skiT7LzyCe/kqYC2iIE
+u5tViIE5vjp5VsNSpyEg+NfZ3RBo04UO3OqF5x7U/9FuJrl5FLBDF3se08MC+4i
VMMhDHaJ+O2GaF5uQziiF1ukeD2xGXqCv8eSGVtY4VUSltK9tZyuO2253vTQLpgB
9BY8fAkWGlMxfDXQVwO1ylVlKxpw2BJ1rmGfoWsALw/BkRknj+R1Ww+wu2UNmgZb
e/pJut7wQyhWv33rnttieGR8kh2HfAK3lT9iR6rtjhoX/Rv1D8MYw6iU9K9pYGoz
/gJw0VwY7xqjYVTmRlwwiYMwBg0wxbow+xNcMvQ5bf5EX95j8O9rUm5xH61IDuhG
JNrhLIDparfS1qg+w/utwpUzZQQGbinHx6cNQTY/QSXOOQUlyVq/HLA7X9CyJDOD
KDXawvDTFNDfytR/rsSi78Yyn19cUZKuCV87oghSV8zOW33RBoqX2NedXsuCyq+z
SVl5eBNso2t7A/2CscbPispSCwMbeLIoc+ceiBZZQtB7o0NQJkf0GDVelabhsrjZ
1qxBxawGV/Pm2H86O7+eeUJm9VbxZqmtkIxyKHQ1esG6OdACy1qTVk91H1BTXCO6
IvfXRIIxtZtN0G0/cDY3Jj7diMe0V5vcf5/+hgE/ppwhdCWxtSuQWIQtsq0iNgnK
RKXdrD1gEQ03VSmmUG+TylOQUNk31sr+vSXykNpiiWIOtSp/fkcXS6VQn8Sj1HQ+
W+u5HJfL7+u98/JHjnCKwEdHaSROc4vOOlyDRvRTLIYAgFea34ZMBMlR3lmjWZXm
CUT0NKKcNwk4KJz4P0eeSx+q47dXHKsNO9OKmvgqvzs6l+c2K5JjP4JYx6odX3ZP
J4EQEVWhxkGMIPZm7w40ULmrYBdnsYYat+tAn+wzbLklVE3aTxBzb7cBE0fgQULr
AFlHG4aBDbRORdD4ZQug4Z3Wj7YFyAUQt5X0yar1NkNfwB7WdUvbMbJMKF+TN0KS
qMSmSkdQY7hZmuzZSX77LNWRIPsxrxUHbHhxHvRd0gSWlI1O0BgU8pYWhwGvRxT5
xt0GQi8lulLyOQzLToQ6rjZ8vMjPgJSWYy65idd2BqO1/6v1Al5CKXuhMsSuEcUS
bV/+NHFm8s8mNtrYE8i+cIbGYqUZjn5IV1Qibdpn3+NgvrCjEE5vL5jTNIFQ2W5m
zDdVVBPd+kw1oEaKc7rb2BWkZo3QzfGh9Akx6FXkhz5QYlvqV3oKzVcMrRDpHmFd
bgXeSXW89vaAdZG/eN1F/Y/PyPnLTlQ3o/CRagRWkBo9mgyKn5y63QDs54BaqcyP
RuVzhMUxd3cNCEdwVJ3Buxw7Yxd6PQWq8WjxfRo43fccMVzwGVtBmY0S5u0T6g3L
RvSUDy4WtXIgkakD8/fyh4fR/g1ibB3o0uviTV0K4h3BsKyeTHZaZRoLPvBRDDS5
qedsxCtfp+ghMJII5WnWE1SvhhhBaDu7/qNGPvsFYf85sKS5Va+krwX0PaTcS+Nq
fe1TPHjsl0flMDrXrfMxtzw4brkjNLS0T7QA2o8TZAhUkjncATOdq+Xh5wy+5GiJ
W2D7f+gOzp/6lIGD66ly6JfE+ocyL3GJfpGouQ5EF6Y1Ue/k1O0L/8p1nzkNr/P+
owabLqjHHWBU9kMNOBG+KB1JiJvgLhDe1Y0pOHRHsqu+X83S+Z4Lu5riQ9brU0oa
X+ZDzIO3QqbPGVRiDOSqxixujHkfejqToQEVe27UsJl/0XGK5YTsjWXoNssr0+/E
J/5hIzUO3ZLmLq8iLcCtGkhzYvm+w4BhhOLkizPP/lD4vG7RDbR36gZlrr1kNP8s
yvq/Hy8JkFZkTrd0O4CoCaFJwe6uFazRq7yYEIhdRtltTRul+2JFDWpO63f89tAH
kV707R8kYHFqPgfMWzxfG/aGKhI7oTYSX6Bq3pq3zmipB4ctloAATAux6j9AP5IQ
1TevFuqFDeGcEhcjOaHRgGlCFr57bSJhpXbylI3nZGAkjvTw4JzutvV0Q8NNoX4n
jJ+CVqeqDLrCOtVxH4htr3NOjhqLgC0VuekBbNXUf2EmY0cEM1EXZYnZcw0a/Dpi
wSlwtw3aJSA7hWAu4aV2AMJ1wpYbnnYM4fwGlhbZnm2l4OGRS1Zza8FhfYJZGBVp
7is2rFnYGkQFQNrJV1W4Db2Nxob83zmIRAZ4T0j7QRoXHtgMIp+VpXHfACRoP5rY
7NNz+WgoXpXj5tRh/NOHt+FjaTvMPc185ABoSv9pnsEGL/XkUTBJvGIs9hI679b2
W/wtb3EXNLyCM5o/4OLafTm52u+rNCBs374zzbhsS3ZT+NHOrhTemUWyan2bfnqT
cOVwOFikXnw6/M7eoIy3PiKTF0Enl0kZvvvV5glvMNnx5vVDxs+X0s+cHQgw+kxv
yUd09zb4SPDZiySHKmbm8yUmJRkuN+nqSSvBEtl0vTKEnUkHTYGWVdvht1+BoY0y
1BKbOPsMF55fxSal11l0cVtLS+Fu+lEzTC25vM+5arTTsizO+QpDLEBJRL+vtbwn
QGsfTBS6uBifNH6XsBOY/WX2PJAcbOxQylU7f0VsHfc99so3Iwk+ovdBk0+JPngS
UUblMoQ7JavN7/FW2WkpqALyKouye35ffmGqAEtplgQC5TeMsAwYWbW5WVEhen8N
09MeV0j3o95GnScoKMxEKsqqkcnE3WsgitC2F+pNJrOIPlqWOjCg4uqaRpsInjON
83ITU4gStuminvGwa4t73EBBEDi61+oMXDm3ED0E8d7MR5/L+hlDwe1EcG8HJOYA
WE0mEgqGFMdGmHxPSv4+RFuKgXP63U2/Y4qmbJWX8Uqu1BGsj/3n5RoUzKlI/YKU
ZaQwiXp7WWdGc5+/u+9ZNd4tjCFRhS1bRRhgYaGYphvp+iM9dSdjCvpmz9j6ueZt
v8Tsz6O2CNz2GlZ2oJqMUmGZes1b9F3YGqDhlFhIUxVmzIZLXkKDuOFevjQVBi6f
PbcIXUCUhOXPCyDrV+ShadlgTx5p2HvHjIls92OYPllIvnsTOueHvXNY5xLI4760
WKJM7PiDSHf/ttp4CdRFffO/S/00uarMx1mZGBMwEiWR5R+O4V0tx/8mwQnlvs+u
nv54p1pQtotUQMrM0DFD/2gutHLJqjBzvz3bp8WYNqkObHiM5/DT2a2Adhklqdpb
KmQY4outd61gqSQ7Ps/20ra3eZLfn6Ix81Nq11dwirz0L3RIyF+CLvxHxwxe1CPm
9+oCR1YnNMPiI1EchyiCm3J3vlWYWv8VKddUHzyypF8cB68zTdKjcDnrO2qzYeb/
+y5LqI8V+8nOzHQOhP+5+WMaLd2Q4V2GIguJ49FYSzM3em7AvhJAdMIHA370O3Of
2W0bluBodpKzCox5N8kQg7hRAig3oD7RpB08Gr8ZIumxsiGUcvRKqfxr7ByLN8lb
3OBFuERPxW2dJ/X4Uzu0yfhmnLwbsjrtaqVE7fPG97qgZs5t+TllmfBCzgkpxwYR
9ea6Lp/py0ajlR4TiFtPZ8dedVmxqftQGbW2na9LEdN+BrT87CcTqhjr5yTi7tSm
l0NPvPe2VvhhkR/AQDKsKc7uhwhy6BHtHwUoODj4p37CTShpd5qhTNfhN70AJgTT
tVvMG+YQaaRB1mWDo2aCOtFZTcjiiuEv5g6pBPBLiUor9irqz5qMFXbDRQi6tEsY
JX8KWKxNDgqMVGzSQb7/Y87HLt8ON1BP+KGQO5X5482zEYR1/Pe/LzK9NxkttuhP
8MoBmGRCVmJvtEubs96L46aiPNZKPIqqW64Vr+lamcYsh2n0N6VYr8TmcHu+S/RV
rHiOWrexCuzWI9vEicnhok1djhdwGLeuJGL5qvOEShPYJuPje311pubZ5qkLXTC7
WoCM8cabsbkAXw5RX51Z0M4Y/VyWZozPI7PxJ06c51nl3f59nG6OgCvTnFQaGogP
5VVW4LhcAxisODsSIJu65jnlzFJpdRw+QKQj+CwjLNaw4RVbmbWTYQD2zj71TPV2
PbI6PHjXGI5jqtZSllmSi1xv5aoP3cZjzbIiDopBnBaxBvAly+L1Cjtvs3I3g6Nx
Q8i3hvtTvDGY1jLdnvHsHsI9dV4EzxQ/WodmhdBx5IGVj1xkpRcWgepNcXe95540
Plv9ypK731Q5nl95RxtpxRGEEUMHzHBn0v2KhigRQQAD286F03/TVIK5FnRdLrL0
5SP/LuV5i7FtLEYITjAqjGSlCMlOozRGZkIgsHhz7K0WMvJYJgRbnTqJcLfi9R1W
j/vnOudBG9Tw2VmBzTJQrrrL0WWRFadLhxi40EKwapH3nWDMV75JPFZAcUoa9Z0H
jx7WNcAZXwXppJKert3hmhUawsXpINBIePB/x1LP1JL3f9OVVtX0yOibNoAVMMi+
2sJ2NW0FBLzKMLm/rhONF3B77GjjmV2f4ZTyVOpZcJoPngXzrp7bwl46IVSsSWkA
lDaXq8sjk/kCK27TmtWWE3SiA7CUKsp2BhNkCp7Q8qAMOwz+ReD7P//MjRRyw2E7
AbR4JKBPSmvGE98Q3u2itPBg/19aVzO9LbDRAamVe/NAfgOTN/db7/7/elUgY2S1
D2plRCM/FpActs+ibit1+q7QT8hoSRccdEbilXjYXu1QIfYkTTb+lqDYRP3RuI3I
25IQroo/8NIo5eDgJYNoYteViEprw13UHYdJuZnWOCxkSKusibzkPoPIuRUmHGnr
hoN8Pec9BStF68NZM57J3PQXDfcgB0T1SD117rX9D8UkIoHFx3AzaDF4md+aHSBE
h0m/MWPAbEh75BM4DJGT/SnP+f4UZZK0X/i7AveDKaoXnL2UKaIymNI0nJkO640a
dK+AcfzzqNUo7s32NPq26Kv8rZbU/uv348Qwa2GHsW8YKW0hiuTbHzBm6iTbztda
2/DM3lI60e7wEhF0Q5imMnWqpdxcNsw0v8e9LUaJ3tanT6B0EgsfdoBc97USF8mA
MCpOeKTe/TIcjBkYU75McrNv1YezIOlmdhAQOxmERc2UoPBm6ewMod7WPEPNcLUt
DCjKZjCUwjMeJjw1MUgcLBcPYXV9tzOVViBAyMny0QT+0byXzqcf7pVZe0OdKTpc
rttq/Ggx6jo7QAONm7ausursC+O0D5YclNF2aTty6km3UCnk9uf0LIhLHY8QIvTU
4AO7Cj8K7NrBaFl/n2arkxb/Dv+OknEOmZr0Au2kCx0rcM0xpfcgPG8YBaxZjGmD
zMOcEWnuYjQD1sPiR6lNIOGZWe+uTqFcdo9Bgc+di3UmUQkp4k+kNl2wgdnhvRLx
+vz32ceFWYd1/5cRYVn6DkrRUoyMc3sT3Fck+ZfHznO2U6o9mFyGWnUHlEwvCzTm
bzJ7bAEOtYoDjt/T+OT5GKMPeEIjMuuL+1xidOOi24P7QC7aKRGlioMkBXMDw6n/
ZcjmtUZfuMJbqYQK8PJ2VtA0LBf5kPtxqNtWk3Kul063t35pSLMdc/zFYaAA3R/4
Dn9h4nAz8X1mNrV9bvQ1wlNRkmngGPUHbuZLXfAypusTB4jl+ypMjI20p01a+Okq
wdo3qCVWeon1oYCyabb1TR2/DUWrrng7g8/6e/nnEYxQ7QxK3oQ/vihzl8F05KV0
GlFSupep36qoWm/mc9i46uthgLjE2GmqKJbwPXMj8WE2jPNCgbIVYUYKmHa/PIRn
C4TleNB6RTaDJg/fiml7Dh+RvDxH7pUnmjZEd1kPQQsMTDq41L1fZ7l3DGF0ccIv
BO0afLqDS6DP/sxpkFLpThDHStr34YJLFXhf2JBMOV3VA099r+4ivZwPlt4P0P28
vlzRv+0irvVXMVM0qt/BtI9pUBGSdyJQJLbcIyLSWQ087F9OPNRfGLaMWdtiCLez
ZymR8XSVm5JiBWAGNfbi9Hexm6mlu+NSDV+U41E0P05N18TwcmGh+0PezIl/6Lxv
trn1g2xwKiNax0t9hPTTdXr6YnfLZrqu0qPChvIkldVbyUFgU4APuVrq7O984taS
V2lb2H6m43GeQwfo2AceNB0EwkvY/EcAalWccWyFTVJL9SHTG13LfkjhfS9oWbUc
0ndOCAqQlooEhl3vke6EBNkFU2aR2gTDLODsGM3+tiPJs5DhjJuD7mNqJeeM4eTC
XbXivW6coS/m+Qs5GmYGPUwm4pQC/NVj1Egdv8Dh/RY8YkyCoTmuhBY7Jx1Lwgsl
+Ft+FM+1O1fwH4OapsO74ZT7R3Z0+L0otcOpcjCeRClMLQHfle/1Qf2jIWzxy2po
+Ao0IZXnIrScjha7bRt26MGgONn6+liML3lfn4NOyge0rQUfFgs8+opIuU4/I8Wt
RQaQz8a89Yw+1RhDHppWMM3mCLUKVGnT0ll1hYK2VnSNprMZbWTWMlfAvEkxe30O
3nzm8hHUXpd7kBwkHua/QFm5QId7us2XVOcsRM7zVhftuiOo8EnLlNnfhobaWW3Y
wvVX8PN5nW5jq6j1w3J05kXX7SPjruph+mj/HJNSlWTiiuQ25WIGrjehOEYWk8K8
JOv8nvkOPyiiNoxn30+is2+6OKrFtNSzoLY957z3FnVbS9UZo7ww3GwG0EkxNX9L
mFCHdrwRvYg8CTLPBaSm3cTCImEj+sLZ27+Q8Pp1Js3QKhuLsUuF66Qha+VexiB4
bFF5Dd9I61Kb+fx69abJV96sDbY3OjJ8DluX9PppzsErJ9EXDFx5ZMRMzkncL5Sx
k1Dy4XrRk+p3hUNdNwhC2XppK5BOmzdeFZBnzy4HcGnZ4z8RT9odKvo6kSScKHoH
qAfQ2iOlxYmgnf101QmDz7Gpm799okOflfoqtlsnqR+QMJeJ6upYwe7ueGFxE2kT
qjXlzLSuh3eCz01g5SjI1QjYnJbFdYGprjCE7XroYLTBGECR2yzDlmRG3tccn4uX
MJ5J9iewdhmJXFsEQJ98f0EKtvjvaR4/FcGoKLGUt21vq/c0MTJPxnCjfMXfwr25
9kSCrQUIB2FIJuxLA+/XpMNVj3yfRLcB4rqtAlLY2+jx9XxIVCvPGiJr36b3TP1N
woUMivtxpHklrqED8IVm0Zjxr3ZPnlcTERdRct90poLGuXrg4PzDdH9vn2/Sf/sy
CII/WUaq2kZmCu0/qbZk0k4KbiLmB079PC/e0z0MEApql2+6fMwRuHo9Z/0ReKo5
nnsrefFBygHo/wTXBoKqpfx+vbEPcWzy79pCC20esFDlb0ZQva2nQXGBLOdlczbX
QngqVVs6U/2ntM4dGUF3nIb7Ey7gion5dhFBCjF1Uc7BUEGkwVVDEKqr9quuNgWv
OnXGUeroU2lD38beg12tONC8i3E3Xb2X+fndk828pWn7G11FDoKbArjO/7xFvFm1
iTO9y+2yqlIjcrcos0et3Y9wSFBLCdzeUkGAIVb4IDVE8r9UBgFQ8cdmdAMJV/jr
3ghgdt5uNq9v5LPv4EiJV0omFksGdABX1kbvNNTvQg/AAB8R5/yHA6YERx38GUig
3JfiAK2kRNCawMDuuFFIf/rzN3Zr8d20VTZ5vZQV0oKLm6QSV0jyPWHy0LMF5roU
l/WkSSWUO4Iy0/PSR/9idSqxd1oRc5gPHWJtB6MO6IlYrDBvZCjGrGpFVhKMFhcm
weAnAUAt8p9zf0CRnBBp6nlsnoXu2hpNTpMaA7xLXtgYCbuWx12q9QMjQiiI5MuL
mxQgABATuQN/7zxSwQBHkQxXWX+bGj33aSsBc2v2cWNBEbLPA76yYmc2pnproLK8
qO78uZjOFWXwyn/wDV5XRhV+d4j4aAIpPqtoD3PVzm/LlQ8ABFSz0TxmmzjtpiI7
2cm2Ept8Dw42LlQ3uU3F4EHsoW/csiJypNGkOGNvFRHiGJb8v58Sfc1I5nsapina
WHARSRuaQv00nhlvos+RvV3UGgefnWxxsLyjVP6xhJRxGcj37+mA0sPIRvnEcpvY
Z5kLkSFnaOEySXugyN/Lrqb59IONqiW3BHDFoz1ijyZed+6j0v3eD7YtkUH0n22y
+9N1sb+hBx9yku/d2aimIomg26cjLdnsJPxZNPmw0DqawEQuC6epUvfKZIfo+1oo
QRX9A0rcpOvpNiALrnOGnAbP1unvEYSmxfyoBFsVwwoA3kkTqYnIkW8p99QUEeET
KhD5sbQXwE7D8516Ag47lZzzxxslg30l/HGTchQQBOYmDA+U0MsO3WRsnHCpi5Dy
cQqCo7cOxZ8wvkVDH2iamqRZNJgu/be2P6nky7zP9btJ0hXLOkOdI0NZ6nDdTOWR
n4dMWmThAqrc1LYo6q4c6V6SuH/tCZnmsJCNce8TeZ02h80LVOt1+sDZ14GPkRq2
w77l2KiTYptl8gQVoHmna+n19G+bEnS5zQYkzylCjEndT75b0Af8xPIZQIXvYOjh
cXdBvpwuElJF/p5RyZvr7ddaD7niRiQe2xhevEjZOtu0036TkG34943NcequGOKe
VukarU+9dYwaVisovbpjquzz6OOv6rv1W2cJjSK/uZVeWysZ4m827aIaxwgu/j+l
G1sLpJxRZHSTfJhuyTin1WU2HvDnCXl5T1eCAJo29LpwOyVxfzPb0HLclFMhsaL/
t0QqP6pz1VJ25Me3lHb++uOgP/+79PbRMmp/PSE8kdwfvTQPEapKFj/WpAISrYta
MVIWHjYOKXb392hjfnQgiz1GBnhiRyauinA8d9/belaXlpQDSjL0liZpJzS/xdy+
eqoSSJS1iIv1iFdIQmbZFhdn6DifALaOxGKxxzjBWHUrzGDjRGGmq5M2JXqqWQZx
dp36hINY645TTXhoDiXMlYlGOdyd/5ivd6qPJlP+AoUfmtIyRecqf8ikN39hxbrG
p0wleTtYi72VCPzdDWu7Zg9VzmElfaP1/V6CmUcIPHNtXrN5PlQx+ymHg8LDimCQ
jxidjeeMQw27tJWYpbIiQukcJSP+oxT4kLJ0Wg8fXN1dL3iBKCTs2PLYATOJHmUL
pHwkBuqYugp1j95HHpTN3WUMHXQU8PS3GDObc6ha5fgD8eRbX6Ph8OlwOrpl9Uub
bOlD1fNSbbHg+e/5PJ+cQQCwG3kKNuANb+i2N8mWS7x8wC6czSpNdmWf8An/qvHW
wSt+iQLg/X5C8qYi4Skv1NHsXzOcQZyAFBAF0Cq5WTLPG5K8iWrTcsTmXwlL2tk8
vK3SyOzr0yaV3n18nwrihdbTkXjHH9V1BTlY0TcOtBgZuJY7hAcdpAW/fOEVIyMZ
0lRqPOmgqK8mMCcUqEWXwnwC7Alzqm0wrFtnZQbkMQxgYo62BfddtEBRj0CF1dQT
r9/moBShAMuonmem5QQQqbvw+oKlID/0KgKSUYKO8b/n5ax5y3tXJjNSfdbeTBRD
NYaTCoXDKzUgd+1QQCyU8kHOAZPQP7Rhnn0NMZkR6IICO59vSA3j4qf452dhqBT1
D5YZhbSux9BMtXK+3CAxFbBBTo3B+IUIGmClkuoZwe9xv99yQrhq4L9X6++5Ooht
9bGSzZyQc3g1sXpdSZnKDboDtObYPb7RDMB+nS+0Oi9ENemZAxBYAuiOxux3gqsZ
BF1yyBVFpwpDRMh6dH0H7S+nKQuocnX0e5VgRj85dMCl333ic8ZjvW5xZU3oCZ4s
TcZ0DBwGEzuVYBMDmoQq/+kOAdmxlaX/UGBMTJNUJJ5TYGcyseFTAEV81h6B5l5P
aE1jnmpZ9Pq7EdWoYIpb+PeopaIwhl1y+gOB1I1UfuOYtSCLNMtmoo0c1zwqKXmH
IdywaJTGnzAZJmqEp8TAYjQl0ONaOjeZw4Zmvul/LUKSHxSJmfvegDSiGNSHLqGJ
O86BUhbDT77p3jcLNMjLbwZY9uo/dAUYZxD/I/HgiD8vESdMZa5L57/dJKtEmERX
/ghP9xD/xMqLbbyiSc7aZ3p9WmZLyGvuyf3ikXGw+wiK3Uuwh15r6HX0RCn58PQa
wHzKu8dLB9L2PwJKjPESr7JiWb3aF9SY0cJuo1EKX1cRycPdUZCAHf21+GgFI6/p
v4rfIUeYPbs73ozZA4WmNryuh9B9YKUYGbKMwHGrUpIbrV3mZ6Zc3f8Aj7o0iPcs
nAM2sVXFUICtOb9TpM9vevcvfkZmDt9Z/NallFhGdcHQ8Rt2vCjsFBRghIIrxAOo
eo3zKGmf6DbbypLZmbXE36P2jORYQnS7dFeMs4ze4/VFzcDb1o28JpRkczCaKnQ4
lI9PACXqiW6hO5KR16uPltNlgotkjhZ1bG0hyOU295MtVUKisg1c+0gndbVnhumC
XaZwjqVsR6ULacNDv2YkJrsqegGvBh4gTSd9XuOTtoEx6h6k9ghOdsFUsPm+ZUDL
uFx4uLfu2mQn9tMAnB1hTSWV1hQXWP2EXYAuNQypBjpUZ/1BffAc9h20yERXZM0U
wfXVtYF/x0O8QitLVZFoQ4jxJoESNpOoLnzG9FU4fp+YNLcZM2GDZIPpUA6nnMvJ
K9JREF9zJxZ7eIMFMrlShB7WrNlgIBrRUhHInKAnzrTy6cTwQj3RVrm0qfSBYl/I
5PHKkwrPdtBGiSpfnw67N1bBoy4AQoDw9g9KDeUG1SLMTioM7pFwKBwgL6l9drd5
P57hm/gj44ZgUi8scx920g7+J9h/6VNxExUS27WuDeMi5qYHr4n+VD+48PF4UaXy
ku3lWR4UD6L8ZXDLgfZQNy/tdqSem/EzsbbfdnWAkmJGr3LivCE3+yT1um+EPIzZ
5bqxvcaiSwnhGxLBoh1k99XHRigidrGzyM5asPVh617DHeBj5O+C92O3IAIoYvoS
vmItoXND3aXwXKk6Sp0lsme61I6BQtViaJWI4Bz2lVw5X/44MrLSVNbsbDQfbnVK
ValbGjnLrSsPTrm5H7oou2FIqgNV0J6eekjNiq/Mp/0mk9rN8NmCeyeSqMYSf9fD
Xdg/IvfHgYXzYwbA6wGZZhqyccL7MThO0qboIBCPej0B2M7mumCe7Gx4U5MY7hlW
yEMzl+ka4eHMU5LkwK1PYMnvRl8gERGxE4wVEP/YpqDGc9voGJH+VKRs0UE0VNgx
GzDNdCOWM3sz7bBokutjbYgNexTtWse74MfgNKdi2L3zYdQZwnjCb7w/+/6QT9b8
RTAsjFeqQFpHwAGvGD7VszS2hHGkeYoywZJd3KKJxpUuQGsIaduC87QA2HmqHs1Q
+r099kP8V0YVBNxy4S/G30M337Yoj5zfda0m7gM2oRkgB9Bx0pdtFHLGKz2KS06F
FIH4tQw+O0ceyQSFiKGNZFg/XpAh2QSFq4q+gge1Z38q3xaz99Jcodt166Q25H/d
Tmut1ujOlFHXgB3tA6ZIpAmQXPhXpvls/3U8UuERCsHLzgq4yh+v7Re4QugAiFd3
JMoCu4UJS8Mrrgym9dsD/pYpm5KEArEUjw9BZWT2JNcTXH+DQgnW1v2Qq+K04MvW
tp1hGdvCMqioqamulRppm3W9bi6sp8Wmwanh7tXMFTjouoJrduRo131EQ6HuJoOO
hnmWB8upFYxBg62yyZgJMOlHu8NmpNkOEiFrkLe3lmZ8rXHAdTFNt9vfBfP7grxn
O4AC/s4xoou6tccvfyTNveaR3MWVz3S4Cuq5AZiSq9SnS1EsU29kfBIEBDbr0PaG
X4VB9nQ858hf/npYeX46eY5CB3qEOTZpfFrO92/nwGEK0krMDtiTzkyrYXKGo4dY
ryvFCZzxZoSJO+957PCSnsYwUszI/xOWW5o/IRMZ2YLErjAWQURPUkug20VFplfz
6t0qDfCzvESJ2RpryZZ6uMqdWOHbIfnbQdsYFlipH63HbFXvcrixCthKlReNyK6S
2q0dqrhSyk28kMdWTGVD9s+yU9t8DOJBFCLUsM23MIU6rRQdgPBJIljMXstxHSu9
pzCezUAsjq8mH7liHRkSeL66qCeQvwaHEb212iDdNe4i10KadwZPsDR8/5CDCW1K
737cFCVlmFxiicf7xfPyZBR+NzxM67fLWGPyv6sYuIbVfooZVbKwhz1A+WTwKqdb
2HR9FFu9SOwhiczttXBuDicW64pxJwHb6Gx5Od0Dw6f+6DSpw/2xxWq28iUCI9W+
P018GIS+9j9VqlqwSbRlCZ3IbvtYA5sHYBAYz4/SntPSQ0ifVDkXeotJ4uAoaqjl
AYRPJudbjGTwIXOhhG8eQXbAZ/TxkQ748J6k4t9n7sXpsxJGTKPfTrBlG0qI+7BW
t+kXVfI186btWgMoIB4sAvJyTh+oh/IRgb1RvCahtVoczm7F90sY4vDH6RPAgW4I
3tyu7vAA7d26CRH/22iSiMOAJj47OwhcOZe8rhFXWhgGWfDtxazRcLq2ArOMKsvu
bHfeA+PYpbr3bjIKTJLeOOMlSpjCZlQzI0ww+g6ewMD2lzLtF4UvVoa/94tJmTcc
YfP6bHd6IU7zVhEYMs5tj9D75Q4+y+LWiwBL02+5Qxejek6f7MY/UJx9R7YlT7PY
z/E6uadDoA/Q42ofPWcm1O59Fbd8iyMX2Ha/4ZqlpdVeriFhzvmcja3low1yW47o
vb8cKZJOAbBJEZyFiVz9t1wSiY7y59I5pui8kzu62fFhFeU8zaCvOc9JmKFvF+iZ
uLj1mVrdFupsR2Eq9Yk2navyEbMl31T0GSNNneQYULA6clIoFFVdaAaf4hizHF+g
qzHc0H4CA4k1BG4webqwfZea/a9X3Dzu2TwKjIVW1DQMHKn0YL/qDSipb9MrH5te
yzxM6rCDLaJsvahMkMtPGwNpIEtVEJLaL562XGWctC8U5oPjovn1L/67KO6YDtAR
FCd3nQXR6xmsZgE/Jk0dHSXxdB4uV5LaQRgnl+cTd+hdCPDI92GIFfBNvTKdcfm3
4zlsFR88RLNXQ9K2B5YFStlcWpEuR31S7NEBrlgPsHxLfejDc5H6h3uyEiJ9WuO5
kDduc43/q8OnvNtmnkYknXr9b/zrdxgC8IBm3FDnxuEc3f2+9rMnYivJofIzEGNg
SsVOiWFnnEDOwUG0jS7RvZsu9YWV0NZlTOe8XiUEgMo7h6EOQZYN0dyOZGRBGbhz
CV56JtWNGR+TrLTUudf4kklqfvX+kOw+nHZ+4SxAHALQBBczDVwus6LN46SeJFgy
nWUXZwcADtORB7xtR3ZtNvnSU4qPtXhaKh2L5eMZasld1hRWKrMXr6CrclyOXYc5
o8uVE38iIkX0aMz54GE8tSICnHsXq6ufIrtI3rTN9DbUmC8znxOYfVo2AakeFM/7
59c558IRY6CqH/4oBQ88DRw65BVj5I3iCB6Uc65QDq1JauQMYVxaZe8y/6nd8v1x
3ZdTWUGKa0l+RNW+YG1xiXgnj88nIs7RM2eWeXMj0Rnra0GKib1/ghHU+Aojcnxs
igQuBoyqVpvscdxlcXtA/9XnlgZUhSGZJ9AQQvOuHXiicdqDkQNMiio+s7HqCfDY
gePjjpnUHrXnVj3Lz+p/A26k83RgwlPO6751Sz17yexrPpEprz/obxmNtIAOOwrg
Hb23hmMbAZdfSheiDWma3ZQ29ZGdMjJHuIyphkEuBhujz5/7Lxin6g+gR0dP3Jhz
RF3f+XLvNUM8fvQLu0O8Lb88WH+E+jXGkYhlUG9F2AEHqjCNtOepSU5PmDfcKy/s
jYfPdcYN8YnnNbmGKRjZchcHocmYq3FLoZ5qNANNYTAc7s1fkvsdKrVK1EJ21S8c
2t45hWJIrGpQvLytK0w9YgidBgzlqNUHlc8ZwQIObqstdrnaYcO1OLDFDa+hZird
StaAy3h4ThGepejP4JUW7gfIvebxAdOM5qZ1YEdyVlcIeYDnHJP5uYMYyTJ0iCkv
oNEegSdC+yEXR0sCyRW5HtnLtlhMiVJwZRT5Cvjk8VXlI+3kOwVGkNe0Xl7opSrn
fQIxjWmDyzDH3vhqTbeKlby4hyLl3P7WGNyoCTG8662XNvkhpjoa7v6NBD1JENaN
hl+AiNVTPokgmwdxV9cQShWjUZHh5d9NGbhMqslokizqrSljkHVE0Jd7Ig0hHfGs
YsyjGLT/wv4BBGBebsGSLyFgoh091fD4IJu1rbc9L4MdmfL6HaNcxQOdCP9/nNaP
raz0etFLjgbUwRta7ywggKZC6C39cQwhIBQGdRc5ejEqs6wjF7bccKLQVNKEKg2L
05K60hzmFH6EckZA3QY0JCG/iz06Vwf/yvxWyoYgXNQ/hZm8ctRa6F79SJvmaqpd
LeTzgZvGqcdiur4F6KLZ6+w220R/qUJWpsEyzKUHZ9yqer3n6N6295Mq1jrMyZr3
7g04i6em1NovMUk5OjXdJjas514457JxBPnFEin3WZpRxA1il2ATe5/Qr3tQ+JAN
yb7jBwjfHVWeVy66Km4+P5ex1Ikorlo2L7gWRFwXJburanJUhUtLk87q8QLMOyGY
gfb9dVY3Oe8YNnrZYH62pmnsv8cpFvi3nRUqi16gWXmDkHzqmpq2w9VC0pXR4+uY
jYWWfQ19MSrMu7F6qSxKKRN5xjZplh3VBI8YCu18RL0wUIsBL3Yzpce3tQqBZ6eN
BM+9iV1cOYYF8LPZJXLfqqtcwYtnexdTkyp7mDr7Ydis/SHfsnqEX4Hc3PfTN0Db
TE3bb5I+yul5xhb+6M4aQbRBsqej77L4pSXpCiFmy+2CLCz9W9s+f0AApSI/bL2B
UCxgdvNwRGIV59jBXxVaXMnO6UboWlatcUWgqyrNtKM/TnRdsh0nadKJQEhXEz+/
okmCdzps75OUJqqHjMFkEwrueZIb3tuvt3omZR07WTJx806SzEjUCAYga27ml+On
0/3wIq1+YaCrgrxI3wtDJsjHAIqs7efa0W4mSHX6lJEkuH5GXMI42BxWmdyJIWaD
TXJekmWUz0d4QpJ1/NrH8raU3E0G7sAIHNf52xJIYVhxgbtkLsGiPyXScS/9u55s
eRuESwV8f66xXkFCc0GYPe1T9LVtQyKbavfy/cwVaSZGURB84jpKnq5R8cq0tN17
4fwXoiEaZAaVQaHm56ZIH6qQw12X3NMFwDmnAodBfjIDsudXreG/T3fhKy3Rnx3u
4iHZSAYQTOa0L42U5eKtlJX3YdF4SZN23Xt0MyDGcP1RvbauPD6hqZRmdDcZGS31
hxsrXHqVqW9dZTv43ZICxXyDWEx9oaqWPdKdK1Fz1nSb+Xv3vYhSl+IqAmlhHk1f
CvFZiDP+4BPbHzX/S/3IKLkSrzPr5x8nXvJdIsQ9BTd8DgFJJ1Ba45yLE8JjCv3X
HQtbskdmx7UiRcW48be9QnckDpDFTrb8ob0EYD75FU1hzbnS28T0bDMwW+sTRgb0
GcbKlRbAnpoklASb9xL7cOKHH/gloYNNT+YWnExL7GHrCnU7gVb0f7peVJH4R4k8
+YvATjjkFlgUYEiRIo73CewakoAv6NDh866BIbCd2M4li1nh/BH9TETo9pVFKKls
9bcbIWpxXlIBH/0Iokqb57EFf8hpPCUXTGfm8BGssrZXgSkujNHXjVvgsk6Jvw4c
LesKD6Y8Jd0dNLC8lw2nHDQxuJrpTFRH9Cqi4ffoQNTJmPnNiFW0uQbZQfANkJj9
abrFgEzM05yCTL35rzzIth/uDo74EBadvvFC5qEQ/WSkvwzmBydQ+bYaTYFeV+z6
0YdkBvHfqKsvefEH+aSV8lxJhEUuL72/reoRZOyVLbgqW8zqKJl9t2GwQYK1i8Pj
M0W5CYTZJyyvUO9F4Va4fb61+W2sdBoVFVACi0OG40Z/EJudQ7a59HtGLsXo48HT
2QU2F9b/LfvABiEB+WIN4HOGI6iBIZIDBaVKT46YKPxEGB+rFADAQf33nVTnxqTn
Tjix7DdmnauC8s4hLs7ArLnudDseJ37mg/+mkBXz53IBGgtv34Tgj2DjZenhnZNt
bW3iPNmLr0FGGD+B1oZZNI3e4LC05EZxnx5JUT9vlCLAACRvktcF4F7Y1HKEa5yw
W9pBJP8jvKOCRySqDfzYkFQLIDZnrhw3jwis1vkKEgndNKZm3B6Jn0rveHp+nAlZ
G+yVzhIaqHFwK4pUN4H93XW9Fvl5vD/UUu3KguEaj9gUpfCjG3eAhK/Civoe0gUh
+A8+e949/DKbHODaYxPERahwN2XEqTkp3nqBWompqgNgLICkrDODkm+b/NRSg6Kl
FpDuQBmsQOi2/fkwEFY7hNfyaKMMeqzJvaTIwsRteNqwEStJ5bw1cIFawkKxiV2j
9WZDH47oiKBeAjgv9pIOGlFRrH4Pt0Y19pHhxGoySHGFp1ZY07ujDOKs6PTrVur1
9UVg16vo/bVUOS/EJ1EN+b+f5NSInBhF7V9k0TIw8qY8MIla4Csu5lbV4OdXoXpd
Z2fJrt3bvGaoFgXf4gCrgt6Ap/srH19CX1FflKOtwWd2w1RT/e3DRudexfDClyO9
+X7OmoBY276ZLGQnZ7Kp+BvSdeC3IunDMC86S3OkyI4V7sNAZHJQYZpCP0XI6Od7
QD6/HjvXYO7qKcRL6tTU/pp176k8VOyq2BJjgw4q+heoMOCQJWjFbl/2zclkSDR8
x3eEsBTzA8YDT7HrrqRiQr0Q/WsIqLcUZ/jc+Ns7zVoX6VZOxQNsVgdFnk7RT2d3
FBQbVVADW6+LgSRRax9ELsTwFFpqDiYFg75mrQ/3GJqW9d6FKiUkOThiN9KMJ6Y4
JVuhTScH4vKvEwdiWbltyk35PROdcSmdCJCDYZKq/0YwLw60H3xpSUinRJvbixAe
MzKdCAbTS4oQNfG7a6BpKeHPtcuRwOlLTIGnmMMuuzDeQVWfWTKx2r162cEkJqE0
SdebPrYP9k9JyndYzVyAA2ZzC1kKEZiOvtSBUpHTm15CdXlQ5q0Mv4aTU3L88oRQ
679lKYoSxDgdEUCdhzmSRyhA6QbccWmyETVi+CgwsWdb71pa6+lL+SWZoKax8Y1C
1DCvDxOgnzzGY990IeYL8SARh+1u3rIgqDRAVwWiR2e7YdaxJOSCxOQoNCEab+ZA
Ls5IRTx8PGTzhGcOm278GPCXXYw/GM/YBgLv08hI1nP+U3tdb4ACbzeFnTVe4DE7
lyTkimmKUi02L2LhG1r3Va8tvkuU8pLqLCnXtYYVirEX8vSUbompL/FIIKmE8gcB
zA7OaFCL0kvmyDbrR/rozCQTfCN6RWDwnj3ilOf3ZtHSw00iPcpUxPOZf2Ww0Ovi
lO0+EVjFXxa900CcYBptqvftZsoooDaQeiUZ56s9MaV4Xe41kb1qf7jbvpan+pnj
jA/+Wf77WzO9ljlxW/128yL30opoEXgXuds+jKSHGowL/DW1WIaMYZqX7Fh0jVow
3kuLgrr7q3JN4aw2iXV3t5dvaXxon9FEbUOXUtAVtP9bW2cEXrSg2qv0mWcnzgLu
uQB49nbrnx91SoZMmN6GSG2oZP4AqMvAk/jDUHG0b0uUbppIKGZ+fOqcC/+D8IuX
48Zdb1r6an4JYtgwyToxJq4KE3qrwXSWuRnXFaNr/2vNqjJQd6w08PChIl1Rzver
eHdnK8lB9H96ovZPz2PKXE4xl/WyIK++5A0aSQbKRnP5sezbSm3sqfa0J3D9SB9a
xvTSiztSZgSq0MKL4Soq3EHGEUFpl7py/VS/1+zS2rbQQzzb+XD6YCIoLnpEPAaI
vkRjt5FtUzpXQjgV/NzzguGQZRWeQ70DfzPuAGPr1yvDUtPANaQ66x+9J0vBYD14
Bstd6QNrwPZCqPhONKccALoitZC6g4vPwZR32aLAJa19c/jQtspf+QsitzFn6eUX
QCQLbnrOMuwxhyH7ydXDi9czhyv8QDiXBixH+gqx8/nN26EtaZovcs+7kcEAJvns
gZEJUFIPLUtPaMRiLvaGRurlehBjbQEIBYwfx+IWH/o3IIulz30pAg9DYbBGvHNa
jRU+k04LUYnJoK8hLKOUUOwESzJ5fYMGDWTCcC4AnyeRDfitOvN3Lf29UEGgntyP
JGh6qWy7qEYxePyhDlZm5JMa7JyV322lKrcSroJhgkfwdILP1Drij6q1y/uZMMmM
77NkcKSXnvO22DME2GTjggrdxzRnE7L1xv2CBiDJvZPKRQ/uaXGtrnjoTrGJNsgI
nLd6TvQwUR4pkNobQ2RMDSYSPh4fUiX7V/iVRsv59006gsH7gh2vvoac2/fl18RI
pBA7yeQPpEDB5IqoWhefjtYE2YtghH35WDUsL0G53QLx9WK1HO74z6S24FvfN3WU
UY41Zx1cBDJDS7E7Hwns05DtCBpDe+9JzWMV87zbnPcpX/Rhe4NjePfRYfYkYDsz
CLbRLy4nSaZbfirPSLisMWF1i14dwjj0wGTfu+84KrpGygslpUJOD0Gsveal0U+d
8CO4Pg89uql2bDj9VsugAgHh46Eq9yyWh/d2VBuCTPw9yaSRmi8bFZb7f/tpdza1
zVzcE3d7HbvAeM9ljbDr79reXSdZjyr8nN5PuIjZQTsI/WGzgMU59HF9/qWrZTjT
FKPydRzrYGxl6jujAOtj+v4JbpJZ33BATvR2hzVPy3CzoDGUI9vc83jEaR06vwzS
S7pNGzS0/Z79zACFJ++AgXANwUKYnANnmEbE4kw61x4a/7oAJ4Q4epAauyhfqXh1
fr6m+OHOt4RgghX8IhGXrWWTzgmrrjFjIiJJfziXkqqVBdD2N4ci4YzsVaPAUAkz
EVxbXNvwq7B0nojjgCh6qLTOuvzhTCkJ8YJ6vDfg108K5VJoHQz+9PHAHIfM5dVb
HRDQb8uEPqix5Ztny02QXYmL+UbrIt77xGxbxLZ+dxJDdKLk3qUBRXOl9FkSrNXv
yTm+wWAtsmmxJXqKMCSFz/zu4u9c5jsiTDU9ivTAm+m2w66bRSztIkQjEPGnM0/8
TFbJlp/+zGa2xYUOSTBiTpfy4zGwAPfsdZMA5AIpX5vLLRV1+7uQcuxnk35Xv18v
5CvRRMT9OVFl2ElcOOpBOahzQeN9CJ8sbnxNavVZCt4jXdcPAJXnJUAJRCUb5Tzb
lYbMw5nhzTudXgHQ2Va+ui1yT2gXNITx1zBZLAg3mhz1uGFjyn/k6qDGYE3o/Vh/
wrLVHe3DGeVyxAfDjYF0GoumjjTs5Jz7KJN/TtHjyDLd/dIwVUL5WIF4hRhe2eZb
QEAVTs3EYMGMHTYxHC5kobxJeqtgIz0kVyG757Jw3gb/TUzmE6ZEH/DtdT21N4BV
y7m5SMuvOAzjzVF1OQy/vmCaUNtiNsr3sF6dpGPyAafPNG74xRj/Q/ckYDjBHNFJ
E/1ZJiTScf/bXNGSINCjKCYjRcALhM88OWlnnOjAOMDtreol8cTma997bYjfW3sY
esdFJuWDsYn8EQO3XnEmkb6fafdN2wpzLJwcoYtZxkRrvGhG3W27liN1r5H35Ajt
3MwiA1LQ7PhA/gC3RPAeOYY9SJbvGPBR5a9VKSpPXc/j+cdd9lsSejLpt8S1xDox
WrdlH0DCj+dJv42PyBJYJeVu1/856NaOZpjAtgb9CbFgmNgAFJAdeY7dZtturQAA
3buybyAYX1Fvn9dE42/Mg9uqhRNcIi+e6MNAaswTT5iKrKkw8EEEnzF3TOrebcpr
kYld+3vf2HFJtDh91xo+UWTYDUFYB7k4/BtP4h3nc8jtBrSgDnY93KVM70eFw8j8
DgWtuZ6qyczeXdoKGSpmmiU2sdWXzqRnhxRUcH/mSsx0zKmzOFeTsdwUu2thYqrl
Wx/yfK1I4q7gn69sbP26rGQXqp8inzFbQXsWPcRpTg0cV9ElrHU7ZkudIy2b0epX
+Y9wA+G1Ucb1D9rQ3mFBN3VE8ocuV6pTPpP0Za8DDAZRPhCumPyrXhHdyvunzjTa
b1RYfziufLDXKbJEFJZgEAmJmXtk1bNDZr5AE654uzJBBuORoXER8yu1D3qe/T5B
Ez9JleVzb6up6Co7J3bcq6jETuz6UuQZID55tSO69P0uRDtDl61hwL2HYeiCc0zh
L/MfsPsnufctlPWG2uXSSJcYiMR9KQs/rjn+wDhTBFW5Iy9XXKisEGaJrR3EiDVi
ciSMR/sRWpm3ggIIW+M/Zblu5oK1VA3wHXX4szeSzKRXJvYATVXME+aGegkOdLmM
njdVxE9a1zkdxvDT2V5swkUXl/Y0QKGmYCmllWHmV3M0ZbRcehPIsyILY+UZbvfP
p6KRU7Bpc9FixKEFLzu05PTG/mpvQzAao5NR49BAqPG6sB5pMkPgpi9Ck2QYIEv8
/tm/v1GLgPW0cSAetilmXG0AnhPASH6HzSR8DBLgUzFtNn0BUPiAlsfegNvlAw5W
lxWKu+XQMge75KKtTwZicua+rlR60E7idRz5lhSd9VOFZ0BUgzHd/n5ECged5hKF
fzoMLu6e4/PFT1/BZNYXbHwZRjNF8vpKTuutY4l0vp2gzzatJ9s3qMtWsbORj1/u
XyoXEttkmBrZt8MqdO6HowEjTfu9PqOtzwcN+WYvcY/jqgIjhjJiT9DoURuspw6G
PkrLtny+4iRQ5RnR+HIs/EkxfiT7B/SXLbzFbCpnfB7pYrXDB7TvZNl5iqidgoqo
q4byxLJKNbS4wczPZM6jFaJVOiVbXg4X9B/HxF1HOr3D3cswyTmnayzdfcFNd+CP
/9bvC0zHfMnXSv69iwWKVCVdbtpjwnim1LW2uTjkC/8Vx8gTrtJFzwLIWgpb2B67
9S6P6uwN0H0//tDl5cg97POwd1Sz8Wk078Y3BQqvsEmATKUD2tLAipk1BCZVh/Ag
UhRhCz81x4kC5mHhTsBMkCbGZiYNONHY1aLHHCpExDos/bz+7JjoRKQcZs8Qgvo9
iF7nvTVwRlwg5vMuOAZqobx8BB/vQYy7jpTL8jfVH5+jCmpPumXqZFB/26ulC83R
ubEIF/9aWuMTnkLTgGWaLMma+ci0U7TvIPMdMrG4NikX8PkEpCJ2nrYthYTkKS8w
/OdpqbVYCZlFyLtK6mQ35LCI81SjHBf/UAcCP1i7j8a5L66Wq9gC/biKxH4I8jTF
6W73nM/UIX54sDND3ZkFP0jytM+s4RkzNtHHv2wfxU3n4QeRijYkjlxjjejEujL7
Q1bmVIDcG4xt4fg6tGCmZnQy0pBtskY4qQNE6+PnAEd+dvImCm9m1nRbSIKp1qVD
8ia/XqkB/CXc4hBmJr4uSnEoosADENkKjPsk05ljPV+67QQTHyJQUTsvkvV7PZoM
GYj9s0j0hioolclE67/5Q/CjBuFA7zX8WX0CqTRsA1vjE3Oj1b8+uP8vZ9+jgrls
FLZICBC9+h3sOUuaX/v+KlOV4SgQGZKIYpxmxfjfuidfVvTQXXF7GNZbuynCg36t
drjNAY/3ja7o8WYLlZM5actkeb1JTmMgwAqmOu8KYpPFzfNne7co9/16ZgHOAteM
nzbOa6PJBhZTaWoidhVyAThcTnAIYHde36yHaO9c7PyecFSw7VB9UBfmFQi8OgyP
obNPHrTQBpLuVp+L9AaeEG4vUHd3gu976lVMSRae9Ah3z/zMVuooWAGjSCqWzNus
UWN71LKXvxYcfcPzGhUytMqIv1EXglbyXTHED+dxRiwHgDtF9+AnmLyQdmEVHXbm
3eg+j679aA0WI4uxsTxzZZRAmrgl9Hr9qbrBsKXxD5f8K8Uq0eFEusy1lzZDFu0y
11KQMLfNPAPzXfxpvCWSukJzt45aj6/yzKyHUdp24iIPWydRZ+sRZRYlBNlwBklU
WCFfTPO0Tc5ux7f2eOKhJKD8UKRQ7Rf3lo/yNNs5lrV0zZ/VBVlut+YNAiq5Opci
lY4V0yAyAZfdz2lSNTEHx/llYNUjD6qADK1JSnlGnusuz9tPZfW071fdyy1/dj1Y
/XT6x619+gynS/NI1jlFlujOOvGEd95Tk783eOoXppfndnwkXKRaA3Zbj8O6pRTa
mYbsFGb0335qY0oeO0mtg99bN/37VtZxty3jZa0Fp32aTscrHSmEB1qyDVDoXmfg
lS6S0mGrDD3X4NRkQFTEp8UCVLrSe0tdpyV2zTWbXpH1L05db8H/WLIP6nRsT4oF
65l0HgrQfYbM+34RMZWoAyuXyNFNQz48t0MGglRJMBu4dhkW6Hiw/rqA+/POZIgu
7eEGQlHERpf9KZgGrDYGLSuQMnyGGbH9XIoEvFjXXu2HiIY0SV9kCUNKZHgIjrwp
QMMYBSwjbPWIjTrbJ80CbUfW3wU0oEBq/GdYI4EmFEqnzxluzNgwEvwMAtiPkSBj
lwdWGTiWUJzVMekc+zCttTQMquUNO4KN8rHkwn/3+AIEog/Xv1knjRYDm+BUaZ/B
FmUkr9RaZ0MSM0cFEBtS+JlsBl2/PTfWNnB+bKFv33wufK8nHXdjdcY+5UyWJTr5
JHnOgGlf0RawrI30AdB8RbOqK+f5vMPku26qQXCZXCVu7rhFlFGHsUDfduzVLEne
HocozsRWt8JGwqZIE0TjruXGKbfYVYE9ysR6N4YxIJqpQRjNGy/8NzbDos1gN1Qk
Y9CngQaPSjXpy5l/7eHkuNiwh2ETzvm/vYAqwAD6pPkgVZnRWAEKiWJA5y53rI/V
st/1sBlvnrdiF+A1yoSxYyoWL/jjWNgEYN7Q9l7Lm0kd4agHb/7lN1EARMcE46+I
UmnI+nFBH6xlKyI2kz3HGoUakK4Ht20ZdFg+uUGHKFCeFUHesCbgtRhU9/VKSVn0
tGEpFXGUAK1VsVxZYoUdn05fhhuJt4ATcblItN4wy4kEVO3SvK2EMaKcwjHpZZPs
7Zp841eB+YHye2ABhp1k6uXGisJjsdCYKTyB6MlDvL8dq5NZTMbGZ4uqmnQYMCZ+
YSjidmouq7hYlvz8lrJfM0SRlUvAZBPmmaB77DBwVYw74KLsdXC/3HYZAUY/uhJK
TQvSNIE+aeVLtBGbF/rSi945XwvevuDmplSAFvGYAbN3HkBMyBD+54MqxVas6dx8
Bt2eag0VipmQFy91SvfWsVh5wLi0x9QeZIgrugf1ch/qETabFu1OGtzEmewzfNFD
qa40jB7fXiNBGCILNK8UJHg+daBbkvTyBHxqShpYYbB63TvL0kU07HfdndmK7D+A
//RipkZpX1yxNioeubKRQNTCH8/j0vLckeHfp8428zBeRenndmAsf/84ndwpWjUR
v2UO8HR9fDKRq/iwPTQdvCKPByVEpVnPkGwRDZCFnw+OaDwDv0gJ0cKsxAbBheoH
MUkkNYApg8lSI9CYcC6esl1drHHJQXZFfYMGnWwpcxumD84KSQwIcSz6j666fYvK
GqsVcH7AgEimgsHxv5X4KW3zcGsDtTeNDsaCJ6jTCEk+g6NyeY9BY9XH0rrxa6V2
TPRMFSbw8qGF2pxFM+UhKYsC0VkwPweMCZSHY4EKMK39Vi71RDDjXi9bNBKoF+jD
33gY0lBOb1Y2NIP/Zn/zabKs4CBR1umlfs10W4rpTkbWdxk073t/O08WEWVMrdyJ
1L2DkYC6HHME1SconpWnLbo+knRAl32YnKfiWPFRBrmYf/pbOkn89MxsZ4WfmTaX
dInZLb0tf1tKEl82QUOEvEvK9D9F7a/bIJkBdVBO3wBCU2t3+M0T68w48EZ9YzYI
CunNhydz7PeNEIkvqk56vtCU7yfwFKXOrcdI8/UELYXCo27Y8RotuO0dLpHK5fQ8
+PkDtmDJFvuJpkmWCTV1EOta3niooMrxs9WKFL+HQF96LBo0WKV65c+PMZOgFHqb
T0TAMJhpcgJ3QUPX9K7eB6tfiVmTsjceVmZuaQQL9nJjQLPWuFi2H2vtv38But1N
ozW/Wtfd3Rd5FmrBCDpqd7jBWy73/lKjOCujv2ZYar+Qrqn2k+RokA9WYv2Vx6PY
v2fLP/O2onH42oqlwpI6l5jlkoj4FZLt0jnEU7GcS5gd/TVM5mSeIIYqZRTv6XHZ
HE2Zm61hEtKMGYBd0V+Ru6z2rh4/1MChn4sFgaHT43rt6TDWqaZDAgsyiCGW2ihK
upISqL/6UBsttagmKyfN3IcooGD2it7CBCYNF0TmWXOqAvibNCH2zxbpz/JGNb16
RoKgzP62xk/ybpSrFu6633gUu+n3ZxcAAiteJU2amUCLjrq9jlo8fQwWQ/J7dSWC
onFySYBXw2bT9mz/B4BfFvmzxEQuamwWz8B8+ezbmAGYp7jd3QxnY1G2iqeVcJ0E
G2Bn9aE1A0O4sQekZnNR+HrrveW8CRvxQE/9BGosvYldBNl+eMAMMSzZOj0biRVq
g9D/ZZEDfCkMvRj1aut1kfiLWQSUsupVDU0fznWaLrWdL4kKXvzwFmjaoFxn64z7
FxelRWqCmjsIvFWLMel7nxwFmABB51feMVwkZ3QWqvduIEuiUpsK//oh6Ro2rMXG
4nAGRnELgxV9CYmxK7mkYEHvHMGYhQqpypNMkngs8XCqEOlN2fXiZF3Y5E1Tx3+L
Zog+3wFB6BMqTmysZHalLKxvHr0vcqwWNLt0pmAN8hBQwJW+Ks/24gQ0kL3kBQWX
NAx0AzBLNd6rn4agBxfFe9gL1/KZuzHftVTWyP+SJE9tM+YZEPbIaFFL/yRNx4Iq
+OfXGqRV/+peJM0T7Jes56F/m2xoDqi9/LZu/woe/6beoqzT1JTXMqC6FSvO8eYL
IrNmvr1C2TMncGQIYUIqruD8G0a/alGF1fx9CSkYsk/hoJiuEqqEAm5l9LBBk6k8
Qx7ZBN4Xa+uw5ebmBfeUpjaSeetyDNAeNSUsvCimSX3hQEZ2lH1t/r6LH8Vn0lw8
WKs7z/lUsmgpIF8rRuzoeOLd8fw7u7tcTO+e+WyG0bFWiO39cffpUKhG/4RGfi6z
AxeRPvPQxyVwKG5Vvsx0G0/MtQCLaxbft/0tTJCeyRXtB+1DDaSXjCyHAZjAfJ0e
xcG36LtmMo5zYhIYgL+oI/kak+0zf/qRHQROsRI4xy+Hg61Xv/M+Q36R+WPrv37m
vKJEYgLa2xPLXXzr9Dfn/9rd1kT84eAqNEUMxvQHDAxDPLmZOsDI8Os69XYVS75M
RUnVuQjeLXjrBPy4WyGfKsBdO6+2v81mWdMP/kayykUJZ/VdG7Iy1eAbacyaGoFU
7vj23pV4KsTRiNQr72CMNM/6xKiJnbaHWvmsniGnMN4OC9KpNd9rBU8BqBvOzmPU
O4mgyF/89PBO+UpSiuKESroHun68qrgOrQXFSQaAGfUTgrFXbDwUrPpx1b/1bqlK
m70mUSqw4vwUwjBmIiOFOTsjmwouzTmrTCIy2gBAPN0UE2QGZ91Qghj4KmBRRSSa
pgNRsjJJGkDSr9c49szH4Ahg4VnhL/HuZYVFHpygcIB6iwh6f+I7XnEw+qhesHbR
/t/hkEgc0sdEfEomePpODWEAgO9Hcy+mTrTs3TQLTD2xcRC/d8xgcb1bIGhkEGKo
7dAyAAaUKlMhrOIC1vg75O9BmIMA+xqPy5EJkQh5LSGEdagW/RpIByS6LZ38trJ/
VIPeMotQ8aOWPdBLOF80GDkIHhx5zMME/ONdbYSqioFefQFOOxMpfSP7mG4KICtT
QMMT4i4ac7XkwEl1xrmgqdVG+84HlDXYYHwcCOhFWGgNyIpCOEFOJ8WEWfSDZj0P
tWh3PTpyo18bONfsjGkds658T4VzEyII3HSdGmHIrKLBlewcHni+F2m7ezHJ50V9
Guf1+POx3mPAVyYaFdy06zBV+81RI3ZOMzrQ07HsQ+7ofbIZrnd+NU/kxtoHUfPT
Z+r1yQ6vPsJILt2uocYrjM9f+fBtI7ZlIgjoxzybgf7aHwvU1dB9nWrqC6TwX3Sx
cU7LYQ8qyhQUzS8m8KWtitUow2xht92vOkmcvzoA2HRjUSqmI0EGQbzC0NskibZX
Ya5t6vSYAsllxbThJPKH5BnVWUCJPEPm+mI2+fYo0xMMMxMeVuimKU0ZLaOPFzpZ
iWE4uwT3PeF24wEMahMB4DGZKjdtT7V4AB8A0vgjZhjRFe5MeA61/O7bt0Xv0Tfs
Z2N+nINuNdoefSyczwRAkBjK1PpPc2+ND0OfTQ0B0P3flsUlULxKUSip52scEIXx
ltQ72a64H1GLHQO8Yc/CsOKXo9jnyEwt1zlpNIGxtGXomIn8mJRWmYIVWVReETVi
yTs81gNzanbMKkPQqu3BTqq68nU+8urzZkS5nOHfvnig6X+jOQzrtpuBBw/pPNy3
asc1T9kgNx0zf7n+Dx601aYnIfKDKjBc/45hdvCPH56HnaZddWXH0zmEfIo3ENo5
boG1I0YNX9cOgrsP7vCi6Y6/yp0CfqhCMBj5S5Oyx5372ADSkbVAF7kuNWrPrrfu
jDn17gqqF0Sq44srJpU6ZqTrbUieJhkjZvJcDNKlTQOC9aaF01KiU1gT3CRsneKc
kQEC/Bi0sUJ5Y2GoUfhV0mnU6wi6dSeAx6mz2mcd7vkgqLlrWi8Hv2L1IWcxTIq6
vxcES3arL52w+t7aRIYcf65L5nbNt2of9GU1DYOLoPnhjHg1H8iSc/yHoMOEXauV
CwOXUKectGIa2WFrzV1E9TS4WN49E7+s8ONyoedy3tV0MO4CPG/+LYuspQVIaH+E
kZ7ffoHsWg9YJ5zQV8ilImBy9zgmU1E+uQXuXli9Ga34ByG19tMa2GKQz6f9Ywq3
nZQEDtqtyi5S5furXqsJSrtKOYR/mH+tFhV681mw7Lt+Bjk7MRo4e+fjeNAuqQCh
iERustVFnk260g032qOolFQjbFdsAnvGIyOVkuWkw5nK+5hFH1JeDhepQ0A/UXx/
IPv9+391TV1hPI727J9+F8sokmpDbnJWnbh76+xpiL9ws4DR4se94jN8YZlWIeVO
UOn6Bh8A+hV9MoQO536jUKRBdLMgyunZ69LAm0KkPXQn3GZjjcWeQcmIP1WJZmRj
vJB6WkBRXtGdfTDQ8C062PmVjJNRX8a/WpTeYIHpzN3KA+rqvF7xM6pCtcblWi4V
p1clIunIWYmbxZb6F7+mbmXPl43j1PEqsyv12jnme+ET0ood4n3GlFgmpNvDOf2p
JOxHdbafPYVvW49msjbl6ChFp5ZzrDMfUX20h8kJitEJODEXf1uf96Eze7s6uQvr
a3EfDMGH/ZRiQPrAjR/gwXdd3cj8jRkOD5yVYhaB/Zv3IF2s+9maJCPEZHwxC4Nf
jUpn0zI2P89VNscy5w4zoz1AT0qSUVKmu4JbG5Lfz76s99ANpCTaIf9Kw11C44i+
/BBy8slWlcyTlnFk8moZJz97jDon46G/sKoWZqe5oZKT+pzBwE0eh1pz1+DWM9vk
pRIj9oAdrbrrnOmM8sTYShNNIfxJsdvsSUF/yth9hrbchuSPqlwTXEswB2ht8kS7
sYovXTz/vGIDqlCeGUbxue6HtS5+Oq67xrWlh1hfI5A4U1p1iadensDnEa6HK3O2
bVqnju0krZ+AvJhYZ3dzxjz4CWsbfMb7v8AHkUVudQdvydpMeI5b8GzbYsSDvsrm
G+MYJe//DEkUPctwgudQA9cvzv4I+younRszCxKupAKS5D37cdyHGwJoKRABhl2L
fl84NXoJM1+UHSaaVt5yfyELVOE5q6JYTQLsVrio+0ickY/UBoOCL7C9mkpw7Gub
QF23LffPVHGNlfyfUNmJfgSHy3WmdhD9rxmX/rHvr5DuYYj6wBblO4gIc2kVgz9s
bdp8a4hjZeB9aPbMhtjd8k8HaKhyswshHQRJIJVHXlYTdC5tjt6TgYmPHALts1XF
I/Rz7oL2W3czDoW4kwMOMo+HFTvdJOHUg9BQX48g439NxocQYGqVR58IHzEOyBuB
gC6FIi4YUp23SwBgtcbGkLlMTwVjfWtE6csdbeNaQNaIGafXzlw/vIh9JwGMmSvO
3OoQi7eBeWpFB32PQvvu38/gz3aM2xhK9WiQIcy8dWn5cLSl1RjwW2lZKfjnCkgp
/jJDFnQr6j8J9Cjqoc0Vpr0woybOl/KhdetbI15eDLcqG37Om3x/Q5m4C11EH9oC
CpZvf8BS19gv9OlSkxJkf2JmK2nXZqskg5WdkB7sF2F8LYMQPS71vHTIYsIEEitH
NvBcBqdxPwPvf0xSzyt3Vdy+B79Fm/6T6tktMr4A3PFVx5XlZkfIFcUvoV7iHGwG
WJKy4LHWfwsQRhF0WdPYxG2LN0ykEeRVllueTqQWWNrSkheJuZ8nL1BBeglJ7EgE
JMcvSJPAPJ/bTCRKwiVjrTiacxAHU3zz/JGlaSnpqnc0bFFlRawSnW1nz2VgiOdp
ohEQOMP2/aqeinjlXKqQ6xIk1qZC6fS6p+DK75rvqAbrJ5MsN0xy5VAV82WL2rjt
lTkNTwsQrN5P57b4xwRhNKDxyQCjdb3OY8BMmPAVz3h1t5b5pzAru25harGLR2lk
8XKjkJm1AGtUDWu1GQDxL6SN67QdFI4rrP6Dc4nLlN6aUimpQupPlD4kiYW5cC8N
w/aYwhNCvfRXXMG/XlKRTYoL4XDazaADVz+LcbnBRPDyEVuXhTA0+w5BiryQgBQ1
qGnqQoZ0Vj8f7zsyrzLKMRJFf16Ji+lVNrWqhdTJN2ArUp0afR9xUx1RC54A5xiy
oaCuX8FJ6QnnFWaLBz84van6bmOHpE+/D41wOsWC0CzsEQNlKDWXCyTo7JaObMA8
nTZkD6mBCDzmn39fhmjWmOiMTnt2tU7ECA5ENQqjT9ou2ofq5e5l+FqaoZ/bYwda
z4Wuo69fhHL8WlaTuPgbkyEU1U2f7sogfhsG0wPiyO1hfelO+v3G2Ng79KDo3uvr
4SkzTP/bDgyeTSZDclx6QGkI0uK5npcGC00qGXN0Vobo7P2jvVtxs960wgDx0i0d
9OlaviA+VrSFAlW22DG0MoV+pH7RsEZT/rCGaDfBRZAs3ZJciv+1182k3BnZvf7v
kdgzrMbs4cwcW/9kWVk2JyvnX0qlAz6/O45gS22jxSY7b1j+ieyiDUzUsaPaW0QV
84eYaqJw4LtAz2yjSeal4ik90J2+Sr9MPa1vuLWJJ/YajMwRmKinEHD/cO3hPtBe
i6EaLDyo8LSc5fkwvA3LTpnto96VUD9X9ONf4NFaiKn12SNDLY63TC8Y9CKH/Cx7
Khetng7IbRP75CDBzVsE0+AfUHo2DXZUp7puCWS2aln/v+hmI0Jw9I6UUCqo0ARi
LI9tmUjESSQQmqyGsVzdIXPV7GTToc4LE9fF3zpo7OAdz4M/L+9ygpR7JDyBDSBW
eATl/sEZqv8P778tM8AM1GBEB6dKYgGKaMhenapjlOOe38PRrt6SnnIsA/WjdbeX
PWBykvAjRVR7i2kpCqucJCLV4P0vU608E1evYa1MabhhOQlQnp2sHm/nFZCMKmA2
cck5DRNghvyu5vfsZbWslzJLO0wZ9zszT3kSAw3K+817GLraaNhR49BAP7u0nA+3
/+einYcFW5pLOsbshGnWx6rXDwCjQu0UJIc6N4ZN1lFcsUtOclx3khKjoC8copV4
RrW8jf6O09elxci0rEc3iufFrHSDjPdCw990dKvkvJdcqj7A1XAeNdj1K/iz6S92
wuaEc1W3sJRjogqpKVtt9gx2b1+V8uh2/C/hdgPZyKOz2Of7DtKTg6VXFlwLIG2i
Ya5uflNDm0bDWtKTBwG/SirYzYRuP4yMY0UdYpDnEBx7aZatbSVYtSktV5l5agyE
9Jlx+WWTkj/z4/erTaqzUN63JLHBh5eY+RhFo4YomCG+SHkTF77cbI4Qd9MuviT9
tOsRE/e5inZP0gkazj3lp4Bmd/35BxcIJXcveGnK7ZAv3iMVxOzUnfwYQZqsQosS
ihpD4mXe7u0SiWqKoH3LGCbd8TR/lpZSYycWJvriA03eIfDwWcDoN1TzcAOwUpBW
aipGSUlpw53axS1ZV40DgvErAKD36NJ4NLf31TAasjEI7YdeqsHDC/9LrM641E3J
OUoMgWvrPVZDorlUABmEf1VHbgjzeSjfb0MDoUn1ukjS/DYFOX9sHAPXPHeqqCoe
W0/0pLlGuvSwqzcSDXgarYUlj9jekvBApZNM6aCRUZ7VfYuQTmXCQsXyYP9G/Gcb
5397fp7bXvg0DNKBTzic7ujhdV5VWdJ837Dpj0SHjlPtcrQ3M3uv4O/S8bz6b5I9
ILhXsu8RAfVnfek0fP7QexbI0c36DIwC0r1IUTxJ+moHinwl8LYGzmejhQRhSABT
wMtkp//w439iH9td5YY93pGrL1ZoOe+dNQLh/hp6UsuHTYnZgtu3crzOJG0T+3Wi
bqwi85OS6BHUJMCVfR44XJc4BPgXGP6LNEzguPqFgGknyP64cT4xdtrR8cqEsDgn
DmvN+16ZebQ5zirixN9Eu+UTQq2EeabKfecNBLnYe9+2uu8JBcG4J4r2QE6Erkdw
xyrota7A7Vl4c2J3jO+HqLxWHHYLJWfNYLapbnurt4pOiayQkbDTKMHM49r+4YLl
gSTKQD2w/RxnxT/z7O1wBe+SznvoKo5atb/q6huL042YoTwre04YClHGflNkYqzQ
Z0GDoM8K+34HH/tCISJVXWXaRl4ceszX/gsflygDqBGpLyVp4979TKlGblDARZt0
CXAoNjfoLZV+qO6IAC3hCaalGEGN6GLTe7UtmD5hCsr6HrnvH/ADhZeCb+NDMeQz
cWsdCfqj54N/MelEjLOP9aQZeFmEnpgGzTIf8yCpTluYOod8Sms3xGRIMXgw8qPZ
HfNkhqqowUFUvfCgbSbIyfrGL1gQ9PDxhPF0u5eRhe/2T1OJxROKJQBLzOw+fM8Z
/6VPVKrRXml1IeV9N8EQGV4KAt60oQGdUvi/an08nbJhZlnQnBWQi+EGvgY44i1G
wzWOv/pSkDMjVJ2qrlq+0LKtsdaMxoiHlb5tECpp0PUcfoZXUS5InNTci14/81lB
HRtfPuatfRZa0iFVF3ZpSMmBVt2zM5KMIosN4B4YQ2GciWcOpUwAXqeeZfvl2AJ3
moB18MnBpAF7H8bQ4g2YIaTfLuCrA8ty48Bn4MpZCFL/M+hHPRvG0/cir4JE0frn
P3J09TXvXOlO/XTplZYnVScKe25YkaNY81aEV/zRKFRuEEnc5bISqZ/scbhhVARN
7MrVobjekv5Fb1cnK3Uin68rzLH321OcddJwcmGAoHM3bmioRk+tDeGSaQLoRvC5
xnj3f8ii77G0ykkoJHv4CXE44kJUhA8R6xcELaumOXhOUL8dzXv7r5Job5mUU1r/
JbM6diRWiydEuRmIPRsZuNqEp5VbVY3YVtaF2/ck9HvrYhkPlDY/+msDnDfqe3c9
LvS31UpRzOKGjKyY08i11Di6sgcyTUbvm8er9Tp6VVRPFYxayvEtLUe1b3UehffT
txe8Irt9Ppfltq3fWVm1HKJw46hb/vJOdiccBuADcJwo31qr8TTMVgi+WTd7xzqu
U1NBCvCAqt59Ibme9dLJ5CY0rus95NTzfxuJsBIgy5morjiKd9sECFhHOQRYbAff
GfcPG5olPweoEMd6oMHKagoAoGyQiWf4/uc2fdirEPFlEgTYadJCZEyLnczGP+lz
dudOH13pGKl8RuDE0zhHRVk8DS+knEt1kQHi4xY+gfOzySWckPr/C1AUlZRqxNbA
iADgIv/LxODyp5MVmRmTEJO72Fs59q7z7w/qCj+tTX2GcIR36D8lDopybvChed3x
a55QnN38NXP0tUZ651O9lpmU++uiRJbcQd/pADrqgKFzC6OqJJSUY9if40vI01UJ
Q5M5evLCTFN/ifH3RaFIhUf+Qxkt6V2HGxMvOY95a80j3b/U5HhRkV1zLCmIJiXx
PXu8D6kJFCrE4E+XmMwdQASXO4CAfES5qbk0cdx2gwXQVRU0RL5ADOruP9dfcy1T
baW4lxxTS1FUN+EnWtFARmTcy6foOXqI/+u/izdXjiX/CZqdAO8iUA/6Q26lukdq
LQFLyhRaSZYYtxqObF+WiR7erQigDjng7XcNtVKSa0Zlj7j0TwbMiA9V+hzJEKRS
F2EaTa3PvEZEDq9kffN1QrsxybTAr1zHU+7kX3qtuH6n9TnQAdp8VOr9qzLuhhcB
sH3St/bziMJopG0daYbk51ypmw/fnyv6Jkos8t3PSBAD6vnBo+wYwXPRjOvHM95h
Y6QlKSMMhIEkVdsDN9FxwnTAXQK99a5ksvaTseewP76UJDyTExfx4Yx2dJZRQ4sl
EkGKWYQKI0DYI9xilAUV0N9ln9LNusp6ihUbUYNUwSunSMhVMTqA2IFG8iLL6GQI
6IsDbzlMVpFMq/xVOtYpnC+gCL4YtVh3Ugj9EjGmJGPpMJIIB6khJJv3aj7cIJK+
MZSngbPAWvey14MSXw9iFTIVCnUY/EpaxmGzwJfbcTB96xxz8zN4HRUSrGsc+tAS
GMy2bXxO184gCZc+UzMZc0G5vToclTbvcZVBJ/Lwt/zBMs+sJEwsvWsQ1rMpcy+D
lQBNCCYRpqCm57GlAJn/CBiSiUzfMGCH7+rUIK+4eXZCdmXxC8QtLQ7g8d62xO4z
/MG2BhvCwkw0GqjdTVmeljLayvj9tj3ml6BWE3FCAUWao7FLRgHkVOgHhwDpfXhM
JnR+vE68uzhHe7+p+04DDPAolsN/cLhimVnG1jNAC30KGyKof/YTAHYpT1JrZyO2
FhBEIjU256ruhRKyLclI838nmtnDnW/I9veNygbB9rdYMiw7U50cfLBP538J3OeB
09XsBvqvvV6T13UCiQhn18BZmzHDhJAr8GibUatsQ/ahRFbzILWXcunM35+YM4qC
30g+X7yBZCTC2hbhSeMPoJZKr9wMZ4lDu6TFSssIW4u0tAhJCU5+MWhbvG8duYdX
wZ6Y1RvSaNT60QeUnMJrxQEkVhs9e/i3UTrY8IHrGwzaKHPP0Jzli80H4Sym442c
RH0oDn/P4DsSZl6vXvr7nG8t+uUnW+PlOtfVWyVXZXCAysB04vMzaWz5o85wLQlK
bPSxxjS4yqdJYnjDf1rRDA8CAI+han0ZY11QH5YutYrEkBINGSkSAv6tlFlRrNHH
roOkv/GZ1Wsd2mtH60MatG2HA8iriMleL3/1zD5Mq4eaqfrr/W+Z/jqNfYXgKfKX
V4/VDzWUZKA9n8ZFovIK383K6f63M9xxH9a0Xc2A0XZl1mLKAow3Q+X4PqVHYqSD
/4YaktuT1IwYoRInoh4SaNrMwoYr16r7jYdtsW0lTcLKwX7HT06/eT9yNztAtPQ2
h71vrgnnQfFR0h9aTkmrZjYMmILvzplpSrNGqlySHPLQOMkhCg6N37hc2TDuUIqJ
RWYujsUs78mOroA0+uX5f7BtHHx/khc8iWvkdH5VlEwKJpfhvQqrZwmH+NQXb2HS
AqGeXsMMtuxbt/a7OPYnpXRTYvvh/PcpfuZFOllUzgFAl+46tvmt5QTUbiUGwL2M
wFjbBELlxM6UisFthhVkjdlTnCCjQ1scvz3TVgAVB7wKM9fpyyYNWfqd4kiVyThP
WWBmIGvzzBqosVljf9tOddZIxTTlcrYSKQ9UzoLm9KQhe6QDog7hYLc0EaG6ND5h
KMRxFvLK4GzR/KS6NiOAIdQ/8m3uXYf48rhk6C2+GyYj+t0Y82vsoXz99fJqHg3O
8epRV/Sna4ABla9pzvJaUCh0KOKNrBia0WRl+FYh09zdBCSc9e7HkH6Qg1ab1Uh+
TLzbvzt+zlDMPeL8+47151exNII6lX4h8gLJJFUJ2b26gZU9JqEJjT0EAWrZr+OD
aTgo6b/44BU5u+FVnbfb0I2CB8ibXr8uUBlnrcb787uWSdwj8YZrWkL5s0zAopMf
vr5sKDdgRG0JOUMnVP0CzmmhaJZcG87DCpf4R2WXLWXgHbeCehXCUnOpp3HF9H4l
b0EymlCSW7fNEw45SMUChSFfNmb9Y2WEcDE507zKo8xbNDF7ZfYfMPdsReIOTBkI
Vy1YsvWVVTYKWlC3C7GNbflmonv0JWqbs/zTRRbVGaYyWDs1WV7xImuCR/fDEtQF
5JVu2YH70AML3YK4K2tkMnb4RIdtGSYeShQ3qrEzKTGfjam90ML2o2dPe41845LY
iRTb1rOFb4EulaaJvtVweW3VpHDNJAjbUcPOLo3ixOTsPJHmgecVIxbESB7GKMBZ
bUt6Uk4Y5hEOFgMuHXTrbh6HJOcAQMMjsvv/zWSkvKs/xOQVzTsj2gc1QZPYmrJ7
TTDztBjJ1S4KVgZs4/wcgLzhrkUBT9h/rm43UAVbzp/WGe2AD6Pm9Gq37/2dQ8o4
YQm/dBAu/cxLJrb7vaiK/6z/K0qjYdmX52b4rF2qsejUmX8R7I3YYTBkbYX0Khkr
gadTppk8x6TzYOgKowFpf9MS4Uy31SUWNefaDZMUh1bwHiDOph5cWYHpb6XRp0i9
Y7ag3KlPofQUTb6gMdq8NDjePx+w/mO3X8tcFjsqUuKms0Msl+rpse9Q1Rn0+g2U
9QuZpudzcbrLbgsmUw4D38JFAzRZB+YCqbxLd0+h6WGINImv3yYjkqVoPL0ihcD8
soQI7G+58UxN51j9PGNdqPrTSEy1+DRjFzXQp4vWA3Xf73i+L3ZMBjMjguKp1zkM
MFwqDl39IHvxxERO63U9TKYx887+jaBPZuPRyG0M0vxYwfV2HqtrfIRlu+MOof6t
EK9dTQwLGC3csHVraBM9V8ne0AK86gklSRwBeh9/TqkJ1JbMaD+XX0vOcu6JYnpE
4o6BbFO7LERAoFz5H0DxClZoQsRbwZzIGt7gZbQr7TbXkT5fK+29IuN28jqGucnB
dZBtrRqdp7Xyf8KvFWYYiP7kOzyi8Ov1VsfDGwqXG7CujcpoUBHkTARujyAgS8bJ
z4HtxXpq5HvuPW3N/FdM2FLdbYp3g9LRpNL8MJNULZMT5KzngGvZELG7C433HDyD
VuNh3MbwT5QJYJslFe7rqBjTZtF6A9jmE1FvacrU2kPZbgbKoV31DlS0FgAC1//s
97rElJYGIT7Ef2kuMNBb4QgItWYihK4roQ3Cg/oIbnSYtG7rPDc8vueUJSpBnMrg
3WB43+aXrFul7Iws3E4DG5TXjkUw5wae7jSQNEseCCh+nw+3VkywvbKT1rMHJpLT
2DcM05hjFTV5bOIRhbSsOin8oQc9c1xjWyRiIEw64P2swxfU7zbO9g3QH9Eh7yuO
gjvj5oQykbbc1kZqTH0br3wCJWP2kSggkDBpgIO4H+UaU0iiFUivlEAV3xw7S5ZY
aSjN+v0tGfPrwIdU6UPqT0V9EqFK3CGiNdlh+y51PXhxJpJtEbEISAn6jnb0AXbg
xJxQCBsDRdQOiIiLM1jr51RmVA+vhIQ3FpVIbmmqk/KnwOHUoofabghwoCk1XjaP
efBvvMWQ4E9L7X1gTTtV5p2qGfzaHyF6oni3ZnJo8+KWeOphjYzn31oq07uEGX4z
+A6KK0GMLyRjJd1M4cqKjAqhUhBdjJSxPxZIjb+4ddht1B9g/eSMMb4xCrBJXNZz
U+86UFPF4c0h8tzzh/c5t1YW5o1IOQtHviww9EwWAleNJo8X3myQPSmdb8mSpQf3
NYD0KuSoVPLn46rFSw8nGsX9Y40FH0yyCYQxdI5Ccf1iT1I/lnpGwvhsLasypXD3
6M6zhG8nvtfFWkP/HFJTDJp7hqplAQxAC15C3mmtbfSnphoJILobGVuOLlmSsdrG
LK+sb187IDCZMVW3s7gqyi2ZKgYm4P2tPF2BcdPG3+CD+LHM7iqosWm+YJIryM9D
lyHJ6z/12lLkO3tKvoExQ8EkRKFAmOfP24QnEaF8eKku+DYKw/RNcMxzfS30FqqM
LlsjCWHiCsd6RSrYyd3lqA/d/b90hUDGlkCJQ7hTrYqJS7pebH7SCh/8p0cdVFCv
ItSLf1d8/eMKedHQmKR+nZEaWcIXg+xJ8eMFdHeiSpYxf8c+pywu6XiWW744O7em
5f7sSvjWp/ujJOwx+lVX1PU7yW4m23yMV595FfV3O7MDwF/V7g1jq/+QC2uFOdOw
FDOVFBSNAPsvHI6QpG8wYycPRPtoxuI2u0QLo7V/ppe0DUvIfMVzS41pvZXA1j77
tsSSwyR7GhBKJXTvqXjmKV3VXJrIDaCAEv21m8UiVZNwqgVzMtYS6Gb1u48jz/1q
sVU4d4yJzQ4T0AuSaDfitXJOZZdCtTx3dMrgahIcD5QHbq/cDtOs6p43l49m0U75
1LaTZSG95/6GuyNYc4JZ7OmjnUnlHHaGjOKpge0BFKIsUC8OJyTm/SKJs70aKLrv
T2zkUEYjkZPkPk42WE8CVlFsedpbPu67Oc/8Q1VOxuPZlgsfWOxIaHAFAvlW4RVJ
mCcrIWO1PJjGDXvDb0hivc2Mxv4rdSkG1xW5afN2AOJPYmOcbO3ep23rlIBSwV8C
snFWVtxWp1/rorUAlNraUOf48yYSY2ngjv0waZCLnDIiZOJn5EivU0k/E0quLjQi
RJQ3/AXVpFG6STgBLlfbaCFaTAtUbvB2aGBQykSWcshaGWL5Rp8O/Gfmp1FqmdLc
HpgQgpi1T4F5DafmxSKYCew5ycWWzsSPNGlSvyg7UAwSn+ynFFmFtMxH3dtv84hv
glRa3lOq4dv1QvKJbJBJ0SrmDLKM2CSSLHDBof8/B+Fk7H4jUjJjG+3NCMs/F4yE
7WnCClS4Yx32Emna2Fg7YSdbviJOj55dtkjOpSuHnNdpLNvBOnYSPWbdHZwKQDiu
fZZkFdOptC+bRGW13s5TPgPP8vr+b9sTb/fKb0ETmm55pJxtRquMkEXBt6W5kYNm
kLFrK6moa4JeXDSp6qtyb8C/HqiFKXjld3nYT95D2MbkRDFsmT8DhLooVjrLIWiD
Bm8PkpSZk7emq7c/AxpowizEpSbMt6PTBvei0pwMy6yEZjNYmaPIdGXwGv7o1wgz
ALrdhDFKXZsHM32UEbYQVceJi5O2vYoWmGMtFUqEareYeKvyQ4UISg8c/JASefd6
oDb7IBB6bmNP4zTc8hb0Dfb0LkwjyDS5lk0fCIBUYttoYdpP2ax/Rgw5xzVKFZeW
cFwoAzCYgTDC4mG5U866n7dWifSMe9qNLuGDH5XW3ks/QqwMmqzHGYVEfn0sEs38
vn8HqcZtm5dB8GD7He76s4W4jPk8TEufc1muP0gc8i/PWcfjhErcNOPTxpFrYQ0L
+OXQ2Urs+D4UHrMriyjMMlFLSPD6DNoqcz4MaLXsbYyGVxniyLK8Vx/gvs9LdCEa
kMjJNOeJPJ8QkeqfYQAyeyhaVY5v1bPz++aUO1yvDi/PZWQFoQwY9L2Ric34FJYN
ygeyypHVFVcloiuHJcYXv/fsylGpWiPrGBQO1qwuZzoloOE3kzizEG/ZKaHirqCt
B4LvgLEcfaqNitOs2T2lb8oHVsQ09P3xwWMrvP93h4BVNIS12lze4ofjIBaYZXSF
1O+ik5jOYT7qP5yI4CQpS2SjXXW6PeHStvZBiSQiMtDAck7oiaYyeya3cSxeo998
lphDY3UfqLmZwdcHektcXf6atKr3aNnUoUcE0bh+PJuz8sWyudiUzZi0IIgdfqIb
igra7LjOwh41tjgNQnl9jYPPn3g8L2JMLgiQ3OB0+kWNlcGGTGWxTNEQUE6ef9LS
FbfqizJ8REY0p+BlzIo0qefN6s+uBNXeN54SuEBW2FJsU9d1K5sk7KyNhJA03Fr3
NJuAPDYIwGdmeBIeYEEstlom7jgMNgRnIL4+XtANUchMy/v1XG0evixVLmhWOABS
X72vsu6GFrYyLzrJQJ1sIos+Cf9WxyiH5VTDvML7DXkABRxTbRgexXlSB9E5wyXn
xUfiEhLFKMk0Rsfh4/r39rtEBvap1mEtB48AGCDUY5Ubm7doro3ZZChz9H70cjtE
61UIJN1NEo4DQWrFvD9UUbAwNz/8R1+M/XdA2fyC+I58qsstwKjgHtIlfYtKB92y
uh/C0UP4s2zzlTfyElceBa6yH8IapX151DJPDtxBD3hp1IOLKs1ypJ2wmBTQNvc9
Lu1EpQkE07Estp7+VFTl2O3r+WxFGRawefHX5f5Vh3T+pxhS1BD+aJE0yBtcg/ap
aFxs9SWBqfh0IPd4y8CnmOY7OOqqdTDPws8oLUw8imzFEUBn+oPgElviWP/ptOjq
o3NfEX7yF0cDSxNOL80K2su2A49B3PHJqVNteRe6Gpuh6P5xcz8hd23PLJyV84dl
clsX/BV2/qPWUfrRm/o29Vyt3wrKkkJsfclK+ufMDVAnPYH9Xhn5ZM/fXeal24Ra
QC5BdKLYf1gnlr/YZoHEuJccY8gsrdDFCWkX5WUahjYVa1mFwGlpaWeiu/71sBck
igzeSgUdIfm8L4Q+bJWbFWJHyP0MdfRFKCNahUZKZcom6792U0sfEWKKGNTioG4h
mKXMmhTa14QR5fc8/7bjGqRO2tttnE83eloOMuUR+Ju8kUXdUfATJ0Eyszg1uAsy
XOoGHllnSYMPYRvBdBt72ka3D0NZxp2qBlYrKowhFbM11/gUo8GQWKVCIHdgkAUR
YTmgdvJJ1y5K5d5TT0UQHP6pKlTK2uY6GWfTy01qYp6026t3WSgJbSVqirsRi7vK
Lyxhmfn8u48PVJdVXFn3S3j4cAFzDuS5OXQhfk8/acFoluoV+SjBWOpEGBR67Q7j
VGjtIG4/evf2JKvy2CssrxUCCIlVVB/IEY2i6u2XJkFdVsJp+byBs/n2q38vYKzT
6O1LB8AFtQfDMJTM8r7aGyC4r/CxTGQJBVxWxs4VUcR8nwpT32eCCJAGqcZywh9f
8YobkCLzpOQoEliGU5xq1UcehEFH46PEk8Dqhwj9W3yrheIGkFLkTcU7gyovHJty
yr12HbxfmWAHRRWLYkZReWS8NohRsKeqDwtxx2vm8DHifhQtwvtMrFmOBk/ihXu6
y+Z9M5XerOGL4wJgCgoc9DU4X9eJMpiu6tQfBwvTAQIVh6MmoqeSpRu2r7+9gsfx
XihGyabPaKLLaG2/NH044g6F54P93cEv8iTFV4ZVsVi81N3XRbkd/yIoOp99wyco
FhEGQ5/GzgTsumMQYp4ICb+1E9tk0/OYYDyjCcXsC1nmC7Wap4dMMSTGkZmo/f/a
vJLY9B1/NHMhYqrN/l+yOqWXg8UHB1fj/IipQSHoO8kLXIFWVgHRvGjzCbzdKBHi
HhbyhKOs6MsDv5Yz1ONljd28GJwYXKsNfRzuck4Myi83tpjlE8z57VrEdjyDK9gM
4xuhv8tiqZaWkjdAQzcSnbyBL8TAt7DvT3T2jC2Lnicx/7AVCRevt+RDsPCCJf5y
slMubfM043RRUaB4VfCZQ+gr/B0zkhi6tSNQASOMB9bEg/IBWPIecaBAsrzm4PgG
Vko8X+RxOvWYCE4N0pwwv8UxE9Ic/6u9gmYebVEgd/4JIG+NJNToOFy2qP9nsHH7
Oh07Q5Pd7MuH7vc6Qtq+9nFE7coOi5oJYKKRL9xOw51YizTRiM4MG0dGBjznsdMj
MtTcPw9OTznfgQNX2dtHpE2eXGjg7MB3wYep8B6KxTKkSEhfMgPWHw7pxmBep+kx
3aYk1ncXz4ss+2KlVMS6u4CzuW4nR7j/FM7pnG7NGiJ5e+KuxgkMqZl8EUu0/rsR
f7ffcQJ90sOHxk7/EwWVnvI+F8AMyfQcwERhN0Ah++fytWo1uVuBhGsfoGCuigZ0
3kMg1m2lss83/0AuENxIF6IlToQn2D+OCc1+HkYrkduyLav+9CUCYCv344smGcb1
S73KHLqbI43ZwW1r0ANV/62Aauq7uYda6FiwPLPqtuOPDfNYzrzwQqcvs2nhXZQW
JNavMrWn7ttXR6fp1G4RDrsbezDFDsyUPz3GQ+6Jit93tsKJ7rxb760Mb3O8O0BY
VhT9toofHT5hlWCZI8Rs0G//vml9rTaHToZRy9PLyrg2OB4hfGVef/tAxckuSyd6
OMVGUaPH30lcfUJ9egGvHh+9TQvmXRG2JkIDNCDBrqnaP8wlH7IJq9TAcXDPaBxh
uAia9Sz+BmDaBEpW5JaWg07e4tsQXQ157zvfDKr5Tf/3JqnFcNla9yz1ejxG9Mf1
nlebCUOHR7tdOkFX+OSlx0sL1xy59XLBjv5+BMlmFzhkrBSv9Rq6XBdGNfzh7dRP
AB7uLS/5IXuNOL9fbaLi5QlONA3haXtOPxv3hNDZIGPLhiqhgOpZQ7uZa+cQQhOv
a+Xl64WFzQw7lNZ234W0azHZmU0FMqMDg6DnjFKbYG474Gx+vgC1Perzts+OjYvt
OltrGEBtp6hGEk9IkgIfO7IJWXgpT2MSGVfj/Vuhq2HEsmI67/YrkNfGErfz7/Dw
NGD+rpZWigZuU9ZJ4Q0qQ/0BDI8NV/8u7BQ/UXHqIe2OGrZX6HwkkdX9K0K4+p8j
dDMARMIoV8FT1LhUkaXhFLB1IEaqyE+Br2C+2IVh8dWXKeiC1qkWn5Q507vXZzgE
S4X5rlzeXIM2zwtfw2X2bueIY8vbg+Bl73zDGPQlb84LiD5FUiMm6wSPqtVROLi2
6RlLLrHVAW8ecuCcf3AIeCsQPDcspNkrzRO+muSJXvnaMXodDWc+XCKTBYZA+gdw
jUaabhXj4sc7/qJBaPha8xKagLfrrlqBWYB8jJ/W+eGRdVcIelQrpIHrvilVc6mn
+AiVTWUzFb8+LGNVEDScG7dK04oePAhv2cQ6Zd5aFOxa32eTzW91tl/TPa87O7pP
8oHW2EKyC64Iw741Ykq9EWzmfvp0l2WydwEt7DgyGYATtZav0kk3WQJRei3C1KMd
4JiXNjggLyHVVBF7BIkPOb68LF9/KiaQK7tG2LRsnUku9svNIrqv1HKjL2XzomBc
3Dt5medsmtm1BEWabq/xsiMjdNU/iQH3rjh5MtiNfLPvCiXnYggH7NJkjLLSs9gn
+gsAFWPSj9JiQmdwffNxzjwAHpBQoFMP1Rc34hZLf1p7oQ5StVg1BSWmIc0bq3+0
O2nP5U81redMGyuMKsZ/BMxvYA22QVtsgI6ZI2Stl0CLSPgZq4hpA0mZWp7z8ONS
N2TsllWBTgzBXWrvTyDPQu0BsJ+URlogXcwspsinP/H81DfeAaK1+411IGcBw6+/
hrx5nA0TVJwZlShpczeyiNhjBGDhgfgZeil03tWsCmB4m6uPZh5SAWpByYSvoqYL
2ssO7gevCtnLJoUyKz3nzMWdjAyBEuCsG4854P1BQmk0xXYM75IKOS6OuSU4wE2H
YWbsa/a2S51Y9jByYq//amYQ4mSt6iWF6mvf2envfLgWtYzUppGyoZYwgtXz36xR
w4nWHWyTFJvyedOB5AlY+gW+W+aRRRvD2L7XXDQKJ13jD471zBwiwiG/v+El98tt
sUfYIbv7AmqWvnZ6UkwDnuQQi7+sd5ueTKaFb7lcQ5YOgle/ZZdMFPb71pi1g1bm
DJGoLr1IUq0shtWzWLfFhCCnAAA3Jdy8QpcwbMJGCSJ8q+rTjqlsoadm4Ap5a6Hd
v9FOTu5QiGUWWwo62cmPyewtnInR5xRs3kz27NHDwlOxVFUkJIECdZhWsGPVpdUS
+xwK59byOWklhJWVlKfgpDA1P2ry0mOReASa4gSW6h1+H9Khpa8hbhtCln35FXJe
gkNr3UGj9lNdZVY07CRKk36l/63Csu3LPXK1DWo3STDQ56MS1IJLzNOp3zLvJvhR
p+Jowtjnkw3OKXrFWrxqJWijz+AdGSXIaJd+V4aV/XOJ+SnLAk8G4V2psXfdRsKX
z7r2xvQFDY9doxmMxyCBCGFngAdtZBGqleynw/VY4gVQWCBuuTDPmNWGnOabYdJz
QzeJb0itrSLVn3kNaHgSGa0X7y9jbQm6EcdEP7aVa+PcyCpgDYcAmiHJdEVBUQcT
J4P4YLO/JNa0iFCcUc5d49gkXKT/Lv4D+01mOcOdOcrkvbNYzpb2USnnqX4I1GGn
7DuZ2QtHGG5abLMGeTP0Zv6Qi5QtwQHwXLgqbIQCOxqOksr6jV7/FjJrEiqfsoq/
TUsX/i+EqjJSRgfAXXG2JF6viALBqsR1e8pKAywj3zNmUiaXdymx6iolqQaZF9nW
/TrLV8sH0eiFu8AWsaa9SOI72qiDtXbU+siNXTcZNNNCC7uNdBYhWsGuaygHTTVP
cPW609f+mGzhfx7EdCSm5Zhal0dRM70Cf8diI1MexvjyDvUi14BCBTaOZFCZzmw2
ayDh+eAiTFjQLUsEp2e6JIAOt+g/qcpUtxG+39SLLwqmuhdHQlwCtjFf4zgTnaGE
Sss76BPP1xJDkAHpAUrnuKwSkBYEfZwdKJajiE4Am/sakt95KLL27eoAwkxl+ESh
b8LH8ViB4+fQj0KcSz3N0LCibv2/jS7u9Y555amciIjXu0wzeEDyZlIjXjKnp4eK
oZnTLR9gv72DTGTyNw8n7oXclrd3aYY/KSgQ+nqVxuz1Kyzq4MZ1WMBQZtaJKNvI
ztO/dHTmAcrpl0ivI2/4EebrD3XOKHlRjFO1vBQ8Bs8oZLM+vP1hz/IxUBb66h7R
wnjwqmaBN4yTUxDeLbXo8RYXgx6vqlKAUCFMCYUvizNnAdN67MHHPQNetSk+aIDN
yMeh/1IuNH9BMti4ZCyZ1dzFrK/AAM5DEwuiGZCdCqDXvJ9NqGt7AVoUIzekqkyi
CFCfxQtanYDjafvtouHzlMd2Ej5AHK5kPy96oir+cQy/mOO0OqzdfwBJ6eMqLk1k
9P0zqRv4oe+sBfYqulG07LTNDBZyvrm3Jzq5n8WJN5nZcqxHImCU2wfYNwVWhys7
oV8vM2tPN5RaTMJ7IAp4ZbFMUaO0Z0iPPhgVvJWMTWIX5w3+M7lNoP10nsDLFF5c
ScNpdoxLuCJ/qLY6czbFuz7H6TKxKHESzSX6oKiREo2HKCqWJSnksqg3fR2TJQZC
bbRT7WkxvufvBqlYNnddZc+ZkHGyW3BBvaxVDmiST2wT+baGI3BUueTMuRBoLIMc
/Oxi2ddBhgbsCRgZSb9IueHKTHPyU61w5p1+iuQxo0l2730p/6G7SYoTnvGM8k97
sRCbbxWiMNxkszMublfe5CJS4OrnoFFN0F8swOYL6d8RXIKUl7ulY1BvWM61JFnM
IzVxyT0UC8GUUpAna8dw6D5tr0wHN11/pgb5Mfd1Y18H+EQiwlnnENal3JvICXZe
i/u+XWUmae+DQxGSDlXgYbTVVRIhxQggGz0yCAX+03nxdAxInwg5kOS6h6wK99gU
d8BAu4YAiB/odlWOk1SQahOE4Kbrf3ShoF/Z6pfFyY1SCAhRiZyb9p6uhez1psC+
4pIvFEi2VHedrQ7gOjIPB5CLpXfVdfR1d6gRBjaOScRjF2uHaqKPGUxTnQw1I6kY
ccWQ5nq2k1ckM38qJyUPJDaxqottWe2sS6jMWD9YZb8QlVIgQcB9SQ5EsaMzVJMv
4G8RO7kJi4uTts7A6PHpqT259AjMR2K12PwM1NaMOFeV14ODtRyppYxxa1HVvm+s
cmfRpuldsQE7M5eiAEq3y8UlKao+ufasCUMLmjxgQ+oO5iO9nkJu4QojAsouUNBP
nXpBjTZaOr+N+gWjwp5WFy0I9ZDS1ELWxe4Oh1urafblT/cEUxq8rNbc6Y7t5Mou
uIQa+gy68K8XT7Zgq3Ev5k4BJlaNzdlCanyT+LLp7N216nmVajBPbFGJu79P2Mu1
1qNKggzhyNC9rm2RvKUheLbZlmkevyWlk0ZhIy0Vlara+uEOrhacIqi+iuoIjyEH
fCRzb5+MvpFkCDdy8JUgfzKw6IToQOxDdTfAVabUcOCd0GuLojVZFP8vqidQifUd
bPbzdRWGwbhLK/VTeNJ8FMkd3hZj9KiYP10MxjYrdNJFWksMcSEWBS1pliY8EAJw
pY8F1Y8zCLVKlbUOObfTXiyFhOYVvBOY+mcxZPV+GGMDKaiDSV0iSDbR6LHE4yuc
P2suAdG5tyV1Ifl+2ibGlqSUyryDw57OMHTQcJp2Sfy5y+njXnKD7isea4NQBOE4
v1MyKLvvbOPvP2T01jYVOh3cYWXy+6vB0hxXRRDcJ9W8Ve8pfp/dbU8DK1eRPFgN
B9mvghhwXAh/hnKuK+N1qX1tGIfsZQ8C6ZptqxvFVq8gu972Vtw1FHYagYSnZyFO
eFlaSo21UtR5chKOZ/nodS5Sjcsnmd8CaR4B0v2znC8qJfPdW/3pmR6BFtn12q2D
4OLpSRKWwtXXrvnHaVXxH5omtWQxsM+FDHDJ9y+ixcPwl86DPhRFKuFRaY4UWTmh
jxMO/I+zZpekCVsUK1Ptx8Cko43kSH7/8sHP187oyB+2rWGtMOOSjgkWsMGDaQ9/
8OG9ysmmqmi5qn1gN4YEwnsUOxMBbqrmfHEN3K8tJqUdllhcctEe247PhAexL1Ra
rWcmra6b3XlJm5KJiooA3xQ+mfTfpvCi6OtWbTFbDjlRaHagbi3m021GZrR9uCM/
1KKVePFNWuw+hBT/zOu3+Yt2hGMUQ6iSIcT01Dd28JGlaiqEtUuBS82whCYNnAdO
3AEoyIl1zzT/eU9YPFHQJrafQozhbD8L7RsaFsNT4r2/aJNTkq5fdj8aNfEEC2/J
45fzCsVx1scYU4CgKYKh1sKfmlbzIYS+E8P43LscnTJshKO+eIDuNKR3bJMiZw1o
vVpatzorThqm5Dppt8GutSeQUNZHaDHH+ZVvAFPEkHYCHE4sMb3E64oZIaIFx8qB
+VDE8OdhjHcqTA4iK2VpDElhIFya90KAvmCOKtt71uHM263hewJmeAPAtzeWUyTh
ULVc8I11v8r/qmbgp9prMm6NrOh9ZV1xHoITA1ElqCWAgkvDDptQG2CspeRzS0uP
THC3qhfAsXQzQAo8sFyFGOdlbI3zBwlj8ielzZuq3EXovSILBOuT/cN6xXKm2MCj
/E5QuBAri30UY/FZJ9L3CnFe7ooIJ2/+y8S7SDDU9r7QMQcv6IHI0cQUUfiOHnn7
8Cs6Ukeh0O3WTv2nRPeDdUuBCn8y1TBuBk7tK18DOSrwbZ+nv7kwzLCPYSp4Ew/Q
5b5VSiqcAIbeGae4iGxoOXV3Nggn7cgfdVtUwuEJ2FM+wI0UTZS3RVhiYIPxM8IO
E5Bkntt5Js1Yr+jO+WOPmSUUJdbggQVwVudUGOhX5n4iRI4kRVdwhyHJWIR080h6
MvznlVTYZAytOt8An7LBo+llp8VRWfaEiUwB2ZQ9NkbcBm4P0+avxxplK1HJ6adD
30tJPwj3dsz+lZf+WvjZrGk/zKMVYpM/i6NkfGL1Sg2Lt7JHhzQArOfN+SRabFRc
GLUK2FEYyB+zWR055PQ7E8OM8d7LUvwxLCj6g1+EGgZ1PtKS90+FfF8ihm8bG8EM
6hXQ0D/8SzrkkZC455RlLOTB6OymcYskVWf9vOWwwnj3J6F94mjfUJeEMks2+eL5
bQ5mA0Q5GXooL/BIH5FeZAqKAhS8uOW2BJb1AAcjRLObF5Q6+udbMbfhjwjHcqsN
JzQhW0VwL1aALaN78FP4Uroc1neP9obMCFjTjS8y31QYfHvKmAlvToNeA0VlKSTs
7ErRgxq4b53EMCY07WYSziT6iUgswAyeYNh3InW8Z6EGA3FASa0wg1RgLo4n1j1Y
8EqZXqVkNq1HtCJ3OHUsG+qM0/Ve3viRQ6p2LNXwAY6RNA+qaUUEdpmqZC/ul1sD
SMBMIF6ZHS6OLBJij0UkohXRCYX7qbfJu6hrfYMvIwa5skkCQP15JgJDnvBfXU3f
j3JEj+Fu1GTtNyo6c1tf2Zje4MAib+pBuFnbAIo8NRjDwymmpwzNT9qexSmyHitF
vVH0hUlw1DiVDzbZkmpkE4ikuUJ0IfhbVazMdEEwNTEEjg+D6WowmPwMXT5MsJCs
y6JTdBccFcdfSRJ7ZcsGx26CHts6+3lEHyDB8I/BKg4ZorDR2hwXxT7dvlzlKILr
DZw7Wm5FUTQjpMl1ORb8fu+ZpDlEMw21ryK7CpszZVNZR4usyzmjQbX4TZC/Q55b
Ei2Ty3YVtWV0uGkA8GUWnybNRY232dS2riZLzCwe6Yi4HM3MmiWmJga7beyHFzG2
ofrGrac1Ty6ucU+w9CSv40RD13OaE8L+PHXM1a/fCjS22S+jNXho5uje4hCXisIr
bpOsgGWrdarEfjZdkz4+WB+I0X5Xf3mNpvahboWQqyTzTJRWbGeedn0H+qyRgqL6
58C5Iskk9EpHX0r5OAUBoZWh73D7DACeJIq1UFSJq20XeXx9+PWvxyZ3rhpP+Jpd
kFsS+P3ckJQcf4E0VVgl3WycyTYBcDvbXKVZ4f4Sm/eVL3fHIa2V4NHZKgyuhRSP
XdIxPjnZqr5pycC73wz7r/w/8qPAc0Q/5F4EnqoJ82p+U2M8lmxNR0IrYm4LDvM0
Cv9QOjMQDDTBPy4jfI2kA3tW+4vL0wdqr+dMJzlyjJfLCav6u8AuJtyzXzOXGUMU
i+EIYydPlGSba/0zP4EwpbVIj0M5TqWiz/ztGv1rGBiO9ixsok3ut3k7pWIFRL49
eCoroCkeabsjUHKWJOHeZbqCI+dQvuxgpvlZxi36aPOgMvdX750VmVxf1ALsibwJ
nsKmYy0xCli41hWGQv/gYONYbO7ubPMqge/pvckEzwDnpLlra9ckoDHntfz6a6cw
ak1X+rEpp7XONtxzKHYsqa3mIkuWBnKtEvwJVOVyBaNOiy95D+e9wPGV4N8eeQTh
LvePkKefCIRpjgN/fXvzG4Ekvfh+99vT0I8qFrdI4+JjdZQXIYjCq0kGtIqB3IcC
3vyZbJg9SgRt7xgT7sK1YdE277kNwki6zkLyIb0cYzIiGuQrPp0cHbH9JNUYH8hK
NQL984Tz1ydFG6G0auK46arazr6ceqVFLR9NKdLauWxRYZYSjcdo0exajaGOx8VS
ALcKu4lzNHp7RVWNBboNGR1Mca6aOGhpoGUQs5W7fKW0ipnX6qZ5LWx9zGaauqo8
URjVtRcnAGyDujzJI6riZ29f30BMazfNCBPx9gVDGWfhWDjC2gEplUYB4bz2eNmB
E6nC9Vn5Xart6sUUeLpQ5wYW8NIUJZDNJtREKtMOZOODv5J7CP7t9MVXsqIrvkcY
TJURzLsS2BoWbxExW2bNbMAehOkoab4YXattlWmdH3P+pjy2aSM/dIg7whVLLgdj
jefAFemwyH02CAFTMCMA94jX4Fv1II4Ce3NE5r3AxsPFIWOD2yGEOSib9Wp0KJze
15sMHuHmA7RnsMAIXxt2OQW7FkX4a7NQ70qQJay43E4WycPdjzMPUmhQ6XGdnpyP
JhNnVfMwusb9KIfiH6t2S8yr4fnWXoA3VEgzO3/jJl9diIQy296BwIuEwIYe21R+
ARihBERgDxknb2LoygY0lToimaLhFwx557RlQmg/ILyYwuBL2y+9jT6V0HN0g1UD
x8q/Chc8SRwVqCkNh3yefuUSN/g+Ocl4uFohk6EBKLBfcZrHZzmKbH7604+dYlFW
bHetCBZ1vU92gwIGwNSC9cr9bJxoAQwIN+n/1LSQEvLEKUzzUmuTyB9CsnVsYgsz
tiTtCfyupkgMsgE8dxkZoxmiXbW74MiffXnwUN8egoYpKP7Uy7sjEPwB67Eudakm
TcvC7QyZMZoMromJBpOvfJ7tj2BuHmOmIVEvo+GSarjb/PujGNDSGV5XJOOFMM4i
i7vz6DgtN8fMkSeK9rkZBjyClm23IQ/I2ZeR4FscwpdP0OPzieubzUN8Fzo9nwuc
W+wAtoDYdTMX94AozX9BPaP4mxTDuPyBIZGg70c+khnnY31m9mwub+V63oiDwuXx
dsdcWKK+wlv+YhwdYXHzs5Uf2odHR8eGEK9hlN6xllX3CJIPX60A/qpVaz1ZzcQN
Zyg0oprNEws1djEwlGPpGJyIIWYMz4iuxKXA9rFL+zXwYXkTmDz8rMs3oNaV/+cb
nA9yy6DZz09IZqKyqlwrD30+PCUgIhJjaz+h1DIiDHu7q1+a/9H20/npTKYtqwdE
CDG9VRo54fSgxvOY18Ipq9pEkBqXzuqjDHEMFIHnoCJ0P/P881vAuIni7qtbQaA4
Q0G6XEckMQq6AvrhpVSE8b3hnWjQ3XGA4gjLO7BxVnedq4GoOokZ62/mCB+rQSX4
nBUsTr+hfqHFnhoHBlG2m5n3eSG9e5OmPUH28kWrUlVcKf7WVqriTrfdxAhmKy9E
prOU+8nhgeugnLpEiZv2k8L/KygaiFRLE9FpSFmoAFJHF+ItcEqMxa2G8yO4czoV
w8pmyFM1uYL+mel9JDac8rCvmrrhQ2hUmxKtK9GPZfW034pb3Jyn0iDvCBTpFRIt
Hnvkrx2ly4/Z7M5ZlaIT2AI8jycVQadRyYiXRjAVQjy7sRX2qDIMvOcm/m1l/B9L
Egd0u0DR1l4GZOCUUQmE/L7szDA3B6YLkjwu14Hr0JGq+wBdmbMIL7Tl8s3qoCVH
mMRAlU8FCtXcMo+24eHIctH2bw/QdWuBGy+IyUt5zZxZM/kF6lZIQL2GU2KYBOSX
G84qwFDqjyRoAVN8mXeqmK5JABFGmugpkTssjdUU6wbvMzNs677SgxEG2xbIKHGw
vN2JlZBQtbmFNhutj3i+d3Iorj+IIRYzrUxqS3rqStm2v1Pwt6SVs6+NbnZ1hM6+
VzfZjeONODrFhaDAnK+u/80tOBUE4d8u84B3xZefbLo6D8uKTe6LlEcn3Q5HjLd9
FUId+Y0G/3kkyG3qYo/9XZm56YJ9ScMYTJ2QZfkLczzaaRNxuQVsrSRNTc3GCBzk
SjvBpzqYAFPSB0cvgCCj6T6K9MbH4vY5ENXXIdyMrU/ZIbKe0V91oNGLfYhZjpT2
qJJ5aSJHz8AL8HONu8/KMXtEo0n2/Bp01gn+CWUpxODj+iBUaAowQwTX77MIbifL
ISc3QzpQGMBx5rl+CRYyxEnbJRs129M+oNgDn7Ft/oIbm9rlqrZc7c32dRxDE8zE
OKDrMY8LbQcwAzPv6rt0qcjVE7m6IDz6xnHVwOX5S3U4YjeK7PJ3VjTsB3w70YAZ
/+ocIwhSWxd4uSp20k+vLg1QpS26DSqr67oqiwvuvMwBWgdYqRd7cfxBBxs4FYUR
Oe0ku6Ii5+TFTmndOx2vVJOlzm9u9G1OUvVBk2kJC/7uUltUIMELZ6FvE3qZn7Is
lCB1kq3PZwv0qby5wwpIyPoyU7qZzvydCBtULeGEvoSreGaUigM1lu6BrI7/3Vix
j/XMR9v/lBqX1PCpp1rxwzJD9I/i2yyH5Q3fqqHTGCdi1Fh31+ycRYzqqCrehkNB
PO8QMPq2jD4k08bBuV/q9mzfOIvqYQniMOoVx5Z0Ea4r9240+/9UQxsITj7yTBfX
pmGzf9KYE1ickne2cD/NjoAZyVAFEZNHgfDzfYJ2VrLIjizy25mskmkuhwcAt/VJ
IRaRNNpi1q4MJc/25Xn14hMMaPn80P1NcdIbooczALQofXmFhlhotnPGKFSyYMno
Zg+woNmeUdXgMSVzC1AYFrAVb63R3hkbIs6a5SXksRwHaIABGJc0xEABLT0JopX0
0HZBOVi7uUEDXiS2osr83UMLMLWZZg1KFssWuSAnJ7wwd8D728EE4IutkpQAlB5O
QqepouoxpDR7NhADblBYkmXPqhEuaFTvgLm9OfSJVJg08m7gYVDxfq5MUXJlD0/9
GLi2A0H0F1/nDSju0AlwRuT+0JgwphByaPUA5o0f+KSeAWXxlbNgOQZU6JJifIFW
X807tPJw+ap4tEuU7rtM6eeklfc8IdnipA07mlUJTcOxUNQxCxI/KbHrD1WG/KQi
URuZapiLX5+s7hAUKvxT4TSnsGepjVL7KPthmI4sdK09/jHmMLk++KGgTQFLVwNr
Qm9c7JZxafjd19oXQBU2GMsbGJ9LWaYB8FvUc9GP97LhI0XW0OmOn0OgMM5vSe+7
0ckqPMjMpKFKhlK4OX471t+EiGWbAUYGC6nItyqYclN9kYbHcA2C1/SFGgsHcjpG
Sbr2KGniPJrH4Ma4XKZQZGrRNx7BReMccG5RYsDKNshC976hkOhH8iCWfzEKVhmT
fitaPYQXZCOZTtpWnvgfbBI+g9GGpjCk1yyhpS7o20ARNwF23ux0lRjL5zC0S/+v
zGVLVH8C+PdMIkQeCT9Xl7uUn3+3V4zdgwSRo+4nMADHu6UUPVFSnEOMOxTWiKwA
Q0McFY4aJyZ3pJLXoF3dV7MrPy8whQYoXV36MrEGu35Fi0j9K+b8O+2prII3Orkn
au3VRNPYxeq0jnnWqCXjIkgOFpu3Jn3+pgJupljWKCmrPBHdxg7YvIvOIAQXpa5h
4TnJ23uPrF1LbK874YSNAd+4pKQN1ofMtdfwTpYmP99xvJqbDqi8SBxzdu4JKJdK
C3hN/cQCJQLK8LiR2tbPKF9xQOTfNrQukLMHNYzSO+D3TBKrzdJcvZlO0ezRGmHL
OAoT9ONi3Lxxp+WY95C6dC8NcAaBG0Nby5AC7zF9MpxZMtVb37R7h2JHFluP+TyO
/ZiF/MH3fyUk4ZXatvFkCfsbc/J0RGQUKKXvNsZ53fe2t5NtWSa7oxqCBotA+ZZX
74EL2K7iv51dd6cmDrvAb1jXJUPFOTlkL1sdBAoZ09cR4JKQ5Z0/voYt4nkR8uDD
VZFW8PjQUnqHxGeCZfOskSCRug0k4SR4KGT4WyeTsJ2Qsenj1wVId8sCypzYMbaX
tIiyEsMex5eU3T/2rcrxOBIl53xwcP7E3fFWyU+vwJzARzk6hTLhYzgA6O4Y73u5
TzGBIVjP1Uyrp08G2S4TsmTfsYrncZ5KbfMtHJeJb3RdwS6AfdcA136lqL9EtFtw
Uyza6qBDLuS/O8ZeFd247abe17PsSas3glKa3iBqWj0IOgQQ1HcVJyjMErtnPCXw
l16sxlP82lfBMC8ukE9H1t+wmlVlH265ZesQmh63BLyYK1ZkBT3REgbESuyxnp/N
uZDf96lJqxicK8ClXScrw74g9dimKXFCMs3ZS2V35u3RIjDKaSG1iclXBibsGdlU
0s2C9Ny9gW2F7uw2iKvT/Imn0/I01LNmwr2xvRpVXLag4ZMZCL5B5sJQiEdqQJjI
w5JB1ynIhw8DpNInFv2uVDv/WGcpf6hICNn3uSKhyehGthuxpgHnLm+GkViENMd3
uZuSO6HWZu7qdGgmXRvngqOeOBhBCBR6d97vw8UexV9O0gJqDkFeTOCLGmE5HaG8
s3CLA7UjVr9yvwKwcnTSpSa4GPgf6G7rLqraGBCiI0hB66UumSKJSCNbSCDEtwdw
fG0NCSph/hdI5NXuIi6Teyc0IVm91P/PVyhNz+UStWA8LCfZfz278hqZ8buf0kVI
P48oemDjWLRvgA3n4JzpvZMZm4x9iAer+bocqUkdesZe/OHWr6y88FsAxEvmLBjq
s2petnWiinyeyvac610ApNoCDUiRvWYv0sC0khwJp6Lg3wUHIcNR+skh07uKRHfi
WiLHCoAjerO4cCxJFOGy9XDgGQNoXFhRZ1MdZjBEI1nX1s5qDxVhNfEPyHzi7EWk
vmn53a6nrGXGO285iPLjnar7UW1hLIOb0rBWIQz7lGWpzm5IHkLR6YjkT1iewlDi
Uwqn2zVeNkaudPAGEcpGhGWwCHtKuBDiQw0C8nSAI7IuXQTfujwrTIZxIzAk9Ame
1mYbI3Q5grWN6g8gK6GHX4oVL4WgnZVGmltVQtORrNsvcoLWsKncQHMYzNOyy1D6
jZpufYFlXoRNBzMfSSL7haQYfZ4Wh3Wkfhz/c0ujUv5zkmY4pr21UpjQnkbdhNNl
VhR6RxYMDZ3iY3kwAuPNXLalXXGEVnJhknAhacV3uZS+xE/PpD1zZFZvlhGLPg8V
HpNxzves7Qxy7yYc6V+kxyWJVxeRwx2iBt3vlb86DveJSMPExsony/7NKR7aEwAN
FiowSgP0YviugCLfnmCMm9RUq8//XXDd5JGwysTem6zeCn8C0SpjowvCECv5sfxg
lTZ63ogwdrzbYK+nKPr6tBfZAeS5kj1EHmBfygYRIk/ty3Ze+HBlnBBw+J0wnkKu
h2N8hqu1bXIKkDKH+i5RbM9HYXGFEjWtezzjK0STg7+Ol1wVJd4wOR9EMd8c/ZCz
9A6yX60OviALn/MGT9sGFRKHROHvIlwxIzFQFg9h2zEy6oZqMUdFPVul7XDmDz9b
eQJODKlGXNlW/O9a089P2Z17H82CA5fukU+YgcnlWfj8Kvlp+ADOC5AQTYouvVVV
N9RviShq5zpKwK+rjjsoECEVJ4vrXlg6jGHqeycBB5BfmA6epMVeFghg4slKCi5h
AnRDEEHDubvkhFPRqsmnwpTPl35d4W2u+dk0nrmH3QiCe3rt2B509lGk2q1B27m6
79zWuFVZOxtBosseLZA2AohIMsGyEX20cY4s9ciYGw8ZDephekKm1/2CHjxcJ3Db
Jpoo52tH5Q/VCcFVSB/4zCW+RbJS5eHfcAmYvPSbc/pnS53mmGNazAF5bRpVZ3SQ
DQ/rk9kPsNWMk87eRc0jX4fuSAbgIxQ5tChbrGbGgceStp3BlnielZG/jc4F6a2l
H16swh4V9DhYXhmkai2HU2dIOMaRui41vurP8DI7cAUiJV6MgEq5TEN5E1accvfN
izGT9xISkJwW13oun1Wk/3uPXoOzAjlKnJ5F7Rb6A+s4l7CATGcI1hpyBVKkf7HA
tleTm5icVNDs5cWGGRqbn8W2nn5zjXNketAZ+1yhl/aaQa2erVP+J2ryL6oLstAp
vBa2VyA2eeYBeT5vlmG+6bqOto01IYxz6jhhUhYjs8vpsKZseAgzkU2pzoz6VkWJ
E9yjAZxYLC90FKWR/n1tX1Y3NyPzQ2SCXE1e7CEJfLZ0OSfU4DjmzF5nTVKd8mQs
FwX/QosT8DBpNrsOX2USUl0CxBsoirVG6evYKm68gJEgEPTxBrJyWqYsWTFOkarX
lRqcm65WDK9rBX3tvwHwCpfZMaO/0eETgIUHyunCGXB5+/ZaiYM4m+YEDbwgj/vq
ON8SMxs42KWiilFNiGRYlVrij/83Nlk8rl/20IrW70b+KhUwCRzr0lEpuPMiVGqC
6gzB4+edeNbGDXvtLGFrt3vaoJOeqYNhff83/9bY3+jWzRAb7NtMkBIMmPhZgXM2
5pdxySWTznVr1zhDXfB1x3HyidrVB064spndR2Ab1pjib0USDaBONvGd/LWqjvTO
fcvf5OTfIEGqhETsv3mF2VYiV/4XHAU/lNGy1Da0hdvahy2eYoRA8EBhO0C1ykl9
lDv+lPXgn8tvcnM0bE8uAh5DrapbbFRQLLg8SLX6yUiAIF0UonmHRJT2wjOs9S61
eJ89ScjZPI2cEY83RwSr/g2s75OdoAbVCPmRmMAdabJIJiXOJ2vTGJVzCNDgkQHI
O4w975LyAlYa0eMZON4osYnxv9W5m0DQoqsi6N6nPrEMccmHJTC+qdqqeBNgi8YL
3Q4nRKvKbdE/njRdn05a5MuWqgmYO9F9mO1mRv/SuJoErAoQtn2DN+jl1wfYvP4n
lZUFHdW7PJukf0I1qCh0660LCKyMPyvpjBLKryDh+t9XAenWMNA47G8jNViznre3
G62n/jjF+ne2/suKwoZfD71ItItc846y5M6wlx17oBWwQe94K0NtTcuc+Nt+szyb
hNDr0Z85nuKd3FOQkuwn17uDXwP1Ock+ZWQFNRy4cWHjw+hrosuFgNdmYSDZ3Yyd
RwXM4YW1wfqYZAz7fBbqPmYBnCe8IN6amieluk1ARfuA80ROIEGs2aRPNZjHhMYi
zqHp3q6lx3BCFRzLW5dFw/qNAiTvIHQRJ65KLQyn8WTC/jsfkb+GG/v+C4UHxUCb
XOXa4ZVwacoQ4vaDSFWeP+SWA5dTqx+3VgRWDsAp48csH7mVQVofpOxyr5ME/p0b
PkEnEsccQ5wTYG/HLyLipQ3PIUc56DB0gRSb5R5JQU7x9a07MlYZIJFtD3fWuyQO
i1RDeyoVk6xU+rLbGZwPXHvzueNEyQSCd7xQ/Jh7Kq2+R9DelRQmOZ2FQ6hkqR6Q
WZfRsXtX0qR5fzTZusbEjxxJDyDyr2LyBDnEC9WZH1hKop+E8HWY52L2SQ3C8Z0I
JcZM+YqpqTzVwtYb1DAbgrTn+mIiKzaPMZn55wiDtIuDvrA0wcW6/IfH5rQjgVt4
/o05zkM8e+As9Jk4ZwDDB/jSfLzoiNOKgkXWFRKAGDllfinzTXuB8fKbJTjA7zAs
s2VtvOkEo1VxlAvoSI7LjZo1hXzyEJKLAIIFuRldQg9oG2IYSc3fR28uhAw8QwEr
FRNRLVtUlkMWOOqrCte7BFGSEONjOVBQnwCsYpVh7Zhx/ew3b4lMHo5MHFFqefBG
TfQTRl3GwwpJmnlyeOahrHNsh8n5j8TdxijBSzbSDk5BBLE/E5CjXnYkHLIs1RqF
8sPFfrHkKC5USeYlquVgnVpynJIG+jrij/Ubcs21FD1DSkwTDy9p5eRy4d/dlCsK
H9oX5S7MtEoYMUqkTltaQW7PJnh2047C/mUwi8ix2GrAmI/O3JRGT6GT+nQMNR+t
8e+DulmaWjHOcbyVCYXfkazIssuZ2qf3BDEx4L4hiPS8pkwWLeOOpEhMqGjbEwDB
/aK9ffdVjgEZc98cybc7rBvaDbIe2KKrKcSRkM88gGI1Qz6MsEgZkG2RTIVz+0kf
GaE0NwHtkzPobzWQiQXhRiG1Q0huSBvrkfASVJe4UX9dfAB3vo+I4+uPMq3PZHCf
goM0N80gmVaACu1vURBQxgAlj/WCcyJWZ40RP8ix8FX6lOHCoRj8TayuOL/hnPx1
Ria7gS5NyaJ9G9s8IbTYTeM5yyVRXwrSIpRjJ7brFf4iCl8Pcs6EsodDoFRfO85U
baRPkW3z5a1e4Kfjossx/6McC8fwNPMIjBtZ60pZrBn9fOnqT83upjg65ZApba+3
/VugmG8qM0ngY1CRcjiP8Dfa2QCJrkPLmm59or9xRZC8g9YQrDNIWV3L/5ymrxeV
l+unXwhrqy9cjy3i+YGySB9VMYulLoMSY5CmLCgf5jwWyc6c7BFl45DmRy+4l21x
rvwptjgeAHjJXfEqzzQUXVkaTo7ArLfs3r/MrKfEUq0JQwoBLzX1RfPDjXOt+41F
5t/KOfPw0mX2J6svUpxEjwXI0/h0KX5rz2K9GAcGzgoL3JDXymAK+xs/ZXpDV/85
SpajYh9JGPe188rzfLVGilIQJpcirBnMFhZknkmeuhg9yY/UL4/lLdeOpOCpKymH
zluxc1fTrHilXiJ9nDylmf1ejS4NCgei/Q4BadYGKMqzmVXFaG7+t7Fee+JaWl0h
vTON//vWcfSwRx+D85BkbyeLD5lMfRPbFfUygKOnSvTIV06SzrvYUVTGB/Jg6Fvg
Z0/0kcGKRWJ3byVDuuQoWyWW+UHZ8h/lyGQuYWmZUmeNcJssiydLS7V787UYKi2R
9fajWqqcWW296qbaJVhsmVecdYSogIqQkraPzE5MlBR3wDJKE+xpqX9T5Xljwf6s
aTZ5hp0mFZVUVBxvqVHUm0ES28ASR1x1OP3TgVql3jzERMl30GjxGz1vT/3HpyeA
PQs2Iny10628rwP7vdssGW61D+zSG6SDYNZVJRIL9g789pkqHHcaVdn0OIr6M+zO
B2kCXY+jZjZrq8ju6LbkEciuUriHHrYnPX1OrskfDBZcpXtSSFc7gK8YfS7lg3n4
FBb3z3GFE2U8Nc0aUzaJ/tNPvw8J8ueWurVs55jMqgTZ6jEpR7HtcrcUBxxt1Nqf
CaDBz2ZCROyzggWiI9qX1jfmnFsBm2TrEFReAsYH1Wr1gq/5h01q580ot1gnUcsn
bXWdreFaxP8wD6Axo6IUQxZIqNAJpwHl8vvBXJJS0zFSGZVU+J/Zz+0hFU+l0jy5
AxvbyD0YwPOxRZymbhSusRWm0nZ3nlYQhLfFmPnTadl4rcIC3QHI10vufIgA53HH
x/EaMABX9eZ8xZXGToNml9I8nWpuf39F0H1mebTC8Pf4cVIEFqq1wOaeOlg3KJvd
dRGbFY+YkqMbL12aFvVoOzeKrf0+OnfKB4E+cP/W+jWmrBQ6BG+qcutwyyJTCs/l
1o5qgebO0/WdSR4MZlX+JcxfiQBsE8LwJu5X7CpJjePsWkbraNxIXKieqa8hfPVP
Cio+czMujRSqxjFfVIfMWmhVF9lcXgoJqqz/VyYHpr4kdYrmy1jPZnXZtDiQjQDA
ms9QpIeQL8DmcMfP8ngshEd3kPPAEvApThUlL/as3SdiwhyyL7fj2YvHhfWWZkvv
5KAEhmBQ1BF90uluDIHFNUkAkb0fBlB0TwCkRV/NBw7cs+9Nueh46Gp6nIgn9Qk1
L+kKwtKA+i49tgJbd6e/p8fgPbIFUMfNaO9skV2qh3Z9I+nT0jodwiSGVUOG4cCA
PB/yLFP9OYGp10Mwjifb4n+Yc+c3GIz7lnMmP01APuArTda9VqsCx1s0NPwYj6Xq
36FIEWa7WZuilkqN7vlr0tEuIhNRpf0PvhsAP9TJvTJSrNNwB2i7OngG+bmaM6Wm
mENaKoTwbwenib3S0QYklPZY/IZ+dd+lTYVii2ps0PikyBppbLjgjfWhZR7PA51I
PHoqSa/42NB4iooLCKKZXZRTd5jvKmFSTjjGe7efHhZXsTAy7La1f5vr9V5r6xUf
e6oLXBSrQgYnW+YZ4b4y2scZopUYoMDZKYG+/hDSL8FIimVfhK6+PqICz/IdYzq7
3WocwpZopzViOO88bcOQjN19mSvuz30owAAu2O85c2kiSS/iSkQdEVd1ZnVP2i3z
TjiY33ibRGelm4v/BZ5RCgt8JsBSf0Gd9q+JAPF+1Q4uNniPclCKwG8oXIVWRgW0
110lm+FTU/ZEj5RpKf4TfpZLfvPsrBE7tL1KjTKQ+uhdovdqzNITlQ8ozCFop6q4
r7MYQV/agXfC/F0xEWN9BmX4QmzSdEOqU5fQ5ePnRHQHtlkNEBgsA1fx8tffzZDz
yQ3oHlS4I1QMReeTMRECYna+qw+kIJfji733TTyA89sUTpcamf6h9TgepjQVqRqF
jDDK1A6tMFVlYD+l5bLJ0LLKZqBSmDMsBPhCObVphURy+yJSMWPkOKpQYswfYHlE
+I7LQbk9IlBp7DdR3XcCCnceNXWBalAXcWYB2/tuA7Jrv9YUu8x+jGEPpdMc3lEm
vCv67G37FtRJuOzwy7qRxPzHGeHYsyJHlzPg5SSwJ65G/5duLlDUJBHP6UIAf3EI
RdilegA4H/opNGqUJnDjbGh5ie/uXfeSLut5EqVreCFTTDUqFXbQDHqZbIfu1I5j
4kHGspiWsgPl+e9mL64rNgxpQYcAReQUSEeG8pTclhwo0AdPzTfSCX2Md+p+qJic
WjhzyiopYmlbner5z5PpjkripM2tCZ5FmFuR2TY5qibmlgPZc7ZQ6+yxO7B/o9t2
ey+LYqKoGnOeaQhLbtPcXuPsQsbwfdzJ28zlW1wrGpreYaCB1/9ciGjqAi3kE+W7
pxiggXnwYjSqFv43Lbs6dDabScnU4Oukg0RCHR3RpCo0fFlMQsy2aQBWsN0Qe6z7
gKZdemoQLUHiMBsvamminfWQYSrbh9fjW87jDfpYj6xrbUCu7fpu5UydRBFB06o0
vFUJ02GGaPWwjC7ajNnarOOxn/sAORhvWWybnYg/ecDPIR6912qvWv3gxE0jgjEr
2XFUB22WWe58RtHsA2Mns2l2nROl0QWPTzcb6Npehv88lFSoc8l0h2ueWrQ9kkqB
2DU7VQSolGlpNAf+f8CM9dnuMESEecTPNH848aidcoPcoOICVspvqFY4QeVRMkXU
YiJBrnE1jthGQE7Zt+NiYqq/W0YxBwd6IwOgZ/IfpZ1qOXUlnGCKGlpvzvqYSU56
frs4gTyMAoJDnEpJgvSrcNWvng+oLH0Lk7rrXhIF79JXJfRJd6Wx2LyCe/Te8wWM
FJWUwwkwDxfIqoyKtqyc6f/3orAzNNgtb4wPUefCimbHMbbFjgsZ3MoQP7yzkjBQ
CSZ4ijojyuBIZWoVuZbo1SQVVxcJ9+y96QfuUoa2SQJ12th4ZUC5aKd7EDz1hH8o
4tdfo3ydLpM0lGN30llVe+34/wJkgf2BWaKJG7djw/H9v1xX8NoSue1BaQc1/Egc
4m5AP4MqIevEW65gLd/zRsnPf/SpPtFnusZ3dVc+JfBqwXDVTsMo1i1o46XbbEqb
yFe4UwHaGS0L0RkxsTA0i2htAn5pT0Iz2YWQvix/2/t6HCDvbUKlbDlBbe0RL58B
nk+CZvtH5YVffFE/xUvTExE9SLqAWxEtPzjGiN3qWQwh+I6/Fel4rX9WLoXOHnxF
Wf8XmaAAKUddXcwaxk3Tt0P4wugyLbv5wla1OUHALwsDFr2pr6M9MT72ZlQIxkan
yU6mvp28dWQgyLfkSBVJ3s7kv3td34pQMklep/+tHcr0pCOBTu05mEBseaEggia2
80ZEX48U4GLalMnxm7xCryE6+UM4kGGZpPxD91BTdklfF+3M525KH3AaGZxUjixi
PQTPDl69dMJGt2RFlDYbR9ZjyZoYMz43S5ecPO3SCy/I2www5lnjUBYhlaStZvu8
qft9GmSgBxwVI0wi2Wyakf/aTziD0f3Ocgw2VG/2Aqd1gfu/z1XeIismOIzwnA48
qd/3+iOVBzd8BZoEAlnZhE+yyKfu1HUrv9LnZHH3dMGzGJYGAIX4zZDfimihuUh6
Jom8kSATdkcBSVS/YbRGOZzvNVIsnuODZdxX/w9Bf2Gs7ZCxWrYMRfh6a0eOOiTk
hITf0/EP9ud5JRK74kHBuAMDiUtBnsfvjvD4JHsh5mLsMVqhqvVCNBV0moZOplEI
okWsyGc3IPf74wHRIqjy5kth7au0O6mxmKE0DD+DUaBZT1jU+QNszqd1qLYn1472
D/T0x/80m2rxAtZFJOQTAoTrJs1T1VhJyD7qEd8rwbYRHeNdNcliAUO7RtJgtEuo
MdY3eIwUjwNbhmeFWJfAaW8Xjh6egcj4Cm8dQMqNY38YBvz4qNavQzjKXR1H7OJZ
ewrTe2i2g1rLR14gBKq29FMRW4IH//XrFvzOrsxBHUGWVH4MrI1BcogEVbtvpg/2
i4+mgD2ytxa0+E3sOmBSSYbL52bnVYCA/Dysdb67NR7FJhRPeNZAVYguuKlvv24c
s6qSUFn90pGiXC5fJL6FlD+q4mrL+je4yygb0kkATIfI88rl8w2DdXWO7gyZB/Ms
DVN7m2Xq+HeLgQEY8AQxoGBnWfJ1Tg2FmYAj8rLcFPapOjH/ZZGBoGrq/wbyqAr6
5nnH9iWzbujJtuho8bOK2JD+b4+RwVT1WqSFG9vXxJHPWolXLcldhyLSrim+mjfX
yVl58cTCuIOaSjl4oqNV0WpXonujg6mp4cUr+UOX8iKrlK41+C324zHXn9h1uFXh
1XOkkldBXm9dOnhutILS2pIvsA308LpUmFGqvSBhjgJmcKJwfqX0ArZTT4VlNnIf
gxsUjo+HJ2KPYe4rCKUd1uxHiUoIeFe1nTbPikDXECYLp61hwKXPn2o9KeToWLUp
VTgAnCtyHk7qAls3h3o8HxsiXWZaKDb0MUr1FbNCnjlAunVOfPsPgzaQ7N6cyTVj
FSt01SW9hD/e2VVrNXoW5+dJLVhfvAdelYLch//OXcuht5k+aDzlxp8ieCQBaPWK
6Ckc6oJL8B9qKZWzdMVD2Df5PVuwm1aWBV+1Orn4dJj6VZcxuZLJfQm7g4rQp+Vy
vH4YYanOnQG0DX/cnRJLRygye3Y7YzF82f1dDhzmjtTIgzKqoKSj0Jjc954iq7hu
VUo9/cn5hSW6ovvQRZC9lUlNgwGVe0x8rNH/JRiXVwx1lKZgZXxqwdCD7bj0wM1F
NXZD0JY81k6cvYhRRxL6wNkybnUu/mw5RT6RAZ1VjL0HNchMqKC/DuXzAaNJljSU
Ng8It67k0pFSVc/tX63Sch6E0Expws5/79lPQRakRp2w0ibqHnQuzBrX8Ounr5v3
OX04srrpWO5/4TkrSFoHX1RRa749dWIp3qfQHlKOZ8TutDhj7X2Mmb/0Gikqxdoy
GA19KYkRBjxkLfD2KtWOZJgxsVjTq3LhBuaKVWSuTEDUirLojmr1rKVktZujQw2Y
gjOv4Pkaarh9dFNidQVslwjJV0QCy/knh0YWtAO5Zr6jvE7vLKzncPPUya3VF9ML
aiUlaUdtm/wkKIkzabugCoUQEBSgWyLSOCGK1MiUTuHXmchcoXTZ2XGm5K+WQrPP
5lhrRrcY4XX+x+8iQwXbQL/z1wbrkmJmqRY9v0LLXUW17anUe/7ot4WMXfqo3z1K
VhsyRbrQnrbCY7WCCZZGwhk/mY+Y45w5gnOO+eAdYXBlj96BGIJ6w8ZRFFw1CdTz
cINPI/cCJQ29KaSrtAJLIhLkTEQj7MZDah3aWvPRFUwNIPe5yvBZm3tBC94mfaQy
6LNneQI2xkyX/l/3Qc7ZrbuK3ohX4j8Z7Z7dXEz4TXOuiPJQhkg/zcGOhk8grGAd
AYfdUnj+f/8L5UBmqkAKLo85mw+fuW3AB98Jgir/Qbwj9bAOMCvLE/5NdwLF5ZUn
BEmeGzL4hmb9GKqgWSl9Z39nvhJyhK4YMDKopDDSepikZ5DvLE3u7c1JR/AHhqcU
Pq1MsRPbYCq2vF7qBgvvks5mbFlo3M2P7SnrYIKAR4+Jf68GEUhWRvhPQCt93QEM
wV9CTDIAu20datAO3qaL+wrd9C+ZPYiYhOSlBeI6hjofS4PPBACn1CmhccYqAQHE
phc3Qz1/UNuz2eeHikqEck36KbzvFN2KbO3WaAzgcSmwAYIqjvojrfJFOBdCEcJA
M1UWVB9J74JIvfaV2YYmaTLQ9Shp6TBELBcDSYX/UH5nEUZAcxp9Cvw3GqIv9OSw
y9qzmhmW3Uv+0SkaUFpAxMaaNM9VZgtuVQzbqyN+tTcnlxtZ4JOjWPFowBmRiOf9
sikn9NFucW68IR1HA7yfdP9+UOeC2VPCJLp6vZjqjBBPKubuBBVTd+S7k5yk/jU9
Hi09V6KpCl4m7LheIKSjBBXUKdrePcYEVBsrIl7CteGJ7D1PRQFQsiUpvsZr/6uO
gMDTyj2qbLORN+/xo7WN+Ir+bUcuUUe5JINCMZ/tSB44OtLBju72dta09NIa38XO
Vpn9XZ7li8yoUIo3UEAGKCct85uPBUpRMGyfI+crv6RpM2wRjCuOV0oSFyTGSfQi
N0e3jALGUGy+NFBkS0AnkzRCSF/g86gh+Tv4Ho03vuWD7mo3WjgIr84S9KDIO19D
6HthjJG7y7ak9h47rJ1PVxvz8Q3w1lYpyt7K2ykPi3cpuJtTI9kvMGS8AKKwh+cm
C3ovVCeS5Q1CHz5hsaO21XSpqJMnI3VnKKAYY73kArh3dQEJ1uWDwvQMtNrO3vHN
y+9xnFdCh+umc+qUBymZeD0c08Igp3sNDbtUA8uYhLE6EE6nmhwODjJe7WRtbb+/
cXt/760cl0avPyQk9kJqCNOPOZ81crh5pfxtD4mgXrqBWATOtZAPz8t7yOSNaNG0
xGpYWtO10SIgNIVay1jxkVOrG0isiZD1fr3Ux0Z1OXCGmTshBk3swpDixfBDgZQF
vLJiPIeZk8WB4Nn/j0Kt8BlRe8AAAM/NXOy5ICp/QhNRfXpPXQ8JPpxpzrZGkfBi
wKQvVbX2JUVOs9v7ZHy/Hx86DZYoqu6YdcAunNdBTvJGdk8F+MgZ+6/8dxTueyKP
ZvBV0zZXggwxEFOY3xdXQXQK6Kd5e3vCfraJYQmiZIwNv1wAtceVhc1aCluz9gtA
RD+EY1cEO4li7KCpA74I+04I/YcNrjATy9Nx/3tPK8rD4aoPswgUls6blPURJnAr
dx1fD0RdqtYWiA+ftm4D11D41Aq2IZ9BfmduBpJsbEpql501b75Jcmx/wbn7SBgV
9oZ3YumC+cxenpcCupgR6V29pqcmPtfuy1FlgWJzavvZFh/aNGTb8CFMT9LzSaN7
CKmUOCrXXCnSr9M39EvnOtT1f/J9w+Ik+3IrWVisdr3ssxObr7NlyB3OWgUDsqM7
ujYDnHN5J9us9QPIPcc/677/hv0BsuO3Kx23sLER2rjZg/ULUWy8f3t/rO+9detU
ij3RtydNbo9fzHDnKULiubAgQgc8Rbq3vsX3KOR+jPhk67j/eH2aVz8NDQCwE4IW
nM3rWhpgJ1NUdyj8h/VYJppSj0Zt18V8yjm5+tsz0mASqiqxRppAn5zta8z9KwPD
ctLCPFFtfIlPz0kMCAd0JcIXi+qA34xhJXfhDLWQrfFAKl6DhoAXC5xt3oaz2zR7
jHhyEBGIZjV3T76y6iGSmmMQsAam/Dzt8XmVUHdGGA/sVmMawGkalfUTawFDGQsl
bQ6LvzTcVdq0ot5wcbF/ETX1vux5IhXFg+oJCphE4RDpeu31Gm+0nVOoJJDKdg4t
9YHaygGqu6DPVSnapmzGaJmfIIWRcfeUvtHUvvkptWon+tkLllyYHpc31Ng9ydji
CI4yH58ZB2chEal4oEQ33LVPO607ZRmdCIlmLWqf7EI7UFovfy5AfP7H0AiWT/0b
NFGl03f6d4jcLqjzJ2lnTqSVPukF8mMKYJWmy9qKWi3Pkk2u4Zm8XRY40VTaBJle
WZGGIYudGolCaAOOXozSe92wzpW3km+uXK9EDdp/M4BYPUFTi8kQkROJjAqWFS4R
7wDWDEhCggq1SAhqElcrDK9Rd72fPE5e2tE7cdR1UmJ0e1U+YGYx+jim6lmn/oa9
Ui1SPWRmGIt1mhJjoBcmSsVWT6jJElaGLbiycWUBpK0cnAZOZ7YVUD6cnMXHunH4
NxgMtiKuYxkIxvTJjFdNIDAKwsWIB3zvOTFyR6525N5o2NzioddPsZI2WIVgy1Uy
XENB+jYsETW9ArOIpkLKynvuiPd8JYpwpxah8LyLPl1JMqjEFdrIXe88M5s6t+6u
89IjIVt88MCXaQv+4+VvOkcLeR4sLhIwXn1NDqvfLKB3YydjWOPtMdLTOnalPEC7
Z/qMicQGnaOaGuEzLdycL5uFmn7PdtuGo4wY3cZrRBB2UtPYFZsAoNOA5VcQq1Jp
6AFRHgmJPGsc85zmR/Bp+OhU+7/LpZ/2KogrHSaM7nE/U5RY+L1/tHxY3wBSKl7U
BlQDeXMJqJGFMv+0pkBvKDUbFYS4X/AlC1CAo/71u9mouRsRZqyBNUS/TWr0uoGh
nOVtrVrhgtIZNLIU1sXUAKDQ+ai1mu3wTL4rIMI5Dlav3eIHGvDI3x7rKAJxD+ez
Y/rrpFxsunL1+XJ/l7AGvpsBo9IFTgXWwtN5FGa1wrElt62R/mrfi+28DO7cpy3X
Nn/TFrzwy/ow2wyhLV4OeprwpY7axtS3YtUlB2LbR6zsBMPfEVibafb3NSdNC/cU
nx2hXXgm2hgIe0Mx2Ni1w7ImuBImfClb+SGUfc14AKuOGkQO4MWd87vc7XfpRN+W
KHsCThMCIDUxb4NNXqQFGdae89kByfWtVZS6msyh6fHtOBy+bz6bwZfchHtaC/oK
UGr+K1NcWDGbOPXllqbmEEAsrNEqstaW+RYgpPIhZQyfbVUgWtPGyi9ZA4QcgBPE
2oHvmbaTtJtcDy2mx8szy4hB8OV9JKwVaSN/I8Yccp4WCVzIl4ZwUD2h7+GGwMrF
q4klGwCTiD4UhDlFghixX21J4zKYrJxHjdCbl1RQgxz0DkJWbSbJXksBcaljwl+6
o6qWtiBHxu9TlU2tvyTxPwluOR0NL0ZYdx1Oh3U+940EJWUmBFekpJmRlOdXC+cA
UmjAQNy8s6OXXG9TYChX389/BLaQ3PKRTNe2CEiHBV2pFDhSXKHdPX2i6jhIvNrf
ByixADgHyrVqHWOXuMd2NXcWAJp/vU5KnDUCJBKhtMxfSWya9yqBsYrEm/+C8+mw
/CmRp65Vl5XupoE9GhyDW1LEb6/5oi1gYrni8r3jBnShLeOtp2b/0cHTUjbNRz+C
Tg9w2Qd4Hjp2Vxb+GdjYQxcWGkgBpbaaUx7MXx/0IsDyaP2WxEVxOfAilKYMax5x
qsnRcFM5tzX6hVnnO9F6Z0vgBV4nrGQIT7ePgK8Rigw59/AmIqlNzuuzYA3aKQjf
NIUzZzEkpqLhH/cpvwho6+5OjqY6bcm7V7Ft2i6aA7q+slj11kLSMaCCuIhc0wYK
2VVijsZiAN6A4fqg8pgX9jkuMh7so9TwiVNC6A/w1LUEKF9lIXRpfZusqEZ94V5G
Gbpa03CG5c1mOIJn2j4P5UhwKKW3csig9DvopKrqo5Po9fj10Q+QTJubQVxW9DM4
Z3EVCN5L9ojqxahyM+xOsJm/D8rm8vhO3bp0TyXOFAF6Y+eMq6P6lQWRUBLGcKfr
W+Nlo+jJGczZ7NjhoPsdZmFCSI4kGeVZ08nYtXEDySb6vaGkHz9o2qDYjWagC82D
QBjKOOQIFI8gHpncD9DIxj4O0qmWvxHeteKv+3yTZ1ECAgkx8F2TCOIMhq92JiPg
WCPioG7Yx5VsYj+OenjZU1kO3njyMy42nX7P6FHn4CIozs0tuSeYl/mpYZSA2nUo
sBUIHSrr51vywbZZkNqA4IZK+OnpGwwzBPEGfT9kSjZrMKc2UF2uPVGXCi4GrP6C
VuJpPydkd7LUzmipYEBgGSFWd2qahAHW+8n8IgM+12IaR8U0zXuL8TpZlrpmI/y/
DvPzXoX6mks3lp8tU1/6Mag0m9xzmBBbgttODInXdtFfVctvRziwp3jQHRqecMds
k7n/p94GFnf0fBJpr7fu9v2hsn0cHrlqqfQHtzGpITdW6LJ6BoNqZBdfAZc6z8qG
aX5lUFIhjacuUqElxpmnX344LPWleDQPkYmv5U0JU56QaSeflzpE/9kMeciFYMIv
dVNOBWAHzX87aoEZ8zFFh32JDAsnJxEM7E4T1l9DOG6Ue+66QmZ8MituKk9R+/AP
3J3fKh6pKHs5j/8OX4kg6NrqlXhdjuHNmw58UiEO/BYvqMsXIu6LEibbMa90URao
N3jfiP8QsKR4q8XSiSDSI4EVAcTl9KCmtrg2h335Hf5JnhmruwSzfxBghUZnagmQ
mPq3t0yJnzxOaVEUrqRbY8Qmqg9V8Tuzc+wv+oHjsJlMuXtKGVRAi2Gp55KqFq4Y
mjZH5vg+jgzA0/39xmVGOP91xxkc5n5rHuPxgb1IFOXfsFOFJaNqyJmd9kyqPdDy
87HIfiMp4KVUJzzDKSvf/2VH8AIxYrNW96XLlZ8c76EJrBvBzD+1hUvUFPSe6Zh2
dMBW42FKgZvL+IY2Lf5axNFwx05E/36eoIeRnRTNcdD1Fmu2ELMmRY44oFb+5J2x
a3cq9ajiH5GvC7tXtt1phjTscsRYx2UnlzCHO2RoAFUwUQZPif2Miq6vaa9UsRQ3
kXX0Udj3QvAUOkdv+nuC9JMSAhZJ1MWobV9q8rRsEB5cXQJSGcN+ME/IlKCi6k1w
zHPC78gHt3WKNRZbkp04nfSjPbidBUMnHXQk7Qh5FEUKcCNvmF6/lsqeB78GdwH5
N9WmVUAEC4SgrWkngyCTREOgwm1OnuJIw4hGlzKnfdCJ2FWfuSAoxGDsQZpEnYDT
VJgrPoBppZPcABvT1k12gRovsd+1JFUl356OKClPk/47+kckh5JL7woYr8WDz8vd
w7OFKWwCybE6CtlXoxytf+Uq3RjzZc5MtmIvrY7w8dZe2zlwyzdaGNGa6iJz+XXc
fdZVFGXxaBfbEgwqGTarSCVbzYiKCyXupYfHv8uUc0ogFjCUD6Ei8iUPuNZgVkf/
cMNHVrxxCjHBz20W2maSKKkLSU/6uCnrCtz+1nvjq7299SzNYOyZrRS9PQYUxt1W
Bs5fuiCHyH1a9lNrxe8bvTGSKeeSVPSTx2r1qabUFNqWXBhGfSdwh7uF2p8rXLr7
qoJ4Q4b+7+QpgNGLJ8CnOCAh8l1Pp04Wk7z2KgKVheRHGwQnBWT3FWvT+TdGCzXk
TKKdJXCbz67n4/GqIlhsKY+HBkJLOnztpqsA1CFF5++OjLdHftsEQMh7qhVKTDmq
rF65WnpIXHmmNiqORrnDo42AOX7ZK4hCOPnlCeqTOSYvDJ404W4s+EClVM6tfbdi
EYcqQiqR0EBwrnZ9DMi2QoK60UAXK786w5joG2zDJ/UWGWVHhOQfMpdExaL8yZ3J
58Tp+JyJYgfduwSS/o03lbr12oPwjYS+NLLD/AnUQjnZ6/3XDvrWD6HqpGKy6BL7
cB+3TkALBIa/rDMFkQw3uBQYwMc4VGp+R/P3jXWyQLuS5mP898xyuBjIMCZMKnjf
0BtYJDI3H9wnZbA5ML0tp53fbk63PaXFT+cHNa3zntYdIoD5SupRLpPyE73iRdtl
raWSvwOWq/MxEdpYqppMhBn8sYaDZdD3PLS9k1tRlkdaSoeWXXxshzob0yj2tlqd
amhy/WjWwwFupuMaidmjiMP86SHmFl0M85lU180SFJQz86bPDdlkziOEFRXaajcM
rNIQ6I7IcdWY/MnK76qH49OZl5dxdv+qf18P2eHAJh2O5sIetbTWJ4qbXupBvJeX
45uLUjs1cMXdPeSbbJziZPy86iFYepQXOv9pQ3XwC4f3AaxsFCh2MDjjrUmJVHZd
PencpphxgNj3bZCNmex0dYsKgNiU5Cv7L3uRhAPktGWsTFRXae+4PGXoV3nBINEk
aCERV7xQN7N5APBU6zVjRVGXt9TlXS/v/+8FxQ3S6ioFx22K8eCPinmqoTH3bcf8
rOeY+k65lr1E4kZ/e4L4Lgd78yjUZiKNbOcGz+xoQjo35Ig3W2k9qK6TF+czCLSI
TNuJHQNLzUpseh/63fEUWPBaYjgqZ39Yq76rbdNDSqTGWFyLgJQZK/LB0VvxSSAM
xSFHMD9wsk87eeGH6q/ar9F/Y6y8KE3h7N31jGvI4dLYHBbqD4Cvqhdo6y0MZJ/C
/FJwmv0RKqx7N+SBKy8Z2O2cnp90qzX7ZO0o6tGK4s1GLP5zAah/h2AOTzZx43ZH
jnR2xpi47/PyjbMWsuLg8YmOYR5ETmsxvLXqu/wYNIaACrQUXeUc7DPWGbEf3Ap0
o21HvrgjUF3+l+YZ+QjUAm+LUvQebrRhbrj0xW2ah85Uvo63reSSp2BxD0tJYSSD
6TizUvjC+jhkkWwV6KLk5pPrKpIpjrFRO9skTB3l4Iq5Kq+56cQx725SdVJAj8MA
0+WTTQUDhw5+SbGHgEIbtUaGVP3/iP5PfYKDLjtURU4i7k4ECsAPy1LZ22YClF/8
vxBN4uSSFjeuGf4c/DQ1A2YhB3i5Zi1u62Hai/F8ep5GaqzKLVc3Ry96Sza/7IZm
e9L++liCrmdA+bKp32YbMwIQnTZQdlPUx2eRv4c2ZYmfzWk6wvleptXK8Jl5wPgS
PGjcvBVVFQEKV0X/atWP5Gs/ACyooidJoiS+fBDMAa8Rwd7SYGv1NKBdIzleih6c
EddNvUKXvoeoWQyYqMre98rHQGbFdN9h90nUhbQjaO3/DyLP8mM1z9PE+OlBeBDQ
n05SmOMHGRkjPiXQKl2Pe8FpxvvfBm4vhU2JgFJFiX6VRAOHch7q9unsZ9h9/2mw
zOZf8/jNdOU6uWdjqBa5zGp9FzV9QJY7memegxkzU3YBSXu55i6tZfLlOU8tH6Ai
gT2m7ts0vZk56pK/K0XZJwAcMQCUTDcByJKTtjaKn1U7yk7NAn3CkI73BH/lL8mn
7Fa8f+69uFGhGRf6f91u6bxQP4khfVMpfW7yO3feQV/9qS/FVlQdBysFHkPMfhAj
FhgX2Nw3qNxeWJT3fkQ0nlBGRrWVUmpY8PRpMBo6SmTMso8HQge86Ml+eC7BGPIY
FCESGmAeDY3kxd/+IK576m9piL4aFruiXj7wUXdW9oWM9/tCKF1mRArkdAnj45PZ
x7RaBvAYR88qP+7yzYhnG7qYBv6e+0vY68WPpK+ZT84EcFfFFK2gIcKj3tXYtXch
991f2qDONPI3FevakcYuW5z5ojKBHNOOPMx5RHkHB9EbEghpXLVWrqrQOi27juZI
wEoiAvWGPTxuaJA6HSr1EWOO+taCJSgBoOa5pObzpigbvaVe+1QU5sjMpiz1Ak7n
njPL4t5q5PN4SoH99k+LuxWWanS4tt9XlB7V5aKIklzLUlwFELBQrDyjWe8gPL0o
AtjdbR/ci/6gMEXok4Gw+M7eNP/1e8Z57Wd2Pidtm2EH1QR5UjdsN4MBk8eCBw9U
OQp5Pl1S+i+htjQg4GOCPAfBMw6rpRa4ax/u6+2OMOFyFP9b91kgZPkPIzXsSoF/
Fk3VZv2+lZqxF5bSDs6BAFENORToAPG9IH+qdTX4P7oWbQawH/OoVdrdFRhVLjpz
JIzKd4wlpooJYCSKW+ceq3BYr+FixlDCF0IHlqjZf7xTABDdeS9h1+TKRV6xpRt0
RQcnfqH2XKHRSK0K9lYMKwTB2r6iybyGJAPosg1uSPAPhHkP5tKPOj1GAwQ+sx3n
2GhsU3TDsLVsU9ZouzYVi9PbCKCAGjBnHZ11U5dqknT7RpInSXJW0Z+tEm7Vsevs
TX60mmoKsBGDX3M5/viapfIZWv3anmX9voL5JzHTHnBdaC/lBZguHGjyjEVx/+d1
YTqkmQa+MO8JnFPTzxgDSuMweVmkTlom/XrCI7Tj425L09pqzGEsgL0OdH9t6S2D
G0zgug1ExbG9l7pyCX3UEvzu6Vsp7hyMeqkRJFD9N2SsTAVMj6nMsoOz0y5iurax
jvSRMPYqvL6sSgSU/PsmoH0doBvKuoNWrJ8Y7ey7oPS0Lp+FdBspIm3kuxOGOLSq
HIVbM3RH5LXvAySqJIbvx91gZFXVX9GiPF1wEeP/2ZoKtN2xzWgkzuagUYJqWW+l
+PgxvnSO8nEgUifZgl2g0XfwUwGlnI7mCXflfxS3AyCtUQRuxrHMYO3dNrotL+pb
BK2GnxJW2KCRic7Pb57/G3e/25Jy2dixKCWCwhoirMjcOmrtZ9oRhcirR+SiSJOb
RXeYQ+oWZzIzH4mfzlJsfWSzFRl74rBrQaOyDi3Xy1uEiOr3xdaTZo1nVB3F8vdG
F6hJVYSRaAbJaWj4M50nzg97dvbkOVf6zweUs0xSABM5/Pbww1LE6ayzZ6KDgDSJ
FGoaTmYPOdD9bwu35MVvhnxS10fbobsrq1KONW03AguJaczS75FEmHSr0B2mrqv6
aFHtfv3eCSD23F4B7mMcOoOEYX6/02iaMeKwF6OTW8tEksSQvlImA6Rd62/i1WJO
MmtZEXBECrC0pkUw+yFMOwZ8pTU8+Gvy+YEtjb4pLMe10ao3ceNhqfByW2PpAVlM
x4j/fpaCcB3vrdCVDfJ0ilxGKo/8LV+uhRDP8em/z6+wXxgmIoXIBolp12iaJHRM
GnqYeNdVum+wL59swosfyFK0LCYsFjPwW7m2Gh6jFv53PvcCHoLGj0VB7kKOo5XH
JzPlrYijyk8e+4ZDMBaUGAuVLR0mAEimK9XdO2wfs9YXdyqeLXlzqayVzza8iISS
NBO79fjpbjhKffYI0RskTnoZsDj0PoqTPq0y2maEPwgeBFnk61J0jMl+q0fi0cDx
5LbvixfZE0Je22FdM6W8yRGVuG8MXx61eJHnp5/BrOhslPt5He1uJ+zg0Y3XE1n1
tLrW8woaNHnXnllFYhTXy6Zd/8RK71nrwpjlZdDjb2ZknwB4pVHan00VdyxmDebF
SSGHKgjQRIs2d2jDUdiFtI6ZQggcZS0wzXXNaNMPyPlgGVwMZXlo7qXKLDq2mEnh
ZwYK9XSLbCKVU+wVkyDGlo3CVOqKaKp8L/cqCmhVzS4Oua7Xn5CKzOLOEQknwEwS
M8uIcb2ZracX7BL46szfAqJLv5lFwgh5zzUs/eQFSi0OOf5UO7ZB6xpwUhjCZqsM
/DewpH8tbhtfTi89Wgmn+n0UikkUrjiAHDZv7NyX/krlbx++9Z+d2ZcIq2c268ji
ZNNj6OZ4Ygilmftne7wUgV6iiIsGVXVbriBa4ea8GTIuVbQxCZC7GAMhHC9RNAMZ
RjV320tlUefU3nDgfg7KSN4wg5teu3vpVxuB7nB5kpfvbtHfhD06Hsx3Y5Y9W8MQ
J/9SQ07fKbzuM2ey2LdxkUczCo6NveNh7TlfFfGBILyRzVGgCO9vuKOWWn/cckQG
8TAaLVVfekKWH99lbXnFSRbZb9pQ0wCtgL6BkF+O47GRbmMJZfmrWgT999XpPDyO
ooyW0pghytyafOC1r8BrNS39uoi+kdcOFDBjNGe/4Gm7is7S0r6i6SRRxla+c/2x
LMUBxQFxMPt51tpWiUYnUzL7cYvi0JVdPe+EQUZoTRxZ9xAHeLvNscZJq5T9ooOe
425GwfQjrAZE1Kx8Oc0K5X7xn5uFnGHXzzBSkVjQIf+Tq6SElQd8lr+sreHFHlJM
pE0rFtGQpLzPEjkau1vZMI77s71lVQbhTRBMbtpJNfuHEEhEkSfobehU5BN953dg
ghJIo73+k1JBTrfMk1Qgc5/Jx+BSgJFTUiuoACCrLeNTi0U1fCONPh/OjAHSVB3J
Y0gFwc7JvoTqgVR9lsKB2qxsmx+NqQwsO4xppoOCoixKZ/hZOdCkw4+iSAie3a6D
E1Ba8qD40ckxuF+pKT7Ny3JSfDkgdobp8hZQyeJRarQpEer60ozhYTQZwCJ30f5p
qaQHXFyniWdKC9BFjCnqGrZfshkspj3UI9M3jXeT8m2jzZji7tbFej9zpwClo/oR
Lur5cDz3Ep7lszXg96j5zkHQjHd+EmBZsRViNy5N/3kDI+5NNLsC43sxKVSZyKDE
a6fj0qzdUPzXNn0eE2cpp+Jl84izZTJF6DXxUGq7UbRTN6mdPbjXeTnCKdDZ3C9X
RgbAI2rFRlSg6G61FG220yz+kPLGpuSHHKFBlef45rUfdCCAoXynkpEvlg656DtL
82z8hqn5ae3YgwWq2Pk8AIAx0zOcmoBFiTQtzxOPZMpDHG62eI6Ogt0IR4a/RJEF
NpmlUxgFj5c8qVdtyXhVBpGJ9fhczVnLXoyMi9p6ab8SNBJQ6mMrTS4op2PnPeq5
MUYao9iAqBW0uqbOzQn8gkwD8u6g0tZL5QkvgUHroGn3a9RbALjdrtMr6UjQ6UNR
81Ib0Ljzsw+qAZDrZ13laOaHLRZzbF2Apuv5Fd8b+xJ3dTzwnj0x6WNv0m6r8d9l
CnfNBMcyEQoXZhe1qFm/B5HGeIkcaDdzv3/qCAciPE6YezUjDp9ZIuiYrcPycRdu
Ocff6DNbBGrJcwCWqzBLz0dp4GJrVtrADwROmaXc5nd7A5pxa7+uaw+GOrEtEIUu
HqnS3x0d1FqwiZCRncu58dCy4V7oBpHq3Frbm4lIMSuEz0AV2DtzVHHgpRQsMb+p
DVv+j9i0CmPLJg3VDLuA6AXi5fsKa7eDIP9LJndba8Aq+c3+jHojw7XkTmD7aSfl
aECt86l0lS2ORsWLgPGt+7KZuqPY7Nxkl5wWONux81+nuKN5BuqqY8AUt4kZ9+YI
2cm4N0RqlVVPFyxAYZU/PDkwriiSxzUHXVL2zUeE2lUtiAwW9beGzegd/Qs/BLK7
vq5YzMxK9owXa32NCEbWl22t+Mh1S4tYwpujg6n0zbZaxvk8MD8un81PjNow6SSk
18okqmJHOtYheYxWWLEMyuotA8QRWpiQakc1iYy//c1Yso94z7uKUF5/ZbPFpsLN
LpejtZoqRvTO2YamyUhsSw01NFobRysBikfLihyPdYPlDrqKUXb3alW9fWR2naRi
jJOwHPhv2Ch1i+9dDnD6IVjxbfPY/GOXoY5DR1wA3L2tj0Sjx9HPC//SUWlFkROr
jszuTNtu7uaTwGZaGgX4H4SBOYPbu3+Sp6BT28HWCxcrCZsFUPAabpnLkP9NriNk
TLbAd1gSud6rfAzbO+8WY2eDP9ENIEKAf8DO0vT+7b7HJhsf++NqHQ3lWbmIeADF
qrNkr+N1tUrSRQMMly7RLC0GIh6jr4NqIZFLiaQWWh3Dr4e4FrcrT5ILOoClBa1g
KiXLt+oaVoZKmZ7SmereBln6O1LKe02lld/rfFU351Xj6O7ONME+W8NUK5tsDBPc
zG+c78h4/hJ/Bat5LjLWRPR1d3v1cfQT8ezx4+evH9aeQVRAhp/kb9zGVHoDw+HB
2BlD3CRt34wkg5E8SozJVPANDQJEhU75sYWAEnz2u21M4UhOVxRlheGOuZATjg2X
yW27YTx2+L+ZyDztPntnghcFdQ8ou/ZoTesgjNp5dUFszDP8E9hAO3w7EJEMIL4/
l/WtPlNStgRxMxe4PGMuERkVa7SSRBh0rZl2Gh/lP5YhWBBINT7kG1JiABGgeCWV
AK4JXmPE/AlbdXlniDB6+nbU498WwXTYXiqvZlw2S8yKpsJL7oQsGVQbKA8bkobK
5xkcBtBxAlVFaEqJ0lJp3oIPqUY2tLzdFmtmsEAfsEbXCl5UVq8E2AudQo5tKg5t
BTL/TY1EObtFai4QKeVuNsyjuHiuipHNs+ey+oQOYNNAJh/z8z0DkvpW2MZGleh2
QpoQPxp19qwP3PpUTzdYeR+/Wi1gaoZDm0nC91Nn6XscCqc9+UjBz71YhmOgmnD2
Zj6Z2plfuwuCn0keKLmr7WBaYYxX0Dih9PwA/70TqguJ8JO+3I1uKOD7SAzpEAo3
z17b7i2IQCoJ4LJ7TTfI9OsALOMrLes8qM1Lg8z78lSyJnjtyT/KAkex9xEBSGS/
LLJvTM1b1zUeuuVEh2iUS5YYQYAo4GcHoGwEGGjFyTI58CHmutPmxVjCAhh2xa6E
+o6F2dn3Yu9AMzTri6yGpU0jNopPV+Kk0hyBt3TpeqT15ZocxmUJyos0sdlLqlhm
hvlUSLahMUyDQTYGRNPjti1ZJYQ/maGsXQ7zTwtjWwWQey5cBLviHLJxEK60NEeQ
TkfQVP0u+htFDZwSu1eVpbCdTv6Ix9k4kmVd2/68gTcJahJ0174NK8LQtMSPW6Ct
AHrXrQ7hQPKMXZtYjY8nDFiaeXu8B6qsOBVWomPVE3Zyhko65nZrF5qV+MWMc8jZ
gr+oTQGpERyhmfoVBtHA8PhqdBoak2FgxP+jcoMU2DLel1ohXPme2FKymAgi2ec1
oPyFgaM/BSqfzxBLNRAwSet0VlKh1x4pQ00dTXQ/0bBrmKX0mxNZgPNCc1K5wEiO
vi/w5/DRXF/2cSwyKfiVoauhu4TL0Gz2IyvQbO/xvcekrkdwlF0ptDcQa+Wl0yF8
ZVZvEJZWjN6XhVyK3Szkkn9vpVOmrM/PK5AZAVV8eFqdJFcMY9D8neu3zrhSF070
LG/i2YzYhCq/4qLA9Vd1yxF0rL0uMzKI49xCI6sH9n1CqKMHTNNUf+4qLD2f5vjS
vS2TtYKPyZFqzxTD+DAQCfPu//TGE7LhZcQ6hn+XGXk4ijkMyk1Fsty1uVVnOQLx
zDTMNnbDoYZ2rL49oQPcjP4gGlPLq6ppV4yhdfpd2ECTryyIrvKBT/h3By7JMo3u
CCMsdfVmgOk4wlDcVZ238TOz/sWdIArUrDDzdlC0QbvQdXkQy74B3YKI2U8qmPzt
B9MTYTASKsygI/k9uZRpFZ8KAV+etGoWtN9nAE+MMAsddiHuPvZ+ng2KUSQszomA
gecL3WQ6C0dPrUBK8hzO0nrsfM53zzELBy32sbvogqMjqkbOJTDAeufZL15AQmfz
Ln/i/kOeqisJWOISO6shWqvqj1ztfrZb+uPxPp3bUZVsTw2IwAp/epWQCDyvlwlJ
cfWrSzfEKBNtmGE+AkQQh0qv5M3XXcelInFHa8b47Ug3sqcpjTKxPFLof1+6INfG
nZEyLRH0RZ/+23c+b/YW+TxTnI2UMwGs620iId5i+SRqhXB7BuAVqyGm4jJsNFn6
Z2t46Gh4WqvNsIdGhTq3w7/d3l7OeoJQ8+G2pv16RzHRAEWXacxlMyfAfh2gdRKf
l6Jky8sov/d1o7LwaEXjcgt+rJyvuegFa6CmygKPBlJKDJ7zDdd3clat2/bqA9T9
yrtidyXOqPnjerMaV8LBIvPsJVRxVt5JC/P9iBwaXT1XE9v0WHFFRXyUZF0rTIg+
KX6OjNI8tSy3MeAhPy+Z+YxUSe8/r8mGQ6fKxOLwFuonlCGjx9tqchsW2YeL9Bvm
gjm8qI6qIc7TdkjcD35xJaUP0clQMgRG4jA1D63wNyBRl/xuV7LF/ly6jI9BJ0mX
wDbs0sRw5gvoIqtUn8Elr43DkjiEXyqqKObNJmlLaqVc0SHK+x0xmV6DU5j2oHXC
EatYgZAEA16FzffJ7aDX0PnV6HFuYl94oR1pG3/NKFV3UXGOjrbT0m6sKj13RFhW
ERMVlOFGfG5YqMzgrA5QBvm0ZY43N/tB9igimw85TQjOJEEjq9mOVxy+LRs9D4Hj
jSfUCa6lQY02oBOsOS0Ll9+hIK5u2M8taQhAppblT9z6Xul9zyOyvBEwT4K+FM3O
0Y8C4ki39RXRlzDpm7JWkZiXXVqTeZTagdMsulhIxQhtG2ViU2f8RURn5a4CxzCv
+YBDS5m7nO+04TW+2TVlBuWeqCEpP991u0vWX4/NAjEc/HlF+WnGWh+2C3uHfj5y
1e8c5T75as+UDNbMme3lYuX2tVC7CQ0EV7IU+Ghq2F61bOVT2cIfuus2iJpxHqbS
UoiZyUB+gX1e6NcIYQSJBZPqCg4R1hR4lN1QLcqu1dxUPQDb7XmqnXy/zU0vJAH9
+4yLQK7yinn+6RZzPBCgkDjomd7tKnUhcg1XqgseYMAv30yMt7jtfbkSkHZ7ejW/
Gq+UcZ4rk22mtXl9qR5erppdEZlBxGWoiMlRflR1Huc8ELvaRCBdFzjqsBJhSBfW
31ptl3lD+VRtqIdQHr+bJQpC1JvlKgI9Ykkoth3fnIafgMjNN/uTtesT/dhBAEjR
BjJRZXEy+xdXlitzkfK9C5d+ZBrRFHts2lrAkZjo9WZGDJfhTxzP2+Oar+IeWYre
+a78cMDuUVznO4JXidfAUv73NSOFvfURfPUDsRPTaAeT4mtO8oPa0DCZ/wosmVRQ
PBq3Rd10jaD7Xgk1Br4hN10gtML217UpS8UioOnTj2AT1cGIcdYgarAk6FpA+M/G
Yx/z2shcF6gaT9jZNp0z4ay6f0ik6jyxtgdt1pFxgz+SthTkM1AVy69ap9UfKdRc
h4P6p/Dqjl/GWt6sjgzj7PzT6zYtKefwGEQKmv06rQ3TMEIYnpjIpzOdhCD3Y3Pu
YeJ5B+W3xwPAmhfAICQT/JMyGmnoWynnD1ixz1L8qXxx2Yc1elmKC+QqLocnPc6S
CBiwZ7x9z8skuHuaLUVMIMDd1oDohEL3bjpjOT2EhzveZfe6nEyYcujYu3m4xRii
5G4B4zxoLGIARQoHB6Yl/1Ni52MR+oq3jAnn8Mr7jzFNjla8qqxhT1PeYNtgrHKL
Ex95H/iYrTDjuBg46fj4cU6vv3CMO+TXTZa2Qm42IcjWZWcjaOnXbK6/XMPCN8Ps
gmyIPzKOPMhSQ1JSUJbJCRTdfnoJWrYNwjqKYvqgMNwxjm1jPe6GouLwHjoxiNTs
dDgoGfGwUejgUT3lIRq796GwLsDQEmXj4NpoFZVEyZodcG9A7s4zQBvRi8MN/bki
xjPM1QKPhNkiUoxCL8i0odbQooBLl50x2V15eQJyLAk4knpXw+fUXap4EEli/tTz
VnvS45nQUZ8xSXxlcC0nxoGtvivo7YauMzZ4/TEQ6/NM806qxfq30o72LL5ac6uX
UqDRIuR+S5nV4muTWNV60QljBipalvHqE7/NvKxb55XLgWjtYtNRB5mIjETGhFLj
E3/tBJAllbdCqFqDzrvUL8V8Jo0SXgeX885jZqYdkvaG9jwXnBfzC/+uQWhUP3yG
MR9tmCju3nt9jLnwnlSiPEy5lvQRi/gcJQGbEKVu/uf3MTG0AkPwH/Z3u+7Gy41S
DhzCClpoJ2IAmGUgMXH1cIsqjza8HaXG7cmtFbTGPB9JqQ1ZIn+HBUo6nXHakeMg
2XxwNGp3t/LpWpUVSDMP1BRwolFhbz9ZIiyqDa7XLT7dc/6KBMJCeunEM2jCq3mI
YpuENzkHxVYbXS6pq4hP1xlnkwLSSLRh5ft4IDUGuEv+9k9TRhwNf/Sx7F57OVN7
w50sJxtGpKUXVOw+u6z9uVUTSq6tPcwr30/nbL80xZIwjQM6AkCWSBWCmLzx0QKj
mEn8rNT5mYppjXvj9eH2yBeWU61uh1Cuopd4CSr2U80j+xpOv7ro2GW+go4XfV/w
3Bv56uQX1Dqr60oTzxOaP+pyX2EK4Hw/rWNNxG1xPmLrVeA2nXUTA80VJs7ci8Id
zQIB4gV6fUNJve/zPOdeJT8ha3iuvsRkgZW+mpynUt8AipP40JQfqiOc3p4B3sGy
2viMdlYE2dttJvW3sJV+v81MYzkwFmZCELw7oFUXD86CpXnRiaP7zKDFdIV6FOBN
Tbf8jlB5BY8iXPRaIsxm7FtRCgvURSFF0E+XzaYSRGr3ltATZpHeH126h8R1LGdB
uRxWmJh/SUR2mnwZ9Yss0gAgQyyFR0fZyxl76cNxbSpCWDxd3AohA67sPIHe1pBq
ftqJCqfl321FdnnnmQ3xB0314OnbjTbZ3Wku0mxEEgda9aK9s0xo8Ja7y690d4cV
ZSHCIC6/fW8vGbsdmOUM+IMBV4IaQT08nCgWPmkBaUPufgCUMKcT7DbRapLnpg5k
DfNdTe7HJfvgNl8bQlPjoTLah6gphfa3vyNXJjHIaAGD/BEXktpA6UncFL8zIr3u
zIha00dNGGzlIfpCG2lCAROELXGwVcWqpZ7f5nnQRM6y5L775MH+lXM1Wuvo+Yqh
PYDf8ihjAc6zDQ+oXb6cUu1U/2eoOF61s3vtVDytJQdftvFyci17wHgVuKiol3XU
yeXhOrE3hPSohlTVgHcV1sCm0+PPJDuG/SxhocqSk+W0FccJjtb30jiTeQtS0jJ5
cXBlE3BmtDMH41xht5c3SZJg5K6sQK/tEoA3nfX+jxtzfOsID1BLPPVbHF2m+KY6
/PXVy/wpP49M2LXeDdJa2fNa16nDbf7PX5XyOLHFDo7W6VojESME3eppl3pe9Zdr
6sLa+IU9kve+2TTBO6LCYfETvboaKF1XP22uWhhZcUbdKRN9P8FI75pSn4kGWukl
uOHeNIwvhzh0eLiXN7TfNELfM5AaS6WQXH0n5lebHVCUQx++VZNrAj5dpuDtwd+i
++1WD8Q03xuo5Pt5hAe0ip7G9c8rnXPi1TTF+pwI8JJS2RUHRAPscvJx+iODUaT7
kw5e9Ns7FQU0f/ky9qMBoKHUfy71eg5D5bVltWXvp9lIQSza8iskSEYosb0VTf4l
x9dqs5L4w4gqwbPcXJJldlsN4ssTBCyGbBvQ9pFX/NYsdwoET1Gkw3BqWXte9cYd
VgXzVWtaUYqexdI+bqBhej5x/o0pxSsfFriQGsIJQ7vjrWsmmsJQCDvkk8mzSyxh
BY1rpzJQdzg3EAq91TKX59qdjd9h3Y2Bw2dLzgIK8M/Cl3jh+JdWNYsu4HTszqUa
Tbh3J913GmYvonDs4pEPvC+wgnTQ7JEDEoabhaPpSjNyqA73t9QMO+ZA+9Zlyed0
62P9SfFSHLYJsl6LnHKCxU71SIVkRV82xNSRJP0x/cMg3CG9UkI3sdSOs61y3ona
Jv/dPDx2ZhQGVYOTYDET+WgWa1X1Nl1zxS0Wm765ZOCqdfqmrRUYfkqwUcgXc30l
LU9cbNFAyx1mjB0aSpCc8ZHkOLFWBKQj7X94slMazWfn1q5OvPMTaNDy8WwvXA/f
Iv+FTU54Yp00XWvxXGls9le63b/rmzAV/0LEDsq2lp617zVhM66/1HP49cz8Kslz
0wWMMu4Eip76prqt3c0/YWTYdleVm26U/Re7yaCleny7kwr7YkqTN9HUBvNotwMc
QBMz2ntMqV2qlwccw8KzmGe9I9kWVyPD+DNTsHDrIXM5p6nT+rLxW9zCrD8Q6j03
hOCA51t0gNkDUhQd0YuesiYkki0cwWD9yz1fqE4zck/5XBbYCAjQnU9vRhAaC1V+
jerneKBN1DV96BLkrj3SbLnPqBN+VbRjD7VrZTDjx5tMg2KiAeyusqsaCqfekduN
STy8xredjAdw3bkOWClhZ6a/R3WdFce+J+qbuH3paHeZJwaQuSmJOH+Glj9+F7ID
lQUJv0oJ1O28cTGDEZHTSYgJNLjU23m2uaRw5L+CR9qTpDBfSsq+M+CcVSaDD1lb
H6G4eZ9iY4XottZhumZBLDzsBQ0zV3/Au5uMq8pXyAeZdYfK6RBx9gMRYHR98hsj
ZGOh7UGDyJqAAbynyhYvbuyhKHxItyff898/EgC+Da5PBZiGtazFqlXS7Ly33PAn
f20odVwE6ng1HATCGlawrt7bwPHzBRgYsM/szwDz+85gG6G/s8tCrmjG2bqQVszh
OwaJBkuXQo3XLDHBQ4LlJwSPeWZ9bU/KmH4Z0XY1dNEUw0pLkKs+RpgADERyXTGi
4aNit7eiRDxG80j88AuCVgImBFNGlc8ff4C/zYL3uBqNGt0sN9At3c6GYgH6lHnr
bls9JC/442LKllWrZzzVqGbiD4vUoojXAx4l268GFGhmqnJxpCiJGyYHZGxV6QjX
rUSv8rNOn/k7+MsFXf89M9D+6KySKvaSUK6TW0VM1QONzJJ/l+rydGIu7Xb9CION
pBlefAr2S6nKcgX9FBjxnniuliiC6o8tVUvUXubMUY1GhXYi350W+GNut0H61nJg
6ciBEv5S+UH7jd5O+Hb0jajQFW4Ck4ELlHQJ5sKsl3REbGpMWeWXDj3haXXRd45a
c/lO/UK/mSdb9chZbAcUchwrLIQyGINj7H26JUVujFrsXkaAVs++Wik7vd9pcbRp
/RECBq5OPbRy/tTArsmzigVB9QQk3VXzCaYHdu6nXlIJJqp5lOd77PH2tQn6N7J0
Y/DWC/KILPygYMreZVPeum4MXCrtFl7jNrCMHneI3m7Va7jth9QGJsHGWzWYAxrg
6wAABWCsply14Hjqxj5Hbv5mmxqij21UteAmtshqRLwtmnZxlDtxj1ZGanMdhHm1
F5CLBnv0ELjpdaQNvXM04gYTctW+Po/AgL6YmTccwE8emcS8ULs664BIHyEmQ+a3
aRzkVjsXUoQdvPxy1K0IdhPTl/x1iuH3Ks2WIq4vfzGcbAcglw37NUs0r5KXTMf2
6RP00o8uTdSAra0v7uFig0lAqhndmWAkGKxnoPuPP1Grj+Wzo153TSn/K8IWqHQl
wjLVYTZ+ETZNOu73VoRA7bz/zKeaLdgMIGbYex8fGi8q8XQ60EW7IewEmowK8iuv
7yuUOCwbrlNBycCh6CiZWTawtw+1ud5hoqLtjbKxoRDBHcVwjNDsfCqP5X6DN0U4
8VCumm6zuH1BU76yQO1orhl07P1BkDstK1Q1e8H0t6X+q4RDVD9FGsB/BsmQ30Cr
d4SvIj26lGtd/6dGsDqLXgTIIQHHc45wfRUkQ6K2Goy4GIlFw5NMgfq4wx/e4I1Z
Tv+wdR7cDFCSvyB5CaIV3qD8+7O16rU518uGr4HYovHbpe0p0IJ0esA7f8IEndAW
k2ouMVPk3i/+G+zigAMEjjoOWK9t8ovV5Dl0eONdGtaCMMky5nhxh6vZGyWlhfxU
FMKTVaWAgFhFRKh0GuzIvg02mSbLdVF4m+vHLw8ZTyJUkKL6i2nB1RoBMvI9XTwj
hmbryXT7EKtCy/8F1QvNn6K8nfj7SrXEEmhSzQu4Ol+464dnb54IgQNz/7GvwMI7
HgJqksqTCtV+kWTYW2iaSDz9ThLfi2YW3N2oY4wPEBYFlwgWhvh1K/dUkSnySe2l
kbDJHDltDNLVYh9ttSe9sChQVs1Eq5bc4ITRUq0ZCOPyDdWmyJqtYR9fZuAZA1F0
daIS7UXM6PutcrnAJBUyjlV4bbvor88nzJ9B7DlSCBZz3Pl0c2E85ppCWYNgAjXz
4CuK1G0pURLxwnMg3kfNY56rG+fQsplXZnzfLBYeWFVpl1VD3C5wpvdAEVdTogYx
HJijH1VyY7lAal/oHDygE3MJjbOOBr/SxM68RuvA48VHI1juHW+8Mgq9P9wZisOf
Qi+DzevZd7qOVO9idDqpx9lnd+FrhqMKokSecdsJl0NwNDVPUWB8eBMDAkTTXo2p
kg1ZTl93B7A7TV4WFs9TOBIJF3cKoa0B00QKBhnGBew8gtD2qs2Ks7m+eEQEJWyX
FHXI828H9+Cj9Unue2F1ilMgnCf6klc2KwqnBIAts3WG1ms8T8068qfTxk5ij5CX
n5NY63dQw/9BG91JXukLLyhqTuMFJGhRhgL0W89rM4jfDY4xrfFqrPIe5M3H2Evw
RsjoitiPscdqCkKTsWjd21/oAGfuQcEbeenGjUI+XjnGP6uMVL7dYVv708UbbVrT
sAWll42GiGNQWLCArPg/FynM8lFo8tFaTnMR3rSTywlVpp+WKfui6IzLiD2syiRT
n6CX0V0MYfwwSW9lq3B21iqvajjraw3jn2fCsVwfK0LW8PB3bDsC5hiG0H/NPx+l
ypCEjU7bBrX1IDooRGfo6ibr976DUwmokAZm0tfONOeZNsxlEvacynaVedgTL+3h
2H7XsgDjEeVaK7LMyFMdOtVC0Emy5LqkQ6+2Uk2YGw7GvNCwKyOESYtn8e0MAQ0C
mHRk0VIehXlQVKAF2T6TCu9KxCLEazxBgtgP31ntey/DmUgT7bGvW42bYPsokdRc
wFeynsW1Nk6eujuFcJzXHu+IU6EDnEGkkPe8HhgXGbniIOWlyjyAKhUDpZkgClrN
CPs3jv2nrKUjnEP6Xl8jadMX26lubTk3m1wdBQUuySigW4MWEo18NWq6A5b3SnDA
DetjsGiXQxmIpVDHp5j7c5Rk3c5BzFWMFnFmrFkJjFSErlgwiaZFIIwOw+QO+xg8
l009rkzXzjRBUiVCWZtNFcX+PuswQRAgIL9JkP77hWcTY1gkE/il7Jt7nNhFWHpK
HK8ZrCHcR3m2gbqRpglhHQM5PlW2Bre/yhlrxjoaW8YEnmSnfqCTGJybOB8v4RpV
pWMTO3mJMb1xhAzZMBVWOEkh73I546Qrkdo/5eVubQVeKQbLgWF5cWU7Q5Oz0yNo
z7O7W1We0VCQGpYPBKthM+ILne1WHcvsRUcJF84mXa/amRmGVZ9PWwXOYbknxvyX
0b6VMYFynqz+LoDOB7PLXIRbOwkLcZ0W4ol7sqWqb+Pi23OJsr6dqKkyY40IIpfY
F3WUW+cp2yWZz5S1Y6w+JjfUhCfglvhOrzu0GbZqlyHvb7eFuHNkboSJLoofUJVx
BOndOB9v3kHmyt78Zs4ntdym1TO1ErY53/rMf2O3qpeZw5zePRB1p0Zx4aAyNry9
9+6CZXpTyK4z7JeTqYFgVhBnN3mVgFl8mXBtPYShQCMXzT4TsJemvmWkWHEe1qWI
H7bJ2CpHhe8xUiA1Z+TB48lT2Cavtqc+mIH71F3onGOk+yHWpul8tih7Vb8z+G5V
hAF9hAonCRj60Q+XD+7S9bZevYmo6R6FmnSHm7vfEFiBbPIxlL7i2AbNL0/Bgd4n
hfcR+8WsFof3sc+7D/aYNbnufs9Z8PGmYgRuJhbbuVbE/TacZPnTWIDRX4K/AUb0
3VwqyDytaoIExsBhTJtTrgluoh1SzAIUtwzyGG9a3dtgWvwvVo04LzlCxJBrVfrb
nJQ2NFy3azlhkObfUBohnDfEf7Klzh4QlwD+UT9hOKdPoweNRla7Zjr/ifUhPWtP
X1Xk51BEYUuGF+YQ6SxCFNo9xf8ZVymfpDNzW96/YGhgy2QLYEMQhiKaOtIEBNNQ
vRrS4/ZwzGskmjNmksuJhACiD5SSQjaRXCZGNhUWPs4i6O8UzyME6HeFREramJOP
rXS27Wmf3H0ixOvDeB7KWuoK0cAwhs+I+2BXvaxFCzFC1AQf34i2D7pVRGUjw9av
67e6+kOCszha/LEpe3uuKglOKeFEzdUL0U/GgH/7xihBHIiVEsBBsNe1RHjMMat9
1RmszEpvSXWeA7sKxU0L1imy540Clf9UcjC4HuX5jDX/v27ANzaOE4YoUT2aobKa
kahy5A6z5MuXvVJE+0juKQ3YPB4rOtfUFeUJugNmdtTJLoHu74WGzRXu30/ZA1Kr
x4YXeqdDNPySUK5z1tK0ewbMKXqhV6xVGICRatVPJOcXqFROzYkqHjtoK3TXNmIC
pot5w9IETWQ3KsS4cn2FmxrnNSPqL6pAV93CAihMl/VimuLNUuSPi55YQewj8/IG
9YrGDSnhw4uoWTX4+SZSdZ2QF26mS+XDLQSMVqpzkLDSaa3Ttuv2inWsxzOGjEVA
jOJDOwiFMdpYF92AJbcgFmUt30+ZdcaCSszRjuAjOqIYQKu1t0BiI7MVPfF12704
MqZcGJ5wcOI4K0djMSDqa4yAnFxLr5lMwZf7Ro2K8py8izq4kJoj2mrBPat+Ef6e
gB3bivGIgN2i7lXoHfq6pTgoGX/WG/gaqq458y5b/LJUshN+0Iv1bWUgIoz2SBcy
cXwiaZEapy+XLvwPCcMhF0ZG44TMMNoLbTh2Yge1SXkXkFrlQkxJeTwO9iaLNQ4K
wuQtohdelxiZGM7t8jpXmCev14jE/xYY8j2s73G4JVfUTTBgkqBgFQg06Hi4gPD2
HpJ3gPrtHPH+UiEFx6LyceKEsYPFJSwxzXj5giG0VE/wgXWl0NWZI/RR0HmEcxvV
8U3AVn36YTRiL1+aDliqolOq9DSh27nTxOZODEXv8ShtdYlttZPR4L5u8B28hFA7
UL0fhw74g6xVi/XwjW/K3Ct5fF/HAbV4GGYq4TmpPwv4ckWwr0VPnBXnKbVxsk+x
XyURlFTN4ZBzefvJ1ZAfQ7VqZrFJgfXbmfEgR5RV4Y9m0/1jtZynGD1HQajrAsMS
ztsF0iduGsiB5Id0heCg+78PcA3Vm3nZcVKyCFNnzMvsMk65veKcfRGGH53mFk2N
jF3tZGiUWF1rCXfSgnPireQSKu4P1tU5eLueD/opKhE093VTrIzc2bigiKxgSYNu
FOIxW/L705/tQWAu5Z2ypIy/n9wJvNOAAzgngtRhlsxtqAjt6/lDqbsy0oPY+hIx
JiAQ41eM8cS5bSNd0CK0P3pZHAVJ28wCSn36PFuL7ZccZiBDDgYIjfGYprh0lZsb
L6UnlCOhPNKbSSiXRcxApH6EHInEdMoevqx/XpIf6LvPJ95veCgRn63idSjiOdNE
qH8JlwcGTL6+x0scHZmOngSalGcsz/iU4xzSzFVhvQ7dsGpjO23Zggj6wnBN+tBs
tz7mF98MNTCO6aYptlOAvClxplq3eDinkcdiWXE2q/ty0J8kVorHK5ZPIX6UwMbY
9ExsAEqKiiW9u4hhlwygHJdvBAu9kkjG/bGhRPgapg2cjlnzSaFIHB0MzpdLdvFR
uJ8sMeoenP2S5UGviS1wEfjvax+k+nSbkcMS9cDfq/TQaenyytQ38C9GabiZ0R/5
OUPt8VwJZChkLx+IwBlMe1ARmsIvLDwBiXeY73aTWI8b5+2c5fRPudEjBFz/VNWM
yiZIEDP4ooznVt6bIQL2/pudol40BU3hH5RA5jEXIyWvjZY8u2C0gP0BIcco2xfF
bWzrpTKBk6MzQOZ8p8UFYkm7inMpzgPcSQQzTxi1jfHFxgKVDgSmkCxp+ubN1bxl
rnRjhDdqEcmochXHTUzvm+YXp7XjI32FISk+B1sLpotYgt63Uuc91tR4MfLMc/8v
WNj8rKIekYlwDZamRMOPzuDiC8l++gWa7P0i5jtd6mA7Onl9fPOgdLrP4P2QPMXw
TWzWfbYytkKhlBXKKsy1+JAP2h07QTFWrs6GLGaMrF9Z+5ZQLuFAJY/C/qn/o4kT
13Y9OGImI6n+83UaEksE/TxxYhjjfBEdAsinGgyQULw+V9TiJmxyUPoBy0YiDyU6
YC0pQmrfxBVpppetPMNKJSDei6oaG4g1yRVupp0TXbgyx3j74TENYUVBV5WwJzRK
fXv8qM15D6vF9D0VAIF+e4e3wSvxA8DBLBLPTmk0oII3NACh5wwj6MeLnIvuvLTQ
2AbQgxMkIO1TCvr3Xmdt2Q+0bQ1inMzzLWyBO2DEwXmgh2Bww64Mr8No87h9JP+k
lLexyp05WDCuOOeUK8fb/jZBmvrVkaGbw+PmPDSKZo46DZ7Sd2TzAdeVeKypRZOB
NGY1F+2prWKjw6koi2NkKX/w6vjhWaB/QHaCvxGKlj2HAnpEh3FZ6NErDnLVNVbC
efyWtUavg2Om80NovFqQuR4qLcqYwYVuGR75maCqcT9qJAVTcEXsulRa65iYfqqD
ryvD+ek5ptcS4ylUgeU3n/22w5ibylleAt7FT5V7JuH7vto/THBybmObKrwwFSnI
kCafCSQtH8OPmZwZPO2Pu4lSUtTJhHMAuXgUYpgbBf52zhCpIsWc8zMwSsQQRZ5T
eSa4KL//WBLqzAYV4QMF7O1vSdHSmlrDpdBeu0wnr6X4uxwG9ChGvQFNbuzcCGkj
Wg2zGiPMyZuTyCSU/nkYdQG05WP0nj8QD5QPKe7oIgnumPIr1ZXFufupAr6fQTfz
zTO9bQGvceWeYW9YVsderl5ES5rrUbiZd+FIi8VflBXSCNA09FooZlpKQUhS9NWd
OczsFfKKTTlJln8C9cbBgBl9qidVcmXQ0Ns4T6WX3AF6VqSu47jKXbpOKvie6Wq2
LDY1nwM3OyqQ+Kjs3YQw8HtlDnGogW7+3I0ArorIBt3qJhk2AuHhtOv+aXK4pbop
2W+7DvAEzISI73bYaJsdMvSzZXc3MP7o9lR4x9YCo8KyeOzDesZiYyqsPjkYF80O
NX2mQU/NL/kNk6Vsf/MvtecnmFlp76ukxQbVdnsr5k8aANu0rPYjYgs0L3OAjNsZ
4ETA5nb4denMWyJriRB1nxaJzRy0/Nu7Pu+pbNJf3k0Mw8fk9sdFa0DcPntcVJAq
5Q9urhnQHgbB6N1A60++DG5x3/RDaRjoOjixbCd/9PSyVcHHxZO+Ro1auIBUB5i4
rtPmbPUX6ei9y8ECtKMM6zbTYsdmdxmT6o1dwNAyTIHYoZTnInRy+Z9wcVTP5ZmF
Vf31VsM6l2QjU1UwSD+L8t/pum/qkgZ45rRu9UEnEPzjjHqr96ZB494RwkBGX8eu
UdI6y2vxClQx+4GlXlnYcQOqzM57NWHviLrXLqWhIDK9HBr75qXZTfWvjHh+f4AP
RYm/pblwGbbz8LEWonCTF2EhPjtcJtZjWEzztYx1y7GKR3UbCwB5kQNeebqxQwjd
YcqgiNW/dRSSFQKxsQjQEwcAchbl6F+05woV/fPO+AFS7HdX51rUzKvO1Hd7tmN5
ppEoqCEnh35UV1Ktqo9/RN3E0WOsYMeftKAA9eS1kgOOqQHbBnUYdmTQR34M6U8L
D0gSm6SxBnC16iZejcQulmsNdYxIRO5gR3VYHS9wbMpX6vtYUdYv7dlTZ/U56IVL
mUgz9JHhGbtBRegLdPvnFm7ph3KB10zwW+gdMZTci7qkFDvqAbdziPu/jaYlFDQU
GGnTPvL8tk2J1XwYNKHlS78IC7GjmECUncuoWGqZvkgx2BrpxOpFkCdMDJQyHef7
1NnXoJkdf3XN6DDbFt/onzoF0w6u1TGAu9dLCZZpDeHrpT7+qYYHgZGpiVYkT0JG
nEFd2Aci0B/0VACHrMq/fgkNUwEpgJSoqTgTjY1FFBUX/4fvbizz0n/JPVjINE8m
CU/TOE7Iia0+Bvr76OoE126idBzw4FaX3cyOchMq028Ql+94fUZjj6ZLX+3mcrvw
VFK8udIvykL6JBc7vyOJwIISIjZVxWDr7oJxW30EkNzp2DpmHjXC6OhRWAQYC1PU
ZN6kGf5ldHlmP5TLkVp4V2W19T6LjI7OPLrVGbZ8j7q/FCLRnfmvLZLiVHaPMrc4
Xx4lX4bMaKw4eKz+wasuoQf1YxNOuHHZlkvFB6ToPnZW5I0WkG4ymyGiIAHHRXBs
98rzYciQb7WE4dWctf2mm5Hj2fA10HvIS4QPvnS7csHW1QFB4MGwEvhzpGxPrvxn
8i1dmY4763qgbNodVg1pFpkWLjdM3KH/d4BEaQm91ECxGzu3dCqUiPmfOJZVonKI
GSH2QCKpbysJEuob5v4oS2buLks/jgTkdx6vrM1Nwp7eHujzMwPDkT30ixS9NJEr
AoM1QLr0dJ1XdkEtcRoeVGVoBY8DEWsyGf032CLufRjcQmLZ1aYuH1aoniAhF3Dd
XJ2kI6DAkF1UP/SFpbQg++Nc83Uy8w/cE/6hrlUnESKGpZDcXclGOV/ZM7usFxUD
SMXX9B+GrhYjnBrQSuWrKCpxqmFw3dF3zQTBeYiru9ikDN99Bz7UJJXS7xCa5pL9
MGJRH92LWIuUUU/40RinXzP88G8i99vWFVO4szFndirEJpgYue4MLCJpD5mGZlIR
BLZNkdvr5chghWlGMggOmANizWUoU5VPHqZh1neGPmKm6RBkjsTsv/CnGwnEEren
I9eyx/M6cte31c1UBPKVeEqJ6Vq4qhnC30r0SLF+yc3KV06V7g8Y5+wOQZn/9Kl3
AfmaJHo0pTDiogSAGFGnEN2qoDS+XcT6W50sIe/crwCouk8bC6XXwp3R0tbcPPHs
0/B3K0c1h+ogxL1jQDAU5ch6GMNvXaoWPuLUmMcsJePIPewS1tm6xlDVc9bAhQoH
W4HOp/W9bZ+lxiVqzx61PP+Lom6c1sAbi1sj8vlStEhBcMgKBK5Qz1TztQZqBlV4
shUO2rrsnNhutiULEMi+PaTZtc4lkH6+TQzS0udQQgMiNs1Priza8QgdcTdTpISj
3henXKF/mrsFCsz8mDrsBAWTwr24I64MMKcmtXmr0oIdTdD4YO0yR4rdWsOaZH0s
rHNM4GD65Sks22N8WBh/xfIxlhl5oahxdnzfOuwQ17ucDSABuwTiF9ZBSb59JHgC
qkC/dYFbbGJaE1y3E7pE8RvplVKQBLAOdOJqiZHV2EfTLh8DePyVUXp1eilfmwIx
MKjoj1yXrrScozb31VxZA4KExKeHR6smFNHfyW9MKwtTwsT+YlETaAHPfXeZ6V0T
gYh8M5oFfjMiKVk+ojvvl5rktCep/knz74PJfz28Ba5QAzQHXxBHEMenaRJikKS+
iZZVTuJqmLkPZl3hFu6qLAkKy/roPomA9OKFSuDyAGXIrBHekqi9nrBHrj4p2HFd
iHOkv9HPyZREmp5sLSayu8k1xzUImxijj6Dyxfq5dd9sUNg75mD7e0jGjGHH+DkP
uf6Pn8dpYoVB4OO7jSVxZwr5B4N8OcIo52K1F8hZPylgWqGyTb1/3x6smsC0MJHQ
3501dZd5NsKI873bEfliD5sYi8YDeJ7FlvP0YKhLIJw7XIzkxl2xX02b+sEULhMg
055pZRvFEd4CwpamySi1RS9KJZ9/IHz8dS8Ir9YmBCAJonazIPph1RrrnGJAOhnr
TuShtuXUdfBTRLf7CNJwZztzfYytQ7pGEz9NkDPvCoOvSJBIsuE8SDgZIBGnm6Un
PpK+NWSLNWI+tsDVYto0HrEroPCt5IkPBtacHC/KkKc0GA/WfdmR6Mp++5S+dBhV
xBUF3FOJswFYsH5JY75hSdsMjqgZypR1zKdvb5f+IJkhyDmIMtSIlJclZQONghfy
Z1xfRTjhQFqXHnS/9wkH7CYaLudBQfJccjvJyKMwxFr/xTfN7qMBjHhmcAU/cdh4
4B9jW2YQrZAuQEB3EJkzZyaQm0+afvYvxJdJ87AeD7higE5cEKTiYFMFwKgAMpo0
bzhpWPLC3u7e2na2hpUJQahfb59YCYfvoXZcILfpP+psImKwBS+RfDiuJSZMzWhf
dbsaNdloWcclp3aP5HIJnX4dLy7xRx75E5yRmZUOh7yGvYTmtvl5zzFt9Ah7YFmO
JPyOHzkRm9Cbyr0OnieCf4MpVO9lvl2YVhT9fo22op4i/ThkhoF72vmJGK4m0gN6
uySjvQBQnImMAGozyAi8p6a+antM4ExzdomqFTRQRR2w0YJVHpcpaTKv37bMXlFJ
w/onGcossY+fejTYBb7QIHzN8MbukIjwyEoRbAO31JsJg0G0m96NBKWgrL+c3BLJ
ZdQZ81dxT8X9oFehDQu64qh50/Ram2FtsLp6/w3cx0sTFEkBFhV54wFyVbGg9qgq
iT3phnYWAq6AdA8QE0MWskvGkchMKZQBHNrAxRGEfG12hPzA6YPTaM+SJDjsmMhE
IZ1JhyYzrgW8QP6xS1YJHU1Yv9fHoloF7xXHdLgIBis6NeOr/dTs4m9Wl6p32ZPK
s5xlNrkgMwKmIYnj/MXaTIRtOa9BtB4UQrMea5fOmKzl0rXBGQT57HViXyr12Y0x
lGtZWnUgLCUdcDzROKi6/3sgO9Ff6B5KkXJDJVGSvlqvIkDeAsYkVi/z1Boyecbp
0DC6yKYj6TuZdDJBU/lZMtfMdEc+JG6GKuIH6KtMfwVg5dz9cPMMS6uP2/FC9o7q
5sMCFrGDsm6pSZXkj97ftSe4tEWjvw7aBNu+f/rT6s0CEYyWqoBWEADumUfmOrLJ
Q98ZFvUluNduRpFZgeHOEaSsTw4xDKVNVXZstPsAhmEL0+du+Zk0kpeoxBdgIB9i
8Se/MxiCFoyQx3BRDNSiD614pRfmQSTjlMDiEgT3OyLa54fpp/5aAv2QI1hQoXJY
pMShr0HMCMJN3TKMioWmj43Pm2jcrPvsFAK7CwQIrlDd/sv/BZS6Dxi1g/FMpP6b
SEMC7TcWZBhyPTrIj4P//R2kqFVN1u9MaFAWfCahdWeHX1pThfkmKdPvL1vrCLGv
HIOPMZKQV5mm8HOL2AEzoNVirYA5vKgvKZMsW1X/Jrd5E/EsY47JTj68Qhq9MOwY
LZZXZpZOcJCziB15AF8olMoMiJ0WeKtvT01JOmVbKnGyWtYJBg+PXza4K31CmWGQ
tW9bJiSXAYAWyy9X7bLS+Oofl5A25SF+dFny1/Aw+R4w0oSOISDcGIbHUmm40PVF
JECxaYwHcna8eav1Eebaq4vQck1YHbf4C9b4CWSl72fOBgCMTbg8nWOfXrS2DVfi
9Yk2k8T2YMe3rZztPDOnwFNWT7rbbRP2Gw+/sOTr5d3x096Wmn9uR6VLeT1VUlZ9
NHxYLu8jygNS3Uq3g1DE6zZKvavGjwbJChglwVhHINL+kU96EzDmUvaWrvHGUYEY
+uwNL+lzsv5WSb0hn/J8/1PFverS+eESgE1mC9t50qlbNTnPnakdhRtUZLSrYfn9
n1tQAntFqO5PgwLkWV7+fqRaowduWgtVs+ctyBLzAsYS99oP00wPDy3zGcm+PCws
ARtbcqtzmo9Qe7eDlpvvt5YnhghTRXGzcYWaRceTRUKNzxsmoDBW7mk4yYdCFq61
pwB72Vhie/yAH+S8L+l/uJSjxAPAM2EGWUGWDPCV8oBeztmzCpR4fYcNdhloDjpt
u93HpQkQGloND7Wctleg+nPVsWn4TSJD5h+vSxg7gAyia+/AV81/X6yZZbQ4ipcR
yEDSmxBP+b5T0qC6lYApbCpi8c0Ut0f/FSZSlQ0hImK7ntFG4+PDXEaBMmDy2aDm
rZIwsGffVyaDoE3V7/dSle4uY6SFMllLn0qJnE7cHLmCg8yqYQWCFCdn9k6nER9x
K1iQunO7dxGcb36cBCKQSrI+eNWwL9TU42Ee5FM+rrR8F/SYcNTRJtKeK5jZrE8b
Q1QkiVDbr8IL6JsO8HtUXJy18TiHfOP90E0Rtd0/qqnQ/9koJpJZFs3vcweUuDwH
o28tw+2U3+ue1X9M1os3wxchJw5RQMVviOGSx4+U6jgu/vLhM7yfpRlj9JehCYHF
MIUlZ4XzhWGBVRaMtk4ASquhZOyogOzjWqbsd2sn7ErEIm97DLD6TOUU4uxgL/v/
RiGHRBitaDxmJ726cWaxUKClOSfE3QGOLbbE9n8FQ/l3dbxzeoMdWPiifaJKmWOO
smxlV60R3Fvyyl1ct7nf6Ydp7l4ZGw2DrS9BXivPUNq7T8mOp98DV/y9vowEAu9/
4j4GU/TemnbplthZb48CwyaXKvq/96bsN/vL84WNV2qVt8f9+x+KU9vRzgsBWcB0
xLRHX6AWu+JM6bKXXXW+UeHeQdxMgi5qETYzZmbjIXkrfY1NCKHguc9AvhxCCEBp
PUXSlsH8Q/wt6YG8KCDCumN21qhV+Zc16R5BGfRuzcW9/C/INJ7BYOV9F6nkKlg6
Alj3fKRenQo8yeNEgctNTeTaQ9C7j7UxEll0W/8eITaddSY9yjbhZjf4Bhd2GVHn
SODhPzGxPqkuv5bCVA0i1NM8MtsrP6GwC7HIjOtqdIRIBmdQj6fPl0RZPOvPBMQI
Bw4H7K/DTQSnrg/RVJYDNuzCVJo4FOQ8V9vzS8b74T+RzPGWZx4m84EpSwxMUCeO
fhklF8TYBb3tUBijOw1hB82PNkxPkp+skJUbKIIcEw/JcUHyztJ+BPu8E6hR8Jhf
b3RNzx084jLRjZc3hNOlDho4ARlmKSVq7VGtAQkanuAixXRqGKqriLRAHDSoFUGX
QvBFLlWrY+J+x8epDNlyogXW3zwSAgLL/jDMx7QA/IH3E8FItYgzSohEZyXv5EZa
0DryonuCmjG04S3MJOHK8rz1AcqA7ncLAbCTio1tN5EbCXRTDnoqEmzHtemXeefB
+nyX1tOk2ht6SqVuUiWZ/q4KpDCJnsKxUYORQduxThaWvmLyWgPZfe0y6kqCEHUa
nvS4hJ29sfKQ/BU6764tA9Mr9D2gvndC9cba7tz9w548jPuHTzaGkaDv6meNtoaE
C6RmWBWFQAe6EasPWXqRn1T8YKi+8PIvZrbfWsRd6p2waMcd/8ILfYGsiyUAu8na
XIHyGTgnMBhQr400zpqDRnlVkUWlWDwoW6GbP/SRgnj8Vpb9yOQnhg7A6OwtIcg0
DvjQplWp98Zn5Io9o8WAuqxClxExG2695ogUp0mBLYrr+0rT2eW5fieckdKargj/
068gn2l92OpupVna+5S7wRd86dkJKuzHv3z1b/H2EGEn9T895/VeRetSFZnc4ZVQ
M0h8Ku3l02IESeXZxwpoK8dx20i6m3rGmxF/efTWUL5Sk/MMi6VDse6gZqgKy1ff
BPn8AqQOwfvs4SjReaR1zyUWDUdMoF9PVCfWRmW1mIt2KDzW5JYMUUgT5Eqi4Gu1
73kK+tUsg7qsIAIpSbDavXzq7FsbrvKyHWUs5F4pAHArSONzBt5RF4K5D3bScbBU
egBx5CvEF/KnWSoNJEO6SDirSrHDbLf93G9IcLf9mfZqVaf+ZxWcjIeIhZZUgA0K
PclWlKUojgVjAyLu8Esu2Jx7JtsEYTh5R0NNRX6AKbh/9PWUSrIh/JkD5Pnu8lVy
w8iOTWK3QjWR5hrKfNu4YGtAZcXfJbDZqYRA6rCJ+Iv05RfuOZJAn8PL75aDMcNU
8FmARKTPeq0Qtn4supp2ICZ4e+D20wAkRwZ/JWdxTX6/hmTxkv7T5GcHmPvNOm1k
jmf3DzFKKYkzqjj5Zww8lWizVikFBj35J7wood9fMjS2lqy5kb4MovAnxtZbg1VN
BGBa8bZ/fVuxJKgB6z3Pcvs0Py2dOqcHnT58PlN0n6B5m0fSj6S25BS0KXLNQ1Lv
0J2gTI0P+8AqA23gIGq6zxP8bLuvHfiM8oUmfDgpKxLvLxCK0dh/WqQUgFUuImk8
ycmSp8lrUecmGvmEW5PvXj4Km5mxH81TIjGKsk2DpGDIBKI2MRSAjuFGEceot8G4
baF2IRTVE7qCJUIuJnqSkPThpGIe/6iyJyJDmN+gzR1x7OS648o7Kx8UTkXb+luJ
5o1LatxTgRvY8icAFDUhQ9u8XZcclwTbOW2UWIacfdDQfW9uppdR+QLkwsTiG8j2
nEZxSx2hU4tHBmw1XgTEagaLfvhU1jO/4SGzS1zasv0uuZDH4ww8/K4ptvklhiRv
KoTlrA6ud8MXGyhfz9yeAPY1zOQ2/WkMhJ9hSQP/uNCj1o+MUtgi1GIMU+Dxabxz
7ahRseMDIZ561MLKcI7TyOsgHrlcv3Abv6qpnX90zbOHnlT0QOIFP/N1EEvW0S30
vdM4x8uzjXkUQZ9IJVh+7rxz2xPuFgHFsWhfwrtg6A/aW9nNLf79qA2p2v5zhbJE
2rcEQfPulFucRhbf0jlMexA2PueXEvQb2FS8x+WqSWP/0dXWJKXzRw/fYbzkr7ve
tsrsStA2aRHdQ67dhaFCmRApLHE9l3ycZbz19qFTDHN9cMrlqFXoX+U4MIYwG1ta
Zmwf4JbpCZF7ia5ljjVjmpcPLF6hSuUuECjzzxarAIiDog1LiL1pXvU0roFghV9U
XVIzxGhi7jqxNUqD7jyal9QKH29u91d+d9hdWab6lGpl3gs67w08WJyWKAt91/Cf
eEFWBx31WGcztV7GuY03horuBDiHZ18xKM8BevMSIox/FU77QNFITbE2Y0TTor1R
dl4f82Z8WNa0u+QIY04Z+U+B7ypvbsNsPiXQ0a0HoyP8UhHHMKvDJAJqAntiYJPX
OPZeczPS9bNs3e4I47tR9WDQZi2Ge/l1MUUPKp4nnaU+W5hJkTKdsbQpb0TRnPSm
uOvCq6cM1LLfB0O+KwUDUQyXA4w0c/uOpMR/dWjXNQ6tYtAlgSlb5ea0fYm1ybpw
s8M75gUgXAGNdDoufVkHxKixoh1+04yyNpMRBdw/okeyz8pSTeqoYHgbQ1xhb4M/
NxUzD0oKjlHHH01iuLCcYqxLFiX9qDz6WmbAGqZ2OGRnwnUXZutjzcDJEmaGGqNv
ybK3Xz8e3C/OvETEGvEd1hTifWFRnodfBuyDYWoN7+iFUSrgcNeLM/6T4g4+xQb2
j8cbR7cLzhE7xmQOKO2ejtdso4+OIzQutC4VbmtUfdCCi10upp0NLQLZ5nUurmss
A7FqxdKRxG9zKjfR0NYUNIDHjtbpw24ZZFq6rDSB+WE05MGGnzjAj8+y+fR6qLlW
8dN+P23XMD2+4u0IKZGxNMkp99LYjWzdpi9Ifr9ZMS3pJ3S6mPcbuUV9hLObqRIl
pldimTo3I/HEIEOkvNyW56AInIByeyA+m/JQbPSZG9IoUS0Vl2m0TZme0ZotpKQb
U3siyemTK3rl3lsmHq1mCiw+IJy1MJxjNQcRi0YjYE1cEdTKi6mdhLrTFJ2XQV6Y
T0wRM9j4xHuSAmbyuZ71yX1PF2kBbeEUi7/VyPVzcrDJA0IkYII6EmJ19OY2M9KL
eqQr99StOijDL7LV+JX8AqkgImZHyICbMWlfZH3hpRLmJzYafqffW3uYyS8XsIf2
Ty2gE8p2a+n5H+7rDxfLf/3ZkExkYsH2mCv3TPlntY/gPOHHxgnLBeWQPBvvty3F
5gpIdeVY+J+UVFw2pYWx7JWWnfEIWPHKSfq13azSnRoiW91yMg1MYdVPrKyNvpal
/X7AKihedAYzmOLX6Hgpxg1dp7QVgGFHbnAEELHTO4facS9qZSyOJtlTgy8Xgx7/
eCYAa8aIqeFuAhvgL7cXg2tTN1GFDeMtehoynZj2elUoCXogGsqkPBSzXTAQRyf8
pz4knRNi/NhqnDg6XtYY8fv3wTtemAzxrEYmJYhl7/vlbAVbCuDWVPnpRz00wyq3
HtAtMpW6546ZKaI6UMr7el8p87dC23fibpc/C68eZihVVue07h3rhSvxKVmLybEq
J/dsrvNmbpPGCmNihcVpEhg/UL3VEo2LY5eb+oZsq1e0GxTvr7VcH1ukIhh9NavI
zEC2JTqjapWgNXe8W6rvV6HXv4zcmZa7cmJWyeh2H/YPPy9ZUsWyXx6pzqZElOME
x7QjhgEh6AlMRSOPg5+zFhfgNMbjEO1S3fXf3YEDMj2kvCi0N08a3YzG5gqi7AAm
VUoZn3afVeqeHcrHnfoHzbCR1/4UZWJDbU1GaOb0wuwPFVS8796xE4rbR9zq2hrf
35ROOCLJyjPmNh/b5CnTphaOo/U2AqPni5FJZrWuvQjyhd1vr0JG+pTqNINtDKBz
5/cmaVsxwO4hBAYpADyBja+vmUGGbYUnbjGWcnNM4yGscMN9QU/eWMftr4sKAZcu
cChFhjwjX1H9JwM/XJZSnYy5P1q3WOvxGDjl5xvf0Yo/oJ8jrlcKv0tbvBjnrZ8o
xqFkh+er499L2Z4xEMJm058I8F4CnFGK6hGm94tAYUJU762XKC5AqKpm6xP4bk9g
gIOkQ5Z+kmxY5VCYkNacnVRwIsMCX1mtGDDa5TsHQdn+1xIXeD41PNbgtddkjJyw
y7Hm6ngjueY3jD4/IRrUKZpX4286T7m3t9ID5Qh6gn1eYKvWAHVgYlmsOeKyqxVK
QRXt/KUN2vQvvDeDijdymlKy2VBFgNcg8NRNXRUnhxGfescvRJ4xshfdDWRsuI7g
Xm8/ESv6wUXnF3N+wANzQHWC95UAGdf+telJYdGPzc5iJNAPF9y5KxlTWchjP4lq
qI/vGeuFOWUnE2tTVZZGUh216hXKZO0SLIOVEK+uOxFWO2kaG+I1G1WoGQk1eOD5
Q0KfYB4+MPzJv30lIqGzUg7SYeri+6iXKSfnDYcs08XZF3EbMiNnVEFjFIlf2Idd
Jq8c+0gm+D/pkzUrbSeV+bBvoejRsvmgVBkBUybf+pj/Mm+doLAfHMEIbeunBz3S
xWqFk/E0AJKNfZnKdXQ6DQEGz/KKwMXp/mDhnQ6S0bCfH5smrdT3IWVkg8BHO46I
4HIxx21nW0CFyDPfwTqAYMA5V+cmHTXbHrkxMVPw9i0sZ8D1kjysInd2p72pSDNY
xqDzaCRCEb9LBxug2AooVI3zKup46g7BmHkrxNV3eL8Jy8Mr51FUzGnWzfnIU6Zi
N7DPhzZCs4L+IrS6BsOpZuqGt5jBIyZ1y5/Kvp4WGjNH+aSPCuWcAqR/o1S+heEx
lWD3fjSEU0QpLXgezkMG9isrBADZsX+dgdMnsVUFJHKcFggvUPAuadXLTQsSZUwJ
WiTOj5STv5rG2F7eHV1eaxO+V5XO7LhxC7HFwNWqzxnZVJCSJ1XZQWKRmGjAw1bH
IQW6ostc8KFY+2IaThkd0OCyASRLY4ztE7unYP2dKJI3LUaX0A9AF1NYND1Ypl2V
RmExR+eZsNAnnl9JCn9U/iNFuH54WqhK+KDGbGKogW8byXJd6fhBGBcf8FPmuEIw
FRQOeVhjMZ9qgXKUulhuJ6J1NmwbtErwKOzhhj99ZpLCbuMcuddBoCgPXb8+zJHa
QsVf7fiaDaQ9ASDpwN4KYiQ0yUiO/P2BuT2CMC5/kKQUwGwfvVK3wk9CboT4u0KQ
qBpwfMQ9K1vZS/cRCPbKYbbzPnI+HvcXbvb41YCbDXdTxTbJlyIVqB2MOQ76X7Gn
EJShx031Sz1pWhwng8ox7GbIqDEh+7PqP1K6wBoHi9Y0JsixlG2w3uCF+ykRlYAt
xz36bw6SP+IPz/vw4ce7lp5DGZ6EE83dZ+OvQyGIrbJHP0gYhB2tB3fiEykKKBUy
ojawm8vHMpWz6VApOJgbDQQmvGTlcVqoY8zRXCzJU01WuQQQJPIk0EgYITbhZuy/
n2naYdTEXreyGIC6RFZYUSKHFSt9C5azqdtfZHzMTQ1GPBaumHNsfF5meSlD9omS
hdb+xs95YdiofID4U8H8F5JYd3svF+cxB9/jBHRDHuIElNQlwpBes/PbNAEeIoUI
JzNZSSEqe1uPRPAKLsiZeg9FYvoKx1W9yUcvG596RoikVlIfRL+Q1jDJBqgflDn3
gy4ahTaQdCgozGGW/Hzo4cw07MD75wY2HwwbA8PG0BSypRHfjJtZ+H9ExFDKqZuF
ZIONw1oNbZHJqAggp3uajJA3z0Xu2+s0HhAfk6GgVmZ2SMBwcCVnQPjYz9R5Xkz+
1PVNAGMzIMEyN8ZIj6TqlCKpHDIGjeb14HAOlGmF4Y9k/BhSGBUCnpuhf1Vi5anb
qKlBr5JLyA6PV/oRjaj6fG4BE59dBZeXTM1FVpxxmI3htVQQsBLYes7jVfoZd7N6
hZr2LVILyCIRvuIKRBmC0JtFKWTghBdhbfLKNP8DiLxhkou6Uv+DEyHUB86wD+0T
55RcONiaz4CkYwGfR/y1QHuG3t2lidsObEdPRWwjB5NUtGTpkp2Q3iH1R+SP5zLx
sq/s+htXcdbeqUwzTlT1u+EKoNTssnzOZPwzHrySfOn/IfX+VIGAuAzWR5H5SBiU
NuR88AREf5++ucn0w6cCfGmQjr3ChxyXy3Mga5MyJvQQERE/uQppq6cIZQOVNLXX
HgVz6vql2Pqs6CST4AovY701wBTQblTLKtjzTZ53DrTGH+rylp79dcjbDv2UaWaG
ClfTmdfGo1hxnvlLEisw47fFfLgPcCMew62YaIL/7tdgn71eui3XwF+6Vb+FhWTM
GB5Ms/yqReqjfTv5OUdp2TTZd/SSQXgvB1gbWD+fjjtopKk4Ep6ovGCs2+Xo9JFY
UqfG9AGgv0l+UBECMMkgP/k/fDGKsJAF0wg6URLlB10Oqc4516j7aD6mbnpQv9i3
JRTxN8a+UmLiXCGsof9A2MrP4Mml1ju8LdXZzadtx1ssf+E4DbSwAEogKMorny1n
W7lGxHNTgUP0vTdnQd3PaUT+SEkoi2p2Rasawzu9iAEMVkzbt285k9mf5FqWj1yV
A9vgt5m69sDDfHCfuBriXiSaKUaEdls0pB+y7oO31DNkiPqMhzoQ9bzNMeUdtzTb
TxYU9nmtQkEdDMHbX2ULhJ3MlC3GbGuQ1vzu7uiG2caGnRqHVI8ABzcskqKzMYTu
FDBt1+n9/D/6UzcR0FtQU/Slzka81wyUYSKvK194ke32PUr2ZGC6LkZywHg06ldg
/sKvwaRrDJTAcUYNAWWlHjW7vUDWTOb2wFCJW0dcq8suMWTi1nk23Mj0fNfkRyYX
7sji7qxU44fEY+GUYGHOwiL2gqbJUOUnyeWqiCe/DXPgVKUOTUY3ZO11HUpqvJOC
rtJjY3mssj+1FVXMNzg9xK9YccCgreJraCjD8g/mUMEVSmMnCz7+QPYzBcQmYdRb
y09GV5N1fQ9zBpqLew5D3Odyeg0XKnYQK5vi513OiITuGam7HpgHALUXcR97rPV9
e2ik69vkblwwb79R8qpHWA5n597t4RJoSShP7oKOIfyznC2R4KDSd0DwnFoqUaom
R7QdD2Vlbid4PSX8ESNzWLa/O10NdqmWx8ZdwJhSGesEToROHdGVHt+TkxJCznmH
RYTvPmmkcQmT7Ufd5mCSLD4WYRP1g+3Y4rtTp1zqQti/d8Yh0BsK4DQRmjmrupF+
3+5YwIFmtIZCOtZ3ez+UOHgFpS18DqF26G4JceDadbBaYCYZ4AS0iHO7NCtpyHKj
QLWhNQxPJoqfQj0yMlM2TYhuqRlWvF42T/+EiRDG7T8/Wd/1xITRF/rY2gJKag9X
tfrfBUGRlQhI9COjgWVPkRWcr2n9KhB6+BE28alc8lTFqxy0hgukL0N9hzNktQVZ
aSCCS93eeqoDtBwKdXPht1gyf3041oSWRtGx35R1mlBPmDnX8q8pB1szYrbQaauG
h8W2cY7JoQmFX2LY4q/T6z788+Ctt2T36lkjV3xG8UquZXpl8f9fw6Uj++pD5qEj
S+fBpXBIYUoBx21Z4/nD7K28Kik6cl37Zd6cp0VSsYCAvKJ0tOlztl68GB+0kUoA
0Pps9lnrdxY6+N4iDUBgfn/fulraHvpYjZncC/6/VePNtZ97Tqy32bd3CxlvnLAP
RBZITl7o+wahJn1WzD+BTQghSClkjSUrz/xjxZhYIGu6xFenIRduyZTRtvO/SVl0
Z0dWpgYk+0aNSejGQgCwojMplNgl3RP1Gdjm7FpdwF1rSBFzmyQo34uKi+APSrN6
zjzI4lWMyBXyum9rVZFk/p0kWo9LLbIgmrdcqQMxeHGtwbVVlGuc2UX/Suzjdjz5
SldfW0TihuY0V9Wlu3oRIrXxZJDnvsSxcjlGBZFE4l09Nr7iIarXGJ5IsdA2EAn2
Sc3W5ILzhNhe32CkToE0/9RDbAJH/yMG4Qa7YaU4n0gPc4QY395to8IFR3CLcKCp
N/89+QiIXqR+T0RVqCYRIC13uMQBCoWbZWsNHF+1vZGLvAh6fdqhvz4kMYJwTKcb
7FEygWqBvhVwMVBYdD843X63C52mHCd1/vY/xh0i6E/oz/bDauhv2Na74jOzEQDK
nL3Bk+Z55C026Ayqipv1we2TkQpXHxoJmDn3hupkQt6r5sIhVpMyZ1jVfJbB8o/g
Dwu7d0L01X/vceQCz7xwYvGDh8eYdsfes9ZKVp6uXBC3STEcjJbxpNHOQDIMra0b
CLv/6wtAFssi0lpdMjSzNCpIF1SMi3+VHl6Y12yblYv1v9yzX286EzG3kAe3p9uN
rts2ew9V/YAiDF7DSX5t7nbt345MUE/dqWv9ORoOCRuUJ1C0JfXZbq4GLMpl9RSr
v3dFoO9FuqRVOBM5xtrv+0oBorRgKV4A5HQQ4uWa/vx1SauBCFAAnH/T4q3WgtRA
EiyR2WuxaL5Zhu6eMzaHH4cUSo7hf+hhGcnDy7eCSrx3LDlK/8NAKZtBPgIv5Pwo
fMlL/nrf1htf+qNfhI6NDAZdzK6QidnIztkN+4X3NNFgmW17aPsRSa/IfINXD7Wf
kj+hlp2n7K8RXoazlSOtYzleQzFWzme0ZBHplJL63GcXTC2KMDO40KmBLd3hlxxi
ZOaHrhq3UTWheMYzFnaSSJqOBpp08l71ZKwiCSUe7ZJdpsCto7sw/VThGMFfYQPm
UAonQOg/Sd2pb0FPTTKInGYiDJL3DG1iVac0rI340MQHro+F4v/jabmfWjxAyoPL
e3lfD8TPoN8zJAsfx0PK08mighHNYp/ui15fy6a5PiJyq8kG2dFuc/EqglY+3QgU
20U9MfPWamqEHLQH6OBneWQPytLPDn9+gvHiOK+jgmcNVNrXkYdbflvlvGAjfKy2
MYw8noCOOReV06R9fXmGYKe0mM0A57pCkBI4cdC8raVeGBngOO8Q8pbfeXI/tiVa
rERobqJwLyYzVENeUc5p1Vk5+TbQnAfGblFq92vHY5ZyekgzDklsW7g3rUJkJpHA
j0AqhutDbthURRY8f3UEjVCTfNd0DYwM/3Zyb4RtOE3zYvczFAgAu9/gdnQudRtG
ty9BJ7vNJHLaVkLQpAKVe63Kuf1hB9O/AXpeFR+IgrAc42QdnQT3SsxaHpApiwc+
KrFjY9nKC70JUFH3JHTklxO5b9i8QPcP2E5TdwKnI0EIMHYBTG0INTfJhHZ2NXD0
14Q6wWVPAulUT0l9i6gSLdYB8LWl94CQ0EbTf69yWz4TPfTf7kbzT9iUsbne8Yp6
445AJZmV9Ly7aj81yUaALtQhbYBYHOCiUOdiueZDKf9u6LogDz/ESRkNwB7WHxZC
FXiziO9lsAFyeQdjZ8vkZZ1V78x8KB9GqXAQM9s0Spoc8nh8OL3emfOzNzrykjpT
rIZNdGsrA59Ep+Bf2fVaVVyqREKjuhr7HEKNwxnhpvNMNJaMZ4aHTaKlZxq3f954
97qUMR9ZiT0AKPqBsKbe8RdDwAlNhmBP1eSjOg5BcMujjPcrVk080xiqJsR0Rexg
dPfrVqFACYtOcJ3a63nrD6CHVPU9o+wWuhzQAIhCQKmoEKc7SyObqSXe1+PKIDgh
BUuN4sXyB4J7VxfmsMpiGnu4yuDBi8h1Q8oxyKZhpnjj2YWKseBGCqz8hYYQSHWe
XCQoon90/eqL1Wp+NChaWruCZddALz58/B2uGomQxifhN84D/Cs/AUIIDpX3kLPp
klitTSqu9npoM65rQr2SohNKGOfls7dCZtBRVrf84Bour3TB0kWOOZFmBXKp+gPd
oJHffiD02bPaAoB9Y3BnVoG6WcDKxh6Ns1D2R0h0jOaNLCTSec4RICTR6VhNKCuO
f536jZQ/4Lp8DYKNjWo4I1bsf6tlQ82iX55sN3fMYtC+XgEHvDyuLcMBTXDyjqsx
4hPQUG3gpyI0QNqKVc0RR9ORJs6QxvizaLcZJ6FE3kbaowycf56UEmx5bPrvFPTq
ITmjrABfUMD96PTcEsj+LyPBxwjf7YzaEZi9mYb0G/M+NNo6eqVVsFZS3dDl7FYR
DfFxcDd828LBVw5E/GfseIaefOnckzG2jiRqS/zVohANCDqoQcmMLMvdyK3h98Lc
MN3xDcpF0GZbEOKsfa1M4XdOBXgWZRGMqfTh73BtgUaOQXkqJc1oNH8CrXtNV8A4
ivPtUm7yb02fIEgMZVxXh2tASnLHzrjQSAcfT13OqgQZPlv2kl7P1TJzsTPj3l15
0cK9KXde6RjeCTS3p/yM5wTp0WgLLjbErZBCX5AzrQGIbJos5UloXb/wZ0N8e2E/
BpnizU9l3WXXpBIz10w3iZLQlB4i/GOWQf3ESUaXH8TsupnVFdWjueZjBUJAd/TZ
kydI7Sr2m82xgL9l5RrvT9EIhk95EDZ8BOTBlww5x3CseV0G4Xd5GQSxcODD2A3g
6hS7ibmG5ylme7QQeOCaXLjd1vwDs8ep0Byqfuce1E0xCT3JOQtkG4bxexVGwaO2
mNMRk3XRsbH2ShQKLuH5vv8bAOXxkvvHJJLJgqQwpuGEHmC4JN9kGLCj7PQrbcLy
QNpv0rn7R6F7PdlTigoTj8Oo9o/GRIRbYRNGRKr8yDcfw/Jy+BRtJgGJSA7FSTQr
JfsZnOfS8m8b1ksR2AOmCl26RUd2HvujcpcKP1viOZg4ER5tS7t0KlVGM0JyQWEK
TBUanDRzWIbAqmG7L21WIC9mEO88QVpPE1WPj6MRlVdovnKTxqKp8u0tVDmEcNKU
KdyP70xn7VTpgH8qHC5kBfoLb7nLx5j7yh3LzySy2HSCA16+ZOkOY1GD77Rrmo8j
8m1E7o9L0VrNYo8sD4e+kFWAuZySk7gEvIt/ujOoOrSV5p01CmoHQCu3XJoTTjj6
+m4rOwR4XwSVbXA9jx60HO3YGjrrxBIHYELKIjFDKBvAeBZOpYu3alnGx/oK8nD/
HAZ4jnoNwKrVid4u2v6Agl97u2utqTnHrcfFP9D50EALoldy/8PAABH5jtEP1uS1
NKeANMCEI7Wmd57CudfFKT5cl8oxO2Eq89plqP0N+aS64jvPoD8KiCWrac08lnuo
ZYjfXvaF86IQgcZNzLLSmbcV4ktQpHzEaT36yxd8OeWngKYEtKj9JLKr5K1rtW9C
z/hEw5jIRe2PgSU1YsOSaLJ6/yHsiravy5qUjSsH+JcpdqrAv9tbeTBHw5iI8yJC
dfuiu5HilXN+kVmMUG1SWUvHoSlAN4co5C8Jia23suSi2OZr2GrkQX8zPznVvYJR
BYfGrAOoWgTAjSA2/1HBiS749MGjgGLXX2rmzjSJ1+5BUdBjW8NgKkLIloGgX0HU
2UzyzrbE2FOsn6XIh5Y/nHVPDIjC50+X5rQsMks/0fONI+5MPqzWS9u0Oc2nOQkT
gYABmK3HuZiRUK91lW6fpUK0QpbBz8wGyBapBbLBkSI4pQKSf4yTL2RV9xStzjuO
86kwv2oCTkZ0DmbicBftBhhK4sZSIuCgbxFIJdyJteHcUxD8DsPKc9tQ4AtSwzy1
0tXxaOH/btf/lp3sba6woJPGhH2KfvFatXeSlrw5LSc+cCiPxrABwtqhEUxTCs6c
r62Vig5hAQ2Ut6hbroLoTN7b+qTmacszK1uLe6RCY+QuEr1ct7dgKSjm2YRCwQ6B
GLmYh4VbgFCVn7WnX6ZZqwYaYo20tkfbqL49RRqJ4ht6sXgUVJEPiIoYh/ZU0Lpx
z2gMSXaun3PIClhByVeF81JJaiUcQI89RU0Q4z/pJu6aV5EwFqDN+BFpDORUcQOV
/ffaKJPL9lU+nKFp0Ryd0+C7Rz4FAjzWT2UrFoGmgoaQoMkduZ6UMpzaQGO/hoHo
tb//ESBKyYMq27FWzPyL6bWO3n/dYC0ba3YPujT7DxQUZm2OpLwDpMzVU4yzHYrA
AIPKK/7QoiEo+KAlagf7LJX8IEsfZMfHcbpNwC/7ChArfSUzre6spb6TRzL+/71H
mEbAnu0wJzSQK9kVM9ehWs6hNwyRyTMs74HQmbdY33YYXI3qRXttIrxkdqCV8A1v
pfETXDKLS8fBXkheMGoJPkR8ca/Q8c52dqeoXU7wYg8Q4Bp2BYd5XwLuJp46ql2L
DiAhrLEccJdsLPMCar6SolUj62LXijTo1ZLXkkHTKpOaakLqyFW97oczqpSQFoU4
LEj59NG40748VifRp7WID32jXks6F0JtWwAH33kvH+3n8YmWTm4TkgFWaSp5ObHm
ydR6R7pZ5gGrW9yPQCjPBmQhWXWPZqFbEhwN7BBa0FyAiPFXUTjBd+eVPKRy1qzw
T1K9ebC1v8LqjvPtG1G9QrNa1VniMSICqswYLmWDZzViCQCwxSCc44T21rv89sGC
EHHBa4MgdhlxP26cQKRNeeAp1UBuMp7IAnATfLs/DMPL6Bhqo7zuJjByhM8LqAE6
0vjfB7RsPNWs0cmNsmkO6ZO4FnaghszViCgRzbwX3v7m7eeMu1cpGBXy2Yv6Zngm
RBVzUntjFSW/eeNXehlEfs6kE90uiKeBjxT/9Uhho/zkgq5l5nlNFXMWUbjjSkXF
6bD6I+kVCiTkL0Hbn4Hb0DxYis0FS/IYzuJfwAz7oATbEVl9KXpjn3i4XqyPzgtq
hzhT/Cfa9S4XizC41hdPnrcrDw+KPueJ6Jv0NY+AEY90/Q0kEoAwZXbvTtWQ7+SH
a8r4xmfF+ihRXSVJDqpJs8hUYyd2NZvRoeCp736+fFBAu4+1CUYYeU2eO8vxsCiy
Qq87j2YwIdiggkBbbP1C3uMgdI+toGkB13bzfyfKgdkpP2MpBxGVh7zdPtO2y1xm
AbKXPiQyYj3p3+AiBWGokBXzrhDDzhQf1bYrXPk9sIWwzsMKByjZjJgVOwPd9zWq
vAZavHoS7syshad91vv/oyd2oULxnYLNZKbdq4ow2YYFkrqSODjQ4PGmeJ00FN+Y
ifKGIbA57Oy3eeOh9aw0VqCg2yPpP2HrlVCrMo5H3YmI9j5RgDZ202ZKBQcH+As5
o3R6K7vj5abmf2+yvS7fZWZosd7A2gBDCTF5fCpE1BqfnvET09dNZuJl7jGcdN1P
CraXvDeesTjkpSmoQt4dVm1w8Q/F8P1wqcdBfc7Q5z0dqwM0qDbGhNACsiLQC76m
b8LTQqrWUXEFTHSbLsvCUDPWei0eCu9W00DEyWEdrz0ihQvGAQJu7gvoW0FlWls4
GUWg+MMN+LR4glSBFNuPivg0LdbvRQpk4PGcyonS2rGPuPKy51NF1WaJZ1dnjKPR
ZlpiQeCmqryW0AfVjBNdxAzwqJo15gkHH3XxUeINLcmTVXiIy1Xdo7VK/2aXUSfV
4+8jXuOZJmyOzUNoX3ZadAyQwHxsIkl+Trd3te7qNpzHcKfQm9cWnDo0m+vx7QnQ
AO3bGWn3vMC/wRwXOrMsYFLg7quxjDBI2eUpYEdNtJF2UhXGhEyPAmlxj9exXiE0
JPv+rb3zY1uxhUEygQudqDu4n/hiNdQyTdg3TEcvcoYuxuiP/TnSi4dqA4t5aX3J
V9Cye5DEPKYfM4uyDKnL84y34zQQB6huQRMPD0Y7DCve1n18u17UcQy5lRnmyKA/
2MR0O0IcfbSWChHhrBhE00EjEk6x0nd5Y7Kd3p+buD6FXjAElurXAN74aHNtMsUJ
5nD0xttC7XgDd8XSwO3K32JDSOy2iLG6pqJIQckEMgQseZZT6/hguBiTCJU2mwgN
OeG7poR1E2BM4DcMGzKw0aWSIsCGAz8mp9c0un7o+7k901oKsTREQ275HB1Vfkgy
HIBhgtKOPr5Cng6+5WnDUilCJR1xqJGeYEiU63jSf4SxtQp6KpcKLv0MGZc9QKd+
LGXmo/FdOpxcXQ0jsFIJy9d8orVdKMtPQ8+wXMaNe/AKvCs705MEWbTNC5pmkJ3h
2udunx2zmEZKe113feLhhiqNocYNIAY1B0KtTuOYj7J7nV9c6Uz3z6fNsUcgE/Mj
JNMq1ypZFSkKSzTln0XTaQpbjZEWu4fk1SCXgxhEHXQE8YW6kAnrZ9V3C4UUwt53
NSnCe4Ev+5ahhCv8gwRwvTIq7l+vGPABTm3PpICjRzwcXcDt3TYx/X70lRYcIA0Y
NzeSd0uB//tGHQHFpWJlAtsCc35CqGFJOKQ1Fa9tYZTh1/gnOCryEyYgTghTWFCK
iKsGq+FkbG7lycobZyU5P71b1booGbHK53YiV3RUMAzVil80DjPtj+OMVEljn2sn
OiyTi6tW2ghVKtspRdhUbehFwOjfEyK5vXmq8gABUnwMHkPQmmIJ4WL8E/0JY80a
4+0xUIQM6xiwSd9z9nyzYt/IrUhcGXReYQ4Vxlgj93XEj/iINIRD1G5tuZnI0zCJ
3ixTgGjNsBH/6SbyOt7UodJmr/0oleXBP4693f4e5HwPCZDA4QCWpn3VK7/HAAKR
ir5eeQTx7wVoAQR/HPF5bM8fRScJ0AE1aGCMQz75sSiYuHg3Y7mFU3SLdYvwRZzJ
wzb5TlcAwddOttQ+75fzXBVFNmQ8t8Fl9iVWM0oMgg5ARypNREsYW6Obv5v2RwvV
J4PRO1egj95XoyxaKAVzpQNAShvTdryFK1qq9Nn5gelSy1sU8pCAgCc7n4i9CAt/
P49RGeK85bIWhSlVSPUopaOowKuZRpPKI3H34ZxMy9Ri6gG603A5gsvO6D6X6eMK
URICiv06qXxZepvLUKLsTMNqR3CrM3Cciv7rpPjsK0Hiq8emAHoOclylW/n3TSHN
UW2+U/BVSyhp2eYEa3aerHItKryCSiCXCrAtMdtoiOBPBZFgbhwiyUJH73EF73VH
Am47h+L+md+3SP8tWblEIXjU21hf03/JZOr0vhoNEK1NTT5aOd1cMT1Sznq7oW6H
ufZUZtVwmBp3+agq5L/cPUtO6a0AGLoG/CRqnVSxv96rCxtLktEjSI22lIl6e2x/
PFFPtG1Oj7URYI1QeMWQxS509dK6AN5kOUMhwP9Db52yOX8yBIhjj10RzbQV+KkM
vB0hDbcVvOG1Xrg4rnD99MvT9VFxN8J7aYtwf+RZ1ENvThJrJ/EcF3xRXUnLr70B
gVAiMzdKSenZ5ZNHPc5S2RMhJ8p1vvcWYSb/KhPoszSBDNeMQVMUInWC7K1QuBpf
WdmsLRrYZah4IOMKwPA4WX6o2A0OHLlyeogNeQhgpQAPqxFdLFxeHTM2D5rao7mK
7gmHcsvy+yolGqlk1FRImLVRNI0VxauqGsz4dZUA42PmZfMYWjvgpWE5QaHnXq8g
GDZhQrxQ/nxgmEGi3PiB1lDo5Qqe3LGI9VCeOY7eTTDKnE6YpMEU6N+H+7SR1UeW
nVIwRaizBpx1UzUwdoChHyr4AC0ll5dzs5Kuhgjl47duY7f/62B7au/JGCjJKx48
7zipD5hcNjpqKE1YhxNdZkE8xlB1jPTYwJ4FmB9v3dEf5tkFHaXVhBGxwjiZrnWc
JDbS70TbjXG4NlQdu26NskCsekzDSFBYkqmzR85DSgcQGIU/S08MMMFJVwskeBIn
gWZHk6SjJdsZzMowBNMmT/6dnesOz1Qo9hhcmNOMJkWMszbeeQyna4VPt/b9dXqY
+JjjOf8QHAz/bixa8sWSHWIJ/O+uxrlFtq5QRCV7kb2fI8b9AcSpLCejB+9enmbK
+RRAwDlQKmyTDLcNXs0Yt/+Ne8Nhc0zBjWv9Qwkw8XOya80UKmyU/Iebq93ppPCj
lg5fJ3EJPtEmjzITAyMNpbU1hgCRDqrqbEWpcyqDOToihKS4ZzDRR8pNlednqNNV
G1uTIsMrSwosNxroD4WyVK3WCKao7k3GzDXEI3E+bIRjZEDB7xbd+0xDnNs2ZGyo
7d3ItackEsyeCDSt61eVOqorp5ThS+rWhoTAtdVSUcw5I6qLUCl+Y0RSxKLXu6wN
zg/ExljOWqvopcio98zI4VP5QAtC8YS8qnbZRGzi9BC3NjmGUvIAHgp7TcdTQbd9
6Wq6KjsFNw6Ng+pblpmsXZeXMfw88X/26qA1gz6K1WAuWOeAYZ9GDj53wyv8ANkR
MiwYjyTuYbE3W7OBZS42L+WMXSWS9YhP9kYVS9YXpoOGQzDXGyxFbyDQzU73GV4l
sIS8G3hbKlgURm9670zLY7le3ENbho6dlUIPaRYpNPJjFagBjRMWTuj1+jNI8etu
YkDcWS3Kfi6gFwaK/nqbSc+a9n1SfuHVnOAxVAZrrl7u/nAMQL9E3GtfysQzv6B/
3JdbMPjqKL1TJ+0RNrWSF+Q4FyS4KGfwEIwm2agBtloz13wVgPSK2rAy9FdLpM33
73arVO1dNtAbpEZ86yi0+MW2dDAIbgVgFegGHuNX2JVfYhmJyi4BMjTAReaQUNuY
V3vnzTFuPOtfqNoT2SprP52fS4llQb9q4fpAV2jodFwuBwXmDJ6ZN9j7CbKVbsz/
DyDIEhg1/UsRkHqZ9RFFhPaZKJSQABcgI5qlO8mH2JzJ4RIKup0Xix+IYAJUj2Gi
RtrlbQS0m7jTy7NjQZJnDXWH08NxOJXyhLLJNEuBDu7VDYFXh2ynbHNRWObv4AkP
LlAsyLURfx5oQeZwaasv0grbhfBPbXe9ZEKKDSCcCJrBGmlwGH+5J3bRJ0PkO/4B
p3wj0GwAIhsZecqW0peHbAhrVPLwslWwjflIW90E3n8wDmoTCM4JMCRjqfIUG9IK
S64Wxo+6ZSbDSplOuOtRY0uPQgxlbt7ZFLyIH1y77UWbq2t/jJfr7R1jyNA/fF4D
nfN0df8Sq+CM+ogXiq6cWXi01y+HNYJ88Cqr+7Z5xAcxJEfj61+kEnYswUMh9T2T
fTctWzajlOFKbkqtCO9LjUhnpRSPmZ2CP3fb4dzq/iFGfBEccOwHxRhcsM+UyC+G
ZFBp2CXJQh+CObUIS678f44GU1C99khOrt2K2AoFBjTSVtFtU5cYuG+Iy0ph5C/I
S9yOJcFJcrLLpXG150tTG5CukQ1jOQR6CM1ufipTDOC+47C1xrbNKpu6A/XPojTG
gtPHkeVDW5VRvlPsr2wsWwp1HMBEKUxXDwytpdxv0RzMVYT3nVgWDVh1yiKgLJrZ
1L0VahYAyvt4gsDeWDAhh6/2MUllC9RNEKgehGuBdbzhNv0AiT+cJwIAVeggPX6D
s8u2FbnXlPPK6VnHJbyhfYXL6ZzdeIGU+P6NTIQbvoVmsUKaIsP99n2HWFpRN+u9
yNJ3rlB9v9Z8tVr2CSQMgOAxzSrQgGSUwQj4IZwend8SW0+vFadFroE9MXcUQlcZ
RI/v6OCHXloOkRoKFPOj+n9Sl7HF+ELvAbmZH3C4EZFTUb6RBNwfzjCRhXIcplXw
UFWmUIkb53PxD6uSSNiZdi4ikKoGWWZ0Yi8nB1qO/erklg91XfBvNk0adbxfDqZr
P+3LI7ZOVkwSKNyB8oEgS9vg6rfdK6QvWrktmNTxyxXYlweDrUlnHrWLPU0Jme4S
ePAA7Muf6n+BbpWhNiwQ3ma8B2ayK0x+OSSCuLYaMhyMWdefT8oLEuXXShGr2Sse
qfRC86lY7JqdeepgUOQadVbuA5jbPCKlmRVk8ViXEKe58xBd40wCM0jLqkdxehWG
UrOyUVvsjIo8i4aoK8scx/SgheKroCxSLxt3nk6WGT9C2xLEsbVGJ/Bj4jNeytJP
a+RMVYGCI1hTnh6Ydgv1DU3CU3pFC5F6Vg7R818MkDxMMC93nUsdwbZA3ZPYtynQ
reIYfI7l6N5wTEvxo/Qp2sMYCKayNbvG0lOQectKPj5lBJKXBeymVjiNlbRJjixA
OwMoJek3TUXfJtjNLBxxW7EcxLnujieP7MgVSDoAFBpYSaZnCFg3+Yqm4W52vElK
HFlMcweqJmhuMM+MkwkClUbqOM9ti0NePcCw6/64mfxA/VWwVNqgZbFhLzmZepK1
2gaBkFhRtpEM08JrdidDRGOZvGR17BQHw9STrQaSEZ/GgMYxjP8CBm4q7KZmQELT
ISzE5CcLu2OrYgdvNOndenrWxhO7Po0qTVYDGCQTKkrjsnpuG+zo6nlm1CxYIZCl
OPsvbZxsnlDhSyOP387LjPEbkjI0/SLQUPlWPsJrLxhau9d/y8V0nQgS1+qAjFhR
1dkHKeg9ZQ8qBwiRAqsw/gIGdyNRv4ZLZO9aYX96TIYOc2nGYqLEaKDR8tuzkcOZ
+fXN8SRIOarY9kqJu/bMpTqxz60azJIZgrgFlHFQ43nlgw0UQD4YQ4o1wwx/qSFj
Cplt5LKVkKqkjPSk4leG1UeEHxLovcuWgrF+C7Z0qBlwVdupjWJtpyhxsBvPyXVj
SW82BvjVSE3wkcWk/qLQ22dQc70+SE8FL9dNo4dVH999uoa8iYiIjSkMxtbYDK6H
1hvk0AfZ4dX0aFxJuccmFpoiCTlNntlnOJpDNIaxs7B2bXk49uBMLrUPmQcWDkv/
JchyYFjaqnuEf5gwcB0M8nnuf2UUTj2SA/oGMtkjNVZUQY5xjSojjvgosJ2h46qm
dl2va6OAwhAp06740gqO8ehJZ5Vj6tqLKhcJZCcF2Nlf19rYc9lAH0uMunA4llas
q43EpMuc9sLt6yxRtEa2v+jLpUho5KMmnr2wJ1Q+Tq/h7RZdc+fWqjhVWSzGHh3W
wzVt93BqADfvXZfWXuWmz32NfsYwjOUhgFJVPyLfcTFcdzRywwTsOUf8mJlIa6Il
OQgaN7VxmFRj1yrkLZ8ip1y628nyGvwPKenA7KObGItjWCQbHpKRllsq+s9frgm4
19LVXlNuG1jFhBEmHSnNBGuR48YP46a6xK3svYFcYYUgB8oE+HPtSCAFNx43CNv0
geVQv9qfvsV7df0ZnUvPMm4yuTBJb8f4Yh3ft8kLRVQ6ZVIo+mNN0il8Mj4F7fmd
gl24HBqFwVisfo1h1yWpzdzFtZaG1h6xEP/u/eTW060Wd8O4NzEKtbvQ0dqMWQTH
wcODaRR42jyL5+KBVWOMs04YMhcNdAbz/ss0OmuzvWKnpQy1gKN0rJYKvE4AU9Eg
Yy7yqO52z+ci50i3qaRgr490wZnlmOad3iaU8H609zkIcsgsnPzAaa6i0r6Sru1z
RmqnXmi3tylPizBVWAbfwTHUS6Xa0hM2hXf9tDjLqG2TM5x+nRAX/ugJDnKmCLoW
73CMcb7/VlP2Y2v0DJWKOtjri2OVNKTek8saBRb+kSFjdxhJjjk+wFpUNZcGghxG
WkYfzKO7D8zf/GLw7prLmz0+ntWrk3I4x6qFdN3pvhdY7Z3ekOsgHyfYJt//mDSp
mW1Rm5A6uvbZ+G70sFU04XqovbKfZ+MIsw7JWgovBvdJUwCy7x+yMI6+StSoWkp+
laNmigRCFy8VRJrFCupzpxQDwbobuyGwwmgM53Ka4S4hHynO8vhszyvv9oR8qkjO
r3bFVDrkFIZQ6aLABBZ+YWYyWn9fG6B+C9gMHGghLm+O/FyfAKg1K0YVTTfozSO8
MPhwbJpIgbUl2jANHXvKIiuODQQYJneaUD2L/4J8gbSOKySWX1ntDWnrw2wm6X5P
/kiAH88GwhTNvSDzroh57jZJK7yOs3sUD+bJf1gUggQNUv8rQ//ByA5hyuBoSj99
r7+3duFM9B1Kkb2GiVrXJ7jxzId8Kz2An1ni9pRug6EQuMnQa+WOr/CjE7sIlXw/
qgyEiRrv6YYvwcTOh+99tL2gTsbnYFoHM8kHcmfDRNuVDFm0O9tRWkUi/Chiyb1Z
rOOW4MyJdUzS5ww/ydgehTknzPMTF7NjhFmra/4MDLgRYBIvAWCGJEEumZrPo2n1
1UvRAcD2Evnm80Ak4AukBu5OCZvjV/RqOfuK1wc/BUTe5NPpadXv9xt/ieh6phGo
W9x4PSEoqZawGAACKDPuASNuH11uoBl8S2UqBiynsOG6UxWtD1+90xIdiuV5o7de
HC644JbmhjoSdkXRpgvLrxc/feL6HgtCDJIPSAOxnZq/iDkUNuLFab59w34tLm9U
eoPggRwNfTkSKJSems/4Mt2PiLbVIkSTlsMB1n9ZW9+IjT2o6PYzTGxtsSCMfPvk
wNquMDgL+3keqToNqOfyPWvgNKiKQ8MKRX5vGwhikiojSAP35M1QGv4hHVrlHdqp
PRFDjFYGpzL3JC8weyNNj6dy3eAo2ZbwphnouH2iux3sedbwALfdT4c+O2mf7s4J
GNo7RD58w0s63EwK3gzHohBUgpN3jmrYhUBmaIBJZfxN6TE91clB/RBDJpcj4t1j
5MdtXnMslOGN7eyUp0pHgsdQ7rpWO4y09WhBjF9e4EwhJ1syvlW5Vn0AXkWqGUWz
A4iaCHi7VvlvzJ/Sfc698GYlV6qQMpStFKTZB9euFK6RzaXScOilndyth/a9t55I
pl4rZ1/y4N/B7EmgwhypDns31Y74EsC2Fba2nW87FwDGJgu3sCu68vHfqwHMmgTI
SEyPeflXwrgZfQMuUf9qpVjf08zdp7T+IVkMtWspUOdb1fpiD2fozGujtlCmPQtg
gxYQDPgJU/db4gfy6WIo+tP0qE2vWOQO/SaB3FMdhTD5/trd1Qo7NyohhM10Fgpq
F2BYFQjf4qGv/lBDAmcFyd+iB6bFACDmvYy15c17si5tzmiQvb5jjUGuxveOa7pd
sWS1wYmMP6Z0X/u/QBWoTag0cRckOrq9142a2GwR4ijIyt94LXLlXJh11kIAnfBi
HxNb2q7GC6Pzq9EToZplyBTd4M23FqmjqdIX0U9hVdp2ZQdOvNoHkpYCZpCNOmrk
QAjTmS7dRgd7P5AgyC+yVqa9GE51US5rjpynUNXIR0akmLPz1sn+TyOTS6jLNmoF
MGIrmyP6k7aHG1R+nI0FspzAIHlDon8lOZ84RRM9ttT+mDubedDPsMCFFd0dGRoO
u8EjTu0B0nPJvckiuts7vtBAInjEo2pJMhsUvEn+kAAlnNP6SbZCHTAkljFs7SPQ
1XbAmcALibJvHV2z+rASfEGKNLG/wZzBbbMkZLs16T+1D3Mhx8Io6KfFaj4QhvxT
h7Zdf6Y6O5KJQY0jJSG+bDmo0bkgXHmbrP4f5RBk6PlAbr0de8Zt1awHTKnRiodR
M1izl/8zTvIMGNf7X4Mxe//S05jMXb89Dz+x5arEjwQA42Vc/szSdLsJIzRouV5a
eZIvMLEyK5KsUSvcnyk0J17oZDoQs5MfUBvB0tJvtpUHNogLLNbp2Ke+1pMast65
RRfpHBwiDt8M5H3sO4gl950KONbrFOaky6kztDFcy/rXe1L954eSkrc9YPFwG5xe
gWSHHElGS09fdfylbyjO7OLzeWfP+7UV3OaL0w21wU656JquRcKMSf8xbFSriTvf
u4aPeuBuR6L1f4RguKl6zNSLyfny4aC9uohDpIKJn9Vea9NK3c2Y49baDwRj9Aaa
kdu4r5r4JrxEw/fsnzkbhHeYDjYATkUKouJIOY4rxVU93ftMvGMj6qPWUfWcB34G
npYwIRXpdi3S21pWpfkGbqnnhycfooxOcWuNi/CyhB+hCxDx0bMs5vTY9w3fYUTS
NGCuFOWRIRn+t6+McZBVnpkWBKDHdZuh0aIqXNo/bK56KesnDpgCiwgM1NiHVbTg
u1cCCfs0Xk6Omx8OqNDSXMAGiPJN9Eexx9UHrb/EjwgQ+Mk/GFOBVmlq4K5E3g7o
M7UFwlRYLQ07OhkYwmGLIku0PVCwHz8XEXvXOsm4iMYJNUQmnemB9oriL691u7na
DUuNBo/VUeaLdQKot3pX7X749tTCt9I/xEv5hB9WASQQlkyO0cBnnJ0EoJ5V9KY1
5etpHgfo8Pddrv8lF7GBYXjwc8kDdnHWKvQLTcQuc0e/PGgn4gShSGD7jEyhCT5K
z7HKmp0xXEZGRgIs/vgwYI7nUO7AqM+F7C1ctTxNmbtnq9s2iH36CTVjhFxShaOk
/BvuOc+iKOTLg6Xh+5dpCSwQL9T+5aLFAQOxiUCSebdsgCo9bZ89P9TpjFC2jn+f
8OXW2tmuFSdqmJn8V2PvDEg0Vt1MMAkzpHIIxAoGrgHoUCXezMBYc3YAvKxrXUhl
Wcf2mWYjNFTNRPlWZ8d7AI4cm3Em7kZo+e44u+eAqqJ64N/06O2rzpwbMupImC4I
LTs40XXIIc/bT6W6OO5IMt700yQRxE2OT38jBfEUY9y4Nj4nOGoAnS8gkrGI7+8N
aiSWFDLwwrK7Cqn2tmorxlwj9iTGOHYADFTXnzvvjikNybWb/RxPkFD64UqL58BJ
3pTFim/6HrYleYgNNOAVvAtS1bfy8Qbtksheyo4Keq+WhzA8A5BtA8WsnRyw31Rj
gMiDuZS2PqZJ20XW1NNtAZxzyLTHo8quCJe8o1ZsljKrziZ6kuhpmlPsFJBuKKpM
HKEepJShmjjz9g2VQWxihgx3Rc5DXJiUQ/yzCGGC/Wjj5JwiaSVN3FO2EyIHE3uY
gWNI7yNg/jGGGmoz9GPVHzu/gyafpKJRKdQdD+mDEA/AT+9BFQXOlHW4yn7+/QHr
J5hto3qkFwbdd8rPLOOYPQ6w1EYPLWC4I59+Aa78Wdf3VooukAzkB+rOwvtLc6Fv
WEj0Dgtfvi2KfIkXughNur/1DPCHaDsjkMcQubIORg1hNMySzr1gtnFW7a7XPhoe
4fI4Da6fCN7OjnFEh6yNhQ35O4MLj/HG2NlaOAGN+pMjhFOXfpFDMBge2CJMHgdw
09oz7NJMJ3EBQxRwWHXHZyUPISc84sU3+g/9RzusFV+X5G9eyzllyS8lxSZ7wbfg
AuWzCDQ6YNV+kweUY67wANhDjzWz+r9GYeVjXRITOZxV4kmi8uAm3wMyfb1TqbaN
iG643FxN6MLkaILxw8MPlgYI/vhNjwY5vry/72cBJfMsoAppWnrV1Z1bXm6kDo9L
nFEnKxfRpeYXdtD/tIXPKLCYtOa+e+SqggmMVJmLD9FHmEoYi2AhNaivD8rB1MvT
obGE80EUTgniJmAu3DOocvAAm3AziOG+BG0XZhWzaTBS/UZOz/FbKETWKP2ZVQR+
LfD+d1twqclHrBlmHaxrpupQR83oTwNi70q6Uo8hSdSgt+s2FzR5vzZh5tyZiM2/
AxZEGVuXilClhlhQclVbA7DYJQF5NkALsHiNYG2kt02juG8FUyy0VFFyTK9XjEj3
3dEhdO3exgJh4SkPYwz6wvfwzdNuW4MYCLVHJyN4ghknA8qz3Ce+xvvbveoqceKI
V+9cXhGulmz1hLtOa0RutS3k9b225yNzbxmKTggmbj+r3QrVMd6IJTPLFYHz3SFw
8r2YD8riQWfYfvViBkamnD7SoJyIacQInLL4ZmfI6K7aCb2yISAS4uU0qrXzCI7x
V3q3BjgOcL4CXMIH+FO528HfaDVZk5zkEejAkmqZOBYQNrP2TQLKUWuo37N+vy2g
b1l/72PRwqOkqeal9QFpnNSA+PBfCEyP6ztFhwakaelxZdMDLzklAdVlz+ut530F
oYpbTNURoSgvbAARnuCkWO6fz5s49BvV/1n7S0L6I8LE+/XqAjmPDpxlqJWHVy9y
4aVD9VZpmVvR+1Qa3y7TbhER6MS6OsiwZJO1MCm+ZspbmpeNXpJTShElNyuKwLKY
C+hamQH/DT9XTMSgLlsAhFpORJZl0NKis9Vw76j77HFMcNznDmG/yuc/i4aRG8Gd
O/j+7nB86xdyKbsJ24jj/bQGqtSehaJm6SsMqwpzodWm0D1k36th8cokBhQ/pWXD
96XP4Zd11v+KjmEGhWxDNSMayDFRt2UlmtQHJPeZhC9x/58WaV+E6eWt94/uqfFe
MgIh6BBwCUp+2iD4SO13ujntsabQXZcCp6MDQzzu0KtffVuOhNS0CeDPH9eYi3Sm
KhlNHMuq01vKlCq9hZ6oPBOoZZe5Ss2Yq0l7GxETdym/A+am98euQ9R+vzq1gFlk
8ETQt2n+vkv5xbkYoSFc3w0yPsbnND072MR1+ohj5/Hx3eWjGfq9MsUpfPWlrRHn
KF0keqWdkqdh1agRCVdFWsd7O/LOHykQMhZuPhXfZyhWHtrONPK5OJ9SaUKLbwnI
W29Zue3Wq+rqJbuhdoYzeUsSfDSKB57vznKLBynACOnXwtW/3Y1V2dX+nPV+501p
szMqs3WfXApYqMws7kWr+wEbkGuUo4Vn6WPHte9miQox5Og+3o+79oZnMyD88BV+
/s25WS6T/Ut/Is5iwFIxfAB89xxRYstvM3PtKZhPSJi8AlD3Nv75cQr2ZdDeK628
1N1Pa7TLMMZC4uSiig6RsnTyUIHUugAbyry/amW+sXdewLrHt6IS5Lk7og81zbCR
clQUxVsphhbGcEAN2haBdQjcu8jUMoEO1JDGDH9ejvCvqAUSyN82E7ubu/HxPTMT
PoYEvXdUSsqrcSXpCbEVRdXgZiPqsWyG3nlbVIgZ84UHarzCN+Cw/E0bUlzHBeLw
k5JzBTzaMIQxhpt7baL0W+WUDk7vLG7e2wS1hF/92LPZz24p7TzD8R9B/N6CI890
54+37UYC2Flf8f966UjrAPkQAETrGPHYKi82uSv+WJozEsjfB+BgtQe3QUnufzKB
EvK5vZZhwoMDezw0Qq+237GY9o3YRrDgm5/VJ+zw6zSL1GsDvwqdov9Z1EO1439K
tx0u9/djw4qb1YuugpaV35tbdhTfsUCiGm8LNz7BYOPFffoDTfetgDNSH80ufuKP
G7PAhjtinTGgr7LfWtmqjIoofVcf71mcI1QD0AtZ6+yCIYYt92JhyOkb4k1GNaZu
pJdhIZg+1PejjkvGNPdrfU40Mtp/ESdi/gyfB1U2DlIvI5rnp0AMhTIh61cvWZe2
4DX+pd0/0VbFBJGaelkKTRjgOh9WrnhvJ27AfeMFXc82PKR87Ar6E/0E3xtszZMi
YfUCKft//k+5itV0y857/IQZdpC3g9Nn3BVNTG+imcufSP+F7INtGzSxiKK9F4wq
ITkSCuui58kgv1tUFgYYCJK49hIXBL65IPZIeBztVgINUFuYXMuQZ74hUp7CMenU
baOLKk5e11RamK1DeEUofx3iK1n8oCtbmUzry67bqvriMQVLVlJzMGMu9N8MPPk7
+swMSk2oB6yCbTN0C17O5gm55TEqv7MtQLqBFu1mBFLL2nN0Q0iM9x0jKa7aPIBk
QAXc1IIzQFoTIpfncDiZt4Zrbvw/YYYPWXUx9Yp1goFZY4zLtxee7UZ88+yYQTMo
IkU5FNF41ObZaYkggvx61dvhhHa88poHiGKjl9/qzrJRElsLdz6gsigfzNdgqAM6
XxMU0emyuAPTYrWjcEcb9p0MkiHmjtFT8yPcfeonwN/C+BFJUv6dObmOo8fV4nGz
PCNJ0Tjv295HprprLdHXa7vdop6B4gPwc5b5S1OnOHq5wT7LtM0FsdInoQVWoLFU
d1VBpzXCUXPKpQ/r9HK+zPuMSuSdJbZjhruOYHbResLNsLs4Sscd9jEsy5JTWhxj
eyf5ztXjfaiTYlIqw1ksu022KLb5Q2zELeHrEeuII+R80/HFNEXhpYWM7dXRtcBx
TM8dF+Z/0M2yxbU6+qS96SHR+BzPnSMI7MifmWTMMSxUIYTePWAkqQzGeXraO0WL
ltniy+sogNuvlTQTaZgksyoyGMuHCbo8Xmri51H5coIb6fRvMPg6QTgQjiFIXfIQ
oq6WfwHSqzuKm8pafvdAF9bB9n1g9ySexo9CIltBMPmOkEypCdSniz1mdpaIBGOm
Mp+l7USkjhwIfmliGVeo/M5RzrF25X7UmJfF4DD2V9pY6PICVW2lzULMJHpiLF9Z
5TReC4VquBOE++WQVgVO+/P6W/60z9GWm8sdnqOpM/EHsMs+TsfPaO4eyYNQQncg
qhibordLRPQZYKe+nRl4V0wRYHynlnVzmnwRKyKElT2yJpK3cptG9Cke+45+LE1O
7KASfSvAhIMgeMIwc2nZLt1bSS2K7l7LL+RZp3GUvIKU+5khWkPIYIkhis5qt4B8
tu4mOfyzxS7KCPbr0fRR8EAqGR9DxpHqerMu8lx+CV9RwrOH6Z3UZUe9SIb7XIRg
T3zcjOFM214jacyP9wdDpDa7/6gYsaj2x7oklYepQovfL995yWHlL4mu8MobcRJK
38XpUT0yO82jC1/tPZxQWPJfFfEzed+2seMNj5V1p7UbxXjjUIrtYopwI7QI7N7k
SaXESPltTYVeuRu+PeONgRB4l+2StXdeQH3gXX1JxQ2TzEb8ph82XVrQroTshFrq
pALapzSkjC408vvflAR1lEjcmYuPYEanp3tXQY9Ib+kiJ/HBqrsRn0+8hGgOvps+
hCbZZRg6GGa/ABeX/lfmaN/9XFpFvLaFGmlLt4KS6YZM1oYyGnpcSVW2y7Q6QAvv
JjWRTCSlboxlHhd6y8grRgYmIin78xzKLzKIRaqc33fOmEhfSE+wu7t5cAK29NMu
Fg+BzZw5f2Wme77FPKrjv96cxaBJcL38YYC5y6aym7GwzoUoUdhyhGtvuUOvxgFY
zj/bxqyzsqHoSuQEnGyTS7MNWN6a/sko27cuZnvlyx6O5qrxFdRddwdlwM5kBiMC
3qO2ACKX2oxvClrINudRKvpZiWiZJSImCGG7qrp2GvcMztujKfC9VhSQ6DYQulTL
aCyTMksgW7+xNa8ePhx+uKwgVVUx+T35H35sPIVywy+dvgyQjRuPHzoSRUfkQtiU
ps0N1Z5PDurXtRpT4lTVkVKgi9SHkW4JfW7sar/51cvOSCNbdXkqEYiAyyEEvFoh
cXqpXV8Z1hofuT2sRfpDa7a3pRB5As8qrmRxxt89ORoDSFhEjMguR9qHEh6d8tJ0
LVcqaguA/R7p3hgtuXFq7IN5OiwL2bj24S7qOlP5sFLOnZgMgdB9F4YO92KF3nKk
HjV0myfWlRxtLemsagrflXmo9V8qb9xzfZIzuo4/TEwLCjeIeMt1brnplqoioLLz
Ix4TTbQkd7/9OKcjfNDiG4g0MyHm6K2TRbiPn9g6/s2/OXMStfxz53xiwn0d2dUz
yhqU/i2BokSzDeRd/jbqNC7ARyL2BbgtV2fNtmue/RpzhSHW1E0Z05tY/ORpj0sC
U4xcIY2ierdxbs2a7NA7vHbuFZeM8K1YktbKjhAWisEOdPWwrIc2lMIgm5Md+I7D
Rjm/GhFbvf7+o0ExWFaN79QAHv3tUagymTRr9+G+1++rz3W/Hk6nBkAh0Z086Dq8
rMlkQnmlJupVU0/LQBaI4EV/RCa6264qD7V6QGoC4hUF9iIbPv8HYghvU89OjGcv
n6Ne8WpuSyBSalAvn6LyD/F1tbCQw4Ic5K3GJTAaZj+qhG2P73/qOcMXNOcj6asZ
+Js/oc7DyRlgfrGFGBaIjWSfmO1AhHQdOvQrP05nlPY+9MD7PA5ZfapaXnqJLNH6
7ThF/7WSZbxmm5tpB9shAaykLK3Aq9GF0YRm/kGwPBNFxUDdgihBxkOCyaZsXFtq
ru+gw+Oj8CzhRS1RldsSmR5kdcVImjP8cps3WYAQqch3PodqrEdux3vJFu2x6QGZ
aPKkQWdbv7U1x1g0Zoj0+CbzcjchzLoBac7seD56GkySk/kXtoQPvWjfa63pDezR
bsQMoOIx/esZQ7dTPcYVy2RpAfQApW685e2AaYBpmWVARMoB6URZ1TQF/48+X3g3
3sdI9dVN4UyZ3Yc1who8QY9CaqyEN/S6aULALiCaZSLTndRRQnfS7yq2Xyl75okn
Y6JBOxsLjinOri6AjPIJduAJtSWj3x7DDHG5oQt6fD7qEazaBvfho0iuxpHPc2hl
6BkPLqPL4X5vrpnNDCfob2hpt0Ii9NSto9NQyNhNF7ViMpH6/i0cibShkP3xDGba
cxfGrt5DGdgANQDZhbYLPdgMQfq0c6ihJiGPo1Y1cRV/JgQ+cdl65B2grBHm/FX6
9EqpoFhLnv3oxwS7Vu+NMnIWV1DwVJBlolcPGvKzJRT8qcIA8y2UeeFA3gudVJJy
sKZgkCr/v7xJlZ4WDwuFdHBf6GQreBM2riG2NDHuVX/xgCNae+PISKtMejI8ibWP
qjwp3LXiolbZBPvf+vamfP/DRLb2ZNCEPdpRtQma+zO/MrM5UlfjNzxyBbV7zGaW
Btw10OP8Etx/ONrbIVkldwC55kCS7GEarKMcRP05CIFS86zqe6T69684V0FonaPE
H4zZbl0Bn0jkSIw5VzUr4hWMtmUUUn90tnq8zjskdk7u+QnPNbDXpdV9yK53I/6/
jOlnGoGnXUkWrUKURlFUHp/aGdXIaXj4E8oca2k7/ZntLZ4mBjnyWHhv+yipTHGd
ALZq+lm7548k8UJLOPPv9hEKwpxx9Kg9CwSQUgKSntvp5Owr/TlgbRkHF2cTN9ca
kZFYj9vgYX6NuGyq6SZ6sHFrSE9ujQ65xYMgNTUbwI50aAwbDgPp571lEE9K+GsW
HBSgSXad96WSnSf2VSW+nsuEtP6rbfdYDSoaz11tONMBg4O2lHGxPwkChVTs6R6+
yZlnvlscaPt6H2TMMf58XAsj50kO5a+xIAL1vP/ofbEMPag85SQDWdgmAyvMz7HU
CqWri3r0sMT2HYD5S9e6tb+cG3AEHSpkf9rs9qSubzxKCdThZf57aLrcl5yiY3wC
zdU5tXSbrpTAS7/J7OMe9teQoeLmeGNRmq1wUK08+KwQFcBdMAbFGc0YvJlNq30I
UK6Vboy+tAmQ/ylPAddsPmd72HHU70gVDBUbZ/57kNiNSGF515ZLMkxfCWIE0Mif
47UvX9jRZmbp0bZTPDZJUCyviYTDzxbxXdXlHfkfH+rFfrG1kGsrjYghhE/eDdH8
/q5EWCN6yfx74KxKdnkZyN0Fa2DRC2t5fXIeYaGF/70osnn4JJkYiQf7wpqw+U0K
rRvjkGLERAY+VjT5/4/yEQ1wIodyqSIG31qI800eZDiX31+lt/TMNOfTWqE0RtWO
KGo+gF4ghETaIWhAUF0drhtbFDOg6r2hy+s0fG+eSMYryAFPZKuqOA8zzn5qpoQO
oo8/LVy7NoZ15S1ctt7xJdz0iPr1q2f2FuzubM5nl9WwSve0G2sUxZMm/ud9uuTh
YYtfXlCXwK/LMJJJc0TFKXMTzO4Vy6BM7f/pM1dc4Av0nkl3fGcf4UCvYambVvK3
d4yNHJcqAC6MJK1SssvM/juLTow9uEvXaSvfT6+1FZSTcrYL5b4YtFzYwhuMzPYT
P5KgDrp9b2qn9vR0cg6VdPH5043BYzM1nh9NBY8hoUUCtbzbCjWrjGWnyyAcwIyt
LQzV2fU4ezGSxYivOHqRJ5cQEDbvK8e25YeE3AycmhxO5xLhjqJwAaLs+JncBrIH
AbDpVOWsuut7rHOBvi2aq2WtDkE5an2GtpeRh9rVGbAxwVAv9RzIp5BTMlmLcL1+
sXq60cxTc3yfgLoYfqdju1TsTtNUJApz7Yaxgl974t1+JIn4gM+znWt9hhizjHwb
YMRJACd1iKfmd9qDkwXfdUm8EyZzvffTfNKOGhDJYdsO2T6ro9RqC1Gnsk5Eaes0
R+GKlsw6w2V26WXCaKe71oiWmMPVBzptM47huAd5+h1VHUGOC7hVkSVh4GSHZ3Fx
Il7Q6MLnLfqjKh3nY2XMOuFbJ2217n5aJrBA+xYJga7larHPn4CVPwnZeYAMgzuG
zQOL+2NHqUpn7QZ4rUNzve+ah36x3k+YXBBE3R2TxXUcHiOZjYJb0D+J7BPo8tE+
9FkSZB/+mF/0XwTT1LwnBE88tKahD0UZmrR876iaBuTkW7KuxVIAO8/piRkn2RMb
wDCVZVHs56fltbF0AmSF9le0aKYLfhP3aiT22DWR2CBtlflmW1oQdTJTlBlYDS8p
CJU6Tz9NTD4Hd95yu8FFXtJ5Ywv+eJpKPikE7RceCWG6bf/hN2Do965xia1as/wh
k0UTI4hmhqf6irf4XmXIyaEWIJl/HzMrP/k7Pg/Fsiuds5SJ3WtE4lhu4bTPDgpu
Jjxc2Svo273xIIApUUmicerxGy0OA8E3NfGo0Y43iE0EdOru0ZDeD4Njy9M97yL5
tyOjWjN1xlf3jX9+s8Aas7RKVh7QoDm4g2iB5wtJh4XUWJC0xfox5FDWDMj7alMU
G8c4AJV5xKPp/C4Ol2iFecvz+FVuFd+yxFIeF/KRRRjxLJeDYnQjpV+O2Apab8GS
DF7rnzc1MX7SbmHfxNbuV0NzcNYNEUEwDf7vVTbKaN+inu0RoVfJm/lANdH7Qr+u
SCFjv1VN4cDi1jcgz0ny9pGhi/mRdiEYMCGah1jTkPJUNKAif7ViGxldT+Rx2ulq
xG/A2aJnr+tuFJ/69rJaB/dYH72iz6lVPd7sa8bdMDSguTwcoG8g9gJrg18t0xXl
JrXp5YJZvCF8WtCM3MRh+teGXbdw4AFI2qV8LR6REFxpmnQXj0Ce0ntvZD7GQ4RT
Uq0kVrFrqHcdHjTwJkCK+XoJHMtT90C617Gs6SCEcKAY6uKoDLrKuy+Zc9uVJ266
oOr8hTqsV6cIzW3g5f5kKP+jhtmXj051qxD74b7OKH2Ech7qaNeMvL4OMv09Gu3p
qyiDDsc7RnyHeealOFJb4sTFQIsE1QOmFaFg/g984V71/qw3aLxuP3Zi+ul8NtSo
YhNhc3ClAJYfTeKDFH800i8z/8cr5LMyXFdpNS6HGnGUBaA/5RwWIygWq7573EP4
7IfFVE817h+6ttMRd7r+pSbQ/3P352J2KIFTr+MlCn5U4tpgszpy4EgL5Bho5R5S
IdnogIco7cTDZ7QuRg4VBHi+CX9tMKPOnvvbJEA0TRF1xXVrrrz2QEE96DIRGSeB
MhbIuSY3oJCQtGFlPX60S6z0dpUA/Ca68HW/EdXu0Qvxx0Bgvi+7GbpO4jhLcWYv
HK8QNM+wdcz7XHvsoFDEO+tW/HZ0Phn3xpyDg0pX+jdHhyB+Kw6zYCyKp6n5+/bU
wARcEFkF1dff6MQ+F9ReYLao+M7twAJ1pDqBzAfd52LBOcYANk2SAYUbZdTmNrOw
nE9GOF+OeKRY1l0sHp+PrQhX3d7X8Qtu6tiKgWBsulGqNIYYEbQrw+P23Dyw7TZN
yLCW61oKVsMWIagqTOtG7KoY2ic+FlE7xmAWkVZjMvVXPZjdVk+GMIEXfZL5lL7s
RC0cabxTAxnCMSqKqqom257EkzKn45uO3jl6gYpgOl9AosynNdepmUsvcEmPZLae
FgCCAxZUchxnASdl2iuqHi+jccl4JY+aQZxkcyChb+EsToFnwZ6PNsM8OvVOd/Sl
xiENkTScYnCdIClGClsPFsxh/sfJiF68K249lonjHD+gfZOCs1j8MfQllXo/88fX
1Da8mUuEig37t+cW5wUPnWE0I4atVd1fwRZzInFL6oWQ2y4TjmUrsl4jWMA0obHt
+jvQ5jSWY0Hu9d8mEMd//WrNY3OH5SdS/fV1Se4k9ZRnqVkVw/QFod1xS7u2KIyl
rU+W0cPPvQGJ9ScXpQBLpuWTUoXQVE12dtW3sar7RSzVmTRCnzKfK0x+OyhPJMkh
BN3wBp2nMwIsycsZp2WqrZ2q7wxNHYidFfaA4hCLLXVuTEGGAYrVl0JzeZf6VZYF
+s5kV0y7uZfDy9kzWVVasip018GiX1cH9Rh5T6MK4OtXyekEBp0x2ZLxVnn0O6aW
Rs8J0wfXp26FIY4YkgT+hxzFO1/9uH9zfgAd6wVjudVa7mLqLdAkpE2w9tBpfN99
4u9HppemMRrl9ytlzrxHETrs5MqH5nGV5z5o4SzS2TyCoTcXlzJAsYCyMSWRs6Ez
q5DDsQE2d744c7QSqFLgqYoJRag8QAPI6xIDTW9inboiyfzBmo0KSOqXC9v4DQGJ
nRgxo6sJHe9YHFijQ4IasQl0yFsNlJu8sohM3tT3nWSi2scG0S56qFBYzcpFf9Rg
7hy0fiqolkNPCy4MKHmCAZS6aL35r3ef78EMgEOZ6davYUJCpfWJqF34Xa4O9a3V
LcwfIvThO1AtlpQ1Xfp3KJ5Dr7KOqU5h71iK4eciAhNayGXHbcHysoKIR9rpq+E7
nDWprjZxxeLU+Z5MdfXbT4bji2IhLNkrcb4KsCaCbrkKZ71xHup9Y6nTsanjkIJs
RzXZ6ghwsPV/4bCN46S10JM4ZpSbe8AG6rEBwCaCLOdtNSvBbpsXAL/PkbmaPIEj
NU9LQ964TRUV0GaZDkCSt6SIBleBG312QYHTzoaikseHqLiV2wNHMJ+mKKSana8s
nFB7vDmf3uPU98K6c115Rbv6+bJ2tvV9jxyFwOV0qQXBXIyAdi/U3H9VwGq94RRp
yEotDEt5VhAUaPAPvK31jrRjCr1Gn1GgHdEgAgKj0n66Z7PK2falJebeyKKPjsbl
tjPafwp72NRj94wppHoaRxLzWY0aOWdVztk4XjOqFMkf0IXy+YrBIKhB+FPWu2yz
7pDguMQcbxrcjT63aEH2+2+FS84AGEhzVI4WVaFk4deTx8WHVxl4WhxkucmyJPdp
C1EOtrPv7I0FhHXeFZoN39hTzYWV3vPSi9mCZa/fnOg9XYNdvPUEDJbXRNfcF3kC
8XOPMjCjVPCLid5PkhtoAhtALj2+VmxSy/DZvGkvn10dIxctrfaS82jijzglvU9/
R7LbdiVdqx8Ac2zJyzHsGOf/NPXEJFg/tVbfdwtW7iNT4/6zu628lBrQMXw0XRpp
sAQ7CPzCm3UKnk0QsWsYpoiWANV08iDQAqKKK5L+i+aXqQTlwBvmoizEP+atOo63
/TwADVLRUTtIt+D3fXcaKLpz8BW3uS8tWZk4Y5Pbbturzoue5LDNrTWK0RVI54W3
YnBpHM8nNEK0WmrUqY9Vb84B5bCi+/jLc1x2AQncsjKqs0JvT58KGnsJPOVtvXB2
kGADMXGwi4rquDwjQlOeU9MhB4oK5P+/ZBijC1pKKU/v826GPySsmXqmsHQDVcZM
nSwOm7rWRUq1IZT7PCBNMPJiHtUeZxuC5PLTkH9jUjJoB4Y50AGwu0wjBbB/Azhh
cLIiPU4G7ZZapPchQrpx9QqyIA5q5p3v0v2q3itUVQ1faaoykIEOjhKqHT++Up2G
HLbeFQEFmRqkcmWerGk4MrDeQjP5viv0SBM3j6fG5imqwV0wGSW1JZAkEhaS9Y+g
BwsTdBsPQKFaOqetQKtrjKfj5ma6k22qtRHCARSklVPxh+VkpIopDZC6MRSRRj8j
HH2iou6IUNX1cwXPlNt9HF/E4+z8wVVC/Y7Ws8qWIqhoNf73Yv/5exQ2wfl5lMlF
DeE6ZUmHDvVDb69MOz4hXwIcspfQIh7GS3it7QCyrA3TkLNfn1KMLJWOWT2Wu5Fx
+TXO9ON8dOOcTJOwKKIPSqclXG8urnjtEnVDSLVdzrXsyp74oYAUgcjrZUNBCpPD
GqrwBZTJKDVCzprfRtUeno7Pz09MqQtR66odUcK9XG5t+nvdyzOWkSEfakDPastw
Egu/kEHThg9cvjToumLhejmzAuBx2UcJGdpXX1k7FnEp4EcPxMXbrtqPUyMs5NnQ
UH4C0h/gki36dALWeExAusX1zFg/q30E7YRe1W8Ijv7T+B/wwtUGzdIOBqXT4RGH
EMjBip7XPDEbtobmCDEWWWd8ZkWiGrDkkQLz/Dm7oO2zxq0nm6ef9mDTH41ncmZ5
O02FOETm5KlaCin0OYlklVAQWfLqaN6OQdjX5f37OQLw77EBuNTqAstEhxCoAyGv
uzhaHl854WB3H50S4tRwwxn+wuxTo/FU5AdBO1AfpT8j49GfEpggBLL4p3jSqMYX
mGZFWPp1T76wehoY5GEKO1JP76C/LNywUduSmXR15Yanr4nTYHScmN8FIOZzptc1
Cqmzy0GFKZiJNhj1cn9ri3FUtrAbVahOpxqrhzCaczPOg11YAbHWxxlyp2ipUcj0
75SrgnTTlUdJ/yb5ayyU0WZvJw9l9H4pT7pylFrUuI9iDQ3xUXTjCpSyqpt+ZA+R
gGEtaQoCk/GDuW14e/nNlRXY7uKm085nQgFFbA1V/0UlGXkLF9IypDOMfczndaWL
ua2/H2iqFlsEdI0DCGBsgipw7A+hGgLrLceOmqX8B1uSZUsUSrv4xSEIyWtr4lRn
JcRqFcrlGK3XCmN5NhuUkn/lHq8srwC26fkll1fLGLN6QXvJ/kQkyqfSlIfVVnfB
Uv7YOgi6FlomMLwJtW/vpPqWmQQ9c8iIAKrIfAkU0qxyDSJVpG2Do8rvJF+Ua7nu
sAcEIsi6B3qzDl9PS/DVfqrM88MDAWugaZ+XEWXXCiDlsHGUq1CUrtEmfKaMVgR5
OEm3U0GsKPec1RH1RVKeFhG9+p+xoRvPyDbUt8qR0gqz2vYC/sZ3JWH/pzvIJ3vP
p1o2bPm2t2XoKKNaAQ9FrpeikiKGvkUV04ou7KLDj5sTnLQYJdzy/QEdW1PxMS8A
wUdDKFqqD8cXuDdAVj0zjtGYuiWv85XvTpbvyDvqst9dgzDFLcRjP9eEskn0Y6xI
xbgqISqn+dA8ZFWpxKgHJDpxzULofLVByFEWVn4m9zZ2AqmnIb+pExduUhfTkuLH
hpwdY4ss+ml1wA+si2wQohkKrAiHYuDqCDol/pBp3aU6GePQYkDbc0Tdv/MD94jo
+qyr9l+Zld6pAaujcqAvTpRbFkYYvG56D8H2b0VINYdX1MsCTW7Oeu/Z6pRQAEdA
MkwuvxmYRhPXGCaOSk6J8IZINifIC6A/hGjWfiotvfPIPnwTEa6K/4sCVI5u2fKO
Yh70ixQMpXMpE6RkmrkS+DaBR2/Ukfj5FLBCcy/iMWPRlW2Xui95xpmAb4M8WilK
pfExb9gYEpXs7M4aJRcaujIs1dISGhnviAcBTYFN3JfIOnFoL/qcFvzRFQ/8AmBS
zYABEpXiCcb8A3xkPG//UASKh65SYxTrSqyKqPpbCZyWaiWk2IK1sub2czVAZ3SW
uHIaTFnkBcwZb0gEhhQTf4UMjvzo8Re2ICfdOFIQJLE79/RbkPf4Vr8BPctXDGmi
In4QEZabl4IyW38njPVPdbMpkRElQNsPJ9ak7nl5Zvc4tH4VbOvflpmpFuEtgUbO
jXXwaJor6LEHOC3FDW0Mf2sfozFla/7VDEQeSOmCZ/9p1k3qSbVr74Qb8cMgyUEC
FPCq0xOGd0aMEXmbW/GSmNlDdygm5aPKYDwwvkWSpuSD2dHkHs0+gvxzVxwsJwbB
iHhx/TzA3Df8Re92jDLpwueIJoGYwAF7VeFgzqFIZdULZbqfcG8mrLS7Ixno+5ZK
LjmdToB5dxsv/CLmYbZ+Mpcpm23MLDxJcJlFCvpp+/X+mz2EdEhUCGQSF6YbXPmD
8PH5gD6wDLV8fbHXauS//RXiBZXzQdt0nNt3mpKFWDZs2ozB+C9fs1k0xUO9Ivod
zu95VCpcpshQBbtI0QhvxL0UHiX6pl8TpyjG+7zd7lcZDKG8jkjS0HEuo/dvBOl7
HuLvAQL62xNmm1C1OippOdjPwjTcPphrOMU4cqz+GZD55xIx2WnaNsJQBYvycdjJ
uKfWk6aTy97QoWbvNooGBxteFpkmT4Tm9rGM6Gtu9SQ3IF0h4OnAWz99Og1BXq/u
h61xS5hvu0zlfNeDsIQMpZXH8Gc2tvGSKOSgRNuJUv/ffdKSXurrofcZB6Op5YWj
jSPdSlIO0pqydXta09ZWaiYLIqscMeEhayj8KzA96/JL59VfPgXL72kjlndxv6Zl
RfkHeDgXAx2sj1g7s8FZsKla6oxNp//Lun9mKyh+HfdfY+i1qY1b4uZp/BTuJroS
jzGypCYugoT0XKTrWqRbHxCguyZFUPxC5lnEX/yQSyjXfJeMv0E5aFXHCqHseUOm
NN2j5pY8XJiPIGPuVG9huFwx9I5QXkZ0QDDDZQBS6Rd7g9lYSUqPfkZv4StCn/0n
SEe9u/DUuEfcJ9JSoMcmZvdhhR9FDMaWZRYwoqKKgg8uch0CFELsBRURX+EBhT4G
XUp6wiGXp7r6EEROQtcghWX1f3RGehj9MRwVR+UEsLzJxo3WJOJVjilWY1YuHlYM
gnR8xDdmdMDs92oFlSPvq+9e4uFBtY+nD4SPCF5zCfvvq1Hnfpb0lxKoH8Nr8zDe
cqPCx3HmoR/O+AE5Z2AoA4dtMEZPwxEv+1XFIa0K/RzmZIekDv1xbTtU+a4bv4My
uj4KzouZWbnk6OVo7eYPqW+Q5ybVJUVhRa3faHVpcZRhdJmQ4Gq2vNxHI5vCJuwS
W835c43KjS5Il0dmtKV6aqitqpfHZf5qFTJHKQBPN1JbJKHGL8w1EQn1YDhagcTO
iBGaecuxPqJj7EWmI/bIGqGDzq11votYqccxr05xV1NiP/fO7Lu758jh+uFTthCy
f0U7gPdIAG+yHtUqJB0bIY0hO8iXie5Z7pUFszhRX7R0YTOWhzOwq5J4lwgg5sH6
qMlcspFSMF0QWfxIvP9u/7GoPr5mq4WaLh68+hqzhSfx2DWpjGzPcVzsHWskPvHy
mhglQhNP93DKBl6gbKxQolHFgPekFhqyuMgvYBu11YMSvubIIbI3l8H9sNz6uZI5
0eat0F9m4zo8zZwWnLfoDfcb3WkUIfDciFI7D+DugH4KCbB0PhuCgv0JAXDhv48E
kgBZTQuQMwzpk5DV05w/B8eUllvsHtxA3Xj0jpR8ilYtqhmsSWdnvxLEAtiLglra
bCGJjr524WlWq0iGR8M4sVLOPY9QmPNNoR/A1S+sao9ndwSqZR+EmKDQ9KaekpoT
yCaGtzV0qn5Yf/mpfDjGAR5IRuCPpYf5NpobNu1wgpNICd7u+T597h60nUn3HfCq
kSembBx/BIq/O1um2sHIvUpdnJPdLUtcfMXdj0y9KCm67RqGnAmBeig1JvYL57na
Roh8IBHJv4eNwexP9ZC1hsIDX2aY1wDY9oW4GoYTThNQB2GqY+HJjI0G0yDvIvfe
tbsGNS19Ah0MjGZEG1pvg+m7l73oYvUmwBB7N7DNO3bzKWs298wGY3S41e0sy4kX
75ZfatP4/rlJMqYgnEkomCB282m7QXtaFLdiI7d+HpFey8Xx/wxxboWaymq4GqI4
PsW+wNU8HKxJquMktpGptgvkYwRKenKfGjjCfcUpMUrOrNRrO57FLqRvQXum19yS
rBNQrSHAI8HBEM7bThGc4v43kPZLH4ufpAG7dN+rBecJ3X65EQ3CUW9Pzo3pHfRK
9q9sHCcbNmUH5JSdjU9DiQHEWnNZRWXWD32NjXH6PsWBfpW4YNCT+i6N0FPGrnL4
VVc+nXbdjIqK2LxmtLVGJvnIC6aabhDaGp3r09YctnKLE6/mtz9L1QAhq4Rps0kc
LoNreFbz6u2cdwA3ghhCxpdgWigIiUqx+lBoxVV8ZcJlzm0lIqcI0DP/qtzzSonY
uJgd0G5/okBRM94tHRkDxzk7gO3sCLgRBcUOzGtGJm0EdWpsPXbORu3o/IB8LYlk
EmPGCHcwwUyq3NQur4kMYmAFPTAB5QkO0FaY6LXR5rdK4A3pNolnIURw+9qfgUz4
6fIGmvAH0RvxgyMwGnMnwZCD+VRe2ROX6NaPnDESzmMnIXJVkXhsP9VBN6HwjxuS
GvUJVHAONjtEwX6EckzbUz4Wb5HKgSis+5SGmI019JGCJiujiS28lLpPkgUSHQmu
76uPizGzvzaqE3aovyZZ+NrotLmpaW5a8Xc0N3c2CNnjwXZtvg2i/uNWjfaZtRw6
DrFNCBU1SIM5XUSKijfJmio1yjyyiL3qn+IMqFzxAfBiKyb8rFRBeb4hvgXB0+xe
eW+OkSe6a3lGh5fDHF1SEFOdlOLDojM0zdcf2gaXzVlYrORhnxoMABOjInV3EIKZ
V52ZoLelq/G5HhpOfUPlUJEdC02SfPs7+vKBJ5b7uxYddZZXVeUE7Wcjf1emFmer
FTA2Mcrua89g2MXGGT1Fmnt6hQZFu1356ZROWRria9VFBoIV0fOQaU4dKhsXIGuB
kTOSA9t90k+kvIPlhIUvu+Tpi056Ztc5xJ1JQoPaWsmgaK69N5MQRvD7SRacKuoq
yzb4gOb7l1HEMY+Ri0B/3ry/4x2SKdDUJsLpFgVppbZGU04XH/8gVJ3hr6KP7s2X
4YaP/aiM5Vtcyie3zaj9dqAyPEh1dPGRhH3IHghYDNPK16URC788U8W1HI03xOvU
1NZoUlUZh1DDOPQu3inoccpypGLDgW+ERpSkGs/ClLrGHpp7yYiiCLgHh6Z6/VVG
U8vu9owa9adGJU7qgND1sYFMzXeoNu74nzZ60qC8A3JMdbcXdFGh5JnksVtPrVqC
ZA07P6Th+cMOAUYHnb2Ghbwmlpi1b8vSSy/gb4699dIasFqXnUkkoKdbQRBKsCGF
/Q41GsHgkvzvpJxdqhq/XU2hJlrPMQjvZSgCGHAFyawT9RjyCRfQ9wuACXSNBw3C
RCctVSj5NF3biIpd9DL4I5kE9Mpfgpw/Ny7rLzZxxsjjeD1k4iHI8rWtUUAXPML6
BLZZFM0Y0vTh2cS0I2E3dIUiivpF/BU8mvuQmQVrZUBtvO3BkjpBPJBt6apn9YC0
WObs2EhhunI7YNJlRWH6W+BaLM0YG+imQod05XiXr5VwLCEIRT/XOgsYRW1iP2R3
SqpkTJ8Tm7Edg5JEf1pNEslhKh4uw9ZQ6Kwm5bAeWRZdiCfyVAAWhf3GW7sdj5pj
mXve3zpjZjP5xVmwA9xa1hR0Dc298oVQGZ+Ml9/rBb6kOLfkEfICW2iuW9mibWqo
hUwTv0aFF51lCX2K+0Xp9TNOCcXpaFrfs/Rwtl2D4CWHvPIXdsPknWsPyqMhGY7p
35kpByk086dm59hYUzRkQWf1yihkPQ+ETCXvya14QIIlvXWBHTvrTD40GlzFjNgZ
lG4l41qOlv3n+syYq/nFxBZU02vO0dRz1PBLkgu7cPkNlvrImK1GXwBpniR882wG
1YKoFOUi+QjIVGBhnkxDfH+eVF2jp7xzpQgpX+Nk7UVsNGXiTQ9rKFzconzq2n40
lXNJCiZX0yHq+BmFfiDWq1klkATkL5vAuqpWi6sYZV11x6sPVqcKLyiGs+86tDDY
eH3giC/PvWSDUKBWJ7iSYnVCkZo0DTzLoZpDuzBWF+Qpp4+HKSVla5or66By5ULM
GaLyghINxx2t2D1SLrAWTfeXQ9ixalwKaf6tjQEr+c0I3cMKaA/rANR0mLHfPYtP
31Ze3wyDTjv3t3XodDZ+IyUQN7wh8GEdYIQ2CvbTMWySdLVGpg2xj7DJGTfQw00K
A2jKBl4W0jSR1f61JFiKps616SeLW+8h/PvmtdCfIJLL8+1TQfPUWDVR0IdkaCdk
Z5UH60MfMdNfnzexVgeSnWvhRe98E3DOYjwaqbuClcwUnNH4q+Vx3p70nItPUaIi
lOeVyuNzUZmwjwKiuYwCZDkweMEyUzYo0lK77MRgqSZaIv9M2cyGirf4Ah4fUibN
XYs0fjNvHuAIjlMYC05LBkqaW4aaJX7eBTU7/gVlxjn2FARhCBxhiz3ZAeUHEAq4
GPjOdxoH801GJF3+UMFhJ0WD2KLO8/zOxSW+1Wh8LhxZiQzXMEqozJZiq6i7Yeig
aOd2HEXf0Q2V2fXo6MODWeZG5ktlVLhzhbePalGtZglZn8ibLYJKKL37aqY2pM/C
Vn8ym5ko54utUb8KAuDje8nGkii/diwc838OH3HKPwiAu896yVj75cm/e4wG5gcX
6ukeQzE1FayHjRmqYZf91hK8UFaDu0WV04IiRST+qPN7NHYQzyn9ss3FPZAhuBYD
aF+nEzIb+Du9J9baHRT6ix9+AzABAiIu6UXwYqrFTVbYFk6lsudw36BcTFXgtAgp
cbBJ2BeP1R3Kl3yCHklzI2mxOldU5NreTFriw5U1r7+XnrLaANQlr5473zJIHS5J
tLv2r9Rr+2ppGT/RgtZhnwY8dSonbSAPQx/8+fxtSt9ShnT3jXDgtNbgHdzznuUg
WDROUhY2Dxb6+6ecmC/5H4RacuHDLSxPtsm+WjmSU5FN9bp9yLkV4mePUAgzbxsM
jvaQopPLKrArGYrFRXqGZ1wU8rHzgUPxQifb5k2u7O/r9qasDHXVTGlr7v6K0iJB
bTAIK2jzS7+9uj4EJsU8JdrFJefYww77QKH9rgY4qo8LfUb+t4n8DBfaVlY1E6j9
CyNcr4dDoJ62gbTOvWAJjRPb8KeNiWTO9jUUpaYIpOSdKRmnzVsqLlw2BzyEBbCi
ASOID4o+WsvRPstaS1S4Fz9KDSe3LIqLHrRCEaC9RGVDVtspg2obKwnV4YRKE/a2
0hSSDV76IfZBLiIuOYpsyJpeM9ERopT0rINojECBOCZaP1ys9Nl9Q4XPLBGzRhOO
Ai/rnGfWGJL2OyieF7JV3jQ0kAJVMHD+8zwffpoRioK3tRZDxDszB0fz4DpGhoGg
HLmb3Zv5V8lC1ydgygB46jgi7Ad/aTH6Mhj1piFvyYYpplx8zrHU+Bo5i5VdmbBu
bqJWDreurnm71qTbueVsafuqZPcqAjRKhMuBBsOmdQaesZreIJ+AVg0UnYdd7kh/
wPSvc/EwWEpue3JUC9Q9thY6G7FGlZTLo80IHVPXQcZxU+Imydf8WDxXdYtqe9k8
nN1Jiuku7CORajliAm9mYfFzy5JUhN+6eqGsyDHUmwCF9iFjHOk85TCP/OSqF4Ip
crNB1S/bxTXkggq5VrS5BQ2mbyA1ZHcnhm0c6cvXduDeL6C2PySQIj89PuowZzKt
u8fkwh3qYAsDfFWhkdOhGsvxfFEYrGBbBRfPZpcgEgxhcpSAH9JIZUjcKKekv9uH
8h0whx02SFZMHSgOXAIDcqCw5iaLzs/eN04vdsu2FG7jt0BKaDJ4hqBpyhnq1IGT
Wqg7EmjSgiI+niaRTpc+razQWbXgpimjYOuxKoUeaKO1eTUExKCoQO4WOnUlnlTf
qpeOQ5cwQvnBBEC6CXJLM1QM9t/MxhvDCfM45sATWZkSoNeA3pgN4Ryx85cBS5DS
zU4T5cUUMNqZUPFM106C7EU0vbolyXy++K1fVNncDJwVuyYeS8/+Mz+16PRpmgCB
hAB5K+XW5vEQVHXQQHiHdY+9eV+W85iZGQaegU+oKSrbNXiI059Qymp+XGW/L3Pd
OzJIczib/x/sbMFriWBPKDkV23wT3LoNs+VxUxVDQCc/HAx6ooVkVhxEPMnutL+5
HxZhkHOQbQ4R2SAyNAdC3LA/D2JQw60gFU7PKBCyAwQ2+Yp5EI1MqMXo7u1wO/Hs
MSF+F/DhSh/lGqQj0C6DbKlObWXQOPbMjnCAWDSab4Bgk6H0qYWCYoRkqdH3Y3Vj
vVn/XOmXSDtTUVDSp7hPRQlBAn1hsWzDodC00BEvQOrdWz2LmJH2s3sQVWprcVEx
DcfaVdcrtG8S/feF+4sqUUmkSko4FLAEcIN3ZZByKvTJiRed5MvwItg7No54l5XP
bzYuj9jEIUjO3BcBIK1gdmaedLeyY/12Py3Dhl7I+qLWmInJlWI5+YTlIpkgaowF
l2wu8HY4G+6zLhGnyZbGnMBezVWJnaGodEI/KgmhYdDEsnLP4I6aarurS9gsQoga
rS7Pe7OyVvUoMZ2nRCTBSTuBEjCndTQBauewqMjZf4y/j//9HMzOlDyGNV16Q0cv
8jlNX6dIDQmg5P1Pfmvg/yPHCojqDsNT8EMIS6IAg0NNx+02MTbwyNbKHjLlqWwH
iNj4hHL9EiVKkswY8VBHC61legKD6ZSl4AqfY8cuox1onlE3WWymuO+Bz8xXFDqE
w/KkxMN/AH2eL7qoYuUbLhkWh8fMvZtCYS2vWW9GcRFpY/46HoU6Cwuhr0xF2+sK
aWNeEPeRzwbWuxNRI3oWUmcn4xZs+wZU9omqQWxwJmqfkxickYKEAbaXQDu3yfVj
54WpdMZiyYxnJywe6xjduvUWffn2c2UnxF7ct+oCDdlh1/Sacs3u4tTFrPbX/BPl
beegxVLeBttOcUDZ42cJ0eD/hjUbn2zwIJR747gUSJNjK0WiTFMAv2vD1IZyB1R9
WfSm0D21oOBBY5FgHp2mAtmA4nVSdlQeE1BtQefRAPL78lP2Y7O+RCHdYqpWVgCM
eAKyFhHUkfkver+PGcH/LH221DYwkQspLJAYaiBlOTVaxysOxOr7YxYL6wEW/2nD
5HAUBeHZSi4mUcvkheVLWfgNCVxEAZLROmY2nRimbUVZ3s8gDAmptale6Ydp8eft
xIhvU6VKNsZdg9AP1uReZXM9hH4GHWp6dmjaPagdtxfyP2/TiMkHrQqWilkMC6Lb
0ZBc6NWeYqEh/z6iZSSiMCNXA1Dqv1q2YgZGIxoXe1bpem7J3xvFRP6sRk1yRF3X
6JwMpgr3CmWhYt/ESP33w1Q0SJ6ZzHCCzTBRuoX5X8k3S+ZJYNuseWjF947oNEOX
u66nQRT7GV3S9SHConwftzYbtYQ6E09HltJbhJUtsEuyd14Y15OhT7GIbIlKhEaL
ReEHYDdOneNTeOGZqPL7z2wiZLJUGRIJzZ3d0I2HuONZtD9jtErAWgC6VLMfT9AD
W4mNCEoGgERwEklU+pbBxL/TjAcH7ifEqSPmsRacYV6BMl3PELY8hT4jJMnMYpaf
MYFi1XV+mR0Yg40ceooNjUIeLAYWewxhxidrHNF/PzTmiUgeThU1x1yOPLZrZJK6
MUS55maAmX955nWuZ38Oi+oaCXNvecnjHp1HA60hVvn0NuTMiPeqjpmgd98KUZg4
hpiIWeJtu4cV7xOrRszMLbmoJt6e27T1khofuJDZcDBS19isEzXrJhwyK/YavJJG
unoqi80xobU1C9ezvqHGuf6hjBQRy11k404v1FWuEGBpsz32cGw5CA5mDPv23BCO
LNxTJR7VCf6jlmpQmKYeK6Ebu9d6zKGYJkACbVJzxObnuvOVHhF4AQo/rk65I0Jl
kejSSVjL48tUet+70+mPIPm4w7ZIgCLlFN8/tY09f+02UULxLWe14nkfv2QMew2x
i8vcXnwmUeirQ/18GyK8HLuHwI/7TEsk3WzM98toy5FhU/lRidP57s/k7EkOKGRF
hipdhm6kHqCCJU6XCWm0/PD9MAvUmB3HsJ2N/Vq9p243313oKP7Fha93olL5vND6
QCZLPZWUJcXQRbCzB3TB59HNyfHwvatsNsIr5mxPsTiQ7AHUAr0hd0xyFDXH2tL5
MDLitoglIYzH123Ew/9b0HK3fBkZE4A6LaeANHeRhFhhTAe4e8QnCyEHUqOO4CKg
5iwSzFpa310DRSswiVKE72kp+IGtVe0Bm568B+Q90ByzZGWvrTuycI8BNnpCX7Lt
ryRnnhHZ6HA0J6DXG5gzj9bpSGsEUZjTo7VOrNo699KoANKddY/RUDkxEgWucfvG
/UCFDWoepruQzGHfFJPWMquu5dTsIBP/2e8mFxqn80S8sHYJ72KOaundqY9M+khY
OpepSWbH0W18+gQwamalnFgSasKzNBqi2slqgqHO8kxlUjohqK2YZwc3edFcxzEC
Y+SqDDpRkZPYwbm7jtrOXp34VF4d2ZAXUTUJyZ7v7v4IBXOc+lnJez8svOKDK+qk
9evCDKSvD9ecsye92yRtTaO1MzAc+NzBa3O/vwkt97C7PFUONf8G0SvVVsWPEBHr
Tm+tGU/6LC53F+h3Qiu1LCE2ingCUWiJn2aVGUCVTfXemnbvNCD/i/jM80n1OmMu
QJnbpz31HHf6xgVU93flAR35AOESTh9AIQutQjTTuC4yRBH33Pp5CXjvQnt5crYJ
xSNfiSiuyTp+WoqrVYnmONCN1DhYXGrZokHYI7bmwg+BlKVMqRfV54R7vtzBTqx1
7ZZmUe2XBUSqUH+5ZwuP6UhAFgYeuLCk4E53SQd2BRAzgUIJWWrB17ZhhZvdpMyh
txbTycKdIHjHHnjTfAUKSBr6KSR4r2un/gXEEL+38jHB0zwBahQtxIfpUXge2VCr
nZ5TZEd5azFVWuOKkWNxTao2kWfm1jo7zTxfKjEHYPm3DtPcbcWO75gMLt4Qwesv
YOUB0BY7r3+yrMmnaS/r3Ir0cInvSaJNeH3XZVS86HjovO0QWAdog3V8lrjDqC0z
CYdSH/AtC1CxtTZbcKUr5Tx9vG0r0BXUx3tY4ahJTVISTJE3cyBpGbEl9von+r+i
fhPT1oWVSJJcTIc+6EMBUfF19agVshZsNc/KOAqsTHDgIWFKZM9DVIxHV9ItWIdX
rhndX6d6Jva8X/6rZRBVnLABvu1B0xmbDZHKWCRKlW75QGKuW1k5yYBdq01T4UKz
edSD1NQkuqTP+fxt54MXKd89D2uH2w59MqkG7rUJ2yKt31y38gsvdvq6plQgjS5c
h/AhvAriDa7RuQLpW6hSKoSjmur16i9jpHy4As8PGxJTYzFKgAi3CpcSIroXLLl3
Jwr9vxPiWapDkz367qoWcW6Bj723fyBKuhNhfs9EfkcmdMujEhS52G/vhpRvrWOE
EI+cEIHjG8MRk9fRcExTmo64l/HWsJD2Lk+O+QpGZ9cP8+5EaurUD5zdqhq/Vvk7
vQzMxVsC7FjPjvQerqTkptmp+6gNvChHXIKSpQTmGXBWao+bReBAKRY4crKF8tQJ
XTHekbbOBjOqfGyNsgDCpKZzRaqNq54E4mIe7MUt8Ms9H+JAxute7PYXSfs5RnKn
mDziPsCwnMHDkrehsidtVpQg/002LmKfvuq2sH5/izXxQ4H5f5TSIjiOmrjHF/ZM
wc92K0K0Me+tJyZHTch2IkmlfXMEPn5tjMJh8tBBAHNnbsT8xnHlIfhisshIx1j5
dMCmfcYPkspSdWzNZG1ekhi7AjAu2Xx/b5pT1aapJsU1eVX/y/6b4Ut1r0r8LTxM
L8zuo4hGnJ2MpqilSAGG3ZREn7F4tUPSPxK7qT7bhod/HBYVqBdZrAJX/x8IWOPK
u/BfWHB2Herhj6unUOTUjae1wDeEhipSU7xW1m+4hkDUp46k8o/CPipWXIdzPu/Q
Q8bT2oKBUHqcHhRswrphrtscFLHwpoLjK2RaaveVjbCRQW9LR8sACXf2NqW76roP
BZb7kp7R6J0CbfyRd3kdWn3c7tmFsG7XdMlcwUix5xpqxe4SiLyhHHL+coeWzCva
X7uLeerF18dGHJg4sGWH/FpbBFHAzJlmct+lxcvh8dQyDCDaV54Hzj+UlMwHdvh4
wDIZMGFrhFvknKxGeivfxxFnQSpyQgfuRvSCXxNtjB7oUFEVO0KIxMZTeGHrg50B
iPnOGWBtl5cTI7wHJms0vNDvpJkvE4yRPi6vUu+EMBOfl48q+f4r+PncFZncvSkO
7OEY6nAYAk6FTKU2ukLHDAmWqRtK9NycUz9fiuhOJ1ZMlaw76FHjTcbwPs0tmeig
3UforIqz6S3dgCRDPSreMOiWS4oGCwKdLtqZnFNcCl9t3eFExv96YnwMOXcQNHiW
C3zg/KXZirXRje3V7Qvoruym5/yoksO6NXH2dSE3vZJRH4S6mBd8EN2syRz2VxYp
GKuSWLrF1A2x/2HLIG45kvduQSYah8nzqVxrzfETCgAhGbWIQR9VajrqyQhaMDKE
CpjtL1rHACdT6uSrsUc5Oq97ggbGaXco6wYCSJcBpHrX9pBWgNMWi8u1sy5fYaof
x44pxsnJyBvg18bgd1nZtwNdnvIFNl9fFrYMrkJUW00MXZ7YksNEwVYsngIiP4To
9H9mX7WoOAqvljIKL0n9YbdtqG8RdgzDn2L9Xh8TCNkqIWMS+j5IqCL1ySjAcFyA
IDHKYQA2sPZFesXI9PWrEz2AV0wU2Thx+ZTsENyBckY6aVFTRfH5HSSydNh9sdQn
KGrP4dS5fIJXQ7SLvJMUGdeeq/EqAyZY/Djn3S75eC3qb8mCbYbiP8ptYa9sx15q
/nUzHPr/K/Cwfn3AwdTEMXj7Ldk1OSVgEFW21v8Ns6LNt3sUpTm+604Um/eUqP/I
2XcKcjs4R5F2XBmFhWnGOMOvN4KU3KuHI1a+gUOQeFj1GpMt2U+aTjJOZxCdQ7cP
M2XKQViFBDNY5qymzlgCBZV2hdVkwoG/qZO/qGrrymgrv8z+hZuvmNwQ0H1OScm+
LPJrUBJbcu3jzsWD11uLaWXJZge3PASLmSKogxVvK8o3INAU8/H74WObruYo6de2
PvVxfg/Rk8qsi37pTtMGlbIJrprF0JRY7X7O3UKuftXkQ6D3hPQOm2AG7G/4tDGo
g7530978gTkJ/8doLaGk8uzT7aA9bTwqneXVU+XzMFWoDMxaqpCQ+slKdW7+UmPp
hh3T5HeLf73UiTsOS/DeOI9FKIB2rkagus2YprppiDfBe5qx1ypGzMaDp5DiQH3h
rFZ1oEX9+Swxq4yX5SnoP12A4gVJV9KF1WY4DoyaEAsbnwy4oMc7mc2018ZYoW1A
j3ZT/pLTMhrWH71v5m0L003EvHd32UGQ1B1ETqksX/fCy25buINkC3C2WoN8/X+O
/3767XD6ONRYjyYx8BYgnEXa/YuZRh0fNsk+PkhtN03bForyd8JKUa0+Evz6ufIh
s+aM4Q2dvCx64saQZP5Samp5BlCSRM0rsvUeyLKe3BOTF80a1aWeQPO6sCoKUGui
rrQ498GjmSUaiuzHUlFad88GVflXO0O11mq7V1TmRLBjjdHF2qHoeYzF6YiCyQEG
cReVHRI8qkyD94KJFmBrw4Uk9hRT/QAKZWg1PjrM340/dziRmboJyUIMq0JcBxuN
vb3gaXJ6CXfqu9e9Eqb7stImz2GYYqlW2DJe/C7DK0P/jErb4oyBrmwtnuWjdK/9
asnfxmQJt4Ktg5VBycsXzUQO7KR58521ExeuKuvkR61+hXDnrEtPwSNAo3PJ/LIo
pTplWLFni69FPy+6xIfE27JDWI784GESOn1NgueRrp0AsDYPFIkS+1ATBVHKhxta
OGFD2aZLK7U8/ofemvorP5GBE1tLaYHa8/taW7o/fHGCFTGeNzPSnc3FyjBqVjyD
8K9othy6kaLWPV3fVJlDzwPYoF4yBfbs1BGjnmhZNQHIPu40J2VMWGdsZzJiD8oe
2CTQPUYcPxvlWsahcN8D+BO89Nd2LTSdmz5z6LU8czdLgX4ziVF1M0jOLDM/ojX7
EQe7ktQX4csfeTd44cuWkjWsfiuyp3M9mbUztLCOuDUZaJ5MQ9X6WIvdiOm4jX9C
ZMbY25kvI5xKcCsJ/bObpRVKFHAzCmnOExn9dTFeRRDViRyWxzxiALXnHd8wcXF2
8NQXuTwjiDwTsTASy3g7pv+KoJTKBtLXIYVI2+YJLvmj8adq8Hd4mgKoi93hcN20
kkofxImIzkSfr810Yf4Apm6ymDNGgWH+Hw4c77oNsqhIndHgL4hPyo8d3aWQpuyf
w8C0df2aYk/+ztWIWnLJCGs1/p2ayOBJwON/mSIzKPL4Fm/CEDJkyk2lR/wQqEuj
VglnKbZTyJZ0hrk9cMofXlNmNTDX4OfTl/7h8onEObMwVs3SMDiVIcIB8a5z8Ag+
+uGZ9XdOHB62Z2A+6dgxzbIKSSeRXetbQbYEuakbFG/Qa0kTvLmixF3FyEmD4Yux
tY7cRZ0ttiwLISz28KVVPfQ3FJkp2bSgRsnAvoiGdeKukC6PkZuUdK/zIj9Wa11l
73ArYmULtm4q5c+5ZZEpzyizCztMZ4nN4hy8aF2pSD0FrLn48Z1wByY7U7sOhuXg
1gjAxYT9gs3TmT5qNwMYfST6hGRgdtaKqlVUmSG4LKRSwe7HMrHC/x3yxgWqU4rL
H1zXb3J+ynt+o3ex22J76+dgjhF+uEqqqpFCM5uqwjRwWXAzVZcy7GUgvf/8/jv0
laYVHeEZua1FF+Eu/7qXivzzktqbQbxNz68YqdIXwnAADy9f1hpZRFqBUGkdtPTo
Jy9JwOSSG/lyVxH/pe0lGGMcqok2j5+suVc7MYbLrIYuEY76UX2+UDD5YV+Qakz6
ghIbuhLn1jRP9YhVtD24vWDJs/T1sXVFUETCHlOL6YqLT9oIFWYjV9NGh+261hyP
mIsoNedKVDpGLIzOyDGuaOKFZhXWWkfNpmL/J5Hk8GIrnnWBaEEO0vTcigVmMbtj
l12lAhYqOVtF+2puspI7Zs28v5tRgqe53eSdSMlo4z05RdF866WVNSN5+3vaNiOD
odJ3enV5ZWJb820C2Qn5FS0QPDmxOyNjb9S5yhxeaf3zTSgrJuKIqv4X9DaPRCwD
NIZpixQf/FfKDN6xXZ3mzmKCPLK3zaAyN0u/jXEj17ygycaY1e+yqVz5iJkVPqNr
cpQ6NgeaJFJPAuWKqd+qhvQpI0Yh30hNiehfq5VPXg2sIJyWa/VHqiRMcLPQZ80B
j8LtNGYlyGUHR2/O7ysmCZSeztldUuc4+y7DR4iFL9pDWmcOl+4piCHB6TftTxdL
liz7qO+ZoYjigf0vX47OTVUJUcJqHzqODFSM7S4CRB7i2SolvcCfSEDnWfjFe3zk
cdYA+hDOJKpDcj4M08ZjUz/Fa0SQ8xcFjEBJr0yefG6CHzvkTv1WqNtNzzIvPe3c
wYhH6wzoT6IldvITftbLGJ0MV8CoO7LMjtYJzWUYshxG6yhoG+YPHlHHs5Xi/dwp
ZKqZTvi7stIcdEMKoAZTHM3itkf599t0EkVpxie+I6IKs0vTH2JIcGsEteXC2X6I
NdFXSCwx4Mun5KCxRbHN628vIiAUuZzNxJztyodCnDCyqRE6yaPnXNZ19M8bMqKz
y4RB2Yn854UmzGBxojSP675sikfH44rcdrEuaVPfphMaBIyTVWcf1N2sk0+5JrHI
qSDMHBhmvBikXnMDATPiO6v7pU73XoI4rLxEu35+xM9wPTcXPzZDb18SarPd8zv1
QQjUl/FQbZ2KP28Vja2cMLSKetv4w0a41vci3nYxxwKhNnflT/a6adhCWTlVHDDw
8g1n9GckyOmjyL+sheYJU1ecMpfKVvm/j+wh95ayYS44NHFqkRhlIreO4+0aUBNl
S13/ReOpg/thKsaoHyMN5RbJahd04koE0PWy3o6xRnguRRst6uUo2n73VNM8XlCz
rfcm/ox8Nlg+/fXksFPQpt5IhN7whf98SE0cK2rtvhJY/vyvTXP2bqPXFb/1IlSo
qV/9khnYVV+Sy4MRex+l4pocrm4SV0HtCHqiGXslHcZvuortHV2Bc/y9TOhj2y6W
eJNHbElPq0Qm/ST5/U7Thbs3eFw3INhntINWnRLQWNcCCkCmz8ksXt7ceZkEbjc0
ufyBdtWqxHIOAzcgJROijxKkr9nfyQ9gScMIlGHIifw+8dm1AFZB11hK6sl4kCcv
F2t1l6yP1q22ASYmHYvw6KnHLmzvdBnBQOkTcFVf9mZJEfLGPj/ICmjwpu17nyiN
Wq8Ppl91rAorwtwVsLiiwJwhoRiKg5NefJnYorbLUbSfZYu8FwQn7xfyrfXxL6jQ
RXwFhG4+91qSttK3DgAZzIsJpsMem7FHPBrZq44jHzE1e3FaZpw4wGUynbJXaAqf
DcNZiBwOdp7pIu45iZh0W5n7E23qMnW+LKaUXm7lG2d0PI2b9SGzkIW3KNVtSZqy
/yS2JWQk6yB2/CickmGliWPksPy7CyuxUghZFdfLmhqbAeeBJSiTX2SBt2NOF1J/
qJCMOfA3CngvXfDTXBA9ClEZC6RGXfCWZkoDVNSz7AWQ3v1dM2AgS048jCMwl3Z+
6Mv42G54k9nIOaNhRzIIXcb9rYRESPhrerAqCUO0mQqQ6TGrDTQ9Qeb25Ixwvf/j
0myhoofdxyEl74SRvVictVCBkrdzcwWZAurAN5mUklJmpBE1M5OeC6F1r/LdTivW
IwNxoBtr4LLB1iErAUrQ0V93XQb3+qT06ba8tyj3u71S4n5GyQ7WhehED3mRzrTD
Acy9bpMd+BD6mZCUAl+G1QhFXVEHOOJdZNNstecgHFvT4wcYbpMFPdSuDOV5md08
2HznuTEhGmE1q7J8dCAjMNx2ugmmkxBAO2rtqGWryw5JlLP2qxVJoENZM22Zj/WR
ZPchSvRmg4jLznhHH/utcoxd+F9wdSTKYckQsXo2ETfhKIhp7Ifq/EmOGKH4QHHA
tfW0jKQ7u7eIOzFw2uxs8jx/Fj94YIrmoTZGOauK6lVlvLnuyM9ewNAm+0CSkFUY
q85JWvDpUpo24Y7qhlaOHGSYURlvkDIWmYQs/jVMq3k23GKiJ/wWZmhr62MOo9Oz
eCITDQOAoRBkJpc/YFNBSbq/InsSOoxKddZKmIYUfYFbuo/O1nZzG0Bkx6RQ8fml
z6kTCW1A2Gl5dnAjsq8sM1haywkxSWs3fHuiG6sefBlD0CTXOuXVPo06Rct3MIrx
R7YD0QDvbMgqEzvvWA/u3v5YJJl7irbsuUSOkHVtYXcPx/VgKeEJ5xj8TqJvIe0g
2vz1x5gv5cx15GhxlMTpKuoSC3oWTyHtI1S8kZ/TkoKdyrBfJrcek3yO7FiL3ukf
uichyoHFnwfVRVoat5Jbyf8/Mv7JdLWsxYuYc349iURm82WXt4oLZDUoAIY+wGYC
eZYz6Ncff2hlqcFVVpEhoN1JgXblqwrCwzWHgpThbX7HQU2bEDDhu7yrNCYlj54z
ejRZ2mcjwWLhdVck5koOShag35fsjStwrzU9q0YaisVpU1kScPf5a2PMjj0YWP8K
88nCNet05qJRgZXwFbfWCMVLJMdwpKqPIQ9DdQAAQ0vIcUgRPiz7ESSozyZAocK0
oR1hp9jTSiMCvR7QmBA0lgxDnyKvaDBZlpfPR1uL9z6qsGojRucsvwGIIw8RGAzw
FSKNhl5AcmKUVKBxHUzJIPk6SS9NST8LDVj9qOOQt2iqm9sEZAWLNVgS8+gSduQ7
lPvODbW5VQt0j7+rKQ1nCTveea+7KtrCNco7FdQZ4l9fxa48jYD4FQ1j2jTAtxTq
OtdaoLDDc+j9GRYpCGcApznCS+06qkohq7j2Ff6J/z0IkhU1gIYL6yuwMHXIkd2c
gFGCu/+4qsGfSzIraWJyqZHBXm/CDwSL1lzdoTFFh9f7vxm/ITSsAXzac/Adc2pz
1WPlVDi/D4xlGrTnvUdbb3bVXflyPpmEGPu0PFZY8z9qDqwmgLvhzzG+LrRkX4Wa
bzFLUopFdDrtYZy9rkwB2h1iO7/kxAoP7K0Ypyp1qoUrQnK3al73h337vzW7Q6ew
e+OPRN4QsWDI0dkJ8R/gZrWGcDfLHgESmzYXTdeQpFtG6Dw2/MIyGNNVXywUX6YR
JrEfM10tdWeF3rIjh7JvKX7X1CSzcwpQMpgtbL1mOWCR4t4NARCZX27bxLbGPYge
090kwoGPyByCLcvBYZ9zpb9IRRO8V8fMsjAUbxswF5VW+B5NPk+OopRujC3pR7Dm
nhJiWLmEJ8un6PftlIXsu8ax1X6d8bvQtAuBEGMQHxNSLYOQMeXK2WYUs/JfLnvM
4Im+2GUg3f8dfcxe+xXnwdKa9MiU1LiBYZTFYr5TK6Wnirb0tKyVfmerNxtIxlzi
lERRdrdqcpYIbj4tv5BgTWS025A3x31hP+zkLCLTaIQKiuOGC2b+VppLzQj0YR/r
FZ1daFb3Q++Xa2h5E5qP8fw4FCsOOruZxAqC6Vpg9ME5+5jRrPVam3/P/0Dm7fUp
4OXDzsHo8KdANfoOmk+J4yuV0krgTIEseYXIxOBQMwTuXmlc1fUX97+0CtT7/57G
OgiDLhS8vESWCn2dBL0yW+ULDszsQB9cesV0Deubm5jp5MMs0144RJ0pu194NMN/
n6WDMKaoc2UwwuMhWfd5zQ7s3fNGd5WZnOheBGKp6hsyKzLn2bmCA0sivOQ027wg
DyJ4YBeTva++9hraep7Qh47RKZTfQSRWd6ZPltujZxzAnZMGkmz7d3ivT0B6WUfO
nwu3lW9vYLypSuyuscUmr08dZ5rMFvGPzIgzy3vttaAwCud083I9EdXZcTjDeeGI
s2PF2YOmi/zf6FkKAo3AKqGLqYW1tJxe26iMxmlldX1PY38noPLKOtSy2LwAmtN4
21KifS3dCx5bwOS/6B5vK70dZxnX08vjCusWsNy+A6B9cacw9uR/fAsqgSHgGMAO
Lu9EFhAti8nQJezCbMRwqzx7gC4HYuF33pLQYTL0uNhOquGMeTCTyJB5npA1a21m
k96ZaBW5lK0+zNQCFrwV2tgatzYgpToCRbrIDM/X1IS9hBLPWw9wjiatFdEH/5x4
TFdIUw2tvj+C7UxB5Co7dxtECPATvcfCrh1cYTVEeFa3N20L86YImrgCbUdeAOrE
/4SnxqNkOBwIlULs9g8odwjwsrv3PC2MpmXM2LKoRFk1tQv4o7T39qw422gKz5Fh
+wFlXo8NMpFgikbC02bvQgECq7PtwVJqZCCw7TFr+Mg6kYsgqhCSRbz5O/P9YTcB
6PjdY5CvFDgECwsCYwzCOzIm+5nr3Lf3UV9dO4soI4yxgXiGRlARP2DajhQ2vtWf
O+iRT9dpViXB0o2+H6SnTye06hFqLi57dQjgd/oCFBnZIkrEtqwnsHxpLdsCqwJY
iX6thtCco6CSEBfrIQ5rahx/W7Z2zbvm/Lqh/4svDirBqq6M2hH+p22rgfRWxYBP
OhEU/egGlBn+mAsd4XhH1DGQkSvZgmSzAWpM9HetlS2KbSUdnb5mNLOgCEkSJDhl
Wm1DOqyyW8KHcriaHM2SjLBTWvDPLoPaf6WwVdKmmMZpt9frXfDwSpJRzpnyDkI9
0Hjol7oj/Ao7ebLU1lMCRUY8jf/V0V0OZzochh7ZB1u7xIMfEUH4+YYC8SJjvOnW
E8XwNrnjhkTdCgIIgQKNTGCo6lO3770NMAnaQcjjPLnNntdfk+Ry9Hs94jGSRo4z
8nka28I6/jO8X0FHKPm5t2hAgkvbOXjtzOOrmpaC9tBc24lR+kotFv249xTVYlh4
oJ9IwNu51aQBfqD2NyP1504hQ/98fgNhi39sJYMPQL+3+phxoU70F2zCLLlNO3ex
5Jf6b5W59w5Rk9vLFW29HXDZx9IdX5mk+QMtvjFGePW/mH1HJM0wtdETr/ni08zk
9a9KvxKzH7fAQ0AjRr8MdEAR+NI/oep6AtC9/CB2PLwIapx6z5ZCNkQQBJ/aAK1q
du3038+Yvf2epCrHjLrayoPC522WCP5G1eNu2QyuVvfaxvM4WqCIxuZdPVRoiGDm
flCTRHAYy+/v40rhkmW6eUDFJ4UKNthvGQ9ebkfw3uIEloRZkNu2QkBKcQHJYntJ
XtF5rSohPQw50wq1wpHSSAxNSnOmMiLZ5r8pbgHxS8WKu1xFzMInQqF5d7JPGTr5
3lfeFO3K6wZluDbAMHw/UqAWLKFooIH4+U7eTupSmSMORjObYYUeYstSWOUlaciR
fP7n7N1BdC2dfsIZ//1gS9NAe5eptZCYHVl0hoQF8Q+DPr3moMs5JxFrVK1lXfcS
vpxmnWGH4vrVg1V5I7CRcm7Ift6P3grk5NTpCFShSmo4blWW7G6RG5ZKqCS6uRWV
xYAek+b/6HupstaWYyw6IS2rJiF4HMMHztf3GZbCvcDZi1e4UZguGesU7oV828U2
GUErrW0FcQ2dHqKqJeM4NnFlx+Or7IXt3oNKoiabJTyWU0R3JLYzhJvDJLVdndHs
oEj6mecgB7aJIVXghEY2CCjv5pKtDZ/Gv+PvWjmjp6lO+zoOaypf0wfMuaAUC1PB
W8dO7lJ9dt04eTaZ1LCU+Xw1h6ZoCafSSYisWvuHocmhhEQB37JBI3OQfEJP7Wbg
3HKGbr2VdCw6NacyVjp3aKMuvEUyEzQAk2E5HV840acSegY8Y5vSuCFYltHhK6Hb
5IUlmMINjNOoYk3Ub/MZd7rDY2MobajwC5CVCO8z48xlmp617wevTDJLe0HXtdkK
no1s3q4lLLOecd/LudD3MlXJBzxjwz8nnEmP/DyhCu2ULLsdzPEmK+G5deqthqrZ
2DbG2Q9N4q1Sjg/8wZGPPBDJNH+V3fCb0dxjExnqB+q+BIU/g78sKvvG4QaW0fkM
QDaPdE4TxRIPBv44qCoOZr1BzQ8ZeCa4lv9lUoXs5hKobY3/QAi24PTMnOHcNJrq
1ZM0N4Qe5HKvsJX5XOr+Jp3uKv+0imwxuUeUm8ofxvYo3yC1XjRmX1xR3FcsyyBU
tTr2HBkLABXG8ls1fbWRFZ2win2pcOOCmZP4Ev21WZCm1ygrqrRnbZSoXTIsYhbl
LpyZu7LRKIkLjagnxIgabBYsY6SrmTHKUTx0+o8d41ckdmGP3sBs47XUNUNSGwOG
v1Kuz0g5nvrNM56/tihkIE9okFuuxVlNzw4/12gzAYS/TldsWa5Kgq7f7pKeXZNz
j+P2iQ+LJqo2I/vWHj0eVuu5uFh5OZ9HpdaP9DKGpdrzKBpQszaOyUPpWIWjeQnw
noA8NLppHAh3JovJ5Lx7bUhc2i5mxD3DUdcW9cGk2pGk6Sb56Q5Xoy7yDQjiEssa
2GOv1vIShxvzzPj0QX3Di29jmvvipmz3aZmVNADb4ewYY6DoskA5ikB15ybIB/Qn
A5iAhCMLQdPiWDxNH9naEL4DtCqYBHACIvPqAjKsDHMqkCGWOcEy2Tqi+7b/enWq
6Mr9jomz2yoSmC097GMrHBQPWHuQ+JP9Vpftypu7fHn8Gh9cTj3J+N0peaAXeqXN
xKQIvYymfHY9G6au+BHPsesoNu7eYyKq116lPRGhsC8HqEgM7eLZxL2JVYtig/Hd
rhXyipaprTpnUgOOshDRFZE5ut1V/mbpt2TPpZLEVoWt+DL0TjpSZ3Pk+fOsikSH
P0Q/FFvRUfYUcUOuZOwrHeYN1GPNQ5HZQdajy6XFa8ikhx7R68DiTsTVEGhtR+lr
bT72J+Ce+aawcEtCIXL2FHzO2Fme5DLGmN2XzNyXOb9EIuioN0WxPLG99idJ+9mT
3emRZXyOHIuwkXOHq9WHj0p9i2cCdfHggqq9UDCf7XPx1BUlR+Nmz3a4c7NYBkAj
+Doqv8Efa00LTCSsfxxMNVLwaabdXxvKi4qHTzya51Eb82pG1E+RCn1FbBHM65+g
I5Pvb/Xhmp1uxMeSw8mLHLZS5yFl2yhN9x+4uiilE7pzrtVfk5c+NDid0WOgjChk
WOM5VX2P7NE4TKTmjg/od0jZRngwbtfkJBc6ff9Fh1YSBARb1BPRKCZCrn9Ju228
JQOc6sk44ndaMiPMVDOIsxjDSD3FUSo6ztIb7C7qLNKQmUUCDp49GEeoDjaArDuf
8IChFdKX+erpfkxnlVDS+2OMhPfvci0ne3ZIjxXk1XpaZUSrp/r1aILHnM8ej043
3bjODkPLve2Yp1BBXQG8RBgXNZQE8ImRezC5IiMfco8cSZoX3eK0xTiZK7MayIzk
vPk3EPIfAYZM1OFom9dTWSD6qXaIbqVGWG5hSj74Htc8cGoGaadiNEUvv3af9CxX
Cj64bkJhoto3uikp9Lc6TCXKeLZ/3Jb/d4TmcHuDhA8K/lUTFjyCk6vwJIXWhqRX
mO5PCMbgFHF/Leqs9/SNkzzJhAa5YgWeaLcm6Mxlcxt6jCQO+sFmGksGYqW5S6dH
o8IZJMu0fjDN2qYkEMjgJZUIa+SB+w39r/Vbuf6ArWLfz1I/an2YX6QOcGvr/hck
BSwFcRzefNDWjnrdRf5ev4FrfdYwOYv6D6y+b2k3feTBtoXPGjE7ipxtsyi+9gic
m7s3P2uwACQBokJW4j8cbqjSScBBl0FGDjrKx5hD5KUwqx0J0JzNkZZ6Hl5p4UYV
Tu32ysdubZzNcltgPOdYo0guB7U8OC7mrd6cN4tQ6sjwrys0VSv3b097zUvuoGkt
nT2VUjgBt1nlmKVwsCuxOv2483VdjuQlNN6cFpMhQzR18TcwFpjI8qqxQYOhF1s4
XeJ4kqppakJ4Ck2IYt7TxEvhwLPZalX8/ysYBXG1vIvvk56tfoM1VFFY8L5gPwyV
EezB/BPop+ylU1z+3Nkl3HmQ7g+mZYCLox1mGJkBOjNC3lKY0nlWiPFyRiKCv01V
j7ixg4x3OtAPFZ5wDLfojXqg1ZCNQvrFqwM7DByx9g4GdxvfyUxXWfCHRKA0TXOG
K9iIcXXPUTla8tIRpJZ0o227xDQUj9aaJKXrCnlOvEU8ur4XaZ96ntInOUVOUB5O
KEJIwoLaXYcaGDoDh/VgnvTWYa1CI+KcfzxLjTvHKs/Z7VQwmytT3NNz6ECGFpr7
jWxgIpexMlMueUqtjQW0Tzj8QUfy4dyW3VTmLxZ4Gl3zin58Zy/7AsU5Am/yT8xq
4+KJcRwvkPQ30CuNJF7TyYu7IQI2mhOegxsYtjt1G9moXweVMpglvMX0nRFjSQGD
Knk4NJHXIFuYcgVRfP19gPm5EL4fMOzotvJJ+W9XSsP8qyadrTYo+Y80QyMToQUI
dEYzrCCDxCyXWD0OG/Fvl55Aq6ZCVikeNdu4ve9bH3fZ6Uk13CNexWq5dnzZKV4D
newHpNd5thtWx7q1Y9mSeo5q3yK25J1Imcue1UPBP/jIOJqDny9DJ6zK5Y1DR3EC
v16v8mSbdZIW4oidAplmedbIggj6LWzdYjFVNajmuOtmqxKRrzrCIcJ06fdszS1O
dY0KQMp+RoPJ1lOQowYZWwvR2Nu/dIOSZlZRxUoxjHnNsfBbnjq37DQIQMxWMAr4
OWXvDFnLA2NwINEvTgrAkLvnYkiHM0xLgBbSeLNPgSCT/pT7ITgDLQWCm+pTQz6y
/VTjMm4f9bCdmwqOz8a6KdsUFefFAm2lpK5r7dxP8mCBWA/6R5WfKCxqJx8u1zd6
VH9MDhM3lR+Muf5LOI3kJ40iCAa4ZpUg4QQb+Ygh9fZBaKKTnW9isLXO32LbFKEI
13HmYC8jXtwk1uto/AFonksHY6bJXubfSY3wC8/sGlB3ENu8wHv2FRuS5Qt9Cukf
knG+wHWo+N2/qVca2wzE93bTzUXvKJFGLK/AFLMvCKt/6F+l7DcMVotu7oNSQOcV
esjkJ03MYVEo5hGkFz/CmAects0Mso0/oQUgltamrLp1tehXU4KndIUlmXk3rt0I
Vsyn0EqV3POUQ/lzt0GoUwKEqFo+Ub2wJSZnlBOxQq9lwaqUyOusCrJG6ezXS/vl
qDBxJtnAwTRzx2VAhNW6J9VG0rEoYTfGxMcd5iD/QIY/5qoGGfvWH/gYC+6Dk0Ar
VZqk24jJ8fZY8DfM/i15VZSyLfT/NeMwbzed6tq7BPc9DXyTyldWL+nuJvTrP84Q
dTzxASnz9ZZKpWxKvEtnQcIqhqPInpjcKFU8MNC565TpLBeSh/NvivuN7GyHNzWI
I9WNgH/XwDtm0x+mED7ts0Kc0jkKasdpbRwKt91Y0Ljjvn59LZlWBhuBgH5HyQ6e
XdWXFX+h5AdW7CjOV26vrdBVtMnv3lxb0/MNPD+olNO1Mmxq0SmiF5WhkejbusVg
roiLax7BR7T6tQEf74vxZn+VnD3JRBkG7rGiBDKvlbT53Wen6J7rVkrv6xcRU9PB
cQn2LHAUhJfP6ZgLd3KnoQfYEky4At4jk/JVoa7EqY1cyxdIhAZ5Yoj+p53nXyVM
bjyT5DgCTSNSkzVkayc9VT0PGnoGvxvpznF7GbP3o6SsyJZdlLCq7aYNJkOuTbPL
axikCcwWp7mVPz65v530h545ghS6e996ew6ZON7CArheIYN07f9Ak+S5qUXmVIB+
SnWQS3Cah7RRg2Fku+keK7jY3xX0Euo0LsrPlVGeF04eAO3wO+mfvFpPPoCCci1L
Tb4pMj8I5EKWZHFQFTLCPZ+H58vhN3Kn69R1IFlNnD78FEHKTzkdqvHwwbpHZm3r
vokKj9yUBrxLiQ+0/yFrYbGhW4AmbwO/kwX4vsp7BMcNYCEvLa6TpckfHoY9z/8H
gv9KsBbz6EFuMmA0wqOMTUm1YZdNfg5ILqQIQ0zRxwKZH3Q/mUhU3SNvWwfQShLN
7BG1cRTmrXChcS/BS75GZxM8IU0D2QMsNRsa77jUnVUXEv2gSDSuQ5ngJtMGkqrm
9Tu9nPJ8sTblxOXGXw/UeR/7hC3NJhzly3BUl0qDuhJS3yHXsuJ7y5Bix9WnUR/X
B1+df3gEiTRWtflXMNJr+n2jf1nBOBntT+XY0jPurLEprRN5UeY81aL7YnO3JKRs
MNlJWJBLRVpLGaITMd+eWlkIW7x5ljZ1VMwinpGhjlG+5leA27iSveMkABr0Zkrx
W8t1R9NGy0AY/FmdGQdKgcqmd6R2GaI48J2rdagXZvAeU7zOzwYHNQQQ9GQ/3Wao
XWLJJKH8lCdbDga0ZHE0+T93wr5knnFZZH8LeAxiJdiHL53b0KXG6nRYiW3ZINvl
fUlA3ohBQoMGpuYgqcnXFtSFhWALyk+9TgJHpWLHEjEd9Z06thHV4mUCfpHHXhnM
on+OCiB46dhWXvLF+ima2cP5h28Anad9gRzW9HivUlOqW8I+hOujnCCdNRgu87kn
yS8uIJwyMPXLHDSdfZkGMsVBdvXhJKwEEYaiX7Fzg6emFUlkk1SCPtU069ndRwGh
7VsfbyKaGhArPRBwyEbl+ppunP4PxHLiima8LIOh4tcdC/4wtXA9x4RvXQIwFcfH
ov0OS6AzTXgWSYYsMvXzD7FGl6HuqPE7BMatKNoNF6anFFXRymruRJiR3GWGDSMe
tln9rbJimobzIXLp+trz63n92KRxl9DDMwZpcq8kUn9DG9m10jsEP8pU25wuYHvs
xWw279XGQrFzxSfR74XgUSBRJon0JgBOimxZksGZu9NlF9/ku3FzTM+TTw1wrRaP
58ppND1XItJXRG6PfsdJwX+y6UNxMNCKpjdpTDcn/e4IpIQvMCHS9DzgCbkF99Sh
jGJy9ompNgkA8KdWPPrfCb6B0Xt02al38oblvTSk4KWvg5GjsGaxZISNIsgMsonn
yVBZelfkNEl0jAv+PblKxbxu4t+hDMRfOX07Z1fSRJBjmbZ2c2wTXfoqd71gBp+V
znMqGOdrCedU02KMWO66kE3V10EE6xcAl9EDxVr/rMPRQgyAkWkt6QPtZpbHotaL
mmkm+3aMmV+VXBHgcqX4xkxsjj+vbOrqZoiWfx32KIcBPC3Hk71vNf7FOc2wy8oV
mybRhRBDTAcLlxzD+UU2WgmbmHdJBJL2V+/Kwos7Vc07KzPrISBHiBDD0zWufYwt
F1kiTR7xhp8jnGD3k/7iEZStREvRI7xRpyjfip4dAQXYZrHh7VA/pNiISVWs7pZa
gDn+45xkwlG6qKou2FGgu7D95GarGGonlFY2xIyVTBUoIok76dizVvfvey0nuC0e
ycHNi2Mvotx4JYw5/8r9SjL11Pv/ED1Rwm/RV93qQNRnt6KCxTrGPvgOor5vQq3R
GpYzdJTkM370HhYuqSH3+ZVtqHEQHT95wQ/XMKEFyOTnenABaawQCfB3Cmd7bVBL
0KMas5W+ThtEBzM5OdcvaYz2w/i/K/1Ct1oBc1IwJS6Absa6vgZZipuD61rZwR0d
aj6c/Wqb5MQG2lh4g6geFVxSAXJj1+Y4GEVR1317eYZxxK3aLYGQO37vE2BvOHe6
cmkRRKeUfNlPVGCjQOLU1IWDEGMpq4+2qfZqsg9MA1xz9DSuQOB9yvsGSlcviYIK
B5a7Dz5+WDT9e00KEG9WFK9vYWXJQgphscoXDaINl1EIuKipk1Fy1iejLalarvnB
tIzIdwiS8+73QSpD2KVeU45yggW9s/d+JTT159qOxzMV7tr7Q/ETL4Hth2/dMm/J
xVnpvWGSGsAimkCUaNe7cCC4IeUvYTQAkeakSXg93MI321/iJiG+bSATHu+C/1WV
3EL3VuuoH1fMVKiWOaPVA7ZfYoYBvq7D1EFqSr1plXqeIDtInN9ONDCwyb+bI72d
Qn6rfNZJ0yiQ8dc/a4XElfqPhombNjbXOU03IEDccSAB6vs8G0ShqBlLlU8EKSZn
b+GJORLojUQsNGVvjElD5aIQc8GaelFD1Ov8D2HxCzUKj0SXboUxJvuVft1+B6lp
tY9YcH4lroa5GftMuA9c3R8VyhOjZQXsIXAOga7KdmlPA8OfrN9QL5pd+M/c70cZ
xGgqmHv6UsrgPEUrh6bNqMp4LNic6yXnysVeaK2coq8WE1WxQsj6r9SpHKJLOk1w
DkGsVFIWBAxCHK1YJeNJmpRz0FFHe1LmEzLFg4KX00ENf4YLlpOESNBCV+7QFu7l
6gpPfU279dSL8HBP8cPZnb8DnEfL8jMAVyJRAH9oH1B2w9rqTBK/D3dF1l9aaG46
I4aFOVwVZH7GzGkZkFuqA/XC7CwkD5jhyL7KfiX4sVJjMzUwziawquGeMfnYFDsE
QQLiXpopX4LimO+0Gya45CZvXqy4ieBefeVDPYewWkzo21IH/LEsBgEvTlYVZk8Z
gVrPB0ZvBdtfXcrjT+WZj6uLt121+y2mnahprPx1Qxue4Gv3HJntwY2WbVrcEFys
wGknZ7MCukEV7dwcBZFYbhD23P+IH6pFzLKRTu2/ATw4S69qZ31KcrbmvSdE8xFe
bRLBEDBcb/4gmzFuh4aafICs3pUclBsaxwJSySnK1w59IXfXSX2asC4MXruWceUd
70xvPja1u0ie1yFh3WIYcYOXsnGll0SrTkwH0nOC7naX14MM6RZBA8jU3j1lOhT0
20acYgsfWomH26EG6W0byIKDcSklCcmBV222blHdMapBcwW80RpDSV68fFSY92aR
HMMwscN9kvNk/aqOTK4w6J/zNhRVnFwIEkQ8VFFhW1lO5ufawMioDP9PeXCi9IsM
LNbQ3QFuBfKetcPQcfSQDZ9YYSan1sP7KcmvD/EZJAhoQYYuFB3MlD6ct/0fgIpl
3p75zFNflYFj52rGl869caEOHgPl2BaMip/ae5dwXTDKVQX8igatdCpprai7HtaW
XLa0JBnXAmRpS2+50LfcLrN3TFSWr6aNwHNh0k1qvgN5gD+O3JhzpQ/xQycOWx0s
ZOnri7Q/HqSvUMZaTsb3a/4kEjg3h6KhpD25cI1SWApWoGyiOvm7DxA9L4eO19Ks
E5vaBd92bpprrzzZsK9IG9igd4/EKWp9sP4EKTuWIHdnR5xTGI1XaB6RWAyMnMQ1
xGAhSmSMiBsMlDodvrQN2jWdjwMdaKe2i27zDq77i++TYUs1ahnzCxuMkrjUZy1V
tNuJHNo0MjPhEz7GX2utsgM9PzBGXdFfDMnupFztnZjLVjyANQ8u5wdxp8z02cNV
oAHB2ARtnDxp7LKxgI7oTZoltyrtO0no070zZhLpBtGCi1pRukUxz6y2wdKmG6w0
95BRbGReK+9SvRvLqw7B/FcwjuvPPDzu2YbagCQ3sHCC9RhoytA8AFTpbRAPxrrb
ze5bFo3yg70Ul/3v8jb2C04JLtbG9WeXOXKnh/jBVMQR+uXgUM937jw3aR+Vk9Rz
xB6xkJHjqy4byZ1NsyVuVoqikmNJ9sOWgi5jFj8j/BP7APYCO/vytOO//8WoqChg
9M3vg4kcASLsAvwI3ztHzSvWs9u8oTs47ajrvWUHcZRGBlX1Qi6xD3oqA/OOZ2So
fu4zYlkJu/zcg3ViGwP811s6lJGOOGYO7cf4qGw/pKSRgnMeLKaO/PUbdhVf1xhk
IxelXkMkZCWWZgveVl4j/hC9mSlTXzmzdN8bjjSMfr/z3CwBc0QmAjlLOr2X9q6s
om71jA1QaDB1O0PayfcUVsqeVt1Cd8rzblsRtiKlMP1gHLx36GqRkvsdZydfHbfV
c99sb7xntFbQ5AtwQHULiLEMC0JFgi1noHIBFgiAXt3JaHESsp3AffR4yCH7xqot
4nsu/4H7wdHzyXxge5EHKzd0kgCctIuyMKw+f+zBW2UeLfPtTje+x3ZZWDmWS0oU
AodhV84SLfXb4DuqBOSETQHvuMg2ZCOrU8cQscu9AWxJ5h7Q+tfyX3wZXSmedbka
Q6HmfbTRGBcZuaUw+aNDe/NGLtIUyNIzpza3QkxNkdlg0VVdmbFkI7+vIGPMienz
XOL1mmprWcSXwvLbABVyCLaTqGS1ZT6IcBIb56RZdq3X1TVopeUqKH29PdXx+pIK
mjggx/8WyLYTMlPWZAL/53mCwzrW2jxLxEd1cfNdgSLuoaX4kqyb8YW0ecTbwEW3
CEkh7eW0pE+ALWQAGBRtJVoFkLDMPTk4M2lImc5fCCcYIBK4WszFsSgvTJy/Oz16
c/Luz7gUaZJif7m4x2r8d59aB2icXRFNxo3Lt6psNIhn7RNEtu/LlKClMnu+9xjg
QzoXdpxJhL0QVHstKOE9SReqhluQwzkWqSiu0TZeE6Twq6NrpDWAPp2ZxnBTJxKU
V2lZGT5zfO9yRCL6xPvk1WdMmuYy1OyQQUsBfprQGN9z2jF4XK6yCOmpmkHshxYq
b9hBPeElqvywgdzpt7AuYmDWahYys55O7lOjwZEZ8xoG/DtTFAlNShrlGmtai4P0
LR4LLID7oTAAqour5mKu+U2HvipsT9HThufulagzugFEC7uPTu70OL8VeA1NDDNv
yPLfmRZ3yoyn3RA0DvkoUq1stqn1j72HHxoQd9AFHkvVZvZsOu0z+fQPb3JvfgAb
E1jsRvEuQacFBUeKa706RowMrklR3rGZEq6cJGuQiXXp40M1XhT+m5tjGZ5cqlI5
Kt+rDWKkPTSBeKktRMuHls6E5mG3VXArk/3EwXoyHn0ztpuQTeroJtm+/rYaNqJJ
meEL54FEyWgQr3jUqiX2LZKm6OWtcgG6Pr7sJozrl1N5//Id7UXSavBPyyOs5buk
x7BXtlOZeDcKtH5RcOXWEZQwOhX/q9yK0BQUHTQ4mcFweVy4BHPVp2xomZZmye/O
QSoxD5ETct9G2rX4545J8eXOoutRdHEwlZ22HK14N2iPWWEvWjCHOg1ugsmA7Eyj
eeSArZZJSOT8Zzf5CqY+fX34jAobm27RBA6ZC04CmKsa1qW70oiszFoURkEiblzl
sq8657iwTK5Er4qZ8xNtIuXDbO2YKsC9nWxOrKoF1um5rFahO2k+XEsTJAaITih3
7ZDYbzvz3V/V/rquNO8+noVjzB6NKfZgIWuBc5F7y/RvjS8mjzgJtrC0LyGIzWCM
9I6cwh8BQ0dcHRhpw9IVNo/Hxf2YRE2wb+STDz7lq1MyF5BRmXYjOBAzJIAhVgKq
NKo1GvQ1rIgSp95tj+mSA5AmkSRfiP/dZS22lRWSZOnt22BTORimZxZP2HiqlPpm
XjA7C5jEVHHPU+zqh+f6X+pvg3Mhh44LazXorCl4PHfIaPtkOO4u0cL93DKQPuvM
b7C4fwoJxeNcfaC4teLj5babKm1TnLDw+3lK7pWttJJpLqXFnKc30d9cN4/eBkg7
43s325GRye9E1Jg3VRfoIoYE4ZGm0PpvpVnVUoXC9n5AyIsoryGtbLLV2atxWq0R
49560x3Fsafao5iFpSRHIdJeXv5fZE43Smkz9G8x9LZ5414kRPD4aP+PNh6UgQGu
P25hioo0yY57yiC1PMx0Z0ZxnKuZq9wnEp/InUSYjAci/krQPXtKiZKYl85XeOmw
qGR7+le+pJ7DhKxQbHUy7ak1ym/XYkOuiuXUy9x1iZ0g7cX0yTzVVzBhz+HsRyZN
x12EMF53gq34b83mNITlhMwA5CigfJGcjOT9JtRu46aKQY4Igk0TphMWl/lwVL/1
rTquW2kMQ9PYTX6/tXyAaHjXQgugwLcKLNq9sp2PtdmN03P/YaM224kB3L5e96i+
oLlhwuBwdS9nkN5xMK552AumTze1szXuqk2s6AQX6f6NRkJ5a0fahvNbNs2iyTBm
/pp8UBUudbxW7F60uFFMYP6zj4IQUVGTS1hfc1hE/HZV1t7AyeFztNfgcMagyhYu
/ELNjngvCEx6JMb8ZMbVY/LT4R+go1m+PeXACtoMMhbIwN7T7xEe5JxKInJ+AmDj
G1bgEHcuX47u9CTwMTyTDN1tHB8kEs8aGQU31LQjcm4nxqnGHY9xKERysWPCU2l0
3KMwlhc2qfCEx3DDuwoYHcw7sHmOSCE63ySybetb2EIw7wFaOOvITiqPzPDXwrHq
tvYkIsoSjp2M34BTaDYfotSQq/BDQuGZiJfQ1jc1ypWywwIQq4hlC7EEitYfuwzi
IlZTZIePX3hDi9gKQ7Jb22Dl+ZGvs4cQZBKp5yUi9hUh3+4yrNvuYRCrXIpdQaD5
+3R8kL05Is7UNenIeWkpW4ubqOr8Awc3Y9BEt0vLKqcujFGRs5BZ/yk81VFs8aIR
uGRCssOWfbtIXnd1BAjyYBlYJe5cDJ4d/Eqv/5oB3ZRu7R+QE71M2OqLoFgaLa8o
LjwqaRWXlPNZeHEcCODn7wDViDUuBz0La1JnqxdbMA+wgH5RnURm6kudHyVMfIa+
d7L/aURVhOFhfflQcmiULD9oDo17aA710tfADXCs08itb8fjJ5+2Ez9gRAO0Freq
cDf2n6wPgF6HjxlyUjqDE1Qmwjd40snEf1DuSS3lr5j2c072ZuRct2KDnEYs36BS
3rxl+H3E4EnjdIhpP5GH7tAI0Tbrv3QlvMxmEilRFscitABMVreCOjL03/jDPddg
mmZpd8bRWpmH+xxOYtnUYlTWo8nwTPQVvGb35BfvNoqq7kDrBlymzsbOlRWZh1tG
qfHsRTNj4n1BQjWRVWzfJGJkpvXyb2lsaNBKwm1eDTddJiJxvYRU6ELj5ssWZePd
2+GkMZuqAdEfFUVE8tJe2puuBGBEAznG0wyQoIF+BY1EinDYGAntHRhvSZm8DwLn
fck3Cql/L+q1JV8l/UEQV2SK1eu8hbhDpnRAPZga4UzaEQ/xYt5IFdDz4r9M4yJa
vw9apOsrJqM5vxo/j9S+ZoCsGIypsvMrh7qib59+OJ1IgfcGp6ZGeYBJzmp73eWP
vBvj7MariC9u1DkRIruV+8/ysTZQvEcBwcGM27UJZDRWrHZZ+kq7dji6mqF7BlbP
Nj3hYnOVqvywkc8lxihjWygdRdsiHF+3ID+mbpL4an2eq7ov1tcnzMuyOry5CgrR
PCh+yDA59pDVaeA+gRosvsW+S8y9b81XgK4RS/Sbp69EgSt4MOBiS3sMaYbec4ZB
aRiH1/Z2qbM/2JSZDfurqx9NZxnFDPuyvT3amoI4WTtkPDuKD4HnCoIl0A2VOAx1
cQu/hzdlR4syC7vhuu1CNlZFUQ8CMGTFk14ff55InUuYHYfVN2rrvsognmF4bzM4
K05m9WtqQvKktRfiRnu3plK6cwlL8IIg8Jrid9zl6GqGFkFqY9c6SQtpn+RZplXN
fLRLyhQsCQy7Bf/ROLlEsPeoPK17Osm2eYO2m2OXuMMfOtHcz0e9MDSnRJaphs5H
PEBNIwMpwwnxOJoOhGIyZ+niU8o4Sp/T7AQUdRZnTMr+fITogzNvPFwl7oArgNW8
aoFozxjHex3rKSbaeSonQ2SxG0Hum9h2OZqTzewzT3+rpUgZFamR3K/Id/ho8uuC
GzFtFovpWJ0sy5KNPD2IakcWMeqB47aTI6CzVQZkvo5jA109eW67bLyR9uiuMa8u
HeZpUzUC6SkxtZdA94Vi3KEEijeRNnSY1vQg3xNYamGdkiodwoC4k1cUTtIpYMJS
6UQHSHwQBS3GdhwNp7xjpfhMOV46b3cgh4AOEHmWK6XUKaUZO7hVr5GOx2LHkqbN
CyJF2xbKX/ARBUpYR9MKSx3m8BKHc57+SXd6atg2/X3tjUdHzy4qTPR4KrzghmjF
41DQQjzLNJ5HOePCpTgKU0dQNsIg6Dlz7ZUehyUffCHfE14sSggE5hYC9Ajun4lm
l4ecVq4hN2E0IAzlhG2AdzpVCsOVbWvoUxONGikTIuyyHiQ4wws8KZzRYhSz1Ulh
MC/UqJPvUJuKNNJXt+gLH/lMblRQ7LJupXeq07JVZkXKD/hSlMGAzLwlA4dBcIwJ
me/lHyDtQBazqfqM1UFiNNs6ch+5M5F6y9GwWpmikkwwfYIQbqA0kP5jdCsd1DoI
nQxwHWV2R+dXtAH9Py7KrPbC3w9/CPxYghlqmNQG2WeZ7Q+CiVwtaLy437lfQCWQ
L6vl4uR+ZZeeY4qMJp36zAVB3GpLtih9fT8GFuxteiGCgQvw7hO2r9YbaDvLpoU1
bfy3PeX004pz6wfYlDKuNCti9Hq9igycO5im+ClMADgyzdjPKHfLvg872RBCUrFu
Oyf5dagHygGsLE68MOWHM2i3LPR0nIQS6BTz6nvze0HzBBSELjijwT9+gTC33ZqD
p6i6Xham8FGGnEC2ylKzF96ITRYGyP898WaSKQBsqu6vQS2feSwuJezPLCIHsq1w
rd6Satf+rcPsJxMylX9QzYWRGvzDE2/jqomcZixsXzRqvd6tDTgGHHBGR+LlAGzp
y6SVGn7DlMS0kEeCIXwilk/QEMy7A4Xy9/do3l+WXiNszfRP6o2VwOGBp7RpoIp4
m0cctgswYYTB+uN9HRuL5/rjUnCVznKRBO9HAdEUPmFhdFTYzzPECd7ser//cNOI
AH8HgI1sFXa422zHoHm5l/3tSD5xRFHnVCM8iNsE1iqXEONXkZXHw7K0JL57NWeD
D9nTZzRFqEno9ytCY5K1P/1yHx8anPmET/wRD9JydBCvrZN7mc/oULOscGnpdQOI
9fEkq976zBE494xlNC5QzqIMxfSQdpfKvJm/UcTlnZ4vebKuIrQe58jdQ3cE5Q5t
PbW8pk/n4Kb8RFSHKaKdYt8CtwuIHW53OR1QyFfxD48oFvWz3/m7ZCydXN35xjR9
LuIB/FpYxm4xIJuhws8e+w/ldplA7NaMItRTKG3Yjc4RRRiB6eGm9CjEvBPJjd4N
eLS8mQRcuw3qv4cGc3nWiMNDKy1LWVM9PjpcCnM9cl6eeV3rSk9WjzZPLjxVIXYV
ocuE3HnUuYzMS+iymfrCzDOFd2RhKlUueI6e0taJuQJOda+ca1S2B3+wOounEr4q
/idFm0J+6QMBl5c4j4qmMqwkxA+TUTD+gLKp9LHdZfnFfcPyD8EnuRsoRa2OFxHu
9becAZ/lOghrXJuRWvoiNiPm2jd4zgHnI5LUaQOgpVjbwsT/pAlDleZeU9iDc55r
+b+60ZLs7DzSixoPK3a+/wtguwh+B/TBV+8nY86bwhUg+lypfWbMI2dTdDcFMfrE
ZXTBrm5grLE+m0BNU6xwzQCLzoEja4Uf+sm1+CKCwM1ukn58zFCtotw6Fh4h0qgC
XYTRhA8I8ECDDuhQYrXH0xrXvP3BIbJzxFUONkktyx1EUvmA9uhJLVgIuRgBLUS/
rYjVOejjl6IAvITqQdG0loo2ukNlYFQNz51VlPdkSxc7g2NmP3mGvFETsOJe+7i4
B/7+SSDG+emtmVB3hK5BmHNSUkw82T1fwJn9IyNLNd/9k52P6Ajl6pwl+JS+YC7w
YS/WixedKkrPHOzoXakFL4l5MllcEvjlThkyd4FDPs99bAMB5GUE6UJWBtfOUiS7
2ZrAc9x1dE7JlW2Ors76VTh2ykK3jizaC2ybZ8xQLz8logs1Bi6AYD59z+Jt+poL
9AdTdcHlmlOBZGHILL0A6MMRxdUX/pcvkEIqiWmjsSO5PjGtUZbVn9DpBtLFjyiY
Ii5KjKgfdob/ZzOajGxwUkDzA0sOfJ3h9fy2wWb9HJwFOHVzEebG8DICPSOs2ExP
py7YzA88D+f4GIDrTE962Uj6uRcGWDWyiW/lo/FR8HP2930rRzqPpbUs5R91po1+
CMWvRTEsxfZjvilfqff6OkteMkWITQ4xD6sBpXNVOAAmCkMnxhcE0Len5l86O2tC
GW4Au8hNEE8/c67eZd+IP5REFUnU9u1oMvmWPoh+UF2KGtja509YA8pXFAFR9CvY
5pd5pLGTeZ2gnPf8pal2+VZWiOLXuVXwNUi5SIw9vAv0c9xowpqMyLUVqRvX7F/8
5YWpljmeT1FWIY3kfBPDlT56WC+L2CPTD81bfLCGcsTiWd/a7jjr9IwWUYjNNi3a
zqf5h51yLe/6CVb80dbVj0BBeNCZS//3EPCkR6P+dwXtc95Z3K7J4mx8Yu3F3rEi
FECjBYws9gIKmox6ucCPQ39TrCU2MRiV5XWce8fDyJQmmoFAmIQVbboBfZH6auPp
j2BEx/3H2B2Y69nrLu1ANEOnKPvYoqeMRvkWfagF4rmyvSkndBkmqe5HbPo+EC0n
MXo7SoZ6lYJiP7YcOnPjvIVI+LAVXUKxSzozliMD7Y1cKyTYtvEq0JopWpeasNCp
RobtOiQ1Dah5kljBnHSE7w3EPvfT+z0tsudjAUxhaoVSSWj+vIwT/lJ20k7fZdtG
yq9ymnL8fS92MTVoZR7jQzpBbmagtaazqkzZUl1vzy5TK7gHUBYQEgZvTPja4sOX
a2YlgtC0C5SwdJOiUg42MOl1/oI2p7BaNWbs/Oc30eO532+3NVfSbC6X1kXD1VCY
TuArNlTfMgDZ/Y8aEqlqnR34jH6Ow/xZsFyvOfKOzpeTFMIsT+TBu2aQZVPLDqba
PEBPOXQ3JsY2U0XJi/bOq7/b9nyEd3eld/W8vmZ4Z204kTNclAHl/n6pZJG0E1UO
LzA3xRN6GUva9Z4rFX3LpsumvXC+ZDZ6JSQwLD3gZsyJRrqLyVJwEp3sVtB/iG6F
+CywpH+By+/n/3RQsA16dBsMmiiCN7/Zw4EyboWGAg6l3NxxZZPVyAMmIVEETL8U
/cuXLOMxSumQungQl6o2R6GdC22oLMVJyZj5OiSYLowWFVcArK2VkH7RRCNLyhbn
+yug2ZHnxVBlOWxvJbHOHoJr0SANYDpkfXJVmwJNoyoFjvgHfikbk38licExbU7Y
4Jr0QzateF9I5KOpogQNFJLsh8P/FLU24WNhvlRV3ODNB5MmXBc2+cm+35kXHikK
BcOk/fsk1V+caL5pk3ZowGgKDRyrqJh/irOFdSx+nAX0k1l+igxho6E0iGdJ0+UG
0kKruQSSRZwafjrAMt069n34seEWpbEFjDvkAMPghs4xlqC1qOiZlFKgbrT/Lxmh
LU2q6Prko4VSegiA2yQ8aF0/GQ2rbF+wlAUx7DX55ZtvcI1dvriwiVgBKLvYLh4P
4/CbFOVMQ5R+u8UUxsf7x7B7yO4b3Lsn7JGSX7ws5EXnfsyDQiTRmMIvWVmZM+VG
7bTRCO471XCJtvgeClipbKJE0ZSjnPvQ+ZwRdLh9NnsaU6WXqg9ZS9MGDqzJ67H1
5STq2AlFL2tt1/m2Fz8hQwCTyjaNCW9Fvhk49Jmj6LV3kuKjC+1mvlarn+rnl7Sv
XJ3V63VBnZo/PovWBfjoHAzfqgb5qXrAY+9rW1nQQP5zcQf8cIPqYR8RYM+BS9yU
NzXCZXNP6qD5kiJzcZuGwiWkr+OXTC8Uoqg0Fq1RlmJ2DLBYnj5XOxuff4pbHnxF
GCZ7QNakXv1NMLoiq7l+Zz7JJ2z/7NXKbz0aqHzq9PEHdr3ZJ615FL9kYhW8pMos
BaDSyES3WO/7Ln3wVEAZKcGI522G604pTCkaI6m+rUmheaslXi//HD43ttNJWm6y
iE9bIVzPmSUeNFSg/JISN+zvumiuP5H93KvO1x+ZPIGDxp84XxttXcGIY0XSyhyt
5s5hUwFjTSalh1prhnpl2zyPqKX0Hut1HNUJMmHXunfxQrTOLI460lpSCeWnHUQe
cRmbt1MZIpR6/xzgT2w0DfyctGO9Qcz5R5QQMRNtaJ96xq8R91Rn9szQ7euiPtZT
fYNIdlmmfArVWBoV3tIOf1OV/p0WLqpx8lSRMM1Y5jjjDN6ZGJrKrw0WYy6QN+Y0
+TY868Ky/HWsfVIq0j5NwA7E9Sy7doioTfSE2azDn+SfnLz+KI1koujHD5qmNUEw
2Mhnxls8uSqQ+uDTtzV0IgabhZSVg2W9+7hZme6AzWl2gOz5YRHuBwJViWVjXBxM
DP76bdk3a/3Z4IQKm+4Vn9qGjJEJLYGuIF1SM09zDYSAlcwEialNdO15SFIBgg3R
VBfww95ArjFI9yn4UyvVlcKG0/ld7WJz31Pq89KXGesvE1AGw58lodElJfXWM8Yy
c+JuqjPaFLzcGq8C1MJQkXCrRqh1XtphZNQwjBa5BKn0kzBsrGd8iP6jt5AkoQP5
nccGXugvhjo2/YzsmsPIvEMJmxRYPLiyzCvsFi2rrGgOW9eLjAvYkyx2SWEh+mi3
JoqQIU/woqz+HFCIsZcfIUbzqn2oq0prL1n4cZFAiMDcHRlN5RZyyyfwt5OeAlXh
f5IYt8bwTKpstqdMW8OSz/ckylXBa4dUIFDzEXLh7GrYFfaowOcy4VDfuv3s60Vs
hRs9zYgyVLo0ZZ2kHu1WhCJkbVC2/LPLCDeitp2rQvebMB6cUTeqp0vdmywuxYJG
6X0kQ8nmWjMsSabceO7JIwUZN2wJ8gZBJpeNultihVX6Pouc26/e9XibG76Q+sdi
rjCFsm01mYamn+wn2nd6rzcNMfu8rIleNnMPqbH8lscUrtpMENkvVcnRWl66Hr6o
pyzPiZOX+dFBteJcuaz1M+ffI4y2E/gsknh8ZMK4KDItRd4a8npTlB91WHX+JXXj
jAZUvNGExKFlojvU68tZlkCXaUsMgyTIqMnUTlBZaDLMnTnOwTR6HfmeP3TRk+1R
86z4rLwBnYrOKASQKDXAMYXWzh0bwz5NNQ8XCRZ/4a+JvLl79eWiE2pbBGM9KXH/
il9O2Cu0RiumwOLHEzSqQ6yZB6S2CU1R1JImyW0mC/8tgz9Jxfc0+8OOF5luELs5
HnkN4EMHUtPUnadv9BLDl+j96OKCELt8e2LCorLlkw74adoptcGs4PYgyK0ysdzs
mXDKoY0GSImkAsD/BKNLZrcCOjvKK1d3mqgvHDsKdiVAuZIZRgpCiH6wC9ZkYcth
3+j1OW5O7CRcLXnOlNvHZrSZmuW9GUzcruTIeOpBTr/2d0h4LmecGsJWOGj/SgLV
v9SDajqhWbJ42swM4btL3uEQba7gl5sFgWlAKL9M+ickJgHsRsZqu6yVlBCMHBrK
BvHZTVbF2zG5N2RX8zTJJTFYn5tCyOTVYNnrwe5Hyreco7b79iF7V4Bn9ANDZL7S
wZgfUHvGRDgopjO2ddn1xoLoC3xeeV5KUTfrfGoTd6xfwfZ14jXLfGtInWW/E3ea
CttyaaOMPe1OcRdrQfgky18ydsiuAM77chRmy6BH/NDKyEBlO+oW5zxwiFzYwa31
oHmT3hbNqLfAgnCox8ZsLD+0d4hCdNb1w5brYCS4ryLA5uz7gxjdaBz9+RNwELL5
zcfT2eIDSZV2PITsKtOP1YrWRPAwCSt5tbX6zNbor60b13wo6XPtZO3nWa+kuqfA
i8QJPgWYZnUaeDW0GmnF9oXlAQv6gQ7jR6Q2IvDJYDxgCylQXTOKX2D3g4SUcBay
zD5QFDF4Ow8l6wcdomUkFA3GUEEbiUhBISzawRM3UrushgRxwBL+Lez/GwsRPwMQ
Z2cte3+HgWgioX/YnQlssqfWF3zZI43uUwGLYnyOgn9OP1BU3mI/wf0UmCB01N00
VnzxQPbSycSGujOYR5TrbJnc9SOJnJe67GxAq9kf32CKlz5Da9l4ndnlNBz4M3mv
x/+kfmya9OE8gQSgAQpGlIBXLrq/e+iD3UVEqruKDp9zccvmtmKL7m25K+KMVCLh
dA4W3qTiK0WuZoSuI2qbcXyFK0g5eXDuEksLs6LnjVg3naBI0zC0VoJXzS3ZD9LY
jxZXNDWWmW5mJl4DLuca2kTQGpE31cXvlaqWunsC2lf/dm2bX8T4ZO0kpZN7IE6+
9TrL5MvHLDu1E9M+cChez7vT9CCfEXl+LLVkOgGQVqdu8i1DeoDsYxoUpsUF3hJ/
f+8fz4TQfJwZuDErEIL6aiuTyU7VSlO1S1qQp1HQLWPwNGHOSRTbAd4AlPpwTx/N
cg6LOO3T0FDHJoJkZap51eJOK+hFow27MhXZHF0YWxl6zbhz53URHMs3oLI6eg6A
5aK9hNwVkzOsDTOYLgaio3LBnT6juWP1+L0FHc13yKizUefl4XLT0Mjd2zoG2bVY
5K6OA0N3lhQEZHO+nNr9OLWw4wM+bIe8SxatPZ/YLCDFpo8yhIQ6a1UqQEb2REDV
eOYGKXSFpJ449Krnky/5pKgvAA3SqRAF3tYTu+VmWkNI9kfiQ0Qh/m0U4/4RUV3W
8l7DWfNpUQokAjuW9RiFszuLOPkOn5LOVkYJme6GcGoxNtQYSr413+JO3MPZZHMt
f/o1O3czRi2JRgk38rZKljMNMtT0MuuC9lGS2T+xjRbQ9sTcYPwkDVYoqJYIxq5/
fHROcb4oDU2kBBWB83+Uwcfd7q2af9E6/TtbyCcbUDWn70oJBzQJ7/2RilFRVsMR
Grrg6isN1FZDLcdyef6h9rdOw73i1YpKo9gGahr49BOsMeYCtWM27W/XfPDWnawF
iJ/CsOtP28g8sWjvWN73hUui6bxb5QcigjjNF1BS3trLiG84wVEAjGsgxbOwJfdM
4JzXlxXYiyGKTkfMnjhqmDm58Stb/McYkBU+ZQFvwIr/VA40NJsaZkwj/pWSW471
aVWgVHK9g96mlfoPPxpEL9CF+L9U1hWfYIpRrokyqEi8QFkY3cVfe2IgFcrK5zfW
IgXz4az/jmKvJd/Z9H2f6sKNT5M/nNrq/X24tHfK9Aq/ybTW+qEjSDSqNMc5/d3+
c87j3/i+XBgoA5o91PthFABG/wRQTaXTAI/BRWwLp9ajDitokGaJQZS8z7biRGjj
oiL7HJYTzbm1ceMKg6xn+20B1WDtZgbUllRXqNcV53LCy9BZuttOAGgBgGk5zmPM
t1uL3IFNLlFohXalsqmyzgL2CTZfPc9opQTzLYdpxG1zTLwmDZ2IIuouDZ/15vEU
WlVj2iTw5Y1aq2Pw4+l/o5Wls9rHbufRDl55lTGG/6S7joZeHxQIpTtbszEbuIYL
zVZBRiWT89kJBrOsxZ4ijDS9cPMzprYYxdoAeH9s2mPM2R/WNjzLAhOVfkThIpy2
rg6ULwkj6el3mS1HvknNK7JAP/wC6wqrK5N4O6GSGlUUz1ty8CKcVesiHuuH4ts/
6eovi28S4CDEQRvOsoUiShS7rusJNTFknjSuoIa/xxG4k1RyP0+oCua7PqeLY/qm
CpwUSog+pYxaDIXCx1TkF2kF/i4pEUMrRI6PCEjkiGV9KjEiz6s3eibe63yobIe/
onKQzAQWKWdf3hf6yuXlV253w946MS818rN+wMwfAWk3tLlLd1svD7CsG3nGSFjK
8f8spAx0p+7aQFyLnb71sGkpYXfgfZfxANObenCRneRieiAv4A74JL3B/5qAYThl
BhSdlX3Ul2ZujlE20wcNNgcTIaEROK4hWo5e50kYP8T3bzUAysZo4ejHKu36VLJA
OOMOgvswFhHeBIc2231EeMV7FmpQUb+AKSIII/1JXrIbDuKtrR9kZyEvgK5cQ28V
/kEzdbbOukDRDHVZIWNHzEVvngetMeM6v9t60XU6ezAVXTdNuLx00j2zR0qJ/5cU
OcVsp6OtBqAC3PyfffcSi3gzsieiwh09Mm0NH293TH7jxE0ca4S4YDwsgxJlt2b9
5++RC7kLBmtwSDRicK0Zaa7TervgD+ifiGnxOA7nzo6/OSu7/pQBE4LiLz1kbv6P
cTeXQ8EVvZzzewmcDitmeCpA1sgsQCNFHFLQL+64OaGC8yZipDdoA8tjcLvPqPGv
roNso/dA9L6t2nqUEG3bvXlyz/Nr14iE8fPXnBvqvnuicYGHP0X4kveHB6ETyHT8
imR8vGIVAMFdOiznm2owlZbollrKwCK5pTokyqrLI5j2CmqAPk1QLlIYp8XRRsED
8w8VKwFVMPicZxXPwnonyE7XSJ7XpImeCzc2WsYdzvQ29ZakeANH0DhkZo1T4WLT
KiI4icP0tCQLpvGnzZ28iY6yTz29z1vv+TcIWEeMWCnewbYWNiYf6jCSCa5N/uzO
qS2SoLr1lNRNBbmIyxre+/CFess0aYBOqJZB0246k5ZTUz2L5pv669yfpyAaU3t7
ozIKtajlgTVkTwvQlMdu/wTLxD85Bev15sHmhVrWjRu8HjLIhtip3AjDmxj0dEc/
Sdb56w/EoixfJLBUODjbrEowXhU0Ac/dMchKNw/waeqwOz58iNjiwZO7K+K0dojm
mXhKQ27TnzOE6FJhIWnjNf5+dC4bMEyCvehnml3B8zsskZMMnf1sKhcQZmZu0NIL
kvfKknZlRvwkSCRnep/xzLWIqihSj4DQ7d1uVyezZT3km5Yw69LHyfXO/+bunXVy
yOBrsyqU0INXQnSk9V6cxiHGOoFA0EU6OW3/AYnkczF80QNG1syjwOSqUdunpTDU
rAFeeZxp0FxTOgrU7n3zOIWr9q1QDxwNAv4hPpfFkbXIA037IIiN/lvudU8U5t2i
mMfd9WJWT5N/Ptz3X4xqWKraa8Em1cV5Ms0vvHXMTxww2TxdfOObSEOKFHp1QZ0y
qjOuqPLdQ7XsF5rouUvz1/O/UrN2aySoSqzWbaL78/d6Rtp3W0fXBWHU4rCXh1kL
UVlCyz7ReTOigezhUoZUZtYf8TkrRmg3whjWVDrihm3q14+yuU2hCk3oHbkxuY01
b+VkjFDMJg/wJZKpuN7vMS4FRtjQ6wB/7gnADDjjE3a0VCIk5SsxxTqi3WcNPlpG
V4rwa5bypa2846hQ5ofcOZ1eH1jSi2t1Mh+XMn0a1n0n7nRD4Y8ejBrABSNsewmL
krRgyiIbWHGDAYG4IBC8xuaxBL+9redH0FBJq7eDnAB51DESatOo5wBurexpnjk/
IxnrWYc2UFwskYaunf7vqW0xug9Jd+56SgpAqLTPwo3LexabTjtFYUrUb9w7bq5V
SE6bbC6XCeA6skU67eJhBZKKv2MA7vnX4ijv35iXezBaxH6jwa4jgSG07dwMeSJV
+fc4IoVkFH1V1/IiMoASQx7Eq4N9gNpPX+7E5x7IWcBEQbo6Vk6oi2emsOlbbg5d
MJUssrqrS0/tlwOlFfk4Hn6ZxW/Vlb3XTHtHfywIy9oZmZKs0CMn6Ii4Turs7z5Y
ihMfVKVOrb2lw/1KJGjzpfP/buiWwt/HX73W/6m/4BuNi4BTnc8jZX6W4i4/UZLZ
1bEWIwwqG9rxAiRqfnq8Z3J0DLa/buN+j/4mTpomvNEQLgiI2aJaD8qLt3JtKxrj
XhU34/ZwJMvR6WWr1ABQtn/BVrqs0d3mjix+1dJB4MjPQ9AQNyH4DybxFwwlR/Yz
FVqBYacAvkydfm2IEJ7i82B2WIebLpj1ROKqOe+zuYtbXNRYSUWTfpaL2koyUmpA
qzPbg3jRJTEjslI/C3+bIoc+htzZAUsXTkENBRfmrjDf/FVlHVFoLDz/tFMnN9D9
121ubGbpQozTotTquzGx2gXzpxGCG5IZrkuSxDU1gh88a7te3vnuV0DhatIaRd7+
cnuhf6k7Caiv/vzk2dVOPrlT5TA7PRO09XjRwkxVHt67srVxSfLXy7G/npg/P8Dv
x0XsnGCG0QM1eD10EO3/FXP9dQ8Oz0HVUDn+D8fnkwNuw9duPx9NH1gzrW0fcRKt
VHunFLs0CM85A3d5xtxQ9+0RcIN9Va+AuSDsWdc8z/QUanPkfO5KNoJ50v8A7NQl
zT94RFzPWaO9H6PHcLVoX0+qeGxh1eN96wq+By9MBOy/8So1s8GAjLpjMDXgK5Y1
HiJOJAAz1FgfVRuekdTkqHax/6vKYkp+yUSFleWlhatgtlseVzKckaX8zETQKIz2
Ntnl4JQkch2vLRyK0iTtjNg+5IDCoyeVCVdLT2l/ZAON2KYBsDl3CHb/F02h0cNa
eGmPD0axGK7Cwo82TjbgJai5JuEj5fkmZhCp9rbasXQxBk9+nu7ZRAY/QHWIkK3s
oh1vvzhUMMUFhBep5TvP+b1OPCIvKzXHr+GFvphjbaoxn/Dux5cddXEqFaQxVH0B
oS9CGlnOA1QafCZQJhrPREZDfRQZCmok/xuTEngh52rN7cQZ3T2dtBe6wnK+qGUT
JZwTIdoQ6hKTgyeq24/AAar/nflCrv5RqwdwN+NhCZ1Bien8Gtikv3RcXS82U6gS
XwkxefQJGFV3SlqNPBmOLuZY8+z0TuQ6YkoWcjity8+SkdfjKJFPESYi39dI/5D/
ZG+HGbmJn9cMajxtsvZNv/SHVndWDes5LUEHYpL0C9w19OcW7RbBwVGq3/9DWxZo
EJe4bOz+Ck3xDiU1nFOSqi0knzMR9AqRWOaLcLE1yLP7meAc4DlEKrGw72fucvDF
ka0aZMZQtjsOPmkQ2bF20S3dXqPztKsuQH+5PViSpXOT3jTtBmcHwIqSYeXkNRi6
HASG9GBARIEfmQr2Eh+rssB+mzQB/kwaVhfBR4E3f8upb8RiCAZYawVya6s2eETs
8QTM66V/19sGK36tUkbID36N21Sfs9zHL+WWSSwPMXhsdrwgXfviMg1OSLE+zuvS
/fOWejb2lSpjBYcsjSYZHTpM3mT+kD4voo+K0sD+hnNHX+NPFVLrH96E6YESt8ye
nl+FMwJS6tUM58AUpoF7XZNEC55bNo1+8tcqd5cZjrMPxt0NvKQyAQOe6qv9PvSu
05DVJhioaJeeFnwmp1Iu6yoMwFJvSogjea6jTOOT77azzND1NT5Ru5Wuf+UF9QgV
6hqi5Nvv7T1QU42Lq6pvMkNGkU0LNAjNWuz+TiNrLdCNAhz2QoWXT+XTjsk5t9j5
syAvIyw3akf5LR2n48BfbMQvai0Ky59PqZRO+nQMEC9Qxh/fmwpd1Iyf4kz/HVjx
wk0qE/SAbcvywA0AjvUpmzJhCkYpsPXL447QlYbfiMYXOePjCI/cLxBk5O+ha6SE
r5pp27Uxh0MdYauyPmpj8fFaT1ecD15tWDOQHu2fmN/yFErpnbozCXh/Q6gi7Kff
y7XKOxGWRb+VROE+pkCPrpbO7dR2mmY/KIjg5SuylCuKRAwmtUs5oXK2m7EKrgTl
ASa7qySNaQtatrv4fhdxkwCtmqKN/9h8sIuWO8nDMJG0+mQBAoJ0gvWhp14rL2si
xjgmv+jyuKtagVaR9dV7sqCtPdUNpgNgiHJl9qlgW6cSkuk1xxsVxtO2CYamPu+v
yiEvT5xyl1+xq0w0a/Y1QQXt5U/sVx/petM4airyLtOlXd8XfE5Un5iHOAl2gPm/
rYTMSRk/oxGmXkuLeHOUy+FJ+pmzZv5S6BlROfrV/tzN9b9cACLJcmH+/qVq1dUD
/mX+CcXWX0p0E8q+7sotaw/Jr/Li/z7DCVPmKOLwvZv5eqttvCUsJdXeNGL5nILC
LjcRbYA6KctXpcQNtR8mgIVwwTj6JYwZZvkJBE7H7SRxDFWuMUmKbDk/chhRbOfH
WEj9z4ghuQ+OwI6HU19II1IEHQQIyYCLZHfLsMXipIRP30jTJpheUjMfACaXPkaA
cRoA3dtCRbpwvpaWp4dF2RnI+fxmdDoUzvmdfRKug/5PGTIETlg3V2Mja0JvdxJW
EWqJwquhNOJwEjoKbaJM1jxLh5NnRKb18uOw/gF1f39fufyb0h8FSpAcif9s2Bkb
EkMXv8Hw5x+VP61G0RFXX6NtOE6d00+B5QYaYF7DDWHRYvG/L0BMlxuwGAvj0KuL
184+nTSbkw5Inw/iDaQa7HqxRqDpa5ESPPGwg5DldpxoxJ8B2BSkD6adIMEmhKuX
LPXgHK77G4aiNto/j/yb9w7WG46vFlFw49Bjb4zGVZRvpN/mM2Ygzj75Xz7EN4cq
p+pa9vRSqvTdmDPurgKYEQsaipvqJc90R27GLJhGOqzd3p47C2n4HOWykrDQ6Yhp
jqayAGvToT5TqluM4WjJt5wcQdcnaCgSMwEalMjsC8zd7IPHRe3zyynOAW8XyuAD
K2jbFoU7xmVK/0BXZBfs3vFGq3i3S/TWdLp/MbBxJ70A3anGlXMvps528XCnUoYr
QRAZuFaeif5ILwTR6nySNCAD4EoPIHksASqo1xyIsAilDdMTBO8aPXXZAutwNKDn
kuTJJ1gkEO8kR509vUuBFhKoijHIDMVCHPRgxHcsJ3XWF0rz/rqc5UNHJqp2fSUY
10sXFh6Y7yYQZRnEjts7HI6+uzbLUmi8IMAboFLmqBNnpmGXObTBu5ygIj1R0JLY
wVOL3xKTAuWC21J9lktvrPzH0XdYRd44hzVuuQT1bTN2AJJvWC2J4qerAgCZWkL+
2tnbT2XJcTdt0pd6bHLzbEHN3S0Srfk8IvUGdev6QEtroq0QFhw5E/eSgV3ngr8U
GnYK9TyVllW4c+BZjxamCd9yPwPnmfedwSbdAGJ82d5PeRg0uaqEw7AAXgrT/FFF
9alQeOMLWDdMxQpxDGGkfhKIXvmlzlKpXkpf1FGj15qQIw339SPz10FqcrXMZhnZ
oI/9DUcTIe4o6kMpynEg1mbycawGkBvwNt7qC2kRqOCEGVU/aV8FyrHRfeiFbcmz
oJHT3eiX/Pwqv6R1VovgkSOYmo5PgezEMW54ogJ9PDf8SX/1jApDNH2Cq1l4Vjdn
MBvhlLkrc3b8vJJZ/el21C/1atPiVoyNGesAQBybgFitUqwRAq4vYHQio2H8BjMo
awyU1ZZchk6HKKwM0dtXSZGJbDD1psEPyX9OXMR0tp2kKq2491xUAFPsYJC0qUs0
hbUEfSSRO37ezCjg50FZWLE/5tGaq76M1OyGIK/IK7C4fwWWzDcUO9dph1VPL/Tx
mPpPhKh2sebzTU5r9gm0O4kHcdcSne84iCGPpDPxiisMZjNxrknazdJX7ucjtR/R
1kZPLz3sOjYpePdMKv5FdYD5vgSE1fLgymQzAYNf4RjusKm6zDXGtFQdgSGoguGk
fz0sP5TgW8GG5Lq82QtMIEFn+5sbrXB/RkTTzKt4n32lELVqy0+oE99Gvh4bC9o7
mn05vfY8dqRNzF9CYgFr1oI1donOPFNn2T7T3LqqIAeMD4qiyLU+yrBOCsw8Fq1X
2kczMUg9so321TKmE9wRh7xotGXN+X3l/yOAWHdaKXgTpAw11WIuBeEi5IvNmwLt
DXt9yN75Q5j4J3ZZ88xglcEW97qZyyDomohQHOenpWOAygdmT5pCd3MxV2j10UsJ
M9VKnKu9ObPbMjNPdQEcNcQhqd7Yyh+C34a4mu452RqLcKvPVp6a38zHbnra8t2o
4C3IddOYW4b2NZ92AVR7OYfofp2TnYBVa1sRzfmKsRERYsLQ2+7THzRQrcyJhuFL
pYFK4pPir86uWDlQH+nl1RtshsrEqkale4Zc+7MAo+RNTRMX0UhUonYbjRmi1Tds
uu7HB9Y9Kv6NbaNtRpUc5ph3BK9hmIddBt4UngISSlOUgc7q/9LGZmVYfvB2NW8o
4pDWfFYtqwguZyx7sNz3ytid6WkDylIDL4hf5WG4mgBY/rJq3AyIocwV1Ya2lNNp
viYg1B4XUpcwsk6JjD2JQivKmoHcMrmRLSGHEMvC3iRYQGj7/ZHuotNUfAJDa3sS
iCAYRvaxBvL5n/hpujPK9xSbn5mynRKkJYJ6R/3z54MNNf1eD/ojGuz6IvqhyV2s
f3H2oQG57kYrbnVTSxhVnovWcHX4lQ+r9OyqyZoUqyB40u0P7JD5cNVwFmXJ9f81
FVWmljD2oSo60jfj4z5gkrLaAv7X+s9Po3SAhnznXTAGjynHjw2JMqbr/LFVVNmk
Bcd7e4RyBtd2+Q7OEtKv+Z4NmN+3e/qhz6/Khp45OkB+nYz5QzqvWP59+iNe0k1b
ugPcUL0GEUjFzr8bJuS9t1i2D/9PBzqkOyFUD/4QiLn4QcZXyyjQPxEh8V2/k90V
LCWLYrXPaddg94YjwW3pnsakgBMg5n/3exMkLgr9FSnAMBMKyaltV8XPuCDIiAk7
YqMdbXVuPGf/KKgtO3XVa+JtJ3MF9PMKJU4WSaPhBQIcUZ4vlNSiM669UEYrOWbi
M5vPyCS9oypznZDbroi3Dr4695WBz4fsVSt/ud23ZCiKLjizXM0SZzAp8Zym/Ud+
vvaWA/ZRwpL7G2GAvFgLn1/t1rPOviMBw0OksXp9pmp+QvRXheLTXV+lZjxgeifc
/2RmfL9VNYgwjciDpl2dJ45jeAQOE0j+uOZqIEXWLh2jMKxtXqtmw3KYgjJ2egBq
5usuk7iSm8fwU3rDPMQewhKKPtWwsQwnuOEwP+kzaJIyGX74oVQ0nYyZELMiYOA7
2Ah9iYBGn2GlAGJ1vH/z1aod94bbymyARaxagrPXKF8metQEobw7ZZPeSLWAWa0t
Z1HJLZLdzz8Fl7GX79xnMi1KAErBwjR5dNkM8hAvjjp4+b8s9LZYgJBM5esI365M
lJhdJJCkNf+sP68mH+Tyi9bkPGsKOCL8naC0X60wEpc9uGrhiV7vHeh+EpreP9E/
IPHWQl02UgWZvwMgOHy5przGHWARYwzNcIg/4pPOv3RAwjl5fksbQsBetK8gaSYu
NeM+akb5RqyGK3gM3204dGy1goFjiip3u4PPG+LCuLB0Vow3d4KwI0EkeuzJSIj2
TYzMpz1eG7PihHQZQbA5Pkp5vkZXE5azRVKYa8CdEjytk3oiRhwDfdT7++0xVU5e
ROtu5lTWpSKeIT+cBcUSmvJo9niNIfP9lOa6ovNt1ABVgTyvkaSWi0NpBme/5Yuo
GD0JioB+dMdIGLU1lRuGYhksn8pliuCcN3pLQcsfjvbKdsJzEMe9P04joIJ4SlE6
Ea1jrSx7Zn+okhbPgv5771u32xol1oin0Fm9uK2X5tEEdaZzE4rp8ECv2q+U9nls
IMbulY58TnIZFQM1QoG8wZSM7/vexT/AgdvAZ6pOlmZszza0ANh7IIU0S9Uyw/Y+
zy7Wa7ihM+kSHOgJbiIHxu5wRZH4JH9IR4FiUGxZjbxf/EMzcPFU7NDj8orWN4sp
eYPQMRa6B3lrRkutO2CQtefDNCy7KWlcSL3F0YSpkAQP8/dHn+XtvzJHtt+IXRJY
//bXvbJ9UXJabGovcO/suySzzF3PNivpFCIrLW4ZGPZMuIpPBtA56tUkhiWoz0T+
stsVO5hAqSQLm89V4RY5V0TEcf49O1TKYuy01/dHHXuTCl3iS9MGMQa4/ynB7ygE
CpreA3JKDB/TULr8fEB6iqCoSO8EzGR1IyAu6E4N4YyQsJiHZnW08eCPXZ5/UWtP
nwZKYAMlD0y6L2KsPn38RMSNjAtlqlPuBUuloLC85sX2gwQbZyjDE3GVd7NlCkZB
hXgYWuWARBO/45qqkSF+5azsAXl2cc+YATOrnM5AGsnemQO9VKzecv7OHrCkuLYt
XxLJJrihcr0EWlQczN+7srvONpTp18OmBrN2+qKgiUVd7wHjSz7UWUag2/2p3zMy
PnaGnWw27SuIltEEIRwG/11vDiGyqWv4GMBFKmbRbBGlY5Q7W8fs75qxRu20i8sX
LtsL75OMfCG0p+/JYy2IbrUETmmveKgiCDdrEpiS9uNhJW1dAs4FSlyftK+xpMNk
DTqOLo+nmOC9owUUeDfAmN2MIn7YbZT3XGrHivet5sbzIT1VyaFBCu12bO5RuX54
rw9K331itUgfntPKv7ULeON6AUtGJV3STRCry9wOwtnqcznaY0I6lzl4Q6PsO2em
doR+fdgu5qxlFxb0lzITXiCMwrJDGqRwAUWRRGBt/gx7Mu6jdgJyvIQ7Cjj7m1iv
GosEeaePUmGP138C8HVWPc+EYQVeSjP0yL6+r5ucF9YRgE2S79O2A/EFjzD/+1qY
7OtI+nF6h4Nmvb8/92h72C5d5KZR0Op8UYjE+0E735/onHXuuZCW/Kks9jHJDexs
+9Y14QdjDnt0070Gbl63i5pLI+QKUlAFSWLWw3kyH6KFrMqV0I2h9DMLgEOlM70V
5CDzu9jfqJ6circbkTwDmOXJS/PHYMR2S+zXxCgCLW7tfZYt2Ua5ZUa3IxWOvf5P
t4Hwhyu2bGogBEmXmlc/Dzo42I491LZW7dkhRl9Wz5w2AilPbHGAesoaCy/Jz8xj
BqxhyLEwiQhbU6Vyv0yldLsclu9POhPEtvSMEdTmZovmMu6fvvq7uCV7L0h1Pptd
GshvM8KBQg+z4wtelSjFsqgyiOjwerQMoa20cUlbF1qt1hXwpXo33E/CygcS8pBu
Q8x7jJZ+j2PFQe9YeSNQ1WX2lZfKt56g3+IIoPh4CjSubCVI3AAC637OiELumyTv
TJsI7adSlII0yxj0jWF80nRIDElBFYQfwHxhp41sXnXWhntnTCnMbLP21XVWqahi
BDSc+APb1bq3kO09BSFDXs/IYU5V713uxEGirFrKLZd5KTge7iCjIxe8UNgTq78n
0aTx34A3lzm+RFBACXfOiqfKmBVWOQ9iGUWM3WTkZIE4F5n1yBG5xI0+nzNHcgiw
YCpfLCOyRbkUiyKJqf6+kzHv7NGy+GhUpis5HwaGZuOa9pua9RKWUrugObWywV9h
oB5o6M37XFYiIgeSgsnZgytKRlmdQ5C6iqH9uZicxbGFStxYrPHOGrCq/yBb4aMI
nCM+09IlRZX+16gLZK6ud0gPO2gF24V9unyzjBHel1jJcWTDzIl1EZndETIDhCUo
sfbxocVKfZ3j7Is97O9/K53GpRN9/m44UtanqPuhJRUdx4D8Dl6oSEIK+sy0/aEf
Lb01nBI+vD707+Ssnfd3qTsKtgmCbNGueQ0nfJHFsIpdL//0GRCzxG9N53Oly2LX
o2iIaMEcHGBk5VePcByFOKb+sVIQJMTOnQ3JL10ezW11oDb44BUfyZtSxchGhsK0
w3CyK3txIQICx0jGh4SobqO7gxvgJwCMTkgCWsXTbqtYE8Nw8bZFkvCBPpzI8ixX
NF7q0WfG3pcYOBJvTYJwCs1Yu34Sk5hBAKFbrUIRqRtWROTw/IQ9sWAAjSPF5sfC
h/jwLsKN3PVUSQp5ZQ8QCGL24owq7NUfjG3m9jSd5ABqCcQMe31GGsOc5melnjTp
+HXMnTm4cRb2lX0WZO3dBWqt7UJ3OUf4zs2wppC03TjWemc6lJL3Sz2ut5Qjw9zZ
pJ0LULDeNgilR+s4UqrmwW0BYIfLY/WcUKajVt1bDR+yrkru0qa0qPs80vJLBjcW
r7uy0/7WVz8Hd2cgPCuAnzp7XeAodG5nSOcr8SSmXujsFtPSthlfMdfeP+O3Erux
n00Q3NZLo1ATvc94p4khVKQT3EY7T/k5MStBPMc3ok0XCry0B2uzsLlsJMlJD/r4
QmwLds5bF0MKKDmXVgGIkmF8wND9b1w2cPNqOTJZVfDgQG5tyPPK605EJQbqrin/
7Q5IRZjCIl/T/LXyv3P0tLeVVPadh3Twra8OdPhL0xC/K7l3yCYpiUXyjIbItqMG
yhWBSiGHNS+m3Fh5MNIQsNl9xOcTRuUOXw0vZkUXtQD7wNTn91PAhJ0phPymItWK
75Gb5XPZN/WjTUhHuVMKgSORX6+79xwfLCFqtxy1YvjmB5ORerhEwfRSuP1NLRoI
svLvHy9mI/rDrhKhYpcqujeiGH8zI94dulG7p6NZmuKGiGJOUNXRXjhLoBJ78Pbi
jgaMULI0B0jRzb01Q9GAMWy+Gp0GrTeHYTlCIojWXNaQwwTrtKxDxSKmW72g+oUg
+gn+/xDWiGTADH7lxCJeShIf8d+yAKESvpEc3WJ03r7qLTz5go/9CE73O9jQnKL/
TqZZYk/V4jWycz75gNpJbNaDaBQKlBdT3acIQRHotF9QphugMXlkt6Y/oCxS0KKz
yDIdHOQkKfPFOP/J5zK8TFSodwEyEuG1lYDd7fj/qwtPpRYibwc7SuYUh16p88fq
8MIHNV5JV//Zl5wnK8ced16xJWnbsHseXv1iDPQWBYHjWgGNGfJHUkvAIXNdche1
A9fVpNlKP3v+BrxF/virxgLSUNT7FSr0nuOD3Ni+CBDlkXNJ59QZWt94G1tECyg7
PPN/X6LwLND0ITTgvvPrYQwDhPp3Py7KVkePPo2pOhkwvCXnwfuSiqOwk5UHEU4F
fh7XYiUftFxgCemHzouMtwswjP2VZ6yI0CCdRxpuJ+bVLSOSvqPlnBC0Nj/O9bGd
jALzE0vrnGaFV28YORGg9YBWWbQe/GX/K7uuedBj/sGGrgL2lmknKnDkPYjs7E/T
vWRVlJMH0XvJBLZSRto8P9eSMGmLSEcoAQd2RfvFaSOe0Jx/gu9b1c8DeV0y+PqG
Ty4BZovGk8TXsVcqptHulS18aoqHUj2ay3Rsv0Z6aI9z3GxyKKB9cbecyXHQkPk1
hZ/bY7oCvXOnqhm0aLj3R7pZE88w8LQo98TnEUgsarrSp1hN3gUb6oFVYPMeIcg+
NR4xdBC6vcXxr1B8nD06f9kamLJLLE8L2m6S5NWm7YgX/leeLmgOeInY0TFkyhA0
Z/zCh/7hU88Z1EYAX8tJFKctW/1CfeYbJfT4ce5uVl+4chNWOao9VyCUr7mFo4RU
EzAsL1WA5Z7u+32x2a5E+eES6P/4C4WJMwuiWzkf1vzuruZBv/tsBzrBBq6Q6Yjm
LmpDDM3Y6vwEz91CIsF5v8WToriDD/VUCQyuZRCNwaIk7pIrnBIcCS2afAZNiZct
UkN/xly1SqxE0U/rjDSIgXk36VHEJAbCuzX9LqdcgbnI5Dp8AFpoCeLKAeyZx4+i
z4NH3caMDvjipDffGr1oNWe5HQI14gu3QRcyD89mnUMjC72IgkqLG2Ujp08W8S3Q
bdFN3BreAun0bQxSEJc7WnyQK/2nuXM3FEpGyUIvmCAt5NL9tx80F5af1SYsFm87
MegycOlAKw1/KGHt3SttFtr8cOFTmH9AX4HCaWWhf48oDGl82hR6eoZc8Wg9S874
GkkryH31hIKM7lsmiJs3skIUVmf4o1PxYcL2v5kEB5W092R2P2cFBxzZdRIbLJFj
gDYy6uwX2XgJMNdwWJWUHbzauDtqnlXrWBI+BRBMdbqSl2UYupXXoXA+Sjx3X7QV
n7FjZvgf2wET9Cg7uyR/mJjLhCM/5xzqAoAdzqy/IJGK8YBjDfqupPZjeJ/EhqgW
GM6hQ6itfFFj8wxhOwUW8V+0LqbRecCQdA29ubBcMbEUmcBW6Fh6AOGNiuOw04Ji
KIBh77lB/qLh6Ms2FtFaHPB8JA8pc2TmdD/Ynn4qNa3AETkvKOKYTLpofJZAYbRO
cX7oGvr7gM8WsatCIXq1McFLx8EFdhE5otmZd0obGTotMG47JqimAv8q0sUK9O+M
g2Rv8zKFNkh3lJqr880UwBZJ6DUTasCXfGG5lBzgTU9FTpM7gWCSXRZYU060VkHT
RSCddc+9xgzN+xwJu5lSsZXUFfffftYUtwDQZ+qBCpkHH6as5rLOTM9UFmmA0txS
LugP6o1xrVuGutel1Ru6eK6DfKChs+s1/8GldNegDdwGxbkkBqrds2/kJX4nYaqM
4UfDUqXbMtskWvVmvCWJVA4CwRe0/2nyCVFbt/FPaH+RjYdZczMJoXLrE25dCDpk
xRuesXyXMaUhd/w/3S5+DW0iG4fq8URvUItCmH2dKMPE18kHY/4mTq8nkyiH+gP1
T/IUgRNbK4h+LmcJYeL9zDRWmzNLjJh6ZAxLmLL+kuW1zEaepBcJB2bJZx5MTNig
w12H1oZvGT1e5PbdXA8ZnlV3oy7tjXG05nnE7R4Ef3E45iJiN2tqFqP66GFv3X8E
YGnge09snDNUqoWnwM4ZBxNB58YDTRd40W3niJNaugS7bzTsdp1xNh/uFSkDTM8d
Ie4lBD6+cu/b/TvcukYbgjXsWvFkJ2rgBvNwQid5KbW5Lk8hLxXpEkSEvl4UJt5o
dSiRBOEdWlzXgzO2RvYPMwNBnUh+xCp0qC0FBembSZJ0bP9Tl0GOPJf4y1R1dB/Z
DdVTfRFmXEXXR6mbCxD298BhlcxUU9iMwVoC8B0sq1+XSqj+8xn00SyUw3gcDw+D
Y5ADLeXyz/eqhSLt7zQibcNcwSMLfjxgMhnIdBb8NDSa6AR48y7vcCfIXNlErkuC
J5AcyckrCdTJI5wokpcKSMqTjz1GncGDIndDSR/00NlRP1jPnQBKFFOrppiqfX4Y
Q/D6uMIMIympAZ9PY51fkmM4wdkyKqPDk2QICLXV6OW4rL3a8LUN7UNv6XvVtPPg
svRkWRfCrqPSQAp4YKxqS3qVcA5/Xa8FFn/W4A2aWmeTHOc2L1nA/s307m22NDwY
c5T/3hcDaKNEfec7POEzStRtJWISp2OJvQgm6DarUhoC6qhy55x44KgAGH+VMwse
zdcPw1xwWh7Tu+YXdyqLmH9zktYRqIBSa536zEzsUczYBAqmdTrZCcLYrrM5Fn7O
De9KaQOWcRo5d6mDTtFnEqRXgTId8AYpiUcl/yqjsjIOB2CiuYx2E8k30jG/HV3Y
uzn2q0SogjgRtQ6IxqsYWNAGBQEh5NVplNvQTIDzg8OsTQ0RIWBF2sVug39X3t0L
bBBI7qfTlEaDPyzyQRCreoSIBSo7GU/mBV7yOGysVRnpznrn0GjWAx7HMNi3BGiw
R7Q7RuytvNa6MmFNmK5LLPCmq5dHvfNKS1ew8fXXpO1JUFe0puwPVF2LYR1XcN0M
4V3yMdEnApF1hxXwSvaINaK71ybEmLKKZnyTYiUlHADA1NoPvQH3TLwYe6xmT+jT
jXCeMJ4WqCmnG/Ta0OY9fManDLrMhQ3PzZS/wZ8VWB/Q3ibRCGG9a5Xm8Oz2kHAe
fOHp+mFgWpjhFLtIU89TOQqYrA3QzWhulwI7uH/P9hIoYoYzalxBti/z627leUbr
uyc4sYTf/Z9C9dBgGFI4Umkxq2VPUDeizimls6nfTBMaPSScyfsk+r35MvxpacTH
mmpde1bL1B8qo17CXsvLlfz6uKyaOKkcYKS20A+KmK8myHbujYEbpM023ZcjvZqj
Ii5k6Rr4pu4rgqk646uKtmPOq1QdG5szgmtXKQM6trHjCyHtDVEgRvs2lTUq+PUP
OlumfkZ0VesqQFIwAvqgCPhGtYHgOFj5aYTb7H0uvnVnP/LJW86m6I2lKdQxVfxX
RP4rRZtJqOEEr2HzNIw+XHl2WDLE7v0ehY2A3Ghvdu3pawkbmLu65/RUjV1LgeBW
Wj0z94dSTBR3zsAsCW+Bk2cL4UklhySo3YirDG4Z2vGa8ZXp9WaniVLN6OpfWvdy
M4Hub6p3tIfNV5avKNFlgbXFkCy9JuXZNnrdaax0lX2rMRxEGDSghYFpcpK/lWm1
P+FgFBDdqNxorrhmQVplJVDjD5eNmZOJosnTq6MNjHkheq3CQhuJbu97IaQ90E4B
UyqyN9d6fFPimCk6cHO7f1IqR8zDpzL5guWleG29dMS/SVBIAdeRwPpz4yxVDcya
G+HznyDtJyyPq9qj/eLTrPod4y4VaxZN64aUP5btwbC+JEpAoJY/4Jk3tgnuqvdf
vUir0d0CoZmwhBZvRThBFglpSBDE3L/J0DIZbU1bhGl84IX5HaU01kpFbggW26jk
JYgkbKtLQ8oUWFA0paZRrAJtfKPUI2phKQrCBbFaFeR/jQyE5buZrbx/rrBjRLpS
m4AatLghbobyal+jqS1iFmgKoi0Sqf1RfGJWyC4Cy+br37i3DUakFzdwasMDa28M
jBC1bUPMSRLd6THGzjJlKMUoyL3Lz+m6Xxehsl0np/TOE8fuK4MCn8Yhji6LSYJD
fvfyIgfsduHYdPAhcRZAddskvHEA5rtawxS3CFhOBvIFVkEIjLvitXR/F/cLXiBx
jvGinKyHjYtIpIEXKUZakltwCA8aBg9HpOdlVFSSA4BfTjqRlMMMt0+3Av6mlx14
K4oJruBu/YybS+RmmFHrE4WVVXiUkvZHBgnQFvoF+9AiJ6IS4noEzt+WoeIDieNF
GlNA0KXr3ZNMP7OzNGAURcLTktOwpheAA4OdGadsw+ZrJOYp6IE0QfNpPOk4iJnd
Axvf3Dyl9IjW4f73MF34YHiCqv8mtM391j8aU81RT+qRBMrkomYtN3M9uDYTQme5
OmqM6wXK6B5UUEMZEg3AHdFPrFnOsrOW+m3Cja+kFzE4aK6NXyXLMeoqk3wwGpXo
j5LmuJLSQjwXvbksSX7K3BISahl628XHUdT8TPg2iikw5bYEuKjR8fMFWVtGMZwI
B7GD77PfccRGiOm80OI/eQQOjuI87h/DKI0K6kQFJBdk15l6Fc4OrFtrddqBPFju
Ok0iTBv3U1M8XawMHtwwgKhIOBIDCb7dMwUdbxogpYTUjiKwsOGpT/aSw7mAdJ3c
wFbP/+9ezZQZPDe6589kv9t9vTCb0HdI7T5hn/yQ4kFOwScWwDl58b7E9Wy4qLsI
aVMQl65lTYXdITXJWlwkjFFEe4/213Tz6QAIueqqLvnfzu97iMkwROrI4EY0fafG
k7ub8Ua7WMK1K35AZ4zmPjSLonEBblUVeBMcAFn/0K+KA89EerK8yC2FBrTmgjLI
Q0njDQG9Mio+hLuPOjmft122jLfYBmA7opwAgZ99vtdKABGYfkHN898lkOj17NyB
rp1G0umdTLiT+/ANXa+E8jYy2lT78bHKWJr+wsg2HWnapPbMXUaCPWtVsfVoJVG7
sVTBl9/sLugJvtKX6uf7NL7qvUFQYzJbwFQLqfjBzDAanLGQUceakfhQlW0F0ui1
zvnN+TqI5fHDWgdXJntTdBwE048JkjN7aq8IRzrqXclcYQ1w4kl5rQXp7UatMBGA
blX/njQ1g6B4S/BBGAMHSyKVUZlPJZyAjYb5JDr4XWYBZ23A2EDdmjY1Apj+iGUY
WZbl8nuhECVaHxsCBvnsx1Q2wxIwPL9WTWqwAf1lc4cXxdco0ho2A6mDsYUxz8Zs
bpYemu/9Bz5d28XgWOFKx16ILCxj72VMBUS38pV+lyLSYxy4U0A1PdSi0D/S5msI
v/fHvhB2c37KpAA0vaPeQleomWcd0gC9fQtZgq/99jpdW9DQOpVF20WO/IKhot9X
FcgonvD4kMBG80PNKQEXK/tOgj2nNNqoury9egIhHLLX+sPGpOzkWoRvS6LXmM43
0uUU3KLbIOOg/2bRHLPBdm2rMdTv2r/Cf38nD94hxNaotf0VPwRkmIv7Jys5nrW2
lZjy3+a5cBsX6aMkPZnv55LNMRfTtJNzoVFCInABoUfLQZPZTwz1EJFN+eY8J9gE
28IwnNI68WLTrUfzQlBcdGMT77QAwze4Ax0ururTgcdcHiHf5RQzS3UwdHhO3nH/
0CODSZd2H2g5XXFVi1J67N5/868u82OwCoUg865LG2EITPOXFvQf2AC7B1JblVAP
IVjqAZRCoz1HOrqiZRNQDQB3tar6TlMhya/8/sZltoQXsUZxYfWU/8Jd7uy3gdH7
rKlGk+VLEBT/Sv9kpPx7Q+0dwh7wTW02OpLSBZlJihtaiBuPDDrVMSqnXyocRCZY
n3gtKgyZiDBbEpI3QpeRoxwz5ZUmER9vH28W2RpoW+Or7Z4njRQB8uzenVTdui6b
CUx6nBd9DNAXE9fkOw4Y3xsKoifDRKL2bWYkkk9x8Ifa8zbISwaEsvCUK6YhJBze
CuH7J/fvLZdufmgdqe5FYiXCRVwikbpWHuYZbqkSh4DIB64RiAm55vh+WiA5mIJk
2f87IlNpZk7Lzl95kO5dBM0+7QESALqzs2JfZ94/PaJob3qAVPBEirspFuCuveSx
5PKqmHKXyKtYEenMl8f9YCspCLdwrHllaXccpxzHG0SNOb8tEXBcX6TU97KUav6z
jC7IjDWPyWTpOwdADKQbWMvSg/3iTLdHf1VqozqyzuF4KkU5nDFOaMsdibwYco15
sEW14f3ASkrrq69HLg+kmwuAbUnl3W/F5P0la8o3nhOxmuDGhitH0asU5AFv36UL
E2vz5WBD8cSUwC3GhdtHor9y9I8+0Fvyq+iy0l7i2X+nhyCz/Aa/deR/WTCXT1dO
HeX3fi5uWpgm4MQ1Y0Lf5kpQF4hmeyChPV93fRaYscv26WWp6JzcIikdEXEUWsoV
pXcFpKyfbUfx0YR5NTCXXvBqLhyYO4hfnUuHVsQ5SDf5GS8dtv6uhu4IyjSltKAo
uQ2OZbjtVJ7sCn3/XquY2qxY0+J94uS02rljuAaZaFwj0GP4Pl06gSEthpkS7V4u
HLW5YfitAMfQ2aBDqgv32Fsl2H+X0QLCS4gZvN0BrCkrb9J8L+LfCYWquUXF7D7z
wC86bqRZ1NMWRTfLzRelgKXrsLO7Y/69uqBrcGlEvhcAi/qbI5zI8C4ba/6lNcVo
3AQJw80ehF48xvLM8mI4HkVGuDyKE4ygVPTjJVPAUJps9lZrQDQ/Li40ybiEgxNu
6B/1/enGhI4Ad34+U5B/9Z7qBexGBr+KuiEFQ4txch7/0Y6nbsSPnXUvAY8SXB+U
kIPTuUwjq1oE6281PtGleJrfp2qdngoi5G4QvMo03m7V0Qhab76oM0Zi27dLfKOD
pG1HgS5ShoNmSVL5C2zvVqsWLilv88G65ni/X+1czXBYVf7V4f+V1152lBJZo4xz
Kh/evrJ931O7H7ntQcFOt3W2rPFpDiln1mx2QibjXQfIw5YHMA33B9REG5C12PJb
epI2oTqctt8nZsttUu5wjlv29HLBB9oeLB2D2iqyiRbT0MfxnNcOUdUIwKu1hksg
8DwIqsydJ5SBWKHEqI+S6k5c6cRRxYIn8TZaV5zifvBqaUtFL2cU/rPVfmP3DH3D
EG+xPT6bmzcv7ctYpWydoNrWWZzxgUBwiQB1Gxj13pMqQeGfid4nY2ozlt3eSE8B
9Wgn6MWZi6eg1jT4ve62P34MYrypJYehrTrf8Ph2xqtaelLuI9DCyvs6Js5iUTuH
i/DsrFnkGeRm2ATGk9hF9Ajpp2Mdqp0Vd7C8QQ3855PQW/MMBHaci/PFcE9dypyR
EgzIqAqetXHWlfr2EYN3SVKnyH+mX/tsOueUkRDyuTiuELDqPz3dvMjSc6Xjj67f
uikkSBo/uUT4YqGBX0bl8v6BWXhzzRQGPbHeqvmQgXq9XfsjM+lT2EZg+HDDOxWb
MoSrsI9vxkdN7KYrrLnUbZBR14oEFCxDU7WchACmm8LeesUnNYYZAKEarno6ocoC
87yC14UJCDU1bFIk0D3gybrE6MiPmNimwN0DB/CJBvH2sxYU9b41FCuvork0UWS9
Ym1RZUCBnzmSBBGUkPPcbAEA259hcS3B55dwxBMqPTuatmgafYCgRLzSQ1yLCft/
x+ZA5vbDULOclOIGYRUUw6ztQzL4TMUPKjMkJyHVIKGhCeN4o+FQ2WoqQG8i33iE
Zrw58OCNFCvwQbRCeIEIqXJReDM9s39d0UeoOUTC5Yymr4aLRIjpMkRBthZcmgjA
4/Glw/Js37N+02GwYg4AwhSdzGTXhhTIOZFYq67m2L6j44DoYxQ5PhEO6Em4MNjw
5bEQ0VshRmBJtyjQqQkDhane+baoHLpzkGKEpPxCkXI3DsombPbaMebqzb9CZOCI
ml1o0y5soR/6sxmYsYnNHSMjPTLl/IimFwK78BdKR+vh7Rn6wzCT0Nvwx9PSVv+L
6LANqNkKLUH08Ng3WMQPbgw4PIYkZzoKXS8qCFJwDTmg3pBaoWvpn0+l3uGuzJUU
EwyiryKwiIh7M6OWiVzki+EOvw+7dOcitj3TPHA/XZPdDVx31C0+KaShbeR9JlXq
TpkvXcpP1BkySubH/F5u8k/GgnEFmERnYQQmGWCADp81uyysLc2am8oowSDyrQyv
lwUbORd2aaarFh11sHbtHf3QceIyph5Tg88j4ec7Q2gtuwRuDoV7LHRKTQ4XcHND
le5+JeeAH0SyW1qdryAqgqjRO58wW7Ld/TgErskyFmwRPjiF2HD3N7dy/OqdhjTN
0KVYvAn4TFl1+RXEsMlNjjYVSXrYt05istT/pdWe8DNhkCHXBn7RCKKhf+PmcSyC
A6ILent2N2MC8k4JItXhRFKSfV7yEitsbU6ESa7RM2YDtpf26Kv+cyi18H7CryEv
/0khjCeu1PPC91RyRucGzlNrEMzDxGccmF65qIjbNpMMU9UNoyd1qn62p9rSb8Z/
f8tAOcYC2DWkOE2pxZDB/HohH2hlcomIYy3hvlMWVDJ6YHVLC+5RjTxP6Zpjijrd
XJL/GH+RBC0arA5n4lXaX4IdBi7iYurHjMjVkJThYQflBS4VZMqsBT9tclNuOct3
AAOZR+hdExdFb8tO/rEd8w3L+ZmU4/JrUvyG8VTfkHXstWtr3AbB+w7OLayqxrmK
4gotuKVlNUjlUWgSEEUl3rkEf9Mrhl8t8knYJxg6wOZvuusKzpCI9pxJRpPtUWRx
/ZX/oVncF3P5pEd4pcFEeDsXC2bVPD8Pqjx1VFCM7B3UnC1EjOfk4kahBtw88amo
VhhiUCcukrs8Qa+VfI/XiSQNVY3C0qagDOlLogYTHY/Wa3Y2FZ8I3DIziLgpA6Ak
WXdRI9BakSVhbxatXAqSzS8WN3VgIfLN8Dy1WC8QjX5gGOi7m0hJuHyGtfgeSXEs
pk6tnZ5hFbFESeOAWJJwtU6HFUTJWyvmKqdMdWMZPb5g5D2x7nmRpL3e6rgf/+Qp
iLCzWzAw2CTLc5IX7NhWjznDKI+8fdBPFCEpZ+wqvO25De8l6SjkE6YDgGfFVN2J
stEGVU17HPYJp6AOr1umwAtyPAj103l1kKhAHV+MtvuumX9ok8H9fruWp2xEjpb3
PuJFbi3rknme3s+yVcLPag8FU+Y8P5YQW2pHVWjNN9S4er7Pb/9Sk05iuzzXcHnd
aNzI9nj5jbFFFQ7gvIHimksrZXwK9UdiudxanXujlZvnc/H6SSN36sZIJSaFwTQn
gCeIKmVujX9WspF5lApwhJu1kO4L/Y5upV6XK9lhmEpep38QDGZgozp/hPUn8fmn
efkvTuQVVITiHqq0DQ+sE51eFPPWP28Ho7H1iE/E7ZUd1WbBQJKg+4dOVfj9xaGc
8YdpW2I1Z9ncOBJu0LcayLdqQ/1JaGf+Rmrt028TOrWT6b2ZjOFmwKqm1yruxfq9
W5l4rvCOwU5vzmDSizW1Z920LE5t/J3StGwF7zcjCuCaExKx/tmcG/oW8TTJFCmn
rVcs0G3zoqx28ZX1FYmVHbLFFtFNTwHF556MpCSgq0OJ5UfL4PjXzndfNt45Ej69
slFfH/XZfBhSCJ3tkWMSzNpX7OWpDql3gCbX1iNBwbkIyKwnG+AANkg4K56AXktF
OsXna2jryuwkG2mxGIDMJ/jpMq9iPAQ+BnOz40qmBk1NohldFCwTxToOCNtzb5Di
P+bmtFli9+DU2O2P2supRNFE11xweUAS4MvE1sg3To+Tm4oRw8kr4KVOkigLH0QI
2RgiIDHIoi3dqgoP01TodRKjQx/pj9b3B1a2k04vVtYl5FMphvGFhwna9VRFqndS
2Mzns3R7qinUD+ferspxBW/8S9H3dBD6V4lVlyeCybJCoxTdabcQVKYXYIb3LBy+
lskohEnFKQJ7o7wGW8/1XfdYmFMPUq87cVJ+uczkZM7TotMKJ/mC9BWsQ8qzBk50
71mgzx7++1tMIgTrvP8h4vg6IAJMz8S8LXIwHFHkm2LNNLJtSrzEttebqYCa2mhj
Lrwu2mU8RmIPZJYj8kjm3zh15Kgl3ZZM+wx+tp/flJZ96XXKZ/F7QcS6J0aEJvwU
ZtbCg/vpEdFbYbi7/JyYirKltGpYTdtYt7dtpxvbf2pucT8I499Tu87cPG+kulk1
sRtMOc7/nohZFqKOMDUaV04v77v0JAVSY5InojuzlLVK3lLn7WAy3gIHSZDfKU0/
nriD45cxEvMDraXkpQyIchSTOJpw0CgsowWbqf2sjYvI6a9A7Vc4wdl+gRFs1TUY
aRZXevCzNPzY+MVzdUyazFhVt6I0Jg3XUbZywFmrx4PFyMBDHHngILEQyY6Cms9C
6xhSD67GNq4t2OzJL48pJGLBk/s0F2mRlvh3bAEqGqh3pDq8n75sD3geIe8076Jk
Hyw6f8XF1hQ1kk/3tEUxaAFf2B/luUQ93SZJ4nIngRp1Bi6ulW4l1mrNanJKrHlD
O78hmRKuKhecwbgQyvgWV2Hgz6AX53hiJYRT0RfYMNyDczGhq2TbvHbauaHJs5We
Hqmgt8g6ii+rdsqoqo5GK/6lCl8PKQWtNkOx8Pvd3A1aijfrFmq5FvvF/Z3qNTvX
51re7wHT7GhL8mt96/kxGUjYrIkSwqJVPWmva77e7Sxp8AeqyItFA8rg2kg61bfk
Kg8NNlo2XB4FiBmVkME3JMmMzKAf2yaLGU/CeaKsM4+Tq3yo/8UznP5yxdXRjl+P
4xJBJqxjX6BkD9GbTv4LwQnu+z2LIMPl3skHtRk5+mTYWwUNaqw3UC22kC29LuAn
Iaxx9ETU0jxCUuKXuKKOp6BptaiUAY+pr+fQSu36EkZ6OH2qh8ExwEo6V4IvfUII
dKPZhLtwUhewnPzRRKMSBEXcSgMDWtlVZ6iyH5PkDCAG+D3d547yXaU16LerW3hJ
56b3jGp6wSxA5QOJpZw41RXAWcknOMah5dcLtuNvCvaXGDeGw7/wRC7ajJuO2SdF
txZFf1mkSKXPT9WHimJRyxCu7BOHR/jICkB40qPjnJ7nWadPzySfUD/ITD1Ob7Jp
LYk++KHnlsBYDXUmyAd5pZPwrKf6V1bNHavscQUxjd0EFvzyylesBoKDWG6jltDn
/mapw/7m9iQhkdEJsC+SVK7+jfaVMazUYQwBI7TmtcRm513Lvtc+cKrzbmDymHGu
GRgKXP0TcgoSfUhGDRPNqgt1ByFEMq24C6CkDD+LFNucKyTr2uA181MDnBH0YwjO
LywOkPBVplAf0YFwIupoDsyX02K8ND1T+nWXx9LcWLfQkFfyMiPacWbxsGpUquSt
Ae6lX7aGl5SxFOaSQg8sRMvzuPKI+j/tgiAGy1ZQAWnohuuAr+KuvX40kFQORTgN
OSgeLpnBuqNuEOVw7Qs1Phnwf9/GvYx6dm7HnDzRpaoGf5t0qP27p+ZlLuimWXLK
beJj8ZHwTTHuFrmxO+Yt7lQSi8reW9ih7DuNGjHMU+xtvRVM6LK93xVlK6iffsAU
tepEHRM/lhrCKwg6nN/j8pBU26zI9tPO9Tnnl/KRW1hTwDRvH8jtGipSoU9eDIwR
BRp2KtXGQNW7VNXqJtZdtplOv0CHjAcX6HTiAKQDqOqULrY79JS3oILAZ+kZ12vA
1dd4JCLhrd3jHPPBMHtv2UBoFTinUuX0soFhwYas7mzrPQdTSoPg4KMafk5HNocZ
5n+p3BqaMTqUaen50DaG+NhYUDCz4wckZuR99Azb8HHakyj1R9M4SoT/3WyhBJ3J
Cgnm2Y3qlhI4D3dgOGVcMcPCwh84DFSP24+p8m4/8CmR2PxgytTOQ5n3+KisvjAW
BzANHijDu69SUBh6PgyZ3Nb84zrXHVpx/ShGlh7O+Ljnk7lINtyByOifGcv2uUjn
hevu4x+LFnJP2Sc08xtBme5MnKrxcTgItY0n0tludy2Ni1IAfeVQo9YOhA1vfA9x
2hProBIw2L4pYsmhhVJjSlbEt/KBiRhWZf+L1wv+fqfuuRgrqDgBK52Kcp2NkBzd
xbFLNjC5RL0PrC099OY875nJFHMmBTq8P/2I6DwViiNXAQZp0jKpzz/8lb4gC0P9
/LngasYL2tJF2CREtFN9LE5HX6cjn7UzkzjToqhS2L1kwQ0D3pPv6XuqUyzZRKVN
tlbnmmW3rqx8UtjkUdyxaadX7ZzRVG2cI6CduSCzjm4zZm7yc4D21QqFWU2Jarlj
SCPWDw88AuT5Z1JYpMGT9lTdSTFItZw45EFIi9hErOY3am2X/c+N8+8m+fZA8LfV
jInEK5/sbfK9Dl9ezBmFwJ3HyPD2QdDx9qN+MyF0WOvRRbT3Ahp7dFlWNsR2ZZQs
So02Iz3scEoIk2y3AVU5bDDgAI3TTrCP1LEOBugRj2A3RJ7iiK1mXI2kbh0t0R7U
sxdM0tCBzwbtUzJYk5EPvJuu0+McaDOR1TB5u2opTDj8LEJxP0kUJCsDw0LaRYCJ
+XCGTmUDgS1Kpejk4JtLi3iDrBja78zFnfMON9UlaMvQLfyRnUa5hWNgdGa8gLDo
8kpUuYSiDXxmCPBNltMDZy6ZR3io/qopZdAWMhUbeLk3xPLqaHOo3E+nPI61RliH
C9/6cl4xHyXJfAw3B9xFUFtuwil6lphR1Ut7ITLVu8FkwhdPDRWZuB6r/gwYy68f
2Yn9yGhJ4Dewu5inStEJT2ro8l45VPSqPTROvTkGq/FZbHmftQZ55ueH9xgh4Y4Y
3Fhr/F3xPji6Yf9akTZA/C479dTH+R/qhK4CxXWOepIEKPJJffi0YifFte+zwBGJ
IhN+64UIqlZamJHTrb7SZMwkfcFcc8saxqXrHoFsAJGGfkP9KyL/MfNnvTnAXIaU
VT5+Enj8dhhEZiR68S28f+QJu5AGwb+w4pMMidf5ZMnlwRf1QhxDPwTqy2WFi0vi
TZeB5kCmjElCxWVL1jjCy3EauLt6CFksfefhuC/5Mu87zF+UuCi16kf5sWG+Xj8u
pS9GR4w0Me/Gd760Fb0/y/zQLev2T4bSbuG+FoVJU8F+ZiTuH7qcmg9P/5DbU2oG
lw68ZziOBoNKif32kfcTnu4dwjJbTpRWmyW8bu5g95NQwaoYZxE4Vk/sdR1SAg9z
gTTmW3CjecF4D0nF5KMOCfgSd3fcsqG8at0Pf74mY7EKEhHDPVCiUsNtZ7gPCb3A
66SNY+vS4QWOCD3TuwbbhShS0eCjkZ8HV3IsE8lr8ariKNcrr2OZONveVQfLWR01
zX0Hwsfb6sL9tBHBANW3ON6EBzSbNnvHlwt85MDLwzgedCdWb3BQ0u4fF9TXA3Ev
8qTsjkfpgC4kv82l+oVXJTJ5LYN/2z3gg2g9qRmkia9BR2t+1RuDFL5SAsuL3o8n
hCjJeQ3IdF5pf8Z0CXmWz23FL70k92xTMG9kRN7/nxnE3QYue9YmTLmzeXKccrTF
H3pRt0L9+lEsiJ7PfsQL7iBEs3Es4a7rr92e3QxXUOuaXuey8J9mnrDJQ+IZubFx
HPz6xKXBPMNDIPEJ6Vo/3ssgQgMCvf3ipq3E/Z4JKlGT6gHzzQCHlamJtks0B0rs
dqyczkmgGEekH9VG0rMP1IWy9XJYTjA0Le1HwLdphtbVSajT+XpKj2ePqXKRa/FW
vcA9hykg8NSwNloTG1bk/b00YP6W/YzK0eJ+TRLiS+7a3flf2+XY4ucvD7F8D3Pr
KQ0eJ3zaNwMYcowq0rzbNE/Y1jwk0JH+3wNPuoHWq/UUni/aujlTesMh+tiMwE/2
Y66s8xlOlyDErmTGC2ZNjLKF3SdSTANR5YAWyVvr0FdKjNsiajdyBKOj+5tkFs6S
8IAALd0QnbTyWYYxxhFj/HfC98H+wjxz+0ovCkxcdeCnN+5pDCVK6oE10KX7hi+c
H7enctGKNI5nK30l26h/8uyFudIGuhcJkEf3kcNWczqHi5dE1oIT6Z+OzoVg9IbW
OrnOvwgmvqxwYW1WI7duCZcjBGoGJcF/CgaHKB3wfe+cLqpvrP31Ew/eAiN634l0
vp+wWX4LfnCSy0A1HJmNV8aCLPM5hUWo+eWYAPhPGDCa2yODQJbMWFUS17im/6BN
cILUSStIZ+VTtl9+2OtZ2670y87fp/BXfE2gpzRxdeLMxm/9cgNuEMMtMXohhv1x
S6LvnSV44TKnHbD00Ubgnl7JUx517EBRVVtVWzgPUE8pYO09QLoVWkyRjaDcdhfJ
1RHT4NQL5z8T6EE7y/7FwugHaQOuESUWSe6yORAwayldjJD6eeYIye376UnckpyD
eaT2P91ylp+X+P1dO23amCuBpGVBq/twZ5vozWKUjKO0sIpx+3P0fk7P740HzLFE
WY5lvmirfcZp4B6jEJJzxSjvdaivyz1aHnyL5nyQZYR2/RTEUDTdJVDnP1Qkcwjx
X/3LbsR3msy/OyIpvBJexxcHldZJNpIu2MJRtcCyN9V1IzNgtq5ALuEeVGUzaInP
fSEpBojHz4eo2gTEmB6eZn+0PCpb63y4BNiqKtYYjA8iVJsnNDM7pduLijyOo9+q
dBKKpI2mwm+SbqEmkW5GJi5PijQt3pLtusT2no7sE+0oc1OMTGMPCaLViH4m1PZT
fL7rKbadvLeszHFR5YIE0r1JopYwW10qvqQrxAKuNfjzZ3AK6P/nzXC0VuUPIgUE
2CKWxwDFtn37YsYxED1HCeKMWwEA3wFKhJJw/9EHOSj24e6xs4weKFFAZhAH8rw0
6darT3jrXz4xd0FuDq3/FeP5LKnv+1cH1++5hOumPhtrL6ORZuQ3V38jNXeY3ywh
jouxXuTrP/Tlt5eDTVXINsqPWlpnz6YNAP7wpowa332efEs7yteepYgpr42cghjo
r8WqwmsO2YUC136WsH+GNSCu2CJihuRJvHOdbPxaK/kbo35IXGPYuDiaku2DlW8f
b3pMM8RmVm6zG/550lGpkIENxMqrigl4JxzKzTzTKPYAQFTKrEoeQ09YTtICi67K
REs672gV+FklwHVm8JvcZSUNH927mkDk4nkZWoqFUYLJoC7VviQzDfQzfuF7Jfbw
/0p4puczEL+uqn8WtfCCHp++Uufv0aTF9NOAt0VU1SCX4MM9cSoB6dhj36OFTW0/
kkGC8SKqd+4ot0ovfUQMRmy4AzkqTAF9npcTG4METJhcp8MaRH/Yc0NgplxSdq2+
zjCcjIsQqC6n2B0WeWi6O85oTU9NM2nbglF8B5jkROUQGlAlfZlao5NIC9pm75KP
bIGy6LZik1SGYnmwPQSMjFr7lbEUypi9VFqCWwXvjt1+Y7EFY8TCsrMuWNUU3I27
+7+VCzomRgT+QLLz4b9gGkz41CASnqADOXuEP9vsBwIf8iynv+1qey3RVTiQaQi4
FM4UkHTDzIwUFodR6lSLBZq9GuTJypKx4AbEc2xJb0VtQ2MpVr0TrznYf3iUEYac
fV1qF1tMkk/N1E0nN9BV2/657pOAFrrWHEGM6eIxqhb2Ew69VgyStu+hby81Yi59
qAzlWt5GIO1BBAxdvSodJj8tusOU9Q9DztzJqF4n/Hkj9C/BobVeLfSIRCS5Iy2R
yVVv0qIaSt2BqnVac4RYjtkjWxxSA+iJQyx/cCv5UMVEOEeso8y55J1uZBCmiQBE
ptEtcgWcHyjXDKv87A5bOq/y2jgegMVK4vfRAmaOKNwQtzmljPpw0JipQs1EVsS5
PHLPO+UD7m2EkQoSIEsbdcdrROkD2QHwEj85ZgSaVdsOn2DyHCLNKI6HQ3k267sS
7yqMM6Ydl7RTHet+PgLxWy7xrILKpO+nAgwXjv9z4iRT/4SPOAUXrC1DZ55slppN
O8DiG2SLc+Z3fLdY9JlWGR+jNFDDHoJAUL/yO7VPKxUpMzHehYUnqPUe10IO2MiB
PihVDRIBWj8iTABkeaD0AE1xMjiXQpRi8ianibWd5qmUqYDLQxuFWl+pPoCCluIt
XRKjEMxTp0Coa5ZWAudNmwg7mYXmNvAsgArGIsq99+O6892oEFVKMkMFPLKD5oq5
z9O+XdEQQVlN2ZmuiKF0YZqISSASy2tNDiE63HsPWREN3C3UKgtRsFrbBiaI/WiK
zpwiBTDEcBARKS6pPRtEm00tSMnKWFOHyVfrh+MlXQ7yEJdCPO5HoIEzVD3wxpce
XJK3dsSolfpkkSgED45tHki2xuN0jrNzsxOcs/t4ZaAo3OZDc9gk+X/xwgHfMGWv
Nvzlr+J3cFYE4UQbwlPD/aYhzgabdvb4Xa/csUZEWFsyAUcHdbCXcGOBEdFXA47V
z9fOJEBGjnxL0pA1WzTEHzr9zvS0/WgpkTCo2JLdDPGdluDDlx5969PTEkME9N+N
8JhGvCArtlQjlR8KrA8T/4wMy5aovyKbmlzWAovx/lwL0xoGmI+4oWu/MH/1rlMT
trnL5eTz11wQ5Vv6I1u6669nZsMxzvek1wEKu2G1fDynval2/hlIkQJcwEeTs+8p
4ePC1oCu6eo/4V41kOjmHsSMLTHY/58z+FxpxaR59AP59VdILB+URVa1QPXujJMy
wtQZeUK8Pp1CssLip7NdkTJ08wrB5gELzuZwjOvyM0qieu2u66MamXXBo7x86QzM
8P7qUzwHN9t3480OZmjqXihl02zot103WC6ypsPbQG6rss98xnBHBUR3dL2nhbZ9
ilLlJQIEHDK7KCBgmhYr4MjCblmv8cZj+J0R6JY4/PyTrZ5/1dFR78naK6oa2lEg
+k6Jnmx/9y3ZwrzbwEwmnAVHJjUTzu4m2MwgTrLjCT/N2ycq0/iDFEyeBGOjVI3G
7ro0ElyHjk4n+QIlRx09sC1TpzcJD8vpwxjxO7QhFEanpwZMjWm/6xEMNNbqwQHu
KoYWqa9U8yL82UwkWuWn+IKOFA14KmOznfP/DFZe7S+X9XtYjldIjDKV6kpbGkVS
J6iMXvUGFEQrzbsuwZLaotmETxLqvYisv/WGiHrxy4wZwpDn7ePFGJ8hRMhlpF/V
bq54jzu64xdnhzpFd6Np9DRZBTnwMbGT5lUVUxXoq3osU8E9Uz0jpqVxNYi8G1rm
n5RrZscpfQVac9FXOqzQVR3m7DHyDgeJmceHx40fqfujJK+tRYmlgzCHyKKtHzN/
4u0Ymr/ya/G0n5VncP9+XVcc2Tl7EvCE5T62+9zBB4jdOFqRvFnyyCLRbcKjq+mw
qaiLb8Z1DECxCsUu2mIoFAC4Eqca4LAk29B62aF8XtKBpn2q3qc0AU+3A5K7SMK/
toRpYHFmJog+iuFfKYmnbiY3J1cXi5L/5I/uoFUmwCgrjI9GnMepKCFb48ARSDZQ
DcsL6GfJeeyDqqpsrIotSkbxffsAYzoJKTEeelE/T+PG48i3gNQYKeDXor47n3n5
99/yIs5mk6XcyyPcMeFFz6GHtG0sLyc2odQsHbfrtaGubS6vFtuyUNGorKiWtS7U
scRnGhQG6QU6gX8yGF79PRyzp7uCN8dUKmw7lV/x0TGnrfWRFN7r/ZvL1iQkXELg
OjaArbDy2eawSop1fKdHoJaDYMeNDkNS4XedugRfPk9R0iAbpwB34JJAZkbVKUhj
Vh2eY52TOHVppVhk95jIVd6sE5ujKHYkTMfb57vwL6JSjq2H1UwY0pB4svXzf2jv
uY0k3YUeIlurlYwDqguCqZzIGciPuDXhoAez3Y369DndBaonT03E87HoIvCcDyOu
gYfl+gU4QctV1Rd2S7cFsu0vsEbeQEqSUYmrII4rUPxmONwlKc1Defy2semSArQd
8BtvN89CFIKVzWbHKmJAJYkENvC8NMikXYlTq39aNsxWAE7xnYGCK1nCQSZ8GO35
P17/MG1gLyhV9c5MBmtjT+yCA5GChSBtuiSMievuC6/9iEGmJ95IEtVlTD+Woxj9
bD5KEaK6ja6u8CUeMclMlCyKSV6xHNrOz8/q0Xts8teuIIl1MOVPqfkGTkFyvuF6
8jndAZefEVCPbcIc7sGCMdYrdgzpV8iOOo8pjBJDIBsWV/Eozx5onLu1BBH7J0zr
3l2s0ZI6ICoA8VAHI+6voME5VGipkzKNUL2F7P+NUhEjmzZgXY3QLuwQpw4c8Ffu
Z7bDRaJ4zyg+0CTdk4XOo5gmo8ulppW8caBeW1jDMNEGn5ZcsSkRTcOr5+2iBAnf
n/QTDRHrirGWRPhBnfZ9HlulEcPM5HTl/GWKG244A5N/vMfu/+AEODSPh75Xi6lA
dWfCD8MoCam1+kQ8kp3KH2LIJ3LwS79erH0XiAY7qR+cTlfu2XTqeAKh8B48pwIR
j87kYiRLceAdqtble7JqAvTVwR5oZ4aUvtesLs7JPXG2LCCUKz8Xc2aDj9B6+AcW
MC0k5tvGNrzE6uL4OfhsU3iM51w5k0u9SPVBeZOvLykLCj4ITvzFBKEw+Hg0LpFt
1MSZFnp4+fQ7bRNwlQ85QowJtfwqMK6fGDb6KdwQWtE4T8zdZ7U3U9ALH5dlkthX
ZnLZLNPYWQqsrXhZoyx1JA6jsTKwTeV8zdJ9daqVungmtYKr3THMhMPpvaMCa+vg
uNYlC782V+DLQnVKmDkmY16EO1xCA4Fe7/UpwCocvo3QStGeyOVxqIq0k8Oqc8QH
7nqBBwgJDGGXcBI8bXqjOyOtHpXbXlwgsHGWw3tco0kc7I8E5evYDOi0ShejOYOw
IlyhZa77F85/wMo99gOjATqZ+wqEAZt1o/7avJ5SKzoKSIeNwyjrX7dwJMMJhFUW
HAZ2BUYUjur1q5wjANzjScsSZwG8ChTyUrhWQkV8ZsLScmXn9CN0s1DxotBgzrg/
GMu+FX6xg/64X0NiNbaT42Cj0VB9ULONe9MHAf2e48C8f0nZS3qrelj7Qn3QyX8g
GtBQX6FEZM1USYIuoK5R+2aNHiiUeSfJFbumnfijLX71+mCI4GrK5fq0OVc30ylL
wuJGQhiTf/Nkt31RcbXKwsMgDTjwJU1qeTArNgzcwZXFTXk2aym97YVqw5WVu5W8
+tT45bHtkwRTyBqCuSJB5TpAeWap1/U/3puBmZx+68+c1qjrgTBAjmZJbU08k5x3
7kTzbs1+qwFgTsgCE/s5WQAjgljrZlLDw2/J5qt/ZnVf+WrxaUOO9/Pnbe55aAZj
0/dVmE2H4Tx46tyxHpF4Y50ydypvjsvY2QphXvGxkashtWO6JOlIvk29zIzBAwQl
vj8MKOA9U6R+lIDIt5YBr1gZ4MVtTRdwLCAsPh49nJWmXCFF2zWuceaMJihR8H8q
bgvF/y5PwUyBPAGIQlxd1hXBzOTIZm4hfxWwiuwdNJpl1XaJs4XTWpw8pJmEae1U
rVRgWTVh5ReeZUm/tpdcC1QrskRf4ECplYKLXcuIsChy4GwsMsJSI2ywThRT0yqG
LbCU+IVM8pJkNTGj21nddq8IYXEzPRDy9nHIzyTBG18CaW1CVLg3THEpiM+fauRC
UVUWQeQxuPf/PlIK1+czDzyHripa57jd6cgyOzGaRdgU4+Qf1wQbLkiTYFPn07vx
B/59hjLPr84HSmvzmLT52jPW0/o9OUyX8btVBKN5BVytYqeRgU8s8S6OvuZ1oH/y
9jvyxR3kBArDSgvrT35JMrgE7pJT9ffFusYqesUSZPNHl5C5gwYn/2rFURJXzF9v
PbMNlLpePXRj067t7xUHgxb/wSymHyQX4wSSfxcIppmNWQYaOyDhEhCx3gYNcm82
P4LHr82pV+SC/lH4gWuFGzp6O9R9k7kA5W5gD6sHJbdwj1JMCIZvYfxYvdaqqCrE
FDKJJcyAovoxhXFuy523nTheTr8TKyfiz8ZyrnCh30g3eXeitXF/svKesMFi99xJ
c0cvka1+ikSIA/N6o3jFSY0wX5dlskOV99ndiK3MO1ce40BHGl/lEXaLVYeYcSFR
ZPpgztdsBdSsfkavLQeGlBxZoWy6v/dQexcJazOmIfe/zyoRvgffmcKCt2O39m9G
QiQ4HggXqnlgkqnk1SAg79SuwZw1nSthZgNrbnAJvAWt/j4qqdYq9YzfANfw5+ME
du/GqKHGZsxACZglHSxagd79+57+VMIgXTIDVImszJBqWhBEG1lr1rVmcTjfwHXw
bTbKLpfklgUSngBf86ogijh8Gza8NViTk6uSy7lPfUUSvkvS128PzPFcARBMZX3V
UEWs1P20SdCHTP6nnHiyMh/IeN+R5mejfZPtmMBLqnWRa8aWjEr3882D9es3mNC1
07ghT6pH+eazobMOLzIpxP1eG43ljZnKsZhI0424oukV+pawjT3bRGNfIt8XORpp
zNdaAEuLGKG04F/T4fm6cTs/6tdYG0qjHU40d4guVnyjToll8kU9rn1sGn8V9JzG
j457TlaT4NyoyrxSYLAC8mHoJMHaevF2iYIJ/CosXtOTwoHIreyI3CulCgUs07H8
XCaNUqmh2YgtaeHsTGdPTZWrqZnxdZfzd08kvyYxio+rRuP68ppjuy7pQ4zQk1uY
woGvv8Evj/Iiiyg1hDSQ58VpSVnGstZ9fa0FCIBBINlbzF6iruZYDqbCtVmyS1xh
ckdoIdD6uMGqvwMN/9rVkMnI+ZVywGA5Oy8mbFKnC+uNUwF2dFQstC4hnS94e0uE
J17HL+h19nHeYvYUV3HJ8r5gHhfCCoaly7QMrkF9GXQ4mTm8DQ+x67O1JGOQScJY
cT1+8Nhv264f26IFE8fupr+iQCpb5IE9bZCy7qQ5Czp1sTvZYSKB1Omtpm2yhudx
2gT6KiLoNdk7rhJPl7dLyzs2bDQEFjOsF6Zkjj+bo+YYnbpcRd4f/Rwwilyyg+nl
HfTcCTdnmfsQ1ExToCzc6JEvAY1SoYrL57lYjNbgRqqpxY0gDa3OjM1lM4fXGjsT
/uHx+IkrE6YOCxcYb9u13U84CbX0N1deo8C7qoywxuPTPFZDRfBh5gWeb7zY4ZOI
RtyXG4R2AliPWTOl/cnBPXa791yDqjvAxFTH/VQpwhvCoxXMUPTEKld9b62S6Qbs
Mn1GiUct02AabTCGPTljSc13RbFalRUq0TDhKHopmt9g8ynohEHE56cPPkAu9od/
+JkzHzr7dSx7wH/eu7E7R9C0LUv/M83y9jb9rFc3VxLS+BC0tXPkmFiRnEsfxhdC
/FYGB9Dl+ugVrPavTL0Gh0mOHqmIhDYNWHBP1aVLbeIatkZaIwQMF2POX2C/2QJQ
dkse0X+9TdZJ/bf6f/QV9vFwF4EaDhfUYSQYdbmupcClYamloavSf9em1aGuxd8e
0kOW7MJ/r/isAFLA7IVIjeKvTEmm0VNNG57FwLKyfb6yRsjp7uKOfGTw/5/tbr+r
Ujxb0snAofSindWvHsFghBk2z5GYdKSvSv6aP6mqrPkKJH1oKC9+53wajPlanzYA
VDcylfZlG7qNtdhUmVArTHrEWtOs8TzPegF05TZ5CfkTmbcr01Io8YxSsoGuRRKP
7SHArW7E7nhh7GLhvS8yjQikRCuRxkkMBl1dWYAtIAPdnnWWoiq5xJ5f0ZpHtm34
nNfV3Zj2Dx72tSTvoyL56qCTXr45BijIk9Dw8i2EG81Vxvf40BL9ylfuLwQJ9/KK
rTi/Wo9G1zFq/NXXr//lnfhGs2ZF7rzTHzFQvNt/v5T1lXUKrDl1BV/kBGkiZRfX
eIv206Bw/n4UG9BpZvCYbIgs1ZHf2c6UsdZDHQIjhE1NDB5UPhKu4ZnSFOvjSaBX
sNDaiAZf2EWLHw8RpxaFJvDWL7HxxGpmqFOp8a/OZGnCk1ktMVA0G4l6vmfTwHFt
vkZWZ2tDs/oEUbUAjHLbTi15U9Z4JUJRs2EWBN06JvS5dAFPOCpMo8TjZcHbRGBo
Fe/nK3UCxQ33ERKxGJyEJCytHRoxZ4HkARJB3s4QpQK58GUL63jnn2skyIoafbaj
d16vY9tQvpDX1zf6Sf21hsgy6+ZucKLNrECGqVydDLpFuwFGhVHnZ4gRkfpZlA5K
W2vGwQDps0XGrvAs9f1FNYS5UtfVPfIKpNIS3AzC7nnQjvtOJbXG5nvmxWA6Co5I
KqMSxaD5yjjJoGK2omMWJf5NtT/W6Ni4M5mxIKWd7Yz9T966K3LnYocrIWB8eCfk
iA9GkZm/TdKjo4/UMZIc8ueq+vlvYypuNvrF5orQIOanSZcWXSQFJF3BAG55NWO2
dMAqfuH2/AR7I0G5L+6Xt19eAQ3qr5itIHxQC3Fz6EK6vrXg/WK7tes5I5LjSGlw
ElvTFnex2aRZgO8XoOOFevCbelG1MJNlQf+nhN5mtyDRQ0nSPSzLHvvoYISFtsBv
JKHauA83ZYPjiOh7+ZrnTFMeyWhPEVoyKXyxmmLdvstXOUfoSgq5W5e46MAK0BTJ
kjRI6a/OQmHR0KGyHeol76uy9S+kSPTxZcKc1xlrbOk2NOb/EgkpoYwK5IzEZD0C
jO9nqmlq31xCBia4j/uMaKrOeoJUIkQ1Qczf3vMop1jz/xshyt0SLkZLd0mycK0M
UFGYwiyGERvDSyWJcnaZaATfp1Q4m5WOo/S7Bps4hFI89S72RgPrftoI2+yqufzD
EhJiFbNjDBE3Pyyner99vjPksAuDbibLtR0IrpXj19S9aFVGKgi9fBWTvUtQH9H1
Vq/v5uNbanEIUMs7neMT5YVi5axh83fa93OqGnjTnua2kH6i+t8c1jkivci1ly92
tUOj03T0RtsYvaoQvRIuhktHKmm5LVQMPxRkiEUMPj42wZbN9mHrePk+TIXwSZj0
nHx++5EOtvDc8dD5Hjn7EraEZIDSl41hY7vd4XcnksMZtMPvpYORs+mxSqSHPHF1
ErEpXYYmfoE3rHSG7KvXQHne5JZUdPREFrIro8HjNW1cDlbG1HiWBcfsX4e9omhF
bJNAGL8wyiGCx0F8XGZE7RDWygPkAmg7yotivGgZj+4lrgtR43U3Qr17iDj/WkYF
jBbXPbL0ozm5nhVE4uJixwHIAxUVVe2ldAVjL8tDaHH772tby0r0iCRlIv5omZXW
kEsAZZdjbXGN5P5zB7Gs5g/hJ/V6Wu+qI017VNR8IoLOyCfLTshGTTbTJQ1LpEou
9Xad6SVjK/oSYm7s1bUMwkXpmCPl2LecL6yjqKFyRVg5AyF80a+S982jmQhMdslz
eayBJk5wlBSjqMqDYz/nUi9e2HYBV4jsNjMwqYBuG35KK8vnX7xpQ/0vreiSrmgF
BNITNDHhUgGw1pFZz0O5/kr4XqxmgOBemUdvzieogmvTJK221J/89Vt7AWPaxg6R
aqmgGjDVnz31Rk0t/Co6qxRkHQrkUkqDSaqm1+CfJ5pnJHO8dmnpdRZU7kgn7LrU
L1SkVB/ePI0baMJFN9U4piIF/GCB7xe+uDWLrwgvavehC4GlLUpCnw+FoBqK0W7g
xTz5Zy6n5qCPUilm/VWQd4Gjpe1Z2cIsfzgdnqrU+jECvcIYBXVybunlEf/lqelE
Ft6YSnmLfFQMauY9g7MG9bROyWJAOHyJnSinOPuES3Isornwd+e1yFi0kwm7gETF
GK8L+XxaOAfeOyWwEu3sArxTeqCcQK8XwHsZzQRhiFaN2Yu/Zsjh30OiC/Qor4Ji
N1hpihy8TmhuTzJnsDXoubHVCOqKy7Z79Cc3Sf5YKik1KHlaDx0YwTH8NLhGpMRM
9oWRjuk98znc7g699NUvCqiLIAMeNIvqxQ+qBIQXO+sPvv4XUGhApY7Ed6cGubmZ
Dx80mDMRNP9tiE9P+TFM9Orqx/UGHSJmH7KrN8mXn6EgBpkB5n8LihX4F2P2+XYb
rnHlLGwB2j0aCtroCkX6gaKFbld2/KrtWlRcVJiuvVtzI571GOhNK5ptFmZzs+7o
jnd7V382Hieo4YfZlp0OwM7Rzi9Kk+nlb0L6iarkZfGFcEXhPi86gG1iXGrUdQBD
aOKZjUn42BjzHRUeEOqgsR716HIG1j5zoEthwXLmhMe2VR9mCuWwzy7mqjq1gVvH
NFApY6gvkYUysuCyXB6QV5UwvWB/mHk4hb9NHj6/RjBgiBpuIEjvE9ReEAkQnnBU
UL7E0SSxcmNhZ7Km6SUQlR6Q3AnlyUaXeU08JcLK6koObTwpE2tWle0gMzNGD/qZ
FylifnRKkgms/fluJEaIVU5KUu2MLuAXHG7vG3J3UbXK6VmEX6EXO7ZTYjF7kIOn
MVa5CLIHPABn7Mp1O81B2hVJX4UOhnNP+sdJArHNy4I7GsS0esJMl3frnJXGXS7p
snD/8pKAdUmKdOrRXKoxCXbPxQrLo9Lou9TEVvLKCyWv2RQ2NxwF901hBTnMDeBB
hLQKPNHoyAjwtf3eWTGebhe1Qfse+0SHTG2A1uht6Zid7EToljKzET9yw/Oma/+K
l/zVjB1BqpyaYJSvuLDlhF1JSOWwA4w4ZH07rUnua4gI6IlZSlGtWW19kak4GFfk
3PwDwvrwvquGV6gV/7ZFEbkN3gvBIa3vD3EkU2t4XHgiBJofRAe7VIhxIa8PTR/7
wk1VDtbKOOXN/ExR2OmOhALXkrudaoyzKRVXIW+5LXc+bkL6aVcNUb/WvxxHvIZS
QEXOz9h5QHGzS4n2moqEUOVyv/rg88Zm4ZruDEUZCvks5wU/mJ8GKT/1eHxUxaTJ
VJHYhjjE6rUashff3D+FtJ/P8lzAVbPrhQM34oSVxlp/g611hlR84gA4xrcfXKkE
/j+c/qCD++4szxCxSG6To3XdFqwqndiRfto0CMxqs9ZDtFbYavAEYmqC+x/O52Gs
rgGdBdokhgXYi1nH+6E1WZYac2rUlPFSGUhGimrRENYkL4PRuicZUzaagvE22P7O
/4zJzM6qI1rPqfyyzSlKQZWqKO2Htun/ck5mXdqLwQvhqDzzY16niAfPZOQEvDG+
FCl/2bnkZcxM1QL3lDQcbMfJ3HGmkTYoTjorZtF1fjEAFb56rZ/L3b2AS321W5Ah
4lPdnbXK6uXTOChDWdrEGntIU6ayDrQ6OvCyHF3kmarg+AZglj7e6YfjxjM312fb
MRs7r1HcJ64MGGc7eJX4rRJKUQTpaE0A1PcKO1KPlu/0RgPOnkFJceCv5o7l1Xs/
stEJ86G/gB4JZKu+HXVOcbC+GKT3Die2viM1YlXgyY/tQJpeyw/2JiqR79sy+nhY
7qfp/mWcoRQ5CK8GAAuyJvRwdJAZVbq1w57Z1WLCzfXj/x+f+Ezm099SXv9bxZNL
TiAmsxCuiP8IUu8wV46HJJytJ6T+HYGa58iTQeqoF+6MWHYm7U53D4YTaWqk0/q+
TPBXxfWyy5UhxnC3r5PDBkyk+4EQlILWOjoDUOxUCQlK1qSHeWSrCaqYr7C5swVr
jc9FTV0ATL4uK/4v+ZNTP7C9riteScdsMMRpWaJbNlJNGPr6XsW9fkOKbcAU9pvt
Qpjapz3zAR52ZGSltwbuPl6K6d9mLwoRimwHK5xebXlNAIqGhw+wbnNhKI1GwsGl
cZ36gmof4NlP1LJ1y8WWFbwCA1y7jmvc19RYRl3INlRmdU7jS6g44XvXzvfBTMFT
1mDoMeYuK08Y+dr6Usmi/mm8xj0OoM/jYQg4qcwIxP/gMblnv3XL9ntZzXp9yBD5
rpamcs6niBt1WERkvZKR0kwSeMvP9Bm6dxPwFnLhXL/x6TIcmr++m+kE3J4VB9h6
TyaM7ut77VY74/cZREHRqIErpKNPLIH1C8JyG8LX306ibuKEGeCazLmlLi9lyn0e
g9JpdTdSA7eIhnfWCC8LU1ClHTe4J+j3ULMW7g8EG9ZGz3kiEkIJGY84dGn/BOxl
yagQlI857cixFtR1uptzngMHcVR/DfhT3UmSDDi8DaZjMLoMb5oGErQ/RSOMPdsf
NZyCYVtFUl6hrkL7SR3utia8lQPGPKBxdqlxxAvoc8lsRojlPnnBb9gMrF6Mmcrr
GQHfrVfFo6gv9rztItLWpdsCrpFKMI5oLAOGjy5sFVFupP+h+XICqBPPy5mkbW0s
UcBsVJ5ycWxkArjqAAP+9VrCtOUUcOWyz9kRoWfn1Ffkh2ycObn11sUcwJH9+yaE
ZDUzNlOYgCDSVO1qUKHTwKogvTf5HXj9sVUNCORvYT7o6HqkiGn2JHO5YOW/bFCU
FPXmb2Lq/jnNwpFYf1CpHtbiKr/fBwwxR+OLkElTOv7/xVPHA4sVUd9fhOkcophq
vL/eCf2BDltFdfQnmCqEwxlg7i64lV6cN+/HPOtaADoDx/NVCfhAhCfbthhqkLsZ
Pp+csshNR3x8TRSXMWlACdUqxnW/otuCUYartqSmTKyvk4aW+4iadPy1xmo2yx2P
G+OVPMfJfx2S1MDgxUK0YLn7gZOm8e7v/J4NlIWlKkzkYqkW7moe/qUBA2JOSwED
JYD9kTrv7JcEEb1oy2Hy1w/QUyef871KlIcGCmQA13sVo/aKCYfNq6so488PWGPL
1CNPhcD5arZXRyYFp/kol61pgK4SMmpbe0IuwTbKi5jZI5ufStMXQ4B28qCtGLxc
Jz6Ggcpt8PIjrDbIOzcGGOAh6M+Lq4o6PRTyFbCmACvr8jeVeOVgktr4OK7nN5z0
e0HRhRRsDhFB/XoT97qerSuDmt3Mcxl3tnIsHcYDVYGIjn8z5BWwy+JFyfK+NGFr
gChq4Dy+n45ZOKisdY+y4hcKCRS5c+pUJAc4hCZs1ba3BBxA99skG20fh9rOtoDf
N+NSONKrzXp0/I+xbWKYAfxwwX8uusGs1ZwyCsUfze/6ZKmPsxdxbdMmm7nsfqFj
RGNplRAyctjAsbJpfZMl9EYy8hCwBz8wcjBld02FN1C4Vo6zQ6cjUuBYlVOoR9FO
k57wYE3hcgPTEhlP6VEXZVV3n0iJlr0yBLtBLPM82Ilpv5dmq2KQyh/s5RZOER/P
IawbtsNZnad3D3/7h4mE8hePqdy969mqxjgnePE7ZySfWtqF7YfQj99hv8qJqFzr
aDQffPEpvpLicZHeKLf7a99eArWZG1u2GpOYT+CsvvBy3+n+4N8v1rrjfS1Z1SJG
z0wlfiWdfQQzslqHShx5pLAOtVm17jlcVQfb38+iHq2GXS8FPztSbMWmSlDjU2/j
PywUfezxeDi4H8EHfAZxRKjc4AHni92QAfNYwOeMi2Sl6bHo2qmwejKZ6XlBKwRc
CUSlV1w6QiYYL6zJLVy1rnbfD9jnRr32r20mL74lMXqZC+9g9J5KJxAURrGHeQVs
Sn7TtfTWE9sAB/eixeiyZuZYJY9Awg6w7wf4HxDE00yvAGXcevzDZmJM2aslO4yL
dIsgiC/OrIL5Vuqi+SgaM3OJCK+9jPyzWAkWajA9u4xu9BXGQX7AQmAqIbYZCvq3
EfswmllzB6qFdNni/nWHUGOSDEnaMOABab2wbU6DTvYO5cDpNUSeR6HY7EkwPAeX
vtgPRLsYgxB6rhu3EeG2sOzM7zvaD+6tv8NnT74hjrjcAHglR6iYhcAB0r/m6tog
gAO1f5V8BxT2SP8fLNcPDsLRi5iIq6N+jPzf0f4VQNOGh+RQiJch7eu9trymrFRT
p+fpAYiqD2I/e0jW8KsaDwRVNqpK9TxiYrEMQqsp8aAAVX9QndW/mNwm6MlhQ3NS
TQcNNt/dJUCWvCO6eFm3viWJjUZ4osWYHq0aActsBI/H3TP1KV8HWgWv4m8HNfkI
D3GVPjfXovhTcmq3kzAdjWUgPmOFRm5h9Csf+Rm5w+EJQ8kNtLGdGfiLht7jBOQg
QE3sDP+XSN2sI02r8TXbgAxT54729bscnhpWccaUNNbuhdcltio1EZ+9eG8leQMN
ef8aJJ0NlLWZGkVyonL6+NMk1stUaK1vhm96xbF6JCaa8Hti/8HEyFPkkyOx1LA/
xR3Wg4nEFK21Wy/hZ+uCSpaaZk106fpCxSl9mQ97uWXB4la1quWvF0h8tZ67dk6v
Uww66rJCzXaLRTl4Y5XQVJ6VxkRqKQKfC9/3XWEu9dpat+bkyLhYYsQOdS4CdYyZ
f0t48yaejWm5SrlD9819apioJN9t8AlyH/KKOQ/y8T2XuI64eTBwo9aw+PyLQEXg
0MWAMbUFsTZkWCKMdf89OV2LRoi1mHPG/MshZhOVoxme0XSyUdxKkzWgWOf2r+qQ
FPL14a8CD7gHJ4EhRzV8542b5mMoGyKcmXp3V1GRbmVhyrcVa44H9iEmi7t/mMxu
/GvV7+rGN3LKV2OipFgHHCfnHr5v45Vxx5n3S+6+ekWU/Fmv/rW7THKdLdcRL8tZ
43OdrdKK1hZ47ElPdGFLBqdbslBV02Fa8O6ZGQHtwKjtcDTeTHxXQpiDBzuFEFDy
ZzkTQD1QCzg+rawEMmYHTQ1blGm2jGmrG6vKZCaung3ah9N5+jXEzq6H8Bn3xgD8
8TKKY2JKUCTuSx4y8W2Zz7Uy/QZvWXyPHJ5r9uJAl6v4s58fA2ehWs/HWnpLF6ix
LqXVvw1kG3fPFgYlv0qgmClmwgjPabb4svlKwhhvF7V9Ilqr5WvFJmqAXH0cRCAz
ZT4UitNiRlr2mMzzd6CKowusQq/VYDq81mUKb96aYq0+efJjqHSpG93p0M06Hh2I
Qwu+JTUytasYAjAqbjmJc8ym7XHJI1jXRPBfVa4FkWDgKzEfefIS6KzsCC2FyXjf
H/SDDy1NJIarW6VomxLzoW48Y4jcncoMtXzPmbAPHO+2AnEby4uvXR3gQrno+UfQ
A3DiHa5wv3bkdSnKdXerY8h745DitOazMUgPpRJ7oWvtjbL2noGqzzkHKu/3e2Ux
gJfrptsOWwLEQD3ldkKR89HX2MMks7Dmfmastp5AOE+ATsBtFN/3Q+NfE504hIjY
ac7su9a3tJOBtZ4v1QqjeckaaB7ihWTp6WDY82IndabguqeOQOG8w2qD6+YOKaEt
Lrk3UVby86kLTiptgL8UUm7QxA0zDiORQer4C7T4xhzZhTKONwJaeKQH3fSG0CAG
jy3lFq6Tv26qXgRTdQkT4QTGIJltC0/nKr0eChuPFkZeswIgFR6g+U9AdfMntUYk
rtJrGShQpvswpqghmlei0qYsIe9SaqtpMBvmF5aIH5vbfFRhFey2EhJdjRQ00CCM
r+II4Dgs0kOjVko3OPVpn/yFlTJwIaiuEd+kTco4B562si06UsPXTpkNi4CKLOnn
NOPW4eE/6sWRRcIlYr7oAdlZuOKSut6wJyupKMOscLvo1wIWaIsXoJf2/1hfQ85b
C1hs+rxud7/fvO2qml6xNJgFTC31NoCbzbmh4PXKQ6hIJRyKLdIGHJQ2WR39uHB2
0nrt1MGqJMFslFc61aoxoNU7mpuDid1ss2LCyf8CIPMCkFYrEdC2hVBu1pCEeH1y
vUGpGIEWg5U7uodlVtldEuzn9BIgnuL+A4oMVYzacVihKOlBviMHK5ZNaZuPoAUe
+r4TPnY1MCYrbqaCyS+/l9ki4YXN9ccCg1mT+DyhJ/OrSIQ/yDLzGYN4SsW2sIoC
9nWsL+CHaSrVCWKa5jdIbKsXeArxjTmrtwK7fX5IV3Ey98oEcXWIyOCjTX7f3xfA
zLOo+4KUXXWnXx2UPe5o+/K/pWwG3dQ8GGVQT7DUNjxYdVU8qyy8vPZQrapXJsgC
5pGmYzgPa6ZbBh4NjsSzOXaq5S6WV2pnumktVHFMCH3aw754B1FnFdZ6dAfeYY9P
bs7E2fAzG40v/v57LeIswkyZttbIs9RQMY3oecRjW5Qy6+2MePJrAPD6bFZdiF2v
LeJeeaKgiPHYzO4WM9VAhMaVSPU/XfmD57mW1FE8v3pdeqrwuP5rnjcT53sC/j8v
VI1ZgCvzE78BjHk5SG6UMpdjpzRuiDcMiIh915gNmL3ZWjPUB5A52I2aivcG8OPb
68GjKf7kPl2tjU0LA7VilE2BPH03QMKPovjIqbrTZ4+FlywADBeiW2E1bo5iJXD2
H0P0En/craqFNQHAPp1XRE6UCS+CP7xW80dmwDiCohdANqO0EEKjnPwhtMxKk9s/
ePT9fAkDPnJkIFuRxAdbxPSf8FNPeQAZNdJD2m3yP5cAGjLWyorpuzlvjbZ1zfll
FmaJvBVkqV9A2Y32wdhD13blh4IBdrg1xS/xVw6jAiRbAx7gpIWvEl+fyIUleQo4
n+09DAh1g9vKkGoMbrbHu4ATLfiFZYdKRR+SVEhzlHxbM53NyEsrGegdFGlurJBr
oZ2bLkubHWJeiVJWT2npmeK4TWeQ21UIoKgtU1P1haiSif3ys770rBOAohlB5uTx
IxXtWymW3M99hncovE2mXw5K7VHC4NGSXjLZ127pIyrmSOZQ/pwJM/B2VppTgNBP
KtKyArwuMmMWP7UaUkvMJKBqzkY+mavFwoR9kIiN5Uw7G81/FiWoNelekrRTdEBx
UPUZt9ICg8A5UcHCHJ3b1ADF+kVWx7g0UZfJMaqxcdm2rM/iUCRRm9F+dFJVH4iK
6h509Y3XtTwd5+7iOrVNCl/pPlZSzxmb3Mhkspv+l1JI37Yb8oEisDZoBNnsx8BG
8bG/ynAWsczHze2shgpd+H8VgDVUOmODJOjh9vM4YNy6wnWchlcf24I0HEc+Vo4F
pj5xhccBT3m5tsbg6hlR234OYOK6lrIyCKHDS1FVC9nHMweaEd01IPBmj+mmzd2u
wW1QUnN8W+cOkrkqPaY2EevMB1iOoOuSVNJsGDjhRtkRmoMayep+2BoEizrtxzEa
wwAI3Yw2pKIoed6dtCDWSQZN2JcGCIRo2X3ZUwWyGtT1skmMnFgi7Cf6NIdXPINH
Cfo6gjhhpbHqg+CYjzY4xgkzFus9ZphjWAzhWuY9Gbr9n4QtbglDesOorbZdJwoQ
HvHyhWQHUfNas+tAOUiXqZgIn4inkQMaI05txWHn6PGWN3577yllvuhfgxFwVdhD
XaMsycmkvP0M/0NApbvDA73UQQprO3FLB78ZQrwoxt7f3RpG2F1Ux7Iu/bOOXa5V
5VednYd0Wjadg6AzZ+9L9rsxCH99UJWVcqGR5vjSbDmp5V2WujRHAxPSikruVZDh
Z/JHu2hCC7CuNMqRBZequ0gCZ+xiDOMmMryLUfPrbaTCRS5019WP4IU59Jdt87qg
EBZOnXmG1UsoCed7m/G/PTkwFWRhUg63gQ3NExcCKmZy+0hviOH/11ZkXyerQ3i3
Cl3w8Bf01bR7bbSSRmkHG76ri/9o2HYEYQ8bIQw5EjsHsW2Vo9OOmFe5axUDJWdd
SMIZC0Y4Dru59SIYJqS1EO03Cf2ApX7TW5JEbU0dH7bEIgPsJS9eUZYrZ1UoPSeC
v5fPgWifygZdO3bw5k/IO41umwh/F+09bZ1hoQ7tH+luXG/CwX83GAyZdyTpNCdy
U7STeVe8HIKDaBxjgr91EdT4osv3cwxhiuN9wQvnsk90WpbUF9uKaI5NE46G0BUL
y4kVmmLNqurZsueReMi6tmlGQa30aQYkwO4sv0GeoPuIpkDBvkLL4Q3o86cQpIC9
8PgW4JwJntbW//IMr7cqcYN+pInc60WA/yaeeHKapoTPGuaQj5DF3kNj86qQZxB+
iFVZasFVBE1Puxjjc5ijeLMM2ah34oCkbeT1ptXDriwRWy6In3KxaOT5PQiDM1og
MMtBF0X/LLroQYbUjaLEfdAOiNJ3nM7MA7ynaLLDk4egKa2bumZeeMCXukfwcodg
Zx604rMvUtdE6v6Z/VGPDbyjO95m0Ahh9aA6myYCYnkk+cLv1eMnN9TjD9LzX7Q7
smdAG9EK4ytKm6a1IOmNulAg/+t9fNVkYQ1g1K1nuKqBJ4aV8CQucaWzxVFvGgFh
ACbJIw82JCvOW4ZWc+6lfBlJZQOBeo6afTirWdiTSepUXGFqsEEATX+i9p4dR3hw
7dyinLW/RyFingcfYhUR9/441ZLax5TzhqSYvITe+rCuvi2bc8w5eSX58gyzzamc
Y//0doJsziBHxjIaQixc2yMicXYudkfr2/d8mIGS0/6tQi4JsPyBP2nW+VQTORcN
SHD46XuejfIBkiZnJ0n2IIds4AKmMGDGTOcHwPRLf0RJwH0NNjpma//TtgceVFEX
2OAsfh1SzYBpCkoVbcvUEBxWF6mdD2pMUbwnZMTDzHrFkUvZbGSDvksAFCeKtIv3
JDLk55Xq0IqbXgmWjMo9DmUTdT4v3CdFI8uaPxiOe2j/CD6n1/y+hiv490Y39GhQ
BLyysEPrgg8JZsUrn2ruDGiTAUSXXGfLID3Xw9Ss4LYd9XWtPCCCBuRh5nSKutMp
pSq9OfnMEuMLqXY3bnMsJSRx+AkqZW4S6AVvF3T7SbFwg9wfGNS7fq21819j3iE9
WBLSWjTxMd7qjiL+gwtb6GFnws/Y2FE5BkJqcbd53sYUf0/Y7/al74laMILONB2Z
D8p4rSLUO9xMKC2rVREI+Dl+QgzXv6ut8NyW5E03Tuj7xU6sA4zSv6txCRNKTZBU
SYcjqp448zt4j3QptzV/HTWeRRy/IiEGqyBCbkHKs54YuYIpx5boha840kPRnqTe
1h2HOdsa4Nge+ikNl2P2nndwtV6oYi5lwbj9LVdXiqAwhlMjZ4B2BqSFR9ZqM+W4
K5WHuw/zKUEi0MMdgLBJuk7SFVAzTAJgpdxY39C915RJ7nUroxLnAgpvXjW5B3uz
J+lS4TKQf4kRblBF1ojXadqzs1VO+0KneX9BegV+QcMaGbtDC8q7exR7kfgua+lD
E8xDZlBaHD+sDzCeJCHjiSmsQdyVqW8ooMbs9lsA34BgR2y2kAj0BnYfRYHnX/Vc
yR0+zWAuLsUeW4+9i8tY0/XB65BoXFkkRR3530I/1I1x7UoBQaU3KJTCaF3aMocG
Xvr+Vbc8kH1e1l212FDs8Rt4LYhJanKHlLZO2guw1mMie9DKdMBWsU5fY/rqhLe8
TZWtfZeOTVzatxA+rRe0wM1qFz20dauvjZXrQzE58VZ7MmluDXJY+L1/T8zFtykq
p4eCz9Fy+vnzWPJkByhsrt0ctXf+sATjA2bbCVnbnKL5or8K8xa+Ei9mGL4rTQ0B
doHdp8QkZSARwwFoFEd+mC9GkC+nUn0SFbsm3RIgyUuwGYSsSWCsLEq8cBxh8GH5
L049v1U64vNyxSK+U7dZY1mHodPK4x8ToZE3B6dZVNxut8TBvzujNRKHyr+L6llJ
DgMPojkU4hsdn7ppohn7gG2SbeBsasC8js18yRwy8TMmyftB7hpPxJo3pdc21XS7
0UXYNQjbARhy23x+FSeP83ybCdH33kmnfiN+9XwcEORYxMXnZlpj963K+2GltHWR
eBKeRZxZnECgpJPHwXF5yRPWf+pAQYzblczI9GlLZCLVnRnk8at+fD9Rj4V9Qaiy
ZsTuRl9j98IGh0YLLQfQghvh0KqcJgRjTS7g9zDWbUCbzWdambywaZCf71i+78D+
nyBLZ648t3Qr5DJ6uBTpCfHWbmtuDubHZwrICFHk31Q4CY4fr3erVptfbqOqFPIf
2RO8oqaZ9ExJ52Bkcz4y8VCR+8Mr0F4RbS2hiUlGVCPtBqQRj6fb6VQgaLxTj6kX
SFRpIou4eVmSyA8TuXtcjIkMvsoe96iJ32CICnRdc1t0FblPwJgeWaGj+zOQyUBU
fShGmo2is967PJw64857YE7yTP5ppEt8JUK0YT8q4CXO8HaheSZ9rJBsmL7UR3ie
zls1pKU6OhwTFySup0zpl+E22tz9ybaZhEvwtEi8FQ6rt9xKLt3UO0Hp8+bTz+cn
/Ec7JaKqM+pqsRmZ2RbezVgQ0cANvuUcp588CIH1Zae/GmdCA98b3vC5nSlHHY97
Pt1ro1znhSHv1yOAbV2iY9oJDNN/ZV4tV84C7pex4sgYEmtWOR1PQgaZ8uOiJ2if
Or79y/1AWbFRWKk/byV1gACKmupucMSN1pcW2nAMOSEy8M5D/cVQ6yUM6Su/996i
Xhi2rvWVeuKu0fg01t/d39yUwJqJzvUwRgZiXvNgx2SuNWGGeGlCNvhGi1mrYeNs
KDItAV05yA5lvrI0cmQjgw4SFh+P5nOCbqlBfk/WsivBUQIcZsyQkzBujG8mZZDR
3gYxl5Y9FJJKVGnPMBYRheySLsRqzOqT6O0dTn0esPe9NJ+05pHXDuTbquCp7BVk
At4dXoRg5B7GatN4cigyIgHyC0wJlc0PSQ5pV5xFih/YvQ61XITNGoL8wodH7p3K
wT3GSBEA9uCSw03l54bQml78Y2Lv3HXq/0nMcHex4LP5tcvQ7t2PxBoRfcHd7Jns
CQipn4VtVotf+0UiDk1bAslUKqpPX2XUGm1cOL9pXHV4H8fOgfsFpx2516ToyvBj
gSegH/ouYfi3ZLmmFPCjO8yA2QFzL9/57quCGmc9meBDmsvCoCLXkdFc+L9JHu+o
Mz8yl1h6pcnFFtpyC4NdHTTWSPkaHg6MphEOFQrJaslreWdYmQNDUZX3ndDwXebc
dCEB3WRuyiae+jQYzQbGNxzQ4TQtcUWuvF/lzeuIVHFgLN/QzJRmTqjsuqt3wQwK
8G4NS+9clu2kUBlz8cNmN3a/hvGiMtR0eCKXzMTSy4coT9EfiQb2QLM/vx8DaqGl
6RzxwJjGVgsy+QraUrPX5CQLmQWKqMyb7GwCljMfJVfPL14bzAyn2VIBWDXroQ+0
rDdE9ZE0mPMSJkGJMMb8KDQcKUZpjkGR8pxO8VseYqVULhDTev10occhneqZIAG8
nCmFXKg1+153sB2A69GDM/FfHT1o11FZRfQDiii2tfqP8xAJ1rVEsm/tx/BjBLnz
NcmuVkwYvKpJSJ9ycel1iJWMdLxhdEOwoDUm2iikhZo3pusZGThljNQ0IJgi/Fod
VwgbnsJgGM0RRauwuWnwZazlIpgaH4leQclLcQ1DCz5dUp1Ku96wpTbHxRC5Y60J
QspNFMUGLk2JlMOBJAv7JozegtY9CMzyNZjeyJsqIbEvVoxU76Qt1tgjfh2X3bTr
qLXCBPPkjZ7FWrSs+b4ELHd7bQCWvUrHu1e3JVU3aWjTDKjCU5DkyUHxVSw+AZFy
9WneSLfHQgVpnzlXjn3zdlJS7ECodrT6OD5sW2zNxbvLbaNxXoQvcHvl3mQs4LN9
VZ/IAol0jrHwlLho33Ef1yHklUie7sC1qPG+BBjAlTJff/g/cELC2/2xN7pzLjpC
WEnrgOhxaDO+JA06LCKZYC+ucmwTNBLHxaY2/sybEJnwu6lo+1l6zXxynkIWCg1b
UhFJttTnCHT6Oe5IF33ZpBI09znC+znNQeZaQpzsTsFvC+VxnVavqvcN4lgRnMj9
Oiq/mk89/2xc7I9mTM33YCqZjqeGWjZtE2r1Rd7DzbkkLC/7HED8togVai3xngpE
9qbc5EVIYik4Z1LdNSsosy+GRjirfbnGH0iei+qlM703uAFw3aef+KQqKuBrTENm
5+IVtFEL5JPKEf/Q7dy3uDPVywBxv8OttB/VRgYHL7HO7vcoba4UTPif+Ax19VF/
/L76fX7ond76QKlUX7hP/xYdp+KOR23ISzEyBWVYrb2NMZNsTUlZx/Fs7iRZQDWI
2p7IEuEKWUFbAyDH1TOtU8MN8N+6A/bHeX/mKYdJrJk1oWsa3EnZi6qK9TgVFJLG
S/vEATV8YDa+bG9tBnxN1B6oUpC/HnDm2J4446aDWGIutgmnbg7zHqSfPvM1ukJ3
nKtzVUp6LojkDAOscn5YGNmz23rKh+gLYYkFANWmiL03Id/+H0gEaCJarnG714hj
yXny9ve9E09v4USFmlyvcVwM6gKRKFDqWpqZdfT5e6zJJEwzR7BGdcw6OVzvMuug
F2Yc8Njf0631UIAAvQCpHsiY2Orzytiz4PDfhiOaF4IYKSeKhXEfYKuHYShwJRbG
qt/XiZ/LyBptWKlcs85RKXeCC64o+mzJiyzxMiLVxXMtF2/nNcDD0/i7clI7DrxU
3w6cDj/jk1hvBdV13fRcNacf2aKY2SzLO+drVaVIEjDEtKCpqRdpsS5/3pT62F19
anSkij/EmQ0eRpWeCvbZ41be+wvNBFNGP5sAnHV9yJnM6adRtPL30nZj931hmOIW
P5a55PFM71v5UoYE64pqVdZW/wmZHXRpI7lM4vec9v42t2F44zpwbHkTF7GJ7jDx
pMg7+zK7y7Qg7BqduHKQ+Sh2kTZ1O62Q48McMcKIghbwWUOjdl9YzxY/5pLkQqkm
4Pmcwlsk87nAQonFNtHUsM6MnSTM93eFQga6CjUIrqOsWfP9K92vk422gY1Bh02Z
55MIVYbnZ+dOT/p21qB7CqXKFH4BhCzReg66gtHeiceOPLlGOf9Ycyb0FPNq8KX0
Okq8cMeMuW/V61uG2QmdaGH1E+b9OvpTNkW9kGdAyxFe0AfRkpW9aSY0EqeOAg1b
BW9pNi1SmoEcdaHN9o70MIkKaFVMdRQzcI9vKfDIJ18HD07aym0t5Nh6Y2qy5MG+
+DJzvCMfI8KGz7SyNNhW9Qwl8JWJ3cRtPDhH7p6ZeLnStx1OQZrlTiBrhj4xdCdA
l1WXMGcSfB8vpNrj8v5p0IzJIu1u6tDhsV9KwOgccF+ei5mKLwXPAkvmqtXKn4D9
cgj9IS7q4IB2291xPqJK1BPnjoCBW6XoPZ+uTsNR6vNoVIvtkmyhwFGpNcTqdNMH
hWyIz0e/shm8CG/y4rdxD6zCTR+ZEqHRLjHltPsK0ofIJNfkJgyoTHDC4XWdRQWP
bLnXlBT7NywDOwNf5GRUeWluLC+lpH1qq0uAAVKmZaFetdXdsefOmjmU2ei8JkUv
IVz83lxbM+gOEp1UK2clVGK6ZP99cLLO3hv0m199jfst53yQmNNA8uJS614bctQx
hw+qp/aq5WZ+qAhVJNY4mMdWe068vd1+RUrrYC4dXh+yaYFOO5Sg6aIm/UsxG62n
7rxEODnm/vTkUSEZtkErBYLVfOUjq+YzZ+YyMgovxl6zJ2tvi8XoHdIQK7e5LFM+
l//BCgIVQRhrp095YCRe32a+WXUFF1HvWTbfVKMGimQz8/F+BD9Xqp/0M+wXOQhB
6VsC8jWX6GGOqojnj+9X6aNk/VbcQt6/qj4Lo9YbHCLGoGXKvzZ7OSSPluAg5Sk9
B7kOmqqShlt9AzCW6GN07Jxv9YsvJU6gRFw+A586t9JiBr6UlD9mAVhlOuvqydXg
w8nwfRDvaEQFeB6XKbf0pn7Q3kuLVbFyXvBfu+yb/bmabVpdjQ7p+lk0uk3isyh4
6qWIKw9psu813VCxDKSx6Rau8FB5YMIGO855Ka/iR8JZt3WPLUZUjcOE4+H/iUk6
nV36j8DYunmvlAe7a+G5p5PN8hgyN11d9SYqgTv2IfVUCp0sgjZbXbLjuvQzA5A0
QuB5pNfYfV07CrIwKcy7yPbIUOj4c2lKA7DMQGVBy87ScH97uZr4SYB2u7mi8gGP
kDRLA/vOSeeCC9kOZdPS/shbsomI/BQLlU4EaIA68uqM7ShSQHPkN4UXmYPaSq+t
CZvDopK4driUvIx7s4yngwOAlZE97x54iJp7DZDvpr8tzh7joZrY4iWMZvExJA+u
+vNYM+QFJUnp3IY0DF4ORXgeXkohyfZiQBcWfsO40m+AEWGQLETcHGQkokwT1rR/
Mcqqio6Eyrv1W2PaXmPaXhrTPPzF5mW2W9GELQ1vAStov3vg5dvQSXgWuNOYynHO
unoORw5q5T7gHT7TRUJw5yL1jgy5A61Gs5UGW9Hx+iiD0zqXOYLVRtOvurVnyuf/
BhEZOAA5aXreWfvkIdOzbhRA04J9nyX5mbOCVtF17u0W4q/wndYQJug0yEwHXMKk
a2blP7bI3/m4iuljOQxSGKGh0vLeht28Zb20kkotYE+SsiUcR+x9yIG6Vg9K8fUO
261i6wf/VJ47I12ChtTUYzNWLXFrlpodgqA/4rWSnzPSONYE3x4atlVw9U3DyZdB
M26sCXvYjo//mQwlG96GhMs0hleXLjOhs8jzeVzaj0Q5QMYrC1s7TSarNOzSEzUt
D+HnobjVkhssa8hxmiK2R48libr4XCdTUyHa9OaQhjEAf85Mp9+3xdt7WJ4vHkl+
v2FeVJ7pzJO4BJp3zDl+jRoxBNndVpmPki3p0fELU2Djnpevu4SZbW1Y8MmW5JAh
dcc2J+kDeWpacScz44YRgepQNaTYuHq6u1DkpmytyLTKboR0FFVBRhkgldRtlbi7
ZaO+KD/9ENWVBODO/ojo0tRxFRiPdyyblXgj/+HSBab7tmylulFhnoVwzSU5LBL8
dLTazZkPSoPwmPRfG2EmW0YiyWUdRCHIZR4hKiwFXM73JxkzdXq7ekD+kHHSiAe/
lAIPd0EH2mvrPbkGqXfxnkXvT1CQRz8Ng96IoWOYpz/fTK3hckNvR4j7GrXGl6n8
cGIN/ixRzg5s3eFgxnk+ct9zP6C6PG3S/ZAiAgcCc6Q7xJTB1KvYaVbzEJI+9Wnr
a0zWr1v7afYQyCSulfXFp5KMDaDm58LHtqiLWre/oLtd4tc1K8vMGUfQ2ZMmX6rP
8DXTaAIotnzfdM7h27igm4ad0ZedGKCHvRDv1X2lzqrr5BDfCcBBA6Xh0F90OAV3
yYBYWujmo/tPhd3SpflUBRwc1m0fuVWFOr4ZhcwPLI/2J9bNGa4UzW24ft5qWvdh
5d59Uln0ZC3H1j2fZsoNKPeclQNI5+u3ouyx5XnlCbbIPkfXCtZPuwQbu8xc5VlD
YUknDCmdS/3AfgwHL2U5YnWNoPPDMeohyP6m+Ep2G4Nb5JVsnu4UZhrL77hkma7D
px/ffPUX+W9TST5vHOdjWPpm9LFX6o8kUblJoaluvtj/Gp+kWgnlyCRUa7hM8qEb
npv4FvAHLpB6r5mYn0c/d8MtCWaAiNSYBqPjyVg2pxKwLYUPL89Xvtjl0CzGP6JJ
0arCXoZLUzgGxZ6JtThdZyV2QoEXgqI9aikmUulKhMpq6YLjJToJvanbmPSytxf2
+v1+f/NNEl1xcGPm0eg9q9L5doOI3IsyTfvhc4HnIJTBg0N/nt7H+fSnhPW9ZXV5
K9IyDHUZSGzZlgHFC8Tl2gXmILUTj43YFtOcDgBYdjk1QrGsesWzgLWFYeIhKnnq
5ua7iA5Zv4byYasTKWIbweWctVCr0mTNhK5nIGwPcn45eUApe9894bRiNMbUAwyk
JEQhKj3JKIKQ6WsAuo2LuKLCSDFOmrVdShriafUua7HHz+O2trbTplH+lhWa2jHn
ProbAN/DqW6Lx2Ilx1M6VOrNx+t+j37pjRgFqBosjaniINiLOfWDeFBzovm8I+Kk
cmxo+KWp5EKKqsvaRZTMCMMPkFep3BbvlQhq707hUNNTrIkK+ln1u85XSxmLQ880
AhHlJbjRzuln5GJ999gQ3xKcDiFihZJHBiBF2ZVTBo57EK7MTdB7M9MLdYZDQVIJ
7L5b259nEzKOlmiO7Dtow/JfcWT1sGvgmWeaRK/nJXPz4CUqNtggHm6am1/+OGOf
UbkqgPUf3KI60g7iIboFoobjptT/cG0MBPO2+MXacpQN6hcLq4TidYAy/IXFEvJa
uansW5yU1633Rt6/uh4DiqjruuH4RebKlRRlUP17+KA2IUrFWS11PqWUBjb4LrNb
s1xaxu1wq0tYG2KuanrH35/GSEGWifgOc2NYZGvqmeExLDBCILlc8+16tawAxBBO
xT/ksXgIzGajO9ztk9bFWB0sYNKgpPParJwcxf7cXNAwJQzysD34+e47sjekrbC0
jG28U8o/QPaZ8+XLCze+5CQCSkWZUpMYPbpPLZZ7q2SaxC4nSMDTXkF+FkPRCu/c
M3QRH8/uNRcz2n2X8XXo5LJ1Jter3nB/2LDuwYfUpYKxippHMkTBhEukEStU3Nyj
og5AGZrDW9XnYxPD9vMVzHlU6evm8EEw+Dk0x1neYsbwWz+zVqUzDDN+WgBG1JCD
HfizikYkcn0Re6OkDzdQ7ehSDNpzEbbvl2a7wvj2lxqsx9/cvlChsAMPXiXKRlrt
eSpuqrKcBqMXwOkPdZ3W3NAUuUkkGizaFukLH1OGonEZGDDFHceCkV7xdUluBvrd
ay51/VahDiM7h4PseFybtVn1XQc3bgRtLvKNjsmqVrLzjZ2JMukI3/jBVmn98LVA
4Dr0y1ARYGdCmAmTL71cqVViedQ814DIA2zoJMi0y+jxpdmYcxGIlh1hZoKi78nj
d23aaZrG77APCu2uMPYqXNmIAL7SM9qpkzJUkYNkMBpVBo2+of4aPUBj5G0LcGhy
jyXtTVHcWvBDwNXXtOsNwxibGOtHoLDYrh+CVIouzKNX8BPyRm5uZL3Vo9spBmOu
vAJ2NQOyozwPYcPYCPtvQtjj0kZyUlbgD6eitsItFmYNV9jnVNR0vyk5sq/rCPRQ
YQMUanP/yoeCPkOr9HTZki8Uw6rWRSkfky+jsHcMlkAQhFQQMK5xzIkXo1rkPcVB
k8rgqu5LPja7F0SmbTqzWSlh+sJkf/K75iKVl+ytSAZzs0wJclbtHv8xd08QI9H4
OBvsm2CK0aUxhMZ3dJlkLI9cHIvgr42EM3pzBGIFCsPXhZMkgAqGLc62kythHHbT
Zu5BhEAJh+7mI0c4IUEvddWW3xWORD731wlEA2vNPELFMu3O/aTExyxoVSsN6piM
8VIBfD2eJhWE2Pj6w3WbfKbU1KIWynNHHTsx2tuDS1ZmSOZ6yyblGrSELNuJgaQx
J7sbhHsQ/fmuKw39KC4Wr/xDrj9oqTPIfiF4sandrWnXnvW9C5N5r/z2ZtSHYePJ
5kn25IaHGul2IXUWQ7y0Gi08szu8ZXCZuG+ezgAP1yjAXTThcmz5bg09OUv1+6KP
0DygadBR4WzAUK1OAeDWfNeHGq+zex6nwTa2fXeI3LGinGURbRbwf9eM6T14Rs4S
dy4gs8RBr+4ASp9dwzjoR24dGZLrzYcgb7R97315WsFQK5v1rjShLPf3Y7pXlfYs
PEfS4lCtnJWrAeE5Nu3JFMsDaaDXefheuwagO1qd+XntjtzK2pTOeaKmHChbxqHP
UDmWHpAb4YQelUaxWAtZxWBzTI35ny+j0/xh/yMAtJ6YHexNygKXlkUr4HAUN2ha
hsRHZL7D9sy4BGJHfgjCb1VFoEdnH4EFinQxh0q0v/s3ZJc5wCLUf2RDn6cW65KR
eE4CXtNOULg4s016c10pDtx2md2C5t5POh+sHYc7cjRBJOJMkUc6F8n7Y7oQrnWC
eOMm5/A00C+SW2a9IGFk/6PyQ7sa5Yr4J49bM7CinS0MiI43TvfLBiJrcJ5+Bx9g
NUA5temmg6FYj9GupQW5FjdcCSIGuIpkt+oo4Q8bMwskqQVKagxNDFpzq8ITWHNe
MyhnmTQRfVmf2thhuSGtgpTUTMlToc3iFhaItEQ5UcGo0WvcwT/VYmJgLyTa0dWq
bRcF/IpyNVoOUztGZeW70/0ae52MadVJeBOXsCXf2PLNx1sJHfpGL6k5crxIHULD
nLt3pOnYbEC2lD1aVdmhNuHutBOW3YuZv7uSPe4qk6kD3eh4CYgIMUzIZ4bW32Xj
l1nYfOxNyskZAquaNVpnsk6U/MWJTxL4SvQr0PTGMq+hrYgQ7m8yrDZBRnKoX0C0
P96388wSBRkvoL2HperUxzwjo1i7vO4X9MBOSG6NTtzNKjhVfB5FRWd4ymq+iVxK
R/LAkjAlkSJv1W8ZI1foHy8l5lQZC5sLNhZQ9vXXq8/UM98aUAnzCB+OjkAo9SiM
GrlcG8puGFDNhHdIIhscU/RnSwEvuhy449Lpb9NmbWAaMNuMD6rMl4ZqCS9BfxGp
Dd5iQ0OmOJwBwdGprSpYtTMdqAWAy/JqyOVyRMh6vrluvPXkYhcY6zSp/MQwLLre
NPhwghCAUA+NrAljvbMjh/mGU+Y7ZOsHDstbDTFKx7P40mCXzahlpIXVx0MHXKG2
zhsZPu8Mbui3NK7a/gJRcoKEBTO096VccamtqLg4CDuaGE9ZcG2OYOdvRQ/wH148
4BMF0W0vqAOVi1VQtSngeEG/lEhXJvlVnPwE3H/xcIugrgPkLCWohnm3hORUErx8
b66JCMW936LNw8jPpb9bmEQ0HoSUgskXMKfam+YKDb2TdgaTZquM+uynSmIgKa/2
qeB84Pl/F4EQCPeDU0ROQx+aQjVTPBOABO3fPHcwBFzmTbkbIu9C4vmRlTIwllO8
bUwncGC3TOhSnQ5oL0xnsAbrXiZfcxz8/AztvG+LZU58XFeC8JaLwPWpvwWYsMqJ
r8PTAdnS7GMDV+u8C8CPbPmBmZ1kccmgE9Bo4CSAOggf0Ihq1F0lqiDBOrJf3cxj
mgsGlelDyNUdbbRIR1EXgkW/fRrZhqv9bVDn2SdzvoPM0TdxsQtX7SBh6kxfvnMq
dYt8GrOIpNJBoEvxsdDdGFDRCeJ9z8I5zkTJZBRHwMFDodHZ/e4qTzt4RG7NRUNm
IcqLk9OanSjjzBqJHGGlicL2SaaSEVnXqpWWxhLUmFb4iUB2YI4oHXtCI3XDCpwr
eLlyY+QHYYECrxXrM/acKGrNG4tTYJ9/chtxFyYdYJTtqV+ztuj3O7o8sYoJQ4t0
RkDKnRBOdZrQy0FaboolAoxte1/yZr6QNfsY/ZU4bWtU2hN2yCnumN6Uj+OgqhVT
yZEmKwSaJbeVptFxcx4IITiOSb3z2ZJEkRo2poiPCwt+0xoIjT9GuVVxR3DLr9eX
bVgKAbbBq1A7FEVrJSoQYGowypg4rc3Qc2QimS968yf21VXi7jbQ5zsbIpr0rK8y
MbDLFwzRT7/g3vIEKY76BNApmOCpJsrdSeZ5EmpdXhknve5MlkCLcHuRZHHFWDQh
YTLSpv+aXUuEib+SunYKboV5yRBLF6kw7M0NWUu8EAHmXsDvUAatanCjV51FCTgB
1VQPcaFxVbfCZ/1JO2fcgkzf9BO0hbTUBNf9AhBBODmhbDGQ/3UKNYxa0TfdMKmh
w/sMkyGn2kDMfl9IBC2d3ZQla9C2cb6xiOHcPpsP7ZHHqXW4vHapAvi1/hZ64oqk
b5mQhrk+m68X2evR75Ho4tAlgHjbgcmJKGrkKOAfTEx9/2ezSK4c/GNKdfbdpABQ
ku+VPnbYvYvhsPpnzj2NFBNsMxe5UOuaRrwofSg0ah+TYr6BNFM12mIjIvBjUl2y
tmUPRh6mhn/2b/AFbIFGa+xzfU65mnoZbT0w/jFgbetU8qeSsjLOdSkiCyP89Fiy
PINOOFlbh2Iec0KmAfe8hKoQ8IWqp7ZvIYFHim5u+orDIKvtWa4T39PitbSwuXHu
hWT25YPHss6UYWTUPTVo8bFlOiY8E096VP1guDfpebIex9DrhTspn9TCu/uiBLHQ
lBpEwXynKkRhSC8YU5SaQrenQbickSpx+ZJSMj9IYOI/N7UJwOqTCrTnywrU301s
0BdSNrzAP3t6LvpDYURySxUF96WmGZnfPxFxWlKs9rj31DW6O4Qglu06UhAC5b6o
E2yM9RLWubF7tawFBCPPBebuier1xzfGoPU1KCB5q5nyGebd9gZJtDebukjVStHy
Xu5QeWk3YusY5NyVf5mNJXXRAtWnTULopPllpSw1aQxdaUpsAzgtNhUNLMrTsXOw
S1agWVvvShxQh+lth2BDe7pd21oD9iUI/CAe1ebLndp/Nk3QP3zgC430LVjGs+lC
nw3gyv463hdG9D3W3d+PjDA7w5lM5WFMxe64Daeoy0Y6zdFVrEeo3cCeF+i+xxyt
Av3qMuTyDmj2nLfOOZL27KHOe7r33q7IaJK3fox0Zmz2IwsCEngokewE7QGzm6hW
Zhx5mJBobr/XhF5jA/2KhKO8iz2quQCL2ACV4Ii7uGld/Il8GlDms1QLOQnSRtDs
RM9pJWNiqHJzfrIt+si8SsKdBzwtuc8vDNziS1pcM3vo6Jo0oafZTrSbnaCTullN
3RtZu9NFOe8nZzeHRXflLe8UxdjzgxJF1n2zYlMcw3wXerwByDaoxRHs/tcN+dRJ
l8HmP1qKODIQwFmzSQE6GUTEyxEe2mSgyBXHjCUBR8rg7Q9FGr4hkuaXR9npLkHS
py8lrZGnpkuQ7qKjPnVALEXVuTqaIz0IUSBhleXESLmEuzh1f+dc08yJAyhIDs20
cCK2X33w0iN7p/fPoSOS2uRSjkcce247FFiKV8bs45qNBszQRVHdjPOcdwxBkwHC
kZgpnAyrNVAq4Ujfy+d2MvkQsqNDfo8XxSUt7Npw1kW9EP+2f0wLjCKET4ZPedw3
n6VQqKa4vfUGjayIYyPRTHuMJcNE1JUHFRfV3NIMcugJArNK2ATbvpbWNTwGTqUI
FdoL5tAozeIoF4XfG/diXUq/tMLAebE3MLDqyRYObJa1sXVMbB27wIntMB6c6tRn
CGoZ3eHVkT17vXrlbRiwMZA3ktXSjbzwihBLFUiSwEPPZ8/uRXLEQYBVP5Vg9XEC
KJL3AuSPAlo+iRuFYvhjYGMpNnZ//pyYlb1jgQZs6p1nT1sZcHfAebjAXMkVnRj4
weiRwf56nYiIxEcinZEK9SnmULPDmPIiCv7ZOPCvztkmS6Tlf8hRIFj7bd9T7Rxf
mEhVgXzRavcJxtID+0znwhQ72GfpNjoaPxKwbv66riowHEBFuPbuUANfZu2zmVNa
EkGBCC0jE2BqoqrouhTHiVuXOWjgLTf3Mfs9LZzIFaMlvKVyqmuL/osBMQ8m7RH1
NaHAUln9x++226llP65MLzLtyfnER7clrnzbVQEx6dJYTh9eHdTeHtG0B8+JRooA
pntcUgGSOoXk4xHUCFwFTqz8d6HuNkkQqO3rKKsefDndZCO8SbQRwFBGhRcRdSKp
qLkgL2lIFzyPdId81rmfSntupehhunoYrq6LAKar6AoDXEgEZCTib1buMpX69cVT
JEqTP9kTKIGZO/gyI4G9+5g3HogeRhrFRKiA0f8x93pNyozv8Y7i0oidECqgCso2
6tacXIYdwtPs8W6MSUnEsOjZvdAXGaermmCZHuG2sz//odcdJjPkBZqgnAdumFcl
Ur88NAApOaj9QlXKaw1NoCX1ER1Ggorsjciq+73xCmAPM5IZiJRlSqcLh9zcaga4
cYP5W0Ca56lTbQeRBpXdBykbSaHKPlTxGSddLZ7DvIZSisIisjV6tEb48SUz93e0
nGu1Ttrp+H4k0s+vMODffdMttn2PA1D6cGJ94BWAfkVXrOCthlJ5Cq+GPlzCZdyE
cgI0A1yUEBhpuevXEVbipZuLv76qWwn69pZ3ws+wmuDzGGDEsPmYZpvV+V/a7hQd
ILoaZPc9+o66FC8hKEkoToQdjXdOvpyf41zU6Ixmu6z32WLbp0uviNZPlmJiUN0E
GVbd5SX2bcbOf1uY3/pAnWZ8apCy3yQfR935t9D6hjCwUTOrN1bD20fuo+9nOCrn
OJQUikEBwz43OvvXhBGjd4C+4UqC3bKSiumCAArDJyl2fBthjOW4Jnaw5HBxrfR7
Oy7yBPOi8hbhWDZPgBHVpPrFlMkL26DT05R2fRD9RrBQEpAbbdbmwuCX4JrNK3jx
ow7jhqsjo4TuTTRZllg/P02KjdQLLKkyCEvUDsMq3QWGWxBNbtp171XzL9kOH7ud
T1aOvjFeEIZWiHampTK3AAosONb1zQYqpa8n9qcP+b10/EVbOo4p1WGGDCg5R8bK
5/8qHygky4E21NaLzNtmppAJbX3qURpY4lcdLMKn5smysn9hYBG2bh0rSgb6JImp
cB42utoNeeqQ2goOuIZk+2bM3SlAN2eyJ9V+v0C9CgSeP+XqRRI5jScyWyGsPS+u
VyHl2iq5AtfaVn4S/wfZt7MtBuGUZSIta7PJlBjCZw6dpY53XrbXaPRQ3lshKawQ
r4koMSLI5EIQOaw5b5cfVnGzdxEkrd63w5Wasw23C+9CVLW2WBQsy/E/cFNL7BCF
NzF+vqEDJRWo9jTpzNRZ9AEPcHOgx0OBMUYGxIgQehhdvNZP8L1/C9HwIup4IMiM
18EZjLFFbJDg2gAifaNvFwtfDzzp9uTISfSEnecXaW5c8ZKu3D3Nk1+zJXXEp27T
32bnIIoa1BYgsAQXyB3vi4Pw3us/S4VE4kvh4m98I8bTxZ4JHb8ATSYnkSmx0PtY
KobFHpf4celAhOolwfQGeAd/RXAfOh84S6LcFI9hBd1fR0QWWvqvTC12J2+WE+je
DM3IOmphlSqerGGBfoXDQjtgCjL7DGbqa2BXecBAs1x3n5J5VMtTz3NdaoHd4lOp
P6iJafeFwUlWcBqSKHYmDHtsrIaG1OHcBJjyJ78Z2aBeVmHYA72q6ZPBMvek/5Wy
RYuLm48F3eERzOHClmjBLRnSfqcdK/IAu+xRiAz6TH1Fvp1mn1RI3D+Gz6RD4NmQ
UxkgTrqiAVFaTlzdM661FX1KkZCfSZx+y9Vg6bHlT410tY1R0mAYkfMblLT15m02
4xUSS93jbShxOWxKpq0/6goPrEddxJgVccBtq6dVLpEJY4By3VXtBc/cGe+5J2VC
jZoO84WqB/Q0Wqs1R4cI3MHt0R2ATtw2Tfyyc0o0DobPerqCg6Lox5qKUspfTyvF
nSmgkwK+BIkEFD+iKsn1NiP0tEDl7RleC3OLzEc7eRnVX68Jrv7GpEsquBM0ACqY
KSndNPDcJQpK06lh5jPk/OZ2SCuElzadWSU3xF+OhRgND4pV56JPcmK06cS/N/Cb
w7wVZe4TcCHHe2Q9wsb1f5g/z6OPivl1etBHpDeHkbe5tM/pxFIGF92llHnLGfa0
UDKtwkZ4xv3XJVXT0C1MlNzKMzvTiMmJ6aG65Q7LUzgqXxA8SUGlheIx1AyCWXQX
0Yq2nTi2Ez9W6Lli3UcOnGWPdR8nQZYdXLq/l75InwWfxalThLSejs1vedxWMU+y
IpXUatUkK5KugYoE58l2lcV8x660FSPY9FzoTR04dG5mGl7frf0NA85se/EZNzrr
05NwF/4mWFLuVu2zTHTkhkeXMM4kOFhmutDedThPBNFCDd3SsWUWkhEGhq/db4PR
OGMeB/1nTz5cdhzgtjGOcFFHSzFLDD+rIU4QkksocBY3ltNQcrtvRsYiaklCWp7i
pzTdGPwvoSkN8iXWq1HG3+SX54tdFU2cyLRlgHBF37B9XlZBLiSfeOfIY1IgPK+J
6f1UCPYt7VdOlAzsqIMbNmVBI0z3NG9pq6PzyOY6Ox6/ztQxTXBdhG8N6yroLUIj
TZVqXLJ54zpgiB1kli5NgWdoTGUgSLN/DDMEdRopDRV9bnKiNh89rNWDkyZdZJ+Q
yr8MVZ3zg574LSzPyaLlHUmrTI9RRVIMQ8fxCsbAUl5xNzewiJ+M2nWdR3rxhPJF
zuvBiyXHOJUTxUpBo0ZEGKKrUyE5UTz4k9A5l5zaUT+CuCtA6FIqldWEZTYeOPhu
yvG+8bFq6j0GNewDX13pxHB7XaNSYL7va61SnrjisI3tIRoilENkjp+i5DI+ghsy
RvhupNG0PAeMgvqOSEglNSBbBpXQcKXvemB2mbh+Bl4lRWpr1m1EI0hl9zT3xQnS
Ax3gm5010ziGw8B0j9OxbIKb3L949Dt775YOncG6uBbGcmFSzfHKyyf3RDkw+fkF
JUaihQ/HmtaImRI3p/0S0/hy6HImTSRqZ4qJHLFxebZAyMbF/hi3SA9o5e/Pz564
qHjnjh4QOos+HkbQFvGxqpM02m/d1ctfxujaaM+KX+UjOtigiuUItAIR/iTLDSPa
fF8RGokadhPhujWVpSjzloSQcQw3IKlYhXWutIYC4Al7rrNW1dSTCbP/OVNUDDyH
g2Egb8w65Ew0E95U5jPn00Y3oNJJl5dvQrgTmdxyyyyYI4yoWosvr0E3rBn+eqOP
EHOcLC8A167AFb4jA/Q/IRlgHA+/2ktallWNjUxgeTK50fyHfgYbmhTUVSuEeIVn
svL+H8U+Yq2WFmfRo1P02hH38qXa2J9OFNasTyDT+hVJBbaGxMZEWK8E6v8OJg5K
gnmo/0b27FVJx6+wwg+hrS26OOlT1dT+cnk/qZNbHNkZgGv2HteIFFCbXwykS9S3
KSu19QkYTJv8RjjxwJ+a1e+NPrXYIsh9R28HHteOg9IUXJjm6UwgOMTmZYt5cKIr
pCUlNEp7lwqEjnNpxc+r4ICy+eFl3DA6GGNpE+014GwvMjGfWu/x78SSte0ZDEaS
LXzNReL/d8cwk8jIpnRX9C0I4E1qg3+sjfkE1GyTwnMKGCwMlAqf+8yLwJ+AfBWu
nmrc2moCP7+jW+Msy4JhVoKlcD2acevqEH/oMZZ7PX7+EruAYmmot9ADbfil1sZ5
ac0GXGcM0GzPh45ekNWt2/o2Fpn8AchFvzga+K+2W6nw2z6GaIYYzw78tWM157nZ
6CZA4qAK6U2+r5mq5LohmTrkFrJ6WWESGnkeAUZoBRFRTaW5uTqWTNSCcYDrzjG8
/abSDG8vNBnpT6L1FgImwHz/KVB42MqHW9jc/+FZLXAZUP2nxvp5kAzpDazcxyhP
BSWdC85vYZZ2bK/ZXeqFd9GO+ebvBNQsb6uc25mMP0Ra2QN28Y8TmEn6CFt5Sp0X
41sjRkeBKm0+6lJyUlC6HDReDEZ3siWyajV98rNyaN4CbcRvB5Y6Tw5TiPZixwlb
IqizlXzxui00jDoMEQojK4nMcY/dcC29bmVbvYhczUrKxU+5PLK4hWYbxgRUjS7o
kjxspx+JaGfNYvCATuGR6jjjb1Xddzeqko5XmtnqIRTZJBfvbYBoxfE3Tks4roYe
APUEoC2lr3tbXbUHve8auiIr6/QINBV8BkjcE7oRiLL/3EzmU/J+xXv0Akh+Pk3e
AUSSNwTgASD0yrCI/1bpV5gU2wS6b59VGQERygEXaAtD+ttXOA+ZM91JhQDUn+eW
k+4AVwNkwwG5duJSXTPGQK1DGSXlGldEVKIzzNZi5FiCaooS9UTdeuJcRZWWdLUh
BFH/8339MSDAlmBm9Tn8lB9aeFsdrVMhDRDPD68098mIfmv2JhLmOOSRY3/e5370
hCjgozIkJX3KZ3RaEN3oFGkU6h0YANWsbrcNugAYBW2f7MzGb2LHxTuA4kNKlEFj
URozY5ozuh4OSpxH8WaWUVXhV8iA4Bf4HGC6Ec4i04v8WAdJY8ayyM8UmeC2I1qX
ApEbc1UxZUpfB6DKSArjipfFJ752RqlyPHbO9O50fAfipRkMCCGNyCq1J1M1yjDQ
q0nh858AsZ5iK5aFutK/1OFMIpiGFgezCO2bjDRnNXNPZjULvsxceR+Mee6OjijD
rPxGVLo/K+9JO9otEVK/YCM9fQSlyENh7QSMMXhdZyZbeWuSmUrf8Ll/dT6ph/An
I3gjuFP0Fhssi1hALk2avuNhcvgK2UFRG8WtFyHS/KKKXZf2H0Ht2yK5P3kZoTGc
PhnWUrN4SL/8BhCkSPsFoCc64IikcwRfUpVdfy3jxGJ+PY7JGMbEWnWOPg3Wwfmy
ZuWdujTRogqezfq1csojb3A+1ZzxA7/ztnFUWvBHY99toVGYrd5chCdpPmZgD9W1
mFHVnREXXU6XlZ/tRAQca1XUuggfLy79xSn7slUgtBb6R1apZcpsBZhWAg8tFIka
UiUmB4KolQm4qCExfUnW+5o5UXljagugiqeMS4i5r/H3eQLviBowhuRFzwBJRwlL
qM5P9LOgxJ/jgaIuB8HmhH0BS9jBJRLFueY3K3PmNS+UCw6ZeFsDWxSYtu5z1j71
yH0Mbv8olTbg5FptfK6XHzwxW+Z0zoB9+UApwsmFm+wNcJYpC3gyRrpXt/8nFVPK
ZK1OeiAn1rFIv7gtMfMyCQMsda+qE6IyJ64KkLU7scrk9DVPsqQ0YCxxbv3UemGg
7Tznis2Wt6maf1yTVHfWnQqbTDjD9yMyoqNxLlpCP+sEXYz4RJx7Ck9uKT0vOBfs
7uOuGYrbAlKPU73VuYioVgCZsviQj/OzTN8ubtVwdr0HNK+hbGl7rzflEKYIdJeY
zk5niOJ/7CqmF1uKegx+8ehyMWA9ZsDpYGWZazMAvqHQfuFZh/nD2FKVeXg+ecUk
WMST892cOYyf1ImlJRjBMdmke7bf989zsskZEcveDEWooKcCMOeMWmr/Ij6wKoc2
eIi0Krogm107ZKIkNpTgSnOJ2/dIIi+Hx8ksjD0jk21z2K40gHp48S4RIt7Yoqw/
KaLDYlmbOMqZ19oJyWSfnzJ+Ub7g3fQCF7zTXkf5QDiDUgdHsxBRnZvMjV4JnNe/
fUSJrBp/t2qNMzzzGt8OOFjlk5IqekFE5imtYiIY4Yeo+4bwuJR5di2JrrE9MrOy
DjvgPGBieC9pwozIt2eCfA9RKNEyv++i9I65qfACg3owKx49qnAqhA0gF3BisNWi
kpXO58ZRHX/lO9PXV3t4biMqpXG2oAaZcedrHUtmWvWgc5snyFwRxcZMig+L/4it
+t0UKRpkOWfqlj5xprxKBelykkv1+w0prqP8MOaB6ejVzoSPgGU0Ppmq5OGWc3QD
ZOKsfyfI/I31o3tnfguDTuhB734f3TJipXl75kJ+FAEf40hkIHVPXNdh4FfcT6zd
/6znrC6ncmFCt+UHaszOaKtRFZrUPNwxU76le4eIrszLz4va8+3ZrFkejiwgSoZ3
0zuU/YxQoC287tOIqVfYOqImxfdgkXBevtgk6qNnh78MTBZxXwQrgdwF8JukNcok
zDDSr0XfGexPdGhM3Mi7e7RoKkuq5MkxbJ7+t/Jb8TGu0Va18cWAUIGixAQ7ig6w
zaz2HJ3jorsJAVZNaIClF95K/3LKvj0EghQ7KMiX7CIss4xfJ/9iT3RCgGGkDLty
ds0lm/NGLDbTZAQundKTB/9MUmPLaes35h5LtAHRDFl9mYOCsRJutXbdx4Bj9QQa
5n0O+6EQJV7FfRp20wgIR1bk5zA7lCZlJ0c/nfFj+X4Vl/12vOLh5Fl5lxrhwziI
2dCUSI+ZKkYKnAbmEavlMhJ5l0NJyz96PGdjWAhynqt/cbhGRpYvQEnr9e0soKg7
u1I52vJ5tZWnB562RLW24MjGgcHGMdPGvvhj5Ikig7WmA6FlTn2Fhemk7R2vlGHO
WWld0ZfUCWUX6hF7XD10ipK4+IhzAuGSzM2zYbHZbTjzCiWZ2Qdo7xyoN4e7Rt/e
4h+2F3l7LGX4Ca13oOY9dvy3Cdmj4DNxt740hyxwQT3WdMhP7nFSxXLFpoEDuAa9
FWkucl07PzT/6P1oCNU6YNwWkvmHvp0fLR/jZLDGvk35YAE1w5H6Q21GiWlrO5H5
K7l/hHU6RWqzrejYv6wxYn0Pji69otbFQIv8lW8cIv7kzAZG1aOOzN4tae0kWczS
NMCZq6bOWTy5m6DA0bR7U5RvgdHCDkXHR4cn7Wq2tMnYyGWOYvptIFp8bz6EtMAm
s4wnI3i9WUYnfPUXhJSbXnc+n1Kn5z7vAkQ4QMv7IZjwgusmIhIJslDZPk29RrUV
ej1Duvrfbac5IiAmoY3QDw3xeFKFO39pG3/mZDsrlZxPiSauUKAkHoXGONke6S5I
w+1eYWR5aosN/Idt2ntGDFSbsQaro2X1+yocrrGLZ3rw1p//bVpqu8G765rCX4Xg
4WkjHabXS0ncgWOSiqedJWvrAYyAQ30r1cjVyztPFOQuR8fzJ/mDzJvqgjlCToLJ
neNaBBJwzcjR7znLlFdy5RNl0y4CxsYSjvDdN1pASIKkVLVl2U6MPfr2jlJgxgTk
rpPPYRkg8dL1cjTlbNMw859aQ1u69Ds5ZCu+YAw1bSroOfdHpsIprddms1c+9tRG
ZZ8z+pzUMrvKaImVIh7oAAFrs0ik0Dq0U8yKWFA6nnb1Ohf5KQCttnGYZfD/jbat
1053ha3K29ktODAccTmIfOmVPdY9qvoCbYHuV9ZB1htTCOXf2m0pc+TRncrbjEDH
750PjxPFUALMcDtotdIDdpnaP3+RPXa5LyNRIFoGl3cUU/e6YGmpZBK6hf6lwgBR
qU9UWy2Bwj3/PuI8dGSmhs4T1+Nn7zSrkFOLyfhCZ05FQJF3KOxStXWYvXgH7aFm
tpao57Z9xHFb7HJfFVSHP5uXLNuBwpSi/STzLyqvlcdpaVZ0np6VsGszYqgboc7x
cJEVAdT+EX7Ri9JWfNW1l2Fum6Jzbvs/a2OkIDSjiLYRxbFcHBnT2rXDGM+xk90a
kHtIDfYSjqQmEWQ3DQwOolXqU9cpwdQo7U0Q6BM5ppF1BwGWMJgDMkGqII8Z1DEJ
5Zlfcg3HDXqa/89WYpq4sOwnBRbJFm2kE23Xn/yOzDKmGe9qihoXmG1xIxZ/B73z
arOR3YZpqGWeuHdauJLFdEFgjb2pVBLuSEbgX6Dpz9bbRATztaBv6Zz2qdcoPzwv
8q0zDiEX7NT66Sb8ab+q7qLkTUpZhRjeDVL+9pqUU9C+BH+F8Tg9BCn/1h8yFPZ1
Nc2/PduH054Weo2xtRZGMasgCA9+9hVvcxudJrdpOhUiusk5yrR4CGDttocsS9v0
Ucdey0uSn1QL3/wMX4rmPs7FcGYgIygTbXRkqG7BKHy7VvSDdKND2AnE3dmskibU
mJntq4pn2kIPEK/9DtXEDVkl7GhpAMPUDUHsp/BSb+uUV+Qwa8MloUDk+iSsp+Kf
P4kpa44HecAzcuE4wCnvgOHwPom3WXitYkkmXWuq5KF2l/0Knp2WeTtn3CShU0KW
kORkGmOvbCf1mKHenzsJb5AEe7xfD45yf93fkFDnahXeBlI8cP1dgfAB/+ZHFN7T
tbuWJ1YYcA2+t+zP3Gz6PaxkG2ArMJTW2Lt0VzbqIMMcHXg8P83yVhlKZBIS1TXx
JwlJddaoOrlr7Be4uvsZyvra4fQ4HQgSbo1lA5gfR48YSJwa94qkLxxNC4D8AC2X
sCPrqwxJXEcP1d28vIKCfbiQ92YqJT8w9P4ABj/sOJsacuyaRMN5PyvpPP9n6Cgv
aCtWmTjkn8+e+QVS+BYsQ2Smr6XqWGxWefyEExdrZybfIG1FAX9Zk3+45DI+YTia
jo877w1m9pZoqHwjN55ljqNnLonUcDPvwuMOYVv2CaoNZ/y762BXcBuNOdMvE7JX
FDOS9PrhZSd43RzuZxszvrrCuS7QDjlMkwtoxlNWrsaI5n+tkA5XbOGFv/RVF9Q4
gYdr9rXBjxVDMuPeOvV2zHEICdf86P+wRb+dXyEg7oM0mYPdhSWgeLFLpYyCInsj
ywIQnJ/VMYD4W5k7r/YFwKxgpBo0d4fdrjEQ0EPK3JYDfxe1pYp7/hRI/Th166Is
CjTb7jPeCtDP1N5BwScUAwMeF0MX1lnaL1D659G/NK5+CzjKgHRn8XqFM5jCgWSl
rt56oBl/2jGNUDCYX2WtBEN3sQCS43s8divq36VOXo++ge3o5mjJu5rRCi4kUE38
FzzTfEBZWSCUlLAoGRPmYWnbYaVUcDklq6zq6TxtaEBhHOp9aLkl8iKE180lwpev
dEP8U2kxaZAfb25ZQa9MhTcV+NMMnaNaSXr6NqptWrJ/+rf/68QDZq47HtCiwVm8
0gcFymWMC96YqFEM2Ci8I0xPk3SonZTmx6ucGWi5zLmKzmlZ0+QRmwfIQEap6iah
nKgvSScI+IwT3b9/SftVWhXmF+AEL9BWW80C6hC/IJxv5CH1S3Qbmcx+6wivhP1Z
joaNsiMbqFFHXcJVWsQxByvpmHmQLEcqIBuolxqhTjDs3TJNRXnZ5kPBhW7n4fuP
mO6IXngQQFenyXJZOWyoWjK7J6S0Kyjx0yqASsXWm502wbdjchUTmeiFFPrWvUXO
lReUmR8Sp74FzcNIDzoCP6fn01QQLoB+7n56xXIyN+d441+2027xU16yE/TxQOJ2
anJtHbgKXlVxd6FgpSg8o+0kaAncO8k+kIVc/gcUBUNdOt5FOO4u0IsAeW3jr2r1
v3uSyM53Fuj9DZv8EhxdI3f5FG3uc5D9pu4stIGwTDg489DYYua1d36+/vDXfIKK
1X2iAgvzYQbgSBG/hYwzi3IQP5T7AZPK+tdAd0bcWabXpBNAQYcM+zeF+wwMq7ub
QAUFfvya+Ond1oJBg0+fDuWKFpoUpAl8hJmxcqH1o6hGzbjUwrrr3iYruEOwBS4m
lrFg3AX6Ww/58+NW7VsumqHjmZO0wgEHiEm/ed0hq101OtqsKTgIP46vEzvWxEwk
sATMHvN0GspSQxl7i+NDUJjFx+yiBYds2JDD3dbqJ/i0Vb2LSjIcajEGPNtnIGeE
ncC16cG9ZaEItpFHpWb4pCEGO4JidmTy2/30Ynn2GKEmwgs/8+fQFTJWilmXPyHk
5hx7pxWhRIdr2KnCVhTzWIsRPSIBYO7IDB5Q5VzFu6ywGLfKmEu0PE84rFok538y
iR/TRXQvAy7dHecGguG417h4D+3EJ1a9fHeftUQE0mfNJvUUhjz3CgfJQJw1msfq
EjpWRiOVitw95GU9OZWOTfSAXT8XKxY5UffUt9PWb3pn0toewAu5gbwQ6bz8sgMq
i5zk6m6FCcbYYzdbWDK163IifbpAw2et9cEZ9/nNEUGWudn2ZzkhXNQ6lmwUzih6
rzkEq1mxpI/vp6G1yQVkmpMjP8gte4TToxoCSDfeT57UGKKVKGeo7SUuxU9lScD7
QKu6kJPTJsECP9k1FJAKEiwmYv/i90Hg58WHNp/MzReB/iaA3iW+ooSotxq7FnpF
7s2Uc29dYUptViwDDdwk+PGD97jWpJuXgvHvQLk6hnSxVTmsc3Oo2cnD8mhhUPDH
jwb89FF/rVTIkuxuyZRQBuLx+iq4QrTN4XzWq3XleTI2udodzjhiN9SixJ5IlNPP
/RBAGvR86roEV5vNNTGpLZTcG8al+NesknvVPWzBixlr7cvutqgBaXrpjhxTzHtj
2tXMGbDMCTo+b1D09Sdicre7o4arYSlxXS2WEwnfI4BkroRmilCiUTnhO+ymlKWQ
v+W4w7vs+kTrISF8uh4NlfieDFe1blLzTKOgbAq1cubH1xqisgayzyoOWQpF8YRW
qJbubQwtrk59iXDGxKvK3zm8GNgrDhB9qeB/5AK/zqK+xg3bFBoN/86luzwswQzH
Dy9rFF7+EIGfhK42RPjK0UEq3M0SRNhw2N9kiss08vXS5fEh3rsi4kcMM0ntGuXo
oZV8o95PU3v9Qb0bIWyjX0zjcwyiIUT19lqyQSoFvZY49wPV56HD+vVN6FNwSus6
mt0WJVEC/Zb5FwhiC2glpCLKllXS7oxlDsoBjfvOd3Iv9zh4bzqxD/IIaD4GnV+m
HGaanwtrRhzKBMpCqS0iStRknoa6YauESCV8jHeKdDmB2ddqxfdg24CPGg8PpyFy
D4LJfMprtv8zh8ftoTh8/A7xuQH3mcn/JR49A1hiIR4HJ8tn79k1LDWLoQMRH6Ap
9FleZa0dkKsrkF4U6yKSZjOen8L/9k8xbbNhDNmcKff/iza2mu+s2tkZ5SXzIlvY
0ej43jKPNAppZu//8IotU16byB6OTDFhtlwKkd4XSeCyqpPhSIpDCfVrelrgSn7+
nvCv8Bosh6iplL4tQkvujHmcVdYGTKOs3BOBCXHU4XlNpoAdkqcCTiD6UOjjA2xq
oo1qTy/v7uZNpPlG086Qx1fV6tcwPX6MqGvxLxlC7bCFzm2T4Xe+S/q/XboE9V3y
BxyB3FTCQqY3SEIoOt9eYN0cXPvE3+aQwJV+VCLwz111HPsZ203YinqAXHRBVlem
2n8Z2Mlp9K1c+QEiQqB7GXXqokFdjCdWdc3UcuEt0Cey8a5nScj9GQjlV+0kEwlq
a7idpjm5oirhTcE3eqQLUMHrmYlPVbB9tLQAqLG6PX4Kpd3w7opk6o8w3YvS84N9
s2yARo6+bKNMllahlrOVzAGXLNarwYG7PGqTTMfgj5GqjUVlwosn3r/Q4EXWZj6T
iAKiayxpsKG70go+bTAMWeB1W9sZTdCT9A4rak0mQ6gJdmSMbTMcMnk4D3Me6zFM
+jPNuXc9Nd5YAANskn1o21ws2Txzxj+nZlcIWPR5nb0x3Jh6mBTluPrZM+DFQjVT
lAzUgo41nsMzchH762yjuMO9W5L6I5YQ7uxyWQY8UWJwXALV3A0olEknVUNEaPoX
eLzPKLQOgicm+kkGKlLuNytqFyb8jK5MCpOJKhsLRvVj3anMUGiGU9SAM74PA6CN
hDZdCPdmBTEIK+l1TQ3AUTPfesUt7R44qkyrWVhWNrXyQn7ASpJdm5IQ7qm/KtVg
nSs0ch7hCka3Pd+mLUNuWmSMmful2n6j+erEHHkF7a2yivaOVwn9cjVN3VdlaEYU
iHPdOA7Dg0YJcz04Fa+faN3mMT0oc5SL2qwFQ4J2KdBmsZXkRbafWcyyc5mIES0q
wzgDGr52EH63xEngZnKH7ULKAOOdiyKi9xyboQd9wkxoFhZSQDKV+kLr8Iu/xvG0
5LzJa1JQRN5gKL/+tWlGM6oxw5FYhs+zFrh9egKBL83IUKXaZxrQIQlZrzWHV6FQ
Dt9QQTUorP8IxOIpMc7uOYFtNbcOrv07+aopq9IE27+3ynsDZXNI0UPbUvrFKzDN
zkaxWKou4c15GoXuEokoXwkv5lryw37jqaHdDIGDhAdxr+ANGRSaxP1n0s3E+/oM
wn73Q6jBgg+c/rTwkbKkfKcCcPlD4BEhk01LrbyU4dkx9U3Taj7FqxNz/Jg5vYPM
PdKNHF03NSrltvCMV8SoRFbUCtJhFLhF45SfL2loGv2r0SUqiUEo0/xmeUkGH5P0
SDSUZZs/CYPzlk8rqUyAMvBLmsTs1mXvn+/Dew9ZsoJAOE75Mck5RAtrhoWzxd2M
gHCzKyGdqHc23BjhOZI2kmsAb7QfLibG9fsff/pxj3ggs0xJOJctq7IuIVoySAks
JSrIzLj9hW6UKmvJFSRYh1CD8IpFUGjD4iwrOAykm4+IptwpmZRAs63OxtG/8ojU
G1PAcGXH2j/w7z3vR7gTi8ARDKA2Hai+Gzxb8PrxOAO5LRllnKlr6ggPpOYaJhJI
WrkBXxmzWHScUgeuBHz4n3mrO+5bLJB0znfQMGCw4a07PPpalcz8dOkN5XuEj+iw
QiZaD/IXjsPj5IbrJby8EpLcP60MUWrdnSNYatqips3DEhQPdIxEDwidv7xna7eV
KhSJ3EVpPnUSmq7zMsdeNziLeDF4Q9bVR5BzPJ122M8dI9H/Hk021SNRs7FtUZKi
YSrpz8QvCYBJlzfnJmWYt39EcMrYNUYbGD12LlPhsz3fvzxilIyAFtwgEQbhQk4Z
74u00zfrb69Kj0fmz/XIy5Cy/wR2ybxgcArZVICq4keUQbebMvOISypkMAsDZurs
Vyl3g9gu0QM9UBBpkWM+wwDOwqnGTQQrx8B9+LfndsBi1/Oin6jqak2XTc+iGrfb
UiDU29OU55R8C89k9aIBJGWpKyE1sTD3kF7raXnB8fPfrz2XX1E106O0OSo7yqr8
Fhsq8nR56EQ/fxfkTgNXXduZCLr8faM62wfO55OW6ZhrBtmH4ZtgMpKHKXeGfWzh
H4wbXrKNaN+uWyKIuTHs75dJbcNlqNbL8rHVSD8H8S3cUpYPIQ4OgDzoL6IPyraa
eEZ7uZiZUuBfPAjkFvB2Z1UZ65Y7G9HXyR5D6zlQFnS9Ksfv8IM/ZoxnjrCZI24t
1Lemlbj79KFwfiaNBu0yAR19TcbE67nXZXuSqKkJYbaCUEaPaf86k01sEZouUc+p
PUnXvJzJqwiAJkdETWHVJ9r1bwYmJbQwefvxmSGM9NX5CawmkeTs9FxlO3ICzE5m
yXQ5W1EZrEL+khnz/rRXH15fMd6L3yUbbaqVd5XGB+7jIumwpliwIXcquZKcJ2xe
Xc+YQ1I3OWquMVWWY9Oee91ajPNyj2U+gcafCmLv4AgkpJsWrDVJJ8f3s8RX+PyK
MjXghK/gmN9n+/yGCKzv/6jnR1YutN/eZKt9nIvbmv61LZRU7R+MBkTM6RaqSfSD
xpK1d+HsiqsIzu7bh64eXCDA+3qxewQb7gD7blV0iFAqa63vuoilK+vXbJf8Rqrt
6jngbZKjNDZDnNVrti++GgEDR1rV2TGsY+NVe2N+jLb3iUarK8Y/DL01lJ0wxkDo
bjxsVjWuj4J6Lcry5T+Q61kwbOhFBMdaKwKa6x7yJWFXbKRK17D+VTnH8UKYhnk6
fJ0Pq2Y2mxO6DzYPztoRjsioZDQZTvJONlkFioWUlPPAhFyXdzr3RoPuSvMRw2lo
a1eFvU98PlmfmvM4EikUWLTA7U/KA41+DF3Toc+o4GfwKMeBo8HrmUT5nbuItf3d
nNaj1UtSpxgbHbC/4zM590gAgXOiQ8WLURMzJ/f+m4tSFZmxJk2NO1XvUKDHoRMU
+OZl3iXwvYL2qVI9PkrTJMEtCRbO3D5g4j9Z1DHxBWb85Amoq1mRHEWx1Dmbm82C
+/5fF3++4b1ZL/4MLMYgQMa7aFgnVsw0vku01/65x1VmT2sjIVJRCVw4VQQoVpvd
L/vka0iSoq5zVsvFKnMm/Tnva1Hsk6slG6+Ixw+nFTO30lSrOBWe4hcskSHml6PT
6RnNNEEiTGufEukhj/zoI7DVqKQcW8R7QF/YG4qUsOrZj0aRjB08uoYrU/ACfUJB
6SF/CFsNJC55GD4eZxu+u9teOk9nLZWIvvJ/chzPihnyeRBqLwCjLw4y9vxZvnK5
YP1reUukrh4HejKgnatf3swMpDtVrEh90t/oBmXmXaCuGhMb6CFPzL2556fklLCq
TcH+hI5Qm+Dmm956tAsr8PNVCCK12IftlDHogrOtZw75BqFW3aGit5ItdKRuXMvp
QMP9PLQzPUBUYxMCD4g9vcYXOnGCQWY3/B0KfKS+zaA90Ww7XSruU1jlAlc9gEsR
Uv/yj+4hTtwO4XKGsTGTjDCNDfeEHjL1xUkPcupKm6ILAae0k+I//HJ7uJsWo7dM
QQ6jJzgZolRneO4rOOjOmTgElGbONXEWTITPF3Av2/eNfcevavE+cG/nAmiOD6vh
sz5Adhm49n/VudoUZzpcZU+WgUTh73EtB/UlNRF3vRMucxxkI29igYPiviKEON65
UkfgF14k62HPJVaIxru0Lj9pEVp3jSv0Z5i5tXo3nvHA2q3gY/tz/vj0x8e1SWH1
rfAgskxH73Bgqz+jeNv5ryyrGyGPyUyslGDj6mmv8OOzhzPl5eE2lzvDfu1bI6ae
ysr4AQY794NpbKv7SZAOIq7nmMxw1F2/OqiJiekenR19pPGfXwDkK94PMBsoUzBe
21oJJDshMWnvrVMt+pEruFd8xGY7Ex+tyFFHGsMr3XFLd6oO7bUvyHa9jzt1m+PA
qy/7tARlEfyd6Q2uORHJ0c+fZindrL+VJBtMuN7uLQTDdpXBaHMWi35PnksUIis1
2PqkbOqxWeSOQego3XfwWND7YvBBk+WG6g79mY0sr8ZDFZ6WE4AJmPWX1wkD0vOK
nZUqabFycwOtWvIblssPLSs7J394r0ZKhrpHApWYZSe+4cUoUQebQA1QvYxLL4Mx
99wmYYzriuHpNIdN4hyESA4NLHL3z0szNzU7aHzlnvsd2ufR0HUUSMNk625gCVra
XvDJrQs09v8okipBbD9EYH3YK80v7OgKxkJZxjEmjAOxEj6E87J5rwwRW9+Q4e+V
4SJ3NGAZiCoWOmUjdv/NjhPHXq9qO3F1Es0jxFCdn8hNS++ojbrlSDjqqHXsMSrf
ONaExNu9lP3OCA89CJ1uzS9bIU99vCEOhi1HUh6c03cNIRaBYrpDNcidWMfkHvci
wdO1IvC0XGWFI3D+/hi26di+wbJee3CBSlJUsZiBr/u3bcp9rwMYNZnS3IeapCzx
jXAUBN7qArbeEvfwybpvapk+S+9L46v1GbBlIc5DDDlDoZKdKpn5eylaaNe3aT5v
U9jyj2481T01AQeu2SlgwNlePpiTAKOpNO6Fi1NNREKXT06ewdgtk3Zo66RXyRmH
+Pz4RfM06G0FMSyWFTrHe7pko6Vx/lwu/K3BTtmycwsrFsxS8IvYjA5mogiVQHCX
Tz9KUzPw3KlW0k8D1V/joYsCorl7AVaQUY0Qnm+8J/ejjYMo257WVToRbswWaFzv
ha1ps769lKoGFuWHrj02CgOfYTklmdVoQbndsGIcaoM3SnfRiDY/iK9uNk1fSZzI
RmuNQlYXcFtN8Zq3Ir0S0DzWKRmKe8bRi8f/uQCnEL7NNZiuZ3WMu7vHvkikmrwI
D5IxYIZx2CMo1Zg+NSCC2kBwyDpVo1KbdG13b/U3VBoaeS1n9whax0gelz79wXL0
ZL9gvfSEHeciRja6rFGo4ayFKBh8kRkuDiO0EAr+4y9oqh5pTRBgV85s//UyW5Ry
pxnEj97qnXpc+Nkl3x7FtRRZQIp9zDOBabJrwiQLjDeMzQQCGkcQOAGWYQYUW60v
uEsTgEGQ6GEArqse5qwNsfzPQ6RvK0uUSpsmYskCJCdZXtQ3rDZuYv7R0BWdSC1z
wLntHn5s1R6Sogw5ioqwV580pNMtsefrQcPGMJUEvH49tIOlStBmUbQYvlzPFdIu
BmMpOJuIDx+NfOTRn06ZC+KlgVVD8dRhkafs462OSPn+OoMd6ZRaaQxOvkD/LZAT
hPB3/VYhbxgTfhj/0gJbPlaQGsCER1EkPyqMQKNuPV1oTutsYq55JxMRVjuJ1TfI
ECvu37kE7FcfQ6uwAzaQUtceqEJGmcv5m25PbMDJcCEY4gtQi4LHCMgcILxKxQD9
YONHlKMk7yLmZNkCvvbTpd2Bl+NWd6zIZ25jfZBJfIqqwayPjFWkoBOICufDT3k8
rla1kW2k1Fh53UlBCj64FQV82tuMK3fPLAZswkGNliInmMVc3j8gb0aJLMrNp4qO
obQ4OnvgFAJ6LiBCmSxJJX3aR6hUkyeWhtohClLlsIJNVG11F1OVds2bdnWIWZjf
Qcobi/tj9PL9tUuosYGvpT+6Y5DrHwXj+3ylTv0/StKEuarKZeLWeVISilnD9CDy
kFkaDT8tGcW+yxO6iETN8tmpQJZnXDWArXiOHNs+vB/DlJCDg+Bebmo9kUiy4w9y
C5vowOEIm7tTEopNjkB7Hqr9uMuTVYbZYSv7ZTjvJxHULQ26Onq4SyZrmVg0eBk0
Rz+fF4uhx/VsiU4tb0Gl2cM3ORhFsHbF8baMkfmZea0GL5bSRFSOh+ogpbMQsOMy
MFVcr9gRa5hwkJx+DSwNaEyOzPEo6y4Y/QOPA2e4c4+Nr1VRybOuYWsGcTBWZQrh
dT8w9Lra3snsDzgbhYfjBCzZbC0li4ktmMEpextiJpLVRcOLk+l+Xb7XuIrZxikm
8vO4Kwi2RlNhOkU2D40HAqPgMxy2quKnwaErS8qARn8+LLTivZ/w+Ov6DiUPA73Q
qx1ofZWbtwFBQ2oL6ckeH9b3mvkE5yXVcF3BlQ5F5yC/+NheGyGNcYp8Bu3t9Cug
2A7dtB7F7zjHWvED9JFrhJFiDYdhaKnHmS/IFoHtQXZW6VHotaxI4ueyBiyOS8GE
d/rx5ogh2m9z1qRyCVIwsBuh/EQ6IgaFrR/4LVFKBIgCkvOm46sO6V3dVt/66OzB
SuK6fwbjF+kZFOT2YxCKOYnkea5XsGqfAiuADbMJnsfUt36cjusSUvecrydi8E/B
fxz+1OFnM56oiJhht4lJxOmKA/Nes3V8sSqTTe2elrNMlvs9qc7fGgbobE5oVrTP
7JSGR+1r/fBBOgjHMNke4nVnJCDUUCQhfOwSvYZsfRfJY9qefSotFPqHC66RSQdx
C4/VVm6wi0LPu7Qkj8n/3i27Bh/55WUNUW6wbQD0qbNkxHM6LHSNVsYzsSSUxsl9
LPQ6osuIPh2W6/FaFGAjLF4TxjXksmPtMSHZsz/DjEXCY2NzsyL60pkNzgMjPxzK
33AV294ESJue0HLWikKbvZT32HeeeCzmY0OfdqYM1btTTzpooWcrm/FK0356OjoQ
e/htUKdHbL0fY9IhcdZWPrgR7dW/mtuKhMUqNU8YVxmidKYNIzuN8ErtbNLUE+Sp
dOhnL7PKH57MOEsNU0fCHQu2sm5TP7wNcNbVr5TBPEc1gnFfu7p+UnU6F8SxuKU4
0ykp993OVicFq1aoh+uoXjsjrhW4CBfdhctoRcGWw8hZ6DxyWnpKa8/OFBC/fAGm
bYIlvr+yACMc1Jq+LD+56v6hbTYXy2NMLCMshmGgYUqxx1Dhelmrkjyv12wIFpeJ
AaTOTx0dM8Ym7oe2Wg40iOeYMG11em4wbsvaM5bp5Ztf7tLWl6lcq0Y8SCZUVHuX
MZAHxA2E1N5sTdMefBeZUHLPZpp9gWKz70ng4uueTZQVV4vq9l4cDcqMPlWZf1Io
a8rW3T8N8CqWyzY/pZpGBDF5cIdhs0KaNvfRlKt6Jln+9bquPpWTvJ5Xfg767c9W
pNqiheMtlqeVJm0TTvmfFjCGy1Mu7vUmDQNDuM4Zq5p5YORkvUW6k7/Sw1r/Rabx
JLsUqKH3y4Fcvo64OUFxUB308Q+Vpl+IoUq1XnzSx5Fjb9o01rTezg6lM3P5QIG7
sJie4CHVEKxfRvcIBbXmKseJ9DTvGve98inQI0zDOs/VuQEuudjpSCe5JhzKvK3y
Fc0XasI8d3JvysP8fhJkgdRU9/7JgrHkMBDJX+LM6Rwim99YcDlz4u62ZS2eIvoE
CtnON0EA8EG9ycMRgM2h7SGvSmIK1EJhj04gcIFhsql2RB+gpQ8OtEINks0G7G6i
gTWb4Xp9RL6l+aIei/Ehil/SturTf3+qyySYSYizW5bmg81PbWTcga9sd2OJEE84
iqQJmusKXsqVKKZTLLcLqoeudo7D7VhhLDbyHWLquVhvo2wsOKlNJ97nt3VKBWES
tpWUSWc3h3aiOERTkdRqWl5u96L/DpNxAre7cLOFgYmdiJ/X/pGNz4c49n9d/D5O
p4KM+Q43VQXzlmySoFumdgGxviW5B8m6I+LbXWOm/rO8VqLe1k0nuFRXPhYVuh3S
KgH83nToscqpxDMH38Aw9i/hlWZZyxtn6dLoeBZNTkjRpHGuQnT7PdA+ldmJrzJF
7ByedU+wopgyKR2qsH6Ybsf3/cL7eUGbZ9B1byD56xxpwLL0Y1q2SBU4N9t4Pk84
YPEgoI42AD3vvzun2KyGj1ywV3ERuQGRjaxuv4/nAG8FtQLHLQ4/4T25EjF4phAW
wQlksqVAC6M57mt6lhQJfQ1FU0qDoVKtjjy+1GAPvuXc/GX+T41qQUdoCBp7GVaZ
vybxXH44GtfndMHqYo8xGV2FGfGUFMucgosO2DfUnakycG/ESCyICkBtoFrjZEED
ayyG3QHzADLdfS3e07ENDdLbArdEWDlWh2VPnN2fhF1sdcuafOQapT/9VoAG7S93
J/G64ZR7gABIbn2VQWjrNPnc8bkwWNr4GsTVXknAiLV3V4kstM0osfwUqLtrCNcr
C0gYJJAunDaJqQjvbQbb7JGfINUcqWyhxZm8lR2qVHuV0AbyO5/f6h5bi/dykWd2
tTbp21r/dHOeizNiIDgEk0rhFa+4vY+pErdujfEkFBsoIkVWKQSk3+cV3Vo2rrKe
2nIaLgkKup0XrNBKKxVD6W/d/y9Vupv3HEVMjmiBV2E3QQyRcMb2M+QY7iGCxRBr
TdUjWy9Zlm8S/Vy4RiBw5PK/mMEv1wT+5tbsUV34cMRgEjiDkGcYOlAvTnuQHp3L
J3MhVs1crgFoMUHiS3VstS4Yii2Aaq52TdJpFdU1Tn8wa+4o2KspElFm993Yj0W3
VQIZsydkshYysNH5wIfGzfhOnPyVMvG55DFyiwrnGVx7eTAHi4lxmbMWrD6XBgMQ
YLW/ATEPpQoyAFhFsa1ZrKNA49IGBFS5avu3h5PKXOGOutpSuAQIt59espWemcAA
rQxRhuYvN1KE8TSrtcsX2+2/xo6a7SJwWCHoSXdSQFIjhayVeNVH46wrLtd+0idw
0wYkOxuhnwNSx+1jUIOve+aeU872SFgyPugCzm3m6MyCa/ZkBmWEcIAKhDsj6JMN
qpCDqxbwXK7S2zdm04Sr8awuIgyTBpW2zHeaKEgeC+1T+re8ghw07u28VJoIt7Zj
2j4uRdKZ8ccgJnmdLpFDc7VICp9WZJoLrBnvieVr+Gz7zFgmT/EalV1CEXPy19tp
VOftXl13EK5fjYqwKfzzcDvQeS9G6bHs5KSfaGAfGjs/qR+wrYI16yfrfj7jNcbJ
tFWvZybARwfGQnnYSxb/FVOcMNXInJCiB3Ij/kqxQ9QfnOHoZ9s0RFTeqRfCYYh5
MF235GWkg/l5xbk03SUQjR5GYpvpwPFLI6D3NforX2CTJf102Z2GDFjUrDYci52N
mQUH+GXmBUSo8n8v4dokPRKusZYEGcRBJIYTjZQKK6RwShrxp+47SDk21FHc3sD0
6Nzuh5G02S0FbnrruRVdQUTkYy+PhfqsWEquuUDn2wnjmhUPu6ygDL7RR6oRjtJD
d4vkvRssrk4j3pLSRUgekRhtcOSZeRvv29m+t6olJ8iDCBcwxOi7mmFL4A9jAfIr
bRXzGQVrqU7IPk4nhmLKPgVgheUQ8ptXu4nwrxXVUOQx5ZnrSTMQnORMsZLHg/93
hk1UYLe4cFX+nhTzGpRHylxeLujuegZxKm9mPdtYOkzEB5HV/d16od0Kj5JAagRC
5erORIefdkQSehTyXVb9tDaf/CrGnXelJJcPkwY5yYbNbP4/dwKtknkYXMlYf0kZ
QtfWxoGgRSsSOB+xiK+TwUmn/+/5/IrK7a96DVhXYfWCSWH5Pdejk1t+bw2VUM2B
KWQhZi5vNxvEApDcE8nldujsPP8dv8bW6dhdDWm1Bei4f0IgY/34v805iRxKQOb9
Y4kH+i5O23Y0GLEP+/Uo+znSZlLwwFHTkXS4VD1wgk0LRj43vcfMoSbEo6wqN8Nn
jZiNPGvff+1K1FPxw/ShkwSrwJAIZ39FMxf4QdMgVyyfBvG4Hiv7ZflUkLwpBXhA
DtWkGAVmxDYpsZYKLtUUtmZ9nrzNJHGdPXueTrNw8JMwE9tQ2rrHWrZdgtqABvMx
Rs8B1tb5997gFg/+G76NCL0tjN2gqwwEjMiqCGe5rxFeVxWNDwPLJ+q8M7FB0qE7
9BMfQoWtktQjjhJk9yPMDWxcvbvXyXbXFlUOqX+aJnT+FYqwiYv/m6VRNplbqzYb
3ZNWubiumAsqWnzC6Zhc1WWCUtcRspl6JHIQdrHST+bERrnfIOFvEoleNv/e4yj5
bmSavjn53nBSVc6sQmIfQBiNtA6H0xzvA5Y7T3lY4rmdXx6rbE963+TjvmjfLJ5f
Ism8HnQqtA9RZvJe2X9CUPfFAqYjWLwfd64+Iybra3dZYJ8uNnbrbwQuWTMbKtuZ
KvJdYoVag8IvvfjTfwiFe4dieaqB6f4rfvUi7uWcCOu305syACzfbQbLmlVrvIyT
7WJriju3/Aosb7myd9ms4Mes2lfFHFjK5vnzhvU+RxbaH/H+QTr2Ely/c1DqK3d0
AD2zx06sEzbDtSFfEYTY5tSSHNMrNpsy/uwp5Q09nFo9Pvk2C9eEoAevxKJQjV8Q
rSTKBsyRhTdiEK0Tyv+d2RFKUCWs3ruvKdQimaM6yHEE/S3k8QHxFpGrgP2LxsfD
z7yPm38W+70PIVGsRjJpCF/TWRczq6YpYSJjJJSk/+4FUp1pOH+RjAA1MIExjz7L
YGmME3z5jBkL3oAgLeLcZxyOO1fQlU8z/7ntr7M/U1ZTS8X08kweBmQCnlOTk+Gj
UrK+caHNjGx5ffQLO28fIrle7gKkYFucDgA+P1eHWak2zVBOYxkH62lkiEU4e50c
/h2ldcBLr+TCL9LrL5zkMyZfYWWbkbiwhM/xIys39BR7opVCgd4ysSENFgcxngAk
YvsDdhbDxI+xdAOTPcgkIhqib5nToPxUPiPrxV/MFR7fzbTKOHSWBJYeOkFt6AOI
k5TGyCr3W0UMh6e1PwlpivZGuhFdDKnliilQZbFPWLdFY/Kt0/zcrehuNYk9nM+c
TJ/3CR+SfL6wsWEaTwUgEwUPK5wTDfuL5uZq0DnSfbB5Z/z40Filoq0TvKS3SfFm
+1xbnvyTaDCBjm9duDYZmhcvQhGy4cGKR6JjLftUTpOu3mF++EFb+fc9nvxKYTBs
kh0irgXjY6JGbVLP4EJVOao7SA0rHWg624qZRoddDbkPeUj9LmiTZlHjAMizGdlX
KNBPZrE8m15nGAkjmfDNe6I+NQdValrvixHpoOe0ID8aPD73bjeqNrDHobPsy/mX
5m/3zKPN55jvd9lAiGd6X9pztnqRaJqxACibslZGLG7wswW61/b/L3cknPD2j3iX
JogVK9IdgQKiijfpSK4P9vpNKxjx481l4Zwo1qUeW1zMdV4427va32GssoXy6/Jf
422xA2SlkU3IvmZRTOMXe6w0T9/TeaxPVUhiqpU9r7UnPjtv1oY4H86SPc5bI68e
jlLFscz4veNa+u+fp6Eb5qu8BAvNo61Va6+PexL5nR0ahWetekdDaPreteR6BUvD
k29drhTyRKtyuGtqfQKiLLoV06QBWzZzOTc0JmPtXPdhe9tiEHZVmY5G+XIUMm/U
/Ke+tTUIDgQkpAxiZFErVIg6iQRenxADTlPtgsDp/D9Wfy+UChMKd1ZOdZxTWcb5
CEoq7zLxsb8UWWFCenSeJDwAj+9QQtfdwq1SB3aA5W+84w8z5evFEsdRRETGbXVl
WHKNfSc12UVTBEaxNRHzTzQ2/dbDSpSAIHzKVoDbFnH4bD6uaNk1W4ujG74u+BxT
AW/y+xNM+uDuCehmpJe1PaP0uGo9utd9IV1afGVYlbpiml2gLkg484LxH4VECn5o
IKJ3lxfqSFUvrNiBb9tuXTPXoLplrGIM6K7tdvjp6i33v1lo6S1QbZfSKV5vZu95
YfZ+Mf/ZyJ/vDcS5ZHqk9tFYvHQ/enlpHe5RuwpEJuDE8Gfi+ofk4UFwgUNmTMfF
+jf6iMvEKMSXHfa27nXsNy+TtlTxuc6gLFUIfh1eo9C4WsISIROdtdseDHaEvqkI
i29zLeiwXcygVliiBlFL46kqydRojWDA+HSxUIgsUVkd2NhPmr2ob8mNqeuGSS/0
nbUsCWVAaaYnUcUTXP0WQW0CpwUQZD05xBj6QOuD6dzQOKqBl09wL6qVm+Ezk4kn
Y8HPe29j7Ali8QVW2cJkaHIoBXDLAS4fSg/2u5LvLQEwQ9FuDQfxf89uIGHhUDy1
/ZgMUZ3fWM6DLWf1mMC/F7HU/USLM3PNC0L2H0DGSJbu7o6vtTFf99iyZFJqx41b
MRc04jhTa5Lqe1ixc0NtuB22oyu8X3au+ALM9PHEipqxpobhaE5cVLiGt8zO/QS5
Ji6uPMZ+xW34K/INs5H5Bi5fbpSOqQ18XUDWJPZp79IgYhUsA0XbynuyWYteqLtw
tDH1MzAQ3fVa+EUHqxQIlNDWUUT/HTgftZj4TutU2DJXXGXRQImJNU416BQqJLX2
18J2GkdZtiKibwhM5cD1S8sLcciHo2xZdf7Vdp6XgTx9S+JTao6mJ1Bma8BcGWka
hPNixF8KFnQkUXqqg0F2UtXOTSqOd8qyaIA/1dRokauRYcU0n328wQYJ+WpeI49q
3983JwlphcxBvmeNrRPkjqk/Cike4S2kk4AZeUW7sKgTNleBSL21qI7toouyD0mY
wKtMClwH0Gw7JL92ztiAyxC56dl7rhH86R2Dxfi2v6NBS7hilpK8hzTaUJB8ypSs
b+hLVTiX2t0HJlYtvLm6g7mnlpquQl12W1aR2Jlcz14xjF0/ncBWe8sWMDMFDTzj
MNWta3f71rnvSH9FqRqLcyW6ormbJRFZ+a/bcjiFoxGEUSWQCWIEJDZugvbQWuf7
ORSHIIKjYG2kJOifjrrlmA/Hi/NDcsHY2WDqqfbCMB2qGyNpFocNFehUNJgM6wLO
8EKyLz3U9WpKE8aBsjLjcpKVk/Bnx0b03x/wPo+UaaBCaQm2wqe9Ko88NgSuSsut
SOZ2xl4PUnAQKNuu7EkJ+PMcn2f0+Dni7oUXeek5NgHGBcO917bOMXUbzJNDL+69
o1uafkNe9g7lLY9Agt4DiQFd15qjNWXh2R1S+2QBr3gwrKYwtlXbxhdApEQC8NvO
wLMYruWcBP441uiyigzVwrS8o7DAg+AXCl+RVF3qsfy49dN+j9GgPee5gpMi3ms2
DPlaJ3V1YhY7/6l+3BDpBeuikKYlMAp99v5KZFfoP0wbH8a2J+GuN177pz/Tg2E+
2v7SQgN+nPTkOJnsAXOcnmaxLfPF+uwAfxxiCoN/MdRP10nB/jsyhVNGY2iA2eqK
5NoWaNSYQOmsGZpD1yJ4nQEjsNw4gr0NbvRO/s849rdQ9vPlrNEaX3eQUF4tfrjY
+dRcIjkayLGKILM2UIUslwyBSZ8/0QQNjAVEcMfzKi1Q7iRBmSPlXRyOrkQn28rI
bLJz65hqZjrsWlBan5YZ6xenFtB/YgyBw2etW3mr/UvD1w0poPKxkaG4bset5v1s
xIxGoOMUymxTd38RfXUQIinOFncJcd/xORSptg+Q4ndslMGEmb5Ud2LL6ZylMRiO
xWlBk1DYoycy+OHoB4/3wZ+Q3m2Mtbwoy2kbJedKsUKpsTVpAkkXQnhip5SOeK0E
jvQb+R/EbIZOtDa7yogF8Jb2TDDua6Hj8YQl3QldOOyrCmibok1kgMsL1IUQ51vN
iD0mw6GsazJUKtEkkUeJJq/V8csdFT7UnGdPaq830viP+etqBmCI0KuYmn/rZ01g
5zyPvNFo54D8qE8wnLG2StKTTROi8AHUqvomaN7pUrDwfqxIqBkmUZoDTGBAY5s4
RYZ+vNZIxoWWHcg/vLE8jtdW9XfvFsRmC27uL5j/S+nkVWOQ4hOfBJ8V1vjTJ1KG
pwslY0ZLmhSEkeZew2kNRobqOABrDFE6+SwrogiWRGoKeMGHvXV6Oo/s2O+yaDiF
L1uzIrITupB5RKMadKl4J+dCVFi+zQ8BAKZGZEiDgH5BDl9/xVxu2rz9Z402tZXe
ekY5TX7eKvkd1vyMf+tdZDDAV+mQoTNEPd/JnYDRvhEa3OTtVXg+Dj/2+1n0tHYw
5SjT7eryc26Nwe/p1j4q+QcYVojfP09yScK0X2JS3aqCOwYhX4WfkFI2StpqRron
iaqP75fGBg9np0HGfpKjf+fspeHlSqDPX+h/MriFe7j7x/47yBa8geoo1wD/uGq5
ZPB4ahWsNT6Bx9tTU4ykj3RLaYqhL/+sqN2Q9QVggaySGZ1RXuGNO+q7686An15B
opHh75QVXUVv55zd7EfyGHgHy27IhPq/XseRC/jG8ErGX5pI4bO1Y3RFjnrll0g6
uSNhQzJTiEVX+3rcrPE4w4it0RbW6Q5W4jbFHJ9wnbrD3gkOZpo6cVaOnVyTOPqI
lGcyQSb9pVzJ81yAy0EgwnP2hQdpjIVypNtFPJvDn/yoFeOSRPJPiou3uRAlN4kI
aF9z1/XiRfojGH07+0wlG0uHa62dahXkBg5zv4CcyKqIPLcAnvMA9/f9apIIPfPz
zTzuytWK6/1Qxhna6V6AVXzlWXcfD265P472gYPzv30rXhgcT4H/UxLG9Kqo2U2K
6ZMvtDAOdATWS0Tk8OeqgAtX3JKkatXOMK9OKZ5w3PXHPVQPVyBfX0AcIjteZYRy
xV4hB+vVHgg2tgg8bOAXF6vxfKO1FuRa7RsT1gywkUIBRkcC7yVZAI7U3E9Ylyvg
OApOcKt1Ppayd/DGbDsQXzMaBRbSvQj3LFZMkedUQ4/RU9ExnFnw1KWli0GVVPRG
1qBVUFR0HKQ6t+4DMjhASKj5pg8k2bx48Txo0XvQdjhkfkPkUM1gOzh7AOpcWbfT
rtUb1BU6VbuMaxvPqRBh20rxCHr4xbWZDoZ/qOy/3uKVid/oMJnA3S3OnjhwjNrq
io58wJ4pMtG3crlEvpGVsQwpmgFVk2GcxATwQcKx76Ql5XZh0SAWf0WmoUauCV8e
PwwRrh5K8DNpSDVgBtMdGdb7u7FL8Tm3+RkF5z49YvJ60l6VqrqlyCd2G6GY0Lq/
wIBfl1yZo7e6ZdiIvlARAq15+bx/gDbKyfZuEGZzOsQMWYJhly0TH9lUKKVdr495
7Bn1x8Z/ZZ9BgrAFpgZqIixZL8V/mvHmDHp4tbwlO4cjCz7fukvssRHS4JtaiV27
Hel6sEmfpHjiYEnXdYUlR7ja2N4/zixXVOLDSJWleYwF9WyDOG8ey4ag+I6ygZXE
l1qf+4cHV2KWsaO14WpJu7zAOplTk5hwoRtOODMPNmZ9o2obj2p5rpwhADviyu8P
1bCMxdFzHMzkAIGruTKO7IwFWgWZqdhuBnIh3Pck4DogHaSENsqbuW4F3xh5Q7gM
N4oYVeaeOSjy61Quvnqief6gnwRkP4F0ZxnUfsnv8FZpEoCQlGNEGrU8KLlwAhoR
YkslwAVNSxqRolDN585ZanR/caeiTd8aHthhTiORFXM9ltHREU4zI+LvVrz2VLcB
VrPimPjLuzZcvNvYq3A8ZG4TogUD7l9k3Rn/ce5Mvxa8flDX8fWMMV+ZX6na7kWm
PmVL5wopYKmnp1PzGZnAOOIkEWTQKgFzOL0u95tSGp3FxSizNeSg2s/G7lvq++1F
P+evq/YqHd5oCcxBSnTJU47wsiWj9o8RohHLLHDoqycje9l2OwLH2VmPK3AIiDXG
7vLwx+QU4xAGRX9Dhsd1D8Zt7Q1MqSjT83fT7JC6C4uIM+Le/NgK4ZuQHgUtTu1p
d//OyGUMkFgmI74PvS2ZV+OWGZKLJp4xrzgIpW5wagyNwiVjb3v1ZdqyUIW/1DCb
t2VA5zI7Nx7WP0DYz2f2MGDQb++vFiRs8f0DuADcHdE+FHoBckB5Xd/lya9G58gZ
oWCDbhRxp+1WgwFeFONkaz6h/4XkHPTRYucUxqkrRrxAhPlPDuLIfNQpDuLSN7aw
Bzm1XGTlwxbWPwNYfQilkwWpQiA+H3LvvTvfII1rdAxvKEagFIHA2pT18L3xQRGI
W9APkB5QxUExeT058NQ0s2iBAi4TNvlN/lcxZRkDj3xejATc4KU9O7psg+kI3+81
SNgorLxmUzDUyi8SBM7ug30O4DhDGBU8/vfah/PEOFRzDeTUf27UlFRBMpDWfP/F
YNbkN+viUGTjrs4qsgsO5Rb6qVJqSu9PxRKfs/vEI0TEOX7mnOZsQsWpWr2r+SCO
v3J81eE8sB5x0czzbxqNNZOCfOssYs+HEYlSbi30CV7gZcE7kbi102Ea5geWlBaD
wDJW2MXhxWE/uF0xUw68l/5gQ5YN2DTJgnLV4pQC0jeOPijn3lEHjM6G3oRc5LzA
WK1R+1yHAiYh1f1VJJDqkbDP7QgeCHaeU3m5XNkywlfyOPay8oEFbzPwO9Tu5w/1
h1taRO5L2ELzKCEeNCtsKc7vQseVcuTTn4P/EWixs2HXy6zGpYEY2/45+K8BGycU
GPPRlFvGtNmqcdBfuLTc/9YSz4rcxUyD51Muuh3cKJFKMYPLZ3/hGTblCg+rQt5R
Y3y1taWY4VcANN0ZhapuXB9ZGpb6sNgKreZn1mwbRuIFNibFJzB/N8NhdbwMoPF4
3HwMyBNCTGQEDsq6bQY4GU/P+eGFDfJCxGmbDJ91QoFKyT1meAXfaibR2KoAsI+H
Ev/h4mVFUUX8PmuydjJdGlqPHCMeEGAfSdEFciB1lnx9M8nWgTd1KZjohkj4qX0k
LBADoIBBX3OvWGKqkYbtyNuN59hBE1hURtPvIwkWoyYFXwrWVZ5pu1Y6kRXfkYC2
XiCe7cWPahBT7vKbhl89RXxdMKJjgbwcWYnXXdNk9N+kmhHx5zzLRTL5PkXmSxUf
o8E305ApRc8xsdbTIc9D4SMUOkIuW59Rcozq/yPN6uPCHgzifxerdbC31wJIbCn4
L9USKowITX+CHs1OLt8uPY3ZTT/dBAhzm3Qax2n7EKMWpMbJ19fQ17sfBF3P5Qgx
WiSXWbb7ib+Awenhzc9qEH42YRSVIj0LuK7DoakRzjUmD+22zbTl4eSxOR1TAjlV
N6X6Wf+YNr/iiJt7X6lSvpQACsf3SdnCXthBXaydqPoaAIv8P1YkWZaGjsGOqFzu
+UQZu8spplwknw9qAxWDjgrSpdyxXFbefnM2cJexdI/UhBlpN/WRF05SHXN3J1v4
zVAWTKocj7xNJHXNeFKoObg25vVMxHqglGoSv70xwDzq+gIyrbrvaCTXM8ckpP3u
Ehwv2ZSYqg/rALd2DQOrgMQXGxvdM+O2mFq6tGQZwdcDLrTVBLiTld7dvAliG1dN
aQWnuEcnNC9NkZ+USaQwscdoGR/m2w73ZStNT7MDYdZwuDIM5BbGZwfw4ZBd1W6l
cynQSAk3KgBscr7W3Q3Y/0CbXTNP7lZbCmCz3BdTYAgSubnMNv7FGsYHkxpUmcxt
us86y44h+6DLS7Ewyo+HrRgVcwqr5vdRK2V5G4M0WZ1iTjaqFyd5AKtMQ94UwZvo
fQLJz76lhFcsRIdFy3PJNzJkcT8qMsf6m8FPlWicLdVGBvT2I+kwZOCzKlKrz9yw
5NetLKeiQ1QYzsvY7tExVkR7vqzkuuFVoVBfeiIYk+hdI546bq66ORdQ9AffQ+Du
gSj/B31D1MDgYZaFkyt6bhXNlngyAzSwJUQ7/RZEOKjHlmb8j1/V41M/bwgCaOQ+
FFeTYW1D1YqbUQ8RC+05TGTfncXGJlUDnQmDVnxXYinVZOcbxfuIE+VqBL9D0jix
ckH6CwB04HkxbXJlbvVYFRz4qL8Y5tQ8OhVyp5b5ZNhu5DPL8iBKOfAyMoJJwimf
TSdLQvgb9DRecr8e8W/a3ejlhrBOiZXeawA7rY8wQ+v+MEuTOfq2LzsXP4XNGU4E
CgqiTTycwWErtoOJS7tGD+0ZDGZRNaFfREGYCU56lhkl2dU2UGUi2tcnOYc9xDjh
kHsRej6gWDME7rHHZEqiJW2mLj1RUVt+KFxCsMQBUs7XX3FTzzdtofMfbzfYZFZN
OzV2IQL3kR8tQXfyOTlkcmx8foNvNX5o5Ynt8LemxZ+PbMTQ1nTrnXl7Seyu12Iy
m+zGMOXLVPUWuYiIqa/+XXwBFrWNSUhJcn6VprD+lOLxKI39mcwTwfNN+P+Y3gCr
Rf194TxCmrCztSn0X68eq+z8rn+NKdwfkFBkxPrWDI5vZWc+qETg6r27Io04G8J8
uFrBGtkkLC4amkhATDbeCpSSxIVeVv0jONtAo6ySGwxBLjrzInmNo/uNrnCcbKc1
TRCcnFWdh+oxUYbPVtMnrykr1cMcltWoTjDc3Hu4o0nD0p5qnmGSCTbAHzyjujwa
jFieev7O+1Fe098HL6S8W8XOEf3SLpWnUrT5ajSssTzvC4vMOh4Q8CZAFAe+hdl2
U3t/q5VfCZLhkfCPgZT0jDJSea2vSsJtEycAEt9DYILT8bL8oBj+FjsTsL782mRc
yq+ZS9chc/hYQejGXAVdI14mOYh9TCK/5WviMZBOlXCpuxNfiMAtGxVd90cYiXLC
8Nx/SNe98213zq9mHrUIQ6mF79j/YPyM8sUkveVFdt4ymVxMOCS70bmtwI646abf
IdnWbXsYmsIpozepC1ghmoRulk0+7N8Kwup4kIqRKnNwe7DBJGq+TrHc/Pk4MgDc
JFp6DGdlOVES/GTwGlW2JsGB/psz+qb3zJUgqsYN2waOme1miUUsSvGBtGGk9QKx
uyroSMkd53xlRhuNUjD8nbMGHU4GazA5dOfv9MqStwcTnDu7GzF7fH/5N4oQTbry
autuCODq4l0yHXbeP1IVRIUXs09WDfK43HGK1VP80wYMfCpWxCiiPlx74JbcEfl3
25Hz6E+ZyM2yUB7n0fLXFmr53ipLrdqW5gdB5tPr1gxOrTa6mOMyar7XoRMnaT5p
fsKwx/hkAM9b1plHUc4By+NMZ9wjW4K2UhCagysfYwaRMTqffNBBqsy5atIbaLI1
j+gF2gGGYCTcdG4mNX34GdAms1Wp/1BKQgM4V9c2NzuiPerlNctd2fS1g6GaHkOu
BG+dHEpm6xG2Koo7pTLTSx9E21ibmWP4WzUdCiZZ3haLuuZZR+GCiBPQYRIfoRKO
QBbBNWnAgQ3Eu9eha4GJca0XhVzv54CKLw4nnr39Bnj+qXuu9EP6do2SJWzlY2QE
9rkQc78w9M8zYM7Vq3waaiEr2EkXVxmDF/2FeMMPGzv6YrE8xEJRsSMTVdJkJB9A
Aq7/8tKQWMx/DCUFgmSlg+4ZuRqKN8R6slYLdyPTWY3zQa+neODkGokdlV45gH2f
OxY0U2fSzc6EAXQFgFf7WAUpx6KEYGHQdQEhB/A8JZlq3hqfxLB//29nVZsseiXU
mMXTjtdV8/5qe1TylPJjk7v2W/MfaeyVoPty74Qs424xKGl9XLGaxg2jx4TGaXeU
LdA/LfbKBx9b2z0/PgB65fMrcjTaXb1F3XAtdTDqTouIKrkq+8UH2yd1S81IxZ07
CjV/1z8Lkv1aJGbG0twTEH/OPF1+uBsdqoyAVnYR1AdMptc8U28ARAlRlZYhw7y+
qYZjEpYs0gjM9eGVtg9oq0ax1ugNBzL8hhrFj7zw75c4A/F6E+YnHq8aiE53B4R/
WxFdWHRRKwZrSga1OXHUB4D0ffOsAMXnNH0jl0fFcemBjEnI868Lu21auJsuP4Bg
uZXVpraOBlAkPE6V1zDq110EFA3kAVeyQzpisRP8qAZgQBoBUlIuSlyh4zNdx9HR
Zr2wLugd6D8cHPdU2c/o2JhEfdaUlFp8SDPcfJDShi7jfH52b6eFadMABa0S810C
DzTZDYH6ztd+9Tvx/hQT1u/H8kmd2SNkzTLMDotppOh59QvEOHH309vx09wzugAs
DbJ4474EtQqxNdmZw510cSaijuJTur0qm7O4yWv8todCvG0086+avXWaZxxueTLA
wgxaqQgr+d+VU1+Lbl8zCtGGsGKrbV04HiFQGBb2TxDSTvk5QagGb1frzbVk6Luz
LfkVnwAmv1I3pFtZmx2yP7r8MMp34snhvwk/txGufbxOsN8zIkmKFrMV4FGS1lv8
f8s8xiwoZLw2rggKc+psDl/N/2TLYUQM8GXaxRNGQ9+PYY8aimgbxJQZI6AzXBMc
TO7+zKLNnUpQIeH4gomMRD9s7KnjYGSvJl7r4h4FneY7831gd1OLea4nRaJABlmH
bXKa7nh9vMj5U+ln+z8AJgohbMNHRtT+pdCB5q3hQx5arfeGj10jo+q3tg7JSSH8
rO5K0UlvqdKvaaNEmwT5S806un4r231vHizxDD+mxZe1+55GagrxDIQzKdMGqv1J
tVoQVL5izb1h3RsmgQ3eAmAKMybGvm3f2dwtDaQ6jPhfyH6ke4CAMhdlbLIW57Mw
f0lUOyxZWwmboiErLUb94FI8xAxKbM8tubtTg2SUXZGphhiLPOeX7NkguoU2F8UL
sEf+P8bUZRKJjsBtyFnxpasoY0fkj1PAEJyjAfpmMdwwIcJ6W26MjBqL1NybwAMy
Jnd7I7NCGIGAADV7Lu0YvnCeloJEGh6LbHBXy/WdzLqY+sx8c5tJW4IaEjIw0PK6
eeU68PCIqdgukUqkIbQG8XfrboRyI0ErIK/kk3j9Q+twGL+h0Vc4DLlt0PIAy9Df
vD27H9dFDtQ1aXu67cPW6NQN+P733W40wtO/6itB6RvRBE8/v9oywLalYb5ABFN9
N4aZqR0oh3jn6pJelU20xaHiFCClgWqZbpDveHptzpAxc2iULTnREEk5VylvFTT5
S/U87JT1fpki+O2jhuAvz4lObeeWp2Pj+I0BXqbL98HutkK+PlNIs22g7CEWvljH
0HrQ5pRbTiKhxDNtUPsoZFqZ3HksxMznA94apYbr0bhAzVmwsEKa1p/iXBQuxZAu
2RbG1GJDyxyJ3vg92Ws+ijaWrD69GBKTc8w4Y2iiFtzGDLBIJc/Fn9sw1TaVuQVF
aiJjFQV22Y0LuZs81B1WfnqK36QeyjiBwqRLnD7WzIQoN6wj05lbGkD4RN5zo3YB
UMT32oA2pTw3pLssnttplNoNEPk1XTqsUzT9oGawWHdnJfBIg5y4yCShYKP7aNIT
GiXFi+qfe7Yb3M3vtMIC+TF6Ss3L9GJAFqrJnyqlR4DTRf2KBcQ4QSMGI5wywk8V
dtDfWDnACrlaeT88+QE/9zJVYyui8xlQVpM+UW7wNDlHY/CajjTYEMAhLCE1uoBH
2eX5qGn6b+jJuVbGVqCmmUsMyJ4XzH4aM06PXZ0EJi/WwHmADFfCGTLO7vR6z8i7
AYevs6rWlNQ0hjs90TlC5L5CbgqQ29sPb5Y+aLPLXQ5u6/itrSSp1GyXZ3PLmBIS
iRNxjqi/GSX7oXf71GGuZYBrnIOgN+G2jl0sYMPNjva4TVFcxfzxUpIfJNBW8jNy
2qd9EjiLj4ID3dbuh9IQsefoRA4qRqCw4HLv0ppiRIT9j/NhuM0pw8/atImLKIvK
cOp5lcq16wSF+G8V8JU+zk+3O/4U4pm2RSfh3/akLZkbq+m4zQ6XkhwKLIdv0uNM
ZTuc9IupXA2GGvdBFdNmnNlUAv4bJzRa7xvcxXzkxIoqgDxolUZ3VYIK9RrGBFRL
SnUYp4jDSJp46iOzxjDcMOP9FGnrmywxRIlMstelPF7nmKptrhXLR4nLayVolHqO
k8XU4S9+JXv1WcaCxTcdb561py8lAzZDrfqIxgfYaEsIjnokxADXRsR53HhI8sJO
0H0bIIGdLAWyMuq+bADM149o7Of9S62SaouuKmL2aa1HwKxridXb3Dm4CLbtzuRI
FPUCQ0gMAuPXrasLnQb+M2nMvXCK6KhtBer70ROytzLtJqNWcEqiLZTd+7hmhmIE
Hc35c8RfKQsfkmZZZvPKQWHuUFdiJBTMw1uCFG4kDSWBXC7BUub3eWOLcLV6JAqu
NC+Uj8o+awuLm1cwq55qDbXmBkbVKC//sseZigC5goz2HmXsJgxKwBdv2lOGzyKb
OQKRxsHHuGq38UT/8tSBwyzxzWDSVg5pwCuGpXKnAV4Pi7TnWQg6tKM5p8eOK+/+
bMorDNIi0Jt8dPD9I4vGXvr3XcIXEgSwAcVfFUV95h98i5FR/D2HKgco7H35g6iF
pZ5UYVO+lsqfIufyHvfLZdvohGPtdA326qSlgC0hPEn048CIv2X3ojnHYcQ2Koxj
ExPp2xX397+JdhSMm77mHYHLGaoUEwYDY82qrG63LxRFQhWTcV00OfR93CawxbMg
MpFfbANLad4zEayAEUCMrn3emg6bg6fbX0SaDWN2QhMkoZVFY7r+U6u1GviJeL8H
fRWM3VgEl1ZtO2DCJQwUx7VSPB4jyMyczjHg4ViOtRFrBPvtgs/IzoEtGFfoTowp
qK5f7o5bZPy14SDU3YHxbqOgXpLaEYPSRiuMXwLRat1+z7ckHt8d8043bni9HuKG
z5bQeU3ubXQ4o6v+Frz9jlIHGlM8qshXZ7f3frZR4wSkq0QQz9wfNK3XTFEgNYIH
OiMV7RTfOCuqTG8Zoa7K+ULSxZY2zR4iAG7wEYSe7MfjHxFAwYmbhUdozUahubsl
AUosIpIGBqQF8W5w1lm1OrZNDYgd/fi/Xn/lk1k4+NYGYYgeVGfqlOBR4CmBIb5z
cV/tB1puiEklnhBIsxA4sU8KSpYRi4kM5QUtw5jDR32NThThr7t+d5HuAy2Q3rJ+
cRRdZtDTLZwZLxrgBio+/tTj6dJdn3afjG766NGnqny7SFY2klHcl/Lu5m4u+NAu
HRS8SA89FSAM3H5EOiWfgiOKtHfFOCPWs8b80pyXeEpEBaScc8w4mTWAPyxdBvDf
VWqrDnmSAtdE22sMajwgl4GJkuFmVJQ8L6tsqc3OTAIJLEGjQ3FpbcBzwapbOtI3
uCAn1FhBPCsfB9pM22bRHGNFlWanBsaXeOjdnBDVagkEyXI8UFi9l2MQbXlcxzEf
TOJWh5Ux08j4u/RxY1u5Rxw9tC4Oe91oDfturMbl1DBbn9YCb3oYokxyJkaS16tZ
FTHhXr2gBEl0Hx2SGbqjwi4mo7kfciVcldMT+aDnFtHycEVNTVAPiAic8o6j4CKQ
pX3VvOmdPxyRFQDotk/wuPHMJXmoycPOu+CBY4Kczw6vUz3hqdmp8TMFinkJOdzb
csOvka/pXy9RzAftuh6boaolC+jlvPewY0P/buBFcn/cs3Z3nJmYbf2Jh26gGamj
Hsoof0YwOsikAOveUQ0tUqTngGE/LYW2heuaflMWSiDabOf3ZP+RqcieDzmKhGKM
2YzFxeG4pOEvFTsiovqNZVOL3c9EOWQqZX4iH0K/cTJSwkP9Sp3muV9tcj8olgK+
Gy97iO2oq77mXxcWtTyoi9AcuL0gSzFnxqbz9TisROHRWZ3Bme33PFg3ut2ONKlS
5YDlkrYtltgcGwktymeSrF4/fH+THc9FmyR/uqxKBmuypr1AVU6FbRIh2g1SmdPp
Ceu0Ojm3d27iJry7Kz6O7vCvihLdUF3OXSSfH7KxsPFCd/TYB1JR6J1namIECOix
xj2lTMzC2T7ayG0h1CU3laux7GrVG1dElPoX1xi2BLWiebqQmJiiTH8DfC7mz02N
g7LdC5Ufk/RS6jL1PB1N7l8zcrlembSB9CbCEu3abQSNSXwH4pCQnuLMoNRLl/YJ
VdJFWNqaT8q5sHRwvDTTynbDLinuvDt5wp0LYR5wDSH7Mm+NP+H246uQlkRbjhtu
8M8vI7zptTNmY2tMTPqe9T1rcQlOY6oytD1+n3YwSW824JbURQJaj2tKSzuB2p3A
PE+QwYsojz2PLybWXJlQlC4dfsgtkxuszqamMdsCIqOnIEfuypdPI9PFypdOhZM5
e4RzMBv32R/3//A772RPVH8TUssNvAapzCHBqtlyllE8ttVwNm4tFWGHvtLde+i6
72Xz6SUMszkHQzLhq2JNG73h7j8B/wsR9l7IEzg4yiKBHGISKAzCyF4vK0AbIZE+
9kV8ENWh2S5gCcD+kUeIsBW0MKKCAo83mSpJTy3al6YL/iTAyhcq9ByGL/TP610W
5wkLAk8IUUkZ4sPFqLn2s+Ui4dY3Ybr6VTIxEvnZoKDePQ00yoRoJxgck53uozS2
U4tk1FauUrdgUbnKCdaDeorbT9Yf9PO6Yqq0ACPe+p6VoveDF/ywjpj6oLeVzJkf
8kUP7msHCARoK/IV9GJel6AZsXSa2YKmpW3CqiS6hLNdZOWRDAFwnLQjwXUn+I6y
gXfn+THtLyY9Kj8pzk03wWMzzwuxVyt3pBOzY1GoV6CMQc126ASH6Mkwt761ywWn
FNNtMyJHl3z/0y+lUAfaWMm1WHgbQWlYgWNYunCAjGgewoHoAG8lp3FeZHrxNN3+
xeY2ddreuOGdKcUR8YSYK08lplJA71r54nijGZgy8sgPnP5mE9GS3gI7R6Nrjj99
zrlP58qfAiuy7EVRxtBuTbBdIk2pgOiwK1Ge1JqD8JRDTnA9PzDLYQTr2LmG8T8Z
enARa0z4h0UbXgEvp06oB5jQA9XaFqXO7Z8uzgAYFNcF1yzpa+viq3FflTWtHmkB
vOSyli2IiMtFlPydsMBX+qhOMerFSiffMoWrYt13fawBL1UI1EHi0cVAz2Qalo6+
L7HjmOdq+8VaHspIGVPyRy9DBnN1055tNyDjuQpbnt4TGRTENS7xhx5D9nFOytOn
dMjZDEjMoaVdZhpPE8AefDNTSXfVo1F6wgny2BZSmkEcjLCeUGlMMB8p2gB046lu
pp31WOv6Ns5ax6c49ZrEKTJGDId40VNdRNDlHubETIrwlMtuEm5tYwSEiIMR4NTQ
A65pPWU4J0xKfyiA2u+Zjw8p4sQMWL31hLlB4aPuyClwJ506PkD3YvhwscuRKII6
hizlG1h2GIaOKydZRxdG94kYM8d5J5zCOpDStz7ASo+dZFWZH2UWr9PgmnLSw2cQ
XrroP6Lhlzx3vlAnOO2zb6SqXHnR9C/afyPKh1viDoLaX2PhstmC3VsPd+oEL14X
kS/UsX8WB5O7PsrsWtTP84s5RxVUIbFhHn4RoYt1YrXvEQz+83VP4fEf7ijT5V0x
sW4lyc2J7P/zEmLF+JOTkD2paTPJuJjqvufO6PZGC9mYA2VqCUGhPOXSr0acnOYk
pkiUZpE7l2kif0FOD/ItBI/fXJrWA7GOr3MJFT1nFst0TS6S6uWTzl8mGnuUAvZE
jL6/SI7G7KG3leR20Uff/elcWUk2dwdU4OXs9GjIXs2KONJdj8PGFrhFImdiMJR/
oDPBeBNkIPGS9m84/p4Ws3GHY2iGEMKbF67zNyQ1zRXJ2FkiG2YBA6r8W2q288Mk
mdXNy6b/0rD3HAbh6NBGqLl/jGJ20dP0245lMsXxG3VWWtI4KPkFmK9hB+Wh4iGa
/P9KloZyujkN4sFny60Yj90OyzG9fujB8XNCAj5JRsHyQuPNEQe1BWykdxpEpY1s
6P/FDKxzOBQVSUsksfp73eBdR2wnXcHuyxqWJ9YMCocChyprtGCaGlKlOfcAWCLf
mW++sdKtYcZf2exoxiMKmmHRjImU4AHPAjIUH7UmTf1yUki5w3ekGbSipPlhU8ir
V99GZ4sfzykk9gy1+Xao1i3bGn6y7TAj0TycVvoXG3q/nzqd7Rk6M0co5oKTZ/QO
qH8q5Anyj6kF592HxQHlopCMLNpCRCNevOEzLY8gml4OTIDYU56D+U2HdSCS1q57
xuucm2Pyo75jS9oR8RqlM9/ew+RKjE+TvhanzbD9eDTmmbajnFdgchacg55SUPnr
GgsmHZthiqA5WwAVbfeqhdlA3HP1cxnpmLLEHb3aYEBRTUf6gi4ya/hpNr8dWroi
FmWAubuqe3k5x+F0VSBdAXCnUc0R3txezxXZ+0/G0Soxd3fh8rpT5Brgua9C2V7M
mfioN4+j4YRj1y9zp5bu3FLmK6cVOoHR1OTgA/YHCOpp9KQDPKbbGIw4S6Lj0tGy
JTs7+q6pu5JkiZyW88JYAVE0YMW6PWWTYBWgWwIVS/0iqOTP1IQ1L/Qkt70nEhwj
255/xIs5QxruTr22ymbyGeJBLNegiKqHCE8fg14+1NdQJiNftV1n36kJ0KTENEEk
+VZm48i4ZS+J9qf4cq7LQYCi+M9lOR8/m3VJz6xNFCaBMTh4wC03yFpPrD/E9SnR
WAdUeNCWZn5gkcbXaye/cTFvIE+QmnySKT2Bl2v0/d830hOAkTT6hxmc0qDc0m56
vG27w/A+joayyc3o1P3c7zDONayFcODOZSCzWI26tZcByivDsNKTKH4NlueEU2jZ
RUItnhzRfU8s+UofBNV5KDYXZqn98vi7VqReGmHoSX5gZG5zgOoE/00RDSLN4aJp
bkbayYn+yBFrHkTokFOm4UEncqGjCl5bOfNLAODZll9NxmQiCg2CoTH2+O5fcB6n
wpwTYq6O9xQMqToL3xUNNky3POQeuVZ5mhpwklNqZgq5izbmJvScgYmRGGqT7ZXx
uHmqxz8UzKgcqsCAgHmLJM37Gr785SVAIH9GG5Zl1cZP6nHokYuiB+ITW6UiCJcJ
6fBpYqIxwflsGm4dOjbcwG5NmCDVnsoKeftcNs5LrSf0kKGeElIQeQJtZkOyGwbs
zTIB8HEL2OrxTIlVqAM6eutsaY5t7ymwtLPi6jP2KohcqjMFJsWwUi7UBwa+A5k0
qOx8yIfhGK8/lApifZzwfrdQ+m7iBFVGh9MTTykWUgb9qXDhB40ASKXL0uhLrYBM
g5PjijjjpNpEO9XLeN/fO2gSNOBeX2ZbwDxIGA8tfsJOhiUGDca1TkBkJn4BMD8G
13p2IPhdjFyYIl9zKFYmwHVoaEZnRGquXpw2FmjMrydMeL6y5gjm8s00FA2leife
Tm61L5Uh+n3zb+pz+LQVpplctCEIaxmBc1DUrZTtY15N1NysNCh44TyI1rSGMSEM
Dyv5JjfpXxbZBTl5DRhlfFuIRnWLFcXDYUlFru/wvXiAJLYDzZixRBKtGt+dPzKK
hoxW2eRkOy6pLuRtv+mnPjf7kRF6QesHe6LNJGPuQzi17H6TnDs211jSU+65PWdU
u/Jw622+9cwuRblg0b5ZZuUolm98Vv6qcL/+5zBP7mdNtZBvIT55olvGIOErksSH
hVNKlAi9XHaU5q+nLuFyH2Ti2Ct3MeJ9dNkLEF1c4PGZ5cIZK/YjKl/e/jx+NUmN
jM68h8NBW3lBHtL3FJuFhZXiAqnGF1BOOLImOBQ4wkAm2GIqz72Tv0g0GvKZb3UG
6yeIbPwwVYuAEW+Q0fnJOISQFv1pw/GQY18SzzjYLf2RSI+aWsqCn46UggzotshC
5oWlNy15Hv913EAfOvzvAkswgKpgmQcYqLEcDNemVlMprrFP3R1ZPQyi5IcilxmW
GQtyqKY5zRe8emESHeHYlKKctMu2Kms4QjvCEhys8CYoTeB6DcOX4CQfyPNtsY9N
uFyzJTHXKuSUJM6rHKyKsjOFwoDDxJ5qemCXnMAyP0w1+2a3mwcUbiODV1NaJgij
vbNoZOVNymB5kSJMah23/fD6dGti1iuR3emuwKHof0NxkL0jxDr8AxaqL4upilt8
f8l1skAhY7/S5q2pSWbogXCKn1qAwRz2f2GBFCVcd6RJTef2AgIfy5jMO3zEbfTi
OycYNBaGxkKkmc6u9wbMMz3nOKJQSEXPn8EiaQehoZiBnzDsesTItzjasf9MQvrT
zHpRfH+kpg1Ht7VtwRdpdYqPL64xt55HEyLOb8mlHJDRVxtARa/8JsPY89PSy8Qj
dbnwagbNYbWpng8OfSuG5crdYSDvrL82PBBw2a7bkc2T0FYFTDPWhw/AzJe2ctWt
XpskiReLCcw6g6p333nsUgs/6YxqQJCk/RmMbWP7riZTADhMIDjYQP0savhpuasr
q0fQZpy/fyQksrSQ/GVlgfADm/Gmw3gsqTstMwTESTEqiC3sOIkvZbwqg6JNbdL9
zShPWiOPxsKDMKkssZRUOFqUt700O+YXICU13SP3at82iMKLjmL28xDCO5JJ2XX1
82+HYL2xP4OUgFqjqEvK3UTdlHLjO+0OyJ6zfln1gLX4QDM+fXwCi7+DH9vQtU+c
hp83dnJVKoNqkWE4/OnA0/pCCyWyswFmdZBvkpZGYP3Ci6cWxBupiYs9afC/5Mdo
L4hMbIjMAP1zfwQ83rzN36kzK5Mg0Owcl7t7YHddbX1rT579JM11gWazNYHoInU2
Hrt3y57cV+ULgCPR3gUg5uCS2EQ4pSC6e7YgCvsrRua8X6qYgXBGAxz9AZK/SuSM
0NIAP3MW14Qaq2REiv59H0ubTL0iGJ+Ur4BhbhAaoweuwe1/El4llwbnxXX7YEkn
chr8+kW2ACEU81s5h1JybsERxsdz+L3fyyMn9U6qKX+qUjcOi5jCHRvfxYsQ9aE1
HAvchPlhP3RBQ3BRinlWO/XhFWIlo+jpV5hwTviGXJZNEDN6ykRAqK+CKMakuBgC
WJqHZKmcgOBNQahLSNPmMtMuq6Qbk7Y3rn/rQIA3dtdMdY70vUF942Mcq86th9kK
/YxeH0en8EZwuzpHlT4OZG5y8Rz3vP+zG+HOI4skO0FsViugwHTZ5HEcpK1YSK49
JIa2inNQyph6hr2jjIhicfVKCVdN3DY9SOYg24wgnmqVvv/CJiO5UtSn8ptGclq+
X06XSXB189ZiBAzIODFYaC1hH/VnydFmNEROZQiU/UjjnFuxSadm9ZKTmExJCR6n
wXJZ6NQTBjHPwyKb2Z1CoI4xHxWKoQaQcnT7S52i4s8/R8ZXqFmDqkvyPWX90xhX
hpl4tT14wH83DUtk/6DosEgW5CnFBLigmoiqrYLKjxbYCiD4c2CK89YueutUlhy8
Ob9KtxWgSUlRUxkorsqZXas6ZvOCS3Z4x7UIsvDs7z4PE0Wpo7Oc46jOR5wgRT/7
V9TTOU0YYhO1NMNvL6OjfrEDOy58nj0kCJocAtY5bOqMuuYR6iglLmN97Vnc6iIX
34ViddsUGqaDgSKgfD8t8DHUsNtzoD2bdFEIToS8eQPTjHSMv4UYTU1tWIb4By7b
mq517q36wFrwu5i2gRPgSXC+OVhIhzvmcnUYBcHlUbHg8QPWJTK32l0sFstXhV9C
VsV6j3ULQvhmsc5lDGa8w71zGLplfOwZ7vJys3OJEM+LC6KFcWUvAJia9JetBFMA
IE61im5gyQSfsHqUhjpScXITvp5XuskM7rHaFrt9LyZupIRKecZD3JSWLluvTkBJ
KbpUz2pGyBbIpy6v2HIQ3xwDVSHPgDOyPqvVwXPgKwOYVdIzgXimgsd75TKydSC6
VpBm87rZUnttrZw5IITHs4b1odKGESneZspE+JmKUCYlahQZz4usPlr1bDsij1wc
LG42UA3n7noFt9CL3tF6sDRZzDmvBUrCI4AjXm+a3+voA4vQpBpYkz8qAVR7UJpi
i2+3Ikk61VtrjjD0up3OSc0qkPvCJM41m0xyTwDl6p7CzAElpaTRFAuK3cFMXSep
xXcDoYCgJtq1UgCgZdPvMXzcVNid7zYIqBzluPws83C2xsUDoog5oeMzZgnmZ7qw
zIepqn2KafmGU2yNlA334N0fo9zkHdpYjT422Tx4nuqg4/ZYLrcy8KsCjbzhKviy
L5R3T+CI9pNQJWqBhfHp4VQRmlvq5sKxoaaT1/jb17YfW5ZGLHaiPEsAygriDC96
M6Cq0pHlR894QUjGDRFRUR/vxreX6COLiRRPFRDY9gQLqxm8qnIKFTFKW7dPdCUa
GAiC2cdXt22ULR4xGw6mUwLQqSb94nEwB7b1Lv0WxUcgz0irMqJICHeBmRrtNe1y
Jahp/kZHVj9s5u3fki9ru5D43toGJDydsJ0yjaZ4NmnLhWjVelNI1WKIRBbgu2hx
IsUyLo2ugfnFtFrXZj0V+RTimSB+4eipZbZd+/7mc3v9EJpumWzQbHd9I//duRXX
nSb09S/+Kyi3H4UD9h4vST0++fcJBHD1i34reRK5OdVEMvashooGC0kEKRTZ7Usn
6HD2VbUe4t5oetbRIG6OB9cfW9AFGg+Ni57Rh0lGBv96W2125SWy3hjKBZDRqfw2
pEsHC0RvlaH6GShXDNnkrPG+ifdthM1ksIOQCvm8+NbylKMMtCpDR4HU1qgUobsn
cEaJ+pumsp5fxTNTQBpXX816liK0EW8gXo0i8V/SNOWDMYh3+k1BXzBJdJCVv/Ov
Yy9bCq83XbMyYeo69WVjvTw6IXCxMaQm9SF9aYKfRbsKdRinhIbAAirwfh9AZE6r
ADBZndZenW+7cnHMMPefO+tRzBrFfqSqNzOGKh1uKl+ce5fZbUqRM9o/VeP0UgF6
XKe3UpolfIM9/J0qpSLBLBL3hxIqeVHBygZxbwqSjJw7w+8ieOrt26mLoGxYeQiu
KIhGXINXY9xLnBsWVNDv7KSkbvODQJ2bcQbyQtfZxNKzAwqC1NGKNb4Hd2oyxKmf
ze5PnSjfgaVQL/cPEJPy1j0N9xSu/jCwOwyLV3UWJzx8vKB93NgrF72Q4gOFDN4z
/D70cmukODgyTUnrgrivXPeQsg4ASMCjLcz0/KlVbiojPaLAOpg/oNOpBzHSP30p
Vz0wtbmGLwdF56TDJgFWuYhMMOJ1NNEJasK0VOwTZSARqtMWFrYfj6YA09P1n8h/
ArurwTJuIZSA8VbFTLfqS4/vPYrDnRjToaeQTGmLMVxane2oLKEKcuDm0zIVr7Cg
Fo3U1GVqXShCokwqjPJJoixeXQtKtnPIQl579OddfV6dP7N5cln4fKOkP28ijQTw
NX/4g/uwBaertcrTJ3Rx6a6bndd3jvT8SpaQK7Lmi1ecRPn3SljwDUYlO2MerN9u
8+kgJvx69Qk+UuQyEjb6VCtUqfYBFD0eb/m9aTCu1BJld3unDr6i8hmB1JdezPnX
HehK10rvtonLaVUtiCCAiWuOkxM1fEE5MU9MLUU0LMxwntOlpj4JBc1O5X9ghSrE
LYYg9rKQI7GYNJZI806ZfhXPOfuzqUhAuET1MtFY7Z9G2/H3E+/0/1hkdkkdoxvU
F/zRuEIxrVdU22X6oXnoUdFsK85am4OObGl8KS3KU5VtpVYNw5iPVvrjttBBjKkq
+qsIX8CGBLYncdx9cDhnxMupgkE/qIclO5ZGm3fY1ZiRU1Vqi01B1WZNI56LtmXJ
kYXnSlLUFb+Rxeswhn/Xj6/fKSLG+yfY67wgRqFMxW2Qxqmx9FnCSgTN1zFFpBXq
oQx44MPO+URKkNB18XDqgrQPnqjtKp1PYiFxhrnm5jiQQ09L+23O1l+m4/0NMRDr
QiiiNo3B+lnp9cz2UuDcLccRkPdJJ2cWJx8ks+vC7tJRHzsTu40eUEG/1Xbf0dSL
AcOFsL1DNA0zRztFAlSBoBzhqZiU2D3C8Bbn8MrVqNaUBcBBIZi02iueo4SgwRAe
134VQhTvmmJwOFMIj5dGbnQfu1JbTI6k2oOVySt+/jZTdag4i5J1j60mfsfPShWV
u3K0clKADvRKYWXovE0hnryk4ZUIuT/Tpn9dayd0xHFuNU4eZtGFEEcM4J92yl60
kHUsLYjQWDncqOsOU1bF96qU0pSfvgbLc7jXdUlrj4/vWkeXspZYfVICoQXoMVBe
ZSpxnT/uU1+0QBh551OsERz1OXfjx4efp0RsxNTU+ScG6q5ThHdsJXvWt1c11f3D
PnmhkZFUqsfaSiyxZcxFw/PJva7McNdZaVSPCNr36kBdlKIMxYLKyFzbXI1Fi+MV
+uSqJwlIEuVckKugCaNskYhudr5+j7p0WOczlaCakRP227FUddmYRbNXWxN760sY
D/JFGQ1yVUv7Eno91pRYTIdC6ytOy/Jzuml1rEDXQJS5Z4d/L6c8q+x77ZrfeiKi
dKM9V/UmX41xRD+jfTQXRaEATz103+akPaHz+upWCI/ZpdOAcVj5IqB11/+K9O21
xSOF25CYtvnOJrCaORHuendSJaeBVaj+cgRhsly5wLWPgqQ4c3QR3YRU3BIqCDgE
z2sj/dEVOHvBI6FAjuX+M635jNrWIMnf6VOGBwy4RlGwVDzcOFyjQAfATtvvHXgh
H0aQPVYzqR62hLezswNCs11AlEx6O2aupGgPHzWk/s2QpM+6/W1EMwS3NyO7B2h3
mCYMI0CX3XhDRZYyR8aAbCnE1jSI0LBD3m2imFy4NsfA+xas9GL7fSVJSfqZ90ZJ
fs404PDFFWmijriZZ5FR2USJr97aPnuB9yfZ8O3Gqeu2bTV4WCquLgeLYInngrWh
cNISJFQwsUhYCt4E0tcvX165v6yHH6NynV2i1PJ+806Yh31GHa1pA/w/6i5QKa5v
UJzOO0s7jD0vjxV/icSxXVRBs2QUD5hrFlkT41HMAdzMNmBIeVQ1scc8TBhyIiGe
9UvviVXE/LuWQObB4RU/4Jq/ZMNJRmgvadkTfmTssrXaVk3NlaeKsxqmCJZ898sQ
X/vUWxKENhd6F5vgJwAMGES9oLmyjQ72FVX5N8K0hAshtKzhpEGfbJ3p/PzKi1nm
5n7kDro1pnKctsT205SqT/fp3bR6X0lwXM+niTIERrlIZQwutRec1T380Vih79Jk
WBRqR0BBvq2bi8FyN2KL8SWXIbP41mnOqPn5CKKyub6CJ+cpXlFBXZshuJJAy+5D
HDQFkYx5KeaLpsb4yLuudf/RYNZfnT7an73NqAFKBySShe6fk8fGvt+D+kuT7JXq
J8T1LTQHaACZ/ohglmA51GOHmcGUm8abC2aSScxjQ4eo6vRhf731XTWJSsKYNaoQ
lkNH0AtJdK7c2pXy+1YXHDTEJo/LAQH1nmULGeEXuicXVwi1seess/rhdzKMt1or
Zm/+Eida2GGNoOVjvJOngEjrBNaZfaeSOc3uanhbbyp619knb483dNXK8XNObWtH
C5Q+8j/0beVFk3YQK94AzgB9tPgrc/oIWkLRf6aBo3k3Ldod5/QrSWoOLDmHMHcN
xSA9mMWSTCo3KMbn6BgFXCcH7kc9G7yLN+x8ev1dSmPT3uOVWn0sksvTyxJsJJHg
brDveAp0ePnMuTFEIsC7KtYR5/yM56Dvk9XuhPogG3Rfp5aLytaK5EjRKOHJAQd2
7yseZObZ621THVJIJGfd8+IcBM2dguWKprKURCtH+bx1RBj+S7cb5lt9Bg6kknCS
Z1UitgZ0UcRskf3y7wu1OVKQtK1aSV5aVYmvR6rJuOO/dKjVIsfR/tClHkhO6GLX
pfVVPaVcfQ/XLKqeNZGCXd4xGrSDwtuHsU7P3ZJX+RSIGNK3PE1+G6T17F+Z610A
/omvVF8lx2sqab+JEzjH8bLjVaS+1NZOV1QxtUdNCNxRw4LtsYWJmS/KKX6/cczS
K6n+s5LAPs9BLTNqo0reMEFKFQB5EUcLO1jwQqKOFSoyskrDANlUxYGqeXlpKDWR
RQLlQxDn7HYQkgy1rjq51amoLK/2BIqn2eNw/Jl05l7n5D5SMbI2Q2R6AnwdEKQt
byGKqezR9h6er7eNCqZUciCctYThOS0oIzK1FnTkUaaHX6UN1eOMPaTwqeWDjthf
2WjBo8cftLtrsiGUvcZZstNSvsjW6wwcJztFB5JrYctAeYrAGUAMpfA/Pg7DFzbV
Iv1GDwsyF8OuIMDqAnMkpYK5ZTToROiYApcUD5OHbHgkF2Jw5jZztLDYIFqogizW
TIjUqSoqtU+QFxMXgTRnSBzFElUnwRAPKCurIh9CVoAO7WlgPgzVBGJoSx/ZFYwZ
irka7vqW3hlGVBKboIXe7RY+KrIXcG/72zmr82shm7i1oMyRLyxawdVbu96qkfjB
a2xElMnag12pd2uK+TqKOWJCZnrQMyL16Zj0H46OOHwLtCFGOym7YxqJ+BRqqDjL
LHfa97SqXdTJV3DlmW/fkTBR+peBJG+APAttSmCIHncI3sBAhQz0DpH6af2f9I8h
KW42Uoec0Rvf+8uTjGeCVD9FN0wUAcQqhkn6WAYPPhY7rlTPUuMPEdyn0k4PzBuj
ub54EBWqTaLETxqv9bwsaWIwwfQNCjyVzcTOUkMhQ624aOeah4BcJPgLN+ecjJ98
kFjz2tNdaheBUW/TWnWdphppOod7BzxuK8a+bVcDJ0wxQ4rARv3irVIipdBBcA8k
v8jQ5Z22Qy2OY/gpBcfYcva+tdRSU+QxPMmBgCPpa9aIcbBGX+l1SX5B3Sbnu/Qs
O7xcH5rkd/h6SuaObyeNV1FfxP4vlbAnvX9tlRCzcQbSjPpLztVqluQSiQymYDFo
NwGe/lcQbnbix7sNXJDHyg6m4+Hh2c4+fVVpt59QJrMY7NbJnjyImg6a28GmPcjT
VFbubS1GA0TKhbzFrDrVKzIbUeTFo8EUt/zVp+xcECyzm8sII4XeRnKsRLZls+Is
bcnmzBqohLRD1dlTyjJdQeVK1mBHJ94jbxomAb5zyJOJG1jxjAX0y3SteipiedKK
NVOVi0pv3x+Hebk/e+TzbABOF325a3Bbu0Y9wyZK6pykeMljprWBVeP47lwGcVOn
OlC0iCn2gXkfYOnirflp7qk9iLa03ldjlwR3JEQccmhLfWIdYOEiUX87wFb+9mhB
hdzyTvCnnjfYhbDPpj/T9AXs/bQNrLmMoCKFEVSDMU96KzflSWWGBW1z3n15meDD
L7gDvhMpqhC4JveqHgueigYmTWRsxVk7y/YuvwCa/Lt6N/SnX3n/EYT3KEW9EIm1
4PvnX133hTlegVtN/T+TTVLUMG0xw3QZ588abjbR4XNDQByDGGkP+C3Fi65M8pkS
oVhL8RqhVmJWscGSSEgowvOW5a31L9LFl5X3uCiV4pbnfWBBSGYs2UEkpCS44Ygf
sYV9OP4rhQtbMiD/P70v9Mxg0B16bai634mvwYQ5yVfJ5v6wgrT02OR6NG4TfOEI
XBOUf+OYZEJGMKurKOyJ8u6UWgJfjaW6Zw9709lD2bhT116y0zF5D0AKD7jFdPDR
nFFUi7ZE2jQAb7iBPQNFhiqG5IqblaKUmo1v4+GIyUQbZL103rlRNm9q+v4RtHXe
zl8cdJF+BQiFgjebJmuwcVHKQKJZTo6vFQTrXXiXef/LPGkzTpXdhHsevsLUI2HN
JP1zy5dK8kjWsJqAXLm4igNvKEiuJeWFjsse6CkTvQHRR/pl+gRQ7HRaRyGcTRkb
Zt0o7f6auUjIoDGbOJPL6ELmox43cp5t3qv3Id/NJWNK/VxcYpD/ksqMbM7u/rE7
oFyggkOS40ifXlvRpbI/9gfjPNLcV02lg5BkYqpadlADGZxp+quvU2qkkvldB+3X
K0QIxc61ZNa8JfUJCSsVWQ5acBst0Pnj+yTZj76BGYG2GeAfc5jf4NRxAV3bQAkW
JRsX0EmIkuN2bGMIwzfMezVEYGV99i6qPP6d0SAlXZMD6WaGYqs5fmbEC1F2+aUJ
i6ROgSBRuR4K4ImgurlIekmwvWC9apSKR0OM6inLtSdjYyPOj2liy5gecyEnhDPW
t6SsxjwSpGEvbvmfTFNDoIoRx2ay9pgChRdecw2BCCSoSdkpOog+5gjugB9oH9n1
KhY5qechIEi4kD6C1F9eFU1koCgCVE18P9ADdNCqNsuRuwkZReTKAL5DUrM84r/v
FPLBzGsAqLB3z10h7ICo6gfQYcEVxflCt4Yw4zqhs0uUPW4NStVrN+ESHei7JZZN
6qhX4STXjBKWhglSPg8QR7W2jVVfPmfvf28RSz21Bqo5gRU8AXbIU2z1+U3aCLNw
xq4tbSZMun3c5FC6tpUupl+JG8O+pD3xgm+XUSCpo0nwyx+ucAp+sOUg4KuOKEz5
QDl1wjKYQ9kGxftP+qbLIGYF8u2BgqEifPBVoizALLgwveYv94Gn4i3CDJHKL6p9
DqwxqpVixoD00KJzVE1fsftnoR/O7MSDyHNZPY2EsX/+P6Vjrm1fP4cZ3dX9bmzd
eTfEerwjrLNK8eie/xGPllqpGQHTALzAfhodum2STuhwh1XM9VaEvjELIFPU6pTr
G5MmE+4EEVEgfXNdtj7RGLSQO5DBJWffkgqSF/EYS7sduhX3rLDpMD0W83gGWBId
j8QjUHAa7NnhwFtcngNLOUG0iEd6Jj/SZNfhRJaGqtHjiRwX1X18uZfFUysDjj8B
MvHXk1LbzuoXBGaWs+jg7m2GpSN4MA3jYUgwuQ27/oJYQArFGiqseh5n6hjFaQhL
SQmXr+u8xO5ovitTb9Rik17HhqJuNrQs2Cd8Cww6XVaTreZPz98CW9hf/hDE5xS7
V9blpoK1JZbLfEtVJvT9JlqdzlPneGZclC6sxdhbMwwxZ3YgWgAi0L/Zd5YeceXp
81IDAQBluofUuSsMHzHjwVi4QrlNvCDMEnd6qhERVfF+HkedZtetHlExIuv+u8+L
YuXJIzDvyb9U/3S5WgDCq0t9FyzgtJgnJqEBcn6szXJkC+lvh8T6wJUp6xzVn2sm
vznpAJmRwKCKJSm7OLWxkKNeyxV1CtHECBSZUpgKVfcLMSuohd6TBnrn1n1k30Ly
F32H/E5gYyg3mkwYQT3J78A9pcE0nH0/tz0GqoTfBZXPAzHBtAGd1Qwi6cV2OhED
NT6R0fnSN068trsmilpUHu1+LATZ/QAfMvDlZjaIYY2JJ5j7HbVYmesvSW8rXBeB
2LWFl4DTuiTQu8Pr74vzuUVIYrTzMSaYzYP5KfAlF0lxWgBXr+c8jU7uoZ5Am7h8
EU+8i4iK2ArTuodopuPhW3yfq38M7yTJ02NyHmyQFx+/RKcGOsn/IKVZA1KwW4oh
XLuN7OTq9y8wHA51u/XvlRVSR3uLf2rg33vBzZ02i/VnK6XGpBZNnJ+KMJyplJo4
S8CCqrFcjRlDYsLqA0uae/5csQSCAanpKjwjG9FVPFFNvJJL7O0TLNXKc+0Wv41U
yAZd6kAfBwL08pbHR2vSQ3PJdLOTjpyskbWIXJvyHs5d47dvzEamE4dduw+EUH1Y
9ZfXwBfAV4iQ4pMD8E4khNaLTEPYquz07h2sbhx5piHBnnXW9cSP/tnfpht0BZ5Y
2OVXLwePj5bPQdChlBmM+4jvA3Ar9BqUNEWpHwj4O+qlv5/WXQjOISMrSsfX24ti
mqfujF557Nxbyr3iODvwRpfGK9R0A7hkpVrY7Uim6uvRuR0OGLeweQzF8AdQty7b
YVWZDLWdRfL7Ce2D+qXtstpQfT5EzoFuZoM3oDg5WNKhj+mocFp6dbUsX4AyGu/s
v0FL0sQbc1sNOEDIxmah1Xxy5SKmAsq4hMbRZW5P2jtwXQOb2ih7oDL+ZEwJmyrl
2fbtf9vkxZEzKK+YGW3dKx3iNCqBtJKfxbjc4EodDooY6MyV3XBKrNwiBh8z4g4Q
gLzwzju/YBJRnQRIqfBUiIZb63VdrIOBJqlaVSMEUiBfBcymfZ08LZDOYos0Fs0V
/1d9ZB8kKMoVed712giXiXqOdVKZU0ou2pxCfQEtMK4Se39cr9qHytkthUulTqPo
btY0X6Y3NcUNtFJDjjxEttYjvT2pT09YsqHngUfrskpJW3V2QU+myByOqJ5/3N1s
f7jMfsVdxsc0rp9cdUyR+D8UftQR2wt0IPLoBfAQR8DYEYy7kduiJ9z1/9kao676
7YO84zEmMeZOzNPFojSSGcLypAFvut0gDNMjoISQQpuLIvsEJcIldWkF4DXv3Slg
My9bGyY5KIiCPqTNAWFWokyNmlPTgFUPZVFY00YCSSUkcMAlDVZAWCLFjJZBY7i8
rF/wWdNp7QuEjitHBL5xlSTO+YzCoVGOHkCCn/pkGNAWtSIcedI9HdfM/02Gnh5l
2hqxFv/FoSVlxCjA6M17DullVr3Hzy4sTYU+/i0c2VHsClPkBhr4GCE3heeHxrz+
+fXUOuDTL1cZUqTUfbjjQxYsYhz/Nph1obTfdLKzHNsB8DY+71K2fbhJUW7ZYBdh
0b9Gy5fWUwYVIsvjmgLAGIUlbOCvjACUaY+GG7zvVCGsRLGqtPCDWs/S7+G6MWkX
ul1nT5ikFvq1QXV3+uJppOATESs/zbpSs0jB7pHAaioe8oCY9iSL2mlHuY//IZJW
0gZsBUw4nP+agk5bQZlXcPlb4i0UiFeSnH6UfeSnbTyRF9HvgDPAZfSq6mVfNPD8
XaX0viG29alUZUp6Omj6BaHlZRehsreXi+l7QwMIOlRMoAiDxG1u0x0aa5+EA1mD
+vvrgU5Nl7KvSFOSEoU49Wg+ct2HZLHNKnU6eSIXUSdKSpuKTBarNdeytlPU0PRj
V1Vbf8KdWc4gOycy7JfwylLUHOwlS960oX7Wr/7oGZovFKnn+FlntFoEEJu9y8Dn
/67Cum9QxG6btNe2vBst5KNWN9grvVGDOblR678PZK5+GIsxzR+EcmCeNy5rjVnQ
Z97bi/uRebC17M4OA03mmImgC5DvKAx5H4nlgFnLeAnVuTc6YJyWUZOHEiJxz1PX
zv6BBeaMwtfxuXsZFUNU5dTE+SJn4JMzUThWGjvqPzp8esl7R/V9GXgNB2P3pwJW
fBzNB/VSr3eWKYpQ+CXVjPAmeZik0o0dFr4///ioKdj95C8ui6LpHYxYONYns9hX
0qacwjzW5xky3LYiouhm+X+Klv/8RA/xm0VjpMzsx0YCcvm3B1BCkLdqX81ibLLp
JDqi1DtFtHpHsQCJWgz8g9ZGDTka433QpLzQRX8XWKE5+dixDemPgZA3R7xbXv7s
e678ZsBvlTqnV9ptDVPYk2W9C87BO3U0/YxQH3LcJjGQj2oRc4yQltO3SiviaCJn
tT+DE2GFiiqb422XytmhMQVCP0NUQvaR4uk8aCfXCo3NLy3etdGCHWBMgQqzh2u7
SZO4vupMCZthFXJVYPEJbAOVgSmLovhUnq7k2QcqD9N+Em2smpRc5xHE+BovTHvj
TCDJunXUdHGXg0AC9cThL0IibAZ9hPMFtDnSDU11PJE8kScwYHOpqDSGgEA9kB5k
MpY9sVmqgbpgDcp5AnS+F8zBaDDr0qA72UoE1unY2OsU3dw88fpGyh+5RYW4nf6h
Akp1ONa20bZVT3G4BzicR9acQuYZYUjVuuK1OZlckR9EmX73mC5iKIBYJF5YgooE
yPctVoqfywgGIN+RAdxFhWOx+pVD9Nrw+n026nTPki4vPnrTzAcZbeVpIKRwlwNH
EuTbsC/BL6ySujqK38pT9ceS4wd0SoQGckodSjgY3Q6ic9hKs5vEaFXvSArrc0GT
4J6AYvdvTcL3K3VCQfBNhDVGpLNKIaCJ56iGIW8iV0jrkQpDyYkhg2ZNV1Jb2Eb2
8ITxbxTa6bpf5oBTHkj4RQWaH4wy5td1EFs98qPmK3SjYSHJEysI32YkEZJHLwbQ
HI5UTHPsRmQjDUg5ONQNqXn9eixj/q55ZWb5CfzrhrrgkgC0jlg1p1mub20vX6cW
+JsoelHbQj3Sbsk1Vcr3WMxc7osVCOfPL9KFqKgL2z8aX2G34frr6pMUL7Mlg128
OGk/Ot7T/iaMfQy4cyq7sEqdabPMPfzlHJJZ/iUmaFU=
`pragma protect end_protected
