// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mnHQyF87nMLSPX1I5vO3KDh5O2MKEjB2HdS3gwPsHqOUvIx4/N1s7LxYoElkYcGA
kUCH1h0nAqAkUXkeFax2InflroeoxmQQbfEkIjBndZ2w3R6Joqs3N9qdgTbK4QMR
btz3UgpYiJF8VRqv7Zz6hKvdw5h6j3V5U4GAmyfvVM0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8992)
J7E5eClmJWm9piOkRwydv/zfl3nH7wmz7r9VI4moOQFHlLXVZgA+yvUgXR+ZdomF
q3Ms9D0avJXlHJjaqJ6YAEXG2PRKU86BuxS6wslQrk4B2YFVlcVBVDijFUtln5Lv
pg7rwwvAXifVb1HgEMHvH5R8igTtjvXcgKVLipVVrOICVQlO0q6V+RnaWWlofEwO
F3eqLHgMajx+2H4jZo1ieP6w3h+RXxkvlFbgmVBEUJh33ABsKNkdnZ/zZ57n/LpF
BQhM0YcoQnq2zvP9Oetd4xGyi82sDBmk6sY/VxgOgREbqqhHOHot9f9Tii6lPUx0
PiTJhk1p0bcNcehQSHe5O+I8vZs0j7/X+mBMAEwurzf7RLwkHOvIZiQv2IPSOKs0
K3jnUC49qOBszJ7mOlmnPjj5mzWWw32n6yrTBCgDFe6DOV+UFEpXR3FN9jsiOkEh
Tcv+PuTfmjkezyIFPtU260ljre8gjQBdDR4jUFh8lyXSzHw19OJofcI87WSekgVR
eAKuF17RPLdbfvznN8ppSCXbyNr/3mjr7dI2v0bpkqOkq3GXYZtsDxpZT61UGy7q
ERb0jH118f1ZkFyvW6RRtzIEwsa6kZx4yN9khCmKe8uz9lBcjZ90dZjjoQzeRpBg
hdUbaomZ/Yv9AiTBJLLKfQLc3fnnGeO0+K77PODlAK8jA40hZ11Xbg2q9Y3rTmcS
OaKwT3Wzud1yhj/glObU2UxOwDRU46ranuhlM6htdBGcUFb32JNFEiQGuWSzZ3wb
jVPd5k1Tr9uPze2Tnpmil1T29bseuYhG1cYsp4YkG3hCRFfU92l+ZGExOrKEGcd/
hlLRY21+NJY68g4rr5+WxeMUwi072fQ8QDKmC9bP/2lh5zUJcovpXzKK+6/2KC0H
nzAMMi5Y+zeuSM2q7MiSA/rCMiOOj9btLsd7pRFn9Qk/gHnLkZ6G8TGSSjTyPyCz
zZ+roTHdgDWLOQCeeEivznhR1dbEMZjV2yhn1vqWOslTK8FHJKldhe2mjOpcIUT7
mI0/jr93O5X60IDxQXOGHOHM8XM9ij+TCzODYfwA3obEBJky7grkihDouLeq8xhi
m1DgH7GKi1AXVlkoUh09O1uIILAcrGSTNWblgVT2AfMpmY0aF+dCcFE3nOJz6z/9
lWXnSK8ViYbrkFaVLJHidxlFsjutqFaNkC0tlHp9eaHmeWPaUXms0xqsNShm7rJg
n5+asGoT8sX4LoK9xSt5d+hIFfqfEUWPjyHs1v1nCN3xeudzjIeBVTUeny7rPRaf
MPjSjrJL2a36Mx9DE0a9Z+m53KPN7LnUASnn4q/TDjVkMehIkphZgmJLsYHABAt+
bVl7ensYoUhbq5pwOIV10bg1NLIxKxjKK7PvjTFTywadQDL2hVf1G812a9hUREFX
yw9uM8vUG8R/VTgo5tt6JCbuNqluJ79Lql5wko0MGcpwlt1XGoUl5kQTsCyPkWIV
6vm0u34XloDrBse+h48LnSokB+Y+CdcSn4s9Q/+nPoVx6wR8JIRBGF9vBPac8+xl
0ssdAjlfNA9GpvFwumiKsseBXWMmyTK1NiLObkaYgpLRru2whnO3bZoq2C43y4z/
8OP8ZNzYgGXk9HEQOoVqV9YDxEdy2ZRoMjMYAc8+K9RfEIL/yXwJxayc2dn2KfR+
kNKbSv+aLx50RyphZj8rbL38m23RADTao6aV6TUVADsoGDxqtt1gaYOU/hVocbOd
NSEIzOUL1m2wHRLyLczwvcjTTfTKGW28Kfcvr7YWScR510e4a0shlN65FsuFimAv
SntIaMMna72+mEiQIQoIFekbsUHwSrRzCgvC7Ac5JLzDwTX66CeWARII9UYUBr8A
K27VGSXKFRohoQGvRHXHHhSlDLpFpqUqFOB1zO0pZI27hK5YCT5HUZYW7wjzdzHb
im+xzkFvNS1RGCS4K1CXwb402SfUHWT5IpGwoh8TcqeQaZcqo8EGYAkIz6SCQBAs
cuILSggVfBErNN5xYTQRhs6jaVFdhUPHs8QuCONo9W/MmaT68oYmyH7z6iamcqhp
gfTKbqfjzHsK7xngBARY0aXYC/sQCIiIna0dnjABB/E2jeVZFugDZqN2Qdp1os0K
tckxnnwoanXz2PKzwh27+FwXodJyGIepcaiW3ODqDUd3hNcSRTRLqfHnMGeesZ8x
sW/w+6TH59xacyshyyV/9k3/q/6hIgiTFzIk//3y0QEexJip9iCWvLqxsVfiyT77
xjnslB2wiyjvKLz1Wu9kAiWZ6SBTqU8Nbx9+5zvh7j0YX9ohEduQRIOSDX9TqEWV
UxvNnGdu3EKM0eGq85CHhMnfbMP0CgEeMu/gDL+U/cYoczhuK0x3mo8PBndzLPem
xarAv66/GIgL6xwgM8DFkNuBZsuJfHxoDZucytTLmC7YB4ERZXT/LM5TIvgyXNIM
wkln4mtNlTABBQMpgJDkb1yOAFvj+d0zyhirKDoCDPdGFhTl2fEFCAM/AADCOMQE
vbt2Ep6vCTkuQVqaahJtyf4qNzIn2BL+4wt5YapIQTfwsyUZHTFZDkqrMVzhumBv
Mc2WAMgkfd6PXteVnoK8IIgudcBZDy7AvANyoE1UgYZiwdrgjww+fKQwXUcOmya/
bPv0CtjRYQCU2E9eemQjuqMeBLIlkhQ65h7vcJTiysTyIy1Lb29km6ogoA+SFOXa
KSzXu1bfAERovWKznK/K7o6tPetB+9DVmeX7JMNY8qRQFi4LNQj+02+rKD43SXsZ
s+WYCQCED2BQXujhVyXnxavvjdUecTydfGfMlP6Hwu7HN0CY6kldHb1gBgERdB3t
VHx39QLTr02+3mDMaUyED0lceReCqXFFgnqch1RZC70NwyzwAb0QH218cejAhtHC
Xnk1VhlvrYD+KlJr9+3SG+DHgtuSO9SGUXcBxq+bQ8OdZjf883+X05hpS7/M31f5
dkuEiw1rD++ZtV2a6CFmubdBXHZ8f2E2IH1AENKjRAAoEwo3X5E+jQ05tFxdTcKf
WkY7LpFT6xUFz4GmH3OycbKjeeQvYaJp6jLzq2nDa3LDoQ49AeniM0nC1AaNBWMh
vx595awVziiEz0SSQy96+o9gNcRrX+4cuHXHQx/nK67ndS4XiuDuMnbfpFauwEGb
6ylSRhG55yE12aF39do64lAOe5akfIEE/9pAzqXEBwPM1/PEQx6sAwImIz988yZI
jcAbxN60hbqaqlVtbTTrAbai2giLUagz87GquY+ZgcRc7CncM9FEXev3CloZpiQP
KAtTJlTeqvLclpHo4u8ZCncAfksMp2UnbLpAWboXMMckCmn96i4Otea/giE671lK
P3prOzzfiMo/dwpBJbcLFcD097espMN0VTPNgcKfePT/WqeYN9JXd8EyY/oj6DvV
qcJvWdi5nqEnXWr/lNFMdzhmnJF8JDykbiOBzzWE7fRnQEQbntm0q5m9waRkhxPw
PlDRXES6BgLz1lvIbxQshhET1j6X3v+wng2xfzDVZsad2DfECFTC3gCoQnZzqpiT
wY9zHxi/Gg/lzHFyQJv4N5E5H7urStBTTK3xeeDWwhC6r9fBy8aLyzV5AbuTZeGX
onsUqKk4FuEjff/64XxczJ2Q8HSji9bIp95tOV9vfH7SAtpQgV2acuAuq9KfxcRA
EKeVaAxc83DUwAYOSLfq7lgAyeNcIgNTyB86H6CLK0zgf/BAwMQ+7KD9bVl8jKHP
REREN4Q/a7fcV3oa8B4ei6gNWGxv7wvGNBXhlusrGtB+f6ZBVLZs7u9GacmMOMRh
jAXqNTgCGnD6tdhqk14Vpib14alXKzeB7F4WeGxO/F3uJPfPLpKrLifOYa0S5tiD
e5Scj5EGTd8YEj39SyZE7oaEa7EbAz3GC/jTopUOdSfrARag/AnRlEZ4DcezmUKP
/EH9lrlRPggoLAen2HJHqLCf9bnCFWok3QZpq8G+lgFgxOzKRiGyIF5BIkKMa5tP
oLcyV7ktSKqHcljeeL7cdnkRXDsOTpN+R6MC0D2o4Fn2F1EZ7+Jr483+ci4EVsUf
zuX7IsDbJrt5Mmgxkyie4IWK0CmnGFgyG8KL9ng6lDFCDqRaLyyiZSJnreQAS8YI
kBIcMkERBmizknyijB4eHYnqJVEMwifxr65nIK9lCPa5swsh2IiNEO2zumfuMJUO
MToEvMPKWCAw5ZK30MqXBoTSX48ZLXwv9fka5/3uUFNfWjuBQyB8odQwYRaQvF/D
/jg6bi/814dF1kcB72XQYt1pbD9Qmvvm2lDmO0Q7ZFpR6x3CXyzYSfTfGiLKYruw
50EZUWrB01FPu3XNhlECKJcZ4h3F6vvHZPN8PsCo3uQCCyJrp15o6y/X5B29jOKA
LSgH62qcA8VL+JCkjgKUc6sZtcHbcqniUjm04QeySu6JZK1BEZPO4ouHzNZZaPq5
YL+7vabJ31tpcdWtc7uJycu4UXlx+it8t1x428e9N96Gkdl5h/ViKbp1LhM1isA2
wpeU4DxZc1Xbn4oK59ntYDF6OLmpIgSOwROWljBIt0HEaufxOzyBfim9kEx1EExA
lSnYh6G/15BggWqWKOabVDjPAF6GXrDpebtirNE/XRENzUNYITiKxLysjEBkVXf2
NMxHu24Pods8mRpCjy2bs13HH3QFlwmOxcKAhfb+IcI+DE92qtjp0/oDgzA3SNJg
haa3vv9EvJjx+q++LG5ESSi4EKSK+ZSfAy3ctfMkGb9+m7uhcPYpkwTWFI7XlPY+
Ue5v6G64Dl5v2hpE7yc0M3IGZPIoikwe7TaJAnKFQgpDOdwu6nAE+ZkRAdvUWZOV
IWdg5jPUwtJgNTLGuv/q3Wd7dUX12ulej68ZaS68dJ+eKpFy33niuOKn5Cbezm//
nC959PcwnNm0jsk9dLR8cNfIl5FhaHY8PcA2uLnRmefNYo32qegIAvEZNNbMTgKG
ezvOFBHcTUlJfSJ1paCIBlCBscCaBzCTjm38lmwr4g7K+zsDfXdW4bmS9gRTVwZH
PjeoYxlDFZSrzTPf+VrPwFrrSRzCyXRdDcBaaw2OE13XkKT1IUFP0l9w/SYzvXzJ
hqjYI2KkVHnEperjFj5htcE4NXcT88Lg5HOuvZemdCbrH+gULDeFdyr19POn5eGd
q1lMS1hGtrF0fS6vfRxliatgOuQtvr/nuQ7Qudc/2bKo2VFXw1hZ+2ow8FFBDtJB
gHvlu2QWfGiK6aRx2eJqsjn02soJBb5ytjBP0XwqFIGvgmbFaaQgYezWFPDtLVZi
H41kcM3GfoIJhP3+dC45iCUrl4/XJerhg1opji+rfnNtJaLn1LdcqYh7NnVlBSjT
HH1rJalRDIBx9QPz3+v2M+A2fLPeJq4JWHoSC75SeWEiGfewUuUvcMtl1HhpFigv
XctB5t8dOyt/58MNeWo/tYMaCslNAO+fhd2R/SngLzRFAiDdyIKShTziwTEGhdMi
BBGeDle9iyxDHrIYS2f5pf66cTBfRFthr0QfXlu5Y0LOz7pfGQigeoqjXMtEidxw
5Mcx9yhEgm4i12jT2r3jkhDgYHjApqJxE5ifOTXFpCqFYeI+EwaZ4U9w/FvtZ9y9
pMjnET5q0Du3M5qOi0Thov2bMXz68GgkTzIcDRrcTPmyvhIotDvX2KhNs7jBETBu
0Ce6vVX0UClUTPB1+yAZPAY695IDbKu79SJh9rglPfLkXPsMpfHg0Q6Duij2rRJ1
X/GHcTnrF/nsj6hUsvHd/blV/CBpQfz7+4hySzF9ZRt74Q7xnmpE0CloEyWCr8uP
cz9nf6V5/kCgh+11DiGpuYDRasUGoYar781JcI8PQwXHrjjLrU92UtR9m111Bp1B
RgaBOyWy5qCrGDnDbaKAH70jMxyV4tKf24W7EfhYOSnQWYgXpd9x/C6FT6iCAzs2
jDCXGQt82lKWlPcUqW9jjCtf4rEtXeREDMIwmsp+IAYJR6wAtFzJ/Vw5TNMOoMXh
lN1epyDD+sibkALIUcddTRGw2+EtUx2lA2eHwnogauttc5rRu2eH+Rl0S01HR394
iarIP/UIvEWVDlZg0Tu1MWxktl0l/XAhui+P1ltadtnQM+1vL/akS/N3tLavJzLc
VMI/Kkpq1KrgCtaCKRhsk2Y0ZYbbXBD/eddPLD0FAGQKBm4lJfqar2CjWkZK1wxt
9xBuowu+9+uJrhsFZWgNW0TPYadaqNLd4yZzZgejK6+E5sPwS8W4dIDNPD4vChU+
5+9+sFf3RVdN5qx/hPRn/1tNO4wduWJWLTJIp3wWklXUik94W43uGwq1wb3uNu7j
9gcPS2PabQpEMXdDxwsibNKhTJtdM3Q2VV70Le7gEl5PsULPYJ0bY1LM6mCUr29E
sXXvB2XQE8CIkcicLGVR0NqPAlIbL/rc6FRPYxtwgn9U1NnY7z0oe2G7MauJWX7F
IzOvJj0+xj3G4HSywcKo7xJ6C/diXzlj0bUoUzLw9SYTKu0KTX3YTMX8Wi5fBCuo
yZFclDfv8xVOpc52pydiT+BDw7Bkni23w7Yo5kQxYx/R0E3EQxFzyo9V4D7d+F0h
yKgp0r+WPO3OifxAp92YQz8Qu34jkrn/l6WsfZAq8lQAb6JMxVzXXnz1xSPUi3Rd
DzkpfP3mrxTgCk9RjuXmGUodJNrJYNHEeRFntnRefbwcn2gfMMPZKNQqJb+TwJoD
uycY1896zQ2bghNtq4JJ7Bu0yv98oMQrq2/hAtvhAQidi7VAvs0ugAohdQkAhZKN
HW65R3It9mdeHQzR/cgA6wBxyy/oMIGFyHuyo3lG17qXAvIbWcqDGF45mNu58dqR
61RywygJXsp3LJUUACz8wbMYI2Llg7rdwuv7Po0HqqOr++18P6Pq+rlZBDbp1Pzi
hDoni3k/U+tfhD9m402Uk56vSFmS9s4Qtn9bxRShxBYUwqcndF8//p+YW2QU8nb9
nb1pUprRcV6AsvPlhv7rXj2jpckyXNaTU9ZiJ3SMo3BnVZD9+7RF87J0TrDK4rtG
BETGQwJz5GZR+KRSG19dVXr9tsTK7Iqbqmxa06vAOqNXns4gIIVGBMw0XQMIFsnO
BvlMqBg8mRsFQNh4Ykuu8lHWBXFM1W21bm7h64HxM+IrDUsUID8mvNCAmMQF0Oss
3v8kTdHm9J/C4xyagH55lLD4yCnmBaIINLHIc53qmA6BFmwZkKsqlrM5+3KY/lFZ
gNUxZj8e49IwmD+lVoWgk8B5gCZNFXmxBcN/elemgX87ealpOxSRXJCp6HvK4Tvx
mysDQAUHsCgGVFOKRJOwpZ98NVDU4eDHS3XOGdvVx4glVP8f5H7L8HoYzs9Qz54u
UuFIuje7tDowvR1ZbYXa9Gb240COpWsastMKL++8bkJkhKaichaLfsQbT2A3KTGP
KQMeisvK0RnW03Gt0+rXLRFz0Au7f9RiORYDc+5kj3JGb3W0nTtYEFfwXbQI5LAf
JFWr5RLld/UOco4wzXrtO8ejxB+31XqUzl1CXqlULlSsbAc5ERrzpvm3MRqEe6Fr
RNdsBTIrlNmhMhiPo4tHzFwcqJwas7CkPB9OPHOUtXtBvt15k/9J8isjSYBGGQd2
eS9HmMeJPDyoE78dxV97F9bRJ+o56KLNmE/o5Ez04EBO/dhrwVt3DnY4a/0N9hMR
cwmDVfe5QaTj35mqwPINQX2lD4GhQGOwF1sd6PLLWBsbNzLPLGW3l17XDqEaVN1W
oL+Tmf2c7BVl8u/+GUZp1GnAnCVxA2wglS/yCmqYrKhKBj0pepLKztoXd6oOZrOB
vZ83kLLfRXw48erv/FF1yPE6txt5s397qqlWMP7s5Knql1abBVJt1tKa/DGpXyXv
2JEg6Ml8C6dri6w8gB+jlBJeaJorowNpVjMLFYr57Zl33OmZS/AA8+HaG1pOLmvD
6F3pdwhoMCMA3hwWuAeENcnraY9KDnMtFsxDr46lSei87RF8iUhGQL4wDHy6BDS6
xbzOpnvS15mUnzL+RfMENZZKRhUuwaxf4ujmSAXJlhubVa0LphvRFFuiq482fwnP
7sBfmiKpJu5UKdhFMvzoBqkX87gjqybm9QV4exxwhfgwZFeNS3bjHi59E2HFYGpT
qKpq3nhB5Cd9XIMjM2KEF3lLY1Dh7rCEkSk0nt+refqltnNpo1g48jVN30SoF5zm
BVxT+7x4EitM3ZqcABLwbTyUhhjdHKjo3aF/TjX/cIqAnEFhzm663d60Z5jREipb
YX6BzsihzNoMYBbpSRQUlXaYxkQnUnjmWF8kHXDq8MI30w7Gp2+uIjZiH7Yr9rLl
KWjRkVdEcPTr1LfEG1AI82qFX2+0x/d7/FNlYlFiMYoYGzHbi2RJjBJs6wQMZdkX
o+l/tmZCz+rTrGro37N1+Yzw1cXrLL+Ko+WQoJq4shzEYeLMVoVrt1rvByru180B
um+ydDr6FGTrWxWuMqJBH/b6Qsw+MC5Ub53HYDrRjzKRFkUdUtupZlsH9UTlCYBP
qbEyWmUkUgnbZDfEHMxxoY5mQih9/qL1bAWOCD2c+FcOHLwyHZFtihahEkZ9eU43
Oujy3Pd9XnZNW0Kl8obbaFhMppKf6uWFQ8LQrrGrkyVOtk/+RwX2KYk5ykivMFsZ
rn13x/iO4HOOS3NZxVN80lfF05me0xmlpfT/RZA8JqURbKPQQkurm8esdlWL8rwJ
SK1GUe1hC5YmXbDhQdjCK8ZjCR52vENIIi1abEOROeGErpNMIPcSWsIQm4F/Djd4
Twx4OJQHb790HFfPovAICk5pReaFh4q4s/p5ELWnMm77pXcjwFiWx7DKm8pLuXEs
NlQC1BdJbMGV7NKrhe4kpR76G+IRVxdodz0reCIdotB17S9JRmR7qU21apkLGznX
LpjcRd8ho4MvHFANyprsZF5cefnOPqOR8LS3cNBIttbcZycqH4VPaNpBXZty9Moq
3XD/rNLVPtjreO7vr9913ZaAzb2YxK2zmo3AgMpaCv8/v8TAOI6nFOY0H92R7gLI
LFpvFaWSDQ8tUnc/Rb0cPifz0eB7YFqgpq9h/wuQu1XIpcGt4rwE3rx6dcHcJ315
GjXafO+Biqo10UM65chzChVbMdyCMbkFmiXTjgnTj6TLty8Sjqx7rV30ZUs8jSr9
nOadpmOZTcgQAVX0s35yOYEM+KNbhcDNqgE4L5cJ5KXFPAtn9xlqBAFqpnDDzXXV
Fx3qsUGZJwNAjRqC+2cgEkq9K/bEig4qbJ8dlqXtAasO88SwgQVmYSTsi7C5RSW4
H7n4+aSItVojOChY/lhoxsLn1kNKhz3H46FdIC87l4upJCyapAu0QmPptOBXzZQr
O2GvJf55UclS4Q7IGgu3ehh9WYbUckDn0UuB278kTZrNetvkIJTgO28uQLMBsgoW
b9CDdo58H58sQ6vILKT4jpbtgVDDUefcEgQnq31jxzhtVDzC29y7mOYXLWiI8bql
iJOyNBXKfUiEBNz3qeIcNrK2RhtD7An7dY4a1Be1o/6D+5VPVtv1KRG29JSWndMZ
AhoMieRwH1jILQmAy+2V/nSM/kvqVCeZY+L0Nl9v+H+UY6jBErjru7wOOuFojmrx
/JcnbqZBZlR3q1t1lEjvl77JSXLDDrdk9vDb5KV29+q9hBl8uwjtB08ZKatxBi4G
9oIjdOp3hKlC7Lx02kjja7JQCA3sxlSDG4EgVd6nh03Zbg9W5CVtYVF+nDht+MCD
0VWimhA/Ycfl8/ASPcQ952EV1Biy2vIBB73BsEDuxZLTPBtWq3LBVChHhL7NjPJT
pr1Pa9Sagx/qhTxCuJKGTmUjw/8oG19l1xg9NQHUdlSLdDo4mYjUGFxEMslQGXwH
CBxsUBwLcDaRWKr6jHPTSLGyg/TBRjVkuC0OCzNzI9/ChpLbQ2KV046XEKSSJ32u
8ZpVBgsheCyxJpiTUIC8UtWZRtxxilMcg9nbfRWTW9IHlR6rIIxFiM+l+F5cvVUc
nitpfQfrBHEj9ovhIy9HRep2IMe/YpjNfVDiY7A8Asn4H0FsLouEg2WLpjlaJBfy
KSznANGv6XhPOaKsEuCH1W3ismTUSfrZ0M2TIDXdQWC6b4Ni/Is/R5BiK4s8+urR
1dn/ibBqRyezhgkpHJj3mlaWVBofUEhQlv+eJY3I6jXsc8jplpGnce4lkdPK+DTN
mGcHwf7KnTHiPDb/SD0mxz8zjoBR27uehjvikfcfVByCgUCCeO4tpphD8k8dLp8O
engAiCxA2teWRplw665z29um3YQ6Ar6KM5JSF6mfvEYUf0L14sRUHI5iMItOk06+
Hi8TlmZZQfmw8va4Ne5rFQQvqGksVvleLHk6dfdXB3QCFOEaVy1cp/WmweUZoaEu
BMVRM1NMEYwsVxcJ4b732Jkdhj0Wtiku3bAbmK1G0Nk/rxbV/XiWwLglfpzBZ7T/
yNoLqEIyUFxVRbPiq8d7v3nYL6zFoDQ2evXui6JlBSUdt18I3fhFCDsp2MyTXmh/
NgLywkQO8u2YkwMKJMlPeyTOlWWaQF6ZzrUX0SIypQwqYtlWlfVLjrmdpINdzl3l
8ZiGdXu82+v7Zg8bIID4qEuPOdDRbxTXSxeI30etUS4fkx6i9TzRnRkVaiGAI6Wz
1sG9MaIZm34ecnWMfoUElC+D2hwI0C3Q8hvYrAA/4/nsSvx3o9Clh1yYqS+lk6sw
BpCfTELwo28A1RlqTKg8GxmrMY/InvGOISSL+YVVPuTrnjRhPiAWeY+uGuNTXoVk
Ah/fhr1SX3+ErowgZONgi0Ru/I/RVl5DVkdh67k0yyDSb9qlV8XYn5Ik8HMeETL7
gOzEIi6rXaqByh+cN72qjGfgReiMW3Su2Gm45R45ctdhWyrQwYn93/eoHzw+6WNY
a6ogjhPEykv7SzKem0ulxMx6uOLFORlvDiLmI7tlm0b2AORrpWk442VVx250HbBe
8H9la2rMz0YT5xI4N/JlRBvGoyHnpLBqaDocBDGRBIQQVQgiQpXWrFG4sV1DEOya
BxD0UMWr1xHOEV2wub3GgjVDo7RKcFc3fA2Q/Y1IVrrFo5PolMCWFvUWMXte/c/F
LV1LjngGA28cM9JNZDzTPlxOPzvba8+I4ZIOEt1/O3rHMTC8NyJ+VZwJktE2/7yD
CmfZDQII8e3i/kOy70liuLA53+vnCPfFgYi8MJiaO4IgBaAlkhUIvQvx5Sp6bHNT
Xjc4E3RhzXhGyQ6b7XCzxXm528yEUSy6VP2mCO6OHS0sLNNodH8vTbDPKoyrR7BB
jw8Li2O11bhBgxbWudmucdbIUsuYxsmtqLDvIRWGkr/TZtiXR1UulIqOV34UYUoL
a/70vuLh0NnhjYn+UwXSUnS0iN+N6x/PI/YATnSbjua/Iqn8HL0qBDq4lO9PcCHl
nR0YFxGoeHWh1HVynpMh2i4JjwvQ+tnZcXsYpx3mKu0xWjxgLhj8cdhRE1PfQvd0
3/gwaE7ebWYDMUzFaxdQcXd6FpZkFSBuiHlvD17vQN+WpDqPOxFL6pfwGGPPBMkn
4LXRbW7+mdTFeCMeK/fpsiGiL8crMjxKZ3EfvWpurhgMOBHRLqtgGBdXo2vFkUUK
+WmBnBXtCXOAru50eVGwDaW+EMjXLfUjt+xIZPfF5ezNXc2Hcwds2J2T9ohVzWzV
+DH7iZdgU+JTpY5dZKCB+vSFSp02ROdRdNHtHCCuWpMR42WBZ8szSFODOyD8oMuG
Ny1P5JSioUkkHqyynqJJYZyfJDjGElBWPNxBDt599LyQI2U4XEQ217W745F/SUEy
NqvS4BGuKHIUcRXTsf2m0REWNOTSyPMhE3ObfzW5WCd3g/ufrkicrlbh8By9sNGj
51+keGUwG1UCNKB8CJs50cCY3+KqI+inCfENJbP0+PPTDAP6/pj8A9k5VaAKsTPc
qTNWXJDdAMhJOKhGC/9am74URa3RjJQPfS67snA4HxA97+8WRGYglBkXg06c0gCX
dLmjnA0Bf1A6s9gH+eMSvbZ++vwS5GN/hpXGvJhvw5PS1IIZUNxj4KZt3ASbhB+V
UmDAQQliuJtczVT9/Ms22g==
`pragma protect end_protected
