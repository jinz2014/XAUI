// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QqqNEVpfKAt+g6Uk+FFlFmgR9+57H/UyoWKx010Ig2Dp+ho/L+3gV2iUg5F21z23
7jbnie0bY75wBir0nCQ7xb/pmfxJ8bvaSPGCIW7ClqPPGnS99869xYo33PAMULzr
k8yfoJ4oxLM3cb+6hXOQbkh9VXDhj0h1EE5rDyr505E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5712)
DZWM9i8iW8uk21DeqrOcfQ2my9a3TXsFESgtYvEPEpnnfN6M29jGWPR/fEqE3zFH
BrTNu3g+Lc2TThxAA6GP2zMh8p6g3+VZpM5KCmp+y+3kdROVGOPZ45b95bQ7GRBj
VmHHpPoneJgwDY92cyI0IqzUOuXD8BY/vv0OoSolbM4LJa7slx7FBIr7p0b6yLNk
/mdwbaP3ThyqWVX8tzdSYHz87RN13vi+P/bVI3ZtofEc7wVabRpYbOVQMJ7UWiu2
IkaqONN9yWz8mHXJPxYqTXotNah12NjthtcHfGZH9pNoisyfmqos2dOcaGmSqB4s
y6CP3IfwxDzCio5CgUC+yr9f0LCyiC63t6fx/Y3UlY7sji19QFxx2G+rzfR6Tf8/
t600pHy+ZYuiWaIbFCJsL2Sl8U2iYnXvw135aUI+PhhzVzykvL6UeVD9ff9LL7vb
bat0vmHA1cNT6umexzqA/GYbQ39QS5wFW2VJmdTF3laAIdfjpGprRk2fE1k9+3sz
6LgyDKfrJa2v993cjnAW1YrkWmg+iXvoACBwS+/bSFEznwGuzGuvkRmcCIDz1TM5
i09fZgaOyT6YAc2DwL5fpTvK5BLl69pdgnHmdlbHF1X/h5Co58QmmhzHRJbvDxBT
EO9Cji5HOql5xRCphFYEMvcUvTJY31zLypwtotQjLHZLGJko9pdtHWncwT6tzLkH
K0i57Z/GRlZqimLYkH7i/0NimtEbNDQeK1jCfzH0NHt1aqvhyr3MbQ5jf6F5Ujpf
1RDBDqr+mdr+TlQ6Js7UjudWj2GRvBigVJKl0Z0BV/wuKDgNGYeUexdi9F58ExSC
q/RC5t/Shz6j2O4otCClLiGaco+uK8mfvc0VoX6jdCsdNM5xWZu5dUDjwZIz3Ub8
rNI7iJkGpFeN3nI7MeV0RK7B7P7uO4bD/DU9v+jQ9Ni3R5nZq3nzJGEhsX9MpdM2
BOnr5EfZwoQDtHgp34b14BgkiN4aFwLcVFQDmGVQPQhEmgSB9FDbz1BbbZN/MHy5
IoVJHIDoIvehOvIeNNbe1lXJ4EiCfBonu4iby82xRbTfjGovHehTqQDHzQ8tpgM2
a9undeGiNjwY+87YPJVKHj/odng8p5WX9VFCW18bbxLLIUwjz5/389j7sldHMdoH
aSEgRpidSzM2UopnMjeN3LXogThxJJhl9hwJFAuXU0Th7NANSaOmAolSYZqa7sjE
Bvr5bkvtron+46cmBtf5F+WeKsLXJmP4aZfgL2kLdf5RoMiCt9GEBALEYo86rIP3
xRP2ROqq6oH0RTx5dLSsoK0Wu4kvZE2avaVzE/q7jHxvXoEO71GyerNbGqZ5qg1d
YAlcwygK2TzRgMtb8sXfOBl+a6VrvDt+vfxw7pttBe3ES/3cJ0LI6dnlfnnNLYP3
GsaV/3zyEJzSLNqLhtcO9YcS01lQC/TULuKkG478rC2d6zAy/WTHyqz5Y0K47zY2
YmDEhkoShDitHU26DhhsY+yTVmviR8O46PnF6Nday8ChYsHlykwIybkjLrxIJsiK
Z7an9mtZhxEOKg5IzI9oNxZfSCrfI/3JZjAmsgbHH49DzRicyNVSEpoUVyqD+Xxl
FGIXetuQv6Dm7dBTAeZuyrWqq9TAGkGp8dq+CpG4qLzlL0xg15mH3U68fKPsUjpW
LWWjnLH0R1OQ7gHXqGSJXB03m0hYtcIkuYlbeEkpvqxtVqWn2HUsLIQogsukP8Cy
yPnMaplLqxYluGwhS8SJANFUuJGfRUPEsFZmkHrkZF59empORBPQt4kXpoCqzALz
uYnmd+SKos7CZamtmHQYJuYj2DhIFgddWuIg999woeZGCnrm91h1cLKoHJ2T1fr5
EN8NzUsy53KSVKItWErbqTZhG8StQGo5r7trv5pRrmIrKpomGGNYjKUuDpDRBapj
dL8G0ZMXGSWrOzOb3pcFWFdWCRRoaJYzvVXo/F1o3JxiwOIbURfr0ytOV0+RMTdH
ZaajhtBBhHFE3xQYzxFDlRprEyL0T2sdQBv8B1EQyvHqbG46KerHxDzI77CfhDOl
dwR78BTWlPPE9i6b6JeiUVzwy29CnJVc98/+Cr/iRr0zbmXRqHQZc1ypqG5ZX0il
AdatIIedBwRJDMr41Ajo7UELyf7WXz+7DgA3bR0sp0xW924M26/4eEJCqMEI2Ia+
Yy+lnAdAR+6fNw2LVx5GyPWXDYe2WC1Hq0NC2s1QbU1ildlb2S2DzdSrTPYfmX9z
cIreD5fDSx1F1U01GIRxYZiSCno9r1GaEl/5hIR+PeKZeY54nDEu7CPDurcFL/zk
TBo09Ih16Q1mpXD3bFWhrlbQsWZ7QN2Onm23fShf4bc14CVrnRNAwp/YBXUNQDYn
R8k1QmATrJmNhhn3R7S8GxgdNgJ00iiv61SPNCqV7Nd/TDLtxPNrOkkVROYNLHie
uLaCY3BqJQ4f57HfM+KBZMPqBDRLTh0VjJZ6UZIX9UtHSUaPLvxO9Ek5nS1iDb1P
g+C5kqGA6sZxLYfxDjrn2QiabEYjW5fFS1hJXovjbW6U+MUNWeomoRkWtsGPqluu
GXMDrO8DCFOD6WH7Fby1/vZanr1VoIcnmVujWUmqCu5rwTSajdtGbOejlD6cv7IE
l3ZdvaaWkgxEdGfnCCjLQdcmt7eTt8HyYvub335MPxJLHlmHJCYFMz5md/d1J+d9
W6MCjsIqc2ctO5xRImAfN48oRtpNo88OiJQc44Awz94wKZuG/2DM/+oxhLxry5fW
mHaaLX/XHRyAmzTZo2O7G/PeppUhf09zm28AHzKljrnVShdT6jQ1YJxqzy3YtOKf
ByTDBrmoSwdrmY25pvwS6CEVwVFyIxoDSIj78YyP26vBq0kpcK1TRMKMZxqjh7Us
bPPUI3TVzfuNmPdRhWWf02R2S7xSrp9m5USetMANQDHpSkPHpJzRb9XkhJTUjof9
haSNIfl5H429Raz/foGPYdSW740nfvVJmCu2uAJSMBfRqRBsa4KoGKUWDQTac109
7T7oo03V2sSo4OOFj6TOtnXGMhetKpxhzkH6Bn36HNMr8n6Ey80+9jmIz6dgEqnx
kxUYuF29OK6SB/S549yecQKvtrusPp9qY9z6/IZ0sxyCPfCjV37v25F4543QXW3V
l/1Ta3I1WVAU2O8SudoFivQUE59+tjNtJWg2CTB9WYciNTgKfwGH1AKK6YIiKZw2
8MZTGj9CM6egottPaoMIHONhkPJrs0ptCrqzPpZg7PMBSOofXkKhgNfSKBT/gJ70
2Xq7uh9vuHsmRWg64w1ZfUx7dswgY0Y+q/Yi72iHCSMxEByQxTTR0E2M5syPQ1M1
YRYXSTlbBR37E6ZhkKUOHAIw2c+Ne2fEV3z9AXWSTyF9hvaFdJe/NNrdXadsbhFq
rGNDlXJAlBVmzHFf7LtE77L9GPjct3ExjsA/mdOT9rwKm3TfeoyZM0mr4sSxwzNZ
T/YeDSfs0hEVKAbVuGYckN5Pus0n3WToXn8U5bNrdIwz/H+Vwt8EhQaAYDl5sGo8
pJQ3fLlhv2wpg6PaZPNgT7fwkoNnZ5B/yfjCkFsS+mlsFxGfgEtynESFS5OV+11o
Yes+azSg9Aj5MAB7GE7dm2wmJKbn2P7EFQ3mHcRoet9A7jAYx7wT52m/5CJCe12p
Fl+VIA6ctbH5ctTvNdsZE1cugBD6rIUDLs0r7v7vdrHWeyNB5fafFarMK9i4+Dl7
z9P6OkAJL+MWLlBNUaTa1z4w0uyZ7f88D2Rmmt+p3bCLwj+kl2u/DZShchw08i7+
hcggfVBK/9SZJG6vpVInLrGsuauyqXfcA/iDZhEahl8fG286xTYd8kbbP5esd29s
1GonyB88KG8zqEU2/LsNMwgD1VIHttbjk+j7IUDnrpR7J2Tel7PCoOdwgcCJLsl4
u9torIr2F8OPM9daBNpOszXDOQ9IkGv5sns9e5hZARKuMXClPpn6Zrs010KoPsyq
7SnUj8ts7aqsHcv5V4qPsnBgcEVI1ZgtQj8GeYgaAhLcRqUBDMIKaiNdrdg3Li/o
K3YMB6QpVTfWbiW7rUlGtVIWXp++S68zrI1m2gAdEYN4Nm7/MG3Fsi/9auaNtVye
nvEVh4p5OzaYyWy04dVAmTCFE5i0lB1sjPV1XFHp1tkYCxvsAWDhVlsFT3L8vMLp
It6LfaVY2/7execE8/0sz2S+8d2L8Mo5bEXYaxwg9aSgnst/ahY8DorajPnE+8t4
KWR7cYGCXMoBoEOdtGbMo74N8FOf0nHXCIN+oAMgYWrF5imekd83X7kLCLuStARA
bzS+QHeE0lbS66ydIb3QIljnNGYC5Iaebh52F1ceLgwYMiBZMoMj6KUL7F7JUIIN
PW1mwKZFCSKyvx8N46gsFxyI26lZsfe1bWfzPQZqvn8BAEzSwVRe9osvYkxlGksC
uIthx3P+ypcllGSNxX0+N8NE/4f2kTjkSHPk/jBeexcC9W+mtiYPEeZdWK5CUM8K
gXavMexJ5QH/xPrdmlMFyOb89t3lWL9MHVfQ7OBHixLy0JndhrODHGyg8iptdEMq
A0wHBKJFgifBQiY7PLgfPWIXwD5MAfOcJzmROfSSGvnbN41WGIaa15ElA6I8MeCo
9admqyVihB9TDcFEF4zcM9A/brMinxgZ7G7zXgp4JEq+VdZ2BnQnz1XQeUDfw2qu
4ce24+Be77V7IQVvqfprB5VXuj9cX3FoU3F7VdvCKdNEByIDnLX9J7/w1xix8Tjo
lasa22LXtFZvvPEA6NXijdBbrGzzbD14Mt4yUZjeLgJ2Qq9Oj4pNbYy+vUdVeT1u
fkO2QmHzKmMNxt9lNoxNRZbaqoGsEx6aHkXX7ch8ABgZ1r/M2oZsrVFy8hStX6lQ
rbJs97U9u/KXb4LXIAXpkHOG4kAN/765YuDmsuqwH6OjN4BCWOITKOiZtMi0jHTk
pzVRZqLG6JpnBssPFt+tPZWfEcdOYFxBXokFeIqLzSnAwoU8yXqn/sSxd50c+8Yb
+wJNV72QX/LPNYqUYuOhJQh0qnIkClBHPJrTKVLtjhvHp0l9hMFvIPsSA5bCPPaH
KFrsFk9H9Ay+LWNOvoob+ilJHzmXslQKQ+1n58G/INYzoupNFPANxVS4nqFGo9U2
5F1h8Sn+ykes9KdXjSIbA0XnJ7VlP6OsRfnGYVD2DylA4Id9annT5TkbEvnaNo+5
nUtw7hODvl5vZCYVJK7/gWYqca/mI7z3sHGq5cPudL6TAOlq04OlWcIirCLmYvtb
Zs8ybq1csiY9P0nlTPOAdx9TqKsNEj3pEgOR3+H812Q8qAvW3MWNZ/xH1ZygUy+T
4uAiwZmtRb8nD8y7FgEWKwHM3pvPil4PPYGEfrjMSQZ2xYIMVE9ulR44uCsQgN0f
YMV5+pCb/21h99psilLIXSP2227HxZBwV+L8HTaE5AC0QLMtwYyiFKQgBF11CXta
vWTe8fxxtbE2GHrQz7rqfIk15dIAAW8w+OST3nP23veLlx2+iaBaYMOQea4IUEBB
n2azn/Q7bAMxefe3UOERhGf691qG94AaBAt+ZbvKT6/3ZWf+xoZeY+EXsh7Ymg0n
HsEnjwwRX0+oiCWLzmyFTzh9XQKr200rI9a5GEmHTYmUvVaRXffYhg+dz21uzEFk
pgEYm6kVJWGY+p40uV/N/0FDH983bt8B8P9FCaOw0XVjyfS8WqMgM7I3mGIIwJvM
/T59d4ZjcuT9wlL6ZeAYgyeZpdkS99fhypmC/9vB3a6c9QM9otrKXLhoTPhi+Y5x
KpETRttF/tCx6KNiH/SjRp9aa6dyvI6eHPsRRG3xpaAMuJ1AVeZBrhDweLLHKUZ/
0n5/FCbBGsxUZlIQKyzTIrflgRjYBAfLiqgNxoQG5oYf2sv43EvjXTNVL55kHTaD
35FGrfivTjfBS1s4kkaFYlTKVAuScGXRYYHcwpET6XRkY1M6tvAyhPtFdTH+QAe7
9nyoA2LYweAZjtQCtKcTINLBpJMVKpAmXD4GZWvhtG70L5L6/dckUI+pFFOpMpfy
ZOSAAt4E+pNQxVJCFGqoZ+GGlEYcDc6SslMLgdwtDDT1PrU8W21EBxiowmAopR7w
OAkra21Y/CLqAWnfyEa2anauKRH/ke9TyizbYoC4VkyHsX0trjmEjmHa7CSWdWoX
SnqhGudzvNj5mSeFoDHvbWWy4lpz9QA3xVg1/rP9I5kWn9KLSw+E5+CB64YsOklo
R7ZiM6Vw4hph0OdipPYGlzPkUsPAYn7W4nxoIkd6+epz4aC6HlhtkbSrT8Mg8WF5
0oOyXh+tEnPiaLYve/U/Ta3JrVrIwNrGVS5DxK3oW5v8PeeFKl2U1seR0U62iNHZ
L8sSxdVsDPycZYTqgiIY7+WbXZLVJNhhw14gS/BABMCY/zYgbj5rg+mVY/uoJI/j
PUyCtNHRD2dOMbXoEzXziwiIZe+pKb555DKQbX5z3GguNJ5oitLHxLMA7GMXlvcx
sHuSMZ/1U9wQ3A0fU7F/NiI35LluKyEhrXDE48TbZeR///75WDoStvApk5K1svKn
HfuGTUZHBSY74dLdJ55hJIyc67Xl402syI14MycW2hbFMqGesdkdRuFcNzMoLXtq
z96XRNofUbzT2EpOdesa9wp7wM370eXTTvAXtn/fJR/wLgpIi5Ot5NVF+JaZlV4J
asLxfqf6PM0K+gjOpYHNyE43AVWzlhc7+aLn/lEnpP8S3M91I/EOd9NBnOaabqM2
dhd/y69Qk7QQc3i4odRmjfNXb6yhzkkrTvjIb+TCC9I8v8IAF2EIlkm6jVbJys2+
kH1gXaFKj4AQmN6joqVBms+MglgKLQcnV+sUxMrIu2RO8Xlt8bYLk52Qo7V2Zrdk
+IqR+6w+Jz+WB9lJ5yupYe/RTeWCxn4/fQ+IqXdpW8z/FMAdjR5af9GscLQECyFg
hjHGksXwbt/JFusg/u07DV3pvBtUkMEg4y/ZNrBuJHVYfQfl7dtMzJ0c00DctkDR
3Tq+Dnv8v9zF3Qev9t7wRLemJmzwGtWd6JRqNUbuV00LNy/tVf4at7azNw1YqhKf
nHczNyo4eStYmPnHlQMbF8bqqsPqvRFM7XirO/JtqF3qJbzaAnOkpcPJw9o+aGbT
5KPm8i2OtO9nJwgE+9fwtJz0CbzwM/Zkh/WiB9bUyvL3wMFCkwwcbX7H652xYnJE
60yGwgOAFlVJT+AW6LJ13AGHNxwTcChm+r6fyGnhkb1nc1ZqlbDUZ1JwHY2QA7Pc
D870Uq8lGhs9AaC+iwneul6RwClYRCCZgx3scF7Tju0+Q12HhwUkH+B7By7XMbYh
RaBPA6VqIsrfP9/gbvrZXzmOFxDrLY/TRrsxCFxNidzPdiYKwh5aW12HkDWF7lW5
XGJhVt9Iu56VZok97qxUSBh+3y4BEf3vUqg35HKZ4IEJl78G3SoDjuitQPMic91m
2RxAnjt6nPrUvYIvUcsuASo3ToXnDo79kMDB8RAbgTKf4mlLY0ta/4/6kO4hWxPc
q8YtrNhWmDSe717PtE3FMXuaK5eb2s3eCi78o+UwbPa2oA6zq5IWdHWctFWePBr5
gDOKfQJ4fIx1ex5Mx8E+ZU6V3L1BFAXtS5mZNtNhy0RVBhrk7Ubqo1ID9hDn4uZs
`pragma protect end_protected
