// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mvDxhy76dzL7xhUZZn8ilNFsclU+wXJpYgaoAeiza434Z1U5itmviqICkrEVlGu5
VfOCkLCCrlFWYL4A0oXiQYKE2Dg37PwOVD+r4jNy0K2C080so91kNRR2nT7XyaKO
SSgPsjk/pOdgzhftfxn0lz+r4knUU+UX4q9k7OU5pIU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10848)
ig7tl0+XavOz/4qYtUDOs22jMXLuSE/PQqyh7Hbq/DHJfONWF2N9FO0Z3eDoBup8
jSEqJuxKcVtUzoTr4xDrPovzbFgCSxxs3v1HIo4h/tUzX/c/6D4q2wLEXKcdgP6H
ry7xOXfWfb1Y1nbahhrVgCAIC4VLra7+62nP33uTb/j3FjEwNSMU/swsDPo2jn/9
1eNkJ3wRf1ebFbWoXVm2FiyQEKkvGNUptBgjKq0NK1pNp3cI/AsKOwnKp0nAyhrV
2p/xAg+yFx0HLFYpvyYGEN3/X4+LeGbZh3BvcYFRqIlaTrsE5wmOcZ9ipisCZ/kI
yG95f704atMhZLAcMKcJeZQhRgFSlmaa4Vvw9EuBttMgFWPkfb/DzG5ZRlmfnBnB
ADBQbLxxHge+RB08E/eHD+Li4AeR/95eVwHi1iKyfJH7zhLDaixwg8wKCHBkekfA
7aegTlmi49h1Mhnn3cZQ4TQqDjcMz/1E73thIem0x8OK2xWJT1snDp4GDpy+BeDX
xNcGR2VGcDiIurypMGTBMuQ7MjDI10WAW6TtwgUnx9aMwBDFTDrC3d884i2M95+C
WUX+dbbnsRZCcqzD/oygsZVnEUguT+ZPVcBuGSJkQ+vMIEnyVxpCyGrhDdt5uR1d
r5JLRwFwWiaMJwVZwbTsX3S73R2K04yXLjQ/wGpAOe6FR7I0lTrCFcErjrk6xjFu
fySVNupXOhY+IjqFzwxQj0VJ+kFgUpvabhuiJbK9G3jJSLLvgY2WEnInqcPeUqVo
Tx+T7uqjq5JGFx6yVEgYnEt9qaeSvPk/TdmDpGIIrKsDvbcKw4iwbnccahaum8GZ
qSn9qoy+tV0+tmBnV4RKf5SewU8V1afPZsB/YZHaQnHXNYqK+q8bhu+HqHhZJHG7
RrHEVVAX672EWv01lYXFHkjSACJvKUg8c0TublYBKdvV8RlC7juGvDatIMXIJAEJ
8FMd07gQhGh8Ifxp/yKe2RM5rlBdSrb2xbSpNcyGpZTlhYqOGtzC3tIAIkKk9e/7
w6Yu6qJkjEYmEdht9+BtCvyLcw9vAZafcvQw7PzbbI8c8q5BmUY7Vzws7vX1OS22
FSagmVmQFSecOyUI5RoS+70NAkJAEvm/OjMetI4VYIGNOd/JqMoNq+tAR98mdad5
iWytDGEJJgisMObFsk6Nu5JdxDme+12cAVE4jC7tu/hb6tj+vJmW9CDeAhcA0MAc
ofbvK0xUeJBWZTxwblCFEdKXp7xETXloBNFfpHlGadg8TbkTy6v4k48gXtg4wE6q
/4kaMt6mG/OIEhBoUVr4GH9WdjsewR6PO3w0RiicK8KzPFc3MdHoSE4qNYtkQCjI
rxqyhT2pZfFUvX2uPLiXd6G1P80vOTWiaJ66ToxLMW4CVgn6IRIW2AkYZIsNHNds
lxbAmRB0SCPfz+nE1Dqw2GtIzPk+OLjRCAgEUM+3LmMQ0B9d5fuduMDJZoO4PhBB
m58tn7Jl7xnI8QFjF0n3cmyOaMSfjMNpZXxYdJ5vlyh+uqsm8tAhHrELJu5zt2Kw
7XCIN7zWfEvaK8EIjmkf9QmqlS+DtVExL0B/Ijc/BluRnArxTxhSmhMJAo7/9Tli
eT1bh6HJC2ljNQAotX/5guOo/DvfzMG1LlcAcYkS9Z3jmzidpN8fLZarWZwPnY1k
zSNgSi24ZSdiqV1+MLDeBSn/WfJXt/P0SgQgp0KlwUEJQ7g2aPEpCbUFhtwXlWa8
drovc/HDmf+JjzMf5hsW5vzMomCtuk1VTLbZhxk0OpKdFdEUUn9uwfEiVmp1+rBY
NYN31B98140Ak0YThnM5hE1tc3kfU28DsWZCjVGdHdKR/91ZZOHGDoo6ruHDHw3T
IsLB69fh/TkcgUevXe2oAEqqbXs4ZoJLnv+QrLtKqS7fBej9OjK82ef4Ks6YPkOD
AaVTvGDF5lT5gJxOPHppaQgTBcG6cyAKgq05ljG/+3vaLJ6W4v10OoBhK6JFE90/
/UzB3ukGKIbxMAdospCmRiRsGPh18bWAQauJMPit38i9UbxAULkGYVGMl7SFg4t+
F2RdEPa3rEERn/R2ObSVLYOU+OGuNW1BEzv65VJ/LQI7sm+YDWbTlAdgN77PjqRp
+FnfcpcQ8iDx9k2RpbSTuzas0JeNuUTAZtG18lmGDsDvP3Qk8555vfO9OVlyLmdS
8sq+7FfhTxnHLCLzyuJ4priDBYy/P55frMEYi7Zw1B+7gKbLjkRv9BoXFeAWQqFt
u1CK2Ti8Q0+/d6Hu0Ze1MILUTcHuhYzCfjLAgXC6kG74qDj/7gyG6oSoyo4SqUUz
WwI7BUiQab/DAcBkeTto6bZyyiXfngebpIHUmYx3AC54oaAhIwLTbeYO/NxsakiZ
Hnc7RtBdVe3oi4tur2JuTjCf7pytJCtXTfJdojZOhJLhy6ajniymmMO5qQlSMb6G
gxt+9E3AZN3R6mAg+8Jfsk67G1DBjyBeC4irVUMi9IqtuZ7alFtJZg2HnaVDCe1D
g8Uw5IprNdRRIDc/Uq396oa6OEJfIVIsvmK0MfK2KahNKQckRGxSYrJEiwV/XKM0
d1qxoAqtmhJQG4nZ+42bi9wd4cPQ5q5ibI5xAzNywLMeG1Kv9Z9LmSi/fSYuwcLT
tAwhQnuw50Os/GeFmiq/CYFuEOwZsrtUZe5pNULLeQo7POYXMI+3RyIfZxpRhGi/
exc4ZYYuSirP+lVB4Pvs8YkF3s+RTCKygixlo/Rk/QdpVj8Fm6VDL4cHjoEsNJRA
SowMxg5nT9MqWytnd2/FgBI7kNlN5fwMEFskHOl77i8INIREq1JpNdLHCM99pyxk
DJRZuPgD3Hy8HzyRvEjQ9h3T9mEhpemC25daWdCBB4i12S2dFEUE7riNff34HEGM
UqJKlTEnVMN26H8Mi7U3pJcofz6WMhiNDfMuaizlme1Q2hk99s3Nj5BaSjiS3pI/
rxwZr8daNMIFBIxM/o6md6M1n90eqxNR/GwSclDLOUCZBVn/7fGyP0hAP0+/FGdw
mUo3b3GXLQFneBSoswsgnhl20AH2Dq7MiV/UdBrNbLnigDHvpkAyDCMa8gl0Z9Fz
8EoVhnojv6LxcetfAoHMUJJ+iMoNAW6+FRAUytTxQFISiv/zSX2dG8YwKWuSdwY7
c7VPoUIRJmWAnjWE+lNLKDnRDke+GR0sDT1R80YhEy3IWSqhCzB2IP02QLT8AXhb
6l+TVEVlukUJclgb48wQAXWopXQsKTnZ5wOh7KFGIYZtZaKukr3Nc/2HpzS3ZrKm
riZ6Mn+/f3a+JEumitkf0H6ieAvJm7xJIvBaIq/39z2KwChIrXnVtzTFgxKP+VkA
BGZad+egEwKFEHwwCfO3q1u7WFiVLpFaBTc/eaA2PiwDqSovjz+k35fiAqBLb+mx
dkgX7HI4kUO9KWZ64BTlJyKBnA/ujfvJDRlfXLYchtMwQNCt4LeXc2qTsY4W9lGw
uZnJyvJG1LK8c0dqh4dNo3s0TLsZ8FTM18b3OmscNfcZk3UspGNREOEf2MltNRK1
jxrq1ICgH9KuR7Y0GomINnWUlGSkHjhZduDwYPk59ondj/87IpC7DnKZZCqjoHBZ
QZslWU+HlgUZn5eRwCziEo8If/ZHUjQ/AXT5oX1ymrfifad4NBmokYz52NEugNe5
dsT/zK7ugBuvMZvyd/tAKuD/OvSddN4jKoRuDm0cF8SeHHMNBXIBUnPOr10+cLQB
MtJL47Xx1oYuBhawbXUQgHCeBErnNZJC82DExLQhLxdc76+6Zx7p9uwdTLi94onS
YGe9fQSpF/Azg8RfbKBT8PFV52yr+29wpHO77fJac599gjzxQZfpz7Hb8sQllv3y
1rhNwq8tXNfcjFrxpv5HniMxL7gJWptoxKmBmjiamPvG+eKTrNZcfkkAC6mgUgnb
tADg2ozIrSROnvAoUEiHXTE9tpVT757pbNh6t3+sFMvYMNepLqb67PdL96S1sNMB
Zc+sk0w7IYvozhVqFLFEkpgywnBJc+gOH1Rz1SHThy+PLIzhX07kfdc32TXsbYEO
QEQcI5f1REsh8CADDyqFZ1ysWHraUAD5U6BpkL9ZFARYxVrEjWG4mg1wJD98/iPK
oN16DCvQNS7KNWOacE831+DQXMv4mqMH2LHNtrcQao2TUN3QMTAaus8cUJH8+Ztr
7RqJCCf8gStTu+iMOdghrexxFT601Dwoc1kRHyVDEnk/qUMyHcBLi+eGh/femkUK
s/v9JssYeAnw7QndMfHX+7ZCTVX3q/15IwvR4lwJ7dFY97qZgurU5+4vO5TgJgYK
RKk/aN/K1SYoHz8tdTwJpKIuSpYisbD3CQMruuSn3KbvptWXiuvTu2kkUMsASFSd
cVLij0qQd5Gq0qy6qbd3PoK4y5NVnOekpoGTY4lvNWSvSzkqe2YAlMpqv+mMHwCm
r0fdKdULYLAGvqcJJW/ABuz7BJXEH6jYP5zjRAwz8qXb2vAjVE4G6KZedJQrps+y
p/+0jFlf+05CTi3YA02rtaB4Cq6sHdjzv+T93EaEPPU+86lnLi8d1NPnaP+ZlRBq
1rkkRuWqduHSR3rvjCdu5Yv14LkOMBaqTc7YIvCy3HMysYhQ0HFjsqSn0i3paNrF
6E+0TR4KuXaCOUCXaj+O05kHaBbI5HuqWBQ4Ux2AICCdKR4/UrU+x5+9bd6o7t5I
Ooqcm/tQAbmt09URO1AS9ouBXAoYhm10Jlj1XgXjf8m56OfPtPs+ghRhIxstbBqn
h9X0ufoqL2Khm2CAt394Dd/wd0UuBT2/1cIwtj3wBQkYXZ6kurPsqhrtp0jrKHL/
wREhG+VSLwqZx+iOuGFjCWUJqR0FZytKOTQflLsfTK7rEjzKFM8d0dGFRIpAwshF
VtdEKUNfH8hap6z1fO2FS7Tfq+XSRGQQkjpUNf6t8KSVoYRmP3DDFc08c30X1Dip
0swO22YMyVB0ksBlruXpXHrS03s/LYT3Mz9LkqSKDNU/u2xMq7maKT3WWDYIFhWi
qWMB/YE9y4xrvRKUNJklQEXoSoKcwz1kgj8/gr4t6mp3ArfDDvhC7EdPD3JF0Ac0
NuO1o0fmtzwZ8c2xo/qeIapjfbUqLPeMWgROV2TIQR/uz+RQICcJO2RLiBivfRVL
ZzJ2jbuQ0dw+QlBocazzCWs9yYm/sylH1EeCvPHv3DyY9eqR7Yns30YDFgYS0+xG
asCZCvFhJfyXlAIqTxZGuc3cTBTKHliTBroN394nGp/dP9kyMQKGkXgqx6qgvP+W
7Jz6Kcv7HvTpTmoBkb5XHE9osq2Af7pwqMCh6s++Qpp7Zprn0/p4grXTmwzh0hWH
lElfxEplOBGAy2F37uyxQ+0p6VjETmeKnwmCB9jdaDXKSHrMuFzPdDV6SazvH8Tj
Ko4jNlqGmJtGb1wuQpjrUVhsgFZo+z5vR6jw1Ez4eydKuKXOS44r0ycAbs8UFiL3
SgMQTjOIzdE7JCST9hCrtzytyuNeKKe0GNlZbvPRNWl8S5MTo9j7+CeczvNRBjlV
XupzWH2d1zLQe0bc3zmBQd1zAGVC/W+vawaQ2p5+z03JSG5PsGXtYm2mg130ZcAy
Lq5PTzar6XV+68hSQnEChnEooOeYEfB0eYRCwerZx9WNHaYC2I6Cm2gq0E+K5+zf
RvINCPqKFyhaLThgeXTW86LlFnkOgjOgMvWx2GxeWHRdLCs0Ha8LFWxF8HtOK6Ll
N3xRx5iKmWS+VFh3HGP0qek/j2oMJEPoDjb6gcZv0NGJgJ+g8rb2o0c2Rf6yn+Ge
o5GzPd/ISqlsqrbduwusYlESILybu4jYEpfHfAnKGCxPFKT/KW91PA1f7TWOvJ99
pJJsYnxH12INq7NpnTof5jMwpy9U8du7cc/heqop66DXY5aaV/Vo6gYumWmSQrRn
J9WbtIhbqoL9xJ2EYkH5Cszku63fmcpPl1P2O2Mm98sZ3WS9Xs7vwzGoznZRfldJ
EH4OpKwKTwXXOWxDdSS87ofaIvjxqrx+rb00PIA4GD9oZKnoF2CY9/IQjiYOy66W
KL3Wia++1mk4w+ad5Vb4S4DneCpKS8Zb+aDBFhTIrcXLldVdA4d3IbnqO7v7LpJ7
p4f6dGkIa4kX4sYOTh/OXrcjH8PK35p2xrfNoFT5saPiBMlN265tK6Wq2d8yGUjy
inmcTPF9WcJXpY7Cj+uHFAUX2oaondTrNXVR5rhYNe2I7dvOsc1Lu+7SK6CGWMaj
WGWlFQsoPn9mNvRSvxdxwRMjKMnRjmehfni/J2EYfuVEdhTP+ixKZ0l7jJLfCkay
Ec/oLJBEgc+fsex9OfuBCBIVyh2qsbtsw7vVmYhYJqelsPkAwxOL/AyC1uoVlHPm
DBqgCxJB0lBV2vz+QocUEH+EIAr3le5SDIEIMWvjptvB/26iqek6mb9sba2x7Ly4
sOqphzfzjhbnWV7BieAZLmJLnp8gfWxY2obwTmX3mHNcQZhtvgUV/Z4eEJ6Ykyrf
Md2+RbGOlbctz0W4R6MOLVdlLgznPYmzGFUYA3dI/OMXBQ0hXsDYm2qdvuN+WZ5f
c/9uaLP/7Oxe24hcO3Ay+jTKUZr0brbLMONOVTafY5MJBM4thZiA7zxbTV7i131w
wkG5ZD7GWFol+EDIU8BfjwrzjKDkMS+HtroLhlYk2Nh/xI0+6os1xo6SxotwasKF
hdl8GlZYJaIQquepo/uB7VQdTd7v5TAHbOCxfI2tHhUXt+NkX1HyVaGVo47Bw4w3
BSC9oLgUc2uo6ThX7ozYbIBJJFW7sBjAKyKZR8/QXXVGI/XodVxGTovnHSlTGMsW
RZdIMqGFQGqlpVrtz4e2LlMHBv1fmkrlTM4A/XlvmFfJn6bwyUUdQC/AxGAUlv26
qWPk4bc5rM/vELZrIm629pt3T5pfZehPS4nOFLZTX0NTx2HWy1Z/1Sh/3CeOICiC
UWEnoTvxpAim9EbRwGTtpJzYBZP055SjJCEmE/O0vvDXyrWolGHL6+a7CAPfnZYk
ypSy0z/n7mdcwmXxYdLa1wubM8CQp2kmPBgURh61L1uf28fi+7cgTKCdku1cA3wD
PIQfsNwhhIv7Z9+gGJOr6v5HLEMvWfmICxHqkYiTLrcyBwvtoNmFGrKfNrNB5ABY
rg5CxdD4DA7dF/+Y3aTE9ku8XUfKMsgHuoJjie2zbHudNX7TOi4WAU/dMrXr91ag
ieLSwjq4Grmh7QLY5mu6BRN3SBzPgAD1OMFcrpjTHC8NIJPGxc9HuSYiVgOIBYHB
wApHkJtm/LC0BETFx2WDC0ROU5V7dWNP4Enl2MenZNY0pabVI+4WRrioZ3FJeUgY
GCyTaKQnpPn7R3tlMm8z3bpvhKz/yZ2DuBaNLBKi4u8Vh2EtmIUDr4ZHP+GEtLvt
BmtIF+tmDk0xPInDCDntREU/CHlr8dDuoKiR8GVJTB7J6oHsEPqpEzXSTCd8joXh
3sxFE319r7E5gnU8lSiridsdyfmuEADQdBujClEHhjTHVrFVMzID/zOLBgJy/eb3
cWNBNaILR0L6fboiZYV0ovmWetq63cdFDlEHZK74EJp7nHybC5E98+VKFUzcSxL5
MpCfLF3Ojl5hbQCBDSAhN1Ped3dZs9UaizlV97ZuRAGjWlhsRrFrxAg6xcXQ5AV8
XnxGe9+D1vc7SOtzbNn5F16hy2h19cDMsXLR8AzoTv0AmAcrIByP+rAuoX8USYaQ
pCVsy7xKcoYiH9na2tmG6ECkfO2e017uuPoVOsyy83GH/5XvQCUpmZYlhhH15ktp
+yQ+nrqszLv/4ISKrBKx66bI5AxlDaMroxx+Sbim4jh6crFow+ECqIPaCdvS9YFV
YEuJWW01O2dSymTY09HFwj8UifLXLInt/Fz+Vbw7zLUL3uVWKf4w2C4mavdHRiz5
cyb64XYpJGpc5nfRQ4iCiFr6tRY6T9FLSyEc9N45w5GoGGk9WptZGaNi3m5MzePl
6oEItRPUd8YX2pEbsnG3vW3Ktorlw8JutPFAARrYiW0+HEWZFZzBiLXrsWgJTvkk
vGBUah0eBjYeUXB2Zam7B1mLBRExtqtY43SIZfJomVQfcidJUFquAfGVQaW14XUV
Dv8Z8JF02vFaccumiWmZ8vjw8Gt2mvoV/K0SMe4nHYTVaH1E7J5GhVk6LX1QtYOT
ls9tlxuhcoixzEu2con8TbLRm/Saq/3YUnKJs5OAgsR6AKFe8qvW+SdqzkFLf1km
o0LPCv378f0+1ZsnV/s1mV/BQiriBJoEF7bWMZtZWAq+40AZiP7vvLnFcyTkCnlM
ToBXpnMoYvTh+wUnLJk/Cg0isdAqKJuYcMBdadQDWoPjBBVFnLqSqvs9+IW4TbeW
3oDLmlLhg5b6oUQlto1VYomCfqxOGbmOKwIrYkNpkspgpfQf+gxkY9fFjkRz1Ks0
wxnCVecmA5TkmCWoARa88h2NVBpruAYeUvcEXk1gc7AfeYyXD6DG9a53KodraSo5
7kWtuS9RPY7pDaHLPKoBSgY6gwk+4tj7ZU/9XwFjVQ8SXjT09Tbn3rDS5/obSP9n
KYAZzMEoqtn5jwQ6M1baj5JTmkcsUTjdgjuE/TkjlNeYCZrUuYyHrEwj9RubDcFB
QUf3IASazqD/O4Kf6yWVFDatWxQnpsJRHe5QQLGoLDEy2Qonhm0wlPqqr07MIfX/
j8L8Z6Akt+OfmE6lNz/J3SktBJ6wjbTRd10ZSWn2P/UKmqOGV1+2T5LtQ+QhKpHe
nRkbp200M/ZJBs3liC3cS/sxOWNB1k2WAqDkW4aarlAs4dFvPgmgKQE8iMqlhq68
GRQxD/vz7904544Gx99HBVqlEyZ8wc7SQVNNPiPs/KcZCoys2aovmvZpMl/iUgOn
zAoehCj0vtiTSod7zbrdjbjAEjGhxJskFsc6DB7y4+WX7hIjvHxGbB5njvgVYMR2
4BxMuF70bCqALJZ5UIpkQ9rlvFfyaDd2p809XoS03mgIko6AvwSXQbN3L8gB7rHk
PHhk8LEPrypC6DOfwQdte39rbEElXW/Tr+eCYcha0uyTwbMMlU0vdSTMEOejYNQL
1LdfP/CfmGQAjKvS1EYjmcdwsGg/rjWn0v8nN1zk4e3Sd3n+z1ZHdSb6nF/SetcX
mdiJ+rVeiZAXr60W4nqp5sj/hgt7/KSwsx99jpca+4+zDNPa2wW/lNSNmrpt00ad
IvvzC6/Hzdq+0tjsSb7kzEBJJDKHX/SoYmez5MPo3SMI9wLwng8kyouGUewH2vJL
aiBcni2T0dQ62B73AYLifmRzeWMIvDy7rNagTbWGaOt7bE45UIzUGQK3DTT2axKE
Vh4eYluUvrYdBHaIfa+5GaIWLPlVSQ4weCId2pH3Tg1SiuhoMUR9znct+w7aqvWd
SR00vVVcEpTsR9rOjYoUrBjp1oWiW8zjdfmquQJVMJ2f3gAjehg8hGQmcHcjcGsm
Vh8yFcxRD4FvBO23rTctvmSS19WWJoANQyjf1MEzRkUDukP+0DVjf036DHOsyjSP
x9Qdakhf+68IDoKJIWMZmbVpGk+KPfrKXHBkLqQYLdgu9QKqCnKRwiqjeVW4t+Fc
D5UkOwxkSoxw3takwKN45CH7wPBayW7s0oo1iDZtvEU80yy5KtbPwUbPsmRvxlzH
skeKEZvGXRFN+gJOJUDxs5eO08w32zQl+tIg+aLKRk8KnWW0j1F/p0p2nWmE2cDm
PU7mNPa4+koty+hos66maATC2X+QkqNpoXk3i0mIl3xdfdFe1/RHm+grSugjSUCf
xF9wreX3QV7ZDU4eQjZgUwL+WexDu6To2PWGeiBTEPFKtypr9VNR/KpwhH4TziN8
w+nH8pTCqWVrtJTxRT88CaeCbogG6G2LUYHcjkiTNB+Gu6EKrKxpfkXLj/K3o4CS
WzgHtosfnaOm0gRUT/XZPOnh4/32nY9ZBCLSz/kFTa0sDv5agAD/ObBngJ5+9yAo
z2mg1gIy1jVUpMvzQ28BRxFZBGP1q1lJv5ckSepmGqa3hlRZ21S98fdgdWpctgqP
CLaL+Rbp0/6SaxoOdwa39TIiqv6pqAlP5E9ttiDcU3MUuCDgTtDs/PjjoUq8EXr+
4CqcHY8blmtUuq7U3ojw+DKN+53prOZDP4387/iMVlNEjmoV8jMn1MhMWITqB3az
sNL+avQekus4JzVIX6+AlsKoKe+4oooiGPHhItFfhHK+Jl2TRWwZ7zHt/NPU8gKm
1e+TaEVVpFcqpcaIfSQ1B2h23dnFBnF+ygOb0gJtIHkNko5bc+np/hZNGdjFbDnn
UMY7QMzaju/t4r2ETb2d1J2CWyjxaOkfLb2SseJa1Rkf2Cy8z20j0B8bMFEzR/xj
64zMfuMB6B2cUV8Si/N1qcdtWxd9+jh0nGuFPG11isvX8U6wgbMFmOLO4YEFGOkI
g0Y0WJ1c7bEalkTcn6wxClwxfi68T7yXV22ZchZT2aKdo3OdxJjQaAMANMUwPMp5
aWToghH3pQOnjst0zbrJkhNo0KGQwVo1baXPGuKdKUeBkBPY9pptQWmKN5u6Xmo4
fIlyfcHYxthZcxRs1GtlAWsg8EwpEZu8E01/Os3ZCzuSNPAFoXrF6/DX97wtCqC2
4oMcySnm0ZthSG2R6brszEpgQCa+ToUQUpvWN/dxSKRgOjc2A/AQSwYKKBoHLn3a
t75bk3G7NYcDSVDcnK0j2x+fATVOTztEfkbzl8o99apQqwQ+45+qL1aTzw30oQui
zoqLsze6LCRMuCLdKoilm4RNkPIcijmyWfGSFeeXN7tOcJFdx5BkeNUkGMCK1bMV
d1wCWfns5uIBJXph3z/zds2Gh2QlS/PEzpj5T92ZDljLRI0Vm7Z4SN1cqRz/7UmJ
2yXxrNc8wZcXIHi9H0sVdyG+1a2YBxCzy3RVDEayzPXyX94ZLi9w5J9+8k+bDHfq
Z+OPZaVu082h+WysAsutNyO8sdtd/YuxkMo5NDmY7zGhvSUWhAeJx0B+EbXSjT4O
csMIpwqxvA/m14HaF63VuRm9r5oYwdpboow4WG7kF06uMtr6gjLL8wBYFmK75JTb
RH6PEs/Ty+rdvk9V7TN8TDSMdWxiYjZHaYesPkujsLuY6GEeo5o1A/2w8VVMll0R
pNB6WlRPi++njVugcy7sOjKDblICEU2kXhiXjFAqb6iPhQOWZrQy4Tswl2uByciv
DoP0n2RzNgcDZLWqZIOgwoGGb2+RRXkxQYeLaz59oiUujtOwJXPJRbEF1rYWFpQv
2pvQZYTIEhF4K+ujV9ZYJwfbb7ptwVSYCPU+qIf7BYz0LS+u3ssiJk4mmSqWATjQ
Bx5nATyEfQNHdyHkW9NYbnf1Nz0rIkS7OxvLMFYbZ88TXKkEQ5uDRcXF3MaYOlFm
OybwfvRZk/jjPyoIA40XMm9fwE2DJQLcCVga5+j3DDKNehA18vWxItB2VVgrBeXG
G8AtoDYwugEhbBsmL3gUBikGI14vFs5bnHw8ySm0jx8+6xu6eKSD7XW/n41uS2xI
H+S3G4Cf/DsXWzlcmKeq1gk4IggZV45YHvfw37vHB05d6nrrIXi4zZDfEKwIEIUr
97gYpiZFfjbiNZDSH6vQjt6Nf2A1izO+SePPkUBzblDa4WsUPW3SuQGeNQwc5LAG
SHf4xXqFh2iF5c2ViRppLQ5sWRG03aVZPzpPoEAaoUcK9XL23ZW0NrA8UPHFdSw8
ASHDZfc5aLO/PfpilcCtkTY/Q/NkJ+EvPQUHqL1ZatGskrjJLTwZZhThEGXKSldc
Mul+T5qJKKITdFrq+p29gciU6BY37I5e7+7ClUjEinbXJm70Kb8TNbateBMDjeeU
erUw07b0HzRBGlnUbl6IQVTm8qpnAlWfxxGOXCT9KHQf29dcnXgvAdyzECVudpzG
K+Pp/WtQZCh1TF+XwJrMYJNKx/ktZQX+NSabXWkQ/75w0YnTa8FzNCyvuyRfRmib
6eWo4WC3g/QYrfu6mSa+C8aM6hZ2VSMD+pcMJng9sW+68Fabqpi6vJw1qhBgaNGF
RcBs3hbL4EM12lQz7WrslzCBmc16Auo6wmQrtFcOju7/9L+HwSoXHjpOenuXax5l
J9duyT1N6bY/p+Glu821Jws4+fXKvqt06Vg+x2J9YkSaJoVUDJ6k9jNPInKzkhMZ
uMDoVOwl7PErVWMmEKPoO2x03vpfICwkYJYO2mqtc5EziMRK/0Wi6Z0dzNkO3xju
UQU2HAcmIl41YSo2G12pJM1bYb8uUwYO9cVYAbtFS9gGhr1xoYGauEwkuhzPZyFs
Kw0oexCfk2QADu7/oHvdlvtx2XBOnS9UXY189QzRETkSr5o3yZirBViZRGZLnqP8
OhqN2TJI7vzWiuc+tCfF0ZYmC80hf7c3Tn1fD76TZNktrwu1fqt2ZwNK3o4Wx86v
pCHxWLpowVZS1LXgJlfGtHxh4QvDg1UwkW3LPSl60Od/myftWtdWZfYxyoZq/z+c
gW+ja5mpCD9ZssrG6tJGT+vLw6aeZ7jONlz52IE/tagjMvxKak8G2UzIvWf3rmHU
jnd+Gk2olLcyhgCVuHJaUH52Zl3YPFq2OKY+wkAfGK/MjFXgRtOjpqZey85NemMi
k5V2JdCGJrm2DJh+l1CQ+cXGD/e/MESIvFy00Nsjyx2YglHkX1ubMqYUeicrw8o2
Zasn77MS207fuZLJKyrDQHZduHOKKWCEKZLkGnBw+Bo0XebprMN4/EArVj29cbEI
ijwxGiqpX/CHcAiB+FEkrTuGb79qNhLhvnJUF2X2nD9dvcNPGTPkxgOAYAjo9FCd
YsUpdPHtHBNe0FDyzRia4L1IrUM/YhS2+gwalWllmAcB5ZSuMbC1Rwi/v8kSoPy2
W+l4UaUoLtYe5GI7yBYw+eEb9oGwSbkEiz52AxiduZag813uW8aeuayer2+H1RE5
Xd7gpbC8MncSQ7p0VF2kKecuHG7EUP44rnKCqJEQGDNiiwg1taDmS+1SuOYxezBk
bCpHKVS/uLq5Nz0bm2h1HB7bhwUif3H+tEnX/+LmN8qkQ6U4T2stJnV1qnJI25WJ
sqRBmDb7VHvKeEagxwcCCQzmEf2hJcLz3SV3/AXdOB1W7KsLmXhFV555i8ECDE7t
dzuglR/oY134mbK+WANMT2nJ4BesCMWeQWVK+ERuM/GiqOJcNsag35/fI2wr7ihB
3ubTOhEYISBA1KIbmZqhbcGDYVudBx5Qhx8XB0i/7AV3MEwWSdW19e3LGnyDRtjR
XYPRJDWlr1gFwOZQhDxpIn+CeVSk+h/Mmu9/PM3+fX6xSeFvXVip65QifZDZSM3m
DLuFQTEOIMoHQ4qdwyvvXLBwhn3AE1FohRqCsoeXFzXWkp8plaPwbQayYx7sKSdw
b+q5kfiaMKbbxFqU1lgwxZXErapYjoLD+WcX8LVjgWPOW+aTDYk7Efw08vwFP9Vc
yn92WSi7OGr5YHSJQBqkCsyL2qBAA2VUAzoI0wxKKck1ocLsQ+EKK0O+Lj9wJ/SU
SrwP/BrBWCxarIWxRtotXM4qZwJUFdb36ayliiOJlhuRzdhZ1jVZFflNQaGxetDE
nZVkzecJSWWZEOWF2vFal+8U464ASbUf9OxEaprQ7AEKgO4A403YhuJfKQbxS2Xo
KRG0vPwPReqKLTfpqzqtV5sg5d3jk/9AH3zjQDCiGbzkOcAr9M3yF8KL0Cp9Dk3q
loyKrQH3PnAyu1HhZMDllo54QMIts8fT2qtchJs2KeSoj32a9X9BzRYcJsORnFRZ
pg5NmRxAkjKGOqyqMB5tuZFYk9nd3DGqzGLbM2aaABvGQkhKm9IiOUlDOTe7a3pB
oTn6EP7BYWnI6q3NAdniyLPaz4+mN5IlT9BTdQkopt7jc97Gkl8oB92tXvweNnqM
PEcEAEuf21Ku0l2wz0reTo8xeocxgvkccJCJuMeluiejD8Y1k0RahvQVjUyIqMcd
z75Psx/qokwG+sy5OmJaTNiJQ1LS92MrHsxppB10KidJTjKVYJYu5dIU9P+HS4Z5
apIKSMutFbm+8s0TIj3ReDfqQxStbUHVZdyXiaRRMT/SYifFboVfkf8J2auB1ALQ
s4KvA/nAuqruv1pS09R4e7iiafHX8qaHC23J2VjWypXwNfsK6gwyXAEbQREx/CdA
CJvtYhQQmWbhfXI4xEeHRN1/9FdkpBt3c1sMQGTbEptvNxwsOvDfS7Df3vTRL0Ep
7BVAN7HUiwlMj7RPS+6R9pGvJ/zAAqkL3JhIbUqFM8T7qnMLTHHLcIZxJaAFnuql
opB1uPDFFF87Z9HbI/FDhY1OQnyeexjRuKLql9t+tZnu53izFgPGorciw5D02s4u
qqLKPW/YWLFgNwNI0yS6XNLT/AbpD5/vNml3ougbkDrbFNj5W4kvBIG6xrqZ777A
a0OPQ2xNleKg07aJjrjvZNjxFafjgbSMkRQzDkda19AwF0cUPf8kG2d85kr8P7cw
Zio0QZNKB9LaxCEh9rhiHkt7wI2WmHjHcDBU67coYBE5AXH8spsvVRTpSjIR5UxZ
`pragma protect end_protected
