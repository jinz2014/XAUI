// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BHosGAhp+keHCH3+yZHXwMPvLpTarbfk5pLvw/BH7iuP5Oa4zv1Quw/pLqmADVqw
M3GRvfAERBHy6Y2OcXMp5fErl/hTrGNP/14SXiDfKpdq1L+KldX+mYEFhWUJT4gP
GnPHeu0RzMB7I/hX1EfgjHO6p0k1xdUIS4bIeWq6Zqk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6368)
p9V8br/KPig3WtFU2okybIUO1610FiNYogNP0RuQzZtrxFohVHHiJKXuGPB3GMOf
8M1v1YhvQWYQZm/terluZzRxUWnzFXcUXnmV4ru1CjYusURUPrTcOmU8zoK+hc/7
c7+6V1FNBE6dLIWJUootl6+KlGa1eWRvon3YCusH5ObB1woXhm5mYqktgqFIyioq
nUmCroXs/YlirsosDoh9mpp4UHD2jrHGjtwQDpNPVpgeHy4lSSBKP4UW6i8UwiZ4
BDrgqreXYmNUclUzYBdMc9O9Y5foTKx/d+Rt7IgEPQHlE3pXQvFUP0CaZjvEV9l6
ik5ZMKiR2NusOIStBX6iSG1QzwzttQU/m7sTjWixR58rZTeWmhCKAP+wreyIZ3aH
LVlVcaKP+V8rYewUawZTPqUIsDfnGr6zGBFT5BE8LtXkAWPzoB9ZrZEiNDCFgkxT
wFOolQyot2jNVc6hhqj5HdKIkB/TWB7fCteDjLCRVZFJ4KHF1vw3GdX8tpSVOA3b
VMY7s7LUAmyfsyIesHggsqVqhQ+lwVUvck5XskypvdxWdizOUkma+bAoLD2n3Ium
LBPUdLYHbk/lYkXOyxV+ABBk2klbzDfAkd8HTQMmAXCG8vT77U5UW4aGorJoOq9B
pPh9fxVsfSg7tc50XncJ+gw9jdRglZIUojDFIK7azWE6zwvyVDVZH0UVu9+L4qFD
/bqJYk++9TWkt+QFgryg1U85YqbCBNMKDv2prFiEQsUenvCcKBDX4GryfuTSRktD
bsBNeGlQ+8SDlUOYDYEdueq/C3uNfDgIV4E9ftd7gc5AG3BVzNoTu4RBUmHt4nFC
0neZljwPpjqPUClj1ZOJzzGLvXNN3jJHExj611EJM/+/zvZ9vKseF6nbD/M6ILpg
vK1GV4rRxvt2sk65uW3VupoJfB1IOyPLb5oPD3U9p5OZo47AAVcq0m4UOiemZleL
nBNZdzNWGdM0EUNg0QXaE8w1I+SGAgsvl4CUMKvVA1Wfv2btimTS4gViTx6zy9ge
9u0CjHXP+L5qgXxZghPcCk0R8pQSEygbafOH17AXx/uYTJy58nsuDWEYb/YGi3GO
33sQvpJPaZq5dWc7ab9Z2uMspQCyeA6dgqaqbbfmf/AlcNDDaTdu/Sm75IWvqhFm
kRZnLRIjmSDWs5fLMKxWFZLZ2S6P26HakR+4P4uWGZMYLyUtf+jjFgfaZVa5HIPa
bEzr50fiTXF90Zcz+jB0OAptMQYS8s3zyL2vG08+TMx2xxUxPKenDUvwTbPC/Q9b
e+oF1kCrVc4kpF756FukoU6Szn8rNunniOopuY2mtAdIryLrxoHR+OX+X7lpkPL9
IlryuKPwtF53DeJRWQt39EYL1opKQLA20DVpH+kIVFoJX/nJDjQBLRqoxo0u1BQn
MUdj+5sQGL/ebigyadpwhfT/0F6BpI+lCrdHl2Z4loypNhiyElEzbibxR9pK1s9c
lg2oHVecVAUNKN+Uj6abBLIfZ78tqNuDiq260dCUK1dM/ShfuqU+Ge0WHjNz/LZ7
OzTqwHwEoM88n4AKORkHRARbd19qZ02DXJw+vfXcJrm/afuCmvu6shqBjxDWh6c3
bdLvqfpjGagDC4lTIa90PUqL6813eaEKuOcsLJrvzTEHHMCSSuDs6aaH3Fx7mFJR
XP0BAQ2gPyyDGAOTWTAPEiR2aDcQeiXoEtpXqvuLQyIyKIK0JyWcgYArK1FusdJ+
7JbzuHTlsTRT8oeIRTdNpyJOl/5MPkhszWAIJGKpeVWvX7xXKef6mgx4YqvzdZYZ
AbyNbmKx0yoY7uiltSUZqi3g96svGl0TvctdMWWpIqzm8HMe/Zb9M2F4GvSfnPse
jMqnZAMzz/kM6sfcw87exxEEfJteDTMoo/eGLzE0miiQLYU4O44jUvhaOl4XWwQy
OCE1Vz0CIzoTLnQl+fAMuqppVCUXvw6pyn0K529VPd1JdL/Dp85gwX/wf4Sh5/fP
ddBssfAPjHyvLPkZ6j1fIKHhIFIBuCtD4mScp+AuN+0QfdxkZRfWUxxdYtCQWp3H
irexGcRk1djYbuGTl11b2P1jsJyoGlIaxH0UBGH4FHbgNXi19ZeaMHkGxwodOsOW
pfoSX3e0peVCnmbQu6+fnbQktCo0M08ugvQhsXcg9G7PMCv9BLegkfFzBHUI0Qyk
jZ0Mmqgj5GppPnkUnp+JNb2bZTFarvrfFPEAOvRufmRs1TiQ9H8QknJJ2yFCTA/3
d3pJJVzY1+CX9fgmSMZhgMl2DDHmESjZc+Z4q7GBvDhc5fKjxf8ccDBbW+04aLXZ
UtG+4Lm1K6qe+45pVk9uQbVtYZzkZ4teFJAPaKhoazFoD9VDK06wc1hTO9Mhr1vJ
u6Osp71jA9QLGBBdxk2uqahXYF0KfKPdlWaoC9qy7CIyykL9ROS9s1u44oXpYbAX
OCVor9MByk2wNB7HJ66/RGU1DWt6u1wtB8oP4wSGjNuC+UrrMRFsPXWSJkR8BVNO
qaATNEhoaG/TfUR48QoLJRYrV9J4hsNcd4HCmfz2ixd7CEzSkYDby+qNzFMywLUT
CPx2nW2BxTpcNs8T9unShaHaG3kZ/f/4X55wju2F5VgFzwtKKK3W6GD2VA4hJ0mv
2VczE7XIrSftQdP0e0L+r8u5lSUPJRGMEEHAow2Ohykni6rIvnxSQIMJS/mn26eF
GkxrGXKfgNZt1RJ3+TTtP241krfzaPEA1/x6I5wJj65zC85kKDsXm3b6s6UdnLhp
ePoz5tfI+PF/Oq8lMAyAWt78f53mmeVBEsPF7F6iHAmpVm2vNg+V9oeB3jMome35
SbsKUp3axALC7R9PCX8NL/sIOFng//tspwJ9RiBd1zK+SF18RjtMb8OVogLmdx07
5R/LwKY5dc27OzIgoKGvR2GTcx43bQvv2aJna/kC+qf/r+Q9Lu7BBlvuXsnTfd8e
KtWw51kh7T0ZO81/ma/l615mx33ek4rWZD5fnnONFqdod+IuH7Ry8AZpZGeJHztB
bQ4DWFlKhI4ONWE3ZsbxehWkwzgzrM6Ksw3xmTRpd4sB+RCPa4DL8ZGu4ETWOmyp
Ck/aPIXNUxvBmpgGDt2ur4S2vUNYTLMMOKgswf2vtqQbK1G28GRLR8BzckZxOJIz
fcWR9Z0cHoAR1uqN4bc3F8ggC1F+wfIoDWAtpEOMTMSs2xpaeUUtb+QclwVlGld+
IbHa3fqZoWBkwB5RF/64B6N8L67MzMrVnIfW5Xs2WnejZE8kFkpVWsCm6MRLTh61
M46TdsNYTA4krudXIY5vcwSoiUXWM7myrSS9MuIUhX/qFbkcC6FIE0BZB9RGt2fL
l0r0BgC84GxE2K4oNxWkVOgpykBB1JA2Tpp9TeRMyHZTh2DkLNUlIdFgz9U6E4kp
2LG0qS6v7g+wJLBxIA1QmXfSwnDmhPe0ObtGI3aOT2abRyI+L5mw4jyrn0Nqax1f
ITFX2nLCGwJYyhxSebyCjh3b2brmsfXzppBn7cDcZ6SvosxxM8O52tWX1b+BvNFf
4VoHVW2AspHLcOeLfx06w+lnSj1Vu1zWv8UFTmzrBaZuEZ3y5t6YU9bJPz2sCX7P
cCLp+Fmu/Hgj4/efkUOCVvo0FIKND8RJJLRWloiLnDDQHlj7+hei92iou4yInAtA
XxXYUqoQST0Vt3aSF9gilLQrOr3SUuS2E0gJzaHEJntK/pygwNgGnFFNz4nec5HU
2R8kpwAAw0W994kU1Sqy23Xx2qIBPbJoKBEQcBAKIUW+nYFl0e2ExNIUtNWDXZFB
nc3qt1QC2kBu6qSzMYMrbi6eDiyegK4hH5/JbIWAZr90nAdBT+aGnP2LAv0Tltmz
IKMvLyWN8Jk29uM7Dvqt2XTZtd4H9xKRA00uLfDyUevqZJlvaeLMt9C+RGX/MYh3
mooRxRpLmIsO539JhJ120vZdZzvF8VnBnmwh/Rld19wJ4tOhQX6wzWAoy+21qkWt
jBiXprIBrsB6326vL/C1yMMznrkDBp066/B5FSvpkDZ95Rjck1HRfRgBd3fnGTj3
zWgrsYHw7jgsMk6rISIDKtOQ0YLZ9lisq1LH/ug20JdT6wzFuGN+abY4nSA9RVEU
g1oP43GfL7ZeOcl+EeSJI2PA38IFSxmy8TkL7aNHYghDE4EpCNi+Sgjy/OEhypAl
5UoYLLdxa2p/Cidw1DibseE6DQNHAQHzqgz+IRsKviBoRbFLUexfJKTeGpS7RYqh
J0cPZD5YUT555E8My1MnKT2Mt47g0wclnSTmWA8xqQbFc2Q+AhjmE4lR8imikQOL
gFvulHw0SMa3wM2wZp/JA+BbCXs+Q0cVTO8+IM82eeGnQh7w+If1RpR9Y7RpCBYy
zHJOuqULPPdt2apcxeU1nsI4mu2GYThfjOXarZDPOEhNrRh655nndrVX0bOmUd8W
G4VNOIgsXQYbJRkMx2k4bsZVDMGBDRod3x7KKfFS4CfwlIMLMe80kTKEHesmgIJ+
VDTlkSJOrUO1odSEltCk2JADUjXq/fQPcZqt2PcVDkmgI+IpOQXfLBj+LK0iBq6B
eckMSivuuzIfoATR3CvxMNdR9zLhhW2yELCVzUUoLvNJ7r+iqXv2SjGGIapYo2Wt
N5V3VmNzFp8pKMK2IKbi8uol/jYzQXpX/Zbkb8kbxlrU0/KXHkIzNKTnA6SF8t7p
0AnSRRdHtKWoyyACBrtWPG7MuBDoUZm8pHMz2U8BU8LR2f3FuX2Z3fCcxT3tew4H
fyvg6hbnFVsLrHPJwkDPz08nQF9pWKaseopQEaKrOUuS/xS8rvLIC8lUddepJWLy
rWYAQL3+ya/ncH8ZFCyo3ZkRtmhP8AScDdN3TvRGR1YYGXKH4qcu0aiSk6ZVLrcF
O6XNDitiJ55lgtr4hYOny09grcY08HgPjGF4h5gkOiJ7WHESICoLHSjzL0pBSZHM
qL1fyN4I/VyIyocXppHKy8p8qU8w27ICdVJR5S0msxIcp8IuJ8C++K7F/RVscLZt
54aHF05l8k1k0g9Gmp99HPlqjNZyQKBamaJQa3Gz1p5CUaz+Br59nsYnEQBwdv/L
YZYTCq5+yuoo2JaUMTI7YINhrNm6Jd+b6cj1EoHKoP7ZAq+ITVvJo9a1/q3aKXQ0
f9JbNNZwihlWxfXugX6SgRXFeekQCVdJ6d30t6AYb1yPX3rk4eY+sjvdWicLr+u8
2uIbIJtEHN2WVXf7GP4bvI8+JSG3OqqEy0+/71rr7q4wW/HTargTrdmeiKy/8AoB
X7ssdexmKe2QVl6Y61/izuVIOP6Iczg6giyzw4GgAQlD9P3rGbCUy2EcuM+B6ujm
Iz4jTq3xBQOUsf0yXP2uSmz+fa6SOvx/Y9WsWfgDq3eTGqys4eunmmUCWOnmfA7m
YwtWJrDTSOhQRh6q9bdJJIXDa7eOHt1EbzWRP4JnQjSlDMuLeJVaZaUN3ttyukSw
PRiDx+pamCX4AnUjtiAE3YG9toQpig29eP5oPUeezQ/AOhSRc9D3pPYQRpwjpmxe
c6MuVvPccb8DTFohni0EJS7JOEOP9NdrJYUmmj9PiLF13H0erBINEpC6x30N9bei
eNwFQWupIZUPbZQGr5ljnJujARN6XhVGZD5hhmMWBwGn2ljUXc6hAnSmtFMtbYGu
kPkQR/NZcVAlgq6R6UzVrUsnOhzsDrYgklePmhh27jy3Xici+GThTNuzzNxE1rlv
i1aC6jAmHuau5QbvXHck7ACU5SINFVab2IL8/sYJFX2xwY6/yPeHicaalJVShWMU
nR40ffrW+ScXIS+p3eTgXrZ9zShV+d0zW+8eX8mtv/FCjcT9OMooE360YUtQWSH5
OXqe0nZ+6LkRaOIbRcURMa2t1YSi2BUc5Y23b4VYTo0JT1/4NnCrzK3za9DQOAGa
q5pxRoXx+zFckKFj7zoFjzhlCEQGy8j/B2fqfktC7KSlPgxeYw9b6V2Y9gACaJIZ
TdgX4xFUW/hLcnjhM3pnGmB6+itTZCR5hx2dyupw4/F7QcbwNKu6JoiP8t9Dd8C1
vV8j5OEv0AKUQrjA8Kd1/3JjxkcbAmdbnHzujvlptGGtxc4DUzctDpuSMHaz/39S
F4CvyKHEpfdgbeRv4x0i4h9vEjnwNY+irp2vhyRtjlamBHmR5fuhxe+GX9B+PA8Z
/p7M1dP/x7OGjKATaoorqlBuf+8mDek3dLI2zPlW6EYrNNkJBaz4j1QFh/Q2DhEm
gltG2Sbn9HDtvv9bin5DGgAKQese4CcPEYSK2JmXEtD9EIEi1LBEmCjkoThWzz3F
8nZu1c76jt//HyrA/Wtyo/2p6616im4scNIRhSOq6kh1ZfzBBbyUi1fqzo1I1SBg
Hue4XbGpwe5DBZ8buCizrRrbXXRPMFE1vczNLKybeEtKu7cHH764ebRFSPcukPOW
e2+yaBVXmo6svjGrtHBrYaGs+8oth0my1m4dLDBV6Fzm50I/hyCxh1bXFinRIEEP
tu9gujL5QVE5j27oRK68IQyD8N3FY/8rM0pCNKb8Asi8MDhardbSTHmbLjcvQKFl
tX+a1lXEu/WSKZvlqkz5GdcTPP0mgx0FLvvmfEHVEr+7dQWldm8l9jFGuTj5FkWD
uF8XBU6+20KknimqwMsqucBIA7ItmDljggXHC8yNYZVExnGVShlh10RBd9jNWfeg
QzY7M0yJtB7EEMG0vEHTnXWTyi2Ru6l/1fWcmMYAMDnQm2luuN9emMUs/zVeX80x
lxg0++TQbwfXJTEeH2s6toDB5uwurrbb5RC+WvlMY+NrAyvkwlo8PpSJCqBVNzpA
+MP6HoyDtQlxkGN4Z2qat0p1U6ll9EEo2u7rUgf8gGt94hUO70cNS2V9wiuQdEDW
bSdE90+M0XOFdYvW63pBXlCi71KgAxbMz47qb3Pu0ylIY8G74ZcbGAF/Nt+W+Y8B
HP9S2lFDnCjGn8VtCK6CrYGJtBwoJJm9utOcAOJ6KnGI+bKgo/sueKz6Q6NVeath
VdJ+VIvtz2eL6XaL2RxRJc27Iab8DTmQLGbJKgtCOLYyqnMypRMu7hkwSxrzCCbO
Q/0LSHW2BPkFY3Izi4Dbcv3fsxCK4dE+P6Hr5Mhy4KwgZ+7wsw+eefKC0ChbpVl+
wv7VN3TSomDuGBoFBcLDrXcaz+qAQ1UWgNzOzHgbI7+0wwh6/PJwzTLHPJSC7FP0
luaDhm83nANUbQwkLcPGuUjYUECpAtmNqFGHp0c2GyKzoYVv44DG2cl2k95dG+WQ
Jq6ezLiAadIA9ehM+HM1IDhw2psfmPG/lq7cK7nqagr4Pwjh4gAMhnz5LxQdHEMm
fdeza7idWv3f4mYx2To/n1Xi3lNg4Lv5Xf4gyFffnJPVRiP23n5Wt6TPmHj9DPxQ
5tRogPtApr7AhTuYRzs8EdC7gXenvl3f+PXMBWtgw0kdT1lq8t7LIDPWE5zw+WPP
+iNhBa16fHBXzZtPrWaoxRaIss8q8cE2WFvcvdIe0yF8qo2yMOBvdYfklCS+XPhr
TIjOwoKi2NJptjLat7p3QUkchsoUUeSJz84a/MFeraEoarlroxdVr5WjBfTa6MXd
ZRdc/CdCYm/Ly2YOJ2YJIxYINI+MxmPWWWHs9+C6y9dMsB6jROK9McF1bp/qbRN1
ayAjSzslZKiAHuaV+MwCx/d9Ws64FoT9BzUfi9P6DJQVlWHn1moR9EgWnaOK1IC8
pH9SoLQAlck6pGebPsIO09pYiOn7dwrMQlgK2/11Jh13iwYMA0OgR7w1TLg+IMz5
Oa0x+6nP/eC08izN2egrrFe4hTWsicMGLZRG71qkZ1XYKUcwkXtGYwEKLFMsw00E
D3Xd25PFSvcmjpEJBgfMQM41BcSblsRnGMXTDwO5eKBWPtKYlfl2iCt9dzSfOJVc
Q7Y+rpG6abfFXFT0DGXygjqSW/1UmFpXianw0BErB40hiuv9S6nDCcwNNXWlYCg7
SDG6XD5JWNDS/kOUBvpfGb54gK6pL4r/W6g2M7IEHu51XaRy7hyoTKbzQdrilXls
KqPL4WsXjzMs6SxkPVL9S6A5l/n1YHEA/cU58/LW7GrC0iL3feXO+C2+kb7JsQrL
yhCUvACEEoq1sHTbJETxpNqq6DeFgWdGe/Cu5wjbKYMCB9ucmNP/+WPpPDSYAC7J
elz1tG0n/KYCbtqDdA3bLvFlYIijplxKsJ9nQ0ohDOKVb2l9tN7nfW3HIooIMVVF
Gnkngtd/ufV+vOBuRqgducBHr7f3lya+dKsEMjs0Gjdn7tGLrPLwap2ZsSNxSAGo
gaD47KobYfmNOh97Up8XRbBOsvslLzRPEOvsAb1XCIPuurJJe8HCppfzGfHgAlDy
vWYU+glw7PLmVFwRVKNPlgkl76fO0E/rRrR8ZHHy7aYvKJ5m84H1tHUXps/vEsSI
JaxDkKXHpnU2VPbgzU0//ZE5GE26h7pyi0VSaShoz3czAqMxRznlDONxD976vFwA
s8k56Ffyn+fIfpGxmssiQmeQ2loD+ht0p1e5fsF8EGc=
`pragma protect end_protected
