// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:47 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Q/GODpXHklgPo/LAcIziFeO35HzKnTENj54/M5dUtgu6B5n2kXwDhSkTdsIVmSR5
guXWlTcvDxD3SCn6upHjW19ZK0WVA5nBB6EgLLJPMItvukZtcxd9Pl12rlo6888m
9FcsPGRjxUCPsBs+Ln4u8OO5bIt6y2IVGolDP785hDc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20240)
gAW5dBodtLTRiry1psgjrCfZd9d67JrQfkrbLhwp1gQV3FNkILweHhDoY3Ho8amY
spTuvb5r+F8QqV1OJB39d2p18m+Z/tqYGpPycp5tjeGNC7YUC/PpsDTG7keTbCwL
XOc+0ARCaOSIrYaBUXwtiV9s8UY6l8ksjfyagfl0m2n0QDKfitg/juIQaQWPwHiS
cfMQVgQDTZDN5Lu/gjV8dvs35xAMQwlAIl9jm3ya8xFwN9KluTLOA+4bs1nEm/Js
md2dP1RYPlgG7AD/do2usd5HTbkOBvkd83SmKrzCRFE1tSAMMMO/IoYNNqzV6ce7
Efj/qrnN3NtPB9ToIuKkuWT6V6w7ORYyBnxcr68SnUL+2sb01ue1GglLd7/scTKV
vhsiIQox9GS36OnvySHehel235kG6ikSu1koQKoCI45KkjbxgAGWiMSHrR9/Q2uG
H1RhDn7MtPXqJQ51bNj3lRoPN5EOK42Gyhm6+8XWBTS5z/xi0iNggkEWxZz+k1SW
Pqs1eQWkzdjGB6q3C2Q2SAz8MgQWntZCywYGkvP8ZiO6Fln8iVVh7TkEu5JdnD/l
AXNOS9EBfyDxfff6L+gPpygGXs0CctfGcd/pTkj3cb4qV/Stmb5f1YJX1pGM7+Or
BwffjqpK4WnbtBEaQfg509O64itfjgsQSEUNxIvK8aNnpFgxY99mfjmXQ71OdQaX
CPHcOl8IYmMQfWVsiIJ1BI31CFa8famI/0OdjoEM6pS9iHx4DhjWyZYJ7rqLJHYk
Ss4XaHl+YG/U/gdnfOyL4e6HzYpi3p9L38R0f3BC0ZC7aghmBmwODSK7JZD2Jxs7
hKSSA/hBnxQRal8ULRRrFxsoPV2Ea+a0XLf6qtnj+z8Jfn3BZspofmEHkPZsq4A5
gm4EJNDeqRwF1p9pTsMIJ2E/g1Li3NlWBZGxMFSGa6+0/nBk9Ut5buBnxQowf/TH
Dtm3ZNWNXenAMV0z2TPmPlwzixCa9/fluWsarS5LV0bSxFit83V/A/46XgRT90cP
vkfis0UnxOqkJ98gB/ynnvc7Q7nVdEEID52hdI8SoKU2NVbjkhDMtI9urDXrl+Vh
ft0Yob8U+PCa877LHyVQBVUrcJAs8NPCZlBFO5jRRwaLYj7klS3FTjqU3qtumq7o
UgnZWeEu+efw4ZbJd+Wg39IFy+MxvbTsGj3I+Q3zLk+d1WCXbnfZp6r/fsEkSOT+
CHC70OXTcPHs8lFnrRIJdfTw4RwlCHFyEErRYktR7fPi+bB5dZjkX7rl1Zj/HbJx
J35LTnZhqLEgAFXH0ucB02yuWbgOuJvg1Llb46QTnuMhG+Qai0Pi8Znho7a4jCfX
4nXc/NCXDVFa/1d6hhTDFtSuoGWukRJOXnO2IGpxIce7kTXzgRtWCQrHQamHE0N+
Gm+CnuzU4wGNp4HLiN0PGx3YiZfHRlNhf9pV1CKVi3nXX1rCzAMgISz0j3B72Nmx
LkADLsaPYmyTHp2wqUXZY321yPJwr4MenEwGCHyRQe6ingVm7l2tEv3LT4qUNmIX
IJxnpqYkFHHoSC07Lh46LcD51mEyxPZw1Y42Xf+w7gfkSXOetV9KDPXxfYkn41ow
IP7GaJNxhmCfa3cE9zImaPKO7i3O6V51w4QyQXQKNj/AW+eyAR21rJzf1tumGmwH
k2/s0ZZg4oYZ88+OW51T1A0aDN9amoQU/VBz8cLn+fu8nIvYCKT4strrKWPtSFKt
FmeihDe9Nh+KUercmdRoVRFrwLrH80nCbBNdPlHqb+cI9lEtZ3isgznNbWj4X7RU
/TFNRg9v1HbrEBPxT+q6idOcLVwLoCdofJqFzQu3/b4KaWyfaiVhoDpY9UENGsEU
2tsxl+w64HMShqzKuwdIBgkjb70Sebm7cCyGW5qdxvteCvvJgJEFnUpuG3hPbXtf
0/dumwaigS/ofwAufQ8Yd7CK5shU5q16LBo9/DoPe4n7f3RgffivKtLgxyat3mdG
DcpmHdiOWfDMDcLn3grvdGtrdy2x3K/QFDwPNYEeKMBtQyRhNhWvaPG29yoa4ldX
cPaCYNlAn5Kba52oKX02+Y66+jBzMbGVklXkUBnoVqkzxI1LAtlNPzb0+hHCYfvI
+AvwRdJqxraFW+hSWimocjldlfKBrOiCZXmP2/1c2irMUfqhVY9bDrC+pvZqV46I
qPaRR+nax8p2Ld7ui5eNUuoGigTcZXbxVK+SYLarcQgsEgktcYewpYy7mNSiMeDy
Oj86fagVNUDFBaGAOnYbBu7hzmXhh50/3jtHpPDKibYBrOQEZNl3zd+7sBwT+Siy
2eWGkbJN2OhynXfJ8acsO9mVr9E1UvyssCEGDKAf87/H8Uxqm4tf5Li6cYconoEb
9a+Hp7EmuY6tPEqlUNTaJlOhZqLvYnoqEzqa7Mua5CYVRPRFdb1ZgkFafwzAmYp3
rX2JE8HkxNp1tF2dBP7aMuzG1w4pacDpojwbxu/vZzvBeuz6S0ix0GbYZL9NBEWM
5zcEKu33dkamA0arTDVt2EZsSkvGpK+OXqHarZLLQWT56Wjb4jipW4ArwF+JvXl7
SvLXuwB7LGLwtjEiC3uQWiWM+d0DQ9DDbOYMPXF71y6HZOvGMhi9weuxvtd01/C3
6Vc1iptYCvthiwFHKUPPN/PuuOxebZNDvaEhifhi8xub5FgiJA2dd/MsRQPz4r2Z
uGAnhdkDMiciql9CF5IKntZktfRNTWaqgxG/wMoPNm4/BBLW2m0qzLpLewKpqBLG
uJ6D4stvLjBCALRwwXRm7aMuwOkAwneLH/WQhByw3xBsGglld3Zv/anuI4M1hwvI
i5Xkq+p6fVcyH7hgXFaUxSU3lkaTaUV3LVCviEtZqlbQgA2Slojifw4wptEPhayA
VZfy9bgD75zabq25TZVXMsePPMbep5ZXEeRBZH6zQN3U3iYcyNiyF+HWbl2V3azh
jrZmlU1CU6cAVtB9xLY0kLnfBQWAI4w8fHRLB9spwDhwHp/ICiCY+z57ksmQpIjl
X9DuO2tsQJUwgWepC7A6Bo/w887DDEPnjsoGPb0lO+DqjqIABIA+ouKzFBRKnGbI
ldaJks/LleR4k+fPoyDPd3i382YIHPt02w6BSK5HasquiUclAwamWH0SM0AQeksD
BK42Lg2TOOCETJ/rs0EiYQlX1MP4Jw6ARvf+haCrB7bzq4lgfyaRzSOB5sEQwJXh
2MftoAVWfY0Na2XDSk4K8r3JhH/+0f2ekszwCT7BjzKE6dBpclEuAFYYJspXX4Nt
wUIG2/1CSCjI+pqnoOAGCCpgfd/+WGWPAoWKtI34TANOv65jz7fJYMUZLYTfM654
xGXEW9cX1ionaH87Bl4X40/PjzfoXaKjjs7AbNdR4ajkZN9uEx+Rr7Fz7bB34pUW
T7dEi7Wes5pENwe01pS2rPzURTX3rdMttJAri0TXwGLCdlqfCc5t8GZCUeVPfp3h
zY6ZnDmILAju56xu8GG7Wqbsu5386jhhsjJEoXPxOIXrBH5yFbfdTOM/EMEyTc9T
wx3YlAFxJOWKvFxeI2nVIMscVfxqsT4Pav5HnKBbJA+7B7I2t51sVYD7xwjaRT27
/7hdbn04DLgxlmcSrUOjwUD55vYI4m+Pl8POQ0MbqhPKpkIb5bLMUjnGy1CZTEkK
3WJ526qlPzeLBeZsXXOto9yrhkPiIlv/psyK/f3yjSCUeU4sCw14WW0Hgt0MNPOA
xgHx3MiwOHegiizoirHzbnD/0Slx2bPKg5gHOmJjcn+Zctf5dZ8PnF6KjM9gbuRw
La9PIrIaIF416G/AFhBEapToOB/SDcyj0KnXtwolSBobMvl6oBSWKp3VNem1WSKF
Uiqg2FtJRqLraqWXBj4QvkGmgckevPEJZye4OvJmgk2rfHD1yHFHHnGbt+bOEj5G
4LIl3SJNlSMSJmwUOoPgo0wyhI/mgSIulyRqu55hWDZwMdiVlR4+Dp2JocBRlUlV
4/qI576X6kufQ9cTuqFA0mFEiCE0wulrzSQ2fZIPv3ovvPKFwCbpKW+f47/a5Hpo
mrhongMuPdq/y2NroAaeueHpmyS6BZFVIlsga3W0z0/5eAUfSUfGrsGYa+fU4cQO
VN2mG12mBOUb0iskHeQs2mgs1IkNMBSEKk3uBXCwnTDgfzYIKYIsFg1RiWiCYDeb
T0I1PcmhihBsHC8aKWOFIU0ptXtpVSBomBEi/Kjln7uC0VebukF2KhPXflsligkg
soJYvulLqwoS9T9xzC9eXRxC/gYuv76TA+Er/lJiVLsmWM/r3q5rwok4EaX6DAB0
PgIpNB7bVBX06vm8z7mJc1+Ci2yooTcxotPu43KSl01jW6gf1Q4OFKYC0uIe195R
Mx7D4TVYoAWr3xMlGDlxq4r82TL0YIyh6iLq2zFaKyldxggKcBQcRUqOkGdQhdCP
VrlcY3CWAAQAmerz7uohxURPsB4npZBMHDrTIQ2bThoqK7ULdXtHqT78WBooEHDg
Tr3lNT/g7SW8FjkFEDiky77yPXxOygv/3eCxxKg8W3MB/Lka3/+/aIVS0pKv3fPB
7bAFJUeBOtnmvfz8EncMp56Kf3NI5Eo0FGn4SrQuhlIZ7rAbVQlEKj0FLgQpfnnP
JzXK5l8SBYWupZFQxTbMplZw3+pAYzVIP6CD8gA4e+EVvw95rSR4TJcOZbl0zi2w
qCUldIHzv7C/z4Ynqb9txYdf9Vb7goTt+jMw+JcPxly/LUqbhxEMmyQ8WSZImQz5
DjZ8OVCd9ovI2Ga8JwBJzRDmjwEZ/ASd56c/+4CV1iip6ydChznJ65z24e2YUcvk
onmlnCO0RwOv3lhUgyABFe1ypYAWkmarPaJY/ZqfpGzdBhGUyUarqhEBX/+pbswN
xpJu7qErKoH9O6dNlJOrIW0Nbolr0UnlZNav1X/p4kza8thVYg7/cM7fHkPf1cAv
UoqZtUjHCX3qTl9gSaXgeoey2kL66wm6bXKadwuBYS489Zm9KaMoegjD4SZf7BIE
EkeGak0+D8xZmuOALDvr4T0T5kohU10JIm/c/1yiJPNRPpEp+D7DkACkJNdsLucT
do6Wh8FVZwtLIElLSwfjcr3w/PVMpVyD/uD/MVIgi0+M55jPt+pzOXwarR4In4da
iipALmhfnO/Dcoq8nUzZDAGDWZUBSlFDrjZC/yenaq7a5RrYFQxYX6Kx2jj165zn
+MxNoU1XMvn8L1/wh7vlJd9Qq8FxgOF9E3R1ZqoMcIzKrouvpvS9xwzX3X03zFVU
RA2XkoRpB7lryzQElOfDP9UAUlD5Sym/C1ynOdjEl5k3Wc8xgqAQvvn/HOAD9pU6
LjLKz0cx1mMsHR1D9T4fIFrlVdsNfQPf8ksTnj/WvvcYlz1JrNx9fe72OuXyPWhA
vxsSCqu0DgWmSPQ9OK15O4E+uNXvVtPrm74pu1v8tABmqvmkhmpV/4O2lEYFf+OO
PPgvB1JPeU6EBN9lt0w9TAV3Vx2xGhbYkltVRlOBdR4RyDZJ3M/FooZdsUm4ZpJu
AtItksxnrrlDYiSrwS78NKjCxl5EJObkmOjPXibZ/YtT3/FbRqzw+CRa4bIvjvfJ
HeRClyx5Ijq6pjCWyWcfAmFsht7P38yNarWGcVE3p++gn0gIAvthremhCI5YVB1f
ViUXsra6zwRC9/GUoZetH9VZVedovuthMvpafM4GEgE3DUVEG6FviSS8Xbwi7CAX
A8cb+M4o0zGutRKTkGAk94qbQKef4Xvkd4TvjAI2B65++mzJP1hNI5pCjU3uyiEL
wS81Srln1Eszkim6TWgg0/sIbF4RqJEZpRKNmUbE0qIyz+6v05jCyiGdFqiB7FCn
jPxgqIsBFkW6Hp3Grid8QPX7I+oVA1XgVzG5AtuoGhUF7mLeZlpuoeHIOfm5Hk2z
UE1GjX7B7Zh4jsu6k+DUpXKItIT8TqxZsUO5vzAgaQPUkLJkcB3fUsASZdasO7j5
tVzN93Sb4wRnx2WynVzGdEbElRCv/6Rjgz8EwdP7y95mIFL8PBpL0efxpWVE7Auy
Qi8X/aFRTNK2vK8BRcJMpdAbmowLDYuJt0+3WTYBRvfy/N5Y483pSqlOD1CT9HQg
RsynOYLUY/HOnDh4B27aIOOTLcSyBxaK8PQhwzkH/GacMUceSIE51wgBDfzxKjvu
+esdZp3y/8XiHNCGb/0/wB+wehZgFlVNNgj7+jMnza5tF8qiWqmprmYNz6n43lwZ
hSmbYsnXRaHdeBx2QREhQ9/xg88RiwBVbO+sWl/WrhDUUwQn+110xTtJrpyGtWRR
wY8YmjBZxTTqBCqDDreqZyYVJ6xblhKVaXMSDMj7BEEszLaWREB2eF1tiGXEa830
VHlz4AlqsLdb1OJx8rojkC0NkmvNjyLZnFXN3RV0GLPQ7oQduAZ/w2NFCZwC5VNv
nuClLcbdBW6/Uid5RX+5iObUcXZ78KqX07JfyujVHBaljrUxQRT5ZJH8BIAwQp1X
CMpt5cEDhH7XjmazRy1LtoKHHwS0izlQIcEALfbd0YPebafZJUwPdA7f2PyKNW1j
hzyvIzTfbUKsnKrju1EerxvcRdFimQg1w0cv57dfbzFxVdcsHZoFgru8J6IVhPBw
1BPQqEans+2DuDbl3JlToDxagLrZn3hmcvcoYZPbeXM0CLFlSMstQ9lvMdMGRSOG
Dtt40Ro/Nm0Fb7Rnpf33triyGswBUtkMLJHYVMVrIFC3lOVl4WPbLWXDnCPl8e2z
kuVQqCUocBzqpis9i8CcX62tY3OrDOcXhqjwrsspwHcqP+2qdasDQWaCskApjfaD
CNfO8pJAnUTXSUxmXu0O3X51LuUm/hQSJLYSzUM+5jvEzSwdqIbqhii4aIlTVZ+c
uzkrEsqOB+gk0eeCsk9gH+suff8G4GOsXgUrvn/GjgFeVDDwBOe+q5/MOcr2+Y6r
sa6rfZ/JKxYNufaX47xZjKFMzlPppcesVTXYbNZWy9ILuJbCaYFFqAqSbDdPLKee
ffo0SVc5YTw/zSwHkQeVrVe0jtZ1pmDwPPheAAJCVAlL8cMpEkKZ/j6eALMaAW/K
KYgkiu4qjbn6DEfly0hJ6/Kp2esfZWelgVbpNVnY58mD4l44GO3j00lu7T1pLyAz
EC7Gz3VEoMfBRCqiL21o/ByeohvPRBTqhAZBylW7KkcyaQfxvCw1bOfA1okot2eq
uTqCrXEj+LgE6xCwcydJAAZXHo9kYew95Aj0zY47nmxUIHBrolXCHnG31ZwIa01/
Fo6WQ+xwO51I1fFZHJYFEK/j+STP1wdCYw/TfgXC3i9lHnOaAKWfE8K19kLMvWdq
Nnc+clPqiZ2hf/hrL3XLlz4MLTB/nqW3NtF3Rc+mCQEeNjneLCkjGz6RMvG4H9pZ
6gOoc6NTW8mHm4cUKGHeJfsHEoE60aDOfyGPtb11G72uL3+J7mRC9tUs96H7E7IK
khCAaXRYCOxtiapWauzDXGy6pxttVOY0/BqnxDS2YrTNUk0Kr9/QnJaIxS/y0HKN
Ro+N7Tna5FCMh3tCOmUNWHw45gv5j+yV/vAD+GRm2MNUYNOOJN14bpJF8crWtCLm
TJpqrkzxPi6uxO790L5RIgnmF057QptH6aleu7HqB/i2xsiy18BlzRpME17sKxXJ
sEWv03JW3/Ybbg1ZL0cKBUfK+W7GoR+oi83zWCCgVV5oBkOf+PHhejgNYlG/q5VL
tYYJ3dXJIUIojFqNkCzgUfZxPHCJ0wV0jZhU8kVt1GWfrFmbRD5WTkoOWzz4fJbl
1JlmTOEUOhcuuexO1QsAZA67ugpLQ7FHUoEDVoGmJCkejl7xnwA7RaLFed49VsPl
EMv2MbXxmEUMwx0dYyVyBLZxJWyovGfY1ttWpeVlgW8RtDYFIYXfGHfuzStbVeqf
Ysh2Q9j4Jat9DZedBkYWOwdINCqytgnzqDTNs3I7p9lLMSuTs5fhHOu8j82HsIeA
V7NVvosAiljYfck0Xg/KHUNxTZk+LknWdhXfdxKuaIPeKg669L/MH0fdwpYt+tUe
6ZKTKYvOCSDDmlnVoXZuFzceG/e6X7+vAJ8hQrnuVoe7mFrah8PFTGQZiaRisBEy
TyNQeDQZoAU5AjeaIHVQnyJTE9c5xHTT6y/+Wl0R4huR/qRFA88MBGmaYgafLrOF
9n8PrjBNpRmlarfzp4+wd+A0dbuKkW56fWtCwx3MpO4inStnOZLfbgqbKp9n6AqP
iCC8DSxbynbCq23V0FeWxnKpZc2seg3LV05dng/rYbN4ciQt7oMkP/8ifiaWrFI4
lNSzEi/DCuanteRxk7jCNL5IX+CW6kwe1u4jjdJ8R8LfsNaL010uMw4qbG12CL19
2aSwDkbs1G9D32cff3zZJj/iiQ9kIw7XMAYwCS4kl+Ta/HGQkD93Sl17/ds143ts
7QDr4N2mebvOZq0uFZQf6fftK4wwWtWLx/1tAgkcoKxb8NP5c7RBedMJ7JIc1Yg+
+ZyTi83YblJUlzT/tIxSwPuxHVyJYB1TgF48zssGO0G1FqoKWClwKtxUOieUf/Mo
GZCzPEHxbvD7VmBEdYxoTE0nVLdwoGQHfkm4LZY3dFepwEHYhEtZTp9xY3dJGIgg
ooCYZNdMfalxJbLc2Vxtf0hELMmrtpi02a31j7fXp2QsRm0LOyCUcjptrxtJqt5D
S2H9CQJfAW479EbOjIDeA7mxKcfzDehT5Kkr3Awyg7Eqmr4s2/on1MmUv30/O80d
7x4nzbnlRWcgN5zOomT6z1ePKxOxFCIClS+9BhHwi9vIxzGf7rY7u4wmX5jbRnxR
uWS/z+Sh6xcLMZE2b+UiBOn9ea+UW6ImFFwfZ1NnQoPMlPsgV3qcESIuGHFv5ygW
ksT/W4+33qHiLJdM5q8EITp85FnE7ojnr3lF0QWb+BDzqrTSZlAWIIva62hQywBU
cMcIHT2nIRVcatSBWQCuOXmvYTJ66CPhud27aJBJ4zMMn/QGiO/42CCHuFHQZR0d
sCGvhMLMobIRRoz0lly4Aqo1HPtunSS/ara1QJS3GNONj5blHvRaXcsNTTvBj16q
CuCYTwUTEVcP3RtUjbK+tO/J6TbH+NMbZfYafxkDLM47kvGkCqQmob4+xRT3gU3r
T6ON3fHscLezdvgOBiekt+OCGODAVTie+gNg99aWwqdQw5+zvE4fEr7Mv6BATCCq
rBdYAt4o2hG/DMAYa5ahMlvmJXJJOlFFa7fY7YsguBUqHCFm6+zipQeNQGR2xPr4
PINdgWHndHhtNOt3R9tUULSfdjPncnqqQq3BkBNZLok2rfgYpxPrqAFYLbKa6o4E
xCQm9qNrTyoY0LKDVA8bjLjYSNoVFkOufFJ5WT9gyF/V0Ibw0pOximwI7hruUQuW
yqNzHtCe4NiJeUUW4hd+0UjCtDKHb8E1ldHU2dXgv+agd5y4rNW8HboYpX3J9grI
Rk5bH240k6afjsh7TJb2D5Y8ILyWmv0PzbwYRroRDIHUMrVQA4P+qHmjQYG4dI3n
Vg+DXucKh8yDza/mYx396F7+vCovCvQxAeaQTp/s7+ndwPCHKfQBgniI7mU10wzz
8dwv+Xy8B7GzIBixC/Nz3wbfNv6eNod8PTf/whsGseuz8f/Do9HtaCPQ+uClMVIk
/j17BSLTaaEP1NJN+tFbW6Kkg/1Wf/87MfQx6czbmhcCudrvCiTGkZjWXc/lQJ03
5tdgZgHLq/cdylhcxgeNuXZOhLBjNwixpnwRHSgX4IMX+PJzkwvhw3rJ1Guu39SP
trshDwmHTgcIvT7Qx6TWiB4HmV6IQU79v/A1NPLR3vqESaZvKhCCW8L/bCv0Pi+e
yYcFqYBs6lHHjwx7mc1DzTNhv50ncJYyOk+zoJM3jeOKYk2cumQxlbEsuq3OXRjc
LI0Omi2VCKmqNG6zVxazD85imwUSDxG7usDUAwEWn12DKtqLgFLFH57YzOJ8Kdn+
to5rIaSpWgWMxOwh1aWF6g4tyyrCJxob7s8CSHTOD8Vvj3x5GWgusw2o9zIVkiMz
nTjyfpZPCCPMLDpnEdv19IvwmpVWitgeOcNCTFnZvICdMYmuXH5Pm2iyg9u2eN+6
OL3Muc+dk6PX2Km+Uw++P3mD9NLp9vbtZOpHKelZkVQQ5tSAy/ZpcLbJSIzv+4VG
BuIRKDjUFUTxj4a8iq49XcYKaghWZcBO+QISqW0QV2us9GHJrK+xWeHaCX5cMzY4
QoxjEEuCY1VJiat7sB+qjiYNBgdAUge0wD0d0BVo2B16i612tZ8J2OGRDPWDI2GD
4cuQNulnb9DBcLc5poeuRz7OXu6LtZiFyGLxKGnOtJW1sforZQSYpbNfQi1Za9nq
2DjWD7NRuyS2S8l07ItZpuWziXiKmX5d5/WjNJGoc6V0WDRoiv3ZN3JzJaTb/rBM
TWrfHgMpg4mvWhjDqJjvCpgia026SchgUfx//k3YBds/njdtnquLx3B/Im2r/qz/
rpF8ambo4D2J9otnNWdGiTHrA9j8D6QziyjrPF5fymftZq1zTdTrwBIYZjiJt3xy
HpDtWUCzpB+wRSwZQk9zsNgcIoRtT3YLLsfD7gy+5ozdwI82NI3Z+EdkXmfIb10s
+zvhHGMNLl7Ez6K/d9iTVEsvEZDsjgamKO63h+P9s0m7HB5Agz41VcHViwS7O1ik
atZFugzuxsZlzrj/DQtDH1oGrBuz1VvZttx/MpLjkLaPWdeanxDfkb7ASpTMXZqF
JHnxThaQKVX5eUamL7mUGQlH9TA+hFT034n+hK5apm2UdZbvRGL7cyJbtswOlSI2
Mb1KhhlpBQ/a+DytCStrTEXAt4mbC3w7lhTY11jW9t5sypjqnimwCfAsmBUQGytt
3qQTODid9q/oatslBGAalFbf23svnebYqXcrAkw7dV3FsZk7KzgmaRgONcYGsQQu
OaMwRJ+KHGKFXS3k2L2epnPVclMLENXUR496SF/92rTeCL5BISQ24SooieoYiLKB
TkQrfZJXj0Rj19KzLWVVw7XhedLkCCbXTN9OcwoiPdpKK2kaeXbJxbA8xHl6wAlG
ST9QgSMn6HCf09Q5rpc/6tcjOLSVmr8oNHWiBAQfxxxnHWHgZLzwjuwd5c3m7D/N
lgAb/l713GRRag4dskuRQUEXl2nWZJQ8oqBCh2ddAaz3c90yN00aZ2cMCvnGaZcA
JNTFyF2+C2ZNR4oPHLCv+9mqGUmC/WsSJAZeIYMstq0DOkNW7x4ikTwtu/IpOyYc
n7lTlVhw7/EhB8SwiE9IqbWHEnusM3vT2s1jMMDOvYOF0WSLZ6B/3QitZxmFGV+Q
rYEa2zO64PUMxMN1+k5UBptxcyZJaVrsTE4jMQoygOwniO/avYowfsAwcbnBW8J1
nxFgXnSa2IbHBbMy3Ant1zdFIvMmEXibKyY0wYiehAIRKjxpKqHDQXz91/jPlgTb
U/FjtGGeLvJI9GTD20U1H6knnHbCksrVX0+j4J8dOwzRD7/3GemZPQZqdGYnUBZL
yaQjwso//e/rmC/LWOGIdxx6miXy2u+VavPtGy3dexS10AIEE1J5UHvrR+SG4tRM
z8gvHn7lIwnfetj6HSGoN7NwmlbvfkF5D5Hhc9vGkFKT33l92RxfoLweESmo901h
6dXUBWrB+RXcKgBy8PKZwXL+t2eDmbZCM/qyynB5jKuhw/jV8PXMc1Y8u8tyTFHe
+WgJKE/4DRsk9salB8t06eOM3E1zyw3yq8GQFGZHl3UQmitJjgiYlDegwEqMn6JP
GF6IpFzEo3vM9Rx3m8///7kLzYCIegRqwMihVUPPaD8E0+IayAW92UrqUtLtrItA
nqvbvd/60BYnABiUeile9dkI1SHxLesV+pOiPIt5fxTW6TvPHwg61vvNcZGOwsHr
8meQ5hWUMbCqrHIN1c8T1XCubyW5ZKk88Qeza2TRZ/04T8JaLNr5PB690MoUvclA
iGnrw24/zOJ2AgxJbbArQMpb32AmgtY4MGlTPVf0MGxxfEhr4y3xPE0s7WR7d0sV
rOl+Gw45dxFTzh7VtX46PIKgAV39NP9AbcV5MJ4MBwc2nX4dAltOEOcz73QhpXvH
a4Hqz4LAFqJEZYbOUpjakj3WAOUayqUMCyTAL5B489vbaI99X8oaDGQBqscxkMDo
mrzg+dxYRS8CCX21NxYtA1QHZ7FPycOOOUvdwxDG/LTffqCnZS+qLQrS9h5mnq2U
K+Jn4nviU7QGeAIfzjAwXW4d/HjdtCxQSKfCVYuERwGne10JFZey2PQFuCRnvbUH
TtJa8O0bpxmy1DsDBqOGiDx5X4aTRMT0g7S+XJy51bddJRj4bYOEDHfIhmGrjQe0
wNdCBBadBP0nBKQjTM+5H6B7iUf/S6eOWQuQ+sUGCzvwzzQk4rWNEwdfNxd1F/4V
9JZkg7RATbZLH6WRPENWfHIEJ9Cu9l0OgcuXUFkcnJcQBSG5h+jyNgyhUiuCW4N5
FI5pQTGYhPdxtACXMWyGlGuYGTBxQxLw1Z2Ips77ErM/3O+Yl3BdQ3DjBfxkvCUC
qY3m+oZO9Zd6jd+TpgWMY87vxl3GBZtHDJHXoe5J5li5xc/dWLmLB0/y+j5DJWaa
XqAQQlYXyLW6pLDjcFv/QlW4gkUGXE4D83ZFSE18gqOA+RGb6xypuyGRyQvdb6AV
S1C9GXdQV+LreH0pB4fcYs5HmvTeN40HPzdDZimFD0ghVID2liOEiNKUL1Uj2U23
TWr1LfZaLZRT/R3QP1OEpCMTVzoBg0k/COoActAV7tq4fLJZikMMzVNEEA8mdjCB
fN+lDwoypADFjYKeFlM6OfUVoMN3cxHPoIPkylW8w2xelY9ocoomYi/Vp9w1Xm5h
CJOK0w/IGQG/at6zit3tD+aTwbUvx1lfqAiaLeeUax7DLFolWTLcRRLaO0lxIHOn
TUIJrzfIOFVi17zo92VgbdJZ8OgPnLfdinCSBf2BSaD50roWvpYH8DY90j6AaLDA
Gm4X/eyULNCDoPKD3GSef9fQ+rXIs/TVj8fdoCPkw9HgF6+bXTSlU4iOUPqMG+j9
yi9bRvRLLxjjnr47pcmLU6/7+8Yj8L2SfyWRbHkKskIBZOfrc5z983b5vh6hFBWg
/ZVQqsHaB/MRXLX6yEVlDtLZIXLk32nxPjPma34iVetGTTKjhM/e+uctb2RMGb6B
ZE2ZIEncQOBEp42ixOJfsny9BezNz1IXIChLfbtQnyTn/1vRhhL1vs7YDyqHCVEa
o/FTznjB1+RoblrgydakNNFu+cjUt78RZDfkpmZtnluIAMsBIvMHlweKvS7pYTta
W04c/bFkabyRPaebv2z5NCAuORcwiU9oxHVVxHfM0uZKUXLMtaqKRbVf8q4OEH0Q
yj5wRIe6yaNlnDR+N1epc4FSCZeTBErDPaf6yd5rp10P2nMtYp5UllOkOpYOnD8v
z6iLpa7iTheHmhhhrFHgl7p3h5H/3xVFjDTf5Vol+320dlxgaxSUgrR22JWgUD4W
vEgsJYtBXYCq32E8vOs8RnBrfn/2ltoeqzxK0MdvIBdV7FT+x+6xVOxgnZxHto4/
SRxVTWxkcvL059glgXMhbXzfmABi2EG6k/WiVU2NsVtiFkuae10+tQuU/Df9EGmU
NJ1w3abTdsDFT96vAgQWIATN40AN4dmkchsRQ8p8NguN5Uf1XfM+iUYHhu09vAbV
lxRo3+Fx8aDDRu3TJyJg0hzBdyjb4d16lLTMixOQ0CgNAtNG36ledUpjVTjUWRbc
BiiCAe4fLbEYeY4xRTrh/wSXdNrUGVM+ryJYlFNPKlhjWgAVuqRamnQzuXX5xcQD
G+qkeIbkcYxAxd1m/CAYKVMRcLg1/0e5Bu0tkaUbjJN/awvIOyZd9A9dH5l5mgDX
YVo7jT8zT72pH5vDjRzrSmVxz/36DTgna9NcEKHmzdZcKKRKedIRMA/QHAkuneZH
waEjdoooYxbD6XIedcKlHgCTH4+yFy3MumqXlTgA4dLAngnDXbciGOaQM0rjhJZg
hZofx3v4t4HKnvTbyt36UslkjeSZEzQ1QyFdkWAQi1okEOziiflTIRM5p42fYxJP
KPGFtsfqwgt7IZH4FWSNWmnAwstRggN0P0ZzbQNlBv2TZegLueMaNAFK9gAMURD/
d7P+xdq5PDpH0TwRytj1PnjpepsGSN9tqnoKAxVMZTddW6TywTml53canVLqP1Wh
ef4/uKkUGdxRCkU0YbMPgacygVaXNJsLM8vXyPoprr4XRoWxPGSFqho1JerabJpM
fSQH4a3LBliz4C4RJWsr+TK9jsnLNWc+LsUhP7IbAqZpN05PaMJcUbMUDG6vG9jF
Rs9rbHZhbGwSdV2zuHKoxahYT/0EHxPhvJH+eSySCiVdxzsQV9ipjwYlbsW7J35c
ajEzuKx1/U6wZ2Nz0QOaRk7qj37JcHPlanZPtsoHw/xmKTmrwqC7rrPigo8fU3jC
6KfAVvrXXvMJFHgrjhufZzffz+yIKFWViRTJsDoRLLTmo5TMHMc1A01dDX/Vox0u
nmjM175Wll8WL4jmuRzR56GNyYUj2iVQi3rDT+i0GvE8ZUPUvFkTkV+wEPhjrFR6
SRjAUmQRESkIRwFlB26smXzjCV2cu9V8wfDEnkKphBMlnUFy7N2jcqGog9Ae/PPf
JSWHsqI4/QJWkvap8l7CK4nTA6+j26b0MPOKSyNWvlXLBSFR8TsZzD/bcH2xLuI8
CKhDwhtVmh+DzkjD8MCEOw9ky6Mr9+JjCrpwLMk1cjzQaRgGuox3riT6ZS31Hgfb
0XMfStNl6DLxF8vrJbvNTAdHxV6d14NBz0xzcvSrfKLs4VDuDgVqSaOM++D4qV6B
iR7PGxaoXc1cfM57WJSS0ra+1icZAtxbpIslqn897Mei19V1HVgmvcTQfWiKyjKR
5BAzo4AYx0R5CLyaY2OD+ysE3sppvDelbahx+RZOc028y5qhi5ZWnnVcMrXk9Rko
vljvhUPGR7oAC0qTi+1+PSy5ep+oS9fk/NdriZVwSwYs2Zed64waRtSXjIXAy9Il
AjdQRjz5u8t9C4Wnd4nx/ZfOPrLvVOwF2a39mP8ZIw416F5iNesud7HsHQqf24b+
bDxB1cPjbRxcfYipSOCaW8Okk6nyg4silG0H0J0kSEFIckfaSJMN7VIhUODyJfBQ
ZP1Hv+Enjv57QV818ib3/ZyjucKzkRQ4FwhY5/InoBh/QLOYyqpeMff+FmqBvI3o
H7xz+7fsJCRgJGGl9p4+nLz2ukySCX6AF4C9qCYNYDq2lNrpuuzhojmnRatHVuqy
nzQlC7D5yyVS2yZ4OMX3a/UUoBrqAqtu8N0PNzV+zeoXn1pa8imNV05DXM3cR+uy
Bv8vkob9hCMv6K2pJA6EiDQ11XSG6xfu+/1JwxjyH+aUYoVes7LH0IzSiYW70Ei+
9gQ+dkh7KEFuthp8MBn3A72QBHFDBjPOnyDRY1ELC10zphwQ/+uYJblTTd2lUQnC
DSi94Gh80sYVUMuu8WEoDFCrPhqDlURC6XCmSaHpccxKwVyl91/hfrHC4/JdK+1U
6F7+CCqgpiP1+Nh4zslq0mcoTDwCyoZJKo9byBwbnNfapFkdw2usSGE73oDJvTS/
DKCrgm0AaVI2FXPyNfTSlWgzTrxYOypURRVFT0tubrokeHaLBfJ5/V6zMOLysuu/
8fP61+4K1nRYIzj+c6lCGH2NIQfqgyBF/lCHNVdYL0l7GJlPcPrN/oETjhMs+SHa
qmvjnhoOZfKmQC88AvsYKVJPGC5M3WMjesBgpCxIpJvpb9cgJfIVdRnb8ma1qyYM
FhEIuFiFjoMt0cWm2w35hR8Noeb+yb+Ss+t9xK8qPNQ2uLC85NA3LZXXqaWStc3q
FM75rxB3lBRdiAr7lcvzhxHgdff7NsQNJmg3HfGC1UW2G1uZFIABmseqTZ+RDQ5e
PEcO7Kn/SQBcK306dCoAWUyko+MKX/oYVPm3uplmxNS3T7v0Qgxg+km0INlCTlCk
YIAOGMGdTx47TNRxfnOzHiRKfPsC+H+VJz251oAhxIqDEw7rIunVSPMvPIO302zP
7bOHHp+ueRx/0/SaCTDXPNdFM7nAGG7anvk/wLm50PJH4lWuV6DZnXTLFtBzeFD8
JgtQWZJ07MyBHhgmaqeEBcuyiZu9dHSRboP7xMLIZDB0I8BwoUVLrOWmnqQwK2mG
6PjfEFTDo+SB0gCLaG5uKViZPUFFcmMOgxuhKtYPVMHTTa7LjFaLG5olKO3ar+lU
vm2NDvVfvxShpSttZLcMUwZihuWe7JO5xav+Kl2+OEE/PRo0Uv1oKsAxN0a35aSo
V3MBq/8DqIKjHnpEtyq0Z0gTNmLT3vIFlTiNvtECfIsO+Qq2naQZXUnMOlocqjSq
b7lkd7OQMxw3y60PtSlqxikMwGCp+fSHLSJSGxLMKT5Dn++7SmYJBg6emxdPai2O
llhhpuM+cYEqsszDVtHpRjWLaXgEBp6V3EwpsR0a0NbRPHnmqMkbXxCBALy7wCUJ
mHEPvbmXkuumvD0/wveiF4Zg6ignudFRDEQdkV+Yn/1yk9PqhL214Zuir4eUmUar
FNr67t5C4v52hPs/hsNoGp1hZWWXkfSScXzkt5Pgvj4+Bu7DTlRwBuur3XpZRsvM
lmOt5z0/vP0N0fj56jkUoAhXfgIFxk06FLUzZ9LcTaN0PlDTI9HFGA4/UvODCE/F
pPm3XC++b6NbeZY/X28Db13d/MXbbwI+qzp0TRSa8oqNYYCQkgxq4XCHiBB/UnHk
v6m7NTQ3BIe7N6NLO01bsojOwH688qXn+aL62Br8R5hWKIN8yXaJQhMtohEAPCcP
RBIYUXy8XLo/B5o4eAmg+nesU88WRB/rNngcJ+P0xxvp38wtRqgAFP4BEP08vX6z
CCpvrsvB7cPNxIWSTvg4qNwdPtZjguqve6eGsunA4DhpoyYKdYLd/sCcZGNQqT1/
qYNQhCqJiI2+p+W8ngFUEfgkrIpoxPKntc78llpjzUI07nGKi/EH/yArJrTcXQFA
oSnQP+0O+TqoMwxN0b667n1MaEmvpkJA56LWaQrXaGwkRZn4FLk9JUl16+SEUA37
wVgYRe5ooqtsH+uI4J2t4G/wGgWgIENuVmBdWwJ0O3G78sxSCh6PL3IZm576iVCo
A/0WfNNIV6S1VcXNPEcT/hnUdrl5aKW1A7hsmuBChxnWTmQ88ct643uXNkmH/2J9
I8zdNv6o4X/t+HUPxYXtlCwMdhpF9NzdiB5nJlyHPzGRqx92hODqvJ19EUimE6Op
ulCU/GvU/UpGmjd2f+rFe1o85l5AIujBnv37XcIcXudTwi+UQ/0Hvp9tMrT33Rt9
aKTPx5WtqZ9KDhY2Ini40ez8k6gdmIbjxYdi2RJbL5ur8In2DXw5gI+4DIBpTP4O
fSamwdCM3oJpd3M+e1ommTKRj/xFL5i/fQYIeSzJx/WrgybE6a/zCrL77cAeB9QX
O/WTWh0IUMMayqvw/dWmcwi4dmhB9Uiy8+xavnFzeev3Zzbei7NvzA05vYrcOI5b
0/MKOH4K09ri48rThzMD8zSkZIXTG1y3Tkw2jWhVIy3c57+uUdvAQK1IjSjlxP9Y
G6Xwzy72eQjC9aIO7iMLqqvrv+qNU7X4zV4x82FfHGbO8i4r5vbaZOfaJzmh+hB4
gzDj4zJE45GCKCXoRD37qMN+vrQ+VB4YGb0yrOiln3koCEMXxGUTdcmDY0lm2RaX
5v/MbUVasV8wgrIv/9Gj8klGKz4vNZ7B2704oWW/B0iNxNjaxx1pPG0MKoiuMk+6
Ulm2mprKoqlbTY2X7/O1g1ZNB8jn3zU4NRMTanSlzCR/PtqpIRiKhirZprRz9iNC
JL0p3xq7kdGmwhVbsbGRrv0dxD4yjM7bSuDNEWmBABAsKq7PiUyki9B1ChV48Qv0
wbgEwDEruiBo/gzHxuzkvsSG5YbQtDHKP9HjOlxZY4dzkmCueQkFPzZbiCNWxsJc
KdVIO07dOVkCEdQOk0L9DYqsveAUwB8B2VZTGA0mbqX5X+Z4PXwTfWT/7tw11T0i
SRHvazujGJzxg4xvoY4lIeTTTCDf6NNeC9RTYvXFLNTapOn9DvfIhxF8T78XECo8
SyXBVDxH8GNSvJ4f6ufQosKJ6+8BuIlUpgGLVY1FT5pg2QK+MAfaDSVMbRdQHW5S
DrIL1Y5rej0JPmZNumyvbjv9ZJVzdSoznT6qIyIY2HIsvt6Hy9Hlt7EbCOvHG+1o
YdI8J9Mgh1efAuANc9C839dGZ83efYSX4ThknDSBJ7tXYjC4De/ix4jHDdhAo9eI
tp7DtmpZ+52mE1DtSXIES6It/8cactJjky1HjMdkV9NgZ7bcoaLvHK8efYo2YxPZ
jFRTu9aPnOWNSZeb0GVmo/SIvYlnX2z9jLrQv9LRWm9FR3YZh2jnHu7crsZDbXID
254y8BVCx3vYVUORtnyVKQgbxrjK9GAY3NKtmxmHFUpLkMm4lXBy8kQdhjrzvetO
gN8X3GDpyxXZHavJ/FicHNVyAuwGX+gDGbcJqny5vA4XpvOQZ+SeRI0ja1iM9zHZ
9DaPHOm4Tu+ULDNNm3FWx2waB5kXrvDZQG5Bbcy6wO4iRsKVqAFPentjo+jVqHzD
H5azAkb68sb6RBlRVheYQStKRE4GlYHyi6qZBec555jiGQE/O1g6WquRnizCgY8S
3nZdat/LkWTiBUstkaiAYTJ2JulyCkf2g14+QY0hCRllccyvvwWCBB52pLbcFe8Q
C1PFqGthhxLeG7bt+w1qakuQfewGfpHCXVYcN5aTeE1DOjApBO/F4/RnOzyRvvwn
dbPtNiWjSeIX1NZkwD7psi3YNg1j/+8UwgTKrG30ih3c5Od7bkXVbAgks9lkjCMg
dBW9NSCNmZipZ/+V4BajbIoYJpI8b9o1eIlpUFWvmDZvtfqkq/P9A4UwMYFoCPyJ
RcrJM1YId/yUwxXM5gebUdDaAh6dr1lG6vdsgZxj6GDkkEz/1gtXBLQlSgfommHi
2aYUUUagSw0sMF/hoNobWMPm9uvTh3jL4UvTkuhUPYJlU3K1BKWvQePwgHcZ+AQC
e40yhK+Gxa4AVLEC1/mOUHzdQHPtkg1eRDR3DHdGWWLBVZLCp3+T+tDNk1i3PvTy
bChx84GDB/PFiDglEsuu/hne8Y1+vKA2qRRC8i3vEf6ux3e+tEsRpBVkj5sF12dQ
B8gOHwFQjULF4krrFV6WSn1Kqm8d2s0//ijH2IzBaFHvabKDnbpKmbAhBX+sBmxs
4suabBpDpClyqKstgTt7ud6xtQ7DpmWpChYZUkVQ8F/8kDNsOiHN/WT27HD5k+Mc
o6j36BaRwssz5+g3lp8IFX6tsVPz6bhN0+ftjFJGllAuntetwNNWpo3EvjZFQupU
5+anINAF89BaYpCNBI84QY3Qst5UbTWcB4wLC6Qvt6E6vzpGWz4F/a7kxyc7ASUL
9vl4ih6N4IOm+5joM3uwPbSYNprcjP3Lb+nARyuf6U1hAdePenPuPV2L4tLErriR
YMrstKdW406KoWRxkX2I9/OxQOxw/rbTf57nTegTYMvH6Key4G3OopmGfwJPpC9E
R97esoLHYK1RD+wx9+Llv5RWrE/YJ2OCHsrl7YEhQRl6Qx+QXLhdz+WQ53E5SbIb
LkK+186g0Fcblk1YdBBSp4iK7TtyRbs6QhmYbkRg4TV1YWyuwKOB+4W7y8iXr29r
bWwPvkKBjLdGliEekiuC3dwgg5ND3DAxIDwmJbIpQ89ei1G+DXvXp0qeviGk8N/6
/GXKhNCOn48fvqEEUqw96bBXyaozBLBsw6Db6sQYsab0iI0diMfaTLPfV5ePlUh9
9p/9K5yyCHde3W5HcivfLT+LBZvdG6rIXAGaQCk9yy6IgnuO+OoUn7ZmLBfFA3fS
4CxI1rJDoPYcIcL6dlFITaM+OhjXtcPzssLCgyLtgliHxICPh1xrCtfMHzvSdTf4
VL4agHiElqEF+W3wWO6+MYy02Ar/ft/9cAwH2ANUeHAJKCYAKW5MYCn6oilESxOe
ZqpLoEBe/JTKH2XT37n3kfB6+soL10Jj+jDhguBf1A9mGus0bLEBempIoP4GMwmj
uKtR8KqSdoN6P7CVkRZaDKjiXIwG5LSr9OVH3dgHlAezvC+jlhLj3zNmh8tfsPil
UGLGxKwgKkP5bH/BhDMBARngz0/gSAdkq2/t1ebnvjgDtXm7CkR0vk3jTxfRl/GG
6AajDL86p7Ei3GddO8w4+jTLlgEWWSazxSD99U9mZu0hscJHAf9vhY0YR2AqA9i+
mf1XSmYrfdBMIzK3esnsi59xLgzk2iMqSR8JeXx8Z6r7sAImV9g+9lZCWC/msuMG
scfhElzWeIbCIPup1Qf1NX9qtcqM6wXlHCxeyqiPRNFnFUYjoOcd5xJOv7ooejLG
Rze9yTSvZ74xX4ziah1x2gQzsCag0lEOGUCQqzWyen4jhIiUmuRxkT8GMd02Bag8
XFRMaBwdPz3OKpAWNLids9TGbjqK2XuEWm7CSgp/t6ILc4rvCg7sH5jamptuWNbD
dZUv2oFRXJrmFJ/7EoNnkw4D3vptYu5Lcf7C+dUFqI3fx8OuEP6Oyp29OQrl8GVN
0IB175xah3TbHqPWv20LprgbMDcgbcNHI+/rahDn8djdMNeromrVXIBU5rl8rXAv
mcmkUq9A2mfXsHLTw7aMbzAZ2jJDL/u1g6/lY6Pnw3CmDL/L8+TNoB1rL19Hq69J
DZFAB3GonmNuLtKAPSsS5FAkbYWjl+QaLVIp1yUIxZOaYqrjNbUFiH2Sc03IzDEO
57yQzwxHBoSF6WlgtG/ewzb3+ugYBS4JvtlI8H2GxoUKim1nuHmqqiFaaNx6Cruk
gH3/P7wbWN7qldOjP9RcFxcVR/3sMuPS4SL9B2PXw+0oCU1Lia83WbcuTS87a2uV
PqHD14vn6N3o67ziNbaGp7XqyRok26sbilAdYbl7LHAxVB52KDKV1uJ0xj6pGBnD
MfKpa9+v9L4B8/P46bOSF997AIKG966y79kNJvfzeoeLt62gnInbKtgAJRnOZlzP
WpPJG0wfP7gT6ewbX559uJH8wFvkMhTATYl0wWE6NoffPYjEy+azJODhD5Bq634F
VWqWilFNYjIYF7IcVkMpGif9EVWpVRz095PGeeCfqSCxxhO7NVsaqkUfxqJHLNOK
RHd3fIShAPltSPhlWunMoW5cPzy+822c9hQhrW7U0i3Z2Z1KTyHtufA/huNf1DUX
deJqIppoXDfZyNI38ugQUP4o32RczOPoyz8+4n8CZYeLLnQpywZJgqZI25rJDtQQ
HBTMuZynxq/0Bkmje074P5HqCweJDz6nOsxPjaS8GAM3lUHlBI9o8HbPK3Dt8gRe
DchuzX0rvBAZW6xyhrEFqVv12nmiKjh7xEtyXuHYI3J9ViM0tJlnNVTbW0foj7jw
TI1aSuFW59uuPrAuZ//2JcrBlF/E3yF9c1FeZVcFwv24xTvfqa1rP5rBc8kpHQKA
B17+xd9/HLp0y9zay+bDA0IduZ3vJjzj97ZrdeD1fGyKAv2mDSZMdCo0m97SaTd+
5+Ucm2b92xvXmyxPTgPL392nSu68RNA3ZtNGoGesrUbpot575dbzqio7dgDJsMpv
m7aSSuite+BQ2IVDnkEwC+EMhdoDQ50NTtH6TcFzFw0YN1hTesah4RqUSaMadtpn
T+DiyAwVV1C0lDZYph1beLIbA9BJl2z3fcKgaoN3E7OrdPmWWLsoJ4PM13jVPt7H
0r0zT8Q6mtnD5bW398FHLlr7UBxOUSrR3T6hlIb2zbbIEIfzVFGxjmgqYKz9IAK6
kNrEdZQEvbQbJ0zVe+xbucntGkIC5ovuWW3T6g28/px18H4gzfa84mS6F39K+nBE
KREoaBbAhc6dGJ8FTuEo6p2OOypzhHPSLtGK5k+VxYk2shVGwWBzH0B9HzF2PQyn
RyHumPRy51Unprm8RDaUdcBIt5Y8cIkwW5YKikhXEByGIEzod3oo9y/5i2Nu91Ea
EAgsxhX9f3tC4eMGLEz5oBQT8LokHThheuPJ1HM5E7sSVuYAgUzn/i915qe2bbOA
PPQIQL4Er6yU3d5DoP3VCTiN9x8viC/uS+WUrBsiZwX6+WiLVsllKxkhvwu3Z19M
UjaLnJecaJS1VaufU5OnneMDX43YbCv0Ouca+/LP2QqNLJN6v2T731C07IqgquDI
/x2YBqcXmAo4NT8K2rl0hYv+Z8GLLcpEKcpkjPIb0NJC9jdBwJDV+2caFXA4HGiA
mBooZuDc0VBHsCtJusX7KlIhPTNlGO/nyfPVk9NdlKbQyC3kchpp4YaWIvAvuVAn
bvCQ+PgKSNIBUPhf+mQXK49B6Q0Pusml652wtQQ1jdOioWbKCI1HILatngB1h8v7
zrbv4xY73WSp8OzZQIGFI5ol/4orUGoVZhX212qaMd0ZAzxKX+MMdA+Xv3S+MKYb
+MGnG5h1OEO02y7PCCsw99JMoa4M0+Loo42Net09G9ThIKsNBYUSuMgkAqohL7iw
rXTxqejbahCIZa3DX3PAqNbsreozclaXPbsi837gb9F8zsWqzQI5kwLJlmkni/eZ
HJ4sFK3QSP+p8c11od7qZ8A38aK0USqB5Cu9HwsvB0gFElHz3RzNHyLUfesLcv8h
352IgtKnyYBpNxftpRILDUY/UzDeN9Wn5gFGCegR4Krv36wiO4xmaBXW96StynMu
SR8T9PdzrEUIWPq7/K9oJmFTKw+IKBIbkiP3NlvbRDJsx7xqInzUnosGCUGXPh30
3zqUqrf/PslNTbccBT12wE5MVYQ0PlQZIphN2sVGyoTtCkSr9P+GUDQtVBH+WwnJ
GN2ixNVRvro0TnssPFf8fgS0kjsiCb+ib0scDxa8+m6sOmgwKD/mT3ZNa2h6dP5F
jYeoxk9xwv+4BdQeQt9aYCRlEm8Uejd63ep8knc3E1Iw4ZJMgDVvtV2a6chg7ULZ
cweGEVTDzvqM/htIIFP3VLAxhHk9Dp40Q+jM1iIKm2Qs91bS8eO/G4ZUqRc/392M
uP59UvXsG3jcajY+cwOxyfFFeJtxpjljFyC6GGZFIlDVuSTmRGBzbD/Ygv3mfjv+
tXWP3zyRCbG5486l/pI9sQIKldTfTOa9EK4VJaWUz2IlrNglSip9b6zNO2yGkhni
Gmwrxiz7wAMdrPmpwAHIWHvEhk+HazFVoED68XoyJ69bFXleuf4ksP+pm+g8mPBQ
1Xkl2qq8IJMKYPO6fUugDhudQaY+df8lAom+F69iHTAcR28LxWBsRPekQrWRENtS
uxf+40SPby/+pwPpnqMmiew/J+RJz/EZ4aWhVAXLYYLprUY7Zw5C/Br2KqQSE9pu
HxaRqe01g8z5TUvsJ4bhpIK6lsRYVx+O5GSS+rTAK3sg0PkG64dK6sJlHWmqOMqO
KYrMLNjVtk0LQyGnLuVZL4bgpBOuHg/FJhS48fr9wj6MdNGLgodn7bzMs+Hj/NHB
cXfCgJtnlRlfpRytxZrQwJ9yfn4hgy7aeox7IkiekAsxQYTqErD7eIUFuTeX9KH5
X84FrQjFNK+8wHvF5OksIf4aXIxJSIht6eVRZjB0ct4Iw7RDYZ84Yh9QvZEUqL5u
q77SksLey9lpS27Eq48h7awDqB5H16a+vAsVCy8lqj9T1by8/UdTkZyBawD5sXeS
BQnDoo1Zqgz0amEIvKmub/JpeMufLmrWVL0lysnNM2QmUW2/84oNPuyUxoavrtcA
pOP9cfXx8C4eDPGWKmA+/AGSEIZkytZVeAva4CY9oru0UOCCo4EzvG44GBZY055/
u+09K7865X14DnH86HGppn/sk7G848szv6D54sJYDNosPRFFA5EqoZ8h34WZjofR
CIiA6w/fPon9V5nqwpTRcHOM1PdIJ4gdhF8xAJJf5CcTLJK0ZysZCTt4I7kLFTnS
XmvZadNn6NI3fP/4qQtxzjv92u1Iibyj3nLSLiCBnIgAQlP1pot31Jam0EGdMdk2
XZRzeeTMug5cJQ67EKnVHaYXeuOt+96KdD+MLMcOb+66nKH8WZai0GYW22iStTRv
LDx3V75MKjDovMhVgxlibEwt/GVNmltHUp05/hbX0MNjJZS4EPBO4VU94OLP7tDa
iDufoeLGKObGToMEYa6eQn9t6EI8oe3D+P5fBe+F4ZvzDObkmsnLkmCi9oxyarhO
q0dWC6ytn4gneq7aQEhHhFFjDIPZWmz9l4H1EtU+lFIug0VLN10b7wG/3O84IqK1
f/eF2zxpgYYYFyJtGkttG44wHbE2LW6GLbaKTvWu/eWLhQLUVNyY+VL1D1UhylCr
2SrDkinZbG1uEQplF2MUVxtyElxLj9oFu1wGj76DU5CRloQzCCWYh9w8gB2RToN8
mA0xWJjmwZVvZygE1v7Insy6go0/IaNjlQbNMOcwddhxFKpKEgOG8JZ1ActSnddD
YqDA5CsKDX4p979vpvh991oTRwxVPz6NNv1m3H6cvsPk4oLaEP0KCjuTQAGan59X
KlIQyPCYgTrsxCaUbLgVSHecKG/bQ6R/mUT5zUKQyFV9uyCsDv/GnUt0JtoUc1hV
YdT87Kj01V77tH1J8iuU/3adKzu0GW1h+Tg6uML98qYBIEUOVnZuK+b/SaQmKFOa
OGoO3Lajjvn3XcrQL63NK7ro34gAYRnbKrxU9sO1g77qf3jRZeca1+F1HuimpT84
NiVLjdA6Asd44FS8GXohvBx5vYq++tmY0rglWJ5mCGbBxXV6G8xGMGC93G9nWJ4X
egaJNiSvP8NpNvzkadinJlecmID+wwnvWVpm702g3NpeuXXCoV7/bW1SFr/T3uGT
3EigtTSJRbCAXnMXp0o9g24YuueiiOpmELDpcM0HAJUVm8JaIZF94DrZBjuUupwj
2pofQeiSt1VpPbxXKMhSLA27wBksEgU/de+T4gl4kmmzFki+m5F8TnOTCx9ZJtHR
MRvZ9Dtgbxw1vGJvi7LL/gt8fZVeC5Ivfm96xiXCWKXY3hFopxHZ003fkqS0P37l
R7JMl+bLir8ri1VFBA3pVR0Pb1L3FOUnGzqGBYPTis98SGTcEhdgv6tFtx6MfPvy
nf/vCoF3OD3GyA0KY4GCv5cgxo8yIUTe7LLtRTPOYQ7T4G/kFytyfVjNmlQ+FY8c
rvIf882klZyHBlSuWtd13pRWf+b7PXm31MrrHCBnlYfhvDYfAHnskoErmhe/Pnek
bkJkX7EZYMgY4hh/N8/KtqevEnmcR7m24bKBpxU11HKwvn+zOUibLPJtVvRZESK/
+Gx//q1eBR4jCoAIY1EvvwJ44bmJAKvcZe/hO0Sdob7avr5WUiMmJWZU1dy4bf/6
tv0rRETBgJk6FGAFjpaJR5Wa5UG3PMI3MApDYgcVCC/bt6A5AIOHEm/SbKsCzcHm
ErS7KyAsEvMPq4IAyUVPtbMSc6jUMSu2/utkldljH6LldEfCM2ltWO82aHKR8ZOS
JRpgzd3Lz7obCsA60eqY3xtTu1pE03uJ/ZDGTNM8cxGN9x/ODjYIcpPxF8f0qJ0D
cS3ila8f8TzXC5QQ1tEbhKlIq/Ar3EOPnzvvwDwvRw9Kn1hteaDq5WrOSsebKD50
t2qK9kDImDbnFBZBLKCZ7bmonRxalIM0Cq0VKtUncpnsbS2BOPeMRlw3vzM+4zkV
Pi5OG+avodp+iHx8d2llrKaQQSDIob//DRiWy53VmRJFXvlmM2bsEq4RFuP772xb
/PDo8CoS0IWX/dOheemUqT3BvWUgEPEDYYf6a/J9c6LWsnKdEsncZg24YH7DHLrp
lcHjXCBdbKf6szZqtL0ErNU3Z2ZlisrLNFan6rHRjZK/KzfIgWu9nYVvIQXyxsB1
1mGsPUqx68GE44wPFHVHe/bYnHt5LBq/wXBe46gjYQddfOF7ri3i92uJCZRdPyp4
dCl2iQqhg2mQkI2CrJrjW7IRsAK0Dl1ZRwaadpfCC06CJ7zA1O8GaHztrwiBoTc3
iYdZ8df7//rhsvMHitqupSPqWd67bhwJl/m2+1SItP71EzvBxp5xMPboHC0U/ge1
K+BZ/5i2lCUPV+DYxraw7KwmuhfMSbe1hoognHiQdOIibp/gWaT/QbFcqBsnju4D
UGrPLA2gcHjD0uX5fjUkaK/A5DEvOF/Cq4dwrYjTGLwWbLawCNVQsMv2NKTO2T2y
8g+aCHvBmxZB+wbqJYbM/X7u45YoWyrUcZJods0vs1isbtAsy+uOsHVfbJGqOwmv
oisHkkvb/xoatcv1BJDwdmu8afYTGYc2F7+zdzYJbUMSfdgmKtrwQIoQ3q+Oi63Q
WJU9t2hABI2EcIxtkSPqLERg+z0r5+YMQ0DhJEb0AG/C2hFjIQSrcMdT5WyhkVqF
2+PubSxjet3yes1k/B/EqhA9+v5nr5XZoGVBoRsldX4knQ36CR3agShA3XYRSZLw
6pm/EkXtW0ReBbyLdtJAHhLaI7f6mCmHE4BYvzmq5AjzkkgnHJbX6jT0O8Gaoa29
jskef3c6r6EDcFs9JC86U3nlWkK6Xgd/YCuuoCkJSpB6l2TTUPl+6AUCShlpLM3i
WVis99rllmIuI20RFKn/+YF02pLwFv43ySYvEVsv9Uj7RSMLMKEmnMZ7jj87b/R9
/lGyn106AoMzcnx6MXUUwd0LArDEki7CG8SphwnRzVBwbA4gEwAtmNenEh5hYb7w
WWhNTcX4eu08Wiw5F5LLyrzDgGkTGjcPbX8bdaQKxIw5OZwEkXL6uyDHIh+lyE0W
+N6iOxqCWVj9QiTqUyQfmMYVqfD+vGDlkcm3iA8Q3M+5azuwhJPu1adPhVD+1GB4
eH9wemJyvaxQwNF2LY1VzgJNvAEkaaBwiNaiE/0Wy02E5FnNnVdzHXb0pAz8v6Fn
k4vBGCVBJdKJz7c8rgo3mWuXNM+XVWRFg4xAssya4OdBd+S3VUb8od0MJLcj4cSl
EBppwCuVHb7F3wAdgQAy7aDrRpp0MJaCk1wjurQRNqt2bBJ+DVYHf2Dyk1fqPizV
hVfEqPnAEAPqImZPzswGeSLmAwypccTsufZNxoseyo0=
`pragma protect end_protected
