// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aiuMp5/t5cCemhyc07IBarVoaOs71QWFPrXvo00vBkGv5BWTqVE8KH3cslHmZPYC
XxXl5pyJoL8lKn6gWD7lmzO2i6Ur5dDEE7Uk5cofEF21FE3PMycZNYKG5e9rn0X0
c8Fq5YkIuU6gumDv+87r6j3IdYUx7yDzqX3O1D6ulkw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31936)
O1NkdBd8iRgmHYkTkEHYDxq+DNGJbHqfA9+F1NcMdPT5vtT5G1VixhyvGFzjis/3
rQuF2fROq+/SSDFH1lQMtC1DcJunQiIf86l0UCEPr6lWBw8v1KXxCSlv9gWkdsF8
Mv3SmDK4Yhuq/zwZtrQbuZVQxbbSqeD+C+31VFf25QYg0XkYJSI0367f5w12fU6L
vhpLwTtQUzQ0+opY+c0IQVwOnO7PnIaFx71k0vFVYwjVIJoN5UssKN3tXVcmHzO5
LCEi6vL7Yw6L3wBJfIIGD33IZg9rEUderOg8jBPh23SMpGXg7uxTYuhlYNzIushz
Arh9vi5L25acnDVU6tjUkRZ9XBXvokv/5MjrhrCGPqe88RcAAWaWfUfzpLbnVTM7
y9So2XXBi/aUln9xX98JDQFa1lZpdxIWHUybPIxbJfNd4P548b1fG+8IO/SH9dae
fRflBjQjqFLDcXs8n0MgACV/B38X9auBIekfSZHUldUy7UrHdJfzRz/6BxLwp1+C
/SOIpmGXmCSUBL6AoaXXF8ueV+WqwL5qqCg0fAROR5j+gvCth427LmpqLbThRBQb
arM5FJ6lrDmxTeBbE4D51nY+b5bxr3JgvbSn7qLVkSdsfXYfVaHfKtbKZhS2SNf6
pDM8wS33jm+vu4WOchQI6mZlPVYzkKt2z9YYKyCNAVM8WQV/7B74/XzdVhZ26TK9
S7OijsjtrPiyhprcGeixnqVmMwWMHn7uG4P7EMiKT86Q6DcQ+TUzGG51ytzNhO8s
d4Rym20N9N+eBaWBu1uwhJb6i9+RLr8K3mWoZoPvgWAifBAMi3Wj5l1MDnkc7qHq
kjzigxZCj2BzJh7GXwA9K1wMnmyXy6jsgcAfy3itJizHDqae5USqbmrdvssYTQAn
E9Cq5ALUGqo9jE156iCezl3fSKOnbx4iJm6be0Cz1OWQzxzwOzR5NjAtgR7vjG8B
oTl/zyfAvU+1sq+/26thfiKmiF4qvXQZp4x6Syf7UzEDF00pIhbB8NajtZvB4LCW
jiSZvmWewl8HyirTW4qKeZE/Ba8f+6PerpSftRSBQWcHxfF7GsFqY1pN5Xii+wet
1r+GhV+/NQi3TyxeXDZpL5B9PCf5aFc2nG2+3Sru+g5khfBWI3p4kSq4cbK0hQ+F
bB7kmw26RoW8g44z4iM65CrC8fUaRY0CyBXVi9BSQB7TqlNxIQv/E2XY0aeKIxIs
pxNBty3fLav7ShddNtPfmYBmq0dp+/OTID8ITP7tts8gFjvcuJ2CHMh58dIB9Xif
FgGAsZfpi/4TU5XqR23nFi9BaRMYaRlXKg3CcN22k47o5pdNnUdI0Vp5+GZ854Eu
TR9LLyd9RNQszbCXbqlhuPE3VlZK6Z92vIjAFelikNxk1YG3KzO58KBA24uvh8dt
QTc/auXgLq+o/c81egh+gUoOzKJYgqzezOKJw3COUNBXoCj7Ku9Q9zG9GnmSAP9f
CsPjCRz5e1Z7FYjPIEdUXMI/z9qmpnU42MOVhhJnWLiFhruD2Cb14LhPxgCfUFOf
USGW9yY9jPxBD+SaFvHEKG3XOWk6jWWWDQdMlTZFkntU8wrHF56awEjMgoAO3Kep
qdA/D6vXdbsmsxX5xma6+JnrejXaGjvV5kKAIzWcejx9NFdeHslFouwOXKJa9X9y
6aTKj8Hv8vef2GnBSFIyrFOa8X+3FhCyBh9t+fLTt54iYyrClpn9+tC1ZBcq5ZA8
3rEQC4OD456UBut1LSrhvBNxKeeaQwSVRQn3irEHTEVWzk/nnaUcwZ4pDZAP/Nwc
FBPOOCU0qluyt7azQqkj6/KyclqouMHLi2P9TOQ3y/GB3uZxxKI0Sqk/P8vUqZgO
eq74Dw0+pSRuEE0bnJFeoYxqtNRWxqPqw3fRP+Vzcp3m1evoak17zcXsGDBEnWGS
5X2PAiAcWNMt9Ov8tAolz80qrI55AwMXk8SJ546aE6ryrpPSVZx1Id8tktyJNaVw
rb9nmBVDbeB2WIoZtWK7EjqtAXbpKPnZVLVAA3vQcBzFPKQCEnXn1nR4FHzu/he3
0XocBPv45lxnpyWYOwwfAHRe2pz3o0ctdxsHmfWCECp8JwriptuFyptNv0ZFx2fM
61sIjKvTCCK0tyI4UbxMJzRof5NtwFOqlDt5zYw5qVoK7T3STH6pzu0QOl8wt4PT
zYqeSZA90kCWyonKAp8Rf1SpJ7hdX+4otlc/oHucYHT7apPnFWRtZ3KlcrII9VMo
3+0H6aIXW+xzDgscvoVDLQaweIr4gTOIBdLtscCfU5Q/G0YTN/kcupSAe996hhFR
NCf1ME+zecCKBfZCJiWNL/wUmLYUhcO0koR2GkELuUmaOhHUHGeD/wNaFMeNvg6Z
TDcV9f5H1poWk4HY2aZ57Nyfln6d+3nrYYJdzZ9/mjoyui+UPknR3cIEVAQ4pFYN
YTNvADzCGW6liAGHi9ViPhtkBHkIsn4t6k/edGmmmCzttK5DESD4dB64hK34Ez7d
RZ/qExdAgNxZlWnYgryRUgzA7jxQGobVue1IMX5VCy3M2cd9BTX21erTltHP1iQS
7SGbw3UlQpPLLR37w+eEYygQ+Lmh3LJ4DJ1ACh4iH5zdCuhO7ZWIsW+04t71ephz
z2B7M/x9cJFixCsU0F+DwX5GuaRBwcPhoNRNZVATcrVZ6NhSRIWT2vfmUT3ompD4
aFBhP8l2yjCfdim22BnZzb+AV7YynHBn02ZaaGbyRslk5kDY4pOXoumQtyXh8XnH
WtV/z2snx8j7UT9fPTq/j7Q/A89KCP0Kvy912uVDghXg7oyLvIS5jLCaJwJauc6Z
XXAQB18SErArcEJBtQ6RecfbLVjx7HP8up8EQmkBpiq0yW9RfiILCdZ39BtK8qy0
wsGyo4GUUt3WgUiFOz2Rhf0I3lhbw9aEEqzfx9RcpME25pJuQoI0faQ5G/aABYh3
UH0UyOm91kTgUTivBWmbHiVuAIzGaxtFxhiGhuyH+HODOr/WRlnC7iMx8F70rXGp
YY+cG0HKHjn+MXW2APXpl+yju9RZXBA2ARrJ/Wi1xmNQWwoXTP3Qf+n4CUZDZVUV
uwLbccaruy55S5jQa7d14EBQkJZ+Sc7SDteepu9jq3AAXXVj4nyYlrBN6oDEW1Fj
mwRz4S0mhWFChiquszKnVG6nt56+PJs9Piu+8yZQAlGblMwh0ZqZCXGJkOCefCe5
JZQWvT1jl53n0xi0/ZxqtjhtubyPfn/t2QGe5Kv8cez8xDoAgrI5q9X6tzSOyvj7
flArRU0An6af4vXtY7dsn7X4rum1+O8uhdMZPRv2cD/+TaeDw+5Oev+czM7ZwLHx
h1ovoMixw/VhMQ+oeKF54d6NYpvkhIDxx0S3gTLYWUbv0RODcXQMj96Z10L8TSs6
iP9+7QBpRlDvQi6fS30HV2NoO/FuDewajV132SjVGf/K33CiSk2zas7Pts7u8+9C
8oOmxnYdzJHVr9roQ+KTRzyen74ZwaiFrEPoi3OOaOOiEcKiBmIUv059yOedzE9A
pmarIhBggH3KOVTjHktpwr85wDLSUIf+jcHmIVw5nvWsc4USca1Kva0+Dqxo6Ya6
QJuoSrtah3R/j0R+2YNA/Oaproyb+ODLdQbPi+P8OETunNbU9Fn91iOIAjmf9n6a
SDkPEBn6M4YALUtC9NwabN6bhtcKlRgeGAi21Qs/6xvVJcLmyBES/QEwCuR5zSpo
T1L42XIudZkhcQGBlSjotR8WCHw2GzWEQtJdt72YOv5fNhZQOgNkgTcTD/puML91
n+4+UUypVfR4iPGLGt5lMrFblr3tyYbXsx2wT8PEcfT1XFcOv9sQj7SUpzxKg+Ex
WysdAtg9LVnO+FqJgi3qz3eifiXFar4UccXm3o4J96jGgTkHKLzhmjBCvfqYh5e9
9ePymAqo6WB4MRGAn41f5cU0zx4UMlSNqTNurUJascMgmlN53yAlVmn2d/vBtWKY
ZDETD0gk62ZvFyk5QnWAMuiTDeQuiX3pPyAZbijiAaUZL8/Ajf/ONhUFHeJbMNWD
TJWdG94KIJQjJMqZkygQYCZtOWxrNnCtyijCy0cngoq6oLiB9R5afaUGPHG6X6N0
CWppA0Foj1TGIsHtosAohDY4ZpbNg71Rgi2hk74Uw5okPHC2jjvgdt3aeRlQQDzX
dqexqYx4WLQ7ECLfn/IrWeXSExuE9/psGS78A15gTHvkT+xpEszZlmYgImh2Xwl9
vatdYyHSKPjt50p/r+cGCOOb/tqXAXUDcMouMpihOXf51Zf+H8Eud48fqrCWvmAf
QmlUfCBV8yjTR0BZK+wOC2kGZ8ow0zBDm2L2f9zUbz2qhuoJvLJz1X2PWrTuy6Lc
CDlUprMG8QenHdVRFQTj35+lRbkUQnUcXeTJucrTS73dshdGeMAuFVmSwSJoLGSi
hYuYj779A56BesMMRfxrn/95WN9klcGckpV5+adv5Tv+l/SnbjgzT7EcqyZ/7o/2
CxWGNH4HspoqkDG9v2xrWN73j3ytOIfFykGZO/jg7kSWjzU91pbO00rIeiB+x/bw
mQLHdPwgJ4/ZWzIH0YfsJYOd77OFRdV481zOlMENrEESJ2GGo84YwOcyGZVr/Ds8
jhU9EVoDnymcwwGGqgcsgDpQ5WzEuspU5JVbEIPW+Ig84isnbIhoeYEJWAWbZ5z6
0smJDkhomEjZfWdsnPS17pdyuxFq3k13U56ZK2qL7qs/JbC2wvx0lL5+KurLlGZz
kTj0LNramd+mWmkIUkqDlcd+9mYTBot2KHWi+K+tm4ez012sYFfbXWC0aAbOcIwr
Chw1mubD+1BWEpt7TfmHCiXL1DbvAu3exc/RtEmHACcd6bsaq6+kd0NucU72JU51
gCZA1H6ZG6lCHEfqoko9J9OcEGdCgOCAWU9ZYRF6y5NmLpfGUn4xE2sf+LjZ0ZB0
o7OEpdOP14Qnn4M8Lt9oW9kdHtXRjidWF8HEdjBNpAZ7Ltg0OcqWZNHzfcuIl+xc
nFZmKjJFAa0YG7M/viX9DugAjO8c4OW98QevgjYjS7pO/ncbZhICw7p3WTUTAOdw
WxCyUdIgcBuaHwvzYQRSJwfLhwKO69IwxLNjTYSkGlZm2x4oOfgbYIaJeWoEzZG8
ZivryGA1VXg4qFU2a4F2WZpsvePGNNIUawmlCezM89VN8W6XIVmc5lZE1KSDTQfR
OGhHUSU4Lsj/wq/KFxdUnJBYNa+BKG3sA1bWLBmLTirSKQh/ft2dinrE2+7tU0jA
KyGpM5JWDNccD6L05/HR8i13nJq/Jdagr6Md+/EW3GmZJGNLab7+5F9xvRd6A3F/
4kqhMWykUuPIW8t/2OoFlOSEvbQChxy0dUnacBWISgSSsl0kuaFilW5jfHS1o8Ua
u0ASgpAXqVXmm/M/Z7UL+3yCQS6dubt6EXSFemRsLpWoe9afvKVjatIGA88vMfZf
4UEFZpDu3T4anV2xAEyqahcLJ5MrjX6qBHnYbtdMmZblLAZuyOrZ0XPPiInntWlN
5Kh4vXKESpKTSm+7S8p72WG7M89Zd3SxL5iojT8FvhweVPAK3xyLxEA8QP9XlBAg
eQfUuK0qVw07EP+6xBjX/2cUr0dr+OiK++ShniCoDf+PuNzq7mRI17t7Sada4Wid
Zj85PT2U51MHYnoqRFPDHUfttM1vzP0OWQHqajYvD7Zw8QU7ZlvQPCtBEkMW9+um
J5B4hgz8E5HabC3G/0uDYXisSx0BU3Ap7qmuFvYF7XRuUDZt79X5RukDFiVPCAya
EYsSM82l6ovwadhX1ajyKdlZy14dg6xWmOmambCxyoI+hGw1AKN6CoJL43F8atBk
KNa4ESPz6bwEQCxin4rtGQkhO2agpnSDSeym1NMTAA9nXhvbrbQhjPDsg8tk9RUm
FnTGF9/yCZEOAtsuSKtIjmoVrs3C8gBzGBDYjUNRpzQXU0n9LtPGQ6culk8M+qBw
oMBl+e4/RblQ28ejVIktsagXKSJBk8cAn0x6g3QXnG+815mjnKtkrrej9kvSY7Ei
MyU2LOk7NuWPuNOq49p55+557XAR8BYAXWWTKeHFTE9FYo5EDQ0NBjGd7HlM8hHz
5J/KdXSgWI6mqb5FRmZFK2y0LbKOoSL2b+sid8OzKOCr37mwhpoUGbR7bQNTabk6
IJW3t5sW5jeeGSoCnf+8EGnbU4VKFC1mhYeRpE6M14F2aY5rBxH4NRejWQyN/Myg
yWO++0xv1unZMwrms0f0rFmhc9C4Ry194beA0Z3ipsfkssY/O5S4NOlHBQ24rGEV
rhycSmuXiAm5F2K8scnUM0bzMaVCaULxp7X++rKxZMTxZgq5uocOtGVKGETPdTQD
xhDjeW2x/qi6Cy+HcKhsbaVK5vYxswtyv8ZeLJkRjqLRNO9edplcodZ011/BB5Tg
EbO9JrfGYcW1nTMq1CMnUd1I8SLmyEAovgx419QbsptKA3H5NpOoHc+ffyX+G/sN
nCrcTf7vqnoCZKsQmlpQGUWZnrDsZ7BFaJBs4bK/HC0UkO++/wQRDMIoD5Xj/xya
caNPfYet7rtylGCR3ew/1GhT5/kzpyJVM7mibNzF+HD96ZfGNyW63SpFIssOklQ3
xap9PPOZGpfk/nlUCpVzcavJM0yCn8as79VHwc15EHwWyVEj15bXCtHp1pfh5JDn
7nJGptp1/otNCvbtxDRDHkZNFhwH7fjD9uy4c4KONbX8nrl25WfsQ3f6q7Zuc9qt
oBbf6aHhovvtm5XU+9OIdkurczTAzX+cyUqWbxpIOJ5+Txfq3HwbEfK6QmsUKUk7
jhlj6HHSO/dLNewe509DOJ3nrV14vW5gTQs+72XoHU3WPePkJ7VoKtZ5rlpuYQrH
ytiI6eO206KKPhMV95HOHV7SuOVYeiRtCI9UAnUpUByB5V8sopRt3OZx6Y6K8FcI
Bvxk8z1CoQKOHksevGb2ct2THBiRXa13KpA2s/0z3DjAAX8PiSJb7jvCcrCPtY/3
lXZhhTYl+LrC5QeCa7NMAfMktCiJrdyLvXw/tkppCQBkj9JLAlL1Mf55903y5630
/Il8ukb8gV1j3MR/w6ckM9WqY1olFKFjgGg6JNGS/kO8GKaQyDfH2b+TBHtLpTRY
+P4ShM9gFkU8vhw5xaFKGDuR350rLM+hJ0HtaAb4Eg5ZJu9ICMy0ga1I6mdL4zSV
xR2Iq/obhhHS7rGxN7KxpU8X6VAnwlpikuFMoL5O4zVVHfrwx+FnzyS0Nm2jKH2P
KNFT1LyLoVmjjOpoHj9f/ALFDpMCAG1duPuONCZ/ESOenqN7iFb9uA9JB80tRqP1
+JH4puIlQzlj3YfszYO4firwuhCHu1mT3N5XW3PS1KToqBxbUzxjs3qNmWdp9nDJ
Bl9V7cGlIxI/oCcdYZ1XYpcH4ETJqoQrDUZXBzLjWMcMfCEhiOCRcJTVcJXAEO+J
NztT2W5M1I8FvnWzATFKfuRkq8keb5kYMgdohw6HxlJK60m58GwS1Vuu3ca2QQNG
6QH00zfZBhLJmFcvYoBI9rREVSDSVC2APK9NmD0Snrl5IDJ25W0YjZjWbhhxiigJ
9tfF1uFZpXBDQbT3j3JFIlv1tYuiYAkGfdabxPFKyzyd6xPNLL6gQ8ZVyIkkQXLa
hDRzfFU0yUcdqcYhYN+BiViRz8nn/SLyVxM0Nf/u63TluQPnvZd0BPJ8W9Fgnc9C
ugSbwC2W6z8nmwPBsu219DridF+C5PGPDnWR0EGpocpK0l15iJtET/MAL7v8mS9P
S4MGSyMiqi6AHNuRXxYoqD1D2FvohwQErbzSwavN+fmlGmwcZv8Kk9opnBkT85fl
Kp8dycRtTHyfJeU6dstqg243EkJsqtBuY+HFCxDIO6+fXq0Y7M9yrn1ha7gEnxgS
pOSLg9+wH67tQptT83vx28d3n98Pp5xjn3TN7G9ratbGNsbwiEnBIpgcTfVayEwr
NyC/TkqTciON64RY47RAdY2WipO+Iko/0MRUhaUi6OTloZhDHsAJc9/XBJ3j5cJm
URsKBEK5VM9FrwBDOzQlMljLOYLq4x2wrGZKKCp7AlpJs/FZsCGGjvk/XmkwrVDW
0DspCmyOBBKgu1Nr309Pitt+Bsl+7ZdQziuAduYBxdSMf0t8jhF+Stu6+ZBS6KTg
pz1ewqjx1LCJRl8iZTu3JzaY8e1InpzQrB98j/0AluuC8NIJRis8stAh+ayHPVl6
aLqpuXx1jA7ynUgyySglNUf4SYlY6LmBJBcMV/sdh/HZB22v9ub0qiS0WQGXm8sC
6zoVSLvwgpuS22unHIV8JMBNWum9x1ysc1/4Nks/0V0R9koPh9VlQEjdspPga5aJ
o1szP4RJjSf1HvHoJovN0JOWgxEuu3bw1Icg2g7UaVikhzmSMioy37w45iG8BLEn
dn15/vgUEPPZFBjqn9DsmdRyr50pLfKt7FOWtXhtW5pp/NseiXFPbhPyE2SjcNzF
lfq+ip1jwG1o0IFov6JhbjRj29Hlf2NboKEW7n+svSevDiNidd4nJNPeWwLYHlGU
B4WkytJgkOfFfrfYnez7K5OS9gCf/C/hreE60hf+DJOFlyzvW6z+tYex9VQrIQ1e
gFe4AKTsHT0wFSka1RLVmS8XQReYCxMWWgpVB6vB3VvbEXzIPaVI0jG8yJFKfQN5
0i3CLThVGV3XTgNUHWP8f8uRkyftvRmVPjM47nBiE89pZ4bKm8oDnqJuZQ64ztD5
VJFslk4MNaETk2Qqlmyy4z3AFFWT9xS+4xDdOY0Sip3/VEULg6bXEMWA79d0xFHD
nSMg9PPOzhYtX8HAntAepD6YNqaop5X+fEukROpVDH++7gbbsa2ElRSALzUufJAj
UJOOkB9cnZ6rl38bCfU8KkpbLI50P88oceaOr033I2A/FWXE78F7U++gyGR8AGoI
SvG5eCz0tD5p3U39JHGtW8OCJqPVoMWEi0K1je7G18vJY2Ya112VjykAfJ8IqThr
34SAlU9ZwlfWySVdLwHl51PQDI5TsWVHwb39fftSRZEWLx2vu1gDI6zm6pYP954K
qvp+oMBivQuhsZk3cmOUvVAW4WUncT8XLhaaRWxkR43SpBOcdTwWSsss913ACtAu
1ne0w8Hp6iW6NcD1gqV62gSTNhIl1+vvceClBjMbOdvshUwT8rBtqakBjeEgKEcA
NTKbaN0fejqlcmgHAnBXqLsMY5MHuLxP3oO0FBQ12a7YivpJ3zTTIUg0Qn4GGlwK
RtN4oxgwjORbiAje5wIdpVjGt59qVdeAlee3D+I3MlJtEImJutIYszG44ka25ln5
Gf9VbTdzs2XLmeS+EdojirHik0x1EeAA4Iop+YAN63huRj4LdbyPulZHMBR9qTas
bjp7fyZTFxA/tSupWSPA5ls2bxxbcKwAE6g1QW6HN72fcU71M9i4eO63fuUyP6jr
udtmOsVP6UR4dFlOgH+u17unSwpUBNkxaAqyao8jOMIaifnnsJZOmFhCEBuZc/Fk
kCtC+QTDLSfTDHFuxQBMcvFQ9GlKFSKGbrqaUreKVPcviBguCCdFYb8Pb4VL2zZ0
WcQf9wSNUT7iOoWq8yW/awStcLm9LKJ30Vy0+M4PwK1LQZkzMqomjHTJcJR9Uxmx
PT5mIOCDfHtbB9tkDkkuqQ5Yf5fSr/tGbfAodBWc5yJc4ndNSPq2XVmVFt9WdEGZ
A+hxHqKQMkBht5DaIkWTgi0TFzH6xWWlphlI371IvcC7d9WN3SqMaTlPgd9kpsdG
jyvKdJ7GoHhOoU5jfDHGogNO9VxHQo7JeVRY+FBohmfA/5efhjvpaqYAqRr8xJBA
KZfkqYf6okeLKerTic/nWHjkiCdUuDkvSxFJ0YPkylyW0v3cfB7bf5q1tKiGXTx2
CvdVrFogC61/0sxopNyBFsJ6NL7tiUR4e6liVRxD6P9CBhVUUCFT2mOD2IPk6Ir1
r3rBoXArwETgLfN9QqaWUUfeBL48LgPo9fDDE/d42xC6uNtG6fhBD78SRhoZPCox
wMcb0z98WjhObzia5jF6PQ/WdTPWFMJ9Bi276cfGWYlS4TyoGmwHKJlNlAPA+LEE
WxcHUjpQmMAE1+JZR2GtvIWMzp8wDTS1Hz+LhFWIBViDU7ATiFNBEiTCFFemPi2j
VTPKqt5e/nU6xuH/eHISfiubJ/Dedg367cE6Cha/ZyP1aNVnEf3SoZ9OhxYs+az8
yH7ZS8lSuYoDT0GAABv4jL6MTi3YX7ELxQ88D5X3LLw3yvrcaDsSQJHYlY/807mv
FTY48pchhiHjIINUooo+c0oGRIWf7H9f1mbmT1eP6Yj50Vi8ZJGph7pu+GdBA8ec
qam4Va0WrgxxjEmfSVtX16Z1JbgwWZxVaajRylHXGPSl6Rwjty46Q/hQ/yO7Ggib
hBYIxTecvZ1W8SE94ap0L25d4WwQsczGg9Uqq7v2RFIW2mpyVZvGEm2F0M+QZEBR
PMqqMT06/R54HOWErQCPScIhAcN9VxFuLrcQgD0mPGc06hU65ck9SNgHIQKTbt1x
hOsePRPAFVrEhuE5L55niJH3HHamWGxAz1Ql8X+QQZGSThU7EUF2LAeO/qPheQ+B
x/DxasrJe1kC2oRAyPTLbt/r3Ts3PWYhmwqo7IZ4xRuIoKLOj2cR4tHlwBYvztia
nHcb0F+RXzj/0QFggmNLtXDE73srt3joIPmK5IGH7Y5YaEZc/ILuzp7RCvbCUdMS
gMk/YDcZuwK5k5k7lexxWgGnePfDvPAT9AORgQy75uJACETaXNhLHWgPwJRvG0LA
WHiRE02h/X4UonzhC3fED3PWHSKjAn5OB4owWBqpPt1dpJkpLlROV9XRi4+XxfXg
k0T2s41NsO3mWm8kl7KdZKQh3k32D3bN+96X61DmIdjYPlV53YUhRf+5d/sv31E+
Mes8rwrby0N/rRG5I9j/EgANcHe1l/rNKqQvHXMfmtb0XGm8T8MGyHjoTx/lscDP
GNFp+xzCDxew3OfA7gfMrIRfvv2PCWsyc9ZJCRIUVesFRdhh/AvbkiZ6OpD2dgQ5
UjCPuNwILSeOu5jbiPGWTwmQx6yPrfd3GYjibfjuAKPDF1tAvQLfeb0iL8egDeru
75ClbnWnbf3HRfVdcHTiT2s/wVS7pRUaryH1Hg3OXFkh5AqaBpVMqrsrbdwkGBJy
ghywrSEs1fcMyPrw5tEVckGWauPt0kYNGdUnfzS+YdlaJL5aJpC3HSqSQQhdXFLB
T+1NStJ4I0D8sG8TqWHbozdD7kiD7MD87X0YyF7BleXFDMKzoHu7ej6dVJuNWKkg
XWyqq1OQUrao3Atoskiw5xnapski/yVlM6R806tN9/setbYQtNZrbTf0Eu5oa+6H
qcg9JqIhQ0MTeOQ6pmy5rCAncgMwDmYaDYPC1PA33C+jMqV7lFc88urbiqnqivDc
LBHq2KUDdZJe5p2+jb3jedDPNyGUBenDCJmndNJ41VqjlZl7t2XtEETWSZR7Bqwj
rPk/9DSAJYGAIkT3WBYRp9EaKAJ5CFMXbpLBSlPUSAkHKxA0KLxM1da5X8cCpabr
fwcSmlN6jCuGSu8+ObWO3gpvmWesSQ39xXLa+Z/JUIHbkHBkquqCddLqCMTuhx10
4lNQeYO/j4VV4hIJTk5IlXaPzKBYMaTIhfqz6XzgxLId/AnCT7iOoB/EwGvZTTAX
BK+o2Qu83pIMOlbgg1n0HJakPjqXtrqC39Q6KYXl3Gj08aVx7bsiJr8k9YGctwiW
VL9UDwNFRlSJ5+yfn9MCdUDAnw/BiSa/lv8UJxbe8HTy4OJKGnzDPqdZ1Iev3Kox
X+z42r+9rrJJooObTvhvDLX5u4PekxnQjaGkcbJVHUx5g4KbEXwLXYrThM1KvWT0
rTinRc8Ant0feLP4Lr4MXZA5XnZ+9yO1XFwDA5UK06auqHAhCHUiCAeqZ0tQrHhw
Xmr7DuNJ1+2yb/nnU08VyPtPc6cZTzbiwtn7GDDgrjwXWbxrwvVkdcJk6hxn7He4
05TV9Iufj1zyApHSv864LVPRJ4HFnw4Ns2T49I9spb1U7+8sqInSczIdVeQYDJgr
SdOPti5oB/wbSyeSVn8/skP3kJ/qAtzsSETTNLTacZt86S6VQ4R3Bl8mXMOsrgXX
jAcke0bM8/aFOG8a8xjK5/wr9qLJG7/iOnH43rPoGVFHsIJayRGYYfPfbQbfi0DZ
oqDoHDN+34uhPoI/joOBShm+DlxtI4soaedgBUEXi7LYzBb+hqTcb2H38gq2dWSO
wIWuLjss5ZVRBpg8Ui6AcmryN6YHB+he3ZdcvSs+zrcGZEnLhOPfk38RDxkS8MFV
EZ6XzOALKXEjhOc0dl7D1XCEbpFCvGzXanOs4LSlc330AU3nr49xHSVDLPMIRk79
MIE5mgVgbn7DMdYANwGH6XfEV8H5qde7+FHtUuYfv85edXKwdjh6IYL3IzFBlBwe
fBpf6xM6mZP5zM6A+H3BySFZDmmxiLC1dyIGtMNouAeQIHlKyigseViqNxdnX0ft
bC227movv0bGGTNp3/vYtsbF57/I9TF9z6g2KPhIiWAeb5W5U3fYou3AQY34HKU2
QW/mtdfH+G0f0l9nDqgzHpFHlr3sVPV3tF0fA6TjrYBk3MXYaoGm8x/oTRufoAg5
af4gvZ5M1z0unNDvnpLU77YTNInHScj7nr2el6NPqBL2MxH40OkZbzVdGGfk/XXa
IwDL1Y7lY2QqEhu/NI/KaCKjkcY7ClQuoukLWKPv+co4z2YQVEvu2IPaFzKBSnbd
msFsdXRHssM3KORC7laGmMheKVZOHB2rDUr47FZKxk7gO2QBPOyl4miyNouVwH4/
oftm5gkU3/znPnApY30rGIjyTJ4jFyLl6/WnBfem17xMuAR9i/6KjnoIPn4oECt2
p5a3ITm0LCISwOAmFXwe/GvisxkHzELLORxvY7hTanUID7HUqQXAM7aGZUAHrHGS
Cwbzesw+4oZt9gm8vJ74hhzRBrX+SAEF231HJ7Th8MiHjI6XE1Fjd8i7JXEbGHgV
DjSB4aKYo1bqWgvmNDh57q94NBkUReyQE6CcefNOQrm+Gd0RUZ5zENoDJxPS3ggw
kzrnSrQ5YmysPhX+8GQPOyTUmuVs6XGWj4gBYSHazxAeSX2zALpQKHUcUIMb7OuD
9T52nUQXOfGcHl56+kOT44eS2569msRsDp24eMqSi9QdrBe3I/h/RKHZ+INAhkGF
PYGEbl21dBk70LkDEpAIl+c0b7twDjtbdeHmvDUMUJTSjAamnQkPaRVTEzjqzPIn
ZAWWNTYn95QXIog2RKTGHHH3BSWNZYseEm4d2wHFwNGcxca6Wqdl7XtYYjrZhnQI
IwJLhWvPGi6hBHySZNsRESRF5F99I88cMvSwMvtJu/zRQwpO2weS9wnQNoN4ZGRh
ulePsFAGcjBBAXCgH5YtZEMR7825lGk4PMcQnn93GVHKYQEMNNHZCKxuG70Y/710
gDYfj0KZr2JroM5VbSZBKfxdKprDnXQC82MU8j9FE1hheQ9UGgw1ileqNI6cZbK9
nqHX28xilnKRatejB2UOlcVKqBHeajfFzoHFSHOSUYkQ0QZhE0bPyk0595d/aSKi
0AZD3oeP96B3QoZNHvMXA7aOrGdZRCvfS9HQgdENk6XEst7eVYoMDfJKXlyApJuR
yvAg1G8eY3WyBiNvGYs6NWuF8ryGVjqsHZkDC2ixRB1IPRBI/mYt4qy2REweHUKy
bFh1UVPzbjK4ZCrIqtXtOp6pO61iaorTiDkBHTQyxtWtE3dxUFpmpT14/R09iIl7
YXKPYIoif9EwmevhDAeQaX3fGe/NHIDJRg88g1VrkesANa2Zr/njc+ySKvMfE3fP
wiCvEsrhnRPFvkAKKkZEwOJyQovO6SJ0QmxJjfaJ/5bdzxcNjeKezQSuJaWmO66c
+KHlGcfU+w4jIKqu/dF2uAgjBJ56UjIoTkhOx01Fza6NzSQm6z53p0d0I2V9fofQ
BX2bodNauKK1IHtbhekvOx1saw/W+Oq40lLsFqsdNUvWe26TQRg9n+t/A0zgDJTT
z0XrPkDpTMcFnQeOs+/IN/0RWS3pe4X0dJmv0B/Pzb0MzUKtWdL5t8JLPQUJ2PMY
gKfOK8DueH22ds24Mbj3dVUBxUYLWYWwYoNhfbOun9CAs1oEMPTE/YmfOhY9oub1
z0GDAloqf86R2d9nKBrNDurh3AOyM5zjJ/xuL9hQN5Sars3ahUDECpQ2kcBgoNxh
VEfUdC0zLKZN196UhqfdipcuJzBmLkr7Shn7MosIs/h7PvY0Bls028B0WdXeI+aA
mz1aXR4P05Tb2s1IuTm5zG1vFZrA5LRYarKsJZpHZEmA3ip6p+I4wNqMtozQC7dZ
JjtKcDqOFubXsSt2OjdlGGmcIwmv+UA7VCa4S8RtnyBssHIlRY0vB8qadeFcID82
ZsKn+rsXTNa0xVeoknkD3uOzlvJZe+Ziw0+px1jheYe52KNzQz1AAo1cbWew/vB7
IT9UC50NbcERM22o0PdhY6Fzux4DPUQoSsjLqnYAyhEU9SxOwdPg36qZaf5aNEeH
QToSdqyzEsRke9c4THEqxrlRJOxmnOur3BXdpTprzRhxWzka4Bq/OfjTnAqNM2bZ
DmGDKmEDnZMvf+zakjDSXfM/0KkUezG366zDBK3+sd+QeIR4QqUUtJLSaCAbYyYW
Upx5DTSZSknpBCwECHDttBtUTuF6qZWBldfAD1FZSRyB+E7PPheaVtJZKL/rc1pp
L2WdnTCIeh768gsUmo6mTt1walos/waP0dl9KKkUIWmkqcTdKmEXlSGUNnw9Cmbg
iNvbJ6e3yXrX9cOyx7pbfJ1c5M2LY8+yUaqaeN3KU+CjdXtG0T0Kjg5vYjoFDadF
HFpDfdf8+Q22jX7l5hUI9jSVEYf73VRyX3hiUoHKEbXDYg39eSAwp0YAOiEU1fMW
hWc2/Q9pAjkqGS9m8eN0vsgGobHZC8Vj9NdrcvvMBnD4zuAx8/xmaDBcXwwlWf/7
08Xca32Hpd7kR5EohO5g6JC6HZDjlx/w9rpwPevrBeah1pFlABGFAWZ2iJGUAY0C
+nKZuv4D6agpsEvp19WLFf8jjGEMvXoqkP4mmvWz3Z+wBC4cnvvjCK5jt0wLTbXk
XSze9+1vLdLMzNtqGy+OOW3XNoSxYqS7meeKZz1eIVzCGiWAc+zdUj49rwxGOdbf
LC7i7XDD2Iz11murq+DTDd+gHEN5ZB7W6tYEL9RVCBWf/qgt96mKg1vawzn3FDLr
XsJBJdTcqvqBotra3iY8r5FeH9xo6PvQQvEcCEcyGEqPUQ22fGlR9FhzMU0ImwIg
OQVWlYhqhwKk/pde8nHxmAZbhmUL5vTRrFIsP/Qtw3c/QT4sUhLoI+qNxUTTn3Jw
QBJJYwLnqQp+ZMLTBaTyARUePrUDYFKeT+CxMRhfp1aHzVfN3/VtMeYZzceHiar7
aLncvlq2BR6D6taP7LQYihZij7hTielR9OEXR/wgbpqnObeNOrSWg+HIygeBv9P/
3eXaqJL8brpheZKneTv+XNypaWMMn8lfpgoYqgYnlmxsm+68hL49QljqUp+U/G+5
Q3dGBWaiMAGEHMyusHFXKZoIMe5/X33HGp07d9dAOPd8SR36X2GybwcijbLKvZMW
D8wOAu3pkzkQ/U9U1ZaGa+0VqNNAW/+AwVzYCjvhzEBYtNr3pdvhqvEMja/hxU0E
oGksrsbCamP5RoeJp3EtzcYwGcoKRTtmDceF2nr2H6cFkDM/uU+Bs8Sl+d7TE21h
/spkuQiukBd3uyv4pPpdPw3WbP0YFidKioEwtQjoLUU4797c3b+j9F7SuDVcH0Bo
bSHKfGWy1w5RPzFM8VrjJHcg24D2n5W2Sy2E7yRJ4/nSUTFi8JcrtGZrX+qKkoFK
puF1PWHhnZMPutvo1ajqlssgrkfFgKJZZB0bkBnYhDooFvmIXnlQZ70RdRbxS9HY
pcjLU6fuWIc2C+k6Fa3gtwxm7GTJ70Faq2DqVmC/jW08tkvX746ccWh5koMN9oIr
qlMGCiq77+qY9efvcLvi8pur2hbjg8jz8q6yTmLCzk0IWHfHCoHTEGxPu147Y87n
kxu9qNdcETyhxv7dThEKQYnjQ12QLV3ICDPOGLu7NeQxq7iy4rv24/ttrx2Oyh88
bnbju58jPrBI3xOYLarM1l1+utvUeif2+hWSxvrVtE8a14jVoEJKyBaH82N15TG9
5HguKgW+yaHuwfN1VHIa9ikKQKn+ZV/f7R80JHiyJ8NNDuRpujvLh5t3JUpA4GQp
YNkjeG1HLvW9YvRgt5dhmbwf9iEi3IcOVuhtU79l+r8+H+5z94J3Aj5VpfaeejEi
cszD1c69qShkI52i1W6CpLR3dNUakxUFGjo8RXa0SlXYOL2Nkpb6QBtuVlmXb6lF
uotep4MtaQsecAxDJGUlnPnE4fLK1/quJ7mYbDhNqGjsmwxGqaCk7AVqlirtFU47
2qhmcNBhZ0queMpEW4HMYXnYigbplrpbbWhsWxVYLx8LStGEDRUBTKdSjOMbAroT
Xn2r+BHsKZtWvlfXeRsvAVJ8JL+SITeaptDpd+y1Xpg3Ibjp0+bcIepLC8uEs0YM
WedRFG1ShAKbW0cq81BrVF1Q86BgoTzDHqKaYjAXhRM6JgwyqmZHIcDsv8fSnYWr
y+uTzx9vxxU1N9tcQd1FJuj1imgwn6Bk/jlkDtesewxhipp/VVQ6UZiXTAz/x6z4
yjGZOcpqL/rjqJCqUh5SFaI3XQK8S23h90gJ6XCklRvc0NcRVPIFPm4evwki6KVG
564P8BAob2lGIULVVPGnu31A+kk2DUtXFblcET7CFnqeTLKKQtJnlnWyDh+Dr0w3
g+Kr7fpuEpieHEwMzXvXI2zOnZPZJmNDEiu12jXANtNpGKU8Duy/uAGaQyAb1KSQ
nsm//oXFnN2kgA5V0f+h49rCNMbszqMKxXRBfRkNF3ex0HM2yYcOaIzvWG4n/eTI
+yv0dzIwXy3ozwCj903z2PC7b0bZfv4SOVx7dCPg9Vnh5gY9JtknYRggKKpxPFuo
IZfh/lYNQdSNBjcg6GH/gBr0zrbAL3ZuDkq2EUAyvu3abNykBzSNC56QBdo7qr0W
p0q/laR9NyPCRnl+othOh9BjFgq8d27wu0HOMz5BY6ZDI5SFysuLTdJxjSP9HWWL
hN04k0nhocdhpiNqg4A67O6efnQm2WY4bdlgCP+5zkhtJH1xXOz4sYhVzbEgSJ7e
gGI2EUJmrNayr6E606kgT3u+9UE37g52hwvoH0QtobMmBmkqq2liacItAiG2UpvP
iQmUMkBiF32ssy1GXNMqbEiOzHpCv77A06y3T06sKG8IARzsB/99S8puK5DnXYcB
O+eeLBP4Fb7ckeuhpZG0+wEvQUWb/4epqXS8Lq0hgoc/C/zauHJfiqp18M2qVjdz
rfQShNmdASnSo/WJPO8Zpu9RNYEDbKqnuDo2qkC3maMq+YVe6AdAVZoBKRZymOGd
tSjWmtkpDVShVgIx3rnsZJzgzz8XuRElFGzSWUO7Jiv62Mtb8b45flonpa3bHc9R
g6Y78A1bFVqS9AP2aCPEE7rB5Pq9LW4twlMYS1lz9ar9ODIZLkt0PiBwf5JGUfv2
ne8sLnfeM/IB14JY1Gd+lMVlVWfNPOMZ26s5zm/kEovfdMZjfcKO/x+HOT5/MIYK
7GH+T//LvGNTrcAXQw4VTSIlQ+u6djj9r3ENBrd6wPLnvJAsY+gkEep2M1fTOFVN
xrhA5wf94qtI2VSeox6t2OuO3i6gUg7PV1UWVhBfzoGVZqsIsFiQt5LllUpbDZZV
B8yNonkrQDAjubady3Nd4KSbOlGIiFY8VsNqKFNiqUx5HjZ9EcaOg64GSMBfQQYX
Y3v2g8xfbXvc+pIjnPiBuYXVDKI3VW5zewJtGI7Vc91N7Jv/4SyLlcp1jSIHRk6Q
b5RvK4GDvundr8EguqZFaXUo4DAExysL+zAzn6i46aSXiqZApY8OIBNwarzYCfSy
t1ujX3BvvIiZ1i8/j9cZjI/BTCIJlvuBMCI6bzur2fzx8uW9Rey9GDTa3fLRuauz
D/qv841kfNSlwnOtCOUPlkwINP3C6kxQ4T817ZXpkTwxr0Fs003KdmJytlbDRRBu
IEWTbn0ETT4AySioIRR7vVfLLqmVEdO88Egmui4jJUu4jjgGv4yBbQi5/qhj9Y8G
3Zfyfl/+w4K9NO/laC2Owh50KLyXH+MLVLs9To0ILZM1Rr1p+8V/zvGt8j3FOH3J
vzc7A+KZMhyNbhB0RVeBViENjBcWwOMDn0gvtEaPnZcNZ7HSGiPzprr0uU3PzlbT
1uJVLIzLoxmY+bN5w2kewoyy/PveseY2ePbx3Ge3BkO1OKTu9xBdSdv74h4y7e+o
5vfmNlVxtHrtqx930OIEtJR0iZCTQb6v1glgcarFpcMjD+ADpYqQMfq/nnMcw7NW
gPKaiq/yPCRhlHtvH++QoykX8shFIZNMbUK/0RXEdh0wz5n+RBzQwvVJkvsVlv9+
oLeFLI7+D306b9mTj5Ugnxkxk4wuHXrKekmgFBSrhy+eKhqxesA2nb5Y+ebGUAvn
Cffgn3xbg7dMZlufCiA+gLlb3c5JANJuAsIGLHG9Umrb5oYTmch9lv7eHLDceS++
tYTmwn8rkTbUk0kY0K+8zsfiA+pqhnL+J5knDL33AZRR/+W3HCWOkad1JATyuZ5B
5Q9uIjUNCPuNhDbxXAZskyuibaZg8ieEYC7sHF1/6/T6fdepJIP9WqBaaevWPkJH
9zPzqjkCDd7vOYWhUaMdUM/OLG0ptv/XX3rcUzQEPSrgA3UaRLeHhDvAN9owdGR8
G26bK/oIADgsDdn1pdlg5QJpvkMUv7xLStMDTgx6V04gC2Q6kwWt6VyMn7p3LGXg
RxRJRbaL49yknf165g8hcB+S9NkVc02w+5pkqLnK95wAGwW+jp0P6xWJqW71NZO8
XZlkLjyos8CzbBgHgXnvGoAoKHJSXN+99mN5TW64mOFt0cq4vE4OTZsOQoIs1DpZ
Z2scpiHaqqT+rF0Is6Uiuv7MRdFdwIBin+Y2+1CDfSMfgKrCl5lLsIrols9s5/+Q
1LEkPRkdDzIQVsr3eWybJHK7QX1gAPtn14WHvC5TgssIPHb5RpUov7NG547z8xoX
pxFkfigNaLnVShrMkto6JBDXthBBbjQYzQL9hFGuNjhbfi13GA9tfYAJhPsyfrEq
hVfziDqXS4wzP4+1Eo9pKvKdSmYoNRRZAuwUrYCGs5bv2UZGmfWXmBDExp79RRCs
qeFI6YgoCB+fh8sylvMNhb1PgKhkTHmRa3RDKeBfb45MT8FD8IXrduuukwoLlIw4
W5SO0BUdyDhlwtwS+IApAgN3REZUzfqfhIglstF3LWgTcnmxIK2Lqpy+VFUeb4+k
xKfTbbv8EaOosZSVaPXByVM7vP1gPTx9JEbMhecrFunCIO3Li9n7q4SycwW4SAha
Ss1mS4z31stEC5GTRDtEbNgvx+wfmm1x7w3kLHPllkW1QRq0l0JnznnHjyiv7kVb
RO987Hfn70JMo3Nwj0rclCEEyGL8EhJd/49/wSAomEI4uuIXVndWu9CMul4pjSNz
ncJdkwtOZnYkmWZGnuRolAIQXcTNVCyK6XYy9SIcm4IfdLjtaU8wk0kcfOG0Ofbh
P3/UtTTZX7ENKAFQy0LsrWVnvSvFYB8A2tEwSvITc2WTjnNdwh0M0En0MUTe8nqS
WL6JCGM/TdwekikOETRvYJ5M5wk44dEJ1o1aPfetBerIS1kdKryTXpl6PPfOH/Ts
H+VcpCPHGpKcZld3B5XwynGAbUZrmYaRchYpcEgES+t6BcG6rQ9qAh3ItQA3Il1G
yJPZ97fJL9X+93kx/2z5etXF/6Dw8RW+K4n3nOze9GDEsXohYi8gZbUqGAfgDgzp
wWf7PciDHGNa/U8D/5kf2G1Ld2YOqNHqL5z9cL8AtnFbZu5yxnylqlb6AdoTBMBO
aInelzvveVuxItbtmlxbzZRo1E/xLpi58oZ8svxgjD4dWbOlscyUZg5cphirGuSi
W4OuLx0AzOMzB9qBOn733zOdSeFTFt2uhNn68v41yUYFCEJmw8XOuqkVEL9HQWRO
WwwXcy73KtTb2frywRXo6q9euQoR09yIcVuexmGUi+C/MZ5/MOj17sLEdu+g3GKl
N3AF16j7Cn6knwdpBJHrRFZO/Y5m/pdRNn6epOFTG12hXEr1vqCbeYin1xYIrwuP
eF9COniGxrnnTwPnQ7lPXSpVxBvw+jeen2Tj4GmYrWxgvvUVnuqU8O5yMj1okTMT
E19+icUhgRMfm0Jc54f1Mv3Q/9/mY3T/upa1Lib8wtPOHOP7he2ZyA833dNwl48R
L5ZT+Sr/TcrKxEx8IllkYY4ViYGaG7L7oTJT1u1rp/Yp3HNIq7sai040alA2ORWj
0l3xBE4DApvY9X9al6Ra5crDiErGezA95tBVnwScWNQr/uJsacPXvrttYW/5lm08
z1re7UIPWQaXKyNF4arGi/f3bkr7FncVOnHump/OM6Y1oZ/LiPKuDVN0xzRDkMUR
yfk6poiYm+c5opY3W6RwHAaiwuMvMGQRgRu1aV78w4evnOTkg/6IlqKQrGbrKbIj
lAj5caRbcsVHvrBlI14QKQ5sWRxJ6wS5lsFo5qIkMBQY+F3UCkjN0J8WyPXnC4ES
o+pzHzbtugNtoWG+ERsJXXuxD1oFmrFYRIWWXYgsuWc/pssnEKXegJYpBkc0ApaN
Jve7am+Ko0vkO3pkDvmOt+od5XjlGXxvNQlkXQFlcLqYyiAWZIBt1yR0mlHh2YrD
qigB4I3aVtSGUvy+fNA8B+fUo6OnsjTRjChA2snkkRa/BhAZm8SUQHeUbRcyCBGC
hrBTv48U0r5nnqHvqHGl7ut29V/arBLlcZQyvv6NgYP2TBYwi2zwPGv+/7VGAMfa
e59CHjUascWfwbYmY2PhsYDiHJ9mn+Lb/o4GDTtBVWO+ytUDeBcNv06n2OWVpgvP
lwW5E/4bOzzNk6jaPmsUOy8hV3H2j2a44xNue4IAggq8MtI1v1m5jXnoEoPIYSs6
mf8bx/NhNzR61qS0XF/iTPzhPzxw9w9a2zFaqdpypj2LQiYktA0DSvMDdpNIu381
CYgH/ISaHwFsH45afVj0cXlMIR5xVMKlPNxUaPzghfpWAbzTNWxYhwvEwbzj/91d
jJkVc7qEWv4Q3V4y814Uahk11RMm3vg2i9K4asC9Wgq57ELquXHoxWn5R8xlwNAE
76ZJZ/VZB7N2UTaE1hpPdNVsY66HHCR/RMD8/OaeJel5u/4p1uy73ox9YWyJzFX1
NTQl/OBlnMD/t5D0cabJPDJnqN9bC0gLMwkB2SST4wq+C9B/oSK1BFeEsWIjclEH
O8J2NbEtVvjEKZXq8SKD+LR92948SH6yM00zq+nnfG9qqN2vOAOJsRctfDI75lk8
Qq5n15i/Uq5aAgvtctVZb03LNN9Sz2wE+BkRFI5aly17lutLNDLBNmh4Jfq8gbCs
B8BPg68w4jaX47SCy5Oxtwzn0+fwxQK1iSafCdhhiFnejqxVwCyRFj/BE66YqPI2
qasRF2qMXU1YI48lZ1C7BKN/MilYvSsZ6/Fj2Fxba4I/qNcfPj5lOd5wty/tQpHF
hbdZKHQ8m67GvXu+0QwcaYuzbiJX8ojFK511U2JjnTLtdMadcRffFSoLYIq40F/I
EJPwIwM0EKyZL4qPagc2Sf+ajavlZAvLSCmQpLsC5+nZOge8/ib00z2I8O2QIOWH
EXReBxqxgpUWkMTdv0wcGFZ9bDgr1pu9ykXLaXns1t2XhFE956dqm8lov5JqPDKA
kVBJ8aKZvlFnWzdflt1uNhZqJ8rr5R9TEIuVdeB14LC0cF5MiqB7VbHw/bEmUvOX
sEJ1kLwApHebhbhy7rdkoriEpRIHOCJ/lUbWrufBGuENiYPx8nkBNUoA+z8wOe0b
GN/AUcXtexfVOd91ZJJBc3OEu7t5oMou53JX0+4pJhJDfHI4BA4BBwi9PxDySaw3
+WO+Bn8YuAHnoeoAbW42fsyGSaEaZQvqSphntdXhPHbMFCeRhRiXvhfrJ8DQnsB8
TsW/JVWgk26xx0TbbH9cbYbLO46+qiU1KXGoe6jjCu3GytIolgZbr1sX7+c70RXI
17abaHihqpu4zLUWPYMZjLzJgcCwaPK78OlY/BbRuB5lLOzButBJ1UfCIur6A4DH
n2R7j2bDpspqDK3ix45DfGWQZnMPyjYD9R1L20y2vuP09J+8ZaenYCDlqqxYxNb6
9FYYGNDNacgt5RHCOhBLAJdfZf4aQJlNhBakjYJGeLVBSKj/jJWq7R9l/+tbHroW
YO+qubZCIhH47ZEbSatRZyEGojFFcxTPdTXC37h5cPqUxBUHl1BGivq7egJakMrl
lE9qO5XS6vacUEeBfqud3FOqQkrZ4EzOazNrJEwO/5i69KYVXys9xY+g/TQTWTgp
axwDg7Z4oj0i9dLOgRUjRtmj7HnQ+ozp5LqqtSlUFCGVBkJXGGNvj+NZVip25nol
wBE3TZCJZXrCrzm2Xb/M75Je8wCx00RJs1dRAeLepHREVPWv84M0M8YQKrOfDX4D
Oz6bF/zITtmCj7oYwg/Tl4jtrs/sZkoY8svyZxxvoRyNJ13HDPwdUI4uAfxOOv4Y
9P1TLYMWoDm+f5rnN8rzBr7OMll0wr4wJXiJVc/qEa9iXqwFGsLr9wM4+uBcW0sx
d4tOq3XlhvYoPfGzjZbs0cgBtfI23sU/Z2Th/jWjnoa3vcw6XCsrQPWYmNww5ME5
vb9tAw0iJ6hAGzN9EjVmZr7CLfFUCNaV2X50V5p80Q82zJMppR9w6f/r7KSdSK7I
hdfyFqn46UrDw9MTHT3plv/PWjZb2KY0jSTVtqTCcTd7XmkoEau4a7jYWYb5QPaA
+4RPE4j8cpGZ81aZ58hTzpjf3sf5mXUArXMWiayAMD+B8xAlpbmITDOQesagzmbT
D3Yz47wRxRhjW/0rVM1+qX03HjDPOEuIx4lVS473h2lAbGnw7PRAElrm0nbMa1QU
isbXBmXwWF3I259F8umR3IYaBcej3JQjlx7J2fBV90263jSQOQbzVHWyicIW636i
UqE3jQerESU6sAZYbSy8TgAX5UjGjZC2e99iMrFYhlNcoUiMWXzcQa7ky0HFDyZN
zxVkWcWJuQzVyXYK/TF1Nw5wHqF5/548spdDF9h4IJgGILrB0TpEI2+xBIg1e3UI
1uR0q3DtPBij40Xh9/PCsFA6x1ZzARrp6JIi81N+dPUi26vQLXMwRwdnM95cF4K3
LfxEfQcYc2NfviU4fJJBsF+28ofLLb4DfKvJiuuBUYcnp7ny+fjW68Vzppkd4M3B
iNyYemrGCrkLRhyMV/nEeUDZtBjyYotQT9G/fXF3e3p9tf6HoyFK1wddJAJIQjSe
KVEdMfQvPlCQpndpTeGWa1cxUEz+L/NmcVeWqqXgeTE+frrE4+9saxVpM6jrMe9o
cpvSu9k9+jkrlX+Aik7HXkqHwmh1xDV7HfdgNkBlfDFzUvUn2O6zZaNjHK6i5MzO
WNk9pO38LTi7lNdzUGKb8WThF5x1fkpGWqmJde/hwPRKYLxeVDOslkZCxKt/0SKu
pnOCkYTVhyzbkRWY49FF0EKGUrrKiWLhrvxjGiBvM+Z6SnAgMfqO6K4SV91S+In2
w/5MQRnr2hd2EHFyxBzs3vX4R0ALHaiIDqRf06217Ftkt2jq4GSfWfM5Ne9RwS4Q
f70xT1y+LpyNUx/Pk41+X/SdWKQKliqf6qcRNMh3sSKmG/Hmvk/l84+JZgR1Ozr5
6cX6t7NrjA/fccXb+KPUf9rQjpvh53oG866jJJEqeVLQ08kMpeHsQnLLo2dr8WOx
j2hE9feqV5ujVwb4sPXREIT9LsY7FMHIrFXSHgR7O5Kvf/Zck9x+/8s2wmi0cqHJ
LFDEoVFCSvXqQ4WF54cdgNpJAFSQ5nQiEmtrwzCq4W87twCQ35B/sDkKAXEjZy78
oEtO1WAHp1wjtrO6xcY/d9AyN8ZAmcaXyb7VNXBFGbnG0qzzvZblvGul4HYlGLok
RiezJufsO7jvRlpboYdFN7A0kVovPW24pRlzNwxY0/4GzIJVg8ATJZy4L2iGW9LW
V+WSpDYgMrFZFtE5FNwg0IhxBXkPh1V2p5HKM7rsr3n43jMy5pStUnRrh5WklEDc
UrX+E/GLIaRv/JeWUVB/E4kem/gGybcw2n2p3VzPNavVE/3+yytLUk9JX7n6H/4v
EQvIAxv/0PA1JCHEXIuP5TUeBtpyF5vkn8QpVVws/NbqKGQQLJnHV1KIJ5Th785u
sYfj3wN5wYZieIBU/Dm+HDmNDE++s2WPwwEt1/yltBmUxnrEb+25bj5Eq7wTl1vz
LyQqixqDSv8Hr5b30ZBwz/7sHSTjc5eMg7MGWjfYBg714sx6DQ83HlqMo/7gwmrX
k25CGbQHWm5ISwiasPZFi2ZbaUhonHJD8S+6rmkKOXH0/zP7vJcUpw9b6JGIseO6
tGRhhZABiWCw3fOx7+3R+r0TRD7i6FjyanoZMdElI8g5GKmUvpqdSk7qFsBC2nGq
S/cHWGAbLvWur7aSegNPNWjGhucKieTTuXlKR9njPsj6A7ls0EKnOl1ZDja0jmVw
mxQeaFXPInBKchimqb6rrrhaXGTx4BBS60hJ3t2HlUtqSZAhzHCa/3BLNLmdz4Rt
cwkOxrNl1Myy664L2m5mJ0Jt1xGvr21OWoZVulSpIN0HRRJlNysCwWTv4xlNGNHd
oEidB+vuR/2ZDsDn+AIk11k5awcSShNWGIuI2BQut6xE4pwv/pKbdKKkpUC6BKFA
K/SB+QCZnmc8f59d/064dUfMY1UqMvJagCNbEgD3q4SLEIv4RUDzP5ptb+h0NKNL
pChW84BRZCgoMYF9gs107vTPftvi0LGv/O1TrX+271ww2oAOW61TxNwE3XcHUOm1
RJGH0WUI8xXmB4Uj6+ZWIw17gPmrXeWh1NPCvATYwDW6isxFWdyv9jLYXVnP8ndU
YuaiwPELl+oeSzh8qNRps0mqq0vizW3D5PKpZxYk6BdDwYXMOtoz6qRA/8ku+C9V
lKDmr8GReQNt0G2azcQZM/SM1FZc2Q9Lb1/Ng+xmS+6geOpS7L2mC9W25aD79iGb
YtwFCaTXyt7GKNmhadsyIDPTFrJBS+t9C7ntTW2XpreXX9Q7vW7n0DepnxMBbr7x
lG40VGAshC1nGYJ+89Q2pbQjd66S5DLCqPCht8PtlKR8BYBvHf25SD4a3EV49xYl
IcggcSeZoW2CF3BfAOTsuS6OsWQRJI+H1sw1j+2Sxp0khoxsZcq82FMWtr+v4cP/
rGpqjhx++hE1bzMUfYfgq/65tX2xAxnz0njaKht/avhZ3+AQJD6cMUN4puOnjGx4
N11yJwyoTcCHQE60bDH+/xcRrt7lT+T3riTDmVf8ZIrtz4KL05HxJMXOAoZc/05w
5sxM5m4WjHEoIcNUsYrMSE9VI4rWC4XN8k0yJmFu0xQg74wEKchpIt4q55g7/Elo
1xL5Q7NGp5YA1kcY4e5lD56NEWavvwaE/YTx1qEVbAcr+a3Q4g/wby1R/xmEiWDa
OqMTFEUtUbPN/Hrh9N3CmPCWEvfFQjGBdHJfObbCbd2r62HQAilw0ZUUYIezCBSb
LPukkR0GDj201HdZ8t1Q3E9HeBVC/r/1ixjaw8264EOdB8ibRu5lhuZO+PyITzK+
+gWnMfK3+6Poyo3JJ+O6B/z6X943lhL7mT9TXtUWKRg7zqBpS3BcUoyt7ks7M3+H
GboveXWuty8iiLEfkGhDN2brymOqIAPKS4TzXUqqGKtA5k5BkhIjBa0/wNForlhV
W8gWO1U2BI6tcw2q/VqK0gjS9Sq7tRblXazd+T4mXHNj9WWX6tsv4AB6QJ/yvrfh
SDL59pauK8kR63OqUQkaMrI5a9GNzJA/rdwCwz1ot89XNyIbF924llPqh5JNSFzj
WvWJyx5lPCVVPqaWt0k9QridFmdLNYOdYrzjtlyfa1+F1FTBSlVlzQ8O1bI84r+S
PrPtiW21Om34CWo+2sicpwhR/sWdHzqXlaJ+wn3zawoITSsoeTfLBtnEBy9Ry78G
eiJqztB5LNxQbaJFIEe59MGpAb84zhMT3ZqELopCXJrtwfqkfJlPDQIHDkwvvFWu
WcpmhyNwWed+GA0KJTsbmU4x9aD45sseFaW3NfMXN/0x0iNzgvCT4Ldg9ExQo81n
Y7clviZ/Rg4xIEqP1qD/ura4eX8gKBz2fqVehfqGLMilbA2ZObPGNPCAArqYn4od
XDDLFab0kd4msM0P12aI92j+3tvb7kxP7vaZ0vGqcqGZHmxo+fI5LLRDDX7zztNP
ZdybzQVqz3gn7JpVlgLS92aaYZRH8v8M7IK+Y+sXTwhj8vRACIfFOVWpVzdBzcyX
rpR+4075qbNNQ13JWdYbGvvtk1p4mvZ2lTaazhHTsfqQEQ1f7U12cQiukVtd5FEL
eqLZifLKgMSA26I4VRsPYdfHra+auwXXRMkIW+IqBKQuW/ozGS0Y8DwDhRNbzfIz
6g1BTmuVoIvIUSjExF+V8YcJzofTYXO4IyOD+SRYaObuptiInvT7/93qfkl9NS1R
4y71+wSt3j8olcYZYNJIL+04nLMowtHQaqwqL+yZO9zhrYNBfvXH34vpJM/E6YSP
UlTwrV72lRp07ZJ+cnrTv4mJbreubQIHwM/tmE3+PC/jwfk6VS0DcKqpjIcrEoIw
8S96UT22K41p3Ae2jV0Tnnh3ZsOxrH7jALjYJL+RuS4y1ws8NpL7MdFTaMLg/50p
q0QVpuXFYaDln0tHwtjhynRkZLyN9cuzbyRo8QNw/6F1IvW2A6fkR7zAYdkbOI6M
vLaLuT4UR7QvVxdneP/4H+7tTDmyZNNdE3mxq9N/Fe2z2jxp6NN38X7gdK2Fqy6k
aecei3kBrT/cDOPSloto1vYC+D6RS0s+pO9EA7lvoAWyr0UlMOV3PYSqRnq1jPjR
0eNf39reUrq6iRZT1gOQrmEpdTWimwm/1RkhRbSUzPMUEGN/I+Jwp9QzCY1dSCkT
Pwvw0s1BT47ZewZh/0hFvo2of6hrlGECRA96THdnKkUntNMCLlWVcsLGm6FIeejx
lxMS3EfBZyItn7s/1DUQ0ZuHNfDrnadnVNO4DIvSQAyBv8Wauqr6EiQB3KtCHZ5c
pli/PsCuIEpXHX5eaurOtiMJVMnSOcGDxAQGlQkqRbPzR/A4Ajkyo7UkS7iA7CKO
te6DvPIwJfyS6wG+ZgnM52WfLK+NAmueYkkkXpOtzRnqoEJ6J9ukcMdSTsPqApZF
QlVN2E7crAKuyC6pe0knyiyM9egPjlG+h25mDo2BFRemhwrfWHwr098i2qo2W9VH
YYXvf15jGuddm7nvNlLAv2NHGttmxVNul1dB4TclrEIBPbIp2ajnJUNjbo1IVZM3
QXp4XKM1EtkAuc4XLvWnPYfscDQ9EOLRVlA6Pug6XpdUD3rB+/sWbEzWGcGE8FwE
LuxppFsDbSIpdgvXXhNB1+GtGgGjZh7LFxgYImQx9/rczxc0QKU+GuSldMImTbzO
HWUjqm1ifkpOcnSTX9+cwCY5qBRTKsgWP7kit1nJCUif+nNVkivDfuKc0lb2aKPR
7F4ySuIEwF5EnItdIkKEm+APXZ5N0LLLa+0ejOFDj8bXOkmTsAPdzPLnJKiEjuf9
I37Gd93pqjA1/YRoLSVd6k0HKxoZ/JpQnRuty3iJgPua82PsKZbq0W63GLR+2jEu
ycFdybuTJrkjpvBb7ZBfWTmOS2qf3TkG7quOsLVVZhL9elAJWFYJ7NvoYC4P/dm5
Miuw7AF+fxQ4snvyHTJPgYAcyjuMtbeBJI4RwyfuZkQg2u7/vIooqOCP4k3qWggp
DIo352npqueQmYFKU56bowrXJ5kIHHMY5WT+cra+BtVibzQfnkIKsScHCpWM9G5G
Ny3duVWZgw6NTuPuclFNKQnXRrIQ13wSLpy1L9ogEH+oJAHx7PG3E2DCyAq+dmbE
sCK+ImxlZ0YtcUt5gFjHnAr/rOl6h83iU4zpG683jmh7dT36h30wI+k5ZjH03GCJ
TbmO8uqcf4o/K80PYaex6I4FAjWCkcWI/7UR5NPQqZBJTNAkCZlLSUZ2arWzUfay
HGNCPiO5OGLLgvvrL/eSn1Khi/3H6LQ/8S6+psPmQYjN9VdqTSl1MYxvcg6QcMPE
1mtpXhGI/NZXniwiX0CI9e88ii2YICGIt2GFDlSta9tR6alZ9//Do6tvZoRfYYXl
/el9G2Y0FIPAiY2PohnatOCY832KO7LEj5/v5Ryv2R2dsAUimce8MNstLG5lcfxz
sjbeBlDLIBo+tELADGQEyvFD3u+qBdKCfq6V+lw/WfOprZ3M6XEyBbE8Ldo9TniR
/5NbHkcTRSKJy3YN3xIm6bqVXrc67o8XtQXiNTzIfzOfc/6yP92dUIGl+o9zoHSb
yHD+W8wpbJSUIWZn2TMDAJevFIJXF69akUhfs+nWl4uk9HFZ4G7t5uPJEsn6X1Kd
E+f10NinfWtTGQYEAGynqpF/eTtEVSfxei4rsWgalNpbE5gFYhN0DVaG8gybK4NP
Kysb1ep+OGWhvPcmhj0E0qQSPd0jINerUcNmUNfcsRUktYt7/+31lNY6/xY/8c2p
JPveypbsoBZ7hbqQJeexD7uvNhYOhZWuLCaytOd8GK4ex+duNQ3JWu++3Syxe5CU
LEOb2STeGi7Tt6bdkj69s88MVU6XF+Aa9wSYBmm0FKvTkRkZR36nyNY13SYixV9o
4dMrslWr7qkUTKOOTtZYHOWHOy581F/ZVokeqPk9AQW8jAOJBKwNFkHDwDBHjJmM
Cdfw5AGK5Gp8mK8xCS4iXpXU3rMbr7gnsF9cFKHw7oJt6BGw+MSbMHg8tcfU/aSb
iIAQ0O1Mc4ikPs3BoJhE0o+ZTARW2Y9COH9qOCB9UWdh2ktYDRszh4AiLVfSJVWX
DvQGsNdXRC+BXFPq6b8z0h8kooGrIQytm8+TgU8q8QinvXrtGjDNzeTYGTvM+N0l
CnXLcMAE4P+kj8rv8ep6eSXfgAzN153dnidxjef+g4QC1FnXPGbeQp9hGzCUo1mQ
fljytht3yTmVNgOd51uqhmNzbV93gZ1BvutseVZ/b/9/KrFDOQTEevhrON2alW5K
cQ5z7OxAbZPD0TLsonbCqyExPBzOw04L8IDQUSPX+k9fGlILpMDN6owCldV/6vwo
N4n3Xj3F+dD8ZEASqgKvsQqSMAUA3rj/ggnekeqxUprnaMxCylF/kxfaanE+31lz
s8oGpZV1PzptcNw0hdUe7M5+6GWPmkVvLLxPJBDN0Ymuc1I5RLYRHWOmwWygEy+L
wr5ddKvyTIKlw7H5NMe6csAx/vv7dq993ZvRCJMuBdI0i8yYY+03y6Ai2GskyrxF
vGZNmq1L11eMUQbB3WcEQzJf4DOQBmSI7MZDLLTdzDjpSbfySkZQPzoasTrVuuJ5
oFt/N1FurVbERh3K53AmIMtFr2GRe4lhyx5WdQyuGj6AELROyxCVJwbDanNQzHu1
Ql2jsZCiML5ADqZ9ZXyOUxWd72F/djWspyHQi+dfqzq5TS686Fl3rMlH4POiIaJ0
Z15ZGfW1ZjWtWePpTHO3CdQhpCinNwIKyzg4ETK4QmNFCQFBT+sDcMtJ3yyhVucW
7MnJ19cfCn7Rx6jJIPDi03grZvtEfJhl7gQyJxw2rARTzzjxh6xsZ862oRFXciiq
9KsZIdEewYfnKJaHwt6GG+sdg4wvlY/hWXPE3TF5xxVKFF3Cy/K8LVQBr5jJ7SiE
GfIqoxuqJnTrvJDPGj4oQut/Ddqam69SgVbQghxKaKD/pXPrNuxJQqn3eFsz6Lc2
hHh3ldD3FyAqImdowrnbFI6Z6EPRmwhdguWo3u0EZZC/x6/1aiWb8dX8yOIQRNQ6
U+KxLQaWdadFOeszX5DAr4z74uKs3TXGgwe5uImBlNq15sEbKMKONfsoYCEfiZJV
2VRRapPny48LIUUgWtMpi/MlpdYwf1WCB2i0yal/poxRcLo4Urh28ayfTBmgFft0
FhU7nrcV9MSvK8KCfelZxYZTxDhTn8wXEBIS0qO2TWGTNhzYpCbfnF3v5DjbGMPi
8BaVpSk8wTnXHJHuYzV0e3oyEMEwweeinFeV2lQPWhVkELJP4uq+f92Np+O93HFw
bcpe2yNyrZzp64CY/FYDzTY0pB81M1wys+w5ch4Y2BRYvQSnNcFR1nX8O8mzb9Zw
YSO6Oenaj8Izp6I+344D5rA12hshZcKgIsdxYTEFrPhv55Tc+uhSDepW8AiBYHCN
ici8YuW6HDqrToJD+8hxMRz63T5/rK1mipUWIX2/61vVdTPBEVmFKJJeZesndERa
CSSCVLORhCG136D8sZfRWk5axJ31Ph8skx9j3Btzrbw7Z06bcTpKtkHOmagmE9gy
mB3Cs2X+JJxwAco+iCG6/4zIl9IqS1qrw1ny/gS7sjAaqNhozhmrjLz9nYNYrTHK
Mx6W506GgC8K8EGGCgS5srCO5DweHtind+aFc1JFeyIJsoe60wdmvg/vOzXmFLkd
2ShZKLOn2GHLNQqspvdvjFeEtZtI2GZ1HHKDxDqvxKmfym6pGPxweJjYc6ZxIelP
GBSBLosbCEPNYPV+Y37/M6jKFNvbvqX9PvR9G4R1h5xgTc8JKA8ayDHYDYcXD50g
l0iQfAlfiK4MRhu9i8tjjOMZko8IgwcdjTpV8FRD7EKsDmbA07bxvcM/jSvoUIOA
65Wgw8eC3p7YrRtvxwOCzb0WpZKWc4rr8Xzu6SBgcaJTMN3Zk5oCr3GYMZrec/ep
UwzHn4gpaLqlnzjSVF8eBsOQnXEGxpAoNZYKDuRTaqllMnz9qMsN68bRy+wcQ07W
8H868PuNwpeZkQxGiwwyT65+K3hdZnZz158kcGPSp0n2FTX/cbt23iTBTMYr+PfP
wgtfeYWdXDLk2wyMVYpUb0ouAPR2xrezq//RJKF1pktpHqLwI7fHfENiztfcWKVy
APEzJdMaat5ahDCmZcwWyHFNsayVGj+Pt1oVL7MazAQ2VjY5kq5t/bCvIA5Rhgpp
kkgdjcDwDhfkYmNgDVK911OPRNweBxAyxZUZfwlBf54yXV2ucY/PFffSMcA0iTqD
SHRIK5v6JyXHyvr0QfOpW3p7yATVJXCjb9RrY/lmok5wPBUl/etsLHP/7mpforo1
nqYNQGdUtJT6meyGxBFWpENcbkJpuwNK0CH0dAUMO1b+bGMZXIPY50K63bdTZ+z1
yzFqEpg0NHpOJou9hqyBNb+v9BAFyyK/4Rw4zStBwrgZudUEvqNq/edWqpkdoTAS
YPS6U9hSj8u4WkT96BycLxfgdgpsaknfPnpqSOCfss1NpN0hcouLA+tNLJglCBWh
3FVVHb336JsJNxx/1Q5p26SDiBpv42BoAFonWR+x/5rUMeevtHvba7l/Bre/imoC
HzlxdiPTdwsNSlIslx56bn8muD1lBXGphv8xaRqR1OF8FaU8jJdfVUJfTEVIZv+z
AjAt7knOIM9A94GV8NMtQVrqPZET29JVaI5ve+f/rnxsWFafT6/HjdLs3e4KfSyb
h/vtzbZpjdhVubmEuuGXBNPXraqQb1xWDKRYYuqYI0ioCTx7VQ/mBOMhKAY1697y
TR/R/tCebVQS1u7HqoanrDLFdecv0CHkuL+3yDRpXpenNDaok4sE6LVkusYhB1ll
g6pmkVft0+XtM9u7irLxHqPY66hnHnwnLVAAf3ZkGCcUfgyRgdD4SHxVThItUYZJ
nYDH6BOc0+1bst3QSlKeRcTbutJ40ncg7kPdvkaBquU3Uggv3RT/Se0PlOjUS1Ur
vVqHFPfnSTKzLB5Bm7iV7mVUX8LNlAwipgggaiwSksjbhMvO0bIPCJrSYDS1PZ7b
+oVprEKe6W8FsCKil6RjKOQyaZOIlA1BfdbkfCLN7ZFpUcROLG0191GIwMUjIxfx
DBLKL1zcZU2lEom55CwDMRf+VQM2pVLgETzR3kiZaFkRMM0oYUYUzanSwNoTXsUT
1ccOcHtinSVa6O2adJF7vz3gRl4Nq+5Lb065yxN+dlGHzN9bHuJkEVc++UVxHpom
1ykypuTPQrKYvQkcJLkw+777DY735U5Q39kC02XpmROHJ06k3vnvNCa+WzjbjOGv
6HnVR9NHyV/2zTrGzZv95QcAcd4F7eEtQjZEKY9uuRsav5oEzz6gFRzoSQWsZNZn
PQIr+bGfKF5DsS8o19buepdaeogv8lnwFK1JYfxiw1HMXX5AfEiwoeX8PGxa5ZLH
DxxNzBfhanLYS6wB8fjsBaM2D9A69hxe69HeU2+61M6o9R5jlDYdjo40MaRRBCBB
RuklMC+bTpO6yLtbDw9dv0nMoOsEZmejmn3JqpqTdOYNs93y57zKU8oDWks1j4oq
MeLafCX8IW4aUaoFO8S42hWM91hHVb1Py8OjG1Y9viZcNMiiGhuILv2103q6qmOX
HenqK7dgrnqu6sy2Afkye95YC7YuDBDCGCTVEvKn1jpZZ4/Ui0YiyKY9KFvnP6Uc
R/zGED12NMZG+1g/q+cYwmNBGPpRCBEgOeGc0x1NcUBUnRgqANgdubWgNZtyUTsM
PQzneZX5lmF7ScgyRE7CGQ986ZxEfFkvIHciZE5MwBa7Fy32uVtUvNRrPBIcx0Ao
uK1Pg+6oiC+10bm7jI8ELBvIOnDrl7JQZhWijGELDDs5vKj+T9+GkTKouCr5ufLh
7rmopxLjQaccxB1ZWWv9w/ATS1WUXW1wVESmk1ulnVCLY/m71u2PpdxC+1YSP0H5
Rc42t4UqXx81SLYsvGlQ30Csp6BdyHZiC+e5AhTeGfUTfQdPup3O/8ZqEgmXldOK
QjTLaaZtO+judF0UIr3DFH+ZveCntEtktWjvtAXDNQWNAX2504M+cRrDYUzudgj2
Jcgng8eKo8OeVQkpxWKtOkW+WS5Cj+PVydhpfnQWV/zrdZBf75HZr5sUlw0puafp
CfyDokXHzBWAUbkh8xzGDNNG1Tdn/WxFJiSlEPprXuJRAVTNyqcb3ZMJkjINNq/t
CrtpZmb1ZFNI8ahj+Q6WkDL5MQohCv8Hzn12dBzt3kzBiBV02ebe5GOkwReA7oVm
skiIeBnLkENqQ1FZxKkycnFfD7NGl9jwXfCc8eKGbtZu3/RkpxedlJo0YNv4wc6S
0W3JBSs+rG2NE4l59Omd8rHqJD96UXIGUs/c8vWT0ZteX20mRQ+IZnIfxHf8Cv7T
rc5wdpWJDdEtyl11LNLzO2SlE031dFRAl/W9DpAjWSdRoNUQXlS1meYrek/Abark
Nh1dJXwZN/xuV6krMKIyoSheKoY1mrVBOcf98aML3iNoCB6V8S5GK0wpwojO3lTW
nb6agolANe/rp4XjxLNXqCqfspoL0464YfmPDyhiYJGLZYaEo8a794sMMKQQyK1a
g9v++9A0W0JE5W06OyOjvQCKJXz0LdK38DOOnvOJFKEkJnCWwKBkoxxYV48aiQIi
1tp503u2qs4L6JpNkxscT+zG2BxGDWX7hUcUWxTo/cVL7ADTcTnpN5rhj5qr/gev
p0+EuJEGSaSdV1eGF9AqMoOh60cV2V+Uo9TSxdNokLWImuyQhiiGPIhENr+WvVDL
dvXcKCTRESyG25vthbRjSPFqkX2pGx5wYK4u7hRacKqbq1o04n2IXou7schHl3qM
IAIQC8cP96KW53F8pnD08EjQmRu+P2sVjXbyDQLMoJobshj74VOK4vorl35iDkoO
In1wrJrkXBU9pgK6/z9w9f9fAa8L8gRlAZ9ZwNfQ72eH9SfG+PEW0T/LJjcSbC0P
3BblfS5omDR0Gsh4QUQYleo5vl+zza3tAcvSnBmgy6o6kW63ipIxCNHz23/xX74t
yodH/rS1+iP8kKPpYW9eLCuEaJON/zOYnmlriZiRBQGVmL27yNqVRPp0e5jOBXGx
b6s9+erWw8XGQ2IXAJMwi8eXMPpcFu6xn/Zl/dzqr5NAztss4vidr+p1pE1aLPz4
bgTw/Dq+fWWhLs0xYF7R2mtuvCKFUXke+z/Sr+tI4jgsZPmBdshYYRgwEtaDHqHU
eH0/TUFifkYeeEhHP/Kzy7jw1lD+UPq2ZvzrK8jbpO773kbR4Shn3aSXwVBosjPo
VsvydmthirNksGTdyC3wIOJ+ZVlGZpptiG0KdeOQoVMBcBI4z6xxXFwzqYa8TXc+
DQZj7FXSiSt2ARJHLQ90bbsG8SvecK7JEPQIzsMwPP1KNFw7bdqujrBAzMIOPkxl
8zIx/9mX8r9jdUJN5to+7ua8qr4iiXxaVP3em5HZqnl1sheDPIW/YxiI/aylaS1t
EScQKiujpaOk/m1MTgp7uMoGAyjiz3nqE55V8Q7ExsXhB8bXTSItYojcMuZE5NgW
gORXz2ghPuhbajYpbz+L5FEvzJTFu0Zw5P0qomyWhNCIsgiUVF6ONwDk9Vb4enpX
RlgP8iMWGiSrD5cJkR2AzxMc86dolLgxTVe2NL6VgS3+qSnQICe/V6Ea+MTmoq8F
7TiYVxMbI4A7cDu94rP5rSx7v4WZ2BbVI97WRQszmDnnc0PpGUDP7evjG4eiPSLY
dobJMw6KqUNi2AVDycTKGiswalGsZSNtInLGXxIe3w4BBsFxCfC5wjVcmRjsA0Un
nQn5MN3Q5Tt2Zg7IROcCBT4jMXB3GidYK1E+k9OzhbZ7QPAT8YTL9L5eAXYIlebT
NZGJbODICwE0zsItL6iueA+lD19rlyeohq9oCbhGWPM/M32+e/R5L6SlE9UWNrY1
pHyJAzpOxjr0rVriAeIFCzRxOEawz2IuLz1nPuXZyiCZD75SsNB1anY2AhmBxN9b
7nw58L4jPoL8BV/fip6/cbqmqrKKXoZV9rMxyTgxW2oq9nbomSon0+6yu1Q9kQbj
y78Kz11Kn8w4xN1mUDOSJwsv08arwYhgIk9UbZAS3R6G2dXyDw0dM25yM/daHWU+
mKG9unk3Uf6mrQJbvnhN6447lU0VSJoBkm3P+ut0uVwCd61ZXRQ8wu7pdOsHclAc
zrIkXHFEhF+8KihrQxU44rLUkUSGLAmebDi/8yGsR9sMbpLzyF0B9WL5dqVoNR3I
sRVfrejXtqiXMnT6rOW+uhj0iv57VyPYtDCURIb7311ZglTV5P0VoXyA5kLlFnFh
7/EVOZrfkqaK7/e+ZScu6x95faCT6PJ0ZyiHSef7DgkrAbCqm9POLhg0PwidwOQZ
f0T9SC/3deKdsUNLcs2Xgpqvc8s5rp5dCrsBTnW2447dkBqlsx6Ckz4EGw3kStvj
giaPFj28yK/pQ5I+qidvmaPLKZ3KUDZE7l3JIEKYnKqrkXhTvWcBPvsjRD4Ji0MD
hIxaJVB8/KO3TCvKCNRNgnq/U/UTzJybixPs9nEOllQnq5w/hj4tc+675xn6m3Lw
J2j1ssxLppfo+JSEF7jGg97IwTce4DCMYclLX7lyvnqzkM98ljvQmCnbzpctGvql
xnU28p/Uk2SY1tdnGc/aCUuDjnPBAafQL7sXbWNyi7uhRkLneuMS4o/eoi8uc+9U
k0tb69hsVfHvTR1/frl3LOHC0RKv285/VtiH3pHdD5Bqd3wOIDugf6Xql9lJJqx8
B+b0g4g6wD0j7bKUADJoaXuIqmGa2OSpuxkqEHMG9Rzvp+wGCuuZ+qvgPsU1aqOP
Mhg6A9BQXnDhj4bkNIQHACDhTyBcQMX6Hqes1U7gWVqfU37TAQzGbmccm7jzv95/
U4lPLQhxyz6DgAqtz+WQaicFtlmoS63Qk1pN6ReHGPQ/Db2psyaT47fnwXdrYVy6
zMIc+IX0zOvvJaBhrDcG5Gw5SHztp2UtWMNA1/jUpxYDSCbsEuXuMx3SBs37nvMu
fQugFDQC63kVvKLHsM50NNWT/svWdbbJj6hYNiba4C+lWDU/YuB2cTApmqqaNpXC
tAf9AVbsU9zLZslMDqVWMzeDk3wIXjHYNc2uYgmmaVskOpRBqVF4BLHdUhfUtMXb
GxjbBvVQHXVpaHeYP616nmZuYV1MH7p8rez1BtP4PJ/rR81nTBXbDSlmzH3R90VV
+2kZBSHSLPUEwaG/hsSQtH4AWvNgT4nuLbkGlSwyXkTdOVvHfW0vHbr0o3t6xVM6
05bqw+1NMeyyK1xYdoxThyhFzFys2AFoi62RAlvVY9ZH0AkVt2GkQSQV0HQL1+0Y
QVNIz4gbY6ufnB3+hpkTk5I42GiDMXlesLX6Hqtz2rgP2R5cWx4yvmHTyqkL/af7
Ju/l3xzcxXtoKum/utKU1UmVidzjv8O42/jje0Lu45vmiQFQZKjXYLTlIFpkTcc9
oE6wasq6TKOhGA382ogTtTHkK6MJz8dvxfi0ammLYo9gCq6ETmt7NmoCj4VY44dN
MEu8Gic3jZzLlGmlKFDreq+qf3hZlVJCv4R4FXclbLWisE79cwJ2a9WVRi6Asw69
zo4C2+YuDvV1E+Qr2ahgPy/Kt7w43fm+cTrKEBIkBt42vSRcu5rPpmtiI7mzO1zn
HSaQ0akvTcS5ZIY8MYBUC9eW2qGEfTflrf9XMjtmZmV0f2h7QNeiR4JTeUoba4qm
EKHPmtPoiLQ3od0w3whC7c68eHp65jJPhWdiAyz/fB/EZWd9GfBj/RSAL/CEDxy/
tdPbV31Q+Ae0zejKSpyjmI8NwyTDp3ldwPA/QxOknupBkiLLQhqnhogN0Syw9DJQ
7NmK5VgLIIOmp4I2vy2lR6U7POq3x5hm4ZLjaCGvibX3IyA39JZSkvmtO+VYbjaF
ej4pw1O9lV1GinSA0yJXFY7ZrpOwaiDCWrabb7YJSz0Mgd7siubfgvvdYglDGBSL
HVw3jsIqseBnM3q8ESCSHfZ1AS7UY8yayKSKnf8Zhp809w2+gtfeQ1w7eM221sjk
aYjKHRxV3Udp+fZ9xIAQE2pCJJ/moMyRzXD3/mvRjAzEsMR+GMlx4/3tbZYWHMRD
p/4YEgeW+yLBcNOpS3ATWpc4WuGCFJU+8Vxd9w1hnPko/sxYLX17OafstI8nPqXu
ZXgipVTrIUWitvQdrQSsdYkRqegDY5BvyXwtHi2yG5ghlwC2300nOMUEDS+/r0Vq
9QrzE6SJijhP485ZCG6IidPVuzoSYkmZvLgVj6sdt9gr9148eKC9Pc06xGFrDMxx
gzYbx3r2MdjXCtR4qOABBNCJgP4ERUcHXbhzq2wmm9EDwwTzplrM24Ws0yqa0g8Z
XLmLVyl69ipDLOUoQ3O1cLfmIuqnyFfDllow4R5kP/9epO8on4QXg7sEpqi3pXoA
ClZVJzHeLkmwpu5aDY/eZUfe3OND5k8wi9AcdQsrqqrL9Zl+jX1/NNL4GIBibtuR
5eaW4Sz3JvkrcRo0mfj6TjmhIWGj5Z5pvneuiSDbPvRUWRXQ1KnbMRyrQm8JjDLm
4TeBW2qV0bLSfBdrFYY8RS0331khkGIjbQkEVrKyV7bP2CCcC3wYkySPwGJl4rc1
X7hw0N10h0PYIUaCxrT1Q1nBls7giA5DHyfGl4Dp0Sud7V/qnwnxNERSISH8kwA7
80zDNmdeE1kWXYBQw77fhq+MDg7yFOSmK6Hqi3KxDDJGub+rUwpLnDArQQuopoKV
Mjei9sMD05Y4mel2ivRBUi5NCF4pbDsYsrgUyCfe3kqjg71pPtQpvPEr48MxGwHE
hG69f81HPwcjEM2hyj4NLVNYVf92RzH4dri2HCWKVlz0Lzzp6c+vYbSQZ5kndVy6
Nz7RgorY82MMQ6mD3fs033rC6GJPcfUiQImGF3VsixHAikVoxEWW1OsIMXxM9fPo
nUgNUbX9uDJYn8cfyZRpsfJyO7pop+RLcdst5zxHAkwhhjOMx5BbpB0us8hYOW4X
NeW95RxF+yS9tEzBFjfGnfZ8JeX13fgDE6Dz87PyWpg3mQiaEstSg1yWu0i0PoE/
nJ8M7+ieyA3rscDbRcu7mz+DxURs1PDSCwu8OeuwIXdu/OMk7dXdOKM5ip6D99yJ
/qE89xvLML/dlD8+qLDZXtGDq4hmITqHOyKf3HZyw4LnEFsVawyZTeN61Yt28hns
GJjzzkqTfbC94NyKJ60AZ9hToUQuO8Y4RiB2wj+IBDEZ6n0G1Ak8TT4O384aM6lw
RyzGTAF3/yJyihoBZJpwshUILJ2WamM7o8sLiwofY1bgY/Eamlei0/u0IXfeKDxi
KiZt0blBQo8jyInvstRJOo78VhubK+jbBMwb50WeyGU5peaXady2LPHEwwy+IPP+
0XkcgwPz97+Idw/VY6HBMFyiV9H8kphssC6jEtSV0LM4/j0Sgpg1jyBwv50PjMnj
i1CETdJXvq0l/vX9L3fAbKxLmPKlTKG2IWmGpBxT54vysZeRR2kWuEZNt3dnbTPk
zWKhmtuLdi+pvmA6/BQ9F26rtJx6UO4un3HH/KXLbEVxIN0IUk0hvz7MJqjVKuEe
qfknMpWVxwhbE/+ae0M0BaZpvtP7QiJmz8CljrcjWKLIcgsqsboPWGH8ttLQWDjR
sTnE5bP0IAq+4tpFaYTkYqEumChDZres87PeLVYVq7BU4e56UC00922XjnaTCOWS
DlRw8LsKbam36OFlRLi25bcfzrHfUNy7ygfowv5i/q+D6oFiKUIKX/wcEuA2KDdz
0M5qFP18IriILtEyb4r1S8Q7fA04OugKUnQZqEn6bBiY0Js2m81pGoPv9pn9uep0
+3aq8SLenH9Et+PqUXnu/IEUFFrQB8ZDsI9ZHa49vtxNuqijgi1EJzSsjxCGvmyw
kuyJLbSuOleaJAbMXmRwbnmYNXmeNSOYSXFO+eh77+ZoQCtd/lXJ2X7AK4KSPVKi
1qTwdce+W+ShRtFiJiMwOM3RXpru2y8ngHuQqjekoBTY8+Af26SodD14Wwb5ymvP
1BtIuZBQs3rkxKCYbi/E3hzb/whdodWauOSwCPR6WZdGhpRcGYfb2tdPOIE/VKDp
H+tL+XVtjKL+VtGMpPO69rpbOT1u/WwaEXdfAx0K3s7+c8z6Km9jJEpt1J6NPcpG
DwiOXFufZAYcK0n35/uDg994WukIuwq8UihgQvuOwnG+igAfC4GCJmkDZR8Ut9i+
mj54sZChoUHRMEVdZ8o3XTA58iCty45A59m/TMyUHhckvE9UvrxRsTn6aWsLCus2
WR8itvSOGcIJH3DRw6g9rhzOmFgU5l1J83ZETTAsrwyIqsJD473RtWJaOBpJCAmZ
0OeQAev9Tcho3Qvdqd+fhEWYE40hh/IN9RR5gJ7KvGf928yX/qEofAvk69rzXoNa
7cR8X5+j3Sa6DuP/TKfTNOQVzg3KI/8hgDKy5vuLzw4JBAOQHtWR4sqJ67aEPccU
Mu1ubZpug/grNtfbNVDcyQFnPu29n4HqEZ06Jp6pEWiNd+ZhSiTVGmfYdfa1qenC
sHI9lWBqo9neAQIUxu3yMtRS6IEFfGb4eEYwYIw9M6QKtivC7mEdeVlVtlpM7ovB
UnUCNWiX5Gc4GCnb8CBhcnetHNgZ/Vu/KYSLnL+aoCO84+E4CNVSBzsE/yf0GG2g
JyJMHJSBtiUKJLrRbqCSYlVgakgou0tH5uR6pvu4T3F+4gGbpTzVJytCQl1yxI5V
2Z03IY/ZVUSkK+deONdMfkLOigm52f5zJS0+paZgkD0BDANdrAiSRSS/3MqJB9rJ
RsdOr+/o3CFxUG66DRPBg1PuKy/TpA434PdobERluwPx+MRMNOM/C2AbIjKGjUU+
olcvBprumsUwGxpMYySuW1Eh0p31hzFtEGWMsqA2SYhoBSzhvGXF7gjkeX4btWvh
DaNkuf8wHuciIMFBS8aW4X/21hQvwx3AuNqvc/DmPQLNq/FAz57GxTBvw4T6O4i7
aJsWF7e4SgJlW6V3Q4AwE2s87tyxXNIUTO9kxBxVW8HwTMwOI1Af1K6sZN4548vR
FEMo5fF82iAc3N1kCPZWdeXNa8ROi0ArLTnLSU/lOts8D0jYiQ3a5CWA9IWoXvV6
AP4RpMO96i6sehZHMWlWS+zA/jhrA5GabOl5Xp/22PDzp6S3IQgp/GmkrDbBZKWH
sAXDCuqfbbFKDxhA0mFJjOlgBjCzHtd0NDvdJLIR6BcT0uo7V2oF0gA5zXzbLt7F
AYhf/R5q/tMjbFI3MehGP3gF9YdpK+56jFFmJJwEJ4Eea/rzV2BR3xaZlTn+FSf9
n4yRDJJlRmZO1XI11tuu3iGpQQNFou+Wps5e+mpeTdCFWQkPR+K+DuO84Uum8kNJ
wx9dGrjuxfNy5UTfQ/amW8thih4sDmuiqymOhtAfY7rZ0HCCdOutieN76dkIGBhd
CFCNjhZ9mkCZ+Rpj8oMOoUFnGeTChX6akDkTMzzNwJ3pjOJnvqfRaktdo87eUOSs
3aq8OCegBkNZ+CwYlJmgNFqwVonINh86NyTFNaGF3BkMJkteyN9uZMPXOAw6SZ32
JNQQktmwlSKQCQUbk5F44ntas8JDZ3EMQ4dGTSZJI9+nQNAPc+ZsElrjY0E8In2W
akXEIWtgzuQ26x9DWmYgjextCTtEcbPMHfDqfuquv3m2gR7DjgKdnMJ9P9NKy6UI
Z3A4uefhVyrnaFL5t6mQCTXy4fQY45NlwVJXs3MQhgwKLihbMOUlkrN6K+Y81r3m
aZKH0UKcxTbf1lwqWHcO8BKuX2DicNFvgiHertfwugNjUQGoxh6Dnjdk67hDJuFU
tA/HvHFh9c9VvA5jmOr0utPUySkkESho/RaQn1q50D1Y7UX+CGo6O2p1GoPNdPSe
5MdFnhfagP3iD1OgnMU5tpvIvhPtMYwVM8V3JTkwpe3Un22VGfNvNCwqF5FPy2b4
LbUkN2C6v49mjmd6z4gDcVqAln+6FjQWBbrLLONmMvs662AKmTkLA0g29volo/hX
QVXxNTfy/3E5o+Sh/znIminQT7A8oOdAhTR3vq/APjDa+sxwLamRM96/cFlCH2bc
XBvguy50dVlvkryPF+lMoukDC7JqtmMMU7XNJCZh4qWMqLJMWi79UixZey7c92pV
+AZwyd9+Rm6LIbijYGOFXgWcl3V3BjJehXAlCj4BmGhjou3t+uFDtqM+voVcpo3e
vPsLjpdhifHCs/nV+EE3E1whF1HUB6dLOZA4ZnDvWOZzoxpioUFISJlwhFeMY+QK
ZqCbOBgt/3+VACE7aMTEXJJJ5cQHIhz8LkhtaxynshMwGaCYlB5vZJRKZLCdqTLS
A+JENIIlM67l3OdLRsXtE2TTGxY1rQPwv7qiVKWzuv5B8fBE4do7wlJzVUv5UglQ
Aq57YQ+qK9vwOGyQrpToNN+NskJ9gzDxvQ3hSTxQmO5HCrL2vhEw+3MR1vnS0y0n
o9gJ+Z/IeKyfKBcUkdQexcIHp6tFBWz9nLbUPbUE5CjxOvOsVDTQetAyIeievAu5
fwEb73MgPAoAvwuDVyFprrks5ielMODPrRuezjcpyFYpAPODWhG54BkHy6+3IqF1
jxjmd3/ZrF7GqhBCGW04SqD1BoCjyowjjPs8h8+rIqnmhhSXrrJxercV6jQmuBkd
0UvqvM1lXW2XD5U8OcynhGQEsJzCTSnSnxPd7hyS/vTWfjtifri2K/ivMlr8qA1y
MiDAh9XgYsV/IJp+/xLMG5Ps8CISUQISzGIrNXKQvvYWFkTbRDsA7LIf8a6ISZaG
XG9fV7QcA+wh8Y2bD8Am/3vEC6/9tjq2lVWcy82kuOpCWu4agF2+tCjFcjiuXEQX
q5mZv0iXUfJDpFba1zrNgezNBM0+pA07YX5kBjGp1buD2dBctGKgH7IJxFuycqVy
j46xfs2ndlhGfk1z1f2jxjsw91sZYhMN/IoGn0ljfRBJyj09sCzRBio10fM3qKOn
Q90H0uACrRx36woKpC+DBd52FeAgJ9iqp2RbBUUU3awrJiWM4ErFrOuWcvDRi6ih
7X9zpJJKHdH8MkBx6aryC27KYJqvjN+TGqp/FCbJEq8EWXlT8obMyOrn8iRohO/Z
oIjQuWQFuB1VQUlpyBdLyJmqG5HS0yIa+PRgE5Go2D1inf8XqIpEFqgaZ/h/vtD+
pSIynrSVJ7jCh0bVlJ1XlYwPsMhd2jhpoi+W+BOUphKdt40LTzWu6v3ePbDmT42e
tj3owoUfXA5TKcc5LxtLVxcsgvNEdWeKCAIReOBGne7MZQE7ni/xgbOZagBFbqAJ
B5mPiNuiLCB/JlWcudMp3BIWDPxrpbFxaoi6DwXZMjye/6h/9PhsVj+kTYQwWRhr
enyb9NP5uIDYu89o2cNel4UANvYhWZWdmGBcTEfwqKwhHDQ0YG2ql1qjyWDhCHJS
jy6Gcv+Zj1WoIPtp8zYnxCnHkELbj/01bq4DHpXjEqEdLD9wihrjMlszP39w0rLz
i3l5t32nmi06quKf+9NR44VChviRM/hgDRLsbtjjckjyf09lmKpeJe0G4OGnufUU
rpCe/Jz2fJ8ef53wyK7kfZqIJujGt2z6R9+Ip0NzCsPHGVtKXzh/BlI43+ELCCvB
ECiGJt0SjvzzqcC1dJI3R9HRv19dt5Kf27N8Y5a0xXVEpe/D+h3rpoQpcX021qCq
6rdTD0EP7sSCuywoMpFGRA==
`pragma protect end_protected
