// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g4Li9WJ2+WWeuYNfA5/S/idgvnkZJeYbZYp8vnR/dSpfiopQm3z1BFLNubjDr5Jl
CivAv146csCDLxXGZX43WuAMzsm0Je5PHuUAhoDODlOZ94q1bCwJxpYsruyjI9rO
J3L2igVJvTj9Xccxr11gZpbHC0orAoC3AFtg8h+UZd4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4288)
WgmZxQxti440ItXwjTBlUEo4yiqvVcNhDr61HvLu+HSw6XxCur9WdNXAlPiJxwEZ
K5iym3qERAQp+SXh8Tzr4yRiSTtXx02v0jPP4hluClfXpKV1WpORh5X2Xkz2jhLo
2KrdRegqbxmetpxr63Akt2UVJn9mZQYJxBYW19LAV9Pj/l/2GlqNg7dFH85O/Hdt
4YtzWH5tDXeCR4lylHgD9XqIH7xnwlgKUpLIbPohxdwVuhUs37W4v5Xu4bNdLgkT
a+waFiZKM4+32cKN9H4HmhwOPuCrvYKPeWtciR94/1m71/y7YC4Fddg6F/GbVlue
YoW+swzMSI4QZMJilXl5bA5tfDMt5jk/7DWXDmc1SsKAx4+L/5HaUlg8rzsBwZH9
ACU5l34miDttM63IKgrQk+btrbl5WJpWSwx0o2Fo1BwPJltYXG8sSKriULG8UQLO
CfNJTN2luX2Bx77VO0fBcZ4+YKlRCdrBGLh9G8m4+3FmyDSiza9mq8gUTEyB49rr
LgrMeZR/hGzf2Fm0dCj7ZQ/87VXau7odtqnyR5FUnCAOfHdKPMyN8l2z90B7QWT2
0Em4AyJFe73LzaGp/ctuIIcUyrpI4Nzr9swUMDXLmwSduowdlYDhryToB4BICOVy
xpWJbSaolldzcvvDLKq0dH/qVrziM/jct8X0y1BeTIvXYUXUi80GL4lLKDpM6l4g
CIj3eB//bUsh1JW3tE4eBrD2HEkV0AN5HKZkF+1VhzW6ycTIL+ehu1cEanCn9myH
+aA2kZBloyN+mjJR42VUmygBJekkQuNxDfyUsE4c3ikjyaMH708mLOzqPAbWsNoR
vmfXRSQ19CbfGBy5Z8SzENACB+qKn+4HcL9YE9MwaLPLajH+fJgRnS/OVX4jic3W
7ZUO9wUI0MsJfFK5cPFzloaKAXfVCl9aTX6vkRVDZ7TGYJAOg7Jfk1MEVsqI4c0P
yCOxnxDWv50ZaW6U+0hadoeMtS1lPIjXkp2G2EfHpyW+zpcNv8wijaiBMLGCMboe
sZ7C1UMm3q5eowCwtf2AOuRiLWdeMC/2ASwTVecN1UfQazaOBsDdCzTFxZkEVPdS
1MxefJQLfml89A8uTTGlZbeegm/we3H0OCGPYQg5AUMa4RlwuzrvHdgENH3jyrin
gqv3hKVKf3rhdj8Hi+5BrbU6seIIHZo4JQHGMRD/Fhnca+V6sTPNz6jTJSrrO0o6
D1Fny5Etpl8P0dSCiABd8V/+K2D+/DZY+sYOoScKzxOFGYGfoATya/dVpwQ96mPp
hKgIAv68kugzFNAmIL7fuwxB9kDLHgq4xYi7Ymbg2+/+qXOcZB92s/AmQaTs+a+Z
1guGDC3PmziNtVKzBPgOxr62Z/l0Jty2d9V9ewk7nB4Ew6SRUMZlZFzRv+MaLPJR
nfiKgsbOMG5zuspjEkN7iapkwx41okk3XT/aiT07aPa9G5Jm+di1agvs1eSCPHxq
tVUBcQlPIP7wvWVE3CKPcsHFTgbXzZRoQCA8OBIBYKxofGhcgF7mk1ryZfiOqIXA
FCcpwcSaMI6hl/1r3kYXPJqzU3TmIYsgFS2J/AIV7/UFp3wV9uoDuVAluoterRJJ
0D5IhP4Sc0q2a1PClhzSBe4x/sKj5tB9F9f6b90HdoGYVl+3JSDS/1wZ1c4Z8ax0
IaHOr3kkfzZsAISJR0YnPsA/PuZkVYNSx/V5ZTHk6btiCyoTEzOXZ/kWu+/i5GKb
wC6HRH6+qlUrabzC6A2v/Vqt+Ea0e2kXoLVE8aRpkkj6U1kZCrWGe5J89su6+rOC
YwmU+EesnTVNnBewk8rQDTn9DDX4OBVnUc6abg8frE99zb0bhPCDWFocpYN02mte
Y2uWlusx8zp5SgD+zm+tSo5rYN6rh7oKTHVhVaCmN02yqiz/IECFwzxguVFCQ7xI
NdF6gyEg/cfxS/F3SYuI2QeMAGjPMoEGpFO3i7uB4b4SawTN+awWPbUwLdNMrAZJ
Lk9Y+/0RwyZ6Ys+FGF9M1HfD82sXHiDySZC7rerfTKpa7SpkYPh+mozoFPTNNbN9
8VQXrJ/6w8l6GddA214S8yjBXorCabJsN13EzYthRtT+RGuoKTGwh5iFA90RfgVI
6/6T/HNxrNhpEE7bOP/01H829769pGNbp9N1CCb9SoZoxs0lgEnSL2j80MmJbtG0
1ucj5ajiERw8+3Hf6U06MDMTGEJ7t0kTIqHt14EnY3KNJDZ874HpFB4ho6c2RDDB
2Qk6Yrwg6QqB6cfmnOm9lgbpnxoSEnPWvfyqRxspDqoVbkH9sUCd3rXV1WBCkGt2
O61o6EF9KU1iyBoRGAZATEigOFvsVUBx7SrYFlo8DgrFewjNQf7fE7ghGUPLKZfm
K99N7Cmc7510U5CVHyZzVrha+0aNPFi5RkLP37b/CmpQq7BLwh9YDRfcY2T/L2XN
YGAyc5osEMSoBawkDFhRV2+VDMh+Wh0FihSzQvETHGt2YN+0dy+cSF8hFIZNvixu
r2gRwsl+svRp4h37yI3RsJD7/dEqlV1KlihlI3JNVqsbTRZM5jLN6VrCiVlBm3wk
40LRnyQn3H1rMXRnHbTjVQ+nb1rzBI3ynSRn5tb05LsQS2UfqiulBzSQGtwpdZq6
ue9coLibeO+26HdzwY0aI7i2gBWPw+39ZHKs1tyAH22AmrhrHC5cKX42fTyL6E9T
3Gt1S2jU3d1XfjbB1vvqr1tginzs1405GO/wrrzgRyTHrxnKKEtZWODL4HSLlxVs
JQt3iyo6eiNku7WeXZ4/BT3+M9ezER5sK7hNBJwbc2cdgTz1IZtFD6270X/2n4fr
lVRgKaWx3iTAdi4N163Jr4aiZdEZT59obHdfCdOI97jMR4MUafqiN1/mFIn/0ncf
81eECjeQMg0sUHOehv8fA527HTUcGU9fu6MYiOoSRGj2iHxA8FCAjI3HFC538rLA
5n1nQs4z5ZWJB+N3cyrEJzTSUihPM/VkrJZLPYnDWgyot8/Pwgm+i/E/TjXab+Zd
qBHtLXQUImjc4yY450zR/YkemEAU1S2I3NPL901hoJGpuUKWNmcmQGyqD01zzAb9
W7Lfb3Lyl8VKOqLHvmliMTPFSE6ZMXEYqN9In1toeg/ZKL1jsyCfdVv+E+QosUS7
f+pSeo0fOBodnbIrAbNbeikbv0CR2GI+iVJw8tVm9qDzvocFS2h9zP2ufm9YUIzk
T9V4mB/efJMmklNTCkAecUcvSgNugrh0gj5zTfuGhcaWBjnaAnoqFj7PnQIWR/CH
vQIN9XvzJfvKX1Cqppd5yVOw0sfPdXv6y3fUYFrVsaaMu9kHYpqfHbpxNhdSAEkB
m8ZFze2VdzJdfNg1uHB+1cZjKIHx+4jwl4ZMw/ca3wDFibdkY0IW1vCPk4qWT8aV
fMyZ/TeAbXftbsEc3GOflKx68LhFbUwl8otxxWkM+wlXHBfUmeua5isN52GuWPfZ
trbeRWn3e2MdBudfxrhFc5NQBAksCeisVYqvXlQgrdMTuriBCdqg/UarhBBS44ds
MJXQzw1ebKpK50flJDqASTPwfZrYUzvqO6iUdTl15tfX86Zpri7WDVBdVsaZx5fs
CaJBvdTQG+skylnZ3T9Odq1dOSafVEdUnxWH0JJczm8ccwDco2dPRf5/GSoj07Xd
P45XXCtS2Wmb340fXKnZnUcGPKc8bqfPF66ZHsiH1qvrH/YdwHlLXIn4M6fCEAFY
/rz/5WTkZFRLXdtCt6d7pUAPMhpZtfqlVY7PC/7nnH0CEoV9GnP0StlT6yS3jsly
D46SHeXcv6fCyzTkUL5BzPaPDoOP5SVmevecQ1Qb3CPt04sQEfe9hhn9gVGAxfOd
dkjF+bXtVZ8C/zyD2blyDpJ3kXYtUdtIn97MaWTm4izOtIiZuxt8tWhI7901lX8c
eS+eRbR6+MBJX1Fe1oQrteVnQWqXEPJ2mL+3iJgY1qhSdIcnvJLtot3fOhI793cF
Jl5SFqzVH6bnY2O3pn/G4DPhKBh3deBwTwU/Y7sWpVK0H0xI1xPZzDFYRld1ABKh
i7rCzhGBQpSYIn7+vmsHgqzdvSKImRNNTGOFxYYacTbENjXzLrQz56TyA3sXB47J
KXlo2h9Q4i0aenlBE1ASB+3RFcakRQAUkWkTAS2CFFcJadPGbHDRSF5pDAGh5cwn
Hncb5gRkGeJJikDj2Lg2+wEKiTcbROHh0y+ps/zFzvoxR5Id+qoq38IvfhneKoWH
IY6gxbfF9t25/rPBlju10bRpjjF+o5X5AHKFpADtGxfliZ47kegUPE5/EFewxXz4
xvPWZ+g9OBRCqGItyH+FkgKIsIjFtM8u6pCXl1SBxQBox/vsBUi36A4lsln1vYiC
hK0FChhp/RyzO1xK9aZOLb32NScyI3oXdQeJ9xO8ix1zGUHqTgytOaPVQrDQpPyC
LqE1Q8eGb16Uj2eB83qknFTE1whK9g51CVcJ+XOXCnp+EKTXkYACFUwVNMtzwh/a
6tVUKCj+XF7DhjXG4CRiv+zVWLfVSOvGiWirc46HS6qZB9kkd54AuORAHrFQCq4n
0QE6oiWvIdCZpLmSruBCgSrDmHP8QVjj87ed9KtYkspY4YkC0bDcyBjybM3/RBgW
jTUf2y2THueUASo2/gc7gniEwVOie3HWpVIqNR/oSVvOCL8tr5Y8xZplTePq/L8G
Kp5QMnM9PhLCX8n+cW+zXWLipAn1sntxer4VRjY0A2aYaR2ElJ/GmjnX3b44ltND
3TurzvKBU5qf1Xk2wqweEN3ckPCeaInshrv0jrn17VO9tPtccrcuFVknsUHfDxP0
yW5JTzXZiaPNiBcdvpJ29s0HdMmTpDZleeBVk+f1A3QTk076c78wfpZPbQT5j7QF
8K9Xi+gzrhZTt1GdPoCoFvLRHFxC9PFJnEWNtwr7W0RiDYagOE9hrXzW3jqbmllm
P72MZmWlRMHqPSUqggeEbnzZYNasBefwPjgkcmepxtGWL5Up1dQK7FrnfCqtJvxJ
fPSrZ0LyV8BVF5yQK9ju9IvhQa8gixHEtPgxaIUb8PUgjQv0nLUvTobyExACejs7
LtOZDG5F9zqCSEeVS3yrroebbfzHIGMcbjeJwGqLeZ7XUEIy8eXEcEo+7iSpdzYt
UeTiMMCFGiv0qehrSetBY1H4HXh7Na0rID3ZYc809QOlMJnLqZP336dREVIh19Hm
V9ugrLYOZrNlmhDLE0c8kFwJKfWhbegIDirwnvCgAoFSPFfAnApv0nkgoFSuSial
nmDYFpxBPi87Zk7wnZV5A50IzUSP7Y4hrj9Nb+tqCfy/X2dUGLCZZ8YwFRK6vKic
mJQ6bA0OBIGWnqRge6m+kAOY8Yuh4JQGFd7IueC0cYI2TsMNyTfW7ri8SDlETO9Y
0nNWSXwn3qsHjGbdDXlhb1OXYKZH8JOhkWpvJ/ZqG7swv+w403JYKmwDxo5i1LZM
Mc1VF5su/1wlGqzXO094b9R16iKfmbSZJPz29QrXhNB1HdxAgWMNzFob57ThSeDb
FynSEDl6nGy4M+QhqNyJ5TnCQ0S4hL8AXyeTb0AzEbqfMSsAChJb8w/nRygpC0V7
76JCz4AhtRNs27427NHnx0KIHz3SpL1ZmrmsIIS4o7uAwFV8S3WWiju6hPmZ/UU2
PsZzHy/ieb2L7OdtJeGZeaC6hp+fkJEjSOfGrsC/jK8R3ojNJo0l4HzTRTs+50CC
9ai/yw4Dxjq97+cR2Vbesw==
`pragma protect end_protected
