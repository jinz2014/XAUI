// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nO1ON5+aLQCJT3zAJubm6OhM16MYc2bb+Ollh9M93GBXBUEggcxAPCVby3V9F7eA
Cfl4bFzEBISNv0sijLS7P7Kv1IJmMlztR0IiXVL0qL7OME4+UwuWe2FmMSOYCoId
gOpf/1lL/+/bEWe2nk/E7pmoj4dERl1XvwR46MW04R0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21360)
cXDd+/5FJetSZxpanrmaI+GJQzBR5Lr7BP+6YzQ+/Xw4Y8yVX92mteTGQummGeB5
7Oo/Kk9KbWQDy/9TvUHJ9ZghC+zBNd29jDp3RQMTNvG6eHwJBcWJQW9zhU2QR5TH
rd0CTbGKYkjnQOAJB1/V8/InZK4l43cnxEV8fp6rbP49cVIivoMXKLhh7FtKcjen
097w8NPyd49+f+7vTDiCvclv/62lUpy0GmJSFYpopbchvyn79PKvH8POKlg4n/Do
+tdGCnLiAfEdVQdFGPnDjoWu/G2PCYqkJSHGxbs1l+gFcfvrLGAbqj4J26Rt0Vxo
D8VVjcL8ZaLCQVRKERyUbtGFgs6QqZykCS3L6mCFwD1OKGrGBU/iQqlewpWW3EXh
cjXsrhcraRgvCXaupH0FEFFZBYrL0rGOkr0WYOopggezBhFt97yyQLK3AACb0awQ
2NYNfdb9lYQkRchJuxAh+fv2nC00P2GtZTy43gBZNDMU7avF6kpVZ8ZCXo6purxp
uAPKEmHOr6RcXEwGiU+yyQvK/YSgZTzZjBo+hMcc5WER0BO6jYfvrBXqW+oud80I
dDa4LVtQy8pt3REfFT+K+wDX+Xh6PlmVyKOCjSsS+y0BwcncQt6sP2so54csr6PV
saMvULFFHstMKwIFNeF6L8ghqiTHxMOnGpmzaNyf1ur7hC8xdYUvlFMlSlFDngb9
jTO9NdpfIMlxrcusaCo/CFplPzqYQ1Svbflu71bhvBOiHrFergMOaamjDzumrtmT
JeDQJ8voFhT4dPIMPlBhYQjLD4d+inEnipYYut0lWaWf+4y5YCE9PH4jp3QizJmt
n6hWFqKAlXbFxB8VxD5v9C5UEnhxlX7a1EqObW4tjEyrZ+36zAJblG2MKp2MP78o
BhAshwKKw1PJyAIgq+32Vgj8m/Ibjiw4thLjmfHwMf3lObrGk6gNYWxJj40TlThC
0ifyGfxiqplgMx1v9Ok5WoEb7ZovY+zcah2C/82+ZVbTroqlYQ8ix4KkUnsy1vcr
Cc8ZSVorVf3dwbHUClrgaCnF+E6eWgB7ME10Cbh4bW2phUhe22DDbFZvdaKqQZwE
rP+/DkdZ3Q3G408RiG8vY/8hOIMuoH88yHnG8eePPNB6yr+wB4KobkRJkApM7CU8
2GWer2FClxeHmpP52gYDQqIXrMs1S3kK0or2a3MhRbAKgFU8S0xh/L1/DW873utD
GoaMw1UCDI7m5vESf2fXpYbhlclmf6q2HWSU0r7HRbW5FqmvbjUaQxzFeoeYihjc
AkITuzHpPVJFRMkEBbVFbs1c+6YPqnBFt2KhjTS8uPtJ1czv8TJTJMGe0jNq3NR7
sK4SHmi82OLRh75JQf/iHhnjAxekBeq0vVG4U24CudLKvp1PnRwbJVNZF9AZZs1E
eNsP7+ukVhLXLDa17VXA/yfhaJSSlMg6zg19iSrvE3Z80waagxnAGuQOTlXTaawT
6QRH2CyhsreBXqfqvgUUKi/1nTH2cyzZXF4UpdbzumtQlTQpzxUlqzOCVF8KCOaU
SQ6k3+Ky4lAyS26NTViQ9FqkHDxVZ70lP33ZJrBzBKP7OWAJqNzV14Qrj9sYGz4g
aOIdT1kqyEikaREQ7yYXb52czof4Yt5VVrtkQEvWKBeyVWG45iDwd8j1Tq53l1mP
dAr3726DCvnWyjuGVLLW/vZ/tdWbqfL9vcWuRdWiPW6XdqBgenrVfzZJGbF0pLyS
tmO1kHPPQPagvV9X/EtbwQiB+XUEoAbPy0Zpl1KdTV4CrAEjz9cdounbKqCTrluJ
KUyCGE4pZfI2XSTsrDXvFcD/JtzKNMldrUIvrUQgHx72C1oNfIOwyayPCDQbkxeI
SPSpBRtrQMUtCVJyMIZKYozr55xnVIDW60qvE0zt2G9FSzGwbM4c9N2/MnUqDnNQ
m6ajmdHw9mcPziVNQEEYDUAtS1nQov9twpYmk8H0Rok8OIv2K3YYYQn2JWhA+Hjy
AKCIMO74IeSpWOfs4g/uLrfwti8hf8oRI8akQv2k7cFhP4EL8Mgr3nEOl19WAV0q
jUvuU0qHGXACUcyWtbsb3BbItg4pjdWRgjYPNsBuPvZi8NMirvon9YpWj5M0LHRX
f+OfW8WF93rhfLjL0/aDhkDlqNBUa/Z2FDh6W+seYs9AKY8FoL/8ZzQQ/VCricuD
tGXvR2DZNyqzuuJAflbF0heEAdfgRMQcbWEZuNHyt5WvDV2a/35VWVRupt3LccqD
WhUINttid3pI+VVFRrbz9wPRIAOAbdexrsNWG5UP39dhlJIlokWMips8JEyRF4RV
OVcTZPFBHHldmDV2Cbv65d4XvewqVH8VimvREZk57tBOxIpPIzbX+I+64f8Nyp5F
BMZNpPqT6LbfUWe738Q6v9+xtWTw6lNWomV7Z1Tk38fZM+GKsYaGvt4KjQY6GsLd
zA3mAgsLNxK0kGfrEw87gSUSdbBPiF9eRkyOk4pazTBZ4s32FdLjGrrNQ430fVpJ
4CBW+YjtZjh2p+KXj9fD7yks4dCtF04uKoKicRAbBM3IDZE5HkRkmMqr0dxNW17y
JBpYxU/qABWjCzTk3X5MdmQ5pidBeIEVWc2X0b3uabcJOiMIDX6ZG3mPw0PgKvwU
5XrIDZAYjkZ3MEUgyaAvtm3Zn5VJY56ZQmhNeO0MwO5r3E6q4F8Dh/fWdn6bgse0
/0N6RyK6ixFrddX1ST58a2J3ZnzoVY4/zPhO1oFRq8SufQFt+Hj3hXz2IpjN4P55
s5gCKE61raNwD/qZLJX+p7GiQHaTWjODkztPliYJ1pXo6WsV6KUK6mCDrDghXiRU
peKHM8kM/vVxcP73pZmVKnbvCj3dhJro94IyyVzeO5cF93HsewPnp6eqNbjo8chm
MUbsoWa73ML7YXhbQxv6XLRenTBNmkzY2q05y6Q056UFBUwDGJt5oSop3sCi2koa
QxhuU0e2pthU3DV8FJnJsMOwkLwVGtKVfj/Y97GEUG1yn9P7OyDH7xXi8TWxzUjs
EQ2g+FoD1gOti1arrrdfsga1uR9GuFMxJPs8VYbDNhQuy5QCLxp3075bhnlYrEMe
jjIhYUsG7Kn2K2iQOFbBCFDnbyz8iBLktulg/uu1FE/xKoR7NBKpHaK4whUj+3LN
nPP0bv46azOobMBGp8kGxT/jL1NwfRO6QW/58v2v5qzJJFxWaDJZiEXU0ouDp97G
SIan0+zNOyqYaIJi+hIMfgXJWwdJdk8XymlvpEUswOAiCZZgJ550kkkk/MKXALnz
N3K2xYPX4rcE0CxFXIQAJXgjcfrLIqBq4UiUNiWj4TAsrut1NS1xnw49hTa52Ann
Fk56tPaOqcRq3sZ3IZo/Ijd7xdQoMT/rDTWt1U40ubOMHpciudA8K0VZJzxjZDwM
JoOzOxP+GLTDzbJn6BXedFivptkn7Qi0GcHHlYsK73x/vDYjE9BXzd2xwGSayLFe
ljVBGDdDeyyDjPCVhDk5JdkwDoyRmCMobrfoRN1mar1nV8PeLNb64P+tBbe7zWJm
to9wScaGxEeRfo1vy3D0/lXNxwslgTh1GU63v5JajI7pFdLYSiJ+Gxx6Qn11/k2p
DuqEmvchM1QJWKOi3CrOMhRYteg06t0RCaifh0WgbvRz9oAON/GjmJW2vLjdOkGx
EXlj5WfLgQPRJGq/KCIdJwwoB5XuxslLAjKqPOM5toOaYbWgpSKyANfRrqVv43wn
hLXCIolP97Ewdb489vZlZaH57uXpgHryUgvCNqGE882dOkg867TzHWfuHAWEUGCH
3nysyXk7jWiX9+rIoxQiQHx3JM/mVA4iJcg2JnTfxuwD0MM7K6TbajPd8yXMMdzJ
jinEoJNs88Ta0qNmUAumaeYntoVM1J9gMBeouO57yZ/svZMiiDr/Eek8spAhMZQ5
Jv65pGnJOf6NBp5XI/eeS1D5bSyhPJob8IW0JoI4nnL8SoMz9jfgzFea89CQDBRx
9Wd4ugfmmJdJEXb6fTMbb3RmD1MxtC/N4va8+0mFm2GH/ogA7baaDkd0hzQ9S5Yr
BFeKPzTINeOoV66oEraOyh6Ne9OZO+sW1S7Al3ODqLFF+dry8Zin52LD6E5ZGru6
v+B2kdvs/yVrKO+KJpwos6WYEvrJmTFecdhSEb7dRFLaks4HvLUSbQ0uhFJzgN3h
EINoQx+VR7mWAhC5CsK3mzRH4ZJmSsNVGEzJZXZ1KAVWNIVu3aIhtT7WpOmwObyf
Motv9f5CwbBsvnwkcD1wSjrLcKF9be9LipHieyijDVg3rC/QCgT1XXjDLSzddqty
QMEE/pmNLUni+Axj+PReNBZ3JFYGSz1t1/Oddz/LZKg1ek5VMiPj4R7mhw86KmZ+
BD6NZ+s5pl7ZIxyzqOU4kYAJHOT40A5Nsh5NZbWx7kuyqTYhW2Qw3yc4syBNrbqF
r6jgo0l1C2bDbOrTCkgsTvs/dij6pgXvDILAL5U1yBO6ADCAIsgoxtufr0Yl+Fcg
37pJYonIKfoIiAd1IqJODK5OH+X5I1Qa+Mp1ZJFaNkOlBAQh5KK3k2LRjTWNTbSX
zOkuplTiyq8VAxIxSjqOmpY3/30jfmzVdWLu8IVAmhgiAmxMOltJb1Y//LNyBI9d
6/+iCw/hbQUu8hMvzAL0u0olj/BlHSfa5bO5/PjiGCNl6TGu9VQK1V7R04tDc94o
qBHB6l9i5AuW9RsgPqzzCO7Kftq87SiF0ZxP+hayiCHIaO+CyYXKBwC6el5KiHFw
1sxAJL+eFJDQKNEEnPF19POIBLb5RC+PWddW/pvIbruJ/uCrTOpXmOPQR+GVD4uN
9cFApzRoJWrCz0PLiUX5zYxHPSS51i6jJP6rQ2BD/bkSLrWTMpUtMFYGnPIJx766
7hiANXcSoG+AGBJXxYze3ejJ1aGNLbDTbYkNXhgm5MGUpjV5e9yCRhdLTEzZwHKM
mmETdw7Lagf5lRQYgucYXrfUu7gWXFfjjbCLx70O+mX2d5qKdtvp0C6R5IsYeJSv
WNaBrmQmJMLWqdl7gup/zqHcyA6M0JsCqHtR3qUe2lkaRazrzy8h9TQkLTm4v1ms
U4nD8KAiZah2ed6x0rbweZx09a7i/ooeUqIHbwINRjlvIgPZaAroU+Hx+9+pvHqP
lUZulJqvqIIp5G6k/INWtYrHKmtuLg/aSwPtHK+xYH7V9KPihkgqCZCVPUNc5KPR
D//sqXpWLLIPtlyIp9mB8cVRlekBwNy5Qh+qp48kR4vkXguEyMyQPRA8bqLXmGMI
cTzDclaqpHe0KWacmqW2wFmLaeESHzreWGJCw/ef8qqZBRA6fuHWpcPGjAs8IgRs
at10geuFiv6dc/clDS5unNZoIGXTfiX/+aPs0qf3BDnQaToq70n5MCKR4ugsSmJB
4b0TUlriS2FGlH7Es2xNahYTmM3xVEr0/jC+ZeTakbUATj5QB3Q1G5xameL1kTI2
Sf0MmMQboXjf8TLxA5+nCSBfvI9R36vtzsWmESZPSmXaqoSGoW8rPoypxYimLki+
xHr0KW2vv32IXZgR9xCFoiPItl9ud/00OgFzQrgrbD0p8te9t4eR5S9x4ZfARnSF
I/KT3m9iWduYx5ZJaltZdcqvmZrOqCRn8ZCEc/k6fcIo8f4TSsnGllMfcdP7TZCj
Pvd/3A0u0SkdAIE6GjERKTxN6+EhmXb0MSnsUuUwvwnW3pBJaxmu4r1CMlHHNiON
kzQR0y9ClVO8AUUdoVwPjxMw3fCMTUBldUF4jjlbMOwYztRXFyFILvRwJ29t0dVA
HPkWnGbW0OSQuFqiT9Csy9QyvAFxombZ3Wcawg54a8zHSrKc9YnxMD4xFyPTqRiF
+XMnoM00Jnvo5QsIbZzVODRf4M0iDb/qzyQIgancvKS4cI59NGjzxjZcSOoUzy+x
AfLCYxNZx/UUzQlLuQDmn9Ahd3GSm+vCgyhvM7uEqBsFRKiLQoTSM7NDPpYBOt/J
gCenv5wG3WmUi6zNWTNK9wvi/nA05Zv3nJBz62PPfynbs3ci5bOyssKSMAVVNJQw
3XnlFtcReR7y80qmdVQUmRDfFEzPRdicqH/g9XG0o9JXo2BwQIivfx+soCRNHg1U
FXy9BhFbDJoM9OwBxTaMQYjlxjL/mnvHaNGGoZuphhf5+cr3nEPQudxZZePeXXW9
qmBucSoF5qlwHIjQsnuy8Z87zksDclHC1kMPu1uFQ7fmBcg/TUM7G0yChB8dGG50
3EKjulFZNaL69lllWCGMb6dw/clKC0V/TOwzloDO+9D4pJx62sCYHNllfWKZP980
gQ5uj3+oCpgT6/Q3UONpABtj7uc+P6idT2yi2Z/ZgRaN8VLQV57L3bMCgllBkMc7
u/0XuYMDpwUlurc/omaolekN6hm/4B8Ktyry51C7CjPC92MmHa5+H0TFjVz1Dn68
3XiQrJNwgs5bIWO6LZW0MvAzPFP2CzOsHaaQouxxgzdhdIijh2pfDR5ISMBANayr
OS35kFZMYB2enFgWE57vs7YTnkFTb5urJaVsrpqUOpv3ILZgG0b/vYBMpQjIOQB0
cEO1H8yWF4VLLpNiLYQ9JlvhptQHX1nHx6VMS5vh5Q81ydS7C8AJuNoyHZmTvK7o
tkfjrbpiNGw+dk0gZHDuJHDHTVEleWGFBDPq9TVZ3P4L6waqX+SW6QKT4MyD2rZp
cteILzuHVXyBor5rQ9/FKMsPYD5B8u0CWmZQ0Ty+CawnEl8I6TgWgZbmOHYtwuA6
wt15l4/49ZG0q7ufg+3fm/VwTpCgGEpQ04Lu393NCzdfZR4/wOwb49NKzhNVSrZS
iMvaO7v+BEPkI2bNAxcHqrM9/NWvW2MF2Pkj+vvpjYL5A5V5vZLEdeAGNf7WH+4E
JYXEgKR8D7Pz9avEXeO/wKhOiQpzEJvN6FfbxSlCCR59Kr/kPvpQeYj92+XWaj7D
rEU3VFhVUZnsUFstym/NiQKwtlAt7eJ0Rqjyv0RhDAkLrGqJ27Qm5cOK3AaIysyY
0qPxe1RS/rNQOZjIb/qbgLjD8T1PkgnWNNNFe9irAIPpmnwc1Vwetrqwcs1yAyn+
/1InxTiSYYsLjqO6GO8vkh6AgpL/qWBlI0QIVwkpk3qeDd76F3vB6YCBLxLwNC/X
+PxvgnRR9kL79Ji3sRQ8yWFkKI5pbH33V3HPomqL3EiIjK8IkAGXS+76cUL+h+Xa
KBbPpVS4Bc1Cqc37rmre3GXka7rRXwlroDainTooXHAu3MXYXBsd9GWXEtxHHjZX
zqAxwmxYKEfiLeVuhH0Kaxl6NUG+bMXXyJHEMA+oPwyjo4/nm830W57c/tHPnbht
FSqcyiK1bfD7mhvZ1C37bVftqBmSc+8a8lZUbfGsKdFAyv0gNAdDAgYiuBgp+trc
6Df7z+/Vro+Gnm2cDmSTt1Ad5EypgCvQChrVcqov+OK+hxsrkeiO/+DdEINtQ1pi
SSU/eQLgjojpSE0Icj1XwtdBCoTXJkmL6Zlqr9i3l0p/G/+/+FIeMk/jTS5Ifmc/
XFiHPOsEK62GWEVc6uW6CCxLn0iJG6wt2XZE+5Cvmd2V3Lm/f6uP3O3cnr0oW/SR
spPTjSn87hYCaif7EOCRkuL3C+Z8yaPNdCswqr9y8w83by4B8tgJM8Kx/8KZa0d2
S/rSyovbHu9Zg+ZS5D+lxGoqKBlTxRSbDwve31RaZyeHXdsZMPedzMYv3JCgdsRY
TzXWViasMIPgWkGWJz0MtgqlASQyAmeEdkTR2nNdl14plD6S+mg5gZoFXrI+W7hL
PJhLktV6jEO0wk7DJywKCBuWNkTZmnRxFoKsk3dE9nnj+Jm7PWZLuktWmC27jwQD
hVKi8+qNEkZV/fGKQg3kim2cN+7HN6WYO551B5hZ9vlbzg8HmNjSgSiAse0HrQVx
HY48ghCqO3j3QSs7vZB7BVvlhgA+/RNC98nSkwi2yQ6A6j3YhQl0Nk3iZVNKmlB5
bto9kaO+Z1AYbJOoDvgrddoLHc4b7ulBzyJAIdnBvclyO1Es66J3pdNfXKNW/DeI
bU7tdQwCSXtuZWD+2EBPNajLaevjHdSNaWVvVGkGsir0N4oQeb/CecGVLoch69ZQ
5xIl8x5UvRSjHYwUuZTRSvE/L2dhgjN38Hs5QJPVVgei6y7p9bXaI0bH2VM4De1C
+5JLB8AGkkrUdGoeIBu+lTUTvt+/GoDHZkkEB6FIbo1AZWc2csxdHJmxcy+s2ib+
0Bb+cUpyb1Z0qNkmwSZ5DDjbrdcdGblObc2eltyC489Sb/VrrfVapBRD6kT567U6
gPWr6V9ajkJFTR13k2zExGx8R1w8zXcX8l8rzYqlk009tFLsBQqJnmaJp0wL/33j
/wDuJI3WO5q8WEzJD6Wbtohd8c5p80ZJtAb4OOli+PhSJTD8SMDV5mBrZP8U99My
tBKH94IHQkhQ9EPr9fHgthtiJIM4AuP+ufo6oUkGtRuXpAc8J9Rjxbsspx7IcUhq
4HpsG8rzy4Jnmh3O7MrxXGKbI4PzQYErDsGv4yM/5MsB/6lfP3dNFAImfS2ljptM
RUBEq9xyZUc+uZykctQ2mJOfUT7uFR5AVOoA3JSIQP4zYUCKyDGK6q4mjuU/4z5w
EkL6UjZJSsrxtqQYjvrO677eEp5iKYq455M6kipgRdmALI8aHki1IL7Ykl5h7GkP
fqxjbG5OtDREAIKMaJU1D1N9iS88H8Q152N6Nir5OjdWVXiZMJ6IUMnIxTRhuBZ7
yi9z+J6p1Cgb2lzuHUgYYTnIJAAewN2s8Gj8Ah9Ke+JDH3ioRr38OQeooPq3aJNN
/2E8i9FyYjHqEe2Djv1ofjm+Q5pNJ4OHGJjO4gTnQnfjAuDFhxI49oePUJHaRuB3
FSfl8KAOY3U1dNHIUkltVgrb+Fx024HTi4knozWHI3qv4dUroeu5Atam2Yt176NR
19cBO0R7iIkBV0+mGcAjcWbZBivux3hCBLAYVN1aE/bVr8smaNtt8bSVrTqqDqQQ
056FGdCqdnaWFKXcoFp506Yz7XSmnRFdszB2eti+gvzdITHnyub+kiUIR9hi/iBs
JX2SWT6W0UdKmPC42X0KjvBmfMD4m/3vGHHShBdGQ9sytJOZpIaWyP1kEbVOmsdN
TTXlVzKf+krE2vLSYZMCZcPEDu46B+TA5T2+5cDJycM5n8e0Vl8I7bA6u4qy5oIT
upeVgkux8ql3f3VpE/J6oKIdkcCGy8H+1GMFk+gaQX14p+ZEF3CvpXWx2Gw6E7Nx
2iO+IROeUCsM6IW++k4+Wi5N6acKzwRsGYsjFTxkQwxUr1FnQakzSlxyr6cKaDwK
Xe5xha/we7dQ8v0rVTj4yJvzLMioLa2d2zSxnc493mNCtwtEEO8iLW1HGSSoH0TE
coOyhnDebN0IWiCcWiF8103cpEZ76zAn4vXCFfcieCaN4PYrEkVbM00gQA7cwhjC
L2ZrZJfb0pNbZAE3HaDlo3T7o7hOyyCq74ff6rWpWv35NqFxfqHHovMXvpa/Ix4g
tAasSShNp22kwUQv1Z7evRt3mb2EWxHYUy0+5HSlWGBPxlUc9Vmh1yCCVltqJwpI
VKvWm4WLC4ieOlbIFHpbiXBOrZToKtRblCXMrQauJSCv6X4iGjE17LVMsxojlLSe
p9lOTNksSutV0P3oLwUNLsD3d9nF6epueyfXGeba131CtzV/4sq06mHhDF34c7nM
cxOiP2Aqb4+uHrJZmDpyayQ6Wdsedthq0pJdab9wtOja51S9dNLPNSRkNt7+Z9np
n8VuZ8jMZLiOL1E3bK3CXoqkxYmjNE6xdK3bXPhzjuQISTRdxl9qLedYEuqeLjO8
ocqvvWh4HO7YAY1UUCjo3sMLGhV4DNWQ7w1EJuPUCHKi0ig+c9KkJajmDyPVoUBi
oQiay1AOJ4Hi7Ovh2Xwbh28ccxw7w4JfsOJOCCfAFSzR0xw7FpoFExKHs4mnRzBZ
CSd9GNqqQhsYfYWTtqQ97Ogv46ebr7R/VW+HtTKmNjWZYf+DyzLZqK40isXu5Z9c
rNGpsnFxFHbyMpWDvxmH+CDj7SHCgGbgjI2T3X9NXdm7B5lHfVhKuTeRDm8AB2pR
80jRhJYHEBCiiYCwLkDoWe/AHM2XSIYZXc60Z/t+yc9pnEi1/eHP2GmWGXOh18OZ
zt7BzqFsPbyXIjrr2CMIHBqHf+0dulEuyp+GLk1JkPgVatbisaPCICNI3AzHkjSp
yZImXqnIzivcm+8ptljAxk5+VvctlsQEuRTndpQ3XeZtGBZL3tfUBFAt0xLlbqBl
xJc1JF1n2qzliiY0G7j2gbfOWo6ktOqtVr0Qn/8l2n3+oRD+OVU4vZr0YPjlOh+d
4zfIYBzQD381p73Yt2vxGpWF9zQx33Nr6asl4RfNb/pghsv20uy3YfRsQIaGpkh2
aWqbWhqyxgU16+GrX5/oxfEOZSKnxI8VeUEA8XIXxbA3IK4jdBAzTYpGBQ30nblO
8ZocXIzxK85OkPhKGE0bXQrRE5pavEGbf2lLtm9ygFLRoue9yMAQpIgkT/5l3Bl+
3EeNG26ogZiSeSJP6xT4JazsJxnPIm2B8m8BNlEfgn8paZtEL6tbuDIkblXbUS1Z
ptvd8boa+mpiydhyNvbP5ruI4ytEJi9ptqvn+9TxETV363KI/SdW23N2XEsfaZQo
e9HoQqc8VvVBr3vluGyvqasAEZ6oOga4lilne1QuqcfHcEKOSjH/ZZuPgrsvLaAU
R9EbdWbSlby+P8M57QIIWep4hN1EA8VdlOvRrcnWiJNWDAGaIASWgzx08rlZuU1G
AfubxJO4Y95BXYW/VNFjVP12lb4w5aeeZO/1UiBjK59D8lR5b5TmwYHpppFtbqGU
7YtTSmuoYlMXkKHSg2eux4OblDtsHztLichiNp4co7Dr8KUZaIWEZqNM1/D2BveH
Q7O6oADKF3Y5Z0gExoumK41OoD1MVHLH8Oi1KAm/cOVK3AQrGDPXcOHJFT1WKijy
14CbPyf9idJcVx7yD9KTV7F9Ie+GbT/vBKmXTVVg0fXnu2ix10MKrOOwv2OxXf4f
HktitOyE6QokTt80ySy/gBFXLEooZ930CRzElVR2NC39iABBrlG6csZF5/MAxt/c
dWOg4WVufB0gkYsfjAyCCd5q31Sqj5HuajzHJ8m/TWG3Ec9bPFU+YmXsv4rxdIDf
1p6xVt/dyfPIigREQhqRXkLgCvUS941kJWKv6zk5oNdXSPE9GVKocLnC5ozj2tSx
KmiMgrSzKi6PEX/92zIZBhv/9Dcjf3tNr8BKvdlQ9d3eYghvVrXHA2H0ruCUZsCN
2sjSvrw9rnn8pjvv1VYdEybRdQRVl9hzgykwitsGQsn4XbG2yX2+07XSfCcnTu48
TH5n0dV/68vwhu5FEGvl+CMEjdzwu9+96cbxOQfF95mgYPPkIxxstxFKuk1HJ4cX
ryrzrhefmoPHtRWDnoewnDCrLxaLWlw7etjPpU2xb/u1MOe8Ixmib9pw9kn4c6em
pJX3P9O7sW0dLguJO16mCQVyUTA1+J9ETv4YbJxOp/3IMA+vdEOdz9QiuujuEkhE
TjDq1MpDYHOhBgD61CTKFwKh+HlZ2ELBTWkPEUjX3bwcVG0OazHhU03iS+K8giDv
bFFoGnmZ9ynUsK5tgJn5IjtieRPVEpstQwow4yvH71b5Eif7EmmY5WeYo2Wim+O/
WVUqqirnheYomu7gATlsUboXkNUq3UzSSru7bQk09eSTalNGloPAGk0u9q8kB1Fs
2vnq2eHoKiupVNTykaE5SGCjWq0WnrgNCHsfBE/B6XYxWGw4c+iiz3dNuvM2eKTo
DljwmJ7qCdbovtHtQj4uEdTGUPdZwASM1/u6Jj14YD42ycNxC3Q6TbQRnL6vfvIl
y/Fc6AY7iBbjbqnLpWG2OSN0nQA03b1wMVGBrQF89WlAxdf9aQEeOrwOos4V4Tiw
5XLC9+CPEajW2HidnsOTo4KBjlNvY3oiSvwkCmVQNT7vK3uPjz7G9Cglzey9JGxv
qcdqjhQbEmJJM6LLLEPRaiUnJNp28sC8t+qEnzle8d2zFG+RFVD8xdu22L1HLnX+
StlFIpAt9G+MV6lRkCKZBkMY3GZAyrMoWN0rhebVpiTQcsbAfSktWXYEN87xRcCM
eZkG3t7SIC2P1FhJ/DMYl6eOkVSIJlaiwjgmfE2FgsC7EoJHkpjhYIOcMKodi+uZ
dxVeiddg53DJPVpdqZZwt29pqYSZotaCLr5VszhgtDGKkV1vfjyM8gmP/Soy29gf
B7D+VkHKP7ovu4XvdV0VUwHRCFIkfq57F9JIEJUOHpF9Etf0HP8SROuihoBGrWI1
+qzt/Yf8X78meIpZihmXt9XI241w+ISN1rnckYQzo4NgAnqkGE2Qa19naG/oRIgL
BFWdFXfFZ5V9NQUNy9W0qG2dhqLl51bP2zwN+gLO7XFoKhauhj0f94I55bSm3DnN
L9darwvow68phSv3qvg74lcJB8zeFiZYip1eYmS361XeWNcnpT4PFu95hUMeiw5/
d6eZvEq2SWzA6iCxF9l0gFm2VE+8FPJRI6j3f4FZotUgOMoIkJ4/KXgAz9NZqlnS
8j7YPaZq/95BS/3KjSfbj+4Zscwdr8bhXwLRNBHIL6yCP4aTbq4jNS1EWWJi4LGW
Jtwx5m5q0V5awlBi5ZKcv5IEJWt2bjl1k6wqeujohzPeepSZI2Qw7DucicQMhdCX
MmrRXV18JLT93gnSyQ+553qJYu6t6VyrR2mqexnk9m20OLB4EHq04o+MsJEfPWIb
D93muI6wXo1vpZ6p3NpLvWu4uYTB9FowWSLaaQPcr05/1SnK2KcLJMtWq5BUXdPx
b+OZmcqFjC2VcXLUjhTZ60lJzHaGcopKeqU9r+L11guq4ay5xJl6gl2iHx7PvocQ
oH30u+dCt5jEGHa9pGPJIbYL3zdMhV2TKMHHAqamBfs939/mp0150OD2rF4hsU7T
xckWqxhlEtjC5sPWpPuQQL45GOYFX6yJwA1WT1XtIUTnbca+ZNQJfKORCx2l8BH9
KPTMhAsj+5hrcQg3S72RgVQsXc9AH8WnFOkkJ1a0RlLfppe4tN94H4EEdnClbzGQ
0seKh1wSEI5ImCtw08GRqZsANeD+OThIHC44nMohvU3JC0W/8vurqLF3yzqTWnNh
2IlFTlvT99isbegLuPDrFe8PGjWikquo1e+ln2N8iGUIjoXHPyoyQfUbU8Y2rwSx
+0YCmyYTKvnoBn2+H7B4bosjVDifqfnV0WXf8Gdfzozq0r7DN4dNebHakZn53OqP
cQOQCmfohrs4MOp6pWqabAakrE5Lcojhia/5DP2z24rYE7i4Et+SYkywTmPhEpMT
8OrLERuP0/d4BfxYoXFnflyb6mBABnPfL2wGegknXTX5e9J0mI9u3v59COlKnAIW
oRq3RB+oJmMxvj1RfSe+dLlHj/Oh0O7UZXTHW+n78nxPbbDi7agjlbNWrQoutBrO
aywRpOoxx6nY2iZK6feVKEiYFWSj+TvFzkMC8c3DHvckm6f9GTklsgMTm5+SFrH5
3dD8zOdF9Iw8a6B6oOwD+1pViHbFAwTqimeDyEV6w55/qmyNF34DdU0aAQ7HuTSB
lb9fYxGCEb6dOsJEZIGO3C2Vt4zgXhmJQqN9Vmg1odPyMTrqz3/q+d9niYoxAHy6
i8N3hpzgHnJ82eeRBEtiID1y4LsABmj4W24VMwAYSiM4JjU+/aK2POMyp0xie2/T
SJlmHkUJ3gSvGhzrzA8M2QgStWrdMDiSPri9/jrSD0zHAjOu/mlmUNCa4d5BDR3N
zFzcxrb0j3ACzOE/UId7vTVK1xxgQy6MVBVoosZ/H3//7VmjVrI/fR3y++kojBOQ
3MENzdbMpZspbtGlJ89F2NZz9A3niX8BCBwahLxs2pmCPFiQmkXGwD25yohATDdK
8QK07+BnNAVw9+3m+Gg8pQT3G2dLrHON857X0uyLiFUEO40XnM8JiLJ9YbYLpOIv
UaUq6antM5T98hM352EjZUSERdBmZF8hnEbwpNqabuhXWGIc4W4yv3z3kxSQ9WKX
cwLmSiUrYS8fG3HqaEmZ/3dvx2xDUcltfQC6PYgE5FgV1znQTy9n3cbuoaAM3LZX
Xw8M6e+10Fd7DjfHpuTF5jtb7VH0OIVgO7yLeC2ch/YkuP42OuM5pCoa4DinIRQm
pnKLbtMJmPTF5+hnCN+B/FDq9USzXHNmzTMNuwD2y+ph6M2cQeKeOSF8FQoeyVcj
ABXYh/O7CfBlK6biWGX95ceuFkIvKcDI6WG08QeDhGWA30ruRy3VFcfaBw8rnV+9
j1Gkf3nByEmK1qU7Og1UNwdAr9k/Np1FTPZNNoBMzIl8KAfBKP7Sz3a2vqF0iJGJ
vOxgxuPB84jn8WK+mM5GCeHT762IHpb5UAZYla77K3qPOszKWeF20+cvqLiHSNKl
eCxtvdCoHN7svKDOkdnVlFDJKMACPGl6ZHeCwYfMvRkz5QHNczYXlgUO3e4vfZhO
8C+KVJLsUImmuz+CbFdYscw3CRG4+74+JE1NsbajK0NxzdOTdJ2woo4TKNEYU6s6
9nOb67im71/YLwxynS5taINTna+Pd6vtxFpNOTgrnXakAAkWBHAYd/1rGJaJmfTa
2NroZVNGz8PawwrsPDr99Z/xwZz/BgsjOp97mdMBUtKiOZow4drOD2PEa6bn+iZw
eQZ//ymwRyXIiLGNA22E0AwVxI90UKUGZAz1zmlbL3MLYr/+hdn8ZD/btbY9GgY0
Rqy+++y7//K+7IZH0zwA3I1Hfd+fRrkdd7lRrmvOQp6u8JglwF2QyNjdi5Usbgv0
GRgANbft22fSKuETXuSBp64MYNlAyb/1ig/Fm7rSEvRn3S/MfLyvdiOe5RZIq/Ll
NkJzqGjbvgikaoipjiNmo8RhZTkaw7xEoFPSFPlXO3Nz93hI2VyP5YTFf36shYG8
DWkJn0Nm2d2hxBpMBrHcfOEqrRJO/xDEiObEXYV36z0BIrG01P3Ue/IdmuamBSc+
Fsu99fSqFBtYXDUv+mLWfnFcRlfPUleaFBR9ZF3hbTPTvvny986KL54ojmhlr7D0
SMQarpT1ldVSGNRx/2IBEY3Gat14qsf87Fkz7pgY8MZdjfpiaOP0ZcUAoSZ+0Xsu
AgNM61eptt0A7IPgetZ2Y04qpAB2m7q2t6fKZZ1paqYPuaNwIA55oyMUsu+ZDNsF
/W7PESbHfzhuD8CcX0z2yMIvnZEtbZFiTt3/oqGGZeuim9aiPqdytlP8KcMKOg9H
WQxAQ8MdBurTl0iUpmJvtc6ROjjvrVKoDe+H5I2KAjdu0eY5yDOFlHYKLFk03vmA
Wj6oF0tiHX+aMWo6Kua015t8pfjdtXqR796G6or0B3RseWqWQQREaF88wADG4Rk3
WA16ooEMjZUX7LFBuboI8XgBlxJwXM3je/ggjZjJpfp0ppvpC1W20olE1bWbyVxh
Lw0FfihkFH74UI26DcoDKFE1NqUDMh7Zdb1mbHNCej5dxev9aDmQ4O8PojP+xAMQ
c7EBqL1IGbaE/r9pcZ1lnndPTMGl0U6mwiCytjfP9JVnWMDp61MOOMc0SZNls0VO
kVz/OC0YSPa4z4krld4IuFtAa2WAZjYSmY9Vc8N3v7msb9xSwtLXd7acpEFC6UXH
b4pymArpjFvAd69bl/2FlactupGcp3j536SjiKUEVQrLWyF+jseC7BjF7uvTA86W
zKJUJzy4in/Y6Q1mZCQQNOta8/N1yBjEdaYIZEpOqqoydcB7O1dJN2FIZW5zA+2H
flb/9IUMXhIInquAendmDWoWbw2ELK9itDt2TomJxcyMAB6JUOAxVj4slZi1zZqA
dJ7ayIpz2pOhyW9Pxyd/c/KF7hpiJIxA0O2bP3l5toPXSrYsRfOquGiVuqc+qaQh
8uuWnDTaddaK/xDAWuUpzLQYa+OtQrf2VQAD18H17naSUttGs+s8q2KdgLogiZeg
FlsXhIqFZGhRAb6duWvquTT/kekNg6T/NI7I5PjX9FPyIWzp22DPEub/Jj16eXl0
WLn5g1Ht8Q7q/AJ/8YDv94DPpMa0wotq56NiL6LJ0/9SVpfj2djBwr8pYc5iWU5A
efNuH8oC2Kh68XXAiPxYREwQqWkedPLxXxcuKx0uG/SjTUE0m3ZFJNVHe3Xt91Gy
A6QC67PXB0Vf7mkc438EyCfK2Uc9rX85kV8or4JxtCCeo5thunwuUCwTtilPQxH5
f3IF79Ux4d488rfXz3oJ8GFrEyW1BzgoDxOW8fogtg19zjiEf4nbKrwuoWGUMZsn
ChSdCS4loJLo3jHgGo5ulwRv9kS0AL5A+xxzeyFuMjVqZ/t6/8EVMep40QIkP6/3
fCPCesH6TewfXK6ZWDiNNYZdlbiu4YBqUdIhY5Rr09TXrCiI7G2XMRQwDXlhrFXA
WY0rHdiBAKQthTSlYHY8vRZ1RZOArI6EZlELK4IBmispt+mbxh1BYgb6GW9WizeT
uTmFQ25TKNcYlDZ2Y1sacrwdypP1hkUX33q9zNHGp3XCbaIwBipsbZlld7ft2zC7
CPDGimBYFgGpWQufyf5O/DTHedp8MOdjlI5J/VsXri17CtBbjuHzbTlbRX0pDaQ7
rHNol1vIhr92OCzJwBaLyNb1tTFbhLRRv1z5E9cFdWlyXuKVmCloAzPyxOLQVhMu
wapR/3j8Ilw5rNHyErgH8KVRXYRxAUwr7MQ11kaBhlIBP9WrS99cTPnMd88au1HS
ielZj4MROgxwtIN1yvM+QYQT/teV7s67ImuMwfg5BkvFWuQ3mtE1Zq96lbDTXoU3
P9WlO3AizIGlZhY/rGigRMtaozSZnvEk1y1bAq46tGjEJCqJ/vevLC+HK8tQ0Yw7
T/Tcoa10fAX7FFqfdFPQRo4E+XRlFMbbG1NbMwGK8VTbQ4J0uNVNFP3L+ndrv8Ge
xxF9HcUHHhjpu6M8F27F3FPl7rDo9YpemTZIZ7PQNpiBs/01/6YWvw2v8IUIKV1Z
4ZYs6vaO2BVZfkXBYOSRXdzZCY21WtcV32caGkYBEmnBZMkYuwYN/JulqlcPitvY
Op7yDhrprzc98TKW4dmW0+sg/4aRewwBtkvrhIgdEdeUQwm8kBwz0OzuUIftjUqn
C1vUlWNoR76rbguOOiaSQ4JkCTO2DibF1QM0l4EpdAYbgT9yBWAvwPxpY6zxIA9N
pgG66x9TIIEeEUo8p72ZIqp9SYgPRlPKENb5xM5x6Zid4UuACcKu5x1Q2pnS4Evj
KvIvmHnUQ7vMZCNHYYjCQZemh1UdawC2/BoM+qIMxnSz0ue/hOLLz3k8J1hWp92C
/xbtm7oqohgZ1ZnhxYjBOhTFVkXTuCsvwNbWp8Six8/WeDORYOSZ+7RPLVySrGN5
fc5yEm65o1yMscLx3ffUcKbGyQbyTK1VpuPYiME5lN4qdkH9t4oLWi91cK9iAHJe
KCG1mFQHuZPauQ3TCau3Ugg5ndL9w1/G3j877MB4WSEju7ZVPZix6hL0uCxGOhOx
3w6UfhpyMCTcEeAZS3zDwLeX9Jods04JRATfnHdRlX1MoSvqLPglbrZTHULh2M0C
Bf3qDNrbRL9R+eE1tX7grC2ETuelGc8Kojaad/qPAiUSzHeom87q09zMH78lnHFB
yZmVtg+4A/k2+xPIbDl4kol6moIG5Lu1tU91dmLPRiU9giPdub0r47aFHzq+8Boi
EAM5RefOrtwZ9JdAUSuQBbYRFkL+uGSTtOz3BWdzq/jBubD/mGFa8p3jziQu3NNR
DCMgbt4R00cGfHuTOeBLX/qnNzuRjzrHFkH0IIVdRW3lbUadQvvspMpgePuzMGpW
gCAgeDb9usmAgdJ6rxYthvGiHGtd2AEuumj/shhgdxHSHdC+6IAGsxzQx5jCFEiM
TabvoyO37Hh1tJjUob0up+sP4htjr2v5BqEpM1Nqy0qBG/i36h2n/5lfDjRtr6NN
5GeJAwErBZK+osGKrPRHn+hJjuO6UNRB5FF/FSewXki6oiTmJ5TfHYMuzbM8FTIu
MDNF7rLW3CwNM0FlVwHkiab9GemUpYUKrtO0MAfTMmbJCjjulIgplt4Cs7DoUsYX
1lwANETXkmmh9V2EYa/xm1w+L3XIXo5ZHiOB3vVLkFTptHVSwOqR+kzjtpLyZi/q
Lj24oekofUw5pvIGXddwW2Oc8zOpwPgWK0GgVN4WUI0ixbvafJ73RDBeVgIwVDLb
HEvM/GeX5cfrmP2yjPfmFFpon7Hextkn2BLFmcxXvnq55KERer3BMJDOspVtOKSI
gY1VJ1wh8Pl39HwKrhYYpfsLOHFr/AKnJInyRCxZ/bTyEnpxS1cAN419LT9teDNH
RM//0KSEXgXBHrNvYp68Q0R+zMSQdYXp94c4qDp6xQSj4rjrJzCPxodER5p+hvSB
qzYdwwZYF56DdOJq2AOSpZVLSFECTTIoJx836eAZNqed8VeBJ9Qp40ZiEyccHhgc
Fhwa1+Vmc5aLIZRddaOhubP2dg/8Ot/Y2N5krXxyfVCX2yVkSIT4oCrmfzc+KpkC
33oRP2u6AWYU9D0Yhq6dBqwSYqWIbsCK/+EsB00TSv/44SjgQE44yWbGGOLY4Wbq
rAcMlDk0QVQFAsB1tKJgYbRX2nq07y3NALvK2isi/NxpLCZ5y0vlkQTtPNqu5Swq
FagVXi6ZVDdoK+QiqBX0IKORwkJbbIzmxgz74ajlP/BhXTUDT5m8JfIaIJaJv4K1
Y8iEmWR7McLUyXGy5O/RpS+njbCaJI/jOIXS9V1TPU3kEaKSNZwcAaMTr8ez4chq
Ok5I7TfXrG4u3o4sf8J6Fa4digBfeoWroj1cax9v/vEdKpQG+HbE5IvhnLK8A7jZ
frbX/5b8rPKzQ7e9wM0Xf7ERL1JTDU4A6ajqVju67bbAiH4sHrB3P0slnfg2Gkub
+Axv/vV6lMbxj01ud0jub3ahWhzrJUnUCvmVRNug9iLoEZEFZ2+4HrfJd7ATS9ZX
itbMQs0gnT/bDoj2YqiySNqU7z5IJkCEtc8wDbZL6DvSNSoYJL/8yzJFeGjfUj/S
F0fmpUO4HKUfv96h28JnVPYT6MZaT9Yavq6Bw8OnBxi6qS0fYJd5N2rQzg1sZc1z
bp/18005RrK/bNrm5fKwf11NjMFRk6kDQPn8zuEeFfBpQw7ybNJwb5bI4xlM/tVJ
IRff+hltswv9o2EjCL9BobB3o66jmrknNjO1fIlemedmtd05ktGlBatbJdgsi/4i
garWN/kpZOCYEUp+myyjILywNL6RkZkXzvkofCjhV/wbTKJP9iHagGiV4NWjC9z5
pM80rL4pvyaFnkPItZznWSqtFqDf3KJPUoPHVHnutwPl/JlnwqdDTdh3GSmu+eXg
/aG3AsrCFogZHCYpiMZl2uos0e7TyIWCUhfYbavGFEhApvGNGWXKHVANf+UEx4sk
a2orZ9R/KngYOcrQNEJaQE/EUPzNduxNAlhFexGCwPcjLJQQDw1oLBAIS1p9T3vg
VnVnAKSTA/O6i5pumcoxeHVGTXk8aiaLvr8nbVqrbfG1YT6bxhFrZMhknsJ8AvcZ
g0bVjkGD8gdMdyUmZXL8Q3PlScO/is1I6BlxMM0J8rB8RgQKkIsQ8XbzkMXfoUd6
i1JV9hgRU/uaeq97gfG+UdG4FuHV7jPU7nezx1DNlFDMN77xaazbxoDzCVhf0R5y
8DrTnKgwKitIFIq+9gyNaL9/7YLOLKRtH366R4zvZShBU3Uj/+nlBRPmskK2fX+b
c83ayRu2YYzTyVnuX5kWBkPCorc+4Sqa9LghcLpUGTi3bbhb8qGFdtdnq5HZlTTp
d2mz5qxRWGbs8L0tPFjcwu3F31ddSWY+JkW1flp5PPFvwSxzCLoWltHlIZqm1HNK
Vrgd42tWAY744zY8bvZQv2oBGqKMImoMyKJS+OiOmNVckwbhbQWSuHTFTR7WXFe/
erH6pOzZnGnEpoUDsuw2stRHtsiB8VAFia8eS8oTZNbv/Ly18QZ29wQe507VPA5r
I+tee42DgSepaNUleCkTVqnucpvPXZslLeyAsiiFiPA2/h8ovL4MVcDgD8Z9cFi8
854T62rTHe0+UH27x5xpJFqgqgRcR2VpAsBq3vg1BVYXeNRvGHcRgCIp1eH0+285
GyNUMI2YvyN1xnsHs3WXnQKTKuL9cXRHk8jCbeb9WYNTpP/aAbE85vg/Q5kUsKwt
zk9mqhz2RA6dIMxe7cPcH7KEBK6GfZzwuukz75roC4vvznllUSnPKckDaD5DNWCk
YP+PlXOndL+ArmuNR3BnSLbc28REn2QMqd4L8kG6Pn99rbUIdRZynwjoCzwOsDKE
QWOUC4anM1GTZLVokf0GS/6HuTDjqiTGV2GkdDYVHBN03ixQZlPaSXFAtGrX8Mlb
AARxWO8P9czIYaIq5hPn//BTtTbjJmo9nta6V3Ovwu3jVw7pOieD7tfZ9chO5ppv
9iRQQk1dN0LmDqeRoOBovkY+L6CR+xYIv14+bZ47mrI5G4MDRMYDAtabxBCp+W3a
9h1eJkZfpyhhT3ivgZXX9P9O6uLGc10pPIk0dctdN+EHgfxWOSlVP0owF8RhWZ7O
7H4dKpGOYts9F64w4mss79N0Mqd8tb0WRgvGLTywFb5Qa1MPDmCrFx/ywJKeVAI6
N2fv5S+NZdnE3myfj6yIItuQb6T1zuSXf3E9BLjNiqBQnrl7WHQNMOzZG4sU0TbE
TKRKhxbdHZFJRzVh18pN7OZMJR+U6J7i82cHkDr99Wf2U9kXg9DT+scv9hLdmpFa
fHxMiErmQ5vgKUsBBqqJqHn2HfyL1P0pSZ8yeKXnlWcCGJS7bXCF0+su6SS09P3r
vXNolIhPaMe++g5NEKHzIvaR511UwGHGl5iQvVtecI5sUNv8ke65OhC1IhN2FPcc
a7fAqVYjrBuNhHJjvotf16CM1L8f64v2A/JWYxdArAghUxHHg+w4P2N0qhJMxzHV
7k6R2TdAKH/s2WC+wclbIc9GLzfQ1Gj1VaYv62mSRKltBCCwjsCLHtUgCJCYxyrX
cCL5IP2yoqYqlVxExjTl31RfrL5wdc5yecJXu3CznOMEVUrlquZD6MVpZPyONsGo
mVvLsSwzGcArX+weRPTgTIzFJuW39e0np6rFji8Us9ebALXMq9dx3QAH/axxy+QT
KezWWjViRS1STksKzWh7uhNeARNKvlqeoZ206f/zEzv1OSHphJKB62eVOLHfaBj9
5sijbyTZamk7LsTxTScx4MYkdc9eBef34vrZ5E2/w9v40IzWgn+70Jj8fT5ddYUl
0GX7WoGrpOWup/xLyB3eTJ/akockK4yK/cxbynemAKEh/TazlBp3DWZNA/HWEUbb
mOU6pJu3mKiOKkyozYdoxRxy8FY6bNUAM6rUQjFjXoxixJUy2IN+jR/amtMNIa/F
C8Fcts5XGdACi5L9IltmbyWnru8mnNCrxOTTmiTbhfVlPbHG6Gz20JGDPHlhd7iO
6cUQ0pMCjj1D2kBVpULpfW0aTgvgnfp2Hykp28WGh/mK/XvWeJNUyLXFN+eubC2F
sm+ZXEcBUfHzNnAWpCqaWUOPOhGeZq29Czl7xqp+O7UFb5FHcYXb8iC6+kLmdQ9u
531/VN1vweLg8B0ITJ70a7QntlZexgwn2t96zSsU/7NbQmiGejI7U914TpW3WniP
D/akuMeUU/Indngjc9QjpSD34PXjmWO535sO/RUQEbYd4jF1tSl+K4TlMhJvvsJs
6qfG99dkqQ4Oq/zwUCf4nOYVrbmqHsyQqnGUJlHF6RaCoBRU/u6edGf4Ya7XhbMG
vDAh9Ewdou9//qAFDgDyEHW/I2GnqPElf7p29ktqCh1+DCK8bzkg5nH8pW14xF6A
xGEJ0rvRT03trZVrCxvYwqHGaW4v8xQlwStESOfApRejW+TuPQlq1OOdCGZnt0OE
IJ0KFNrw7RR1D4til/jEZMtQZL9sme+6znj8UCjdRrQZNGPtiJFTeGNXLklXpdzN
OKX0s9AR5HdxtbFPnGQAtOzkS+if1Vc8gRQ1f35KNWPNcoqqt+WGCZQpXd51TIwS
to6H6E+K91425+HQz8CFytd7OLvLnI965rZ8yXdQkaXUusO0X86YpgZhH163ik2u
6WfcW/5ksNHp/Xo0HPkv8V0ob7+8KJo+UL9fqLdAxEvogahCRMdgZlFiL2GK/1UD
zEMDvgEAgTqQF1IphwsqTLQkkRRHFJ5IWqHhJ77+yDrW4XC9JiTpQDHt1jKDcK0L
obIlQ3MAp5W6JNRqgD8vtH6OcgOOPBx+nch7s5nNKz5xymQGMnqrfFm2aj2YSuNf
pU7N1X4+LLWsvCq8sbbxb6oFy329g2zzizZ2JNJSf1f/9n4wmtefG1l3rkrQP1ZK
YZD7HhcpmaC8LsRIOEmyP4usfKAjujsKqIXQOoUe4YpQ5D+k7ko3rmSi8PmlFyfJ
dGqbmRtJ61tPYI93r2mGfzmKBdkBaxXGTs4x2L2k+417asB/7C9oRqjEycFMTlOR
mCaJAZVwretUMkCTYmTrMjbeRYhw4/P9ZMHWbBSpwvHsqejqk7SF35bHIId6CsiN
GweUI+J+9PQZE+hwAbMA5FXokhK7roG4vq7dV8/l+LcRVkr0wgC8fpFpEVFfwViU
GQcaQHpk8A5T56cX+Tl/MRpVn/AOsh/MgdPqc9ps9LdcpQGDMK1aFpLYOpzddz/c
dC9JWuXD3oAO0ZzKCAWvkONQakRaSKq01y6syPCCn/47vAKUncjDfMn0bHLFsv2v
Dhp2n6fXvQcD5dnogvytuLZgl0Vc+V9JGvFMrr3/GZ/8ubBHHJOLbqMns2ZW+xdH
VQ3OfPtRIW2lrmXM++75Mc1/H8tXHkZCR3apDhdmOrfbneSUfHT00S+j8DKM1/wd
Z/Mql+sqFW1eL1lvPXUjLL9E1RLj1IeT8YiMXr3DZRExVSzvmtlgJCWMhWgfzlKR
bGErElkVz2yn+vKedWZ/UV6VSjNeS/7OMylfxcQZwbjQXxPwhLLRuVTkvJm6ycik
P5riND32pnBM6ZO+pAlEMSkAPP3pIsrHf+Xi8S2qDew8S3kqfGCe5SplvZ/ZFm97
Zsu4yW50AmCXlDPdGPTClUiSynp67ywI+zae4dDJbgCeVKa8rELYmMBXXtxCG97j
1QW4+jyMyzcsYZ13HLfMGM6pAyP9NXZ4GOR+w/AOPsi5Vs1gzx+KRc2UFrQNYTIh
rVe6FE3C5VbZgNKEPLvDVnFwRZ/3yjyAtGNjJL9UTeRPAGMDxgvhbWFgBZRNG4ZM
J0v3QiCgd8bmr9w47wP5RzwwY5+LQywpk9T4ZmDcMRpUUllxcqkXvxFNbEmjD0qz
ORIn3NBu/eBOHrnfgPVzNb6PjqeKKach/HQ562dy3FV4HK9p6A97IVClkNQJ4m+z
rCIYQTYRZZwa0TYHhaWH+21abG+PzS2M4lcqTeInhvHvlkdA0uk5Rdhp9Ft+NGOg
awnbob0iOStW8iZkHIaZHkkhWMRrn1wtR2rJo0JnBKZuO3RB2uycU1D7SWtpFHjZ
GpLY/kEomOKpG8+ROcHFVk9IerWvFKA57IdTf8Gd4j9xihmD5NGg0mvX59GeJ/tB
YWkSpTca7XW6moXEjrIFBcsIsMxRzTFvVeRUvvJUGhCbXRuDpko1t5ekCXmgRJYo
F7c3nVHICG30i7aqcgqFxgds8uTyQbx24YL6RgqXGGa+Ozqq96zxtTQAPWShhnMv
6VSRhXXTvAS5HXxyYL9p6SezIWxNJCaKuv4skKOE+R8ZSeRe7R898XoOHXve72I8
uUMaYuiLy1xcA1LbLdlZi41l5q3exKIef6U3TK5v1nodyxyquhFs/WAHEGy9Vbui
EAi7dopqciW37rqGf/EJ2dCv2G321dtdyooAvVDrRfxf+Ysm+mMLWGmJMWf6ao5e
/JblrlwH2t/GgJyUFf+xekfDh5NwZ2Nw/86waDy5WCQvOPfD6bKUdTc2aH1VyVz8
dydPfn1jV69/YZA4X13WvT4BXX07hXoGivfkqb6splmATmM4zrW23fIu3CMabZr3
1KzsSumv53IAs9imugFNmVExsZ6dVBkEX+pEVApp2pjMoH0PdMbIT74caF/6deto
a+31uPhtszIPZIqohqwBC23cLrrJoe0kcPGwhWXSEN91FIvyAyL2BSLNTWUJj9kc
9G4HR5y9Z6dsdOmm6lJnxaoDmXnekLNLmRjQAUyHTUEQf7DOELZuJWmsP+USUMna
diDIZl5fd7xSW3pUZlkgSCjBwLMJWM6SBpAXGNZdMJxfO6IRadzbLNICZQc4R3El
cXgwngwF9UncU8RpdJJv3oPn/VIYu9IUczUmwtEVEUqau2p7ImxVveWmkn3KUU2t
S1fhwFLGhvCQCM5H/115StXitCqWnw4Ok1e6jgbyaZa4+an4lu3bKbtthupRr7qQ
XdVzYqS6Q7GBkAze0Ru9n5+osT5EYpp4+IP1eCrHfXpWkBebMQeHOi4uSOBYPSoM
cDMVrDdttHlg2AF2nY7E3u+huZZSbl5jX5UPOVQkpFxpWhaV5t0owlusEFxSPd9p
D0myfPP0YZ8XoZUunJp8yQj88Pq9yKpxYGEUqw6862dHw8RijSwVIl7XdJDt7eht
YV2K0pNpqh6PogcaVYt6bB/Vm4ouFTyxVJ2pPtqVZ1ekvBbxzd/RyHazfefee5Mj
w/ugMCb37CRTk3LfJdPI3gXfOH1Dj0lcgdjY8kQD1rJh+CSzQPL35aOb8zBLGaJB
CJGlhlQhA2lne/FacS5R/hGtpq0xRVQx/ZrnNVwta7HGnwj8zWGOF5S501cJ9Dzu
YelJ0U0K8ssYsIi3bJsvInd+XvoaeJUBReIPT4RHbE6hf545q+c01oMcG/+Y8z+U
7K5o/heEoi9s4HmZv3vNkHJKSQJtBqR+IzMBnKwW8qh7kJVjYQNtPijFHqCc8maK
zChcg+vOdtvlPyf8sQgWssR3PSH/SyLQfbMylVIekEGpbLo/KQbfGfcY1foUL+/g
oL3cnroK79CBm06OFIxM9PyohMKbiedW+t55lORVBwPPOZ8WjU3fC/5M/mNX0t8K
3Y6PmTeTPenIKFW0+T3HCd1f7NVfkX/I4OM+XUVKt0kHP2l8aF2prHnOQvqowhDC
W5ZZWHCMqop3xIa58gjjZ6THslgtUK7ptcNMAtGNxJRArI6tzuU4jjrnpuk7qqdm
aVCSQyc0LVhUza9NZkGJrKRNMF+lGDWLVPbuPmbwhR8GQsWrzLJCmZIK+kbRl/16
+EIpZZdSPRHljk3LvxVD0licjl26A9V0DWuFkhKHVuztH6g/C5gtAUl+8qh9A0h5
87O+7vBt75Gbe2awOe+yKBLOkFKEurvn0HGr54X+BZoSJdLoCq7aLGsbI8Rhyf2+
jHcruyLG2oNhYcQI1ZHYAQmGUOejLI+EQxHuPqCN0Wr5ai102ZPrRIUgd1xq3yHb
u+ohqvyq3q948w8QFTjoQs1UyclSLOV6re/l7taObOijV6k78Dt3zJ3Wihz808VR
C6cg8tPLvXutU2UXiBqZ7O0QGKyysiyViLK9bm9le3+/2mW/vjJc33b3XZgbhihI
uxzSqfAdxxRqT+cwqYanIsqLPfQ18dGWxMUw+0lCs5OTo0EPVovOVBvOzuOcH8Qu
dkBfRmdflrNEs+sP2Wa/ABmHhUfKll5xM/DxayKqLs/mEZO4Uu5iQLn6hM4+535f
dFQdWgvA7I2gopHMl0aoNgtcM7Bb+iuSlEbPv/oMGIzDd/8XYClrH/OKDX1GJWgB
5DVLeqZH5nhia6sN/7lmAQG8nTX4LQW98D62YRmFHGGloFBh/gErwB2+ZZzBENvz
fPErDdi2lfW1eyBn7m5tFt+22A+bP42WuogyZ4UxGpZj6NoTXxALAx0AsM7WdOML
rTvS2k26QsOQUd+4w5J5hoMfdCxXE47fM9VO5HYv6UYTwvvWgDU/+x69jWY/HHEb
7WGhO/RuF+gjhfZRQfq6rRHy6UmxKbftX+ujAnwDCYEqhg5ZFyvggERsxmg2v8Ui
8ZlkpOU+65Kq2Q2ZP/ozf7Jn9rPtOHJ8B7c+jKUnlPrSOIiLpRAKhRaYund2/B8W
ivND+N46AFavo2CKmarKmd0UskAxG+TvVs8tGC/v6qxbomPZU8QrGJL7fwn0osXn
4QNQcBCh5iaPvnMy87Ny43ybrJBX9UQC6f25gtUZYw9nXtWAbTyMMb/zNRdPCa+0
v28zP7y7IpVumrxH+8LoocDYxCy0Cq+9iez62vCTUZedyeigAbCaGb9hjpmY+1G6
Pwej57tyCmeTeOFDy7+60b8wqqOqppx+qX0qur2aY6hcmSxIf5oHHY5RgfICwgtY
GevkaD2cRo2x0wQsZlAqgqH2meClwOTGwI/h1FxzvorhGw3YihP3L0aYCEZdSlAy
EVLIv7JmtSVjiB5JrnrEBbg5/4I92aWz/5ZYyaQkosoPCfIgQKZtm0KWA3/Hv0df
B/tp6ruG2w5nTMmddsY+xU40nAnOMF89wfgJzHtwIH5u92XLJIcugmEjiXkhj0Qv
HNnyawhAHqzmCjf7OZGp5vFlFvKgbCmFz6yqPTa31QNLqrXvoyTMsrblumuyAUTG
RcCCIrhL0r1v9snaJtx9XnqqlWchHUGL5uJt5K46pRYt8gJDU76eMXctaqQG7a6f
f5sE33N6lb4HPfuU8PJez4K8WCWc6lsx3DXQtbBpC0/d+ceEEI9GjfnxjUswgTmu
aoqkLpdMftr3CzuvngcwkyPefnJULeup8FpQluFOOIpQJCi71Oc1zE6qRCik4u8a
+SMejuHhwbRyamjmtkXFKAlLn6F6ombvSeDRJaU0XwwpNciU56MXDnsYPYpwS7LM
agtOeO/r+RadiOW5PKMdR3MI15jUQNIGYqh+aa05fudethQqv1yHNrOqJgiPqt2X
YEsGV7jE4ZV/JjX9tfLpKtJ8nRKa5LQFLo0+vWLiXSA9u3rgdhFreAe3rIb1EnCG
O+3nwjiVZCJb/MhxCeA6uQDbmnrj6Aagth1rQtI3JWEydApMgttHYK7ja5MfzKLT
P/YNLZuTM9fGfwk6yd8jIpm8hIpKsV6pYQ0nOWPYP62e4jKEe7o4FA03QiFUSoS/
m/PLzsCd3NphkGcaVNPhOAh/H5jjy7f8BswI+iuoeX7Oq+I4zbkpJ8O5ItEB018q
6iGJCmZTT3BVjvmhZ78BMhUt98T7KuIy9WnnY/KRHVZUYjyxdjxoyjJICyb+rTgy
ZFVKbvrSphu9UZsYrdXwi8DA4Z0SH7u3dNwEMA6sdzaNilnRwroE/JhORC9GXin3
eEw8JFko/KNL6kUzjMPDzdoID/5sQoADtvFGNzYQBsiE4bEU2wQPbr9SuEc94m17
Kdmn2yAY5/c82e1fMOw0M04yZTV7AuWrrrh2ZVnv1H6GqmakwzWTI1fCc/5dkl2X
25cJ6QfKAsDnCMEb8Wwf4xCHKAhU3TJRAgzXV8hRaLWzN3RM62euIWXwXTREOoRd
6quvhpMenODh4roSNNekEWxXR0H/i7jWTskFE24ErNrGIOUNS1DQXVnXpOE0arJ0
YweeEaaBaZqUg3aSpthR+ZzuIkAzIVt6yGej1s1nsZqsvQao++AG6g9XrEqAvMdP
gX9AyQ1b1pup6nBUixx6KcqYQp9C2JTc93XRrIDdXgm8fJkWaIbLG9RJbVLOqLk+
kPqjjeH+lCzDNrQcAxoDZZ/khdMIk4TKMtLYja7ef6iX4nx8XcT5jHSDD8Y6Qbx3
wV9XU29VHJ4FnskYyvk6SScLJLg7sgAlEkATj2U+Q+i1zwJxvKKwk4xg4s3W/9Y6
wD4nIChMslAGF7OC1hZPL6LR+WoUwRSdAT2jY4R68CT9GeA9z+YkfWoPPUnq/OkP
9SrO/6WILrJ/aJe7iFKVj+1Y93h8Gzu5/m044n1CqkT/DuRhwzVjXfvvdOb0hwkN
oyvo5uMyEhkYWHIRCSbWq1r03MNetX2XueTlyjylIZ1kw08CoJM1FOxp4oYH81Me
wHRoH7r9TQ1ivNB1nZMbnO722hQKj//AV3d4iuFym6I+/eqehpoVZQTZy7fw+ZbV
VXSzcT8tnttqvwLzEbC1+Ev2pdoQWSDIf7ZdVVUxxhYW2AW0gM9cTk03nogCgifJ
S7jFfA26Ei9HMxYtfEczkWIDHHb2hAl0FaM1TmZQWlmpgSlgQ8y7l8qHHa3fcN/W
1PX66aGkZvXUN/suaQ3HFK/BFya8Gv9et/yqTi9QjX2mQ5+EDR7rSIX3gztO82el
D+F7RpeAvuFsVSXMftzTt7xxW4E+NUkRiWl9mZQDoHjjOLw4t0e4D1+exOzdhi8v
kdOvgy8wfEPC4l7ztxnf21wYFWlFELRF+nkTCSue8OH9z3jxKPcw6glfs9bPU/y2
+CajJ2xBTMPoX7aOO7Xx3/ptCc+G87B7ouHFoQvLRQ3JIA/TLXp4anSQn45OUAeg
vP4M+phD1CnhUto4iMu10ERHE+2WUY0kCAHAO8y5BXTMVuZEMV453Day4bfHmOzg
`pragma protect end_protected
