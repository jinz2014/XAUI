// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YD5Jy4Tsys89tnvE8+9j6P7lZw8sms8lEPESpHqbxTZc+rCHbxx3nJ7+5mnTk7GE
GQAvdzGUvOlwANdc9rb7nbFKPWUQlGel5hiZm1AHWK/4NnDENnNEksxZuct9gHmZ
JQiVDZmgTQUzslDKKzeqCun8FL2Nku+8sXaxEXOVE9M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8688)
qBSDtMR3ZiFcC5nQL0CTiMOeou5mmWDZKYquLGg/vs7sXHAKmAZDHFUfHw/zmdQr
9gaTtWldSoYQTPcYN33n+eg+vOUhjAUOyJuNv+yXBmUEVC367tPJyl3neP+J4ED7
OEkA4rJyuamOPsG0inSc/XXROvl7zRxK0lFd8oU3T9o7ljKA0Seua+uF4ELkMw/h
B4AYqu4VY2SkxqCotNf46A9HiqvxWyKIBap64Rrzt7bCBgkcL8/oNtmDVX78gfw/
BTd+DWpcFhId+cVD4ib1nWiRX3qoMcV9AOaGTcea0h+a4jZ9pnrt6FdRHRcb8Vsu
m51Ldqyo827ol+Ks4VDxi0o8ZueyC1S6DnSb7h0jqRCPFsLMKkI+yOroJ0jHRMzY
Kr1dqQxdBBE6t7bfN5zvJg99T2MYfmnRS8saJ7E4FNwxOjgCsm35QtxdLQXcOJFr
XKKX//jSjo4oYt2bIP7yTKCuXTTYvK7d7EtFLn4zpnalVS7fK9VBwfmqlZ2BDK+o
Or1CfADNs0pVytmir5zTt1b9qIcKBKuJXQnUmgnaFmOwAfOHlzfoj0BhDBIQgnG/
o0LYXCzbpGWT5bI7OuNOI1WmGJZbO9aFTzZeiTA/VEIS9hPr0wqJwIa9Jtsq92Ac
4nIyBnrG+V5sOILjwMLBFK2g3LeYl6loZIUjOU08aVGhWXD5P9h+CVky+wRNODcr
bU6iplHsPH9pQd84qPvsJntSLuie6R+r7nfOdmLeUysshLF/I7idOw2p00ZrFu78
AKoCrrNXlHYI9MLGeelRuhnsIm9UuBcyuvlZeOuhrpeo2zRz5FUGnk/pMVQHd4ZB
7exDQ9+uR2NiQP8PBsVElxsM2GwWEYo6c5B3+BTSsrAr6aU4ZZ7UftHDHOxciJYY
p72VW3dlFr+C/xdQoVVF54elz3syXOXCTw0qLXuHbjgEICctLK7K7qqXffM1ks+7
pvB61oiPNK/QtHlUt9LkliKhzfCIWS7FzWDNYyr43w5AWqw17A6gxt0GOe8xvo3X
0PhbC1AO6+tvXkKrEeGHYcyN5xRSvEE4eSoBz8hl2NZ+kUYd9qurT2MeJsrillhr
stGRt+1w/31GO49vaM3tgPNj9wgqF27LnzVK3U9G763hfG5gyuTH0/DPTE3pU5vf
QW8sRpnldZe4GSIBcFapErfGw9MMjkiXeTVNmlksVbVRmR8oSE/8ApJ3T8UJULtO
DSk2kOKHldBP1kAq+m9TP4+S0IsTxEB876NX6heImyNh6121O6PpOAiunJQ00xsu
m5q8FvPw7V1ZR0eq+3dwsSmomXoyhZ2dRNfgQqZNNFssSMN6LnWDFx751U5/NjBI
jyJS3263stfgwWj6lr5PCQxMTqLjmuSu+DX0yF/nsRwEPrpKWPGbQDs32B9ty7ZM
8CRjCSNuw4GlgDzGNc7qyh4ZFS16AEoyTZPRv4X1PSK9VjmbvEHMpYzL6fyDL3qz
fH4iUf0FI+3ltBzDufQiru81UK6mXIPvQaf5kkWofgRXDHFOQ6K9cvGI7yXCHxob
eUSDiKd8D+Fk/RDDCTgbdXkeee2knEyLmYbjfeGOXfCko5zdzpXXJuLgCosoGVGn
fD9GxtPbw4QX84JuOuLCS2d5NKRxOqcrFBQBzt4jN2LgqIFDYQcShsx+JvwnS8dm
AOxC3C+jGRh9MfWoETUW1J5XuAl4Cg+UegDET+Vex44MzIgD2ZnUxmu7MPIz7Vc9
DrKZ2reQwdn9nCdMA4/PNzXJl+1pIL678znCY2/9xQJzuLudKUX+YYcoqR6NBzbO
U69JOjQ8edtWnHTzWNzmj/Sh7h+7hc7+R5Q3R77uxHSk63IXNGkejBMEi7LfORAe
FwgMPnTsVOoC15z8wpbY78TbDnnYXTrs1lOTJR+J/9z5PwSAz1gmViGgiMfUKO8b
18wNsKFWKcUfhuVKF9NdTUhoZvz/4EGWUmPblYJVEL9wxfSJ0RIpbWH+hecvzKM1
O8kLP0Ofuh37PG69fdklnub8UOGi7MVBXSqBVtKoPsDOKUB+OSF611HBt5Jhujxu
VLsTjHl1XImualN0N86xI3pUcVxnkYSCawVYIqa6J/B5MT9NJpvR+55zh1YjVNra
RApXpishPvPxZFS0CLWhMI7oME5h8QQI7rhBTEn+TDrgQQY85PCpIlLcEM5cc2Rt
P/AMp1mb7xca5UOksRHrKYntSdaTipIxeqaZ7wPOb6z20GVFSg3/yI7xldps9W3l
QURDlmEPctrqiNvDvKWPd/eS9s972fYQaSciwtNk8yJcFMKZWI5JuM62XpYEUV/7
micvpAcB6Vy60G5l87YpKhqgygoGwTlY0lbWBeIeiaIcXVu02nDvT+tbE8D6cNWD
il4dRB3/69pfCRmiwPrp+Lzd5bsX1vvKy6TWqcmLeTRd1gkNUexhh9gFtwkRMqFG
BrKovGSZL696kN3wemCv0FLWJA3Bvw4B7UB7zus9DtebcsHgn9sisRvGBibmRSbH
zak8OsK15iiGJf1u+e9OKCe0tDelY/CJ6J8/ajhDBjTxrDRsnOzjp6O/YrMnU/v1
GNWvDj9EhmWLGAaPrHOTJgHtS+BYLLr/h77ZXyBo+g/AX907vB27nAA0brA8zWIS
8tOUoFesnnnYYEdhkULh3jZboSQMYRGXwzxh2le4kRJUjHvRctZGnOp+3zDNjEIO
Em+5207QJ25hTtcdE1BbUeE0iWApqeg9Fcw3ZfDv2dl97VEzIj3xf0XpZp6v8oDe
BsY7j1UNdYondJAh4R4bw4WhjI83cQZobDrKLZSxl7yayaw3hLc3NkYU5uzEmoT3
kP4+b2UFdZKe0N25U/ynF+Y9ZqIOw7dRZTNLS6lfxYLFCWYLRNK+8CCR126j02Y6
qBHWZUW81aT3xH1Fg6tpJ13iclgfdw0WnPEi6GpAfLeutydVNTcpX+E50COB+Dti
I8SVkf9YQ0nZpAvtKybZ/t6tVlxN6aG+ZlaU6PvbmyiOMGDsqua4Tge8Tm9PWgUK
4vhj2zV/ohuULATy0JyiemAYeiLruEVaVibc/9HtYI0sgup46z+nBzYOHAFMaJdQ
1K/JfLAYIsszX3gjAT5Vx36oye7XP6QXvPF1VOTbw3xGDNt45XOgPK/fv6kwrlxI
ir2T2HcpiC1HOEQMSw8ktIYLJxKxzW3ePY59z2L2pAngltNSs9QgEhxOY1aLOoPW
7WAXlZSegtiIpjqQP0yckKdOuu/oVFGy23wDOgqH37eUpeODZZ5NX/92MeLOo9cD
zGzM9QWn5UJBnZxuFiesH7GlX8PO0AzK5/nbBZhPIGZNmQ0VMtRz7TqY4AHVnIUX
lIHfCF2zycATQ047+3LILkIOZKVBGC8IbPMxgeoSidnU0y8sKuT36b0E9z6IB3eu
LFsegMLcL7AzHCf1BSSQ8NdMcA3WhZ6/xvxYv+id89/SrI73uqyD3UUSgz2lTaD6
xo9tsC7fr8lNuUv8tc/z/6VBaYLVZZJwQ4AWOOqp2O0zfFLFZqULEvS06I2XBs/8
EUWa+1RC8EzNBeu9OBP7+x8V+QwI3R8Uf5cwnwT4j1KxmtN1/NBhkRQ1WB47LQZQ
qf972kYOriD95Z5jx6+9tKdR/8xAoCOpP8Wjak5VnouMOpogZy5NCqZ0tLye+Wph
LpjU3ApIIiaGDVjRYhCBsSD6RSym5J7oYhbzCC9tK2ldHctdGop2d/EfcnhCMbk1
BW43m5kLdqy7HE1tSMb0tSAVnI+Q7Yu1z3yWTpkY29baknrGMeIEgAJSOt/gMK47
NsorqSxg6EDah+gDRhrtSfhsrfEkKT8LxHfNedv3PRXbQlxSRxrjMrnsqDTgoZ32
CpP3awghMGhUJCEDBElv/Dm5yKcLsMxmyHscPYwuHpuA3YxCASfH0YuhzhVt0x5r
KNAWtlFjdAqLVGc1NRHrU/ORGBmZmzlfIQzbeZLusXU4QzFk31O+1u0kkKkK9GWe
EbfGd26GUdaJLfT+2YtmcejJMYKTrKhPfg2E77IPmF6SHElaJVjQNg4wBYpaPNDJ
Wd/4IJ9y8CspGmxD38t8hvO1CbUsO+UeJesk1zVgGqAK18yo3SvM/WlZr+u9tyVi
kVbYdlpoqE9wTFN8/KA3pSjoKRS3VmfK99LclVziAb71nI62K65WXo/46vOxjMLw
RXPypfDhjIJCi4+XJFd0CyIs0Lp5QgfC9nGcjSMq4g8WEO+43Qy8kCyMHfcJY/Kp
HMnIhXcQGmQSyBpZMWs++COUmyZRr1CYr1TW1DagZX5vyL1he3VuPVO4fSCMImU6
35VYaCODBiXnt+8DFy+s0rPQkN1Pp3ba2crLd48hNJuDZmPhhqh9xWeklfJVWYUt
y5LtjRsuvaZ3gvGXcIi4RhFFA0U8aDlFpaGvlIPp54TyN7rtH5vdWpiUmjSa2Lwa
4rRlfLA8+2NNmKIN6ERdhT/PMF9VR57YY96Vrw9ilhbCB9mk1lj9AHiOw2Qj0vFe
dDZCc9S9cAfdM5rnD0KJX63KSvyYD+zHHsaReSnHdNH+Jekz0MvZdKl8orDOFB5T
wceKF4d0Fo8KLpOV7LPVkryERtL4srL7V300LYnU+htHnVh5dZl4lw9v6OGWyQom
HmLGLRthFgDEyyHzIXzTazGxnJP2/LAmGS03hy/88rPFeLuY4Z/Pif9eCJFaX8Tj
MauZ+kp+mnF5bb2x4pmwwwYmg6YuJGAyUQHYw5bxnhEF0mkrYl53q+DK8lCc+kZ2
phdIyNy2BomXwzw89ydMkD38d89X6WNPiqkSGrhjoQ4L55Nep+EGigrhoLzwXC07
bDBtADf5Cs7wCg8A8DDvRlNar8xq107ddK7JAbETSp01uSXzHSlfmrq8iRt5za/U
BGAXe4sFrUF5I9IvoDYIkzKErENAJBV45ILK/gTM/riTqqK8ltXS02UX1QsFC3wj
QmvlKrgPXYQLSpKAMrC6E3EWnDBgPy3wUSPzwt/RziOibnw0C8CTcPCM7813wn2p
GLCoeChdC4bjMHY5IooKrupHPsEGnxE42PA1DL2ugh6sE6kJOUHW7UNPABLVuWec
uCttAZA17WJq+14yI4cDL1Fpg2HZdEAdeIhMkzf9kg8JmLjELLyY0QRSa2RTHFoe
DbnZit20NQD3or7bTqEMnsMMdSDivQT6bS1T7EaBMf1e+P2OykXTbPgtipqi3Z4P
PELbmhK44LEYCBzLSN/dK/ioEvYOgOLwi12RJnmKi/J6G4Ow37RwvXveohgnDJE2
lydEcfFcMLZSHsp2Cz7m2X5sjNFQfpPvjAcZLN1bL8xf3dte/vNm/ZWU9lrET9tN
UE2KDJMvol8AHsBSAGSA1SezE7FsrsFTfjwHNb8EiRtazyBjQ1jzLvM9PK/qBiZ5
0e0da43a6D4NUCnf1hKh8mMqsEmUot9v+TIzFtft5CprytsVzNsX8oNTgXLlycJI
BkWnpAR8MCTbGOR7KZI6k9aiCoKhL82ldYPMKAfCAL/QhjiRD/3pmB0LP3UDh2Ux
sKnFStWIVkjpON6+Mm3SxFUXfXgL8uUyTWoDWwr0ukPcutVeZLwW/pvRiHdKf6lV
cx2QktxaqTdjXet1Id0YQzrKpJU00fL7AI4+Ku8VPNVDw5uWXMvkrSeo/gRkEMX/
Y2t0DQQaH4xQq7/oeGuYrEo9zWM1biqdM9bjicfWqnyyaCuFNpl+PNq8vMzjX2IA
9jMWiyfcEesq2imhAVbUeoIF9OfDWP8VIewR1Nayi+mA+Bi1/iUxR0bVXo2LAvLH
Pvbe4qMJLq+Il+9Iue0+6/SHZMMvnYArcCUp4ehiyYJ8ik+YWbddnLSSL5aXUtz4
4FobSMyR54NrWBurBIuVBwmkxOy9T9XoKHVABjuoXh6NOS6O4Hkx0G+/0GLsxL1C
iSMG5A9OJRJ+hN9eI2AKMpFxcytojAD9VhI/rtM9pYfmZJh8Af4vy8YaP/4zzjG4
8vz4OVcCylweN3k56I41HAc3Gq7Wc45dmXUAMROm6A/7hOll8IyahyhxTL3vhPot
5MBtHtUa1BsxiLWevj1xqLb65rTuRi4IbTl8vpHY7g0IcGatVbn4eHSVd1QEM5KQ
lC+SRt3dBvvlVfTqdWYz/X1H5IqZu6DE//bjEK+4DaLZG33eqGZl14q5NAPqU6Sl
0kr79TffuUPiZFn4SPg4tq+e/sBkETuAoN9tT6OjPjSoiIhXe1U3j1JdMSM1KpyL
aHfqyc/VD1p1igmS9shTAyM2l3VU5IwUnSvxVuYWM2UPK1t238UGYikj15gwV2aF
iEhe1NLK0ZQHURu0/J2bQlqRARli83VHu6FbG4A02y2BQ9Qh0nJXiPPSHgZxLlal
XF0Ig9Z91RhU3ZPUG5own3wV3hiUV2sMq1opFH0UcVKaZ58RzxASDVwsydS3U4k/
hgtbOkA5T32Jmc/tyB5KWawlcYx0sh6Uxw7wi5ARenwxv9GfjKJdc/gfBbEA3FVB
2q+3LA2C72qXkJRicZKPOdu7VAuSeAe41tAbW3UY6pYY2hS4q/Fh83rPhOcXGeL/
PpTjgSUzQaqmAYg4AXDy1lPFlGrD5zban/dDonDnp5oVf2kRKeHtadOxMG0Suvd+
n/xrfMgdtfxtjSmbd5hnuBLfPyaIWH9ptAxdul57WBTgY/fPU9gkjkKkpwNlErPS
FbaGu4IRMkUOeapmVK9CSLK0ItWNBXo99QU9r+ikswz15CbQpZpTMIfjVzUDyPWe
Cw2FBt7Rb1FVh8gGjGqaEo890Tix6NY/3PU485vXL1A4zIpIIT2vt0+4Qu9fAUsO
WxzsXxi15ZwajwPwhNDfnK6dT90jTn8cMvKtyYNghzXWVW+1s/1ZhjTyduUmhus3
ksRd5Gt9XRPxc6F1QT0de2EBs0otflDfJoqrL29ykTyxtg30327zNbvY73D9pGas
mAyvWEGy5a6X1Dzl0/ihD73Y4pwYK18v2/cyq7P74O+tO5YDC76pCL1t6n6Pd/0t
Od/ascpuWwJAX/Ou2kRvZs+IPUDYE++HAZpNssaTKFjaDxcjuV09d+h072Uhcw1I
epIS02U6I2wKrA4kubWEhsyaPp3DhGjV4nJG75FoCGcHxMzlJfeHuEJjp/iAPAlC
K4GOtZ+aPM6we3BMKyH+zjR5yY8R4PzBuvIyaBZo+dC1uIVR/0S5AZWhYY/WqxAi
VophdRYHHP7N4beSHdpP7DwzmZzRDcos/dAGvGYhdIQiQZ95EVVb+yTJ0QzrlfWd
oyvMfZbHPagZE2C/ZIzABUElRO/oIf47BrxlGWJziwDM8Rr7KOSn8dmnWOcCHGBg
yqacx6PcVxGYplr41gAhEhn3qASRfe1J1Q4JK8kOnPHfaMqExF+O671SIoLTiAUG
l+1b84rqBYhVJMh9opaEBRUsBY+1G9izEpzT06UNTKsnVQDDbSUKX6vzt60bczDt
w/H4MQ6x60Na0Wmj4TasUELvY0D7t60aOp1w91wc+/3MRZuPjsWT+aYQ9Kdw2oKw
fIha6vq1f6E2V532YycGC593ZV4goNUdcQ/pl91DeXmXHcfSnTkDYXJUTCjqAKaf
P74DsTroceapHwQ5nZdNASSg5sMfeq85SSxtTW/fpZO7U9fEYjzkYOaHZl/pYRSB
XS8c26gFJPH/dm7BvIJyRKxv3Fi3TCwRnJLXU1+fBF3lsZzFJaewpnBDupyuHL3+
EE9IlDBuZAu6xOHDDGbnks5QC3s4OzAh8v0mHOKuKzZRWmt3q3BIY+ya0NNG6Yww
YBhgGMVyyiB8zLF9YReOig7MrocqX28PNjdFBm4wgR55Y/jn6JqFD/sOyrWKiVYF
GlFV8teYur9ob1rv5stsOzk+mCkGrQE3IYCFR5zmOTRF86gyhHaSTH6K42c3Pvsf
lITPh9FSfE5a1IvFPVfjjCjHG0qn0Coo1fxGIaizN73Hj3bxR6Eh8mPKdoIMZSP2
0/BacnvZYs/ogAgiLl0xDB7I9RkM9hgWntyyQhxYUnVY1IUQtvcCe1ZKKP+BWtDZ
AXljrmdxuT2EMlWV8EdLs8JDNHTfyKRPGYzSggHxVlIc+eOGl6quWRHcXXD55ZwC
jvQ/DS7Dck3ahXzb8qo90qpdTo5QmZDqEmhOeWNYaamjsmrHo+Y4J3KGN5enbNHc
+0cwyzzzecuEJ2YeY5kxXw9Y8VdXNJz7RcH4gEMzDdMX7iTiCp1/E2UFQmxQF19W
DiQfj4jOtDvNzKCFEw4ImTzNfCbIV36Si07KgWCb3TsRcWhzATMZb0+fdbVzEoQ2
pQoQBcCoNGOhAc7ue6JHLKgZp+KMzjT4HXze91sSI3/+O2rlWh8wJPbQ0YSrodM9
AOeyq8lw3Pvu9/6g9qsnNCLVLm0f5mG1lOjiotNdCxYd83wv7ubYQ+1QXzdQrxoE
jTcYP8MGs7KfwTxSrRE93Hm7awOpg7kmdzpCN/Cw8ayCGZj7Fn/PFJbogbm1qUIO
2bqBzdGq0BL+1NR2kC+7qNbjxt7opbchD+3uaWpVFDbwM4nzH886BBiXwIYmFfPf
nl443GjT7/EJ6duVOEyBLSZzU5qQobaGdWYpkaj8jWTwh76kCtkv++bGDQiYyd2S
35NPL+bXTzKCftdzXjvQWJESFemKv35QVPqF39wIiVikfdkShVnWaVWnCWeQAXDo
A6vyd9/t8D79KtI++/+YQ3l6V1jX+OHKRbRmLw0+XF7FD35wp0bQUpiP1CI1Koew
zJVTdx49CfbMhKZFsHIKtdX7pZETQH61/uSy82l+K5xRs+tcTFz25efmDziKa8hc
iO5unW53IbVHSOyxS+0uHj6VR1E3ojwmxi+sQG5do803qAR6y1bhW2j2OoZbZ4wb
+vlTE6rywU11Br5SwX2kfMu9LmKMDVmGKSb0HfYhF8AYLyTS36tl4j8bNIk7W+2w
pG8omBu7BNBCNJQb9NUeQqMa5GoH/+t1lA+d0NK7VieQJEvt/OduMEg/due+4f9i
403Yuon03FD3QjtvMuwln0BTvzOrMcBVBFWr58szLdrnySGqZfOcflRPbJTGprgs
dBxD14pwR9SsTpgu5Akvhkk21Z477VLdzEzr+loO88uUuE46XeHumn71sA5hC8jD
oWwx73YxTunvn5Oxy6RZk8pbIp9lJTGx0b2LL8vNlPYnjqpckskKg4k4jV0eORXt
YGqPF2V+DMVuvFgJ+cySdado8Bbb9AA94jLtSlG60BSAqiAxpI5w1w+sTzXId5hJ
Le608uBUjvQDJfsq+9y3cPtFMvX1NpbSIZrasK0AtX95Rab5LecDUnbbMZT0WcZy
UMKDxumn9RsfhtENsQ2Agsv53LOeqRSnlRC7kYbFd3Tg2z4Ht4tOObGncccJ3lc3
lbnT7OYftj+uyQO4CUNrZo4Yhlw7yuGGNUpj3/Ej1KXNmJ4OjLgkKdt9hWCdiSeP
NBmWcadFjZn98QkXxAq3j0LHnRXITGUkeMvxXEfm7lKRGlHm8ok/DvKnKhmNEA2j
0BjxRz3/+i+aPlpGWRSHQLgq22vawxhG9anIkgCajCabIEjgk7jbLcpIsC2U0P9J
UmO4JKz5MO7ZWn7JuUrrZLUJaV2lUTyCssUDaYN0KCi3/7LBXcg+I4vJwVDFEgjU
VtopxmQIixtaTTBr6k1rYkf5BSxxMC+G5stynABPCW8BLrTIz0ucYmqVBk4XPgXC
Mck5Z1rHuGmfcP9LfuQ2jC1i9UEIrwBEA2NStN4J0yQfaDFwDVCn3Fu2L4P7bO0B
E6uWc11OLdGMUNOSYJjtOfy6ucwRJCeBYK+L20DD7mmgcZdUrkZ7+7uo9J5T16sP
Yfp29YG56++QDhu6S8N34fDOQQm9plWoyXqxpJNOKP5w+7ZWrfTfJ3CCazo5X28e
QCX4kwyFxA+6Qo2Gqi2KtQHeTY3CgY25XpeI6PoekLV2EWx7rNtJinudEtyTva/3
yBipeD8YmBJExmuOiRQ1vjbOCFZCFmsDXS7MF+37jPrDLhdZA0/byP9oKH9N0zcG
K1aHDL+fW+J0+2TC8XcTefILMOw25h3OYCiy5VVYeDcNqjhC0ne6X2dnYRvdGt9j
FYCbUjaRqgVg1HI3xxJGRjKLsotwKePV+FtuQkN8ROUG6uei/M2a92pAnZjXl7B8
H6izrMKUcfT3vRjTEelEfMgCLDTCFleGNn0RptC+LV7WN8D5g83XG+APvkIT6+iV
vXiJsEag80Yu7SmYdCX7gwCcPasr7jogEe4VrryS7AHOgPQdOrDPozWGXsBuu7IW
54ehL90rhL1qSZECCst55p9z52tbUBfvZhvoWlV5E1CSqsSWPU5F81l3c4i2PC4c
pKkGQQndjWf1EfFE7VxJta5JfkZaQNtWCyQ67h7tkf5cZ2egfIyfPeciahARbQVM
U2eE4u4azaSd7Q150ZlWqTtP97l25kNKicXX/642CTrAlrISC0VYz01qCgXfc0bp
k/qTOrOPN1TSMS9h0cbL7hV3mwfRWs26soWs3+vWAtGjf7Vn0nYsn20rOoUElwCO
/BUGYhflhqcBB0DEpv/lWIdYBKAm/DGt5uKoFfGsoSbXGVNOK00n5b1haCEioJYr
ewCq0PuNFiPZhBK9yl+W9xM3ZKT0mzgZ6FZETtZeBk30+hamb82AxNC6LFKlycD0
Nq2xmoUVVjnkx0syIEG/2S/zgKxlj6P6YTPTG+Dzxbv5L63wxqfYBMGWLx40cvhr
8w0vESQujBTzyIAUSxEVrdt5md5+G/VdZlOb290EsW4WiDgpG1juwaCipcweec5I
HpfbcvlzrKNUOnL5+sbHyG5B9rCZC9Ob/ujRznqrPbFQPhbW+Yz0uY6fAPAEY78t
GrUngVqNSlYJNMbCFqy9fV6uGyIoSxYOumt3wRAI+fZ0nvXvpCKs6qzqwIUphNK0
ROCi0pM4CpARhwHdhIummyIVz4W0VmTawIgVhR72FVYTbSad4ftFZp2z9rTp6y8M
WCwwKMxdTQKRf3jPjbsDx+6ROdDjHgUoWL2DCFcpBvPwKv4pBDUsiuqs/4XQfrdT
oxLmtZnMqyNdgZaYAnOubCVLwjDNZ5STcVNY3BMdKPotXjcf9MIhFeRxTo+jHIae
Q5yiqiEQxzXWjnnV8QLtSl53TqFx9FHMVOUYWSEY7IsANkDQ1PeD3uhEocBOj6i4
gPpi1hu/o4qgUZn16Zd4vMEhuu8faciNg3PX8eNlYa3sn0luv93XT/YAtAU3Ydnj
AeCWPSZFAB8tRdu9jk+HJr4K3QwKuu5G54PMoeMuE5aSnpUvM8lAA+gGphXi1izV
/3EG/ynoMOtPM1x82/O+rBCekEU0Q/y8EYD+lxr/1Qx25ObIzCRp1n9d14mREYh3
6mBZuL3fst7ZazDtnWtuvMj0k1a5JZ+9g3gAhOcIw2HsDXROU183R/MjHXfGZV4x
urjoPQsSxd9/Iw37XUAcP0CYha3hPE8fOxiGYQSvqm9cFPYcCRgzQC/npr2EIooN
C9YFCVPs8Q02YP/W3mbhJ1pYZ1WwmJ1KVZFzzLKBaEh4OLYALMszFBtkuyVegD7Z
p1XILQXJKHNngc1o88RcQe4QzZ84dhraiZw/A/qS5mLNW/tw/eDfFooC8/0MbP7b
`pragma protect end_protected
