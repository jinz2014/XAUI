// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kiKnQkFS/xGgybOBkSpMIZJcDyjumOeSwaX9u/hOdSJqkNFRva2Vy7iOtpbxwymO
mFjXxpkv2k0v6wT6igi9kaHeBRNmvh1o9x+Kg86NGCKHzNOArkRi0ivw1fBMGraz
99zGhoBPutVjOEYyq3YgEpFtNGg0QI+fGUxB/Sw3krg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1536)
2i9lhS7O0ni5brOvqREScP5gxyBdL5dRn7uh6Ge2xovoPAWpOYM/rNhLjgQk0WUd
zvniAvQ+IxWKxguQgggfgzQ5rpegnoUgF7n31rc5KMpkYgT7WiiyA6LScc/Qics8
IkX6hFSlUa6+beZOEpxOKPE/cXEy0vcvYbEGcaVtxTwls8JRR0gNB4FgJnKh/1qN
5Q9EiyRXHn21RWMi4684/9dE65JA8xKO4z+USPmxVJuPElFhhvyonvaX6UD+IhGA
GUqh4sr+LSkMBcOBBFsqY1F0JAaWWr1GrqTUwEjwmbXrLdRZDK8bI9PX+0Z2PbLT
UEFlYfphDbWxBF4S3OnDiwjn58Ip9iJApiKr6l6Oq7VZggafqNI+CsvDt3Jmb1Sl
XYnmVpaLjI/VxkFgvqK5YdfJ8LgCIJQATfsni4Hg/xY5jrrxzbh9BFzBgcJeYS5M
xczuwFPC8OFs5I8bA1izc+HUzFJmTkvoACvDkpFHaEv3Z26gvK6KSUT/vvxUKKSG
XHaJvRf7w+jS48i+lk5L4U9cA25HRA9+3NPxsnnrFMG0vGp0F2kdpiz07lUGtzJO
ZIXHjAvohbpVChX8xgNfjlf6APD50s4TrKgnWsAAwU5v58pAxofFrwzxhSPM3jfD
9eBqbLXoqb2rZtcVJ2ocVufvIrlp+YrSPxEAI65uH2MKGoOzaVUIFB1AWgh1jARh
DhcLmxVbCeyAWFdD/Qtk906oG1X6G3wKvYpJZjhELUZg0CSy1NVUxFOYfIc+k3pd
xJ6kx76JVXcXausZnMVDBjn9aHE8PfnTrQUSxuY/AreeMLckDa+NPNBMnyVfqHyB
33SsQS26HRIB1uxGuVzThQq74V+OuIxKMPq4JE6EeubYjc8Yx7L1zZPdg7kU7Uc2
hRND5BWCEGIpoaMojMwlxcvQcMk5indrbObJhrPz1CHEaKKLVLR6SzPsMRFLYkL5
OnfzNtGo+bFOGwkGP5Ze4SdKpIZ60Z0WhS/nX0701KY0jr9hTVN5InGruWYnSoHt
Qyv1i+hZiAmC4o3QFYpnXmjKwvcZ+9wWZpjxs2mnXm7o5npeoYNgIWRPfvRk/xCj
uuSkUV/8VIjfAS5Wr9guUn5alCkHaOSgsQI9+mqMfOdYd4vbLsgqpsiN61oiwBBb
VmpV9W4BDB6s51x1OZ1UgqJwtrIQYkV0qyxyPRnmL0i8MtDeUtJnWW2o2NITjwKb
trekMAjFTEfBtxdfP81HmC8G+NcQItU5MrgNK8rWRDBrutC8+oUqb0af1RHQBojV
+0vZa6zsuQgBUKhRPXsIzu5lzLhJmxbCIXxptIVJ4PA0j26WFQHMQc883w7Eht6U
NCZM3xwHuStVVA0+TnPMdORAXdlppEsIkYqc2rfRnBAcNfBW3D/5qG/dhM7ft2J+
boBkaHEqus6LWewptXQQO5+QWG/nOvpW1ajnJxRHQmO6JYfzsRXiGpLuBz2l2mZ5
+wX01HWWsrW5FUeiuq7THvkErk3bOLsv/ij8dILHfdS6xUxMAUnKtquqaeEEX46w
L8wnnaEiCoqAroR7MqEvVflAKLu40uK9RUgFrVBdeBuIzeUogt3FGwjrnMU0P8hD
LPGwrUmSHy/BndITAgxusX3l0CZcroM942nalAS6zQNRCTf+aM7sDxN3MuepgiiN
t3XK0b1RAIjc4qcmbuJeit+f1OfDImqZW4gyqXJFVegohH26AEZVCKuRL8wj17Tp
Tb/PCo6jV3fzSAEgpuv38h6q8LhH75cS/QrUCh+ivfw1zJ7N2TYTXj0gz5Svpuir
YfMINDLI+XFW/D98dJQ4LdbpNg3kq4iS8U3KsiOn0uH0j2fphjU+vi3EBDal/z/6
yIwjwUcHmIEuzYWLfVdFH5sS1r6C6sMHFgNSf5GXFsOkoD0wn3pQJC8AhccUdAfX
dkTw82zFiAXqQTsUsrWJvzvelS7u4fkZ5whztihze7ztpE0/IGYklVtDokLOc05P
wyXNHclHg+h29qIcq2FLRyxuSfqxvrtaOsaiT3zS2uDS1WeJdro8lunCZ1M20iEE
`pragma protect end_protected
