// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fqFKy8HfpPihJBdJlFv+PTBpsMObmmYCmyzk6l/io7s68Zkgp0r+8Q131M/NFhz+
LNpNw08Z3DV8y1MybYy/c4KlXTGNLALkAKh6D4dE/HhdHzfvqMShMC8TfLz++hoo
NPKvzT2rK/KZOKvO9npZhKNkF6+Y17tYYqMu7IgF1Bk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7744)
iI7xjkv3sfSp/MwQ7XewFnlRl2fwmtGpujbWUoiVpNXnUlWcqnnOBbVBvVWKvEbs
hlD82FxNOAFrv13q9p93IeuhkwwEKKOS9+USqeIMSIi0/JvKGVblpbd7iHTzzN9J
zFgoN0YyJhPtzXHJQCnfjdd6tQpC2yotVubMw3/+XC2zHvZ3cZxfM75bQYCbwLbk
3Qi9thbf2IteTYFwC1t8Vn94V8He1BEf/90+Eoma9CRC3j83QnWMQKyuLecVrY35
Bhl8ZkrfLYd6NyXf9WYBq4IIlHx7UzSpQkc+ZjgnogE5wj/IeDAsMaU96ZuS3lz0
koDGeaqQtxrF9NGtWneuEACk3OrgOTFqLtWmcdeqQuc+J6YHq0o7aQ6TCy5ieYI8
KGnY1eMk2dUq+JtTFy7Zm+nWKSyAfVWpUXOBnaHir0lt0L/tXYmXy8O+AbIsJaU8
XdXaSlrbB9pCToeYwcUis9wQIktocgmJQD80/m7HDyYM8k3GWkwLRtEqqegX6PY+
fl1PkMB4vqMGfI6HpKwSIM5pSDykBNcyP5Q2WCAyVL1LaD6e+vDrGtV0j/WLmc/r
pkETxOqnXkCtaA96oQTQEnOrJulz4iPVwUY4GrDfLYDreN89ydLiACOEyOXW4QNE
oC/BaX8nY7LgxEtobWnQC0R3/9MU/hk8KWUec8W+ewLJyFD2LPOmU+aXaKDaOvWR
V20wxmypK8zVSUi9lZXgMbIQVCnNpNHvhrLndRHXECYZshdJaj1kDNx5Q5HIQ3zP
lA3YQfZFBWbWZ4V2ZLXf+pmsTqXNXvntnY22lpsx3urf+U7Dnx46KdGZeoSGnDfe
+5+0LBL6qMB2QndSDndsY2sWjGx6QJiR5dp1LTToJpH9seVHWtF4z9kQaxOvjMUF
wFu0Lu4HNFzB9Ik6ViN6VA1Hp4stiiyssRIf8LBOy4xvn7oyCYsPgCjHFpFWqWDg
w23sIp0kmOX+bJh/3hgyHtbyNlr/Uxa8gHBqUlK47zkGWuQnNPSwzUURELOof22Q
eFZwTKQahf5QlLxxVISBlPOZTgPJDIhHkciq7kQhujxP7WfKRJ5UlZNJa37cM+ED
dH88jlq6nKJx3UEgx81/hnPwRONmy+C0mN1RZDjqmU8a4mJfNuBPR3OGwrYaaxAZ
q6xvXRI7hTwiusUij6hLVCMhS7JKYN7C4lcXhIW24vSmivH+Hl6QOvAtfKLxSj0o
qMv2Qx/ngzJQFK7zSTpxArygO4T1GhFg69hpLlYwsHTKg5UpiHfq4aNFtWOh+AY5
rjhBMeuocXPpujxS+en8PT7zH0HvK3yfd7q00oDm4tIANYBfcw3DMUs0ez0chxHI
GoF7w3avk9Yc7tPiZdH0jWDZtrUYWcKMwyzK4Ry79gGWDJmUmnV4ctJjTpiMz8cU
HrllyYqCXjHhDW8yXISCrodfNSZJJUYcDH1+EmfpM+WxRkhUJZzsFveaDMKj34mt
95KlCZNYlOTURZ/aSoV1UMc9BGKqLVfr8ZIfqSjYUqR9bgdUyeggu5s9mi0Endgw
e4d6t05T/ziZF9I6jcPerIMVWl9eIP5ospJ8Nbxp9xWoMLycMsk1DApCDfHlmOJk
292g0ATxQm4GvRVgV6Q0DUYQE4QyWBM/DzJBEBuMxIArm7Yny+PgV15ncFsK/fP/
ibuj8jpMBduli+uA0SGoVPkNjtJeI6PgW4SzUjeOxRp7w8AMiIR0kJkPf5Q4o8kO
3ov6EtZOetHM4ZoWYpMK05iw630e1JQsG972RkGURgd10t7bXYkC9A2mnDV5ngVx
e4t7fiwLANV8idlSXdBBnziS7sZdB2j0N6VjFMlZlXPYdKMjSvmF7NOY8cpIFSpK
GG+SxcvZLWOpSG/X/T9ng+IVvhklhhdmkLPftWx/QmhBPGCzsGOhSJfS1/zlELLb
RztxIW7f2EZR7gOCUZg4k2WSHgoZNi2e1KKTpmsqTCWNrWGnSAYL2ua3eN2bljnz
oEClyI4P0dh8GlK3KJAeDQHd91edE78jBNWus5eqaKtXB477MyEjmt+klS6ycd1r
/QuNoS177Agmdsc6/eJ3IZlpTXn77FTRbYj5sq2h8+tr5iRvF1IdA9xusws+GUbd
nggoOcOPZTa6KwdMwfeHZXk7QJKBVw3MsojumURzMdfrF6O03uK5cinQLSdp2ILm
l2EUAAtfOWIHEt4uY2Q9ED1dc3WnRUlSlAUFP1eArihcUNWszXgeeCt9AvqJwQoT
bFrFcUgKRDu/FfWC2C6xiF25n1KNbCaliqg+TZe2HJJw4tuJlmWDJZDYJjED21+h
oA5HECqc5ocrNbbn2nkt3nsRdkMjLZee1aa8W+cCFNZsAx7HXsT0zANhQLJ5bSCX
vmydib81Gaah77JNmA8ml56nta1mQujjzipeF7zyTRzaxMm0PWxHFCPEuZDsAD3n
bIlXcx2VM1nBvRJ4JGIOnjhfg0+PxHtxMW0EnIcnYaZ9amhirJjR2UQy/h8ww3JU
c4hwqMXRbmzhYnAkPZ/Zr3jAKqw6OfB4H8Hp6fLBCTaLBgmH4kwUO6tg5iQoGTeO
cOB6KmMkdl2bnwt+jwLDC6UTiKRNMs16SmmoObo6bIJslV4z2gzpmTnqe0Adz621
OaJ7+bd+c8k59Z7KGKRFZHCnP0XKaVvtwDpcTfaftIb6Lx9BB6e0m9TRH+6N12oz
FBHseIb7lJJw9lfsSEi1mPqPs3B+mH12oJyfMyqGXZb5/YLEbgGqZKcE4FZd0nu7
W1ayM87B4ehbQjvpJUhIWBz1x7S8IEVXFdc+mkWYvBUdplVoXbZspSzVR0mmLjWg
iaS50LzwqPlywodkm7igBKVo7ghv0ejlraVirNKBgQJ8Py1JaDOGHcji+GYQTipl
AwwQh/Mz9HToPqrdbIniz7tvWkRS9tCUuCPQ6xt3hTdZ3O3Bi+Pp+jHr7SvyTjJx
eT6HYQ09OXHvK/NY3ynyZB2mWUnr/HAYUfApDg2xMt9o8B3884+p/48Fhyvv3Qyw
VDEaIG0SAqEFRUSIWQc5zzDEW3ynF/D9y5DjMbj3MxpZSLM1fBp4pX+4AT6xesFI
llG5dp7HoGWB2b/06Z7/LEOOTbbEng/iPqSFoU/NgRLHrSW6pzjaPN+YfWmKqv/Y
klMJJ2HVunynkBoFB4+LbucPhZKGQ95mjDOiw+d+wNz2aq24AA5gc8nEucifhFtR
+9nLyn5/2tCB4Gb50eDdr/JxRtjbTXJVpD6WmocBmO37a4pKBGsi49qVfpneBeO8
S53qJQ57BjXiCSqZ0pOx8jdKIZeEuReUQHq6G+OpCSLy1TmBaQG2zUaiufLPqEC3
cSMi0fCUHjxmfABXUYuAQd5PgXejQ2FUTDR8YuZZJ4rUKMreTFfxY95y3BOLMUBJ
3HO2cHPD+VkzvzUMu8+7HqYyWK1GHmPMQdo5WZ03MJoquQFAv651brqrlHTcuGdo
tivzyX4in40r3NDWTgGgXl8IYiM3uTti75toFRwuMv3qB+x0vSwFMQbprK8Z0qPD
uMxOoSXusFKGclpzNR6FaQy+IJSnihhm+5ZVBis953JleMSME6UzkNyy3Fvvl4FC
9v3L2dJyHOecflA3AUGtmkbPQlBlkZJDj9dtw3stfmKC8ofMGfBnbY3ppULAdaBR
xFHcAEW8UVS+w85RpAxFhVdBU5oVe0vlituOsMhJLWTNLbIHQ7FPdr8oy2ZQzXZz
s/iqXOQA1fYN94hPRPrqBOdXT/YQyk7ZEyPzVCYx4OIBPBxvD0UzkdB070RAoSfj
f5SvJDDHRTx4wXlcs7XdY81H1j2ekMO19t0J7icAmNH67b8vhlQ/gcnkJebqpIHe
jahbLsQnNDUGhLs1cLOmbmfeH+v5+M35Jkt2jUzUt8ef+P5eDL8mf9MelVjhK2Jr
nBN7pILzlTMn6ZvVXd7dbpm+0w7RVqF54MYUPmabah6PJRUX36mbq0EiOOFK6Fkc
VhG4Exjr/OxK0TITba32DLTIQhSBU4I6T9G0Hlk6dNg+i6bMpn7k5d0xhHS7pPUj
l4ub3TuGFY3/xwlEKYfbHqBHmKHWcjE1npB/rlSHoESpIBfRlM16s3LbzlXy4jas
hMCKi66xmc3mF32CrOBBgE0QJqjvOeqpBIWsw76D4OCILa0cDDPWSvQWQrhCKuGJ
sFpBOSwe8yMvk2u7vqNHvOREd2dZ6mGRgmvIhObCZtcyHEf16NCdUIjRc2xiXZIO
4rrau90YCnlYSG3FSXl3DJbuuYvAukvLul8xfdmJdZ/RgGRL2eI29SUUMho8W/i3
oycq+wk1WG7EyFyr/BfTwnYjux/0193qOzRlwmGuZzFb5e0NzDOBlA9S0ZlAqP4z
BnwEKRW10Rrr6F+hk9PE7z1q/Vye+5fHKpiGiEQ4ls7wD/PnBRLV/aYAC1XtVxiS
oYh5lwp+sHeV4UgF+Nk7N6KaRoK2QWOHe3nFXes45Mb510CVGS0NEzIOV7OclQA3
poSW/cii/JJi45STPqJsXvAszLtMgCaUbFTqMGGhQ0pu8pYspeX3jkw3N816DB59
Nwr4YchCOVZv33sHqiTwYfk5dIqayVqB91Jh3N2hOKL5ogwoDwKpW0pBw7zGA1oh
4Hf8vep6B7nW+PgDn6LoDwPJi9U3CZJOKn5yIV7Mob9gl8KaXok+nTSZrDEQ7bsE
wcTIxyVf8jBRZ4o9+BvGQlD578q7vqxbUgbjaCk339AVmA27eZsK7S7xyBXNuFCD
OsYWm4SSQ2FlPRqlbmCdyFnJ8yfgwRTjgj5RW83TxqkPHd/4ApnxqgTl+xznG/1p
ZQhqBuowtdeZ5Bb0N8A6bROwvwot8SqUT9FZgUjIVLHA07VmxgcbL51a8rBgyc7J
OIyCnWXlVGCq1O/zbwZ8aXi/xbXe9dqIEEJWs/Za/47F5G1AEOy1cDo8SWLO9/Im
4Fe+e/GsQqMa9/jMzrvlOo1nUI2+NpgQkuFc1MBpfw0wZfpDsC6HnlD2krn2nGl+
FZe1qdcArCJlK2hfS4YYT00XpulxhflvjXk+B6w7mq3F1YIM+qLjacx4kOchdBCs
JXln3TC5eIHh0SQtdQo9eFw2ZyKCzVSJxNWrUk4NlKft8RjWG6llFZLsIsL5wNjG
KwOdtgjNQI3md8RZnFADSbq272WKh69SMVNNNjlIc8t7bF7TykwDRUXe6buOU5N2
THz2nQdcZ63/IyudNRt9uqxpM8EAy1JKIBPpxn6Z63H4JQO6bPfACZS4JR9ICC6U
Tg1KgwseDXIroQktUWKRrVps21UIboQVf3u4K2BVm2Ltnw3O5xXCFCktwKeCzF9s
ZcA8mVSMCmm3ql8okLRaJ1g30aXrEPemWLtHOcZyc7ZdPrUcXxqUZGVFNjzxn2lQ
PnjWa/DXbpPqBNeV+ksSgEQq/XPl8uTVsAcb40stvP5BQASuJM7uRdo/J7rrrg2y
DnivM8wF/xoCDINyxOL6s2PYj6iOnAXMRycpGvLKMimkPGZlH+BwHWwivzeq+/uy
cHFRk0q03DvrO2Q7q4Yc5nBllGG+sUjnAgArpKMj9NFjVIo9UI3U3qhPoaOWcK7Q
RrkLpLfeD+HDF0X4QGdKnbDKkhVFMpweStH012rTar/IV+oEF/gzjqOHXw0p25VH
iKBZUN72QdjkXUveofaHgor4guapm7i58npUh2jG4r8eyfYE/bVFTrESC7DZU5t2
6Ch/i5rrwGh0cKUoisZ0cMkHqD1AGyXQ/psGpaU1wwnyij7RBFH9+Bycbw4LOxQR
1owNX3b3qWdnX7Bkx7IsHFjjvUP4/DkhQz+l/sji7H5/tCqVk3cF5HgRFyPwo6CC
rMqFOEQkD1ct3Yx5wpwqUryVJfEYeqE4NM3bYveouxXPT76TZUfSmWCDZ6gYFwEB
dSNvh23wqFBE58dhgCgOIvnCcfFS+ImD7S70pWuvFhRK6CaUbFSUQBq/8M0Ye77z
RTGzxb1Isv728JtRwlRytysnyVszKyVW1Hdy28PZFrZpl0JMVnrqK7jp478lxdf+
3AZOisheNI+LIL/dBqIp0DhsLOrICQkmaOSWluAP6ug4UYs0DJXTiGcR7HLZZFr+
na4fAvOnika4UTwqE4o48L4l0mJyBjQRDXPBonyuS1wxlJYtynneCrA/lKtUYbeg
j8GBa6ExI80hhtRvYXbv+vauE78TNH7zEBNTtnA2SyHsl6zs3qcgMnZcSnAF4O5c
GhUt+Dvy64Cod1SUeI6BqB3tFdc7fr2m9WyIXfMRY28ShtbGYAWIztgss2J3SBpE
JySlLF/aNUUUKxFENmP2V/7eL9le6BG2yReBGnKbEBfVe45XyFQVuPG2AWDjUMl7
2BK4ofWuR9H305AeyVRrI+kpwSEm3M5kWnIgVECwdw75jxLSKMyKLA2pfitCB4vA
Uke6ddyB/Ce0cAlvj2nxDERC8PYS99/6JY9M/vAGFbb31kjPanhNxJBzbJXLN8m7
2WtH7rOZPuXRvdBYiUWo2WKNtrkmyVuXd/xsBOjGDxvqM3b9RgFzO+qw9ElBqXng
WeD1eMYp9H+80OOe9jN3NKOs7VPFmFp4nGzGO80U4ceN6J/hV0FVPZm/tcdBkNt2
hQ2dpaMnE9OD6fbZ+k1URHZyEE0mWieOsFuuJTsRyXAnIGQwXv+6+enD0WZH6H6B
mhtNhH3pqE69Bi8fyTYw1JOyraxTJ30uq5Rjt1rjBCJf7c4yisSQQOWfYvZW+6za
RxZF2dPnXsygdsAXkUB5mWs2WIT1dnT0jkdBWny8YU8GpvKdrlQDCy4J0bwbH1KR
1ZunF0uKgU+JY0o+qt/WakNfFAqq0UYv81xXUFRjdpAiqLU1FrVYZzgvThjlc4La
4S19n/tWQcqkKQcl3AhSNv53EOFjDVfK5duTghAR7DYqk685kqQD0d/H/PS0og+Q
kqioQoW5+V7IARhUez2ua/oQgeVzIe9NUXoyIP99NwLC9WrDzbvW7/8h0RBoC6/E
/m8BOxllih15KN1SWXRQCqnM2br0VTWFv6LC04b4ynM9eTaY9Fi74mXl6ZOoLMOy
1X6ZRnnW4BNse8cKMK4EgyCV8cY54rdvmf12JspJrTGotMuIaiMb5LhhjVxmuOM/
XibiE5OBl635zP02NVBMYqMv5yFbXPzzbGlKbMwyRZalGB6mo8jlpgqdQnKYQY2X
0Ruydd9dpVWX9QA9clf9irc5WVek2LXPDca4xWhwcREeNdUj57KbXVcYrYj/tap1
O3vmrm+Lz1/LZFzTj+jCoJEZH0vw+VODQqAi/kjjQns9kX9uChNN1PBnPzu5Y7c1
9p1v5jPPifAR629l9V+/DJuNMzpv0mv+imnXP/TRCZQzRrF3Weey7PCCVZHyyQi+
LWazDu10/kTbVmvVYGP4K9D5yQ+vuwJv9s+oqw1qxbb2TutC6ZwHjE4MDM3d42Hx
b7bK/13hiGmSqHgYmulScrQRBAKddCSkaRiH2xcjepA/AZJRxvIKNXx6GHtBZlZy
deq8GPTgLF30CBhmpiHlgi32/9PUyGLgxdIh7+L279Pjin63jqUWFgiSkCartvH+
41VJY+/FSxA93eZ+XyuASxpK8URzbnIdlUGEVX+44eAmOVTl7RB0esB9rOwKbfBE
p80WXc4lvdEd14r6h3ynT89MHVPz/7e+lCHS94s9vViLIc25LBaR9EhGS+ar8AGQ
T+6QNYwd1y/ITAG6HMxcG2sIbzvVc/uKEV+t+LsxIDWBEBTlcLcZcry3aUTZADcA
zBNLt/xj4zhu/EifKrbzsY7qrVVIr12Rbq+6cfAvhWvcp58mS3asvnHfDLU29dBV
sw3tYcosE/oA6KNHY3W204OnBnpL+i9fJmWq443bT8HhMD7gYyGaB3rbTq4RrqHT
FtB/WNS+eLXr25cuNLix6CeLPvpJYLb0S1rgfX2MEx1yWE+W8lZc2eri0qQVuP8w
juo4TM750enTeIjlrHDzRG2/gnvbB3FElog/ChkjQaGmAv0znqXaSpr0SvulH7DO
nrwq3eBpv/LF+grEJ+CR4ZZXUo1aBYRwWgCblsHutsAes7KVKUUbURpdVA486xf2
5G3uFEk1bSO04Uo0DGI+156lu6ts40UHbesg+H6hNMf1YN3CcrF4vniSpSvFRsPc
iVAGf68e+0kcEsenhfuN2wAKFMq3TbJW1OOORHIUgdFKZ51lfi8Bieid7clrVYlB
iZL1q/QbZDBCUkxBe4r87FCTtwRmWMx/cJ39Dlr+WpKruaP/KpajykpxyFOi475Z
KepLcvXrkFoaXst9Tu4nmW61LqwCqD75Yz65vYSabtvMvhvnjITYLckm/5nK8X+N
zsSs6Rke5EW0ZaHPnCBqEb8x8tlNfTdCiP4E4uJarCXTtSzkZoSsTfWeBBxEloE1
IZPc+2wA52d5iE57chY6CM25WM7p6j5dqm1rG0elyhrKw6cBefrWwI+a5MUgnzBB
uoaCtTGCLEMezXLROUfC1Df06iC8/9kewCKKtvVmD+UskoulY22wzbmlJPUOwsTA
/3XFMxSixlnb8c5y/rmKXfV+apAchjql8tGdYEUVVhTJqup3qiHSMqvjUbPiCVlh
SJs9qjgu4WyiGlThjTwEfu2A3NNolHnxzL5s7D7Gjom2vZcQtcO14t9bl6+gmaKP
1rhQh2cy9zfCpnosDtr6bbOu+wEqGJoPcXn6dVa42+XRJiBOZ2v52i9EBM0gEgwP
o+cMeG8XGn50dE/IzE0LkLT5cvL5Pr3t75j9YJx+PO0giFGIxESDxMFU7mOPr8eF
+Te2yaf5tF1rTYXisUWEYUa4x25TGbznDegYGzIRqzWPXGE/KX6fayH3ousCXIi6
zt9+I6uulRFvW6gFPDYGyXdEHWssX3ra/WmQW8wXSJ/e0FEdnUNEzAWM6s4V4SRD
oEKbtC8/aK7YXDhD1LI52HDlswDOxCkf+QkmSxKaIjxt4r4Xsz+gMdSRyBVP8d0v
NOeojs5wJKHHVEx48h/1Rql6rbKqPPt1MCpyAEgEgh/2TOAIakWQgCebCOEq1fWp
fIP9BIXvDVMQbbp7HQ4sOC9ANX6XW9Mu7pKSSfkEfmcghNLFdNAkttAp5l3KoGNU
2U8QrITSTHD/j+MZ8vwO4cb/IXSvMIMxck4OvyDcYd3KurrHI0YOUcysg/XqGfbY
mOt1ZV5BSQW4vsfWqw0iDu695tlQaaGnExMXjvp24i3CLfX5FGIkk7+x0OUjU324
yiu0vLscyxNT9Lqh6+NX5gGWcQp0Oz5MVRK/FsQKeyqtFgxYZa/b/hRrdijU2Npw
AdWr4mIJoIDQ/jViUvH98CblVH7lHZ+164r4h0vVig5zHD1NZLuBpM8wTygvF2EC
sc6G/JZy+jahTWEPqlQ8Aoxc+s15TaJ4vyaVGfeStwxG7vDzICnQYGARiAS3nmJ6
B9QlX+egXzmW1y1f55dhmpiFzGdvMGXZSnt/o2YX281BgoXQtHbZXFqrkydz2dGU
92xyGa1rSG0sE2SwVHTWB+a3icimleDTeyYZOYTLVQagZcwdaxJoXJYB7Z6owbtZ
CEPuLmtIbTWZ2kvkrR+iBPYr+miCSzMb8vZrHGIL3JQR6hsScjZnqyOXpfnH+NL9
rzLLpJp1N0PDhhKSRK7ea4JMyGPHt55gvCKbKQvWXXqdrJvX9r16QYHQdI0SN08V
fFV1ngZIRX10ZW1R+VXYqosiaRJ05M5liSb1UR45eZ8EvGEmLCt9O/Zm+rsescNt
JJU+jCSitKOYzdg/tBSZkJRP4BBhf8Da6ifylzYp5Gf9H7iuIlwO7QcnK4abiFh2
nNldNY3A8OuY0tRNqmICVEN33en+DqlEByoNyXDAOiR1MskN7YNyCyzSyCrpU8ge
ukq602rcUotusWml+WSgqLnFnLAYfCSmis3CXxq85QvJHeT5MI9ALFmlJ4K7QaZr
n4Xw41c8o7T5AiUCcnIUklooOOQEVeFo34xtPnSiB5HnD/6we60/q2uYrK0GZB0K
7KctzjEKywPHYjyd2nfKjk6dHYeKCrbHGouwfomykaMJ98PeSKpfh/PxzodudPVX
QyBHfiusK81sDH8OS/nYkPaWEX6ugzeVT3CkGliE/kM1f2foy2F7p8ekO+98CT7l
2OGZOE+KD31Q4JuySkgfUnLAd9nUIpXEtZjrZQdxta5kjYeiaj8rzKdZP57IBDL4
hfZS0ZAWfl37xWtDCeYELQdgdhkL8dn16T06GFMpErEh8oCrotMij5VYf2pKKrvi
T1ztnAJet4suU1fyFKG8EGd337jEcBhr1XLmTkD9DSmpipa/+3/XD/80/NHOyrUr
B5hlXKSuhF2D1N98fo10LA==
`pragma protect end_protected
