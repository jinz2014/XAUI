// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZKUTDTjWp3xxWSt20z+eKcelpkGsr1IsgWMeXptUTYATGMRxmBevt7RNvYVMYmcw
ziwYxGZ4hSni/R51yvlX+9Gw2Lsf05LajpFIy0QpvsGrlnoQ871z+LOg1+CB1K/u
DT9L9VllV+02H0iSuFcMxwpoGAVd9bg2Or608WcjWcI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6928)
CkmgjYkMoATIm2/ybC2NcCSwKz19KBkEGzkNtJ7Jt7W6ZWOzQC42q1BW4Nz1GUMN
J61v59kf6C6eJG74EV/a9vNJ+6WfmolPKoM1xUeoGstvHRtkpXaAb2QvOFvWjxuv
4KtMAo8cpSjQ7FSeNikuS+mt+PwnmlANzLsXmHInt+KaiJq3RWQlGbKx4ay6yhh4
tvI/YTZlACs5uUQ9NF5geEzORkfwsQ5tH9GNNJmonkWjx624i2NQPfx61pzQ5ksi
etFGerLoczLtXUaegc7vzSa92MnSBdQYZJW8sBldq9QepQ2mBPUFzbjVHZhin8+t
do7KqWac+TbCsKE7nrN2DpEs9venTf8NV27V12Rz7M6zaViLQkmyrXIouGv3yWrP
c31jnZWqSssexUHliShpnz8iAqeYFoK49edxoalc4mgojy4xwrse5tut9Ybcbpli
8HbkSNa0oD/gEpS638oxbHvtVT5H+5kdjjGtC7363O7iBdrXiCmdudXphkCRriu6
Z03uwN5gpj6ei8ExK0Y1CxXHofqcAq+drC0sKbc1Y9MrUmJJAU1XZyJu4AV+7+CB
LwMQx+jnOMA+eQelBWId/8sOjrhAT5WteO/pSxHZOXquj8TbT1KDF0sCOYrzWeKk
iFsSaPTHQ5LS6+1nkVBq52FaTAmtjlORfaZmBjScWgDBUldl/jao0GYpBOXHjxop
YXYaDGbWrAqswqtDz9NfjZxONeAXCBw+sga9Zg62Y1OguSbyPnHbxRM+OoRz67kk
CjiabsHZZhmIK8pcszAGfK4GzmTkRoyEOeawCX0hClG9vmXf3RWMelr0v8PDdZco
k4aSF9hUYJVnDF45Noe90fk2EganL9QS4TUMrywISbTR0M/7/bBPj+CD2TbvwRaE
rz3THAbiEZdA/9h+fTjUUl63W4+w9CM8iYDXx3GgWUu3ZbN+eeaGywwsqqC0/i5C
nK8xAAUuk1w6p6rnnMGNpT1W4LTYr1zueOe0JS9zFITEN8OwSeyL21PZP41o0iuj
NUICQ7cD3vrnvTbfG2CUtyNb6THqXLAWVUKc2bopVWfZVRtDhzxat7Lmx4c5hT7h
nQBcj8tqLRg02p538P2cZ6eGv4HzQonsN5SwlyQRMXMR/CCCWhK86HN7dCNk/G6p
CEYl6/jTyWGmuyg/AbfWfs6KHzFv8Dh/l42K55yIBMsOGgaiFXZrYYG8xYuM3KAm
jFL05EhBBdcCWfWYVysJdB9LQ3ByttTgkiQ/m93jVb6qtGMUJrnrJL8VyH1jI7UU
AGx3i3+zsHDiq4Er52sROSXU/hDWfCmFT5dNB6Di0dcTA4OeGbOWjU8lx2lniybM
1TPgya6wiX2XbmxVo9l63B/ivjwEA7Jx1Rp2FmX1Z6dEwB2dcWkeQy2dLs7RwX/H
dpygr+MQ9vPPrCO2uxQjs66nk7DrFzZctzCPEl7zH1qns78G3ahPa2011Corm9RC
Z0U77sQvSWI6ylYk76GMw+eVtye9HzB8PF9b4D15miVoHYEHHzHmwYf/KxbZAqB0
fEnQp5QwPO2xvX8mncVGEtRmHJnWYj2iqPMPmI+iO1G1IoB60BvZUFk25xEzen9W
3HqeiRPwLvsrwnShWPiVOoxZoNfUmYgaOae4gWvvm00cn5lsEdBSF4vnUwCRS+/n
yf0WvNsh5FwUb9rjkuRqJBUBITwO9fHKMHOCuqsENf+JVIDaNJOJ+It7poENTFLk
Se2LlElZWwUUprGRcJZFV402RaPvsHDr9mg5QBD6ie00zNRKPVkDNlyrEVmFxgr6
a7P+3wXc3fFw445OzVZo7VcTIAwny/ws5SnpRZP0ki5B4rX9Qq4ipjpvnr1FLf0a
9tTZuhNJz5wHiXjsx8dvSrBO2WmioiIa15+Wd4wbgp1b8PoFE1PvsVPYsyPW1Ufk
zUil5dotYoEma6GYyDBMx7dHsVzL10zx4iPe6XMTb2I3HPwD9zgPEJ5dAyBR1rsD
T46+Zx+ea44lK7KX0QLDXw4pj8lAUnNFm0P+Gy9pJBXCA/BDUgguxmGB3YTSOwI6
uwvItcJxmJxGA4zeBAE72hJ6mNzVb9D+puADgFMiFsec3uoqfoWF9TzHKJmp723T
BZASAvun7p65NYQHjhrW1sDq0z8G3MAV1rdE8KvL3MuMIthLLU3gAD3pHj3jsl8u
3FotVEeArgGtxOOBjg7DOhLJHVQXXrHHqOSkabhR8PG5n0IK/MuntIJUzm9D8hcE
SbZDHHffLc1aFSxqLZ0/Ovq/UQcQCxhE7sl5l+xoIG7UV3QeP3myQ0jlqzbahYVR
EPfTVH1A9Lj/Xjjq+y4PCMp0ficT20egwQMThXz/T6X66zXkbLS3jJj4ysCHMNIv
V9C/1XlP3FjW45Z08WLd2BGsYjGwwx/56PNbp84SMQDSqMDG/97Vt5pNo6hTFduj
ReT8WjoWL7ddn87pRGu+gThIweIyqEwFDea3kLrYeymCv9Y7/XzmMK5hCQCsifZj
lUliINuAaEv2NJlrfIfpEjqoDk6Lbb6uKgq8j+7jjYROWRj0mZQBvSOjR8mb1z0A
RXFQ+IJQ2/Ctvg4iX9lFKPK7Cukb++22g06lbvk39ohHRrU0hU26j+jNfQGhiiCE
NoXQ1Jnz8qzMvp+9rklAUHJNRAGMT/ocCCMb4he+ydoOvPtXWJhpNCROy8qo/udn
rah0CcoAsdyRpvhruhnngFhoSpWZTx5YtvHADIlbggiIkgAn4ixaUOJCAM057D+j
TDyS1yXiplBRALN5CXMsiEpsb8n145r4n09BOwyZbQwzvrA37YrVQQ/hvlj81H5M
jhx3TUn92in0HYuYY++a8d2Nvus47xwtXBUf50baSyVn9sCvEvChmj/ivYzdpvEb
reLqn+d6Ej3y4hsYYXCldNAU/J6tn7tQ/9JbkK8XjiPmK5cAd1UFsGT23ao6oS6W
krys8th4I4Qn6QsRUqT4731LeTJrBs/x8IehyLy8Q2hIXdveVN/wC4FvkT50PcsQ
sfEZ7hWBumlMSaivpgISo7PRpYyGtcOmbr15xeW/7UUOFa0K0TDK5jG2WSrzwLpp
QYDGoeOEsRDpAeINJGxQN+HhpemJmQ6A94pSJUEUG3j0EHqLa6apB3++QGLYpzz5
c8VMVRt9P1Cvtt1hugJqIC5w3AMsLrNmIjzVtv+IIC82GLx6sVyv6Qmz84l/z54x
gJ/kB34fgqDrU2186zfxOQDUdDvNDc0FW+B/MoRhMAGLs/p+8YWKcsXLnVktjK2O
The+SDV1LB/GzTAK7YQayVP+rLzYNT+ehYyWXAQiszKx7G0f1mxOSUbCVcTQ9KdD
FX2pchK7pbON8fmMGzrocbcEkMs+FZL1v8Jw/q5jPkEfxSKf9PIwf/e4+P5feljv
ojs+C8c4BNGwad1AxM92epQs3kAhMdnjZHpSEclz9j4vgAOvAjDjhKRHAPVL2zr3
D1DpLuxqMJviXpogWFGDRvfCWqZJ+NvopIEhVMVQOPD5W/IzJOfNzt4RX6hQEC2f
VcFDZyK7QNPFrhdDIYgJffKC1hsf76aEwTF69EVh3uDHECW3Mk67UMVvX5P8DY38
2hlB5WfK61n0j0lQzZEFS2Q/jjVbMrUCTYVywGO40DuiC+ElB47HbyB2laxh87gN
8j+f/dy3RXBnITCImzi4lr/3dtacKBtTId423tcKxSbIJMzv/q85QVfvAMkngxQ3
rRpd5E18WJiE9w2hd/Nl4VmRRc2med0xvN3i+IjWBuBPrsJbdj13k0GNzYZLSscN
U9OjIslBEfvMt3+7h+bsI7BYVvkF4oNqGkB75GCwsS3RiUPAidBZkIsEn1SpNLOk
EMepl0Kx3DugyrCJB1HQE/GEY4b2LEWXa3MgduIcrDqNWpYxRoVeIjkOxlUm9Ii+
XWE7W0+q8bN7ik15GSZiRDZJT3MflPMq3z78oVd2C8zZUknqRGgu20scyiiEsMbn
wmOe80VPJZjDwCSJ3J/s2rA1ucksOgulmYhsCatJkc7qqhngsmMxu6qVEacv/ryq
ibkcl4d1D8ZWRKoonmoGb14r64jur5tojKKe/co5pbT7V0XagSP0x/7tLvNQmWGK
+Zx2y8QCtQZE6ENW/Aj2FztEUVfDZaELTuCC/KUlBaS5T9Zve6bJlv8LlMLlPF/2
Fg9TrUocG/Bzqiw+evy1v60zopzMX/AGkDpgzHNwgHnO2S6iH4tWq0XXv/jUqpIa
YR6YVCyqOngw2A2UU1I/AcTD6Zas1wSawf3JrhMWHcTPnCRcQ6f4w3ADObcTHlm1
INLkEVYlzAoKiYUKls2enufF0GpjceCEF/MRu/j54LwcKNZe+Uc6fmndhpKtImkM
d6NkO2SOkFCU+OSRe3A1FTo4R6VGjh5IH+RQ0wPYlXX61q56Ze5vGBmionBVWF/v
zZhfyDDR2Dz7UgW/7buL5NULw+1o17JYt6hQtAPjKVzTeRkDFJowbLoTQfgPQKln
9lut2soJdxGW4p2kBbEtPGBiYTwnh3U/8q4MJF8KAPDObA3V077uz2HkY5KenvJ2
LFf4EuvNiRBRnJtYmPr7j9kwbrzae7kugonpykEYO5GVdtJYD6g1rozJ4Qybr9Tz
tF5E1Zv7wEXIiABeIl1QMBh7Aw0WqyMeYy2SrgEGaL9RyfjfH4uFPXnCDcNZY5T9
64t92OqXwJSGCMxcrKnvfInwnRHmKAgXFuOWqygz9YfexFb23aOx5VQ8A0U46lWc
EQ+e0rIdOwtf6i+8jFVZ07Ps5OLde7AFRQSYDF8JaQM280T14Aj8N1kKBUNvrM3O
STdFZ6LxrztD6vhuVs6vcQjviDharAM1199G2wF+ckuye2V/Z/upNBb/3YQ4aydm
hmRcLvwtZPLeonckPHxPvbabWVt5L3g9pntg86p2iPMsMUMav7DMXfSuE3D7Lm5y
GplbASg9d2RflDEz6UIEXuaroSnScj/1JYhgkdDfnHPic2swDVyDfofnJNf0BAIz
ztPBi/MDH0N1x8YBgTKs8pZ8sxBL94i3/PFkAzPmlfwaSZDLfxMGIUZXuATivxBP
VhaOAm05Bgvm0uADJYT1OtKzVrnXIaf7ltzjA0E1FAlbEkQT2DXbOUZ2TvDe65Ab
e66iweiqwCJkdTdm4rDPJ2enD85JiDrb9EA76kf1hocsW70GknLdoq6K5BF20w26
yB3vw4Ug+Jjd5qS/0/zIQYw6cSGRaDqkd7L5NluzpBvV/NKsc+ZExjeC0WMw5tui
EdiiOErhzytqXbgx5TvPCgGtLMnBFoWbLWpv1n1I8NzRoGtuzDhXyZjugg0bM467
p3KDEqo4YFSvX4Hf39LgKpSKdFAasfbltq1Kc0kbnmttT9Z5pk/RzG19J8xmzsAf
1em1p4SKRPY7RYL3EPerNDmKGFmD3orJGQq/Ha4wim41IUxDiX+mvy73hPPQJMa8
ON0nJalIuCSguQLfDIQO8oTNCWPVGnKw0ELj78OYRQxzxylQP8A+0D95YoMTNm3O
fttQwhNUZ0PTR95Bl9xNqgWj2VFvmB170NGqFHTaP0VOpheq98HLYyygZDaDbcqO
PmUE6h/l7idzy7RolcdFxiZ7ToQyjlEmR63vkfU6m2NYLYj08BF+/DQ3YC0HMEZI
+8bujd1y2RraLEF30/ImDJbnxyEkJzLJ8n0Z3DSpPpnVaKzkys1mMNSZsvs2DT/s
WUNm2Fcb/ZzdvxAO4FyW/BsHw4FY+rDfR9X27fi7eaZNSQB9nvHtc34Xg9rvWgPM
jjn22mqfyJDJOHu97ZlATHrzn8TWLS0MO6gNZcfMTPRGSzoj2XP18fWrm4N2+lwl
kB7+flxWUKpLMslB29AaS73FL4uRpJ1mIN2v8Fm0qzLUZVH/nQJFoJ5SkdYaZhjT
m6Dn+l16muro1L9m6TOWUZuFmTSGH7GiefY+heLeeS18TSKKlFHsMnF6g7YUk0kX
PR7M67Id4ZsBCw3Bo5SODLcDFuzcW/GhJsr/Y4JA/51QXa06wPqYrPgxjrR3ihZ0
im6vMszffUO5F76RfyFD+9TXC3PAuRLvJW+7ejFdCsv7nk+6u+6OxvqsbHWvhOqW
IM6xbcq3trOvaBfiWcyn4CwQgEWBNdWB6ghJo+KmIijr60VurRxivDY5VjHEKgmV
i7VBAb7HQkpwy9q04yDNSIIdGbvRXkjTn2xtjwOEbI1KD2iG/Szz83WA7UHW77SW
hHX2p43QuRDW0EwUM2jlG52xgBJotU0cO4d2iPTdqv1tfKKQcvm2eSSLR0M8Qlnx
bAfw6iuceneSJ+tQrTPVnetYfKwbdrF3mQsZ9WT4LL/mc4dLgj6pmlBaOPN0nohN
FRDjA5W2kNmkktBx3R+REnrPNY0HQf581+LRV3CT/nylZc6GgI1KADDzaV7CVRg5
bt0+JdOG5Wi7qSanvOUSy6b7tz6URalm1SSd/1EZZXbLoK+MSHeK4jJE6n+uPMvF
fAqNmrDCO5rff7CdM0LQdHsqymCoP8d7pT9V2Kg8EIn4a+gkAEupJdiAYkPG4CMs
SYorvbDwDN3Fgqi6fUf5GcldWCp2BPRAakqlRsNErfKj0HLFM+1Sdm+nLUOk1hf4
y07Dk+xX1JTr4UOwsCDrGgfTbR/HOP6nQ6ZMuHhJNcu4QSW13yMrQe3CVHJGngYS
3upWPyrmFdtG4s2WCHC13+KwoKu8SnXsZXMwti7yVOSYIAFGC3QbGjxO21zSVlsc
iFRoXiCvfxGXpG0SDJJnNdJKEnuvOMr+HMDBw8ebsC+h7yTCCXytzVnjciJP7vFO
ARW4dqjF2EMgzmEiUj+7FKpRE1Itlg4Tqr0lHnRjTf7TF6Y3bHypCmCGAuBSDygK
+C46bsJN8P+lPJjYmLt245HSXgyMW8GpiwSzQjUIuL1vQJ9p4eJee9F71hZUbt1l
XH5vVPRbAgyFcosOQ7xir2X2YGky29pQ7OVNn08VxgppU6x8Q3rK+GaequsPrDoP
Nug1aK2soJmokFo/3eKBSvzkGeCeX7kPYUZ0t0/pjONDEgDPasStIsbm9a62+l11
vsYVsnMFeP5+TjzRYe2yqt0jpzzK61xFsxDvuDKiucV82sbdOZ9FZ/uYaUO+SH7p
/OSNGS3V42Bc6e1q1LR1TyXmHfX1q+i5Xl+LOeV0FsMSrPSlxAYs9RRD90gw7Ylp
JODuxn7sWNdl598Wn9HtEq3q00fj4Lik+dQ0gLd8JpdFusVDTE4w0FQ9n4w4cnMO
3PhrY3EMxsF+la7Vuno+YloRDvkGhY1NKL2kg+9fKVyk9c6swTrTbRcpJC/H9EaX
cub4L2rAYe4gF3veDSX5HFYaQyX97h4rh2EU0FIN+gbzV7V/ls5NEo0aNzjp15HD
IRnpAPeJnoafha2V1IOy91mCzfu9mK5Aq6yr1BhsQGyShIy1qhM5omrKfuT9j0Jq
K9Q5b5pPjJNSd/O3zWdvGfxZvqPOCX+TmirKHChx7Ndd1aClkjHC4bE81Ymyhwx9
yNl17RifguMQZPE8ugkygic18Djt9Kd6wRrB+9obzudqRXgejUMvNDUUJzpJWsR+
MKzQYFQifEKuOEueUuwbYtDWwfxGN0s7pm6te9JqoC6nyECR5CX6YM7CPxri0OxY
gZWstbrLfstmixOa15LFJ/qQ5UHFX+GXCBpFN696qSf1CnVNMCmcwb/DBPuIjakN
2gqugkMJTYDXVCqVxDO7jmJsRKmSxYwmUp9t+kmwIhaoxCZ2Q/bL5S55S+rBY8IG
+KLYOpQjmF1Xupn60nWTsUd+19H2cCZDMUBZiQzMgWct5oV0jw0CAP89qv9zbobT
erGob4wlVcbylAJ7X7h6Y2PSiWmnKtie8k3OG2N6LTWbUlu9CC+3iNoej4jDWvq5
iN0Auqz2vhIuTe+aDpiW7iue3pAzQGJmAW5gsfBLulP/i7OEHz3OhhtZRN4cQSWw
+N8JbTCGjJtRn8wlz5IqxeECIRcAQYQ7BypkeqXcBeJhac15+mQC7qxsbyllAAa2
OLdzAxM5eZ4qu/IRrCYOXb2gX6mRHHfNWylzxEMJX5XKyPw1khJOdKDZnORCE5us
c/TZSfiFMbvIUlh34yoEsczFfw6U8GMehovIS4V23SKTZu54OT7fSnzRjDcZkz9G
oqRnPPfYHqceNXlxSbx02E1HZui0+fPFKjjJzucYAFYvTxK6RQW+S6DX1FtSrhTK
pUePu29iNcasA4oqEyrw+cNXnhv5HCYofNE9OQpCJJ7n6zWFVvK2QmzHLfnzqlDo
guoaZI8mmGi9hKW0+UFqZXhwjr+6BcHUa3zOyW0eIjXd0JVd2+HG1gjSVepL2MB8
klDBzOPWRFPj8G6wEpO8HXPomQswmvjv0NXK6Lz2jNYQ/3HEfUVDdIWLaXkml1uN
p6SKFZqphaMOwfQ/QHCz835TK4jDDVehvTLuo8utNDV1vHI5klK2bXh5E8tfi+Sl
SOmYWeNGsg5dglIadOAwtcChIY56On6O2irvDOyFklCAp8Dl0cpKX4gzeBkrtpk/
Mip2/9McaU46u5i3xqGmdRHt/j0hpdKcZlPRlVPk/Sef1xCWFx7hkVmgyY91CE2/
ppA29wJzg4NESNWUJtElbsEQ6cpS155xjxlrqkToUi7VHfPEQmwkdmlValmEeMP7
TmKSON/wk9DdzpmokF+qZ5aRYuEJplbi8AtWIIF5C5pRrZYyvDb+78xNwig1J0IA
HoA1sFjOL9VTn+7C7pZtMrEtjFyGpTWpQJF70EG6dMeQlkBNK0Iugc9LSusPsn7v
oaJ7i9RuBzE+bWcMpOeD9/+ArzvH7mqsocZrRYPAEuMmmuQNTaFOUMn2D9BoXOaL
kh7wc6Z07GbtJpUhEqUOwKP7A7iiuIvmNP1DtBSfFfEm6NELPudNVRWo9jUbQbOG
+aX8Etx9qjUC+9kENDPusSNI+YzWgGPn0nxo/6c8G1o6FlMRQrIDCEqM4rD3bDSI
u2husdW1Kg+H7iYvHSmK1ytPxNLMKjnBIe3qE5rl2HWAnpj84R6ZlHgjnni+VUtz
jeE0eL//PINTzO4PODuCbLCl0HHAu0JnlxngjSEj8RtY0zCreKeDduVt3hoROC/e
cu3NSdGp9bmRVzdsidWZr6nJV6qjU90kzyU2T9ce7RA/WFOzavGEh1cm8kRHDIv+
ealPmRvCVlazA0ryHm3/ja4hhXkRDcxAhE1kIzI7IKDK5tCjLb+5q9l6t0ccOFih
7TKlugZeXCArUILZgLXRqQ==
`pragma protect end_protected
