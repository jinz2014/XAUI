// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DFmr97fSXE02R++pYx3JyzNzKhsKjvJHm2khXR3K4aNWSVSeKU4NHg2RkOXsyksJ
OZe+eHaRabvA5UDBLBHuTj/PTO7ulCYn7mQgxEmrA3/0D7Nb7iudfRj9SUT0Ytms
cE1QnZ6J0DHs2/S+sPKzosjIxdK/SX6lka6NT+Msnyk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2800)
tNqWhhB1wgh9MzZhkxlObIp81lT/wCx+JQYYHtBcNUufBeswpZXtyInkgDNvOWm1
P1vjozsINZjueGRHMr0VBQvvJTi2qqlTB3XAiyw1MSP6A62GjjO663irrmicujWB
RDPfSA3As5Na0ii2MlGWTvz6t4kHIaF9qTjZPeksjZrGHVpiIQ2gx+3UDdj5sfj9
SsSf9j1ZXgPw0UoBFCTOd6r0BXxi1frklxpuDZHeWv0WMPqRq/wTWpM5cDwoS8ch
Ldk8jF3pt3C7bkKjqoaq+/DXLy85BHRb5JrhEB7semDRYaIxw8jhzx9DySfgox/M
60kd3BHtsOdwmO0feZF653KC4j4zAEA1Ua6hCzQ/nYOM+AbClofMLHCi+8L1O9f3
qBqMr/YkenlbMj9KdM0VObLH4rnLj0xpkqELkMi2jZ/eCxbUgTbqsrqvComHxA+R
9iV/6L2KPXefdFQ/Yt2Lw/EqXwpxBilI+zasj4AEF2btIHf6eNHRpOzmNHDdNa/m
PDE21GU1taPfELfhtR9YiGMUkzLOoo9YQw6Rcb4PQe3TuxKczqOequTZBebac547
BC09m/fGQEiSpDPEXm7fBHqg/rwU2sCoc/MDqDYVF/kuVXRxrKPvv0knD0dwGeGA
oVmCdUmm/VWShVmyLGxdryLF7EHGPT3sYX8okBL8wfIunmulAdctfgw/UJ8fGoTr
aV4sVy8lUm0hm70nqXcn4Tq/QGKrU3KWGTjTaudJOEbMyDt0iMTyHRlRcWnQd+8c
V3Heki1+32VLN0zsQBMlIGDIpgFKRrCBn9/fGAptnrc5AOel50izIoZU6YURZzSx
Jy2HOyYrBzLO5euKqWY8hYMhsnmKW6qXRgBnN2mo7JlkJUaJySeRgUWH1Q+x9B4o
CEbBYjy3B/uLzmxCEYvPZ9G4MXeQLZKauw0+ILVVUEQbT2qOEVLqbn2n2qAqluXM
Ms09qJROEymkv86JFoICd80MU8Jognjw56iJDMoPa7HyvL4dN6628PpiDhjLIQRr
NMhTi1LQULAJAkA1noeQxWdDQdj/apGbPhalDKTC0rp9PZ/ZPfan+tWXgWMK/dFi
IPnAd8g1FlJ2sUn36eYkBh+w/dRvMoyLuTGGKKmKvzTPBZxWmA8mdZbRMpbBPvXQ
nsa/GKmb5kakqjj3qwdfIUeaRPi65CSaI0nJntz2ImmE7ORd+LzphtgxHRw1E5Af
ExT5ERUPKhAodczni8IVohWR4aubpepxSggV+rnevEo1u+ahT+XRskr+v9hTRIFU
8C/7q0YYQSI+O2vgao3URoSekZwH1wG4VNGkOR0Y/YrCYSmdkLVOFEgfwtls9Hp3
k0cMbE0yRAIUDumYeN5UaSvnPHw3DL4/09z3WFxHkfzUwGhA8uS+46bl5W5F+6G0
ohb1vMlT2NO6XHW2anZdG2sfHIWckjBN7niCBtd0GTEi1+alj2IZoKQ1ZlVHloXf
Y6p5rWrZV7tmIaSx0x7wTzlQYs09gHrDa5t/1cXTk8gD2aONgCjjel6uISlJLpl3
Uh1Xl4q6a//VHg5gkev03D1Xba+IDyIzhzDHbmJpr+ZHVcIh9P+71QPINPNdXcVT
do5qU2F95qXGBRdeJPFk+XbnN+FBP7HSEX/f7Z3LxKhkWyza8Y9CeR1x4lEMQkEA
NzykozLGBBEO52p1tEiQWN6f57YAEmwFh6A111PrYl6fEXS2ETq1LNKabiOKb7v0
sCJ7bLozpFUx5YBboxuUSAxzBDPxqrxB7a0tqA8slCfV4jyfYjOZA9wMQSIpwv0D
MwJjTOeUqrnTAh2b8sjOmYL83JEXfNDor1il9XvOxNjR2QnfqoSvYyyLIctH0jjX
2El5CawtF5C9xc9ltDDMpDczW3p4yW4NwhUErf6lPh2B8kW2rVLj7GxrMzJdHBY/
nqRKRy/8RPTJ05VLayep5h28mxixhGFExm5/4Fx51qbDfP+Zy0VErJ6aiaF13QQI
usT0r2P7YRP2MBXg8N+XpbFVYkYT4fHOoOtxxZzu9ZRjLjDypB4Pu1pPR3j3TeyB
ba6ckqKapak0VJ6MZjqg4kH57s3L5BKke8b8R4aRRFiCfsHH8tIGBmthj3ceewjn
zx0YQTVAZT5qJaRL4fdhXswr8i+pPfdj9hYg/wjo9YtECEm9+nX/PTHq8YaOJeOc
TIhnNDOCYKbNOdc+rwD3t/lU1BmHP4iEZySmwrWa8+fEZq3iJwE2TgsB0ekjjKG2
w21/Knnj40M1Dxdf4S6JBJ582/y0kLCeCZMiHT9SYkeTUFuxlQJ3kOWZN9lTMl0x
b1k+3nSo4/2SHwWAb8xNMjsF6MoNIiRBOftM9jQctWquu333pOnasi5vnM1We83R
yUNq2vrxvlmZMShv5T0Z+56DBLP0ZQxo4+tdHkMKJcvjIEmcbTXHQnXX0NbbXfrz
7F9jmt9MWPdxaz6dcGP9I5K0H7Aatd+b5SJe7dwNtmSLZU4samR6vVs4tT5cadQR
NNK9XKuSTnu8LzhBL03jALBmgphRWCPVGZvy9o2H2voaIFT+s2Nre6mKLds0DuCg
zfFgIGOKpwRdV/wrfn4UZsxR4zHKS2cK2V3xqnE5iauyi+hB+nJXwWY6RNH0GM1+
XFvaDBVeo1FmPvMCIa5nYHLIepg7DG4UyI4bM6zjc5/+xsf4xDvbijDP0HR5ly3k
m4L2C7k7l/bDmK9Fi1ELfLxvojZ5ceAOQrD7PZuduy0O8Ik/DsvvyGhf1N6nH2ep
N9suNIrUBnxtqm5g29pOYF1CRgLDeZzi/ILkVTC+seLIjTMywH61lbaUAhDmxyG1
wW0w2cE7cxJAQY/DuhUfx6fJ1Kj6Agz4wHH4idAs4aLZeOJivRPp8EU2+/mTOddo
ov9qd7cukQ7mLwROEH80oOVqD0/DBBMb75YaYE2XbVabK19dkH11yVpRTLfX+xDQ
zdFRpUlXBKbeTvIK+f3Pu6FbXEz4Jm/M1vmEoDPxGjchhOR3lCgXQUzWAzLQnLpi
c40nHcdv2krogKjVJhU8gx3LXZNS4NbsFDBqOdyZqsmBgIzVxPx7Fdf5ei9JLeUX
+12F4fSSxQC5PXiw//X/FLHc0na7a+eU0xWPpsQ6hAflZnmA/k6so/Y2S8+t53uk
OV4NYY4QDpmif008ryg6U19CFfeQZ9uULugI7OFD1RaqkW7XLiPT2VlADlzXCQ+n
QZyRb8xDVW3xEmrBIpHPArF4XABer7SvsqL+ymsdr7U82qhK98b8hPT+i4HnwqsE
z61ixRjG2/i7P8omMD6e2fGztI/ICbul+mPCp1/r7R6QPnrKmXYQPXMe8g9J6nAM
TbZTxd9t4lo5CbW/n1O0uqxVyw866/HkOmn7DPt16mr1fXcYMeEtLjs+NcVMPLjz
cz83QypgfW5l7chM5DxoomQlXY2N1K/J+gwKuSQsvNZWIA3arA/CcvNgqNQXTSjl
dSJ130QD/ZPWHcqjpl+8KnpbP6MEWjrLyXZHqWANVjdmDL3daW/TwADUSMT8veZ1
rk+VpjVjFnFrC+3Wp8GoJzXZ13j8hOXa/IumUDAucKvuXIlz6ePiDD4jYuyWVvcE
Sv2PkKQoVD7l+2IY0+syjMWi+qFXawJbXXKIzxdoS0pEK8i0fcenZCQShsTjAHsK
zGuJ7cAZD24RzmkRUpiPbbFQ2JGzJVMU2gSkstUucbyUFFNsr5M4r0PeLP/QV5dc
Djcaj7D3ONdihcaeySY5mg==
`pragma protect end_protected
