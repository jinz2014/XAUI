// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Pq4Z+2jnqkPrbGV+hFceeEMv6Ss3tuUvbMLshylXwOPbL1Boa/RuPSlQuHA7Kahg
n4rpLZnewe9pYylnl9Hdke1JfnUIrmcvmt2n6dgJ+qnshqp/c1jx96J+ID0a30ZK
rfgsv/8AYd6D8/F4Gb9t9kfNg3Tux2I6tYeHchULODw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10320)
O/CqoT9SEy0QhvQQFbOq1RQV8shjsAmc1ubWW2kkGLC1OdqstymzizSS/QDiQwN8
T65eBcw+JN/lsyEd/wpF/D8xJj7AfTal6RSi5xRSn1QjiKuzQzknO1HBcQfd/tr/
kZ2H+sIGzASOzDDMugTj49BXyfQVkASwcvPttZidBS2WXhTBn2UYlTmsOV1EkqOA
lm1QBNAOVzNyNNtVOSbKdlqDSNSCslnwpxVbQld0dXqnixo3QLZfmzHJhkpt90RZ
TCDIGxtqnmhZmjS06t6izh6SmRs1o1eSYGtCJjP0QO/+NUZTs7TiYWYg/5VoV55J
ro/jTLtZQQMdDdRGmH4D4vVz0TMLgIThYZhpDFh/9CvSYJBa6uJ4C4EB5/V5DCyu
x+VKl7cY9OcSJWq8mG5/MD0JjAn2h8YaXEc0bJpMp7Vkd5zvQwenS1MB9Of8vMng
Diyrz67ucyvr7r5e5ipUPJcWtpaL4K1ZXiTL/N5mmCpXqL+8l90nkYKyPnkGpOke
NsJ8aORDaeWlfQvZ0Qww296pEHL/Fx9CZqI6ysKLjS1zEvFcS/2ZkVhOoIZz+7Fw
27isOvqeXXu0QFI9VxzJH3J/56aHZraMxX0tpKXV2KJ9jBKdD4qMuXjHBfmxm3x+
LaU/pCX9jvBAFeFNAS+8xOCah5OODZajQYizqoTY3NbuPAIUpdzHVO/IjBsnFxo2
+kt2uTIQBdntRIxR8G9053ykeS9VBzB1p70hJ1MEtNmMgpSKLionHqgaF8GeLkT9
pFtENJdp8efG6/SxcxoCJsoYMadalAtsHy3XYpUQZv57SzSMYtFeFhg8FY4SQr3J
OOzN3rl2d5dpmC9la3ssIEZo36JUDhi0djMsuW+N3Z/L+CSocw2r2hHwj681HFXp
G92QsSvq5rvyy4mffbPVzhPW/BsmoEdOyROAtBSQV4kI/BDIfNRq5hi5+QXdBggc
VaDEQm4x0mr57eh8SsPgB3Y9vvRLoXRBcb+0xszYJjnn1ZQJeGtCIZFLr6cYCm1S
6l9XO8fR7YicZ1cqaegvOxa4GzeeBxTZ6JkuhNcNNcOvuNoqhCwVagdzOFPQmmSR
wOlxVb9vWbo0BAKnWR/I4T81aaraRUaaUBL2QyXug2XN59p2VkTE+bUodFnKUu12
Oq5V7LCIxLrgbeu2JKTvQzelACoTHAhPtPEqb2F8Z4m8W0HU/zjCjYvvpG3d6Qau
IblRgrvrAtVc2amHGJ0DmcYuX/zk1uLJpxdI+sFGqRUo2VgBiyE/AXPlP4p8sI+k
aO+81SvFQIpLSsUd4ULKx9LCtI6N/5h/o2KuXN75hZUat4n0IFMH9hAGwqn/mQwr
KVTOawyOcZjoUTT9wnEg5CYirpKXu7vtKgjpVd+WJWm2gLWw8qr8WlvT2UqNyYks
CKKp6pacAMkGWDJ7MubK0ESK3TAiwd4vLPBWuN342YyJN5rPw2iOl1obIkPyaFgO
MST6xY4zb/RzKb+cIoXAOiOEvnScSXnk4yvr08pemnce1lNJmRNB8A/uY0aKVD96
9Y8Dokb/gdfzZ0wy/FkED5Y7+DOvAv4OhGdTyK95kmGZldgrNhXSSXYj4fEQg5Kg
YbcACDLoQ5WSKWQaFNvCQq1EiuGU1Pb4sneIbUOh4O02igXBkX2PTm1SoRyAMYGc
q2L0HzuRnTRWCspiEtmF8vVu+4TWUhDUKL9dD2RPhsmBARYGR+H2HfI8bPrO5Eh9
Xx7/JE83+h9WAE6g6Yqy9XF4zyHBqdy3o4I5FcSJ5AMRWSJBuFHhzbc3MV42Rlbh
oWTe8G3s9HSuxUmcqJdFDLPvL3pmknz6FF6Kw3APLMslyjiS/brkMCpSm67WoFEv
ho4iPhI8C5GCRoru6qIMpX3GTFR6YaxLz+Y5S08udfObrqMVp8YkIln8tiC48g/B
1ryvpDkFqr9dZz3BK7Qg+j55HpVlKgWo5G/Rmgp6tIIUKQS/NPuso1WlQ2DJrkqH
EwHWH6Uu5FDtoSpV1wewtLy15CjPzVUPLFtjPu3xOQ34OCjbA9p4rqrRPwdN8mLX
9OUdPIr3/KIb4929OHfUOlJQMYbGacQlNM9XKCLvDMR6jERvT6iwh5yGn6NRMXXu
xtr3TNl3UIPQ5ZI3yYpYiaICa2zCepAmbZQgYBbj+KMHWE0dL5r/MU/kOYEHVvsT
14o1be7uI+d+M3M1kCvmjJ+vOf9KRIGN/qYFRqJ4LXZm++5rKBm10H/PmDmpQr19
1jZuDatHl/48vtmbWTOQKi7W7Pj/RiNLCJlrGJG2MxrzgawdA6yvt0kvDc2Y5bf9
LW7CuzGxLPSmAOhU7BunKoHQYFOBPsHTw7u6dp4+2QCkdMup8pcQg0yRooc4XDJ4
xOZDMKftlRFed4nzYKkK4SZNqHk9m7mTZjshdR50orNoMBT3UYq1d5HHfS91zq+j
kYKeyI+4scgpYXCl+olR/mpOSDr7NBIqguNI9OB73QNIVsQgdyJnYHbNLN85qHne
l61whjXsKFtYUArdbTnp+1KSL1KDmjPbIwJOkOpxrEnxq8Gi6DH9FszldGSbJEFQ
XJggCFcKGlT0QNL5/sRsGjlHN8xwtzDl4Lsq2I1m/a/XL4vChO9dXujKgIlOSkVq
3iJDj2iVTAmX/Vi+xnYxbDejhb90u/tqqjUF2M5k4IHRAgGGEYki9n/6fRXWsRs9
hdFmXAg8XPYBcjL3JqFxYqK8xPYb/Rhn7O8FcjZ70Rpn49DzSkBgSCd3JN7JvK3p
RMkkBMJ8MeeGSUuVcUo1IO0L76e0H9sP09juuaWaWgW22OE6J+03RGbkRW03RdUo
6/6WhSZSntGmBctW8v57cEvFkb+gHQErTZ1I7NnPBCEuwNZGVXOHdWBU87MQLo5t
ntgGjR8R09PHXFA1g5bQMjfOzIqYhxlw/7MIa55oXQ3WaRxmXYR9Li+yrD764fkg
dmhclolUEXHchI0N15PKGlMnA4U+27YF9Ye2g2gmbRiakS47D2N5WDqxX3ZfB5Tv
slQmthstpGQzkBHviFNGTok+sIiBf2ajpyPz0bpRFPqBtik/EQQG5SLA9+P/+I2N
Yoy3NzHSH4sir4bAaME7TrCx8fUhd6O8PQUXpWmfAl0kMtXs+o6nW4bGIsWq/MYd
27Vrg+4g2sZMVvFScdGHYh9JM5c46mI12USFzooaYucZOY5iGjVPubCv4OK9N40r
qMrPi2nR8nmn/zv+PqlGiI5mLcsPB6iU74PtlrGeI55HztNt554ng00DzLqNuYEe
hJg6yPUlUT7TVzem3gYIT+kwaVTe8GvUjlzUVPHHrC6RruTSST0YGR59BD02f/bw
pLkul9v4gEYVlCmoq13kUAsbgl+g/E+9Emd1Nc0po2h+n+dCFzAAO0Tx9i/+T1Zs
YQ7dIkZ887MbtD8WeXO/DmP62QbIbFVJ8lMyiO7KevUC4Yc/ruk6zTT9+Ic7sOdT
nxFiV0HfZzdCOvk/P9FNVizLV8b/ZFWUWCr+Pmg5qzZq8hJCFpeuqwBhi4ZollYK
yRloR2mcZsubaHvQtQsGmPED076FV2nWcjfAuWlXH4iGPDOOJ5RI4qnW9ucGnZOz
A9GJ6B5z5zuEYhCLs1bJ3tfNApg3CJm2i5x4JH9GEWVs+llAx+OxcrcBvlw+zzLx
u4UVquzbfIFLNLc67hJIqze4qAO98g4X9HPWXR+S+LJHnG9ZF/BlbY3D6VLw9biX
SO/18j4sQR0KnNBhH3OR7+B7tKDPHhRLf12LQwpUzSel3sQWAMc0yzL6QYTfuRf0
4UMdKuwjNCT74LRCSRhpwNOrYc/9goter4cUH6br5YkBv0e8PuN6wcGT6ssIVK2n
pGITsZb3OKTZNkkkZX+VN1HurEbVBanty6OHLbRMmAN16UKxRQb+dJbE+Nt2xAux
w9LXPoxBxLQjD+doR5ze3YDNsI/fFkQV2lHArTgxtiFrpl9YIbnCLPkPHWzG2mUm
3pjZcDoEHyKnJBn3VK/CIcWIVWDah0XokeDYwL3ArIzzXcxt72mYhebHEFuPS2cI
u4ff1fQnHTTOj2g2vitqnStMXWvKT7KKC4mJJd+CEsrROpWvcbUOvsx0g6KhRKrN
A2fNmNGHZ0PNe9BD4RRmgiGUoW43Io/H6OnWaoNLQOaLBUGkXktuD/awWjqba+51
q+ebPljA6M6LSwRzR5O42HW/KOVnJJjlLyf0M4dCcJFJJYXKiSwfgigq3hYw2TCn
4ai8OFmzJvuoFRNcNyUqvCnZF5rMzFzw0W0bKjBQU8mo3vMRUNV0q6vE8/yl9y4e
cqg4RWpTJjOwIzNi16oesXrhnVcvMkL/HFf+uNM0/CFMpZbSrTmks6qDUEC4Q81f
IURipi5FUIUvuFQOoiNKcRW7Rs9DVuBirbfeKEvRpgbV0BxX85Ki+2wIGdZRbuwo
1d8c9FfKI/mlDr5l7+x8Xz1lB2z+25pvbyc23oOXbf6pXa3ia6k6/ooxL0YaHJm2
wKsS8/b2r/RCAaYmbsm/21QJ5j41vP5xesoUYI1lJhSL/3sOk+za0G9gCmCqVKMJ
GInybNvUjZ9o6xgdfE+ApGGkM9WBaUb8QKYfr06jEztOUhKG1O45WCzav8QsJi43
cNE+8rXXOK00LwIjZjzGTqO7yn3Ing9zMwm5Pvhd/Y8+GijG54C2GjMxaqgGKVry
kLOOsQvX04/5YNL2iggrj/FL/f6E41MFflXt+rO5iT5/IinYXA+1jaSBlnd0DsAg
vK5hhLgIdw9T12FvPB7f04chEuwO9+oxrqxurDNoOhZgr8Y1nm567vO4rZcKjnNb
0BA+MKsjqfNbq+OeyXKeFQ8J6EV5Dleqf8ytvJl3C5mT/nZIhZ2XI2YYTU+ha7lg
4OwQ43E6PimwB37kdynyiunJdQ5GHCR3wFf1M8OJjZgUgym0cD+HZWLpejEqgIEj
Y9arKiXJ8iwY9omj4kziJmT8E3dQXzXBnjDj6chL4l3rJhT+6kObImoEzJxHZPzP
ufRh0yEWJqIQsyW45K8Fog5p0zouy1oLbSrolspT+j5wjPmoP0/2XsWFm7FWg4iR
h0x1Y98a22rDt56YOZuoa5kNrN1AqxT/g+qN4ortiMafdIAw5xK5hvLuuND2cpaL
ayO90T7+PskR8whGxsu03Js41pqYqkcxbmVEM63hDC8wO1V0Ca30P8u8i8OMtfbV
VDuLe0NmJ5G9nm8ChgtpTWO7Vv8q+30j/FBFTX6OiDJFFdPTWEDPnqk8WxxHXRQJ
u9pFY7IWMXeCXZCW7rMT++UkHCvgOB2aPowbo1iYQzhRzxDBSMVjWrRXO/laKOK5
7OKJ09ptiGs9s059WB6/Skq1qT9khueaaxNTbL+S/++xbZeJ3pK8Z1BAbHEndq/p
ayLuf7V892LDLtJUrtxHSaSxybIEEIIq+qXOt18Mz7GEMqTD3jUsI3AKTDko09Bk
srOo4cUsAZHJO0xBJAfLwVAAwoulklQWO1sC5PY4RN5/eQWSrRPplD7d8JDfGIIa
ITORUaSEtt+PFB7l2TOYrUzfK0JOrum7q6DxfJRh/gUMqc3uk4zcUeADES5uB8t6
5xAr8wtD6yexZWS4NJiPIr0EiFKjnN1szurlrp3kp2quTGcvoTtv/Mb7+7dCd5oj
zI1oREezvdwtfcgK4prK68DNwgHvWAb7tWM3BDm3sVWLG9dN1EYfYQvC5LSYzCwA
WaYF7v2eq0RhLZhYjTlNEhdDhPw3tejMnTdeCdYo7dz5/QmEeV6C7+38UI+OCFhR
gNZ3dX7Qu6TXgGW1VpnBvwRNGmN1c9IkxwJO7cHIoY9tUZgmhe/y6YiQpgSANvDh
PDc0MQ+DO8tgxYyimVw9wsXvPWpStv12A4A6HNljYE4FOZhAomFnSY84YOEkINLE
+Ez0UMYtfn3i5Ghhx5DxuThXiIUQVGaqL0sf6LpSYkpNPKcHqX4HJuco59z7ahG+
nrO2ui+3lhZvCl3rIs1HSwIBuCid7nHelD1lnnpPSn7sQOuiXKwInZctWmcrbmGh
EqirR0KWpealO1j9xjtrz1m38+30zZHj/DR7ICiHQTwMXPaSBZPTN+AZgPnvxMSh
TxYwniN/2plKiQgsdIV4YqvQnB9JJpprhKKD9uAddcGVv846/53MRVsP8Haxyi64
wh11PGNhgbHnqgB622H9N0q/6pn89oxK6IbStf5Ya14vHq+z8V1BBo3uFTzj6FNt
zmBdfjAyXiwV9iUYhKIGJvOlYhU2NlJB2biy9Sk/cbokCsYPBNRz1cPWtNDWwjS2
itiH8vYNIm0QXzy90SkeKQksoPPDclB2mFJ4N7gNIEV6Tblcr8v+6UXWaFMBibvk
cX1Y9kGEzQY3PzK2bjXc+sJH1bZwAlH1EdUmb8aYHT0Un2nAUfYUNgtEFLhjjqHt
+JZiGI8WVL7nm3CxhqSOs39A7FCid1dligM7HsW3LHH9UN7CBR6HL7O8cS/gjis2
D8pET9C+jUpuhI7OAfC3insScWsPedPMN9njyO00DXUBywsjH+RApnfK+7dEuF1y
E38WIa+QA6cfRyLSpXJAzjoIspOxt3Bjf7+rMotNicQruwfp1S62WWhezFnQzBS9
0erp5oftxqIBEs0UeeDlmo2ddTC6gVBtD4mSL4+cfsIfECJdBtnZnu8ne+RRoz9d
r4Z1BudApqhRHTv9dCcEACkpNnk2oK191f5wCejbn1CsGgyoeRv8dmTGIerNqjeX
BZkkCgodA0uiGY4c70NsS3D2bPVDNTdWJdFmRbWESWpAWuXpLmg62T1Ig8Fi/BlT
mo3YWOS+FYLEs1v2QZjuCBj2+Gl5YjO4OoIuwyGuZ066Kaaa9ouQ07CXgXjIMuDu
Ty49yShr2gSj89KmjEDpZv9dDmnQpVSvtntW3A1upaf0IHN3FisXD8HIdXdUPXp3
IbkqdGUEkUpcK8Q7ta/44tBl9ChDnsyAKGMDTvlt9CkClGmaxiVGYzmvDnfPsZFC
G2GQWK8Fbkh42jmfnZxWF+b7gd/9B5yTueOS+F37TTefoLmv7+QlL/vwJIE0mXuA
gpvEdZIc7VJWgN+qIdyp9weeAcB3B82MJIFY2evieXEEXJ9CYmWN84tKunPXSS/Q
EN4iDPuvjX9q52QLFNjlwnxZ0wOqCyU4cFnCuFQ6K+BNPuIqCMwk1RqOzvt5aZKG
ndWWwqS61MXMn9lgP6BjjmF93LeHZ33IAvILIPr8rRKH9XMLnlZQLe7hXdgK+S3X
rNtXn5eItWHPAQOOlWmW2tsyOtIofepMxR5I0+tGGEB4XFl2i2E9f9lzdyuGnFKK
ffYv70U+RvPTQ0XTkJl8g2wjkJ5plGfQftzGr8Tw6UbVt+46ucffcJfWHT1kPtRp
1JRI3VEJUOQRnY2oRHHwhNyBhUaV05LiVOgt6vMYkiVZcvbaRP5YuKTWQxk9y/pP
xY3pjsiD+MPBOq1/ECHJ8PvciZ8G/nCn9hio8TRzDLWjDf7kU+EF3VNNLIccqR/k
k8zlqaSWAk0d4OYcF7cznojUm3JUjLzTw0xEji4+1r3D+X5doc7a+LnPEXYXmRPk
2ACHgKVEJQmAeNVIUMASP62rx63SobBgydo+7uG4tbzKq5EQOF5CKoYXww47WMkk
AMOh0Reh5rWEvtGa+QgPnOfRlVhk+fsa0fcHQivFF9QcJDWdyOcHB3W/wXKAkvGj
8WuQTYDvO3WnP3xIr3zFhwHTvPnCzAIaivE+Fvb2ly5TJQKAUkF4+GM5OGjJu4LB
w+8Fd/uB7oVEUDzX8HL2OVrhzGK6eer2l94W9Nh/EQuACgizgN5Aoz32MmUp5rtr
AEkEd920/g/bwuLrhLzZdiSEpXLt4O8ivFKJ/1eOEFcyy+3znmucyWxAbhN6S0ee
xbal54ciKOeMpzk0HfPb1hsXh5X/EirscIzj7uxTdYEPuvnTvLdelDka9/Fjrvco
C8xmhrI4N9UcBvAXB7Sgt718cLU+QuR1uex0d0RJoXBbYi1wM0DUXfgA/A2PC4BW
oUYR0hYcSEPPA8TJNCTB64/X1eQ5fyey37bih0MNXJz0bwNGBUir+StDGvEHzpzK
iNmKXyi2iqY877hmMonlDR4F6DbL6Q+oUavKyWUjJ2iIhkJXbYF4mwuqI6w2BtO7
II/z0qgiIIEdRhKFnWrnjUYQZv2gzwRZjWtED5VxqLm6fU21U+8ZtfYYamh0bw+r
eIaA34Q9creGEKTQ0x9+JPij+zEKIHyQdjCJnRhOhlR7swmbLIOVRKxCGyC3cw2Z
C9QdUrt6tHMq/2mB/4O4npyKX3mmavXNLXm18zNKk7eRuthaE4ms+376ew5llrki
nzlUD7S5UMqka8pytTHJRZhiKB4bxV27WAfNp4hEcE3L/6ffVFkKG041tOGlRedm
9oJ3hRQGHs6f8Ojk3xcZwFyaS/ktX6BX2Vi3HTm8W8UFQ+TBDm9DR/rBMEuTCtFo
I9HzHItxlJceQcudviRhfg/z7DPiYfSMc3B/2Ke4QZI0e3eJONp+Vu+YJ7K3a81W
Uo7OERfyfb+G+FJr2QThO+iefzXiUi/y7tAT8rbSAXlj+xyZt7plWBRvpbWOsFjm
A3XEWrzFixjYsS8cYl70ktA2M1+SjS5oumdREWxPgT+3/D5cys7R6XEt7WGiSO5U
Pmx4FjnzscBSNxcjfh5Oi8j+OJNBZ0zVvqegDdQAgN0cMMdysZcoKVUwtr6mxPn+
n26Q1nixvG2BVaV7+nueAuXulh0anPvQxfPOR+2d1kZu04xHNWu52lBcfijvFYj2
Vb8WQ7piEdYDfsU+OrHSKKeusmyzZh5jnAoKO1P9Pq6VG3n1ma9nzpnFrHLi/kkv
Bl+ugXivtNE2VnpbmUZfrIcJyEcIHyxkbyyD4aQhEjad2DZdn5QP5QaPh5KZUdZY
DPuZTdzQZkUTiLKYqSFbAafyiBe3gqzj1JLecb3Y79t7Tm9PV9w4l5+zkdmBVAqI
gCjNTl6j6NyuYO+E5f7zlKLeUr0U/cUos01Ickudk5mgS5GFgUfPqvIRDXngUNPP
7EBBUb74mcgtAWJCrK7UHY9WPpW1pUDCFk3iP9VuV+OjZ/54fGOFoh9WKOsILBuP
Z1XjVOt1swynXrsp2xT1hU8Ix7hR1H/ElG7EQ+aFOuPMn+BenOg6gx+VygQa//b1
wvWvRdTHm+eKp0rRCWhna3zQ8WkLPO7Uk0qNZQqesxSlxLyNibcB7BHgDH7PV1zQ
byoso6sWkfp946b9EckD5joLDXK0T9vU1fSpwceLWTYB6Y6dJyQSwPrF8NqRWJja
cFsLnViUiZoyafbWDTrOyieeMvwDiC7h5F/g2PxMir5yQ9dG8S80gX9raakLFYgE
nRJyZh2q1BMSDZxw/MBuW7K2TKh+g1fggRTgbY0Ik1xqf2KD7RIhw+nAZTcBhiyO
UCSo6U7PZzFHHU/lB8nzKFWtT49vRmsNikg9so+VrcVaeNgJpYu13T/6LUVbLTl6
8at1p0biZYfh1GizuevlpH8OZvv7dgoSEMuI8gplY6fLegIPQ+MN8Dh4N6PTdYLm
49J0KKuPNgo6sP6JV8/gsdYYPTo0HchHV/LU8Jtw5SRAVnXdVaXsqn5xRIhYbUp0
XqrPmhiSavfyIWd4GkeEZIObCeWzaVV/dphh2m3Xd4GdT1vBKjKjIiIep/s0mVkz
mX0W9V+d9UhScDv8hGFXV8M68MKauwuy35tA+swJIX7YXJhUhHlUTnYlpa+Pd48o
cPDOde7JB/L/EIj3wVzpNuZLhqc1m1JpZYZ0vMOUC2b43tuVWtYrRA+/NRAr/HU2
srUglZ0VfjUfDOzn9v1aS4Uy9RonodcZcrQ2ECVfM0/XKh5ZrH3iLJS7YOOMjz4v
ef8EtBHqsM0YZeRx9b6V/Vrm5GKnICuMb7VSJKnF4i7dUSE7QbhJTxu4eXQGM9ES
6aXUdM2YZUZSQoypHr96j+s/RQO5PBQgL+PrMm22FGYfVVx4XVRYfATzOcE8tsOx
9EaIKowmSuofaJ3nHAO+j1dH/wVFh6UgI4Xpu+el0KUo3vbyy4P1U41OF1kng7Nj
fH6AnSQzQjachx+8qfF2fCiL2Ra355lyz+a8kMb1rWJUkQiRogJaTPKEqBqyt7V0
/TPlaJItY61xoCT3EdLyZgUk/7Kpn58CkZAvaMIIkYvWAAfGW5ghZxSrwuMdG4eI
ID3G5R1bmZkQYeOPIe9eC59e1vGHsrNNqPOqBRQ+GJPGOWnRQaZ0sxC0/AJx5Tzj
F2nSeH1odnkd1fb+hu7GrCC3njttpfJmpAFYDUkSv/hDQj6j65RUf302iauulUf0
oDpzj3k2pv7PC8TnyQV++B5My+ThIg8tffXzmydi09Bht9cWxKStExyupDiJA/bq
7DHoF6ewK0z7OU5KRSZyJ408qwCk+mQMZp0rJNBH8gpfT8uAeD60HXDIQOTm2PvG
L7lRDE/or4k/+TKAHwJwUQi6iSpplg3U4FfXTN0k10cegLagsCqJj4GF7gFCozAF
txEoRXCTOi+jSrcEcVjGMsAqXwGWv9m8bHt46G2q0pG8Tc/LKgl3vGIDHsFB9m6i
ZxZARIZ/Ez2gs9FDkrBaOR386q4j1R1V1ypYD6MGOJVRsfmlZi2TD8KzpiWvDHAu
a/LgFhpH0pWdkSJV/RYiTOzKPmNoNYcGhBRS4BVlMHBNlwnf9K0lrGJQtXyx+UiM
Oiuyb14ZDrGXWtq1RSyuT9uBa5ikyGqKeGpru4aTDi+yd4R3HW8TkIZrVV/WU82o
uizVikpzryyhc7UiXyQD8nfsMzOgdLeQilAOBPvkJkowQbW5ULzVDBtDr1qLGtVp
VW2FmDxfoXIAQSoKhJzpv/Il1me9xkRbQKLYCan8PDVCE0WFqu9KZeLjmVYjTHXn
GohzgsSwXqggoCMEAI4zjlq/fkj9XJQHaJjaTu6bVscvnlMvk0SK3F3HOwrl9JAN
e6RpG+0hZG3R5NnzJkB8p91ZqpXf7eGaMXoIuAkKRCh/Zunec9IVIHeaV0K69lj+
GGHQnm8NZoogkmGsrJ2KpwaC0ANg716WvnHErSbvps1/aX+vbSyi5fnGLKU9jQR/
krTO+ffnvHFGXF3yA8jDByVezXyRs9IR5ai3RhdAlQoiQa3Iiq7tioY3umTTteqx
G88ff/4tG4yJruHldGlG3Bkd2rRqXUW0N4jy6RJlpqMhmN82m1hrd+yi2Ic6/JmB
5U8cLxu6NFqMYWHV5OLS0rv3IKHmk+120Li7rBjK150RUxfT27oyi01xnJy5mxfp
idGDyq52dkmtAg6dxavUyxtBKQA0b+E7+ej2jyQ0kQAxywXRuG/WCq+ftVAXE9CZ
1APaTj63+Q2om6GAAE0Lp5z14T4A+7a8Rc8oPtp7C/5RdEHocJzfRFvBgxx1Tu2d
gU+HJktFirYP7QiP0kRA5/R/f1NYIynDQz9AIAHZH4GcGgkmIS6D2B6HGE7iUC4c
IcSZW6z/7Xh/W5isWkM5qwGsZ1+DzibGCndHjY0PDqr3PMZMCE+n0YRg0AWUCr5f
o98EFr4fvSAsJng4GgePOJsKmJ6SSFZEqKMDySWCKqqLwfG7bHC70c1w7ztbf8yd
NrrqGqCCj93QmOVDIjkrvZbbgTz1eNIL1hjnTCCSsfRjS+N6+kW7cC0aI7G7OC9Z
f/MNOwo1ZPlQPKzG5k3jvBLFd6hDwFks76+HchuU+bPyDrg1qdENk7paSWed+GxE
Lux4euHugE9ibiWDZZHB0UYFROtVpLPFzgbYqDJhsD1Y23KfYvS0Ea3KvR74y5Yo
LXylQecXbfrW945hMwPYUaApQCX1hc3MLecPLi2mN9dsTKa1sQiZmMnDbUiIS1GA
idoAXlSn/Bj4bjt/USTvzh/4BXjXSzT8aLbfHuHIlLrrWGSwtHQ05p/uaZ7gm1mI
2GOhsmAFqTvX3oprtHqgBcHQRCxwEqp2nsvkTcujfBDsjHFQ6bMvRbA4Zm61r/U2
Zs/MnL//Rye1fFDoV6Eo4dLQYWRp0aGp3sRF9G3HguOYgi5BwdXoNvqnXb91epaY
HWJS0kbVJ7sghf7y5PLUrO89eXHLHZrHEVYJ0WIjfG3+lZWJo5HJj2IbrogL+2Wh
t3t0FPNBUYaEVa9jDQpIY30m6PtoSkHRXDkNpuqIPxSlYJbYsEDUw8akRcVxUyNp
HN/yhgCVqxvtTFz7l5BkOAjD4Rrxh/p51mFDPmpcAth5pTrZSb0644rgtsR/j9yS
8gDqOO9/77oWfDLCiNoEDUg4s3jlXlfveU6BdJ9Vj1VKTgxnb00Kn6LzrLJf7OtH
yL35Ud4nVu2UwGVXYX0lpYPdqXmPWaFZliN2S9hW7hjL4sudNED2YAWl+mzPZWRH
Smq7k/0ySaqwNnF0QYJkgIl6W2FPEy9vs3awNuNpsgLwBfx5YW86QouUOjuhw+O9
kwprM9HyDq+BE8E3VORR7ntvL9/x3Vmm8lFzphZvR3rAAqHI8ZLeP4GnYVTvigqj
K9lypdeLTlDeiu1JppFfpT0eNAfUxhFFmOD6u5fkUsbkj28JfpFBh6aL/O3d218a
PynSMgqplqM2YuTPEQ3OpAbYKzDeP762tuZKSHCWxzACWmPsJ22TuoL5piSC41yK
m5GDTeP9cZxiUbxl+Rw5QEoDZE6+V8bAHOluz242HAXUi+eW0df2IrJ8TJC2zE8z
nCBMzNE9ufWFRiqWEYJwCYe9khUdtr3FzOxtNr41E7qi3cDvFbfY1u18XhAWtMl+
oyrjcHrv2mSqD9sTD3zOJOUGAe2DSOCg08Vl5dXVwqjq4EtICTSOWiJebREAoGjd
DrkEzpvT8W5HMZ4zPaBLuwr52xggXGyDnpunSrP3wip5tOW4EncBVuLJ90dRX7Uh
0slj0G9KZHqNnvBTEB8WfaxNt+/j8ljLZTWm5C60gAqPhwAVsWz0pSCxEYPDJYwO
yT2E9GeAyf0yIszyk392VUPcrUehhjBYH1KmRoNa+Ma1gVYg6C+2P27iP+WghzY9
eE3yhVL0iUg+Tx09JCi09/0Xs72VVeJ4InBuj83ZyJIJwtaLKDJjR0wC0nEpjqpN
hBktBNV3/hZYjg/a3mT/Zx4cuRgFvGm82uBwQR9/h5rYRSyfQQF5Vk4voCSuLlC3
lFjOc0hme03WgJRwOG7evBi1HT/oVm9E/wzmuuhciLJ+HWrQQY3rJi48X5NdQ0Nz
l3iwau30Uvc1DCz9cWNdQd1tuK7dPr5qi37PM2j1/kSPvJEYEyfTyWrKWM6BZl00
lg85/mOFtYiXXMMUbDubCi0WtT8Wzrd0oLCAHQNCVI9FcmLpAeEbkzlRTHcwjlkg
Pn746rQ9CPuUYk+5DWyG9GkMBuNuK0ewVx0YCoLWDcCKeuwNHo/e5rm+w58oqUcE
IGtEhGxu9i/SXaHCpfGq9KBb5694hMHIWQdATiQPAl+u8U13oUX//8ksgjmTNoab
fvyCFaeJdjWXk4yAJqVkYxvE+Vp2HgNWNcKkXQUHuTIXGsD8lWvy941pTKCeIuBK
PvVDmF2ZHXe/6WmTSwo7n7jrE+VohXmacFhX+Z4SVzaLCLhRLqqcTd5jC2bwEzNs
UbAkfGXC0XEiBiaQney3FijHIkw3ewHUkDhc721pK7VG59HkwiWm3ohNpMhroGxQ
jgFEdqQE5FANHTv6mvDGdh8c51GGXRZIKsBDegxgpWwdYQIghYs6p1m66i9m2UE9
Di7mehVv2GwrCJuTYL7CW/DhzhBSfUAGiTapY0M7ghQ2yIl1k3fXT1MJrsbfDO5Y
`pragma protect end_protected
