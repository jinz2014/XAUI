// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mEiBusjySmxIxWWO3VPxWxvwbdJrowRCGBrD4doIFV+jJLE9HXu2jrte8M554X4F
Ev2u7iTjIN4FiXBsoWBlgu4WNzwtvryjvp1WIL3am2PLSje1xSnIl87rHrmut/LJ
ZO4EHq8poddjjrOLAy5va7QQliUkDEelkNr8GVj8v6w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9120)
TDp37PQpbEVfGkfbTpUmGvA2+Budfd5b41rLGPda68IKX6fHqwOIZ7LbkKqb3G2/
UaZVM7gJwRwowRKNz/alcjNuwvK8xKP4QLbFSn3NCQGdzCNNpXFiLJGNFojiNnkV
JWedmFZWPaYp1Ca9ELwu4hkSoeFIZaazcV6wNryG4OOroZU0xJ3mCxNrsjdPMbJY
SN1SDTJnJhE44DvR6uFJV/np/I67aktW2R8SNv61ZIj4SAXz+SmmEanDqsPlUnnP
GBHgFN+KX7zvdWEKrsOFrY7weNfVTfc8DgEYwSre3dyiSkwnwoaCN4LqX93htrEh
22eUiSZp8UzEqu7O/mAJG593k5xDCo0p5BnF3hudwEXPUjQeuJPe64cNqT19KoxQ
rqPyoves4zoXfgGprhtTuAuotPYoM2g6BWSu76/aDVM2ad551r9MBL+oeTNuHHbp
J52cBgqvg4LEQxQ7O+Oet6j10g5EmUotQ4ofgB2g7RdKcyA1PP97LuAIKo0nsAwm
+5yR8Hga7t+6s/NMwjRH3kiF6DpUmfzKVYX3bFzWN63ltPeyV5dXSUH6Mgyvs4LJ
xGBlNbhqPLz1E1vYhk2ViWzCx2VSofenLFnzyoGCeA5fHtuppohFFcyP5Aq0E9Af
SpgbtSPtshZRlecCIdkUmjJvraE7U56Tk1Zylad5JPbBdGFkFiTkV9bU9vLFXeJE
n5wxHSD8qKUb/BqVYYicl1r93c2k0rnxDkfH+USlG1qfZz9Ux16GhARhk1Hu90kC
ODC/mbd0Y7PHhPVUP6v+RATAbgS07RyB3kvIQpj7KaOMkn3l2bymyB4Glu8mRL2T
FX2I0CjVtZuS9esawCmySGpA9ia+6Uvv5oC2zMPEQq/BjvWEv+23/PPEs5q9K8RY
hkS1JUqBvbzjmzcZER2TJ0gRI0YErj59Vl6cXFXsu5Uigo+jbbBxqq6iGPKp3cuY
ZlHDBWMiHTq/DcHoFokwpyX+JwiqQbKWAP0v+3zY25aqVx/5CNICMabDZnCdvdqE
+bmRMEZcE3UXLKxETAShPHMFgDmlQpOFlirCB0HG8ovpohwXvu3agKmrEKOkvcBu
hefsfiypUX2xLOCXNfgVC3U/R82N/QvfUqGLkFNlrYnyBRvXX702j61UKXIphhfP
mhXZe/Kivk8DlHzNAbmSeCemhKJK5Br7lJEsEmEgeXuDnDjln2gikMyj+Bdg0fQb
Q5+PxFLkoDo5k5iBOsPb8LY5EYT3V51cF9NyPpFIyt3YQKyFkIul+eLHxMzdhwS/
a50ClpcdAN/qXntmoK8re0uw0CItgRfG6k7byTxqtjqmozzbgffT0e2jNQ/sIfOv
96MtSpvH+7hU5v/D39992D4R1F8b3Qn3C9HchmmXFaachgasSh9MI6+cM1hzeFoq
/nCZ8Ds9brn+Gbu3cO0teZRff4VDaSLbJBjI6vX121Ed/SgdRhEkFjei77Kt9yaE
km3egYOmt/wbLusJyuEcCbH5BHB1pqpDDba1+ViEKuMvErrx8f7NWayATGm9rBQj
G7y98A4ZPifkVZ9WO1t7DxUshwSSvYP9VS5V/LS2o3w6gOL8k7KZb2hCELUVuMUF
bkEgAbum8CskYkVUJDdzUUFzXd/4raa5YQGi6jFO8dFS6A4rT7r8/Oc3igtLN8Qq
uc3w8Yy32T12RhxFKblHtf2ZQhEZBMj59YoVdKD8xbGqBpqAmppeH/IpTX98GjDN
SWPAFYNAkZzPx2a7qcM65ZUPdg/uX3bHKsF+XN4E74QwXExJMgJngkXl2cPJUmjH
sa8+GWZhyumv1GThHNn55aBH6GxUrOoAhrqbdzVevqEGWo95kKmUMXi3jjHUsGuo
kqcf7+ZfCzQA0KVSx1bUO5HUZmg6t60jBz2e14DKFGcOhTDQr3YuCubQDwqJg+WG
jmAfjnXcx3EeWuG0+YX4yxSm3KP1NS1PBLz8ImoBAddhPgapQgXh/z1DLHyf38eo
NaySeQDII8U+1JcixDTJyJL5lS/TjUaVi6IG47MwlZkN7W1gd2JJhe26YBhoRktI
WhI6+tDCKYDzXlBL34Xu0/ebUgCl8yTskCor1qzbxsgXrl1X4dCph2pCWx5lxZee
blNkhYZsu1UeP+fkFzjfHLa3f15jjvBemsvCvwbXCwio+kfpx00hvlo7vblebKrs
3csj6nmFdspcwYO78dnXs2NdXnxIG7hy0Toc5Elt90LUJWNmYHHybU38Af9aeZiI
Iy8s+ecYo5abXymWZZma9fAe6I9/B5F67L38zyjrGO5p8eNYmdytlzSqRcSZsoFE
Uj92EOgers0IaLejL4iNQfXAqoUoT3xnFbkbwGFvy1HgmSZQ3Jm6QQrFdrqUoVT2
TIDSwZPpO5sQS53ITs/qNmUihdMFceUrMHcBmLttR3g5cSFmNBmjJ/aWHYnA33Uq
zHeRw+aHVeB4VqPQTyJno8UIukc4EhBgYF0JgIJuQoiPaz48RKb4OcR0Lelv+Imd
BElA1mJumTwVoHw4kUeJL2X8JUawM4bZVICbopHGq+vFhIRoa69FU2eXXR46qFvP
ooWqlke7+QMHPNR4Va3MD/z/vvBHiMAeacuTYpxOO0x/ziwJoHnIsKtqt8at7jht
NI7CjMF60woMY81cZsr3ChNGIKmX2bBqNp7A+LBTFmaYhqr7zLTJ0wMQu6bPS5z/
SF8QDiaHYec5HEucYXspnSku0qrpZG918DYSpTUzPAddSAuF42xnQDLwTZlbt/22
9fStCJ/I4eZ23afrTyVc8CnfgB5/o3CfqusU4+fTZ1WdNPJPEwrj55uB9YLI5joA
s9lNyLq8eqQz0CaQxzphc76iF8slXvPaDPYw1I60wUlkt45dELqbIU2qEkenxQ7n
dJpFnHRj+irzf5vuQhoWiZGIWVy1wpQTaWft9F/W9MPFBuc1h3Gv2RASl+tTfBUJ
BLZEQmkfSwXyiL/A53tIU1vwuh2fFOzRGg5nrXpiTUXZDF6aC/z35BDxLl47nb7h
kA9h8SQcOnp30/RO+u9ABUD/w34Lo/FtjBhi3r3nJhQetuhbfiUm+RqVmiBmW/lg
h3LRfjGZy+DMnDEBGZnHGYXtBGILSh/0s1RLca/MJ7pwuAxle1fneCm/TxmCuOa3
BzLKJRVi5l2gzGdxf/eaChx++ov1XVrbL7EauhAogYELt/V1/P9BeqHGGGnE2eES
kLedtQEQm2m2XUQH6sistBMtJTBrjWBFZX9/ltj3UFSy1U044XwPMKQYfbPJk7NT
AOBuYuoN/CAqnY6Jk9MEO9Ek6krvzi78Fxl4oiH2M1abXdSnZGz62H0IN/9kJoko
SLI3k+hLs8GPZui4RrjWosXyDwbrwGZJPE39/N5pZatqjkfYzXiSWecq9oo6y/c7
FxSj7ZMrA0yo+ZtMs5iTpBPabIiHFyLy7z9YBj8PN63mifSEG1d7ipunMgMMVug3
CZAZDFi7F3+VFhvGWclBAApLFmLasIKiJ1IYFGfUPoyKJARlc7++J/PajFbxfQo7
A5TWqSSJS+x6lVRoRmGxFfW8hPrBxwjG9UbAzhp3cDSxRDVzKtKQmEIRiddJr2Ea
zXhvGwAZEO5o9VO5vHiTncC08xQKFsEl2eK2GxRuGKNQnpFu+/ZkwlaVTHcx4l4/
otyCZ3x/odptTIRX3G5QxR3aSRH5xXlR4oQiDQnNudSPklIOmqJ+OkN9ybIkfgwH
QyDsYKH5tgcdbvm4Kkbfn3I6Gu2nSa+RK5ZgPtkupMLqUmADMQ5ReVcOn4CpjHTK
E2gNS37WkesKNnj9mySMdK2Pj1UPgWC7ZEGi1fmMkmNGTEnYGAJXRMFU4TDN0OlE
gm2Dyg8R92VGcwWG5eMOpOm6ibHinBmGih0iq4bcFEHTyXxWMY+GGDIXe8b9Fm/d
HCWVGNGqiXK8BJpTMydRVVVtfpMDOxFb+9dXUo5P8yI3I9IOiPU8mSwdjz8waoKS
PG+5a26bsUqJs5QyyvjXhuPwLmpYF0Sh1wMmDepRL0UrBeJZuSNdcfjqTZzyt35i
LXN5kqr7vgn9ayjpQz/h21EPuPxkatD8YyhymdGTVx/NYw0Zgc4kt1qdxofOc2Nw
sIFwgcHsdAOKkLad5JXt+NiMXkM0xxILgAeNXQRosbp+eXqLyIW2QkdCXR7rUz0V
5oDgEIe7teNyakA5dXLgy/60Czcwfr4Z7xaiPGiW6fdtdkseD5RXXtZhgW8OqA2C
gyGgehF2Vq3rI14rGo0YgeA3ukHLrsI0ip019ygfvg+oXk0QXHevC5m511N7tC4P
r+nXS9oIdKE8sQMFZfJuPE720bzAH20DDZGX/IokZj1Mdv8ZdWQMczeVP8Ka1dkH
3MSqZR2JCiXPKl0QmQeR1I9Abbpbay2x19zy68cCNCWjti7ej/iM9HADv05MyKM3
IEqNWJHPez+TWgt6uUbMye2RsjEYundihZ7junBAj6bu+UKZUr6y1iBwM6Tlfn3N
zc/VspoWss5WkATie/INXJXObCXwehQPH0sKPmCwag4ljio+oRBnDOTKylHDOsqi
I/KNY6tWaLJ++ZPqLYDoiX8rCzhruh6ZQnuGU2H5KRA/9w360Azxzp3V9hCPEjpC
Y2o3usnovc07X4rYW3XJPwvhVTJ1QULAI8txVkl9sPntBSZcJP0Ps4GyKFMY23E5
ICXfEaHVZYCe4yD08itKQosTCRFECzGLbc0gOdH2fXI/5g8uzC2UbemIfj8KeYNy
pDoKG8DQde1QQ+VoUcPUapU/6ksOdQMgIC/eD0wQTDdUKCcX2ke2xnbzDHPeAclC
cu6gtV8OfUk5nHoYeN9p9+0eTk6j7G2TF9ext+PtNk8UANHZAU/4ifABNZN+tjGv
WTmMc0L6omvRawiFzao+mqfuw3cSuDXL+WmQOr4Wc0F+/Rt/Rx0F1nvmUwxP4/YD
+4Mf2xRZh1E1WPtCecg+tx1q5p83lH2ZspoMVC5U330SXh9J7tgMudzLkcXIw3Vi
xvYk/XUZ49CAoVxdNplt/0GEOZtlv2FH5Tv1RmHFPxR+C4+8zdfTk3bCo7ZpoxtY
nda4bpoRlcxgmId1lsfZSMrN4Io9Q4XQG84AtS0NhjMd2AQ2UvJZQczlfXBK9ROF
VlK4mSJdaj4dXaOhpBgxZG6nR1eWe4IaJEkqo79tZ/t4+VdSAUKWDUEQKEYwdSff
wkh5DKLL4C9N98bIbVKgJFMzf4ZTaZPGNZ+2fDPnI1/Vufbh0aJfWXL843FliaFP
jjrTkO1P1jVm+uDTyUaxU286UB4LNyfZAqgSEK04o697Iv6VXA4FOx87G1VIZ/Q4
OuKGl9GORq2Ksc1NMH9tYV0+BwWre4JXS3PU9nx9VpFKkA04ydF9y9DhYi6Vd/ae
P6TL0Gf37EpOSgNwCySENYGhJFUJKfMThbRrt/Kb89qS3dU7CClj106ELSFOY9rJ
2QYil6p9pMLvItfjQ7JuXOdRCk29PKJUNsvjgDLAjOUmp/QVk+e09pDVdjCW5laf
rCLMBywb0FunuoPt1unV6Ie0S8ZSgEXPcUPlzCVX1RSfx4efEv6Prqc9JRXQZrCQ
ZLN5T1QbbrN1a37dc0fxzyvTLznAqMnWTWZWxizRyg4S0PECWN4aD1UxDn4aDmW9
zWUcbXQb4vWYCjCr7B/DRUBvcQj0pkHQkAtc0q2OF/o5pvCPXABpR5RAusOdVzZp
Qy1aKMmApwYGvlXJxKc4jEizJDpZynp89CZQ3ZDemRsFdyJ3Wo5WeeSSwSB0YL8z
FlsmU6aYeDM3Err/hM8Pinr6AhD40m2s4INwPYUTiRHd9kkdSWgEUxcREMLyESaf
fBT7rlxN/Tpx87O75VEkWno0H8yP8ivHy7JeN1jXyGc/lOu0Zq+LVIf3f0QIVYa8
E5i99owGEPX3v6veLUxF1adVtjWbQ1RC94Z7OghL3gSEf5JLYDhSL1lpPsmH+wHe
yBSQPEz8K2rKhIYDh9IQFMRC5l6eX8HGxSDFxDW5nqOBSgpQ1MeuRiSBwXDA19tD
F8u5fyG9tx8SUwTN1+IQPBPac4nBEJ9CvJkIb5NALR0TohFqGIq3mlp1rxtWHoU2
MtR8i54iHuEl0PVvLSpkFepD6DmD2JuO+p1KZfyxPtqaEnXadkharzZa1KuHvtrE
7o5zoory4Us1RQdBvKFgFCcQ68AYYwZOFiuvVDNVHAWB/FvQEYO4jLPAG2qqARMO
8VDSWu/F3/UdpcGk+ReILADDtpQ5msoNih6dRCrAs3t4yle+yHR6fxsIhR6NwPSY
S+OwOFOBFeyVbtyRsqfrG8Bo08tvDRoLe0dbWSJopvvO+ANXxAUmCHP9snYiUDsL
Y5XCNh90PA/3gP/uluLiy63LWzCHLb+5zRr2bEvgptQyiNM4uBIP4xvbGzOQdBoA
3le/8c0k9id3JHOKivwdYKgwzaO72Yb6IYHT9ufSs31P1je+35JMSf9VsG1bgq5l
03JcwG8+W+BoBM6SIBUsasuGhSLOWUaDtvJyN0xOD13Bd6XfcKZsczFYc0ikAbg9
7Ya292pL/mEnG2XZ7eDARMGIZp7A/KaISNUCLry2I0Q2TLVhSq9VYirCe0GMzp7m
bf2TG/kIcUoriPY7CunR7DEtZalYFka9Ww+hlbaOpv/I47zIf4A4334n3T9oENRj
Gas0qINak/X+FScVAbED7YhcpOhP1Z1slHI/nFS60+gMwa0SYtPe4QJddJIhqC1/
7DbPhi/N+vtlmB0Ts8HimU7ZidxCoOXMzCinLDS0uoKJN9gI8nmeCkBYc10kf4lZ
FcAKbthSzYTB9GsmV0VCDywBheDa6kfJhh0at4kdsbicqiejE6b+j9aiP3ek14cb
4e5wvmtSbGdGSTK7sOOl+k5rN/n4lAq140afOsN1NQFZUX2okBeQtlJ4S5lXWPyN
cp6FWiWopEE87M8/j7Muq/i+c03fkrlzxA20DmZJjPvf1iB0Ve8nuPrBNGNi6XHH
AHvYFdVdDBZO5Ecua/e5OVwV0I7H/RoHDGJeCb8f1cxnA7vJvJ3qmq3MIf71Oww1
yn0gMy0ksbjj5WO+llFf4mJ0IRHzcIBd+ziuddAaJvn2DZJY4fQz0u8Q04tBXy3c
RKgDNSGICwp+KpeHsfYj3kjZ1SfhHIWhzcB64Cn2Y+BWnlRJsGhix9Bg0Nxvou38
4rvYA5852M77wwoRCb88BU+GAjexxmfxzGgLo7cK++3+B/NCgFNOKHQpkUHjus2Y
KCXKx8FDylyhguMsEqG+90ZiyZl1H2vwvTBmGtxHRJXz4otb87gj7LHqKwhj0Wq7
GmdfK8bzo7PXFLzlJgLPY/zfXKyCNt3iD5il6yugC/9VpzqgshTmsJAb/UR++CcK
fWC9dOXiSpQsgUEO6ob72yWr72CBPsVHjHLnNfymfxr/K2rO2mfIPYQ2AAgE2a3n
c8eNJ/f6VLHQaHrWzDFVnMqvYTRd69ylJGsvCovJ99F2k2+Z6PZ/zj8u3ezJ4R94
YMBOu+uubk1rx7srUWdBH0bVINro7xHbg0x5UKMSmfljXIFTK+esK7QA/vQjzRJd
uJCa9bEb9LrJINaJIBF4y8Zkf/WR9OsPVzaJ1mZ8OoX5NkZ/KXiew59GHdo8aJ4z
gekAs75Be6iAAZl7Da9UQOgpT7TIAxr+U9Pi+AyNgzsKiZcFdabBehKUD5hpD4DW
cl7MaBO1yRux6c4bvv23lGlYIyj8q/qxprHFA+l6I0+QEiZamCIWCIcxZiFGOaDc
DbQzvC/w48KgQXmrSst6q7dg3zM6H32vCSBZBBK6i2IrubsQoJWO6XCbqKSMBzO2
mZWF9zfSb17VHWKT+Y3TK6p1Wl25TlBTXsG/IBNEJQSkh15W3iL185t8TfCUhY6J
1/So8zhkAq+d4dzB/6Zuzt+0E40xiE2OzC0kJcu25EqCvw5CdYeqUfU7me9Po/Dx
akWz7x/zwZA+4uVKqAuR26kEKIdNIG2T0LP7qv3LwJDj6OwHatGanEcJAtoIjCqR
mEO2gm6isW7GtXHkLC7B5eg2/zEqCEoSsc0NdSwJOT7PoEl3XkISKn7cVYtXyfmn
wGPFktC7m/4OySe2vaON9keXiTdxiOJNTNIFFVybqQ9IuTHC02spuCf8KjMJXWXq
5uq+CBu5F9BNHf4xs9pP3WU/fJB4a4zpDTTQaB8WNpTop1kSHw/1wDjaCoJHp3lr
v42pPIwyONhlxbIahpA+Ibi+bFuI1IRep0tC0/Ct8pnISCzLEnrfUWNxiHhj8p43
nSjgmSorLgyXRf6qu3YPnaQ4PQdnYsCstlN9CnUHmpEbT1H/P+T0QhTywf92bA8m
bxidaBdD6elDR18gx9TDTs4RmibXRcX38TG5JUr6M3mpQDIjfyqKcKX3RyOGLBSP
OChSDCfWqL5hQ1uxAlLiYKLV2UnNFXWO8q7VEsiYf6TXR864kAWimtt/R0YZ3BAT
21U1kTzxTbgcHPqqtoWIKANOw+WKmg2Mywe8rWOIG90eW25xfodkeTbrA3omiymc
5Qt9BPjyr9030ecLscsh6kZgZBCbeqURAt4v1MXBig78632PiYadoxOV59AVBNU0
I7Hl0oqafOeuxGe54fVOvVm7Z0PsA7hy4hFXZY12AS53Tz+M57u8Y6ay0eUMN+tV
iWcrvkNSkF2TuGteIqGW11ap/+Z/frxH/xGdZaphE1Xo/6dRRn8HUXx9+eTtvGHj
HwuP3YKdGAzPc7wIthnZQ/hhTRJaO80QB3xkP+uZ9mMWy+3mitRLAUJmi35TBxl/
koTohBLw1qMbLNqiiR1Xzx1+jNDVbex4w/RnflRYw/64y3hCVIv/6CkP5AwBTC+F
7XhaEaCQvy3qV/pc/ffO5JtsJ0v3PXb1WZSiZB4eR+NM3ebr5n8WBDsJnHaTg07K
uJctOgQvPirZPRvZ4BKBb+UjrUfTguJGbhDUxVMwiogj1AcFmyVsX0N16VJKPhL8
cBYsnL7NMJQNyOq8haYOG7tgS5b69T7Se4ZeI/8Os0j0IzfgiVqCI6BA0/D2vTPA
Pb0zMOw68FCQtif49JbCReijNahPZIA06JDGvC2iC1ageZSHDgWbiJsBGw6ZxGDS
Lshtja9Q1/nKBLJj+tBWXBljR2iIcgtcFH643kf7PUSFPof8hF2Hfxzey9LB1CIP
Ekc5jBoKsjQyhSjNHta24iosXwRBnUkI+862060t3CaiOqB5vO/b0y0QdDj/0NWM
lQ+jliTWYzVujVYUvndW4W9AhvVrL0zYJx+Gk3kyuB7O2AETyXddh9hsLTDlsyaE
q1q23qEdbTOTiuO6oPZWqDrSXUZSLA+rCJePdhA7+60Gd3w9pQeFrOfWRaWANM6s
7PtiQWsY2VUPGUAJbwgzcyMdr7WAH9dAUwm8/1xSR47WwqpypWhtsBZJYGEEFR59
1pMDvyzZWav0Vpke9CtiFhjmQl9I0l2p4w9ZCRkWO+7mY53ju/IWPWZfJnfBH6dr
vCf7JQ05Z9nvcPV7eoNDR1IGEo4EsCGpUJLAAESK3Cc9pac6GNjEELWOt3huRoxi
+sEu/AgUgRFauFlG+CQnipo5GxN/Ox6wYyIE6BqSFuHVhymG+6lklDEt+cqBy4UG
n1g/6dkMOspIpjLypisIz2OR3WKYLrBSaNrGZTiNvBeQPPRpx35itlYcBNtO8f5H
K4F4SHLN8guPtT7akPuELsLqu/Mc7lFlYHNmKi0iQ6caCo2fvfpXNbrm9spXcj/k
EHtPxrSIkgFRU4nvlPzNYDuCi36U2h23Z0I6HDZVMCv3k1OJUc05HK6yHpcXnmkV
ejenBUcKIXbA46FwBi4nhsRpnqtpnIJe2LtXS++tbMWG2hPvs6/n8xaY/kdQeyhX
TwVHWKAZwtXBeBAKIMv+1sdl0hokvtQtq54b6lph3szUwLqic3Sfgr1EjUxB1FEN
2HvzDu2yaw6vPLv4h5yzcqYGuPxeZ9p9Pnq0IXnpQj0Gf3PjgLVSIRS3X2JfSTV1
988lmBumpC2vvJZLEyDtmba3rmOmX1WVqbZ149HRSC1EaWXOMsE0N7ubIo4QHeeJ
1aPXe63SaUknSrIhaM5suGzHcmoULJsUFd7ERZy5dc9Js07fFh5kyvkYx0KfK6aw
KBx+f0NyKw3C5LHGU49YRP90rpid1RmV7kAgg6MUr/71iPdmXzkFHJGvKib0bOxO
7PJT9ywE0EQsXlPk1i1QOYpPMgfDNzNZ3z3YzPsbIHj/KLhkFB0hzeB1tajmSGfs
o63DCKkdYnnhb1KiwMpblfBrAEEdMAva2oJ+yaoepB2ywsJtpp9iW4gEUCXF9UcZ
4wxpUAy6MvRArGsa5dB7CQve7N1ZU4aO19sDfD3nnKAkyRJ9IJD3xJ43YGW/JbeF
2iE+aBxnezdmkFzCQBlWUnFAbCfHUibi9B6uWXtuPmTzKGLVbbFViLbKcw8wTmiB
s8cjY1nrf2zaumXYUgzuhhh/VRMVZpy5tZsvU80Tyg4cmkJY4eJm86obQCj+6jt2
06iYnbppImjIoTq57TLAmyIqbaO0F3oFufh5j5VWGWO4NUgqnyIXXTAn5gBjE6ek
LEpxGFYw122VdVZG4T5N2QNxoP+pkb+PtwHX+MOPX99t/nV1ItFVvT3vNBMv485Q
pnCTrbN1fMVDYTQErz2ueW4L1L1lc2271QicPkM5xIMzUvdmAxuWkoFjntWmv7MI
4QmJ7RJ/GPMckT5jNtrPiiy+hCz+BUw4Rs11nShRbwEFWeDieGRYq98T+ovwgq6W
aNjRt4muc1wucAz573BoGityH+pPsJbPWejbH+JLXMMvy+NaN+jy3fqFSOtUTgE6
A/wuQIdugKcI+IO3DG8tWXf71cuarpi1M38thj5mL7Ru8e7BtEqbmWkWmRv+Eb8c
h/hKe/xiLl7/FhO3k+sMNDzJX/K5KihRbAIgg5mc+VcfHNzJMex+miq8yuipl3s8
qiG6a8kz1R1XPYGnZVDuEYBIXq9QWKKNWcAbQJh3ZLnFATzz9Ikwlqh3UP+CVC+b
08/k53hqbQ7abYBN/oux7/FiXqi2F3BRHcFTW+9611QRjdVaW3NY1xBIiexrIJKZ
ZiEr6eZrAthqR2g3bEMW5gaZf61imirKVEKvPaIUzrw43XkUEKpIB6Xn/vMTpdQE
71ZrG4n38zpmTpsJW8MSV+Xt2MJruaTEgVmEO8n7nE8EBrSTL8v7Y0DjmnZHFQZO
wUpu8i07SCUmtuhuPEviAk71tE1nFw/CRbvgCVAXgTb3dURA5chUh4Pf/sUObl8O
bOBiuqdPhbZah4zGRxk6NGEt46uVdLy4OUdvMMyywctmOK3mwS8u/t5h+b/VSG5K
KRNf9thH13oJPoNsD4x8KHMZSYqW9P/0Qq9BoH5pSSxzCSPBwLib16c1jYmKK6ZV
aFkeP66kD0Zg3rSKUwN/9OS/Oug8r8aSZQosaGBDXxQjHkrkEm9FJhatrqmF936c
pTzNAWw8G/OkXjyGvARFKYJD5NWGYJmvKGCvQjg2QuTsCNZ9PIxTLQTPqjTkyvgk
KlhAFWQAUqb5idXj/J16vR/2sIXzmyIZ5LYhifa4NiEgYEZX67bTr55sPhvu+sne
ljB26jczJHJzERDHdDIkB1eKrKG591/gHQT0F7My3+PdEZmDF2tYtMblvmp9LEng
QiodwUmRn234ZdQb0Ip8o8e1Uj4rOUigbOO/WFblmgGtNm1HEEk9VpefL8XL3DRY
9qy0/DMuE6XUv6Nc0EyLbMHU1sisBQrwqi3iEJQF1HXP1KYa45lCKBIlGwm5kJGb
iJ/0IYPcbvnqHD3U9/aEGvBZjBdvTVsMVNvk+KJTz7mSuvCcd+1qU5VaFhny7zfM
1GuyrgpP6iK34ONJGJIsmG6UfIlqyaQko2GOqUrxXaZKU1ODgePKx5rYC4L/mMsm
T/7e8SWsaU4kztc39wuyEZ7MvuWRlsca8nlP/r0+vLurYBVuL4SMnFc6vmgJ4dsk
/aMrEyEGenPqg/zQqdGenBYMet7zzyUk0nvy6vjODKYi1nY+10dKOSzhTGWGG/MO
AtgOpaUt4q7ru11WMhljdoK5ItpDn2BLe2GX3jwWUY89IavpFaOxFbbdNN2VlsiP
hFwPvCGoyFfbqZyjEE5+h1MLENjOjozhlR8iVaHTWMhouc9RJLh7jvu8da1jehnn
`pragma protect end_protected
