// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:31 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UmRbARGjyNs2+WUdCg6ugitR+xTOTAqY5TAuNqqmquLvPPDOZHeD0XHXO+FZAOEc
IlHG3VIwA0zmZMI0HM3HsFs0ABQkl5Oqtc0RbH/3HD7Y6UNi7MqN43+AfxUuPQVz
k9+f4CUQx7UYeBlhR+dmnlYFB7jTpQwh/uH5F0jLcko=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33184)
R/8QXSj+55a71VtQgzdgLg6eoFzXuJ61rEw3ne6KB+EY2mq/XzCqY9TQ/LWHAxEu
iqJ8rSW14N2xt9UemLXjz76xA8rR5wYiXK83R4X+q6iX47uodiZGk5YHix7nysY+
ONHZoFVrQ9BOb5Pv3FlGFFZX7Sf9eOrdT2yXBqhy72XgkdF0FcZtfje15ZKAFymw
gVdOVmgB+QTebXburUY0rMg8MYHZGIcHeYzHER9+wCb8PMB+ZUtpP9zFw1QnOU7C
/qOCl7RhZbh6IqfGsx1BgB8q94VnKPbaV81kgZwWTl5r8r2j3cdeyQOYexb5EWtq
6I2cNwOO7SNH64IB7kAGqR8FHApSkZffnBih34p/e1xLLhMzYKV9W9k2GpmbSbi3
WGaLV91v3oOgCxtgk3+kn4XHGKVMs8mNjJqsvyYYUJYImf6VW3Wd3UM06D4BpIs7
E2pKuovG6cTXfa7A0aae84PmRxE/BbsF5DKDjaLCpuhUzyXEU8i3qjVMLMr13oWl
kWc2ioqVkAHMUSU10m8au1ihSWBn6pZUDO6MlDZSdNESES9NyciU5EHmoQ2iSKyX
xMGQMzZj6Oi48GnXpnX4j6p7di5CFfay4KCx1slSapRCm2M1pB0pkeFQKHh2N+g3
uu6sf2Prp/SwSZ5KDzvSm4wiYNWhPUf00VrP0V+ruD1cjqPZGnPoupaa4lzIMsxJ
UadWkyEHMz4S1PbRqGRZzM32dve16AhrTNAjsgFkpYZ09rFeD2I74D4ePEvSllz2
/po6cfaQlmhGAmXZkXVMcme2inbnJ663LVaI5tgSekAlnAuzBcaqsOmqULifGSi0
0QuxRp4r/RGIUelMGQhSd4dnoP83qNaC8ab/b39wo9iwllcuYbxNiU5CLvZ6fFwo
BkyG3rv67nItWL9tW4VAQA+nCxaOuNFJqyFBAqrzQavEFmuIYwJWpRa2NrK6JhlM
2GSpDGv5Xp73kY6bFxkIapLXQoU2H6pf1BRewbMKLZKc84LUt8ruYj+dH1P/UZJh
3a8nfJzkvORbvfvgci+duXf1L4XkvOR4AgBwHrZ1eu0N2QTE1062KkzkX8BLi7M+
7FxTcocAROxfZqCm8l6ZeT1CRTBQJcquqCM0p7N0A0fATfwCJTLQFE82TkfqtPap
Cv4UGqresw8tYAreJxzWH2KVPmhDjgvnOstREuop6uAve7vdj+OW3WCNFko5mVIR
Uv3C36lJ/fMiA32iyuj+Nk1fxfCzdUrGE4YuwG///b13Zoi0JUK+M51YsXc0J40d
K09dB+jb2LbtoaXTZ6ssV/SThJ17yHAOtkjDQvm3G9jCIEh/TrkSu6EpHpJL2Q4g
/5XJE0Pq8St0JdltSQXb/cb1rqA9Q7f7krL4uJEQ//ZUAKNUg29IdwPqgV1RZU0A
gjsQjW2aC7L2O+9C+a4aamb+ndn/RlsjVmjioZ1skL5BLQGVdg7tk2IBzs9kMKAH
3f/AGa3YdtBk50b+Vq23V4kRnP5we+y63rgj2cE/hPDW1MgdL0SpC2U++u7oEBmQ
4wOatSVrLLeHMcl7wVZrhNK81/a5J6jBkhjQr44LEYlGtdpaGxgNoBWMxUC6NkCz
4VwNKyCQbVtdvKzP5tqf5pZkbt6PLTTWY5UnW+qnqPhecg0kK0LRg/EcAyzIZB1t
xJZ2pCnBMLxRv9rofjXyTbVnt6mrM2Z25Zt/MD010BX/1awJ1sUw64QKcB5oM8/W
sRlxVQGJmac2q1lc0QTv+ZHr3aeUcsRRB158cCkfIeFzS3PEBiEF0NJnW9L7A1BV
2SvJcpUciOJQVPGU+WijY5GW6OHetWhgwBuEJn8sUI/T9djfz3mWIAPFo3PxpB+z
/BR0tJpq8cD4awqVj/TLBsJj1N/vrLZ9VTh7jIrXYpbZuxFi1lgH8gZm6BFHt2Cw
nuZmprU2BccFlVnYwxPKIlhXiV3f3mATqikN8pkclNg6Y6k1K03lQFQNioWj7Pkp
GdiKmzP4bz5N2nG3q+2MgwA26ksCCKAakkOlwn+VVu6r2CbXLSJi5KYn1xM8niIQ
cEdkqVc/gCgVXY3aBBAY6uQOiwb8Dbyynxf84z2FiH5H3senleiburpsct54qGkj
u6hf4nGvu2hhCLGjEMYrYk4taT1gNWhLo/idhJlKlvqb7BQHDcGWUpV5k2fmzD0j
Yqtcmk1dU6Bx32ziFD/NdQJ2BrIRZAvgR5gmF+33WcNKnbevaTM1z/Uga7QmR4MU
A1PiTWhsiDD5nwvxuco9hkIR0Z6kDVnAKduLum8lfND2HCrbfdVNpjwDu1UZalLM
sUc5nBkxOQz2gk8+k4u1vRIhZyRuHBNHDI7FdEFl6oFrpfzjSmrRPpUmT3iNzLTH
V2/242XLOIpObyTWq8bSYfTOeG05FFtO1lBgwnXkg3l/Q/KqwIIHdSUrrVbLjZFJ
QBTy3SfjLpZjvv0nAv6+a91DDkXmZ6VaOI+aBAh3VM8eiMXeabBwaW6o1hSy1qF6
tcDQV09JWUmmvKzMjLqYLafoX4YTRcIbftJR/ag/5g0NVw3mMq/va6pmeZG7RQcd
AWHBTDwlqbADUF5t1AHIluO5FUUpZZ9cTs8iPFd9qQjkUmYtiPk2x3t0e74hbC5G
SpwQcKLQS2c5ac0/r7NZeOCw2p7SsfjCzG6QKW0jjKBJotZOnli1qIGl64UXkSLN
eLud9yisYCf4Id83KAcMFLzYBV91JcbwKAGeK3QHkxA666BpZAJznYZKOb3zy5o0
D6lGtDidep9hqtESx9M9lKjQY6IQZ/nhjrCYyGlhM25s/ku9NO2lWWx/bSAYJhjb
C7hZj5vLyusn5r1PXU+x5gG7Bpp4orQsSvLpkDuhbot/x9VisePJRzCcxX7Ejjme
p2Wc0eVmnXiEnPSytew6VHXPL9b/Z2NuW+3hsWBmp8bfmbPlVefgFp9oPDp3WhYo
WdPDl79DWrb1odnxclk6TJXkA25QMtqoNGK4nToCKsLWhc/oooDboGQJcmW7D5KT
x2XcF6fwo9XFdQ/1HYfljDBiCRVLh5WF0pJhSY82+AZNOY2MWxbRzt38IrqKwWAX
9+je+mOskFaBNOAEk2CStj97QWqKYMNPcuchk1NemOEcjTlEKCj4tvhUDec0bJgF
fySZv/1dMK8Cg8rnr9Nr0xFggkwvU+nAAAoAdzCB26wifXXr0kMVrx7P5wDzd9I2
ClS4kqUqaJlPlXb1PCWv8oS5cz3VAfLEr2zqJTA4DyJQOukOictfkVndkuDWyq7N
ijrDc4wX2967sgPOSGkwlZ9YIHYXMq6AHIGjKWueM4jkwCD/aFlsrnWOyCUSMXg6
6dXl/ot7ZwFlpjwWpBl+0JAqNylgFQKrCk8yRTMkF3nxhwXd73ZykaDg13WF7ETa
vAR/9hdz3xAV2YEd4iz4JTPIBX0EedmjHyqzwQbHZTHxenOyNwx/rMN/rVMBxQnR
yhLrAm2/n3WSf5iMoeAbROn60RFJOk113I3sGawGl3IH1wgzIj1p6i188LTM/R67
nunI2cQdXgMkGtoQOAXUcCw4AF4/Eg5NoswjOjGAQMfAlKPSbBJ8OkHhG0orpmw8
KzxjLpoY8WAfru56GwLFogUCgBxbcCDd3enEis0SW2tF3Lgk0GVJXyfiMGu1C4bc
KItjjYBdqYh35Rh2UuJHurPsFY92IhlZGOVRuPrYtsRol5o/Vne74z0EH0ky4Lq0
GcJ3B/K+xmt0swStGBfX5ya3k6hLcv7YDd/+qMYiwTbagIJKh2srup5LTd3TXHxN
gCrmK7W8LewBhVhZYlZLDLD4lXKB21f2i79IHqgflw2vmc6itrDMciCWMtcp6b8E
KvT01k8HWfad2W+LbJFxAdYwmSzt+OeG90f8QfY0Gc952N2/EacFVS6LbKLFq2yq
WVcLT0ilRByClBplc83QQoo0s5769Ul7sceL7QkOMrWp0FehVvbCi1dgZTLPX830
kD7HtEeDOt04lI/MCx0QrIBv5UlSRShC9d7zivNEUTTUJEjJunlU/eT24LUCDPFf
lMfmQXM38d4cUk/jWACrw0WMkK7LOyIxYqjQRe9+0VeV2Sb9NFLxzi+/bw9nYBOQ
FvMMhDqdvVxISvP8j9/VVOf8Gag1FVihahNRjIGNlBUmx+WDFOyaD8F6W/geHehW
gguBDnedMHcmTfM4ihhjqSWuOiNcOCG7buSu5eB5+BZXcxr3MXdR89BIRfSKL7lm
CeimZK8u4+y/WGASz3EyHQ77ayj7J+MPPtX7SCp5H9dsdy66rf80mdUt9bb1qOz8
NWYRyx4h1PIqL3N7M63X2K08AKkVW5Hm7OJ5oDZafCs/nkUwPoL/5tkcmy3fxVTP
Icofw7QO/q1SeQM77osTbM9Xzsxt8OP4he5M/bn8rh9SSyo+9EnnDdTgDqf1e/qN
NTATf5iyMWt8UisAekGg+gNgvtBKGdxCdQImkoggtGpJw3ZfgoqIEHN9nGhbnERH
PgmIErRKIunvzYZlyVmOCvPigILPcCdiv3hrvzdG/8z5HA69OkspZBcY9KpykHp9
uOEBB+Fj3DPYyIC/JoCm17ZN9oJGRmkdVOzz11iB7OaQeoOHdaO2yQDsi4op+7Yg
kJenu0H3nOF8p2uOfnsd3UoEATJmirdQL24oXG+cQy0KlUctjqO0+G9eZUSMI6pr
UyU/7epSCIVFZmt4tH1Pcox2XWO4K+CiRtW3Iwrwb9a4FWEaagcep0HoW1IZtagB
ljw4EJlp4uUkqSs7Z/+wX/xB/kWB5NEDlp4LlUYFgKhJaAec7oogsPkSV8wr5Nxm
FHAvcFAMi49ugpm8W/w0SZBPgQ94+7qzAR2oq+FEthLXrHThxvY9tuGKEkL1FLk5
DzZMy+hFtIAwo2Zo5PWqmNO5XN5cv3FUGe/2P95ZP8m4Yrq6rWUPfPbvA59PSlKy
CWQ/Uweyw8N6L7GPTRjLqEhJUMEtDQmYNbiFh36/ZqdsRgodf3HQV8c8tnwWC8M6
A9+vBRXDDUFU6Ec+nwLLwtYU7sWGsIOXfh8fE9Kk0Et5DZY83RcYvAwqZ1xczJCX
HY1nWNlrd8jRalWVBpxV42aZflSCNzjMLGPJtbPmXX4jXtoGOJRX3LhsJMAUW9u1
RLCLTYiBqQpqKCjdoVMbC3zc8oKmoeNcjoDkzFB2O/8OHahmKwqWOoJHRm3Q1KAQ
3sNq5b5hwoYKb3mwpx07D2o5sSkbk72JoDSOPApiXAWC5BPK/KGUwujWMHOoLJpK
Ifu+X/N1sqboh67M4g5qCiui8Tq1U+Ijrxf8LstEokU6Anf+qb66LP8H69wvLshD
n7OfnVXFz0VLbf6veUNk8Qrlz4Ok1703MeyHQR/qgQvlV7K+iDp0dSxEibhjxSZq
VdkLbAbYEyAmKrpiqPruEUmMyxBT7vlOMh76sBHc/VqzFfHeVRdfhiuoinecydER
dU5OtPPTh82JNSqFd1qZEZ/ihA73vT79d0BMq+SyMrMFLN1QUqNz4Jm0hhLX94vc
a4WfttjLSezA/hzak2Sc4hR0xbtERwCFng7sjECGm9m9AXrdo2PW9pykOCFvDiHC
ONY+/bymDOvY1XNgpZn+6emifGWBna46ZSO4Z2fGdxju7SXewxdmvViVt9r4i5Rl
0tYZMZtBtNyMPESNUgQirYrP93z2F1a+N0ASu8n0d/TYYekUGuPzBVFxubbd6h2C
On7LzhMRSR3dzRYna3qryKYAlLHbNKnxLwHzPaBb2F+/nhxZJWxVjzpWnHB9amcb
kdrHB3ErLVKvIDn6b782zWEgHO6OR8jeEPMeHZmdsfe4DkTGPzcNeNL7TQCaN0pR
VPfmBX+/T/AOvq7NvQwl5TvSHg7cFpMl4OlMCqY7weM4MQ89Egp20yOHffPJDxgP
/v30XFtp2iKx1OBpsYVrwPSI7Cp5OoIo6fZMWL69bGmcNd++o1y1JvC8rVP6Jtup
1VdDRawaFsRc1G2XNqJe7KlDKqrq3dNRwYSg5mrTuyLpyL+g6xLxvO7gjho9kBxE
fT/VOapxJa0oVCatuvJn09shB8RWyzsMCgqz6QfAGA0mhIsbz2fWR7PrpahL0ctb
ire/q3ZQl40U8+GcQfT9VyOseiL9qYxmXnvGS09xLctk5vFl2fjVUcZwdNmoeV3y
UlpKwTYt/XxMDvHV65Opkc4TJ9rOj+4TTiPtNA1k0HsEL30m7xoGnHlQLthZlP2g
eh6MiorZIpGyZdeHnScSPTVIXQ1DqRDQ/RvhZ6oc1qM+C/vATkrR4ezPYqcHZg+c
/1xtnl7l170Mk0s0T7A3KolTVgiNoEKqS8QizukYen4sTOHS7p/HvjIkeuQwmQM5
s2Ehe3vpTNyyyaMYvcKgvlk198YkVMcCHqPL1X+orcG4brEfN3+YdDh9JOT12GZ+
0NMT8y5PEGHhaihPGKWf+BU4hI73G4YGXPkb9e+O6DoYxQK/MGywf6/PXcVCYMWG
sHxxv7UxiuhNBIH8qmuFvjGUeZpf/0/av5vwYNfJSJE+KdWFmwC7tYsvkUdVQltB
DH1PpHswwSuWSUwcHMjIRbxRlV/mu9XHYaqtd9MjofM88WdaGqtfsYgqCgmqWbh5
AiIbq1J224xnKNXjddiHz53gXWpN/P3KuWwqqJLKFzL/yqNPjRC/7yrLwFMnUiOq
vNuvNwlVE45nRJPdwVpskFcLz2uSDhzWB1rheOBUjkuhlW9dRHiIKcTOMzfPbI9H
BI+Vg/TSnCSmS+Wtt5El7xEpWr1nfJR8JsMWmELI7WnIz4LYd/GWdJF8X1/2QMV1
HVlWQByMb4IBlhVSwsXf8e9n6Cbdzv3dsq68pn/NKoNOT8Q+4zgpOIqfRtB4pbgN
6xoIbt/wrHqComb526qolCjrSa/iJ4SfwQc7dZp3sEDLmU+gByzgzwssY7szdSsf
zYnNK/zvyPlwrHpA2icj1yZZQ60wRWkVxnjJBmP1609WXVPck7lQVVxGlHqy4J+s
6uSRd/lgdElNHJo+YaP3ybsnDX5cx5rHWEtk3UNeo4J2ih1CG5Ux/QTzy8d6Vm6w
DLonygJP4B9ypaJXUveRylaHsYL8sbQczFAdFpEkHNr3OeMgtmzmoLbZu6Ob7H1L
8OOjx4kXr4nxqdCt//vX7udnF2Y/Ll9q6C8z9E1rh4MJX6cide5Gqr08HUGTd2iQ
H295Tt/IyTumxDZPzytropq6rabynNHCGMfAEP0NhlSWrz1v1XUMV/LfX0Lk0wcb
4rr5l8K8csfg7va8pcFy+HbMVR8MjebS5wog+NlAaHKOQCsuFRW4LTJcqOkJp2zQ
uRW31EhTrz60uikWDtdQ+unatwOmPKX2egHThy1Wwu8L8ER3cSHY69jMwjbbnQQ/
Zf4PdfMnbiR7hfTy+REo4N8izrhpF/8ftzp+VaUR5NHzpxAqeR0JYXPLEenjuDVl
Ib5vVQCzT4yU6HLYXnVb8mBB7KFjvnOm3KKW6J5tuv309DDG23e2z4KEZtYLdMEV
SXFTdKP7cfqr/CQbAbmPJfNxuSEeCPyQjpX72mGo12zZ0S3mqEfXpOjpdwkpAY6E
XUP+Zh/naV+0MVsSd6f8qY8u30IxPefnMknGKgMyrVy2XZTB60hAFLrhs/rK4aYB
bvTUH9GfYUmqIa6xMv1UJmUy0EXlYXlCtJyOEPbi/HUf/mL0WgqxPUsxyQyvjCbm
M5ZmKzuWyV5iMVHZbz2ub6ZwBOOih60dmSiKaQG3D2kltdFLfWW6K6cf1idEglQf
8E2dcv7zTedgcmwbsC7fE43k5+XlRHFvykMwawA3ksRXimSlL6goEN1Z+b1qG6yR
lonp17G5ZFMLm8DUTn+iSYVIOM3BpBOpHUxkIqKxoFFjTVObxyZ5FG7UIZqwBOw8
K3ytCZf4Ww4bE6oDcR+lQkIB2NSr176o2sZFcguDvicVC1HEbSZws9Ghd5Mbn5CB
/8b3JLgqj7LrhCHtgUOoYvnXCdJy0ji4I3Mdnb1p5TTCVyymItt8E+k/jE9rAPh8
hqiuGG6qV7ECuQnPK0bylxAMslIpKgcSvFLPDW2yDudWYeBwFSYKB+ypUp5oW4Y0
Lp0lpUpCJxlY3kFV9tFwjuz/UWfG0QFs4fZ/D2BH1kGSD/pjwIW3N+t6ibXYpuug
+gbghO2SwWfIyCgtE3Bdbv4fwpl/PPWcK7HJzi/eEuFfkV/YivhTiHFhfikr5ZAb
Kn3UsK11RNXplk6xJolV3YkEi1vEjt2skRoA8pYK8i2pYyXZfxRYBtI9GTjmoSAl
APynqZdW1XXrj2ceYwHNrJex7MP4XjHaANe7dvSVaSuug6bHgmj1MIuXflPFsWx5
cG3b4JaE+WcIHBbZQ4NZ2wCmGwu3HSXoXxtnUxRa1KuGT+OtDMOBpTD0GFH9rSH9
k7bfEh8js3l/gtM+gj9XZdgjt92gYOSoE9YjhrZoBznRdicVWyKFy3ICyKZUD9Fl
ZQRe5IxO0sIfgjLgChN03iPONp9okXxc71+UYybsydF2raVUJuSAyj8labLYTTXR
CS5wUAjn/PTZ1K6Ig44rBsoc8okQHdvNmo3ANu6wk+hAsr8Gl4zmunBHNZgldRh0
CmLLKKiTn0TBMKMJBRXhRE4DHmjN7jCBbxYzkEW7/6bIyz6cEdZMCANj4QpFj1iV
XNwR+G4Sd7+E/6fQ+MxiwG763lFpPMxywHaaB2rRB4mNb2QO8NpdR3w0wCc6jTaZ
YXaR+CyI3IR4a0HmfvTjALfNpyHDBRYTKuwkDwn761x1HSg/kVGdRk6dVqANFTNt
HcgK9YJWCtsDIKJZUzoLFDMZ8j2eljjonCplA0mHN+22Z9lch+QwAaTC74hv1cZ/
/4ELQZl4OWPgNm+4h9dTYu1x+gacrw/MMtU8qCcIYqzOIQCfaRG9QPbFSb6vZe0G
e+LcW7n+XmwHO5uLTwjWc7+MX5OGgUzrUR734SU87eqny1s60rX236ew/2zSGR0g
LlY4/rqhj2VvKKQC31/vXgwew75TLFeZc7SrlrErS5Ni467NOsqd4Xj+rlCrZSf9
I8QmpNPu9c4bRCe/RNP87wDzxxLy7+qWLR5dls4flqOVFEpuEL5HnszwikQ6ejtW
7T3oFbE3xfJcHbwtslprli6IRd8uQUDRD8b+iygEzxgDMoCldRSdPQXDgnBXst2L
gyg4ABXOmMBCbqRjMqbDRo38qfkGgIPsjoOAzn2amzQWu4/yAAHrnFZc8wgapZ0o
2NR4ozRJ5/clYs2x51Mf0wMJhKEWJbZNMiDWfZSdS7YGyj2nYEqIfv80KJSwloqd
1KzJbVYGHxcDiSQgco6IvqFtCdnWR4z4Z7ecIXqGN3uonewUc2gFsdSutZMV8sYc
Ao4wQOxNoDgmLVA8wKFif1VTa1gQojr2WM0i5ErhrJUgv483qG6WJz8YadzVG/fS
1rrQjpqAl2jBlA3lrV3byaIwwjWbjIn0ednSqqO93lKXvINIzcwm3da/hKmR5WMo
+PR1/GQJpegfryShrdjl/+AULvp6sTazX6p0rfNlpYRk08YSyxaBiK7SmE0SzHx5
EjMepTdj58SAfXlQFCtqfXcNS6B2+V4vtiA2D7TfBjOVwFob/LOcx2TMHBnsJfzJ
HDs1r+dDsMqxrM2DuGmZe8pggYCCaychYAKVIePAyI6Wxlf6/ZyUXDckWBnk2tOZ
/UX9e9aB9Yslu1X8OvbMf93xt+2NW67q9Z8w/y9zbVgpj/WjOIrpaSlsL60HViB3
wauUjs80nirC/9wI8mbnebWzxDKqV4DROpaTTIZXsazJy6HweUhU12NGTvkmYStC
21J932YNTwGlZ9IUSuPw3EB0f39kdetYErWyk7fjowhFq5gZzobV4x+RzUHYCpiq
zAewdIxfq05iiJjwCy2BfkAGAaRzIXhGHfPAMRVRGvCRtGVGx0AiPt2a1+qmgU2E
tvD9adwUmjzDywiXGOEO+xe0snQmfX/GfTdLAz9Bjh2R75mWYZG7qZvsyNO6eZDt
Hs8sKBTOBCi05LzZZfT09buUz5XoH32KlpmMQFtxjOb0du8iyIpfvwNLABA/XXeX
Z7R/zhubw3IJU9vf8nI1TQonqQA5yL0B2T/2L07mOLEwnduREhgZowJgSADa4jNk
2BWX4r66ooQkCY6UraqScCgbmlqFzq7YqyZLZ9rEHZhgOL85MLpa4rpHu+buaWgp
P/KgH8JLAXRyxYc4ziaW0yHyKDqBpQuh3DTNXEE22qicaT+ss67X+bCEaWnkmS2H
xAgPgUNEIHf8utrOQ94r2czSGcxqfjSfz/0ZGhQdRft+3CQQP3HPgcGU7GQxNGx/
6TXX/rgFA2wyGPWhqG6iuPe5k5nkf/dSJ+Gdh3tqsYC6tdLWbfISjbZbhK7MIUOA
R//3AJFOF7bBeaWvasXnSbE0uo3sU6muh23YHpZJE1IGUVL2h3IXWzmlwPGpcW/y
+qiawnrrnXxuzc8mWieTJGj1qDGBT7pFm1Ya6L1z4JO0tD3wZi7S8CSFYf1PmVJ+
FVrShybo/nD/kbZ7VtIoxZqPgD4z9aReYPvJQxMpA4Vc8fMjCUHMAMOwEj7ZDPCq
rYeSdxpKB4MvdyR1CLGOTlgVlDo6RbztT6lWmpJ3ZCG89cwWhOU5zAysW7RPT6ch
aE6jcTK2CtW5Az0K3daAfuCYLboyRB78tr1wyzqV72ImEneCSVvHNZClLm6PekD1
b0gjGZ7C42sNgWLBVkgKmyREqxiNuC8lG9Kx5yAJjs6RMjWNy9gtXF9B6vg4JVgs
f2Lf2IKz1q6fh3OscZwV/FohpPANsMqG9tQ5rP8+kBtGSa2bnz3Z2Hw3zwyMJmxf
H2UY14x/b9t/zxFXG6gEurMf62IEgEdMRITxRK5PJIKX367ZWADOuaqFElAJL6GA
PUGRbF9wee5Jci1AAAmhBmwA0yU4UGH9ETk4rYqZr6SjK6OAbYXkwsDdhQu2bWCa
jsN8rOXh3bfesm5BGLNH/9T4JgDOax2blYGw1WaLowRG02t/HgOdKV73lT7ZDr6E
IZzHRipRvRv0aj581rdyow3B1a6WMZKID+GWXbF3FLFVrfZOONAC5hNkAZwxR4sF
f8l5fj/Z/CePrTpaBsfE1tAiZzn9YY4XRkESDnEBRgty0JtewU99T6JSjU2E+HAU
4UBZKmvfeyBKCMCDgPuxngy0NQiGzNtMvZy9ThkPAIGccGKO4JUGoSJXKajtyp+v
nlv9qj7QvlSnhyE1lmz+6Jww3CpMTagE5Ij5iwOiqLr+2lptstVdXNexCgNqs7AF
cN5QihZc+kUHtXrLP8/2/siIgKUReb0F7WtHQjgprEv5DqU9WcTTvkqwYIcgkNO0
LrUc0IGnLDCAVm+l5d3T4QnPIWsaclJxnGfi9EgYgJliJ32qsTWcWH2yRcjdszh9
i5neuLE5gm7DQR/gLu7TRv74xqiHhaxnQUlhgxqQ/C0CS98eZYXLyECmvrKQYVso
YSPcQFM2t08vcxaWBFWIS2LXymo61o0BipbFSr4vzr3b0TTauQLX3EK70PqU4qBN
RpThiIiMqs1vOZMtIHJkUXDb0cL/zw5I3RorZAUUuz7lwd1m6ARI4UchZqtlJxn4
TQSvEt3pzLdXDLyP9MrOTVVTIpHYfQyFvGfw3AgOHnP4psXDlBRlxux/9BcuTeWt
mGmvME+kjhpA7vvSNanVW60KOqsSfyibp6Vstjf1UhF7CV+1UuZgfdjtyIe5ZqQt
nmHFlNgAalxVLQN1LOoHdAGV1oq9YRHmMm9XG2ky1JJ1GzO8CYVZqEmi9WpeL9Ie
iylIRB6yFMyAcMQrke567Ebny0JUEsC+kXfHeE4TM9VwXAJkPyDYtqgVRhicJ+kp
S6T1nbypc9drq1VDg5aZ/Mysc5LkDanR3snblLaeewnELP+jhl8Q+uP39NxaQDC1
EsI8LZqERWUiN5eVYTi21A8jo65Z01Ofc4VQGeTevN1rkwHpWwIP9DQkTwG1pRXG
lPdn+3lWGoePscfB/ihCIkgrGae7tRulFLTmoxS50UXRmwKs0vVBKHzy/vHW6Dcx
kcqaVeFj27FR5uXys4M/ucx6r48oK1ILNrKXVxRFKYNPeqnp/z0Q0pAd+NxDOGS/
C0A7gQKgAJakQu2G7bK46UbUnN10pTe72xnh0PQxqrAJTXdwEUP3SV9eaUHcSI7h
w2Bzwce0n+8JX4kqnrp8WAbAepN4hnHlNPRvpqL5XfHEWI6VV8URK+sMVUHZg6rR
N/mfOkB+7VSXd+11hITMZP8XbYnBe/O1h4N9KMSOJFqG4k5NnIL4JqdMTRPDsWzx
tKYG++6rrFCfFeRh79wpAKDhTDwuZUd4fcztRiSckZqI9gLftEpmVM08tMhAXcBy
SxeUvlEbIpoFCPkaDYMhSHyV6ps0Nk3Gedqjl9Vcui+eYyc+OD2ToqPazpA0Oya5
wdTbq7+ZuKLq/6lBKfxAmrlxA6/7qWwB7g+K8hXjWr+RLpy+YP30+kVE4UKHQe2/
/vIWN0i+hYVB9xipg/MdFXszjJ8bnar9oen2yNpZs+Dmj6lBTZihtF2uXvsZOkDh
GRoqvkw3xnQcd28rAnP+ZHKh4DL69WVwwu57NUfgzm+0ZyMv/m3Xv+IoWKUXQoEH
mS0x8Ol8na6JoGTGEsniUMVSxzIQoPWwNsWa9pkfCvE4Vw546ams+TlYU1q60U+h
lvATq9BEluDoF3f1S0Kh7f8MJy5JiarW+DTZ+rSaQPmXsBDKQKKO+Lh/wTKx9EM3
6bcwkvC84sfNCsTLv8L5Z+unVJtghyzP19+AdMJfM6BV2JGTO71aQyVvQ1EblW57
iyaS2lnnSISOse4nWIlByoBpw9QO5nCk9anyym7fGp+Js1A5cGzC/HVPTuUNJOPm
3BcDLMQ15bdTQjwJD5BeDlGtINO0HHaPPicXyaAj8NcQibt4M+ryxcrR2c9mo4yM
0JvC8y7omcaW1x3X4va5avGMlrgqQF/5RDtAmzoECiPjky+loYkI24S63Wfr/Ee/
Sfk0WCkpkj8rlj9/BcNHmwhp7eYAZ3jZ/3w+UbRNEhpdzmocN8u5l9/YXxVZcIbe
xxMhmWWFaImC+wXVqXKGeD7KzWrwBLkJWSexxe8sQvv0TKeQ7izp6g4gcLY3s907
whRSoS+bgKLeW2EPts8LoNS3zGI+Km7k147RsENnz75yQQhRpDPnRom0Bain2/4L
nZdq19JqAEGtnN6n+RKvanee+G2aE68bXFvOaP2Etc40ORelPy9s9EWh6+lxWRtO
2y9FVaBq6OCydfjzk+XZ1YdPLcHPKsHgjAqNZvWxJKeubJkzq0AG4SGTa7JeHq+1
HjGNKdd8NdqVHT5D/4j42T23zXlIQFaCWd06KeIMLA2tmm/dkUcbXTUbO6+qAGzw
QxiYB2/NfI1V/aj0ykL21IbVkhXW9cj0onSgtMISt8n7ZbVXklgI3KHvaKo2Lzlt
yvuS2OFik0+SMQiONBKiBnz7frYr4ClC3BzK9xmh6HZ9KpAWzCgj2qQKUGoEgFv3
bD/pkb9PPHa2PLNm7YpHUpDulvc5mS/JkPwzaPQwGFBLVGfAqDpaM3gteJ8obBVp
URFRgeo4PQNaTl4ivPJVfl7naZienZp/IrcjgBldMtADz2GaVG8TSILc3Q6mls3g
Cu5AodpF95Btsd5JdFo/bbcX0U1vl1Iqf90N+IDHqSMGbr4o7BBRR7xFwTaDZA8V
tThMAYuLby/pEV9qkLDRZed1/7h75l1RQ4PLvWHPoZTmdD+FdcjXJYk5xi6qNAeD
EGH6bVg9dy0jmCVvIjaCv+JmKS4OiEq6yENdthC/THGtut73rgs9DZSHnZ1eofEd
XywE3adRjrOu/mql2Tsq+qZfB5pEji1NIDWE/udjBXgQP9ZZpPZSUmXZgknB7D1b
oa0lKWsohxloAV84qiYIgWwUhVBXXaklf4cklLXAiTCeDorxc8tsWg0EVXedE/Tn
6k7s2zWCA2j4yxn3BWJj6z48lT0NCj3ujup+R8mOvJ0pr29iWyKY8dbPtOKZLiOZ
DHz9lSXRYCTUJuMgB7gJRMocHBrJvYirsCG85PsgsHcFGwgc75Ob0MkC51siimWP
JX51bK7Qm3Mfd2OCFFZtkEzvfJVPrQ64et35KO4yxFnMSbTYJQYvP5xJMHqZsuH8
yHIJl/ZCKD5+RbQmDOJUTGYwLROGPrEvT6IVN3D0IJnxpPoCcOhX/QBOWKaEAHog
TaZyWMH4EV6JbaC3yhwQjk2Ekbe2qC5tfuRCQsEzV9goHySsThTNFtHtzNtEZlTk
a+g/zMgGdyDTqlIx8B6mQTEXBDWQMXE6Szpmw83IOYdasgInfMcbIR3ITB9BU3jc
k0Ygjl2Xw+Ju8RNjNWVb5Qenxbc9IbALhxfMrjizTUv/GVJzPlhDvrckj/TCCl27
eTw7WUiN9MCRmab0tcv7bmfYj9EjikPIgmlQbmaPzNMKlK5gSZaFQtrJ6dH23xn2
6TVXlKE+GXGQG2j5B+EJZ0JRvbYppInb1ygjKQ78bbAGm+QxG2vBezhuu6DMjoYv
BXd79mQfOT4NWhaMDiHHVFJjMUaK9r/ziz/+SV/KwQa9GRxvsNvn2U/RpmnTKzRN
KIDXA5KGoabjA0EWW9gy4FEVOtYJPejIlsDSaakmwmRTb4ro7MovYrg4QZTxEaHm
msAWjGiCyTmjv7Et14Mi6nQ07IS3VgqoYhHRjmLd6TK1cjH8DLvoNn/fq+5o4sIQ
5MjlRwJ7zZsPlJoW+foofIOEEz+wdkm1qqGHDmq14PNQZxPinstvRucWZO9FnrEd
l733H6slVmPzpKhX4wF7BHQXaKDmqLuWi7O094rXcJFsRa+1uwdmnCYcZJMqj70y
CMlL0hz1endmyVTffdHPU5AZcZCSHYvaI8RhGwkRcBr+yqe3biUBCfcro1A065rG
jelSrOWP3/Kxc2VwJ/8T0WYa0pwJaRjQOGGX1x7PN/eFNahACVKQ2JedJFDf+uYn
m/i/ogGO7sszOEOiaSE8vHqF0S6B4Z6nwo9Y6ebfEU42FmwTzHwVW0LovJlbK3+p
iWw/BZCMv/8XyWXL9gSPF8GuwC9WuDMaDFLvgZrD8950kRzhTtIIY0C5dW3z0GWz
v0n9niNUwEaYnFg1C7U+y/Huqf5Zxr1h++odADrJQEZd7BinOIh2ZJaXpAZ4Pj5T
PjimhGoQvIK18K6iS9QGWhs032AVFzt4weSZ3OUcBl5yx/ekQNqAkJH7AerQNDot
tZJA9fD4nCgaf3NxM1lL8TK68CYGAHcxc8bfCEDEM2DRhOg6icaCEc7AunTH0SWY
tYYiECqeX7ri5cRKyF7oZWYKpw0gD6HvRNjmMqfPpez1znAMBIhkhicl2XlxcgMH
oyl200d4H6zQI3GihaF8DeDWIxgKxvz9eDZzrKA1tMYuRwHhXTX1DouiOfYkxWUD
sDNDmBi8iiudbIHwX6pR3MEBUS7a9+3l6pKcCLiugOJsmF1Q0yeIXLhlDbBGySjX
jXR9gOjPWZw3BIsGnICGW5GcotQEvUHkIIzRwTNM5SxxufB9EmTQ0NbYLpyPIJc5
bdiyJBoJ/kgTUDpM5eh6UHBQ2+fD4/9hZvxP863k8bx59Iu4b8LcyFqX225v0FGt
YT4GOP7erwJFKMqxP5okAt2Ur6GbrUdqpa78WpBsVbIhKeFhRJlz2FRv9+UZBlmI
aU6DZkoCw2K9xmvv/ybg53h58FZDAijhjHo7h+Ogq6MK7YH18L5s2DUqdwa8z+Kt
sBN+yw1X4KZPkzdpiJP11ZqLGz1JB2HXMWD6aI/3+2yGBNbm0CanAVGCvi/9ldS1
rNn5Od78A14lAZA2iAjpjCgIOalE/MWc188Qg2QePXHKDaesY4LtihgJ6KeupzMz
E71983c4eIoTSnTrmEo8qt40HxIr+5d126VkYFuDjFe+5Arf39ZspD48u4SvyeO/
5SxrGpvk6xqHJLVkzUMPOsF1k9ptYXAREZHf7wAe4OeJGk7N5nS9tHXB8kUTmW5b
W3aiqgFGiMbuhsPxWLhO7ZFCGZ/RCSiCXboz1sg8L7LyWVAPXM3gJ3wUZd7ncQWc
53UUYpptf2sq1jKVykDM7EGhbGHxjT+mdqFls5sSe+rO3+phMykWhvONak2wQXdh
8uVSG3husuVQK5F/mEr0VAtpSxqq7pSpkoVr9iUeBWPQLxLCFB2oH3lT2Xb+D2Tl
wkOPbZTgrRJwaiTOsuQxs48oU6NkuJKIwl1+yNpOQHSs78raviA49TyEj89O1kCY
Xx2kZagMYmDjqtGlwKfbUTOC6GIHF395nlX4YZseVyv2eXDoftZKN+2EgrvEMdX1
6Sj1Wa//K3MHWkNq39jW4ulys8pSe7BWFL1ROPuh+o0lGRssrvrrtAoa+CxVfmCd
ePejy/KBuIjjZ17Zy3LOboMFzJHOMDdQ/7IPplgUAGpTXLrdfpq5NrMTJC+o/MVH
j9g29f2C+h8FH0gIGngHtGiF6qyIELZPqJGxY1rZuYRNCHaFeekbkfCiHcp+5O+P
FwdIelqDZmDs97YzTxyok4ekX+M64v1Cius4A8sziVKNgsfC9Z7JfqvMLM9enMLw
O7jf50uYKL2sHQ1cHA/FlsK7xpbMLMQiElQvgwjaaQu6K+aN5lV5ITwFMxyoWQLT
PC0zQabGfr7EM3G4MaeNPzyMfUZvFxDc+NPmEbC1x4BbR8PWABtUzQe0D6DB5CDG
mXaZkdVQdh/pF1XtzmlOOEPlxvZZepBbe0qAveSN3uk9SzxbcDbfY8Hufhkayagl
YEvtXqI5aF8F6bYixvBrDc2XnOtqZ85dJ4B1uLBpn+mwdkA7eu/Ifz9tDe6XKkp5
yYU0vjVuvwaAFr6sIX6AnF9ql3+vmE7zlzkuyu6vgr4NPwDOTS5IyPYziJzwmhFm
jQewKc5bk4tkQ26QzVIjq3scCkB40T9WB4PBBBW44KvbrqlrgVhuwltkCo3SmMm7
kSd47KjRVQMkUcbMb6eTpf6yfvtBX/4Qx/TfLx6DZSEbMnEIbh7jfoQdxz2DouSg
07xwTbiPyDwEOsX7gj/oX05KTQBGn4RkDiqY7hc4xzmslBOwkNP/ky48vsNMzuQD
GFKTGthg5YtPP3hp1HdCtaB8+BlKxs47VGBELKVELg2qow8QFlbPmFq1X9XjlHY7
gjF974yQblWPKATMJI14unVO3fOhjDWCdtmr60WTZ/Euh6inRDDwCx4qGLYJy+tH
Z75zAXEkCjudf1M3/ZjqntrzJ8rjl37Xmlv16LYYbXl7+Ok6E1Jsc47zDTeW5uFk
utB7H5Wh01yio8Se+HrH/HfhGzScqIJuk4za4lry6vjXrhn0O/QcoeOAGxUwxUPK
3ljSw4C/a3mOKTw6ic3DtL8pAyal7ptNC1PivrtEHyEF6HD+G1vwSb3834Kk3GEg
LG8AyLOTUT9zRU5Mqyg0bAVTsnVGKULT/YEWldrFLF4nECB1VIECyPZqu61mMfDu
rshHF7W8AUGIdWf0YXl/inp/13Q+eMS3vk7H8rxCyeutoMhKWP4j9Su3kDhXYdI9
5+XF1kX0zb3Si3px9nbriJKEdnTpHRAF8oAmKattDLjGr8PhVdUh8xdtiY6mGAN/
DUpoxcri6oS04WlpDvlRpyAr5yoGOJofmiaXPpIZujj6mB7x6XKTEzxENyd4C1ni
RQ6CjVL9g1Zlb/hZUPVMVHzG2MKaMuwggyLavZxVSMy6x48yWFQO9ebFm58kdD0W
I/KF5yzRkqfNDAoLf08Gfbg/vRpj1DgU9Tb/IY4MyAnPP/qqQ0xi8Fovv/gKL34E
xgyDv7uzVP78Cff5D0FzqmtgyZPCvu1NyyyrA/nbB7TtV7eUPy0jpq/AJEQe+jwu
K2b5eTHRzUvMtUIspiqLVb1le+dnfRM6AvnEat3p8aRQyp1YgdN6wzS1yl82CI5E
YN9rnk7OI4F/1AzExKjmt3Rc4r+xUEpq88oKB4e+qJQF0TQlxzBkUt18hwqiHNFJ
Jd1ai4gWVGaeoi4qN73VNcOxQWWKIZElBxt2cqVvub08M6ea6O2V58biQRGonH6e
OUutO835obxfIaiEzJnjngniHRttU6YIhYvG4kCW/Z9LehtQLZxQ5BBlKqzZYGit
PqBZQBOSspvUnRbjf0dH703cjcmigdzd5nku1Bn8MUvH3Oo6tdtZYEv00oK4fkMg
gOZzqVnmBIq31c4sBWTzJ9aZVDAxIZpCmzmbpO1bYleTHY7E4bT/9HnrMeU3zN5D
Yf+dGBLzxJxPh+oOg/z74PCvGG3ywCDubXONpIJC8v0WOg3NwalDNxiYOHVBKSSh
MCgbevO5BNq2Kdp3l64qF914qzTgTfaQLgLbZlYqGt4Z4+kff+y6DhnAyGWd8JkN
iK1rHhu8oT+Tq284Zd0aprFud9TucwKAxskOq3eLKwo85Wgnd3R2GOThdcVJVE+P
y4o7Fb+iwZFiz7rC6e6+lZDNyIhQhoc+4onG80eVYNwngNY8StZ+Ett5bZXxYY4/
c4dSpbCGM7+aRtCxVq2EU1SNAsYnReLqwb4YjWjPzVHdUQwYsr8ub6CPVghXubwG
jtksVEjaelZZcrU6vkeXTt4E2uVL+quBw7fEf4HwIk95/Yua+i2JNxU3hhtkY7bg
UBeG+vEl5IHcd6t54wTZykekMcYmrBKKTgWyjBmiLsw2KTe6N9QcN9B3+R0neNlI
NanD4P94Y+P25yGD/53SrxCDgzVU++g1hwpPdIaItRITdmGp1xEN1DZ8HuGtUF1Y
djJxcKNavvpvnypOR3pdtPolBFcORp/Rer1ZcBq5ZH4WT+HJjWlJSFI49TojomCX
pWmo7s1lwyS0x0EaVNTWGRZ23yA4G3C9BpXJVeyo5Cpc/oPsMSGA1T4UsQQsVOou
KyK1yBkNjzWQcHwEygNhRabLYpJRdc1Rd6p2YvnfPKYG1PXszplMhyah8jjW6y8C
bbdshXrsDUG82SN2Scteurir5OgFtU9vk9Q4nJjhX4RGiBX/QBUxSFenCI9PezmY
8NeF0lmSDfIbOFJN5gG/3vYR6T6Hs9uZFEbvfgZgjjQDIdDZ7qUL4HjU/hMRpiM9
iWohOqVyl1LGW+nIayZCm80uWxS0cYA/l8FXFMUiHk57nvuVsXdd0TE4vJI5jvJ2
dHuzUP38el0u3AhqU6c1Xguhoxaq/xIGIEguj2QTpS+jBPqCYsn6ATtYH3RhRORV
097IqK5o5s9q5eyNXX5z0kRMwTFojyeXwUJ91VcYIoJYSLLYtwP/EdQpv/JR/U6W
XpxXzMVOcqCrq46tbi2LjcAIXpYj7IiWWRr+QqBcp9e+bN+5JLH33j9MEabKDEek
qrUggl7dA5/6cguvA03Xe4Or+CV878R+S25zkyTZTGwKMAYvZdGztEV83xc0i2tf
9Qp20yKf0N/6stzSl+mlBNdVj8QwTtYx2KOEKc3LhojEZP3zheM0zqTzbl5PXbj9
OAxySLrlg+CX487DLJ8Ghf2S/iAvy1KNqkApsxnws/++Y5KX4KhouhT4ik66HC6M
kM9RBfKawdHVTdRLm4ppqt8EmVjqu6iwusMTYK/btl+mHJASQj4BZDn32hNXjXyU
kzf0qLWvhQMVO5QB0vsJjZnkBRozlttiLF1BE5in7o5Fni3H4zBGlxUINK8fQc3w
ilJbdHSdQRvGO8Wc+HSqpa/LMvQXbHKABD3uCrnE3HM0SOrwmeHuefvQZ8RIIYlB
QEB+t9B+6H3ahonAE7F+VhD0973wy5IKSy8gDlq4w+ZG1LUJJDBJXzabibRh833l
VCBUrFlEJ3zA6+zxA5Fiya9SaYecapocyJDpMunv/sg5pRyQDkry2j4SAPDUtXGw
EH6oLnx+xVDa7qQ6T7P/yLz7giOeAW/NjlEXlu493Hd7FDKmznXPvwmMnGyeJbRt
PLfzs/Q1b2ETtZdzB7O6UtLj5MUa2ZGHkHcfVhz7iit61snyys1gcE3k6NdFfI8k
YAclbwIDHVLHhsmx5y5JsSbZRZYHdJw0C+GgQTfzmjkWEYWaGM8Jo3X38AqRJHQj
bRSx1HDc0lCddvkosR6RPaoc8PNYb/dweStAvDXf9bzNQB159IhSD61yJ48bTHgC
nTmiZ/21PPlcf3gsbefq43Un3KVOBOex2Qfo2e/m4T6Y1OtYSThS5IFe4B7SqGip
khCMhZXY9PkkVBLZ26M6fngIZOp76eduPxid2pYkw3FHkQK5Hh4OQa8NU4/TUKdu
h39huJ4bXkjhAsg0vmPE/x5bg6H/FtoZPnRBHtWxq3X2Xs5MKB0BX8onZDozkxCN
UTYMDuVg6CHKV8ZC5zndkgCaEoawekldT5GL6Ubi6DW4IK0U37CZRTDymfD+DudT
fjmpY4m21CfqBnnO7jgG7ZYfQKEUhGbVzJeEBPuIMxHHDXC47b30b0Fhb86mhgLm
OtaTaj8n8BF+bqBwOsYm/TK8RyXcM721AhFvksWem1uJxC3pNsEnIsy1NoWtUZYi
ChEUY6IuboRrlIWhQx/gCagxt1X9sM2Bpald6lAutJN6YDQ/5bfh0pjIZKZS/b/X
6zXxzfYGMl0Ez8Cl8aiICJ93MvF0+iMqZWHlHiED5n6u10RQylIvhVe3iPAZM5/t
8n5GO7Dn2jsRaQ+hpYngqaLP7m1zMMCkTCKAvKsovrPS+b3vYmiikIivPt984mQZ
jTNaZxjcSWvnQuFkwyLgAPUCg18Z+AK0IjnNBI2goFSue0L45ixfDMbtNN+n8c/U
KnG8r4v3fQYQlOPtFsMof9KX7yJdcqJOtXL2GjZsQ2UtRJneu7tf/P/WEV0Wvffw
gOyRsu4Xgfc+SFuEH7Hy/QIK53cVlxgm6W3t0NcdwLcRP6jfx9rbI29U9+Maj/hi
u5ixzQ6fm+JNXlGgqkMa81csOY7XZ1dwDB+ZG/qyXt4Y9AI9vVcNF7I2A/r4bUMt
XkINgMYsjfgkZ+Z41pVLQVNME+vdb+LFeW4jI9gcTzl6LZ3m8Ug2LyaAVXpIXeLL
pzKIqyp1alUY68pOLRIK/6D5SQcp3YIRYufnBEP9dPcvGyXRRwcbY63+QJyeMzJJ
9Ph7TAUrzan5b4dFAQGyOSIu+PtGmp+HKVOuRQiyvfjbMRr5IiB6/cefkg4c1uiV
fFiDg/Aj6L3/qWM3p+s0iYPQFiP+74ZHT+9b8kOQhinE46xeZRAMc2qqS2bZawaC
Xhf4vSOWXgBy99+SFIt5dXw/SOEgIqmj6nFYM8pLFmIaopANWcA9EV+o2UgpMcg1
lx7R+eAzTZfKEHRleqF61XFHr6+UPJHujx0nNJFO6uHWR4Z7WaN7Xvv3KSujTPSF
DJfHuf6aCC1sYPVuyCOX6nMxUvOVOpImvVsVgng9x1k//TkJ2vevQvt4sfA9nV+Q
3Xa1VNZVqs4REvpq/S0ghXML35zt353qBVsyLbWKbqiBoP/DRV0QTmNugTrWijT5
YzbkcJ8DK4DKWV1DGUf3+q3zX4MiNXjQa4XizR+qZV8efgM7uExEpRNpuY0nAnzV
LQp3j6KphCNCP9mQx7gn+/aqjEV65Sf6fupJQdG5r8BL7F8+9In0M4kP2R2Nj9Ec
fHdb+6LqrpHON/VZWDyYInj2OfnPonxPF58UCsKBZcxONq99Cy85BHl00FC7L4lQ
j554hl5LiY13N4itye9YNCZJWa4hSJz9y4m5FL5KsMe++t74fBlGfAIn5pPnwRuJ
e0aSRHjSzCZ+o1Yq7fdS6D0KEyZfp7f81tEuqxDwwtjz0wEZVLd1Ttk9JBbByJSa
YpVMwRTGEwGrIHnCG2pjHZWgBusMRvatARBhJehUUQEjYQFf940dKPo2155cojwm
egJbMsGk1ybGKKycGfCe6vmV6HjUAWBdsmfVnTsxwPf8bj8riBmaWiL/Br/9H2TN
6sd4qPj4/15jUcRFg6pXmDzDJ3XSBzZLpSAZFPiTxR4DCt2tPOQVBUuqsPIhfoZM
P9k9x7wsLn4Khu/TjMCod+PDH1IMNpq7ydb5l+S2GHHkH6gHyP2IrwGzxUiIyhdg
um8/PQRYZ52crN9uTy3E5Vc7OGPOC/SkHqpBIAnyN6fAEbQL2Vy6lHG1U6nQo/LD
cup/95qQCkvw2vyboIF0oXN/SkTJh3eFyfhAs+cuil4rBwvWjN8/ZApiR7rdZmXk
hthT9cVZ7T+IocYkX75gGg5kgt1Me136pyXd1rYH8pC/P70GkrXnL+c68SPfbkBk
9BoF/AIPxgqUlAZzvQZVdEY6L6eIUJDcwTv4UWRxmfJ916GQV378MsaV4aIf8gEi
Dp9sdwB95C/NXzsj22LwI9eZwilU7slaG64c1VU0ODtLzi/13I1uqK/IHkL4Lpbe
9KPPwkNHah5iqCddQvYeMmfs2LflNlIXtQqgt1iww7de/HvNcjYff7Dgm9dCjdAC
3XeR6Uj09N6ZqR79DotVOF4F2cIyUGvTPyZk9wA0pa2PppA+fepo0HU0gFrBuL3y
E1Y4EhtBUrFZwhG9AxOlq+38OT9PpWOKvGeitRSpjgaPwe7CwtGshWZ9LV+NEtYW
eAOnKB7JOC4TcBUqei3ozbzsHQ7BanvpY0kXtERW8Oq1B2afZVjoFIvZ9qV9BcOL
PFfMdoIqoTrVM2SaaW7KCNYXf0nxGE3PKaZNbjtb7oRPcVK1GgSPpcMzdPcGvXHI
5v8Wo9g5zsswTqQ314N2fYR9Xr3JgNSsQQimneUEATdNnev4h30XK25+kqQ9mQI4
/sdESzDNwyE1FaWOamMscXNRoC4tsYHzfgcAzHxhCWRivVS/+4zyRCsGJAh3tPWE
2vg9MDQ2k3e867emgubI75T99m/ucTCrI8TQHnof8dIMOqpaKQ24Fq9PQ+ZHXCuy
0Kj7/dzFFcytjrjduy4xDPweKZJugLJmdkE/eBnQacyzQ7mvoJ/nhpqt2howkXxw
lrMobUUmOuZDmsTkUj6C3gKkBYoh4HAK9NwSoAlALr1pg4V9UUMcNXSDtgyflE2y
+NTklWUoZ/eWVAbo6jeGuiPXr+zxhzHOzvXNRon4ElmuwBV49SItxgYj67s9lAvr
9ez9POGnAZQhYp4y5DyTiuB7bH0r9tVJQ6Td+2xxk5otzd19wDCvq8Rou7WXJ94J
B4MLtNnCAn4LvuEfQN46TMqThBeT7zfhCN9jvdi1OlH4NmS/BWOrUXLml2cTVA8k
9qCjEe9jt4fQIHccQJnIxdcWzoUM1mpUh4XngtG7xHW9XHE7nhXJU7mVWhOqjGaC
TLXCWvjGrTH7j+nlR1o3ItIuceSacViw8Q893z4hl8yNunPvCzKG5bgW3DBw9tFp
98tF1kM5KsIepUGA0z6Pj5lcLUZiI68oLWAha/MHp1f55zp74odBKiV9MLFnV/E2
G2GQ2ZckSK3KplKoicGAyUbZLE06S9DnDuuXqO1ubl5Xji14esy6RdP54DUDDSKu
CJDJ9FmIRDqTJKOSFPvk54UhUxG971wMAh3ZvIveL6EjgDJrj63QOKQ0jh3yP7Hz
fp3rOVCVTR4CEXI9NehJnebunRm//OFZyhomQ9sbS81/LA7FlEhU6dKD8bePS05t
M9DSYchiDyARq+KbeqamcEy+qbA2onqI3MG/baBgdE6+prWcnYmrgVgyvFM8eEdm
i8wImAE5Co0sU1XV8Y4RXN3yG2ZUIV6RpMX16lk0FhbopUUMtfRvM6qSyelRTT3M
OxgQMD7elm9n0s5ns5Ed4kgXfjO6ezTXGMlbjx78P+M61BKQG5a8iQryWI5zeS3R
8vMV0QHSveg4mdQnQTclmXXEZGZhtdvdPndoa+JlQFjUdzRKrQpJZy53NMkDDV3C
t9q4uVaUEWFS/E58+KGZ7pr5oBsg69MTw80rCJo+4L5/bkPVhNsNoOpa+tWWARDD
v8c0akQKOL6bqIIZcnwtJYhVLziJXbrFtXvEPkH3SaKHRyBaJS8OwgHqomntxs54
WCmEWac5kD2LztKQ4ikafaZz1oYZrUHw4kXefAZ8DS3IHhqN5J2KTuYBXnLAPDXr
hjUf4aeOa/Up8jMZ+f9pdki9f6xrUcX7R3NuL6YX+3h4Vabby9Im30faSYBQAOtY
d6A0ZiZD34MqJeA2BprtVdXsmtJN8dyBzQC5ny8zl/OTSJVYzUp2dXXcPWDbb4qX
TUNtgIqoxsQH+AqOJhWTtMNIqnuaR7OUPiLiNyY5yWU1HH8ps/s0hlHSvGbRyb+o
eokXgGKiNOriMQStilRNo4D+6vRRYDxEL3yNtXqv2u02oCVaowaUU5uZmvpwNws9
/PRf/Mm2rliI1FqCc+YxYqBTilc+eL05Zz4EnHyF7O0IAKDB7iAgAivbYzU9aQwX
VubIXUL7iI3t+/93rG53od3Jj1IM8ftQd4vObVaV1edPeH4rEQDfEsXSH2q+jZn8
cqZa4NMjuuqEodKaJpr2MOOXJRQa1SerUYPtghDZk4ulSRKjAS4eeR2+pRJz1N/S
c29cj0lNT04TyXdRnIbmavXrLBpe5cDbxr+meoU6LxM8CyPi1NOlHbDgkdlsnV0U
Dwf3LxtoD8Klys9KVz207VuvnG/u/+4Mpn0xY4mQ/uL8451rVIN5z9+dE1uH/blv
ftlpsVpKBGx9osWW5bc/XqArXJMieD4Zb1hY2d+49Y3IHeRJxs6dciRRp8kJOmmD
nUXhLbHM6RDSquwumhnVUjxBhSJOPSmrlCgllptv5Xpb4RftkWI/tX1Kdv9btZyP
SFpoiFFvPo+iMjtAQmEnT3h3riAZR18HSbcxHqSuSDG5+JCvIv+wzyxILdyxMJlE
JWUlfSsPubq8KUXaO3VRPumFPC7MhwOxmGnJpWYsLevmCkrUfOxXThzyOePAGMt3
a4H8q8aeZGszR5gDvKatcsCGSqCdZuKnOlmwrCDa5YNYHux3Rz7Jf4gk6wk1dgWl
dMp7DRA8xWyTMkb1VGL/IgCXKrBmn8h3TEJkHuh3MY/oq1aBAxQwjmNi+qPKKjuC
U+vux5NRr6nc8NvFBB6JJT7qu45K4g/2t5z1BFmGuD4a8WAv2pfZBvqPFF7pZXKZ
Mxp3cQSQflZ6766wTDuyQOdRnn42oKGN0IRYGG4TxQDE8M6+Nn0FSipEX1AWAIO1
Nga8WOdsPXmZJBwBqqUWUgDrbRSMBYVQHw8V4lIiMpX3Ca8EphuTWMo3d6HYh/kj
Hb49JuKfocSoRtkPPuk8SMLAoU/3it5x7JRc00cSXHrtBD9+dzxLmo/ZzbgpzYiC
BRaK68L5V/+t86GRZqY3jPr06t5PWNf1/Au/gSlFyZQ+t35NXP1pINuGXAWxD/D4
gNcb1L3TFhGxp8+RF0ubcnCC0aAneWbHi77Ci2h6QICEnY2aBNnjg2whLrGRjFMD
lmdEQjvlVkqPcIwqC7BGYSfzQjWsss1q15ypt60FH+KOBQhSP8HTDExRsmJDURa8
1B/tiyvyyG2ZRNMWY7qh3iXOI+olUVgItiSFyY4NxF1N8ZxtN7BYvZypazGthxtK
U5ifTDqW6mx1p+CGZVx2na3uOn50fRTegON38SU54YnBuBSvwGqnsvj3xuVSrefi
Rhq69pappdQjHxXvibNOT7S9HmCLjuwQTfbdGY8wrPt/vwkUdVMx1jWIawrpSQKj
ZIzUEkBBrkMkrIZswN/7Kpp6/FjPQ8RdEGcObS6LbaSlkNrJqzDKvuweXsePzpFX
/QREHZJg7wL/vkMX1KByAJE5u8gjGbiq5RWw5Grv77vE2p29v4SAM1rGBruF7DCP
FWyH3xGaVaM9jxjnOOMkPUnMxd290nsrkRqaVxHogqnGHrV+PfRxirctuI8Y+qeZ
nJwVdjP+u6lLMgB8y9q6G8eJ0g66rKY69yhxBwUB6avXtIOhUOFkp2kjjq9hFaeu
O9nBsFM3XOhDQaiMYJsSxTnqO0LHAo3c5sirvskK8Px2JbLmF4/59WP/DdA/DhkH
a/Qk82lDr+A8x6LpEu440ksg2J849Ybp9a/Ugv58ZoHHP169lnbi0kUbyffWrWqC
e17y4/qz/G6xflnI0OmTT5qz0xxikYhCY88BuqkXn+q5pCHd+2xlkA6V01oFWKhs
5Y7qK07DQSGPS4TN4U01H8ECuvlUlJoX0wnp61RYSnqOJgiaeDcZGMSl3t296DU1
FHQzKc08o9oPhuDdViJcx3hLRnHVbeVtquWmEalgR/XqsJp2REpqTgJPpxvH9Uqi
qaDu1nLbUpT6hOE2M4CkuXhFtPtQUsMkVIZ7O+22vVkiDjbjitgyHSStzQz7JP/D
iANdot03NxECw+WS9p7FsI/ddOfOPj+yxXGY2DZZHJQx0et4S6GEMPUXK950TGJ6
uLMkRSAIU2JDZK4xhl1Dkv0cpNTZ0QFNhyZEsbe0TJGMeDimWToRQCTKDlvb1wp+
GBDuWhX6nKrS3DAkKx1DvLHnB28sakdpUQ3nLR71i8nczGMdXGU5qBW8+7Tscqi5
5ieDEDY/acEH44W9fUgXIm6P393Bm6n3XOVjVGlMG//ro8vqoXry7imWlm31RuOr
I43gzpARLCIaF2SWkIoczzjSj9pll8LNBc2WzBPtTIB5niR3HmhdCXQmYKBJSzC0
Tac0+FHSjr4iJk6kWZOyxXkuWAjJYHlDttkMYHPUTR6RFR103DMHz0xABk13qJ4k
W2JWmfRUafm65Uubjwkj9sOAXnDRXosVZtTH07xhzcuoLsX/DHzNcYnnmoCA2M8c
9GT4Xc6gqwYG8axrE3XsQDJmPU5ozNUiku4D6RTl/eW7YcHTXhpHUoVdVDXWcNYR
lOxRppjevB8dIXdl2SPhi+dMk0eSHA8RMqjQnL+7uYW29Mgr9lNXv/bbF/4PSF5H
P6yyF1bc9ptd7+/DzWYfnUxjtqPJzBXjie1am8viHv38MhOjIL4i7k9hZuk5d6kg
r6zkpqAlKFsGps0o5VA43OLZ4WUmB5XA0+bh0g1qy0NnFIiF+pj5ivBlGuQkemQv
A/N26ImeV/VJ6+grcQxu3UlSgsI5yukML5AX0pWev5C7B+EtWV8e4rhSJyOg9O+j
gVD87udGVnILu8Hv+ASeedLagbAOjFJnHMzz6rm199oRXZZJzBHp/J3iJx5m+Kto
coTm6015RKk52elVC7Nwf/ulExYMzrnkI7LLUgy/JyP1SgPRNv8oBKfNz5Kwf11g
w98QkcdJnqfnzeZWhKvmlsizdCf5Lq0x5yah5w5eMCJj2GYvefdWuzBrFnEzcFqJ
GDphq0zhn6Uf6wnZ2eullBi7e2asp6Cg1Pf/gfHsQ7SJl+vaVOXs4+bBEu2luHXV
u+bmdPXCQFSKbXZgl1k3OB6osFQLu/ZXlbHvPgxuF/53hPUISUYWzvBxg/ngbWPu
4fNmxIeh9qJo7dnvzsqWPSbt8bovKT1AMaf7Yy6anmqauqmp/dAz4L86iO/1Jb1h
6ZCtz9zfLy2NI5YjETaJ/nTI8zlh3nyUfvPIxs8UfbvR6Cweih8O5Ogt8vP3Fn84
djSxo5iL8QF/JAwpmaU7aVoyq7dr0p/DZtswfrIVz+LLwkDQeSbU6RU2RM69pqYm
2NYZNucb7sBdtz+hgfVXckkxa8xDCSqzflOgdbulSzwzUxdAmfIaFL4c9Jr0L2f9
ZGC1tYMNGwEiCSGAcUlhJgia6bUUP8xgKsz0bQpaheVC+f47Gj4CQnV3An+ZnXOW
n3oRjWpCQ8wv709/rdgyJlnE2KvE2qeBgvMQHvK8eP0+n6EBanV3XPa6gPAyMWQN
3quUdc0IItYjdr1RZc9oOwbyhim1KHjBuilpwpE9d0+LQSGKvpw1fBUNq/xm/EHt
7pCZ+hTzeUKbBcaGV4jUI8mUsCuPWa8Iz5cjT6rFlxaqwYjDedNKo9Y/q4KCTh3G
1Up6HbaofpJFDUb3yLjGaXahH+mpTSncuPU3532Vqzp8DyOm7Br9DwkJqZdKo78B
HMUUYXnYP3cnZgaMoNysaQfRPLKBVr+7rY5KgMjmMMIQFZ/MsR7R7T2ty8WVaqb1
/GpkGHSgExbNXULopxmHldNlYt8ZDLLXm4opoG+jtLH5Zfihrv7Y1V6KzoD53/br
gnhqOKJb5mIHbahQ2+G2xD5zQ8remEXxuG9wcWTkOHE4u+jo23nqJ6Hms6ElCG+f
vC67ptD/8LkwdTpSgKaU8pbdJkpDEVPx6WusyBlB4AUcsjaTBQQwsoMy0DpugBfa
soiP1bsiTLw2riCHwI/UmNtrm71MYkmSgo1J625nHiClssN7wJJNAVLShhCMolLv
Egua7OGEpzubct3f+ij+M6Pa7v3rqgpX36w2ILgaG02MUqd5RFzbXeRmLfk56+9g
X8Oa4wGIOWnYbAzKWK0Wac4EEUg9U3m6+cqakBZLwNprurLpAwtgqTy9OYAQMcOg
qAnfmhYTpdcNUMBzLJzB8TmxkI3dwMxrpvsJwpcEJCPMMy9Mgcv/rpb4qmkSWBm/
sq2JbHyiGtBFr1hOct6arduMPbXG6hOa1HMNeDFpW9TyC9tCx/8oFD3IsprBCGok
pyc424kCL2cFvp1RqCWB7i3FJEr8OHTybTjmVyIxWj4dAUzho2YjK7cqpSXrztgo
T5M+45dzdVCWyTX2wHY4vGYQVoM1Ny4Ir2JGKzpnZAtcD/SXc6JcrpQDa0FCKh2c
GJMUr1kqSO87oEX3Zhfi6nht3PGBKJJ40nyapS3TzkiOutmoQFKHFOvhAeX/7tY3
Ms7WNwHDkiQqYkr9x+8guu3GDVuFXfGGa/s405bd304jAmWsWg4/NwCgUQPQcS7P
pcWz894RVexfoZuYoozOK+pSRNW0HVyqaCw8bjetUe7JsJJ2XdViRj7QdE0mBR5F
jCH2JwAmHcCIvXVAUmdV8KcZhn0HkzSGO3HlgWwxZJa4aMNjAERrt11wQYvt4m1F
2TjwvbkAyCh1q1lTKZTz5GXNzx5GPSUXKVw+5AO2smoCRpsWQJVp7UQIWGjxCk3c
Vh6sgh1JTp8Zsnx95t1YobaloG5MjrlPXFXBFKqqX/5tQ4Kx846uOxdY1lsvabSE
mWcD1l9ROup0NRxycXIboU+W7MmI9ocMJexyd/C9iKzuUujVvV6Yc/GmBOYTFJHF
66Ai3e3cbzw1lx5Hl0goKkqoGzib9F8SZ38Fh1k6FnwoZCWnW+aHnfC3N5Jgi40A
tGNzgrTPi53qdLPYWffSoHBgwQFPs63Pr/+x3ZyZyklEcvj28QGjnD/X80kB0qFI
/JuHz6eYMjkDrCBgg4Ogt0N1kl58XHcbFkkyfhIy571wBu+TXdff1n6BzsxE7Nup
vtL92d8TF1AkNNBnmITZdCBJe6yipPWr4K6FHCgYGZIQVV2AwhdrsoJ1d8huuuO9
3l+OLnmP9QpzZqyrOywgvIqZNSQRYzStnKMMkU4UkttF1Q332I1E/D24+mQoOw26
QqmqTs7hiOs/EDim9TMcnCcOXs+6h/PqACCdxkJXkdhtUqk4s+EtMa6/16ScC6Sc
BarKJJwUTYJUjqCiKAPkxdj5lVftJFD39P4HZAg0sNDYNVSbnhuZ4Vg3taugqaRN
GhAG2dY+L2Pmi3FFyFoFeJbxy3Fy9zr08bfTPDdgxxXtu4VlExzh/SbZT0SCHSkP
QspljVZLKDRcKdQvmvOWTK3w62IHjo7n6ZEg9MlgQAETXDSxeVZeupG5nof3MzCa
gYYp7NwEdFyY4E0bmoGcB9NKCdQSHvJwscIcusePgwVbKOMVxm8Dw++1UJVt6igN
KC+F67kKNOLWh1EkOKhwJP6ObLc7rb2IPb9rbMvuvEehb+MXv2zSHV8Lco7X+ZgS
1nIDBVbzImSqN9lzrClZoc3jJ/gVh6SSD34JwEPX2xMaLwxfJZ6NprSlddO6DO3K
7uJzEgLtvPqLcERVVz0++pWByI7j389c/31IWfkE/lk4Ut/SIWlTBLUq3wRMACFc
pWLobv4fbVWaItD9tuasT99+G5wshMPX5U7rksE/J00GySVcgZR/d33MFCZJQ1BU
J9keYwJfAywOifP4ZYlzbNZgdzpE8PpDoUXcZhnlnWz2cB/j9tvC9sn2yzEtcN0T
gsBbDph/84nJECtLO8kdxUeN1yobjEKLBjCklTwDCjA50SEGkr739wf6KF+pKR46
kNRDO5A0OL3SjqMPywiAtp0qg5fXQkHk4JF6+B7jWyi9n2uTmSsz1pZ8wxhpb3je
WP7eMNl+GE6GwdcboOenXYkIK5XrsIwhUZMrqGPbrI4DpcRRMPGGXSLwSAnMLJ93
K2jsfV7PdFJdvxPtJHoYzjbS9p776Y5NkFHUUBfSHlLrKT2qwSaqVMrU/Jlh2Xc6
EnNgiHMYFOEY4Uta9D0wWQidR8zqfBPEojntWsz7WX8tNGPGyJFhOe0G+A8R1/SL
f2Lt5bgCQVNwdSmHojkEJivhhniGYY6IhR1bmgvzGm2+ECMpymdzDfmtWfDmR5yz
SHBSVNCbXNwdQ3i66wxuqsvqm4hsg9XJ7K39RZYXRH5zG0rDmB/lRuNlA9B9u/4R
MzWcGHv8PDq6UMMw8H4hmZak4zuGo5+I6RQd3OB0gtpiBH60KgMoDZuRTEy4a7Eg
YPbyFwI8qN7VRWtYG9U6teTPNcPJTLbVmhTuWDdQOLVh27BcEGMBnIM4BN5CXxMi
mKJPpyUf3xW4jc+mrPQgCJFWEwEwpvRnbuU38sLGvUxgbKVUgDt8/sMe51Mh0dor
L7o+r6+o3eynlq9wLk28ojpN9A5WL71QW2zKQnvsVCqBX47wCWIwJ3Z54sEZYEZl
nrLeO8fwKJWPiHWeID5w0V05k7hVddWhjaciBu/dWHTfyDxOV1AGgxthUAHs042x
Gy6XMVXqr8K5mTwKqZuT/nRe98m8eyjD5dYTgWoBWfzLi+h+IaI9lIbi3KLS6LY+
0u9au8IfQToIsfqjtnk5O8Cdl/NYm2KttpXWbCSR2ZFPPEvZKk3tEx1VSx4T5Qna
PV44Wkk19J+gffAtVt2GilZZemjLTtl5KdCIdT511xuAY8I19fGVDJUmlMsFe/FB
iPAnMgsBuPhRYsAZvDYRQii7bACY1sfTlSEFz4IoEQEL0JZ1D+WKngJhh9s/Z04l
9sO3j7jKEWUH4YrLcWMqXZxeedstASQCLq9SPXdI4KVuK++G/K6dKeb0SqoBCRJq
rckCXp6EFM/XyWcK2+Foc4je72cIQATdU9IN7QaHG/3XplV0F7dg323VyK0Jnkxs
/gUIODviwHKKterieJbFh8u3iRNRf1232mMzg8jY8qYhWosL5u38yGa7Z41DZ7ET
0Uren04MQ9yhNcc4j1OgNtjIg47OWTz2h77UJ9feMtzeQj/DzzCzMhuS3oeDj0/O
YmfHbnqCoAlLcp30FdXYe/SbjB6d00VApQ++UP1njPy0mS2QfFRm+YD//eJ5YFTd
q5+Un0kL4DnOHTbCYnF0UX29OSerWaIKlgancN1PA5AAr44ndaj+mAazmBDZ3PhT
z12XLTsZXYvrVbYnr+lS8aJ7iXHeun85fg7VqrifFK6AVgj/Ui4OMG11IS8eZy8t
RDdQhQHdWBy8SRcmm0Sq3uYkav7y5TLey1dvJ0BCdpUPDUq7Tq99zvAeAqu1ITQT
eEQCqTE+SHNDjv6gEk58duJVcxwzfVrEeQEcaG2b6XqjrmA8zPdG2iJLViDdoYs4
hm8C4288wESdENsYSXNYgPNtdY9p0nTq3HErdz83pMyOA4Y633HUrCogZrTLQnOz
tlpMv1p7q3cwnqIrovKFBgSfZno1T9SGdZz9D8bu6YfJHPbGJ/E+5DfIr+nMuk25
ddcxT+20QJqUHuDgSkkfMUqRaHfvZa/yDRgsBNCHL+fE1NntbmC9G4x2CJBg8URq
66gcqpVByQsY+0xwZ8VECvEPK1ce3FuuxKlB7ZVht60ad+VTAofUPNk5Lfchj2BG
a0LfgJgireIBocs4CjgwSa3+MnJMlZQkOVAEDNiTwRQCQGYgN24NRL9qfQuboaVs
GaZ1sfodRcKVq0MG/rOLy9Fx43V7iqbN+bXc3f1flj8TFreTmnIVt5yQWJvkeKHQ
fK1YZYjRfdL4IVxy6WodXv7qtPDiIUzN3uYk53U6sySuBhfvxGNS2nfZdiC3d1IJ
UimdIKyoUhIUcL2Wi0SlUDgpEA+7d/Hn/fGjZGoi89zPZ1b6UleAnkwHzjav1Fl3
UbMhwA3i22nxjBKjRyEHqChYGoDIdsKYi8lBqPGMc10/+O81yfpV95prul13OFmb
OKfPvoditXNI4O0rv8Rt2fM19TmhISMHN5BjDTrTFvnmlYPmRM1R0ekcJ2GU1bI0
6kow4+2Dcx5ndMiWnD3WOu5+7HylNfn1actw6baNCWgUugK4Efs4extINNVZxCq5
36tB9NkqQKsAaxjmMBMSpONps7scnSeDlDV+UqkTYqPwoHFlAoWxxURQ9eRNIHdE
bLPcMdhiJwyJwFmZYcwxaIB1jLkie9aRdpGujcgr8l36JCMpfowmW+4ruxovSMLk
tRVHBiySd38twToWRC//rtZNcu7QFOWQUkEU/ZejiEX3kMHTkYoGPaoBfQagGESn
HxQw5GXmeGbSxuDA4+daZlycpfcQfzOhjU7maMTtxZbXiA7bPC5WCAKb3g95yz//
2H5SIrZ358E2vRX+OeLmbgNyYt+YX9MioP6PC95q8i62u4T9mAiOeUu1k00460dZ
HUpwpYr3Rp+ercGdS91JJTvUfslTeEFZc/YglRypnNlRU2+20+TNlQyc3RK0Ogmp
ECAmgjbKLrVOBbc5MSC916rAFajz6PjapjFacTDXwZk+eSo2n+Eg39cKdtcyeFEV
+qf3iVBzY88sGIws2uFuEaQxjM6Okv+dd9cb7ilRXUEb81WO0g5xFEruVUnBoRX1
m9Y04kgMRmISlEobiSH/2T+D5xClqiJA9GFLX5X9os5SrJkAYVaZ7qLu6Wtgr0Zl
OOSD2kbtnAi/0jy+K35taVQo532Rb1LWqGMV72xUBnyLJyznGGK658k2dMxy76d/
Qxr6wSSDQhfO1R9SJko64jQEAsIBYjY3uJCQIMTqN0WoEzXS96Y4mx4it66pCjm/
KlLaaHVPWazFvVhfqEHDoh6o5s+CpcGgs9T1nz+8sJ3n4jFY/1heC5O1yDGww2MI
thDJGxeXhPKJH3nRW4rCLJFVjFk3ctxY4h6bJFH1DgJy4XwvyurIYkvxcg9pvBgq
IQC++/LZAgcJWOkIbihwZ/Qk8lrr9pazbjygD5bgeAOa9tY8e79s2ugmCnxWO5Y4
EOHXS9N4ayEfQAs7SnD+fsM67XDoYzj5om6Yl5skObal8TS5Nx+P+zc9Zl0W1Rrv
fa57CG1gl2x1sKlEL4/H7FEzK9Bnpjg2rw4d7KVCqmipGKJ6qom1fVo2+afe0S9v
Q4vcbSTcmt7/A52Ep/u/xZWUPooGTZMJNU4su3scSEniNJLT51OKgRtYKyoIVzI8
UtUAGd7roqogL3uD2+20PTCt3IMveBc9RTG91HceG1FXe/jkHxvMvYxmyCRrNMcG
r9TIxkUdtzg1F4uCK65S/AykkroC2P0zfzjCVCviQj1t67GTiUyExmN3gCdGAd60
59vLvdjBnN2hhYFPaCPCwtpF9KIZToXdakCppjkmZThwk0ZctSCw0Bj36PBTwwbH
mUoAooP0sMud6t2pAukrX73kvYCgdOob20AFyXLrbBP8z27ULWPyB55iwx3Q+IMS
khmkXL5ZMMszcdQ9w+egI3wkJBUOtkNKTkIE/Dj/mmvX4ie7iMkyjVl/2W8dQvBJ
YwbZCVYJHyZ2/RpzCiw8AulFHLhJTtqRLdA5m5YqIuveL/Yzv0BzIHUQZUV63cIT
9kIfTRoSF9oNGPMwxpunjO2qCxbWMsljgrx5et7iO3ktbBN6tfPK4w+Ofm8MZIwA
AGqXBOHp94VjjPqFHOyQGnWrWCphhK/HYYG2gy5JGf0F1+TYpJkP9l4AjX+cNM9w
aWRBzRZGx49QD84+7rXRN30hTQtyY6DJhTabXyHMvflUbydQerPTYAZYBXPO1DtG
8G0gGU8u8jN6ZpvnHSWukcQ7+loWRf4f3V6NoFbPFHq/ZmcxFjlEGYKud59wgJfo
t78qGvNGjOOJu6pYJ7MdIxL1/EEsXwjSXTgPc+Ct/7GgviN2Ftr95tWlz0BXk/Tr
OJ1uwxRzRtd7LwMtWJaVKWZlR3q8w7ti5jXZN5bjXZYhc3YTYjO+VZH10Ify8vah
GHH2cZRfOOHgtNwB3E/k9DlXwx+t/jP3DPiug3yh9m37lR2deRUpBfV7dM8i3jqw
SDmex6yjQTkkPTMSq+Zy1mxVWUbfsJEhzMA5Ybohkopuo+pHY0foFMcvkuJZpyGN
lc6vYbEpoB6D0hbmixjFtBqcOIGmruQGo/YdkvF8xCSk9TJg7XbtHSAPcPMwoJil
dXDPrIoUxam/FESfMh5vzhCgN9FARlPcupGlHXManHsQS3yiQyjZH3WGIDoShJI2
xcOq0FZbmaTZGWSwIDHxj6YDlOWOSWM5dDlZvDg1kssaLdGzGATG3aVmaljHzRmE
eqJJrM+vYIrge/f9lYjZPRqCGLwSh7OEpZdVnalMcTBHk7fXLiA5bShqOtPaIUIc
/rUUuOfBjqCHf6n+FAqZAeJNGt7x/emzHtAek+6CVulnTBkWAPxUWXWqbm6GpWmb
4PTep7XSLP0A2Um9Y4+d3iAnEixWBiMar4mTe7vzICntzVSIMCJgq4A7PEquholy
yMB8dv/o0bCGkg9q2mHTVi19vjCT0i/awp/43Rwt+cslGDHppdpgH7uqklEfQ/Kq
0/WNuxjcugHYPwBQEztoYa9EB9XygsZ9Ua5yLoPxcxxLz4ETUIq1JmxHJk1bnslH
i2/ZhVUnE+oN8LA/ESZszCuaayRFVHdZflY25V8WVNaL8Mn6JaiZFdZ9wm7VAc03
DfaS75mdOHo5lqrixHPCvMVm15cUDVPj2DzPEuYD85JhOISCyA+lV3zOUoUUYp0x
FZ4uhjq5UepFsZ0bFNXDM0DdlvBFTeRzuG1+SMGgGAVN/RIOlOZTHX2WGofFAOUB
n9cbrS14Ci7NNioUcvnfcnMmcrBz0TdxP3bIZjhyfGsaGYrrT41CfIiSs8ZCeV/T
dmGFVB8GvO1/Bcr47fTvyLyy4TDqCS49bDbyROzHeSJsSGUaBk3I5pYVwHL+EpNp
6Hm1Xl97fON/+XykpoEXCfGUC2cTBW52jg2FdqInem/sjqcmyRkRDHWkhRV2n8UA
DNfUi/WMEQYK3I9aFu9jfyDzMMH7KsVlQKfaCv0PgDADFQm0GFeRtlpd7eeDJfRQ
yns7IqWlJx2HzITh9OhWUaUy7f7WUVDyJRef6TPWY/Zb63c9NMRmfUGPcBmWaI7z
d5lQLH41O8SFpEL/B3PLmrUFsTQX4/5h9s0tA/Q6wiLlilIXKbPpuPwgkiUyGJkl
X9XRcKuCbjUEtrjR15N+qKoUNFBubp181Nc+RTsmbM8e/PmyYzYPvLADst+fKKQT
pCl6zs9F7P6a/V06fqM3zWCPLGjUqTg3TcPBDqAlP8m+v+RfkYNhEtf5II/qdeKT
cq2fYnsWVh9lUmD5hQPR4croQLNkrYkdKdtWVEOLTtO1ZDoB5rO9mJFI+P3PPonT
Ccp/+seCOzFc/stQivJADG53+qsusVAHi5JyC1Ny8w93XOVOGSWjxJT3TCT1TrY+
jUrHpPrxEMc4RC8jdTZyCMYty4vuKsKh7PkUwb076E+ssDarE48fhB6acNma4o+L
m2VfzoghPqpYiwX2WuUU2Pguy8pqR4HJFqTZdqqKqILv78DNmPvGwsxI5TaeinXw
1g54eEjgIvVd5qYG4nsjL3GNXXRSB/qMPUnZop8P1wXBmHddN08Yhlq8op7Diej9
toRxghY549hpPAxpydOrS6JiiyZHpsekR/Ijw8FeGK1TivSB+6IV4zZbvatnBc6r
J1XkFsJY/NE47GuG31FOvpZRNOEcbqegHnB4ejSF14OzEvDTppt8YPZh/5ni56lI
mfviZqa1ghB5O8EvXxJ7IDr2m6i7xH04CQ6dkaHDGoxDcQGbGazAe+2eEXAvbJnu
M73cGflzYlfUABIXHemyPzFROC80RsReVlJfZwoYelcQNlwZ4ZeeyazxIhNgcMZH
najNquYcTddKWiRVDwrbRLmxiG7y7dvC0Bk9oLY5r0sV0neFnGKwTPb4LOFgyukB
aRrXw9fNQn8ww+UjpG8TCq5I2qvxt4tNORLalIeQ+oIPecqQI2Hz4m+4gAAAMDJ5
SvXHIKGiUypDBBJYRy39uLmkaA5vyhuFasXdmBwLAc6Bb+LWamE5vw95c2mXwMCy
t2o2xVErIDnbyGhZ1F1LGPg2LCZMxHA2KCQv0DvSh7MJDjVdFLKqJLFbhrS3fgra
xE+H2PyGM8oq8aCMQt3Pe1fDI1HMTaKJN4gXlYKkkbcYEbtBEQ+tw7IKLg7Mp7ZD
mo2Vud8Hj5rD2HYjn87O+alzVPDkpJ11mMUeB8AabLPjQQCfX+TLA2qjPkc3+Try
/B5DUPO5WisVHJMsGLMz7JvIYLcZOSE+32ObHUrHP30TZcTdvt8Vlgp+i7TU0vKX
jorwA7as3CGcxah9wiSHOWhmpZP/UNrEf9TlEY4Xhr3laLLnNjU72AdT7QEScQSW
YjpTOp8NY7YnGzF1LxTVHf/LbBA/PDp8vtIsAT7rEWSeRZiKCzXYbwLlQIECHyGR
2ARiZJzU05boG5E2HelJceqSHAzXNW/wQ40a34xl8v5c8KaipyJ3iEEQStwQaT7/
FXFlyYjCHOheVcAmZzGPEmf7+ftyJh15VPR9sj/xnDy3F0Qt4KPmFRcnu5QfXRhR
GlyrpaQzf2cKYQhT7jE1nnCXo4p4Hinpg+0GuDWADFrBr/eWpHSTLi5eR4OhU7dq
48N7aGWE45pxSJEcNDHrRnaMwGUguQ5OA2hRo++31tUoWrN8V2+tn6ufrLGXh46D
Tl7x7BObQ5CGp08WKdqQ/O+3Cs+y2hR4sI7J4K1EvBuRdT0YbpWuJ4uWxrfE4ZX1
vo8eft+++I9JaeFL+Pkir72EIRgs7z1RnDBo4u9LOoH6OuV3wmpIF9OZsL6VJH6M
oB1cwWmBdMuD0BjKdLkIbTI+gJ11+Y57gJuo+yFKjMeSTKE07wYSxP8MZUwyF181
EMMzpzeNd73JkBGYglSJDYQwFoIKdHqruwTNhWNh5QVrRHB91GfcFdAhLS/s4Z2R
oQtunJ6Wb9BNzUatku4Q3c6HLYN2Y2qW/nnZnVPJxqMPKpYxJvP5JL50IWOw12a/
20bh9EEKGe3KXFl3S9tdQGiST4YahHbuMyl2XlKaKLSlU+GARed7gZIz3LJEpItO
4ZqOPFNURxSamZcVFJh81ZGo0WZhThaMcMde9Rtpwhl3uTrsKNbMA5sU2N6Ia0PI
48dZ1/Eezhmwo+J/oYHqQjp2+zOARS10oEq15LWBJVZy51RfAE7plx4Tqi0XLYt5
H4RxDSEeMz5d273AxloIhJ+vIOoETz92f6tOhbXBbzXonPBd+9YAow2eMbiy1opt
ECo9wDZCrLR5BZ7zzd+gX6BmjOttNn6yfnsPv1hlI4gywkGe/K3QnhO1Lbh+GHnW
lmigjs2c22ULjulTzof8vJkb2Ha3lsn1WiFYDBA8UHG4K/NGJoulUFtXQWFCTX8J
fQCbTxp9YWoH/QBgfN/sPlI6xwdwoA/aB6IYl4wDgotguiL9pBLQPtxehkGf3qGX
OieJUhOHFqQg2uHF4uPhSxa8IHmxqozNRym0mUC6HYCBwY1ApqcIicq0ywI+cnN5
6976cpsFu30y9Fza9/tXQUPfxIKwC5kC7QCrgmN0ikQsp89h1vY1rRPeXOFY2pW8
23DdznQrHcT3fcxH4RqywixtymMqGr3/MVn2J864O8wATOdiG/HAhuolIBHOL2HQ
CRvOFjBPYd3nQKt141UyoJ1FYudOOltpPO/ln7VC51Xa+ljOTWqOWUIFNwYhoOEu
ELEGLeNlHo8APmnq2VB9/icmG2UFHEapoLLYfJWtY5ZKxgD/oExJ+NeQSMgyAq/2
fba4GUWlrjNUF8lsyPmqKOr2/6kl0TEXWO/Zn22b6iZKM7Hb3em2SK45OLTDPgMj
H52+/w5kGdXAM2gnZPRK8SUzFmCY33BIWuu7Qd17xTjeM8SLXBHw4xI43P5kQ+Fx
CYgQ3XW/e1/oEoA0rUVwT2hCCbxd74sxCqbIse9m3JWiuW0nMl7KSuYWO4856vML
N6h3mZuP38RJqHk8O80QYW3QK5907gYkRNBZ3xFgtVk3JiDWCZug+WU/evpZSIef
/c+0dxSdf1d6EVOdktr+lAob1+lQYH14EWGOlb9nllNOTyGnts4g8o0RVHKXFw11
r1BjeotNN6myvau/1An5qp1439n/J1LFCsf2YJG9PNpQP4dpJSJV+HYOFe9Wtlxc
HvsbPCbZ/tFrFspLcv9hb0ph2+4kqTrSndoTIrZjvHusNQb5rBCttbw9kev43mnP
997aYKGo3d0y7qYZu+2s4QwLvsBgjXWwib3DaREJkBD8ff0V80uCqDvieWd/lDtk
x4RsSk8waFE/t0zidHxsaX2Ek9b7Rsx/OfULG7jL9euaEF/PMZps8xPNcoPU7a65
KmrUtUFxYz3LyrA1HQmnDZYkHUVavIKzTklWmhYAZL90p6o7eixJTQsIJckLXIew
A76JxJ3mjoE2jfF+StvIvV3UriHqk5y2wDFzANMwuEvPzSXAV3S7s2OL6G0h7AX8
ZL/xT9joU9EAms92nJkgxPYxuFDvshfnhBtnhvwBGdemvGiVD0wQcdqp8KQm2wsa
JLgW2A5XUaPr0msVg73T0etFj1xeJjyfD6fJMymHpsm5N4OHbwi9nLjL54Pkjz0s
wzzQD5/FixkOpB9EY0I7D3WJCYYcuVSFlUyDhdSeykGyd6ElwhKkE58ZjKHvGBvI
8+dUsYOsN5apDa8ZcXysajpne4qpmcjJk6CnfH7hUSG+Fihdl1o0geFYOle5P8ej
VBUnYjk4gj3bFcQxn7aNElKKW9TxeULuNlLmywOOa3qPYijc57t6qjV7cbaK0xtA
MmGUJSYUwmAZlr62mffYF8aDblN2pbJ/tstW3qNvcAh6Mwvbyp6KFaitXO8JO1R6
/9CbdDnJSi+lS/AUlTGRlbh5/D8SV07DxP+ZhNZ0sb+UTOLZRmstuCNmu5boZ2xx
5egZNOyOn3IY+UK94/oN8l/HOXfMBXaBrHdej7g8ber7UDTDyKMUHjYgajeGjb4W
UxubRjMD6a4C1WexMbtOK+UI7AZyqTRzF9rCh9qUOkzmZyTRTx8FGETcA5Vz8/7f
geSAaogE0jPGCzeg/OAUyq99KVcePfX7og08udm4XMEMjDUYOBSOxskbRLb5AgaM
Nrq8bXMeD1bwa8665E+NXlB4sR9zo2Kn+azEwAJNRA9+9DWTLNGpXwhVkyVTdH+Z
b9CX6eNuLrgehH0zHizIFMO3+s4hw9sEi9y395gN5G2UqZiDh/0oWx91oisTEY3N
P8T/Z0D1WQJXNB/IXmkPM5emR2Rcl3BmV/XVN/b/PDkAUUYQco4KlZL+nUvlTokp
owk6zUp6Bl6dM+0cQdTJdTEUrOafzkffaV4LgzKk+QK3Fj2h/d3khndC2wQoTlmx
b+Fdbu8OORXy5o/K4Htbdp1MHrNqTy5TeEJ2UEj7RUYyCb6LdN1NkFQ+vB7Bhm1I
DGaAIBxMleAOdKW6VwiBG7hjYKp82v+bpa6KC+8znX0CbnArMabfXwblMhgXSapI
AXZerRePUqUAjxF4etskU0sq9Iq5i6SgWd3tT60rRT/zjb3eW86g3y4GXALg3E3N
ls46SvaeMD+3Vy4/1Ski1ViAKTRxuJl35f/qR8m7kMo+B5d29dgi0+ITlNVqXe0M
AISASTZ7iPNEMeIWpGy3Y9JbuzXUyEOZECErxA3xnjJSQfuv6MgLIsnHNLMAnrlK
FRcHNA4TECpywDw5KxV/ldHhMEKnHUFsy2SkGOWssLjHjAQtGAgHUzJZSR6YmXrm
EwtLuy3M9RgPpDTistbAXTtHzlxpG+lj19YadQWGDg8NRjb2q9jqFwUauYUPp8Xh
ihl9+h4FSR47E0081olGSF0fn3voKCHzepsYGc77CLGbUHOTIT5t2jOfP6wf4p7Q
Q6c9W+9hkuurjMHBFkRoA9ryQuJRt0ljQDV3Gq4XU9hUFKGPIziz2eR3MxS+wf0r
qq70dlr/r/JD8fc4G7Eyu4ctZ8yOFQlubA7Aw8wEprLj2SvJ6Mly8qwYVf9LeXPE
yz9YlSoBZAqjliUkUpjIvEHKXNRJMC4SnO7Jf1mwnTjkVJzS1d/gaZfmwMkjvUnq
Zv5Yt9LFQ2J61miG9PxE/ksOJQVelUu6GzGepF5lsMd1+qrC60EEZ3F5YdMPOp/q
ls4kwvx+5OKveDBnmdxw1UlaSmp5c4nb5dv+mStkiCS6IPKH9HNu/Wtiz2tDjiFd
YICOCalOI5U2HWEQnLfsy1rY2nPMUOINl5NID9Fo1sADHJn4FP3kUqcpq444jWNL
iQ0Kya2C2Tfs2tGIvxGywrzvarlIgkkTVgv/i901CqMXI2lKuG35041dFTtdn/9f
gPkxLcLi8BMoHdHib3g/BAMcwZfbNYo25kPA7MGxx48d93Y6Cz70P56Z3vmihesU
yiaMeCcUwU/nT9H5YSNelcdeA+VeYRcCl8s0ld7QCQD+UUCB9yEAeZRXAv3r5VH0
hnMvA1PL5zlJaa3ovviwpCPXs35PGXG6w0VtnWxHzzD28NcNwpwcyllYnP7rmLXP
LtkV43ziC3z3KJV+XaKzCUdE5TQFXkjuh4h0G7oujHd/+K3coz4cWZctXJp2cjHc
NqrVfCkH4BLBRS4cLSafoFJyMyHsIrinmrpPyv3X6Ueb7A7rJBR2Naq8PzhqwCQd
M/z/vw6ibIYE83VyfDA+WqKWE+oPjy/wLM4NL5A0C1BA2dY28OFhh4LFe4d5+kpo
Kc8/wuzL9Ro/cGs/LfG5YniRJGfxUy+4aRQtumyt5ilZ5hPtcYSh/z0qfOzJ7ndE
+7tH4pIzUW5HjjUOLmwH1pHBmmYLdlyzPWksj2avMJBvoHnpLuu6RIu2WB25lzN4
TTIByyfYl/R/PF/LgbHXar+htWu/MXVzkSL3tIEonkcvBD3JbnEOsfFlov7BhZCh
K2fLA/8X+e0uQ0oPm6dtK62JKKWWir748Dw88ABB+2XQrSa8+eQ+uM20ZuPDm+UI
755IdW3ROWRCkHwK8//qRKkiSEMYLVRZwnTlI8HgSXbgsjxE7mMLrXtTf1VVrWni
X38a0zac50fwHriVEnG2vgk51455B/D2tm3UoBV1z3zgQKBP71MpITJ97wX9Kz1s
OtB4+7Apmjr0oVHfvI1TEntf08Q0zBgScinUIYH5PBKjNbahwYfPWjWm2qSEni8F
dX+oV3+OSxjKa/6mOMbnXAw2Jq/XCGyRY1T6DvSobi7p5V12XlC3DuAmJUHRHOTY
kQN7SSRWSLAM281Ot9CnJ+FgArx3PyCt799tO+UQu1xPlnTtrnZBCySlAS3N0R3S
ktcKR0R/huuKfHYmQ9q2diPbQ2VjFoG+kZjZ0lCj7G/wYbN/yTjGK8gKCQKWcmKL
LwDZfDuBpfyRIiTyB/iPQ+yQcIrT/W17YpgJEw7gmqaQ3pacWIb/IzOrclB+SHqE
L/LfL/qTJq+yHh529JWO3JRXUJOLA31X/Hi0lqZb3n6UepT3O+5MvQWcAT0bDYqp
hurugccjU6/bmjVQvOqfgw+SZr8VduggYbkDea9VQXWDOzC3NsohTd8nRcGTNea+
tmUkexjHDOOcq5oHy0/UETJJTirCffXeV7vPNXT3i1A340lLj1Vt0M+Dtg7uuhYf
NTzoUbjss305Y5SbNUj9kS2LaTXpcE25mCxSg3ih/ieoMGaxiiHJSGkzdCLHZTN6
imqw5EtXeR4qdclpwTF+gRybGRtUaywYCFmhRCyhI8ixPYdL2gNgjI6v4Ayiib6r
61JLWvmimnEPaHXHLiZzZdAdqunTHK87+XbVRJpyZerK2XYYCHaaq33WTQiZkhlP
lL7rkwvBTVYeLgpG7YUC4n2ZZP9P9b9dEeMhlQ2YhdemHeN47+U/Q4bdo+KWaw2B
WLVOSKqTkKo1FlBPg/a74dqnK91EJjGjGOzKwjyIkIya1zXvIbyUze+WW9yEQl/y
ziDWyKRGtDdjaBqZd8uV29Y9QrQlK7F9Iv11RX+Aixt/gTWijK5rQpk7dIIPdnCN
qV0Q7NiDvaHNBWFo+qNDufHOZSpu0K2+K2kTrC3x2WP07mE/PnTM/39B9Toudc+m
UG0aMYqr5xFriokqA6DN9GGtfkymJA9fllWIG6pJxXNtXHl9NByYzznx3PZ2LKl5
1nU9HIIag29lAsNdRRVsvOlsRIAzY8/XRwsCXxGQYC861Won0Nbgog8AXTfF9kSr
XrE41iDoAOJd2vWxBpPJW5l+OR82DLxRo6RN7jvvM28glU6Gui044EhsauGMctwL
yH8DRSrT5VbXgdvAUV9T12XG30I8rCBTIsUeWkUrpZH1nObfHkixFUyT78qUJ0HF
tv+zXUEmeIrTKiNNjG7UDWUnPyPKB3DBaIBbqAgSfSLr4BWB9kvUJSDqhOnwvJyH
aX5WpfLG7SQtlliA3wMVHYPpwsPQDrDKRXNtCkzIhmcQOQux8bl2eYqiNLE4IcqO
RQw17L5PPPtFO8tP6eMvpdoY3PP0vhBJ4xOWA6j2phxhwpo2nn12btEe92XSo3Yx
D9c4ujyJEj3SwCtmmVH661yB4p1XHS8T8v8ny/Gec/GBWbd9RMgtV15OE9Y5uFGu
VFwSwwx7ybLIUPDMxfNOg9bpNDbE1ovpYsz8aSjxH+cbc0ZPAK5bmVppuam2dolP
NJrwKrMvlZGpgTBB2n7ypxry4NUBYMST6zrj9CS2640uoyVrRCdbvl2G+SGso9P7
IrDOiZVDtZUH+g0yxAMR7a4OQKyjuEdVlZYRmA2vS4fO74+kIqst/vVe0psn7zj8
/7XNf7AtJ58a9IsY+0L8lK1dE9jbYSrC3xlQXhJeCOynYOMoFZMOscHUyX63af7G
zTQVaKC0cAEOq7Bn5lnAPNB4SvJzX2zloV4Hlopi+QPnH+uXIft8sXyPJ+H4YIH+
4M5U9aZrbIl+L76rUVw0lQlEfLcTSfm2PiZ/6eQ2TublK4UzB2dAEzedChTS5IPB
cWjtKesNkSGcUyhkKVjxL7xqSWeUGxgtz8N0sEChk8wZrGY4fiFpNZXahc4Mp09n
pbUQ6YBvcYse+fKPRGYwlcBbuHN4Un3fgbJKhE8qVrYRRh/6jS+qDkIKANRy7OQK
U/2/0+ncxdLqzRn0EZHTfuXg9tYB2/0IYv78/VAVwKOKcNAhrsN7t6w5t9IsM/vF
FI7mvoYGG97gcowDQG7Kfg/1LRcPI/UnkNjbP0qXdzPO9pUTHgC4ZKe6fcPqjieQ
tY+LowrWEjYQnwj0skwZ2a1wACuRb4wViNaRL7QswjLjJNfjEly9ogF4jFfRuXfR
kpPANmVJU+rXTAVS8NJvlVNQh4FK3/vLmGXSGGT1zIL5tXXYdJoJZdJMWSWsk7Zn
oUHrZeHRi9LWU6azC7XwHP+WILn5qH8uhdg4SyH9H5tH7mMW9I3HOB9HOWFOhD9/
XxdD4Fjv3YqBk1+2/KNjg1C7bhPvRGckRjZq/xInfgVpCLqXDRpUlNS0W2lTenMx
cdv+nqsTbGNJKdi8KYSljrNkq0ElY86ANjUQRSw2FbdQDxTnGkmleoOEf54iF3wn
XzatOddg1c8mYChmNUW3oky2rR4Vn1dPB5pVkgZeqJqmd3pwdBfF7P9GpCkaO6pB
KG8HkBST6THTpuwyJRSAm4LUa0xaAxOB3IQv9/6lel/zePPISTQgI8tJ+Tp1jJFc
YY5CmWXSS/VxgoZWx1XtG6l/hHS7XbDHcrQdB/pvqr/IaUtOKSu42ieNULlB8/Ys
fx1ApEvFcJXEQwQWBA084YcPFFf6Cvtc4CNVNcnfKVhg1/wtqRoFBHUsVRsuKHxW
5VhMgzz4NSEthvnG8vppJM/oZ3sYlVttOn/GfRR1ImQdyT2xkEwvT1W+lbEVEmuo
JUhcBM51WyNnZCI0EYiHVA3A+GfJ8B9MkbjqhgdPQ9Bjl1ykweHGR19h7IuRUXCb
Rr2w/0mk3bMYalLBRH63G8GtaY5mMaVKSW4qzxT5pxnam/0tJM2QYLVOUa8+XcPk
M8h7+wiBBXQyvgEEHIxyuQ==
`pragma protect end_protected
