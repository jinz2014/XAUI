// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dqc8VJxBLTD79qaKqZeCD9liuWGCr5oM5KDMHZt6/7Sr8eT85HDktgVkXLmI7cXd
thLBBVcg9ZB0oiwUNFFnfXcK/jZoqyOt/iZPliRcUDnH3PoPO9BZj7ZWAvVeQOWP
alq/+Pkd3f9VqnpaL+VzgdyIWBbnDIbDVKyUU6rLEs0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28304)
bMJLmpz7mkM0CiQt8VE4et8cTdzmfqOx4Wvcyw+3RF0E6KiFFjHUjTH9BW04EKBD
N+y87GUbL9ClnPyYj19GSc7lNgax/m3ICueukTIz07Pze3IVi/esswoyR6/+eg2i
dzROjg/7flljJGSuSOMwWicONPi9tqip5o82854egCs9TXl60PRyBn8sf9b3WMpY
GFA98jSaY0MZtwwAdP7OLekRVrdkKGi3epmwpJDjvl5sBUEcGc2duHuRLFmzzxst
tVNIZEX/4K+6IB8d5C2x6kqtV1AlzQxLfD1ULu5aobPIIBaqWRsMf0KKpL1+HouG
rm4Mxulmn6WspiEfZBvjAkv/3yOXBxw3rQ0EpaaJczvp9LYoyTyfZWQXTDmzXwjC
GWfhkk4FcnZKagWAgIXpWxfWZXsdY8uecrBouRiGsAW9RNoE1MenvQRs485mS8vE
c34OweUrVHMAr9RyOT0yoymXYyDt0zAmFPB0pYdAWlo9v0h/ZqnmBMuFFEzrhdwO
I0VExcUsDH1kxn69nQn/j02Nn9YVkZBz1SWQX8+rg+HnnB/PTs29ARjduNOWsAW9
Nxxr4GeuwlMFfJkqQopqKi3t2vzBMB3OUDqo+/8I2oQacrmZ4njW5KIb3WjN80x6
fpq2odjWlgd7FIE3zjIRG6AzisYGDT1leSYpc7jxJDsgFF6trO6Hx93Xs9M0GQVX
USlsrjxl/h6ptO44CMWgkCArV3hyRTMgfMoYOoJSYfia1UQTzXn4tJlX2IU6euug
OVIZDnpKyksO/eLN5Ci9veWKQWpzTIZ/YKWQKb6dcYVniXrjLMUfX6wdUGL7zXRo
g+AgLsVqASMy+fBloPEsK/GSE+x1c/IvBQT5Nvy8QwFt31XMh51THBDo9lrqGgw2
vDEsHot45gY7iW5myHllYr3lCxfWMqh/M86c7dGO9ZXPXW0tR42HPXYj7mhY/j8Z
QxKaQZtNAj29tfPtV/2tdEvQsM1IsUaCjN3ZtA+sb/vNomNRMrxfi5ku3KevX7dg
muYRP4zZutOrG587C5lJXQh8dxXbhhVTJzKOwOGIyNaxeqceP80ICnkYGfWt5O8O
ZCmQoDzEVDsqMEJMpNKhJUswv8pOKmxc+a0pfGTvLZLK5wK3c1iDzTyhitGqtsBT
p59Ld1QiMa750VTYLq6Tmi9u4HR7dm4FVLWBmLkVnKylsJzxygu1d5IpDL2TcLsP
9LDaizA2WI2I2bOp8gpJYq66VpW8prqbL4NAMI7ciL99kXAy5va9Bkwmf+HfqCpP
Tys8UKBdQg5fTv6cd/XUfiUNCqwuPFeclZZKHQM21A81SrR9MaEG4fv7bZCtI+aK
zocQCTZ8ii9rn04hRxXfi7XFvMZBH5ltyGyv9pe8lNg425kCDCrZWzctdOv5Rc8Z
MVJQMha8b4Ql1h88sUIzQcNp7vM6QvqVc0Yz7vhXeEDWunsP6rfNOwdN8tihej4Y
cs8lWbUiK7rCI0rShSd+gnH9xhqtaKfFg8xWtAUq0wWvFWbc3i7uBS1d5qEoylUV
heKlorldl4akFSMcQCTm9VjvYXnN7Og1nghE+i3OB+2Z30CCDE5PrZAS2bwlZSQL
iXJZTwzgTvObEeNBnYUcDV0QP7ekaUKks31ONW+AmSYNNA1IHSlscGdyOvs5BZhg
hp6vV2PUrLxbrP6IgDMfdUcwX3n0Lc3EXLEO+tVhJvG3sPY+9bbFXcxbHwhIBMcV
7GfKkp/ngYQQa49/gh+y/iFPHj6Tef2vKbBTt+QY9vEepNjebu3fDAWpAWvIj0Tv
wQkwfvXGtD3HdvBw2uTMnzUIKVOtPoeU5VA0a5U7wYtnCX5x7BrgHuGqIGA4AVgV
WNZg7zaeQiM/DA9vVx6oR9C1hjs/QgCCJGDDStvWOjkA22Ibv9hZQpLzEDDVOpFz
ab5Ib2ax2SfjjpqbjgGWt1p1FttJfiCDuh4smfF1GEqHc0nIYvetjLHJPSnDePNQ
k+Nwi1l9VYubvq7TxFJ40i4/BTXRyaSTWZOpOHl9axyA6dSTvta2x2xIRSFlN0Cb
NEdFefZaYGqYaH4DulHka3vF2Im5gAFTVYttGY3YEecy61UkzzOxz4r9Tja0ig0i
nbkH4w1YGDlU/VL9jyko4a8TVCaEMq370ztJCsvk19Vt6z8DvD8zxUtbsWHpuRrC
IXCmnUwMkriZBHfhNooPN+Bq9t3KGcXNNDhb1eDBY+8AZHPPDUzK2Ra304a1POZM
DHd5XEEHv8M9XW8szob5h0IAFyknlIK3IVz8anBz4cBqrvU8CzkbrFLG/jpWNwa9
CCDMv5Sejjg9vU3XJDEBwdqwRn4Cp9P7OKRtx7AE6qLNRJ1/sGX2HJ5jMHK3xXOd
dkv6kcMZgeFz/fmICb6whyMPIIaRu8IgmG2bWIvor560FjkrrJzvxVD4EnPAndvE
QjWEMYLJs9zDB+Uw9J4fYXWcy/NeL1oBD6yM/Ltq52PqCCi29ZTUXoSvzD/DhwyZ
+Euq6CO4O6AD3bryw5HztPoqkHp7UxGeOpqUfyBF9CKqUtJIFneCkfq0HiEQ6fZU
H5GxRlDlMVoIHg+3rEwUpIbAOQdN5yBPdpJaneHF1MFTvgllh548pOJ5bC8CRei+
h0oA9GUNGGfSXLrA/v5A/8DaEUY8b+t1vZpyf4e+2eWqkh5BgYcOpWxk9C/CY2H7
RFOUXUcBL6gPMV/r2ZTh3Ga+3iVna7jeCtfY8GNcQzr20woOunCk20vBEdx3a+LS
RFLeygK0HfbMeq78LDTE0D1pDRvVObW0Ut256bb/L4cOgE5//PmBWTVWyVptFocx
57GSpcADUosE/fIBhHWOFo8zbz4q10wbD8hcykzaxOJGjzeAduYDuY9Chs7lScwN
ET+TH1DVwymWyN7y9Xn/Orm/5TG+5vR7fXpqLfKq5zfkaiWK42IHxg9vzxuhbq4P
UR5dCd8MQI52qc95kjMKXlY6uQFM48eTVKW02hbTR/JPcBzUdC18fBDEEPPFtDGI
4ArVzd2125128Obw38dr4aOPAawWXscFXTXN5gSXnmqs4seYqmBBiuGUDJ7fiW5B
s/iCfnjhdyyKi6aJVjHbIzk3erZTcAg43IqLHQZ0vnipQWCwd+pBNtbQ7JqIWAuw
1V9H6HcJwp7FloR4bGSw6LyTyOkphwaPsjxCYql/BU2JOAsxAx0BLwdP1ieCC864
K5T0nHunr9aNUvLg3jZdF/LOVyYA3RCPnETHlvUgggYRA6syNwGd4MaBe7ZALBzf
yXc7RGLI8qpC6hmflEuXjjgTnL0q/w/JqjS4gaR5wxgm1gQG23Ejlun3pEK4rfMH
jov2UTio66n/2wOJtMNMGGTsHcfLGewB02pY1PoY7ocvvd0p+Bndd3AnTqcTCOGi
apVV6XWOjr8k4oq+Ta1x0PbWv3VeR0ZFiPqov1j5sdGacTcF4zPqh0abXn4ZXX32
pGSW1Q37Iqd2EcaeZBp4Z9OcCrGm9jp60Ku5gqzn6UxLerG80Sy05CHCgTDE4cpK
EUBxuUHMqgq2yHIgbKzCsEWU4a3V84oox5pywScE/L8RugRh07OJqMUBYECkVmsd
sUnmMWLJHXuUr0ukuEdcakWTdGDbDBjdJMv1lUL6W1HGFKzbK7j8BrkE18yBrPLC
ULyhFjU8b/3a6xIU8pkW1GoiZD1FKllsYiOUcWdUg0owGLtABixObGnk8bsQ8YTM
vMvC3SjcTxM7i3gilLBI7dwJEyxGyNauy8gGDACx1J9MuckbFiBEiXTqnGwZ7MvI
g7+DMVdbbvu07v+r9YBOeKAUKCYC2rRiPgC45txiziz2/bsWtI7rxFcFUzN3jrvO
mNCohdTOvxnuOTbyNJkzDP86BLVcFcz7VqUM0HbVG4ACKJZGvrQXyC8JXo2GGO3r
ywk6O2rQot59uOJmxGp/ywAqZaBX7UWaANw4vCHHK5lrC0r8gQ/kGfjOv/UMa/vV
r/8u7Kw0Wb1D+aP+vsYz2CKFnOPUzWM9LGFYNnlTogtrsXLxA3S4hwEyo+CVGrJ/
BM2c/EUU3x/XiDXTXkwRttXLp4wLLGi6mD4yK/o7+BEzCZahBVIUlEjJuyONQCyU
Q9YEPgNzFC5fJtOxy8i+Hfadcfi1dFA60gj+lnkt2pNeL2Mux06e9f3LKeMZKJrD
EH88UPZJ/nhj897pRiNxee2jlUKRBtgfAHBO1NtCHZMVbTCbJpqzU8+DCp1UDK2t
GFTHPL+Co7S3tkBoA34ua7x9taqigoi1sefpocFUqh3FFbr2WzogyKgnkBUPRhpJ
gVcHiVp+vT4yTn49Om/6i5HiFCU54hxDJauwewfCYIgyM5gnWweMNxeQpsgUC2cD
1wP5C1dM/lwbRAvn221JuUarDJj6usDYjsqX8P89JMIhBow6mrgeMG9p6ydeBNiv
0GRmiabyjlbZbwTQK1BfyqaG3ZtxlgwGvFl8lRGX7pkChIOeiO/E+86XludLb7bA
qv3MP9ESWjppkpdkVc0XJfY89nFL5QbRjQGDtParIu6TE+xf69FVLVEw71Yvb9UK
NFldaXhn9TE02snyFAgK6EkUaWMP7Xap9mg+w4GPVyqSHMkL+8MfXCUXb65JUqP6
NUra5g1PYmicA8vWOA2RoAdEqyVj1aASMqTmp1zJ8Zi35J9bY7iPsWqem6x1M929
/4iDpv71vQPTYOvTn9RoIfqqiLG295D/ZQZ26S+uGTz651JtpNSoswuOK6Q5vDVZ
7uL6uXplq10JJsCQHe5vlUI8XZCyfHt0XK4Y16iKm3UmvBuJ7Z5ivRyg8owwcLtK
wK49uwxot9J2xigxHmV67qiGhy8c4EjV/3Lt67NysoIjfJ/MuHVcs9iNSQ7W7LPK
kJgQ50LxfBLh6U1TgEzn05OqMAkN98BVlf0tui3LjpF4v9FusgHM7duvrtuIBfzW
vO7V/q6NfNxEzbNzMwPRgaCgpDR/xDyMF+fi4MgG5lW16LeAWGZteDqbxchdlQKt
Iu2hyv5yUUbhbDfaL9scyE3ftpx2AL6dBYWc/MBkf9CRD5r9Oz230u9qJEMkrxff
W/sQ/PPskeCaNzaW8fhInGgj5i2hRBR63r2AIXrTosq17lSBZ9YVadQJ89Rgbxse
qWaHrZcpaLkium0KRuCPhxaghwYixkoXPuIQtCF9rxTgVzoGDGyCqZfXLwqZF6SZ
LHnZmnTsRS6tndEBXWeQEWZSC6Io9tpqBZEuS7q4U2SLyRDqkjX7wuZh3B9CVPld
yHcLrcsnOo+FneWMIJsUA6niZ3YfN+nRhRmsVolYXDM2++aQu24fd1mVAisgjTnr
Fp0c09R6MIgTz3h0liqxgP3wWIZX4oSa8MYG64yzwo/bOxpXvMbEDMNJWF3F7Vah
4Xlms3QOaBzfdZBS3wvzkTe0alpfWLn7o57SYWHRW9RLNjjDeHyMOpKDWIT9DRzU
AsimO4b3rZZQmRaw+9equSGCCIbeIZDWJo0sfYxmw98FzknbiGL4DWlBVTCo5kA+
qp+BNkAto4DabY5Nmulmn941dQwREvzF/gRn0WZcRNUNNn7B0RnGkltsqSTOe1Yx
WEAAc/V/jRaenH+A43VMnTFtAyLt0CzbUzryUHYPhKsSm7N27VvaR3K3pEbcLfc4
xuaYOILIsFr8oWaoyZsDtZLhMNL9yICIK6fSxv4EgGb38C2IEMshdZ8ls5VgXvsw
PV7mxt3jEcGBv7oHDfANCtr8RpcNbF2eR2d2x9XHyQFgzy19aBmhCtqa0Gu2ba8h
F/ofmPJug/DAj7I5ebllG4eHhF9yssX2Sdsmkae7YuNwWDNpDro1eM630XI+GSru
CBWmPhmJXOhiLBW178/06on7/3hDmeyTYIBI3Rzi9SgFjRjAQEFOqV3HaW0w3HcW
ZOTkL9hYZayKlkEyb5ITXJQIJErVJC6qjtC+WLibr4R46mRKQqJ/viZJC6OrmSjx
b8148UwFwaI6qukNbFO/YxL6LXF8BWiOVdUP5Yxu25g5ifE6sEOprn2kkBxflyV0
w29RlmOFtybO9hgh+wjRHZI9k4jqEhnvbcm7CuDfXEOpnqmBUfqxdEz5EP6g2n7G
jWqVsxlyTU9VXar8qALBrnA+RxC2LyJH+jjFF5lq9aN96OOT5rF439SvqiTBye8Y
p7appMTL3v4QDbBT2XFMEZAQqmEkyKsRt+IrMUz6Qs1qdGo38F3nJR41DSnLBpmV
ZxGIPsntYJl0RIdgZAIybmXHaiJweNYl0WRXauNG54XOTOqPuzFGWIp22sOr1AV/
0eYJTZWoDL6ifGHF5cllh0i/8rKj0m09M1wK3Pwgv/6WwEvmOaeW/bvSps/RPSHZ
WgNHlzVorYzsc2QbbVjMjNhLDM9B7yadY03RPKI3jWDN8VKYRYMH7ohSB1ubNoL2
Ujs+IvbCI38c/8ml9rp29ZZhYnvxAJbYdeR6gG+Z8FAv7+u05uFO36Nw23rWw1XS
p+BWJSOjwGcamKFAv0R8igZO3Kbf4r563/s67tTgXlnrGDTIWmQj2l/3QrZpfVA2
6hllcpecGzzu1CMgyeeVF9xuuSiBudTe+CE1/Ciwpc/aTH9ieNtEl4fzikgQxcVk
fj8veQe8D6EEU3zC+rPxDzSCwa5kO4sGAiC1Q+HNHUgiso1k3lccvF+thjX73lms
IT/NMaDNxtog8jpgKzIF1qnbDFysQ2AeXTmhqjxl1Shi9j2+yHSocj811MmElQuW
Cx9dAw/BqwfPB7DGqgB94H8IFe6W+Sv6uYDWjKoVCYzQ6B2+DRKFimcUGMI4Yhdl
qi9M9BLvGnVKA+bax3OMlPy9dmdWF8Q5fuC0usgL4k3Ilkv2XbI6xGhHb2fHy7vU
BwbjMu5rTE3YBJlHwAGFDZRln2f9JdDmuKBO5o/SmqTHj0iFq/qbNCzvSS9K+Trd
fFK9EmmL700tugBQfCV41ElcB6VxJGtHzT2lPJ+VNkHM+XryyB1Y3KaZXw+Bs5Yw
RIeRmh+AuXHsnbYHx9n8DdPoT9ihdYS9F9aCvvTXQAKcLZb7n7wv4j9lifvfPXQu
hlaw927snvSeJ5sicTg0cJDQL5tDiBOt/jlTbv1JJAuBQ2+M+Lwc4BmVvyx5a2Ox
Sqbt+yNXFkn3KI+YnpmcEFTTk90o+4VgUBuFkAZsfNP8i+8rXxm3ySLWTZp3mVhm
UsixjLnBclc0CO42/DOZ8NqYePXip68D8ux5lzLEUXAvmxHK+RZ+fNv4f1E2SXQS
XMfsvHFvbPMJIQJsJS4rRZPKDqUru4mSZ8ZZbBeZs7MexZ6eU0ti1XhhTsd0KuRn
iKGj0erGLOxm+NVA7eUeYFj98fZ6mde+ReS+FJRm4eJf5s8vMJjUa8KlkYqfFZqz
yOc1CWmWwWilZP7VPhdR305aIyiPnyVFLHZwj45Pc17fbKfw6hBZ+aFGHKIu8lpj
qgn2YGADW8BX4RGmXPeAyMS4TUcUHyPryiqPkjefUaaJ25z4l8Wi9oC8a+UlXXra
LF3dqe4jjyjwjrlh96QBvuM3QrZy7iDQhgSAvZi3OQ3GtXyS4yxW3st/WmwttYle
sOOf1Yd92mLgXayRZLvcsS4jeyIqlQCl6CRzA0fUTffpCAW0VL3SnvD47aJs0ZAu
+kVxv7CjaNIt1VUURvaV/QFjenClafNQSv5IoTac4AzkjP9DCoCkYWLZKFmHqbEj
B+5ylI7FONYuPFuHTDJtVwd7WsXIx5q3MWWWTueo+EjLX01wUIUTSbwWpPAt5/xa
yPzAhTKTuqXbDb34e6YlS6GSbWlbhhJrXiZebo0mrQEejOItM9hLQ1QcE81RQFN1
nCXmNUszwC9HEiFuYIiNJTjrbtfZAtr7aZUxdf3KgGzn2nUx6tz3TN3heDJu18US
jJwdsKvwo8WkYNFrT6DMzNnt/65RRTmDWztsKchlk4eDmzrk523VxaJCETmndsvB
iFfzj0brATDZwL6ip48dWHHs2oTQ2U1H2JHKTpgNjrZ0pVYg+zp0NDlZQfJ+ayVa
sL7fQbvKJfMCheJ0BxiSG67OQP1wyGo5q6K38Y+fbGsvi6KkvCwQpA4Ts7zOH0XD
55x7BMRuLKuqsLYeijqsVnkUPNJfmou4fikfAQGMubJN1lK8CpYt/RMSM01Aj5d8
Th37oA2pBHNvv4kT5A2fQ7D7oNo1ZldZFym2eyegRtu2lFm63P3vr/pqikKgqleD
k7DicWKFPHlsT5ZCiK43LpSFYMh9CUV8xagnc1mnIDAedg6t8crScOK1Bd8Z7Nsd
OXp20OWt1W0KI91SdIY8LzZQ+ixLsg//SB3mz+1uIvs4MqmaQhFSgMeVVL0dlzEf
Oal5MnAFg9TOC5n5ggwfLsBCxZulYSaZJ+YA6J0rIIxd7/LLB02kNwidVPPd7R9w
u923/gVWmMnclDTzTxCTwdTc0/yHHUzlBI5Z8uh+FKFh429Lj5haLoOtPIJ//KA4
DEigbWUCL4AAg6OYij9GJlpCAu30uADrC4iQDL1hFqv9fpgCFmHRrL8HdMkuBnqJ
VT2gU6MmheW7m5wA1Ux7hPr4LNE/YjCSh0L+5KugMGuhebitpR2PW0yofq4PA6Hu
z/obPEfMHougxFivEuykY19Pgtcn4gbwQO8rrU+Xr/kyl8ps6JgzknTFYwHAgKhS
aL5AYlSiHNoXZkY8+cps5CKRKgtD9Ej0qA+I7x9NxGJo2OIO8OueUrwg2zq1u9YL
WJKE7+SHblc3B6InO0YzFEs5RdKSYTL38QlO/ugXpK+RJhdOj6VNrSnkxvCzEwPf
atlJA5E3Q9YbsnY0ATrz9HNk2/RI7gaklrKFbqSlvzjugjO2I1L09vrLpX7cB9vU
JOmuoVPWP8ZrTJDsDFN6r+zQqFtiCDjVAO5ykzqx9zFua2fX/iKzrIquMk+R0G4t
hAtX75mM5scHURe34aLV6MctMWfF5XFjq60zVGiCCNjAeyZk11ua6/uQUpiffbp5
EH6bOnL5gi6fLZpb92O/A2DnSGrNz0dOQMAd4oPK9hWjwxArm8Iyo5j9wiQcQsL6
pK8eB5NQgWBwPkj8JpVXGjfC1yLtRCWP5At5ltuoFAuQ2x4rjQv9aFXtivflnajL
khbEudCqPameZtL/l6xqan0mG0Zw5ZDyXcRP74QSxOiwPnykBjQShX3JFCtgPuda
oesOuY5OdyIhdZVLeoZ7Szdr28h2URJwTg3ztFawT23qo2KMHYRIZFmAICtkjUt2
VYBtiVtQ/EP97O05bs/JkZeBrxQERE7PuFbUkI6iwUg8alNs5se1FU2uobxAwz/+
q2NAjMWOu8T0zqErLFjTwr1Cvq81FxqsJ30Cfnaw//gyWV34eKCLSb/V32Fo+Ulk
Q99zifex+oSlig9C6f2b2LBlyfJExcZorDvNZpIIwkRNq8OkKKo9VIsQahaNV+yz
Owf8Vz5dxQ6sswB4YyRXWLexWpArf2DwTB3xjynR+AElusMH8n1RHMwTE27UAKjF
ZqLw77BFG1enCAAs3MuKOd97436do43BuMwq/vrYFSt9eOgUK6MxZzr3zHNSVV3Y
WJKuVYrXF16lodDL5jg7rOlULsbKk6hpkin5It306e22afHX3vbBeMjXA0CFSSv7
OSNYXaWqfElQdwL0zL5a2uSMI0uQCK6ls67hr0LoGDo+WmgXw+9tvDohaICIPdg5
OaVNA/nXYdp9CXBs7NMQcEUXd3x+guX/bJm0QM+/ZkZspDJRMtP0Uwo60M4iqkqp
88InBbv0IRLw3vrRRgvw4Jz90eW0SnWqK/VLmzpaoI5khZrTFnmyK2I5UUUi1q+I
jgWzJXtM0y0OVhEsg0uSjysd1TGH4EJmvvn7r46kOX7QWOsw2G1KRhVC+mfUF9Jb
hB/jjqZBOiM7TiFjMFVZO82WwPZk0NGNNZfTlVfsoiwlO9GHVBGcIlM7zhtNqyLb
M9vCzrmqiGjtVSCsfaTNy+R0SwilBNsgF76wprlQrRtA9ZbFc1EkoyZ51mf3iSEO
kz1Fk9vhcCFWRRoPjGMyIw05ntlX4w9jhYq809P9zJHso1eelfzAB+pQUTmndWBB
LSFpM5q6/1y6TQCwafHJeZVTqWsfTUecRKqSTlZdO+AfltG4Y5pim9XJWVTvdYap
Mh4ybiwPekhAaXeVFTOXRH+ZazvJniUZ2VXCaKLQ8xsR4zHV6QNZzK1aKjuUAYJU
kgCNyq7GYnavN2Vgco8K8EA/6T0mE3o6TlNJfxDDlW/6AKaGMshy5RjRl/J6a7ba
/01hIGFV+cN7OwYZKCUw0tIcOPQfcAhgYHzCGCIODwGTydsHXVncP7ta94yBSWn5
Xv6+1G2qDOShs8aeFdmcLfF31jOeDEUAhxiOiLWAtUAuBC58sx1rma9jxMSVR4l0
/FFAoAvcsoqFH8RVyeuWdUMh289K7S9FQcqvNzlN3VsYWhDcOBLlgopgOCqBANei
fPek867873WMXgrDzztLdMZiehZ2tbAZ8Uu+rh7EMT5KeHGSTQkJzxnGNcrQQYro
wAV88jIX3JauS1+Vy7fZqIY4sfGhUQ/OBnD5VCNF22BF5ykM82iG5S1F9oJ9N9AB
GGIIFRFGA6Ex2Fr2h33gjfnrpDcKPcTEkYrAsx07jl0UD8Em4WAOg2/M3GrqMepS
5l/loU0RT465fFtXD9qMHB2jXXQKTuVp1YUW2jXN+qKp9ZIq9CAz4SfXKizUbDJi
c64XsiWDxcFy0ywdGoZQOqGgDPaWfXv1ASF7OiED5Wsot/r7tQoDQiGMSY35k4Pm
4is141169Lm2X3OiycqYkRGDpdbaepT7sABmupmg2DpFxVwgBmAAmapnZHYz/pBn
pndFPFY5KLE1TqPnnWr0BhcIvtECBkpI9PzhpO4ZWiA3XjuClQApCbM6sfT4/7s9
EP0F3yXfeweWcQw++VYqlwtJpzXfgUGhtNj6GMRV/Am9kHpMuqiKJL5edVAHxmp/
4aC6y6mpLXKCBXp3JNg/+1dIg/mbzYQ9pGnzPx6JewTcLVpKWN45nusvlbfl0etI
+QHBW3AFvHUmILBE1rSOaXdNnS6U54YbU7pYcBSvOhuiR3/73HJJxb/PxZtOExyo
+TREpN7uocZ9666QMWfjYNtv6TvAnJWRTF39nI4qCfVtrV3OvXqo4G2KtE2YT52w
47Rp4ygAc/1/dwyZ4I2Mcrf9z/Wd2yjEbepLp+demi2FgAyEXg6VEyMrczQp7WY1
vI0jRxZfh4PKxJqgj1q9i7Pvp7NNW2IbDzim6U8B+XgCCU8AcgWJ02CXSBIl65Ab
ToiaMsZSx7HdU7Lv/PtKiLi9M88a6Dzd4JYKTN85BB1dAp6g6Ap70yh9HkwRANq5
Pr2ZYhQJUnbGJAMgHpD0D1xr2jO0zu6W9xm5600MbrA3meTm1GnlpcIR5B4JHZ58
4+FCvM5c/GDoLC39efIRTYqfsVNsc2FrUQ8JezIUrXAxklK/h2cE7PsDQS1fdN77
Fp/QfB5V/qPg+wIWgX1TzHg3YxvU9LTyPoHHk27AmujCurCiFcQ0AEkFWbmtau/k
DObOLA9fRjy26xKUks1FFlKOoI5+jUv58op/t9zkkyNrkD95+eXmzh/OXyD8mYYj
ZXt4TyFaOhqvdt0sZSwuwpKfE0Pry6sg2YIJ67rpGwvOzkc5cRPf/a//EfkpCuZ9
s94Apbqx6v0edMgbhugTSkbxhoABkAvdm6Gb1ait45L6dRR04NSDdmcvP8bqLAYz
N7HfREq7Rxp3bse5wMCpybu8K93ceMpyWLC1BICMfnVhLPxyA1N5lG6OlXS6fJYW
rdFkYIbyvG9oyI++CYa/R1ZmOclxiuQEMWjDFx2QZ/n7VK91VaSCI5dsbze/FSjs
8Ca52BC6u4IUxCeIsNiIdEB0x6n35rZWV38P+Py/1dvuTk+esxTvMDWF2i7HZxjF
4i3diEE0wKcd5O5m9ST+f2Bpt39GaY5EVQIQBjVC0KcY2POPQPOyYbfBUlX2T4vm
1Fjbu4tOyQxQ8+aYwUs/CzDsCe279wEm/q8GClEim2eQQ2FlPDWWgd3P6iCLnbve
OZU+cIs4ijGtvScRjVtxkcVFbeX1MmN3r4dvVH93FUvQGf1Ceh4q2k5p1bXFj6St
l2EPZXZfDT2voJ9Drq8RTaqaDqf9f/x1SdJHyzDuu1BjTKu4yku2Grk2W4g/MSfK
bRquKwwbv+4IO1MRvGAkeIXvU4MntWeoexsh5IRPgHAEWxYhrrQtNiGoE1vNyLyh
X5IefjlHt7VS2xoNzD97AL1XF4hDYRpr8bC08rxXKaeTwBFOcl+49CS6OdBfNOCW
7imtojH/+4vKKeY7CUO+B0K32MqGZi754lLAJJCRapirlaSYI0iXkWXqOVlYnO51
IDP51fSQzv83G7eZV8ieQ2o6fSlFp+poVmbSZRsf/k+1W2Nf7xukjwhFlPe5390O
Syvsbm4UjtG1G4lyFG/5Lmb0LWD6fnjgr7YCtooQKIe4num5BqDuB8Eg8ZB8dggt
+1DKRNtuYBKN6CgpzbIzd4KuDQabdWdAZsFdgJGDhG+SWVRF9eeDzS5GAWGK6ySj
g8hwvsBI+8gMgD2KtvZUG0YC0JH1OeG7u0boIE78ZnhV4TWfsOCD7hoMDvCInzms
TFSqr2qbI1XH7LxlHb6B3wqWLxznzHulS3uXIyPgy/zdOQl2Wwq/X/fg+OtbE7WR
gott9Q9+2/Y3Avn4qqp+Z7U021jvG/9LBPYyU1hpqb7API/8i2HGclD+ePFXDeY6
FPpwwHPzLrTuhxYTV36h2qG6NZf/DQuBIovggWzdi4CFWutb+acKh35n+Gf1AGQc
tB1VJiw8truUHE/pSpITrjEZnZiH7TC44ZLCCH8yktBjMAD9m7ty4sJvd42HVD13
dJOGjjuHd2VOF/5pXdOotwkoS0Ye9/OkU20g2WXgxRA28/XLQlivWwS/HC8Ak9Dv
y3nXgSoXacyKm5dXnOPOQwf2FjwVLF2aOZpq/hTXjqym9GRQEqH/+aen3/qnBHWE
3aaNQCHl5cLzxZgSQBa3VPGwbd/twCp37w/RM+DQNAuPtzGibz3l7trhrXCp11n4
deOrxrJ/slp6EISO7pv2zVg6upwwmtlaBZZqrj/efA6O9exQkYhEvf6YaSYoPSOa
RaNTUNSlg0wq+8ZsBJ2lclAu3RFXvt49f0rI3s2EzHVNWwNTxlKdG1NFPqY7XYZu
DNE1sqWputh+ZSsAyeyV5CNM6O7MTcrMzgw0qAgJ2rk7I8uD5fj2oZ4BKH5Ki/dw
7IYp8n3G3lws/CD99CUSodmClZhxuo0BR0XZBniEkNt+EUSgRCZpS7GpHDNGjLkL
hgEQETFqnI7KDerAzEWUzX4gQUlTcfc+EAp287HcmYGsJyiffQ3qy6DieiHaBmzM
NNvUrwvTaS3U10R7Lq+GdIzpq47Z1spTi4ZQBpBs0aCCOfhwQisApGTazq/ZSA7D
w+XNgzUDz6KA6ae0KJJDnp8wdkp3/VoH8/eZ36in+EC8heLwIrQeeNFNWPFcMxjB
zNwV4bNUNIYf9OnivJ0Xqrtn6jVH+D8Y/zpExxfSG2uktAN4FfMMWMz3OYBC1/Mo
8b3ReF+BEI+NOiKnShb6m16FoIBf5dqXqx8YsdDXlzg7uixsHOozxH8cuwUAdMmz
C+4Q6YxVphFoivoERZk1W74km/VzD8rSTBjhAJikzVCfLVtbVqUz+K46srHdnTkS
rhhGWOxDFnqdvrhnkE/mzHV5ozRSzUA16CDQDTHxA92Cg4GEUGBNsmDajp0YB6qW
+h2sDtc3ekAYcI24r3MC4CC5fIGZ38OYatx9eF9LzqXTbRjSGvzmNz+lndkwPnlz
sO5KC7zMHVrMSRjD37LNpJr7zpkcRw2zfatG2t68SWw5oa06jndaCCeAgnlejlKV
wirjIIXJ7iYjSe9cfvO1nGd8bQvRH1wqsaUHdsHLyGZlbRwACVgWQur/9BbU7JQJ
2QfPe0Zx08OyTKYCkJWA6hWU54u57lf2fWYc+wSAJMDq8cQmnwAxvJIAb5ouYSzf
ViBpXrbWgS1GEWcpXcb+OvTIgPEV4Y+qXWEuJRAq9Re23OiQehs5S7ale/oex2+u
XKNPNiWhvf7GjX8bBVZwXLCF75CdD+h0CT8VFJK7qTN4PYDNZDG7nju+VVGRHz6Q
b+xIJcsageAlIxv0xuJ/1GE7an3jrmmIb5Stt6C7dQGDTo5z7QfYdBfnvTDsvx06
/k4kBrhZ02RQLj1MsJwtbX6BcZl+U2uGQ7w4KMfE9AqUoog/YPVDFh0BbCIwhBA1
+S+6ax+dKEVtOGZpl2octB6d9H676KbMmU6qyC3p8ot2j+UkcMr3cueDFZQSf9I5
mjqgAH2zKAkdUXZdiL7jhQocjVX5FyesYcq/3obCqn5BniCB8RKQI6w1pOWxH7H0
KtMIviFQt1GQbck7jsRGuRfAzPsQsFsIyZuHqrU8Y748OgEd/5EIadlqkcmxn8Su
7qvSfqxLCLRVtBUfgB0Vr9Q76oWHjkshQrEs/zAgmgScj300DfmgxVF4PBLwwzXU
mnJbBaej93yRzBQJdj+BUj9pGnL+gGsxD5D/35Dkntf7OEQxre/qG3ZEqttL+MPS
Fwpqe30OYFmKAYe4VvbH0Z9/wqKInJG7R/U8Gc4bZeL+Nslic5LwDs+X2K/LHEP2
Plx1c8DhAw+qrDE4oZbKCqPjbJlhHwtB2CJtqGuTKc2wteoJgnugsRsNIutoXJ13
wG/B5gCoCdNxLlEIbbbP9/D7Kfo6t9SF4a3eH19NYEiEYHyPxqEBjww3B/tKYWTb
LvCyfdnNnNt20GR2QgzvLHHqzatawQ0nCTGuQPNsLYRU8eMAdfLABLByxrmV82ia
F4E7fKfqKLuhF2H9B7wd3vcCGE+jjmkfRtfYcB+bAq88tt1LLI9GluJksB3fUDgB
nXKfGlLYd0VnNK0GbnNPrWweRkJLKyYpNlzfyuNg9HmZAkDJ+Bg5tDxWpcJxL7LK
r23dZ/OlBVU4b873zEr8UaQe3k1gususny4kh9YFANWJjs7K9SNAp5zrQbL//Ej7
vCdC40YktdvTbVEBUfyIcRHfBf5UY0JPvAHEeGYmzfV4p0G+Y+pgpSmZNC3QyTGt
1DYT+yZ3hPlleejzgNDA4Xa2+W+9VOLcvt5Q7jyJsjVsby875MYCa1YTrYI/MnuA
C7sbNHw7EAimL0/C7E/53st3zvuXyFlXqs4Tv1Sker3jgdULBM2hVBitpamiLLgH
dclpvkMnbwqeSCyVep/vJ/jrjN0zfqKokZxJwXk66jtwk+gMkEa9vZEAoh/8C9lr
CdFQondFdco2AOaPwYCajhFxoeLJgEdrkIGL2W242sNrSJqUvewADd0JaSq7/0Ca
jn/ciDdAnFPfagaoTZKPJBuBYPJaHGybznlhXQ5VWZZPXNrkZkOoSlAGj/EX56qQ
+O2jWfG8+ywjMds6mnyNmabui36k3njr0oLsC+7ZWCe32qEkI8//43k7e4PYkKSv
0JO2zur8x1Y9CS8ATUDAtV+2A1a98dhKxEYpx8YAGPSPGGmKUW+CQMmwihpSwPIN
LdMJhS+lqTPB57q8dv0P4xz3nB4sjdvIYyojComFFJDwx2wCV2S+wgmwttIBPATd
zTtZOBBbmgbViiQeqitZCcsyQxzfY8j87xdE3utLuAmNvxCULGAG0KxwigNC1ocY
1Y/PzI9HSiB+60aWrV1eMrybXSTwds96SHTbX9sxMHnRh5vNlCL5Io5BfFZ0s47S
6TdGhliU0yY0AxHpX+BHQiKJ4bGgbZAkGYKyHsNr4yymVCzS/BaKCqfnd+PX88mZ
K2LHM5SoNs5aHfuFE64OO7YUxsX+u3MbIl7CcXgFk4p3i6kES76NKQ2zW0gDLTKo
VkOnxeUfe7uZE784kBQW6BIICM2row/KqorkW8y1E/86She1u8GafHpqyYt3yrXp
qXukIxU9KUkGyrilsHzQW3n4H6kJXfCLxfX3ZA6e2/SXPHB4CZO+zORgAdnwKtKb
oN1A/WpAFWGmMbhg0cAhmKXRvsXgmcJlVzloDnzG8MS/9jXG+n6R9AIUXkCa/wrP
iZi6aLDpSr1DImdagujOxnqgBhXLUmT5taEJZRXx0ddSNIdkDgHdQB6/M+xy02J5
vMqi/U6vUGazBOfXuS7SKsaO6j06hjPuOqgu56MikurLJT4OaJ9xmQL8YTg+hC1a
bSXawNiNxVRVHfBec30XNRNSdieBTT2TRDq49cIISDCWi3mTVTMkoG2dFdZ5jJsz
vmcczCKoEv4IUoMm4GTYUvOCv4YjmbHGz3hIXeJdn6gB/kghkUudjAttNRRv0Xkz
vUU7e171hjGPmuAvc/UwQMLPI94DemnoREtBCwq99zjrPzrz9nMEaUqGFsnYFkbS
8x/GXCKhYQ5AbZY3n6wfRQcOydKQxk2A0oy1lkCXbcB48+jf0nqbkJbyCY5UiBNc
8pe/47sLcTYI69BOkD06b8sTWNRrgUkfaU1RnaPCjRHMRCXm7qSOUDuDbvDrBR3v
WIuVjf3pWN2NrQWuFt8rrRRN8xtPIlnszNqIiiBnf44p8bdvhZY+QAdCRblKNdZg
VrQmn4CZxAdkL4Cb2CPYhW/X4my4zm0dAn/gdk+jUcZmDt/U3lxrBOdtG2Nw6iac
DKiztvelverHOrrcARbGqzupzlPqIKraeGpLKoZaBGs2acxB3FMvVX8YwO4LLi1D
sID0dzix7R289sucGty0bNNnzypmL19BDr2E4yEr5Djn6eYz9zR4gyPh4oBVCi31
5l3tsVkynXgnky2mUVzO5O1wZpp1cPk1qFgfi/THqy89aej2sO4yEXsZ2mLUBJa1
aOTP96v5V3YIliMNCn4KCl1k+qWXPJ5B9XcJ+1F/cWTe1BzSbtW4dUrknK3nQs1k
HZ2rJJyT6ks/IA/N8NxeMR/kR4ybJR3/4BegGDwAGbMmGNfeRJszrl7CXxeHL1+h
6dg4E87EroYsevnAUM5AESL8dUNYvg447QFWA34pT7YRXtPfxwcdLVbuszI46Xlv
Kyi9GNjLsuQMKqfrUeSnoyH9fOmu39CoDAup4bv2wipWGreYliDf5uQI6WSXz6KI
k95EIrFmXn8lkN2SZoEVMb8Cv6PupVFYWk8i/c33edAnSLdYkrtDcbFP/yWx+cBs
p9LLO3iIsU9V8Y32Kq6tqQxHhk2ZYu65/s8O66Uqgrvw/HpTIRO59WZ8k6bTZKdc
1GnkPVQsIt5S+XRIiFSbm4AyA0TnE0cgR0+J8Ma57mHt5I2odRujfbSftSbuNSKa
cXSkvhydaDDoMF4x6TkaKIJBosTO/MFFg10QyXzgl2B4FS4M7tImmT2DnMEbT80U
e8nNFI/PXu+Ywvtqccm5Y+adTdifIeceirY+hvKAgt4NZVt053NNty95wxxUa9Fc
Z5YNJkkePrh1ljP1+0tuAS9oJ2rZ//9j/NgzK2n9ff5T7hfc6shQFH5+ob/CwnOq
BPMSf4w2GGZpQDBPVnWpJuiq63byxmf0nrb0KTA8ri2a5TigbWvv7yQBbzIWcXbj
RFhmoz/yWmrXJhxzZFpKNOJ6Ns9G/2J0YBSlvjz1EQg5iXdbyaOfJcbodg6ITbdc
xtT5tBv1zXk9RvBn32Y4scpU8jtv4hfD6BZDrLKcJhh8Z94kKsEgw73awV/AI/Lj
9yHkVPLY3OX+3+QA5tTsqUph+YDmxPPajSiJ3fqHgPITdVcOinZihzNIkE1d+IJ0
9mSwvf0jLNTLhnATbNNXRoFisw1ry7burlnLijeiE5Pzy2GTZCBieMgdGA2o6I6s
irwsEyw1boDOLt7/F8B/IYb54ul34hmgRTETSCMbqeRl3+dynYt5CnLpv4oWPjh7
reXNYgPtfYkrGBE2barHLcLnwYEP6S21OKIazyMqlvXsbYsVwJf6KKTC/UOopu7/
H3uRX1F8Sy2rGjnoRFC1wrW+G/TliUFVHFTni392jvcRHm21i0xZ/5pVxQDAUyUm
q70JN6BAKuBnlSYDRfwnncEuuiGUG0dAdenSL7ZKngjV1nhb+LEcdFV1jMIi0rFm
VCDwNakMAipfa4GeMwKloQTdWzbWhH5L8aPOU8nrL3S6WOALTTiRVxMkO35l4gwD
DEu4KqUUbAvnSeOUdwjccYAGPcNYabwOamRPol5RN5qJrWF8n0bnJO8Q4xpYH428
Z2MlG6WdUqlfm6OI3jLnzT8O5BPAYuVrU1zbNp7pMlLis8b0AKLBIJKhsbEc+rI0
3Rge5yFFXZL5cqVThNOuYxnYz2t102Rp2O/8VgjaX2d9935FPi/ObpON/btk1O7w
0txAVcWB1DjobuLZm0c+eYKoHdGVpBR5TXFWw6foRQq2+2tjiu3vapCF7NQLm4rL
qLAXx0ADVZp9P4R2j9QO1RjcOV8ytvrW+Zl29EChCU17ZxwHwpjo5p+YVCDH9PKS
eeOX0uYGuNlnW0pA3gzqhZI53AfDVC7ubWdR3Wh79jz5tVYRGItOv+YL9oR43tnl
xwBN9+SK0UsKb8nARX7FIfbg7sTxqUudQLTiRs6FcrPaOYtuxxkPymUJO/+SB2sj
zznG4CRJgOxn3/dUksiTwUWqj/pmj7li4hdC1z1mR/WG0KsGWSIgBFkAy+ZHaoU+
UWHSCYpRJh83V7dQIU6uDkl85VNgtPQAKIN6l6i3Xttno9x9wAP6Wf8WLBHeYy0k
7EJakkjxEwZDB7oogFzD5LGscMcDRsXisPEUgmqYkWHF2tiHU4kJiIEKQJd+onY8
fq6/2kCNHsW0J7uNDOo08wMjneLkRsh7qmxxuo6IgoteQS4upotf2oZxzDgvE53V
3w5iSg5oiOROfbJcVrbp8rw381F37l3Kqx3Z658r4iY9j0/a267ORSP7z08ZFnnl
zT6WjBE3qVL5OxGNp2NwX94jmQmDZCeu7c3atMHn7CGi4oP1kuo8z/pzpm933nT5
sIBkDBKfhqX/q1sU1V8qpmEYku3YQENgVMWNLFDH4QXEbLLXMD4V1I5s5h6PTVaQ
aPtnmiqlwM/6gt8f5fXNA/BWyK7dHJPBzzzowMHUMMB4vJSs3F2hcQutUrpnMuY9
oDEezdktvWVW1tUSfFrwvqYvPBooNZry+HjIAVFsl44/sL5boitiS9RU7bX7SI6L
wpnW0lq7rp4I25hBznF81x0PtPKjJqzUgW+lHxW7aJv5yAuNt+6IO+qqxMD9tX5P
lfRMpDB9kTw74Kx/dEBY36UkP5AzDyITxF7zuwOuLa261EHSyzr9O2FXXhsR/+Uz
Ne6gm39dcMQejAO62GO7dubVFbHvZqjaysiheIC0c7fXQggLLi1I8DtDLTvcJ9sc
zKc10RYR4HhegbvfZ9Fpdtanx/uxjHwoCRQ0EnWul5pHVYu1RbqieeWuSu0ux/Gg
hFBxDdAvOtj4kfR/hAcA0plogBdyO/JwhV2JYRgaCBFiLyVf8EWtI1zaO/yeAtp1
T3GfWk1e6iy+lXcI7LvFtc7QHhc0+xfwUl+IXKbeVHFIbV1+dxmi66HaFtFhdF9s
dGfDfcoZHkn6psYSRbuJGbsZVkH2ALBRBXsnZ2R8EWxXyKLFoYkYZe3a62SF6CVX
3zj02uBeg9v6BG2/jeC9pnPykBKN+Wi5xPaX7LZguobADMY+wDQDAvi0fVVoQgFc
YAjQFh6230R2m09/ODJtYdSj/1pInS1F1R1O1MSNblMWpfC5xRa2mftZOx1+5Tzv
ZLzAbKHLOLwU/iqzK6CWsQPUJ5SEpE7iGVebLlx+coCltoKlALurd2y8/EgKjM+8
8/nXeaFc6t5sPQJqtB+t8aJSTDq+2bshOrce9CqFT7gSFt/IC3/3HxlAazMGviQx
D5vjPLn/ikvHdlkj8S7mocUPYif//d76x5UP2Fk6s/8kBg4X9KfrsxjMvCe4dsrt
cWQpcK8vOorOKS6/pSmBVndJ2p433Rc8b8gw9HsAafoYzKo87CKldOYkYofaqNVg
WBgQILVSstaExAZ93aF6rSENxb1IKaUIRl4YIC5f0XQawF7EJBJ5zG+RxYYv4qiD
nvhOwsWnBmIQMRRhxgl+ZoAxu4TjnGKFiTi6rPrp3PruCEmYBPS7rXS2pBRbcX5w
ZJ1X1Ga37QHAbyJ0G3sTNu9N9x70lN3rSqqNL/h4hwj8U9JvPRyPxVN+/MlH7MAl
kWobhL4wd3zLifZyhMifBVCyK1BthDhFW42rC3P58YfyhDNozzEhTnp3xDrFxyxt
axBDo8DljIV6S2nElYXNcs8ktrgAjrc2FcaJdF+9Is/KowFlq/u982f9cFQVw54U
ctLRboa3L2ywjv7PkDS3KCPFxxT2XE7EWKtu1+HK0ACWgyKISW9qgaeEEWX00KKH
qOuvVSlPFjiR70EJtNxm54c+FlD7itM9C1uR1FHBh1BcwCZZ37cPkCPCPB4cyOpM
sLLTybR3VR5105cmgXEm5cFHihtdtxq5s2nprXZ/RlGdkdOstGJlXIphSrM68meM
ymE4bgH0tD6XLKDSM6eIx68nRsl8fMIgLhDIkxeki295GAmE8G9iaflj7mDxPxsJ
eIAOxKim9PZ9MfNkqHgNquvXlWrLibPYsijNNLq99LiWxRIzd7uXHO5kfaBG1CQH
1es1cxiaDKei9HeFrApmA6rMhoX+P8VgdlA8JLlms3T3L6HoWR7MtVK771q8qRRb
a36muzAlkrfIoSZZkZtC6BrfY3h3JR6IGIYsI7/xPO/RLSH4UEV9FMIrRD4JJ+fM
l/r/9Z6ACssBYjLAjK1aw8gWs4aS3RYroUr1RiGyCq1UtTuNpAEerzuBzXxSxdMv
CqAM8HlMoVb40KOXCVk3MKmyB3m7MZsIPDtqx+NUMTLBE1g3xIOLYBgHFoUts1mz
cKGz8LaDEP45ybbyTT/6qYryqUbvRzFRFbKVKf4Zryz2CnZj+/qKW1qb9GIJoAE1
3xz7h+Fy5cFlih2+yPgXdAdYNs1VcYVtmcKHpE5LwjwkZLgoW6B3+KgIjUT4uFId
HpU18Hubn2Q84gIWdTBMOWHJfIu81PEu+u7lL5U8L67JazgeIkmp3KbWRby5dGib
25/GVCiWQo3MOUj80QKlJPEsXxsQEshdvvGIr8FNZkrUIkUZbbqE7ftUkQIH7MhS
x2o8gG3uCF5Ye8+My05ka5w3frFgtyQA9BGS/UX9UP08GIEhfYu2I8qVB/w1ZkCo
crieNcYkwpC+zelOjRGG6AB5pTMXfS3gyl8wz3D+2ybNhRiWf4SDlhXlpRod7vsr
BwvKh3hLQtiVXJ1PJGjlYNHjrg2CkNsggWDePV6NmfTHbf/N5QAu2ToHAIF1yKD1
tIgpZME20wUZWlyZAMx2lpRjTDUdqKUshZFpf0qJge780W67kbW5hxMNKHIwW0lm
ZEwaL//Q+gxalTNrWMNCjfcu6QaPbXPmOw7x53WT0dmj5Y4KG98SYBFsuFlVa37y
J5aT4a35951vw5YFUfleaj8h5hX6BN84xzQGfBCNNUSwwI4AqT/Q4sW0n285JGIf
AVh4nY8NgKCT/xlVmbWd7qDz1spC164rkD1sNBZLkwGtVnJ7naRmH54r/XYtrSZE
7FQQ7PLVb/UFSZPWYloApkw5QFTVk9Fh9FkciRpcoG63z8Y1suTNQDtLORAaI1fa
YBLof995D0dll2ZhO9mD0eLWDyx6dTt/MrsakDImBaDwPXCvdAcYCXM3CZTEy4xH
LFu2YYxg+BTEE/udRvVXuj+Qo3lrT2FNOJ69dV2kZR6qO6INgyZlPUKZLr3qUQ51
DxmEmsus7VorVG35AwlSAF38Wj1VMEOxXW932FGjcvG9u+/iN0zIK9iauHOAz5aA
lz73QIm1CA3tHP4zStwbKhnnaYglvI/n17F/BDOUUC8nA+sGjsnLDMXbdr4a5uOC
94La3mAPYwub6cQrAHmbGvCczbQwC+kvkemQ4KnAsWfq+DIj42MytCN1ixDvwdQb
Bfgm9Ft7w0gxfScPTng+KuB7POBbxxs8C8Gk/x7h/55sprQeLXTD2aIr8ER0LMSH
pUrK50i6f3n53G5pKehYTqwvYVjwXfVvlcmKIc2vD/YoE5xXQ9uwOW2nqiNSi9it
Vz816XIdXf3H6ls8nGV9n6UmL2d+PmEu47NICZeDCw8hhDxDdrt9q4URzta3bXy5
owPdH9CviNMwbp8LEI8wfuVh6l5cuMKGTnwyFFlJHO6ynkqGOwdfCjLeRogYPo0/
mYvkbiFQqrI5zcPyb9KlfwyS9si7od0/UborRPBhRlo23VvpeYpsgVrsTkaCY6fM
JOlXKweHuXLCYTs54qO6lW6z10z0p06NwsNK/n04603pDbLkeQzMgy92wupiy226
6iuOeMTHjkr7kC66gyjDEqFRrRI3RAW8rY7RdHLtMizoPfbAqnXDWgjOTsIKjVN+
tFPEWjV/xbXpFJKgHp+lsj9Ntp7gAU3wQP9kWFhyLeFA3dZyu11Z5RRkZomN2g4n
3Ei3F1tQnYvnc+s7nW+Tp2W5KNP+cYjNCwSqOyQlEXuH/aJrF/m4+T2LfMXMhmpY
zBLH027CIbzao3RtpUWTJrE5kLe/k4/ovVsMu0Cs7ecq9Jh0beBJQ/HHzAqV1qqY
cscPaw5jnQAab6gcK9AFBg9cyF9mGEAe9ZtrZWNQ8AEw7MLs9i3U+mVyiEAobfyD
a0u1nALUEseMzF6njQXpu7k35SfOH0so0cKIGTPxx7Rmnkafe6wvCtLWlHoNyLDw
SkAUoNhmGYYF1NIipwZ2mbLjy3jQ+hVQnBmWug5yDqF8g4plarc/NUqWedWOXEmL
roKZZkrdcmUip/seUtxT3rwQajRHtnodNJXML1tZ6TiVxT2VVFH/9LWn+wGOjNb8
Ec++UIRRdoIbi7ZrDFsRek/CETTaPKGdgkGypum7RoaFuq9i+Og7Z4uQn2OawzZ/
Y57KCNQgERFE6IEWlKxD4oqb9bJGeb9yDuXQupLKzEcoseDVrWqUBoALzgIeomSC
zECHw4tLXeETzeJfrIY3CZqskdoo7hFqZ7ZV7PNRgKMs3jjEORhB3PCVbsBufX4N
HBsUh7mmgPTy5beoE/2FEDL5kjDR+qrbw3qZKpxhMY/5zOohgD5uZ6HMwNRw/jd5
URKXO4q5iZsvKw0CJNlGDoNqLB+sy8VXXAxKNk7zZ3AARqISxjUiqcuwXEXtRuK/
KfNoufvLrhYInwsJ37CxHK/lBPacA+43c0ZbC6o9S8u7WVPc9zdpdTOQIIBNIxzT
GWvWYCReqdJaYr0wQjszcXC7CZLLY31HjxSrUZgr5ouJwCK3dFeA2lYAQf+rby83
/1DHa6/PrFte9mmxEaAzDQ2HyKyPuj3SiWwH15uIgrrNKBxtSgLgiS9EQv9ZJx2S
zpo58tN77CnIDzFcClP8DMf5O/0pXqd3sa7RpW8sDUvSv6YdIg0jkpavWwtcgbgV
562UXcQtPC+/Vo+1Do6ueaS3FyMMrqxSPVCcHA3irAxl0k1L+cvLoi4ZMQDpeyaP
v9ElXYUyI/CK9qcaUq4n+aI5cE74hPv8wK7M+HO6n/GpFTKZkgf3MJS9U1vCcB4f
bsdrAOGgP/oWoUX++NHDtvifG5tQJyRb/2GnSJMsHYIirqjjoIq/if1QfLOV8w3x
XiYP8JwLDEceM39HOEjSljZtki8990r6KVZGzfasGOKxGnApNQIKUjiKf4lTSGK8
P4Mg7FkadeLx0cbyW7MAsjOfuQTGykUl45F36tcEXEPnSlB9HGNFz4HNDacC1Ufk
nz+G2m3O6WRZdMNl+jL5giheYvAq9d6lxvrMe7VqEVIuvGW23qtUF5CFFMn/7bHN
re4RT3Z2LT4camT0XHpU+YdioDRMwniF03xy7m399C71cwfS5cVc7kGUxE8aVN/6
GQSpcMwVxoSt2ISSW0b0HHWf1FvQiyWlnCGJclPuxGltGLk6xbPsYBOAwp9xlYSY
K2ip8OijIWOPIfCdVrw9a8NG30C5rp/z2yFl63utAdDkmGr59TgcAUmknDc7WkVh
6Qazdbsm/wACgdViovtXTVnq8mt3k9B8thqVv5kmnlSp+L193A84KepEjCVQ1oL1
iuD/dQ1001uMkpw25PHSbHmnl0H91U1dcbcrKqNupA+h2m9/SSaOXYMblFalHl3c
G03P+4xTICgUJhuNSC5HSaUdLn5aMmkN9of9lX8ds/uJXQSZfbAm1CYl3QUG/pXr
SwbM4EzB/x+1U8iOccgIy/sviOQtADdYJCtvMRQiF8TU/pMeWcy9h91g9Ec0joEb
T9Z24UvICrFervuELawqMZAlYR1aWaZJ58YT/mVZ/AzqYj6eO5QIFEuzZnPuf3KV
n9xRcu/aatE7DB7FLHpBiYqduPmrdWKpg2ScNeDQwhpEjDfSwqonb8WWMjzBk05x
kwE81DibiPTg9yTQkh8GLkT6uz5Y2gMtOwmGr7no+P4uXUge/T8o5ZuIdPXuUaMw
IP9vCdQ35iBLJ/4cvxPAWzQfMiiyjBIS4KzU39lOtA0w472AnccuHVYhNbpYvD/6
qAO9lW5jvimParxuc++kd6KTwq2YWnWRX5dhafQQ4RpE64tCHs9/LWwpABMAp2oV
LYj9SXVtm88vAbC4gMN8wIutT5yArNvGgZ5WZuW1VqaDudlsXVuSGHt2Vs06/edJ
FYNjVeOIsloNfCqEEuMVwFIja3ZCWYqfZ28Rwpr4Ctaus77kJpZeCUaUm5WzVDJp
633IJM3mlARwHW8MJ42HLuscSYRID1Ia0xc0RUxLhYc5PiL+DZP018FDGiCADq6M
uuuGjBB1tal+ZSuVAJqj+wDR6yiat9nA5V+hk/W7vE5bdQoO8x6kbD2ZaTCcR84g
HLp2lEcOWAMJc7QIPZBbtY70/lHCx4vFo//2o9SZrMFgLz6kxWDZE+cQqEfoeOCw
rE49X9WDXaoEiOXdNbslk1TEWVBlj3kiHZ3rHFp9RFzOEGuB3JDa6gl/N0CKHf8q
ESItQbkLOwSN5NB+XJejfSx5HhZ0SOpHiLb1jgUcyT0ieht/1RpDP1SHzmTdo+KR
wVfcHoRhrQdCUStCeG5SDX7l2vTzopwo19MbF3rLaupgEg+Y6nDTM0T8lvIhFDY1
KQeGkYoP4Ye7smJ/ul5mCyECqIhGKNLxPa7H75132Jj3trk+wIpKivsWQPgST3WO
MBgt35d7ZYLnJUi/3shEw9MIud1bsmEL/m5BWSEfscrhuGyFFgAFQRijeseewwaX
D/JWjLxdz2Mm/VAubmXp8UvF8CwqVbtN1NfB+sb+imdbMIEcOb2f53nSNgujiBOo
yFcM363pEg+uR96tRD6a8t6TE5RgVuO6vot0VgXxgvNdIgM4oXouITmYVlx6zc1L
pFY33KJwI4GqBZ4afUYlrLm1ktfmfrUAKnVRbaHSwOU1PBidM3wltof/uupuD9kH
rgg7/o89lNpTe3ppmldxvC1Smg3HTpS/tykBioGPQbWbssng29uoKAex5ykRfX9d
bYPy9EpJt9p+vkbMMaukhVFP46jcqjmg1Vw6dMEbfUK8TgR6PdrmSjR2SKb0uQ/4
ikH6d/mGy7avx5/ISyeSORETOqLcT2Pmfoc/6l+38PUU5wx95JJpXJ39wuoZpUhX
1rV1l8orYv4wKqnajK0JeJQcNpDVUIyB8i7zVvE4xUb5jHq+ILkJNMSrJl0W4yTS
CQKk13qUv7u8KyDAWDjRkSM8Ohv/MviKnKAq71XfaY0WGUzVGIsaM9EoYnoHOMN/
IwrwJ8q2XSMeRlba+HTuwiBnG6EXoAuSCA9Iu7U6wHsd0vea8tQ4fPhfITQnVJI9
JjTfafMa07APXZ2GhHv+oaofkKhvmAX1/w/jPeHB0YCFJi0wkjgvFz2S4a1b2Dmp
tu1efaP7sAMfg0AEeaHs+u8PyDYUWxPSNbb59x3d9FEeqbTBYYsiP1/orVmJsYdg
v7vGoWLkMwASJS/0wKmdkUMz8EjyfKxr3p/hsAB65kzdGdph6PyAlPtnvAOULymM
xuylIHOo6Dt6osMldASDfP2KTfBXvafg8gwVKI0zc2zU8otFB68x8f6aAOqmkYsJ
Hq0CUwAf890r2eFprlhYvjPLLSVe9MivRBAInNDbsQPm7fmu1YsYujxjwzlmY5us
uH1ywKXuTnDR4q5cq6bJutRRAQ54wuMVLDlXOCi15jq2BwaB6BtwCuYDqZGinUYR
2NPsnA6hoiM/Xb3n5qmw+xut349ZEbPsIcVEsmjZnZ7LTidoWRRIkzyB/hvmWwNx
JJN/Fc45Juqq2c936LDUKyKkRKRgFMjv4XQ2nARmBAnISYeUQmPKZfxNlUuiQxRj
jbYk8+NTdWw9EgqSvHWMpP/5a5wkskQWyEfcdG9F25BM+X3Dglv17rdu4Mv/uapN
D9i0x2ycIEq4hJ4WWqPBP+9NFz1eyBF9nAXUSy/NWuOMeAw6dB/tzLVXaIr3Wd6J
UdfhMouGEP+aLgP9Nc4OkmByFgM8DtG9mAqNqCa1IRcgwBlI1bG0tLUpZMsxwgkv
QCAR4+jM98k+dC6wvfW0pYcFHc1cXGBEObfk+TxhXpGMEGzOmEHF4Gju4CV9jUmJ
madC3bUDBVPeOyJ/qSnAaZBLqfAHHKH80Fa17dt+SBaaAr9xPICkd03q+Jd8d0Fn
2E/ubeScsdhlWCo+MHqgPcFCq+lFd/T/ez41DFHFZfnUwNZr6rROc1iw1gG5dVlC
rYlp/1VFMSblcod+PgSSm686Pf++C2cGK99hjv03OaDEaKOLKhSgjSLTwpWu6nrf
E4ptMYFafCgs5R1rbvP3WliuG9God0+oFnkW/dRiQkL4ulxiorX7JKAEebwFUlnd
Z8Wt8A0qmODuqvb1cYmyWZ0lw5uZ9Hkci1j4BuDnarpaknZESZKFQYD9EXLsVGkI
bUl6rTXM0qHWk+hKJ+HhPuiNaXpw/v61w9mKvJdlQ+hwq+4TnrmOk8lt77QZxEld
nNaI26cWRtHe2AuhLzYffUS6QDvtEiA5aVJ6HX9/RXsJIVmCiNcKF6ozmN40H1tr
TfPsswVAFBlnHOHgAPD22z5Y7i+y+Xj/YukTPiXvev6LVlCJLdYnE5PGUjN+SMMT
dz7hvnNMGDW8Ie4VzDlYk54/Pvchdmxke20+Pz+f8EEy0u7Wt8BeU+PovMPp2pK3
VCNSSgbGt2zGtVMcQye0T2krkGcC9AFsIMA5Emu/oyAOhBRpK6lyVM9JtWcvZT6U
F5cBcdHgw310k/u5lzm9rcOuRCB+csBnrTQYn7b1kDmDtE3n/C4FpicsFLza/ZLw
2Bu2z0EeXiIcWD7zcX1InaagjLl7Z1Ur3Fe7pNG9kS8pfzclz1GAwNE4EiT+ViyC
wDXugIIxVPpthn8xftkk4PTyOokuwK75ey0dkNwQmw5FC8dhVjZYAgDRZhxVPcTL
rKKqe6fPS3HF/znOudmtu6P4vDSK7w3HmVpbsErik0fNMfMjVkvHT1kj4gjlHvrM
m7l2LXhuHGLqrH9xw/WLcI6NTfZVhQ9xExqb3naVyKx0GKyett39atJyVH/M7m63
ZEBU31381gKylkwzkKpDWIa4KkxnIYNKPqHFRIX8UwqCHmmZam9JuJD+IHv8gIzG
ZkOJTN9Jo4NJldSDyoJPXsbPgoybxgKxroisNnqhtc4n2lpmW4xn70pVzoMW9a3I
2VCi6ph+/xaKOf4Cdr3zLM602gCY0nRYLMLl0MM5UyhRAHd7e7lJGnl0Cfgz9ZkK
lp83Ztt2MI3MZPRGeWbXBJXW0NHX42gweRCNhY49OOF56EUmCNp2hKiU0Xf+Xclq
jk0Zly+kmrEdSZVvjdrN5DvYLyMUpFi6QcZoa5+ZVBE4eX+twKc/ouCXuIUnqoZ9
0HigXlLCqKJJsbZo708RNWw2+E80eRDIxLaXNNPxvtdQNv5dtT3espaooLQBhTRk
4yr1u3pdq5+QPfVisBFlJKspTVCiXzetthQ1x2c/wbGxCUqkoRkEN3NxlM7Ldy0V
VzqgIzyS3irNogNSYquECxkQ2EhR9pTBHdBHXCI7//Jo8zF4T6AD+0MihDsCTcCm
cXoE5pa9gPEfoELCScBLIcmB3HMWDopYwrHAcBLJwgVHc8EmCXl3pJmirUnh5Cas
gwdY8oNiX+kifaoDFkUvnPEBL5sSdBdvo7YM/pp1EBRIYL+mau0e0dFyhL9q0I/v
ARq2XRJj+mZJAkqp5HjtYEic+/ZJACkkcsa1UG97N64kDOf7bgICnxSpaaQaaOIu
jzCLCR0hM1gAvkXVKV30oSn9cV+pb1o6M+a7I+ENYKHrz8OnuPegNzoIE+wy52FL
VV70VTt6emIwLs/Ky+3beCddXoFzKkIhRBSNYzxVnWW8Nsh6EwbndShCq3Vw7tGM
EdunIJPpJ21upRpiaTmb2XBq3dNGVKH9xB+Ye/6yu6cVZZ+jxag+85g6hQLtoaRB
gDj+IjJzyEkWwNpj4jkFMLGdiR+KamFikzla0Y/G0n2E1DVDxo64jn8gawdHGl1Y
7APBXjEqwEOWhQF/QTPZurja0elJ9YPR4ELIr/1yVcE0N2Wgi/PyXTmYCszgUnSy
Hc3N44JyQxytf5edMOw5tPhZWocmtqrySgpJGiRNZD7/3586IrQzB5Mp3flNsJWG
EkkjYcleQfgGwS6IC0qAXmPKPvs9YKYEynFuolE6GNqUjvvsPs2ZGOCPM4OAgLAe
0tAsxxpsdhDhToH+4uV9bFtqK8focVIObJ5zhtW3pDtm09DABCUMeISvSdpDqITe
G3/xAA7OOxy4rjDtOXkDBJzVPuCu7mn8iUrjx3YoMqYJNDhzyLrkup372lDxFy2j
PMuQFWWH5cQg+JTPu3rTcWl/VzDrveTRQX/MyoMwawhzkCrBk3sfm0z2nTcWfZ4w
uUkdFGzFGfGfwG7xmEoNnK0nJL7XC2C8L3KY1qKbHCaOE+lo0tIryW4S6ddkUC6F
G33xLrXFoVs1yCQjNbHNGM/yMLjGZbvtVQvRUER5pWJQi3exxUCe2rhzfxt+UHir
gQ/c5HFyS129LfBD3sJBSnRWnsVyKZqppE6ppznUPv1KGJVxcuLbhpLj913DzF5a
7js9qavkHPwHT/KmhxAB8cIiEdKvzcDlpVZtwd/B1SuZ9HOVUOZ5VbpnGb2gYIJo
NnJ7kHKItxpb59cQUn/7KQfsj5Z6tbvcJxHUch4MtTHx0oOIUeURMBiP0ye85P4W
VJOVNZNKBjZWTURtdZYRfPIyraAJBf153ENajORstVis9H6imGjoija/EBtvdxXO
W01GyVT+Lb9KyKFhc1DDbttfAb47EQwmqf5CHhPqEE5diePkklQjhbhdsBkSxuML
ZI7DL/49t0y4OSPBoUGeEjM451sr4JixDBK1ZHhEzCVUmYNk3ZbfpCdrCA7cO9l4
Xs2CmdrtSKYWbwGp4qCDQ69y5CrBKq9seqfcamIQXFeO43whwe7i0y/NeEzjiX0n
JZ5eJb15qbMuI6ijfEAFQnuOP56tfaoyaHc+mYynjjQjKbd9VSz7txKevepNFqDK
cq+r9yiYm+pbBgCfpbFnoMu6K+ZAQNBQevz46XZDrEBmWRfs6osz+V+3jK21zrMA
xBD77Cb0XBHE0T1L26nR93Y1HxAcpTGACO84Fj/kvFjOrsb7kS2uVw8D7aFWCyL0
iG0790Y/Fs1QU/3WazzE67r9OMVh+qDff6cuaRqlY1HxW5WksK1tu21dBgpk+RTR
LTAJud4mLHIBWiZpXtEZ0DmsPVuPzPp/4NmPgJtfkLlOOzodI3ilb0IaRN/pQ3Mb
FHDOwDUi3AEHeRZv/neSnuZeA7k4b9cYBQndF3WTpZTltT6EjQPd/bEdyj1NANlt
L1Nv4re8bhGDutifQXAStL2FGv7FAtSCc34Ew9/OHsktzWzxZAInpqsi4reOZ2Sh
S0a8WOF7Hd+v12UoX6jqLJ51lqdjbi23R1vxCo1GVybRZMUpLOyRzeWjUp7AV1Su
IplJho1zyqJCxohNDNUIiL9oeUBb8Iv9JnHG2USWcJ/lRPfuhi7AeQtK9sOYVC7x
4xUkhdKlMEuuqromwJC5FyXYUuh8+fOcoKhsv6T3UNHyAQaYZhqa00VX89eG82bJ
AKfWJcJfrEyHEd8+B3O+PEBuDHhk2yHqJZUup+nThL6eKd8lnZa6b3O3iKFulHXT
Qp5bbqh08MAIOw1QKx8OpS7YVq/Ik4sc9DlgMhzPusc+Ce1euZGGkkdiwKjwTci/
AfajoDIKTphiURct6ur9S4dxB+QVB8nxd7Apx6vIDGlD+8HGG+HJEoqRSkVaz6ZQ
SIyGEmQc6aABWY+1nHJWJFvzSwgfEcukYUiDWJcx2u90YWxhQp7tPayjMktwhkRf
ytbWwh09rrlw9rRfqU5uxgFkZ2f7Ei3y3IqY29XUSNUbX4e0EKCDspw4Tsy0mUNQ
3B0nTOzNsHdDlm+1QDc8b4z4LlY8q+FE68YaXplu2rpSXYPpBYr0+9lPYJtvBpvt
PqwxmWVitcf2jGtB+XqBYUL4pPCBzp+89TcHdcyAVQlANmXafWEEtnemnaZiTgbQ
dy40ywxcfPZGTfDHcRhKSuOfg8jJBKqbuH+O3IM5bXJEHN2phGZZxCpzFf8SNMku
e3VXGtuWiK/i0IGHVBQIu3hPs2xBlYPPT+X6vLmi7q/cxOwr3/c1E6xPS98LCBoW
ug3sbQ9C7AiojFBlPcrcWW6f3dkT4pF0K8R6A3WVqJDQJrFUghJtUUz7Qa8LjXBx
Jh2GsIV8UMRxCMO0V3lIRFkyTOf/xdeFvcmpkZje7F0EB9o7jaGNNAwuRvDlArua
xYkw0WCgnLmnPm6a6mD8Z+nNa+7GT9Dj66gcjGvs3gSJH8GsADsZQOwrlKFxCn4h
zJ0MLvQ5AwqMayTnfFBaod+5LYTtjx7ZWFr3YsQb3i0iyWYtETX7FftmEaeuvJFN
eJ0yeVBYknSORP5/FNoNf49zwPIGWAVojlV2aqwUXMyuxBMI57RVOW/emngjFH/V
fzLSI+P3xjAkWuJjCrmctzlMtYuEyTiccfHqBLKPB6kdm3s1Za9jF9/qeLxB/hFt
AcAGU0ByEEEdhhtVJ67eJ8bkOrMlh4mjHZKpB7vt3v4u5DIz74nzUOlyY10DnGlG
BXaPZEnB98QmPI8iEM1/IHPxxdfsHyqVCXx3R4NL0/tszzP42GIOKpo+y7ixPVXS
5/ZeHlUJYGph4bT+15RZhx+JnBv0Bmd1AuJ2sEoOBTott0jKiNpSW5GjarSQknk9
klCi7DfkbBzBErZrfRW56DoUe2/6sFd4IdUN335G/fZ7kEU87APmKtosHsyLrXRp
PJ2Hw6lB7CUBQgeFj8B4pwMLVpDDTfzdge80R1ixlPB6p0VEpTwvw3dSKrIEFnMY
zfxGEtlLOOKNnB4TheO27g9qsFwIa8oDA3XHrZaxWueiJejfW12aYeqZZ8D+KWJb
o9nJ2/+pfOxxi76ioG7U44lrJ0fuLFdNUyBa2RB+fVhow2cnqaMR4yyJwgTi9U4/
BKuDh+JYPiDox0iohzlRDOFmYKwl1Xc9yEOJaWXUO1psrfOAtXlke6Z2vnQGkXAZ
TC+87HfREeeOj5SBP0QSG35I+6F2PaxwMz16Pqz44tMIg/Rm+APH0UMm2C/6WEzf
2sFO/TwGElU/EbaT1KKQNOmhUaXcVjoCGDcVp949iyCzcPolXcQvz8UmBwp6MW/L
7dMFdDQSlJgH6hT3b5zMf+c0/SdF8xKEQGw+B9k3hfzJEt5vGYDDNJCUnqr5E2ok
1TDiA/ti90CAzpNM+DKfvPbgaztIUvMV7c+4WOc/4FwyUXxc6eu5Xgzb1l6DWetp
OhCQnHASEoS6VcaX0xUhq5DbfDgNrdZX4QdTzjGSVjwJvx6MqJTxXF8tsyT+f5HR
N4K1xW7qYPZ3UDrh1bzta/x78bUT2+j2YPTDUZNvQABmmJxZPS8Lehso3Eeenjkf
uSTzF5SjwG5/8hHZqHAJ7Q5CC6d9SDHlNuMK8Mr/hEL0xkUEAFyIM2BBz/tajjDS
HOgqT3oQoMU603VwJB+tmBLtHJ8+O6bDLSu6OxLDkMNYZGmkqHt7rTeu7JhY4dmd
MM0extk+bQtaF2+tvBGJcY3ehjX0FUD6izmdymZF2hYlfmGvmgOT3xFVeyM7MTtN
P++5TF1W1E4EPRU0Xr3ELfPlQ8kTDB3EaxfSc8HjHolvPFqIx2g5uqpNpdsxrmNd
nlXY0/ORs+u66YkMvFQzbLV9kAn8NC8KoCADIEEGwpZc1DlExYZy29R2OvGWPdIQ
3m5R9av4/uIQ0wlyQ5d/lrmR8Ojz4dHcC9AXDEFtplcsxp5ZGeu51h149aMj4/G1
3Dr3FPlBy1aLDuOjhbF/4YAqp4Ek3NAGuXADdv36obJ5ZSMxmFt8m0aPgOuumpQV
mIPpnzpE1b2fjv4ssaTZ1q9/jM++KKLKdMhBll9Vv6J6ul5CJiQVBZGW6+F+UcNm
ub6/Qz4ufM7cAmr7Lpajh4q1CwnL6NaiY+s5s3rMotI3SdtlYUIFZooCZ8KIFEnE
pNAqlUx2fWebM/trqJVurrnSfSyVpD9Kqje4x1V0c39KuSVcT3Gzgr4gKwPpjnKP
YpgqdftR3mcpgYI+HJcauz7MkJPDTdLjIrkSd2sLXasJBI6zxmmILrUCRFHl10qJ
HHzST0SFjxlwCk5v5SKi2tehT732ykHcSUjjUuxKOdWY+Ez9Er8HRutU5MTneFOQ
eRzG7TfUDPId3gd8msVqNGqYlwYXBDJpTEWdL7ynXkokHpvCtxWPCan8gfV7UUFh
EvHkTg2t2H21nkAhvMActlVOD58KsxsHpUMGN6DZbLRimcjnDrr0MzlM0w6nOLNI
cvcp8vGptmjvoMNSlyOWhum3hms1gbz/PdRTscqoOI3HGcv8RpDxDuPPktEe33uE
iLnuCIYSAO/Ede6W2iffSfJR93hXZdMtHQQ6ZQZoFzsbrJifIEW4wervj1mQDIv9
jLCsbNCgqZrhkosLWVg5wKs38NHgmulDVD78VFFzYcs82gD8hdhdO9vdVWsmH8pi
GQA5tTE4mEWNQGKLSb8wyJviMG7XYbI65J7gJkE+DnRhJRpqldijWGQCpwTi0mRW
Z7rk8edRMB8r7Y/8GT1+GxrElf6AisvL9JrYb+czDj6B80C3NQQFOOUdyFceT2cK
7v0TdVEoSsjRtgXsTM1I+HS/lRJuUJGwA5q3+fxwS3P/qbf/Wv/y538zgC7Q7/HG
klgflkUHD6SrcM4XIigHvMIZOe41uI/7NvCdl+SlPICAD2pyEnnx2cqb9YSOVGJK
3jPWqGzRkuPEoDctiRAOzVFVl8VXnrZGNJbYI7+v/R4kVrQYYtvYNUItRo/7pHyq
AbEh0fjnTn5LPGVQ89iYzt2DnliVv5PKysetXjgXEdxlZ43Q6fSETlRmunfB1Gcr
+M7BFugNpFiOZgPOX/PnWbVDvEKH+t/QMsvwypb5xSzuFJ9isZpEftB9CK2QQKGo
0hjN4VMmma+E6O2dgxO3/B6Az4Qi3X9qx7gqupAK2oMzqF9qvNAeRoLZEmdQ4MZF
quYd6A89EQmwfy922A8VDYQYzZXyNL5lDNAibSrJmVudGsowmWnWAGTah4HYLXYj
MGfuZlAOWs4gqcEKsXWKmebnX5N+agVak+0S8WzfZnLY2JzTh87SQtOlqpODDYZ2
S7KNPcryOyfoU4s7UQBhfoJODr5lUP2xaxQamc6+yxKSXwlTRQdYeIlbz2Mwy7fr
s4rI99SR0r99BQlTijiOBQSozORN2NFzRBZGHTRZb/GlG2aCMbXrteK9LJ3dKreW
/Fo1xKjQBZ4p55mc7H5JWH228clzV+oecj3pVRO1mXEUo4hoTXVkzhdqINoidJTM
mW7+jGU9Eek1QVe9GZ6kl2uMvkPwwIJmRVSXRHufvQ8f58gv1zE7OBFUlCZfxc9H
2Qixqtx/jXKgQvOW40imYUY6QXHTcHRmmYbycVeylyTX/n2vvK5/PacTadQ3IOZA
BlSeKuU0SsHcMTsy5DpnATnD8qp16hIScsb9hp084uU9UVII9NtJ6Lol2p58T7iF
BvvF8Slu1f3Z3jwWFFrJC6uQERfJ1ne1Bwzt4dg1qxybzkz/BPIfDHHt9YrVuh4r
vYhfpzbP/uO25QGAWZGVCFt7dXiwSzVsAJMQZX27Fl69S1EKDSmA1/b0qhz9J9wx
KEOiHACmnvlBbdFIWa7d1x9P5BfZRcSta4eXqmeDrYKw3boqpMphMNWhRsJVicGz
C28ZLr42zsru4PY6HPpMfgSlLhJdIeQT3Z8CkOTyltYDTzjCJBdLRxdW/ADJliQt
EEUwmVE+NMyABFbbIyaUfFLOprYoWpmLX3oDAWqgVmwSh5jErpEMh9gLVVe1dvBX
iNVhD14uPAXiH6TKPFRZb56fdfL93VbbYNRfVJkN9EZ+L+bi4obfqWdV5GtEvLNy
ZSsoC1aWYcC2l0cr7jUK9Zvrdin/fDVKBEyn+TOPn7v3aneUKEtZZeWebGWqMhy4
aS/BEwyviKIhtcuNsIVuMJUxbHLCIrNScVYgcIoaiL34cioZS0e0ptpXR5O2Z/pm
x14PNwGw+oVDR+0dkVL2QbQK2ci7rQaxjh6J4tPKHpDgiaqvsxzTU30D9JaRAvd4
GSNKQh/iREObXU07lqMzQ6kBjn2Ro5itI5pglAlST/ZnMx8dihF3k1fc/2d1PzWM
8S64BqP7rr28EDZsSqdiK1i9U/2QyX81hRgktlYNbxRlEcjUsG4besNhE5OI7OnN
BSBIGLHyM992iXg0uuG+CF17g0/2sQg+Fm8bGrm4SKjrrtGUdqjeKuTEnqZs/sIS
WXo+02isWrATNU0aiWEAR1yooAQnSoyXM/kWb8Con9+3t9bVJk+uif6VXXbD7Pmx
7OsO93bOWJlaOAzgyk3+QsTFm3GpL/+43lQ8t7iiZczCAK3Zn4+pdqpsXH9LSD/F
1WsoX1/yzlfxHNXy/gdgB4eknuFfNpwPGi4yl0xwbvGWxNPXq0+ILoZr4FHO0ghK
INRHB9GhGQwy+jcQ1uKI+i5yVhl/kZydBbkEKKe57CwtqEvRmNhhEOUps3Jw5prc
wBP9fkkpWRp1DOHunknEx4UYYjTZuXZ9CGZd1ZhORj/Oy9pUvewN/Q2+h+5XFw+o
lEDg1jw1iCAzELebJP4OE9m988ms0c3whhUP6Js9aWqic0Evr9Dk0BaPh/28o7sv
3b92JR2OP1scJRY33f/XCD5h90Rt1MUSNgSYfQ3s5y3WytYAd+Kz8uJ7/v/ismke
LY5JO0Fu6DGxde9f7CFxgljEvXGVaCkUYpovOLziFecLRPi0Uro2Y0kDFKDXKf1/
5mGVqwO/PLODOWMo9tEQzO9wVZy0iDe+ipREokh2Os5pTfLWl+NWOqFIw+VoeX0U
6pXxXw2TKAo/nIMg6VhjYINUxWNrw6ft/U+kUDT5/TAZTGVO7v363h8YMBmwDb6/
3G8dTa8ojToO7w65XytVCLHIb4Mouq4LabE1il8R4aRuy2FiT+YYiDf0X+43OxhM
3qV/njmW2/mnYnO9sJ/XE4D02VZLSzW/mV8zLo7Q+qI5fGw1PxMiK/kRPxxwHKMa
msvGVOVq5iuSDPouby9weMnmOeW0uMSoMz7VNzkTRbJXXHidm8qCwv4gZlhnXH82
f7Aoe0JRbevBAWCgObf5JsFyoVVF4b48tO9MFsA+TWzYsA27p+82hpMhpBlIQ0GB
+UxcWBXk5JRFc5x9QTghxW6iHRH6OQFiceGfE/C51uKUmWHDmvFPUD99TQ+frGMP
IhXtuIZvbtmLZGGkTAINfcx3OQf4LE98lfzVCEIduKAhLdi5u2W8oOp+iOATx+k1
eHZoaYSdypCrtC1K1OV3EzkBCG16VUhol0TshmIlPrqFG4oaMoKtL2PQPvEsLfwc
zLmNr9lZ6zdSfAIRcqsZbgJ6oYRwKDzf67vWWVX/iIYGoSZCmTP8Ol4e+bLfjg9y
bDsuLYhVxVRvp8sJfxs4wPcrix4975tEV0BlMUxL+3mdHUaAPqfBy9pvBCbAotLD
aHPm7Y2rgLiA+yZB0q84stZ4P+rAznzApETCqC4Z2XUbvp6dQ3QOO2CaRGq3Lv2G
oJbL13HTB/I2LFdXmp5vc0DUB9od8LWaM4YjYpGKg4avbAPagoQEYQ0U0/4Huqpe
Rb3X8KKuuU2VA/7D9I3mo7wIjf/WjRtIbSJVkuy71luY2N3hZhcAyVKMnZ3W2Hz6
3UtaYbIf/z1yMZT89BecRIM9EuaFshcQ4YHC404BNOhAEY0K22EDAm6BcdD45Zmb
zPtGTv7UEJGSFzwZdhLwyonWS/vCy4GS5FC4mYiVd08xaz8Xiz+iFLWvZjih4ypk
nLV2cssfCZQSPUo2q9wNL8kIfyTecF5CgTDjvVP65jx91pnaYTuPq7IrPZ63OLjs
cv6wcMbcl/qodcnAkkjjSvkiZVn9z8eMTb5y38/U9i3gpq32bohfTAc/kTKGbBQ/
x5iRODOgRXV2mVae834jEcPcibA8vyaeJAcp2++ZK9pILTyj78ifWUjSSXdG4LGs
wEagjGLfqXMONZQQa0fePXuL9YPe/qspFs8V3WfTNmx+QN0qXCnmdG+dbVoa681f
IxjTesdcEBz1RZxn7Mv6wNiJ/cgSmkTBrCe2NbzqI1w3GJ1HI0HvSTsmyfT7dKF4
dlim10cPfg3QW45HzJzG270Cu/qWlJLflN33loBcQGRFTIBDHbUUSDvHD0jV+jyL
n/jP2y6rKKPlmBSUHYHvLItIj1np0dYK4BHcuumdLLzw869eeDZRv68hqBhc/uSf
Gcq5mhma5wtXcWpQiZQNUwkBYeR+DQaiKwUzXFpanp8r2d3AG3U57nmII82KmdN9
WQlyVbgojEX5M/muDANVjm/tmc9nB6lXhxc/uVq0MFsSLFuJ6qwIPm/j5R5bKkWH
90LBG5iDanauVlTRQ7VnSyApJ0N2Jz03wWACCZhy9cwg0gHxK+6YbGuJi78Y+Rvh
UH76ta0aHUZk60v4rTSyVe67JX0CrXWRUNi2dEmrihLm0/V9H+xdfBdHzUt9TSGO
h5zUkkyMHL7EkO8u6kbsh5/rffeLNfErG2SKEnAvsoVFVnezMMc5xHtNUhB1rDAS
m7G35zeKxqA5RPCpO0IkJHOgN2C5mZ3KxJI8/CVcGOy49vInW4RNwGTUALAI+oAR
ZVbMpTwA3OBSjZSnsHNAMTGCKZDg/EeVrJ0eX0GBN3TgN4R58szea29at26042Do
RXWeJLB3ne2tRe05SHYOI+hHmGYIRJ9lf7mZBhZu/k7SJ1rpYHr3+cnRtbhuk1z4
5S7cCFLHrKqd650xmJKgo2XTW919KSgDAdq3eOboEEBmP/6FiY68oeTn9UvmWIj8
TGSxB8blT9mNze0oRpT4aSLEdgKmeKgdcwratc/9Stq47Gor+SmXg76eRoYLp/Wv
c+uPG56vvSnQKR5dce2gL6FgIE4m/VvMvT7fTyj1AA2n6k08qiZR6H8vj6vjmfwx
zzFHNHWwJ/unL38Ewoqk5gG9xeV464XjuuzPOAfPhBqlFKqpFRj+azal6DQP0kBk
BxLja0e+/IMPrzpneohNijoKkEjczdCs+6Q8jH8CqtT9D9fjdmNyqRAM1YJzrW1y
4b/+cu0WkpryaypABMxrnK4qTj0ZTmgMZDFHiSoIKzw7HrIf1HMeBsp8fWUFpEyl
MvqZv9A9IS4xopBEQeMuCVARptX2/PGUa4BONkHDnF8=
`pragma protect end_protected
