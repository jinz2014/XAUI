// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TBmHPICb66fMrpuXZAXzFeKwkyA5f0ogvFPDurr7BfEGSUFAlAmpml8XwC5DjnG3
KwdS9b4VoX4TIqEkYn1GO4L6GOr8jXK61EXBmsIebKGOiwQ1saKRb44k731Kg30e
biLa95Aa1bh+pCZDBIjsqVnyykt33OM9OEV+WhwII9M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6992)
bpjXMuIm8JGzThsIMXiQqRYp7AK0YVhcn4gXHrYIcQoqzbIzJwPhEwGMCWkpT9c1
kht6fd5Hd1ib+dUFNc+covTg8RpEQMVQsDLWhU+6u3yLxUwVRxJJJ3aPD2a5UfbD
HBKePr8HmtjCxNhUuSTT/UZR83QwHlWZ72R8yqlML27DxiY4sGwLXrP6SMczoX8U
pMerpMh/5yEG3Hmr4wI/KpakrmBYQfiSa5tVeGPPtco+B0YlI00ENRyllkQkPasa
/jpqvK/A0JojxLslWLOXtF8XhBWLl2iggbdgewgzw7g4TKgTwxCv1wUsTwVsIz4o
TY2kze6LnNNnvuZ1ltD2UfSfl6C5mx+Tt+rHik9TVkrRCq0u+4J4AWTl9LMQDkRV
Qk0W6i+ytYfTKo2lYIcN6eioTWFIVR0T2zBBjtzYBFxxMbph1a0mlf2cJm8nJrf0
gKI+Vl6shhU0GNuWeU0l/fErW/JVKsjmioZE6XbNX6Erbbe7oJ+14RO+fMYR0iRQ
/WPM6K2gj0uroLQHv71ID8gG7zgQ3fbCUB5wdP/2QgugQ65NzTKfASPA9hAGrsHm
ze/1whoOjGj3RFFbFPUQhJ/e1WuM62wde04PHVeDCVDhHc1JX+IBaUR0AmEF4q2n
nQSI6KhdJxCwGSEjr03U7dHGV0JX3TuC7Rk/gDFDlCntFokhfnqp1FQWDBgrpDbY
yx0dtgDosK7E/CGVAeBJB5xzxv2YhLTAgcqtwew9E3gM53NB+PxkNtkMmzq8tSA4
PnVVkG6fhL5oyaAqHGlDPkVDZEcq0WAqSuarsmBLBlKcere9UGYXlAiHGxjJyOp4
cFbF7UPdoJmkKfwLLNHljdeyk2OuBLlhYNn6Qbo0oHnPdicsnY1Sz4+UsRmRjZ9Y
raBIbWDQbczURFbd+Z0HCRJKDEnCqyuuntjGZ/roK/DSxiN2AJF9qxTMSeibf3aL
CVF5QVRqL5H2iaflVsgC7mqwDdoVpmZYs/lDMA7KhwWTI+qOl7KjWL6dKhYIx2GJ
1zY7qzmGtkPzhoJDU+SFaFm7Jqh/MyZWpKXkvHG5QUZyzNPDjKXEMLuIxZ4vrMXZ
9xhrE7EXnju0m1oag5/pnKqUdQgRmgjdB56cCt6H/pZ8H0os/AFMoxvH22y9ROfU
sDp81ShM2oqkea6Tq5cim/XvXBIdVw8SyLAT8SIkpZKj5psIgU9TGXjtvsrfivkm
5TnHRFEBDJkQC08IL/OyQ9pO9TZOpKk7sNjmPou8bMUywqsadF4l+k5y4Rmv0A8t
QOA3tl9lIDkZ7c7O8yTtr8C04Vu/BasBJW6pMtKskDE06FvHmtpJ/SU3yl2XeeFD
HwVSMl/km+F1kSVvDlNk9AuldC6Oe11NZd9gucUWEdTod3tSh8iPlAdQnMwR6vSf
UprzMdJwtOdlXujeWBmdKdwTnjVknINPV3FMqpaz4POKr0wPi2+aGkj20Uq+c/J7
3+sP/5IZTBUGeCH1rEMvOr5w9zmnXUbpuY1XdGEjfJxKeB6pkK3g7IQ/ZioVFOcH
xjLMjApMxfWmWrT3uwEnKLSlCKhGDYm4T8BHHxJhff7X29135GeO91cYZuTOJcvc
E9xmyDFZLcLqvQhpfgvoaqcjRo+FdvAWYvENZuBf2gwds8orNVUp0Gb2s4CF4DM1
Z5G7m5BTUZRYWdF48jvSIOMoSUfIOlLjbcxxSJDmepWuhzgmqcgGUgO4LaMjjzlM
vqF2P+MZG9Nv2NJASUfeulYMiHadxenmdabrCvHe3BprEvL0zadYRglKjd63cElC
wIUwl15XlMUxAMD/XsFpIkp6/jOsfjuSsN0qoNw2qZDbtahGQ0gQMEJARU89CRWK
uvZTD5pVX2JeDOm/457F0P4ng/EF+63HzEza+rMSccxn9T8PnMRe/XBi4TDzH/el
aVlfPQ78tKpNemp1QBTdqySaE2zuUamzcUITZKpWmZxvO6U0HVYAPB+b0MsmH16y
Pnwhf8QeBlvRNjai2x16uuCwWM3ADb4yK5xSAG6nuDBQ2f5vzfMxCVy2Yot6pGiU
ziqei7nP+gKN9kjuepQ12dECg6Qd9iH3KOmv50s4rbCi0m/HehdRIwODd0FMRhN9
ysjoF5hhoaL6mtCUaA7ZOkDLaMQJALDh3ywBeCqc8iZXxrR0TUOVs2GsEooNkAtM
EnXAZJqtraVEb7C2FtPmw9Vb0e63fziusjqDX4uvRft26t/HDQbPd8LNCtBmtuhw
5lf3GlRjK1Ku73xrMnnGL2y28bJZPM6Wv0vB8eoWDTwj56XuTqULdupKLgum5Kvb
33V3cqsrULVg0g5kwLNLmhPMaEknB8hxgpC8CeUSLramustCF3Tdc5RtbVS4GJWM
tbmw/i4eOqH6f0ZcsyCiSGOqYUrzJDC7cl1QqwSh2CeMooAepre+l7DUIm7X0Mnn
bKfhXsKMht0RJbVWN52oNVlqYUUccS5sx2CBuq/LN+CAVTT2C9tZnukCGE8wTTxv
222YpsXNyV6iW2fi8cPGI8j4DUdeCg3HV4AZeea2Hnprhwzd3+UhKA2I+498Cb0R
FIBfd0YnCsKevPCbrYwFaQXXe5+RuLLsoGyrJs2IndOa+KKF+sQJ7aeHri4x4LOi
xMSWDPGdOEOsblLsvvJWooBIP0A3jsNGbJBtzk+qsjZnhQDoW9i+AlOVurnBPqtt
RkEu1YdRrn10T15zK39nfXHW1TD3ZfLESRXtAUpWKItrzdbVNv+8OeJywY/gnmGS
jZdux9gciBf/moNI1xv8GC13aDlFcwXlmy69qAuaXqgGx3FWpPDIJBelS1zpX38Y
o4MnLhunvLgfbRFmVwuR86NhSxWSIUj/HV9oza5EX2611+8P8sDA+tSacwAHz/Mm
d0t5oq2+QfakunxdPMXiJs4gcvvt7/ttVSIZT3QAOsdcnmPf4Qww8w8m78FkJodh
fBJtd+KMW4SnVG1wqp04cPCgB1vrvf7/NGt1DpGyjFAwvKjbDv7PgqbNzgMAAfKS
EjHDy3kGAfYrGZ0fRCdKdIKXbSbvB6NFgYW39KpB7hcS3tS9cdcO9L+1mhu8IYRr
ubvfrvSaPivn/30ZJyNjtBiuK59QJIrDA9w8gTQad1K5/uNBb9BGrsKzlucbghk5
9YdBcyWi+9tUL75rDBPcSj4hbHMpcF2w61ZioTAXQ1CiTIa0vUuiSVeFtL1RCkUO
RE/VHwd1+3QN4gf/J3JdGhxFeNUk7IFYpYsgoMVaruwk2+8z25TE5bKcGD+DqGZF
+KVRGs2tBVVhFod8G+NkDTSWR6oUs7OpjWphRiJWrOoKgIunT6JmvJ01uwqPwdM5
6qldTHgd6TGsDQ311Yy29bCxV1/wbIF3QsNTKjhJhKhGpzFlBqv5QhFHlDjr43bq
UoCtyoNAAtx9BDGZAQ3J+FFGYQnZHJk2tRGRNuutp+XrNg8QEx01NuBeh0y3I4lZ
SU+ZYkY2P+7g2t/r4D1xQpl3zMuN/MTD/xVm9lUATVPcf+g5JQZgHdxx1SSpLhpu
ClDfcHaXHqZ9aQWi4PpHApT/rfHHZGCvLN24Eer23WWPJH2wF+tIgLCFjU+VdWRg
aTnHltVZIaNoQqo22vOUSQdpHQkmyzsNGXFEi9D5JI9NmWFfxPCNqaANsZc/qXDn
xrwvWHNqqFS8swG1RUaGrErfonMuft6TM1cyNF69EPk5YWmF37uyGLJSkOg3sH0r
kodqCqVYOuyht1ML+yR0UcGPkiKRsTj+aJZJmL1nj7TGQF9p6p51fyK93fRCBbj0
qdX0Zaoi4XPaa2jpJ0Ro2rybS3X0jDyMU3k5yOax7H0sOLfeRtDcXWY9N7XLxgUx
A8oZ12aj3bYyLlqSedQFn0iSPh3wvqYUMQZeDuJ+Ap0HkjMeu8eU1AaObUqhDpn1
+Q7jzv8CpPEUtJUQX85Njw/JR6FeqY1KiK4G9mpOXS2Q9WSpIcz7g/XfJ5nPq8ku
dmZjr3/xdLaEKXl4YwggrwN6594IywqV1vPTWc1GlQ/GZ8dx5kgXhumXCuvwCv0C
YLcJtymQ+AbwmLntuEjXHUEnLm1YG5pim0h9mznq0KY6rp/uQ9yTL91bhul2lYLa
YKfkm+Z/0R3gW3tAwkwI58nZOLEqkwEwfmN6uJhmxx8SHX9Jje6xxsYYX162lIE6
qgegyfXqxOs5p8IG+gkBp4WgCsdZmMFLl0RCtFAHdj/ziJQlHEcadvx7SozhdEbN
93Se9PdhkwYUFLBbhbt6E2x7sdoITqhD2g+91oet0KwbWxcK/Sr7aX19LaFeH2iK
SEY7beXvGh2EXjNAXc8PvTlMHU6aHs2L5BlcbS5c1Ezj0HCnD5nx7l9+ji4giZ5q
Y2Tum0DpcbNzB8wkX8aQlMqWv+7jltYLJTxU8qMj9cZirV0BeBmkby9ExdHEPmhh
ioBXP1QkvBHCU93KJWtYUkxKHnClUh6mSm/R9qVc9FtOyzr6KeMPMWIG31kixf9l
Q2kwbd+TCHY6J32CvPzq1pTBSo1MJ0TRi9fOV7YN5rkA/klMZOLkKHuEipSbEVT0
yZ7t/5oFcCmFeym1mBT/3yOrHNzRBDshHjEhfueto9gzE16dCv/BD5lr1bd6G6tq
xM7hdAI9+jS4I75pWOr3kbTBlluuuUb7psnJ2p1/CUHru+kJKlyaVmJlP6S3OHZe
+WLJ1OxOXxIUqh2tnKKG/aO3WT1WbmoB+sOsLaL+xFYnf+fYwKn70Evr5QLXiBvE
YSkprwYVe5qG25YAw1SrM4HyocJDLM4jWexIDy9S9lsiw5nC9dAIp5XHg6hydfDB
GjlXlbkDNw6tn4cm62ndFVsLD4fyf5r16HK1RDth4M9huwv/K7c4M11AdqYksovI
l9XA1+hxWbE9YQBDU3IvZRSK/6Y+6lVXXuU7sEfNe5pnlnuWI16IRRB7zD+cBoxG
YaLDbDYAlIudANEUHLKcDdZacpOjIp28oOK+1NJbEAFZooOUTzt0JgqlYvKl/h10
AhwBoxdUx6O0DpdHlVP3xjEBWShXJGu434NueAHWsozgjI6MJ+iHtN6oDO00Wmce
ZCbneHTTRqKPH0NwBPl4pgMbgIaxCbtNbhRBDe2M/mRJQ0JIv4jJowLAIvz1pUu/
rXibv499DbGp33L4iXuSrts9y8mTyicUJUWqf1Z/3jwAxdCbf3ZNIL46cKiZrgJ9
mx8Ms/sBju2oDFuAKTG1XH0CVutEsY6LvBI79U7GQ8F1BDPQbqHuaXpBEncI0U82
ruFVJz0VBvPVaWoT46690LJccOaGp/t8Kwd5BmprsMUcWuh7CEVNBSB7VyZsFc/5
mza7VHuLi/Dc1mYHOxN0c9yH6HMkoM+dNwdwGUPu4RypjL0gWr/FJzVMDx3b4u4t
4T0R+JHHuToF7wRyATT1iFWnJUnOKt9N8b7Df62cWkNiFREYRLd7q+rCCGWNQxLU
qJ8ATigrStcjNG1DNDvdwzk2DAlSxINtVCzq//0Ec9Ni9R5kl3w/N3oBeBYwDqFL
XYgE0qM0ckXkK08Eb5HwRtVElxIoS6zTxdNDmlg7kjmeL0NpMvvKMSKxqavqBaRc
c1qMv2sSFplg6fFeeM4Zz0CRmjHNpcNV62q/DFz7oo8MeYJU70bEZKx3NUWo8OrS
K2TZVFRdd4sUN5QK5xBjVLxefLRhoQAOukLgbyTdoTTlUgQpVqh/Lu6B7X0TGH3C
fRSVmINUJUZNBm7IklceBTcAkDJluBMuYO6FisSHyEEsEEfah09esP7tOOQeYV35
kSxm51c/m/nIWLYpz27joiQEW/HCbHNEx/xr8MH5Tns6H5Wj+6yYALkbLFB+4je0
TuhB2V+Q4wjyRToI+p4Ngu7choDFbOMZTfX2Gnm3S0KWCZ/8Z16KFwCGvljmQYB9
dUwdxFMfv4JipQ8U82+zw6GZKdG6GQneKRxgQzn4Itu6tk+Ip/KmLyfZGTOFC6cr
xzGbInstSpo7YTaDF7qgeIjCJWsOAWrEKFwonYfZkbRehyfjj6HIeOV3a5gVOs2u
W4aSHQ4mZSs09JqHur7H/TWS1mtDQ7aM6eQef83247NlWJQx7fhOML9Wzi1WQ1lK
IqTVwmncFnXOfq14eSYSqZbs3UxpcEYlSvEa7s0U5IMCnZBdlJCBDuSp1U2AeSc+
c7JP+gt2/CEeXLQji/HiGse3DEtNus7aiWpiUej9kg/r9vZ97fs4IHfGuUDAcwCI
PiX6dT6wPG3SMldBKcGUynJliIS7INpm4x2gJPwIVES8LT18MyT7813of6EZPmrX
SWh0Iz0H1xelgaO/oNHTDMaykg9OppuJzgQD4bPMPjT1vcSX6hy7gAiryEwiqVpR
TS1pcSd7qta3dztgiyOviUYY0mgFUo0F7JDBja7ax/CeRO9hLtIeRCYKkp/EXkoy
VhVw2mA4mXfNOxIPoiFnQMIA2mawIlrcdU+1Ek3/OwWhZSueJmgoMVO+BV3tJTbl
mdIKrOkBBhLQxaVKsoUnjHeX93p5pST2tXlB7VIUEs9GlejLnCJErfUh+3XGdism
S0WSn6es/IVhhIOz3vfGrlmCi0JKHdFnYhk+WxWAzxpTvDCnMrtdS0ihT/kMkjbu
d+35zTRaVHm8PCHHACn4knXDJcVB9MT8MQO4aW+YEZ0xQ4+3bszsQPMu/nXIix0/
o7GBiRkTgnXzrN/SG4wG5wR2h3m/gUP7/ckfGQ5Y1+HqaLyrO6yv3jk3a1E2U5so
ksFlFkbOPcNisJqHNe+M2oQZM9Pe3Te9EccBzpM5VWUMwNJM/mlfkZjkmHCxl4CM
uNl1n7vq356TQ316mCw0R0dhrVdvRQgV6NNJaqHvCtavMn1SHzoX8SjChkhjuW11
T1nZplQaLjrgUqzXTrStFbNC9InUKCR6LXmDyh6oizXN28Nw2sTjsRCagLGddApo
tTvoC7ppjxiNvI2V/MLEj+wfe+IEXI9kpTfIAdTktAnr3ClLOzVYdxETM16lwnrs
vvFpmu78tbgwrOEgT4z9ASbAalASeiXs07A2Ml/jL/2TULA6a8i3OqnE9DZ0Sov8
StU03z6rPFXRWheOeFk8H+TyiSxkz8YyybokYWCW8CHuNa2DiL+enjum/tgGS8VZ
ZcKkpWfeuBDip91HLVWT1CeRUs/XxwFn3HNxe+9CchHe7yWWEMnyq85Fkm4gC8Jg
YaFnjFVtNlMilTSqWt6JTCRy9vtH+FejBSqhCTsHPD0Y7JzapwScwVvnDG1HtRm9
vCUWj1PRh2dn5AcSHM2Py9Fi3PJvPO++X/aZZZl1eMSCsSrUzYMv22hZlURJJ652
CMz2nUojLXJYJEPlhFwgZqaWlF+S35OETroeaD+N4bOn/6LYkDh08fO4uwnJ0moT
f9/3oTu/HzJvqPT7SMQF/wx1y5fCrQBJjKMTZ1jGZ5Z8sEicypzflI6P4Qhdw1KG
aCSOLN3neMt5VzstQwbXrqN1NcL7kjqqE/tuLxVW96VTCV//zaklFI0W1RrgfcXG
KzieDLGZFo87jktrBeUsOW5WRR1fkbmfT13Rtud2gxfHUe3ej+yvm+U6HVIVzUPa
5TlxONTw9TuKfFNRK0ytum9FFw13HMWkUs3p5vj8qCXW6OlBvbI/n60oGlykI0mx
m9FiuPM/LFI0GPjmcFOC6xYcNUmsMXNCP17l5csmkTzm8WK07VzvgiHvgPxO6nZC
zBBK097AQDyglCEDy1W64dVa3/AEPrg2JCXb4DdhniyeoIPMakQDxUHGdgrZvnXs
3Sbwv1w3xGNWIZjkcFU0Bnw6W04LZdbbo0Ccr/VrzF2+15aShv9uVarLbnCDHx91
7AwV8ne/KU2FcHAEChwCzUGc6ZJkHQZnBLaa6F+OVWmjGo5IrxwUSUNJbCg/+iLZ
Kw33l2Uh0pS/tXGsUQk10QQfVtwalgGKbgiUtfJrt29nfM6Pq7XCnbp8e5CM4byX
gpIaUAQT87k/7fexOrx1OBkATCHz43nBV33zNw97Cl73M64DdnjUCa0/Egd7O2+K
h8RRlHfSfl/nCZ6tQ6kgqiuMGXcNYgCozki3wmBvRpWyKiv5hHeJIp8tmW7UhkQ1
rDsGDLoyF8vU4b0ebGsbKS2uf2HI4deSADifkGaxwIkBgsAoD0jrSm8YIaKvvhco
LHuf3KLfqmsVOwQS7o/fF47vYXnOn7O2Afz4l6qPsr4is2Jgjh698Ik2DeE0BCgv
T/MkYRBprSg2mfz7r6j2yCIjgVtK+n729QtXhpfYebTGLzlHOMI6sbxkvM1xawOl
DvoXeV3a7569LZ6AI5o0SDPlFsnVVGpqmwvFnlUJ6jspMD/rdnjypGxqa4KWNXqf
rYjH2khDhavCySX/6UBsjpfEUjm3zeZ8G4pXCmschchFRJ0oDzjn0Jtdp01wAcRE
mSDb9e+epV7I+Ut4nyysobYU4cSxuHB783id6go6BDyrdW4ZXduzsxhP30JGRV6p
QpUcm6hX/nbMEexCACTSQbZrTH2E3ArTcmeDlzLdn++QkoiMysGimfI0ro0DX4ac
7VkNxjrokuJGD7RFa6s9LkpSxfPxKIKjpxMZDvn4rbSBG6CxgFZRb6GAQv14M/IN
+3RYWfFaFKCocrgc6TMaZ3dHq8UHmGDm91/8D5RlJrJPqCNqw9O5bOmF+wEbyPQw
5VeuTNawpMugtU1Wc0N9wJIqaDteZZW2keDE5KZVWF0zJDISBOL216lErRuy47Nn
UdZ/tERQzh43MB5yw9S351xmbQwPYgsMQLFh4ofLodV3/jieR89MsVao8t8205lZ
GIUjl/myq7IhQnwW5LRG3zbrclwlOKGfnZYybfgKzkCtXyXFql2LwSimtIOHRuak
Oeymigy+oluwVGlXgPdUuUW3kqon3kzPAuyk9XdnawOOsGgHnX95+QrCyNSPlPyX
OSLGbuvJkgDs9ozq72NWxhpmotBiMNGweOqe2iMvGAXQmDKI7I1fAwclAbKlLBQu
4L5tjUWEM+WO6kh4fnFI0IpblzugsiMcnFcpxY0kbECqLEx9dYmoj7eblMwwTMZm
PzNKHt47MTNfRfDuBZDsqCMbbnHNkSynpCnMqF9cMTZn8GaXYj/F08N1BsLNp/lL
OBDaR9FunDbWT+3QW4bvMh1UopXGAiBHAl9rMlrGhpR6gVuk4uKd4OUNl1mhGNqu
3p4yoFJHZAdLrSQJpiahj0mmmsXHRg1ZvcXltctot2w1mFrYB3Bqr8c04OrGZnVt
JSYGvETWlMyc6RXkt55a+uu65CuYIjY2kdOWgquYEYsVtnNObyxmSwqsqqhmv5bJ
29H6807Q8gkeijnqT76sCuzGi6Y/iWm646MHa5ceWtY=
`pragma protect end_protected
