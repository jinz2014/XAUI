// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hbxOAen/HkseYrPOqlVdXZtaD6rX+0PMEMblcNMehOc1m1asKRg/NhxsVJQ3to3O
pOlPu6wsjrCO+Vn4pgyhZ2ALvbMRH8/MQ76znkiUDiGJ8i9nAV+y4XG7FtTV9/fw
tWWG21NeSQHFI36zQsc1KixjKU5N0h/ujvCdgmzbe2w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17632)
ZAWJGg2ylJqxu+ENd9Pe1T285VuHfczGCHN4OhX9+nhnCRpmIyGBGb+/i1ty5zMt
S7QJu/Xgnqp4bX0z5CvI9+ZuN1a/osSj1Xl0PckyXXxnzV+de5Fs5l7/myfHWEfL
V1dOzh2qevKCNrI7AJBj63MWrSkCuXwkJbG9VG8o5rW2uabmBM/gseg4/zlys9D1
SUKueYTMPrC48K4z/s0zylfGKhCnmJ2azn7EYz/qKGb81GfmDGZpJeHwOyjYskw1
WbsGBP8+kXcLPB4Tsw8FE8MB+yXShnP4uPqbUfAWp35+MuUvBzqrSRSD/X3VSS7D
N+X0bbHpl3+uOKGUTawxSQNX9xx9nPsBgXajPu8MSUCmNg+K3CB+o4UCcTfxamVo
UJM0dfwY1feORoPn9Kjaa7uLquIN89vvHub5pZYMRm761fti6A6h7nQWtnYfyijg
Z5SKgqGZjFIe3QeZAWpSkgqwLaQ2AkhJHZoFkGMxoY+c9BTw3poK/Frz/pdLP3uf
1Q4UOBd5clxWRUBRTXiONPlIrQL8ZdiANJTMS29Go8sTqHW48lDpKwW/iplgio16
hpS6vqL9NVkxrnK0QWPPaxHedcxaBuYcxzbkrpnJdqF5JYGvbnVG84weUV3Fich5
8WBPn/mODj9MSeqECwMJeTDfsfR/JWn35uyXw7vXbTVk3d/WoxGxXFco7eZ0Nvw4
HDXmkPehEjaZlg4dUms1zrRzoDLeAbALDLlNTI9ssEkUUTxnzn/dzEYbcddSqHW+
AIYGWL50FGP5hJ4R+/J55vGKzO/Ex918x6gb1Wz1Ag9bnkgSn4zouulydV9EUkmJ
KZRLBsyarV/u1+l0bkr6nAugnrf6w6lxQe+ICfGM8RLH1RAIqWZRVLvoNfxVr9nX
Z83Tf4u4WoyEgg7bIu0TfIGYvcy1UNR4AMZyt+DK+UEIrGI7tqUennnN6Tqcy2kg
QnX11z+9AN/s78rGZrE9ae2DyMlhn+WfTLQa0X+UE0Y0GgbktUEhlYTl7dbeOUim
RUh7clV2pDIyhiZ/OwVnO9lLXkN31bforKTES9Banu7tdMNsVX5dql8/TGY3DZv8
wkHubyhagg46Ujz4mKXutz1JmBUTG2lSKy0Bh7NCjrWRgP8qXKggMHxeldc62jC5
ZX47wISsUZlwH9A9WZ8VwsQtgvrowqb31aIXhCecgDhmJiHwRcKgq1633sZwfg6W
mik1ZYuFgfTESISKszkmQJfU6LOumI1mb/njzx/ky0QL7VYs3xZY3+rNqb4i8EJr
7xWXrroh1v6XRuJnNiKu9Vdv4BRqSGGxtDhnO6mrKHuZtbdMnhufarjVOy8YO4V6
uF0uaNU+sFdjeP+nYy4IyswpMZP+RylRoun7sL17oq3SxqrBtH2TYnbGkjxNbN7E
n/QoQvqncRS6AeAFr8GSCOuIicYGYGEREZ0gB+Ga/i+hJg6AlvGGTfqrhc1TaeWD
QZouKcnrA5qEGaYfsd5faiU+bgMCnnPiXevAHlQANHoP/WAFPUy0kqWpMxO8JaoQ
VhO2Y4IXrnh0iFQtJ4QLMRPjrOYvrvSYLAu3rVGSKNat4eueYoPQ8D/NzwZlvyOX
IYFVzlxutXTPZjnPWdrxSaKyerlMeOZs9+Yqxz5BKYlfT/rn9qE5y3euSxBCB8zG
KZ5jtkM+FGLSNi9l+br14cQoECveVZ27EBRbjaGy/rh5Go3ZAxQuDRP9aEc9/PWs
amQAG+6KRkA1uemYFNUVJaavUYrgR0ee9wntJdCyesOmfQRIqXfntjbzUFCB+Z3H
NIqJfyb/Z1uQhnkH4SXznW1ZacvLlfOGocubw/qdOM8iBvxEhSai/nJTwZFgJDVR
Eu9Inn42syf1xXHWWeLRJL3N76y39jH8WrbYpLS1xX30ypa7GaA5CFc/JfN+txyl
q64vJBeV+hGxvZgDA25WN10bybyG/TDjPS7T7kX8oL/2RhTeUHDmQcnUGOhm8pYL
6qbyudGx8naKSeOOGJmFZ0CdrZ9kGmcxO8aV7z2JQC7cZpv5krfGjBvCpxhN0oyF
8wEiYCWlnliT1y2ijpo0f9LZeDDvQr5dqOj6l/Mq/CUxG6jURymAQXW3KcdRKnl+
ktPL3YOkTN4/xQ+TdokVlk3pOV8WHuVPNNX39lBHJyEn+AJGOh36EnuQjz1q+ogi
18BxRpukvA5wLupyoHJzUh7oG/1QNJRj7MspMZci/vTMWjq4kPo5Nn95nD4mcIEq
v4Ne0F/pOQ5e6PiHFMkXZ5UkHERrGzlB07mhuKSmC5cwg8SbZSxzG5rBO/LlLHve
ZN/rDcgqE5HjuwcV/IjMeTEbsFxqDXZ/If+pzluw3BNqbaL/P0AbpUBztRFfGaMb
YLPervxRmzr6SB7Qn6SYolYsC2eZnsRAjnWrhXHH27tT+dPfYZIVYWZpQIoVcNnJ
hKFqCgnyZsYMwyuj8C8DD1J1XXyOROuT4WFZesnOWeVmdYexQkFtgqckuzgcXQwF
1IbKqi4wMX0U1KMz6bFUYWqRXnYeVdVgWG07eWgDyKX8XBg6CTG+qwOgENZkYtRB
nIzHQ1geH8+YSiObF4SDqddeSgF7d7L0Gll5Hz8yV8FgptAPWnOqE0lq64d3dwou
pK5Jx4LEukR8/OvLg+RJbXmBbqwS/U2b5xhnF6U0i+cWg7PUs6inKC8yT+140dpb
//3EFYtHPBXYaYvoST0i5I69B7QTcYkLlyJL1FRNY8nTpAGhheHicpJ6ytPO9jF6
/+vAyehhQZF5ZDuFEkDoZLvwHEEOmFUkIy1Bx6YjqnWML1WH+SYfdg47M5ofmcfq
b41VXVN/0LypQ3dMy+Kdm4UfmNp3Nq2G00m0hjPsZhfszCnew/AnxguVa3KSQ7M+
clMCLBKtGjGRXOpu9YeyACyRCFohRUduTvTo+VGnbdj3+2agfr8f07X6dg4pLBDQ
bPTbLIKp8XyikhfpcAfvzOgaIH0VQjWWl2jSlrXDse4qHFzYW4j6iPWSA+kNbwm3
ITA8QXXejpROPdE48eDWfjUn6aFeVhUM5b100T6ZD4dtFht1j1Q/YhUivK3Y6bv/
0kLgJl1Zon9TxJbK/cqoTNfgWe0yHPlch3tgEuAGLMrFSuQDdt/xDakJHSOkTbTv
d5mXHMQ3/x5KTL/uoPHBUfERTXyfSiC7/ApDMbgc9ahnG8kyI9xtzo2gog+4jg+0
6m4NJt2tEvABH0ZM27SggpidzeHWqQILtl5zzAMOYT+p8OmqWBuwSyMTxgnWX3wr
EaUGFz3cpKcHJqCyVr5PRSxsLGYYANvbyjMmE4hapEx+4spY/uR7fYDJTUaZyDUw
3ql10GoSjTrRBeSiMWfvv1wT1Z3lkP4QwW6xHdJBwLwHWRqmzAWXlW0P1BzGJBw2
8n8xG29fht3YM7ovuc4s5WJl9+NN4Y4E4+9l/C8SIysn0DSfjHzjx10GH8pnSZCR
htBk5gZ43cwSzrxjJeGrleF7PZuVZb9NRxcm7pldIw/966Iihu614WDbpRWDYCmr
cNnmuegJh2QUtpX66TDxS1eVp5nKV3FbqBV5+y10U5bH0pd1dO0RdJHigWRexbZJ
I0T8XgmOO0awiabVC5l7Ntl24BZvRJTS6TcpywI2K6cTpIwNipF2V4Zt0jno4p6V
+tMSLuCLUhH9i0Q4Cuhru5MpG2GP2refZ8b+IIdvLyecI68g3sodEPrh4ZJ0PeMa
9Zea0NRU/aKwIMu6Ih7ljqVsvaKm51856mzARntyZkKK1aXRpri8LYOcqdB3Cxoy
dHuJGoP/fpuU73elfzbgm/22y3yG69oe4gB9uieLZbw7nLLmlFWamgCdYsDn8rUc
Piv3nwwb5JyfUG+yzH/zy8xU8ct/Zc6iBnwM/stLqLeAIGy1rIFIM9TA2W3EoXRJ
C4PCC690D8kZvW6LMD8TxfYT2DYB1nQPVtBz2qxON1e5j3I6n6hYQu8rBLreR0Jw
OA9FNo77ond8nHIo79ifET+EhtH1m2XqluvfxpU+ZvFidi3OLgiafFb5pQ2RRqn4
LbvuBvIa3N8DhdkkDmwuSEr0oeuDsjHgoSqK8tYfm0B3k4gVpPrQ9RW/U/zShxtI
gMt/L63qKiDoDLqG8dltmHiExIvlJedM22kPMhYlGxmG36cN9hx0BrIw1D5FcoGj
++RhUeykM0rms+2impv6oYSAtlWtryh8u0cBGzgnuAaTLuh4g7C7Q7B5s9MDcrKh
P5MhgQOA/I5Iq7iNr+RFUpaR6DMbiZTBy5elIgT/dLnVSoicsTKmmEjvLquyOsVE
HYHPNT3ZswztJEdcVemJUITL5hO7kG8RKK7fh0LbkjpHrTXHfz2+ipWz+A9HAGKJ
Q9csuyB3M6I5l29W/IVST4V/SF9Ne0O7G8TbOioGpRY35+urR4U65WSuONBOV8iC
PooXjGGudbukOPqFD5LndbzRifgDu1vwPxe/znK38jemiZuuUgBMnpLCyaFBWGBa
VUpFn9gZyfH15LORmhLa3rl7p8CkTmfC2pkONJndtDqVs5hrwgXRknSE51iXrzNt
7Kn6E5gmkoj/jTYzOnU26QtNCKEbWLggh4CRNNkTfQmpMPTbRKjt0f/lJ+hpbUu/
tVBDf6SAwbStfuwxVddgi+IC8ESGdB4zF7VXdpNjMqq1v7nLLjmuPMwkpMr6Pvzl
tDoAgcw27HivEZ/+KlExnrYki1AQsyy43tLu1uOcVBYeSqGz7ZEpeSj8pGhPPF45
nydzX5nn68k6RTCVwuht09cSf9PVVUMhgE8g6drLCxOZChhDEOzZ8ywRHxxy8I0m
ZEF9MsuDmDoXQGW0BcAzvANtazuAudS0qMCZjOQ5Mm6S0gAD+vFokviJ7J3+qA6p
9puolP3vDpdif+lJLACzNTDR5xGUxAG+akhmmEC+LCdWcZzdE9nd0ADtNItwjMfn
G/FuSxUtv6nuWXnU+GPPt5oyBHTRgJ+X08tWPT5dYbOAnvd9zJeQ44cgJXf05Y3i
eExdSf1cFOt+mPSWlUuozXBUU38dVYb8TJc7X5o+Jmx/nQY1bkS4ONtNndxNNWK0
GeNaX0r2sfThRoiKb13Xbu5yhu1w8CeaGGFk1zxCKX1WCtJ2xHO4Z5+RhqqxmZXf
sbSj9TZ9Ga8tDsm4UwsLJJoGv64Q62iKm/0bsoL/Q/qZOCL6a2hp8pCBufOgredh
izwks+3Jc8Y1A03vgh0GCaNG9mA0jFdbrsQBBuNZnqKIURi/BAqQ9VTM1NeKtRY6
Z1YS/gyrb6cDzQVFe76IqtVbwjPnbv7YlB3QLkzGCSZi3CHRhhKgXIvy7ZNNYHYZ
6kNhh9OBr3BSXljxNpswax2h93ZiBONkwVyKcmUZU9jensguvxPvxJsY9cmi7myo
otWgoEHGsL9fxGbSfCyH63o4ow9osK6a51hlanPIeisNzhz0uENG2v1v5QNt9y9e
SgkqrXIHs1gUSn/pdVJjMJKz47A8XWMJaKqn7eNQoLA1cD+5rsnpZk2dtmO3d5Pd
ZV0p0/IL4Nkh53IIUOnVeE5XiTsIoG8U0J/KNzkU9PMb6N1Fn/5D6UkBowTw3DpD
2gs0OB2AQmyqjVT6YjOkKtVfGEvtcw3fwvcrzAeIRVbrg81Cwxvl2sMibVB+Nnt0
WILbi7RPEXkKsmY8OenwpzeWKC4TGbnMcCOfvbyEtap9z9r7vrxZM+xDKxKC58yN
Qzbe08KxidfMjhwl/5AdjQKgJLcHTR45xq3D/dzI1Et19KXPxSo6zpH9iiTCCfjn
MPG7+WVPMZJD5Z06vU4YgF/L71vgP04tiNIQVPl0nzorsDi8vxcRRmXkztulx19v
TgEWvmEetOBvsDAHiOa2G/HD4viYnOfsmphOCZTFS/QRQJ2Q63/QVNzP7jYii2EJ
EDKHxZvxSOGzG7SfkheZk0vjzUadCUtPJr/G3rehVPXw4nVY/OssodtqXfHe0OF4
omjUV98U5rCeyHYLdJS5opfTfhuigJ5nCx3Spy8qLAvhP7HO699XtDdHAPeqekhb
zwZ3lhRg+KeUgIqViZOVwZcVk8OpMdnNCeP/PtSnJfdOJXIUVNipOuzDukXFhCN+
Udm9WO5Lt8ky7M0fyOu3DHQ+1uEKqLbJfHnDjKqqCoDi2X3opXPFTH04KcjDf/I/
YDMoof3zge7YrIVy0ochZgObATvP8zgOIwxcE21ahuFoFGdaGm2ncNifdLRjawrZ
6NzhSsuXDDrYvRsAPWNWvwfQ3bnlCageuzMej68P+EJh0wa2K8cA3LKzfoIsgh8T
CwIDFY6zd/3IZMnwy9328avhpkDWHQFloSTLmzJSgoXTnh07UuTB3qEg+jpvx+GY
LsRG4FezeTdamaOPXnCck1Cn4adeyRBMxnNS2BEOvP42kW3ieIS3G8oSRURsF+1P
G2yJ3oLdtCvPuS0o8jk/aNxgCEUCS8L8y21BExC26Yi3Crwl6U+2gIcSaz9yM+GV
windC+R6Vy8LyB1QW90YYIG7NfFL1j48r1wROaCNU09RBEIJl0jL88wv83sqr53H
cvs4Zbflje+nKPTOFqJTebi0zVluW7YQKFsWIrxke4gv3y8+fWuUPNdUC0K22aU/
PJ16EyUJOWk5JUc7VrKh5EEh68c4/Tb5who6eJrXIDEkl6hB8xP54/xQdMCRBvN8
NZsj5+ZVtnUsSyvd0frpxh4bP23SapI3YSsEfFsocIhiRYqtSD259oObn4JYnN1q
yQY1V8WnrFCXYVdqbJRHGlPBtm2RndTPeuNXCbwNUZ611Wlo8PFGnbRo6teGAg5z
iEKLpKQZa5+Kg1pW2I57d6HswmQf2XMdMlZ4ariiPaN0WtLbd/t/ET0O1ZmM13JP
S19612q1UusbEysr6arEykYO3poA2Wa2WiUhdGxzETDJdAZFA+fne4+RrnfgxwHB
f1JvZKjJFDza3hdn1lvWfq3RShdKm0seGOA5vEbxK8oVQfBY5ZH1FhK7x8pOLKnJ
iSYu7DRtfbqOVAjX3zk3x7YXb0NGNAYW5uB6MwylzyjgaIPDgnRpHi3Z8HphU25o
GrigG1UjQE/G9+DGIJZDmPY0e5qX+t3DGeSQ+3QR3HLGz+A5j6my4hxBn6fp+dw7
1rltVC+4LFeSLuuFg806e+wcPSbu8+kmYZewwJttbxxutCpHG9ES9V7Sww8WVLok
hE5sLtkCKfi1CoVEeCaC+5/+VtSaN6I1AZEQP2yGOnavankCfbKt+cgxMVqImycT
+6sGbccwtOfRt6jFS+65LEbO5ZDRSQgHh30UM1S0x9FydBiHn/jPzDKpQ31Ex0O+
2kUx7JhK1XZ+JijXI9jPR8WY+Xeto94JznSNTvIaoKqbrgQBAgMBXMx26VkGQL45
7TkyO4mxuO4miVY8H9orsNXPgbr0chE0H6ZV04suDJVtWKEml1Xkk4AdiO7g4/JZ
Wh0kuQ+66HxNf4KvASl5dQf6KeBlfH5PR4zpEcLgvn9akkMEO9bRQgRqr5CYAEmo
gts62JUzkFS+QGw0o9UFw4Ds572I4Yl4xgOboje/IUO+sQFcW3LHRcQaWzfC9lfI
WIFhfA0EAdNq+qejuWoxBzbeQymCR0O7B/MeN+y+dB5YhzZ7PlBBH09mRpXRw/fJ
myp7n63rq5UOr2tLeJPtmPAJD1qyrVVRSUjZu1WyviiM/gSzSMSiLVhqe+z14zCn
2T4kZUYVDG0D/FoEywTW6s0ZUFIygU1ugFbmmIJcn4qoCeAKsEV2UfdVumyyhxRE
2v/yvGZn/sq0EDsk3gmVji9aUCE7dPhPJiGInb4uHsIWSfg52ykdtvEVnUCjsGMS
fKYLc0tdgOOQ5Sjq4KffCzQf7Skh0u2DC3aMaevyFnsZ5jIjFr2kygQdg0A/uN+m
MKpJ40FVj9AnoITBRSKjh0tuX643bsbFFK/X6lJgu/foWMPCKDGAfu4E1hsYxiKO
biUfzEnP/Ea14z2cNwVims5GgI00yiHz9qvjrUX3qiug6gipBbmNr399PAlBLLdG
+Q0JaCOOrarRcnfwFSFQjGVHiscAz7PA14Oki8dTeVVHYMJhFIHu4aGel4lh+oH1
4F1Q//l4PX2f7rtF6RkE81yEaCb6g5MYzlRCIvLwo0ggZohFZEHu8vUStveDdqQe
0j2FZcDN0sFGnvMkWWbYsJ7wKuslkzYD6ybIyq+JMvoHGGqyBVVW0ghhsIXLnguB
cafNShJY1pKD/5h2q1S1QB5BWSnl3neZPezIoifvW9qmaDFfgFJ6WfjkRdBPhQjI
5iSGdg7xuXJXn27lsRuITI1BL2/55tOjbw1DH5286/3cSUDeM2AfH0gGbPfuC46m
T69Md2mKN5P/jHTt3oc25Bh5Y9gcZ4sKq+Lb+nxH83JK+ZKRw5Gukh4W18ImQ6SS
hqlewFCeahi1ksdn1GG3bz4ibbSaNDRsPVfgUerXa8/d5iVjMMMbFs8XxBzyB4HD
dwd8rJksCCDW1BpJV4HV/w/QGHmkvJRhIRROL6AoJd1Sm0SteZCqt4b/uatDQDgD
yoLsKu9uAg+460PeSLMkRhGTAncFM2z1B5fAsiDMbzZjkAwUtC1dzBOI5teYdzKj
e2EOzW/xiyjpvOewwog7vwAPSUtaq6wUv0EOG7g2eUbkej6urzwCNXruA76YFMQ4
HVFOkphdYyn+QyRuOpJNsq0ECELdPk029IZp4pAroPGLEevuwTvWx2lfbKfx5ovP
ZZhCkw4YZckXldW7gPvmwsUM9v8oL4VwaGXG7WHBvPGBj3yy/MQDElijec4edeNr
OkxtSy1wo4x2fi8djxQs+CwlFeQGWCavcQNjZKJMjoVIAvnbr2WWX5z5IrwQ6CUZ
rDiqqaGUmMOrpwug9nhnc+vnirERGcv/5CgQNXqegg3U6W1iWl5OYLdwl8u37Np6
FWMOM9UetxoYOvfo5b0GdL6pEfte+pZ93lu145cUgdWTK+ic7sNfCKoDWZecyRU6
mtAPUw431mNGQYHgJoFFJVlONNGDHgK6tuGzcmSFkw4iqSicsQg/97sKA0pHE442
n4GbSPaA0P5qLH9z2N97U+ounnXYQXKNP28E8RJXKHQeYXOWZfkpzynKFD/lC7yk
Xgs5UM9gCelZPt6+L+KJk+sjqyIVrW1HE1trWYyJUmQsb9SOx+iZ2KEdPeSNO93B
5QkiZwhvDUjPtYjrP9VDALsTf0OEEf882ujGo1SO5qvPqUjneMCycgV2wwJPDo+T
UBZNWmUDJplOvM3NOB9nUl2JqkkKsh8JpcBaUSb/FRbASgP84Z6aDOj3Etcb0Fd9
SHMXlzHM2tsQ7YgGnd3Idl9uPkQetKvUebJWhpvzS1vMzMJJZ2Cj8PAdnM7o7U6e
o0P1NJJE43eOyAaJ727lzAn3jP/xGxBBFEbCDrYrH8gajBkwgr6Xd7Ojz+6Yvko8
kBXVF2gYFSskNV3Y7uwgo8FrOKkmp11ZXhQs+5oYfVNoV4O9a69hreQ8ObdF00+X
olVmzMft6xPTKEFs45pPYUBbGgfOIOp9tnk5Uat2hYJ1Dy8fK9gw3Ex3ACYe+Qyp
hTgikfnhUeD2ktKiGZ6n54jfEN3+ijyJni6Cbzrfmhr61EMXxqjzOqv4XSN2kc+d
1sT6Ul6iRfkoVyFAKNybf7XOiiQJxfk/suz+OswJ3keBZDjq9jUfug1kp7rVU2pq
kVIHBr0dWwhhwLO8VE029rNK+i7G2GSonDonDte5/HESUpBnvM+Ror7Ufe2Dlan5
2+2bu7lFRWvIUTV0oODQsfVTqI/oWhjL/DoAYaZACNiX1mEVWIRegpW6tjur/ibJ
GOceHk3SaHqW8We5X+k+3ABE4mYswCLrCQsJvpT3pSxcS8Uyg7HpZJ/rey5dsc5I
Epz4CpoSSDVD1jZVZUSvNrx07/NueJMlZQqUyI8MLwom+k+7CAB6sUVTgYYOyYqN
Kj8QjVSsll3FcUMe4O6xm1F48gy/cc8b+TOVSPiIfnChJ1YOFTMeN9QaC9JBGE5i
mawo4IYKJP/KuaGI/rc45Ytlxypae8kD3Ukk9LNcHnrycZLskoDCMakC7cvdYvvJ
f1f99DnntODt12L5j8j+iKiYSNOfS2w1/yuoCuQLdpZ90b90kEdLsw3cP5zLMEvD
bZGEMBRspL5lRSwMfiAyij4Uo897kBgvrfMQs+SNInHeONBVLTc1aL22SLFQ36Rc
N0XaHBnNFrFE1Z0E5DS3lldHZxnDRAaa13mwSuiCrzPWryhvHLK66n649DnvV7Ei
Xu8IIg8kiPuVm7NuChk4MikGby/27NPCWvGUd8qq4r2+dakD3ZkZJ5c9mMUE9OdU
E3pDO3UjVGPU6Ee/o/qUXnElZ5+IIU6mPYxJzV//Vi9+enc50Ya3KpDBlSOdWg8k
FuRRCo8U6bxWbWORW4Ii2m8KA1BUxGMY6uODkUj91PfZ7iVNnmeM+Tw+WA12LgFS
5OCfv0OdMW6MenzG8dR0Gngi85YjmwtcpBHf5FJER5PhzkWvqoiptu/8Y9HC+05O
fp2cVjVcWvha4fBvlQuu13+ZyExDOTcI1NoOGkQDOxEwbkZEi8qn6FJM3Q5V7GVq
KAcDz923r9l0qbOajF1WL7K6Rx4uG8TfbDCPY41hYziqiVQZxWnkdqOgiGasHrfx
XCSa33yIPVFekrK0hMHQtgN/AVZfMTxtoAlUyHfzc35/UdJsVZ+/CbwZQMtWK/aa
TaioSi7xGwUqeZZZ7F1LOheWC0t9yFp8x366ABV6ncQVC65/e3GDxjZGd/YOswWx
kTCjUHxhi+L8qvJdrxKPCMrO/r7D1+dniRJCDEO2ZouzNETRBnhWDWykhGw4mxid
EuXS1CPuC0bA/uo6eQ7ywB7E064JJXxbF4cHy1oNA2XXJr0D5jYA38uJFSnMd92n
HCn5XS3v08S8ueFNxqjK7/HLRCL1pJWLUa4CJWEmDDOCjDyuI/iPZdmFfBaDjyZc
HZySjWYzJeqesUExGdGcae0ogxW2MObe1syam1pQzo5YyG8HQg6TV6lt224Z81DZ
NHljN0mbjsSS//jqevyOA3ErL/Sf7UAGxXjgRU7pQCuD5m90tqm8O+KVHbYEXe9I
6PAcDpp3FAphWOTBQeBdaKOU/asABQaXVPCK3kFNCKw441tNSNSkrkETzkN5fyI4
pvlF9Pu0PuQtZrK2+2LWKXb/e6Ojqv/4QSIjUIN02d5SI/FR8TUE1HnRTw8eNXo+
uR691ILZGSahbi5oOsMzQgxIxwJZcoU6w7iAicW5LiTrFII0aC9r1xE+uDExuLdl
OyamLUk95kdHNp/Y01cmZaiN3L9wFXDvoai7ROWF6xmz7NRlTNO4uqwk/SwDqerU
sr+tmIyshOFHiSNrEPJdIN4xGkeeutdEg7jDxkPpJz1PHAIdeuXIcqhFoMaiCNkr
DECpmzg4yn6hHX7sDbUgxGIO+AyYC082KnsWt+4W6ojq3786tJAVdRF4pR7mfQBi
lHISAa4PSmSinor0CnZjdoT5MJ0c/4Mb+iNQXa/FA9ARFkGUtt9MCaC2AUeCVkh3
aD7jnF88Aueqtzl1r0fhDO6qArxV2wOkBLEBP030nulsa1HZo8H7ARwSAtcey1yS
pLDbwKSQv/Ud2eqB0iAWX95dnM5FyEc6FM4aWMf0y/z5Gic9j8fW6I/VVvCmvbd2
od3IPFY+enx6OFbtZVRDa+BN21MseXwx2Q+wH80mJ3l89xpaVdoSj6Wq9ZE+Xcc1
2sp8QaUiugfUGqTz+s/6xOAY62gBXY1ucBv+XSVmkTI0pWNyhky8i7haQDZTpMF9
5ocNh7Nh38+tyt+2d8ukzIXvwtH9DAsRrUVB7PoeegbA2KP6BJcUvQdE2IGuTa1j
L5N/Wy0DYz2xeZ4SOtlodSxakICqO181ZHUPp5/YmP2/6buo7Jst6ZL23+mek7Lq
WGZxX15t2va6emnBxxvRBruQRe/rpVYSre9aqdN87WYjLlq1z4nIPWODvgjJvIVv
RtiJ+xKkUqFsJyEVxz1WrJD85sqsqbwVc0WygnF3wpjppb6EUMAkpGjnWhManIl7
Xmy7U68MsMkbhj9Htd0OmhvlVJGcWaFPux/MAKuTARlAQpAiFmfFfqnVWkBwXE2C
shUyYoCYUUxFnzXzMwUeTpAgIfR0DzokYFab4vaN0tQuCCsHz8FJd0VbmBzd3l2z
2IPaf9KA1U+K/Q3BCF8MVwZTfrM2SHAobQAVoZ9yGbcPFPqHTju/+cGspBofMRjb
7gGAAUumJzCl1iekjeYYzGs+fmxnXwjJDjk7ezob1ahELr2rwlww7V2EVgq0LZF6
0SpDXPrW3N5SDYvmhLJVW7A9UnuEznu/DVrKrt2X1SszS9PZjvOWnJN3QkZoviSX
vGAwCZ9Q48rDRYPJ+r9A4kNBzulyV2fTXpqWMr7mG8qT8VHqIOxBbpM9KI0JLXnV
k9RJ4wkBD/KugZNca4XibrYZOoW9rtS7fYfbGNqp+IouEsqQYaTEZAuGTPou5jI3
m+QOx96glKO+v2oONytfYWqI0cUUpos6kOk+mSFwSubHDtXwhCjgnEmYA1LX+YLX
k5ENcwvFp0/wYm70wzSdoHU+AzT2PZ/8e7PjfOdeLlfjBVQmuQVmZJS36dc/M7hH
j1PMlIpZKSU9CCx5totcaldE2yRm4SvAc2DdWzuWLGqXf/kg8sz3msLcs6Sj1pL4
xeiqVd6y+ZHHejvT54Hj5OGUrXMb9WJfIILZ3lWMyhvRqY+oj3HwxF0G88hjGWC5
QrCNMI4ozbNtKN6BKaRBlhr3nqaTEBLxRDi6ImYenGHbd25t6mTmfrgUwLp75+/d
k6YOe45LwxwewmeBeMpe9n8axfXXrTcEnGlovsGxxmvsRFU8Uh0XyJIJcnWwOEMp
OQP9HQ/JzN6PXXszloxNIWNRykfcHj4MmPwaP7sm/tWAlFLWhxfza1DwoH+KSwlM
6J1B6ys6FLOcODRlGHl4MZ+46CLXjQBeHmG6JwCgZo345KOqK1B7gGEG0VauP0o9
s5a9M3z9bQNLXVVKVy5TimcKC89xik8jFkakEifAnmU7A4GpwooRIQoIdOdTxieP
bnw4tI2yQrd+2niqOOe0GTBDd8HNfURadTMiVLRljgtYM/9iT3H6XAv5Y6Y1+E3q
u/5tom0IVjYDyEfRiprnQxhZgPZUp1jsKaRrCm1oUKEnnQCvSv/BnksZb8DmbE8o
cMhRJ1buByTKTdzq03HUIQ/wZGeR7xDyll/zt/eZEqjGjnt/BWpU3oOI+Hnk/uwE
M1eWVENVvr8k2jC7+ju4TbotNaE6yLHaqQwSeuZUYz5VnNqodvMi70cukuicewm9
H3cIGXtm276Q23e2UiN5dst46uaBYyRhqEbklvwb9T/iFQPr8PWv0BwiEBtW3MEW
NhyqUE3DtGzOzMS6EpcV9SLgGKAezmHXRUW/UY3LTL8esDzBX8GJFYBi+25eWj+m
wH9K8rNOrs+steY6RXvjGWsOxKpqA4mN8GqF8Lq8Fvgos/O3ToTgGne5HsGNY8b6
gWm2grYCMJ1NBF3EK1h+xEuxDWZHsyu9TUCgxTxWemRprT8bHc8++KwSc5Q33Dm1
EnXbVNj9S+zZovZZuEdS8Vb1IN4uiXkzjC/vK7mnohFoKfVgXNlHZLsTlNV/0HxI
YFuMGITXm1Qq7UKs0G+GtfAm1dnUABUMhghkcjbnNuwammYgSEKbogeS65GaPEc3
6vTc0V4m07AKDOIr7CJ/KiNHmg+P11LoBajbQg7a4pfahCXbibsolXOfaTzsUbWG
R0VhENusI4vmVPY5Hpk8yZEJ9FVCxEmwItFpj97APnef+O7b+2TKTerOgfRdv428
ynDgasTJFY9VP3MtQhDpYA6U+egEhxRnBwGK6nkWcO2JqQMD3b1s1gyRkxDOIRMq
roQvRC4CUClOgx0DXBj+CfQR6Le8ZTrt6Yxf6FeJhwuKsIGZqsMpuzpaBp/PXQqB
mZXaR60VMtp5OtGUyIOahCvPhlV7hw7NL97wIQBl86bjpby7KclzI2VQPwuoqu0u
XXiR5JJko2SCn+Uah+rzVcQzYgjZqa1VTHgWs0mttXmRUkuPhLPGCb/l5uR2qiEz
Wdsw5uee4k/D6iq88E2y4OsYN5stYkGuWnEFNAjyPxgX44eFmpVcuOESICh0Pmxa
R+49onJ308QzL7TfiY7eEPbtOpLvCpkkyEsq5+EN+vXburIFwtfK8z/s18YXv0Cu
7xYURGBT86rHAORsZUmaiCsirqxM0Zd6DOFEbK7RzRkGFlxRxP5RfL4BQI5o3UWr
LILLUB/N9J+xGGetot5G3AFhh/RmMA18pPNUuLf4nMdgVO6Ww3JBowjKNzo6W3jP
7NQnBNTkfRbHaoBwDvHRCyJ+GAWJBXFrFzovReI1DZ1RvkIm3kUnJbCq2nFlZB4n
4yRKs4FRweN2bnm+o6wxRKWr7c45lSgD4zMl2JsYEUQhcltiIoJrWhia9lL9YKgT
COVT0gtw+YSZWiXipp9VZYISoizoCIA88zYaeDcjq64R5phU03NiNdYaIVKNFd8h
yPf7hfhxWvVL8Oy6qC5se5wfjBpvF5glSDhRJFYuNkq9jdntmyjhAagqZ0Qa1KpM
nQpDLg3PPg9hDCbiKzrzw1rPmc5z0bueXgRUoic5Ju1jFcuKRZLY1AW/ETM56xT4
060rXD7akvA42lBGSKe0WuDbd/Mb3klCUVl++YiMqlVC8rSW8Vmb9FLuicuVMcsB
/RAozePdUlx50EkKCHrBcgCmL9S2Nfy1s9LggqCc5byazrOAy0A65qFjZMNeHmBi
jFN0r+Z3VEkINvgY0nJOiWuak2nSvJki/WcxD44aJ9dnjGFUO000femgB6DN+m4s
+Y7emguxYlTTqWynFRklpKjtx/c+O6TbhFWCnf2vvECp145R6CPf1otu1YUcQzb/
Uu5GrtRwaJYwtz3demNvsDs3CtzgAvolV3YmiFyBQaH80z1BH2hjwf9Kj1pmBUUE
Rp3OzEQT+QWWAiK4UMhWTWL54ya4s4XT+LQaL9JujK3zdoPb2IZTRXGDw6w2hv8T
0hHE6/JKYdfPvYp2wCkfII6lLTvSknL8zwEdvECugIK4oeemAk4/Rm+CD6o2A1R5
SfwhMOJ/RUxCj4jVbvJpYeAWO2Ua55lA5WxsITtavUIcbXzVP9ozoeNFajbQb8ur
n/6KJKUtmv7ifi9H1yi+AKCZU4KpC8SmIgc3T5onpN52YLT2cP1AxgMGrt/R6FD6
XrFi+Ozl8l6srVEvbB/mW1krkvWqM6nxsY+glavfbuxA2ViDgObNUwnNsjojrrBb
Ri91/2wAR+e8AIJDnMw7yb5w1F1tWgXHd3wqvPRW2RKN9YSh7eHCDzrJLXmzIK7X
NRd9UcyCup2I3/RTfMDaDyV/GytXcR/mHiXFzRYRu69uYG6DkoXpErB50sdAZzbO
92LgE7Jrf8qFKSUF/UEQkLDeAsL1nF0yw2pwdsuaojUERBG4f8+qgPuJtlTXq9mE
IEyxw8EDYOoWlgmnU+1drclBKbj/oDouuJUZVfzDCN+MvzqQ0Das+MO0C4jbrC+i
Y3o6Wm8i2z7lYl4qu1Lc7i7pRHR/poYgrbHQ3nnCvEaih2vk8HHN8CJyUBys0yK+
StP/jmHTUCW3GH6VdEmlBageNhvmNS5rWdYvvTwiIatPjS5Niss5xwo6GWOPetEi
Hn1/gxlp3G+EO21mQMnVusSEdusoOMUW5yBBebJF6z8GwFx/H8OfaPwXjJ+pwptb
/A1yzoeGKoHrtEH1y9IL9/dXvfC8SqKVMJS5Bj3tR7CHW8z1z4I7K+W6yf/eQhWJ
nfP1Y/CfBZ8jeG43CphM57bIc8XBoMd8YqfCaHu5L4UnFQxrNqc9EzaDtMPWT6LU
6mm12FQEfO9ehB3ss/40b1l8DCBdja2bJmMZGkumO9Rz8xyQFVgPRrhfHwq9JRaf
dFRYh+Z9LA4V6Q7gYRENUijYy57qKAtivHt8v+n4wP2DsPJfNZkfRqT2mZvWPcn6
vzV4m1uXT/E7KsKHdtbe9r7z6njPQR6lmi8e8hkWKbufNzSr2mbgzFKIBTlnioZe
q9Eq8f5a4wWvUF/ATfOmmQfoA+d2lmIYCdLFL9mQHZSPqWSu20MS4tq+8g6oV4dQ
3d8XDJcPyVNAeg4QfOJUZ1UKWc/fLxdfyN2LXCxnmWAWG5iIaPvYjbH+/YmH5ZkX
hFhrDVte6xCz40D0FgP+PFvI3c3ZSg3RJOFSBLU2KVsz7V5+s6GRw3WHFQfmSv4w
ibLfgvZBKK5Lf9Z4f7ROLb4vZ0V3LN12L4TM/tUZm/aZSJB/kA69sjjd3NrdY8s2
avX9JuEqMY1YN49aJ1wfn+J2hr5rMzj5DVbEN/tbXw/ROTqTbNa/ZUbywypxLP1M
cejXdoqmknhhxzGTCDp26dUBUf4UcUd9vnMmOa+E0QeUpVIQyq5yEIwFC6arNcZY
NooqhZn0ne8NMbECLbZk06Tys0cP4oNe8By9/Z88OU+5FfKUHegEoDPQ83c3rVo9
GmNnHQlidJeUUw783pDo/a3zevco9xB/RBTY0bRrXRXyiH01U41hLlg+vW0XmpWc
RPId7KPGllYgMXM+xuIdOmZnpD7I/aj8RMAgo0yS09d+F+0QIAbZgVX4eHi38GTu
Yllu8oPBpysMfH+fVcwWphNbS5PQwJENfrNggO82DVRjOW9PwUfnQ7kpUn2snkwd
fqV56axyBb8yXOInTFpbMmStonUOyqqLMOAuWRnOZZqktkCSHn2wp41ugZYDBTxz
oT7xEJ4CnQXw8qCkoZRK5JfXmH+R4L23EZUa8TOmlRNz01FbYiUVLnnW/VoJIoir
o06KcYVitB/G66RTHV5WEOMbUEjCuqRmizKL+tMSTE+2T31f4/jzRc1ie4zISdAV
1Fd6810BE7EGSYMZngBnDvg4OIW0CZfIzdJhpkk2ekVJd7HeShB4ZyLH8NCHJNHA
uR5VsyMWfK4+c0Cs/CqRVYVpkTMaxYhzQA1sPLWTwkb3Is8+XoEGeKDJTm6m06PP
OfKO6oXfyW1QcSU9SBP+UAwHnBCjCmUETWveMlkC/82QiXlTzuh57YLqZ9k/k0ic
drSlIHayItOGjnbCkfsyyFX9V15R5r7e8t/wCmzGSaX0JcePmrY5AzzyoEBM+s9I
Nrp4qde3D34ynW0zcpJMtUQx5AA+BRS9ynr4iYk/6G4HEgBM63AkLtUNl4NF1o3W
CHqZTiuLDYVRc849oi/3rPDBShov2xzOzUl+/vatH6sentOgnJ6k+Bem4HrgI7VV
Oxe0QggoKmwwfKINI6k63Ljdx34LsYrYDMgrdC2Uw5U+j9G/q91mVhr7ZXjalKjZ
AtJ88mpvXH325U5PVmWP9ZM8bYdKAD2ZiVROqbB3qAF2JpUklZVvE2bIz88s9z0b
mIFIulu2Lz+jNC9QDcIgTfslzbR2O29eJWbaVO1RSfzmI2Arz7XPf+704eZxspHl
SVp+5lKY5uDf0GHsvlWysvcX/4DQ0NMSHCbSdrntpqpKwI1S/gf74yaI3QAzGuCM
teoH9I8Vxp+KIcG4c8HBSKmNz2NTGbdhKrMXYU8LHITmT6OVOaW8HOZqYvIm0EQA
AMIKr+VHUeiSVZ0YoVB/o1ui//FuDWnZXjT1Xp4EdYdNN12s4W3mH47VO4YexQsp
rskfXVF1YROAUi264qE7eWG5YgyY6bTrTGAQzNTw1BZRI1AtP/3IeKQx48dwfJNP
SDl2ATHUfWul5AyO6oTmoyNKGMXvZybfKS+Zmd+4vFifGxTo23h+3FqlDVUcoCPk
2iMbMtzwkCXssCCDmZxnSOnLhBY75fe0CAvlxiK5CdHlm1zyfpiyRHe35JC0kjNT
+Yif2YuOHibXgC4aKK2McuE2KI8FLrifj7asGRtIicuJsgknC0m8a7bbcmF4KM6e
K2NTh+/bjFO1C0ksbNmgjeu8ypbVMJpZqGgC74xR4hbBlGcmyro2gJuvNpoxPIUp
hyRjDEf6u+xwwR6PoIJmWOXiuPAdcbYqFBkefKTda2zszNxHfO7tM8hnxFt3iPZg
5fqXmIqy0B1toEwg/YMsw5Rfm0rhLtfa0VlchziPdCcH2tZCFFcmbMwQsxB4uu0H
zzayTIHbOHQ5meRMMG4gX5BVzmiXoEk2fwjGXbkJRyx9Kp2OJ3SMb6D5haDWLk2L
CM2wZin6NpGHugSMqqxUhwC5FDRELapcvtLEmJjIWYuqLGuYviIhRo3DzA3MCD0C
kQJ0aeAtFNyJpPUguMrDhvK1b4qZ0FBptJ4EalTUSrCFCa1UwGnpOIX3vdtAVCmS
T/OXmrtrX2ifBcrYcvXPybNSlHfS5+bFF0i0ykeLwWPkEz+87EFRAsV+vrm9dVOR
kTEUOgi6UxB74uqlBM40drnPH457B199HZGyyjLWa4CB9/kuxAK9UyycgYBzrmhu
VXwpNXIVdhIKhCu/y+g09KvSPm13lDc3XXRvVlhR2IaKmE+t2PbEyoDfZ78n09pH
cbFyDZokZkm1NgzsBX9hkmvhfjqQU9l2p2kO5y/0aPdbiIP7pzOlT64/ecppbzyT
00IDhuZq7jf1Hj3Og6KdALJUBuaf3nvVCc/6c0oOd/uQwfAYByZG/aru2rVTAL7r
e39CluhF0uHhoizG+UO6pTwAb5YZ3qcNmEot5NF+9agNDq+1Q3lAo/mfzkkFizyl
cLwYwG2nKkrCn0CnkQubu7PdbTgiOxaw6Fxe6fnhven+eY9Sc25NIFuj3oJNE6p/
mq+8RN0O+mhJ4OS2SJq8oUj1xyfeZ+tI+/dF/cY77UKpWD4Jo48Z/tDWehWUQNl4
NVinODjtxqU700n4ngkAx79ZvXgQlzEqBZy52lYDz0K6J+AnRN4NFgqSP9m53GE3
fKv2clUT1F1+UEuCNV6I8LAhs5aJMtSE8SLAgvj0ACtUlrHj17iW+RW6llQe45Wb
HBFbGRn7HBgRD5AP5bsuHWzRCalsQ6hY++STw7XTfkbKDTFQquTGcx8cyMG+VSBA
n7zrNqAsdX3tYv0eu2CM/RDd/zpmGmEvghyWUi7x03Wy5pT/nQkAF/N59Ke7LisV
dbWybOUNO7ZXLf6b5PBam3YY/pD9ojVLrWwtoZ7c+FsD7KKCqwlWLdKR0M4wACQy
PvgaP+bQIgKhrG34fx9lio/arFd1PbQphoyWD0bGVxG4yCHnqzsgtoQy1TdCPIoK
gywkPzqmuw2NlJOL6nNxeDG4amt3+rB5g2cxKON9DZWb9z4st0f8xTmgQ7QwdjSM
NN7n9/g485GskxDOSepuwdWtRZNTGYk/eV7vqGDSbbNsFk0tI899pO4lJIlKE1aH
SM/KvmBYOqnNZK+gskcEVVbnpaz0iiWMaz/MH6GECvF5LQauDIuvTVbv7qqNgMNL
4oUJUJZFPbupObCsDfKjEIipy5yS3SiM3Trc83xI6SUZwrqUwdkKMNtThwFqmd8o
O7i2mx87gxNxNbB8O/T+Wd+jZrT4if/JBe0djChGXL66a03mnn59xaaP5iDuFyrp
/lnJae57I56Stf6ynj3NroEkiq2K8m/UAkhn9s2vGDTR+B3QE2kgOUfStuUTa24M
pmuP3dVY4GZs4qwPAvV5ADGggtPoqx1wRXK1x+ahlo+rfR+kjNBwPyWPZ8+W3os+
hCeWGlYckiITaemBh4geJ5bF3miDQIRm7gKqHzSLwQaSUKjG5xEzXkgkrFR27OPl
gYh3IbhjZlFJUVvHzQHhyL2QnjVpSLntQiKaeEunJP04haHPuQsyGYDCYywp88/+
bGMdlk4gruHY189gesvWcWbt2xBSts6UQ6AwYvciqZbS6L9jN1jQgrzwwendIQuO
eN8TFX7nho7CVHnSLId9wJaAgc/YTun/09GR0PYFEc+8gYtJvi+89ewOE1nR1dHA
0Z4N1BhUqBIbkkUU0PZ9hsSLrjAP8GjbIX6ehLDnrRRXzrQNX8x3zdGFBudSRPsi
SSUBS8OtV2JdfS3U/yiv2Sgosz8Ym26C9U1N29X405R6foH/M2HhE35m+CJOwQx8
3yfm5dUO6GVThvwJelGWT3YBHt0pvK04hOVH/MkuZJq/7cuZe+ZQ8DAgh4mMxFYn
4IovNWqd7SWi68JylrAmZMlDFBAWp7B7oyJvFNWp/yunSlFFTrFAllyYwuHiy+Ko
fY++f4cHyfnh4iC6e4K8F70Ryc0qRc3/W+TEl8VcyG4cRhkCGIKopbn60ITXq1s2
K7TMVbqwtinX92wGeZvRBI+/KpKNN/L7j+JddutU5cvUuXKhcat4ZYaoqLV5UlXE
SZTEcff+0D7TwO8qccv2zemI1m33omxGobp8gY3UQHWEWwHJmUV9cZHfPxRC/EZd
55/eK+8Gl0tBvClyXX8INjJewCps++Vp181wxmE55AP+WJ2n5qAtb3tp1UodUfc6
I8npF6vBe6RCu4VaiYTfdukJJyBim8NEnhgVr/o/WVXaPF5TBJb7Nd4xBv2hOZ2m
RhvdeFzn8lyK7HxHdqJkmGHF/T9x9esOZNeI1kyeMFdkiV8+jQ0beU/jaDqvU9Ki
DHl2xAMxzv0vvdujV3puzh+F6WlZkjRlmCyj4g3zjUqaPZHjp8oZ55iqCaYaIyEp
acvmxsarxXojmBJQKCLYLk44nBQj7xU1IdEBrNl+VXoB1WdmkwUtO79kGUmRXo03
AbuI58AVgFUk9Wzwx29L3hbuG/dNVyHFhOL6PxoQG4BvGznfEiIJRiYkPCfNai5E
gDQPvZs0pLXHGbTWL8D8FL15lWI1tRUormhwWfWH244MxYgOGU+uzDmamCiKFAqU
PPlIfExBxYosLd5Y/x5RlgO6gWgszNIqdPvHLO+aPi11xnhSzz6SLW071KF8yI/B
83qSPfi4bIc67PWfDTnss6m+D7vAe9RtrGU4tb7qbSmwCAYDbhOmeqUzxDdJXGCb
IgXI1M2BOr8vLW1NS/CUntB7xuarosu9MxqQkaA8vGzMm/q/4g6d224bQAuSp0o9
V0ajqGqn+FGiyNOD/K91I7zZ9GAq/Zj6DoUA08r3oxqsJW+75x3c5klG8IjFZcLP
DpC2EcrOoW34xwRz/G8M7ESsOV0NKNZC81fS5iFQrTkoimbXYVQRjCwXSvL4WZPI
rezZmCJBfglMK9o9i+ElSRQZ7riYW09ZILgW77o9XUmFA5qmNS4dcsFG67obwXom
IzYNaESXmBVBa2/8Jqf33FASlkzKCH0unx8cmF4rMUxW/eio0rcGQ77/cxWUhy7I
PRwkZO+s0/yAeqqFgbJiyvzqC26ogaCyDUuwBcyuXPdvJaLELenrJA4rf6c+4r7y
0POEquVzMCw0nMrxPDCDKZv2cZZrK6SDT8ndv7otYC25FXMgc1aLKhooxfivKNda
MXD2DrCeN4bRMFE0ZwcRQdvL7d8e1q9jjmiqoa7COVUxKZSA57KTxTWrQfG5L7lq
U/KSApW8b9e+sxE3g6QMJkMty5APQ/ovCJb8W0srob4z2LdT5VCbGWB50bItFiWY
TJcs/1SwoMwvKZFF7iKKfVbGvNTw4lVejqJcEeMi0rYqICLzKpkPby/pxvikFiwZ
wzY0t8OnXGtEPFdymFK9yaDoulB4SSFSOU/dlLIxE/512FMsbGg1B4Ixkp/NeYri
jruO1F605OlFMJDwi2JnpvFn9aqwrwUFHWCcn4ioy1h1iU3q7mlJkLkBcYKHxxH1
1qgIGc60A10GzIdYJ6OVbIJtS1VvqpiSGQFaEWqQnL8VokSjdW0wU62Xv2VcpHhA
uwWR2IjXIgGnAqaXjeeAxXTtp69HAiPDT4kKfP7xvqTl2F4qvoBWvx8KcZoveSdr
4PmjDq9opFlBPJlOGxFvihrAHIaP6SgYB4gksV94dkSuZRxxCNi8qSN5YW0Xp2zs
Cy3AmdawZjIazA56xhHL1isY0+FmhM0M1IjN9qt9Zq9gtYNQXDixt4CLqEH+18JR
it/Ql71YmJ9JMr2gNTm/aXCWj3lgUoTLGi8Wm50QFwbkhmY4Ae+VlNij7f4YJMxO
1PfBMV4HiWajRNm4w0pGj0k83sLW08F/6bikl6bpkTNg/2TzfVU2nU4zMYUOW3jJ
NEF7ciFKQ1QT+FKTVjC4HQJS4bovJjODDGh/0yviumZhQNtGN4ujT4Mk23UZZRJd
m29rwN87nvk4rLER3TjY/NO0eBWvouvMzakAn0h88tqZqAjiNHy05/9hHyWEVMRl
m9mO4Z9dEj3ujtpYyrVcUkyT3qb2mK1Dburn+zARtmhaw29Q5wOXxnV29h4s+Sxr
Mlv+W5hG55BzBYgxV48JAw7M4L9WvsLbdJQt2w3RFs9RlSXtiZ3OC5bv7lIm2Cra
bLRmrO5+nqyeRhfJG4a17k/FrrU89dG2C/VLg3e6G//UdE24hVethMhR/WadYYtu
RKp2VQaYMSFlM81H+4F3+q8Pdj1bb9xzKmXjn/x4hk6UldfnVTeohfIXB+BOTXwt
UH/oQI7iOXyth9OGj/TFwwStMa1cHjTnd0ELA8CZM2LXZmk7mawNrmBME/D09hh5
MZxK1oFyMrnwBn+0IiFjs1JEcYDmHqjraCg3cKSfiMU/tqn8YpWiohtNOmm6+QFo
cw+pXttJkaHgJqEgK+0N90kGPSMKQHkoBWcx65+Hh2htC7baXSVSTzuhdtJ9zVpO
eEirLy6BCCAiCnHOGgmckxVNi/2u046RDLRDv4UL/hfvfSmPoDTOYfFSbBwUDnKk
K9dgjYYSP+shuM2rOTOkBWd5fVKHnQnbU6zCwW56c2mBvacaECF+PTYDN+9d25O6
+sdy5xIV+3iMgvyE0396893cHd2BnzOQVT+XON5yUoU6fBh3hmvo8KYmqY0PrsbK
uvBcqBRVsoXPdXLfuUmXG/lyeyaqqfmpY7oU0ua2S8mgN7aASejdnAI1+iFRB2hG
q8r6s12EpwjVEmKQUaCmuGI+iIes6wO2hz4cmDRqkPMqXRxd7rSg4P31uMB310VB
tZX3MJAIK0WVF488mhQku3G2IZBBUc3zBy+rWR9zhKVqVTQSxQq3jhbtJ3QUpvBA
94WNkbgGG5OksM/ljF5YMHctiXrdh8gVJhuByhwfVPrNUaL6FTee1G6co4S0o1iu
uaJsaSS7GTmsQHrV4dTkOkMSlTPClaK8w6iSLzkp7bJqFp6xgwah1CCULZWc7fM/
SGZVnKRECY1DEwVFxDSZdg2C/KgctG8EVWNPjvGzQg0UtUvBSH//3e0FEgyY3ait
nvCs3dMwnIspEr3906Kn7A6YP4+oSybaE3h1K7Q4wbEkWoEDJvY5GHJE2f11X9kO
zAnfp1C2bE9qSCoD9aYrnlHf1t9FZKD5SkzIexRa69ihP0dIjYrPYu4ECYgR+an/
OJnkrThrBswt4VjAr/khKQP9w6/DrVgzN2PTw+ainEBMJfhgtxJQJ9adb1vQj0D1
n5A0KWjVpEc/3KLBhm1Fpog9g1ZGKUW1yrwi4EEn9D/D4jsc/+NHUrYvZFlOAR5K
fw5lsTQMe1uOPIkUJWfyNw==
`pragma protect end_protected
