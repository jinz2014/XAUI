// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z8Q67+zcmdFrqZDHfpz2DahpjJq13bjhzxZgDxbFiJfkCc4boqEW151uDNJ7ZEnm
FU/4TFQ1tQYPkaciwpjEWHHI1kT5Ix2QoNI7IriPn9iabQLdRvMFmvDPhqg8Y7WP
uxThEzG9t7EX5m3T3aNaaik+kxbBeueJSQwMRdQfZHI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 50112)
SfBJ+38kIYSI4lM+Xo3XDGVgxAX0Dn8s2nyIK1g7MKurxewlEGxKKPyRBNIf3UQ9
3UsbG9qp093gQtDhUiJJ6whP0+xS2FcbIiTZSccnzimMZ4DYkLB/qCCj4qrojQvB
IGozOQ0Uk8yiMb1JISAT9YxvWgYZCmS7wpXcblVlmsydKDxoEoxZRhibMVb23Qj+
FgOqxbKdhtbtcjMoKszVjE1yskZwpsx/K1/JnhRqh66gvurn5Fapw6yvXiFtOsO9
06nsJQBoex2AQYaqQtJeNDGIbEX25MVmcDNEB4VTv7im/mLLMjhQLD84xy4ldYwZ
SfsFe5anF8/Z3kQYm87sPsNWoyzrfAgG2rgWKyN+Ijpfy7tsO4xy7gwLehtd+l8/
ImUZoQ57uHpDEyCTI/hC4SXJUtC09XH+rwbtfHlakFbhjLAUwz8e1VlwaUAGMHj8
UpOgIR1+oodPrfS/jwE11Z6NTA2pgPRlXOeEGozMpc5BG2ou308rI2ePMoc243pN
CPkFJ+qzn+Pbp7cpTiR9jJjQf9EMq6OSqBeQjrP5OIa+++4u0STG78JmCf9125Vl
RMBROf/ZF9dRs4DjmSlgCSINgjVvEdjHGL3JF/3xOxGY7isXSZAW8t5Kcsj3gcK2
Jn6VcLgGPbZBcy8VhNG5vOUyAgqlyWl+oAO/nucTT+ZCZ3yO5Ibxpa4FpKJhRd7R
97EO0Fr9nSyGpGk+zzX+mMSrbkIENA93TWXohONCYWCFO4wYzMAL7NYnjGh5Vncm
Oiwu99hK5pcpSKBTAp8c+NT/1LeIek9gtw6lqxWQcRh0h0QqkVLhW6EMjTdbtqfy
65k3nHUQp6ehvN0gwkW0fkW7E7jaR5mjdoxk5Da1i9nwiOhWeoCrTQoM1CbLFakg
/j5RnTrOZE+yvkk56bJaIUFWvJ1/8kyhXZqCjkSbd6mHCtk1v/Q+6DL9UcMwb6tR
6UE7olIgyY2Fnhu0dGlTHw2yRhZC5WShFP9GTT3ZJPpwE9WEwemoXqqnDOrFaFAu
ZCt003NIOPiuBXlaaaFZXJukaBs6wrYVNUP06//hhkyszlUkjrIBs7OSx+nFeks3
wR3LGz6zPFYTDL4KT3iGhcXEZ65xZfhToaU3FOdoZG1DvkPe+VPAo9q3Etf0XMCY
rhzRg9q6rln/xMCH/mC1+SsCjyaJHrwT+IPgZL7vFE7bnG8ByQ7IbFiGMurDDN9F
sCg4imQUpHKx4xusZUpJM2jX6z1zh7nKpO0cEiwEJ3USxlmdowncr2nyrVHkHaF1
rhiRAPWhZFNQLF+J1eLO01Mx1wVcC6C04TIYMzS61wEfESHptwi9JdCSy2WSfz6X
9U7wW9DToCl3Qvbv4jVGTAQy1VNe3qBZcauKm/Jq/8QAVHp/K6Y7xC7UjvN6p9oO
lpVMEHcqQpFM+oP1HtX6+Q8xTrv5oSKWabSSp+CetDzclKmbe5CJcwzyOr8wbcmP
6NeATCHZT6YHtWk0CKgr1qGo+Nd4cqdKb7eENWw7QGzhh68DW2ny0z8/5edzEW8R
BX1msqSUPogZjPFOCK9iRBiq8Ri7LZl6NOYvkP2p39icIxzhhOhA7qR4L5XeSREf
Ims1sqFjXKZzRXbBfPiuDcVgCI4qLDYQAGZRhQKBxuclv0BsXKgFSeTSpjuv0Tyt
WEjpG1JopxSaCeTFU+hXX5dySCraIJ6dAQlU7eU4zJMQBIUv5sEI+ZtPgE/+7ReC
MK2tQtAWWNKD7ikuS8THI3qGv9JD9xi1psMmg/+R6cTuhVAP1HDGtq60wwgeJlgF
Q134BTBIgPGnE1mCcglBE5UeMamiMPFstj8c5FS+kcBQipWpv/N7vMudzMIX8YFe
i0/rqJ/VvaX9kfLb5mwIZOgepeAj0wRHXQQQa1800gS3gk1M+Bzx5DtvT/Vmyg88
zhQaRZkUdhtx55oePn8EHiGh15impc4H5IGp2/T1hbydh6sgit4RykQjnnZesE/C
YnqGWrMU7J2cDlMq/AI4ylYLsoSzHyHIoPElvPGf3n9JC0UwEZybvimdhG9X+Hn8
6Ovq+biWzYstFq3BylL17KlqdMd3xFOD0RCqbS5XYq+fDfAVmgrIsqapMsQYlBac
lUFtlwgK7SjdGz2nPUc7aayhHam6H4gczvSU8oBBDAdbtHel4LSpqEtE6/7/1Xo6
2rF8OMU9K/zHI8jkPglbaClj1vzX7Yf4kqcd01iOkY5AvPVhCaoZUGmbP9nN0D73
F95FC0y1PQmFd8LjIfZ6rs4LsWwG7NRzOY5mCLauwXwhTeWOpYg72CfV+Svm58/j
EU5fIkxCfBeZB2JUi1OaOn6zbI/EY8gXTI9pIrMiwSk+DgdFlw47K31URbXgq/Ys
Vsoclcbzzdp+LUVe4Y7p4o/bFmiAgxOl4KYBWBia+3NrhBNGBdBIeMnOd2NmxxUK
0A3U8sZjHZFiT0WyfjoJbvjAYJNeH3Ihd2MXOww3RvTde8K0dvih2TYLv7avtlYi
1RBgRjT1mOuJoGBXoP6vitjyVq2obnZtTvGXfas4dI2eOXeYNi3TTpadN3IJOqnm
zhs2wLKSC2sko/GnWv7UENb3WihgG9I4kC/QNaspKhogqBJ6ZJSriUY+juZ9/JmE
BWerdLJjgtdCZm2i/fMSXeN1Uaa9dkHyW89dSfkeDBFckPm3u8LVNk7PvWxLKUfe
O2TQBk4lLgxkwvaA+zMJXfgjK0+V5bbJVxFAQ6wL1x5Vi2ObV5tG4tyMXMCqzb9m
RWiTTm1siGtA4Xw/mPCdKlcEQBmjz2PSs9mk/fl3LmGjFwq0PNy5+m4xip5yKPkZ
H1Z0V7QSmErhI+ZKgnflakO9VA7ZebxpV2kmpBZsMZ36BqRGkQ4FF0YDcVgEghC8
WZR6qQkqLc2WODXkmL0s/EZAsclIzkONnz9wfsmmEvX8GVaF9TnbL15lqm0R51Fw
t/eK8U7fQkF1U94kXkaEtpxF8en93oeTgx0bA/6PGkW54zdDYpNqC6Wndr77nxW5
XGMFsp41VZPB8r7DNsTN2igDNRZ+yrIgrcqxBDfEE9ekFx9znoMzK3fyFgxlGPv4
HzDvP9K9U9Rnu7bvKJJPvhMwFtnzUfTgZdElIjEGlZ9EXY4hX1mZjgR4ZWeIKTNv
ljbvdQC0e4wnCIeRk5FaNlgZa6bHDPZZswEl23gGk0eK4Akg2piKAZ+b/c5lPv6g
mfkP8N3fqatvCWCT65LCs9g8fBOVZJgT+A2Rmv5r6YZnco4CAi1gj0S8FTfctKEV
40sJw9GwtBOCSvtiomcv6zkdTRydqDL5CIgS1YxdBEqMVfm3SESnQSnkyTpVOBQT
vYls6PGzO6+coExYieSzI58iXANJZxRz1lSqWepZdXP03pnpwkMt3x7TtaZ+GYNR
/RIj/xDSvLvpKHnKKwuR4ooUxMMvThNxQVUcHfjKPFjNOIC/UQbbKY4U0iBcDTFo
OZRE4PD+UCDBG6vvmNCaDAltql3tK3RAXskvtynapLbN+dpXYQh81hFOmm8xtf/B
W9k6Cp4Wz6qNRLiHtyE/HmCt0/HdjI+fSk8n/o7nRBYXvXJFOYcG/bZaL84IfpPS
wMYiY9f55/hYw71nDZHylRNvBtXcdV10RrlN00X9djjdBaHx7vV+Mze6CIAewGJh
pt4Bm4NPxg7HKI8Vo75rW3ZZi4d09tsmmpWjEytuH6S2DkbK9nvZLJxidTzBapxe
fV909Iak8hskfnrhy8p7qpPJpwcJv8/R+E2LwkoG43oERO3lKsbbk/QRSM4p0099
gROVDAxo9yUwhgzn9BPKmaAg/y1HHHJbd9A6UBcUxYkYaMeDdxGbdoSKTCjLnUlE
8b7ZoXYYg0fSiO3n1YbYOvyS5tNOMLmc3C/vPE7RJu48r+g5ZaduVDnhbkrmpt86
4GxtlWzD+68kkCxkjME76TJR88Z/72sKNozSGqZIYF/bOkxTS6nUJPwXk8tdHXmt
q+e48FffHWOvlfIT1Q+Pz1tdD76lLPBQ5vwQJZs4cRttZBlJbuzWCuxVgutYMI8w
q3thy3aRGSvVPzFJywSOrC5/UKMch17ye1lFVW6nW0ZEPgL6q9fc4vyIoDULZuf3
7V8bgjQCf3FxkIs1kM2/mCoo8XCJIcdyEOO03Vkaw90QabENX0eXa9xHhYKAqVZg
n5QGINJPcYIguiEPnsjulCIo3Avb7mLZUksmzuNzbsE56xlcCDyNi/Cz1RBvGHfk
uSvUae+wxRDyQhHNVpAtbqrd4qC1QEoYhoblTfcQZhJpjUbod58fp6wskF1Y1+e5
OeyuIojzVRkVQ1mmI4ccK4szpVBJYnnbOmKwm72hEdr5psWnclnVM9m7kJ5W44nB
/zvVD83GGH6Ok+YfYM00vhRHHL9cf8lxDGt7AO8X67fNrpr83X+uRl9beOaB+PPZ
jApPtAF+DrAoWScvc+aEeTvxeDhyQmMmbbudDaCfrPS+W0xKDXVRcOSiVd19Y6YQ
xxbYwzZ0TRzlismxhG9V4DKLTPCtPFTPxqpgmMmduATC51HMK2CurGOFhD9Gm3FQ
GD0fBlo0439AzcsvoV4VlZ03LAd2g4/NpyJuTjacPKk8j+y+0VGx+wxi1LxNeaqT
W7jEh8rOanTFS4egxE0+bJalUjUKQXG59eAYWbfa/+nFndfCObeamYVnJpEgpNNt
NP0gtW3tlXPczf7A1DEg1jAUs6RXJTnKjQZuYYE6FJVWKUTR+bbpBOTv5XSje2cl
whwMnRlD8TQXtEk/rUIGY45ao/2IKi8n0LIeiNyvamylKgwnpl1msFslLHwe02wN
DuzfBqwU1xJxgOgtXHPLim+VGMmQA9qFKj8LuXKnURLIxkhCMpP4XZ9A1joxvIKg
eWrHk4lEnTxUAzOAz1SkHW5uUMLoMio/INKZL0eIQY64BIpcGVE00bzpvHA6cT0Z
Th0NmcgtB3gabt2YsMHVPnzbBieSA09C5wznQPi6SBaSDALaiWue7okkZhtuZTfX
9SZOUpXQ1zsWijjQvglQejgJadik4CAWdBhblhxqiQwd/F2ug+izU5vY39h1xLZY
b/Uzrc77IbXXQZ+mjcMBrsVnaZ3akK+zsAoLZmtWpK86OC3annWnTaC4itmFQG+0
NnRYptTDIsFIyfshnyqxAolOfQGxK2iB1vwcle9uLRJzUhDwxj1TX+Fwdk7Fe0E6
qzit0hzKjazKApQNW6z/SykeAtkh1uhnoSZmGiX5r9S029GFlDbzu1cKtKaaHodj
V/x7oXjqglTLwsoavOmQ5mlQ4pVjLu7ctEozEQGTFb91IHtwsX95jeulESBxB8mH
71pD/qzcor2kudGlHOSadM6rtKZF71Ozb2OV+p74IkmWefNMpI9mvOQ6nrV97Ba7
7J/5UIlaDOkiai93+CKcizAnKFlBrtvb3rrbw4XdXelcPXJt7XEgBuhRvrzFGnm8
KtWDTqwGjNWLjeE40vu1+FOaPXzZ31Qqwic2S5wdPXl54/0wx1nF6dapnk8LnxHM
betI0vCjZ0Lw+bP/s6Cv+CNPvv3yW13jNOTuB100Tl9PDu2G3HBtVKkA/iaRk9XQ
4XVoeF5Lyf+v+C8LD8RTkX3ceWGSB//4kPlyjrMLctgbhvwN67AyEJFQ91vH4M1s
HAI7cYzxaYIFiBnWyEXJlwu3D8rf2iA28FV7OYR4zAANrwoC0LP8rstNOS0ow/Zh
QHi7ntD9mn2EvwgRj5s9Qtgtg1FF0jIHf7IAlxV+AJAPHU0dImdtQdCAhixpvoDh
rg7lNi7ZsVGAjZ7FFKauGsA62upxL4L0CJ+X0CShfmtLIMRyteOL9D5Sgp1J442Y
DnYm4qxLEJs+SiMylZ896B8NXa34pOZ076jamwMff6jybTrtWElxq7SKQ6vlIhDQ
Na+Mj8+k1BPfZkE3NqmtRI669+OMe/Vgi16qG22Edq496OvcVd97Ki+YQZj26oaT
Txo0x6cvdUfxmd98NSZBgRThm+JYsoY07pxuFW9d9oIznMZ4+i3Azz1Ap3CE2/dQ
apyzP7q0xXV/5+Xv1yslFWj1r+3x7lmdN+rGEZT7bKc42te1l1p9y7yfXtV+oT9k
xLWWBGulfS2j3g3NUQ9IBDxPCJuf0Ax9aUyB1xWxeO7w8exyFTmHl4hqL+iyjF4F
gkS8a/GoL2bc1vu6kSsQYiTbEd6fUpWD5iFPMmeEg7rbRNB3d4oebsyIdHoomybB
tGG/OArbYBYCiiDZ9F08mmYP853ONpU0VJjqopwD27bmuedLNii2D/cG5i0K9Kp1
yTvobeOl3g7YI1igTe0+X/t6BXSF/CsX+XNdN+Zcj0orKGfGZt/J7sutg40SufXH
AMihEnjeTaPVxAd9QGXyso/wpmGvIlWx3aFcdeP/kZMSFNpKDRzoC/Rwq6owrq0d
aDmbodAMVH7/ZkIpIeLasX1wJ2+4ZmpQdpR2EgnN23h01c2ki3bZuNs9jI84IBbC
3Rh9p9sYGmGFzyp7BinPh81whiwLVxnOmedIMl4zUhDFi2uxr4aTJOfgwIQey+rc
4vJbuootztYEPZ9UCXCNkJaDpQyev1y5KOJlYipyHY0+hs9hkNBlleNWHBzppfSe
+xns5xVY6Yb/ASEanrRVbIQQMPqg//8uOC2hgAjO6j3lGgngLF4fgXl0nbKgtLQY
EoqZbi1QOlQK3i/r7IEMkraHRvNcKC4RQUb9Fh/pjcP9MvN+rNnbSmxx2+i0sTJb
RO7tJGEbp4gBk/gQjauxGq4d7661mkAcTC18P4A6u3CThfT2LGFjniTWZe/DIf9+
J+nL43cPYxgG3hGBUUpsuso32Y0pAsy8HPWkfD0CqZHxtVvBialpWZug/++MqA7f
J74HMpxIn4hLXTUUIVQR1WCCuDtG1ViBDpam+mRJkg7njbG9M+5Hp8dFx9eUooVK
l5hng21eUPEXO+d8X7A5h1ap4AAUXpLLCmke49YcZ9eloasDVWPr4OO2eAe/WpRP
WKAYqayaWR8rhYPoxyA98xaGTzj5nlV3/99iXnwrsNaVtK69Jbybypfny442ltjl
LXaoIWebkqQVwK0RSCvIfQhMDoeSfZebG3ADtl35OyzU91Mo9KeMyAWztggIb4aZ
diOu+FQCnMyZ4+2EBnN2sAFaCz137/3nr8A95p7xTdQJ+Tpy6rIxoOrRWHZ2Ytk2
8Jw3hgVyYyMSaUJJWMHWT/JP2XBMHOVfqqHyWL+ztUR+qJtO/aSvF14SqZYxLRgT
Dhj1xuYDtCfLEKkAjv2UE8uYrpSSDXMt7w6WjpbvpOCltaexMJQXtRDI+cIu6PgP
7qG9olKjnDXyusrMq5/Ki1wxYVjgR/uTlfwcwMsus9gzTKfo8lk+UL8WwciHT7Rz
FoBPlbkqLCDlPJ9/elVIVtucl5BqDXNdpS/a5+ix7U0ROW/eUZiu0pikMbtOteM/
ZRL6LICcO4U3HM6vIiDvM3uB6QYFTVlOsZ46yOqN2SSZ1rryZyW9vXptaZ3sLsEh
19teFpf0UBPrcCamWNX7lZcjVDaRutO/E76k8vV/MdiH6KdFAp6LaBhY8RUpa19X
CQJoq12TDfU+AXwKBVeM3cTqlsPeald9eiWfbabdfJM/vVPCiDm9elEiEMVonwc6
dtemaXZOjEC2gwNMQ5Amh3sHXdbgOcvDxSVGBYoepO6xAdP2l6ROu2ZViXx2Skfv
w0uzUicfzVOcMS8/UGz5LbSbGeFWnUTLalUC3i1uyw1ATYmjj6MYg76tspIBsLVP
3iTa8uWQ17Kd60+DqVihHV6kSgv8fyG51sbDqNUxh1AuujZuqqvoZGS9Y4rWSu/S
J6YfKy9FAqLuWLBUNpEeqHfv2Ku6BkwRLPlRYrCxO0rmkpl3BWVAY4mvRT2z40FK
KCd9YMmQ+9fMQk5sogThPvFXiCYvUZEioNtawqPQdWerJKpAs27MIlQWq69BgQ9G
7bkEJp5w3OtqMi6dRKepZ0lJtOySDm1AaqE7w4rpSaQEIdf6wX2hGoaOg/dtDnQN
Hzh/yd21G4JXRGCaHctmQqE7hZ9u40/lxDkegEd1x9lPsOSfpiPKvjUF7fg6W+rv
UYW/YDjZ13Y765Atc7f7rKWgLVEq53Ina+9SxmrL3Uh1PP1JOxfc4Ym0B7G24y5d
ywV5TdwvelkLEtpsIfbCFmUT1jUDZMfMPrkmR3w8D6v5k6PrNfhHVr1VMe9+JmN5
c4tjFHQYCB5PGvBEC0rdoPNYxJpAu/QHQwqZM2r/SpjEpwlPVgRj5h1dP3a0Ncc+
aIq1B3atNnDnQDOEZPgQSQXS3toN27U9cGj6i2S9TnRoS6UG9QyJEkFwU4S1QfI7
pmclS47rMNFyw0QiqvN97ZybSs+aHD/Yc8QIEDUnZF76MdKW1r8gJBj9PCS9XKxV
yHGhv2lM8E3T9GiHVG45HWo2/sYXX4LddlabFILea3i5aoDIOIJgXYvX1EtAfmLF
2aSa1ppdG57W/Z3/P+KVGvODSViSJ0o8sMvIAnvRy065BV6uOl1uw2SiI7c9U9OB
YStRvEBp8rxQUJ+qoXWxYFdcqPr0PqN32eRM5MX+7l3fVFYkX3VO0bDQ+pggu+uI
hAu7j2FnNtj3R7ixaxglH+py7JZJVJbjG16FWBzQl+iNVO9BbHoG9YaAhE2iNtRb
QwhhP/7BOAn8XyLiTwJzv7Ucqovn2nEBGmJfD/4c+ITB5+LswNK1Ee3SYFJ359CQ
DV83rxxpCorw+IYcxQKxI8URMeaYpcsyMJGHHCvVfTg6o/LmPkgCdtPBsUc+loVL
VA6UtNpQR9s+WqbKy/LvxnM853YvcalSnIC1auJlWUVtfwX0/koJFSXNJ+k6aPmP
1Eek1/I+MpLwmzM7V5CRT1FF62f6UekU9LtPc5U0JFzV7A8Pg7yAOpE2XtOcoZrw
08y8tCM87EJG4glV0jwxi6dEhyJ9o0QtJuJqae3qrfFrc4ib4pyry5NDnn3yg+Io
kI6j183yojrs4aAXwC7G9Cv8WJlok99lxattfroVqvYq6pkA5Msjt2r/zR4aGLzH
ymJTMqobvBkLT49tf/pNWmsVxgp7iYNC9mNdrtzpi6F+w1E+TqnnkXZ07I4Edm2L
WzGmlbSpbRGKS5OT60QTh7o6Wc5ygGiEMgj+Z2To4WfGIQBBNjTHedrbyH4t7TNR
BYZmoMm4flkgp6CZcnh0KAVSGFEQ6AO6EeqEp73/CejMMWtaUjK20UlhOP0TnX/4
qpP8lZ68EKMhKDDFpBvBEPi8XzU5CzGu2wSlZl86+ySqqxAHSt1JAeB6N1/2zPF8
O8iFK8BdqlXjDDJ2fTnYXtL7cmiI7Daw+EqvpR/0D9jiL4n7rTl80CxMkmcSvN9n
xtbqGJ6khN4sX8kfT/D0U0ioqj87yaHf3AelF9KXxxF6Qynz01beU4Pcd3jdJnX/
e3q9CfSqQLQQ8r0DJWybrOFaUUFa/YVEteZhJFCRDeHOyR67UG3W1ibIiR6N85E3
yxTwCOMuIzKaFBNMEbFjH0kgfmPOMaFgGqku5Smz7cnQHRLuXU2G8F6+xLyV9o42
BwPWV3lVn32CazctHSTW4coDWQpLyV9nD0jU/yrDpZmoTPdMv+BWNl+suTIUJFAd
zQgvPSQZ9avmo8k2QbMJBO1i+jcIuN4gyy8mqV1pIgO75EzpfWM/NEtHF68tN+Ij
cYCK1WlpC6A96CTiAwF9n+kVU5OG7INJM9li3dgo0OZfKyOFCkk4h+RqvFdgG4E5
rmtXDO1Xje7MoDLlTJXjaF/kJP4IUo2O6ouAJdek+bN3MzYBDBe9cgbUY0CH1XiD
PROxOwlYatWslJwDfrlpCbRSaYIxj8XuKjDp9NXz875eQwWOsz+KurR2R/cqeStu
48TiFh1sOmx9/88XH8tPOcmZXxXPHI9dg8+x4Eazro0FKJbPTumgMlb308h7V5mK
p63bM+1Lgq8C2A83Q5tzN2QSeE++x89oKgZENiuTms9u5cTtmWG1HvVFPGRDT1nk
ktK/Ofa73of2zarmsNPAGjejWhneJIX2AOkcbTUlBOJ6bwyoGyhJ0YX7wo6a3xCO
W4mQUZrjaggNKMXIDTh5ydXa28I+sJId1AS2vpQbSEKoQuRLM1julKnTnbpThIG0
9/mAtouhlcs9QrP9MQuOne85sDk0NDQLFyqcw5pxbWiIifD9ikDw8HROJ3RcG4Ts
asMS4qUYo/osiS696evw5RS9sVduqqMD1xIoUYEnFWvnFAca+2cvcgBYPBM5ZZG9
aiKq3Ul59y8RgHS0wNwt9ZHH5a7CbWHtFjbCy6Lfee9EOEjlvA5AgFhjBELlNnIE
GJCvgHlABfgpFyfAqZwrteECQif6xfNwHJ3xCaBMD8da+7TVo+MkWxT9m1NMkxRi
L9p4G92PsrITYBpqmG7IEX4bvG0x6Wt1SRdDOvLAoCIif2qvSwUYpQ4egoeP27z9
ZTMNCeuN+iRUNy7RDNVn7wr3qyAQPoDmxhJXjZUtTPjW0D7aqxHUgElG9AjIFFmY
0K9CqYWV5WMX4dx0ACIZ48uiEImd2wSrZq9i3z2gJSEziE17q2r7ap4yluxPZyc6
Z0xpTFZFt7Ui996zImnYCaEWWj0KHVMYijULvhdIYrQJVK8sLHs1xZikONQqY517
JvNDkgrKsDiN+MZe7fyRTMj7UmuH37NtOtZxwLbLqGxU0XaomfrFXCVcv/VrnlIT
AIAtnRklNmdtbsHXmJvZysl3oKaTUWgp58PaSIDt6EyK2mKTIwcrQfM0t1ZRIQIM
jfh4uz73zN1ffbCpl6LA7TeuEK5tvheoKK3z1sR+6LIqRPU65WjmI6/fcX3qx8mU
1vvarBArcePqHeIg8x1oHb1XcHQ1Y5mDOMFP5MXWbcj+7UkDMDwqQM97YsC/alP7
Txvxao/6SSFOiajXf7wJSgUJy2AOddwX9RYaJhajiy0JDOKCrh60zwbZzGkfOsf8
W+2FZ3b3OI/cq85OfsZ3GPZeOOhZCXLjrkjdzpLMl4fCloNWNo1f5B+Ke7fFKUrV
8I4pSxrGpYH2ljiSKpRqEdSOhBW2j0tOZC9xdzWtmDsP36Zf+hLWbwKQYFQk39yV
iPJsaRW9Cq53zgK7CKrixXWcMfr2/D0pjvOeo+OUkCE/6w8eVXg0tnL0eys6uJtk
jffuInfAGgtNExo/et9P1MhThLyxP8QI1xw6j7zv50XKbqHouVMysfqSld+BZ8r+
K1iUd7Kzeheb2nqz+1/yw/CSBKrchK2O2nvxNL/Hv78RveuXmqhIzUIH5dPu6dh+
MfmZ92A//5nrojX3k/9c9hOV+F7FIr4KZOfdIWqaqC6sjiWIqkiYiFN44OWNhTBj
fZWpUE2dbDiZ7vMCmB8xVDeypIzkVsZLZCUu/XVU1LDYqS4QnUMs078a/WqAoyW6
BwHi/T9KIZWLicbmT2dH2RBnLB9TPf/SyBpdgl55GQfiJBMkQ5lQJG8mv/v3gubz
+Mji4zz65KdJRKrF9QOKmqoZh7PYC/eWNcM4Qw63W6l0SV3A9r/BYFHGL44mx+CS
pc3Z4eg7Z12cWZMkNfEzKEEmWteV0wpp/P59fgeJBYIhHCb4SdtqQBT8lfx/u02d
qWc+4B1HwWDzqMMX0cZ1IuxxfycByz4k5p2F4tlqoe4bTI9fYik4H8tpRbUu6U34
BoYs0VKGmmmEUCbt6zDxbnhfNM1ucuE8gTzag/0X5V9VbdkgLZowaJEWW3IbotKQ
iglYFaIoBviFCKA14NRyaxbd6Xrt0eYo9Uly5ZUudaKOZa1zYWWrahv6gczp//Fk
Vygy6epfIXkq6cItJ29XjazfG1XGhtiBYuA7gaWC2X+68Cibe44outDIBUEI5F7i
43EbXxVxhS/OzuknwIzx+wbWolBCvy0Tzgtw1grwTbQnlnl1m51z/XXeHL+ZYBTq
ZhI0gEHTkWVKFp6d/9vxZiLOqrVPmbXPiPJzQE0YUSMJuPvgCSoVMsBk9Orh3WMD
TLDu2+pnPrsJhtb4oH55NrCkS949N0Y7MSylgur1obvk4alHUe71AQDw2IG8oR8g
f/UV2rRluI+AlKzChxy7fGqsfZU9WnWylDozPbdYAclQnONFCH6kBVTKKArMmTdP
VnSGAJpSJaelyxFKy1rGOf/KWvQb5jMQA18QtbyDysX0ERXJ65N7POjOJzxQ5JA5
7oc6+afN1sO2l1/8U6XsjFci6yyDxtnwBiV9HdrX4HIvqOxFihgsfWDJ9Zn+bMvq
/vAkmdYcC2y0/fIEnDgG46H0/SVmYPg0g9NDMllzv7PD+hWQlpMTIZ9ZN2DPGcOB
goguAlyfZSDNPI8H7QWny5fYAg1+NH/EoDba7huGRtoWxHBcKHe4NNfeLigExb95
3LN/Hgk9iLDGYp3DBdEaAO0Vh3K5c8q0mWLjftKhX+JLkpT4pO1pLI0duqrSgr1X
3f6QoXiEzK3PCyCYnTgJjX/HlAMa+xoHysTQ7FjEW6VuvUvD42aUO0mt68dibUPe
ZffpLTK3ls+s0LnFhPjn8zYx4/qgsIrIGbK55OIqoQzuUMELInQAwcvVl2jJ+qu0
t+bk4YpT3Zv7BvI/LZOmpuj5HV7NYQUBBgKyQC3l1OpKgOZ5VSgKpfH/JF4l0/4d
cw/WrDyvP09lSiGRUrc+QfCwqomHWoLPbiwreHK5jHCYkPDyl4DmPccP9jhqkEkj
laXp4mNFugmyEOJxuy0Q+i4wU2fVDrizd8gxDsRCqIwtVimXOzT0fRlrjTLXLkWV
fkiO76PwfpBl2AIoXrSM/69X9sR18HRLZMydI/aX5AiE2fS+yQfez3T2RWSZqY7e
rK4ZMIk7q5mpMQjNJrcmrXwSMkoOK/b0u7dySQRyMTkRQcs1x+9VDhBYmlZq6Qh7
OhiimVteMOM2fJ5X7WwbSt3ylRbQHtspS28xy1NX8HgHedOOP5JmdmAmTgpZwY5u
6usAlVaQcvBoa21MHYZ900DLPVXy07gQW+d/piTU6Zrzr4ovHK8YHtU7idcgK6X6
UVOSA3lMB7/n5zb1fRLxAgQYoNNMuIeGuD43zhXx4fgtW859Qk/apaT4aR53CFSt
j1cNTGa6Uv19SIBFwz6mULGCwmelOQCapksfUADR9JF8MZXe0yxrAbp6E/tVP6Cx
hqFcd4xoT6bDHkGq5F/Ge5bf9yitXxt7SiNksd6AaAlOZRdlEsBvaXtK7WV+HDBc
aHK5OHJML+Owi8qqCUHHxuzSbxPcCwsQoyV91NlOnm0L+u0YP1BGbjbzoBQ9Dbzh
7jiLmkZfj1feQzDAqRaxyEhncElkwJDQMHRNLe2mMCD8hciq4VP5d01pahQpAz74
tDd8Nsr/TQLutfgPkqPYNWorTSZ26I5L6XCYs8VLvnWGYGsxRzBt6UedY9VJV34Z
VKwB/AFw2XrccwYFRCeqzxsV6NS5sWwzpatJYsubOBhVM+pTj2iHencOUbCeFXrW
wdFd+Vk71CRcDGsrHEW7YhJZqV+IWnwQce33j4Hpm1pmukqFl9ROThByi2TYSYt+
SJmF35uJjxp8arnkmAu/h2k3yaRy3pfMTxESZBTue0RTu1+4ZIc4Y5rC1A1/2RDR
5g9LiDyta2n9vBYn1NIb7ZBlAAedPrft8Pw/m9g7fObPl2c5407xa4GYnhdLVcl3
Tbz/bN0ti11j6eOQj7ECoEcrbe7xCMHhQn35ZetjfDYcdfDnbrmsoAYrP+UC/oxU
PKD7Oklp+B3rT7neP+XRrqk3GdXsrq7JbV3XvAj5hKEvqAtmaHYd0iD+DRqZdBbV
8yOluhMWPx0p9S14hMjRYSnkV1/KORZyxffAutlQzqTAwmgKxTH/XquN+8L6IgqX
pRqG0uTZcEBDeiu+3bIkayaa34AlvHdCVRlmAZWeBa75XeFC48eG2EUEFdw5XYLS
GOI3wbIoH1i/Agk6fu8MGUN/MI9wrFzjM0nB3eGjJjkvWm/LfP/H7+ItTv32NX5j
vjanZmkKC6DkGPA7tZ5wXHzhXjoyJ98XWLYrrwLV7sDpF2s5CDyYWMPvKAs/RX2e
lKALEOgI25rS9x8daT/7ed/wRuXhjWr4Ft0fQEi3H6FGgK4LiYcz2YU7X0DfM368
Q7pTJfCSNK0oIe9UYBwhMYZSyJDSWz42Unvu2cobn48lTpI3WS8DvPzQR1KdZA5y
btmgbMRQYnOvVwDiZ9VGv2IIwpmO6meUkS2Cq7xJNJIeaPebUK/iDHzUqHJ1r/Ix
NzXIHDfOq3h9HSA41fz/zJ+6lS+Fzv8JxsAxMurH+ZBye8XWCmiMWWR4aC84GNSo
7Qo5v8twCT7DOfretmMB/ZtXui/JAjnvfTd4GR7Y7e5O9ShFxmIXRw78GsJ0oQj8
tfaKfuo87Kjtjhk1XLqAa/5gc0hhJwl3/hu1BQfUh85FJCOK1ZmbwdsRbFxN/7SL
kdBHztnOnU3+nd34FiywdIkvV8Wsy6PAjmmmbxO7AF0PNMkjjjTHAzVBoJHojXED
fGj2l6Sq496sEbHR5/BRvQT/oyPsaIgPqu0HxVp0O5tDIALiTDpI7Z+kK8p9f8nh
XoQqHPSdwNihEWIHvKdi1UC+G5FpSQaB49zyQUrM+mhpPpkr5OUa4QCT0T23HHu8
VIpkb9hpkA7yxxE9xQ51tdsk8z1YJQ1RYAUYZzLYkj0Zd0lo4gWX+CrjQ35SSsxj
Ag21j0EvoC954TM4HBT9q7iktuK9EgvC/mGhjKwikI2s1boXesfo38GLq2kYN22A
zEdzXbfLVnl6ul1mO+R//+nHOJh0trJs0wYQAhZjP1vuetxOcP87PItL6yJnSPqT
hGngsgAlK96r5+0JaMMow/vPxLgqydEDgZliOkd1GopEsZHbyOiu+UXBtsd3obJ9
WaZKzH+UdmymFgT3ffRAA7lSDHE+L/7b3G9ITOIuhNrmz5fVZc0awjgF+KkK7Nka
dhEbpUssDXuBqg+Zywm7OJ6LYVFmK7NwXdca1SfCKtE8OoIUTg2VhP0i05FdoJMy
DpLb5GQOlMJxWSN1TLczH6zI+umBHFONImR32Ka/KDJt5KSh5GCBqJeLVY7equGG
YzsIw50WGW858rdX6AJLalXc7UzK48YwVuXv2FB2h/TsA0a23TyS6v+UIhwM2T04
IY7j939woxGwTW0BJ15ScgC8Vvw3FHSnEXvnvF2+F32B9Tby+VcKHeKlELvcNtYe
5p+fwkamawGVtUL8ACnaspfMGVJmWj+qAOSBYOiuf9XICRCoEf1fzSLxYoKy29EV
RA6uqGqYyFzIm4Gs32rSxKRGByAuDJaftiBfEtrvEsxD+Ia4p7jEDpcHoRtgUZ3h
iDCETKk34im586xs8KFR8arMDCCCQX+8fZaOwlwrplmQBtbRC5XGX4kI1LCiqubL
IL70GBabX0bjBxW3//nLEcqmfZZOPJXgcn1TbdoJnTQoqt6ahd7rLtehDnRB3BKI
0tHqh0jaMao2SbDbk1P/gEe5pXDkXudkgzBSljNAhxMQE+zid4/6SQB/OCbl6nxD
acs9PETEXma5WBVWXwQdB6VoU88phyjxTLRv5bzUK6VIJFuzDtB5g/u3qayzTMgv
Kr3B1gEt5oXKdqiof9BUG9JFit8ZYRBwIlpA24OFWBdPx1oN9uZSOiyCEFhDt5bW
lqo99T/Tw3hJtfQ9Hi0bTN4x70f3+M7iXyj3eyKEml8n+9HXNABloqXJC765yG7I
mU6vYJA55v8FgjW96M9lqiQAa5WVPsoIH3TkWL0my0O3YLWsOFadYLHDOlHXmKFX
mtXFlRz5V2Pgw/A2WZViez17TYMrQ3u0s5GHvWaPZ9y1WbBrtDMpNyA1jBoUMjp8
0oL+yoB9LFxSwJ+3n6yO4EZU5CQcBzBUERcPOXMr/KGRTtfVDbqB7HfapJQYn4uP
HZKMR7H3pRlf+oeDW+iUPoJ/0pxCw8lMLiz4piAFNuyyByf83oZAzuOLb/0yrb2T
eUtkYzG1GvcLGvJtfycvXnddGFS6z24Hd9DDkbKKKI17CfED61V4TL2cjXI/BN3+
mtG5IlwelpHMPALl5PD/5unBnm0XD1NIMktSRh7S5kEjwRkcuwUbDRgelDWr6sJs
CpHRH1dnmclXz8dmIKQwZ1dQa7UJ9WTfjZC5QInDD8eAEOr9ggNBjELVr4rtZNCO
cP4HArGyPYI+BFbW+YwnSdJTDxXSrQ7g+iJIn7FbMYgPpQktKW0DJo9eSHzoYa4Y
FXlACMZzrkYJ4TlIISw9Xp5+4ap9wY4V443kniAm43C0R3PnUs3fI7hcZBHh3Qrn
O8rhB+FrldknK5doTD5uFrZhqHkPdOJbKCC1tSLWWVuNBO+ifeXgH+zNttBlxC0L
EvKTrObIi/2Ydmr3lWkaETsUzoNxuGd89IUxbSNTeFso2nsSdcaWeJ/9WmQ4QvVo
veh9Yqt3l9/Q2+pTVDo18BHGX4rRRS8dm0+LLUvzZI029mNZ3jDlI30UIKYUfB/L
AwAFe32jL3giwjWlmoSwt4zv76YzvsQ8+DZ5Xm2oNCiF28QHBWi/BbejceugSkXB
4ZZubKmrIf11SBpoqfh3XGlsfjS+MyGeHa318LEp/3zSCdZ6j3z1vQBT0t7y9ouS
wZVzbmCXWUVdMeAvX67vPfYGe/kv4VgRZE+zYqxL/pCDCvByPFhwCXx/e0ui2UaS
yoJyq0AqePYEiUS/5ie63LzCTTbisG3KqI+Fp8oJvGYiHAY8AOdtUUK0myT+jb4a
/H45HhcTDBZNhVBSowKo+pjgVB04EbEOi35+tRZUmOUofUEy+BmO+mIGhXOfUk6X
Sx6SmjuSZQ4BwQv18QY90XIFDpzE5Y2YqqqD3DXRz6kymzvTVDRf1Jov37WrCiJD
f8sfMlxZ0w/rcwqMQyKgzut+vZ7wtCcpRo9dHf6pcsKGIFhDkKMg4ZUa2/+zcuio
OWVO46xcJHtqKG303EDNU3YosaIn+KQMU/A2T6eCwqqeRUNmpnySUIBxTyPVrqs6
ZO5cfx2H1b91y2vyKFrJCgkAyuaZPj2sqAbtmW9JtpY1Rq7wcOwWzDDSh1qfV8qe
KZ8xbdEesn+cGlOyw5EhhbVSkwjbpLIgni2qDSwQGpcG51CZlZwv2SJgwuTsbXaw
Idqen1gaRJofQM+eDIb8+qqBkZPGCX4eBUvsbzAo1yQoIpVG0kSmZYUZj9pAmhDG
jYGaPBE98LeQ1pOUyuYZN0k9D8Liv2Bl/9rVpzPe5TLnOJAjUMzTp5mx6QbiiOc5
CleHUGC+fZhjqCu4jwu9Aa9c+iDXkAUEz+dRKrBr3q1BEXMdXLoTg4ZIcFScFuto
ISAzlRHyQuqimXeRV1XLAkkSOgBr+mQgZk1PKNWoO9yOFiPFPbwqaJo489OFBBjg
JibQNbDSRKRfBpjtjR5DqXlGE5TgL3nZpA9tFX7clAHBjpmLppgyGVKaOuItQNxC
u2ij0E4UHRkffciH8EolJf7mtG0EyL5YXnA5aPV+DeNwVu9OiPLCg1FiIeXPkM8Y
eywGZrJCpf6A6v398YM9e1sc85x3PE4N57WJSrVBXFSXyTDcQg4Vcv0PlUqC33qv
zb78aVy6s3prSy2oi/09itvuH/xQ9P//HhGRFSO4+SthTOmNUi2NpxCggAdyaBaN
gEejK1WBtHv8Y44PZkPXBtY4gEUqXMM/7LCsstQ0np//aGnFgJqfhmlnGfWGt7Le
oAzvCZFdvGDj+DvLvjjzVGBgTSW1R135y6zGIOoMWw7CEi6M7Kps45PgvvytVoJb
xIwUQY43gMqzNDkQcn5x27KSOvmyJq+VLFFnFYVimDVBW/r9vKovKmxSP9biuaDF
LJ20hYYzw6Gt3KdhV4phFkFG/eGwJX9Oj7V8XHx7avtacmKeF8ykDkKiiv5e2Wss
RSqVcU9URuQ0rGQ18q+XVNTRVSsfY/IF+PFdhajDPVyjB3SAaLh67YWh4MjlCQR4
gEjalE7UwXRjH9xegIv2bLtkHM/aH4TXrf/OLH7QKjAMUaZJk1U7gSBoHrrJh32c
Ciue8FuYnHm0wec13eizMTsCW9AcFYkXXcEkN48QqI57lez04hKKpWzyrY/jfVVc
/IO2SMH9ke3BQ1l2Ru1V21+vOWpu4xuGFzYzM0nBHnBN+41+YvyfesHza4LHLwsh
Vn4/RDr82ZEXju020qDDTxDqDOErz5f1kKqS5FIJFLflrpBBYkkPQinE2UjJCCMi
ecUyaY8Z0Zp2Alf2WOS3t80tc09sHes60YgQ43D4ZdzvunvzMqMN0Ujn7cmWLXP5
RT8wISfWgy5urfj0PVLUvdm090wSgrEdGV13gBPKSGNLhpJWLatyTnztdMyHPphz
yquP0HLVdOwGXYo7h3gts3i4Qlelc/e/lHptpdh4D5RdACzWG6GW0gGdqvOD/gtY
owgGIUrtpe8ADhsv8xLQYXvGQaqPmY3pLZur05vfur9DMrbj1XqlrRdFRcONjbrH
ld+LhHfRAT73fbXGMplr6sPc1pqUWmDPSA9Z9ZcfZbdLMtVwuDlC/z2+MzJNGVR2
RcqiJKlx85JTe9h7ykoEezm+43xy2a77PPl7u+sllV7xCwLOkyOU6yQa5zSsn6Y0
ksarQzi0aTUrcbMUEw6wwdPlreMq/RX8mO0CYlSxKYjkwf97AtSkMovE6ObyroZ/
e6+q1OoUZa/U7VBGnc2q058A5O3wxhJe81Lc8vZS4P383UMMSe3BINzY4RSYA7Uj
0Kg6OjMtuGytN+xTmFYMcg7pEkgFya2KrmX+VZ6dKb+wWExUs4L63Sp6K+sg9Vu1
66G27AqeTbp4Ud2D0PoZahN9ZYE9jKuUwkT+YReRf0080iYNp2Fpv2Cl75Y8YXVU
4t/nYIVwu4xAzkmwBoK4YuREk9/ESQOjRzALzhLoaBCQQHtnwazJi9iIloZensdf
1kq7rSJXUZ7+n2zfnCMC9djrVYExZdOpsghCl/FCPXtCC8FRk0hKnyaIp0I4w1hp
jRzpfPX95hL8fLqAkk61AbOQ704M7IDB5v10nGNC+xYqwVEyRWBFkC3hsaFEVxvM
kT4h3Yf7bAE6gXYwFrqb4LsSpdfHCANQRO03woG45c9RiTIljYrB45JYwslTJL9j
4geEREUg1C7EvjA8/ycOkfKbyeHlWOd0/Eo6Yd+NSCXpHG6AWuxdCV4KlQ3MMjIx
KVtCVG1qSQ/mXjWwEOYQYwa1gqTOOVGGaC4OkE55aH2LvXarX0HjkAuSss6ie0DH
wmA6DnLk/T3c2gNQKeS/R4bGDVD4Jzd87ylmUrvYvrDtSZAc1exvSTLc4oZ7ufGX
Xf5OcXFtaUtgfthCQm5bha+iSThHDJYymUYUOvtV3qsvFXwKV27WzoyZj7dlgmoB
NEjtau3L1Uu3aZNK0Kx0EYkw9VOmKldgtyK5kx9cNFKhPXrl3rA2P2WuyT6YNRUr
+9qGE7JT7txR/yqVukPU1k3oQPa4BVYjFL8xahHo0CRBdjE+9ykP4mQw8H1U2UZL
GVpexsEiGUx3sYcPhtGG2TLVRRh8RcaQBdTnTbT/t9P0X/a6xRE3NQPMmtw/h5ot
Zc9OR93sai5zKi3Mn+CXEE4ydguhVwjOzjpCXZpHZmar/uCkJ9KetfYJ/hMW5QSS
govVyDtKr7RvxC4dYE7lDXEYMoVAvzt0qkuGzxeN38q1wrHAwxIu3/ZnGAWw4MbX
hRDbYmx8N9optP3x4q49Y312XC3+9eurHkKBQpFRSXWrQmnRB4L+ArEozgrAuRZm
fhAC7UbCYvi2gZzO98P7OfYQc8Hjl29UsZZssR8/W3X16lIEgoPWrgQ3xVfVjJPH
KFAc3NvAQ/D5PpLsWNUbnWscUc9FiFOhYJFCeI6sRCqS6CKNOJxRiKx0BAa9Gvwe
+58jy2/fDRS2iO5xiLgN6nZs9h7kY8Hf4YK7+Q3eQZAEXZxmGXuq7nGJD/NJQ8ld
4Mfnz8r7ObCXzqdrwU2E+zE7d8HXvzs5NLM/Fd0kmFWc0jWzQmwwatM1tgJdRrU5
jNN1BTfeVfOU7CbxTcOC8tsS13/J6xnrtG8UJfgzgNvLPiCAa+cHYCPXLPQaKPGP
SI57ur8KlwtzKuMRx5VUphKCxm7flp9RrHgiK4wQyApzAFsTG+/nWPliI4OSLzmQ
gw+nXeeUccrNOnReMupFNFgntKS41C2PqrJNMMHAQbQbeLhabDdnVGkeyfoOXI/g
IKCtoj03HS/5581Af43XFOirdZSibWEFzN7QS9/+/EWSOjQKknL7hLpm9IkEni6c
84+PPRM0KR3KsSDxs0+wTHe06ULpplhCy81dodGhJr5ZdHzmsOjGnw7HGS9RFOWY
LDvN0Xhf0HFZKAROle+TPzrQ47SBNjuCDv1ffeQYRyU7C+ic7cKfPt5QeCyOnO1m
NqRRi9TaI6LoxszbFxFr97XrGLz7aKd2RDbzfBsdA/mk5QjSlxHjVrKg/LLGC2HA
DjpRMF7ypHjvJ/pzJmAbHFLmmscp7yCIQv2QHrF/7zfXxr2TW9iFFlJUR+VAtJu8
kOKnZCLTeZeFiv5XMVDMwuF9Su/LQ82kmk0lIGqaZFPEOnWqKU85Hf8mM2Opqzrv
GKyjV6z/0W7GjwYmFN+L32JofdyL35b4AJoKBM/3r/qJSVZwJnvBHNLnpi/jO3nb
N43xt1QqpLVfCc+xeGo9mTm3GOHKRPNc+vJvdNjPuySSIZe+3GLQ0eAXJvrjDqjZ
nkosmzcUDsenO9G9iGAJ1kVdSpm8t3om4Kb1liQI3PRPwH+b9HtJU7VbgPrYejO7
aYy+YBM0KH8MH/kInYEv21QrEDlTmhXPU2MDjxC6oqihLsFEEK1EIIB5YndN9F27
hHAKFQxF5O+ECDbxin9b/gMmzXMRJszjuMUxMJOsf3eYrdk69s80667GpYAj1tPD
EZkTBxdQiYUVND+bpoUPV/eD0cdcLuSXm1kzyvA87vY8W3eiivCi7pBnzuW7LTDR
T56QoYR4cCkJ0y0Z+yxl5/OBIdT/yyS/yYIA8JG5dmKNPje43dV96Ac50LLfzsxY
QdQs6Rh2/Dk792tBfH/QD1DCw2EHvyXdx42vmldrTz/4GfUyIvrLL6bUo1rxZn5r
0Db73gLM7IQpNYsoNts45djjrdaKSgKAp7y8gY7TK2Zz6EtqP1UtmhiGIndOsUsq
cYZCkS65uUoNRiIIQ3A4GQ9lSntEbwC+P0z9fMkVaptjYQ+sJGPavSGlwhwI1M2f
eMM5X8Ed8P1uZW68AfwhxI6Ct/ZaYfT4kiDqU46dtQ9iGrijdYCay1D6AzeH7Tt4
SVFCfftln4/fKVGUB3dsenZps3v+wAlnaJmDwkUeloUFJfKDVqcRWacpH7A/iGRo
serqaIewrKWrXgEOn4ftHKxEdSIZTC4m0xxJSHNP9gub6784s+iNikX2BxjES8bb
OeYAJepz9WGkCFqJxZKY9e1G/vzqt9nMoW2osEll1V0hjrMQFm7h+0nuobuq71yj
1JzoX79trot8ukLT4PF3F7vUYC/5XPDeMbtO7ZxlireU3IwDOUtEkAShtphZrrWa
i0U14/fp6aUXUSHt1pnC05RuUWSjKpC6fyNth4K0ZXVNvVxv/XLMBW/PWpzOgHHU
vNzu5dFqvqLRRlzU5UN+nl5zwg61x0jOIgM3LFhOdfdausOS8wjkjiA6xl4KbgTg
R2J+EpPxshNgQI3W9cCndgPGEDpDkk0OwK3lVL9nLsscoj64aovUx82HoxS6vuIF
DMDZIbZiD9bV3m9S95vjPI+Hil0pZXnnJgUlC2g6RGgS4GQcyZWCLYoGAp8vDs6O
EQKOlNC3WA1uIS2+GxeoMkLkqqbMQZJvgIvYrS6k1KwX3ON/29i2zhkdfEH+tzKK
Hxwc+LPnGU15FngfCPz21D4ndDqVcXF9mXPAA0MzmsNVEJFX8HkJ+4yWmT5cOiPg
YT+qnBlSBwNxhZYOFtMtI/Jbg/bcoe969zhasYiLE7JOeUTFlt+n7RGfFLoUvfk0
Cj+RmAhveMfZC35GW/cLd1yOADivUekgciurdYLf5P8wZ8V0++vQyrhr7fcdE0Rh
rIj+oYpk2GTdMo1NSgad/9qN/Yla9ogBSpNkgg6Gl1CDS+PvgYRhSEtjVKBlBviv
lJDDuDRwGfi0G5hOxbxUIHd9tbUoevWx04WkL2qhMJiTrSJohQNuekiju36aJZys
54ocr4PRZMf46ujl4r74XagEVr/qwQCOEsIcUBQ0dZBhQBPQfOOzvRYUWtSmt8Ev
HreltYIjXNNIeNc16vzeLEiwbuXsVMUycuSTHO/Z+tezipbjeLpMgKe3a85A/RmQ
lyAr7F2IHlvctLeipzbBVbf+XJVJuF5qMVkEs4cfAQ5SSxFT+OJ7AqiM6cRadja3
AgBe1eJtQp6K0XxN7nECRV7x+VridxkGREb6wehp+4rMnI8eXElUU4xetIUlHpof
Lda5Yl6WHtXh+s5HIQlMmhQ6Uf51DCfGDd/+3u52tL6RFZjsc8Nb9FvZ0AwX0px5
b/XnZa2x1iapTBelWgd0j1XiDK+D68HOR+bf/Y+SWw5kjALJqxtVoJof2ShHlerg
rBkoHOT47p5UiW+8NwzOfD+SIsGGdbkr8cUAmx0pv932+Pu5H7M7aNLGVihvg+vZ
PbpmCi86m0rnVf3vrAmFbaFbfBUHuE9UZqGkrb23GAwnAlqr8jrhXJC9dzawPEFv
xPnk6jf4zz1bX4hoxd6+ep7QT6tcRKrbaLSzfMef1WHjsSlkTRk8VKaulqJ+MqIO
q547tLH/JgCH8mutUcGuaj9F4s2AX0gORV6epRnB75hmzca7rUzpfeFe5RivckbD
LNs+3S/5YcROBpZ4XKY/pfRGoT4SeuAGpwdd1hDS+XJyO6gUaZf1MKYNJTDj/Olb
VbmBKgfHkzLNwa852Y55tIvYMUDv0eCYSeChWJvzdcuuDE0CePIpSQ7YQIDr+m7b
Ao+/WuSJbjXlWf3AD8wcCttN5T4gWyIW98gCEWCbWfWPPY2+mv5G1/0LyzMoYZGx
R+/E7+hZXHBFpuFfksJBMLNRlQ+/DxQSCh1Yur2tVfczfkZfXUTk0iy2R0UWAqQU
WtmQrzFsdJvdFTYG5eyGwQF3Wt8duHMw0aNe9qfAx/UDvVfdNvQqrMEA447OK8iA
WDTCikxl8UCJcEN6rfMw3/BEQsYvMBDNB/gzx3aYaf1POxJfE6uyIL0Jh+2ZYJig
1h3oaVxAVyUnAF0CtVnkVnlte7rPF6bxiVLGlD3yJo5b6lxeT4od/EHTCpR83z8o
6O5q5gNWKLyRIcTyED/kKgFKShDHX8sFlLXuBNfER+2y+HdFYJm3qyzKl8B7omJ8
BdhxGGPfXaM1tMfT3WqdbvcDnhqn0VJg4mLsoKtvNSMcAlCVLmB+/cwKUabV3VcP
i3HMTbsk7kCqwQV+2OjS2YjoNrOi9j690wE8bMoiq4eSPiO0EctFnFXKVdwk576L
qHukTHQ2DywnTVUwpsPkVH1JLNcejy1vHcFBvYpVH31w+drMztXXssDv03VAno24
7wJCrWMZoDbQ5BOO/NyNmOGyJQscli/z/JDHda754D3SdREMSL+d67IzwzT3tDol
Iqpkb+kbNd7KCuuB+I3RBwm+U1rmieQmEVcaDJVbdPGzeHQkc2UCb30RP9qpvK/0
fYGfpmfbUVdwf+DevnatRaYLiqDS/2bppQyHJcgBjIKxJ2q9det/Ud4nopBJfO/E
VWGCNvA+ZdkVHPC5zYn1x/3QnF3T7uxdC45z6DOYdwjJFmCXkjJUunrw+DSf8Btg
BgPoVpxXX0uTIQqPGWzgLYHDUyIfpUCMa4cqKMaoPhdiDuWQIEm3kLaL375darFS
vdE2fT2FZTPX63BeXZzKog75R3l00kxxmuCLUtEre9hXE+q7D7jJgV9JgC41Pujv
r1z7bWqd/ee1AjuNCLhNQFY7+rb/+lKjWwWpfbzsfwvzcj+xZ6je5nwQouo5p4ro
IzBYBPBWcZrU1fslsUIy+W9WYFIvfKYm8rejM8cW0liucRu6IwB5Vpj+k5KjTm++
b/m07cvkrBiZxp4Uq2+5BDCR9mifGKPQ1UcLyRaF7sY2r2F3Mp5HRjUqxOpKQGFi
kZi/g9alsS0HleiK3qwauLztNN1lND+41DaYnuZ0by+muci5G9n/uazUyXhzdyV7
75ZSmvtljnqENy0Ot/GyFWvcHVno/WODBucygY0g3qw5egqiDamPrztw5FgKgy3x
zhX4/kzYJtaoiFPKTtWGmgITNdbYHykA//U4iIKAAFuhI5S+QZmWVt0CvObSSuMs
rqmYaQ/S/feuo9B4OwAu1VqUL2L6Z95a1c+sB2yhrViER2TckskNwNCDQYQVWm2I
R9kxYhW2OlKaTM+SSq/d5ajRolofUn7fTXcSQ47NNYNksRbTYySjeb1/eR5up+Fe
Xrlr3b4ve4LPyxv90ZWJHckvPOhjf8+WNBduwRwhD+jFTayKGnDe/AkO2hce/j6a
lIn3gJJKq35lIZqFKEQeSZVpxHZJkT7PzA8uFYfgqB1UJcT73vXhq+rXMEynOazY
KoU6bEcFF5ieJCKao3iIKYhLdQTTSTnsr1/1IIcQUtT0GVM1aLJWjPdS2XEJJFvr
1i+uF4y9gFoNMLtk63hf+wNGkgSmNEwasixSdPksNwzipBTCQ9PkBfjLkfnSMT6Y
pAEU6+CdAxXCoMHKbvcDehVw8npfCC6sKrzNeijDRVnwJx1FXsIZvBv17gVX8Bp3
lM+cvVFxFEZLvEm4ICrmlesIJdsV9QJfUk5TOGMqfLvojefZmjpGewNLfAysibeh
c3qgMSasIJW/MV0L2GTLJImxjGmuNXtIOOYChJHF6+hHps0VCYP3+eKjgaIAB/1R
1wUje+sr5PR8uqem/aLBBBFD1QNA6J30b4ZjyvwSHZ2G7wjdRPpwPzwt5dP+v1/V
mf6GSaMKGEqlG+pKCfe4H72zbM4pp97JBhIkeKn/McotJMAbHx+itTkFBEzCxo+P
+ysLC8ZApEC3cQCBErhXPYrooC1qQ//57nRXdUWvldP5z9dBpepuwX2D3K5jTS1n
pSzzjhDOldOmutgmo+bbxlJaSs0Y01CEyzaktP0/wjwoPhFgarLp6LbOeJr1hdG6
vDeu20OCEpXTUIJ0vk2O8TZbyXZa3HkAJUtk73LlPjpgeYqWDBHlqyYCrPlDtSpc
we6dyNoei6ayYv16Tvf821UdhMPag+xt3RJa13/pFFoiMZX4q0jpTn5/2MLyquF/
pJuiIftrClMvov73FBNm70YMMHzv/f66r6DYeujtdnLxqjfk88cf4S1dlY24TSr5
PZuyfS40pLQ9xZ43HrrP+9qygi+iwm4O4CtESmcxZoAU8AtqrjWDrV7h8Grdr1G7
dxFcqe5AMEmxszKMEz/AtYGT5XJAcsolWX1p1SVVJtTkJ3fFnkrBqvxVbDleilkZ
7PKdkO79IqZhgLDnBfgGe20EEyYT7d/XpQzz63HRpeDDnRvKHn3UCa8qFDQM6Kto
aA166YLIBq9Jn4qhJnQ29vi9EtVCnk/iGGtIF4MSfZSFlTrBJxbA+jsZYQPbmA48
d5b/ojXOw0K4SOV4XUlHdFa4rT3OMnMAm6utK08lv6q2CGoBwkKVP4yPHSpVvH2l
HCckz0qpJxZt+GsXq4nFbTl2vW4DHY32ulGW3beQ9ptL3RLfdwvX0BpV2Rt9q60Q
I8gxOGGphv8hdsi5N4T4RnEmluETTDoMFGZL1oMWe/GD7nLLtBfOk/0dL5k7mAav
fgDntKNC7B/um0D0ZLaPVHYHBgVfObvV+cSYFzcuKeLZCepM9aKphKjc+vTZQcdE
azPX4NBXM89RLZwHzgGPa+NtJSXaV7ckijYpg2ght1DmaFOjaUf7edYjESzfqtXn
rCQi9uoRVkDsdsLC4cxbpPPsWBU6OdORIPqJ2krh2++4YRR59kb6aLOaCeU2j9FD
ewXq7tWUF7AxIgUzAaKOX7XFrY679NXQ7HvSM1oqso9jsvFohmdXFpYOFda4tswU
Jbfz0vzMGKECro289s1RJw4cWHiYt1aKTEH7eqJYurQNP9ik/IxULFY2XacdQRaG
GNyeWjzxNi9tf0WxOJWS9PoHG262N6GpncfYQ02306tLgbfnlbNI7S/zWDR7uPLZ
vRJoxqLlmZX6cLFZ2rhz6X6q9ttUDbOVMrk3LcPhSKfoKN4Sg2jWWdTmIJb98zsc
1G+I2+EDShCjnzrM7W6gTwFTSmcawJn9kFu03fb22QJ4InCdLrVLRAi9qLvMVrwV
Axk5YP1GFKvoL9bU1Qv59fKT3lCAOUTnJyabwB2hNxi4gIS4d7tZUI7yA1AIN059
cvdo/QT710X6JvGe3f5+NsCfl1cuKjikgQ/UqS8cqqyzrS7ODJpddwmBfq8D15Q3
1NstCpQP/DPAFpfXVxtmAKtOjhqCqgmWot8RXVmYUT0xXrN/QgXJQL+W8tmK/oDn
ly52mk/hHtGIq5LDfcnsxdPYWpNmTTYsAM95mqOhHy93RkKJB3sxU2Z00naJQ0gs
/E+NllMjeVy1vadWafvot8uB0cl+8gxM0sHQg18aekIcC1SQnHMndiYTEiigxw7E
jvoFWJ/fb7V+d2QawTcgvJvngw3x4KKDrMcmahIGMEXzwJJP+BvBsRW8TrUWPX6g
wW6W1+veMG5S8Pbd+42KlJcE5VZAiIDzudOT+d7M1uflnZeP2lr35F3WA4GovNUt
PbLJ0FLuONRQ9vO4nmgTZ8Pa2Uq3Q70VscaRsphjy6x2VGqUDJc8gc+M8kcPEOf7
Xne9AZ+eQgOlVHyPSOsfW6AaVSKW0x8mqEBfuTJym15+oQ7W/ZWEcouEJLBw+JWm
s1COcJEaj2JUslS7NZTzuJ39OMqhH+7InLAt+hVfM9TVZPWpBsPg0nYKjPn2M9Wb
xpQ4ObEU+0ViM3cw1WrXAcctxuD21ztUfPiHPX9wPI+RUP7EWG+77Zf22aHmaZIK
5EjKlbvxqBvTmftAK02TQOJHgYS5PNZVJkQ8z/78zJSh6Y1ndBtIdyaMkVG/ijkJ
zMze8zkwsZmkpPxNfEDcvotkZNv3epyCtUmIDDZq96JEdTINEyEZbbR2u1HdOKIx
/k+cv7vjlxXT+ZTtjh9EXvqfgTYDlC6bvPwHk4Z46VNwHJbgTZdX39KMwMACzEvV
ACwkiAe1oaE1eEgfQF1/2vB6kSA+jLShEwiBGkbU03Y4Zuz8VLyCeq49szSdorX4
pezFS+VQ4xaADU9bc9CL2pQGMO9VOZRmscGj/aB2JCP9v8fO6PiK2zRCVihMshAX
GiywMTDUqBT6UEPRv6f17R2o0eaf3HKFhTkncdgepQZy41pEdn5s9Ys25Yns3+2C
r2GNdtey3RrBIzEUfNJh9gdskB6lA/HHOtzZDmJGJ233O52y9bACI0LAaidHcH2r
r+fyR4BlSJuVHRwAy7uJ79c0vvqfbrZT9dunLPTt7EHt60IF+N6LY4wtqN9Djhet
801IM7NbRu9iwXLn0riHDsi6LSRa7NYAnYTRLuQFaPcz1JwnRzp8yOvZ/W/A13Jv
4FVjMbBG1UlcKNakz1WBfMlGQw7G7zdCBCcLAguWRDhcAc3WZh0PH24jb6n0SHX+
IUMriGedLy45h5MwPe/RWHOfRxIWPNms1PYQreNF38Sf6173jg20FqFLjJ9HgYzj
6x8UwRdaeCg0Z9qkuuogqkdOEa6JsY5QencdCUpE+HPKl0E7yzfG7cf2h/L7EFKR
GunZARZnDxJQo1EvM7VBE/tO/3Sz8P4L6DvvcifFQV2KgRC80/gWqrGujtG5dSof
pHUbPQR+6KnVgqaOglV731CN7wgz4nx2LK69UUEh7trd8YXSf99saLB3tkE0FvhC
t8lvW6aUwxqmlSCNuS8LbhiKIX4xJFy4ng4N+dxw56XjRbvFbVDyBI2UAqizjdW0
gRuSIQRz9lb9nuB837cPnKq1pXg4AQU7lpG3YawIiexgqxyU1GdVCNi21D6q9UYt
77TcUR+32TvaE1A8ASQnFSIGFppFU/Vmov5H7QubUJY/rCjXe30iF3JPVERGUL3b
PBmXwjD8f8tXuQKgDCelwBFzrRVJFloqbD1eci+lNYLxWypdpnvtFBRYsdt9HF4/
X6bSfiNudbaTg3CfWpJQ6XKZhIyX6jmsWKYqUg1jfMrxJhP2Y/J7eShIPygnnvGv
WrRcfgPOoknsJA1XGMmV3z23Uh0zC0tKqxsD+jGmcxFvUQgplLIXPNqxmxivH1cQ
C0DHt22IXzdUkm2RukxWYUKF2E+AppcqtCKwCPzNy+nN7Bgnqfg786JEMSJb98IG
mZ4eUn2rreOW4SuTb6UGzUGZuLGzeV5TEEZz3GMT4jWHUvHn19V7qZIDfh19JtwL
2Q/yZPs0ogK3+J68h0zPtEjJLY9ME82M8Bvlo0IAXQEt5RSpmT1a/kHwc3P+jrjU
JpdBLOYuqNdINkkb3F36iAhptDW0S8TrccpXVQBAIo0zuwp6G/UD2hqDFb338dx8
ho5kTlPjCj/dvU6VntSh0q7vqlr6eSneXpmS+gZuYErXxzWH4fHrnWxluU6jLqOX
68SFXzC7bB9ykS+G5c8W5HfoLhvBkk+XOMOd7xPhz5VZ0ZCePTMKkgDGxnAkf4Kd
6xFCexrEnGdwYj+EMYElDMYb1mNz1fazFLGVZPzHvPBmZ9T0T0YNZrcI9TWOsTyd
KDa/qJ6JMhOW/2DcI7qyUnJ0OSJQxq/i4JiAajVGjPnlSQzscfoPRJjkX071NHwj
HE68SJi8R9eUEQRQzjgVMxzchSHANt89SMKvDSWVEWsYcxa3A63AVVaZaIBNGDQ1
Nj2W4Phzrs5NxZwgEMhnvodzmlBTeLNtp4+jhgo12Ps8z/vnz9kadb0De9BVOYsb
8mUiLaVTq5O7YGiR8xZhOwTMhgIZBNmjyRAyDjZXJY+haX+8mgukW/yHcttYSF/q
ikw2No1ujNKVmrYtVyGItZajnZ0CQ7wKn+MsiT/bWrJr0VG050c+VPp3qfIpCH/e
LD5l2BGgEyZlzaftDw1BH0TF+fntH3yMLmFGS4gSsq3DPD0NfcnI1yN50LW7BmjS
JPR+0+Td+6CQzusDP7GSgf4m6hkL0/2oRQBJQVS510srdqNyEWs2Pz/CdofllxvZ
gPi5tGG18UUFyV/uz4Ezbiyhh2EfchHtJQ2f29d/hWEv43WlZ51wMoNf/ZlpY1gU
zVRG+aAvrBGuLLOPAozUua6Mxp+CMMsT3U0VpaumYXWqYcJLYeoxvF8R9tJn6BP/
yNkksuQB7qxhTCxxM7tx/PUGg8SVK703rzk4g9FZtWN0Oe7mceLZ3QOMdVLmz0i1
e3Sy3baZMd+1ty2QcVe9DXqcloO5VLpLWIsa5yGmbRZ23IMFYSIgWyVFT1IU1SPf
SuHmO918gVkfg1ioiZO3s2tmA9/w6V5Yw/IaVMqZTrtsfb48cw9KZAWc8yZ4zO5L
zKydjtyZ6Ump+5mKWPSFRw0VZ1QpbzPfVtMuRRAdQXq9v6f0DJsJvIMsIHZJ6//s
zbY+fdM1N0/P6DJ1M8HpgI/O4whK85aRSUbLOogjUcfBqUbKUwKMTOob+906cJyQ
JHCrPUtvRGSKzrl1YUqx75th8lsJQ3dN1DR2oMug/3372O9GmtiDmDw+GE3dEfXu
Njy54GncWDSLWle4tcx8wNYlTS7DdIhLqBK/txOW/qKwxH0SMHOm3Qe5TAyi+aFE
bX9PfuOAVDg5kq+Lr0OlRZNt/qs7leli11drldyLL9iMqC3UTPvLsRJWekQ6flNb
zdZhibpyNJOoldTJBXnin/1bvK+NA5CECJibtOCJ93K9NbviTlvQX9Ef4bVc2l6u
zm1SJFyabR38rmhs1uoyI/NFnnOeigvAX1SkSoILQjFYmCd0C4nc/8geD6hKp6+S
rogiyNuLnQ4PYwMB3MsMqiYUD8zaGPnJesGMB+trxOGGrejJm8VGitRAjumxmL5L
JRdPgxJMNlN9lQLDRICDGDsCnHpDpIUXWv711380cpTjlEDHcIBio/fY9u6/mq4G
T5ReZ/qNPYSSXntHeWGEJfpyXCcEOAr7DFzf3cjlQPgl1ZsHS3PAg6aC10nunWtk
/uKr5+t2fkLwjJVQ48U23mWndKSFgI4WWNr+PhuPVPVH3iO7lytfm1Mph/cbRjoK
OjWhnQt4B8Hiupd+85cUtLz3aDmYbfoEuSU0idXAUWYbooMLqApEY+6tuo31wRei
wzUxHJv259krt0TVIe/XFQ2aDZLIbrb0xMBB32cgUbUbDhp8vxXWvRvC2gt3SbjA
wUEO144pmqC1G7Sd9wgQEUxyi3iMlI/nuGBMi55hVr3QXpHyXM6zOX5J8Scru0YZ
e/2fvVLI+0GPuzyI5am33q6J9d2MRstJo7IKrfQhP/qnyzMaaFu6rkhlh9Zh2CZd
GqjA5iGWoFlHZlCUAy4nJbc7OQMnpdW37L9hE3Nx4fiL1LAwxzSZEkuDo+W85WLs
vuzqkCtOP8lH9MrGbUOu5vqrCkxvWSMlUX6I2XHefyR9uvuhX02D/NBUoISxSpN/
zAaOn7rFU1lu2X9Zb6M0EJNaT6EsHDP29Cq8T9dEMJ1YFzQaTjvSNTzA4KaIAqwb
ZKWmrlHluZXO3X2Z2QazaRlL6tb361EMmwdWoTc4nmo4DOavTl6vvx1oR0uLkVEK
43J+FJ4RgBmseIV+zrqqE012bqAVOY52wevFs9WjDYA9GfqclA1r2sO03jDnkSfh
wi3Xakv3Z1ULTNTMKVTeXixc7G+jPpTn2BvKg/e6i0XYwP/a1m76DS4bDg8dPZ7p
JHL5Ix1fH8XJtE8DL4gpzBTO14HSFmbgwybQ6N//d1K6FqjbtfWKtPjsE/seWUx/
Uqf2KS0qJNWlqoYqBtDMvToIT8hoKQJ8a50xYLBFV+WYqUXR4Ca4bHZycZYAtYLf
s13rOXXTlz+0yk9nKaM1IzDvEsAO6th9JL+pNPcHo8RsUNkkdDzSjIPZaDVQcl+v
EpHqgwdvEsPYiePC4De5wEoyrtFzboKf/pygX7pPc1Fbr3Hz1smZ7hZIaXC6203d
kNWnmoJmIM0qa+ecyaKAFIjPv9MyoGNcZmQsYRCwInyd2OygXLSl/8OTWJk9D6zl
2dM4OiE/H34v6JevwqbLvHyeAZWp6nSW9rIPCyQdase/gZ1VSbvwvf/VupERppZe
ToKce5a+alv+KsOelVyniFN5eUVGto5Qqk82RHThLcYK+E5mVkpxlqvkMzGwb9+U
ns9NULqDeI6Ny/47In9uevoSLK4Hfd/XAGTYNpkl4z4vJa9BDKhcJYYQ2Qn00JYd
5RZ4UynKib+APuw4Zwaf7Wjrik2vn0XiueFe+5LPj90dv7ZprWI4Ij5P3ohwvOSd
ULkABfr+aW95Z4Ch7388i0hB+lCKuwHdSLxHrM/PgBBVHQCXrjuvzAID4HXN5ySb
5F4gHztMHMJzYmvUrUYIVHbSL/qqccMeb8Xx9hgB/gYLEFLX7XqSwFfmqc/795OV
qijNOtQG99Xf+4LvybvaZSlmd1ab54Q4Atwye/FS4WgMTFzMkA1MA+tbU7ifbkzV
iV9FdQ+oORu11nULN1JDioVRLI1PEJ37/meiq/o6XtDohkYva2t/QYCKjjIIimfz
Ac9RlyDQbMItynmvHenbThRlVwb3osNjbexh6Ow7pny+M/TZ55Cwd5yiUKZNk5b1
HnjgBqnviox6QwiHLPQ7r8fKcVDZSlJ6ku7yXCFy61U0JMyBEPrMZzpvg0jWU1Uf
ozT8o5tz9nyvmBd58qPPc/DPGUgwhfXNGV0pxGvttkdoT1ipmPFXngcqWlwtiYQK
KpPB110awdUYtN53oenH2f3ygSzX+CwCYzB30yVL2XVVPGJxxPW+AdhkAbDgRHH2
zf5q2GjSbUwiyEsYh3+voLGL4CyZA4zPk1MhphEc+RuxrQW4FcWf5WLN4EAy1fcc
/OBuG2rHCHjwccKjWxlAOzsGoW2GpC+ALpgxubrD5vEHr7/ZOj86cktPpEkp0WPI
6HCJI8jrBNpdHA69BQcf6cNXtlsNGRWxLi6CV3drjvxj2TBavJtoDpjZ6E00JEd1
p0qLBueK+jU7B+fShkIF1Qvk9/LuHU4Jz0F2wu7cidxZZ+SQ4+5W/YnjrAcwI5bH
DZHF1/WQAmISZSIECLUaNelhjkWFFcUE9g1gzUVUsmkQ631j4V1qAbuKIcowIC4m
qJi4GkyCInOuuYTgHEapq+OHrvkPArjUbF9JzcctAyQ9S1Jhc+wG+QhUuu3dYLFO
ZL78XhQBpXizO3GW1G1YmZXVJ/sPqVsQoXCH0N2LeYlDjllJUCR7LnQxungcuewX
v9W1wWp3sjyFZ2oDTj0FRURRrPvTvs6ngDysZkUEXjmobhYAywMuheuR/tpXYTA5
5vx/fss10M7j2ODvIVHFOabHv+vE+NFyxGBm6aUBmsVpAiwiFay5QovbPwjIhp/+
i/bygly0Hoxyh2lEUtnjMG2HZaOQ3Ks7jgHOBZSxY9aT6Qi606+76DfpCbpfRLLZ
QB0x3P5N4OCoDsDvhOvITUX18nCZg2FGjZOO43Bja4jS62zgan9wLTwBYjefZnKM
NSGqTzWMGoUUv9Pg/xWEYUBnwn9GTYBNnW5vmQ8GHRaWFweGAJOSe9+SjoCPHFfg
CtIiuJuLfXmIfItj6VCgWA8oTEhOb/oXkyVBtcygZg7ik66oeDEl3eCvbveAMqb6
LzN/wzT3TFwBLEzduPVV0AhR1khvVbJIARrHR31ii2JNiM7aDNtc5++ILX64EroF
rT3rg1sEgqMEO+B7MAEDQIdp+vH23u8CHkYzCHDEFxn5fykeL0SAy+oxZiWVOXiS
ad0YObhXv68PMj9+Bi2V7Gc///92xOCSpl+pAxsQj0y0u9/3ipIf05BydcguJ27Q
jrVlWSPcF7gBLtGThSEGCRDDs34NZNw4/2Y/owdNbf5YHFEvboj6aSx2yUk3+25a
lXF0hLacfws/LYPAHaZX2owUAb8CJm1R8Ta32dGvtQwPJCOdQNXzCBI2uux3k67T
DlfkjCTzn76dM5i7Rx3ikD513MsyOYy69NgOMSkjP7WQWg/eLlcP+UB8LAl08aa2
WsDdK+bnnj8HCa/yjozniJUwFJOnicqNEC6KN7h6wHlVnYbnc4O5S9dZD9FXHGqK
lujWrR/ZIYydOWM7UCbcnp2MqDFWjpAkkOSuu0pMRZGWTjR2MgnJYK6Bno1ADrJv
QDqWywkx8k7CF6FlhHu+BxTtumdAvo/lLpTzJXK9Dj821UDdlHWFFOc4zqpxdLTg
B6G4fDFZMcEsl2nowtqF5aaEC9n30DSKu7n9UJqLMaKEfbazqcsLbGErUKJPbIj0
yWdVKDoJ9KYRf6VshtOPWXEEhBTW/oDBnN2n2bmggeXaTdWFFG+kQeaEyj5NLVU8
Hp70tw/pZjXfWsKPilaZ4JcHRgmcLlheRCaFkWhqcQh+yB1YLMCHqSsH8BvcmQ24
Ni6QSVC9SSs6iCqUg9VaSPn0W7yCgojJEdR9+mxxaWKTF8iFP34ByqTOL+fH6Vwq
OabKvYnuEriua/7HDQ2yfjL6STZkPBO7krjC31xBQLKj1Q+RQUfHBPSjXwXoxhZG
acIBa/dydTkjIVCAOBd6/S5mP3KmRKYCzMw/YAP2TfB4GMLXBiPnI6KAHqKX7iOl
Zn9Xd3PMLcKx4eukMaBuDETZfULlYSuP9CNZu5lv3j2QKjcD/Ov11t8ry/tiIXmb
Wo1PRRUtGv0oXhNEgJdNM21Fo87ZQ5DMPDHf97MyObCTrP1beAu2Rj2YpkT30teD
TlAowL++4esfABv3VgNL9miC8LT0jyb9Mow/fR4h37lWHLtzApNBBAO9WgXjw8u1
WH1wDoYxC+rLLo7BZmID9wlkSp8T92Ylu2TzjVmpRqNOryK9q08KaaeFj+fiNcWp
ZAXkWZuhzfrxhp53FD2VqhvMsevRqBLDGTSfZaOsCHKIgxhTYzQ3LI4M/DFVNZhW
dWf5FtdifVqNqq0ghYU27nbYC5hX3vso6iqX3GE6WL+8LyxaaI/n6H+IKJrTlavn
KxNEOClGrgEAToqk7oqLBjWv6yO+OSTA13yMXhHS1yiioCP2g8HrA5P6UJI9nHYk
6yt2B5PolspKyQfAvi1ymlP28nfQYAKlcHzYRH9FEZYsPUM2WzivEr6cMZtzTdEZ
i6f08POenBTjER2ItRrxbN2EgF2b7knrKQJgl4XMjAmHpTc2VMEavEg+N4IQu+1+
rdD4TuqRcak0y6QuXShlYEtMctjFaNDFXCsmuMEbtp+nDTBn1hXDgjJlYTAt0ovJ
wetS8GEGfiQhPbTSIxpaOazupzI4PrR+gpR4MV4mIeP2CSY3Qj6RNt2IOj5xkWJ9
xorcoDcBUgrn4/ViUvo3uFyLwo6BnHmy2Ji9fPXR/PPeGV78du0Ssu+6HjxbkcRW
WMfFcK6DiWEzIImmIOKXU4h0pOWf7a0AbtG95pSlMHaDBqcLHNl7nMsQnBJPxti5
pshH8k3Na1j3tX43g4BZlvxKnN3vaxcQ+osalsCg7OO1p5D22pmMET3bY9kj/EPf
6OLYdhvca/Q3QlW+TLxZh6XORmhUxdbPj3ALC7TzlIYL60zkx0FC7q1mqbfgbNAr
nbK1Wfkf8uudVMG+wOQO9de11anx/f3FZAgkBGb7Bt9aH9acFS3mXr4Y65wBVR/1
Tx1faSmeCxYXPRc66a8HfGiXOu0yRfuyYe+51a6dmEc2QFujYLkWIb38rLYu7Nyy
bX7PYpslRqN1Kvut4Tnt0jHrLS/GwjZf5/9rTnTppTjUOU+q83GXyO2/GE3ix3e1
OEcXvJsXIsY1/zvPqVUDyA6LA7tU8C5NzFtg6JZ5IqJ6oaDz++umUPk6bX/0l8BG
vOXsZHWrcOeIgJ/SW9vzYcgRdNucmhGTe+2W1XlTW39D+lZIdxbX8Gqp9U2/NOxE
52gJEaVAc+hCKBJT6yFeLUcgknpQwRVGHMKGCvhgiF4ajY+Fx7YguGE185MFiSKm
XWvxwwabxByABZeeZrb4wCTfs5pd+Yv2dbRyRe7aZ6mQBdVMoYcjv6n389jVgg20
bB1AXlHXPAEUJXCjLCnzDAflufj5kM14Jh/03/T6aGZ3L85Fpk56uJE8NURlBkr0
rAxjwmr4U+GCRgcbZWRFNxFGcupaUDmLFKscuFoMLw93HXdwY23jHzA6Uh+XRji0
C6tQzggNeZXv6ldMBv0PNQ80+0kTsmZiZFbrsdDNL5PZ9sVU7ihOZPm5RwJrvqu5
Q+hRsfHW5WTtAXl7bpZMD6jwNydWa58/YRLDzxTUQxQdV+ox4Wj7L4Y9TCtD6AXu
RsG/Gar2ct7kgHX1MPEFKJHLRC8au7pCQnJMfRKsfwMuIGg0XYsbjv70Z2pm+8WT
zVxapUEhQTIknVmFt2OXfNM+FXwMsFXMZnoFEkW8/SH3mu+SjchB02wZzUF2Wvct
JUor4NLdHP+PrVU3/xmuZl/upoWFtBn8tXrs8BBW9f91FuytZCgzc3FZ0tj9pQRK
48f2krMjiO/9rb3jtlzGdnsZ4PlV0OW5flqhSVDNKaj5+jgXG35c0gIvzqxwXCmh
CzP/+JXOTs6Oan6+V6BUJMZ5r9CXWcwL0BoFEcsIOQzO5fbXWFH4kOzhP2gjPrrU
3nsfvNmkTjOzNLyW67Oiy8zYGSGrXCNBc6VShUv1MNGnJqFhUaLRnwmH9P+rsBU9
luUdLFJeTn6IZFFoua8n7eWOKRJestkdYUA58s/npngM4pf3uEqvoZS/R0BqwRBs
7hS8okRcMhllNz1guHHp1XmiibFC2/83yJWuRFFpc9yCZqFwbUA4/gggD+xWlFNv
lS5LYxH0O/GvhCBL8wpFetRDIraPN+3YJtKC9Vn9GhgzBHTVLmCIIb3H+BcWAse8
FAWg7EdLTtcx7488beSRtmDvzD6IdEB/XHFz07ttjDq9H+2RsMDk0N3gUBnley55
YImta+GexBQNpvnTcP3w+FkA6ezH5iu0oEzetRS3lT+SOK9sw8iDBrihwzpSN3q4
m/8n1IzvV2NzlonctZllsp1u82TmL8/lQcHSGB5izuV14QYi1ecCX2TnGcLKflGm
hOx46yb3umZi1T9kdkWFNpOXipDxfVRbzfXLe/BVFtE1Fj7HUU7Ak2AEGFdY3QcH
qoScf/pDQkHWb7jCcikSSN7a3uzEYTJSV+F90P3PCpUG/XbqDAY4PN5e5EBssjwp
EGuEwd2l9199z0ZPDk+TsF1Oioj6lzJYfSGjkceL6JxGNVszS2ahUSyDQriNAbBw
mcW6fqh8wVQ+RQaSlxjTPBcQt3BKWRoV2T4I5kxGh5w0tDTYoVdQvqxcPYCibs25
MXYjkqs98HwEraeRCjyU+J8il6S+gwaPk8wqxlt5gAZ4juzFJtiZS5dTUcO4bKmt
qiFzy8VORHcHdSKRB/XwYTEEidvx/qCefEfsAWUD5DIYU9Joa/0EZJfRTPZSAe18
o0B1Ua2WfM/nBcIs39aboEdop8pf8dCchDIZcnwocHkmFa9tijaQqs1FSNVGmLt5
Rub1QYQAyCJgPl2GSfc+3/i4s8RBUccGPU/H7mOVFnUdMAc8GqpmG66DfHURWuQn
iZ3gh7mhwN4mBeziKY6HVYhinVRzZShkGI0/JE11lUyCnVPY0+lCDafjMAmMP6vj
9vbEPKN8zBLLkepkQBkI80Dnr82CeiFQlV0Thmuf9IwhELYFWlL7WZM5KQrIZZSz
NwPvHp1l9u6kLrChU9/Z7achd9SN2dFnac2+aJtp8VRnU8IFf7qD0YiQT5UOYsqi
Ip2x2OnuxRJvkCoQRBJLMSl29ogiJhBQhVNPP4f0ZMn5133hrJL/K62D8kMGd+ef
JChYHx840qnWT91NPFohyHk5Oct4dUCZEmpp72tFaBzoqwq6PcoHphLW7DmzKtPj
HAChvq+sL+px5YU6sw8SyrrY4ub0htOG/2MuolD0WvCOnw5BiRmwCx6WMqj2AY/e
3ou990e0ofR9mlCd9cWX+CSNvKgHGMm7l/Eu+yQs3sdOM5Kp2u4A7GwBOTupVwV/
qcHsgv3F09k6Hics52WRVDcZ1LohPSEFCLREqfxNesBkkFu7S0XF5NYP7eOFTkXs
uODqciInEVjqFgQ2Vh677lFxu5pK1kbZ9X0l8bJYIE4IX3taMtDkfgPN1sj0E10J
QmtvLRoF/VZPeqZ0PoWtnfNhN/1UxWnaXw87lLUpMHj3CTcudxDEkE0vYtkqYtXX
WugiR96/d0qo0/SL6Z3SS8rBykkxW8/5a3E/++PKqLe5B0gYLUxspi98cMni4tvM
hC8o3QZdlPxoiIRGI/aCRV0/+IsEINNzPLWHUEDOnqyBn27MGaroFtHbylVYrnZ4
jEh/HAn3nkShB4ZYcNBE5Uz+CS/mz3h97o4i3TtpZshUjznuMzJ0NLXCEv40ypuX
7RXQIxs9VTG2Fw4hgGs4HyUdHpS4C8QrhchuF5MREdKb2wlbgGgOpsEfeKSd3U8M
q4fdA5h5PzSeZBVMwKZ25MdS/VbZWKcqfyQ1Hq2FIAmKCNE41AxhU4amQXrB7DYM
+VQ83ExnxgQaJf4Qauom2AYKNgIH43WmRo5deQleBYE1LoiFACREwtzlzqQ+FxH0
ZWkG1J1aHFx1MqWos5xrFTuByeGx5OjKE2H3DTYXOR5WAb6BwW/FCbsP/a9DXUBZ
d7VrO/KD1Gq9tdT/j0n0MfjhA2SG4x5HVnTUeB9rd2n3bcac0CFuo/lIG0oRYtXc
QhXf3gA/gHT7jVfGMbwmdEeWLicGQJGoSjmPgyY66bbYZCvebdJ7JemWVOYcZjd7
/c7A3rpu19zReT3s2ikrAAAHTA9xJWm+7/q/KDf77kPh85YbwqAMWuvmBk9nQK/G
MW3TTFw6UwDCqrOpKu352y4hcnZ97E/eblVilWeFqJ60azzT//GW+dbKdxdql2f4
THLKpqO9tkzB61qrQUMqOVZPsOab6o6QLXx7Pq/FeMbWaGxPzGHyLD2epSpRzI3P
2EFiuVfE9hOV/cLOyiaBUgEZcyT9sazEgD60pzKlqlKJgqBiz2S8745WcadMU+i/
o/Sf5jFsI6KrL0bnOMGE9bq3qrVJCZV8Xb/oDY739vOyi2w+KF6AE7WiyS2m7xZB
93m0gN/I7q44oS5UxSmEUoKBQsmVfVhvipuiA1DzcoD+eASZlPlF3bIQHltdqPZY
kWJpKJ5U2jN5VkI+AS+x8WgWx1Ai98tTGpoJsnLIxqKlL+Qvr+6LHO45vu9xwnRB
L6gua0E5SjcuQZ0goi47PW57bsivUXpMVktEe2hM3tXS5s0myAB/O5vBGlLqk6sk
lQhGr/JY8JZl2fdYoHBeure9WC9/ZepdCw2W56ezJLOx8anwUaA0NRTPUY+whc1J
SddYkaTdh73lsASKxgiXkwzlKUqBCzNweBLxTmiumhGJWOrZaFbJPGXmB3TvqoDq
imKJ5UZw0bX5vGnmmNhCTwAddFFNeD61dFQ8xl9lyOiao14uDAI9eQ40+aCMRjT7
A4gGVOjzR1GzDXZgqO8WQ2RgUIczRFwu8FEXmpGnqZEob5mAlduaPGxo8FymFS6q
lV7E+yI3YS49q+b71s/5WjtdZLw6zamfOEWAZ54DkX/la5khVHeow0aSYmV1fhP7
/hRfJN3TnApf2v+4nw8JFp7jt7mjqcJv9ETR+oZfimv0Sv+eL1/EZSo72pbmc8kB
ZhUg8oPk1Pra8V/7DBdftWVhPRDdqFyVZDpxxMbOHBVzci5S58sFxV7OUuqElyOS
0Mq5xwfxKIV6yymuu0kIWud9pGEwV3NZ5YSOuXuo6pvK9Qb9RVQF01pnx8YE/m/u
aGZdHlDV4509yH5+83QstXjRT7DLI94RdOSxPaIjzjwOjHl5ytb9uAKrDYWgSDrm
C/cG9WlsOHvpiJY4wZXZuLq8mO2BOm9Zrpsfdxo1sdw7A2F+ExLkseswSPOomvWn
9Cug0o9aCcE3cH4WXwNEzX04Vt65DZFCsh98Atj7UfghXAla+nhx642egbXItP8u
RUfjHs0Rbo5EYhDNQxEPoV19BmbFyPN/CQzQjXOJtUxjbgxx8VH0VwKEdUiY7iv7
IssBDJk7VMK+F2JeEaKA4CV5Bk5kzxyJliZiNBRrILgZMhOdhJJGBSOXRJ1o/cvA
lc45rlfk1XCLJcilGPJBIYdqEeYvIIVFvn8H7DwZ94OGfF7n3f4uIb055wZ7zCSb
S39kHT2mpyuL6pp9g9LjkgzczzxJdI7YbnwKL6prt06G4qDMCt4tARSP5Eob49DQ
egyb9/lWdCwIjOw1RSKc3Rj6Rqzyld9BLmtgz+g3PVkB1I1Rlp2immE6hLIiHD0C
tWQEXfpHeK5UroF0a8odfcpcYFlHIbfoZpW/0pbwyh5bL60yr6Bv3DlD9DoZJjVh
yKoiWQiqjIdrl67HgKmOhgfCDhdBSuQWeLW7ZZdvVNWZ+5RQe3wgNPtNe91YEFKe
mczsYZHX7GGSxL5TKXVpCBrOy2b1dTmpoBcsdyq+7cMeFFe1KKeVFRX/H1aoq5wO
0vlQOpzGWhjY8V5oxrAW26u77UkpEXWMIRgQpNT64PwD/ggnlaJUq1Rc4sT8f1Lp
2S2/V5hTgpW0nenJzeOyEYC8Z6Liztxg0vknxUhZBlnMeJfhxORtIVqTUNDEYK58
QL6HjLyugMFs0t2OroiHC1Tf/mzDXexUHWD42V7NQkPh0/84Pbq+p+pV0T78clOt
20Tupns+kvIysHLVVON1A+9YeLNJLInGxwK6s+KygNYAKV1T1efE5RKH2rnmKSYy
2SSXruanTRNuaKuq9vO63r9fyqUAEFgsECyblXKKIslsX1Lqn3uD0Ak4a5Z0m4mZ
EMvLNbLE6SL2JWAFv2EnBO+7kvbZdq8RDy2cWxymqhVZllIIEYcfo3vs3/z4CaCA
IvPeEU+Exb407Qy42IR26AweWo4ZKNFPNcy+VjyFzy7TnDUkr0JmVYyZ3l/A98mQ
Skvjkj7bb7tzuD0bLysEMEcXqtYJJqbhdtW3tXyW3aAHdP58QE/vCWCqJimkPWgM
ZU64+d5iJ0qYHEbKxAAJPHCnPeW2zxkIJZ7mUWRY9nIt/eeMoLnyB0OyWxXV3aAB
BvNZhtshmlWijn8z0dPa0GYiyd7u071V85usombu4Lyut5S4eXi/NODqpK7yvEoW
s9pidGA9dE9DieE7TuDHshbF5Tq7+SuLMZrCdYJhKMm3RooOBZkFd5W98v5fVRXr
iAdqfg7fq7flj3puhNoLQ8Dn8pDbt7DCpXwyPeU5L0+S/4ijWm7vuXJ1o69F7OXQ
9YAffGep/fqrbc0D54hsKDDc0BDgSu2ANYNABvRf5fv1kWi4iaN0P+HyeWgvY/A3
bu+WphtpZb6qlq40dCzAoszY2z3e5rJmtj9y8g8zYHZN66PDUSwWJdqaF/z/fPpW
oaqSn+D/Dk2ss6nwmAPYRLqCxCw9pHxzUAYQ4eaRfobeEZJsmN4GnaNjK0KE8704
+N2kXosuMcTUv7a0eSsdFqFY7Ib1FyskrPRnB4pfzixQixnmKJq2aYytSH8F1GNe
NNzs4QwISGjckzdpodxlAJ/DKMBr8bwEO8EepvZfeOR6ozU0nQwpppy7hVC/hjJ6
BNsiD/NVHSIX4zkjnjIZ0Tuou4JDC7GA97OeF5j6mJg2M4pRq3q/72pR8g386RNG
HVsyDnUDZO6Qp+19u4BFnAxnviTvB1qMkn6+7JCUufsEShr9MY623JI7Chy/hgbZ
gsv56hiYrVuZWBpFO6bvx0SB7NoLOxSOqhmklaLWCNFSu+TixnNe19NVsbBKxJ0L
VLNPGkPFQGrO9KPI1mCHIUIEubTykeQdiRISQfDtoqjzRKYxdmZ5Vq+dSYxiIaDO
HZTG2MMmYCJlBDierHxHKkEI+FIHlPcDxyKD4YaiZlXiKWbRAMfv2zX+IwuR4B6f
w2c83zg0nAJMXEKYwdDGcZFZAiKbfu/qjLgcqZvyIp0CHD1FYPHRd4alRAEUKm0h
2SePR1bsvc3BUYl+goEb3uLGVq1ClN509hxCLWN1I0MH9mff4o3hkNscNjGNYxlp
Svx65loqvKblNWzTqrPUzPixbzdXTYT3MPOCLr1cGS5mTfPooxTqTpJvItHjyTqO
1o/D7Dn8mqoNgkv1NQe3UhHUM7I/euP9mchLpik7dsGV2LyjaI4S4VIlWB6/1MVU
MRvR+hoGVnvFfdZc7rGqHvZilgOS9jhGjrJUIcbrLnJnSMvCfp+DNkZtImnoLfOf
WuW+NcZdDZOCFmwk2iKaiZiF/+m7WNVeWGcHuaihl970ZaOuLIBc07sMjD+Hz7eL
5l1+lJJraG1M/s/Di1w7voIJr7enKBNRxaihGgGrD0MoVdzEIZamayvZobW1sNng
nvtz1k3y+7btsmGl1lgn+q3CcV2/b3RbGVKf1beI4DmrzzFt4igBt0jeFqXT25K+
qbd2DW+EgAFZIa3ewslWTY4YnzvF3r2NW7KGixUTHfTodFxDA4oA5cgmZSh511AK
RQVz7OtHM6DJFr9v7TXWlmKq/rheKoq6m7BFswCHhFve08YlhV+81hcfoV5pFLQw
eGW5giBiCXWHrowiLb8xcagDp18tZ33JmixdrZykp9TSzHfMaB8LWYLoyQSqQ4Sx
OrJegb23kjp++oMLKKTrQTH1/PO3j1jaMt9v+tiu2VYKyXdKabAvkb5mDgJT8Slo
CajYoc+eKJw6pkDr6DRAdzKgWlLWrEXTavYNg+zLRaQ2n0QLkmih0+Q4JPcbqKgX
8YPm21cRrn6Ls8PXmD1/w/9NP6GBujorBaVKA8M4tOjV5d0aBAZLgxVhvp8pjF9B
rseeTPUpAKGzI8ejCNO2hPc3fiRFmwf6jZuLMSFEokmmNcKwZskc/TRdSLhncbMb
ncnNixlc4hNRW4IaRSNgGbMttyive1KxggYccBlOz/Ljj1dRt+Gtqri0sPI9c+0u
NwOb4vsQypMS2AcM2W7bZbckd+kp2+hzxfXgwfkHJirMC4gTxJVpTXFoKZsUbCkT
ZXtVib6B26lrmv0M6Cfm+Ukn8dj2eKLDVQe4eFax7mSlEVpOf/oNiaxR0isuaU49
KVESqtNG9eYVIbzEI2EuplVdJQyEmmLPagYB4lDhaFfX1AcDxyLlZh+Cvkc1Wpzh
kpHPBGkyzl+qAovftjh5RyAIc3gz0qdpXL7l4IuGGDAr78Rs7KRssFYH92o7iKij
QerQ0SKf6NrM2VVXqUlujzk/VdbvqxrZguonWCfA4+KdztvzYvTDfAmbZtB55f7J
pjO0w9R/g7S2PBunVGVY9423EqRR1pRFZmywjvYRQP9lzLH9jsxAF/De6KYA0LAq
uP9VEsnD1bUlli7RQbqfWfHQnIBDWwXiSsaYPtskVLRC2/hilehjTYd+MKy+Lz81
7eA94oLsOphZB49K8LpLpHyrbo6jtBIOfPH7yjBizIlEb3qUcmx4xPZuo6IgnXYc
PkMChmuTAQ8ho+6ibEkFaeAKdElPtu0ZXSEnygVkbVw+IpfOrcOzsj/c9XtV96/e
dHo0/s+79FfBPaxgNXQtDiq5wCHlycpROdUynRsEsvK6H8hr2OML32mxv3HH9KpH
Zzy9g2fO5Ut/sEQ+6dP6g1ask7fqVzUyTRNo5rAnm8SocfAYc18HDMOt7qA43sn+
I6qmMJpn1OW6ZKyQwCJCn5ed7mhhdO2pu6YvhBWr3RseRgqeuQH93mlF97yR6RNG
pPX6P1Nq5Ka4frrFIJ4x37RKBIM8Fdt0mwZKTajHT4qC7nuzlYYGJzK077+z/k7F
9mIit2FGntSzdtkkD6P9Ge9RPTtnFfNVVdzWAkR+PT98F/JacM3yGBdM4fpFiEa5
/qAG3D7SPAlks7cmPG0bu65yhNLcqeJD2TuDwyKtrCRjM+J67MZ8czH+xfwnaxyW
QLt16hKhubrGsXrCKCL/9b2xg1f4soCAidw2/BJKrXtm+ujg309RHp5tq4Yww7xe
kHFSt6whYNPEaj/JlwlJ3BqKgcLPkVjLF8Sexfi3oGVafvZ54dCfV/vYoywVw8La
/o0Mnq97xVwKcgbNc5cTFxH9qjaEwSobs1zX2e8g0kS7Hbc68Gaz+4WBCVSWtIyj
+GiwgGWd6P4YZrg1cLw+SGw5SJbdMW5R0jD2yTEUf0vDx16yX0OC+5xPbAVE5b8P
rc9DTX9xtb6g94BWjANu7BHh0EWQa+ju1ZT08ZVX97+L8GZbNZYQ6yAnSUOAQtJG
WCuwU7qfaQ6Uf0iSZABFU5uvvM1oP16cfrZsGrOQug3g1CNyUdIX5sQkSh9HTyYm
EPD/+iiauJnYQy00qXVSMwzm1FOPNtz4Q3Qg5/ECEW1sxcSwQTyuvHXnKmbUgHtI
dQJoJc8GMTnUmHOfQ9fSPDKemOTAkGeIj2jeWVPrn/YYzgTUYjhu1qJtp7j73x7B
7FKL6lmZ3g8Hr3hDP/CTar/NtIoclcxY3iUu2fAYHo1Jx/l9krfEv/GQWLnkg3Hn
N3O5AoQ9/bmVCvs+0N1ULJosmof0tUe5JrqZsOVutWEiZn/44ZyKQRG723Y5HYDw
2RP4TrrI8Nbnz5sM8+kf7ZIXrhUJ+1LwnPYQC3cG4g7O642B3V/t8bD24nTgID/Y
wimpia6GLlZ/rl9n29cH3yjdNbL6EAVaOOKlbNXvQ6XChhNRKkAHGyJ7UHL0K6tm
tBDrd0XTE00QHW/0LBbjEtnsXCeYNPsy7AUk7InfARjNOOML1HmooU8vBbdDriHh
ywModH90PPTSFWq0wAgSNnij6lDnlbn+QBK8ifnUCoiyA1ktRBYUKmE5z0tqpoBe
ckEX6G3OXbSDil1ma4pOaW5XpAZsfE6c7jSnEuONqf6jz0C8j54jhmnAh2/Kxbom
jb2cHRf/TslzVpi1pW2SjnX4+o7S1a5ixiDGmDMQd7RQwI5bM1hayg1IV6vfdApj
eTt2jDkELW5DkonpQb3Jlx+I3Cdr13mfmfFMbqXNGGoByLc81lE3ehINFxdxMVb5
kvO2NXZfXoQH85PXih657NUKuz71Aq+Zy1pnx/G5YBizBof8gEC2QsoAkvjd5zjH
1AXaAkwWvW12jrVGi6Av3A/BnB30Leb3kMKHv4+BVwBboXQFRQemxNFymSRGUEUN
oieX153koe1WjxQL4KXvvlYXL5+K/fqpkrpPVxuVVVXCrcfuzvF5zMT50XFf6ChO
RMR/q0MmZQnkccd0o0f3lOLzPmzqRwI8Aa5oJ4AjC6fg0o9Q3AhGc9ZB2CXl2x4e
7eucCQ51/7lTjYS8v568Qiatmm/kLbsEU+IZ3VL07gO0YRPmI/8I4JK+/dsld8zD
y6uaI5yD9FNoZhHZwlC3Ryxege7rdSUofvoUbkcJNsOEBB/4IAdeu+UBi9C0hUTy
OmkxKBYpO4POhZSIOGThvfEDwYK6hqIooAyV/7y5WMapWnQ0TIJ3vXY1gatP+ztP
l0E+zMDh9VqTo6t+MfVQBHN36qCvGKIjJKhB7GIJ6o/XLlN8khakxA1sKYj7PX4Y
xDwHCxwcSG3wqjkbs95PLsPFcRDfrmtSD7E+eH7nYQfcIlrq56DCMUX9Gv1gpwqV
gkmyb9s9EmErVoHrkELkEE4d+FWYoJSCXlU41FHiIeFdz7kT45djyFLt3xYMpaV0
SE8hEcTRjJW1Ge504bHFiioJoMcihy8A+6LowmqidtQ5n9KVwMOyS2NQ2e6cufQr
0FUw51N673FYqqaHRtdUWbSUfHwDmbshCSkA7ANp/9eZg8CXsJm+rXBtORGE37v2
enAxdD1RUo9D1PIRAwiOZeE+xbmfd25uM/QtUEYTSzkqUQQ44rhxPdcYsAG4AVgz
Jvf0e52gqgI70ksnchZ90sXDT3FqzIwLnMwAIGYkn4Aky+XJYTpWfoWatB4YZx31
ScWAA3mu8VyfaTDiiZ/9X52IXctkpprlgrat59VftDxNUaZ1Noyf5MrU50SbdL0X
TWj4Lnei3/+4aR8Uhu6t6r3qFP3WjKdHdR6DFpcjiX62+oVyg3Q1xqT5uq4Smbe7
3jrth5LmWcl1XWAn8TNEQUMbCuNGlr3/cN+FU1kKODXiCZ64GOErq/cdDwyx3qSt
X8YpZcJNc1exwBEYu3cbaaupvwWlMAdfJGjzsIaSy1HwWRcsXWHM/+TFAryIsgoY
UGaQQcFqDpFEI/fEsS6BKfYlO29tUNEhInGWQpNbmtHp6XbvLmIgt9DEkBdZKfok
v803Ut7ukrviN4bbjeh6P+8MXrBh7XStVqGotVNk63d2k8YkEYKLQswmiDDk5GYf
401bCXY9Ua/WL8x6r/oyzgsrBsmk4Z9kkqWBfOXsp9RTn+NvZXy1Q+MkAg0iuncI
50gTwHHkkSg1UMTLZeMr8V33JW12FVGL19qcfaSJC5vC+ZLwcYMuqv5w5vf5oaZd
sXdHF8mtjxExwY6xLMDO9hnziqsZYewwCODOOaxfCHxppnzClgul7UPH1UzNI3u9
0xZVqQ5tbDEfZa8VjSqM9LUEqgfi8bI9ikC2JNyBMfwosTnRWsVzypQmdw2et4rT
UICclmfhzU0JhA6srFiDjVYCgK1+OJtxjbBmC9Mz1KPEsvZWMI+WMOOadGNWK24+
LV3d//d3Wwjbj/Hqi45qajvUpxv+TUuFvYDoc0Gmfs8zcldR5254MiRqWZZxfdLl
RfWZ/v7Ud1mbUfk2jy03li+UKQsNoOsfMRQJp5AEAHbyi6xnHxS6fo94KW0ADZI6
v6/1Gut65BvKavW7Ne2LnLchaFI++KOOpHarMvXChJX/yQIb7G0CWr+3T9YkFmH7
5GBiU0H3G6Ovv6XX7qIbC/2QnL0OrznRI1yq6ehWya2dSv+qWd5M0tjRXEtSerh4
/6sgYW844oBOZyY7TfDOo3p+0nld7Tgfz6CU0Ld+qAo48MSGQ/WYTIL6OgVYs1Zw
+g2PA1vjiLLtmwrcvJ9I5+h3wQaZlcCNupVUy6YINbZWOYlzQs/DYZsbwKWDGJb9
Ci/8ViK+K3eR9wjCssfPOxsnr5e2PsBNzadpnzZPPoBOLh6D8m+DS6hPlhBMmOz4
dSjMRJjJTOyZezT4iIRPOaVBfD/uItEcN07tL0TmwrV9tWG1QjTnfPF0zhE9f4F4
kkO8pKBnxaIEUuKwq1KCwwkptIdrGAKPdmVjpThQtDy/xJutsrY3IXk1nkyCQCYH
1pSRnvuC1cjcndsejJ3doLaalNZfjozCvyPqbAy8dvl/jpIbh2jn0BEGazY07w7B
it8mHenGmgx/YNNkaCyKbOZxSwp+CJwjPbHMwwlzBoVfRqT4r/j4z75vnNrW8xI2
gNXzrNUM2wzvA7DJ59Qa/USk2aNUw6aoFrasRUuSq19CUw/5T+F9XptNIx1sflKu
0fpGO+PK4mscwakcDtW1MbshqhHPSPhkLyBm4hYlb05OEc+h/XoQrtkddjmbbsto
AqnxIqwf0oJB5PKRxQNM9wQsEkAGSr9tvo+KHVA/JVjMcb1IQDyxi0Z8eon4lgRs
Rnawc8BSD2CvhRgKySeZ9qa53LvjucQImxGsGUyShC0SkfO3P/dterNlGSXeseOu
VFqvx9brCkgIvMY2Aaa14FPGd8JfelJ+tSZfeWGSnRS4oBk7FZiek8oc9Sgt1Ykx
sj437oGSA7Kj1+7Jmn4arKHs2e9ul3JJ2+QB33yyzoscrbdhAqpPX+JPJ+8gaTUc
+Jz3niTJps7vgWSgY0pdgtr9R2fwxyLQMtIXWflJsO53TTiimsfKTAarM8pghW4b
kWeMS2DON2BEht9qWeASp13/mZNgrkaEask1t766geHfThvb8PKGjXRgNMiVhG0/
JkIqCsa18GkB5i+NVE/gg2AWvu/TBB+uVvGhSyw/mgN/AHkbGPbtCmd5h+v66yLA
XVxEq/sHjUHVbw1BhvmmG0WXlFjw+s1Pv7H6VTrVVjkaMBH6w03ZBp1OoDfgKDIF
iFsO9FWhVWMQdpelZLlWQqvzuBwfRERvhUDB6opMNv/PccitylgOAEu8ldQOFtUg
i9QcChiu+LUoCoFFiaadcvl+c2irtnCRDgXEqNdrfU02SP3LtIzM7/k4yEZwwwHy
WW6D2Jph/mpgIDK+9K844aUtOE37MjwOG7otE1XbKGEJXZpHNB5Bd9onyz2hHHp8
USHs1pzcIAdiv0beM65Qeypb0j6smTE/v8ei55oMpkrU1PHsDxCH+NeScYmoCb23
VHGQFZUpTHN6M3UPIEu+3CWmjHT/NglkBxQsvE9QT65txQgNgileNZELotyH2ZaR
sEYQvbq19DJ3nauQeIZ+0W3seOY5WTvKB0qF9F818CkYZrVXc/dNS+4EWbZthjuR
74J4Y15iYLNSQvCdxUlU7gcctvMEXdUDvUPUdDOIaObjn/gFrIBKuYYESBLPMUM5
CWUURL3Mjr+67GSgQS2yfC1/TCBnL4TbRJgk14Yt7mA430FGd4pzgw7V+pEOgZSp
c9sXr1NKwAB7QY26q2tgW/vA5JWpdk1tCGx/QBL0rc8HmJxYeHa2qQfunKog7QPD
YtryjpsQ6wsgNuJMktgJsOYof2rPx6yjeAuAO9F5ZuTIhibtnZgOXZjxOXVqtBdQ
4spME+7atwf/n3ruR/IwKz+FNuoIvHPFK1OrIbSLMS7ulJFvR7oZ8yPHNK/lvDMA
hty8nfbtnjm45KuZP5vtUmsnl+rz2UyiqKAa6h2LyNlTqBPCwgU0KzWr4w+Pu0HX
H503yoU1vbFXi4U4Hf31JiaH0BS1WUgDI4cecm4jC9AmspU3lGPdJXIl5P6RhjBp
bVxAa0y+h5M8q3FYtkHGyBQIFqvetPaJ/Q+PKuso+ocYA3dCEJiPZdTPCcuva8k2
S1zxGHRB8ZVQovOlTi+HMohwAoo5w7TG991UTChg4RoykzZq1XFz8lIY4+8paORo
t4mTRZFprxz37LQinu/iBCEIJdAjHBbehOCy29VgJQyQURVXYIkWM8PWLQcJxkfp
dA6y0RtYPTmeOTUBzGQSJi0F6vYcmMQ2EWKiZYsEOwQSKhWWhbGkkq2v3MsNI5W1
U6qcaOGT5qSwsNf5SIjYfG6+oTc+lX48gqHBiqZu6iupx2mJNFcxqAqvdCv4m3X5
h9nKjhctc3/G1aPklJRT5MwqyF/BUQSIqewP3eME6KUFYm+nLvI4V7+VX2I8WEe1
GmLDUeVeIFBElzLbpcd9DUPgkVBbTEbMs3ix14gYy35gSJMhJWCy+BNITe7/X3Dc
jIXYXuFDu40llJwaxiC6yR35FBLBZe54z/Z4KBoGCViQIUCrzi3GqKyFQfGcbDqq
bYdWQA0EFjjphRmtVkULkgzRQ3iRYUvI9N4SWJEvyc1VKFl9at2ot/+lrjR/aEDq
sLaEle008MPr61kCv4zVKztSpOF85cs0cMR1G1uRjH+OVshJdxsB0UDKh/Ywfks5
HgDBwt93WowHgCDrfhStp47h8p7jJQcAN3u8C3SKHaKehipq8kBMatiIJBzO6LML
+EeVUWPJEoEeROZvBlq4Lz2wy6xwigGoS5LmskwefrmrPDie5DJ/PVAAcrKXUPtA
naGlQ0fSzLVz5S+/UZhqwIXXxus851SW3C/7Yk3h7xK4tvkmfYFuBNB5MDXy0h7d
6DAB2hIwb27OBi08GhId6TwmaGR56mpuiU/WNEMAYEmRc8izYHh31K0F+FgTDufB
QPUZcSaOltDB8ESviUEi5KFpM9tw0MUoHSWJeFxJW4ItjRB8kTYuLLFXy/18uk0z
GS5YN/tcJiO6Ue8But3rIEAHnSP9DEiE5T45t983h/O4hrYvFDdO5FS7/mbjbbqL
hp/O9I5K1S3GXZmgaAvSj1brT7opZmtQ+qwRimccEA8XDBq+Va8WDtVlFpegIVyW
MSmv6OUv2r0q/xEwqxgu0Ab+yk25n7Qcp/0QNmXMGeVfNw0KmZp7+p6UMPb1AX96
Lq47pn0dCt43vugtdM9VLZqrlAKUxGADi8Zx2Nzl/wNz9sUGt6rArnABLcUlMjLC
VJwdyH6jWm1vak+Z353PVSLQjHHnTgFFMAOIGdDDoDUL32WKJ0A6/sq8HHDFjpEs
kjAbq6mdfZDunuZ4Y1qikAwyvpP2c4PD/Y/JzdGffWvB2BsJ5dF/esfGIt7+rkjg
QRKBDVHGftWiohD5mOkWc/JuQU+CEe/db+olzTIcOb4a65QAI6cNYw4V1lR8HwzD
RjeJgzJ+YKvtKiN2Ajct4ieUgnVeSJxgu6bNV9EbGqA7zZKESEVc24Yk+We5pfnm
P5ODacuwLc7nBGEHmsmgBnBezgl5Z9HLdzNr7X+qxnBfbSrrZkYfi5cKgU7W9un6
K63DylsNejrt7422/1PEKccIR74pe1pnMm3Kj+loCegpa+vA/oa1DgO5RXw4ETJi
mHf9w/AHEluuN2I9INYDBMwsSG91mPUU/HqwrSimAOeQKR4tpGHMqNPY0VuzauCn
GACbx3Z/piFFwDy7RrRoJwwAPVMVpjLsC6FH/rOhc8zNNG3yPJ6UfWOczr8uxYvg
wStTqdAkPCNLAau2ScViagiB1TLcCLq5RJFoJbfzOa1SAPRkrh974eeQkuEaOxzX
9YFJpOsH9XG9NzCYfp/9Akau5568A6pRjRnQxZGQ4+aCsaoRXjNzYBnDJwhIySUN
iBzEWUTlLdr+yrhGs0QFzJSVObe9dGk6rBzZcYKS/IvJYzApQZ5xdQHG18T7brj1
KmNo67HB9mqSrnrPNK8JwrQPpqTEI22DsH4vV2PWFOcmJeRD/yFdYTCvj7V4NDro
hq2dcqBvaq72E9mg3VJxHK9tG5/BTETfWSFlzrMnO0A19LUxzbOUKsGTGfPjGjot
3fTw8N/gcDdKmYLMfuQuxAE1WZTv1cCaMsdSSwUP+4dpJFa6DvD+QJfjSCihFr5e
iU1QXHXM3SqJS+0j5DTUFDzAKTiEDI7oYhjmtSPt8E6HtdgsmQGP0+ulDwUE7RnP
++8X/gzR12jh9KBPYXwkoU21/zctwbbyoJVE5KfV6NWsRKgHeGuwaj+N5hXYLTcp
jXTewuJe5/okAN9yA2tIJuHimhvo35W7xukEZuylwAmG/NDzvwOHrlDJPnlOazpD
pQIMX8Sr67+/KlJTvf5aZqxXiPSduCpVzCoK//ux5mhQyC7Ofl462RbW7Qz967+e
SMcgPpmTsYnJk4ZLhRVr1oaqXB++ZQljDA/6qfYyfdsZgsREajMzlStJaW9FJVIP
bJ7MofHGmOCfK600x3g+Q/kJpP9jR5Jo4/6IzDM1PpR8ex+SJ1Q2IcVimXZavIbu
yMU4BPWrxjwbl/UgJxPqx9gAmw/4K9ravT5xysPOvG03wd68SooANuXThY8oIGCG
YOqXTfZllab18tCfgkrwc5+EJFegVM4j7aoDJIW6ucVq7Y8sn/FEaDFJz913oxiG
lDc1fk91JM6FkR46+6OLOOpOPOCBt8kybyUDwojmaR85ujRvPXv+Bl0LIv4oplOM
F/O6KuExDgjE2ZqPOUNtgKmGwrtkdmdAOFcW9MUBGb8Ksn6CfbR4/pfNKFjE0PMN
qI7qzC25Rd71GSwNcATH6AfLU4E9MNWgJ090xku1bRIPhI/7KNb+39aWHK4qt9Ha
+CwO82/el6nVJW+SVrNhj7w4oTUKRicSsdGaLJIaeSALA5/mCA07zvTvlHOfHyxh
0pIN7Kd/vam7pmy6XbREzFHoYd8lR7fmfjG95Rx/TDMVl6w1JgwK2nMbbd3iuJ9m
WrA9pbnqAsVO2MwPAHFHPGaEZakTC1VIWGmkl/ZPSp7w/2NMjJERrMJ7zgthBlJF
svsFdc9AU+wXoHdqMSrumc3lssWIsKT3GGoAIdkgj7kXRGdYLWNv0aOJKj/G3MGi
6jncRnqXfOIwjLzYj0hArFM1q9lmlHDTFhXnxMrvlGr329jJj1CSQnnEbHT/4dOB
fMl7+uP6ePKN99bcbk94C9verPS5itrwiZZlondcq/ScaStZdPIUaQ3b42dJk/Wa
C1BK7WZMapGTsFuNI8sUQFg8MXdFb2moBau6Lhm/55PN1I+6p0+tVabvzX867A8N
2LnWget1GImk6d5syQaLy+dh/ubq5yWiOpKLQcfCZZGjfDdr0in2G05U5l6cgK8W
xNC8MKkl5igzhQyxoX2mtcdLtALXJmniReYwgmhL3emGLBCjXOoc+bqqFmu9VAEA
imj5ISO/O4e5XkcTbU3VUyQSr3bFpwNUq+bfuR+buSI/pDf5an17qILbLozUCvGO
PJ/ZtcKDPjV+n/8cfDTwCKlOQzVC1PeaiyMpHyu6knrhqAEE/R3MlOiv98HoNrPC
1k7yqchdIb1Q0KZGBihiLs2bN4GWxnzkbw/T3r8jCrTxZolpvDoTIXAYCc/jmkfN
RZ79/XrB8WMwfEeS2Unn1KlmwM33Nh3ksZZx9BTuVY/eGbpHMWfcVDXQNbAlAIe5
qyRUAHrjObhkeuJ9j5NDytRCiwx2AEvtOLXXJr8IAut67s0LpT6lVK+lz3GO9w7F
nfMJ61Jr+jAcDnV30RngXcjqneqXlaRcaP5RV+O8xZm+82DxTf5Aubm6E2IeBeug
IOHcM6jxKBv3XcJxJ9cxLRwKIvmyXUcGvezDH7Oq9QCwHvEf/wa5P5xDBgTswnkr
pMmO5CFIYpIzGLEQ7OX91LSVojUN+vpAKwdA6yY3grmArTAoU9DtqZ1EQ2OGcEmP
VsWRSLFU6BlPpFrT8yr0nj4Lb/kUt6CguNNK+Eu0tkfC2RYgGu1j0ielWi6mCDxb
7Sis6pAGDaQ5jMk0cBeG/ky/uhL1zASx2qVItOyyZ/GqzNz0HdiiJ212Dl7I8QT0
Zxu2KcLrlZHPKb1+4TTxBGDcSmZT3V/VYqFgU14hU5NMPMBbZeE4OWg9p/lV48yO
OYCWvZb31ix4eGf2T5ZwR2H7SXBOAOTkGQI+424DDBrxTw3wfQSgdebXCUIObByW
ewXnSuA7ncvVE+r8hAdoGidoGXiyUk9eaC3ysO7SY1RiTmq9BhlkwoGqmIsWg58l
Ai6O3j1460g6AvUSkbvCI80/skMeQsNXhyb7/RtTL9ns9frtVb3xA1fmyiwK377L
c8NV7liRsrsPKpa7W83yCT2INGX5806ci/EDnvdN/xebWySgixFIFMQII1CzpP7C
rY5BwTkS9qgurCHeFmbqyiMEQOPGgcCKXzkLVohL0CXzdakXKJ0xn0zXGMUZpFx/
34HUh6ztf6m+VZbAkdTPSzEuFD/TkgLTNgOk0yBYmfsDVYG4wJjUT98hAfdaknIa
PLLSnw0oYR1YKAE7bc6D/uPxlhClsW18VA4OXgb1v2c8z9EBdj5bB9WJ1E7+poTb
HitXHWos6ngu1MOfqHY/ctVMpTdpW57a0hz4sAomMS4g25mcWl1bQS5nJBpo6myI
JZdf7F1yX1gygaILvhllDf+mkWjMNuBZ0uBB/SBPYu0KTEK1m6RTyzu4JjJAduVh
D4/DOSyLmcKDRYiLQc1FoiZ1dIpQh6DW0gUQR3kLeJPCw/aAMpEnod02R4UO4xyH
dx7QnvnEa3uGXQuQc8JycJELvjHBZzxuk0xF7/TK+m0rJf94pVT1qWRt7SyPXnoV
mr/b9rZDtYwgwQZocr6FV/9fhPr6585YGDkxe3fUgX2VPMQ4OgRj29IlWkB4Ak7D
EM7jqo1vsuuE0KCZ+4K8rMq5PRWcfpZpg/L4150ImA8CUaLUR4cBE12cL4oxvGeJ
mxM9D4/ArIH9xVDX2manh4yFsYqSOtCT9ioMyn8wWAuwDt6jTZ6xtq9mYXOAj5oj
ECX1Ujc4lnJH7hI4TVLZ9iwVWCZytwCNtDDnTI44KTMvL0sjkZNYXs/sQhp3VOiC
NqUREMLxX0GPvlRw1BZyT1OHlwWHQFQvTiaazUgdwLy7TpdriR3dK6G2flO9N8d3
YqQnGLULqchIPColoNoIdyqy8TQVHuAV8kzi8F1HMR7bmRHyesB/8gZQUGa6UwlG
dCb4dwVMYoHmKfP/Q7d0CFsg9X5LfafTEs4CRSlxx7x1Hh7rry2x9MhOSQ2wsnnb
LHoVUkjvQIULVn9JcEo1/6dydV6A7ZFxoq2zsv55FhFgjIUMQ/RrbqUGkmPejw+5
ZDgpKwCEqk8tSc0SbMk6okkJGUpSQ9+8UDuD/JbIeRWb9+IP9fGrjzVklvQkCZwl
Dlo4BJaadsaSUev5XKD+uCX8DRxv+ZsO4la2ifK3TQQNjxYWjK3tFfKsAiAgECHd
Yn7jiS68wGZ96Xqjv1yh/9jk4ed+6lJ1LZvo3c5bGwqupG2/oqIDUeBvEwxHurlq
a0OvD8p3Mp7qUg8ep0JDX/4E2SzowJ43sZiWahFkcviHPFFBdFfbPd5alhKQsA3B
Lc+JGLTu6dZ17InZo/KhrLk73w2oBJUHjOd6drJAZHkLyz3tQQ0LA3ycOBHmWNmR
LrIk1nNg6SjOXA+C0mKKWXKeo+GWf3JaZEE84g3QXJD5f6iwvcinn2Mycx00vkdM
F4DzQwVRZbfSboZTtSXp3ryczGoZOGde6qpT+doIfRCXLR92hQxYNoK/YFoDoXGE
d/JPqUwEIDGS/KA7YE79LugdFRGIBi4cHfaMgSHq/BLs36UX8STmffNKZYTkqPVb
xGtETKdnGpP5If+yVYLN9bsxGZ/nRHgaraer4wrqQHatzv2hd94MYH7zW4vb40rE
hK6aAzVP0Hd8f6AuQzYIoOl1tDRJGDMd0wKkGM/MpMuVVsT59RhdcggyTRbZA779
Fc7z+UwvaBuvgIMDcjq88nXElkSkkweWWdUJXr9Yc5hg7wYrYL5OLyc054zegUKM
uqMQyJcFvFLq0K5bUQ7lWuss3dKBnlFitsp0XMVAowqc9/vuGr4JhLozq8wnJKql
h5O8c2OjNjUO3g7r3l/nBbMU6ZrQTA8EShV7YzF/43e35OzEhaAly6fOjZqEOIOS
cMzJ0QFw0JnLtjGehaKSB+RzhoMMno4N2n3NYz7e+gONaaM3hSeC3TEEOmICBpf+
QmpHmTimwSp0b4DUoyoAw/23QjiHf0BO2oS5XKlMVqnMSsDEmu0LJ4Y4T2qfYFYx
dUvcwlbIqGxEtvyWKW1B1GqxnhbHCZkBoKYr/B6HXxhj2a5Mgo9jS8j/6ZeCH0U/
iW33spRmLifd9Kz/EKEL9zwbdBmG+zjSD1Lzy7HHCSIMqNFy4JtR5BoS+7oG0QSV
yV6tX4lAZ7vC1Xy48fZqj08cQ1NCkdIrFkRM66wruoLRQ4B/lzxPpOOxEBTKH/w0
uKx/F4/i8AvO0fds9Btc9QYJqWl3ZRB2xVxqEBLqn0isQPAf83NWB2Tr7+Lk2qK0
fk2dlHmRfFDurwrt47fPaBqpEpEFGPUTAo6v8au9lMLWKZQ7nBbWb3XsLJMgUAXZ
6xeJvraFcsPMUu0gRtsq6wmkjrbk66IWYh1JC2GuJXHKGPYbqAvV1UU2pwntXYGY
fR5SJ4W91AXyoG2bwdW4VelgfR5RwyDaUpu2QrNJL7BANrrASt0jPcOKlJSHfaZP
4bhEmyXGyF53MbdLire1BSu1XLny8d/VpI09j0Bciz/+f32WnG3vNwcjid36PyIs
2e2XFQg0LChujynUxn/vQKJM/SijKe91J/py0kH1Ob8sw2EFLNSD063eC/UmKdEo
/wU/jhozZVDKRkScwuX2DAm+uUJhOqhjJ/OzVfDTWdg5TUd85MQ5h2BhN9r3I+Es
GDbOOMvZ4VuW4+YitX42koJ6iuZuzBX5xCA+tk14YIMchCuVmDbGSRV3T0FfiP+E
cF3jXrmjOcW8lLOj4cs8mCZnmpiJtHJd6k5acNuZAazHeyutuDiszE4ExYTh/1/B
WK/HR5zFobKX/RTvDMfaH88llqi0wrUQZEjzDIGQRjiyrvrv/9S/rWmcRkXTEp2W
t/tTm/hC1eJOm8JQhqHE/nS+OKAy0vN+cH9TTEWxnZquA49vqvQ0thIt+fcLlKlm
Kk44wPZIAk6gvcKH6CBYJnbb/p0IdVRlX1GRtrNCUAuzq5ylqLloLRmWSFKSGeUp
doKu/ZGMEsnLro4rjFA9Vfv07ze29sOoaqAG7ug1/bYcNI2BRLTuUntMLkZK7YKP
fEPzKCR0ageVLHjSHiheIw3uF7svHVtiSHBjd2FgtogFg7wLmsz1QV8nrm/mNASF
ixlR2RRqUtBXqdrB+8WI2PCPBYjpWS6rr212T141ZL9cDUphgwJag7j9OegHd69R
j/zG315SAPaBQ/lRRj5LiuaCvVlyiztFPIic4V11StlVolXE3/Fgl8TMesNwg5Ni
srxVzSjytkfXdKB7opPvkbl3pOt6WqH2UfmwWDX/OuVJo7sMhK5PpyY0TbAzYjyf
fM+olNbixsKCFUodfn19zgooMsFMpWpKcJqaN1s7xWQVklTOnMpbpUMrIui6IF1R
Tpu9gxfFEIT6pLJT2l4kQG4mq4O08Rul7BBBLVKSz6gxHrv1LhHC284g5z36cSQH
h9wDuSj6/po5C72T27gkaFMdPbHIZ9lbbqiaLpWe+X05rUsWDix5/cJMhB0D/unK
k/JpOMjg59EiQh7K5cf5LZiLpGwYgYY9Hig4qi8GJbJeZA+Z3nYcwYzNWlSEMfjC
t5SkdWHkfitybmAPCFFXbIGBP/14tbA4iT0K5GA1LxM8TSAxEo5iyTkWfeEhTGNa
yBN5sVDbiGgKuziqzFnVikrtz7fv7u68U2n2Yx8jI/fEsKdZst1r/ARZUl260XEk
Bs+mdL2W/1YB6ncBIVWRlhsuuif4DUk2J3oYs1W2X8sEoYERHwyxvvEZfztjIndI
P26Zmw5cAG5N6hWoTcAa7dX8Wv7vb+h5/WsheZgMC9zJDWq1DvoK+4YcXZQdYBWv
uhDsyFrln0sXvTHDRxP00fKDMbeNr69iudgTxqTEAFCZpqAf1sNOu6aZdxfA0kYL
sZ48BRFYzMtpgI38bOM1Mv6ugA8UPEgHC2uvZ0lsNQLQ89vSC/qbEDyIQU/MVXjz
+ndMcHYmIJDv4/SdRMGITzX4k2aRLfh+A++LyFSZwwV29aQQ0FgMf1OQiL24ZJ0z
XTtaFg6vTuZTnUZKAhlOw19qG8Y2sQNIysVqHiK6j6Fhf9Ijb27vLsWD1aPz8cy7
t31/u3bzV25VhHZyBAoEFlVINY/Zwdvw13M/glwAkaM1MKudtY5Vha/C6FBuwbQg
BXqZCPCwHjOlVF5iQ51ROpUfKWpUtGbwBGXtDGGK1+wtMRYxyByxDgOybYGzlNSP
QYCFEJuLcaeNMP/aQbJTzzUSm/8Uya/dCV+W/2W2czKLOtucA8OZi0uYFgwGO6ef
5sFuJ8PTjsx53qeM9lsDh4Y8HX1Dkk6y0LIFzB/AnxZfdZA5gz4juV1+UfHS0J4C
OmzoIBqS/GV/uHn+OZLxakRekgIN2Lrsy1Iu3H1c/maa3UaGtV80l1mqO3T6IrV8
d4t0v3Rv+bzRDzhvjxHSDsqfN+HM3ExkdQ5pACEeDgqMg3D8GO6C+YxAgkjSXlFl
WgXjMelN1hJg10LPjJZrVh4CqyIKXdfsmi3aZoVGLeMu1GENF1llfWRIT7eKUBuD
yCqUoi2S39HWBaJbwh7nvqXDcKRVBzx+AEhUV6xtYTNnm2QaTiXTQBC8I/tbWI7K
gU7gAQoRPAUZLVljOyLn8Cq2f+OudOtgGSy5LXX+rQhz2BkeMTKJUu5T7hW5AoQv
uxtJfwju9bPxmFaJqBfsy+Gh2s1msIdRusm+tDM33LoRFt498lpt3HhoZoZDkda3
ySwMCZzKQCCHZ0TBo7TihlM6c0SpUUBkzoTT92X2SXJkibuYPxmcC4cO79h+tKJO
j9G2JcZC7Y1NhM8ufJNCNkfXwh3BOPjXR9hC8xwCYhXxfMfsViqWdcxm9+FNXsLC
IWSR4ZQqRsSy9UfcGNEwPVcJB/nbjditwwgV9vkWpzkfyr9GNG98naJSgunpFCjt
ZhYMLp7an4OJhGz5u6eJp5+mVCnSkRIaqj7O6CqT2Zrp7MY/ho5JIpypjPRe0HEf
LMgKjmSMIVwrWuwu47oz0K7ZdhvJr7AtqaIj/sHjjINwtcTM5PK4ch2UEeXf5IpD
iBuqd2vMteXpaoUZWpHi++RZd/AThpeLaagPjWUO01H80+S49DZWJ4wf1TztAFQ0
QDJEZ5aFMOUZOQss9R0Rbe7xvZo667UBNbSUMdVHYL3/FcuAw9Z/HSf0LNX3Jagg
ti0VGIL4O0OdYZe9TGz06eVtlUSY3AN/fyHLxaaC8rdLS33X+DIhQPJGmfbLZzL4
y4nBOJqAuOumjLlJnUCZJl4k8RuFr9EEUDwYhSD3iDjbYWls1jsXyyUa/NHmfMfF
Sw9m1vYXPxEjSSM5ElEThb46LpHuiebnZsqWfNdt096qdWNTb5qp8cg4zb8ve0gE
OrVfTzAHNd5ndjzkf55virskaY7HOp8dqzWQ9qLenj6363OVbs3kHjPJlZMTu1VR
9v7rZGfc6cPerWS4p7yfOKfN3P4jouzWxIlez/qrJmQ1MXwVqkajYKlbt+O15F9D
uauTz/GAylAWDjqUW+hjKgQzQg5wpY3mEJfj5VoZs4X+58PpvYVXtV+O3O+IIJZu
R7VQw19JE3FII4kA5XnHoahWySjWKjHpCxchpSSXPtN6VlavX3n+wKKa9QftE2nM
aZwHRwJGF0bUpUlM1P30RO7zViVj9dj2XlgyDW7lIaBoSJKiTxRy119iO+4cYAj4
MbzfZzseuQAtD1GC/wHYOi4qBzJLXRTb0EkffxvGxnc/vy0sNe9eVfLE+iDoMB0X
rN4yMBJ37z/dsZIwzx46CfwTN7cyChbdlJ7c3MRESIFc3KmA/B7BCWd7Qe5kJcID
bVU+MNaW3ae3gKjGz9LG4PKHm6FAUUa6Vtc6GOFftrfp0wMsUskIvmgMAP2kt8Ja
BwbRA5Pxo5C8Vwj84icX7pfqYqHAj5htnRrf0xcoctmIhK7eF6bavgHdVQy8u00U
L0U5SW4n7kiJAZ2g0bckCttcXhQKObID2fi4TIFHH+ideQsYvt99+8+OttRw1fT8
nRGhKdSzmYspPRuz6v8V8/P7WlFs56lPyCDRuoFHXvIeyYttOrvOe0qr3q3rqgI/
6eFJeC7USBeh1A9P8egW4i1h2+/njbUZKE75+Po22z+m5YrDNpzz7lw6WwYSo8um
Mv34B+YIddFVVnOEDi2SIindArprTcME9pB1OhG3PranDMx/QtoHhPprNC99IUMo
mhFWt1OcRXE8ItDhSvqeDGgF0lIyJ4y8KIbsdwLdFLDng5Ika1hhRQ6W20t1b23A
wbXAWWExLHIr2pQ/LpBAVMSsasmKxn2TZq2Pf8Vt/sRRJYjQJB86AOPnwSDXfmAL
xXLUee83QpVFOXvCHTJjAKF44X/vC6SfN/8GgebrtoyetjinHGQkZ9HjAI8rbxGI
7ORdYDlFvonn6YYxcpnAvG+S1u+4NWJJSt8o46uAXxRSbW8UyMiBlX0e711I+4ld
GjkNYd2UJ5IcELHKNpwPWEUXEuT8dUqI/HhKGH+I/ukIFuR43NphsQOkn/7n5lgg
NANtjPFrWGusc3WDuTAyZzIxRY1FWpH9L/Neb1KFZDVfRyV2bcip2n7mbj6ZxRB7
qCjHqmpvziAoqfarW+RpTWqTEhCxARYz1MZTA8nzeofphvA31qiQtQQVZulLcN33
tu/ITn8iWOob3m7crdYwdJJW2Bc1JfknVmnEIGBtvptsR/6/H0Mz6nQjzpz/YTSH
sd71zJJ7Rd+D0SiR0MwrSzbSm7y6WdFLR/BUj736IjHTzAzhFrmipwVGrNxpRMoH
KIkCBIdFGba/+TNdxh1Jw8Sd2ndD6/SGb1aFZcOF7V1167c9eiaH8pbf41G/HMO3
DUh7YpIApQj/Oic4VeaWAWR066bI19Zz71sfWPKkgnT5z0EbDwU9CNOmWrGHGIoS
D/5np42D7a7sAYup2zEAOi17mpCh13SQyuC0zm2TaK/S5A1UEo+0ZG8xgOA5bxus
ixraHfDbRNlZxuoOxwUlMNpK8aLewZznSG9KzVOjboffjYu12BJK8iz+WdVtMFYe
LgdxxTLCPgQhvCXt0JM3J6RCmK2XG3w3NcFeufvQoBSyIbstOeG+AxZxx0XDXbCW
cVjbZUO6Jg4NrfXmbnNnKheI7FUZupVoRktb8ecEouPAZCo+j5rLzhalKotylhj/
Pyo7uM2X7lhhkfnVJ2Vr0Bz5S4EdYk2lII+BzettamWBgHOGtgDJJsnqDt/nv0Q7
6cdXc4BBvDwZrvMbga25k0b/Cjl6jDRwfccY5VF8gdTBrFhMFtwSeUGyQfAEEFCT
q4uqf3kCvDer7mY0a4IkxQa73BFl+xk3iPUPsmsSM74VzScN4RK9RdDqUJFKSgzb
2VEv5oGECVHvIWS6fe6/uynftAvHAuzhKD6pvx+FuAW2xeQ2xpXwikYsC9hAGZvC
F3wIEAar0BP/VpW/jrDgPVkJPUVAd3diq+/m2H/7bejBHaULNX5zv13eeHrjbiUj
mLIBr7VumATDN7rLj/tdroYuPaTe9zw+7k4Ldiz7u33NjetKvtbMk4v/A5wm68Nb
AdjaQcq5DpMfrKImAJOkKy7XmMtfZntcfAe/P4FHLi3RI7qqTOerSVkHbWzM2FqR
uZ5fmyPtVRCHVBmv6NPtnd9QuB7DmuJ6z2hqocWv/J3OnNXF5NPRWs5Kq9Z9lky1
6NT9ZZoSSnd+Aya13DgsxBfZ7gxoDy11udjlQbtepHupeAhrDDU/PbfJYGNG1kji
9l41OvsNeBsneXolXEXHoXxTTckOfx/f4jqkKKBOUue9q1dTNE77YOKPnUtA8mXy
jxx5Qvf/vYSlmfcRP6yBy0b8CqElsdv4OZNeL0A/QGeoQOkPlU8MyRsvvuL/8374
uvToyq0kRjghp3/fKsbZt8wjeGKIlN3htci0l0TkxiFlRSdUITA56bcIcSd0xKjw
jyUftIz9BZbf7uQK+a3EI5dTaKDDDrK344m6paQQB3Dfph0u2JZd3+Vs/K/YOSHc
mD5qJJhhv2QBF/dU5rPZQDr9KFdgS5z0Wc+B1nslkar44rD/lq5a/5gX5mFaN7rZ
3pFxcCJr1nlTeDUan1mHcYTJecaZHHdr+otJPv+1ORDc3rdDW7dTxVWFj3gwoveL
jwM0lzj+zbnsUtXFxtNkZfs/alkdkc69bgjyQJvMc0qlp7B23+57b/bNU34D/c4m
tuXZrbBKhT/iiIMlhQgcnFq4wAQJj8GXAttR0Dw16UaRGiol0JX7Dp0cSATAZ9sp
ARD8fBY3RnbNwNe7k54whc5a3kYQpfbhxc1oEXQRTb95zBA+Tmm7ctFYoWLJQsjj
T8IZUKm3UDFsTLTU7qFTiSGYF5h5GisDzuNYVmWyr1McCx9WTkIa5IZevaPhQdWA
T3cQOAiAmQlbaaR8Bn5spv3a68HuMd8BUfgj9j/MRUsuWvcs9poObaQ0gr4WaTul
XUlmJwo4Zlm47VoJ2Zd71Q9NXO3aRih7ngm3x7CU7WXgDoe/Qt4x2U4Rc2tK8kTZ
v6X/UoCNfYqyTklk1fuPGgeK+HMZcaueOekBKqN+mgikT1WMHsp/6tnO2FRPcMFV
7DfP3znMrnZvJwn1g/uMESID8Xv9uVQK+RD0MPOOu306+uAWP4fqwy6mqHzAJUjQ
uqE/jIIncXwsjwbk2tP9tEYlNj2YMzzdV7sV/EBUKsFgeTie2mno+K0RLaOa5C5H
GP3uCrh4tCzLIDmo717m757OFTDlBBYAclP1mkTNAngk5/xdaC4RaBmIP9XfIHPQ
lEwfhu3mPy6nTiMAzx3Duf+M/37Oi4FjQox2n8mCsQ6IhTULADj9EdR3ljhdklSF
9hkQkLJ1vfmsEkw/lOee1tkaNW7JC33DpBIB+r2Gan4H93FSwLVpcAmeCWATnX46
NysYB2pqnJ1yl/pfvCc0nUuUMqssFun6V6oHmvFVm7NcAJcDeUhRZWb1CQmpxCeL
K37W+b2ZYE43eK8ARy4cExVXRmCrtEPdYIuJ+ZkbF8uwUz5eNW+cAiNLVuAkDIcU
a+sbSmLZFYOG/S11JVrG8d52ue28a9xC7cHbSj59kxWauQ+uxhviCQmHPl09+ijO
w148jcNzPEw7oLJ7h7fOm7YHeJIoi+dweAskylPPRnJHGhMgq0svVm21V7cg1tyB
7exgCGTpxvSsOjaUiT53sp4mVDa52ZF3or+6ZkJsDb73ERM42up31rmGfHUzSGpa
YDAXi5AmcLlo2LSvN22jTQ+NMAS+RrGdrLTB8bM84Qut6TLw9hGk6mqbT+7bSgr7
2o1RZaanafLQlhTQkleb+KSoOYRmlyXZTF2+I/1CQ7GwlyQDpcJYbwteOTGpiNhy
MFonMvaAoQyjRwABpibWECnZjo+/UYabDoSjs7ezld9LuGZOl8Td2f5zG7YTzyIe
mPMXSNL0VSZRGroMN+Ha+YK4gdH8uljViJDWuAe7dkpAk2KMQo4h1Kqq7ylFfhwn
ylljuTn7q9CqNBR0sTswpyntiJOJhOcDmk5zxsKypSJRRGcCk9YEoXCawJ06PWrG
b8nP/mOGgm9wchX9IoqJ8UJvZfvX+LYoF5DAHJu43WeY39mRlkEIfKABZs/ltdUn
K8p9ibEeVq910PUdhFxElahcd6lUji177JztgIHhD0AM0bc/6NyIBCfTaQadrWQk
HKfzzpzJfO/hx/inLWYtgQEwQY7INM5/xXSWvBZFZMSjVs8vm9QBGJkiR3vHwN2H
4bvCVEkoyhW4ft7RjuDJA8sjuFldnSvbEe5rNehvHKerWL1O+wt9qSrms7bMfIzy
g88bVZs8Om9I4FtWjoLxub0MiWBuBP7pii1xLWjjmPZXKHHCx7i3Ofdem3UCdAii
uHoN5tugB36QxpJ7PFho/sHsDSdEeMXckYE1nOSw2RKyh8o/bMqpTqxOIT9yzEXq
DiW7s0h+iHsFF2Ja+8gDWPabRqwiqT2FUzGOXFjUh6zWQgitlh554OeHyHix+xKB
BAx27tip49XUTfJjoDHdY6giVeIl6Pz9+zd6h95Pj6u7Nxhq2JOHgqP6VqeuRKvP
3oxhm4IMEx4bYPYOf1t6iL5fiazNCpC2y56quKjjQ6Jd0dY85PKERBNx7+Zt1zo2
sXV7527WLmP47oGIdq+23E6LNLwnJm1Z10NFO/niaf2YdhbWV2fndlSVs8fFpDWF
EEPFM8O8GqxdkgApDUPh9pTaIV3ChjJtfD7++k6yKCRHR6rQyihvnyBsUvBL8vDB
UUx2/kzPVUTtqRrGmQ+sBq/WFc2GJA1KBBqUV3716OaN8hGklja8w4npe6OKgeNF
4C3Ac3DUVbyFtYFMyPo1N9LlZYxP0LNxv8B1ARWWezEJH3b4Yu++S/seHFMljZRS
xrkEklc1zbRBOE/Qzc2GzLAMVwCIbNFEwOSZ4sXR/nZTaw9h5fl4PTT8BKqFdxAA
YUuzzSeV5iCC+sXgZ1hSBtyXccdD4MARAm14VgkbzX4Yrmv5ka/9eQFdUfqz2B2p
jyz8p9r5CTPxP3O8KfEGBhqiIA3RdyvwYJpuBbo3OvNnc1JshPyl7rc2orTGnNHe
cDl6fWcOL7d0PGXrZ5PcHelutW2Jee2IFkZhdP4HP99Nn8rtX3IGj6y2MWJeN65L
BcEN3FOb6fLke0lDbYt4b7eISYowMu6Zmt7dpmr3/JvE8DLtbyvrDms3ckQef0YI
eHeB9RCuntyFxfI20vRFnEhlqi9hjuIpFnTjokkLUJTO3E6T11DXTMToiyg0uAYl
yGLT/7sKG1LlOs9IksgETl7ehkMK7cyVtSKerxYIC6P3LYJf9fS1eBXACVgFDm6s
jxKINwp4xPCqtZiyRx8rJ0Ocmz80qCmN816E09ORhwc1+62fLwllWoTIa/e/c5y0
kc51I+wn/0GbnAo0Tu+JR2SrmJuJkIgOZWuBYGJzBLgZ3DL8PRQjjYFgh0/JpAuK
3gSKTF6Cw+fPkTUWq1KNx4tMkl1RtxJ7PEJEOmo4+6q16HGQTLNWsrGXKk+3PhUF
A1XXaxezOtNZ4zJQ+8611XvRhQS9ZoaNeI7PA7PVxhpMJsXAMmYBxa82R8mGSes8
XRV05muD8GRm2bhfeaznAzQM/E6zn3Wa+biT6noZn093KPnsXqk8syCxuqitZi8G
QpQgHCarkJoL18pYitPaHCwFeAa9g75p9XQsb9DI+KfrbArPgFhw22S491+KU4r0
KqCZPQAo/F1LvzLQDGrE02zmxmxxTzWrS2eGt054D30dq/beDVLxR+G7oT3jRL/0
eQXtLMMDMUDjdmfuIa4ywH8GBLHOJR1oyYqxBZv76Oahj+93dS8myPf0TLxFjs0W
RfT4jDE587nzaZQ8iQE0SGTRf1qrD2rICLFSd6Qjd7wHVmdF5ux6uqsVmD9VOIHk
/lgejD6Vezax8DHgAkySr725hWKdvFEVCbJGY1AeZrdmq9KjsDNrCiTHe7dIgAnh
VwPumY4NuMqkYhXNMKXDntqGvMI0gQZ9ug2xpHnCoiI6WtOBs8vKrJlZZegxMIKz
C/PFhM5gwTu2lWvi8jNFaPjlgXdPwB4HbAJx0Onc2wDP5sxh/OCEDckKBZS6Yerr
aCHSBCto/Gp5Y1E9Nt1HlxyijVyOOzVcK/FV/vDDyyjledpJAwP3IELJY9azGbO3
oQHd+tgZ9cKwDiTNglUc0skm3zozGwGb7k+pgkKK3FnKvBkzI3fdYeUCJ8Ehhar1
KRhfTrwdKzyqCJYj2/SxQP1+6rig7NrKo2aKg66mFNzWgnMRK1p2WCLTBLswBCNo
f/1Q+0ODvhp/JD8BAAvuWG1RMx6MshsLcT8UySWoNaeUd4DwNPUVe4EdQbxho5cE
bmarBWllWDiSuRrCubfuCu8KZ1xy6SYtqZ5+ehK+lyxaQyD04Do5U5/AH12tN9dW
VyPVy7JjbUXbHsl4RO4zR2A6mF8mjtNIj5EOlBUy2hyZ65xU7sO2HW7k9k9rUAkv
2wWRrutnCK3+shwCEYMGA3GQNyoyKSRWx6rStw1wvqgIQpd+oA31fVnTH1yG64Fg
EVDOri7oBeNk8Z3jJHzC0YdFzRXyhmw9rW0CDyoe/foEthg/bPS1+r7Y0dDOr8vN
V/GxHml83tUDD6NQkgrYIpQNDtDc9flAHns8soYImRyGAAk1PpU0NqHsJA9UsfTE
NlmWWoFkFzoIxccgf57aKhjI0bnHsfPDCACN9l9XnVPSLAHo/8LOyOEeVVzQ7IEE
7c0BsOuYEdRWcx4s9e1rhS5YJencZ8YkAydoRpP9o2D4KWRtkDAnzuO+FsKN9u9e
eY36D6nVwxvBYoMOx/mdqzpfaf0Ira7Hr9Uc7FmSk35wTxvQH1e2jTaYIX976X/m
cDKwhOWdOzbQTLaWCKcx3GdegMLJCWUwSZPPiHAp1vKZWr2B6Ppawclqd7cEyt7A
cs4VOvo8kUYdX208y3WOYy2YCiZdPW8hC4mxt96NHIPS3GmoK5Phs957JC+R4pqK
0g2TBHHPRCY6Iwmcr8S4k/X82IaMzrwcGRbvU8tr+R3/VS0ad+bGG1HgtmUaVDY8
2MGEntR6BMotzTH4vyQuawCU3EQ3IBw9eRYR6wyeoMntWhXq4MjFl5VPX2z5PzfI
b5egZNSuyD6yk2Lm4H6plFOFdXvkVAH5hbUgivPTuiKWo1jzwNzJyq2zIbRazy5C
0BU0YVPNPDhyV26SwuXFitNgwRPWSQAxD+Vu9uqpIw4TsTVdquOSUjFYiavTMRL6
RHFEPggIEnacH3xCtaFT9f8BlXSguXfcOIaz6guH7CUJsSwNyBL+5eArCYxvdCTD
qiOK9RMKuwR/y6D2D4Ej68rnXCDjuYoj5lbgnTyTcZQv07xBrkmCgXlhV5F22cXs
z/2+1lc5zTXEhEsCF2UnVAInvgJOkh4oWCAjyv7TPT51TJBSdiJHcBPQ38adqCG1
SHNE9RnR0JoRzAdReSXFKhPCoRCQ0yVhN6baCpDHcSIGGrAV4kdIIOjbyvyjgN3y
woVZ2rrtqjFyyo8hOrmk2eWBLEsLpLjuskj35cC+PpW0EmAKrYUCWtz7/G4GDfPo
GoeJ1NwmMvrCuksi68JLASZL57pRDlswOMIwpv9S8VzL8QPvR+44r57bCCSUr0RT
JCH2bSa6jJ7c7XpqgCUVY28KkHdpch7FL9R4Hu2kwP9Ae4iAzWRluJXd7b+4e2Rp
0/xdIu9QcKDBYKzB1GmPKD3sb42P/uRG9umaWKES8SYhs4VcNHj+W/Pw5hRI9NYl
dBuKzbg97QFwFHaz+VAmOnoA8ORlLyruRLGrvJGsD19QcNRrAzkB0gcAX9srVXsh
63dUotej9IZp+eVkXSOF8OoMFjUpgEaawbFOqUosT9V65XWRTTO8r2nZNL5+Kkmz
jMoXKR4ro/AdxyO7ND/VFhZObtIZtI1rFd5sndjTtbPRWsE5MQ7e0Zska+PRP24g
9Qpznt8ADkoRLBTbwi51tvsV65aYAFDeA7D7kxhyqNKKXM/YIG8BxFdlPJQLw9py
AyUk1WPR8TDDd66aEVmNljaq8KO1U+GbfQvDfT35ymqOEv+4k0iUcXsLEmqZe9ZD
0tPrP52jWCUxu6nSs9hHommgpfTYkFoA3E9Sx2aolDSDR4/WagTeJJ4gBeOTABM4
qBP7rwN9yzZukZohByHamb2OqU8c/Pb8/W+fsJPxGYORw5bQhPNIg+s6M5xrTF8S
m+37x0sAetJOhAICFW0ttMiNlgzlSnXNgNL+pirlPQuJntm9fF/5lXqwxiY6S5nu
NN8QUOgL2DjKIjqsmoE2jaR13zf8xk/flJX+8T+9oQf3MqFL/6MAbJOU306cUJF0
CPVQVPuzZRQ2CIGlfScbxOtqa9yhMb8uNsC2frgG7Yg6oMvlEnSzXUVXLmnDiYJN
uqWLFg949w+gWcBEibrekEeg7DqreE1k7z03rfyQI+JK7AlZAFEiI/0Qiq0ORe39
6KmzEUok/uU1kvuFh+cEI9uCZJKm1MNq+haJjSNBBUQtvdXqXEWfZPQ7eTRYZqyn
0X5bv/OJ3+npC4mLoqYjZkd/gKzp0Q/h8ZlMQ4p2JBeVNwmYa/KDf0NlmawMUsUp
N0WlqTRak014zm29ZYHrUFB3eeYU6Ky2SEd8Tnt29demvsB0SfICsGqgzZVQ413E
5v1dwK7IRq60IG51nI27aCFM3MUil2Ui1vhSXqjAEOEmPBpIdM4U5zqbdl2prgqi
TC1eVc4aJZop+pSe4zHf66gwOYbQymk08fVSaCQEadBYxWSr199CKgZ3Y2JaU0Bs
R9bpJMwXBdXuH1vLQZ5lj4uw2ypZ/jSFTB1Xq4eWuuPc3Lz/XYmX876tnzF7B3C1
cv3wIbTHh3wFABNsMqMAWYSC564AtwMayFehar38NyjMbnnv3LpZxKbUUrPgfJml
5Usyy9osIq3Q6TTHOwidVnZ9fdGyi8NLcsMkEuUc47pG9WSKnXdicSKfcgEcraRq
H73wiyc/smO/9CP81oXykNc3+MlFm669Kz+UGQEbk4OzdEgmDD6lSnmlM9ahyRtB
nIHv7ejMODs9it2YEvkyBhaBL0qDV2OI0k2gUYpvi+5Yx1Esf2z5MIcov92+EXur
ONl67qyiro3ysBa8bck84L3KW89YnUx39ypTD5IO/tuR00KAzl8MT9vmfk6UKXxX
TqAHKxmxAPsTNfksOZ28wDLaHGMb1CHKzX0yGFMSB7QLlbVQtlRHaB6EiTGuoZ3g
TdGEZdCD9Mc78fk2Gm1GF4xuC7FEYtMd0hIG85CFcUUUn/VJZbj+zIuiEC/IHZv/
`pragma protect end_protected
