// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
f1IG3doeYrHavJrA91RfXEdm2F5Q7VyK36vSS/bk4sLMnW1HEKJbFMzCyTIKnv6f
A1qdgVBN+balwlimOuIhAauEWv4JIVI5tzfT6IYb1nu8O8+rM/4kw+hvOS1L72Na
JmEk7GNETOH1txMReDNE4Di4g4jwzq6lzI0k5yZoFJw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2368)
t9/Dwm/w/svMykLqSaqWMdGD1UDVeSTmWeYqKcbQgeEHqGuQ6tnJMhDJ71Emm0ok
+zZGiJw07TJbT5CwhH7ePN6N7Z9zZLKtW22T6OIEtLDyUeef3kqoptb/841I3fGz
JGIyA2jXH1yW28Br4JpHM94TqytPr9pgVZOpoI+DIXwjFOhPf6wMUX4mV6i71nIh
uQqi65sSze3rFpVU3e3lMoMhj/zqn+zz1VlwAtNKoaBAngF5/l6di4O4Pb7m9niR
eXl/8bfY5ToXxriyS/wh4F4ipW/T6qz7HD+egErn8eZvptYGm8nqSIFhyclPkdsN
giVHtk8P3+BKdA0fFKsujxUfjXK1oMBVc7Rt9K//D3rHchTr/4FIZnJzMuTWauR4
ng9VeCyHt7AC9bVpZgqBW1a2N8s/3Af8yaOf7RAwv6qXTYn6zoPXPsiZpURV7NOd
vkuXxh7GDyRc6uLu5+gBy0VECg+/K9y52z9ldiCgbVQ328yT73dBURkFp0JNTbIe
G1oPcOYLP1ss73FlDNEz8/xXprNeNURHWXgPnel8LIK5BpL5uh4PUeNRWxxV+x9f
XVl5d6igBBO+fLP7sVDclJ7mtt35euuwPdsK0gfAwpfikTJoDq5IYgaFHID0o8NJ
IJiJQd6xAe0lUBCIsF637StQO991ur/dlVwPUuswBIQi1ruMEwwQwvQIJTFDVB0p
eclEHtVmeZX/Cu+gvpPhyTOeJSbgJHJz6fGpklzwWBqhTTFM0yqRK3qUN97KlukV
FuQzjTCWE+d9DefAhQGMNBF5I6G+Z88u5H+Zas1aI4c2e5FtjKtP4A3jJp/M82JV
WjJxLBO1CutTgm8MoPZ7hibKjxnGASHOlSQ0CbLGM2FXQv3O4+4r3NSR4v2ht8uL
poEAOFjk9/VKiHQjgkV+bySIpuGWx2FpawEt/rXIet0AoNQH2O6j9CC1E3QjtYmz
6N5vmYCP18fC+F3QX85eeIuoBnOFwdUIQOrfrHzRNT+1lykyl2wolYznt6Cpvhzo
8eWbbezVC+B6jtugOtxKYkzKwuoWu9eJTEdh5d8NsTEnapIfB8n3Ll38rEphppaX
Ko2ILPk1ufAg37z0dZZe4vG/39xMala8KzM2Bh/AsheWo5chjZCDvDg4g6rEoML/
jrWWDClEN75KPQqH97t1u9/VLqpA/CPzCD6P3YZXEnCdo9mYLuiH10fzsI1JQp8k
jiibdutAgkb4RD3qG0uYmGPuquPw8jX54BwA39JWqxQoRwcWTYHlrAcyXXXEKjX7
9svE1XHblAXCob0ecGwGQitqrzjdlQvYbrjtkXP7OapEu7rTKdMEd348Q+64z5xe
9SviYdWhTSe9JqdEVLYzqkcPRjc5wv4ZTO7lnDhO6RBjYQSnTS2oA7irwPI/YHhS
RpYcEz8mpvwX+T47g4SPRf0Av9jr1JeOf3on6SUP4BxKWx0ND9BkaxPJprUV+hQk
OPLXHLNkhr5pfzjmBd8CEDVDhKEjtJTlFqHtadSVZoJKWq7e1I1kfRgJ3pXh1FyC
80mgm9Bl6cMfSzUHCQJLm43XWKq7Yp4IR4lfo+JD4vpJAxsVSe3L18Z3+O4XHbuY
r4BOrB8i+D4SST51SF1KZ+NffFtpKYnwLddGVvG/XzaWGYKCjLW1jyCFzLJoIUol
HJ2oywbKxJeY4PjkBIQ58QrIY5oeCccrL5g4C4lYdFWe8DpQOb0dvtPArk4DdaaO
bMWVvsLUrD4sLtC2pZkRxa+7W3lalpqq88bz0FBM/dB8LOsF9xVynhFH/jyuJFyJ
TKJ6xem67VpVPSO67LL6IJl2oOhj3IJSS+w4OkONxbsRCLozqKlOcHy/nZ6WKrk8
8yjpHQEYLhh1md1nj0hGxKjp2xKrqEHKga351sPCWvPbBBsLoeWwlCvJ51X6YUPT
cJd10U7unFSvtFA+EH5X44tyakKpEIpEuctfitY0xJUIPK8gAZ+k5geLwCtTtlW3
Zv6/yWj+GreSCv8XW44zBUKKCrfQNGRRZkDCdoYdpKd6C21sgmlRv/DOJgyZ2vv5
DuX68hXPZE+WPAt3pVAhvD6iPyoJRRZ47G95Uucs6wJ0jXZdiR5giyl5WgM5IdEr
8k/Y5/v5reTIWGgnYXDswJsRGf1UqNgKjkMNy6FqDsjpFIjfp3pX/eY7wG8pOkI+
eKyPrnsnmHIbazY95wLQi3Jd1j6TBv7nVIUu3TleO02wcNK+rD+v29lpjAus9ehN
oD+0iLVE7abSHomKXFQNS7CTNqLl5QoXWoN2fLKZtw5fvlwBeAMYXQE26uC1iPY5
A0x2W+EGpg3RIzBi3Qz1/KbxkTWCBpZkNiHSvbvD1lDmQAt6PE7QhR7PhBbgx5jX
ztXUh92LdeeiI29EptkEJRyP4hgMJGSwXuMad67MS45F4G86ixZ9+8FsL1XH4sBC
qfTkZVaFO+ZT/pe19jJYSPFZ8KpHhrbzwBExH5F83GygVuKL41LvZsy9ye671kLo
GcxobZje9SNhLyQxjlTJemclgNw4NqnGqmxI1LBbDpqKLN1DC7YYVgH1hadiq9zu
cGc+WHRT5yM/pCqXo2OjHfhWOmK8G+poru6zBhSDJ0HmbknIv1/p0uMmhFwEG3ni
faqde57HyUsuew5ofmPuJPagr19Hs+LiK2x8dUkhTOA7XlGFIbHvkr2MBmowX6tq
liOCgYbPHvOz6S7LcaE4jEJ5jFYjWyvC+WVPAYLjeqJs9r8q3848PkrMbFnWIiJV
cE8qWltO+KNsisf7/PPn+xZQ8pNubvQjbfEW2R4PguFC7A1fUfm0DiS/3oS8pzej
PF0bgaMzA8/kmzkKCbXZkCzNQZRmgg1mmKlGMHJe807kphtm8F6QMav2lUjXwAEx
/USgdd8docoKMW84heEEoR8z5DyjSoYexVZZeuEG5mqSWxu/ldQgtT8ptc04uqkt
P9GoTiSA3+4UPSMaSkW//HYtPahBlePSzGnUJ3uw7NY+QkLefHEuaPKWXw88xWgs
Yi8B7te5t88eumtUmIZrefz9bJBsmgxAwSh5JGUJwyOQUzMJWY3L45oq9Uwn671m
fRCHbWE3PzYjbvWB8Q4mlcCjeXR4LsX+GTrSD4AmUuP2+IofU0nrKim2jmGNg/KU
LG7VcvLi7kSTUdD7L8zHvw==
`pragma protect end_protected
