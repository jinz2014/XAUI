// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rlrbGLNoKqgJrvomhIaamTc0IX0dyaxzEzyMH0XUJcBwCkXKxwZI9cJeXE/K2r5S
RNbkpBrDLxB74V/zYOLHdOBggwbP599skUik1nHtPDq3cLUAHgBVxkmQoYyKobRp
/SeT5CebT778Fc4VrwZ1cHpH5bpfcesbWkQ9+XbeHtY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 258752)
4WMKU63OvMHBaBB/xfIFJwrjtyfbmo/X3XxxAIxifY9T/qeeGkRIx8n6Exqaakwv
sd83eSvY2+74f3BdaFPOytrPRVKcNQVQJUHXrusXJrlvrHVMgn8hkRnltniWftDy
9keDzKRaLOImKJg/EjrlYVJVu58SEHHZvMX0VXim1iBXL6EYVlvDYk/iPaiIF9Ja
Jx/KcBaiU/ExFh9MF/ydsG0C/4zrgmANdWqfVuDVU+cHdZvzwbfdEX3JoAhd5s4k
w8erptWe77ZSqfr8AL+Omo5LzwkmlaNTflT12CGJBGHpxFwBva7qxahvj8Kp2rPr
tjHlBbdJ/eKxAL6LqcekYijB4BoW/ShJBTfjtsU6pyPl6bcRnyFJcD8Fwnzw423B
m3UlEudkuO6j6xnfbB0rG2KM0emNFebWuE/8UagZV/mnJ6trWtqgUBnuALO8thLV
APl5RA7s1u1LBClYVNeMFpeESNUs4EuqluYSZG3xHu7074j1Fv07RijFnG1rHxSr
wsKFiOoamcg6t6YiGojPrd8C8t91ilabY/N13z0qxGbV8LApb0Ej89PDgNEbyoBj
tAwFgak4suBgc1o3Yv0McrbLUbUT5eqJw/gDg0GD+nbKLad3K9Vuotf3Xz8sG/qV
ec5t6Q3ThitBl6uSEDC8mKB0RDgVJ5GR+4D79tOWrNxQgpiAXVIlFC4wV6lzOjlE
zTEyewXamAMq3awy5chwAGUsqLHYIbAXzZk3olaambxDI8IrxAXSD5aO/PVyeMXm
Kr8Fk6GBnN5o73A1alOteoCVvsOKfpPEZFtRbVusmDN1hnp9XmdoxGF8g4EP26L3
9jmiVYPhlqdxEnkjprFnKQv5rV33RoVfCle7SRJG7FnzRa5RaOBnhCDl+PZmv3XY
AT1zksOKREmI+RUNjI5BpRbOB+0f4kWYHwUrHYeYFfdfzXcBt5Yea+4Z4GH36S6S
ke5ps87qadHOjiV0YXkx1sU7+saPNJr6w4HaQvWxJKf7QfY8L+pF9lx93U/X6xPQ
n7rbQPQiEVqffd6L5Q/s+9V/Qq9vCu1ztAEg62jE518YrjCj8olfjE2RKplrEksJ
2/dLd+o8ydWreCJMflRbinE8NoYL5HwAj9ZhNZjh78YH7WjweuWfXOqrur4IuN6C
piljdyym0qr6Bz5By5z1oDl1gdSSq/XpD7gg/C+yRIxy7vkqnitJOOz5huFIcjwV
fkjp8Dm8TZJUI8NfW+HNWhzFH3cH9g9ewqc078ASOKf/dCZ/dPkvFd8SBxUqq9Dj
bwHuFk+R6KZKzGQQH5Hj5nGdxnf4WZseKbG3uR4eb4ovpU8AnFB4BBBoRH9fQCcv
K+t62fAS1irk2lObWCegKqd2kjz+6C/38corXbuGfDCoLw/zH9JPPY9+1Glg25X+
+xuyIwie3OM1Dtk6ZBKoNcO8BK2M73c1zb8E+/2l3a+tqhMwHx58EM6ltycGgEA4
bbHKn9QN5oYMtjyThcUikS7+iWBCZBd5lorWKks4kuV+iXZBVy/d8yiEsw2YasGm
7ygBG8yV4jw3jDRrg8kLFedq00YE5HIS9zaq1Q5QOO1K7cxlEoKEdL/uVnkVw3Ld
Q+5cNjwFULhQAUSuoky62QkNg7A0VWi+6qAqdUP8c4F41pfj2bLfovtBLvJzMeQJ
rdUPYiCC41CbEM56nEF4NOdaFwtG4RdS7JXKK8S8fmYjd471aWujNHzXqmcMIQ+m
UBAC6apb4cpsdQRG5aQCUpi9y5wKC7PwFHUsY0kZsip7dXw8bvrxvG0TXZGc4q9O
DdUNtQBkoTCClwfR4O8nx+gsgQR9L4u8hKn1XBxIuAoAS1CXZlSbeSM/fYB24XPn
k0B5iLIsWYsSho7T5HY1b++2sMb8lMO7YpptBXRVW5kBUV3kGcDiZGgq5vfmVTBx
r2OODgzQQItSenmfFzfr9Sb09LR76RLZXV0u+mjIysWwlUkB9Qb//6lMnrlIWQ70
xAYxS7hRhXjfWFkG1A/wg1KJTM1Ia6ce+lG9c3V9YXiXQ5Kt3GOVx3N/NQjMhJO6
yD1NCkaPyooKUp+j4wBu3SUM1ni4EP4CgWYso8TLt/Z8inz4eZ5Ynx6nekX6H+rN
q83Kfix5MXHSIfQbwk2Ybo8/+lQvr26xzHvH+rVjn1qFnR0aoyJti07DvXKmPILe
EKw8JaMNgUCKaq0+KR3ajPslZ++Ztj0JhWeqqiss9ib2lRnMmxLkxO4K54I4hbd5
U36uWmYzR7WEHwERfk5SoVzFkJ9RohDWebXhfZmheXCIaao41PJP/icJmoQxz2nN
5jwnYe4omD8Ob0iAC624JtNjoRuUyEJN5cZYrA619vZhCJL2d9JrN8S9wTgmGqWR
nCfZGQEjoHwzFRW1//FSMpwujbBIRiMi+rif6Rme4RK8BGpV/FQzcDfRFrawQqVi
4fDNQLUYQ4gWENs17nxQYEgbxr+pNlbE5gmGxbSOAJx8jdTTTY3ebWv+PudWwNaf
Y/+2Cu04dBpff+RWP8BAd1OKPRi/kf3TsegSP1rrt35c2rg9hPLeH4OHJzEVlukd
5BrJY/7rLnrNdAA2kQtVsg9UYzBDFS4lzLXvSvMq2ItIgWqFu6BrMkPRjfAa72AJ
L7WNq1+FoNWd0l3DJQ0obstIMFSquvoAA9/A33n6r06O3AG7US8jkJodjC1DrtK3
G1Hkehej7kwNNS0AItHo1xzHTR6fjpGX0a3jMsAAr5C2F/J2P1slujhhkBp/wU4b
zLifzqBmWTMC1FT91kGF81kxvbn8r/N3kELzZ+9s3MEMee3LO0OlWX+/m06K5qsD
aR4WI6uNnE8ddURQpf2GfyN7O2fdFr2GijakrElBqNZXCvaGYfz2F73CxPwxo/GZ
khvvj3iD6LfyMM98RJrr+x5d0VUalBo376+i7Jo2cXzZNqdBZ1r/W0lbjxnvk2h7
cKeFQYRKj9bQrUzj4mgRcHcW4coMGQhamuEJ+SfWaRESXPssI5KmV4fT79IzvSaQ
Ztc7SGKqYZjB1wX/WGcyzVtAcrPk+WOtOefUASEooKX4z5e3d5or7JHL9UlhRy/e
mxhO3jPquauUXMaiiEBMQZC7D4ssU+9eC/cBaDhL1gKySMqRIrwzKGMd7rSZJw5M
RIvWgoGwl6VaUX83pgizazRXazIIgmVOlF+h6rl/FKeLKbVY20LNg8GIRMaHHlA0
BemD8J6Ob+jHzbqfeVfM+sRKV1xLL4y7AxdpHkGX0RN78CJGOZvidAvW1yy6Pl9V
Xck1b5URs2gO9ut+wjFp6GfkVMO+zlPQw1JM6ojhNUIQ88qsx+KoUKSgXMB5HJAE
MTuAN5NUhkGyP3+n22b63+oiJKg9pOGnoYZWkrTWxNSfeLQ11a88pu2eUyKxE2Fn
9kF1pdGzJwzU51IEcvMfHQUZ3dxhljcZ6SeXftV5ktIUWC03/L3upjIry3wPX3ih
LzLbCGIh02JCBL9Vy8wfFnLUEsBvkfXCdmvfXi8eVtY/izWEKfKEJu//iykaFW9t
XTxVx5LthMf3sfgjSJigdN1iRJEZSq9Z1AGgC50K4/Nt8mxO7G5al9QFGx79IDE4
equ+ubvVw0Z3mPXPlrK8T3qK3cNIpL7GZwKt//jQT/ryhqg8dHQBYINrIRg3OdqX
YwGhwlbERvncJxbnwhIR+E/ZiG6NTfqum4y/nliCaGQXak9qsXWdUfejQAh24yt/
b7LEJ+izISix5+aTQtIUZYuzOt3kcgB+TqxrU7+XjDPzfEK+zGoJYGoo0oqy7Dhm
9mnJpE2/kigfO9mgh7YF4CX8qLewdLjndQ3VWpOaFgSE5U53IJXuZVXzJV8P5zyN
0nhPLACgA2nShURLWumrYQcsKnc4EkAEKwm+FHYJ/q7ZZc54puSW6QsngBACGouu
ourlAZvyNZ2ljKTQEydcaQnPLRczrjG0kJ3u53eczD7Y8IPAGjz003zecYKmd50J
emo659FNjDNhOHTfHooYm77H9hmchDpTxnCg7cWseLWceVS+72Qejya3nqESOp7O
ouYA/PMrVuGhNXfebDcILONFzsmMdKWC+rrdXjcsELCpO4ZUnxaTuC60psudC8Zb
icP4hpv/l7gf3b5Cikz0EJBOswP7/09POoGkxMDY69e+oBswEYV7waIQILX4VeKo
2Aaz9BEzkgBjUvMedAlDTpdsdE800G9tUAZf4RqlVm6bt3NkrnaUXUq9ona1ADt+
5y6ztvcBhkN3YGA9Cy7x2N2MAawmTMYwzt9cFUq9RTAXNSWHKTdo4N0sdshrgsfO
ikri8CJI17V20TCQB+c5CXN7qQKapNBtlX+6irsLgNFE+fVsWHlAUZ5tXaBNUBdk
jG3MXXSONyixNU73Z5diZl2/EnuBvgIu0PB2A9GklI2pTBoWtHbjW2cz3jX3pWrW
btGa+WJA91qUryYV5KRUgvSDoEANHvrqt3O1+yK3ooyqPyUY1wjf6YyF1ejjS3pU
FYkbaXvmpyarQcNTryvYKUNvBAgklwKNNBpaOBSK1N/aPtEI8GNHhyVyB9yVgTYF
+GRbvNMIBQ+GL6I+Aa0rOilcnqZQHx6MudURHm5r6bQYp2F/ZbNdYieOehzN3H/A
MF91mvTCCxW2o0UGFrc9T3kh3ceDJlhRI6h5uWNFL7R5UVA1Q+eEtk6Tli8sqeN/
MihRwUb7GHvSco4mgbZIZZPHLjeRH+++GkKUl87iT+ZDbwjUmU5SFNPnzgF1YbOA
tethuFc++822OyMnI/4fbgQiXR475h/85QtmGFWSICQYTLq/NGKqALpLObOsEazu
J7KVCuM2wEN83kUlXet5EjnFY3bDjw4yi2GhMAvlmBr/EKaARrX17LK0epEttp/a
tH00XZ1LO9Mrx6SZ1K75xTvM4rNWnFe40c2mw7i+hM/ZvRbSIo7eUEBA33Z9LHAb
G6Y/y8+c4jyRpyeqjsQ4LVDV8Q4rVF/jsAOyc/hiKrIv/o9uemZwXJUwRous0I5w
iqqDkSg8QclFfU3bUGBzFicPWw/o4d3IcwWuilNGfBbzBZBz5oSnVKv8PowrTDtP
IhY7aXjRsBFHgCDOmYcqIPAQYdAlVMzTcY8OA9ZH6ENP0gjz4pz7uZcdYw4YonSL
5TBVesOjCOXShmMmKnZFIIWbazLg6tV+u5x6nyx0gEZTWDnif3wZx9v9aWCR1XfD
BNQn0CUGPWaY8B/zixLxLODNob/qRH4OZVNzUEoo1WW/mXW/R19pzunbe3uR3vx2
PgwFblkTL75ynP48zq1xQOpMu8Z2X956UkBkv/YGZX6VPR3i5w0UXyyb36hQhRoy
Z9s6RGfB5NiSKX2xQte+HkV9vESDtsmcovUesPlEt2WrcIdC6zuU98WTAqA3T3jB
KVmCWATIZZlHktYReXNr/Ti+29VM83dJmBLbfWGkiTQxGFazfKYFVraycRDtXiAD
zl5uejWUYYCwqfm8fFfmUtwZqAEANT8IhQE11+/ZsDmq58ogywFze/FFm0s4qma8
cid1BiMnKIT4QccSTmOZEjDW1hdUHGXXKk5Vcn9w2Z8ovfk/BPsjrOWn0i4AYjZg
ixXsOzW6Jy7qcfnBZZHCXH/MLXEZ66Jk913cDdaFDhv0nZTeiirbpaOWZ7rKxc6i
ArvvTYaICwFgz2MkpTkpbKXfDWV5Gt/6cYxzyxOUXHIIzENJ4F4UcD3BcrBJdUZU
PtWmQlBrO/GAdSEI9syuXODQyuqCuMa92Ditl9Qbcks195YLk/YfF9yiDw6wlqny
njxCvXupP9EJ0ZX5UAL5rO+B8zsy9zWL1tG44Ft2vXd3PekBWU7Y+iSGrHyLdSlV
fUOrp29k5nZpuP26Bks4rUhXClREz8tYD3HpQkUR+2RaPmioq8MBtQTBPIRmaQk4
I18MjjhxS/CqPXClv5zrMQYtdOzEJtG0tEhSu6eAywMcTXZ0p8yMMzK6mkOS7FFa
EouwI3wRF14WjQMALSFD4xsw6gz6goCiMaOIdnLeibkyOAd3nC6GRimAOga6paZj
oLGJuqxvfEpDUi4Vd821IC08PNeImjwZesBh8XnuJSPQR6p9mrcCHOx+oNid92nc
hqSzjyyplV3+VzNl3YkLXJjXnYLM6SYynGNUriukzm9XJ5INWSPm0nnyo3Z065qS
4GYN+iwyuGFWsoo2e+xuv6AHL/COOQ8PBLy12CvFUnzFuqQ9tkByL4233aSie5vs
JXwW5Tc5oWjuEeudf88dDCjhk+5uO1xoElkGuG/1R/TV0S7J1k2Re4mjMF5AXzEA
T3DB941M4tWPS0HwM1xgHN6LOMWwp1aLR0bk+TqFJaKAfbiXI9rueEVdjDwDnrxs
4ZbGfxDG93yvuLm9ZrDgWBCtpHpTvJmElcw0ENGxGSKNdbodi4ms3kGDQwxqYw/m
5AG0zzuuNJwlyOsEcDVM5/wADc7YGZdiAe6vDhgdwMqglN+ir3mKQEsmj59VB7mO
pSHFFxQIGVWhtfGxgfQPBSZjixJWv0IuCICYzm95sVw2TndLYoJi9Xcg4l5eyys5
FjhaiRt7km8iXa6lGm1WhKAe1MsjpwK+2iXlJ9AKssalrc66teK6+jHd8ox4pWw6
8DT/XbWDsKJ3P+TajGjb7/nfgZVkdqmQURVfv7K37T/k3//T1avnLl16FFHs0qjR
kO7/bohhbd1JlpKpknJWgJlJApq8U1ZIIpwO2ei7pjVNO+0KdVjQ1dFfLLNo3AZI
LyPQOABDsL4TrN3joUtj0JcvzEh1wFb2U+vZhExczVWQEXY4epn4sek9GVaJeiel
JgTCaasAXKwi5HTxQ7VCjNncktcXHjyUd5banWQ4+YmtUaa6YnRuGpri/2JCjMG6
Bsh1ek0zHHKtW4zEDUrrIdlLYsR/PwjIAfmno9ESJ8EkjF/TpJji97m4PvlieHca
O00Vnlr1nOWetxheoFCqY0kY7087SjlWWl+7eiTQ0fIqrNz2bxAN5lIeMoFozHkM
SoR1nHjrDzm+njyimKr9LPkeYwbjvHhFgDKOMzuYpORdeuKEkA3DX6XOvneLQKr8
Ycy3/PSjtnRxvqJHmIbrrPKZbHt7gc34x8dwI6r0wyDaCuh3A6yc3GBMm4R2J3xv
ZG+7GyEbNipoBwSmxbQz2U2Rl75QZE4kVqiwTsbcgjih7xAfoEtLD+l1bMir9ysO
c9RMvLvvL5ITBnddWTz/TikhRVUqh3b2K+sg6a+0yMeVkqJOkj7Q9CD/J27g5rxx
+g+WBWKI3qN+JYSwkQ1w8cJX9Wk0E78/A0tg5WB8WfFCtfsh2lmVGH08QQsqNdgH
cAqZh5AYIOpIkARTg+m25SArQQHRRHw8Y50RWYftULaxmaiEH3Io/P/z/rb/AUYP
7bf+a9H2r9c4lE4gNdDLmCn0OmNnWH8G8+u6e0B6gXQrKvB/EMy2xEhGrCUwkGKb
+nyG2WsOPsydFLRFIgkO8xRABe1Ajs9HwtXLMQG0NL13lfMsN50dSOgoICuhrfTQ
dK0maute+z3zDkps4/YG8YGGkwj3Czz9OFCYTRoFnOOBWFlY7xRhYSAnDydqXrsp
GYgqlxCIQxePR2c1Q87Kn6JB3PJ089diu8EEMwYZZxMQfWf+loKyV0o7C7/2/8iY
AVHDhWGLKIoK4LJ0n03xOagfV6m+IFOcK1GosrSy1J4IWzmEkIlx8JUf1VBnSYEF
MHUq+DwFkYfbAWwsy2Ohrr0O8rCo3lyvzdNophF+Vm08XbX3ps3jL+5PtPLpXFf/
+d60KbaeWSDqldotk5yVttp5HjfIWoIRGzF97nq5vFRce1EiZOlbPtjid4R6S+gr
yu0qzOLH82EnWNzH+t10GUHOozzDPNiibY9JZD/v9ClxeSDrBOPyC71+y5z5U3JZ
x8BTZyHNOzPX824P/rWDm8CQR12VKghXvwX0+fh+tFOqLKvZ5OTWjtqo2PapMG1A
Ol8wIzL0h4JgZtMsPJL2Bnt2cUlp357vTwoT5XNanh24PIu7Zal7Jkm3DZ6u3Qmv
OTG3Pbfq93vYnaZ3X42ngX0EiubPMY7waQQSVgeJiFpWKxK9ueiLy9cbrWXijj7W
BT3uCrTg9R6h/PWonmMufhendXHriivgmhr1bvPTCvlDMhlx0TSdP1vds+AZCHJY
4zwLSHHKAYCpwPI8hOA9QKzG3uRasGeWIrL+7ifz0a+0ybqtTYxs43Bax+8bZoY8
ajeAIRBJd8k2+GTs3hft+IovkGjYw3IT3sGnQK2nRVoiJJXjSFPrVjw1E4ndLtkV
Rc1HPI7yloFctXXAGZX6FgbxJ2vlUT6cyFsmJalO4gdpH6mYCCEG/S1oOMx92npJ
KvDEA3ZpcS8Pm7+9fAq/rlAr6uLBn4Yio9V29e7/o82Y9zWDh0K3ARZuBg3bGQ7k
qF8gtGnukyFhUzH9GE97UfYMRkIqd75hvxk6s4j+qpJ7QhUd9pz4mH7+LqhInjQ8
QhOE0z9NrdVWaAE8mItDN7qVJ1rXn9yBPpQCusDiThfuwT1D88HGlDktv3w7znCX
jIsDXmCltMpL5I9bxFGwN7OosLhdwpOH2lAmaEmBYcnKjvc5WOk7UNgTieLvDRGH
hmrK2yrR8yPrw/Qb4+yHFWLdkxzTOLj3STw5ABLuCGnPAmhDwIpsWaab5mB4eX1u
G10Is/ytWF4IuqvwghNuSwYdPIyY4lnk/G2kK7sGYDaLrpvqv/yGrxGaF6yRJDyK
F4QrRtTAedY/Y8cjRoIlsw/Yjn6f9p3q8eeeJi7EqlxQVaYAnZRn3zMgZH3O7X5k
P9kq2eDPMpYuLnqmjk0MFxUdSDV+Mf8poLE4vkj7PEQ4LFFEb4gnmFivrYlq+p/n
6vvtAfnj67Z4bkzmezzc/K+Ncd43UEy0B2+cEQvPgyGqo5ahMci07sdCkIXd8ZbE
57gE4v20vUIKPMqp4F3uovFh9t4vo9j6B7/gI6YRpqp/XogwCYa8viPnIO/dXrHX
brIVllUHsyhiS78J2vqPeOIdYJWVHdiJj0ayZkcioKNEknf0S9mQ/h7K39RBiP8q
Oeomm0P8yvAejh/tonPyHFOlRikrGwe6tEdDS9eIIXkik2c6eNPiGJlCFGQ2Qh8q
pPlKVmYrbBnSdrjngqid9I7B+0gF0VTZMgGZZ7TXaVZ9QM2CR0sKFUxCt2GwnXsu
SeH6xTnY4ZpyuFG2megUCM2H8uTP3ow+B5zimZ7GQroAA0ospdd33PfJJS1KtIWH
iRjBrpxSvEXqaOQ/9/gZFrUSghxnY7B3lXlwsvjGwPN32/KAU32MPqQve6WSvaCn
oc79Hz/PxiMNCr7EXyP0haTjBnE9e7uBCubHxmU72Aaz9ovPzH3WpQC4BuPYNN5B
ZJGWggJdrAPDUaE87/Ujd+lGwscGgLa6SH1LPbCydLd/W/Zy8PEuO4vlGPwY2qwo
y3LAyTbORZKwv0jkvdtiJYrGzBEtayIQN/Xl3hwILcUiQ7kO1TUpTWIjVGS3GE6v
KzHgeWq6X98zD7b0b+w14gpRVr0QYAeS4Or1qdQYbrJdf8vjMmt4ju6qXWSpcWqe
gSzVyj5G/MLjiH6otrmwawC5pBVpsXEg0FYJy2/8xlPBA3g5FsTL43H01qpNRhHS
UkRJAaRZOjsnTFjtlmOAf3j7ma6PhfdsgXIGatb/A6isU7B59nFA62bdURk8ZKo6
kOP9rIrYyxhJAjhzHS5Ut2xJ4ykhVia6W8KEvHoBNPWFN6NOwUUmD9YA1NdhsWwA
6WAy2KvZClxRM9Tmpb80VGKdUeyyo2RmxqGpSoLcF9ErAqsCENq+FPu5yYPhPJkJ
H5iOs274TCKsqjAlvHtyKnmTvc5QrCBpgRF4rLOsx2gNKuR12fyksL7sk4i/l2y4
wSHssAXsMkSwrg6biLmu0jm6j23p/qmTxR6l6sGILHT4T/jBHbt7O8eUS7ngEoDj
LfcrtqKn85ZQWu+xRR1DKdbWrFJVcFHHLkywxO47c9SIL0HrVwsULfNuLlSP/SpM
HcBOC7bzxJXe+82P98Tpk5mH3P1BV23FCI6zp3w7wnCu0Druy5/YoH/MsICNScRT
D/pQmLnHbjtQxeGxH/4Iwu6sryZdlYOcMzqcpmtpAMI/crFB4SdZ4E0O/CapaWwR
XeGeb5wbQ/xWDmB4OlsTGZmWJZO0RT8SdMcjDw3pdy9QamZz8dUAnYe3zcspmuAU
ZKeQNfhcKupfypopMB6qn9IDsyISmg60ZieeF2KMW4KOubZ7nAP1ca27IuJ0fuxx
mJ0BlECVUAUisYQEiol39QwJOdE0SLohZELxIS6f9cHhWpjBxY9ACtNpfUxVVS+y
R+YrUEJ7gB+vSlHwL6HTNa0waoD+5PspLG5/LkmQB60NbqXnLdkDH+R2jANWD4q1
jELO7OrYTwz3W2QSU540/BM5MExcqqR1wytqEdw5ltNb2xRRqxUpedfkymmmaK5j
5SpUdPmwRyE9mfOXS1qRt6QWAq/tD6n0mv3Ccf9L4kdgk/wVFxCFcv72V2tfuN+v
zN0hI8X6Ex96IjtQYtiWm4BGcm30D3C9QKO/HWBeJ9pRJqLc1C64BQTO33fuXwgR
tLKMptI74UpgevvAGAL+pHLXMeO8yVvYB/Qo64gPXn6dD/x3zhdJdMsOrhozpj6A
rCbRncq9mnkIZMxOJDfaKAvP8HERaOWpl+emshwv/pgRbiidKFd5LH1Jg9bKDlLQ
8NGFQl6lJ3GsPYL1PsjBKoHXPBwJleM9o+LFpW6hDJJY1sURvy3mhxutb/NOOui8
ZHtJSkDF6KEQLIXtkEoKXr1PJYAJP3c19t//Scki9tPmWWT0dwVU6qf7mKzSVPQt
F/rtOzGJSh/hfOlNZfcEGuoVPfpuYQf2DXF7zKzku7qWesfP537ssS8gAD7JSCCk
+Y7eHMXFppskNjmGrcJtcfAhaxvfvbjl7UrrOBSYpWPCA18BnMMcs1o51Y4AUhAZ
EiUoCGNbYhILKi5hbNMP+S16Axk6ZlbxsuSKSi30o0BEe1UGy1XudVCgIcFV5u7A
iYSKQlnZfQR6CXEm6mGuJyzAapJvmqJHESGP9PWcsYv/KeMTb80+4V1bWBQIxS6G
ji5ErcI77O63z09ZSCQDTlAEJUowz3IbxJt28y7/+CaxsOsHcdbdgEErxX9IChE0
R3vBngNkbQNHGD8ndtPwoaxTREedcpgdRhCPLrmMzf2JF5kC3rZM/IleIiSeVXT9
UrAcJG9OGryg/Fqy4xtmDA2rGfOxkp3g4U/TjeVwMhtVMRKZ2dPyG4aG01f6++yE
PNIlsU1Ct0KRmkATGFZjwqiS7M1XD28yTsK6TBFa9P8BzzLHqY/SUTTrLVAfNlQN
nmqpX+brdg/mMxrwmhSDykZUw+aawPaVr3nCyvZ4YeMg44mRt8Vsmt7sj+dvBQZd
diiOOIThgpYtow45P1RtiaKTgrN7swQoGKCK5k6f53K3/vBiBjxsd0bQVaBw3V3h
lGKgJBXP5mA6UQ2zxlpmqaaJthvdmmCGPHFGqNYTwkDmG783o1RluDJQGvAo90Gk
i1kAlmpjZ4HrvXhFiim2v1yQxpUTN8My11GRlZfqNbGeoGsyyhE2W6ANVBl9yPuo
EQKGMAMP0MofOsWfmSkUDiU6fta0H/0qrpkcsI/Oabb7QwAPGanhG5g9jScMNTSQ
dmM3YhyrRcko7ANy/bF6rWbSEoY5P5bn1/OmBB760H/Cpz0kaACakl3QqRUQdi1Z
T0qGByYM40e1u9p9I0MaYyTHCZsQUQkNSxTkHOIyNQ8LhdeTDCHDHnt4rs76sBtD
948SCpMNjQ3nDV0DvH5xC25XIykHKGe2YhADQKfL35bkscydQhEpiBKTjnuahzO3
lsN6kKcELCJcetzqj4TYZGN80q6Js8PzuqINpbWWLwyptZBcIk9PikKYuXv3JmmA
X+sxVzpxYHeatTlI743Z83XSnA3c9cJ1uubgBh5elRoLGOQMsbD/jirxmxMXt6ki
cszoGdRjn70YRslXuWTY3kyQI6XUPvE+s9Ifu6jVao031XHSSOY2ncKY4dEE01Z4
FPtSDI4Ya8fvVmm6ME2wmgFQeg88bW9Bwib3vCO9YFormo7OvKFqE+N3VmZDOh4c
ONsrQrpghHLT/wQtyApG4Z2SXXetZHKaPDEljhE8RqiHM3tIhkTQNqQddwlS+9e4
nWIDDhWxrASYix/foO1W0SA99KJPBY5sO1pzmCc7qtk6TtO4b+RA9h5FLs7mp0A2
58wAP/Mrl2qvCHZ+FxdFQevP7QaFwggubPfWK+UwSeWG2IV7wOsP5tXwiOcjw79O
s8p6rnjS8icSzvvTXjyUoB6zdKKyqxsR7UOrzC3qgK47cEwb67YpyBZAJkw6woN0
LX0IIIPy/2p2hzSr4Q8O05fNbGVKa+xK0IWx8qKGqnctA+leTmdNI2gme2JomKJ5
BBiWX6Cuj95SRtUiJs3MufVQnJhZsiR9uBnrQfCebLSkgw01OViKTLHlpV4TR48e
olUniZ/sTG2XprfNFfm6b7i0/0pPhX50ovXT9sEoXsqTSKQIpIGVl86/XF6h2+Kw
HI36AwBqhBKOs5R2KB7wIdEpaHV8cRhozN5I+8bD1SQ+/oj69q3Cm6+iCeF0Jdf2
4eVkWF1Oyss8D44YuItYpD8Py9F4wuWNb4ExRSAPibL2WSNQwffmW+RvVi+nMQtW
S8vAuK/JWHdxwxFbwMb7+twgW6HV85fisvN/H8XwpIkHF7brKInx9buKkVXnlpHb
95XodtLDpFhDrnkREjzbP84ANdafR4U5bsq4cE+hTawuRGAuffP5zyE115nwzPCg
z5hb7sVvfQSBfPLzZuqFB2pU6ATKyM2hg3WlWww+DgG6azRVOypkSBU0qgQNYh7t
QbKvu/8rPzsAlAQAudxUMePlbWL2uPkImKnXlC74IrUA9s325BejeO4LKMVhyCbC
p+9DKtw5gtinanpCipx2dfttMEMkB8oajZNqAoWo/zrQE6rY2y8HQJTtDUE7ALbM
Y+Om6BTyxlV8KEB6I85xB+o/p+EAt3jjwMuL1OEgULfnpelDAFtKnHfDggBCvDUx
nn2drZs/R442qPMPAvEtr8PJyLmqzHGCkVcQDc+XSjjkfJC+EPRfnqGL8SF0wWHY
Ca4EPwkSuZPGziFTMp18ONQxivotF7QoIn0YN2q0Z7/POp4VVh+8GwVIV7E5YDvc
ftpUstctrw1HXBbLAZmFqsFErAQuSI0ZCpdf9SJroRWsDKV+r4AFA9s3u5iHjlS9
GQyCCsgN1TBEgQ2seiHUWKGZAHtb6UHGWlSwjwW3drxT/vjZsnrmDcwFzE+ole++
cIWTuF8sjExmNgkUpqkstFhh0wp7OivhZeQti5BcCQWbynfg7MbMoGMGWyTJXT8Y
zksueD55xOZL9bKUFDWiffVyxs33oJD42SRR/Gfl65mRZvp4i4O5Kf7uEV4tF/Tk
im+3k6fqYf70N064V62Yq65aZnsJWYzlTBaJvFAK3NMQJwYh+pWrItcAmI047eQO
ji936uVJ0Malhcb1Cq22P+exids1qMqTE8XVAAYRqiYUWY0QF/8b6Qx5qEkw17ut
ngERVcXbE+QSCi+vi7tgsnn3McAi5wdVJbYQWP25aU90RbQBD5U/NqEjzXSOzP+I
6UOwalC6L7RF7DlNSXF5NNCo7u8iI7DO66rQmJJ/Av07PowFPYyHmsoZGfTujkwq
aPQnfUvWIyzIVOMk4BjPimM6tKJHKpyfyQfeRdfCJvXfk1X2RGE5l7uNZUJ3g+7m
476zjECMYpAtGrIqv7VMRfnt3JLwxosxvZmQWOGETKBgB8M1vY4Ok4tu/SFRupK4
ERLeCMRaQrRgKKHZu5f7lbv61YlVz1HpaL0LKX4TO+3Robf9xDwBQIPu5iUDRBAv
ieBx9qXJGhhpQl6CgWmSNAyWzN0pkVXnD6/DJ++gJga6HhN07bi0Eau6r5js9i1P
2UN+0J5OAl2c8gWDwot9/XgOt/2cSv00X2aBRyIiS9YT6P9u/6DwL11S3/646ria
hKZSH/elv/4F6+mC35q2BFZqrCmbdNJ1K9TCALBnZkb7ooo0GxDwXA6XiZIxpt46
o0z/rzKqPAinfEY5zJRngHcmTAmzH64F4v+Owkpk2lW9topxutk3GrMJffv2OtBH
nPgSFWpW+j2DVocd6bl9cTKGcj2cfjmBmOdmZB7F+B/HWFnTju6mMy30BPklq6KQ
htOtofqHdS8Lu/S6X4iKWpOQvk7u/KyXWeHYVVZUzkUeelJFbnOAXNAHO68+24R/
iOcnOGppM6BNG4QwvJr/1FvN8fHkLI3+zKtJIpRAP8opQ8AXBgtoPtkEHxZvRuoK
D8Rb1rKveVTMhzHgSE/4gGMh8RieREbnaJRJzyIVRIPttrEMU77K7RHsLEwyEwVC
r0ekWmAqwMdGGucoDC13aJB5z1GzPpuJ9MnnXZmkJO9BiQXWv80Co1OJ+8gJUntr
7+Z/o4w8+p4JgoifyXTiQs0c/2aZsanipVuQQNnecJfBXttQWIfUSJiWGOc9tsx8
bb8XP+wYqnUKCWEwH+rK4qovcEYB1kklWnzy+a9D72djA3zgfPuCJy8TaMMzRH/Y
h395HdM8hDMf4EzFziqpo8feMi+uk6Ko+o6BgAChv1W27Anx58PWjJrxZslVdHd1
onZ6a3bzeQhXWpVFSH19n9aHdQigYTlDBBoaV04WUBO2wKyGiUGB9wPL5Yzc4la/
X+oH501ZeEqKfmdJ7L2S9CoqAMayQ9A+n94FHFGSf7w/FG2o86Pd+F7k8B4gYpRS
iaQnUSy/KgF8S9fWZMvc01bCPtJFFvcjq8sLOybFkpzqGtabZR2b5PgzjIHIEWrh
BBtLiopBYtjZWdF2SEXQD01QYT8lcIHb1Neiy9fNeuMUBtz/jjfBBKVTA4J9FQN+
EP4WaXcEojJLTni3nHs+O/EWmedCnqeTNw/Kc4FZ68Z6Ls1cpNO47zqaU84gH0aL
Kb3Zfm6DGqoajxtaQs5xPn6xmePFxnIZEkPrgEsTXHW896+hjsiW3A6dRqOu++sE
PUFnBr3YoW+g1YByM8NkCl9M3Yx3HXzYo61HGOpadGkq4gsv8hF6HRuW/RkAP9wJ
90Eg+j1in393/V5o5tI9igSn82LwsgeIL5BsiQ7gOfFtGN1cPcm6K0yMC/YQwhvc
oQp5oslQIR7oOHoI5wfcfvS9GQhTYQwsWiDKERXdVVblDbY6cfwyZbKtWakjJSgn
2IaVyMVY6KGAaPIZZj1C+rQZ4xuOn7XQGoEbeSBwsFC1xksYfUi2ibRJA9mA1kX9
Smd/j7DYvc+I7AsjAa2xo2yW5fUBs9dMxpzbgkZaYZSkiBACqI+BNaghUwTaEr9U
rP4GoHd7dciQ4SKJzd50w8aGVXxKL1Q5NEZWZjk4KMSVJO6ekseyn/ZyGLE1xya4
9Gr4p88hjpm2g3LguMms0hcLt8TUZ+x1HUFtWbHJe8GNbDjjmpDzeWNjqC82NfFL
ip2Ffs27qMOaut0SB8ejz3JHoqjqbqXp9BiV+yOmjglbWxPQ+B9QVQyd8CsyeY89
xOpdqGJBkyuh9FCfKqKHK3wG9eWyDfSxa16VUtj+ajPMibSy6uCcvw3nJHznDTw9
BjQliCPLzQC/3ugdgmSgyvxRNkGUlJRmu4AvQXdbrFm8azLIe5VduYmN2dW73Koc
dBFAyvBsOgPhMtz/AKZkrauLafy/ZFLl2qiDtFyNFmsKpb+BZ8xH/XygPRAzT3ou
AyXsj6ERmn5LctT9K+v81vLKi0YKbXaNwH47lPNhMq35u6o1MRMjlaqB8w1kKoKv
TjjW5EKRwOzxY8RJq1XEUgZpCgNThqjDlZ1ZXxMEnvJWIzO4LdZy+h9tq7xxQSqK
b7CsAr27Nz8bAHPivPwaRmwL+v43n3turQodnZ8HGPP7924zcmfINRrNVvEFM6G3
iWDKSjnmoHcEQLNUuFmjUj9+V16DD0doooZxTdmhF3uOaNenzmQ+1GMIWsaSnZ3n
KpdRbcVpyU/S19Tao/vn0TMdXJNOIHeMdVZd4xo3BHbCJGsWAi03gd8yZm/OsjDq
PnTvJ3e2oTJJPm2GXqusNYyfRJYXutEh6kHVsMY+P7ZvDoL1J3VCHd+guuf7C1rE
OYrE3IrEzxrNys7drA05ilqOZXkenuCd4Z2ogBg3NHwRRpOwWjjVlkpgnyyW7odr
J9hX/AIF1Ry5np9MSBGvjyli0vyLABgKS44ibGKw4XXNZvwBGigafacUmT3IUgcq
aFLUD7nKdtlEncF2A3xsv0O42hWiZf9uAZXBbVVGG02QzQyzPMA7QqGdPAeY+TAm
t/mkWxkBH6uPZ/rnxsYoEsBRccpGul1E56GC79H3GRprrWkVDukspzzpinNVbGOR
VlgpDcmshF/RJTVawTl2cxrrhh25YsPWM2kY0hJ/bRA/ersYzGkRoglbKt7WiNvu
luxMYhSXl7Ask8FaHLchHjtoPFGWN1WoSrcVAA2R9nX4YhRVqQaA+QGKY4tkn1sP
2bGB4/+A/CqzFNVvBsSfb8DRyB1rNzvmloKQxHVxRKI7fAsoLyNQMChs2CAZZ2qa
r9dJrbbTAINxDWVVm3LutLGWl3dXdo/vE4tjf5pGjPW/MANrJSjlJy5Ip4VtxtQB
WzwDIVcYsIOJpa0kClNGGeEOueD1IjrrAp5h6Uso2Bu3itDnof/v6f1UxHEe7Vsi
+5DU/PI39DrilZx0sT6z2XH3CFK6rp45NjDAjDTDZFchJ7zLOvAqa9LIA0kXJpfl
fYakoFtjiHP6VHWNFWcOpo/mDXITmfFaSwgGlh3A7DY8Hz/GoQ7gWBIMk+Q8cSKK
BhuL6Gv/C/dbPGO34PFroDzw/40o1C/fXU6nloHCrlTgPdgHwZ0i0J+11Wlgq2fJ
Uf9edtQAVHLfgiUhQYuF9Z0oSkxPDOHSyaRxAcHG0krdA7JL5E0w0zjjAO3+MqpD
vrplci2i9PLZ5jzWQsI8Ngu8EU6WLohbbZLFsK6Wz0KWhxyC/tucnHihIXAWgNSA
Ncnvv/ZxuWiT3edC9ntYGLTy6t1PMg7WHI0Nawn7Pc3ex13KJoREo6fJGCUKt4rd
erBxtOBvHUrBlXFq3INWBhKUixr2fYZ3IBgadDk95ePd29K31bkTdMGDPx/15zhW
pKp2Ii9n+yoIts3VdaTMVuL+V7tYpINJgTiqOaeXIXp0/RmhIwDCb3636kDmJQFm
i3DV7/RZatw052tkHpFOfluCWzkTe1IcSgckGerROaFOzxlZMS2HnhhFqNbVvXlk
iECuIo7NCUXCLxyWHPc1aRGhKFR3QUFEbtuNFRNXD5QdFZoV9OBBzwPDPwmNvMhr
Vok7+uQ608J3MDoHZgCYIIRu5yRj43EBeoOApAqhEInOXqFLgiygr4jlc5+ZIdG1
zVcmEu/yEeQ7i4XYUXsx6yz7yDao5mR9nc24IlnVwCG3EvY8hHTw5PiGj7m8N412
SpuMbKDt3yyb/8hK0TRCn5tt9Fn7pBDeL8+Kuoz9yKmIwucH+Qfux9xRsHvaV3ZZ
SWUL6Zo58QMgI51w1FIAKoJ4AchEaO2B9/90tnpxCHm0fh/9uRx1IBRGYluIc5JF
trBapeFA7Qv3AR0jEManG+O93+jxTWAqwxK5uPeIKJsfa/GvtlaMvzVncaHYMVE5
KN5xeVAAHPbYEprS9fiHgBARIzpxLOP6nf6tv+Yd3cY/52TsjauHwHdJ8IStDGML
3pmN5ONT0En9tBGxUnDqS7Uio99mKhqyGV7bIzmQenFZh+2yf2TizV4U/mL42WiK
rOt9rAZ9N6U+sr1xBHd8PNllWqfC50xs1KnyjcM4yGWd6HGOUbXu8XKFyf4GzUu7
sCvgf+FQPwIscghD8h/yLYpcdQRpWS0RkMaLrvhYHsaIbXSoNr22oa0szx6icCVh
6bvXUVg9Qu8NudJF9jttcsbvdJMzQzOi6sYXvms0a4leQmEiqr4XA1/dWZ8f5boR
W+9nr16s50B62wknHxtzWYpmtvNN3+Wdoo3z/H2Be3ico8rXADfeU6LGBVjsZuyq
FvF9c4/lcZ5x9yYohVcygwrRpT3/yZYHQqsD+sb6Rl84OThScedEr3Emu3r/LJTP
sL4IiPSF/2tTOFiFzRwAnFSaKO8K2Z3YWlpCs7JGs8PlvGjn8AOIUvebOJLY08nP
sKcTkFkhqrNb4CoUsKkZnzhUa3zQbV7qTw4cuz2atzp+sk2E0ktoCZA5j+qUcKVB
mBXVqQFN618fHgn5jPbOg1Mo0DPPWdmQUdBPqLvX6ofVlE+XCYQ8nwJ2kwWspHzk
/Yp0V8aAP9+yRk0lW1xXO1Vk9yu0cLEt/hlRvJpOiDybWKfyNA++lcrFkoVXt0IH
+FC2bCxEsjxiKCMlf3TLM/XB9GrqZYGM5+SMjUGSILpIAtUvMH+9jXAfVMhaIPam
Xta5EG4XDcbzvG4fZPZ1YRXEju9E5T5KOHitNb0S2Is4/N62wXVeou1qDKcK+PW9
mn2m9LOp38Hd7W29+UcbnEAhea7PmH0Rh8I5khWsj2ZzqNw5ZKccI1I3pA6ZCYVx
kWYh4ynhvSpqSC12UfNCripIUkyiyICiThxi+mtW5K+01yHXFgGnL9P39cnLSCFN
iN/ctrzIgvDhRODu7pIDnXfYOw3m9JMIKTesFFI28QX6MlAwCiRwSz/qD5nAdps9
vJMl0REZm0p1Jikf163ErMI/ThA3EK9OADchFuA8AncQiawoCUB70ZOWEdef+Hgm
apukQV0VKKBdbr3SQ1ie9T4EdDwlYFsvAGo2VCaRmFLKuMG7hCia/NAyJKsNCydO
Jllj/PhRQb1HJLrK+L75OZER1P6GKmTTwZFVYX0pac+RTtFpAxFAbcS/9oEl41Sx
HyK9GzjPXMrDPn9oFZ0S4LEnkorkMe0/wRQ5ZsTRxApZWRRX5omsfukxgteu7/pU
rfrdLni+Ifjve8Jnmv+K6c0RxG3xGM23RrGmqmu5B7/ZSPnHtJ9Bs32ZQVtWq7Ge
OrEVwfgHOYNwH7fz8LGM2b6xN9iEJFrzYVaOkOkOk1rJ0WqCHy6zlmWb72kmQcya
Hc6cfM+dzEtazQNqNXNp/w7MdgQvH3leqo/dnZvLno6GcZJKWkArVx0GFsD6c9ip
01em4wTtdDaH0NRLjLpTyDC7G2m7//NUN6n4AwrKxDAgAL+EwhZYMBeoaFNDiA2m
LfVuodHfh4cHqGnhanBwJY6pmwNcorEESnmrZEYvQS3iraQKo8mOZT6kcRp2KkQH
fOf/6Ge4jR4D9Pmo5e0dxRdloiYGoSBf/I/Hp8n4PRLoOlZvUorMDL7L8X5d97+f
Vj7q3agI35nXySHtF3YFn2LvnWvaso4MwnOETax1dLSvCjnkRRtoOuhrlRs/ksbz
kGGxdBVlovtue4xCTJGy5sswxxXcpeDwBUyLV/HdlDI3Ls22uUzp98cNXxgmpkmT
0BAzRqsenEe2mMlouX7PrMjXBZmV50wYwD4czREatm/fZXDauA1ZfDvjBkQSGq6Z
nDiIKffcTttXinFfvudJaAgOniTuFnwsj+YFNuYznHtkBHB3gRyQoejApNbAwWmu
aK7FChSpAYcUNQxwDuUTuJEqwk4USXEYEziXNRwS1UBI3Og6F+sjPojXLXNBi0V0
5ctOHSId00Jmm+FGhrPqgnLi4pQ1U3cc1ru2C7+X5tWNb1uusA/lI98ydR+RIGWh
iBvY2krM+sKwgsJaqtVZ9Xn0eRoLoZ03PMmesfwPL8RcKML7TFi6qdFd+D6O1vEN
coWvhf8zaUtm0Dkk2XgXv89FlnIWSvQ+QmlCFCgb7Z6DwXfBiHb4p0KZUQIvaTn0
zWySpp1xBooWarIzHjZbwAyZJ+RJR7aR2/dmviZgFgrF39WebTxRtECgbaRYITti
0x75KMwn/4QBoR1RomNHpxV+Qtaz9UWqttigSmBG5aTndK3zH9A8Jvns+WlLhFeF
h7Uolc121UA613GyywaIbWunfGZiH6rTPH8zpdDsAftwZ/us7WkdCTOoW8qSVcK3
ORhWZDw1wx1DGmuTiboM1f+JnDTa2TaqF4r2mXzVE5rtsqjmrLSq/90h7tHjWh3k
IqMG100aoglWypkp8noK93b7BfrDEB0G7P82pdW2ltBfT454GNWoTmMuFwrVj5Wl
TLOr3EC/SUqbSz5VIrYO5YUtPV1vY+dDwaN9chjY2zm8MXR2zwesuOYDUetFnuwz
w0xEM3cAQph0aCn03fMwNYcY49zhg9m/FvYk3VL7kzNBvXrnXqGBdmjZ7tQB+ZTB
oWhDZZfELMYFof/nNyFhfdHeGu9+z+6og+s6ByH3yqrGiGVUdbyr8gAVGNtI+StH
lHqv7pHKRvrRb0ZsE2zGQK2gqpb9p4FUdWNOVZppSAD1D12W9E6Q2ymcMvX9lNCf
x9LjahYKuWJqK85YiPcnPt0buzgWpuUeyAizEBeyrIdsb5xqDNCy+2KueyPcKCIj
1OES+dw0wOGLsjFZf/DwG7LNBp/ZgZ8t11oJ8yT5vK/EtJ8nlfGtj8seulz2YdG6
xJaAv3mR8MXxRIF+Uo8R8znIUqfsIBl2tuS2mb8M5IU4QxtSPAY3SYfqBjI5DED7
wqcqgAeuwKndX6utXsX1HiDT7cMythdE+evo7f1mxhGcfMA9r7SEy4sIPn2wjTts
QsPPPIWqbSqWC6PPwafiKS7nRrosVvu1SYX9Gv2bkjmsDQbJhlSgea15jMV1Wyhq
NbDW8nJ1W75jdGQlEk+2EbmHqjQ+SajgfWtgrzTS+BsnWavqvjcDEtsApuZKqcGD
MJC2emx6omhIZanDUgM/HNYC0v+mCXSQ5Mll/f4Lq2eDy91oGAkEy6n9z2gqfQMQ
04N/kB8tKNQaZFFnz4IZCOTW3OISO5xVs8Afv0qSZabe5FcoWWeNv+ZL1sBALmb8
nwKfpdJrqp4Bfw3yLMktHBZknPeNc600XTZgp4vHBuqcyUA1DUjMwekAaDlWSqu0
Jx2pHDGluL+52NzDoV31KX+oV6eYClNezpio189uyGUbJe4F+ufBvxuMxbnZb6zj
1yWKBqtIx+bPz3b0Wa4qhWr9rVW0b519T5xvILrTTkvSkD63BcDKJCTmMlk8sXkB
3v49a3AMFgGgUeRbAUyqVsLleixi2N2ixRTBI7JhQkOYBjKL1kAo4N4RZfSzyTuw
ilQpJpqr+Xu90x8x7GWJM6xuAaCu5tHROT2WbPBZHxhyVQHb/DHj1+ucuKoBvn3v
3iY0T7cMiSMvLgTNAMJPb3GFHIKEw1h7KrFBoFTRM9QmfqPvzhvGv5Mx8mcqgqwB
aa4GDEdR8/STvA98mPIklXl+HejrcHvi22qfoiSplJ0aWSkj90tRnckLcLhqRRxF
QB737kEk5ado/eQa6Y28KGPNmfzmdcJAX2GxM7hEqxan3A3VFAmtRDjdA4Yl2QF8
AExjO27cAptu97q+xxIVRPPJiRnFOXrg8g3I8LVCkFYxo0ZHHR7UarTABIMvYO8i
jWMO4/N9O5NxNCHSywAC4lKj5diPk7C6CgiULyElaOLKkRi0D1ggfjiYym3wChWJ
Sp1JjOGXWTJO3OElM6FMLBHWZQNkwPmZms9s90RIHtZ3Eo82cg7ZrOfEZEP8SH3c
m7sdRy36TSZ4KDmijaLU9hqFxEGbM8IxnkB2CUB9LyKuUdjhf8Op0AiDjY8XqpC8
oLu2UlJNZLQJ5XaNYgIgNvKh2gqcwOk4ISZD1xCWx8FAOwdRySe2Fs1vgsFXYTU2
eairkNUsX0x3fdOngtIkro15mu3cv5dVzIjq/ocGwQXqnqLBu5S+D6tM7YSY2ZJW
RnzVzgbhv8+mQiUNK4fTKOUg67ATG8gdWr6JPhV9UMn7wVT804kUuUti4OuiHXAa
uH6wigB1GKVKlfsCRrMIbJWMqYxKtK9HygbOuY3I/yOLyYWFurPpu2PDkuOyaCk0
EKXTCmRxXx4kQRGjZ5whjEBKF732oosFRDPfbcgnutsWJLsEze866lckZ8X8VK31
qOZMYv6qV72tB46Bmj1vICk0Q2uhqJpd0fRuK8BKAaMqevQdSDXB3JulkesnNUTb
cC/2rHVGMsl2nV3uvHWeq+uGBk9h8xzDYLTCWujHIq6BDHDhan6ctCmOvK61BvwY
qJUSEyhpkuKLPPf8/nlMyrDR4tJ7NF2RZ0D5X2YrGpSO+ahxplaMojxybM4JFCFu
gzFXAQ3E1NuvolKoY2vVc55CdCpdqULfHTjh2Bk2nSbsd8RSsRo1kKF0AytaNqAM
YI6dUtTJ7BINMICF9v/Axu+XoxsFIZnJurTC+XpDQsreRSxnn3iKlRldyiFe3m+6
Mk1SZIlMBcrX1R6QE0/BuEok5BIdxaSOBXiOjBviHlE3sq0N77lnbcphPP+mLrSP
jjY+1RxY4wX4AkIrilsLDbYtrvE88k31pONjMbb+EDhmHnur3Pi6abVsMagmBREQ
xixEr9FISVCAKRfpcFmOg1eDquSkUz/g7rnC5yzvYQvjeIdmpH/OSLN1EoCDjD/b
B7RXFKE9SU1YZzJ55I9+XPH6yhbLXAU4PkEkfGGtmpQYHc7JcEBrziEz9dkD7Crp
gZluJN45wxSML0KnR14l5+kCvwTKu9hPnWJINzBdj0D2h9d7PlqEbZpwCfk9RRUC
LID1gzVUbMXA237KfpPY39ZUvp1WxiTWPLvWHqvvAgT5JXS6GjvNfDBAfQHx2GIP
CtthY9g2UlZpCtfV9B76OqOxDcwx4zxaKhvhVFykaThfpC+WC1FJecF+tGEs7Axj
XMGmgvfAz0Me01/1kQO3V91ieooShueNl0QX8aR0sRo7DEKT4PUoQWJMPr0EIx99
dXM7Fgs3tHd05J/wpERjt4MrtIsY3md/dgacez+/XpUlvwh0qK8mX+9/opCwRpON
Ya6Wf1QW5uvEJ0a4aNGt7lu5CXCnopyRxAWttax5RZVdYtfaa8GM8Wx+b/u+XxHT
amyYg/6jgC2I9cMJ1s7sOvQEUXkUWmRZxsVGPgFcXpTySLefaHIJpkm/hy+9YCy1
4RwbIYniTJoOqzBZhJ5r9+XGl88D3YecL2SWT3Q069qCuanm8KGXf4+kR7KuD02P
Dom013k/qcOBrs+JN9nXYtX0I0ifQfnLPT/W10oHx6Y0qJ7odAQqxqOG+x4Cd6O+
2cCVlNc6GTQ8x0VTGGPn5HAfO//rHDpgUnilV+y9bVntqywww54eysCDJrRUpgZD
C96QOziaZYRhvZ+JX66MBnzrh8UugLkThaG8dbo+M7eLDv9GuRiKm090RdD95+1w
VcfniE6aJdtF/O3AP0NpqHmCsFApUfNLd6n5bNdmt56wIR7fy5y/ovtf9wNU1J//
RvSPp+yqHG+vTl/zXuvg7zGoWuX0nFnvkdZIPWm5p673hSo9nJDkbndpAQbFGNkm
YHiNf/ALnE7e+Rr1Y/AlHr9jXTkIi4hB0YKS+n3ugXWpdzijdsb0cG+lxApLvxlt
yZfBiVxirOzwdPANYsiVGMJ2pNitEPSRwzi/w/Dt/b9Eabg3t4k9tgUcdIMyFV1G
dCv/QysvOnTwH7XWUA42Jq3edLBlxERlcGlGCQeH4Gu7SKx0XBrPTYmExIjRDqB+
gFOEoon/fDfx+fgJa7PTKFR31ld7JwtIXusgsgnUDLhX5hbMq546RiZCVLdGcbII
FysIxapNhONCFoLWLtu99tGXa6DbmzVlOxAFbkYft+dtfarcqdgdoclIVrXJV5gU
ezkfbpKgLXFxm8e4SCvV+gkWJI8VUk5NiXYrzTYt8iBUFsgJv5DLKhZ8GjLetlKC
SlvPCzHNCk7QyP15xchZ+b4lpKcDcsfcOU1NZP4jsxY81Vgx7OAp+RZvxdxIrgn+
rDuMFQi5dgb9Q9XOH6hfVpMJ0oOA8NXh1/wHT7/2QhC3vMuegCFfkBXT/JWSY+5G
wjOFJTMK1VF1nsO/pN8qqJ9/nlFSgbdANB9y6Q+KiBL7hyFDU6EDJXqWaqMqqajK
lZ/lKucix567gQfnYN92L6gmWh1lmTIENJzZYjSJAPD56JXax+FHxAIworRI54i4
0zVtGmRQJuh5naRToS80ibWdwuJXbu3/+ISvNcYQtA6J9nfUlCSSqv/tLAMaQZtT
IKvN9LMAJv6jwUnj/MXJqR2ho5ntjmwdd28c8BQVIQXE3dUPUBn69BsYBj47i0mh
3wrFfHmstYyl40RjVLRerqvn/UIjhMcspm5KXlIDPZQAmxmB+/uPBXgkQSIikCoe
rNjsF8EcKUcbwLxBN4lZDdteijSdA46nTYXZnWqhApGGKAWg80uEaRlEvee12Nnj
WuQqzfjv48rH7Daypc5PUMulqteyeHPrtD1pID1Hl7DOuN23Ie+dEK6+Hn87gBwB
6LRDaU9LFti4LNclchq7+gFXHSWGzqNEJCfGhhk0Jv6pPko8/V6KeQ3zaq8Kfl7T
8zAw91chVdvdJzuA9LlY7o7BCygzejE+Hcka2DM+ZhmsnQlSQXz2DoFlLgXuuyCW
6G91XY9tXJOOkHpwKt9xjkFL2plWF/bQdrN22JJYWUrqV0kz5yAlIYO4uEp+vAo/
hzWW7i1FiJCvRFopE9DFZguj8mqjEyHw4A6sgYRIeyjIB1FpKmqPRjyWWDPpsVyj
qWTuScJOKFEOObz40aq90gkG8w2gs2AYTCOFfECzB4QZnuVjyKzICGu285u4DKvU
jDOr+MKvBNeOrZtIdvqlRFocbKaUasE2dyHGODUhqz2a1EW3injAqOh2pPdF4+iJ
74Cv7iORxXvm28IjaKnL6KkFl+UzNydQ5A5nX2s/u5ymdsvafy9+z1oCWUYS8Oli
1PKMvMLCVIN4b3V64KYPlnGeqC/grftJR6Ozo1P1kK/BXTWQQ2siZRvvpDfk0D+r
ar+fRQ7VTmO1YWphXl21qqyeSrNlvlsX1sb5DB+r4NJPTz6brO+rtO5CghZwse+e
efbb2+jbSpa/YBhbUAlyTAY3PhF3vRbsr21fwWYJNpi9TT6U+fSscogLhIgdmWCl
eADaZ/jrIUV5+wLAPnuQsqAFHwA+tzb848VBQ4BVEFZw36cvTWRb3rlrHReoct/Y
+izo7FXllp8dv8tJxKq5RqKwvJAFLyzeZDTkpzdpCiUsANvBaepq+ViHjrq42QGw
+u54VU+srHsBrcx9Yp9lYzmb+F1x0CnZv1iNfKckq4sCeVMM6B9Sse9GLDscWMOF
sn2zS//rQ9I0IE93xfLISprGYvPPYvV0/eH+Ay8Mhrc8kDPutjJoFUbLiy9uqErV
rYnTiP79w01etGseDa9axq6k3O1dsZf1IEN7nxDirpO0zQwowXX342RmxgMkCykt
s9o4j+ydi0t+LfcCXHzoYajCJ0GFOGTeEZKG1gMe+HXzzq/DEWCnQDx41uc0PB33
nOy5EIQNlVxCtD2vTz4VDA0OzNHcyIH6tLan9Bc7+ERh5rc9nkjxgN9FxuD7uZ4P
M+GXJXpwllDhwGagbsU7++hxHnAw80SvoYJG7gJ/W5FFeqAke9AuaeFr3Hv2AYZE
uODVjHF9LlmU5YmYQKEK93tkDVydneQhC1vO5g8UB2hSrBqssn1UapFhZdAFBHKT
SFzOs3Y4IEyRqvcMaBNNVSQBEycBaC9d+CZ2TNUwPlE80M6fyoY7MVDndHHt84Dc
sK0WfW+0C10I1ug4uWscNx/vzpExTzg8X97bqbt4bJQMuHNxrGcjpq+0SxHh/tJ9
J15fDnmSLfMHbcQf+cOy4Zb0pWk+z7ACJse0ObrLnu0mBccjTFUmtQoCIND0tWin
o8sZk1KyFEDFmtBu4c9qCrJbUwuBYA9uM4AJpO2V/3hlbd4eo6LfftmAk2Dh2GrO
6AtKG5mTgBb9BUnq6KiuUSydKlsg1wowPRJPD3Ys11STLBcJBGht7/B6EidoXbpK
KFkOip/rIM17Bk4DaXBpltJ0NRpIzPAhR//hwS9RUvWaVNRv7QPPhnx9eRuKByHw
EHgIi6CIfJo+pOm4S9c6YZQSjjPfVi4I6vOu4UmrCzYteh4B1VGs1Prrc23esht3
wD/l9+1CfLUDdWpwgZYQ0ZXL+7fevcaVdJYi8hxRxNBs58S44S75OJffiSeh8c0F
2RFl6vE4nDZ7kdg1c/AyeF0I+83gI7kFSsp+OguJi8RYMD+1a8QIE8RSnEXrSMuL
T2cTwil5ZUInCLd9frdcb0ucFkIkpOoIlcIceJZOtZAelJBAy20okZxMGD2Qia1n
Fcc6Zh2bAqaXBOKkSP3iXEexUz9RlS3ICUbfJF54Q9wWqJuJBrZx1NXPWqGI3Yi+
/Hy/Vbqu99cqD/vH8+pDz2bYiKA2EQlNBXdZSAwCOILj73ZZPyAUn3uy3G0lganZ
YwEiPESp9s1gGsc5ugjH+MOI2cmUguc5pZNKAivp0Gf5LqPSqwi7UjpzJpYcnJNG
OM9GyUr6Gck+76EPUTcyZyj7gADjTu6qQZ9+3iDvbOrcPnwMn8CxO4qXYXm816CU
L/fQ0FANOtfJmL5NkO/8Y1Z6pAdDFwUFBCwSF3Mr4ZIzqvVi2/5rxSMRHnPPZ3ZQ
BHgAA4pwhIOnAR48SSO6Uk7w+VZL4gRXhDN5HTp8oCaYbp6Z1WSsf1Q/tkDcTEOI
t7G1rh3MA2+XfJBVC4L6ktR5nbM2j3HL+Q1HEGFt36tGx2LWoP3DYfX5QvRgdOPy
K2igYXGw2E/z8sslNqUEKgWQZQ5je/AES+LvzDFuTVa/NXEdsrrnMXv5rVoxo6Xz
uUQbESVa8uaGLi2kUtrx08zuUjZa/4gPeA5ldjj/Jofs16UkWEpXKWuw9d9OoO04
DGcdKHc56nyi9BKsbI3KNARA3ZP5KOaKS+Tq4O0GSaklV4VAnpUWsZpEMmguvjXB
pjv162hNcMP00aXTchYhOx4qPv+oOCZSEgy/LELnb9Yg6pGeA74v3tU4zO1rQEYJ
eYo5bagRYe+ggtALvpMjxowFSRgA7XedAkonxxj7cnrmuKl+Dj7uOQpNzD6sh6Cq
SboPLx8517DHC4PrjXoV3PVEFXPl4wNUG080KKcdcK3rvpEw4TGXJj7qU5Qe9498
yRKF2VvwE3N5wqASGmNw1rOPvWM/nBD9aEaL6ff2gEs5px0YeX11fW3nVP4UclkA
JGMJ6SgYzCDngLd7pcQDT9NrXhyCITyzVZgCqmiVvnagz36ylMnj+sBT2u7YSHR/
8rbCqOBetUqLNvzLLxI2NUgU3RXsfSUaop1gWMv0rYlJctV/HPUNtROo/lMTKnXJ
5wDR51Or1KTwZ8XFbe96g0vl6VLPt+thuMG3WGUASa7ajXTY1fb88VJYpFdDMAl/
BIK1OczLmi2gkjeHmFZYrbZULhUqLl1SMC1Rz0BaDadMG1wL72H7FPeprnGFtjbK
YfDGCYZkKtbLwtY1xTEkVAdqbavs2F5rSZS0m0PdlA/zGI1uZUrtPcDV4g23fifi
FDhWABvs7TwmfWNsJvmtwUVh5QmFtiL6snWo3uZ8ChhUpARpFNTspPs6ZFnTYxcd
VUGGOknQssniFenCXuD27wjrQoKURbqOel6AOHwT1RxnxsIZ1z1WK37CR30uoM63
glPlhTbCRcNN+J1JsXhytGe18eQy2aJi0FgZE04EycLVKVx06sd/sUvS83wN8iJo
URIrDAeAbyhtxb/0irS1/LYe91eAn8BceqQxfDD55o6/oI6xs4h4TTNKGY18YOq9
j9Lss6QdFTIUyZrwauNmWVTK/2ua3pDkfKZRDtxbtcPC3Xn1y9t/lN1czEhqizRi
FkwZoCbfU5dqs89nyVpqh4pmh7q0R9Ka9P0YPRrQaEYoWhEPqZBnznA461M/09f0
Cbe/71kM88+ul6DkIxH5l0o/DnZg2Q8do6cRctI7n88zhdrzBbC0LVTx7EYk8iwD
MuYtQwzbNpuwg1rd7SUZSt2hPCxLyXSdYsB3+QR58ZFC5OpuqeIObM8nr5fXytq5
Kq5guqSDktImfbCd+NQxs8CGaGYPIYeyhEpsQmQMU4rFfA017SKW9XA4UifkX8+u
DZ/3mKKRZBX16Y7gNdlMVP4X6Tom1hpQfhr81Gszs2FRF9iNiKl2hg1Hi/raI8CR
iVsyFIYeldidrzw3cLUvGDUXzjJsl0G70bjD2cvQP1rar9tgs7H9Q4Zch3HXKz+3
+t6An0yWFUNAN0yOwClhkozH/67HAmuW7vTlpdE1VpNnFNk59+tgU/t+2rYPNmf2
RwHeYou5BRhfhq/40JbNo93hqGvB340QzYw0RPiQgOtWhagWggiOMW3HUKShYT2O
TsSgyFjZI6FeeMwXeDcNmxfh14084ZbxZLPQkq9C+8wzpEwwoPmY2yAFEtctx1fm
R6TdFhGCQTndLMANJ/3CWBjd+icGbSdXwFWywuvtEoh9YhL+B7fPuH4uW8lm3BI4
5fxTKce5xfsXyenfv1WOdAYo8uq092PXlmeiOl+Hr13eCzpsBvTJGQSpBdMWVnJB
/PpcIYZrv/UTrsTGoYISbBpKj6+ivLhXOUykW/xn0Vaw5RNfjvwkMfKc6S+5pzVF
juMuqRR3bXBl2fKO4mPVu+hnxWJK+XOthYFJdhO8y7nwpp1HIAQGP2ixuDqtEX6G
if8gwis5SXDhh1ezw6oq6OUdGyV0pPgIYv2I0bXSP5umlF4/SxS7xonTou34FR1K
viSgvNt77s6OLL9DuO9z++DpwpEy8Wd1jk3gVj8ZkHTwPuUIp4PWgLO+XT3cK2y6
lXgi3GSyzEV7rq4jtJjOUoN0gOsptwstuCBU5k1N8akGsMwxU6J/wIHxSwS3Md9y
dvgjdLJ9rQKGEL5CHw0jbSQENBzQnXD+wsck9lJaDNoiNVkWKnDAJkMMSXoJZJH4
BBlME/Xymx3JTYWlGv4b9M/uatbkXc+Rc9uZpOTppDwpNCovEBzLFCDb/BxNLL0C
1OcPZbluOPCISp9eSfpaH3vAL++3o+QGbq3VZlEBRDCXLT5uxpiI1DglrNUWUOaz
ffrww+7CBdSYFer6XvhTUdh3TveuKOZ2JZB8fHPBnRdh/+j++OkqW9hnr6voOCOG
QLovTC503D4QwgKf+YW0qF1JVsIo93ZFXcvJrukFOvbvPWH5kPD3kOEZAKDmhdX6
idg744BIlsUtl5WCY5UHIuOGUhhERzXJbOB3qDYFxkmw0ttYWVOQb13WeZkrpYSa
M5cCiPu5PCvAtcAil+qOkhXggNTbgZwGkjqWMT5zch2DNixneALx6qWNE5r/q96R
lURPo3/mHpIFwpjN38FYXeC89w7zJ300Vuwj/NkWF+WKP2gBfDAe2Ps41k6LT9om
3HLAAE8UbzQ8Ve7bSUui6hCxc9L7Y4tDlz8dxzQCyCmH2EdQbxsbvWK4+yDykf50
iqokS7XMfYnSMjpjvmwLLY4mm0bvJlXZfxEuuXJoXAf8FJBajAO/GQWXkNjjP1Od
IuR9VCm+gBKINlyDtogi1zIXc4Q2JCcnJA1bJhQcco917CZyzYgz0MdOsEVmQp9o
7uLs+uzSYJfb2TvnigzhY9PwMVZgt1pCaJR397PsLBQ0FqdnRqZWOXB07N3Wf0SO
EOj++WZOKbwlBWJnPkSKBcKZ37Ls5pG8+JTrcMCl6648UwsGWE6Ng9487XN51vWU
VxEwE1n0UZ29kk0CPuVadGYPwyHhLEpHKAOGDTqEkUjuAXX364AW5Zeyo3OUwfPd
tYI6ql+CPJ8Sj6Z/NKN9FJm1I8q70AKkNfNiqxALLLPd/3v36M7k837lZZpEC9C4
AFJEwNmfXokpFPNjxJcQQ6YKRs1mp/PMRBNVcl7a9vlAsgttMpBH8zXDckVWgqrR
ueR5cMGWf8wK0ec/yIYsyqBMh3RKPQ+klApjo9MLF6C/q3AgYMLH/gFMDpU+aS4F
blNsE3aN1anE8LEYxDrUedUgfO+usTC1D+yOg/UJFQh4dUOH2iwzlu0oSufaMsPa
Z9YggxM5TEIG/fCe4hQrOctM1qWzsiKnBsvI7d5C9WwvmtoXuXsUetGgvZcL2scs
9CrRIZXnv3JbayuoMx1kCy+/XtomNG5y655AS/M7D1of83MAIUT8FYN+xWKagAYr
eLWjee4f1nW8V308K31QB8XLN62l9FXBMKkMGCVZ1oPSDwLsIi1Qo0sEZJdZYxII
JntTP/MUYUpxokrDH/PUZWFxn0NyiW0jeEQrYxgS5Lq+EtK8Byci3eV0L1si1Sel
afL9/iNxnO0ZxAiGBrmmWXlOqDRrbF/o5UGDEODQqbYcYoM6UrHqhKSlArBv98+K
L/wdaWTXDlOlH8XY1bi4hIHbvOR0duOpyM2smDUSPoXM7NxZazH9fpHd1qp/bFdU
FuQgX4kL5wTg1/vZfnOcZUfxriwO2VyRd5QhJRiuF+aFI2ufGdnLOiqA7gypqlVC
QAQ9nwtfiESjDIJWAYfdiqhuInIRoiQd5MOtugX5dGGQpDcI4dxFKqeKbGH+E0K4
29WHnzgAwih08Ks+NtB0ZqpMbIYCdIor0V2rrf5lAmBBWanVEg9k7MKsZwNFtNT1
DyEZnbk2ytWeMkLb9wdyKBCg2f0D9c/whBCZE08CchhInSkpbA44hxdgktbVYl1L
t7XzXoPfhPbG0Bn+/qVW4dQzA6irIRozxaIislo+jySmspbjvKxREJgS6h9vjo4A
a4XkN3MZWibhT8Qmoe4I8AbNOGYx+qqFw5u/2njL/cED9RGzwPRpwp8KFVzxr0eC
M3UrKbIPZTyALR3gQk+Nvk1NDs328M7wP/hSauEmsHt+1LMLGtxk224zpThQ3fz0
4pSpEIpBg63UGW2XIZra4L6YoUb/tC3kvVrANYfDaPuNoC/FPHoWdMAsOWWD0Hsp
+m2k2l96WZL4bNvpmVXLGeaxlr9Q3fey8hmbE+KAQFXR+9J6f+NE6mOiF1QaRKX5
uihA+L32cAF0cnD02YYitHxWG8g+aFUthOnfn4hoUfdvVRBtx8HzEB2I+8p1p1pp
ezIVfENSmi1Zw0oBDZfDqdZbVwf/CUOr8nxnOa5onBM3ySunoh6bPZpHNv3TtlGP
Zt85cw1C+50ojtKmA4ydUgXPPhhribmFhcZP2mNvVku+pHSk+rtXV07CR/Xh9YPe
KL+eOZgEKugOE/3d0YF9Mbmzgt12Y17bOoccxsOfGLFPsiL4+Box6bQcd2psKE0p
Jpmfa38VbiuE5w0jzF96Iaf1aosLY3jy/1bL3fgrgYBog3Yh9KU5IW5JiMtNLeK5
YznIfaT1O1pH+LGQZ82bKmn1WxPPQOf8ttnyVWjmIP/ZoZ6U7cZFNdZf7WL6v+UP
aigryQJLHG8etC2QAZPFWX3o+4I1MoSx+c9NpnPNUprmk78pu+Evk+D49/vT/rJe
8K739nnkELw69fZXA+guu1komjn40r3sHAOORL8aIH7pnAZJcGXEYSCqto0dGFZF
k97gaXHCUWNEcJ8GHidKYGfhhJ45oLcds17164iRDq0KHHhZvJdcPI/VUbwx9Nbq
MAxxXIHKNZrdaVRc63gfd0ag4dgBMzX1kPbe67Ep4tC0y06SrATx2WrlAjLmgKq+
mRs5Gz8PlDqYWBq3pIGX5tJlFJ6EZ5yxBoZ7E7MklI5K474l/BIEE8ZPc5fHYaiP
ZHTx18K41BWNB3zKZ+UJtSsKA+cSlefZdwbFDULu9spE1G8AOEixrw0+pEK8Nf77
byTL7DAiCMQvjmZDVLWH/RZpoMTO1T6pCdg+4g90yWSRCe8eof3xyv/k2DJyfriX
oWhtIQ5RC4AZIuCQT6fYEV0bIH7OWxKBWKBR/hKIywEQD+425HNPfRtfRPfzfrwL
oZiKjsdF3AgiS95my79Dt31rrB1XK+6JU/WAMoW1fvtxzxzcO5nMgPHuXKmfs01/
sc4RtrPIH7d8F+tolPZewR6nQHvAQ/Z+AgF1f5lgOn3xIRwMRtO+Dtde8vF6WrPl
h3iP839cc7KirWdJN2WMMaSolG0B4i+GlTWXjbghQYxh/U3LRO3cTOmxqPL2kKBq
SzvLWzYOOS29tkeDMoiFXCec/2fgfkruHBL9r7a2BdH7XSa0NAP/oqwAtmXS0g/W
v55jLBrFyHn2uEQ51X6B+HLcBBe0y/mLki1UY3ShSqCjCKyGASZK8kTbFHRbGH7X
LYulaQzYUrd1OdPBYjNa2WPInPZpIzaz+t2yFUDhdEdXGmkPk0CPb4UbbxgOEcPB
1/YRuA0f/2pBcnWPzVE5ja+5jJ6Q/yocN4s9bWwL/YCpvPBansb+ELyINb1aGi6p
9JtTIjwQOM3B/f1LAIW5DRkU79HH8kBG2ZjcySW37rLLxpYmnzN/HNePwepH/X0/
VzuCen51V0OC+sFeTC9jHUkZ6wDLPrll6yYXh01TQpzc4C6A1Y+pVKHqWx8vpAiN
ZtRcgtBdi/QNnxv12x2pYKFUyKuLS88k72gcw7Pi0qHIbQMNaFy8u9Q7/HM6ZZrh
Cf4dtzJV7Amk2k3REHh05u0mM1g5bx5qFd1xy2x+/E0x1R9gBAoYiHp6xmuRYUOQ
PFRHEQTy+hWF2FV6+i2CgJo3ZlfvI4cToh3H94hOAo3pdFcj4v4BmLsbNB4T251U
EBW5rYG3JFcONo3zM56QVbRIyyFL2DeNeZ/A2hKgvjZUy1YE0zkWiby0gyeSbuou
0xPDZERCfQd0YcIddkOuHD88/9gyEtGcQJjDDrhgTKbynMO47zgtDjduP68oknr1
ej7ou9pgM+F5iABLU30Xi6GPIrvD6MiiFfsov4v9WT2L7GcInr1QI5g22FCrzYdJ
9Et7OGQiuTmDZOTeSD36Z9iIWNn96Kxr7cTQ097ye09tgZlje8G5lP9hkanaRJK4
LwcO125a0ockYeo08uKteTg3mtl2tQfYA7FaQ63u1hI08pe4VEQWd5IxXPNHM9y2
gxzLpj7h26ps4wlLK+Y5T6wj5GfTHbaRIsPmkGmm+jk0+JHj8Bi0zKcEEyVEuAUo
0qs6wRwD2KEH4PfbGIUAdnkKGo43DhtFNOXZAtrAxGNeK7DrxRtX8i26eT4ZZjIb
5B1zwdHxNa+Seorer86QWbjGr5G4Gt/O7kuPG07Av5q3FJKv3DNB8MRjxY7TtdmF
nUMqqkksixBjkq+sSZQ54b6YHSA98tkHhLtlY5lZLpKKEsZlCFtv4XoKbJG1lwng
rBzap1o1cfuik+Ao9vPw/M8ys/o/5H5HZJB9iC1tffWfw86Iyk4BVJUofZayN5z9
UOXqyHgYJU6Srs3+d259Ke/25UvJMVOjZCMYWIfH1IRtdY0oLd48uOysBJt/4ZSY
9usFRg2AwPHs7+6XE2v1vIsVaCdPgxrJKOWOfV8hmO4GbJCNR3qHGCrrTdYjeXKS
esnbKjH+wSQ7Zw+iM1w69wRHpmRZM3fx5aYXZmu5IvMJk+QaUW5CnXOnY+vbcahT
jK0VV4QXJZwuAV4dNvuF9B6IYG8HyIY//OIYUnFfSizcm6chbF7vl9+aXe+YgO+H
TKS42so2dw5E5MOHjHKT5+jtbkqrdKikPm+nKVbmxhoR6u1VPYsgaXJJPHir0nsO
3CTdkxKAS5BieyV29XYO0/su1R/TUEjgcqs3ApN4rLRF4yJn4BJan6mOTjxI70ll
yxLaznfbY6XSHmzX7sQy9aeHXKAD4NFy0j1o5jk+AGNCXryjjrgIcfFwkQ8Cflpe
PRKojTa+akbtY3AgN2w1gKJPIGckVmZf5mqk937YRu1rsiwOtr2hLcmIZULV/vKu
97M6ravyusGBnhmXkujZYCToQ38W0dYRlON7suDO4ZnCUaQfx9Fj31NaPTyDdd5L
GBxFx/+K7vlvrwPhuS14O5ZaHt6rEnSBv+yIjE6wp+iAqfb7cNRZJ/EphVnFgxO6
wp0H0ZAB95iKtPQioyu9TXFYoZC+WWy+1bOeo8OkhXB26cUkT6/IMsLQVMPRj+kW
McMFNMkjsCiMuiDVC7MAePNBfrNCYB+YcYPXKeMOZqLCX6qL+MAdztMuFBohsFp3
fGsb99lACVpsey6+xYXqii2jny20QN7SRxIQ3fPoXYMWRjiOyrJJe2XLlJqerV5u
OuPr2o0gtGTBsF20cBu9NjCtOQk5MZBwi5ZAx5mvF2M9b1Au/O7voXOjlD7aTiHR
VXC/nAY3Zt8sskyEOtoi9ft7LWNEf+XN9xMdunQGFhZ5sRetOVcZeD/sUAd2kxRu
HSZ8JocbskQ20KPkGYsykRr/a9dDDnrkh48OtoF4nrcKJsoF64+CtaWaem67IVD7
kWCcSNow7PtgjYs4C8AVBvNjRHnBU1re7TapRo4clGx32cQlao/ZuomuYCIH5ijj
M4eOkZYhM33CM6OhPl8jsLqXkOMQoNXWh3oRahSBU7tnh9NPtYVa+R2pX0VSTmNc
qB2S8rzrX8WZtKTSqcNI82LnvaLlybJKKit3snDJJpxpQc/pEtgd74+UjRt1TQWz
4H2BntwSLF/9cy2eXfhS8Kyajy09kAUK5jpr7b5hdm6Y4GLKp/WXkOdu33AD2qIS
+6m5BfXpk+E2HhjJhLLMNjORkkrPfSKNZFYhd1k5J7xnWYf0+xwxFSOd/1Lx9n0z
B6bHuRpmabQeH1QnY7PDfS4kVLJL+GeIdFwZPRA3O5OiyH6SVWS+7SSCV/vOjTtc
vyFIw/aeIJYGnBLLtKy9LMDIC2df98B3AyZr51SwLP04FQnjUwdAPTaVKyxU8bL4
R7X+ou9pIy/89UMPpGBui8lTic3t+P19OGRFKEUcqQoJfO1/knvn1X7Lg4yw9J7P
xSPZoU2KA8y53MqgY5jpmq+cq3slITJmKemQhxYhfux7EERaeIRYMKUesHSxZ1J6
ZPv9bzXw9gxJl9LSFjolfBV7nUMnyVEgX7TOA9o4iDQ8NTg6EX8pL8SdeyH5vSP0
BrfJkkoMsJNPXArINqNNV42JUGUTIZ5HaHuD9nqCl+g5QvsXRdTt5lL/Ra/p6TX+
0hXfOmH1T8tOFWkFrbfiChHYDvwpsLTRkdHdo9hmwBOlvb9tbJcaIGACPL0lVXDa
Sq+unu8D5kmPrnrLIOBLcWidOSd4/rP+c9gUw7vQIfIhSBo3SaBweM13+37Ga6Bx
Dn1jzKvwrzr/X1wprVwlZYfrjyjIuNTLDNDRpYsLNyMg67hnmt0WodPf+ufQMBtJ
w60Vhx4pDaxQzacU+ST4t5e6h8ciLdJ4S9fgj1pgdilWBsjgRejH2jGzDawQ5Q+Q
wN7EPRQxbVpDReArrS0qNJ9Kf7SlkiwEP77uxZJ++1Pnfj9EBfW6ZWQzgkCF9qE3
/5dd3FE7D4sQzfvrdygKAxXO3GYuDYXHD43FFZvJd/4d2reU6r4guY/zvvrRHLyw
HO363yRcIK/HfGHZEHKsKKvZ9S9YcAEQreiUt6T66Z7IHnLya1SUfjSewn2F5GmF
Yl2P7nkhs65iM0hHthCc6wUYE/Y0FaBOn1EZ4TwYKorD5uqWdIHkRov8w3n8GBTz
MzWoeFsj+g5w/uspRXtuIEfZavn3ukHapeL7FEgQrBzKf8vWXlhEQUhZOFX4TDjR
NBNvYYVE91mjwbLHK2sJCAQMH/T59cGd2UvkEu9wLAfW5Wvl5/sHLqQR1zq0dL6e
VkdPwoSkpxQ0Lgszq39kI4g974g4lxwu4v4f7I9C3e0V9gXlvgvhN6YYS5qwd9YN
NS99TmXtfi2xKJwhAkl2v/glvwD7sBL/9oL7nhKJVzx9OYJbu00kFg+CHTM41C76
UbZ6NDo82VspJNFvWYbwRFjMqw/sJ+3QYsUhFDa9H5JWTDQBurUJ88xXBrJq41Ty
tm54oHnrPPOUwW37F5TpO0HXZI71vJHRDLd1UebHXwbUFITI2MRrBP/Tnpe0DD1J
rFTeoPunTY8qHkpTkuiQ5eGagtfXpvWFnfdHOdaMBPYZiYkUDmOIfjkgsViGWhFC
DPf40szOfiEtYka17IMs2Li3xewN3vcULQ3ZfswzAPMX6zXLKEeanENzVWEgJ2cX
F9hXlA32yxdmFi4kHLrEQNzXdNeTqNHXJ1msJAt64ULPUznBkB4q818dZEeY34yg
q/y4nIfi4C/si8vzjxOdB0aDJdDfsBd1+kaaFDqtiMBwQlipLVPC73ALmA9sJ8/0
SZqG9CnL91ClDVSM/SWm1vaYkOYHhJchWfR4Q9wpVH1xTYbOlCtEJlcos6zmz3Ek
LCf2w1ERvP3/zTkAgHejftBz90sDj/qmUZ8IAtStmKaggI0ELRlM4xi1Pm1ilfXr
LY48cunbB3SQPMm9rEqnHch0bW2vL84yh1JfwavQzy0H/x+A+5Ht1owvBVZ+exRq
GGAqvsWfAcQJb2du82N6XCgJMGi+DE9vPdm5mMbs6Obwwwof9x+feFUPONPGp6Vy
0cYdtb22GwpyzadtKRYaRWuynMbfwVvkudHUXg6EZcu10zaoOTIqOcKTChTYdx7Q
jm5j/BRs+ZjjDSKRrOsNDMUq8qInpW5Wo9MflwXw4oHF+4nCOSW4bskbse3EBJev
eBX4s+29+owTTqOTO2hc3YXJnLI0J3xSCmtA+6zNk40aZcccKrnOwAsAxkgF3wm9
5PoDgJblAxkJbQymfpHsGhh3s9voldTZvG1ToCe2pzwPaEsIRyqDDVrmQuOMEGwN
sQ2PahauPVtU0YrYLaX+yha6t3ECraf4d0oaYJ48G7MQ4KNw/SqssExrnouOVxo5
Qjw2xWHJEQJBXpBnIbNavf34B92yioLtdBIxWSca8qXddEjbz6uDbz186tLfMPIr
5c5ia62VfnLMpxGXN5i5cL9ln5sw3eLTxaNpw+nkXvyiQdJjhroYZ0kTdz8eCgwB
sqlGCDjnvyZFDhiLQ7lCnYyXKcBD0+Lu24q/Y+CWe6bR29M0sVQ37VYMeVyX+brP
OqqD8KeMPUDnMj67/mKnEVP7TPcOlTPmg5Ik4zkByj8fAL2Tu8XFZpn/fZcCYNlX
CzpHj+zZxdfJWDgqGR7y2MwHzVIIZ9lVUdBpYukePH3mDhGjpjXEES5e8+rQXQMh
LWZWtReFynWk0AtC5GuC3D1eYKSCZ23pzdKELLCuZeI+zXuLcOzU3szdh+O1YEx2
CcL50Ibe+6GOraom4tK87Jf8IJfVGEDvAMTJzD/XIKkE3Tz36yAz7LWuFNL6XTUb
xG40634kkk2aRAbFka16ukWkmkmB+bIR/485WDPglBiyEe2QRcGT3190FSGOwHEo
yt3bNnQdgXU6/OtSHfiiAPWTZT/Qw79q1pDr8bO/4FJGRiN9EkHd590izHTntTK6
A2DC7mKHERD78izaBmYayenaRXhpqqMNS0pZLm6AaYwWcl+211azMA3H7taEKjq7
25NLboZddErtZ4yfw0WUCjiP/VImA0sHk93Ij5mx2/zghIi6xHPKJvyGuRvTE4zJ
oEc+0qAFW8C4QMBqf7xstUrrczgmK6+bbzbNjxOXePK0PGQBLyZkou8lwaywZaWT
m0ZX5RN9owNxEQq+3fLqSb4c7S4kS6+fvG4/yPB1YkAUkctVhaY+O4KqjtmnjFNc
80c6UwzCzbEuMiCJHWancBzjz2sfDAEjq3M3NJX8HVOUx21TmgpS41aVKeNUB9te
gqkWjEtReQ0C6A6bvoEM6TZ6smhc/bR5glA+eTHo9G+Ib58XTwa14LYGl/ovzV5z
6PYCpPZb0d+fIVb0MdH1h2blyUEDjLCetipzhx+nx2nPjZa9F9Duhp3E7HME/jxz
AqRywWDTikkFl1sTZAhcHcbNabt7yS6WL2/BJVXPEWaq5e0G/0i0C4Eo1nCMnNzl
6GwwjTfZsxu1eAFuS6YKgSj+vMYuMGeTlo9LmIJSPFKLV1aAT2UD1eut7TrG0sgL
r0YfqXgDDz9n6scOYSyM3qRn134mPB4K/Dqc7UHc34VK3WAyNYKlYEGSIvX3+vej
eqApw33PZp+OzK++pjAwim98CoRK7hAPIrkI2lr9OMzYn+n3VNha1aS39kqOianA
lxVBUlB/ZZsg29hKM94hy8eUFaDLlq7ZQmsjf5UQPVghkXol2DMMRAG/1KBeBq1V
D5GWJiPxFwTweY0vqEtIJn+biOXIaR3yBmnVCCi7L82tuaX6vEBeQlyux/RVGjK2
y77T5FMWSkcvsyLnOVwgfylCyUXLYjbT8j3MMHQEc91n4elVvjnWtXfXy3uSeALe
uMPxwZpI0OYit2Bn6f27+tj3yP8/MLkPD2yJANHNciYTGb+znkZjZHo+e1dEuI+b
fOW9R4WEQ8IWjw7ZCLAMkGiq0ny6JAF2T/510GCWAyGckLYl/USP+ZORZxwwI8qX
utZOnQ3j9GkbH4oifWvXp2x6trx6xOMzdi6aqfAQms0rh8jPslVtGUDGcr/8s80Y
m/f8x6Ljy1WAnu51VYNwwyvGftA0empzn8ur/2E3hDs1LnNObb6qiYbGzW2Q8dHO
JOdvgoXTdxzXCqTnITPusWEJZ4VFrIr4C1D6o7OTd2Q8mPaIPP3Vs3GZgQ2QcYQc
vpHn/DKLy3bZz+2ceamT6pkAbQGp2h18c8epvndCx2CNfprYd7VnRwKjrzMDyt75
b+sGlTh9XiOEFwFdkLdd9ElVLRlCMdRrbZuBm92pJjhm70ChdtyjO74PTRz2+D7M
r6K/5+/kwCF1gisaWnGTlTuEnrtm0XlOs5YoQWBNrlsPIOkLwcQ/ZrSYxuicgVtS
5oQ7Z51iAiLNZriCFY+3FwnhX2HKVqZnCMv6xK+92Tq71PhWy4Nv3kQ+7Clb5IRz
cNxsJzEbtLM97HUZjHabNnb5RkKJmAqswH2M8TIufv3vB6Qh7JPSjnfBlZfU1sxf
5/0jPCemttP1qiZD/AWb488LmSpClLckPMXJf/IuT+8/aUwlVdIyfFeoRpEB0zkK
FdbFAJqmo0spatZsTJUtmYHcMGydNC6wBj20V5PHofEEutvnuknxGch9NEr9SzZo
DxWegSzkLvJ4mYubdBrrIrDMgve39DIQw5AfCbxocmNjXtIxPSUwm5k7bUNAnqgE
/R6msL+8nCmywZwXMcAaxA35/Hfek/OshHTrcoYQmDSdLiktnOTgk2dSG+dR7O4b
9irIOG57iGCEuvCUqZTQ3BMC2lkaiNq+PJHhI8vCBvTbwFR6NihFC2J2MMtp93Ap
tzXOUghmKOvXNVCK6FcmTn8U5T38qiZAoi59HFwCK8SSgaYiC8S+paqJx11xJmvt
T0ifjEBWfjznXLv50eQk6odd5HnnLFMLz2dGUyZfnK0IA+vrAmZFAo6UIJWVimFt
bQzP70TlMOJdzUxeZtSOdjT3Sre+ympn+/zSvKlmctOo9lbLXFmxs7uCHjMcZT0F
SPKfmVgxTT1AlZtGdZZFk0qMXvLlVaT2hzBt5IyEQaE3jZXzFWbB+Lyvttk3LN9Y
Zp3LTOxUM+0c5hbX20RAr69Ii7pQbDyXWeNpPJOfiSpmfV1TKrMxf6izS50kOj+a
I943qbm7IdCoBRJaPzfW3XOD0lxsfepwHcQzwXd0q+bTpygKBGWr4U2xvWDVz31z
wtYAmi6UIn2RJT7fMkMdWwtuHpOYwrz9q9ZN0ThyvsxVL+LnmE8NOmLdqBqJv6KA
0gmVQs1wOSq6DOjFQMMM2fV92OVXXRYdy7hWqwX/AhcML7uY1f38UeiYojj7u+JV
yqEqobnLopWRD5kzP4XfIqpu9uIOh6Z15m+DjWUmrZIighOcA5b7BXexefoqd2zO
FBunCaW2iSRppDtO3kTE9IEznNc2qBqwcvDeEo6rCWxCLTGNuzx0EHsGzzDQyCo4
7J/k+fxpI/TM6yaSGclyBinz4qS/CVXLuhTOPfjVzKDikkW7MchuXFqnKn36yL6I
WWgOlouxDJcmWWMuOUyAhEYSVa/7otZcu/xkq3k2EoWNmQcL1V66N/ito6C0bhMF
/eT7o0mX/+YlgvJS39rlFXtPYysxYZF7n2HwEwDXpopxOFR/5jbXAX+XRhO8y4DE
gKkyXfnsCGZcdyPKx4MQW9ITaWXGDIDxJD3/NYcPe0yIAH5YGWVsH3Hqm415dkux
Bq+Epdi/+M4i3horhL7dQxBG8+9eNju32pBVrk5ddMUGxhIPpwOUG0wrElmRxnEo
PdBaqEqABrF3VxLGqr/Q4obZ+3rL/rCG1PEKPFOrurMp8AaVmr96ceHjAEBQKJQk
gVCB8/8+FjHFHkHqJTBAP5UXX5AUw6YVDKxIIIKkWHuc2jRzYiYWwc0hHfBiA4me
7YXlhqPNk8NRbVNShjJRjqOqdwYANMtTgE0XAs2/ySUBSVZd42WANmow7n5GWGnR
dcCmkV4FEsWpSNhGiPvEnMHKggzoF8YRG4+0WQV4DqsP0NOC/++o3C2c3p8jBj4m
0XGK6duOXTG8k/CTd7x7bp4XyOf+N4inNYUBIj/d8wwndZMz+jZPqV+3dPF8LWUJ
lTKOGhBrtzKGarpXmcPSKkQj7dyKF6B1MvV0EB/f+s/yD55k+UnNdCztJsCxhNXR
TRMvmjh2fWF6SelucZ362gawf0Zioyr9jFkGPG9eHI7rFaDNTmkUNqbI6qYAqgp8
lDxCjC8Q74TsMUd3aVHSqb767Fh/7YsLSDZ4VenAZG2nMIyVkjrTewycU43Uekfg
NuypG7LG+XtevYJBZOg/c43TenxKOHX4x/tWQXmGL5hlcC6rq2hVloJx+X8SVKqp
IJ+wRdf2JMBaAUJ130DXrHpNDTf5b6+liXxH5DGkA0MuaCPpHyBdxm59aTe/OavJ
1oqsI1mTSbIJzDX0o2fARYtjaoVIutngm1cN7qzr+7mJynMN6c/VGk+M7HzKc6WH
uLt7tXZwaOAq77PgsXqHUr2DvLzQsV3zMN4G+cr7ljXlYTNo+ofb/tNsMaqdsVvK
ywWcie8vtCoxhh/45nB6p+2z9uO+x6HJ7VeDFt7Z+KlH0A7N//azS1hbNmRRt9St
wQXW1CAhT+NtQ+e2g3e3Hfer13iTQyARMRIXQzk3fpLzmnjzATF2dGTk62XBOCon
LqxKktnevoR4KonYmdVxJpCMbSGK6vwvSYZskO5cPR6CGZqpO6MD1Dz6395Gwu63
U44JC9ilyKeySqoegLkB9zweiZ3GKTI53PBpLjaBe7c5F52wjdlapOkq02ot46s4
9YvZdmDgnqWvLX1AE3PdJguBhA0HYccCriv9zt2gATFZ+hEruZwslFDiq3mFH9xk
1SsZaxNvt+IE7xaL8fyRBAC73KniDwtfzH7jfuQ+RrNJyqH34g3Mt5Qp4MYJMzaC
nV2/z0+zLWyZPTl9pxg3X3+9Rwbig3fgIsHjNHuj8LjHz6PlAuPS7qY6sIbwAPVP
maybDUK6CD2NAA9k/mKaC+I583k5bYIHr0Y0G/fGhg6agZRjsLd4RDpIQCVt9xRq
gfg+KIvo0+R02KGk4M0v1SUFbF9APshiHS0u22fIQmNd/LysS9BbzHyi1jO8/NeL
u9QRX6nQJP4cOtdvfqcdkK8Q6TQi/i4pJPhiUj7mkyfeAUwqlaUqmlXaTV6nJ1E6
5xQBoOzddAysKqdGjIkmG1wtEo1mBvmIsDJKCmhBZjPO1V/OKSZAX7C9P41/v9lx
yC7juXtxVI3zLHJbA50R4F5egdM1esPRKqXqFPBUG4LKaVcr51Yy4eyjYZuPWjiY
d9Mf2LImfeP7q333bUkGIlJr7DX5Q4nsFPBVPokHVZgIFdKBLWaqCsZSt+5GzcLG
I6Y382lvVB7olFUhWozLQxA28BmO6rP66Kn849UDk0MYfSr/dtxVJg9tiQv8NTcn
KJK5Ok3yyEmO4ZCV6efqGf1ASRIZ7VXCqx66fYiBKE+Mc8Gz9RlgrYB4PjdjDriG
prnk5WCALt5A+TNSp5UQcDJRKKwPiCYayJuqTRySQHpVvX9sktRbemR8N6O4C9tS
MByEOomCi9Rx5nMyGQBWXwN6LXL0GYeczA7/3JWvkI+nbzGKyoGZoxP9SuzNLAd2
vnfuQypEi8Zo45f+URs+hMI5GXtoCb1QnvSQKbJqSBbd0XfVduqPNB/FsStwJXkJ
pE0LaN3zbXsUVxPXs6RZKaaUvVK8rSUAKC/6kURX9xGD3upsza0i7cXCZpC3Q6KR
nn4OIuVJw/Xyzg9uIo7eget3lVhXcvi9NaVaAB7tS/tUSjEsdYrn8GMcEpNM083E
kov504hebjmG5vr4qUzwoMQcLdEvrP4fdcjR5fLEhwDkmE8UeHeba18SbZDQ5kSI
IUORdt48DMBs8WUdhdGCg7WKEqUKE0IGSwbuE9hJLxX98YykuWKqF/ZYNL2/tw4H
asRQstnQldyUlimOdrr8uh63OIydHUKoX9ZLIKtnFkBiz2v9zS2oZ5B3uL6ESQlQ
rIpDhNLwYrQVVg4O1JwRLd+BV/J9qyaRpvWyRGN6eVDtPgH//hfXwVsRsviOc1gT
IhomRUnP9Od9Siu8crBb3kx6s9IlyjOMbnlQczDzpkVtOAn5sYQyF/bz6VPtpklY
shjYSRnkiSWK5R/iKsHVY+soz6zY1Bh71oQJkWXvi/MdlhnGMoGBlcArgW8MfDFH
tkvlkYATN0Da/mGvh0HmYn4ylx7lG9qm11R8+DvW+IzH/z4818Ni1WSyyZlhbzgm
hXbDfWkJOH1DXdTKskSwQtRT6WHjWNWflhSa+/5J0bWJB+klWN7wlFkjvcQQfoQw
pAFLigyPDHdsZintAaFLY/zbAi2Sr7tXU737Zx14UwvLYSe9XnXAMkEkEuCHgJwp
nuQa8bixl6jshkHMY/9eRjpruGAIKwpObVqKCYj2edjTuY7gWInb4ODQooSg3KAD
dr7qooYkiFIF8tExuES/J+Q5QU7j/foKz/W3tzqpiTR+TA9pSxaI+KMz+WL1rpbX
MbfyDEyAkCU/Mi8GvPaXATFFeEK0J3remYY34Zw2OERyjYxSm3IveV1AdSKgdoCb
fg6oyiIf327n2IhhymNkTPKaVD/nQtgAoA3IUYcvAk99TbKHHJ4KQ7ioNGZH9ew8
WTzebKZrz4ekgN0ioOkkAk58Fs7a+mpp9aSdgTvH3vWNOGi26/qsgsP/KF89z7BW
QwBkJtJC1JFYbDIV74hv5CuXSKpQmNeNcIxnACJopqOcWGgxkyGtknm49qXvYzOB
2WSNO/2bHaYP7TVFk1dvAbmbBFfZbSkRU/Htn6RHUH369j6YjDXD4sIewdbDORUT
wMoWHbq57tWWtOcUk7z9eN0H6WKd7jTmfRtJkzi0ICFSNkCxmiYaBJQ3k6fBm8FP
GKUvx9T1Rl1CovSeJITe+UVl2ml4vNpI5gIpNyUMsuyQWOdaiML+yV3TBMVz9wIP
YBhGLEcoBekT0aegNymbP8jn76n0WNi6qHGSS5vfyWk7X533oQQiZHPDlUXcmtJU
JM+juzzv4Pzuraza9LH6qQ7YpyelcpLL1y3EoCejwjP4Li/iQPVM4Q4Hgt0g+6br
r1144z9HpaiwT6DYgGxMcRKTxPMy6HUY7uNat1ToPz+0kjs3crr0xHRSRTXpSBVk
kUsEXEQAkMJuRQNzhSFz+WQL+CM449Hp9Nlf9iIUuMgBOj0LN0t5r4wbLFjcNlsF
FTmn3rY25i6pQy7WEq7t0pFbbqZFmyXHiwZ6bYg2nDwBM6r+pbk/6qrqL0qRhFy3
rbnXhmAFtHx/psl5rTu1DCgNGEcAzcIBkNbdQja2+9JB6QwCGYFBFkgWNDddjw12
DGtzIyS8Ikrwec6NVZBztmY4w9UnGGHxzWDJONBKZse6QPuV4h7bn6va+3sSLYNh
E8eb5Egmxp3F3tCPqCnz3j6i8+/uQHRTfmGHGv82lvslfjJ1qHLUKLmJecqcK6Dz
PpW449n7s8s18a6ij46WIx7EWqmjMrwnyR7oCfVlVJVt5Z8gpgQzAGGzsJXwXmYK
WsrZS/r5J+fi7Mq6/Y5O8hC5cBpSrqCrJolqA1T29+2TwgAdG/BzaF+Tm26+aeWC
NiNEnsYlN9Z4/7bC8J5ytvtKWBEVtyyWOGzCe1xlvGuTg1Otsu2xF4dwzl9WUtQ5
sGSG+YuQ/t0w/H1M2LH30A0ha3gGzMstUcpJPk9XSXxGG2FTJN5h8qNyOlIlg5Bj
E/1atRCryXMO1IZu1KnS35eyQzPpo9h8BFucRjVoYlNpqWLo7Gg9RKcKB+58edAj
Fi7qwpabOzb9K9AC3XClzv85/rieGfw2F1I/Vj5QumuYUIun2sRAgnWh++nniBr5
JPQFirTtsAWYiEzzRjdeEjTptrBpCAaBiaBtqrNPOMFnBQNw2Jb1M8aBDElY2s7u
yHPPp7ZaR9jxkLDXz2XifGXz+GHdbTndcsr3+qiZ5WMj8Zr81EP+7kc64tqYIXBt
Fn2gCBeW+ScAOOgabbhGxhE2BHZT72YYQc3ftlox8jAXEk0ofhLmyEDgDR2V3jOv
Ex0ApYmErdfKCaaLzN2M3GKP+11yh8zq3jlj4hwA2wpOnigPNJiwBt3fKTZfJ2Z+
gibw+IR4wV4K3A/S0Fb6v6epi9m9OiX9Ee9EIyNPIqK6H2mX4hWpKbx3saOSqwUr
i8pjgJhwsG2NQZWBzCkUhozqLnYSOoIN3wB3GGvPpx+oamJJ1xzpPDAadcYNP10W
O7Ez7s5AWimwDX3lkSdgsRTRqJgpH75B16hwYK4brdQ85S+KeJP6nRrECM1hBXBG
Al9AX8GLIfukDbOsVh24eVnSNsWP4Eb1bSNDjlvT7JXssw/YfKNv10iPcyQmEdrM
DDy0SAimj6PeHpZC7KYJLy7zFCMbUUNR87M1n1AS6oYJ+cjfgXBiPziiHyI3AIt5
h2ZlI1xWY6M/1EGyQ/RCx2VQhq8mcjXJE96+5mOI4USGu/O2kH4Rk5a9SPHWrrAh
q7TDfU4IXh/95lK/+Ky+TUirzfM4RnAA9mzilwfT7QOS55yECn920PreBbkl4HZ7
rkV5VtIzYmx1IrXEMDTA1ykucZj07PERTivzU3vFRAvg+eDmL2QtY363OceQPIM4
P8f6LiPZfgdun9W2nyAn8oeDLAQm7LzHKJypjLN1XjI46G6m5Jn9PQJCIAk9gRqZ
sFrJ3ofTbQLNWp3uZDu5+g8XFyo/T3Ada7tIDOxJJuM9SRArqHX9MPqqz7trf7E4
Nix+0EZycYyw+MiqDtAzk8tzSTXC2RZ0U9nFk7LSU8VnJxroSQssag7mYo/EfYAh
0nwlCCh6YQiO3CGppEbwyDTWrz0qHaVvQBzjkCSfCrlU3XAbtzJ8j1tDBf6e+kqu
hQ7Kt30JFHiKoPvcd3VCKgLwqaVJjYpXpVx5Yfxkx50lIMYPQdUkBGf2WJ1KkVGF
w4GHR0XvcwhH+fGDD+L61OlawxPzGtQ2ruDPdE5dM10qh3P8Ee9H5nB58UO9tTR9
DUCBO0g8ZIOy0ZX23pacmdegTEzcG5A3nHaszISe+DIHg52YEHWPxk2Cdftu97HZ
6m3qpIZsEPlUzNmMXYpx2HNIrxAUyz6lJuEkvCaH6YtCHgy8txfcRkbvwjkgzOhc
RZGh+35QOOq6pjrP8R6DiavJWk2hw8wWi/CEwK3tG7aHW1a9x0mGPojciSh/gLg3
l5a7/Q0ipmI5r+PD8qO14xRQHzHuICBRzHmojtSQSJSYiIZ0BBvlTCK97CQM2/AT
X+/zwBL9VrrFv8evh1az83oyEJcJf4FNPcFtFSjVPyxm+eTxmrQcAdYmu18rEUwU
srw2mh79Hsz0nLGiQj1+Cy7pHY4hxFkVZeJApMcJOCP/Zpkg+ufLqfc7nmCMGZ3K
wj73CowKXEby37s0UZuOpkSCOpTVLtcqourXGNlYLPJNQKJ53EhEEzK0gni7ebc5
cAtZrBHhmGBsOr4f4VvCANdfSXeT1zqrCFChTC+1BADwJ7A8+eM/06Ci80XzcAEp
jV0y8ryGcuqSsl37YneJcA4a8pNxRj1nUF0QApJp3mL//euoPCczJsyf1WE0XPvD
4lU9NAPucxjhnucQq719o4HbzT180frO7PpU9CtO95R1p8OF0a7UxrZfwqydO1sL
YVI79gLKcvpGuWF6WPJyVn6P6B6Xj7qFTmwATCTRNLumlQVR3F0t41agQnzk0/l4
Wvyo5ZmJHLoweCcvid6VWk58BbCJL1LpGq/3jfaomwPkZqBZ3UE5Yb8fT2eLQ1y3
v0PNkkmSxo0UzthfIzbIScsqfIoq/Lxj8rBgrghXniWfagWRcsiNiPELr+drJemY
+AwI1z9IycIGESHfvXH8EC0dJ3Ltlnm3iO9Hr0fVzzvHMUE4Xeiqdpxg8rJGhUno
vgHmNBkZerule+16fewAkrguL+3jBGbCnTr/eVFmR7rbQYs8fxP0Nnyk90vuuIxX
1kwm2i/vRbh2MnCiZG7oLh5nIaBcgEuEJ7kXwFRKqx/Y/vxEUw+s7A0MP9PiexKZ
CilgsIEGGXc9b4CXgxYsBlFIuicN6K6g8JykKVaS3duA/AGAKcXqBgnTWfpqeeU5
nb+3Lnm4R87U8Ju2+lVoHHNSF5OoAsMLMeGBk/2q6lCO/ZxaMfN3jwolTTLYMTqV
cygAqi3DMloFfS9sQnd8YAr82oWu+rCF8xQQ2O1USGNzbFoKAmG6Q06evagfQmOV
ATScfFo5cX72SKv4eVLfrCIghAsKLFJKqbneLkRyEsWfaNENTE9Te75OqctpuCq9
iRSXmUh+WxK4SkMLWXRx3PCFFse1NoXLG5PCuQi2JDoQrwIZeQjT22tiG5YY6Y35
dM/Le6gziM0n+3PJLWEFL4sMyvyrZPzg1/w2LHQbco6DxLuuwQEEAViD7+/nQqst
qsNruGXRlbThkOZshl6OkX7dd1HDaSX/W98Zp4QAFuddOoGn0YlO3yo/+o7F4TEU
X6iTM3TWEWkF5wZSZImNNF9LB+qgPL2QK+8el1gg8THX/+TWX/38R/ROA/SlJAbo
EIIjQHIfXNkoOT9I9lTqfmbFPUl2v5ax4K3zTMHMewr4HI/8Q9LSloDzavwwBII9
Lg12HIckDby0stFjjjl1whzsggmNX7dWVY5B1F0t/J8VAJFlGDUWKLEhF0mMwp/0
6w21RNjjFzM91isVnsUWY94GxbTmnrOUMt31pRa+jAZb9xEm40Gi1eCuYmAbtQ2T
LGJKRke0fm68A0yL5Cu836hs8Toujp4wvHhnc2xNocXPcRZfiU82MgVrS5kfk+Ud
mSTIjZNl8ASATdc28X+6VBkcI+6d0rGpWul850fMavI0wIwveBgMuecUr/Sl/NUl
OqSpY5yO7i7DwyMwfkIhdrInr5wdORUdL6ufMtvKKO1BQPzasaWPikea8oah7+p6
pecOrjJdeCP+yfChvJ8MlySPYCz//Q87OFzqleqi0lQsjCoIqw8K8PsYZBgKmJQR
U6806wzHOzbCBImeHSpLmF3VujnRSy0ThCqsfCH21tJfP1dckn174EL/YRnUFwJR
pHJQVS4/zp7W0QTW+LdXx15y3GJ/kLu41jEwIomD8XNV38ioSoM+wsc3t/IoZ6gu
4XjBNCrhJsY34OitPFuoffWJm7/W8YEjatmNkXWijtNFqu710dra5Zuwmr1FB7f/
5ZrDUxE9s/CgiFS6x75l8E4nYG41Qf2FPHVfIEYt8oHxAFd4SNQNlK7auwyU1hz/
1XeMi934Q4Hj+ZPmKrRROAOCnYANTA5P0AxflGmZgS9ZvPiPq7lBFdt1QtjZqeTp
WQeJ6pn/qScz2tizSGWVMPkptFPDldEvrgSYW/+FOqH/pXhsUBrmWx4Ebwwi3qTE
U3ODlK+qmUBBrdTjlPLr0jUUlhXDU4tUr31cqK18CXrnl9RDK7DREdWHEKzESiOJ
fiGBZphP7xe1V7QrOwF5YIrDjXGXFZKInaF3ouKHAegafJvf6bx+EUP35bOg7/Fn
j/+RJpIbavNi/Fe2Rglc9wHP+xEZT6vjV0G2GQYGCQcsXeH0gx/14jWDifCYukDj
B1AA80Qt31lu4SUpUpGTjqJ0ImkXAmU9OHnYIq+SieJZMDy0UjJ9EBkmnQprMKwS
hM0g8Q9RS+P3gt7PLF15hTp1dCOVdPL193L97CtZtTmJTRII2fjWhROIHdSAfY8Q
6PVaxV0GLBcO2D/ZAI848mjRdKe825qxsoyZjwBWxI5MBVgMyatx3F6j6bBVAdHx
JdjbeQrNwgoFEQWAsw5bBAJivvE9+jMSDwPZgMTazyatlee+rZX2YP1p1vn0RV7a
QC1g/M2aCpQ/7U+RURnjIAwpK5MdpxHRnTH/sShE2jP0QGo9cGk8UoIwQIjUjkLu
9aboCmiWl/nt+znDL7VbwaeePqzWAKfREWSMQFPNwDBAEz1cDFyRAqGLfOwA0Ueu
5Q4i2Rfy3oav6RP4+5JPHsF2dZTy3p1sdbTEl6xz8QoMu8X+tNwMfk+Db7acbGh4
u7SPFiuBK0g0NMMe+HcKkhquliPQoNOWrJviS2C7DwDqsSdyeBETkcqKJgm0/qX7
WkH7NAb/3TRZhqqLd3rKwhbz1FRIOE9VmcZiN/AbMX2w1b0N5y0H5o90/7zMcKTV
tgA1DnVYOyCB7nDNMlgoFG2tQA0nqgegItMaISF20AmjD2fobumBPgVCd4EEGM+1
pRi4w7waFzlgYzo1KEgj7vZySPBAU0xSLb10ZIRow0rz4fOR8MRL1SgAfPrcao7T
68Xfk94pwuuRV81HNJLjCAGeJrIDUew0Kct/JW0LqOsXoiW/tR/BwZLxIs5NRFTp
xabTJuauoDsTQv1VhdllzqtPRmJRYS9qmeqd2gtw3/+OM0TgAy6CSmFEo9JWbuJo
wROxt8OBeC/ouDlDOr4qS0lJcYI8NKKPWn+PNEYS0oDuWvIQc43Eas6sExueLL9D
26IzL0nGm1VGK9PFDm+wPjuAL/UNkKllgce6HsxIA5x6n41pmvbztR7XjL7xPfQI
kcK4O1V1MRX6gpcV/40D2xirMIQczFYsb3xxrMxj89NU2f6wCljrOzYA2iuTW6DY
XxcPpZF3zBTz7eOFJOoPBuxO70Nj1Czrl4Ber64NRUqpg8IEjJcV6sh1Lyiw4rRZ
6Ysq8FZSlZut8TK8fDN7Bh7rn6P/xf61ekb5urJIgwI5rTnz8wSgT7MAD7W4GaAw
8bpvZjicbLGiJi0qaDsR/IYKUw5TRjdtF9lv+lTrlubVYjhtwoeDgqk3GwSpTMpp
bOrmD0PL3xHkNrWMlR8wE/nlYJ5ClK7GtYCqzbIwTokzfXMpyCgHSzacbz++suxx
F/YPOjzWGlV076bR7PK5u31DjWERveJ9vvQhKUA7jseVAM1AoXaYN6XmCzfCKXfC
wSmYUibI63+7CsvXxdj2Db3XKgRbhcYhKOVkn9/ppgtLnVjVPju5fMwDvsIV+6wm
gsYIlJKDnVVA5PBEi48GeHJ2vCTHWoB8QAuxgHrmBQ5AnZaVrtgLxXPnRzgq7nHd
gVCVefyQ7RjiAR7I+l9unBPJmnzq+vlxTyEwHEmdAp8ZzF0CCFgzDTaeff4I9N0g
X6V0bfnwMnvdY+a3c3QcP2Plcthve7ExTL8sfyhsExc0DQtUgdVz/uxZ8G4OgyEb
Wv0mX9G7YxY3iz2PtfpEdjdb0tPEen2l0T5tsX7Py7tkYnZx+K9luwC1axg3O0rj
nLhUN9WbeXb7nJUOejDOtlOR03QbnGm/diMvDETVg4bC6DtuyaPh6ZQFxhU1pTRP
pVHqqZiPHv4Hsu5UVBjwjGhNBx3fqv9aZMNx53d7gqsJs8KPweNJylT/Uo9Zh7Eh
DTkY8FFkkyca1Y4BjPuBGbVXVW0uxLWLgyeNOQFVo1agpV7EDNk63Z6GfQM8gK9i
3J5Cck3NvjODR84lfbQNNX6LEtwn6h2gX/qZ4bRh+KGtF3rUEGZpkB5JANPtkYbC
KEynmHiZDrkK4WMsUdHgckE9Hp34y6jbYDJf4bDktNhbaNKvuP+Cbtub4iDfMcsX
hzHWOiSue8RIxkOiywsI6ncB3NmDKz7yev2OBcZ5k1gQsuNEO0TZKjYmstmwFm9W
5uofU+OVFQl40/md0bC029FFqhGZaUGKn/wz+2Wcgqu+f+OkNML1BrlaXJb9lSkr
rIIwPeO1Rn3Ae1eeoxtTtQC1bxFvOACuPb+e+YnExZotw6kZpSaZwQqP9SIJNlo+
xU5U6JH0v10PhlxaARmGAbc3ibeSyhqrQl4fuLBmaW+YA1qDmDWbjRGBiqWCBOnl
G/B49SSxKgh9R6hNR59LDlG83h61eYOydw3sK4dXooGbTznhhLfnMdflycFCohUE
4CwxnQ5eEtOScCx4faaTldv3SpcnSsUjRv56MZdReP8HS2z2SDwm+VDvzejMeDIu
9Y/LOZGLuF0LDo0o4V+kf7aMwvJqa5MRr5x8i5Cl7Gk3jgl+qP83zOpJU/aHUmpH
LA8aR8g91CyAcfDw739ewA44kR6EmcQeZgwFmwg5j+qdsOhVO6F7lG5RipwdE+/g
zBgT4eHzkY6Q6nKph6ulk7iE2fd4K93XvDBrrBHRIuEwdOAZTUpg8jUpH+9oSpvJ
UGNVTL7nIEK4c8wbnKqWAzY4r7SJzsinuZ0wT3R58R+XCUviS+nwmJTmDm+CO3PC
CNtqssYcwOFPnzpj+lvl1LovLilWezyMNzgrVGv1jPEhXOCR2Lx4Q1sUtpFiJVgi
3vnGrx79wVp4E7skHfEztcbaIKlxltg2TZ7xfTPDwO8BopKQ9XUFvSZHzreIRfMZ
jbpm+c9AOY63l7THjgsunKO6r4Rd+r1VxK/QWbme8bkrj0+l5rDaZDHVHg1V4BdW
0FNPz4ML+Q237tJE/fKJ1qGxUFHbK2rUQdQfWz/DYKZs7EYPNF8q92Ejhq+ItEBT
1HxGsl8erLpvLH5IFwd2f1uF8Ak+pYm07yw5EtyRh6D4e7cjp8I4CU5YE6pUr4FZ
TpqzUD9trg2IEIV4v40TcScR3cuyxePtKPRnP4M3RG+TifyPgiCr2zEi4pusl6xQ
/JxOG8ihwa4jZJs0vk6D9TWM3EFw5yyzGLIAgjQkxuz0pA7Fwv4BEfYWE+eflY8q
CRCmAVt66sVK4m8vsymC4V3qJBMb1VuBz7xtEHpVJXIPIa6C7JDijoEfrsjlHVU4
PhyX40i++okMrxrV3tb1+sZZVEO5jG8RucbRQuGlIyMgc3FEBTH38usjvme0LiXX
43ypr2UyL/XMt6YLKaPI4mx8mZI7N0Hl/gR83qunRNgBbfDqH1r29QBY+jzRddCC
70tvV1NAYaXwcLDGRxQlRkJO9XIeXa5UWTuYQihFY5X9wSfE1h2qfv8wS8XxTerW
ch1DS9f8JZ1i6bf2fpdJsQFVHVBaDEvppegKvuswar2KAPAdH+R9OiptODJx7ZKG
rcANBl/3tw8jOjTR6+dXnf/HrbyvAcYCNOLu7amNfLHNOm2QDyyIpluZ9Li0g+Fp
9h7RxvGPhPNR6An4Vm7b7u/+XFvTn1QidHgZdhkbI0HfjEgpJsRskoezIOy/LdLD
dhmJXJIvOUnZZ+yI7jViObOTAxg14T0+PhK2Ua0DpKkNf8FbYuLHFrT0qMQzEsN7
yMKkMDldTLt4nR/kGx1MZvAjCtgjtWSyWvP2P/sGaHJlqaEbLOMGfplib2IBwk2o
2Qi8spkQ1A/mNm/OiMyxBotyGGF/PE7HXlM5e0fC4OmVK23zNqq/uRiIft7JiKIm
a4OgKD/JxViRmgeFn8pygoSFxDM8v7QChWIuAelrJOyA8K9FEBNrBowhQfTVACP0
2ugg+d7R3/Qfcf3yV67YCEMOPK+LpQ0hcnhYRb2sdAEdaVaESMMzdNXvf75USE/0
zh+61ElsgxYpfA+SFMjGctjUHWgpH1pJd/LQnoyiRlFlzu2ZcyYS/h9fRWO7lLj3
282SgIiBwRWMk9PCKILzFl7OXY6xE9WU5lStYFg8pbbp6uuP+A9NT6I2iJutAsCo
WaL9P+TW6vWL7b00g5T3iMl+EWm/78C1qJEh6XWvwNLoZZl8U1R53sivlk//MQZw
iFd+wLBBkhc7AnWy5cR+psYZDhG80S3Pe/FyJ9fOKxJdgbdWtGqm7uLsrwQbHLD3
QtXglBFWBijLY8ZlDY0N4dDJjWzGoxQ2duWxB6kqdAxtfSmNGUWM8r3+Sgii5ZtC
P7aAY2D0ALiqCYa6Ny2Pk+4IfJ6BKkEF92+5kj3QKe2+M0wkVYQglFNrg+tp5k9R
1cRWtF4mg5tk8IB/rCQXdaK/ynAB34jVVYetgrm3oITh9yA2I4lq6LTxPVTvJuFx
KNn0mbWUageJiv2SfMISKNVtHYFj7mer3+wbH3FcOnKeLizn0083BXrPzgDcxp8/
oERxmjCsmLe0Nj5TVm9APtdRTk4FFysg4x6dvmuv/9xRuPKyUuiOID7nzVKc/gPT
q+pMwBLK5rwnpfl/hNVef+qqTkHv06BJ1Q19b2/hH5ZnFo3GJtoQNtzNYl46Jopp
G11aXWMADRacx+oVy60OJR51gowumcmwj6H65LzM3V4d82Ma5VBiZxpoRjDtiXxt
whKumDqsz5xFp9p+GC80Re6pTaCd4ImAAmaPv5kdu2R1S2+8EXhiJSMqqMvvn63M
of8ok8mmAAfPtPWwQITys4NWOkGPb6h88eHrbmbYLlPH8M4Qv/yrkpCWPRe5QQE0
VFjmGpriNNSRh/K6QOZZCLAdFiA5fYWsTAd+JHChp5fGvqTPToH1GR2TrmMkuEI4
I6SJHnRzzH8SDfasFx0Mj77U9Cn1js4wjBOie5KutgA2p3ax1TolzjLjGrK1Jb8l
xgWWiDjU4LHpiUJvZaFG0eCcWi1dWJLJfiABRzs+H0K2YuynLmKPIiB+vZg4X4Yx
u6CeY0oS5+y4nBFypDymAv+qK4w73B0y+i+moJOJmqolv3C5InLW1iktwp6/mKwW
xdVvYBe1oSLam2V762Fnadlc9wSyY4TDz+7iHdr2EWCz/Caj1StJvzq+eRD7zM8n
KABMxEATlz7aKqS01Sp1RwaRZwXnTbfwXeuIKZT9bB+VbGx6kyJnm3KK33nZ1nnt
yeAO5IT0WHbv5+5+F2jco+HIOQ1FHDhoiFcGj5pbbAT3WLKNgv16Az5BWjsuxaTy
YbHOGM4nCz5BGhgwRMWkSmDVdL/fQCiO0IWlP1mLdWwqTT0Aj43pNuynB0yHPUGY
Tj3ta9UJl2P8Q2TUMIDmdaOc9nmGrbuXpkjNXRbFUdbJUYtI16omY/byLP420t/I
TpT0t1/gDGyZbGRgNf+o7K0lxMptZftq+yAt2hXH8zl6GhyZUB7mpdWC9/hNaXgY
uY+J2lG1XQyX28g/0eAyenP1Pwe3vXu7urOgFkLbyfnoTf8LrIxzSregI+HSXeMc
68oVERLgXx2I00pXW9FrR2e2hOTIvaF8cIL62a8zUoVeaoNGyO5OISAJtA+x5XKH
sk/hlTWZsanAlFwQqfn/D3Hglw1UaoNHouUQR+nP8J6WUI4UaHddl0/xhgPCySMG
6iIsjT6IqPHElpBDliWvCZbIQo387wUY1ichfRs4DEqNzcvn7EMepxVNbn2IkDJ0
wz4FOrYM7d/wc1jEnHxWViocCIOPj0egltvz8GiaOmHhgOIKzClbzNxN6dgkcQTD
fhtBoROupzIsPHcIuGOVUT/XG1nhDpFmTAmElm99KXflPIdolt6/vyA+0pafbGs4
Qubf9yXp1UCMOfLXC/3cAO1XmvuX4guWE8UFRg9cv6imxDvMbL/toaYm+t/BOYdJ
cs9QNBP1BxzxclrQddyd0fTXOZv7aaHelytv9k3rVeMRq4rJ6P0GFxcGnuT3ozNj
/LHNWA/1ic73F2GHTFo9T9j9MMrn2oRx7y6i3v+te35Cti4BO5ENGSRYynMRTycg
05DMsT4VOepTxkKUYfooc+ZvU4YFRpLd9ggpeEVrTeSjmEQQ7IEn2Y/hktYqKpVH
pS4ouH/AIwlfWY404B+Cf7tICeeAbdJ25RrobpA/WsSqSMAwI9iTmk1qq6rz/+VR
bPtJVKKrB/8OCjkjDLTGLapzwquFYLsZBh8I1GehempKF4F2TK5Ttkn+c/hoJx5r
uerdWKmbaEYY3cPqBMfnHZyesXcBJL3C10RcHT6QHd/Jw1tzfE0RAiOiHXqsYBh1
4P9h5myGWMwljPUadh7yCKeN2TU9m/F6khKkD3C6bPa39fhD3Zgy7QVIUXH0MgXs
QYfbGVCur8PNJEa1yXlSBZfJ8x+2tVT2Gk37C+WlQ7/asVmh4aHPnl/iuLVQ4aJv
a8KYeAmFu3xSG3I/wUJyMLxGNCl0vRLmS01k8+HTKZ16fmE/vnLQvWbZu7hQGBrG
U4aqgWOx5aIRp795/+okX10ObYZdVUl3csaaOFhx+Z9s+HtWfkSyE3vDGH7blE0P
7h2kGEr/wv7AqMFaIVhi2zHMahZrHjdSbsgIkxv6UiA/ernuhkT6NZv3pArBk84o
2/mJXpM6kTVkNyUJstElyLJrcMXhZtPz/pCMsyHxfF7XRJ9hAnZfQFK7wKee1I0a
sNxL0/kQbmJbjaaQ704qJc03tImmOH4gNeDlM+gY17dNnLj0+br3M0xqn4QeXTiM
TF3r7TjpszEd8+WuUnCSyo1WdeaNoDuTEAHkClE3Q1wujOGWM+eYaf8rljE19xIS
NW5dXrAmgzlsLZuzglc7NG6pYxGGXvb9CAyUPQkbRcJOn/MVhxjDc5xATOajxRv1
Cnuhk8LW/02pHjoSzDbmugKG66YlzDCVaNyamV9DfFUKcR3VnIF1dj123XcEyDyw
dmrQ7BRdyOH8SHfGPuYcpJC/YMMQSKygrFzSmAYnZT+388MHheJaAiXGkk6k3yJQ
YgCXlG6smGDc1RxpZGEkf96PpYBk29mVjeMDxXezjhR614UJm1n36V2FtOMQjZ5+
+K1bKAUTFc8BdQJMICyBoqi3vCjrycXKq30kghoOAdbYxlWyv2hSF84ZLIu/BkN7
tcZH8lnwjNCq6Rqk+psW3wVbJiXJQW5PS39RddLFVMVjKK/cPvn+upqIw3AHDlRw
zmvjBYVBK9qfF7kR04IH/Pckp2aJct/ZXrvb6QVWpzedQ1Vur4oR+06RKJlStF4L
p+h53ru2xvcoxQUJnrEN9QdmQW4LuP3p8xIgoV8UCGSd6PvwhdFNJeUpRJ2pRW+i
tZ8TuDi6/hbBjGSOQqgxtC7nVxgHUnJ3f2fYCCGq3nIDBic57bexsSe+WtblOfeh
nzqxY5+xnDAf51RvlIjCQkMLS9S7RsdOOdpVEm7gA2CeT9Tvjm0+DFtgPfVrdsEx
waP6OmfQnFTKRDcBt7esF92AHYMu0bh5Z5LS7rzfbxvlPyGM7OAi/W+Zmg9uboLH
HNoTqOb39WjGkwIkbpD5sKfCvrDQOHFk5TvIMguk3FY8m5lzuttPjKOX/0LNK+/D
Zkqq7dSxFfizri2S2V9QVxqyljIF9Nc2GkeDUX7L9cDDVjDZ7qvpkv6PhlsRWZzU
Aq4YEGnkv+ZGQ6j10EJ/Bqss1ts0cMDWWnXb7du+UulMd4SQk7yD3uNeKPtvTwwd
G6blKjewHbs2ZfYvunEGf702gPlsJTe9SN3RUbxyrm8V50XbaC4QIrA+CyXNcDQw
SztrJKE4mNSvjr9FaF+8l90a4492Lo4DRw0vxnCPL7rbw1JhUyxJn3v3t7oDONTL
Q8r5ozaTAiUpYAnnfjAbpJqw5LZjzCQDi7vfl9sy/9pMGtWqROMr66Kg5uYI5X0w
DicmTTJdnxHNEP+R4/qsSx7xorr3ckK5BILFENW5drXra9MWhZdno6UjVAQHCgmi
H5n+UZIKGUHcpeGJEhqBTeHZhiW82llDDBUVt0FBg5guyGMvf9BpNtBzCCd2lfuX
dmf8sHoOxfg35EzGc0BpxEOVf+4IQahUjcZWHOdFtZ8sC9jJag3tQyd1qs5wOBOj
QLviI411Ww62yG+GGyosQ8Ji46MUe73wbEBj8ejnYslRujocIfMYle/0fDMAZsgR
CMv0eulwf2NIazuid6DL6xBe4Q8vAsQBGMDpBYrUgA/yktcGDQAof1ovEX9rBZOr
jZwoW0dfyAl6WC529ZKhVar93s+Tq6dK9grtzGi7DTgtl6oUXqxlvEVEEcL2kqSj
GfNwNwXxdap0Pxf1glgY0tkOKeAC4AS5Syp1K0MRuZmwzPmwq2cacSxEF0ho9cd5
OxpNbQyV3lX21424R977D3QwsABq9H7En7EKLlXO6Vkz2C/02PvebDlcrRZtL7SV
/seafzt/EACl+DpZ0eYPM6P5rV2WEoWDU0TyOXnfhRAHM/XCzQF2fiBebegPbOZn
YKJ75GQSfyt/YGZZCSdODOktWgHoPJr3El6uyOtaeeHNNB6pPz0ENoFriupNsBRX
GPM6vk4XR/crxJn/ggg9CJrB+gSsh1LxFanwgZ5j+h8TVv6HGlI8FkZ/49gz4DuD
Q7xs5a4hueyT/eslBFWRgxpDPofF6WVyyXjd+8KFmgBLwlJ6zQXP1Uonbe5nictb
LYChGLnzO05XiwudePsqFVUPbpnZO/82UE5AKoNlDiBZ7Pt5gbY6lJ2CzoKZqlTm
JMNmrRhTLllsMbcFT4EHUbtFjKZkEf1BPx4t/eW0qkfamcpqzv6ZgkWSWfoXrwzh
bKEcB2lFSjvqaWUlcbxM+OpIuUQ+NdS7dJ8LswRruPSNJCv2ct+XV0xPIYkKglRW
1cG0mu/sHE80a46efkQmBWn8KKptSs6ItER1tqiCoquZ0RIgnkBf/x/Gi8V2GpyV
hDjwhHuXnpa+8Jbm8rIZGF8u4iiG+Iiet9wbUTcerSUhgztRUbBEVlrIkrKp18+U
L1U52IzzB8xKhSI5dpYmhvWOJOqnHXmIU73KMyAbU9jor74GqwfbQ88iqaN/DOKo
vYXHfKi8+OuZ3dPEb9t/8lIXd62SAUJsiMzPrkd7x+jbKC/Y1o0/YAJTDh0yPQIQ
WXy5MT3keqXdSZ868FLbGA6lUyBv2Eh9JFfoj3EWuEln4QD/0Xf1BbNNQzb7+uJM
1srycKM9bh1JtKcBo1bCb8USJJa1dRZiRV8iUmkvr/lxvZNfXAN6WIdA5LqtPfPe
Bm6lOx63OuLoUtMXrjacqnYiEwH98jB6BjiHoqPs7sd6sJZ4UQkvleyoZVglkY5M
qTRPCDhLYeOPp+Z0DJxFgEnxrjHQkAaXyKiLPpSj6F2AAD1V6Sns9jWK6ZBBs6f+
2pjdLq7vhvTrEwpk6H/fvoShsGVucm5QLVi+En/dzxJoGxmdx2J2cCCDn9bR91SL
b1d7/5bHizWOO7cph7Z6rg6XaNje/CyWnM+LfTayfZPpnT6v75EaOlgBOjX3+lAH
sXGscAM+UMPrj0qIiNhIi1aHg/GZB1WBnHBmmqGv18lWI2JRGvLzCLWcjJuI/dp/
GYf1/B9KzvgI0rGLY5odkh2EOi9CzK0qLH6jjr+/GdRl7GStcuWWY7Bly6ZiEHiA
hwfWU1pkwDUznTdl7GDgRu+VX0fKZyZtct0t8BWuGKvu6vvDCTKIktMRY4lA/ykY
ys8Ihb2kDP+vJWw/ohA0566fs9TMjQPsNzFg3h48vhRlJmA6xMC6RsSNq2yHccNx
RlleTu53AS5i4EqGlxALGpm9NfqXBk6609o5/UuWdtnwZZUlqa5nT1w5APK19KSK
x1UodCZqG40Hqld0mj29c8cvVRvASzTMtLpsxfSJb8egr9p8mqfL8ZLF21eMbyqo
1Y8K26i/6phGZoxFZUBV+TfHG3gns0BeuWnpCFy3chJ4MVcA3LIl+qtIC7wCqgzT
m6RogUxPD6gD9OirBM0YthqFAUEyctshkRAhTOjALjSOJ5w9f0dDDp8YIEFXpa4v
wBpsg1TFk5l6BP/0dd+dBb2/VLzoX6MT2OhndGe8v0swY8dEX1rIVvZ9YB5BPSLT
t522NyzBqZYidHekZFgd6KuOShMam68/WFwVcM9G52FdbxW2GXK9XTCLuq+UN/oU
sHzkWNFYYv8ggCwMSc/xzrHrH0gbwBvmOjApo3iwxZTJO7m+zOmiBgGVdNY5GyTU
NwDgKhbLGjyavqvBC/IWsw4dz+x56q5hlaSII8W6ZvYPteAXvU5HBubYasQj30xs
3jrWUG2Skz/B9O3eETEYh1AOVFa0BHjuCUbmWQx9HtV5xab1OG+ccAMDz7sW4G2T
07JIWCiRLmcuM7K4sZ/NVvnAeMgj1P0zXFavXxlv4A8f58vof+2JLzEnEDL1KBYY
iWAPO3i6Fw3gF6eIV38HkyXATTm0ye7SRHiGOEkj/nHn/xMXBBfalFrvu3ysro73
o0B1YJm2yFYDsGZKPWg+pZ9xF/SoIvx6t+IyvdTki0115IQBGBl2O1ecGZv32OP7
2FtZYCs11Mer4Z9fVTW5/KzvsLDPgrxr5leM3kfdIosDvEqj3zlkpPng2XKkw18C
D0v1E3AEJFbCuTNNwVrl+DYj7iDCZUc8VPQd+BvxLUAmRgITNERZrCRiUSKzVZTF
DwuRZE6mM2w0NU0sczHLkfwFfUErPH8EB840XAlM1NXjuzICOMKymMhwUW7so5Eq
4tS1vVOeacGdZINIS3bsFWk2JXfR56CIlXzBEPcdg7DnnNFa08t1LGQsu89DJGUm
uOwOj0gQIJEH20aavOOK0J9X3Ey2cPaEisC8FMBYJR5woeUv0yCcQXyxdChO4uoU
nj06FvChRprTHiKla4fyx68psTzqANI8P7wIRjUznaeuHz8Ly3hFjTzKCr2r1cOE
6hQQjqi8V9EqSXyR9Thxxh3itGXevuB9ZNl/FuXcd4MZMTCkEo06R4NDFSP0trTY
wy6p9n0zjmg5/7iDFe+o5QNRp4QbRwuiElLdrY0oD5ojrcWbCh2w8KN0Z5qUynjV
RET1Qg0V4WnMNiwpdUkNQq9j2tYD2Gb1VvsHKtRmjWLwseuOstZeXlJcIH5Szmlu
cOFPVYLqtCe3k8O7SPVZ6RjPQ1L2Vo6YXrvZE2aWD37SoOPbRkZ/4CyFcz+6lU12
iGgtVXlvFJ5VilSAv2n7+5iTs1S9DKvkKn6b1TX1p2zuAoXVSdFTQmJHLQ/HlAkY
eTDFzlNquHP2u4UjQ3Ocih7insR+kPLZL4lJEfWGhZJOqRu0vgC5Lx0kAe6Nyix8
qQUxbvneYTAmLuA1kAhgWzeDdStDqQgo4U1hEEaQ9adkCq/OtfxsxxFJ8sMW+rdJ
KYKgERj1RQSijjOumqKOu9heVYt9piasiGvByN4Sbeg5R0Pqg8MbQk5dT6Fr9kMD
YhIs7QN9D24KbJVkHZoA6C41zBztlqHG4Qm8Oy8YTFbk9qpiL10MIt4EjsE3KVyk
qdUVMxaEtXo7lDTNIDIsI7HksjQQ5R2kZRIM79laDZg6dRVlvHwPCNQklTwEPb6e
qSTxx7Vs2MJXeaKWMitScwT1jLngSpzC9OZFLekzLj+w09wF6e7aqzBAFHo3VLuC
KlHLNBLif2/Mj/HG5yOIkH7IZUw12Qzb8vWNbR8ew4fXJBVBBD2Uvv01TU9N2MGE
CdzelRbGMnOgfFAgE1dJtSErK5/uzOyBHBfLhfNNxSKbqA5IIarhSm1obhswOpBI
2BllYVzK5lftPB00/5f61zhYO8NHEZP5g0Oxn48Ogx8PJ9WUlwYeTGa1KOA0a2Ou
Dym3crrT2XVIHsmNAk7MQqKfFzEq+XrouqqvS/OQi5qgthdSvedIwUU+mAiZGXv0
yAvdjck2xsB7CLeVRzon1Fb0IgfKtrp5pr/KkJycjM1cXdbOvT9T7mnlXi0TDdtW
VmJC9rDRrNME23dNTVcCifrT/fAUXeKa8vkaVR2I+4/tdAHme7Mi1LUrxeIDiFEC
0BP4KX+etriDpKl4wIQiYInNkhXUZSsu8YX7bOmUWqowO6zqSnW6te+LMMCYjynQ
Sab/KSQn+keawEZJG6REwO44mQeYVHTQia+7l1PLdXCWAG3lRoAwZ7R4R16rrsei
nXVQgXf+HIkHaSiBNWgDEVndjCjGcN+k8U9NCiGV7PB/gIJxTGOriQUTi6CzOygi
5hQOrsWpn4W4c7OsUmpDQrPwe3MyEzZq3vewfCFq3G1h8+RuJu1VCkja7HGk2+vq
0pkC88f8iHw7YUYBIDDS9NVYs2ZgbgZfkd7CqRp/lVHIBQjHSgEZ8DU1WNW4EJul
wiWKr9JZLD/iKdAX0c2bLfc4sw9E4uaacE+xOM3tElv/GyFly2J5c8vbIHkp8RDB
fFq0BvTkzzBvy0JmJYuSdsFEa+tPQUpqQJfM0mb2n5cVqon7YA6AKEOT1bi2GfqW
M2Mo5ne0TSQmvIme7Y6I8z3EqNbQtieoRMn+7UlRq0cvwNAR7wNuDJvWIrVvsAOw
J+g5qcH44aoaEHXBunbV+RdTXV0wHD1cZ95chPAI61QdiMdm4OQ5ES4c/qJU9zZw
eEBu9WaBwGZyQCTPIDMep2RIGt+lDDO6HmLjdh5z1wtU4Ohq5TtQHiSERpXqLMqW
MpkCZE5P6IO0+ZHr0d1wipXXqWM0dmKYamfxkBTX7WIx+1GeQ4eF9R8CTSx6jD5U
O8gkzCp38sIZCLrZ8EenmLigbqIP6EsuLI7TZrguT/VCDFWi8yyPYM7iBeth4roE
rw513dqFqhXorAVEfW2A6Yme6vzBGdTKACzlvCnnMyAoq9GRPoY+q+pOz0k3k0kX
jW9jHARrdx62sqzQNLxlIJA/Wk7/jVyMd2M0KJpb7Kz1brEEM/MaTePDM6At7l5I
F6ZZf6GFgpGRVVyz7Nh/2HcWM6B2mvLf97Ne/W4/gXe+9W4iRYw9YSF5//pBKlxh
7+ItmMj3GbTAEjfwiIJy9umvAHlpxWLJTZgTXmbJLfhboS20stdytitROZu4spxB
K0w/lY1mYHcLwzIGekvGANg19r8FshVa/WCIJn1CFXHAT0IcVUlBxfsY1scE8WPq
LBu7gI+YDUHu3V0zUvZPzfqiUQgvfnLLPLTsi/24LFy3xCyELtUnGbbSbgQhg9F4
irtyffO+uQ7U1TCh796/Of3fFIjtq88FfB1mWfskMU3LUrnjUTeoeH1dWuZ/mPdY
Yq337V0UkuP9OF60l91tgi1pBhf1B7ZAsFzY3zmD3+/uC3Bb2poNcP1mrPweWGfM
CAF6Acm7o1GwtAgCcOFQOZtkrlagUfchOzYCa3PNojXQvr0keRVRQGDX8MD+Xkmm
iEqJrceI4HmgP16klRhVLvFC2e2upJ3GeeIYP+vW3UVglNEzDmbGMMZvnDXqlcGe
UiHojA3mpKaoFu7ytqfTwRMnFtFTg3tqlz08f5M9p0t5Op9zBvbzYK9SyItvgSmR
Lz/bX3MCHmSuRv09NVrcvLMQOa5mlhdN7cgCtsc/kDXSgDvgSn6+0Vq0Osexncq8
48hKYBz/3f4CRoIjZfVPaRn2COC/FLRHTuGpIyp4J7mGPzpYYg/gB78ILtHi/wpR
92KndG0UJa3OvsMNVb7KYMPCtsVld1umjH8OINuJELtg0kIV4v5QLzuyutKAbaEw
GqjMVWIcPaZrHuUcfnaWs0wvNhhZv86/lGNAeSBcnIRdPSh0orw9mlUZZ/N7/0Fx
KIv4TN6+TjxSxxuXfllvj0h5KC410MBE8GUgYVNvCHGiO6BmF8+XZ6ASm2EYG5Mj
GYlOxr/AN5riFTUeQBqGlMOEksB2Wfz+CVTCUN8Ap35OpkUIdkIZGgQjnBeu98RD
bpivVT/ECrpVb7fOw34UjXHOnDXOT26qM/TO/5ui+CTI8RBRLPbBTIBrkNAFQxlo
v1+pahS4ngaLjrUvnd1GLendBq7hhULdimQkXNohP1+EEqov4Cz4cSp6gZGBvd5x
+pzX8MHJwG6HmsYifg4qDvm06NAxegavxzcfuA02YwxjB960/U5Mp79AAnphNM88
YWG8FmZ1wGIWtm1zcgNeVeY2rgNJZhb1576HbFsr/8zzq6H4vS8h0vzWnEsvaKuQ
TLs7rxYTYXWv9U0t1x23WPOy+w/6mJsq1SvM1+Hh21TF0AOmTYzADbmWsxgjYm4A
b3WK4Ql2DJOGt4Xq826+/IxtSuf8EfMB3Rt8l93HoKn5Xk7Jm0ttH0f5rpfeygS4
pIdguxipk7etaRHB+AiNA6fmGr38LDoAMAfrr17V2TjZvZV6wnybot5jguc96tmq
SUnIgyle8AJhIoLxD2a/dSDnHvtKAVNFpNrKlncvRcj986FVbdxkdGA5gfyp0TY6
MJUwdErt6xmaE/gt3zUnyO2PeqtmEyhg8LVT3g78e9zo1Cw6WUvFA5Urv2nKRvPy
Cy9V05ymTK5qFZfdH8xDqDF9heQMId5FdZ5drdZbcKO3/VKqV3ecyAVf02GFIuaA
8yLrD0q64Q/+7L4SJJ6/L4LhjMH/dxZ8qZJEGHcuZfgMBSKpxswFPfVztWyvU2+m
oES4bpB5jmsW7EaBGy+Ult0LE0jU2G0rL9cBldqmD1U+F1/vrl3/s95jdr9+1XCp
Jb2R0jMDJVeQjdPaS3tPmLM1utmpjVyq5We6MVH6IKDKqKxT4BV9G9ne6XEfqjxp
q5u+2/KzwXKaiZTtatZtd9qyIK2VkDeCWGrZYuUt9ApHgGACZrwyeosWIeuVKkyT
ajB8uWNSvnrVsL9hIm6bsciIl7KfLNzqVe8JHibGEY0bcu9oJMzpVDNRyM0zvP6E
lI63LTCXAdfpR6Zq6KC/WhtaO217dXW20vZ/cb865AFWe5b8NZYW/PN/aRUJwFru
4TWwjh/kMIa+gcoGz8V+yFWdQPwiqAFK8tWBJGd2mDkZXuKuGnz9yFHx8ug1PdWi
NKNiqAJg5GLylyhyKxThAV8+tQabh9EBGoqMN8msal37pt1exVSzaQ5dPXGvFuKq
dC6b4w3qcK4U+MXgQ1BR2GKKhJoe+glBfahdiLOUDFVnRqZw11c8MJiJ/jY5Cwov
HTUPklpqZ25PsaPBKHxP6XFJssMl0lvn4KGN5bGUNqsVYTtBf6NN2VSzuWU13TIU
OLf+D/zXYx8n56jhRZQFuLlkABYS6zYc5c7dJMN7cjoUWYiRFwvL5HDo9AXVQZMI
RJpdt/Srmnd6us2ipYINzgFd7XZI2uTVW9beUbysEH/Rgm1fRddreuKityyDdbE6
VyPxFkypBQSzODK5mHk0wIP9oiiz1/HFkwZyHdyB0JNyRUiveBLq1kz5CQTQDIJp
9xFXxi/m90KgSlttN0SPLKqswkguxE8jNDmYU+cPaxkP5N+EfBy6TwweRBd5Jnb/
KUfeK+dKc6O3HsmyLaixaYKzlASxoELmOiP+TIKFc1OxilIIRLodx+9QoOLqWJ4w
8V4uEoEWeBf+uUNT+iBcpPNPI+GDAda8/EUMgIMii5/Ou/Tc5dugcr87dbWnl9Wn
FzzxX4jiLYlDc5IbOyD63FQWNtt2diegM7DSaKE+fyKt0dUQY6AyTSWHbQgDagKc
WyPgIbMNg/vOKgNu63/Am1fKqpXzzU7womy09snUtLyj6nkQLWItWLiATAJeiN0w
QLrfVxppMlBBbLjW/UtegCvcOl0tAwdz9pg7ST9yaq7czm7kYuTAz4OjGMIvGmpc
0sy2GA9CjjbUYybChaHeFYI7MLvctZ87/OUvKiC2IEjLB9sk+GMX9sC65bMWEoGm
g5y23dTW1qHK+LqdE2a4TxdvD49vZl/dLPW75ZizSndiyE7QvfByhVX9UiizGWxp
l/kYrBWjnYEOE98GJj7p5PcUOW0uFd6FNAkrjGFqFJMaqvpBbxOyAwmZ7PMRwqKy
w+6RxMRIOAPj/befEchdSJgt7Jo8F8USoeunW6NrlenXH9EgieheZeUg/x+5bkW2
1dcZI9mk6+noiT9VCsRhO5DHoAIOReN40/5u9lyBCqK1vr0VsvIaxClHo18bFuMx
CxL9QIngsk+GoNivAcW8JHAl86YF3Lp5lg4+CHpz+jrV9MXQlj/uO+jwSF7Tw5ie
27bSYSEy5a7DlgyReHjQzOrSCjOUv0sL5BF+Eanb9cDOk1avxVZDQqp13Ty6QdOg
AO8TK8Cwjs2DBckLswGYTIh/OZPJVn3G9cnS/Qs9DGLz1EOGFoTUrgFEHP2+IjfO
Spx5PKkvrV8aGfAcCHFdRQSPoAgQ9RhXHE3fe5BUVzXrre1GAYWzd3sjBt8MC8iJ
aRmHy2cavd21ZtNGMkhohmnO6S/PVc4PxNWpgjb7STYlNr2jrHUK0y8eT+PDbKQv
LWZuKNVgVHmlM5nPvhGxQCXQBAFZrpGXOCM7cctjnSB0LMwfIsI9rn/b4vUPQv8M
X7840NipXofU3NN+OK5xIjs7xg3EamgzGlNOL5KDP+vG7e9QzMx1i2r1IYmrAeIR
M1TaHD7VHwGQ2+PYEgnH8QGR+qA9y6nMnH7vFsh+vwgOcj8igFegGKLQJcOGAFoD
dVNY+GDJafBHDEgih3M1IGH/CLTl/73t3Stm5m00ZTH9mdy271N1UNa7PSU65VYU
Iknrh6x0HTBu7GZ4OLdxj9lvc/3igbpkGhqwjH1r8OLcr3dBIDfLMoRP/vyfnrIW
AQr6GkGjJAxP/Sl1cm/0ye8xX6WR0tsrPsy9KQ7AmVtxx800tXVTw/CTVc32oc3/
nQ/jGYlF2tLDvmrAH+vR5OP5mRy28I1Kb+ouk2ER2oZ/qBVjCHRO8DWH5SFe28Qh
apY4iBTpD/IE9+CVaTFecL7ckmRuh+cIhOgWif7eUgouBp046Uio38UX5EJ49Y2m
a7946HwP3CPPjATir1Ce/iAylDDFrPYUdYpijP+RxK0+ST4nFjNH0HZt4vL4lo01
kqJ1UaFTh7TzyPmNsJlcLQSOBg2lM8r/DY4z35gdWlGXf7RZb6aWx82Kb1eNYNYg
29eCrWKQizeeQt12ZItScgSIX63vNzmuOAavzWIObxkXdk0MFLHKp8NknRzcVOdN
t8k8J3dmWgLjU17vyG/AzB/ELWkrmqfyR3pP/87MHMVxVRz1TITi9LQiKkBO+sFI
LITEaQLSVjdk+ZVCQtg+8ETkULOEbY4s6hxcj5blWPdd5jmy6JzKAJQXWv//v1C/
y5UY7xZKxOCvc30Ddt8A+g7xi0LUrgV9/47xy24dL9PIXBPeT8p6KzDydlGWbdbK
nhbB/ZrBj35o9CXqekwWHFvpIx9H8pnDldIHQ6hckmm91mudhPDlYqW/yfJ2qZmJ
Fz1l6k90C6GZpmEi6NPt8NqP/xjaHgIOw1XKzQ0vtu4y+8m3DEEDSEo71rL2chww
wN087BjH6bfvGc8y/MTMK9nBtV09+AnBr9UdNIPKwOrolMMy1NWacLiRcuwUSyHm
gDKMUmRgB32vt4FP0RVVyvPtxLvzb5G2El+rjCe5tjMC7/AsW83xh8NI1zUCUHCw
vCp6h+zm3RbUILKeB27hJPsBH1Le2a3KVqwi8gwJSgDyJ6Ou5OM2norK1VBZnKYu
Y1NmXKUlmE/PDL/yJGjj/FYd6r7KXDh2qJD3Lcwt+da2pwQQ42ZOZVxmAapOyQgm
ZrQ3WIVAPX7J/HRUONJtoqoMOfWjbtgLwcIbaJLUnSJdRMFXAVrBV0uQZ4/dxi0L
saqHwaltWNw/y42nN9uKuPTAABSkHE9ipjSNCvHhBUsOg9JmyJAuoF2HwMe86ZIH
FdqVG9jJHLinCrV0lk1OYbBAs5fOWbGMeFKtIIcbC4d+gV5kQVuvMvADXlDR9nK6
qbKZHCUaDPoHKB2lZdRolYGesXw51SGnYtPYtduYtHa/nXflsK+0a6RD19dJo5Km
NIZ7WRljpxD4OYayDvbmCigeTicUTm75GNRuXPIoxmpO9xldYi81Ft6VqjFvr2Tz
WhSKmOCJ6eTffHddlcYhVnMyin7e0O8VkJy76LlJ+/HpcZN3EcF7qO5KlzjOFg5V
aoxfDVNZbsJclHiKUjj25ITkMc7Rq30ByHRGvNmoscbNIAVfU6ikYLPfXTZYfmvm
6KPxat41FbHdTF9tYulo9pf+LRarKes6h+xLX0QrguSEcGajX8e7R0QbyagwSc6O
KdSVmDaJklq/iwql/eCbvSoqCprrO0i0IXGQfqNHUNrn828QU8xMDOl4TE6fv2sY
CZ/sRJzGlg+z7F2d3I1ad8TD826gD5IzM78JspTVlfMdBnFkismXfOzfE9wWP/oP
n3/n4aFHe+XdjiyDsqR/xFq3Lec8af3lQGAkIVofrOhxYyFrZkMoQN1mjXdIfLX5
y0JR5NG8i1DVqT+qjQ1y80VFbYnBSWOREpM6+hLQB3mjIzliCDUnu6FKm3XL8ti3
xJgdAyzJb6WaO6P6kv8aiz95nLCp5EVqVlMtN8FOZQ8K8Gfq4PKRWHW/Fn41LaKH
BmCcHInF8qbEDjG3jmm7H6Ed8FWep+DrbbT38wmweRzn5HKp13hLvwCnyPpVgBP+
TL0uGzw9FIbDKM77yvuZ3dYWVtu3l+9M2T13CFCSRc8dttbo00ku3fuM/E/xBBTJ
FSBLI1SYptGD9ELR/etZZUzmpup+QpDCo24Vcdq4URWfbHS7dkOfkBfzU+pOQr4J
yTvlHltpkcwWr8Qb9AgtHp8xgU6gPDgsnJ8YUX3t8IR8hv/Ns9fMtkVhP2T2ogoW
B4rHqrmFsIWNLAHiWAnSrOjJtgu0K9S0/VDQJ8ZmeotGwX4yZT20kRx+/bgHLmET
o/zKFXg1s3r4dnp/r1pp/c2Cv/AxTtg4WWbkCHPukuxc2q2kbYtE95MsZAjLpoyd
FCfSLKJ8CcKyQJMRB/ABtXv2JcyiIQAUAe0eIR4xt2BtduW131LuQn5AegwX4mAy
zjxDc8DGL1Hm/CF+tl72BYQD+6+6TjClMqGI24iqt+UCNZ9k3DOt5KrbdE7dBfJD
E2v958zyxVOATEKkW6xH7vy3N9zbhXi9KLQFbt7YZ7dvntbobcyL+m8MCgpQTaHM
cvCWNgJgaw+4uT5EXFE/4VjpunOzZPA/BNVCPazH5xe2cSY/IGVP/X2issSY4gaH
JXSIbn8rs5XfhOKiyRD1PEZR5Kyn4kHqVqkiGCE9lciHJzHeFCH3GlD66CLrFVv/
LdoQoTvBvQHIUpXz8kn0dzZ7x3p8huuHXg30DOR/x0Jh3B4kDFPM8/xzLKZgnnj3
HheJB+v3MLftksuN//JUwzTx4VIb5YtnXh09WDavQzGmcmTAZE0jFrVr0zSTGL9+
0Gna8Bds72ZeWDRhOr5n6aWQy/shYBUXDbxr8WMuml+KW0yCvA56kCxJrS8AvkHE
4KSdg2P8tzHNQplg8uoIBQq9wJcevP7te9sBOBsYDsqUakPfK5P9JVAyXsS7+z8j
jiOORJ0xEF8Jh2Cas3+C1yWaP94zITnAUHdY6mLe6h8FD/bSYgCwQWRmOsbo42aJ
9sC0FkV7ROyDohu/AoEP1EZDamXnmnjY3ksyB3jczZAbOiVbhsymoWUDJO37G5Mz
jM4SuwOq2pH7jrQ7bwGx7HVyDUDGnmfmy0KFfl1ms/zUa1Tl0S2RpkjlrSHuHmDY
lsDy986eTm1Rd7WgjVV04w59+7UBWOt7JEAPSi7rIQprwlKiI5Bza3v4Lsdqmgz3
D5+kdl/5Hk5nvY2Tn2AmFIvNlCpmvKyQ/J+PhFdFo3oAPRybNBD/rIfFmT2Jy/OS
JWYR+j6WPKdSmUXhrXjI/38dPheSeeSLx4EYLQTxXqMsuVfk65xwP2Nwk1XOy12A
BKZrY8VrvjaD3vVO531kaeyo630ngTG31Y2bT1uw9KTBjDtukfOzpguvuFDP1Bb6
Lu7ZFRh/HYv/WLMikxc/PmnkFjfotpkkUC7aNmON+/I/9roXvheJ82Vf5MpDTQp+
2qqha5Uep5OkGYH91rlxjzDaC0HorK3YCwrrOH8WJavEJqc35AOGwgz1AsKOXcdv
wVyV32t0iF5itTAI25zZaUka1m0pdQ6MATRYGzkNDpkHfLVhnegkpYVaUmhzQuq8
FT8FhNnmnSlRabKZ+2T+9I8487ow0qCOe8Q9Ro/yPdlAmtkWIcagP/ynfRwV8pJY
J8b0Zk414bwUSMcMhDaqEeXtVGtSRt8uMBgy9JoUwg2EEOTlSpCIx3ouKXsBVxgx
jrVdUVz64yBzYSXmu4taYqV2VMcbmH5DtQkif6SI72KlqNjle3sTysXemS7UiFjx
IZG7P8Y1cxyGrpjnzpC5QV/XCWuIp/GfLaNO7n9nGaOl6rxXG2nMFiYLAFHx+f7M
olfEUgwRMLESwo+tKRiBLmfX+HPKOVXQbbCvktFC4qiEj+xS723oFeJlCUSSrgOA
UdxKjxvHEKMhKT/vMMntElKwWEGTWq4UJCqVO1AXECr1yn2e4+K651urevqEA5GC
2wT9E6aZUooG1WKx/U4buqYzTc2kYUtFnBEvOn9paZTcu1MplUYr3tepKEY6cqBJ
yS+PtH+AsApearIzTLcHtcTupRN8GmFgTRsOU6xdQM/2mmhyEdEUqt/i8Lb8fTpj
OZX9LT/xQStmrfEFFbdJvKNB9+2inHJdI72L/38JHKH6RwBtoMD8Tzlk/jeRHu8i
Xn5IryDdWb4gNL63J+Kf5r8nRM1S7O0Or3KH6PzlrxgzZ/HCZ3wJcE4A2xsjhUAB
Kt5NBUMgbkY1BA0RhWwfbxs1tl0wW/mY/pnCaWvkOUEP/1nED1jjOGI0/Sw3OWO3
RbTyFo88F76mY+IPW6rXZlBQ1Jv6y2Td2d0heAn9EVybfb6lnxE/yZyW7D/IaXKg
GQX9zIe5YGh9Bgr3l2DvNO6XRWWq/NwIip/5gq1H1TZXJ8ovR5PzmFGuigeXhqGq
eV+m/OEIXcHSrxLqzRTRzhfupvNqwm7wT7AXOZSPLhTAqg1QztvzxpFmLE7Lvbti
bau5RlmZULHwBdvC0oVGX2fzJ3iDmiXlYRsWNlZ+2cvc6WDJIC+cub6QkLgFYXRI
OqlLFJfRkBTqjq+PW6grebqcEigANAVQ2pnSDgk3wWBCvWM1qijBp+Lf/qXXdkER
yjj4vhcU3MnsvL8cZDFVB0UXbyDfmApvbGl6CfzCYkeSggqYIYFjdbSungiopzm6
y95qGb5alVDj3y+o2Qv3Uqh5dAjrs5qmOq7Yk9WpotDeMvqjZB7YUJf4J2/0xh6P
QUrCR+ilI2UzVyLY+CBHvCc+rEhDAsuMDJzqN5Wuz4r5Yof6rKNT3uPVE59UJSwV
BSdNTSN6qVKrt9RXy3Psv1k4rKGHFXUFe6zebhVYb5mvCXIzSJ+4L1OoHh5NRnZH
SHScPpTJv3EmuN2V8Dr9/NPWZ6khGMVAvIvPq/LRHqGN4y42Q+IerjXZ1R6s3Zvi
mrgdJNzRbjYroKXwBrzDCmyH74F41eIzuNhcksFXtDLxVrG6+qiYbVstlhiJrduS
VhCYMAOUiyO3RsMSFGkSihhitPP8QFBEq4Cns57l5hrx/BbWpzfWKv/NxTNkv098
b39XvDA8Pa5CDAQz1z1/0F1fEhjCoCsCfFXiObuNxRBpR4ChCW9SNradGWCiIM2q
2ep+vpNknwWYEFtzXhfSiKnO5RUUMD2phFL4e7DMKStVP7q+4Lrqc7PbQ7gR1RdR
VvRMo3yNLlFSD0Ed+BCI/TQZhlmjgJVLZj7Js32BSDiPnPqZ9eZ6FkzSkeYp2uPc
UQGFrEN7n1Bm7YOe+vt+R0hulhba2izAuAJhq8Uu3c3uN980egu0UnYOD+NE3NQj
hwaSMDZ564jjJRGTttLSPsr3NBJxRXae6M6eSWoYPk/NoH2w5nc2ch4mUrnGxs+W
k2ERCiI9x50gNTb/SqVl3WgMocrtLuHWm9ob9fRMISxyv2M2O/orCyKoH7P1abpc
ppBSDacS6H3bi3LMembIpoAXmvxsndDypAA+sRqSyOoAbOMJ4yRAvh1GrSYWxhbu
j2LtXGxgLUyLWpLCVOcFF4g8YYcgNA2lN0R3oT6mlGsTxCfiBTRzqZ6jYQWawCrc
Iu5PH2FHuHUv9exk97JtS5M3kC17y5JgSuX+i3CpHowYgB0uJADaO8SUr2EHKsPo
/r57dtCqB33Ks07gnD/RihVVKDXR1OfvmzZoORX9e9zullsxKPyeL0BIWLu18My0
G0HSzrUq/ONdpVdLfCj6IPlIEuLA0IIuPALGy1xLWJJLVmx9MCpBI7CMfasFNXsG
P+r7mWneYCdwUuXZyerXrUA1usNXc6Mcm4MEYBu9iR3WQEBXhiPKokarIVvQlHtd
G0Em7JLUuGkbMUGbzw2LzmFkJqsZmPZP9ueizuxiyztgyVeTGpqWaNoqHnf7Z8gQ
vtbQvpM5zkVBsnWXOHiEl4OcxE+rWtDrsHMNvA3lKXz7G38QYDUrmvi48BkX/DyO
sITm5/SPX1bn1dan7dVh2iQDUc3xo/TnmC8zFn8lfEcYWBtainyi/t7RZpMKE/w+
qXJqyCpwZt1fg3YeOjwhxyFQqKF27zSrnlc+rSWUANs16HnjIoqXIqsP1yHvhtfJ
txotQdLXJJmes04LskqBzwmbgbCjojBAWOjATyqBpna/IFQenj3qXCV35NKnQM2w
qYqjuJO2NKArDkLzpaI/eoOt1mbobAq9Eve1cwQQRzzFh36FxpVAMbWt/5m0Nh6h
EKDjGFmV54LEotVEaVtPfQYIslt2F4bpbjcA0BnVsTTRQeTDW52fsPelQTv40F/P
jtUl43NYZ/ALyvb3er0/4QyXfn7auOSrRAdzoCgQCVzt4QdQShZ75ojCgmLqC1UL
n/SNEA9yy9KNDaoN8j8UZ/mTo0NdVtEE1ve0y9+2rNfKgTRaIxSIUmr0yU1oXY8J
xIvEZakdRfHLRQo4WJ6gpFdr9KyAo7nV0NdLUEBqXlR0loXTvYFqkkSCh4gT6Fp5
7uPnW/hwAS54s+uiJWXOun3Mw736gb3KKeRc1QI3rfFhSXDwc978dg/Trxe0/nOK
a9w9EhBG/CYlxYNQQ1ORNvZc0swaNHLrlEwoU0+BqbgZ75F8gHkMTBNYTIFRAXHa
dbzXWQjXyq6daMvZ0n+IIIpxktAsWEADzyN7Jr2UsZgEaGO3VA8rSkR90Bg5wLSJ
RwWqTXTwUP1pLk5jKHzVNbEs7XUS3BwBay/PknWdPWLKhOz3Ebi/WlRKxarNdEZF
/r8KP5qc4gCXqFYOuaEypTxzneAh34ScrBekl22U+8vDTv7JPqXBz8FMVe/UbAHx
r3bHlo8+fYJuuoRP9W0WLHFtwIFe0oXcovz0TtQ0OUzPl1DlnBVE+EJje2cc71rI
6ZgZ/06MQvFsI1RkLn9OMMr1i4c+15msFVrlKd2WUJYyfLsGgHL8xZso+rUdleO8
HxInZ3Z0RbYUuyqlcX+MZLZYtdEMEcrp59ybotTvbF7d/64g5+w4aG8CfrwnGqCX
wpzqfgOtRkABQ8CdD0ccY+3EiqdVTXr/rhRN2xJGp3KJYVydGVk/T6A8L0TlCXyw
CqVkUTEN/RVHZgoaT3dlk6GUQqbBk9EhrNbp1xWr0epeJadH6a64xTeYtUTla+q5
7Y8K03PAsrloykGsKX3svb0prsFrv0LrZIx1Qia1HvLfuI53Grzb/pPNeWL4jrba
JXnvFLqCHo2E+NvDiGKPKTL2tDundqC7qmqEL7+nWE93xQ0S8IwfoHCxfP3jZNag
UThHgELjgHeGzkZUFygg3ypuuRkcRj7siCx9cBrx/87b2MBmTFcTw5d9TKOng8Ls
2yfCWgztmXoEqZk86zlBDFbKxK9KthSOx4RaSwpalO06xqV6+l9uKwwjwIg/z19f
A9H17Wwu4RfALWb34+7K9AIovaFdEzpNnuucM5aYLhXOtoy0a3ziRvjZgR4JMW6W
3hYYWysqYooT3vd6Ksq1Pg7FlVccGXCZb5Uv1rCXOMryr2BJxHzCZN+BjrGD1PMh
hgkR9uvJP+n0J8WpQxQ/JXQo3li89rgw37CYnnw9fNqgbqql/5c+h2oRzHod4qKC
3CTpN2MR8dmv2EnOPnGu/E0INw87N7DrvJh0LCKylp8U6dAwi8Ll4lvsShKiqxA8
pXYBJWdUSbjorkEOm1tE4FEG2joSl3eHcxtZFDFQIZHiBlV6k+kq93nCEbszHyy2
vM1/xrj4SoeR4w5zORNVzL0bjf2lcSLU/vp8GbUpccNKz2wziQnsRRgYmjtbPVEK
aA4x0f1Zjfw+hCINEaJZw6uTFpgXlFiTVcBuWoMKMRIKjyhUMXdTUOWDWUxVHvSm
8IHZXsPYKuER/ht7IMElTKJmZZCwhBq4o1sIIr4cHy+35lmsil9nEZsgk/RDM59M
+9UtP2VtnPcaN1O1P3Rrrbzvl6GmRK2mkkB8axY2QEIF89kZmScjPVgxL3KbVwrI
+U64FnZ2dzHMgzT6sd3/hL5hz4EksTitRtSpAjJj3CFzzRJFw/F/DmfU/d8TGJPV
hqU/HVsVt5/RIdoqDJsdE+27KT4PqUMLsDCb+Tf+NeLowGZpZ5JeZZdnjj5RshoH
YuosmTv9/Di1gmeKzInV2SKKgMPIN6nuxkZvfmcnqPHTFxFH7ZWnYIuuvSjF+nO0
qqm126+MqpE8ZeFUyCgZYw9G0vSrW5T5wjLHWhEXHHsn7XanByyt16DbdbeCN5DG
uMNuwsAqq2b73lzwTxYFX+Eb4e/27lrDKInd0hpXnbWJFyI1rbcNeIiBACd9HRH+
R8XbzbiYR0qi3CzXtkojX2kHMoKw/Zjk7ajQm1H9Sld7F2dwE7UF2rk82s3qLSa1
dj7d10QupxZhj1SiFb4eUkUpLlPy6J/AxSP4Bj0WJeoe+MZvzkdVFd4i1J8LcMH/
r0dqYHSxujxVUjSX2/n4SEYyBfTDXHKkwsMzZw+ufVRZ+XTqU1kLYBCfITNO3+xJ
6U1nHCkgEzXEQrqfilLdYGoKk8ZjiNnrCuCT26BtnawdCEQ1niTdeYwY244AJHpc
Y4COtsrKrW4y5oAjUBhIpbHMIzpE28LAuhubkJphOuH4osCRkPfxkDsd90vUHGg2
jvEHk9RQABkqmZpBSy2e1ZATdWCr4kgIJ83UWYvXsiWIoJb05yw5QpNh/K3LVnXc
MAzs0U3BNoC7kHhByrMkz8uErJkD4hkM8+L4g/0GaGCluobwUTMk9iODKekWz3ks
UnpsZn3exc/GvRsErnwTWPxfhMpSO//czIGIfimyNriC4ttWBfy/o51HiPxH4fne
dc2pSi13nm8iVpVlFhNMIAtOie+24J5rWMAwINy6jeA3+SCUeqSwS3EuSuw/bNya
eSvOzxF1ewMW3vnBJ+F0Hf2NNLxXBDCkwkYjC9VUUcfXJ/ew5dpNmkUwSjZce3I7
Rn7wmY8M3QtkpnVF+1edrCGkP7dRkSHDwXOx+KvN2g5y2+RyHW6W4kpgweh6uYi+
NWepHn0ytUJI0Ilqa5e64nHVPvZRjmLsWwQzOeDK634nwYEsHZfb0Yy71/eEG6J2
zugb6SzNEB1bpUs/OXFHPT4S9UAWl1f0pzvP08v6oJFO/ljdcoDN//e8UNwCOoyG
wixGkBf3AnV2Z3wOFJfVpHzH/LCfD5CTukXedKPbKqqqlkvmj1ey8ZaYA2NxpSwW
LuYSQ650I2GVHS73S2NQyHGE9Gbmj7dT8/3887yh8uBTK/uKHyLYEu7HbK30rXFj
v4yJdP4487005Os3RM4JRlQK1VDbORbDyXGe4UrNRGqritCJ0cQRBWVUrBDwRdd2
V099FMMbQkx9I5WJJmbLxLW4CN78ZODGi/ZDSouEY0o6d71PzoZPbqwq6FdFoScK
KqyTFS5k6tTpwm/Oo33TzLSA91PvYc8wZMgw3Xxkq7BoeqPxn0xx5uihgzUV571E
1Le+r728OLNP9afO92Z8psEZ4vwaIIVXmx5yD/bio++ZOLJfnsobyzB+xGcsbcv/
omfN8fIBKNnBiLMikg3npt+e5GOwkO0mceGPCqsZlwL39UE5AuZU5qxnMiMjxHix
3HtokN7ccga+ZcOZUn9XP6o4F68mEQdfmObGdjHSMLsjA+zqnVdcwO7HnsFESZx+
sXe43l966tV1AxssXNLaqIcOe79q9m8BAgl9YBJS7TMtMHi84rfNfFzXT8J9p+yd
KM2JlDVFsHRHXorZHE3Wt/rj3ikGs0NhaAmtOg3adKnVKQtM42A/AkIYloz9tpi2
ys6GsbEyy7vGBwBq+qwom72vwmiUA2bv0Y/3v8aFlRBOnOy8IG+nxgZqa+YVwMuL
MSKrQFR8V1W8JOOsoyPp3LonWBb2pRwF3n5kdJ1iu1R2tr7dDyycKj5nj/atDVGO
CHhWnOphx2+HbxnBzTYxWb7mUukNqlHSVCrNifEskmaKs4Kw8wJSa7fqbFcI0wl5
TlpVxPFnwyrUPzp1mMO3j9snXl0fG4q7wg1hO4axmDsH3w0drVB3tv4z/julBnnU
nWUO/vta+NJuLXmblBkjaQosvnIPy23fsyHEn6kS/KHKUF6BUfoL5FvEpIgdBIKZ
gAjusbxD05p3/C/EkCZkqxmrknPrtZwxMacchuRzP1ak4S9ZCRNgmuP5Nn4rB8Hr
yQvDt1/l4Ol3aXr6iEbkLFQzwvLbFA6ymjFFBePPc/Knchzh/qX2ORUN2dT8aKQW
0cCFuTM2MdfdxHU7MY/iF+708hRFa2T8FlGWTvvuWnaO+qXWRbg0nKk4UzsWG6C8
PK2lQ1hvcxi/NKI7dIWG+nJGQAst0n7QWDTre8adFEW0FLO7Jber58h+EZWnRMoo
QLwfCBiO1I8TisiOG93lWAyOjLc3ufVcDOEEfAYBI6g2bfpxHzEkQrewFiuyMDl/
VAaUHsDnOeT4zM4f+j2oDAfiAh1g695/Y/MRI/u0beAQY5PRToTqdKaWaTa3xIq2
D+glZL1YZrJrWfgUk8CJCQJ1LfFiJg/UEgQOPCuLx9zWmUwJqzD7qz5RvJehuTWB
VZ4F9fgRX/KBM695hVevRVucQXSJDwxrJKpTX0B61Iq5buJKJqEv1plqdbmgv7fH
/U+QNvP27E+zQMEfwH0tgct0w2KUDV9Q/oLzWF3rBMy2UeG/4sTF9FseKPMHe1i0
WJztI3LfSiFLH7LLJBs8crp6Gx/IQt4isc50EVsfHrjvNArS1G7b7DbZlAtjCwYl
yysNzm4OQKMHGSaBDK1lAQi5KrkYvj1uQGmqCRE4hnHH642sN3skr6yJcqBxX5Ux
JTk0a0I5z/9WWbMqu7b0o6BtrzetjSiTWkxFT89YT8deac/u0eccM8/5QPmx3yH7
DwpGeMDtwoMFZYSWvQJj7rgf2Tf/0rKLy1h/amaO14mgvaVc/X6jvSJLhEKLJn5i
HwNH+Ib713ZNL3CQc3KxRXICC7Gu2Ll/uycMbzZ0q+n39UEWMTqr8BuBHxoLy9le
dtbviwMqU7BVBAR3yTlucPITQmeuMTd71EUJQRwUa1Yf8yhENU6AsPg2rDufeEr1
MoUI6A0GvRxuRqyJVbnjXEOyADILPHMsPKZE5vvLyoBXhILONNimpaRoserDjbfZ
M3vIraSFAUn+4T+9NdizQaYRJSfTbZsTaYW1oQ5a8fBVygJgKusT24MT3zuMDvjL
TmqfLUk61QJ8kPeekEEwOjL6NzshvJchL3Hr6VCBRfsZ3TVWFWMLDrxeZPqlPZnd
tVM3LKY8GGJaUsrJkCSCDOeant6yo2bisCeVYA87fdgpWXuakLqPx+Phnv1MRsmY
1wPOPmt/KR0fVu2gb4kRb6RlX8EDR0X6gAO6Lgk7CZZdbvRuf++5Qig5KA7RT57A
OyJJX5jbHojseKnDR4tgp84ZZsGRxRu9QW1rc24WZ4adVQk2U9NogYYGN0V5zIGd
NwsoZs07KCCpwXCYuHz8YHl3ln8NvFxmvzchHP5ar86OtiLRUXGjs9bt7QcWprNh
IEvdFYwbfkfIRFw63i1aDO8zFPRU7EARuQFLowiXXwQIuqxeQmx8vOO4ZuhybXE2
nZp1lrwVKS4/Lv6Q3xJs1aCj6iMzWNictnNmMoqpqtf/LWi59eYtVrtdyGg1hF0s
iPtAY7tPExe0dV/ZVBfhti9FCm5PHPJ44hL/OV1JD2TRd2fWg0hbLIf7WiC9S8B7
BdAKYUKMKY7/wt9oJ67Ni7C4nLgT7drrwySxs86oo+zideUlffbdnKqPXjR4IFPQ
SUWEgRa3p4UHnuWELBd8iMG12lfzDgDoS+AuvNQ90r2dsLihwt8Mg7Bbea0zfx0x
oPHRziap5bPzE96A9fyAC/WJx/sm0VJJxuz5x7+XxDDbFuwTCH4DLxkOiR409Wg+
v29KnkxOOvMDdOcmq1luPbwSK5/2eV6bkWq5C4DeHSvcnelE0H2543/pHMT/Xhuo
fhMAxeHf/DDkeA/BvlX9G7hTFk6rLZRPncQfxyDddZXcbVgRil4PC8O2NqksuXP5
AfYvg+XXkr2nlnRJngdxgR2sCOZUQTDaspVcIadgxP0kRa7bYPQ2uMuJ3SyRBLEr
/KrH5M61479cKZhkt9KPk2wjgNcWy9V4okFFvSk8Ule9lqI/JyaS60KXi7xOB9oG
Z+JvDBLiz8ILL5NsPQ2cDdEQvdJmP3cqozFa8qstKSiPK+C4DuhFiwRIpFdXuxFi
BES+qgeXl1hTLnMRlI6ow/6YktS0v78GZbB9xfXg0xlQEf5AnIvQOY9GGPSLoRMl
DguaRpzJl+q6M+3nrEtAfVafGl97kXI7JOLfx23fw64sG5gf8G57sdxZmNoDvsi+
A6aD54yhom1lQcxJzvR4Zjv9Z7X8JmMb8eHteQHQzZ/ZQZsnsxjdBHNWYleAw+vK
5qQS8oVUbaoxN4oyGXTBJ4VufqSvJZiuP7sANWtsteBjC+k15NxLg0jJhJg63fTA
9Cgm6kRfiBL56KjQy8jMJcJh7TnPdk5GBws/HC421RIVLGskqL0qRlGt7FpYfZ4u
zY64NHiQbIxuq3zqPfHUdTQjvMtPLh5U58EYptcQus4o2oG+k1bZ5k6MRW8vwx4+
Epu53RTVamAVyr+Ssy5RnV1vAWRKX82A+gg7w0WT5N5GSyrCoKcgsUAqTUd6kUZ+
iYtVmNl/NKCM+eyfFFv5KOvphTZ/kcEYf42Zx9rYQI8PS8m6J2JQ45zKWVMnPljo
VPFZyKv9f2j6zuMbQJ5lWQVdDcnTLG3UaskmehOkVJIhICw2iAscx3xCdehRHBJF
DFrQN4qFD5yzvoKkKdlWWwKhSH74Wdc6B9Wtgj2XzERJ4Yxv20+TQ31/cMifZoqj
kD5n7r/IWmPq5UQG+TU+WhdPF1rS5yjB5viSVEHEyT1xGn/skCQMH+df6+VbVbMS
xY4eT18hZ6VFj+AucqiOUvxQFX51CLSUan/shIBTOXCuYCeq35gSjbsS7m4h/A8F
tFZS4NoA089YKZP5dKVCxKJMWKVNuCRGv52qMpTMcNjzrGHqfscdxbXyQSnyQvRN
y4Tsojd5ibc0hDRUaqdtwKbaRgUy8pPhP8rj9e3sU42ZbEcHY5yCRjl1WYTGafDG
enQdQ7Pr7cr5CJ82OAmWjyCvAifgNhE+Y6S3b5322DEhBSJ+owZYEPskdui+FdEY
8yx86wl3RPBEH+oqG3SSGTDUGf+3vER5EGIaXjqR8HcQzVCrh8+2/OzP1dxISvxs
hSFriDINXmLxm4vXUmbPnM+Qd9MKP3dhBgBk3izWoNDLfm3Vq6zXb22l10mxBjHf
67/51Kuql6ReDGqRxoAWLGcSxuJk5q5mpTAGy0wjqbNh3EDJ7hzEFoVEa+9Pq78i
lnyU0Lgu2bk15Kb/anFSd8QnPT8YY2c8Lls1/GzxR9B5emvwfg5BBkMiKwCh9zvn
u0gd5yjZkIWjaBEr4UdJm15/bzAoqPgqQlAc+dqzoRJqdHJ2HYit0FZJ7V/JAz65
lfALIgJlOiZae6Od2UeN6vujySwB/FUzGlh8EaX2cN4D/1378KNaCZJq0hsiOn4B
R7kYtOQrhWEjmxRA5iMwxuQhPw6M9mGca+COK24DjfBiDSb2xwDvvY5WnXMI6AqW
gKtDLou9s5Q6t6TdkkNcP80iJtMG3wMUfZoRR7hqzDsPC+BSctXorwKd4cKREmDl
M0jitaTWPHoPw48YB2UlmVseaSAQ6480smHmUP2hVQyjrhygoKU5UKelmtfGTKfu
x/1YW1llmWmF9TLCFArHQUs2w8vfwNTHPyW8+xNPGoGaKmX5T/xR2iL5SZDFYdvn
kj9ruDUILg1OqW5NFHi0b+jn48iykiVLNw/pY5fDGKC/wq0y6qpH34U76hI3EwYF
+gO6weO+kV394GFcGDtmQuo1GSAMAAEh4kUe1ikbwR9/A6Kiepf3JSZsFjp2KZP3
zrFzLfnPToeUH2SbMhHSxvzBuBuunnZRNojxQbYs7UfMVlZshn6MNw2fiQB0f5wz
Cvp24efhvjOGTOMNTCvS/OGtL0hrdTPBO3aSSU2DtBZC71DIhCyblfsfWxK5tvHF
Zoj+sIevXBNkflf0tGEY56kZsNtVkdDizbT6m44WmPaGPq+Nd6e7eQd2ZtUNpgzV
nUeBW6bliV7PFzNHDn1ncT0QNF2zqXOUeD+xVjItktFJRY4VVKPaO42yPB8i3BEr
PtqYyFlZxcLZMUE/RsQpbnkwb0cnrzQ+555MvjxsnjMHZHXJC8oj4DOmHCUhDOIR
G/QmbjbQEh9If0x/nq2sfTtozgu2JGkuEfCIOh786FIX811eRG6i1Xjiz+KxeNXr
WB7z6kN0G/mFfrkcdYVVhiz+NuKYIrGYP6gm+rX7DQYgJBJ3swzMNC6VetnhgD41
4uApFgn1RO2jdBTu/CWmwkDE7dv+R/iY9AJ0mOrjdwM0I9/wvnzAzpQ5zrfVaMbt
zLk5DLrJht7Sae/yzFrp5TEKVWfUShh7QuMlITMhWk8tSgMz4Ob89ulQUpY5THDe
F3jCLqyy6520SAbhyEQFB4KmuGyLrHiXtHoe8RyyQUX8rmH5ly/eDPIIG0DIMMkr
OedJpUISv0c7B80VpUe1QwsN+S9GgzRoZRqsRTUQ2XszE5r77EeMJQ1CU+jLYqgm
UyoHpZBJnE4U9shEmpDq4rR96k2JF1mwv/sEqPY/nFBCyYdp072g00Qo2rJbEA9E
7XWjyYIX3LwlrPDpQmSqNoanKiBUdpa5kNjbo9qB39UifiCgYl9tIXoUei5OBYCf
7MArd7EdMX6PFXRVo2pfiMSQ4WrWh6Midyp1ZdKWeyHlHgjLYYiIsY/6eteLEFMH
NQLBG6mS+XB42GAJq3S+mmtHjcsPbqjoj1Dv0uxknfcN4Ld1GUoGp2hcCSTq1YAu
EYgvRPyOm+7Dzbq/kmlBWo8GSlinblD2skH8yM7bgwx0MzOtXHzop+/Aa/y/uFiC
PxUrmwLWlZ35d1cf8pT76qmyyPFm3+FYpjwBPeZntDbzgtY2TGP4IprKjX0Lp25k
aHq1xIokawTQ5S/m4sEfQ032SSQvtlIn6qFaOmKTIHQZ5A7PWIkqm24eb4KT2sLB
3t0t06CUnqF6gWci2t55CxC2yRtHbjRmDZEEuJVTSCsLlweBD4hoJbfgpJWJnyfx
NBlMOb621BnZ4nEuQOPgUwsyQYLWWxas5m/WzbU8C9l1S43+FkJH81kabT277x87
lTmYwd7ocYIbTk4ZpRIS3XUIqC/XS1jWdEHt2QD1zVUNvUobd+xR5dzRtH8u8zF+
di9pbS+i9SWsZYf3chzTWUxv2ZMUPd/+oysTy7Z+4wWHYdfo1ljQclJmJDJ24Ghd
z7pEbvdAndEmaZJp7hA7k066G1uLGc6mcjFBBu6QgxtVmKOQfcEff5lq9L9yUKL+
JTwMCvTMHUf+C1Y+frWcj3SUa6GF3ch+xvzMQM60+jW55QvWbkDQD6THs5kPVcqG
lO1Ux0LvKhol2xAfdcTTCaNLX6uowQaFngijghskDzqwH8bunYbCqDVgMl5TlQDu
QkXikU70GDOzDwlILOJRnl9ijyiGJ11KvQdxM6zOjQceIxtuRAoGxk+YajAmr+vW
nfigDpvqPRkVMWmad8gOy9BW9Uu9R4p0/Lbi0qOyx94Da3VcoEzNhgtFsVt9E8jc
gEuAlD1RabdQE2h43sQncSA/2+obAbzFq98eYMvv5xgul6eFYmWDIAOKGXyO9N0b
KoXNgI7I1B4Jh+og1GqCWIlkZrxhb1nJLgnu4gTmy963bIo3d1zH5ev+mW6hhI59
dejT7lb0wqaOlJ+bVkG9C+TczWk3Fq2UuFTAVScyy+dKmqgJ3Rk1ZfK2dX6/3I5f
hrmLN0LH9mZ+idrTToWMajg7vg+VEFPvpu0babFrLBBkip8iW5PhYXaGOQjWfNI8
WlrjUDMgtxCDhKYlds6M3PrEijYdoQXbgyuO+fPCxVD2zQMAWTp2MtNsInJ4yDgq
8MiVZbYjSaHkQ55dS+q0nUXxief+HLRCWAtZFu5tGQLFQY3YKipqM1jNMd/S1WVL
bUbzJiQK1vuHWAyx45e8GW/DZXsQHXC8rdPNOnIncK5SMo/DW+nNiPTogWAMkcDS
Nys2aP9ilRPwRMD0XJPbFudp4v7nLU2yvN7MUlIhF7bllXzJKoWq7ySI//eVa3Rm
3I79li7F2bxFG2WmqyRTN/0bdjsHS/QO/G9cJOe3z52lky3zLQJnYBxwk+AVAFeR
uOWrWLxGKdB0oJ72AW9CxbJMorKV7MS2O4F2Pwz0sHlGOxxIZT0CDzYp96mP342K
zaCvIx2CJI2oPJjuNASDUmk4FnTw5dO3LsOubuqUillOzMjOCtVYBEsJSi/DFkax
q5C/Qcgd7e50ZyJfOWZSOlFjIqpKsfNa5yMS7hmQM3WeybixNYN/Ojvw2P6ZbghY
AXpUT8pTbY10gLvY/hoR+P+MZOOCnBfNmFlgvavGbrp/uIbUXg3CuhIcdmpUduwi
sE6fD3Bem6mVP2J9mQiPnpDoHrioE/umRxsEKhLin5+j1Z0ayQzTdxWIHcxW87p4
8ElgVTUCPMPSQr0/m3jU6Eq7WP2w2yAbLKqWHubUMFcxQBYtzVTkvtvqtxBDy3PZ
nTi2Pi7quJMKHFWKNzpYMUaTcUqAThLarDwTGd1X4GdTbbOlbvigr7T9ke5+FDM2
fHUTsipeeyoEE1BRzvzGpHo/R3moU/siur0uYhcWcaYrRrgGU/JZqFIpmyPqEIcD
JCyNJhJwlqzqr4f6ZYIb7B1d7GATiQcYQNjQYloOafmDxrKrahcoqmmMlME0MPqg
02KWv6LVOtpLlHrBEcRcbO/26jsv3WV6muXoGGH5WMnC/Nau1Im/yyJ4uy6Z2cpx
FNI4HR6HJG+5e/D1aH+R3B2EB4EnJQyjmz6YxOvKUejUMCShLtVEMYYPXgt2JDf/
p/W531k3dwpbZkqJ3HPXtOT4R7kif8StPEzlmU0Ni5SpQbCUgk4UD+aN4wv7TgGe
rvoViP+NYxvqoL9/UN8FyHtBxM4liETM0bbRh0sS1ld50sX+HBUKfNnjzdtehD4Y
6QgmTJ63kNwz7hIQxjjKaS2VXQVpp8WgU4S7QiARCJrP3wjnRji5UJrHqKecy7Zb
YlfB6AFsi6KkygFrqMouXewUDGvldzTcZIm6gDEkBPwQY6CfsuiLHOR0tXI1DBE1
tjq6JQV0p0EM8G5lt7mJ492jKZRBdVjOBeN/rXNn3Rm21y5avg/NA8mYPXPUKPAQ
ydakGSF5bTzCH/nYoVsUQh+SyJObTD6wE7DZNLPAe4yMyVb+LXhASYhexvFo+QvM
5E6EhrD9QE+kuCuwOUxRpHnt9bQJIp3FsE2uM+k+Uf2MRBz70AYqQAYdIzU5Rp9c
fugNCbinAsIbmmF14o5/qPuR3CdwCdc4J6V30+IEES8F0ZTdXDRI0OG+3K7Qfz7I
ubsLnk9m4YmwhFnM323c7fl8u18tW2TihgFS9eyIqKDaht1IFKVCqnbMpUdIaka3
uSEdTfyq27F2xpyGHo8lXmGGS5L8jq8XnEQkaVnJin9JHrPfIrqos7GCgBsg/Mcf
ikPdqG6Mwz1UFY4kKWkm1VizNC+CVvOlbBKv91BHrTNg9VU7nTw5UpUpevh/J34j
/v436Sb/SpvUP71oiOr3y9yLol6mjiRd3M6acrl8RsT3IG/GhYz2pDYnaZzVlicG
yOePQZoT7f73GM9EB58YoHIC4IFQ/l0JqVl4z/UqhttVgtaCbnKfzh7yHO5miRLd
VK1DYEF4e+3+M2wbdHOOMEMpQvpLpPT2XXfa7do5/jRjBJW/0gUnN3gcpRifs4R5
3E0I8JQYNqjbwIU/Z6xifx65oudWCMeR536UA8Io7/BjS850dCnNOxgo0EsNmehp
ysyl6Ha5ok39r5ArZJrirf4xRY2o0YBvg3mi4pfM8qcgmi7DWaWahhUCtXsFNAKS
yZ+HgiERL2LMZev0G0PzQA83FEXFx/cYx4f8lEC4jGa0MCcF+3NxfxlKeH+Q6o1f
mWEBtjEmSgBGP8ltIRExKVDQkhc7WTWBAxWR0Axd9FIuiwC7iuegaMney3TuB69A
7Nshfml2kQJ8cC8Dh4xMwlDlqEYteq9u4znkmz7QoMzDbViuaQtH+pKwDgG/sJsO
I5bB6bsYOi9ham06cC7y+mEuKj4GYhmGo1tzm5myEhzW5iSHIbfFyXL14wX+4EUd
oPPmkdbdBaC6c7LX7pnx0RR7YwnV24aPl4Tl70cSoEXRI+tKrLhMjww5chevlX+1
938m9vRT9TzRtD4LdnT2yAXC3dM4p/BJ04zJa71JY858EKQfEcjp9qC25L+mKftz
qt6rW+jI/u8nAQR/aMvuFR0aoIS+JHLI21SZxF6h/oI5smYSGrR53yMhrL0NhTKN
K0a0IsmGQankfuNiFUsTug3TwmnrQmGv6yoxMMdFXke4BLcxiB+TuNtsJPiNoswC
6LhZs1UKNl4qVNhQv0zOSdPg6sSMhoYOEnuNirjVcx6QBwJF3LUzF1FUWmlnOxvI
D8SdDCp/+GA6GM9UdFA3VOvURFitxLe4WjdT6OwhPUwLMN50FONPNlWykfI/LSLr
37WDLLIROVTJ8HdpAVKgO3AtocQqUvBejTPF3WNbLZje+ko+dycsthllY+KBZVTQ
EEQKaq8q1qaGCTBgefehQ0MWsTwphlEqpLViYS0li0cUfucBwRQQLBNNA5PEm4VN
khR0I5I4FKriPkkLtiJHHSIIEFO4SATeJd0CpkxHh9sqESDg0fqmShH3RdcnErLZ
ZOHo+BzzdReTFGKPAYRoh3K2+rA+KgtUCtQfuTDAlwD+Vn4UVceQFS/FINDefY/r
aOCWfI8GxB2BfrqYMsyyhNlQ5aScuSrpaiLJ3R6P9H0t9PQjRi/3BwkstXviLLzf
sir8FKdQggv3CNo+0zkAlFyXHiO50oHyRHBv5l5ewRm9nf02xekcntP391qxW4/d
4jwz6j5taKiCE8CzEz+Ya0JvxUNVuxq/MUPxyjDJMVQY2vgJ0WCDRWSS/pxibQt7
mvkG34A5wWurcuSDwOGKzXEfpszz2gL7UJcfX0dzJ5jBY39y5W1fEMEtN/ARI4LC
52U9ony6IVaVusnQcc19XDsift+DSxy7ztgh26TgFJDrahRVmPaLfFQ2KQNVglK4
CQ1PLylcsAodSQzHbT1j6sTOnpfSJbMecBDlsxp6hgwxQ6u6FZqkLM6m9R4WILby
MSZC7xrFIRaf1Wlw7abPBLar3WB+oZULnv8VipLGm0t+WpEY1Cawstzx6LQ0ioXr
TqPkcUdUrSHfAg8MReuVytfwZuLpAdMsqMQ2dULh0T3P7TCE9YBNqG7ohtSjkTud
y5qoogq2lfCl6fkJ8R/YofJ8KbGY8rsEpKb8JhhLlUEVfG/Dhia+Yhid6WKX54yp
oLUqxQqm/QL590CEjk1vH1+tg0IEOhLm3j4svFLPLRVAE7VdfWep50DveTPO0lhN
8hWAgOguHXZye9QAaWhoVk6vaeR+Ct2fngzSl2NtI4SyTkFHCwc//qDc65GvsuQw
DDKPUI/wmVPzOusbCrskNvia6+8H9QLdKdfP5SnZtlh8bkMiT9JboKwewj0c2Gfq
IlTcoaaf4LKrP4WzQ+cBrvYJ694uuNIkQrBNJUv8XJxr4NymrpBt2WNF7CObDJ7J
8fJPXmNy0I4HKrzFCVCld1/HNHCOs9fOhavFJ98cXfgcFvkRbzmkXFsK4NNRHUoj
B7M7LHNn7Pvwy6fkVAsJBPWWzRDr2RnoOkTYvpqaVbw++uJtwMdaDfWXMr0EAWv3
ICseiQbjFlb6mp7+SgrZnEZIYYjrwMNI1Jy50g84BVC/qNrXwA3MFOaErICTQ3sI
yMbmGwCw6/IRBb9QSiKf7e9njudqi2M/HD/fbtZZJFxahzq+pqN9jAgVVhA3Flgh
FLfmeNNt5NI5xA3PFr/VgLbYs9vmEGM6ZU2nDhDQl9fRuNxwvPC805FghGBnLvCB
dy+APrYBfcg3h1P8WS8BTNbWB6YrcL8hYAdTQso9PvzEBGJuWt1bzts35IHLOyVr
cYLd7G2YvNpQEOSsKPdOaRj4HYosUufGEilGSRw8aJwNOW7vFG2K9lDmXdscUBA8
L5QxvK9gjoOiJ34nVK5L8/odWVTYeY6Rtx6h1O5vNRn36QpWL+iMXw4LC3StmOsZ
bjrjEXGYeFeJ5Ql2tvbrt7kQg9tD6aLSUrGRDzGmd/JJO5Wflueu9lKCzc1M4pBz
Vk32hse1mnxq8YLvH0JQZIRwuudbeYDPeHf0f2rbHTeGqt7TsfnxR8Uut/Zh7xzA
HburS/ECygor71GvZ69+ZI6vHHHlfaXAO/YALy0DjZvS+/wrJlaz3uCwlnEAsykc
/whUjAFke7u8EBk6BtKCc8+yICWb84BDXuYqa7Oqek4YuZ0C+xwGl6n1rm64ZIvq
o2hcXeQvAqvqS3DqXPyklV/sELwt5uzc8tFI1vu8nfLAenqfLlZmoGc6jOoQEH0S
ZHROO+RMGFQKxvnSZQ76hYg4q0Ge5vctCfGAAEpBa/1oAXXMYKDh/TMcaVw+CjvY
0eMarkOnEa0U1YKDrV6FBLjG5YFzLN6p1udRH65u/4ghCH9dQjLtnLM60cWwS3N6
L55VKAhLbHMzMyToggEFHdN1Cwtr47I54Tf3BzrnhhTPWb0Kbo95IS3fbElVo0lB
sGxQ3CA7Oj1TryKs+3VzXkAzAFKC8/LLTzDlq2ZktTlkvZivu7R/StHYHToNVRQT
0m90pC/ZZWkp/RJLOdVwx+QF8aiuDh6RMwQHs+vNo15uKkOeHUHVOUjpWgBg5xJf
21kHJCmPYJPJzS37Q6+AwIXpf4Lu9k6P5cYERquW3nlqdA9otSeuc/SgRwoZjiyw
nRmc1WxOijMKk7zeRdjMk+Y8tO80pWCmnDvJrN3W2jEv2QvWrH5xkLz2GQHhrtuu
t8H7abBlwbJVxwZlqt4XKpYteRplLDCAwZNSDTbSewzs5dwrNWiUjB9GoejOZ8Iz
i1sy7JrVrSa63sZV66vdPnF/kMrBV8PUi9GSsoAoy1vyiWYX3XO7vohma7eERsU9
XwJ8RN0x8KEwjd5PNg1HDp734qDE6T055MlrTHnQZKn5JjE8uX5XFmNj539A70Q3
OH1YBpj7GXBUXEUUzZwgUsPzepacbhChmiL118RVfUqmSXJlFX2JvZvmjwgkXAff
F6wb3ll8RJZgtReZE5jKiN8/5wdR3kJ4GtCdgZpeoq3Xx9cgvhSBAKTWT9QBV2CW
gV8+nK1XA1Uv2uUaPfJf/FE1PL0l0yzvMz64m6BceZ4ftxwLFV6RKTqh2BtFbc7W
kWpLloUf3TfUo6Jt9Ap4msJIztUaGTLxzW8XZiuyoIFSbIwN4rZnyMlCfXRLo2wk
cakfPO6R3HGqcUmiH/R/AOriH04YFRZVuSlFmcDJRDuLYTnPAOwr/Pkk7JO4Wb7Z
9hnfIxqPEg/Ol3falnBsCoYDVNHqPQKb09gnQMjfNyuHoZV/wG7O1JnR24iDLCsM
XXc2a3izvDVN6EEUUQ3VxPgk7ow0tCAnQGL8JrQLUVDbdcF7giS5D6/NI9M3098u
K0sqUNSASVSSMbMwtIn/8+WNKYiBNM2wmTM9Qi8DFv6eh/H1jEQqG2lysIMYv9ai
Xn28ONQt+sJorkemoR1nv6mgs+1fFOjK/7zRhXdAMy86CVJh/88ZOmnyw8jjMUyx
PFJrcrivwpJTiAXmQoWcPfR85+l7PZyz4o4SDl836PkswX0PcAvnWbEzwClObr/i
LpDUutBmRgJSR4ALTDJLLw5QCmdEgbtLPy3l8jogECQXmqlDxEtA53fVqo+VOxbK
Uo5i+eRhtLty+9Tl/U+TGIV4elj8mcQZjj9GBr29ErFe7fkbyC5ze3ASL/wzIWMN
4eVJ8DagptT0AgShJpnT4g2jYy2gvlKPCIRNEH473lZ9EE9+KgnPZ561xBuIPrr0
G7l84+qStmCZgF1qDE0KZMFLfZwEbl34q4+h8Gow2G4TjiFyyi3+/hq6M/Q8Wqi2
5dSsaLLrJNWQ+luDcCkukY82hKyf+6wVd7HeKxTarR5R31SVZEz9o9gdl48VaTNs
lW+9UXiva77KpN2oHf10pxZV5JCU0jZcJ8Islw4MWYqdJNsFxHxyIgk2CzcdFrS7
moWGvBvNyDd7y+Pr7uFn76Rrk/0CVQVLCadcQDQ6sI1CqvCIfi/gMd6qZdBFy0zQ
UZPzd4XIlxFWz5pYtS5n/9HCGBU+bXjtkqcZsHFGht5uUNVKDCL2W1BtmkG5LnSl
ZeKV0rT+jB5gAKjJG6B/M5/Kb5+XR1PrGNd0pbUQ8BWg3XFg+L0zRmFKL34e2H9/
hF7+iQdQT6zfmX3tBabv1aTrhC64ohGBPnfqEknhcUUCx546PxxU1+SBtBHfRHDg
G//tRGHCuqzvon+X9LyM40y71kKO9xPVr4onMJuiBRTP60SU2nWPFu++x8j+tmKo
9e5/+BshKL3BDOShvAD2GY5lbCAxPOcm8e7l+2/+kxiRZvmuB0X7LTaZu9qRfgjG
c3B2MdAUQtPA4iTH4lzbPbLkag+2S17AqJ8ZL5+7kA710H6RzTSuXv7vPkQpGIdk
Rx3fgno0YvXkaK2ZTd35bMtN6umB+obbfIH+G5XCGsj/64CEPQ6dsPmXlvLBaUPO
Jb1GKb4pZdX0i7c6jIC9SY+f1CObo8nvGc9fWZjPzM9msbtQiDVfJwSX6Uqi6yWR
IZD6mK+378ZGLRyF7zBc/s9qXUshMAbhMHHgUn5DBYBupz+ikQqRQmZ80Cnt/SkM
798D3uQLzFLV5cta7Yzt8bcuRIfl8c9kaMFvhEwR59+6sM9F5agElw7eMnUdgIeT
PJKvnQe0CXwp8vIe0wH2rUhWhufF0Etk4LielXyPV5Hv7slSlL3H4dw0WZaJJgdx
eVNu9hYq5F42Jdt90420BQ2PtEXqwVp/tsFGK61J3QJX2B5rDzp/xNpId6dFZGoA
vsuUQZTirFA9FImBVPqdzZki8EupQFyJ2ZRINf3XhzSYTc1Wlv/Ze9DSYplCoiw7
0M0r+EsDObCBvdNHhwsC9AwtD1s0kD3odgvu5FAOO/mmUwce6aZoSjL1nMJ8YDuH
is9bHeBPqV7euzP9KQQzbtDacgCb5yVI/gCzWG7kD0zzudnMQ6dvfVUReyM/MWs+
ZAcvWGSiZ6wa8OvEYlbK+CSd2TyzsG4Rv5c3yJTXV884rXjmRlWnKhLaHBvqzr3u
/5fDvWXKeJAFPM2y2hiiECVIcT46zvTG0nWlPaR/iDIH15ISlSWsWSkimnzStZl1
xa9nuXf35oodKTknIWXhyT4zxvGpJWTBBUbkkRzmil4bFN5vBYZV+I9vOlpQ0xIA
U544EX7rnVSqkiMCezf3dtvo0maN4nljOWcqlQ8+tyB4yhE0fJ8ts1h9rWkH3wcB
VvghciYQ/9O2hUaMqghdW4bWCtQqu5iPWM6Pig/sJnqFWqcCzEHlPRR60NSen0wT
qCmw4SUWsVLPE5n+/WtPoP4NjXYRw3MF/4yG/CyJA13RsmchjGuTK8USlyJik1nQ
pH9d5GMxrHOBl7TzUQXLjEXYvzOIe2Ot+wZcHh4KypdGvIs88TO/nYP8bsDCBpaR
rjHYJ0+MwUByQtV7Qe8w3RQq53TrXJ4Svpbkb+/7uYvF70+PhgCmTr3J4ihBCqqc
9IQpOmggb2Aik5G3AmkyyxyHvV0VOS1sBUzQKvCRY1xygyShHcXF1HvRjJM4mu0b
P97fPk7DVPzPt7HKa8DJs6oAcgfZtxUmt5/mLb1vmCnerFSlD03zQrDce7mDCTg+
g5TIwiSV/qvf+akVu0At573O9tP2+Qx0rrBPH8QBU4QdF9FZubAaEOffJEwVXXHU
OLHppNGM1SqM0JNWlzuF0tJStFIox/+fHRPxRxlKFx3hF86yfXq7+tu7DCZaLlGE
nf5H8HsQKEhdmP21bT8HQKwXvqOmPnB1Gq5fm8UC16qthI5+D/7VYqjQpIy0gjmi
cbeNfigOwcnrsWULuZOn9vxUXFidVVhbjAlnZqsKL+1JP6/zbLC42mctQCqDukYZ
MQke6fmjOrJOqu5zTM4tGh7z2/48ouRxgfKLHew2YNDWPdO927x4e9wyzl0PRjrK
0SwBxjB22JHNX2ndTmN8GiojOiWlkikl4CgtFn2mfF29PfNaFeiiQBVe9An4iSi1
898oq47a8EF6GMsYnxfLKVgqwUk0C6Bx9NfpXC4B9tpYczcH52k6nUZsmYoPAaK/
G3nW8Dg7l6cZlX1PNGKgzXi+iVKokgVw69SZgPcLmXFHzMr4DcVepJCIYttZdYBy
8P/Sq9VL2e/LzuMVDmTQX+zKofrrdBk6yE+hUbfdhlxLo3NSGqn6ej/xJebp7m2X
rLUQ+flFmQe0uAAf15YbKakzqgv0yYm8WbNyCeFlpemW4rgnWg4182Ma3bZm7/H9
G7fSKzjhKIS/tONgiYOV7c17r7sxaOQuY9p9Zykn685XTwo/QJFEQ9ocPwEj0JB3
bri/xFsNpzgXXpF9plP0eiFJYG61bWjUNfb77lf1Kn50mhZ+pwhhDOENvDPsSX5M
/GRUyUyK7NJPVn4wub+PRX/M7DjbPmJ0fmsTqcAq9MNDR7z5ccxnGzhpqlSgL7lb
IE2wmgw6ENYtvugXyj3VdQVO0ZMouL+RXT8iHpMu91u8Gk+RwCtQa47yZU8m2PQq
2S97bGjCOo6KbNNgK+z20hsFJ+knx2mTIBJFlOPXuky04Cq5dEI+JUJCbYQ1gJsE
U7GsfronTAm7TpCUUZHFGG2z/jMoCC+WSM/My6EXP86WA/XE/fNt9WUjHqwmilob
3NBLFDdb55xHrEpNfwyhHq+a8cvMtGjZb3OmU+HQnYsFtT+38+EOH9DnBjHpP/aZ
PqGtLD9axJyfGHXaAszMSEqyw/Anr8So+nXbdFScAWJz+RXNJG1r478XV1Jf3+X7
yq7bNVwNerW31o8sSk9R9T2kArrt8v7O4MunOnbu2c4N4Umc8MNySZlwBZq3knpp
F8ruHoIjVN0s0ptw37Ylve+6gZAa9vQlRsF5Xq4qENFgBLlYIFK055tFVRqGdxjD
YZIVZ2CPG/hMtv/25KjTLSD4SI0L6wngJWtuPK3PFQy0l2nRXnufxw8aiHusb8DN
wlAI5B9sT2BtqMMLx4tC1JbfSncg+odiWgmwhH+Xn7/f+rpBNU/4oB8gbDHZ6Qz0
TG4GhmWxokekkeuMHvdN98r4W5P3jiYHPQgAMovLrszp3O4vAjnPx2UH3PLneQZS
YdkLZXx0Fz420IqYCVq/0iIBBttyO1CcyDyGlb5d/sxnjpjedTuyRlWGgMK18qJ9
vKfN/InnxyJYzxPelftL3E4I6p2RngDLujAYG++YTvjAasvFtMNDQmWeQQyXc+oz
ExKYfN2nBBfePxAY63uT3Rh2qS0vWJGCiwh9AyR7X8kkcScxQ/0aZ6J8NRYFBN78
NZGxNWxxbmkup6cBAcpFipXencc4hK1TrGeMj+1TtipExSnWoR41nAxSgBsnfRNk
85/1qeRs2dp/94YgfKk2FZkELV485MEMpJ0RBGQYOTLxnuublw3H52INcqeI8rHd
hNXFYaxMsrmAbvIgwqkzQfRryuU0ww2ENGTHC9eyYjRiZijhRSo9Gp8rVfleuf1D
8r//UtTb4N51XCTZBd4w0GygDDRrb/4V8VxhIqOrOTYR2HH1hocCoizPW0OxohCG
lNn7TxgBsUlSldnEsPCpudy5FmLfMM5OXiLpTQmOLOW3LI2CGZnTGke5NKO2TjLW
VnJjrlkesvJ8X5/g02NIRt26vjMGJsKwqdGPjwXg43FmPFE+3XZFJsZH4Rpfh7BP
x6zQ4NFjmWr0kwO1HOmEhfOtlkFmfzzH4nKSLn+yPpTfLuKg5/h6IHDAH3mAxjBx
6GRaYHXQt3YD+y7dWn5qjCdepZQIDymT8Tc4RVRsAPJ4SHW7rvWVfL85gVtfaYlE
tq2jeUCoJTopOJMQwP4KUXFHtDH1Y1/tjCAjaIPWatPN6P328/JSwtCfo0nZeJAO
7gRwH70RNGyFiotLaW+cv6fYfwIa8GVqHG+u2E+ohVZqVHRR9f7/CALksZFQGAid
Nb8GgiMgpKNoX3rmdA+SIRfi4f8R0Nja1XB3dZdzgIl4B2+JWrAxgXyQH+mgiUn5
YZi7H7ph8EheWu/wopWeyThnzLluADtr6AqXecdS6sdtcUHhlkdytQVqVEQ9Uikf
peBpYN2HgO+hO91FyRoibb4p1PvSr11JKjEhAKOq4IfzsvnGvXdJQ/6ZTtAr+sIR
k991xWN1WYFqsVlwPOjQg132e86aoFEHQGw5cLT7TVWNCS7Hf+L02AQiEWaYuTIQ
Jd9C7BNaT4INbowU+q7VENSNuCj/NXRcNHTaRr6Pd7m8vYSiclRvmVz96PMfceOg
6d87xoaqN7k75nwxoV157dtFN2YVEEyW7AC5jqq2ZGvb/FHdgitgeJO/SnWK2Z2N
RgA7op0evQN2r0iy5ARBGiWBsx2rQp9PAuB8OO3Sy8R2XuIweybQF6hw1EJ+IuLK
zTMCcQig3MR8uBW8ZcPIDsQkr0kJUNI1Lm231yJohS/lYsAIyXfCGKJQypjJ0RVd
RTElnvbLjJfjm0ymLtPnzecKQZ2VZkIVcPSwkalKdRmmKcj5Xtaw2Fd2UcvoHOMQ
oPcYGbAD4ISX+BfhyPzHqxZPGubHeUdbgCpFH/pCbOpHbvzfUjN2S74xlgYoKM0f
SvNI0HTqEZFuRPgzImBI+eBWgAajsMrdtSO9/pccBxUUfnwk9yBZGmOMGvIpIdwW
M0shmtJ20+T6BF6GqvSPHCbpFO+ve26aYu0Q1eGFIioH86xK2zUvqduxjfdNWCil
bPKEmXFrMPWBps1wtMcM9P1TgrpC4Fspmo9XiS4FVl9W8uidI3xrNK6RgtS+RoRw
uhnf0vz8IyNye4mt1wuqsy/X/mD6BUnmaIczW4Quen/ZypAX1eq6ADUxAtgoTiQQ
PFGYwmQdeAgzzhBo46C77urGP67KsQtTBncK/QABoyko8fIS4Hn4NWK7U3oIBfBb
8R4JIPyqRMZiXG1USvL/DTvdWdERBNxgrFdyKgXVz7Faxd6tL9NlSvY7dabEGte+
52vCf0DQ3MtbGl15tFeKERCleRbYDrJVi7pbybXWncoI8Pcqqr3kLFLQEI997DiR
QYhjdnmAqNXyTQ57LyaIwQBZzKLZF9BwYnrVQL0cS8TFAMUpqHEatKfaa0DQpUfE
+/Qw5pdL468wuj3+5Vg7W/D2G991sTp+P/+WUtgTV2dpuZGZgJBFiqxVzLrVw0ai
1RmXXekUEhA/Wnu/Gp55HHhCsqVdoy6vTiS/2t9uplUEpRE/HcPd965+lHqN9p9x
czR9vzp7f/uMoaQRcb1C7jSJTrTBXyKr646jtQOCUbpmiNzK0s+btvYABxbCmvwM
i3YhbHN1/84tM4/yaZPOvX/fnbJvR2pj1r6oXYd8Xz/MDiA14/zoGNg6Fw1yKR5b
2VX9OFXIBSCNZ5nA1MpcewaBE/9VzxiDzP9aqOf+II2/secFKB+Fo1xvMx3IbCFc
b2IeFOgUijo1szNnErBUiWCwjiqSIsxZL8jg0pU/Q0yCzJEFRa+VT/XBVr5S31Y+
kuNCKhJQv9jiV4w1kyGM0awJEQV9yYczgTaR5yvYGaf0rPbvymnPr3im4/lSmkeF
32yHn+DtQOJ2vk8Dr9R8oqWZWb62g4mAN29i8M8jX1QReo6hBxiy3Q/3cOazQoiu
eqAhiFKM05Qa06IVyonAXPWpm9BKfwkeeYnuCGPlSuNmfwBqY3pGeDHePgTlDLdH
rdLVwt4cIHEMZgfqzGA4fgo60OqcoqCL6kYsuthndk92fwo/76pgD5EXi11hp+TL
TDDqBpuiOWku7bOCefFyKxCgrATX2bOu6W0hQPRSDjMvBBwLOOeyqzWZSjtb+zy+
zgvydwJQCPGpykYe6XLEmHFcYWE8n43qCAZtwPgH0p7p5ONgt2SqV/+pSTcGCS4K
IxFVFsGJEecBs9C86JjFmA41YatcIaXEnO9Y71pDWj8z2IqSkO5ABHNoBW5cjpdN
bl6On/r42djaXEktrsDly9pWfhFeKHTnr9kYzG9MGFXWej72CtAUE5Vg+MRxwVU+
06KRnMgxsD39N34DJHxbN02J+/3Ycq94ADf0aZaXbyco1fg3pUDjgQzr612Kz6My
wcWf7mh2iUpUdq33UXqiYVetowYFyUbS9bP62yqwmAXSENIKJPB24Z6ODnuAW9we
wDgwW+olYT3JqLdRSU+EHNv72O5NGgnQ9ZLYKL1ByRFRwQ/QoSbg45NGAzRIjxFc
BoiT9LFAX1m794ymrOy5s0YL56JwH/+an++JpPiomvTwyyFwPMukaHpuXHqPaKPE
GzyK35unbpuGIdmyjgSD93DpIdeovKP68p2luT+pNum6/PoHyc8soHZRNHV93vB4
PIX31WJH55yS7SbcSOXVg2RExDVsakemPvAzca8XHEkSAk0Hva5SjbvS3L/5VMZs
XZjnjJz61Uz4nkib/Ur6vvzz/7xxgPgld2SvKXkBoSQ8gNNWOR870vcdnmcZ3RgJ
JdzLxD5BkkuMre81H4tzysKvLNMuq6lAL2s5OJdedH4iARBQxA255BCDY0FqyEBl
ueNPXAszxaP3NpbCsGBn+wgP0yR8I5zByV1wp/iUk56BPZwYx077Y9YXD0Kl/UaS
EBlzQEsg9TWpqhmdUMTlw5cK5Vr/H2Tz6ALsW//7Khm3XTMLjwR/bwjQTdMK/Awa
/b0LHpqw8W+W1K0v9NvaLKSxCy/ARerYddeumSRb9pP5kn+HWPxFkTJKZihwjUc6
DUq8LafL7H7F2UQLuj+6O4//7n/KZ2GBopiKmKqS0Qv7eZOhONugSoJbuEg3GjFo
0xQnWq3Wj1PwyvFyRMWN+T0rmO4Q5oUKzgOKTzc0Dzvls+UiGPetui9zoC7ceGr4
yBIqbeRGXqtiwAwFXwOnCHQ6XZbFLCSEnsHvmfZv4MfT50X2n2WrThz5hwJNMY0S
gouwORYU7XQm9kK5tU8ZCEAVn31tzHFgVlR1OdPtHUtLPS/eV60fNKZw7LExzKfg
We96EXm9dGsFimYO8ZDpRzGEzKB7mTGZUfkfMr+i66DTVaANSUAdR09hr1t6aEQm
Y3H9iXNXR3XwMmtb9LYK+zUQBmZhIulvrL+NTsHhIiSzThGeFt2RNkXdju1pTJuz
z7+RIaa7JsxfMjjRkrKbcPwZo4x7aYqbo7NvigJ2wCYq0e44d57OH5Zls0nQOM5E
7c92RPr2ckFsJLsqXN4WJk0YQGhCMwNcqZDjD2RAWaeeK0cy0Hzob8AW4sFY5AG9
kc+3+QUxBKehZNerYTKstVZHdCoWiEyuptyuEJufjzJ47vSMLir/CHJA8aUZpCW5
AZpO8fvolzZ4o76ae9Z3zrFWAT4Bu5Y/ImTkXAb4RswQN98L1fTtJ8Ub1tOu61lh
mureQwBa/QusbNvOACmMvFpjIe7VnHJJQlSr1Daxf+If7RH3VfwIzHUI2QtYqj2b
Mt8flEynQzTz3aPpfBNJEnysuKoor+XAa9jadz270Gm3JXMfllO2TZ/3BbEqRC2D
e2a6V5P7cVx9GBkmCVc91HR+vQqrduTWVEeJFDN+QgdjNYEsAIg36ZmfmPyLaLwk
hQhordtMjI5ZkTP+Naq61IE6YQ5G7SGkDr8uzyjQWiZgOHdY1psHIjVpCa00xbzw
KmSZGwI+lO2dlTBI8wXILwXzi4TUeYz1lL2YEL0HB78r88EfKCaQ9obxzY9vj9Yo
/huzDE27EO25G8VFQ7qutrsby1z5BZP/rhnTXyG52CMvo7EwAQG6RS5s3+bVFf22
5t+H4kXoRsK+xcWvZMBQgBv8d2XINRIJvp5l4c5rHaQUDFxefwLgXqFgteEI1o30
fL9sEcKvaGhMdsExgn83thkN15DHGDghbPgfQ18V83obYKA/kByHEpNe0EK+Boid
G0dtXFUMwd2qB/o93R6w4/OtuFXP84ybm0AqfQEFfT9N0PkWiTxzS0pB+AenIstp
O5zhNeF7ep2JSEcdjEuvzvRukX/1dhtdhPSXq1/bBFPYONRP2J1v2F4pw+h4qYvW
gWU5PU48rSCHBHNZm9beYjuTGpZnoC15B09rcRdd1hxVjL/EkILhW0byvaj2AOJh
8q21d2iu4yqcsbbBbEBmRG28phoLus4in8TxHt7jAGXDTE2nrS2RkaAHFjQ6wSDi
XSpaL862vf2mAr7jJ48Oga4LWRhtO6n8Rdop9mIHVsQKyGZltjfXX0olNOk6qIEY
whSNfYXqeRzANDl9vSVZBJUBaQ7nK4COHcvp4eKjTIzlE/dxqLg/PiLND8K8+m1x
NyypRwpbo8nz5L4p/XNt7johAg9ow6l6lGmnIEvVeEOnYHgLk5T7xZWZN5CMjY7G
ht26uokiBZ+FUvcaU8TrrsChevn/U0xiLKI6zDN4GH76GWtk/yoi+SAE0Nq6xdzJ
NmMJRL24Haigu8pQMUzuXn6DQFeH6W8e77yZMjdFqAxJZicoQHZdCEhiIVD984St
9Tn7MqJ4G+4aQbZLSOuV5inBaki3/mwVRwxp/IF1H39EMrLsaQnkBgSTR2+PjnKM
jtdOdVWJp5OmxJzIXsdmj2EjvvHKbDLxlfdvpbXUwuBoSlUgZWelJam/hfPNmY4p
35kzj4JkxBYwWE1bq0NJgyWfYAuc7fEIYSMgIpiOpJpYtN9OaUTLHC9JfEAYfy0m
1i9nG841ClkpPIPwiK8D3SIG6NC+/zFA1Wpv5/spiTZdZiruWnAQkstMg3pmeJ6u
Q1pG1cRSZoR07Ju+RLiLNzHMuhxSlECByMEtDxE1FZhT+VJXqthgqSEkha8ut31B
kKOyI01X4ch9jAcC8sk4bzFjcoravEPP192YvbuG0uFOp7VxxZdfX64eNqHIbHot
ZFgGJmq7W386IbdbQc8/h99cTvQqo1lRCtTJSo3EYW9VHVU2VmqqViRFIHp3FIB4
eUn6/3v8L1d5WpUYENlOQCRbKZQdwV82izvwZC+5EH9aPKiwlolya5fDHmk77Knf
N63MneDGM0lCtdx5cEFkoxHz5XHKWxuLRbE3yz6dNGtSFx7D2QBUr5umWnzho2oB
9vsjVxvUHPloSm3ViFI0pmbTwtS/cWUUoojwbLAV+BNufbeyHwT+LTwe7HMgVMYu
3yaTDpamD6hy8lA25oAMKweLtjOSKqpJ/6BwmnJA5TGogRL3OvxhS58jUlwjprs3
Qr8E81WsPI4Uv9RPy/QuGvPlImBMxp7U9IOmM7YdnWWxHb16VI6N2BuZr4eYxExs
E9bL3+BlrIqDjmPpUn+yL3fR+JJKA2RRoO9hXMItLvRvneeQuyPTst2Lk7tW90xz
fqc0y9dA0wi2AU3jPXTF/Y2hiJ0uwtKgqiO5yFMos/SBYq1a/9HrFuI5Q31Ph+n7
8TfMp87efzNmzIRErsayMVAKcYwF6phl7kM+qh5u4iuKmVNpeTrw5Djy/W5pR0s/
ubmt44ak+UpArdzahm7IlN928j0GAfG1VePkY2126QJAp0k97jJ8nDUQDsDk+4ZD
4fQTVRW/WGAgG/c6LHq+5twGVV2TIX8GOD0v/0/wGfiWj4Lix3Z/V9gXgXsi/e4N
gA4lkJiwDzksB7f9ucCrBi1NCSkRaEgIyNuwQotWL+an7riMHx6QDCSPhorlM2Xu
C+ubPSlCc5rsh3sXFgwfEpz58P9Ov1FOa1uUMYC24oB8dyCJ+c38XTzDHD7ILqnG
A5W1nIVdUAnlNADrTHJOcJPSzknFaS5UcbsYsq/Crt/bU4UAVMptArKDJsyfj4Ck
+Fx3PUgFISSTTLMWOHQial+5OwYuuig2HZXneYI5duVC0z2UXhC4hOHqMUb4JHb/
Zvu+FGndgAJRliwthLVQ3SjoRojFMa/ok9REORzsPPM92R4YWvyXdjYsi1YAhrjW
8bjWMDZujn0YiMuNYbFOhzowH1Y5nHDsCgaWlYhl3YGQDmtf9lrotd0+5Eadx0Ql
R0WMsOqKZ+cCjjENNBrf45awY3GWdBnm4jPilG5noZEz0qR6Bkgo6xGY5yvRgJ0w
KlVr1weeEf+cS5nRzKR4G2T+8xnGtNK0e2/nfPEmNlER/E6pGOWpIz7N0PNUm5S1
+qLk9OCYtbWemQq2BYOLd4C/6OORF9iA0IQ5etwKPI+Ar/7/51ZWqbC52u4BvxsV
CFRksBElxSoD5jblzqn2Nx9aC3pqwyR95YLjleDNO3dQBEg81xFUe5O36tkvCJtj
FtpbUaqt84AxOZi4O2+EMmsoE9C0XwQr77xxj7PDjqP99O/Kk//D8moIIdg9Z1/B
myJQJ7lt4GuFUiABrXjlhfNXo2/prMb6BrNQNkjKt9kB5+8UQ9mJM4P9vBLB86RS
AfgKiTGywNIqJsXdrXJHuNrIsQSihAOGxyvXCByFJ3CoZL2uTmrEiJNgbPc8fgiT
D+C3KbP5cb2BnUlhF6HaJrtLchfA2hDZdflHwBtF0j1/Ae7K5Z6BvcyqwFk7sSsz
UjtE9b7r0KYxg8lXKgKslAIPShEC3FUmn6Pa2KCz7CjhaqfyXZIh+guYbp7F8gIH
1VtCeasauH1BvFmIc8L8soFRxWlzYGjHq1cXdvMm+t04Dqj5wWQINtO4AY57pS2v
SG4rf0Qtr5wR6KuhOATB+xjFImVxr2hhbmnq8om1Xb1GvXsflPe84pm/hy5uxqFi
LDwqotac7wagYoK3BW+gojkLRkHAfGIYcjv4o3cSnNtBMrlO09ruNvAhBH7vVlLZ
RCxmH0fmYGRUgFzoApifwJQvoblLJxo+KviAYIETJOtsQiFiWPXBLUagChBccVkz
/CLb8o2z7Wd1FJoxkg8HP4NYQIEw8vLwlZ35uk95RzbsE4DzUhn3zmvHb+68XnmA
svRZANP5F2X5ZMqyrFSJW9xMY46TzPnIUQcwN9m/bsE8GmbldRjFom3HbWT8qs/x
bHIfAy8Sx5KYMYlEwNQJuPru5eJ5JZhSvWt94RhT+M7k70QI8z1Pe6AbxnGlN/LT
AEc82he6nOxx4m8v9zlq+Qddn5zwz3eRCooB4uLkNtEBa3RC62XmMUU7GyGiTUMB
HiDLWKVDHROf5w5KX9vJP7o1WenuvNQgdmJHtfZyjpuyZTThL2i1gkvBwrnMKuLQ
lLiZJS5UtzpnObCrZ4fRLMO6dmJb9YL23K7x93c/AR5rFJuFxgQ8ovKN5/cA4qZw
fUNY5MM8eTr1VXMGVPyrL+g3k06is7ma93ShpzwCD4VAbdE9QCntzNW2cOSKuJbr
t0Cdn6Wwsmz5ULvo0Nv8fFmv/f+CDTYkZeFO1FbFyGZHnTvRuSvfGThl+pdoPpys
Eq7l7v4bmRcGpGCVOXDnFLe8tv/ScVAQNV/SPHzNa+bSPe+6BeRG0ZPLVZYd1o1x
TCBiVzr7A/c+ywCPRQ3HKeWtBsx96+DNyutUPBWR3YuPR83f1ru7Xsus8fHlxEOf
qidQFDLmCv5pAVgKUsjAmFv+1pt+P93e/8rhYLD8AFCOK+NYZNHbJQYWvkBA9gq6
QX2wbbGQre7j1/VbV7Mu/JBnJeN4K3w4UUo7XFR4BF4XVu9mOWJkGQwLjyVTUSgd
IHqw4TW3b+PMhk7XzWWFnTIbRJPuGOTdbKf6oqt1dmCP92kLSzGO8Ng0eJJZIkK6
ewZ9CcgAdK3FeWaaKtUSwMMSH9G1ExgPBsF8+ilJ7k4Mo+jR40LGhGbJ/Se5iZXZ
0HD8/dv9pWqVjNoJjjjWAvWnq8Wq+QWZxVfxhoj6yst/UGA6mr19GdeUTLg77E2+
XfToWf6JMr2PXoaSkIHhmZ6e9etQ4o8n1pEm1yO4mX+cJRHZMSkal4Jy8Bf23LUE
cTszCGxvBvxwop7+ZHe5d53Lb4bw3urlen9kKbyQDLAN9Vh9IGP05789uJjcDSaC
NrkdeEN0R3l7VYknh0Q69Zc/0FlQlGTFkBZ0s9JkJAUqQidieBaGp4Ifc7vVq4BD
6rTVR3FpR8betanHa7AFwXL/0N7aQ2Z3JT44uJDsd6hS4h7L/ZavwM8qIdBlEinK
yWm7P0UtzxHJkijJjFURgXLlhdj3chKs69zs5srmspI2svYcYQN12K+4Ma4eGpoR
0e5C+slZZxND27Hc8imnxe5/L3G+MNyNF9QvMx9WcuJy1Sg0fxIE0QkLNi0idafY
aJ8XiYluunUj5gmHhHktrSeEh1Qj85hSp48GfKkdcmhmjeV1PScsgfRaUNaqCOf/
TzdmnPseIABaC5f9ybCWOo5Ha2646TvctRIR4b7iFaiC+cahRjUAu5eCTJM1h17T
ho217qPi07m0TAAnwzjOpfRWgs/hWyrgUDCaOAtDFD14zf7qI+MYEoZA8J9TwyP8
3XJSWSNY5hZVjPPOKueIDVHBq1ppBSPUDUeJ5xt4tXjTYummHGwT4NBZTTeVfidQ
TC1wxmVDPQq02i1jxeXyDwVmRIml1o6f/DreQ3WByZe+PRbQdGsPtbe86WXPcLEh
aU4LL8gpIHgca44H7WMOGvRCdrXIIbkNaBHfRO1naKzdNn/z8WJ7aPdcKT8na+r2
+oH002as79Uy7M+r5wlWtu1d9qGa94Qa9NIRQuO8+9n4ufWV895+oyrZyxpQaMf/
5nkUJ5NYv2ZEoHuT9CJIC9zgjnqA2aOtPq/0/aJ12j50JTHJoyw3XEJjJOb1/K4D
XaoYH6t817q47hoROYn3o66gt3d223kyyvaF72E5MdTuuyvOZe5ttz3qKaCzS54t
sKxZ/TiJ4VZt0RzAep3WFwU3nrxW2RlaPr7GDBYzeVtk1BZZmoSe+c69ei+GYsY7
H/UpwEerT5j/Nm6MyJSaDxCbzNSw9rWV4UZhWhYQloCpiQtVOMTGcQX5WyJKp+6U
lP4ee4YHEthTeoOz+MKiLNoWychTO6Xqjp54V7wPOUf+wU0uL9557DqbsYIU04lN
LEfKEdfLEF6eoGrSf4opooCnnPHrcIuFMj4wqh0kJAZJr7iYAkZn/Cs9nJRHCFR3
LibCuOccxrTH+b9dzTvPfOhuGmyj0W12aZ/GL3B+P2XeOk1h0ZBDloRhfx3kcdYb
kXmUFT8XV444vYGUMAVHyoVVPN3YTYFJXcn/xd+4uuUonXdXxibv3HAjY6RdUAse
iHYd+bGi/JrTsndDk/aDapygjN4vVZ7S2lisH5Mkywg54JXUXUrhPzf0c6WXZtOY
5vY8KkOGkPW1QistLm/5zgDSbHbm3FoQOgMJ20LTGK6SKFs0X71I5Iy/1Btk6ABt
iGVnc0avtPDJmK6DR+10jOyDQRBGCKboWgRkzr++tXmYFG2/ch5nwOV7VKJQN4eQ
zfS3VLaOhD+isrPLhZZRR7x3sdNApb2Cg9cp82oc/68u+BIFoYE0lkHMMtuZCfKL
mts7g2wA00wFH9wkJ5JZf9iK/8N8EjwXzuQzSG9ideCBF6yloC6uMb0bIFOHzyHH
YTHNBTPYEI2SXkmns1b7oXa+EnGhbgv+9rNUATIMhLaEvQ7TaCA7o1YQgMAg2j/Q
0HRrIulLiq7ExQfr3/KKsa31xZyUadM1VAf6+3pDa0lOm8A9c8cM09x/Z9X5rhVx
lUsX6A838U4HA/uFq1W5uI05S9TA6KMcvZq9yvJX55r4sA3s0KZzityUnmceQiyE
UuJNDl/SEk59P4veM10+O84MF80EXrKGEdpoH95QYAOYdVww939LCrFa3rBP4yTY
UXqOWqiQ4Cmq3TKLo0YXvq1+HWT1vup8MdGJUNx7DdkhIkZHFnDg9d3QlkDuxfMD
EG38F5JlXPusu67hGSf5gZKyK+B75OhuB+Ru3Kolfq50JG1ZpYn/0LytghQR/tgC
2ximlOEVOlvSI/xTKzbniz5xDOcgTfw82rmrQ8rh9rQWrCuM4+hTIj9Ec5aSWwJO
E3adkkRfHJLP8kKFSP+NwCz0+LhFwcnhItblVZxu2TokUc4ue1rRUCCIvXzc9tiK
g7e3gl1SldkvB/ZEPVMJ9rtQtnxMmqT3Rv50sMrYDogO7uC1yzyuij6hBWmsGn8r
eLPksX7Zj3148O1swYaScDkdl08neGzo/AcYosUl1UIOxc8zms9Dt758Oky/VJr7
YqHeGaK9SR54r5ueWdU8Fs7guuEPbnD2VCyaZK4iLXx6JuTOjWXJslq50NwAreXm
3wjRgezuaK6BFT7pJ774yuq7TGBbHcsstHV0bSoh+IphzL8Y5eVDZB6YYJeoCAfp
KWNskcHlaV9+Gb46wOfbn9uyw+xOGPhziI+Y5VZJyqXPael/vsrSDzPdbAwQnw4v
I4ROOX2ahg9cGvfFPeV5ykiYyIErHxap5xs3j0ngkDCrCCfGAqRR08W/1rPEo+/p
T3mz+a3c96GSHCu4QULN8r3cdmEWRDeI+H+h8y2EOe4/Aii2iwuFjyZEkuOGmXhV
WZLeX3y8ePs8QOmbE5n4qdR+7raO2ID+KvWcHsKbgRqes4WLsAkAw/ELct4pPqCp
gur3AUNACcETRComMRu5x/Vc9cbNphksMUeUR+s9LCvPwjMRtRruzzRZo+vj9fO7
ULIpODiXyUOjf8wAwc6jPJ21sxHtfsmZSnSEdKUvHT+kU7We70M+1dB9tdHvtClg
msH08YbMj0Cr7iCkbIDS/WfsMypQBjki2lMX4UYKHGC2lGIvopRWn8EOMuZu8KaJ
fNAwyCLKE81/rrk4Cn3ZqHfngkGjHHyY7G5Xy4A9ubME4ZorlYgDfvKmItekpmvf
z8Ue2k2rUU8/qIz17kM4Jt1LK76aFIGqQkBQlduU+LY2eWZLGoCnGiyId8W3+0+h
eKZ8zbvG0j2wwcpxETfUknh+OFP147BPjMia7SW1bkZ8MxnVvgP4Lb7ScvAHOU/n
gg7E6UFkJ4B8s3KJu29ZxuoKUrN5JLVb5OhYSQZFIwYrcfE+1gPodUbx6VHlpjlW
7ije9pij7iXpD2HsR8fyd9mKbGzqoyZBqRCGiJDbQ/fu4ZfHjUJ8cP5uRJzyi8PR
VstPQCY83FsReezNlqd3e8TuxnT5XpCoOC9qG+MNBtgrGk5uFpbb54wMetlujc6Q
pZ4Pv0X+PRUSRyZM3IeX1pzSzlon2j/qpmJ9D8pbmct8GUbhJ/I+GYTadAHjndk3
7IM4y8BczKkA49+y1XryVly8iS8EQAnfcXugVM0D8BNqYpbcpKKblwkoQmxTTbjy
66z95P0HiOph66mv9KIkRrNt9fpmfQGeRK2Laz8Ezs65gd+Wu7jxVJPxktqK7dyJ
zQvV0kYvc8tluylMI/SM1GzuySrgLqltmbLJaWEQ2cvCEGaGaVKrhyBVdzTEOiK3
hLBw+I9pn4F5R/3xZqLX54p+cQSUu5/dKAu3hFu1kqZP95RaGaDsdvwD396zVN2L
sXEelkLwCukjRdD4Tnac7rBudUvzpKBGWnLsD99y45CLcSc4DAie6ob3jqyQWgkk
tOiK1fshPnSaIvM22CGBdW7svsaMwMYFjwSpFgXKsuU14kRHcDj0MEo1HUR6EHqK
ptKvphIurXVF7IPGGvknoo7tVDetJdfMLSt35yliQGfVHK9OC4CfVwt0ue/QCC0M
Wvk4b5iuZHIanZfq6oo7ie6qS+ZMz0F7qu34Fa17YDnWU5062hiHSnXPHr55b1DZ
XxyiAZQm5U4NVx+uY6V6rf67Aw8O+ZxyaRUaUu4wUZ8YGVCHolXSri1mLZYg3Es5
aYlF4O1+YMgNlnKffji59a4M2fovMK9mS8kNtSO997RgAAx8tcs+BvsW9+3mtnbi
hWlvFCDLyRWe+Mlny7GMHdwAvgMuRf9mTvDSM1Jrx39Qv1PLpXmFead9Zm2xpqA6
+PqH2CLP2uVJg2my0b15hN+7KV1L102/WGLN4AKOUSMFBNtrez5T+/lTznPBHA0u
V4djqpaoIMypS0pRgtfCWUsRkoTd4ZHkogVBFS5tXju6zMfYxm+AB7eoq3BniiW/
cxq5MG2RJ+oB0qNPj8LMWpANbNljCl7x5SJZWeaIjwWYa3fc6CeYu0Y6ZCDK2aK2
qy4RXxlkiqy8TkaEdjj2CPYjF+ZMxsyOg3VPgutDfdcgowN2otYLciXftiRmsWT/
AWn2z7CpBar0//80yW2zmc2RBxN6zSuEdNuTMr4SLDfX+OjZx9YweUqLRQRjHw4K
lccEH2DDWeY0k4ewnx4CD2hiZK3/nL6c8AxtJiuFBgU1bNgnMcxCrAZrmzFLLpey
r6/SQEnQ4Z1q9sT8WiQchH2QFMbTznZ2IUznUQ27BV433mTbbOxLSdb34UwqNlLD
QqP4nC4YSHGsSFx9KnMwtRkTEnNFwMQMXj39eVxWd/Y3sSCdZKojS5SAxUf/WKEq
tH/8SgvUfh4PkIydtYxQg6lm4z1TF8CIi7cekOl1mKQVT4J0c4th1cGPxa7wB98k
O2mf+/N2qjNKSPqT5ZIheE82zJ0L1yyIUd8HII5QXoRCf8rT6DJI2/+laTO3kKjN
2NKJ3I0kmORmNaaySX0F+/PIQAXpg4OLS3oCCNnOcl3Y7b6OmXdeaMgwV07hHzSq
GswqQTBJhzd9C4w7+evLj9xAuhkG7IAinWMd1peeRTc1mH6Ik28WEXKxhtQzSqRY
iBziT9SQQ7iEYPywrGk787ZKrQLmINxU+xXyrjgJNka6tdoY3GM77dEWsv+Ww9wZ
mWfKrbxH6V+L/e54Jge3yrnZTC3rMGiAkum0kKggKfCYd3Z0/kmTsK7JkKkxuBhu
Idzfnv0ZECujq27RcJGL8Wz1m4tB0kWe3uNFjgJ61H7PldWz754iO9fwq5SguKL6
oFbevolG3UErm4XFDUl/iFvMU9PFubelWFiPiZNKvSwfaTUzNCZbfxkU3GrLm8ll
DfUT8q6hjdBhoBkG4DlCwv65fsY0Q5/muVf1eds2kEbz4Lldgn4dTyXXzI4sJzgc
dC3ZK51sfDxttX9yZJbx4CUwmFDXGgg6EZC/w92/ph+5KsiSzRDI2VLReks//9HL
k/wqlrRaJJfFyb0uHfyhTl/2a6h0VfjoLRWvoX4XJhTBr1aKJkdAu+O79lo6dutm
3vwWkTVwCE4IYNThpjjIzcs3h7dmXUjtaInyFymHIJl+D9R27vcn8p4PfrkR5UCH
NG2K7Lmk5a4Fm5Utworq+TjfhsFYtQI5ZwmwKlWEcrM2ghqfLXp1S/G6rnc0pkrO
7QBrmQ8jsk/68WNdQ1wR6k3HI3bkdT7PA132TLV4Bd0HPyvejM/khh/MXDphrecF
xhIPcS2lX8Uefou2Y8wrAZr6KS4bkZeuVJIULa8nHQPfCKdTFAtRk6wAtw/5Bo4N
7Dvj0vxhFPIBJ4iiQDETkQI6OkkHBT7Qy93PBqu0RUTo6kbxrS4y/jP6oJZWTNyQ
AbTyW0+MJv896QBQr0ToSTSzSuti3LHqEJT7c6JnIc0GtyaQKaVukxx5Vy+O0Ja0
ydugz1gNKOTjDjVAlBext+K2x5Gj7U3szeifkZZPyclpb2KhSHnhPN+Qrny3l319
QtgC70SW8I4dVFRUxeMQwdXCtpkC3gd+jAf/CBuWqowQstkH/UGDnxzvS0DgZ3wV
rQX3N5hs+I5emmzclo6OFDiQUK4lfu+IJkXUgZtLYqCxyDNM/RnYuYYmZwPJsAto
NLjDgOgyUM/JD7Ss2rz2/ZIxEZmutBmiqNtc9idIHB/s++2mQNzLQgVGOgWXHQ6i
zw8RQfemPvGXIioCuiQ1WyGlVEUH4ePx0IaFdSxEOaHvQ36VstqGNxa3ssyrK98D
oJeZ/jc65xobWU3y+JPz8gz8Lw0kGhkhMs+Je4G0vU6kzuay0lgtB4VwabWoi2r0
4rfOvrEbijgshN91+wjD93oj6d0zWzJzbRMFOzBDfzxDTc317LSgpkV2ne3ZIKB2
3Deh8HM1tgsgXCuJq8ESx2bOKf8Kpk7GAFQEGunD276HN7Opybv8a5Qt4hAq8frO
7KFXaNHIX7JM+4GPks3kLQb9+6NYaMt/UobjGCLTdAK9j2J8RyVlgNzYl4jY/0ln
R99deIauDZnyzkRhaG5VdSTc13f411XAOMmYFvlejEXYzjIfRBUAwsqvu2VebCF2
yYc/rDyTJM9Kp4cMSpyaofO1NftFKlU9tgqQdtTE+PDTbpXcJtD93xqAcM5f4iGg
6G7cdjCcdpE0tOqD9DR9SXFkMXHZ1EG4emh15C+pOsiXGzhMrfDHPUunsSlRlly4
khNGJp7lNQESlrCLH/dZgS8D/9rWye6tUb35j35KMf+vZrnEFYuj916UX11K/am6
FsaH2iCbka8ApkpnEFvBTRQPKc0TC4idR03Yk2Zm/EjSTbuYKN6KldHP6YkJMN20
2MJxrjqxKEgLbkUpZovs7dV9CN9ntjtEtNgd8U1NMonYANPKtcCkG3NuxEIv1rDd
F14Xx7vo+0oOVIqWdqkXjDYjuR1YhtzpuGJcVb/WC9ehoM9uTErdrwXGDbAxgBfz
hsWC8anbFlqF9jdGqB0nErCgAyWJDWyaiDEj3jjbyV3n+gRMAbDWE4RZfQb/HVd1
HzSrTieSLlKSu1VrQ1/UNxQZpEaAu99450w1b6dibNSM3bzczQaHkRwAcIfT2CxE
ZJPuS3x3ZzxGlBlLibxSs5TLGeouV5y6y6cjoBCpybo+1nOnw8Q1S2KJ5lWfvw3o
FA83nYVJB+5zzfGmlt2GNRmgkE+hzaQKeRuQ7tuMSWVI1m9mpCzdmy7SPw2Zg7LH
+dJrI+p6Au0cz2hnLSqXGEWbVXd7Z3kk5XAidBeYT5lOLdul3E+wdS+0oSdQdROz
FmE1NM7+5JenI8+vZahhycCYiX3+3wn7Hmd541Cep+8li2VLBaSETU6nxJrmolgI
63GqNd26xywgqqASEy3ann34/f+z52FeRNZ/jcBOXfmBrgnBXJJvR3I2Qgh3H7a0
8FNbFBVdeRupVOzRjEqy+VfjtGFfMlnbW39cAREhy4cMZ3Gv3TmDPQHv3wlIcFEA
5cnBrXkh/tnr/KLZCk5JmGN51Lq4cYMDwukww/lvLXtcfnNyV/DF2/Nj43VWbt4x
JoqD6yYvK/z9GMpWoRSlDXIzG5TBu+IgcJ9AV5sWG8RVg4xWCT0Poli3WjSnAyDh
WpWj+zhtM6rTqknCqgCxzFnl8Mv7TbLchTzePrie5IF6xYFfdA/IWulprnpiBVaE
P8GgjaAfXkyMMaLkOtULkNMkDYICwlXYYCMnwI3Q2we/w3NUlZgTXFXusuX6X5cR
qcoEWD3NFf1mjebu3Yboe9W7CEq8sism9lC7BlOQQu+C637P535NcBkYCYPtcBwW
Q3H3jpeOF52HX7DqWnYoVhP78FKVff+dVKfrLHZNKTKSQ1YB84Ay8Z7K/bknOxfv
hPMZBgdV/p+GZW4Xqfx00KBiFlzA+GhKAjJ8vBzLibCrvLeNGETzYxrvyoiwP97q
dviKlcxlkpmwnJT3r8ptAz8YQk4ztKYoSTDi17Ky5+wYq5uZwQW5au9aOJ5Vpk8/
OlxyiXGAN8e8YGbPWu9P2oasAut0cGko20KxQJ82tVDWqvjOAkLjhwZMdWFm82jp
wbUWM35tlEglpbTvdOqChhU7Dxa6bY0oB/BZrECZhJOyfQFKJwA+EmkY2DSMb2sY
SWPr28IkjuDvQWavJUm4WZHOv+TISNAub1SXcqFCQKCzz6pB7n92zzPmyzi+GYjm
VjSfy90Qunh4x5IYhVwoyoCWp5OmgZzVfpq3ixHzzFv4hXTX2JBgP0ILeoCxLmpx
udt8Cb3OHHBzZbPyngQXgmQ7pIB6WUG5bBiqDGHeTDGeFUGtPuH3bt56gbx5t9G+
Qs0xrOtpzITlhvqoFxvqnGa2JY9P+6DR86TcWADpp338O7lDJoTANJtr6mI1JQTW
mw7gdN34x3kx4M8ZnOzb1w1zk3w19xtehmTINfs4IEy82hQEwbH5+mq2lB+PaONK
StuLINkyLs3o8B4QUalikQbAOr1608I3BM1JsdC8YDtCEBEBlaiyP+ShlHPK93/G
m7UmsEK7dnPyEVmLXXF+whabgedV5XrxMWvKqlMhd+AH7579BvcmXbe+yvdIeves
xJsBQ7NDE/Ozgz2ISPf5ZObvSiobS3u3sPHfXT29KHUOsxzoyN1df1X/5zrCaoGN
5mO+TVmh6o+7DOT+9hhsBdjHgLdhlRImK0D3kmKaIG0kRs66m7zyzJX4bAKCTt13
pTJVMsGuFZIvi3PWZosmd+psRIhwJDtmwZm9apkVSuK1/1bj6ZyyB11YTsTNYAi1
bpRVXfEGuq5kDEcu6foD3nozBhnB8RmV3phw/Mbe7yNxaDqkmRNMDr3GnQmBGEAh
ymXUtUXMQDzfawO79PIy8cDu7/vnaGUi8qYyMAcAyl8d6xFrvkeRxPB/2Got7E7V
C2u9Qtoku6M1GDbT5BSi3o9B+zEoOwKxcVyi6PMsuaB5dYMIPevAsyXR44m8CUxE
jkVTqd5PIqmuyN/4+8988jKjRbZ9Hp9AMbNjcCagzm/JDgdHnYYMXdyn+DUIipDJ
9mnThcmn4yQ3wOYbgiSoNH/mWLPBAefMb/KVIPhETtPQV0ixebgwiMTgcw8HD3p5
9o4cMoAs/fJDvgO58cErUB6xl5L9rna72lU2icH9Xc3PfFkmcOdWSquHowVZ7miU
otsLuYtp8cQiydFHXwhuQ/+n7wwOxAoUg533YBYQWPW6CJSHcL6ht11FOyWhp4eR
EqRBDch4ehpspY0dLYyATmrSBA7zE2viabFzaWcdEknLLwY2/R8moi+u7W4xuRZ3
IwIwoF6fuKkp2NemjXXKdP97SUAGcUziXMd83kjFt2oCwdGHN1rmTxI3H2yjUsDA
C0Ag3wELkhjzEyHghDRZcPVziybqv6ECuixFjPN18M0s3F2yHy71uistIWZqhYJM
6rzprSo9mELtxqOKNVQrd49Oikut8VV+Jix86Z3wa3uGV/7P8yPIEDlnT+8mlGf0
GFoNk1l99qi9kTyyYvm5jDwNrbG93LZrThhngMnqNxyi8M6GwlU0tubkomGOa+ho
VTaGLf+ay2qwyg1lGjET1g1jfuaM287PSSiiQbMrlqmTnR4UXcs/HViEQ8AdNY5X
oX1I+UlbzzSha/G8DozVd2Nr01r56hQc1+sE3SvvtYUpzRDtjs1zoPz5wEYZojNM
LbSlN5NKBOdr1yPlPeghLUmMlSHV+yt4aq73u5dI9eotPvCyX/Jktq4jb5D01ijs
JtH7tphVz5Jeoh3YeuuVS9na4z/+gP8ACQH6Kh6YNbrPCxDZOE1TnAiefVwNcshb
TBoUMNI4L+r+7Ro1cC8+cZcD+I+a+890uNdSVuDBajKfGRmV+7z67VBFD+KlIvra
TWW0hHXcNa3Bp4Mil21dgrH4QUV+I3lNkZJZfnE2EIMIU8IXwqWz9ewXM+GrRjoW
Q3s10Yy6X7QVkGDYiayalaqUtjZ6R5GtFDvP9yMq1eL/rh/IURBauUuicmV7Ft39
i9ug/F5G1ih528nDNZVzhCp6fgh3a1A6mTv/W909WYWXbulDJaC+IAFk7rLD91DZ
M4doB2P/MhncKQ5Gk8VQgM7qR3y8Okhwwm3+XsjSVxsIunF5d1QBuvJTDGIEYiRh
ggp+C80zhPJRCH0RPTn7CFyWP5lJozs/WTw5L/1pTPMz5XoCrS9b+Lw3vX5mIu17
gjne0cSpF5b66wvzD+62FqHYt0dn4p+9rD1aGI8gl3yAR0tZdRG11bGmHn3RIM3Y
sdHqhDx2tNG7RkeGf3rTg2rfq9oL1W8WdOmVFqy1xCtvR9GaD8MxaWf+DxzZFDsL
+/hO6/a9Phroq2cqsTZiORNDCSz67rz6/+HJDqkt0uA+egXlK3uDZLtD4U/RZMG8
Ycj20HrywO9Vbiz5AH6Sw7QCoWNgtMa4J2u0HtNzdD3+i3ZtqkJsmMU7MMwcVOss
ZbnQE7BjY6yXYzlqOCVXH1vd9rYtHUAFe8jxYdMxuVMxf0CAtUpofM2FcyKsYoJ6
amtNi8CObUqbsDpnGvi6c3RyhP08s/0yOO/2/vcH18bRd53wYqok/MAuJlZe51EP
zaofIZvEEbkVbSQG3aW76FPDMsrNVTYTAb7lU63Ysnjpffu5MoKqt3rnudHsS9NK
eTNAmuiV1qTl57NfoDAXHKdldbUcfIugeCU6bV0okwWjjGfq9RyCUE4gEmIwB5F1
WXSbKdvhPigvzjf1bGzKxfayR87wePbJMAciox8nQgq6+xYQ6vstuLVtwE8cezUy
FaHZXea1ElzeGZS/QSq6sC5JyAiiS0nEQKsLAK2crnerKrAwNan/ewKG+508FPrC
T6BX79i7qF9VUItRmvhA0tbW8e1yPaZU2P7kZCruJmlVYTicydxC5N9Z7DMYdfqx
PeO0GZtQUSiUPO6EIlua7E3oBzxbZp14nvyUOMlcbDbmXrjgY3aEgM1VIGZ+gMxN
nLoeHl/1sPcQ2y8KRg4KmpJHwxj7cwvgWzeNaYyLuAW2wCLu1i2xbSJjvAtVkO4S
jszUeaMsbPe3hVffh9eN+pu852Rj0cqsXSHGqx8ZakjSjrkIyE4T48VQaWnx0p28
JOhcxv2aaUIpjRcLtViZ5EZz91NoBSUpjOMetlz2r+q7Vl+Tf1gA5WEwlDAezw1b
MU9YOUXiSGCybkIAAPlIhtddyhMt4cErjQfcHhzkuW0Tv3z93Qgihkmc1HY0LTTB
H6iElqNBxLvDxn5fD+UZyj02J9G1rm/KTq4U174Foet4zeajzVUn3d4HMQp7VLjH
xTK6SvyzPBpuRgj0GqjwCpjMKwx3lMQxzA4K7s/iPufS5lGOp1qds3zissIYwyav
HaNoVJyVxuzdY/4BbEvM247PgElp+dL84kbTR8V0LWiYuCEBHsSoRBnZSnlpIdNo
p5QD7JIy1Dl6RomFo48m72cCHsUcRSCHHQyIdItxpskySfAYKUXLq7YNysjo3MzA
3JzSitJS2dh9OU9rjty/sFfRGO3B43EaH5vn2KBsU65CEppKiJ6+0IDDgvN1aSrm
G6p3ggjHEq+dClJ5rXm1qO9K967LzuWugzHx6j4Q7235ZEnGo5bNRNhTJy7zNEhc
mKlLdmwbR6z0NTEjQXNPQdbDLBFmOJPxCtgsykaQJVvmtcWqWCfSwZkhbqolfAj1
LBxE6Ab+CGxrjRqmGrmBjEvPRpbzIn1G6hSvOT9yyE1tZ8rAkPG5EQqO0u6YDogC
kXb7vm6I4FQ9G/cDN7xRjeJCwBoVU6uxNV2iWh+jdUT/EbBIY+0+QPoiMZFR7x27
Vj3b42p2yV7Ye7g6MIE7rMRbAt4MFe6/SQo/8ytKTlJKbE2NT2wmccorJZ0J+9f3
ssdYC2KrlU7ZkiN5FNrzY6g4s7SaG8EdbdMS3xN2PDF0xeQTi9E2MoNgmbSLf1+W
FkC8p0kS4nwPty+a4F2N2sLcpzEQ8fNs9gmVW+rkSvpHoTrWi0Sk7OvFRI0o82FA
qbNcNlM08eU4XWHXJEuNlJ+/Dc82bHjjsKkY7n2dMWslvyFfUX7aWbw00mgaJTcF
muTchYU5+wcjM75Jmjz26UxHrO3sG595d4hznfAJrvkIVg9xdsvASEZZYuh8/hvP
QfKYvjeUDmcKD1EuEDt/xOY6p4oEXenh/MN9PLcFH//SvGbDIhfnGquoTcMAEk+3
++eVwVMhZjFbnlfesml2gehdhipEdNLwucXG1xZGAIyivHBesg4DaBQezJofysLZ
jN921uUEuKy3clXZ8i38zxYH+DgeRC/8zHWEqs1adi4tq7cf//OVDDbZ6caI/P0m
QAv+JkkjxAKet4DvKKhdZUUh6r5ijzQ7Lm+2B60+UA4gdQ80BcFFhLy0Th5x4Eg/
Vg4riGiLSIChhnjgvAmntWSZx7Hkl/SeATjpNARjsRuyVdfwz5r3d7spic5Zjs9g
bBNNK2k5WYOicdDIabAKz9CyfONzqI/4GNemUGcZ/3Krpk9eY8N2t/iHQKkCneKu
QAxueTLVw6vBJk2Xw1Lw3Jk2GkrBpzRlpvcdHcWcNyU7UoaDF1FZAcEXBs2us8K/
N1D7tLeRctFCk94PWHzJx/lLmH85UYxNTfF8oA0zJU8L/Uf1qVM2X0FSPX7lVraI
v38Yawm82jF6KkezJRk+3Z4oXvt/1BlSQc2zc8VZpNJ/N/Sxpo4y9Cm+9flgFNey
wKff3KPytihICckuNumZlnKC3w4S/wrQ/ypMYAF3aGqmrnzRDXmVviu+15876PKd
ZxP+DaZ7k9UOgs6ttA/ARp0JleyLYl7kvv70JiBvmPtwzXsPHBVDifa8nDAEQy+a
gcwGSTIFReKleSuN3aekQI/PaHMywvwCQduc55ez05rx4QqFBVSvzMx/qGCBAEZb
KfNhgtsxs1M/ONP+3oCfTrJP0D3lzF9swDFLKxtEu8hCYBeBsFOZZdHP8CaIOthB
ZtfnVCxCsXK6WlyMvCUYYrzebcaTS6JNO93DilR3Wq8ehNuWtbsDi84/7zGD/Crx
X5PmNoHkOP4RYAj3a+nJqtvy1y3T/eD3ayY/kbvlZZEkc8xSS16klDaYCUM9g1Ae
SxXnky9l4Tlcyz4TbJvVJnGkOc0bjew5iRMzfKS9WuBDLFKU+858ti3Maon4v6hA
4KE7lvQD77xetpfwNnFcRueiU+G+eh31w9R4IPl7k8db99jgbZAVeD7fgXkf8X5o
nH2bhbTCWzwsJs17B2XcZgnBp16YTuO/ZUHSDJWCVtCJ1kE7fuieCfqOBpi2HvQY
mRURBsn+fv9FiUizGvX168PDsunEkTYZEhs4wqPRCvvukx9Qn3AG/9GXINYl4qYX
ptykPC5dIR3qgwb8n1vz4xaJ2hcltIIOjxUeovJDFnOFmzaghBj7fpmHNDhmBql/
uB2eCrUdr2u4gXYdxqoDI/VxQJ5pEDZFK1lEwkoHLQpa/5LOGov2Y58vwFj6ypj9
sHaNnzIhPgpOFKjqOXOsUCFYxxf9onbOb+rFcdpu89lQRm+6p82AFpAywbc1tk81
cf0Qk235lnERR/JHX4Z+ZBXJ2q+lqJGNLgUPZ66aH0b/4Mj+Kr2X7przZKduqGVP
hf4U7mvmyaQq99Lq7JOajTMulXLcgj/PM2WsRRCSNJjAyMqNM4qMrO/xzYltLCUG
0Bwu/QqCVpiGWhQX8HbiPSMQPJGH3XeKe214w+aTfrByPOqqB4Hw4JvBjUsq8RpB
x0js0zdXTjN74cpZkkmM9UxArrlwTI91QsfNg0g/klMXEL7ZjvLIJTbmPPnWvw3j
AdU3FCgt1te/dXYzbSTG2iPh8cp16KRtt9opYNpvL9fGbOu8G48oC5D+MKGxVQ7B
/YbrpC7GSmjfsNQYFJNkr2PS6k8GISSyzGNI/YY+Kzy9HbbtOm8l/GZea2/aJB5J
uZ2gp+qrf81Zp4lbHP8YzxlKDIncRiVPElUP+BuWuGMlFqJ5Jruh0Uj/L0Gh3Be2
CvCWCrU2EgwWcJilJzfQvCqQ3g+5QrQ+5sjM0teZMmiufWuwScYB8Si26jHu1ZBZ
c5OITtdels0JTMe4j3n8n1bPbwIym0nYNQALfLtfNo14KiOtrKQXlliSMSG94Uw2
iD+J4GR7/ULmnybeWexKzHl+2AxyruPgSoX6kHVE6PlK3cSGBLAofu8Wcx2D4Xdo
nD4L04SMRNBYd84ZogGvBJoil9ozDMsXrNqDsTuV6AIcewt8mzuSO4UGZiepRkCZ
CETLuvNrqfaiJXMy7w5Uc6ZTz05i1W57UGBwrb/tIxNJR3/7kHXpaZqJ5BXOjuN5
Vhp+eROhrAxSLYQ13uUwx4ZFnpcp9yAYu1nSSwMdXFvnjtIsI0wNJmS33qG+DgxG
3zyscwASugdc0lSmlyq0Py0QdzrnG9p8I6ETrb71acTg2e8eQh3IuOQYrCGGpJ7Z
MnDaH2aznDbHKZ38S4wV2aXb5MyvRssp5XHzen7aSxC5IcRNzkBYQWNXvRKycEgD
O7w2FfBloDQEue8aiO8SPI4usI8do6oRNFugi0hBK4ThfyTvMNImwSZ7471CF5Cx
6SrHlCoi/ZEioa/1QB3cr1b9lRqab4NZiwT6XOBxsKYvhvZCpfO8y9bLhruJax4J
aD6O+nCkcuEmipb4i3tJZGylHGaGqu2YFnGkSrE6MVeWLueByZgDbTpBAQe9bQPS
7vhjM9BW4riUIieqDDH0rbX/FXC99EVEE+rfTzr9Q9/2pE3U+RnTdgmyOp6hB1lS
wPkXDJZhEFI1tiah4DUaEufoIX1JgLRbKQRo8fOe/Zhaf5dUQjeZHL/3vVmEB7l4
snrCxwjpTOFdm1nypdklOFDHFCbojclyI2dMod9k+nae+biEflGrbKCzyLt162GN
k0lEsI1sCdUjA81elKS7wLgYDlGHmseAw3OnZlp0KN2czmDxOJuj+Jxov+Mkv128
Ptp1V/TJcKfkqympZ+fA+ThkpKX3IxIgMP1eheDqFWK6PG9Bro4yumaIQdvmZ04d
+1aMnOj1Xhr4nj+7C9aeg2uigCPwvcIuEKpUf5Vu0Qar1DXtofXWsSPpVTDJIuY2
/3CN4HdRFXV4/ats1HQhwKs3c4o054QeHwZ5A7NbH1WhyKG4gzRPTPzOfXXDMuQS
pyhi4xbBd/xTCYNZQvPlKPHF/UMX879UyKpCZlZK3JsHkgurPecG7dETF98qlcBC
DuEbhkvtZfznzREh6rAgIcwIPqvHaz4pZIMANIlxXe+3LskQOOId6C51s6h/fnjL
uixBCbWJP12KA0JH9bbp7otmD6LmhZuwOUzY9Zr5TcFjzzs+f4H52rFV9VSDT6ix
cEQl31lc1Ib2fY0Jo7Ti/Iils4ZGaAPTCd/WaJ6evFaJYGgwZfoGoHAKOYpB+nPd
Qqzfb6Vcbi7qeIcKCIGYWPT+y9efg2apKEd0KbG8s1fSMgq3jGaSW/NgX1rKwB4K
76px/6+FHMVJP7V+HVFmrC8W9LaRn5GdimqiKLHl+N+3+oltTRsGJKcKbpvgL3QF
FYqyFr2kTWdGC6Ij8BZ1H0VOKUfriCo7b6tdq2Q1RiWFmvKOLLVQ9N40j+relolp
W4GgOVUZe8AFZU4DCX8SANcUWhDi67087dqb55p0SrJMHs2h5nHNWSUn2vrnDUsI
DPY1LGH6LcHo6wLfebsNMpo/yY8AUL9H87W5SOlty1nO/cfLkxtkmLd1GGYeQVRr
PPt1SsV80Z+IoS2r81oJVjcoFIf22B6sdKtE4wAaEhcQGY5KPde1yEZEg4C+Vf1c
snM430pHI1GWb9oFA7cJ6BVfSpRTevxg2d7VviNZO4ESeetHxFRpYL+vbe3Giuhk
HzF+DHx7e2iI19BDUuk5MFr1yAKv5iiIxkKfhfyufyGpmGU8lJTH4XKK0v11ZFl6
J9b27R/GqTb4Mo55GitkY0JGfTkkNxktqtT+advhTz42og+hAaahmVGyVUeh+Iw7
2ZekAfm2hzoeDHh50rL4HEveVitGZZK681sqGfALxAzAboXQZjiMIgYw54qhaTrs
OYi1I3aZIeo5YC5BoxSSknQZtsyAQFiCddrShcawahbsdcmG8tYSQWBH0fGdW2qc
OgiSzFNXLN1p1xeyocPVCh0ufoA85+VxnF80qInY0JsDw0Krovz+8DCyioTSusMq
kuzWpgt0vEDBLKeYYKKVxKhWx6mnl1eOENs0Zt+Aa936972Z2VtAiq14t3z1KJK4
kQBDcspm7nqPHucbfukA/KLOf2z9WtMj77PwPPe/aVjx2HyyledFI9zzj/89FzL/
dEgoxQChsVPBUmq+qau80yADPNY+CWv0XQDkHUloqOcDgYjCgm1dwPlDvf7UMf47
uS48/vXHUSyZe2DuBuAk14rsXETDbZk11FHSOJ3+lsSGRVRhR+YdSeP5q165/cJ+
V/oFhs/RdWyTN5OJJFYaT6TkMpPG6s/YUlmdk2LaORFn0PKis8mAPeDxLwI60gzR
Flk8yckNWkjz2EONOd7/m1Q6OZ53zCftrTFa1+byYHA9DeaA9sVhVVKih77FwSza
/YXDmDppCrCi44nSwX9xrJg22F/4iZtmW3vJJ01TTLckrstSoDTPwcjSU13QPxvL
L0wMq1rkU4x5SSSilyLuTPz7JMxKfzbjTJmGT/Ok6v6bYISnctQRB0iEtyUmYskB
PyzgB6WyyVzFIAm+PSKHUMK9OxsvGXbJ3qtgnkkM0J0LMZ37puRZynadBIrcwfve
qj+R0sAwEoQY4H76CDnycHMN8iJE2A4crri9/4SaIN2s3XJD294nscuthsbb3iVm
rois2iZ93mQL9y/MSWodJaU9cnM4DmA6+Hp5P3XfNN0npmU5UcjPiOaM9m2msEXi
Gz9KgwEQ/dz/admeuF5tmPlQUfXOQmB+hKMG25FZAKPKF1eyNJdIe+NYA1lRNPp5
LgWb8uMxZ+tXbE0lQYvhIjn/staOCMi5HhnUfq8JY+AwSJWm/5hY/fiy+inxvKi+
sB9tJkVcjrL1p923OQd8oUQQoKdOyM20LCdF9pPvuFTAqoWW/Ic3KEHDTxXTtjUc
hyNwzFh775QVflnToGPzmAXdBGxPidGKa0UMQsq5ijNplFZFD3Ugz8c6yljik85y
SYYfkS6/S7evhqXf3kt4OortXOH+50QxEOosAAhr+j7SLkdEtP+XFi/AsrI7spGo
2PWb595bSrzgxHmPa7OODbVhBTimBAmygILkGn3Vh1xJPyXpVdP7QGO9g9NwcU2M
Xy21RO/vZBtmnxzbOLfjDp22uKzmiHbh7uFSNyXmV83xSj020BuO7TfrPW15KQoX
d9E0/v97u9CsvMH5JOBnRdd9SDgW3o24Mi/HP1M4ECVvlvHZ0X0+jfkZe91vurv+
Tsvtsu/WmJxf21RKkDF9lWU7hvNuY8Uvsw65xhdMimD3CFyZXOEmfQOklbwKzQ83
llioRs1tpn6d9z5rmYywfzG49rb4trNpiaO0GwDKkb7lpfuU5PujtjYDVvxQt8OR
TAeOEQZP+cTPkbtQAKVp0bp4HaLxjo21OIanEWDY/eEeywrZf5/L8uToGeXOlXGq
D1EUFlMS+4h0cNHMtCWBoTJqs6l0Gfr1ikpwswvlIUWJfJPGgdtlBWr8VoJJtFn3
LV3PfJeEX06RYZxpUA4MjEBqgwYPUvXGsobNBcdojy8JQMKYJVwdVj8RB5mIhnlz
STlwRFKXLzN/vN+gpRdUmLIEz9t12lVIHPYANKdCMW3aV4ehUhffJ1hYVrR9esTt
APbuwE9mOvM1Kd2fHPAT+v5Pbg/46ojzKuIFdF8qEq+zzr2ymNsyxAxus35H+MKN
sQJxAiuw5peCILvzhl7iwJWP10+YGSUflb7yG/hgY9TXnT1OmPNhiQwmPOB/IPqm
GXEd7+CT0hbnLw6oNjs4gIf8OamZu0zs6y0QIGgVGme3B7FauPDzA3Ejc8pH4X3V
L5xg7w54RivB/lsScMhgf4PEKRUMjDK+0RrkwGGBxezPCE2D7UOnYYpIhKSWcrEd
Re82uue18ei9F/jyndvVgL6u87r6Y2EuSrGcyiq3ccvpYA3ZBJIp6BWimKwjH8ML
2eYVo2Rz3aclg9RLrDwJhM7wLo5DGPFsJupsjogamYic7zrQIGX7LRmZtB0LPX+O
TIQgL8ymGeX/FGZuJTHx+0s5b4UdzsXtffqLGDxF/RR10lQh1rNa83oat0H23o1p
IRY2hH1Wp+Z9xkfBgKsmixmjKzMSODcBhnmexksHCW2/un8PJHM5VUgnCf+fgY+u
o4gfYTPgq08VH6c1LwIHE8hWo6QGVdI0h2IrB/qruzZlt2BgRQBtnTDfCVBTKK8d
ADRvaygUBuGtU7FbI5ES5mv52slu0UMUyWg2d14PBbdFn+mzEB4ug7Mwra5zm3WK
AwWaYYlm9zHay9t/ciBsbMa1zfkSy9glMgPc7DwIy8NTyiqu630qmHChpXQZvNL+
NEvZIq0cev/swdcPrQ/VjbXYOvyF3aIMb9Bp/TLl9U181duV3/xJkHIWp/5BjCyZ
b7dd3EyooC6ZMsUiVh2o93YBnHLlfMUSCD0z59WuuLgSPrsIXyu2n565dTMn7+Cr
y1CMui77+CFHbyo+9HwJko++9mMCNnMIROiQ1OxLOJxrJan5yG/EA2c7Eb1sGsOi
6OEXoQK4uCdy8qmzc7e+YQ8c7snjCMl5+zRrQyfBswQBV++LZ0MoTxgTdAH8uLA7
qyeBGHy3+tGWXIh1RpykHSd0MzcVv/k1kIlMmFlViCv62iRx03WxNyAzwCUMOlss
7//fh0lKN44HCAi9l22PReffXWUpuSYZHeGJ3R/Jdn/lhJmha8R5hKeLn8rt736n
9Vv/N0QdMyXh8rlnIEU6XVNW4OoJipKPZu/AQs5xbOFFiYWVNqBIWu2s8C0uLyqm
uhyOhDgv/hSPYGx6w2VirKIoYFk9SoeoHxhO4Y/N6G2DnxUUTBJwwBBC7jIlEyEb
/jRPLOGSKKMZJkttLYHT/iK3z4vEbqda5bbZQ9e85gR18Oq5RKQmAKlXKABI0P6o
l/7JXYfR9Dk5lCafvXPixX8f0k8qgm9JCKVxKgn7YCszjKzQqvMMuyYpwDO/pfnk
9UwyT/5rIYiwSoymdnPWRvqV9pUfRrlyjTi6Lw3nYLxnM8MwEOqA8EfnA2X7S3/p
+/YXCsw+QHtBiUEzjKrhOjdaGx3RvQkzsoe+OLoD02BRjWO1pq6c/oF4KUZyblTP
o63tdq5okCTtL8P3ZlZiCmcxivUBKgA2MhHJ2EZRLuHNvrirw8M8NUmeX7lW/KCJ
fxLjTD0ZPcPWTj628YGVBsK8ah181BqgGOKYbg30CSX4++k+D0UvAJBY2zn6Hx87
JQDgW4o1XhhsXUYRXEx/JmTDFmuBaq4+ozaOK7WSdP70/EmoUhcvQkM08Oi3gX4q
DksQttsRR97b7KghdZDfBBBEYtoprsfjyx2E2KxdyXKXvqq89YZQ07EvqE09riAx
+/p5iKM7cr38PF3PZ7DZTj65nirnIR68jDLuZoBjQmxyiusBZ6kWD7DVG+HeKIHj
SgarHphubP880eIa5UjMzbELfwkMoUP3ZrD07iH7vGWe1ilMyODdqdq/h514J7mC
EHnqGSc37vrDKidXr/bxicUePkDmews/ZSsIk+rI3kC35JOF1+FQiqhQjw+dO/kJ
VspfKqfd3LoiL37OQESSgdCHqMHq1l9mjIBBOWOsASrdz/j+dHSEhL5cmmDttoaN
pvT39hx47fy1ftZbLkZVQbTOgdkxq16E6xlUPvgpP3FiVMGfimXx6YOwCu0m1tPw
88s8gJVKa8qZGFs9ArBJTKKwEYICGLX16xzj1rXGVlLsASyvi554LHFFsC23DAeF
p6CDKN83tX19UUpPtr72a9BjHRb5V40KeZcroLy64kB8KZYdxF7A78MK46V13oAU
9/jaIjd9NScS0LXo54omLy/IdjcuCsN2D3jMZVsau43CZ8i+e0Q6KAQriZgfT8bo
WD10iEpBM4qPMuzpXXE5bs6FRSrfINuCInF/Cc5RrM10MRzHHOoLlpeclSXokYXb
6vSrSNtEH3Liqw4zzI3GZxwle86S1CYdzMpp/MZ+OqeCzfL+36aNGUWe7AddGwIa
y4u3o6bZt3aOU1EYo7ttztsrTFyGHgnJQQkr3kJPRVeNd8q3W/uTSTLbMYRKF+JQ
Ic2YJKZXwfn0Iw6U8+DNty2yiZku4TbPqJYX0nln3t1/eJ1fy0YVUy3M3Q5DyQil
m5RsDbWROU7h4ZFd1vUF4CN766rLIWUz5kMFJl3cWbN/w5vobnYKBComWuu0KiWH
I7G3wNOzBZAm3bfz+PlCr7Y5Bhk7Wlox7D5DF2WWamD4pGcwE/jjkTu4JtYkJ15N
zww3xUEXbIuj844pFam0Q9zjoHRBNAYPgGRqvYeQRIf/6wLKNo4LkMT2/QEmBHxs
VcpfFUXi7tHsdEqySZrxr7i7utV61JOAEDZDYRXsNwiPBA4GkdvPTXDb8hrv1U8z
y46x1IoBRiaYqaBLpS2HdpGhaez5danD5eE2Bq/112sU1GhBpLqvXBe8GYyTelSc
Q6tskEoIwesKcf+pYpiYuhSoXQ098VtXY+HkyQylrv9R9SjT5hJFSG6dCi/3UenR
ig8MhnUxeZwTlGMK5JNyWdqSVPL9vcqhemA+JOA2E2pNcuKICGaG6C5WN15qldcW
ObeWv6YcFWEeDf5hFeQDPR9N41ZYDbvOyQ6/MDDTbc6hmENSpPBvDWWmeRM4lxSt
lPRVwZeIpeE7FM6XV0xfHX+O2HpHDRibk4VibhrAEPO80jC5aibr8cafWvtYtvPR
hIq1LrdNl+UAkxAXYOilHIoP/12hjvUYc78JXvm43BLiPrvOFWuOcFH3vNVaupKj
Zdw60NI+wMM6xlALAj8djtbArhappMJCPdUbZFWp6EL+eSiEFwUKdt6wobluVCq7
sPBW9Mm3UY8zQfgOUH2LfHRUurSMxqErwbvttt8nPXEDnSyXKV//r3fYmdAvTctW
zGMGTUBnblI9/ODHU8jQc7Tm6LjtYuG8XSxZfiqUaOTlIhjjgvBvOqI/FS8fL4Mw
gXLKb5EmVGJP3BFD6a2rEAvfiL+0lFKksk/I0KFx3kGulg8Lqyec0svaCtxTQUTK
Opa0qcETwGi92PCC2pe+5VDl14AWcWWfGDMPNaoHPHO8fiSUhU/Z9axUdFSNYMBF
IfnEe9eDwoZy8MGg31sqVgk3ryCPNOZxuNa9VPvtybgX2goQ7j0IYb0pouxyrgCE
vz6e3Fw191XMgPxdjanzW0NuOwEr8Zdx7uGun+xbn7VrCCt3SZze3w/y81KIq5uc
PQ9Pe+yfAisJCtv7T4oMLz+0TqoUDMQuRQNglBhiqy39B/RYo0I2kiUdRz3KsDOH
kDlv2eHlNBbZSHEQg1nf+RP3f0D58xHgmCVJFqPpUYW8FCulICTA9AqBdLRY+2TI
G4+uH4T/xM/z7BJQKETFpXfePpul8ZNIQ/Ojmj94uY9P0papG7zExO021tQxrC70
walNywKjkpbA0nfaCSBK9HbKsnNTQfnFxkI87Xm1Yvux+8PQ5R/OR/hf9e0Ex8UQ
EQdbOMuRc1HkZ4wP+4UNT0vCvOg/XuPbX+fbjEKo42WI+I9xXkc15efMYVijJZYY
BXDs0PlUxDFvZ0le5TEIllq5opjtm0X+UIf3ZeBBDYJMRt6dEssxYd6koyv1k6qU
Hq51WiGuADz4Y7Y1r3Pz4YQDIivD2+fzBCnmhehTEASVawL1+Orl0+YhuS1IvsII
U4bcfB3X3bhEOgKoZt27ea2S+cP0R1IP74fTuag9esOXXClBAqZg3xP6hLXkk6v7
G82tdoTJLIvcBh0sDXi5C2C0dCIMPblP/dH3NjhTs28QqHrED2ztbnKVTKlQl52F
HCjM+zi1rmYtPs7f3nCDmPUOV3BvVI9MnefdD4wVvS330xsrKoR3pDDQP2p4bNMi
3tidNSpUp+1KcC5wEExJizt1C/+zSTvhWbWGUkT3eYOuebNA44CeNwcUoygwz37G
8QBh4y7SafU8a9EEIuSAYetuV3bqJ3gD3kYQRvfyLbAux9a+EX8q8xton2mBRBeG
maRqEW9jr+QA/HIjLuPaAyFBiE8rxUpCvr141TNd1kWIp6mnD7BjdMtoDqMHJrWM
NjUe5mBa9dK5daamb1Z//T44WnJZlJQ3RFGfQ6+Wp1u7MXrLgvdkN+hEc0KOAbjT
ErbN4bzMNjJBPGnZwOoJ1zuLaC17xaWQcUR4f197hD9oqJnfAvNkFL4XaVg+4mn5
FD96voNycBR4kjoH3HXPmOuQ/uu1CsAkSTb6iHWasq+MItKM/e9br7gJgJmYCxje
caCmsmZ7tKy8wa9OZKVm5jAs//wjWg6HsjxkhDBeTOIvHoONPqoKorj1Ok8l2XjZ
CHEO/ESHUiZkQmIU3Vmo7qKt8m9wS56oAROa8TAvIQ5pXdtuqadQxjCz3Q2cLV1p
5qnTmCfmOWt08sd50CMT8fttH1UWeF7km2jdba7F7JND7mXxuPuwlDUIQgYN7Tit
z9IPenuUh+VdcY8Jrhtt0BbY6sZk6KFnQNy29NdAGFRjSq4ZWIu6DrVbSsri7f4H
0T0wHHC+QcdRqijh+YsGQCHgms/NKjkJzaFFnLqJFzJCZ7j2aYdDd2tfTfG0il3/
/6r5iXzAesXHnqASlr+r68SLhcK2opOWhNGdV/oZfGdBA77TSaQuAN0mQNgMen9M
nNtjbq4stfqZv2Pi/CuNsK7ugkr/NOvooj3WzIlns97dy2QZjxTL4XNJiQrvgBXI
OWUUOMYWHhwtahwHWMv26SpMqfBWd2EFPbvPOkYdBdfvKok6zjHRmVZJ/B7g9iC9
z4Dp5oGvbAzuMRvF4ZsdtwpawPXnlVtUIyjxongtIDhY3lC4LGjmwFaBBsq+PSyW
O9S2cPqK7y4JOXZAnfNOaKklcEpRMxvB++O8Ebw8RFx7Eq5OE3AO81kHLLJl5TNu
hajQEHfTF3ptdam4W0LEPwrK04/7QH6Z4dERrkDeFjdQehYupBtblfPGyJLQ3YnR
kAONfqWetmfsqU/Qn5WW85CqrznakGaHS5wrgY43puE0D+7dRsTzGpd6K5b5L28H
4xP5r062LXS4yRj81X66mwHhef3KatDcqX+AwKC82Tw7YJBXLWawN+f/JD6bTT3g
DO9JPaMAedmh0JXv6FCD1pz/26gSDtMoNX4FAR1GBcXmkUx12ASwsX7VKEFKa70Y
zbWdnuwmXo0tvb7GIitt2k0jaCHVEHEPsvDj8ZgHqhOmEFwUUuc5bteVlVoHeyt5
YwKl4JykLv43mI5wk9UEdLFkcuXlW281WRnTW2wVWdYU7RARsZzydxAxnQaN8NTV
tK9tUv9gHtYG8y/pHV1kt6JMXQYIr/Rl+bJBZsfNgB1MCPDDzkPZjb87vbp312ZI
HkfZ4Y3HsiMsTwZzQ9Sa24SyGaqWbQMZD4v3ODQEkC3RDCpa8hfJCKgNYMM80jxT
rqCNYO/aYrEjpgfzUP3X1TZVWQ+c9vftTBfukB2iGsy9YW7/RVpR2PvgEn24CLXE
8MFE38EsZGz9G3HpkTjSD9ghbKzuHSwqPGabTEeQ4kriLz36GIFFKGmdLliu6Yq5
n2YPjbfA3oDrctAPogNV8g2Mu1a510gVPsdCzfWaANPKgBhZzcJSnNnmk9KBjtAu
NbZlVMvvQrfJmcOfyVcQxFgfi2eN0bPNd/H+65TDEIFpG2VopExksPB7q76bvtIN
qp/Q1zyO1ZvAGrPbDJLZlq6XxrhZzzFhgTMthXJlCnsX2sw382BO6VZXEg3OnO1F
/gVI1ctaeSJz3YYSA57TU568Bb51klyVn4eOtQ6injcqQM83P407/CsBaL7AZNHF
lav2jEuWxcFBarNFNW179OlFGmrwiiXTgzB70ning5OvJrkpcdT+Mh17GCV1qeOK
BiTAuAoQWJkWFT8jrnf0N43ZJfIGyMI5n2fYVaiPzlabepdm/o4Z9zaf2B/itJIG
0vrFTDdiRigglbrJMeOsW6Doo2Me9SpgNrFFOhvo/AkV5KNXKlSerDjV16BuURwe
ky2m7hS8Hn+C4PPqrHtxKAqihM0qg2VjpaptTQELzb3lLh6RiO7KGjbZwVNFeqgX
HFgZysiOF2fU0KHlyUBpedkdqUZcMJuOh4RpHftmBoxHc3zrSzfKScZtXbtH9ZFC
Z4Lx8HQDX0PWb43Qy5t2FqUc3sAQVfaUKILe11+eoxcsptLuDDlRw/cFZ0fDZtI+
xXzuGaxAT+IqGTy0cLuzlFTvbhqMn7g0qv6CnW2k9km7LPKR0dyKjC8EXz2roLrx
Ebjo5SQN6lB50vj6FJj9XQEwg/E94ngOCMTnUrBcKdt/F9+1XCDB42HVS7RjtsaM
wMbpVtVqwB0rk3e/JYdN4ZujQgXD9gwclYoD/drVH+CR4AvUMxc1XRjQlj0Ltk4d
ymbwgqHTNGglYG7EixKZgPAdz9LIZDRqFoRSffK0WWaHGgyfi3e+kSwSxyY1NKom
Lgz6jh4O3V8KCtXyuCoVXUL/57EHl01pnH+sRyqtzAyPOOU1JMfoJhHpxRUO7Dve
Vrh/s5gJaOtnX5qsjLoLrjbvG96/q4JCsH3uw672isKNIriU5XilvTxtd/051kJS
3KGFjBl6/TOBHF/EP19iDGS1taH2+W6m3RaWxhj85rutI/xsvz7j6zFe1iTnkOkW
J3YZJyAonmk3lo53imKkW+wS+F1+HAdEXFTVkoqBQJmlraz+w5k8kQe5y1BkQgdy
4H38+7r57aBsAurGogvz49kB2FPE5aZ2uaB64pUIKgNTNqL5WJYtyCFcuTaw8vGL
dB0QLGGX3EQtVB+kZ+YUih7RXh4+0OoM8ip/5287xA6AnKyDeOgaJAlVMNBtP8GP
uGWq/aBNlTqjbatMRD51t96ljCGgzMOUjQiuVOltojN1PKTWKRz0vwzFnaLiZLL7
YBjAvHB7Tek7/7EHdbsCQANB14nlYn3whoKO2T6p5cYSBhihwwzOIXX6vjd1ejCR
QwF1/TK7JvGHzvnqO4A6ASk5BO7E7LCWFKp+Tu9W06oYmu3PVZFNwDHrT6O1DSVM
kIMIPf2iqbeW9NHnrUjMXWwXvXcuDsLq1nHyYv3aT2HuF942i1co0uDQu7d3c8Y5
UybCQHsX6q8+AUYKKMZZtYGZX/9wrRgx4P1IDilNqrWOXydASOxYn8YzXFj9pHNA
iOIZ4DHTptAGx4bQNktmiQDcMeYkCenFzc19cL0K2auI2ip7fUqZTTPjuRjktdfX
DgbqzyENEr4VqLosNlfel3R9y4Sgs8MDmTIl6bafYfcTsWiPe6IIGdeHzriE6jYR
ilNH0VxSEb89MOd+AMoHh6wUwmYVoXuV1R3mOTxp53hQ+lNyEdd+gElv56PamakI
naja80H+x0OmnxF43ZnSChujvvY5NDPnTZ7fg3U1vs58zOPMQpkSDKMYMH6fUOLH
HOUJghlqB4zbyI4P+r+nDFsz1FV4hklzO4Ku2OFVMGNc8oj0lvIjgrfVKVV2tkCW
0w8+O+CUYNsM6gI84uLVW7hXXqWpLJ183j8eT+n/wlFTYlfKi1l5dWeDLOK8X8gF
Mm9sf5VSnFPG+WEKCkaksPbCk95A1oOF7DN2+dCZhLN4hWSnu0xneNnjscj/9mAB
1lytmzAqDIdD40uiTaNYlF6xwWTyWImI6g2NJXW/XFW9BUvvAbenrWIw5GJo67gq
WHb1MFVCW7iew6KapFiA3ev7SdydJUGTLY6UImUrT+K2rtVe3kb4OYJRZJsLWz9M
wRXsV6T0zTVfUlmfcLkJgVlrl6D3RQwL/cxhBuoB1+q8TKXyfuEpDlFJ7ftACvkr
Wej6dVDZIZqqL6Iea0ux+opC83TcxnrUWZW9G9MBioOOR6inaWRGknXlEx75UZzF
q0qbNsy1YGVHlgpD4O/3aVnZr/MBVEVsoz4XCYniP7YiXVTU3l7KG4us822BDeIv
aXcKhlGUzQfUPlx/YHKNEdzpcWU+klEZyHa3sizYZ8KGFPRigRq8seVhp5dOZ0nl
9zq7QTc7uTxyzSe0FJoDdTb+qaU5RbXyT4g3l1VVJrltehuG+RwSi93qmCAwqrWb
ZThx7UIxf8arYqfyumrDL4WX3jFxkBT7zj8yrwuGz7ZDUHA9pTGTPsrtLGYAhUUf
eGJXmU5wDlMmW2YZsQxirUHjtWrMKkqIL2jwhCLbpichiQ3tdIF+BwnlDc84dZrj
QlByRg+e6Dlf0VFXebsiP8DbPwgM5begEYk+ITkN9WyFroslTN/uOxe7DAYG42Zh
8KUkM972njKQDc3LxE/5nrQSkorV4XisPJQZg4R83tapfKrgdaRmw9T+FlnYAYAv
89bCp2L3necpRbE3hAYOTCwCiyi1TqBqNo3yvB2ewLcuBGy6IZxFWbSW5PxWfs0w
7tZUhIkSvK1L4FyB+7yLCR5YhqpzVXxlzDVmWLG0fR/2w3pdef5iQszZwo9D1Nlz
0cRGy9o7qYh5ZZbT/BWAYeB8amlS+UdYPv9cL1JtJ5nuOqQ7IrWMuBKE/cPzk8D+
lh4lYOQSzkv2zD6HS8w4+Gs7dwwGWgj5+ksFNz5gFbpjoU+2QPsXQ2geyoZ/Wa7p
kmwMf16Jpm6eWxTCOQzOGqgmbmzMmwxCwt2MsUmJXKE0rB5rtyTglh9rvCyBsSAB
/d+3MDjQzzHk0iEEvvweTKQEQyeXNCQnS+6GdqcFLCSife/bUc6u+T3SEX0Ezwob
PLs4ErBWFWlujtPNbkUWyEs6CKRzWulSMJwEVhXF+8+WkADWg5LhYIFnrWiOmZty
A7k/qExauEh6Vv7CeiZdsSEVChcjv9jyTfrT1pF82NcWBEu2vEOVP/yyAWCXoy5m
pW5PcqJz43dVjZZcIz1cD+pK7Q0zIE5aqHew4oWtnZuOIIq06XDD3k1redmo3Ouu
Qgp8VlLnuW02zLqookqm5po3rNqh/EHY4toEPfCiGi3JtpW57BLD11OaJTXzaZiH
5JEMzWUstzsWFtFkw45fFAsagEp1AFcYnqBUKhHc2ftz92R1qWb7NvK/BjDBUQs3
ENRfId+M32ndSxeEAFR/ER2O9pAQNYoiyLd/Ft6Ul2tMixuP9GfQQkIjNncYoNaW
pn84tM+VA8Y01SdqCc6pM8K85hWNyRaUG2W+6HkUnQp2R05JgO4mNciBQo2TEZ4w
TUFsXZtKzU93hlZVvpm+oQT2lwPRRog/D2Igp5S1YlGJ72LTV20teyPqi7vDCw4d
jnjDWX5ToKC6aqNbI1dtGXDVXlAM10irPwBnk/hxntLfi6k3zW3FHVHsaXS/2OeW
2D9+K5UGu1KFNAcIgNyfiaD6H1pRXbguiVPnPFWMimj1TPGwb46Sexjmk+LI2x9l
bT+q5regaTZfB01RNr/RqUQGFBEoC9gTPYFoMfrncgfvAEUmU/SwUqt8J3G39Ph5
+SNtT3joWYhnt0ABcV2wX5fVuXu2/Bl4jctYxJa7pzwHgafy32dl1wVDw64pmvZS
WVIrnuVwMmDx3sTH/xsYDbphq4MSnkbMklher27LMgQio0RH3zDeN+xLxBgo5UW8
D+qC2QfU9u+Wjjr7mFaBEsc81UMPmZReJfdsf/Dynl7dbbfBQFPGQMarMOL3z2yY
dZBA04lL2cMDT90ValC16rSnqIOFyXbClnvVA7meCl1Ow0pvplRnWPpRPelHm6bJ
C2S0RTfQ8K3kOwQg19ZZIjoBb+N4bIgQdrCSTnE6wuokh4BkaQ8tmjLRIemfqNRN
DXr/mJFXGTChoVjpSBT5y9qvHAOC2CO89MOjdb5Vl/yS0vFoP7KgWc/fmSPzo/iD
Qswftx1PlGjwoJrQRtysvGNiqDRFzSJkeah89cj+XPGmEzjdBuj7sIGwze7fxBIr
EOHTjnmu1zBiAaeOhc0zDXR0CaK49y9lkted+KQndi9LBBVXuIPibHr3Cg+BJZ0N
QaKSTgYYwlAu8e2JetIMP2MYDwwUMrUGCijaJ0O8ELZU0dop0xr+qOLl6mCZu8lY
NCszaReasrm0arD4WbHVAXQ5iPcRa10eUGPQR5SEMGZA33LpP/9PiwGZZOrEaxzC
vLPLDhp1BWAKIyXVq7Jipk4HtFB6KbvJFlMcIiaW+MGALrg2XIqhBIrf2JXuaaFI
2rUehCMunXHkeV6PHoLnjTHRzMu4QmaTbVUxc7y78g4lXbmOlic4QAIfLn2QZsgU
uiaW/aqDAhiSRpSDrlM7muy1DfyUzEeWDg6NaRcRbavh0KMASSGw2djs+DQ+Bkvb
q2VacdGBwHNrmitvkEgVdOFpbmhmuNgPXgtdvNaX1eYk5pnmHJicyTNSKgzMFrKL
yOAhNXkZEX7Td5FGFXqyK+H3W0ClxRuxfp4Dmpz1d28bsXm9GvJXupwsnJeotypt
Dvtk/70M5LXVOrrbm7tJyHyvO8y6N+PnxB9bEM/uy2gRDAQPZPWsm86ebgvGqqF/
s7vqA5Why6Dhzsw42opLCDvZHF4QRzrIpsWq4fiwcN3d9Ag0IHYclPxF7Ja/AGYe
HDkSq0JZj0GYMZzecm2lPBQYMHIEDf0fAStWwHQtkwZ59vLF3N0nEdLQbOdN32fG
xls9uI+IVSwdT1cP4vDXL8tsAg7ZD+tBgqniDdyuesJntS1HTX2S6J1/0Sg2p/pG
JZCJpx8ESy0IRVMqEgrhdNrcKsdMB+uSGTIaZL8s8BRzyCpMjgacepQkVsWKaHh/
7QTbkJ0ZR4q8W3eAJCwg2Ik5KlNsf0rgSfwbSo6stvhqm5IW4zDAy9vDFH1HZ3HH
/FUa7Jv3nikB4Z2idaOMl3g4D5XI33qoziTNxc7+qABdYdlQGXVfsk98l/BQ1lYi
Bc8tsRiN0490Fj/eOWdP7RCt14Gg8po8pqN0fUrUE01I4uHVzG3J5IXemqY6hCQE
j8m7C3528LyaHmfaigiH2hIKno7HU255Yua+kvFQNnqIPpI98MTimsm+qBl0wB28
oTSmqaFTajIBFZ18VPjYNyGofbw1Uvuw3szz9BPerbvnPkLSozzBNNyCozZpPGm4
EqX7xxBeuXc7wotc54yS471jm4boLsYaygkn3NnYOSPhqJdi/dLxFTf2Oqg7uHQX
VjFi9sd//4OW9DqtgYEiFlOObqNy9d6kj79LcneBwUlfpSTUx+LujCZ+3QUl4FZp
YxFNeLYdqnbRtQtWpQ8MqfjSZ7oapvrSilRzLgU0I+qU9a5sBBRn3IBl+cwQoAu6
ibdfomnFN+ypnT11/DxP0gwXYAEvQBcQPkzRDYeia31+Rq+2RR2wrk1Ita/K2Yzr
8IQFnwfM6rwtQyZiImVapWn+2a55bRMIIc92YZj3x42DRAS7chOHKbCQ95hjjfkA
3AaLMAArhirHR5O1N3bs922kZGmLKHBrNlugt9S8vspZMS18+uE9yvwREIhibO1e
zRygIp8At7MRzuoH2DL492XrQqewtblSA2O3zcTKNT4UdkrScKeqxfO+BlNa1DGl
7MuU/GcK7oCOMsTvGemUkN3Qroc6zrVGr5Rk7X/wrwDY3615EvHimLa+gzsbZLSZ
Q+9XUBiZvgH4AFVbbmtiX+zJV6UytFF2Rhs56EYXkjUKbeeTTlr6CMMmN5OanCqL
EnR3d+r7UaEvep5cUqv8BIxG9SuH8h7FNQItw+038KI3RPTQUNCJ5KbTccRNsBBp
iBPdjE8vMXZDFg0JHM/Hq3+BtuYe/1xaF1sX+/lQbxnLqIdB6gEP1fDeW+DPjYcY
6tB+WrCZWGSLCuM/+eWn009If4Lb6MFtTNHwxByub25YL+7RQQjCd9CMm4KDiuMC
bJtO8FHIMdWl7AmJ+LTrYoS89VHOdQOoDU7aKvpzupiGF4N4Im5nvd57Uvq7O09X
XxPuTKJ58sOZrTUUjQGiMWFOa5rRxGUqBPvLbs0oZUTRu8RHjDuQ0cTz/8GZP60r
FbumO111WNgwoZZaOFY7fIesCQxyHp2mROJSNURNoKxr/zubSIKyPbKx0GMe3n3V
QVboxEFBendwavMcV9Z5pjoFJkMsdD2QsohiScudSDWegdYDLoPx/NayDBf9ksDM
BUkibIG8vsJsaOd/zXQWRJuc/YyGsi984iBzhUMwzBdJ3x2lXwdISuhTEMDZkdWB
t3S0yCaCE0doMHANR/RsaJa1u/mmJILo+/cjn7dXlYgWc6DsDMCZh2Qm2GZi02MN
cZTKUBB3MglXKJs4u7YGd2kyzTRR+ls/QdgIF9YcjiG/Ck28TcQ4wqJ0cyy5sj39
+wTfkujgglXfuBXZvVBbUSfcV6YwmBSJOiBs4XvLtAokQpj5+OJlgc0WbAkLmWPp
s6Ncri8A12O+pJYbDHyBg+UZDlKYkuSjYFK8nTqJVnm+Xu023+oeXAfsYnbDfTC+
npDIi6H0hQsfXZj5gzDVHEoMkkjp/r4b1ndd0jboeeRplsWeCtM9DNUX+Ws+PxLj
qXCjxNHcfpw0F+Bn/N9byiY6Si0LsUfJdWUVEpCiO2PeZWqEYJCzPkhIafRjGnmq
xBFGBu8SBQ1AtV1hCqbL+SQvgtYmGe2bVM/FsZbTKzCL+OLtw1wVDLaqkqFreTDN
PfvHJqUi0dJkpuyz8IdtWbzywlfmvYoLJAF5Br8I8Pl1/ryanx91CI6yJomLNsxK
/mzBn/onlQdhklTtae8kLqG1p4cNP11k0C52AXUDmM1WP0C2b+CDUlcJGA1RGwLW
5CEB4CtlFyrDtt6neuUDZXi/q4WkVaG42ctJEAyheAFoUWmixyg4yF4LVRIAj6n/
WVCMM3mPxxcZ1QTYeB4IMuDToX3i98nHJU4zcLZ5k3d/P6GahNvT0WdYldbI3xO9
HljXHdlVQ0sD5X809TPfo+ITsDL9Is2nbHzaLZMG4+kRYdb40i+NvibmVtjkCzMU
bDVw3+aGekwmLY0XcUE+Vt9UrHHNS1NNf2/RhBwJlekNBi1s3IIo2wdc/YV1P9ud
PwKVzVRyNNHr6zUvJrr+jikl0WcP5iCgQqVbGlj3O6GsOSaBFVcjD3MxLRVmLemR
YVO5z8NiMGgLetQLkqTqhTlp+ehXsHHYYhdAqGLMjgKT5EU6j1T9T8TuuJ9fDgjX
1WBW2SFxX4Ds7l4408aIr6tD2qOCaAm/gARQM9njGTlghVnvqnozn8suy3XQn1M9
wvjDWW1Yzvq5W6R6/wdl7un1wHTaXsI6dR66FVnRUaz8dNRQ4JGgvVuak8+HKoS/
VZ8kfmtcU+AiRHb5mJdiBD53SUYCqHTx/BBhmXb14ZMs7QPUQNjX2W0rfhi6OrQ9
rrzL2NMqHe91yqZCkTg05UVDoBl5YuoXzs6idgYJYRfCUft2LuqJ9ABLCgFAXo1K
OIYYBH/XtttNzod2k1eHOFhq8/Vrt0gs957CKa2lWjuEgX38m6QsGx//qAVmmPxH
5kSWNw3e86GVOTa2ppYVLIWaGiocYwOm90umCGCQIZhLcPBoXB7axErqj7sYjF/G
JsRPV4OXzsWtZwuiHzyU/NsmCj/1gFAg1f5URwiu3EM8G/1LpFmeMT4EKt7FrG60
iyRgePCdpOowtA3IE0dXcQnZAcfPdw4SceQxosDrlnatcNnqay2E9sw1rEoKSMz7
KXOvfMkTRfUXKhhS/lEJeYWgyg8GZPfsJ86HDvhH540Hst6uenTVCHlznvOpipWk
mKU8oAeLdJv4wJEqX3Mu/rNjxUlwbwI4ahiqW1MgMWZf4IgF4VJozytZ7hzYafp9
Hh9ANoDdaXFh8u5fgoJO0cpTWDoavsZjsaOZb25eYuh604noX4C36keO8uMEHG9B
HEUWjUAEYNzLFAE36SPeP4lnqKHCEoWb0fVd7GQPcPVh9rL7tsZKkdN+iHYaL3Kh
JhOXfhpfYmE8DBj7q2klZwisCSX0XK3x2YbPRhEQRgmg7yi9kAV3OssfxD0YSKkO
gyh6jJyzJEAOSICn1Xq033K1U4kvlWdFuI4j7XV+oMZsl8OMUXcJsolmiSDNWSS8
qi+cAODKEn5GigwRHs/7JIVGEehVLgkmI4rHijuqRIMKdmfeUWFlUIpdWYguqG/r
XIpI6gMdBVFdB7OI+Y/ZYuqw0MwLLxcubCFKWrZYVZQpickp1ZSKlcsUDyHqa5mO
QWnImKo+oHdbiu3QtjdLx3KWuFNUIWQDZFGAMecCKySqPFJAU7W4i9c5dmXoNo9M
PVG+EryMePI6fNkogHRvApNQYNQK3ykpAOKnskoKsuBCezdHbgDDmbfMMEnnfL4z
6anD8QqgxgLJHDQqOERcbZImhAKHKZpezJ06IPPrkvP97fP0CvcZGJde24JNa+rN
jPMrqTjreKt7VwrcpN0X/M3NDYMD3b5KEPY0DR6hBpcMKb6ZKVTv2QnO72lfIeDC
IcTW52TQz7lhPIPOImarAyE9sogEL8xzrtC8sx+XYf5gFBF9uhYC/zfZTSZUD78Y
VYpzuzuFrPuD/ahyCrim1UnNsJsTdEpTO4YVZYDAhmYU11Ia4acMJLnt1Q5qG/6d
+vFebopWY04fG5toZBh11pApTRPqz0xnH9lw/b2tI6TMudAyzUvZreqDeEXW5+q4
7o7nVyHF+uSNjO28mGge5A5qBZabQX/htU69+PoE3Yuf8XMwpZScFfNZBc98RlvS
uXcGFm5xx8M8k3NkfY0Ky4nDMZDn7pB7asHkTzkO+XL1OmCHwsoh3YztWqbhuKH/
utYmK3WVMeXJmnflZJItJM7z9wpQZB1ywQET1VeLsXGIG3gLlAf0VIeOfki0qYoT
7sd3+qZV3MmNKxmUoF2LaycUZjS1z18ErwUGQ9twXRLZw/ExvvWyd9BH20W8STrz
5Zslt/YXWCAksGP0S5ln/n4coMa+/gZmuZU4YSLQVg+c9172K9Fr1by8O/bKEEza
ydrN7LGJbaDlYQE6qO7imxthxbQLSbbms48Pitlq+xfFKpI0dMryui81rkxtAgK9
94AWaQPT63XH79wFBX6zGyc/nTZccUy3hs/RVVIdGEQKh1yLdSGTcqjVpCmmiG28
mhcsSSu6cy7dAJRRlZbcNIa92GXjyuui039ZFMwb7KTqZg6p0L/YPz+XRizazeuT
BZcAVPcnHTZm2SjGfcQgEP1SwcJqgzoyhviRy5vsF/+K35yUEqfCKJMIwzSTGi/l
LvpC3yb+RGnzoFsgLkh/Tw7MbYMDt62diIH4WgXIvuLZXv5g6leM1jaNb+SCsQdC
yMX7Ftx25fI3qSB1si1bmkJLrCUXT65VNaEJPas1/Cmdq35YxF2ZL5ZsbE4rbZEg
vSTZ/uN2vgt7KSNOnaLYbOXRo8tQvbLsKpV8TBAJiMZ7OT0pgZsq00XarskJ/Nbs
5+gs2tDqV3ESd79pIn8IR0cODjQBzSoO8Zqw5u7/tImNjtK6TYw4b26+7ICT2rGA
epqkDvlxsbRpgfJhTA9tQVz6wIEfbXdPZP1yeoEGMUPLjLCmWzZz1P7wbXbEj2UP
PRyHeQW0ZYpX20j5q+mtyjHY8GgOqh0owlHJwqyfm5Nj1PvyQ7mxCsroGPu3ASZK
gNTyaEB6cz/SrmR8QWB7MFl3S4LMeB5eKhRf77ivx0QllGkPmHg+DtAc8vLrhgqx
GPMHkeqxN/lSSbxER8o+f0HYI5HdODyL+KxKCikbbyQt0gkffbvmstP/lMc8VGqT
qAdkA35afAl4OX+/+/SpeYL4ruQqLX87InWr2LmCGcoZTjvipTRm2o7VaA16oLx6
n4QrARAz+5lWkZrc+AsZasErI7Wn9lUfsU25j5fn3Z2/txnNnTKDyYu3qTQ/JPzw
7yyHNtN3ZxMb/vW+S6R4n7NppB53PmMOlzbBI57brReeMyY1Mw9mZFv637RbwWpI
rgLhFy1ji28UlW4bO88ryGBYd2z1qvZAfS5je/vH7sobf0HHARZsO7rlGBdhRrjp
1QrSCM6Mi/285BWZOvPn5CRnPYA3jRwAwSn03NwRsTw/s/vyB1dreg0MStghpjOx
UbibNRWRrI/M7dZ3vAS0Ma8BzM3iOzopQLIg5CDH1GdL3V6bTZcOCklHM1YkNN8J
D3Kh8kLH1jZGt6iTN1K14nF6Fio+WVDoBL+fZxLmQrtoRzsBAMVrrpaFW5QE0ePb
A7pa2CoH9+FQMjGusk2DHjCi+L1q6+X3NXSl3q8+FzucIfSy0FyjQn4WOX6rlb/Q
g4oQwSNswgwpHz23zuPn4yvhDKanl8qL/YBPcub/ucnYoZGmZSg2/A8ToPU0rtbl
MK9vQGd4idhjTEyB9NzJsUF7GF1Yth6K/n9gOw/sr5YnGRkfY0ExKa1rtcWBeLP5
+U/AKAHjJRRKEnEDTDJhSeXJQh4+XvoYKQoYXhoEyk+b+9L1xUpcc3I2OOoWYj58
oask+YG/yMVF7PJy0/QFHfhWyCAHTUX7XeO9H0DHnApRZ9TTChPP0HuMS/ougnog
CRjxILR/rQAzJqudCJVEgwIn8MaciM8NjNOFp9HM7V0NEB251nc+QUZmZTeuL0zt
EJoFAKZjTGSmy3W8atC17zBIPCmXDx1HOxuUlrQlELoAmEfJ/GhphQR3AgXitSfl
4Uk+WTi2A/d4yxplPAuzV8DaX1dmyE1OZsNohXD9LZWPt4uujySm/pRLrCE7EhD8
Cdx5xCeJVrrLWJvYv0DjuTYQBb/5CUwmn7uC+X3Y8fqv56tz0NBqsOArdkBOecX3
v800NXohjCKR+lgC17EpcRD45mBODmmlGTrp63FvHF/iWVLvFqHUEd27wMGPkRxV
hDt3XYUVKOGfXdyzttBHFUhb28CFbZjn9RSfyc+sOLc3DEvDQu76rTDV71bJbQY4
fVCp4O7kOikxbm1yxsRpNXxEmIh32T9VEU4b9ZraRiEdO4Q7d6NHisnSSXOo0FEf
LchZnJ9IZH+cHro0dXUeYgT7vBNT/8b/lLtI3RV+y3j5S2i9VPZLy+cKCt5rm13i
2abL+CZ0VW6DjwKT8nCaLIEp0Y4vXH2+zLojZEXx/uO1siu8YJk06anKufrghLae
Ht27OH7Ye2eolb4eSiskLQTpOlgU7qFm76Op663IyPSoeL2MpDMzZoqh+ixj49yZ
2VSaRt6cFTV1eGxG76AvivciU7Hff/FsoqfTdSHBt0jzZ1rNUgk6beHZUBkytxWI
sUCUHtP8ChiBdLaOspEaWOgRMzy8FKY/SQWwIb4e5O8xaU+G7/Y4cs4Yu1oNgctP
BLNMjpN9V/wOsxpXfZHlJZVnRWRmf0jornUN9rIFW42z+KN49ipeHyYJLjPKSOao
XV/EBjpwnVagFv8xqa8nAdAl3wXOn+qECy+2ec4aOR03K1XQrOmRVVSqxhYMU9hV
2WZvB7Q/tyw4J4ixV9tc5ymgG9gqG4HTOlrtrHRtTGbkrQr41+NyISG7pQyi1I/m
TBWwooak8cf/okzVXcToarME5mstxCEAVzUkRqL8uvoVxPvMabsbNlrp60hOz0Cc
YOMKiq09k7Cgo7RVSqHFKDzxiHaH+wo/g+Dthgd7vVPkFwPbbcRBcVVTSe6T2WWN
Y7uiyTX5H97KmOy+HhnusVdsfaTY8umvYAIBlOLmMfZH+eq93khlJsV0Rk+oVg7b
OngViobP/IRLfs49sfO5Dln3Jcbb+Lzox4Mg9Hs67POLfKqUZmTUhWt8vAgRdNdt
BTdR36PrhcCQCmBmtUOCwNeUXCgZM+IELH2PvrnL+A1QVRCrU2zsv6VLuf44P3b+
jMu8AwJuYtPapEup/RXcMqMC0FGL3mcu8A5mUOKtj/UJQYUq5HizuYi56KDl26Iy
mVb6AzL4OeR2+RFda0kzw5d4WcQVB9Bicv3Re0m5sThfFuR+OZa7Ph3RiH8aYmYz
nIauOoverSX18gZe6Etjz7etd+Qb3Kfwz+fUtIxxHEsHq7cm7clHi2tvyaGRSrvC
j8yQPwTMaphTjebnDr+IT4GJmZqWjjm/imu38MIgUGmSII1SjYwu7qSNSTBijh1T
vZ2fukvA9sD8IbLUdqhb08kOgd5sAntp68bYsx9lll6yfMbPwJNf229Z9hsMgKvL
PKJhMoCFj1ljx211aMASOFqZ4BjAHlTJAJRmu2jx/hXwD3J+bnDBIrKAsReEDAFK
PFvaATos0+iXHkaELwHXPTPKz070+cLt/jZEXQUFuVw2z8nPoQ6se5Mfpqye/ReD
XSok4TVVWPnaQCGFmn/HOzwStv8vjRR+Pc1gSqRF259y1crwPAYT2hE+ansebg6j
gL/sTcXk30p9JK46j5MCtv7XHjPj9AoCja45skXrS4EE5CjGpGYjqUtFV575YjlY
DSuVZg+D79Zv8XEBrQR82HYtKyjfMQ/ZE+hq6QLRKo235DY2FTFPBCTnyrVfGWk3
EP1CoITa2GPmLpZoIIRh4pJeZVtSDLxeR3NxHF5rxrv6Rm6h+WG9iI+MG2ZWhmfA
wyxgX6QW4QK9mImmJrB4IvYfBjpXrx/YosTFjRHaUrtlQF7fIIWX1+R3aHH2AWJD
gXpLqoUaezAxwMDZpmCscHYQtNkD31cPh1k2VfSRPREugvHxrMRYOsLXqaQpJBEF
jCltSh/CreL37bF4grAvCgnAbUErd4goayMboP6TmaAvOQOBak/3g9OPtx328MpW
ckBMJCVpYs7R96QF4wxNa4NegIRaofStlpdr4xZipQJdpAIo8S/yIO3fj5GIsRKl
oN8AsfwlRhbtBz5pzZjDclo4xUDTY/iNherRjviEu0Q/YaMBVM8rLA4jcTNfxluH
0nv+ffcykinX5B+9aq9eljNdTA0zIWPiFxJYWFOOUyEBEdi/xjd+Nb5ZIYJfJNjI
2S1yvOxRkTYv+V7V4wf3rUWpyw4sMUnGFS2BhztBRnxTk+rcTYZFNqb4J8wuoMvF
mp7Gqk2rNLzN/5p181YxWNjZAbCGz4zbJk6KzNnjlBS/LOrQIxRIuaTV80CHSRuo
CaLVavnwRSveDfhHJw54/1RVwh2ocKyUIITfj3lIOjeziJLKtfB0v4gweDY+n2SN
X/LHXxfgTDVZKjj4n3uXyruI0KZnFB8sURaWYq6nKOc9nV9KLIlT8LTojFxoM4Aq
dGpVudCgLyDS/29nyRVPxpVVAfBDGdo4U4z/F9gwOW6eW+CsHtlCYeZ/AOixcF9B
Ly2F+kf3P6PxRJG/lxHI0ceX1+Ew3U7qvdfm4t3GE0Q547vlXT44+pWiquwIKGau
+rtNGFrWmy5KEf09s/1yJKD/fAghSQ3ZBILFBcBAaFedxA+kqg6OxlgACUBxYDvi
NFexirNSeG9LDYR5g2Rzc94y5UytSbgnFEkiB+yOrXSljCDFqDqK+WSxrMbC/jku
kRCTDrSacSk5Xa+jTfeQp5MzVM++ZNxDgBv6zvi6rnf/AW+oB8EIjBo80K6w55fr
YLh3nHMg42AgqYqAC9BnodmVcX02Q4Gf0jS7R8Z/jMQhM4jbiNdOIr5NAHRxxuAY
l7dwDWdtMinKP0R//glKtmG2q/shl3UbOVOw6imE2u9XtVT12a/3fRXp5DCq84CP
C9bQdD72ocqNNxo5FAvd461sFLB8cc95INEmgliQ9KrFRVdsWZKjk0tYnomcCFut
wox6sfzv7bOHVjh9YHYAWLuc8m47C4iAQW37iaojAC7ic89QeWk+Rdrd47Tcb7Ww
H/IQVp2g24NLKhSIYlp9bx1jyrCIL8jDfclkn1EuAvpjyVBFW+5wwyiFE+3wK29X
pPFzwxGOZVi10WV571BLoV1BmzXAUXF40T0faNO83aT1zRb2HFQq1zQ+521xExi9
Wb9OJDG0NFmgPQ+pq8XSuYrYBksu3Mh0Lt7q143OPT/tzMPfccURfSDAgqG77WnO
1vctHFhoMomj83I0EkPV4ZI6fqe+B8NEdpE+jjxLHlazO0TfX91JOntLTF70sHSD
6UgidC0bwmFwuGpoNqkXt1v13aqNqaGPzhq+NJUIEXjQwIRtAaYlrGlvJBmQkehh
PtvP1uJI8Cg0v2QvypK+Kv74WM1GZ3Wuyp73iWc9ROiCZynK/VjVKLvFAkEx5CR8
vEwlRDkiEIHlxdu2pNPaR02OC+Lov+fpVM76rw5MfE9gSZxoiRePfZZY7vrIxU4Q
s7aU6+XvNoYrLPf7FqPbwbjOinp/H9ebZjCuiTK2VZrqlrgdLpBrttzvToTKz1FP
22eTVeb4gy3pUEPtQ6RbESBAPKOohpcFuxttadphdArTPxsVx9ttikdfrW6r22/3
gb8R7JxtioJ3IBusiUvr8QXdEcC2YR2H6gt5fnbb4OxisCLxU4Tp1uN746NElUJM
ldHA6RKXlfNLEuza3SAQjpp56bWYhT62/dPsJCMYNxQWolN/RHZYrtm6/SiVMi6+
KH93mQpbGSsUuiciFV6G8GZ8xoWazhAK99YQz1OLAmcfGqj6EMrVHAIdM28oDoam
vsygj81Bj1e3MnHJc7pJ5a9oahn1b1ke8mos60Ry9yzxqi07Io4Xptku3VkxjbrN
rgbUUNBRjJkryQ0anLQCoL1cFT18YrsXujrCm6wclg4FB9AVycmSitH4/1Hutm5r
BpJ0pBxWUO8mIjoa8+J/uQXkxZwK2doHCBB5HhPisoM6yTlSGll8BLG8slN2WY+j
QpaJkCmxNY3mNzzGmBYG0OwR+Xplpic1+WC0sqeRnlfbefufSf31t6ZmxiKNE3w0
FaMZMZCtI5pBl0IxWS9gzq8IdajaYCZMhHhUTD2iyEIbjprcSq8/u8OM9nJGwKbC
Kg0vGGWcxGuyRvL6jWLVAG9xZRbOoXQfYH6wvU7FlMl7bCEgBEnTeXCbTlwMG4Et
O9LtUwBDMi4OvDhcCyWMYDssAM6DCQAC7n/Y0j3MUBhEy6cjf5SSszJT67Mb8AcP
hy+wSZVFJK+OMrnXn6U1QuBK/u6V9CNK/y7uhonve3D0HH7uQj4V8St5npkY4v5j
VrC673rBV8fMSajjE04AJ2A0S93KXHiq1fu6LmOYkxR+EVbs6k+qf9Lqg46Pg7At
LWtacesv/TTaXM+vYI69/OlMF5azYZUO3MZweADOBtFBZ+cBKnJo18AmSjmfBale
iC+hjHdbwLz+ThSrrZ27qH3k+Cyu1sIFB8jD1HB4nPZzfDb12FTmoARhk9T8hgAE
pMBN8t22qcir0//WuVsTQCn9Z0zPuG/orw4rl8pzTNjDxnhQvnoHQbGj2EYZcmoQ
F1k6iYsVnMhnT2kzEZugraqWw7CoVg5zFalelcW2T5WTVYAMGLTgzXEq8D2h95tU
vbLPqcI+mo0BiqCPTfps4iCIpPp0zrgl7+f52yHHKeyk56BYhto4wXJEFnlXMrd2
kZNM5adOLA8tuja70dpNnRFquuLHn4dR5y3P5+PE7VhRp7lfgN7wSSqhDYmGt2rl
By6foytdcUWHgtOyvYU+QPd/erpRX8PSy9NVA6xKXbPZZf/1lu41Rjkunxfk3Z1x
Gz/cSU8vydNqxBAfQ50Aa/R/Np4KQg3H8L27X0CcaLJ8oQdIJtsjwGQIi/bXb7PI
cvmlLaXK/mVlHNapgPpbagk6riG3CMss02bbT26qlCrAeTx3bJCOr5jRelm22p3M
YLwGRH/602ABuqAtotL6GqQvvZVpYj95Vx7Bgb8PBMLy3CHsWKb41Pqq5p4QHP/5
mo3EKR+LuuC2FYJK6KVQ/gSbKxz3T7v5iKsdM43CnhGVb32CilAlTUB9nXKTNjG4
fKHr9jnENN2XCc3b9BpbzuWhGfN/YgKTryLQo2+T5VtHv6CRLc28QykLRpAjVji4
HC/VeLATbsatqn9thcMyqX1NXjRCcLP1HiWzb4dRvhSp+MMCS5vA5a8ssw6RaLDb
2olCLYtJ8etjWfQbBv4RF7x25/I+pMYOZgEQ1y+uP2NBSrfgfns2p9v6Z+PfdqvC
L8xPBiQDaByEhprg1ObrGfr45G+AFT7CCOyBMTu+0SOtKh1632BVSpqRh90rXp51
cIr7226Wdz9mZv73ouzu/6Lp0nHaOVkdtNqQhY9CHmSXGZwXWiAtrQe81VSTJSlF
0oiLgTWSSZBr0iMrWnGLvN/nGdaaHYxgnbzFERANU/nDvInRs+DA3nl4aMbqP8GY
J/pdOmf5hp+OQX/A/tQ17VKq64w4MvROilAvTuBdLnZagJ9/XmVS3YmYbVhIMCdL
fiJV8a0AY7g0VxDtLZCUWcXABjWhL9OyL2Kg2z6yLQ7BsGqlqmrKYtbc293N3CBD
/7uvj+ruk/CvCQ3/zkprtQUW0BDiDjrwUzxIUR826eGO83BFDRzcWEejArPzQTCF
q9DoYmPk7k7IKvnWli/X7Xj8tR6Tot3oMuLCOTD4+f4czzdYzA+LpfXjCEZDRfp+
e5MmgQ9GRy0TPXpdwZ4uUuvZ+l2Kq16OkEBiK85QrnQd12Tg8xznD2IZSzye7T52
NvoU4uq1wtml+D7dZNqcDTWoHtxiHcEA+rKb5vfiIt/pNhU6iQvHKzn+g/YLlGTA
JSGxu0P6p/I58UTDl652IDvo4rYVzSkXjBLy9hgffdlFazSkulhR/XRRdER1aRoU
SI7otTlNsImpAwyIYnRHaIOnwoa+yaOw714KSid6eBARuPImTDTNlbECeOU5LpxR
SrznyLkL1hbb0xRjtVK9coBbmuUbgP3mnFo4/isqgT0ojL8Vx07oEpM4fQq93d0S
Qjw0ZcCxsI6CNQHEtEC104B6JCQBn2hrBYxjiarmAvlnFQO1FnS5Tp1oiHHtsmQ3
p+3lj5P8OKOAwU8sEIMvg4W5z8zhXhXLo/H26jPdhi9f7uDkmTS735rpwchoUYqE
u9bbkazmT6pfEA2BsFmVhh6DrBSDxp3bcoTFunvfwNITvJagnkvhAb9g0RbxdnsD
uqsYCar7xwfZSoCOxV4xvTHQ4pG02crJ+vM4HHUaUUiyzilG2IWDK7V9Xi+x2Ozb
P+KOyGcMstwMeXTM0f4Uetwwf+mK3094Nup+41IopmcsYaGA00GhHkKauiOhPZeh
bmW6icbCqt9mdB84gRKYbuCT64CIzVK4Bx/AeJXFm/Qa0yfdYEE0Hy5IM7K2wBPz
ps9BC3kuRIqsJMwq19ilqHQaGxFs9u/Yzs+5FaZwXG6O0NkkeAJtWA1ranDS2I/q
8cE7BM/RlY5Mzco8PssZkcwsH6xxvsxkybOV6mMtE98ChhN8kDnqItvUn8RmgcT8
5cM3Hr6et9LCAWuXo2Cq6ceSRgkSbq4GMftmQjeMapVsIdxlI5CMjOD7YOSf3J3z
xiOFu7ibe5OKzaprZXnVOjJSJgrRWCrKC9Z/j1J1pTxUZ4h4jxF6Nv95/Jdvmb2U
Y+8P7P69zTi2Ap7dtn3UiTppsccecwNoVtfJ031biNw8rR1BWjdagEpqDduoYUO/
Vjwn+3UokIxc5kb2zG1Zma7SPJkgYRfZtziJlExsiyhxM/kGetMZIF5PjUc9YYYF
y2OH4zktE6b2bYZI8eHKuEJOFrAtMvD9zhMu+naZu0slxlhSqcaPGA5F/JtBuiQI
WaC4LDcAhjfBt8G1PUGhK8O3dn+9pzp37ZCBQ5fwPfo832VTWRYpCulF3QJ0Jtc7
QJx/7VGHRNRU73lok/xGRtWTnGXUiQIq6o6brTO/ni6vCbB8BO3WJG8BjoR4mjHN
gRO/VurQn91TZbUuFO2xAb4XoMVLkIFwF532fuztcFGIAivMttF1wJ3CmzwdahAI
ChixKlj5HB6JbDikU6UhLHGhTFpW/Ztj4PQv2WulsrmNqSRD7xaK3YAu57UKZ5A3
Do0NiaEImG0C59fTDcNbDi4mydY18Gjmhq9C9gM4ScZnqHg1CtxBBojHDYalREkD
oKqb9YHi/ex29pVjXcP/RWrxRpkX4i1aRFssqgo3ku/SusM+i51iqm11wpFPVMCW
f/jx9NafqbTceO/8AVJJmOQ1O8q6bbDwYzVWuMndMA1DhQ1iZTtmn3S0NfAIbm9l
s2oqGCyg8mEiS3gis6wMBwwQfUoh0szwGLVsDrK+rTpc3dKoHHWVieOk9FBI9Mc1
laOQUI89APpemNXhpztVJ3lZjUzFTN2QTeQ+OosIx77uBbx/suI7//5tIesZacHT
RnXfCG4FptV2pw/o8FAZ2mxQVR1YQmijJrKcC8Qj/umtKBeyN5jfhGUH1rZyWEOH
FPpU3e9XTjeLDfRoPgG0S/Nj9oUVeNTnxBGKhk/dZWhfFU9toiskOGjzjeNYsnIm
fjmWqnSj4iYyeysH434epTLZcfRGwkKC0Amcee41bxHD6XsOujj8PVOS1KP45y9e
OJ3QiqIQV6uwLiXr3x6D5EfXZp93FSXJ9r57dhVhmmCMxPjamaDGeIcWYrgH5FSC
qYULAqupRg3gt+JDStqFPnfWFsdEMlCJXOzp2iUOuYy+NgCQYJ5f2HNvEzR/yXzo
nOnmAjdITiBG6jzbWhmDo2+HvUX+1C1iESJu/IDcJ0Ug/XTpXYms8L+YwnfyxpsD
dB1bADRbgYdsAvAqpxudNpnVwLtVAqtpfp1sE5XS9poabtsP6+kp3ACFMaDGbTh3
hfASEL/DnJ1AoDFWPg9QqWMCw/cNzREhHeA2xmhm1wqJrAfVwVjl8+zBrbfB1sry
WMO+qnS0fnGzCTNnE1kIN3uFEYe8qEs5O4ztsLeHAQrPHlk3GlSdQU08p76hg48J
gruds+RZGAYmbmBfjXONEsvdPIvHdOzouWT7reGUsi9Kz7mcMnaBfaS/QKKw8J1r
IDE+wekTtzFmGi5Ey8vJgtkM/qvAgEgWPJ51qHdd3pnDZxuf2I1Tsrhn40Hexklk
Ol7fELWsK3ED+Lap5n8A37RKgZ7C6mC6FOJO2zRpkaGCQ8tR1xpN8bCSy0/qegcX
14LXWmNKDaQ72NcNJJ/kGYHEFzcMt3l1Ye0hr8f4w4JtXVPO8Ki66E9QWB2qwOkB
orHxI4lN9NP2m9Gd76qnXwLbX5SUZQLVRBYw+lVYIz69qWuwNW2suscD7vaHVQzS
0dCi7rzDAeBaEGnQhu4qCrIf70tzmj+OsvuVKOk290OPXasI9WYZPyiET/Mftctb
13Z+bNP/nX4NslDEuj2rdbhUhZsOhwOI0qj7gMDkTOImWy8KUSq+iQi+Cm8eXA61
T0o/V25a9KnpelMQRya5Y3nwlqWbD96SkRKjyQF9BLlOiPxJe63p5kicdH+WqP48
9DvlCnG0NkPjS97GREUQudH9q9SvlKixD6HUVZtm8txuWR+5cr5EEpqkDXF+9tjy
nZzz8ris/pVegTVb/xgE7CFydnGHNrKZmOavyKt32FHh9jvs+0ARGw3g0VIQCLgL
QtBkgMSD0wbRGX6gZbqpyCLhvYP0+Epssypc8Bf7VsZXjmJ8ZVW//v3iPztujRA2
gJuYz1pAr07DyUwJ3xXYeZjrj5AQAE4a1MTYbifTsnhwP7rDcuUbrfadpZ536mE3
RGCVxDPVZAGXyOX31MzX2Ds8wPNpt2NDdCLmKj8WlwpC/zPh9huSum3DWMZfshC5
auvhwBYGgTFh7T7mOwvaOQJSjlIH6Uu+o1sAQiC/vmjS7KWPklP4/ubiV4XUvtfC
5/w/uhkPQe7r5AwdYSR60rYdc+RdcMo5vGky7UImWVHR0GxnaDZY6UO4IrnE39TJ
anXUgk+lnKefnaZrqCFZefdwTSHUcix78HkxhhBRwvba489DACQJa9EPC9Bf2ia6
RicVg370P0629tJNlRpwUKDCn4m9f3jG8+5hSpstwUrUxQdL79vC6FRE/+imCkqw
VPbys9I/qhRfO8xiQCFgzAeKmdiBLQto8QwWnHnJYgIM9M6CK3mgOa/Sb/6ik0bI
sdMlYzMMZODCI+JHlVbBR8T8NBN5R5muczWZEUiyZ+EwOg+C00SFQkQ24TIvHKJF
OBon3GrRuB7Um1hAeD9CpQUarwHeRSxKjilLIuNQGOnrp5UuaRQ6+mDZvAfFvdkx
hHDrdr7Dw9CVLzNjku8h+H+8d02CCsF0C+my7SZdrfisjF6Q10ZEBFTnI3pCwga4
9LUn1h2J8bBhLl2CW1qPq2C7oHC+n1TveEs0hptojefzwwdRHfXcq3PLigveTn3H
oBQMbMXV2pc4oYazQfJZ+ed39DJ/fWJ7RJeOu8CTnxLxD3wSrdXJM3teX2/P9Syq
85riDS3d9gmfVU94zPekGUjNsW7a/UuhUyUDV4CJTks5FMQSXGnI+LZZD3TYqrzz
OIk/zjVfr8Fmm6oPzkokCldu2iErA/lB4mnk9a8KiYxRZUnSnDT2Y95hDOns51Aw
KZSkOSB7zOgN8Rpq3aWJ+Rtg9f4K5/kDa2wkASwqE/y1ywfhad4K3nRxMImjC6yr
Z2LzSLLRAl9SGlPyiR3ucBSdZRT9LI7rDcWIRQByHLkrwlZtzPB+zlHcQv/VaPll
am0jvAHMKxItgv9RGSvqx/q0EtEYXQxyVK6HyAOQ8pVce1+BLU9ClRk4p3ogArNr
js8vMZJwZBi90JP9xlGLrxc6MzoeSr0w+aGTBoX5Ln9XJ5YKfyrVFkJV+zVESTpG
obAwM/cFtweSvjV2MlgthJpc69eGS2rD3GEXaPKjELh36W6L9wEJWMvNoRIaA81U
PecjXLVRzOuUoyJRmBj6FIgZLan4nMzbuxVBH4tNB7FenUCSgoUa9Gawd8Y76vKZ
TnvMAwm0vRw8fXCCHWE4kDsV97GcXs45IWH7FD4fBHVs6xWcRKehlYrQWTxhLBun
WooJaVGt3etlbSSF1vLq+IlbqWXjyYOaAznPZb/OKjAzxvhKGfM+rUCvWtYwi5Qk
aD680TBJBNe5s9EzI7uQgMOgxCi7C0RY035WKecO5BQR9iqSxlTpkOfEkAnXZ7f1
MlGxRE9AJZA9cr7mrx2pvtVo2jWpMjW58kjEwO+Go3BKdKLhlXiyrrzcvceFRaE1
ejEbGv6q9sul+DdiwHPalBw1TtUqRbRIb4Jvy2M+WCstFlOSGPmlF2bYx9puXqQc
m5uky3cf+RhGezH71mU5EbhKVQw9vL1y4nGxLY1XuGyAdLne+q1EsyP4bukdSrwV
mxdx1XtGL6Exs5qTnvQFSvsU7sQZL2Cd4X1l1xdWphapHYc0NVltnojuBXNJKVA6
rTnXrEdLjw9n9rABm/YI15ZaS+c5vK9dK3Ihmz4rYQBswxmRkRYu5xNJ0CbkWsSy
+kvMmOt3SAROIKtVZQSQun1lFD/Opmf+stIw6LLTN4X/U2Ne0QZpFS/9juDou1hC
plNTh326iPW3V8mbabsRhZsHpxz03WaFZFJd8w0uy2+QrPfzG56rdJ2GmruiiOZR
Hd9Te1KE10HaafFPlVU4AVRGUNliKpSTdpDVa3KS5OVOqBvNEizmU74Tr655foVD
cPsBr3o8Sc6eyBivUUlv6q5yZ1M38KAa+vzLhQHTWfSR60S8dWeNwgrUKzOQ9A9t
WGs/FxHfdSrm5ZR2saf/dIJ7N/xp4ubwUx1fmaFhlI5xeLYUQgstxfUvMGK/N8EJ
l2XmN2Uyx5GaaeEicyKMVOrzzV/fk2d15oSdwlUlBuuX8X6MAVi2Js0kMqK+84lN
/x0DgvAWmJvSnpVPDjNmru/KYRTXLMj2EUeObqg8XkZIbxWlBPA1zQOQ1vCl/TnR
AetSRCiMItN76OIlGe23Hs3JMxai9FnYccS9gnxBC+i+1GRLr1bJTnxVbWdyCxsX
Muwfg6OA5PNMqTo3OSCgACcfoZwmrbIO6mrU4w0/Ua2hzL0FwpGKSJwUi7oKyXib
50C8LgYH4cXnEiUrN0YNZvizfpYMIzFN8Zg2WGiKBsYbFlZblJaj0lrSaC5ck2u6
qkvfaMG3LxivLZnycDQSGvKXQQ+RWCCoYJardzWWWEp8A1/yQ15EGSafVgdboZ8Y
ZEpwlaxONTfZLEfCBODsXAmK21Vbj7Wyn/i9Ki2g6SkKivOwfR20/ieENunq5tUZ
UmAJyImuvg/UiUqVM1U5yvFpsaqI6GGcajrNGpuNWRHWbMXoL28ARfvcZiBtCjdu
80SsAOivNAn1hpZh+trWd62tZYNqa8XfPAQGo2GAE8CrMIx+IzV6IjhfoPudDkh8
tn9CGONj28vZmVtp0mmY3rzv0SnNWSjV/nZ6ToDz4vpzJgyVbAfDQM1MoO3V7q8R
2Khi/++8PJNY5cwwo2+vzA4jLFWH1afkTyIPvLwE5IvSBAnUOXP94KLmAIAvYNsu
g/3CH+IYBFYnSsuo4I6fbyKgvOH44nCuN9CdXUOGC5Oz+jfLMEwJGMeGZkMHZfq2
X3eW57WTRvkAX2RI6evgsp2KWKBSxx9KV9uI3MBou55VD31FqRN2AWh7mvacHmdF
SJ097Ww+OB1qNVwrBSaYzLAz/eDCZdktdkEZ8LRxN3/m0fczu7g4hOJo18mFN8TM
a6Hj3oTyOtXLzR28BqtIZrg9WGjzEXQ3rpY7eCG1Qd/tHEYqBzE9Sbzo4mjq4JJN
376Q+ly4UuZfy2j650vJaQxUuQLcg0pL0IfH/qdDkFW2RsUpTEwXkJo/qYjvhuFq
IZ6XoggCW4kIsToD9AQ/CI6qagBeiilw5wONtHJkPfmICy8UXmcvr/ASLPk0DFY8
BN1wgm01HHvu9unaOdf3wAlquGYFyw8a4wrBsCMvED4bMEym1pIodAX089lXz8Bl
6WYn+T9ZTKZGLNvTa2N774vTrQ0YrGgLEj+vgXaAyi6wvSzZl8VDvfKS6Kk5vQVT
wSJbDDNIU3XCKiN3rW9rS7bKpU/WoOykeniviJDOTgot6hvBJj81lvrG5ldKn/yY
DIdb2f+HDlqYo/17c1ECGjFjUfJpKiChsHjxCtmUoJ5E/YLZ5tiVUeIggVR+3d81
SScWn5D1YdGN5rU5q8/3S9zQq4kodk+29keuoYX10ACmtRD/i0hJbgrrpdRNjyg5
ZY4cs86zRc9c++EKJnCt1RHBShMsFR0YHNIbpwQN/jAW/goBAuQR+BD6FGJJSeL6
4kZNXI8k8UJPZ4C10c79tN2aTnVc37jCk326iGl5D7OxUUXn2Ol67RJOCpHjU62V
uk9Wq+e9LcNpj8XdkR4DZcatQp5ndc0JdR1SrpQQJ7/zzkuZd318C+qFyReZ10YJ
0RfOCc8xUGIlFBj6WEU/Iz6OPf/bufQlbgM7vFssQTltxRXMKe8xHuiBudJV5ayN
Sm/wBfdBNClDYxMaQKLiEDk5peaK/+ggk9Q1IKPBpAGmQA2lMEM8ZOAYAzZvyl+9
2R77E24ttjRmE+/UzYEBGaE4Cvx1Jv/lC0F8pUQu1h5XTSJN/Il84dhGE1GWB919
4Odpih5sa04zLMsY5a/YFpUSt8NQbR9/yuspClmJ81Q8FjOJE9tz1bIBbsSXMYFL
SHP5jTTmsMTAtJA0GbHEfgLQYe76pxb661ZpvxQl1wxBdATbG3kZph8ybbC6m4x/
+YvFj8a+dME0+wHKi7DkHSAUjo9qLh4W2nzzVwq42DlVO6czk9dQ/kYwJ3h4riOL
8FGhbRPyJqu/FYPnho6KeOM8yzWfQqVFVsbs+OZDVncx4QWI0dDLDYYaEP+vBHwh
F/T9Aok7zKadGTG+o+7ysp7/0jZwZbnQE2QYHuPqxaaMmTADIw4m/xGDEX5uyab7
FLOJ0F3v8b4f+i1QNbrLmAM3hdDU84O5a5kth7RuHwy/FJ+dwX5F9qWLTMYczKJR
t+WihW7BlmCUzLDmHAuTkuBmGQQIffUdM3axGR2FRjOg8bImQrjp3h35klTaYRqm
qh7yGu6suH3A1i/JkCWNGtSqBNCdt9cgyavRVjYXd/A1rgxIAIsAQGC/4myKtp+Y
A/CXGlWiCoRDT1l58kCHMbMa6pBRUApU9GZ0mc33lbAs3OstPTn3vh0GyX88y5CB
yHiDS2GCO60Q70H0SpN1dMvcAZJioeJ6NgfQH7bep00u3+ezNSFVR84Z02FPr1se
vyM1DVDSfEYBK4M8fJ3CuzWZUgDhNhiuuWhDHLxlFPDDDmM6xO6k3UQIOVdKe5xL
qjvi6QENyhBxclXD+CRRXcOi1jqutf2ua1Sp9zn2DNQIdDlfIO8XEFKooOoQz7Zg
tRM1pN5vR4HCf54LQ1XnhNAioxQYTcqt4C1UiTmUbiOWMh3A23tPwP+wmZs1dnZB
+X0AzmN0uu+MhNDkTmdOx+DuQwr2L/pEYRE/l0dVaI7GPxYXefjxoWpWd3sG+cNy
WqmloJMKDKZ63JYC/+XzRLmh/r6kMClBwHR+I4hLXe/BMWZUtI/P94CfadTOXtS7
qnxoLcpDULAT2vuX4dgwLAtG2PM8Da6QfXqdg/YUIJwhjp+fwcVB9NjQKxO9oKIW
AdI+jqH+4e1nEjnwoCPaQ3HYWB3W/f0XJmmXjAoZkSYED2qn4gHNtnAun6wvMmBQ
DZr35fsNSZ+2HwRNzmIisO7JQ3pb7dFQBocz6DDtVXJw8IorJfm/2nEy0duxr9+W
DJUibrNAUUdKUzFQh/bvGwbNjSl8tM0IlhOlrZxi8DhYy3Zcfs3X9YXGJdR1MiPa
gnmJyEh/OTYv0is/eyOeUaCgE0VjUvSFVnQJCbRZCWwmUgBEc9u7SM2q8GRbPdyy
3xg6GinLyp1+/QUfBwY/PajYwjNC35x9ij6K211rdkn3/VB25eKVjWW8swYZfvOy
7usY1zw9aYOtNpDJn5Zm11re7gFddmDemxv6+GZZKOR8BN68Ivkig1k/CwPVBxiM
ve/+9QheTjU67Oyvptx4kqzZ1/4cRnxdsYVhwStdWWupAqVuM1PEzpCa7bu+pFpM
C/p1IWcoXtUIK3sFGhYxuYnEaTNkw272VNTCcL8TsiBihOioVvGSUmjeg/LIDnXA
gwZ4hQQW50r+4yI4C2MvBenSFoTr6y9+m7Zbq6muTQpTM1EGl7HMuMYgYSv3Qlvh
7txmOV246nkF3/2UUBR5YzIZLjJtm5BzDhhqqbH6Z4EkHsye13F2hl6/Z9dppkBR
uwT3ZQBZbMtNzYoT/daR02UssMe5aUY8ggWAnmTDsJychu1eDr0MPsfX07Xxg0Cb
6xEH2gQJb3rk6Cvrme4waaeQJnS8zj7xIKaueONmADz6V4bozGSpmbLbxTykqPbZ
r/oZji1V449l3kS+RyC72LbMvA2XLPlNiVGk+x+qzuIahj8Us4cDdhN2SU/iO3MN
oKofkEC+I4UZVOQCPQHdUNCZUqbmynUaY6kUVrUqm9bY5l6QLvFqTHVTqCK6qhG5
YJyFDbl6LzxdVaqO+FYaqjGveNyyPh+CBPq33vxnYcBjX7dAsDFccNkkxC9039gU
8to795qXemHL2ipqz31uP61ZEjFYc0IS1HsPtbTRrm7gU9Gk7ZJYfm4eJlJCsb94
JF90QKz0wKu2TSuKj7XtewAaZUpGQWlLolcpPvP7wpJiEZXdutK60dzmQCsm5rOS
qOH2gDkLnb7H3+AFIioFK4Z+YLcVVtQ90mplbfEMTgko8xkHSrfoh9A249k5M9yY
PSN2zlnxBBN3s1t1DbljS9tFmB3C8bri3Lz3hYhcbzrU4Ai80Fo+NghxQp5wTvf2
LwnnB6haYg9OjbagRWpQ5xyCTDRDVNcjOvTwpZrgIQ66H6AR9JEcQpjgri5Gp8iB
Z0XwEM7gV5N/F44JJEUczPHTYpbJDJXl0Y1azorJkapbDSHT6QI/cw50FSNW/T9L
udr5yawdKS4nMPTiIuScPBjCc/1ngQk46JV93QaqFSObMWe6OYgz9gSIhmahS3sf
EkKOwZ/+QG7TgcPSUVt95/SYAERynCOy/u3TkBMgbeU6UzqUvifTSBzF7qSCXo1p
uuI0uo9Y2XaOHWS3uiRR/Rphj9yJl1jOSjYqRPr/Ox550dRCGSZ3Jpy33XVFr4N6
N2Mm2/6vtIxSNmFWUXSNin782N8TwnXzKD2RdJYJr4ozkynIakViZmmqufY1KtrP
n1x8/wVWXO8nEb0metIDxujkqccN7NcK3MLsDnl/TOcXsCzKpXBhH3PJkk5U6OUv
M6TbqDK4p61MaL2TLmJK9C58mJboiVM+nGzSooxfqW6bQ/PM27Wo+9rd39R5tdXK
RGI1nJgkOKfwF3CMlZTMOFerGnDRMvzWhQMj8KKGMJgXakWu+3ycE13DqFTbP47a
RqnFVFYrp4neaI3mwYohacjxt028UmYIy1aKL/H1eo/+26c/6ds7sH1XwiWkORr8
i5/tZkXOI3EyX0otpmgr8Q675/fh3SN5MgXGjc/U8716JkNePRMQ5uA5N9RAElXG
GZNOmydKEFPEcFoKZZ1dFrO9M8//hwzte1EYyZh2lntIxk6SBk+/hnHqilr+dx/T
qPi9OmnJypm4JuXqkfxEckzVpTAT6JZnR4kqq3ZAFzNpCd2RUH7mo9WzfuY9JHNh
cbC8+HXBIsZ70rBie3Dkg2bgeYYwkezcgerVkENwuHYmGAdqifXt+7RrvlnR65Dm
XrsDlKLbprmM5ikgWTqy7HulSSgAw1rOuwiLpbUeDzGK3GvDlGgliACXxtEAnNRh
+nAuO2cHw7SAlMUePDHhtBs7r4GH5zDnnG1wH+AbZm6C7m0+kmM0Yz6E3Z2B13dc
e3vO0f1mYif1bbwsdhbZWx/+8mvSCJ9n2SHRaMRlHYwJAsfbHKyAtStCaDm8Ef+b
l5FTXGi+d37Ltj/CJLyvbZraZTg9Z4QXSb66ZUaV8RUBBj8G0ixZ7Wt2biIGPPJM
vG0XrBhBSAQeYD4mjNxy8RMwhtOvs3w9o9FB3zXQiUcE2x+Dl339deRG2SAolHj3
nelUIrMg6eVXvoxRC8RucfUEKrIEegnesm2IRXmPEhb2uV9awuB4ID01gwpB7+8I
6ZtSlXKeZDrngjImyr3A/ap2x8rtmzle4P++Tz1TPvp42743LVOeczdR7CGeZLha
laztRAIQvz9GWN4VUYjfTYRJIdvhsyX3ahft7qeFBB7i0My41uOGQC19eu/FZ7cS
VsSmPtLogGTVXuQB9Xq214WfXISmRtMTaDjQDYEcZxSVx0JcmUZ/rE90PAUFdDi1
EETE3yeTxw/5qXEut1Yk+dQlRtHak6+ZBcpBkGT+z2CTfkX/FSEpRnwNkkMFqO4J
X3obB01n04HS6h+5wz4I0CJmklZOH7mqLnU9DeuzS8mWwVlZgFOzHeUc+h/UthZl
vDRr1u3ydzmr/DppsYYgtU0s6Crn41Xkvw3I50e1AE4OqTQgGu9Lz9xmAdxdD1bB
Bi924+erlHCVqAW2CZHPfEkX5KN4Ssp/DJw+Sfsh27ypeiDlJoSb+0RNwxuMP+wz
QWG/vwqlV9ucn9Clh3nrnldcqbphI61zUXHzjNRm3sB6PaKrC5S622GVX9XbT+R9
tZ9NqM3BsHsXOW7UhAn4AQVikpedIX7hRSmLkFjKZ0LsFCCm+u8RxgkXY7WIK6HU
0DxL5rO2PLZzrb+fiH7ARoUnyAM+7y4hAF7xzlJ6iamDG1+iDdPmMtGfFZU4n4kR
UR/aI5erOZ/dwoJ6Yg3LkLZT3LqgF0NT0Lx+4+yIE/75Dtt3ri0tCURq4cMqqQNk
tnaadCTyfnuelIAUow0UQHnAz2rmgyZqQ05gYB8ik1Tc/Ke69094TVMLow1qFzB8
O9rYCdrWGn9d8rDe1qZRutV8uUqleiEtD5TOWKJQJP7v/EwDXZ8mUWKRIPMragM3
UpvAXeFOjuQyKEf5fKKHPsqDvHNHyHQVU4ZWgtLzITiRzutJ9y7s74UtlnvyUNB5
gN8HvhqK7rUtoQZyDLJL4aH0uW1OwuFWUJdrVDQAPR/pdlCwWqSoQvTqtMiySWcB
1Pg130KSeKYl12Kw71eicYbDW5R8+a1c8Ndcrv2+P1pgk6GHxm0NjVCZ5N6wmoPZ
rudWjlacRd7ZKT1aXVLvRTZl2V/U5obsL7R1jmSz/GZ0bDgeTiCO760R76IXdP/9
7cutFjghQzk9vYseyR582gv4d+xwduMridzVYnKnHI8JaSoJp8E8t/aLnqDm1rxj
vZDwQm+ep4qO1CD1hz5kN+7ISa5KQA6fCa7urWiJdFBv+m2dX8I4ebwW1UlAXgFm
8oi4XP5otpbQyWv2ZlrKo2AuvaTYfrCCQPM1xPca8t5VYaXJNMbJwFd7pzMqGJV7
vOFSRqk4OqpDGwpkMfoHqtrnZycc2udC6CJuDjHW7Pyd2oRjzlxzq4FhV2ZvKAm9
TNzmjsuHjN+A1j+Kz05R0WpCjav9AcO714eSk2zpiDI0AM7itj8tsmSkT9VbWmZQ
pQh0WECACJDmzzxAyU4IAUEYrlXOVx2XmG2QT1gG95uEUsvUCy84Sg7/XO9ohTiX
Hfdrj+JIkKXsrZWLpKsoVCtEwBKbvUTVdyf/8d7U/dSClS/CprGpbF6vErhXg18J
yD3ta6dixj/9f9DluHD81tJrV7jbQsxGLuaYOvTlK8AVxIi7cS/r5UsZhrI/ONuY
WlhkdFce517KYSbmkc7w+dEIeMaWrDHa8fBzK0yMJo07Lbj1O64lIKpLOo7p/40L
fzMs4dJhp8VQg3pikXIV4wLnIgdF8OAZC4nphuUC8EzRMQQzQTb46ORIa15/m+7G
Xu9/KtKvE44n0DDtHkGvXCaj3/tUhr8xUYkBiuA+HLXCDjWukQWEJssyNYRs1F7F
A5/SdYyYzYl7QXtFae+AeMJ/Nq0AhFn1cf7yoixVMYL606iD3SPUY4Zmk9jhNnxn
/P5bZ044w7oENIrbWw85lF61Tt6IB3m/HwqXfpdXe6lzVWvD3LkdOlLUiS1qJnJL
ZHOX6GESdU1xr8anC4HD17UJ3nsBcyLmIGP1fPXvHLqSCBrPGw3h5DRjC0z0usVt
jCYxIsZKzc75u+7KU+X/KDdQAqzameuk/PmbFYC41iw6csOS8UGMOCvcVWUBaU0l
lf8ozS1CrgWz7ve79SNsc2TkhFn2JHyBhSqU0S5Uuw4PqHqI+LEG9o9pgpUYQYN+
sNfUWtDMNsW+lySFnuqwIuVEXgBSS2CncOgtJ8VQOJOXWoEkY+PEzgbk2RUqK/bO
s9tV696vbyOavLRVlA2cKh71iRi6u+dkx1vfBb3Q+9hgKHyL3r8+d7SzA/fKcUmk
mOAN9d4QFukhzDLHJ4ix/oKpscOifWDUSh2ZmbMhOXdZDpUHAUu9Khd5AWSMspnU
H+1sCg8vBqqWvo1Hf2rNPgoJSnVuw15+FXK2QKjz+0lG8pXJykU7KRjFuJcFF5tZ
7yeik5NezTHBH89+ymU9oGbGX9w2Z01EjbdOzEQRxLZs9l7SPyMvTzvppN0R4doO
fIc4NkbhGKumuFWB0fUp7tn/BwAgusuOBLY8Aa2yw6YuTGTXW5J2LEN/jo29J6rp
7vmjM56WgXyh1NStzzXX9pT1NRd+GxmUiLJTSjpVF8NdAXR8QUZFXzEF/opU6XO7
UiwKmN5tUA9os6XkBwvyC5gzhJfOq9R3SdhyO6XeJ3DwwfB85uwX8Rg9xxzzn6mV
x9RmPeQs+3iXViMsGfa0IEujtawdNKfZtdLE/ZgxOvbbUT7aWwV/BPJRtFYKjHpl
2pYsaph+3spOt2bl2TDnVoaP6PfZ4mEBkfUvqjlnlqgQCmLXef+PUVsgasJYQSa8
0LRpBW1w59fRtzhaWWgtbwu6G25JMR1cpJYh7zX0dPtg1HHCeHoPUxWFCtyzJsBQ
3sOCP2WhRGZFy/b4rmUERtNZgmMndki07lFB+iNxRLEgzu4pwmHK8/6AqgNvB5C1
OEJNBEepc8nZQqC2M8TozOdwv3RaRdTEMiuw/dLzf7aFXrJS+lffx8C4GNT/vdDb
d9vvYVyiDVptQzv/N59FoQmF/3U9RAywWKnTQzLnEuZhcwHKI6eVLSveeP1CGWat
XTb6sfhCoWFqe84HMaN6nBAzeUoLOipNVEJ0t9YYHsooQ8MBCrzS/YC7kMCe1qDy
Wpa7mr53xmq+ye8hDPSe8aG1qlF0DM4jwbiMkblax3NJ3UuwhLU23QVBQXR7HWMG
ThnF/8pEE9aSfjcRJQV7NpvUcoNKYRfrNG1Oipy7NrB5WKDFt9yd9hknWvzjAnaT
4uvDHiIqjUavM80nOW/YCNuUvVjkDIC8AxwAbCKi2YrB2TN2v2TYZqZdw0WdXxZ1
MG9UyfzdMvj7JqIyuaIwC8+RfdozjV/rMNfhkmvno3K2g2aYQZMUJPP5B/h/kHoA
IfDdprmi03e1Odpblax4kmC3oDVmyKJ4va0WKH8tupQR3WBPdputCDRAKwO5UYNi
97eeKs/CWk/QN5DX1YFVhbi1vTzY3MWLXbRgesmPQFmnR87nbSKG3ihqbNm/Sk1a
PnDxiWdg231mon/G328wKDcWV9Tst/bhuo0GxZQixMtMFTZPe++hDF/3WccMuo10
MZlb0wMRh9sssl1YlkI517q1fv7hVKxtdc9YThDnZw603OX4ZkUugI+0sJRy05oO
DNLXQwHzFx7jksJV9jcK6hzYKpPgdkBe2LoAIZ1P/pcGZKebroAlgtomT06Q7m18
R8Klshw0kKCyNh16Gh/aq01nCr2YRN8DQW6LuXSAQdSY9ZDvCvGlhi3L8lDBD6Pc
mrWMdlwdO+IEIm9IkiG4/kjlYZYfEV/gSyFwde9n6MsVQ0/WczV34lbd/tax+pr6
MvKMMn68GZKr792vWMpyqb1VHTvHdfjcpBFrzAz/WTQB9ISyCr5PtjoIAc+ApGrQ
4Gr/2B/3BCusf0wO0wPwcdFi3zEc0rvbtbQGjsIwmBdo+JfdLYJc9kYXm1TzK0hm
BCYK+bdDMbEU84lWAfO8ZfuPxJ4+xr8OFr/lbMlmyw0EIdFJiVjWXWfuZcUlxKVk
Nx/dy/kwL7oCfm0gpYzwBZ9Eqk8JoGnOF8DNE9HuVZCVgSSRj+35+bQXYTPO8LAg
TMVU3hLK1AOR77TikAc1084QVcXQwcHCwBkpV/i7WA7NhYLsNW9k8VuIsAL7Xgux
SGADkYoTVhmfnOPD143NTvSr58Sn4DVrLDkKeIE9/fvgNPfnf6VUChs8PqOXtg9D
q62hHQiHBzSd22xlJHtFqX3m7CE3JRwfIdDB4HcI89xdBsO3j15gat2Utyq5Hs7E
nGwOYCGtZ2a+i68lliadPjulx6DBxMQjZuw5xDnwQFhB4o+daPHMEF5bKaSOHfZi
6Uw81dyulxLlMTaLojozgltdcn2nhz5M8uYxMtsljJKP+zMrF1GE5IP50BsM8o/s
cysUSFFLzi5UMWYCqMYcpHBejavxH1LBTGUWdhbSrpo6LeBri/nnh1+8UrN8PAFJ
fy41B4VE0J5jy3DtKBYvdlPByY40MylM/x/1IXAH+7yC1jiza/6iTd5+NTfCUhpl
/vj59eVXsEJaV2tLt9vGiDMEma94qyXtrBpUJZXOCGuW8YxS9NHHYoTVvhstSi0A
BIRBQulYWUkQPIwj5xmgAv0dqkFhY4DCnfLKvasrx6LSuG5lW62+Gd0TD/l8mpf/
OhBOtsY78vnz2fJ20GMcEI0LDWeUKj/l9TrW1jThtB7QOJLaGZBLdLTaQJPnJ8Lu
Bo+5/8uvkBqvevFHAGvmIXCvKp27K2M2A37oQILHKPdA14INZxDXZFQVXZ5xAHky
wUfKh9CwfeEpQ2idFh6re0Aw49r8MvchL4Zv+oNN7NkmjWJ02hkPaSljTZP6aJVM
mDmgZCfn1QpKLiyPMMmaDPbfvfxhiFCN+YxANi+Q4NcACNGoWbhwODmYYx2lzL4e
oFFbYcGqX2QSkDCpmWcUzgeo8IhMfcSfWmDIdWtV+38g7vHgzm0SJ2ly8MZno1Sd
i4EODQULZR4msInkeJba8MqWkMN6rXk6j1cU2gQlGnrC9AGL3mwBiH/bCv8LwttB
t53Y0ibGkTeQnXg1TJqNO5QQ/VYpnOjicT/4pc/QAy4giWB+PZWM952ekxx/JQLQ
BmASmhX7g5xm/tJwhLm3G3bHiLMY6yyG+UK6rWDhQBSJ4P0fBHOcwq5M7rEobSI3
C1mzhT0gO7Kzg5TOJ11ReawP+fB9haL5OsgdRXzQPtI+ig/1exU/MF7FxK+zyN2h
tFrZjK6Dmm8Skka/A32aRgS37N0wvbHt1cMUf+WSpooZVa7RKoDLCE7+i4r3G/in
G9n5cyw5l9+hMSf3d822iyHodk6Q+1DEArq5QjjHGePzOErBNW+YqA4TMgWMQ8mk
b5kwt6A5HivvjRtoQHZ/EY/acspAyD8r498lz40T0yttDja2dkkRHtpCC5ZLG9Mz
PpHYM3PTKsZO1rabZnsKFUC/j7udCrsZOahnpA4NkQQT/E2RWx4NRYKLZU62On5G
a95uqQ0UsQNb0TW84gVzow5+DywDkHsAS1q2hryrv0HZCQ7kMdqrBtyV420tFbMd
cgfrQcaLCTn/RIDSh/LPrkCbqAK1EgUaApn/HflkXjRq3cL5cfmoUp2YwYPqMrT1
Z6oxBE/gKwM6IGb+/ka8Zc7U95zmjdPjAOz4jsu7tUYYULGzdgvBhciK18x/TGer
OPd3mLEnOa4261VPGtNpX48DUgIBioZ3L3j901XWxyMlGlaz3xzzisox2DwfoV61
0gO+5oChxM3ahwwR4NdDnYnGV/1vfukTskIuMjWNip9ktyOAOtzVCnHYC0koAqfV
I+JIuWaSB9OlOK34RhVIBSo1l1/D8o32hPORWIMaiqgdIoV3HBIW9nY1h68CBW3Y
78sej7HYS19tKH+oHFSrEx1HMIOCGDPz347rh9ltjyfhaliUAyhkaA7QNEsH3HcN
ANdxzgg6qFO4ikrDVtzEzSnUSWYxa00fAgCBalbz2luhaWhImwQg/4xfMC8o5aBx
0ykitUKDc2hLcWL/K509rDBRRzw8uKbhqQ0tXUhwE14ZSdpZREMYB5zIWAeEl3yS
9dJ6WfzYwMD8bgAdVMuFunmvWq6W/arCuRSk6HC8UuSfAt5i9g2STA2kbtsKUE9G
GddSshLVLbkRs6o5aoPVi/iKSmWqBDIRkCU9vUC2vapk3eE+w9nGPHGsnq0PcBzq
7BsFQxCjSj8EYDoHKAXR8//fsMw2fbDBAdTuhJYwjBmB6L1rBQzi2qhV6YPYmTZU
BMqBjpSSIUhwd7ANPnRDXfzCX1ZylqAh3CkIecieisq4Y/E7yparr9wqzGR5fYsz
EdUXt4fAD2oFjv8/giM3DSvjUxQQaGM9vFOAtGg8LeSP1xnou++3wMwbS1Ge2vKH
mm+1AYQDl/1+GSj7nrzmb0719l+BsQSvnzKPrqjrN+Arz9/dmQOk8MnLsjDWUVMH
slJKw0a7DnrBZ27qv7iNA+f6FLF4sKT9ctmEJW1mcxHdFKA0XoMTO3eJdts2qOnF
nCuOZMDoJu7vXaCZ3SdfVj0TVyJS/eW39ATT/qxTn3N2uw5DZ6KloabXGuydSXjk
Sn5D+jYQmqo2yKZl7DK2wmKQSuPteUvBpVQrHJmJPghmKhHpHgFBVZk0HGjcsddy
THlu5NUeFotWvcYVYdpUlqhV0ivtI3iEIsDmB9q7bV8yHPgUHC20vomQHSV4DW7h
4DMDaoIIlUHnYIJCxtxPZKVGfV4eFdDwphc7JUrUyYP6cB5WtHMGpdyUTI8lFrz8
7wpKK6Bl3kkQj9fjhOXN2+IN/Y7PPasgoT7mwlbQnRq9rYMG0mi1EyCNhveVoH4H
i6181hP83rJvbn8GAeTYLfN35ZqlDAG7FVS/enXstjH2+opu7Q534vD773UCFWIE
KCkogvelOfCRux+4ZS9F0CvaD1CLfAGjd0wGC2E+3wsFBxA0h4wnAfZNgK7w1BLq
RZq2l41fOZe9bgpsABMdJTkZtIklNNHUUBO2lfIZpDknx7z/4SF63o5h95GVRKdW
Mj3AkGKOZ8oIQLnVt1NfRKaQK0cgqyYx3pLu9fCwtwrJyonJJSKdOBbcLgE7Jwi9
2Z1fAi3c/zR6U4hyn821/rbVRjqTFFPNfcxqXvLhjRzYAm/KxO9ogoAMsVsItFrg
jAEnpLGHuyyEswNU20oZb0je+LPLECSyFYH4lIk66amGRmTMuFz/FUXdwEby+vaV
Bjmgxo7LFMeP9kVJdv6+I5kRk9CVOMTf034ED2WdLH+B63Xy0z5rHmbjq2Oset+h
dl8uyf+t1keNXukLwbFBech6DpKGv2NHjuBUh45q0DiA9/verENCZY8PSxab41pK
Ya6NZv9lVYzvV15JNujvT1nncK9nWgJFqQBxn2iNDSssNdiYOIXCHQGcINS8jly6
mmoBiW+ifegibW9a9JcBtdVpxpXuBinlYH//iwduN1UGW291NXd6cOjMkXTK/ynW
QGi5uEgF6MELjanMWSxdE/K0Dcv/84Nf/dDOuQX7m6nWqLgYpEMA4vPuRBBMZD0r
BdRXyQBcOXL/POCMoW2XjGrm4etQy5jttV5B6f0gC98LDP9Zx3aIJ8zoyGYCcEZP
85qBU2nUg/Q5m1oPXdeI3uFm6ijyvJQ8NCRf/LNhRxVv6BjhcOcFZUyVdq7BWp2v
2MBbvHD2eeTbcxZ2ZHzsRCGkYY+6ZJlo49wOewpAn8GmdusgjP/4G3/aMv3Am9Aj
D5xu3bKttPk64ESrhQ2xzcl3JOik+MW5swsgOZ7nACOrTiJgV6pn5FnwUhnzKwJX
JqoRbDZ+GaMTxTcQwqQEOnDsrQM/BD7ZqF/Ja7erxoWMPLN3thU5q5VVI24MimAP
ATbeUXfsHp6ELQPM0WhxP5x1JwVWyG7fI54AV5st12QmATP5oos3+PyL008sAIWe
/VKGFBhzFMIOfpif2fb3A8RRd0734xS31bAMYSWZytdcONPQH1u5zeUtjdix1ne5
D+wtNjExKt5aSA/1Q7cbQSD8AfRKehW7ICjK7saUCp4nYANpg6RAtyNgIxwdXO2A
dmGDpUC9GQ8rD812pOIFLVbpK6XiVAP3GB7xpHVMrBuC/LETIqd8/0fjVPaP1T4G
sGGaEMjvS0jy+ox5ifG+9dqHNLrUNrnId/FmxORZ1GxKo3uQmBEQHjcEKdFVSCNw
rfiiSzzdXuGts/JTv4EcBVDEk3mKFMap0RQ6bMCcGXyAngpPGBOq2vCBYeIrZMnk
0GZblYSU+EsjAiY0aAZGqRaTJ181p8X+QNyDzb74JRDfhwVdgBzED9aX0Xj3Vvy3
bEsf9g5szFsPVOA21mP7RIPIhoaEd5D9Q9suMB4wRr5l1x+SUDQ2yjAaKBEUDZgd
/C3x8FxvttlkA+eLi7F3QDX24Anf58Q7yH6yNnioV7S8KJd0SQ4UUjW5PLjYlezu
K6HBdfLeJQOM020RKSqhVWe7K0YDoNfmY4xFn8Xz0MimJyVgYEwgElLn9ycJpivC
SdAt2upxa+YX0QERy1OTPZY4/EZ9LGaN9sY4Fi2S1r7epOk89VEdxpKXyqiQLabb
abfSIvkz9yf6FPWTth7GQLJ8IuC1b1TqAWPTiq1DczxlGQfoYmm4lbfyb1o/qtdo
1crsbLSfKKoDg5My85X00PC7ZMs1l7I2Jv28IA8UtEyVIQo2OPYCUtQ4vnQlO7Y1
5TwJuYmqYIGVThweCPUjUuyx5hxqexHVdGgPuM+txfmWTS0WrUi4AXGzpvbGUPpJ
IHZ178jC4h6l5XEOKnGJb6M0RWp8wm/GNPn39lXaARl0/x8JobGFYy4mVwYczPWm
CH/roHea8acJ+iUrUqyBaYnivyFXAF8vza9fmK5sk6ywJbgePZPGY3DT3QKvq8wF
+z5wibioEwkoKmz9GOomcV5kn80W7g+9Zd2XcBBg3+VNNna6oEL+fW8OEeHK+LZ+
ScNejXyAgW52ISc2PsjOAmE2I6xal5lkPrIX9wgZWkRJauxQ7rAQ4qoEsh/i/SvI
AEicOKdlI9FmmrbbrI6C8gdHsscPKw2lztOL50FgW4nEtJ4R3SHnuTyUCC+QbsQi
TF/tFofshRsIoAHP99SgdYErM5xLQUByyz5EXyvD4UjrYAFF2ViCo6/sEr1wfmyH
q82yrX8YccJ0P5E9PyyvFJm0jISUmyJfH0o3XW7975HGfAZvNKrddtZJw8eZTh7s
aXyxKH11mH0G/aq5c/9MOlQL1NynJhfQCnky50o6LgxdX3weZVsonL5vuL9cDc7w
5fkh4WpIOxAtR7gt1cVVCxoIBmTHwXW9sE9IuSzvNbtAAaCf48LcrMJ3XGVQWCZt
XW+qnn/JR6Pe45yLCE3SG0WusUwai5+8EoKPfMFaFl9IDWzqn4xl9IhpeFO06kCy
UJPfHXV/W8IUb89ZGxwD2+lxxwd7UZK2zLW4ZZ7x1DbfLRkrsSNmzC+DHTOzkt81
XYfSTWM9mkCKD3NeFFNohUdO/9ONbhRS0xqiCMBMdUJNITRECZQtAbRIVl7NvyqN
4ZY/GFFv4rR4N6elhjU7SjMBhVRVFqZet7WXAOAthoi80zV2kxlu4CEhCAkjbDfh
KGOfifsj+sqfc3ZUdgnJK6CjRzV1EhxoyU2zvJXKY3RaKaqMYtNGnMR6jDAiDabj
sbwdn5+wQGqXEJ9fu+/vrh0jVELYvAb8zWBPtucVVylJWHXvMDPuldkYeLA+fcvv
KeHqmsAmNMGu8XlC8mQIbuPI1UKfrSGLN/e0PWKti8bfqCdcUr8bQIINaruJY6eP
bzOsOnNhsSYq6yWrRJzzxijLeFiHupBXvhbGeaI2EbqKI5G/0g8YrVncKmLDiloq
zWnQuslM2kIOT8U3URUZGNazcqdl5su1wD6DpUfGBeb1ao8xOcY/ElC9AF9Fb74E
brqKhmyTwT1Fj3H+BwbA5g9fA30trL3i/OWMIG6AtPka8fMg38xipHOWA7KpKbmQ
76zZun0o/l4T2/ELYZpNGQ0510dkve91TSTTB5DxmSGlpByLbMZ+kHCFoOmwMmGv
EvsCopj8LC02Ky1vNSMhi8gw6Olw5a/3OW79ff35IC/HJXzKfu0g1yX2L0z181U3
AHbUGMdpXr8pTiBxv8qopRIas/VVLlk5p5fGbzmxD0V+HE+R/3MvjmcPonWxX1Lh
X+dYGPBtLbRNC6/HqmdiyZcHc2cWeXdpkMCQefdiTn1ikIT88CDgF6WLg5/Djvy0
+jrA9RjWaOExQ6mv0PFJK3NLjJ3JoRqZRc7DI7/4pwvJJKej1h8RFjqDyHI00Jt2
t3DWirYJCBv30e9Ykh4ElwxDjuY9MajwzMFfD/2vh3exHsv9ekGWybmWyzGygexx
AF+KaQYu/1mEHQm6kNyWKTyBCemyHDbZyYUcsv0nQ6EsDUacrZujOJjbjH57SFBR
6iBOo29tWi7wLm40TI96HgYHBVIYyosI6YHWVG5ETt6l0J81FI//RO9jjQORDXbN
DKQlVFGi8VYuOjIL1t5ZZ8ZeiBMQ6dte1qBo9I5Dao7UE0cNA1f7gVayIL1kAgSv
lOGhPDLyXoxKptFJ/tpciS2Nc0vIGYybLQ5xHpjOH4n2gO0nHPQUBmaBpPiqU2yu
htAHtjF9TrDX2BJl1AXrWfNEia/47PDSARipeIXwBBZyEmB8N23WP+5wRlqO4T8d
bRKdyORkdnjlPu56t1q4rT6aD0O7uzjHYSqfVYyIZ7qdTmPHxM2NYx8OiYYRga/c
9sWbKBJeFJkrCAVXpIaCVUVl72rnQ65gFKVpNjTa+AC0Rd2oVG/YqnPzvvO1hGkX
o3UiLp4QEXhFnFszs26dL+6hQL6BNzHOrYWAcZCXanHxWDkb0wyBm1n3rEf7Uaoh
Wjyffsl6LcpJA6dmjYVQsniN7IqRYaId5K/Wjwqq8mz+35DD7GBm5cA9VRn1Mtbx
jANGNFA9sg9q+61Jo5EZibZes4xFv3xCd9gk4Zvm1UQ/krZjzV346NVQkZHUVmyd
8EGKDUiTbOPBtyT2aO8LGsk/kZFabsr6+ry3+uihE+f2RawUsGa45bqQysaSpW4S
HERksTrsXapIIZDEShf61LsdVHnuHG5kCNbZn5S6+cqvrY5JDAxSl7aV93wYF0W+
ZbkZ9Rb9xFB4/HQqdGXip7b5Wx159bMf7IwtfNDOxIp7FvjPIrdYIbcDPrd4IXf3
Sp0V+iSae1CEFQT7YeZJSASVg4GUR8mNrPiruxbG9D04M9a5CeY4zRtoCazGTeuP
XTSCM/fFSOnWIqFm/i344WxhiihbGn/IrwNAJWxLVPdAP8fSNeuLc10TJty2stW8
JrxAg4AxR89tnT4Vy4kusIaqMc3xIZXROpGfvYu5KQiCI7p7qXOx4X/NOzBkQCPh
psf1h1ai46dGneydgp67+t2Vdo1VBDE8QTv0liNbaeLR407D2jVg1UG2F6b2orEg
5NL3R13Cph2MW6vpp901FO6WQx/u+nVyevZRQjIxvzgR1tmW+VFkplp4rY52xQAY
zQEagcdJFamOU/EJGaipp5qIo5qI/9YohOwSRjXx9XNcE2W85r3fuUyCvshUQTjS
ZlMh1Wbe8EzQrbAf0yIj1EYA6V4URA+BPGicU4hTqF4krLncXUk1SaNzLgK6zjyl
unNoMMGA+HP46EdrZWqMiqU2sT+nnxl/yDsXWjJ0TURCOkFF3HZR67pKb7HhHaNb
ceLC8cwe4w1VZGrEDZEqi4CtS2QebPau4k5AuwSa2Jl89woaC3ZRtG1z0ExvU/Rb
Da8EBtyjEn8/BPBONbSknR2Evw0W+A31ynYFiUBsqykOQa38S25jsO64CI7IBgwI
MKrGi4XaR12hyuw7Qnj1hTijhilAVSKsvZh652irD0blOyCvB6yLUodoWjx1XE+9
MByDjDGgv9yfTmxFTYQscK9kOFrErVLR3M7UhGtidTtYLf2pTezY2k1jU6vzmdCx
0rYwSFZ1/cce7+7SFaQ53dHb/pfivSgy8WrToXgsQTNaTrGv3xq16bDuT+Tobmbe
Ivii9wZNvoHCRToI1p+vIwrYXTL7jjMFrLgoVvofULMuhSwgMdrVCln0ZfqgdLJ7
HSr3xokzFqnSC5lSixkoa5ugK2NIqhLqUe8EctQrcugcd0zw3wEHQBbkm105ZCL2
wTWPjiuQ3PIoWy4tw/iaupjp3nGR6puqPEb2pPxeaakJIiCn1K9zoZTDtVjp3qvx
T3xPKolxEaacuvt1sGDthibJhrJ5yv2JGvbBeEVHqp7Vd9x6DiZqKelmEzNVIJEW
5PffeZW42oKKsPS2FMBBOK6y/FExLjACXEWpJ+T0rij+E31C2a01iY2b/TACvD6t
iYsGEZNhZCRa8oWRAFJ3VDZl6hB6v0EwZQnmKLRz/RMCLqUgpk1WtQ00dAJOg6kC
x3HNa0voqRLTBUKW/9RlGXd1LnQahscN7qjjiYEvRrqpL+WaT72GH6WvCcO8jPMw
eB+snNcuxgOZaGh8aIdCiC0zAQO0U5EKbW10WBdjbabP5SsaT4A/9qrzdWqoJK+h
ze4iWwV5CMFR9sgrtnW9wPMIm5jOgw+Cls8Q8BeFrpFLWcAYaqdHLYx2tZPetR73
+9MVMf8ZAJkN/iXubDYDlYMToNxhZjdu0dLNPyX2vIO/wFq2TAB5az5wGeYXwbpr
2W2yO1sM54zYn4G0kJp28+aFta8EIuvodMEMDisYEYkeHlBvOn9dG0MA7w53oExf
+eKFbu44WviHXVDRCvy2ku96OdYmPYcN8s8lRgSPHniWusHbXS96jlxgKj6LGCve
xqysQp5z8Tp5N+eh8dm06xPEbUE7gHVKCH+44iqrvwGuVICjkOtw/k8HGPAYj+wa
6FBOe6ItM3mkReyXM+slT9Hppa+FPK9X3yAkMX7pso7//+S8y7HrW2OluZ7AE+YV
FpDPHmR80WG9NYDVIuqhMg80ZXm356zsJljsiPZoJ35GsOUpisUZ8em1tIOhDLSH
4nZh63gxhIsPqlpw1/4iQXBJ7lxNEtJfum6zPDz/N0LoKeGaSdZXsHACGNeOJGoT
j7kWLZSBkGHpp07oL/Kcl976NotTFCrbkUkU3MSz8vQUg9YwyLnKzPIG9V46CZFu
wSew1nvSeFknugO0T/PEJyxdWN7nUPtZ2HHGfN32Nhi6xwi9milJIDrbkEHCSk2Z
1BzrwNhsyR0GujyffWnXrCnrk7oOe6fTJWCCKny+7o4j3/N+6hJPVHQuZDB5LzDC
luidXMSV/1FEfmKepCqvMrUapvljeei6N+8ux85eEkDWpKEGUaXvi73+uSZY2NV0
DVh16ofLJtmSGKgc+E8oleAmxPDNrPuMnF2Mi6S3V/EWjwR0xqKwMNP7nha6Urdp
rm7WKXBBy+gP1GIqSxFXTq1EOo5H7KlWWY0jae0HH4hA6KWPBs/5j9Q34HEf8nE3
GkX6S3DmRDUMWLHgw5ExlCyNrEtsK+qnoZWlTDQrbXhrHttMsIKX8tsQ61JKlD0L
HX+7rwa5nMCDHsbh6cZShsPkQAp4N5IAtwSpt/kcEHpUwpQepCgw/Lt9Qqd+G/Zx
f1lsymOQWwu38qsYOJL4dMHpDi0y0j6Fk5xTyh0Cdtv2cB4CJThQ6lmNa9Ua2bpM
bMJaMkgFYmI8D6hwlaWHogY9buhR62gN4GTFnSeSkpnKuuNJWmN/vUA4LhwjOMZO
sWMzbZkDVrJCK5/sg+P89mXeO4TZjsZ+pH3PgX1VVjiHhJCCeVJbG1XliRMFtI4c
nLi3QAkmpSvcoV0gOfNglIVhETsiGXGS8xkADNXyMAwCwS6SJWMQepcEBigvEoy3
jUqkdPjkIP6r/PNYKT18/FNUt/PA6wqm+WJOGVPrR3aqCo+wQT/gVE+7KAyL0oeV
6lHLC4MdJpySAlhM9MB9VxR3UBAMh2zKVd/KyYYf+jl33cPmZvuKYmrsMmR6SrfO
6c9p73VEnOXtnaGj51u+qhx1jBGInv3hLZeBvTlIMHmscMhuYXxikIDbRd1lGouo
Wa0f8mRELS5LpDKYUfCsQ87/skA9HQ0OWU8QTsWRkor05Klce5W51DXFsbsdqxlp
Tem+Et8XaJs4KWPsvAqtWvAqCjOdfDblAgAEAwr4VwcIwkl/qnvtfY2Ld0ANBS/T
+8oG1uveIbGsF2j48/gi2JVM6WkrLc1Hnd60WsOzs8gAHudZvwpaC+rTkHjcGoNZ
+4/z/9aPu+AxnkoaQMrf0Nxr2LsheAqnwnzKPngl9qDS5DSW6yIohTYwUhaP6p7L
BKYAt/MJU6a4IX/jM8jj2q2rldrlsjsqWJmsYsMN9fvyWu/tmW480yrObiblNTQI
G7/Co/KIfeFAjuW9Ybcnq0/rEACGeHgXkENmr+QeDxjsNZBoZAHrB+DiRpld2bDe
OVuIweLDl+c//ESzduvgbsxTBJrZx1R68anfQe+LAXzKRaR0mhXpBTM3C/gwPVbj
+3nsiyU/Q5tvIvwBqKwT6m32l3nfOZ4TTOoKd6nnMTHVL7EbW7O0oe7+05P5p/JU
3oBO98QFH7QoJpYbBkdXoDfk9Hq5JhTAZTvFqGcRB7HqmFhDoxccGC2Nx3jhoSTQ
6ERtMOwCITSNjoJrTEz1f9OB7ModVYSdgizp3pG1KcMepH+np1yti0eXiMJrJGFQ
k9N7RU6JmMwDLbEkge1xWOmNP46Z/xoAx8gWWpPQ6B90FBi8hYW3oHlOInjh0aX2
oRyhUvMP8k8+Uj69/LcC9E7PGyszU2J69HFQ3cPvAZ0p8c9rq2FBk9tgbafbNVb9
j7G+xTGs4Oaz9hM5lYOlV5m0uoz9NiYhryLaZowYs0xpBgjiLPNQSeCVzplq4/5W
ziaz8MjHIP88khVzN4M0TjB/2A3S3OSFXTWncFOeTjcUugpDo2OCzjNuLWmh47gK
yR5oVqc5InYt4wSYQNwKYY1uaQAFb1VhcWt4JQWxST1Yz+ZXCsQLEw/341X9ppLj
NOzclxiGB4PUEx5aaZVxfOE4IEdbrsunyhXZqR0bRJzPBzzeooLoJFyX9D1UEh26
LSe4k7052KUsGcyq0AHANASPZWiJ7R3Phhj1aoWpJmlM7ECQ7znu/aM+1Y8dqYc1
YBJzbJvSnAedMADf87mdEI7mZuu5glRMjTdJC1I7p2wUsOLmPgQMOi+dR+Sl6K8o
Q9tBhA/RNNapW3whV8OFRLkiAoDB9ymOLeCNeojHQ6pLygje7l7Ca3tNsRoXYTwY
4W/L5HkLdA0HvR7xh4sTfFCMOzXx7FBLwWoGr8dNVF7jhzYYtxnCvE6IcD36x8bT
g66bmFYn/AYGPYszcU2gd9szAXIOAWHYh5ElEVnFZlkDuSbOeLBQD0kXmfMOEAQe
qHPVIgEz95At4PTVhgik2hMel0hrc246xfgQFemcCsirYCTM9NdDtkXcJNjnklY9
wpLQhoxrPGwlcX15QAD1NIyqGFM2QF1WomoPoRhYUu3Ls130uwj7B4C/3Fqx2Grb
+Ldp4ZuBlFNzyDbNYYrCwAGzFRgkN68aeCCfqPgdw33MVjfvSz8O9jkJY9LZ8QbE
mLLjwZLyDlpckUWO+y2JDzlIrUPPfznb0oFgWNEqUbybaJcEVKGNrjwD+DPzd1Ie
qXbDYavADUYh0rpbfYwai78RUnnXCq70172Lo48Q+J1Slk7PqsPt4V+Q27CB1MrC
D/Y6qgXXEzDQt4SuiJcYO0d1vy26E6xxwLT7zpwiyASAj0qLFj7APiWKbzfrtGDX
snWrHa+Gv32rNXVUf8qQrCZxRjPwYHq6ajqFmQkVIAFks5IDC1j0vj9BAI5r698h
bYvsPw4fkRvQH+drriJiGVDtAQoUYr4/u2JMb78CUAxO+fzVzkgIXPZ0oGtITXkJ
DkCCt1GoVSTGhDvBVCtFG93wjIYqk/PoGaUN2P33ACUyz7MhFnnPJo2QHlOyoeA5
t6bjg3wCYTObjrQwdVrr4qPXCUE85HqxOzVRZhRSGPGs4roel7bPnMBdsTVzM9kf
4MxSKGRNE6u/xZqb3oZpyPnp6yKsQlevSkTi/i5VX7yBecmXSlGT40VdsMAofgeo
1MIc87WyXv0N8I7yM/K0GXv8OpEIpSU44+6lS7AlxZj47GyrpTdGraSTNVwIUVKU
ynD5/qgMlt9wouBbdOklEnARqG572DeM19jIyhjVUaNm0W1eEHiX11hIfSiSj5gz
hApli9Q9CL19MR7GrNnPw5Xn06ajijXs+qoH4+pJbB/OJLzQue3AuiZLMHi0fdCN
pFJUdgtAAAxckw8iksITzOixHJ0Vg1GfZnNVqbYgIb/VhnorusQHKBk81B7+frpG
BfNbJOSdmW2bM1Y1/uuZzXdGccYJVdLBENHxvipkw2hYcL9gjpWx+fnnMmzzqJ5V
U1s1wwcMeKEm6Whxn04HBQwj4+GxqTRl4Q6DrEx6N6MAyysJTEwLiHiCuzlIS10b
8ppGYmq/JxKZxTeJ1cS81QI3YtcxCPGvsUA8+PUzH6PRlpUORnWOHP9KDELJXFTd
fVMeDoDhXo6PFO81OcXD8MJg/HV9hPY7ypvsyQZnR7/e+SWmHo4tl6C5USFqeFBZ
MFDANn/8oWFTuOOkLiUFS3n3ilMBiNj7+197EOTz4txVPzmlG+NiiZgX6cMq1M98
CUtHAK4tHQV0oqztJIkZ0yNBwhTAC6FJNZqC06o3LWhp2UJYmanMUwEgWNvPgR5j
XfnUcW4ov6FPdZIc+KRKHtGpCNkCVCZ8upFMfQZwTFEcmrvmD9tlC3bltit4dU7k
/jh9A3RXILDJLPTuZT7GYzEB1yegD21wvWVpBk6CULPdBXkpu6hp7SA4PvdCv7f3
6PRoa2lEPO+CL5EWWWglCKoOOvMVaipI/Dh6p+xF+275YVdMmq1CgAdTBzfrmMGH
gxOvb6LIjmdwQJcsaOUpfP3f0fx2J0ZgOXiGVYBATQpLQRlUCR6/DVkZEoai45I0
dW2HgBRqc/qD3cA7MtN3QLIIbDwzGYVf/8trJlOwPCDWEPhfZwXjO0GUYDX6A70e
5Wc7jJBu2GfZGsxfVLnQpHy49+oXmFcFfpWcHd389jDyU9LR18YNi6C+sSE0ZlcC
vsKKptz3yd0zVatUPF5nDlleZONlgbMhcbChjcx1vmUnDZT1EuMdX91eO897lONH
d4cDQsNOYprAEWWhlDDWUdqvCnj6FRBmBPTUbf7ZOoGkvrIYSypX5acsYkXOhWmn
wph1i9LV+CsuVNTVC36/65qCKEGEC69KzLc/yWZLRD22w2lUpcZwUcepKuqq5xGO
/5enPIbxHxe16NKizgrGo5UCYEur12+v9v5rwInPva/J/BnjqeePOuxoYsprzg+3
ZqKIcXZmUWTpyemkQs3q7iusiPVCdffffofZ7xORL8BTz1P6GuTfn1KI84xykYmU
/Ecl/ErUSu2+Be+7OawqpwgbEM9n1K3MaiEIFc0BWk1MGHR8s9zLO6JWXCVC6Fwm
+ZPeF7Vu0Em8f2nodsqVZWqrf0wp/cphqTRb4Hx23FVAYrVbqVuNWVJPzBoyRvRa
y08vtC6M8r37tXSeKzghHSpIaASQmLrF8p6p1SWtnrbFqn0ohBYTNq+U/PTClCSD
qXAhd0LSBeP9T6iiMg7ZLXFR5takLBa38lnZhmwdNIYJGMxyoa3T7STqZb+vfOpT
4CYO0sbuf4wFEJXET+ivGJz1ga4fDPncCda4msaDpT/jdEiWKiEDzgjjO/5Zv4GF
IB7t8rNWFQMfjOXBlS4Mq+In1ryCObzFsUEdNzyM6O7w99+vjnDSGDluKjTmNgH4
3+QNON8/bSmgdaFJVtsIB6yA6XTNDwHzellAk6f5rPsymTyo0sIUIuUkYNUOMaMz
WXBMwvcKusl6bJirpEbu4zcnBFWq5x8mx7gJyoRZlGm5fzrghPfCNAAtk3mt6Fdg
uMSmRkCqL5voCmPHq0Axm3ZgqYL1nfkd9d9+uevk6XTtasIii/w0C3s4eUUcPUwp
yWGsE8OJkm7o7gALKEqXwqCaXot3eX9JQ4SynyGftnC+kitkOooRnHZasYSlOQ80
tUciu5d7LA3BGsZax0aPM7Hr43qAk25u9W0gY4tTyav8B5oIPbsGriFsvkmu5sED
lzCbSsleFXqrn3ga5HmvExrUhwKFLuze9MRe5+HV8Q7SgFtF/fCNehZwFWO3sO9a
M7RbsyhtWMi1qZf5h8QYd+nvQbtTaRDbZRUN2vpNK9qQGtv/NXVZ9lwdSIHnW9EH
IbYdufAk6cne9r3y/kQVL8thYutXDbmIVtCIoQyLASxuxDs2CoV1O10944GcCwDU
1kej7fs6Pkx8xGypcajNZ2JcyQq2qpONJfL0CcEQOcbYfKWJuX2R3gQLohhwtWfj
V8eW2eqVuXrZCNjl32ZdxD/xa1fkV7+WvApQrRJvz3EDKpsrhEZrwV53Q/CW/YW4
4+SO/BLcbxDhCXvrlTiwrc/yFzhVuIlqtsnH6NEuka3LUUdmSYj2BaFGPOhKF1SF
21SENn2RJpS2solWsWfC4e4XGUge0pD0LxKjQ020/BIPDecauCGls7qq8k3A3C+n
6LbkXhKdX0+BfnOtgV7T+UNaZ0JNOtLkCFkPzSY5RuY+gUDoO3mS6o25vghXKqH7
wDSVEyWj2fn8/OfCXNcAhXjlcCqqt9ZENB9+B3y4LdLnvXXkJoOHbOKNCz6rfqXf
5P8q/ojX2VpWQMkvpVm7pxwmQnVsZKb03aI8+v3jZ8ElviHuJb36PlA92cBn6A1L
CyrUZlCgbBYgLZIxTkNOk9SDrTSzPFEtgHj2F8YAm1FCmXUI5xNeIEbfokxIYrj6
DuA9gLXo/TZVzU+ynAjrbCiLb/FyshRyq9aUQRu1itBpeMrb4siyXW/v/6xPwYEb
KP0QJwKgh9VVMnvZpRs78cfPOPjr4k91cExFjAz3KFdujZIS3ZgUsBcoaSaF+WTi
YUEEWk7KQeKwkxqV3m4W+fUfhzx7DKb5BPsff8WjVvguUt3cdzyRPaqRNzk8hRxa
612DdRVcl/PsrJNjS6jOIn8ISOBtw1fX24TsCgbhL8XIjYck5bQGajsD7mPdxDgH
7jTLRypyuzoKnbRY5dfDH6BnMPd0z8x0TzWonNrY1Kwp49uGg1YK4VyeBJHZmPpz
osNrICrSuzA6Bcx3Kuzv4t4HqCDdy8GB+iQP1oLs65g41LXWgUCkMRjIgIpqOqmG
lRjFrDt/J1xEIarVGWHRT/vazol+SgA+faJWn+uOsURDKY8qCtH31XJGf4hGdP+R
Y3Vz1NzVM6t8ewKVYZHhkg8ILTsTykP3Tv+jpHZghxZF3TBZ0rfCO1G7LxhazdUV
DcewY9cTLSTCdsW8n3hpCI+IwMMJRsC0p8iQOQ7hMjFE2seczG6OTuMyKpee42tb
IodMzVMv0IUAft3S4A32alZbcCXmUGvgR3tw1rAwf0WBGuZbNVqRBAPChoygPL6s
UiZpY/+/QIJMRM78Y00m7dfysaWlP5J4/BfrkKUm2R7gMlMs/SFNyeUmZbua7Rg8
98oeK4cKoQunJ93GMvEe+WXPHdWXWFuQ1dqEh05puSHkoCFkjFZXnPxZBSPVZJT6
clbxB0DoZYK1kQvFgAGzFZ3R9lJjf7g1zkRKC+S5bdtc2O/utjz8nkJPLfUZsw/Y
xtFVgR+8hYHhf6HCjJMd595gnay9Ks7g19Hfe9hcvIUg8PNSyTleXj4u0Wv6QOAx
n+ozAzfjw0XJLn+EAhWcPQI/QbDhd2+tJbgMJnGNoErcr7n8NUAyGE1sYEIVcR+z
rV0VB+SoQ5omFa8G4xEv/+OppIP8b1nKTwsdP1whzalLgKx31i0Ute1XCiXY+UcC
/mq/h9DNOo7CPN1NzUkwh6NP8OiOudp1ctqiuwwz68wH8fKQxeXEXC7hj4TpZzLW
HdQLy9cw87bH8vs9xg6oa74UsF4kQd63CnSp6zmmFGyW1sIbeA0n+zzSFmRXvrwF
UdSi0eFuG+8g/xkT3iUPdhIGaGYZUykLRg0sVGe2TejdJbKW56jcX3IJ2h6+cDxi
AlWuLTpGHDVfFEonF+RXssy6KWt17GIg4pYxrDQUpiD7jSi5OqEPARLgNzapSeTA
yTiRCmzeMtU9juPzQba0yAe23mbWMgyWV6ASlH0ciO/KEGVzZ3I3oI9pvmeXSNoi
JZBnIXpCjZYW0c9gnIY/KP5xXG8xg5uTSYyPlHiZBEmFSRvQRn9K2/JQRPh48fUt
p7z3V9SApp3iQPhgwKwrks564gcBO2+LrBdDk7+FGiM/TJkkiA65G5p/t+D3hmm+
0Wgp9vXDECAXRznnBmoYfSGNdytO0ar/NLWj5lDJ8bCKRJ4yciCE0QHoCAH/hWHj
HD83QMNJ9nVnnk8DQmnSwqwiZjPlQTtLQpwgD9Ob0bgkq4TcS9cRn0XORGg8R1Lk
iuj9KoevhUqesNTrUKhowRn1fzoZh7Z4PewaD48TYRxPLQ9J86kfkFxNiT+5TNxY
BZflD9D/G/HGFdak/jlZa8N+HAU89C1g/WXJVDr4JnEBImtxAfHa61AxYRGcKqYb
QTsgTEF6czFnZsnPK+uLkIt/rkXyvb3wQ2Eyk+3XHh3Tc5A46OZRmPKFBL8YtnBF
j/L7sA2uVo8kN/jpmmOFwshXVJfRBvYAIEu33HPiv/2vxOjbN0FKXvOJAiinfqou
xpjtCi4NXRT+XPSUGJ04XhTyXLPdSIwR1A4gQ8WHVhsYCU0sWJedadsFN23yatFc
Vdhz4si6JiO+bzbcsrY9FA7bfZHDRQ+swNzlZF5N/deOG1YoX/FxxuHA4WNSDvhR
iPucHzD57LNt3ugm6GbTFOIJXC9k/ah/sOEnfj4P+1hfm77uYN/STJZ2aKZlPiBZ
Wb7YaTr1yB9EtR3Hj3NjtRp/xOGVUsgY+3EDHz7gX8e7W4YAJOsLmxHFaqyW2mP/
tagIWyBfJcy1dX403BE2UDMi5CtP2TG2KpFbe/EQkI01fa6iKhwja2D2vTu4vagH
9DI1sh/UNVD3BaRfICJq2Frh1LgdEeQe205Bw2srbSfhjVCIChNSIYKMJyZKQhPE
mW3tN6FRfCKY+XVOy1xvYlJgByUwKm8y9YTa3qIjYl4wt06YhJdaJ22sQiRSmMeP
RpSKb4UsWSePoAs7JWHhrycgV8SC2sjnVoktx/IkarOKYXZvbTwGrA6fmMf3lx6O
AQfk7So4GeO82NnPdnlgBgBQs8XUs3aiHee+bkFE2kqzBqZb94QaKZ0Ue16p2Kp0
Xd+bB6+9n10aU+Zsi7UezSeOCV1fg8sZv3OBPsReR6dCny0ARJJKFkkVCs4pl442
k73akHZi9UiYrjATuxPFURyrk8104rTc+hpavaZEJbTTaIxlvrIhN3YCrhpV5juT
TESj/AVr/cKB5rlulRZC7ITU21/bRc35EM2QL7SiN5MOf6gc8kQsYX6NGBdO9Gff
AvFzTPOyLiA/2iKnw7lK6tjUmi+3cJTRueA9sKU+s5RNlBGGySRjYv7US42FtGkk
Qk2k+r7fy4EfOcDzFKPetYVt/bM0QdSys6jHpxabXNJ81CKNb7lmIbAtUxmUT1Do
ezun0E82I+2VVh4VFCuZyWVuTCX0bsVZ/EWHD2L67LQ1nvFCJUeqFNnwvDwX/mD2
WOySslwDfedBERrh5GRVJ+2IBfdq0muVjJOYFdiFIMvRc/QTdrrmw70M0yvSf6AG
DxVVR59XDgGzvasbn4qH5rgGVwCXf4QSCsumjdFWksgJNhUzpRn2HrUmHLVlZTjO
woCG+eFcL7XqhNIFvgO65p22JgfZ997nLLoOz3QPaeO+RQlr7maZyzOMc5mgRJhM
3Cn1Chmrm1VqJUi5ac3Z9P6mV9yhQ+4hMxvJH70iF6k83JNyoZNQ7br1AyBbM47+
T6haNLQDaE0y+uw14Y6SALVsGYOaycsvYUn1Yt5Ba4fivt5QKwXSVw9wTe133Ot5
36KnVr4ywFVqFvWKEI3UIAN22zhaU358ojKrEgQcG8JJR3ETegZldvGFiGypL/Fs
k/jZcXwJNXCiTwugF0p13f/tTXiWxoJ8/poWEcblHZbQXaYMUAbIQqW3I8Cdrdwi
r3AqA2yB3iOxzJGuDS+avIJKS675DwMaL6mzjKy7gftqJEuDHv9FV1igUY843LZZ
D8MTIwOZvhVdNid1C1BFeu5IpIB/jTlkygmKfuG8eqBhaw6uIrF6mQ2ZYF6F0QAw
aNLqpA4SgWwMAERDPtGda2J7gdrLroFcd0Qatr9uVQYLOgKY/1wQPLB0rQiaNfOL
RwgPY/lIDnZT7eJNm6jeDixF73wE+BuOBP0EM7YZTMRrUzTajvSQq747S96hUO1T
u48gt78ikgiF4FOU31VG5poeyWprUVW5yi3MzmjQEyZZdbJrvL68H8evzDEQougR
wA9BGZdB3NgwmpBkPr6eXHAEQHWYH5RlUNg60jaPATOYpCV1og2i1gsSYvGr4ZkH
80VAHtQ7IeovV145qXX1KiyNKvbkLfQMK4QYeq/4N+PS1QdGxsaroDy3ZYNYp9WZ
KDFkDaMhAwXyiVCK0pDcVpXqI9HAjCErOeQvw3hE4EUQl5zJv2/qMRQwJ2efP8+M
L+UHwQcD4vVuQvNYBuy3vu5R2RwnWSfZ0pQGHRc7zIaOqAB0uC924XNk33sKryjK
vp5xqrIEJWUqVToVd3Jz88iQs8NsdhJ2q6cRhlDwiSn/ZcWg1Pp78snZmdqxVBF6
cndwCi8kNFVs1DQAH64XUpV5VJLqNQNi3v3NR8UIlZZoH9UDYak67iJ8tMTfqXtH
QhKi3aYrEx+NpvgFUdQ/MSYHxwycEUtAqo3LYSBpHlbjaQXGg/PGa0gMmoldLR8M
JZHibYhZCWDDuhcuDXe9IBAeJmR5KZM2BTVFJxhgf02QWYrr4AsjN0SqiO4ypKwu
tDIfQflocJK4G9S5tEUwpbfT7IOvbglvWC/PwBxVXhvxCB71VcRdwAIcZhRx9DVQ
c503UecedqgZvr1h4BEDKTvvGbTacl4867nm3eEYpJW4GFlexrnfymXoht9CXxIg
+gsIaL2B2Jl70DBiQkaoFV5NaCvGkXvez/6nZlHiEsejFLAYNRz3Gy+Yb4/8MEn/
aq5FjRhxLhO6EIKDldmkmfuibq60VHGD6nG0Ltdg7sFXenoXbuHocUXskty86trt
T2WYqOI5JfIlZuSgVfuufxOZdGIRaFZQ4sV6vgdqaYk2mNVGSRb6KXkRoBbhdZAq
GmGjcNUY5n7dlFUNzZY5OJOosGl1iSo9tkJb9p8sxRmRsXVuVy+zGYENwLX0N+39
qrqOsVSL0Se7iLo8VHtghSVKrgIwcs0v6d+hci5CLfnvYKtEP926vuEor87C9w5A
KU3Je1a/KDrHQcOsld6fHi8Se9VKK3NYKprdDY+YAPONoPKYLtfBFE8L6HTSAkXn
dw6x2SLiEqF+ortO+5+kXXkIMfZ8YVHKvpk4AJ0SOLW91k+Y0L334n+km6zSp0Z1
GLsAXxPhHMFALbkh8Rwgni3fQ4D/YvqqVbXJxmOF5/Hq8hmCSPMk4vSU5/VDqY9T
D7A1GzRylX58rtiuhMn23FkJ/NwppToajkO+f5BEpbfvMtqKr3k2l0sdrd98vmQQ
6Bk3mbOHnrq7DAL91+V/VS09lN7SQTtRLTD1vmSkBT+oF8R9kGcw/iIruERTJGG4
wrBji3nRlJWtTXXzmKJhqPB4+14c3vIT0jqgBhBsW1hdHl/eHuP+jCAk+mHvVQ9k
5nCVSr+y/yfpWBLxUkWU/RodQGG3ILkOzHr2HSgKiJfyCNagEoiJDM/qsC6wJqAo
giAbzJaiupsahoTd6pYKAGryCE8cdhN/nQQ+tdSF7XKh6OgkHlHF0RAhPbMc0gLz
dNovQQgSN3L49oEH0+Hf0+Tw++7wqQxkv3adjL0A6JOEVCj+PJGGmnOKn19U0BCl
ZVCPDYXAiv+PetQDjU3lXrlh+gancNsKxNlFhwcDR3Zw+h2/xo2VIctF3TjlYQtK
e1br9Z9aIHkvRlrLMCcPYDdiCn023O0tqY3hrrjvq5PCMVY7z4XrB6aW0XYAdIZ9
p9YGQpyGAI41YzY8X/dkBGa3Poc9CDQ8KEwLaSqj7eE/iRsjQrMOfy+4mYHG2dvc
rDwC5mpcJeU3xBhrUpU+D8KGtzPp0nusBpY9JEq7dapvw3v/XbI5QQ9gSSHCjSvt
qeB6IQG/gelBDDdz7RZs+p7o2IOJxRLUenvYY9JRfGzpuI9SD62bgtw+UVLTxsQ6
3DaoVs1QzJnvXDVToOhNthfEw/Tt5TP7xh2KxLLiaZb4buVk4DQ5tYlRI9wqKe3L
Z4GIzkSaM2GMh7aqwIhwn7VmEzMLdkIpOZ+W+NKNQnDQ0uZitzIAyGqIn2+mYOiH
g3/Ujh7dxn0uF5G6VHNWF1gDQn3ZfaKZpGC99p3dIwrebYm96HDo5hx+MOrMAE42
XhUzlX6Qk8UcXcY3VcDLJtvWjom0idang281+yNIylLy4xvSIi+14e1gfp2Y1irW
QCTIR6ogjEEQknAdN0WzAzQo2L6qs4n2SAL7cHLG5NEH50NiUp2qfOLec0cRQ9Rd
vwBGcMI7kdMATQukYPQzu6FDJs8pt3gyMUV/Knom7nqcfUfd83COVOuqOtUHZKoU
QcH+OAjW0lZbUE+N7Zys5YyR4UMkGdA4tot0i2tgKvPZ2MqQBPa1S+jmn7+w1EdR
0twj7zZ2xMLlZOCiMVx44vYfy21PvBgcaxW6U6ND+9F3ZYsJva9chkbLPoLWG+cR
mZXUJDJG0Q3FZEe0a92+Ag6UJqG4Die9r0WfFSVFyGgO1SM1Qsv5w626ZI90zYLZ
9hggT5diysZbZCQZiSvmGsbi95sinQbZzgnuzTsRQueTGZiYt9A+pl8WVpycYpQ+
1KpmxUS36aTxRegw/byJeelxPMrr6vsMJZfCvpVZcUuqf+s1ARxJZva42lCHEp6S
TIJv6gslXZoLiK11GlIAOUFUuOyyIPx/Duel6kpiUOS1jH89RDkVmzkrFxa6D1yL
52K1WH0wfZl6eops235TlBlJRISJXJXbLOEV5c0HBH03ypEBRBAVGki6i03opm2b
/n1fjDcalElG5d3/GJdjaG2ia1/z1C6Ye41rCaqP/lfzy9/BVRnK/3+uQCGWoam7
GTJ6dnQ13Lp+NfbDzKihpJZZlGp/KCN6YgKLeKKHtN9pOHQ3paJw/5WaD47iXagH
6dNY53aKoEyxbxTs2IgN+h0GgRDTWGC6NkSZIBOzexyPH3ebWJqClRece/j6X4Er
c7kvZRtw+SlTZPOoMEj34RGuigS9RKOikDu+Ax4l4Uu6oJbI3LlBnXh1UF63spdG
3zg7RjvBx47oy7fu+1B1ybI3dNVZMoM+VVul+naTGmjemjkBGCZHuVnzYGBx8DET
lU8mgj7jOCUVESJnRTfC8Uy+LBNktW0LuVm2nX4xh7X5fkbA6FMokevcKJo72N0d
5SQa62IvektCOfEBOjO9zm+5unmQNY/sCjc+609AS1ed+lyKx+quKRneJOz6FlAV
6T4iGxKkJTD87yG3w9Rl2CTDRIZWt3MBA5/j9RtcEfugAJ1QdV8rRaMi4mNexSiV
WSFnPhCXehOQGCp0/CsN2C5w7Mw4OzpjDXRPtpbg0iMUGHch8vH/v9Mv5vwxgQpJ
ChM6bPDEo04v41kj+1QAbf0Rix6wCNoQkOW8QQT48SNWelBsdl25e23z6SQ3EDJS
xYyCsHXz+JO0PVhiTOowGQnrVt0gT7y69O53ig2itfPdwrJsLx/fprxAZbm+1A6i
TV6qerESPNG4E9X7CZ260OdsyAHoCJmR2goECrg5HJGai0+gm7dPSZkHeWyWv+uV
Usbw1igWEI9/MrsT8CMygm3qW56zX/qyHSYtxe5upGzNv018EgM2r1dh+VlZQg04
XsWHC3PzuvhfbBo3ZSmfxpZnPsKMQVcCYJdkkGP41c+fEVOl4snci7E0XptMsrN8
Rr85/mi92IetwSx+2do4GT6VpOexOxmfpTVt77uH8D0504svFCoVqfuK+mZ8N7kW
MK6h2ysZnqs3PxcPWkHRjMZ8GMWU+0xuALjNDMZOABgDrq6+fMtBcU0Iw9GfsOm0
xU5BvizxzZMHGV1yJ8X7dbr/hlLTWngf9Npn7hLabP/pE4xbsHKIUsMU+DiQj3JE
c9M9rcYJ+CdDObjH1vxNOKiFgq5k0+1pFfO8NCT94iGZXwBelTFxfS0dwSTWmFY/
86YoRyshiK46SLzgjIP0jOLs8QQ3KhESBb+LvGBn9bgP6iZA9w1sb2crQQ7umqVH
abCVBLtgu1BlIiTLgbiK6fvasRmsAud3L1yLOzY0kE/Jw3uHELaAHDKOIcr+I091
tiwH4DkleL8+vXAsd/d+TDzgUl5l1j/WorKiZ8gpcwZIcsxAhMX+6hy6TYVZjvJH
jWDFQGjghVVUZFtAch2ijPquu1h3zfS4d8qM6xSPxJWkjq7p7+Ucjz+Mskhry5tR
Xs9SGZ22ZOBh1Ew5XfjS8OYdqiNdAELAtfaF6RHhzX/yN5sb3o8cfWV2XClPYcMm
1F0SXebaMBu0X053MTCk3teOA3zvU2vx/cjtcGijPI9xLADQ2mKc9k7BAJCJozpF
p9mcufp6dfVtfgQ/WQPgMhRICiHatG84YLvyq65qgVl5sWxYUDnRnbx8noTuhduq
45Cq2BTLWC+cL2it5XKNyN/2Vbx3tmBapwBOWprJxsTsaAKjYnqL/g4Lb1UQr21A
tSpFkcOAD2pEbJh7dQTrAyx1BNY6vcJPxYHMQhOhRpvfur+GRPkleliEGhEE52L4
BVq83lJNHzEKik6YF4uhpdYATLqRgwGH0o6S0NRLZQ2AdnrxDFZBnuHjNyoFqTFB
QV1pGdxlBr8Wsv4WfHoLA/1n6/jhdv0I0B1cKkF5jUBri6fBx3HlhgQWk4SeJCa8
THjcxUFHizuV41cs3R7KUro/Jx0oJOFwVfxD7f7/UZMT5Ckw8Sfo6VaaoeGzSjC/
7a3OPNfxH3HzXL2V2qtm1UXUysIHVdfKleUeNkWQrtHVUvBqRYcEp2DIxGipZgU3
Sy5NJFNfSSZXsxeUVtHcCuulhYOpZUKO99pG+ftJ/I71i5xaMxFGx9QuZmxOCkvk
DPQ9FtSMYzvzyPXoiT0lJLdE2DWDpT5PdhsTu08y2cq8gKT1WpRq/lVEPQs94D7R
fKMpCDTe6gEtS4A+vjiPBNWYCblIOLkY1LYrwASJEkGJ5qV2kEFV/FC8BdZv1KTD
yt1IMZOBnljbvBP7Blok52cO9Z5jz163BnoH64ZMeJc9amrVT9vzebERutKi72XP
P8OXRPnIoLf5uzcmw47TjppkZ6eUw8PQFc76PfwpEEZOkUS7s9shzC2JuwiGFqr8
jy7SdwPwT+IStnwJiKXlk5H2sFxzxwHDxkPRV2sfIZE44/zPj+VldW8Eg0aFkFTn
534V1/Ue0RvrKS3sHbSaGPiqqPp7VFEHbNtzioGBqrBP5jHEIOe7Uue55qiKZQvI
NVzGKC8MIZmQKkYlLEEcht1r5exNfdPl5SI2QZYfpDLrvKoqz+u633AFFLK/Hl74
4ySNHS+nr0KRu+s4sw/d8q9q5ZUZNO47z1v9Xzu9q9N+ClmoGS+KF/HPKUJ4UcsJ
63teb9SOGXnj4JOc1V1sm4byNpsDnsWvWYQ739qo+QBs6eH+gB8fWuWmDSjwfQOu
j86tDZ5llUzq3o2cdhpexqwUGq2xA/IO1TiI4CJc6NvoX+k0Woyg5+J9O6i5+1R9
COJ9FtHbzp7+e8dBJdTBYiCjfcCXPlQh1oE1yLqKkBfgqR9tfV+tHUiCEM+h4oHK
Us1AkmvIWXiaLooHg/is10lrvOyEkvgPgpamcUjdVW1jyi8RwBZeDPi8ljO0yAYo
Op3qLCRGDRrl1xi/2X1og2gCM14TwZNVimW4wOXiHfum50CiW34GHOAFwHJPG4BW
8zL8XtYcm77UM9qg7HrTADoR8lpxYioVftThBtpXa0sOTqhiCEhubUZM0yOsFR4/
tREOMEquZXB//jmUuKrLx2eiDNZXJjPrtH6Ywfxh4pSbFNhYQD9gunJHNNKGDsmX
MJmSaVNUcjI6O/iQXuqRs1nWIH3UaO9+IUJp/ExklYv0c7dYf280dnYGYIkYLVvP
DvE11TmQ2ZTiKAERfYZ9YtO336fM2YeQ9EUd9qgv0O2AsvVSIkL3usB4DTodCVX2
9gW1K9w8TvuyYCs+7kp2llQuVK2rdt1eJ8gaGxIuqd//dVwuRZjnwjAvqsHvmtVr
6tqgekVeI63Dz9bWFRghDIggWsk7uUgBvVDVEeuoaxwM6znhy1MZ3vPy/WYw6A6j
45lY8E00bFDyLBCtPChjsaWA4JYX95804n8DjXn4dQJ7BNW6/hGwl6qA9syRIEsb
TDqMtDQYM7dfKgBcFW0sDEEZgsQ2cxvF36Oxyc+PiDXmqaw6uVLyM7yWMqP/vbkA
Zi+fAhLXaF2V+XM1ZyFgT/YMatu3Itj1IDtMx7k0XsXvNWLQYYVBi+BbDbSyNCQ2
fTqyt+jnd4aTL97F+nEgDoqffZuXBUqhXG6rqz/zn94OEguo5n7I9++InnXA4peD
UXXVur8/bKMrLhcfb5HnF51BV97rBvj+K/gGQHea+rPiyjJqaQkMmHfcKL/jH2CU
v1/oqt7miYalQDfrMq/UvuCus1ZnwAM+eFxXUlVa5KA7hV7mzCjRbzjposWy/COv
h1rBwLPOcz4K504e8JVeTLzKhm44k1yuanogZd2tmHIf+k5NQXCdtHsdX/lbTsES
CXIY00ZsWcWX0qRAS//Z1klP5+T4Cqd2oG79DP2BsFjcMXkGViy5SYGjfVVOKEco
uPtpP+J3A+IKNz0bpg+CwwMYYtkBWkaNLe20ruiUN81FAx7OD9aXloYNMAfBpHuy
+dXh43za2mkFqfiFXrsA03E2Wwh73U0naMMgxTJlNsYnz2iWkn0vICGEE3rGswK6
g1ONugkh3gS0NLU6Q18w61FwEdKH+A+ck0zcyZ0EZrWYfaXaR2Trr5d9+0Nt5ghD
44cr3dZaoYPNgyyp0EjFJHlvLbmtY6vLI7BpkbJGnq5VO2+5tbQP5OgnYig2Yot4
btD6vXgZlLWATj01fcn/QolsyFgXepdaWCLHkGIEp+YogZilDo4IApCaR3n0j4CZ
AFWWcClMjRx5arwMAES5ivEIKOcTkOYecX+NdCkFC1pgFhqbsiELbL9lmB+0ExEI
TXKJX1slVdCEemQhXOmbxoEYSCopxpnVLo7NXTE5zudF8Rc4R0poSRlasGScfZE2
DkT0pt5mwY4rFiV7qtrAEOguA1yP5KtnNQ2dD4K3GUKg7HeNEuPDSNUlcRnnGTtA
E4V7e8E8qV9uQKxgUZmfDh7/DAKg9kU2m0pKfQTufYfgLt01Xi+PTKKcin33Im3K
4JzjpZGpld6C02vE2OuPAyhVgGDXvcGKdwpEgjSGMlJ7MnlOTNr5BpYaTxDiqEtL
Hlfl2qcv9UmdbgcuMFNO0wzDoTxsk73SG5F77JAY+6FCS2/6fGvb0Jj9q+is8r8i
Mbv6L/7OEin9n2XMKGBoShjLZH11p4ZvAD+o2pSA+VgYJJH3vWn6vpo4cVAXqz9G
ikW1LM+3UxxlMSuBOgddC0tTfiSawXM8V4oUrZHF4xCvX8mFdRqs+j0D+9Ji3sMF
U1IQmz4TWRphuZvaGiqA1TUfIK0u8WqkLCqZ6vS+/gxuwB9poNbzTqI7HmdY9z6t
7zoCVN2hyoPKmqsfEfiaidaP5YO6VLikTNBktJWsYdIsTgRyQCVNNAtJ1v+1ANPF
/VKCS1AeHYuwuBLoYe6Fpi0pfSIdoPlNfXtj4INtIbEOomFdZtNAle/GssX7aPU6
h4kELBo5Vuh6lCF8qjXyMkx1jgYk7gv+qCifFPaCB2aXPa5Oa4LuwMaF/zH50Vp/
OUYJ6zq4GJUtJW4i459yXhlBbvUu3xxRzBRC2yuZ+AALax2itnJ4yRxbfUsey/cu
l0QubZa/d2s/5ZU3TvvYF1yfwyv9pGJNo6G/7Y10Kx0SbU117zU2DTP9DPMTXFWx
VKl4TBxwJ9yAZqe9cGnUP2kb9VBCVF8Pq3hkUl59p0AU5ajC3GfxLpkVAyXRAz7q
Y4LBmuxOHNwiJNaDC3QJ5RcbFee/keDieMyRxlol5tdBbaQWQNtLy2tEY11CxHeN
nI1xLnSOOsZpgxb4D8YTuHTc2X74CQr0miGGYyp3/Mx2+Wrzj+ZwAdjPHAJfqSzV
k/6OuMgsNlf4ETN2R9MhjZrVBwoK0vJF+N8UojhPH3xTUMxSXjl/eXOIl9c1kjwz
pQzRSelXjYNq8hvJepddi3mKe4KbpBUt+bua3q2Mc1K3xzj9BIsn8xgqBX1+KnE5
WNQSyxX5U2I6UjOx4LyKqCKe6EacxB0TGILQyIImjqFpGpSveddu7wytIevjp8oY
SQ8CHeOj50UnZ/1e/pQSUr0xBGRSi/+Bl81Crd3qxa+gkOdYHOVK0RxO/g2UOOqv
vGAx8unHnhjoQKzHKA6B4ZYwO9TBDJaOGkvljDlVrC2umk4Zh90yTRoAm/vqJNIP
1cGoVd9859Y7IQQJXibD3A87LCBBQnlRVeJv+SGPl1qe4+8KyT2WLX8GQbPb+xi+
1LT646pPWuGrC5EMYYfd/vH/D62yYS1R3NctsW3bo0kizO+xEd3AfFNPuQA9rKII
Mk+pnMLd/STiGjTnf2b6k04uKrhI3GDmf41Ic5xd35GmtsFEbq49ZCPY2MswRBCa
e8MTnLAl+sd73rRSgup/0R6otf+sZrKNvByUrRIU+GJjr9eFoffxLKMZwjyyN0cm
1LObDvLqd6UvNQ1JrY/+3kMZDEzDrAZRgMd8rBJ4ZQw2gskLX68+4yD8PQkzpQhn
i8qhoj89VBhX+pz33ZFvI9AOkMcVFfQ7EfCMOApmuK7kgrL2fkRhv2Gn+A657qQl
jfuCHInmulZpROEjUgSJImvIMX1aO1rjs5o6IMWfIZh+0Y7eBlag0uCoH38hK2H+
MtO5vMHO1rJvzWg19KFm+L6jlXqKP+rn7sek8IYekVPXfF2b+vsq+L/36CXTxSM4
hd7SUmcS7aV+biAjvLXqfBaKYbnHfpzp7w5C+X09aH5Emmppz8+qhOGfgIOBW6Uf
he6Uo+aMxusiUsCgHsTMsaZKGJouBDP7d3ZDH2B+ibJ8AqQSw3aQrGZGnLUSYZPS
vDmQTuGOAnGLMcFfdUI/sz1dZoU5V5XibEg25SwdG9C3pLSM1P4gUPiFy2U+nquV
ZsVUl2ZfF/JsFVmvnbeS8QXMTbKY+Vf6g6yeas7i87qHks50j2mUxY5Zws3utAKf
4kCJ3RGsPelp5iX2qFEUx275y8pkDYUqhhyQg6geJ1ekEwdbbMeTa5koLTIIhEuK
cwOPadII2Gq74fO/7GaR5Uf/MRPuWzNRpZGW3+skq6NwUb/FMBYgvdwsxgZZieUs
nmId231z+z6wfsFMZmzBqRXZ9f1rlbeuRPVFFI89Bo1ZMuDxwNmuW2DcYAWcuPqO
eQXaqOhc+Rj+U9gZReW4hgG/RDBazzaFHcG4YohIrKvrYoSYDqqcey7zzgK/IV1v
qgxc8tc6wb6ijBr1O0L0uilH8Et6VSkNjjJlYLiEes+nS6qCSMoYMHsakqs92ibr
k+XRn1p6UhAiLlFo++y3iCYNkl+K1HL0nLOu0WSmZ0qYt+lqGYI3X+4X0pZIW6cO
2Z4GaQxNcsoWUrP1u6PRrpI/Idt5NCvgajO2JkTV/VVJeMnCkEyUyC9eaBnV9mGP
ViNuIlMXm2D45cWRoz1lbN2Re3C6wfjTyygHk1e3aVajOyMqR++SzIupv7iGXz9v
R+zIfnasdfQFgGL0VEDYvKrLvs6Qk3XGi9W/FfeY7/xVeRjl8hseO8N2ETEBOTpS
KBKi/w/EaFXUwf0TAzN1CWIh8IGczrS+UVaMR5yKyFjFk71wmnKqyBuyiMuSRgXG
zV+Gz5XkChpHiDJSGO7CBicRF2hPIvlYHWtJv3njX0Wm5+6ho7UaHNOu+i+LzkG1
LdHW6NGHLi7LI0rZZI/eDzDmQ/zs7U24gCgXWmXFlUF4+SafjY9HVCcAVuC5kk3D
K5GxTBtk6bYU7Hgf8sbGFt+V1rdsblQxZ8sphesBo+gl3hYCmOBo/lnCbJt0W1Tv
JmWVEtugskkApCshQ4eLb+BahMW9f8EUhQemVmgPUrsa0EQKqUklS1Os8KBV/VcY
ETQ4+NA+RAiIsHSFiPW7uNTUvNFqU0JVDoabLsADl8cI+StnZ8CmWgFRmOdZUuSC
qrRECCVHQry8WLMiZEKbUkNxm1wm2Qs/qSBSyddRNjJctuK88BB8k+8upzafHE50
DthOMxX+FoT2SHw831WP3R7OzubA9tn/qqbLij0hcDXZjIQq1eC9E/bCBhXR3u73
IJvp94YiPCWIrOnvBLS3CsUpX+thXmzcQ+BIgXPznkQh6Bn+D4vb0s3FmPFfQ6l9
7408WK1/HtyHWmilp1X8eESYYTrSUGpBojiB/eyZas+3AiRfHGSOV9pMWpk/S6cs
L+o/4wO5+fm2SWP4NAu3pND9mEehwSbxJv1MYV2a4rUdsmw/NvOMMwo/iOeft2z8
Ax5VTqmbFv5v+luglBDoRhyV/SPFsAVRj53PHGPkl+eRec5+iFju2RzFhL20PqSx
kmmTIxflVfTRaQPZQ+AQKn+nY2797Bp/9BawDZ/Uu0tveDNx02w0k+Bf3hhpBou/
49rVPQ1V5SGy9XXtmR20W91SbISLEI/vfzBtsRROkNIgWDWMFs6kLV+aai5r8hif
Pb4tZVuGv1UwCcQcWi7hcFH358xHcLcknzhevqgc/848ayKK1rIWnfyQBBEmp0Rd
bBmi8I8rTacG1oNiGPJ/QNPjl2x1R9JMHL/Xx2sdNI7KLjiBOzTvLkDca7VU8FWp
cdbLZrXgie3pa2p2D/9HKPV/oW34FOoHGKEQw0q5lv4lhkBIdyyUOJ84zBRgNcVg
7dpToxVI1fs2iSrOBsirli0hy1a7EPqlyRyCwewxOHHL71C4IN0xxv9VeEVmK3NX
yL6A7MgXPfxDjLNe7yGMLXfkDwdKd9lJKAIKvbfRThvmRCdB6EQMTDQ2Cd9BVmgv
RviteZX5edXNctwRV4/P4hv2qqdgaxgANhVsqVwsuhZDWVOWPhBBsXdgIrknXcJN
77cO1NaZqF+BDefolLQO4NCMXq/c+WhMLtN1emOeDUJ9G/I704JOdY5Kz3EYAXCo
TAp0wTsEY8UlDHD25nRsVwKFYLqSBHomFVtIY+cCHqnVI6pbvRdkfDDMx5hCP2kl
1EoXXB08na6vpgUGfveuo29JquWn8xXRrwzeranJ2mrM+6j9d4WmRQfoYTbbqYwI
hsOcx8OGayxZJ2S9qj1E03sSZ6EwOiPiekJEUlBQ0Ppcvs2suRROHNu46Nc2yiAV
7mv8ejOViPMtPlgFCUD1pIuT8k1clSttyHzBFXndFitS9otBgUckc0VFVBNOZP+0
yxboAPK/Q95ZzZ4sCXPTc5coc3Hx7L2s8MY5c755ZdfNAjZWlaftmbQX7XBPcb6c
8zaFQXcyCrECk4fWmMY0ZGXC+dk1fMT6sD2OOGmR1bNaVQjRRpy9hrezBAmVIjq+
u99UzZLMs+X5pJl6dMYU7tzYlAy3MtmvQ3vWc/sU9gcTqQlnYKejl6h1paa6T+pP
u6pbZXtdxxGQGnuUAeUim9JPeYOwh3xbdpVm+NgEr/o6hzgDEr7RHGnM8lhMWdh4
tTNvoU3Auk3tteR07hzAypbryJoX1zjMIh+t9IL/BnIcN1I0RO/vYWPGxAOGGMiM
LqwsTTyBsTMqxs5wC8Z9XOxFNPGPdgXiSPVy/A/bCt4xYRT9SCllNdYbpduyrq9H
PtVU7m93pWU+af0XEJLAU9a9mY5AYngBn8j7oow4H3XVrHAqhCAdTqU2dMT143rZ
Fc/rZ64/9XiA3bjjQ4vbYESWQvbH+s+EBDQ/gk5yZRO2516mgwRBotsSYh8BG4Cb
hjDnxHkh4AHoDoAc4YK6q0rnWjof9RPZS7lKA4C73FDVNSQbkrJhSjWUjRJDCY2i
VBxx3Bm8Yc13pte2VVHry2egk6agRDXvryhoO5l+7sw61tmVjdihMyJTv7CqIaZd
wkGjIX0h0zmF8Rwb4E1TzpekTlGpy6hv/TozH4XR7C6YflI/aBk8flHrNyV/TlRU
XPPIBuOqg6DLOw+3m0dRlyt1D4qz8VVfViervAvw7AJ1l0nY7w4x5kmGuO+5YRVj
cV98X6SKBt/v68dWVMOkuBX2wtr49dsA0a6TOYBmKKW9r57lxu7KaYzTfqlYRGzy
HiYHW45rHDe3WpIfEz7m8AeqTxw3lKJD2GIBDE8mIoMhYq3ZkPQy/Z/fiuvxWLQP
F108EGaDvqT1RhuXBUfb5ZNIOgj1Q1iIdRh5r4NZcbpG1TVM6w7VizrfjjS3oidJ
J1DRB71rf17HPRbKSJi8tZN4yUqeq/+pPaVjaIBGAc7HJ6jX7e4SEF55nM2DYvXI
gSju7t4auic0eE3SaIK6uKWm0ZDdiiOAQpyum+UUnXFywBtvNm2iq55GELvKCkKi
sH8HBld9OmrSbobzDhjuLkVsGjntdlmXKOJRbk8eSZ5I6h/6n+mUwV9afeHkXojs
qtskFUdVK6n5ZLWeF6NNTf/QNiVeMeB0o4YlMr6w7qsQ0UeZKXWS1C7O982qmYyI
yoJgA7uy0IYOJFkX3SBTmhYPNkq/r7wfwUjIFYv+GguQiE2GT9CczG/oyk2T8lqP
HryQGKV5GQOZlq9YeciziEcn1nU0t4ANK1f1p13ZgPUW4vycr1bsJ2KvDeoj0q/h
kXZXv1l+jeIz+dFvzftxlWItgMwO3YC4aHOMjoHiMbFAEjBj9180JA8rgrpNDSGB
eId8eXkEVqCT3sd9+zNPRcK/YMPOk/c9qRQZ4pFhz18cpBmU4FYOed5F/DbUJFpm
f9oprte2nyClFQLeSBck/9eS/937N/hnT/sdP2zGNLzfeTuLMCeS7iC08LRMym6t
3RtpXD7PEIBnJuKp3Xz0lUM2aK+0oASRXer4Oo14yiDqgRQD6UFNjAZ/HdmTiHDs
TurVocTZlITcJy9wURHU6ePvISQJTL3rMn0lBCH3vwkigmMOfBUfL+5fR4VP9iSX
Si/Gqm64v67w6oLhmc1PcYyLQUrGRhYx8wLJ6XcqhABoMvUc0621EVOoP3i4HXsF
BuY2f6apXOsrgdjtJKUszTwyBxModVNVZLFJ9Hp61q0pbZbqZVEMd4JQXEePsJQI
HZ29hgXoItY8lYdxXVEV+6TTI7156CGy3IUAKDlG6NKdINum4CqfJJ+0SgH6ycK4
imWmxjBEEO1iwPgFlYzofhUNhjelcAmYGBYb22xu9PhBl7bVRsiJx6PHcmwIBbIq
c8i99GwkJl2CEXZn+t7h5HP/WBX8yFhqG0Dktt+bZ7slrjR2A9RKw3bjtizBSAR9
q7OF/SvRQGLhE733iORHTCQPEsyiU+2U1gfXlGIV7qEG5185L0i2mGHmgf0mrDEm
gfaldH8zhGdiH2HwJO4VozkXfB0hGk+9iNeTL1rySjXQtAfIrV6cei7B5IXLPksj
zl1zOr23x7Q2L+q5wsvzMs8hQ8LYWC0hpYDJlp3sjnSSYeTlUiaTq9EjsnmWY3R4
xeKVM+ls2z7yjXuTG33sNoue4PzEBDG3eVtDtf0V5vhUYLpL2xg/ENUEwiSH5hES
qJRIjRtFYrwF704HnV7TQwqxahLlvhVyrmODK3k65hjFQe/sG+gpcY9ulbE1MDNh
Di7q2GL/vID/BzyM4Oqm27dkL24YQR7X8DNaFM9SEj3NecuKY7/w4UrPd3ibRO6G
BboPnP/HxZs03syoiQtwIIYJxHBmRs74vhpHjKqxNrz5abph3XttQEyrfjYrHotm
6lBULA4q1ucX2rOnAcm9X2AhXjaQ1KrVOnL0BuKLlg/HrRVC7xSQAeGLDghHeTcD
rtJ0WeNTUs/VsjiyRlv3zyT3DqUxxVdnRFl1sUwnn3MK5W6uJ6YUcyaduM1mEy4M
ubbSn9XMVScVPSGO8YtjivnDwMbDURniPv1o2UxNGCHT+uWIOtzPcMboT6xiY1EB
6QnJypX2mEX2YCE4xeY/4+8faCZqFzCDlC56ApEXfiRS+2wREM3+y4zEhPlhfQqh
20Q1JuodUyZh5o50e/gkyyhu9/SnQnBWCt8KX0JslGG4ah/WPBwucUGnrIj4yAPr
wcZXZPDZTXEEXhK8h4IZ85H1mPoOKO5Cf+NHN4lFHFNJZ7IeTNLuGtPWNZS/Xxkq
UxK8jPfeyxUkMTSUg7yf1Jwr2lJ9f7akM+fjCmPmtTRFriOelQ7Yc2qzgz10iohI
sL5HCIIPtfRE/R/EEyCT0q1s4HdRUEdAejU8ETYXFzwYxfOwiYVaLdfwyhOufIeK
f5AAYqAMAYumEDELJ2XHcm+Jok+PPuC1y+Fcx/+l+3RTCuWkZ1Vt4HA6w+OXLV+1
rUKZugmU5WmbGwu0Co3xUivMKcu73qR+RiJJsXQh4WP24pV4rozJdOHZNO1aaRLC
otEUp6qSbtMu5SIDmBt4SzPP1YRKDGovh79vh6xjMAvSKK+tAFvUnH2R1rz3Tdt8
VNuXsVTNURLzEDgt1crIRaI4vt0W5yQYfgMeTd6Dkfm7OEFbX5pFXZdTYhIata1f
5DOgVcKY8ekRU/CesbsKgcBDt00j2hPFI9c2kBihiCLkkp7bXht1r16FUqzG9xCT
bhwqxLS85K/fkLvFi/ELE7by/dERgJxr3+R3Adjo7GCod27JiGhkCvnFNc/2cti5
U/c7/JdL3RxmSmSEMQeGpEsstCpPUx2MGU40Q4XuXVt7+0q6mXegrwFW+qvnQkZp
x3YnhVtDLWXvD14qXVs0q2E3ctAjeZDlex22ozl6+8gl7CnXnzlYFqEqAVR1SNMc
EILZNimJcFKoQxnDN8nb9AdlBiQ5iaf3VfUfyzTDU+PSdDTRodeDbUK/TjimLmhj
ndTekwZmsPk8FO7m3T7ta35BmHvdLuBEw42uIf+3p1a+xrnOny6fmo8SNU+GJ5MZ
WA38WjygKbpAPAMIPRlZVVsGO1nkr4FOAPXOufVr+2GUuEUcrhEnHvEzXz5j01vI
hZNU68lj6ar2RcUDZ8dbMqrbczELX2sFbPfofGq/kREznxzYGEasSrl0UaTcVWp2
scFTeYpct3JFfXAorxG1p01/8aZ4zg3nwGMNYGhYgHrPhn6qc92Lb8VZRlU6iAoO
U8W4dbjuM2t/YsGUd/V+1CE0i/MM2LAbqSS81i+DJwZhIQI5GGCBO53zhXNysazG
YdDwPAOcJx4JrL50MQJQ+bYqrkfdx+4BIpamV0eRT9ZSREh9XNsZ2peTB5MSbSp8
ZmRxp0tL2dD+UBi3rHkkZLzmWLCOaOeP6RHwfXwqesx/jHGUNdaSJdNxVJYOyk8X
Im1LBCG/M/bnMKU2SFkpa1QIz+3V3+HVhg/E5PhuZvfHy07ATCeYMUs91LP6TSoL
hwRVLdNCemgUwvHRsv/lN4G5D2/Te9iLoRNU5KK1ULXdM/TKr85I8I3hEANy9t/F
VIvVxh9jkegIu9pexpJRWGH+PYWRb3HvM5fovw7l8U5sJNmSm0dF3UJbxj1RH9bu
o0NslyZec+pgn8mUj1P4/OcCFCyzReZTt+thNCoMlgK32rMl+2SZmwy6f3C0PRu3
6vw5MnOArGHMHXmcN4JS6uwqiMDY0PmPnbn5LDAqkhQvohLg6vEeV7dDIk1NwBqR
jar8CRWYb1EuxzL+u4nD/BfBmJT+wyTMTe7BfruPK5tDNvtPMl3mqq7UpPPlqK8d
HLtgpUuu/w6oT27h+8OxRkyH3+7aJkZQdz7V67lpMQXRx9W32GZlBPwzFUDuQlOx
2200NnKuYvUvn4is7fVrt0hgmLWy2mkwc1qP9kGmkLG0cM4TEDG3qOdd4fSmwukP
MjhHC3S0JNgKZ+NnHo7fCAl5lWGuLKG/Wz/7AMGQC9GOpTjd6tLlOGilHjvHH45z
8q+Y3xN7E253eP2gCk3ugU1zhVHnQq3gD4KHLvARU6mlG7rHQYnmxKoJTr6ReGJk
6XeQlQzbGonjW3+CO9Imy17BNwvaSvaSgrWiklyIZTADnQG/2BoT75550fnQSGKh
KbyhRy3dyiVSWg8cAXBOjpzODEOy7XGzfdvvhTU6iVTXFsxjyVoB84FMjvFKXDTC
ncZ2Sm8qgYczhId83LRdsZ0StDxj0v2fF53Q730RZfAgei38mdroFX5lAMEGfaes
A6ogPw3ST8KOAUKAyLa5paKNW3Pss+TsgkSf73mR1mZMkFoC9Fgq0IdLV4QFpJcK
kcs6EKK2fVryYzLuWkd5lx2BAyEIkXfDjAIRyqWFe2AO3vaUnKrnFH1rZ1VcAWF5
5mKkVZR3/NoPznEi+JtynrqelQd300WWGYSon6+w1l1R/8UqJLlqgYx4NPgXLTTF
oSYVCbqNHpVpopnRh+kzkVkOYDFuIUfrDch612wBntjlIS70W8Plyap+5NRNjQb9
g2oci1Y/zNRdhhyIS9hPRMuk6QN+80PaSftfl8c3W5hzcfPaatA+OhWXImzFrG15
r+BpgJzy2qX7eDJUtnemmyKKlVOEF0gGu8/zWla0OrfJvU62A1+lHngIH7bKzYIQ
cXwI33nf7GkeHucxYPc+EaOtt7nCeKg1ht5tdnf+f8+UizL2oCufqX0sdDwWgXJZ
TcjR0Uc8rCuOObvW5kjJ49xA6SSnaNizRzzInYKDbK5yoVU9yqW1hY954Vhc4rTP
7mfIJWKxny82kNdLkR9VxlkImJWGPAq5eD4rZ62xfW3opDfZlo8LOnP1+z124OWI
A9Z+PCizl0ujatWRv7pARk22ItDisX/BeXihTtRE13IVznmu2KRKnaW/P6QysXjX
dkgxUqcQqe/RYmTjukEhavfZN0/N6SETLSnCgqnJmJXx7fqvDR1KFm13IxVsSasF
ya2COOU0S9gjPgFsjsc39L6dbf6fIFTX4jTo71dWkV/J0cukWxDJmFFpVCB4rxs7
ygRRtz+hxfCVvWO7rIxqqgQPP5iFRPc56ea1tRZoVOnB+8H8sSwRewoIh30QWq86
16GupOn4tjaz0gtPr44kgnrTzv2mJ3Q8ZSINr9b3rBLPdOkHbRqDhSdm/A2AgTsk
GlBLRDTq99g7+DaZbtTRLflY/6hgYuXj34/gJbLqi04yH+q8fgIT9JhDT7EenC4Z
NR4nbg8xBVv80XTjWlIfy1awXDqDHGSYQl32AUHADw4peCsumuhufaOgIDLi+PIh
M5MfWT9ufGD6VzcWUlK9b47gTYszTAw4fTqS8wtHMNVVEHB5S/N+YeajdpbpKYkH
qm2X8YuPMyH6gKhfgPa1ykQXmxPY82iMTSOzRbHGdVw/JXMidmgr4MN+SDvDh0N6
/JTWyfTU2YOx1LlVRtz6FCyGS7NDEm8gFqEXPoXWcfP0SWhgtCehJaNZi/9cXY2i
lTXOzZ5eHvcacw1EDUekfD3IHqI2fuYB166NlJ1I2gsVgMdMhqyM+gIDwifuRTt4
yKu7ZEQUHetd/TdAUHC8nhetMIXDolvfOCkp85pTDbdx7EoDbe1yRKOGYFKb1ntD
3MutPLzbb6n/ouLzOthFNfMt0LJ/xfvsIwjEzWfq8b4kLN/67RcNR/JKWKAY8dR0
9VYB9ubLwNPfeD9NYKzGQpaQGUANpViYUDOG0psLLkEhVgC6IiQw4uoZYR0XdEfH
TtC5zQaN1rzwvGX4FBWXwYlky2ALXdcZZQPvTwj6XZZwSj2A3ZXyS+/IVEfhOsjx
CWgVScSQNs1F1B53EJy+qLETQUo0NbXp09GRK5ROeFSkSav7nuQwolMuKFtsxaV+
oyUWKC7wCougF/600HBuQaP6qrv5eF7qs2M/qt398coua/PX3v8BczM1X4UA9xTq
SbOv1PBc0akLUo08jWFaSom2M8dW6BCstXgJmjyC7xXH5/8FB7K/uU9NlDehxeZC
pLks2eRCqe/TUE7SVi7yll/I2KHBOM2YNHnDPbNFD1HW3AfDPp9vn8XPZzvUsCWP
q62rlX6/AjpR5/cd0fmuF+bLow1VkDX/HHNQDiZnmpyd+MlFBWPYMhufkMy9+I3L
Be1Lqw6KiUyfoLduf09qwvSM1ps7FRRGbL4fSx1xlI/ni9ztgeRqPKXN9poAYabX
H1wFp14F9q9v/i2VRcmzbf1CWKNN653pwq5gZ8ob0+OfhLAWqwizCt6psLNgMtW5
3FJnzUVS1QsgMUQQWl32JNBoDMgIzANTUVPHkTumTFSHa8rnNZDfKeAKuPzmuLBu
22TukPdYxScDFTnKSUbMtaFPJctBDsqHj1lFfp56cXBjat1zBysqtKVPmvJW77li
ag/dG+9m+xuEkU0ILlq7af34K0L9pGFGN7xP1ednHJEBfTfkG5XN+a9xxeDnyihS
1QPkEw8W4/hl0xUUFEc/6NtDP5THdqumWBl0gm/FGKYDetwi6ceOOBkX0zZ4H/bW
5hvBpbGjsOSErSrP6XwsDkY9yHJXn8c51rHGXIDPGjz7r2f+mCSkWUMW0eYsu2DV
6FrNjNhhxqXfT/dyUqXl/j4JGoNLeRZDX7IsbjgPCPatxzMo4F0E3hLHcvGmJ3td
qLY/cZcTWkU4FZI4DqF+yPumBefHRGluq7uiM/LVzcvkKwy2F/ABWVg3jS7uOiz9
3lpS5XaIkMRYOdRcPY17pVLB7pC5/cFnctqKUGcOjn1A9f1JSIC1HBkdZA38QA9A
cQpS3Eu4aMQ/fFFauM87UXBQbAsoiI11W/JTrOOTyzwIumWaQH3e7/T74Hbo106Q
3PYNxuV5intRurYoWBYQzzxi4dtoqJS2fOWRO2uNxpH8JN7fmwH9kCFf+c6B3yxB
HLKfH20b625FSHGqPbiUtTcgF7h0Ma/Af8A6isp1VI/33Rk6cikI4FqxiRcsgPeU
iDiWMWXFp8gV9n1iOedFCKfZzWu69Nvw5cDvd4pVxunb2INTU61zLZ7576jMZPeB
WWsmjCD5twrvHRP02xFW+++nWCMe0L08SzfHaaHcsproKWCZNT1lqMwHdLvgeojR
ZV2EhsxOyY1lffjU6kVxsyBLv5OtheJHFal+QksMWJZz636+kCJHEcLbTuu+8pz1
6Ba7zOV6YNb0nsj1q1njBj4Ctfe6vv0KcVyWUq3vswgKe428xtB+b9W3deFUil6i
UexRbQbL+lVFRhb/GK5EhP1wYreKCdnp5FwkyY3NHn/4HR33e62r08EQhs11o7s8
e3PwqqjjJn8SSA32Mc9BLqrMdV1VYVc4kEQclXYW26sgy+jLjkL5VXTOldOvdVNw
AD6HlgydqG2NM2Y4xjUVLlYjFmQhstUeF5NJA2f5WF4zEJXRL57QjUV9olnzgwCq
Ho+poRKwnKRE1RBo4Iu4fzMp2NrK1GJxcqS9/ky8B+xqWvL0X31h4E9PfWoeM+Ky
DkAznnGU5KqZxdv03PwJ/vV4qFj/5cx7u1dNZQI9H/cdOLoe3ICbMDfQeLlxdOTk
Tkv/wGeU+PNKbynxrWChmdOuyNZ6Jfy2gs0k5orJCev/crI08lAOkCu9hd58MgGV
vougJa3HUGOLRypQEB9YVyLUh2R4TKa34d5wu5gUvWNVDUGPjRJI7t4+CoeTklrJ
1KYt7KBTBG/YtPdOIW4UyDbVsCH69H+RapMTy8YwdNe1kPkVk8ynbbbGCeMM0jXZ
bBNELs3Qs58ArmoHN7/rWz2qwe+SyOZjuJ+4RGXS1a7Ati6Nx/iJ9qTfjdpM6h5Q
UAEQbh+C60hdz+Tei746wS07uHqBB5fwM3QdBE5Fsi469zTqpsbISwgLXU/mpRdW
4Izy1RFXAQA/iM0EnUf0SKyrFIsiXg5NALNvAURg92YyMJ4Sb4quV/eig6KigW0K
tNV4P/Euu6GK04WE2ZslQnPHproS8h5LgL6cly0QKyLeAcIe7pXYBgcVjrMfgXWA
HPs1SZSZl73U/UzeLWVjNHk8f8aq6lFvl4e9KpPnjgyCV945HQSQ7//Wf6MJCDbf
XqKXWANv4YyY2LPg4kcAtGTuHsnF/TW/FVcDrSg8U6svMm0sj4YsssVwQtGnoZDV
Xph2ayzjNRhsUqchTByUISdeOJkxYqO6X11dIaFKAHMIpwPV4T4RSBvrE1mOZYxz
5lABZWQbayKyH1VoaD+2Ufi+uU8bIUWLEEWGxRh7vmt222OnNXG9yeDQD3IClgbI
g8qqBsb7Arkm9lp+PYwP0E6UovbwgkvIZyWQCN2vj8oXfpV4XpPKWWk1PFqIFTpB
U8ao0pYUwjEvANxu30D1+YZVb7T0SrtB3hXkjrslOIx+aGgRhH8mjoXsveJHvpXh
YU1a4L5NjMcWETLST9tTJJcblwYsxjlThsBzE0kGFcRy0x8/zqSJ1L4a/diSblA9
wKmAYPG9rQzyDHFsm8Z2kcrHr0IS4zY+vNZNqQFf8vpfPKaqTp47K6pSBJokCVMP
CM91rw1wo4VGYmDQANc4t0PGoqn67fsm0jPty/vtDeZkxPhqSFKmtuv/5cdps1HI
gTPeFlSA1Z8yoODtHpq/qQWTuh+M5CZWXuUjZjuH2NuyOhDvK66WHux0lmlPK2UH
qs5ahybtClaMcQPTcygcU4AlMj+kWQVqZkYGjpBERUPUVnxRmnb0x+IDdj4nbetv
tfu6e8Zdc/he+xB/g3josewgjyyJbvWSQkbTMSCxJFYqnxDVbcaZFPxbui99jlCX
1ZAR3Z6OvVG61bxIrpL0woaI46osDaR/AApMbMqUBrUlO2TLaVAx0Vg41ymhjkm5
AwYKPHAcRNISzbrLdIqBOcLb1UuREPwADhZavDOGvNxF+LDCzPzW+wZfDJGDJVZe
DUfnNjVl4ST0SDqIuBczfrDLtQiMZZt/fAH4UoEq7uTysIdpxZM8+kzkEZK0Kxk0
vWvS4C0DNP/7SwEmF6dPy6urxL+5wgXOqlPvW0MyMW7Zx18j5udrpqEYh/etopAK
dp8A3XPSyy8mroG1JDahtiPb7rUyUIhzu8su09tc2lkdsZdZYvebskTjNn0waRPx
5Gsps5lGOny8+d5Nf06SC9oRq/6ZnDFxX+U1Md+te2UMr7YyOPqdx6nYZT0pUpTK
QM5UmtTBZ/FvmFzngt4s1/fAAmrM+LC1+XSmwZXIi5gVL7m5pOf3CMpbum6EEhB9
ndvoqWddEItR+DpjRNycqg7n1eB8OwUiYBf1FtmPd7HbUnIeFpD9RkkuJxDZ9PUe
9RygkrB4l4fHYzQW2KGNwqom8d7P3m9cKuQmtJbZ1R8yfYli4SSsexxtfP3WOhvF
LckGmqsmpWny5TIalQjrpAO8z6JT3laCrLBQs4z8TXRzeoVmPhv59PH3+BTy7RPq
AGUlR4UAmuOYBOi5tcHPWCWjT6aEB8khJa1yOazJC0z2Zn0IeaMtsfRl08MZRyWl
NXBCy/Sx1rDTYcLJ6HV8aG0CAC4B1MhlW1qv+DWqWga1TUZ37HjlAHsiwO6nhKEd
+8u6OTG3X35GQ64Iu3sfLN5eegtQJvYnllu9yJUoYn/kZvrP4olCVcgPQKWxiFaK
8eV+HYJPRmgDSGidgAV8GVu1t9GXzqxn+GbOoaP/LOw3sB+QVWFzoJrgf8wA1jwS
10AzrPavsIT9XpXJkDjFPYRCVBRU1N8ZgVuhwje3ProWuz29DD6Nfe7nexoynTTO
sZvNnm0cNWdRjRYOS7zGn0Kk2hIh4Lldq+lTNgDjs+m+TJfoChyrgJ4CjbwCkB7W
2H8OZURJmpP+5oizIj8s0H+fjwS/5KTb+dSysFARpCetJaFukRLjoZj+RvuvaQry
upWKbO8byeMY44n+visQ2+FZr7QqV7rtzSlhja4ZMBr8AgL5YrE0Zij/pCI8uWe9
MhGaIxjp753/C2PLyQAPHTYK+sICoPE7qxsFoWYUnCVqDedgWIF4xpysYSWPhhW3
TpMVxBHvc5m3GXQvX1ZAEKfohCw0oS1O4whik4yCAYPOekFlejE/80nTE85aKA0/
FRtmPOJfSFSRLenuND8CryqpVNY60J3WLkKRCJJZPEAdLU5xLt/G9tWcUG6MrLb4
FRGL8tpTBlvdrjotMqjDwYiPNsT6WpiAbwpR3WlnOKbuQF3bLJBV4vpWn7CrFg9r
MwvNos+vCt1nojyzG3wFnD7BazJ3R7N4Job8kzNxR4kwqGEXP0nnRtxUK1yg4H4W
oWed4XV9ZljIYjARPjyb7tRFxaole8vZH5/JG9bdulvZk4Q3TW+NfwSYwxsoE8iY
YLawvH/KtD4OQtOun6N2ooGM5/3lk0EpoI/IrJP9tGbtkvCXWj5+0FQZt4bZPJrP
wIIhvSENiKdjPFYFSxE8ZkqDuI7wJlWooVY9DslsEJycUveoLHLLhex+Cf3bPY8z
wy8LlU8VOZ8Fag+os2fRUaAO7i1bQHPSNdlNQuXTI5M/JVdgD1UuhXetnSbQGv4K
VMxVuJrgma3LLWv3dDxf0JbXVN2o1n2nuh0GUmsanf3HHt+ak4AcrkoD8GqGLYS3
FrPhoSuvL0ngfSO6yvW21IzH//hzdWmZjAaFp13gncrcBEnzm6UV7aBKfuiDG/rL
4nQ0Fq7qptQxFwhTDOkWR8xgu+v42f4sMc7e/clI9c4VCmrOlg5OX32HUd7WeoZo
vyeN2XqOCGA9CCDxyqa89Udw7mcBKcEWa9KCLebkSWNN1f9TNWLqolgc9oGUDjz9
vISdu9zkHwgRTDUY9B1m7itpplYz1RgiKdniBK1dVvA5odLq53gTCF8ijv1mhY4j
E/IzB7tBjwF68FUILhI2amBZb/nIvzsO9BU8aPI8p14P4K+4un7ToxNUdFwgjimC
2JKnUb5+1dWMfMD3APgZHBsZ4Wi/h7iajmSi7FqX+3+kpASR/8roJWPz84qXvauN
K1nS1lXY6OxBdYbdMDWr9e4Yfum9h2q/x71dXesP/4G45RsT3XmG0tkmEU5QS1Do
K7ldasyImx36XKkxwiT/rBmEc2PAd2MpRnmrOiAM4GK8UNw/taG4P5twIgwqw/Ni
Ckl43ZQ8b60XZmst5nsNeGC75Mm5QebNfDrzKnBUmCz3jf4EFNpxSt1n4BV4zyRx
/OLBaPETMniYzvTGSf30rt9uqMdhDpzquND4Qkltl2OouKHu2Cm3Xs0TuMXVcLyS
i9RFDE0tvFw3VcK4ywPSczIHpUZ4Y+IhGabvZqvX63Y2TPxsnpTgv7ZsIAjYCoeE
iJ0OWKDG6wTioxxyORtqrI4VSzH4thcsEP0RH9ScNG+/7BFBUsI+IelpaJ8QuYcU
PRfIIbhfQZRsgRmDrmqQX2ii5WfdzQjHpUr70rG8t7RZ1OktrzQDlcfnuxy/7NCr
q+m6MVGGaBg/px3epelhVfYibONnBH8umA/Y4dOYnekeLDosQztHW1Ax5SlyShEB
pBMJoDvQt4f4ScKjEReHGfa3L13JSo1MJjK4sUss/940SEGO1wm9hk4L8LS+1ECs
1QOEuSpdb2Znz67EN4olOHbIogsIGN4YzRMX3hU6f2bygcP9GTQxLB5h5NIMz62g
n3/iylKZc5X51RfL0o0AHuco8xgsi3gvJ8esFLqF7lkFJ161SzVwCxQFKcc4JGzM
q1nAjqDwNhGhOylA91gOykxl5KZpjXoyZJDqwkuzmxJFV6bkgo3Qp2jrfD1uA1Ui
a6XsT4lUBf07owPgTdHINpqKeCrPZZscP4K1AuSRMXb8q1ufQImSgenSYc6C35Gl
TmU7BkaxyO7cH2REbcnyxHbSHNQvmlcTMcJGRG8qdrQDsFWCnBtYJ2Zxt1bPmXAs
Oe+acdJkQAIrxW0VD0MVQUKt5PMRvve/jwv6yBka8HoEyl0LIkyG5LAVyHYvTQTU
QflmdxO3pegzx4hzYFLlp1hhEkcPzyroz7VmgKPIRavexsYocggACA7t3MYzx7MC
AoQ2b+d/ErOzbXaCKeFTYxPN8BLnAW2uJKa1fmonnWj4pIbMW6LXIeuIHun83hNK
c73KEFuZvmWpE0Rp+FbAOTF91e+1W9MP6MwPqvJjofQBiL/TZ73IyKAxV6wLJZ1E
JYX6QXakCkG0DWBS123WHf6b8QzNJY3c9Gcr2EFqHaLrtZQnJX24gm3dB7IH2jnM
xE/roHnFCPvFw2JCMrG+3ML2/QtEvY8NYEcyndBcLcCHf31FF88EKsROUmmXGLVL
V0qITU0YqlnUaVHeV/zfsBn+ZicXg8b1pFHkDLAdcqUcwIFp7W1Uus3zbuUv/8Yk
BgEXoyPS6L90CQHlur6FIo/vLY6+Tca8yZJPg+ICm6urZuPw03N+ix+aEedWHfUk
OMOJNCYNAxP+HEbvIlHhSP1Thu6r9zHXItwQSpIPcz5cuifG7ztYbMkp6umqAUJ9
2YD6v66CreBGLpNEYQHr0N/JBEkkwJfbpdLgqp+jBMLvn5lHWwKnY6EOK+qpcNSs
nLAakSfKGxEKBv59/eLlXuxEAg8kiT6qN30y1FyjQepi6mVuuQ0CKp0DZjNc47Be
/4BLqzWwNzB83vVYGD0LjaBpX+3pbxxDWoLVOMGvnK9QquYnhvW56vD7YUTkO5yE
nxJaPXGsfb818hkcrb6ChmOYubs9ZpOdvtI8CLhHAqrsy3+3+e4t++TfX159PKZA
BKEZcR54V+ttQbXh25iKMMoLI2c5HeTtNvM2uxbr7GOrLGsGhHqRzUKNK4Q5z7G+
tp0AKG476x3gPUp8rsWloKJPzKbnCndvukWQO6SBLycUE96Uvx21J071U/utSXu7
PXHNQhYFBDOZQvHvyrjmlew8dAbRson4Fi0d0RF7jA8XCtJTMmbn+/bXH7Fw236k
ED/az8Srgm5a0Hsgn0gVDJbEeNr99KYNWgnFj23MlUhbiyonvz+GCxAFpJzjpMVA
9+CC7UrInrHx3lUC2zXdCusAUzxn1NuJSGdR6JJaUaKlKAsxd5ymDAWggJsxscRN
xuUCtuu01sfpxjlJL50/yTp2Fh/eMnacm88BFP4aa8C1EW5ow6WHMOl4sqyNnSiY
da3QTVAPd+VZJHC3sVp+R3/1mNQAWgEN4w1NyrA7+mgSTWfil/tbBxvicV6x47HR
jfAUjVBOlBcIjvmjL1/fHcVd3Ta8z2sLBtXo/bIxfByyLw+XEYclVZMpuYi0C1XU
TiI0DI8r1EBDavuC9cBMeG+PB9zIvim1uUIyCcq+bDE4xMaen9mty9zZvq76vlje
Qchoz/TW3hiKVat0w92b7NrpqyKgP5Pe7aOey3MJFaCNJjKUM55KrGr+IlpkPFTA
Bslcq0oUYUBtyn+3N+FIRRZiSlOnwiQgbHo5QqQMuFnxmWhp/kvQUlzqBOA7/b3K
DrEPvmOBqW3UKxutSmz/eRLX/TOtS0Fuz8xRwUE6+0t5gN22y0xLdF9YCTdm9wgU
C02OJ89ytOjc1zTil9bN7dUUqfueerL7kI8Dsk0AuXEHLJV6EglkBwUOvwIgDhXK
F2g/dEIvf3yrh1U6kw1wivo8COjNIxDjpUy6M9nw2TH8hZ4yJXVBEdSQa7MrRq6K
wweQasL9vtQg7NAjOOghZzgUdCxT7p4QjJRArzYbaxKQfjzZgwd7N5eZw0h+8kFa
t9YTDmRH+BPBwE4nqmST4EuV0NZ4f5RvAdwHVAdoaYm1LpJUbKmnYxznA2MMn60q
gUBazpOa3kUG5HLwDV6PZKu7OljjGCr21HapQsBGCcuGxzOtALyRtsDA1O2PB7ZE
oTcvrKisC+67jVx64F6T4i33RtR5b4lq1gz2THePcSKcGjAze3ElTVVacLQyVbOX
eFc2guPwvm/gyQK07Azg0b3OXzL08txxvHRnVTJTcmKP8NBV7xy4CzeYpd7sWnu5
8spzL3Ohib3hEHuWr0LOEvTNegiCLkbkvc0ChFhHzNG1pSU75+hRfoE9wnzQrEW6
w8vS5ePqH4Ua83V/2jkEQR5kP57g53j87xlR/TDxvtrBckIt148Ex3KqnJ0K5M0s
Rw8jpxsBLC6PMCJN4m4Tu7m5+J4VfdCWkYIsBs9i5OARNOkm+l+ShOReMNMVnEJl
SYwN7es8I1i5n4NLNUZJhM0AcKl49Pk/cD5fl/AbWw+Fe5bRr0xK8EAY+ggCHji3
fDKZRiDdgo1mCZotIaMz6ignIiZmFdjBljvF+hlA1gFxk0kp0TL62r+4ecfGlCXa
CJq4Cu15n6JD+CbUP9Swi5kCUByZB+DAyPnKsnAkQn02uHKeG5TJX+zDmpDQZ0sO
nOqShvKYXvLM2V00OZYoqKxkR76QNTUMhB8a3W+m6LoK86LM9O6Y8EDMPMbpHkll
PNjf83rtzEocAE7e7rpTLS3IcPFOMm0NBviKG1fMwt7/MDVXNuLaS1c3wElvfAf5
Bws6zXn1lvJtvjFSgoyTisI6CTno3/aNkPsJ9coRw0X3CCM493dehQaiMZZADoL7
JTKzZaFPJAMv/N4lG/3OsZ3GBfu3sne00xEeSGzY0mS/qdJ3dOvqJ+qDcnYykRuo
g2UOJ/fyTAAGkOzuzhXTeGoVE7PIgvWuw4LQE56NQrmmivvgUS7Ml9IpPLTowam3
DBpwcge4ZSP5Aeu/35NpEtMn636HMXhsyUr3/Joz6VdbgrFdskhjGqG7VYVCnzbd
K9cld2XdVXyHu6sVNC8NeEo7bb8oYCl8cum2b1CF/8T9qgOJgNQCq7KeYuktfXlQ
WswwmJqJYrbktroDwr3oMWIiYeCGOsWX75Ps7/W/UiDaRmjBpbY4/lKkZ6lnxVGN
er9xJsWfe9Xx2iTsTmibQs9gthJ8Gnwf3gf4u9LMexMyd41dZ7aGu70+rIkTcHBy
iAbBVBcAWbqQW1wyVGNE5QblbyuGsR0rCzH0x7WK/FdouBpQK+5HbgLum6DCTa9n
yDEVgdKDhKAoRpGfG8bNMOoC9g7Q13mnS6z85wtxivPp+hd2E1nbu+qJ6CUEhrh8
qdzBipG1w4zSaqGuU/S/XSCAlKZkXzVWJVV+kjCfw8gURiC9g4hwsKfQW3TuA29t
fUqhTiWfJpzGimE3gdbAC3xbn8TCXtr1FMvgv0ljuYdw0Iyqt0VlYSts3C2BUrlI
UaXNAtB+v08puKc/tr1YjBtiLzbnGdvyxHg/jgFYxYWVPXeqDDN7ZBFub5L712rP
gkIGb+hizGslgld1ir5oA4IMrOCezvJ3mafa9nUz6ZqBAK42Qz2tmsYFHbJeBvAj
u9142gXhSHqeBUCdw39fOhCU3o32Syq7rl2kO0jw25TnAaodQvqacMFqfbNGz9r5
Vh7H5kYgnjn4e+dv1Hbs7iBsCmF0I2iUNAQCEzPNGf5R/ffTc1QbBg07/rKsuIqF
l+CCvUoc1wzy4HQNTrDl5JDEC2ymFLTWmBnchbTEOMZLt+PtITYLF2E32cLPmajf
W34oa2nVMd8WelsrG4Qf5937tdCNC1tMFmLtUyNyTw8q9FiuMrBWzmH4S8Zh8HXi
aVYBd5/rMEp42OiwdMbFTCUbG1p6QK1jhoxL2qCdZtm0NrKp/Bn8d9c7iiBw7AR3
1D1RZm/BuDiWKZjexe0VaqQaoaF6UIvUVKn26I9+4Zi10F273gpYuPM39V9RoaPx
q28/hWKH11SQMPfImYNHsDN1xi/wIXrZkFO6uxPMdO+clHnvGzL6cLyrUaBs1Znm
AS/3FtS/MyAzzZzNpvJULjMye2Rbbov5in+xzjba/zcF6YoEI+nf3PD8mu+41V8s
9X+ewFhHVIc1R/2MD4c3VSroH+DkkhWGiDfij5kzFNmw/+MBFAeYBcS9+CQxjcT4
ia40XBPEbLkpJ0ccRe/EMim86kS6NTKR7Sy4jWyBNWr9IKr0ZM4Xy1yhP2XVmiuB
6a0BDIXo8VgYvGp5TFJWIh3xiC6Xp2AFxqb2YIlZDjjQ3KurOqrbQBJr700eJSLd
BFSrr2sG5uUhQ/eCcYFCAfnsd+MRmneKVbmWSJcze21Bm4z+EpV2yuAjEw7JewXl
1P5Vd4zbNFvPq2oUUo0co/ckq+9j9IZ8jxZxBcPYKezwyZruvgK8nqsrMcERGSYf
De/1v7GntgKdCMjqq39t5Q3KI+ZDGH6bg7WwBYUUQhmPYwiORftqWJfYjVovVSxA
Mg53pEAeyQr+/zKYkmkjuYCA38S3OpMecwauZmgKXO4BSt0gWo0zDzcUVxUXZC4s
z3R4orE89/Pw38nNjDFe6wj3e1txEU7HKk5gFlnGnf0o+3NKaVDnZrc7gIASfTu0
TtOoqsGkSDa+yat05tK9b5CjJUu4uBhW+rg1MTmLgxDzX03KDdAvYEl0NMwwLO8f
UXq6NA0RuiHQGPBHu+UaoR1W1xdbuwYC1NSdpVZ7ON/TZCGJ82OBaJrDiu7QK9x9
Qe+TgVFkfuzqe+46nsqF/l2VLSebbB2LJewlIJ+w1dg199JNKBXcTHsaksNAlv4x
bjxL36jHSDOgurNhGUVFOsI6av0jSvCQLMbE1Q6u2wJ1xBVw81Zjixs6H//YSoD+
uzxhN+rbg1nS8YMMZWOYMSRa9Jf9CTfKPt7QkGCbgkAl5NBCXxU6fK8F5CphCAsJ
MTr4MPEDpQ9eIJ+F1Tjy+ZVOJ8tJBs5K/rrBll0xEp6K9Y4CAfMnyr2Ord1K0k+0
GgxALcZLRVeHLMp+WCyCirAEJplaiNQPiIkxumE0C3qZdNidKSdVYFC8HVvNDNPX
82R8e2pWdIQU5Bg7uuZywLPTFQn+zJtXAO+Iexk5UhCBTyWgI+qOKdHxHGBI5dJK
KepqVyWjT/CjFQWN5qaAi2lWURAvIaeTTf3IvhtPtEXp2s7cPc5VT/oTd0E1Zqqe
U/9meviYRQFp1d4CTwH3cBQsHHwmcaODn3n3FlB2IPXMefelE5LLeIiLnFA/xJco
GWbFHRHKLCr6ELLYx2G27Xk0/syCdVMM2kH59bshiOr8tuco9xDeYimchb6cJWEl
Hf3+x/eF8ig13GkYpBaSVOXkGfZPevTEKMHBp6XM+CV5wZqs4qucq4Sccdsmcdap
h8ceZDQc2NuU5dVSXiLrwWp4iCYXb5Q1ol1a/Uyc3Wy2D9PIe4btcK5MVTiyKlzY
xZmaFz41S2tllwCYZ7Ipebbep5VwEPhVku1AyPBooSQjdyJNh5gLIyx9HJY4h541
YaWvYD7f+dKasCiJkSsZN8Jc+oA3XIaM9VX/h66Ap1ACKNFMGur92M616GByNLvg
XP3KXg1J3cLHygP8VuacPE9t/Rdlb2tAd7XqPsVtb7rkF9tHhk+KGsxRF3UBk2Xg
qfz2jVM5P56LbNSFzG160z9g0uTMW6ZayIk+EonfNk40HRRr01DJYgxb8Lh8XN/1
KnOU3OxdJGkNzz+W0H6bNjjozD+uCjXq2Nun7DWxZxz9EBIzctBznP9Eibcxe6Q8
Xyc1zsUXc0tSFIkHuwiEXVJGycDjb0W85u3MDxn94FQ/m+TJUDbpRe1EnK0QZqcv
28re0hva2eV7tXUxLkNO1N/y1I4se/qbbYdM1rwywZBxNwJ4Rz/rlEmLIKgkCtm0
SQFCC95kWni33D5yFGdSl0BixgE3em2AMho34EWLBTumCYszx5rS5L/SIK8hnuQs
u6X95S/9RpK9a9K62nAkdEj71MrPfpWAVIrfkVvSYMea+/Xx5H/cPDUDG4XRi1MF
6+if2GgLKncqTjonj+t2yD4KNdEOq8A8rmz0kg8Z/tDq50uLPhyfKadggJj0cnc8
vpjafYpEoSZ57cDMsqMMSNqc9y/WfGiZYAamRDENxL146xgv9CE2P/Np3Z2s6261
2ec5fZW2hdYdlvoMWRmUM47HZsUK+D5hL3RLvX1zytUeZ7kT4fOTAtCacw73R09Y
eIEEiGap9Uac+ews1k3Yu/qV+84VV9Ncoy7BfGCZDM6qytrW97lUhy0mHj/5goGe
Bs3CMHqLFBoM3ml0ymfYEvWe2314H0nB7xpu4hrTlAxfvYC61OlIq6EJlmqP+/fF
UKby7AbgfXZhN1Utq0nqelk101BbvVlHPo/BSrBdVPjzrQEEORdf/1/ONHmEIZl3
WzviNcra5CgZJNgwYkG//Gc3mWAOhz+U6mcPn7cjGFaZFwblfGxIHqh8FV+s44GX
kPTBnaCZDHNHD/SMzM56zCb4AxCuomDY4DRg1wGlrVaJ7WxShSxRBjZfpcQD8Rrh
vJUXayrsIGaawECrJnZ2wK2Ov40+8VlI3Vrgwi8SwNlwHlBDxU0/+FEhxtwxoHhN
5HtHBxkn7+LPqDBPeO1kb/5oGppsBTTEaHB1i55EvGheqUAuN1L0BQuTnLLJjGTp
l1pKKPOpHJsKsil89pA9pjvaCxbkwThF3QOlPTNWFTDsWS8X6mPLGLkZUl2CObye
0H1PSj5azpbeKfRE6ZshKcG55F3dFOnzwHouQjxSAqGvFZ4zfpugejSt2VrNvJW5
2UZArnf5LkQb2uRNBrnhiiRG/SKX0PeQxk3KH3DOwsKVtxR4ch/JuanhbyhrfM2m
p6JMmthE4VBnvaTYtWwl5sGOjw90bEcV4/UwChwe/CAV1keH8VerZHcnkVjZ6fnc
nHvayodqBARct0kHd1NRJZuaKsShWkYMJawMKJxb5G3A+O7dKc5tv7/fQ6mQrn8C
yuLRokRAnVJvbeR/lu0yH6JwsgfLybXfqCaFzqB3vnd59s6gBGenv6Euz9Ep7Y1S
xoJYXHPWn2ti1IlcZ8LaI7WFoNMejA10HxBv0pUTSMUYK1gvynjTv/cAL949eQZ3
lA7qyy67uqJHwsRUGCRNxVlF4NPEA551+cDCwlz4OWA7PDa3e5rE1y17ry/FPrK7
sYLNy5ulYXuslPfcxPoGrW2wGKNpZWiJJ4UXNNbQwTqlOJTEC12UCKgnUqLq8MOf
0JdIP+58FzULPnR9bPpt/N9t6FuqEsPSbqMNfAQgp70wnKciuD8bNMoTeFXy3sGa
a6l2hq3DXJM3waz70zf9YLSeyxzK8S32OOvAaF7MoxCJyJRL9jtRlmzdHe4SSShf
zdqpTSdEJNO84FxNaf/vps404eunocrakWRq0tP7JpJFrcs2uGogXCJYBS2SCOhd
koJkbrYXxd8e4fMwK8Rr1enpcPUTfFP7DEOzqSizt3VJU/5AizfIs6jvoy5gaiTi
pNge1N8YJ7d07rFClX3L3jMXgpEavkrTrenzEaKVr2NWFEgu+EvTJpJNMhd+8wsl
msZAcwjXQ1ID7z+S8nbXmzSLLthckNXnT//qTJYQO4apJWDiY2oZiSUyA4oaIsGr
JjE+lxTyTcnWpExsseug2xzWBeKdO9LrycaiayuZWeHXwwctJi0fIr26JEXA4d2n
4YY2FlvYXJYxsjdgdNPWY5K9ZfyfPTEi7SfeDBRvMn3WR+GFZjoijtqD7OCfRn0N
1Iz3pZ03l+4dNpv9OcZaqVXpdx/vejILCceNI14D+rMsxIHtH46Vcz59ZA+Hw6qg
jKjSU1RrpvhafhIMFqjk90Eu6S8Nhv6MnouHsF6OyPpeXB3PEfBNnUzuUHUKVA4v
7V/VDZErSyYyjFW/EhCb+Lu4CtZJkNRb2henJ6EYXZTyTqMPBB6usd/wGv72oTej
Fbt+eEYcYzeapKq4OiQOV3ZbtaYRIitNXCw2kp4Wct4yiB1iBBPrPAMz0H6mBAxw
5/LedhcM8V/c2EkB7xnPFGBtdJa3fvEBAE3IK4ssskeK+NSIovaMIn3G5hf2bNuN
Atw8YpHGkyhY6pFn5/0HHuXWZGaz5yQ98LuHUt/mJ7Q/gmILfih+EKcX3XRALrei
s/klnd7ksYUmlncTUEA+KVr67zXTY1PA7ZMo54nFSnI+ag3Wb61B6QcKC5ySrV08
n5P7f2Epqw1UbuEm+cJ98Qi9TeEWIAi9/YdIiiFfHy3tRa3QkUNCxnAuqB8DCOVV
uwI+uLTCnnNw8G9b701nAtZe3jyhpwsa/tseQNXm65ep04iqkc9ofOhL+bzCDZ97
2TuluVXyKmy12BMonrtTgsancYdLMssSFW8xC1WW2Q/FMx+Jvc6xkfdUwVB5JJ9U
5h4g7dWp+/OJMid6R7TzXoBELKJ3xB8P9rYeof3b9hu6NNQHbIXYDvFO4/eHdI/o
EHyVX7qQIZaMZE35F6/TYGIvekIGIWVUA8DN7uVv+vUu4pnW7BP+FU+JbmiSUouQ
bT0bPb8CMTTTfLaVqLMqqbvuCwyc31B2Z9S/ro7qYTdwICg69kbb7JhQtoKNcdPL
hhBl/o2fEqaafqvxCjx5PvhQqxnXRzRJEf8M9O7VZUvb2Tagi95PhT4XN6vkbM8a
v8hqdVBCtKSQErRanUcD84Kd4fWelaAHbb8660P870ZgomqXJdQpR/0mZZEwWiZ1
7chCHEmzd/pXnllgXqWvOHoAvCcvzj+DKjuGesJ9n6znBwPz8TORQKx7OaSb2zC0
TpNaG+evkkucdcb7gEYNS8YGfp3YsYqy1XPaAWwCsne0Xokw1zTDed+9903l/RGR
ld0Zl8oi6C3ETtPqBuMY0r5KjskE2Tpf0YfI+nBouxZa8ambYej7fbo6kcCKfXOE
nzCxDNbhAw9S/7zCoa9XQGbHsw6DIQMAc6m+/rSwntzqU0n9uCcBBTpf5aRK1l46
F+wA0X8u8W/Ih6c21+6Dl0/p3SuxjuyUDkFA24ms6DugKcbSFkK9H5Xo95LQMRy2
++3AsJW0o9VcnnPzl+nvpgztGCrLzkwQkepW69BY4jHQMikB+EIc8QEaGj6ehrPs
5MarIePLqlSPfh4Px76zkyO2pa9lw0vzYsnULOp9vD9OfdUN+02UJ24ISataXXvf
nTCUkwZB9Im+pVpepjufzkWtVr1Eta1XPNso5Fm1SnsS96FNvHYs9gmKKUOIokEr
W05HHIggV6I+ym6QRda0UNIxzM2rMUnMtJbYUT1z3KV0mTz0X/OH3mYUu7FGOecS
q5W8v4ZVHvAaAdvY4rNkT2pXovpZ/e6ggFUvA2xrlEjQH2IrzF5Uuy9GPZpRDNau
UPPZXdCJsjXZgQu18Hu9XhBU45hH1Gr21q90ZeYESiDcWdgRgeg1ilVTY3SVahcR
+kC1+hi04Xqrfh0/WrA25SymwEhU6korSgFHs1ChlTIcg1GdLf+Y8w/jWp1lqU+t
jK+hDEn/pFo+dDt97WWU3KQMtfufYpIJji+/V0yEsld9TroRE9NDL2F5gn6GcCUp
MhnpxWuagAeD+8JNdIyCQ4LAFIT+J9LVKy4MBRjSiTnwkeC3IWavoc/6No2L37iW
j46+Y7uIYWg4V+YEsIIt4weLI2VePBMXqGAuHgyeXJlFffGqlSvBQ9VpHPpyFcGf
PNAB0YAB5yLUCHZ+krk8/7isjh1sFJmhD9BBDXf98QttP7tcWTFZ8Nq3UQsTyd3D
QF74+VD7/2bWchHcE5kRNS0n1OGTWi8Ov9DSbW4ToRqCOmMD4SD4VJMScRfUx6l/
tHlwCVNpV4H/U9LkLpIgYKzTzfywncR7QaditKx4M8Id8megrYepVoiNUsm4hudx
xvRj4ApmTVLqpE0KCYBzANMt8fJsGkk8bk9I4ejG7b6kHZDTwV7W6RxqQUSLmdW2
zVqrGGVmhpG2Ta4xKVb+f4fULj2P1K6TLj+dcfSdhWqdzYlcQJQY4R24/zIq1uT1
0C5c6DuclA9YmMKADoPEEROg3S8ACELVWkCF8ETc351jAuWC6/nFLFMgMg0tV6G9
w3+opdJCMMidbDbX08Bek8SKsWaU96rfIJMiGVRcDzCx9GCCwkJaFwK7YIcTFSJv
gUNXZDaT0m/FkvYmadHwy0O2KI1cGlRjXX8+7Iz0kz49uViypXeSs8/M32uazlBx
tUNjouTM2wFfbTFumiK4UIWxJuTkQQ+A3F8PHapoMF28x5xsfhakS18IbC4Ul8Un
jN+WsCOScBWdVZsw5B2Lc43sJH3Z5I2jrMPJQm5KeqRyLILfEvKu1q++xloS6Q5B
RzSRQQ/FvqsbJ5YvmNjYhqTrWRjTOm43OQGVGYYz5v2qX8pqEDHDjz1onumnY4/2
rRx9edM2tz1je6Ickz4ZJcfkPZeSjiG787lNG/7rQWS2lmxR5s5oT4ii+BCtKtg+
IPWvsznUqCj2H1AipoZtHGpDagltkvn0VDSam5/NRETB+gmWwuvEktnHkHrqp4qk
mF/2ScmoJKgcfsh0hWLY11rmgW0RfTWrW8yGURkHrSKgdKVJL0TSGFB/RegOyKRQ
/wEy/e/hpOlx3sZ5hikZ5eLCKXbS5ljwMNNyrTnGgezSS8v1NH5hzMOWAARdSBS0
YK79kLap4sDHbzloQ7uRLxl1X7v0sBSZTdp3vTdRF5iHvAhE+ke0Y1QZTj2mxHYe
gGb4PMbThgxmKnf9gkFOx6Gdn8eqWr+MLvrWWa8HJFZG13gq608mYiQ9JVlHQdPa
jJs2Zn40AZt9TIj3sj5vGRETDjVa3QrbfTqP9aDdUhB7rRBdjOQquYLrlQLMdIY9
Ic4VQJ/lAv/nkquUkc63gQJ7EW+YANlZwzXwxTczg3Cp2WPshhAtJ7AFAbt0hn8H
/JUbtkxYBYAM1EDPEvhRHufPuWZux9jn2WHwT9fuEHTRvxfZrS6u6LRBG8FbHTG8
XrHwHeMoN2twJspfm39SXKUxSuLNsLCGYvEkmX53DtCPRaN6L/3oxJ4PNi1StmM9
iLpzb+7gnL54EeF9ZnZ9mmuOVmKfjClt2SLWv7K8v0CfPHO6ZyJIi6tkox7hIqAo
6tkUtRbie9YYtGHrgBLRGmoGLq2HnxJvBIeCOtE22jNG38kfj8GNPetU+b8TbN2Q
Ge+Dcb8PgxRi1Q9Sn8hU9+I6EIHUFPOoOA3XIWNkC5c4mRrEQhCoN/Bvihi/hlMG
E+QLr8cCURtMoH23EdQpl573zswbOlvjbRvb8pCNfgefW2KAE5sSERivN1l89BYh
hnr1HulIS84NBviJ6NhAIz8lLQIyABQxE50b5gq+ZXtXq4fX2BSbXuJeKmu7BA8M
DCWmCJUP0FOH0MgsMp2JxhurlmPya2OaFf+umVUZvhsO3TUCBVq/DmYgdzmlXhAj
jAqkgWG02wzOPRf3q9ieaW2b7ME/mAezkkKBziBtNba3tRp1oRQ0Kr80Wvwp1xAA
Nu4FEipmIsUTQXTwh0+3cku3z5bNyFVpTMC5okTA1JuzYlGfXSp52eTtkJv0kwnQ
azynLuALWqriYhH2NqplPHed43OikeSeEG6mCB8uovwigdap4kKVCK7nhFuyptsN
pdCs1WHnU+CzAvEMCtJoG9BaDU6y0+Z16/nd0hdbk0NnsHLCwg0EAKIaNUnLDHpp
u9uhx0hJiwO3JptDcYHwXh9G8qt7pCe1AfhdoPZUGU+YMzq9hT1ZhVn2rubuAe06
pFEYJDoK+y8wT3lgqucqNWPTlQJJeVHyyp3wSQIfq4brYZ9AIc55ZsikS4GY+beQ
In19oNs2Sezw1Q7qvNYBDx62vLJGsEkl3lKvtyE10MoeYd6RhUjDBYG9MBZ0EFL0
eeohjwRc11rt9ERgorP3HF8NT4d6DOXiRrSPViD7Se9bh9f0uicbRAPXwppTrp9W
MDgNF7Xqy8IS96cXpHTETAfHrji4gtaCrnlmT3/hKk/3rYItGTQDKRS4bFcZiCAJ
ylGvN7vzsqV4L2s0liXoK+KsTT3A0PaCyoLkf4MMsx76myvauCRqXgJa7kquQ0WD
/LORF+qXShxql0ooVerahSQCMDjj5TIn8ib3piE/ZtF+Wwr4nLPogbgHguKiAQKa
xOkqKLFc8on5SN46Asoo5cRAPtdtCguTCSVOBBEQsXXn6S0BpjPcGX1C7l01vInm
NyMHJgOXBWhW/srSnJ3TNPX4qrXxThbYznJgO3+phRkj79/6wv8KUmb6wqUyZCGu
XnimbqgyIKrZh2AjZiSYfvVtsy0e0zsCr5j7d+hgvs1fKSTZ6CotQy6nTN87B5Rf
Rd7OIXopRdGq36fYwuUfMEwrbgvIPNCPlg+RYgYB09qcinHuQ3BbzTK90eY/LcUP
GuU43NtPT8iPR3U/2SczdsdNfdQdpWMXMK+WK3v0WN4c7RfeG10jnJrtLWYWya9b
xSVByqCIsB9M4Gxx4sbCxLfO86/ZBMzf9yrCSETYgeQElDzlonm6hXCH6JiUoOKt
3Q1E/WakfhC6tPSWqf1bt8A2FEpV5Za1JuAw/0qrnfoJ02XGvIC5+/k5gQ7Es4Cl
fXRRdUlrPqi1ErvnHYXebcv5S4uxGS0elOasE6mvJezXSQXmAjMQ72cbCJxT+lg1
DgfEgfeWAKp1PFhDoumV5Z3s4L/2Hlc0vpiB3PZfMXRsFuiv7MccyNFzAAxjxD/d
bqvhELxnomxrzQPmaTJ2fs34utZhvo+gPAUwDMZrlaaMJKSMWQG/qobShIjOdh6T
EFYv25SaFpBjUnRsAqUKN7dymOF6dGob5Agh+YfZtk7aYNovwidMFbfNxi3eycVm
9Qx+8nvGrRsIYbQzwJ+e+Y/NAMCjt0q27i+HLGKYZ+DVG+rzBoT3dtzMGKKBYbcO
kE1Oajegt/01pTG6nyjMDWlFzpqUkzPcdex7QRf+Mp8voheD9fAv2KIy/6eIsbrn
LMBJ/pF+8wb99EDDdUXGFipPR83+CfF0yisllw7CjpsOYsHtXcDiqlTURQ0KybF+
uDJlrDUcL3gE+oGy/l9B74bSVKCIXn+emZmSVNQyEDgJIDM2PFy8Y7JuQIWFrtj6
ok+OqALw8fljmIx14S6eW9dgGf/bvLEKi0XMSIZLAHIHzFv8NVBL+Tx58iGZ7Ls4
5hY4JYsCcXDot9HmSiu6+4S1pgAiaDR/eT8oLWfDs7VAR5ZrDodifPtb/B/ixrhR
ZuZTcw1zzD+ffMwkpknNZOqHAiIQ4vXLV8jX4wmeAGvEp+7IaWOqOzXoYea/49JH
UXYLNL1G9cOWyEZ/34lBwoUbI3/F5gZo1FsdNEID2klQreOvTvScRqHIVnB7dbyy
lKFSbw0hLxq6coEsgFs3TiOO1yJ80I4R269Vq1Ao/vOxzgH2sVvgvS+G+/xOQiQS
ByU+Nv7YnAcszHVjYEmD3WDmJAh69m40z+fvaNwaBn9Ju3eG9BoDYdq5cQXziN6/
jvAI+ohFx7cYCkm0t6Q+Y5Cj7vY/w71TQ4ynyiiBqHmV3ZFz2QrHHCzCWoEUoW0M
PrZASaSTP2enmbGP6dM48fP4ubG7954HwmKvw3n1RGAYrSIXSLFFkq0FeOKw/5XM
k7dsONKnk+M0z0/7fLo+hFnp2kSD7QRzLnxEly4SmXgpuQFWZhTFfmrIS+b4Phk2
XDLu0BcEYoF+KWvKYV/lDy/2XJqre/0rVDNeUAy198xXQOsAlXe+yJPEQKMED3fk
BqvCbO3uaLESTTZF8WJcrM2XX0uWrcPxBZ66XymMWURdHK+hblwktEnGEllIJFJp
Ee2Uz+jZ2sEZcX10tUt7QmS/jtmqlD4H9CWZvho47FXzVksjJffuydEgd2v4chG7
e1YWWrQ7ohBwYC2jGQjiZ5cgqp+CzYZyRrkeeKHICoje3EPyULCpRYLSqX0rJh3M
G9sF9Rocd7uWheMaa6MDvbWjCAMH9DaGQxvUE6PQsmZAbsWg7a7ea71Iqf3b5wMi
7zl43/JndcOOUMpDWMYE2qavaE7mDOkd7+P0B39OgiZ+9Q2nL/tfKoXt7BSayYxd
agvI4jJUaVwCAKkcSJHrZm1oxVlXy+vxaOevYudvdTxHWcKvVvyInf7OHhwDbQ5F
RATgWrJbzqiGDi739mton3T+qeRh1bFSG59EwuXc7HLrXlUKxjK50W3bgtq7uQgc
OkILki3YK5R5vl6Kix5D+/Fh9McjX1cij3Q3lXNi4Z3cDVqk9Y3iAtAecmfNmVBR
MRdCOWp8hZXUIDP31lGMsi8olHYo+fmQ41ML9yoNo3Vx8pgaY1zsQps5nuqSasDc
VnFctrxtrA09OouDmqkAtc4JLzFi9gjnMIyDDYvLY6pYczhzGUNViVjsf9kL28Nz
+TolZ4f7220xq5rMBHN6aZ6X7lpjILryaYTAJBqC7yK+sz/9jBPHoNDMbeuNBc4v
hfyBYPRbJJy3XTtcvyXUJ6t3Mmy1ESMh+JLgMo9HrN8SmrERiiediYWcnfp8W23L
+V3StAwa78vN+PDJDXOG6kP/FAP358LZlCxwK9zYZ2j743RP3uDUkIp7AdAYxMGD
uWT5JQzzh6ikRNLN49fyoFVPAutFavauRkMz4BN1I0J5W0tVLv7XGgc4+4Zbbrxu
g7Hp6Q9AlynwQpMwzGEk/ZVQk6OBYotRstJCIwEitjCMQKSwbmM5CJ+aW1/1ZGlK
euBLqHJlv6KyMIDuitEWdqTxFD8fHLqAfr3JG8FA1tqekIOOvyxnx209NrNmu6SF
R5yfxQdq2jXrVCShsOxqlEC1W4jI/YIugMA8UZ4ATH9QN4+7LF25YXQO4pTdS/4g
ObjP/vQl2kqJhznmJRzaixvdvpNPezspYnHwwsEx/nz7C+aMoUKVjjF/HZY7ES2C
rFFNqgvB+bvD+7JnnaH5IkrLVXicTFJ4zPskaNtxaeDiD7yxoMCily8k+yoigEwm
h4puiZI++8zyhpBhynZeoMipCHlVWEXqr+JJ6sv+sYZypDC88iOY1d7kKBBxsjg8
0bbAm4e+UayySSeI9JRlocXdrz0ZT+gc4HzUaYNXjw8v6QjIEArghYKi/8d4Hir/
aNE6xYWnv2xPn3uMkY+xpUHwHb/eu0XybgNx0hvCoIPlAUe+/xnQImv/2LIXG5hK
1Ipjt9YkOJYaoYjGbWPVrV4VzWPUHrU90M7rPQ2a3fI813wE4J04DtPzXzdREpzw
rEy64kOz7qGSt1aT30tRoqGP2fVj0tRJrRwtNA13haCLerzci2/PW/DJOjLCDFaN
s0jxHXhvPWWGV8fvG0dOXYabD2vZVknUJIYjVhT8iMdjENkJV4rkvrkgv0gJEfaK
flCBYaFEEk/24w/7chzFgt5/X5l7oNK5oupYaBdd2UTF4syg/DEcRpow3kDpiGV4
1XrhT5lRUFlB8uoU/fgPOZB3RVEOppOGu/oPJfw4xH2DWMmKwmjO/ycKH4I4T82W
6T/ojedt6yblWaJVP9STaWDLOJ8+a7RNEOJo7cDPecvhBd+EoeU99UrLhoLrxLML
8hADSktuqn7ffscTOdd9AGvw8+/V/LfTCE0gFaLBpVQ7Hd2SaofHBX23+1nWXV6S
B4ESWrl6u9yUBAlExP9IC7zbva9JnGI64F4TLb4JAyC9CnXsra7HM3fc6V/9YkZC
8EuK3EDC04xtjgZVi2rQR20T/V9jnVx4DXADB5OL7k+U2W8EboMnavx6frPTI4Me
zDKPSIMEzC5tJ8rHLYb/v1zdTNpl/WNRW+RCcXl/kYLY0nGurpqxZ5Kz14sJaC2Z
HELGb0XrY40Iqoer/mK1f4HMJvTBQcyaqUbYB4+xZzGhF/EVCaG38J31y21RXry0
BXL1xr+JXvJszZ06Y0A+lZXY28Hty0kJiWNEQzDpmNDSanJZ8SRPIpSiAhZE4HVg
NTQ2ea7FA368LjUoTRSuierT6nefCnDn80XHB3VOTPGMI8mnJQBgWvlLIjYet7QP
hJodjhJ5HYOhX/wXQDrNtmOXbtwAwBEP0pa9Wytg7/NmbftJ0wkNwLL70lxzyAwP
4UTEKpzWVzuTGqunrXjOtmg4TC11OhDeVcE6KiEeTi6463j62tYKZg2MbyS8x3v3
+LL2f9DzCNZnRSlsp0HqSp4NL3F/Grge5tWs3Xf4qRVvIh2j04Mk+QAWVzR2Taii
xUNNnckCIRjaIgFPFbLpEZvZzRfvz8MAU025DzLp5xYDOonCZJebXD2LEIrB+N1u
2BgS+o/sPyHFa5UYJbTCib3LZ/o7UUvjpDdyiFR6qrThmY/PsKSQvw/dB+RS2RY6
BN40YmNbPpoVbm5jdnizaY32xl2UDNpfSSuZWWLj+NFAfMOkWRltSLH1/WEf7rQM
J3WQtGLPczPD9rdLStsVAj2bXXvyMZpF6uFaQCeAK74iKVTlEnN/5jwne0Lbobip
lbdzInvmLJ7fCXvCDMb+afzjKLjkClQbB02ux+2z0JlxjV3PN/weNkfXfZFJp9lT
gkJAyZbeZbCtVmI20gK3IxseurREcd9apMc1lnMxGbyoD9Qxt6wpLKR6sqdNG7Pl
NAfPUgwGlqW7ayhYf79iCtuqAFjtO5BV8l3JN2JQIcm++HiD8vKnDqo/rhtUPoDf
LCXzdirbkj0+yt+QljU3lN8qo4syZ6GbfPJRw7ivJgBkeKow82DrT+RDVQYpiAY2
iXyvDeEAMDvG3jnkyUsFaF6VTFt9QGwYvpQW/g86QQAnGENNuMt1KQy/WR76DDrt
WH+D8WngvvpMD+f4GlqTOQOrIJsYetoCWes2H69aiFxb2uabSXzcvHuVLc61sWzE
p1BJcsx7rWInJIIItc1U1F1YAWeCsIgwWaatm/uuczAZRcWdt58iBrAIQM/a6YC3
sGprjCm/gg+KY39tRpqpK+xSZ8fhd8YVlVBvzEgngg+KlvrCu83wr3uhink0Ph+b
hgvOkPK3rzJSz/uL85kzYSJCnLkCct2F4bINePtyJAF9HA31RpsVTITgIYTKIbER
JmfCDow0TvUHGB4ElVv7iq0p0bQkXBKms1Ys1Lfnz4lCst40gYn+LmOwvn+RpQHo
dKSUwvb6piGRa9BeTkGP1SbT06AucOXmsgB8rUWYdEYYr2MMGkmf5Tr9ASKX8YjA
UYuMkAb/YNcspkZ8dtpWnX1ak5O7iRmLU/Xy9Gjlxu7Y2EtNlKk6SUE5HxpK5031
sOCU4p2bGt+gQ8haBCGKFSDcjQ8vZLEqOKooNrtPdj6Q5nthojwdHbJ+YLLhLDpg
6ET7X5WXUSIhBJPOAatb/JyzYlm79GMz2hNJCOROgYIUdsZ/TozZZ5giIgVK8RJp
NTutkxvW6QUIOViRo+JEQk6yLzZ+DzeR6d3zIr+OWUfOV7BOX3BxmqyUSIKYNp0n
WQmgicNRI9uKZFsbEtF4uBJubygnJpK4XSL5idKjm6tBPv+o3sUSvcrHU7E2ibU1
Wsicx/UsO/MPNzgw5RBbfbXjwTZe00dmabvG2WONdwux60NuctRAeBuU+tRMMztH
+6PI9UrC9uAvq3W4uTJdWlBbCZkBZ89xA3ebJaowNQ7NN/u6UC/LA8xFvOgLVzH1
w7DdrF77IHTo6hHJ4Qxomac3fjF59sqxTXvm6MR3a+c/tTsPh2cHsivW5WfgjCGE
uzPjOtF9toRKyC7jfoV+GUHb17LdehdieL2Y6p6E6wjMv8aM49OdCbwjlrhLPPQr
DJhd1tyL5HqR2soDfzAR019fExaHzRHQE290zKri78GNl7C0qYTeAMjbcWwhtWOa
r9SVrhjUTtzuhdBjH8ZDbGr2KNSkqTXlQKudRUzYlmcmvQQPjy6bxlzcJRfLSFH7
RiwG4NmlYlEWkYZTMTpG2MMo1zX3hkRY0Dsm0vZ4xjo6xDiJcIEdJ+lZwF83gaqi
GQtGZxs+lxVPzkrxo3fpkmfEAiuoEYVEmpHllyuOkqSEFGzPuORfxlPeM28SOkBf
dYOdGD3C+yzLPy6Zc94YV4XT1+xLPoRXE5ZzJdCD8XFnRsk4ju9WNvRQACmATLgS
suZqQsE4TgFFg5A6unmNJzPAQupVaAVCQALggDgKzOy3FpxrQXeE8XfKOGVOUYyb
RzF9wrCvMqhA4o7O+8dMpoAmA2iRbEf/9EoRbd0Ewthw1A/goQTWZBNK6l5VIes2
WaooTlD4yaXNvK70wSRedWlN43nf9Z/p6/ds8AuqyoeWLp4940Bslb/AzG0hSTde
Swa3MzPVuebEGhi94ONgc3CBiwLVESWd+EsRpxf7HwItND4hkW78wnlIN5MJ4Fn8
AvoUNYvduzrcV5Pb8zga9Q3lw8P7Q6HNQwODCje7CVmiiEn1cNuiFj3pjwwWdl15
acqcOg06mjhjZJK6WN/mS5kcNIMRHfgtK4w/RWSpIVXfuqGcVSU9725z/MnIgTdL
QNGczqj+KwIfbGtXZQq1ilyuLa70DcbS2mbrQp5EsmaVaEWhBR/CUgvsYvoF5l9o
cDQCdRzAxPIsLnAOq68YQtWplyDjplR5gvWRmPXHQzrtmRdZ8b54PJ8fOvZB/TgR
ZdMdkQ1Z74lRMhX6R7eBmNCXZh9x8i1MyFjD9pZhagVuU+f2mqvj+0eggapFbmb/
1yRIRZlaryMspY9WpOwGv8fiU8emwokXCS6EbCuoxJ3XxBodi1vJZ+8ITad5daJ2
c9FmiveeYyBQBUFIB+hIa1lH4A3voTD5ae9K/A6z3XxAV8/HaHdWIybhN8sAjmcX
Dje3uJUBrDx6vPKsy8/60b5ZTw/8RzsEj4fvhggRdV1Ep1QYJ0o5pFWGGUA2da6F
nJlGfwEIhSUh63LHrr9nNZwCqUsB2AKQSkv0pS5SbmCyssrs95aYbFTqqs+QP+O7
ZoIhSu3EMsTwMuXaJSr7B5IMbAHnhPz1voEwFybo40JZpFLeSKfYtCJu9y9Ird6s
sflXTUf2ecCGrmT8fp/YvIa/vEEoC4xFFwyilzvjSNzOKpHi2x/0jydwzTURzkop
9G9cry6AzVbeHwF+Lmm4ZlHnXncQlpqiYMUsqkneiqA/4rUbGTKOteBrKyDFy2rk
aSb3wj0obHMQoibmbQn3E7p21lmNDrKujH7nZBy1USpmANTV+CNPMpUVt1HHjDah
ugqHMRXdG7XGMhZ4YIRvMexutRPpV3eqRWGi8Z39Zb/zOvI02FkE4xEAEJn9728b
350u64bVZzVsPfGC5Lwq3/9f4JmkJAOVe2JH/LASNvJj5xjoVJdxF8sNZHmueYep
N/9y/biftg0YF4c1Qi23SE80UVrhKngnDJD87//K4Uo6RO05Oh6nkFi2q9ZZjgyN
q50uvn7qG8iFHNA5nt9BwT4IJAd70o04x7j1kkjMhs91cOWOBfnNCWogvj/mi0wt
r7z1YPuLgWgcLCxpU0uPxuDdJvyytMQ6rUNhJDh7QgoV/ie5u3pQa3H9klrxO3ja
IDeO5JNAw56CGNpN7ja+yrpXPWAc32fx+mAkXhrLnFZ0aXVs+NFNj+5lKBnRWdSW
DCTPGRkBXoD7mha2tw+6dBMQeZ9ToKRp5WcBgvoUeU2JqyQwhNh0SLySWLNc3BJY
B9nrfww2gMGQhSFtTR4XG4zDIVIHbYycqS1BiscD8z8+YEjUeWdiAsxkVnoqAt75
LyR674am0yHRQ5pITFySEUL3sjw936sxadnZvlHs1f/B65Et8SG/vyb1M9INahFq
o4VjCALap2PDwv3EhCgBzjz6dePg36orFTcA8DumqpcTy0xqgQoON91gwKOSh9gG
0Jp3Ch3e9wFJTKoKey7LEU5e9lqdQxWyQpYw/I/PT2tNH/l+lfYMkBoGQK42qgSr
FGrd/6+nRGm4XKyVEnIQrNS2t97r4f6Fo7JuHwazmHCszpSZnAaywexm2al7fi+I
J0HP9X92kKyZ4m12XGjwmPUTMMKEMlLrTB7Kv31yhVsojUqgBKXy2ZcVMhSWpq8O
erC722dH6SXWvBJ/aZ5alCTo9+yuXdLruX8DHbSlddkqY1jb/w6zbAbqMIl+twKA
OQHs1v3yws7RR4MN0b1olphylz+M0sBVN6FcamXtx+U5au3JZn/K9wYfNTY0bocN
UwcjkSCH0sLdfRuIHxy0LzSlPossWyCAuzNJBLLMZ5gUvb8+Ow/CMh/RzMupZlkh
q5nznVMPqDOoVDMd9lQ1iMYm/9LAlpLdmDZBDv2Nscz5/1QsO+idh67R+WERXcGP
8ox2X9GMOAgYI1hpPlAyTyhVbe7ZEVp9IiMAq+rPtLjmNAWDmVfcl4TIVw6Ytnh1
BauvZgae80fjbP7qDEpZxJE1OiwakbecKT4RhkIdHZZdYWWxzbcnoleG1tDT9IjB
A+aCt3s9ecQpJshEn/j1hgdRlh2jzMYMI/KRPhbg0l15RXML+/gM5qq0NSj+VwGY
d6WpvAcOSiGIft5sKMV9Bqa257tmDEXiF1wzTG4xUcg97MyMSLRxBAFkJu3SB+Aa
PGsHq2onBF7/un784nF2Ub11l5XnzZY3EdV3SzausmSBWVNSxJd1v7cIqxYU5Xk8
OdG4lvy3bLkRH4myPCGxjllQ7GmMNwZa8N+iEJUyIT3UZVvj5fxfAADHr/RlTLdK
udQ/uzpBeJdWoIzH2JEIoTviwI8OqKYCji/87oCAcB22vAFpm+cBz70uHN3ULG4o
WBe+bN8crslUGWnJDBfHpmqDJ71Yh0izOYAL1i6sfL4GXaGxRZOe5ZBMeJA5p8wd
NbmsyBBL68D860aELoTGI3JMcpe9b6MI2jyqsBQQ1xZZwy+bix8xukbvwXUTbLgr
CvygUOjFBBe2Phxa3qbPoMj+nsIZDVlUEKZo4H8tNoMSeLxggnl7T42o3GeomKPV
Q585NnC6yFGaOWPWKnMzV5wYj5+5f5LJKfZnLH5gY1VSdT1ZZ00tDCZUVnEPzf1B
18CTgLD8Fa6mRld+uNyRgEldgpsUTYaD0663dyUuFMy+MDzi+ouWf2fmaJ1MsUA3
nZYQmlOafZ1dO8jAlQqEHV3IFS3hLF2Dgu6qsuzL1IDzDEMRa7LhWTYOUmUaIauo
SCLFmSIP1Pl2O+iPj7hsOMHqUXFcN/GE9167wxRNL6IeLluFxYNvEh1fO494KeX7
8Ie9wMbApUAdg6A53TP1ySrNf4iwZowtgAzkhUu56/kV8vKremndM/j4YbRdcz52
ieLabTyC6SxEtE4IjF09DKGY0loQYdvJxh1Qdq1jI1/AZ60aG2Kd69VA8Bx6fmoW
rO4du571Va28K0SKWp+KMBNdpecNb4KcLJZqH4jGFuvdsn+g/LjU/3/bjnYBGuCj
RCjFiPPr98yStaH4JyeAh+3rYz0uQRrPH7aZd9ej7wL2cM87eDm2qiaora6Q2aVC
FZk97Q1HsY5b5O8+leMTe1TjuArxj52IiH2As7tGlq8BWMBAaqRClUC5Zf1xihMD
gXf61kfbqHyteA9ZyGHPraQDIN0qZbayxmmv4rOiaPmwAd6f85B7e87mI/CfAvUh
1EZq5XwMpFa/zhlWBK7pirPlq4ZnOYhyi5h9fb+4WKLPaGcF7HJrTqUgqI4/TBic
jNbfhWB9SzLazNByGeY1/F/gOeij7xVedtPHPLSD16lcKveYRYVCnVrjnTd/NxEL
jQRLUrPaDPFXqB640FNPdCtLptq70/ZCKpitBuo7U6om9a4zQIHDxY+bnFOSYkYq
DtQhkJQ36Wxx7AmBGy7DzXJNUsowJHjfvmfBujRBm3Po1kpeOmV+AZrHcHcEFHX9
tehqLFLO9T3h0aZFPTyF8RJuWPVFDPwHF7XPt73+q9Jw+Tu8hHh9l0JR8byr48pG
RiAHq+L9sAIRmMOSRsn/x7Jo1btmdpW/ESt9Odoor5a+DuZje7ogyfnuKvwM6Wha
X8BfMmTMZ1sDaCoN1xrR1ik+S4B7U48xQkuqFxs2Oa6GVNIx5tlBhkTC1Q7BCOtD
nqY3/afwwuuGdg2x3KIZZx678wjwgBIwny/iytGrnQFw7p7265zxQPO5z/9Sqpb4
UGPJsX4MsF4nx/Jf2mjW+/d4QwpkNRDAfj7/7Ks+ropgaswQxL1glZgYB+w2kXVe
uUSfgrtlgvPtyV9iKj04K64th/I+x3ixVX8sfml7P0LKpXqOGcdTSdkqr86wzF7V
3l2uZ6rFRFI2oG/dp4MU/5D2GsjEj8s2iRNdF0dnWdeEhhEiGGl4rnC9aCSiyb7Q
y6VmN8OyYmvmuOqIcB+UEUVktUB9FgsRWu4c4JvFpmjiwjAXORdwEDK04eEdnT0J
0NAmF5vN5APbKLCsW1pV0W6K7VurdrgP0eXCQugyCF2d3Or5Erh5kIz+OMh57KFj
l4OIAVzr3p+J3qFKYSePLgID1FVIkeH0EP7eKjTZUtlHNtYZsHps5t2cuQC4BEzB
5uFWqrOH06xS/iQO+KOOobfWwD9WXR6xIZMN6BXbczW325UVirdPUEYihUnUDD7u
sKQ/wDdDdhkx3pzwwZDduTkHrUtFHMmGMteKxt13rxFWZyY+eNKuVvRPr0wUedpN
hZgyfI7Rc3myF5/YkNsPAkCLWI2moCqBn8WfyRa8aiCm+gHdvYhBN2oZYrNeSzY2
WuLDMWDxzwnaMUKe/XkWF4KkGv527vGgJ9FHUK8L1/Zo9AzuwGU5NlaxQ9WE1iT9
uicF8Qso37JsRQ6b5m28WcFgyjbXI0JaAaDEUYSv6hdy/8SMRM5uAsmK8CtGlMxJ
587Ai+iea+VMKFGflynKv2pgcJIGziWiyXq+lr68USY8R1FeEUc/9xfoUl+q60gG
MtCpzbM44uOTJGqvH/XjW5QLDsu3jcWrN8T5NHY6/8DxlNNZ6LLXEvfH6bMSPvYh
HNjg3+e4Ykdt1tpIjvhgzYGugQ6zGMk8hI53MrDhACef33B/DNBhsTFwR2RuFtFA
f0FiejWGM3sFULhnnPNy11mTQLVp11tX2zAUa0Hmfm4F/uSxiA36BNn3PJwmpk4a
S/QSfxCv8Ftqa59zJFpW4I1RwWRJ2G6XVAWyfqO0Hh7oZuP6tLv0jAbmkVd1puH1
0lp8ToeLkrStsc2toFRJUZObrrn6qaGu4cCJAtwZ4bnKXR3ECgeZfrRr55t4y8SY
mwxM2i8rmeK5BrrjZNTfvHBD2O30lcg7zK0Hymj1/uHDQ+aItdmYTUikcbWOO+zO
ovQ/SHisdlIJUgvHHwvXlcbGnzlINZFNXnvqE1R/Q50YDkjwXmgCI+v9LJ1k5kwF
99l1t+mKvxfGIAaF9BXVst3NyYWegqv+vKrG17drsLl9yWmiYM2KE3xXAIJRb0Ln
/SDmFd4Hv+TKos8a8+Su3We7yyQdtjswTcna6ML4x4JUGnT4IDwD9+zp4V/ZNl0x
pWPXrDlMU+G8stRvEY+b8tluwwgxCzCLHyKgZua2JXI5BWzB2cXZRQv+gclHX3mb
4fYthCsR5T26Kq89cxRdH1LmOnsZYt6XJvfgW2hEs2J/G6OnIPzFoySSsu5sYWcq
0fc0oJtx28cupDdh1f5GBlKhMHw2iZfOXyDRmdN11SE3RsYfsCv1dZ2IWdFsEnoo
WD5QnRJiyH6QvqfIYaDIRNYfBHiODB6njeqMA1V8N3LDmsCd8fVggoiuN4xrk/Je
dKIcIEvkZ+6ejEhJbdlYcDeF7zKLwgluHEuw0e+AGoiKm60Tuo+feulnd/ZTPtKX
b5TrJZ7sckiUSkIra+M/Pf6/TvyuC4pXqo8c9drns/twmzOLo4rJw4INxcajwFej
aBugYzW6ReMs6i5Q59wSaqIa21k9fKs7ge33N59GqhCc1Iks/KkzIK1deXlsezbL
urumdWI+o+az1ygsLPSUUvRvt+nFV1E1fMMvU/hFdqpaRA/Z5t+OvNlJKZGGG+Id
eoRR57/27aM25DdjJOWnZYhMabWipW1zDizDCkAyLBaUIiqv2xZjq6H/7VYoGEes
OCJkz6m1Zc4H/ZDRFLAP0M2j+ieh1y01+AalirT207qqxqRRZM5UJoPRD4z8MagP
6iCoBy4uz6Y26Srg9p/UZzYUaE7C+jxYHfvpVnIumXQrr7JkScSayb8cVe65ErWU
BtLfg3fFCWTpfcdJpNQPqUIWpEikQIlft2Gv87aqThTIQz3nrmCVnlaWM93Ei4qi
w19iOMBjmdaUy1jZu+aiUgHePi0gTN+5QXhya9rU1QsWXkDXeNOQRU1T6HGoijzO
g0gl+crmjoFTsz4WW7mE5PPCYwacKitlbziJf9QQUbQNhwseIeB7pr4J9h9NXRXy
94G51nudlPAk5JNLCRe/U1E77eqrm4rag4sBL9z7ZJ0y7ovfsMveu55ZpqAlPur8
Auw+mFttxbgx8Yvl7WnOiejtzU16gLjWNAmz4Cn11UAL7+CrXxlWA5rKWzVom2lc
yQSOunpA1qHy7zUcLyJlq6NUB7g1gy2eRlfuljoLRejjxLi2mK1wZlOp/+i9d+ch
NY+tA9LKE+Mf9xhZpZxkkJqrMfN66u7iCuMaltAAeXOftfWYcRJF7nvvwNL+HVJq
+VYh9Fm+/d41+F4Psipr16NZJ76/FASEXlxKXETXoQ88TVOabsSC7xXPxJEOMV1d
4R6DIDVweXFGFOyXpCv+LkdWpNvM2O6ETodtmshGcG71KLodc9/+sh8PPqzOQB8F
SxT54idHScj/C4m4uSs77aGLg/11uRS3Qtt8PNEgzane/WvzQm6Fbxo2lYYsDc8U
npAQzMzxyhsaMHkerLekyw9bVWrMM3BG8PmsI7giyuoyZrscavYm+8vYua/M/dkx
vsAzoys3gB6wnuzsrUi78Z87v1tTnKG6A/TWifWJhnT4HB2YOYInyXoOVWa0GjEP
Y+odSJHrfG3L4fxCBVGpnR3AZi6sEKs+4o/+tsiVL15BXzFeqQnx9s3Mn7z6P4JG
SP9VhkN2TrBgytOfzBPZ/Q2pZHUXg+K8XCXzqsHtMPs6DQIiUKRCRA82B/n5mGMx
Kgp5YUoYlg0C8d8jXqvSQNgjfAPzQLbfyPVFoNXdezr9QspAyZ0FvR/JNL4JHWdt
jO96WWBBTiKZ5iHFUkV7lymTYxqKKY9S21+tEIIUFFq+jt11oLXUV5dgXD16nI4D
KErTVcTcYKqXDtNSfdJY/5uI0PUeiGqvdew4bTItFme501UHkUD8VHqOkbAHlB9A
i3+NjQM/nVtLKlPpCDm+kPnDgX2/Z1J1mbqVmscKlmLiyI24UkZDVyLyc2Q8wezK
W25WcixEedFWP33e5IBKsgOUIW5XhYpXnDsDDq7HKZ/I+zznlt9KPLxidSV1Oi1W
rVVbdXP9NJNLes92cyCFroGDSiFeZdQelR9ZVbLZ+C8DERVTMjNcpciXPy0j/rmy
D+1FvvJTAXsG0GDsYdFPcLsX8jH9WEpxIkL/b7MWlgKUJLKqIgJUMsjiPXfBmaa+
DvHrq2a0zleUTidweYB93xcQ55nfbJYb2GfB35o19rBXlPRBvs3M700/fQq/FxWW
5yBi9iJyTAxGkgeWihN3Z+V6zj/4ZvIAivWu1oHIdxPrOP8spA9EzNF6z24mEbNZ
4MhI/sCdYm8eozAhks4GFHHySBYHnHkv7+o4uklR2KAZ0TFHjGmfXjoXAADJlM7A
J72m3qJwohhEisXNoZdZ7VHz8onH4NTwanccDgaHmRYRhiLQRwRkd/AprT6qZ0tP
h4dXMzMYCwkT+gR/e5rp2LTxkuYIiZ01CcuoynZDCGo6IlCm1WeMQifKcOaO/le5
bV/b0ViwRXssxI+9+Gao7UleP0riypwozLDHHLigBowmOkkw1kF6EWmRPaO4auFO
dOt9WDVAKYY4WciG0qdDu2O5oKrQro9HoQYF2iZK3/lIU9huKpOz4IYDnRrgWm3b
q8GFz2NMyy4m3nLhYpYRjr1rnWAUOWBIMLzevMrWH5FlCNCwI29hYrG0AQePjVHN
HGsRXGWUkTQbmzZACNq2jDDfSDuIEAxFOZm8+JYdrFd04NjtSCrV6KrFplbsmxiZ
Ivoaz1yQpKyBSVe/iX3Y2qtc2BD+RnLlgnRUAtUI/hXRory2XDlz6Lw9k9AfnWfa
onWK90Ij/l/VXuvz/Lyr3khJQ1lyhFGz6LB1RpyAfDT87Cu5nISs5OULeOj2VQmg
4+g2ppFel1nPXG6e4kE/jFwk4+45tpesqqVbzpckDpz4H0on+JxUKB7x7CRlFgXV
igftZChMNddDCRuW6c2F3Y3jneDJxBaU+5w8czs+HxKlPTZYcmzoL4gfVPIuQsr6
JAAJwI3bjksMcJe+kX/mfb9euJsglzhZ9C0mGvBnwxH2CSa2MPvjLWAwK4OTALYk
bHslr0uEV8iT6IlC+RmkT+1uiXS7gAy+Hy4EGnqaoWSqIXEjg21i/JUQ31Bo29sb
w+2wg/SozSEwKqBx26Oip0co86yrJKFWM7JUZbr49yPAfNbWxB1rUx2xpHmWyBfb
ZE4T5/tRSEte3O4TApdyv3hHxd9schmop0IJj94KoJUEQ3piWAJ8QCct2oL2p/2o
VJjdsSbL0gdxXOlnVuCCw92RSS62F59JLYGqTUkqT3FwOztDiLmBFKulBKZgV+Qg
Wsm9OTm/u1lrLTjQDLELqzaGqNMjsK0olVtuVzbh0rT15mHVdsgyMem9dqD9/xOk
rRdMrT/ro1d47Y2xPpmbZKv3IByCKAKvns2ymPxv45EAyf4eICMtTNaIgcBEYqDq
F3CuSaK0xtLCmnL0HnV7O9kAornKviDIgX10O1f9cEobHYmz/3EdG/rNiyhdeb8m
zSya7slW+UmAEPLE+XiA3+qvGiJBMJpTntENLe+CYrPOG28c+S6jYhzYe11gvSI/
IeYv84pJHAmgoqW8zfw7HZXw7uMPMQjbcs54pNmK00AbTWSfjZIZllqLM/fH6RjS
2p1kyHyjCa2DltqjgZn+5t40kQTZ/YdRdc02YzEormVCKMVVrioakfPrxZ2vYwMt
kkULXQl4YQMhy4zr+2KZkv8zh+E1CvOzBaB2AkpWY/RRElhBgWACZuhz9J49x54a
tsAoD/2lpios1KkflGJlTFX0o5X1X8+zaogASVOYKoFnwA6t4yVul2TKCBrfumOF
pPQxI1urxD9theLIbH6qy6Vaw0gjScicdXYqIL+J/CVCZw4MiyRRjS7u0jJnQM2L
aZFa/4MSS8p5jlkDYnasQDHVAC/Gs4yfEh5gGjLcdDxR7A7PCFoM5USkJkCEcoRb
y6QNuwrS+J3/ikU8DFezi8A9NUfVpwcr0IdTZf84lRK4gFZ2nTo89SUY8hilMoyV
32JgpTKkr07OkzEDT0VX0Yk4ulDefu3TNajGeKPm2hUjbTjdQ+oLsynek2Eu5kDW
Z5QEMgZF6Sfubvoq1XIukHMphRDQArZBcQfQwanO3T1hhPOCVTc12HeCqolP6vWH
2lYhjN5QRdDTwGtvEHSFXQgvCk5HgDgiITxoCklGh0bQCh1frtBEM8H3OA9spMwa
ohYLY+EdszHRVP05p7XPNMk/qFU9P6V47X3+dIICtrxyECywQflBwASZ104ZLjHb
WXWNcjCsKfEep49NIGhLIQc1Ul97SOUtbisevBycnb73DnnUVymnvGyjIEgJ2hQ1
q0pul8DU3jp5yv/y1tZqB1w1cgz9DoX2yibKjBs/p0E0RBWCX8USeD/Xj0SHkLeb
//W0vy5tojX+FE6lGmmFLFFeI38XYBwK5eDqcsixaOAxFH/wfThMZGP6Rbz5AUk3
ZGSshcJCJ22s7gCfH5SHBiRORqefL6Y/vgDYiXEejZ15z+cn5lBeTYBl3zF31Es0
YWK7D4jeBeN/IZCwPjmarBmwzyQJiQaIKfoRmiQyxhdkEKAZzMl/wD3Ryi9E55NE
zIfB9vwvxJrjrI+gKmXv86eRaHnpU0NuRRVeu3vLEwUY+B75fa8WVLp4erjAkA05
MoIujPJ6ouejtf9Dk5wR5D5NCBgeLBjL/O8KAV0d9vBZSs2r72qJL/1+7oWu5MfI
+0XllreXXytS6+UoQxYucaZWenEO4dBYAkCZVzd1p+QkjjyTHEVXQJa5Cv8kP/3e
kEQ8vSEVs5I7PgvWbg6VPoYUaXOzeT9v0+OvUigiZVeX3N86IktfFR4z4ygVOlbu
BslBczlrMEBs11og6ZA84SH4NEYzw0ZYskUiPx8KtIS0ypfA3ZZTMVD6LBqjR0qO
3d98IYkjHn58pPtIglXg7IuIN/OIk9SInOU1PnXYFthkwknoAvC/nhULsXN9YNZt
Xy9174efBN62op/LPZjpEnMLANYd7Vac7BuCSmXzhyWf8CBYWvA3hR43KfyNtvWF
Vy1i4e6l1ZlygPtxLTLFvyLTHuMlHklD1lAu2fT4soeIs+2g+OhEruTkNWZYYqnD
a1LesCFTQACxProUXM3Yg1D+iuDWpc4YHx7hugnIDnAYwOOiBmYiT+Fr42toC7B3
7FZL51lSWPQDpdBklbkb7UGnQk3W9IHpw0z6p+9yu/hpd25m7nbiIX2ysDlDkELu
n7HQ2kJsQTcrWwZiyJRHsMG+6Swz7HhGrbZKXk9Ax+nTAGgOTBniyTNqsuvEq/MK
NZfN5SvJ3IprKhk+5hwGVkj6LJ9ZBCrklD+MbS8Aan8e8/Hv7g4R/dyK5Qudq8+B
oGoVWEZZuNAP5Qc6eSLUc/nOWxwVCqLtbyrd9ZHlTlBEEAiMxAY893gJCySTeA+i
kr4wU4K4r2NNXpZYk44FL1OoU3xAk3LIABaonBkafIkoblWlcXZwsYrF26IS1lyi
b3CwUN0qoaOtnOsZgXzeVtnZy+qdDnDv6kd87fWhhTSmSNUBxdipaF7wFA0LbidI
K9xzCt7qxQ0MllDUl2ijtn2h38jwxqkskz5mKDJtMXsP8BCAMMbjXTWh7VxsC0bG
URrjC7mNsIIKy3vfebPhKSwR7bY6b9d/JkJvDeOcE+FPvzoi9xac66YjlhqUdof1
WpBALYxcB9y1KX3S1GzIwyW+J5KB8O5nqFYRgvzQ81eT9ZHI4GYmCOmd9AObJzWr
9uVA57xp3O7/cy0+u3RG1nkbsNYUKtEg8CcbqQith5pTlDV+9FHyyDQMb/n7ufkp
hsfCFRp3B494KOEuHGhIDFnLoDKTGpYH2XSDxEG6ehXp/+Ron2bc5oDZ/GP6Bcrp
GQ5NR0Zkas9jKB3Oxoj4Ov1wlMcB6SVfFZ7dsD4UykB3ktZwe5VrMdNXseW5JwJu
hw5M8sYGry7kgZmfbrzA4uUSCnyYfqhCfgkBY9Iz5NhRqTe/wuvLD93FBc3Uvvf6
3lYTdJrsfAuBZgLRYeWkvEckdWcSh7J3D76Bh5Rw3wQDm8Y1cXcbN1/YwaNgdF2F
JuWpQ6P7eG3Z+dMBp+/QAdJLAr1oEttqwY62oKGCS/GxgOGAMvSEc2J7V2wgfSKX
F4GglW93HSFghzO5djxO+L3WgXQcTxz2NgpXmoD33FvzYnaJfgDUUZneLIx+bDQE
eu9ak/0tk0TFOby5Xu2I9+NfwojoTQbDoQoEidqkzkIhjlDqflZsqgw/2t7kkrRc
oQrsfzQxeCr+B0vrrJmYx0diajwXJo/Jrok7SDrTqKV6dNovMbrz0FVQqCa3mDP0
QzMDtjOvryqjK3SEsEer/J0XX3+IxcxnVnhzMx64wcP/IY06u8dnxo0+FG3QQu/z
5SmfdJDWOdc5gfFLjcZffp85+O7BjFJOrpxrPhdFFBmsV4inRxII5arUFzHhlia9
HcjvhOsYnDevWsQuHDiXwiOmVupsVWRR3W6Vtc0u03MNEgFDrWNGQqC6WJ2KsXEK
pRzFzzEhhxZLI/hAWZUcWx24OR3WY9qSumewZONMxJs5NCJnJPWVQMo5aR41xZhV
P4RSoDaaoJAoRX3PkERAzdSAEoFKbX1VgANutUbQJIuq6sIhLDSSGcm+NxNDqWVN
jU7wFN+cW+0/vi4jH5iPsxA/BNCPqJ01MVx1XXbccA8U7nvSAxyo3suHV7VHouPX
6UgcI9jS7GLCl4U9ljyuSGDVFglifusSqLCuFKD089f53SQG0I2yi3lWNyJsdI47
zqIdS49LYYEE5Q4v/8ifHOJKvYvZ3o9ZV7gqa34gRkSA0dwG0KE0C5ojGpKK/Zs2
AzykEbi6/VKfgVFtql33FvKybZmRFo6gMTM7EjYFbUVeZPmOROu63yT/KY3yiJLo
sjVL4agnK0rESROMPkkkI5DehxelhxRLaBogDPSIBK/MI8YwiR4V71++c0CAUoGz
vipsZA0NJDsk8rxice41U2tz7/totkpTzfeJm9PfhtcIWHUrl/aVAk4Jp7ccPM37
FGkdhicZkrB+8WgudJmZhXIz+AUKb8NWm3xV8Ylra3o9W2mdztc6h6+FTsmHhsQM
qxTQAicHBlhXjp59RqQ5h6v37Cr8ZWwgOBTw+A8iTdVRsljeQ9ZpYFfEwrqh2Da2
yzquoNPuLmhEEgL4IedRpC5SKFKLZ3COUkF+wzNcOcRPrU5iqN1IJZvzSEtduSM3
qjv50ry4Ho2UHSWvPkI1OUA0WzeBPY9ZyoIU/XJni3zoC9AYUEfc8xZzo4oyLRtw
ZKh014NpaRhZ8yaxAIadRi1PDmBnDlF0vwXoZBWq8zSRXi3htZnKmze9jGzF4u7J
yM/M0caqEH1T+aP6p7u4+Ui5LCiqR/uaTfqyE5sqHv7Q8XZdZeNDJeAFxxas52B9
gNK+zS/YOtXoAwrAVqEi1p4KQ8wmoHUkDCbdL+45cREx5nhzKcRt3ydnRpmpnZuT
vN6/8NpLIhqEJA/3b2dbC7eQqk2lhYA/n18idghS2QvvywzcoQOf2GHB3d6u0R0o
LOkdIbyXv8Ey7xngSUom0px3vpGayEqMah+NK8LQJsCsOz7n3lPORCi5YLAG07QV
RNcm/qbo4UHzsRPCT7dbxxLh4nl/tVf5DBwR18cPe+lO+qeVpc9pK9AOUV9z6JwP
iiNV+tfx055wMD4i83++XnA+qTa7jb3iCM/bhDsusrS5yiL8AvhV3q+OAhmSVX1k
DKG2AYRvmiZfYDKRiXyMP/OD8iRvu6DxIgwNHcXDrbbuXnJZvPYUn/pcRWE1YibG
o0heRWp7cdLXnLhu9MsHn3XHfdfdpzO5HkjKORHzX5TOi8azIY4XbI7bk2ce1Tl+
eX/oi4BPZ2rbN0StTDPd7jOYzDLm1mXEIquw3xdq6F08zqmMUaSeYscsZ0o72bNG
a301465Ix0HKqQbh6wCW+6X29weNHAgnN4s1wOxOYUiiO2wXf2AZPacFH0gp2Ho8
rm+UXiPWg0SkUlhELaV9LDz0YqDNJO46VmzJNJNDknseZ+IJvgPBxQEpS2B9qZtg
aKgYKJoZLtY3KfD8ecO5V+rl6Jf9iB36QU/WSqcPpbVnPOXgsIr1QU4HYAVUOknB
g4XVKXLcxhmnf8Y+cpBkAzBS7v2ukNsfxNn37iMcTzachzwC9UsPGDuW54ns5GGv
h45mTBsosN3CmYNnkiTC3NjeKW/9NIBAIGyKpy+8IOdBCmmBvTAzPXdMAL/CoUj9
HqWcnJo+i7rQ7DtsLKFsd2KqzFPhpiqW67zB6nuJg1SVSTCJ8enfyd3YQgN2jDF/
AIL5aSG1sL9/3R8UwZdNKP2eT4TdGfd5tASH2pQByRSVdWyEoQ0rc03rc8Sh1CYd
zg0MOItfYb0MnieDXqA2KUhvM6X2jc3/X9E3BMwlsNat/LDx+Sdm2WaZtMVcPVGn
VXdgNiUhy+mwhp2HgqWdzEwp4vn1Cxph9I6IgYBX4Jdt16u5caLQkUBCLGb/Bhmt
2m5sHiqgrTInk6cB3LkTFcVi5axC0s6CGqoSpKVv2kR0fAFwJsQnJVEuAOqIjXAH
eXOAdQ7Zte8dDwOxC3uV6a+/3SLPjviNwMcqfz7WBtoWQY1n5AgUaHenjXl+/ztZ
OUju8Olym8q5IqDBjca+O0h4Wiyd8QNCBtR3+2I0UMxvGVT5IPvc8JXhJjZBM2Zh
YPdZXxVGsgt2RP9Y+kUVkQ7UCi8oIXcjPEmWsYHk9MmzeFv0po3DRI1sEg2FEaae
zuasufHfs4OCzqQcGWsP2jA/5qRpzUGTq3F+6a+8pC0X657v3dfDnep8S6IuSKrW
dNAIJxBCq/lNQw5U7fWTuILkYDCvrAje9jQAZZ4n0chCDyR3LlYbJI6Uetib+AG5
0D5b1sd4u1DMOX5s35HJ5XAal1qQPsk3h50zS2Rn/cOkSHM0SQFJt/natP4mlNes
EojEqsZ1mLrbEIpHyodPZlySSNPgGJH/SNcmBlAwA8g+NIAWWUdsJnaxNYntjfLa
OMBGox3QZNdrknz9JET905+TZ3D9lOdB3obk8S9ls8I1KCN7YkHiU9eg8J5BRjZZ
yWQTgYQdMyCafHYLyJq7bOP8Ut17qSSDo7r/dAs4mbOj5nFVmFLZNVIqYVRmnfll
HIBRwAYLiFd1jVhDdyq+m3ifQ/ICLGqfoZzpqN2ElTPZSZdMOecQlZ4wPdMKqffy
dXPB/Jf4Arz3x/MUKf9vzNjTnCapM0tXvZ1GDQOLhF/yq6BIh8AtLLL8Rt+LhArc
8vsvQ3fahVw49/9MwGRwAyYuPlU9mZLVd1lSHc7Gu4tKuUh8GB4qQcI2QMbCyDA/
zI5HLiyVcmble12qwNSCxfB1yeq+yoUOq/qJmrmQaWV/mWipThjL8wq7PprIF+Gc
+Of25BzWEoGMyj9fUWD6ksNfsEeSDAne6ixVYY0JWWT8Merjil4gx6a9/KrB3w44
iQ2PHGmx9h74R3+M/bG8Z1k/QfCRhTaSCcPBFwQdXjNHk9UulCbiVTrvquzkjYMm
2gK1gR73v7yt8bDeQC3Pkwf6faWZi1/2beErXriPKpkM6szcbqyuZywrT4PJzLnw
41Wy3oE1LZ6z5K013lA+fveeNNCuj0t24ypCFpgv1vN+8DN9GxF6fmORxCu6e/U8
4P1ChMkwOIl8dCIehOmde6nVeEk8wYeapY6HxI3hWebIKB11Q7Yu4e0qMMq7pWaj
YAHNoJQbpjUzfUGLolZjnfN7mSOI5/WrsT2pYBlNwcHhXzy4HVndNeK3AoYIJWmt
awcini9zBlV1fLaJ28KCkSJ2yB0jHQYj6DrU4zlNcoZ1lskoOYaZ4CqcgTsYYpAW
nr6Yh2M0p3yBqndEG/27m1sCLMAu+FOIuwZqyWaNNJDzfgDJnNgG+8hzNzxzogf6
sCL2klXKOSoy1mD26KpQuSiWz15cTyyN9CFG4m3/B8v9piHTDY84vmQZg4HIzWrf
ebvM9eldIEEwuOzwCas6Cb+REpakpxF3hCCoWOJsahpqa5hpVhN9MiO08ZYsNbvq
/tlyOddUsjDHfyeR99aja6+kY+/DqwvWuBtL7D4dQp7hY0sSXF0JGbX7e5eU6xcV
uxS9NbPIWxoJMQcoU5nMNdP7tat4wAKk+J9dpDU9z9Lay5KSiKZ23n6P3AkVKpu7
O9dxqBvqjywMjBSRIYE54c3ShZCE5QaulEHz2V+K4gwy+6wMHD2WZBFS8ErjxRvL
UYgHBqpWLzUN5k2HdfPC3aqcoz/AaHTgf6R/lzqdIrUKEJfCFG9YfNvqeIZYGq5Y
O3jkQpfVcDFHW1Co0q4UJ6SrALo0o7BOTIYNuPpRsT9h755Su7KkDqtNda5iBW3R
7SevIohTnDxAz+dB+xy7n5Ynv/Z8ix8YhGIhq1NDtgbHqKOtrsXeEFdFMY1BPUQ1
bUYLYNY1373YK9cz18BeoAkFp9AbFVrLBBFPlrDLNZAXwFeM9na/mZ5M4dhWgzu1
01uP6RDeiTb2TuStVulmLhrV9LGVckBB4rPMrR9f6t2bnEkWxncFTmThR2nZiy7N
bR0E2+3mrCVZmevQn1qKxiIJQPHXnxZeJ1/okeLoJoZ+zAN2iv4HcJCcAB08+Np0
Cs0IdifB84t4j7c33NnGIPK4jxR/Pyc7SH3KRnxnOk0OHgVU7rTw5uiz4csaAtmd
lm5/UGhM3Dh0C/e1Lhu1QCcC0WX9o8dY1kTwuQLDABcwJ36U0RmUpEyHafO8BirI
EXFEdUhfoqzrLSivV2QVjI3UeYb+qz8dEvHD1JPkMs1av3tDSLJ9lLVp9mxxyp4v
2rX3nEBgqnnq+KiPeJKCY5ABoC9KfSe4HpiUK2/nN9mySwZ0VZCHiwMnsDDK6Z8W
QAuzLHv553bzNmUBYjHk+3SVZlrCJ6yv5ScfX8tlXLINsvFOnjzohw5wt4C8olK4
7EvQ6FI59Jy7Epa1t0GDtNp+qKqOmnLSMoWnGxQSgbumhcARF+uIzMiAPshmdPJA
hFQpKB3GqMjY3ugFOIRgvTnWatam8ZZv8DjUIEZBBwmiBgGKmWO1yS9UJMxWWpeu
UWqPP4AbBmbR9rnR7VvU/awd4EHp7aZOfvjnQ0rgo6Tm5BSzFOVDsorOzKzHZFnQ
1zZ4f4wyLV9kbRGlHav2wL2xDjBseGUJkaet2IUM3Wah8twmxOkxmUFiczrvvJF6
03uFWhtL0uX/zZCeAIIVQl2+89Gb7dGplNwTBIf5OarrYXhiJ6WopR8+vcDD31tb
VjFvwaDCTvaivb7agPgB9wzu+sVzgn/AmuSp+r1cmwBIaRLgvuJOzaEC3GMuYe6w
vKGys/GYo8AIFQgJzZbOnHt5zOuvtp7rT1UFGEZwScAVT2RKdBZ0d5REhk3K55DG
Ly2D6+MOsdF8vOrc8G3ZYpi/IPcRMjobvW0ypL7Nru8ZZJO8sf6y3nMGXJQNzBAM
JE+sqYfbfuqsNq/Z5SKCsT7E7+4imnjs3mpsBNvC/vaPK7Hf6hlqZwO8Mr6nz1S8
04StkM4jCqRCJQTVS4hb+l3mE8dQAAgYj+xLi7Qn8p6RnebCU8cDzB5AR8HbTf71
liRt0mtEsQY00WoOP1idpOvGjZoQlq7CbvwSTdqpPHVba7scEaCY6BOaAiylESyS
q9qEgtvb6RVc2KosJCoqgHwTIVCCZcd3tzILzOEu6dUgrxgO3Bb7+QL8G0a3DeK3
UQBzUl1Y3+5FItelOcy08HgFwbGA6vWpdk1tzRIq6k9DgGYPFF5chMZx5Z/DFxEQ
mAAcTOx9S+eNGut5kfD22XNSAJJEgYx3O7WiaCVPQL1R509seAeyvG5xCshipziN
fNb3eRNSWrykrVryBgkqMCnsVVSWJjp0c3bi2m68uSxva8vAgdEyZcATwfiW1z5k
/pRNxpekncucVfEgTAquIswR210B1GISnVciFdUozFKAEfu0pOWjsg27GjQDWVzf
lc7NLFVQ+BxngZAzW63AgFPFF9zQUeNfAVRJkOUW7wUY+i5cq6atUGGQ2s7Ki8gV
SgcvUB3xzD8m2bZH6M3+NDB1RkK/AG8fP1k/JgR/GoxVnYYz9MGjc5Q+ckxVXzSH
ogBpaH7+jE+vE/xwiyADKVdqc5WoGPTd7WK6N9Dhp3hVWu8g3g7ofP+xcKWcHb2M
NsL9lcnm11xSxi/Y1W5oX3rbQ+X/42kh7A7V7k7NXe/Qfk9K7hXjr8SKiThaoY/C
sI6zscVHkTBeYgnqEA5EayeU6AQ1VZEqkI+H2d84s964aOjA5F8qbLCNlDlbHuYO
1kkyndS24jWq/AHbEEXWNyUSVHE3+M6DLt6vA0qicsLPs4OvUACA7QKdZxE59CQG
/Oo1ryTsegBKI4D4Azc0fk42py5SoV6X4hpBeNxTDKKd76DgqQ6U5ERCyOXFnD4e
6AV6j6GQQQ7yLFhut10lApsNODnVwCQ+LdIIlseI9wSnez4iZO7eppshJllw7oLT
pe0PU8X1M8vwCrj+dntvTXI5l9xEBkOsyy5oNL/aqX+tEofMOQsbOmYlvyIDXEH5
m3dKTPLJBVeWUEf1C3aGiPfOzMjb76Y96xbBY0A59X70DFsNoWwfv5t9nXLSQgP+
4sErQ2FIbxWvjSdssU3TUpw/AP+ZfjhZ232vFtduH85vH4Zz36kM0WIop4zbu2Ad
w9Pj/xx7Fnae1cQht2eqSAfZhiI7ZTesYLXj9OzTg3FkBB9FSc+B9CWIQwF9czNH
/uJ4OXszGweacqJonZAbb+Hx+KRQhy5t0mFYMHEFbGaWwS/jIzxKu9KWY8pzQRrZ
TYKdpeOoyFz7fyZ4Ai42x2AJjIvWfNGfHqBt/GwEi4gTP7zrueXfwHcmD4zz3q/E
cOsvxOBNRkl7100BZDYFCC+dflDltUWu3HfyPMNCpOp7jn72UH5i5nt2hwy5kqWJ
24hnAGILypXsUJCJy5zvqcFCidBYIpexmKa7VIhzekj0XxVEJkGfEczD2BZ3wX0r
qzxfqdxsmtPuDIJ3MIaqcpSEe6xTbL+KeJucJL2sFFW798yJ5BSXNU3C7OMfrtxj
CScF0gS8HT0uPCr3vY58kfrD2GLkJAhwjfWp3z+eBvvJD5UqiOHTS9NH/b+F1+rW
X5BOmaFfu+b7WsxkSRULdgniSFPveu2dbSfZ2zHhxcFOqALoGIRz/EFuc90kdRZe
l+hx5NTAbV8bKv6Vl8FgG1DSrc1K8+FiUwc0BKfW7THGKc9AIcHgOxpVt5AycrBO
qQEt9dLbM8EFgTz7hWOUXG56bffdlCvVj1lHzJkz8ubHX676pe3UictOXOFKxruQ
7Wbh1vvyB8aBeqvY5tbxFSsvKrsJTX2CI2Crj7x4wYFbpnXFwkB8Kg2E9WxEw6Et
lJly25B+wum7a8TYxZ6sz0zqgp+Zr084ucalSTMTPW2vxlWYJb17c4xbn2P+IuLH
GfOKl99JdqW8BvlOhBZjG8GtleY6WAR9N94pe0szi3dzs2qwmbt9oIro0D0RsLZn
hBiTKWBLwSV5zD343qc2c0R3yQaXKcQv99gv8u7WsxUGXoKCTi3Y4V0oWhFMPKQJ
qUDW+OoPyDlBbZVuCP60hL/S8b0V38CoCCO+zsrWFEmFRZX0i1T0aPohxZ1Jg7Us
0m78r+oc5t7PPxCgXeIxsc07Z2jK9PIdPAtrm1R4zpKMzshm1oRaKcEjn+mOdyfj
VE5M8C9SVqy1YvxJ5x+ZSIhUiG9ISkBbJaqq7nRtqul/mju+NbjBkVbm0vhm3CvK
kD0kUoWqXESKHhbvhKfxu7Gnjo8MWXHcDjqceRC5eAS8jOWbREAcLX/lqm1nR2gv
aKDeEUIPWucn78rXl6yDWO+dEIXfICYPfzHC3qpyoM/HFoVXWgYUrhvJ+F1EmEvg
eIXvFjCeYpr0VfiCPZgRJGf+/5oruIBweCq/T+MEG9YIButYWffAhJ4VEky1Ceqx
F3gKfHDPMmvQ4C9GtGio4KyV5YOBKe9MFAX2EhHZPUkQd9Gg7RrRswHztiA/TNHn
wWpuGe9SbMQeALIM4CTN4HYLNk/m1TOE2lnme4Ol1d449JbzO04ONArOT/MH7QVT
JweAxXRAJhi8TowNbc7skgnJekaOvKNnBtPutpiTWdAzzj7a6V2/BbYrzq+1z/1P
YGj5uFNCwpKjW08fhXkNckKQa8CU9WrNZ4Koy5tdp10ib5FPJj88VSntbQ2N5VCM
78fZAo2RjTnMe9EX61L4FVA6mWDKFa++ye80YdZZhsQBweLAzP3xwbpPmCF4zbi7
FJEzYD7Hg57kWR5/gekdJGDVrAqe2Xgwk31xAQAemq5cbHUr2zh+lxt+dLEHQ0S/
BXEFSW5hfeQgdCHBwtA88emQcsqrWivt2T1nsPBdUWO4Fghre40G/LlmZum/j5XR
ofRxB8jLAHRXX48I2vFTmYPp/4wfwRlRkmfORrCp6LfHR1KRdXWxGQEpLV/TaFrm
eOuavjFGbggTYohfMIG6Q9CLVVBx6nDNd+3zspTpcKof1ppjkmR7OrX7zQJZY1Sp
s+SRhxP19iywefXpMxSYAKtXt1N2SIa9KawoF7A+RzvBRx10qOXaQr4VrkzUwx0l
1zMZcBKWL0I7UDJBjMy/UbCq9JEy7RHEoumFrLCYUl5bjvyDtDUQK4+XFVQ54qVr
9AJDxV+zadlzoa6D2V/1P46mQx30KDyVbQ675WAnOY2OEOjfMyoiz4DpSc6oE7at
uVik0K3xPCv/b/rMzeGPlWWIIXrEOt+MnYp6RyXVObhGhqoQNe+DtZ+PMykAjb7U
lIUDSDyGpN64TqsnHfe2Jm4+lS6dGLfRbl7DQDNqBbqabJRqfzJxf5GqJ/nMjjwa
UDqekfmjvy/kjL6OrJPvvZPY1nKYyItpvBx3F9olJR7HwKUdVVJ4mi32c7Fr4CQf
UMmKLpXbWczigrs/KmRu4Uo+9dNBpTgEA1KCbF6bdOxh1N8eS2RHVwzfF8isMRFP
qL9ZY/c/gAR1gQekRTIgjlzuvsuOL2TksF7hKiafG5l5m5SirUMBtuU7+9+RwVxY
H4bTBPkbxSqFkGLeQaYjHKpj63AuseYI52jwFJmmRMi6ZwOpUTLxVxIWQHhZo5Ua
T1d5NBUdwJ5ymUq2/ll+fS8PLtvuXroMTVz72/b2OYtH8B8YbTSTAEJmihDj9Kwy
3PNQPyD90EKzJ8s+JuWeBUtx1xw4NzAdnZFDxbxCWquLHJrv58wLJNzztsDUl5+d
CHZW/KEU0HQH3r6r3d6vhs2effL5aP+TAEUQGf2KHks/eethHRtl9fAdsKheP9e4
engGvgOllGyFc76UL0vZsoJexOwR2gT02bd4jOlKEZ50LyJ94HgJ3yjCc44RXhOf
hAvvx70QgnTpiVs4AW3hqyA618ieQXqUnTf/UNUpQmBpAQfx426JYAAgr9Tnav4a
/7eYOTXen2cxgtGUMcBdCQxhLq+zJFLduChh8cBBKVFwqEe9cbh0HYAaTgDn2mA6
t//0oHcrUPCxZCcMnf1kKJ6VjwUESYruRPiybDSWg5dIEPqM+OMoWoxLxNbiobdV
DsM4a5mAQuqJJZSxFsCxVAI3DMOnNXzEP3DXwX5WChLV4mqWYamqS6cvyHUaIZb9
8SJsIEMwfqBIVlne7gXhJt9SjALb4dItjte4jEWeIbKeyIAoNkzE6O8MCTzAqpNr
xVAX80Yaq9ZTX9QDuO2zhuWkUyvKjh6wZrs5W8o5fGGuwneKTdrpUhTYpwX1LbUb
cbWd04sqbj3zYI/klAZNYRfkGlwgb7RHl+YGTrCuyx3fWnKgHMvplPKAQ4mY0bqA
Q5nl7e/Jt116dcQxUDsVTcIx/YYfRe1a49/7FIJQmaJgRaxNlXDdRDLyJyDcUpPR
G9rxqD5Ul5R5JuKXGGf8joA1E9c54ZYJZzspQg4z0a7jHLKpXQsZ/xDNnh22nCrz
DaccJfbpl4LBnCYzX66TpoGh6S0+ZIkoWcDLBAE+aVHi7PKB1PI66zLACh/oQV3k
NW3vV9hUcCko/0Zyysvd9KswJ7vVOnN8/XP3V97ZRcmMLUeXwYTcC0X0fxDlQQhQ
LF6xhvpkcMIXaLyH4P0K/WRHykhG0AIz9j5PZ6e5G7vOVIC9A59DKAVP7JMSj1yR
b7zSxvNEeV1iu0rGyeAO6CirAXddUlHe0XwG6u1YgaZkT2Cy6dhdLeRiw19LXVPy
Ed70EL7v2yhZAwKkHtBjb6HYEH7REBMDDMFj0hMHFg2CXqlFxB3FO+DTZi0gu0vO
sKC7K9OvLgXwgAo8Yn9boBxm4D8xQ2MfKKlaga5CCp9tbwkGFxzfEdVmGtbdA98i
yQLDVK52IDHpMgaGYskoqx+pG9DcdQ4gmgJmwiceeWinxQDyE+jmxnBo51AlSMIw
q10aGxNups/D763bav2Eon+bF0KCGomWwWN6mCz83tagoFyC7/ihl3xhrXoF8Oid
Pu1Tt4rLZvCWfdZUltIqF2ntzK/klhCf+NCexoHrx3HzriclvMawiUszWpMK8pqI
7tlFLL8pUSR5P3wZjdyMmmKEf2ykeSGaH4Cmz36r7txA9+F+1T3YbwmilrdyQ/K7
rxGhypgJvR9s+ksScJeFAl1j7Yqeeqbu/sIvk7iIpZV0RMS+S8raEObA1uqo+slm
J/4qQcys9QwCdYZ+bPc19wMIKkCXSuaPwoITNCqlzh1cNzFUFxqW7iz13Yj915R3
OFf0Cp3DnNJLPMwmD4wv4ZIIN9E9D9R1fzDcu0/EyLpxXePn+2SmdO9bHPEaCW3g
zbVnXlfn1lrxJtNfM0GzjEJLfoWikqTQq3pImQWSv8mH1HB85EOJXzMAQt7ZpWI+
Thk1aR+LQBWNumr4B+P1YImjILLUL8mphVZe8JqICvusp4+JiF0mktglh8Uzmxq9
juL8AavM5P5FxGNm7dU+Yt1vhg7/hvBQmjoRhnLzPv5UzUiJe4iqoQYgCVrhzUv8
S2C1LFjwYznFdqHmlRy1+G+8pKXctKxc310RtzuKONSpr0Q+eqo2+2lq969GVpoU
zrUV2KScVujgf7hDl3+IPSdSyVswzcgvDfaw8P4859k10Aelvn4eol6E/c2IAT1l
lQUtVOu31yzXYxpK1p50S6zif9fuRGo4Iqbi1q3w6HJozMnZQx6fBTEs2PJ+Dzqc
38anUtHJDxYgublSDJcYpPX0PwfbJMkkCaqjkVdE2D/b9xYqxxW2UORFuUR55BHX
SRIm5NnxUuW5nr2GtuSB+Y+QTb6WE3JNWM4j+rMeYAgHKTBf5mLVkyfOqnmucDT1
ppmPcZ1/szOyU4LZ8IOQtnKZR0u9wAVzM/miFmFEy5W0V7BdMQKNfCos1qD9YMuB
SW8HHxTigkHzwLAYSnOONP1sDsveRezQq3dgy/lwIrsRDU4PzOl+tI/BtlDjE86N
YHB3kg6EfQnZ+X+XXPX1xKkY4H+HQyJ8T1qXz9WF5B7CrXBqjGWGPX3clFr+l4YC
PoUzym3GKe5vg5PVi5lkAf2nkFOMhIOA4j0NETaTSNJ6MzIVF28HcneObf0iyb/s
6YNXzd/InIjN/oZD1Rb2TDewc4VfzLnExrt8dYVmz2Pudaf8Ng702fMrTAKjIK8e
BrfXIZyTmQwIl2NYCehckoIo13GunddF8QCmxlWOBJvByM855BWdjMwHAXneahj7
CyPALS9ol+/0x8XXbo/RREx4tQSRkUmsWLLHrxIPe+mJAfwXJBIbqNskh/3sG7ar
JSmlazGCiiFvnoZ6G4zjyRRUgugcCmroB8o/frjxe6TMB3DEELt62hdJUEi+7Lho
sl8ZeJH2QJZutVAgTnOJ+XIZ5NRDg7VmfO8VrMLnFSyVIWu4/S5pvmVc9v8Q9Tpf
gXqN8pSowcD+CR4f1kOPnZ4FxuHUO5dRPkU7zmb7mdjTgrM92eodV3MYKAXXNQl8
44eR0g8s6xLxiA8jvu2V+Y+Pi0o7ssOKnhFyKEG6EsnpON50N+msfeUaGcCm+WQa
Yl7RMDy+qL4QEhK1hmqU2f1FawarphuMyJDO4XsMw+1RNL3ii941ylljWddMfUgJ
OEjFSJmvYzyxY27i5eLOhVef3e4112Vxq/4nCxh9dg2JoFxe2LKXSFfus+LNbMG7
p0nncI6x7bP47zyb2D9tgSg8zQBRH2CqYGts1W0qNojR02bEBBernCSvN21+GcPp
sSaEy2HFGPiEpAThhCRBJU4zmSZQLxIovQCWkrKTylu1g4j2khhO/G5z5xQntM5q
XvrdiVJqx9JvnBm/PumgXEgmEVuuFHtoNPjiuQ3xyTdNp6OsDg0g4OrCv4GOXNHg
fkZnjP5Sw+iSz8OmBMEN1t5B1AL+tZiuSvNNMbtsfw3I/XME+fsJQAV2+2x6H/5W
LcTqGQv/2gwF5RRdjzGivlVg3R0mVSyvYTAn6H7UW6c6UnstXt37oFl/RpdueN35
MihXeGa5eI6ubF+VVLMEph+Bf0jwexZyKWO0vOoTFT8KUu3hgD4tZ35PBAcmT5LN
4lj2tiNfA4tnt9AVw6qQFKdATSF8IqYaD3qcdy6iuwZH7Iamx7oIKifmF//g1geq
rivXB4s1sx3R5aGlReuukmVj0+ABHzoJjmiB/z2uuHFRz9uBEbKQShm9Q3ahwHfY
YJVK6XnAHhe3wiK0S00aQ1OiNpLQsjuo+X8lZdK1LTZ3UxZchDCpr5TtlBRSO6he
DjYMetC0XHJeezQ2CB08VroXR239xCUmPkR69JJr0YRXRfGsgP9PneSjWZKO2xfW
dBFr6hDMJcvDcnj2PM6ndPQsWMNEwjaHcVZdYE7pNjEdSy74V4aqMmW9W9sh5py2
SiWS3YUnUWq2PyWxKrIFXUBIVq/QhDVwmtYfaQ9+tTTPd4DVPne8nnBM0OCPd+n4
lgOBLs90/Nf5j+P5xLg7k7MbQjadSR3LmJkHZPFXEw0wXVnmkHMw4Tt6IR48l3LK
gld+Per8IEDAHhfGC7v5PQj7ObKRI7Ndbp+DDyAPYbXvMWUbIuuPW/gL7S1/tduT
0DOyYvB4VVOwzNkKuG3mWslwDbn2ID3c7FfgjYu5BOIs1Gg5/gxE/QLTVyy/R7pB
VoYTaGX8RmLrzYen4BsTNYq/uiP+u2YjPOmxxbHc5ZbVLPcChkLzoX5/Te8TZATA
BOsb9jxcKN6JMA89G6JXHDrpr1jghOotzHb1ygyqD65ZE3dOiSkNwe+OCis6EtCj
ur7I01f+9V34fE+tC/ckOTGy6GKeh9T5BxwD3XCIWKFFn7Ms9KaREYK2zeHmHxBb
dhsVADgqtJFx7CqQDyZbXBrWIWtAUrqjlq35rKXhNf9nP3oQ9x6yJLWAuctgIKqB
hQPD/NoZOhD2KntWXDwGIxSzQXtJUPh6FUNZ/RKrO+OisuCLpbttrA1OY+f2PYMK
R33zfU9NPyNtQkTCgkQM8ik/uBaztigR+bQkbwxprFlM3KYx3e7StC3hj2PztvFE
NqeZ2EaHhTyvhvscHtSXSamceZSg50jUVunNnJNYU0e+Swf11GKtL+WlneyZq7d3
UqUTmAMP7w9kAOa2znpITwqXi3203ThUkVHCGGt+bmA9FGT0sfaLpg58Q45DllbM
zSvbREkUnxrDKxPC9A+jsyTZUeFQNisi2Nj/ABarHLj6xl+tDqHcBHdFMSCnw8yz
FLh8hhVJfFmpSUjImTgXEwAJPmGl6fwEWGuz6AzN9QORChPTekNeb8dKDBq2asTm
1zjZHI8+hHkeZCVS3i9oWU5hVjUZoiazbWK9Y7jKG5S6WiEnEEAw9JAv22b2b60U
lbXs+O4lEXuEjq8CGZlymCo1jE28/4uT9QKUeerqfa7QQJrFzo1FP8Ar/H+JpHEO
XpLFrjX17GhH8kIV7PBDJZtmsaqvfRBMLMUW2jDyi5y1k8zGceL76AdMJ9EmyRX+
raXdckhpTGKIluBu6GL7gcztehpK4jVvAAH7B8kJnzqaRzpQLrwqq4dRR4/mDKTX
oOvHZM/9zns9ZRzO4rNO27vRfs7KtEQ0LEL01YBl78MdLEks0VHjAn+dESnUtje7
S8ZB2lA/eOz5kbFDdJaDdOaVZFVWxH4vguBsyY19sZpte0PGh2W50EQlvWu3f3Zg
HM/isezK6UUqQEWlvTKYzS4HRTZX+jO8FLUfcUs91hkIuvsGUPBFqIFZN3VpDJEt
wsrojx35zAkvvBnTFvVnNOsrMuypuuYTBF8rAx6zV7qpxIM1b/HWRLOVxrE2V8AO
pVXh8h8qYVZb3ebu4J7g33BRhwBG15D9V7DCxkCP6cGYpS1Q3k85rM11tyVHPr7m
OopzgD4dCMacJDle3JjmcMVcx/pv/RtC+XGFWdkdzSoMIIcvTl9RwrQGSP+m/TuI
utGxiuiTeIK1pJkO8/ZxxTTKCwJoHA1N6CH2AbHLwO5nIPVA/6uIH9pKreyO3iJa
AaXRCA3B9y3FfhoSjmb8lxp7QorFAgPjOTXhD99tvGGVwkJfFeNTLZRZx2gExO0W
Eg2B3Q7yeSG9wLQGo+kH5DKYljrfrniSh9TD2pXdkz3teV/84Si7mO4NWL8sAo7W
CbbEfrXHfqD0ZaFj5vn4aqRyetvoP6/DhsW3QRNXrbDqi4FtPQipSvCvKZGcaE3L
U6RbPJ6K6nR5qG2AxRr8xfVUU/0y7ej32rxLddU+oHHrrkZyVwX6VcQ7fZ0xHlhv
K/sl2DSPmbvxZuDerBvaxT6h/p6k83bUQitOeRGaPACp6ZcBCRVT2icLev4tZkJY
NYhK03UnxWjawV+3Gv0FmssmAQcRGh5aF/LY/cMlP+xxm3UFThlzmaUbNJ/KzAWt
0gPTqY8ksX07nl588c275vxqYvl1byGwvL8Q0QVCjjA55OADUyjwfz9Lvg3qk1Mf
dMUx6F9zvaYL/OKZusSrvjT2M1teKGk/b5LYJG/FgztMGkZjeYVXDh4jhqf1sjDS
F4C6iu5mcF427L99nNrM0U7jp73vq+02A0lxBmSM5swsqdrvyrFqeHgKPRddFSOG
C3lgc90BGZvt1GKWO3MGauql8Nfj6FKnTZsjkaZCQ+jzn6FepJ7uMPtTa8Fe7zLa
AAgPmtyXKP15PfU12sZ8KU4IG+v1LiLKHmmZdj8UZl/ShCt/HXAArrLdUON8I03B
PYDRwRP4z2h7yHL9GEG7WPv1cwN7gYe7B/Z89Zai3XCVRtikgiR8UoJp3zojiVoq
8+1bo/c7oo0lAi1QB2QOM3bev03u5adwq/wjl+SJNZRYR1Y6LJxyl0bSrieJ027q
UDaFqxZKsIFfnQ564983fFQLI5oBzNevieIYtW0EB+9Jn7azcj3Kf23pdXmAC7JG
3Y+m41ppG5KaO0e15K7z0Jh30BzJtyArkYqbrbz56R+4DTKxNkJqV351gwy0h7Bf
yqF5LWrqisFjL4inUUe8WzoXc8Qd86p2nuQxitYlIppBfkHFPpjlyq9jTcUIUbYZ
tD8OVo5pQo1JC1276Wom6EjW34CnfgiWD/7GuE4KX8gCiaYP4/4jGnam1YF4Ckul
HMa+ZLEMFIMa3TULuW56PpxpfF3gqHeGGeUUIp+siY3y5RNir2jtcs03/J4M5xWQ
X9GSS03gzXGZmyS4YNafZy09in8gYMaTlxejUmDksPjiImXGVSHl2EQsc7qG77vF
/H2MmjyhiatNsQZ+cdThHAKGFT+tjhnxaqohBNHF+7cY885R7dsfklVoQ6I2NMfk
VrVA/UvZN7hKOygxp9oQM2iAWaVRkqqfAjYUhpRRr10t+DFyrFaHX8dqQFQimxgQ
lz1fwNhLrwpw9Ove2JGUxVDEfvVEIYwuyiun4lgKymcIjC72E4/FzzRm0I75vwcF
pnXBxDGhD4mSIl/ncP92XALGGF+/U91EBLkmpuQS3PC6x2q8W/WWgYoA6vWGRRrX
nMUzDQOsWmBkjJG9UhG8dneVyeSWX0SYiGWlXqpiJ1kivVzM28WY5DmAfbYx2CmL
7WSC06wzSymI1yFPPCgu7IvK3QIbFt4kCT0kUkYOF1XCozjcQANnKciOgJgHgAjn
eNtpgG7N2puov7uLL1dBKuj6IhXUrexY+K3Nd9E1Zg2csJNqgs8HnMvYXKtRHUwn
xcFMl87nx84z/6LvwW3QEccSKU+PDJeiYlHi9s0dJJKtVJmYfzi5lEI/6bPdCOUk
hqazDaOw3JF08QOJq5Y1DNjD9P4OhxbQnHWhkvn7jPymeWgcxoFK7D7YOhTR4v/1
UN+cfnKYPv8EWN2TmGSA3TxMuTuGFHrJyWqV724VdYavzfIGK/EN66tZXMPkP1xY
ThEquS39p5yzV9bamMuaSycpDxLQReUdKTYlTKru/vYF6XUgAal1IvF/ZTzHLAsC
WkGSnIdShbNm+SL5LZ2LWyFtjzBQkXQFYrOrL1kxDzIiztXmqL8ad8ftzZLEiJBC
Evx0DbpRzHZUwGlzX9sLWlsWRfntR2j2++wDe52nXXAKjdxRCCXbZv/cET56SxxF
Q/tttcE5/5yMnU8XDD47El8s22kCN2nYevaRKiBY+4Avlt1uXNObQufqH1TIiMlO
TYXww/wbcLBukM+ACwGv913SpAd2XdYgBua9f9w+Jbqb00cAiWFcOz44U9Kz82dC
OJ/gGVe/cyw/PUWgidTUSSf8PljsgEUCtgrAdNGJ9BLEwSd8IiXv7z4WMOfs7UFz
Zs//9+JwHcrkXAykOhqBXZ5w7Unv/foJUcK2CjRSIs7zCZ5lPpAnmQF+ZNVoivki
w7QzpRc31DHddyEZNOr/d5lVpPgS7RiaE0Xf/LpNpNS/ODG7YhXJE7qnn8Py4vIy
wrvUt3OMbFPN84t13uTvpznQ83rAtQ1MmeI7//guA37nbglZS6gxXGZ7QGJyXhZf
mT45LllCTQDryRndvFeOVe9Bymd9z3tnMrYsg9GDVeHF+ZVtXFpbC3yzCjWPwofo
UbmR5Pk9JmuglPKOW2ce+cVbfUCNlt9Sfb/kK0bQiOYspCS2ZXXJ2dZbburEha95
80phJ2VlZ60XwsnZUrn1NlJjNlIqsei/RN6vX4dhKSdNN02FuSee/LgUUtyf7xSz
DulOCf+8D8WO24xS+BpM/H1jPl+Plom3BdaYrLS88WtOX6J2kLWGdjpkypO+fBUC
6eVTlre/Gp3BTeIZ3qMJBpramJlioN4Cn3WA02bglPqJrDT1vKEuoEniuoFAiI6M
bfBU29ti9qALiQMt5nKkDNldpjHVAOsySB4547aaC2ZwmKc5hO0tKdjcrI0mK1OL
8T2ua8q4RHW2gvzqN3IHhJvdWw/jz7gLVVhkIIAIgaamYr8QjdJI7DRT9HPuRhqC
0b9E9SpD7adhQsfchVyCZjgMS8vYP6C9y/Q79czJ9vXT6sLDrMltokiRx0XzH4uZ
iBJtzGTQhLN2fjgrJmlAbpxM7qRvounBq/iEe4+NeGIOM0HcauDzBtMcEGbF/MiA
cVJbxopEXkzLwcxzMD//l6TmL9ALjyeqtTi0j4yuKXymP0z2vlOP0NxsX0fGjhUe
F0KecKEDCjgNOFQ8y4k1N/vmRpwq33t2mRc3Mrnv6n23+IO7KbK4hZCMnaUL9wXG
Dhiig+Ox5xeRWIjfMDCzocZqaNnSJYxlK2qcecf4p5v5dxKmReVOm6Qa0bPQjqsE
OEWQrFI+Ah8Wa/cB+ahHnEjynRbfFb1huB6kzSoIBxYLR8xFKD1MzwHT2G9EdBOP
MCgMrq6IOa9UK2RAdtf2AoRV1TimIky3xscIZ6Uew/Ibu4Yj1/ivOyihVhniTxmd
CxiBT/QKSVlC52RVRB3+n5uuEb095IqcbIGxGl+qlrIH09g0jSGmpt4AgHQJeeq9
Cb50LeNSsmBW7DMUM9++puLn0w5M4G+u8yfG0bYj/HfcTtT0XMpdEjq4W/6Wweav
VUe8PRd18gktTRS7oG5JU37ZZ8MmaIi4tWPQvsOMfq34p6pJovd4roeQEOsraIeO
kDMHBGXFtezW4FsJmjcfIUc4+Ix+EUGTdYQo1+7q6sZoyQyAWq3kRhAttlXa2W2H
Uvs3y+xL+tJNJjua8AZTJdpRrZcMZwsIxoj4Dx8a6aD0G5vIzL6Q+BXPF1SsR5Bk
WNXeziA7X6OugxcT4eBG92kQZAyyWTDHn2ZZzL8kj5M4f6F8lPb1HpX1nTenimca
MuX6ELtefk+CkxBikYAkoFDKfSU5XbBdif2h+5m9gN8hy8mRUFbxhhaEAFgsI9sD
RaVbYiuHIQu33838dspz+h04/JG30qpwEXLc1/0zdnNRDOuAywuf7yJyG+roNgsO
1NfaDOEYX4Z8HSnK2MNhQXs3xIElbHmrxhPwDFakLXHucM+glbrW1lPD9PKOhJMJ
MzWnkBp36lzz4bkSS+R2zGxio5H7WkpcaXw74FwCp4y16TtL8vO27caPbWrkGt5L
vSOd3pOnNMgOkAxoktrOeo6+Qt2xeT0A2eI/lL/uqGlGjDDwHS0WDwQfSA+Gwfw8
RnJkO4Yo0lEawal1T31go0+BoKqwYEEVB9HPKTS5oKEODSfChjq9L2Q7p7bNNW8R
xr9BeoUCBxBl1iglcP6Z7zZV5dWfmpjIT3Y8Jx+LA75XuAl1e6NEE2PErhPWX2go
GgmhonoShLsPigDlwC9eEWElDfp8UOJe7JgaSzujH51r7C0YIQ90PU1nZvCm4gQR
2Q5eFVZ8RJQ3y7nTaGso0W63qzhtifDrAmVeZSsFtjRhpTJ6jrnm2fOkLOzxWCRY
Oe7zp4ieaVqM29FBW+3l0TqXkTFveag28BlSL/nhRoOeqYBNS4Hw6nBI1YRmEy6S
EYTqryphLTfhYlEJHswn1i9QKAbpy1Ed8J3TNpYeFXofe0CuF1A/6Aecks6g5/Wk
KNd2/LsSz+gn3Mrbud5HmYZQQPxZTPOQMEHRGtpgdhVAVZ8CnXUha+tMMSnLc/tr
1Ml4e1qlWQadyHGnVIM1++K/DctV3ZwSdk1LjlXtmXEd1l7JCPsg1ETMwDVwCRuK
lvGttr/d+UaYUzwu+Dod4YWa33fjvSvtVVz/LWnvWXXg7GgCWiTv+T9/hpq4cAB2
vKukpi9tQ0hoImpjnQyAvImLz9lqa4JB29oN4yXRyT5EO2nlqELW6keZO8WLJ/zW
OPVmkv8BpZE8K4wMkgW9jnFlz98DTWwrsJ51eqKcwOsJHjFi0jqxMd9Pa75zKBVe
9zi9jnoqmM5bq1PS5mEOzFuQRVY8m0vVZ7MukIDl9MYpHFh15yQasKSHXMtvKq7M
igfMhHBYS5dpxyU/ot13uLsdD426uNvUhsXtAT9K/N6rVqeNu71HAQW5bzMWF60t
X2nz0DsOqMantlFjWEW6BSNk0rIoNiqOJcGmnBp8p4INwwn7/bYLr1YVU3EiUO1v
JSWn0CMpKmg2uDg8MCyQM/C6fGyeyENJvlcIOucETntb81ZiqEZJnXLvUs4ZMkSr
+e1eOu8JY1GS1f5N4KTrHZ8chbeLYidVd1yMjB+8ot3UrSWqi6ykl6PPuTitoxtW
aKf/XatZK9fTZuBVPeS5ZmcYkecHTrEvqywZ8pTLQyPNdBQ+DZcyVLwIUNRsVtHF
4KTYYPVMM67T+lwyXD+29AifeISCE4QUCJjzMFbS570i/cFAYkf9GdGcbPH0eqS1
vCiKz8uBQPiuzmVhL60aTnmY0kw5wilp3piIkhNdummtx9ERnEh2QqNjpRv7on/O
9GgDS/Z4Ebxfwro4xNcqq/dpzIm94gfSe0PVfUzvOszNXxQTcD9hUylTW2NmvJdP
92JExUesrNwS0nXynwaKxfQE84sItiExw+WQn91L7D2k77RWOvWKrr8F2VSBoYcV
HPq3U3zq9ofrf1T2MUgSVZ4Tfg2zwrnvVQYOI35GX3tXMU3jTpCIz6OcIK6xE+MB
31KIcyedylw8+uJaUMLloiwytKjyOaNxP0qsioI67bNLKz3AwpjeVmCs9tjf+tcz
IGaiDvew4519e1Ah8/OynNStyk9WLFs3oEBUKUK2NKPDNOJBvzTLpHI4//rRTN3Q
anpO8LJmLNKBs/ilknG9tC+kfNKQ5+y5n1m55ONlgN7LOC/DbtzUFveiLXDAcyvq
Sp+homp256v3Eshjni13fUGElTgEMb9GPmDRK2TWwaYshDaCiVixrVjQthHS7fq9
83Ic8lggMG0djY658oDv3wZ0WGl2zReV1auAAWaoNDmhWLJIMYvS42qxbrTg1tpU
dOB8d15NVHXGcdmwteFrL2+X1mXjnGM3jYynxc6Ptygs43mJ34DJi+RrmWQueHXU
Rgrq4ZGYfTQ/WRZRXIGXAL7eXj0saCKNgR7zwDA9T+9ipTI9k9tdwRkIjLxh4V9w
XstDDqG/5Zov5rzh3S3w8sct+7txfSByBpVmE2V7qY6ReMMUQPud3J6JNLVE+ZtP
NafC3b06a22D51LXSpurTSsCVfBsQuQfQRVAO0nabn0iMoJExpdQPOA2sGg0iPVT
ee7QY1yllaSwGF5YybdXmnramQbpbkgH1LHkhXen72EJFzWLhI20r77eJ3648Ihx
6ATMrj3BRpyIwfsraBuhs+L9wQaEwZaLEmzYXmj+hm22eAQlA8u7lTfDSY0zrOJr
n9SEKU7gVVVadEdpMJHGgWONUAUvcDDy79udg0hHqOjHZ+72gegxPAGCfI8Qr3V+
QlTmF3fl40jKVvuQyOV/67U1rg2i0jmmBPpdSmIDsxvlYvdugoVfBL/kFs8qGF0b
jHBKTyWyX9VwM3FkA5ECfrUemg8q9Lssg7ixft3o+Qsmzsre7ezx+LbVqSpqKdIx
6kaGXEByHFrzbKcVGpKVsoJmlnbZ4oUDOsaamHPE3KyIaZl0GYc0jtPJU1b9wVHb
B76RNFoLcYiG5hw5Z/J3NcDnwmdhdtvssRuoJx4qQxgH3RIf/R5DlxHSuElaeN7x
Mn4G6PLiMnz7Hqxe7PIY0QDehb5fhdkYeyW8MbZOV90i5SriLHKc9/2vuVK5oKHI
rA5zlIlJwUNA7VjdrTckSAaBlUAwNoSw0uXGbeJZEIATKaZlelPImnTOvcXgiobE
MGjwYD3C53rs1LqDMYUeBLDzFz2tDiVDKJOdt53J/9QH6U6QkvkynnectIDNadQi
pdr0xw7Su4F7Xaa5ZL3JP4b+Ps8WS0yu4eADURhWgU8JXgBYWU9YtYb7lqdzi2/s
pAW7Z9/8sOCC8FJ1mkX4tFDnNUqkA46wpnYMVk/+vkPYq3GvSK7ZkPJSVMwXv3Pn
zCqDeX3Z8Vx5vR60UVCtKWdUZOqvr3kvx+4v2ASY2vWFkGMjKbealsDao8H5K7Vl
f3awh+ocKezT9mnTn6aIz111V7+dxLX4KurdKk5vGOjzcrLLabnWn1DgkKBaecDN
b1pBY8IhUHY5PQg8FrdOOnZws+ibmzlf9VdkiI4b9gmGvSqj2GVD3Di2BCUNIgFq
duAIWyiE+xHiavX2ffKErK577Rqh4uMavnDrkR8d/ET2BE7JL2JeUnrL2lf9/r9u
yApg76uay/UBfLWXJU6hoI7FSqgYKG8Tfdne3ICG0iiWCS8q36nzukQgR7iw9936
YfeFdXF8dDkdFPOri2FLsipPDAasNVJqX8lmoWGikuQOIAO4EwEHASfdj1rPJOHK
wO+znDSQ0MPBXteI6vZB4wUIiOo6cNnL+brBFFrCRUZM1XGr0wibMAFzl/KxAbvL
LhNWcdxfK0OeOkvaJ/ahS8QBJJyd+5BpFZEz1VTsuo6lrzBrOuCFVRthMq+YQ5FS
OfLvSU1Dqgpi9lrcV5it8eRcF9ssL9WmEx8DGa03qJ7QKKlYd5xiA7Qw2ERSN/l2
R+SSO9k/uXch3rp7+ulAH8OUFqaC1gBybgg1I8LWpBvjxqtClbHetWpo2W93wwqN
GdceJ0Y1dDfAHjo+wuDSj7aGBAm8zb3Pg+NHPTtjNZD2H049jbiECk7ibqXPOMBs
PX20ooZA4cTITd8oitQ4uOA5znbT8d68f1HE08rL7h6nzzX0SR7grLF6YJcG4JG5
erIPeetRN0NacoIrNXgOlBkLxoKAW5bmUj4Ti9x2ZPAjK8nekevUZ/BdFbyRfX9L
zFAVkwTpH+nB65X4f1qZ2VNgKmiRZ535TlosSvXRG+wYPsdXiykcOAxHS6GtAgSD
hdNYwRW9bRdcZ48tZl2+1J6ns6qWFNAPKbvnST1MregCU8ZSFKReOVWJX6wukZB4
0NDaQcwFm9aAHq6TSfH6QiP7u9xv9OaiWSJfgexZqGAqU2CgpgHrBky0MwvKHAWM
5yIQ3zDy5AsCZ/QZBMioh5XH2hIk2zIUEbd+1UPAP6T793UlUxegPmr5ZXOCbe+p
wIHGuZFHJ8Kd41aGtA554/GiHijQkFUKoqAsmDhYvMZGzMrXtQ3WOnQUdL27n8Ao
GD8GL5b0+F7A53OvBqWSaOrw1GJBXciUSM/pglNs1iwd6+QdOFwtPTDXtj3D8mnS
EAmCQ7mZHixZucEIqgH+aDm+tcltdzDYZda1wcVHwCM66IvaZs+P4oc3rkJb9KjB
1fd2T31Ui/lgTV4N9pC2EOUodJ0RSqk2v3j+gG3vtULyMYXTtcFU3TwKhbA62B7E
MvOtvf+NycQcS0Nc6vVs9O4ABLXa5vTjpHzJfxlObh115uHglux4csyr/qzxIcWz
WjBEIdS5lJ30CLyk7HXd/tDzaS76djXB+Ul3CsHAoL6aeYEvqE/fs2U024TF7Ebx
znQA0oAx/CETktPZZefx+0cwbTHnr7UPCQ/ypDRC/xjo9pm81f68henUecJ37Gl6
4xy0DDVJOVkluG6d05WxWEGmSdkrFnhHBn4EwcaT1xRxelCZ80o3ymQ8oTKRj9S+
gEiB/xPQXWATcAzBr1YY29ALCItPETlOGo0UK1GgjN52HKbi9T7zoUMSPxeL64Vq
eXp1gTNlDddJWZn//MAXHM4qjvaljmzRgHRQACxTor0QJnCOeutM/MFRpEilHtaS
M9KfWZZMlTv9QmYaTs1Zoqi9woMTTaVS56zQHQq28gsvXbHOkPbKHFRSOH0eImef
GlresBOm/rg84sgD5INZA6Oao18jGML/f8C7LGYHu9eZhmOxAiu9bVuBysf4f0T9
ZaVm2sgUYLrTzAwa4PskFJVYw8gkX7Wx0Vhk+siJMItZe43qfCmFznGyCXierM8Z
HD00CdVuQCyv8dnI9yIvTq299Qc8V4ildyxyAn6Xcqo76OtT6qYpvJQVWbNklefF
vRND/R579zRuMjJr0oCg4rzET7MDJVqWVmGc4t7/GkRiT20ae+6fSeVeUbsGWYi6
44N+KSz2JXoyytd+BdPycg/nHdHQizoR8SRwFY+gW557VvsPnd9UKKiz9hWFRjGO
tivScU/mpbBbU3vmcwxYPsl8KGq7YN1uXTL6hGA5komc+IxZRfDivJL3NhvSzXgF
kjkZtkn7diFMLVlTyqdEPuupl6MUcnuXrbj9iEg7o9BnFC5oGETsbdf/7TGH3nFh
i3OXyvL/TaIOyKZ/gZNm9jmQSif0XMie6wRM209feg2yxsXzz+PO3mzEumROrg/g
zdJyhzFXzBJYi9OTwUojA2+ke/4P01DcroQlzAJlSU21jTTXl3EAIUIbxwLjLS8Q
/FFkGTTKF51IyNXXKsRCAPlVZgDpEQOcHwm1bKQlFlWVYoHhDZnvGEsC4oG4dpvo
WrvVYmuY8hVx08R0SOnePwOXC2HNh7qxMrceUNx6ufCJOE4EtXVW3Sh1GlDQP7G7
3ihYZ6u9JevBsSSLmvIPaS6q6VUWBGL3iYphlgB5XyEZMmxELrflLxwlK8n/Pz1U
NWyNiRHrkEljeThVkI6boA6K+1Tea6findMJ/qV2JqjMFfCs3hGahvLJUlKuFSXU
bZixxuIcy6udGLZL67Vt7wddJAfO7kr0T9HWezwazYmgUY29l2Kzm9SUniHzfsYd
Zy+Iu4lqlOs/koci1nVCUFx93Vums6rsKifrYK+LtTmkQ0HRtcXzXLfq67iXgQPE
CF/jaOrKgbOdjFtVSak/ykns904lnk5GQwLMxfOuHl3F6pIAuMsSH4wH0w8Kf+mL
znyJtl2c+w6ER84eQHrJPXi4Bzmsjk40T+PgEvCnIzfs+Tq8osnijXGwSmJ/ICn/
rZ1LsNiwDO8kqMwnapVHoi4VHW/s/zs90U309H9ACVhgcbCVK/o/CSNxCtKwMibe
qgIDi7TL+NUl1nZM1BWfRevo6w/+NFipndjxtc7mxrUwNN/1+kBQqnB5j8pLiQpA
vSOZCSsvVhasguN8g8gQN+VVdWU2oDfRYTLADvmDN72oOspBfxPdz/y6/aBlIs0s
AT5NO2tnPfjqqQaAKJKjvHiQOV/PjszI/AiH5eqTtj55CRw9uwD2rlmuGvlCxRCw
iRZ2tYNtiKf7OEWrV3A2Yr5kIlyS4IUlpqVbhF6FI8MoXMvT7snZTGzclHUNVAVe
nee9HEhZHNZBFof7BXQHwZJsOIYtfVeg3C45GsfrSkSxc6huKq5fRc+rRPuOUiZW
oC6lHZrf1boMZRiYIB2HbV1dG+KGBIpGAXBkRsQqj75GBHFsVDqimTDjtVnW7SnA
9ozTPOYKSWsnYB7cLFV/WobeBcgsySno5ZCyhN/9YuGpwUMMNtBQfNMriCwqf62b
rYauMr46sLJbEwT0eS96zwFrAwobKQCyXKhJoxAHEExHLh3K7bEqWzkhpUvjkTMH
LiXr+CCW37iimp6C4bmpn5b9b372JQjeSZYC2EMm9jizi0KrKqE7ruyk6gBwe/lT
zafqSIiuiiA0+Se5YIEE6pMO3rpVoodfsSF+Bg+hzHUtIG83vmz0JNMeuoZuB8fe
If0GZREJceC1ufjP88XVZk6TbDkoxCh+4XfxQjVT4oTitsZ+v1Nht4V780B0KXBm
SEX78rPbpyvq2fjdRyPxTFCBVlz8Ql8jg/NU3vbCyhXS9QacicbGstpoRwNfOVOY
Fx+73h5xzEy732M130KyJxriLAxSstb1X7DmDvYGbkspklZ//YG+Vik/5bw192bL
gZcjcgRhM/xnph8jUJb+VDOvQOWZRNyMwz8SuSEMxawu8sDiKootsuyGbFk3Us/L
VPyrPoSycHMU76icfQjrkO3EPpR09X3xxHfkBxWfuHuzaTyHK8mA4KZ0BbKFQdmW
ZE53tPKOCCrCFBWdgTlxvTyy4R+zyN52YqixcZ9RRsdy5FN2rhn4yjf+uktvcY4U
I5biC73J4H27Dyr3DEfQmXzm0chrGvrSgZeehuXJu993mwSFh2hh5y/Zj8UsW0td
DEPheTdm7E1MWxmnuTykPWqtMEvIrWmjw94iAYQmiBE8OYIpnrNYhnS/unPX45/w
papmgM+Gk3pYsTtvqD52EpjjzZRj6twEu+8ukmdxUkPMizuVrNrLAwsBnoZYqX4n
mrL0BYMI0UB4e6LtHaNsnOKABv2T07MmSpz7bkUOKNlfMWSCbOdzFTZMuDQsxSgU
wAEYgB+gMm37c5dy9hWfTTx6BBTu/XVy/9clMPQohhQb23Jbpaef6GmTt7Mggs5I
YIvDtca3XVnK6Wu7sYmA2uJ7X8ejlgqBXt93QajBMYgZXF0hTTlrgainA7KZ550h
by0pL1NlDNE1cP+lIQnH7DvHsWNGNeAAPN0Y8eQj1b3bp0MmBE70qNfAmMPMXOBV
3S6elmrZih7Z1GK7rwh5fEOxRpLzHAW30UWH/Qq2nkswdM08LRaWvNoNGMGRfjA/
e832HRulHVHAY1DhR75ucz2z20jcCjAMKHcIQ0n+YVuA1rkewlF5aDr1wqUREO0T
cTO50yZ5g8ybySxELEf73Js0n95yEzxvbcvChrs7IH627mQESHoNcVbU21v+Mqi4
iIwOjoN1ffYVkYLxIRRYCpNXI1kXifllJeqZCVc+MJ52QIP4MUC1fNyhDP86fjbu
MchGJqfZpNHKfTXPTt8C7MyZ9bYCBrJ27OaLrFR4dooRq5DPb+/IKwi/3mrpBcon
pXUYkwoQuq0H73GY7mqKWaLa6BKJ14SATmtgXN76uPa04qRvEw6wDFN8Vsz4WoqO
+yPHz4M4+jVLd5og99UyRCZoLf9NVtHN9X8ylCRDdi8nOzNlgYM/eCcksUNiP2Z9
XjBRzV4FgsYVbZhK1NgDPSY0aNGzRJPfHK8zIRY8d8bcs/qK4+S5q/9wls6IBwyO
TfUXHiXzgaGNaV7oRt7m6sE444OO9Pu5f5Z0EGen3nz5DR+7Pcq8ocgp3tZNwphr
KoR5a7PEsuKNfgK43HIX6lSktl3OYjTAPlsSwYnqm8jOyclTtx5+esjtCr64ohDq
lpHFoVcPM7biROFZDE4yVHna5eojglAmJxoTXtOGhEprB28fF6B5YWDa8fGp9Dsz
wLctxq3TRsUPVuDTp1CUWLAY1id1ewkchepv3yVkcBeiJus3ZeRAQxk7X8UPrGvX
7/3Ioe1ZfXxXY1bW5bTo5v0kd44kx6rS7BjXERgqDyuz6uhMcOQRQcZQb57lzZwK
0hhj+rJ7uEI8y5Pu3qhtm2ulnqkEx5faa+OHsXfcVIp9LuKMAb8NZs+TpOJIVpBa
q/zdKvv5sDmYsLMKlozqFhMrr62PpuiRUFTuHFmztrE27+m4XxrejocOWaTy6IRx
BrPssm5/4+14iAo2DFkA0uQ15dlwwjBvvDOUNN5LfF6gfIUKZQl8HxFhZEhHqZyJ
s8Vug4yWJN4J9EeTCHMfobT+wrSG/ws0gWWdYNo/SOABuBz6cC9dIIXtLNefEf55
YBfFpsTyovb1wyeHYLkWHYnMe699Q5NNCxRv4KKntk6tEgcjReBwUV9XMeWM307l
eRjyxqNQfD4jDnaGKZlAebJ096raVpygaWFpy1tjYuy3DRaK6jS7EjHdmPCY5mYq
iB2ZqKV0OcJnwvTDF3Exy5eEzl5bg6SVx4l11+5Cs5hb8y16rpMAAviMG++goQKf
W6k7ugrbkISivm0rLH+IWeoriS18SOAQVWVs6Ti3VD7U4vEpa+vtWsdbQzkf6km9
A/rieUB6PRNK/crFF3EqqaTPHgyag7WQovmsIPL/RtOjsYw7GhX3gDgHUvb9CByT
nnGfXB2vEvV5tceFG1JoFAY1fLzmPCG/fWuKSO2uZwQIc/2zLRtMmCDFUkLr79ho
pCyxC/Hdsn6FmKKNdZCuWn8KPwC+iFt8rWq2tp//Q+gxirViHkVOXvCLDjk41Pqa
aXzW2YsOCvBV2lUPBtCYDy+hDw/yNIcIFjxHHvIWp5WCjGYR1p1aD3xsCcskZpLT
SU2zlSk15FvJe95ID+kBZi1vv8VaIXCe3rHGhWulyXD8aaf05jmdR3gOdCMvR2Am
uj9nj1GE3rrqf04p2mbaaD5dM/XUjCryWp6yHSbR2hxrdCo5R+1IGJsxh9zJo8sM
9f5vMih3TWJLzFpuvdKPDd7F0MKW+/3zEdq7U31GfPzl3rOYpLz3YAbEvJwI58Wd
dZcjmT4ChtUIrN3TUFxG0aJAQzxaN+sWo/l+jLui39OI2dmGTFcldqP8ywsCzryJ
pk/8pJLuDMkQmzqNsqOt7BSQEM9XgTWu0mcnmBDQIuR0TCaTw+VPZN1bcfVcIE5w
7qa5v77oCQVie9ZGg4htOR+a+zlppiWSYjHp4z6zeDbGxmTQiMRfysEcpFROda9C
IZ1h5qaJfHDCPSbG/hr/g9qjtMDrpf2Y+wRlebxI4pXkQwRzyHhLR7N1GGSA1Z3M
dVhwjV3S4zDmUVH1s7Bvfr42I30CWPDl275C19c1XmlCYoifgnxxprJOBbqFeNCV
yCruZ4NP93ft0LxugBzxXilX+OnpH3hmoae1LcWfyzjlVNF7KB/8pHnizQk8BGJV
f6zucgEqVQMK0tXM0LK15LXwnwkh9sVNfJmBoGuowhHdXIz6QHAfJjAreOgjs51Y
gGaoXkL2ikdNqRm97LnYctZWo7R/I9DPIgvQUmjbBlP+udQTjLPSVvp69O/79aKE
0WTxysh0cZMVhNT9uJd6Fqqgl3zW6gRlG+oAk/b3+HJYraePelEW5O0ZeNB0fOMW
m6ICwLNNrL9PRsosmHzTG60oZjvZcK/r39ACjCuRtHdtZ17b5e0NijjdHKxtu2FQ
lIz+r10qhvDWJxjDIyz7w0BjifsTghLb4UixW4vvcRcJjLUoheeuA5JeQWgKOxtP
mgpXDJgV1On7ID+SQq9jGmGOyj/pqV3r969dBHH4+ek/JSn7zvVnxpziVsGY1Y5d
D8HvDYNb/K780YpajTYWFN1U0efinoWpWzmuMKTRnqUuy8t/Fh0Pd+OZysvQCpnn
KRRaYRoTAagS67SZAiWb2qweKMABJEGh0yjIbAroMYouVk4Z96siWbz9DE3ZU4TL
I0+93sHJ5Rk1uLU/cVYj0c6QI0bSv+FwIwPnd6Q5evNrCRg8iJkYaYyN8QNsTftz
s/akxVkRVWLXJNeTu+HqodWQPUDrThNJBioMzora1vPZHKcg2An77oqmRcl65xX3
KW7sAGEqH0y5bffOmj8azOns3J6Kmti/nj7FqYUEUhHt2xfJPIOdXeodeDO1ZeB7
yapLnSSkBr3kcSeMA+HNslau/iVpGM5dE6Oa8d2/7qrMHsqSF3sHgMQzBqf1Su77
/Hh3VZYc4MBKdr5FJ2IjCsXOu2aNQB3CvtuwBNxZrdhWRajwJR4+THZczI1qGfJo
fb9x8biq7t0RYZzByr51b+Mm76MTciIB54/swmJDgiE6gg7M/QAazLpejbfbjSzL
DUHV1dzwJ+NOkX8Mq8ZzMszGIvJ5CM36i+cZS/ggYGg+sPcx8gq8yTRJ0RHFC4pg
9lMGpV5CuF9nqq9njaSR016FX5Svq+AXYTrcoh5egj2DIbU9BWo7o0Zav0ZaQW82
ihq8KCngm1+GlXOlWbTFlA0N331QxlFCrQR/iW7/OX9CwJ8+N80vS+KfJe9rNa7H
cQbRoniDdBfo7d8LzvXypegIf92fLgI90AkhUuMyF3iPEP6NCf5dOmYwmiW9wp5k
x1WyV3m86Lm2VrP4bqHE51D/w2/gVm6rj/AjHt0hlezCrCvWfQBJAQLy3r3d+dUB
HjxUo1AG5kq4HxWJZ5SGkvEyXkqT34pC/QnB+XbTk8GBv8daQJ1rCNw3UegNedzz
JP8lvqu/Ee4RUms3ioM8JtojAaeNU2vtk9BlEM4wl3U0DXHsUUUHmsS92sk9oTbc
HaoFe/VQmvaoZNBWFeFObqncvjZypoOPZAgpFWV+56mL7qWmd9W8Etty2V7JghP7
eTPL5wMRmoxXOMfwnAQJUry7DJn5op3ggxdZb1QI3fDSYact7gGG2dDgkOkubQqQ
cWSsDoQGWhtFyMx+t/Ig3uPJuAcsl9OHGwrnhSG2w8ZO/7dn87YTwiuqYt4A1DZr
jpgnNHZT79ZeXhWLTnpFRP331F+syaiMJAu8pBq4g2kQlg7jn7xLiQxaH5VAEVK+
OUpSu05E2RSiWsQWKkzU9fuigLilHwuiJShyT6VMmfrmONxyPGTebdD7FMJ1VkcC
cVYx76LkXR9O/pJm1Axfct3eJCmkUFVohSBThLKGJBeJcrx713w14GplqmKVGz+3
Mjxt8muBPnGN3dD32fg7rwdxn4+cZGiPp1KzOHD3svW7Ii5dPweY7UPmH/Odc+r7
wdf+SXadAI5eS+2Lu8Q+tozc/UIB08BFGSG+YPjZKTYakDJSyu5yTrfCi7WaZV/4
c1TVvfgqGMcsua/1H/do5oB5zQWa41+adsrb0gbGCZS0hVMoLKdHKe5ktKpDXlEC
fdbeDt4uueYGjSlKbEdebwUbHNaPY3nb4zR8zz4BstavKGc9WFQ4xOy1WRP4Gn8S
UU47ut3ACtGrNKmjmgjdFhDJTToXFyxo6ufFV7NOqK+HYNKyQw0Etg3VpG4T48Ds
g9UMSmF7BZ+Wg1X2M4xn0ODb7lvBez+5TI/ihASRBWAYOrJ2Pjd+/aQxXNRhCs2h
m8bqP4CNB/HLkQaTjr/YI47+29mR4jFGAB/R9X5wFxUuWH4a6k4jdMr83Ym2r0wd
uynr4d+8+PG9saIQ8YmbOm0skUfYMs259Va1VG3RaV2buSrx1jB5n8FYhcn39PJH
jDmlBac3OmotV6BAZC2ewFusITbuOqYz3gKWP8TeM3E4Clj64WcI0WlB7sdoqboi
cdVQYONcIVG7I9PNMh9lV0oEZSc+BMZL91RucpEoAjXvWlsHgVpFSjzTtNf4PB6Y
05zyxNJg8gS8VC4xz52vLZ1qc+8LQ85mn44ugYM8RM1Rp5HCP1vIfiFUvfJHVo+p
S4/JrH/eKLOmpXlrNmlU68/D3tbUVIOWukfp2FqZRvDIhqosn+Ix/SAkvYpPjDyD
NMPXqSYBRK2kePeFXfbFLETF8Cwk/etS+Pr2IvCDRiPaxLcIKo9cZSdOpsje+JuS
zrPleiImaBW1qBZfTBIKBBq/Jw/KjqVIL5x0pUBWyLDvbcs9mN9xpQSZ5a3DvVQu
NuB/Axo6NqQH6RI78pubkkcls4rsGZ4dxEp1GZokoJ7mEMyk/Ug2GeimOch+A2ML
AC+UVMG2F7xC6nYm3+iDftTnX/Dd5ZtskTEKtH3MLYW3FmJARzMnRsvjMBZ2Cw04
1padNPADMhrzDE8+ox8Kp4JPDbjjMskdLFIj27Tcuenz9/vbBorYHLd+F7aGl/49
dOvLY5q0pFW6/YMgCCWfzUqeMfZXMn5E0Kpnjcm0nWKrZkX7wSUaPsEHavsCVJGE
QLRlYplCO2/Q0whGWfQ7AqoTuO2TGWdHjsl7qMZ88mmvxb0q3yiIv391hfRizfLe
LaqVVc7DQb4rq+PDZihsxaCkF7RIoyk4XkyhqKsOBzlZSc/jtZ0EFGtTto+V94uh
HQp5ePjDx+gB1XlcMz9MAqDXez6cV5gEAMsVQxdMCMEp4mRRJlYYi2cVLUfrtjNs
7nxesyrQkt9Dc4PCJBptzWDTkei44DLBzRbfvdU5zp5jFqFjOtCQzLbDAijAQXZR
sm7GOp64PQhd3Obmnz1EvleHLHISV3+b3FhwQQOEg1H5GbEr37QLf+SsOM0qtZR6
Yi5GMVf0ngWGvi8BOBN3VBQRZL7AZKaGS1DbEi1mShJjHwvI5SXas0p4+1clKIxV
a9vTeblpMm6D/8yeLoZ65HW22zntv7BEsGHSe0BRjW8XdQYYN7SP1WNFeieVkujV
SHKIYTTpcDeizb0LJmeJ1F2HvpBEwqiCqh0Yot3I0x9hNWQxcAo7vcSTnBSpIZ3E
3lzn2uhjpzQNhGH9p9o1iajS7aolLoqAu6/LHs/+Qli1eQTyg0xnTerpHkGpyE8i
pnsTK9IbsNKI8WazdM0Dig0uQQS3bGn0WJTs0khgFjPO1cz+MtlO0lAKKLKnSNRB
0HDRkc1NtPfeRlAbNbVV+eCHEfn2Ma5mGjmPHUfNSEWln773+EauJBn2a/z6ZZX1
gyw/6KepdYHxv5ls9nOtk+04lTi/bH85Nk16CHDXRVxjTmFgx5m2Z+GO3DSkHlne
mFvYutKg6uppbluXxvR00JLqbOKmcXrPN5mYkb8Xrug7889losMBTqiVengKE5SA
aHtELcZAKLBl3t8qobXR3lDDtKK6cACrUtefo8C4GYS4FSfcapncehp8/ZOQ69DZ
JYWas+djfsmZrjAaqENaJZRyn0/mkwqwKVNsBT23XXfQaX2zKTQsKJVMSIa9uQ+t
LVr2LQDK5hfHREsRCB+lIncBqSGjOs+mmIEvWJy2aIRswn4J2/KtHqwa8WQuSSK0
34NWiIFEkzl/fyAlWMlbZMV7gG0HzWVWbXHIdiTY8rVJipRwbgUHUFjYWVIVgX85
fVe1yLET6sFWToaMq8/ZyA3I1ikHr4BIXUa3YLRATuucLb0WfX4ZZgrKI15zGIof
exK2uN9FowrNtIijDf6HOWe+xMyJuDV4NQEuVdYJ/TkkQVADG6N4haRTZKN2Oonj
2IGIWLa0tU6uD+yco2BUTQ2fDrWmzOR/ZnHKMSHeICogZc1jMnMcMBQtqQ8KCnw5
vSF2yam+2lHd1ewHHQtGlobzWyjZKquxjvjOl677xCjYEAeGncLhzk28qBC8iXyY
nx4juyn9gcIG3PU1dshv/FDLDHdLzTzz/JI4CSY7pBZ+JvJGvcabhCJcFd32xVyf
NHswahZQjJNDoF5JAcC0L776LmEcrysSRjzdgGi20SCiQlRYHPb9B3HRim5roJ+m
aGJlEeSaF/EtFr6VRKR0w62//WDf1cSOCiFjchPONGWzlcYQacB5Emyt6sxwLw3k
mI+4V8YESZ/HFcVncbrp1wYwOWVzngxVEJW07mdSDDmu7s70AzwdwH3+ZqPRm0ZX
6iUOaDv4T8CeGE/+RJ2O1Vo5LJmAaSYTG5P0JdfNKEZ/P5vIWhfEqs0Hu/5mjKON
FiF5dNFPdAJ4Ed2NAvWZf3YQGUElUje+WAcIiu4aOGAwZGqp8HEn0wZt8P8rlynK
8kmnTlqa6YSi72bGk/w9dzJiX3QOZG57EP1LXth1HJz2jHPXOUN0rTeiuB6/WznC
1/YnHthc4D/6ff3AWo1vKbhuhtVTv3EJfr58hfH4ZMTFjQY5JuNmUF4EBWeqhec6
OsjztVDHSoXllqkAO/wM1XsqbfbhD2PdH4ejfzbuFPntdrzGG2sGYKoogucPu87D
ehS1id3qhZn+L+UojK+Uavy2RSK26OIPaGn1J4CQrxrjxrYqDdElUWw32YkQagFq
1vVVIiZpXUc/Zg7PlDgQkDoOh/Q24pHsbGvRwVkXuGU+wFSFVupjYAxgfbQpYsnx
ViqStVqQ/Uye1TIq+eeTLnKv/iarhWU9pH2fQd8XuuDBMyyzwkCQe2Le/RxH9g2p
osDil4nRFVhD4kuFXdSf5fzCJzonGu3xAILHdy/sGf43M9D/S0rSAis+4sTQA2UV
vUE+hK3d8hBOVeglqc/YwYpXSz7QRteImtgtUFjm/rSB/oqsIf08k8b3lkDIAAvU
fb1c0SRXyEQqHbInUu16tBOcoJJpjZVg6a/M7hkEj06W14EbSDborQJS1WFW/PGE
Rt34IG+RpkEb6vHHYPL6qn6YjitHW+l7wjbeUCLqnLb0ryXTdThn9NupIh7DTywP
JAI5eHhKqIIjoFemeeOqm8nYw0L2n5eI91WjTN3rPNHYf5O3nB8HHy7jRoYTQDgx
HM7xekfynsE8+M6jI8EBzlZIaCpbeKjsRubRDV3uE9/KUgHfz9jSbiq336w1o6f6
DJOj9ZTL14mak4S/cse6p7RvPW14jsmbG8kh/TldrhmP3c2fUDpClL3q5NQk05jo
H28rnf2HgCaTN8QvdoBHH+Xi8cMpHECQtS2QlyxbMxe1gAcxKr5W/w42VICoOzPQ
yzC5wYJ636p2t6SDT3uimgggX+HeK2T/7Sj8GBNLflo5C8MaynpiM0yRTyzkKzjO
5hZT/aQJ/PsRQ3X0OzdE/9Y2F3ZQOgfsoezYrRYm97qIwqT4+R2RIFmStBT70Moq
gdjcqyxunqyk0RWWeeZxoj/7yiI37G8llcppQkUXIO/bocgstuSi3W5nQc55EO8Y
04S3uWx9kjth6mpMmb/zK57qtLu9/BN+dmWbKM33IZABKHgqYwzRk/CpUyKDF7wu
UnawCRZ9zy9ooJwXv7bRmBc4mZBA9TSDfZwAa4kX5OurJEEfHgEz1QNZDTvfZgzZ
RROQvmk3heHp4IhAc9W8BF0dFeFyjnFsHJTJppwh9jYieqJ4tW60K5AJXMzLQVTw
sjocaLU6l8pA8V4X1uStZwTP7hbU9snWewP7mLUCvxBlGd5FMMUJ7SjkR/j8lWCA
zve9uV3dML800AzHW1Pa3YDZMTGTqAXAAsfZB8rnbqZAHBQB8EzCb4yY2BGvC2xH
ZtdluVaeQ7wvH/8MF3qKZY9kxi786LCp82+Fml7oLX1DGK9h83wnnbX5YLsr/gr4
+rrp034gswYl/IWKj1MRYwlw9ddf/iJKuHiwnZcmQ+AqwlA4L9RRXllT7rZgdeYG
x/j1DxH1fHkbiamYFW7IEhxBstd1CJyf0KyPaI7ttW6CzxWxDRMcl/9H6jmpCl15
KhgyAA2tHpjvmxMG5mhM4A9BzhMuGhprLPAP7pCBRgA0DhPr61UXuRd8wpyQm0L6
wCbabz0Ggj5c/07G7dgyul7aXrDS+9z+9icMV8Kj+4gvo7mh8Z5LnNACTYRXdseg
t9PUfq4rxCMXXTEkK7O5RC5JYrhxSPqzoLcqB21CtATReCAZM15UWEO86HypXuT3
QiYxWuFAGJd1s4GXRflShufKe7y6t4wVSfI8fAzzBZwdj4clWrU1ag0uUxb9QHlp
dAbeMFoF7j/NVH3wWBlUlD2oGkRto1NCwoUw7xFzvdcX3v34wUOSxeB7ERjDEL+q
Mce7KjfM/G91oaHKTBMEEbwSnhpsWyiqgZE911BYEJrkcRTTsAYzuKxHYlhqRi1o
G4KdE40OvvN/ZIcM7fiz11UvhGGDWLMIa3kSlBvbRlg2frLIuINC9GPah1abuTdI
hoMCc9Y8MAPoaxbk006nn00/oTMW5qpI3u9NahFJSgB2AiWB7gCwjGJsNlMGMzyl
bT3RqjwNbTelhM6moXP8ZcP5To6dQhpKuxmhoZ4zysZ1XwhlZNeGMFXDA6ij9Xp7
PC9NoWK06EnDv5veXbvcGdeQokSz3+HvDwawChWtYWTeggZBGOe+Lufk2yyOs9zX
VRV4GOqgxXYBGIhM4bB/d1vAlQe9Z6CME91XhC/rgxmcpFDGXwpfocr4Dc1dSBlE
ave5T9CL5ulxOzY62vbC1Sz9c+8vrrcHQzrKa9YrZZJv6p5xl4MZMDa8RN6wghrN
EPtSV8SEiNec8ZosehqMrwjN0LeSj8rBsDy9modYmktZYYBmOzelR6Ioy7rn6A4F
4/UqstMCA3hXJWtliNUTZT2DHU70W7zPxcEbeqQ/xKku3S4H13xAHLwJV9vG5U30
HPoiYJ4L44u6SBtzoJYvALWfysHjXXMopfJrwuJbGOkJyvGfx+fHQo85TQFFWzDv
fDZtyYVqHzDveN+RCaTPMZ5oyrPqXEns12g2PeGxLxBDyuTYhxftmzr7QwhRlOZa
3IjibRe5XA+9CPi37JZQytScipaoySFYoc8Hq3ZIotrqMoahLihMSKj0JTdNR3XR
WviPA9TvtEqGvJc7fDgt8A4zgw2MSwDGefPUEg9sV9xVS9zKd0nPWPPrVkVldZyX
9omUjdJu7pmI5sRtB47NUmThRrIWdYE202hZsQJmfsSGjfq3AKnCuSFI692UwMxr
DOcTtXepwe0KQnz4i73pIyfMfNu7zBSK+tFa6yLQuUDW81KCnoMfLMEbORJCl0Ao
pBUHqoxWROd1ET9ab/PppA+s3nd2esbBkblvQNMBthiuX1/swQNB1Ea/CqyT/DGG
qkS0mMvYT5KTo2fb79I7AaAaohkTEp/XXHwR6UtUPBliJH2n+VYoLbB44911UV3m
28ep9qrv3EJ4ZwSq9EWhqXxlusohGZ1qumzv7q3yBgm6QQ4FD7gevODol0V+4Aoi
dzJOija+PvfM4FNONonL7nUuwx6AVuMUqCSHhVQNYXopB7DDgClxPOu1Un184rhw
mbwZuGzPXji3VReUogQCYs9zc/VbZEopXG1pLMuiXasOsRDy4j68O9LLWj/VsZVT
/YozW0580VrV2f9lW4xGNAUZLCQe/Y/v0giLBOfrjGA4Mit6G0C6I4sIqjGm4aNn
B8VVSfAv9WOLWXkcOhd93Zl/UzExaRoiLVQW1gv9oESob4wt1dPyXe9Bmh/xbmfT
kADdIPULRdCh4bq2z2sWmiZPgbOut6tuNpTYswrH+FDECkJ6PVfRVnZ/R1sI0VM3
4dsG72IHvS0tg7CwjR3pswgmuqjim6JxNl4GTUqlBYNzIVnFz5O2MAO4Uuceur3H
er/MHVDOq5zgeohJnqgDBQPNT1DCf+D9vYibNOUJQWFZTcfBupb+ggGNFd9hZgk7
sG9aRJUG5QnQZQ1+kSQZiELAS9PZSgKDuV7ttKb/MbYG9I4TKMrNXpBecNR7H6eZ
eP2BFcwICQ33HJslUOP2aGX+/663RCKEPMLyjamHwKuSZZJreUneY/CT5SdSkVXt
WOBhzTqu7Xq+wN9zN3OXGH85k75dWUBBribXQfbB6A2ckcHEuD0FKoUbpW9Xm5sO
V34bnAj3cQi6NAIP4zUZFaFEq8+BSfmDF306clKIO+Air17iKu0NYTrOVcArpWD5
9QwxqNf5V9sI33Ip+4ITOsZGlfRdjYiP1C+TGRzBwuSLwjNO63W31XleDtDCDguQ
qAdZpAyz3ne9KmF4bB9zmI41kBCzpNIn4Xq3DmKdKEOwG278VIthaaAo+K55/wtA
iSpVUBbtlGQvB3m6Jzh1k4tbL8QR90W6Fj1O0BQFrIxzM+uptycVHltP2NzUDbAb
buVJYUsOTNEc10m1BjHO2fc7e4ai2inyBW/R9dsEKFgQV8pAmtkOuaRfc9algc96
50MhuCxVV+aHaBsd3m9eECByOoZQewIpnsr/+5Mt2PZ/e4pOP0S9OwXAOfUZCVPf
3AIhh5USvNg20HByqsX4VszZegOWHxPYqHGGum46Pbk/pEjvCmJ6NIKONV4ndtsv
DNaVBQkmo20K6fK+IuFhKJAlUPEdejV0ELgLha24yhlNYaFcPic3hQAgKgJYvXPI
ccUWrOORVxdBrXCiG83UmQHrJ2Ad1PxIkI2NG6BiYCuDNxZ3aOmXv4pRKb3DDPCJ
Vn1NAVhRXybaY8gjDt8eExo55mq+eVmWeupIvarPtoqg/YHRpGeCqbe/pgMGB5xm
9aDFViB1e9Kxrmpk74c8ks8W2EA8PXIYkkSnd3/pmL/rSvlXv6qB6fCpxd3I7tPI
xfgT/csirSCcl3bwVoq5R9LZUo28e66leaEhmVURlGmW7MWGYwNKJYybzuy77hsX
yjY9RiyujWQAbdk7v33URVFc9wydQJPilTIAceDFrxsQ4JIaAO+HI4lczCwvF9zo
FBP6klX9ycEcxGm80fpQLlsS3qAk9rRzB5Q0v99e5O7t6ZeTDsc1zjw69nRakFTu
U2B+eMaApoK9mwhiGaC1v6/DbIcek7T3BPmUgXSdNT9fkhmXMGp1JDdZDlRCCRNo
A7231icbYAVXW35xV8SystdRUqo2yG3yQnvmdMi8p3T4I6s8d4IJNw57yGR1G1N9
gX/CMpmMlACPS59yFqs9hAf9TPjv1sRQM0QFcJN2vKzQ/CKAygPLzVX6oHQKp4Ig
v4r1Odc+Vx4B6zKe/xAfggwEo20htm3+qa56acUpYuNogoswqLXe2tX9+WNYdNGZ
2UKYwwZ3Hn+otGTK9mGEhyArRfsJ3SU8DS0sezZojkrg3JHca1QuWKMhIJ95Yg5v
4J17SDrxId4s8UVqXN5gIFb9pojyJ+/Jmyzp62/kOHmAHUtUHNdtl39aabben6sT
tcFE2KOrJ5Q+3dw2xANfoeL6bVh3+z8g1hU+fv+6a9I/S9pav6y5thaI+WZVemcz
QEE6Dszx0pp6UjQ96Em+Tixk6wTPSpfcZWitE0PHT0YsD1XFIbQfOh8ySB/T8lm9
AUsczZyeicSWu++M89/INGsKsg89934bS8sdzFpfqlHk7sjoPzyYfTAWe25Fd4di
Z0oEpMg94RfD6QTpnoOzCBsEF0v3JHkOq6/hFvZaF8DE2q3KfgG/AAlPyLRkSpQl
1gSlgB/Olyx1CyiRaCpVLUa+KmG7LQ33CFDAtDP9w8yQBa0ghCXmQ9TKUiuP818A
mMijvhGvPsp7sGcVgHH5prho7Ze69mDorOMYbHneHRZ8/SXnw1zzvwo+LEseGAqq
bm/R68bS3uumU9yfJPW2MMvs/9MN3BM1Y4cUhK9rbksILzoYp3tHnQKboGG1i3Qh
mSQzV5LPB7HxlJQEGfRKk4+jLoh08S1O1FzqGQLyvW2QskIdWO9u/lvQAovVXElX
OZuuSXL65VAgtsmMSPg7M6a/ZVCvc70FQlnq8FJ4kKstptyBJ24AnnpseGBzA0Hg
C8MxiIiaCEmuJnDHOriaIlg+w7HW7J+Q+zfKvT6canZ0S/fAhrB4QGpfAHO13E3C
m7yFfXcdrERx73NYNc0BiMbETfrDC32wtSyhiQS8X7WOU+vjP4SVBsKM8XE0DIpg
Pmhnq3ZFgCf4ycI0VqTVW0PCuIwFvY9WrrAF/oWf1pzuDl5kDSz4d3wRMDmT+3kp
KLPQudses7Lpd5tKfwaYeqV6WIp8HQd2sFxJyLYt2IC2KUiq3qlUYb+ZNbEHSa2y
WvgxIGj56Vf7LjD3D7ONBqdI215pzbd+lcbYe/c7QU4UJx47kUzzPgj2ixtMlzFo
/B8+Vkbk39lGlEmsP383Mjs4wqH2dfjOS0pzKQHs9G9giEmQtzBxiDSp1R7DIok0
tw2JGhsRZLsADBfQleiGhpt0GCgA7J1RfQQoMtdN1GzLJomY8N0VSDUd7C4QEJ7L
Vwb7IdPOh4L0K2WWCCd0UHDEYIYL2POuef/7iUgtix8oQ+MJCkrOQQrs2xBxqWhf
y0JgAADUgoayBGHOZ/EoukLRk+Q1sGJzzU6ZM2woS8XBL8JQHu73+iYzj2qYQKzG
9spvDSmudlYV4jPnItObG0Wfbi0BDbbKfKc94wEBUx6lVl1Pf7Mlk1+ybLqFHPjU
ZQ+lz4GOUgO4QRwSf/v+470DKGLGSHOk6Tu7ddgInej71Zp+hrs2Nn9LhlTuTfob
k7M+ALJ2LVpGgIP+NnV0Ij8RthgU1rp/IJ3wFT+os6+mSQzpEiWu2Uu17BQ21yA/
2LdGtdUbiXbuzDQmOoX2XS3fU0NzBAABahXSaToTvAqdjn+sCICu8a+l2KR8qG7k
3I7+57YYASXT1KiMn1ElaG03bKpmWKNHEQjKhV+EE5aIlv/tl6LAFo3685Jvnzbo
Tf8HqI62GNMxAXTpBbtxjDq1Il3/JJBTDRR3BhWHNqpIlOqfRAkNybsNlVITUoaM
w2ODsmUbMfleR/9edQkgdQAjinQ9dpjPhUx+OucDFuHrITDqeT0s5teepFIT84op
xl7GkY7B74x1GIsrO5IE9T3JxLWkrDS5zEvk3p7kPpXS6Q7L0k2hXfh/SrjIdVRF
0Ud0FddD2ugBUCbVxbidrJQsAd4Th+At8nhObfhh0rNcoc47rhABmeMXoz2oN+21
hyLVPZsEVyFRbGmt3qgAOuWIDUfeYjzJHj9+1lMgV33j4Bk+rQq/1uDQ34L+bHnR
XFnDUuWD+SSujCngLueBDXRyumehxyq5+mctTtNCTYgeA7f2ecLd507/Zgz249mB
C0pBvfQIto/8raji0UO0X47xFzkgQP2IzDnRXgUNdx8tX4WL3BgrrQVZtbqBTO2K
ZztZ7aBpDnE74RCTGHvNEgJnZiyIGvFgqXl/F/U20GE6kusDl/z5XQhs4DLv8WDF
NZFaEX6MEseVDhQVVHIGYi+B7JWoDhoU9Y7ZTOEINIccJl1mz0punUi2K0nCVrQL
s4lrXTO9kKu5IjWBz51o2dfppHI4emn0eqpgAMrkZcCHc2XG9va/iQ0FO1xBiZfC
x96NcRdSAMRI+HuNN+GzthL0W58cAauffxZMdl4k0AMz65VoButggBy/bCru2AeC
U6Jz3Id7hWqU2xMKaRgEFh+slpdGQb9Z0OcTTFNOhatAvw9+9lg4RjFdGxRvyfbl
oc49cC5CSwdf+2WSD/CsHueKvcKxwTRRlP4YkJLgwVdUPkgZlGdBLIqjxzpoyUqZ
rChsLFrTXA6dLxCK07AbY5GSsR0RXrNqC0UT9wNbZxTvnU6UbZvYCZmPdfjElZL4
Wb6jgsxPDBxJJp0DNgGlTR0ymx8DVreVQKORCE6a//0/JCtGkm7p9quKG9AvbxH5
rA/oLC7b0+zUGlQKQ8UtcEriB3LcKaj4ZtK/ATLxvMYO0Vsrpe4PE7pHaA9DYnFN
oZ441xfPUqd2zTJWNBBohiUAzUPgTDeQSjB26v3Tcy220NKaivkIFK9c4IK3Nslt
n6wfPTimF1peGtHVIOlEZAxSNgwpWMCMyB5WUsNqJ2ysGhxXj2DHv+s8WAxdmrkf
4idzLiy3wrJPVc09510xaAMmtWADwlaPDNbiZcOGdmdp+onhUt6CeOapSZgWt90y
24M4AvvfYElEuD9en/pZcS+nls097bM1ifVKgbAR6T8puxBBXXu61uKfNpTngm6I
HHtdoVrwIYDQyzJLlQnTEIKhAKfZ5O23fr0OrEOg75yN4T3GN8hVtxIqeo/sELrE
eDBWXOFMe/l+NoGWp7U06RlEe4osKiJ0jo7Ic6Fj8Wg++X/GZyq+Ez5q+Q+800WS
+Uunu0U9tS+qSKngVsJlIhHnJiUq/7dGDhv2GTDM0wHi3S+lNHlZiKgWoN8ZTEwd
/ezu6Z7NVGeCOwzziJ5zCA49XvUY0gujpp9fBpZzK2CqA2UmFTdWV2b98fTl8SeM
GQiKUeAFyrsIxh5SUcr5ZDviFfx71gn+MUUTUTSkOtSWZYyTB0d/VXi2052KFPUc
F/5Oir54GoB3+qJUyYknX01IHdinXku+A34P9w00CucbVVZCs17ij0rPvEidEZEv
+GRZnfBA4PygN/7YAlySbwqFM3v20tyQysUVMObsPWYIcnuyR10seE9I/Ol6u9j5
O7vb3jGRXVpvaeqJI0yShqJ+rmsBqgIZmjToIzvpk5H2aOPZAk/hyIQZfChBbGNF
65gddejMMImHAfhUil+UIYXggTlmM9sdP7BNb/lrRjo+c8iKxcl80vEcZCELf0sm
TUdsSyA7uTYqIi9UAmPdoABzlLgNu8TeO3LOQDHVdZ9KFwgXPXU79sfJWv5NIkL1
XT8ODX+rCqWXz7T4OlGsxp9fMu6qmFLljTto800hvSlXARhEiJnFhYdJBWvXfKXI
TuC+K+SlskeKAs2wRIwuQo3f3yBvDDPIz1pY8j6COXdHzjEYhG/C/CpVrkGAtW+c
rqF3VIWpwNl3I9EQftZsGc6sabH/DM28+c0ShD3CXOurqv8NDGc6JDNCXA77xsmE
YiOw71FpG4uNOE8P9I4V32Tr/WTZvS6YKO+WiOpIWWxStvbxF+4CNcO5p4fuwgEk
bhcekcxHa8cpMG59l2Zyn44QGuXZOvq7mVQLQGqZ/L7p+rnyk79+8rQJP2pCIGQJ
3y1p2jnzhS233mR/NYskaR9RKaE01uS7spkHAxw8p+i5obGynGaXiZlhB1fadh7P
z/Cc/bWZfYe89ZyfzOr7IeGuofpoBOAFUUjroSp6UBM+16DUVNJTz2DO+yJFfzjt
Bu10MtJP4zngObg611Qr7A2+tXxWnMZhMo2un9fsr57rMmOPZBBhra/l+CyxwiSW
ZA4qmWyrf71nTODGvApQCmm7+pyS2UpJAg4aquEzUYRHLKNLhcvZpjv4cthUmk3i
jY4p9QPQHKO/F59UM5uMkPuBJh9Axcf2UGIGTIxtz+O2ifzDT/4/v9UwQO/b7MU+
jeJbpC5FXM68HbNAIfa0E71YT4olH0/R+fG6b6hvij2qoGg5RMyvL4ukE8EPZePY
N39B0O1sQZjEtLL18tlhjMoxqOmvssoUDSbnHvDYVuIGVEQMRRlg0bWMHb1HSezj
dm8MgQ4nuJQpxr5PDc02klWY0aoYYXPsKox3K7AkPnnc51BWt7T7PhtKtx1FOpJ6
B5fmTNcq1XUaYBVV+kzPfYFEAn/4mMOPjA5oMw9fMvHVJYU4I3+0GujHXljLBSu3
bayAAfCOtF8HjhZK65JfTpav5HL+OZ44pCa/2h6NZGf1CgJ/OyvBX4VAPt4YDbcE
hYbYaM0Ey02fLXoS+k0vjT8w3643tKgNxQ7RNw02vIc9OywFzkKj+uCeJlyT030N
WmCb9v4Vq4miC+OdSoqjbFVK2dlYDKQ78w0upH+ZCshsJm+7LNNwpjaJ/tl7QwyE
jkpHBpiXYpKvjSDgNRyQhtqw/D/ZVjnEfHm0f04zfI61P1U8I5Hxl/i7f2C6s4R2
ABBUpQIkK1HyRjIWMg4HT6i2Jn9yBW+1sg5JrarkX6ARyNxKC1VKlHbAwoV31CkG
6AX/iSHHFKWYQR+5A3dQEhzMKFx/ztrCLe7pCYETAHSTEv3dS/CjvQx4nWHbYwnJ
sJd5jAhJTqL/W5vCb+xRrsd9xMnIZnCmXHdcLi1emLPXPAlTZs1w9Wcy8bfWbTuc
+Ciw0EXAb2zBCD/knpCWWOQg0CtL+2dgYCd4M17eg9v0p8nwcn5qe/bV6rVBRwEe
jP8/kqs7RJ/zVmjjUy4QulzPfE3yCXqauSbowPNoUHlQNPXTbP1opCorOlSv1fhB
gA0EEDnvwIvF04gG/i+eSOrRR0Civ2VbNiYl3tUOvOziZRL/M0H+hV5ASokGlUJC
DC15X//GwlU5JRWENRfKVBtid19n1wpfcVtk/f0ZsTZFDfT0Cjatbv9kTs0UsP2f
/lX/62XBsIW7ksWBd9LQubRxfuUze3wA4zxbSDnzmC0Y4sZjpEn5CKOqj8yuEO9D
kGSdzoo+EkvGP8zoeo3rVelfSOl+YhYDokRbkJxU7E4iSzF3wVX0ryd69AwSk86b
576Re9/DCTMXpVeQZwpASR8Pq9ouBSbOg4xLidX4em0KkgIzhQcxD8PFMdlwdSga
qECfYCoGhJpqG7TVWdeRqXyyRtNi1/1dnrihR/hkvUDh5NjGdvfjTMaqKTHaHFFO
1NoXkcMzw6L+GjpilHb5FUODcQ+zp2MCY5bA+kBDS2PaVhGed2CfVKw7989x0CQE
zYT4xnsZzfBCibDRnYIWr+LCJWwfV6NsKi4fQE11v0nagbDZ4dk9xYFRiuuXXscr
ZPcnPDzSw/7n35SBgXYpneq2IX4+EAoq2XUghRXe5FcMoKKilZwjx8DIRHp1weNq
3MOSaanCoBLD/RjMgOQ17KfuBq6mPqQwTkkShpEWTzMPCvOGLNr+7ybYqc0zDZab
YDIASQCAy5BtSd8QCsZMROy9u/EZn+aKAg7q5LzRKsiO3uRW6fqav0fZakaaD8Nr
BpELM7IYCKbxDBxut8mvliBs7dziAuM9rmS0LpermWwoE28cPVvLEkFUppKBiVzA
fPZKaxKZI+JW/RKCGxfIYbmFPE0jFZjbfwuB2xTR+NaRphJje3M2sqp7DGrTjg45
aN7zqDpSVD3DCtzB7TkPWQTgAF3A6B/Jcn56/Z47Pqc+PRUU6l5UIp6vh5TibZHZ
JCQ2G62Qns81QNF+Rxos1l/9T9K6S8XD12qWO36jJKUTcsGReM+tgTnjSBy2ulEd
mxyvkyxyaF/YYXglGZlPQMpJBnA4sFWOqn7XdvGsvWH+jZGPxKmeDHACul07/eU7
AjU++VYuhYuZI0fyNQ4JOCZih5QThzlIKthr74JpZcZWwVbSHoEWhRTZnwYQ6qi1
sD659x4yDzIpZvr/q96Sl7IQRHo9OB1HGhjJ4cCW/zxOetYPrR5yPP1cW6VO5dz5
t5u+sDJkf5Jf4ubxt36t8BSrawvX6ShaGIpY99R2nG2spS9OJQWwORG8ZrOt2Nir
tc5DN6RPrSDB0AGwbbiTi9h/BZH+q/5pPSqyej3BZ0japsGcY4rNIQVis4Cvwddf
CGMtuGl+VoRMZ774yZou6OoNspfm3UnvhaK1rY6et2yRbX/JEJS7z6D3oLhnxiUC
j9Dm9tib/sr9BWiXf10lMUylRjih2a/uABTVV72q35u7khD0i2stlwP5BOJn01zg
EoARHU+IV8LsezwvGg0Nl0M8lpnJJNd2TWopOB0045xn1FYI+CJC6CiqI1l2iia5
t92cKJZk2aa2onKX4K5BOjdUQQ4F6n+EgFJi+kDn7iWAzlnwP4Ee/FSgWm4S72Ft
IpjHpb5JzbPp9pZCiDW1igzDVkJxpjZZbB/X3UIr5AlOA8y9hPvhZpjCfZ7+SNId
u9zIRQ2jSuWZtLQAfxqtJIHeEuyjAF2/UdRYZQXJUmOnfB5+0xypt8tItRqVZB/F
YesvyFR1z6guMMf+PrlXuUFb7o2nbFb8RWH130hDqONd993qCk5H2f9yhtrmuUcN
eNVkOJmkPQkqLlugbWEpvWn2WnCbj/+j8pssBDUBRwjxBq/kpwO81xaOf/59QEb5
DAUsSEdTKnz6vtdyeFhs2UVifWCkuRqmUgHig+72IT2l79LoxViLbduX2F0DrGV3
soMjVgxx6uSNwfuWYePjH/XTKjLEx3whtyBRQhZyzEXeD91Erc4VYQWgKWFBLbAS
Pj7i5I3F3OuD+2QUBtbTU3HQpRXLXOAj7RSVZ/GJ8GR1d1odD4kG+iW4vAj0FBsb
lRDCO0/eXNPrU8Eu6bhyStqgwri0TLOvQKsCVrA28fDC6Rr7uyD1rITs+qpldack
lxijE+5bqgaT6E0uI2GVsbP3WIiUZdAiTcZMeWrCxu82bI1aEGnk6i3aLQh5iQRU
t4Hnu/61BinzFjoLaV0P7ENjq2hh7BL2zXX05ViDOhaTs2UvnTQi3djL9wdzTWrh
cwsNEdJZbbr64MgazZy+OFTb8qE+Y/wsE3SP0yitqoyq9RaafaNEMkJG14ravt/B
su4BXt83DgWIb3w0Sz58+7q+Yejz/eVATM96JFfz6rsD7cUZgbayB/+asixnXCHE
5IqV2XwVkzQsqTOE8dPhq/Gn5f9Sp977PWjeEnySp5mAjK2OivFi3uoVp6QmXosg
PonUJzAZwg3SyxEVeInh2XmE8D7vurNMNLESmHbowmQH6OoE/RnViA5PMYzwL/wl
uWtPs4u5nRkC1EN+tXE7d7QNSuS5Q2oz/hw56JDkzdHMI3BZvXYanblemFlehqTE
AgUQJVX7zqjaLalm3JOFPV3aU40mFuKKPvo6XLZzZ8pDP5An89wLKsG9NhtUp359
aboI4YxAMCPWmyNWFtyI1UKG5FuEMMruVX1rOvnqEhICGW+5Va5FkiF/ml1nRZol
jT1dcd64G4IA6qfXt/fDwffggNrGc+XDJGS15t/v6TnySQfQgVnFkpMpKzVWFmz6
lhU5Czz8g4C14ko878tTRoDmVVj4Xx0Jo2ZLUNw/U1a5m0tmDvEtuKofAKsjTY06
YxXb6xXV5VBNusElkojaZXqFt+WHHw76t9bJEo2Y3SJK6UyqjAIsNI+A4GRABm/P
tTCzrYd5Ba/LRK8NJTLAWOolYWAa+Li8YqVMP22nBQzeZShroi5d/gjLaAb5zLy9
oFjHTmpIgr2sSIM3dKBwBA/iUduM8j747xaHdmrM+PME37JwW18M6NNDfAAulrIz
LUrujRlM3y8++JCVGb43WG/9QhIwn0fDEp8MoxchJyqgztPh+8Su7vPuJe9jzzEO
e1YEmanZIVseA5BsnpZghHAqjUdmFvJ1bOo8D+HIKoz0Y0nxwsFIKiL2jjlA8PQh
DV+0lnSES9QuxZNPcyIU5z/z+CCcVsSWJSJlbxYCyDmTXU4PwWUN6uZO59nmLIfc
a8Z79LF3EMUcH6y1POMhcqzTG2wzJkdYQf3BEfqz9iDfwx+y2wmzIA3q0qP5K7vN
APdgwRA7Zt+SL5k8L0k0rgTgVU0Qnsb+y0mhYbxFohZX/c1LuDgYfeNAzhlLQJNF
mRqbrlOQ8pgC+N2VUrBuq2qkP0q0A92DTQw5TNUBN6JvX89ZFLzFsRixW3NyjdA4
ptE14gTgqT78PSkFTVscCaExJ5uFqsfWtKb6M2k4Y6P/X6i5fC8dlElmbpyCjoDL
tWnwNMPEqehEDkKNyx6AUK5XXEt1xmlhPzEkShfzR+WN6sAtbjo4UbHYYXFFbApu
pWmVNxYq9UUuP/bwT5Jn6dArN0+R0vEhuVjQrDCTMs5J1rTbknMQ/8C+U0MpHpjX
0max20/Z3DS684sDrgqpUJ0rWhfgNEnXetpRw4DjLKXW6BuWgCf8iELdNcwYbCgU
7y2pg2jItyBilN4MJnWpNuNclnhowuabN+cOjGFhUEgqKUyDfgLC6idp8zyHtxXH
3nevYetj7wo+qORroTo5rqjTS2IKPn8BTE8PR++rOoN+qwqILU4ZJ5Rg8nZREI4q
QCOzwl1u4mziVk+eCrUlkg3hNfH2QX3mv/BgUNBkyNeHZfjzuiLBSG1b6AonOsL6
SRdRU5y3+4CziiuxdRsE+k7CtWEAx8XQOzaymkP1BrnmNSNg+MxhdfDHcSvElC8a
ql5/pHZaJ3ELiUZLLD8b1tESGiY4ZNQG4fqXS3/jCxrHrz20JB1rYSENiP2fEcp3
7fXFYZpM/a+f25JDvcTinWZvSTEsEcmQhVpXSbOip2d5AK7Em0s8837XWV31ZAWz
shukjMXWXGNK1aHPr3hTnT/G5Igu914wFF+OUpycJswIwKeSSVKB4kv4wSZGvYC1
TIfAupw5iX0M0DvelKFwkIeaWLG3pxrmgrhPBFwuXDmMa8I+uc9KJQbsJbd7aFJE
dErfT/BT5g8ap64oTefwOfCLhJV8M9Gy9ypkin7d1aHmk0DqBjTJoXSef/Q2iQhq
zmRtvk4NdXjZxc9Er7PGU6tCf55sITLVLMefBiT/ZcvrHELAv1TYstWYJARIMDqI
CBwDy5aZqQTlJEiJ30e3uU0LaJjufRMk/WAcH4HyFM+bJwSUrKH7FQsbNKO6n5Gu
9sDx7BccjVE2YXqL+4FwbHOb/a38u6aVsVc8nYw4wENcYyWlihaGQ8yY1A8qNtZH
31dqXCIy66SkvT7AAh+bX7VvigYDSbihzMRN1pWTxNoZXoA/Vx7ldptK4qSxcSOQ
acuwoETo+vls0Jw9t03iymdkXJ4PeftWMfHH7nbYnCUN2joQlwLYrEMomg0dpaFA
CN1ddBFD8UBnaaaxsBBIDTteki7MjQggkiqXndJE8IXNJJtYjvATcrFMwi4NVMT9
7IVWpbTg1m30uQZzzkHg9O96XiQa27wUiSJ8qo2tKm1g9T9h/Oya2+pTypdBJbCb
AdWR0IeiEV+0UWQRI25gGLjBTerHU+B1ltNh0hHsYiLJckQjmRt1jZE//JFsjSjI
d6hqDAUAjGfBg8H1fvf/V2MJDGjNR+SPt8KWPK1ApM0yME0PCpjDEybOe9P4tehe
f7X9JYqP9lyA5XRukwO0IkNf8qASZAQyvCpz2a3EbLkmgKknSv9v1TVxBF26uLnt
yJe+/TuyjtPsTiST+GITTg3PAIJauKTyH3by4CldzUVOD2VDR4hJm4iVQQBzudRH
YpJZBLnGQKVrajH1kKFe3ktjTW2Q2idbs7m4kvVfaoKoWO1D4Uh/B3CDCHrk1Czt
iVzqTUyLSX9TCx3VIqMQhqL25iP05YHCB0dkG1mtnoud61OoSkIY9mEnIRtfP2pc
eKwZXTuTydu3w3OBUKP9I+y9L+PFDqfE7/yocmNBrleGGFdLv8z0MJbr9pvXoyYj
SM+b7pJ6ysoPvutebGMw6Gz5DS86RhNai1f2dh0oomo4bo+zEJo5zfoil+u71nXs
UtddLvuwW/r92o18iG2Jcb6InJVQbsFj7bW7WyUfniEIWlKKsnYzDliltzHHQ9PX
Jil2+lEYAYyGUFSQH6psjEf8uHgD+Oa7kAojfURoweJst75MBBXRlZ1VaOy5jpVu
BQqwjTC7aZQjumJQhg+JJQE2lwEs2ZhJf2IQRqDqdAdxd2erISViEpF814JjunzZ
4u5u13ovvoYzsIov3lHX8G6ca0+UOZfLhY5p20UxsZ+4l/4LEcanKrVEYjTbjm4s
qVsDVSov2hACGLMrTajA4FZehmVet3xtPPCyh/Xb54pJmJxSL1nfzPP8p8l1+d9v
GQZFGeCdrpYHSN1dzxw2AjPwJ+F842WbxJSj0FS1BwSowlG25l9OF+japPpX0oqm
5BNIDqbnMO5ZpcuhIN+MntHrJTHKXPfvkugm3+TSmwN0Mzi/QXlqRFix92mZMzwx
H5/ZwhoP39c760E9duedTS8xWFGCXl0gnM/WoVBPQC8ox/XisEtoAOjOlBuTdl+I
lXjMRLK4EzVsxtXq7TvOpAPl9YL4FyHFsqgdLIJckKp/Rp7nRZbwbjG/4wbShejY
hW5usDcYmVit+mmBFjU47kJ+W54LHfwDu8ddyL8qB7NQLzB8oZQrqjGYM6ZjQnDl
z5Vquiupn4iVe9qESeEX6EEM5+TgId9A1t7TZmq6jp4b96/uu8sgGWd9F1HN7uDC
a7LR7V1Rk+HMFqhNDa1xvqZgeEEWUWZAkZvUMgIWFh3u00723f4/8zPMc1gSjCz6
CtNcdmyEFaMfb+ZEO3Xy9n5T3taYvHw5t/KXjmIrJnDLybhSwiFn1pXavDvAXY3u
8NlUmNXfLZz9qO7WCmysO9ad0YQlNBEvTkDcNAV32uwn4gB12feeLoXBNRbbQIA9
ncJYf7693mZNUlO9ZPAhoNiGuBIuTF6IM/YJ9fbo9h1eDj83y0EOxWhsewSk5QIe
MpjTl5R4cJOEGd69VpChF9WSbHRNk0jvSGAkibgyS77fFD9S2JXPSx4OzicX9OQ3
KiDTS8qjLUFDrkGiPJlKN+jeVeoIHK2JDTeVx1tpbgpIGyDFevf/xScYRVCZWQ8A
x8hlLngVq4PQpPmVhzpvZA3CagaLby1pWabkmONAn7efUVBMC2U/IfmYJ5T+XkYL
HImRiehJ2b2nUFUZPnMkSHMLN64pF8y3LMRNYCj1Dhl3b96z6UE95j3uMTkUSRsA
uqPOO3Kfl2iWiZH74K0948L50jGyQqxFjGIxldKJU5cWYDktpzQVLBllIOP9/31T
pfBmqIfcoMWvyD7OBoGauECN2OhIl0bhk5NNQhrlET33SVmr9RXRZVtvOrGyzbIt
6bT7NNnv6L2/ElCD6VsiUkpuSsondBZNjBlRdAjhM/ibdxyxm8Iw/HqbyXEAPfWX
SN0yJ+RAsuYmWIUT0vWAAvSgvTUlLic1zKQTDhu7BRDeW0AXn3SExUoaPTBkbsBU
gWO6GVGlL1sThsM4aZPI493sWfK2BHZUJFI62R1ORznay3q2nXl2/FibPoRAvuOb
+kcRZ4XvtAOwWuNxDhakyfxcFC7faVMj1+IS2+2F0pBVxHj4CL2d1UVqMQ6qd66l
XOGZp5gkT3o79LpvwvGbo3SAwoJmR6zZ0aryOzAFpF5ZpRq4rIESILFhGikX1hmd
6mcm+2a1Iqce/zzbuoboiltPKvZLeW3n4nlrevEteiXuHnDzoeaRRBpvcJXa5HpX
69Zr0pKXjxkoyFet3lLvWXsZ0sVgmJb0Go0UjDDht+yPYnwRcWCISCCJBfQZvacA
bvl+0fpCAzdRkmElNrQFLLSThHcQGw9t7to2uxAnOcyy1SWR6S6TnGo2jowp8Eu8
gxvPzi0BJecJ7gkkBxd9oWy3EY5wGgRsHtuUz1SrUS2CZCvCimRCfAztfC4Bj622
Bu1rji5g81UtbTYIZ9LZpdIWbP3TrAWz198w2FIxxCWwS1NKhnZ3M+ZdvhRi3ZQE
PYz+ID/hjbDGSXpAoQZkeC7T8dUJiP/GeL/wpatm2U3FEgzl/r2wVRdAYhckvnT+
HDNuaJTpK6TBYaRGnAcY4ZcgrcKbKOLt8+XSHHrYoIDagUvmhveaGLLv4YcTBtlA
DK0j72/QqlaBCExWNTJkxLW3KLpkstj2F4qH1K74EeMGodbtjw36eradKqxTN0i4
ITn1GKTfR9ZBmz3RXQYp9lb+qMMUU3YCQaJbhfPIt9gV0LmYKxGS6c6198HJnFNJ
Zm2nPyVUPH4d/b+DMLSUpK0wIlKy1uQnbgzCUleviI42zhrmCRdgHDkZHxTLjRjo
nOAlgc9x+1Kn5S7Uaafp0NPhre77RggcW6tWZuadDV6XE5LVrVBPYzTCpxe/r0mF
FZ+XV9GLyI+iIlYJV01UfrUBXLquxSINh33HlZ+qz8wLD4YBxnc17sD/GUfzXKCQ
74icsOTjmFA/5r2kzjsVRzA/RkM9Cb5jscWWbL+TVn7W7LebOWzk8+1PG7gL9eV3
9nTOwFweyIAfoToJBDw3bNPGpGGei8i6eUfc6vFZEYc0VGKfNMv3HAbICxA3tjMO
BMqeJ/7GEe5ndNx/aGzUBK7rOno/xUWhAnE6E5GqfcJ6F5lBoEX1T7SfwtuYB+ea
vPo9rxuwYLRA2+Gs8hMn4116pHOKCy0AxFst41t3JmdbZ21TG5DYTnz5Ya3YBmMo
OSVe5P27MDwbXUo1spTRGQ/2lcP+demNuUZl88jdY/iJaye+9wMjaaryFIC+DJ0r
Tak6/LkplsGUUf4ZAlboQ6Wb35jPfL2yC3f9/7vbHjZd7wFKMkMZRYqq49eiRoHx
ydqy3HqdT04ZAFAvI6r6qiJSSCfXivcOrFxYMgdnPd9Sbz5T2rzGVviL2WHwxPEA
fZnDv0bbewsqsolG8dA0rRUjLB/SVInJWGn+1V5/aasoCI0ycyMlwjtYWIwRdfUw
0RxrRK1Qcd3akTS4Bvq6Tq2IgIze+5e+n8bLz0Q+afCkTV4CEyJb236ZVW0YeKE4
uwUKbqZJ369GWqHL0lLra5kqBjbu3nzRGQNUG4LdGS/a/MqylD7QH6po8LSPsETr
5t1/sZ20G18jTD5BqC+ZHF45tqwGfQZOR0IMCjt41wURHd+SBW5Ti88nJig7yDlh
HfurBgljZFhNJwhi1eLeJXmTP9FGwqmh0fvfUmonY8wjsYUhvyNW9Bz8cP8tb7ZA
132jMhN6A7WP30E1AZSVzM5HgVaA0lbQC63BuooWhHUUC8U5YF7MOZELBiJSSpow
6xAJq4M69PNg/WaI9XfhNX0aPOuP/hBzCHWcTyFA/ka/qFvhsQiOXGrtcWnNW86P
pR9Df3esDimZmCjIiQfOKNovBvCrdql5EfI/KQq9EjmHTuyBNn+kRXBxUSFQHKLc
qkZzI2hCkGjB7hcuiZ58umk8osDGA2x+MDoCkULeaOLHRCd79aben/MqTRvAgSs4
VpwuxUBjddkKt1BGDR7bVPKr7ts9AQN6RBHRRos/6FlDTZfM6fmD6Rpzi9df5Nh0
09t5Sfwh7v5P8zC5TrxjIm/he+/oQFs6vSvTycItbSFVYljBOxnxvJA2kGi0JHQu
DV9GtOiwlOjolgSVs+3xmvK7po6aRZ9lO62aGmb+Nj+41NrR3pJpEraXdEZCscqd
5FLcR86g1grmBGWPbj4Y7bq9HYN6C7nQJ69kywpzhAe3xeVJl78hsA4tRaJOujXw
r0d/pjeOk+1KLO2c8bgrCSMfkQc5PUdm21dyPSqpcIpY3dF+n01Vr7YD9OmypANO
ltYI3qMZJsHloSx7ah/nkSLToutZgmfdAPj/rI8rafQNVUgQTLr9YFPJWc5uiVo6
VA8OwNOV+BMBJXvMh5a3HlZj4NDgDjhfx639mHTsex+ItbSBlHQ3hN2QzLKpLjtC
n9hWaudcVRClSMcEn7ZspaArHe0o8E75DucCJ6XaSeThIs7wJNm9+ZMogLN8Fc6u
QpRd7l9+xzkt7QUF+t4Mu3byi29kMQcgt96CXRMsxK+zJA6+DQKcz7J9S3a0jSbg
7DDi0UE7T+Ku7mq2Qlqcou3NC5qv0c2rmm4J2Qy579A/7KfJuilWSrKZ/mEsIHDZ
P0zn4RkPpChN8vgFEdF4hnExRVGJb37Q/x/n8yKNwHCtdLYrAweae7rM516elNs0
35LgEe6HuwNBegrCU5yx71YTwcsbrM8/NcRJ51gbqzR9x9kSKiXBBREeoG5mfDx4
su6ybiP+rApF9OqDA+fyjKQqIWjEy1MuGfxByH6U/ep54LCzJBtOQurHtbZKZMq9
ta+yJ3oioDhP6Y/lzTEg8R1IEvi3WGkdBHdm08Lq9WcJZLLYEqzRtzAKFDpLBA1W
MUhtDjwCtZ017dfylZCay2X532AbU4GaX5begfMTZs88qdsuqz5nkL1cXAHr2+Hs
oTyuv3LpxXFDh5ddE+dTAPiaA7XuRkjZd0HVxWK9WWagI3CR9LH8P+XgopkxaxWv
y+uLMm1ys6yuG1Lts4hipmt0a/fHJD7cei8w+ZZZUMTPV8fjkRXIsESCsGg5T5SO
AYQNVfHVT0X2hvr/7TAMyqYvNosVIOLy5jkoI1G39zp70BMW+zHoeQjUXlkVNSN0
sn4v8gYO6nCp0TrKOWoNCh/s27TOvz7y6MmTyKCLp/GvIRPshrb/o38v/GR4BGz8
hvHZw/QxBXQDXlp3gFwav+lEgtGd7n+zfV/Bj1EAgSk09mHbDchWVNlAVR+b80n0
Ko4rQibTF5WIAAcMFo3mljTphIfd3ohifctmT221tWaO4eRk1l2NjBwtxZOA187F
oyyKKE1GVz37X6Wg7rW0zxY/TKHRi4DBVe/zrtCg4Ro3u7mz1g8sf2JxTsJ8uFgN
HhZfkepiAoMz8/DaMEUAHdD4qulZ0OfaBMpr1riwjy81CAb/7Zt5NVVBf0NwC8Wi
2zb14DMaN1QvCegqAMOOFi/YANS4Z7gWoiiEZ1uiVgob+adKAa5PuBpe2TZVRGUs
eHjKwz+gpTAR8gn71xp5lLf0QeyGLZV02E1SPq4TC1+axaRYDwOhZ/OdjHrFD9pn
6tciBdz58SseCEP7zaSbbui6tncMODJF0F3cykNmgp3/UbCwc8dK42nL2NWOM3MI
m6+2gsD1spSn2MN7Ojj8khf0hVRFsLx++nSIptdjv5e8Dta9DbPa4LWrveincoLs
PNKUCcL4CwwJQOwiCC/WJJ3AF9j+d4meW9F8EVglQPpQzznYfJ9bHRxyCg7cDw6W
gr2J0sZzdy/yVxd8/4UOMsjXxxvNLAXzzfQ9Vi3qAl0aUrF33oNql20dYzMPDr1R
l1G/WDb2RONuoZqZP7a9raEgKGdBdKpXcHagWHcHGtiAChwp5pLzTLoI7b9bsot+
ZZWnfXVltKH/sCmtTVZraifAz0JXazE0JrsyzVDWZwCm0/T5o665xydz77QuaYh3
q9D3rK7aFAX6x4ITcHcdqlHvg+5UtP777MeEfFX8EU8KBqIJgBk/IaS6fe5kzQPd
5+sqi+Cq6LBBUfYvMuFMklNvfScnl01zgeeKjBFoVC+sMqZeD8uldvVj/IQyNrxV
uuKjSfyxw0eNGRbTZXZN5TtH852KxbmncuE6Gl8KuQBeqqsAWFBaRHAlSeLBo53u
X6Fsw/9obTsXf/aSfktIyN/WgHx1QQc9cZaH1CRMmUgbT6rZY5bmLr5FNLtZLSmY
lP3qkd2nlXzv0mLpsCROSJMcCy+R/dopFRbgsOCwQxZgUj6Am/JkN/rQy1i3F5tz
1wUkZrecFTRKFH0W/F3vb8hwBEdGS2/HUIlo87rPOkAnaT432h/RNc2vZbnXkf1R
dh5vKQa9G/0ZBknY0ZKqFbDk2bCZzNGwtUCKxchBKkVITGh0V9pjXNqwJNAon8ZB
R0R4yBm4yK7iWJilxnNAAZTdMPDmQRcvwHrtCQsbsT73xE4Tttbuoam4DnhwTGUL
kf9iUX9WOqTjYLfEJkHrKNBFpuOl16bWk6UazeR2dFVkH9ecN00/+2vHOHLNNg2y
M3Dcr/g3xo3d8jmSzGLFEuyqQG0570iUX6PDXIWG7f2viNpchSXRxbr2HNFr+tQ/
pOnRP/gjRtY0+oNRBvmVf7g7fav+03uSVsygYS1kY6Veb8r+EnkJRrOhqu5Na7IC
BGtqBFVngYpeL8dkxv6NNYF/7XE1SprytS4Sgc9dObXmEjBupQ4W2lfBw0i5TIaS
9OYPQL5GDm3MUo7/kabu0B4omsZr4jRTHi0aaK/uqAAUC3Ei/kMw/sOaj+StpnG/
SfPuBkqXIKedJMeHOwTzjxQTuROQ5te+VSkiGUWneBMVTrevlXJzpm2I5Hv3QcxO
0vQZD8Cfn0snrLAfeOkfPY9FaPc9iIFEdjxc96c7LcLSa1U+KGNnOic/psTr7QzP
mIH6YRSEvLslTBA+GSdjRv9f8WwlA14tFT/U3uLILNhZdWJ2zAzQq5qdRU2nm27F
WJhmBo+6OR5BgHfpcVdRCFhAJCMY2SSC52dMLnE0oA27A5nG2zczhz4lfB/tBBQG
MgXaSZ7NEfGh/TtIjj7W9XPDyQpNYhWj9Sh/HrPh6GxhbT0NxQ5Jdlhucvqe+972
Ci/ffd9Fu8A0XhZpz6oqn9P4VWqvR/b4izzHBtHRg8fiIvwrqczRoGATd92Kmo8c
h3QHoneu/pSjZbvZ2c+kUroYBWkNDLCyvjLlo64qHaRJnr63W1LMgh71kIdi9KHj
lRHjmZB70TDSkgU+1/BiGJMqQS/ZpTT27MCkMBpHu9VuT+oWMQ0PfujnLQ0kYzUq
iXGx0IhHyU80k/fmo9/3EjpuJqYPqELvpMFue4fzXBRtXqN0Qujxd2ZYFThzMAT1
4pr54fg0NTcUUK/RVnsWZdZn/gN/WYmgj5rI7LmOsui+AEcdpNdyaLPXB9Hyk9Iz
pBDvEZ0Ua8cFoYtR6LAGcXRNb9ng3ql6H68lXweXv6ls9wwXFwBpLPon5ZkA3fvD
GoDUZ3whHvfX1kyck2Knb6HLGAJIFSQxDGj9LOYBlscMYmN6pS2l6gD0opqHJR2M
fucdzkbPDBv/oOlvY8+ymmqms+nIM+D/eKRx22ofsh6Kexb3jec7ccLHu1lUU1u7
tJD0rManX/a6VQMUO8ftghpBIScXBSps95A5ldTcDb5ddHUR5P53aGcr45jxqV+v
bF4C/qQGHosyB/6QYWPylzC74wVfKGCfSmCBwC3MlmmLvqD1XhUTy8NYWFMzCWsS
uwuSqy+JS+unKcu/1QxRitlcVDCSQbgeLaRRkoZJ/XlRT5BcigK9WlP6NzYArIIt
yWPa9iF5mmMxgLWQ10gNe+8NafvNXyh/YA9wnJiiJiwnECvrOq/Rj4/ffuzWMrgG
1xZmp4WZ9AYWcKTVL1FMtMNyl1q9+AwlfrAUqvnthsQFGYHPyNwtCBAxYKgeNafl
HknP4z3/b1X+1zg5Awiklf3Sp9E0kOrEVnE1LXNdTYa/iq6U0RCqGxsgwtGOp+KK
TQBGQj+w5ejaf6/0Ly1UIdKzs42esbykna8B7JejjiuJV6Reqjj84DuGw10orHZI
V/hX/B30Zet2nixCegtT9ox7VDq5mrjz4pogzHDOsZ23Alqyc7tXb4vtXObqU9xD
cQEDpFPaI38DEofV19CnWgCYLzYe8fhzVJ2r0m26r+637i42j158qfcs/dShB3qy
MeyFWxrTxzljpZoKqgOtwTa6OxaT1OceRKFKlDoBYeAFvgQyvNOc7zyMsnWa3BTD
bsnHqLgyqQptsfGDMpfm6G3sDq46tFt0Cg2DagNHq6Tk5gRMZgAdp5Ei/1av3ePO
iPxP7MZIFPTArFpwzJrYX+xPXHaHhQruhMLcGBShKPEGPzvtP+0H7IjojfUWkgmj
5xaHPiIRrdPfs4NeBMC4wQh18AoID5tm/1rNq1C5taYhyrpWMbJFMz5bsJm3CJ1/
MsXYiGneCpU4ssVbtCse/KjOUTwEzSbhCSTfO5an2XwoZn/Heg1hVh8gWtKCZvIL
KtjMT8zXG95MQ+LGEm012xTbGA2KtAjKgQAA491tGAOG2U/ULxN75XQikb7ISL1j
6nZwaalPfbMAN387R7/gpZnKbRSlerBl7zO/JA0BM/Ytndd2mDyruG1O5HxkAxai
bY2ASAmWiRRjyH5WgZd9u6dw89cVNagO79bhxUo3SZv7y306HQBFKUx8FJ8zNCm1
TWX4eQJWi/BvCqFSBkBhz8+93qGK2dGTnEefeECPlpiFU8wdCJoa35gOfLi1Em+9
rX6ylRjN7Eb7nOakvkqWf+6PzjrwOcE+cqzl3NMT56003WQzYcgi/z2cH3gDvxcH
d4yiC9pY35/nyUpOfDVGAVypp8d996kPVFpSBlQKyy7fqhWEyNwSFDw2nomVgN6m
tvuIHYnq2qACWXzd3DWYMe8knutZ283CppXpa3WwqdKN/JVCVV9lzpk+u54q9l8/
eD5mXnpIZdjS361Wnp9yfd9LFC6Hs7eowIgtrqqqlKOrPT68jIy3MNoD2YLCpXN4
Wj8NbrIt2w9YxSr2nrFFauHhQnyz8n8MeGxHIVL1PMwTTsyAs4OH9RKXTCnYZ8z5
kt6VNaEZO96vZMbdBPOoPWwpzb9Dm21BGxxI6RLcKdyjUmyZlF1GXGZ2AzxyAalB
VCbg0F3zBMyYrSOy5X0X5RRR/i8a0N8RAQ42B4KikO934NrMdisDqnU28Wm+MgcH
LADJpBrb0JlQAlt+3sOXDBNpJZdalLNxmDqVlFHeTIh+QAb3Fo4uaQXHnCL9P0RH
4AIOxAu4g9hn1FHk9u0Zbm33aWNeykZdBdnpQrCzG2mXJT813qdb2SJrupqev+Sq
8oziBxnR0lA2oLw4H/oqy67x3HgP4HUg/bTPtEKNDPwxvUucjPngeeNsvemJbwfc
HaxqTsspTySWf/X1vkLeoqKMB3gK010CDwMRHTiTEWp5maFVahuHokCI/ht0RHXB
ihluVH9xCU9X/yhc8BwDDYjj1AZD5K5FB4ec2wG03nXNilB6RKpfrXgpFDQ4wG9q
WQj7qB0KmUOtCcFKVX6oO1Mrf8GzLL7S/oac3VNgyeNQyX8epRAeMrLOrZSqdwZK
eoKClrJ/OCSQF6LzGksFRm9yhirZyFUOV0YR9xj/PvQNlasZxoRWijDvidc+mNZH
aw7QjmqjrO/1/GM9lOPUtrU/0ZMIhlInY6uaDBAJPQAQLEvzZ3nEN1pueX7udoZo
ruI3heoW0e/Z8zXqfbbvfHDMf4YN5JFNnfUOc0F5kmFgIv8JTbSgY+ur4w9BoZ5E
gEBTRl+53m84fZltx0juWLiv8Xut/cAj3LNjTV/DmpEadWVyksZoy7t3S7uWlpko
G2s40M1vA/PZhFGoNnj/t0Y0T9c/zTINfTic8fbXdZwdZoVX/hphzGA6P7IWK/u6
n/79Uyv/e5RBC+kNeXnfdZQbrAreKgqglfWpGwCfZYxX+pBoyxRkpWnemOAOt0OT
jSMG0ZmJUPNtbp5syWRUn1Ez7X36D088ZD7otSVUqllGAQ+tU7wodGCvqc3Ieknc
fCogUoDZx4eVuJM4bhxcp5cpj5aFrwmERo4cNmR7J5obKam6K41FypaTbe0GXFBa
Qp5FhTaKRsOuIeXKm5Xeahtvzcc3v6ietht9FQ5UaFnaDnbig6Mznhufby88uodk
vPon1ct62v9ZKawsgCIKltdjEuT3DrXiPMka0JTvIN9Sfz1ByxRJgybevIehAr54
jb+/uhVU1Yrpedq3FRDpEYvKgoaIfD7yR3tAfvg4ZUq4Ns3/GzdVOlPGEJNYrrxO
KToJwaF5Z5nOq6d5FhQBiakC8jkNp/E++kofUJlxpJlz3ca60tgCDifHXXtsXBKH
pYL4wwlq2G3cM/u/3FJJ3G0mKVLwE+erpy3AzUuGt9tMH9e2ORR0YW4Z9g42XprG
tRkAVIXo0KhMJQvRWpFD71svut60vKOMqsOz6ZmFH76qPwY2+lXNsB5oGrWYkRpX
uF9lwRBXwx/6TB1rtDyYZNjKwS08agD7g+ZDmZI0Q2eofXqLc/yEUHtmXbgDmsRZ
xDL9YT71oJRr/7Vxk1P6ZahPUKMsTM2QHmH26CuQgM6vjGzPFeaAAeNczpQTdJGq
fFAip5FRSSf5kbbL35fyWAGBLiEpFUk+ATN2+NHENpaMIig3UnQh1BZXvOr9fqV+
4Ckio/YV6Ljr4nWwRowESr/RsxHENnbPREkCfa5GahhRNlPpuhTqTcHvQG3vLGZK
7g+vRoofIVlnUyJ2p/gK0vI61F+e/Iy/sHl/QQF61YIjVLLwusFyyZRIPqh1as5Q
ofG68YrJ56PLTmg8JF70m5YQPe0NyziIDhno9KJVJHjpU4Fq82keaT6Nmt9xTIV4
5RgbkQc6cWpGv/8WBSUSl/l117vP2kxglQ+yGTAhuDdhwnC+OIxaboaBkxvY8nm+
AeE+HKwercqLp0mJlimNzvwhRq9N34nIAM5hvvG68S6OuLVDUFAg96cdX+krzk0R
PQHQ129YHYqE2BXOkH7FuYpEm1XnzRN+EuybNpwlaB744ED14slczz2+QOQUGsS4
+x6gZVEEx4laHRa2tgt/1llNYYrzWdOnOo+P6S1WsjYfnJAj8YWkLkvd+wbiLnl9
YSa35e5Vsec6VgTaXEDAzakepjyx//KRd2NiPMiR0dSnBl7yqATbBg063WZScTPH
O+Z8rJjyfPAAq30D5njdQYZRmHIeu96vDd7fu1R536iECmrSaJ8Y5mhNfCmvsBWh
WM2cdb9/tvZ6BhYUoLSB0up7vr3GNUqeKud7LQsryCQ/F9J1ioIEhnrfYD5JalnI
wnsPiJK2kh+MqD30UsACB+/z472PDCu3DhWXh0pG5ZQheZDHkz/ugOleDZKeOkLg
o1zkPwq7A7DaG5xqYsfmwQpZO08pWFEfdLgWkfo9pG563QZgxNzefF/i/LIBK3kG
waQURjDysKyyF8SsMFhkvdEp8jJBn0pGIsPvmLdq8X8OZa/nkBxy59YXqodg8Ipi
Lz5FjUytibsFD7wL/VmMKHxslLOvrHJvB0Bk7VNmVCjnUt6w/qIbCTX0MY+QvkfF
9yED/azayuMoDTJg2t1BA0ygouexcawBJa2X82OhMtOSjH6+z6FRmvF9waodxeOa
HHZj7yFLKm5RaPND2UMHEFdDTjCUzwx0lZeSklnsH1fnb9c9J3ULeYJmhUTp+9N4
4/RTl/qOApNyY9+Wt1yc8+JNx8thrIiEr0Kmp8Dic2IDN2UyfqDCVRHt0PT8pYVn
NvzZTWUMZHlYt7ybAE7fo2TCXv14yMfOl1MvS9LxqjzaURaIekjLrYWagJOKpJ2z
cddQlLmJEPogEO87HGCw7bt8krf1UPevrbzRiWMeyBgA0C/NeajD32Ytj7IsjLm1
CAFHpQs8fQDiTkdNS8K8O047xrL+qEDB9MKXpumy6hQbsTVWKQ0L3GGXLR4wxMp0
W++qDGoOe8vlEtUpnFxnsPjcQEhmphTvXQIWOeO5Q/KIufWFEIDhKc9Jlajur2KT
7CeNi0HFs9x5BLpDFYfkm6aaFO7wxBO9zkEjufcZGJ4KfJcJW5FDqp2+xZUtYYnA
C+FEBAdO54ObY7PGAyCL+dJ4tV2DaTpj7orHJ8Xd73DFvVkaWFGHYGNY32cD+B3J
yYTzL2KekxXf1VJmBzBnewrS6tqwUYo7Fr4dvkXZVYXq86jV20KbXNy3beel4ywl
XUkS3/vA2Bp1eQuJj+LVNywttchPUaU3RPOxincr49u+04rTpCzloDpKDmRq3L12
LBkQghMqiQgW42hdOTDU8dE9/BJXM84cgh4BIgsJd9cm2K8QhhefGEK7Og1Cwqht
JXzJqT69JaB4lcuZSNvW0pyYDfyAT4Jv6WydjiuMtOUg4g0RK1yJWll8WT0OzJy8
CqP57Eh4Zfd4j5Ujt6y/aOtiTrzd/1w1Adfyel1Hma2E2cLQK3PrY+4bvb/sw9Jz
1vjj8npJCL4XcwQ98r1AjnyUHmWFbQo2BBvmIcQVlViAkWsKKnWyl+XvSdhobki1
OTCYOL4139Fwit4lVd5kFFsDlrdDUW01+zZT12TqQSiunJ1IC30qSEO519sTl/BN
oLVyJ5pcOOU9VtuvzBT7rqP7NH40SgI9hgDEuqAQ1b1rykOW1gDt7+dwyTRUz5We
ydwtuwZTFPEOLkfehdzCVcjTTO/PcnVrwR94nE/kQFqfnsK4poMks6XtfbXGqUAl
84LjAvSV9zRYwvHYrC/eACBdnoFpSiDAdMsylBmFLzjnC4/FHVvj4tCU8W5YGc1J
VQ5Fkv1xN8gj1fPTEu3TyOoMEh7mku1ttIvr6BNuglaq8WrXNipIucJ9Kx2r93EG
3qYSZDUUbQb4b2owyGhmXpxqEwZbHkYehgBzApXJKNyzsIrloFAx+HlY262P/FNK
YebP/OfAe3+gb4ih3D21j4tW1MNY3dXIyT0qJqHGnWMpoRhevYJgfrj39VcAsYVH
ZobjB8AEW996SoiuSZPNiSIjXEcrkLTCZpdrZXM4zPZgMQTAd4BsCGlRNAIo3LXF
VMPCzW3XmkOjQI52UbPdoCfelfWThquGeMy/7Li/sn6rEzS0MJAqBKpf07RjQECn
fRkGZiENQQAlZ2xVPkY8Bo04y1kUw9vFClw9AxUCLy4MORHgLIs15NqDTDpjN3f/
EDSjpaM++3aVcBkf/xHCJ31xu5Xg99rwqyp3tJA8iJSM7ktlAIpinz4cwB6L2aAM
URw0srrZnhoyG3Hwq7kgXoqsX7lJbYyRJUsM2E0g2H3MQp48SroIqUxhrN63Sc7s
A6APoAJjx7O961mTUxrIro9abeGWmda7d17rvcntsUZ6Thmr1rNCtJTNEGMqfgP0
285ahHx42JntIskh5C0J+hiUFBvh+2wnDNGP4yo0eJk/OdL4sY4RRhfeyQ/zBHHq
x9Lrwl3klcjJ8oC3aeJm+Xtkw3DFhyNY8H46oqQ6hrS1/25+6/DYkx0YX3tyozfJ
XIX+maMb+5cGxywxUiv9CTHKAxt+dzTe44ZGLCvPAASqzQDTC7989mZWhBn0YIJK
qR8GMDIoubULG1rFkO8eRBeEYX8TMuWHatNspNYIaT/Ba8Obrv75CWTNGeAkbuYZ
Rd6xolLb7Wa2eSBoYtPZxbuvVYRfy7GhvY61UDMznm0+t25tVJh5gOEXcRp6Xh9O
lstAfVAusYPTK9Tk24QwdxympIbC6nJF0fTJIHiWOaq88aFLs9gtWJDjpHnxLM72
kNx9rtkPBBP4kzpJLmdMAXM8d6NPNKA4MmcAHEAvHR7wEW/vkPdy375NZZxpnZnB
lZmgc/lGsH8+tY2lQ19BOp6ZplNW8840y+8bGGE+VAN4QsMUmscE+mTSvTD+IY94
Gl2rxuaCsIoapWV33xnpVavwrrhKny6zCdgTAYIJOY7J5EwEEQqKKOrr4t8UoG+8
CbufxhsATSjLVoz+SRsAFbI76WVxAh3eoumJDLDFRHm7HuJekgzfEtYr6kc3gwre
TMcCkqyp6Ok5FsgSqPXXi3gRwmOgHepjGP0qpC9P1fINAOLBk/8xJl0qaR1brURb
2qAXSYHXm4BGwWE2LjWf47SEgR1ojfGhvNNql79AonbPsNRFy8MYm5QpN7AneRsM
kWI7oXg1asJnkkLJx6ZmGeka9jO3Rg9j+sM2rMrnLO+ms+fONco//0F28faddW1Q
008AgUHpsnafouKFC+ydlzM+n2RNttQxwxRHf97aophiLW1/8lcRWkP7sEQTdXMw
O0+IzJeFy9RNpJ50sL2pWkZBeLc6ut57P4msNl7zA/g5IpR7xLX/g/FCp6+suMDt
+XJXZuJXdVRurUc9nphjyXapUFAivINnZVCStKPPxv/TMx7R0MMuv0JVjNmaQTLy
B+heeo45pFobB/wbpyuGgAjPWO7Gh6gGkZp4s9OhJX86m4qR+UmbtUnaUixRxxMi
l0GVYcp/+Vaagh+0w0Bemb+YFpHLG6pUJNXeu+xvzk4TdJsEFbR5bxTxfX6gyBXN
ZOPx8wIOaF2ABIblU1aZs8FN99XLVOS5gg/93003KpEDmsl6pqH+5r/PCrtdeEjq
0FfnkbEM9Vn8Tu7P9gH5Bwus51nU+DA3/LUWbBrhWjmOExLSrfGsYIWzigYVTmtc
3mKRDlic/hT4xmAuqhRBByO+1fRuidVgnBKtF96irPUptJDTKJGYEedcOXAWrb0e
k5pLiHpJidvZTkcgVX/g643ei5Mnu738NvkTTPfs+ksV7n5UFjxqD+Vt0fvLiUm1
wsQca0Wdw+8cxbELDkM9WfoMZhuwmEz7eyk2TBr3fl7RBeDpvul9RxTrUuVwzKad
kUPBmq1wdTWIm6pzt9cf2nXe1BGM/+3ug1d1E71SbL8dMpmoJdjPKaRt84xBo6sr
sg95dU6cFCHguFWBnOMEzPRurK/d7GMBOvD/HRsI52HIjY3XymcxLfQ2SS4Et4YG
8z8LQea/jHoqTDz0hZsbYDknGlYRxCmfUu4euVLYaHzbwf8UyVWSnUD4dtvQ2QsE
ATgHGCW7yAl2wZaA6rUR6MU9T/Jhk6QUOo72KATIO4OzEFPTfqdhvkzU8iFai/5M
IQteJ8nYEVXI2xyI5hlxKo9iRu86wSSI1c8VjlMRq4fErFzbZSeTMoQ0wlYlLhh4
y0fLyJuKJHU2C1Q9QFmYZMQdybfAjGmVGe7tNMqQcUaLBJu3U0dVrndCRzyvLRMM
6VLcyuAz20RM6W4aXtit5F3InwBaaxVCtTV7QwIvY2f7FtmbJMRsQSVrLMf7vORt
m4hJrYS5ezJsVYE/Y7JVKOyYHA8D6saoBwxNF4W0vm5uL4vkiu9RY07U0Dksh1u7
RN3QWPLsE60uXJviejKVNBHzimahZgxoHjm65bycp/1SNIpY8DqXBTZdP3C6Epxv
fPSJD5AunlOkjHl1tGN2GI4Q7xi3sJCmsAej/yDcbRaT8LatsYm1++JU1nkoRfUl
zYqS5mDFIFJ47qNO77gIOsnZjxbSdbIq+0crNS5WNTjhSpdwQlkt7n9mu8xMrJlH
vFlQC0KW7ee5xVR3CUlhDy7L5rRg2//U4AsJ0p8Dxyx2kzoYsWUX9fqvFPcadcOv
S8uBHgg4JWjVTYPjt0rM6oiivrwaoHOZThEABZziZ3Al1tqx4Dli8G83C+/FghTt
5MfR4UJU5hCTrT/dCvFJdhqtt4Wdxdoj4UjUA5C1z4nPtdwCkVxOKSuldDbK2ovN
p4bdZ3EYPzdTGisamkHcum9qb/X114wucLg2y0xVAqlfNdBagwiXsvQBYL62dxDw
Ep7aaoMor2KKG+nKKuPXuCwqrNmuIn9IqzFmBNJQGi/3LcUMCLdtAKLyq3auCcon
LUdtkNzN+6UBOB6BokiBdM7t1NGKa+72nJLp4eBfx2nrWN6Kfsu0/W7cSwxxvTpG
f4GcXLB5NReOhY2DF6e9A58O2vX/gOcV8QzL9vQVk3ActPrVAgde2N7G+v8KHxD1
g2RWG9XkYEeNs31RP7oK/UyNAyj/T95PIEMKsDYArLU2TZvxsTCgbqB5uELlVkjb
iZGpL4Tj9mnmzjGQZM3GfQemUNj6YT83si580Uq+00sYwLPdv/5UGp5X9YgmfWnO
rovPVBxrqFZbR/Mf7evcVjFiIe1KQc1nrSK3cn4mMM8kDVXBUhRYY/9rvG2Hhzyp
D8mlGpM1kg5w4bjq0tIPLHEikKspIqdqMjuAR+OqL8yhhna460pm8YKIKML0BXCl
OKmG3jw3NpBQovv/ubazD4SYPrclULtc7xLVrfZAoAQF7G0vqBKWEZAsdHYz+Qf1
JZZ22kcrtZd3+h6p/Zic4R7e9RcqwKBDmmH0yJdEEFDaBTg4yF84RAqhofryZRxK
yycV8KY+ndb6xYsj9wz/INsiE9d2KA98Ht57v5pj3ajUlvxWYEfbChtDJanBNjxP
8uns3t3Z3GtAN3CoHbuqD/sASUDUbKB/EM5qk6URAZprVu2Vy48s4OvMWnwTPX53
vFJ9lSTKhrQ+Kp640UAo+7KBKCgZL0cmwJSyCSuDniEnZ1yQqjjSepknxY0pvdSW
m5bdy5uJUxrjYR5mQF3+2u1ORQVni05i99GoiTk/eFhEyBeukddCX+PeIB/cU7bz
KS1g9TTE8Vc4VJEnhw32OrkZpdo0OqBReWEobfuRyYM2Ym+c8b8dCeTV3IZo4NuE
lhlhbPCmiX+UHWfTc7qvxbQgQWzFdR5HP5ubKnE3+jk1oIkpCfBk9V9cFf1ivDmR
XhzE+28QGbo0ENffEQuordFGjOdg5045RkaZ2GHoNGHgMDYtf6lI34oknRyjdIWi
skfCsF5zI9UnzYZLYC43g1WY9MfNJPE96gJBbAPvvYUp+a8sJFodbkpioBHq5Xsb
UIgdH0atWetnD137bPwfrRynx/kgWt8788/Su9P06r9KMzeQ4NR62Di4p/6ifENq
ZxQub43RRLH5UKhnN3rt+rG8RVgETzHwUIU5c6amxCzfGHWFSxVvfkUyVLzFxTI6
WdlN/iyer/ecTQ1GX+aMaH0nj7l7BbWNVvXBN/Z0jWPmuehsttgqGtGu5zyu5Jfc
XhU0PtqDbbE3Ctk5+a0xyUVD5jBA/q58V5S8nxSEVAs3/tRe0lAlvcgs/oAKm5pG
ts0U0u9DApKJEOlt0Gva2XYlabiUKGvIIgtfbN/2LV+US5uEamZSS3XsV7kh/ffH
dRiOyhEWpPoVwAFjzzPJzrd0jwxQ2koCl4EvJgPAW/q3mJvnGF5dYj2uTbTvfN4h
IFMcrT2aA+TYpqfvqRuUgwg+SJ47sI9WaG7UX+RW/O6/89qD8VQaOq+eFmRuVy+W
osY/WOcNbX4CU8fHxSgAyPdRjnRTkcOAdz6bNR1youdMdiUjcX0r82yw1MfvgAYr
3FxGAthJHw4aVBe1Xz6yHmZkwxIkVySuPakLy5pHOeJn82RWY4AuKH7kshGJWXFm
OK+S5dD523BoVckOi/84+VmcKmwLlvhp0P7rMc3zk/POHbu1wUt4N58OokZMICuM
2hO23bPxW9q5SV9u8l5tV3Gbwl1sqTLa4l3hVqC2eLN1/8BGuHRSjF3KTnp7e1dT
af2j5sYsRtQoUi7SYHJnytc7OPzRseLOnYTHLb8OlTsYDH8Mts0H/lhVO/nH2tej
G5qJNXpvqkQt8oZgJxQWvBzIZmUfHd0ZUmPiEfO1cckKXwnGre9xzrdpxVDHUiie
wp7YZUJlYj+3c6IF5gSOy4nSUzp4/W1WzbQuIy9vUmu0zEEmRvNHvgvTd/8Eq+s3
5JV8zhPCZ5pmbvlHUsNBx7/Rnei6gVpIVNyyZAMiGjprHipq8SwSA2//3EQgWwfv
xfDO+So5kP+pFakZYQWIL0hz9tOMzjXDXyVG9V6/f1PvhzJmysnG1S8nModdgPnb
bWkgsyLh8Edb8HifiUE29c7n4zcGErq6ZMSyQ1IlVgEUpgShyRkhciHhgDIHIB70
hSTIGdfoOjOE1xKmOj7zUvk/9Yxe6TOLdSgSV4IIaU25vXOM0/pCvkxbkjVlJfwC
12rc9JDwIt7DRG4j+eFdpjKSdOlcs2GoB5urrQeUfmpI7Ne/8HtDHHjGvVdWBsq9
yXo5FQ9BkA8a3gE4o6y57qb2m4Uz2HNNkt3PT2HQOn1AdST7hwIjto+NvXMJ6YB2
n6OrroiDO201AokAAmUjCkaObKFWSQkvHUd06aJD0OXs3+WA+dUkA7Ci8EswG0GH
WHKo0EEbnpJz5b/o7I4+Fc90AD+ifygZJmCuOrtfYhdKWU6iK7+e7+fSdGnaJzKU
NFtQTkeuJtCumA0tPd52inegAyaHOElFHQDPW06GA4/EQWwAEW2LjVMpQS0kJqYC
Hd0RcAFmZ22R9pNlaTTOF1dQVjExXfE7rzZfhreS3YYLaS043QeO50Z5GisUri3V
YkASeRBoyM15vMh9QoOtWKC1gBMltHXVLI5XXw18UPqngnAoj5PZrtDF2hxD+7ZK
cmMstO4npT4aTvKo2s8Dp56dsFHNUc6KoK5Kid/0U2bala3HGHYzMrPaZKWETbP5
terHWcTlDOnBjj4JwgxzxhduwWWrrONyqaMXZyM6zY6ovQ7/PSOCZtwDBrd8Me1p
amtGDKwBz61cNdzebZnQlYTr/21FtxXkkQ58lWPoIlTdU8GTzMa8XdJFHP57xIS3
Ma2UHKh+5gNavnfzQ/68pLvp9AF059OKTpEpA7zpJb0EtWLeK+1A9GwKL9Bpwtih
W+BuHPXOf8qt421feyySWoZPWnp2eKF4V7fIgKWkq3VOUBaX3cu1C8bllE92U+Ik
TauHdOwVlnBZkem5mJzOfQHH4Ice4AajahLU3MH5RixP9C5ZGa2e9VofJBQK3WuL
R5pP9ZY4fCUwsvDB8gmVqv3eChv+oXWBmra5t3174zsAVCgHU/ir83xtCUjxuIBt
2w5Lou8AEM/H2E10GEeyvd80vmLjwjHB1RXuZWPqgfXFAknoiIvNTbYL13ewF+wU
5rp0BXSOfaDTxFsuUNu7BiBfH2TnS1+c4pSftGd3oe34Z5cFvH7NtbqtOCE5XRR+
9wMTv+tSJBc7wnDsBN3LwdN9ZFy28sWY/ToYVy7P3F5vU+9saVNkNDoIVWnSyDFi
xFp4XfXLbVdoysyWkX+NHmqQ/jfgBjTskXrADbQj5fG8WqxGMhhnZ4wi64QdINGz
ueH8kmTJ6hOr9JQAiVNXoiNsSQaeTd+fvukAS8idUH6paD/takk/l0sQQ0CdjXvp
76pA90VgpPk88Y4bv/ldYo7A/nMQOv6UgosNP8QO7c2vPB9Kkm5W2BXLgtsGpDFB
l4uiM4cmw9x6GkmI5DCI9LEvyx/cVaWRnOpBrBKgEveQ5iiJ//LfN96bms+bt19q
BzqeTMFgDGGXzydL6E7Ycc28Blc7LikxbOyLLKIUOHrVkzUUHMWGlqsrmyvypgYu
Bsr1jlrlUgvs6XXQqeGmr8UUsYzuWPIOKXSQ0XDQvwfII9QJvzqkjuphsZQ+A9lD
jvgeoSbifg4Kax2LsMn7j2gmlVnGvB6KMRmYS+fmFiAZsquyZ4CMtmr24PHaSsg1
VgROVeb9dLaye3mRzp4wSqvYXl9VrlBAcG0IZbnxnV9nnW1bCrMWdVjz8mDCAj0E
+zv3nnD5mt/DPQIYr6Li5r4hNYSzdaylY+gblIL6jdkH12/yhR4hfQ5MnnLtKB8T
1mPfx0gGYIXCqlFFvnRrT+gSk1AV3kVxlDeDDjX/mGGUXQZ235cevBE6oVSkIfiu
R64HfDCoLOrt6alc7+eIwx3U5B171CIi0zo0oGIg2D04MvXxhVqm4CwQp+mRzHfY
sALBVfDRjopx9rJZOYV1UF11+9jBk/lS4g44OgXRmTrnZT1aBRBYXfnaLj7l5t0t
LsuYpX+h8nOQ5yI7RholTnCp/0udSEGPhibV4+9Snu/frJuxpbdXglQGIbDEjnFW
y8SdmiqbRmzsdwkCjlaTwSew9xHWW/Sadaaj/nK8htfsNw8UkT3ujia+ChyB3gWe
j1rwLpvzeTFNsJ/O+e+ferVlA7xpgXXDsB09l78Gwg+7PzaXC7kp05buH7uSOEYa
3GRYnnCfLUU5T5TxhZ8oGZYbHAZB1QlvGRbTMYatqmhFnhGVOtITv8NmxS9ZinIP
hhdOKXLYcDRZHgYKMFC/Gy/92JD1sLcNBSAI81Cc6WGBSUm5Y15jFIMofVbsNA2b
PzcR3yRVCi9dEKjOR9ifSKJD0/94fYhUGQzoYe3IRUHL5uT5ZziyNz16kAlvJNbq
JtXpFesTtnn1dT68aF/S/Mc3q/Cfe+VZHWlzqhY7kknZKcg8mkibMY4SxP9DKxl+
w6ZBYz0RI/qCZJ13eK5orqG3FNZHypAouN5lWq9wJhpjI05qkjFn/VXSHA7Lreg3
3J4blQXFyM/Fqd8L+qtGzqBU+4NZ8yxpt/Ya9T4UisF+/NdYdKEfEGVHyMWq+ftZ
XZMHEp239jeU9ElPfb8+9gEJOVzuguoK7/X5g0Q11kTWdslplC+GMg44xhu5K/4L
1CW/wK/XBsGTtLLDHIrGL6IaiETKCLKXpu1YyF2tevmJb6sH8pkIIIFntHrqaANx
TAIfBtVTx2Vrdm9yPbPQLCWVLxbj4jBIBovT3fY5BRkBE+kxtG9W3aa6y629hck/
2p+uswxCgLwO/jxU78fwJ13fbnCWiRekJFxj6lyoTILt3xT5ieKpCZfw6hJnOdxZ
bkbidaY8TNDrRQwiXdYQ6Wimol3WlZPBnODGfrpwkLVscMdatLCP8D04MiRnFsa7
IbRlaZOiQyhY4zMnrCNDaGu8+4noWDYcHncT23UNYiMp/61taSK1kplwamB07P/6
0XfBHCOZZLz2bCuofKXgFPigfSb19vZ7JSllPtp9gk0VqDiCwnsFSQ4FOJfJDcj5
WKp70kINlpamPA3qwD6Mo6EcYeHPV+jCJ/pFQwVMaBwwSnrlW0ipgm0hPXbnFV4R
7TaxdGFRKw3vq03VeFOUU7n0j7pb/HL3M3+UeoRlZQ9pjZuclLx3OKMeMgOkjSQp
toPD7DlOfZj0b3lTMtwQ6/Xer2iHtd/pGvHaHUTG3hym5PIWoMU6iQIA6T5gnWWF
ssAGb5WyJ2grH7tPhhzJamuqmqa+YrTfghSmWNyvTntHl2/h9EPS9k8hIBpVlK57
fuXm0tLZwmOMEoBegJnHr0Cefq3CfOeMNbHHJWvhh7TkdMDC9E4lPtZZjORpOByH
oGE6f7mj8T8BUXXhAQ2Tg840hlcUC9N/WuVkRahDMlB3wFTGMSvGLdfoscUssZA4
vs2BGhe1PB/kdKHNgzFLfgnmun2sdvFuFGhHVE/IlXn27EWUuz3SzIecWT0FO84U
nq1IPtDWTPnwspsmC8L6jO4L335Jf076RGOpC2FnQSAE5u3TuJ4IEOwq7EPV8Q0g
ADHSL7hbxasTZKxMCEdPcqz80/Y/D20WtbgW0CbdxVRGxWEWvyruAy31le1mXeKs
6Nh1MzexpL06dSe0AFJi4ujBxkbTHWy2jcGK7dWsozbI2L4rRisZfGvpzDdgdH9s
4A9Y44NSI+8mwX/XIaGOBSw3gvxAYTptmPZMIKqNB7EJkw1bsVjVy6wDo26id+bz
nFEq31Lw0XD4Irl443XC48deEjepnsPj54LzE5BzfPbbT2SsUPok8iAt6Ab6nLde
Azc7qs2qNbd+MH1pNBpAXR8hhvtmcUYwJpbN2Kks+u97PkUxr3xSJwBSeV9tj6Wm
O/3Pnqwcn2uztrTJDZsCfAh+mVaqRdqSQyJnorxRymnYQkvIcFhlTlGzSHRFSbL3
9T8YZ9CMlAAAmpIRpg5tjzPR/qX2juN7/X2OC3S1GTZJdo+D9e47gVipNeXGZaGc
AMG1+AoA8qBB4n7+eWToa0s6PzNBdf4jk75NIo46H0wnW7HfgKBZUhDtSsRKau/H
Xuhgd0v+kcMQflCVtF+VJkB6ThPKs35A9DKXzqj4/JbY7sEhjq1M4FCWsYHKiESf
M65UGPnCGkeAQx59Xc/2BD0hamBsLj9NbA+TqL+LpEsruRlpypJ/tcCBpNQT4Nbz
E2ICRHdSLdST6ntILElRA8DoNRwo6hr4KMqkShZyxDrKIqKpiwtVi/dgLjzhEF3s
vurEy6JlJvwwfArmURrWZcrb2bCodrQocsiHPGpOvFH7z3LQPmyIX3GUs1xBTriq
gqvxjCj1GxmiXtJ3Y6OkN0FpnkVprQdMWdS2QHf3lQiLH2eT3xRiuDMHPqipKBYg
xM0G+/LFi8y1qDFMq1G8kqIH43GBvNS5eQ5/3DcYod5EWQMH/4yQX5QnHwdHg+JL
JYn8vmHymfdI7ykrHxFjoL6xLmbc4fP+z+Mk0eB5fROEFJmIU9mpinN61wjbXlPy
0lRNfo0+5oUbbLXEX8Dji/PlyICvYFtTJPI8NfTkslu3ann14O5W6hUDKgswKSjJ
N6EpTkWAgVrvoPC4FrBQXaDUvNUgZDdJ+2AOT1KbNf5TC2iNxcnpZRHC2fpanvH3
3Omu4sKAlOHYmxEwlTwJPuGtDShV2N5IV51FZV7RoIw9Wsyk+lZMHzNmEENQ+6Ki
4D9K5mwfM0IeKfInJRnVjFP7g26tnhNj8404io0k9eTeB3CS9fzNBnTCkyCEv0RY
k1TIrxovmTrtjoQwVrdXEKMhS4/RTP0yPNJRw+ehTdAlXLjy9c7R6ZjThbbq2hqt
/Js+d/QoAe56TEXPvFBEWEu80NWFRLeizKwRn1kl4GZZKpxcNsIbayIaB8v9j7nX
fbcr5FkI15t62yRTfG48YB57mEvLJ0LouG7M9/KCvGKqgqJgX3ljJHL1ws9uG53v
i5hU2jwcLUa1zs3z2Q4eIt076Xo6H1iQ6YCcq/j8K/usX3XF82ab4rcmt6BVo8eV
bGjA0bY7XQsdvzGjWGkpJMX4yP0eZiji/aDE+Y9rObGHjqUXhuK+gCSpDBBUfrJd
UDN+dVVaK9llI940XR4rbvBjb8eI9M+r9UuSXhd1SYy6Q+2xymklmDLWcAUq85XH
Te95zS7SBhktACFu16dUxLf0zaaM3sGBn1abpcwRXc92NwbSMQ1il5bQ3FQJvj1+
e10IN85KoCH5BjEUPZdoNoe7fIKpVV/HE2kB/A5W9WpG4Wp+NB9zuVB7e+AEgTM2
+7JMgoPWCa69+3lAKJM+TSFZRNhFTEkx0bOy2ovlOjEgXx+LXZgDNM8OIyaNemP8
TdJbDzJAIUagHi3q3S9SGiHWhIdjXxSwUZ1P6OXTPHiSC3kLpD5vY44qp27rDHCI
vAEb6KGp3kowLB/C2bAPQ0v88pbKaSrOCaVYd2k30Bvdc4acTcqHkOTkp7icXeC9
7B658mvQtePkocgToJQpaGW0bWKq5VYwvIugNa/toO0puqdYYX2ANYTJXAYhE9Z+
reJBJvb18Kzn02KkMarTBoq2ZfGJtFgeFbY6pN0ivK7t0yosDVXvy74ZOPYtfU3d
w9lnVoUhGuPwDnwYM8bfvQTz5TQA13Mso4nOSkd1vVUkcOvHvsyNGCgn6jnL/nkC
0lGAW8lFDFojDipiiac4bhqRi2bBfjtsfkfDkiWMtEpNvu2ADh12UIT/XAWQLBGg
po1FL7APXUCSid4LLqA1gYLCn5hM7d80IYX4fAtSXcrDhXiERXrl9p/1SoiPgn/p
aodnZx68y5anOjNk1byPslyaZBav1dGspWLwP9KAHstPg5TvpBy99U16UfYgPlSc
ymM7tyblMdkn22b4iVxk51tUbu80VcqqHMrH4KZpXelV8IsUtPJ1fz57USAK+2Cb
JG5Am9aKP1/ox7jbVKOSfCmP9bu5vII+lEuwFcfnAilt/zEo4pF2mkpBgtS9ORNn
q6nTR0KWMm6PSWD6Gg93Yl6Z4L6bWsJ67Z+2g8cKU6aiFcOYuojGPcjesJG7uWoz
o22TtGUc75mftQwizZRaFOwfYsvpeCssEFe9aqS15apOxY3aGfBj2Bl36g44G9M4
WZdlJrNYIRds4HUDt9qzuXovp6Ek+IpiGoz2TGW3FPXMlupsaJ5nMYppI1NEwiLh
3797OWrPQOT7er1fE27ybFVRW6ZAtFxXarsMoyElizsKkKj5wW9ybVVu6Urum3Kc
viNrd6qnCTO/nZre3J9AUZCPJnD5W2A1lGEz1JOVZUZfTksr/bQORpi5amJSSrTT
ZX78x+CSEr5frlUlTbwRRjMh1I79zUSzGh9Rn5abMYKWR3I0w66dZTO9E0W7rzU9
aa8FfLGm5Tdoop76ZMHK5pvcxtxkAZaSgnVsVVPGxXA3E3TKxoQgM0mRT2GUsHur
WAOXygPMivInHkrWwEmVMeiOVN9JJFrOxNkqvlEOGh9Qg38jsCTFMb6i6zyaW/sC
DwFFz8aVEK7OAgFqPr3QdcMgi6q8wpAGladJE9eHLhj3yL30GWyFVQWjqEoRsr03
b83b6rm8YdvGW1oYVxFPmhHeOONwsS2zGvKV465IOYB9XdKPxi5i7FWd7Cw7KnsI
al9sNup2aJWuUjGp2jWFgYwNAjbc2LEQkMeyVuCqf/j65SNKu8DYpbOeTRjXtf/r
Ntq+6TqeSLi8KWwDadKyq6kLWFlTrSyPhml7WXTM15H9bJtz3sSxluQ3+B+8p0DY
/t42BByIUfxaXtO5b+QJqnZHSxzSyX3Z/GHW+qYsP1G1MVyTT9wnXLe3x+8YatdP
GnsxSq1UfqQm+ei6pdtILUTFf22Anzd0+duxi8RcmN5ORVb8Ccwy5v7/syBBE/OL
MgKQpW0wkTLqxIYiOye3pqu5twH2R2gQjmcT87fDt03CJkatUhzQ9qbLo7WuapxO
Alz6l7K8+SzEo4PXe0vIpP9Mp7J5ny7vIBslyUAiDl0jOi55XMnQkbxninXRFo48
tvtEdl3xtBGcTb2ac88KX3sFdlQnz4MQMnFUB2yPqc/h0DhYdoezHH0HagF2KDdx
j9v+Jc3eis8/nI2Yr9IRcAm0FnVREjZlCpkfU71QsdAhOjhjVbXTkckUfGDqEAQh
uSb8pcil49+W0WP9AI9sBG7wq8KSOn43+BR4JfTAXsRYc8XtHWT1oc/L9UN6ikRr
PacVv+pZlgf8lsui54h4lmTCw5+Wet2olr1vXLCeUJDYfswYeLYI1z18YcObe/vb
pPkmYkrZjKDX7BZjVRwukAr3zAEbqg0d/oONyIjsQ6oHzRHHrwKrECSmHy415k6n
nsf/pa1v8pGP4L9VuMEA8irW2y8OB2oc3rtWYIiCp4LchScmFrqscoNxzVQn9vLY
8IYd9L0PiOYSppZ+cP+ubIun59WAQ5PeUmw51PkaxbQyxYpUzHBdzX2RJhR1p1JU
SPxvfXURMAP4BUMF8dsrmxh8kjqTmnZb4rr1lJYArmh82q7d+pywJ5bGuczUYTf8
GPPvFcOtkiLvvVVbRq8sZ555j5AS6fyLGLUT0iBYRhF19X66VMSD3S/MMX4GZK9d
8AOig1RvTwo6f3aoTjfNyjr0OPeYRysSYUMEV0GVGWpF7by7LqbqNBlg5g+5ktuA
Hh9k2OK6lqwTzUsUVQJCy3ngLQA6fz3ZMG4KAfwGOvwQknzWp0R8C1C5HcIh0DSJ
+htbS1Fyz0CbL0nlgxLbFhJXR16pJxtod+RaQBGCtSHZcjNE1osdP5/8CztgKtw8
fkps979YudmQ1leDKFQQ2OmRS+0SXKHGjPg+mcPKzahPAt84/Bvw87aSYTed+M9n
+7kAiqElL4GaXjDAYTbaASbKLE8/oskMip3L5ZS9N2NzjAyBi8fCmuvelLq3abyb
7bKBfK252ApBy8JAzrfttZbPqpZT4tqXU8AzTPgMyl1qjhXpv4mMbHZPTjun/rWN
9SwvN4Vc4gZAVanD2EDykafpb2IM9NZFs4M2TT61vwJNyAWLfT4Haz5PQe4FgB2A
V1Ijn50uPwyzFvo3V08JMOFb8AvDqGoCJWikVrjp6uxarYZ7BIGryeubBmTr19xt
RgiG9kkeGOTcPAdviDgJExoa42aR1FP+EnxXqmEj8Jycl4EDCEaY+94dUm+bHnTz
+98jKCEBdW8FudFlXe6PA/7Xy6yQPV29ykBtUfZ0C53LOc97Bd0Pzbuef0JBaEyX
zmT8Z3uIVMdr0VbsZ+uwgU4RF0JRtbGVJyQ6WcbEJe/gF7kDy4RDzRvD5DYc/hWz
uotfpl2+DOI256f5ujgeKKIgj4lcgxugC4/PNu1rl4FPUxwR0xvymD5WPfXPtS08
oHhNMRH7HCkT8NWKb6Lwn6wcekyJM2YJ3zZVeo7LaL24961OdQD0wIvqsf48/lAR
Oz9aI+BqH8h+2YiJGuSisFA3BW7v6Dmwm00N1o/tJy+FmA1KuAuozcKN2NzWo+VG
R2UvaH5UTd0hdbhtVyTUrqLtBxT2hBr6YhZsS8ZB2cufD2TIGMu4YFmSxt0oKAxM
LRQCVZIlPupJjR+WAujBVbMCNJ0zugjz4R4YGEx9IBfWFr4bQ8dR2AER7OrDcz/+
AHA/oy3rGAH4lrqSsoaXfXB45NQwAjck/Aw2AD+SiXOW3IFqk4JGr3nHlXBpYvSe
LVh36cK9eSGHvpdOUXWtGMz657dAGqdGMcSware7lAJjcLBvPyhE4tTMyUmh2UNy
fOxE9kL7nToKUN856Wja6KTfIdozsrnmreSx/vohkQBQscgd7Br/kchiUrjRagiV
Nkqc/dil/er7LjIrnwsYvvJdaQa5lQPRp8XPDoi1oY/ZEPB7Lknj9Wa83Ods/LKW
AEiJB9Xb4xSc426p/h5GIeHSaF96XqN0KOUkLvSZDVEd9cs216Id/P3ZMo3jOveB
MwKmb2Z1z9JFAf0bD6L5uzcCjmJVGO1jgixqyVSCY+ShIoNaZ830Q+f65gD0BBY+
3i6LM3EJUE4shTpG6ZmVWgmzjLjs5YLbiEN7zOMcNsiUZimG5bUUIe4fa+a2C4l6
mXtQ6X+Yhz0P0UyF0a98iz/o5M/Y4Bsy9DB/cXVmISuzvfVxRBTE7ZIDm6zLvtBN
/u6pQ0/2ewzmKKsX/jNGGNsArqPqJRTpWSqT+ZGgoGSIO5SZOwf0gRNhDxImhqAS
uKhxte4MIEGgWvMYGrwZ8XKTRyWw37NZa2HkCgsTTID6/LWJTedQ38fsLv4TxqJD
I8GVYcfka5AAcbU0t5LrPJEl8lrP63VFKic7SpFitkbVksvKx3Dl0Cg8Xb2L5Iot
xeNPDb2LIplgm1ehB2z/Z4U6UQZBK53LEYgXoG+Pg+1s4uY+oPpIFXdipSVx9GgI
UTjJTdelKCbMYQv5io0GHTF4QlkL00LqvzodHkvb0vQxzlcv9w3sua9FdUsJ+wms
VDZhDSoRNRJNOQ7Puiudob3Thzink7g3/otZ+s9rIwKdzseVV+rNXC3pm2wa7Gp1
JP6Aarzwxg/xr+DBWTyCQiwGEYvPOCS4Khk/JRy8+tP8cGzK5vMEwKmesbp/4TQf
5R9mWJCGw7qMZj+FkxOR8CDPA05Yuyf2aW8XNeQkkp2U2UDpV6l8I9/oDTIK1ubR
IlQJvIZXKjNPWYENmd4k6tLi7BHoRtpcbF4KMvrRMifZapIAY0WO5pvjHTb8I6Ri
ApM3m9ZodpW/MUvJU7zwkKqY5Y8vm0gZejQe7lksuUD+wPiZAy/Y1AjESEPa1UM3
houELXHd6Pp9rQlFQwJatnGzlYpmIeY/Qaq/nYf5Cq3zMZUtyFcNga2bt/aWB02L
KEa/lcJIkL01iDcQoDBjCi8H15/x2EmCuWeF/4giyRPZ+YT6QFzM5wuC37IiiG6j
vlnR0BQw0ZPG3Uax/3DR/D3sJF9KZk+jYIC/jgQTIhAPPaHm767DgldJaCRPi6Kf
qqAPJu1ChdPt9jcgBi0SExa+BotItjbBEkeYff3CGM8LqWlHKnGJ8r+ZRTrIyBz7
zK39jW/q/tX8tgYTJAlQct4FIz2TMgTZRzLUbbnEloSs15sDJHSj+9yK+iOyrrcA
H4q05kS3p9Gz/mR/3Ar6cFeQ5vXAx5OQ8DDCPaJsT8WpQpqX4aUr/5TtPR/eHzij
3wp/OpA4tCaEACN/0Sv06bQQJAtrwn2scYuDRZtjtiAI9ZzRxLjW8KnZpBFjood+
GgmHrsK2HJ8Esx/hczZ9pWA0BbnAImU6DcMycvTJv+3VrhvxoFp1Xwn0zy+tsgmk
ob7P2/8mlLy5Z/1cXsRjiy0NxCPnvrY+quEECKUH2vaaRcIRh7zCPfGJaWo/+bMY
xhVjOUHd12r0hkyYTyfhuRfcBDZmDmTVlwUUPurwaVQlnwr8TWuFQNALlbsASe3H
JhDzFUSh450YbZ8ZngnugsRcQCbJ4WLtY2ufroPmwlPelcf/m8NKteZsS0hzs2Kr
Pkz792WklvpA7qpdlvzpuTAX5Io1LYJkKl+rjRBqz9tWZh+1MFbS7/P9Yp7O3/cB
j+goBtw2asoDCrupGHw57vVid9rnm8LuBoRJdeg4Ii1Gy2zdrhJt5MEPWn1HyOqW
OZRDttw02NMSnrFVXkGUijbAz3d8E+sAP0goeNkF4Rq6FYZKbtwS9H7blCAstKqC
rk6GVnrl4zeyqIyiaAIma7kMavwFkVx20I35Gvu8TkCeHBOsiLpwE5SSsGw1OxsI
6qARKuibxjSg14iKCA3lVgs+A4HcI7O3OYTRSrU4F6OyqUviOZ2K9oAs/ewIRr5i
DdKndlft+pyS3GbXUfvXdCwJgoFFF0JUvMWUDZezU0RCNXQJDem72fsK6nd3Qx87
Ppn1w0b/RaKPFPhuIFhVkALkxMEWQukpZX5rtsHCzsKy0/068RsBqOE2AISpou0n
XRaJMfR7CEEtLl+CNJAwd4bSX5EfIOMD6T2pCSgDI+rwpkMnGpwr/ZjqHsy7HJlY
+7xYp3yX0ldWQnreJp/En5B+6IW7MWHa2AtkrMDgkTmIVF54amcyjHobhrT+pUbg
hj3eIV6YFiYxAfPOAoKjBITxsgJbpEWG0jmCq/orF25vweyhNFUvsF3y3cQ/bPPL
9L8Cuf1nRqXuF77EofaqQZZ1JyjOKGAvvJrvv1/6Np9q+KQ3bFI+O1Lcz02O67Fg
kTY8gozQAKy46oLinbzkPGAO/exU+85yt5TFeyL2hjeoxkGj2zH0fgdTd50t4T+w
EZlKbupdg2iUZOOam0xZ9V/YfJFynkMED/hdmh3Q+ae/WCgcXlZvnZyOxIjAkgtW
04RfwQvsHJKMZiu6uEwAEzdNNzF19bCi3g4rJPpBJGtRZHBkT5QHNuOR2njlWyt6
ypCQPiDYxQZ8IU2ko5lpmele+dKvBS4E40WhsSzbAprHOnxYCrTaM9/SqhFGFVGn
YpyNdbLrBOu3jt5X5qC49RGDrM5MOMm2/XspX/hXjPF1r52oZNb8PWzaf/3eBZFH
gdQJgwvFhqPBO4+GmFlciXewfMHjTjGegSDbSw4x6Imz4YQs4iuEC9UB2vcIueaD
wFiTlPwVnozLoO3Z3YFMoFO1apQQK6TIHs5vlhjUQBPAI1RFGHHV/gwCLNLj1jHH
IidFMkWDZou56EOSuA2dZPzshlL55wFS2OJn8i17se0wXt5eNgJTx5iUl9+pH972
0b4O+AZgUYg2XUIgnqu3dW2QjwwTfaCyfzgMCjNBbVWMxX47nN70dQZHxjzRvRk5
l36XsQ8uLZr/eMRtpUpHWMAWrvQ0RyKLGlW3ic4WnPpvi8y+B2BQEH11e6AUPChO
NM3wYFBGwDupGhrzdZ1BZgFHew8f04/AYidwnagkZj6mLI3f93o0kE4k/fedi7+A
3Zl7HuHCxYEZvt1Op3f1ceVx0j6YtVFjjDAqXRRoIoXlOfcLWOVMXQ5WWMlDYCsX
uGP0w/ikBDZqrfKL5TLGwkxSG5J+koN4LUBNg1HeU/GzLm2M1Gkqyt8+raWDwmHk
JUWxZOm3VU85qT0kqK2bU8j+Hi32keDdmx4Sn2Y0Z4xNQRH8yX5nEWZM2Ok4LbGC
d+nCpuEecK7633F9v2GCPG+f5in6WLi5nAIHR2U/EgL0xdXQqOKov+OABRBepLfK
vixhTY1qqPFK//bEE4GwxLdCq8HKlT+QwzitOoL8JeHQBM1bLZ+5OfpCW5AK/fhy
nR533/n6wSBQUJHzmBFxgEFVOUQZ12Je4A58uya51abb+AX+iuGbUkctpI4rYxbL
sfDn/MVGW491j8s/+6jQeIoaDQ4mo4My6hddwyUGZ+bvSjcXWDhECdXreP/ty3Cx
zgb6CPlCZfri//kFG3Xr/EdETWii9KXhZ5zCwe30hjvY6Bb3Mo2K9/l6VUboSe1M
ihby2QUDQwAI21c8r5LdPOhP2NEkgEVbQbzfauwc6OWPjGYCYQQb0WdCBLn7IKu4
gSFnLfIkga1uYq66zLo8wwvNl0Dj+iNaMm1FW4FREf6wBokdGWtbCyZeiDX4Pxr6
g8OyBC4hDIoejttAtCr28RdCXFTlbFh6d7xhc2sEyqFvA/8VmobIRvqTvGK43PGK
mkygs65fWUGkP46WSWRBhFyIMhOXy4Z5I9u8cMG/Q+qX5UAx2+gMDYyamr8Wc28N
JRU5sxAT7k2UBFGf8EG4asSjeDEDa+54jg2IEBddmZwEC2HyUT4tqyh3G2Lwzrtn
EjIwZtxmBJJLeCgELFKBLEtWic+bD6YiEoQSA/RsRZHi34PgTP1bb3fflWS3Vj2k
i0dyHjPC+om3RUu3Bz7rezLUMhvw2r8cS0JA/2/tQj5fivdywOh34RMGPwTA1G0d
HrapM7xmJgxDc8lTd+5Pf/m7oY2LB6qSVWiaUm3A28k+TckfXbLh/th6UVEANZBj
UU1eyDPhM7stTFlTJrG+K9rrPWthuxNjn/CQbFdxwzL/3oRT6aJ/RjzhCwG0oBCt
vIvQ0KRu/tFSnDtQ5TGq8wY6gcG4jspzTF4+98uwJWApFTgbLqQKOWM3OYCZfUub
LWTci3152DlWysgNPqNlibftALdLnX4XnGFim7aijEnzzl3WuHlSeROj46DRlPu2
dbD8QAu+xu6EPMbshWvpmF+eHTPWfChzHzUVmsvyRV9nz5fj5bPjJHe1ew5oqRlB
KHp2JT2wl6tefLwGr6MH3nxSXi+11MnYzwSXmQz7+KchjrYCbxP+4ETbCgIKnKsM
MHPby/GVSeM8V8vxaT246ofdunoIqdKQ70a9NRUHTWXVsOKQHnKLJvi8aEC9uu2X
iMASyDrk+Fv0A1MiKSydlmwQKoAgQYw3gqQYBHSV4D6pT2TV4k3GMwafzgI+ZYM0
mtls8WarmUGSrcbkwx5jAo9jWS1WMz6hPWWvG9W0Pq/Wj34j4Mbfbj945phgv5zr
2Tk24U3WoegJ2L/NS0nyKwt5E7FEhMOJGu/2vbHyqpfDSa4YI1FfmU58VunVqgnG
Vsx/8q+tiDRhoaaTL2RUb/pYcdgVegp5XegBuQYifCq4QlLNGq/SjqbW2n2CpN69
wOPGCUEr7V+n3nS0kwUQ8CTZ1OwEk/kivuDefKKvW8Y5hnUFAwaYdMuaaTXsbp5r
+coKeTtV1ylLBqfkE+nx1hWlaxA+Zuq92fqG8qQBNMptyFQOW/6a6U6QrXKB6v9H
KCNAnYE+XBlI8zQkNlF0KWtlPIQQOmcxLrC1KAlHqmogWi5UxLSLN/sP3evp16on
SN3iOvdGPuvExDQuGDaWBaUPi7B4aojreHSryZXRoL18JTG0UXQLzaspurZE9gOG
aTrayuw+9wIEmJVUN/wmUCP11Tazua7RupXoMazxYf1DdNnKP/MOKH4DZyeJNqd6
hkwSPLj1V5SGwePUoGBOK2QrvY0pjjejCpmJOlNeRMzrU1SHE96pOCp0RBKzB0se
RSWOlWqP0kZ62x4pSrT+pPJRyhFiMpkTI2kdP4vPoR+M9hIpPOpBqsGMaVCth8n7
2STWPMSqCLXJP5dCLrNH9PD3GWH3m2a1AMZ4xEIUodVh3NoNuZh/k5xWt8v0ixbR
qx+4dduqbbHDW98XfrjPa5tEUd9NgYjFJTVGQvaUqHO6TYsUIaRIhZIsK5y8ChH3
lQPMqCW/oAnAMna+UQTxabpkbq22RMD8aRHMe2LhM5qI37+zK+1znbQPsL5EIEfW
AY7cLgy4gvm+UFIjR8cRbqjsGpQYspN+byrUBcLkiLDogLRBBwHNq7sbjjdNCYEn
6paafIXqR5yXqz9xcUNKPVQJSkgOiHIi6LWbWlvTzTeuu2S3JLc+RjHIPrqjrc9m
/SH2ivLG0CCE6XRqtJnJeDEWcKJT0R57M74OxKS4eYV9UBNOyA/crPPUat/TvXsO
qQ4UJ6t/xQ0UOqC/DLVlQ6QpaPvVGp2SmcAFexP5yIvk+ICtO+rgxYFmyrRpR5Od
HDh3kM5ldRXYuF5zXXu3SX8Usg01FDFx3N11rtwDpmdmf01GjJuXb/dNjVhLNApH
OqwmUWwScEXQqDtxpRfYsmBqXN5QGAZ+UJi6sPRn6CDDpscUulRe5s+QQHwchNNT
oTEH4+chIIHIQoTNkp3oBJSVl57SIBRQH7+24hTUKtQZvn1deyMrq4XVGqjbWg6R
ce/FQ5CyriN7sMvq9OxCCllgREcQwp4gPxstl7nQTPC14ClUxzQPWYt0SOTNKp4K
hCw/iVL+b/oQXpXvKF0zTK1eS9/Gzfy+iJqoXRpoU1m8qr/hO3e13n5w/OEWF7Pv
/R16pR4Tw2ZyyHF8m84FOGqPhqsYMQUPdK+G4bCPQ1xVGJHL/vOtYYN5yNeH14dq
jHb1xABE+zGUFppJLNknlZnasaQ2cDqfTalqo7h4yDJpSGlR6x3ocedqq7bEEOGH
t73tvOGy/CnBs+UdjdKDmWxkF3x12RAO9MYXLOH3f2fadb3z5uYOIUkul847NVac
rdvMp53AYAaviheFnae7InfFg+B/JzfW/A6+DnNt8L/gh96WNzYEe7v5/dKsaKtM
b2GplsJKsiN6iT7ltms3REXQQfVR3y659wfYli+430sGX8Z13D0Ap2FRlxbJn0ev
RNzg2cvg12VAMQvBAoobb8mCj0B6y7KsjyRIBXjqJhW0hIKVvjm3pT7ynGG/DmPe
tX4m9CWzTOwr5CJ6tVc1Ms491tR6oOmM8oBMjwqM+UXtH6Xr/xdspzHdNW/Bs7y0
WOp9uAtNsC6xKY3TEfkbTFLKLgdMENSxY/ieHe0GlZ2TwfKnlWkHsthmOeKW9j6a
5f/jf+cgdNlJ+BcGeTo/W8SRattA9+sZxsNETE2KzPez8n5QuGGjm8GTfhVTYVZs
9YQo+qZANpeRrR6/U1FbE5CLnyDzM+5mIfjcPk1sU7siXyDiU2t2gKRGygNMZPvG
DLxWSMgFqnLIF0on04b09D+f3ZWR90Anj3BlmJAz0LgvRrPQU5mI5UiqdmBgsCJr
gZ43776xEwgrdHvmdENICHJzXdf8Dp1+XmvREtlp8Lh1pGH2tCgnKSycZm7In5wg
InvOFezhoubZc4eUJ8rugsa8Pphx4NbLH+JqHqmmFUrgL/+CGzzYYLIJs2KcP0tC
FqJD8CFH9tNhzJVHYvjxk1Oipt48vpz2rt/Av5wunzWTNq/eKZru97rQCOZe8Bq/
Q7XZK/Pxn46bDYJmIo3k+L3Don+zwFejjMVOcCDsUPkNgOwN/bWHyHjMm6JYKG7d
yxAuTezgcro8CmKrtEMkIjYtZlKN1jf4vqkzzdHYhEXwUXagtfoFL3/2Hx3LXapc
Eb0WBz1WffhSiFDwnFKaZeesE7O6iHMKIOK1OImrtw812rNtqyI/+YfcrTytp7CK
ZopwlhgXAh/c0cZZJRGbMqgzZtNBEWQ9fHyztucZ4F/tGhcl3+AnnwGfIDOdkWbP
8wraSdw7rORYLMdiFV8239sfUl4KuAG1oC97EFp3lJx7dp0m7gBc9MjHMIlALXK7
A3Px2FH3Te5xoFKkGPIF7p6MlfpLLJZm8tBt7zbBME1a7ewlpwK5vDuI4Ody6qMc
6bCe01DDwukRt3l9dqg6jKrHTjr06sIsx1uSrJyeRfmpPVSRZlMwYbneVHB8TM7K
J8D727gp8NR4rzilekBj9d+NiaI/rcUzUtbJZsJt/ca2tL4fgCnxEMCtFute+9PV
f5qiASkwZFmgEddqaSxyx7MPKHOQ43DvAIR7eycdlkTKbJP2EKSYJQr2ggLEbPM7
ROaTc+80wGJ4bATtS9jttMtvRdBPIC29AdJVWmBBLalwVjyhZdjaRTNhCpFXBJBy
jxvE7AmVaQ2TtXLJ5h1MPonr+EIly8+xwnr/PNZpzmu0+rJDdo1RAt3E0P1RrZZ8
bKiUWnMPdSeUknYLj/TwGsEXocM19nVREu5sMcVYtXjDjTR0UHDIilxtNa++KLsc
q1UiXWwGPSjbzHM4HpmAefgPW6ADfeBle/jETGM1V+sPypKdrgM+8YQ3t5HVYdpA
BJOuXSSlY32vVNwK81eiaRrA4xfhI82jLdK+lQsKIsibYFKnB+lpb0NYJTZbHQDn
f82pQ0RlIq0KemHGitYgw322vpIhBhSzgYjic6aXTMsPGv6Sf2uICw2pB+/O8FRX
JZ2oTaeQYhKQAAG3POuwZSIE4o3KsfbNYdpv81+mjtRbEXysJH6COL2o3/VjgVi+
6ur4mrmdUwXgY4wJadCPfyga0Y9e7ZYQPpTz03KBodkoDvIS22URgw5kxjwHru7V
Cje1CSRDDmG+0dzUMoV6aoUnWnioitwWlqkty9AhLpsX8nCpgdrCVtXiwsJABHP8
In49LjcRcwxDB2Q34QHbQGt5lqqUHowdaflIShlaTS9w54lJyKcPlgcZJmdt0its
M1QJo3E/lkj3b3rDiKl2yqULPBKCDl0kWcAe3BIelvGJhIbbdNdoskZyAcx14mjY
IfdboMb5VopCsqk5WTCjH3pYKBZ3WvH5KRIxTLTKj5l15e3T6UXBBTvn/s0tMXO4
zwO9kPaae1gIofmkQv2B7tWTOVEnrMCos+KgOXDKp3bPzgjr1OT0tP/407S1/zeU
To8NulkBJ9Q+ABBSs/YfybHggLrH2SWkYMvTTY21T7j8gJXbSc9Grxun8Xo406FO
/j7P0Us7UnHeOS83xE5UJMAU4FdgykrrXytrgTNiYAsJetIb2t44VXrfc/We0FCa
6MEyTkqcEoMiYEvvsBzn8jEHWzs3YA/YX035Vzs0EHlGXrQ4rmqNAp7dWEmt2cL2
6jKhx8RSUopUFVgvm+YYypBMStDLJftWcyxnc9Mmk7hEzFESk6zyIYJOHCJ7cswr
r7AH3Y0Or0kO31uf+ZnwGQA7InFLVKWP33csvwdWJgwJ+BP/UAu+X/LNDj8mHNmE
o3X9fDodRBn3IblegHyRHfYrSsemF8dq1vxMQ2K3OGn0vI6hDtQcqprXeM8xDmsp
GU71uM04sw5IrnTZ+TSIK6iMWhFnJcH4DCWZx6govj+A9A2fuUq24U0dMAWEnZ7y
//CEaY2cN7cnqa70khWGqxwUitaKDs1Gsgzd6K4UeTt/ZdNHpFqjbDu3eNS/Y4ob
w9zS7jEDE1+jjMrLTz3R/P+WZrOJ0rVu3CkBlKpLHHEeoHrFDTB9YV44TmoOrqXp
cm5JlYsxLkiTHgvBdMRhah3ypEe4jkUCfc25qwH2dgsb158SNyu+3+Dq6Rij4nx/
TxPE6B2Xe7jglGY251lJKB1Gqxo2si1ubq3vNVcWs60vsBXiAgyQRB+Jtw++lX6E
ln4IMCDIz1Ud15O/KNfB7LsSexVopYk8xCuahf2vVPOE3zX0rpkKj+RiW0AH/U4k
9EEXc/cuSrD27XdDLRt4cPdo7eMPYpSu4V0gqKGNCpghZbxqab0cjqAkcr4dkNkm
PYFrtPVNFd2rRAkKyDfMR/j2Pp6DoXXy5eLjoWPbIbJ80zUjk30mmeQ4gXmBRGRz
EnxBvw6a6SM1wI+xobUajsaI8mAurJrTKdr9/eP1lgy5IHzws0rDv971xns990C9
ePKxmObWWzvzSaiIzyhurC8BAcFRu0c2gb0hgW/DzHfdG5sa2H/vVK8cyGOLoMvl
Kh+EXQLTJKR2EmqrOPk7cMUbDYRHGts/2/DA2W2ZWH9cf1NFed+yEJEZot69caA1
T9hBhALLdfjAmqZbdVzBzrtPuSJWEE6lq9lzM10UHSFiNv+IE9XDih+Ug3huXq0K
2e6A7smnEnrsuUPyG3ZBmGoFms3Or4M8xh528g8g7WsjkUEi3lmlFiDsPURTiuCA
iW0jafhvzlCqtSZqU9GM5AKXFAKyE3d3qmGwOwbyKkE50HC111JgfLkCx/FAlmRW
XKS/q+NOCMzjX3Q4BSUX6EghyUoFMCKzLrgVTi/JWhvJ7t3/VcIA35AY7KN/SX77
8Q0NTFNkn1CBSVFCZmLK0fHbTJCFD/j94+Ufha8aBpAaY+9fDmdmrDvNyAX07Uwn
34SjX/VKMCiVBONkuB6GFnG28kWrP24Wx9kYCMe+dnQ1O2jOpvm+z+4EWOSLgrIF
AjHosaZG8XpYsAKDo2FnhYhrW/btKzi+ftO8FyNucZ0uZSdr2EGwnJAfRDUe71Yu
XJOGBWeyxnLDY9gi9kZdTVolBFITaRX+cZR2HMnwfWsvzRdlLiro7pd3C3BITD7R
Ep/M+Jjl6fZQPiFstofxMFBa6uofqK18KQU0sGWPbK/eNpo1zWPWc9spxXHrebTF
pX/MzdLQjl89SF2FblxW1gekSfcZsTy3gZUTvDJsrYpT0N3j5gqdMRWU1sL4SafJ
gHuSV8czYQfdB8UurLG3YOtI/Cb1Hz4EJ52L40bUFHJ5QlYBENWSYu75ilesQk/f
Jcc/mLcbedBmobmsICVWMmSvqXX6TfoMfJidRbmuDwyC0Ngw5gKHFAVDq1+U6fNn
rpf13txueFuTRO5/Abdyhgmq8evoqwj01uDAAXZuFOuhre3MDvlnx2JrIKDSEL/K
yHi2jeN47tpwl8w8fYATIOTXKGKttuG9T5qFdmp1KUXax4+pa/1/6JYUA278Jzqt
5C7EYBT91bSUzjtHQ2GIIP7INu04rkRbTGhKwuS08irPO1QU17KPm2g5EFf+SMd2
2WMtULlnrfFH83fJxUfRkhw5SVWjx9OHRDTrFFwhSMcf++t+nS6J+smcXquhu/dO
tHGN1cOYUEu0onYQjcjrl1YIKRi9nXOu4YlcaR5lKO0l3/REH/LSaOBvjAEVP1oZ
OyIphExnnL7vHO0o0IUGGNtbQau2dV9vea7kpaJYDCkrlTsMSiqWeZ8HWHDp+Zq/
VVcSNWvcBXfD6l9pvE3WjZZMp9DD309TaHOfv9Qk8RmXkTUkFiE1/oivG07y5iOw
NgGMBS0aa2glIsbbWxU4DT9HSXI0R9c16Y1o9OP8UFYHjvdqX3zPR6hBSZHGOBlw
Py4bRdwNNb7hbdd9SZzmuKCd0Hd4jzqrL0UjFUM7gJpavdeYZ2uuOilwXpciZb20
TzHXLy2TE69c38lxu6eQ8XEO8241yDnDOIhDIUCf5zcWiRACxPiWd5T0qJdEOgg4
S14ZjtNMkKi94zCueau6uFuyPHnRFe1TlxrEPYaCppCfSZlvHdnyIjasfQ6tNKPs
26EjZrQSbQ6/CC8yTTp+JIb8adP/G4isQFW1iKPGBZeXsjIWVP/kL4ikkAx7Q7/g
gPBQd1Rx7FEP8A0/jzNVpVXUOlPLLYNp/mD9uV6FUQ0VIjkV0W6mBIZU/alBZHFe
JFHOqKrKMg69Zd9kdQ4rTZ/r1IZ8TX5S2/aT3hS8TNCzfXvQEtCen9So1iLd7fdI
r8JXPxhKz78ZxhQWZ/79Cc19iIJjP/AG6RHTeTDqoxBGcOQgZriNM+vQOSRILrpP
t0BvFl14pXsx2IZaUGuWziO27eAT7TsgSdg+Z56RPi7BNqDlrRMn7y5SiHb48QNX
r11D7eRE+vZc2hOAML2gN4/uWaw0puqEgpO0w6XY28uZrLolW99cQRGjGqSkjr6Q
BebUQnoGRMmpFAhJf1wOuG1VCtokgBLhsntPhybTjpoCve+vT+ACK6CGOZvgVHrQ
7N6CmTS8nbVlGsaU9nLWx2jqCe/9hQzkkTwdQPswuT13dRJtHZyMRojSGrTZUPIx
B/+KDae3J0J/6sVRNYw0CnXlX3qcWSEd12xlx/9deWGFnsIbG3NqqJmVRpMaglNv
x9blpdSc6hrFtGdbTJh2YSfqUqkfsl2FB5ixX31/AlAtrVXZYEDocR201SPtKbtb
Kohp8Ald4CZHiaN4Bbx7IYAIloh6Q0yj9CUMjXNg++D0q0724ONkj4CnjEjRELNy
vcdMyTmcBwBpJX5cmqpM1HSwiUhDQoLGGmw07usxBODUGFLZxCmMYo54EO4Xr4r6
HFTtyOziaVal2UhrSkh6M3oF+CEiPHLBdAm/hApU2Kk2e2jWGEwVO8G+JfEPIMIj
6Dt2nn/hhOU0ptlmOD5N5tmKOup/aoxXYXLn9686+KnTNUDu+DONTQt5Q4KyiIsa
VO+twLCxv1e+Dfop3vK1znSYAYYOg6a+slJBCo2wc2G/+qEVRb5uWukhPHB6JDAN
WGR7YBIGRSCncQJIHYMXAo+4ZdkSwUyHcb8QasF8iavLsySDXF3PDbmY9LrKYNCt
7cviYd2HvS15Div72gBOdlePZZlTMwTFc3PUV/iQBdAIpT8l4vbm5hXNTt2iiwxK
79t6Rxsx37tiQ0F1wQfl2wxw/OX/VcWCVNk+94b9xm/pd0G8tRZBq7Wz4vg+DTWQ
d36YfXLRTXLmolwvDwQIui9brHvaZ4wkJMt+8BsxuUHtEqAN/xUANmlzTN38yEX2
owZb98MumQhugF96Yyo6Em2gdVazpAhzdkp6hQcVufgUWzvjXNwy4SP7dVQReTAA
BRXXfG6FEOROtDNK8oSJmgUrTBMBjA69DEK59/b2u8cgFLhpSgyWWTEg8+FrlRln
QvAEJ5Mqtf9TTN0pWGSuk7336PYT+vHjel9OnmqRAJU2feY4kFxCoqDiRnR6WwEU
8H+fZNWRPKEqNdNDmFjaXs9lGIPFO5NgtdND+lIN0Hpt+g9s5VSuq7B6hYJh5NX5
zbTD4xk6GMMIopmC3Cif9Dir9fbL9IHru0SpJhKGgzlj1FP93PnUop5O0wPHDPzT
W0dXDZ3eCdSdl45LJDH6QV+mOrtx/3igJbkA3OedLot2EB9uYdQH8mVRz9AS3dqr
pilBah0P8Yyz/2FaRzCcA6OBLQWRe76cySRQkB8RX77F1w5X3s7QCfXRzU122q3q
y4V9c4FV2FjLIt7Qc5+FLqWtun7E8xZ36zxa2hYuOZuR5T/Qr6YHwWSEeROvw+vV
4pYd/g8S2uJMoCArj8OCH93e3rEQuxiFKGYEj/Cx5QV7D8dZaIQxuJpET4yQFiMZ
MhmETi9g3Z41ED8f4h0bEXYnoDGvvHIxr7UP+gRh61tw89zfIfdKVjtkGQEzJt78
jniah+0SfZl+DAb3Gs/9mcOY56N1clxMJ3E4TvpTnkNtjDWotzqnjsVWTlIg3ZwE
KY34I1Y6nygRGdeqyBSZMAn9fA2bV0tgghKRGcMs2N2E8Z0NV3Nng1nKVnfDdOeG
Qh6zHyeSrFUCHh7lbZHKZA0JPjFNioq16w/eA8oWUG2xu80Be+ky61ZUQ1AiP7Bf
OUJ6uaXxnDXmZbvrx+g2UmNZpgrAzrhL3EctFw/vnBk6lkAWlFKyHkKPds9bzs4R
Yj33MZOayNedXOQjQLFfCH83202IHPyRAZg3OPSpR8644DKO8JrdvTyxpnTNgaK6
lZvVhynUhJWNdVoIDW27tdHjZ1nKq1xpLOkyEQUwBL94o2PSf6orOFmsoX8pP9qw
1BQl+2daUZJRs1HcDdGECMpEjjHsonbxz7YntkOSa7hDje5nqLFqDk3PzE/+h5Tx
HMyQXrcZaqlcTZ81UGY9dQXjEZwNquGGdS6RXea7MnwKeUZCWn2ErPxuv74CnuoF
KBmlJ2HEMDCxEsRz60u88iw0JTSxAtXvX1PHZgVLmkqDFwBYoLF7lG5cAYK8dfP9
nsvsi9AqPRiQ82e0JQI/O7tJM83wSvOmGfJXBZw2jXj7rAZn5jAXc8/7kiPfyRB0
kYPKZXjShP8egubBzIymZ/PLO/2Wa8jl6Wa6NHGZ5bV2aE5Yu/QLbvSciWnx2XtY
z6fM1S1IxjZpySnk5K9kkKTB3sMHN4ucq1iThCJNeRm99cxeW+13iRWLloqB5CZW
+TfLhn+5eyinLE59R6J8sLruNLCFtJMQBa2z+ZGN6PmGLUrehgZ+n+pVuWagcH8K
Za1fGKTa+BK5omX/cAZFjHj4YtULXNn9NTT0DOnyXcoDcgLf97U+W3a/AqYquPjb
uWErovCqDQCd5BzAuOubCZdtp/1MeTyW5VwPX8vNRAjvZYBUOoikCHDlLv5VFe92
Lay7ET6h7bhE1IQv97K/SvWPu+cBp2Py/abZDJX1/Fm9MyaBKFy91s0NJE0877zo
cMukzySfGdSM0RmCHrqwNq4aVGFA4ImkfyQzMIYAuhVplFmPtxq+7BXuMf33m574
NBMXfTK4mJUAlP9K4JhjAZxXhgK+1plYqhGIz0GmIkBXdU4W2R8v1TtLzrv/GopF
A8jIslNYFfPARb+IGTieI4EMVhvMdQNSaF5oqqpYF/cN0wkEubh/r/XwdAj54yj8
PpGNdwWX0No5S+CavFQhzKIH53JfwX5OtTCzo24LPfmlTuDYWLxfzOYNMnUuNMbb
v1dUBkNAzqe9XFJx2Y7aIObppNAWetDSKvV0ZKXYc30tJEqMl5f55mio+Csn+vW3
27q8yYoHzH/cwYI3K6znlqLA3Ld3QviOY41EINczEXtp0tmnQvfs/0WljFZTN+Ys
u+o7vPGxgZOkE0Lh4pH0RutNWxD0LytUTpTwvQZuU9ftTLACTGCalf5QEd4tiaw0
R4tWrmaJcP2w1uRHmmBnLzotdeaRZYhYJ2Q+3/3RWPWg106Bl4hQnGqR6eYNTQEA
liwiTmwDdUVye8/GGWStW+DbP0OWAhPOCcYBTUsvstN5J3h2nH3XxctC/0X5kCqi
kEYAX0r4BkE07WYE7s+sYa6X6AX8hb3XaVurhOK3ExO7wvdiQsbuoXqCV8dfJljJ
saPiQJZ2eN/IwvZlYkFRzYB0OP+7B5kJi9yv6eaeKDytjQnnysRAeiWBfV13Yrbo
B8ExuVJbIXSPDYYRHhCGR22QtGnxnrjWH/iuFphPiNyBw+hs8/4Qn1sDdRUbKrhc
jnBIWa0LYNyR8YTpqX9a0ZF71LBfy9gr9lq/tGNolhMoj7nEDW66ldC7VcQ8Gn+D
MmtXzUXGfQuworKlct7HGxwfZ/Vu90qvqcToxuodm4Dm63R56CSpdDttx8egr7yg
Qx26bRHNORH/vEcamygJQh0RZpoJcN+LNun0pLbXaUCXJugnkirYYbSlEqZEB73V
Sb09Cp9XW9h8idwE5a4I3h0xc1et2GApkKkazn3yI94ZJV1TAiZ43qU9KR3e5x9r
pNas8FKe8xx1Yp//3Ok8DrtIR1cXllhJzY5PwQA7MZvcWL8klTksj1Non8iyTFcK
WVaqL8/YojQNBq2srXSuqnu4WRPfrFLSYqnXiMkKwfyj+md4YltPZYKYtkiIxqq8
IhfLZ/gapgQ6q3lwH3rIPZpGLp6ad2w8EkodQaHalWEPlYa2koi6JvL3KWL345UF
CA6N3qOBnGglYZewNMd9WU7CSb/vywZC+pG/WnHi3O2ml1eQJKYdmZNIqnPFOLE7
0VVUdnOW/nWs43XL1RHeJc88E8uI8Ro6nQpONRf0WxojkzOHpczUy3Jk2Mq6m03v
bEWTOnfvnwDymAAE5iaqEPjIqAJzMs8aUmYhuIeO+Mtt4akrA6l7lHrCkvFy8d5z
pcl+p/LMut4ZfZytajqNE1AS6HIkFJwXk4ADFjsgKvFJHZ+GXNLyHoX4AtU+/IZs
lT1sdQK/5yMLeUBipaWAZ7qW9qeszRlM86BOB5VXY00/xM7MV+xvFaNAiYWvEUCy
SlFkchns5KfR5rsOKS53JyCGLGZg8SFn0IBX/tpUP02s7mqRYjBCE8V6FuWE8/VE
ANqLCZNAGRptHjyYj9uENH95vDVOnjxThk7dvF3vzh4sIVKp9Cf2h5ZAh6pQ/56F
Un3Dp5DloxhQWk5KvmNku3nAUzHOCzwpmHTwptU9RPXhjaqAEavJDVg3pekfU0ej
+Am1l5/pC1tb2/6faKdgjhJXXEsmaI1BC7STaKTUbu/LMRpI/HIgIMdvU78u9/IS
ye3Ls+uMz51Syg3gdONCwZ7CbJDb6VCtyDWHIVZAW1SEOWRjCZk1weBebEsIVVpH
Kf05m3Bmvo4SyjMZel8XqM4PkDlB5ILKZLJP3JPujWj5qS105x/1bavANm0mZYbl
uEAR2jFMUQUUhKjUlQPSv2Z8muAsbt3p3PYYMDRwRmLQ5oocMUmLXPbcOmYPJB8t
JUysYY4Fv3MGLIkJ2UAultKUrR27fABP+57m8rqYX6RxqI3Xe3qUtjB6skYECmQe
sPxxKC0+CWOd22z0zatG8BzQwhFeb1YQRyqApbOueTbOaIQHRp1sZXirWrFS3rv6
1rPnV32yai9r1deW68DPbVujPWM0MTnCTHaj3cV04hXMspwhRUU+dIkp+Utd3/HM
xikHlWogIONw/afWnsLipgJ9kZyzxtcqyZLK3PjDVkhBP8aVnd3D6hJLe1+xTNuE
Fv6CePjjqTpnoiknDI6nW3zL/CVEfmoa5vN6J8zmWGmUTEXZeDOtsTrOqdRTzBEp
tuV3sEtwCBOZa0UeziL0mM0/h2igFKVXlk0MvRk5zPRNFOcxXFCZdq6StvUrgZmZ
C27pNbhc7VNF/XIw07iReBVNjHDTM4WifqfC7+Howqc3t7zqUHUcmQF6GgrOurN+
qVHgOef1YpTkMOHSR5IC43Tj5BZn8jA+ikKhFabIY3XPhLoQJadnQ5uYaVS7Gt7N
hcac/vNcAOucGw/rquYCuEwJtOVcNR24XotrwZi8bsB3nt/xxuKVVAMxAp8/ELpJ
CukNSioVJ9TgS3UX86NHG1+flk+lUsjj4SCNvLkmJ9ZEr0i0YbbU2qBdSgFP6njf
rCCBo3zcg9u7rWvRfB7MlEfu2eSkGL5tTEefZ1yR7hNzp6NfbPWabDjT4oxGJACc
AvDt06NGb/cig/6AAvMxlYA5sqlO/9qNdPvTOnfXwxlbqJgc13PLrmPWAWrriETl
gEdk6r5TqdNuYPnwxAnD1z+dpLIhNm6eYqqqWakvSS9bXKv9LJWp//Ro5QUQO96V
nzF05UJoxU/IRPSbMtykM3djtD3dB37/5hen9Udr+tgAP8jCUbF5TpXEDs6bZ/uR
R1V7oChtY4PlDhChCrKBp9mRPLCrxIh9ZsBkNIQHbRXO88SOOxZT8eEDjwi6+O3l
QwNkrv8TYDAop+O0foTt8HIDA+PY1Sakkd+oshgkiED5j+dYzI3cjruMW17AUk0c
3eUhF3AA/sashjNDEjPZqn6lf7lXN4YRCSfiL7emVRsGZHqWNuicUS6+f8fw9VdY
sDt8noJB2fcvwF562+gKJWJ8rI59MuqmLuxpxEAAdD7YbBmN4AuPA21Geya9XnoP
HEJRa0ugAzSWTdWmBLP9/j4FLL6frYZA+kqpoUjrHpAtkj4OYIosw+gwV9DLuiht
I3R/0nmuhvwnJBuEiilMT9c2NJ6teE2Aj7D3f3HWWneBR1QdfdAVF0xBnEopeHLf
NzuRRmvOGdIPWt5k+J+uSeAYEpzzrTECD96ofxoTNXyGSFuVDnPKvcjrerWrZLjK
+QHOVExOLZXk+36qcexuMDYs/LzV2in+j2rsEqCasLJ25xsh8iS0DnH7gysOVPjH
WTKPVuhEmRs3Rzg0Tltimal+t57bHJY8SxbVGDz6yTRqL7AI4W6aOmeArZyl3CYP
+EkbpfhzuelLvXf0ExvbTMQd+M6v+haRVUhC9UbtHCJG1vDf5XloyiyMbg/+ObsM
HZFLMN2byD4CRFjcAaCEdITT7NrC28fimsiqPqMbdPx98B10njmnO3v2Dn9DutBp
zmRxmssds2A/t4gWPEXQ84naQ2rfRXunfs28sWnya7qFxQnPM5WeK6gfFC6j6MKR
3nZ7iafoBLnYZZkoHQ+dawcpQur+dGEZKglhTxpG1oCI8f/F/yXEQ1ItBEXQp3i3
NRtT6yIDZaccyesNNiRSq18Qn44B477rxyquQm9tN34ExfTFrZcrqlwEk2Bv0RZB
maSP96FGQwu0p2DOgVKmiO2cv281frRlO9vtUy/HgCUTLDkUGuJjAThOQhcs0W+7
EXpV6jYMACEvYbzhTPrvV1eV6inijT1bjswJfEFRK5m51zTX6ACR2G81lXzc6QVl
lkXNBIV9Q63Jxg6QHFABplrRlvNHLvyiptyUPTTyaojr8XAEgdtXe/LlSWROjPgV
vC09ZuW7B7VPi8Qt8cDYXMFBzmDGUvhEhTQA/dnuzEN9pgaFxbdWFUmnMkXYnGPi
a3W0mnWPDZscsPGK6H1mNbf+joRAUyagcBJ8WOrShJWOY5LR8JyuDnWDpcn80a/7
ABKJgMHuzfDl2W945WwRDLR+1LRvZwLejPMZ76LK7O4HEhiW7/PQJHjhtIIll8U/
2QeHKFFyjaSUbt9WXLFobT1eKSMFy7E7CaO7THDH0i+CymEt3U8YEtZ163WaZblX
EsPZAB+Vn6X58XIQNlkkKUiq0TJISHSqdj9x5oBWbiXSjdlYqGeHNIAZaEKSqmP6
7l/jWTNWCyR/rjPGffpXrtBHTRDf4fVPiNFxx+lTtvsx21zui8MWtRDjscDpLpNX
0rDe/ANjMz9w4W5O6T1iMOpSZvh9WMrA0vFGMM/U1NHzYj9KEFear1RQuRux+RG/
gayxOtw8Ketcj4B9e4uYNScxcn85rN+sL3n4zfpFGV17UwLMero5SV8Ie5HgWJKW
4b8Z5kYEUWhv7JyiRs7IvUANQpAcvWVBnF3aUjy/cwsF+LACPBj03u9/S7Xxojyd
OzS/abSt+m5LyVaHeLYfqcPyT3h+bE+E7lPHXpJKS8lu7JLJJWnLc3k97tu3Pzby
/2pG70sCcmD0VIMX7y05udKUSuYkOzvwdobnwPRvY90Tk0fc/ZUm/a9L+VVgFNga
HCJ+3HMi81WOE6txdzMSUVuenuOtzxz37jf/e4UxbyFYf24FQqtH2DP80EE/FcO4
631whtuZdl2zGySxUibvR+Rf7dONk2N/OIOOrtLb/ujtDHgL63w/qP//1YxT+reT
nDOpgobqmwMEsF7jxO9LPSz9hDEHNnvDg5J075o86VBWOSHtMw9YjrubQYtAqOTu
5HHOS/EoQfMtcslZ/PZXr1IYPSjHRhqfraJeswOPjdURliU2IU5vL50zb6N/QqwL
DOswAsh7yhUhKGZCl2FLoBteIEJNLhvftf0jkaAsy9cqUm3CUB32ttkTnHGNtn0F
6WgKSVp4CEYJ5qUPiVfvEteJdULetaMw/b1D8zQ0mqYJaMVYWwQaoQbbr3k1BXuI
uEXptDACbjPzx8wvQ9/VsKS++x3S6jmAIYuvDOrlIFruNXYhfYqFNzx1xmz5QmCm
RMGBYX/h+q6kyAQXSnBOgkNvBVgB04dmePwuDTcZTWlef2SnmTqv5t1Om2fAgMuT
MxsdMlssJDPxkZ7sv0smrR/p0KObJWHLvu0NDTbojZTs8Ljy7MZw0ghypgliN/Lt
kk5GkX6XlZTi6vftOY4sgdmbVaWenHODA/8r8Mqu9H1YDDf3DFo0nqUBAa3RB5Qz
z1lpqBVPDuVRkU3ot06m2BlUuuqskk+5LMMofMPNMwCkDJcpC+XetnuJyq4GpLwS
Hgk7NwWwRuB9+nor1R1hQZoS+xPYSNkJHyng8nFllUJikU33MVtrTycxrDyf4eMo
gvmUiyQxsqO6QvKr7V52ZQEFYlwoEEyiabKTJnzpFrCCuQ9VOCc/0JpMbDkqR1aM
IKqCXYTKLj1gWw9tMZ63roKEZmC9mhiQlL0Ba6aOhpB7h02BjnbnxnL7G9ONP8dn
lxp5Wr1ESE7pn9GOCJc5h22LwX6oQjKCEc92BHX8wAyY4wz9tDnfWIoRsE7eLk+m
AyQi9mBzFMrJAtWC5Me2SbnxbWBau9ZmLWBuGtF3idIP4ZTzszoR+HOH+FQDp/CP
XqToYkVWUMsJzynixpRBZnCBmOyo6slO7nHX3EOwRS5qK5XQZPKzWemlG5geP8Un
Fy9NgUitkSbuC3JDVMEfKM6npJ43ZKzF64LZs+k3YZ/x68RDmxRlstkua0kUnF99
1kRd+Es+8QjStg+vHVu7toANpco5saAa35N4b6Ze7U5ka4nqzvg4g2HUIi+q2QFa
l1xzZqbuY3yeg0h+BfeMVxq9n8dhrIf8g1lgXGYxX058gxbqW5tBjN2lyvIbAm7W
lc5VlHakCVbADFM7VbZgUKQjo5O8BEvEQk9yI2996STezi1MYNQ0dMsD6Bb3Cf44
ZZmRr2QzgJMaOJ463yipOAgWMoinH5tVwi4O86vtWA5hvgx3ES1siKPNMgpiIXD0
q5VlXcZ4Pm/HpUaElKK+zfwBIfxBM2xE5Cz+MjAY6SlCFfXyxJmnvIhZDlob2x17
qsO0NQ8M3zjTlO7lUk/6U8NISGt2dbG6s+JBaK36wIRzgaAXNOA9aX5Xhr3J0h35
xLovpFMmO71cZMcHJKTC/gsCdsJcQAsP2vmb085SO/QdQkc6aaDWIgyy7dB2296Z
0YB3PuQU5MzA9jcMQGJky28tT2Gl7kW4GHVBnZTTVYdf5zc+CTNkZavA0LKg+j7N
mu7jg0Hr+plsNNInNOjCdz/vplcNtAuvzKtf1qmTmj9tZ45kNISLN74Fmx7Ik23v
iqteEm+jQiBW2e/2KpMmS05lNeEMsL0DItXcfAk+Uo7oIgu+/KtaUjKhPmJv3A13
iGhrpDccfkQlCXH+e8woSbv+OdPAOqdsSrpchd9G72XfCYC4wwNMZey80WeRYStv
YhotBzGIHoWBBarccmo5bB2CZ6R2bHbTTlt6gytc3BOdDefHsrbmmERZ2CW+Qqlx
lhP6HyR/9bnbE9bujVwQUBWw7HNPp71XQzlXU/6/rUBi3IpCk9nrntjsJZtAO24u
IYG4OujYe/ZtoMvn8YCE7hGIYWD89yk38ipfF2z3sPeXKSWD0BKDrHIjzYZPwSEO
j4k/DvvztHVg14wfarKwdRxv+JC87c8HVbNghJWKSV6RvBj0g2NRjIpvq5RwgtdY
5OvRWv42p1FIRZ7H+BVSEE1fLYtt2mFk2W3/7Sl2jvFlvK7lKo/1X1PWJ6623tfj
apFAQ8gNS6kp23REC9ho5TVa6iWP8jNxEkP4eZ7xa0gNEWrB8QcKfLObokSkPpni
nz06uIlbgPtElFbmFn0Xxdz9HoR48PrztfeLZkQyO0sBgxQFP5O2CiycuAV8gWKw
6PDQpUIiG46cCuSyNred9YEsUT7Wbxr4dxYLOcptLf1FAd7ectFpG9h3dJ7XCIw+
xW+fHIZdRnCNTt66LDHQ64ZmNzhaxdi/k2O9PoZEF+4u5bkFgBTIHdtSmphvMXZn
UPS0u1gVPpQpJvhV5qPKC3W0cUqL9zB7EcBIApme6eN7CsqbTbfexMX2kyaUNSyg
EaddQL4ZhQjMODuD0XLgbgPPE1ADBn984tE/ANu8QvSfzoY4weNXQZ1ZpiFxSPpG
LlNO4rN4JEvtKAkPgSKRMDDXcXQyHysg7I0tF3UDWw1YI04Ua+s1/z33oiya7/zd
FJRU4nvRIpfY6wBEFxbRp8Me5tGZRiVlKnZMwzFODQopvElKaOaZLZ+qIgVceATy
1R4nIEIAlNdmJKiqHeFapUJ7jQexMEokUKxUWxebn3n7QAp3IuU25PoP1AwZyQh7
v/YFk8GLtRbZBtuI9rj3cg2jMHuQVeV/oU33W0odV6OIvEXtSCkFg8vsK5gGQKev
q+Ugm1vL574ClyzIZpZpuIHpOGHhJFeSUxibdeeUOldDVTjcJJztbq6M+wuX3yNd
X0836c9ps9IOOEIAdIfJ0jDx9aPXNrHcvu0Zi0lPsv/SF1pbHi6NbhEBNfr60dgM
pNLDjdawDb5A+RepN2MsN3De6Df1c1l4nLE/vB9x0VoKw/pu9CJEzSA73LPzUeL/
nIiTwIh1XbqEk6gwtBG0hC3geF+8g110nhhQQlwq7uPZiDVxS4SPVATsk4JY51cN
zCL8jdovwx8tUdtnl3rftxSsp/DHHnU5QOhvN+fvYdY+wruqqj6DvakPE8BUmwdx
tpta0OYqODHcwWS7/9CI0SBAJZcRjBRRR8VcK/flKEx0N0QiR+j/xk8ajs01doRz
nP8AbOwtBFgSkqqCYkfQxaF2+N+K44+3pGufBepwTPDZxqGmPBL6p282wYGbnc1V
61QKrKhks7k7/UzIFbCbt0bSkuHd57DRuuTON3mjmTTJZrqFJh32e8o8A7chrAQS
quSP5zMgyWveugaab07NyWeBOLxSwDFW+3eCJCkQwuvmWTIDI10pApWaKlz8XEg/
fuGxdsSFA7NO0BBLql1JV2AZTSGLpwayiOqaN5GCUm72WTKbIkjec2274HkLKWTk
k0ETkS7+avmGF8D0KS1Hiq06Qq7mAd5NOPKnZWR1E+jJwdIDQr5u+cOCodFFgf2U
uyYV9VHtJNCdgiAdj36pohzP8yYQbKNzuTfd0WFM/kK4sJRYOJTprTF75ZnDoqkO
oP5RpJb2digMpAVK5h01S5kV2HL8iYioCX2jNa5cIKuCMjNH58hC+TP7m5pvS2Of
f14igLrNDLO9AyX1jMN4sZGxD8yY6hIrkNk+Kv3+ImI5RvD/RL8XWjDR5G7k19dv
UrrOqnCKYFWBGgY92aWA1l48VTZ1qprcsppLYwHAdA/eBcAqnYZKqbWSycN5MTAZ
PxRYWbgHMZYgXlqVo7t6MBXClDcvKYezc6xW83xqHcHa9iHlvGWFSXkpRdPv1GRt
C7AycjbMoi1naB7VrP/2y92oTdbZwj7DkuSLAJ1PNqntPjT6J0Lvb0zg40UBo+2s
Scm2/KMripta/JwYSkjsw8wB5BmEaTmgqpihxviaVj6IkT0orWaHvXd5ayutLtHa
G25iaqQv7N+01l7P5tf2pfj6FtNg3WatalgQXeNgMpEqIWna5ip/AF6C0Wl/Vard
jQm6tUbCtbv8Ydar2PUy4H/RkbY/jPxsV8Q8lwvX2191M+P1AP9xPt4/W7/NMXmD
E7wxbdzvb1fT3b/iInWFpiafsQsHilv0JmmMR/3NQ6eUppoujJUuVNGoOzE7Ap1Y
INT7i0UQo64DiQH8ymy0Izo6YjWeTgRWsiZU1hrZS/xygMFCGmJlmIzvGwwycZvw
ZAOtl5Q0NceHRot/NnaQ6DM7lGVUoPvX5mMbHfbANKQwgNFIPTUG5IQoP8GojuKj
w7K6PGKQM3PxqflTRKFa6Q7S/ksnj3IiFYtH05EKUIWT79ZUKZCHspuqoWT31IYw
tg18l01F8iYyMkZLgx+uyA2EwJwHnpAtYHJBpGFwYbop+Lso7BR/fx3YINq4nk10
WDtHTEJS31tBRbqAOyjnR6alwixlv2KLRNY7dZZRci7oLXpzljWUmRAiB4cA8DO9
oROl/VjXVsZvONHB39OlVzbLexeugKTqXJZl87ieDrCno0GGj5MvmVZHdGsb/Pn5
hdYbUzoCAkLiuUWO4EjbDtA2UCwIyOSd0DYtBbcbieBI7afwFkdKpDSe5KIdf87K
+C6bV0tpMrEpKTtKKdVzpgAzeaxEXr8UyMlkUyL3d6dUnnmVEL3OD8woLUfhCsTk
KCioa9tYxjQC4Lgk0GHbaj2GfzKCAMwH4BhzCh+OgqdkCXpMGLxKzgOgWEN61wY4
uemTw0Z6bTaQKGDw6SQvOSrPeBJeriOU7K4kKJZzjhJ2ZQFhrvBhE3wDuYvdsIkf
8qTG5fb4gqWtqBN8DLxYbmnfxokLOCrusZebWEhlRjm32VdURYyt+mm7p2f33lpq
Y40hiy5U3tPxEVwzj/79RHRxibx+Xl7BKislWQMmp4QaV5TE/TdqCwoW5V50ASYR
pU9mmpPtFMipbAYp8MmLxHyZ6yK8L6fLuWSiW4QY7RPlb04t7lfrzHDU9F7Okg2f
x4V4a3dRvr6iaoBWhIFYzv5Qx4BehyV3TT7yF0ntGKoEa3dVrs2SNW46KKsO4w3G
CmcQvnOHRdyBVIcOFkiBQDok0knAJ/HjDr1x/wDs7hGWD4NkAeGTfKWLHje4rHSP
1e4I/6oDwzB5MSEHuKUc5RLguEHo8Sa2BZtJxMBIMTdQnUk/YuhyoTRwT0+VJ+6m
AOlygfB80k3A4ystvw5/4q7sPzT7sVGg/xe2ULZ1dfleNQTYteHJ4PjzyX14HsG4
rYVgnZ0Limq25FziWN1pe6dNwyayPsqJq2MhiABOd//K8ky5IQhto6q8VvAH4Jhh
rAEtJa8ux2vKSQuDyStrG4qSOrW8kfMeqHbSSO1nD0tMsRhKJqWKYZ9k0opWh6gn
fu+2mX2eTiBPGFEYrc9ehxXUp14PnWYUnzM3NFZBHWNSWfI2oZpUMjJ9siuW9adq
zlwGfY0TIm8WsruY9cgYN5gZ6WdS8tHw36sHFfa2mGup97i8OPVaN0LVa/GyzFeB
rr36W3UiFt0BY+vhEkcBPhXoNPAU+xThUeEA7DavWSO67Px+EOmf1FyFeQ+NM4L4
DyMgZF2askKQ5BU+Jl2t9XIYmfuFKE4GwWex62Wh99RRYGUFR5W463a+U8EC4Cm3
mvOVcxYHn40il/sgq4ytFTcHlkfXJtbWLgD+2u/UKZeQFtr8RhVRoQWH/vWdITO4
Yl2KqzUayelGQjPYmsVfM6uyJF49/k87zntD7nm/l0eYj3WJ1WZdcrJ1+ie9pMUe
Fd/JAftvzdEaLol9tl619sfcUxRHMKLnJGP/qOJTbc+pyf4FBANa0Em/SlhuBJLP
/1KtPNC70qviZx7WqdIxKvvAk7/DF3v5R6DY4mcZGqm40VDzgkftFbOCNZ8wPSwA
MkfqpoShe/pyNyllygzDPyRUFqimVWkwCeWwdKpFXGk+qg+N/qWz1mperJMYwYJa
jnow7K+5/SoEC411/NcEnaRhcQafaFvr5/xQgCdwhE4zoNy+bZ1r/yL+Ufdu1a8e
mp8BBiSYioyIt0RQQ5cpPGBSi8hLzMOlwaSpkF0yU763tYg1BoeQ7jbpsJYW09fJ
pgpA+4Du4DhpG3j6PJuU6d2xz9RPbMUEB0FofnaE1T+EHa8i0imJip8roqxx2BBx
tv2ZetIr7kQ8MlQynIx+A0M+UrVPPvBjhp313BfO+vBaZRprVoXpIMJ+1siRAqjQ
HvJCOfM1kfa6+TVyf/yqRVH/Z06UIQA0E6PHjSZZwRe0jU3la8aIwr3ZI6yoi85R
dc/kmBUsajnCBIGK2LvF+1PoSWfugrbipR/rPvuhl4SM0EHuP+td9WUrb51kXmHW
XceYHADQ7eGP887hr7ojJfFEAn4MSqIEo5n8QH366kKrRRibNvHRZs2mwtWYcH6s
sk794kwjDoQcFoFf8lbXl2DGbkNEhCAQDDrTTHtpxPFV/8UKxibBq8CjMyuuqhyp
BpmtB7/sBWoMzu98rupBr+B/P02yWWofiOz3w/vz9vAVkvBnkk35qKRyR6fAO7lb
RxMGGMlP+2UriWJRwJ3sBETwvooNy/NXRMer9Hbhv+eFTq7CN8oQhB7fqODllp6u
Mdb1U6dsegosoNYcsHR704BlQNQFF1Cj80xaHbHnn1rAygJnC82rRx643n2RyuNR
G9EetuusXkKnoTGxCgUHcQyT2PZmA234Ww2vK5HV9wZhXQROwAuTjCrEgJNnDjUI
nEVgP9sAUSpP+udSLw9npj+MzpoddUh3KrB9qXNDKjkWeDngvvETNuLTeGE/OBRC
AaijVKSlBygp8Htqqg1pTS/T4x6VRDHWSjClLzXWVmqdu8niHMIISBJVEKy53BUg
Xhfi3SIcX296+nInzerg80+JpC5dPjFleJwSA69eAGxuVBm6UGBSuDAvGevUg2Me
FbgMr33GM5B0+TflzVLyGlcZLloc+tJafGdlCt6z2JcdbVXGlN2bhEaSk9lAvSN6
jm2WG9gEr1PTyTaJPsG3iT0INMwLN4fMKauXJgytEvnN1rXRDxaxT/0G17Njy/sn
49yMtIewszfySl4/aAniBL5qBc9fQQOATGOgca0QJZ2AfES+sSMn4aKv+dNmah15
9UH3nBBaCb73I0xjd4XIdNwAB9kUDdTORqFuOS97+h8wXnlRbWU0l95q+VUN00cn
pt28nib6qMjaRC54vcHDzTUex299wit54KnpG852Kogx65y1nMa8HmLmJolq7/Pu
BP8v3/ZZCNt9oEAmb+/kQpSGTqfEiZZs0piXOiqW8v36tSiyGsLmvrQF4exm9uTk
XKrGJUo6pBWQPTVRU+omu/NCQeKJF2DNvI/M81oDYEiwcZyfOsNBiV5WOkIXjZ8t
iTvUMYI+1KcZywMUlra4C2+Z82nDvB+rPABD0F/ATNU3Zh7WhMBpffE/KU9JMHoO
qAy88sx6iGQvfsVuEt3LiP1bH/oqby8JlNI0fZu0jmmNQZZj6kzMbiaM+NWMjjyY
YkqfXmYV6QTdgkbyUOdaJWbrnwU85eIqkWw9n+A6EzQkhbFtraSQ5T3U0cX0qFBd
J4Ze7ManNyvG70/PSdE0YXD7eoeRBazDceXvbMQjb6C3lMYfXNHmSWlD4kqtQpjN
Jew8TzrmP51U4kS3oD88dGSyO9QNW13a8o7t+eBHA1/pDbJMHpAk4V5gTnYkLeHL
+Ea2QFc+rom22ZpKcZTkS3+f6SuIBrqQzSrAbcS3MLZfnw+aiRizeg283lk9DTy5
GdioYEoCk9athg+VmA7Tn/JWO2IVvyk/9rrzbbF+YOOvQwzcgMgTL827eeHqTn+O
upRURt1ElT7GMxeEeznkoQdB0/uJDba3DnGKYU3pYT2Fv/d1ivAT/VZEY84pgrqf
XD+r7YqrljX27ua8ROcMeOIybadHlxZaHsy1wdRujE6gGVh+z3t1gQLogLXoUt1P
w/ZcmDIVA3/StVEn80tAAsOXofPkNXUMHFQChItKqmhANw/5pxmQqzjR2hbbN2pV
B68gCZhZnsmrpEsMzfVR2N3fOK2T8z7/oSPGPkLuLVktrhTW4BIvjvegrbPUud35
nL1hS70GqPnoApUKv/BHfeJf/ycOOURd71uq0mAPyZUACFgE4maXCNHE94i9sgT6
58pwEsYjCckoKnqyVKZ+ws2R61jceCF7xLq8uOTrn+NW6VvP4gfeH5LH7V+PK834
G4cutJ4afOKRIScAOh3EbV9Tnjk0NLbvqaTQ+d9dfFrXfS4SlCRJNVC5SFyGezD+
gXUD79pOQpD4ntqI8WNJyICNWvWAhBu98M4yHELD8WwNgver1bH6//1loG4Q4x+A
I9Zw36MS2l881EasXjZjc8HfFNs+76L1nAS3wcIXvlA6sqgTWfFBQrVO0Jsxerdg
7vCUPGGrN/mAB4e+yCNKeDXXcsYVnHrHa5xqdUApDdwA4pS6Qyf1bhSvn1od3O6Q
DSRiACKEoKLQxoKdr7iOBDDvtdJck8nGCPhtRlenSGsxWbMV7MBHGw5+wA3ZKzuO
sMO51II+lgKQApT1CmQwou6FLLtJY4Bsh7hez8QB/+QqYPvlII6Njy5LIC1NVQsy
jyx3Jb+R4IzO+toaxP3Ur9LsillgexyjosbtRhJX7wj89muQwdNAQtSryPKlS99N
sjgGcJ0L+BVk7zeEQDH1BAlaDEM0pzVY62M1P2U8sHDLA9/ONbFFIwGFtKHXmudS
nhVZW/B/jOFKLqx9i0A6WIkPbHptroyoNWoFFR7xxwo03eJQFcndFABmLjPecUWz
FKeB9Si7HOOtc81tYhE9THXAFmUjbvGzi2O+x+a8Juuy+bNxRkxhJr29Fencbzdk
0jfzbB97G0Lt3DaRQkUVoaJ5lHqnwgKJ/FYR8a7aw67oUQt3naZrizUywHofa0zd
WlnnEpGRj2l293F7+IhyvTX7ds35QJCq4KexhFZuBxkMZASJRExBH+E0rYfX1rb4
Vs5hRIYK32OmtQPtQLcbI3fbce1d0ZP39do2VZ1Vv6APJypyCDb41iwMa0XXqN1Y
UJaTdgXovUYQvkuoNsYpu4AZYQt5KyfuPWZ3DUhtFN+oI4jSm8tqGiaMVhNXQwAm
EV2aQLvDshSFpJuAebONXpl+WvA9qkB1hDCkcDMAJ2NIOryUsdpHe4jhlSlVDSEF
BsZDxx8ok9lxH45bheh97VAhzoes6rCDkpPoa3hDbVGdJ6tzvLup5Ji0uFd8DrUK
2Yn/DDLkuJ3R6hDDxqGBlbW+9L1TyBI/vBst4cFvtir/qyCIbwFyrx5qUk3Mya8/
SaUxQrBvmjyXZ5J2S1U6IbnN8NET6VaQ7pAQ27Ofz7uGTxlg4bi2nmkd9Tnt94ip
EGh2N3teH771J66kVHfIF+XxPGh6os6By16EMl3YNiz/ikwwgEUX36tT8yKgRYBq
7EbSjEQXgYUD8yXPuEvHaPc1wvkFhIaCyS2KzIbSqIr0QNm6RgkejL4KdkIWr0/Y
g4yb4arEdAljttORjO0YANPZ/fzqpou/W2KaeTE8vH8xXPTMx3Ypj1KTqyU9AqLc
iyuofBJ/F+fEduKj2fWV9MLvzZeI8dHPB8WNeYAz2PDguXswxTKxXU3klJgl1hHn
i3iUICDI8OW4sc8STspL/Fzz6rainpW31kUGPKe7WCoXD5ROy4iVXz7sp74ZBiu6
SpFjEabSa9dREOZZx+CGNpVfA2IfuUeqkIpfK5PWgUYWYa5afyYuYXl5WlL2WrA5
h+ahBuLAVT33BHAvgnyyypBp/BosbOOztynwO2lxQ2lF+06Ns0QfPIsP5C+q5+0W
skqxSn4DTmf5wyxwIhnLHUIDDMbCgeEodkDl6n1miocPH1tGUguvm4iDeAYZMCic
0akaRJ/QVMzyPkEzdWt59nz0xKkd2Q/hv913tJPeMsYz+mDoFjM6h2FNavvwLnnt
D/9SFgrLlZlHJw1WuoIqp2EPM9232kXdbr9Kr3oBIwmuB9L8/V5u4NnaSG7Kc7Bi
mTTWpZAad+KM0Meijuo0zn5Cht9RwCaWD8O49vEIQek+5czq6UegrjFYYu7bB2kI
YBjkeVCd3FDywdexXGLb85YVnn6Ll1+FIddTD37SfphGb+MGoQUa8Ca+jkBFMZEF
6TnX6SdgYh030vm+dUlVhkHJRzdM9zMTNkVnPgQcIQbxVWIqkUfTmRFfOrF5TfQZ
eccDzQurBA64URjm6VznC7dqA+U91quARxA+A1r5bZ+djG98/D6wziU4BvTIyJTp
iZZw8756/4ppj6rBfC7E2lWJItz8Db2TOc0GKWvFddeOssIq7P/bwEI8PluiK1Qa
bx88R0HmDp3CjvSs2kjXLz2waNg293MHeGQV6T5Hpglv+6U/9aNaUHV2yxPYwrNW
ME1rjdEVUjEn7RA7xVxHmGtxcLiMk9hDfVmqpaX3BVvCoXvAGDJc7R7wtKZFHL3g
lHMJ/sJG1mXuFmz3Fx8EdIYBgjw/EwqdULBSKzOZYulmrVYDhTUJA7pOIgiCHeGY
Scobh7F4C1PLHUoxX+ohml9vGqFrQWKoLhHfb7L2ic/Vn7xXgs950KXsi8pkQGAB
/kDRilPjzZH0Kn9zpe6M6bzuYN+Gh9ZrZwuzVBY2726Z9Zsx0Vilyl/qC3ZCxW0W
8i6Bwl23gaMXW4+ac94A7+tkOeLIlmLlOkdgbx93pUgF4feTMVX7Lse8nTYUFUW/
0WSQf23G1ZQqYik/S5jcUqg4ooypjyn4qx3+qLYJ7sxeeNixjXs02mOlslWZjj5j
OkH9Zg0jCvs4uDikAPte3IlroxUi3gDCFQ9AY+NaVCg1L9i+ogzpaB2/BWMl0G4Y
TCTMKwp6UxjVqcxc7yDmefv//nq9lg1Ow7EcphLWb1l95IYV0Nq48iD1Eh2A4eea
CHNfEZrxdowMvClGZC+lezahIZu5/2+2O4gCr5Lgb3k6qJhsNxY1tHW3dehHnT04
QQkOvX2Q4/sUoUzlCg0yCg/H2AUjJwmpkBR2ozX7jyrj2B8KnQ+dKqE3hDfwrWaD
0XQ3nDnPNxc0cIhYC9M7k2E0F0FZQ1oisIL9SnNC8RD/TDZzKMc4Gne0rThdgDHU
foOLT2aPGmEQ9lwM2nxBo/sq4ZNxS7lvY3XGWx5e8EDxdWNUHuFqlENn/ocLH8I1
bWYOrnkD/xNjI52628J/8mffeWUSYz2dGXkkgZAYlHQravS4cigr98lXACMHssRe
lawV6DnM33NM6pmlS3GhVB8MxQ4Kbthrg5zKFl5SZTcXylU9pdU/FFB7AxqEr/bG
B/N0+e2U+7fbUw8PLuXIco8Yuv9zXCfJpKLaSg0WXIRKr6VcWv4hdyuiOqygeWCH
dtx0GE3cmnInvn2Rc4K22H9q/wiOZ6ujigpXjaMMBvTRcipLdEHBQGIyT7SWcTUi
XcEtNr2x0R03hFhLQT7GJFlRF6tl/fXGoYkkp+vhvbut0+ZalXYs/KrUcIMHojWN
Jh9W3bkfC0au4SkTbNCIfUQ9/b1ZiBfhltoHPjUwrMZW4HxYKIjdjfuIxeP30Clu
Ut/bzfKaQGBQxD8UWBDpnECuflAlAnhfYCYHFI3XI2DNnLUK45IwrqyfNYmboFYZ
0uXWR3KNuPXYeD0A20tjON5OB+/sDNl6oDPUtVsOHOvteoWaB9ANBVRfChtfJrRs
Yxs0qFg04o59xrSKdFhaJYAVYE5B+66DNwebUGEshYUeZKPN5ehJwemYWKUIyq0X
Tv8JJrWEg+ikwd5DtkwkCHjzYhairmmTw+zDusMPjR8fy5E6RaZ8kuawUtOB0HCK
peQjHXqJ0OhzQ9KI5nW/7PKqCtodXaSWDv07mTmGF0gG2jiqWKWlqtI864LSk9El
5ND0z/Gl6DKQhDfK6UpO7a7ADrnQicy4XwwhhTZ2ANNtbfjDA0oBghtEvmcm3txm
6oSgZ+Olba5ultRAJ/k84A73o6NRkEYwr7e+Q1ybU49iZIutGRfJaT8QinZQSQGD
fRto/2ZL6Jz4Lswru1sIEBrgKu227AlNL/XmAVSRGvVMjawujOvNbdP8ABSnWovc
Cc+0pFvN5hNfmd7+gSuux0Hs/ywQoIsni9w+wJKbZr9VlATCeugh9QgThkfyctuL
FVe3WgFnhys3aUJkI6Y0IRJZCh/jwFrIxTr3TkJNWUoSxNHpv15ZMigvJkMBqDCq
nTvxjE3ljz1ljUhKZvCbtt5xTt8o+iikTuCAbns9ndiT9nQhNjb7+EPiDh+3pTy3
emcGCepmqGOTpt2+eNT/v3zoEYOjGH/aMrM7kN6ycdW458KinOBjb3uTJuRT2EIG
o8YrluBAkTxEVRrxIpx4efp3wkMd3eWrl0WVudSHmeE7ZPW3pQFpK61L2POy8iVs
wtHlcd/Y5KQUP24bKmshS9kCbnMAwkvGKxx29THnxGyEIv9fPvEiXGqvUoktIrzc
KVRPedgQpC5cBXx03psV2v855ZJ45LBmeLno8oXkc/K2PCFos+d0zLMnZ7DoCpMW
IRIDVvgfJgrpLF5W9BFIXu9O8xdJgYfG0Cdi4RNj3hIne5JdjyIT6fycdkbWmDYb
ug92mWPLO7Ntl1Ccb51X2SDmB6HDlsXld2ufsdnexv8WvuWrlTUuB3aClCpmUSQ1
RNFptIlMkkYY32Z7X8jEgNOxELrPL2kyu1WzlD+3qnOlsJr0VZXoinYsHU01gimJ
KDen6igiA7H3pEd4nMX/Mb+Z2Ie7lh8Sy6acmYTy6wD/JurMeqvuDVBXI25az71i
pGM9yL+O6GmBhC+/NfETZHxmERQoFwY7MYf53hxqOAZ5RzSrIQ0f8FXPdTk9eZ44
8kgromC8JanFV7IfqFhf2NyKdsfZ5LMVwmpqKRvhyC0auvbY4wpewQ11Q7Uvbdtf
a5WL8mWtYl4B0m+ukKWuTus9D+2UgxSx30aSK82EFQk+hW8BYOd7L2Semdmb8Pmk
YkanUeRZuV/aggo11vsxWP+COrKDg4FEXIRzw4Ioyf2Xh109kcVdKXnkxpH+hXKI
oUCComCTX17bzUpPu3UOi0EjliAznP9C+ZkbULjcngjvz873m2Ps/YYrzDMxMBNp
hvkhS8oFCYChS5K+93YVJ2iXSA0G6RlO0CVKjH/LoqTnvdwgjSROIWQnRVbcVV3a
RWFi7PWiySAhKc4fRxgcV2t+R3FWY/VfLvt/OL7CfNX0q9g+Ar1wjLit0wc/wlA2
1PPSwsPQz2MHamxA7IlWNuOiyicPdvDK/5+M82xb2rllO9l8Pz4dzH/yIGajDWYc
oyKB4MNwXJSKOeyRBqEfWxvJMHvsG1ik6du12FCauRicgZZJafyJ3feqTnp7dEsS
v12oWx/FNq4gY71i67QXl33BChmJLx0ckx1q68tKJ4XJHoWTt+zB9fTHFi4aTUC4
mxW9uPZ29x02IZEHjqPErJn3dOAd4w6SsM31ioIzA4FG96/gp7skc9BuMaH5GQLA
KEixiOJAvCjLjRVqIcDgftlrxnH0/oXWR+rxYX+1r5jkk0yP+SPSfmxh+iDOiGyz
STti/FGh6B1cY7a0+r8PqY9j62Zk16aEPgrJ7osexfPJ8bh9/2DcTbAjeI8kaOhk
xZSMaP4yDjgC8fPtqgtRJ7iP/tBGkHmzwyQ8nz33Dq50fXMfoRYQWfCBXCje1Uyk
2huIYnkUWeSp8083k2S6Iq/wFGv7UhOIAnrMZhDOwfG5yyqxe3JaOlRGvybnEK+c
Sg8ETJCkWJuUOHH2PIn+3FB9IB+IpCwihxR116wNypihNBg60bXSLCKfaC7MzG2u
vyG0Hur57JSsU7Eqb6YtyLl7k9bu9h+jkCZQjUbkp+H4dIjT1rTZpasDEM2Kkd6m
D6keAmXk9N8cCXpDlY1mTv5TXBC42FqcOaa7FQHwwX28oTDpLWGuDPaM6Q25Jj3+
WRjR9jhslcbP/eieLpttL0UbS9bNW5dFIwODlW8+GSLN9epl0wxWSolIgWho+0K5
Dj7t62fVshElnsLsaknyWDVc4oUrCRrYcmInZlDQmg095AFN11L+E6obkmrFcbak
Ixapet5uDpQRA2K+GSQQN+1fk7sCqcy61g9S/wDS/8jyeZ63ptejf/Zvkx+ql5iR
P+CopMQJeGTCI0KjByvdutgiKhc1a6vMCA6P82cBkk+CKW2/frmXJdnR3W+n8qCp
WdihiQNW+FCz9J1j2/JAMcAoHMMMQxowM0irEnKmYnOIFvzq7eRYjZQVkYRnrpEr
/MH+X+4AS6jtxpBGB5/xyo1DZhXy0MVSckb1PzsR+re0FMF3uvE/jr9Q8WL+HaJl
A76tne6QeM9e68xIeei9xX4YQE0jEbDpfHxyrn5pMBBXXkn+sFdYWq7PRmJUK9Zo
Eww39XDpKV3xW8vMcCz9BKi7a/LUlTlEVC8oZsvTCiL34P56j9Ezdm9XSKCTRlgc
c/30Mc0frHo83Surs6CA8TwJ9oMfjnMv4NHqme/o9ZyyfkRIU79/yy/rxvVnd0F1
NdnT1hjvOooI6aF6J6PlbF3pa2jOJ0m2IQotG5L+HrttbIofqJLQp/Wkv+vaFgaQ
brllHSC/z699HD2ZMvcwkCzlRD/z5f8pkjRroKTlT/nLur+Y0kLmp0spTjAwpWNF
D5XnuVzvQwK2AHb9InMwWv07gGlyTq01XKj2gvlnjj0OEoE+Ba4tXjM73VdcYAj+
3nsH7l5CEsFsefCOYLdwlxt7uLzdzJT2LnxwASGphrWwaAlo1oxAES2ET4eTre0/
inKG89smzyRFoI+33bsJvEgUZcQ6dsNcawoNAuXbicdYVdn7zPFtvom6qoLpEOqu
QeUUQD15g85jlX6w406Yy3U5WXd3ikc2x6ft5Su4UPNo7HNLqcAnr3lDFDQxghXg
u+m2naDFPW0OVamAo7jaCy0wQskCKB98yhrpQHj4FM56PMDgDfQbJpfunzkp2l4/
B1YgLKHhIkDvAfLcshXbP4d1LqOfzZS4J/ep8lsvJNpOuXxRsFQNHZ/OQu3iZLJ5
Ct0l/JxP8+t0arEwupweLka9zsd+K0wyIBRlfPdtDUIZMjD//xmSHjcZGuRdUVZm
t2H1TeXmmLRHjuvnH68R4yMb6Ewfd2H1Trzeb/btEDIz5wh7Cu4egYuyETepSXFE
687gju20dw2sv/gEdj70Zw1ADBDJx1LSOhunDh7cF5YiJTqDHI2fETL4GsDICyg0
K/Cs/6llk4UZ/LGsJXxZGP4IzmrvOwBdJQzGz8mWBcZ8g11kYTgkw2vmbfeiobO/
CQCI0tHe5I8B+sUVt7k3Dp/dHqWo2A1exZDjrUGO9VwVezrM98+XQL9iLOjlfT0S
cfBy4kREoicMaHo0fnIzicwXlZqY8nMV/kMGf/1XX9gnvQO1umZ5uflbeFKXj75/
GAGH+P8dTYraGrJCfRfxwCIbfk8si5vPqJwsmOCw9Us/9RO+ofTOVMyscQVVLVv1
igHMmx0563Xy9woSP5KE/QgzAdZZRTXRTZgyxkad5DqWPjOLr8ddUxSXa5AjxStC
mzF/kXefRxGr3qwpNlokl4WVFDedqtnjBunwexsbF8rlaJSJKwg0IncijEwsLHJL
lWoGfD5HauFiPqPZW5jxsB9kZU5FYIgP6lkOtDRss9EI6rIhuSZA45Ose+GZnRjX
F0r7sxVD+brC8RwPxDRdW8jAWt7l4HFy2B2nDNhOXLXLL9+ChgVsWBkGRv687Rvf
8r8jYfff/9FBIENefVddWp9FCMvKCqbGJfuyQLZWIHeajSOPu2X1Qv1w1s1Z6ssB
aQ+Bq5BzB0uZLLRgArmyC/CX0vSFLnKvQs/NCxv7cRltVu2saeoHChoPmvU5/b+H
PFZo57RUT6+4FopfoOIM8oy4HgSAgMQR7+qbqSnLv8miB582MDx+O73SAWMTs47k
LyMxQtEoYIiwkjvv+QqHvFHp/a3Y1ttkfMRn6QyJYxoqSzMZB1mDzdfpindIohHw
EISdULarotEGtam6zr9zZ0H5HbgDh/tZaXIG/41qx5j2WE/l2xJ2FfNqiuUG9xd0
NJuQKc5uwgKsP1qAtZgi8g5pTQybh1EXW6WX7VBCM8ZK/3MPufML3SAQypMaamqR
xlgfmc4B13g1SxcamLA3d9OCKPoq3UvoeAU3BkWb2kYUoTlgfrA7NTKcvuW3mK0m
CXU/K+hWo3sXDOvhIdLgRtJ0Mrd0YGQ2wSD564AgsHFzRvtVHZoae44X6Hjf65X7
xKTu35iVQlfgi65pgnQkPV35mR79GQ0Qa030iXI6Kqc6a4Fxt4rJASix3wLuok0Z
mEI1zq9EJj8WjswCSp99iwdkH2RVHB0QoiKcIy+cL01xBUPq9xb6AyLrDy0HsK/U
hdFBb5kxS+hL/zfznGCYYBZBHBarYwTeErztAZk+Li4IEyA3bv4+p/+UBY+7twYF
hCqzrMLJ68VFtiuydc94p74KBncGqH460a12Wj9QDZdBWVSFPxkueUc5LmRA9BDk
wWo80wG8Y3vdNW86Ljh1hSmCNn+1XEBVV+2CxxJsCsDVAgCB1g7xACYHwmB9wi+P
ihexkWsWePilkVTVo4zTk7tj0JLVJrZS6qr+fSq9GGTMN+noXAp3QwnWvLrRKsWw
sqMRBUc+2DZLJ6fnRwhtcNoEzFJ+1ZsTVvW3s5j+1mS2lHvhypsKGls04TyGxCdk
hTpaMZbLbwg3nwqbtQayc5QAWkGuqHzVjdYFIVnXM+QpiBbFsVkPYM82trmbkm1+
hgRrprI0c3sGQipTY2OqBoa8nxr/Xpg1/10wqnIRjHz1DpzqYMbg/8nlGfPIN3kl
3qWYtOt7ZwSSbXQRHLW6O4ANSefwEC7U8vKImY/Fa9m85cDLhT+5Dy77io9idPYZ
G+uuJmzSCaBjpTWpZbbmYZcm8Tx7s2fPGwVYKbf4rg3awy/qguT1+3Y0VX/3oKrM
Qp/2Oet8qPgds7LjCoAmt8EfFiVYxZE4lHtOUQ71SYYNy1hE5c979CwiI37C1Y/i
pKJ5vTrbIaBxJBCGL8k+qCPqx2lJFhhluipx6RYia0AMI+SHN235NAUrivDHPW6b
f7WWkjlBHDVDtF3MTiH71wt14beLbPjwd4q6nya+dfQMjCKrp9HAIMWAZkCvw0gG
Fk/FcG3qstMD975QaMGy+1nnjf3MVF0y8qOtMm+zRg22YG8DeZyp90ChfytLFcu+
qbpyOyrGhTT+jl/OSUxyOBX/AbTGfGPwFgrGSrr2qZhLMbw7csq0RVTEeWsfkti1
+Jgb/vNCv06RtHhezrd8nXVZ8QMnFyyo+SzxwrF8IxJahzXJ2skhbAOh3/unK7kc
nQichoc+kmFHiAf5NK5UMRUrnorUhok40hUOUZl0OAJ6vWjn+7X+KBCTlObNistE
MBFJgyV+0HEW6pHYkPfRrUc8346JvnGZE+jjT56ZAfI8ICmBzycP46grWD+QSQzI
cpl/XVcmoi+R/dQdwd/E6zndignBlmdUxVIFk5pLsGohvlbFdmY234+9Rk2P1JEO
JROlSLPStzgrElo+m4uMTG9+beQS9qsvHHm5NZhHqNRoxd8pdqltHwRZlTZ+Rtxq
6OH0ej6cbRLmJ1h3nqRUAEvNc6+L4DO94QqqT75dZuT3inD/sNoCKvf9u63VaEiu
sUBEbtY8TGbLpNbBwoMOmpijM72hOwgONQvP2C2CQMBHjXnQk4MvuxVL1ZWy3sA1
SQwshUZxE61X/f6SKjAlCILyZZg11+EJBmzbvXNEz0phDWFBRwa294vJY4teVZR6
nTbHs7JiliUvAMA7s4EVVZg030MXwJZg9ZCnkatSADK+iDVhKJK9EGqk7HkIcMcM
codQ6bDDHW2zrOcPC0NUfXP5hf3ifJw+Xcogg3Aux86fPNVGLoGI2ER1qcgESSBb
j6iqTNCkufwGOK86A1MlA3zARHqXUNoBsqLZd1kOmYRerFQIxMlNNlOjnI9u2vhp
Qd0jLrfXbCK2uTS9Ey1MKY+XhvsIUzT2BGHBCYgEeOVvhFR5Ui+DsNs6fcvCS0mr
naeozTrTj4Ip5KGGbpM+JdF5ZrbiHlsY7OJSnbwAzQiIZNqy5tM0llWno6NNoxeS
j4O0YQgDawwHh9aSFCGtyJ9C6o9L4bmVsVSTN5i/agXqo4Ftezw8RT/BPGaHgtmK
iRk5h+RWGMpt5J6N2m9DmTRSBE444bP+6EOic6XiCBVrqlQK0NC4TatBiQKQi13Z
Q8FPCoUw2lO8ehC5uqApTo87zQDDp9N97ey3ypLDTZpzUfKMupCd9NVzJ3bCqM98
LU/UJhRBtfNM2M/PUSqINcYy50WggePb1tClxeejT0qNbn+kM+ES13R6waf1+Z6j
KaoFqmSbIf+JC+R+2H24vB4fO1GGmN1Eadbcgp/KtIWgTgNcmRXoqqeLIx/o1DNi
flNrbr1Sgub/AlFN/tp+yLLerHDGgHFWkfFBdRt5B6L3LtocpTLnVWKj6KSgd9Yg
5Hx9s2tXzLx0TeZGi7cPsIXFHvM/+43To14sA4otYBnT+6k13EfaHY/hDjWOOm+f
BoGLHm+s+N+ru6///Q1ADgIVdgRttXpPdl+69PuoYj0r4k4v+hiWXbfVZ9p9kNNd
jlTwyafA61Nx/GfqjJbunKwJe9KTSiCV32eWvGFkGFkyJwbBvEvPcxwtmWzD4vbI
q0wH6QHUbZU84L0VP+iu2gyQMeo6zugYEmtnrCBI8TAXFvP3apV02PG+tfaSzfCs
86fQKXoYaJJ04KGA12aYpF5SVS0ZtO37VkyZf0v6PCCr4Hmku8iVUNKhopGGyi4f
GvA2bcmdBj/MnzMrtT6yPcv6rULcOMbZZH20MkOYofP5SfWHP8HZE7ws9MtQTkey
m8r9oPlLjYUC9gUCNfbU2TbaR9+ARF/4cayNTsgvFljumfKqHcYZxLCuen2TQEnl
6q1a4xQfM+hZrEmStGDJXh27jT/VlpRZwL1ykk8/Xd0q3/irAkKoBOGMv78U6TRw
ILkeZqXNbQg/4OPQMzljJsWeC6pxS/MMO8CXWCVHDmqFIIMO8cP6pJXmCWeYmqwb
JFhpS7sg7yb44dIvb/lSzcjTBenYGDmErKZTEjmhfjlhE3zoOFr4KlRB7pMpBEoq
oaAyrhKpvuWthu0Xycpi3TxHd7Ggc20DyLnJzePY3JvM1ZnwnPhMOmJ/K4NtHE99
tjRM0tKRbMgCiDz8z7tsNEp2i3ohH3KhyMR53tgpfYdfDpd0y7YSajw0FU7xuaBZ
Ax3aunIhVrvO9lGa5dCk4vDSyefUoPEAAyaVcU5ZTJKdIHC0lo8SPygE9pKaliEq
NdASsDQyRTcw5foZXsLLOJxhCTqhsoAtiGgrYjeJO9RPCgZVEsvyhx6Fpd53sNYn
pGoUljvSZzA58BQSHA1EmAFSs0waG3+5hNoVUUP7g/3x8r/3UflKNB0ryJ5bCP2P
xYrFnfpt6N5PE9ei5FF6OatUGeIzutjlJDe+uSO9HcUsu+jN4wPUi6i8Abk6+eK4
siwAWvaEEZ4hOpsPEJ23kU1HRwy5ImgW1ny/9jtTDXlxx570nRiW8Gd1+LqX/Kfu
i2FOwr/ZPnlMGyj66yuP7BpbKwllBLBAyrRjSNfqyw9WFcy+h9RymEzS45MhgTFo
nJGlabSwf6C1O0YS3elIRA/4gnIYilwOLpnjWfAOzQFiR5sADsjOfS2qiQb9hD1J
69yklvUY1YMAJvTfHaSRD7LeE1d/9KUQvrkSm6yw5laT3lLhXWxX4Idyj8Quq+2E
7lcbmTZNzXr+zqFFFkrCmKxGm73Zi+S0F7unMSgsK83LcEOikDQeoM9SrUrx3+m+
7Apo0UQ9Zf2ze+XyVWVvhEduDo15IMWMXat2Luti0SwE5Ye2LskFAyZxhQnUPOQY
MsGHNgQG4Gi87Mwt9h8uDOfTX9vJQN6ged0xnhmGpDhN0EU5OQz0eg01HWujecvT
Y5eRWRjqCEFv20UVT1yn++sYir7P+SMnmSGupp1MEZF95IxjGXvrlT/4Ltl68UWW
OFBDvmmjyZ0S3rKyYfF8gqdCq8Eh0HaX7aRxJSVUp2+TPYCxOLI5wOjl2b5VB4fn
OdniR6qDe4Kti5UB8RYZb5arvY2ggryNj2Pd8MWqiAXUaNH5cHkRXs2Mh48Weham
MKqaiy9+XF1bO4RDD0m6Q1sLtfBk89IG0/GjPE0IpK/NE+7jXqQS5GV2a/Za0qa1
BWWhDLlsjGTiXTID3rdlJZ5JpCw8GzmDKbXLvxdoj5dVFRTztp/wbJ3LG3k6yz8R
D2D62upfryH3P9TKEU9j7wFZHRSTS7NP0cDjvFGoZfsYhTk1GzxwmOaCXJNtCq7P
RHC1Z5IoGH2E5o/rWo7Fbvex22XvR1E4IYM3oKEZV4opoUEJdb/RNJFBG+MElTxr
hcuyZ3j3cPB0TvxKKlM1HEBmW/tu0iLJNtUDtp9gC3XRXFgRyrzeFa8V0wBMLtfr
u1aPag7McEp7WSNl02Z1UhFKnQ7z8BgeFE6By6HyMNs79cViK5bfn6egw/f8c560
7fQtrbyeF2IwUSR5WIEKu05949xWTyHDMUgY+KGtV9t9Y0PTIR2DOim1YawzXPVB
moBvLvgoWuohWE3fkduNxoloq4ZCsIw4cOOYeC1htFrXk8hQBDwCWqQ5qEhB6uJB
zYLmjTf+cArAjNLDMNpXrxzMBy4rsj23vqQF9Sd9QVvO3QoDQZsWgw49XBtZHo+H
XQHTtrvIJKdVTxyOgBattXAS6z1vewymMyn2dntK109feVrHU7htbn9KrKYur5C4
XGE5Isw9qBas5oI2WQdzEA8yKQHwZhCC/0INB6m3f3jI8ocrNjvHfg93PgAC8mZD
01sLECMJF8WYoIX4UWECtKRGXE/7lqq0I2feLwiCD3MLSqh+OiDOjSH1UhQsCsky
TojdZ9RJqrtqwUGHCgOeN3bqZCSVDvf3JwG1cFruNE1teggRzwAgW9/BOjQfDaow
bsD3EsbHhturTdnyoAM/w37Qm6FtfeDLV1bmiGf2E2+eZxuVIagzwffNDqRwXdYl
GrY9fllISJ3GfqNJ59PcBFLDgIO6yp/AlizbNODDD2cah/fgU75wu5n/2NwWIy7y
RTjsJ/QvgmL7F0LDw427rVwcW71F14hbtEhxUfAowVwhQ7lmIrtRWDRv449KhvxF
86AHVDHGGXv/+MIKTdLxxwpSvKT6l7CY5o/GUVTzZ2832uO3o3KekCKaBErytcGC
eovGLIGiTzuVCI6y0Wg9LUUl1DPTjthdpQ/27fYE1zjKA1H32emCSAjLb8eFmkcg
vxjxqoLBkhihqjptSoz0ZGrhdkWxlEtwKItC+WZ7PHeSdlRJWfFnDj2YRyQ8UWOt
BjwluDAYSWvzSYD6N31lpD4cgw4uZuSuClDCkQpVKbPRbQPOzoAoBwtLsE3T037V
EVYKi/ATYyGIaA2jSwdRBiBw6rDuqiMDaM5zJD1DPqIVg/XBR78q3xYVZCe7FcyO
/EXa7x8wHZuOxl6IknPQ0z3HRcidEI4Hlg7tGYcpijh16xckKzDI9XnWC+ABH/yq
hEbqBRSHUjPFlrYscm0rXfmAssjpAmpyV14n1HUvMbZ/9Vy5K5dZWfgmA1s/xub9
Vkfg8BYIO90kLXqD1q5QZc8O6JMIZggQsp8j0AqW9dWSgjbbezHgASSQexSQC4dY
Sutdm6IA0XH+uH1pn29nKXD83njuv+Ys/DIr/GP4yB1/0lOAhA8pWSIE6uQ0IO8h
SXRp4R9AjYQXdTMKpMzcsnZPWZ6RilnqHLtq857FZrQXMI5i8xUhxcEhe423U33+
CRsHbvVv/AhxOv9jvsrTJT484Yqkjyl7Edyj17AsT+Z7OnUvNsppqgRFb9wAZ3UW
QRPsGIftBi2/S1yGm6j3kLPXlTNFlYv3XlApOacWS+lmNPbWZUnrzdAuTD54lZU7
HWIDupNzgSlAl45GaXhKg0ziI+3gDAd+r0Ri7vaQAFGjcLtdTE1ZVXnxBotQY9fc
LXXY+h84pGWPogIZ6bLtrB/eygbFmaAp7TBe2MFcC99Ndcslbh6VslWpmNtSVmOl
bxTpkPSTyUSVD3jPkLx4Q7rYuoMYZgLY1sUP1XyFMdls+hE1SJR7hem/e7LUdxOk
cVif4AaPkKnIF3xvzg5ynU8u2wjq4oiRrkqeXqNczPTa9V0Rxgu43a45hL0jbLuz
IMxrlYPuD51BACtQQI/DQ+uywdu6hcqfJ+BRNYQliCXuHwcM9+T291L8psCgDfzB
9koLRXwnNwgw7Zy3RPxPtxKhT5mjPofhEEiIKiPjhWHLUFQpo4Ygee8dTeT9z2Gb
L0f9ZATEFCF32EV25FP1opcjWa71GZ09veittdDtH1YxALK+STEB0LkP2CFJMmfG
nQHvegLF1qKk1nzpV+8xPkwpefHT9zktzpSkglgcGrwHGIziUnGruwrWjuGMFTFk
XwG7JjZDytIVzSAygiqPIgG9qz1rdwaDW15QYmcR+uPM7OZXRPVdudMiqloWv/QH
lUEhETu3R4n970XzQ7+VRLX10eVE/1hoRQImoPquD5mX6Cx3KKOWO48Qtpb38WzJ
E1Hh7lMdYdQEuOJl0IItWTxuZKWuQBYyLSEMWW6CoyIpctELuiu2XfJg1HKKYBYG
uKp/Xx1+1XLTg+rlncgwOCadvN3u3VoVqOUh367YZP5yF5cjlH3pZYnmf/G++J5k
qwvrCVH9AaQLA92+FK1SrPWFfZCgXkz6oU7WiZ8W+G7P7fZRCxAtuohKjVzeO7pq
r1EsjPeR6QU2a6RnUYophVGAdQJ89fAiYCRadW45zo1gukFxQMPD0vbTcIwh7s5X
7Pjz95mBqV/1JCUJmIH41WPLbMVCgWwvUqR/oaUo9qrHxFvgRnUXed7YuEls4a8A
4sBFHIzmreioZf/W0VcKROt3ViNLFVr79elYo+JqpkKGhrnMe/2fYscINzbzjT0m
WB0uqkRi6lltjI/laRc+4XUZ1KTQ1GfOLI2XVp7UVbHSb8tfeP+qXEQUBDmnOjVX
F2k//aYWyINs4ewsIkHOlNP39JehuXf8JiWp/gWxXZjazXEA/7zCbLTmJGI3mQzX
/62TMytPo6C+4LrZvR0Du1IIbJ6A3ESIiGmuM527jbjYM62ENF+KXxG3uOb7eu4C
gFGD/hIWPNMqP6f+yi09+dj7j40+i0dNbtWdbHxOnnh2kPZvk2CSsR+PwTLVCXH9
7BdHx/za7knqTHrDQ2g25Kv54SsSOiDhYed7ZwLi9oVX3q47pGZv83D62Tth6StP
UqvIZzvs2QAm0sJHmV+ahbYK92PWvMfRMf2tUk55FxmOHypzxCYcX65hUWleOtZz
Z2dQSTsy89LYhSvLufktCU16mJbEPF4nblUHNcUEpAZ5t5tLH6qlggP21w937HCk
SuJDgRgkDJUYY4u7rNKd+BhrOTWdMLQ51pYQ13fc5kAEESB2UPix6EDLD9M6YnaK
CMR3fBHPX775npf0+k1CWz6zm+yPlqlH2e76Dn+LxqA8GJCdW9xJK9z1d8/TV0Pn
usHDOFetiUAR0GyZoSyz0v/6Nc7L89Ft3SjxjSGEtX/tglHbpkfY/j249rC+CFUp
2MCOi1NryTqViakme5KaWN2CcQLpLf1GVQewm5crq1PDumnGGizLuvY5gf7nbnI+
C7mKXHWoTNNzHFnKVdAxlj6civ9FOmmUIRb9wTUL/P66UnblqxD1XkpAjlio7JBP
OYwmAEWE1UmgdL1MHZXLxrR8wmxQYbzGy7jsqVZYhBjZDioU+xKBrFlfdWeen12X
7DeSqXzGJn1d5W+6WZkFWU/bJXkJ9sF2bOV0cPvWnvrwdR9BxbeHRSuKW0y/laBk
iM9AO6nvWG9jx9cbjQa2l2nmWhK5DeS5pbOuU6iJi1zKET3n+dTL2mm3HqlQrnwd
CKo5vq41JkBZvt4BJITYbfJNhtUM7wZbUEyTS1wlJxIDO9QgjMfTKjX9thbmyZEw
/2a5mw1sOzEDc6tik/f8wpIaO2LJHZuUoIsC5O8kyHS0ObtfOaDTaOn48uM1jSxq
k4SNP81gyF75xwnneHPgIFihTt/x2ae2SOS1Q6BK/HWW4pHVZOZg2/Oc3tLccmDn
ggWkywBUEvx2Ro6E1vca2GfHfBQSIRuQDsvxjD9OLnZSW0tBFim9y390d/vWbK64
CXhHIyxHhl5e1qXozne4JP0tGflICZ/lwmU71H2bD/b0IWomG72kWH/6FoGKjJZK
rSgz06JV0gN0nqv1SNxNCiVTlKwoQUWsbBBMsqy3rqMQy+Pn986PJbIVPzwZ85dp
eM281SrST3i18Ggfoqh/+XQxL2Pg2x+kdgarwaRfvZnf4/LOWym0v2VpX80Xfh3d
6ONnUwjfs9s874puq6+XPuIlnam2W9qHs6VGdKUxidpOgbG+RQB6QlFN9k52RFq5
ck0+H1WchxO/kODs4D6hWFru1WiegzHuG4FX7PZnO3EOvHZHdAcCoInB84Be4caN
j/s2r4zRORq0VvRzhEs62Wyxigzz34a4qBy2V1h15/ard9AFS17VcjP3QnbsxoKR
1YR2vLLwvXl0gwzyPWVJ06LxGDZCazr3Ns3esB7J1i7pqas/IVDVCkA3CLLS/uSa
p/ICGMnmNS0LKbubDW/IEa/MMkGX9vSRdhFjFDlCd22qeCIhbabHfsB04y4qyDsa
LSgGfR7e2dCBfb9c4VjbjA5hyjpBQ0w0hPp95sPOUVXKU1qz3UGLEPO28uP8e+o2
rGI/fxtWXPp9HXy5Jp0GwCIyt897MfX5Kv/E5ZThk+akq/JRRmwmluilKL57uC/I
S3CLzhh9bySVjTzrRlWsKkkklFqp6BWtk0bgo7yhBHkdT/IYGw49T3RgPJTkWBUT
kOvfdRrnV/8VPYo8t2oVTex4j5dSkkbgI3pl3cnZyRXfdwcVTlI7wtZAv39Ob4Yt
cTGSoSKSVxa+NE5CI0KGzaLp7q7ZZWKHBL7PHXwm3ImYYbvG2vfq+56fg3n/wHq4
KpvFfGCByvKuQYYSrmM3Lw2r9hH7iBJhMdY0qL1aLcC3ZLDG1k101tTKt5p9S5gl
8FSVUB7RzSyzrEsfoi59lA1GTOBhPOAgl7FiN3e6lM7kOuT6Ng+U8ygYjj00m1qU
WhM907/KOpy8kJJTP9co7++iofiQalyQ/pRiM8gre/NhK8d2Yw0e+0Z/drWPmA7R
pHZklDI2/jDqCiMJRmPt524CtLgX9+0Tv6SIw5FCSd4KbtbKfkqtPGjyRYk9uqu5
RMGYodefx7/QddmfOQon/n4Rrk3VUBzbl2uSlLLs62+sokhiIv91a9yOmteB6rVD
4rV8Hl+QYNu912MCfFQM+yEhWL6oTxNyeDg03u8ucvVEIU6gM/Uap9LfMTrgY66T
cS6YmhSK0s0BF8rd2vHdAlxXG0jdJhImmFrSfaeHwJVYKE1hQKpzWbkCYXErILWp
rzQNm1polU2iv9hbOnCeffiR9MqwQfL+Mf2xYmQ33r3WGeEvyHSBuUPLgSaTTNtE
qNCPBUkR9z3JNWQ/sv27mREClyM1WDQWPpK+a8WfPBe8StBm5p93qilRTeF3f0Ex
/nq6Udo5oxghHy+TOA03mP0tg7981bfHqsJSMIuVoPFVYoLUvtJV1MnBO6d07lcM
YX+9DpVAVYZ/92AaJiRjuPr2KBcWSpCzHR/CfViF1FJD9dwFgYQ1PfQiu5TqpS99
uwjaesEGRiXTqXwMMEonxKpUlI73kxfJ2QFcuy3sZBpMXppCvnL+Kl9NrqqFJmVa
XbFE8aAl7sdvJuOCS6p/uJeVW+knH81sHeZLjych0LhIqZ+KAGGU/EF0cpWbO+k9
Gkdws1eufFltjVURMRC8eCCq+OzIohRl97pv7HYTyydnBjBRD1BLwhk1u1nNJjlZ
Ir7a6kacC/WUL+YUuuCH9Bu3oZL//mwUufqIMZRcGRTFC3E6BT2L3vSTrFbG48oN
s2bZmi5QRNoYy8TtsyF0QrwavOzfq0OAycRGo4VN12iPeQbn7wO+MM3dE1VdoyeA
VFp4kW01ir0EeQmeMr2JCXLRChwDgyM0w/vY7c2H4noILzem0yqfB+N8ul0UraWT
U5MKaFo2k/RmoTHI4Qh15JjlSV7tkk/YxhrtDdwcEBH6HkwLuw9bzwgNhkztgDAL
wPhq/3P5AjbMRSATlsJqFk1wX3XhTlk8SLvufiRkDWJ9J6n3iY6Orl/Jnh6/6xnw
2lHu/hGWejN/mLb005DeRb7gWEmCszePjNS7zu/QIX33DqqqPr0952PbkzBo95cD
ilzqcjTaYJTZl/zOZ2CQqkHmnE8t2/xOKMnlUlC4K+rRdfadtf++2LrVlgE1r8rL
vIok2ddnWn3m/mEdRW2HbFtgfcGz3kZeqH29/PcLPO0sTwqixLGP7QlnwB+vn5Ea
40mluan0zEhpGik4CEEH4Pdvzm/bdz/IAqD00N+HBNF8U/cOLVnvjPXPQsUp2LUP
KRnT3kLFCcqCFalmkDQtc82nLjaETEx1ejV3KqkrDFXqIQv643J4OMTWbywAHwye
Xtc2NEAgR2FUbE9zC6LjBbRpzM0uSCpF6/sFc+q+GD+dcAdfLL2Zs1/J1sEkoEX6
GNn9VCqj5pb20OkP4xCrydzzhn+LWWwRWEeEe7+2v2EJGnqBxW/6hW5pKVfbwnVp
k5Y9SSqYdZG107mDoZbGmpSwD7fhNoZyK8Q/vbSDz/aIutTxHyNyQYkonw2K0DDW
1P43cFXyRczGfEkk9QpOeYeAjR1DTeEYi4fRsJhdtHK6/9S3CtfSWgYfMJpqg3Ni
xXVTrkqALhpJho5ahxYWs/ejcPppVjpR5vl0GA3W/fP7oOKwpesMHJOa3naeNFvt
47+KkCquJq7c9cWUc9FbPK6fWfOyFcUNTambG+CEIPCqotEhPliAu0kExWAvAOIO
xDrbHEXy9NbwO2Y0V4PYuaSJYgI7kAXOehWFZ0/bJaJNXIVZuEmlboir+6YnCzAT
ivRk667uESa7mumx5qfJBpQV0ytpni/VipNNqrP0xXcorHb/BpthxJglHrEzDjlw
WPMgXvjF3bS5o4jFcdxTWYEkj65mUBG7oRFgWe8nSqQsEQ2Rjj2sx2gPmUXgHLqk
wHhcXlHhC9n9nlPb5Lnf/cb1l3hN5Dkj6AxWmyUjc9g/LuYRILmK7yfrvyZc7FT9
kNIVn3IAo/RDdTI8iZ+K+HLNNklMRIlgD6gT2qAh4x6uMelzwDhq861Gzv15Jmsn
YMkfykfsQXtqxrtd8jM+Fr+dK7G5gG5Vw/mHUPNAu/rLhfXCa4VOw4LZHMk2TuAk
+eiJVIKEBVDrMvrmqbHR8/Uz6qZ2Evv5rsFBn4zTr/ITB9F2PExa8/Uj7qj9A4No
Cfwylunpm4wN8sofW3vR6T0VSHtW6AF7yNKg9LVHIEIhHOnTjBhuwurwHwNSEnSf
dUcISPXyfQGiL7hU/fwgiUedtcjwfTNpdpXBs3mySK5yl0WmtAOK/EfKKTrs47WV
3J4d7TM94kaR7iwQcDw7JPd0jkt3pV/eUycYvRFJViKuPSAwe4J5Ktwouqv2a2aZ
2DBiROfTMwHABMxxmbfqaH1Gh3MN43xEN03hyuatfWYFGdIZ0F/GjLhWQJB7oTBJ
DxskMweKbiZn5/g5mKN08DJjtMRVK7cra1CvxLsqD/WqpgzmuXLFeKbYxZ2Thy3J
6KCekb2bQ7fmv2iL16FKH8nto268lJ+q7JQIwfmOtRhu0XADS73qDHcnqLu8NgQe
O+3oVxLgZhYzzWos8kvlN+Fzp5UBYbTm56IYeNLWlNiPdocV2EglLnRmPVa9sHVE
LQpn1VRejI1hQjSnGy6Z6yMAxo/nZg9aIgzRTubSjq3jbU+l7PW2v6tnNUsct9aR
7BxX3DkqcZ2HpMRS2/bSRBZnhHPJoiEM0KQLlxgLcIufeL8dtMr8ILh11L5/Cu+H
1clWEKFSdpQcTICPwHMRs4p5wPb+78A4o9YCI5JRuXRzvw3e0WT+sk0Tg3IvHMJm
udRVgSZurxezcgAwKCQIfjkBQRcH/FHgDW1SdJ7GftTeJcuanCO2YgHiAUNNddfL
qR7hbPm2UMAUFWBbE3xUeKesYA9i8LL5f6GzvK+deWM2GD9QqKAwNFF9re6C5euZ
aZqLjfQDQXUBa7N22DWxJ3OBxjU8mbYv1aEX7CWat7sUdVvOLrvAIDnVU6lDc5Tf
rzrsVPRHroRE5faXw8CvESONKEzuFzWIazGVW/H7QEgTngWhmNbmxVjTXKsHOeKV
7UISOdP6krdvhQx9XkntUYCr3123cdFiqLkmGh6pr7OHJZOAAtoOUBBvG53dCP0q
Kbt6gc8XCHsaaP/gZ4E/2UUlHZ4qzykxiGvhHNB6Sf9QidpjJpRY/EwPifl/9F0U
wrw3b1yitWJ+cUsDH2GknfAAGXY28UqjPkx0X1wDQHTVL/XHr/7gtlU67XM17vR9
IeAA4n267KVWtDz/W+PWrWEU6RqRpvbgMJKEdEAkGI4Qe+J5XJPK8xDVyRG041iD
9ejAxFxL2LvrAdtIOVF+Rnbxi/w/4bR5hbliDWl1ZxB11GZZxKB2axK6tCIPsvFs
YHwUdzelTUjMD2NXACf8gcFog7RGahoktNtIUWG7pSw3U2J0KKZjPVTzQ89MK/ox
/I8KGuj0Z0VMyIX6Cc/Tg/wT1U6KQuY80nfV/zRE1XoEA66e5ywARYEVZcFDymRm
09eBT70KYcy8J/+DD0ZAWTwE0IGr1zXkpFJSC/f64cuBX8+NYwsVRF03jVsj+pud
ETtcLy74UZwUz/C1rpCyI5bLf9XNseTwR7D6tE8Kvg1PagE0jfIe0SySXC43H2Qe
sS8QAjmbroTHnwUh8QGzSBpMWXGD6UJAnSpVwC9Wi4cth8n2c/pQh80tXwc69f/g
eMpPGw4xcvPIBZN54qXiwuqtujAqi/YbJlk3JUABUyVthfKaf+SIup1Hir/nW34W
tPJG7Q4UdpdW1SVjH7HbTYqZfWEcSA/OSGTp8Qf6YUwKgCxm2Jar9zAboef0N5KM
RgY8J9/SiYH1E0KBsyuFIvoeupklneUhp7km0aDRSkaNa63PX5fiHihs5Dznz+Ql
ajH5BlsbH6ahDpJP7NS4KBE83IBzXkd6H6kwJGYhWEJEgQjv3IhEoDE6VLSc1fKz
32sCUIo98kfy76y4FndKp1UBZfqssKs1IjZJDad+ra3UIOpxXcCA39cT27utyRQv
4/uuE54kvIPZd/p46Wxl9rt3Ms3I0o5tAwGesmkiShEY5EqHX87JhxGc+9/2BgdK
4rDX/qDuoas/twjOhPBkvwFQYXQJIgcOY/5uPzx3/t0OgAQ1X6e6QjKsqEz32EWB
X19UIWD7Fl2l5/c60+X3UAT+SXZMi4eIIp1OP2XfeWwL8oGzgURpPLtZr0P3mce3
RGD1MrUXX5gVPy/WkQdiUZp1IVxsDnqZHCNXgfWp6jjmZ2h+fqtVJF4X5dzdfA/M
WRYJyMksNV2BMgg6Di8nbYEoTBn4K8tuS1DztQRkkDlNaoTjhdYSIobcdHmjcFGL
7QOlXlzaibR0bXmjwbGsl9tCFy0I0fyLom9fE42TvzALeZQGASt7WGVv9qxYoXIX
eT8ki73WmrQpmWUEKqnFeYJLGW3EsjfD+kz/PwukKogndS4o+L/pnwwP35pi7Pcz
qCEqapZiCblgO3JeQP9U1gG2fMOaMw1ta8Dcf4lPbnVzV1inwP5PhDiakFoJRjj9
BA8nHkenfz5sMuC3e2wa/4WvqwLhtKMretfzp8hXP3lV3Nl5Puq4D98pFkQZGLMW
zJSL9Z5TNz0YHNIIthwjbG5pUNLrwbyIBPBRnv1pcS4=
`pragma protect end_protected
