// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VqZjJhDA1ivAd2Y+LQrfgmc9pdSJfuNau+cHBhHH0VdN5X4Te0yoWpY5/gYbJHkb
VI1ZwMrS8uflAVyh3ykYIDXQPruGSlmB+q5lZy6xrHeP4+cjr43T5zjZRUf1tdCC
AkRwyfqMRHDjhqQCQnv03YE2C/ATnvSwmobsnyH8Glc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7248)
RhXu+1+HoHJqsrKizYnA5nDjf34FOOi5LIkCc0CZ6L2CqMAOPDxIC3bxlO4O66m9
17ybeuSHzx1Dr2rHdMoQTfwe+JMecC+oTCzZ6aJEDNkWUY6gPwuOKzDtZckFDnnr
ERavIeGLYrr3hqrSXM8OUKU16ljUI0zO/Bx8Hvi+hk2vQ+NPd3+hFyUjJ1N5WkJy
OmtKeqfvAMTt01IDHwAQo5TrZlhbRVngehdUqgCIig0TPqQQPE1DbRUTHeGsUFmq
W5D7oiCswu21Ofn+FuJaa8Zpx2XopmRv+80zueAUZKIEpGmU1lJ+japlje53J9Vw
ysIFqaOfJXmf87HXrsV6FWIjgAbAhUHI0DWa86Ene1lbyU2QU40RTyouhJFcwfBQ
9WYpNQTTxs4RCVEW7D+Mn7DG57tOnAU7BbTPhKFEiMHk284Eu90Ap/okPkDWw8kj
umpwzH3k6njqG6n+v6VYY58GOnII+8CladKFZwyKxTE72QqIm6Qs6p4HbDaY5uo2
asnz7IRkSJY4LvK1ozB79EwEzNXstLx5rh7AOZH56Mg0TLeQvXw0r0Kh3mwlGXXA
i7fU3nZUJL6f/T2vBU8rW2RZs2d5VbhdFq0RLsHmvvOjj26Ewe968KAl+57q3pqp
hopMqv1atStBRgTztprUxEDDyR6xQlJfZC1WMcApYnXbHVMU8SgFH20QZWvN0RNd
06q5SaXEAdgGcp+jsLTAxMHMJQNUWL1cms5ySSmm8ZLY4cHXRshGOzUiIhQdBQi3
dlqcV9BZG91dLu4z/5GnCWArQ+1EccRSLDRcfR573ohcSixrAEHkRfWqyp3M6nyt
/H1JzQk0wW+JV7N4Z/984I3dNaJKP+e7vNXOZoa/Rb0kVOiYXZ63mGX8odSCJJvB
Lv6HTZXL2a+g8kmXcV9K7XJCQJCkXWSTmYohDiSNuz49YCv/hjd8FQr2hl9gpCB/
bAVDe/atG44pU6K8qvypwuIG5ZHBYSix1XIkqrDkslZWfxk/ugTkYGW7V6ti6qF4
PtDX+UJRU4sr9lE8rvyn6PSy+khLNDr2gfwj/lRuEx6tU5sJQ/U8SohnDyTypObl
YJbQFVg1WETcIwVMbGo7AIr2uxo00uOQ84/9JzpTA4WQJaDJRhhowniDT7pu+7q+
yxvT/p42mdAHilZ5C8a/rWMV1OxeyyCOHh66d10MeD1aAWGWYJ/neUbcBTyVqzPJ
raWK4BLw9l7hikfD5TO0QKwGZCqfZGTyfA7lM1nkCoFhy7QJlpugfl3D68ioanNW
c8PqJjMNryChT8y84pUkz6YXpdMqAOaG8W651ZtSRXqQLsiAAdj5Mg1EyihKUP16
3VSmu/J3Hx5X59/OEIcX+aPddpH1VGFnqnFqeEtjUWG9k7fDmgRqyKtuIWBowHif
9m1F2WWv35+D6ZaFqRbP4WyR0ATTBXHlEoVXPLzUZccxiPsPaRybKx29MfCWDBJd
S4oY/H9Ib8MN1GKRKXxpBWWF+/w29htwbwVe2TnUHLzjZWgLSOqjqz0Z/p5ABPTN
lpwt/4aEdJ6J6FrQnsOoVuaAr7w7r6As0kwuXXMwgw39xsZbAwaIS9HwOuKj9nRE
XgsqXaujMlvKMgf1QstaJRb2R0obH/C7P930kAE2KAsdHqwye/8LFZ6+S2aknBpy
qIxEU8p35P5Mwwnm8WI5bP0tBZjq+Q2DGT5NuYh4nd8xMltW4vngYRc6ckTrnNxJ
/5KD/esZZPYhikgX1A+eGNWxzKcE+ea/DsF4Q8bvr1tiZEs0RRGvfDHux2Tl7xgV
emJX8ycdbGlABg7KME/woi7LKlTHJ+SE8/Ps13hW//KHKZx7TxQ9t5jCeUfJiRpA
8DlRcyh5lbCv2BB77opjLDywVho/c7j/hvskt1NiLCznDu2cvCbISzYPHCvUZDZ0
+n5ZbMa2JWhSMX7mW+5u2EzBl84MB6gXf9Rd44io0EskpN0j39ERHWjMT7++8DoU
b9LKJJBRR1eIrWNUy2X4bViqyDQFL6Jxu3t8gBdeqy1i9y/B+jQ8OxZBS1MyPLfl
KJnQtnaIQCfnVbhZJDjIq2eNhehIrM2X/Ct4Y6rbFQ9xGTa7UscbaTu1ukHPNxUN
1PTNupf5rTyVnj4M/HbH1ugU43a61rJ2U3ZQ6I7dBnSYwYgTjB2QRCpT/MwVD8dX
RG0yxvjyIzq73Ui01Vi3XEFNrdqTgMq/HTn3zPtFpejsGF8t/odRBdFDdmyB0rI5
xBXUEjf3wR1muPO1S0CiV202DamP/PrFGQzzq8iwIzgbbtxU7z3Li4mISvrcGlIc
2Riw8BgF61h+jHmPDHN4KYTXW3USwMM4ClmnaTN3EBVIvIHzvzWwzSAieXvWUqtk
A/nn8G4IZtIPnzQgNcWWrYW/dzpkP4ESjf0QkkJyWs+HWM5Gt2k+/pEgFjfNjbiG
gjieRYOIxo6CzKU6KQ0Hjpy6ZkPhCJC1Y39p6WgNIjkts9Nk6ckPhvkmrLy0W4Ak
OScGrsm1bWmRVz5jujLN5FbI55281wkgBpD17St/8fyF8lb4kQsulp+QOQ9DXBsM
LlOJ+zBYQqgMlzKK7OWVrZxCFL8HTQqOXYh9obK2zz/KMyX0FaQkw4yJ7NNq2wxR
Lk/Ir/MjDGFDzY4M21iztCYAQAAOrpJF8hLei2KCdpFWkvRYW5pWENYx/jJwqdQK
30v7RbdIoqknfMROfod/9dphGkpq2Ws0o0yqCSpH1jWadUpeR3goWuD6nCcvtGYp
PhBH9t3iHbJ4zQA6hUEh7oEzWfVBg/CNxxNJzR2LRsu95FliO1htIrQZdYD3AMYc
pn3KYzUKIX+Y940r8K6eaMSmMQDs5pXmbNURtTKo7k/3mdJ1dQx7nDeBWX2SdtQ1
jiocqfdecPjaMKamk//9v1g5NsdZpMTKDojknDByeGB2RQQwMzbzSqPPzLliBiYV
uAMujmS/z3N/YRT1pMsxKnctA6qEidYr13p85L+P/uMpBKDEiMaozMxSTT+tIbKS
ivoh+4tETwBSCNRLY8TbGqS2mL9h4k83zSpz11WXl7ONGBAg6zn4Q/Fm4Kat4wLb
TcgQR/3ExI7DebTSWJUJcICbjD0vj05qQtzoIsonVgvn8DD8tXszWwEt5Guq4xfI
qlgJ9r4fe09AZAF9I4IdDZws9NYCZcqavuw5Oqkrxdsl8friwTcfmxKuUetJi8rX
Azn2hop9cKXXidRMb17kZ3MQ8QgPzchJvZcxMPUxH42B8efqr7ePYnq8nFCrRa7e
og89C8fQN9LJWc2zD0BLRbuEzrnEKqeaVm6mzhAAKPQvSQQZT02DEEQt1ABiMvO8
mAlbLOfgKse0meJmWfFkrmCP6RNgnUpSNrovwHJ3NRajoGbtm85sAi3Uq+Wivz8k
6Npwe2XBeus8dRgS+WlX9IhpHZ6y8YRQt9F8FgSm/Zs8ioQF+pd6kjyx4gBMsDKa
R7F8ZKQWR4ZrMM5hgaQxsHG1DdMGoY6Ufbo2huN4SsOBwmBgiOVGpdN+aH2m7dJI
x42m+1lKe6mSNkHR4S9i/gaYibKjPYAJGwq9QO43l+d5azv/DEgm9/jqMGyjAmeV
ES9pqeUa8F3048Vv4qmoH7r3Fy8YPFmEc8UZQXqU2iE+HLnZ4IEKT3vr2XUZRwSl
wcuPKQxywTz8Cr5K5ZDm7t9Dgn1fWBYgFt5hCJY9FAEEvA3EoUkLQ7XknDkLgjXY
IOONVeSg5brj+owLqJjo/JClF8x9nXyGE2bu1fNTZej/9z8GLLUHFU2JUCamvjGQ
k/I5I8dbQhjFyJ2LFIHU43dhV+Ka3ibB2GTj6SjgfnFWEXKbJUYPDR5AiW6cpoUW
P8ZAcK0AflH12PF+9GCyretDYh8WUEN5Q5yWahoTa05SkDN8F3P8gBEG/AIGQ2kW
eBG61k5ohkFaYFy6wpYmuaajUqrmYMjqOxDmr2wu4X4rnC2QC5VMTVhYV1WX7qgK
oKFX9iRUiul4AhaewgznArx8IuVnAi+xwX3HAv556ITKTnZGze5i2iEQmiZ8O1lI
Dz82lJZu9L2G70hhD2sAamuH4A0pPWaczAXOsFCOeVqEl51ORipOfiKh+dMrvxKB
AON35FfijrEwKkigWMsvTxr6ozvVNJsjG6eC+SfQmXF19RCsePuAeQCphGvsvA3s
ZEKDUTlZodTxu52FyIyfG3M7sfK/liv29dMRyC0Sv8dBVdlKDz7fZ9qaHL7uDtew
UGsKlkNm3kZxmiu/GC9+zQNA8EaQ7zbpinABVqEtyjV0Poa1r/mH87tfq9s2lARb
FOSirXWkJq8u84VMzbEwjWaXdZkC7LJmYXI3Khfu4f4aSyUYTxnQl7lgxArmzoH7
+W6g2S1BDPwyh8+OiKS5FQyA5/oNu+XLxA51+ZEpkCZSFr6Q6GB2HdIC5zIKnX8V
FVL3d3IxLrjgp9Ewb0WRUldrZEQJbY3YCGK0vObx34Rphk4B2SYmAG/U3QidNcjS
h6XSpoKo7uqi28fpA3NBz6iSO757hiWbXd6hUk6IdKQ4MWP+mgm0gUhATLYwVBFZ
mjLqs+MaPHk55KPrKZc3JunFfnd9wCrkuScEcuEQb3RvoqC6Te+D/HZVm1jVkzSs
bV2L2BVPT56ChLESja273GIs3BMBD7KqHnZgexHH0dj7ny3Gw87I/SYd+HyOSAdY
c5NNkO26lJvL0CHYrxvOHLBbPFDXQ0KK3g23HueoMicL1XbbDL/Srq2BLOQHg6xP
7WFTVJjLjbwzlN61xh6DDAsp++OCkNM/cPNdm6Apklj94v+nnaLoHFAB6DdoMr37
9GUDJ1lycu5UbpUfQ1mS+iI92/9SOxh0CVqw7UiqWWaN0JNM1a3H5QgZLQaQgYQx
WjmTyXhBGKHKQNQfthjvpVDqb4R3x5avrDtauU3f8o9LkmBcQX+zOQz+WF1++dEq
poyGd0np6g3IU8trE6U5Keu2BHeGg0dT4nVXdnGKts7pvCOx/ZewedeqzFClUzzx
rNZWvESeW8SL1nK/1RzNMz+NMvI+MDoJ4MOasOgF1NBSdXhwNXvA+valCcWI0Hq7
tbfx062utbswb1v71PvPCX8Oto9KvzN2Q7dy1Ck3S+skBjXh/SJW1Oa0nvP5/i/R
dGEv74b3RfbISva9ainWP5Il3tLNCsaWBLP8huKOaBKj2djoG0kI7tZ0AGBmAm7s
wt5uTYBF1GgqQqjN2UuL9r8lVWW17jE3h6n3liriCOSzec69bt5vv30W/K22l+Wd
tU0Mjno8jzNSqAVxZnvUiMO0Zwtu0fBM+EhiVA/Q2uiW9gu2tLPvdbJNhKHrRDK6
naGCIJdOaRKVsw9qJ/Jr4IqMu1Q5V7MHKS/y2NQyWj5G/9b2XOcHFmkZQDdTP9Cf
oY50ukKbigwDohgjMSrtn25CXcm5EG9cTX7souAPoGXKh0E+ZutXwY3vY3VveeU4
btf+Pn6LaqD7Ns642sg1qNnse7w9o/pRt2+QrUtFTRpaI6O+M77JhkCbuEHjCi4v
mqEnkXLuvXpmLHuReEc8tWQF3L1VhE+DQwE9RFFFQc22JusdCyD8rs89kdUotIQo
wLOwWX4KHGxkowUa+/vzCgdQInWVRYg0DXFL8qjNkp4l5uJ0R+0jay8PIO0vyE+W
XDSGSxcCxZ4qDXAr5gnsiXJGl5EyUA2akOLfqFHv8hakvBAUGAPEkuB8gZqpA1B7
j4HkbDYNynAVzldS5L9mHtxC5GhcxmVxBoQ85wlEmpiyAA7Aowpld2zK0HLazv9P
h3+zFKgwkT/sv1S/QTWLDKYveoesjGgFRVYhArPBu+DaeTnq/hhcjLfNmxaX6v3O
nBZPplAoAi2BagtO3wSKj/FwZSxeLszaoWlyiVJ/A5LrRvm7bA+6BQWIjdHVcIgZ
etkGl2nivt5jdoKxm5oZotjVhl8JCvpoPWY69TG3KxLwMMcIp3gIwPqYj21PTu5n
fpaPdCimShTBgs/5FWzToSUF/BU+fCDMLwY/AzIR8tYfcsmSRQ7+x6jzKdqhFU+F
9lQvaHkrDXmow8vZeI3TZpzHjf2Pp9rXbmHUOBllb2dd/WoXevFMLtVc3uDN4Exh
1n/1t3Oa2LmZnjRsLfUC0sSkVj6XHOzT7ForWRsHPdIeCsYQPBuCuB7ItjxvA/E6
9fy4s17yHUySEPckS9aV/JN2q0vqZ0/pFT+o0h5Bwi7J8lbJi+/PmlmpAm7wwP3b
0pkGq2ilmUYtB94jjR+OBUNyTxOKmp3DDNK6SOA1MgsKui0fehScoS4pO8NOKo4W
FDOm2zw1vCZleI1J9IVXQ/Ux/E22eInunJQCVG9QRDZojQQVyy6Hlzmpj9RAYqSy
8S48pQ1V7vSJeBfBekZFd7V+VpMHBO9lFcTIDxmCv8f6e2/q98Ru2kCngbKGMTOG
mLInBQSj9nVXt9HF2ZN+iD9zs78N/voJ9I4odbp9nvSo1PRJUFJ2beA6/lxuHVqt
FO4/RuR9+SV93C4nVvOgK7ZIq+a9FonU8AFYloZZ5uY18psK20HT0/8GU+9ew9q8
z4ykl7ohH9ZuEHxIGb42dI3yLL9vOlGYUnu3R9HQTpgky/wuR5aENvzUQ5gq7yeB
ucdk9raYWVrz5goG10w3MC2Rgc0Mptaw+d9Bw8v78bTe9Ss8tf3OANrIezou/i3F
idQV53hhxRR89KEx4Y+3qiT/KiVL4kABMYNwMnGf5tIlpEEruyhixWietT9v1Jc6
JvR69p8yRm1BcY2229urMiSC5qzewi0OqvJV1/4YjANljlaNSHRRbnZ/9HaSjyDV
qMvvdvruFGwGLShvKwhuR0p/+fYhtN5sTtKEvVszlq7WqSB2qi/R0eFIRqU+Ns41
eF8uyle2GAqfFuAgJIVrwbNCQimELuITiqlPtAcc9TYN72ParE2zQx+jD4zX+XK5
p8bWAC/OOKb2jPdJkpyRt4P16WFrsBXotYp8YDHVtoBy3itutqrOqdv9GbBnjIpf
tW6ZmSy+y/57uTJMw7qsoyVY6zg93mDIqvsoxdcBGp0S7sDGVtgHJ3b4UGGIbeah
pQPJwyxfoYSb0TWfC/txrwSrms26XlRDq8qx2FmgLfPtodhjS/0+rhEMkrcusYDz
O+GmRlc4UGqML0avrhm1GLKBgJFZ1+orSdZ4MYiG7ENxKPmCkjExI7PRcRcHuLXl
emgAOybEIuieJfnt15nlJYTcWbMCLOw3wNJK1jqDG/KOOr2YhXrWwFfEut9jmD4y
OGBMMj+I2QoJUrBVkjh9YBg32AGUxsHXdQJPI9UDNKO1n39/vKurX3qT1okQqioG
XQo3AheNqb7/SOPo4LGUoGLyxoej9n/qlYh78rb6r91cGeKDVf+W4oZ4dwU5KPT9
K7O6rz5VhEEhI5u7NNaQ+FJ1KjG7d0/9hIpIyvX6TJlwVNaBQNWVMpCwCPPun+p6
18rgMXMTsC9eabLKcZTpcjIB5LtQKleJLY7Bq98CtiJ8/8hIbu9UIlyvmOynbmNO
XxmBfSXsBYO5Jpj+neP4vwn1jbed0xL2oGcqOeCaqcd1SnPM53b4Nv8U1itk6iT+
c2nHPGHww9tLMzCUDHAZDCU8KQRrre/7MmaWWte8ROmugpvBpKAqjGc8ImkfYfSE
BNuINB1+OeaS+J4ZrZdOvtsrpJ4omrXsInLrRV75H8BQcJYoDDmfiSInKFP0vfJ8
JqqZa+UFQ4UeFwPbbiI0bf0wTjn/GIwNhePRch8dOvyxEJGBSTsDZASaMRPr79/G
ZP02BZu8jHkG7vQpPisL7dmYV2wZBZVQsKP3YpA1eBUonN4cU1gQwXy/IIsLOrzI
10rbdAzdd/WaScgQAhhPp+yN0WA6IQI8TWfx2U/qeCMnULkO1gf6NKhmg3N9+48P
1/eJJQWFfnZVwcJ6OviwYXDpRGp1Mfo7fLG9VQp+h1TaFRoIXKUDayd3tUixN8Ll
ALft47emFtGgUCo3HBj+bZPIBIYGJwF5G1Yst3qz5Hh0lHjkYJRFhCEts2XuAWmG
r7MbweHFli3+DTDW3pevPQAvDSbe7+0WEBU/Hcvj69WKeQpoLlqvUbY5L65jM/u2
XQBm191wjPqL6YAxEylUU1ghO16wxmuTq5ptgJVVjpc4n4E6nPKezjnAR/GdM0BJ
QGhftGiKmx8RAHpNWXxV+7m1s83LO6PTAOheHdF92LqjuGlPx3WtOjY1GAR2CuOh
lZovuZXW2KXgeb4Z8ZzcOR7wb3xuyCqMcz61xlMEMRKiVlcrZLL1ra/yH11+yvOX
W+uupWqI01WiH4PUT74ffDdi8/R/MLFgQwxjSzWakqGRstLPiQHjQpYg4gR6dZXZ
CYzibSLnBF7/w1jyqJS+AKSYw0UVlq0y7J6fVTn+1HGkqZ4c5j8EsM8Zi9PbhVvv
+8Q+giLSTmCfffHvgRsUznEdXRPIekcANWBqCVpfY8tHZiWlhY9r6Z6GNuhY4GtP
INF+NTSzJUXBXuX5QQVOmkDRvy4ogJUXA+I2LAxbmwL2nV++iZ1UvckDlqUWNQLC
ogSQ0kZgy9bi2tcCGw6CA0lc99RlAWIt0zYnOh7zhk02nkMQPmApe/sRfCrYugJr
w0qH+N9Hv1MKfz4aIi0mrfjh9Yk2BC6ZzqINHXpi0tAETv+0UWtheTrkaOhYt8U2
uIqZMoAryucyrTdiwow9RlXBRlyXphIZ0ePCz6JU55d0jWdKD7yOQkoS2c0ysxgi
uzKWlt0Xtg1jZh3lMcXjnHGWAEVOFfDZw3k/rBvNyk6+A3a3xsSgU4khnZ4CLx2b
wXS8ZKuL4r9d3/bAVIgvs0G/G8OS2CY+IWI8MmXgqGJ/5d+SiZiJi+9a5DMxygKO
0ZDv6GAzx/o9ar5BGaBBdc9YKmM1PRSLg91prpCkt3gryZeEdQa0BmsN9ehmDf8v
Oa8OrCncQn+MjricVr4eOZhhmOUXz4Slmct1McJNYt6yp32/aYp+m8hCsBcZrrdE
Jk6Z2FA8xkW4M1gJFtSGP24HYX3NtnEVMIU72q7g8QeGUJjvkDMUXxrAVjudOdZ7
BEK1gmGcNbmjEZoMSVdn+KGEx5R6OAgqBuomY5ZxtZ4x/rCjN23qmxTrzfuCn4Tq
mFLpc/aZRPBHiOK6TibN/PTVKtzj+G+rF/X/RAwsR5jNSj3pet5ByHLAzgsKvPRr
s5lb5y6x5ga8kRwpeTLLuL922R1xosvjq18J5a5asgA13FabgrzdGjj7siB7ogu6
4hX3SS0OE9jMdzBUL2wyYZItNg2z9pLrk7fkIqFhuOghm6IHlTvTzPol/dgrlqJo
dWEoMfz772+29eOuuCTkpD4FT8tCmLVeD6cwz4q+i3fb27LTT9Vbo5JPA7xVBcqa
K5N7yoFQlJas7PRO9xK+gxQ/ATBsFL7e0g5rq6RA91LhyGeU9tYB3K+C62/wyi9G
eceZaMS+zN62x8uLZCDGJukEZOY/bEf2A9COkEl4dtc9V/9RgPZVLt7OtPMyvjdw
A8PhT/ESeKO1xrHoNF1r+YoudjK7kCy4xP4cdYYAWOals0jqOuK+oVveCN52q+e5
HE1eDw5SKfjhkaTk2qVdf1ObOxUF+eUZBsOtZMM4l70p7tT93fWg941XZOdfi88T
mNAn0rHxYxPeEWmotQmJVZ9Tmv8QalvyaKji+3eFLB1A/sDe6HX1YAfyRRn85qad
`pragma protect end_protected
