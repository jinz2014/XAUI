// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:31 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TYQIArn9Ib4R5uW95zN+nunPXtTTJbtpu70Il9LqokLhcWsywKBPAkmejdBLG48V
El76nTEODpk+AIGNRNhhTYY9bUV+OAU455LJlMwA8axixDC6LjswZuZsM1z5REKU
yO0hI1mpLShVgEpz2OPRCu+rEHzgDgDf2b6y8HPMxco=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16400)
3LFDjsJcaeHjp1Xmf5d/qRjelNwL4s1TY36SqhtBJWBqAi8hLv5yua0Q3A9YlgRf
wS+ivbfci6gxtARhkqND9NpCjEswME+7laanPx8BVaS/idKYNg5eD4ymgUnFpPOg
NA1OvYuWKibbNkWlobqYurXiDEiCOJvjvJ6NpvGZbYO/taNJYfTzYjavkMpNbSlr
msPPIqSDcnPe+jAKYqWskWkl0qlr8G/aQHIq7nU3TULqLaUlzaCMQQQ0m7NDWuFi
PUTIolTDYd/kZqW0Ys5YL/I5+1e7nvwj8/1T5jxn47Frlt8YQOtqsz5FRP55GYbs
uzfRt9VT2sIifYLMpOCsctVkTw2rL89ZRwbQI37tXLUulAlbKX8fR8tfFNq8O6jT
Dllkw1e3aYKAWdCCHU3SMDcdF6mYxf8ow0wXNupkBSAG9aK2jQ0tmjhwVVqZemCE
84loVt7nun3CZw1B5eIyKxEP0r5NZLwh8j7FlaOaW24iZZ4miCZl1gyb3g4rC95J
iltVPueddwJT51GljdUie6PD3MYG3LpdDzPZwWdZRJK0gT4BsZDmsrFouG8EcKnI
8CSY3c89Z52kGMSH8m+gyqfu5m6TgXaa2O/d2KawM2f0cT6EnzdeB6Cfjjz8E9m5
Il9p0dSlZrm26CWzxoFxhqCtBgcmq6MF6/YugqpgJvqlYXO/aQXEEQvvwrs1kW5C
vTa+j0ONNxkfCGt4dcMSs1JneENqqhQOGWI3IAjpUe0RFg+5ww8j2GujgbcwDDh9
l+k0iiQoZJkigzM8Buv76SYHoqrHILbLd1MDSFxraB9TXQTtL3VOw8LtzZx8acTF
GibH9PK7inah5yYRek3rgDrJLCt8SEqO17tYWJfzfGkLQmJmXrkm427jxjZKBVsR
1CIk34E2wdorh+vQdk0rjj74UEkJPUwA3chCmy01sDJIyL1yijzBj0P853ZFH1VG
1GvT5yxWb5VzYhItNqndgM7dFyLt5/LcqvrZUay1sRF+dlpw0Or7478h+A44TBP0
N6Es86WYmj81hzd2RAFOvl1PTIZAihB5aMcNixWcCJ1wqlisOEWgYPD8h2KaKvFY
ThRyOTrATMJEKup5GqD2s9qoRM9EJZOl2tK+XfsBDzlnKs0DBiVCSi7P80oWGfnk
mJEVqCho5W3AX+EALOLeGFQR/b72Spkrg+bK88uzcLF9mSgjB/R7d390fo7wCneE
H+umOagmoXY73+L3vqjwGuSoZJw/JHnM82E9BL9ji+/J/B+GcednI3VBw8jnmcvk
jB3Umbh+xY1xLkD52h0Tq2TVPlsAVBpi+pqkk4nS3G+f8giFI7cGQ3hUN7Efa9Xf
zdZhJh1xf9i7Af0iSgxkrhcr4rH9mQ8WVtyDKZVirOZsrY5PRF9FogjqD+OYo5wG
i5TgqVCBP5T8cJKPuHulyQNlaY7hF7TvZvsXoS9cudjDO/1LPmUtfNxz7ntWGPim
hmifIGeU5/HBCh4t1dGgRn4sp1crO9/hm9+U5+JzKg2Vfi8Pzrv5Nzey2PjFqgPr
pUDMLNRJceU6IRnxi8cBDFkVK13Hc6ZVTa7ySdr3VBn09g3zR+axIXyxuK83UBFj
JHL7EysgTMzydlVZbhWwp6g8RCXNNtYONK1fF7u385y01qm3mvKAegcJcOlMw+GI
6IMD6bRLJZGrDizd/2Keiog49r/ubPjRpcwpEUrwgSAyhgol89Cvv+Wb7CFcMYYZ
LKKkyC7A5CXukK+cumvbdc9BsRtVzh91hmu4YZ5Mh13wfhcZ5OEWflQ/ctQF6KNx
vlMM4QX+ZK0wz6K/e85JEubk0qNi9KVk4LhqJEpXLcYKML92Jkwf+rOKC+CX9ho/
8SQz8UblHJb4cFmHC93DlLrOFaBd/nVdJx+3923YX+7rv+wyuzamB5Q75Ys5duOi
jsSOsVS3evtSNzo6cZDHScqxknFRWFMk7oHxJdFOSwu6m+O+YQYV70Wwmy2j2/oS
v/+6XbK8durw34FflTsT9SXQhhQJv8fDIE50pwMXk/wgrB7ae7+c7Djn+X12GL17
TWjTNXPC3FhWbN8P559j3XUm1bb38WblpHoydSF4kJt/JoU+aCaElq3kUVCoh54T
p9uVP44L8+VE4DaY8sUSJxd3B7kxZOmAamgmf18ChX3OFT21ayjdr5JQ7H6i7JVn
nskecdnEyw3p6Rf/mhTXGbAMGA/9uiB7P7+wit4ei+WpxoBfvZNhzFb0UN/bljYg
TtsOtQi4hu9izrJh+QYDovvQkIW5EZkPQz9t9oZx6hGjnLPfI801xdV6svJj90zj
W00rMNaHOr8/SqAuD7SloUGLmeRWoHTxjOszYyU97AIvvgSZnGN0CXfd/f8uWcRE
/gNloUIvqlDmQt7t/gKyooZK8bGP2zbhSXFgpZ8gx37HUmf+LoVanwKvOchfMFQG
oMmvn8sTPf0F5xNNotXR5MoncJsqzVASE7Gu5WH8CGYww+A0V1uWjQEbaWbpy+5I
ldwdpSo9Z7vHJhHTDxL1KXd4zA3z3dTZaLzaXuM9Rs5Dr3//urEomjac8ZqnPc5J
ODxe0MXskhu4OX+eVQTd3KAJFRfLTb15fDtcOrCWE4PCSwXNIyNJlD5OxAy+TJjr
33KWQVBVKYrGb1RqhI/xDFS2fzwkZ/ikwmEeDQDGVSg/kmDe6h8eQUcx1PRYAQw/
RzUfUYQmZUHw5/pZvRNaUn78zuqkMfi0Q9lmC0WN304GcDyycN50n/ydHtJMVReP
OLpBRtlzlyfqcE/NQMWrqZJcxZQdse6I0JKieC0wV5BR48h3eP78BsW0NjpI7m8/
cBNsvtk0ey7n6oyd4/FjWJMocUpEoarPBRPKZONUGTd3YYeJ8khtrGoTD6Km6HaF
3g8Uq9FrbJ1FLO05eVyUghBPAcDs/t/2QhbuNXro6WHKK3aDIQwoTyg/I2rs97kJ
m8Aq6BOVz4KBnhyhdRQ+LzxcvIo5UgRv+AuV9lyJc4C7AXQaxYglO/0YUbMaSS9H
TtUBBORtW4MyhQev2titxWfZsCknQ0MX5eKSU0m1WAfQJ/EagD/aIIOJ1uwb7qI0
2ytXTaWMYCJaYmP2YzfJpUoPQxQAB2KhrM5f1ame4+RocTErotwxrgRyn3rNpHRI
ecdqAOkVcdRHy6Mp686BcvQH0ijRUJxhCBkvtJE+HvqW1sudbykY/RuS81gF8rpe
n8PdC9rMKj+DrDLe9m1SesuREXD2L3JIWw7QwGi1fTCtt/YMnx0T94K1ODe2UzWN
uGIxlR3T5cK8PAdC9A0nL1B4PIIvSi0SqW9toC4vmwt3Y92o4LMU65DfSvKOZ6yd
Pwvw7dsHkCf/DwGXFGEyDPBQKQv4/94WmuO6xdunoP0HpU0+Zor7FoUimA5Nt6H3
UgDmtdUpDvCJglEXU/2KUWFx8W11t2diDUveQWvnie9Xf6RsQPPnOpYLpQgMMZlQ
97o+mgS6KQE1CQHvq4jcUXYdyDxFBGIA2A1cmFF1aKHHOrjRXJvk7Tfg8qcVXucE
kqjWegVZd3hgAiQ47wlPGI9is9HTArbqImxBzBgBRKmTeQNZRwlaQMzD0FmWLmV+
U5EEM7ekwWz8k6mhGlz6psokDJ3WzBILB/CCCUE30oe+WaLWVEfJgeWrbFqbYsFt
pT+WbA50ytqpvmrOCX8LU5lWdqJDSzU097WJNlFgvVuD2PrDsYhcm26n2oTvQ2zw
8lQvhKYxAbvTSs+pJJJIwyMtScW/n47ArRB4+6o9pFKyLtJ0twt+UqKZtIY6BPu3
73W6SI0cCzf9Ix+7HeugR/QOZrthK4QwtEYDZptNbKhX1SJWGCBDdoF83SvJCqq6
xJaBbkZkI3rv00SZQqj6n9Bv2qlVLpPWpx0h2Gd1pMDc+P07Bs7ksrf6eMv75LHB
KO1tKRE3/t+P2jLgDxeNDqU8HYOsqWgUStBsrLX5eFhpcHWJkYoxHtA5Hg8A1G9Z
7mv9Q4V0dGUazbmq4h7FjNvZicTEshqzXMd62mrnX4tf0H50DcJmvMVICfLxcQJQ
3jqkVyZ0WQ2A6ttTkQwNIc6v0IlSEfYn3vogxbihUSvbzvhUnE462al9vdUs8yEg
EKfmUj2urTPWDj/XYUCOJAZQ5zcu+oxnCwzlg8X/45JJtH5f5TcMZLte+g5RSXw1
pSH1V2q92eOhSZhH/OyaRDbhTe9qEg5qyiBKgwKMJfGUBzvS5aiQsnMModOyIFAn
UirjMDD0gXkNO/uiNmFsbMCKnRvd7uKkEIMvfxu4niuYDtGZFZ/1IPhCEvHOFvqQ
KGaArgR1l1oXu9Y+UNpCco6jHTxcy5HgieXxL96TgVwX6ij9vj7HYPrHjMK50e4+
BJvSWLWN1G6Y11cmyUYJYlYj9NJzVXK9tzAR70a6FkUAQRWVZQF65wBpXfOYwr5t
qj8mziGoRNtrW9kJX4+uGE1ySSiE7P0Kep6dW/kThpzYgIqUr4guCKm+EmtWMUTM
TOdJkriaL4UYMTEDvsBmnM29wMSDExeOf16kq96dSlOfDjMqYEo2ZxBz396CCSSM
WZ5Ay0Fh5ioVu1k8vyZdhaDBgitGN9NhR3CxjXvnLYXchIzJc4ZF1hfCnTQOTZI7
g4tgKvKk9jdCPDFqkcRXBbxbSiI6rMw8/sbWyi4Hgr6e3W8/rm1X/aPbgER0jKLO
8nHXyEoCBo/EBkBSHini3TKjBztQ9uIuqZH+goPj47+QIIwwFPvav68GCRpwInFu
q1Kn0xjPLVAfxVFf45jd4Avm6usI1ma9Z0ny/sOwef/XgtbAlW0CGDuI8ifO3AAJ
giaRYR16IywQuNeBxBIkA5hzOTOFZg5LYHRsb0ljNG8edEEytt/nrF47WEIxcROm
UKPVTZsBaahaHQL74yDgEx0WkMcaaeTkFSRNxySsFmn7NhUEecz2VFucGdKHPlk5
VMVxsbEvn9+3q2WwiHaXsh43bAPnGINHvQo9esaTOAz088feSXaRcZncLw443ZG2
qrXsrxg0r+VLDjDC7S/GMp0cyYmZGBN+BXtHGfzhUxUmZPVwKKMzlzTb5f/TE+7U
YqJf11N89FZKmfpo2a2fzU4H8V9U+xafZhOAT5kEzKvtj9rCTCoSSALCJ+eUwtoT
bxt4vVbC8OXf9QdKJRBwmpPyayZMO2t5nJbjJmUI+z0YMyTTsk8iLkbS7YEtiaxu
hROnY9gUjOJ/jH8GSUwCxoAsiF/holhGjbslojP1iLgFbaC+tDsasS4yWTzgh2MA
h5rMlZtkbgBLOfG4LS68kBrbArZTTkmPPoecBAKNfxFU2FwZPgDSUUdA35shd8k7
YsM1lNgjxKU7dSfHirZhAFnWVRMBpgoCtSZzCm59UWDEhqGhvCTvwssm9zAyfawW
tl9ZhI5Z/ER2+SpUC23AqFBnhkItiNLrrXkQZM+dygR76XAXxMb7wIUpZfQd0eeW
vBsJDouBl+mfXbfePwurSsCN8AePbltwCyqJJn5gGInkHdtv5zxMEaVvq5fn80Sz
a6IFchx4xKb+m14ErbuW4EMWW8a9KIZ0zfaGZLEcnSMLD/YQdwzX2HyzjKyLjHmd
NNaex7FqIH+DXk1ozHYQWkS3/v8kKkFRAq9TlkQyp6f/JNxvVx7ENDDDSwRSpFdk
thjMK1LZVIOA24lMM6t3fkmt4qXcq4XpChwMZ69VTrU1/NtDbyheMl04QDRcaKBD
NQBybrp6WMvjsX/cNg9fLr0PPERwqOmm15tIMcMKD/a9o333sbggVuTHPb2j2uUX
yCQfYVg5OITBHhcWlBuZbMkRtXxVi89Uv2UXnLdTXQ6xaz9dJdZ4s2GkXcoODcbk
JcZcYcG2zuq8zS+de4YiAg1AwkAbYJgwFONVZHRGWKXcsnPkSgWuFj7ystQ8h/5G
0sNEutnZ4OBncduRKMChtvxU5LCjaP+xPyjY0CAmr3yB1dScJgORquzd3tQg394M
Mn/89DrVahmReBGhEIkRtmVj12+UlqEmxVyoROuHWlr+1I5RZY7ejk2sdZlv0dB8
BiWQ2SiGZH2bn4Qup4+DCCMaWhEjz0Zw8u5jnm+1ybDlOn4tG8vXe9qaFRkLez4b
RrH9KeKFKvNT2qnh9mAxuKHezt+csh7XXtoRkZtJ/hKN188mZx5NooV1UK6HFAbz
B+6fXSoszWuZQJGp++p25wcxMuq6UrMIXGsUbf/t+aU2ZWfzl/av/C94Ows5iZZg
MqAE1wmbmg2yhOCOe1t1dDXAi+yTyCASL1svpsY/FEZUU+tMSTaG6yWv8OPKSqmq
rwVGtcNKzAWnTce6bufaK9e7Agyy2JZsM6ryPFwe6CePpGb3yDolJ9efAZ3ZpcL2
LmTxPPYdH1y+QyfyExI7M4vbjb6D7jL9u9MHhasFqaTfyRD36zXJmSvyDdJzU6Ny
qieOqUeER3aiUsLckweP5CuUp4iFwU4sR80e8SxoXrMhwSHkDjXOsOYBxYE4PrKG
bajJDfav7APJDJsug5VwNZJQnEJMBGfKzY9sxsquW09GaE1jvQrzUKw2fwdoJ28z
gkMlfgQ2SHVSGNzkOhp37qMBvJDhtoca0KX+tPg1evhTfAFEIdsAoA+VyOjAcFd4
JwAKTeJPR6YzSePCu7Li/O6/kWSJDLvGH6wokWvtEEMsJPo8uxuyo1GMOCw9Ojjn
M9tWJfJ3pZ0yWLA+JrdOzzCnZ+QrnE20VmFEEzH4ATAUsN7qJQurSVcBxgdpD9jr
I5laEf2ZI7pwpVtLXzZu24fdELC6jrljWzTfHBZ2SftBQmG1+zZF+Yyr9YE2y69K
8RNIglGDTG09p/ExT/VePzpNhif218YJETKbBD+kersZBU6R+JZXInlgv4mZMkqp
UMTA72CMz4tn08rONDUY1OfzkmcZmFbb162GH028geYCcJ+WspxP7hdKc46iTa7c
CvZ+W3WeBV95cyBVAbLLMWH2lAiUtrsNB43NX8VhRN34rKYV+ntuJzOJFLPS6chs
PgKObyQxS7GS79TDfAHJg1eTkwqTy9L79qgayO2+AnqjNKeeBlRypTCoIaCErAX+
hPJr+tr+Txz1ZkZbMWu2QB+gxwDfQy18axVL8n6y+RSkOf9PTYG3pzBJube7YKaR
4FC+lIwEAgwLqmWHwHEvQIk3oAW7x0x1gDVCjgljlVZM1KcWN4yAvOaN9V1VXbN8
Qo2IrHmmEuWhHxojA0Zoqrrg7LR4TrTH1hpWcp8PtLgD7coUhldCgEYJKLsQynZM
hMu3fStqvEDX/quU1BnGI8d2U4TyXkobaQLQhh4poJfWt6X/E4GXzpgAedO4p5Gl
/zsLR7AFHL2AZDA90msRguV5K8seltk6rR0/NMbi6jY5/JodTexhZ5SG6/l3qe60
SBB/iAuPFTmkkQZ4wqW56RQe8dIs5PU5YS0ONhgLSjnMwh4nboZpOpat+67zJMNl
ERX39NQMd5cwZXlBhEzrtGyMhma14DHRXtBbddLkDbkHe7Az/Y/2WBo+6faUvPxy
Lzsw5MAs+hI955bLUtuIWAWcjsKbzM6Qjn1n3FZV+zOVZuW9oRlKS4h3pYnlOC56
As2+Xo8AXveFXJ7lQ68fOstbFsmOEOsBBg/4beYwTKjPdiRZ+Pw33HUYxAwquIhV
/yopDs57N1LGikncQiRxrKuN+0fpVD5+AFS51hzDTKfR9TG+fItFqcesy3K3IYtv
mJudCUxV/pYaKk5KUtXnFJkDafxJgDWqLdhbQRSxkHswM2SOU5Y21CjwBhIOJcNa
b9XWhCY+W5WpNc05OiiwfWz2dSr6snPg/nq55Q7vdLWRq1BKMK1A6n79tZg/JCXP
no+ASlBmFtii7s87OLnOh0PwAqIotEBVzY/F0HpAq6XP9x4Jp1gYs8rAlSBZ0yI/
3mXWyBUw8/YqEIBlB+jmq//MtniDocJaiwG8DEvKNNbMzIZ3i9UuLCCa9zgXiaC7
q514+dPSkS3jF6xsiuZknhYl/YtxJ6fdyrh2Y8SYD8pFfNJnb7GisBqs6VpQSlln
a0yC6yiU1KK5xRR7h931iwYD97HkGb7xUDhPVV9jxHNYyXJTHksRMb4/kWIKXUev
NaA+PW6E7itu2O6GCLVAAH8X7ebliMJ+7FoRsvwl13jn8Y7OdsYbqcOqVl5wQ/w8
2NUDCYQ0cIi69byAZPvD43hrJP6eJ7vaZHgldA/7M64wY4uBBWJ0cBl7aKuUU2JS
hTRxsSZxDH/iOYKMqJtso3Cl5xj4NN8u3Xfpdq+yp5nBeWxVqRIGnHW11sj3DOpV
Va02n+fpk7hQNIF9cgybLDY3ESTxVikh12NMXgqdLNEx0yQxY46MfRPpzpe/FxRz
71fXdtNp/dU7urTlV/MXA9IpYsg5717fBSUeYGR28XLoSA03i+8iNUc3aeamMj/l
okpNPwE8vYp+8Jy/oOfujZ4q4KPgkITE7Pgs/st73atCHmF4vg59hmW9/6NjGTkM
/mjNEb3Dders7+y1SzuX3zfPg2s39AHuhLcgaXL3f2U2wpTumNPHd+HpoxjOMObT
QcfBok2/ZBQ3EFG3Uy7u0BnzUuF584YSuzJx+ELHaVO4CmSZi707Cx7K+6B0hXbS
Rat1PY6NA5hNhQBvVY+H/a6AU20DRNdaKVdbf1qnF/eMC/K6T2n2M1+2P2XTLdW9
ez0YM0sNb+ANbsM9mp4T48hbdpi3X9irwTsRn0Nnc6ckj375I9p6v9Ldrbt83oGd
WPLba7daAI8ZXCMPVz/iEhrrp+jbzF8WWlaBlcoIKSBQxXShHhrHCA2VQIquEUXa
4EA+4Z0cQTfOQC8DB9TrVzw+AZSRnebJmghmWGuJAKRCasI2U9LGhq7rINrQy8qE
KnCGUJLOk7QBTXbCHTXqIqld0KBYEe9omGiXlvPVLzCotNtU/ph+Ga+MXFnMtJOE
64qP+E0IzwmZsWW3bwwvashelDXiFz2el6fWkWhVVACt3wYn04Tn42uTkgaOeygO
HMunJNEuHP1XFTTEEdfxz1twapTkDyUd7NIzi546ndBZ4Bh7RiPvJlDmWSNiYTX7
rIXovm+hVGYMZZXLHlYyPz1pd0iuJtmsphifhfz3TqlQKwItxVQeb6mWyLAul2jT
HhC60tLnMF2g/JFbTjPrzjm6q+MyN1nggt5iwJBCih/kfGBuzqiuHmeNojRa+rm9
GKHauLeP1Vu+puAx4D3DlDtossH/BRdBbX7AdsCUqeZk0p7jBg2quqtj3Xm7y7Sf
ngtRdzm3PUOAfcQR6Ukw5hN6ZPTxh/6QdZ24wIjZtGS/qnh7y71PSsD+DTh3VwmG
FUrAespNhGtuThrxZBRgHvVSWPuDrf6AylW4cGz0U85sQAmR/XB8hyl7s7syEgGz
VZ+0jkx4memE387dLOJgYbh09QjYOP3QTHNoMj4GC97sPkYyFb0vUPpgMmJDHQrF
YsvAOwK8S7ymCFBoeNqxpuNGy126aa5thnAQIibYorE72Sx7XIXS0bOQ212xu/S1
KSbVO1/B4Yx/s+orjm04yDjk4xgg/9ZMqi6vbI+/KGehzepDuvRpoN2rf+560y0N
u6t5Bsjialik2AKfv2HdQJuGDYWNARs5JWoodTxNjD8B4C4SLQxBnTI9NmjopCOn
s3s1acJZJzmSmJaiq5Ubx81qLNqOG8qqZ+9HnqDbXSqQj+EQdBwKT5Avj5jS1Wh9
MemoX4xh9d8VWgQHoboQIzNjKsczHhPhwVv1Nhr3WRim269kgrrmxF21YPHjrVo1
GK7aHOe6lgBomzc7bIJrJFdPk/4Ggaw175FJWl7v4ityea9vmjS2IMHZSnEGkPct
W2D2AXhzhw8lbiHzJ73tYc06giVQ4QByIM+82fQU8jCPeScJAT/a2zQ7pCoxg8AT
Gx3VAQExffhA1TgY6uWW7rP8DR8Ei1i/9yDGH3sJuzreOTFA/pRH4Z4sT0VY8iiG
Ti9iavZyYd+LIo9hNMGQXM8kYkHfY/1ZPAl6zHkLX6XHiKHw9kkyIrJ/X5sOoYHz
/KcrfzbcP+64URPXdUCvvW45SBOQdgHG905jAQSSUZZtGk+VvK5D+aspm2yS9DJU
B20snGOWNi8uMnstrMXXUkR7s2BoTKUWgWN1kqNYYK2JRYgCouU4qme0tgaBuYNy
g+co8dzn6V/X3uQGT5mUmBRhA1yn8P8DIg3n4HZvpndOChFXv8OJU9Z39R9BXorp
1K5F6hu1LrKoZIMqZkK8ZpcRYivgKtFhoaTw4XK2q7mKaF14V1k3BslAdse0Bkp1
Yo1dbg4tuuuPZ5gHQP694Db4JgYNMW9xAf1DAQgR6EuAbCCsj5anuIme/navqklD
1pwyXo5x0BzFhYZCtE3rKd2kvZWN/Fg/9dJF6UlpzLyF0zmZ4wTU73IneG0z6Yty
pZtCHQud2vfVujM16pzekxqLOUi7dvUZ+mwsS5oaTEe7KJ6HRiLq2LfRrBNGM8n5
ZVzhMFgTO4G4VZ94/MlPVEiqVY4Xt/W5HciU7Igys/wZgNN7uD/v7XsDsvimW50Y
WPs3+KN+H7018F0sASebVuKg+SRkefJFW+R1lnbtp11GIR1YtqDMLSfCcXmEdZSp
dIs1SzUqaF+4p8BVRHfU2+dBWRLf5AL5zESMHzJZdsaHLKkvupX+TmFaSsx1i0m2
G/8a0ub8vDHnGI+ts8Zu2gJrxWxYCVsDlf+cihyvzrNRdwvWJlkWGvcE1FF+JLUo
gdC7l1RpnmTQQ7Pn7jQWR099i7+3gyHw73pOeMjnbHwvMmo/iASPMf6RAcU9xGO7
TkGNCSXV3EinzUa0iyQJuCa56toDjIjO2TVk0QVQij1a+Graj3czMHXn7FK7Bota
AUETS5/FebQi5LBsG4gbHHIMjIgrhL6rhW+faFCMkiXZEK6ndBwe8aO6PXxBVk22
l4N+Ju5vhcA86vpaKNwCwSZ4w0tJA7I4eOymEfhmf6y8ogs+eLjsnyeH3Tye2fh6
a//ByNuRp1Kh5nxI7JyIi5EjGK0adrKoXuhnP5+LXiLgvv6XzFm/qtua5oiJvF0l
IMcYIQPze6WRvgjYBhAw1K5hsZNGnEAiFyEqh/NNw75ux6Y3Lf8qyje3si8yKuzM
Jxsev+uiAL64OamUT+yHhdiEljJ40oRHEKsLKOcgHykC6yA7DAi07j73kLvVdSiu
Qg+2JL47KplyyR7YBwOM038kEUdv2xtcR51pavz8OJr+qycVZc57IxtpMHPvdMyg
VTALVYcZw+959ORwGrgGcsaCDOZ5ExaG7KSfArVkXKKNjWQcAei43kkdrWJ0PGnm
xiepauXXkl1Tp6Q95wS5gUe63Mk09pRXhnibooJkGf4I9E9EL1r1EdSQDy/20/QL
IQXVG3DcstqU9Cn/jihWV4h70nba8x44WD4tIzTRct4Cb67RZAzcFpICCeQyjqfi
O2++1DZHM0Cwo1Yjatn8MDF0ZSOrDtLYegENLzCWPxq8/ZeXSnF8nl4o2GMaDvuh
EVCMy11Zp4xCmxpF/KtR+Ph14jbWUCqnpATvNFMh6tdltN+XI6yf1iMgUB8ES9ni
ZxW4uIZ+6R5454KsKW8gFa66Qn7EXh+Ri7pgt0a/NiXk1e2S/b5HU0ALx7ZyzaLR
zXkdUNP+rJTfARUzVuVboGidfd2N9LWwAEC/MlUUiiJTEGyl1wrIlE8LLlCeMlCg
PfEAlaInPNgeJJRGyIbatfOpwoyM0b/+xzYoEOLT5/cKO/aAVck8rM5TlCotIgVV
sFWx9+X+yCqerVmFOebfKkClHYyisnFLCVqEbRN2644x0H70aLZS60tEdJstKYL7
yE/s0c0mFLu6GqjGZUR25/FJenbppZfjrSr9hm7hbC2ZjdoMKx63HmN1KCV6IBbf
sy6GV05XBAwESzAQWicFyzf1uqp/MBIk4nluZuc/isdbKWGtnLWKGZXkHWQ1Cchy
6apKbJ0wm2P6W2IiZDgpI0q1St6q3xYfun43/2MQI+hP/3CfvEI7cJg/oHfgcoyT
f2wF8clB+2BLwWnp2CWwY4LbfRQAQHdyFVXrqSQxQoU2R50CFxio9otXSo2l40cj
fZMd8TO6IQWVEIFxqWi4zZRRDgcbAo7EwmwBYPEplNmXXSu1KxzQlairVl0K94UH
aZawat60m78tGg7SProBRCWbCCEG/wBgfuyP+F88D9cphQKZs704K7lX5QVMjdAk
E+bwbj/5Px6opFuVjg03X1LP2pvcPav1FDhxQZzjTu4Mn0YB3UJYVRcZgeBEQLgV
QPEDF4oRovZOvK3qa5ckG8yc5JLEXZAxMYhPMqJdUwzX212N8v9Mq1OoBmlFxVDf
t8szgOmUtqlWHzBIDymilxDqNOeUP+d2NRyLlJin/6GF5P9dD8iUyzzAGJcChQJz
bb/M8SY7KJwYsQLMmjvKpDtgXv+IfewLfr7aI5wZMeRag5ciNUv98fjUP9cYivK0
v+A36ZqJVSAL0/6CaBUvYURTwjtH9cBOW8oYdLDp3p+e0W2YKt0XSAtN7jaHVddJ
fLsZmrIr8LQOHATqqtdBfn+U8Z9swV5V5j4r3D77klE4EhS5Lf5lisq3AVpqGmc6
vwHrsgLfQRIehGqWdNefc5pOa9c/qXCWpOI+IlqyKYoWzgDhMWpWC0bIlGmuLhLm
YORR5S+yPYndvkqWObnHtHW6oZMwLWDN1Ch2hjFkko1e2VQuxeCPF/dR78Bb9xaA
FIxjehJkUglrZtwQPy+JHZiYdOddWIbX7PjKwRg6+i0/d8eOHUr3zJYMuTZhSjj7
6liI0OJf0k8DVXntNY8jheL/Bd61P4bVkmAPdwm2wlTS1INW9cfZ8qT3gUWavZrb
I/JtfJtxj0WIQj1Vi5EUE2rmhkYHw9EFP33ofebYhb69wFXyqCHtlJ4G4SimLCwb
esCLhAgDvPAcMOI/m7vQEivpsafbrb8ZujZBWdHgoKaDArtz2+8xd6sdhLmAibSM
VDhjfYyiv9MZ1+KbNj2Gm3FoA3rBbuIQvIUN10GqnUB+Ct8wrUxS6Tmo9BzBmIFd
/v/cBy3SG2WOZCR8kWT9FiMsy+mOBaFQ5DcC59SCuHytcE9tonlpSYy5oJrUvArX
IibFCppm9SMkA/WMKzrhNLYTEi3JdTOmfJZU7gxC8D/O1ccmDq8bFhZA+WV83LsX
Ji5hIHFAaSJgAr+CDQYyLWJhG98SgJS6LFcQcA2oEdCHdHlgHaA7Z7Ks6ILGcWXd
NNKtjalsaH6QxDn1lvhU/8NtuDZwtrsMn9MdFsBZw3R+6O7RjOEMprxMeUrjGHWu
fzPAxZ2kMm+hjwWVcxXM2Vhp7qUyvya0LtFL7WvJUDCuDvVChn1Faq7WI67oDGyn
z/Y07UcSoom7y7a9O0EokPUHiK5Xy1BPjKCSAOoQ6J/L+wehiV2sR+jnXpyjXLJH
oBcgSAO6ymF4Pz/yzT/vVARlKpN1lxC72RGdOsVBFCJkS9ME/WRKh/mkWBmpfSzH
Ou9OLFCJHemhLvfG4gkkLJdM6YRUvKJKVw2s5PfnwaLrG1xDVw8zqB5/JsnCBFaq
Tk+jtPrRwcPT3KrVcJWMuU05blDwT3CXuMPNUxPCKQjNmLLuUN+BTIK5CdvONZGK
haii5nM9woio5I8jw2Zdlh9AFZk5TY5NbXMacbM2jzbhJvRvlENF0U5BRQHf4ToQ
RhTdxWbNpX5GVc3y5McsEfIil2xm9iE9jGw3HgEvp4yc14UrKt/bDy02FuI8RpaA
lDR2VthK+PsDJAsMh3CHKUX3GiCMs24M7I9waycRkP/9Tkdj9VkLO0fhISUBOrCM
deqFTXEcHTfHBKGiOOKI45RM+L4rNeia+sgV/HkXkQBPC2+ogchww7cIygWhPgV5
hP3jcZU7WChVu8ikA5bYxceqgDowkNltCjX6XUvbTJGZgwOhph9LXYqPlEGxiiXZ
lcMvAniB1NWdnU5BYAUoGC+zUnk2kRyS3CAlLs77DVOsulZrRJ09vUXJAUBS4MSO
iSmtVRE50Sr6GHVlvHqXqGZ4txIRA1fUpTMLc8/yB852aDjl805VL9y38L8qWDu3
sJdZQ/M6VeLWBdB0xmrTk58IiKzE8HsZIziL/QX3fTE1be06vgzoJcMECC1ZnLPN
9tdK7ImzPfIuKnWIFmCrZK5WMNxkXTbB5WtR5X+5Hj08EKxYxZl3nwJIfklBHdly
MK2Zts+fL7xyKwbFtlTiFFHZSbk5pjVZ7GkCmA8lSwQHE0/ZxJQibt0LHIHtN1IU
5KVemvF0xglZ89ctWLl+K7i/FWePtuf3P+aC6pRAjlqAEYA3JvZBSDSiUGrMG2Pw
qNPXIPchWOF6XgRTfA10INaS/JGyQjvTVJ7UsZM+rHq9+aHwsOGP2+1b71DhlDUh
EXet6nAV8aWm84QXRJU6lDPEn+dNfy9cdtGtwvqQbgH0qydFnsSYy0ve5WoVDoSe
jfDO7IkShWaL7bYfINrRSf6GBci6FVOyuvM2HcWL9qaZSrL76Wr7S+4xTOfO9uGD
piE/k2TX1Q13by7MdgVxR0Alzlrb4FMHZ10G00c2yHkKEY4FsOpHrch0CXGDZOVN
ekbVUDK0i7qjIYufyswfidCfoMN05o8NaIs4vJxQm5mcoewm5x+8fct5UNj5ryyD
tGVy3pabujOApLi4KVsRIsgbI+RNR7j1zsk487I/9mpxu/Mb2+Wgf85wRM6qEpSf
jC2lTv3XgX1zv067QDqbS1OzuQTuq1W6Dkaay6n0byXkzGC1he1NEIsGhkFyAEAj
DjK+QCUYmBbitqgmSQdKqmrQMdHrNr6UHUTT3dbQW3LQt+/ZW3PqK1XCbPj6gqCd
5DA9nQf991RrJuUySIGVZVIVZPyB0EWaPYZ62W/hcJbRvyA4Y7/JiaJ9AR5AH7Hw
tvmjuWqZ8Vi5VneqKl/HBb2CsbIB5FR18VVzpv2O5ghp5kp/b0yOlwXao9t+QGv4
sfnbNRzMT9mvzJ6e7MVpY7UHkB7V5nYiCoYXpLosX2nQHDdMoUi+Qcu5iNfoaxd7
+eRZsWfV8zcp22hn4wCu0WGLIay1tm1adZSOksoqNm5eB1y8VHsATtQNYDfPwIlZ
NySgpm2u0WhgmxUlQ0tF/VEW4dlbnba5ZnKNXBw7rNib++tIz+FAgZ/wRSMhvpUQ
hOiYwDE4VkA+ReFnh9rdvZmAOoLE19xAIsOAiY2s6IpkV0mhWlOSqa6x0KW/oGG/
v3mNc6Y47QZm53kaOB8IbNRzx+hiy3nNSgFOkfcxREmdjdG6Iy73nFurOyWTtiAw
eTNZIQ4wizuv6VCvgWnF7g9QTpEE6r6go72D6Skvv1JYJqdogyK6WMAZoSfSk9jL
yg1BqjyMTQQ8k5ZpuajONsLGdMvIGOsCo5fi/2vd+9UXfoMF3pnBBjLeEYQGDx4i
EER2rr78wrjN5rkNNTj8eNsPHVbeu/aIGz9iMLXpUUCdsCbqIept4Jw0gBONhqXu
MOsvD4eW14er2+3JJCAkojBgEb1oBC145pPXyIrKRVPzmaxThUL7J6SaT/MwqdAM
v6UuURZv6xRNHrwgQSSeo7tyMg5Lge2i4eNd5c9U8vG3pWImynXwuLW+SStXkjS8
l5QDd1ynq4Ax1Om7AjBoAf4XwKWJRRZPyFomsGB2RHObzzbdM6Rw1imfGADueFvS
szDdcS9wC15DOrlCYvngs7eHUMsf4rgT4klE2+aZ2gX8nHaySrEY/SvUckILKbiz
haK6M69TMQrA8q4Lb5NMz6MvQ8h6Br/eWAoXswdyo/qoavkqYdEeXpj6ct5Xlhl9
CYLVsKYINN6cLRj3gnAmHAdADAaAhlrpqkksUKc0h6ZcGZ6olDiKPD3pTpimEUJx
NT/UkTmdEl2p9JgNvP/jzdDz5/0ymoHr/IF/txOowtFZZRNDIs2YU1leYy0aIXRT
lxR1g7zyZucooJfZ0pYQKAAKhhkQvdbxsTHH3/bJszBtEsS0GvDeBOjCTx8KyZSX
mvtEfZySdEPOGpbDd5nQ1nmqvwmcj0FqzOsKNZa2nHy9UGJrjH/rby9y1EBT3JXP
cK1gn1C58WkoRh6L1U/3b8zsyMh9Lmj/RzTQcN43tjdhe6kngBJaF+oIcphlOXsF
T9p8e58wo20mq1OyBhFGb5hg0zdA1+oLEJ77dcvfCWxBtXn62jHq/JU/iGJf4dgn
U3HpuDnakgsD+FNL+OHJtL2GJk7yv0GDERRBu1uW/eMSrABTEYhEUf3pnENyI/L5
6+KoiFF+doEAJXIyukG0t31BXs+Vciuht6kB93kZUhjnW0xbofgDuEyM7ANWRVEy
Mp0MEMgnZLg3OVC//3Dz/7S1VI+5XgK/1PCLVGd3MJwSNtbuPYFsi7qvzNQnCC9/
Z254YsA8rzsz3CGo3fA5TY7gH4LJlvjTfiIxUGzoPmpI8TiVT821lun5m1Ir/TLE
UHuJdVUYFP0K8K63NxChJa2or7sFqEFNhsi01Ms1i7jC26ABwbju2YTUyWSSeg84
icJu8Qi1QNwCNnMDRe5sipabrRrk1EUaE4vKeKoV/lPmFC1kzeDPaz8i5jIukk2l
vAl59EOajNpwyt0k9L7hQe/icwp8zTQS0Mugy94alSobgvZwRTtdV3piT9zkgiJ8
Iqq5mq/W9CEahuKHgJDqsCtz+jy9+p8cSDFxklGwSBbs43pG5kTNRtIs9kGwzB6W
na/YeNmPruhpFYQWQT6SL1fci1gr8bE1PEjXHZVAAVWGXa14X0V6zmkDCbHX8EEs
qCE3awmGH8vnHQCHCFr/a+SNbbK8yd/SCC1jFMcIwry7CIHqXWa4/K14YiCeahkp
GrqYq2BHw9oA0fp6qKH91WQP8QD7Av2wMyIJf5pSn6uDVltPY8ZNwFGoaNw/LWr0
DPrrWP7W37KiihgWAig7LiNd05icJz1MVv40jhRvuS6oV1j6hw/aUuCkuZQUEdSq
CecI2OFXJiPVKzXvXgX5IwJ214oIzPxmKkVp7qfk88CuS2atxddlMSuv/OkGgZam
bhA4NDDHokyrzvP5VKGCNTrA6d1TEdJWe1q7v7HzcxqvZ4z2eGaTNknZ7wLA92pY
5m4hlx0goxDiympQPE2Il/7/1W5DnUjM9Lrv6jdOsj9sr61HFgxUiX8oYMxvfk6N
u2hWi1unhjkAg7P8sOxH6ADcD92ZcmTlBAQodeUjUg/z8AJm923U3UACrYyXTiAJ
Je8RftB3p5vrl12UmR4KxQnNf+DDinD0yfNu7IA10as8jMC6UuiuyQ1gruUg1ERz
c1FCzeWgTqLXFbDJi2kEla7caY6Mw7+5rgabZiXzgYpupxMhTRL9RYewSfF1d/bG
84na2dhy9+YxZitVh0LwEHmcrxsew+PQ6jU8oXverl2cYn1vTjUZ3SEV3mne1spx
c40+G8vs888mAFBUHKTBclAWfxvn9KevboCUSR/MM4B9/WiTzURxOTIVA36XnKY8
qzY4cmUVUF3suEmiMqj568iEKf8RIX2iFN6mePfcxSSv2/mP1LMrjbPxk9DV8cTC
ZKZQV8WLsGiGX4VRtLphPKR+A+ykC78Xk3cnJxHgoHn/4oSZHS14MHWo+bi0ewBE
/E0TFV49UWQ5liPleQjC8IjSrWKK4NzTItanh3gik7GHKagBON32pQjOj6UkQHYk
1JMyXnXclh4y7RRdK+sAKLxz8SNgwkRHWJ2mAeCcdPU093c4X14Pd0ye+GWeaLjj
Vvts5mclrvQeDgASXvFUz31nKoteBthOEqIwRK2f9kcEPUu8sBgOIYOAjQZdb6KM
JiMCaUwnnHAoNQFcYED752tFFfhAWFTS1XOhHczfHsHx9yGZV3/v7LvN+3sw3dTc
YSB7AifqeSDHYNSmehlmfLLS84LpyfHv8VXhgTZs4ir3Q3QrAwIBA0MsGNn9B8qV
EkAWHP6R8tNuaQ33qVPKUnf9elv5m02otbSfHIy44NM/jD0eICGEe1j35dwhA0Tm
gnyPYjDY4XAGjdAg5AH+QW4b7R0aEF6yBFKB48jE1vMe4jfIx/f4BpPh0QESRYYx
RTq7TnCvPdrQyo9iJLbpbnw3VNhjdR3RRZlc5wkzF+ZhCIGuSTvuhltnOOsCzPgv
nScfESKCYVDhCGoto+ZXCGyKMH2icWPAUAxi9qndZ4n4f9Zj515SvGg8+YaUS877
qtW1v3Ck7nvVaI8QXBD27zrPjDnjCH572RTlm7F7JMELGYDy15STI/OYXJOBcfam
swRdzxzxjbyBNQss5SfqGmoD4bpbd0u71KcQjqonXdAoIAIWOlfv0/R26SG54Bkf
UIJ/GIQ68Pc164SFFXHjx44PB3hbxHvIz42qWffkNEoTs2HRy3egOpHnz11z5Ww9
hsWZxpikQ1BAuX6suwrDlcW+nHNtGEVEP03DJQesnGRKRDUGWZrn/50nEDZnUoJr
jZ9NVNgnJvPHzisZIoHEZTT4ziUOHafmxOCTuvorNwSNFv8aBpUmZZnza87GK3GH
6MuZffEIN7z8jil6bZWZnv1Lr2wKY80Y5Fc6A5/mhEO+4TaEggNF3xhRmXxgO9y8
cpumIqR4+z1fGN5Pg6dRr/3H/yjrKhMsfkJG+qMmhaOER3xtKS3dCh/fFO/4Gmue
Fs7T2T61/kT6+s/zXZdTemTGl8q2V5Jwhy4x7uEBMjayVTXbQeEWFCSSxYXWH+rx
0mJK1IoEopad8UY2uWrwMeE2XJrAZkHXbKe47cOKvR8r5tHqyXbyMpKPcwKCwuoQ
pB2mlIq2jKWksZvISwnFmguQsiIBSLkM6bKu6fHcp+0FCvOewDkSebuCBrbIJUj2
B0SbmTMuq3JOFdBz29PpfhmIUoF1jty2HDAd0XAa8zOCnarwzl9ZR5xppc0PuLCg
3I85FjsCtxcTEB3ldjgHjHX1/JVwMzK9HMtTU9edEBE13qhzcTXi6HYGF/QCA3bK
6ENYFnoZoxsJdfu/9ZlmcHW0JfZjApwyjECaCmER04NNqN3vG4ozBfNcPeS+rPA2
G4sjnUCtIlbBIANKrcvod8lyG+M86MWPVp0VB7kl1dTT/cpaSVTe7yu76mtj9WL9
pPINk+7kj2iYorOebPx1ZH4sYOHHQuKpGvEttX1J9v4gSo+i0tLE86LPZ1oZVk+H
6tlQIxgAiaSb6wIKLJCiijXzxJthjwy4U5Grc0d+NKL2BYj2JZThF/9Y9UXgFTz3
o1WtFVWSBhWpigN8hfU8JUfNRIKcm3Jy36owuCkd6vKvWxLIWpsS/a8zfkMfnOWB
N++NfTsLOQXjzoB8sZnUYMyB+TCL6jjuOeHzo8OJqKsdaUK11ud9JyaSchYOG3Bq
68t7/1YgqbkLbkxFp4cxGYdB5DKijkCHcWHny48SqrE11omEfDhNyyQEx5OUcJPn
0lvOmnpW81zY/hREy/gRZFwS2FRltH+JAskuxTrg1kdKqZGzG5k8/hybLpwrqEJD
qrYIdHYr5lvsrfvi+otH69nWEdOgzObSlbkJ8u4TKaLGhQkdZUZyew6o7b/T2cLN
KLSxOfKetR/43wLEGe+iXTY7OvONzDjAYf6iN4acwu0JOp9mJG/QR3O20DB3n7F9
BU5Kq9NueI3X1Hamz7FEg/EJjswWK5vhf/g2u+Bn9pj56qmn4twIx8k+lSisWICl
HoX9wSaWi5nwcc2NTzfmk2UMLxN79lmKx+Gsd6vtVxTG31UjI0+27xzM2FgKcVD5
xbOvQneW3lrGuE9qNwA67u4w3ZX9K7t/dQCVi6HOAwxgbkzBqyEJX3PZxtHxih6m
+KoW4X5WgFY8fe6Zx0LmFBUzLVFf1SoSeNGRX7PRPLL+OcrXpuFZ5Wghz6L5RIQq
F7hAtk9ZTOVJpw7+5Nt8HpGmObYZw/qi4sy4XOPOa66zn191CkGjbpE0B6KjzsJM
YuwarbnPq9i+OqIh0Is7JHAcA142/0pH9hC6y7bGl2jxZ7agK6oHxpQ2Y2rFPf2L
07yQT205oEK/KOd6IvhyHNV1hHTqyD4uhzbfZbfgLKS7bRrJg7vPF+brFWIo0cS7
2pXU8x0udpc0imm8DnYn7G5fBquHpTRYzaoMyOd3v4ZD4FqpfQsDvW+l6mMGwR7i
IT9Azyx/USPHHIK60sooQjBlWDAS5TLHc9niqrbRJQQMxenIkqzc6G9fJX7pSnmH
rkgZ7xMJLNvrfnR3pLi9oZ15XfGfwqNMSbvxt1dH8UkIBxA6SjsJhLnyma+b9TcS
+St/8u6t3EHz8gZZNCfsi36UQ0mOvswoBgcGrm4y9AYoo31ahg1Q0lTiZkuaywQ4
cyx8K8d4BfkFHxii2KNf5Mr9PepMueKSveoVidDBH+JpJYi49a65L7RaStBv+fcO
bX65FBgpbMxw4wkMGm3ql9W7FSAk1mcKUynRqtfY36k6fE8/I+982brWpAFBYNP6
kOizVsXfZD04j4fyP5FzphLtkAt+/LkvbjKDCPR9R2F69oVU3twUgaeoVCX/frm1
1KNn+1ryks+4tv6tkT+nIa1bEJw/PHaLlkAX6QRDUAW3g1DJwHi82MV2OX248xko
UvL0a9ga0fi3Zs2PjNmvFvLq/+Lf3pUIiWSKdqe5nW8HzcW2IqI+6m+wnlyZMmbz
qp76nGnKCBJ5GexvG9B1I3I9kU4TTR50Bj1ALe9lesG5zBqt/EkEv3CUD/qiuuhL
GidlyVIItJzQg1Ekx8/f5MvntAW1ZwfSE2m7BqBM/7jb8eMZfI99myiawJRn9GjW
8uE92nI6DputjjUmjIc1RYgsihK3O9GwPDSk8hpL8ZYSfNuKamvVCS8bgBAKynvS
axDYF3s0cDzayfDBVFWjYwF5mtm7eko/jhrOaRngyRPEHvse8JWPwabiNB22cvb6
LBC5SGy9TerwGNm8XywCHFCNsqT/2SLvZ+V/csxPa8xyKc21kkFULcsuySuIMi/u
2+35NbaW4uZuRw1vu2zYFUQxZOh9ggH0QWS49rgIRoxXtE7AasWq6GEHbzbESgXC
oU8UTQof7McNYO/wH3O7dMmXgT5ppQdTRrKK5q2PbD78VmaR7A/YAsbWqpCfGdPR
ykGdKgryZNboDkCb6Ne4yiTdKwTd2mP6aMrv2RQvaDgEPGNpBc0FaGhF/eP97pL6
JosdBxD+hQ98uU/SuUgYcpJjFFCXPCDw9qDUiYOm9sosWSV5GabirJJDuLkT4oRX
lkhf8PBGNyga5PC7ebEXjQcHSTjQd0bdRjmt2mIr/lFy8HMWikBrMhJjbwAuel8+
UshwdpvPn7/lu9N6Mv4iSNMxDpIRJBMxUgVYxQ+c8S/YMYeqIiuuqUSAaDkTzQUN
Toh2gXL9yJix8+phb/tqMc7fG57uFvUglV3QGDwSdSiokFFnBaxn6BFW5Zb1zv8X
BCJsvbx4Sf1ta1mwpoK+/OGGU/Qid4yJojgP94jPKM10L1FhwJk9g/7+CJfeL650
emMIIQdSrsl4bMpBbptJtmd/7CC/3jIMbjmSu4XYAAWnN+rlRtUcSgAS2ZNDu3H/
70yv9FO/TKW+sDoh+vLePwY5O5NxFIzYOhVKRKvAxkLJcb7DeAdsxa4xAKQ3PuIG
MGUr2moWAUR3d5mnONPPnEV5/vRq6NlWaSFtTLALlEkA2dbYyK42w+aKEu2x5oKa
0VT5pUq0V7HebCrK/ugExmplSknURwhlKnFHlqC8F7r6NNvvT2CQ0z8qE3MmR26F
0NVfU0Bj0gAKca9ouf3IfBXLPUczLe+xc2pwjVcU5WR5mtMafpGXac2JHbLoGYj+
2i6kT4OtHbracTmwhM/Nx9QpCHLPnW1ShEQWbIPL+baao2+9We++2aK5pCnQ6yHE
7UYSMVZfpJNTFOocQJ89t077Yu2IYM604RpmjIlcjnJWfpexjcUgAuEt5y72SflA
ycAY/4rDR0fjn3xYjKPmZFZWf6TZXAP1oFcVyKLm2EE=
`pragma protect end_protected
