// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KjdM0izMH/T5c2JM1XJNF15GtU8+XmHN/hYihtVcjlrjRBg8j2OIh1oHG/71unfy
ngEcNQUU5yTeCI83QWhO8Cq1w7mLGDRhnkFt0vBjq6onQDKWAxk+Lx83wWkkAtYn
IpKcrX6SJGq4t+xWZdE6icYw2ATERoiSFhE+5X3vauY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3120)
zJkKW+1SVXwyGQUW/2eQwSkWHQhbyd2wGJyUFuuZcE0ewJLZgFbrppvkLilSTRF0
CVj9Rw0BYsefyohpITUOZENexDDC8S+/2a3ODf9/YNcZOqZB4XUZAFqoEM/8s0PO
ScBQZ9JMs0EP7RxMpmn91pOCcbc8ENJT2aZPOPKuqp8eJs+BsAWSxhDjAoWOyi6a
D8F+C2L34qtGqb4C1jOA3TxlxD5zs1TnGLWIe/NFXlq4c+V/tB5eUeRUwcz9d8+A
LGFlcXDoLvPrgzMnXz2jUkHN/v+Hh1IH9BtDL36dLn1nZsEl/C4I9HdWatAvBWy4
fC6me654iHaHMnUU6BV8R2gt0fZodH7Z5+SeqZLTPtFTXlw0P3hGvaYsNO0HTcDy
2CKxJQ/SbzeZFx6K9rObnqTosEpGla8nUhc1OjW4dQh0XDI3ZxLpCq2Vto6xaJ3g
DL2Yjo6fSiO9wBIoo87yYjfuPXBCpWhljQ05mqpYBOLh6WL1rTnKY804le+uW3Wn
T89LMYnMebZO95xf7ygiECOO4ijtZTDnJxBAiD2tir4045T1gWk2EECIO2bdiZHw
4QvohKnI92oV73xgdc5V3jjqifuOLnI5CAwxDoUZUbK4CqoWM1olzvAvKKv9CIKO
pr+nUxrA/9bgygPhdMEnM73dnbTyc4T4wF/0OH/S4qZcJIw8y/bP7hbamjxDYXvB
6K9JDN+JvGaROgudBGhEDP6uN8G7W1eiPa5ovUaOVlVe8YzLfmfTaQ7SXP03ZSVs
m+biwKfKkkk7x5tesr80uHdQaOiyrKn9zSubwsmC2A9/f9GVQ6YgkwdU06/2ZPXJ
RQlv+xbX4yAiasOF6yvd9tk0ySDRFuxb/WMlgRZ96LciwGT9tV8SKL15wMG56Z28
zfchag2w2Yj1PwVrg/2AYkTmsSiZ2+T82lJmBjrdZOfgjdsy+ey+f+6/Y7qypy1k
CazZFtEpXSm/1frIgoZ1M6Zbp6JHKxAU2ZJUbWjmwABUdgsmg4HZZFiqXg0Ykz8k
HcrIyhSRIHDZ4geCnyToo1DCI/pYm/JmldCqCLuKUz934VT/qoVArCpwbYwqURat
FFuid34BB5iSt+84TkZkHbTP3ItHNQ3wjDOChggW09Brnu8LfkFJVkbiVgWtbtJm
JFjcRvkMq2T8IMqK+WIMjBh9HYchfKRI13I6rBLm1JZfKO76xCk9BIhh25n0oOFP
wKnzU5pYhsEccPu/D7ryPubUKIsalCP1dQ1fKDN/pjLlPsiSGEeQWQGRZ5Z6AZpy
EKXacmopH04EjrqlaNiclArppgZOm7gzEQVfqoAiwMlKFRHkkJI/hpr07bf2XJwl
AmTJTSfzStbz0z/qs7nJ2pl34a5r2mAsaODvdSmZkQVdDYEoQRP8XhZgZ8NIigsg
7DnhkHombpCCgZyPCOSLpnO8D4s2AYPh6/uqerSj8oc7p8J89vLLiksZvHLXIX3h
LHs4bt8Z06drzd0aAkW7ZYK3k6xJuTtxN8987JJHvXGpDIKYEhvUsnpHMpUiXzmM
gcMpqrpAAj2oRSQA4cRpo+xFIBKEk8zWi0Q+ha4VdUq3KVEFzzO9curDtsA7Ar8y
B+YfmGKSOIWVhKbQPB86cTvqH4SNxFUwDzhKpXAlFG/hx5f+oiXO4A/DmPBSTrsd
sW976HaSam8olkOLyXpr267Gi6QssxEe1gbRnRJo4FPBZ7nD3Jda8huq4ww5gsFb
qEuwPuixO67DbK3P9zPe/8VjnMr2eZGwz14d5fruoQoio3rc/+q2aepSM46MZQZP
ZxxflwHyXnm7cpVG6+djXmIgUjSQ+WF167Ajhrf5D1gakL5bB8L7TklUUfksFyAR
kOZ53au34tJmLX4L/cvnHKhbO9x2ZwxMJv1Hr/yYLyWSRZX8pCTT5IRU7TjucZbZ
MxKytt3SsCUvuovLxRQPfZqixj+IxY2LfVah92nEAi7pie+u9NsJdgPBKOdxfdTo
RTBpxtOVh1MbktxcrXi7T00QuQsY2BTo1QvgDCaORqAGZfveygBSZjrW9E7PPPhX
AJwNEJ6jcPUIZW4a+ov3EDVfAWXxgAQ9neCEULcju6X1G90u2j8msOjEG7RMmECz
MdGa/JcLcDyWALl9734e9zHItaziM85LFrGpCzuy8hyDSN16BKqxaCe+OZxcWhb3
4qZf/Q++SXANMsHw+PK4UT4ngBPwpK2Lh4ggVm35E38EdHEhH+rCTwYUHs9LFhY1
X05T49ppAII5cyVtYLJg5fXhdFBNTkYXFqNZ2THt4Nd5KDfM+AHtgE8qCQCar9Ow
8vF7PNtTbiDFO+aahfn6jXpZs6kLncMJaBl5Tnsin4Bz0kUE1vH08gQa45TeXPwE
xcTWBJKXZmz8INrkIk4Mq/7RUaSig3r5gpL+lO+B8vwTwaRgq60pb3S2u2udJ0jP
D6zoDC0LEBQhpAMX2d6YdwRn8TLRdE5hmWIpTvOW3Av1tZ4CJEzdyGvTsR25uqKK
JJ4m+0BchE23Kqn3tdtOaDMe4PBhZwSgxdwDajvmEVxxefkTXXKCrL+m6zSeeYiV
bAMp8i2Op+vlXpYZMe3CUh3XPNkemOMsYgZOCKbDGk8y0vGnVpwb04sWn2EorWQN
jv3nb3X5jZ7Q61J6JB8mZvMcn7nlXKhF2v2ml+jcmyeQBq4toHvkUhM7zAHr/0nV
7KQADobOSGyJnmhIOJMWERib98q+Xn3Y/G7zlSldhuuKkxIntZ5mlHhcodRwC3Xc
nmF0N8QxPBlU+Nd22PaxEPXLBOC0jW6n+gvMor2WTWv+NW4hIT06LAi4zwtlgN29
+cs06D80zxdpFvmV32rX6P7n1rLWIX3Uczjv0l5WySWgcLwqWA9LsE9zrS/MrUX5
mouwaCXjf/3sxzwhcWfZquVmarLuvaKfm30Yp2N6pxdIx6DcTafcLibMKxcU2U8M
TtZNcf/3Z8uGG4BqFwMjSkznXX18AktTnXaSmofjPlACS7sMm50bYKo2iF8znz7/
+sjC3rY+z4uohnRCNgkVmM1excStAaAzvRgaKdWzi/SfbSloTyJNljOWE/7sipvN
B3Ya86vK5C9kXuzqQY6niSpTtr8PrnL/YGN8E0Rv8Vy1RZTKjgDqwjy/aPl6HIOs
dYHZs0UQc4K5+OWGLDnrtylAL4h52aWDKiRCbBIopc8T5LCmF/6OpsIJ26Boz74s
d6BWWOEqr02OgCS8DJXE7mrZ2m0dd1yQ7JhVNy0D/3AO810d6kzA4yjQPp0xfp2i
J7WT01LrmwFCi5Dj8JvzlYwBR8s75nSyF/9e1VUX0le22cKvKp1QTG2cgst2NHqx
JgW2fPPunnl0CIJ85VFcIGw1jPvoItiRwzMggLtt7yYwijP3C+MscnrDz9t0I2Pk
WSxwCE2z3Gr/TQuGy1qNxDlURB3ftwgrjb5MNFU47m+1Egxh+serrj6i4femmvgM
itafsldOFb6bUUyxQjlZJheZ1s0i6YeoLBL77Gh6hfOlb4+WcDbFDZiOIQ+pDRbq
E0Pu9WgJyX29QOrV8pnnZUZWqq9FpOBWE7vfT+3bYg5W2EkmduFu18t/YqdBbQDS
+hEE73201tPRrRX2MBQQhIc+T7ykqEBhr6s4FoNp7KFNSxq6gEI6J8anEX+uGxXc
7Vyd4/CvOTXxUh2DzwMl69I9G37Y2g4IuY0fpDCmBO2B+XZL1aG2XgPlp5EJyi15
H4zh/kYYCGhoZlGtxsG6KixTcLizAUQkjXZi8YscXy74HmaP4CutiTIFcusjCRWD
5bDAUD0vEbUAcDuVeBFVGfygqIp5YFhUwex9ygUAwhVEcUfvmhDswc31Gb8zL9Wd
IZ/4ejwXkxtn/PO4KTmYkiYBppNgH0YZO5ueLJEvXc/UQHADNvzvH7Yj+MubVJQ4
Vx28itzSbT04Fv24uaplF0+P6z+DLGQ4gTJ0WtbsJkL6eUDbVWyLqSHtCKO/BhxJ
ZuqJaFVGvqoKYhaMw1vD6EkxoXnnWfPmHIsDS9JkuDHL7tsNRwj2RjylGUogDR40
h+L/6XKKkMvAMO1PsQMbRLMuWHWdXphdpNSaL1L8llsjSBPCj4ioa7xYPMT1nNg/
31l/NxJL1vXH75bRmPrf6cxZkP5keFfvR/U2n80SPhu9rIrLrcI8HeLcwa6mueNO
`pragma protect end_protected
