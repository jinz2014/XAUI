// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hDm/Epe5UodquO+7qd6qC6fYWY9TkqW5WKNzp+Qxdh6PHOct4lRCwC4+7xn5f6Yw
SwjyY+MKjfFBggxyul+CWyJry9RL8LqQ/GBOdmzolQRYT0hfPDbHnxypB4cWSFBK
M8GleuOBDHI9ZIwLKJaZ1h9n9xg2xpH0+ru6KHXQNVU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28144)
/e1pPrT42VYZAYCGVVXcp/TpTJkr78iBD6UZamyL5XZDkGcHuPWYjq65wqvUzros
NFu8Zbzo3YPaWp9FaIio5pomhbo6EfMQd6/wdGoRJ0C8sHLlep+VL0ZEd+6Nsrfu
kTII6P7cBRpTWT8JLFK4u7uudK1FIT8xpHg4VeBSae1KF4keB5ZTIBlZGjZadDUl
OX6lvLA3PKFWEip3mUZQ7W3hzya4XZu1vD2N0I/rfFaRt+V/JbLz68ukRAWhcyhu
uejx8hP72FIjAuvWYFl1fTcbpLVvLWq6241F2hwipDjch9SRm5lUQYKdrCmnidnq
MihbG4UKyKfXp/8O+FdEd6FmnujNRyvDGX5z7X6v6I8lIwdrDUTFt8BCZMAySuj9
be0I1kZAm4npkFqS+1FWQVUpicddfb8eSdLOGGiGRL7C5tJa14TiOMug/87xWs0N
pEXZPm2vW3jqTOh8UJw1WiLXwtRjCdMTqCtSsDRmNnCAslRfpx8YXz8dfBktNpVj
lErOfYt08dilhilUkvl0vXCKjz/kkGkQn2Tbn6MHJlriHJQzi9VFWfpNV+/wVTW6
dHBo9y6I3fn5l0uYd8Vf0JB2guVVLEDCPN2zqEJ0euDNXm8q/zcCi9rluIZQxddL
jwMwR6uvTdhw35SXLe5oogbIRgv4ne1Sh8boSouC9xKwFqwK2FfNgTyZV5BLVmwZ
E6gpFmcgvfzJI4KiYuBF5hUOx4E03I8yw5lv5QKGFLNGL5DzGnkT8f8GKw6ebnA3
MfGhNv2UBsWl+G09rMJLuOcOILeNrfdGWK9qNPxSE1n0tvc/XyAnzcxq86ZmNHXo
H1w9sfFSVhMJ+8FkxD9oDhoFjGpjIHNPLpkTCfYEMsRAh7YaTYj2lpxeJB4Qo93C
sUWgji0RSv49a137s0lRU2QiR1w0FrwiE/8mLyYGAmUAH67YSLBfarL/1JG+S6Kc
QYPjGK/hq17UyjJL3JZTBc2s8LSgNELZDsqJ9YVO8oVYxd1idMP2XAEOZbD+y+X/
bOxhgw910MC/P1x0gaL88dt6OJlL/U5UbbwisE4Oi8XdaNgy6PJE8JSF15vkWeLV
drPOz0LlJFaAZ8AkmaNEKrwyEYSDPDor85/qMl93IiFN8ppRaIif1nuoBy10CRGb
jRdAp3uEXiuAxBx8K0YHuvcHG+tt1cW9+Rb5X2+GdH5Uc5fIpXgN9Tqo8E+nINYK
REEGyfRS+k73LrRs1Hp52h3jO8ZN4SgSAzGQzagKSfMR7S8nJyq04eRfxKY4kWw5
aCyW3UkGyX1p1ixlQ/mKOZSa37/EG+SI+i4CREverJePzxyR9/EaU10xU92H7wDt
IEfBA6cG2BdppNx2jowlTrrof6d8GXDBZY+SMd0dD8JVK9jb3g94Z1f1eYXeweOI
V4PgMrb5VFUQKRp7G5Fn5er3BtnLUDN/UXtenyIrtat7+2Pwfg1Et79ZUDRB1Uqb
447ediDzQpcM7UBe93rHI6d/ZLdHyEu6RMy2DimRE38BOjEsefWw5tlgI4qCofbS
A3GFVetVG70PeHFFT99vMxtd0kvYrBK69kuksiOB5XdXEJiyxzkZaijClIo86lIm
Hagdf1F7eV98o9K5/jcNeiNbkArZdC286MChESqvIH/ycvqR8MsnnaD5uZMJP/wq
8eD/r9IhUOu2lU9x6NRK5MqUks+k7zx2zXay8X4NBxF7GQ/VAtsX35Ag2J3cuAky
1yHNn+4Z6MQSSArCJNdCGNosjgP9f3n4jq5jGIAA864THND27ptlJGF9v738tmq+
zMIdECjCEsjpCjdgTEJfhdObzRWjDXPyZiZtlVGA70aAcdxY9f+TgDo1nFVWuP4X
IZGPrRhglbIPI5m6htEBkaZWVFV2vo3n6oDD/FPJz5z08/Obj0VsEWBc7CCijuEf
nC/bZXseOXaY5KGhXPBK+QYNosuZH0Hc7OQbBClLaMnaTV38Iuv+jJiHV4l/sfsB
tT7TYc4KsDpi9Jxq2qTx3+YqSF6T1EcvHUt2mqkfZy8gwsilZT4mx5OlztFairy2
rARKjky5FzRai8LcTlD/yHzdycGRiQK+IVjSHbxuLGIh63R29th7WUUHMiVJl3Nm
ZYCMuMM2ZTNYTBlLykcSyAUQMiW94DPgVG6pCEHzDdoub9n+GT90sBXYOPYab9nZ
yXyBFSB44dSJjgpu/44hhwu7nMQ8NnOaMPTEjaOBu2Z9pFJo3nuxcp+FaU9VWQSS
zj9I7W13sC6ltHWdXrq0dyj+vvNWy1cNoxoPUoQIQYw+rQo37itXidB8P6MYPZi3
w+LS+QiFyB3aepYjhUToaCm8N+qZNZlkwEIM4UeslL/XRzgUqSPEVjl18Abos82p
4giElIgxw+FQbjEOL3c3lasxtxBjBVT4Jf6EK8hRAyUgEHHEIWyxW48iBJ0Rvqnt
sgQ5Ngoc4qfNEhaMbXpfGwkaNY4iSabldSiYOj2PrO8Dm06xIg+RFKY03DYQZ0xz
ovjK46qwp3JVYAjVyymsQrcAWbmOvWsKnjkwvRNS6AuoGCsfEyo/Z/i/MvKoDIuE
SHQvN1GzsMKWqrtpPH3Gld0BvxUL787cEa05grfXjNAAtVFWf4U/ydp3T65jMmo0
EApAxJBnEh7Eghy3NoA1OhOJks7B+mMTS7ChEZIToFbr/uY1YuWnwC9ZN09+b7PJ
c2LYlmRMtRzhnG+PnDbY8oz6gJoYBSrvvZLVUBDMqKDt4xSPttViLIUNRo6jaEZP
TMBsIc/vGSo5K3J+EMHRhPEGrCq1P1ruHyftEQ7djLbvWN/FfDZzvxNm7lkhbXEe
Dss2AtqNXtyaZHsSQk1lsFKxDh+ejRXA8enm1syoKMjFCYUtYlbtt1409Xgf4m59
jk6ZAZdP3DKg2HYOyOCXkEmhigkkxKB0kaGTMiKFFMl88KxPg67XwxpzPMq4lFTM
AhuWxzpu9WUEtIPr3jkxz4VyRpzyFEjF/aMU7MtevbyAKqehmNrSX5HIbI3ncc80
Wzk3xv5K57+xqBjFg2pV/naF7TD1C36j87c5uXaT816WNk/YEFBspaujxWlKvhAC
zzVsDkoPp8+nqcnhxbUl1C3w2wTM/6V3FDndX4JTnTFn+Jwv2Q+QaNEnqLv5dnVc
V0JBu9uab0rtLLg1qvAk1WmxTd09fLiuuyRScZrQQgp6C11MNY5sZIYJLBcxdWrM
kUWR6HDrAXNQklHKa3TZQL/pyMUU6gX+jlYdJR3mqAwd6tV3b7l1Sfd5u7pPM+dU
9AnfMtvzsgTpyFuGsmITkqZwiNCWVyiNN/ju1pHzkxqqp4pDSqd15Xn1Mngw3Ema
vR+2vhsmIbjETTZuK2/cP2vgFhtfiNk8jvwUBXb8V+M45YmHW6r7APGWsy+bFWOY
D0I8KmTlHrh65c1vytsdfpWPR+wWTP+TfNio1U15Bvd/AgHTaZbcqC5/IWpE/R0b
BPo8avBZYyXLdZq+juPHpYZ8UOVOPZDaAM1SXWGFaBh1k7PC9b9loTuJACzd/qQF
sAr2KE2/3LYKTSSmB6TQf1AYE0AUarvAi4NEqX9VI00gwslIJ6qRsi/LQp62BO2p
iQ1zjTDI8RzRF/PW78ZF2MfA6snHbx1ulQ+AjTOG77DkOr9IpOaoRSr/lRMOisiD
e12eO78Sm14ZoqRkSQdv/pvjdgC6wje67RLhhwll+9Q0vuUNmQpgEXIFtyPh7C7E
tS/nOigR3LHirc7x/hU1E2gIEBC+YWlg9IsTM7MdU8kXkw3HwZLnIjkCRl2/TLcB
fRsWtmIPB9+SiokqFrk3Ca5oRAtV3j8++cfnlyJazcm0ufSwsqWvN5hBY14gP1xn
P331a0ZGDDRwwLQFb2Gwpxy86wfwr0gTuAmR2shC34H0OkmkRVA4W9pj5/oWn5kd
aaJjkuLL9EFgt+HrrRrLjw0omuXaMSYajg0MldmXu88oPCqXnvXOtQ0cVcYfLTaH
0as9REbosGnxI7ECQZ3EuT1H+qYWW7/fVBR9t96lezLds60wOFZy9IaGKK93qGOf
1PjdWdaRlxN71uNLtLL5mcFI3+HmSWNUEMZhTbaUX8eeq3dfFWbg8uHTjRmpYfGq
UWOs0XHdm0Wbt+2PELKqfSwESXGZ+hLcCPJ60GNxuWPiSXUCkK6mW7WBECrYgRe9
fdN/uJCo7QCJgKRf/5w/i7Y2jDuelHCu1cNxoF+gobmtqzd1lOTr4DYxMXI4rHzr
ef22xQT5QfCLeN5JWyjXQKgxasdGnaOuHPjSP1d3NRYEyqyOYDf/xX+8XIAy4FSU
lsTzyDnC3GI6LfIfRieCBBrlNVDncGhpD/HC9HEuC1zYckTWL0zeJZt9OiD189/y
TjidsdpqLZf/3+9Xb9VuB/mQFfTwidoyvlPxAxG1jQVa8SC+pXRkibne6P1Q6J9l
7sonGL6hsSlikkbeVRRX6lubjaB/FxPllwmPPyKKaAI0f7ONXrkGBDMyRiTW16Tl
UnYtThuCOfJkrVb92WCxcBsOVsfTxCJuK+T1TqVwdG7blFBWOL+iskYaQzpLl4uH
osgKstLpF2RduPndKe+ID9bLne+VdBjuVIJIx4zFdshT76V/IAoauwsWA0P6jK3L
gdzeuT3VoA/9ZhbTmoaVOb/nOOwLx+Ig1MyGKvenrjwF8ThTe4V+rUlGKwgQqzIC
WsHBB20cxU9eCJzeYUxufVGz+FpunEY3iP0E/0AbKVlCshAOqrA5OuQz00tK/Xj9
d6zAgWExXz9bh9HG5E6Fi7wBIQS3LNg/AhBypW3NehF311Xg83WkK6c63YUYaN4F
Q5/X3W/zzjSmT3q4Bv2j4ePyCVXAO0atOSdP9iCc7kxr9GR722kIRyQe10ZYuzW3
nSF1cjjfNSQF/i1yCvPVmPuAkgpL+YcyatayPaygs+qBLjFyoNvoJKgkYYSOLeJT
Isu659XtwrCO57IYRcgFHtbzlY6KrU0/vxCleN9Y3Do1wIF9aPBQi0fOsF1oIZy9
E/lJSkZxrKBYCeqhMBigCX9Ia91HaFbQFIIU3ksIN8GY6tPsSvxba+bfaZtosowb
dw9EwvIQKIQoATWkNKsRkKvSGX++RtdUS7Ky5WK/AyCb/gKwkQH57YOpUT+JNM5/
lcDiOLnMdzHmcPOCoY25SbBegA3ETxTVSjiYJRR3U3Rpk2iNY+/sgCWoMrDkxHIA
4vdzbZ9NukkCquX95U4dhd12pEpHxSuEYP9Th+LHkubw26x20CkT+4qzTX64CKXf
9GzOvhQZOGXqPtWABko0rQqyVoSB7TpfdzZyza3K92rX/Pfz6m3YQXe9ke2RLpn2
DeUs5oT/PeslxArUXSJGwkxntL+EhmwNoJBC+rx1wwSHke8FDnox+QeQa+AXsr5f
xFv6vdeTF63Y+kYIFyIDXwjl+m0I3k4Kt9T85/GxR0AJUWFbbe8zy3zMVcLyV7V3
YwJjJS63cUgUYA65pbiP70bNU13JZQ9jBmiuynICzRNcZEtoXpfpLXicSEkTLB6f
Td2i2LebOu/C68nwofX4jdrJ0RpEP6IkM3lK6wu7c/CP4eFbFJkoMms+vSZ7GfCV
OeObQ1EynL+cYaVECrj0aske2yx/x70Lg9amp0uNnoPSoNjo0ZgO5bZ42Dlybhde
fz+8U+RI1JD+l9B1Ctrj99hkPctbZdai+5asyZfilMj47GUQ8EtSJjzXlwe46mW6
cVwoTs0zZtLyvyya9fd3dGg/udsBMs+ahPctTs9zcV0DYgGP/ZI3fEKggJfAh7Gu
hJ1QMxaTHkQPUaCpb1Cm4tukNqO+eFgH4rXEXlAHvn9YLQmcOjAvb5Ev1U22KX5i
NLB7saP9B68mtfajzM047XzaQwOelnW8CxdW8JBVpFPw8nB/QASILRlVFLn/YgmL
NTniAdILOy0NWKIcStGVXg0VkVF1mSNLPGlr04fkPQ4T2mNanNI2CWW4uuTyG4uJ
gfDNrlKSQnM142ifLMIi6nG6hg15J2tFD+pcKhZ5JKVmFK9uKIJKa63v2uEtpxKG
pA/nvZLgcVCoNCoTahhdPubvCftJvoWIuic7z2x1PyQJ3y+47rOAW6ukgTtDiNyu
oF5DbkZzDwCW+4h1awFZmJk1cy3lo/iWJ7uRPCBKWphiHhLHTbC5KfTS4Uy6uLjl
8D/k2YzctQPi/5RJIxch//SRxMGENSGEeP7OsKaHhdojBY1UPn4AKHWwVgivUVpa
nnUQbJqz4nhqIv9DBvdWaNqWTIBrZq9mWn+3+VCKyfMJ2pnDCtWLMqqY+FCm/7gi
c3sNclzilRycH7dOrEtu7HGYXDguD5s1ZIllJmhzzryRw1RsHdbBPxw70FE4/HTM
di5vQW+UZeceJLB8cA1HddSnfOIDcU18snXuduX1Eh85lhVV4he8bgmM7e7qQ/OW
esQzzkf7ESJxfVl54A6bvByWX3Fti6pnYsAWRttMHxPSCcupIKDOAdUDVcl90ekN
02Uj0Y55V/uI9MpuTL5xxcNgUCee8P5CuBSZCeJgsRcCqZRzjVzPe9c2rCMZbu+r
bVGMNZGvTuwmvXqc/BkHuY2dRELB86e+XaS86FG2RlqyM2K0u0LNMkCUiYtWXCgw
/qcgjZutj2t3yOkeAjzwZ47N1YisygAMZo4ACzeKee/e42ffuCqgvGRuFt4AmLJq
w9Zsq3jTubHToxeZI2RAL4+saRl8DAc6Ll2bCnAz12QNbVLKpAvHsS5VCCF+Bdty
Sv1gD4dB8QMDQ+Juabm05UK1X09jHK2RXBNczgM+lu12I2gknTfmHjeF1J10tWY9
mZOMerhsMaANpZ1dHebmNnJ3MioEzzKr8NPYpskJg/0L90okb/GVFnp43QdlLnB/
bXrycTpDaKpp02LPtR9A2VgvT3MGh9R4aLJRo7dD/tTW1pJWYng0z6OOogOmFw6O
9oReS4NKtxTzEkvFHYHmhXcpf8GC/D9F08gGbbYyU2Xfp7TKr3nkGhFTsSm5M7h6
BTzLfBpbAyebCPcam/jvxO4ab7xddA3RzyjLGkuBezwpSkgaXiDXqhocW+Aa9eH9
B8t+RS2UUdC7bSLWIf3sbCPX3GEEQaDanLsS322H3s1g60bEWrqLiN31BWS0j4eL
NNPyOCul6boJA9K0id2895nbD80v0jxEaxMOAYZJ4a9Ht2UdDfNHON2cWFLaoyoX
/pVckrdqiuK5o0awfmSc27jOLcXpTf2rx2cs+VhntOPDh15Qwe0bqEuHQfaq6C+b
JiXSCWm1Kdq7wJ97ZhOetVQezbHlgBeUTdty0X27WtiiIAdxv4kXKGTfp6uLoar5
59QUaOEwvhA4ZuuSfbHIYe8qcmxcu+5uotSq+REuwsprmk0HJUYso1Mg50sd45pc
fbanLwJacpXPka0e4EGs+QniByQz+yqaEqZW/ylXiBKj0Rre0cWDZCBb9O+zxhSE
oBJkTRbJCxYg/lneGc8yenozsVwfEaU3XKk3Mr9DUqEOnMVjcuUzaQgmlRs058jK
dZI+I52KGWTjJSirb+9J0sUmC58x/1gmKW48zWTYb9v7IPQhrLpPjy/wOHKwFdx8
3duZQ6/k4gSCUfkZ/kzURggiaHoc5aFe1ztF1SomCBZRP9+teMyuq5jmOYIFB7kg
SJPn8xy2pgsLSg4Cm/MhoV93asqJlU8IJFzZ1cZpvzKXMYsKiUz9uLLj6k48o4i9
M/GrTYF0YrRH73Eh51i2pKBhr0ATAzZPSpigDX4fzd8ZXcE0XVfrbKU1/SLl28VY
nFrAs6wrj0SKQDqldgMqjrQArkNNxsrUK1F/zofWIu2n2waGP3ECAWzmwQ4WIpmq
5bnZC0dv2ROs7TqFMckoqMvbFJI1MxnXXn7k1jexMxMB6ZPqubQ8MmVKiZfqEsmh
hyNLq95Cdrc7qFw7Ee7UVawWIcukHc9kqqyXUWKwH1vR0eMuD3cqkix+qnpo1E5W
p3IaPcCoctGX3wous78PqKBBC4E9oUMRDBle/2VS4VGRSQ4LUFX7N994UGR8sElL
xmfNmf+YAofXSlflBk4GQM2SuknT3Bfn8JHDRIENUpc7DvCa/vytOF+JLp4crwnx
sgM06Nf1R2eAXHgsYtV10ipXvbLbiiIqi0DKtJ9FNrGf1rMOaVzJ+Q+hSHHSWD1U
9MtRt31D6uE1DXV4/lEKthZ/9DfzdAQxJn3AlsUioZUZqfOBioqL2waqRIl9YFwB
KEVBnWA3ozcbKLDLozjGR19mDB12WBRvzfMgmkJxf1iXZaI0FmbOCPVOdad6QvQP
9mqzLKWIoH8dRQOBo2n/zRgxEqFgFHgV/u1VKwgkMI6YUNOgvA/uhKhMFZIbe0CL
3NLpQr0iwIajw4O2APbEeA8nhrpYtNw/pTvasmnXG9RvIORlG5DgfseCszv3sltj
9lysuBgquUJxSDxf1+FnSjumHSPKNw5179A3BcuKEgWb03JS8wGNNjhiMS52o9fH
Rw5UX5yy3T+hAtKn1C7yD8Oi0M1Q1yiG6ZmA2Sa/tkgIcIPG3hG7qAa+4ESZm/8e
FOYLutycf0g9Koa0fMCRM1n0eX42YT2GkchEy5nNSOgacO55vBvjOc5VGqlqnfXP
No4ipTwo0CuqElQ1LHb61AsY/8yHZUkMFZ1JsR4+rVLXA65atwachtUXorkN2FEn
wQDZ+h6zotttTmV4TQakd805F07iFrESlERhveeMeBbyEZ7u3UbtGbBq6hapqecY
ImcLZ8+gzsl6U2LpMBHSMvXKtzNGstrUBRtRDc7qQJnokw6ZWSxQHA5btjdSRFOq
8upiqbgpyNAzH6XFZLPiw6GOWgfmSyPG0tjWZZIR/+MG3fFkJAW67gwgA0hnL2Lu
JtQOcXCz3mGALW9NImNkcyTVQgxzMIouFdcZIX2Gm983WlJgLaCAOVkUJCNRgUFT
Y/QoKK/G385w3UTD4iHc9a2CSxHnnUVr9+elt8085ifm6os7idWjQd5k284/yYha
YSWWqsUSM1gsIZq9TmjTvubf0SCDlHhz7wLZ0EeOByKUfYuaPiNg8ze14NH9bHql
tbR0qj3zfKwU4VAWdkbFTSzfO+GgPsJrQjrfOFTW7Tib+8M35S2gX1HfQCywdMwM
IQrhueb95UKYkVRYFEyJXR8b02+WIjmtHxLDoI5YNlcjhFNUqtQWozg60VZ7n8dH
rW0WjiX2FA/EQOENsGfDHBWiWxNzPDj68J2MzCM6rxr/v+/HyuUg3NvAHjbcEeIK
EzAUsFDAu1qIfP1uk9v3Tu+moPVRA1hfYXba0r/90YRIb8EoCm2b/3rx+G0hf3eF
9DfTl5jNLIGcCXRjIq/9AEdeNutNxux2BujWED6EJ7D8HL+TBq4Xz9rYmIWqH63U
w87bgWpZMKIJpE08+JCpGnsvqODERPQ+5Q67QPZlJrjQHkuxQLg2kclj8cIf5Er4
Nu++gVFkeEvPXCrnDHpf5Pa1HPFEoteFrkM5tRa/DubnA0xEdgQvOOACCSK8qEPw
907gQF89l3GfQOVQe9EiKBsbDgNddCT8VUst52glUwZDcOt3AEFLUS8JMAFcCi0F
dbI2tcCWv2d54VXWNHlxoD3a48oR7xKfZCX79boiwqUFFKxSN02aIJBl0yMGeos+
S368WfJ37zCm2MBbgTTpENq3gWyB+V3i2AlC2rYUKeDIdCyJ0flrP9TXAaFwGLN8
uSH1qfgJhq9xaZsakFddwbkW/rJlxioYMq9hslcxzVIwB5AylkrPJ5tyxEcznn3l
pI9m58qGKpBJErPlTqSzlBDTA2RfJtu0OxM0Pg3TR5zRuonG8y4fAoXno4qpQAOt
1qRwiSmy0JPZ2keFK18ImwHYhE1Egu3fMhJ2hMcZTB+g2GgynYKuVR6TDMwcD/W6
F0zzl+FPZvBgshNdxKc9fn7KlgQ4fNxiSucLOW18kq7LDdQwa04rTWBakI5SeSF/
KV52Wcqv++MRuF7czaiyblbRngu+UlxqTMs6pJNC5rRv8ec0Ns1mVGF5oE747eNC
DcCOoGb7aAU7ZAnD+XRmjOS12DOzpCyz+0WYWWQv6/VUrJ/lUqgdmVjaoJpues4M
9hN1u7RdTHu3GgBbUdrVQZHIqvQYk/OEO+P/zoOD7ASnDgS64gnE2+RWtAs1CuTu
ydPhQsDIw8N7LwTeESb1LWcenvm/Sz71kixIZ/tQpbfbwYI2bnDES3mV8Gm/vzRh
yiMRnGOZxCDsu7mOa1/Rxgxlx0EqcV3QDSkWLuvUgX3ydvzcTQ0CGjcWJ7aP4fl6
+7pRZBTZmMUzsYkDC3CkB2qZ+nSusPwzzeyzw2nYrbAqjDkuFwnBp9JfoH/eAxXi
dWZflUQJzNsEjuyKgHo1ZQAfzUWloeJHf+82P9UtoYKhOHRgU5oc8pRIk7g6a/Dh
HHXxuGVaq241wvhVuQSf+uLdqbxUDFcYLzsOG3FxFxXEIjV2anBsBtfjehs3ErVB
mAW3E1cRuo9yZeMFyKw1gerxtgOWPmLulI9nBgvPmhcqlDy8Lsg9Imfpl6/K9zmW
yIstTthSu746ZdCUSJvd04O759z/9dI2aa77F+m2RPxuxEXWR3MJvm42CU8eldo/
03px4oAbSgTG+CHF345tVXLpkom+0lyn9/OMomNL3rN1czTJqSVvrIChQ3M1Z07H
2A9TGkWRwS23SSNx9oLuoIv9vkSaTA6ZaDOCqvT59TbeOhNl+5bRr8zTi83hEAgM
Ka0HsvE5Wn5HfDbnW5XD6arWCEkuVHyo5uJHhCHwhWcs8MfOAvU2B8UkKU/21btT
/L0GXkAdtp56p7k4BAiS6Tj7y0BhizCsWatTXAKCZ32HzTXCHcYrxMUwSOTg1tk2
p7LhjZDn2ykxoYcLAVgecfRvNzlCAQTYg0hjmHO6VdAwL7vPUbGfd7tEh3WKiXrB
esOMyhSYzNuZjLtWwqYZtbTcKrFeqz7m26QXLqhy1FL+Njhisxr75z0WyK1aWZF1
72mCZ8XJBRuAqHqzV3oyDrgsL84RdBqitogYZTIZqkjY8CaXthPzu7gyMPdAnHV2
VtTVcM/p7XGeJRE9Oygam3sNr1kPlDH7JfOaKYjkMVQDycpK5jVp4wd26uIoTzdm
Lo9LqgeQtWdlLSyAX+OPZNHT1kGHuikHRsWVQMYS21I39bkDhw6CcWlyz8uCGcbM
Is1vjT/+KOXUiF4KJoC6h/l6kz+l45O/8SfzTAE8orNqpa0fX8Bly9Do7P5nghKn
bu1Hzo/8M0k8ntCSyQUXT3Vaw5JqWfXf7+QyT+LaZDkHYtURFFCi9aIyy1zrqxof
LL6ZceABon8GgisBYEh1DvYHe4iBm8DuPkmbJyFDw4OrwpNU/5IdryhviK0+SDf8
JUJmAEsfeoSttZzbqaWXNXq2ZkDxcmFieGi9PUVAeqewMvP/uKe9JONV2lGCVK0F
HH4s2lxC11BY9FTf2mE/LyyBUQcR/lKqSjCuYNMwcSLZgE2Bq1UBbWMRA6bPWzyv
ZD/yB6PPZj4bKDYtf8zPpRG5womVWqsmtI6tC6X4E6SR9MIKzHCzP5wQKityXDyC
t+zv+NBynPUIB9B1IkhKJGqyd5dwbGiud9WPljeFoKhJ8F+DKUSjqs+wTlnvydF8
GkYtSkO77SiHUQjFa0Wfb4cBzCkquA4PwhnN7EZToqrOs/4RSFA4ZeEnkqOULkD4
xEsiipHG7WfaXcEnEdq41oZmipniUTTwVJyaiUQAM1YjPn1RiK5H2ugbvMiT4WpJ
eYLAUDiFmBjgLZpRW+NbZ1B8OGYjPYwfYk5Xzmigfe8G6ijEcavAbAgZjTuNxVeP
aTVINzPGyNlKDfL/0whaB+E8gx9VPsyFfdzgpTL8jr2cuoTGQqYe8QMRedNKYDyX
dDJZQGxXx/XJkeDWyoZsVN2utFgIwS5NZ4Nr2aSDJljg+u/7izndUt1DWWb4X4cb
7G62SvhmmvH0RwncK9MMWNwfGa336SiqdN7hEP7g48Fcp9mdGm5NqNc9/L6KYW1e
Dk3QFGeycPo50Q6rR5Ij/thwctq+/OUk00Yz6CXIEAiSKIxNEQHLa3FnNyuCbbBm
JNP4emyKRZKBsSlprkNMhy66R5FEnQjYIEVRvWfj0b/O0GjpmotnwWYOxBP7fVfY
p9Xel08BWCFZZxlJyyA23vj0VfeW7xBcTzdoMQo4xAX47eh8KGBkmuZnsXBOyWPV
YVzAouRlpmiQrmNmQdryo4CLop6igr1v96ZJN6aIARWqwI/5jh59EuK1c0CBJBt5
q/08RDlH1/p0gxpf/CYoPO3xF334BTw8RRYwjc1cQBCKq3ts4Xkzjw48rMx6JGLY
opQ1pEeHflxu02YpqeN4iX4xCYhzXojxWr5jCzKJTvW48UU5ueaNkEVHuLmGjb+z
G7V2cFabuW+St5gCqxmq0Yqu7bPCeIg6VG6hGBvUb8eEOmKHE8dXSvvlVzOPNhxw
XHFv/N7bAJ7mk6QVjmUJbwYSzczcYKdF3sYWKHVAB/R4T9d+q8oKNhpAsDeRmfTA
6QdeOFEz2ZfoOqpcuHa/2xWfdk5SUQp/WtrwblKRM20qaiccGKcCkHxW3jSWnEdM
uir7ApQRQ7SAN44ur5EeH5j3kSGMuvgdSRU5SHYsLe7Yz6jWXN9Mxtnsp1m2TjYA
BnPIkx8PJVKmCErmFTBX2eHYLT7+QtOFVCF1sWSAnPw7gkO6VbEABubeAxzhxNoL
oCnecIP7VVmFfzJcSqeSrvmCQur0XPBalD1dVBp3zGfgvrilnQ45MVyXWcCl7Biv
u84B5FHz0OpQAt9oBhPX6uIFQKvUNeqNUYCqJ6LSopZzx++jH69DNACz3VaeqBg1
kEmxWQGUCPJu0WQGrj784lRzd8Zt9+Ajh39Fdlz0gWs8r6+mZawP6ZlzGOH9B2eC
CXTqskSB9XRya0iXHVsOHgRVLoDCoHNot8edHObfbmvyjLdKCbeaY/lnv9+hk+3W
NJCfZ9tCm8PjABty2E4QmiUe9JS5O8MaQ+U8dMf+hA77ClpTmdnyxcxbbCHxMMrp
RmujT6M0e1jXofBXlgFgyqwt1M0RnID0U8Z+H7ZZ9y8NzguOAdl/Os7YxDT1ItB9
JNe21p051ycmq6W5w73pbF3HcbVH5QWhdPLfYjWwIq+yHeKpBAXcJW9kZYj6pnu7
MyMN6cgZD+9K7E/y9fZv8DrcojrYcAPKAYkP1TiXR9QhyoBBgl3v68Bz5kNiBnWq
v6FIrP+034QLADLEZDvsZZc01Im7TBCDPidHkv0/lRW8VrQq4Bi0PA5YnoU+gsU5
Wd17G+GD5Pi2aeYDr+iKa9Uhe+RwxX6ancnNBR7jqlu/WC3z9LapM0Mx2lG89BsV
VNKBgdp539tVxfhF4s7Xv5FVi60DXMA+GL1udsAQUMBcPzIpwSfb+ldJOG0bOG/L
3nsYsc3pLlo7BeB/5aLxYfo2LB6N9+r0kt5TtMIny77p5o9AruxGoTuEzdajCN2J
1+9lZwdNF0oOflZjeDBfgsJy3PixgY2/i8b9EBtyEZoXciNBVDAAIVV3OYKae1Qj
ktxoVAIwiYTqek2OXdrq/VLhoKjsUZuoH+061F/9NKAYncAJpGjw91WprPE3C/yE
yGofYvnhE8ob+Cz/0nMuXPP1gSXSZldEFs6KXRtrUOTKTwW6GOaBEk0m/eqa1SS9
FGf4IMqlg6L4NPXaF0x9Qmo/3V+EwcdEuNWr6F9JR2uZ3GpP9ERtsCzADWB8GW+n
7w22a/wudHujKBAi12K3X+5seGc4WQ93QXPxvtAOZc30c4OhTeZic7thux9vKv04
yK5zwfxxMnQdYHRp2OhHDGXWHSRGvg6QhfdprPltKk1ftVG6tnQCnRfMLDJj3Eag
vPYROEwUnV4s5DXjbsCmxI1BIpgj+KMQo5gV+Or+GShUDJlCbfm2neosEQMlgYjj
MBWOeI5mOxECQPCyek2kW4NOtcQfGDIi0UkLeBWTQD9sWkfj6rORnId5hMuLHkjw
dY9lH9vK65lWcI7QslOTkJertLtqDX7Pu3SA0/eitFoViU8yLgpXdK82GwdMi9zl
kSf+0yJnrC6jMYRRLe0cwZiY+kNqVdprVeUXa/9upXx4eaWGiwL9kVFoSrXe2dbz
YNowh8EPofmnBYDEAkP7PddWXP8uqYoVbY7SJqlHp187PsFC597+YTEWkcDkg8Cs
2SRLpdLbwRDsfLB7ZKgP24IjxxuqQUnVRUXTfjK1I4bwjudgrIYSQgPg6/OYSJgv
P8ELw0nnNQzFpK0yw/3vPin64KkrJAWOB1Ta2HSL+gl85tWPSBCfTuFwD8dN7Z9d
Tfr2Y6qXO/6ce+0bx94Pfhhl1TSfwEMZdal6YY+fHi30kPrtznBZYrhBEyhjYd49
YQ9u5UHrSPL1TlNmHVs6BYEdB5o7kh9CKazmSiTOsKFWZYhOcl8y23mAph3ezSWV
LUNkcUK39bTJkSu2YD6HOH+o6bRQGXbzKeh/VFPySuUyImnQUJsVs0UeNPQo0BaM
uN203fgLWDLSUcvxA5Gx7lsLR21SNWsxUvbPRDtqQaazuw/8vE8Hkc3wuYsHwOyu
2/FfPI3vMfZsrxX36uH5wzDqJnhDk3EzKbNPbvuhQqZ5nDX069HUFrMWQriIBGsO
f6Plf4sLBY3ZGwPgP1KOf6RiPB4/M/JcBUcCBei3DinnX34vx0UFDBUqN9h8ygoz
VCGjAehEjVWtOd2ms7FBlwKU7WCwtFEyWUUzsfFczDTVQlKLgSe3hk4A/2U570Fu
Fkr/FUiN583FJbfvPXfiRwu0F0jYVwsbCUW5b7yvr+1Fv8cAwLikL5nV2fkQPJIx
qQAio/kmTrSelh4M6RH8mA5d6j//53dggi3p+H5tLkY68VXYXHX9mAHCGrGcNplH
PoPdWfDwFb/CxKxDKVPa5DIlPyas1748h+QHbKmQ2lCt+aPrFGfme+6AIoFwixWS
w6965zr0lDrtPiblap3sUP6VgJQTdgOXuN5ne/NI8qQxdltYxSaXh0Q2BphXSSuM
OdHKfS7Y3yUjEdxbjMHrd6/+eNk1HTHARtxl/UGr6tBzJA1Y6WTzFOL0d9DxtoUE
QF4O5hx5PpQYpWbziY4y+qw0xRnhFD1MiMASKDzY/c/jWuWSgvcckwG6lE20HHaE
7ufNcxJzTJrEfrGyPGYzhb9HZsFEStL4F/cj62NLpTMIpf40+gFhtwR7aeRDf/qO
Qs/JpvKwwnDat0vZ5FTWDkuBoOhaOCF7pFCCN1pXOqfg9/+dqzY9ZV1pOGeQeifn
iV+d3HHvrw9rQflZxU/DbOgm0zzgirDTwZd3/dhyxFhDmYvFsI1LdFPi5sSS9qqi
BoFcpsUxSEAE5gDkzjTMRVrY34qlo3aPUuQ08U8knwBjrYGq5p0LOnxDlyd3Gn9E
Y1FyK7pjNCRGtyDezOjm9iJTZNR0ZcpuHdDQPwErUPswmuuraoh7/vfUrM8wl1Hy
TmQQscfQqvJ5aKZrAxC7dxgb1NDLZNKBfaUWdP8GIL+fOS400rOE/cWmFmflvVS7
CVlYeGXTD8u0PJTXW/iNZDsrZoE+OH3OXIKIjfOpAEjSSQr1ChEr2LpgpqK9a93A
RMN9L1tlL5+5Ae8bTPpDbjCzS8kYAj8Cz0IrUUrcY7d4g7TGER5GTf/XVp5OqKl0
GHHS3B8VYpIiZgBjrXiXE38xWcUHCEPhGxP/ILXVi56qzwiAb6Yphsl/gtpsaltL
HJDDxSlL1zSa5iAzMt7SdsNVrJllYpwv5z/trhbW5S3Biw25Y3Uy8HQisrSjGXdI
OIj/kw7S9BSmCA0DJJ0NHH68DvNK3yXfPbyHVVWnbtisi0GG8WytzG0zjbdnh0wC
sNyszVcKj/H0aPK05XoIlyh+0q3YuAve64nE0UJxxTMydrC2JTjw3uiJE/JNl94A
VPopzXH59zJmOuy0SHxMMCbptrGXWq7CumQeCFO3ZSFMqhjuBh3m6Qo/eGaq7BNw
TOTng0vLo1j9x2LdwJpwc2dQTCFtfhC6Osd7MEgmh2GY8ba3xFlnwHRigc7Ee1ga
+RtdvfjiJEGt1ZMdfclNfAyhvOydQhmfgN0ozumCKG5f3totnJYSbTkzxOaWJ3Ck
fNw5Dnm3Jkd8S2exuNiaA4hu3K3Ywjok7y5VDJaqy+48oYxgZUs9F+U03JTgrAVN
oFtWhvYTyi41kiyvRPNtcIGuR4ubyTjQnSnUosoTIDlyZGSv1xxvo2JUIrE/e3tr
eIxnibMq2401bEfiPN91lS7dPT645GIGn8kBQH2ORgEi/gdBLzjH3xTjfi+2V0h+
q+t3obz4qI8y2wvQaDLY8UOrJjUOSF7pzq7jTjiLwhh82z4Vpk20VKXrwsddXMpX
Fe17PKbfTxxxWaPdWZY9TEJXCnbNL5HsUk2pLiq8UWf6iJQ1g99DoclCEz8p5vEg
jliyPHiV4UPr3wg+uEs0Q2U4Xc2LJVfI2f2k1O1NNcuY9xUMkN6zux+EczEB/9xa
khb3WHqr2wUUvcBCCr4TEE0RMpDs9Bl//CSJLeQYiAHTjoJZGhIwBWL2mkCNZ1Zp
qpn8THVrA/Cpb4MT3Ws0odm3uvhox1hU3KwsqQf8FfqE214NEKu40PKAsv4GX249
2wtCCaITqtAx1+B1uHz2VA5wnZm/CSheNkVAAgTxFhKLCMMRmILVTu7TTlDE6mW8
35ulodFi6CQRN0h+OS/hvLKISz/8jVYCM7CiIICWffAI4nWdW4QP5QRRnLPUgnnQ
JbIOk8w+omanyp5qxA98vT0xd4a9bDdnvZJJYJvNwUNkcAhHE8079u5p8W6bDINh
CwKYTt6v7t4FsvIldF/5qDcxQLq9uFVubfkmRyuMLfjPYgW+PddAuIPIX2sAa3y3
M0cR0bLH0RW0QfGNUj5weFOb5OxoMsnUhbzI0+ajaSWcDZnOIjxkYXm3wL2JFthB
NlIdhFVoZnBVjdeP3whe694xL38Pe9lQPXyTYtYRIei/wmp/FtgWKJRlVQtpVS+T
G7MIYtvz4yP9AGGRr4m5pLXBP0BafWZzkak7DkXvckcqP//7/P14U1QCV8Qu4U6R
AwmOgWajaONbKwCKAndvU8As/+esirQW/YMIogspWSKZjdStpE0SodfyoblqyH4C
9X0Ka6kTw0tWAO8u+gzaDBGNhswfJGBVSltJt2Xl/pS2AN+0Tr5EkU7Q4N+dh2wD
Jk1IYFbsDKwuG4qPr03Fx4a3z++uuaSTDzNRQDqNDli5ieNz2jJU/2U95vaGr8ap
Ld36PEhy64DqqG86bL6iahv3JxZRIIR2HysG5FSFXoaY1DKnDGiNXcN54bLpQurG
sZYctq1eBLqJb/s9nzRnqQD5N+H4Tdf5kAnSlD6oah2YJiUKNNsG7Fd+SiqkbUuf
kquVZt6T3trh9NCg2GPMjgiUag4w/P4bAjvIZwZantLuy+C8FI42Eiy179A+BPae
HR/UThjLFOSxUBtTr8qFbtaVRUhXTL7eJ/Kgw8zD17qmalIFUVZubKOl8I571Fg9
iiENxoA1MZ+BTsXx3GdiDWNfqAZatZYHrgbZsmz8mrIh2hD0UrxmrraY8AQOydBZ
Mu7fdNqB1e/3IyHp0CoksCVJFnzjULqJuCTHx7/g7zyjLYJ40hdTzy+IygpvyUmL
Sn4q6u3gHcSdEKjnBnDAFXvjr0zzP63Kbl6vt9iZJnG7t0n8SwGAoD832pZd4bdx
0uyykuiuVuAnbTRy2qF7jjmdLiK8YSeKdzzC0O7ImIhjMimvMv1jfj/U4yY3XE3l
VR/6wG7OSiXGvkyB7OgOtsWN6i4GRLXb6iRHLjId7W5myMLv/O5578hmm2w6+xoS
SCgtjqZ8k+m8Uz+JhzWpMPDpS05HFHoso0RsjelQcaZo802TOS+uvD/IRilQcqzT
fdqTau2UEybOwSUKzwqMBfjAz0yyTn0CkEhkOEcsHHZxINMen78lo5CoHeZT016p
cY/ggVyd4jvS0Ih/uPVmKxLjE8Q8rMGRmj/DUxpQW1sjs3M7HpGRY9WtDfkmM988
uvwesdCubaQ5bbv/f9MV86IDffzjg6n9LL5UHCoCsE2SUiOZPPIgqOf+a+qr9B1M
LZTgili27gL7mXBogcbUmoFyXkxUTWtpHEfigVcSAUXUMBIpSRn5noshozzCEUkG
cp3xr3XLSHYhc2fZdn1G+5A5VRtUNmxu6nLKb1I1fbPdL9TQXAhJpobcgwxqgTF7
gIXLc04hkF0nRmtaUd19N7GwsVdxHomJJY7cFE1zgfSy3WtXhjk1rHRIPxqboCh3
ydak0Kd0TVYlE4yx/PT15yJqsoQn7NzgU6LF0CAlOInqEPeZu12riBDeQilRgehY
NaAMTtjLSOPAoqy3Eb+yCZ5VPTESnN2IwcmP/lnkQu/fwX3lDt3jfjoxxB3HaIp6
BUSxmrM37+NPCFSPPyBNkLDWrvhpKS2dwYSjH3lezxuSa4f3Lkgc8sQoS2mb6Pji
hhDkrPHTBJs5p+XJSrHkXb3S4UoKpj4V1zbq52td33NB2Q26GVYrExD24aUJ6JiB
0acyTtr1F+HqsYoATgCnUGa133WbIVxoCfQQpJbFbcI12xgVBFEMJHkZKrrfx6tG
cPlKUnZjzO6h8MHF6ZPfl1bGcGv69MUJ89WE3V4TkrzVg6sLjrv4AeeucZ4HL5aV
pMPvteeZcU1a0kWSpO/v9TaICejMz/bxz8qiVKMHoNqV4oEnXGOiIG0i/Ei7DnWb
Kz18Alpa59Ptx+uXAJOqK1UtT5j3/qJi0xYIXj8JD78OyMTwPSCtH9rXWSDqkq5s
QItKC97bY7fYuV3YdeI3/705O4FXbfoHam5ycUKd4AHmfnPKGFmdMxcVRT5QRNPF
mD4ZHIfexqORuzUpE8RzwTS3fQ5Yt5xgA9DIENKjXLKXSKue6vDyFA53zIlXC5el
CkkGOy8NyRRwUiP3XfUrECom6zVGBAuBoG8Ahca0Azi6thIh6C0GDK/ey+Y9lgIC
1zClVA9fb0r+vgAncPiooWU4vW6G/fL5IzdoEqAI+7LOssnetmzkKA507iUK186L
4mHfvpTNXoA9+FtxzMkj0hvy/EYQxbhrY6m2l8R5NIOJuX5NNlfTpmcZkEbofMU2
Ev3vbtKACZSzwuKYMO4NgW7XEmDIf9+jmcVdWeZDC+qGKG73n0+MC7qiKT8mw1al
zXBE3IC4SWgLNIux+UgAYDu9RPNaCZyG3xrWv1BA6JwDy4197zpBX7mXmnHLkcAk
2tFM7TME1cXsS7W77O06re2kVXSS6f1Na6zvKiq5pLnK3o1mZmEFsyvahOSsF8RZ
irOqnCNthDNVg2k+KT+6VycDR0akczzTwwSFJlkIzQKiVdNveBoOfe5n9iyorjO5
ZKWFE72n9gbX8IBHB0cNGLSZlHge3cvQ+CzS8RmfLFWJiFsXJ/9yiOqRLSLlrlN+
MLD+x6s7BwLrzm9AlRbgXEYMZdbZbvPp+zRY7nHKAp1+nN9w7e5L0/4TCCkeOzWs
q328XiNCsvrNyQ61G5umGmGS2GwaKXQcbxHbSxYATntZ+inSEEQs/mwdJyXxNsv3
X9WiWe3MhRTqDp+2E0qqCYdLvK4ablkG9kFiwoE3orYo+IIgdzDLtBEZbUsyozBr
rwiovm/RUdiCS97iIkVwaQM6rsp86BpiSigguZ1w2kEn1AZzdSsY4L/L+Z8zpDwA
FS08Le67/njnk7V0IW+PpJAFmOa93RcpaeKyZ7IFJ/ef3hXbMJ/ZMPP+v2C9n8BI
yK+SdOyEXrp5TqtCfgJZf7DT3Fo8GExzT5wMmqFCGvwwxc/2djtMxBUdZBjhh+2C
8RJ6GVLZ5NMq5Z1V+SIuIbp2Z4iTCE5CnodXR1Hm4wq4dCQJpwbp3f4usSCMMdvs
x03OjDQWCpFgU5YUCbaL5Try8ns0B+eMrHN4Wqq+8ODYi9KDVTk6VX04ajMScJvY
JK9zTUZMFD1u9BYmR3TuS/xpd3RNx5b+v3HfxoYf/KHaox4uJhqClLgyfANMkf1H
evMY9JyfHMjEqkYQGqu1LhbxsWGt9PrugoqXo0+i8mUGr8mpjoMiK5wKrEccpx8n
d3Ht5MJSkQ/l4Izv37koQzMoJZSWKUasWz+nFvBBsDTInugwrsJP178HcKFk9YvE
FBvjCl6JjWllCt8RoDHNUjI8KEBg9tbhDbdfRkxQ9rn4tkDDj3QHzt4sDk+tkjsB
3Tc/oB+JnVtJgcDPwVSyzVWglaUDArq4C4G26fRpLtC3Awi3+r4tld4jCw+Vg0Ww
bSvofWUMRbSylApwRgUwOQZWmdZ9T6OBM4msTmyZ3XdpI5f0apUyyttGLjd+4PgV
vt6Ksbntda/A425teXYLbfr3dXrVx5Jarv9aptu9AR9iX/0DM454zwck+r5XEifQ
nq1mIyz1dKhb5Rq5lx+CRLnWOFRWEIuTyQYIIJIwwMbv/KekuBi2gqQmz56WRgTD
EMIh6oTss7mYy2VR6UHj0iAeBEmsZkChHbzHgJT10zJ0EYXuKP74T/VVTn2SUh5c
g3E3cPmaoJ9FiBS6AaYgcFy7fz1A8kH4HvHTCe518M5Fla+y3Psj5uTpy3sYRymD
b9r0r/WTYa92q3vgAWdTXbs1uLnaUcpOGvLdHczW/dpxP9IC08OtRaRB4epfvsV6
+cVu1FhHqFqpkcRia2w0+0iRv70DrkIpGxChumvht3dt7rjg8jnRpzh2vSPhF/uB
I7OT3pH2RqzgJ/P7qReielL+qTENlZljoz9aw3/yBz3TvwPu3tAXeL2a/GdTsxIp
pXuJc+Xr2/yTCASV3C+08zqFMCIZPYpAW6hkPN4Z79cUva2jMfBFtSnbJtZHQ/jD
9a3ykpUOMUQQIXJs+SpcGgYuOGFuk/JQH56nfRhO9aEWtsgUF2aC0yJeA480pZrs
LI4hEL5H9uay1bb13PkEEqKS1kWeTGP0sb/ZiST2AHPUrjpeqn45zG9JobRbtKdI
6HvH5GcAJHLJ5w6LesK5GYEyUQc3RNunWH8GejMoApujsqrzR/NuRPvRBrPCPabN
lkB23mLzbcHMAnfFzn9vcnTuG0UPFlIkH7/iYQaYCh1wKlxH/o/mvDJsA08VE7vw
T7uPsxwdKPHPY0x03781wKI09XINN6mjkCSlU+YTjZp1t7KJmXlLrOQIoWVOYjPo
z5rbAb3WeqZ4wcQ7O3XVT/fPM6OI+AscJwY4nsREZ3lJMkhq062To3kfEwh3VVrb
cJlx0drzObxx/2iYIpV46HlKV6SLJVIDcY7HB6UokysWF6zpvOozLbflTygNE0It
GmWN8qcMaVfjotoh2inz2WBHjQJ4BTCXKCOwv3FxL7rlnGaVrDDQ6T9zguZG476y
ANbKHNA/yBKZQBkFDcXhEyKz2RLvlxQWzZt/4v1IgbBXJgRlHlUB42dhdBq7FNxA
9b6jhO1vIdJy2KRhCXQ0X2TG2avuJWECr/7Ke9EWiZPfBLex3SB0PBjDBa+K+ZBa
yr4xCoP30PmX8jvx9Tj49chcavYVzsspmzFfNsU9xGH4XKI+xAUW3NIKv1tVpYr0
e8ccjW6cru3ZoFrTq/tEzY5h93RZeV3AebvhCWCdZk77s/+jWypzeO+HmXJmAWOG
GZ6REfEbIR40OjOo9IBJKmx4Jg8NPH0ebC9i8ARyS5oQXD34EPg/qyYLTazf/Jzx
QoJ/Z50GlFUnMmcGGSo7a7FN6WXrfV0HJ4Aa2gVMiHPxBCfzK0r5vpIBMYMt+REv
lAIjpFbgziqt8a8uhO/4gFkWsKjyrOlPSzlPrVbc01H6z7JCdLflCShN+cuRy8mi
2Jjlc+XsA13m9dfVSSSW/UrH0vbVZ7L+sUrbFe/bouHps2N147Dz9GNnYl4LAcS8
V8zC9hsLDsaDAQmJGOKkgEnLQqUIZxRM6jEAUneQH4k6iQhKHwDCn4kKmXo6jL00
55vZCF4KxpSDzBw1ghye00pZGZDILiVwpPApW4H/KOvv6iFTJJYURPKysof7KJ1A
7IOijy+NYQcvMHJxUctLGccCKdbEyrbMTNZ/5k7eD2u2UkP6RH7VPoE+MSuIW6ZC
Zcqi0+Oyb7OC/lffFyXWNI2N3XOxz0vU/S/PXTPWRZqv9Rf3Io9pv3uyIxylyimZ
oIkU6Z4xvX08ckKTHXqsVvuu0knKPBrMJaPW88Y2KdykJ26shihiZF5gQHJ7vKPt
7ot3xvhT22E74bqOi+Z5BzxVmri5ZFI6agCwRvoBTsfrOVd6zvHdj/KhnhwNDHBp
pb83iGW0YYlHEAt/dD8LL2ygMsFLjsCyc+QtlyLZnYczprddwJFlwYdTO8vTIcXA
PrbwFW40R3IF5dBN7CjkgDtz1kKz106FXF2Lw+x/JpG+OEDaI2YFbW7y6IZC9tKM
klRKzh8qTRc3Z3df5wqENQ5rGt5Kte6qWrAZ65rOh8e4a4L8HWoiITOsWpPlyVcS
nyPyWuoe5yOGcIuF44RMHw7fQVIXQoKbET5AXjiWDapdyVRJ2jOrkp9ZSiozeSIH
4Djc8qeOFwg84U3EapEjW2E72LmT+DrxlX/fHcmO4KFJrUnDIBMUmMbaDsJ8BvIt
VWoG2C4aNxQz9YM8XOmCwatMA68+y7FlbHtKySC97Ssi9M0qX2MtPIQhW+ZBojh+
aFz3kyS/0FqI3OyWTLmbnTTwXL9PwP4zVCnoBctfgiA7fCKqSqlyI7iqTZ56jnln
NW0HWvoxc0EVcjpQbx7LWa4vdpzcE/nSJ85t4e6zqcjT5ZnqOh2I60X1KIEASBAQ
9S2STkb3d6Zhqgwu9Y3hkGZvnLaR2EZqDpHLOysQbeouvseYzZ+jZ7IyEFKZCT8I
wgW3mitv3KSp/3nkBRPQt3OvLiNoaBGAaK85KSR6/Ns0FrvD5KEMWnOwJMxUqHxr
JliImUDMN/oMCBtiAH5amjf+RZR9mUiHN20qIvNVx7vH+Nqg4bFMhaJCrZHKcFEw
ChYzD5p6p4NlshBohbDEsCZkWPu9xXvoUeH1AqLUSEN0W5c8fzy7DBqt45bpSzLP
ETTDjSgeV8O2cwQnXkDB0BRDcoQwInOmRDN76zzMVklnfJznaLMSnFLqsDY0f7OG
kYFGVz183t+XZHpmtPDAa0TXSzrQTMuYg+af6iyotqJveSdDWgcY1iXeqyU4iPlE
pPpJZ7fHrGEooeeWaokhCyGxv+Sw+yzj0Lhdo22cSTYNQgdO2V58YaY12B1NS1xw
kj6WA9F5pkU47+dq4vGOVXKh2myEe2nLKGktem8la9C9/WBTbnJaoOeD/JokruJo
DuJS4PqAZpSZSMEqpq91Ia+PKcym/+wYq1CFjaXAeeu0Osts/K3w0x59qp5M5/5Y
H674Ful1ATzfyk0VRo7fSJySyrtOHY8wDMxGm1aKctSELDu0TkTdoJupnBmwu0kB
k4L6KEFnXZRZ9flZTgsRH012LPo2h6GApV6niAsfYvD+GWtKe+MJ0TRFyQ3xSijo
6zU8RIpD4tSIus7d9veuSgw+hHxScQ8HiOmO16dTc/29PT09AczQi2olzph9/NcN
dYRr3bO432iddEKwBQvRr2/a7K0e4pjO2Hsqn8sNvrN95QOMwI6pkxhoPy9N66II
0OTiqYjzRhTlUquCSYe4NkpFqerUpvxVzhXo4nn1v+Bv9E8MjKo7JDMQSrQe6IUK
mrX1+1WU8mM7Ou/87FKLlGAtW8GxwJIWEbHw0j4xecGOIcl1r2NoFW9IcAMeHrh2
rb4rjsRN3zDKmBp3nXykz80Xy/2Bz5O2HbHQHkk215yWt4vJoWmFPE2OAhdMQAPz
kcUfzOzCPY8FB5GREDgbIxAmDzoZFcOUI/zvEkl6G2QujcPNz63BA0icYOOFCUMQ
0ivEOE292MdMzGj2l/yB8pNZNw1viJfwElCXns0dDGkZlvQu3vRFbRLsipSeA6dV
Iz5RlDpLojh38BRDTBNc6EiCPn8UdmmGthZM+pvruUUFUNvW1xn8wjqESXlv2xHj
YxQE0PbntEv8jW/IQ0Mvx69jbtGnDXCpiMbr5MRvblpTb0basuMR7SpiofhQ8OuL
bXFcQRo28mPVNFJXfJ+HTvPcSn/R+aNuEdA6kHc1LWPXS9xmJNbLglbu/Fo7H34w
G7um2qz/pGJ24zhNJJGhsdoZkvzgqyQpBK09bSKWciXEwnf/IxMExvA0IL/TKrOg
kFSMFLJtAvE7Fd3o+OpY9FDD7DAh9/CPPbmPTd1sGVkWbwQVHm+ZjS/UrDItftNB
LHYdSONDYbfIOABAGfBdlsOVdIKla/TpY842e2ACizY4rE+8ipCyNRBmNYwTTZ31
3zauNrDuqsaFqqOFIc9Uqb/DdgCp+rCXKanr8gdjO9F+xoy/N/kxpN+CCZZ6hbNI
vmq7vcBQ9bJEblKmRjtqwDc7UtwKdTdgxhyG711dAcT3GC6L/hqQbXb3XAS+x5q8
Fb/uy4CfpTdoA6XVPkck6XejMa5ICltAp1lJuCuK5KUTZkfVdUDvmlOn/iKUjhPr
YkI/BtsKwWaQC1/aKJGqracMFniMS+ald5STawPhEgjLq4Sp31LGcwn+MoQG3iRR
vJXF26aKCcc/wRchlAof8560zBRXKCbMpMA+I8oe+3KOqfkYwLWN7KsOniedSnN6
4AZE498Eaq7/bWqoxIWd2mmjG35PWMiZ4eEcZIJ20+B3yPHmB7XxehUUpPk/ErZD
6xvi9vqMasQvIOQiEwVfEjO2xt8jmt+J2ada88GIQBd1Rl1UeRzn5FzhRHZ/8NBJ
eakxbnIgV7ktfcapD/0WnHdvkGO1Nr4cK4VNdDdyoUwiMkUXZKw1q3RTnyKDPSpp
n8eDT4HQJ1/mLUFlF0TeEhzTQEY5aOV1u01+++lyhWViRsAVIpNCmBKquiDDs0jH
dFm54Ng++ZFQ/QKh2yxUj8f1CvQ7QCMu6xgHMlka12X67xbZ5R0dbwTu1KMhDV23
iA+dDNKJn78wsMQ96jARlIE+ByXv6b02THiP+6viijZPS0k8JGAEqqHMgNm5Nzxm
NrPL0ykSYf2gDbfEBG1cRBwaWHNR44cZ7/gVLWY9ZYjKiwJ3pwwKIP3waDhaMEEj
RdTJIFuZx3GJIeoIC7OGPfH7qq7GTpjzKIc8SlK0Sc3kgnmZIZ9XJz8aB37MT8pM
CED8rqE1vAX1GVeZF8eoiSmiWQEGv17R8HXhs4zmQC/CJhW4PPexjr/+lL0NbnOx
0oS9Y7u3Vuw/0EuU8DWEErZm9qBfOW5/nsxfzXNba0NZdXJUEQNYGpbO23R/lI3K
tY14BoqdDiWvwfgiURaXyF9fpFFerf+Pf1pe41/GCY46bxwnffqW9vuq6eFvK/oH
3gB1PnMmp13r5YNgaD3hUJ5NDb/We3ZjJCpJWjlLm+4CRShlAo7N+1Wd9xJ2zERX
uPA1wAuLD6AgRXR+Tc3rufDKFm+JhbwiM31MyaTD+YPAKLI8+CVna3/2IZ4GfhVX
y27cckI8hvuXkjvW8J52j4OuMM4rJ4XFx5f2taifkY5DiQh/D+63dUpuEqnwOCav
XYbwqZkNlz6k6W/hZUlyrrSV93ZbAVs2xN2EfOjXObA4oOocoRLVQ+UknrWdKRoY
DsOxazdNzZmGBegLzFs5PdT7PVGTI5rryOg/Ut18/DxOkU+RBxQstNTzaNdnGUS8
zk4X0v53bBKScrEsizdFckqc/VmuJj6leOL+nM3PA5Ey/jQhrbM6V9vs9ZjSvjxR
UFPUjfEV8TN5Nsm4Yte6pQzsPs9J0PreUHSQy/w76L5NMlkIfEI1vUKsYGtyTaJR
budpQJ1HeO1uzNMzwRrDgibG0qxQz8ZgCdfhBd2TsX8xkbM+k2+VKY0lPUvDvDT+
OU1gDHgt1VARfPxWNdxLMN+Wc5H5to/ZDB1wXey1t/rGqKKwfK95Xge7pLeRFpmo
LClgQvDkAk3Ml3z6ALGrEUv2rdBYuBijwIvTQpm65qWyRGJlpvfrNHucc7Zwa6Qs
YoaaMGEsLhMOBS8iCYICbmJtMNS7vIvsWuo7obXOUiVkN/QMv5Ogoe9QS5FIe4Cr
XJjsmUv8IbsVyRa2jHfBqa/NM3WMDdEhJZAlba9T7gsFipGx25JPZjOyLGvRfs+J
einJkf1JrWkjW6H/HE0ULzhajbwOePYUmO2kgYaytZ1APw4Yg6Zd05fV8KwIuOol
o0q8HEXiSNOFRDhoIuUWYWi+I0So50mkKN8dyj9knTsn345NKZbE/AOeh0ZYY3xc
V2p879lwms9a4q3MmCw62UMZhuU4O7om5giLelsoiOakDyl/BAuK8H94SKorHPey
Cyqt2gmBT1ubEpGmoxtoF0s1vbTdMtjCpUpUtG3unV3Oen9sjM8s0TNfMJ5WZB7T
VTAkOchk/89HxdwrEhbo84jIo5NXaO0lK0oHc06zzyJ8xl2NApaN2OhyFHJjcJpw
ikhH8zCYALc5DVmd14QwCNc0Vd8pucJQxmrwoBimmbOpiFP0w/tAV4xKjRXKWXyg
FT23bnT6zsQUT/EC7H/g/UF0Z6gBccIuTJo/3Un5QXkVW3z+KanBH+QNTUC1Jtqa
fkwlOaeAIewsmnRGYOlwFOaVC03mt/8Kkzn3jkFtTqbFtUhaq+xZ5Wc3q4InFuG8
s/kQTfX1SltUbMdc7KXoFVZlzdCeyoPcW3yTMiBqmlWVCPQc+R/bOybNGSeYn1DK
uxw3C7nTnFMZIHPiGs6Y6PkN3YyYO8r3BstVcYC7kuxq4iSbYhdwRMZpKfotCU4f
Lk23IXxpN7uIh8VutREB+66BIgAKt4b54KWhR3Rdw4lDpw6l/2xoPoS0O+JO6Wpx
N3fNP+beV2HbPHLSavGahJGEiFDbDQPDgk8Np+6+uLd/g9pFBXQ05xTYG/bZJXg1
xvlY0P0J7vlANQBOLA5J7cwDWVWCossAuQ3neUoccaMMzL+Cafz4oYbGa0KEAZvv
auUvqabnP5t4HmYpHOAp+0OQ0M+mmWPEcoSRB432aruRjRwx59NspA23GawU4pch
TgNrKSPCV55UblqGYp+T5x3xUO90VydUL6srHWyr0XSjFR5xYs5DgL1xfH49KUXf
q/mknCvImaLTmP5NWd6rpXKMwbGRC00gjt7oc0q5as7E3MmJOsm33gTMFSRY3AdL
mDgqAmkQjT1coDLtmrgxaKl120l2mhgYXv0cxTa4T9uwgbKMCk6xc7lRhFuqTiGL
aqzD005Wid8+zszKhD/+/i0fNUBmsKx8bu8DKm2s01ldjgAbYVRZLLz0bDyPFshR
I1rOcxvqT8+WOT9iRIEK/K/O16oOy5YiZkw4hK+Tnh7u2imWadtNptodbdwW4bNg
DBmFRcLpBpMM4YgMDI7fNGh17OX4ctdNeVPhoeer+jqbgZseVGEfYqNYdAtkeDUd
7wDuSIdZ3loUAySdfhnP/dAx3O7EAOIOp7sBYvd7LpbXqVpwHwwDa10UvNj7kC2i
qhm/i2KcX16BAka9SZ2rP0f5LxYi7yiUOFhkQ69tkcgdy9kMWvQfCNngYa09lo9d
18wTnTPI9G7cjqAk9O5vj4OK3016+83gCdj34vBKTrq7xWpgmsL1WdZ0erp+EN5k
SsxAB6VBqGOAu+1pV/1wPMJ60fUs0XsfTrjL41OU4+7/MW0R/BQhVvPJL7HFtSlY
Ib29yQyzU4VUAhK1SYXCKD9hBn2YfUBPsg7i3SZYHoJBH1PPGBK1mhx3StVt/ltO
KEPvjZKYaKTfJkRDM/fY1vgSjsjg6slsXLe5p/bqSY3EUPCCoim+HQewNIrhU/Nr
TTU1K3i0MHxYB7zjSgeBdz4nJBvJZ/IsPvhY7hc5tUGS2a0QUTybG3VPS0vwcQY0
stJ/oxl11eTvVB97j0igA3py0sjYmBPPSW83CzFTHDagHidnCMdREmp8E3/NGQW/
lCXvz7sjL0NALMWgUOI10grrSLyQhlANLay3UfoMcaJEy/g6Cp4r1yNG3JGy1LqB
zZali6UUm3G5Z+Pg6Ne8nefH9JQjK2jTRzDTo8NbrIMF73tNqi1zbANAA8I2/Bue
6ffe4m96PUeixyjcphu8bredd7c9EErRMjmiGdZvOxFkNZHyMYG7E27T4CABI42i
ncBCb8/M3q8GR3CUmfEbDnpBejstHvEFogdkMtdNpc/PJMUckocGbhn9QSRohrbD
QCi9nVGScBaeDU1rL6Bo36HI78FBNcOxUAcX+kYSsXTXvtQ5JsbHsbb+Ks/apnN6
gEX2b3zPNtYi6rx62PVki2YuFHCALIlAitgadBdey4V73Dg7sgMc2WxuwMmw7Nas
AAl1Fw2zTGk/Z50WCwQzSsyMMfhLZGi5UKM/9vjIQyBT1oLpvyy0YJC4y+jKqZV5
7zNlDoyxKhsZC8VSo2AI6snJJM/Yo4WSnXWXqEgUHGMTSsugY6l/wltkF9EWElD9
JZ1MKsjlanCTq/qc9ulS5th+SzAYqU36Npcx4qQRGmJSsxmNswoNoqYlQznXC1R2
p9xnn3lCXiqA8uic1kZpEx+rOhpjpfYIZxwXQbADr1B2uQKwvc/YNYy6ev5YSRto
+t2olOhz7rGXu+oEk6GJJ/af0xrK80/J8ZmG+SX6kM3ZNl61xXzWtX5sbgjlQnoh
UVlqSGRPFljsdv82wwo23AY+UHOmxbixrGv+4ohisP3u0dYREUeWJnhvNqThGKDY
+REvHklJLKWI5qRb+VTZ9ZkAiIEj70fTK3c1BjEidohL1vKl6YfW6db97WAAMn2b
jwx6jp7jdZ17vIXZUAxol5QRn8ChLXV6lFTw2HFHoMEwwr84rYyfETmFX1vsGRvi
hrFnfkACATMdfxR1BX6qq9dGJpcIEEq6tF76cUoUm8BoB28buN7b9Ljjwaquk2II
KbhbejCYSx3JrodmMjHUBL2TdGsk4Stb5/epPrLCRNRtddKC0lgSOzw+owQcX75a
7NctoCJmUVQ/9isMs+hD+UDSdMaiwrV2YVuBB6jAxVqH0X0muSeg9oN2CpDUVUz7
zoiWvfpyUF+1ouZWV5Rb6G9lY/k3JD9iPSrkk1HfRGEQtvHNV6R2zZXewlh7CTcD
+VJBnqAwyiBqqJeow8npnMYij5x4ew/XwM6oUq3yL7DNffGt3V/hLlkeeZ9CfSbf
krHOnRll5Po3LrpS11GtQCSOuBC614q3t2Zfo3L9XjiKiZewHmYEYTTk3/ii3wdy
jPEsd1E/oksiIH2RvEXLvyWa3VrR7AUs/KttoT5SvfatHL6ExeLaKody2NOWd9Qv
7UojHXQhh4ASzH68O9DSXIaUoguKv75uGkIH+IxMSHEhBmbrJ6hArKWy+K74WBAW
HU7AEMOYNo+Uh5kuMuYEGo1u3f1PzewD4fqdWNjVjgKV0bvZ9P52E/NNVKaRClIp
WKrcp+LPjjVpyy6a5wIRDb1S9/60SsQEu6IUbqH12tR9+I6XaZpWzQQowDMBjeAr
ZwgTOkOsGhl5Eb/PltZhn9d6xbW+PZ1cm3HPJdjI8mTxl2iBDshazt9LFVIoQUPt
rYNHIMxNI9VNwpSYstBJfUgi1qNkXw3YiKOPElFXxSavM1LCIyavG3p/+pGr/rIg
uXfy1paIRfrXd8JT8OJ+RvIzsCJYvJIqL3E+BLa6kqPwvz6vbfoDPH3ZyR31u9bA
lEv9tZtVk8RKpyAkmDRw8CVHXTKmoM9/JUHvJJVMP4bGxfvPFgxqbpEosEl9iOot
uvvZgrCEok4ysesw+hEpxIC1RB8Be22KZ5BHH+DGINK7rxxGcPLWN5d8YevlSvhf
0Xah6nq1/M0EBEYurnw+fQjPcjY/Q4BJC+XD6c3Oi8XRlKTgNVt40NZbs/MEkT8e
EoyMqFJhmWNxTfvDkRYFVFKkdofPe8c5+jfUetFV3OnucRK6chw5EMVmVGpwcO69
2AJVzMOWQrTupG1As2/GZy4igsIdx0o+YB8qQZvrFge/vLlFH5Rf8O35DCvZj6M5
x4AUYbBGH24kHXppmSX4oea5WdsKwGuJ+4UtLuNBoALsvB7tFXqBnVyvDD5OBgaD
7noOlZdR9vOt+sDMNWze/7ZN1ztvE9y04BEwdVTQfPkLRwXoLrmcCZ5GpxkSeUoz
ZUTuUo5aK/Tm58hbT8cIDuB07toJiNa8bYssoa24nmbSLO93U4e0oatwWUFY8oh2
7pY1JcB5BDQumfk2takpoVj0+hWcCI6k4JQPiEoZ/bDxWsLOKKISreOZ/VpR54FY
LMsrFv//D8J7E8tZCUGEpNrLSNYMJzkxhTICNCqJjZdk+ON7OiE8TzpdVlX7xsKw
E8DHvV1vf0S+JIUL8b1uBuqEGVNjzUs1hRFZKL9e1IlIx2x/1ASn8GKvn13cnsxs
hKT9gaE+cKHfTCHxvPZdvC2WCob7STAANLJWsoffzqkBllfxoSQwzN/xuXAT8rHT
rpAtCCf//s13+WORN3iOOyTQ3+56srJ6MhB7Ua+PmO6TQ4sE1WFavF/lABVUuEUp
RiCvx6EOiQEssGsUYdhBNCl6iBCwUpI5JvmeemGHISiAjjFMBRcgxqvqZo0ncAWh
bgAhXGavKq63Ybu8vRRyfG8xjT/zOYW6XQha73L6h0RM0/szDKGyjBo+MXIvU+Py
rlb5xy3mbZexBMLeTj+hgmD3CWjLpeHwVGISX0SNFI+7KtoLlCEBeowFzeDidiSC
cpD7UKdT8V5eWZdXIyLlcDw1ckLJOigTjujz2BU4zzskVBomUAC/gTzOHjKDMQWb
MXkksLFbi0YOY97r9vWhxgdrA6dmZKrM30/wXVf1XKei88D1NgGQWgo5zS4KCr5/
ASwO5AnBFQjplucERyj+/zB66xKLiV1sXm5I3UeEd4wrh4MI73MJ9VGRzsqjDOhl
IoqTHyv2FNuo9Vvw8mZYNSqYSNSEDDdQJMbyRiByySKgFcqFLerSEZXvoThixZ1R
HTvvm1CQD1a2O0g7QBii66fTFgELyrj1Lw9a7gR+Cthn5WciP7T/bPLLa1b1T7Zy
XWasJsLujQNXGe7GIgER3jD8+mpulMZtFdcEC3Nou2WO0Cmq1EhglYjcHP4n11nh
LZLeEyjcB1+QNwuXkufW2eMOED10ab3bEEt+MVtsLF9hWq+4Ao3IPoPq1rx4ZnVe
Hp+ru5UlQVcYIw+ZsUB4tpj1ULR099dL3Bpqk3oIWIFzwgYXED8bXvJlDryuWJ0j
4TtAkQH9iv1DAT+Fl2pSRR+rrq8a5J7X7CexWw9ekEvAWgZAr7QFdz/QCtQ5jSjY
9/1aO6kqu++d47mbtFi5zmXLvEOGryN2StrSP9YdJTUn+ZymdYzZ/7jUNCRqXbSz
eUpU1LBo+oOPTqs4woGSzwh874W0fP7FMOEuPlTDXP4r1TTb4f3SC8EflootLs59
eewCGOLtCYrqfK1yoVSvQyeAWSJCDmtLKVkHteNd1uR0TctrAhRJwS9RXu07FX2/
gZWQLvGSXDh1uEMduA6+XnpJ4UT+peILsRsftWsa03U2uPSGc2JjHAz1yllBMI+h
ubMTwydSkzxkesOaJrKm9kUSLM1FVW4GI/IWdAPOYLCjfQ+T53QEtwmLBjs85wfK
8yQl4xAOf/WxWExH7xM0bwDV6qnsNUK5usselyZt0GxtIK+9wQ2UIdwBBzUEVoDX
jG50aqOh8pebcYifBbU12ue7ugYV1ALI8SNxhhnyeGvoHIp1lNR3YcbfZEpMtZya
dWpRLRaSrJ/SJNgkbl3qE0Gf4qqva9SxRkFMde5xbPFOofEhlhU7wvmbfwfLcxOf
SesZzVSP4/6ZUli8hfWy40l/IPqtZ7WPkSwA+LO5jC5G4pWADUlIBQYoGJu7P5Z1
uZPcXoKZRygF1lPP8AzWdPXep1BDVSysBiRJMPsTZwhDZvrs3b2of5ByVHdReiU5
3dkf0iNIgIKPORPOnyDrd0cskzGvRnhHZ149sICVXsXXV2q8u2DyxlRWwu7cYSAl
9g1cCiq6cGrHE5BtwrqJW5GX/k1zNhigdiJCRZs83IVdEqyzum72dmq5hLPiSO0B
1PL9ZWPBpetO/iT9FRfMLWxX8Lj+V67lK7BCa75buxTk8WrykbJ4mAoEV1h/LsW/
sUSV7P7EHjtWXbA3wtjW4l+imWxxPzYXd1Ztxzq5tOAZ3HbVdKm+9HIgNHANaLj+
donMOB5DbamKRgKU0luk/CAQjZoDdXE0uAPtSnxbeHVyZg3LfPr6kLUvM9m/3Xz1
vE78AfDJIC+VR6i0/zkBkrx61eoZ2lAIUEr0OXto9mSz24SkdavPLK+/A3HC+hjS
656+ictP4MUKXsubuf9bf9biMhumGkJzgbQvFxak5HNsw1SbLXdp2L+3i0WlHyqV
56frmVk9mRdeUqBoYxtrid4FzF0Vpqu5ZUQbTvivL9TSVCP5xbYUJOEHF2ZEImTx
NCuvww+MRddzdUz1osnSHMX+fZe30gilMAVucsGrYbXHvKP9zhQw4URfIAwEllUy
+VXhHKfx/nPX2HdKl5hWH81qiMYUDU3OEyXHM8b1f/EsCjCduFxIKvA66UVFf+QP
YLLuPy43l24Qt7i07Jf92BWSFDZmXuwwSgd1h6Hu7XiJmrTzWnvNSVbkB8EyVt15
ME+BDQlxtrNYP4vEDiyMzQhqpsFoET4Of1ldqMe8g7QQti1fhZoetECtOhIsz5je
RY0ElsVr0YS1odmh9j6LDwgXoEPor6E5Qo2y17YR0GQ3hAzKmq2teGuIBhgp+Ij4
WfK6PvY8yNMFll0Uh30wU4FvNknEfgwXyWaV7B0/YhhG5pmWDR6oH1X+jIz3ok/p
ISlncHWl+5s2kWK2p/M9/feu/24eNMpfyxHfks3bnRVAwdDcJASkJug9ABb/qrt0
9ZcarHWlIEQvD4YHgssz6+hbNn/RTXeohBY7quMxBKaS3k/NPLHmr/+i/wnICMWs
gc34C0p4DrFOrnOjxM9CjgsCAFacnL7AhM5xxb7vzW3plvUIMaY/TeQYU0VS04f5
vgt6tNfhA2sv5ENYU84gqyOkFRwWw9jFjc9YCo+x+9ezgCtonrnQggLISs5U+tmU
0uv6H1gy9PH2GNpj4xkIYocebx6llX34EIdcFZ4EdWqG2/eVoVaGS03dKGCVK5XM
B/GEJvZG5WROePjBDCTl+xTFlELPpy0Ia56o5b3yhzl9fBhGJlfsLkCagKGjXxLd
fCy9t+mdQ+485pl+AXpG+uIxE7rz5qjP+PFDjKdJxZJaL29EZ2/DrFmPsaaMdWMQ
iGkNW7tbJC3dpJupI6B1FWUOAFVJPtIuOMvwqMzTqOJQq/jlNaAbFZ3wJxMIyWDl
euHTB2i2lpwl8zL+wfSDAu2RMtJyCkgbKmpvr8b/ct0lfjFMCou1gBO4A8EILjxk
Vfcu9s6//8eWTuLNUxVvUigvJ/pYYq9Fq7Mt7e8rRieo4XlDWGeK/LNBr7VtKAEa
KDnGv24IOuqiB6OHgO+OOOXChcWZsQZyKDS61EjXKq8sbvviDyIqulGPzPUFXBCk
Q2CU4TmDQvcp9ky2JcD0OjsHxm0uLfDMJmqj+Y9rKUmedywNtlP7lzfatcFbdat5
EJBASWK5cypLw5h7TGdo2GH9DqnGDhGdaVFtWzrfHP1bqknJDDA538Rim7UXDSb8
FstoSdvPCZVcszpuDfScpTCH7XXTCY/+FvJCRGB9MsYyqsHrW6LWWgDMGgi8bkFw
e64HE2T+L9IYYmojeqE1FFLIODI4NR8UsblvfrnNqVKB9v9LO6SlR49XHk8BDtcU
oYCR0TActQ6oDPnNEqw0sKkgO2aUQ9sU+6aA2/LzUngyH0cFCeEw73X2m2prCuWX
JPvSPvqkCqMYYGYRDJoperOE3oLA15IXIlDvNh3kwBCTtdy547+1TmzwHj81kCiJ
euaaYlzlVekemCvPRaSE3k+8ZiaB7bkPkqwgbq0Aql6GVJvfXVAzutXvs73SaC4/
V6tlmsWQphdaXUF8QE8uW4PrjEFByiV45mClaioW+AMEsFKOD6Y2/5OfAE9u5btp
Nuw7YFJQuriwJLmyJuQ92oOY6q4BL3NT9yRsLxaWYNxW5MwDblHLp/StffnSl0pw
JN96hGoVO7B6VGU85CAfnFpY2tl/px2+Zi0abouyYn7EhTp7+iiKLChxggOcsMfo
xJgRFn0hwP8mn9WNPTWA2mktKY06QNQtqGfufZQu5R3tsEzd1Wpas979USsmBFfc
3+CFSRyGvoVPhrV43d0qnyKX1VADOjoVCrrYU+51gjyJqDW4vbnBFIFLqVwkYdS4
Dj2T0KfUALsZYFMv1MhjOlY/3pnGxw7hRVQbysqKwM7wSalHyreiN81RugjS1qIw
FgROZ8maVUqNqxF28gAlqQq5hfGmMFeNzaKAA0U0Czf68V+I6LEgza+CBnzCjhmI
AsLrHXDcNhHYqLyAdhT4A8xM6YlAw/37sfIdCn7s25fRQYTDdgFpK4jCuWtSNKmU
EWbWcwFSFAQOMHFcUZwYIQiKy1uIDhd9owWeALk2VBqFHMfVDA5PE1G9P8Emeezx
71JpIt3LYjKNZxXUFejlLhvn1TUyUiQfp7lMZfaqG0RUy2bjnk1s/cIthdtk1KNh
GdZO060HIqfyqXdhDpEgZIG5n4NXCMoSUDBMpN26WH2pO5ep8sETKtbfVfttHevu
SPCE1Q8PA7JzmIH+QK1E8c75ESwxl2WSlxVvj1UR5SG8DFysBLWnZcB3aXaxaPR9
ISx89ZP5KW56AzYOxTnpnv2jbLipfDj2Nd1Aef/EKhplEi6gPH9HxZxYKYTL/7Rw
5k5a5AR+h4QeXKXiY+0T1L3TKkUpomNUBvrOzx4OkZgFNutS4TnIUIN133DJLhS1
TlChEN7e12qecAVBEGAVsLjyg9ohXbtfAEBaTOV4bFdfi4qUoBi0MRvJSr4oFIM1
Tg/O4VJeG16MUWwS2SQpP3Uen7fMPRGk8ei0mFYgjS9OetzHUxLJmxHv4Dr/VBkX
twgsWkFhvmvs+foG+Tn2bjGx5HaqNH2ou+FR2KR/i2Er9udI0MXhrZ3EyStb/UpT
ucYBdWjb0mAvrnO+ILx4anR9JPh02n/ywCoxyIK8AjNhopCsriEM0PPzx6UOyHCt
mC7u85VcWL4uOsAGcybLtN4DepxrnE2xrUtFdHd9mm211tyd4qbOstktfKKXqA1P
xhLl3sIS8K2l0ADtfsMyjbLqGU37b9krle8Z/RLwbcXZI5LbxdCwOMUjRKXjV2AS
t1k1ACHASK4i+XxeVogJXx10M3jCPlE3o/jht/LeYmbbl2nih3hZ2VK8E48krB1S
Zl3LiIuKeKM8fG9LyEpwcSMAt0sqgN1NDsmVScB3tzLkCV0ksL83Mz8HnCOXxhmD
GrZzEEXvZHzB2gQcTf1TOUWdJ8pomSsqOPbY/IXDOeh6l0XJz2BhodE7AxxG8KME
rT66ZqnypDeisY+wniKK8pM3eq1xgOzTv1X5oQmVaqiNT/mZEPFYdUW8eGgWDem7
sABKsnwOxygBLSMK4GhU7VFu/FgQGDZYLBhKcaiRWCD6L0mLsWdRxoKNr0YpxJA+
E4gRtA4ROyFLiQthqosLhyba/Cf4xiD8iV8xt//903vGzXm11RD/mKBQ1+jS11Sv
plMx+JG0eFVzC36BOy8NCNJwxXGLa/drWEBQB49JFjyMGrY8gx/U9UAuOMWddvln
yEq5HreLzNF0dGZU5giErJ9sVy2axyEFxNx0KSM3gN767HH5fVdi4Nhf5kSP0Fuc
D101+SIKpKvKDii2EwLkl8/Hk6kcX62dHEWrpFzIqDtvFOgWh9Hr57+4e/P/7h4M
NSRpvUd6PEmW1I2244ODXwTIhyyvNNClnpIe/RtTlDydQf1pqbp5vWqEAi53jq2x
x/OrzMzZMtkJ8JVHq/SLsaLJP0oa9U1ffg7n2nfCsh5xQXzX18jqNcveWsI648SH
eC3qloAjcHYBp+nftll/ez38FDNrZDMj6GCT54aspRHQ+g82iX1mngqhigKz7J+t
PkoEyj9XpqGsgI7kT/m5gkyA9BjFiOvVwBg5+5s41NNoXhscyBadHK/Wrn/dI/pO
zhNB7mHGRlyLhvGroO+qL5UR1GGcP1msNc1iUct7UeLgYqrZemdtLr06akwfJ6Oc
BunPWsSVbth6wIWspq+kzhsKHm0+uBYWufP7cut5HkBAGjpJ2yrig9FpnE/poidB
6qQCahjsw54wrV+VaxlEW+0hJ4asDEiHhgexsLAgBhP/qtlCQBZLlSoQBUklT6GM
NWUgoCIXqaAz2FzaF+GUiMnQRszHDta/mRCppPL9NZPSjqAKuxOyq18IKOqvob1Y
NHdIO4A1FJSqQ3niniMUzAI0Yyxbfmo3VNGeYVgupguIcSS53MFC6RY2P+opY2hb
pzUpiUWtVwaZmhJ9Qd3RNUO07NF/lD/qr+s9tSIUI6XX02umI2kRwdaEh1U2UlA/
vg30vaz+NrZxrvc7xGyWxKOYPAP5/mIJMGzoJ6Z+3fxz/fE38nv3S+nKXKBNBJLM
vjL6t3pRHtblHDeAFefAknoH7H3RiXTXrW6HmnSlXv5viAYCjrHt3YILTcm7z/j/
hO2T9a8eyVBnolPi7jkaLmcbfPBsgL/oxEerHgd4OS9hFHtB8im156/R8vo2ed4W
TlddxTEPkKBH7dBKx0hkkEd83jo1f2lq5JF5l5b5T8N9mBnLkeDrbCO50WaJxvGG
WjIYU5gdLcnKoiCFnsR5/Zzvh4gpogtdJ1W3LmmBkuyPJ7qDYO4C0Use7NHvIR6s
foHc7Qg8uKE99m+QdAjOO/p37lG6Sy61zQ6A9rZyJZV5P4sryPHSXlIvNnpnLdlk
cWepsbj6mrYRP+WbbDzY7wuNmxc8orGQhSPBWjcO6yByLh0/mZhmWGgjZAcds2pZ
JBMVJm3l3IFLJDSX8TFxWuwQjF6H0IjFvd/6IwcjteLIlHn5IUYwiGuPLlt9gPQM
E6vabXIRfav6XZB3AlmkGcFC81pYXRwg1jS3zM+44onDWt2at4Wiy6skgtd6+sJV
tErVqtir1Mhp3aKryUD33mLyFe3sfPIxxAvSH+N2yVhe3/bJkfJuIY8aTkWAhsiJ
K6zdLLVrIPqqhp0vso2ElZ/F0qahIlFBlqSgTIICuGxXwlGKnVttGwLYuOQB7ids
yAEozxu/wwwo6ifg6qoEPiK8w4D0b1/fe37Us5+68HZ4y4UUUGmMepBfwycUy2rl
oGl6Blhl1XtkTdQcJn4pEICbaCdzQhlvaFza2J4pR9AzbtTiztizulKCxQgkv4H0
o58RAf5kp0og0jQFeTgWN9zKI31vPtsSLlfIvYHm/PZ5z134SPDw0ZzazlQPA11l
vEKCHS2fCyWq9zlhpo+QM3RELW6q3i59z0yYsj0s7RmICx9g9uusyGYmJbdmLAKa
BXQO9DOlePmC5y85hBZyF/Xblj9fbzI8fFko8eC0UAa6sRBVHBBgVJ4281MD97fH
MQGbqrBJkNWM32xLWTn1pFMC6nqdKe1FR1tmIlwMi31wsoXQUk6opL4HH7H+cAtU
ePtxMK4A04fDpHtXSl2zEkCHTyT7i1kGlHzv3KOCssiGHrs0CGSlrjgLkUr4PAN4
sn6hI+JVnkFQx27HKwyPtw==
`pragma protect end_protected
