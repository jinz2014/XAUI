// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:31 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FKcemiokW1dqMyAIvhzANVpfK2uJGzTQxGvvL0CPHncC0kUnX4M/XmSAT7QCaISJ
+2uqsNhz19C2/u+j558KMvysHq95OxTDkbp17NEFLCzWMJx3ABUpGi3ybypU2XPd
Je3CReyTXegPs8BUG2CXExRZ1KnCp6enTZY+9zrbHuA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20336)
vNAdCQ8PBOO6cemSmswAk2plcuT0fU4bw+ZKc2PaYY6jm6cmgK2iAu485TC1iFLA
VEnGu8IJcqHM38Gq/ogYccqcQfvXJbKtyf0jTmJnvi+13Dtsz5Ff1cocCs0DjQDM
KJ5UojMb0NXegVYCeBFcG5+nPQ25C1BqHRp0bm/oTVwkKcmXGeJY21NdNKcsplbu
/udtUADFBW0EgT0AEFNLOwbnWJV0/o4rbXrgVUIy5WYpfCj6KSrNdeMxDHnpfTZ/
xc3YzWZPBUAAuFZ+FRPl/KiJKMuJiv1xdg0XFvdd6rcegdRhAYKCRx4jTl7FTDnZ
0LTD2/3pr9hMWPt08aRP3LRgWPOKsZ6L7Cmv8KYwHcFSB/yU5u3WsJNj1ysjq2Rb
yVWf3NVMgB1mRWymUOkPBneixnK9VhTpOVUSO9CEHqV+a1uDipJZujTVHMYjd3t1
uGprVU19C9qCEkvyGVqHieKqO+8xqlV+6HSvapqNPFvPBUYOG4xk0xKuyva4u9mY
rAOR2gQjE973SMoNbijGaY59SkwDy3VWjL+cNMGdELoTVxd15He0Br9tFs3jOKXR
a06LiY2o8ieZDyEOGkY04oTcN8HIolAPd1/JWMqjsnAVLzyUock9U2JV8L4Di9xw
+6ujGPVuN9chwIXI4KfZK9NbWJ9ZjJALjZq2945MynmEXpFVu7dphkf0paV/lcJR
zKy8hKyi2g2mVd20A87F1LuUZQH77Mdx8Edo+Yyw3A7KnKtK4DmzL9L2nWWbB5Cg
m6/EXB5duRTzIKxYd/jc8zOM2JvpgEkYkXN+XcaIgDwINsLHUUiG8Rn2e533ADAt
DgF4mJhhEDFbKe0gMGmlMSOFl3e/RcEJ0YvKIVfKDuvJSgGIksto0Lh3n1O4Bo/C
MhR73RSqNNcRfmiGvh8EbAKFMPYMGDVIFVrJbpwwkger/6VVFnnupJxO8NzKuqLX
ZVnkb3iycR6LgwO+z4szG/cpmuj6Hl+0K67l57iBCpOLVvzSiWLF4DY7CiMSaKLf
9G0pes0RXsQjxa943GzQEtyEBREIp9Cix/uavnk9TRKdLGxqsg/AcspxlgHn/NhM
qCiE54sjNQdqamHgl1628CJsrS6k/CdlgnzPLCojSbkvt0K2JuDqEnBRz42qMeCl
7hPb0DTU5zXjDDN7k5j9855VvukMeCSf6UgB/ki4hbjz4kmH4BlTA1UKRqS0UEl8
bGF3t789bFY5VO4eEIkvD5HToglvAgz593G67u32f6G0e04j3LTOgn57DRaMULMd
WkWHODgnaSVoYNsIrAd6qvu9dOwF79nj1n6VlMq/DpNuQb1Q6iJ5HNkb7b/c4TH/
OdVmg7ARYWFHM69lWrHu90fbR4S2yZVgr30YLpz9KucBMUtzQDHd8EhSGQG/PZt5
TuY6+K/6rHoi4lBSKgEINwu5yHay8O58vply94MsuXs3RwWjnHN+3xV1yGzwNfOu
ObPjxsPng4Ie/up0RXD9sfSMRLDIIGq67fJQBT8pFWZ04G4sDDMne4GOUVlecZh6
/DIARgzPRolIiA2XIWo/TQKbLcMuQ1K+rt56XuMQJ/EB53cGC/jd30gCzMwqmq7l
MGpj0ZTtxz5jfPyCJHIytCAdWbSOoa49ClwkACHfTRb7Z5UxEW9GVBdVEf5Qu8e7
wExmxNdv+tPnUbVikRC0Qsn6g7Xcrfr/BNlN9xpnBy1Os4dmMei9fcmMWRrO5Qt4
g/k3s+zMPjhnUWxmoFBZSyphQNCIal/yrVVizrp+krl38UJdbN5Z1apJyiDxmrQe
meYCpMgyGQw3BCsLOCaJyeZjQQrupc17OXWjkmIkmFOmsUQr4+XA5DmpoAG73JFW
P74Ccn2shYjLM2EwhQG0LWvqpeK59KGDfmRoW2IKVlZLU4sCPBTw06g/TUTH4fOm
TYg14O3puJuOITbDm6/2StkJcskh5pRmgCESqqpaKaE0rxy0tDkytycNdepj6MZe
bIGf84HgaanKUH/maOsJzE3+bkp02oOHlFEttMbQa0pMEtavsuvOK2AAp5jjiJPf
bztpC2eeMZTe/h9DXRmu06vna/KflVHfxpX2vz7vRWX6JByhZrvpuJIMLYWhPRjV
QiLqlNKlPixzsBq3U/OVDTL4tajO6jJDOD5b726Ui97DZEmptK/QHKdFD3nvH/YY
hrKzsWapPitd83+WepvOYfH3z99xbl1h/lJ+PmR00YWNyHIlZnHGKYVmDkUcPK6B
8lVnwksOfbumMxPqlSgn+2JMoMVENS7TmhYYkAkhqcIyqKoM3F6F7LY/Szj6tc8w
4yfp/3qYQ7+HDDt/ZN7sIPcdAXxKLjSBOwVbukcTznifUKoxWZi6cXsiBkIrr28e
lKXS2tPGxRGvc0R0w77uCSlJ/ygxr8aWYoWNnwVF6+MV4V0FTaFg3GvOe289kJRG
pDsP1J2G6CbZYSnfyjUFIClx4T6cbi+NOdUFSUGbwcoc712PdlC7GOtu6QQj0inj
JuqY6CNPYgZbUvKK/TcAW7OjDRn7Gm4g4mMPNR/PD2pptUb0KVac/4sE9EjOQr8w
fp+YL5Dq/TAtrqm3JH1Du7aQgOvVWokJWMkUZmungrpfs9Tr+Vea6RE6a07rGa13
h8yCuXHA33DJ4G8PCgV4ZQ5e5YKSCMINwgQRqDAxHAxg2qkEPCm7spyrbIrWTa31
Y5fLQxw68drQNQVVlMirR0IT+xnOCuFmTtISen5FNCZqUe6l1T2ZxpwjSsC40ZTv
O+zNzjnsCta5PmVoX5E0PtucOfCfmnvPAejhfOi1tvjODRE5M6M+4qhS7F3QrsMs
hI3Ov0EbUHM90eMCshIb3Vf/f73KYTj5ZSOmaMs7W+yK6VTVARz9BiX6iTe8p+EW
xApTtWPeu/J2UO8/4BagcwHplgaCYcAwzhdHjU1lfCXbwq3tlyj7lWAH3mrt/nvO
MkbvoU0ruCmBCmd+FIIgPKdirllxk69ukGEjCNgzL+wRIKo17w+ldJKQpi6tTSF5
UO5+JStUoHMLYADfFV4xnHtmpm4QO7LNNQngIOd1iFXZYX9nvN0ADN+osVLn3TuO
FL+7WadbOn9oHCddlLztnPJQaUnMFnlVIZTlWBNn/6c+JAFQUrDB/waF+CXDmx3a
tbgSv2NKzh6bqp976rp83fN1qSoDQAzATL3Ch7F2/KUCnN/+Qp4tYL+uZHceAVxM
Wz6gE5Wh94asw3gDy2Sql02EuXWDNKTey3gC1ZUUYjmD7S6RbwI7J2nDLnHb7nlF
htZGpEgP5x2iPQv1sgC2ANsmnwni6OVP1NvUwawSdM9WuvMYUm1Jc0E9+4s1CpcN
0yrgpjz66QA5cbqMTCxNkC1I8RtDuUiv+J31AOQbume/dqWHzl2kA/A535TGMGdw
fLgeAnbANiRuLZGJCsVIBeZRy7iVevDwI+l5qCutuQNMZxZm7WkN3TCvbvW0mpds
OPNXpt3rhnJbmxA52+KKSZldBflrwDuY603FstXKlEt+8rHKNhYXsQGFEyISYzlT
rY9ALmSZAwtdn0StD/DX70IVJMI2VDIjMVNCWfKRM70cNeG0NIReIVepMUU8KQCT
A3qELzvV07NjLQisjE4JsPPS2n1xvZcOkZkN2TABZ5nInXxQSJkCO37qcoxiFvey
7VQMvj3KvdNWv285jbix3Cd6Ukxmwm/b8jBvXa4nIFrd2l6CQMc8JF6KacMvtJoN
GB9fpeCqT1gmNl3HrIe4VOjNHz8J9TdoNfgqiM074wzvSzlVjFourJNHjVnZ/C7L
d4QCYTUkwnIY7pTkTr9ZCO5LxkAb4t4w8F9yjHiYN3ahLQsVaTRgPkstf3dBwHjv
AxLRESOKHgIFHlWSKPOIwKgSpX0ifi6BSNcuwZuhIwto52WlZIP+YfHU5auS3L8w
+WLB+FhxaLoJeRTYnvNJovDtVF/ULfH1VCcYZSEqpFNw3DR8Cit+7ng7TiCN+8B0
slJzh4FhMZsRYM9qsfx4/M2EUOwj7qvmN1gy+yUXRtUHmLr1qlrAn0bxH5Z6WFNA
qA/slWYN8bGL69DQgVcsNDUPgIqTJmIJp1B5ymDO7QJhfV6R9PHGZpa8x1I1gI7v
viBL9luqKHY9qJPD4N3w8jOSLAnJRp+G+62wLiZU4iZgqm5MD0YNUxoEBA5EO/34
7lCazen3Zmfwpdtfo4L9vF5VxZKq9VKqdf/8MsGxOWWmin0ddkbpKZjqeB/GjMTn
l+9kVVI+/R+gt3saRjKxC3JcHQPMDS+ip9bfvbg3ndsAnLunWFAX8B6JgjVcja2Y
pwB5LPHN2lTPowBNv4B9he+JykEkLIvLgIKTI55g7dQ+4eCkL4K3pOx3UJDhvKlc
QV8yIOl0nqJ3k3lhbLT43WKF+tG6OBGdp9LM8ZApqjL7UPnHOMPlGPQ5qiMdrBFn
pfW+AgNEymUbZjOcRYI3tGHOT90ABx0Kz2FmbPLe631g9aVFWPrXNStOvYS2b6dF
Pg4UHQNsE4tX6EIprL1X6CeHjEAw4mKFhei8SfwD/FvfmqVOO6HwcBN0trrcgVU0
iBpRy9LT42B1cm5JTkaStEwdqVStFnml9A3D1mhnCzgiXwHKceakM9KG+h/zBQZ3
RmfjnKT7f9WQ4gHWikTu6SL9EbO7TGhF6iVRHksKL6lqhNSugq+LJC4bqrVqRrqZ
znUX0bx6KhNjgkVFSNp5NrrtN18/43PIYbaLI+tn6Uz7ZgYwPOEj3+mdpwvdN0sO
kRTWstMompbNuBHWH7SPbREJLZAgbuCTinHZKAgOZNkfx0dDj6LcxQhGNZB8aEWu
5BYnuSslQcWIQetJv/SDeIUpd0M573GGNu1igh3R9mVHvryZY6i3u5Zt1QpLqigd
teb8BCesP0heycbOY/gdKmtUItrBjvr+asnpHVgywos7LtP1HAcIVgbZqDO8RtwS
vjHRUvG0ovhzcMhuctv0rGFMSR8v023QayvO+IDflyFkdmmnGIAx7X6K+9ddHG+h
6a9F5nSTouom9MenLjwtLOwxCmy2+t5eW5xCHNWNS6/zrnGMS+ttEPgizDq7ESLW
uQ8dfo1kf77ELeh9VOHflDqOPmjQjmN48BR254vIaQ/2xm8xO72bScFWrI576IU+
NdvkkzEFHE4tJC0iKJ+tkhvU78I8WiNUsqh8egAHhup04mo8NSZk7lEITy1U8zCI
fdFY85LshYDR7Sagjo9LZ1IfRcJfyUuF5+mgH63HBbg35DF8/3kUQRtYuvaSPJ5J
lqgvbls30j+Y5G0sL3Vunn970fmYAx3TpNgK3KfV0iZ+hpwFO/3OJGzphKq9gbNw
k4R11NSKh/RycSARyYHL/u/1VIfKfq2NP1ccpqPii3LQVwoTK5Qpi4sHNdVeR90G
KXujNYVIpDPqCNQ93ikM52G4Q+OEX3NoxkxVPEAduErevV5Zm5EUbNlZByGa4AdS
kqRjNwkBVBrtb5i1aKYq7vML4EzSPjBzxHicJz6XtIAL0iBtoVK9lmF33Lg3CgUo
MzYpopvnwRdVH/MkQTGIvaHAPRN8e46OKdW58fagf6eWFC2LCFXU6oSP0E66488w
WuFkufVur9R6qQc/xtmtUakohrRrtqZxeBMpX5kpf0pqDrV7/O8/f1RV96lHyA5q
56olk7UD11bdtqv8mUD1d/WiHP4oQyHOqCgzn1cQyN2dvtnGz/i7D1i6goi5M7Oi
igE3Hq5Vku6H5ULVdaKfQAZTvO+B/e1OoDU6xXgZ798e5UP6izJzJjEuv5mDYUtD
m7rILCWZo1dn9H/UOEuzn6cWo32phvdjN870skQAydKAwOA+qVCRLOB85ZIdlX5g
YLwmamcAMRVxcBe+7eOeQy7BA0ldKbk5ex8poMBdgAGYcXvx7raA0+UNu9ey/r/K
AlPjoWIz5V0XK76ITRtYnS2vXW6hR8u5PDLgFmdqgB9mrlGgvOVrbzc22hDBweOB
zhij35J0VGRimM4w2M8KphYZcY5WJRpqOM9u6dvoUqLINrTB+kZ+0nt99HZzygkX
gbHQeNfN27IW7ByZK4RnXhQECJI7YDL2AoUVbGDwQ8mL7tsf47Asl6eVa+fGIRbD
EQ8VSbZ6pCWhfFsGTRDpn/4K46zNkEKnbZecMXwd4Bfb+l89kkWxgyIxxTUrySUs
0VWOiLWtRQWvm3sFgbKQNxIEisUrvFHy3SU8ERORcC6AvjWo58Ebipe+8w0icVMF
8lykxKgLGLw6QS0LJx7UneAEnz5KULNd8H6ZkK3xEDSxMOTYGzaVE+n+3fbYjFgF
vtBEMFUOg4imyA+ATt329rKlBsOU2nuqpdyfm9et5KNcpV77PVu2v0ORb1VLJQNj
UEmLYKNieWNxF9wZngfS2SPrBd/mhu1yLWzL3y82swCOLlWNc3tf3Z4R4VBNlFOa
59tr4ysTAUFhPz0ZDX8kdDLZByCy1L9V/5S3AQB+6ioLVU1lY9J4vbJIrzpSBoJ/
wMnKRgcCEeb0QjyXeOQDSLTJLVrFl/m7Pb9H33hgo1ZS/yaFHQqIdyYt6ygrCSCb
/CPF8mWaYbRRtvx9jfY0xD6HBhatLBoOOzq+Z2CxsnYuq029yuXymgmZErD6VFXV
RlI7PxFZMk9rW2vuTI8xFcjS/CJLcR3QIqZKFQf92biyfZENX9v6CJXOchgKFxzr
ADr2q/DYcr+QmWnNQQA42JKgp/BQ0zD1lRNxnP863EFVj1xbje1Llopa6zsbqI+L
i4Dr1FPLWT2KkvkcvnBukt27Gqgif9PSUNiPM3nhadV0YDpNfAzXJBNteCTGqdkt
i3Xc133F6wNPsgj7uiM0F3voHRegl2NtmLj1C3bbZG0+5tiAQFvrK1IXSVBs7wew
njqOOFaC1KKyhYfTL3lTUnfZcvMSqmsu6DfhEq2IapH7GZ3Q/0nHOQGRnJlc92Hx
X4HUFnJCh7hgiA3n4fsr83aNJyljA94HFyVDuelq5uUB1/ll1tDUXkffSGO6KVuy
Mf6j+aEBguOsZCX++5ORjJrsNeB+JMJDfcAyE5BALf5ZbcQwu5kbwmgO++2+lf0L
Qy7MWlBanKtBz5q2a2YXGqFgeoAqLdSCQ9C93M9IH3VEnwD05LBjDqyF+xyP4LHm
7CRUU4OLG1vlb2LjYTd9gr5JQzxb2+Kt3AgHY9TAkKlUjiSyGuYPdaVNhliZ9NY4
JqYd9bJv0fERCLcjrSdAw9IWR5rVGRDyPXTB2Zg8KkGzI6+rhvq2aQDJaGEMZPBG
wtORqxLEINs0XOSw39X+G4x/ijIA6FQ1/JfCIHwAMBUIO2ndj5+Kv6KzeUsSVcbx
xP03EaVPIFNUj9nOVZsNW1ogLeGsPUPf/jT1oC3NMaBs/D/8ZewPsOEnnXPgIbPx
5XPG02NOWG7+htR9tyxvdtoF/OrNIsZxRIXfL+4BtBhn9O5XLqTkNXwC9ufdQVAX
yqQ8dPfYPlwSXtxJBHBTu8ZLj00YBWke4shOLC1gTRjChuxlU5d4EWGan+p5Vawa
mjvY9szh+B8WlyLsjg4Dn15ZqUJbHeS2QTl4c9yyGi/79bGhMINvcshvwgG0SCpF
pCKAjD7L/U5WJ45W86tog5JbLM2Ivg8Xsa6NL47lo4L4ApDYPutSCJ49K8MC0snP
1ObYgNvYUcyCxG/aJGgvy3Dlh5t2Xjlyp4DIu67pfcJ6Iatozh/Zt4cMAVAEpAk6
X11DmnjhvX04CD5KhCUb6vj4pXtG22CR6qzdSRQSEwrkk8Ip+nBXPrR/eQKzWO8A
s4eEGK8C9Vo62QtFYup3OwcE5Xkpc4UM+OJ3Ps/IU7OPEKk27aC+sCGqTF3W7tFQ
FUKKuwtxMWs7zBxvzZHCBLNqGw6fbEe4m9fdtOnlmgZmcrj4GPMBpoggnrfIh/JO
jbsrE4Fd05WORS0wBPWplIt3Wa64sNDMeAzTNGZMyhlbMzJ9cYKx8sEJkgb2YWLk
OK5bL5urHw19xqBpWGYeTfhFr7mdOiz1ImFiC1Bu8u2rt9WJD6gSiD/5zNgHYygp
5txI5AD1bRNBHlZ+WLjh/9apqu/a3FSW6FBnqS3eZ8elsV2qok6j37O3rsbIeOXf
C0sKxOyatcv0pT1Fq3BRnAXyDnIqhG/F0IeJ1yqsAS2Bj6hbd8CytuRaUozEEy8+
BlnD16hW7/Tyk76KIqkhV0FyLFdn89swphhOQRPOXbYxPBupouahbn6KBr7SlJUW
+utOftQSX7cecAZbRfGJy0FEhumRwFRUby0NLaoNts4az8t7v74gTkAp5BfwNsgn
FxKOnhkbN22fsWSSedhRQRHgASrkprQgzv30dL/skKYEE9Pd7xq3vrXPUq9KzeQQ
awPJuRGRJwak3L6nAuYGwmbwml7iAbZ1YRGOP3ZvdTvFqofvtCmCrx9bmed3lKhn
+qee0IjwDAh561FnAbdPmtMPYhEnzT32ELxImaC1DY4MsM3JR02BPsb8TbHdsjgN
+EZKjR2qWx2mw+/owJ6EM2pqsXf1YR7M7eJ8EC9c3yw6SsHyRcvgKJe/BNv1HDwM
a1x0Jwowjj6VAgA8ISJdzCouQ2FIyo8JbxJXaqnmVWo3eQ5CYZ5OH2qbC8LX/J8v
AuxgHbHcS5eKwYchZWyHGDFJnOGhfiDCHCTonqJFNGLhWX7Bs7h0nPxGIgmgQqfT
Dwv67Dl7CYyw9vnaiksdyeoiWzVoaOnBhRLCflcSr4Wwvlatcf0NKqBld0IWsPVj
eI4OpESuDICoWwHYbWLLA9DvAZz6Tsys0Fq1a8MvrwTOUnAmnSwz9NIMNUNq2EvJ
JY9amM9M3p3GoXd4JP9TFr91Q9L9+x1ZhZJFttrUXGE6QO//WUwa7h76OLPHFCLt
YSIs7U9HiGBoirIbZSxsplbUC2yuvXg4CoRkrV+Rojvv6b4Xs8G3V6qIKs8S84HL
zj9+rQrudr6qlLmgEsUh0KbF21PutbvNGCairlk9yG4Q1TE1XjvzKoF84c/F8nsY
P7hjzj/PiHRh2jy/QsTbBOsbBmS10xVIeZTtg/mzXILKMGFg/mtb6sbN8VVTE9qQ
aJERHRfjrODR03aCPBK4sr9VGJfHdyBgvySh4MeXgKFIbwE1TgYMQvc0KLUgDMvo
4nXBug7YvtWOtKQn1yYqfKX8TcITn0SI/RCnFoNjN9qlhLz7U9I1MsbY16vbRBCz
Irt+CKj1XsCake4ixVkojKQLju6FpUMmnNtdkdYhwml13OCU/UVoLVG/ruYVg1K8
sY5mY/AXikCK3E+cdfvKYkLzed1c/KAwEkwjmlXUtr16qI0J8kSKDSC0gMiMPA9i
HDzbmCa+xaDIjVwLfsr5EGJ54nVRMduiO9qn63SuyKV+EVShoo+cXP0/f5hOI3sN
zVMNFz3gD07trk5Bh/Uw+lAzeBfg1MUljmSOo8FLzqGvc/GsaTEAoweqpi+BHezB
W0Pu3QPZb2n6OcdGFNuZGKDkFi1FIoGtHe2Z1WX/kw3oov3OjBmYcIU8f6/yE3EE
198j5CYej+T8KqVP8iNKA0vJBmsvki4RMC4c5X5MegsKPN0eD5sYUPJKOgJBM411
4aC+qxsuvgMteRJM1yYqLt0O8eRpHhoAK2lD/K2Ixkp6VZIC5pDfOtHzmXfSjVMs
8XidjiD4FRaaE9LXM5ky0fMkQcocGJES+DePB6OC2Hk6NOCWa3iOUzZFES4UYu3C
niSNP95WWvQLbi4P0y1877jJIIRI+DL+QX+loZm25S2ptEr8XvkbFYVhLEMakpQ5
Sabc6OX97ZmxxpPBz3HjQESAg1aHxihy/orlcR0CTMN1wUM8p47SDw+y4H+wPNsm
ZzctPUCrvvqZg0O1LM/+TArqB6gpWkPJ7Dx9aKjIzg6DwOhcDmF43UDib7CnltsA
PQXzkKqcwexi+c715eXqMlbyzEjRuKPN7eDSLlE3qtcgDRgtGhmoiqHTUF3PdInn
oPdvwJG/LtgaezvDWQw7ugH0hkMnCi4rGkUE02t4Wj1af+rSyzLy9JVHnjww/WS2
wRZ08+9WY3lqchV1mSTEvMg14PTtRQoPLztVJ1pFuhBbog/GMFuASg9R1j/n2AHy
SCDk+IkwUCDYtzdKEG02pL1lWjmQph5BSy+lZhOr64UeCnBo2ud/vqHetso5hl7W
NXvN0PQqWUJmn0AdZxh8vEkwawAvtzR3g/fs3r5/E+yDgs4EW+JpvrDU9AA7O7S+
WAzz2YuosyWu9n1I+Vxwi3WTyS4lmkZY48Ep5chjoaYdJKqhIF+CUuP4S00dJtCv
oHWjXgpVd+fu0gTre7NVnyC1EJDbOViK4dgJ9qwGH9wnJ8HI2uFBTY5JSj2b4++0
T30umqfTkQkxkrRg/fFUR3CmWpmzrvOf3IIv81D/WG4f2M+sWKPsxR45aDiuyris
MlHsri/CFdHdAcdXl7zrXbl0V12J1tGygW1cVp2mUPx/j5QTkQTBsLfRohTOG2Cf
JoRyUte2ROomd1J0PkpfrFKYhugfCBPBUK066CYyADQoo3bp2k70c5tsqOfkiVkf
5J9UbUBBtIbok699q3qntvDn4ZYsqsxjxK5vk2urk9Yg/Eon8TUAztbPhbGtY7lD
6fdMX8wRS4UoWK03kPOsuRGEDgfR6vrrbVYN/qpqsLQleHIyI5xH9b5HbaNa1Zm3
pkhr0Ucy1Fqxr6lGgxJLEXXVbFaBk8BRk5OrsAf5trrpAVHKq4+k+jU6VbzLyIYV
GHceoc1HZeURn8uT4eaE7CqOraLLc7OXC+D2u6JSwj8YKg8Krdodi2o74GZds5Tw
en4DW9qqxWsceaRX/dNme9fSD+EP5FFE6byg2jiLosCTdsgoOjyHNK7Rz5GmRb8n
o4ne6DRnmoO23RmJJ7NX2YDNo4pwIKKe8Tgy4O5eZ6c+ecQvbi6uxuVQ7Wgo+BGu
wmUvQjUKaqXyX0YBb38rhpEnFktt7buYHpPiwWfTN/5ijCVpS3jXnSG77M1ufeRa
XUXORr9xQHx9qFu8+ImkoGDwSj7NGppK/2cJAhN65z8jgS8oLO2b6IqxKoQ8da9p
PrtlICgNJLlsd/e8fIv+DGReSX8ekZ3pc9Bo86s+/xX/k0RIZQtJkfl7te9RyA8L
Vl/LETiZhdu5v/Xd7KrkcrzqoXVIc1fO4ogk9wKut/44+Ys1ZyuEXiRjRCdrHEL5
V8KshWPyw8aBuAX6+15jJ2k53ivFQC8XfWKhCgmAlEZx846125XMJEZlP1wJuzEy
arU67N5rp7hK6Jo7FdOGbolJb+LsZy/GQ00HD4VfOU6Xz9xwU6r+Vuky0Hd0T2By
z2agT1wq61RDacK8vaTOjVg/d7yr6xyUfTu14srDgFWE+DdBHHE8KRQMv9nC9PeK
ZkQSJ2EFp8KqxwyZVnZsMflpXusQ2lXIcr+LeIl2bM448cK83NVF99eieOCz3Bko
hA8f0tRt/ZXiIM5VLEFPYM9zs68y1ZDqvegiTDO6d3S87QZX+5YwXMYFnNoxl4fu
taasXby35mcJxnAotOZeDRS+F8Wpwv5/52kx3Sz4Aj2c0y/Rh+mMzEOr7YWblDZr
mBr6a7hAZCYULj/Ta8DS1lpWRKTeDifE4vfX1riAbe5wr5VfDeGJFM4375xhSxuY
1qzCDN8+hsL1DtZgk7Qkni14O/5kgu5YOKCVSjgvTEvw5esNourdBJ/p5lOi0b+G
R8NTBUnezDDxID+qEgGm1r2HhBnwm9mNPfkuUHP7ZHBK+8oDoR5wUSECvUAhCPzz
GdSltw5OroqiXIJXgjW30+vZJiN+zTmEYZUdyscyt7D2dvcgEXyeBr6YhkeqRoUN
NtJUwpDi/xMOaP1bX5UW3HjuhFzf00hyL0r4f+2ZwEkBtBlyCwsyM3ID02Mm/y/U
cRui2W1AVKXPdZaWtcY2nX0bjea/OSCguZjR2eSgh0NYFi9GOof9SueWi4MNi8+4
mHwyBZw0ehteaI/mcMn6Z3+hoptA/10UNqiSGPxEQ4Qfr9aaHjGnq0/I5Jtkpp+p
pXe5gOu/Zpc6Z68Y7WLvXpA4Lx0oyqXfV3jfcqE1iq5y1/L1DA4Xj/H4b7E2QO9E
zZ/O5F8uVuWHzMdjLyUxOwscgAbeH9gV+nQQMJwMIXddp5ZWd9KVlGVe2hg3H9FV
QSlGtyUTpiXsPpR2RsjNG5ALzoj0+5FM4TQPNPQdYFH3CfZprHqShHs85BBw+/Bg
6p0EDXRLwgug1GT19fsuwdDRZxU0KnVcVhhpacBgy4TerFcvVlKPXB65HGGZ2KaV
PcyulJtgOkZpneYNwciWRR6TMEhHjXUarNaGos6xUdIK8lAGxohPEgntqp64mvBl
Qfdb4PCPwK3VPsoGHq0YzTg+KMYasbGuokitCp4b35jekzUho+/8yzL4Jpv55nRC
BGg1zzL20pprScpUkdMGr/+huKA6rWKOgoLIRysMd1cLj9zJLKvSSobrikYfx7vY
6bOohUcK9n/DQeLTFNQNrCauBqnxPb9cKjP7O7qvn8Sah/8UYDfp21gJCZEKokrd
fZw/VhmpkzbgyhTfYG7N8E1tZXTib/pmqwbvYFiPbkkAIAHHdUB3EzP2w+jn3xl1
QIH/8bMqwZiKmVV21mxMWIKNdy3M5XquqhiFNMpS6lvTow3JJtd13YzULVtnW/3I
xc6sg1kZXe+X5YLB4nGYDNTPV7QAB4Jyb/aBdj5wYqAOQQWJ68GaSjwZm7QMHRBY
Szk0i37ahw6nAvNWbCgVvmA1A0IXMsvK15smtdTJZYdYsKDFU9NVmAWqqysYd1D1
y65kq3LwqyZMPIV3/+Y+cylbj0M7LvbYxdTmguBQvismQQcmQnom2rIj2yh44a3U
9afAAT0+IddA1tY3DUvup3pNeR1MKjE9lJljsfYPbjJmIb0rr9pojWTaxjfbXQF6
+5gpR4Fst48tOP2N6if/6chMrx6BgycLCPVzzBVXKLfq9Ql/XjzQkLVAVOEFrT8P
ejQTWtvvqlYFtQ3yHTlZwwYw3UupR2CtNnnpJsrnRTvYuHAULe2G+xJHnOxeDfFV
indjxiFEvwZK49NBXDk1fxYv8A+hrOwb8tNPqMm8OlDjq/Hz8pm09zH64Z7svhuf
u3/3fPS8RKeBJrynnL6Va8w7k3PfjFZv9VjDi9fPCB4BLTArOFXm8xDvfdnZfo4y
o9GA5N8RYt+scde+3xPxSFe3L2y0c8Z6CU5D4FPv3A5OEIzx3tF5TmfmvdXvmpnK
jutf3g3c/+y1mmIoCeurxAxn6/UIZ0DvOLnwC/MWV9YAhVD9aoxDeYmTpJci6iRi
vg2OtuFH3uVZDurK3WhtLK38kjRBOpJdW2/6pnM92jpu1X6k5qi8j1OWREa7p5vq
UEFCgnqXjV1pS1PKF1c4rlIyk1REkjkdSifqqHeb6XrJzgb1URC4CqJTEwo95ibz
g1Oo7l4DUkqo1PKMx4OiLEIJSVe68Ff0om9UwCLYJLISCHIyPr1rzJfb0+XATjkg
yAdxbhYU1CiWVXbjloZZCrsXlr1QlU0NSqKrrSAxgTI9C0NkxE6J474HuLfhb67o
RUd8OQhVDcQWRI57D9WFjNQLF8CxJ2gRjM93Ds/rdWPM4pv/FlMJQB76z9tyE/B/
uK9wZvM/Fhy+a0ORNYy4eqB29DT/PB4nLtokm71o8wUdD3Ob69m1XF8R5KEbDVNh
dF2HJ/KmsfWcLQSZ3EAGaiIK2yKt3F4Au3MKmfn7BM63ZVKYl6+oorPxCkH02QiK
AqqzU92QxdZXDZ5x632W4yLP6pCNlt7EUtGhyWtLkxKMchL3iW5AjqbnJJ1+dB3R
swZUTfQbVD8DWJL7ZKxQu6ONbQsSb6ouEb7MTIQJLn8+dw/WvIDw9qyDOKPZIfLe
ZfsR+PjMkhVnQ8/gJzhTIzSHqUngYznBPhbl++P/ukPMP9bUWfOzwfglA6A5Rc2m
9m5M8Izq2dnyWzC0CazQJF1FXJEPiladTiSZgrotkRQbdrKddtlV1qYqHttY29fR
qXKDhKcGgavA0L5hk/f47ddx5UOybH2hMuo4pVvoCT+n1aJWwCQvL91Vko5mJ9K3
zlIzMxIW/niPwqpsocdfd8v4r2aUV/QRNNcH9Zyem9PXjq3y6chTKqtjfKwDLYx2
hDVs6G5qvjuEeY72E0JtZXT1VnHBNwjvzzpP0/aR8+8INwl0BS9g6rx/lcSuVKX4
WJ1Yq2R2M0i8fnSCTHIpmbDFxs7tUzgm8zAZZbEUDVJ1+Jckwv+mVoHF0bANgBMa
iAyALsVsTnZNdyUeQidP2q6VnrEgwKNEDV3B6Za+ViSJYHnD+IEZ10qFmWgPYN18
gl8gm5xV1uiOMlp7vFfXPna0dSkBqg4sci/dlanhAUGY1CM4AYOBCktPMLhcCz5F
gTI6Fw9eGZoSx+XF+NvWQ8AdNxPtOSyncLJxrPv0ofBrttbkFizZObvh7hWcWeZc
jPSEes2G0+rqsvQD0AvNeUbPhn+53hMOZXPzw/cmyI+LLhXBdmeE+AhymXzzCKhZ
NHfblRdbsK6Ath9K/cnwJEwdA9/lAka9b9sACVJRUT53htBx5P292q6NAapxU6X2
iD4bv7I4Kf/nNZH/U1dJM4B4249TsE6zLDK7zafhUxS2zWHBve0BWf8CO9Hw90Tl
6L7y53NQAF/Lmjq7i7XJ21ykR9YAzV9KoqBCspBGzg+IUBwDRMr0HQRx/jZiCVLR
IIqzZ/PA/KVmcL4rbx/7bPpa+Gm7w3e8nJQ4QMobWbkGrnLSHWNAP8P+sXl18Nts
665fCkTZNvMhwaglmFUoeSulWJUEJg7RLGL/fN1f6CngXjnPd4enMzYOM5RN2Lz2
KyyuvSES79Adjh3isREL8/nWjIBJ99l04CfdEqXmQiF9/UfVoEunFbYOhH7ogJYy
rDUX8Tq4HEeGuXaoRU+VhlFQ8cJrD7aip7pNlFtroRai1WiRsi8LSxCazEHhk1Ke
XzBu/5D2CjN6xcCCz71hMBaKBNcdpBGniUNX801S8PISkzEHF2teucxBz/rUlCpV
0SdkLIv7DahNcVoYYhMdWJTSt7QQ5sF5Hf5L9FMS/xeo2kDJqKF88X9VwayZABxI
dxyUsuxdXY8amlTAKW7Hmu3UlTZxnUEMx4jhO2V5S/8XXYw8aZxzFFRVjsnR6UGp
1HOTdgYY7F5Sgnywt5VBc2a1/8NiGXQ4bFiv7dUxhAp1PCVbvGZQVc+itb+VOXRZ
k66ulm1uDBCSrY+LLXGbdUEPB6n02KiKdg4UQEV2hffTFEimdGcrHBilTCuBRYwd
D0QRQsKwTHOk88DULdN55VX7qcy6L0z8GGIYxuSLBn3+z/WzGbYieWKBNyy8DVN3
X4MMU7zFqwJoKs1YYwGy/ngYJ+J6pd8yxmbkvhc39R9X77UVokjctGLRrOkiu5iH
x5qQAuIbrxrMgUL4bTvoRXWnJZC9HpZBA7+Xj7eLs6eMk1z1//PbrH1UYOn0DyqD
cXJXXoE9DDGbhkRWzPZzktz3CloYrH/Z55aw15N9qaSzQBw0Z9HZFfA8TFAEDtfB
VImaLNp2eT/eaKjzgp+sCNvuRYIYOX2jIrvaJabh8pqSYYeamIBftziTZtxsME2w
EDvLT6Qd4/TlEMLFihrk5+suJ3hdSR8jTdIngryCfiDWllBeOXn15PahbkVJ+TEk
wX9WouAVA5HIn2nL7hbRgNT+f2ZmiKsjMEWh4l/U/UmdklIOqTyf9C92K3vpb7wg
EqJCrFi79lWhTTHSUoFiC2+y5CJopCzWDK187yWVpoORhsNqXLYj/oj5+Lbhrz5N
6o6ZciVq54FrJ+fppa4w0eonc/dCg5L8IwO1SjdfnxkE2rCgfqTs2MRVWaBkdPJZ
hL0rDC67nqaNtKRfo+ClQ82HGCm8N7ki72FFHdTvehbhtkOe/HA6gpnvuj+4j6Hk
C51XksvB6Z0+eV8kgT/y2QTYkR8ibwc3fFUM4hH5ts3WuxWflGeBpxtRgIMDDKYd
FjCX373rDCMYQCjzGU9gpZRdeIoxjyI1OdmpkJ1AbFBI5DX5w1/ewwwWG/B4v8Bg
dpbjyeZ+Mq4/5Uz5kyaNbLtqO+i5uNPuuYGrE7k2Jx9dr6ld4evsyUUwLKMVZ6xm
kh6L4MPsXdoonn3loGc5uIUV9xHC+z9WfqGmnM9oQhdYXhI0YOMHesWEcgPVyzhC
HKGLdakVjTy/7IDO2xCpPl4aNRgTSEjKvYMtIrFkIwLRVZImjAx//FirK+M4EXog
D7PWOIj5tT+NdN/wpwSLc8hpYQspkiSnCPOqSkiL74VAqKCsA7t6u0Ffdv3RwhVo
GRd3XHFSfqidQ+M2IoGWPy6K96D0J4fsTMP9VVCJSVffzRy/qmmjPl441C1wSnjE
9Zhdl59tCh4LRptcP8y3vyVCFdQJlLqGpOPAhAP6TNRQbh2D2guv/idaK4lT6hfU
OgcM76UXKXUcdZZIWyCtUhUlKLj5MJIV895SFgRt8/v9pOJtGD1KDwHE1nTuASce
+Mltg5IF9F+Dd7jbYLgt9uWLvIu4tiYcZIgNMO0RbG8ONYL0+DOtTZacafs49S7+
klXYIEWU8/4ykyYYGba+pcHZNXXQyCj+K8SvAdFQ8/jMz3TfYXtoZ4x89XU2DsVu
Fmshg3euP1BUg17LxUD6FNt/Vo10taFpbs4tCXoqw3VzLjM0d6TtJKbC7pK9zrXP
rzKISE1/+bARa5udqnnxD5eXiF4JgwP9upStQ01zpH/fkKW2S0dPkmHfrzkZ7/J/
xf5qd5ZE7MrHKOXVkhyqUD5teuIWOfAk8HMRUvaxuwQC3h/dBuMs/TNl2nVw060g
zcecMBoYAhBR1dux8okHTKC5Ezh6GwtoAq3AlcbuDzHWB9OVXEvHMlo6T9oNhlxu
EG8LbC2QkDTOMoAl1hZpc4fPn63VqCaa69q8mraOGCRQCTAyweXtsMjwKvk1MOuw
zCcUJEKYfhPDAWuALfY5IjFAUDVJYnnJ3RN7jhBfWvv6OklJ1daZ0trkqLVoL8C9
pj2gHr0HoGNBzJWv3pSoOoORViD90tc9Gd3I0J/nBAFwscgbfHr7cNP8cVb3X6XI
kkVoH+L9a5cYkItYXummMXYUmnFmkt6m5wMfk3brIZ1HB7AEb8OlMDRBm9xmzXHC
sMGDTOFZqOyhg0VNxqZasjcNmbSqAXM6uG7MyS7V9m/AfPJujwN6eUN+ndFy+5vt
lSkIodLtAvrTEMlIHjSj1bps+Nw7iS70GuHqnjX5BK/saoWuZJ7Ae3YCHxL4ejgp
kHH5KxsUJJwYbw5tC1Qazh8cUn0KEYEtygbKy16jAhKK37WP6z6+36B83JOgC5i8
/NeI/jUHssEgNMUFMBGh3FziotW90NFn1dQAqNJ4EQgPyTXRiiWHKW2dYNoQHqAy
Rbpoyahi3YGuqYQMSGfzQiNWEjDISPRrKpsk3LR7FoebQYHMy5IxiitmJrMlAlMa
Y8y/cEAv6nt0N2577RYPYRDiR+wrx8DDiKipGbM4L7fVe2gZvD0FI+Jj9vE3PtFx
iXIAP69eiMVlHJ2Kt3OFUTzsZXrqi0LbaNtr/sJnmajJ5IdvMSrM35PFWxbLGAWK
oaBu4nTqIhlpNnvgdkjWUdFX826hZyrQBwFSIjf6QngsYUrQtj0PxSl6N8pdEzZ/
sqY2IxDOY/Mz2GKW6lD4HL1q+4i1y6hT0mCxWZyiVEOfd3CwBfK/xSjyqRul60gx
IsQb/34zCMni0liT9trFEXed2adzNjBk/gXTrHJ7S/z129soRnqKO6H3XApfU67X
kNk3TJd8OqT8EZCT3vKF4P4IQv1eUFST9Fd1K/G+FmNdAfSht5gdM3gZIV75bLnR
Cd/GOwcyKtNhnirtk9XLDnGoSEuwVZJEXCTBgVePjZ+LmHPzO0wlP9arK4F1DXan
jRrBC7E5MuQ6DPcKwZHKbQXQkuDkSaloQY1TKye3jhRx4E0l95mc4M40xgvOwcja
jFmZOSOCr5wBrnbDYESm5yvb8yNMbPUS+LtbwqQcQSNqwVQpphAVBX7TeIXw0E7a
pkKZdRv1v8mG5Wd3827lyii705bkOHIvDP1JYWNQHbtxGggBE/weKHlrzbWQPW1U
MrbKykcXLLE9n5R1p1li8FGu5Qb51H0LlsVlhjwhTiAIK815qQ0oegTmvoFM5CFu
TitmMmDyVdoN6kwZpEph8LG8ZTmFkwPUhqbwMTAMp147g59ySWcVHerGKXW7T0Cl
hOZcK6DYwmEziHBy0H9k6f6ee3AdW8p8qQNQT09feXU10pj9Fe0NSfxgt/2dlpxJ
o+3BSO7AcrARsApAVrK7V7d6VgtgSTEW5czmMHg211Gx8KufHhmS81tvr7sn+KcV
AMNrZBxJrT3U1foljt34l2Y6OKO4WrDoFqJSQnCA+MH69xQdhjZBxvUbZ3gW/BPm
SdSiFFIdLbi65jMR5LrPF6Mr8MUKZ4CgcBI0+DXGA0RGrlHdfD+5azvOa1Ngz0S+
+c+dfcQDf+umHbrVbrIQvCBIl0uSvxRTyqGi8zi0nTaotud5hIyF+qdTefvqbE4E
zFbG4w/o7KgDyHaI3lxdG9Q1SNIF5z31SeMXro2hVre4LHiiMG00rw7rNoVJUimd
uHxfL6Vn34F5SEb+3ZiBmgoZsJDbWrLv7Ir34+rzzHYlnVAqxT7cNLegqLeTW2Kq
UkmclyXW5pFXNr/UdXqz8FC//ES4xh6HoCb2Q1Z97HmjmAMoYWIvhY0/wp9ASHEN
CkhR7yNZ0e3TCRh9JZVnsHw3tVPPhSlQcYszryfA2dRxRvRPl3P7wh30HtY2D/2Q
mDF5QlaM7tVl9l98nUzk4aChlYZcf8DKZEvdBGVQHm/qOVJ0DNefelFIQ35lrNH0
eGa5nX7iXpE3AGCopNCoz+g2qDSITNXktbU31H2eBRazJRdFpYrYZTD2aPbZal+3
eLzJzWBEAqae2WDioRuChOdsn5QlSNaC071sNQEIBnfdG+MJdTvJ0x6kHn00hK+U
bhAE4ss9RNEVmLCNEK0MI5hrzl0wPpOODSnzesJKBtFuwxg5J5KIKPFgD58EXEs1
HG3VdClbC6Q+kULTcsNhvZuBaWnWkPQBQtDG8iPT8j1itqLfBta0EtrZTZLiHXKg
Zr8vWoo2+Pz3BuJjIjIRrbac+xbD0TXvV+p6OadBTXbxcqlcdYbuqhTtrMm2AVnr
Ilodq/MVLYZBmp6MlHj1jR5JPeYisvhybyRj1f/JAkDDp6w30LLyrnr9HVUEABvo
2+E8OmYpCqA9EKhVVBVdEBgbHNCVtspWFt1jSJIdpIb2KylGgVGWfsP11rKt7vGb
/D3n8ue1vPV1kF0mAPxOX1dtbYls00GHBwoHLUhva+K2d9oZGZgyVztg56oljpzh
KX4yxugt08ul/WMTRxj+sIHJUfSMfctTW5dmqLX/KlS+UiuZawmenUge4IHoeNl0
V/CptoWPorZJFJ+di90Fvkj5kw9vm0bL0ETd6oISPUQfxMqbWgW63PzIDFYpJ5w1
J5bLM/tVxYfytFXtb5OBcmYMj3KBf3N0GDRQfsWbYc/21Psq7SBRSlNn+/Kbyt7k
FIYN5MXChVn2npMKtUKEmAgrdAoC0wenHpnH32Ze/IeW2yM7GryEabJdfgqV9Tz3
5J9ffRN1z4hWKMsv51Lpthu/KHQUkDgIgW2cg9ZC2Fh1Rfw1ieNQjlPpr2F50oUG
c0xG9MEAUy/K4EhQWCEH4T/qttJ/XufZRF4xs5oSRh2yGyG2tdqKgN8Xz6d4s8br
x9N/7dY9+964e0aTR/WsVEPhkaSlyjjSnvkmEQFhAtkJB/ZYJEuTCggGEe6ia4QS
yH1FH6W0K3SNW4EZz6w/KADveZ8LHOIJgtuhecMuz4Aay91hglHH3XGdMNKDMA12
CgGt+0+c6i+nm1AeoZLqQaGx/VWBbDG/hjuwpRUSlIxEykvGYQqeiC7jyvVNMaIi
+NaH+pRJxNTMJIJszbN9WM75H9QdLv/gr4WadFOu+EB0JktwQHo2DE4RObE9ZJFV
SDCkTBlaf1SXZNvzMU8eIFNgRzSXTTR0Cpdkq59lbSui85ZyOO8/S1QekRcakw/m
ELRHHBX6lOfn0aK00HivAVCimW966oq1d4vTrj4GLaYIMzi8QtyrgvmN6p2SJSJA
05WRYmQeJp00rKDsm5XUpx3wuELhu7cuE9FqgMAhLTfd797ubP7YVN3sraPNxbxS
solM/E+GJecosMS8eiJzeMLZl+Sf8dkc5enUtsJC/d9KEfRPoAf2y1wIipbF5Ph8
xaf/oTnwuy9120dyJgBh+mfDEqZj2tRKJUkxTWeWE9uvPpn5nU3YBpqXAX1yPPbr
5SbR3WR4iJvQqBewZHPlhtjg45rCbeSMu8IR5p7YV2Ihv7ekxQrq+QWAfR5CvRiT
ZyN7ycYpp7okvnC2UdcYLXIwo9ogBOUIWO6duP/44mIoCjidjlrotbxJ43BCuQ6L
oWqfrXT1No4GLqE7Mjj+NmKmJRZrm7DyG8NfV2RtfcYe8EODE8gqNtzoe84lBmj0
SyHPUzNBJBoeE1Po+guFZiFy6SPEWT6lQfZv5AFWPl+nQZ2uJc6NMrnYlAzGjwQv
yVALg1uWz3aTLipy3321fpNNANLD6NOv45smJ7WrRloJuM0AouhxDoKXw4LLNR0Z
p3GrRh1IevwvIOOplVgb1kdj7E49Ea6S8mYeurFL9TGDBCLTULb+9+ZaEu2SF3z1
7NvFRKdJpy0JkDmI4f227044qHQSG8wad6rrbzo/ulkoaHaiRff8rWb3hqafSWu1
DIPnkWaVAt11sDDX7J7pBxufgubmdnLGgA7Cxi+BIBBLK8wzBFDaNlY8XBDgOwYt
WEdphas+F+Q0ExLOQ1LtCOgyrHv3zrnU5M+dQspPd5icu93cvr6C2ybaYlojzv4s
w1NgXKf17rkW3itj5A6mSklDA4TwUbsTCb2Wkxk+L8WH8FBjtsd65Eb6CocHh4mN
Y6cMuAW23Q9wlcMyYraiUB2I8UWa1kPyFaGf+tTUzFYrt2vyuxno5SNy3H03Sdx7
ubpOHbRVGkRy7FgKuEx2XUCdEpJMkfEMzVSR5sKWBp8IhW50GqJ7YeGaTKTqedmz
Evz70AvFS/yeeEvtk+hBAiZ833vwUVWFp11/Qs8+3b4BYZhuTce+fQ697gZ0h8On
Gcxj04LxXWESceB7z0MzLbuPhiB8AzrRjfFtKXUXvN+P99anyr92vG0vHcnOlwb3
5CWEWAf/qvbbY+ZeFGQ1hJd79uThR75G0GJtrSm9VmjrBaWSBJKyuNzQ4S5CbVLL
0JD2Lr0cstNGyzLjsBwGGKm2jvtV0LsPNm25lg76ToqdOAbidb+avK3IfyaPc+YY
49H4ojdu2SkEObpqriviWdnY/KHLjoLQToSIpjDHzGpCzHuxNi+F8A0qp1xwK5jC
RTIaX0KEea2lE1Ddlx0dZVrKOTZP6eywK7q2ZhdtGlugR6PUvIgcCyjc+RO8S1q2
nOw9VmV/5yfBEryxBppasbPgGYnuIU7tNh+uQxfejmhLf4g9w+qo2RaBzb5EDuJv
2XFcNN+UUi9PqB4o3m7n3auZV+I10PTLslk9EMWTCGjsgwTzujEeGZohBugRMiFR
WK4YtuBnIIGqBgEKxkcmLyuQceu/7xDu6s7O6RAczzTfc8uniyXCXzYYkSb62IOa
vE8ZSNrqByp7uQByG9IMsd7vTWKPJOGcNrLrqgxfvWtQVV4A6q/E+setYDaay89o
5fPtgOPYlOhAkUOcCmw7vyRP3VW2sGIQusYkZDe1m7OlKXey8uUd6tLSLxvBU4J2
SJCcxY9DwGQjg6+i/wj3k1OrsgVA4CowJcDbJI9Nam9w9YjwIfixZ1Dgq17php+F
YXc/9a2nJIaqx1la0KOw0Ln8P8L39uncOj85SU/sRi9P71Cg0f2wIjv9/TAkKzkK
tmA4Evs08d7On3i3JInI9uQYoH3bmhnj1Nr7j7evM3XxIgJdm3lIYI37zEptUpI6
giC711yy7W99pukKNKRskmgUqJu4gxkRzpL9n6utOjmThyqX5XcuftPsP/DSF8Th
irXclFWr/UEwgb44LU9Q9upjpRX4pBX3UanIs5+4cDHfdkW2VQBTo6s1ZVlpUvtO
161zE8DfJHDTZWtCcCseOZ0GjqlvUUlm+Ja/cT2g6zdNggQbUQxaeR+8/qhbEPZL
SWuyCBvhEd8MSJ6Io0dau+oxcrSOr6KJw+jBarSaY32ZK75y5/NKfMoFP4++UfOO
qjVGQfZNBC9oV0yE6b/3gz818WJ6Ly5fUyrb8dqfIPjpJd4gbQQmBS4hU2/XjdwS
HVZQQXLZsLOigewU6xyRFSoVgVKClVOJkkFM8yOVZJn55S2iFCNiGMIK0RC+fYMo
rigTyekbqBX+dfn2RYOh1gJN1Ox5XW5h3LzPhiRaFaNpa7D0/ZU9+wUjXEr9I+rI
dyFKXEzr0UQELdhh5qDuOgHGlUfVnVsBjuW1MDCjMwrFy5SIaE0ZNW0zM9ATcxlN
QPUjFX/wAl0vUueyD0Yp2sjn+MsoeBvIeTGUQRizOy1jB1oSN4l7C5G8lSe7047J
M7L1DgnGO98mIcvwYiH1x32+6xJ6egk96XxmZowkSXPdD5sY+P4DUUhLe9SRvl/I
WksFQOEVTOqsLpuiDmW19+g+ypj+S1pMaToApHVCzXajshepO19Og4mcg7gGiZbe
obQZy7YFVQmOQh1u51elxeenY5ojZPCwgVzBUQbP+yls1LwZPhEfBCqIyksjj7Gc
pl/9mXIZTIKufP4Ni8ExmXDgs0Rg+oXqLec85/5bpKsQjxCGpPE8YRkiPOAk19GP
Kv9iJIOO/2QpvwWBEhZ0zQO5KhQVGKp628s+WLRn/UqH463tS0j5eienBjNmifBa
TDAbpVdxyP5TR0B2PDjNw/YNdZRQeoMR41xh21YO2EeIK+QNE+bS3JPIaw/MxMH7
aKmJZSgJm5/uvwVvl/f+eTZeIexjeue+7xnkg1FwY6uHvF9PletVUiwahtwH2NO1
u8gp0FVeFDwp0/av15BAPE3qW7Kb0EA/Ps+xvjIyQFE6jTnUp9ZJJx9A0dMd/3OD
jy+pL7N1a8rTwtZXProUWbDNJjx6USY22/PpbaE5wMbUgdfBuoaCiDgV5uvItnTp
w9nmk0vnqd8B/TssoJGB7141adKRh7Yfm/CpHq9XMBT+dq8WZJJ+s46YKoOHhPKz
ggFhitQg22lKDKUVuWAphyFREE58mgwzDTPXPUY2UH4oi2Xzb7J2clUtEEoylKjP
hsYCicQWhyZZ+YOgUJy7/c53PAn9tPSvCFeCxs8C9PdeU5jL41RvKtCtaVreUm86
5E251kSQbac380fCPXshXhbjUCcIDF7VUiVqq88VV9PFNlwK0oaSYfdJDS1n3as4
ZTIwAervzfx9JOFJuP3ovoZke69H9r8rb74flhl1U7DC3MsfCpdF0qhL39tHmuHV
BSUAjeb7QKYhEslYHvLpml3tfyx9WID6MOM8yUD7uMEA2it22sbtoHAJW5Ftfyqj
EWwjovqYIhOvLgLFEMbHtog1bUjtz/ypio3NQfQFvnxUdmE2Op8NhR4RRVMNJ4Co
zjDxQx9McsbQW9Jq2MKWQn3mE4hf/uQiN9KOEhvlqvT9SmqBiUh76Ti/34CApvrk
uoguCf27shIHf4XcWqNNiWQQh1PKEW48KnQj1UO24evI9UcLeFJNNAD6C6etsrLz
J2vZSy5Y8KlaVRZ6jz1Zwfv42Bcf/TBgNu2EAdrnrom2xJvRmpg5CAOm2jSk0+WI
1JLTvp9jiYleJ0BA1d/Di8n7ZvRMf1aDRvQ1g6TeeQpo1pn66ci2lIhrqxjW4aih
MqQXVq8KFNde6v5dERLewVEzBEBwlPX/be2/3C8GSlE1azcI32385f2MnzXpqEX3
KI/ClxJsaV20fTVFuwBACHhjNQ7UzBK61x1OU7ZbYnFSYbkDWYqSsK8ciCMp96I3
EwI1rZ5I8JvOe94WLG7h/bTqHw95OxyMpDe50qj/HKL3mtIlnNoB6/bd91KW8Ytx
pvU40spwAsAgfVgLmasRdqArArXUW6Of4+u+Umf5uV4rxU7orhn06fWV3re8MS/t
SO7uIgbofccLBvBaEKD4V8nXkxCNFOznKTfy16GAWSS0PTwPHif1zF2lBBvDBdbK
XPk5nc7Gp34HMLoy7mXKIE0Y7QiPC14gS6nU/MD6CkKoBg8qo8G/6o/NZh/FcNoL
Cw8Eyyw8NXWEBrm7Adw2EYg5rMY6N1sMoW74VLWrtFNRuS/l53g4SGOoI31gbjSj
GFgqUAu/5rq3xPdgnqGLRsfjcpYENBBKIAkxmskyYDOmwctvEa/Ib5a/Xl4C7A/4
/qMaf5iWp43FdiPrUapz3uehZ6ecS+2g50lW0woMfDgLFMb4Vtv82gAf1x3ftEhB
oQP6AyAG6t8tRmmSO57J2twRHdOUOyjs8TXcWOmNWqwsMfAmfLtB1m/u+EOgOnoB
Ll8AbZosUFl8yaQuHBdX5RP/dgCgj/X5/jHPxwgmf6sTO/tvPmiqJo28xzgx8Mdh
7unI7hA7XE81RQIA6nUyYKZfOzWENjDF0JOjo0lelIWNOECHWkSw19dGfrJCvVCr
w9tUfu6IOqmq5FfuKpIxXMMjLWGJ1/R2as6gwdn39tJB9OZWvhWqvAzsNqnFPgSJ
bX4oNQeOhO0sxOLFvPh84WAM+UkpiXLsVrbCbvvsJ/s/VzzHjhrK5WQ78xSaxhKP
O5g2de7J3S2fH+J839HnYO2clGFHarUBJS1O7VPNaBAAv56b71t1kU+qHmmwNAWI
S2GYC56m233WCr6vso5WPUe+XOXkDtbwKv3Vidob57mY8DUnRmcV12xcTQaTg5v0
eLworq2gNSYQlmOFm1jOrDixmprGA4flTdEO4cv8k0iyMofR6Cq1rwL6a9E7MWe+
1A2lzNPbOlrU1j54OO2HWczljjc/hd2+A9r4YCgyi8sXx4FDHjV9BQmoh+B4t3Z3
cIRBy9jk150J1PqhA81puza3pPI69VEOkxhiGESdKNxjJI84pnd8xYQoWRNYjH4R
WEWlBpuaz9p3+lK1St+4K96QdDP2kesC6Iaup6NjuiGp4pkbpjlzYfJmPj0azzvJ
8qyRnnMXTZpUEI5IjME8e4rutXsgTMgG41VquQT6XhfucbQ0DqyWI0M1sc48+n5P
Lsr1U7mSi49RYXPy4Pcmj/a04m00E3tjxilJp4ICRU7Oz1uFLkVvByvWDusc/5Ro
Br8SrsKQkYhnip+DOKeDexulFOpgd8a8Wi6FfKaOXfZHtUJR2Leu2d7dqWbM6o11
I6IaHAof+PSKn9A111c3nHIpS/4Zt4mRwETt4Nw9j64hdcXxO9weN+ycGlu5gvsr
buAw/MhyOcGJpc34H4nh2K+rZAlNdlKdzz1BQN/P31yXz7jpHBBDAqpRfXpvbGjf
IP3//L6mdE/S9V2fk9UM9GSPqWVJAxAWftgqetX/cTvscbqXalwqu1/Ei7R7V57t
a/pcpVlgoTfkc9vHmO2VfhnuN0T1IS8VZNg8qthC5QlAo784HgG1Gh1f0CvVW4ST
FxHJpDp6rdkNN8ItiAszFeWnCAZ/TVJMDDVJeBK1CbgeypJ/aEQG2WAKwHrS41j9
gN54atIERFeyejIpGwgILBmIOFPcZNyQbZPsFgQ8fgiJpw4UgfscU3LvpUQ/RV8j
HMOYBsOjfjlhjTGE4myfQlMpXVlQSyNsEysq8P33WynShS43PKfbZFQqg0aatUkC
bY9WU5eGZbDaQ7Q7HZ6mtwcl5giut/Va4FzfDXdHtD/SrSpXe8knjzgCpp7ZuwOL
McmsYzEq5RbjwxzoDIJoQKS71r0ja56qKnj9ylS6UaVKDl1Yq++XQfNKmzn/AkM/
C0q8ydQAzkPd6MjcfbEB1B6yTuRALgk29NG+Y2Wim5uamvzXHD1UkBwQtPhQvdkx
1Wa6v5RRp1wqYPl7q2BxVrCOEOYaXPcoI7F4trtHTwrHg4KDQT5STy0x8qvOoWoq
gzo+YJhc9b87FiecoDEJBjKZR6YJIRDLhvJ4trzOWHGqszx2OZDTMofgz3DFAUZe
uXnv2NRDChuk2/sjxuMsg7UflCY4AfwgSYDJiL5JWlGiaDW06CEvDa1pTAFpNA0t
INO3YVzGaE85neAZuxNF9p2HwtsnU/HSFsYdlOJMfYqlcKyeE7T/hqEa9hBHwQ58
8642sl4CZB4PjFzGmXDCrDhCDT5p9r6wfPK7NckiwzPXYkFlbuurNZFtj9MJx3wm
6fpK5T3LxRp0kwx1PJ52Mt6lnD7X3n2cHrMT+vtCoc0X5E2PtrN4BrvzdBJLSDXx
DFxB6aXzjSW1LJPi1eYx62bYklXGfoamLnGom4mRedEHdlDjJR8HdvgFfn7ROmPP
y/RvbOY6zW/ZhYPw/ebj5DS2Ztn6cEI8JPYJWN5bDRHN7lflm7dzckJzKX8sWNCM
5jMtfkoeSJFzaPxUkrLsF17jcV40OV0jb94Va6xtb5DKVqQ9cVo6xLXi3PFaQ1rC
kYJ8vI9/PFcRgB8/PGzGuFnPOYpSx8pkgAqZ+iK92GJx3RYvIDZlvIFJ4FXz6r85
4eJcr1HN9MpLBjK3vlZJLK2oKROW/r+JSf34b+UlyRzdPtw+F1kRbW8qmPt5mn0n
y+27TWxiqmoZCvLkh8tqmez2Z63utSdfjdJ2DGuDUEbdLk8xFRMjc6Lv5oXiNqXu
stKaRC2sOI/xDJ+NeBDfuZIwsj+Q255oGiDHlE4GTCMnn+OGhkqmwiSa7xYCcT7R
mtuaQAy+Wlj9jkINBb4qIrykDtjJkWIh3FMPq06q/nNII8e5znxSznSuo7FTa1GO
e3780xULC1dt9VBE0GUFtAPASPUws1dn28jvBz/W2x9N5DLzKv0Nnr10O9Z7p+I7
ypFCJceXUcjHuCGV3WbIY1ICTEIyDXfXwsUmmXxG75F+lFL8ryuwg9nLesLATe7P
1fdBGC1zsLzp4xtdNDmMI5SgpYryuXoId2mK/OcahxBOU0TwZR8BUSFAEBWCqK/t
ZnakKtJC2FEbSpT1jn5OhjvDuHbk6mdCc8XWIMcIwztbm9GQgmqEIrZVecsqH6Gn
N78jJiD7NUaKVODwJiPxVj5CwWk59K2k8sRrVBtJ/2Q=
`pragma protect end_protected
