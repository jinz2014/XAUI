// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TvGnjB12cQDjcIw8p/inpu63LKrZS53GgMLOCYLjVb5j5ua3+C0OwYtA24cyC8X6
uyR/zQfn/Jgol9vXu7Y8ACKFV760OoLdPglQE6PZoPFHe3vhfDUsY2fiVS/A/1Or
m6jL36oc8I2ESoXXF0SbEfjaXl9TVJjA6UTkK2k/aSI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6080)
JJqdeayEYkWPZnAdiT89OB0LVnX766e6MQB8MljxH00e5/1rsVEH15lDcJlUdj3L
p9G7YlruvX11BeVGwIvpdxxzWrYLHDR0m3498795qHS024FH5QuGsuJMIBbT/P+m
WqR58Ie9mAUi3w5FFYi8p0GxRbehEWemGsVN8rWcSQWI5Tm5V7voz6bwjTTlUh8p
okrZpbjIq3etEpQDMoJR8Es3LY+t4JulPtY0Z+cnrCMGVvhqKL4MvGz9SC1dDgAj
Y+gjrned+i2JsNdKT35FsoJZNitWhC0vz5f2FyXvbL/qc2Sviybw+BiWqm1TvQ8T
6y1WbxdHUzxnJLhc2X3ID/JBDryzuFz+Mx90a1Q2RGlNiYNXvbBDwNRxjYBQwmuW
vnc9bdtjW+VTm/zFEp3q3ysEHIGzNY5oNrIuAqRKBJa5eF+HNwiFc+O1/CkB6eQu
l6z876QR3JFCQqhmYfA+tKZFyXMYIBRyzYaP/uP5hlN98H+aD8DBjn/IUZeBq/3C
I+YLStxkBmRWQ1b2SDLY24gdr+HMBJ6zSK/DZipTdEaYYoeIw7cd12KZ+Z18F1VA
IGiaNKNfDQdgjHIvNHkagnSFEH2a2xH+YNe+ar8COj252Jd6Y47glLCVEd1gYuex
8CU8hzlX+Os+O5jJ8m4YNagUg0tm8ero4OaR35uL+MFr5UmGAaGUHM+kRdaDc99u
jzisONIlwZDikfbD75BvH6Ie6+vYfiI5B3FxU4M0tuyzbmJThtRJwN8X0SIjaMrt
uoIUuiU/yrNz7CENroAXRhxmKigFFILNTJdF3YGS2NTz+HgpBMCiPKcLhbHiPyQb
Y+9ueEQEEsaDDKrcWvvz7EWLxltVH21BQvJaUa/inMEZ6aVJDnc7NL0Us+jcp8Ie
MQ9Mk4WUeGk/y0YKfo59jJ6leULb7dQnUisDcHoson2VPavxi9JCeMhBDV2LK5TR
cleBrseDwq2d358Z7zo9PEHMAuMTpoKhTvQCb0oIVt2PDqwOZ1cnMqnu1eRYwVfv
wOs592ygpiTPTknhIx/1qAbv4Sr6u1/2SNf7defZZ8EvtdtGiwEqJ3Jwsy16HOF8
DKOEX77xVCSTSKxMEIvkLhViIFsgvY+ptgJrvWIficZoarHWhYq7pi3YffMalZUV
p48b1nhYsXLfqXQSXwAn2zWt4/WJP2md77Fc9i/+EtH17fzrf0OoNPd1fkNJeKyD
OPH4JsTRYG5uSgkd0pV/mZixTs7cOdH86X2SItkwtt9gvcrLeQiRm4MSPjMeWh4C
pYi31lr5+OeTuYndgWxBaKnW/Wf1Fmn8oytrQfXq62nGM6SdZflkVjledMqKzS9T
A/oGVYjR1JVLwhr8kmxCn7dL5/KHGGTjS7bmbDqkfv5/zV2hDh/izGcVl2FxnrVN
iUvr53/L9JLomltpakEeGyNbvhdM9aiIQYP+CGRH3XgKXSXtNdILf3I6fUQRBS9e
XvCCBwJFHVN6dtp64rTK4Z5mogdr1KVWTvVk1wbvvI0Bz9IH2suDi1CDRMmoK7WD
4/W5NktXnPuZNBB0uWXdqDGzf/zfG1CD4P56x7zP8YUCBhy7ZE3Mqi9xk/ARwPo1
2jheo541Nh0nAk0Szga0y83VLbHsEOOy/2woox2CPWP0QGvv7cgYLh93hTT4C3Y4
w2KvMv4UbKW/Z6aHg22YwvYx5efbcxS6w5hKbJbat1a7Zw1vYOegytdr4PAVIWwk
/ZUZHfEpW/IOr0mZFoAjqBH2d9dDIaTDm21r1H/Tq77gvHFtbXLKSKSDq63Ar4ok
/lodQQ+2bYE02lswRdaZKlW00vrxSRocLw8Z0snGdJnr9NYQio8or55ALP/u8uHi
HmriOHj4qYVnhtkK8odeHq4p4itfDCNY9svCsNBu04JjME/JCosMVF4jNmITMGrA
IE7HR+xjvrjyxekdTbCR/sq24B6seI++VCJaMsaRssp5eSJuvXlY+rBbJwzOlL7w
KqomCbOTDLxgJpYEiRnk8+IEYBWh+nf9csVvYd8rsgkz5qb91sgUFey5U62VxN2S
ijBs3H+Vf+kI6Rm3WQ/mxuacY9REle6YWTw/RS3kifvrEds3XvOsyX4BrrncCXqw
SETqB5vzpnUsYIA4MiI7vXDtlcV0X/W7c81R7w7xp2SjV7St8jRSMoCNwXHSLymc
vizi3Uml0H3HqGk/42r0mF+4lSr3hLu+4TArG85nfAhci+rpThjuRkgGen18ESw8
ZAN0uzu4n+KOU1YIDkkmEll/9JF1ozMbN1W55xaB2hGN5fitKezRMrO0FpnihGy0
0OYWJzkpb/Td1oHjWkCB2fCTywCd5C+4s+uTLGWeRXkUxCwEkmTdBlelewV5LPkz
Luol2d4sbdgd1sPitYdM4tOAV1wRx4E9iaSioIO9r9ohQRgC+tVfJ0zFAGP1iTUs
0sU3bemK0csfQbcWPQnKBv7CBeMQgedSUKFAkoeQHYECxqSPdqTRoKyWcId70N4S
0jAJvVthWLD8LWGKGZ4Vnq73Dcyenl4BO9YUVIwtrv1QftGBHuhAqTbRsJCzXPES
XbjTTjMW/HOHVRw0hJgJvyMH2T87PUDs7ZkrFX/xZM1MKV93U0dOTE8F5TPDHPWH
AQK9bj4Y1nE7OJanYPOsYsRuJr/b374ASIRklN4VNFjnvs+mCzrXmG/hLcd/4DLK
Lo5YiQfnkCnU5kN7sjHnp4fhHOKedG7KUiRoO1wxDjqO4NJf4JO9JemswHDNdnkE
B18wIH4giT1peAxCHBSTx0+QscBxLjIaqhHbcXJOesaTG0mr9B6vJX4yUw+Zmatq
Iz/KK4CKrzJzsEsUispSd+MPd2FSQT6/DYXFV5r/1CivdfkzuePSqJi0CrUYuG31
dS62y4h6kCp1JHE2qDqSLtPyg1deN0e3nHVe0FmyMH9kEpnTypvTqSgyah1w9Ucu
8+98+/6+AJ4E3AlsBPLWGJm7YMTQG5tk2r1b4kPzFgpXVTnyQRh+4UbFE1s9Y7SA
6p1HKunVmDGB5PvPLbPSrwax2rGzpSf6463NfP0NM4C+WpA5EiQIcg3PE9M1MaGq
TLrq3BpLEZqWqwOZ+h1Ds/VX5H/ODwDJvsVxsNI11JQ0n1SLjlPfu3x8qPHDDe3e
M1N34EVJTeoXNfFmFTmbwvRt6Jq7FxqO0GnMl6K8YruqfUjoeVPiyIA5dZVuw/cR
oo3EYXg2O7kcsjsy+E44yF8cp3OSGCC+QdLb/nIbqq4lUo2AnpGxUZJE3ZDLst/x
g7IS4aEvae5iGBh24viUoT0a3sq2wDtt3x3MwJ4AiXDFP6ZX1jD4Qq16xKg9DMzm
YwrqMBMANcALtMLe0rVjxQKod/uS7VKKb7xZrE9FN5sO0S72pPJHtLrPoSSOwkLX
FYioJXnzViV86Pl+KdCLpvyP+eNjPE4oXYmD71AfLM4tZMAFAvQWoLERU55lMoz9
8czVZ88URz8FK7VNcpfYHyq7S2J395kMKSYKjNi/frQD6proBnJddmgjWZCOB6Wa
ZNUfEgfaQ+XSa/Wt/4Yf5os28VEWpuE7ZVL62+AnrI2950DkWUev/AdmsbR2hGTp
MpEeBqJCgEdK5KhYGW8LQCWoUk39fTKcOhfmkl+EjYhPH7rXASKf2W38+dP2wt12
S3JBJussX4hF5xEZGy7UJQJhwzGecxGauHeZJ84hzb4XtKqa4xkNbZr3CcdTRw+g
okwxc1vloPfmjgVnEvU4B9hEo8QpRTC3PqMNOKq1ZteKgnRNGIyJljyNkCGF+mB+
PXCTomClV/OTxSTGc8oSKEaMPNMAPi3RDOgdq1NQlmsegmOsGYkrHQIC88jPjurd
YQj65BttlsNROVos0Px21n+1bY/bGfw3SLu6vpimlY0qis8N7Y+5ujnG6SEBTZnN
iGHcwJKSVZR3oQewKz5G7UQRxzEPgslE8qNvUzX83fuaWEGMQ0HBFSQJNYgdX66k
hDQHC9sv0jSXIaV4P6Myn35nlBe6InYYHx+GO6MCSIj/SgP9FnnMEYs5MV6SRVF5
l95n0yPrXeCklS7jhl+g2ahZa4GmbEDIXzAkP1HxPc5Y6sx6myfwbPkkh6ZVnabp
WZEJ/7i1zIrramDcVlOq4+HJd8EsJ7nWAPnPbvjN+AZtNpwRz4PCg+7PhOqfvkrQ
Y7Gq4EZPChsAE+dLrEZGav1dGPgV/BcylOHkf8q5jFL7qtcakE5lLHxovkxXgwrN
1NMdiw/w3oZXEzuVPnrRXiSHaz4z0rUTvElCX44b5W4ORaXZIgW2hiHhrPpn9rbo
tT2Tnj557kSPaMY/ud7XAVSK028dHFqd/NSptHNtDbAnW4M0sHjypMmDVhMD1Zz2
12DdMLWQseem9SvOSv323RQPJZIAIy0QeGRKw+IUKUKNewffiNie+zK25R4zzcjl
kfbELlfMwHVpeFN6I0cbPVlTVnD4JRwkKyTvKlJDuyHluKJQuiTX6Xf6lBh/2fZF
iG6pVdOU0KAkzc5JGo8u01ci0s70NnC/vI+yHeMBL0fVliv0BG6yS3kyQnfe2Gfd
EwQ6PDM7V+jTqwIOdWFZ1ayG/osKmds+Un7WTyWJPTYP5VYC7D7YQqDkP9XDy4R5
d3PzD9eYnHNsPN3Z+6SO+lea0E2WsDQ5sYkuAHrL/lQw1g0ImEedKgM8cOcRMwtp
hM466H46njSiAf/V9f550iHPc+mI41aZdShMzjUSg3AQHj9G/plricqjxBPiLpZE
K3dm5CYIIKu0agLBwXB5hEhN+RBR7jqbn//D/Ykb1GoSaAnV11KCd9auJXj0+Wyj
nHbmOiOkAw3xINrK2sGV5hRWBKQiV7WfDiQC1iot14pAk57fgHNWV/dASwGvrvk2
fawwu0C+7czPHWw0oe88bCa4ZBHYKkkgoTp4UmHBNqmMx84xEei3Uv2PJa9M2j3h
mHji1ZXP5iyIRV9WG4hmxKliKGvyAcmb5zyE1SPKgfhiGNx6lgqM60G2VnW1Ants
fep9pZbZsWxe+0vGgHZwJuw7Y96fCkcofTOhDBWjB4WFPLv9VtBRe+keBvjUH/OT
X1P3Um4k+Zlf9qDztWu9rIQkMRYnYTl7Do55ZresJmguWfOl14p35ucaf4n0ad+4
dqSK79eC9HwZe3yHIzWoB6kmptQm5vSpiOceYPpBJ1xdA9+XIuSCRC5szsyGTWgY
DbprmlP0dEztC06zuBjFfim/9vt9iJ7Gt1U6/W5FsRJlp0flvAj5aDUo1gx3Ydpk
bi/Tow5epS+dZAqZLta37ILf7HUa3VDDcxu+STmgGnkzJTdq7UBxpVSnZ5K1XzSg
xgV1ygwzXerlFMdW3M6SBNImHEcNgvkkbOBsBaP3aPE8uA34R+wNSG18Lax89tdH
zkcyE49n/nZkKUKUn12MMa+G0QPfh6NgetHv6nFA5tOg/l2GyanffVMUqcRbfzUm
6Q/1swn/Kcb2QYRuxQQbVsDYxyHJRxw8xI7ONxQI1kpwwAMKFt/BMLigTG7zjAkE
DoyB0qBMaBG7WkToRR8QeRSa32YwGXQfhK6YkIYXL0gDJ1s+Sl1CB5mw1bzfHNS1
AT92rwyJMcHBV3BwbHcCaID7Gbo3Z4fODsA7hXqo6g4LQEysTGxVqCNrQ7N30pX6
ELh/eBwrerLPBuG07/JSWYd7MVzTxQKqFAeb0yLYqu+C/KJhxHf9DWXxSJSsJH0c
2Z4zJHiEIdMZahQagVlWI0t4XeBxVgD31kVX0JaLEtcilXBupXsBAQ7DLgchneoP
HTYWLiI6MSuo2bHqIWnLOBGE8Cxsz5BhJYpQj595tQQYEhQJj0qZvIGKL9Nx+XMQ
+cfi4bglhwbFr0hmheC2HfM4+0hQTHPcyg9PSdxg+8XcquSfV5pztz8FqdTbDj7d
+do1pXk4UlmuHOufVJlnayZsTp/h/t6LeMC20Os+6lmcUuhLwWUFfEwJGqz8RWF2
OlSToOPuicK0daTcilzdRrieUQS+S8JGZjPEqewQ6w7bHircaLeIjLlsVLgG8dOr
vvbZXBw/mFT4/0sxDDnBMPZzB1IkCVjzV10tVz1JkBf6+WNS/eTl3REcOJJ3/no3
0v249q4pNp2H8kIdknOnuFYIj3fld3Lfic/bdX5pEovxwt7+z1k0OfWoDPzloZvk
nhpS/6tJMt4WjN9KO3S5mWnArtSB9IyAAAG8OJRmy/EiBXJEo9+u5SkDugGJQsnz
8IqB621++s0YnFr5Gj3gnrtOOauIHSMAmPDFi1CjvIUi5AQpt+5bH2llPmba6UpW
oKviAgzr+DQ5V88WCNzfTCBTDDUmzqWqfWYGY6BSOVSNPGpx6AnkoU0fnKwFJi8/
nPe+57A9x7CFOoPrzzHv0d4lrA2NRTcklW5/CWZ5pg0/sy8rRC+xV3r/hqXgivNF
9mOT+zdUqeCcjxisVjn9cqXQqpZ1oC2icucf09Q+JXbmn4HfNFb8Eg9Puj2gm25B
2qPOAkAOWi8tSl7y2/WU2qhpNU5xYn/oDPzFRjhjqVGCWgpALPhyo8t4i6V5Je7R
znpeQDI/MpGH+plECVxKSNKAEvZmyEcffA2QzCcXHMJ1UZKcHRu6qiIBWOTNddZr
YSRh9QehOvbUORP7DzSwbrVaJJscAEFAGzBRZfbkcTpROZbFiTMtOFZgm32Ychz/
rkuxYWCkJiuTRfvY+CK0zbaUH9zuyPFUqv9FLDnjaxmrPiyHDjOAck41cVG6+mMY
37fFYmIRfXYCK2DcEZk8VqTTBTS0RRVXaIYmlCIN5yEoeohPpFv6SP+Zu2+tiM+r
7FIvIDDe0n/I80yEuMJF6dQqaY4R7eHa5i9jlLEUzbJimKbNZia4ERcHC3D3TkhD
wZCpq0ev3QFYfzdRaFFjIo2rLZWLveEcRZ4tBe2NygPWy9r0KuJj8UgRiJC84pcJ
kNIDi/QfxKOvzU07dU8TKOJCOWbD0TYclWfOGxwl+T9nU/COhgqxEVeMWiRyi8SK
MjyoK14axQoNnXKjLSxcqW/dC4Rj2/ogIRwKDtKmZHj1XBFNaNc2NVt+lolD5OAn
uzLBOR2JxnwusWPH7uLJ0b9WjNNRFqa6mT7PsTwQpTwp1mzOjhCd/Sqh1zNV1AsK
GQ7hXdZC3ilHLwDLdsg3UZrFSLLHgmq021oLC3wWXV28SDKJK/UiBJmvAWXbVTOY
vP+4VXPQ6wXA05SRGVwOO/xq9SaryOB/BTQDgXiOoKsXRFK+0vJg3Dq6b/7rgNw4
/dNi+9uzVIJlSvkDY6yvr/OTP/Q/ZaOsAJHoeXTGdgY9iTnzvjqV8Qc73aCTDZd5
NFjc8aZtQc5yfEcn6JoyQKE4n5PaPwZLNPLlBET8Z63tY+NRUsDSZgy7Askh6cnp
1NmBm6gkoTRAdDpm3eDejp0degjkNVlU5NUiz9wQRrlyOcBe0D7vxUs6SVsfGiZ2
xqvhcGWXRamCJoyhtl1TlcI2GyI5xj0TqU3x6iW2ApKJYOBYTboZo2c9DZ8pZYz6
FHQYCbhV8QePJgwr+0sTsO28yk8RY4Ud6hNn3+aVfL+5PbD51Iegbtt88NM74CDp
fsmz+qew8VF9rp++a9PEKI3EsVfaFoi9TRuEe/QvA8S0Dz9sCP1SxRIrqpauneIH
ssRppvWahwXklKSaxkV0K+5RcL37fodg2xerTCcpVtPhLDr9eRkrlL82yGCx7yBg
+1/xWzqdyJ9twpxnX0Te7f+Knud49D9A6c1tBHqTRoY8C9hQQHnpnbD122j/L800
yy6q2kFGKMSZEI5gDMk604YiKGfB/Q+jgu9Gvfrrf7eP8g92SC8R1f3eiYRS94Ox
tOcrg8s20/woRp52KnX9aF/RUdg4L8Psz9tBGsLtsq0WO82Tm75JpBjWNKU5+UnJ
xkBSruj3Vui/0xkdcRgrXTA3X90IwyptzoZj+zP4aT1CYUV9xQLKWAl6/G3p6N2u
U3JWvIMhXvNwiv9sMDct8q6RQK1FcbCEpu7tvCmUo0Ik2N7AhnLb5+taKGBg0+1t
M1C/XhF4z5Uh7htNc8Jpy5Eg8acgD1V7itYt/DEYwdfjNOkfH1n336cRamiVDrFJ
b2svqpsfvUWEHnNU73mSJ+g7mqorc1NofbNxMtMqO7o=
`pragma protect end_protected
