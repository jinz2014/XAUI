`timescale 1 ps/ 1 ps

// 156M
`define xaui_ref_clk  6400

// 100M
`define system_clk    10000 

//===============================================================
// StratixV device
//
// Latency (based on simulation waveform)
// From the xgmii_txdc to the first valid tx serial bit 
//
//
//
//
// Note
// User cannot drive the XGMII txd/txc I/F or serial rx data 
// right after xgmii_tx_ready or xgmii_rx_ready is asserted.
// The tx_ready and rx_ready status signals are synchronous to 
// the phy_mgmt_clk.
//===============================================================

module xaui_phy_top_tb;

reg          ref_clk; 
reg          sys_clk;         
reg          reset;           
reg          xaui_bit_clk;

wire   [3:0] xaui_tx_serial_dataout; 

wire         xgmii_rx_clk;        // generated by the xaui_phy core, frequency is 156M
wire         xgmii_rx_ready;      // xgmii receive i/f is ready 
wire         xgmii_tx_ready;      // xgmii transmit i/f is ready
wire  [63:0] xgmii_rx_dataout; 
wire  [ 7:0] xgmii_rx_dataoutk;

reg   [63:0] xgmii_tx_datain;
reg   [ 7:0] xgmii_tx_dataink;
reg    [3:0] xaui_rx_serial_datain; 

wire         phy_mgmt_clk;         //  
wire         phy_mgmt_clk_reset;   //  
wire [8:0]   phy_mgmt_address;     // 
wire         phy_mgmt_read;        //
wire [31:0]  phy_mgmt_readdata;    //
wire         phy_mgmt_write;       //
wire [31:0]  phy_mgmt_writedata;   //
wire         phy_mgmt_waitrequest; //

wire [559:0] reconfig_to_xcvr;     // 8 lanes as specified in MegaWizard
wire [367:0] reconfig_from_xcvr;   // 8 lanes 
wire [6:0]   reconfig_mgmt_address;     
wire         reconfig_mgmt_read;      
wire [31:0]  reconfig_mgmt_readdata;     
wire         reconfig_mgmt_waitrequest;  
wire         reconfig_mgmt_write;     
wire [31:0]  reconfig_mgmt_writedata;
wire         reconfig_busy;      


initial 
	begin
		#10;
		reset = 1'b0;
		#(`xaui_ref_clk*10) reset = 1'b1;
		#(`xaui_ref_clk*50) reset = 1'b0;
	end

	initial begin : xgmii_clock
		ref_clk = 1'b0;
    forever
		  #(`xaui_ref_clk/2) ref_clk = ~ref_clk;
	end

	initial begin : phy_mgmt_clock
		sys_clk = 1'b0;
    forever
      #(`system_clk/2) sys_clk <= ~sys_clk;
  end


  initial begin  : xaui_phy_monitor_clock
    xaui_bit_clk = 0;

    // wait until xaui_tx_ready is asserted
    @(posedge xgmii_tx_ready);
    @(posedge xaui_tx_serial_dataout[0]);

    // set the clock to the mid of the tranmit eye
    #160;
    forever
      #320 xaui_bit_clk = ~xaui_bit_clk;
  end

  // initialize frame
  reg [63:0] dc [255:0]; 
  reg [ 7:0] kc [255:0]; 

  initial begin
    dc[0] = 64'h0707070707070707;
    kc[0] = 8'hFF;
    dc[1] = 64'h060504030201FBFB;
    kc[1] = 8'h01;
    dc[2] = 64'h0E0D0C0B0A090807;
    kc[2] = 8'h00;
    dc[3] = 64'h161514131211100F;
    kc[3] = 8'h00;
    dc[4] = 64'h1e1d1c1b1a191817;
    kc[4] = 8'h00;
    dc[5] = 64'h2e2d2c2b2a292827;
    kc[5] = 8'h00;
    dc[6] = 64'h3e3d3c3b3a393837;
    kc[6] = 8'h00;
    dc[7] = 64'h4e4d4c4b4a494847;
    kc[7] = 8'h00;
    dc[8] = 64'h5e5d5c5b5a595857;
    kc[8] = 8'h00;
    dc[9] = 64'h6e6d6c6b6a696867;
    kc[9] = 8'h00;
    dc[10] = 64'h070707070707FD07;
    kc[10] = 8'hFE;
  end


    integer fd1, fd2, fd3, fd4;
  initial begin : interface_logging
    fd1 = $fopen("XGMII_TX_IN.log");
    fd2 = $fopen("XGMII_RX_OUT.log");
    fd3 = $fopen("Serial_TX_OUT.log");
    fd4 = $fopen("Serial_RX_IN.log");
  end

	
// Management interface
assign phy_mgmt_read        = 0;
assign phy_mgmt_write       = 0;
assign phy_mgmt_clk         = sys_clk;
assign phy_mgmt_clk_reset   = reset;

// Reconfig interface
assign reconfig_mgmt_read        = 0;
assign reconfig_mgmt_write       = 0;

//--------------------------------------------
// Altera's XAUI core
//--------------------------------------------

xaui_phy xaui_phy (
  .pll_ref_clk           (ref_clk),  // i
  .xgmii_tx_clk          (ref_clk),  // i
  .xgmii_rx_clk          (xgmii_rx_clk),   // o

  // o
  .xgmii_rx_dc           ({ 
	                          xgmii_rx_dataoutk[7], xgmii_rx_dataout[63:56],
	                          xgmii_rx_dataoutk[6], xgmii_rx_dataout[55:48],  
	                          xgmii_rx_dataoutk[5], xgmii_rx_dataout[47:40],  
	                          xgmii_rx_dataoutk[4], xgmii_rx_dataout[39:32],  
	                          xgmii_rx_dataoutk[3], xgmii_rx_dataout[31:24],  
	                          xgmii_rx_dataoutk[2], xgmii_rx_dataout[23:16],  
	                          xgmii_rx_dataoutk[1], xgmii_rx_dataout[15:8],   
                            xgmii_rx_dataoutk[0], xgmii_rx_dataout[7:0]
                          }),		  

  // i
	.xgmii_tx_dc           ({ 
	                          xgmii_tx_dataink[7], xgmii_tx_datain[63:56],
	                          xgmii_tx_dataink[6], xgmii_tx_datain[55:48],  
	                          xgmii_tx_dataink[5], xgmii_tx_datain[47:40],  
	                          xgmii_tx_dataink[4], xgmii_tx_datain[39:32],  
	                          xgmii_tx_dataink[3], xgmii_tx_datain[31:24],  
	                          xgmii_tx_dataink[2], xgmii_tx_datain[23:16],  
	                          xgmii_tx_dataink[1], xgmii_tx_datain[15:8],   
                            xgmii_tx_dataink[0], xgmii_tx_datain[7:0]
                          }),
  .rx_ready              (xgmii_rx_ready),
  .tx_ready              (xgmii_tx_ready),

  .xaui_rx_serial_data   (xaui_rx_serial_datain), // i
  .xaui_tx_serial_data   (xaui_tx_serial_dataout), // o
  .phy_mgmt_clk          (phy_mgmt_clk),
  .phy_mgmt_clk_reset    (phy_mgmt_clk_reset),
  .phy_mgmt_address      (phy_mgmt_address),
  .phy_mgmt_read         (phy_mgmt_read),
  .phy_mgmt_readdata     (phy_mgmt_readdata),
  .phy_mgmt_write        (phy_mgmt_write),
  .phy_mgmt_writedata    (phy_mgmt_writedata),
  .phy_mgmt_waitrequest  (phy_mgmt_waitrequest),

  .rx_channelaligned        (),
  .rx_syncstatus            (),
  .rx_disperr               (), 
  .rx_errdetect             (),
	.reconfig_from_xcvr       (reconfig_from_xcvr),
	.reconfig_to_xcvr         (reconfig_to_xcvr) 
);

xaui_phy_reconfig xaui_phy_reconfig
(
  .reconfig_busy              (reconfig_busy),             
  .mgmt_clk_clk               (ref_clk),       
  .mgmt_rst_reset             (reset),             
  .reconfig_mgmt_address      (reconfig_mgmt_address),      
  .reconfig_mgmt_read         (reconfig_mgmt_read),
  .reconfig_mgmt_readdata     (reconfig_mgmt_readdata),   
  .reconfig_mgmt_waitrequest  (reconfig_mgmt_waitrequest), 
  .reconfig_mgmt_write        (reconfig_mgmt_write),
  .reconfig_mgmt_writedata    (reconfig_mgmt_writedata), 
  .reconfig_to_xcvr           (reconfig_to_xcvr),   
  .reconfig_from_xcvr         (reconfig_from_xcvr)   
);  
  
initial begin : xgmii_tx_driver
  integer i, j;
  // send idle 
  xgmii_tx_datain  = dc[0];
  xgmii_tx_dataink = kc[0];

  // simulation shows the data cannot be transmitted to the 
  // tx serial output when they're driven right after xgmii_tx_ready
  // is asserted
  @(posedge xgmii_rx_ready);

  for (j = 0; j < 3; j = j + 1) begin
    // send valid data qualified by the control code
    for (i = 1; i <= 10; i = i + 1) begin
      @(negedge ref_clk);
      xgmii_tx_datain  = dc[i];
      xgmii_tx_dataink = kc[i];
    end

    // back to back transmit
    repeat(0) begin
      // send idle
      @(negedge ref_clk);
      xgmii_tx_datain  = dc[0];
      xgmii_tx_dataink = kc[0];
    end
  end

end

`include "phy_driver.v"

initial begin : serial_rx_driver
  integer i, j;

  @(posedge xgmii_tx_ready);

  while (!xgmii_rx_ready)
    rx_stimulus_send_idle;

  // it takes much longer for StratixV XAUI PHY to be ready to
  // accept RX serial input data compared to CycloneIV! 
  // repeat(1000) is not enough, so set a larger number
  repeat(5000) rx_stimulus_send_idle;

  $display($time, "Sending data");
  for (j = 0; j < 3; j = j + 1) begin
    // valid data qualified by the control code
    for (i = 1; i <= 10; i = i + 1) begin
      rx_stimulus_send_column(dc[i][31: 0], kc[i][3:0]);
      rx_stimulus_send_column(dc[i][63:32], kc[i][7:4]);
    end
    // back-to-back transmit
    repeat(0) rx_stimulus_send_idle;
  end

  while (1)
    rx_stimulus_send_idle;
end

//--------------------------------------------------------------
// XGMII TX monitor
//--------------------------------------------------------------
always @ (negedge ref_clk) begin
  if (xgmii_tx_ready && xgmii_tx_dataink != 8'hFF)
    $fdisplay(fd1, "%t [XGMII TX] xgmii txd = %h txc = %h", 
             $time, xgmii_tx_datain, xgmii_tx_dataink);
end

//--------------------------------------------------------------
// XGMII RX monitor
//--------------------------------------------------------------
always @ (negedge xgmii_rx_clk) begin
  if (xgmii_rx_ready && xgmii_rx_dataoutk != 8'hFF)
    $fdisplay(fd2, "%t [XGMII RX] xgmii rxd = %h rxc = %h", 
             $time, xgmii_rx_dataout, xgmii_rx_dataoutk);
end

//--------------------------------------------------------------
// xaui tx serial monitor
//--------------------------------------------------------------

wire [31:0] xaui_tx_pdata;
wire [ 3:0] xaui_tx_is_k;
wire [ 3:0] xaui_tx_recclk;
wire [ 3:0] xaui_rx_recclk;


genvar i;

generate
for (i = 0; i < 4; i=i+1) 
xaui_monitor xaui_mon_tx_lane (
  .xaui_bit_clock        (xaui_bit_clk),
  .xaui_lane_p           (xaui_tx_serial_dataout[i]),
  .xaui_recclk           (xaui_tx_recclk[i]),
  .xaui_tx_pdata         (xaui_tx_pdata[i*8+7:i*8]),
  .xaui_tx_is_k          (xaui_tx_is_k[i])
);
endgenerate

// both clock edge
always @ (xaui_tx_recclk[0]) begin
  if (xgmii_tx_ready && xaui_tx_is_k != 4'hF) 
    $fdisplay(fd3, "%t [Serial TX] xaui_tx_pdata = %h datak = %h", 
             $time, xaui_tx_pdata, xaui_tx_is_k);
end


//--------------------------------------------------------------
// xaui rx serial monitor
//--------------------------------------------------------------
wire [31:0] xaui_rx_pdata;
wire [ 3:0] xaui_rx_is_k;

generate
for (i = 0; i < 4; i=i+1) 
xaui_monitor xaui_mon_rx_lane (
  .xaui_bit_clock        (xaui_bit_clk),
  .xaui_lane_p           (xaui_rx_serial_datain[i]),
  .xaui_recclk           (xaui_rx_recclk[i]),
  .xaui_tx_pdata         (xaui_rx_pdata[i*8+7:i*8]),
  .xaui_tx_is_k          (xaui_rx_is_k[i])
);
endgenerate

// both clock edge
always @ (xaui_rx_recclk[0]) begin
  if (xgmii_rx_ready && xaui_rx_is_k != 4'hF) 
    $fdisplay(fd4, "%t [Serial RX] xaui_rx_pdata = %h datak = %h", 
             $time, xaui_rx_pdata, xaui_rx_is_k);
end


endmodule
