// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:39 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GHRNW6wN1JCuMhGHMgqGplMCsm08ifwVZxIk+Zd3oLXHEvQ6DZoIQ6WWzGy1C19o
Gd7Rfz5bkpVGFaH/oAbTxBaKt/mGwfnKwDPoEz3L+l7BQiDMkTh6k9d6BpdO7i/x
nD1NiUq0V5V6IdxNzeYMmNNUYrgj5q2I2edMm/w0M2M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34608)
+aysxnaHHyy1a6s5P+G7x3zHrMwTwDltxHVpJuW3LZC17KZbKpSALSxT6NldNzLe
b7eilD8H1OsvbpSUFPM4MjfP9h7C0m23OKQGH0NJ2sScKJ9+wDVcWavsbNTrJNpj
v5rfUjVGIvOQxr0iojH9htOkHS7R1K6D3x1o0oY+1KZdjOLXCWR38PVRGYlbDQby
ESMIzw+0g4YxKHSfVnN+wtNq2RfWIjVyPTgXHBNEjYa4zCf5O8wvN5VQ0cZRQA4k
I9yobt1Z3HpsL5oriVQZs/9CuEfPcTXL5/xMfrCU5CU93xf5M2sqO8QGhSIOpqH3
jVDyaG3efNEKxdexW4N+PYvYXBRPyBI0BBKd6lgrIW0axQ2s5cjXtvCBLQI7V5gn
9CGwjUy2JV5MsBPPYXFS5n96hBde6y8gfMRY3q/Z1aTKZDPO6ynPyuzybQS87OEu
OY5zCojQYxR40Y9Gapt5G4ha72cv+zbOXDYzGiGr5yHf2ro15fUvaXaBhui+R8+f
DHbuUItVoQWkI0HBz7FyzmWXhhZt/MEKu9jlwnaQbRifB9yZcD1iRIHTVs89e9OA
D1OcasORAP3uGRjuT7dxDxrxt3gp63FyryRRdD2AbytEKPVVnkjRApKaxW2dSoty
29JW736gMRqkWvuEvwi/NsttiYpFdpHWkMv3e0FPX49jvIbThPH2NuyRRlNci6Ra
z5SOkru76EEIxVlE9/CeHEzsdza/G7KYMJJgfz6EtlE9F06Dxb3+CqtMmf0J29wC
OeZQaNp+oPvpxhajVIa3S0F5xv5u/ZNkHpuLTLbqZkFLuaNsDP2RtEU3bVPv1AHc
Wg+/8OdvmugtgnBjTv6wfGOrIaCmvZo82VPFTeYDoNNFP4HDfrthTrgfA0JZEn+N
gNiGHyPv2WJZv6/IuHZbEq2Ta/l8xsjMJTm7lls5KcqoFs+ip+3lgp8dyzD04WTK
LYYo9dedGDHqwVHg4X6Hp2S8KSoWqtk53MEJfCMgPpZ0fNlmglwQMGNTGmzsFlul
igNO1AT2PIH2ZcIcrw8vXTxTc67fT0peXyxWsWTCcuoomQZ2lwoZ6Zj/aFIVxF4p
XXBwS7qT/oFzpfqEsy84kMXPTWq9PDFgHBj/cqyGZrvneJlw61N3X+UJF9UL+AJ0
DknDh7VmqR/xZVXRgDGCA11mLGD4d15s0HzLm+3V5LDTOTwibB9ru2NNrUsUxYw8
95iem9Xe7STsYIJXSZPk14WeISUPrqmBh5GVud9fN5Kr2Js5JT7df4yplURqxZTR
hCielQNo7PMFvcTGhO/RyOmGqN/NNHRQ3tEH4ZdZptnGnHmFQ5lRGu+twzgr+O6u
PfE7rOMUukDLKOEFUBzijubj6wCaD5eATmPlmg6jhPMtWGkRQN6qy7ItZiUy0aZ5
EwzYQglVkye/aSPjb5jjDfwPyT7T0edoEWPWfzbe2d4iHv9aIzhRdN10Iv17dLPD
0U1VpcuGwIx6dPdgwBtF93nMqEMe6wPS6tQO/35MTfoPJJ+1VFlXmL+qdwdJyr+i
yUP2JOjqyLviyEzPRK2CjOa5ZZGB1lwUqyMER2y+UHeB2r+FeGN1Yt7B4LDe+TJB
TvyYUc49dT69Z0JP7HxcOQ+8vClnH2QvvLYEiMIEEnhbb4tDRfK30eu/NkKmigf/
FepVMaXb5vl4GRRh3XQJ1XFGIdNnipFVe44/zTSM3noab2viGyDNiuyiKTWdf4hL
zQIRQZ6JQV5rUI5paI7tlfIEgNi93LLUKe181eQQ8G6hcp356oYlzhhpsbuAwosO
12Q13fYLhYvEfSU+rifX1bVvQ609VCq2cI5ZqzUdiI8vYu46w4blS1dVSBcxLcr7
t4T2bKehaAoBaHEMEldd7XRHoLO9MrGNnmpcSvKnqVfuOfRJUIf4Q+Llyr7wYlLQ
IU4e3uneuXWhYO3pZhIKqnrNxX5E5zZzWXrIIfULSU58l84OI4kAW9tOay3+im2d
UXyDq7go2PRSSFnXY6y+CLJnDI/0cujHehSM7sqo/102bJlqVdXG4hBDHIWCHY7S
Fxc8RbxluyH1JAMrE7XW/VGvQQF9liUAOg6qZrMZE7nk/BZ+ClJJ1vcO4cj4r0Ot
UOKiqaBRVMpt26JHYU7iCRomCNZT5A6B93oCvrZO+Akfunp88RV1s0RJn9DJa8n5
akUa7HfkFTemUyivQbjEPF4ZUa7jW+5UTeH/aJI9Cb0FO9tkyuS6O3n8DsLP9DZG
1uyHjvKV27tjAzmXwQro+A3eNxCvUIqqsiApes/AAuSRmfCNXW+jCkFhqUD7tdfP
nT1IvLaGcFThxGj2Bue56/9GPwVUSBJiktoRl8cDqkr8xNifqZdxWqyHIfDlzj2H
AbrGLDpglu4Rklcw3qZCPO7roTzePwfoMfE0w6tvju+aQgwd/EKfPgM7a8NeFK5R
caCCrVShWFxMjcZzx18VJE/82aNSY0Nw4vNH1bs+SuTZNVrzNH1JTV4fTr60Rp8v
dIPJ1dmC+r+NC0qRNZ2KT3SDJ/gwqlLqTIl+fU8MZYuuuQM/7FCRQnLX6oro67Fm
B7RuMKkMNOGZcp8KzCDTxiqFhiEfNcVWq4EyxTyK96/qEB/pbFveXPLbbKE/O9Jp
DnAXmpRx0CChM3zfd5JGh6fMVqEo3G0Qp7ev0q8xkT9sW7/mJPETYNeCyxKyGODh
52/OqhxFyr+MtHWim47H4AIS0IQAUBP9uf8kombU8vRm/lEGbbOVsDaRoY3VfCH7
7lH+0yXuvZ+37wIudCEetNrE6t05qGoKqrG9g2wHxRldiCOZ9bT/Kc3t1knZNde4
qd5Njn3gXJuEEXURD/1Rfjk2SiM18xUxfoVfuTWzC8A9SOvsfcapsGgbq/Bhi6Pl
I3n4iG/pmSTifGrK8gSQt44o7VBzpclVVXQK1ijp7SMygEEX2UXSuSk84ICZvXQu
uxYWAAp5GDmj69kKQRIqHc8FgI4Ok30XTMTOLamZzTglIHI7NfGCpNbewmAKfY/J
27KmwFQxAIebXYGLFv+I0hUvWTVNvthVSqWIzG822EqIdWGU4J19i7VssmnImSsw
/nbfZFHH/zUhcER3jhQEEczRurQDG5Ue+CgJG8FUNfuDhBEJU3S68AxpD99YXKCD
7IMHuHF9vEhlaE+PsIm8OgXHFKH0Haku4MWaeB9tLs2GxJbLKGG3q8JDZ2G/F1b1
3hlb54G9SCDEH6p8QZ/bANyjdkkb8k2SuYKvF+tWZkIRk1RJYGbRExqjsZj3ceuK
uVvGCLroVjrbfYpGWl0HYY1+mDloFnl260GpXNz0/WExbJPUf9pBdmIleS6DkHwR
xwHrYsTMlXhyTYKmEPrObIvswm3vtzLXLfqruqPXA8RA1fu1U6QMVB+jDHdSLQEa
hfMzhSfnLwsl3eWGIoYrZ4kg+26gDnkDuvRAwOZ2ZYs2NHuI0BpDWnITgdypthl6
2NGEC5fRct0kRQ061RpMHDRSDeEreu1o4M74MeKYpYsjEl0kcuoHb0NW6LjfV7Sc
BY46r+FhLiLsNJWXNYADHBH9Rhn2pZXHsgoP9nvquniTgSF54YSpMV2x9ijQtLki
igD1iu7SqQudJ1uEmsF86itaO+YYXcHapC7lpSApGe76Fkxqxkv/JK8Jj2jIjho1
gzE/14arhoCwuwJuO5tKuoxlh0PdUhaXfnAoMSh5KKqs3O1aaTwD9mG5hTrI4vHw
fUqMMLPohxrPZMCv93QbV2cSU9sYHBCwzHtogX4nhskPhvRIeWk82AGGHCLg2Vej
VeAbg/uDVQo7fHbJ77OjMiy+3chrhgddQKcx4CdzxXPog/yEw97CH16saw5Wo8x9
cWzijxGFzF/7Tw+JM3lqQBmEWMPIm79SEwS9paUA49Q/wE0sW5+g8Bak6yjCA1QI
zM8XANwP/KcoOfyOreggR2to5IMnNb+XvofLEC/XjJp4akNmuCsFIbyup1BY+lKS
jMBMRQSXmNYz4gd2K2l9cvgKz+vBoYMxUilkTSLdmWpGPTMoWKQgAY3YWvTwnhUw
gY+S3Iiwv0EuazKvr+0VZJoHwEkIo5JDYR+7ECkEtWKo3OJVRmw7CYpy488OQeOu
aZujDYyUR4zJK66lojSJFXIFtmj6+Tj+Cs/CmfWlDH3YiK8HjVUf0YY57pa2SukG
mt+yGgoFCzRxjhr4D56lvTUHBkBH52NxWM8Jj6zvUDYZ8ZwSlzmJYlQJaAyhHd6e
NIbnnHB+LcSgzA3Gmz50twEcZQnvPO7uI6wvZJgyPSIJZ++752TDYnpV7/KnjjrB
IkI/rNLS15DiHzAqwbcfuOCDxxhBUM7mInRANhuLxCltr98TU3rIOHFAbUt8e/p7
3Z9GOId1yDcNVkybVjoGQouCPjO08amkqXSks5USjAVQrAysh2FVBgLEWYX2KWho
Y/2hmYqkCvTBRc1RhJHEi3qYr0dfeoGNXzaQ33q2laO+jepcSnkajjiW2HYE7zQz
odAWEDtmDwScedPE2GjcFGBY/0kKj1XvMItUzB3AduA+JZHZ+ew2G3lXxEeETnBo
gT7Hqfl+XmmFP3VPtPyHNrMKn+vIW28T2fGPXF1NDnwkpyehZvcSsj+bZwt6WN9J
OwEuZZomCaKu9VPgOp5i3kWZmFqITRHcz+1PFrkFrfGpI2dCvNRZsimZU9ctvG8F
3hg4oTg9urjczkgCnGfRHOa5SwZKLPwCZavfdMKJTiClXSWi1ZPtXIolrUBDyqtc
SBaEWISgjU79hWVo09vkNoibnSyfq/USISXBXHDD32HRxomoY42Si+0P6vAO9ebV
FJ4juFTCzgXtjp5l34n5aS6pLQ4khs2OMa+VmxNbTsxCxuQMcxZPZEP8jZqArIgy
M5Ukj4ZWE9jw/wajDnFTkRH/m3GeprIz4/zvA75xUJHdg50piK4htvqzduYyEUYH
Yh86ganGBLOHB6OeUNv6uSfT6wnI5ezVOGfwJWbc0Id2FSxfR+3a3ump8/TMMTGG
9tWYJ4WbTfdCzw2Ro7ubvgrIwvZZKYWnHPnF5r4dKJbpIQKEX/ha+MwTKNCv97B0
oJUnFkeXedAR1tFZ2LZX/axV7OyoRprT7iFiThcw6fb8eqDKCalIWdiON09k2JYR
Ekgy8isgBGACWxYha7mzSfMMpwZ9lRhWNS+/GVGxUPHC3Ofg0iXkM+PGMJEpp+M3
qjFe5UTnbdYnUwtbF4qqOCat+j+MA5Yb5izHX3KRJ7ic249r0S4psi1gQLgI/4Ig
XvGBhEi4nY+dukdVnvPZyErtU5ddHCkR7bzXtHJJV4hQOIBo09RVqML2HJtVYf5j
dZInv5kvFQ6fiqFNK2aTHqWGqgivi5BALjmihiIVr9KY7CXEIhGZ05/oh2US/3Mi
OGttHsB1CyPlReKBJ5H2znbri7sTk6lsi8tZ/LYipDS6l5eKN1i7sVEbhqwRlepq
weJRHe0p/rQgK7/wxJ1BiBaNkKyQw1kF6w7xhBpNGhVAWO8jxephdtII9yO53jh2
RR/nNrGNvmrzHIYkrQZ8zRU7JYmta+IAGKpktWvv93O3yNAzmyeXpIp/VO7OLLPX
cJdVl816OR0z1NfsMep//0pXy39llL1jdsNLHiM6+VznXSdIsKsnZbthnWNcYAyi
eR5TCwrxeHVGyhkBxcW8CEE1CZAB9yvPMAvmSMS4Du7yKJKq6f8IeTxXyB6J4plf
ZIRAIbXjdcFgpjYDJXcZLzFZrJDNakrxn/qJMENkj+iUmnucaN7WyOZbQaGkZ+H/
uKbi22WBUqraAddvObEMNYrNsnMXXHAguiCxAjD/PQfe2XaKqgxgmf4TkV2X5BYF
KsLhHCRoy8O/WWnCiAaM/Sdw3bWDX3cbOlA3vxO8mnGUEjb90P1FEat9s316TBdc
utT1iAzhIeuYTYXVJnwq/8+sKbNWdy1B6UeXDWDyuxvBHaCPtNSY52znqa39av2s
Kdzb0WGdl/nKd9mpfGtkUIb+h661D3lAG11hkuy8+Zr0fmCqOoAevvAxkixxOaXB
LJKNc2nqY8l9Qc5upd7d2J3ng8lZB5ijt5a6XSl2krzwPuxe5GWg1iuQ+w4A7Z4J
0LRuIGoc1kzsjALuwvpTIWTSRYKFfgjtIOk8YTj0evKhLnYbKYIB65B/tZMFEDag
DgRWq3L9OTQYRZvYaI+OeJ4CrYjn9l6WFgXuYbSbSl8A0SxFEW/L+T00Kc42HxzE
OVrd524lqqIhlWJdB1BFk58q4mIl3Q8RYvM1939GXwkhCNqp8Wu7R8cLSFS6HH2D
jUoe6xTRbRaqjLJTYB6vXseOGqLuJRIMaMaNzKHR2WsMAqJ62hYK4BdrYcWmWjlK
hEbY8U4Q53ZDK0h7K/bWJ1ZPXpqgKnKRQcHUIlXT3UB/ZAMTrqb5cYiA6xEi5JLa
2A1J41XDmVS1rHPtY+YUa7G4mywwF9nZZHnPD0chzYJl3liIvGNj+e2XqPj+cKUZ
2Ej0bghf/ganHdDKlSGdaB73yLq1pJwOsmQvY8sMYMeQ/OOVw4LSX5g773k9mdBf
hOKz6sAKelVN8FhxGFygMFxmS5NHUZDrWee8OPOVXWF69Mtdwjl/RXabsVM/Azez
J+TxtVC++zQMz5ewJoJM3CIDiNfd4Owl2awPTcaQ5Q8s3kKhRLGtIA0EIR9CyMFb
+8j9dWWQMZmC7PKv631hJ1TfbQXIKYCu+9Bk4FUg6yRHQBLdAPSyTpCKWg17WsM4
ecV+f7NWC68kxn+Hy4rAGy/zUy23+ZBvNxZuNFmGsz6P8N0TV6cqm7w3Mauoh0wi
Bc3Pe/N3UlbdlSwSL8N/86bLcdZeOp4x/d9y0LfqPj2a2hhRNR6DhzeC9+QUrXqm
FoNU0no/kTaXwKR+2OGpRTG/4TquGZCae1Ag/WHdixeCAXz7nP8j8Pd+N5RQJJEJ
rvuvxdnnakJMTbDa6CoIIlPFehZUJbKZW0a9rtgysHEjeO6TdckvNhhe7mykTZwT
aWuU2wuPrqPMrKLN7Eb07/myXa/Q16MKIYeP3Dwqgt745mNYlEAa2R8Oq2cuma8U
SDHyWjcj6eptJZMLsZqFPF5RMrGQu6sdCeN1s9AIa5V0kNh8rQsjcMaqj03juY8R
ycVKhyyoqPFAjjiYSX8w80lv/KzAec5kucVo+93pPs2OWPND5NjFu3kI4FE0UA2s
V/T2k89AsqCxsF5S2ZaB4z+U9Pqeg/rZ8IJNW9RdxZu9YU/7kF4a+ZQUPV0tlHF5
KJ6nPwB2oZJoewKYovH3lhzyrngaNRSgznxRbu1MzpqNPznj1xzUXC8UEZhwp4d6
L2VxLi4CNfyfZ5XePqpTmZp+zyLCiGduESluvIHz4BJluW73tlM7NDEpNp7I21AK
F+9YSpqPsufmeQY4Ijpabg4JQYc+veIsWw0BaNxHpbL5IN1gpHISdzNWPK02V0MB
eAnu0wqSzkRiUauQEe754FVQJq3uBBqzrDb0upzaeEGIIPBEB7oqJ7Gn+ngdJSvc
WDbjrSEmJHJF8orsJrzNtHw6EkpgZXCARSfdiTvdapCptYp6mxv9f4E0MMKq/z4N
ENCBqyooh4QVd8dzoFPuYMjHB4gHXpuzLK56kR6fo/dwA1oCCsW2WgZVJJ9Z+Qoh
NLbXjEgCQ23b8A2NHsDK4QGdSuX/jt6b0TCyuLc3OE0+1bPj8lxxWqHszyOC11RM
nAPeMAIIZlvjgx6Ap0BaLMC7KCpEyE6Cy5yt9ijUpdwOEaHQKLLx0rHFTCctPLfP
7kikzgGQSDaxCdUmWPqU0wZTN13acC+c8fLETKdKkfk4S4dUP86uF9xk1NajallD
sb0Sj+eJVvPyglgwvqWZCdW6b9zqATesAbLYf6BArVnRUlYuJvAgATPMUPSO4IbL
oc6mGT1A/5H8b7NvgmYLMhMF/TzZuzgLAUwq/6pBKJLbd0hMb0axSLL+DpbBJexs
6Kjltc26TXQTXGjOI857Ae8E/cID3opEbPLHZSIETL5TBXE0SPPlAVlDXG+M7aDh
kr9L4jIf1BW6GSR33YJAK2Dg1vpP2sTb1PTcHHDOKf04JLxSXAl5UXePhVN1YbPK
kfmMFRU3UeWVzlt+R6a9hgBeqsbfRJoDDCDDV5ViXvNYL6QWHdAuLmMHYqG5MY/n
9zcA0HzL3AKNjPTfING8i/ThKeVctVm1n8egt4aW3TrHNv6IKqG8tsmVVuPnONef
DNN8YFOcAQsq+tTaq2lGbv0dpOx4RfqtsHeUc0muHMq1VBH9c03MjcuHH1HTvWH0
UkvPZVYR9EX27lR5dhNlwAVwo2sUsLNUMmYF9ipHsx9uUabYpX7k8jDYM2eCrCvu
exUNXYNLftHV1SAU6wNnGJqArd0+gIesbzBlU7a1+Rh73Dc3ARUgHlqJMU5Kx+2q
YSahBU+tcSHvmYevwbwr7ZMxRzIe48oPST5xA8BFG2Aaz4TJ/cxaWgbxtkcqaGRO
jrmYXhxexnyyVzjad9TEHY+crvlsucc81JUDoQTmWqnLZkrNNuJQumTXdwIQre+y
cB/GOuaNm34yQXJtrkB+6fGVT2G2WQIuh7BJSwr1MDX7Iz5c4K7OV+cXor5aPvNC
DICtqPQMiWSgjheqXRaOPV7c8fdOOn7+Lha//lj0GH9qnjGj9Hwhm26XCG+Y+hVY
3quRvTZQY9Ka2hnBDTzzM/nwB9rnIvhwxp6MgYu3MyEjw/nxY/rOcZJ4NvYRMYuW
1u5fGvEx2tQaOWOfDa83rPcQiLfOAUXlNPRJ3AlovCDc8bAL/8XhcKsq7gIj77yM
odLUh6ofLa/Or+rPBB8egLOTDunpX1Trh/dSYMvY2kCVlhC8aSbJFfcWRfUXxZ6d
pS0cXcH1UiUAA4kOCtzCZd5f6dzrDMwBSKRCOZ3v3FAi0o+wSiX0fevnOk17lHmX
aN2QvjVOMuI5VLOhpKZ8kilzjMghbF7vTh+HtCItF+xL5Fa7s/scnzjuDfLs0Lhy
Qo7DfbB2626k9sMo5CllYjHvVsXSG4JK3gNBfwTKOc3L0tCagkhN9rMkGDWL7pNj
G7p3xOBntTMAMbOg0THDDttIAKvirQhI93C1PGDKmw3i+Dn0lnJ0DWDb8iX8jBPu
FxB5QhU7dnROoAkb+CIsve7hrGxIhSrSRnkCrEk9bh886jw538VyR9MFD0CoOdxp
ay2HJeB2nVq/d+zzE9d+s6qRPjGuOqbvqOZNA3Hypc8rvNChCjITIRPms9cGhKBv
87/AR6GN7bvSg7Y2FyUAxYq2VTTjnKWVORW5KPJJQMoeaZX4Hjykv2BgNs2+lOJ3
6jFnZ3Oo3k7SEicirYwPb3w7Q2HdGg7xOM7GK3Po23C56EFSu9tYlbfdPe0bYJ1I
+K2WxxNu5f5mAabSIpaD3J9gcu6FABI5Fu0VOauhDsiclUid5VjFPLGIbMeC9VJM
iOuYXtA1ouP8mBNyk25vnRYCONB9k3XttDUPpbOL/AmJTUFjaagKkIPX6Byb7jVW
abn8j6DbhSI7FNFYYVSiyOgRYf2ua5Sb9tpOTO13BRLt9QHEwmeJ83Zh7SQCiXyf
wVLt2LWNm+18L2PtVg8n1FKX7b4JdxmckmqdAdV3tnk8Y3D6lWvY7oZ1+IM0lNG5
Q/rTwtuFcu9GUkXFKyjyIbijKybJpkGd/escOl1/hAtVvWRbsDFZTClwkwMaqLNH
1NwY8WNw1NsCzwF60+VniyRLmU6m0/F/gp3VqoAsAxRTWqQ4Nbpo+8q1o0Zu4wRq
rZvGngGT9v6BgmJoeyFZL+dfwEJgGYKTh68bERaBlu371KPq7Lwm4fa1tpqUT17k
eNRghXF0Mk7kDOT3s8lC0p+yf2VzZopGRJmq18gCn+PvFM0vZgJoFi5J7ulzegiv
I3R6H4oNe9JnbUt9bI00N6qv7xxV6Hns0fFf3n8qiUaLAGnywYTq9q2k3R3aM7LR
psCEi8w3MeGPFBxkuPVIq4X+ZttdBgZ9BeXpnnQAIlxf+jUEor9TSwBM2PHP1Jp/
LcRuXp21mwB711xWgBiRCYsmoxkIYaJZMghuR/7p2jSuObFUcmcglZ7AZk2/tS75
4T+aKCR+4lWU0VUj28gX2jYeEzCG8smipyHn64+0ODVJlvApLnuGyDA/OX/uyvHR
Aws8OjkC8B1pJvsSm9WKM12Xp7OtU/u+Dr8DUx41qJVij9xBVO8vhNQMNLddRDEi
LVKodlk1cQxBq8gNwywPXtW+yTYoEfyxd63DV3pTBZhytgOM0WdskbdJCNEOhDEQ
OVpWBgoqP/bKqxM9DmzVXAnK/TLrv5aJw076hDyDLZ4vE8iVNgGvJtp76DVUSlrX
QMsC2vwhxhGu/fWUAdGaORUs8wzDFYXo0DxBdlBhD65ihJv3LH9ywscu5JiDimzB
OWz3uwXtzXEGYa2fdQ77uy8vhQVhEjrhOgL79AqixymXNQ2xDDAAkcv7dB/VbC9K
8o59Ix3mE9H/81A8D8cuwjE1nWRuXXROtItvGguXMrmbykxzcFFE5uxMeppuGlxR
nW83ZC6/NgNeDTtJ3dUfj+rfk6LUVQ6UmbrYg3OmWckdfhLTPO7epw1W2drkBLVS
ykDcvQvgGZYLE4VxrObZRcIJxhlFf4MxsxZSdwk3l6mp7YB/4zhyq0qWR/qFR/1S
a8GJTgTejKq0845Iq1HUju3ZbiYQltCmmcW6QC54LHVcxtTpMjXfFR4FbqUT9mUk
J7qwBR0CekbAxrWE+rYuTObpGFvDyU4+Q7FCUxevISeqTnq3JYAJIvRZbaUfuPEU
oN5q/T+RnzrtnMB/Vgj7fwJj7gPpycX4MZuEVbhyp1TZ/r2sggam1CNvykzRxrCn
yIrwE2vhkczfn9XYPKEB9+9w1R3urxSzKZpbPvyruL7AY0uefG+ywEnXLLnWhBFQ
fhdmj3Vrkmv4HxCju84lNqeLAv845kAaIE4mhCSN0IwIi0Z8ggmdpZPE7tRrZ10n
dXKVM0o9hpi5Zcpv6Of4/4lttBwoIAbtPhMt0CWQakT8Tp85uLyLuUzaX6IIQPhB
k067408stXW1ZRAcf0zcsji75XPELNcsA9lGK2AtyVbv+BlBEdSqpTfvocGO0lzX
l77wTT2VrHuLKFxsJ5F8FPcrckHhFqQ3I69JJ/YeVztWc869h8arg0iwJ4MWgpoL
hyhecmjdmg96i0vxp8ifXEV+FKk2yi86dJAeGvcu/ZZWh/XDLoQYAiAWtG/5eP+3
1E+BN0vgCT2vEOQe3prF+olViZ7+29f9pW6KE9m7Br4+655cCC0vldR9PW0gteVA
5UoB7o7a00b3I8soquxXW1dMPyGHRbK86iRdfbOi0iAYbZ2pwQC+xBNguT53R9sX
El7RqMKqkyp/gFvMHlPyfdABWbY7UwP3obcyCG+Dq1MqlZrV0WJJ0U1SMW23flqh
RhaO/VEflGCNXUjxRwL9tKLXii8wWUUSrTWMCghvHMa3nOMy83dC9acj+bGjdr/U
dNxwgL+B935D3ILsnyrei5NT6xY49Ea1a9T8+UOKvdZL+E5uCGHuqVohdLWYXNB+
FKZFpJx8hFz0V0xjr5G0ADHKg8jOjvH4Xbc3o3Un6buUBYGRoemCJtKU9qb9NZSX
XQmVS9B28tix4Um1PB7GFiQsVg6P2Lle7fqeJQQcmXFLHRJrvXiS1KRfxU3Nak0p
2mR0JK2dAapumDPpHYVkg2kRl5lW43vgZnhTQhVQ31mOZLvV/qLaj7WPf2g1zKc+
L+7x3MbmeMFRFp6XOG6XpcSEu1ck6qz9TyIJPWA1TF+WOVYCIM08OM7CehgphwHz
+66ga33h9oj+QzLJSI7l0Rpt0Nh6wNAWPZWAepCfTHv4MbzvVtPdDIdplmvH5BEl
FGY1IxLqjr5Tq8sYqE6n5qARlVN+/HQKPDuV0U/j0/HBIoQkgxOSQitajWB10z69
2lGcD8oR4DiwWAyLaUi5pSwgTntWUAjX2OX2GWdLzonGf9LZ8ZVN+B3r6YF57CZj
yjo5CiVQs3jyOu8tCCAhOryRcI4yGl6DcRLQUu8WkQcE1msSeOG5lB8TC9mu47SH
3voIxtlQoBhN5v9U68Ru4ixKellLi6Hd6P3DqExN9ZhlPBoGyknM5gHVkGlJDYwO
RGEjBLj+SC5MYjkRsF6LZRw09tsc23n3VJYDgSUNs5q4JNm47VI283JGb4mR7IyS
Gqdt7FWjodhKDmI3K2yV8ZGHQFJdLwCBXL1zrEOm9qQPUbbywyP58NBtu3Oe0n7u
2Vfc15O3QUqhhPtUGDOT2CxwFriLC9LhvikMuhtvNK4H3wXno33pLa8ACLp0K+g5
3U0AGu3R2thB3LfulS6CcKWgQC3BgL0eVNpOfS8/DIZJVYmxn6Xp+eC8Sbu/ZOIK
EQNBJZYFntw4byi5nE1SexN9AsZ+UMFukCrTC7Z2r4u7qWaGgm0Qvddit0WJHbNZ
YVso66yjCBgU15mT5pn4LbsMTz/MVm1sgxW+VliGSXAUSJELWYgt5VzH6RjnHX7c
rsXyWMGK+W5F5/+02CVx23hl3vW2l5UG6YBKumiSvJMPp2xNOd8aI66VkKuV8BSu
MrzE2FMNBTdiwJVRPgbPzkN89JisCNZBrFIfA/LOYa+D2bF1KIi95nPXNkV5XH1Y
KYCOQL/rsKdv78B+SImEMBN+tZjIxoa4NrwPCh/y8ZdbLvY1rN6GqXEl6J/WPmUa
UeWrpWWpZ4kEVqSsW8aCRbB0vkaJqoV9rYG1aAKZatKbXXXDGQrDxhh3/pqnbjd2
vX0EApJMNaRTUd3JUo+HIjp9tgQQChXRVxwz9EGof4z5yFULPljdMrG7q536Tb0e
Rmdk3Pfso6plk+Vs0oGdui7MoQpf3eErVM+cKWYZiXqzaSqKUpToSUt3yzwrDGu9
VW9UCjTMoeR5zSAAY6dLt4zu49grWFKE9qWtckTfbpIwWtGdKQwDSxE67zHgHwoD
8pSKuTC9lMIbrlofoKTq6wQdlDX6dTOIav6pVXB+NsVu8AOHpGeBlQtA6ThD3bll
4KbuwmVI+BEqfAcqexif35vcc4uVMI8OidRXFVbeG2kBwG70w0/ZMNdSVryIQUvW
D59+aP+eC+K0FLekUI6RSYd26ymtFBEyBvGvinEw+K2S2c8uCv7wzy+9iwiczug8
LTcpD7ORQvj/U+ECCZutL6GPplSxPWHvJd16riGXY//blndpoWXOAzciZROKuO7A
0Ql9I+Q2dONDUls9AjrKkxveXjdPpF9fyYD7rwh4ob/1dgxQXCRSRvFrfXSqTJL1
Ldd8PQ03uJ3Y33TAB9jGPF5MeCdRZtEWsgzVpq+QrW9s4iPE5PJTAfIVUK16NIme
LEZ74298TY2Vhimy9WalG/eNNHie2VQuLc+SOeEjd7awvj2qtd2zTcoHSqiZYq/z
kyxz/JCttmu46UH+qF22AZKY0JU64VRdlTCzeSYznum7k1Fs9wsLUO/0qv4qLdkU
ZD+W4aSuuQimksp0MqiPQoODERsA3eVRBSpcHoGkEw7jl2GgjO0yeIN0KniZ8CMg
8zWsaNh5ak1g6uptKsoLOgmpqLQ2NRqu3hCF4izgj59rSkUgvipnYMDijBXrMpUG
MwgAu4UOVT3TQs+Hq5CBsu9xP3Edzs7wfwYsFHt+hZnutYW/i6gLrb0x1m+qXgLo
5la1APr2Ah6+00L8/Qj+z/vVwLxSrPNrgxiluzEug/l/zr3rzlGz7ZTwUD8ZowX4
AXbtS6YWK+EjamxWPZXX2k2NEmS9SKcvUgD0N5iYgWJXrkH4BT5nApUFS89beTyB
v13sLqd3YHfoU+aS+kY1gOM49+iv1AkaxanbsePar3U12QPZFtveRRPeEfwzMFwp
Ec1Y660KFPgMhDFGTUtufwBMRLdx86GRaRWZ+bo52bIV6WMwEpBqbDiFJhpGtzNv
0QsMwdOlGJzoyQMlcFqWN4gPvSYfw6VXcIMIMxZt2hH3kHkl4v9euXbSn1dpwxqx
lY1gCyLIdSbJm4EJipt3uoO2kSC24moPO0udQFO6IAhPkIGgj12ITG68USBS1qpc
0XeEiWS62/NpIG59aMabuXSEUkR7VRNLTLmJekTYuyAviYW0RQgXejfynsIQO/Pw
9lzClQLimWBHWd7dgu4GoaK/3VzKv3GRHYHzP3GRUovQ2raeYr8OtszRQB5pw9Yb
nzSHRQd+ZhLdV5cR49CNcEdg+XY5b9FPIwwB02yNdwY/gd2IcliPTQE+7dk2ALf1
IlfBw05JgV/WyoaebSm1clEwPWWmkP65Jli+Ri60unhnnBELUAwQX2xi4jEcB4ML
bfJw/2lqXYYuP90HVxtqRqmqqj9Dq9XpcjMLzBBGUs0Ttc+k5Pm4wiBtN6X92BW5
O5C3N1C1e3w0vvYPwVpGCH+EsGCQu1I139SCPp9IvMaeyiOXImHQoxV1Bq7MUKWW
Obt8yP7JZsLJHA9UsN11BK5s2143W80fQqPgcHCCwFUl7YDMGMg3JDu45hd5upT2
FyyqHaz26U715mh2aI7zlUkhS0AQk0IaARN4/7ROsdowzIcCJrlIcp8gh8mZMjSG
9cI684A5NGDJLs9D/SErFmITDsNjEEm8fk8cRrNaUEVZac2mHe9MjCR59U6t4jwI
fN3MiwlRadVpEi++9bXqIbtvfoLlPgcS4Dlc2SdeRszYcgPyrdbRTplcfxXQaBom
ePNMY3DRyTFtCXWAeA0I9prmPfppa4sIPPey26jHRU6OxM05yEZaM1yU9KNOUGAM
GzTN3N9GEVw1X1AwQ/NLVwCLCCxtHCcvWO9RN9RQlgFJx/Jrj7tWPFQm8DsUa+tU
T4GV9fFhoWvEp4RH3goR7IuglMcVrDScePXJXgIROpd0OBC6G60BQII0s2zCH7jK
6Kjbv7qlkO+B02/p+duLpnkvRlNRdSrqkZMBsMIt7aLRsamlmnhNpfP35kym4xBX
l9uXZdULAuYgSj9N8TE3/lkJBRN+ynH5Wb/HFgW0B37FJvQkTFk3oRt1WnJIxNtO
esM65vANYq7skhmUMVJLoLfckIOL0vYVvz3dby8z0EXdP1CuZgFw/SlhtQY0LshE
WqN1nNIpwICrdh6pzr5i3/7zIyQHyUccr5Ptzd92iCP7Q9UCVQsXPvhIWGlMxY3I
O2K9bU1S/VtHX50On2Hr5Fl2HVy8c2ewgHXF+dW1ncg+jogeOUeqv7o2jLp3X6Ug
I2wu8ascAnQEvulgDaKu22waxXuNVRJPiEjTTOY6vUPfMxeq5NS29SlTt0O+w42A
wGSH+Cbz+QI29goC+l2ckeLSF4E/k+YHL++7x3i5APR/GSGybaZzZAEttv1N0/DG
9HQH5jhlrh3PPEyjxdB2fS9kTYIT6eJ6biRJvbxT3aG2rAB7GJK8Y/LjtFVPXclt
EoepykyYp87CNbkRyNlhapYmaFX4ksRZxr2wtM1K+NZX33/wsenc3ojgh5Z5d/Ra
p7WToF+LFt9+uXtmWeTWaRcH6MwIImf2B4jl3mJ+/JxkPmT+oiwfzChwQfEqbIeb
iz5RSCz83ye30OjNEZssPF5lpKgESnDNjNDjG02If7Xer5BQIXP57Tf9z/PVjkF3
3P4vPuDk/YyORvtgL8enCPVYKaMLB0DTY0cPnH+4om/YhE1uxA7Qhc99KYbrkXjx
Nz4HMqDLTyRQgKrowfMh6KigqLjkkxq6J3g/803LhDwS+LHwcan8W3LBcokYW1ur
wkXMcHIlBaec6tsMNrdovzIJvm/BXfEoEwAms02SqckqAR7keQszaPG1/zRc8vJ/
TMJLgYo9V6tyigTfRtixQ4vODBxfY491WrSvkjkGdLsyOXOUtk69J5YcZHQrpJYM
KmjKFOTNWJ/r6otMZ49+7cO4f8ds4We8fEYNT3Lx1ZvckePmb5WwJV7ObhkQmOrP
3KzFZbU5TfpWO70WO7tLxm2DAuCH+dJ+aKHBAhYTFoCaDUlDgfM7TClKN5sgMYIr
RtuIFIPyCMyv+MOdBOofjCuapJIztpNk6MEXlbYZgXSQfYkcQhX2XxHcg/9dyN09
aiT2cENalGoj03h3WgZyqlz63k5wCNk/gEcwap2Z2YlDu+5BTHfcLuptWmqSk5dq
bklTzUs2rQ60JeqJlZuyUqKb31Rn5dfkZicZ4kFaJsk7pZSfZCsYncrp1OcPy6Hg
9jcvaeX/FQ4SEnExymPhPGH4rYs3jK3JPNfDLmUw9PCPpOf3GVbYAzr6ZrpFSDRv
rOXtslbTzc3wjDbUGEwPS1XN10J0t2t9lIVsiOGT9Bfhb3kmMS1huuwUOEMVl74A
O8p4K5eX3KmTN+085MD1pBeGCHOCKOSzhIr//aiLnM04vF2NeFJl2gI0Ai1JFi4h
WdYblUSj8bg5MD5oWGVF8O94vf1cns3svS8TriS4rvyGEWPbvec8kuaFi8RncslP
y9A4y6NcLEba/OUqCeBtiSBOmTxxgzrVoHQwONyEQHcMxk59pzNmdupuhSr94Uri
eCOf2b1EYRWHoxJdp37DVmF/naWfgt97keanm3bCy4sfqGAMJFH0APGQTgxW4+Z/
WBYLIN7el8RUjNpHndH8KfbUx0sJax3L8GP1XRSydxVVXRWCsiknJ6aQftmP+rqM
HvBzxbP8AaeSP/aI2aExU+7hNq9uVXzp4mXmIQBXeUMA/TtqjL3I2rz4JmltAGsr
5+poxEQJri6DO88npekly/cndM2oS4gJHjT833+nlpwjHD4KgP6uL4zwO+ogIOhf
qSggaaT9ziYO1b8/BpATvFgIpnhSybmMPmndtrqqpCxXckwN2e6uWtaaL+2PL0eA
brR6jt02VAhmEfs5KZBHXjSNEdKF0+WNZo6rKMn0dlEEQBsy+DlIG4UM/R1IbzzT
kco2g+S2JrrBlyjulsR3EKmprL88zcYU27PSnPRm5dRVtKTL7QT9qZcHDNh9moiq
D3nebQ3irGLTx4tyYr4rLMkgp3N4OUj2PjXVtrkgOgbXxa6CtOuhAWbyMowFfG7U
PWlkWk2E0dBw2ojdP/3X3oluJyNEOctXw/k6gRfw8+xUBVcVeidHFBLfArzJ4qjH
eml1P7DJRBJaVxBkSdKikrooqiKCO8GiI6S6S7pd8TV0UNSTVhsKNvBPug8WORCN
MVIC7g4HHNpORVbRFmRcmL8G1bdhxlZNsg5W8ite3P0p3pd67iMmriqFF8GOhDFp
rpKpDErYo2VS2OYs9hyL+4cayfksWJUZk4gWOqZgctdsU+IORq5r846TMRLrYk52
ayI+ZOyYfEfv4Jj3GjnSMxF5dkYoa8Plydcjp3Lv34O2SRJKmqdYczlTi+Mo81A2
a/XrWz7jXviNqvdVTglpFdIc1Euc30JRsq0/JYSA6nEV2D+8R1fkwlLZ4A4uqdxS
gvPb6Ukv1Udmox7a3FeMDP75nZ/pxHNbC3YnYxKQIRtNQqwnZebqoeJDgk3TebmW
x6rizV1ubBze3jft+qY/x+OrtW5iKEGs6Pp2Hcw+erODcB6nmq3EU/1dHgyfqvnq
P+/BFk/q2Nk5/sLpjUsj9FmzTp6g6U2yDAx2dyMpGL9A0A1v4uOUK7Rt/xLMsbgd
STIVYt9jCh2OUZRi6dWrXTvAghG9SLqwCmgq0IBKoGRGnG4WKeZbC+lnr9Dk4yR2
crRuWaiKj5eP0Do09GMaeLLtVVVJoqbqRztOmGyiupncP02UT222Z1YthCB24B5f
vKctMMPFqyYjuEEEysp0ZLxd+/ZMDWgfXG9RDk0G6ZlJzh+DngPLuzTL4mpLsx6R
0DdBMVVEdRtgU+y0OmZ4vFPRIjkRrGp/DFYm9q0K4R3wTxa43WdTtIsBmK4RWAI3
5XibN6RmATpPY2jpE8+8oPfrH21siMWyiidC7kMteiCobv1qpLIrQb1RxkaS6drG
5Oo6fj3fcGP9cNvZ8GbBSAMn7NqXc9od7sFwuS+hrT18fq5iUUciqdH4iMpMc5RW
d6AgVhXDK5QuFUAa9xARifkdoe0gYSkjdnKYTZSmR6SZPWk70i6otJre0EthCfHz
FscHR7iIR5JwGDBgLmOeszc3NmVfUL4zpCW62rlNCVNoUH0dBOGm7uWCrnkTKMlI
Ty7eQiBFI1NCG/kbWsHk8eQydh8z/MzwiAn8VWxlt9uUHDZXf9+OeEbA7+5G5hSk
4C8iljF9QhdAW99C62KG3E1FJc63qofjdcvIVDeNkW0yKE5VYCmed9w3CjZJvuE/
/NLx//9nP/oIM6znmSPs0Bbm3OPAstojjIbLDwI/iW0D8ed8NiXV4s4muAbIw8nz
rO+ts6yPOB+K7QXt2v1ZfWxDYYTVwWI6G2740c/hE952MkKdja0GytEBz+Ct/nYc
ccKwsK0lwWHNiUSfwGt7nfChOV2nIJU+4HeIodQlxNpGs50sXu2JBVC8n6C5CaIm
kxHU9dupj5nL/87XY3cLS2Is52hN8MSm6z6lbH0OnmEzL9IlO+/EHumJ8Ayzq2Au
QAt9Z9XeuTKVnH+VtIgLJVN/Ukp4rU1MIy3mmN95aJQqefgptk05+Ki0JSIrSqQo
uAc4cYdkW7DiwwKiY2Qx/2eWcKR5+AGKMzIWpRboc2iTMCibdF8rgO7uLcEaE1kv
pTsChlkABRFIAu/ahQ/OylBsuqpBxGzobAHl8u5am0dh5jOYBXCyUUwVf+9mslxP
yx8aiglFUQJpy9m7PCUnwuHecRQSomNOhr9MTTxysQ2bvF1hZ+GfMhSSKtxBH5sb
sxtn0EN8sxtC5fqWryZ27/0vKxPKMcn0RqqeKNec7HgmaDR6QkGqd7vrt1PT/p9E
nJm7DUW5i13PPH9jXU/Oal+viFkluqKSILI6N32PjAdrFCco6XD8fY5YS+O0nUw1
62dhfaVOc5qcwu1aJUI3lR2WuCpygvMFmwTbD3nLFB4o4uV0dBYSf9EmO04TZZJ7
WE7z8dc97ugzkumic81uVZJTuh+gRNXI4izkPq5UfRjs4q69SzYGoo2Id4nYDLHO
SoLzTUWKvjalsdAEcUI1Ckp4BFJqI7kLc6cEAxywINvoJadAgIwBv1tlwScovvuj
ZA3xdXHRf41Rl4S0Sa5kzlNoDtOMpjjqfQff0/YpUzwJLOBaNzTtIvDq5bMagLql
s2C4gaoZf2T9RDXel92zY69q1WjPWnZV2+yH5kgH6i2k8pwuXseOs/+AQ7OOyUR1
2ra2L/JSu/VyVUhSmkzWuglvGEvzjNH5OHvwUNP+zSMP21kkKZoviQHLqH7sk6wE
t96b1LuYd4uQeS5mztWDAPIyspBiLPcMU8ub/7X4bTwxQRJfPQH3rTnF0JAKTaw7
k8FABKF/GfwrmwFQR04v315n3JASwCcFwnku59AIdOiUNGg9doF0ZhmS3F9+tsqk
nd7lBPKx5S1EzpdmnXRn62qBVlmO/4/ND8JQRakd+sFzTgq9QOUO3rQKYwYV5tdf
Va8BD8WL4UdLPTvdGJRTT4UNirHhEDBmu1ZMjc4lYmSPng3u4Niqhox7o0peWBaw
zFdOAQDBy8ftSLeKDwrQH0Jsz62h39VsNd5aqE2zmEJwiLgUWnfr2g67bUNcAWTu
w+SDOdJ+c+ETaTf3S5BYBVtkFcAfEpczGpTLrkOA5Y1D8zCLm9ztO6megFgXds9H
nZfW4Qo9yqlHal/SMso2erX0Q35FDHANZfLescI/U+RSzHbG3G2d4qgG6nTHLk1l
XyOD4pjxLJFMwHZoEreAwW9cwBAz9KRRxL5G+j/JHKRfZ3bfkxmudfyBGjQ1D12P
xBcNPKjcj30bub4y3pL+d8KSiBUUIof1f33XhM3WOvTa9/Hp+pnSULihI4PXA/tQ
pfZwx5weAUhuRDykU9+8InLNa0qdEP0fEhHKGoUsOtOAYEqS8chueQhHt/hS1gQc
BSqh3J1jQVW2SpjR1buYuTugsJn7zmVMgNgeed0hhwe/xULff2ZMHE63D3GlYxOP
qHQmpN0TyZ037NvOz35zltni3mlobc3MrY5N23Z4nRcgOnEtpsTRYsBtYOnBnAGi
fo9R1l1z2IblJM+ZoGRMvehCSxhGHLMHCWKEJ/CEhCk5Jf/m2DVpJ3VB+n/M2uN2
/EPw5at8almVcGDs4SIt5BL3AAvguNLRl/QAsTCapLmlMfdX4h0eHYnmGtpSCOZl
w9CVrblgCgJQ2fml5y0r3AQaoUDOMmlexnMUBS4A2Ogmhos7y9pP3ptgdf4U52ZO
j5npr+nKb8b+UZcOkJptanvgeaKtegDL1v8TEHJ+4r1j30FxxSIfkH5i276Wocsy
tC273XkS462RqUGVfURjOnzpXb1W+tU4H+eLWgmf7whvHhSVtg7EWytk35x3sPYQ
KdOESaGmMsIffEQhjPfRV5ozLO7jnOMEr7EaE83gdyTlyyfGrFdHL3IXccl6B54m
r3eCdtaDdCsToxtdh5/2rN1WxAf1QNZA5m3b5mf3qZnwhdlvzyR8pT0gUjIcChgk
WhKvehFbd4TWf5Sw06Zfvnl/QryrSTgasrPZOEs5pi1yFGiyCXDhCaO5EsA4Q/2E
LJhEbiePgLi2JZxsr7usSRJumMIvfs4tCo2jEWy0rnWb2qUQQw7Bo0c5xW4tbz6Z
+odyhJA/TJhnFc5xV3i4hNLGqkgx3iKk8IGzoxhzztrSEhFJhsqFr0Y3spwRJg0a
vmltar6ANYTXRas6Xgbrj89orEdrWUgarmkhhKlXmG1eb7JHg62a467lB2oVek+0
ISMqoLTYAc/nZtzJCcHVM1FKZjHOfgsvbT3vmR50vhBRdkxjMHNzJMnVHPgixmkF
I6nTFwWWrIGLORImeAoNCnYLzKq19GJLRHqbh+Tj9hPaKVQVOm2QndeLTkBD1lP/
Uf5Fv8dYk3dFj77sG0jvHkZcLTi/qFD4S2b6pHc8zSU1aoAJky5Fl0ay/m9rb5zJ
tqGgFNtAa4taqJCXp86dKV7Cql/3XnnmTiaJ7k7PLftVO5rYrXbVTtTJqARqu0SM
PoEf8d3ImKGiYmlP2uQVy1IVRrmXDJO5aRIL38emK+h3pejvGMRdtWlgxkS2UN5g
RN8r1M4v3qyn0sgRM2kjROhWPHYtsoJPzddLURjBmLYESKKZJ6iQXOS7Iyzz6KaK
9PAFmssUB8lTjPQr8/DPuKz4qc+2pZEcvDfwB7RTES9gOvh2+MzB/9DMZsnJ18e3
bgllgjAZPLqg0EyLy0pB/OXArUXrDbhCBReT9Xjh5/uUZ9QUzuTWIlkjHI4gTkku
b11PGmNzyKFInaFwgXoFZMvBASK0FC+PBIbhgCXrLe40jLEgFmFAMz6zFK8zroVa
viGhrjNKV771RfRhnh9dVNXR+o8xhHcR7A1MMewqF9juivgSxQQT3vtRnicSm2DC
6H8CjA+iUKGrWrsYtSc5iSyvZB7uCo3npuz1AfAIEKrHy54DpxNtY3wXBWtQoyx8
3Dki+VgrdfG/VS1VyyFHXWasmWJ7VNRJv6LLR8AnFwAFcez+ri91m6asbRocfDqp
PU2QuNzoLORhZ7XfN7AbpV17fdWCROEB/aVDIiWEELSrXgrRbXeGOoaLXIiO8+D8
SA10U6pU9JjLxl7mTR6YYk5mbb3fjvEyS1z4zajOZ8eqPI0tg7R6ZK60lTaOsoX0
DoKTIRZ5zNts8xCZPDuUQ6De6phM+5zmpRhGdjJAFzZ0G6QrVRLHg+NNlgn5VN/c
OxTIJUKeCMC3gPHDvz6HrqroTmXeuNSQesAlA0OZ1CRuU57jpnTgZSAfywhLMipm
yLq9n3cDyJ1eMM7+TdZvXiWuQ6BjHYJk+edXzvQPXwG+bhPB9OYzxWuIlqvWmcg3
0MhZGQNsQVLaJ1Zd9Wt5P96g46pHHgxRHtCaQbGRQCuLBp5IIaIEo2oBsYRGTfqm
1/qteD970HnI0nwB4c0AvY/hog0cBiOt/bYGlJheIka6Jy1FKRyoLlakGNMB4nea
m2BRuqPJhax8sUKr97yuqGU9THjfSo34bbr5mKNj7NuAaqEs3qoPG7lyPhM8Q5VP
XnmccBguzisUxhMvZ+eV+P5lXFR4YyKzH0mKLeAtmpVMATUVetG7kVINGBXEEXJ1
goLIaaesQgLExT/aENCTbCd46SreITAFC5pCBh3yEbyxi6tJ94yc3daw6vuMirex
36ty6GTwSMt+Qx9RCGHDnhgXPKcSO7KSuIFlPdVxbztBA1RK7no+IH8Fa9XwDFQN
2FEh5ID7GT1pWRQoMxUMsbCXBbnlHTlqqh3qA8HILL9BGFCA39xqtR1K0gVEG+eT
Yv73ySsi3DHbHVjVwXsHYstZNsStykECS8OXhB4VsoBO1NY/HKPUk1nlbMAawb4O
aX5uUJtWqdrc90aJqGZThGLCfRQifmAOx607auUmaUm/In9RjZyyE0kG+XNOureF
G9h2AbCYNvaKm7Fwh++QUSLFYUdRuu4Hd483PLIqpXrZ7fvuC852oi4+ebFKE056
8ZjT+2z+3o0oz4GalLtPUvKKj9/KQhBmlm7Nd7iSgkOjekMvr76Ybkda6gAlQlB8
YifCJ0ADGiXcbQaqaQZ94IUQItdM+gZz6dei+1OfGESIrDhkelAI42zOeop++cMr
Wf997EzT8nckr1w5daFT/gzLBjWe9+ZBvHwRJiXLgNnSUv5xcrUX+gEcWzkfw3eT
OkaHw+hdcXGJdcOW67AdRdWGzpCjuPNR8rDjpf+9nD/IzLkS9jKaW5nRGchfl9Px
WcmbnAlH8+jzaEZSbQx/We+eiUBI3hUXRdabSByEAZZXjonfBRnb9AqxAjM60HIe
RVa+dsAzWRRHSBjzA9pqlNYvodxYVtcPg5WTe/D2jxFs3dvSWfEKOB5a4orugh+s
ApXM1Q9gfXFfPyZdDvMYIhqakpUClMTJ+FYcbBfIGrclRDEMuGSwIG4gHfV90Qzp
eD6AMLHvx9trzKeFHFQlfVRqcXdRVwz7cp2B3UcjzFNMSwVRL9C0EovnKTHu7mp4
0pFLIzjO+zVKlfkaPry79JP0qeShgzLLJdb4qZ1N5A9BIuILViawDaADJkx2EDlS
2Jj5AeSMWnF6YbDI34NmfRzeihrJGhwjkXbfJw3H+1EcgACvPlK32AQt38jjlmzs
xBvv7uHzoAH+pMvne9W6Npd+Pc2xVYuq8Fg/1zBSg7yK8GsDMZD9UAZLYOPL70ra
v2vY2hCHUsMmF+itu7blCvmRTAroyUCpchVkSvmgB+mWvC5NpTy4Zwv0uJYzAIYs
hVqYyPnNNwcsZoqk+bqU92A13nGlIg+KUb1+85U+nthroxv5qLaxMQfES9Xs67x3
GlRwhUXhhPQYdctWx25S0fIhr1u5mC+QJur2Nb191bHusGRIwM8yxJmEdVFlQ3tC
FSEIPcU6w1aL+da7nsKaO9vf/taahwxvD54OGwQ1bjxOb/RgfMGl/c7ggvh2mOz8
2OGVN8KrydqzqvZc9wR8MHRfPnV3zMSgnCB/gLihZyAilldC7M73nl+IxWnHWsx1
M/5kzqW8sA7reW9OxT+1rZ/pGWUNv2bD5zxmgWLC0/jCCS3sCgzw5fBUreoZgEAg
IuqPOq9/7yDvxjEss8anIpvlHBXmK0qEY7pjhVmMPdXNovKVt7qE+fK3mXZ1xdg2
pNNo9vhHC+IkZkRGZFjEY84Bks+gs86ciczkUHTzBexVDi8y9uUllY1Mygps6zax
cZ+Tu8q5AodLe9CAAwdmauk+FwVxIil6rl55fZgZz6S2Nus/YpKJwLBOHin6uzFS
IJh8yHis1Cc4vB4eBGzRDKpQwhQf8yZVinv4C6CT6SNAsOIx314ZU7rd3kKRKNBd
91Knc7YSEh7+gkju2Xnsjosdgh8Y+AtRukvnGc/eXC6nR+uspe3TBWb8KSxdYE/H
PiYCIVqWDdtcjmSQ19Spx1Ol+je2t5XqD9Vh5kfVSaBPSRiX1R9bD9tnlpvSq0Cy
hJMw4a9X+MmwUXBV6PbA+ttAIP7gvTgDf/C64VMeT0CM2Y88QtZZFdRimWChvBIv
GVbzGVsl2AR7Tze+8cMVhLbhWFFArKPCtLv8uqTL3ZZGX6nsUqAWbjPDV4kXyKEB
XnfBjOFETcens0P7edPrucl/hfCn3ETUPRe+kzN6bobBsYBDBwBYjHXCeJaQtAha
AkG2gVFbGBiJiqhgLg0UUw6dWG3FeMmC4qF6o+qtMXbu8vuEbMYHQwKeHOm1Tsin
P84gEIpfpKYgHNaBAoMSjGDOCPKCi4mkVM1m8zsWi1slW8pn2jBIC8B2fmwqtTM5
F82WzymhhwXgX/IlVYttaMZQc/oABSkvYGDSEkesca8kIL5PK89i0DyoXDrtAIyX
xcpcNhrazmLtgbtnkrhOlDCv5kvbHw4Y0qN4Odva6r3ux//e5nHYg21Qg3e39DDx
k5tySqx7eclV69zCLULO/y4SsRUdFAVxzVWQcIUGsUtAGQC2VkYKyMv/5LTB2LmS
i3WTTjciNAhcYJBHrHjyp2m61A3JY3QsZXqSQ7Svy8FTq4+TNZO1hzN3n++6VWEC
380KigbhEQcwlpp55xI4HhzbHOPwhMLoPsJqoTvzWfx8mhkSVn6zNcLvvVA3b3gz
Y9w8vYVVQd8vSGYGGEBdYD/lECgZ7G4Er6MfrqbR16EUtyPjR587enyX8pBR96ZY
L1bLETDPXAm2Ldx64Ye1sWJPJHgWUxbHbzQ4iNf2j14LZ/PD+04spfMuiJ7y0EZB
0MVZWdcunQhJH6FUXwtOckKg4uucdkLHXKjj7EpefBTMygIKC7ibXMBxpv08E8fv
gvHrMur+VhWYYM2+vflxxrUbaGFd6mudbem6YEASAnM0XRxRHXu1V0vx/8MXX48l
tDGocbRttw2CWQRNNLpaIa/sfM6j3TZZp5AYVzBx1xXqkBi7nw8LApAMiR07BHTI
MLbPfhtVmGqeaQTbz19rjzc3RNvapg7l06oOzfbHLL8bO6T4YoVNW4eHdQmmqfWj
KpN+G/k7XZclidD33a4lBdExuu0JQBPX66+ENeYGlGrhUHTYebpG09sY/7FE78f1
QrLfW0WZRjtHdvUIF18yGgaGgdymheXRW3PDI4jpjmwIqFGYNM7lEl0ofwtUZLa4
jqcNy3/tIRRovOUQY639Hn46tDk/sQK1iT1GWUvCbRlmiuA+3L8haFZXAJFjwd2m
npLgaRM3ISdt7rmfXsu0fCzAgtfOrEfTXSwYUN8NYG98weeVtWMsvTmCKrXBqWta
Y/cdKm/waIShr0K9UBFUY0rITtjPE6FJZW3Iun54TkZzyXYj5mkcKlOLMVVhiVrr
kCVcRHMC+JSAdxl6jCrHGHH489SjAUZgI4hXQESgFJvqBos2rEljxsCw9AbW0bEO
RNuLo7Cc+P5B7DLydEmIkDzO3LSsQ9+VoQH0cZex6/Ni+er2+mLHasFmA6L9g20Y
PRPqt8SdxATYD5LLIaGYaWyXJrFfb2zHEaWv8kKOWEExTAojtG6w96PFECeN1di+
7NkFQap3xZV2SQbWB+G0av4DqmHdXKWni5Lq1yzMtMo+09dP4cZ9B3Z2adq9ofCs
pAk3W1l9NlEsl+JndcT60Cz+pTZrCn0nrLBseRPeWkqsyi2ORO2ayfkysxBj6jAG
BzxyAMYXx66kkWxbZhHVYpVOsF97dNHuug8FzY4cvCv3iv2Y6fmngdKFEbnvuZ9u
jVhdmRubEBd5ykisoVVI3Ox6ZyqpeC6na6pJDEVwFo20f39L04Cclol/tlAqiIKB
P5ntJgubOfFKZfxPvr3IhpQoWolUvQnUiSSka8DCk9W+sJGfVEQfHqFMoWiBHLnp
k1s1xLB5PzVTMmW8/5vcwHKl7pC5bqfeB2l0QWI1rqiumrHQxwjKtXF65uLOkXIf
XwkYGS2GxeTzOxbP0O17yrFhQw5FCPD87ejQfjNriZ6M53dsF9jpxkfWDUJxAAY9
l0b1UhtfAkOYphJraV9ltS9hr8IaOTFvnF7w1kBudhPIZ5ucOjOAUqAbQtadPTwH
7BnpjoyXqHaaXk8epf4D3SIVs2mEjYAUqV2RiGKdBSlPXnX1pEqNXJ8fXh7ByvBf
SqX5SLRwBQQeOQzSeApIHU+qIQ0AkMViVDokbSuDVUYveEzfu+K6axM5SYchl2sF
fYJQKbeK7ctbv4kluviLa/93UJ1yrPVdWTKc0mVOp02yDR2YlwZ8sM3dA8hSNE6H
ndf5FzxYnfoiVk2PfbvrWUB8bdXk49UDgTHte6SY9gw5a8t5u+2qQbwOP9GJiRlr
mV/OxaDS1CBf8XcfMvji1JwjyyfCNHkh1gYouKzLMhaF0F/nFIPRhdMfM0NY1uFc
vreQ5Zqj1PaobYVBQyF+/tMDBoAm2aUfXk1TecfJXUW8JUL64GEgtdLteD/xbnrv
W2O9DjSz2J+Z3L+jnUVy0yStleMkqQnFmPppUaNcBdSZpfvlnNUtfi6YMYpE0U2/
IYPUtCzaErqsmjnHjxvieV7rZdhY/jOcxP/0S5dssSsV1g7YosuX0lUILKJDS9Nc
uElT9B/+B7NzUDtVXjih5FXnsEInoz94rtbuHnD+fugNR1ZbIL7WDP5jjQ3/ZVz6
8bWeZJIfPzkKZYkMQYOvihsYj1uW41LjoHQHBLKLvh1zTXGHqIBHIYyVCG3zMM05
TS7JQPhuot3B/1WX+p8pk68iXDTl7EklXasS5gPUxe30+bcPucUmT04PeofC2ysF
v/eMNFUxAA3Rka+jEEjxIpHvcfM3PjZXBO3dT50Qo2/Zd4MzE8olAXFQY870PA63
3Aw+jmDRzRZCrhPVUtr0NOpQfVBMd9MIjhX1QyDbPVYCA/3uI8ze4YwuhnKl+sOB
Zg5hqPY3hrlU10d5WTa4mNyRiFqAVrtsjPGL8ze6q1Vyx4cpj8m4LHFgqC/QO5y0
Y8JeWIl4vc/MkULDEJ0yLDpsHXP9A3JVs83OKEIMXPHeLcYylFPrALIKGNzbDDQz
+V6eUaE0E2sZ05Vmcrf3U7QVUR+dDcztuioNp92t8omAbxewHB7VKa1XbLHqSEzc
z4yMKRiPCm9kZ4l9xP3kLbUzldXoLFFH5FWwE68dcybxpUNtdIoLt0+uCtQ7bpwn
LuoMLIVZSG6PijQ3G5PwNDUkjZm/MSklHoId/U1PFvn5I41HNM9zm6tdtMEq325V
LyleVoFubTTEBR3UBF/2UTpkHZAZAzNpjEYRqQZPT5LTuYHYvf/StzHygI9Ar+ka
OlcT1OLr077QAyfsKQc2zZ5BvZjZrzjTkxl1mtISFx/5WyVF2VzO4tHOZUQoIGAI
0Fsm+fJZCZnMPKZBLUJ70kofCWCJtwlRRyNbemYR/3GVAL9+baWj9swmS9RlP1hK
KdcY9uo0FpOz6wg0mAFH6AGPdRc7rXRVSxsOTXVfveJXmLPnz0DEG6W2Agnndpjo
PvRA5z6+zwMvIdys15nzTgt891G6zjGsDUS7T/KQgi3Z7UuELLG9v5nBU+8f9IPn
kDbn+sagD25b6iYauoeyjlF3bktJ4km4c2ldxvXePCJR6enVm83irWHmgPHBeJzc
wF2ECgIwNB8W0DYsrErOWBXKYpgtD96Fhu/BZkkbolfVPODasdUUVgII4wR35aoJ
BD61NxAn/jqxuu0zzuUzgFg7195+svy5jmw7kyIPr34az+ovqe4e42HPn8fp5vQK
nY79h0EGaLH9C8770+VJDANXRpICRU77+tKkHv2lJw4SSllBq5AStYVhIdyODSCp
A+QjMdh7YOG54J2rJhuiOyJINw43l9vZJRys+stTT9r7V/N3bRLznl2DjQfPAxjA
q5y24zSPBJKjmhjT1OZLO4BJKG4QqTi+/Uc0EQr7qzzgQ48vK0LWQFgi7o7DvFs7
ul7TSFMjXbAllXHAYFxcPHWl9ZyYwuTWCzy8eBsMoClvYMi3blVq4b4fG3n/Kjdj
1qBL67XKzObsSv5rSRnsP5r/ziMobXfHtXfeYN+nFDluxBRSNbax5ZyL3WGj4emB
hkLytSXTJ/NtAHb/OmeF+n69Q8C/5LEXuAZU0KAKoAVf6iPrdnFnBMcTlYRiwWm6
dlCXHjlEOkKgSRvdbCIh+EKtAhrwgslIHKhy7Mj5uwykbShOIYKYMEICtl3ckTh3
Y1pLLj8NC+baVfUzrScb8xtZeWEjc8spZnghmbRjLaZue+MBtfzftIdRA2vgDH33
HVLgoon0asU0hA1fg1ur2R8+xS37A/MZjU9rLdd6orvWEYG+oUnDCws7buvYrGxQ
ZpCL0vKEyl91FBkV4LmmnAKkbe9X89twJF/w6g+W1Bxy2xQrMuuDtFwTc7munLD4
n3RO0dLlgL11tHiQH8yUkOCU3YuUh1vR8ssOnPgBOiYmlbwawdONoZtGoEqVTN+D
3Ovff5KEwLTm1g4wwse2Zx5wCFF/dZ34uHjTyd7khc7XVWrx6i4NjHIZxBHE0Nfv
YFXd76ZW4UWNNy38NZILNN+VDtU+u7BpRigcEy4bt3VYjaaHeo++STUYnytEq+Tl
PfZtdJVQSuR8m6LESbvcy2EfgEFPPripiGf3JTrMRurovHrYZjMVHSDgttYGt8ns
QpW/9ck3YuWs9Emzst/dWQdFQ1jue6NZlOSUBiJ9J+IR1CPgm2fe1cZxm8sUfR31
p5K9x9Sx56hHdHDHuQ7Djg9FFrjmR0SROab9HOtYz9ONXWV4R350eBEJAjAVPINs
IqfqTTlzOr3b6mbVxMJfDa/Sewzt4hbJxv0rSRR4vcQmvKiuhsrCqhMt/SZOu168
21rHN3HjFolN5y/rdvsvisGivIfFMpzm6d2oa7227m0BymhUN3m8gLjcNfy7P9YO
tSXik9E8vCSuIMnOxHXVl8c1z3+nRAckEe+asXyQjEjkuTEFSpMWA9ehbg76sqie
U3hZfxVqLql/9fc9tmFwCu7C2zjpiqKhjQdwxWZSBZDPqe266fLIOCVrynUuQ7mP
kesZJomrCfzwikeZvN6c4/FciVNE3QyG931Cedb3FnVJG0Y4W5hmuIlt90EAWA+1
oENWUzy4QVB2KzpBEWMchUxXtgBeKmpudT7SFaANwI7q7hfTup3caCpvKZS38TrK
M5F/UpOUDlH4fNumbyUX63CLkPxJBNieROzp/wDkHh7FEXkehwyfZ17c1MGGn18Q
3gXjzMkljADJDnAvX/s9hdH28oOcyTHVrw3PJHB992hNETom3WQAZQkygMKi52xu
uAN5sBwnccOZDRrEdt9mVPhdiMo+hZyhYkf/sCtS7HYfsBoZ/CaYASqMijt/in/6
ao+eBChzZ4UvQnWxbP2kf74YuAI3Wr0fTr0le+I3IWjUG+AiSw5UU1v90aH4aA3C
uPHsZkq9vEBjalCq+rflluv5mXsUo4iW30wYCPrxUCd8o1tZJKMRWtDEgVyoY0l2
3uHMacLhrouQdUpgagI950H2BMtWrhz2zvNouH46OGW6/o+28VVNMQJz+zhCnWVs
K4iVcwsMvHt3ikIJ689w9uAfvUX+6ecn3e9trDMytug+rMrg6BTz+HfUarI2tfe+
6p1xHk8yhyUhHdl9jy2/ATC3EJKiQHsZAKlXQhF3u/zMjLbVNfMxTHgd7JJoBxd8
hoPqw4LBSJe7iIJ52uHOpoM13QZPjyc0xbq52gLyeezrRHbRvLZf1YCXYpYFTT3I
ZVHQIRjAgHd7/diQbdrWZeQyJVSN7Usss5tYzLjabCCymIxPkiPqkJzr92u30uo6
gfol4MJ99/GiMzISk0u0/5gIWewLydttm8f1AX8ynaw1N+dCfT+EAc7o+PNR82Mc
z22uyuVwdFrbyUkP7idKxxPZUw9mU4WxbDG+2RmHb0RZ7Kr6/XZReRGnawQhPpEf
Eq2qUjzEP2YDQbAe0uTaVSItQ9SYoSyWH1cz6jz5A3HdeVPYTe5uZPouRTy00k2C
ssvID50F3IZHJW7DsevcxSNyrx8rx7/AyhgoU7HDdH2ndn1Pw8vm6dHgjzA/R8bV
zFKHTUqUQ5/t13lw+tLut3Yv+iBh4PBD5b4ZtT7rffVqUCA3vZWoh5s32l1Jxpvx
b8xKd63f38Awgdsc8MbwBkSbgQOvLBj18Ff/uA97PYzWLOcCYCXdD2T5TTMyzgeU
Y83UlpxWI8d6SRxlZsz3LoOHXnfvXllMH5ArSBsUbfFbfA1G1PGsU4iY9A9KBzmU
ZOJC6274a8qjNkre8I1B8r9s1yGzNOYWS5Zz7OaDlTjj29Y5AdcoJ0XEWSgWSaOq
Bs7XkxeIJy3uDD7er3M4t7Zl7fUyfVZ5dJlb/qXB/Ddig1rnjVSHtK6ngRP7VkLz
YXqVeVwB0o7LrX0/oCcQ/WMOvtEw/CrKIruCAKlTJpe/mLH/Ytyw7PGClB975Yer
7kAogySxIdXr+j3F7JljFhLuB7sTG5XHAqcVbkSJfHpjcmTh1wdRQvk9nyYOKnXE
BVTONRhR6Hj//jv83vAlSdNSDhUYIlAkkhzCw9XGCC5MznDYWqGFMmAjnypnKM/A
JulfKqLFvIkz7Ns/NZyuSGuNqqzfZrg+pD4fSQhb0u8JSoaAj7rO/1iPduBUnK4D
a1a8EPvuG0xj3Sqb+ttTUyniVB1Eh4a/6PzrAHH5L7mSHahF3z2+outq5Ru+yIa3
yr1M7cwsZJrYk1+x0sRGynYor2U/93xYUmdJRnnDdk4kudfC3VBA/pHv5Ie9X4kC
7OljhaeoFJutSGiIjA0QXHnGZ2GK3c2V1QvdIysgRrHj1Z3sZznPYYT7MvYyzgek
k9wIYn2V8zxGUR9gSoZJUhCSdditLqv6yO33pLX184hykUm5Hwao+AQ2c9GxZfPy
0pVv5UFEpeGfHpWDZe3ebpHKP5O+QskQpbDR4lktLL5vc/C07GkAgdBr+G4WUGVi
PC31H18SqIGXVzRCLm79CdrhW0Cov5x/p5UMlgzFdlnfhWgBsxaW5XhXIS8Gg9/x
cvjOq/Ighy34/nHWZyj91mIvaa9EogjEmJOKM2kpmZdCkQ9XJTX/4o+A+NRCM2vk
QDhK518VddxX/CRONzjcq6UzamzkAT32YgKpx6zUBN0okmLwOChLhoNQAnNAHbIt
6Z+1WZPPGeialL+LZ4+TUvJYzocgiqGN4hm9jZuJ4akZH5opx4kt8q0fiFbUdk4H
snuwqWkyDQD3L1uM/+uqiLaos0iuVJBnQWSgbBk6PQtj3JUyV18CSaUQu4jip027
JONh13EXuyDNIMzBehd5ZIwM37ys6E9vYmYfkFJjwMJS0f27TL9qH0lmVcglIK4/
HGpIUI01+WvHQguYy1Ra8zj8vQ/Zvf505aOqCz8u/bkAveo57N+4RB8i6vV//6fg
S//G4XwZmpY5hqrhTh9fEg/Voc2nxuatabE4Io4i37VzA4Kl21FM1liIkdQ/IINq
XF87533z82med/lHv6OFZFQFb/Sju7hf4GwOukbG2WL+9ZsENuByzySTy2bw4bF0
yaZfWVtvoK/gLJd0rnEkx+sIlspUXNR78wtcEeNTGDA/htYsx+WuEElw7EjEpHx3
0yipIQdUccsmIVaTb9Y5p7Bc8bHxZ7WoJKFynjv+47Bf3OFdMlueVWORGkTmgJ1m
b8raiQ5JUjUUcEvpCM4cIG+WgJRoMD8RjkAjAP3tz6wzjE8hlQ2yDW3YxJ/g3tuU
nFAXx+o5EKN7MgJmuwToge5KbMFFpWhUfPGTRosNosBvrZO7QLGW5jw2UgJxETip
OEBillQhKy1G9S2u4pvu5ck3zSojKsJJvp05U732ynfG+k+2R/zJKWu9XFNX8PTl
/pChCx0aXx67tk2HVg+pfdontxfGVqBOHbOi6VTXITH0n7HO9E6dKSybluedMTHj
f9o7hdk+QK73BXFvPDaNSutDWOPn8P2GMTPebMYT6rXP2xJiYZBnjM7lO19/e1Gi
d89xjMqfMX1D8PVKiVN8fKebpMxPnGXKtwI8Dc6CwblEXzCM9eaqtkl5zyVX9hlm
mhyO7dT4C4/3PbPzhfiHdREATpurPXL32hZiXN2WV1319mnB/kgrWeCTQAcCFjSQ
AdXR2/xi4Ku2fePSbLfYTQHRfx/PQwcyA/pKjR8ZR+3psW0+oWIyrDBJ/gJc/pDi
/QGOmdtCcCEfmleOXJ8lj+rwRaugBDE3TPMyK6YTTZpegW3dRY6X5EFpQDr4uumq
hvDxyyKS85QplWHqTYmLvMOWAou1XfkHYZVPMaQLvYWvPfxwwI4llhSliGnwtj/H
HG0A7hNYe8dC0q4PdT73VPBb7dN8NVVHVzraUdwwLEgNASQ+P3Np4mfDb6LKJX7Y
BfPwHq//CtXaHNw6gLeeyjOffrv9UOS9sGsGM6NAATl5OJm0OxSsBnsaivbpUpOx
Ej1FVSZkUiT1kP3wqMsbkj2cPZDJ0wocB2uTrzpZMxqtFe+PnG5bte0jmb/k4CP6
kgM7pXsIe09VL1agCURgSqkBtyt1yYDCbVHf8Is3NM0SW6Q7a43ZHpy4FBD/tueD
fLTCw+ClBQ1zDMHoXr6tyBF7DXehjZzIuyeGDu2Evj8jSaHhjXNp05JM11TgQSnn
zURIJxU4iKhbw/4xcCYr2RLqU7ahjyeORXxdAcEbKfVwEKtmLUWgdr41Fjn9PNx3
PpdbXCpDlmK/TUjdKBFtiMIt5NquOuLXwTAMfHLovwzwfiKdGrVVv8nUbCy24qwZ
3E0dc9jvMzGPJKyuhF0YUO5xHvoXTa6VyNHNNzoI6O8IGJFQ394AWVGjEf1GN2Mg
YupnCyL4fW68m7clGRQn/dx4PURMKEh1cisUvxbGcXFycMBNHulUvPwgFvce6zAX
x7p9H9dDeW/htNhqW1Y72JbR1fRTBVFAJMFzsq1msfUGnYqVMBQQ0sAdiWDN8P4T
VszrLbvx8J/Wrdg5JwrOmBclt7N/g9I4Xl+tsYRblLOiYbt4rPZYOAxP9bHVMjmi
h5Wh/AJCUa8jTAH1YYlmrxQmGcDGehgMk0yUQlhm8eU3dcuNdHDMBMxoDdXK78VS
rj8lck5fDBmJvgVot1aZEN5OPxEmJRE/i3VtHMC4GBzU6DgyzlcUio96GeDO2ciA
cWtJDIN62GPnEVQP03aymOcw1kSMNxo0smxTzO8sEFNNtyG33hBIaX75fy0gZc5F
eWqy0amfJb/C+keA7ReglGsVSO/paGUUzZrqBvIBQtKlqPMsi8u19jemnzFCkhCZ
+O0QRsJPbjDIXjo1TDND8nEKWUh6GArAHrtfm9prOmSFpg0UGIUTtkL8POi1Uy9X
g3CSFqJZxnfSX1eht4Az/pF6PMSFSfJAxVe1I+hzQLnp+XF6ueOe/2dh/c7WbjXU
SJTcdZDGSQKECvu4qdv+QVAwpVd5se6pcm8JjiUZqM55gJkveAWsSgHUZi5Pe9Dl
57ah0ZtIohWSxHvDG5tt2JnC/yFi/0tgDtzVvvpbvMyGfJY3tOTfHHOVWZDFPrKn
ao8nYAnC9h3ziqVsmYK23GwC90FS4tzYuyMgDRs5G5p5eCTpG6sq7iCHgpQ/zxEh
FxlnCXTSvn0POBLlnMuvsv9SFv03tuDPR2VmWgq+rDc6xOfx/OAEDzy69PwBUFzU
cOUptAkubChFjoKIqgMrL0+dytVVx9bOcUUPYF76XaO0BGq/U2j5yXYtQFFY053/
BFAhiRHLaLiZhdtdmpweg+XFmBaUvR69F+H33iz03Fp4DbRg25VTgB/qGGFn6IwR
3ASmOyl7zfo+GY525nphJhKOJfuuXm2G+cztNd4CpCxwVLouJnMjo7ffY9taf4mT
VJeBFn4jplemP3SLiG8Pb6PNeDkDZzNJSQAINMd3Rq7l8Fsty/Miaq3nu/AoKt5x
MPuWvHwrrY7Su0lZu1CGWRdB3PU9gxSQnThgieEhtERNq2hWTIOZn50OyNeYZjGE
kInvtrftki8Ge92o+IvN4aQLURjeu2ccnMSQKMjcE3H/ppDDNoGekSnUX6LXJsZ0
44xpm+6MJgV4Oy/NAm0h4FHqjQZzD12yAFBC7KaHw8fw6mn1fVtjHIGLTC0R/tn3
dkzw/Ecu044JisW3ohoN0ib4ftR0B07YMzbsMlOw8xkHiBb+mJhyPlAbBtgCEzCy
Z2nW1SlkSFSghUUA6PYzQyRMZLUj0uLoqAAoMkJy4EbzUPwQv36YpV451kL/OwSa
akKf9Zua4bxzdLeTe00cfBi8rLdhf88xPhjNZqOZHBPxwa/hRNs3ieTcLMKZQ4oE
YzDjWRbVZv/zncg/EsYVJpjVV2zVg4AHHO/+UX2f99ueuc4Dsy2ME7JGBVSmRebX
/LP5nJFxMX/k1kNCkc9akVW6if+DjYGsdB/YcOp7876zmsCZhLDA54WMgHgV0Fr4
t6vd2j7UaaLF+rtMyKx2ksR1i1pqBTZ8DiHp+3p+GFveiS1ZhGL2oL43DoxILIKU
bH5YSirK83RZDTWXQnRq/kFTzj4wjpZiXJCjeWQYlGYMLsuh//eqljtJ32U12bIG
b/Cr572Hp/E0PoLnPc37+boo8VgmRUztk7OMFslArsAc/nRcp9SRJsG97JO+Ctft
Ch8AX9nmHN4poDHxgXP1Xx0Mcl4doyBpEGmwmE1tDLZRvjHfJiRKPxSNjye+vSmv
NMUtF0fZDFlGQEcjihcaUZSz5mL1jhYToZv4nKl115nevKn5c/+d3JqognGtzj2U
5U8hJ7D1bnbeiVrBepPG/4zM6rdCmTc++/IxWhCevMLsXSpH8tlSWkksgfAfApzk
jjNoklV0SYQ/bVElWUyslhNQlIdIQaNhDSyb5sgoS7uBWiofHebNSbZhWrANDZLb
ome5rWEy/X2XIZFf3SBEgmBwFQ6sxWouhNJZCn95VOsA8VPPoW4h1Fiz2fXEoYT+
uIN4zot3eQ4Vr0bUnxfFjStwU4WQGZckrq+GGyWSt0ojy8aT++clCFMiy/yeOKGe
6NeV6IT7lcGybETynYkFicBAp2ebbcb4zAbbwiTFN7tYZz7gQm7+GmD5cgFrrYac
P9m5lReRp6QJleUqR+IVuGbfVtoeqejkrtd+2jM4EBs2oYkvK/iTUF8Jb9iY9KDI
SSKU5spcb00y500epITCvSKio/AYCtFKJIjBi9v6aIYmbSkXjdtGf5DAsc+0Qafg
iHX098mTd42o4pUOyeuAZfUAdTVCgfPHWiQNs1s11ImN+lbRejHXy7xjKPmZyIbZ
wjiZ0ztfxYd/5aVOXpV1BhrSOyOZsv54PYtrDtPE4X0P0PfMyo9t9VN398VPeLSm
OgcVvLwQuYba0keFvlpSbjitI1977dn5l8ZI+sWSwIm9NoRipkakLGVgLjBw/ABK
UpLG04KXKw/RD6j8qiAaVH8o29+3z4ydWxoI0T4DR+ZxOcjzC+wUd4YZ2/0Aco/X
bfzOyTZe2pT7neXvE0RAHhX30bTDCikwjBruTzYZn1kQrDlPnbAyFzORQWh9DIhZ
gz2pbZiUUxIYSKfuDKHDH4fDjnjqTj8urWjisrYp5guzgoVuauZZrIxyBLQIBQE+
JBsm5ROkVAn154pK02A26Jl4Nbl+IUIirchGoJVm7LNcop9MMHFdZGhy7h8hn7d2
YMFVNxN/thThLs6aJqlaGHfF3P3kR5R18i3qRdaJy2dTJDeA/2ZyGizD7JzkEA1D
fLuqdFnGaH+ET9k7XStoKdLRLIZJjVVlZRVI0OdE2NzNtm/g2ku8qUFqnZx2zsLN
C6c0utsB/hxXSf1XR+wDgXwYyeCYxNiOw4liFsqRPR3jRKbCCYu1R9Z3LcRQ84fS
WNHkB3xt1TS899CCUxoQz5KfoV/hSwQqtRbJ/Zcm0G+ADbP408VQ5Jhgsapm1WWj
kBfoZcdKCjeDZVk2r+PEWTeDfJ3sROcKjI1R0NAoopMlo2Pz+bsily3FBSyxSD5e
pukvWVB2UTBuZtGbEgqV2t8GIlSTXwDP4yrrn4yRmx8BOIfbYKl9Vnm7tasw7Xyy
RTXYl5xsOBhDbvsow2V2Wbw0VyZd4A/8WMmEdDa/DTeX3gPTGtYZzz2fPIcwVVqk
PnxTqwjdRb30cTsofey7ncgqXr1l+rlfS1/f4hUHMFqnY6lo4cDcW2/Z6xuGiycL
UMSuUt6w4WFBxAiwWtchbahdlDii47n/aVr6cnxFypMYngZOIvJpK/p1mY2DqnKZ
YvJF3cyHnxXkEeuhZW21c8f4VS5IWVdlzhS10+WRKnK4sc1tKQIwaw8q0jdOMZA9
LlMsQef+p3gDtEPWiPhUhhgxg9CxnQiOUNQ/edSgVorF4vYEirvk2SRBBVdG/0qT
tycdSfMfl1sPlk7UAJn1nz1y4xdJJR7pbUDyLEaq0OBg1BfqJ0jk2idHQ7MFfYFm
b2JH4ndwMeeUuw+D6yS/6KkX8w7Hq4oktM1KiwtNodogQCqQ0xtLuMnqDgPzyvHM
GtfYk0XopkgjCAoZT35DQj0z3ziwKmNc72Vco7UV4As5sCKK1lIKUHP1G3dW2kPV
viWJZ1BjfXgwuo475wBBHjmaN1t+6IAvy0sjBBcVvdOPJfWJuePqdfjadnTKl4O6
gVOq3QFgqgdvHdgRVB44jFwEwJbNQB6mTISQQYm1kqmLVlygySOlQi6qgKoiIf0k
EZMRKyg/Guh9/wnrc4IpcZt2cqc0Qwrd5z1ikvK/6YoNTaIZ8wtraGpym5l/JcpE
+Wlkt52+qB6b7r2d9fCs131fT6Hat+P0YVeMncW1Pve+YjPs1Vz6qpPvdhOWNj2d
O7DHOZS6Xi3nor6Jef4KvYG4VTd3jRbwJQd9MFcuOkGsFfH+mzxG4Wefgdmy8MI1
UIMJ7vALRQkk4PK2nofmwBc36y82Q4GRQ4ESgkUOWoQ9ZTn0eCshmYIgCTKuaARs
mq/YEqDSNPGXGxi8M9E9ACiw+xRZOvYQj51M0yuXp7It5o8bfxUth6Ki+zcb2KW0
PH9VI/kxQMGBXh7gNaGB6PZBUk0RZ5kCRiED6dSAcTC8Xolv0kqN2I200EWgtZhM
Uq9ikd4gRJvwrkE4eEjfHtxOVZ8XRPHRqkfwZF5fGQrm4cRXO+szn2pIh678HuBD
bSPtvaEG2USNNIeOP21d2H0+/vyaMl1/trdnK0Re81JnGFpeU0pIwHqu+5SN/xpt
iwTOV+i+ovsP7fir8xIb70K5v2czA5yNhZDCt8IzbEAMDlpcVyu6/rbm3Z2L7y2R
VFqbs5bRC+M0qizPM4YpmrDDrotBkjxvT1i1pklDkVjzJBAu3rQbiDsx0W7yIAWj
UkKL1e4m2wgcsC0g/57tjPhCcchHve4m6Bs8YXSIQT/TImEzqmD/YnmR2YDhw/tu
V+sweP2bj/EizsF+3e7lD1OCSSNiGj0tgFnkfS8UGzmqal2i6yuX6FlneRy/U9Sr
LJuf6YQEvQYDVe1CF0LlpuTZ48+Oug6iLclj609ZldfQCJJIqYFPiJye342LkpEK
mGidnyILr7/oQdq6WsZBfsF/z3v6ZPD5WsrOF4N7W4J/RyXW+N5fhH/j3gK5kknW
HcFX6FPFwuryObemzdvSPTsBs+lOlCrGu8Et6EoOEkTJE71k7qrVR7/SIYNQ5n8s
XGccFpPDkMwIyyRDyD/l3Ck3e0oMvpHkcn5JYD1qmZ5nqbIgC2/6oKolsFBfLWOQ
kZ2dz9aub1CoVgPeV8xmgiQIN5YjeBrjL90vEIIDF1ttyR7kWm2m4lIYLVWSqtaB
glHcBjtRSVP31Zqgn6Lf4x+wSAv4AExRnXFngPy+/LWkY+59nxazjZp/cMBc5cDP
18zdv+PV7sJejFuxiklWBqn+eala+eDmBFq++Zs/cP4+qofCI+pECed92FNYcxJ0
fuJXWvlJozk/d53yD+N82vJza1JFtdBVcRAkiQsvUdR096ArXdnWseSoqlE7Y/wB
kvsjA3goL2vbC+VaQegrLxu/rhgij8NcbTbYIPF77HR0SnceBLYsZsbdHfaMpdbl
AcgcwoNEGUz3qDTh8fjrK25vXPenXSfx4Ehve26Dsml9h/pwQ6Io20l9mnBF1Acb
ZBtemAYLcP9Mfsd5V9lnRGApeo1UTEduea39gno7Vu/PE2EK2q6CBdk04K16j+k6
t6B6G07DEdVzGCvYjF+eI56mpAdgdurienBKBpLa6VC+Uuicf1xNWjYmvu6AMU5o
Cs7cSuxwRvHaSOIOiOjlqff5BMafHTQWXTMcnQwZ3WzYXqmQgZUyEb4CNSM/Qdl+
6vgEy5pWUcJu8d6FRRri8sz8g8pCBIGd9aszmV2hKuds6lSQFfxlmenk7xEO6bYH
oLSnapxYMu/KawUjNAz+SYI3iFxxo9Qfommj2GpaYcjpq7Zn5nAFwXXqHLqB5RiX
byz2MWwzNxJ4Ug0npK/2gibfPEyPayXhe5z0R1SbLpHZ4oj3UFvtVigGyeaMYRmO
IEm9z+MgNHKOdUnqlDW8PVUfCN+NdZkkQbef62eVXjdS+2NYWI4H0MMnXI5SalSw
ZGbZVuR05NqmmmPmz/izDQWqZC6vVPDZwZy2HUbn4BHR15MJNLj4ATR8VBem2RyJ
Rq6Oc3jMo6UkV2+cQzRhBJw+o0kQo8I3MnoNHgCdWrLx+enX7axXOBOk4jufgEyR
l92/ztqO0PwhnhGMwTXT8pJdi82oZ6M7zff0kJU7J3nnjwrkVGeFNGtgrLX1RDGv
AC9CfmyOTJGqwt6p66wUGupDiNbFZNJFDNFHuqUh5hLOlANosNiRdnLG6lnave94
HRGxbF+V9lI8cQ644RZwC8ApkJ+6rBnlXOmYpTiNwK5ou5BtNPnSIrfTXRa6f4zB
vQvWlaDiz2yDE1BHnL4GbQtG1KBrln1pKfRxtXGAi9kGBY3N1omAUia7POXGvOHP
ZHIZRg+fZlickTU5FDJe9Bpr6/PVzI4HKA72bUQptdBdI5Pj8bzV5UADUgHlO1ug
3FpewJxgsT6lUx36ePNcuPHdp9udGW6F+7Y7Z5XZsRODu2WSVFnuMauIqbO146ZR
FTIcDPzYWRlzmZJKZ/ReNc3ELj5miwqeKMCQ1EYK+jsW4cfjvjS4Ng0arpnAlTER
zk2UhocH0kL7kNh+YBaGpNeXEdC2c6UXPTzgCk6X0n0BKQiE9hiUXJ4sTXFXGU4Z
P/Z6kO8X63c87vzj2yuGL/wNZ2vAnheXBIYcuogK4aPeawo61NXQe0NxMmncwiq2
jcTuXXr5VPYiOw3vFN6Ut6pDdMy5jv3y7+OqayoJts4EwQcH83/YOf2SfYQ7ZveK
aWEYjTk8CSUQ2Wb3EfaDo4PbhSmh8dDshLosKQxelVe3bZsqkgtScJiVBjLVc5me
1ce+3g2EosgyJ28aouV6n9Cz40+lnbDxj0o9YJ9IKXW68huX6be0gBtu3IPkeRyK
rPLvoyoSbsUr4c7o9JLB0oLEgPSmNFdVI8i1lQa+p3HIhvp5Dos0xHn303RsRoyp
w1wv4MeJjeN0kd0tZqaIX8+dy2xa5AAoSahY8ztWlZ+HQSvFID2d9VqJmOjv3cKh
6/ycRigO4SRePNkzu5qKvLxyLBE4aRCUfWYIzUvCIo1JGMeyuefuCXwksq32a5UO
ZYOhE7veouOBm4l2qJ3vV95uGVlZsUhe74AftfVO5ubVHZWaDBTdBvL6TTAg2iCU
qskEEKQLfL//VG+oInwHPB1R24k+nPnpvCMRsXLu2clLoRZOjEHp59nvpNWMRG4v
UH+rIzFtaNN/FFSrQmY0KNyoUyD0pBdSFG7CLcvQDdWsHh8U6HynOMsidWqnsO96
bjfzYMG0H0JZRl8xY0DAWUR1c9R9f3ocdgrhPLAY+f+IVm7MfG5fCKIY+3GFb0cl
7LoD97GZKNtiUeJ/Fk3nNUSITZjMksI1/oivsz2tK1KTnZsbLmAeG4eMk2uEdFq7
MwidBM9Vln1HYEVCzsIJCLcxovcY4BDbYeh1DXmMAT783DhCq9WJa4+IxrbYxgU8
GN6FMjhOsROx5HKnHyRKaUd+2/nK0mP+ZS/nJNNwpZL3F/j8qRnGies/Y64+F4I5
dCcBxdHaCPLxjG5/baNbtQkBAtk2jg7EL0+vlnkZyqWp4Gqi1BeFBmVHEurFk6/w
vjwadAhwU5d3SwU4IAA86qgXwbqp3p5F2kNhwJdM2oFyOluZNXhqN5R4oKpJifhj
FNvJok7ZiL6G/zBHKI0Q0dSKf6sg5FvRA29Cj5hbqVmz4vl2bo7eIoV6W7ZX1jT8
GiY1e9Dj81tbICtqTPwLTzuc9Uii05xOp4TDqMjtBaVucK+et4IJkqkBsJ/eT9kH
Tl/zeKN68gcm9zUoiReVEbjGlEkeuPtvq3Uy/tqvXjeE5OkzfckhMUt286wiiHPZ
uZyk3kfGTeDEzbJeUtSwJadGt1sHSpWGFY+/BR09iMAfmzrRM/DpDA+W9n4TqIh9
JP9nJWqLfyAnnQRY+DYdlKYnWJR9HFJN4GUvL0gUIM335K50czwOIKYWqFiEQc4s
plSA6L4X8jYpJJpzfn03q2Kom/ypJvNPnlp19p5QwERx6E6Hf0JAsHAWKkJYpJlg
r5hdfX6KqtZM1ZdGNq7OtOh/ZWS6XI7vtObiHoIsN8p+U3lYBuiRAt7IKyO+CsNG
Gw90BCElWBUzWYXWI4MaULy4BLsxwcud6kAGKOe4t0P2pFw9NVAQwJ3DblfNZXlG
LZKOG8CfwmGB4ahFzNJOBWYk0XI9lnj3CzFxNHL0G0ygU/0kWVBLSZsVuaYbeIf+
Grcwj8uC3sBmEwETUDxNWyBblpNFxzQ4zO8C+PTbrJYpiLiMBrONY7kmb2YbhHBS
8V4/rwsO3m2I7fpJFvweZ49jPjU19FDTvPrNWQuthWYBL0cdBc0CzfPD7qRgQmMk
i5mdFGrf6Wsj+JGSGV74lVQiuC7eygWTx9Mlmh2RoUtYtoy5c8lfj9n1w6Xy57QF
KwhTrKfTo+2LarwDIPzRqCfPvlK+KmTgyKie4XAgjcX7KMQRNgghqpyZbWeVhQoX
CuH5q+2sDIRw9b8OGGsFvQJSibGBkfCk3INMZKlfvkI9VA+UGQIDVQXSaoetC28J
QLpUkUA+mahFvGiBs88rxym9s12mYFa/kHs0uzyB4o/ohQp/2i2hE57as4RPyMlf
NELmrTFradSFW0tk2NtgeDPBJDMkiQKg1ioeEhVBWULXSFRfAuSnbd/zWmADee6y
bBKq8alzCkku1jKfhCbGT+zgV0OfDDRgaT2NWl6Z35K1NN143Jws7KnDdpqJkq2w
/cHjUruknsshXgN45lV3BVIFSdy8lzZCwESKDJHhcJ1mdQgXf30u3Joo24kNXfa7
YiHac4GHzl43Ld2+A7D/HbkaJWHmlfKhfUGNoXdErpXajLObL2bVNuglPVF1Y6iW
msujCTl/MSmGEj4f1SZlvq/0gi44Tb6GqZL2CQchzPj4+wcRVahgw1LRP3j1K5Uo
AnrsaD3vscskQC+97XzkK26af54WVhW6yjKrQzR4JxWHIrcoz+qPaS6ijY6TSOyX
mb/bEBryRkuRRsbq092Orxg2bsOHYjnuvMNITfEuKUzgs396ivq+Q0s2IttTd+Yq
dtywYR1e7W+zTY6E6jHP1rBktug22H2hLSaFrTDFPhB3oEEmksLB5B/nx/wptwu4
oPCsW37aqQJvzKGfhcMhsYb5oKmjbpYbQBSuMlo4JTYAA8gkzGC95TTjZoNBZyAk
xEWWZsAPXbj9Me+9zlVjjS/2Z0pJlWsrSSs9KsmUY/H32cLPnQr9dXVTrcRk3lgQ
FJ4xv9Y5vBB6C3o522WWwbKC/AOua9z5bdwodW1+A2ri1+O48M7+DkeC82Zxa06g
176k+G7DKLfbRNXTMkTJeTDj14uP3gTzINOPeL4yw918BqQ+NMyQH7cKfyce/pGV
u4p0grFJFXeqyPxMIP2tHjUq15EaySN3CrQOsoJPR7JQIomPVFFucucvSyR/c0pd
Z6QbfWQFdw1ti9h+pt9QCRTkF5GGOjv0no2jVPzVXIlPfFj23IQl9uc4GCGIq9u8
OnAySGPDdqKG2sY/jkbSRe2obzdK+7rvXiveo3wjzndO5yiJiGT4mRWk5HcJK6ia
xD2fhYyPJCoH+nlLLx2Op9nj+bZXC35aIeijI8AT4vwUw8s56JRMq0eIHiv/DxJt
uDGafxICvDff56xUk9BqjBMq1u6vbV/s5HXPQzimQx/61bw+jkFocgTALuV+J0BX
PnKpUL7+dnZUeehGZyCRGa452FVTi9eB5wlxv1uzhHZgmdiSp/0jdrWyo6MIgj0i
5wvqdQDRXgfFC/GdXplEX4NEmh8GMwtCKFDQBrsg2e3cbA+hKsQpnTiSgrGPnF5F
Qnk9sDNBVWFSB3UN0rP1iQNF76YF7F3SV7t4HqJ07mcecJ/Hg5uOsRQk+ml4zRMS
PJQui/1vSCMeNyj9eHbQsmE7TgUDJrHU2EYchULzndkewWtmqORIL9SvyeCe7cfa
PR9SPVyyyzbWJ2eh1kN8WOSZYxW7yQ3BoW3yF7KlEr9rUkyTJPiJnhNNIKjnogAb
Xj7I44ODjg4EwXzRJIWMtx0XOAh5yODQsUkoqHhvza+T0FgdXcRARelN3DdMx2Ja
2Bt37W/J3/WBlBc/XnHYjHYfbkcDvr2TagqnW/5o5u7C+k1HWhsuVOv90j9iROkS
liVD1nnLg7zO63DxwfTPbTl5C0xzmt6xbcj4lIQWb7q4sV8cwB5cnJotoF1b6yxB
LgsKnmtrqnjA3SuzYObN+dpn9MgvisamPc6Cfvtg+z1SAWjraDtrJMSZr6p1+J3J
n5cvOYF8DJTwc0aw+a1IA/xmJRrDYhJx2aF++apvZTUloTbUWLBQZxyizjMxnmWN
UvJ1/ay1XKQDEtIxfdnhsTmzi2GjD1oC7sCgNYr7i7Tj+YFlDIT5897HhiBKq+sN
H32NGT1WgHvhG4RlqlYy/wQHnpQCS3weo1o8fV7wQcX6kwi0sKG6YLbBJoG4cscO
yD8ZfB2a9E5WR2EtgxHtp24vBGLdNiY4eKpN4D4s2fwTd5c0/SNGF8kfMrp4sh44
tY8nDI31LeC8P2LlbGC98+DAu3jiReoIwj1XoR8C0qv2OtVMmx3vKSLkBWEsziHp
Uzq3AxdQb+sj/snFmecCz0wdoviUixOdDYi0MBBpIAmqcDdkQMGfo/8pyGAzBw/9
XJ2WEL4gG3xluzwsYzqlUEwYfGR6b9HEpX4rN9WQwQYEcwMG3NvONtvyCKa4llch
f/h1+X7QJ2R6HVDWg6FPOxPv3XO0Eg5oJP2kfw7xq7SDEzWXiTcL7pocK6J4QJTd
1ZcHFGjHZroL5kSqd4+3GhdLu/rqNWn6REbDpe9tu4+1lu6/BO33FJNTQeTTFsV4
OcdXfFO8Yu5qKiLvKguJHXjIsiwx8Qy21sEZZ4PGGzzDQ48NVCs8TFZWBJ9RK+sV
maTs3SCHoS0C1ez+BfEjR1+4WcYsZ8pZOY62i+IqYPET1J7qSaVUfI2T46TlesUb
P9qL+bV02IGfgpE+zrDOTMpv4s4Jz0aqrpg5c3xFrKebd9E6mTlk94CaWEJLc7tP
YGT7+qs/3rHd4lTIyrhZ7NMj/i72pqjxdT44KLk3CGo8Lu4CcBSyzPdwPpnYvMYo
VS0rhq4yAh2N8eAdQmRmFKbMzdcm0W84J0tAz+8ONaTQ9eYnq/OFJAOP9cePa3/G
P6J5Xhz2++5dtjELr84JWqbvGRTsHjes9zGNNxbl9io3iAYFLGfkG6spwUV5KD4R
BvgckitgDGNiY0660i1oYU2dbGyhdiW1UyF/Ni7bawbaxUXEDjTDoKimvU80qUD6
H3LBLUDn0w/y5RnTKhw89Lva8HY4WsSm9Fh96eAoNI5Q10UunVBQDbsq+VGfUSHi
36mM605VjE60/AOIODbbBkIMBDpc0CdDMT7x/nOzLkmiUOx1bKKxVXWfF4GTgpuJ
gYXWUz6gTaYrn7xQFnOR/LqXpZpTfU8RahJhZ1BKaH+R1d+ihu5nGU0QobRXJs7r
s7n50ZGIotj40mAcyso0PHkKY1IajTx6gIIcitnJmRmW9tqbPMleP7t9DF4Yw867
wHAU1nz9xrCXn+enR20Wg+KOR1d9TmGzym/d8hjsT2IUDHP+lBUhBim3rYbhMp2n
vwesPqKlYXjWWbksD2NU0+NC4fduT/VDUcjAl9IqkieOwKKjqVQdDXxAoFAdcm1g
VJoJ1m51LgX+CD1xpVuHf2Wt+VbLgNgPAy7IlWiQkwDbNdHgzgp2eTWyPpV5adM7
CVYVmCeLuAwWlF/wxKMLwSkWOEqdZ66Q3uMv2T61ySIrctwg4FphCrkDEIf+IMuw
mv+adxLl7QXn8poH9TtYhe4h9+kSPqou3NnlHbOmnnKy3670xYUn15KmPUWTWbbc
gHRn8Jju8WwgoevJx9Mdw5Jt4W2/o+VIcrT4Ahtltiu/ThMAkxaWiEvR5p2MhcBY
coOemdi3zvvhNtdzJoAh6qkOEYTwVX0MZXlDFn7WGwDQzljf/0OHKTccBxYW5u+s
eUUGOJbNsD7mqqPNwpk0ETtmfbUpsNaKEj4TTeOc4klGTlA83PBz6n+sADwe0/yh
umdvaiLCffyzA81IDJX6sGTR8jL1q6muF/cw2HXUOtHA01DmePyOqw2SykiYiHts
pOgBiDF57jlCaGJhwGTZW1MTtgqL/WASACUikt/b3duIb9RD90K88QZoq+oC8pVC
FXQiAJSANgqhpDl7W3L4frbPLAwrcBb+hc4yXc4jhIEb/5g1IQfr/zSina1tTLOt
SLo8/7uG/Z8tJrsK0gF322CkAI9XXNIQjcwZOvOiLcPc2bzhEe0sqc4wc98oqqMA
gczUhowVUz/+go8SOwZ8hG9nAzuOfgurW8jVmmKcrnDiNoLIKT2sGO54hDhLi1Dd
BIukvhlLOyAAX5UKSwb5+ZVUhY3NEHyk+77gGN0/xxGYpDVF6tRG1DzcngW5FNiU
sPAatOrqBCtt6mwtsOEMPARH0YcF1CXSJifD/Pu70OzM3D/v2HmdHpSuOUjTDkpT
ll+AVGl+lYMGD6wGlfjogoGf+MPPy4vmwCG2ZUT7JB6V2g3/y4M2vX6Ne9LafBFb
UimRvbUcDplexxK7uEXdXa9PPA3cdyP1EuPGqMYChzmnWcqJq96qmdMat60SSVaT
JRB+d7oO/tqD2w6zenWY4tpHg8kFf9ZscX5z6u+7FK3w9Jx310pDM3JeF7fWzLrh
8l6eySW2iFWAYo6aLq7P2PzAyCXTylGC3lMSSAkxB0DZFXj0FoNv9XH9Dts1/Ls7
7pyDDYwDI3Zco5bMOi5DtCJz2+6Y1Et4r5yZrHTjdm8PK+10z1vt4xQBb1/rOQX9
hnRsvg9w14DKmHEdvCIAX0zvjeWVBEsvr9DZ3y2Z6MWElFcenAF6ubfYCYt5Hhfd
7dzSLhhRYHWBrfHpJWfTnRQGDIY/QwIdHbfeVgPZjBqAcZmcqbvJJx2aVGNO0Ig0
5lYMo7yP+yIh1YOaZIDj2DiyN0r/Yu+HOoL7UUzapXZwxeM1T4QUaXnQF+i7D0Mx
BJapG/mMc3Lz91xNlOHyleleZ7EKQCSBa0SzgKnHS1NpLa6lcuF6CIUgJfDnnsFw
NM8gu0F1jqDI0/2Otw2nOH2JVazufDWSH6xsa66CgWQBCKbPND/8s+aatOFF237c
VvC42SF6Ii2VoWppJmXEeVW0ufXzfC1kYxihO1/6ruJZhcgVHyxPlJgpBIhI5K7J
DcWRf8iirMSwn04/AdMsMj2399b9p2+qgrUi6RV/u3W5bwklvS2c6ZkTnl7zYR40
TnN58w3dqg1nu+PdK2VSN407OLvzn+JxWrXCgnDRlsoT1XB7T104dRKXQoFovi4T
Jk3MlLj3zDJttMI4bC5zqjNPNkfr8kyOCoHn80TDLz6p60I6mSmCs4nvFUJsLFK+
Dx7cAGNSOXGmzJaOknsHt1aEj13ua33Uj4gE4wSNW7kq4W5LdW4tu8R708UWi51t
nWKyBhm6kIYibQihN1872+iIOcRM4TEsPxVVMh2eg8bZLKL7uNKAR5x6M09+AVnr
eK7V0TuOTE6KriuIjJEAxbneygWYt7bXnllFotU0/RGMLFnmjz2eC7k78pSjMeQv
RSOnddNhrMNfTtrgPL18mH3UamqRtdO7IX6f4q8MNKsPOwY9XyiWh9+wPHldpXTX
hPm1A3Wce2/voB6Nun2ws8Sj/25UoTNvXUi6PdzNSYgSUZSQa5rkMGqR3aBMbzKn
+Y91UksAVkwSqEJpDdrqrdesGx5jgmtE8Cj5BM+bnMhR9scOCwjKGJA2830fSvXz
`pragma protect end_protected
