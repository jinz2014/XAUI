// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
psXPVgXzKxuOr5PR6fe21EeBy2/JH+xsF6PEgfzVlh9xLBfX6/PZjN/GXy+rBU+b
A44ygn8qJcmRNkdDOuXxQxBm/5FVyM+7BjYux/3JD92cLDiJZQGIihrNSnHVBAWm
DX8fWV9Drn9BKDVv3hBuDb0QfgZNBmFkVgTWmjSnJzw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8592)
Oh78XeeHGUBnONOK2hKgOhjHkoONX8siy5TlHKI6NvLJ8eMa7OsoMS+PqzcXWeFb
0OYGIMYft83qLo7slS+0CigOVmrtPJ3e5TQKWi9z3vidN9+QliDNcmlOBvK0JPLq
cBJ6E3f5LPZeN4NhgVJIEMphJzzGDqg4w3Sl2kDtadBMlPnlS0Abz4A9iHW12l41
6r2jtau2ehSIX2HFbYL5fMQjNVmIeZIPBt0bC3hb6pgwh/KZKkNWtKD8GgNOFw3U
L3hRDQyCVdPDgGsVoUZuGc1Gp0UuV2vxhcnEsCYXz66YOBZjnniFGFlk1bDmn3XS
s0TleT7HmnT+uB8H0mrq3qT5Ysqzd5Ill6LprblBRwtIFv1pKFJiHNeGmBB9rQ7a
LjuA6Kn2QGF1o2l15vYCjX/Vlwh4lBeHfVzdq2EhSf2UAztZv4ncP+XUIWLjdXQE
K5l2HbXZHkhhueVD2no7dir+6a0BixM1PDit5UsG1SZB7RhKVkaZLlOMOJiCM0BI
uvY6eqpvWm8CqgGVLaizYODNNP+pcif+3wwMOBgL6XdUw6OilRRsR0q91wTYSTok
oOMDRFzwG+dDqoN+48Qnvb4ZfZYYeMeNEhDxMwZI7no+oboHuKw9ZzpOVnrHWtew
2aJ+iUcmAGlSpx4j9VJqkyxkK9rEPieWhJzdGdnyc0Z5sfXIhAblUYuKvGhXjf40
V5JxDoKeUxEEvpKoc1MwJMPGuGQ/k+WTTL6oCWV30/8e2Lsf7Y4ov4ShyW8xd8Tw
bBBTILb/dDNePDn1SjYep0I+04bR8UxuP+YTMSM16N1lEiIuCD71pcL2MnW/0IRg
MhqxHOShGVDiEGg1bAnfE2alB4r9ZcmPcLkn6N33HHevVkMw9bbHBUD+bdvFqKSq
lYDUfjL5iDXXUL/re2atRRpT9Vha0jnXusZaydBGvt/ZPin9DjeJ3pqPfd8HpSyR
2XkuxZq2KllFkh3Km7bUOw0nowVoFpK19qF+DQpKoMEDLFTWs/C0NjymJO0hvzd1
sw3zJCay+G8YRu4K1ybjht3LhiAdcbx0uPwMluHq2xP2mMFLNmVNNF6JtRxUCfkQ
wAV6cYcDK7SMYS6r5Jn7Puy/NF3rQzqPc/1ao/1HhhhoZ8ju3XiCk42w1ORjTnP6
7N9LgbmFdk6hkWXVPgCYnC5A3TvHbECrIrF7qwCz/6hjYpcuxOfgV1o9/x2TzBcD
r9h+QhaYZGEpkp7y1oMhnkg5FniYWcmJMb8NQP269ulKModce1dcW3UXWsQJN92A
VztdCqX9Gp8CyFENlWCGBQqGrF4FgRiWy64j1KTFcChOfnbjgh8Exsinb9D3Cfcv
MFa6mOntX+4qUQUM95r+yP9ES0bZ5JWTBBoGajQ10aO60A2fCnJNFBknreNbvsGV
Q8kQzlVbnUIBBSkSYVF/C0SBzxZnr9JNDsinMF+BAJKRqAlsao1DNqwcrkPejOZm
Zwen3nAwnWdGPMybKudMj/U/Z4kTAg8hzdxHB/Z48XJH9CwB/3imhBoAxo1wjEQG
xTvOaQg0CSUIDo29FxBOc5dfcQEup3LvIBsaCYriQek40xBaBZgN7eMNAKH4CNzz
OKvNECyIC9BqnxTGp4vpTH25AW8dBMFzVyr1mjrLlNCxRd5Ju+4lRwjR+cjCgaQi
FhKtsdrBlJd1+BQvKAslupOGC/GuOOlHJZ2/PFPSlFvY1tz223cm+THJEJfOSgV1
bRddNjWRSGU4x5Bp4q6xTS3oUflo6QHYcz1i7mEBfaeBTJ1nVPfP0hQUobkzeumi
oCbUrrwk01IMbuk6iWvQix7KXToFLv5qT5v4Up+HgrVpn0MZUYtzyqdI8tyjE9Si
rG+rHCnjuyeHNDNG4Axz2yq5IOGga7lpzf5xsrSyipnhOdNxDrL7Gq4q0adJUz/e
49CSh3WKYw0BugV2Fmk159dZd9iNKKwZ9GH5WCsfQtdCV65VjhY4SNQROkYSBltm
wcHyf0klczXugEHDW2XhOHfqyzDdSgYaMcZfayZOMeHfzm4RM+5G/L3Q4YsoneOq
fUam1UBcJvkkH5cGTCuyYnr1mAc1/JJAG83r83iM8s1oNn03Io3rQrJvKZvMt28S
EON31taGRIOhmkLAy2x1OvVaiTQcfU6/msIImkCia2sZvrTbELIU/Q9ZgEoXDsLn
9yi5F0Znk0SILOMANkdeT+FbICk7aryokOh5k7ZmhiLBx047qwnCNP6NqFZKLRPn
L2iz/vci6pI2Ho/59L+IRXe1Pet5C85o/oUYNLIppqypWP6yBXKVSQyNbCdZVg3H
Jnk6+gWjwQ9IhWDgskxvbFe7pookwFeWfwbXdbH1LVSRdT40pAL/MWrPZiaejXu0
DJPSSIUP/wXE/MJy1IrSsfHAI10GyZ/qA0/642XaJ+pQOycXdLUu7K85lHl30c1i
7TfOgvbOYFUFChUQo0EE6NH0BOUK2V8PScG0mLGxYe4r6Z90zQZNeuH8Y39+eZ/g
ok5tbsecNZ7+HmSQZEF+ys3txV5KNzpOMwNILvaRftxCRxnFpGBD2pJoz5SpkCJV
jGgEiwYvi1K3gfDSnf58uNIaqeVr68aTIvR72eMB/Zvhcr94CpxPqXGm2cMHSxzW
A43TGOeoIEiqnj48LYSf4YPfcP1YV4aXkxcQyXrsXOx29s+6jDfQKaHsgd+hFh/w
h003DA38lhfB+GmFNUSy5l6TcMe4bLv2mIuEsXWfjwJmrR2yfekKmwNI+CqZsO4M
1FccDFl8isD3hJRF4alFv5sj5i5WkG11KHcwf695zTOwC/dj+WtZqrTjhTKZ5cUU
AHc3G5UuofzF/frw0sGuYze+i8AFBB8spxIAqSy+oUyOjLfhHYZk/LdSoj6XoIaU
PoNjiKn7GUbUSPRHHhTrqKBmVVTMyj0DuMmZlj+rTUHATzEdc9sVixyHc63njKyN
yXKtMrVqhgop+f3c+BlTUO9C4D93MQNhtsX71zeDRxXRvdEiVdyN0MxTg621XqvV
tZUkv5dHkeSb/hEBIBD424i/Bs5LOTv8yTeCLIyNDsg/4XVWQERcnPLqL/iVnFqg
+l87AJgPhJgJw7eTIHsQz6wxa2Csw0vmDfpmbRHWcysh9UPH3C5ExyvItIsmrIsL
0HoO8SPkqvD7fJRx016CKYZOd2yDwf2htx88t2pHYn/D1PebiLVbEGLOfciQYxlF
gwNm1bb5Pcy5N2Xs4lySge4MCn6aimQkNdNhNWEUX0YNgliiUUQHRW5T1IUXNiDK
KIZVQidDhbgnpujQ9oeM6fUtNLGPg8ERE9wyLlAY9Wx9Um+IPrp6PXuaHRKL9vNZ
Gtg66Ubn85VI8fHOrQK7unPEptPBUytw4yZrXeCEKZSkC9/65A6RAlzs1gqkiWHh
nMECTPFef6XJLe5bO36soLVM++5segK7R7JswRv5xLGeentjR6vb74NKJIVRCxXH
he7daAafVoGesJFuaPKF+odT/C4M29+56pZEKOAqQFETdsuc2iwH4HZgY4UOsGZs
hPGWKozsPkAM6UNUcz482kEvYynseQpApRStf3Mjr+mGXqmT3zqUutJYQkCqbEHT
1cNKyQPeSrqWuitxUU9HKJMjon0V7p4On4McwlPOq55IqzAugIIoIEgyRY+B8CX7
W5kxkH6THqEv7zsdc0ssQ1IeZY39XR5HEyvJL+KyJifByQcR6DKaORsxxUkj6Yi1
Xs2N/Ok8ye6K/NgADDKTi8Iie3+62Rrke8IZaqAA4ftABV2DI8ufoNpRqgEwcUeP
cJcoovnA87dh6Egyys1mOg+DAkxeNcoxOnkIKzs2m3N0riIm6KSYqMhk/14/I2f7
8saAIH8AUtHqiK4a6xQGjbRKmUc2xhH/LZ2T1eoa230dPjXw7EwnF4vy/vqnQOLm
RuoaW3Lf3VpQMJmao7ZhPeTHoFfSyvndwWvLHyrFV7iRJNH1MFJ2VR0x4z68ma82
o5OzTde9WJ4PQntIUCRAPLM69jv0ZOSx0khNHlLsBmfSKkc8bnxnrRSWMChCFbSE
NivBRO4p/91i2wwjf89RuIng34wU7DNrZCkpZbqjLTAeRgJDEtP/35+SD3jcIwcw
whXwy8JKD5CQZIsJZIUKpOc3nmS2chGj5BKT3Z77b/p1WqFFUsjEla2OUcQNUN8g
c63pCgn2ZpyGv341p3u/lpw0etySIBfIwUV3gqDo0stwabPKfKyZYG1/BbQjznnd
aRF/Xk596Ix4bBPpcD1aFZiGJrBrj2z/uHXk5TjGE6StOYZWi9TCZegVW9crbdw/
LjcerAZIb20h7MCW01AmbTY+qqvtm6BlFr/TkHM85VzXWXh+ztiRZU5sXnM7nY39
ht96dLMRWexgUxV8RGDFMJl2QiwMhpSwg1iXZIuyx37KjJOxK2oQPgX4eddMLhV4
qkjRSN5vfT53OZ/QpvL4nf3zS/YQucfc/AaFSCKM1jbd/o6eN9TJCT+yl3OTPPYE
NgGpMK/58AzOGASghAiUp7ylGfhHVw3UwIkoj5cSesaPi2tRmPJCdBhJusPiTQaQ
P6Eevp2efa8mRGKJKSgX9KtG43dUecb8cdV14EH2TV6DOx7nJDRdtZg/QeCAXaZI
I7XzonlFwdvEktBHvn/xP5iJuiC+c4WXRk1n2Fi8MTOkgKVYSBpHJuR/D1lrnjR0
2SOSxx8mwH0EKe2rmlYnIiSAJqmyUSWe6T9rNdcKUV0M7Ug61tXR6FQYrDL4zKp2
2gIWnb8V57XuRMHHYOIDKQxt78J8fdQyTzukcVkPwxMIuU+hDmQuzDaPltqCBP1u
n/D5VMI/zHAvrgnY8kKmLWIChznoB4bhZ0Ex8ixGjzU7Jj4E/Ls5rrL4uILem9Sq
BDcVokeSv4uH5V7Ad58bSmpUn24I8tUkr3ifXKcBmj/jo6EZGdSEA2ivjZOdbWAg
GJjypMk5KHGdyrqRowY0FvO6GDmfCCWqsIBttl/TGF4wY3ZNmQfWu4LVGQ0gqPOo
5EHuDNznzczCoH3anFkwvOpXL9fAJ9dXEkw7W9KXxNHJcs75wC0z2j7NzVr/XOvH
7UhUIorCWAO0MOOx6UuhsW8VIokMaMgKFxFCmZ/iIAD6TbA9tG5scmOtIX9l6D8M
2Zbmd4LfMAcIM9RxQlD+yDmVfbayYKTGu68vMfHs23aMkkuKqeSby7PB+bOkR539
0nCAcCaxbuL6NUCQfuQX4StEBGTxVy33/l6lvLYD4Y+WPSa7NHXOq5NDcxHvwTJo
GlikpwXNkhSseuenahUUGvOZG1tEMVTKLIIi0j135m+Gw4KeRm+duKKEAXvnwzTt
r6pIe+efyIWFer7wU5AFylKbcRr5ab81+nu4E91XeMB7TCNUmrEa9ubypTShLNzM
yUpHyjvTTTLk8+JaSO7vwbIdPy7xkCIPw8sxhLLDkynAB/HxgYkKHefQdK2EA6LC
5Xw/oPeK0TCSw4SH3LZukAaa51TKpaARcvb94goKKSEVUuq46emGLfsg1TUbdL+d
Hjwrmjdg3NFTMqz7DxOzC9FeWUfX9PWEendl70uoaRLmG+dS5lpYwetxVVTGTzGH
gPXxiPo3H9uaWM/aVsSiwYKQfkbkl1eJNVcQnznoP4qeRw9z6MDhg8hU3SQ6BYq3
e1qBS7aiVW+HQFDj8NEBbkgKqfX0TTEBuYum3dlkjZejuRu+sSz7gkwy2gjX2CSx
o2IkzG9StX8Huh/VxX0ZGg6wxCSCiYNzJTa3p/D/NDTFcKN6oqnwc7BFKQSrXHYp
LtUnZc7ZAeJbZzPBrEhX+wElLYXzpCJpLvFPeLk4vNDJCgrLCMxTa6n+XihVSLQV
pruUTVYTljE+ozAgrhPNvLJAEOslg+Yzdl+jascTRV0krse9ZW4uU3/HTwbPvttT
wHFkmNHecLrgOsUIdECQ6L0iBPINPp013Fg/sB47/bZlfi63ZBzm6wCMSBBDiQx5
9spK6LAdjB9SM36/gxPVdnayn1dMnj0DcpuKQYEFYodw58N5JyLE4RW2Em6G3ECE
mW/G8HGVocY62BsR9Nci3sXqQ1DHAtk6+ZpXCUmvlz2MajT2AbwKvtVC5IF9BnwX
9AUsSdalX8ICg4repIHw5OP7PW+WjDeKINBeRl4WDPStD+I4pO0cm/G/wted7Jdx
o9dk+ctyu8R5YCxEDmKJ7xxZGio+Mke0zw6bhF8VT6my9D24cg5hNfBJEJ7+3iFC
xKqwj2eBR7CyjIia7JErceB+kLlKn7dK/bYRIkufxOhluRKc2HjIB2oM2oPv0E7U
3y5Zg2Y/ej07h90puAWgHgCku41gKjFsd84prMDzjehMisAv8PSk9vRr8C/Kgmtu
qoc/w7Dn5y0dSBOT5ZdcEU+0bZxnVtajRj8z7Dm8qHnarvVvbKYOxSlZ7SIsfP4p
9ykJCxKtMgnNkT4a2VMLhS39QmcMa8ojporoiKg+MSda879oy4IGFnoAn78Bd6bz
4ZieBVO+m3286+cbGe30xXiYFTmzFWVhHGl7XCt/62C0go/cbcLDqawacCPGmNpq
4W4xk4VHqOXgnxepSnYu9Ydad1D8Ebo4DH3PAoCq+y3o6wIGqWXRfmgkIVcrDVxU
tNwaEFG4JQt0bqZvnqrqskoKNzTDfDJpg9wYxR6fiCVUE6Szr0lRXHD8uNYYfr/n
uOc3QQyOc+Q59/zQhSR1O/xDGmPMDO0Un274yhn8yVchhfbTJFV4MNAy4zAZvCzr
Q4QhXrMmoZlj1D9QZv3gtk/4M6+oYbPne1CEm1UNH0L7LAGZtskVtNdFlFWm5dZt
YuqHKIwvs01eNakWem8K71xcVPPXR3Sx6axEfxYX+YcuicSBCi/ToZCm2DxcQFrc
YRAj0S6iEOr1ubdSej6lVdeCxLvZafsx+E/KU0yD54NkzgLrK/uwadWGHBPrqQaq
Kmo5y7y8H2yAHVhY5wEqaUSodNDt2TtgwiajO+HmlICU1Qm0JTke4maIXL2nso/o
Jzcw1pzoYbHN+R2p9vMslhDz/9uzwOHeRX6dPAMOHMZ5cij5SBNWeikQ1NixDu1M
eKQjMbXV/lYqLwQ2pZkqpibYYJQWq9F2KZGOXxI+Lm+xGaqaFOksdxfkrM3O8/OZ
m5XnzirYeTKLEeEHOhQHsR/JPOW6sfrtuTxMZXlgcpauly1H2scHpf3UPgzxL2eY
LraCNTTG8Cob+wm6PeksotZuwSNlej8iFv3y5M4IaINsV54TyEdGgBW5M4pfLB2J
DbChSUqWKO/r27LQSelZ6Mt+PKLyjwSVEUJwwb0CyHcr+f5a3dju3g9O/3Fikey0
SMPFKHlX32N+/Dd0sSFjqceeDZo2UM7pUnX79+bwvKmIEPztK00PaWL2qVNl1OZB
hDbEllj7kzRLMp3dhHtkwYZkrry+Pf8VhcrXFwwAzvdU3jedD8gLDqvjjBHDkj+1
M7L9HXsz6MVphlGUaonwrPzeNzN57H6NaZnmOcRW/zvB6gJWDAxZOp3nDMQ0CUug
H2NE/ksyVoD5VM5CWdgmzelVLXej3HY+Ni6qayw2aBUhGVuO1GUTrrXPQUcFkvbm
78mNjVGGYVo4XNN5WSnqes2fxqFYLB1Qm1J0RFNJwhKhdeFCNDoIKVwkdxDJihho
Rcu8UCRM1yVBggfrgPdOIZIMnaGhX8eQmNfCjq5nTeaS+S9OHuL+btDrlklTeGuG
NKbkau5UAvDvhViawNXlS3xKa1K/Cy1wWN0I4jBB/89iJkUU2VVfPCl+8qb9gf1V
6+L6SIkdXm+GkEuPX20zE/zE+ma1MNc0FJhPlgGY0csT4NLmzXqrMsKM9toxhB7B
dUScEC/59+5xpWanYP5ai3dY1tVEr6/u/VUs/lVvDoOEpscGUmMWZWFLzlo7oI67
N7iJfLpgc/fdom7kvk4AAj4pbSZJefj0P4XjCnSdqbH+trc0oZPrHgI9l9RolCNi
s1+wEJZvCm9lW1UpwIenMO3KaPapRkU1TpO25lfxt9NRR4g03Q+WHnv7mmWz0VMy
hcs2kHh6zv1BGC0bOa3CEt9reAPDRt7z1F5wCMAxYqEoiPdINe7jKkYmr7Z22vg1
wqziMw4fwHlHyVU1SUY5pTIgQe7hh62+H/VwZitLzbFbYr3s2SzgiG2gl5YZFuKj
4jwFRM6CiS+yRPKe5yfpnlFB/neNqDBXSB34ZJLKAfqiVNjlG9Q329PAYE3yEUwK
WOYyPZfvXp0ReQFhPtyEDfvotMwhP9alU99oyHEZz0wcK/w/KLZuRnz8jPCAQA28
Pd/DyDuFX6LWdobR9Qq9WubOMfMWzSRzO6cAbAd5mErm6KHBvL/kNPr11O8E87Zh
TBEUgltOfT1zjmL0sH5vmrvqc3TduEljT0Jzdg0uCzchE8FQAVnuO391uV49eg4v
U399Jg7rFDFPSnUcugN2h1H7aqft7PzfPb2rktC3WhUGM1+5MEf8pJF/eQQmLSSI
Ybd6ZAtITy8f2QHg+l0sL/GfZyWG/7u0DTqiKt28fdx35wpNVL9Ylsp6HKO92kKG
uAPsxaX6na0KHlLLa+nuCg57L1d2pvvEOcx/4ccEjnTX6egpDns+vaCGyy0S4/BF
PtK5wK2BQ+eGbVp6UkgturHUpbefwblgbjUZ0UkYQIL+p4mvwjXVu2hHDn9H/4NJ
rSNPyNhTpx5d26WE+IYuQ/uwGw5DOVyUmgFRtxJCi5ZrwlkpsEWeXfEwYUi3ejss
lLpIuyqUw/YMSBF/xI0qpuRsFlGgNCtF/mYi9xsU8q/W4N5/bpSwurkkd6EMZvNp
2mrG509kPhCM7QlxEuDzxyWB7QPauiSP1R8g4KMpwk/WeqRFtF+QRMZGVOqFEn+L
1XU3JKvm+c/Asw7dsM4PorLvCLfQrlQNh+0E5Ta09CzDmmA47JuyIk5HTzHYj7zX
nYJR18fgWSCq2njgmUqJc1qHWShBuaCXzwNuU0Eov4QJroOJJK/U7akOiudRules
nLo/X8ARtLj/7KXRDumww31XMSCosezDKTN/O7uV8t9hUvn21p8iwFmwR0XtdRGo
HAYayNESogYQZvpaj5kpWsZKcM5nsDvzN3epidtfr51HUMCb9hE7lbPoh/emSUoj
andOepcKnw0AZA1AC7nQRTjKnauOioUREFGld5fwVZx5ltEheeEdu6Y2vWcbF7gu
YhyT31gxRaUkLFFhha3mEzRvX/XiXsVxd9vtzyTIE9T2bRg1xS5fod+aiVRnkVOX
rLIhmNZzrk6O7RSutpQ4QjAH/5ClvTUUg9QGpjsLRQx6qeoYwtRUl5UkDURiKKFd
47UKttkP29dn8exmT+27v6PQYLzrsm6pdllkgf+fnsfFIyS8EJyBk6HbbXnoAalU
VRIGcy2cvW01mklawgWwUxhfdX4FmXANqpOAa/SK67LP3fxOW/r6YuQVNMPQs7MH
MwnIuSs6za8Cq+egj8EpYoTNyTQz8qTfTBPfMmwJk//0W25J8Jt5RVVBlgNAxito
34C9JSj+uOxbcZD1v8ctU2a3Dk0eL069m5UBJtBfrk0sm/qlPjKIyF/fGPXEoNza
iGSYR1po/uNMskHtGvPSLglCeAOsF6+qrcGbbOYbBKTl3LxY8jP+zcIH4tthEFIT
beQZBHgSQi3hdGarnZFG44HRaFNLBLihAR42frE8ChdMBV4m454BMRHpjdz6B4pY
tbeuUNAvQY8OvdCdY+wt6bSxhHqJzi0iVb1SeFrGquSG7IzRLHrrKAgudncw9onH
rWd6N7Ch7Ka4HPtOWK/CX7bPLgRKl2kLp0Sh9GaaXt9jG5mvvNEb7D51IdxaJzq2
4f9O7WsXGmxmADR2Z1iiJYGZI+7j1DGy3sO2v1w9hRh8STPUlAERc+fDqniwHgKr
MLXf4WUSs9eBSrobK18D1Oh81rL4dZQRJ9ajKagl73PJ/hDWA2+3PMDbpxAufIkM
qReD9ZQC2L7oZf1wwer1eZjoMN5psy15iCObXLi0UIagI5Xov3EVcrG2vcwSosGG
gUhawx365jm+YOw0lcyGxdWCGWWX+GTE7UCdGwOnDNCDpemelGT6qNb9PE9zU+al
6USAd9xWJQfCSOIUgJf9W065N6Va4WMAe1R+amFO7qmofTgzmFbDw2KmG7FZJMcG
25jeU8q7ObHEF3kg529zPaGRHIN2Bjhn/Xkmp13j3ybDKHkG924EBmjPzRy5NhfD
hgZm+1F74VsuNc5YnN0URENWLvNxS7DcSNj/YHGV8AmA5c1o3j2h0MYuPnt3f2tX
F1zjZWGLQLY4eX4gKaBmcGQWdSNx8z8FV5Nn19MZQA1kr18A4B6ajiLnRIDK8qrB
gMkrnm/H0IHoIkeVWVEYX99gfK7Sxmxuo5otXMDeN740tNq84GMQZgWuOlYiTZsh
n6UbhNsNMT1k6DbtWKrE182w5aes2zQ9JEgyJGAJ/Ou7SotM/JTOObE4AYr0jo5s
hy+6XM8aSINcHgMri2SjQHp74P8okByppdX7J83WQ1Ni2Rpr55DxhPqoWpdkSuF5
i2qlRYlF8ZLu6YmhuH80k2RutYjMXrd5ae40uiog4fNG9dqdKNOti7Arezbdo2ZZ
55FO1kIWGjOolWSIHT7JiQLatfILK5TVdPIub+oki9GjKLTgscQYSddbx9ao+Y2i
Rx3Xjdc2Ow+qmMp3X7qpEpl7v2RM3Hqc7eUHiJ/AMJrEMaQbCd0247ZNMm2+uvil
I2R0jkZI3dgAQy3+8IKu4XjQ/+ata18QqWSBAUEQzrKCpcF8ybD5xIULLIUf2bVZ
/q3ZXIqzW/mBcA1ZTOmE5uDqSzSozarYj+S4U9pRAD6ZKXT/O2Ks6CkXqL882my0
vRU1x+lxIbFSSoRAVpGZcAD04y+TXqHPVDUShGPA0nXqpcloIh7LuxPX/WAEpHxf
fwNzhKbNowPUW0SrYz4f6RoHUWY5uTKyQNOEkOTtVV7VP3k9aQ+OsXKnR9974NFO
cFwXB4/vnhjMy9dRDrS1ib5nBo/wDdRflvoC5BrDS1bGDq4iulVI+D/shZlb2zHz
yco4ytRmkuDB/Lahj/074FZw+ev3ObMvEIPM13sNMmdHZ05SoqQyMZhcrWNNwv70
qIuH9mEYeUIVa4NnSFVQ3eyJK+Kyg777y7Mw5WmD+fm0IY8NRHvkFUiklTpBE0WX
LwDYSglWY8+RWUwmolTDfEYq6rJsJJ/1detNcfn8brUVO+TN2lrjtd1fUyl9VYos
+9bcvC8i91992+jlDFqbu6ypm7eBgjMeeiIKnBBdMPAq20uZEDHaE+6POyslyiLd
z2DPvnGNc/kjwMcmZn9uiuwHCkFKllnFU5KCdYnVBjGR5XoYm9z1o0lROZEpF8F1
/56BizZN12ufpULpPLLH1YLGusYj7rWSTDZzt99bgepoUaXRMHAJaeuZ7gHSTqRA
ZmdBr1a/L8kuDrwvrdCPlc6d6lOiOeIS28URFlX5+JpPvdLDZ1lVfP1UIJfx3URk
`pragma protect end_protected
