// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sO+OWAQBhMkFL/L/4aIxWgOtiUx5883h0xKxmQcxOSlTXcpaM634T+D//B8ufeas
dxRhV4SoEn2DGrCYvsIEaWXRY1pJAoXHMjnthj5TqRJxA7giAtpECsLU1izQ47cI
Cphk9LBKCAcOzF7qwxU6FuaZoVk6LRR8kh6RBisQDRw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2272)
1nJLEvddSNoIsID8aglDDBzAs6CUKl/UcXQHnF2nonbHWQLh8ok7pJtVMmcf5NU+
X4fHr/U9PmFKNB7qjcw2aDgrWh9wNvMxBal2X5rjrhFxpVTeMCfJM9c4xinaBzOs
x5gk8AjY+y/025BHOX1mB0wnFt4WLDzlvUavf7sSzHqXdYfT01qxTE/5uyozApeE
xBdgmm+7CfNit2Ox14AthKBGGwk1P1pIlKOZAwx3svFP1D3T52otIxDfGCaUvppR
wJV6zc9iX4gMedQiJxn61kUPy0zm6ykPGjgiqWmfa0XrPb8ixx1SnCtGGry1w6u+
QjsGrOyPmOqjYZHGwdjHzLxjCREseYpUnwmN7Fp2Eq78JMDCYDJbfXeYpX6j2bSY
0GyIrhv6bvyqsgclEs7Uhh0TUOmm9/xKF0SAbYDX5Xn3gAKY86D8NitIA4c6T/0C
IOKGEKObKLGTEaYqUdXxTWoVh5cZXv241hOCF7JdfUlkZbO25XNPz7gvt3LO/ClL
qpxfMMsKljSoslzDhDOBHKBkQFRLrqWURlY5T2dCwD5TfB6YtZHsVCaDr4aGO6o3
mPGdkcK/9Zm1VJ5tUClAWy1o90A5c0sCnYcXRiZusJMc1+sk7a+Hup17xMVLaQ/t
lgQhszi/Pnxmk55M6/hNIT2w993cH6QDw0F6FcUwsjZXhYy22BNSjPY7RlPF9acw
BTQ5SNdXyDSgi+clDaqZBZ4+sDxeQDFlQStTRJ3kbgf1FaQs/yGNDWE1XIP53dcS
0/B2v7NChQb788JFKn/YhofhbyzcOxULdHvWSJ+ZmMwYmMSX+PTDuHet4qUvoJG4
MP1+RR4qHF5RrkS5uHxDP2odXoKExnpFoKudVwosTrbPg5vbSjN7f38OXTFlOH8C
aDlZLbo6M651qZyOTplVkUervwCmaUDVtG58KyzsWuQpACFFWQ3f53T1s4HgrsmM
P6LQhkbE8jn5bROxo6WvXYf8gUzLk9WR/dSnxnkRt3avfHqKkh0kyDe9vb5ZMYkb
vg9PjzjqbaziJbqBF1poqK76lsP0vbEEzuzoJJudeCm/RBiqOSBgztYWKYpE2dbO
cjQhbYlZMNxHooRN+l9TicVbiTAszfMYRsF8DdtOsbwnBVjSlRCPFwD5H6s1fFs4
Y5IvjiJ7jrUV1tSExF0o/cLyd888y2HWJ7mAe87e1G1qZetXdYHz64j+2iAXQq62
lbDq4Q6A1AHp5ZnXitub1Bifv2q2dZJVep0wPhocj7PyvyV9ZnVt5oSecbL33Jpl
6ls2XStgBqDdXX2PHYIhY7VV7dbpibFvs8+HM9lg/0zDgoPDGI37hO/BV5RlPJE4
B2iDWlUTwDsnJEleYKUYX831jgSNVtLW7mlraFUC+ap6EnnHs7avjiMT/uPKQsvm
2rLaXgKpcd/Joyyrjj+E2KQB+5EPRKtBgBDel4ESDdzqq06xtrx0GBZO0WRvH2/W
jAzz/bO+X5+ZOoONEfkEeTx1TrAkgfQSJXjHjUm35i+60b3HYwtmUBDfFEj/o/wl
8xyJ+87vG7nSWuhCMn/X/eOxs/7Kyz3i7NzHLAA9GDGgAbDDYs7jrJD0NcmZ0yhY
Gu58qG0wHz4IKPxJTnVXsL+6wROtPQwVzzMXJQIW/1QeN6M0lxaytSkuX3kAuhse
gEefZSiv7cWWqBuGTrQmmfi55lke+l19NAujQuDQZLEJxm1DqbfUp3nJ7uUvvLp1
9sk26ln/IWzpLHq1Tbw0zPhHeOXcyVETvujD5ngmEIHcU/2MoGyv+DTSBbtEqm95
azwbwwTJ+T5xNIEklAJuNuGKmWDhx5T+QnbTzpgddnIwwrn8FLfMNt0Fn9Qv89Kp
zzi8m17efZwNRu/yeIToJIIy4mbNUvx+sdyqTgAfQ7xjSJLauJBwiWzj6F2IzKs5
IzQJo8gW7haFYnnz/qdT/22AfcXrMKZS4L+kXPXeqtspKvkrNc1a9kC/IHvBiwk0
50LYhFejlapORKaaCn8n145/P58pZmNT+E3vBNEPlIx0PckfVvYLsRhEGzcv7nMx
Jz3RWpU1JTWD2q8AQMiQPPHnRhiWjsCcJcCWHIXlDiBSAhya1eDpoOjnKbsm9mrM
puO5r9lekCv90dwWIoEjeRWBTisMKcQlcCsvPH70HPNBNLoyQI2DBMppEPHNjwxx
a4z6nIQLMMyiwqK7AT5zBc9RrL0lK668kzl7F8d/4jSwLMpgXcZoz+NH8sAp/er4
wZXoisxhUT6WR4eF945+/k7J/wPOybnEsIC6YcSKVhkMFvsh1TMmgWvEpPa+P9SF
jdUq1MLRdJwkrLH3/DRKqk4yv7Vas5MbnSe9B8+sz92aBo+Oe//23QRLacMNDVpT
rE0ZWuRANIoDpoccUsnQ6WnxyBbEtnpgJFqtTxDuOIRZepgLhlKtRQfxlqbUxhL5
QPDuomCAyio7XaBJTd01U1B0UoqC3HE3y74mBruzihFBKgKsHnS2we/bh0HsxGqU
pVSDzo63P4P799w/ETIogXg7YYtt/0k20AnVj/KfT5rxoGQAQ665b9cGYHdRM1r4
fBVFUeRmD57mXxTDvYTfjHOOBmTYg6IsgLApm9OAf/tkIoimhtx21O6OKCAgkha2
ZeXiBp1bMTZOkgWAUjnWL5RBcia3DWOJbWTTK4UJ7DK1mwa+NIaciyrBhc0r+pvV
cf9LFaB7sU9+T1lm2lK1/Vrmqngm+8mYLogXYGW6MxDHtKS2xKkfffCnFcpsfTdP
4l/6c42+s3tPXAH34QacvRiKNklbmIn0+RLj3q8TDDDseCxnbtqJS4yC7tFeV9gp
AiAPNge+089s9c7wOm6AkI7K+Doj+zuFWpmsfJMd3rrGQYTIXa7BCYRABMpLtfJK
gBa7892CnEoaLKX6nWFPKpQrw3Oxidy0onkmkk6fmVOiaMA9nXWHVzmy4vhMphxv
/R4NBrS3kY6Npzl53gzfj3CgKPGbQIHGOf55p2I2m1kpi2zAELuFvmCGxbs1M6v9
hHilDffavprEJtm7wuSG3g==
`pragma protect end_protected
