// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tJojiPY2FxDfLJ4Hvd984g2fsY+EOK+DIjmX53I015n0EU2inmnHda4UHzGS5BkP
QCSn1d9cn517s6mxV1Yh9rUr8XsWRPOA4OIdt9RLOa5IuTDE/M+oWlZkv2Rtwqgn
Xt3Omjwbv5cf3cT7OBZGHM+yIe92xY+UTUxLB1k/oxo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13040)
MkZVKtFcjaTiALZHszqcN3z6zZTDe2yFDpAgUslU5pffmeafvumirLtm9ox7vbqT
k12XHnWlGIaMe3SsgN3wIoU2T2pV9EGbyOjBrpSIRufvu3TUEm0XQ1mHPy3U67Lj
DmaM7prXN5UWMsGnZD7AaloEkTioxp7cyqAhvBWtYPuGAOdCpxTBixRA2l+0fAYj
kw9sPx19GMxz3Kwtt6wdaIVreCmapEIKmwocYtikvdMIYOrmStT2NFZTV5HY99la
d7NGmn4Rvz3VqcIl67lgJXlsPp/yfTi5CovbVnLmm7zHPYPMaNulSN9A4p6uohRG
yB2vmyrVgsXPN682BbQQFLqfUyP5+LSGTEniQ9ncf7unR0HaOfChaCXrZfZzjWwu
TlfU09lfIIBYztPHo9h3ippBuxdMM6TLicGhn6Z2IuKYtcI7VHugUIdGfEgkfy4N
i2v7m8978OyeKI0xUPy8D8axniJP8SP8I3vCug/1otNtJKJovN4TumzrdX/Bp/BG
ZeHC8fuFP5Q/ZGAgbd6/JcJvVmwjXIKqFTIvViRP2rmAZ5sVwwZmGabNErxV2eNp
XHnzkowhHhjhIEh/9kb/OX3hcelokUQ07Q2kAQmMUa+/o3rgcnhbdw8bNVOg4DfV
3TLk7OqHiagxELOxCHLV4xi4mhXYyhhkd9XCr5+al9IY1T7h7yAaRagrfspdEfZq
0hMnIbZThoSziYM03ovW6wSI0m7I2V3hK8n8XRxUeGraH1ideeIA8LLBc1LSfh4B
yuJVpvBj58JDViTZxywLZJY/Fp17kCZpsN1XUZaszQC1vqezcvyU/do3+ptaia4p
mqNGjeGmOd3D9jjyCEn9VCmAkkhZc17fKV2OuSZzVdg+dgIhurjWS8ZrbxNZOjLH
o29tgD+2l/mrS7yUz3y2in9+C3hxQnHSRlHKi3FCt1J5q6LgRCmL/S2MiIAGXNRE
CuHw6wCWzJG47n06HFEoJo1iQB6Xcvsns9adoGezGhZXsJwsV6nygMV1lUKxDWjL
AzpBFCwkg2bB0DrQO6Lf/FBK7oiCHm6GZ5uIwpz/Vbqi9rWN8qibYiamvTY7t50v
9Eq1E/NYQXvI9JVJsVqHayhvWZ/cmQbAdjEG5NTZGYBLfziWrZnrgd336nS1YSuE
kS3Tw4GEEPQAyWghkg1LJqb23oxYhp5WDTRIN/YhYhzipaPKB8le7CkVzDQbyf3E
L6NjuDdzzNm8X1fQi9DeW1lZ22/iTZaqXSFCp9VF+xLU4GG+3sbth9tau1/Mcmr9
Yv5vbnA77syjIb3lgrPseVdFqK2hsHX3mA/v481TvKCHNdvnzEtFziHkV1yMDMwi
9zno8xhWT9kCiQnVtNI1+bLHs/NK0TD4pyERsNNMUfKMXNTYjCeE9mnIuW0FuxTn
gDZcpMXXkbEIwvEvKid5jFEydn4LAPcxB1TKxhUEh6Zr9neRYdUhC4pLbh4RR/qL
c2HkhbxNupd6wys0XNGnzE54q2c2PvEjNzL2JUTay3mfCGbEySteKT3IWGOEjCII
5+kt4xVje+ABbL/SGeJPAYl2qn8u5jW6VnwMPUj9KFKlubqf6lNa00B+QvLh60/K
MBjuY7yBpF+3tWGSDB/0468bRzwSjV1lu7f9cDB0nOWWgaZOCOeHNUQx/ObfLKX2
MYYKL4DShn+LidWOL1rdtDOAkfVkMDdYHpj4JGqg2XkiRhMEQnbMQREQf2pW9jSC
jJLwCpVWLsDD0oIUyhpcEGSo+8BGeOSKrnBNkDM8rN4PKBHDkRmsUFzMWOmiyHsV
WkJSxS0OSeMoSnDCn7CDv0Bfa6+i4rPixxh9qRMQ/Am/me9MJx2wt0xNrTVybIue
xYe7ztHcG9KKpUZKcNNzw3TbjJ040bjV55+weHlsr0KuU0lagQAYqpe9OolK/uBB
LGj2NZ9+t4Cqf/Uwpfz4pe0r4GpT9XdGW4LrDHBTpr6iC/k8glEF+ZZ7GCiABpfe
eCxAPtd9Ycxy7g39sZhgLIwWrnNNSbC6IX6ZGiPXSHedUkd7NOxiJp+2gnNCn0yn
8Jk3lsRRUrf1265HQmqkNub36J8ZfOuoJHnefFr48REIB2jjkPXjfsoutSxXR8SE
qG7au53XSA4rFicWghGNsKzKkt5RTvWGfpN2sjpVRYokRL7wKo+vdJCqaLmsU86K
fYOZgD2qIy6FsxnST8xdmqA3+fMw5/h+De8zwkZH/D+NCi7/cJ7m5t1boXjhPbO/
6nxuoxJRGj8phK3LXomOxyKSKRiIbf12oC0DAYxiT6r9rELiN7vUbXP3pLN0vXhK
EHYK9Mk6H+u38TP4p7dK2YpZFjWlMJ0iW/vpA5t79zyZphPD3eP5BZEOpEvJeRDh
nL1u5G8cbHe1PwOMThcztSddwbYGZRzSyPon5Mx4R3PFQ0BJiufX+9bcXQNWaj9j
FT3P/3LOUtVXxAGzyzCx3ZqLI2kjq07bw6gM2PvU289menp+Hsar5OJohGzgb9kJ
l97K3ikfpIjcCR9CNcPWucG1Q42w5O7vVpneO+vqH8gzQND+Q39UIGhbHlytMQ7U
2KuMQhpJzNilos4pdPWW6qIjPpwX8qbfPnPzg/mRZseU1ng1LtXshp6+pwVDvoOD
JFVnUy92bpj1Y0vqp3kuMXfCDwJ0q2WcGyUTd5K55nSYmHH+QHjI2ic+RdRDJJ3z
00IKfGtEDbgaifXuuwoMSr2UTQG7XrE/UmF1dcdi8XQqTJqVhe9M8HbBXXYMogwl
DvY+geCl4hvKSkvl9YPlZEH+Y8nDuqUFBp1mUK7u+rF4r0Vzisc58zgXnY3kM2Bf
PbiZtWpSnuceYr9s/swgHDpQVti6PV4qCxLGWG08cTxtL1f+FB8ZcPDqA6mdnV7d
EnnNOW0fGHRkjXFPJvA2/zflm5m/75/FpQIcVSJYrO4qKs1umnwcTMlQTAOw6aYZ
JVd/WBkNPN9sZ/Q1lr/wF//som9bdgOsiRb46y/pEK5xS2T2tFy/JK/po9uwqRQB
03gWoG8WZ3s5ScC140Aw6zISyK8uUnY9atwRSqqrdUmnFZzxpstGd+tC/MRb82O1
F0zY4zDnWzyetId38tJS3CQiVBS0sN02x/JC9tSeXIIz51nid5VgBxzSDG06UR36
VPRTBDmcTEHUt2j6R38XQRU8aILdpKVb9FhLQgdsS2W5Np3p/oVpszkv9zNCC6I+
/xgNRl/W8i8puWQz03/1gVK77EwDDDuogf0P1/HoRfE8fA3gQp2tZvhlhq/LrIAa
BxwjqOEfCpimt08u0U1YbE6E08JZaxxpT+kXBFNXDGgqIPMnLZp/DlCTC7QP98HG
iLf9dMrf6QEzlAgHA0fLMK6lNr27RjBuWEJea47nWzHIbtJIy+QZeH7KYkotFOIT
UkBktO5Fk2CpBccKWpdrG2Mbp0rb3oCyJygwJmjbMWYsbCK3EA8rmNXcmkEz3FG9
SCsgLK/cZLGTZdDF1E22fB2fJ4lfGxAK1FxWgstUSSlZlFd0eL+RB3FQAvEflWpa
FmI0zVMDQXHcxwmmqf8HOxvd/1NDUgqx6QF8wlR+D9xMrPRSufZ0ssnYso004FxH
Hjr5ruKb0wMHsWEed82OylO10uC7KGK3gHGM52XqK/Uu1cqMdwXq64XIO4cSOm42
qq9opre8L+hy71Pchr/dazbREtS6A4t0D+RIotW0LrY8fjuxiB6F6vgRgUvPxLOs
N45GlW47/zAMWqrKlcEnKlFMG9jK6fouFAZEYj2ntcyYgPXwt3P4U7ZrMJLGK5Ga
8t7n4IYpypn0apQlJWqRYjJJjn9/6WlWySTEsfE/KDoYN+ECaFggCLsgaFsqi8OM
Uzc/3fOslDKYIvtMIpIqejuFlRi1HLbIRaoW77rX0V67AGc9pAGXtIJS9tw79Xct
TNiho+iyNDnxb8xd+uzIhs2sh70LyZ5Y97eBnQ3Uak8Ji1I8YZRfI/LluWaulFqQ
5Cxh1/unZeNQmMsQ2l+U1IpSUUrsPehzZusTlO2OvAW6oXOqL/Lo/y3s/JktT3xc
RL1mhSUO+Cl/cE1MpBPF+23fjRiFDrp5AVYNgcl39wXOyBzSE0b/jj3ygqotWdkV
jKQE6v1pfNlgiBrHpwdt+UbpfDP0WJC8ISINTngs2Z8NQyk1sKSM7Tmcm7T4xn6o
x3Q4KtwwKgjCM2+auyJTLQ9fmACXme4N8q+jJMAncHkIIwXdf5tRlMnl5m6l8SZH
TZhSesvdKpT4L/kDJ7Q7x7kRle9kQ+lq1+YkCbO/hcPe9IvcnEoIQbbdcB+7oeaA
gIWoF1xjsCKqM8eICTyA4HyA2wbUt5bLwjebMxNfQND3Utk3EucE9ho7ixmO+KKg
Oc1egAyM18Ue2WgHvdIf22nX8kRU1m6N/GOumSf2ArUxMMQqYkEADEljnpxl3hjv
3rc3Y9PyJVDdGNdcH1ACqk5nw7EDYqyjKu5ptLmJs0qpckoslano3mRyT8ZQN8WL
bhWGLUCZ0HEZ34GCfvoxLWLwwO3Vl3Bf2pomiQTmTlKbOvGbnn+KZ7iQUxoCOMiO
HrCKNIGqNri05Ds59N+DjP3K4tDWx04PfK9kt1F8/5QWfY9bg8w+2e6VkRlLY74t
DYJLsNj31NbP1NYQPA+x/WSqcWwg5X0SGLpC1PPEMMugnD9LLu/yJ6JOVmAAb1tl
Hu2T76o/TaBujMjI4huz/g4cg3140NFzeFKIi94yoRW1LbNZKvx67+ajqj6hH58m
MCLRRaSJ9adpumtO4uO20lyYYsGNPhByYWwOWHWDZjVAqbU7X/EU/sg9jY6YzAn6
v1QsYf7GW5FhMXRdPjCFTZ0ZO99yxzai3s4JZmUrc6cGOfzo//rpATUIGh99QK8a
mm4mBrNf1qv/nMbWDhI5UxgGBLVP7DQ5orOGRqsJPxYccVm8QHKNF8uwyGltQ+7j
xgzxPzLwC+Pm1meZclZ6LuOvodY+6XXQc3dusrkeoveeCDx27xKiAitcnmMXtaoF
36km2tgiSClIITUIlO0UM3ZJD7H1LTk8fwKnCjuMsFr7/mLYyr592cF6MxYALSci
cpLRDl3wrOY61pp7EeEz64sEczfg1Z5O1CMY981o8OEMmUC7q6ddboXiiCTD/JVt
6mryBGTXxyF9ppOrWbRv6AehD+oHYJ0ryHCWKEfhIbXaaMQOW79qSZ45oNi/j5KJ
F7kowplZU5enPfDS9PIArkDFTVhttD0Kim6wIBVrBGsChVWGOyC7Sms81CIOb6uR
tNAXAqqUev9l+tolHuriDSYXs207tMMPGRY+Q2eBA1T+yGhr1YP5mzWZKMerVeoc
BjxMtcK18OdAJA1m5e3sTW/qABwq+RFYJAozHJRdP3IS6A8IjETZbpBoOPLjX+7C
0dfk3ZHTJVwQ6/5KFXbrkQxIKpcFRMTyQHjZd4gtv51p4TP3xGIpX8MSbLq3zCVU
869qTaMOcVxpzigtC1XwKWOkJUoFrppi02FvozcmBQ6O9+pmyNtcvoMt42OM9+SF
0cvWEUqXnQj1WOymH+X1peg1AWgkIq3SBF6a4BkKp1qCOfIqDujXyNDYg7df3pS9
c9B/rtP/GWMCixL+HXjgiZHiKN4k6W15Cd7a5xgjYMqv0l4+K52LlZ0olInNH+iy
ULCW6xNWPeFr5exuGu49+Xd71k5vDepDAsZVRjrqn9UIRvaFcKDSent0rYdBaTVw
Nr1C9+god60nY0M7ShmQDVNapTahow2iJTRC8tYHlzmXiigUWrDMJY5EI67XLykE
11j+AE6uJNebXHfBix288bGeTPpV2zojJENapOjNEri+KaXYHlihkQs31XDXyC4K
uIBpqbQLLYDz91EFcn3HJiZxV8k2bnkVznH4X6+T2Cj3wa3x48jX/PYh0BZ4vOa8
FnFT0UrN2t5EEIKvNZYPTJNe3Fa20eHtH65PXoj1FGW7wvRIVg1sBEmTs9jwYL7I
HvrBmo5YsXOAcQ/3E0FVK9iHpW+6VWz1PjA8OlRrkrIfJ+5B5t8QzPv43RLSW2Z8
XANEBYs3QGRSmfItjeD+1p+JW7sH/t50Lq3YI8zUosArCscqhd5raOQXygYZ24Q/
Vy7h5KCKZ+1mhl41sk2SDER4QSBLJ67cIOQX55NoPJ80qZmX0K6WCKPZTrgFKcpa
zqs26c4nJDjiaHqOMYEVt+2532Wo70lK7wjGf/IzhWNx3ZcCsV0f2huyb+JMKZ0R
0yNd7ez71YtgG5V8UIaX1vV79Q4vP0Ds9wRX2ylPQfQnUp2w2boKz00GN1QsbIIP
U5bjdZpbO3qgroL9aDOD0tUd5FBQUuLxKy3nmTdJF4y1LVWbaKhCEXKhbMp7S0lr
Wvl9CBsqG096rR29Dro2G/I1qRYa5QUSs7TumL4VxfFVFcTuTPNLe7ZjJB3IEf2F
e2QEImLXnUUTQwX0llDLqupRC23ESk2HTdf14klGqOsspcYO6XJIIIoEsVcALwfN
rGH4vhy+QzFJ3j0wQm8DElHDU/ZBeWn6zvjVgS98sAQAMh+LpPPDr/yS+mdF7keH
e4xLqTehn/B63mjWv6F8XvFiTeq0VKOmk1CCgyfXhfPohHwrC4KVbxo1K1PuMPNr
6H05jRrf0OJ9S6jpSgQpK4410IMCgB221LA8vWGESBotn6EcSob82gWFf6e3KWWw
r+GC7sTKTAzu75CPJVbCPkIVFrz2qFpE6geWxHtBcRDzFBWESSgKQZSstgZ3zCdS
/a+VZqQ1rrP6XkyJNjZLgheR8ygfwkCSX1L3+tA/TpSd98/IT2k/eJ5SJ59QkQD6
y22CBlmxx3TZbUSG7fZZXK8xRSbk82hAyRGe1OVk33vcSLUXThepGwkHwU7W+ghF
vsaYOn/gXwmYQSxmtjLzLY1Ykv3O7qemDdOBZU6OGTGV/HfEWOXakSIszhkW+fkC
/lDXtRmFNQOkeRlz1f3kLSEXi2Do+yftgVdQZFoX4s87Ax4e5oK/M2ZIcDeP/DLC
myKgw+wjMy180MolaBZ3j0S+q8ac3UD/SM9zQWaZGCrzIVRaxS9I3Z1xfiEWbDID
l1rc6L+oc+YQT6TwPPjlHqyFr5GTngJyiY6TPTVQ7m4665acUqsTQcup1YiJ9fqL
K0THBFa5RCYDUTvuh1aCmNWzpjN9O+hzvdOYLkFtKmDDWcCD3HCiJ4hd4Z80J08E
MX7iSKVU/B9K6GtxEXelDDmMgdHT1xF4BjeDeYZZ/TiBWgkGdPxybTFsTMRJs9/Y
KKq5lOAJQ4Xb6NZ5htJqGFfhUMYgClKRsEbZ5HqqQU4H78wa69UyNF0fonZk3+5H
dZsmEWg0kcTa7JJqgDi7RFTquwJc9kYfdYX09p65mE/3FEiorAUoTNvqxcJhMTQE
p0mSvtvxSLR+gGEpsdp0yGmErWB3aOMKwbrnYXHJusVSqyFavkmovColcFFUQZZH
9/oixP4iMUS0BVutb6J2+fMWkV5Qecy2Kx4M2okkiN37zql03v70AKq+hru3eLtY
kTYIgAKTJRXI6TMVa894hFk1PjrXHKUH1vUAhEcOhuhOcLIygDjCqUKUSH42gy8S
pxtVhFHzARuXJ8zWE8EOnWg3lkfMYKUM8Twv1p7w7gNjT0YcD3wysBlHcgs2YKAt
t0dotbDdvNuMIitdtsLA9PqpJd+YC4QZeiVw0lP0Tgj3ENVcLUJVZFhlz862q0Ea
E7g/b4ZdCAe1c6D/csdOb+RbVoFXmzoGDbWQg+7U73q/NzqLAnH2mXRsBFYcsxgl
FLhnKA8C3h2wPtH5hkDq0g3iE3aSH2+B+C1RP00GXFGAc5KBjM9YcvTwAOidOjZ4
lMXqkpCA3ox3h+gumPRWjzhKuEvpXBySeNFrqpPpUL/tseOiK88DzAf10IQoHZAk
/+WrOObdD1CZi8IhA87cwfUHImIjctN8hpLiw3cJhkyZ0rf+rF5ghrrQWxy/+h2i
HHqzVAaV5oX3fW7GQfBSui/UjFnmxS4VAOjPDI5mQAFdo/1ImLa8g92XWbuzGr5i
bf30b2hj0WTzRwdu944yb+BcODhlMR07hPOyR6o/u3JI33/2/lHVQ/f99y2mDFS8
5YdzIlxJC7w8OBQyce+JvtKz2PxT0ar5A+iu05wObjqgO8W62n+GR6l1A1jAS99O
dqlSC9jwdC1wMTc3Uco/8sVtUJ8sisWFle9UGxL8ABA4XdzgJ3KUBYP8+cHbubMm
owJWpQLVHx1+ujAEiWJBp3E5EecTwy9WbtJRaYkoLxkmge25Sr5nBYEwxPrJDMiu
Jn8F8lvZ3Ufd9FjMglmBtwSGwHl9Uy9+sdYQkVXu+sxZuZz0OVEGLxxdioC7fWSV
tfw23hP3iwDDxLjz8KYG32yhgY8ciXxHc/Deaq/MvoB5a3yUQjeyX68JAE7ct/yh
VD2e8UUgFV3IQbDFgMKFrnOea0heRC0o8B73ondv5Pbos7VbBe3URkV16JuWRY28
D4l9WYVoon0tJdvfcVTyN1bJ/zNSBpGhYQwBtDMQEhhXf+dBeaz59AOYVWJUPn5S
9cTQbAS2XDm4fylofIneJYPQK52Dx4tO4T7xGbq46eIj8E3X1U0L+GSGd3/vna/L
D7LnEjyJ+aj8GOCwTE4vTKKxZb1XBRoii9zLYwKpeuH+2BuVlRNoep8vSUTrYCUe
pUQWWX6fG3S9fpfj5+yigwsf81OGZxFx9SEtYwU8XWxzlDyierQHI4aGUyj2ko2J
BaZAau1jiiDTqGnaVYnNyN5murM+Kmmo/nvGTTqBaURpZXiCDaW1/v6zPl8GaPMf
CON93wdf/YO5H2axwRFO2IvCf7nO3eP0yUVzMbMluNOV7tIhx+7yMW12EakTYPfY
rIwBkFzQdsEfKRTjTRlZbYhxFTJe6NyvntX05O21a8AUBcn8L2/OQRlkIw+os0kj
iaUQey9fnfaA4raEMovBsC1OBLASncYRI9n2lO7kRo63zPp0v3fpPvIc62Cd+Rfj
youEbUH9rduUzAdPFOgHkYxWYsFrRWEUUzE2FvF8quvaz3B9sASLQN956WGZUv/U
bJS2yhVn277X4YuV0XovgbSzxnsDBJhF4rI9DwA6ExNe7ZuPr9Q/hhkVfTeY+XTA
BmyBChN4Nwoqamehn3B9q2NqCwK/hgZBaQZkt2FL+35UK+6tkXyfvaKUPkA7HGHC
CFvNkgtQbPiKAXzqIPpy/T/muI/4ULyoNAAb85sZ6fBjxIMvJK15GKR5kuFSDtXx
wNjcLpvWixgsoicN42nxiJm3pGBdSYyeTidlA1OMY2gPnjK1/sC9eaMqKEOHHdPS
baybPWpMqdtYNI4YVvRcui4qoRQwd6VUjbRNTG4Cy7xIOWt/EvBJ6XabwMNfDQeJ
tA7fzWfl/XG1gAKv5GO7HWbU8XiqPYt1wx3SBYbuBtxMgr5wqO7ZonrjShJyl7AW
mdr5OOvzewSEcokoGzyxHcLMYfImhx3rwDFO/1ZQtXC/shpbLXNrnOk2QkAf+k/z
j8CfQV5mOEhwx6oI7+9dKm/qlKrlCjDB1fTAvi+xV1eaOTiB6wvxFnssfAqLjLOv
V/K14EOBmHQUEYFEDO58DPcLjLwSZ9PYZBQH6hpngM4db+EoIad4jCIG5cU4t0sJ
4KPVi0PocGK5JwOb3w51yedilVao1QL3f9jgM5sxbm8/I4lEIGUoQWc5IKdwXzgZ
XkAcGCbYRvulmEJpMn2Wp+ZG111srg+V4511rcTyNigjDWikP/xvda5+Ue9p4fRO
OvR+P0T1gU4Ke4GUyIfwni0ggijdBPu8ryUnh2wdIDzrNhOhkMCvVrkPvIlcLYKJ
Tx7ONSyFvw5W1hxPfgGnduOMDCotxyRtebjt2jeH83Q0NSpRXjSAyVl6uczn89lq
Alw+uChf1V80VAilU6PSIqoIfR56ddxKCTuwBfXeJlhueWoLPqsgY8UOk8Laju3U
ceGNBFcfdCmWg9V9Z8ROuhXdHV7U7UwvJIusio23Ecv2v/pXMWhQwuAu69h9k+q2
/CpsCQcEjaH33qIhZjf1QZQM9cNmwLwr/uYkyXafdlPiIgVXNMzpGrS7esz/7wB8
WbQXoxiVgZGDX6LMDl2pUDKFCzlocriCgS3eDvVHeF+wfGwd2gWt9dcvqSDneC6Q
ruZJhAbXzHUeaTZo22dNoO9nr5Rv22MPCKJnr1QRxkBDGRG4e9e7ROftJGlBNhJo
mt5Pw1b0t7TnHGTWzb4U9rPqFWbHkCK34596UXC9MBq0eBolMabL0mXuxowW9bP8
zdfQwggdaQNUOzLMKecFxEKBokFrg5Duv9tDTUaC4DArL+qy0M7Joomd0RyBzgWj
rMBR3MRh/2SiECgR6wgbDPXnq79jv01pEz++IynoysuMTykxiqpLQtfsUv2VzwIu
ZWtdA8A5N+K2tbDAaRS5fgagFMkkFwEs3bCtj93cQRGg//yvID34MS4jhx2j3Qs7
DOlN097qlDFXBKw6nMT2qJyekSeeYUBEzIK4EhJCyeZWK1g7A11GlwClqx8NvY5/
uxQ6KL6R4JRz5dbBgygPAZ/Fim3SWj5CVmWsQeQNTFuM1ZCFWCKmnAi1ptnPwsfx
PyqBwoX8lGThWMkbthiaFobRYu5s6eSTp2eUHIrGuHGgWctxIn3OHKX3DrN7bLVq
W0aYXAoCrlSY+bLLgtJwLdT1Var8AgXoY2mYRt877drKfWZ4/6nOa4E2Vtrufjdu
lEww6GqgdaBOJLjp+8H//F2BpFv5nc/u5woRSxYwZQ2XoAimg0OwZPJ4RDSLg6CY
VfPp1FiDKoU6iL/ETzkgWYshHJalwUym0LqByod8DHWf6muGXvwC7l9/ixHv0XLn
ni6VxEoDbEueHKfi+onaeuSPlzMUsYgOUrTfg4oW4y1EiyAxNQFJuVHNDT4FObTZ
R/SQiiTB5L9JeBJPhXqr4fExU36ilawOCKp0k9n/G0ajZbaRtX0t+h7ynCe/GgZ9
elINSrPMjwnc37WnOCLLSoXr4v6CNEgcnhCLrEFWBgOPyHJW0uZVVi4ypVvlz/A2
nRh/zCApG7vzoWw2sHjqhhOf3gVw+7qDbqxxPx9M1cLEL8Rhx2cS3s1cVGdZizSt
oEMEN10VxXk2wMCmU4ZCzxf7LfZ3GL+gaCnXDjnN79v/X73S2zQNooRHixnjgCW+
CTnfVoHWYomEP3Tlmh3gAd5PfwPWrsxwudnE/bBftV2LXPdFj3Wc/3sj2AweHqDw
2z2MkgeU7Ji7MS61mJeaccvOGDsK/cnYSczih8hdAK4hWNhNeu9JHdQRaxuHzAJp
F6c4eSTVuVHFTbNlkazj9JbV4cU67tY6vcrTkaMccQP3b8ynI4uhY63qM5wkUEMr
u2VAwMACnBkBiznyW6/rSgmNbxB1vBVCv6SCzLvzNSZhzwsfIdB53w5feg4AiD+G
BkZGPlaCWoxZ7IKgqVozbQS5cFCh1R04zxrRFDKaAjzk5vPfzLN4gHq5/uQb7o7I
zNJE31qlAAsUHRhbyvQVyka25BV+q9ztKGo5jUzdkolQk2HL5pncMVDdW8QTzlxI
z1PBOjceovZv0JfGwXX8NTp6aM7EawA79hpMx+hQHar58Zvqc8VRWWjAZ77eyddb
/BqWCE/TJhIlc1f+5isI4hZc0EqwDfwIJ8AI6yiOZozkwykO4AWzS06MCb+k0Zsc
k1K+JayBHTJ71ltTiG8/SZz1sc/kDq1+3Gz8+Sgo6reLr0PKQqA3GUua77vqudkf
pkzzW55NLXzXvF7eS2bBRL/u/2EemspdbnBpsHyfD3KDsevF8Pyd9YhZNw3cbtyk
KsV4sRDwCLlnlU9k4itPbXg/EjfkIxMgnQa2p/8q3rtPWB9iHhyuGR9F0YlkTWVg
gzgFCTwOoKEY4WzJf1MlmBuqJM4NuxZvZvZh1Ww52l/x7yqG4aFipnb60XUUCThr
05Bkh0OzjC67dwLpreFXnnDhyRsVXLlnbm+UpxHjHjsq5lCMZisneQLE30fJRWeb
1zq/cISlEDxsm5EUgYntHUzvq5GlG3wMDpOJGxHnKPx0F3O2wNYttxj0a9KwaGdk
IhbGcFUHYTLKlHF3cYAboi3qBUHT52qaAzGSGKN82TtoAlQKEXPDcZPbsbxJYI6W
ruyE9AuoTA8M6WnLD+5rxFbHpislokWcLYkDFfQtuRjRt7V9houSGMDo67nf3/6l
u47v+V3fofHx+98Ng1C+lk35eJnQrXXm22Ag/7Kp4Ur2D2JAO5MD/aZC3C1aaTi/
sMZVLMsjlxXbOh+9rE8Uun/FPXcPNfPOEGuzKZs8Rdd9rdEL+4bRNqhjC5GdBdzB
GnczCmj2jRtt7LODuOraPNMKwgrO9Sdiv/qlscPgxmz8idog01AYeV7n8v92QiyA
nMuBT7gSuJ0PgiSmfpWAGNGYjxBCTC/z7KmSyqMEDdVK0jtZgi/F9GGGMr6ja3LR
0EUmYJ9H+cwljztLHajjzo88rUQahNvSYM2UPRU+4uhHHuHKF8cv5ovq2Awgxy7B
gQxF5bqjc4axZR+uLKJxEn+h5BtcRW4aEdIrgtWQsI/T+AMEb4Yk/xgP2rSkWw2o
9vR5CFrsOlNVH7e+JOLLQND8PEjLwv5luX4cAlZLvwWpvb9wWNctK0Y0My4g2oti
vgQWLTr5IEPsPAcXeErefTPaQXbAAn5/G3+38ZwwuMI8FnOmu9zn9zurblu2Np3E
364l8/ri+otC5Ln0/o7lgEoOjNcQjHi2rAh9dJCoOO+EHqUN2uT+CTLXgVCZPefB
zgadoQQB1vAMZM/CjMbB0jAx2F03icV7U3ngAXIJ6DbHyzzHsnnvQ7OdV8lWeIJS
cPRZqf615H6iPZ+ZnwEyvCARVzjKZwt9iGGMcdvo2a/2fYwgv6F344N/qKCrgW14
kb112RAi4JhPA1jyiA2wQtko7D68WhH/mKl9rA+xHD0Ee3hokeWNWIU+4oavWvit
lT9/A8hywgL4X6IpQ54KJ8zeuXMjnydC8ZrirGoPm7uB41uEbJmOWIK4DDod206g
IVH8+CkT3eljWf3qxL2wxEKcieMAQpMRFhIlXMZgCKU6/pbXDqiRGIxW/7qgBAwx
segqAN39aznlTv++l63hyTbHbrG8VLRw5ZGUwdOMjTLz6vGTPCZqNe7szNZntoj/
vsSyBOywVe2UgLd0UXtWaSjINdf2wY3VloPUHiwe4CNsOIH5FKjs/Jh101o1gAbS
ItnUPNXGw5yEWP+r0UxDjygEOEx/HJqWGLPcZRbza5aqmAfjJN81zBPVJlycVcZB
jLS2vSqYCXKpe8Eg7q1mxKjyG6uWsTt8acEBFtOGPTZ6ch0iKLRYxHzYyTGEYMor
ZKHIfM5vDQsdhYhGOB7b3K8vwSPu1eDODxOEnXwvh8+Uu2NKAPs4ZGmFoStZVuAJ
iTzxK9V/Y1O9ojQpnBcNvcfAogQVIvgXaYyFpzU6pRdr6X3NAqJOrrW4RqX5qEJd
sQG895OX2BvJcLbA//eBwrR61xd5UtK97zkkSBSOcNnCKk08DY78ADmDVmD6SPEf
2Iu6oyKE34jMu+lVV77MjZp0G3x5FblP/WP5yPuAgb0oiwh0YlAFy0tGG8hCyRcy
qWHi4rO2uUB1/WpS/l0tHX8jKYhmqA2BbDwm+xzJKBh83nrbiaa0ZL6cEV833Omd
fk9HWiN1aSaJMio71lB/A2sTF5HamqnszyTDTd289SbQ0CIUnyEP1ixMrZuIKSE/
yD9xcIk8VOMH+iSfbLZDVBvbqE2KZmxEU4fGpt3fWH5+9IDK3Cr8OhPVRXDAO0u+
RCbvwF2DL06SXrB6F53qogkB8X9lnxPz2GTp4DUOCfn2Nssl5+MfBs3TtH5fA0xI
HYD99SU1dhaF+AGo8XPLwRaG+7tQGh2Ykbv4QznS5YW5Z7jkmn+OsLVs+OyYuIbP
WcZ0yA60o8xBJgP+ZM7XWGcSPQ10zjH1kFsBbXmjenieq/++2LVaFW8dSjTaRQ18
fu2hFO3n7CpG9/ldNXRYh1luaa0F4t/xoZ2zfIherNhf/nuNiKeeawUP34fnbDFP
QBetoOFkqBnHy4DHIWNRnagl0EbTDHvF3G0TKcTA5jK8QYGlt3R9KlQtfLKPMUXZ
N2FUWCT61J4az8zN2OvzSXAe55+XNFZX12t3Mc7glFPDUMZGlBf5lAfrVeyxmgRL
j/JqqtyOVz+DenrHsQS/7DufBV+0YeeGOUiwPiihBOQCbiP+0QmUi8iSHRx2z8Tz
GbKzJxuxVOYPaJKrugH0GLYDwNcbRTJ/1HSa7JhZKaL8DOIFjTo+6ptIWmhr0Ris
dom9xfErE88DJKhJ+oCm32XxL/SCjJD7O4pmdD+aaWkAx9ZTCsbdTtuBl5HLu6a7
sqJIAgXv9ZBeYxmbMYVjVu2MrMjs9EmyVZF0HGVzNJy/RDyCzf+disstKT70OnZb
UNL9cPPzaB1XVuKF9s/dgjs7IqGdAtbz0hivsCkTkOxWFjMb7Xd1HVl2r5MPtQtE
Dv2Qacm3iBTGR7pgKLDLXCWltUD8DEa6e7EctjerDJfCyX5gLny2+2WSKs3I5N0c
VQBXx/flw5aKhrSv7csma9BfuMQeqWsV02CfwnH7fTngrTA2uwpJuPn8kVWkWqTY
Wj2xXvbnY3lhq3kMK9GziSrSt0SwL6JnfFkoHomZDTfLtgpHB1D/foTyA8KS+0Fv
oNjUhcF0/NJ0/YHkSxdEDMPesyxluRhdm8WhBid8qbT56lUcHfq82ESd6LMtl5nW
AuBIzn1ctNwh3oJcntrOeBlfwIWAvBEsiwLV8miqicPkbhwEzeYfFYvGg3D8ujQE
fSJMaAY9AbTnp0fODc7KgyaT9iwFUgXjklH2TMJic+jFPPR/4SLfzOghVkxkN/Q3
GExCOoxrPdPjUsi2M6x8Gx1Sjfap8iuOyf9ILEAs1WWvPMQKwfRCDICsIn1zP0vq
ugbW0iZQ8+TyPDVyInl/oq/XzmY4nhKo5HRjxQ/vayv9ge/oc3K9vFER2UUeuJ5y
ViKh+hj6Awbxaub96k25rZqScB/r6SbyUkgSpjLBCTz/nzDF0igBVw6VpnU5jNxy
k4IbS5tNH5/1XGycNY2Qwqzz/onqrM6VuwcUpyo2IVZcKp0ZpPq8ag4/djehUIb/
atSQsOakXB/CHDA7VJDJLKZx7gOF+VH9ohgYGLPR/rwTYLIMPMBrdO8vjQjF03QL
uBmw4I1yN4aYo96j5BSynjEliYSNnwddXd2fpdx2N4WH0fO0SGiqHP40N2DiL/vb
VybYEspemuaEJhvGZtTz7NCNUJYrD4g8zJMfr7NsfnZwUOik46eZmsF2zDjjWW74
zSRIJwDaxaSzsNtHaFIWTJGYU9SbejCZj2IT09sILaIuOqNG8JBsFWiC6EGeo7W0
du8LrY7PnDM8VKjqpy4T+KpMpnWi3F8EekEsOeEiLgUUKjwMDe+Kk2R3Qvq19f8j
/0A7aRuSAmQ3/l9kTJos1MWAd60+ZfvzOoHVJ5sDfRxEkkwVGDKR3GaaTfUTJjp0
kb5O3dZUlFWIXRKXnZAVC7gmrXiib1Z/Ulnbf7vsNWYWq2fOLIWqbYtrN1tp8Sru
UGlftfkStTkr7GKcwC3dIusaNGbezdWFsNQpqYyDh+qRRrNrubuXrs8duAtVqWQR
28kP8vAf/fCC/FIKyT9kPfgKPmmQblVB5MAQ+cnJbv8UXGzwIwSJa5jk7A6yk2Zp
WwInPV+eiD8k1mgIx0R0ejOHLqRAARkXbA/PSkeUjyD3b6/drcSoGTaQWaMb/ig8
ut7Neh1sE3dxSosGgEPHvKGG27DwEZg+MCL7N6rllz82nCmifwiPT03fZBMTVQ66
FXupaPWlQZJKYAM4lq3F3n0jOtuTIEBsXHmECx5ZhXZRIcedylEeB5cQWY55OYfm
CikPsPiCI1az3dbZQusAOvQRMeCwu2++WorwKQmC33Jlk5i8pDs/MQ2Bz+KzlyRu
UlysVhWTReMX6RuV95jebHEIHd1fdr//rvR0OlkZdP3AUmQxna/ZhMIxxyDXheZT
wp73sWtt6n5DQ7O7JyR0u7bxugi+OdtkFsCxFFp4YflgGw4AwmWjYxvSsLh92L0D
uOSXj5hbOQcQnBV6D4WTZFzF7YZm9oUw4yJwHhJkWoUoTmgiUSsrGIih3wy4oxgz
L3aY4hoztpKjsgEes6XBylbaZj/VyV433jwB2A4jlRM9q1CfLqWbeD+cFb6Vtz0A
9j+QtHMUQnbATG1GpNhYeib/gZlRkuM8chSNfmpdVqKdl5Suy1njZUUUuRjJajdU
asWPgV0eNALH0hgWli+xFJbMqIToIqJou47SJPLhphldXBT7RwE8KLdJlGFdhIzA
NgK84MSHQQlMqySF1+bQbhKevLhDiJeuopImZ4r41uVrmFCrti4tiAAU8coYP+Pn
C3Fy+FH7DsvJ7ggxJ8GMKy0yUEtIjWV51zStQhDh7jqQlDZTvAzhix3KCXAcPSSP
ETaNs7S6Yjqac1yrxHAwcrr0zljH3SCCRKCe9oJ6ML4MAFrWTYwVzXimpDU2rZhc
9/HiWMRrjp5D+3H3gnbjaunk0TJG3knja7Y2leE5eAPIKcXcVb70o6XFzpAjeRu4
G8htIO4h01qJa811iC9chMHnuYAPDb/1/ZXg+90YYZFHIh2h4zUvaZ2ZKXoubIHY
g24TvImGz8Cj1vAY9iwQY9MzsYjKXVRpspKLzwL8GQWvzjNWelDpoEIHhP6rjkwR
TfapLcVLyFJj96b9QQU5q2v8GxhYUCp4gR+YC7jiqVRxdCbgSnCD5PcJTOg0ivSF
4U50NSyrEx4+AGtbGk/pv1MTmiSarLGdm4RvA7HSQD8pd3b77TgRWtFniVGUVkAV
L2qdVlyUeHFK9zshz5fOnVJYGxIqO8mgrGYcE6Bu8ndQEZkSgWcdlNLOAZVx9g2p
f5Nc6DMPOAvBxo2qM51FeS3EKXK+/OY1q9DfYC4DDnlehWlDsxRswpbUh2mwLVuv
t/O8qFWL54MVdE9x/A7BwcWCzO7UUb429VIrsWhsQ1pUWtaf3gjcp8+hHCUPXw+u
9UnnK3dsbo3BvmtGT7F+UsfNXfVjuppOPCWwP5d27dOYhRDuZIxWjhJKCXKu3XQp
Z0FQyJR93/l1AYSZJPJwpLOsMm8fQtRtZ2JwiNarzD4SQwJCu99yz4ieou6LnskJ
+d9WB4oCuLdWIqSwyIJgzpPLwB/aQkrxWyjVok/vw2Mx52TJsPdQCpS6LMnxRxH5
LkjbRrVhmH1+0Vf0jUzrZVMdvZ/+kAe7/lULJs/SNcjijmfQwl4AXaiExEfQxWo/
c7viYl7O0PnvIL+2KQ0mzCPlT50TZpJeiZ6cZ1GiYkdtLtM7KJOLc6ZBUSL0BIXB
l6+RxS0rD806W9nVhNmdgriIzLDSmAepWevQkhceuOM=
`pragma protect end_protected
