// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ElEH3UNnak0E3Vt1IUIBZo4dwSKXOfq+WuLEFh94rKGjy4snhgMNt5MpojRE/HC1
2qb+vPbSSgGxPzC7K/6NpPiPS6gm3SwVFH3fr7vSWNGuIubTVKRL2Ik69uzrK/kw
mEXiVKt62scobwmksEEU52bgRSTAqVAbeVLAMt22Iqk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9776)
bUfVVtWDRcR8qOcSHuCT6GnGUq36Dz1ar5yDye2MitoCiNpOLkpP8ZxLR5hkEgRQ
+nH8k3lAayDxnjGWltoZjuTXZE7AxpNRW5OiUYcdexecWDg0UU7O3pZyx9mWe8fw
wtEBHaHTREKYGI2pHcO2YuQN7rjz3Wu5NF7u0ff6HIG/4e8MYtzNKYhFYT9102Kw
H3sIyV9hclQ3IsP2vYKcq8iOs4+iot2OU7DqhuhsVQn6bPIbOQL8K+ca4uaSSc/e
MQ/too4YsZ2g+ivcy060VQWFACVyV/67+13NAXV6zYxQXM6j1XLoPD/WfS/q9j8b
DndJ4nXAYSLCSw1bqlAQ7E6gvKl2qs8AtxIuY5Uh/yZDM947wmFuJtqp4nMPI5Lk
Xonl4NkOsdwwHVQ+VsSQyTaKyD7AF5+5+beagQcGRBLSrbiL46i53FF44j8S7bRr
swE3jAVhF1zBkpfxquPVdSH4CeiZ4mFpMgOgAidgZM5iV4qt7ndgEnEgmuKAT0V6
JpqpunlaRg7Oc7h/9+cQovBia/TB/RwU0hjNvNG3rFWiwoXVIMfCDYYv+wPsRRp0
mMSwFowweu4MauRk1CG6VS/NMOy9MSESNzHoEvvWcjMNXLh9e9vCeIGdMJzkvi2i
b7N+Es8PZ4d7LnFQNYAMLcsLoMOXuvUOCFyuBvNUq+XO1lX2qlM6eaZ2CDpm0HmZ
C92100IzAlnc88Diu3m7RkHdLUpzOOhfp4Sv3drCZbcqoE520E7AGLwxjpwlBreI
bTnXxbm2mDdzZTFM2bi3aWhcnrN01Ux0YQQ2sMBIMhh8xT3Zz7CXi3oHFLbeii0B
ERlMEFFg+Xcu97V7RNQTuy1zClCsHB4XfZ3upHEYIWiwn+ih2JH3ktD2H6h+dnah
GzS2vjEeTYJe6ible1KrNfWcanNqJKCOS2PFhkO4rar8TBYoRhi5S0FiPcGkL2sk
HSG2YAVCLRHGdrt8f0jxfW7FWQJC7jp4C6lJGA6bOtA3rpLKV1AB/Wjw9QcQqI6G
yTA8xB+XrkXynqT15HyLBRrFLUx7ETh6jg8Q5zbYcG7yrSXyoeiuA7VuCCI5cHOW
O6lU+zZ9bCGKatnXimChAyVDf27Vwx+TqtZZB7f3zXia8Lk91miNr0TkOcm2e2Yc
vvGcA2C7zGbYFz6kCz52u5nG7CZInScujSqQBW8CkoyagrbsKPuspIJhPlNNRdDx
6YsIR7owvcde3x2x3iDOvr9EKKHyo2JpdCwPmKvEPfgufvRChxm5kVYkEGM3V5wF
yh1+IGjL32fkEFeMq+3RSB2t1cWBuxBgykvSKtvBhHDFI1qDsOFAmcYwYDK3YIPr
dr+aEhkcFzRp59HeArsm1FAp35EE2xCtxjnbtjHr3pfIdJ5HkclVlHJxy4VUICd8
WUcWDKtJT2FU79KIKHLD1Z7VNjBnxfzepYjhUlCL4WRYq7kLVwn75jGy91Bx1rJZ
3khqdh3vcuMTQCM9ar18PCtgv8kS7GpRCmLO/gmt+7piOoNxPB5KF7AYkyWyMYYk
yQp5tdbO+p4tQyVLYvGIUwAnrcHQXVkUViqVDrd4J/IvdHJqnarfHo9KsBfMkWNa
k5tE6pAkHfzRm/OWJzPKh1yfGuVIljL821naevxEmV14wWP6ng6KFvcTOcqDf534
FzTpb5HgSiMuOgHwYo8JEWnfJysARxCeTLi/juJEOc6WJpQPYtgumOHn5JhYQ5Nk
mFqqOxZLtvPszGk8Xpy4erSR86MHcQTXu/4jqZy2YWMlp6juQJlRGQvejIua9rKM
osJrHpeyRh/b0TER10l7uJ+mIgNavaT/hDWK9pPU10oiS8/FOjfUjq/3INpuimcU
x5OyqKhR1IrEf+3U3bJRpOPsRNX50LcH+fvM/cf3wwu9DKmXC9JTpurwqYQdpAf7
clDoV0RriXEiomlyFmWD4IISlIwyFt3z/U+4fxfGG/AuWR9TGkwLCOvGBzM+ChVJ
BSx0PrEdaUV/eWHB5jmbTCh42kOVxR2jzAOgSsf0Duzm2VsMDOnC0TEqYKEcyIB9
pOyZ5j6A8mfJAB2lASjRdleKv4/lYmIijkQLX9q+Ih9dqYdCA4alIe4RPrOrRQjS
nUBWx96CS8rXNfgZjJndwa1TcwXR3U8BkMzcW0OHj/cLOFkLF99sE0L0BuhGVc6T
N287oEUR1vV+CpEvO1ee5m5O4pFYU2r5YF6dvVpGnpFTc6AXWZymMPsxxjuvFhJN
MZSLXxoMWvqN8+lR83BocM1Z/t4rsAy52ec7hF8UzW6kh76MlnHJF//XRzW/zlAP
9wuXVk+g2HH8qc//v+XZDUksJNW22u0F3eGvU52PRpBYb+5pNYV/uwJDetPHFaIz
oUand5pXHYVj333VhT+S3arUg7Ru13sfw7Zt/zHb0HeCzUXooX4isqQj2KSOiPH2
9vJaq0wvnxRCrbAjNxMfMO+Liv3i7evCgyJuo5/2eGduAYCWs9tdsyW3R0jxiw7+
vLjggUTEv6FaMShN4avcJk3ccSkVqny+xE3MgIF/8IgVrl1GvI16HN2lWaRlyMYN
U/osY+X55imywcBqZCeTgmO2VMxiDlrcOZbgHCwbX+AMgOSxbDm0QTe3Q0tf5Lmj
xbSUEGhAl6xmtIs2E88b/xRY6ihqwtuJE26Jh/A7jUpJED9GOnGej/jz9rq4qPWq
5JJH2kWFnmidnr9K3E409NlCfpbbdx1n9GSF2PaQAZvfTiHLlJEfpom5gqQ+t3ts
UNDs9Wd8UU4+5sXvLIT6iiqYg59+/haUCLi2RKkZkoTMzGh9eg616a5a50wWGTMD
x4d9CVqlaK6uZ3cp2FqeEBRpOk8wQMPdl3EIg+qfy3gpWCEvKmgwtnGT86mlMlCL
oNKJw44UX4OfWxahIuuU4DbEmfq5t9z2j3ULA1gbuNkqVo/2pozaOt/EmWNlAkKq
PUnHD6Amj0WsphTrjlQu3ik8+X9j7h1x6ZThRzspzXDRSKN/2b7JMVuR/1eaHvCA
dBH+sKYC3XcMxYGPuOIZDJrMfj9nhH15Jc2mZzhZYU5LslRX+g1l0w5DfeKBbxLn
hbdUQK+JlMVL23sJnMPA1LgKqJGNKwPYLdeJRIeq4/+KALt0m7DyzOVVDUMwalzS
Fx/GrpQU/BFvRIpmAvSWW05eXZzHw1F9UvaxTwbKDieTiZ/xf8oAcN3yLWxNIjIM
AkFB9yDEgLCrihPa3Krevj4GKTYf+mpoi9i6to303NJpcphxclfTpILhPnDVHUth
kgf8JCws0yaMaw0sr9NWPZ899y78ZAdnAXORXTAkdFfTP711RLrt0xitECLLkxRg
vTHn0QswtH12za89HoV00biR95T0AZd7p02ncxKmN/I4wiJR1Nx7oS3k3VAlfDnm
vKT3qmjH1kNaPoTw/n8j6Er25gjRVZi7rnuq3nJECp7buxor4j7iVH6SOdud9A3F
jwfeLDTW2zDqFF/lE52QSEgLYUq1nPq3fFThp7TYiMWYNtwmeuWaAe8LMN4jombA
e3FpVeihAKGiWS/XuBo8Wf/CwTo0VXH4HnbCOv9dSb1LZutWFdNtER/tTMT/FYYq
VjJw2c8Eja/ETADPEZnwRGpXZrqqhgUwPAbVYhlx6WWogXZkn+JUzbZRuHBZmW+L
0QqGInkW0uMIcolNjll/8KnXWrfi8xPT8tLMDx944/94wHK/agdZYUNUr6a2gG+u
AkPS/a+/7nG1/tiBfHb5ZLFXP4wQblUH0YJFve7K16si+qDZ7PiqH1sCDAFf9SFd
na/E+WS36mBcOYz2Vmw/JhVgrnu84GPwmkpSb+U6QVpLvUa4NIZJGopd4UluFCWy
WqYIJQUW5s0wyWgbNCUBrKaYf6DX9AHXKrfVNmBCsdwP4qzrcvKp4snL7Bx8Kmg6
9dv/59uV24DKfCq6LnRDTrPZIKwZ+SE7UYHrdDk475tg1C7zGODIgnHMeoAaXZ/q
hPZS6QoP2OGPPeCghkG5x3s4GUzMs68+RfWBQIOvX1AYQUPYi+d03zYZtWZykrsR
fLyW83L7w0Y/fIZ72yLQM+vL08ERCBjjjxLuEVWLg8SasQSGyzg+SB9Yd95fOUv/
7kccBARK47MLl2Qf6kaiXRxSXQ9+/EfSh+MfXb1Rn15DxMi99+Ipot2GnqCJ0wYb
wqBgT2YYVi0JLhcggJ9DAIA9m9IEqfilV2pDtjnpGhRg0BhZtBR+47Jq105eqI/h
dcwQB9wf3DHe0+CvfYcKBWGInz4Sf78nSRnYe2IrR/GoVmH0BdqbmJrVljj+lTMq
iMii7hEkIcmiF5FJvDMmRl0BHoUI4h0ka3WEw+JVhxL9zmoP+3qy+/ePfIsR/pqW
pxLxlFGe7vNeOn9UYLlNRK3YAGo2jvMpiX3M2ePQRm5wjW+ktcgZt1P29MHzwQWZ
l3TkoH/ZsjgGjUpb27B/J/YOhtrO+hR5lbT80njSOKMCypIDli+zQW7P1VlVvyAF
UQ57A8X8LG9bORUG0sR/eGIB8UEB3vYydMdNOm25iKbC4VYS8ftP5juZi37RB40S
RV3/XVG3jyw6iJ/HDWPdVgSM9EaKRctf7qH8dMgGnArHbHKGAA7r8RfwB+7o9Zyh
bJCFs1iSUlInkT8kH1Rg/656NM+9dPgY3cspGm3OGd1BVvsshUZrtapC0tfagR1r
SQC44qkzsU40BHTPKp7dao0kjk7i5kTffujl/uIYBwtdbHDBfAPMr4iiKYbTU0JE
d+99hg5hDC/XLnKkvCZTLL1QWB+NVCh25uKdCOk2mjI2FBg7AByyr+8C7t/g6/6h
ecKTBSAPQbKGb5dVQVf0vpPpODWkOEcByYj6AsSSPw7klVUv5eUciTjj6PazgC2f
icbxeaA5XDcuXruaBsTtIkiyNYMuSaKtoYYOsLRqLuUY7hgCm9jpzDG5n8Kb9q2e
84eHyOMpIbF3FCLrODvPJqNprKZ/wrO9NUpIvwsq7jsdLyAEzoMs7dEVgQtgFFtH
lfSJGyiRPwUqevcWL91K5CBKH5u97CYD4C/G2kaTCWRrpJ8uqHs3LQby+2CnB+Xr
gZE1+qyYoiIGnuUzK4S9qtj4Gy5tmZGTHMu2iscT52fWQMZCd34EmyuYEhRA7J5O
MXe0g2fyDcQyiZdXz1p2sGCUfkmvXXhxvoV/m3CPlVjwpoTvKM/ze4EDTvOU4EI3
tHahvOAB6kZX4rjRGwrWYBfvKAdARO4zogzAYadlxjWAoHy6UZoJEVCHjnxS7EHo
btDWAYAGCj//c5Sg7OLGMYFMGNkvOtsdEw2upI6JaTrYSoczucY764a3qLVCIEEm
4EviWt0t4MDrCfy2BmTl7/hajwaY+HpM22jtvhjDNZKQZkCdT5fw7I4uW5gniwv6
gMOORUaIqrwaFcFDZGBzXczULbYZMRxI9fRm/W7W7FCtAqOnxwNKXysY5WO0H0pK
9eTSUSsNri42qZI97BmtQezB0fqa4X5FvzLk6B8oiPOtey+BpRZh3sO96RnzLHcb
rYFRoJK8zlOdGY+c+a06QkQ1gyNowU511ZYZakp0gBM8FtSYrqJu+FJHN+7QJB/R
Oz2CM+8NX41lxw3Led8DfboCNOOMd9Ro6VhJj8YnN4Lbac9oGP4RSy2zlFrTlxZo
5t7mTgRbj2TQV9t1d8vktCJQ7GzX0p0v8msAbXCPv7jou48OcliPVEVs/2MnYR66
7U1OZP9UzP/73rVTUZDufLjSJQZMfUduMzk5MV1vRZsT/bUJ1Ln9zdwe11MZqndY
puKlkMejLWzRdf+7wLGYj9YeFcjQaiEKq/LGbQTAPpNfBVGo/zh1xx5/q2IAYRtp
e1mIuZxianRSMQcQ8v274XFUPrm52Ty/N7cQQ4apl7+j/tJsTqq1ODaAfiQsEsrj
4Ev+sS6vzCWYb02gjM2U7l/xPtRXtipgAfrsOWE/YtFZBX7JgVDG80V6Mf6f6Zk4
hDyLPpl2EbCf3oFmTKwYrRi8nO5tJyQ3S+loP4wP+pheJurHyDdvilI3UIG7DcXT
+ypEUSUbuLrlTxeZtTJsv7neZ/cG6LvYpHebF3ikASIanE2FBRRqa506iJn7M3lx
FqUn0dSo989fPi5laDMymJ5aEJxRitXTD290jfLHeO1SKWByosNfamFkOlQmwbwn
FG1s88KViuW4aGihuIySeHIQR18MyPpF5o8WEjmk8UtcPG92orfkcL+5EGY3OO3S
/1ZJaJJJ09vFbORmpLc8+/3a5ou9LbthB+Eka/Ki36S7+H5vY7oViilKe0izSiIp
wzO3zYEVIYjXMQ88LvoYPT0AEWiA243rbj4t7Btg4pN+xv2S5rIKFx/LUzOWlbjO
PAEjbgrtt43SGVoZtuuBwlMhg7GXH2SskRvwB9LcGcBK2y4+4xq2saRkHAlvG7s0
7SCcjYzsqiRsqZikcKEvU+rD/V0SIIMHspRWX1slLvrp1NzIHFkOdP5zkpPdIwkB
bwr1zlaz6fZ6671hCJAhIniI3+dPb/njv8UFl5keQi+h69xpHXo3uRts5XkeY5UL
dPoxOJoky7Mf43aNhfMabeKbUVYhVkEC+A7FWBpi3t7siTboHi57vd2AsYxWtuFt
aP73GuEaPg/nNSzJyOUONvN5LtYL0qLfBEFUyVlBUMII2aTutEPaJfjzthr11VGd
vPlofdJOVD/iEvM51pPZUAFVLXpQGZarIZFHEqO1ILzZDzzbv49Dg+KRXyo0xVhp
TRBcWMwnE4fM03v7CplkdpUZ05AEYfVx7GeE5u7EdPBg3ybE8me84gp4u0JOz/gW
UI+2zZTfaZPCSt7U3k6reBx7NM9zZX6xAxeB1lnMbXFq0aboIeVyjd/nOlVWTFQG
m4JqKt2pF0A9rbL/hFJQD+vTDkY2ClNIaUUEzEoTBS+U84XnWJTobnk/cAGyvUmM
qdhGi3POhXMV951JyL0xM8ORGdurkBRZqmikG8338AKkWwRQAYDFa1YsFW3WsHer
N5ur7OA2LgSBqsqNymzLhy3ZX8nWcNnujMvE3EZ++u81ai3DSgTCf3UvptB+dkEG
/bolIJL2uSQmtWeWoBkyYHIzmJqS5uBSGKWhE9VvVkciUgAof3d4bmygc2leLpcw
H+g0smjeGgxf4vbXiPcDm198By3cF0qpp/TCnpGAUaBz3PZTBuVSZUESdZhEAjS5
Id0R2zYwmSW1qBX8qgCETgXIdvZD/RlU26d98Jb/pb79KHs70HGUnWcp7h3ZLVP5
g3qqwWCl1dZRpKq9K9UR/wN1EB/SZ/1oSozDZ8A0BlYWWJq3hHVT+7au6O71bp6x
v9ykq1fA5pmCepR+5Ue8GtlEc6Ok4fthbMddUfB39kg1TgbxNabltQmHzWRuOboY
uM7NRZRSBkOWYudv8t8kMxvSPMY5T4eIfqFuvPTNIgtdnJCRoaULTNM1oTV9oC+a
uy/rYClGKYWCGdQMtKuPHudEIXB64fnDRU9BEESb52LEgKfd+9NKmfpIMoZDPlNH
5QhIagfoiEM4IueeD9EQf4Yf1q4f0UDxBmX6oc0vfVFZeiC4FMUrFAZItwRI+Is8
OyA8sR6gFsu7CyV6+YFCpBqgzoFmbTpvAUlWch7i5Q1Rn+DAkewwFD2DPLDmkU/0
hd0D3dBvA8fmlTenfSyw3U30VuYPB4OyzNrhPGNnEeLxO2rrWDtTXbaLHj81LDu0
zoWrkJK5A9rKs0ZsoatBUt+taUsq80XGrhXyV2y3GsbuXaX4EkD6fa0u8iAwDrlr
rmjwtgxoE4IXSVcncHwgMNhcw5ECDDfe5y6Qqm8QenTnrsEaMDiOTtAWHWh3Y1KK
BGWdfbUv3POqFeXL7x4mWyMdLRLbJsukjfEsX1sRY1tFDQVwSPqNl8sjrnMojN7C
xdNeaMw6hgZVRd416vopz4+Spk4Uu7yYdn/H7w/Y6qr7F3bfGzRgQGq1YszhcrPf
XUANBsItp99al7LHHBClzKw0PfjCwi/NiHwgXaZ0SiJHnlyED468XfJoKav/EOV+
cKtplLGb+8xnYXu1AP2ozRoS8Jjb14jbQUx9WlD57vdL8tdLtlnaYMRPfTwGtQHs
YZhWjZdt/TfP+6xod2qZfpIrjaCC7bmnaCJ8pDr5j9JbRzqEX441+TfjkmV0e/Vd
2iluabZvHy85BYFBYGGMnaBEGDe2EGnrMnYV7oASuXXQ1pDU1lHQFpwKEeK2LWhs
zJAdl+Jnf/uSYoPehBEt1lY/jvEBCJ55KqtYKG8ArVeDTNBmz31oHTSrAe4vXcWQ
w0MyormcYwU/Kdb36EmM2a9quEwuOyifaLlNcIkp7aPUgWfJy3viYg/0oIZkwq5W
T8TsMS6C4zgmv/RrlME3VLDy6BP9Vjo4RBQDKHAJ3cgfW8EJnKpzG91+NcGrsaMU
SdNbGDt/HjI/stsd32rhyDCj9UP9JNwVbE5cfCseG/+CNTLqF9iIhSTQfsiTVfq0
eBBDF1O/BnO23HslU4IyJU1ZFsSC/kgogJQHTHt2Cz062pfdgTOe5fWiVHUnB4xA
BWs9ZWkH7j7IYukZmgwOwIHf+gGJENsPjrZn4BmucAPwIeZT8qU6+nrMnvZnMuvm
luAE45RnD7erAUx+idUONrSVdMcDx2UPZLALUWlCZexwqRDOB8DZBJdddp4kdGIR
bd0YZ0ejXSFheEsEwgB96Izb2uVVUR0MHai2aSPLD41Obb8G2ihFs6KwXwfgOzGz
mp1bqbc9n0xcccvBwBfkJ7SsaTwqFeLEzVCal1zVchh7xpfVKuKIyG3NLf32efEi
Z3YZJWixBkRI+Cmh9Jik2WaV4pKbHXUjqZCyzh3NuWSCxDu/dvtj1LWQyDAhcH0Z
D8gncc6qMqsUO/9qHvGUMKCOHtAMk4jnUBJeLXJmFbVX7Qlx1eJs+iICEK5MlTK1
ZKzpUAARyMQY0n3pmKzHR9hts7eErpR5oDK5gG7opYvrbdaTLrIh5xE1VQitGSx6
Sd9fYcyb9ZC1/jpHZUBJUE89hX9QM3RdBRNUyYvoQmDOhZuboiZGt3IntbtzAkQg
JL400klMpMhQoCRBvVHrgpWWq6IdvM65hWupTyPqPY6LoZEdsiv11K+erI3ieLxq
cMfOKv8KtT9pA0OVoHSLi9/iUE71CvR9VO/6xDIzWj/LnlkjOlVcyHYuKJM5qZFV
MEyld4Hcnn4zOO2KY3kFUPSoZp1ibNfPAgcWXsQz8aoS6BjRSCtF/sP2UW1yfoC6
sTgmE29a/yvIvrKJW52lAY2nyn8Y8j3cmK3AtYM5S5FoEUceqhmm8hkdYMaKyEZf
jMS/fa3L8RcX5w9u63T+HxYOCfQhULiS35fDUKxzWBaJGVD8F9kHHYcYplBEvfjr
GOoLIhR3XebE0fnGHoPr2UqnNwMoXXI20ElmIfj03+4k5S2+26/NwCjupIiB8tcc
G9QtaiIbXNcec+2Ej88F2LFiXf1ApBLwUGDZEZjENPhsTkBrap1FIjnGtM9vFymV
LzjDvZ2Hyzq3PWLehhwjWjb8pBezbqimiIVWlNOR/bnUKg4mgekZY0ZpcYYOSgjr
NzSe4oo9WNcip+KYZxDd4conkYLiKUJ36d10iTCEpDun4L1fxNUeJOIfxQTSn25i
rR/wy7WkSCiSkNe18mvOxIbB9Nq+wuqHHzu2dKizdXCDOkD0j6r/SgRnBURTt6nG
6c8Eb5Sve9uukJPH386aHtfB+X3PEfh5GJMEgH0m2VYfsoSnyROCQNbr99C/Xz5k
JZk3iKPVPLGKqCIEO0J0nO4GfAeJHUr8/oVQgGRmAKZpqiurDrjtjpYtGqaXyC6I
/fwZ2jPDdWLQGu5urHTJGiEqsAECZkNyq+WAoQnjrlZtWmW10mmQFv3VNO5bM85w
SFSuUjTGELsdqK2QbOEUvz5gm0mMNVTKj+FlUkBdn4uNPy2rvE+8dUWb/DTIupZM
/Zp1Or+nLQ6UDzHmZ+A8aeY9htxNSIyAKxugVNVfhKguXRLf5Z5pRyUmIhT+dePC
IqIXkdnFJcBbNglJrxbT4z4maVRUJGaF9EOgpPasIRdBeHBFGNB/MP6GeTpGM6e/
AJRwq1QatXXK7/W+38y179mqVyUg6hrtmQLY6B2eIR6YSJXtg4JitIDw0HBOmwNg
vZEupSD4W2jVOnEI67CeL6Y66O43OzG1RCWeVeE3yVPL4RDRphDXS2HWDXynuBRN
WxR0uH/J6lecv/ZOd82C8LeEGm2I1m9wWp/MoKkbldyciTzir61JFQpPK+mutNdS
Fg9zoDa8FlNI+NVRdUTJhyJeOBj25ioMgRa8ROF97Tz7zwnxzVNSGLGd30xqhcYO
tixvm7rAMIROwZ8L6H/hOGceg9mR65TEuN5e3MZYhMFQfWs8bMFr4BxergFDOwu3
M5ggL3HfBmeRTJxPgqq+CS0Hw0Uv89dunTDIdHXqKTCms3LUii51yN+S1EajZcTJ
wi6A6yrimJvgt2WUA+LryPxTLX1Jl9x4BcDlUILMRg0jkACoSKwv4UubYxX9Gbcc
TlzraYYl3A6DwK7Zs+GT8fGFc2Sx9lxkcZQti4xVqJfwjy/UKpn9iVm5G/b71tVG
DOuWOXFZhEw3LgQiWZOJdf36/+RnQ/G0al+naJxrPuclEVt2vFt1wcVWiappZ7Nl
xED4SgpMnALjFVx3ULPvEcnqTKhIZl6oi1t0308zLjif/gVXpev8meJlKPudQ8xA
KzobCxhcE68Pylg/XbJfpuYBE7zSXr0qhAhwJ2e1B2Cmsgmcj7MlCwnFBZNH2eki
G6QRf12sEBKuaH5UCNexXR4eFjDJfl69ykdWiKayuqK0QJCyMIpDLv3Y8KexsPY/
EPjScmnoFgBui5BOdcpCrRjCdT03e90J7p6JoiJ82HsPazEqYOZfaxGitn3Indtq
GQrrQi1P2LwQs77FQ8wu3h/yCe1uqPQuXfFGNRznVr39D51RLghQnlfqEHmcZOdq
lkX2sTikKlXW9cCBHuqKRIba5kK0fmftVdPWTYCiXCZmCgMtZOKlrf7mEOc29rDS
oNESJ699hbLb0Z+QSGPVax+rYIUlcj+1uoqcw9/+BgoWHCfB+LlJ5YquSgzxV12o
GvOYHkGo5MW5HmQpAn+eZVAilXffNQBfg6yruVq1SCxUWr1R3Pqly0eCwwWqWDFc
zUH3Shf4C+6pDMP/sgK67jOkCt7phMap1MWjtjxeiMdeJnx3J7C4jQ6McInjOwfQ
Uj5/5f6TnKEd61/tY6tYx3LNzpv0uX09MceahPIng5W89qak1VG5Kfqe3jgiq6So
5vx9ZaWaaTvknFWIAK/z8SmTBQF5GjaqpQ8sx7HDSvhTgLEjyEfx3H29/htGB8ub
jo4L4ZyglC97PG9Hpcypm6B3NTAhQOug7H5ukrQELg7jSTlg+K3D/xJnYLitp0xc
t9VC/e+IbefLNd6o6lAKjzxNRs8v72cr4UoHkVH4Gx4fe0eynUmdwMISGyyW+hT3
jKvXVRgQQWjKi+iojvAjzk77l7hP+4rW4JC6VDSsE4XS37Vp4Hv5yFyT1JWGrqps
bOfY6e+ULd33Yj0TZJ4XUsSpzf3yYdFUK38/O880ENb/edmaoqR1XRj9E2Lpyldi
SONgEsugBoxCtId40W+fiHwf0IUUVpRe86Xtm8noVMpSrYoYPmaKNVsK8SjXFgvr
YKeePiplPo/8fHRSXzExitDABaKPSMZSZ5OvwFNlTeSENTZAqmY8nTM0UExdbVYu
xz/56IgcQcs2JWsfvS1CAoyQITaVM5av63iKYH3VQjLxLWQm/Of1eEtOH+EVG3Kb
Iv2Ynz6IN2ZMO+QGZJeWm4/KoKqye9i95Zm1oC8z9SAUu8U67RwHKU4WFHRJA0m9
UaXMDkvqNxlauIJK8FiUyo92QuWs0f2jq/aNxAvtdVJPCQ50UVvBaqLSG7jI/lU7
WTiTMFsyMRvg/c0F22MUjty2xbRI1MvyGe4OUdRIc9bh6ztmN0eZvQDAr2BfSXLn
yeaEzSTld+RQY44wN/Pu7OmDGXYvujXjttYafpO+Za5GzeDGsdBJht4NOH4BfDFP
w8ILdoEGZqh98Dyqs/TPL0DqQqWoXWgDASp+JqwoKlgJ6O7m4pct5CvsOiY0V5Vd
o9wuEpvlwCcrzECjwmiUZw0cTj0hjHUYiN2vdi3yAzZd9XLIMzUd8SEWjYFjE+ON
1YdKPwiUKmtlBd4jx31filCGr/Kih8se+6egZ874Gtj5DO8UKQck5ySW9Olq2jhM
H56D6AeDmyRzwAhZCUDdUZOMR4IgrLz6asaRh9B2xvkLwthPmTxZwqsTn5ItFoiw
OD7WbyMM9vJijSfOrLybiTzgoiwYqhjdG/8tN6F8QZALrv22wOnxY1/Z5ILnwrKO
6kijKgQyejErAxTkGepv/CmZXqCjRn8Bt3sO8Ok/4+kiaYjnv+cuOgAqg3bUn6bU
9/SG6PgLlHhur1OOtDY1gQWtMcA0Ykd7l9GkcXc0H9oLqsLS7957Ia8eLifHsjzK
aiHoJGnz1VtSsn67G/nT3zbdayEBUyAorJNrsPOElELSXC+uxityx3vUP6BIw121
GdaaMQpzcpxv1r1qIidgnqHQIgt2K5p36BLnJlUWrWEdDFjZp+8GTdzwnW92ZvTl
gCNpaVRoy08Lh6ymLjmPxFBAvbgvNMLAhtEMor68UnfD4Dn0bvi6Gqwb2t58OUYZ
fZjx7sL9H38hh1Hr7R8okqCiX97OkHOPiVuUZCefQhXO8kIg7SnmD7jOo6bv9aW7
VMD/96SEXGljJwQrArfCH6MH5ul4I+d8tWzM8WlOxyojgWg8L7/8CSMHZmLOEPdh
5pobJxJB/wgB/LITFvT5bc1Cb62W2s0qr0GX6LblQOqs++7u5tk0YAFTHbK1hxfp
E9darPVvXi7KAjfP/hUmblWUIJ9GVIB9qY1m7/2tViiMDXSRLmUzzifvlIJ5KpJH
gvFx/1M0T+Q8ctnfY4EgBjYi65SKoTtQyLyyhqSSkmSSijYtiMxTJjsS4wwo8yTf
s5/MrzXjJ6JM6WfnzZXMudufXK3QtnRpWetkBr2EVjQ=
`pragma protect end_protected
