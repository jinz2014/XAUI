// megafunction wizard: %XAUI PHY v14.1%
// GENERATION: XML
// xaui_phy.v

// Generated using ACDS version 14.1 186 at 2015.04.07.16:24:55

`timescale 1 ps / 1 ps
module xaui_phy (
		input  wire         pll_ref_clk,          //         pll_ref_clk.clk
		input  wire         xgmii_tx_clk,         //        xgmii_tx_clk.clk
		output wire         xgmii_rx_clk,         //        xgmii_rx_clk.clk
		output wire [71:0]  xgmii_rx_dc,          //         xgmii_rx_dc.data
		input  wire [71:0]  xgmii_tx_dc,          //         xgmii_tx_dc.data
		input  wire [3:0]   xaui_rx_serial_data,  // xaui_rx_serial_data.export
		output wire [3:0]   xaui_tx_serial_data,  // xaui_tx_serial_data.export
		output wire         rx_ready,             //            rx_ready.export
		output wire         tx_ready,             //            tx_ready.export
		input  wire         phy_mgmt_clk,         //        phy_mgmt_clk.clk
		input  wire         phy_mgmt_clk_reset,   //  phy_mgmt_clk_reset.reset
		input  wire [8:0]   phy_mgmt_address,     //            phy_mgmt.address
		input  wire         phy_mgmt_read,        //                    .read
		output wire [31:0]  phy_mgmt_readdata,    //                    .readdata
		input  wire         phy_mgmt_write,       //                    .write
		input  wire [31:0]  phy_mgmt_writedata,   //                    .writedata
		output wire         phy_mgmt_waitrequest, //                    .waitrequest
		output wire         rx_channelaligned,    //   rx_channelaligned.data
		output wire [7:0]   rx_syncstatus,        //       rx_syncstatus.data
		output wire [7:0]   rx_disperr,           //          rx_disperr.data
		output wire [7:0]   rx_errdetect,         //        rx_errdetect.data
		output wire [367:0] reconfig_from_xcvr,   //  reconfig_from_xcvr.data
		input  wire [559:0] reconfig_to_xcvr      //    reconfig_to_xcvr.data
	);

	altera_xcvr_xaui #(
		.device_family                ("Stratix V"),
		.starting_channel_number      (0),
		.interface_type               ("Soft XAUI"),
		.data_rate                    ("3125 Mbps"),
		.xaui_pll_type                ("ATX"),
		.BASE_DATA_RATE               ("3125 Mbps"),
		.en_synce_support             (0),
		.use_control_and_status_ports (1),
		.external_pma_ctrl_reconf     (0),
		.recovered_clk_out            (0),
		.number_of_interfaces         (1),
		.reconfig_interfaces          (8),
		.use_rx_rate_match            (0),
		.tx_termination               ("OCT_100_OHMS"),
		.tx_vod_selection             (4),
		.tx_preemp_pretap             (0),
		.tx_preemp_pretap_inv         ("false"),
		.tx_preemp_tap_1              (0),
		.tx_preemp_tap_2              (0),
		.tx_preemp_tap_2_inv          ("false"),
		.rx_common_mode               ("0.82v"),
		.rx_termination               ("OCT_100_OHMS"),
		.rx_eq_dc_gain                (0),
		.rx_eq_ctrl                   (0),
		.pll_external_enable          (0),
		.en_dual_fifo                 (0),
		.mgmt_clk_in_mhz              (150)
	) xaui_phy_inst (
		.pll_ref_clk              (pll_ref_clk),                          //         pll_ref_clk.clk
		.xgmii_tx_clk             (xgmii_tx_clk),                         //        xgmii_tx_clk.clk
		.xgmii_rx_clk             (xgmii_rx_clk),                         //        xgmii_rx_clk.clk
		.xgmii_rx_dc              (xgmii_rx_dc),                          //         xgmii_rx_dc.data
		.xgmii_tx_dc              (xgmii_tx_dc),                          //         xgmii_tx_dc.data
		.xaui_rx_serial_data      (xaui_rx_serial_data),                  // xaui_rx_serial_data.export
		.xaui_tx_serial_data      (xaui_tx_serial_data),                  // xaui_tx_serial_data.export
		.rx_ready                 (rx_ready),                             //            rx_ready.export
		.tx_ready                 (tx_ready),                             //            tx_ready.export
		.phy_mgmt_clk             (phy_mgmt_clk),                         //        phy_mgmt_clk.clk
		.phy_mgmt_clk_reset       (phy_mgmt_clk_reset),                   //  phy_mgmt_clk_reset.reset
		.phy_mgmt_address         (phy_mgmt_address),                     //            phy_mgmt.address
		.phy_mgmt_read            (phy_mgmt_read),                        //                    .read
		.phy_mgmt_readdata        (phy_mgmt_readdata),                    //                    .readdata
		.phy_mgmt_write           (phy_mgmt_write),                       //                    .write
		.phy_mgmt_writedata       (phy_mgmt_writedata),                   //                    .writedata
		.phy_mgmt_waitrequest     (phy_mgmt_waitrequest),                 //                    .waitrequest
		.rx_channelaligned        (rx_channelaligned),                    //   rx_channelaligned.data
		.rx_syncstatus            (rx_syncstatus),                        //       rx_syncstatus.data
		.rx_disperr               (rx_disperr),                           //          rx_disperr.data
		.rx_errdetect             (rx_errdetect),                         //        rx_errdetect.data
		.reconfig_from_xcvr       (reconfig_from_xcvr),                   //  reconfig_from_xcvr.data
		.reconfig_to_xcvr         (reconfig_to_xcvr),                     //    reconfig_to_xcvr.data
		.rx_recovered_clk         (),                                     //         (terminated)
		.tx_clk312_5              (),                                     //         (terminated)
		.rx_digitalreset          (1'b0),                                 //         (terminated)
		.tx_digitalreset          (1'b0),                                 //         (terminated)
		.rx_analogreset           (1'b0),                                 //         (terminated)
		.rx_invpolarity           (4'b0000),                              //         (terminated)
		.rx_set_locktodata        (4'b0000),                              //         (terminated)
		.rx_set_locktoref         (4'b0000),                              //         (terminated)
		.rx_seriallpbken          (4'b0000),                              //         (terminated)
		.tx_invpolarity           (4'b0000),                              //         (terminated)
		.rx_is_lockedtodata       (),                                     //         (terminated)
		.rx_phase_comp_fifo_error (),                                     //         (terminated)
		.rx_is_lockedtoref        (),                                     //         (terminated)
		.rx_rlv                   (),                                     //         (terminated)
		.rx_rmfifoempty           (),                                     //         (terminated)
		.rx_rmfifofull            (),                                     //         (terminated)
		.tx_phase_comp_fifo_error (),                                     //         (terminated)
		.rx_patterndetect         (),                                     //         (terminated)
		.rx_rmfifodatadeleted     (),                                     //         (terminated)
		.rx_rmfifodatainserted    (),                                     //         (terminated)
		.rx_runningdisp           (),                                     //         (terminated)
		.cal_blk_powerdown        (1'b0),                                 //         (terminated)
		.pll_powerdown            (1'b0),                                 //         (terminated)
		.gxb_powerdown            (1'b0),                                 //         (terminated)
		.pll_locked               (),                                     //         (terminated)
		.cdr_ref_clk              (1'b0),                                 //         (terminated)
		.pll_locked_i             (1'b0),                                 //         (terminated)
		.ext_pll_clk              (4'b0000),                              //         (terminated)
		.reconfig_clk             (1'b0),                                 //         (terminated)
		.reconfig_reset           (1'b0),                                 //         (terminated)
		.reconfig_address         (12'b000000000000),                     //         (terminated)
		.reconfig_read            (1'b0),                                 //         (terminated)
		.reconfig_write           (1'b0),                                 //         (terminated)
		.reconfig_writedata       (32'b00000000000000000000000000000000), //         (terminated)
		.reconfig_readdata        (),                                     //         (terminated)
		.reconfig_waitrequest     (),                                     //         (terminated)
		.tx_bonding_clocks        (6'b000000),                            //         (terminated)
		.pll_powerdown_o          (),                                     //         (terminated)
		.pll_cal_busy_i           (1'b0),                                 //         (terminated)
		.xgmii_rx_inclk           (1'b0)                                  //         (terminated)
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2015 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_xcvr_xaui" version="14.1" >
// Retrieval info: 	<generic name="device_family" value="Stratix V" />
// Retrieval info: 	<generic name="starting_channel_number" value="0" />
// Retrieval info: 	<generic name="interface_type" value="Soft XAUI" />
// Retrieval info: 	<generic name="soft_xaui_cfg" value="Only Soft XAUI is supported for this device." />
// Retrieval info: 	<generic name="hard_xaui_cfg" value="Only Hard XAUI is supported for this device." />
// Retrieval info: 	<generic name="gui_pll_type" value="ATX" />
// Retrieval info: 	<generic name="GUI_BASE_DATA_RATE" value="" />
// Retrieval info: 	<generic name="en_synce_support" value="0" />
// Retrieval info: 	<generic name="use_control_and_status_ports" value="1" />
// Retrieval info: 	<generic name="external_pma_ctrl_reconf" value="0" />
// Retrieval info: 	<generic name="dyn_reconf" value="0" />
// Retrieval info: 	<generic name="recovered_clk_out" value="0" />
// Retrieval info: 	<generic name="number_of_interfaces" value="1" />
// Retrieval info: 	<generic name="use_rx_rate_match" value="0" />
// Retrieval info: 	<generic name="tx_termination" value="OCT_100_OHMS" />
// Retrieval info: 	<generic name="tx_vod_selection" value="4" />
// Retrieval info: 	<generic name="tx_preemp_pretap" value="0" />
// Retrieval info: 	<generic name="tx_preemp_pretap_inv" value="false" />
// Retrieval info: 	<generic name="tx_preemp_tap_1" value="0" />
// Retrieval info: 	<generic name="tx_preemp_tap_2" value="0" />
// Retrieval info: 	<generic name="tx_preemp_tap_2_inv" value="false" />
// Retrieval info: 	<generic name="rx_common_mode" value="0.82v" />
// Retrieval info: 	<generic name="rx_termination" value="OCT_100_OHMS" />
// Retrieval info: 	<generic name="rx_eq_dc_gain" value="0" />
// Retrieval info: 	<generic name="rx_eq_ctrl" value="0" />
// Retrieval info: 	<generic name="pll_external_enable" value="0" />
// Retrieval info: 	<generic name="en_dual_fifo" value="0" />
// Retrieval info: 	<generic name="mgmt_clk_in_hz" value="150000000" />
// Retrieval info: 	<generic name="part_trait_bd" value="" />
// Retrieval info: </instance>
// IPFS_FILES : xaui_phy.vo
// RELATED_FILES: xaui_phy.v, altera_xcvr_functions.sv, alt_pma_functions.sv, altera_xcvr_xaui.sv, hxaui_csr_h.sv, hxaui_csr.sv, alt_xcvr_mgmt2dec_phyreconfig.sv, alt_xcvr_mgmt2dec_xaui.sv, alt_pma_controller_tgx.v, alt_reset_ctrl_lego.sv, alt_reset_ctrl_tgx_cdrauto.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, altera_xcvr_reset_control.sv, alt_xcvr_reset_counter.sv, alt_soft_xaui_pcs.v, alt_soft_xaui_reset.v, alt_soft_xaui_rx.v, alt_soft_xaui_rx_8b10b_dec.v, alt_soft_xaui_rx_channel_synch.v, alt_soft_xaui_rx_deskew.v, alt_soft_xaui_rx_deskew_channel.v, alt_soft_xaui_rx_deskew_ram.v, altera_soft_xaui_rx_deskew_ram.v, alt_soft_xaui_rx_invalid_code_det.v, alt_soft_xaui_rx_parity.v, alt_soft_xaui_rx_parity_4b.v, alt_soft_xaui_rx_parity_6b.v, alt_soft_xaui_rx_rate_match.v, alt_soft_xaui_rx_rate_match_ram.v, alt_soft_xaui_rx_rl_chk_6g.v, alt_soft_xaui_rx_sm.v, alt_soft_xaui_tx.v, alt_soft_xaui_tx_8b10b_enc.v, alt_soft_xaui_tx_idle_conv.v, l_modules.v, serdes_4_unit_lc_siv.v, serdes_4_unit_siv.v, serdes_4unit.v, sxaui.v, sv_xcvr_xaui.sv, sv_xcvr_low_latency_phy_nr.sv, sv_pcs.sv, sv_pcs_ch.sv, sv_pma.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_rx_pma.sv, sv_tx_pma.sv, sv_tx_pma_ch.sv, sv_xcvr_h.sv, sv_xcvr_avmm_csr.sv, sv_xcvr_avmm_dcd.sv, sv_xcvr_avmm.sv, sv_xcvr_data_adapter.sv, sv_xcvr_native.sv, sv_xcvr_plls.sv, sv_hssi_10g_rx_pcs_rbc.sv, sv_hssi_10g_tx_pcs_rbc.sv, sv_hssi_8g_rx_pcs_rbc.sv, sv_hssi_8g_tx_pcs_rbc.sv, sv_hssi_8g_pcs_aggregate_rbc.sv, sv_hssi_common_pcs_pma_interface_rbc.sv, sv_hssi_common_pld_pcs_interface_rbc.sv, sv_hssi_pipe_gen1_2_rbc.sv, sv_hssi_pipe_gen3_rbc.sv, sv_hssi_rx_pcs_pma_interface_rbc.sv, sv_hssi_rx_pld_pcs_interface_rbc.sv, sv_hssi_tx_pcs_pma_interface_rbc.sv, sv_hssi_tx_pld_pcs_interface_rbc.sv, sv_xcvr_custom_native.sv, alt_xcvr_arbiter.sv, alt_xcvr_m2s.sv
