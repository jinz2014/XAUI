// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sGd3pXYGKBCtgXDHO0D28M4v9rSDbIhpXZmcZ1HGFJyPpbfRs3uHSxLzahX5lA+D
qxNJVaHxgGrB0YmUDYcYEdnY7L51nUPsnnZCMJGsH8PhsBPQu21Th+b4XtMNBpU8
ZGATlF0x6gmFgNQNaQDOxxTaf7yhJ1MUJ4emIIeSdGc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27440)
wIda3Kz/9HNYOJDKezMOIM7oTSqxoJv7oFlpA2OZ3dZrl/FdzQ8S7CuP3O0OXYnf
t4N5Wb2N6YzgXg4EHGbhm0gipvZpe7MiwE7nII+/kwbt1GubZcp+EKPoHJVMYYNr
OgbZymi1eA9ijWa5FCaoD5J0G0h9WmIyL6OZdT6eYHfK4dU6VTwSK8oe40kc5tgC
6pk2S6Bg2HjW4tVfNdwyEED9CVtvcOQH3dBo7n2dMgH0Am9hKHCdeyVAvVi2541G
PP+1N/c9pNOqItVwEYA6pU8+pBL8sbmFg2wV8les4GfxSLptNDM/5OJ/jucB9U20
z9PQTtXtkgibDmQZuD0tZJOO9a78BbW14wBznp44qwoMZOeDbSYlTRr7U6WEVKLc
rZqWQLbETBq2PQhGCp/NMKWxhQEha+L24JZ1r9x0aLeaPhgdD9W080XMdme4tDmR
OHiQelL5O5+PufNG/4OszvMtnMDefOUPYhKJ9xMayChKui2GJyq5/cyndpc4okI6
PXF2nv4bMU4+Jj2h4G8hkoxsH3fs5LdNwUbM6g4IfGkI3brSZnxVVi3eL7L19fCx
DmbW2W8XIoK0Ev/dTQfJYf/oTJp9SYjhAyvPvLV25D4/rhFb0qSuBkWks80xfnr+
W98ADXA7XFe986DJe1saxprJEBO78cJacc6EuYhndCeA/YuvVm5XtRqOUjM11eL7
anNkpUtSf3T+KV5DOBNp4z8Ey1eKQKFjfae7kjXMU1NAfheG3gnXqATISjVvbp3w
vOIDolNrVDWkTuXfixb4sLogtntTcRNeR1wpomuKA3++28n2Nn2A43N/1HtA7Y4q
Yc0IqST2DfqNj+qk5o7HN9uIc4vB1/VhPxhyKc130x098XFnWBjkPvHz8bFj40gA
hW2cFlnTPHT4HhvkP3PJPARYArwjDEX4cPIV2ZnR90VvXsr72OMJPbiKAarpok85
H/DHTCgM6ztjcxo1Pwzil/co1mym5n/YUbflasv79JqokUSmyoCObFLRfO+lcVzN
N72D/D1JnQWfrvID9zZweByvSgfMjP2QMcfwOUDv4tF54NH1qQlGHW4ID/XbaGBQ
v337XAuO3/Zj0cetwb2ASlmO/qk9vKrYkVThGrstFnJZGdP7hqJex3ma/OakDqLz
bN6uwTW16HU3gXZrd3Rsyx1n8hesJsd1tbS/K6TaOFc09AfoyV95a+ogPoKryvoP
MDp4vbn3Zv5XNWgMhusktC460qM72D4qseQ7ZdAcw6h8Weo3crpnTZOS2HemBn+o
lTMkdUNyXFqRDe2ql5bemjgGZ1fZhtKAOomWpxh1PBJoEt3F2o3+IdP0wkETbwIb
lIHS/1Npv0pxbL9V1ad96EK0MpusSrftypUVMBaGNZg9RByaYZ/cul5NUYMPg/NZ
RQo7MFYYFIh7XysvvO6qDb2bZ1h7Y3YWwWDaLJxuQigs+lpkRQfpOreDvgIldZfE
dPL/K8e/cQf57KVUINq5n5R0fPQejbUTq74jEJn/xdEX3InD+R3A36YQrh22vKkd
u4CWg6uyw4lKsRPuqdonJzoCDP53IqDcCD0O0P3ZtCbYFYUm2slrW2i/UikRCDNm
vE0wBpQvv2iiUTGYujK3/B9rux6l9V5LNXzAUFJP0vY6v+LW7ezy8F1LaNq1o6PV
p17HhAuRhYfjAWSceqrrxMMLJpH88Rv9/1YxhbqPG4a80MONLeRUY2Ip1Qfnf1Tb
45U8eYD7Hk1agYi92Tq9iUmYw5AN2/A0fe/eiKXsf5rDfAXiooX2zJNy5nSu2PLb
50oeXv07lIEbg3XIsADA4+ZRVnbBFjRfx82dGsg1OaDYnI93Nb7d2Gba7LxIxo4r
XkLkm6/HSNex1AeQMJ/lSXIp+c2sTHNc7UyQR+I9rKbQYOomCxTfm6bK2DGI4rJb
pf3Z/BsSXkPehwDjhadzQEi/v8V3TdOlyaHKioo3TkTbfxAC8WhHQsq1bummR9J4
OqEiMaVrPpKhS/xagQbiCoy3PIB5ajHvpr7aNdjufTJ+C6RHXY6tNYv6JAKGHI/L
BPTKUXxYNtIIsJD+ybCFRGI+5P4CyPD9SoI9098OsqJuehRaWWJmJyIhQvpJIzHs
FwHt6lmx8jDlhvU4Efr7+LO3VdGLRVW1kZ8o5t/OyC+VORWXQb4CPSuUp6JkVPf8
WGeN5+//3OPbw6sxPWw+IGEe4jhChpsqxLbTZnYgQFCt1k30W1mhn4xeF5q+E+OM
vJdGleFi4DXD9iDO/o1zH++2cMjNOosZJsmWQZBvKa6h8KQetaTLM1lt+wFgcRWL
4GGmjsy4B0KSEJlNmnDJFBQS2ZZg4V/zLU2vudm6Jb4YzLut3FmLMgqjgYTpqHNM
0kmGwcTats35oKDQb3y+Z1qiXpv2olMnoo9PaCJoMEafQsU0ai8J+2LL3ZNt+stX
H92joFKjq4xIJWrOWteFwispU6K9pZHZnLe9AfFms8DqCq+A6dXohpiVvOlSkwWB
qeQhb7YcQOwruUXFjAAaaugb8tXbVSSoP5T8fC9P6NcyNWqfDFu8LGprwlfheLHC
7KHC9pcMBsBE/Oee3PGCsbfO57PRdKQs7HOy6p+zLmGol2AI6K0rxWIG4fOHA6Ic
o+CpRY092kmlIFWrmTDF/4uTczy54Tkvg/RJkmsTq1Xq92s2fH4T3IXvrYsWzu2w
KUBL4JSvJs+kN219m3CMPwvtSZSODrf7ZrwtYe8U7F5weQ4Ph0jstKrRShGchNbg
FDS8RTzB1dzDodHv+zkl057wVBH7DXjMbNrpMysrSSlbepOPQ792EZJHH+/RuZmS
hkUF0MbqE3zU6FeUqpM/7AQNg4ffI071EvCLna0gN2YaGZIxXf+lY5VLb0AVi5tR
pN7zC6xrb4aY5+0V4K5eYfFIgcaxQpluzX+AlLRb2+zyA3L7WvnOtaCxoJi+w1iA
o/vGwL4n/WbkusybkEdcCZHeRBHox+ZECsV+4YTL3g2Egt8pOvvKcSBK0Nx5C44E
uF+EitXfU1nc7px2mS4jOkVYEXd7d+yGj89wJ8Er1HelYhDk3346J5/gOqm9jTQO
KkoH2Ik33ov3h+FHkKwOQthcxtLoiJMGpV6K43WNhqTue7YqJL7Xqs23I2jqa0fA
5GlpBdgO/epnfpiOSp2YpThc7xCZl4va8CsJf5lslEnvPnaYKgYQrgJ6aOF89Mcc
h9bjiPRusWSQxzzAfTUTsfSFCsTPw4okMEnPA3+lILADM1xa6ucAg/8J4hibwPFn
o6evX26APS50MXNyMPZXPzZS694FLsw25NYs+Xh76ePDm95IIwfHkkberXwEthhE
8klrvYYeSZSSqoS5fMDN6Adq4l7hchSwJ0kbY0xi1upwOn/psjW4fyuxmHgSungw
94QRJy2iK76IVJ84jE72u+npDXpQlAfqeIKMqAYYHY4f6ZscBwPZmg0kaObojlFI
LEqMA/P+8Ky86VE2R058EHxf6bIUGmxtT5uA0MX4AlBdDZ1xL7knPl6BWvqOMCcf
VW/LsD4+GrJEt1zG/xNXlBZ8kVBeZzI/W+m/3F3a+hIYFp+yWfx9QDzxaWGkZVEq
yym03EKZbwdzzuAZEhgqtopabdA3+dlBjq8PoGCtNZf92LdVuDi1rJW6kRjfwdpU
kHDBVmZJRwMWblHa4N9g8inQH8LnQjqnNwfQJk8LfQXGYK3uLHmBSp5P5UNgWoAL
bPsrE3GEqJqQQd+drIdwEYvj9z4X699A2ru773F5XtAx0RZbi4Lo2QMKdqPseItZ
wlMPy0UJSUCC/pOkOYNDDG/vkChspFzxrRLP/6YBipXNBzXpGj7oau6o3yaKpIYM
jzG9IukUnm6mgdvvMVJHt8w9Cbx1iplT/XzJ7l2MRhtcOtgW6QSIjSGQLEUAUge1
DHzF9/ofkaSMo5orANYAT9LJI2th4x4tfwErRGTu7X8pIk8F3DrZEZjtBNd4P/Sg
pcMm8dePGtEL3XtePsI1g/Z19u7rRGKR93n3nmWYVd40hmxoMTgowSqlEa5ZW9wf
6181lDjdg6RI9P2QnNaJJQjaorvOVLmRlRqgtnAxKacSjqG6gMjBa5KAwUbd6/+g
JuWGXgrjiKNHvldG+89xdhkT+3vJWw040+9NF157kHiOBt359FW8hStLI3Qn6u1c
TZYO7bfkGXJtax3S1rQWx/h4dlPhd6ZrNIgpv7I9Cr87o0vJ2oOwIOmIT7w+OtEg
WFBaeLdZzX5iC4zKvSr/IE0RjSeTFUpvJbW48pVrBTY0ru9uK6RqyYRA8aJEg2z7
ifXRH5zoCGEPGDc0jEtd2lqgtHrbfCA0tKv4vsKoMhvQgyyprqhpAjx3TfIAR6xq
EfWfKTa4gEM3HpC7CUTeHJKLmVmToAWUDDFuVhoCPiCprrIJtG08XAfwzKPwMhaF
NUx2vnHOVl+uI3dzxIfHqmw2NAbadJwuRZzeDxrEskyXnnqE+suiwoGcvsg4T/jX
V+zmw8eHP6leiilJXTTv6KWblzbT5raNURywvd+FPXIBMaubDjuwTJuN5dldmj0b
ZnATv2b6xAKPQYb3ipx4MzIOdZciFQRppalijquL+/DgdsCsp3Wh4pHZd8WAmMCy
lJfpNoBTac4tV0eXTkcDuVVYBbO6UzLNR5PxKaq//7rI6TVhzon4DEBlL+bp/qLn
WLh3RsaHUYe4TuwVAAX1Rr8vYyuTdzvZGOnDHd2rdPKuQVJ89oJqsAk1YC7uXhh5
OASrGOGKQBlabY6K5nd5JI+3TEpfkPLLXIBd6RT+SwwUPHoNRRiCPCmbMq5TjJLJ
zU44Wr5L8Pd/wTanMVw5rBUtw+2HEieXiSFwtC/mszo0ITVjKxdSrNEeoW7yXQNn
V4G+/w5v2p9H8e17ex2WI229JCDOJ40xwQC/VuEWtPt9wyoaC9Bt8vfT5jjl21D0
03ze0vctUnfs60owr0QNbx+PXxZNZ4CQU60RF0fR5a0GHClCeElz3xXxy707r3Wv
QAp7fBjK1b/uzBImPCdHnD4zJOJOutBffhdzhlZJOhnH2Jv8hS4zCF9i1c+e9odT
eWLO7/w9DXeKXuLLq2AqVGTao5ze/PAT+y8oRwbWTtMStgj2yBWkjNscZlifUBQk
cvJakqREqiqn3sUZ2PjrX5Ov0MBfSgTCmOEhJltXJ3aEtIxqI5igm5CFj/YeCzeS
2C6RR0YG1SYjXLGrv/+kiCj+2nfCXuLHhGyprbrg39SF1XeS2Hhun44nipluvjef
QxoFsK6ZvVZr5g/0WXXdDBhjnZyNfjEN/bq4Bz+xAHcQpGiAsLFegrqRM0aBJhq5
soMtpSpWtlBDPa06A5oJvYYGkea4oOaO3cGQ+tDMDr0k2grjLJ3eqtaDv2Foe3xE
hUSJwrY0mx6c1ygPTUGVzSGJ5CEXf00m1Hn/Zg7qYAbQ4NzpOOQpWPJWSfc+HEkC
9lcrrLmzC70nPH2J+rXlJvT/vY0KfyUA4H/uaxnlTrZsgN/kxyjKKlRI/5rpTGiv
ItlIxPWWMq70zuM3YmJV8v9q0BH7J9lR323HDtV+Hsd+Yfm2xC5/gdrJFASCIgDc
1ZerBYjuIhg675Unr0b+6i/yLLttnxL3cHOV/6kQCliHDjMUcVcWiiryA+8GXTWo
4CKjkp+a++5lJpFgpioD4brggyIustW0UkNLVn0AQZreFrOO6/JvI3kO4mG+rkrv
S3zVXVCn36mo+QzxEuBh8hl7T/OzEQO1tYVzRkC1rFd7UUAKB4Cy7hVknm4JjGDP
PSIWTf+XfDwULoOa6/TpfWjOmQ3mHFJin8PgVp5jhk9aSrhRn46vX0cCvr+Bw/Jf
mMMlIF8TckoblwuhI+cEae+ct9hvksYSOp9liHzWhTdN4QGKn0enXQz3h6Eip2D8
tF+5IQ1cINsou4JijXa02iGrnm44aPuzF3exiEdPmX5emfQR/3s7J3TQ+41ydy0N
wU+S4YgIegzghZFjixcKKK8LNURc1qPOJzgxa7D0tuII8T7wlOF5YCG+mmSALpRT
g9mJalAb+usOMHUUdtEnrVWouddWA2tw+CpkSaOXBs7F9IzV+RS6XZlh8PnYaIrB
Mqs9cSjz46s00mfYZsX1wj36Ah6Br8kVbjBU/u+YGXsPkeLaviPXWC4dxgOBlKM1
bcYNbhJbvJLcm1UF6fLxU0F8M76yd6+abw5ho97dfCD0Nrmh2cPBuzuNZghKYiAk
zughjYIZy90bD1BOndv/K3iMYX+AXLrTSnEaBGqMgD+acDWQUj8ricN0qcmzq6O8
RH2bv6Ybwzm7GYiNEWGYodefdZNDESg1Taabs6anzn6XKoOh+1j9uXXdC3rJoqkP
59zn3l/TZkZHDXLgsQVN0FI+ivFCmZ6tG9+5RC7/V32rpCN9Y/4JSbOXqiPHQ/ev
pz3ycp2i2xXT1L+ZcBuowFflzzf0tpITkbvsSq3rwGjS20cGxGL5UFEFiXGAH67I
BL24ovmhScj/1GRji+9Dzi6CMnKAw/dRCX7cxHODw4spfZm7uFS0+l99ujvIAAq4
2H4y9IyXbk9kvSbeP17j74ohV8wSuLP1JpuaLVlWwYLCj21VJ6PX4QsvV/hergFl
pq1sV4LrAnVr4RH27NlpVW1q/nMumNk7YCzMayE7MbIURzAKuFHUMZgAHTeA69VS
vwOtrapYzKXXOOZ0G2qWcpEATeCPKL+ypIS4xMeXeWXBhId8fyB2qnkk5dhtMBvc
2IpLWf1VtRuCXTfN658+cn9gjhJyNdD23843LyQ2E1Jh96pUyhf42RByynM1IJiu
LuNYWwbyQgIkg49nMdzwtr52hWoDS/XKyGafOC26LjywBv0Ls27w3xlTa3ahYAOn
AIlhQknpV2YMchwtIZ9BPYFX+PPjevWa/FQCTOgjwNBBdAJTj9UQH6FHMSKpbilZ
ZCnckUY9Oz7Rcvh5o/IBdke6UrXOOrsnxY4Mw6p3Si1gT2VV9AQF9GChNmggOSu2
aosTF1c4M0BzkDPA+IjQ7tGhn1vb4Tre8WvRyccyjnFjnBC+Nd9m8qBSyN0VJhUE
VWY/adSQrzbWHDVelzVoeAX/QC1uvofGiliV4InVRRckrc5iwzE4y7evyCZ69wG3
HFm+9X/Aolcuodz+F8Vh7JVG9s6Aw6GmpHsmlmFmPtkkTG4DLDS19PZeyJ1SIDZV
Lxk46KVBlYZIYdM9IadR3YnBAwQoZKiEDGfTMh5lz9A+3gyXFMdzLB02nnR2HJ8h
7DYHoN7bZNCaSTYeI3RVr7pbRmAH7J/hU7pE3fdrd9qNYO6nBVj7dOUDdi2gMBqP
6Wt4gsqwQ0DklHdJtN87jBFeli5dLvUd944ZhcGZ1/FXXnLQloGBKbUWyo8NNMk5
Ah+VBEIb6YnmjWnCi5Msi4+JMVxTJPvZwbUj9UN6b41Ef0XJJOPb7tc0aN0couV0
T18RCnc2wcUQEILjMvsKoQHVkd9Dv8HBc1kkJqjCoAB6tBOwKJbP5VTuiUWx3Snk
N4iWJkdvM32tl6+qWJ2QHXsT7p8kj6RLvVL0kK2vo5K4zHlz9C/mbrJ2PIfZPWvE
FhA0/f3IULXqKx6KIIE7ktnhlPWpfq+PBEx1xsdXqV0OwrmkgwSVUnQGSQ/NCyq4
GD9kbFnETox8w8awijpxShk1T26HHjPADt4XJUZyCU/UqQptrsVkGPaZ9tmvMB+W
eNGzIubEcdLSDexp7zZeBd3mhog0yLeX0n4Ewa++3omkSFmjgWSYqrE2EXD44aCM
pLmg5H7S4GtcUDZfsrU5r5AoaYIXwApSvXMY7I+UtlenkECK1F5kHjH3W8xYMIM8
SOPvgwy6MpQjd27JVfV8+OqbH5f4v3TAz/CB2GTFO+BHnjzgAm94pGENnez56yzs
1BW8eX+NJ420Ve+VDJNafeywDqdPRG0AKOqh+P5xuUuSwFQzz7+ctLym7DGiwHRH
NwwrNyCywfvbDhjP2chSN8EYAaP0WmW87YBfdk0L+XoHYQkXR+HndqH5PcMOLdzl
rPF4y8Oz1zPE8DCR22SNCfcy5e2gLTE5U8gMjJZe6H5zbhXhWEbRDadELRhbII/v
+DHuwZHvOuMQw3SiyWoHomQQYSywphYzk9ShhRqNurOEJcS2kIR/pgQ7baekS5oO
Papgx3PMV/TdFcLbJWsQ+gF9WWBHls+AHuuiqVylmxz9MKWDA9r4EcsNRn7dwuH3
gf0fj+DvQ9LmIFC1ltveopNkyIAfT1dCKfPQFJNg9+m2Aw2lToH7ryewphS7oRH7
doS5bvbecQNxKVmZbFQIGtfaPCxTIMHGYnjpgs0yDALxBTGXUX9ObxS6UMOGGiDR
ayndWCUcDUmvUsg6aDx7jtqk+0JRZG5uHAC2iRnYjesO+35mLnFY99AoPN7WEiGu
cjrETtHHqUChY9idK/RlREEBxeGiewO2mvPkp5LXk99nYzBiwuOUhs/MsSzD+boJ
ekPqdptyHLt8uMa3iooxG7A/x8v7bEGuEaJAtL2uL04AGF/xzLAKHl8VHG4VzTDS
rt1ZwCyye6u9Clt8RUo7h7TZQFgOtZo4h73MNajVhvx83N1DEHstIjkk78gufjB7
GFxEO8MRN12R3qP72ICDVUE1i9gJqIsfPOKLGCUWygSZTtBSQfHrPkumQX2pcxXp
remG6+jEC2nG2rQKrqYz6n/+bN+7jNdZYIryHFM2DwMh2VgXywiK1tB7Kbkd1Pyy
jRQOeymz/PArcfoHq9dYBIV3z+mb0/dIMSt4tAB2F/XaeQqSPVCKlEFXvwvwgc3z
KYMF5FCsud6VncsAJ8k3P198YwpOgOQDq/hZU/kuFYhNd5+Uw05NvN3pq5GJhx4P
UWkPZ0wA+5SJNANsqqR8tI7QqKe3rnkuvBYF+ze6xd+pOoBpwQMvlD0+sPdFSkoK
x6EjbW904qRXG0qfKur4p3Zr+Sx1EKwVkdApgHQa+JxVXicqlclV0j1JuSoI2tor
Cnvhmbo3ai5sS1F4yfwxq9szOjOj5GPSAWsc4T8RMMQkIKq5A84+4sbPaKdh5ohW
dAiNORSSPn3DiIDekxLjwHxa1sHTzyTswQdId/mYa85qoBnvQgF5FQgFLTqENa6T
tyCjLei33mYVDkg0Jhgh+BEZFdazeD1DllacxDy8xOqZS06Iy0vPQ35tbMxcGk6q
T0+VvfwSN7X6N0vIIZue0oW/WAjAYwtAiYzyLVhLkNIexzoNvqUNOaBoRsfPqTcB
8743q+6GnlX5rlZ5UJmdJj1NjR7iY6a+VEO2gxh55DMhXaZTe/R5iYzvYjJd+IpY
0Y6Qo2oflYhbEHUa4Hq1+0WE4GRraeglwN9dQAL1PnJtooLiQ4wPgJ/Za6TxBqqK
rTvKh0iLdTzqCiGFdts7fJun2+CekYkQ8YjtX7pQO0a2F1JlphgXt6NJsKQN/pNx
0OG5u7OfPMlgSV1KMyBfnHUDizHYoNOPOl/8sO84RLvKF7/MwREN8PK/sUAUEVwy
ot+6IlRrF5d8o5GAvZ1nyOJbNhhNu1FRsSCzZsx9aEJbXpTVlxsNhNlYvPIRyaIy
snxwQw2c6VXgXtfQbmRITd4nNo9qzrRtNHGI9iLRa3+uEWXadrsZHD6eDjLDDYAM
Uz1IpDDl+7sp1+y3hcN3/u9Z/Ug0utElP0AsE1FtYcFVJzShVtA6XmSltfbeq/Wa
CrFn8tB3IFbyA+akfXqhXp4czM7p48SJtHkWXDPTVgoASxg92Z7AcGOYjrjxKIaj
sdSSO9g/bhwZkaDLkzPa00sfSFWHAiHe/PuZ+XCPYUQnCYdtE2MqQiwW0UDGT6rG
k8WTPOMKVLcyrQHxg7qmqL75TP3HkTr1H4a2oKyGVE5R7JkLTS5VAQixOOKjiJJN
oeTXVWUOe+FgfN7z3ayMRttnQONJpLn2ZKvH6+xJk/IDy5FiN5XO50gkk3nWQGby
rSSOEER/aTWl1NwNNW+SwLu5a6OL9ngLl5tDJfs6UT5dT2ete95F24gn8ZMuiyXy
iRQa+TfGRsYHroRzqm7AgJCRbG3j7W73cKEwRk2jqgNQnB2qDgMmSqnrtsA9AdT+
PxX6HCttnKtdvxt5ofmQjCrDsOPobTbmQtJgmbmCw1yc003uDkTMj7a/9mjuhUqv
0FNsK50p51j9wmNLSjgFWu+yW6TeiCPDN5//tQQ2AdxraQTrZvUyrPfD+gOslSVj
ZVOCWMv9U/9dwiWPVL7Hf0q1lLal9vHGSWlT/lNbaWkc52Vwnf1qAJh/GTxivikt
G+Ju3UV8blOx5eJN1tDvb4+oH/wb+nNlhguKOp4sy7t2+hiC8kfFOnhq/zuUWJwA
XBN6fr64x0joxPyb+dq/YjMcKmHMGO5Te69bxSRO6V9Tddtk8D0WkkDgfFCZQ78G
7EnC0JxxsXE2yJpGdxOK5NiRZgnv+TZgcdU6acvUEkK6UnECuUkU4Us32mg53imB
Ux3VOFfRGcv7L+bs8MiTMCDe6U3sOF+hUJqUjkM558vaTTvD8uJUDxktjbK0Dwx+
QLANt5Qm89Fixlzf2oNpvv52anDm9K5SKlF4JolWfjjF6qZ7+KYpeHNKLfUIjNCB
3Un6s9MgANLAIUCFtrQ0r3PNX6q56NcptTSjtsz7JkACY9Jab+mNEghqGIKxYIjx
YbVCCR4uYeKVJAU9aOPIgIqbXuBj754PTRpn2CTrfU4aiyHR6bH1zQTIbDwW+cqo
YUiTR2V9lfIEJhqPSoaXPlMY6zUOKihPpWW+TYjsnU6EyCwxhtUneJwtgjs8K0c0
QmdNaHWrXVwHIeQLJsSgbPoBhB5ki7MVPkOQUDUA1E7GQOva8s4I+Bv9wlDP+3IH
VDyuzljemo+qoQKXzhYiJ6B9lBknkOV3mkKEZ/2hCixFUphYMRdsX9OhsSTuTIhI
lbnpACnMN7zIWDQOtXzr2k/pjeM0OgDLuBWmw26zk6UQykmUlAzgc7ToDC9WGhFh
CA1ChH4EpUSCp6uzXSTGgQx5Z7Ya/MOPNiqIDqmG44Epee3D0kVHVwHlG6jU9Sm7
pD+GAGrAj28XRcCY8PetE516S07HJxT/glbONjCG2BVFDTM0bQvDsDcz+AV13Tgl
IqZyeUFBo7zkAyRnw2fX2ZRMNFEvDw+IdzSQsaKW7z9VTy+ZbRZO1rnfHOtjDCcW
JohhncC7PCn+N7+RPFnyPlC1MuWWIyHJW+XuJTwsYkGAr0rg4v8PPbckjlski61J
dOxuRj1X6hYIdGGaHqLdIkRjBbArQfiLWFxBQff+gzEdyv0HFZZTpR5pA+QI2fr0
xo/qU5DAiHqJnIwuYuVm7pzseksx8+dk/m/FcwXT9EgKxY3FQkTNW4x1XKviPnfi
kFoz0Pp05QbVrYSfmdQnH9llADChFAd5JOdS7oGOYiIA1W+FOodd84eTHE5m0syt
pGKMNo52idQQQU98/52GMLDik8T5zBolxRuUhxNzhd8itvJznCA4nTWuabAkbJhA
ZhWOKtHdYk4H6UdQEt7Bh2aeBUUHyDtX2ie7FreNED87lg69UXE6QCHwKVk+Zl1P
RYvElNvfvKnVq7kQxckcAVyCFt6NEVBrRcAOrcekGMWwTzQxj51mmohzpXIu9lSY
Sjj1XY/kcjUGYPaRQf41a8tZ/VUSWr1/KQKtNyBbDZBDtj8sGODBn47ep6XQycMv
bO9xzTZcAKTiwcu+65yRIklRwhK6+DlG+1b2F9LzMPzj2O7R5qMkeg06+9+H6Waw
asrvpf6ZTRhDHGbNHPhD0ZS8GedzqT/lrZ6U8gbhFfx6C+NtYw9qbdGJYepvp1Ph
MJTgdLEK3dVOfB+LFueFhxpcQWZoUmnMqBmgfGKFJFaae7tz5OijE3F8rQ3al2/K
tMU04e700amqvQurFb5eew5tMAptyP2jvva3iYUKPIIJFGWWB+Ri19GrM6hzRjyn
ZHzZ6RShdngFLgf1zu98IvA4xuIdQuGWiKXlZJcRCZI0tzxmrc1AsySmh0B8vJsw
a5jnBxgKnfli2B9HXJ+ijRcn0hMreJzu+mm0+lcC2xUA4OgXQyt8m5FO5QEHY+mq
hpTXqqMyfQ0c4/pM5Ef+VUqAkNZazB4/DFzVYp3XDWNFbdqEfy5lxYXjA0nkhcQX
nDEsMxu2TBBiApzzzdxEIuxwiLHCZQbSpFTsW9jm0fK02UG0f659glpkstEhQ7Pa
8QiM52mOTf3zBbIYiXsCMN86CU7zFGUwsVCWvsEDS81Q+2QXmiXsFsJ1rrgqKNRI
eT+X2iEjmhErlFELmOwwQjwSSYhy5TeBz+wDEaoU06t5h9nKhGkdSthz3BFwE/8S
pP15VQu4ncRxc7e7V8JIqxzooj++/tFy5fKs7iLs+1jGFsRXWFStwHw5bZiDWLNo
MYgLaH7zIbHHP2fPaTjsV915ZCxXXud85Iqzt78WBaSf+fbdlir7hu/9P5cbiuni
VcbkhNIBaFsMqjVx9G+nKVN9LbUMAN9VUcv0Lh1ynqQkbM3rhe8x9UIW+iyLrWLx
kA/cxJe+e0SD5M/N74iXz01VS7L9PBFBesC5tAi1QH9J3fffPRI8V/Ooo5U+Yd5X
mvfV14aA455XWQDiT6TATWroc8UH54KXLv1qFPvsBLggormG1vACsK3whxML5O5z
4zS6pmHDlPCfacqHYjjQbs+eiG7XXuqxxbkvfvRD45ZpcUSiubQB9fUx6qfppoR/
2UuAG/LhDX136D95yrW3PV0kdrVru4p8jq2E9kQJkZq79dCvScs0+YzXJ+HofQJ5
n8iPJsho65BYkp0hrSfZtSidpcrYfcIkkFoiEZLQUKdznbfze9l0GDDvTa9ncMxr
fw90YEIgab67qd20EHLVfiozpJBU537Q9GdlRomxofab8/1h2Kl2g+nDLA5HetSF
z1PrWL4xXDbqpckHPMwc/g6nz0Z1f3l1secgUIrFVg9gXSedMtPMRILo0QhR5Y1h
m8cdMTJCyErJzoXjgyycnBTPxVy9rLVLrTew9DGxpIpWBMFYERsI09MWAo7mPMUP
ra6fPHXHmou6Of71Xtpc+l6rtzM4hrFHIbWq3QOH3gR50v3d7TrF0rkTX8D0Xqht
3WOBsFkH8OvP8602zOcDZfNrNCKdLBNYKPC1Zk0OeoFggnJrUfmeqn5xdeHo3z04
AabTVv+ub9Da/hm7RBDpLM5qeabWmbfZzBoHCAa0IJqCFxm5Q6XRKl2O5oVEHc+D
J2M6Rezc71EFa2pttm+m+OMwBqwjrJrOFMOHmw/1po+ldz24brtG7gQO391I8qsg
44hJHDA4PY2+EBgU0YDLhZxXqQWRxk2FMTlr0wVkXoB1KrDvg90eHC2+vj/lzfbo
D4sh9Ts+gmrBYfBit7k5LsiWvC7bsGGWO5VsK8lATgDu9DR6Mp8tpZoWbIZSB4XV
Z6LsJkFW1poLz/NEehyanYKU4e6fDUNvIvJW1NGOBSrK2+XzvAzNFx/G2wB8yf/w
pCKVHyLNgl3BTHOmD82NFy9AmzlL0gti4EnCkq76UwqwKKfhyKITrJaNSdRTUS9C
nRzbpmnVv1A7j0vmFPVeh/hxIkSQfPBnAzIxkEoP0hC9k6tMPulekALntN8J0p2O
mBVauQL/Oi5eAWm99Vp4ulEETo13BAdl6Bu0jgtKnWu44SoTKw49eST+q7Svmez3
51ZRx2aWpNmGdjTe3Z7jAaxzgLebh+HQTL3UmniANvhYO5metMR5uuMEPWgIoO//
E/a8E7sIX8QnCmNcdBOOs2XYuzpYVnXRftZqnzpWw/W0juUzPjsCHMYSEWL7X+T9
wDyuiWdcqj9dGsCMdmXfiWUtrYu8amS2Q6DLVrBFaAcOYHAyVOZ7b4Q2MpyjxIjo
bMoL4appNCnif2816V+pB3g50IJ7oClJp0TWo58OuEHDAiOrFoEvJ3KT51w4GV2T
JfD3bAdFq79ZhkT8kuQyMjACEz690olHyTHPBBzRF8xw0DA4sznCsw0CCaZ7u52q
PYrvzDuGZVtPORfNpjS/gbzHh5KLw11yDvj44MOGFgm0jzFvtn3H+LWN4E8oHk2u
s3usHrHah8jGmPyQnc/B1LeaUeWVkKnEp69LPgwlGAulNKMRQDphAUH51714cgpa
DDGwbrt7hWNDUfnb5Y6YnSYfvBQINznuBYhJOsgsfFHay3YIPjhH/W/IfnbtJGaX
mNMIV8YRR5/LsC59aAsROJ1AaoHVlZo2Gbkj8m5L/IWalGlXt0068lehwuMcDyzA
A5tAbAscbvY5QMPD/ewnFZjo8qsA6fbmZWpCioz9Eaf6eN6XqA6Ds3w7KY2fK8iq
tOCxyjarJzWZlZ7J50KSY+GyyGP9c4cU5RqIgoPEZ8alsPUFv/Dsq1j0UW9UqrSj
WLBbhKdv42vvIyV8uH8TsQIl53F04uQS5N/a7nxqFslAcplx65WBxGGbFfMXFLeV
tjcdrpC5cfmrZZaZDEO8Cfb3UcyqX6uTncdOpWwT3vtaYl7THiqE5gwiETxNNMfl
D+lpbrC2Yl+kr7nu1S/5Upw8FvyTHQ+M/9e+RqfTEgnUOMzIcMr+KIeKfmtdxaU0
oZ4SYE8szYHEZm5wLdetFxrVhakcPrv7acZSVNUXxcUKlfoimlhlMq0Q/LW2BeUv
er6xvxv0Vo0iBLug0jKX4KFJJyZNYPDYcqgWRj1lYpfsnbx0jR0Y0/yIekV2TwA+
OoZ8NAuCofpphmmdwgQxMnhEdoqohCN8zEwARKKHq5K3p8KO7EvmNXTURirtilw5
CcOslQj/aP9/TRnzEdT6OTCCZNYGQH+AqCIWFucSgH0KVslyo5eUYahtPWTwZoqP
WyKqGHcos93k3QoGdC6RPuAkR0Qbttt0j9IyscfGQRnCpWB1lzPm3hHT+H5j5o+G
4dn6Jh0bmdZ3uBMuUq1kTm8JNj2YPfEj8pPxtBU9OwNvwu34TkXG+DPEBDj1W0Q7
d/fTTfw3CBF2ucEThFODLjgUbUsJh0isa1l2px2ZyVzCJDHvT6ubK0BhYPnWayUe
jU+TBydHyB36U16q3P6mQ4itVVFlwPAhWhiwAepKi+gIL43XVLwdaj0NidA261Ys
JIhLQ5p1EdyGnhyL1nKxWTdhzP+gNQdgs4WVaREyW1uhnpuU5rHm0y0R4b3oFEQJ
5U5uAGL4wcJnkG0D3tiAnwRX2JUXVAW+TEgqBOTlaGn7G5AqS0bcEnSQxdAAd5sH
FHiTh9YByqNYjobx0Fmn77Q2N3ytSssCzYH5PFVQH688JlnhZRNxwzr3QLkkT4U5
CHGoimTwadJgPFfZaUcnPbArzjdfRmRKGRIYjp1vycul2dvX3z2Bm4F30SghuRkr
M0lgVv/FZmZAGmL+c9Bxm8/xrm2p3jw2GIvKAQ053bOAlf8bI534SsVBuU6JXHWK
9idNZ765LRGsdwa7WatkO0mxoJx1dlr21xSLr/574jfkopHdj6JdGLtAOZYzNrmy
C3v617IpEwmcy72iLzKTSUwGXSLcD3RoTgXvMTyzbyF8psbZfB02rpWtLCfPOZ4t
cdOy56G0Z1U3elqfI9dWbEueOTTkc6WG0vQfrXXhdfgYKFjw2b2gNmtPNq5siiXI
B+tPxjMy9dnLrAS4z7+pCUPEKDrYlVLe6aCLvZa5Vq1cTdUp32gjnaq1E0ZlaH0P
ez3DNELYnK+Kn3kbODEPv//3rx5Pj5sNis51QUlKW2GBrDPyX1nk0jYTC3d7Uw62
pB6QDdWp3lulcu1bqWZaVjNDpsEELlQAHfXRxkhYKo3kDA9bZ2wy4D8uU//JvdKu
N0GCNHGlQtCrQ01HqZggvQB+duZGZv+OKZulFqer0so9PKHdfj6oq54HWrM7WQn+
/6AfJrFVXv6PfEZBkGJQky8cKKsYe5JHBagzTZXBimSzNJJI8NtLmE82E4JyWNy2
28cPtD9ZtE+V0Vl8jaSNA5ypAd0WPGHmMoznIjgXr9ltS0aAXL4fRyY5O7ekKVKw
cvpLRXDKLg/eTdwPbW64XNLeY48blMQWIqMjh1oT12K3mTt68W/qbRvlHQRQZAHq
nkWJacZifZ73irZMiW9C4NIaMWW5t0G9zUQ5UcWV/pF3YW5E2QLwEAXBKFqcnJpb
/t4+/4kykv3KGhC9jETs/OJ2wcfsibZPjTRD+roKIfKu9JFqC1i3+rh9iaX4knKa
bD44KeaTHmH15Umilg+3U50DK6d0TOYJ6dNObRWNK+lgL+P3gU8ksDN0+RVK77K8
UuovqvnCZdg+dgQNu0WKeosSCuTLcvOYl8/Hmk8vzGpn0g0nCXrT2iTzA9mdJv7S
q8bqGndCwoiQuT5PALW4R4zdBCl8kG+Sv7YhZjhlH8s8pWgf+vsu9GXheSRgr0Um
PyCgU80En8MIT89sfQdVJTP7PnMpl8n95GGybIGqa6g5LJNoLTgcFD0xV5mHwinl
qPmti0IUxDtSQeWQbHguU/A9W5IUyWH4xfubWkIAb6l53T4u9gUgMEWiFFKNtLKb
ne0hff/PXu+A3YnI0NokLGn05PFaXA2CfWuyEWL2l8bb40kcajKi7RkhXlDHBZLj
wKI35QKfwyZd1ZUHhkpFkkhgffpnPgaLpvYrTuXMBj64xv3SvM7VgtnjCPRaPWdZ
XweZrF4TmLM7xnVKHSxcJd9Fu4RquxcUkZ36ciRJtwv0mLz4L2uUHpv3D1k3kgTm
mZlw0BkKyeftbNFhX2omY54aUVzsSQxDFqBxtzihyLB8Tzw/31CR8OC2HnFg4S31
+jOexYE1WmLT2iLlgfCmLeno2Szf759jVG5XC+rlCH8R1ywudzof84nLTXOe205X
ArB3YxLKZTOzA/i0S+ms09PMBvVdYzTrzGtu9mKU3OxajXza9SprTyOr3TN/o+Ee
/zmVUhuW2I+VOO9TKepp845XEgFjlotEUVrNUkwDNj7XxBobnlXGMxsr+m72CrAc
J88qkUTWgiEbE5c3IXnXmP81KZ3gmKvFrpx4Teb4hYZK+mEoei/CIfHWqnWKKmvS
0CEyH6F//hfShzglwRx1gUfXVlza/SQRPag0BrTwXWSiWVAxyFnh29OUNXP0uz3D
us75XQaCxLWeU4/HLrdtE4QfxWjpYfnmuexET6CsVmlv3r8AH+3kqEaJd95hxdaO
BPUcqoohaW1/9yWf36j9dSgl70h1HrOJZ5Ru6F8QLh3JhnMRfcmyhyFVNn4x5S9c
za5nCVpSvSAQgWib6g/gYGmUpOYt4zHB/l8aBmgJ86pXSqIgxRt/TT1/J4sSpDmo
an2IB0QV8/hUC1sZ/un77OaU08noPQtpxLQjEPac38916aQyYKZ1u0T4cJVhwT+w
tXaJctiMbtVn/7H/GSCaQvzB7X5ZZXL83naHchsu+z3eepGoroGijOscc9kk4OjJ
kPcX9SIHdmnGdhHOTWhZYrMq+KdC8Cf3tBROnS5ePRjHZTbY/p/i+JzRiMpVFrci
5gdsjmMY8aIBo0wsV998puaYUZQKmpMQ3gWYfAoCA40ThYaylCb+MUyR7QUdOAfY
udPO0qzfvqmOWIEG30Y6u2MxUGhzGySlCOJ32nzFIyhd96bmdk3K0yFqK95bVh37
UFhJfcQtAU06ia+vLilHcic4mbhEWmWgxvJMZ5Pv8bOPUuJYwRALFnbFYmMCDVdZ
GRybfbW9fNIRagvBEA+kvJTnQBWetRjz8j18+2Wuj+g/6at45fTHQp9njNdjPiEg
suY7APsgRyKIX6A+vajxyLN41I7ZmXZv4WdlFi8VIj1+WqnFd4r10e8GyjAfOw7e
68VamMF8DNe6Tv8LtlC8SHexNZaOtsqDUCR3ea7wEA0ZRrqSJ37fINcUNiuyTJ9w
LMcW8OYYgVl1I2BoK5gLAQTmJ5Cf0VChhGG5KVMXc2SlLN+jEbJmduP1Fnu3VD/2
auwt3EWcdrxVs8cZ24hwYMv93nPBPIxdylUb0N5bi7jDJ7btnkqmlltVKwixlV48
OScXu8l4MaX98d5IjczbdsIS/B9r3vB/ZV/Jmbzax4hue9tTGFeihwJXatcyw1Rd
5AI8Sd2PczLoD9zJ0yOW5uVmq1cmuhRv8c3l2BPHdPhGg057W8LgEMIP3WpdgUnt
V8RYCii0dTVDd2AcGctgElAhK+O4X0xnlQlRhO8siBzw7AQ4/q7ke8xfSFaywDLN
tfDp0vpRILyjPcvJFyKV09PUdy4Af9WgGhJlLRJNvzGtAP0dE4Gji3gKUs48QKfa
cmSByPSnaW10UINbmVHQfAIGgHIgNWOxSI1R3FIiG6dCSsX7QDNKZ6iowEIN4isY
/ccvTZHmlq+TpWNm107jdSGUpbis6WGTuFHMU+JCn7wRdiAqW+D+kWZWO1STMLjV
uEjich9mKvH6pHWMW+aKJ1GitI3A849TqKCL13Y6T/o3/mWRyfR5Mq26YXprjcMI
aZKoww5JpxztfBHbf3h1djk7s2Rkrcf4OwrSVrl0Y+dXiU1f75X+Tbh8YhvYfxb0
g6VdfsvftJpak6pVvI1rAkAbdLhSHVP7eVgdwFbIEp8T9MNFjKsDDBYntiZKwusZ
0emQ11CC4qg6DLhbQKdZlXJ4x1foNijGIFOmQlbciGDsDfmKZWhwk585QDxMmE2t
g4GbFoAMeSq2ZKxX0qS/HXH0W1fAu1OtxtY0Xua2P67lxlGCduO3ORmYDWHdUvYl
92oRsrq2d60VhgA+6knLHb+/WoZWXm68SP9yQk1m3t4EaWmCs1V2e6o/LK1U27Gc
C31SmOdi4Q5kEdtEtrLgCTEfNpr+HX8JHEk0Om7nuMn2T1K60wBWM7VQJcHxsnFB
mRHiFhrGyJQVlSqMiROMTtGrL20IfpXasLbt/MUbuGeKG7daW2buMLc1FoPDaMSy
rkI8TgMoSKw9/JMDsYt8/LNrd3h6zMGAULspAOSaiEygu8gtX0syc1820rLwMYIP
wncsKmCMzUt8kk9tF3QdiBaASvftk2mIV49cXiOjxZb7JaIIdiaEAV8szC9Ktvqp
oZcb74vAwfLgIpDFjb7Jjzw77G3JNAIFl6zUf8E1cjeIcw8EElAuL4ZsVCl237aL
r38ygcpn78zxGChdYIJbLx+6wETY8Xn2e6ovXaWL7Zw+Hlaz4ljSyZI/nZfKzxxu
FUCeMxwu2WTwBm/tjHhnudt26oChoLZsMMQaULR/IIQabub2DnvMT5qQsnamhgPd
uwE9hTPR8h5oY4ccDXM0UB5InxwjcVxtqhFfNOloyoBhQb7QBOhUbbGZhT2evV/h
Lf/xzPdoFueZMdKZpABYS++GHqN0aVQVHSh7oWqo4CwbP5y0gBNLCcPysa8VS1Qf
xW3JBZ7D/bg/HQjuB2iCNS7C1b4Me5mb4K+YU/Cn5pJ2ufdVzAwrVF99lpxFz2ND
TiJrdk6dbmh2ccz5kmzfPYLqedjCfTNRDhtdb366Vnfu+6y61eAA0k5M9wr6+oY4
PVCdNvhOV+CeSYxUVPzH+w/aoPa08PLuQuBO7WX6ArzkR0Mf1/LZPzP/8XEs1iKG
CParMSseRlnjzh0kqLbgnNeiwrZEd9WycBc9bzcYlD/N0lQXOEMt9EuUs0PIIlfl
yh4W10VoaGtmrFHEfCCysVIWbdY3ifHHEbUybhPNCrFUJGDflTJ70Yyeu+fafR4x
bDxXd9mULWDGv5cskE41bE9/Joi/40hgRvNZndjxBLmNefyRetKMUwVYeICGa//J
/FRd+cbK/dGf0c5vQeROZk/tv0EKj3IZ/NMUr3VdA/R9+nGdzCGmA4nj/0k1m2tW
wDXB8sbtBSEXUZhRLgaPRMy4Y6znlwYONjZBKyBDEF2+lj08noK/CRXjsaM5IDOU
zwDyfE6wxyTw1B6CLO2Cq2Ghez9HhgRvFMiUJCo3cvWO9Gi7IizfnIN8VJhSSMLe
QcwTwycrBnuwecM2oxlH9Qv1KpuZExZUT6Eey/UVuV3l/tPJXF7/8Er1DNW2MTQt
yOJPgE6KbDzFIf3yHovnGvuw55miB9Tj0MVQ7cGhU2PN6Gv2POffUQOB6aaxYpBL
ZrqOR00IYuV70L9JOnASqzj3AGISQYnycSy7ChDOADf7QB3Cx5FIg+8sPnAKIbPA
F5ybg5s7Eycvj8K8XZDBBmKQ6nEsCXvaacPdGGCEWvwpY3IT6wZ50q/7finrDLQv
qBt5rRYa6lqQFq+Dy9TOZ8kUbvDVR3WuYcCmvel66RjErWdiMBx8stibXxyNgnf8
Qzr6i8voDV5GAouZ7als2gJyIemvDX82zTkKcgkTFnm4HMA4zgPYhOy8d2rg/enD
XuS6SFl4REH7BEG5B7udaRYsUzSY1y4XX00K8LuuuH5JhKYASczE7ZpMQlzongWv
bE9CGdD8VERWQ6Db0672zp7ZtMKVBqX5EOUMFWFMvw5+OUz3et3L3a3H5XlnXVS0
Je/ah54pEvMQ4IRVHvTYA8y48j1b3oQ27dXYaM5HbUmMgSo0kWXx9xXIdMlSZPhB
v9ei7FnIE0CqfW8sZ144OisfyrnBcwkG59kxTJfWFBDuYP9FqomXujbcbZQkvQ4q
Kp68MkLS9fmD5qsIITpw0SyNx8rWvprp3nFs/pYfCc3DRDo5iRFA2sA5nCopBJhZ
WjPjUDa8LL6V85ZDQ6xHfBJJIKCpAEq4gzNBvS9nYYRDfanZbtJcdEdFKREySzSV
6dKhTSXQ1dCpPtuFsuIsruD/5shPR7xNj/Q8fOr8bXtE+u6Jr3dLnPMEqX0EF4J5
0k3D0/vj6aYA+EJ4K2LvisiwjiSrJ8sljFhhIyADAgm7HVTsqaOgMUJJ9CoDBWgY
dlXode3KczmdWD2MCDdsYhEhJLAfXielP7JxFMu4S/OWrmlULJSqID7ndIh8z7by
pzFON4gDLHmaZGCWNJ0cp0SpzuX+FhJWFuCB6co1xxvG/tYZQqqdIZ3LcQgUF0Of
k7MuMLDgVXljq6761MrhsyhTOb/QuD7fSEbMNKZDqpZnoH8fbYnEtARn/UYIMhnU
EJ3na3t6h0uWcJk1k8qtfk6N1Iyl4R9DS+QZKb9vWnGQfiLoB5CBLz47OocWbEP9
CMBJFAYZ3LWM8WwlXHef4/L/yywUMyaph7rN3jr0tlCQIOjBnaMHDgtMt4l+K53f
4RlU1ev6O5oN9mInE5LboWl9pDmBSYMsbLXpNtcXuyHR4KQqgRBopKzwuCe6zhE8
sV6YTettCC15NyUv+AoiKrseyERX5xGQCCSI4X0My2BPUQ6Ng3YXz8lKsMiBhk/e
mXr9sef967JR0wDGm3PffjYzi8p2gvyoQsR1JZrIYjPmYYm0iZkSee4AXOwJHa3M
4Hd17OCNoRP+n+pCsgyhEUrdqPtDCI4QtfW0vX9QNMsYidl2hT47VXvalOQj3IfP
mBG1hN2XKNu10TXu1zY1BRjyZnmvH4r/iuTqa8xbVpfrXU+ze7yGHupw8uoIeKtc
ShnAhdKcaHhOvtlJhCAsZ/QJPvl/MR/XsrNqJOkQh7izkwAaGXRld5GbeHk41vrq
g8VfGxH4TcVcfjQAY84Mc976nzjGD0hd0uHMXaGqW7JSs+DOxAy0awCiY8Ypt80P
iI60Xe99FLG2Yl0UsF7uXlZfaQZypcL1vrVKmZ8a0zQv5p+X7IeSSHSOyPk7Frzt
Fintak1rR7KZSCxN0M03kF0h6SoxPFXNirqMZH8GkVR5PVc3xlt6otySwG5kznA5
fpOODNIEob+4kCOoMrVPnsQf5o8dSOGAsWpJekvn6UGEOILKk087T8e39Vk6UkvJ
dwV41bwUrBaZ5nLsm0ELLQv6NKKrcaLpXCO5yWY1hCdcVqxxtvjo9M7THynU8mbd
krKG8N3UGqTU2H7fAfPbkcUGXTDRNN01PE8twg/HnKIfd/4Z92rPaMtmhSSe2cT8
GZEJsGGIb89WvfkehoAYN2UhFKn2+TEkhQw29OmbDGJeBls1n8bBoLAQ8RAS3Qjs
ImppcaE5l1/WAbiU+TqWsuvzrYDcv1hyfcljJLDoI5RjvV6SgX/NfulnBD9zls0I
gYTmQNWltgFCgwU2W2dOiKbE+Zgdikp+bqXrCzku2v7UH7viCAaL+YJqhweec6h5
sGQuoSbOpmRC9G1pNXwvVTVfiijtKGQVsnSWogzP0CwN7Kzx2s+xi5RfUYDWEY5s
E2x8OsoGO4m5oecuCvXE4iu6ty21hHlZ4WE3Rk/kem6LGuCD6a/Mhyvv108tlSch
+knuxFSmFH1U+/W0V6aMNCgw4aQQWcTI4OTWhn7MzKAcea6N2ITN0QvZCdv26P7j
LxjUoMjCTgEpr3JincDZcoESuZCpfTFJPcgyfLAhP/HsjGoqYQ4wr7jIbKU3XT3x
5nCtAuJwrafwqpy4QpA4+NvPbHwyxWcgGJuXs3RAFyfLjoVkkHV7WAO+5nzKkcfX
qALqlKkqf+zJlb5r2wVPlVLei3qlkhEid9NCBuf/jqAvWa/NlbTOmbuamdRyqlh6
e7jlaBe23xQt5JGYupRi/t8tYdy2faj82unHU2DqEICq4QCQ/IAFqMYCU9fi7cLb
jnptfwN4w17gV3vm2qa7N2P70+Se4xrZM61Q5Ka4gzGEeHabN0YEKY/1WpSKCAS6
41Z44Ehcx3kVUEMgMNNevb4ONUN4Fi7EFK3IBaHrgOUC9GI5E8ecAtqUMt6fjh2V
rE8j5Oj6I/PNjx8G7A2iio4G484ry4usqDyTDjTAbfKDEzsJm+LTiUMWTh41LXwk
ZIZns4Mj1ogwMb6bPCgAEXvl5jQ3j21Duu2WYFeg80zphvPXJBGwFm4FfhgEceFJ
VkktX/kSIHWTpnBl/BXyDQmdcWOYjpBYmBCkisBDg5r50OO/h1bREi2Rt+kgTod5
mbaXn7DPajDAo9oIcb8+olOSXlukHgV5zWqjMj29wzex4rf8R5QJB5ntKsUIWWvr
tCFDf0uR+OYDpfMLetc30v9JWd24ggcNB3e769Foh8PvcPu4UUpQRQsELO3XSqgo
2Q5U4d27c9M226e/3WhW6sRi/sGZDiu4YeLQ5WqmGrZBOxtmLt2w8+lDdZd77mEc
vbFImOKp9eVp8o+EnpAhYZmWPNeqtaxLesp5P3mwTPGO0VJ5FE+mS1XcWEz625LH
JCMpgEGmVT+9x/YtKZJjYA9E5A5ahs98qoy6tj6mJpIFcCxYLvo+aQmWX3wg5zeh
yONFynyNNCbh1/2kMQf2qlgjk238u8BuMuU6C4WCRy1q8t0lUldiDqi7iQbTre3y
/EWMm62MgqXi2eBjcKq8Xso8+ql+95NjEyFO5UqVDnXIZe00ckT5H8S1xqZKPFhP
Vbep5ZM7/ql/jLRYPDq+8nFx+7kEB35ta0HgeC3CHewsDuFD/qOtamTj0LmA8rdQ
ENPMl+MVZojgWr+0pCXPxhEUuIBesJKuj+bc1qKECQW+vCn2xQy4p3cdTn5kH9PB
9WzTt1/dYcfXbXSn3biZANWixnSJiWvtv3Gnejy2MuV1ZIjO3t/NRtN3bvKtnPMT
84lmOvk1fabHHZO+JA08HlhHZ6YMZAVxKJXF4NeVbAGlGzN/cRXLsssU2PNFc4Tc
sTDpJWTUWQKMe7EhgG3BOAeMwD+8zNgwJKhYQCE8yxPvtuGPBSjot+C02F9vheCG
4bWOnxU8nmSi57dKld79yaBztoFxIXa1YBABpq+BspFSIx+yxUzrtHpxThJtWdTj
GWgVkikKAHRkNUVSmIw2epebfApZrMtGVa15U2rOuXcRI04dlyoOYX4opisVoJ5h
zOtoLLleUTzqkggpG0UnnSITkqHwp2DmSEYe6s5crENPISpdlUqEX8ud+Kb6esrU
dQQlKJy53XB4vDFA/RoI6snCUjEGVe1OhbYL8lCspCOGSxY9fi5rf6XFkvRe0v8R
VvGrv7c0O3kd2hvPv7406JVAcavyVefH4a8uRH8QHP7ZZ3Gk1ruiOM0RrTS3Q7j5
/E/o9DZd67UYsfiV7hFbdHpPi7SqeqpWoduTL3G1a56uwKp4am4uafjE0ZPowQKL
8C+d45TqWcKGZSFfgk303pTdeN8wFpjp4ChbomUjfGTi1JSQAThFmkEokEvvyLpe
guXFGCrLgnWZuPHVLc7xXK+v9hxpDU35rm22p9uy58JY27HfxQxjoEb1XOFjU2BT
+t/En/8Vvw2BOY8T5/IZEwb477hPAmQxm5lIOTCN3nA1GhmaSzXM7tEMiS68NBo5
TZx6N7GSUFHa9DnynpVZqlDkka3W54w7DAyweV1BaBcYaXxzgh0i/KVcLugbGopc
T4zT0OhxXI1MV1pmTW1mnF0OkKM7s+/JXAmAghgNpidgZQKQNJ1t1nZYHUnvmoqz
e9dlCewYdGSjnwjR80c/PhjBpi67a/NtMlw+PJHP1alOezhMMTUneIwRAu6aZnkh
LA330cMINkhvIFgwBFuXVLoP+kt8LuelxHbGv32WXEPY0qGOy+XLemgmF4bq8dZw
P8TlCUA1nFuGgWRH4mgNwGFx4sazb24NXJNFuaK67gip2hVzWLDnI/JkQ+xan71v
yOhfwYJY+ZgDrFrHo5bbn/RUL8Ky6+BcoYJjvZxlHC95cQIm/qI2tVkIzoNCpT+G
YUxdECy1gIJ3Ev5lRcbnZoA7OwR06WFHhTdwX9MqzyO5Mj+2/B+MfLdiNSihtZcY
iOwtMbHrFzHcyww/sTuy5lReKIyPoyYgEkJjaoDV/LOE8KD/N+xZo3XLYrEu+/l8
ww9EKMY9ts0UmjJdP2kiBRAOzX9O8ss55xHTGw00R/J4ZjJdV9u+fmllj7Hjf6ET
xTQ70CZziKYJ0Wc7IACvFstAbDHpZT3sHpf7mZVfwBrimyCd8JeEXn2dB4+qS5sJ
2eau9kYfD3TSxsQJle0wp+Z9gFHsbtVRBlPCGPVfI1OSRwmexPJpRkYXabkLas28
iKuhln1DnEmE8y+5ga2WFylOn2/4ro6F6THuZN63RkUiFNaU9tBFwvE1hGIW5ry/
Nj890ctrEP0q/z2hJWPRyo24pD5Zy260iqg93kAIIg4vssszcue9/N2at4Mo2aIr
+vyyEyzkarWpdxwgLEXevfyEJxQ8oMkRJ2I54l49oYzFaMQ1i5yQJXaiUVQ800s8
T0fqXnvQYtIp154CQ+G4szTJ4S2TKCF4Jdl2pGSh135VvOtJ/4RCftFAVmco5cNA
La968FPe5t8pAaRM1HnJ3ePL8YqDnEhGrR1bUrMidPMPVSBk+BssGOCTu9CRLxbv
TCj65R/BCbmMCn0aChTK3TF0OzPDPm9sF4wg4e7+FehKOC6dS84fmtna00nvs3Qg
7+8uwbnQ1VZtjY1yRWtpHk6LVzLEkZZtRX8/Dybj/XdElJQSi5Hr1WhcWM+eRE5a
vP6RqJnzTnOUXkUScXok7kIf4OfDlbAqPSYKhPtdi5xnZDYyogbSZ/YXVZGERQRm
ylVsTIFGK/UZER8wioyC3wKed5MCIoEcjc0q0DhPVI3fSgtE9+nlOCv+JfLDPoEL
cpv7BLqJoHNW+gkb9yzGCmi8vcwdEc37N7LEM/fI2N5qBi2zCSv2EZc2HVCoBf61
VccnWb1GmVO2tOuGsntXCwDOCnfyW9vxGCh0i4eGUBWAXjhSmKMJG0gyghck7NW0
TxB7lhtOjLjzsUNS0Tvct+gJgcEzYAMZsLlPa6SZr1rZfNML2+mcPaBfpR3KtLTL
ho5+xeDjdsM5BB+lEkQRt4wX41WuGK95m4W0oizUFtGzOzha/fb+LdKyIHxgoebH
r4w9DlZrQVhviqQCQPb+kqg36jEJq9xwA+2j3rWzChnNkOdliJ7DsH30M7d8hX/U
CfF9uadaaV1231KEePVgCB98lPb5G648InM/Uwxn93Iphh/QEc+YNJ0fevlDvt5C
w3fn7r+O1NQFqaBgEPyITaL6zGrEdz0wp9pGIRFIZ6Q4trKZNX/D6IYtdeVbO6rj
khdzhIczeN1afEhuHKz+DaOgMMS04xbZPi1ZFK3erRPQO2RQsHJva8wbxc5KjPEp
SFfnLq89J4VvuRkqr7eO3o9xp1t+Jc0WNym+5vbpc3s75CHqSwn8FJNmDurQ7ayk
1HukT2qKigVyXjrfM7nkh1OT//U3dyjqiPkCORa6G6nZCThF3WDQbIlh/8IyMBCK
7KY3zCv7hqHNHjSFzL/lJjdrN88rCAwFMgqxT5m06icuEnolt8+2FkMLbSH/N1oE
e1Glt5RSwoI5OlsF0230vk8s5NFLDVWTZGx8x0ygbziwWHhHY+oWeYiHA6Q3SGw4
PESykwep1ARFlXoCysVXAzbumHpJz/v+moJnlY6po2ntpFWKH6zOhAbzQ9+war+g
JolLnO67wCzqqBKYmn1n6yuqM7E/9YTt4bJwioXjc2HYl90XBXJL4yHL0mZ4ZFU4
ah/qWwZZrTc49n34PbzwKtZ/shfGREVGZGRXIxhTrpz3qnngoYZVeYsC9l8AEtek
baIJ72qLpF+Tv9Dfq5/XG/mVSFbz8umncUljgJnJzqhB+bDceIGU5n2kS2kf6qQn
ku4FoFr9MK1zzanST/7aYUKpm29wMA4qaO37VjlLXLViNwPb6mTRQPvhkfzhetg+
IdlnmeR0KGUb+v4d/jmDala5sJOaZwfrbvD2S+oxQE4PpTf7ak36PAaa1xpoO0nF
Gq3JAaVTjswPDKu6dtBWtZANC67oHowFtC1t2lA7sez+CPd9skFXu5wCh3MxiNc3
UX7eWLDd1uc3rGDhMORCdUOmKwefwP952KX/0F2FBx/LuxfDiITlbOFUDDRV99pZ
D3rN59Q1iA+7nbG9wCIiLGIsabC2Ltbp7BsZtiECCybY90dP1+sWlxRQNzIUJGSJ
h0uKDmuyThViDP4eA7Esd2Plxk0ZbrsMBZnZyjar7fJB1eD9goWr5bVaqzLRgMJR
FxkDzmF8daY+fi355x/aw5Gk3e7SiIEooxQ4lCAa4863MnXFTRshvWHBsoISMus2
YNDnT+dBJCgnT09t88N47n/hvAg56Sn/tN5kYC7hpzEdzYbwZGKrgCWJDsoZ8umN
LIEq+ulRQ1Bw/8uiRwJEYzTo38nG6Fl2buCxrKnwLSpzM/feQMDrUGuxkbY/58ni
9fCB3fZeXNSHhgpaOJoHb3ccRGqeBpp9nuMBvjZ1nMsz1pk9dz8E81/fskI2YGUp
nIcPQm5+LyNJrdRqfixOpKzo7+zO/tBwPQ9/yptFjgFcpuEEdL1sAFvTv0i0YD/M
1CfXAQ/v6tj+6kIpHV4r+wDcJcyySnebvfhCo0UyXSKrSdruKacOFA9dyjVJqxCE
LGerI+ERSFf16NrEaV9HPnKBUo9QIcqT5omYta/j9ndw2OQBbZltMii2nuQGHMB/
dUz1Gvj0nc1HLh3sVfgcRFfL3ifWS+awGDlSUtKyV+fL3508S9nwQcvaFKtI9D9q
t8LIkNtndWADYp7rt1QlIAnfLfCuiiFTz4x+UDEwtyGq/Qs/3KnRwJO1KMwNnDOf
diQjT4oI9PZwsQvjyyfgSns7CsyFTYLWIDfRU26ny+rEqIjM/u0JUVYn3vT3B6qb
SOABgfZsnWL78UmDvh16M2nkS2TNIhcxM9t121t5DJKziVK7gWCKE43aHY902paA
yzgftoiwV31qEIR68pliPVYLZp8y5ZB3rgGz4BxlO3TODgqzMZtdDTqF4CvinaL+
PLWGCGsMrM3VVn4BJgm9Vw9kXhUHU/StZTbmwY1lB8WnDakQlDYQF6sual9pL6ZP
JZ0iqMP/TGX3+Kb3WJsUmqcwayl8D4HiXBaQM3e8y7uaqmJE/GPtXy+9y4r6EuAm
7atmmcnWH9ZDfsY23Des/MPzQ25E8pL0ubdym4kWtACLFOsrtklbpKjjYiOdcMb6
Y/OYe3p1+HXQHiSSsax2EKrprlDE6QZfA75VIW/B0pAKRhmMsuJspWhKf5ZNBT3A
tNdKzOxri/I71Kb80UBCtnC9NViqHqpPqHCiHHZoBNGo3SCADVqLVlvXxReUVLZ/
iNi1BT+G7gtVJ5CHk/wQ1NHR2mYH/edfL/mIXlCoNGre2CX3HttGP+hMjyUZTJOt
HEb07BwLoE2FQL+xZ9VURh8QNuifNC/d+ADIUYmaI3tqPNCX2YMv70OEl3o45Ou3
Ef+2lALDHFNOrD3PgKOJfF7TH2YuWdQMhAknu7bmLeBn6ZYUF9XT9A4ZT3AXhWJr
fHWH7BwMo0zRLGLvQ7806rFtSWa3FZvmg8R+s6e5QVOH9pn8P9GmMXkhT5B7ltmO
/5uzN/dBJcm350Ur417BNyZZblUiJ7cAEzWgQ2WU4c/0bQ2pH0RrKZO3Q1rL0CTC
kssblij40QN8e9UfXrq/YBUb8LnGFf+v8GU0c3muEwCymFWZH73gZ9RralWJnQ5E
4Hy9bUZtNZZW+UgOLMNHrC9piZNDFPtRC27JfwLJ1xCUkoNS37RsMu/j1nU2kvjk
AbkqnMxKxGpImCbTb2mNYbwURTB8aOk/D1WGbhSTESA05bSfUgxY5IFuz9Pc4GA7
/mBjCRSqJ9qn7rug1+Tq8XRKT/JGJI2u3C8P16G1/7vncEdm/pNWTIMLZGwbFsKU
yoYBLTN/OBk7BGU9eF5cvtnZS+wPRJB0PSX4BBUAFxtm8QbQYuictjxDKmc+LSs/
GNqk3PuRVWydO7cN/AijX9zy2gggRUQl+zd7EP0/O6s5frYwy/sIHZ0L7ZOXEAZM
1etFKKizdy4AnHOPLu6V55mVhb0Ox0zZw9EpVvGB/EUSpyRK2FI9haH2jc2MYgDu
UJqELdF5PElewa4mXvxxDUhJcSjVd+E2nK1gQDF6f5LetNLfDoQm41KnC6GkF4Oe
luDucALf55xNRKDq9TiPb7TOs8FQ9w9lH9Ug68Psjy/u2j4myVjwuurLFVkKDdcW
dBG9MZyHgUME17rQ59za3diimGbBc1eOZfVn5ES2b5IxIR+zPSQzAepbjWywnjD5
DAWrKO5l+g1VhPKqyh3b1yRWZf2tDWtVzFySLLuWXhNMJT1FUtGHVSPV29xGuGmr
/+bAK97i4X/O7F0B4V2nPLV6qX20LZd+70ppL8E9jqrA7RY/UkOUQxf3BYWTsEQF
lmeci+QdFb0dFfSAcXI7SN6GDdAPlEd4cSP+a2zoGlgsFhq2c2dBAblJYFrJrL2x
J42wbpM/1Lp8wtipHUpekn8rKx+Qs7Z5wBjYj45ER1XpoBc71i29sQKKedYwNW+y
7UCqwey0cKOREA+F2BnoMYRPt1Lf+cbusMkoxoAdstp0Gqs5v0YpLVyIcIWLTzED
m6dFZZZ/8s7d5gvs8mMzX94x28XT8wj0hUeshiHtgKr+Z/dXYU+339QjoayE0ERP
c/8WDLNHv/ogkXeIanWsXbIt7NLuo5/Yza5MU260la4QIXGq+fTWOaLIXraH5hWc
lQZe2WU/Qcz200PpgSEahckhl9yLBipSk4MRLsbU4+KGd3pGaUO9jsyPKTtsD5sG
wpfiyigdppD5m5jGs0gU24xYQWI/WbEVt/02mwz6LKRqFNw9rOU5Hp3MKEn+/Aul
J5CCG3pQMAdP4+I+i5OaqsDXM6lRQXswOToeoyniyXF2QuJNIp8NOOOAqD5sM37j
+kcEcPzBmi5zGlkStmOgnVntf/X7m4UUE6muE1eY0u72949GMJUcTzV9aLNVa+Sh
6Gi8s+tV8xlDyeC1DNRgMIQ6fCxuhO9nS2ThNoPuRvwbXlGQrRW4Ydr7/3U1e4iE
rWoDHsW60/HEHwdaDIMv7XgchALR9iJ2qQSfxd/tzHVsJyCzFXL9JvzicQmhgazl
mCOO/EQYetasAuqNgFodao9wSWuz07q7vK7pww9oT6bCZOR72Tg70AfN7TxFyuvI
JMQ9F7exOIJQnWMaDSmjB52V4sjW8DZls4WWOyViVN6Yw+WstvSJUJa0FhMdy7Wz
LtvmHoCkCw3Jjd1IV1ODJPUj24Lk8DDbS9zHxRPRIpCavo9pDtQCdrvvQtG/DI2k
7EaLEAyw3Knz6AyW34pMKNph8idexRNAMdLXJpfog27+Qo4rclhVZrBjktFGFFOw
sOAxicdy0unRftkTszfzyZsPksLPGTo5N0xXI73v1VoGWxHDjy1zTlFpLlWMzBy4
Fb3CsNKwkcvfWYbTwj0hBNDNuuAD/l4nwM/os1xwFGf3cRMgJwfIMzOE0aRoWOb4
3tN4bR9pnEiIy1V1ssV6uBS/xtwyrl2wJ8Ux/G2N0VcXbpJBRjJe/9/wPzbDguiU
LXO622QXcPz3bYcd9vZGF501yT3p62jbCy9IDZi7iFrpbjEU+zeNJymM7Eh2DcjX
wL6/dd1bsL9w04zzCxXDF5EhRVhaxMSn8j7LUy3SEf/O3914wtgC0TZfnedllS8Y
CNBSMjHiQ0q/5BtAN+e2wCnlC5UI4/EWYw2B7t0YHsnya7Hwt0GPV5GMTVZMqoQO
F2QlqlnX9Q0o5CZGTotVkN9wk/X7LZ+O5TAu79puiaSgGy65oWlVga6BQpFLNHQE
HMurxFkaTrOrrlRad4UzYEa8QUtXzwfDFSq7Qk/nDM65Ahfx0eCZuXvP8dZHDawa
blfPKi8tls00GTK82kgV9e0MgxO8y0QA8AmXCVUmLKcTFtNkgwGFXxbS63trEm7I
7x4aaQHxJyLeO+AgQAH2Tl2QnCdbARRsyMSq9hMlLN0gCGzjo4rvcEA6u+07KI4G
739T5tZcEmWFgdLnnvo8BSMmPlxcrcGTaE+letGu50VjPbqGXouMtX/m/nzS6I4R
U27cgsBLK+CmFG5wKZH5Kv0qUZxOuKPWn6oP3mSZlXFcFAy/9wOGTS9rnpHfIaIn
WykjJu8olGprPWpRLLIw48Ekk0BDg4GyXtjP0pN+gVpUcjtTAzeSOEObJdEycSan
AQQvzE18zE01erk1/bm10mhBSnmvjVQUn8WFpDgM8oL+5Fq7XL1Vl0MxdftSL8IQ
hka3sZIRrFQgdWqYa0v013xY3CUfygRv+i4AxySrLzfh+LbOGng0zKPff26Hz5At
SKrRpF5mmLzx74Woi3m3ZGAp2xDpGjgBIN1XdPqIlmf1iEBQA+l+U8HHou4NGL29
pvCSsiZIQvg4WzUUgBbt7n4TxRixrZoWGPrr15gybKQsVE3riF0/xmI8a3NMIkn8
ROA6XhMC/AQj4H36kidblYKqnkgdlgH3Sy9lkPX5dvyu0EqcI3jFq78ZVR93nHCv
c2UR0yCquZ7BF+66kw799rpjdOrjzXPu9vVRLcNI+Qf6rrgoNIn9/MT59dR9HgQB
9z9y6g2EznM47TXlrpPe8s161Kfusvera+a+C3q7+qzgEDHKO8BMpvc0cuigrEyZ
9N5UdIvDI/cozni59Q4ro+uFbB6kLu2pvia7/MCP2G1Y9LYTV5idqyR5ahT3tKSe
hBboGjq8rDYifU0oJ6pdY6qW8EFzYWiQ9GB8CRI2gF6M2Bhh4HiKVbf/3soUchE9
dNWuSsKDYscSJEu2DQDC1vANdalq44I/JsbEH4kvtxs37lhTNWxoF4Rzkh5KVur+
2fPFXLMKdlK9PspEhNI1tYGYbWZsXjOihcpgv66ug3Bpd/gYJKgQlpsqC37VL8XG
//290QaLhEOEy8dGnZUo4aKCK9+pLrXIkvxbXcTN4MRfq5i2YBVSenvF0GSemxQF
vGy+YWWT8/4gLr/rPeGN5mzFCffQQHbGmFAl1KWy6duhyzVhImndSN+ndgYW27it
bABtbDT47Qa77Tto98nIGwRUMEBPb63RFqAliGxlfw9bWZWcmGhQ1JTrgla1GdFv
j1Zk3Of+W7jDqCPriao7whQBylP9XIwVUS8lGHtmXovgG4kdtNDplcTfT27DnlDE
6+BEHjnC1Q+lRu6VwdZRfKF6wbWdkvPH0gCgeSe8ZAv+rAlgYSNTpANbzHz1xr9V
VnesNlgT0pM4ZNEu1QBzCsuRSRAT19Bl0yFVFcn18IpmtT+S5UCANQ2otvp0u+9X
+7dDAYUknzAE6SUr7+1pM3Vo2E1btd3B92LhfBHLvto7QpV8hFWbCADkg8O6d76/
c6l3x67IwTQWVB89UgiVSzaKq3FRSZBqFODgkC8wybSRIplisn5tqWDFSPRKTxQ6
YQabDdGsOKi6qRXoLYgWSCkL2trx9/2F+zFRryDugQ8xCuajlSD9O6xVzhW9DsB8
ExdYSXwoK9D37h9XmYmDxdvbEAg49vVczm7/QtC32uAC7fuGUAnuUBt/106Upad6
6EuWqBc7iln5B4Kpkj0Z8q0wn3y0gBQejbJqvscCZCRMjFKy7EuV4XqIHhrDlTxD
+8dTq/FVnvvjwRQ7D1kMGe8vXrv91UUoHGg11ydhLp5TaUZi+GW9LbuQXhW2evqE
7eQybWGIszE1suaPIkbXLPDHSo3oT6e0cJrI30gJcxMFSLOPWe/qs/4gb25zDQjb
dIBCoNKOykcExJ+ibf4vJeae4K3xT6hfAZelOHPc1gCgjHxJWc1PoQgY588EVL3a
iVwLEnUXNME0bLeImRIM4J9Aq4RATwlPe9yAhpNz3GqaUrEDRIlYMOoTZ7xIyOwn
P8WeGx9MC8ZtKqBz6XWTfe/Tuv3sg5wZSHpHc8+/aRDpg9r7gtNDmLW+mmj2krv5
ODchPGbPKJgIEe7yFB3vapDfso/knSnBazTBTUURFfeMLDBmUXcAKEmLb0oAi+Jw
zNHvDq3rf3hBONy9xfPTyN7AWUuNY1woGBvtaIbxKzknUtD+tqts7QOwiyhpBR9v
uIkJagggm95xNapqkXLs9A5xzonTFuFIMb6A7zvpYqMTwerbtiQmyf4a4zZ+Gw0J
wfuWpPE1qDT4MgBMkLO1FVScCmkldhucEw0HP1KkIrSjPWzmGYqnwD663FafC/OQ
k+LY0O9s5EPIKg0fi3AOj0y4QfUSyt1ZcykWsWEULBRGzQAdIGYx+GZhw6/e8oJp
FgOVUBhKMd9iUkP0cBhOGEZmaJhKzmhtM2btkO5Wk6V5XMiPGus+PlMZVnKngZP1
02WyUkYiLHeyfVHgCjsOZHnukMhsgqUi8d4lDsch+n4JYPAnsE2LOlmXL/OcSW+V
HD3MUS4xRexJpCw4SCakAeaynpXgv69AY8uxd6ov8x/Mvby4/XIf61mF0GnLjXEM
H2Mmv5F8lcl+4prkK36DkZtCuz3RbayzZHhmH/gzm3gRpg7FNAM2gutvI99RLUai
9lUv+GG5gWj44/YhQDrHP8H3Rupy0Vrpy8Ziz0XzcT+eenOeNBp3gEgfLav/apjY
gxqUGrZJcclxPg/4am0dBRvs0p30zK1HFbCETT0BakLtwyyj/v+YtCjdRPt5+R2P
Zjh72ZDl9VmRA7Xgin5o7AHTZ6L5w6eysgLI2OMpVLhcrmesqHy4ugQ2qKk94yQp
Na3o92zL99j8hIpDG2OXUwAy10NkQk/wumMiZZ8+KnRgKxQc/B/6ravdmyp9cpyS
bv3ticYeJa/2AxUJFwx7R2cZzMVzVQj/0vQOh9eg9ZbuYo7erHVQC5VXrWtPa5Pj
oBPvS7hZ9BOvVQ/LyAdTPwijVVWFy0owZHYVJz9DJCPEcsGFkmPw2y4qOYZoCnCa
JqWcpphMlgh8/fmMjqewDKQ+Cnwm4RBGqWQsCeeWI1nuWPICQb6ZwdD0Bh/o0TPd
TL9bkVNxzQ5mfjJl6e/DsdjPHMCTE25ug8hrvW8FeJmmcS2B2nMY+04NkwxTUKe2
kHqN1bjAgimbTpKn5gIOWuL2CxviZQSD1nyKD/oDZghIkKhoHhS8d0BxDPcIYzt3
7nCej1EG73kXgHtnOzVlTK0obtGtVou0bSg5pafuRuxSBdRmZofNaXy3nnJZ8OCI
GhqLolvz7trcDDlnDUxpaKKANkMdMmrbbjxF6SdDf2ym+Ab8P0i3e63WJgh7a5iv
fXpwkwKMAjctYygJPh80f+2DWHrMARbBPHNe9CaykLJioBubJpSJuR7Kt73X1FOR
iSFSyCcrY2Cy223RTye7nFN6bQFXzH/KX+6TJqWSXzp0ip99wXQwVM36y/uCcIfG
8ZEmVSArT6YojIjy1ylTyDd9sbFCw2e4sUDe+UiAQ9e6U9JVC3oIA3AA2GSr/pO0
l6KZj+MN4fwGe/gIXQBuUbCe4kAP976CKpP18tEeDazotSd3KYFq5pJbC4i+a9mZ
DfipFI+Z4Ji/f+qUIGGypnYCdwluCe5Ws1HPLSS7XBU9K1y59Lnq8UjGIWDtYb3x
/bN+Sp5/8uXjcGrd3BGXpIkvXAiHZ3PxkiYnNBGgeAfi8E+JPFRHmSBW8S4bZ+NP
xeQYhdy0QeBF8BTbs+Lhwpoe8xy2K+RXvA4f1YSmYJ1So3DXARAvcpvCIxzoPBvG
dqqLSoIqqxTvVXCcyv++6wtEJZogZ+dIDS9OVcfNIP4GHdgmp3AFnWRwxkFQcibz
c1zV1l7xq1lOmj2h7B6sCXAUDMevi+qFZXHHSVCxeNvaQ5O/ZghRtSJ3iOSfBkdr
10gBRukaeoozORDmI1dMjmocyYK8fDjzNL5a8R11Tg6aMdGPwmd0+dfrkSah3FRl
ckZwP2H1Malg4ioQ/ZS1JXfkhs3YIXnMhY11nz3JjUO+4wImGt/0Ud32csjTM0Gw
qivuD+2zbDsCHIM3Fpr8ANVPJ0XmWPs7YklM0GrSG+WVOtL6k0Hcnt2qiMVdZMKt
DZBdNiKJ2Y6xbpsJsGw8slatoMq6c0rfCIB/+AFS3alBKBFpQqkebemA9ZEEtrvz
YQ/SBJ/79MAWuLObF4cFWj38zsbHfMmkIKQUuJ65RtpAEQOxj3NGgBhXCO1T7N/g
AnUe+dUOnWFqLCIKKhhOLcztE5OMoOhlz5g8OpX4TuZgzVKQvfiCWWqSkCjv9dsT
8fMEzUrj5ClFkGGdpL8mxuLIuLqRUfs0d/uS6ToVDgLi5P2jkUZiMba86Ex/ZL32
Y+bIEotNda54NyjiBMie3L9IRgyPUXUSyFvM/96HDc/D286UQ4UTczFa4dyemhkA
sdtyDuAGtfp9pTkIVrMHCPCsEoNU2isFNu84036QBtTudPQ9LsAKKysvlzIOlhLD
cbR/XGSYy5QUwQduYdSJY2e0Tn2jSxtnvEweI48TjZwffysyf4mILNNIFLW+zJwM
x6HwWDOqEasu2NsIqIl5TjVdEerMOW7dfQZDUd7czBJgnQEewQtifZWO5pL/+5LK
mc0uqPtVN0TxoDoOfmXDChLvXNdTmUT/xCQMZ4ifkrcgklb9R0OsgD3T+65z450/
74wJ17KP1JjZ0xXiFpBjqiBgZ9W29dUIxnJGkaDqx2MWNtHsNOHzrKDu3BnIkCRa
fsY+T7FpVGnrJhiSGJFUF+Z9CDt9tAlgkvh/qIMkzt5uqf1of4X18af8Md6h5W1c
OlJ5TFMzwZ4sIFYrldLgnH01t98Eu/3hqIzaGfHDAEBZ2CCC3MRVcmvXkYCY7+ll
iGxx7A0r4CKyWWe/N5WZDtYP98GnB/CfazsxbOE65tVPsFVJMllQ5bAg/SKF6kb6
kEAYhqpBpbXVreL1saMXYqu6v1XI22D3r16f9u4bOM5l2EN7PmwAe9LCMFQ29Rng
UgAfdz9JK+kI+PBV1N5ugX7b3dG+C06zQ+Pr7GwCUYUBLsuMatmw5yE/2PFKkZ3B
FMXtkg9e9XalCDfsT6ySUPn0ergM8SXr2q/fbMDqXfoWQnL2ooroLyf22IlfkgK0
N+L4LZJsZCY4JVg2rGpdlYfcamPTLZaIdhi8YvEAeyKL3PIN4ftZY1cs1vSsaxQH
vNKWQyRVmM63AwLGuBycNHyc/YpmshR0bWN7Ao0NJht/MVguXnfxHRRRlwyRkiD5
HrlkFbWYH9DOb5nhUETAvF4vdAAVPm+fmv6asG5rUjPAOScTSBytNyqrAYme/IYl
PVddbkdPpnaet1Tv6OYc+6PsnwTbAF5V+o0VtZBN5YfISr3LKy5iKiHhTbrranY2
v/srx2g1yhk/tyJjIa2ttczCpLZ9ES1LgnaB+hYdTk8ffSOJvucGwyML9EDdXU6X
LpVDPv2gvTzTj2+KhgxjeR5IB+QY5WZHtwcLbrdios423J9l354jA44p7nmt86xT
ISoC5qi1mXt+gKBmggzgF6P73S8ir2NrrSlC5AiLdpX6GY+29fmrJTzPA9zWh8KF
81RvK9mI7HY+ZsD2VMkpuB+LTuVIsbou4krUQs/dL7jn/aXXCWlRVb31Ph2CngUY
bFy2wMCLbtvzKqkDaAEhevBBr3Kf3ifNJ0QxYrguiaPpv0uaxLGx67TLiLI/rxyx
m3z6XrJTwZ2U+kJMRDhkfMb5cxBZWSUTGqUVvTsaezZBX2dGVR1On//VHrZNao3e
DP7ihwXbsG6jtb78ZkeGq0AdmtvfKG4HqNbtWoyL+4vYLuv5LjHgaxztOUN+M2fa
PaFS+cZYjjBdXdseQh07H0tzoHdjCvV1hAzgSK3LROeu2/30TAJeJD/yWJAViaT2
r2adDnklvWEt/3ILah4ccvqH48ssnB8TxNTOwAr/gV6ApUMOFcBv2inHn8zy0d93
noFUEnTC2vsMFUaM8JYOPJQY29YGaM3AXqqnwSxVdOPj7WsBpFKyAZKJDMwQaYZJ
hiqBiufxvZnNZWhDBSRAPNShT4MFGtpXcq3OM4fgeBkOGEovdTwlcznyDY4URDm1
ZfMp4iiDpHE528BE0VqDLisr+RimfzpfK7bGhReZNjQ=
`pragma protect end_protected
