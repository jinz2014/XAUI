// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ov2v8ZHXwwhlNmF44ZTDlaZSA1pL1yS8DQa4OHcifpmhrXlH7JkI/spz5mlvdcZX
KcTIwYZgiKtkE+tnPNTumvsoRWz16g9DzrbQNQmqTNx2K3u8lOT1GlEZYKbo8y2Q
wxRwJkfPOGDQkmD+Yg+riv7phSNGfDNQIUpvErV3fG0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8944)
iJtvUH7dFmasu42aQve4WsGLV7JufqcNW7iFTniiytSaqk2fY1p9oQzrg2xhk6cW
ZFXuEUmUjuzH/nR3iT4nGz1i12NsJD0bw2hNpn78E4bqFC1fLYOSRJDUBVYqBVne
MuqS1soUb42ILWLPIusLX3tbd8HRx2HsDIhkPBhBlIx7FitbrRo2RQvNNywVVAU3
6MFQiClqQXsWi0MpS9MPV+B7smF+vtCRYOxv3bNcHXodh/K/KtfCK6MV7yhr5eFo
PXHhcOGAIJkNlAhFwx0KAIfQKPajYQngqeyclKbJ/Yx3JBXqe1nWjf5vy59ITGIf
G+qxyLqekaar/6KrYorH+1SPoZRi7gI8h4BwuQkwbHkhL5ZQDX1kWNYeBnZka3hM
gc2clDWEFAdvRQOvRQfbiyfCJUL6uZaWlgAIZyGOgFtBy6oxEj2NI+msrSgdKqeB
0V8PzCQ1EFeYf9BrGbo0o0LAz1xbo7fZ1EhHdNepXA5nhdc+LGM1PWDfyUPzcP+C
DmllHBeJYm/MM9PIJE7o05TOxcGfwJXnRWoLbHVGuIZB9hCsmIPt8e8gFN4Oi6Q1
mmFuKOPR5GNd6dNq2fSX+Yrs06iPcXuOTwGVqxAHqVOSbj1VVd2kH33IeO3/dFEx
sBo9l5inWOrs04eQRJcu9Zkt9MQCZedmEU4Mm/9y8SZCCSmnfZuj2kfGApdBBQLt
jQUKQA/nKoAJDlJXtvDzSQeogi3i1ONapOl4/iDa5zRkMLoRN+1ZEWseVYhJLaD0
+0dcBcZQpdkj4/UD3ImSm13ryNklk7K7RT4P5PytyEDfKBBKhCAb6n6p//bAOroS
8t+RYBLBBsyG4nsJ9OwQruFNfI7CZU0O6a9ZUZbOEUWqP7VM+4exuNtqtTTKZleT
Cf5sCZNma17KlOYwfQ05aRwg4XRpI+Y6VWEdwqEb90U38qBpdl5+cBPEa89HCzKd
YtHvd9g3qQXHtvIrFCDRlu9cs17qZfUp2BdhB8ojOUfd2boFDJCAZSXZPcaWYqB7
R9tdh3S0ILw1AQIKR2B+DQH+0DnP+g6kUd5Pdy8lpvltSi3e0F+FkB308mOfPEse
BHFk6AgDXvMZy7k2c8JNBnv0EhnFJtmP6MDzbjwlmIyDcyYGRXxCyr9HvBxkH8BJ
b6TLHkGYIp0HNhuhRH+oWnEdzxS6xxjbZk/YtA6RIztOCIldbvzBnoCQ0GqipTEf
HHpc5vy41Hn2Px+OMbxx+W9iPsiQ2LBtMi/sSUsa5ZAN0RQIBYJj3L1enrCI7CqT
CqWqlrU+Xto5uEb1Xo5ZiIJKvoScyapUJGAxoZHyYe12kS+56ih3k1nMG1EJwsuk
B4f7WNGujHhQKqZdUX9ovnw1yCdAwIK7NBdijZ8rLRkSTXnE62MxNkHMrTYrPBFx
jdp4jXGu7w3qmOp0nocAdWjvYp5gb08EetTRN0ZFIGBwcmYTVBOiDA8irK2fwXHF
4ipm6fMScTK+VRCH6vWS+J6sHPqaRG3Cl0cjhxW4kv/BtXv1GkArIP4IMbREK4G7
kZK2c+ciVOLs88K+8FuyYtLBSA5Qk6KgZDackHIEwuiEyjKpk8ApptCLqZKgmgHo
byMrhxpHQuIfNCTae1d+z1JkStQu/cVChF96PVW31xXrk+RtGjUOtKdPEU8ltjQU
589CNolWAaBECCjArk1kPAN4hucA+rhbx0sX2crmPTzKLph2AuqAE51vSoXiNFCU
2/1QKyWheSyb1esm0WnZ7Yg5xoqBe2Uh0QSLFfk1/+2iYTF3HrFFe2trutaTTNVv
1HfUddLxf3E5hsm4akD+kOFTSE7s8stCdT3E7k67ykv17T6TT7dcVOTCPqqawHAf
deD6ZRgDyNlqbFbXTTWYOsV43J1X5eqB5cTwjWnORzf0Hk2hqYQa/R3SDaHHWPLd
W6ot2O/qg8WTIXu8yUlhFd9O9yoVRTN2qqs+xaB4yZUehUqxNB80uabI6HL5VB7/
z4ZYTwQFNxJt4T01klFOFj61+QnAzETqvVWcM1wgtGcvERp410rMDj5aLF7L/i2t
HTzaP1DBYSBPeJ1F5LQI/JO8JAVpX7QdNadR6EN1cHn5zWFOJAFm9tpJMNiC7SDv
eOFD1SWlYBFq9zUOjpEF3cyIoboBJNh8Yl6QS7Mp4N1sj0iZxEAwBym1cbSsqV+1
z1TCnA4suqEIoD6QQ+khbLwRlznxxR+WPaR8mkmsYsKIlDnIK9OGdr7thjuL8hZd
qbW8YMNbKhURre00BGWAzRLdVwd6+e2f/AdMNEu3X/AhAJptvG0qtYm/D3uRb5y+
WGM99Xt1txWm4Hct6iJ0pc8FY+nOF9SBZmJg/rs7gWDjve05Tu+m3ScVzKZLgXFE
ftmHtBO3VP84aiPaL1T55jeDCdk5LTq0M3pqvo3Rg7cPh+EfdVDHfXJnm02LXHym
6SmMNwsRKOlI8SSxmjOWNcvoy1Xcd7Ht1re8K8kBSoDoU+og4bZmdni19kZT6kfL
ZNOsPqZjj8i3IDIOMu63ePe+JesIFxE+uE/udJgGYj/u64c/YDdJ7O68SGpEdRJV
e6J/o70u+50O16VtIAWCSuDkE/8KeoIVPeaO4ttcTc2Q3PlcjJZNEXTh6Myd1COS
kA8VezmxYUtYNyyI273vyWK70IzEa7vSXfbhlwJcuCEteGmnV/huTAE+IrLemWd+
yMs7HhZugQaxXdyGFz4CmBSf+/LIAQGWJVB5CYAJohFLkxz1CXMzJsIAQjaS0ITB
0RleWNXSdb8LC/xbI6fjtzK51HBEPtnqxFwJ8QDKaETcm1KSezdonz5syOoDAIoF
F2lIbDFmXBiwOdr1t2NR4LmzZm2V2GlKqdhne3VpAQrJ1iPBKswOyIoT/r7M0xwy
Bj3j6lxapV8rq4t1FYTMFBUJiLJj3vCQB1wm691NIoxouIpLZyH7lTH3esDyC3ai
OMDuBiMdaDs9ebkG3ULN6fsNKyrEKhx2oWEHsncan4G+EYh2vVnFlFUCrf7JrkBr
WWyaYTzzRz+iL+0/4mGbTfVPtWP+HvUdj2vCRz1BO8dbYC5z3fOC60ARXK1gOzRl
YVfKCEkcLASLErp45Pj5qaxx40G6yekKWCcEj+lMZFjX2Wkc3Te33bLJBsKbyejl
S7eZSq2Ktj5AcPguZ2mXSgqHt/z4hDMgMg5TScea0LrNy4OUi7Lg+HdMZ5rJuVJV
dTL3R/TP/kkKyZNiKhpvRViBwwVtHUezf9OnGTLXZDYNmyzDp1Kc5PTJvbOT9dPM
fxTipPm8tHAC0lsgpnXQ4eH9DjkO0yRdzOysy29R9PUVKS7JzsLRODczWsMfw2rE
zNiRYtmhsCIEpki3DDeYE98eG2/8fX60FVD+JQVPg3pL0uXGk5Vi4UH5bv0V4wxe
OljmfU/sdh2OnnQMeT4C0KM74TgDQvzwHB146sKwun8DHX6Ka9yNRn9bnP+GMnBg
FRjTi5ZF015OiDwcaiHJj2/sV0JRZ31gIr2rdxNWlgnxl+Gbf3g24VxRtsQbXLIV
IxWKGcn64RKd/fLhIR1wpEzEPtOfH6QAFT4Saafq8uWhwBO7mQuatFUaCIz6KVif
uVlhKrWF5XEEPj04pNMBwxzEb+g3vEeb+6t94S2h/g2KbcLoL8FdcclQB1bDbRgh
ObIplpMVYuDccFwisQ7f2quIhwfcNAW6Pf6KiGTxfj3dKv9I8nKBj4wj64vdLBsx
ds3XXauq2lnMvUqqJzma5K1p+x0vQdtAguTA8x0QLtq1a5XGhOtSGlFjieqFnfze
LJd2D0qTd+k568WNKaNHWOI1w71WiBsOICeK0HH/yeAKgwl+hW6XDupiyN4uhxAA
zxm6sMTNln65xyek5HqPhKzSjUspPrq/uIZhMCXyU05Ko/atEvzKMbGbVzdz4rgX
3eHSz+wziV24jAIY2PDero+5a/d3Y/y5r1fZTnts2drnIPvayhq/q0bCOUz/9LDm
oRRBx3QZrwOOa408oXzanoc4LX2TLAAayjVpfug93NCLViiUr3pshy10gYNmf5W6
wU6ntqTcFNTg2sFn+Sbx5JGHjyk7WxxgfL+GYF5YBYmXW58hMhhxQ48xT45KOjnh
UW7yjQfoUiwev/ggDNzxb/xqRmtpXg7EOYr8JkF1bp09QWg1j8NTS+KF92zBFvmY
Budsh3mcEzHuO5giQ/wbcUwTxMwa66qxn49S1f59pHcmDHOwJBrH9xQrgPoNQ/bW
1E6e2yXSLs1aUGq7NwPijx7HWKcR8BF0NOs6tECsrt0tLr6dfZRzuirWleff4plw
im2tw/31av/72PK6Fv7yuzRjvM5jekJNEqcPreGQjUG7wDeQyvQKw7n14FQnsYVN
8jpDzHFEzvpTH0hoILeGorj5ty/1iVVj4fX0B725U6bjNroPkVTrBu2y+Hi8SCd+
ys1qNZGnUCegKVS/VwxgKO+Ct56iF1cKt6QU1G1SZGXkVKcaK4QXrzlJ3JskEVAd
AzhkodSSSO4FlAuGbJU0eUMQwy+Gq50QL1dx08ISmCGCjNLeZyIaIhg5i6p/mVsK
1aRezUGv4ezHpEsvpH3hmNXKzoE/RFBNb81UsynfxSGaL/i2ZsxEthlrSMi1B+FG
67fJsodoN9V8m9PzMdaidkyWZ5aRNrZ/sAuxIzyIez+g33tghzvT9/EB8IA9X2F3
X7lQQvA2wVGqDD9Q6tW3deGjOzVfYJSzUn44GjcSod4oJMbn+7Kj1JebZDCt3oEe
HKKOBQaxomlul1NmlZf7eLYAxBZ0HFSux7LVUVOX6IHysXSGQEZ7UxBuZidtXBfc
bm/9QzmeabgEiPqYWc2BswPCcnFDjgnS83kFq1cbHPmhlWixzX27X5P318AhFjAf
uWrLWrw7JHsr/BKm1GwmtIBJlfYxY6Xjk0iXdmin2ZywSeY0ZIVmm/bHxlcyCuF2
wvxK0z/tyb21HezRJQVmKEOW4AvF1u0ohM/6X0v8mWY1YN2jPTr5BTgjEZzmbRN7
xGR+FvlcwZt0n9FlX4bsZozu12dPNlTSosMFmNECLvNod7IELAZHA0wtppnnFLYm
HBAFUpvk9wVI2UVqxfoj2cLeIPlN1HsJK7BVJGf4PBwKn4dG/+O4gio99SAv5nvk
AcLHKU3t0+xIQGzYwHAijxohsZwmd0HLhBfWW+UE20OxaY8FPLZEyba88xJCzmN9
apzL+wIWFVfQipOtxeIOGImGbzTSYE6+KRAXlU0E9f1EpqaTxkV/jKMA3zMilR9G
AZlefBo0fyuazMwhz1ZAKNxRXQeFrhZ2roKs6gGD4Ex1VObKwLTDJi+1CPqLQObh
2B+dWn7O8iRRe6Yb4DnBM+wwlb0OWcbmFbirx5tgfpsq1rQYNfDbdDLB1KeHxdhB
GMB+oDwFPGFv5krbsLbuRBmer1iZyPxjq2dNKX5pEcyMRpSQyvzqdYYiHmvoJJqO
aXkJRvqRATRFWVC0F87xv7vqJQObFuV/qSaoSKoJ7QL34zBTkg9YnGXBIGG/sy4z
b/QNdv7D9dYeQMPeOYrcF59+GFujmas03y+dDZOYDeq3ezF/QlzhX9twgVZQXyg0
9Xz3EbUV7Yo1fKeWDXz9F4lN3UdGsNJnAicsB0Tkp3mrVA6SGJkH7ZKhciS9KASg
JIOD6kwwzM6jGvq/fERN3HHN/Y+0nCVguMP9MAoK0aCVJyKrAg1KjlH4bQJgp+1X
U012MqgdL+2AzfiQixYZTdjsdSRaNECd78LtJF68KEqW0RZktDqacR2jdtfxCPVw
m1Py6VBNKXm3qIQVdNFe1k3BPV+YkmwM6La7Jo98pEHu6gkzmyFSQuHajhJmu1vd
GHOiKtT++U/pj3fBQe5s4EJD7F3fCkdFGXuzzsVqW8nWZTUBExJLQANtojqKbmLd
/mumHALKxx0MFI4jnUeuGp1bSq5Wb93pcqaGMX4w1l5lCq6VgwJaF9DQCBNo+YCW
36+tYwEUHluoJvxU8bUhKQ5JiPTsvLM79KsDlLO9cR4pMglr8S+GEkXsAFtB4IcU
G5IU46OP1Lo0e6xVySrYk87KudqEBn7Bp/ByldtS9ptdwAjO/78RI3m+SlFJM1Qb
CsH2Ks2er6FV9ApRT37gMu+vpg5eQsO0U9YNl1zezt65IZmbZj+m3BhQcF7vjb6V
7shnlEBFceTOqP91AIBJJt2Jkc4uVLLvHUghuHdS6GcN0hxkaedSsfNJhVgjZVFU
a8HtX1snJay6zn/zejh14DdCaSIvCjO8sl7i/rq4lOa1ntFP8xhgLKLai0/sjGM0
uThAZEde2pWxZQOjKJ76mmU/R5/wWjclCRPSvHLFsbimkRaAVrWX/Lp8kpsygwn8
7x1BukPr+hmlkmVILMVfkwBq8s1EaZrehVDlYZ0cuxAs9GeIFzxRozrc2BG/IN7K
VTtxhDy7teq4fr3alJdCts/noYRNQvqLvAORhve2yRCs4J7VipOVaqgQQ/eppc2n
vf2rPzyHpjNYzlnuU8OqE+vI5UwxySo9OMwVne5bKu7ntLr2OhqtNzAjzbOai8oG
o5L851Fcy+mmDvk40+cCdRPjGhtaK4fTUEuDuwus5UCZBVhzYqctEpIFogQYh8+4
sVyD/hgPdx67mJLYK/o8u13ypp7EHwnE+gnoWBQJD+5+27SSekAdH08/UJwI8I01
gGstn2M0GSU3t2ItL/Ir6nORhHp2CtfLbOQq4abGJUu842fxH/Scv7VSyHLAumX/
zSAtiPFSDXujJZa7OJarHF5W4eQBxXd2hnjkcPpaf77pGH4lwH2QjBEzFJvOJRP4
UFpYbPXVMTtllhTs+1bEzg6KL052pA2fShVpPbiWwKnpK5ptCYRFH7GiQhgYD18n
fxIAeFHcugc6Pflzl0tyT2S59QVNcKpmzT8XdsbPcFHv4a03Im0DemRSm4qEDgbg
jGZ3W6WOwIgeXH7B0qQo9WdXs7P751zUQ7lL2Fn4HMtEjdMqaHYiWDT07TL5rlY8
9nRPmObtUx3MCY2Nl0Mq0B2QH1zTLOOacO8Tid2QvkAJ0jQtRSotFrqi9aHKfLdB
UteYYksYwL77J2QlrhGuddumeg5yA+NZEyJbD69j3pr8HnmFMiGlmQxTdEJcn4RZ
qKV2xx5B4tjIut+E51C3PzYVJn8kmkYNlmvN/g91uCq8/E0odWioxRNlpVjr0DMd
viH+ubXT4otm8oqXHvkrhDj6UW3ueaxGX/f61dkpnMSdoh1YzkBOrlgpnrLNIBt5
v8g098RQbZCjOwfzhsNix/y5KZbrkxF8sru7OLIDWFtN8+q/c/FxYvOtRIlbZl1f
nm8I2FhVMp32gdL8OJgLgSe1OLjzXihKI06wDs72D8QQf1NZK7798qvy478UlVN2
aCStSs2Z+BkR4tDw6+7LNjk5EuP5HX5tRMyRtpNlqRYU7rI7bDfM7Pep/plvSMEP
S27WiWbHqdZ0t40zwnBilAX1K/tqnqIxoCRCoWLezw2B77bRELx23nqb17JS9kkx
DG24IlDjeGoclwnp3Vs3tBreGzFzNETKkU9800/t34k6K3tiiZgbWv/LkuZiyq/g
fypsIrlZ7VMQbwoQeSuhZTrMNtGBsPfugmKrQQXmCC14fykYZzClk10OckGsZ05D
llai/8O6NoukZz6B900YUt2A//4zBX3CofasDjpYnWmITdhZ2vbmgjrcf59xFl8E
2Y4cjJO+JEwy/90skT4Le0/RC7EBMJKhdO64n/57ptUXV2Spm1Pw4UcXn2bp26Ht
Xis92A/Tm6OvuAKKildQ4kKlqY1bzqXqAWaO1SRyLyeCJVVSFxIy/GX040hqnpih
5et3xvKzKbmXAU/NBicKPYjouSlT3H3VKa2xR3gUsbvp+9LP97Y2VvKy77TaAyD2
FL/XLu37v5rZJBB9HPItZ9WjBV2ZXbINgVuGejP0OYv7bKwAbS2EDw6f+zLNMdiZ
iXfqGx1vo4z+DLsvBa2irHAcWbRXNNzWF+ghZCFsEJTNRUVuNd4ZQ5LwJKnABU6u
OUb1da8Efl7PPvrRfTbKhj7//5OudfAbh3RXCqmR7ueOxBzFOTbPhtQgT8EYIh/p
bGZwd00flKVgqQ+kLdWEMW3goijunFK6TDdPLWOCWKWIMy9MOz/wjEFY8PqdMeH7
IdIud17VYRFBcUv60jeUrQUX555AeYAUvfXKnl07Km6hNib3uxqApR6B8zVZJUo+
6DYsXQj+zW8fh6+oGO+Co3PKp9w3BPIQ/XxwLpGH2wAXxlfzs42YFZ56puuAQqh3
8bpP336u0F72qSfjpUeDEBw4CeWRm2HwSx4saH3PlR4I9f7WntZBDzIHLV/0T37o
z7C2bBw6ERw/k1M3U+mIpitpHq0CUeAs1iSFkQ5imiuXlKNH49CERryEe4YAfpnZ
FrlW6UoRZw+89GB3bmrJRODQg1HaPS6JHw9ROvYGOx2sD5n0CcBR/47P98YsjYB8
FsbrMoBe7DvRslDQSSknaMEnuTOSv3GsAoxQdCSC3E1D4ze97D7mHUhkLRQ6N70m
Y02KnkTI4wfaoF2dkspnRsozCukBY8M+G7maMtlMKsNxoNY1zkhUrTDfSM3scGwp
nojNB6pbLDlDhRF9Sjtv+lwk/1h4AGHX5OQVBM9b1BktkuTyKkTnMiPppsG1QbwT
GiZDjsL/hZW3m8DkBSB+1U5zrlTLVo7ay+V+SjvuCzB2IxGkALDhbP04t+NTYmBl
v9J4xx+/MBEY44/rSdpasHMYVNi1UsaL9AyobccG3azn/A1BexTzwsHUop0v1ome
ijP5MkfQ0S5zxi6MmcoFTx+3Y4/OUcBf7liof7e198+9U4FETnVRpaoLCdI5WIMF
kyny+FKicSpKcFCQ92TDDZiHLFLyE0+c9Q9ULb+m5ApdFbIqOBOTS6zJcvu94IPg
Ya5dCnbe/MH7X6tlcpTF3211OoYtipx4WMbYeaHSh90cdGuuONL1U0aFyFCsLEx/
Aqq9LFbiESUFGy9A/6hhwNh7TJ65K8GcoGg04jxetA4Nl7zTrkxeezWrg4GEXDzD
TuULVVrVhS3K0kbvDrdDy3QA5t9lrc50YODMvq6fZhws71Qww0GRNdPIfZbFdVu6
N7B+dzzj/Fo5YVGX0sReVV0w7m2yY5X/Nr+hdSZRSJHe15Np5zA7VO2uI1dRdZ29
NoHHM2kV2TP4rQ6cpaz4arRm2E2m8u5HNE0u/gilQr6jiNweGkytcyVjmrajCaN+
CnVxRCMWWBmu413Z4WHAS4cQAGzyq7BsUM8V0b4A+HMOyxChEVRJCSehYQbAw0dW
5ZR0EI1WF69fkI71x09h+PHdbt8RkWxBHNmw7t93Bq3ZwMfnQqy4I+kTaMqIco4Y
U6DvPFdtXnoU8O0UBwG7uve6u0RyasbhVhqtgkRuUEjuOlYykqcy1r67rvlqImqZ
DZAsYbvqLiyAK5OLOWIW95iIHd4YQzY7HaryyS9TLWpGn2KDUXqhxA+S1Yq7+e/+
0nZNFBOled3Tce6CSEqHuX4lLyGomidh8ELVeltz3egUzF6k6Be6A48haEoBtluz
zHYMV9SDSRG8F6JtNb5P4wocix99S6qFm+C92cw7wiVLOXb3piR4Oi+M9cehT6BD
J4/0QV3tz7wHVOeG0JHjWassG3yCBTaMyEFr5YgeHSQvIik5w4unPICCx9twcayn
FwNSPFhsPEPuep27kGpH2bBByznlem60OyxTf8Fp+bAIvwf5X5iGY0bYkwB+b/zX
JeW9GDzNVMOTsmEgSkOFUBG+Si/UgW9BH31HzXaE4W1YynivmulaANbCnPDp8pwC
Udlhg39qh0Cds//sNNgxPjJik4hu9RVqDnCj1mGPD3Ug/tPfPSy4ChI6c8cVecea
+UB0QU/zgue/1IAebGaUzGqd8EajVblRSqzclLmj85yhWleCqfO81oJ/WuUBir37
6wIXbwbH6eY9luAglLCM6N7KpNFJluXc2DkZhFpBLmmjcstIel20obojvzimUrh9
rZjLZdeccnVCCabkPucoL9Uk5SCYRpdC30a6Jo4W+eEF+aChWcYMgTAG2fUhmkpg
zBan/Pkw848GHjQ4DYhK7qxXE3K2IYIIKD+1BJlJEjlNYD/S6Aim0Xh8zU4HHF6Y
ldmR6H6l5Q+5VSvP8UziOvfQRMUPLd8r4jpmnhiKow4FP7BFDvECBIe264iWauJp
8MTkcMX048+1OJSHFkU1L30cnps21wr+ziQY9lcy7rYx/gKPweHnJ8WadFLfQK6D
jEM3kN/9lI+ChPdLns7HNTVMP7oJuVJColY9dajznzlFawRL5mxdk3n3dNq84XPT
RqyfTwhy+3cK4vfQHxMFj/jNEKxEbglWHZsFlBjhKZp8l4rbskRvkTTpHhSuLEd0
AZsT1N/BsU6hwLH+TA9ycaAflX45mvjhDm29GYIQICK00HCYG1mn+D0MJ95I48Z8
wAm3vhCnQnpBJ16Oz2jKDX9wiyvYM4lpjnD2uqRkf5c+huTzm+FPjDGSKz4B6SQS
vGejzWlCHHwB+a35Jn+sIpbPt7HhiHtUURh6nUlY9EQb4sdUsWoCzB19sQRrlQwO
0gzl2DEDdPs36rVALHO1OBj87yvzCuAAg66t/KKApliWOB+l0XTAzPHuvScr6PVb
ozkMx/KV2RRuD+CPJ9pNKbXQMB/jDnK0fb3N+PCwuby1x1XBgC5YCDIGq9qUBPh8
phvoDRdPjLMZSBHxW1t0CBdlpgd7EoIXSi3gCoSdetxxVpVQq9spn4cQI1OX+t2z
yORtIcdvGH0IZNTVaZsehe78dVTPRyFAEetuVXO+AgT3j401GEHfiq5ws4hvmsTP
vXPCYjYCMUc87Yi37Bh2T8+z74y/PYp3nSq0P3QmxHET7IZL5fYCUZ5k2gpzQ7iM
q6ArDSSkx81tZt3E+CjKCA1qxR6Y/PD0kpcAAPLfIwoejc7eVR8oMpQzKH6eVwwH
2/977Z8xSVNVnfiyejJqCxkelLX4dfIOVdiCWU79QjD/FUiDppMzTVjrIoi7p9zn
+8xLFHvED9xhwPsrJbdl2eqxHl3QQp2j8Wrz5xhXky8ErRLT8EyPazomrN1QdcuT
gN51ydIm7/53SFk3rUSG3Z0JoYdxi5RUGbjOhiiomU6ZvvJLg323/RDgYEIFee46
SoTiGi4mXZNTJ4UXJsiC3JDbQ5S929m827fROvw/rj5xv1GP19DeMnbNzDs8T+HN
GIsak/FPLFa1uUKcD5alF2vVyGLqP1nY6L6AGnhzWqiCX4jltHsIfU+EHOzcFImV
cuv8dOCcFXepMo9PvEooN/FsEad8zBfKqKoV9XxB5ypFG5yP0zAkmT6rmuXRu/vo
TDY3IX3/iBJKrbxx/HN1GQGlvy73c0IJ/w6FuYq7BdI+EaJ+Z7YRVnq45RNPmcbq
eSbfLUGZpqB3o7GC7p6FOLVgu0PQE6DVXUvuwotr2InPe4OEEDZ0yboDD/e7EMzm
dEnc68TJMm/TAMe4Gj7qje1JJAYL/7F+qtgLBrndxsJkMViggrcISMGiiDFodtSA
2YcEFmT3tEhxpX+FljKfSeRmQA60hbHWyK5mgOsK3lQazm6QbC8PFhwyQUZ7cweR
k5/PosRv98/+971J8nSWVE9v1gWmKCmXXBaw8Qji9HANoLnX6r8l6pRo6ZLqj27i
1TjDzgGxS3fC8vrbBtBoo2194foOimQVwiB4dffNwR4r1YeipHTY1yewWcoVO19M
PnzIDxaSsW24WnxsKtyHC+YYSEWY8rgrJPHku95/fdHo8qnjT5MuQzBpc35dEVYv
UPKYfi9H6E9RBXovSTpXHsZZaUOjUfhmbbdsh3oajqtgSRNPPq7CDC2h5g3LKYU+
40yZablKEWbl2HmvvLO1boLj0VvRf8FlRbsrFvxnwaXQzwzggixMS8FmSE5nycZo
u5/eIB0ntt1VVLFAgJ4tUg==
`pragma protect end_protected
