// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DRbNONrHHwMnb9QbXX1ZEU8t4m6+kK/4STfIzkroWdMsDBzMCY33l5rF5ER3ujDJ
3lV3dgycvSG0O9G4bnGiJLL8ihB5GPvM6PeQcQCzP8x1U5KQTBXF819Ux5Tsh56u
Gfk69QSyGL81MCC6+iOBywaSNmBDUBsETI8TChnYlew=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21168)
LPo7RRNePPMdsdYQK3ocUJHEJvhnrd/t6a+NBSZfjNZdXmWlYaVv21UmazAuCnZ0
8X9f++J6sm7Oc0d8eT270DqCQqq/R7j1he/e2ZGcRP36rkFpvWQvfS4MtdEgRFCB
ogncvtZD3RQXA4jI7ZwFoLRip9zBNcxXKdmnwETLrDRLIn5d0QSqrbm+6eqN8tfD
eNma/evIOWapPDYF4/1+QhGOgZV5sSfuDLROlvaEkgqYEtHkh3ypL99U/HWJ8y3B
xsHl3ozhbhLuw41je36zKtF/obtJ+FGc2Eb5IXiRoAmJXTMmSX7dqDzv+KF/FMWu
81q9vWgLBvW/h0zRfEfaOAx37/J6vl9c4fE3kHs7VP//IMffpK9o3hfHJXrtSBSD
oMzsrmrdTMJ9PiU4BrnOUv1a2I1W45wp+pcY+HLFFT7Jz6F+cdTV+3LIqeQnw+Zu
z93lYlpNjqUsl6EswUTWD4rJHxTkSNZcS1o3+AiWYm2dKx9PyovgeGRHwk+o3Ink
qJwBW8zlhFIUnDTyI5ZSgMTvN8m3xCg6N5UNXpOFK20MLKYdzYf3ky+cCMEjmW0u
No6ze6AjvBrCB997LhpvRZ+Z3aGVGIWhVdvHWCvEyThvNVfQMWoQ9U5cWxcHWAW7
CfqfG5S88Z2VTvT/OolauiPZQ9gYtH9LYVvhhN+eI9Mu7iGDRNf7C1O7BsBY1CAr
jThq9PcPY1VfjX3NIyoxUzs+hOmM7psWgjT4Y1mLCqFLaCdQEzVaDm5UFiU1aaab
RCvnDdXOOA8bjuuJbL5z99MqCJhUWL0rbOJKmMtoOvYROVrD392BVYFHjVzwLDMo
e4Zh140WHhE/HlsONv4U/R8iA/52fockDimwQql7Y8ia2DQjKCp3J9fjxKA+92N0
lFnQ2saWD8GGFiAaeeP27Y35nfowXYKFgad8HuD4JHd7DdKP+wBIQ0d3BgrnHfIQ
5oiic6SQIBBs4rV2mpe+BVgUczTChC3XosSr9FoJZdaj2UIoAgzBhV114s+nwGvr
7RhGkCWOvCLrDM04xa1cndbqYYFchWxyD7l5jUnmg1+x8KIJYbOt8Q0gh845oXx3
Yh5LpujqANQ/rxF2GE2+mP/cbS/R41GIPwmU1yvdKRCfT3vgypNZKHO5SB+QNcm4
1Cm0I22cZogv45z9qBQ60NA7TFn94cogyXGmkJonUDqzDAoG2I5mXoFQ8C00lD2v
VnjejyoFPiqCJb70bfaurrLCwn3uR7sFQ2Y/ERsr6OF9EmgUhGUKwouJHLCE2O5V
TTV1/0J8INl99ozG3BzYeU1/1+ggnfLh0lB8m5HS5FG7OPY+1x+QQVQKWjC3uAKe
GJYYN290hF5yTqOC3o4HIUpG1ngxik320sbYhGZNb+Xj/4hZqnMeuipMSqIbARgZ
ZgMI8lAp9LeOhK1JZnOUAmlJBBbGb/0KIVFKwx8UOCB6oAkwSxuSUzP05ckKg8rL
u66dLo2RJeUWT6wNDHIqTLqFMyHKtpwK/QRdX6CmkbWyMeF2SQLxZw9pqZ2BDkCC
8/E2El8MHFrJvx8NCbTyQqpeCRuCuvGgB6NfWtdvoVTxoQgopl2S/FGwAudoV0hE
e5uc963te4YBLmgdN0kaUpBWtpJ4LnQylgDqbtvMv9gAIMlytFG904IJgQNdq1XE
2Trc/FFn/SjO+g0ycYsY/hxetnp5vdp2Ak/UrfBlERCkHC+5LnoRw0b9oOsGhTo0
r1BPK9+Uz/h1SffojwvRxW8ZYKg4lRd5MortqU1y4eqXPQUIZ36g7Zvz7ZpErTmE
7GYcQbn/ipbMni7/7hro4BTR+fsjhXkjHjqdo/AkJTtvR6jGTc67M1EXsJzKSb77
YCG/HAqzIZAyFyI8BFHZAxdXb9bjHbfTFoPNzHEXAHJ4U0mRxxGkiU7rKqSqlXSB
WFQMc6qZ9qfgStfTY0AKAp7M3I3r4eNQWq1yPEwX0H+UrJKF8/YraLQy3cprU7eP
4yInB8U4XykJaWzMGWVAJy9P6m8ilSoh+T05buxXT9LrZB9OZsq67m4Q8OPU12PY
FJ14e6M/Jp+4zSWjPkQemhChJI9hFHT6h/RaszXzIHtkAT27TFo9o2XGzP+jCQHT
bXNPZSZJ9xUrfp7aqts1amhDhekhpU721ODgp+0K4DOq2HvaQv74jxGymrv3itUi
Pzai5G0XT3WFPB0tbBNDXV+SlFZ91ge8aWq/in4fySxxgiVOPIgtQKFuKqwYlphB
xRtFMJ1d5VzNHVdopuQKO9k8d5SiPm5n8ZoMcJQeeLvrneycXwyJ8WI08QRntHkk
PfKPvxrv+pl5MxqGV8EKyJOcqqcEJ9Mfh4FvHucPC5KKcPVErB7sOPZRyVcIYnOg
w0RcztEyr1O0YBWueIpOLHhZjZ45GoPesSKec8inLGu9uzlLdQjc3WVMHr0ar3gn
JLyYG6hrJvtOrzbRFJW61v3fVH8AGdGgzlBdbqWEOJO8dENVvlSpi0BcTJsj+l0k
r3yHnpVyp3xLAJQ79jzFqVDObYHjHCDT9XCPXw2zSzX6zBzkEs0RqHZ9TCamRouf
remADuAG+XYZoMh1vB5+OplU4jwT3dGPZ/WLW2mYyet1oI+AbdOhvDnIgmqHfomW
PUO/oISZMs7eLKoqKo8815plVuqYFAMGMRFHqk1bLAKabnmijYHATisj3nDAfp2D
qsFtPoFlVd03nRG5qAilzYRqC3pvADxGnOPlADtZkKTcxN0hjRSAgmf1ha79muWB
yjhGtikQ9al8OgqvTlIcJgjYSbiESOalOTZUEbP4CKl/bWdBas3qiDW+hHuYVS2V
k2dghHxsV+/RfcQPeiDmckeVeeOkIz7rTkEgXjX2ERRj104OdtmYE7zTZhfn/5Wi
XjXoac0ApitSDzaUgtkEuLIkCfLGcP8wHAu75kbl3RrBtvNQfA2zwwohJyWYoGLx
6ro94UHMXQQOQFLLi0MCDpuH2goo8lV+k+RTq8Oott2cHTdHYW7u//NgQ1GHYMr6
FWF/7wQO6n4daB6fXTvaUyYkJnG3QxtWggkSj9mQWcHRlp1KjzTRTJmnv9JNHZWX
nWSNMGrBl7WW/9JWfqPaTG+Ox2kAmBsuWilDNZl1rxXsV7aC912pyihIMaOg3r+L
sQQ25Y2rhIdodvkPKiC7hGsAgszYi6N36iKm/9RF/917k/WHbAEJYXLO21Wf/Od0
ClLj7Xrywk3MeNHKLC952uU+hmAmrR10j7fToRzRNF3qeF3p9t03/v4kPiHmOvCg
hpabjOZPD6sshE1pm3PxrdRT3mzBC28wcbNtJNhN8n2dyABboulIYICQbq/aL0LK
mzmh+OcBUEvWvvddMPdoIMuwIFXj1JFwjJlC2Cg6jBK202/ysdlHZtYkK+zTYqGf
1D8u9hQPksrkOhQRN57E9Empc/SNDwC6kNyWeDcj0A+eouNbC5AZ/q1MO9tAMnKA
8Pu856plzvPsX2CIWvjJTe+14Js1RDY0NQUB4GbUn6CgF0GKGSh5+P8cUrrwy1oM
JZWw1rSXw6RnMSVioTKM+F9JvBQTf3WcMBa1K17JoVDMAs8qxxuoCV9u8HSxOV4S
vjPCzFLFofVcA1xLMeraJQlw9iNQdyhAjV2OHpLB939dJo1+lMuxyR0ou87266BC
GAsXsUab68DVzLHgTpp0ZYoCQj6/aqgib74WLGaNB8AdN9ptQyhKz0mtKebq0ALR
dFsnJ/7G1/V7E0UPxV3SKSXVBruxOrF4yYq/8ajeH/uz7z5UsIKMCXVH+zi5f/87
gMvnlTR2VeXqDhVsSTE5YlUsoLm9KJP1ts+2u1ppT0kYbFh+ao6H+HKqPVEXlmgu
1Hrko0mHjCkjyBGrN7QHOZrhWpF8U41atGzbmk7hQD5tdeQ7q27ys4syxE7J7LJa
cD5Y+QPzO5g8t0DWinnvCVReQFIA/RhbW7n9Mgxy2lDjyD3PA1nfccJJBTp6zCNt
0DMq52nkS3FtNt625zDwi1TJFCqtvOmnEAGzJFIQmBwV0Jt/qaJ4kPLr0+YfTnkd
RrqPuVzh0HzmUG6+rW5oqNVnIAUNnaOfkiAW2vhnQdgAto1jSzLiTbyGemWbC7NN
kbb31X8FPJPm2HopkHcppmlj24n+rpePbxMhvpvvgPEIU4tPoAdW77HomIzxQ8II
j4Uq+M2RvqAzULVurvejkkj88Ct8Z64l0RvDM/u+sz+qnqR+iPF/Hk1MClzxDdIx
98OFWyIXGvPTJ7oUYjgwQHFKEKjRWpLwelLCdkPxvjqslSZsvwRs1F3TQ5dDAX8H
DnAq9rvFyIIy6WDgCQJJ89h1x2tKc71w8D3IRIiHF8YhVFavJf+/mR/5q1RgZ/sL
N5xnBWx2cJ0QNjTIzhaTKw00NzKk9Zh4Id2l4379K0KtRLd8/MyaNrCo+iW8hKWs
YI9AkUMK6wprrFdKbhe72eLX4ohyLJq+/NPdT98+aAzqTO8QokQBLzLHWcUI/5R7
K0M7tsDf5rfZ0Hn+EPbSGzy8jFX6Yb7qxXE4mp1if0Y98xK+zZUG6uTuLWpgmWii
Zj0rxlhO3XU5uJGjlwWY+d75Rqy9Pi48z3l7VfO+3MEfE5xuh3d7lHKgsg9irrzr
/EpzqBXVOy63zaw+HdGjkmnNr+sRXJEDf38hk/h6KsxYM00SyY/c69oK/+YVuqjE
gDBDicbRy3B0xIbXuwPKM9kEdZCCQwUKoUrIl/nmJ0ccjDoQGnJ3P7mUzlYzwOKq
JzxwOSwnZBH18imKIYPsrAbyJwQvV0mFNyR84NM0HblVA0Mc7wYo2WXZLDz6sbYI
Ev58Qx9niDyoJoaRatYuQgEbjkwWq2XOXSUyKZSBasjuk2sVSvd9cYbJRLCq/UPa
r/tOOMVUH0qnfbcDXBLOw/fJFuubHgTmaYOzDqqCu4damodWaM6GRae++g+W0P81
0RUzq34IGDXM/xU2eggSb5RkvqkUc04CSCz7xDDdUqnr/w/wVpdHuYHh+j1fOQcl
ewYjEipOjkkd77s+czcjQ9QBXqRdKNzKXURamCl+WhZq+XJpI4bU30XCTaXuThtA
5frVJnVne/OFHnbyd9oM+ZsUv/1qZtEbKhdouZ4FtBTEqpttJSl5yVakCKu7GH+m
o24ZGVPngIWeMd+vCBEHvBtTxJyhcIzDv4bdY8ri30cK9/tK40pubiVBTu/lB9hp
G3wRdHe+iu1IRW9XcyyBVG/3w0mhkn/S2cFiDDZvz/0uBtGBzNNo+uMa4YdEH2UO
5O6fMNnZCr14mfeU509tuivb1XANMrVhKTbjmDyJrYID9vUHmUIWY39dfVj2ge4R
eFD0hpy6dMj2iOsAY+ywWf3OUMVEG3uxz6TryZeQ6sShb5k8B3koc4n0qy3SiR8c
owqTl1+HGW62sdB1Y72431A4jl0pRUBBizxgr2Cmv0neLXMS6EWNAP2Yec//w2sq
qv1RY3JMZc7zBpdiN8GCttzE+aqcGri+eJ6iy2flISdoVMyOuNEyeX7zQoiYs1ZY
CEwXv8XXbtL0+ddkxFawOZmls9pJ/3GVWo1lXFEM82MUDbojUYu53+jY3pd61Ali
dcPjFbbTC+QL/520JL1kX1+u61opfPnctUZMncelxUyyPd1sjXWWGZTLveRZInbk
CL8nnxSXtbIFQ2dhFzwjmYxrIgvZSohouI1TPbimHIIP7zJdUGKs77cbZB+qw4FF
bgLZ6qYfPQDVPWjIBROvlUdMmDsvMawbvHb/QBYhDwd2kfjBLap9iRGzXkQRTOYO
H3Vg2HwTik2MFwx5hTWbhIciXLSdKxo5dPR54VjZ/G6defATbNagSe8wya01ktg2
HEwY1IECPEx22qfXuaF9AU/RIwBQYb/sk/uI6xl5OA4/isv8eJi70qhNvr37Cg0A
m9S87BtHZuDgOZLZNHSVdURZIkDSjhtK4afARRRLxS8JYiubchHAnJ5QoaeIJz0B
gWbLEeO2TYm6RDKMc7kCROJ0uIMIBjMKLc4045SOl1cNGHtmV6pfS41qwD59zEji
oNcMeBSbGUumtHgADn1Vx3wx5iC1JEz8Wr23PXzN8nF2g+CDPYxMi2WjECuwkbHG
wwhLDcjAgXWaS8J5imU0b/LbO6ax4hmKqti5t1XxFv4OSXLNKpqTWykGwENj+MsW
vgWUMq4BhMKGrthVHi94Jk3SQj262lMgRbRgXVDOUQZpzmuf2fO9i/jETupk0nxz
47gZXSDkwwGL3JS+CPhWdoCDCBkjir1EKA6TKU4rEQ5ZuCIsicXPUHEX+p1aRiHj
WfybOIO3ZTBXFuFkjQk6l1hd3bZy5HA2nrrnsJ+yA8pJVtJ9vv5bGu64eDSl+Xid
AHCD6yM1WW1DbyUkQuw0U8tdnzlac1X7/It7d+jR4GrlzbUAtpRsxVpPeJ/G7B4V
XRQxIbypYJjN2ONcUSMiV0MyKjpopdO3rR6LWXi6jqGjeP8sekWz4kFeaYwUt7GI
sUqHjwwnBdPQheHXlu19UVi3o3mJE0G5OqSShPAFOLh2PstOiWhNptSZzPG1UXV3
YX8o4NHYmqKBxtlYQiHjdBvx0cEii9//P2jgUPIUeToAbaLbbRUYeu63TRiMIZc1
AXdchIedASpEUr/qUvCJpX0xGzPr6NTXPUp53CH6GEvjHE6rkkdZPHLmZgK925tW
gmQ5f3mG5nQtg2fWIAG9cyK09iwwqeGGDn16MrIJdhMDskko6zPM/4RDv8P4wh4Q
LRGZ5TqjX4V0POWZbhK/f9DF0WTE3wHEiC3G9uD9LWNYukz9PdqCCriD3e8vdO5H
1Dzs0GkcEJCHyWPDmPyjN8xKezXL6h0YEfXk0Tz0topXbdYWrHVAMTAmxal3fYiZ
ktOOCtiJE8sZqCCIXsp65KTfJQSy0VnlJr9+qC8ZhXa7t/WOdcbzN0ktKfaFhoU9
Jn2I8to7iLeYH2QI7YkZVljyWvMKxIS/+kHmPdhJ8fpIPyyTw75zKQrb3CjI62oE
DE0q+4XHDyKTN2psTtp3y2LzBovxn8sqAMT0x7xTrfbQ0/iiRPANHs0+4pEHWJDz
R/fj102dp6XDs++kDArltU88Zgg7dejCZYhqZLWBBvUDHPsk7XRbQXK8KNiWTPNX
QrGzIgu/s5SFV45Lw5XirCXWjcbOJmSdiCZNbPoc/utreBeO5n0C3uTHUoSeqUfX
s7hgTi3KC+kFNxm8GKTGrAh8LsXzL6eX9fK3KhwCtm/oPKvDPe3tHRQeDtg6WNek
SW32zfb6HpeIEcOFRUKVlrJYeKLTvCsRoF5O11LyvM50WIo3KllnQLLS5I+fuy5f
ppzEiePzCIxUPJBBMZQaWrNWMe4yavvYBlx6gbj/vQo8KNOkg8x/Kw+SvrxHoDoF
qCLY/i8I+poyLMuuyKDs1yyCYOrJufB/F8hdVIWs+oUwQmDzc8DLhk7hPDtv9LOD
lvgtKxb790xqzUShLsmvkycBPOcfGxGnC/6ars3k19V1d7ob+H8iq87OJhWK2puc
rHt+Wy6XicII5BjUkE0ewLn/ubkMNe9w228fOInY/jGw4nkO7LsI8YqCic4IpsTZ
l8dEHUKqOJ0BJ8/CxBT1C9SI2odliITsqBrbHD9YexMAt7TKUj/GX4IJ4s+ipFYR
2m2UzgC5J79rJmGmiHRBerUpzkl+pAFHCG3RxED9kLcg5uLmqX3eUojTyjhs5eu9
nLsULP4dqMU0Madj5v+VEVNbLVJ3H3m/rrBxJwpEtTjRnDewU++G6zUpUfbFdCiw
N3PSZ7H4O1rV8D57/4pzJa4QAzhmSJtRPLWQ8BwhI+dQ9DE2K92mzY3UmQ1i9ELD
ZcommhK/zIrLGo7nsd/tZ98QNM7GATC13zDU61bAuKmVt8QZ9G5xbE7gioOr02zL
X0w8T9E2YjOgiMJHbm+3KisSDdmc7mp5l/d557Zh887KoezWe8bSodl7ZwIewGIc
mDwULs/3l0AP63P47rCD2lh6poHoLJVJDjwWL6/FJVD03nSZlvrv3sXr5t6utX71
Q6EYcum1ys7QLajJu0rRiq9mF53zVKS+F0ICfhnc+9K+2v79GHJhJnEFBAXSvtHT
lxRfA/AY1hVHkOrMy2fzPPGy/6XJH/Y68O2qcL7qLNe5AG6kmWeUxe0WG7GHfTXP
hnVLL0DM+mv90sZSob6BqQgr19Rpd87r0eFBl8r0cCq3D2FGBmLCdBXbzRcKGgd7
cgyln48FGNMGotSILa03VD8/OVomFTUuyEQuMCGx+RFlTaTzrG5Qjk/kmOpDpaGP
594UXzAheOM+yP/UI1T78/WpDMskapXVhdbHOlSDrpH2dg+d2MpHYQfZFZnk1UT3
pCIvbGGiQdrT9ygB7BqUZ7QyGpKzb0t3TR95gwVIAVeDHKZc94Rv120+UGnLvQ2P
klSlNMnxA7UAk1KUPW61VXQ3wJlUcNlwKnTrkoUPWtxxEZvSV1oXIFim8GztEs6b
lXh2gny1QL/RzLxM3CeJftaWQxbvu1VNGEZ0nPVbbbv/nS11cqUJ8qUHqUpm4BAs
A9Chgx5c03v7gKuRPEhW7LFugwvP1Lptp2sgX5NhNX0wioJ0gxw8KRGDvONh9vrT
bZFxikoEVfUMrkUHhMtYKrD3hF85f+Dr266itlJbo8ojc+wbYu8UU4PQOVvmUhgv
S6lDuYdxWqUMhhE/H86L8ENuIpV/zSv381X+Jsi5/VMvv1lg5D53OvARhDYwuURZ
sgiT/f2VqXFy7xlBPGjmDuKNh2i8gGMB+hmdis7nBS5YIXDrxf/EvkWn5kzBAziL
aZmjKdVgshvoJOzgeHpbUx4ok2u2rF7I++j16r3rvbWxSptzYuCGKfN+bb74ZXYx
rz35Qbz6zVB1cdfSs1yUCBmSwQL7NXTMyvcQmidkyIzT/QnJFFf5qYiLaMMsi0pP
wtswPYlcPof7o/KSPfaDEwtScstHBHT8is90o0WjhunprG8ym9bkWFLPhWnfNwe6
Cl48+8RkUxLfye1KtsgganSPGksISaQZH2jxruvGI/q9GeLRKsrjUfIxUn3qcPfr
fJwKiz+2X7fYJ+HUOLZWGPWSW1fo4+yszHo/vpmofqDseBTZuaK/LhwQLniuftSS
PJkMdqfAv5F+r4/8jb1Vy59K/4xy86YvKlsFDjA23EPfnotFE9yZZqZRKBaFGkNZ
LwpOy/Czoe+9j3ARuKYJvTvEpYwMj2WJjHhGFVGahlfR10uOCvCA9nTBSXWFPBcg
f8DnRfl/BmkGeXA3e4XpnvLvUkvykLMNoEw4u/RF8J9JfMKZz7EhtnxCyPuXPGeU
t9UI6ZFS5m8sWAVEye8DaJr7acaKLBlVZmziYG42J2SQNuHTgr1IrZxJpcKIKpH3
u4O6K1yzgr9CgYZ5VAQohWoTWda9JqLKGed96dipRW9SZKK1uFc+aGw5Cx4M/Wae
yPYksgjrMEkZ2fGp9B6ETNUs5pima6lofyelLeAM2KgHa/Q0M+Usrun5YX5ueuKL
+acYzcwr9szkDDyw+WBnFuMyC+Taq4I5xBvcQuthhQFzov9ahy2fkc04IeDZcERk
5+/Z4zdyT4httvfRYXr1kKbWOetK+Hf2AoTKxtU59MZljyZsA/A5xUfDb4X25qiB
WOi2R6Bg2qKzVBWF+RTBkd4K47lBTtdFt8wQf9hjBzbPqQahsRc6HWVJ7wBR/MdV
70AjpANn6744WORbnEQIItKgO+GaidQ1B0GNpghg4EJLLw6jcQnsIQHzNDlWRldV
LDmTiVpz49VbiX1gWFjHgF/NDc7ZLhQVZVSrAOEcqsJehfzZQZ1AmsxD4imt9rjW
xNkYTp8sgbdaCmE/rhHR5/pfKe3Rot70OJsomTn0jbMvbckkyf4rzFcALiwRQpBG
E4pv5cvc8yNyjilAsko0WQR2fwl3cb2KfYGMRz1HstdenBTSrJbOwwkB3jVk+uF1
7uH91oW38Fzv3OlSrE113FlDOIMeRjZnVxTSBMCSfE4L8IeQc+Ap9hdUUQECI6b9
/O5MARdiwRQ+dyaGKGMc/aruN+5GKiDccwj9AlHX2lA77Q7W4GSXH5vlz3mKO2O3
ywDfn4GbL6UgJbzLO7HPr4j3yQPxYDaRoyD8VDrUJJzeXjxxGE8+guAqlH1yFxAc
psO2wc4ml78DpdBk2Yq7qxxqJAI8/5eFNUv8YURHGsmHY7RrBbYi1a00EngQ5WfH
GIH5VQR+YjhI1OOWaK/3NyPsUoMPT61L8qBCYQ+Z6FKr2bywHdauthYgzBpaPhi1
W7DDBzAqpuSv31y4YyU0CCnhAvOVchg2hk4U1F+2q6n4+UWEw9QHD3pVFetcY6U0
kmlOPptQWp1lzHBGSX5PK5q7XVFbFOOIJTlE+ky0BiKOGvpVBXb2WWh82g4MO40s
OrRjvyCJs64MVblxVNr8ngcZdWqlNzogjIqNouebGqCFUStohlHczSYK4QM+4bfW
JDxn6o94MfVtnZdgtUua1A4LDwraecAZEJr7NjxhFdCpejkMbseKfZz16zNFQoB3
p5AlgnnflaC5Bn2LAlBQojY1/u+TdqEnqBSVOP3IahMnoDVt6y6AF0Z52OuIpPDm
18TIkkN+Ppg2AP46AAC490jXh13ZQYZWXn5M9M9ycPSpuyLfqqJyNRXeLZtMoy/C
s0jPob+TgibEbAwU5d4HMUDwpnK/0SOUMJ6UQPoxdwVImZKnoZUTKxyEiYoCoXOv
J4OgTVR6WD4yZ5AcorN485/m+DxopBmzQXiipKR7J9Ck9qyZ3VqVdlIQSp4s92Em
h6LWdIfePnEIlh1hVHDBs+HLOR3zVf9lyLJghwxikOyUZuZ5epwLqhJkGjgr9vcJ
ydvj2JoKKxVTwjGiQpfaAaxA2bK4a81u4dsN3S9Yu60L3mzDQ2uvjMV0VaPF+pG+
vRGBNqmoOPw4gUcWL9k8aaWw10q9pR/OJRuZ+2ydOorhwcuUWI2MU0Uc1QrPNPE+
x+xUeQjT2zeHzpN0BJcMw1eNCFPkkO7Uk9jlQFmkO3NcsWohYxw9+06dSW9tz4pC
0E4wb6JW6iF/b4ZyX7MVW2TZr6KTh+dJYyFhcOpZhSvTDp+m9F7OxqVh/erXFx2a
crxWDSfPdqDCF8nJOcys33rl3rRHtt/Kk2uFB6eMxNLQgCT4uOpEIo2uzzOx/yu5
bhwWZ5irBdtzbFf5r6BPBsX1In7LSpwBl5tyn3Mnwnh/gy10bZtj4y2Pe10vwjDL
UFS6zJuZWofcr30/MZFNvyvxkNqpu1whC2Ic+SrDRbg3OSAmURdpIAtvEfmtzcoy
5qPGGKjVfjqpfRKlP0zdLuTMp/MCmYwZeXjoLjERDAWLxemnwz+47fR7kh8ijtWX
CdEtilErdKvspX5dlCvzdZjKBWhGekzTmK3ZCFwcxJ66MNmakZ2RtXrQsuQryoEc
iH324KTzLddYAmCMYg6Mc7QaJQ97iNc3Z66+eyQKhjfOrDMLq2XbJL/c21pS3Uw+
inX2fSFru6XnTXiffb/mv2ziqom5zrqWauJ+mmvaesxm8V3l2QBSPQH+g4DkiuLT
H3z9TKCzhKBNQZVn+YSFpny8Q5n7fSxwsisUNBMSbJHfJ/jrDCnxcHhQFDFGfEHk
c5oLrA5PV04Hau+rR/07y8J0Qj+hOZFH/rms1wD8K3Ql5smU6Z39bOyHmRHADdbu
ugFnbAxuHuwYUawsiHiudVmjbhgNzrneuxF3TJHA5nHba4ui61FEur70CdvjEk5N
tmD4/4hxGPJ6TfA859cVYJlZdKZk79kSiQJ5Ph4h8eCiBCYl2p9w10c/ZCG5Lufs
+9+L7QhJU5qbbXZaCUh60JFxDa87nUaaI6oQUWX9kljD6V7TcikaJ/yHEDSwb1WJ
pQ/7lUYen/A2FH3TOLq6V/du3xrUHRFK9kxIeeOctyvu/El3NZDYElZxqPfGzyme
fW/7GIYelR9XPU7P9EcgjukP2fP0P4RhuHTL5KnzecEZyvbdX3kOyEQTAmjD2ZcY
+Gjb7H4TF8FVTlgJ92Qusk0gah8FYGFQQPWcy3p0AFdatwoQqCxyGwU09dvT18l6
9EbCBF1AMDg0VheWKpWRrzOVfDseek4iAyctN1lIWbFGysiD8He38wzC29zlbmFA
v5gL0EhPg55zJj+Vh7RMzyLGEvCkusXowx7LqfQ2kk4x6L9jeWZlacjxlarWX32q
Y117B2v0aU5ZynCUa/pVCq21r4ckfDzCeM+n28Sfb1mcLllTyB2UnaQkANlW4qvn
MeF4LL90bRYLdGZ+4B21EIhJmzEeJRgZUrKPrQ9JZPnjBIv+0p0INVqLu7tadp0v
S6pdGhIxYIeHl5JhHeNaGEVc/PuUBu2wuk6vCHIpjSTF04wi9pcmq98LY7nLtvil
yENy0dCLJ73A4BWPMxFJG7JS/mwDV8H09DOWEvJSwW2b9EQhD3WSpZCYuyRXFSwT
EadTGL+w/aB2k1eLYrKfTUVHKUmi2yWN9f6NL4g9ld4YZdi0JBpSWm6TftZYS6/J
RPzDekPNahzGUTdF3azxyAd6l4QRCwzol4jyQxoPE6LEXl+gxBMhqPH/6BZNTSPq
oJewYpLn5FXZ663hIHuUrhzJj6gNXsQjFURNHmhzedMLCydXNukM5wsYbCDwLWJq
QZz9XuA7BSutwHDH+5Fx0oq6VWM3xG4oKpc80PAWR6n3AFAnbNWhtM97bVorxGcc
9hlecl6HbPySTkNTZKIEM2cuWkcbMBC48WTaIARGTursU9F7UknkaFdPPNwo/ILz
GBFF2FpGASZsXCdes4HslC4k/rz+Q+zHeata5bfiiE9doATwARAuOgHBM1+qzKqX
kvOvYxmcH9DKAbu8+TswIfHcAbp21dW7W+rEz6/Fq96lq+kDT+DzGszq7x9+sb3m
ABw2LNc1n0A83mWf98chKYqN+vvUdIHXZsW1F1leTGzZrhFop5+5fNmzpvwMD1nV
tVERmNnkid2pDV25723pkXmy1b8opuBW+Pyrp57McXHvg30cnjalKYPlv0vFWVcb
jTNVfAPlYpmS8HVpIG/SJV06/GxRqbUJ+xZVveD5RSqmDm4b6leWEamUX3QL1OdX
hh27VFq0sxO4rDtPa8dkt7vEDbh3ieiaU4nkEBOkqfsT12lo1oI4d50xdSD2D09V
xwRcSWzjEV2Yh5hpaSGuwQ3WSkAkoT8BIJm+0kThFsnEIX7o7wPNzzrziEKCXkKY
tMcKTnAFdkChDXsIctZYAAbimn6F6gA9ADs7DEZY/x3GF5F2DMWMuzC0tW4EXsei
hRpn3HS8Jx/ITxIovLghyOpfIvCK0963J8GZ5wcx3RMRgdDbJRDb78l7SK9Fkqgq
cD9G6k4q8unMKmu62ybKA6GRnRdhp+mRKZ0U19PQymPEKYi185GpLJpJPC3sbXSo
1Dh1pGm/TgJELjlRctWpW3zKc+RnP4FmF16VgUUDpiaG4iDpHsz9DoUZJ5dQT9Y9
CW5E9HZlhqUB2NS2B+6Bz/f5BoLZDRxe6r+SOnEG+1uFhenHA9hQXrJ5GV32Jj93
7HW1h6PgXXkltnyCNnnevVslEyidnJ44kY3b/6fFeoXhr5LAhdNPPVr6j2sUlqkJ
2pBVgN/kL0AJdhzC6Cp5rEHTw+DRQeFp5ReS1sakZ9mUk0+guWID8jeNGkwHpoFK
11gTbv6CVsEtrzgUvWvCTn6YL2FBTE6+hBRA//GRBhlefidSD4DfBIMIdIhnwps3
cqB+rSohKeWYA0C+IYavES8XseAjkro7jR+6vVHp5DwRhiZbgFOzBZlsatiiepvt
hRUmYvnAUqV6NUB4OdevGTsPhf91rUpFxWWrFVRR7UfkMa0YA/UNDVaOUgbyLL8+
k2l9zGs9Fs8HMUiAFQi4olrMd0zQDKgBPXw7OFJ0UXInckBSmfupfqJ1BcSV3Ohf
49VyleDASwkLi1qDvzuUA4/psmxZcVkndau0bloeIG1WNQMetjB7iz964SwJkSXB
2Joyi2Z1KrTyiKWKk9Yvk7ucctekPMQBNYU2ySv5rJfIX1Y0j0tymVTC2WkyeZl1
4NGDsiJfzrvW+g2xpS08Uo63DM2cQOmLjjSc2H5WECvnPCXgd6PDx0+HmxUiWP5c
+34zPlF51YB7CWxpIh2UWblpaKWYfJcpgzmET/DD0OXJa1daMEP4v0eVFbfaU5cC
E1cRzSqHVoBcYkxHSnDFMh0Rxs0RfAJmC5hOwigPv4mRw1kCJ+FLV4ZDFMP05ekd
WSPfyNXBR3FjvWdGQ5ExhGSC9lkL0mHo8pSMVRz68b7ZFU9S5+YIvzxYNdyHRXPK
TnRm5UwqqwZ0YTQj7qa95on8aHdPjBbbJMom4NeHbzjGJN5Ycq2FP8ttK09ura+w
z/SwVKPBNjeoYV3LO+nUsyVFNq49Cm98LArghrbu1GoESKbqDYR4dAnR6+lQjhei
g0LzZhVTO7b/Ta10I52AaAHNwjSvn3/YpEEKmgQsu1+TDfLZRoCO5fe8TRGvzz9x
hbeoc91iwnk6PrsVHWJBCBu7q/8ihFXrnjtEJ/yVRntOrsmMu0LOHvxVJ6Dpq30W
xBIeG7SvRT9J2RFsacEldWCQIvad2EhTPCW4vv3untvXzP0uoJP6ge0U8FcX/nUX
TYCoP/7viE1c5OR1gq1fx81+Yqfdc6fIa/kOIYKMNVunuw1wRZEt+Hb9QQL7j4/m
UIhEJMF2n8DA/UBgxLcj6GXX4OxxTVJddqjEwYzySc8zaF/9PIqQ9LkvwCnTytQ1
Mz/edT8S6ZacrAxhf/uVvyzbPqUW/iM4lit1C0iZGFbLZqmSHC0l+jUpq57XD+UZ
Cf3VaZxWT3P13uOFz3PSYfmi3GpTDIXVFNsvncMaSv9clJA/NBO86o4kZBkmD5P8
exqX1aIxseJM89Y5ztvf2+t15IvDD8qqDnAxw9K/jNGg4wTVAroB8fztC27JhVjc
Vtc6S8v17aI+e+/SN0S6ix3cYioWq+iBl3PczdLrmGaa4iUxYv3iKm2YFDD3cZyP
TG7P1OAqgqylmajObndBs7PmKVg/j/vy6YnkcS31Y673VXucShf01x35ewZTt9up
wtUlMV0nGXlF5GBuWfvUnGYiXb3UegtI2U+iEEYm3DndAnnC9Bqkrfuvex8niQXA
7gwF+ZBMke4OSVho5GAwOITH8s+SsRTL5g8ZkAfL0Gx7ON88OZmdtcAHMW4wcN2r
L9ymJtT2lVQL/ck2nl5+rORhYh3N+/hOc92T5UFwXmxpAi8ifqwHK4ingjz9LWCx
3d3iYR/fHU1k+MlxNiJJMqFgw7mT4kF3CTHDa8RQVf4/n5Nut9nqBQBcr+Ep9BSp
q5DVrQcH+1VLBPRDWGqOsYNfBDYRxS6N3cRolcT/92nL/v79zMqqk++HIwaqUmyc
u4cFLW/4oDTJ8h3eYSh71Fbwi/V4jm4eUj5uijLiRA6O5vYe4SPsldo6H+afzSB5
VEAXvQ0emaSgfI9ExK5xKdoVzbJa3vsgZPXVxZktQFWzoF+VjQL6c8HiUx6MjK3Y
lDdMqtXUNmYuq1WJ46/fZFfkMLlGP25HUgegjNnfenO7wqkSE5kF/e29TsE/lasH
+xsxg942YQ23UdOW9igQcw47qb7otS7LCIkd5v7MhxOs5sH+4JTHPrQoFyeg24ZQ
TSi7X7yYh0mt5V+P1y+bLSl8bbeff2AmJcnufsCghLic0nE20bleqDtu+C1kcvVo
7XTpFxAI/klYlv1Er/wo+GEAjNtpkoG/oVhesKWdHqyB2KpyTaRARLxaA98gYtlL
oMaa8kaF/CTDuehh912ioMe452fkvGoxv2mNJPE6BLXsmBveDXcgGI28rmyPBoU5
egF+BGG/iKRbsnFG9S/0pMR4qywFZfnFMzEpy5OYqnbPrPrP+7aR1AWa2o3+wms2
zzKVKn1Oh6EXrAkyl5UexPPsTN2M40VqHHTUdWe0A9yjyM4BXATceIgLNvcrVAN9
OfL9jxI87C/st7ch1DXC2OmKtCFAmfTE+Z7sf2bt6dhNtDHx8aiOyP2pxOpG+4as
z37FnfkjuLXXj4+QbL5hF+OG+sg25vdyTTDbvWt7oV89tl2oeqhj64Uh+8+uWnbf
NyzhO2yyFSm/NOXaZ58UQQMG3iNUH8XRTLsekOYEiE0Xx4NLn1X29J95qcV+ewt8
kRaeXG6p0d+GyJ2RKZ8Do/YR7nZECsXPmdOMKi203nX9piPG1F9j77z0ffXByKch
mpiA7TLI/3alDdiAdkdUZU39sEsuvuwB8NXHuwDKHPoUmRWJLktCvCrMPODlMU13
hrtrG21uwiFt/+dlZ7jhtbMyVLOZ0Ilm484auIKDcxT0MhVLIbCXUcfmmlIdC/36
fQ/9Psb9+kswftlzC/tr+CeLvcRDxCOD5zUap9WFuXxJ2xTEN3Eg7YPyZbdvsZc0
m+1UqrLHwPvbDI36iHIoX15Ugq/lQMEaQ/POjL6DTv3yHcTKvE7E8e0RP/pXUx7J
YiB3Yk0Kv+xuVtuLyVEwWOKpSt1YVfaIk9DKNUdw0cGSSwNe9F6KyX9HtBWJ3BlB
owUhneJ1ssHW60dGCwXmcI2dzOG89Ybso1vdS7Q0TUlsNeX8Xlf7NGARtyucWMxs
ZfJJ8QKpU7mY1Mi9PCJL2Jxw6hR/eVkt2ZffCbfsY1x3VtxcGOu4Quv3/KQwbxtF
+1k+HVurTdvXBFXT0+Nd8skxPkEpO/Q5SdbJSD+HFO0yH3HGzR/5v+FyU48YRbab
utGlv60EESnYyxGsnkq0BEaWlGZiwUtM9tljSPHKyZGuORkdxOFDx1bKuaxHtIRl
LktIsILoNQ5DDv52yy40LgmezyaTIM07RyTNQYJq6bFnFH0qV0JMaYX93rr/1ihT
5YpxYkC9hcr/DfEZW8uIECc2X1ffhQr1at95krlUe4gUG7yLc+6KVRgfAd1O2eB5
lTg89YcbiSt5E/p+FX3Y+1s2AyNwGIcP6tFO7Guf/qP+XW509seCdWvMTKPj+/4X
5xFbjxhj0W8z3DfOTPhLofbdJjbCvTE57SAHm0J3aEzQqbsWGXwZc/TTlB0jF5Wm
zxFK4gScRYQgjgJ3x2rSywbVQa9OYGJpsNfnPvgS0T756VTcmfPXsjrSSjFfYrJV
W88veGJH+BSOdyBb0KK9IFqATbBrE35LROKy8mCeOZmcaZW8Q0zdFoLVYV0vuZH4
1gYKe2l6Mtt0RZV5eF+yLqHvd13UrUMJLml9QRdMUAL9aglgySpUa8TrZBKQT1VQ
kBFnK/Vpijq2Vwyi9PrchlQmsxXTvr6ZJqDJxMhadnc+oHBZAcIUBsN7p/zzgWsw
CXwp0GUgiKlNmJ1F4sBXdYxHcQ5IBGM0n7JWutg6UajtDmBgdisEYWk51rBOOFYI
aSUK9wUIF8wzggkI1/U8UyE0/w3Vit33LY8VDiFebPc20je4ER2FUhxehvUPomIB
/bFmI6+FqsvcREJcw9HeLP3iMX/zY9oVyihRxrz3yg+s5Jsihdy10kMRAybmomxp
Nq0LkB/P/IhQOdiXDtFVZSw6WqZEhM/OzDrdqy8x1/LMFT/TEMklsHK6f3lSMENT
hU0EsJyHsjvFPLpNNR/WOH2SEHPFK5S6Re+5ZFQqg8sfZKWaRe/F0Kok98FVBg7t
4YpQsP4oIENMwrmgwGn+O+zO/RPVnas0mggz9Dg5Zr2JHi9joN0MPHSc9hmlJTw3
EDQ5Ehqpfsx9ZL1EjhKf1CHSpuWzs5pdgm1mxl6k1dLiRtCFek4BlIICzmVDfCQO
f7cHlbyiI9BxMyaUTlNUf01m1GIo/y+s/QDD6+4dt3OG0b+wAiw4daG4sSgNkkQI
it8flrYGy52jXJGWfrhqRseVlUHkANPQrhmLk2f4/2UffCMjRqSeimD7d2HfASNo
/qOvcMIjLmq+V1qyygLpvUMkWWMTnTS+fM7f/1wijubaDz3nDi3daAdJznmGJujN
vqAQxC5yFgHZwRjAtGeqbHtrmebSMlUD+Sg/OkuOxEKuEkI/vjoQJM5YMwDhllup
/iNXh6MbpmrM3ip/5kG/qlYXiLdl7R0IEA5EiZHk1YGbmKaT2AdrB1pwgLOD4NL3
Jzgeat4/LbP7Jx+dn7r//VXC3UawSzdvB/IOx0KPMVk1vPLzc8n8iMOUNwF0Decw
I+2+svhVXQUJEqd9ywbY+XdB8SAOMqmZXNunljsaE4VjcBnbsY5qZAHJZ7u79EzZ
MDs1n86JpBQfMoLVxHu1tNb9immmMxLDqzfAMMkjamIzBOo3mq0hnXevz+MUR+Ii
c03Li+Ea5CAox3ZNUfzQQV99z78bX+SHdc0SNM4F+z01JDCBdhnCtMaOp0ZIPnnX
8B6FDMatlp8EzWY5LnCKP1rpcjKSfQygcp2aVHstNIPLLXjA+0JikpQUnWnvzCwi
nj2iWeopq5+OiLDdxofUcjEOhXi9x0LRcyVFR8l0DmrD06pBXa/ECUkarKF7Rf1o
uukTMKQ/fXR8IDT0tc/mU2I9TBlTlMf0otchXs/sDTtaNfFdyIRyZtxX1af6Rd2o
wCt+9Urq78KXtYHtJ1Bn70eSOCFIrmLIHufYDhm4IgrpCbnrXHwA+KdmMnD4sCjD
+P2dV5zHZveHmykOVbm+nkLJCSOeqoMFkB/WiWY1MA/3b/Grdo8HuA2xyDCdnBgi
8eZ9kCWtUUZYTK3g25BoS9JJe9gmGH3ytmTdvLsyh5vrPeoPXxW3MmlipQomUrVm
ej8TDB6e4DdThS99PZo3LH4erSc4CcTFAEGlkZrH1+IJ2hR04bTGlZnpPeFH8SVo
ASrl+Xe/HEI4eJRPXixinKDWwXD9c7d6UTXDrvQv+oLNZOsP4XQ96zl29UIbM98i
RVY9NKERgVr9jx4vfOj7y6dHTpQBCmDQ57O3uI3fImdlwL4/ala14hqd1qwB1LuN
/jQA/lDbCmv5s6kpHC8Q1aFZsilCAVLEocc7qryUJ/hv9w1hm0VPMW96MCpKeyDW
iFO+h92XOSbMV1Kmm+YmoVs14NEdBlarn2W+KNsrGCKowFNvasATRts2rBYnuWIG
CuRvZ7ntvk2zUjgwkTvgmlFw/7X/oqBWQpJg4l+12JcaXxThrgO3H060D9cXDFt9
4QEYOnZvPFW3Qg6/2DDAmo3U1YKAr0b2R5h8KVl4ymL56NdfXkW8JzbJDX1Ktg93
LfH1hGLrIyuy+BTCRXP83X7Ksu7kPSGckE4HPrvjpwlg/++VojhnI17h6X8OmDmV
s/VP+5g7GXX5lgkv3xIhLfECax1y1VghsTju5mljGdMc2cTcmeZkLdjuROg2dJzM
Z05bGR5NH5UdW4abJKN/uqwwnmpZyEs9HGx4Bc9TKjC01bi4Jj0zkERehYc1lwDA
BlLNf6C7ltJs0xEj4L1NGIFA2Hr7+26yKapQ3gtRiD3FJwPTeJbJwgodhIwQYdWX
pJyIiiD1ESWNqdzKqAeaGgnCT8XdoxATodxNMf43OVX5mJR9LGePqLfVKzR8Kqmb
QrPP2dREfOFYzqplMR0npuANBrFf4L1IyAtwEIvmrmo31/t0UrELyZi4ii01HrEK
ErhGCx9VhRB0nJE79BD+pcpkt+SNz5vualCcMl+M2ejt9rTRLCzMwnQWy199YZyK
Rrv3/rOQjkanie0rLRePxP+Tbn6T5X/CTkfHyde2l+Q/akbOtFgShi8/h2iu2TpX
hlfzlyPHwpGs/kkox622J7pj0cAmzv/5Tm2Ok8GOMRhxhGA9/cXj0JojxKlhnfG1
rJpoEz7QU///Ug9kdONTbFATigJ6VUH07QgwW38QDijRgz3giw5TWc9THVv9WRyS
bn5UyhpjmYwTWnnqeTBd3FE395HUSRFqvjn6SipimS7DVvF1JsZNncvuNemG5Lbe
FO+SRVvsCDPL/shs5JcMDroUIp98kx415GdvzBBd41gX+g3BGkT8BB+FwJOOWPtR
80kHDlvSLNx9gXHmyAijL/IGV9+hb8vP9J9PaH21KOc0mR7UzDetXiVdp6qvhWD2
2AFbLQYsan3hHFgEvVaoX+b4/+P8vn39C+iJZO2VKkBVETL0OB4YkrgfXV+Zao2r
OB0/xaAbPHRf7Epcp4GfodVkh9GmTXVuTRJyQVzoZskQ/+0i1DdSmJUWR7Jm5v6t
GtBH/plyaJVu4dCk14BB5qLg0AJlrw8RWcVzFqEeD5/SrzjOQ8EqTz9FbHqsM8kq
JF8N22IZIeIDG0uONHW3iGuvehMDA7iij8lCORlATbckTGkSVHPCdZ57FhsBjAO/
8eXWp+Ahj4DClw+hbXSg6oD/Y9QxhdDq/DQRE3/AUIvcan4ibEhrtgEIfW24Mfz3
7WzWM+Jhc61Dz8cfc4gKzWFIKT8ZBYNHufigeL8/zBw24kB7GC+blPK+cNUHeA6x
xW73e4KMuPqj8WI/4gWe/bOOPWBK4Fvc10+hD93bIt8HHlBMcCa88vhtpztUxgwg
1up7xtzxb48/LTQZR9NFaKWsZRDrcfO49CY2/GZu2idzDP/woZIh1gLOjbZUi8hS
2flRHln7kq5eGWDYuT+VE1UgmdpYDWcNpX9TgN78rgJLkABHZWzq2JNYeSbXKR9m
w+tO1n0j0CarntHrZboBDPO1qABqeCq1F9IPDgV2aVKNGNUHiNCS4aAFGvc5/40z
f8ryekPf3+VResRFU0lvRnvZ0pengnzEBq2DlSowjcVJPcR2j+7RsUQa+ktWJfBo
gPWfyyj9n8T7sBzEMbgOdOElwQxaLfhyXJrIg/cQfCYmamZOfvFGrBYvTAyHHRPJ
pjzZzJ6SkjigJCpFztUgoc6NubsvgTSh8qux3QwQIWxDnecyNxSDdBKOO9uhX8Pj
C8Ums89BdnelVq5ksNGFyFMuKhngu1LIuw0vmpef5suYj5bwifTmgdmd4+bfOZCP
UKf/vpV0/8e5FGhbVIAl0PkYFGTZtQRKI5QbqH/430+dUVMtUo9CIMXichmORaGk
4KzqQH875pmBlH+pw3ZdS0f88Dmm4O/FRbaHlHGl6CFTql3Rjl1OSISD3nN7BNW1
OsuDTpWd2Jod00uIHR3e6u6MCFMppsAWk/FXQ3L9nIKzPaXvbnw73ZyXJWw8SXID
cp4R5RLIYvgHNgi3t/C7T+bYPV82Kr7gVWrK9BbKM4z0Ht6HMj2H0lekiCS40D2H
+VRIXMJ0NvnxUnQ/L3YKZN7haOMzJInghlx+X4W6e/xZ9b1eXmbT05SKlsDWPsvJ
+zPCZCILpj9m618WCjkdrngl5xTj0Ol0DB7leY5M9ng3U5c+DECcfwgeKLgWXL+T
MZSAtzyYv9OcmEjCbQCb1FBIELUkkvdZcpjqWcn80wsrgVLRgi8tdR9y9WDND1ke
/zDQZu8bvbsdtQNoQ20HTK2ceRLoswSi+yWqC2J/Kvty3uGFU8mm4FM4PCYGVmpK
XZC7tN5DAtuI6MYvNTiTvpYdIWCiUbdSC9Oqpvr5PCQWqPAA8GEqtk4oh3HHuFze
xow6YTzUEB5shg5AddF/E2DCmHykVlzQuf/0IYh6jvfv56WCbQrKQiFpb8znXW7p
tEmpaYbw2YmDwZA5kRzJRCdd+JRSCbLpcxvsCZqtY+vZnQeGJ1OFiohKAYd4AUPY
+ttsXRdgs5lf1nou8pznkiZFAdUh3MUCKV19TPyIlvTGTMoGeL7YFS3bmmDTk3nn
MDWCgp0/Wi3MSubQoUKintMl1NjW4POF4eJXDqW1F9K4BHZ1s4bcB9f/Iu7mAnj+
cN2q5qXd829oJMsXBsSntZpxhvWughZp3tOIBKJrONJ2YXqhwvJoF+uyCtEkNBvG
oi9iiNHPeHXkAAZ2njhiVTjUWLWu02MW3Bjn6UkMF5EavPDy2MUUm+g/PkIRhwzI
0EgYW5v+4dwF6jSAevG2mRrogoV2SIKpMlU6UZ32cC/onHUYmjUA+Jn1uQj8RByK
ZWfa449nKrYNDJzWA0Ibs4gnStCWTkJ74eoOB7zHSKQA67ly1o24hHJdcu3od/al
EYysMP8SrwJawp7Y/9xePGqduFogNOaUfq1EnNqCpeQq9gSrvoMzyskUpEWCdqNY
YK0xBV50t3VrbW/jp+e3aC0jvs+/caY68ZiCIrYmCXq5lvRLe2eCCJpGhv0oXjuY
X4h81DG2v2sbgKw6hN4bmPPlQx316FWb95MuQv67sooUOLd2BeWfAgdo/HLcs19D
iaKLDDqawF+73rBIpg5VLyYrUF6Zr4apoWKh8XZJxgTe7+ywsXToikJNiW+MP+5I
WgfoyMc9FIqrSaL9dWxCBd/LCv2fEhQXNb3+dtBVWgjYW4p9edvg2vqht1MGXZh+
hKDCvaWo70udL5xPsbLgIFXitC46xXcm5F9TDtG6hdq6jDd+cAaVLnu3VAY/DQVa
CUtSVi5T8HCfvCERC84UKOy8desj3lrlk/jjFseS+5o8Oht94SNt7n2ULASEt3M6
Km7TNu2UnLwU/qaDdY4GdhQttm6W2zcnBuQsowcdMwDvU2ADlQUHmPCKMrCuXWXI
9BZlrG6DqsskuaAL4iUYIFLz8GGfrAecmVuiNY1rMhF//LG1QxJ2gRsAT01yha6E
Bj/koyPF/kZzBQXpFt7Rl0V8CWg2mCb2a5oGkLuRCWYxsGgMMYcAgafLEQCZ0TK0
sgbT4KPI/QAZFe9g5QbAFnWZGBARCDJgap7UHN/1g8FVZBiSf3K2wAPlkMHkNDQs
M2DA2hcK0VcfZSinftAENsSJ6cSeMHABeiA+JNd75hP85R5RPTv5PXiZh6g3FwpN
WDEm9ajhC9rbAK7qeGk/KnrSDKsV5K3iS4xZQY4OKGiGZPykPvujoE9lzopDQOcF
rYYNJ98+dduUeJm6VJJ2M+VfbEAUxJzM7Ei9QsmTiks0yMWazNp0AArgy3r+tHRt
w168jLTpxnqePvlAwqRq1sPlKeEPgYEyycdHR4/9N3OJty6SS5bG2YHP6Iz9b8v4
lPr2ezpJRsFKPR2TA680WzE5nkOAOcSu+bsKAIrz4k5ogGL08O4XiItwUNp2NiDP
P4uXhcGdnE8kTdh25HNDbx8aq2fznesK3ST1hsaAbCguE2fS5v/ndzlfolD48B8F
yAwZC1I21YKgEKhagEHJ9Aw1JGNYbHwCbxOlEGz/CCfiYKyFOU9J7g85QO4fe961
QAz/lSaJAO6aZBWZaCLmxwPB18AyITEAHD4i9ygQGWhbkBCTK0B3/Rj1V6sGYswY
qvqj1GFvOB97lr59a2/IFSVsQsGi83SZmZXj9RnRukZkNPf5p8BNvwlNqOWEWXtP
9FMO3IAPD2rEW8Y4H6kOWdHRNeBDMNOTOZQOIXMZjtAib6yL74aU17OjkG0z7ABM
G9l7+3JWTZxGKOM5ZTIU3HD/HnBnbJV1lLRJrRQV/VjlQsS2aa66k843wN766lU+
t4b9AW/FxfsOEkKL5Iosnw1ttPU8xtQurrDuTjNGjHr/1JWW8/mcOawFF9/EtWrc
PSCWwqDGf8P3LGqJQ2SxvtckcBaQFKQiejYhiokceLHeav5/kuEGGGf7GvivdFtH
gyT1rDFR0RKlcNJdIWB+esoQ0jge0wiYpA1lM8+ojhHUfrKTIMavjbNIbpLF4l1v
vMSChRSCfyzMWeEjJ8UrXCmhl3JS91aSS2LNg+hFG85SdN7a+JYHtj+Xgtje0jxq
LILVG5/POuC/dr142I+f8TnQVh7s/E1riupd1ffvfQ8+JPuuhY0ea2jryu89uL1l
rOhEa7QP7+T8tBIAebq/CcF2eD+rTwPytM4l3gCjKpqd4hngZoCZHYGZ62+UK9ez
y3gX2K95vUZTYs7Lk17+B81CqwaJygcWtL6pfyr7wBNZa/weilZO4s2doiibmJyS
T411tIv8Cd0vXJY/yCaTSkbo/q8m7VM5RjIfCuZ1clrDkKsvBRp3JpWiMDN9IYUI
WVfbcLj5MM9a2tNlsKrd3lr/Vgmz6mmGGGF78ZjFr8xlKqRry31eRkYdcQ8nMc0D
JlqVNlNkMS1Tr14mMvylcalwpUE2y1Ai/CtQz6mnIu9qEKcqF+H3RUoTVw5C+ZLi
/IXsJqbDqRMzSgICxJ05UcvoC2EuAhUQNVkjCnr04Mw9qUQr3MKgPytbwPKiF3dy
isim1+AARfA3j2h84cJFXqtsuCxsLhjHNI2PwVBlzxvGfJAKIg0sDdGVrlu6e3J4
woubeonVBpSuwr80fh1xfKKU+bJ2ILVTj2JEtqLMZr5T/DuNWFi6KGS053kU2n9d
E4V0pp8FuVMJp+4eK+nXL4i3DW00KqWeYZqr7W1c/PRKvMhSBty6TiZE421NVDck
+EH9nu8nzgTXLM78sLSIClmACkR4gYyD7GeQoO7Ye+tmYym7qiRQWlh1MkFriUsX
kvgHb/SERVpqMkOnpD7Vy+Blop1jPY7ZOquaLHphUIm1y8WTVEhJSx547Db6Jy62
PUXkeU+63+pMs+4Y8EOlU235jO9YpHNG8kAZQvt59XqpP2q3SCGYmhNYUBW0EdA4
dLaSUpGyhIJLDBUVRu324Gz2ntWWMv27lV6O0xND3YwM8IFPLzUrlvDI/koDMywt
fohDqrx32DTGEtwh5/S+88YeLbDBfXKBKU+R7it8nb+7U2x6kUO/feJo2Sr+B9jA
Izas9B5mKMgrfqv43H1CGsuqLGC1w39Y29bpIsNv7NI4wgS56X0XdepLWy8PRHp5
syA6nhLHx44+ZyR7WXeV5Qo75e6FSf1ZMZXm7d8j+mTJs+yxYlbUbm/Xsyl1vODs
wOP6ip3PckGMe7VnEbMMlAIZQc2Q8OjSpKB4RUJSDxc2zCc3dlzT/HONrm3efQ8G
rpPc3suHb8LAdMKMjjCtGhitcIyWNN5M8k/ephUEu7cQzlHDViC1o4f5xUI07xEJ
N4hBBglBf0hYwJns/F3uIIZ9Wt9uQlZqIHBCq7+mNZCot5FIG2T8NwWdl0Fo/qTD
lXTBjFdG0RkhArY2YHZzGoYQDfXWm2m8XvlB5PXgZc6g7nz13bvMIaMBmctJ4wXR
OIyXNhJ1924E6brXQ+GXuq4kJgTsWE9WRujYXxou92U3ok85Bs7UnFlJ17m6p+c2
fjItC3iq6Mh/QV1822AmMEznkTPhcd1zuFfBU6pKKP6dDQt4GVBQxbdqD3poko0Z
m7yOF/Dwu6LW7trnPkzmQNsXORLF5lN2TCOeFHSd5bSinvhLpKzkihkfC5GmoHLg
gRwjfuSaVzDa7GzcqYqcD2M1+4518UiVWhwsBmcy3eb+/S7Cu7vzkYWbXyKXbhYx
toqj1ok3r2NpqeN10/gcszBVaZRXOg9qud+aMcZ3qPapWMh9eeHBeiras5ZRaZKE
2iiY9Ce5Zh+9jHtYxDmsrSRBmjVgsuZCsFk+6EXob63B2UE881r3EthDnDgMYSfj
2M6Rja6BD6jMoSNA9PWc6MdFmAt1AS0anjLchvh9Ko7BW57XdppJe8E+gBKOaTNW
7bI0fobcIaUsGDzWd6gZD4W4S6y5tSBJ+aebI4jDfBvt0rdxn6ViaZQr6xcDjYJU
Z+2++bZG9NeyVfOO5ZuiUyqVmc2fLmWFCPGQ+8zLwYYY6rCmF3OrN8jP0e4MheDq
Uz8LeHspoYBUX/O0BttKpDuGdvWrzV5ZbnXCFUpENUVwcEdSIkkQQ8UtqqHDD8Ct
UAq8CzwNf9PwJndjk3aH3V58ECpDNovbuVbkKLgQMb/GdtVrlnN4VR4k8TwjSReV
jS3gTqxQWl02eqJGlTc9/PCuQS3gJewwRpC8+PpNqvbczKL9T/XtNa5/W/jzEBqk
RHrC89JoPblebB6dNhdWGJhTEsY5PfQMBBY3NEh9QAl7CF3v/NhlQjvJN1xyH9lH
Ryv1Ry9nCpD5YNFnmu7kZVMd8Voa2QwF/ac4wFuVBdw0WM7qt6EneGMoCj6do/ux
XSKS2wEo5Ab5gPaPG1wnrNI8HKGUG90KRzmofIYYJAmuKnAgw1c0BIxk4RKzt/8G
kyOEm7ZRQgbsSb5JtYkYs5aRJWCH47EUqIm2gFHNvmccYrHB5Gp/bE2O9JVtHisY
tJOF09IaMFBnSl6beBb30ZfrRf5NCllAQbI2Mq4owiWUak5iVZtbXVNva22t5tHZ
pl2hSeXoVUlOrlOsto5yx1SJWTgHDl5W/I45ppXrOY62DXNvtQGmLB7As7r09oCC
HLanRvSeQWyLfQad1LEMSFM9L4mZ5TZp22VYD/LM5Cn2vTHNYy4savRTEaXc90J0
ROczEWeB9DlQPP7qgJIzXlbXHLP5C6o5EX/xSwZeXsVpdl7e/nZLmsdcqYuK7vy0
eap4Ej5ST9D05qegb02x0nw9z1v075gVtHDx/ht62ooixM9vZhPdl5W2+78Bvt9E
Y8jRHLztc9mZKPAEb0yUtdxgG/5/So+EPv7IcbUepvBmPNpapIX1u/ukVRHvw2sc
lXMRHpVLckcnO7d6xbuH69/9LPcpFU/naRyrkjF+LBzZ1ZPleYOjQMuurJ+zHnzC
YOjVUE0lK+cXxtjglaJG3uRhuIxrECzIsnWyaZfEgC9MA/RJkXgl8lX68AgjvhsA
QOCy4hGcjlvtiRbUUAMWWkB6bSJmY4RkEOArnr2ZFScwG+Gsz46FKs8JGAeSALbF
4cLgYEqUkn7jUDiZHIrwIk/3RnB5lsMgobJUmkvf6rzKk+7RGoRtbYZ2d9n90b5t
VlPmeC8Kef7GUkEWMJdBmIeTj57xqGMamVRRq21RnJlR3pBW2RRp0W9jt7CXlEnY
+qPf46YBWjNVpJlZA9ZWMz3AUXVdGRzU1Vkd98aP61bRz2rszmWArwvLHjtgD48G
tZLIW01SmfCD+s2/6jHE4t+wnGwwK57z5DAUKX+x8P+jgemnnj4RQ4qiKuYWz2XD
pERrxB1yTMuWOJmhTjETnX4cUbSrd7QZQSkYlwvEzAesF8A8RVF9Hk7bQwD8fNNO
UwIDuE/tnCiYIDFHz2eUpSinICaHiekXEwLLKB4L5t5NRRQ7eQ7vh7uF26b1tDSa
3jfX8XhJ0ZWnxvn22afIFIg1wy84jh8Q5/OsS7YIoHcRb0bdLPCFvJSBvX07d/kI
03n9uagEN3ADT82zy2rQKMElVr9PLGgaMW12rY0clTxdLZdmhZ0Jt4jQ0yz99abO
CX49YANu+HEjMbNINOLMerzyZxIHSk4+3qRA8j1lvQnrKiJknxhPfqp+Gxysut06
+9A1XZ54vOoQTKbhgbhlkRLLgPiwKExrz3P0/Yet91MIVsal2uXL2GhAR24GQToM
7GYNeDVlsQKA1UbKrNdkKRuoCTq/hrFBvfDdj1JVeGFDSbTShg1y5kGeoBIaSOW6
/+f24jjBJzOjkUCERlm1Nc5p4grg54p84gPB/bXb63HuO5f4viVRvSKUKEAfVZU+
QGFlF4KRaH1bcyWvfRMIpZ2gijO4h9/i9L4DommhX2ZxqNzVfkYP6bb23kTnq5RY
3UX6R1TKaE31cKMiaz17rFnznyZvWz5597fNhFqM8z+pnJ621HC57vNGWuenQ0O+
ZbSZr7lYUNE5YtoRat656qf0+qVDnNRz2idkQu/7FJ5dn0QySszWLUyKtPYAcGE7
Vp7sG5VR4JSSrFLXZZjd7ANL3TcuoXNJHWjn0zgGQmJeMf0QdIysHNqxLC+9Pfxi
ZKET171KTmaZQiGNHOyIrS9oGItcPo5jMULnYpbx3r9etgiQXM3M3hYF6SzHrqYD
VvUJ22rUm6xMVVlP3WCXeuiLiQ6RMKNestT13s6/XLVD1kok0YNGbAYiXtWj1pGM
1HRbjt5eLGwies1wUQ5eQJVJdSbFAnHd+Pd4wDdqWRREHBgOwN0l0b06hI3qXYIJ
orkJfNkb+jslniG7GHffgVBzKxbDkfhvAN1zjCv5OxDPN4PAqt2AnC0Ms6wAJxM8
HvF7rOB/XnA2RfNN/JbxmhNsYr7Ns/e7Kh4vSvTatON8QXLbro08TcU7eBxOSUKg
Ck8DqzfcQJ3wKrdf/3jkciX7rnTAf1jCcQ2/2B78teptrhKno4X5bXdz0NDvZzIz
CtScx1hZ3GzOk+KIgMwhYx0nb3vZBStK/taX3usibcldg+x65PieQZJY4YZsV85y
zvDal32qu0u6llFg4pYsdv8VzODQAJ+GXla4MC52TSWqw8Sq+NnbJZ+jvA9/WWju
pfSHpKH07cY6d/DH4GYo4G8poWWaLTp6lTP7om0kdQxXL8NIK7vFdIOeF21rRLMR
DitibI1csgpJ6LWB2eXvnG1LBGnF9gZTy63zvlmmboZ7sXXXEFXx9A1YrAvAbzpK
`pragma protect end_protected
