// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IhCR+b8EBuWC6swf0QOjAk4eLAdp5BsxPEyW39dnoltNr/yZCQBOOVcH1TmlNJED
VWPyb6qetECGa9C1OW5UEjh/evZHleUiTwAbTI3lMekm0EQXKIjuyI0PKxhztT8b
9h6J3lW09dgE4WZL13xxNa6BOBYTxRDHzjho5Dj0IiY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 133120)
3freSoZJJMk2rEK0LXQmNUlH8D/cOzeUc2c1lAXYuzeIifHUbe6OGsIAUkfUuXpa
QJZQl1jr9eVWSng5KdOHdEb+jRexoaxoCKIya5K7Q+BgsTipjVGi62Kw2EJnPsjl
DOsnD62VBFkc0qDKxkurOVaauSnAS08SmhrU8iVb7dwvDyG3fVlcrZo/IP8sQL4R
YbpChyeonV2N2pCeKFaT3CE72DDGH1ngqyIgnbx3q8y/fFnzNxdqO1rNNW1MEc+x
LjcTIakNJDjnt2h56Xe8W6PUQy2AW3HHzG63jHGsJBn02IwZGzNRnqOKvEvE7IWG
2X6nSdZNHI9B37LiM9IDQjWq6e7YdeJRF7FOHMEm28x4d6ChDljFa1+d692p9sux
/lTmtnLmgpiTRhnbZuRny0/NAewZuShb/s2XrcwVrpJAZbUu/aidOUsyZJyIILwZ
F45j6bsY5eQf9mCJ3h39UUbr6rEcPvW1I8Lru/ynvPAMqlbh83ahuAXPjYGyee05
gv46Mi11U1cVyEC8FuMGvjsCFWbP1t8prFT70S3j18jbHjoNacMb/VmYEDE5W4Me
UvRFug7dMpsCBwiNzb++wi6hRg9kMqQf2oR4WxkVeszmq9Z/TDNWpYdkdZieEytI
CU8anRSwwYIx6Cq9sZMA9VZZaXkMzcsNY7DUetC0AW08JMxzWiKAXCNLi4Ov/6Op
xCnQy/+0IA1k144UXtLrdLJSaa5wlqOZhPGBCIWTWlZQ/jLmoKYSBlvuSd+2FuP3
UWVVf6tURrQEv98aAviXr5U1yZZ656Vrfx34BdYZEw7uNrkbpRq4HkEKZV1rU/95
NQjOQAakAqAW1Wkr16ACaV2GSAyMszTmpELmsHEYZNUdjEWpfyIjzLIMNpv2Rep9
kC3cMphFQUvn5iIIPE4Wlx0byakipWYEbWNekOMLXMW7OCgJYtlE1JWoEUFwDJg0
v9YBB1ov7txXndCkslVUTWMPQl79fiLGoqP7H124WE0lFVta9WRCcwHx9jthG2Am
ekLCciHyiGzy6oFS39BCKlxt2g692R3zj2cCpArQJO7n/J8B6dMJT5l7mTwhO6/3
N+kCkawYVVKFammmFY6/ZdRGCsHr69WvAYQXD01GyJ437JyAMlOTxJnmP8lRuU9b
w74YW9RBowPhyWVcUB3VVp9XfudFwcYpWea5FNS24xAiF9I2jw6pagepZwkiXNgD
pFYKFQtLocXfpZjJk4ZnzBbrxCP6yr1KcQfcntEN7AXmBitDSvgtU9qqs/TUbCHg
0oin8YznIKoz+3E/ypQGORAx13aO8k2vTFHKI4EdXOT3GO+Cc9VfUbEjv3+6Jn4F
CzrUyLZ2NP9suZxTG59RhL1tqPIudfogt9NTlRrTwobalmlroNH8qrqjgsm/JyQm
D2DintuapqD8VuPrwUAlG2mQRvlv3YInbVZZEVBcQoVhnHm2sGGg3FekKuWgYAWF
hEEjoi3G7KDGyU4USmHGH9bFqlrMfbqB/gIBeUYDtYxTUIsk/t4h+/G49ZOyXn5l
rMdeKftuxr2xR2PathOr5QyVoZpWQg0i/pkbSXET3Bw+9QtONgY9VQFxegs+Uuid
YFFiCv0yOY3O+26+GpOlU+hj365TS6kB87B4HWaS6qqMciU7nltsDFmFH1v1CLdD
kwTsxV/HiSFm4MGrUkT3sh68VbYXR645PIxyxB9fcun1zYa1LC1ufI46w7syZqWP
TU4TN+yMxR8GEd/eHxECMRSU4rrBp8JWw008erZ2cc/0jvnk9jvbEB54A0nWiH7W
97iwO+y8o7B7xcfgxx7zXCfyaqOfGA1xOJFfKp/qZXzyJaaVvighMswq5G1IBRAZ
Btf6vUJqdnMdrjxzmeoAGuD9qaISTL4M1gOZEQzH6CY0lwzOkIjND+IGGKjwyxTd
aYzdSI5KpgRzYDZSJ8TiXthF57Vri5Kk05eXVjnruDmaAllu22drIR9ggpss44k1
PvO4eBAram7pDj+qgDNJxAr+RW+5RQLOW/ihvmbWfuOfyULdMAGRfveCheNHZ8+I
Gi7ntp5311H8qILefaw14uHv9C0psKGHgppcg6zPSK+0RayLqyYM1WTEeiAdq96Z
BxZCEtjOx6pLfJqKCuu9LUf7gFVnU3xZSTf9Nbxtv6FqpZ3OhTEMM79wWKUjfVFq
U31ayl74KMKza5OhjA+RzAEaKM3xA+u1L4b8iWl0lq4I9h6A9M09C7+DeczXtjtk
U+RZ+c3gL7ULimrl5j1Cf1fnWt/cOSCqJYbcfbjSikjfEfrDq2W2VqTGK9IDPWkD
BOYwzCYHRK9YAQqFttFfztZJvdtZYdkMJb7rmtUgC0C7J6uhpi6XVbhoKCe0MxJN
g8LBP3urkYOuvW/knfRPmVC8LsE5bj71QtHGnOCQ/CVpSHbJn6VsJlvn4zXZXnlG
1JzsuJHVhD7tl1okvarMFzY3F3v/eoFckYuEfRvfYioIKUCqTBgWcnKYw1pAHz86
uMfA+PK2g+AQUoSvBSczzJRcoTFfgfSrABjQzk8969QuYgHKvDaod2v0aDlg3g1e
vV2RhipRlDnaRsmG7dJlaMxytxTXFo2VAqbxkJWl+GI6D64/7mf1hP0yBsFjFvc0
W694Z+qJhThFJXT4Q4/n3RK3ZM/0Wy7LOdFjrDzF6X44lDrUavqFtmC4wykRTlIt
oVp6BmcrQpDYSdmUl9levw4DLk7Y4kr015ISGlIeNmfTuDPwlKRhVz+BYShuCS30
OJpdK/+640i1KDA7auWt4+nyhF52hCZvTtWXI9zcHGB6dOP8ZRRUYGCAWEp9fKOb
/os80HnEfgnqH7vi9Y5Kq0Z5SoQPmyICl8Ux9pCimiFuOoXnu2sRoo2MpTWH0HsV
XQd6EOtMWAvsrBHLd73u/pLGnswD37XSDCVhipWc4I8SZDikCFWrg4NiiYJAxjxu
JDyDoTXaDm1M6J7oarRDweCT1dCcYycZiEnGjuqDNk4ylyZZMKwbSkRHZM3OTZdM
FQ+JSlweVIYXb1JRwymIRFTfSHIuDRSFEvVSszaspzHsb6IB6HhAbE0cFLYdsSwc
S/yNbDmsr9s7HloNapKZ9l3sya5U1HwY5PEtzky5iXpwkYzA/nrc7BV5cV7RqZmg
z4TK/U+mmTh6BpfLHzyytDLEc2WzPOlxWK5uYpgjPH5qzSWZ4D2GwwecmhQ4qifC
6LWkXUS2Oxmh4yN63Q+LqJcLF6TENVWdlzRo3o4JPgxKBwJasd5NHTBuFPiozRth
rYULfXYv/PHJt8PeAsuHGJ+/urIN80QGcPLFh247nknpElikF+b+jEF9imlmlxrl
QvKlzrF4V+v2GgHBN0W9y4Mpuctk/Zi9lmafWVA4V91Pay+s7igTxGzYqdkGIsz+
c1/AfjkRsE9+D7lppTxAqfpCxcrFSz1+feL+7t95DQQQxzM3HBteFFWp9B8QP5/0
n8woOLhICZf2DwAnRMU5hM8SPR1dleYzmyDG2sQYYnlHVnRABhogSsJwwzgy0deQ
XUU/6dee3qGpz2zZICWRpSIFGmmbFGkhHxmy8iWKoMQ79oJpX6InP4Cvcb1wZSgj
v+drdsMb7bQ9Ni1gYv6wSOX+zBG+zO+CcVemgBGa8i22QZBGSVCUDB1BYWo01YVr
KaOcA/mDAR0j1AsZTNvP4ygrO+gMngYRFf7Cbj/sSSM9pr/RC93NACraaDCB6LRh
6yKJ8HMgkKM1rt6XnGB8RjHSscXtkdLo2BGNA6xpyTGC63eA6CTnq4qAiTnWKTaj
wl83Duh5HTZ5dg+u4YSo5q76pP9lVyt6Avghf5WDI8A3H2mHD3ZvGR61xPW65DVp
VMScdgVg5ggleFORnDXnZ1n0/qYubhGgow/cn7bthEq78Cl/WF6QyvcRclNCnSNx
BbIojN7V6W6Fv6EenptlSOPEXQj6oszwj8wPrIBP0aa0GMOk85oSjD1cGaOnkd8f
0+OSzVow05rmbiJ/RgSBhBV3hdshjoUwADKbKXB1jjIed5tM7vh4j3QsqvdcHcPs
sWbCrmu+pB9iFXFHYDi3+NaY7J+pjYShN5vZNptTrv68aXT7koqbxZVQ/bMEHlrK
14nvZ6Jp74ZggMadiFePcCHa43pHn9SorVpZTn6maVvSws2d/nZnCUHH+5oPbAuq
FZyCbd7SHHVXXnQFw53J0qctLPPyvrymahg4xT29V8fFH4/ajg/54QTa5dPdyoAu
l81jAvbmxgX7ktDjaWx4LusCmthvmZOtACSrjttI67IXB7C7WrerfARH1lZRBylM
tVa++xVMJ2kovuk9JPKnfMVlyk3bcg9KsxGwqOYt/QQXLZzDc7ZBer9XPOIPgctQ
dgrJvdXDCqVBurfRHZhH9aEhWTwmG+ZtahHKvRDm7HfcFaxlRgt9PGkxO3yVWbrA
4QZ5LadmLXZkGeLUInwCWCCUj+H4hROMr4VU8cr6zyiT1dfplTZJE+xJD+Url4ev
76SVTqcidsM6M29the24piXoUb7JnL9aD1W95PB2O85r7a6qZ6C3N+amI/Z5mE07
yezKCdOQ8TKJ4SREosuFPMIfrwp+E8Nf2AVKXNaC0qbEwXRutJ13x/iI3MN3EYti
sDZiRfmkYVzHFdMcyDmUkcskgGcXFmgA8woevF1VphfEB2hSZA2r0JOF5c1AanYY
M6LGs/bqHx1qIuhNehxJhmvrlTI/MiSkUL+RB6Iyc9LgXRHkaHujF+ppEd2Owl36
SfKjy5XjaNULUaSDhWDqvrzych8fHB/ETBYXmomjjjqyhqhX1K9XSTz+IbNTGZmm
P6pr7eG222BdUQ3JLfPtpxVZWY5Em6eCWS70UbpUIv1uy/55Olcc7ag/6XSqXnQA
fSBeLVhMFk6yiaIUIAGm31CGZYgRehPZ3zHVq0mUH5eWL+iaZplqN3uG9QmCrf4D
WAAwM/HbXjALYjil1n94Dtuh/Kk0m6ocp3A2mPq3tRVmw/JMav98xiNe5WPfqj4A
klTSxaijPkZ0PIg1f+HJttUhtJuSdqnj5CZ9z2RjZBwVcOQEmDsD0X4vlEKAmrVH
iopa3gc1nP+KTTBhmN6eHlV2q+NJRcfJVxkJzvc3kmY+zpQFOxrTBJjGPsgrU/38
zqve3Ozojx3jodRmZcVVNLYfyMPYtrWt6e0bnUq50M9EFUSNNzd9LHQ+E4onoSYK
FaCPA8sNrKqz0956FrdoROnPplepcYAvPcEI0I0Vk1BXt/+fz345wIRPluAU6BJQ
xcKjbmMBpgv+e+zD8ua9KowAOfw5DUzoSXJQmaGvljIsOCpG2puFpU2JN7B1wzm8
i9FlOnPBCA8BEp1YL71mC7runTw87xSXiemDJsUBB4/F8v+cM+lhHp2xN8+OxuD8
gmJ9HJjovxvD8jAzlR/GTBJQS5Rq0nnKaEN2M8Jki0tVvnPqyH1eL3tNNeeygnuw
R2VykJ4u0MWbX6z96ulKiQM5ELEiIM7PVUgojrhhKddIi92pjIv29se52b9YlZeT
tEgrDzFnwN1E/GxVw68aZB4AvJ7WQXHsmlpUcXNiEq/x+F6sy3heVtpAeLlq1AKe
MAuHJQqX59jALrOr1DX4mm6cWEA7+qErNt7a8DrqWNwCldzWwnCqQFifM80PQ9Ci
kY3eJOKEn/w+/Bb2Ug3mdtvmquPC5sWT1WhlMqZyo3k/w1ZFbCZReLSZGMesESTC
AgD9qM4QCxjeCZIKyojZRMuc4+RI+qw5tEKkG4T8f5U3T33yZuz203TId4029Glb
NXYaUtcWdqFTxWNt8yH+RghN/ALfWFjtOcOKl7q40Yg1EPE+O7l2Hc/oMAhaBc7A
IhM1O/0VHabQCA+ksufUeAUDMVmilmZAOgAkHnxS6KsEvDW0EphPqgMeRx7EFh2F
mbFP07qyriG+NPuLwukzpxZdDkIRJerTbf0MLD8rcTnSOYckXKiOayzioYvans31
rPA6ZijuiWCP5ma1/Lzw1ITbGPtCIG/wY3ceqI0COUCO8PvuuZynxmXWJfI3hWWm
L66Yr1uc9T/Ouovctv46WH/QS8ZFpN0G4a6/1eF2bZXS/uHOVFI8+xbnN9SWIqFs
QW8AgQWmoJUz1kqYa6OObUqZ7Qhv1r89T349MM5Qmu8lBZn0Rp3It4ymGq/VmQXb
EBdgRrYS5vniB0hfjugP5qiLFSVR3xDiTj5tPSN/Mqp6N3h0yj94+1ao5dVfQFtI
hMSEzPwyA1R8nb/6DE6itbk8bX6guf7NjTqQn4jNjcRcwDSED1iPUT/1YHyxEKwJ
KZyBzlOvTCHlOvSukSN7YGPlWTB6GFUm5SNBI0A4dCZYunY35bcLg5xePs5XAWTg
df94lZm996YKJgSUbmgtkzVMIDXcu16/mFJBcdxj2fZ2Otm2n/A1vXkQZ3+ZZnj7
hja9V0pf8zQrhHfcxENqyKbNlLrQWYHjGkGklSacRxccHiYP3vWfL2/HzHD5dMT7
AJWQ+GzkwLoqHdlgDw6C8sbmyjMRarzzV8eTGCeQziXTSzTJYWrEkai6fi9pipwG
CoSOLZN3UtO8YvEp8BdExsWr49o5np4RfJ9xvwpPrWst3dck/DyTap5wBeKWjI+T
zFhXQW50uqB9Snpi92Hn9UmB7cm9VPpDn/M05idv9T0jbxCDDLpgZcZvBcbShGPu
H8E2HcAd9LHqf8vjCFFr1leA9RhXfNkXyzYMz6B/v+QLB+uxqbX0qflGuGP96dvb
jPKg9TnctLjpX1QCgiByluTuaUGFjpd4OtO5t03V1Um6Oavk7t0MeZLNg1ZOcX+4
ySceY/DnYY51uEvCuG5m0WjojajoXKVnBicqK0nU0v0yN4JY9Z/K+FnTDHMe7eba
g0n5t1gSW1iu3jgQGKTwxB96iciXFbyWi0DpNU02gpUR/SPnpSuS7t+0cXsHlhi1
2YRbHCMY+eJUhDb12wUQGRqoKW+SlDlwTZVPRkk2g6bJh6wd7DIkeuuXiudNwrpu
0zWCLmoDux0LNek0/BTCooI00isCTLWdMhiCyUT12igQPn5e98642l0EwkJsPIie
ah8KsTilTwrsAksHp3+xRdB01AalJVYG0Dj2PqVDIDYEebRzmrnpuuOEVB53LeEA
bAejddUjkDBCtW8mV2oTGBDjoiVi8qri53KqSs3YscwV8jqT/jAQjYkkCBfuuOzl
ge84ZOs8nVcd89ZlWovMGwRbiVubbmrCfiLPzB4EpAcuTxLN2IJ5gj+1TxGblGQS
MaME2HtkeUhAiJTOYhNE1kBTwvbvlv7O67kff+/Qb91iyT427BOKA+eDoCWh8TlC
lWCxypRbUKeOUxphjKZmy/DhSNXn+oyCuY+AK+SmF7DzicZrtogCC0W41RQteWrY
UeeQVMuy8AEOTNbWhVE5xcELuMCeaovG/ODCjz3y7OE1D1O2NfArDwGv0Q7GdIIa
rl6h4EhxRy57wwsbihd7nIcMx+nIDnQ48Q/Aqgy538ZMd8qghluOkD3KhLhFA2TI
DEZoTEYHohe6frdXFk5VfIblEdG7VjTVZ8+Mjg4Z3WB+ZuCZ+HHHpnBW1/H/Ys2/
lEPpyHKXmSN6LYopNJN1g+w2Ge961CmvEpDV4A1SgioNRARa+zThgOb0e9ROWLPm
zgu8pbtG0GeZ1vFj54gRWzQDtR9kt6eeTbM75Um8CSPgwscV3raQOVd1cmul4r2n
q3glVHTOnSqMPdMh/C27pmYe0zVuRqnsn8wQ6Fceb6V1O5/mSCr7AJ4wYBYHneTX
24q2pDx1TSLxMAISIAH1UHBVL4Bccvo2sZkdo/DGzL4JvKj/A8ZmwWJsaOobqN+q
l2SHvMGBZXmN6PeXIRyiGl4kHUhuzeMsG6xZLXZ60eN6Boa/kiN6YMwXKFbf6EBf
sDcswQp4rEIxVNsLa9790ghrtGfP3VhvSg7df4eW6Hq7vrBOnMgfp5jYj6YK9wtN
xFN70NtMe4p8IkezwECLe3jgeV/C3BWfoktVs52PBOs84xRBYqr4nMhv8vxwPiea
lnH5MXLs6u4ZNhQJjxfG4Fap6hqOJWGTlgM3C2YFFCwC02eiqD98TEDiqnYF2EO5
MIcKa/eqS/8tLSGee/7beYTVtPP0x0Y8iXrEk0Yq3EDDt5G+/tzBy+n6fHB7PUE/
tDkvqAYSy6vuu+CD6gJlVkB8oX8uRxgVQkyYELbA2FPtNNE+1vg2Vvp16gN/2Pre
ivKuzYQSyYJNSdFfCKkhgD2f+J+TcyoVJ4wbjNdThOaw3ZeCJbkWYxyK5DY/nbeu
49pA4AhmghiDFOZoVxuPhCBw/QEwFj8rwJ5EX3tRpWfO/8OgkqwRY2nrmLermnu9
3GGilzxnagiPKyZ7hxYUFUVhQ+YWqSXMQ9PvCL82UFc6zxatuaPoCdJSrw3lifs0
PsKtoi4yOevv1vLyJEG6BB7+mZsDeJn39mPSXMesdtjNMv3BlHiWUmK1h0Ttzsi8
uNrFBSLCOlVqFiM7q5LozvnHGLYMe40QKJvPBuvvOqSon8/q48GhmKP9pFbC/a7T
NRlmaCrarOECRNgAGNXzsFhJ1SXOJCFjw+NekmEa1dO9aLZCdlsdfAd3c1CZgV/Y
ZYQKSo9eQCGYROFKmGocmKSPK88hwOcTgkdNixAh1ARo8HJtDpEVf8HuZs6zqLmi
QbjFBObwwQutFeurFXNQ1yX1b/gnyRDXwkt08fz4CWIGsIKBBP8swKgusqEyO8bq
DPHuLd52aoSTcFZwBFq4hNvMc0rOm7oqU7gQVS6oaphzUMq9RWcuiQnCrjdlAPQK
FhV5BF9DTb5G89sE9zCY3kJ26cRI21LUUZOYhc5MauVUc5lBnzF0BGbbkUc4Yhy+
ZtddzNm3qDCLGFoJV5wkz9p7K09Bg5OMh38Dd6SJVCMkFzHa8FBPH4QWpepNauZs
uWdK5T+qysFCl1hxoyaFWv7NfTgZ8SVo1L7TuZbLGCv4OU/ryhxlwwYbZpz7F10x
rzFh30Tfw/E9CYT6/r7pVkZNnt5KY26lX9HOSaYehSA4nRlpKAy4GrvKBg/LFHcK
JiAkP3+VeCSKp1wLglVYexS8z3VPY59AAki7qXn/AfhxcJW/YjqjmZjJmSG71Chm
l8rM/0o7nG+gf4ey2hLDrk4cNYKeiHZpKFUxRRTcLWaoDGMm0FUL1H0nxQUukPhs
l7EusgMLT0aqpbrzyr17zcInOboFBmYKssFVlBILpqLeNflffV85mH6W8bbhFJiU
jR4KIEACTT6XEa5+Oly9zZQY08X5Qf+16NzG2Gia65f8arDvOHCSxGlA/0Bzuqn2
USRK+2UfiALrjC1ZEbBBTSh1AxZL8S6wizZw37PWVw9d81QB2LxYvslo2Q8w/c3Q
W5Rtv6c1tiS4meegX1dmc9IeK+EqHD0XXbU+8NSz79J1a5p2PXvWCj0DmGLndzjO
4ytLHnDK4295YdYmhHCn+0Ft3IRfcn7UQYZxjcTimISwRPCqxSfvuHsU7M027vGC
qJqUYdWEZkOtnhPkUOaRgKRu59gEpJSF2/gaNVFbpfW5E/4lu6Kl2dh1uDDhFWN/
0QfTFXkrvdOhyu2nkvQ2YyRV+M0qAN+B7On5zv0qpOvR/waYJFJRpoURCkcB4ysU
F9m84dSwqbfSJbbrVrKk2xVRAyGy5WVHDBZYSacEZTRDFa5bfbCaXL+Xq1sh0/2c
rh3moc3FuCZ07imTkfJSRNof8vdxauneo2fAnWCVWaM+p2eq/NBQoIdTKLX0hYVp
R1Z3MvQyKMqJ0nvQSIHS5Gwfb4m0y2GWOqY3/n0WZDhydLzEiWK72nxAkyENvf+3
ANgM24kKFm2dUPpJc6ecIEgv579RxfHZ7INMVQpecnNRiTjeM/OW9rUdaLh6C+4r
/w9qxUmAD+YVKZEJAUT9kC9K1Q8Az2S3RyybmkNj7JI+3WX6/5aQkXl4ARftkzNQ
OIuMhVIzsiQB1uHLIi3vGNzhh/PPrLDt96QjjfRWHxKjik2KMhPwpzroS1O9x4qt
tBo14RNmNo72dDfGaKHbfCuam76HkxDEY6ZR6YaHH+2VLJO2/hFfjNykq6f/GOEP
Bv/u/BFDAgplE8rLOJykYLLGJPQIrbJS5dpLGOV2A8vTs4IuZ9vbw3lXW3ouguKh
KovnMYa+c+1xqXFh4MWC3376GgfOqpmSQhceSLbyQ3eXFWQTQ3Yv+7GpEc/gOAaq
Axq1y8vZ3SeJVt2AOY35IibqjC8MS1L7n7qBU2+0cRgPp4pOFeugzw3ROSlFJddO
eZ4O4l+F/sWA1HhlwD+2/l723nNNBUR/kOKhW5NhqVtJfzMSxo37YJcb51AUlD7F
0VexyHAyoZU7ErHxZ8FembOQ+KdZyEdDT5LTLp/VwAus8xWCczMbiyC/HY+z/9My
VuDJqAVhSEuhpiMaWksObMDBQqMCykckSMMvpaqdabN7Xi53T0EDgEiDxfr3e5+d
L5yVXVHw9MKjgnqrAvpUT70WV2LTQXv4jC9z79z6pxNMS6C7d1WUykn8oQkfNHiw
L3uR10/dUr8M7vqAHNy3hUEkavIy+xZAQRFnP9aJwUMhtNl/8CEScNZZ0JSR/wlr
+rPEjV9e2PLix364Kit2M+Q4ZhInDB57QBxKt2NutiF2KlnsDwxz7c3VKCf6K0u6
E+Zp1mMHvLK/WRhO1fe42e55rQTWWJVPa3UO51+FFrdS9CYZXS0MWvaR9uk2eYF9
7LVTw9iW5uHUWngCr0JNmDBgzPLM2MgYgI947AnnsubBzKY+U0Nhhhx3I4ENimGs
/RBT/Ycc3Zm5pDLHlyYQFnLB0erBVoFmmo42CvhORVZdwtL5ys688bpqP6+htoKm
B5JCjSRMrkM+FRXWEUiieYX4V9fzS1xDp+y18xfAukTUQ7L110rdNXA+dR89iP4r
lhIhRMo78rvFDlsKBn2pEkhsTVVaWAbI8Av+LsA+l3+8Yp+eboz5k9cVQl/j076a
EYh0868+xQmYAy+1zFDrgMGK8gKPHWytc3K0Js9lKCClFHOVM0ynkdSJcxmloEEo
Y37J0NDjjo9MKQdGEIisA7/+72CsZL2bJQTLfoHOjUIzoqNDQ2jI4rgjCOn6/jj7
igRvuLMupQE12kqrcaZZvG7wz8cDUrGyvYAetI0Z/a//zQj38n0wauozPw4ZpLCo
Abg89vgs5wzWQkYS4mQsatMcYy3ulwE1HpuaFvlVJANZznQiNUCrp7/lFjwPxjoT
I08S61KScJjDxakV6vH24UYRZl4N9xCwDx4Yza+vB4q0teYMLYj+vmiwG+XIv31H
SRRAf5sVHfH/2z/zvZfKpeCo2Qpo7eLL+WwSlW73Tn0bxZlXwayqwlTHTgWPakLc
TlgLJye6dHC2ZpFYw46F/LA7BvNtZ17Lw7mE4XKVkDM3jfKILMs8+M8anLi1si7T
cf1/Ur09i3VAZe7VHFUpAQm/pwegbGXvF5toHSLNSanTFuMnBtWicL+TkgmctNfv
oEVdHb35EHHkRGfjMtLwbBYAFOPSUSo9LUuk+muX3iEtZs6SxBza5p2yeheU8a04
EbNW7bRtmgiMGbxiareRc/iCOnb96GWQRpNvjOha0yxrFEKrQdbKuIiToKbHAYgq
ts4nctRh0d7bEONiE3FGVxR0DMmI1T9uPMlVgWIKgJAzSkVEhpb/1s+dnjggklvf
gkSCsE5oIcbk5e+HfXIf7u029KRGlB9Qe0AyojGhKG2i3wvJOUaLYtmD0+tDVtCx
ArRTWbZTe5AfonoULe+AZSr1E/FhO9BBIEjigZSRD6haBbdN1KwGwkDoHMVyV17z
lMdyHv8PTR/VB7IQzcH5KR9LwJwODkohXpkpoVQgEH7QfAkHxXHfJRQCD2lnGMzD
kq9BclYhzjliPmAOjjUqhbmTfZ80OwK7J6Z+rzLtjbIPdnkificlmz1Bvbc+D8a/
zm1y8vxFYWaRPvgT1NM14WTgoqwf9edavOgU7RTkAUQRwzqwKh4g03caicEY8L9L
K/U9J/OWwDKy4qWZMiANKKSDoO6cPg8veANG8y9X6yPY2yHt4Xx+q17eep69v6nG
b8HgGZbfDg1SvcPAZZ0p7NkCaQvteEp2RYiKqvIQ4I9wSyuX2iCWV7G/R/UPovHH
Ifbip/rytyZz8Y1BQFlG7nY7LLgHC353WNuO22009870OI3SXlkf1jIvyA1n28sV
SjixvnxpU0M2nXndMbsfsG7NGmKEgG7MsGTKh5QVcK7nur14CL6wUA+ZTlZOL4tD
0WjPbVU4SNOcmYd9DB1isemXA+wIvqnt4OQayRwZJgkgoDcOF509SCxTEvgVm9tw
zmMMg1RMw3TeAieeTV2Z5N2/eVxLSzzyDEBhYY7uWXx4wjGAfgw/AoXjJeWket/Y
5UbNA+0N8aFjeIkB7rgE4ZhgDEgNaMLrFYWG6v99X4dPN70x5/v/w715Rk0np6rw
L5h1mrmjbYOajSN30y9Pykzc3ALG0bSQR9XJIdpz3AQeyqZHgta+4bv0km101S7O
6XlBWlTvxDEVYkR6qMBhv07nI8tz7t9NUmsgpCy+Ko3Xbg5roLYdHVCkwsRzc0Kq
jNxithgRwZR9YBkzNZcAjVhflvV/7c+ThjC4d5GXuwnMGoItCmCxH5PnZsN/JYJo
3whj9k+4OsR/pFo8FHY5ppvskXAslTPPhPEymnsz7CAGTFNoYvWDKW3IrjJsjYVu
b9nwcV4wfxuk6W7lwW9f5KAmNwR2sq98dSG52i4dZVk3qnBdvzPRZBtcPE7iPVlF
tXvZ8wNlp+lM0Fdtl0+RdVc8efO3kSY9EzfLY7UBS/d+Gtek1HChTdEbe31tvq6Q
185vjgVgWf7DrsXFlWiK0i1N+EUDYXd43+gNfMwhywGf7c9Q6YGFsCaHboBLIuLU
HOAqMHnmVqD4m6qD2s1ui7aIhxz7GaggHAr1XpcYF4Dv3fqYrRTCY/AlCaRhzf9k
oTUZTW1G7nUlRiJS/mquG319DODA1MgQ+xQESEdrGqPWAEb4bVuwSGrDmfPsOyf/
IC0/8NLx6G0jy97/kPfZgxVGJBYnlI4aLaCnsBshwVX0esOdtYOMVLDkqNuJhLJk
agH/RSmGb3VNoUxTN/tesTCH5lzMPosF1N9LXrb9/hTXD8Ob7xiZsl39pgQRPW5B
fSDWCiYl38h7a4vJjxULXnF3MWggGVrAikyUyXN1DUBwy9ojuNWuqdP/gAjglFxc
Qsor7h0iRhgoK4q1l2JJPtQWe/I7jN3nJwWesre9s5ww3jp9C4YQEtexp/5wmeCb
XdFKgTkMi5OixP40p1TMppubpm2nwYpwLPtJX2Ak91VxkDFlxfHRsNjkTBEP5Scb
N2ZkDdhM2anPqsiNaxAyblg6KzEkSu0adwAzVVMXC9sntSjgivgyvGJiiZOMUrKe
0kKBRMkwXu9RroAyBr9mIk9JhazZutc8iYzqJuPL73LYXU/C1r8YxIUrKsEWDeo9
1fr/ujrCyWsZwsxiis1x6t3uXpdSS9l1mUS2xkXx+jS55a102yy3MUPXNCE9L3Xr
130zvQ4II193RpHR2HTEbxhGhzIuodG3WUPk1fek8Wl9W+N/rXUguQljX2P1Ww+I
G7JboSuaTsxeaIktCNP0dIaL9eop4qi+cn5bd4uJo1hhktS4VecGSc6o1pgrkzfh
qyn+x56cuFPVZrDgZMFXZ9IQTp8PT2qwLH5e3pneWHXFlMttMJAxujAMvXCVrsNk
aujNcZJQEKsVbV9/uCIrV5fhkDiaZvTdxjr/tUXw+2sRfWrnEH8kNKwh7D2PYMYB
Ei08UkxjPCLDJOHoAiGdhGumMqjyotOT5v46HAVWd62bFp6PHQ06RYu/aH4fqTLC
q4QvgZo/yi4RyKpUwX667//93dC8i2KjcZZG6oMEgzSMe5ql5vmaz6+lBHKIv7o/
QWkOiAAHgpKVsZV3op1c1JCZ3R0ZKsaMT8MgAKycQynnV3F1a6zPRXkMApuOOD3K
ZRvDxlxJoFypGTMvRHfR3rG56p1IrleApPCkbdM+sG8atdOPx9IOeIrRIPbMM1X6
WRRMTNa8X9z/rgSrB+J2d7hCuOfW9hF/wC2vUb+OTUMLL6APW+eNZQuOII1jB3ge
hEG3mWHjni6h/xQDzFeK7CKlzgEFBpqsodgwBLNDFmysj3RPqPjK+D8BfoUTlW68
sMYIAtCgtLhZT4mX3uxz1k+vVrRbINhE/8JAEH8q5ikY3p6+R3YcsGHFm+IjCYv7
WeAYfKka47iN5Z9DjR4ztxWa2oJtCuQIKkrFjhiPHbJvRjJz7dST+hvKvZc3hID3
aXQVEZzol0LPxTwHEBnnAND7Xe2UciXuDplxzb5eSN4tQfNZjKcoFMfhsUoSTvHy
afrHPWMN4+90oTnPKo7X0l9UOl+msEvrrMnVXvEDp1UPVTzgzxvNBMEtFZeVflLG
zPAWL6Mgs/7xvQQ3TavSYWWbfwPewNbDpEn6p0dUdCr6NBcJ7E9M26e7ELJakKH2
sJo7eFtm9Ge0wae5phHvSSFdnXXRUdv3xh8CnYVrWzOWKaHUjvkYsnTVy7eIRGv8
JI1ne712DLxc3ezN7B4sQRf5gCkghFSBBQxz1VQz+AZ+WyLPkTYmGXgwvS+/BeEw
cnSwkjSOl2xuDJw3/VNnL5Dp9qzBZjjzXYOK7i+pIJQQZwnvSkNT1LRTxZ+18bYL
u8hM/3N+5Xq8uf5ZedCutLUd69SioyMyxLuZ4xtVwsF5lPboEbjrTGkvZ1YKxFVz
tIP8UMKuXv51MY8/jQEkaIaHu1bC5dHjUMkgMkr8YSsP6Jkv4+yNJaxGByJVGooc
ebRI5IbOMhGMtD9viP78x/U7js0UGLLxSGJZeHHLQ5VEZbnUUgalA89zh2t3pPSG
nSw6fJJ+HPgLjl0rAM7Ymq25qEv1sm6THvBqpfM8GAFFDkaWCQD+hpdtqiFC/IGt
rysMJFbt4q8sFMMl1ZUWCUXBWSbNHtuF58Eai1RbcVF4u9l4m9cku0gs1eOHRTyS
1LxcP4h+41pVWAzhA3fhU6CVNthQNHTTyZhQr/daLJCeAEA0WihwIgjqLQz4ah3R
+rupMvK9u4fQWCUncatLy/3exDQZGm/+OQOGUj+/R5f7nQi6OTlBqozUUKp2V0sf
WAeXAYk+d93ldluEkdf9V7T3oad/3GT1E6T+lr1q2OGoaQr235qn7JjUKaGFiXdB
u5thkj4TV3khwypLQeXYNpyne8BxDfwcaHmNk46MzlsBaRw8HlZFhUYQSrv7EC/L
0Ub0r01CxMmrKjvCHM3fkoXtI3ezkKh8SVSC22soRQkhE9M+cJoYo+HmQ9Xe+keK
OYWbbyEP/Q4WR4Tv4cotpVXofAQS4SGqrun6j7X2apUJdWSGew2s0b7pSOgx9fRF
l10aobTcrhOX+2RB8yvcLo+YsNZVRyU48C4MPlULbq/tO8HSWV5GHtGfSTrRGRAC
8yuWMTQG38lyqeS/AUQn3Z6yj/WHpIZa+BCQK6dci1/i3wR+SHEfT0ouEcp2jOfP
vCT2Dlv2iIxthE1FU9Gri5eOjyk0S4F09QCIQjr9sN4aOANLqHSK28ZlaWfmoglx
YC0p3556Mw2i53NmAzlwCmt+oh/3f4xUenofb8aS/3BvmIVAGqebaEsWHsJQLWqg
P1RAoFl3498fS1dSTAt7UlIJZasighDM7Vcx4wpFSLW6xRWA7gwZhlDqsux4DQPU
+t89+8ozHiWH+kAA0AlyCyuK2aa8KdQjOe8/RfP+d3OS6AnW0NbmSqdgWmG6lX2H
8OSvCuqaDt97nJ38ZkypKG3f7pmR8aHSLc49T4jAphZ8f/BTTSAxw2tJuwcZXk6h
pkSLmd8lV7/5z/zZHyD5p+G7f1VzBsCSJRHaMgTJDdKtak49TF5XOOD9uluuWGOp
O0WpRajMAjMdWMXurqif5Mnq5I7fNyerNgwgLVSfuLCyFTXyqwKJ7U/TVdvYhStr
vYPtpjeYL/1vhwb5cBa4aKtoNcf3RbBXe0NhbOiYonW+kI1QMXBOSZZ4g8uqU1Oj
0zO46a8fEIrUFVPkRgDdeMWo+zKx76YwzLgglJJ55tzC+N/ZQlq4EMKbnBRX2FxR
IIVNPHZIHEPu9zCmsXE0cLFogY5BKcG2Gc/pKEDkRDQvB4wa+Iyj1gDTCrr1IkSh
bvI1WUowdoWOA/4n9hJhEYLe19G4kk9pi90lnCZz8kAB80ITaEwT3EL1p7KMdT+Q
uD0jjRHBgtsLRrVShxO2F+6JE9VdBapQK2G8aY9ihSIl+30mpXEGashLRUMoRgDL
YlO6IlFf3qlv28XAiCdHJ3CjsC5O56kVGag4ao1laRRw/bP/sH4N6la/1mhxqNOd
oaxW5mX+u3KqazS9wZGycCryNDRHzDhG7rhaL6dZojgcrxwxUp1Lo/cEL/lziHt2
3dC0JtaPEktm0v32hAvZII4tm9QW3pMfVbCiiUe+m/PVbz/WtzWamvESAkTvjuy6
ySnf1vE9rv2nGSRUOQLhJ1R5R0Nqga/yRbPGasrxOMCwiKwpR1mdywyicb6OvUIo
xfEQXu8i2ZM25wxytKr33rADgEdi98wtzOOADxi03qwvLp6MkWBBdGaabSMdYqFG
2AxFaug5KNksaFCopy5mqls63ysvirMHp4MQHtk6RfNKyc27eFOVeaAYgeKs4e5t
wqrgSBi2X/BTen62iZ/226tkZXjjlRyC3a/nEWrOluRzI05axv9ekLMrbxEwmmCn
6Pn8PZNLECrZat2ho7r3u25qAp2CzXg3CWJk5pMwQZLNLwUdXA1gZBr21Tp0jMjK
gRQMb+V/OGMhg0X3aphyExy/fT/UlvkEB42JNsJ8zy8kZbLJ44yLL3n2KxKIYQ8g
209PYrZYVisGuVK/JyZPYmkRzZkI8tvZRIi/pJysZbRfz+dInP8BNjz3GBVK/kcI
sp+pgeotbzXT5/4c53xDtIHuBZQl90Xi5eGN1n5gLjDZlsjfMJYyWQjvoeqMq5Ql
QPVtWatTR+8VukJ0xEqGmNwq8VyADaZYw0GdTNpaPaa19A5HVwl08dvFjJNfH3jz
B0Ab8Q1o9rkL4btYhLQRlEnWcmfzNdCpZqZF/JtYfl7PZiL0EiWtpnxog49vKQco
6xBOlJhemkN7zdNB8nOoZBR+bGddH5tA3bJmDY0uL1hXf3F+gGAcSbah6hnZSa0/
JYkyTJJM5yckYrjea6MVE21z5WJmzFwxQCWR/RdEp+AgR9SXlJEFZ4I8jOxWG6Tq
fcAJGHQh8mbNxMuQQNe8mnnUbZ5AK3LFkSJUCYEXCoYpCxA34sIL/9nLV8OSdwdz
893bE+maPdvi8AylEz2CFYgBoAeI7VsmVZHp6LgD59kC9P1Q/I2n/cr/a+gkNkuu
ZxR6XAh28Ol0v+Onz30+Cn5Gw4P3rLO2c+D+Em9uEShHjYFjVo80qiLqGZWH/9Bp
I3dJ3EW4pp5W9z+xtdz25TVyoiKi9dkhMs9tqU9fU7fCIyul+gMKmHVnkEnt3S9s
HwCWPpUQvCH49P9ooH+/ZJWNlpO7z7od/b9HezXkwG/50LUaaxX7Tn4tNv0nLzXd
B05CQ6gB++4P9FZiICiGDey68qvrTPqQlINYmjuKseBzrMyWnd/EjN72/X6mUPz6
TlN2qCaLvIqzR2Pk9Gccytwz2lwpyNwgvNH/w9aaLaNf6D9iXemYkj01h+MB07Gd
cmdPl4qim7oBSnpu0/wXsa3KO1r7pcPBD3wtuYZUQaMqU2AXPIecxGbrzP6Ts2R9
3LIJYkYGV4vXIzwWVM1MDNmRM2wcUA9DkrfG5qkyQ5n62p5r8DinIEj+uVACpmAq
H0Mm/XXdFaJKanfwBCHmjbdG5eepPlsaYDqiY7kHSDYAl1iQnRraW376k6Z1KPD/
EEOR0gFl9E5GOzlFVD4Ps7a397KgXTrRZlbwk07YmAqqcvI9p/KM8MqKr0sGz32M
7X5KqSovzDG0NGgThXi029m6WmhIBKHXKFLt821x9rT6QtsyloOq7dcwp+thsP4D
cGrj0SfKbNvEPNROX4D9lfAqtAPhVzznl2Q3s3tyQdE9DLxgrSfNqV1XTOHr9Ui9
XjRgsndgZr5GniNINRiZeaM4yM57zGxXhWUdla/HPNmj1VJ8LPPGwa9yXXNArcQl
hz4jAWO8IospEtdusQKnFe1fD1m3vU0YX8ffPGugV01lkYKYlU1JuAE5jqxHK8tM
Hf93YV9U60eKTFtXpXnkKWZgvRnRcTpZ5LiJy0/SX6s11U0DXSrSWNOrWgRR556Q
fQ9KW5zmagbP9MNQT/TbPr3Go/rMKJnKA0clLBedV+GL+mNt+iOMyWArocHNboRC
PObj2NR93pYP3jm2AMnVM4oN0DgFpZXVnEzXdW8+cDPP257J0KzSS926jJJkCAdR
O7ktMxktW5zTomwclfKo9ubYz9+fq8q+RqwnMoaPVZmWeSR0drGVlSK6x7c8Ou2q
WSkRqEixT3vrmOLJhmv+ZKalPIm7qdtkSWUXnSxkkJOJqBHqHOG5ink886haz7VE
wD3bicfFVdi2KryTl3pSrOsXorafWOYtG572UQ/bITtp6aHTThAl9qoGBMzbq1Yb
cxfPw4o+a+yk98JTOkT2xUGFl3t5FbFkmBIuePfOpOCA7x7h3Ko3D4bQOoo04nvo
ooPKREw1Y4LwnDBv1F/OLy2MaWMvV0Rs1le8KVtWNTjgXOoT6Jt4eGrHl2tptbp5
bMzVAsUZ0GnhqDIzCD8fHAWu3aZGBvAkExn4v12xSK7hHUb78AVLeMjsq+uBG8JY
T+mfFZOdEUbFpoigjFOCmKmTisDBCpQc+ObINJ+7I8L8mukLAMiegBXaroxO+iwd
htXjRZ9A0KA21SuLV9KG1tDKaLWsccpq6EVYBAm/IogrfDiBwucaxne7tPiybulq
u3JP2Af0D9GkfGKgmYTCdgBg3GZ9XPS4jqzbQ5yF99TnXuxKXilOeOjJU9XkW9Wd
lkULqAihQQD2aswTXEQ5g/knxnHyIG74wnjTj4wu/JNEKIM3BotWFSVfv2Dsojt5
S2VKsvQXwclnTvPm6KuDw8Xp8KVhzO6zibhd8JNMqi5icHpnPTMh+lu5xt4uZE6t
usnJ4z0AOWBvaBYNA8MO8+7ili2r3KPt9BodoWkm19o8Hnb1QbdEBTm60ss7j1Fs
kMeL4Np7geBllcueDtUVsKgyKkbuXNgOlo0V35OZQ4pTlZ6Rnj21m8ErbMaJdArJ
lR2oIRzekf5wOCFAnXwdZPhlzHJ1IKMZ18JXHUcFOzmefDwhKvq9bH7IUIRoM8Nu
g/djxB5s+9/l1C3LdWzubRb0VSwr8fLw+Sq0m+2VPIOrgAo4L7Sk/7bzcDT/ldgV
Iu7+MduCpqBxp5FsQrpMVcDZHOrw3Jv5JP7DY1M5wc3ruj0CrkwuWGxKoR9njQBT
xEpgNDSxTbM3pDJVa1DPdZ4T19n3hnu4DY7iiTqg60caYrHkY16gYfEA2u2TG8/Y
uADVJh3r1V1TDsiLm68WuK4ZhYN44mzoZpNC5Fb1Xm5XHoxEUFYVCJ8AHfqR1WtC
ulK3FErGkGUxcOpgow/ZzRxfHV5sWHJnpviqjAkzXRPWyF5CAiZaZuc8BdOSCcAX
7qVQ6pNtksx+Moz9U6tcZlSfwb9VrZWVZHQ93A2iUPtDPH5UWG5aZYmf+vbNO+5L
RbRoF0k+y+eeA9YArSBk0wKAuhfQe2fYqURzSwqnDst7ghEX9ZHqYdgWINch5I0B
/J71bRhB6ryFmoJKqlmKw0CnseNxC9BlW5l0LZh1FfjFxFB8xAE3jKplMKJiasTE
ToKMFWCt5Sl8uhF7FaU58xh1nCFPKYya8lNg9q1FYdtH9UKtrYKvEmLIwryggbTT
SKneeWXjt/tqzjdgPn7pjeHKWDDHCC/71SaqAOVaCpDvc3xtwF9olY4/BAQORNz3
XpFBLGlz1Wh5p/Fv5g5VhtK23GQ+b+ZLr+7IRfp5bHAigfC5ZdmqAv45fhGAPIoZ
xFP56Z84Iuubo911432zPxP+8plBuPCWVMw5Po+Xc+RhSLiFdnes/Lpse/11Pt+b
Q7sEpuMmNqnV9DcLwudX7LUBeutCLmoG/Xxc64Rq7scHCu2EnMU1NtSGYDAKv/FK
w4ZKgGWgOXyeaW3ayr0QsEQu64R2y/Zyxe3O6KFoDVOX/Q+cljFRL9Uy2Sw+nDhF
ePh9qrKf7aA276TJhpciU1LSCUIQD7Rjl1JfFYcgtNciD9yqkwfF++kt7dRxxVDg
bhc4NRP6jEceetNa77E84ifas/RB2D+dkc69BwZfOyxXJb34pnfAxicjzL6xgyHJ
rFKNcUvmrpXdQUqdaO+rRjjYXwyq9iNR87zBYlPUkzXUR9GLMzDCXseg0Xr6vutc
GrXqA8pjyXtNE8/np03hA/xAln4Dz2gFx3+DBogOW+NeKi1uwKUKmGyl12w1Zce2
9N+ikKyRvQaSZMiY7HaFU0cznu10KRAYR0e0cuzwzDXeJfSQ4EHqDDagRo9PTwao
mHxPWbNd6OISqHptVBef+kOTdBkpgn3aTAzmfHS98Lq6Y7RdF5qrXNlrqgy651vF
eM7G7DUyR14FZ3xcQrgm/2KYkbSIqvS5mXOnrhqPDrsuD3N3z/raQNxrAEo8Qfa3
qpLJdtEBSr+QF5ZVfLKvOpZlXAZF5h+qB07BfIkQq7otMdKEiw1uu+/BKHwhCTSm
QNoosK2Zo47AI0bLs0DjDybhFkjRaGP60RpGLMmMck0MBVdGrHBocTGd86xFZ0zC
Mp8OL3LVkXJmF/RAzC9f2tj2JTPR4kMQEtnbLcFTqpmnimUyZS1Tco8d8VGufluA
phZgDsLNxxF87O+DLdVQNNlLa9On62lrOKWgQspbfCNZ0UTnB7hOXXm7VnJyT4LC
JhCCb/TsbAeFizqZTMWZGWTLHa+ozjRMQP5bXJS0NiChybIjK6rbGFucseuJjLe0
m6X2ZREfhsiWuBjM1eA/hfJ+AoIfy9NN4m2KjQ/fc6+bpdK3GpS/1icViuWGxX87
gsUyYhadKjPOx1YSAIixglcSQmPzS4hm6xd539IWvztI6kv6ismQnf7Hs1s1aEtX
SdAJL7j7c1GP8zVynmLM3piYmIqzoL5U0Ne5lOFaUbjzDP28TlNQDDYJ2rcv0jAk
XXbTkynO+dK5RSB33PFlt1slxrFh+WgOseeI9GjMmYo1RiUwnwFJKKG7qNAlxBK5
KTw2a21nxYkjaDxz2wN5Bs/ZoDfbAmvQ//yB5q6CCKLkyjs2/QR+XG+VMyl0F3O7
F/J9kiQ2VfEaUCpxJw2+TLmuWCKqyMxeNDNIhbJY1WPELH49cyIxHhYoRHFf3mi8
njCT7NcF2tRjZoJu0eOCbLCKaHS1Ah+etBIO039ReGAw5qnH20KHxYUA8woMGRcA
QnutmlV+NuMtGH3Ho/hEzA3zd5aZCVa7GzdoE/Ye7malwTzmqkcdmv37WnarDJZc
3fdYRtKmX2prMPCyAeDojMaFwjlywJm8gEGiJ9/SGnB5kEz5/sTRm+AM8pJPYtGW
mRHLnZ+gSNVEv4TSD/SDdPtqCjHa3BpF7oSp5ncVNh0VVldQwj6BtFplvuQvdfpF
ntcwCz3uJWArMhZ4cTspBQcOJCvySHv6K+vocg1okHUBYXmM5s5Up0UX+n1UEjVS
aNIqnH1wOKpFZ4tp6GFZQo7hxOQ9EMbJi0KFWMQ14kH0++kLK2SwCn1QmnE8BCyo
p1gAsj4PZs5FCno6nvOwGq/JyRkvpQrJA7fF/W7qofgOXjeDPbEItEp+/jSfvwnf
om4zdOw7Xs/hTJ3CA9Rp0gwsp7tb1VDUH/Avr5VXR1zjIvf1yTYMP1OpKJH2S6NB
Uom/8nhKK0VDhd9t649GeIQg2tLXfZenV6whs7cufa2IJj6WarxI80mJ+SnAwONk
U6YTeUaUX77ecDezuo53YiaB83Bj+ryviQtQBioaw4fs+UvH4whMQYPcfUb3sMYa
M1KC5xBEAR0V7RXPN0OGtV3sfaiPXMISR0i8nQxXJsxHD32boOhB0pMT8kSCH3MS
Yf/uXtStDvAnzvqRElIFaEjHTQifRKjT9yaLXYgpBGdWooVJntB+AilnLKG1nYjW
Un9cUuQTEudlsFPrWqPCamjgkjzN7vXz0n2qM7gWtEE0A89d446r88nKTpkYdkJg
bqEiJwW0TvG6OQlB17eNwIQGBTULvV+yzUx0yFAG97UipDW5e1NSMPpl7pI0o+1H
dcIvFf6oAaj/DPyCjWztRApKZeS3S9O04TgIe1HA36TZwFB6D4m5RMu8aK2KjhGE
JLOGxpy33tKFcLNKXfSr86Z7v97/GJPHyG9BH6oS0oM9fN066ZIEIayO4QDWqYeE
dym3ZeWt/Fx5YCo7WFgniz7ZPHZBh24wn0J9XyMf+f1s3WBOXtN1iCDdoE0qQh+C
yQQCMfNjG8Fs4ce7YyCsfcFFfQwvuz3+ECpnhdYQKwYWx1HfiAUwD7ckFrM7R7zE
Ax5YrMaNMQGC8m9dBfl6OC+xBUOOJpSF8FSBLWkL5eCbq+15mNSeWkA4S7x354Eo
tgj7ybSbiz8azbnqDc/3Z5UgysVy0AC0eMbZ4JSlbL3Tk0dVFYghSMGrqzJpoyR5
Cq/GiW14sPC3XhH3gYJBNl+3uI5kPsbhyxjjFozgzDiYvz6c6XKF2SSwOWweGOXs
7U29BU3nxFq9s6OCa4tJZcqLTl0IVxDedISZarRJE8mvZj2AcyGbXx3+9gHP/n1z
NlGQTo89sMrDVsDPjSQLN5HEgeoAR9TFcaPSaymsbkQkoo3F/c9ZNqj+Qk46QirP
GZr0WBisADNOGdGpVbode91VDHuusf3E7GeMl2MfEOSAFR7+t3UsHOuOADJ5vGo8
2MTEE8RjAtR6VkiAyKJzyF9Jko5owyZipjH+juH4kTjLwVVJhOk8LBlTyNgq3Wgr
0TJHcmJhjV2IHH3wewJ5ZJtvnEBnhQ7CeGhEeuFIqwX2Lha9GcADbHJm94T+a+y2
FRsWK1PsA+v7BXcoo8BWkvBv+Qba2qqAtMk3EgJPwyIua8xm2aO7pvS6Br88zDIb
I0j+b6SzplWPXzTE8wxNwdY7f0CjH3Vr1ILZcHbVoihEJJIpsFu+Q6t88Hs0V0Sk
QKDTfhPV1tFu4nGW9WD2lygkuvh4yscBGcMXxl23InyQObY8p58nYd4b4By4gcKb
AJvasRp5ZtNArZT0c1RPpcw6DcXREb3BHPt2nIRe9/g1b7cZiiIHReolJjtz5m0u
LgZ+68KOwvcedTIUZquqZoRo7XPTsGOQ/pF8SYu3RqLnwU6ErWgzdSIty53Fk8CI
pj1cAwGFUyEUh8pCpETCPeIc3EO/F3gACJ0o1F14kqgFSiOJ00DlnVH94BZvFpeM
ImvSKxgTvb5ISMGwuUbd7fxPzmbcOVHw0qUjF8ZwHYq1bcp4DGnhjqLo0z9Av6dC
YikPJ7Sx4ccc6gA4AtqzUTubYXL2mj/HPyK6/dQZsNGyUotuQSKJZq64GwufKPIV
k5wy5jLSKoLF4DJqo5TrpEklNILvJ1JBU46iwDA1lrP0Tw4lmjt2p06fmBw0Joh3
khrkMNxc1abrIUTg0NusDaGPJbRL2FjJZxGfInArafi/ERc3Vls4HauivEtCmFeu
WHF1R0SFrssNGf/0z46dIZMqX1yGbVas92m6UGOdiBYsaHxbC5u85C16wkKkniZE
IE//WHR7WYR+PWtWrPabYD6qdeSUK6jteqWaP8PpNUwExl4x6PTcsZIwzeuQSrq4
QgDUofwXDzrBpqKg4obVYWmQSoeKJwkqmh5n2QW/1/wXZi7nASzG2fE0GxBr61mS
BUBRNLBF8qph61p04EWWZiNNgjL0X060An6giZ8rYTZapou7KYj28Mo1A2Qz4S7r
82Zxtpjfv8dfzF+C/FPhy1ttoz5s5P/2ENgtcFXtNBnCWuxOtXKhTUdwVRa1zq7U
N2e26uOu19J6g8KwwnxcJQW0R5Y3GT0t5csb6wpD5TMh22Kh9TsXdmN98za29q7Y
JFJcBGyynohWxucgt8LPwtde3lWQutgAax85p3pAON/GPUGFu8zcZtYkPljhapFM
YxwBpXXGR2ShpHnRvaxlggbsTDr9ZuVfznYpJdLQFUvmOXzupQSRTv+O3th00jRs
BrhkRvb73tn6OhzkZiFNl9/AR07C9AxXa98dkdx3Me5CZen6eCwSF3iy6mc/lvxe
1oNApWJzYJj6LDrZb/sMzETxigJ7qwzJl6Dr+Y9yuWqnqVXJrGB72bb5Vr29o2l9
F1DAZb2yIKtKfrNNtENbuM7R8h8eKLcps47jP45u+MRRkSV+6A7twAtb8XerByq7
LQW3l7E2LHMcFCwYBnRuC5fH67D3f0fFkVoWs5BdVtGwgG1cbnD8hNV+ZHY1JD0G
MjJajgQ1WWZBr7BXvbAna4d00BvtOPXbq3l+CyAjuMVnlx3BVLBxkVbUKpHUPhII
I46/9J+VU/qOWburn+tJAuUUpCo35+pqIskEELAky5puiqL7LVf7XfBOsNhhPlCN
c/1y+jR7iQAAAPWSpAxUlkY5vUa7kosBp14ZlBFTQlig9VOUAXqgFPYReUQq2vYc
1rkdmr6W0mFd1MfxtXXnWLVssPfvpmSmGxZs0nBQoYlujac8lx9WGx1naA4WkdXh
NXQkDxXUQgi9S5Vv8A0hFkQdRJXBSrnpucc9+HUhWbyi1WSVifI0D8TIfWG8z4k8
2rfcS9Xh4p62zdwZAU1fbLJRTIby2cmbBpxzSgFPyxX5quWswp4y/dXLlV6Yq4HO
WanUF4qq+5UeTDE4eBMED0hugdSj6SyktgB/CKozkc8TkuBnQecGg0mMFPoEHe2+
V2doprtEGo8Qeawyi8VMgNUd13xafOopufscPrAhOjBhljdfTNNXdaQOLa/4x095
4ohJbsfKlKOHc2cOOjN14Fs6/bjk0KNgX0qulBWX7wUTPB390RsQVRIpvRoVSzle
1dGwQE36KOijTh0oPSy8DNlT0ekOAC6kjbhRPlUbzgl8msibW4JO0WAU/+NTncUQ
lEdlj+to2hoPWUnn1DK7d/R8bLyZxyK1X8Pv02QYIhya31MW+FBZ9rTIPlWczpYz
LUX6YDJIPg36dOQVjvKfBNxuZlSUJ2xwVnhI8PvQqsNqSo+VUHl41oDnGDtDDAYb
U3Kny59DBBC7KbTp21jIL3o5domFJ1DmyOVvsrIuz7pUWUGVH/LIeePI0HHQHiDF
Z/zAOT+G9NYVZ2oef9kq9uVrjPLzGuhtBf69JOgF/JDcI75T/PNXCX6jq1u51Pho
GGFiQsIhl17ggnkBrUprUmTCp80jhEJz9k1H571xf38nu22C1cSDOzEQw275ZRnN
61qMpji5ohan68RMW94DeA+q1VJJ6n1UN4pQH1x2odLKErcnQfmb8PtejYLOJJKq
jrL7UW58IJ2tjvJPIoU1jmYwxkC5JhEHcx1JiA2WAI/XAaIWhP8KMJ/TlFzgWezN
1IALO9RIX/1maZdxrIOrrtL7ZK4bbLkLqObjlJLeMz9irPqjJd9m3HjZtr3D2D2E
3NSv4yj6HCfzQyHRY7WM6YKbg2y3VEa9mRshRNmcM4pgr9CmG8SRg2Mx3vBz8bgi
hiFpUucACaz1Bz4j+ukDS/ppcmsDAjKIjYqfOFPGe576WRNyNi90o96keApKE+Mh
krMAKsjkjZx4CmOpXEvgpI6wmlO9JSHXv34K44FpozfTxY1F3DSyI/RkQo2DqiMO
55AwcuGNIeyRC4WBkS/IPJxUSMCdDjCtVc//TKWZgcyovGKPdWJ7Edt2tmBujkrn
OoBBmbCLdanlYUwlr1VI8zecvH0vwHrL0YDDo67Vt/dlqMVGqNEn2UnXFdroGS5f
IzcQYJ32GyDg0Rf6kDQlp1FCLQshiFPhuc+wh6R/CIuNYgl4Z5S/3QQw//wbJwUR
6cNxUikTc/4VmtxxDSb54OSf4vlxUMYkdi1bPrw0OMBsOghMrESlcohDYMOZq2HV
d/wzaCa0ZIBLimFw4Pmt5nX+I/iY4Hap/idj2j/4cDtF6slyS4onPeQ6hjJokoH7
CjFNbxbsb1qaU/NYfcDgT1Z5xaJBiiF7kHEo3+so3SgEdz/ESecbnhfBJXO7qNgG
PEu2Udi37orEZYFCIXUzKulwCNkiyCOinTtzxScsUZtTXEDr4068GYKVaVeA+eY2
Z0RD8up+rtTxDJI9hr9g3jS+2Kre5JS1/nyZ3q55jujz0hjk2zsZvaFyfOrkmh6K
GMk6nV2L3IlfYUg6Gm/Q8X11aaZStcIWNoy8Ct03/F5g6I4B8TkZChBXkmilxTp+
5O3zPh6KnEwiajR2XEhUY9gVEpnKG7c6ViMmEqJwLl3YBg1CwkH6BAJ/nN11sHCn
NJNkb2RZyW/25sd8sN8zm5FefMTwwwIUTHmxc22XKoWIi3v1Ay3PzyolJnbB+3Cl
pW1XcDUfR1m+tvfFzlG850QdIAtQdQxBMdN6m9xB50Chq82FWkHXN2oC0cXJLlnd
Tb2V0s6gFXoVW1e+dlDBPVqj8zp8/6wkjFRq2jli21t4thnNQzbZWq2li5+5rLXR
MAqHgQuB+T+CbqtwxhqyZK3Svu3TwqlWX4dgnfnsx2NPr8cQCOOi6BD8zbnXP0RE
OA+P4FT/7esxr8LVZWWOpa1/aHG685I4ElErP4AJrqpQHm9LpAopXnqLOgWrNE1w
Omnxz5e1rrig/KZllQZVooMAHCHjuzARioWlDSE5ZG7uJ8fdK/QkXiduwYmmsvuk
8fm4AegqPH3606XOb45mrTsyDzy0fat3fYTqw9k+iGprHvK+ul0oUOmnhl1RNkpm
OJLJ5Bu6iPAZ/zzfm5/Lx1xtullnuMwKmZ3jEKoTUHb3oXZZwlXILElZ4iKA7SqJ
rZcxLpCZUdCQdTEQVnYPcJdIHkR/7Lbopi05ir3jGNsuI3BnrdbUeqyWbOnjo7mZ
+1kQA7PdASEjrCwM+poKm9eKvXUTnVbPOviNxFiJq8vPQ1NEuvPJN9RDFWijvJtt
7365wxyKI1DtvNRXDpmb5/pd9jU9iRFZBiqP3QeHDXroQDDxbCOD17vu3XfS+ZTz
/xUSMXfKsfX2K1/+Q6zegUl8Jj6zcnp09CoJZC78l55FkapOHhjQcA54syWYI7R6
XzQWZZ196ukZHC9/lEnayqiAtpse3WMpt9Yeyc7CLyby7j4DWB9qmEfybQwBUZJh
EXBm33a2SroHKQrDg6656ljOpgvETshkHH9XEU3jVvYofOKL1EUyzmm3Vh0fYG3C
Vw/AeH4rnyioCU1boj74F57JqQWTyvvv1FkXcsljN2DfiGhXNY74xjLHRPXFaVzC
AnRMCMEDtxfIBw/X9dq5A03VTdzh0ndEgfRhdihBMNm3owlTMd33qkKKwVGO1gvw
XFNGVIRMm7lYFkWAgIQ8CmonMWTo0/dtMiDsdfilsFFMlSDPjK1CFu4IzHMRw4xb
/NIiw4eUr2X+OApkdEhv7GE4gokU9dHW+AyMp6KZbTFYhtGC4kmpdcvNiSS/LRbO
UNN9zq5b/MM2WMxywlVSy4qGsBJKTy4TJRFJZWA58HBCJbyLjQ0muIvrw6P2ozrP
Apr8TmIhNUn+BTbxtQ1bOYposiiyZt9fWt+GGUJiYas/zkvHT+s4/O1OmT29Rems
VYYTkkqoPVRQS2U7fdgsVkCy5rZmlzh47sUJBdvl2bTIFWWOm2Fw/cgHrDxv8s+p
WxnYC0LiWDVNFRjobPD/koXsrc8P5pXW93VR8q72ec4SoNa9ncyYL00k6nUu6+es
9NGKqdNUlaX16+60hqwanskjOK2D0grYNhEttjYCgOkxWhO/cSeutAVcee4WnPcn
3v+CT6ttrNCgNFU1rFGujLYj6Tw/BN1N7TzMY1j+P8+iE7baSgG+LlX9GOtz8IwX
0AxbDpTH8+191Mkas/3EkY8cpXkY+u2iIU2wMpDHSAB8fRJn7JmTudnetMBA7uiu
O6hc4NZuuTN7cucfW/TCKu9HaO/LNNWX7l50QUSIUx1PSk7FcaQg1xZNzgVhOGuf
0zYLfy2rewmLKOVCFU7/dyi9DAbw2Rvl6ZZtuKks+lzrdDGHwskVzWSzIP6duEoR
Jqcn9vBK8rruE9gZPBE5vQDWUayN8p8JPF/YFB+320VMTp+kwkxgCH3514oxWKVR
Tf3PFYiRPhejQB92Hhn3FzbBNTdf8GryDRUfU65NIvmotm08hUKmGzTNCC7SjR0d
yFyXWMwNRnM+DoERYeqkghluJL9XethMXXXEMVECOgkE4GqZ6T91gCdOTyQolYmW
mcy/WPIpWNu6ZDtuMsM7Th0eQeyt4G2/RssOdE7Vf71e8zGpOr6w6NPUlAxRHBEQ
qERnitrCTFjl0NXbZapAciEaRDMG39534zQU05s3btjBjxyeLe/UGp4OA72gXAMl
XnLTi6XRncCVlr6PXUd2jQZCyOqJ4b0TL7ztbu4R+ugCG+wXQ10SCxE0o/m5mX2E
BVT8GgNWshx77sIeKYUwSJdDHHz7b009nCUt5KEB8o3sdiYn5oebhUffn96TztFl
DrgIf3N8i36C0DFyjhJibqgAd4iKVPcVVhYl5cSnKp3SmmnvtLKii0w7qFEcV4kV
vOk7mGjz/KtfhkvQixcp+CxFWnRdTB2xy0s/VT+2vN5DXPHPX1rbxNnefC1MFq81
uvXBarcqguDSYRrMjUMrHISBMZy9BfjvbV7jVniRLpYOhFUka25r70FH9pzAtMmR
ODGgOqjTOdnHRI25NDhzf41nvJB5DoMQZzEi6CoEl521RaLYXT78ai4b1oWDFJz0
R3OXFEjHNi9NHAgMwK9sYHKC4sBrTlCgmPVWve7lla44dWzn472rlYSN5MvG5awZ
bT8+W3ycVW89r0EKzE3UzPSmq01SZBBxsjOmeQDeBBsiYkR+NSNYvw3hs++pt8sq
6MsZriMk1AsmLYb0sGvSyTuw1JSUm05P3eIW+9meFu6Hr/y55aQiN/zlLoB+89LU
4/GtAwozItMu6gFJPoRZ7GuNfen6Pdf3PIrd9o2VIrDTiMfeNPoOk7PBlz71MqDj
oqWwU74x+tx3D8XVS5LfKEeM9+UwkZhdq58uTF9gPi7roJpixzIRV+EVKrOjt0vM
/n29AY15uQTFDLOj92fqWfFds/NFKGKGpPH7H7PDsYtCSUsut9lAowAyvZ3LUWqv
pEqnZjJALmouhuhkeBzFfOpfkwuLpyZnZDA6Y9CY4bxImCtquNpuwtgDz0JFr9zO
0NLeTdsOYYhVo+/hHdAoP2hBNNAlctMc6/JnIz03BuebBuiVnXqUgv6dfg0BZGs+
lHlCZ5JCEA1h1c4uYSxfv3OIe4JtDclIOG+NQenJdRFCLAN21HvJjW/5kXlaI/Kq
zAdt/v30Rx9dOKHHg0SSW4NivFd8STjjFNJo+Yl6zfnS9wDE0/n79/r8pJ1Oo/Kv
+3XITdCOXYERYiPBZevkZO/xF5JR0uWk5UcBOjEveqhvCgDI8sz2cvkWOKFz2nuH
HGTBxQvqvlnbXS8Ni3fD6dVY2du3LdsFe0Nm1udRTpEQ4DSCOfJDNjn8uMnRhLjq
Gzm7ZH5SBulXDJg8q8xTBq1NkqqWc07d+LztSjLXd9apJWc14DH69TEIWwtyz4jq
w3SCAUSlyCmoxwNzhVef9d4voVpEnUcNcDVAtpkOSCbMq0+21K/nQqfr6RW5ArPH
tnFe9JpJlkGBsFG7gFDZov0AfF9IRFXdJsZMn0eBEfziEXZ5LkT2N6hOplN09POu
CNdUeArsZ3+d7FQJOcCjbCrA8hRt9tB3jnMOpt4+hZTlpSRFPRP6PimYKMW0fu+y
5j2r3W5nCS9PRml3XfXb2wvUuzNc7x1Mo9AZt7nlyX3gjDxpjMeUiFbsU5VLJaol
PAkKl+AedkVlxEc4beWCXDw+84EVUuBL+psEdOs5s1yfkRKek52pNIWRdrRQKlRZ
iH0u8f2dlPeSs+R2bDJUTc7FWwkIn2J2pfKR4i1YmxKynI9p3Mc6hpPE/YkCFtEP
abpJa0PO4wwykb8ENXTDznaqSonQzClQN937+naCAmJ6UgOvFSajshHmt2L3jv9C
0ERAJCIngPINXliWor39UexHJjkXMuzwbZn+GpHQE13t0PFyFi5MvusO27iy93k7
RC0vq9Q0EgFFQMVNa54WIMPtmvVeWQVaLMXcHdh0BJHE0iTpv1E6i4fhX6pesX1s
q0qNDektnAgyZ15uwMeDPZDqyQua1TtgGjiIwb8YaywyO6RMfuXj+HZ5L8rug1jp
5x164StKai9JJ69FHaKdLG118FCx16xXzjNiDd9OWKrvaGa7jJR2wTTOoE0XvEZQ
fEK693JjYw08hWTjqq/CRADvsJ9th7FQuwKdVTjC2XSeS2yEIpOyg0yRF2s8A7Ac
vXnthp8ccWZzDcPFapc6wQcgyO39A4Yz68pqMdbPM71KT8gx0r7QDuLkprz9g6fg
11/jDZjvfmHRT4ntaW1iNw7rre5oZHaCcMQaF3wp15iyivwKWz/FWvjbHTR+A0xX
R2X6ZQYmFmwWn9Sq25Ykkb0RisdpmrdcfA7AH7AHg7fpIGeV+TSOB61GYi7mWAbX
mEvNUXCPE6YFLr6lKtq6ls4D0FB4zxW3TRBQmxXK6+IOuzU2FghEVzSMHrpQ4j99
KnIGjLdSprDCns0i5tgCii7fQrxccXVx/hs1O5U8xx9xmR9OtMUV7qCItypuB9aD
8pUX4PICpkSjResrG+lo8mvVZdeOqTet/LV3PQkIwt6fZXJWbgJq/Zf/c43kBFOj
c5LQlZo57q+vWpd4Qo6cYZGlrrx1UZiJ4c0GcpOVgh/X41+/pzsiPSOjqq1W7AFO
20c+oxGE9V4i1mrWkDOtKDtD9eEMkXkTKhe7o8iEvQwKO7Grgesrv65LY0OjhFAn
35OufsWg9BscF1zDgq49CwSYgagovk0py2PcHKIlR/VTclxmTQuI+sClV9URkOAM
4MwvOeqG4QpkI7qV7xhYCefUxNOkW+4bx1v7mo6VFNNVYR9JZacs6wF93IV9hV1+
ol9w/VYiiCttlVDHbVWLeC4nWHJezDCJAPGOGRiUAFbfzKHZZXmYZ9iBaTnOAkOQ
hFyXxyV1lrwBkrsX+2W4sTvRuWzjo9is8454zu6uVMh1juLi9jY8rO488FWCBb2W
mVVzKOMUgndn7eCZqj8u5Mrl04Yy2wmBx8nrZKMOwh2vZ8pQAt6SlFlHcuOiMa3G
1/4btjGp0Xa4r0w6EaBIpiIBFHfXTr+YBw5QexiE5O+Jv5N+NuofWcVQgKrh4bAg
2H1ymuJky8JR5/6AsSJR9lKYXQS7tw/119pj/SiTFEuiup7bUBGeH3V2XB3Q9EuC
gbGBH+Dyxl1eF1zliC4UPuEyXt/Dlx9LqHM55Iq64IrM5jen+tjaf2Drhy2tv48A
zyQpXkWxnQ3mZtj19MnFK7kvuA4OyfRQWb3lEOA9au5q+ZKfGPcS7d92lbY5EXIQ
rgCrmxxlE+zzCiKp82DsP9y9laA6zIw0UzoTL3H+wMEx9EDZNY+Ide4OiWBh+0t7
SdVptqCKGup/gjl233YYcPq0P8EnS4BvGCRNL8PXQA08rZ0SzbZI19zG5YWPZSGX
QNMQiV/lnNgS12Qv0f1vI5mIbw6EhIaPzpGaJQa6fVlkjKN13jlzePxj108R0Ser
cxmXPU7G9gkz3Rl9nc7sKoGlcDpSBZ9RsPNfvx0KZiuuiFrvjU510rQkdt0c3HY1
eT6hfqYLNS4eAXU7P2k0RGirt0GjV5UirArb6+YK2IxpuKcVJR29iGgm+oiNtM3A
hDJqpDavD6+su8Svtj/dAfkwvXXNZv2/u/SgJrSygl0odQP/QulIy+fTCnhgGvhd
p3sm6maLA9aDSTnV+d6ocPKIj11AKR8wNsXfRKIPV0rpZasYecEllvcBLbG0gdMZ
xnyTTsBdutvSMekPtICILj8/CeGk9l/jsm/hZBfYdrbVr6HMc94ly9PcwyXOMGNA
ndZxjbevCn4yUUaEYaDrM0Xqq44buBL6VnXQvhxDt6S7RtbNPALuL22Uu0Nn3PFx
6IHrNVtY/6gmtFOYoNgCoKKA0PDj5T2xUpuhPo2EHUAKUfc5ok8+yZW0Xx5Yfbze
932v1f5Mb52F/QrfcHdk0ETeC3uqYdyDeZdK7rj8BjRsZGES3XInhgUBuXt52E+p
sSgnUOLlE+9K9YjDAXUidipWE8c+UwO+N2+bbulP3Me/f/+9A882SRZloqSu8/jT
IYUf+K++y0bZ6bbCyKs6CctBVHKOocshIq9zIcBtpmy1w7PIDAnq2S3ObPZUt+lp
FCZw1pS8/PvSmPuEj4GESL1dc54IK78zNG4fP82GQZLwHIIev6q8NeeXzjv3pSLa
fo+jCTZkI8XbPSlALSU8E8WJ64d9X72f1m/bOMiqZalb7EYZR0nRzpGehfUE8Z2U
q0p0fK20Me+AKf2xjZFp1rBgSlTPVNrtRjBelyzlBSjn1aiJxSh++zxUEjcB6gdK
ozgOJFK2xBCn13b8atu7aWzT4JNpGk74gZPV1k6BJ8SaYpke5COY3MCdUce4l0c2
pJZ0CRJLMpUuIHf691wYIwhiQnqkOzWinu5/tBcqblqSGQwOjCCnP+KKPsvAtBxg
O3fRXwcGrR2O4eMcqofOGy7roUeWgI/SOzcczVy2PoWhq1khqXtL7pQRKTmPGHot
PHWro29zSSOxpcZBsDjoFTj+NfuxYP0q5yyyNRYjuZfFWts2trMcM2IHPB+kkgCO
l8wb/xYj4/yczkF7pS6Vjq1KK8TT5bYa813YC02v7mZg69LK5xrYGTRsftg3lsD1
VjqZpqRAlGJxiZW2CvJVU4exucutjmT/3dLcRkU1iNlYV5oWdkBkHBuK94fJZL7P
ZlJMePU5/cXBOUZolgYZzkGM9y+kaJJRGNAdSKuNBzWaCxwH94wNOdZJI1oHfc1U
6FMzHzBEYiA0n/XskRj7+XvD57XxmiKRS1goo9uy5EF+pIvudazxNKpsGYQrE+jf
zf+I2hlkTlElD+p6+JYP2rTpjQiNRKj+g2kE67mKGCBGldKnax4edioRHHVbgF36
Uye0nlWTUA4aES84WBii1qzcTMg2wNbxPUW9IGIsSPL82dwFvkYnNjIEsSqCvGmi
tsTGS/61gw2/sWiaURb4HfyVdqnP/x02QOKww2lqxhS1MgsBr/rsVM4kW8JRKcKU
aWL6HyNhHodzKl0moJVpQc2dzw3THm0pzyILlIYkD+IXvqifiPZVeAzqP6FA3DHS
+lzoh+ntDDYw65KsrUnmhhNw0zIrYHrsNoAY0dIDiFG9Skn89hmNzbpMHrpS0FaC
Zz8O8F2n/OORJuP25X37oclPSAkb/7K9zNxt88NUrXDHb89onfrJBhVkGaw2xIVP
wmUsKTpWfGQss8V1ul6JVHB9M0IPuZzwb3v6il9GyE0A7pCOwFYOGnMQMgDK4Jh9
YSHPEFDt/Eck34a3B6gmIM99T9ZqwHIl0BEWrXaz1109URv9dqD9CqXOJaO8GnX+
1WbIpQlFwBkRGurXaemtutBr4PquMVFDyoUYFmGrD0PxBUf++KQdifH5HW8a9uyz
S2yY2gHiOEZMfyWz8gUJJYd/apkPpxBNd/AL7wbCXdSlrp0XxBqWgS4pU5188RS5
npvhuEVnZ8XBc9NtHTtRZXTLsRcBfkZ2fRs/+qlywt0qum+2cZFxGvlf47HKPk67
DnN2K+ml3qDL8urWeusr3RuTFCyQaFWDCNm6rFKOsU4W0vV5J8xEPTq0e/Dzerqk
bvkffEgoWKhQxMwJpCfxJKaxjCkX2jMgkYfQc7IQpQz2COzmcakG2fLLeiTbywy9
BsGBtkyMmqfAxr6ji8Di72IrrV5MG7rbpoHa1XaK0piTSuiBvwJLXIeF4spXotI1
0p9E0+PCWZUvNyDywBC7eb/2NgMPJwDckTnmNXPFQoCgPK6rKQ8LNAYCd0z+Cpk5
/SZaYrAmz/J0cAAIAhVtUo224A3LMhIAkuAEO42ixWDuJ9B4aDWI2kCrUkq4qpd3
8V0PshhcRkmlya5PvQnBOak/tiFE17NDNwXl8B1bTXx67rGk1aAdzp/LVrVcpBy5
4eX5Q4eiwwiRgNqeLrxYVA0777DomcNUuHt0Z7Wv+P75ZG0gE8kMuErs/qdcpDbd
FUsjnKHMLmiM2yAAPBIHzV8qmxBEL/FEiHO2Ja2DCrnbMrY1HzJkUCWgyIbRH3XY
juoxWc1m4JISKxGyPBrr9RQFQ683hkKYHgKW1ubkyS65dKORBLGQkTiaVXawCGaf
m0p6m55+OkpJNAo4fjOOsbQDxdgyi0FvE2iMjLh0fiSVlxEcb/xZ1eyoq5Xd/wjb
uTmg7G3MFDvQiUCZFEx0H5QNTHk5sk17AKbguu37R9ejy+6esb8wF6uV1S7RFHFt
FsIY5cnfWHCG5w4yW21d8OocT+rv+TNcznuaNmAi8sca5f4FcjV3gaifx/k/MhM6
aTq2wLjvX/4fS6/S1nAUZz05p7GWha/ajE5HzaNxYha33q+NVobeurrOLKrsoGCl
Tgj5bXetGT86+p8u9ajJWbDRuS/cCGcN/LbzcG5JP3XvxhfVPMjhkTdE7CASuLBU
Q8evbcuLgIEnQLLS4KT34o/VkEKU3mear1Ie26k+sQF2UArK8NYsUPLCLLbM4hWC
ud0hLohGsQ1z9nz+VH70r8xOWiT/17AmqhsK/kr+9x6mBVgaBrU2m7DsqKvVkrt2
ZGAZyNy7rU78TmnszuIZFBKJ5kC+KYJ2ap5AisAp6g3IW9pVMxcDB/gjDgTnZ0NH
W4NiJX2E2qrNF9err8LDraGf/a11BWOMsnHiUJ+nfhgA2EXZLvZHgdp3usjIJ2Uz
kyAGGhuBgsB2upofLhAth3jahUz7ozqLeWdAEEzwwzFpZUOIKm+5AQ8sw1U88/AK
vZX+ppP+oJGeU2Rp2ELUNaGy4iUL39K1SQlwfQdWn7zLnEV24PI0OtYrkfnqLm3x
7u+vcZDR1P4OCCsN8HQXa0WaLcyD9HtIGScjP+SaVWJnEp4v5/0ZUvf8LSHWB210
tJVJ0kO95QmNBnwLoegNJSnX64YilNJZ6YjrYeuvzrrGPWW7L1QIeIyUjQunqnRY
cTD76YDYQ3n087jFps/ZLSH+zG7dMDf5k1TQOxKkVAAa0q8ELoBPr4vKBZQnOqD0
5Mr8PJ0y9XhczzKRYwqn1yPi5kWUzS4r+eBUn4FJr/t+Psywcn2XR8AXiZ61RyM0
vgnIUWC/EDccfnmtvx2DfSBzJ7gE3Z3t56p2ZFDS27CCEoK+trHC1cYG+RSoyfmH
b9H9ZsgYAzi95crDc0/aR8W+SuIhUhiVJNHRb+F1FO1ubDkU1gFqC1xpLjPspm5w
bzdA1VAv2jAfp0V4T1Cd5bmHO8jkQAQwMNDc6YtzcULcbqVeKHgYG2lePnBbC0NB
RtbtHkm5UpW9aLG3IN+HtYgPo4ChSTPKipAio0SmksRxE14Ms0r5i81XTW8dipFI
UABcLQjmcbQNDzlVm+EZeQRDml2EBVh8X2P05Kxev5oqFwx13gtOBXlFwysSCksB
4cJvWd/2jl6EQYPjJQCePCXX5lRKbK5iyoHKlryP5iyup6hT6YrA9CkUbas6HUn0
fl0SKNeDkJRJ6gFZ7vdAJbiBoTbhtEZ0RLTxOshqbbIVwS8pxGez11QM1KDCnOcr
kLeuuvIxU3sl4arQVsnufcZy4vE9I1kCkXgcD7PX18Tpz/cChHj6jl2PLKS4JnOj
E6i/N64XWuRnqaYeBvg7Dbe7e1+JWPAAu5+U2cO2yU0hDUmB32N1+z+Py3Qa8EGT
/mnFZyw1Vb66+OuT+Gv5PJHogWQ+09WJIbiUysL9xMh9NcgSWGMvTvDPM91zwOi6
1UR2ezoPyNZY4c6qWgh7Ep3UImllPdiruhTDF5bfo73PMwV7D02YShK0tKt9ikDT
T3TwcoXaa1Pg2IrqzLz+fOUdKwcDoXj1MuKnzpEUe7plXJVJOir+r7Bma2tgkG8I
edlrFnxzWevegOr0ixp+OXCLjFGcH82qtZnVxlaVj7qDPZSc7WcrkTYtIuD6C3GA
v0be+024G0mgtmER0tRmTgWv7iGfL6EQ5uZGEDmt9qs76rllmLh2hJ9j/EitXPtl
A/EK762ZEPOpEIYS45SWiOFiX4bLoinKuXwN5px5XvwiIktnm+8nDz7Mnc/bKOEE
INCPPrHFf4c0btHJ2YQyA2jDscWhCMN6B3D/UiahokRlU/Hv0Hb8UCRjbHMI6mLW
7fJdlm5xQPmx85LPrNPHW1TGPUp+ZWT7634JXRBznh5w9dez8yBg3Jcn+qYv088e
Us6zhJuyl630ZaC4OnUP1Eyj2fRtpCnGJf77rT+OCaM5DFSoEwVF9HoueBtsTCbG
9CiKjYNTHpq/0pvp266VBILeQMOe7r6d/oX8kqzuQUKoPxUEKzpyy74Z5V0o1rPy
QY0gKm12aknJaxN3DPub3kG192Io4OPsKA96cJ6te2RW6FJ5RZU3VjHwLg+H9+gN
9J3Vvx/NZqyd3tA/JW4q3MXwFYdl633oOj8f0kS6pufEiy0W0TqZU6SE/yFCtqGy
YhwhRxT1xY8qS4QyWz0fnmFexrtsmz6zyjQZJQST2YVmMHFLaViao7c+6SRyf40Q
VmPbcqB29AbF7PRp0a5agHV75Y3u6eecdAKc4AQ1CoRJ1w9naDYSlvtJaEF24fUy
QOl/hIr6oP4tM0YnKOwjGB6rSgDbSFsyCtZ15DEu+HbgSzzY5gClj125qrYbugLV
R5jxDQ5ZFgIfWTvxXf91mOp1omolr+G+GiSxJQvDn4okcKhe7dPWjmUBMWmIcyza
5BvquX0FBJcYGMaCxXpTbrt4328MJY1OgTvUdt9xNH0kfahOGqFhVarO703Qm5qV
alrEM+jv/WM9XSG5GpsNHrXzSCqMA8PI+wkCeecviy14m4YcHoToVCowGxYQ46tF
xqqYBXz3OuovL9oGqao+GjFBVR48AGyNN1uLyaJ9Zki9Jmjgce1J4ZVMMF89e5gv
NzLyZFTKR5BNKI2HRI4d+yKOY4rVtGymQLM5X20pbn409xuh8qRz2NpEr+I4GOLm
x3dbsA+vWqvXEEqLqZDU82qbCPVdZT0KGQD/u7xxSMhcs6uPlQcLQ3Hn3JiLgtqA
DNU84Eyb9AYQDJwstXpvX9Vb9HDEXJZJRUMTZ6ENaQgTikZosvlaRO9waETQZAwN
4FBgyDxzNdwsrzSgKqD6F/TPI9In2gIG1c3x0McYxp5zv99OwJoV0FMpP8PVW5ij
/mIpUwrOsgrkrYYOGPY1nofSa9VMrJ1EuPD1FBgEbmvCR/LI1GCP7jAqA2fG+DXw
hAtdOnOUhEiqYXUJqC7MSLQK9Af0K+4CscHMt/KlxcyqLBG4QuMbkiVj/n/1CyVR
Uprw4vKnZ1t6/JvtsOTbSdDF2wfzGwEZsKpZSuYpxCx1Wup4sZdTu42TKPsUFVCQ
QywJwpDDxk/n2Icqk/Jdo8rUTmL6JtSzLLA3QzlJwODQv5zLnzbheak4DQ1j16k6
qBf8QC1/mpnMaC3lNHpxzm5Yn6Z+l9nkgD/YuyVgfc2aLW7Voxf+wYu1rVtPxPnn
EzvJRv1UloIu8tMGVpztyEXjUlWVRZm1wueiPYyM9+77HvUpINXJfoGz/q6WA6G3
Nnf3WhgfF4enThsUQ5BEiF9NxiAZDQcl5V64Y8RKLCJeBGxyfZMgUBi/VWXC13uB
zFXSvXIPcFtweGQWAQs7xb1wEKkA5rniBsRpwLdfe7araaHGgSLakEJwoPTH4Yi3
POyfH+Q6T2/lZGzvF5njls2w73tbSAO7yG1FC9ACudmqEpZ+WgTvcn/aeulE2nsa
hA71YtkuqQv2P0baeKWljRv7OmnyR7u2EV6wzSHl+6HaAd0gEQjDVL93a2cPt4BX
HzfGAouTtCg305vLz1p1ujlS74QFRJwhqSSGxgdD//1Lp7Ycane+nhLXoJ+JTCfy
Z2hAJJb9SHIL7/K2h9bg0Ti2TfjI0cFi9JxuPpr/tiCYZ+i0UFL65z2HbmLvEvhv
WG7Ptu/MzBNrvzTFDkb6JUTVpFPsZklA6F+HqcsETrTh/fIdXKGekWYZcSNCYG/3
BlS+38YrjsjlliKUpdT8G2EX1H7kCPgdQdeV6pQ7QZpIwZSFqwhmLbdruVhhLQvX
g6Ley8OYpAA66YD5Lxu/3vmX2gehb094Bd4rDP9Jlvn5Izn4eEqIhwt4jtlILf6V
6z3etC608JrU5YGzI6Jz7lTeAymoZoE/44by7PCTjWZlZMygoLBlb5pR0AUAw1/O
SvdhVBqw9q2g2fkne4fmmCt3uaUglpSFe+ZUQ+wAQaqaOaf/xU6HlLeQIFV+IfBJ
q9OD4ywi91LCHk/eSrMKvsZOT00ygZAakyokFSZWx/AHEUlWe18E0O44U+6kAVxx
8WGg+R0HaRmp90QkCs6JKWFMJfu2GsDZM6PcsjnqxigR6gyDZ+XnRbw+0iYfisaU
dY1wYpsRjVb7kEzd64q4mmpk9gptv5O5JovPkSU0OasXtf/ZZr8vCDzO57v5l4RG
7Mpef1gJjQO92hzsEkS2mjtIoeh8Z2XmKdxxfYAFQYrfAFPfjQMgr746vDwNQ+uG
sX52dUlAl8i2Lz+vnOzbPHmFEbCNY5vjB/iC4+sAWaelX6Nbx+Ok8rwBk8Q/wDda
up5gf5MykBygbl/S2Ck3ZdcHhnwF6mCi5wHXZpdcESIjk/eV3kkFwlGqsW6+MKjL
+ye9/wC+BpnJ/hxn0PtawRf3tN7/8b3uOuVJxLxV3hq7bE9Kc4K55bAcime5Zupa
lN1eWr8unhCJE0/jLmxEQDWhfoykqnArVdWKntPOUZ/41JA00NQn6RdXnaH/agi3
T/toJ24HYq47s4lZ1l0Pe+8pexPfNZpLXlPZEi75S1iv+uWo75OB1r6HhgVgn0zV
ObOa6nAbcJVmludAP45TM0VMvNwfENbiq8CWisKXEROH6uOmFP4k99wb8ToZL/8V
Fe7OKAg/sbKb6z8XNnQ+NSiVss33tV1NYVPcMDTu4Q4stYtQWZHsRlrrAC1B8YDS
O/J8hdOuCuHiRv8DxdkXP8B0+TfMSFJa/9xB2UChtoC9NRWosSrwftt5SZ9tOHMs
7Ut1uEf3tUYpMtsJRQReIBVV71o+Tw0ZZ7c59O67QwuiQLD+7VoHhQ4eEekjmA1/
W4kTBphY+pq/HJpRha1EW8Aldm4HDxMBtUSI7PUbYziz0J716lvaxeGl4ns9sNRh
/y2SMRVA469Uc2bbAwsR4WFvvBuhG1vBJTtJnGK8LiK+WUg3vwsF3vL0k3SyCq4u
LGMLIivyHhFoTIKBNu4vqq2S8VUR6jY5/Z3FDKPGV5E0KuZ9QpwRj1m1zJKNmmdn
6XIg/AzCYhvtODPipFkiI74xxD9BDT2JM9QcaYRj8zji0evB+wTUfa1PnTObAYGc
yncYcQAtVXYbcDFXRJGqq4ZgTGeY713sC4FIdfQIuA0iQib9pmBjQhQdzgOFdV8T
Bx+WaSiVJ6esjg+GlpJlHS1RYC6cguPo2heUEnYa91kHnMgo5csghCfveRY7tykK
M+zcAidNVJf/QGU3zWazjINclItsUXfXEkTVb5MXhS1uIRCP/8xdZJy1Zz58JBPp
5wPRdeBszjXF5jZekXuNscLe38Qgl1ymHC5WMT6t1WfWbam20Tpf5W+JnCYS+mxx
fzhNDG5gfbo/i5458dS6/WRyrkl+6eOEzqpXYqKl1+UhK4PxoLsueWLcm2lbstcB
PTKqB0XHG0+XT3lYaxZ06YUy/z0Ozm0yL5e5Dolol8Li9FgOBCGnTVJKnOEITwqL
yqVWyXR/eI7i1XTmigFaOgeGRqy55R9FdAivHC9oN7lPQzBHPEMMEAe14O6EaWbu
7z4aGpnwrOgWP5iYFG6hYLklexxSodR2nh22eepgsrWuVqrY/mn8iiTkYnRTu0p9
e4aa9zaJaZybPMNOXKUM1+t60U/CgAGL/zKwR5KcmDlov5Us3Kaj2UhZPbUrqq19
680aehypi58C/WMZopYtgUqp/2eewZz4wy9S6AeDBaNomhMGuGnCodQCeLKyEYLJ
QlHvSwAaDsRcdBXSGydcpZIIHfPwVho+vQirMpIS2gXiDNG3uM1rFvo1SU6EJ0ku
d2tDZAISDqCRa7Ei9t/wBTZqBDxSUbNtbi98a+DMTG1lmWhT1Qx9yauOmMzoK2cX
qj+QzlfKYEGukO8lkZccQgMYloUXJEj7rk4sPdB6HdXT9/uPRQ7suduAknYYV3T6
pofCxhoG4tM463mAX50isZ7BgkmFf3J+KFsk0Yu/laSoGvkXXHjMMDUBlkOJI9Qp
QVytlqf2mJIBClbtLCXzPdX2d4X8zBKv5mL8uMx5rKQGTFAYKnUB6fXg862ebuXW
jB0ld8eR/Q4n37g0C1Uq9CzrRlSCa2vbay0BoANRGB0iG6H/+cZVCexol4UCTa2P
1+jLgu8IEuyAs9a+7d5cjv4fNQyl25J8OWuL4HRr1fOwUWpFxhqx8PjSgROZ406t
jHChOxu/e0vHTRjuL2fa+YJq9AW7ZN58QScE9OtkBMY2soRarE2JiGmi8Euiww3T
C48atLXxA4CKUtFT9BkfZZpoyRo5FD7ioGqc08DyhrHjmUNsA2rgU5Ql70P+ZDug
TZ2vIiwcq6xT3YcGkemELaldMqsuy28ub87dkKNc+eIJ28bzwEnSCR6vKwTjUybs
+TAYu97/82n/1tHnwPhh5jooyDJO8lnJ6dQpVFfcXlM/iGPlu7VXtulzmYhycHoY
GN2bc27RACdelZfMLtcE0S6Jf9D5++hBPhNkJMliph/MyoSO8uC5g+3+JxG0DOX2
243hlKa6HGNdy1QX+H0RlNDbxV6Xv/0onnK8sXC2tfziiImQiJ72jHdi4G8b7gZF
HgAJoddlKgUA2cQU+bt8prcw3CebW4b4xhqKIpq/g8FB7iCon8dX7P9xDtcLYxn9
z3Va3m6gPPzO/1ymz+xOfCQ/LOUrKyFZWLOi2pVglUoYN0/owNddLkf3/JG0TnF4
IHqVNTNki8XCASG29GZnXNpOazj+5i857h0Sf+/WlTF0wi6MQdTEPdKcxL87IJxl
ijC2deFQ/ZM44yPpazXEaLnPmTc5zoEJk9GiXnnM4L+8BW9Nzg7tbxeqOLGa2/1o
2ZuLAdM+ZTDPK562bYRawPgS8h7wDd4DvT1Pc+f+yMjanNnI0CpjYBmm5T7tgstX
bVKq8EpAGh5HyEUyaXqkM3ZO6QVlzXb2GS6XevLegO9dabousjCZQy2vKLGcbQQS
SHHSoVId6Wzcji5dqOWY8Y5xbs5eBp3E1LqqpZD59ksU90Y+wHkZ0vaBilV4MIeC
h815YzazwFNqPaDkB73fgs/IvgS2m59QxdZWM4EzL4ZCMZW480wgpa3ws2dDUdQg
CJNdV6luSi2AHehY2OBENea0IKExTaJ5mLGznc2xYYD/ncNZNSaxD9KYbkqELAtL
6gsSIXu4PxKAncm8RbxHNBbTNqPmPZ173lat1g0GRggd8hrwNTWGTbUvyFGynMgp
LkWt2RkBpSfkFLjjiDHsnq4axh+zx3hmboj5b1qgaCPKDYSzJ1qdIbI+Z/Eu5/kX
crnNo694A0/wxquDeQRDMhDOKLHVLtPYxeuAf8zC9tuJ79q86OmgFXBjN/2izqLK
3Mc69w1PJsc5XU6wMfZCRIGnuYFJ0cFZAxLGXc1surPrvVhxCxFcxNsqtCCo0BRs
SlMmrbAo5LTUGeMRMUrFtGKSaCDBNEMnXe75uUZzPZT4fd6ySiHz0ms143CGyU0b
9INx7i9KlUyFnLztJC7yeIhH/iqCg6XLC9t4mDP4gGUfQHru7J5dx3whMkHCcn/T
qI9AGnSbrrbtAk6kIOPaAekMxblf+CmyqsKfB1zapgg4K0o4nu4Fs5TP60O+3188
g0JbV6yVz7nbAj/ghr7jyrvLJZisA62JOHvVfFRYvmX59Vz9AJ/E/OxsTaHA8H07
8m8bxhigsht25bQzO3i8l5URqKcHpu8vbyw2qRYSdjV08Tdg44R6oaPB0oGX+bza
xIxBp7wYGakWRTZtGR//CM/fD/xLGq6ik5TWwVILYU0Krr/ZeOW757BHkDQFurg+
pPsos2/f3vL/h6dSQ0i9AAmXepGyvMfI4A34QRRtjtL7UDmyxd0v/QHdRjUtX5ts
HT7U0I467t8Ee8seGbq2MrOf/xSS879rkiDS2qAs+4igkNAagfkfPwzrCHImgruD
XuH9KMlZWeQNUCQaS1mRIEoh3DbsHJhHuaM0LsxEeInzvpcgn7YIytaoJ87PBaCU
uc21ASIcSMtlYDSN7J3H7py1mKG5iUHL1vg8iFNKtGwQYVnnCm+NuQXaXT2FnYIm
K+HChjS8mzxgTmzCNonHE4aAgXffVdSc17yv7iZR3FYNV2pWnuBeGUhBlzvrrZyJ
nRb6sPmugyAROxGLcva3KIEihsmfWurc7WtedeRgBgrKWGny1kFTw+VZnEFobHM3
VY+e/q1yn2DsNl1s8MDvEYdZyLtheJ9L4ABPkIRL82oWh6T8ol26WiPvdthGdGBp
KeABCZW3UhctodFr0f7zRpP6fnjAM2VAu9jh10ofyPZq9JouR7rZF+REkRfvcXof
UH/HwF/LZaTB71ZLbpf5BuyVtyXCUAi2+fuPijlhsj6QsjWsCmBwE2VYA0UalayV
wpI3pPnpcQfBU6ItKnH0+H1sRuGdHNG2VjOesYcoVnb6Ka0DizQFTxh3CJOBnEBh
KXeRWEdKAajol7y/94WBEA8ujZSMrclZZshoTAzJRTZ77yJ1eozdAM4Kd31PU4zz
TvMfQQZH3rhkKbpFyR+3SCRKI7vxIK/E/kC7iyAtq2oNRd15Uhc7eDRSisdpS2pr
IbfoKueOUqvKsr5lD6+tNvBMCH6Z3ID5FrZ4nTCLt4t1RCwf7kokmavBtk/o0Ies
oU8WE05v6yeNlsNq4BhirajJmuK3/F52FA1fi+nxSn2sDcMQFqCTFbopzhGozxRk
SzuovbumjWy8oemBxrqqcvduSmjgzZ+erR39/l4kKHCy39SinMNxjZx59ZEYW2cf
kkYlw50j6vxaw4XEOQY7Q81DmC7dkwQVNXbfnhImzwBpveMuvyqb6TDfsVjmURNy
9z2yA8ZjUbAikUYHxsQsfhqyV3WRz0V/g74ZvaCNjRpK6uvvaB53omGle4+wP1JR
CIweNEZRete5/aLqK6rtwCTw7wlGwkwitUMMmRomUsPfQYz/oxTvexDODQSOd9eY
QauD8mQvr70yE4xLNX2oVHY3Ul6MfnJcjva11yEFGbEhfDuH+1+Cop+OS8o+D3G2
1p5E+dZyEzDTD1lEw/sZhevlEqP6XfCtpL8kEbNivskPsGYo92kXK8m1GiKx0uXa
ChViJNG+dZAzLyOe3Tl7wBU9l9t0TmyceqOuxKuFxj4Rn0/rUJkEs9Rvg8I1ILZe
VqjkN8/SjiEjPfWYwyyIqFxhFF8D9qL1NsaXhToXV6O7IVnBC1HqAzcspT43cyXJ
ByXCWG6aGUVFyTyR1ZSmkUfXYVQqZ5CZy7TLz4+cHDLCWdn1lTmGh6uHHIJw5o78
r8ihvXERH28KDIySFtmuz/7Bl5NsGNMxgwAfEibih8LeNUYqv42nBc4n4AkjF7D5
ouKhlqW0A+/rUvSsvazYVr0PPhtBekWp/4HXVq2d6dMyRyx4g/5yR6xOvKBWodEc
1TJKbzDejfFJLaDOQ4vytgS98DGUH4lig+a759zljSu3VAS5lDuYpBDsnQBScb7H
ASIk4g6X/tS79vMwRnmEE0/RoGn5i5iQPxyAD37/IjpZuYuZKfyfNajbbGu2b3za
yLkQh6lG7t85RuKULfueyIE8fOx5mlM1xL8RGRMlOLN8obtRTShISS/qgv+c5aV+
TrGVwg53UPJZzNJ04XUhCv0S7iHwOJd0a1PAun7BpjUnNKEs9TydroiUZaIdnJ6C
W4N6WGrhBiyWkW+n6VwVm3pK74Lzx6RPqtIG/2dwenR+XS8Brc0cXjHN5zSHHpTE
qsdn0oeLW+/qf+tSCcLdoAlYGdKUoQx6v4TAP4X6FuDg61jqrQEf74AcW9h0JtxK
MzJPw2xHjiQZBAlouOxOdW4TDv8EWzSQ+AxBPQwg4hbc1ezAIHImjJ+P5Zh57fAX
3qALNJE+N1b6y87MxWOQcebPxh5kWGtsE9MPPFDZgg+PBNfGB3YNlt0uVW7nHlHk
XUcHOTJD8MuddiKkU5ZovONzXcjDBRFdH2qHNzPoh19K9aMd2YIupJEAdWPw/Kh3
GFnJwsWhXpHMjt9Vuu8sKXwXa7wMNnu06OirBD/wl6/LntOZooD/JGk6K6q0qzql
lC5WzEJxZClUlfJQG+MkBLaOxXobFBHlHclAjInMW58Gx88TyJZpeh8WLppS7M3T
0ATVO2gPIH5v0mftxOqkUnKACqvSfxUS0VWmKDbh10twlTCRZqCtjXlcJ4MEWCGY
c0gFkWV94n6Ejswnq5gbRmVtc9KKKKsYXWP7eEzvskfyrl7/mfk2NvS/X1aKJoNT
dQnU0l7i8S8wk0whK4zz32Ab1hO8HlCceseLvZl/cVYY63n8urqgldSFdnDLcY6F
drVPCa0erXE29FKkgZ3u1Rqe2aNLAwUlumEg/pbIvCbjyUZ/mPD2ClFgoSKC8+u3
+Pytqwq3d0bJ4eVyN3ybu0VU3+Mszzur7UTeIwd4z8B+uNLPKAIRQ37Uhp+fPuzg
CuMFJ5jwtDD9KVZscW+IVOZMySFvJlzUYiI7tJG5KA+J7xe23ODlid/qT47ph36F
AZ1DFw//ka3iX/iemVPBe48/QEjQfnUTUTefDSG7lX3IZOCI7zqeP3qcLDktR+z0
n6iltnkO/kKjhHGGVVz2wQDFAXdtTqz30UA5mz0va4MG186LDJwPxILGIaoYCn9w
/YXrH7GxExZuPUYbZmwWxuivf2YVYdpS6mBMU9evbmDlCtvpc/1wuV1DgWeveIRR
X0rmPeO44ivXcGtH0acKmd5CHRnAn/6NFlMEO0PrNBToj0uh+g3BrkTRDfKsLt33
zW+ORrPhzSWU8iRgjPjBIFpc7AGWaFJLCbu575P75nEMZ3ykw5GMYWJf6bQjsBnQ
+Fb0dYMdQfat+fYTscfxzm4nAyWJWvRofto5H2h7BRvTqkujNxLzx5pv1Cjd2a/D
Bk/XypNPg9qKPqhj//8fFdJhSqRAAhgA3+srCzDYsRGMzp11uMdeMCq1lo379oiH
dz9HXs5Or8bAAZKSV8FrSCWNooMsG+Z/DqUNU2oDvp5dFMooNuFps5nVOzCMWolp
QnMhjHXP6Pu22ROaBtVdcjpObYcgBmxVi43s50iHe38B3XoIuGwn+JLKFZo5sF/q
9jmHi9xmDhLietynSDPF5AhJo5Ee70l9No0PTs0ZSbz+8KBNkINr3jlIdYcbVOw9
TEC68DeP5GH8PyNY8+DbEZq0Av5qbYqrm792lhpnFrN6Y2CyDpA5ZKuRkrl87Yqu
KqtRqLI3ZfOqhWgg4bMd8H7VA38HM5DQqpGq3oWo/3GmpZWwvN26kmWAXwcbCzzY
FYkPWLSVscF+CJ16eMWJTM16oNNJy64EF7oAzvDeDEB9PHM3WEjA7+V+kmbXaHdC
Ulwx+n5ab3SrRLKXBYgoCc7LAbnxh4Sd9J0AkUk3zYTThcCtuYJwjTPwo/ZAzrNT
6J4xa+alT9syG+mm4bDVqxFub1iW/SWw/vDmI3t4BsZeuEh8Gqe9LgwQtz5RNO6N
A4VlzR0zJhyPPzM+mQXswT2ttNvCBqkokSsbX3OxtaKRCOJV1H7SMtbKW6Ox95oZ
qziz/EW+ZhqnjuC76OiYBmcBoUNFU4wpnCrXo7kj0NtHBL00sYQV0WFiYjDGVP7Y
Av3QAgCpruuAOM+8x/pyNuu5fK9cRV8cQ0RHWrdeWfpGz7MAXY5kX3y9XLENOQ+m
JvG4EKDqk0v3nRG1hrBDIVEOyyytsT93pvn9u8hUSsGxF3Mr7E/HCC0im2tF71D9
Uji/YsKR153M/Fza7usjE1flrSkQUyuzIBMQg37OS+z7/i+cUOgccf3FUszgD521
LjHv4Vonf2ygMlgxH6/iB5mIicpZMSRA+EaVaSkscQBimUN5jiKc4iIYmx/Iu47y
tTz6mYvbdtc6dxnt7wfYVLp3UE45HTaoxn9fzM0pTVmUHgYMGHVqgWXCsc8SDvYu
B9WELsj5MLanwLOjbED48F6oqrhoeuYuf9h3NXxRl5kaN7sgavSemcVKnkxDnkeQ
q/Jix14yZUme7hBadD4m5UfPFJyPvHassxFskAtOEh1TV3T93J0DovFD4b2VwLUb
5ihvFvorDBU9ZuNnAhBTGTK8jlak58f9HfNbFQvdJ3+fJXZfH3jWtrqcuubfTAWE
HEDugn03eTmXx9M5uEmzvif9xqUcsrZqucYPFt8ormBaBt5IppDdVNUfbnrOrNHO
rxX7+9PZDPxioxXkTGFzMDud1I+6UHynu87mzzKJcH3P9Y5orzgs/PlVdH+jp3mO
MnW9PrGzyk+IZSqZZQgKzX6+IUL/HDqyuNEUyLs8ONAPNnrSVKxVrrBpm+7DvDf9
+ZDNOQ16C15kRAE7YQjFx34omzOJDE+NWK7t4ckZCucqqmzeTUNECyefwDxPD3is
hEl+idYHsx26mY/etJ7tlmnQP8rKnIduGtaI9a+rykdAl2/o+6FveC4JSRIAGAf7
OVN2a7uuLB0VHR35EZLBchpnQCr08HcCTsHd7UBR6lJ+TJe6mPTQgye0PTULeSgf
KHNXRwRNY+whxJvTtTsc6ZDPpAuWFge+v4VsHLb2AQRF7xyJUG/CluSLpuy8gcLC
pJXOTxB3N+NY1r3rahyu99xkkbNIVfKHrW4TYBSROsES7YbEoNbM2rZIjUYU4yPK
LaiRQ6EfPgwaNene7OW3xVI+duKLB8e+HVHOQ0mUYy/q7cZDw/tvmy6m6iEuRgZ/
wJ66DFFEjMd11JNud9hSO+UnI4ujibiOHYh9SBgAFNiwUoUrRNdPERmMjQaUE3WI
H2KTK8o1gcx0nWXZkZHkxtQY3SXow5Ao6Cqw+FDEe39uZ8xil8mg5EvkVMgkMvky
JLrjBPRdAr569Yanax0x1F1SU7X6ro8S03U8bGS90MAW4ZTuubZcZTno6jCJGUTS
c9BGn0DSvkgEYiaOVF3M9GB+WjvsfvUaLYgQdq5v3Tlf0RjnwPkIdj71j653w+lb
AZiC1x8OiBJLb9EHq97yoNBc0ArNqKlA2rcdRXYpuZVnjdVZnS2K3LI2XD/yd361
5l4iQ3C5HiPw5goTgdu/C7bw6pG8R8GmB2X4YgZdeRFzbEhBXQDLb01+uDgtnZs8
+K3goIOpfpK4H1qylalR9frYIXvm8a37QPz1IP7fPTrDKF+U5dMUbU6/itfLOBDf
xTefUONqTUfioF+cRaaTRLJWatq149C8UCAt5PbH4eZWMK3Mq1XxgqMnu1S3gMvI
wFSWdj+oBVU2muP4hrLBk4pVUuFDMI2XDnHOip9NTxiq4nHihSnNmCUsjxb8VO8K
pXe+8NYWDwcOI+so3QJUvKygOwy/25Xmx/JuB3DzEOMKi0xuPngd77gpNz+alq5e
OXnPtSCEyAZ466M/TbiUS/9Oq7FTL9BoH46zSINhC/bF/Kn17rHUfgaV9O4puwBK
10Wnzs6bnVXtWjx2CUZob6nUsxLkgwFanAVcNmJKQyJi6Rf96Kbddyj7kE9vC7bi
aB1l4XbyFbC0ZWhHQxPCBLUb5mIugKnYAWLRCBIpptxzC/bvMOTC447+l6m/vGmC
yMxUK/Nmc/+OS8FPT+T1XFVXWE+mEydjKbgkGPm+XkmOScgrGDdor9y9B0DyMAaO
ZxuauYkLG58Ez3Q7F58fcOMhnuP7xLnARqn+FPP/6I2ryoOYb9K4luR3uajVw6Jh
gxOVENCfxVuZFSYZdy8CGqE5I9irxhrwowHHceDov08xMiv2jZYBoVkp+A4106WW
gPnfgSNN6AJGoYQcZtur0TSpS+wih6NNxzudaRXVLGINAqnZO1iEEi9uvtPTR9Gi
VUyZTxYoRS/gir/cAOYY61CcIMS74zOYamkMo+cnAprw3rNAlEgxaBntG57/ZG+L
Uh9GIZBWEWeim/nXOKjWtETkEla66PTzSbOn8F11dOjPvlHM+Q3QVPdsZSMdn0Nw
t8tyC415qS11dR3Ay0/3irAKIcRTOGNkvuvO19XCHsbv1hQbcPTKjfZMNjGQqb6Z
Ui8sWms2WH9/JvPmLTtrCk0cUw/nTFdy/3LKfiaTB+055zaeOESjecmrdroahbXF
2dgRElWoyCmiV/6jeQZ3zK1ppuBc2Hz0FZRV5v7AH5jDmg+172AWftTustqF9aOg
35SLS1ESugjDPWAsrC74nBjFKDBM4gtlehtlW4RM053v3o2Eb4OJbqqvqSueGfyR
oPXXWN2UftV8G6W+WWO72Wbv7O2oien2tjOkrm8RY+PxLvq+s/JUkIVlY/8i5BmB
XNGlDvZ/hNac0e3BaRozGXmtO/t/vuWXNySeGix7Xy+46g3dtq+Li3e+UktPn3qB
c58ImR3c2Qj9Dk5r1f3YBY0ZzA/xkGuaNBiJMC9+lr89iuIzemmqYzzdA7mxyTEE
1IGzOtnE6Q69HZIGCui8Gd/vPbJpG+ctxQVMqBECEzJP7HiWlfrmeWTT1Q88N/DX
tDh9WHvb5Vn4b9PIjCZsEQJRSU+QQFvzF3bilL6X4ncRvV4C3WGTdatrYGsIp+77
8yekH2Et8p5usS8qVYTiCqmzmkMCKwjX7xelw30C+TtgTVrRRwPeTaWbvnOQNbhD
85cDr94WHzHuOXB0pG/7D9RcXSEnkTbD3NjNaXRgCw93rMGwBsAxXwJHFMHzTnnj
cjnwBcCoMdzEyUzGaxnYTNfyQ8fGfP+QXUsR0auTDMeXOw6biU14EvdGjmQaDrET
nx1EReGXmh4+a5S+XtrnSR0IW7MV0vjcEilctLNFE5IXqA87h31R/4D78aQqlJF+
YH7FxQA2wDRQoR2QyYwGLOcCxPf5i5urhw9IHPjcL6rpYW1rwXLdM8FEfVBToZeR
avL2N76Agk1Hbe4CGrJH6mMPfuOKr9FInQdI7jxFJ71j+5ZSDdSepZq+FgPRf7iM
JuRWR4H1SI87R26boxZ8vt5/zVHPChLiBgzvnMz4Y09gve6BSWO5kJ2rxqDxZI+8
dVwNUNU+8uH9dTbHFKMK/myEorEJQSwbrp3hm47LoOGPwgpGi4ddX+iSvnbAQ3LO
qeGUjp4DWEnw0YogxC3HWrnsp5pTWYxRooVkROioln2U8yvoMtuLeGhQCeYEwEVt
BNzGIXnWvJJH0518PZyC7B5rKfWUQ7sej/qloRuUttu3MvqmdGhfuuOEJDEIPJiM
0YNJsJHF++O3qNsYLPrQHCYBfPIRhCtEysTEnRdZSxfr1B+ITrs2nNTmnphW92Fb
wa6Yd0j7f4MaIT9HpqNRy1eb/QTeclSQN6H2go9LS7sf1LvciqWE4egYDIFjDNKA
FcpMjQ6wq1rJNVpkK3ghKS0wSfwHFsEZo12WmaFRnMWdIyKd25Q50Zb2zNNYJ6j3
fFHFf1ZequXhU7gIENyOwpfD5EOcjAnu3Nuiyw0MsBnjNRVwxkGxUpY/edcngw4a
5ylDJTgjyEnNfn4GuwBIjPEgPYd+OiqKjTCMWLSLtvz7fdvDgvAkkpVIO/e+42hg
upPeC0KWN39OQM+MOyb/oKdaaWEy7J/MRvbeK1SfrmvEAoWIfkMUWcPXgX3tf3w2
5wE5/KHlhAggmWp46v0zqSsu1kYmF5NLE7SzymuVt46M8qA/6ULfkAbQ1T2+9P+3
MOq0/DyMt8oHAw+Wp6/4RZrwE+hm5iWnaGnOvVRIRo7MjiOdFMV/iiyVsM3rL+l7
raTkTraCSDrKb4uvxvJnZbyhww7Vw3jRJRVFf7BV91QB/vmyY/BCybd5ZClJTuEs
trpvBFX34vfXCnKRXduk68v/+XGot2yhhj/erR3SIN6+9x/COnR04oYSCndtdyjA
matgS/mT+jEl+REKx2ieyb8HpDWruYf/24JYAXtzMouSi52Koi9lA3hdrJoAK7e+
8AHdnGQSE9aOj75xsE8IQ/zyyiBgGBleJQhoUKpWh/j24FSKYd/28Lxwwpj5r/h0
/gAbCjK31UUoK+PUUchRiglv3y0XJvA2Uyy6AZbXNACS05dI14or4Yk9wIbUKeVp
3S6htVLO8OKT6Elyx7U5zQXpDw/W1WPrq19/qhgAjbfvrk3ulbPZiYzxkR0uMisv
KjCzzN+XwsvtCVC8reQDxTj+BXNf/mp309ydZfcN3UdP5hupAQLWz8YnE9GOH2eW
lEchQHf8FKnEeGe4LFFffUiWJKwfUELTmOH+CIGA2wXTymGKHmT/Fku80sDMPAbh
PAGpg+NInKXljTVtakPKNBskPZ6Nr7U6CqaCfOlNxA/YDkpfdEwmnt6oqdFWjYjn
cPyp06ZDuZKvmHiJFJFMapDvRpv1ftapXoI20PRWGfAf6rEf+92Kyhile+keqitD
Hj1d2pl6kaD1JPl4WP2f8C8UVtoRSwC2snFNK0sTiqXPB8os6SbNrPwvBveS1zxb
Fz70ISofl8qhrVbJXySHCUUkishDfA6AI6i8DraOCQAw9EN26pCcYjcbs9s6jkYl
2Y3ZsPZqlpfYk7Hu7uQ1byiFvB+4AfIvCJsUZYPgORW9hSouqiO9AuXRlLL1I0i0
bAXr/v6he09Ud79uO1S0igKZdxBpLsNZGIVmgy6tSpC1gniwdilMwdEiHIuu0Hab
EAU66WD3M2q5zhLf68PJFCCSjf86D9TDmYX09ZJnHBBihXxFbwP7drK1DaIM5zNL
LoalJwIJcMUSNQHcK3rwSfmVpaJXaasgMwj6GDSARdJaHumjY8KUmWTYYY+ufcg/
c82VhUi2/jm0W1u9uthlGFTwAP4fG3YdBOSrV9O5A2g+wTayE2lLZMn0bBXGiFfY
PJIJTGfEIH5TLEsEPaERc4sAct9kUDqIB7goultpAsWCZuWj8QLY4UBRZfPnXPvw
rABv6aOqDNNz7uzlBDHymiCmJXTZ0igtVhB7NpxM7p/RoMPwzSffX0rFGDniPq1i
nG+vycc6Eo7tOqk45y2K+vpfYD2YO+OxlbxL9TrYfOmZkwJyk88IavpeUOglXLM8
/WWm39/Ahn2zNskoGBscdDiXUA280dJ6qiFe6YW6ihUAx3gHVZ81+/zzlgcrbohW
0sNbOOcbiSij+vYJjnYaoCL1zDjSbf42tnI9QBr3Zdz0E3dtz8ecMXQqdeRAWP03
nHNYulcNr6To3fwShl2KEh2owozeOXs3E8bMl7OoiK4ikoc5XnisMNe4qGJYDIeM
ia4hY4XbKtdL3WMaG8+ZQhTKMAg4BVK/U/pPhTfxcJheeoLRIR4ejDj5kpuBdSQJ
wv0AM24tVtufe8FUSvgeByRA0o5URctevQDbN7emv5uFfD0USos1qRrmxxBj0huy
3Xpy+v+JYIzKkpVdAd+fgxYduKZ68ebNCQfgq12op+FSqT52gUieBEZKbxJ89rya
dncJF18FzbyjqYjNENsS11s1ynHh3xW0BIumy5pZNSkW1l3Dc3dw2CQmLKL7TAw9
IDx33YWnTM7Lm1aHTWvP5ujIdfQqlBasS85fbSJgB/vqbYaO1YyoOIb+V7GvOMtH
8dYy+M9Y1lg8MBXE9KDn9kuq97XnjgKbSLTFTVxXHkphkqZrq/xhVQCXMJM29xDr
Vt25Ef23pVYy4wXM2fmLNs6bkYxJK6/Ew5gQXvC8xQtBsaBrtTfGMzTdhivYxYWp
fu04EKF5sNhi5+SDaY4cIi0QfQjdrwfqaCje+czWW4OLh+w6z3MgiZrAIRTeUH3f
OgdXzk3z7O4hWyinza1b3A7rP9N09MPHnmW4cNR24/f/I5AKCMBZoks12sRuFfib
B7t10KiCohU1L6Pu8b947MRNODGlQc4228ipxWLqOULr/YgTKaGR45sbViAYchU9
ZHw7pT3egt2++CKIXUaXg/hyANq6ol+OnWUGxrPiUmcQQnIXPpQ9xoiJ2jESbuUA
Rg062GdoLqVgbW/mYjDfN5xUM7TLg4Vx9MxSxkBC3Q4EjfGnko7dF87+tNnPfg4M
FFFWdIqfajhejnV5ai2FSiWh015IvfojfqtsFnUfykdVy5mY9cNNze6sivbJNGiU
p5P6+P9rPHuyxPowfdSEczzJe0GdiXHOLzyl0lYXEuqj3fkri5tbUS3PGQgm+w0Q
DaCQ4dGO9QUY/sm7bsIqW4EHHBHotOGa1LigSU3kbtu++B+efaOfp/NCjbGBeOjL
SXswhDwkvm8qyw23brJUApqU6VJcSXDh7oLHF+2fO5eiePBqC+bNE9j2dGOhTaE6
gJVqyzTHn8a2jGQGsoQKRmD+pLY5RQYxRPZvlf5B/ZSjzuC9Aup6iiaHPRItVo59
XOpfrv64HEbE2MyreYUCBUJ3pAYcivzufcO33bZXkpx9YTeQIW4ZnKOldCcJSZkc
rfxNBXCiah54Qj2ao85ChVctK556Yp9JahjrP5+PwaOiPVcDmfhYsYRIXE2RNHy3
2eIvw9jFLZSgj1c3VEiaw8vbF9bzOIrY+RePnWnIvV0ak4IaORKItjCXufjefnUl
N0/7jd6dZofeC5MwTVGvcMJD3W/6RI32pE0Fm4Gwd4xYt4DWc7nU+LbJXlCW/jZ+
teV7dkU2n4kkvg811nmMRoBBs2MaulOdxqYpPSyptPyPPPB7kX6nlWhfrQ4QMcpm
2+KRGIMEVkOEopDsOOaHIfCeE3FkZjBJvibcYUPSSuovigkb0NNrWnJHDxQerKdM
uWlnHy2BIopTQnj3+oN/Bry/eM+BT++UJgxjEmP5EEavyFjWJtyGev1uLssH4RK/
CwOK6KhsnnvfPqlpBXWbl7CHvRJuAYx7tGrGSs72DeruUnJej4kz8714BJcc+VAZ
mo6xTo5UyBKXpz09pm4rB/yjce4kkupazGP1B9vm6G0N2To7bI6Rm6isBSPSVcFi
whfR1iBiPpO5YQJFvgyGKmLSJXRcIGZqzdLLb8eLuZY+ZQhLYCoCo9EqxRDlOOun
wV446+1lbG5/3sNuu3NM9YdRN096SSwJu1wEfeDdJi8yZq8wLjCdgHCWkX9xEUl8
yHUSkV6msEjPDh3Fp4sP/MMYaBUZt9UxrcHKCv4E5fmF/PI0dgdbW1sNvpdta0HA
Cxxfjnc7mig0SHxVVTZW1zKlvRLG6kAMprxPXhqeLXcR/x0I302TJZPFQSqhD1aN
w+aL8kaMZsQqHqbLQULjI6VE0J8KsKv9XFwicMKGHGwF98fmnl/Og8CISWq/iXav
espw82t8c3sRx3LyRG05lUSUfDfw7KxC07f6bZcxNrcA3OfUbeBj5eehkWKyg4X7
qjcaIqSb6uZqAbklwFL7wdlPWUuPhmhnIHUuzJyvMkjeVwZhlPlmOspuwm+KNP0n
6RcXBeRJJ3RDqrgQWE2UBew/Xz/1mxZq6/lt5Dh57exPntlzqAPWBomYn97/FmgE
NSfyhAj9EeZOwBRkIf4LkczpFTKb8ti1wOWNh6zBj+6YSlwJP1vZHXjnSxscWu8F
kNNK9N4C+XToqqOwLYbp0vcrW0km6XZ/3aDcDvF+D5BkodU6MfXDZQ8H25nArSI+
sFdN9hAyOdv1CbK3mGUwLvmofnivF40TIExrkWeZP3A9ZmpXDvpH+I37X37ALgnR
y5g7rQ8jokfRCwmlDh9RmViArHSIlMkzafKD68S6nlC0DP8bI6AmSqwMUcMkIWbM
aGt9IHIk+xQw8bHUXEDDvVdhez7C4xejtAeQePk177zxbE6Yz71XI+DWltiw1Jw/
qUIKeMnTXnrFaTGJIEGdO+iBizH4DHphfhGhejg1kZAWAP1TWCYPTwb9x+AYUVJU
42uQngUMtZDZU9xRX2GCk4/8sRVbqRnAY+yp4RgnZ6AIIt/hhLgLL2opcLn+wbAx
hBeep+K8dvY4INlnWy0tHIDa+fjIvj1NlnIWx8D7xU0aiA9H/a127GPap4utKwDn
N4c3dY1cUf4oylPTH4ioOGETtXrgU/dcW2UFD70dxwD1eMFJPC8ydSLxQKQbQKDT
eR4huhy9seOg1uY+Jl4YTnR3qOBbrAUBy+QTgrUsdBM4RI2igFAOby4mqSononVE
4l1tzBaRsi/Wds+xyl//X0bFozYbUkP+R9sWb/YJJ4J9dGuzlMq3xIfgP3+/Akwg
op5mytasITwsHO6i/Nsx9EWd/uiLWH15+1k+iCkkXfHxSc2oayeBkhYwQQHPOT79
nJDF/ZNN2jl3+OzvIaNBkHSWJndw6oNhofbe63IqKxVIWsU+SCdeQrtaG5jiUJPW
LkriXQ6FcXZtAJVRuxXPEr7UmPTnayJPaEfgARZldL+v847V9NCD80jpdhn8c++W
JOmAR9nlIpKNIO2iMp/wLazuiAJKk6likzUMLn22S2o58agke+rryJGMYBM///Gg
Mu2xo1H5MB+66yHyHkJrUpNeJRF25coLb6Dbd7SYVAhtnsLdvI1LcPsiRYRikiWm
0NI2OSjBAm2ChYZH73RObpQBzkiBkMSDA2lrh4oQJu4lijxBsA7kpqhCc6gSFknt
h4w3qTT1Eb7NrFpTPUt6c91izDvRyegoJoxhtZgstMWMtGyAfxBfM/BcHRd27GI9
K/7GmZlc38LhS4vxqZY7TzYaTwTSymhjNBkSfUIUPP/xLMu0Hm+UQCSRw3I0o6Ax
x1949qaS8Q/5Q47xZpL8+y6AJq7boml5LthSLFi5wjiE0nzMK1eVnR3/air8N9wQ
eOxXT/PaBhDKPQXBoMhwC7BXgukUyTL/a8QuL/gn5vUlMvDDiqlpD5WyHkYxP6DW
auzd1QNiFuaHZ1lArSDq+Rv94mTL2ZAkJwS3Qi8A0H5fQkMw0LViiDK0e1Rfl1Vl
5UB0eGdiG/5stPymsDvt0FTU7KTneFu+yUEKpxvwj3I6ZQF/bHtKtLKkD2IN/BZa
OP+WkIEIVr8B82Etg82XYdPBgEK2gb8KLgdFYczfL5DkBuVH6qgST8UhEVmcmQ+C
LBxiCJAoJVvgzwd+8WzCFcdz4sLthH+pZg4Z/YqNm1pjTCqK0pqZqCekq5BXVYgI
X14jXCJr+M0mnBSYrT+TfVIVVvsv75UuKsEB1xqjJzIh2xPQCnrREUB77ofhy/Af
hv6g2fXghHGWsjwVYaFVkZhJrJCflvUgOdyluYhf7QTdYFN5P3FZhfR7VOfKwQAk
z+kdswyl15Nu6zQbg8Oryw5YkgFiUOlMMfWmX+Sk5kFOoszYVEzRznjjk5R6jN0a
exPc80dpuPcvf/9H0LauYmYcE6mDBIDwCGX04HEPvrbvT8lXpzexQhpTRssYvpMb
J1BWngT5sbxq5FGJ7PlW1U/FHwvbxJPz607ZjLctVN6Ct26+uJvHG/KuXAkgaIQk
nd4ddjsojQ0DSxqVPYQL+6JtrYZNqhTDDLOL7G5x58f+qhx2SrqEK0skPoqigC4w
fDqj42G6QV4PxNV9wdtlgYVw6L7wfZqBcIoLhNNrJZXcnrgQvwP4P/bvlwWz8cap
vLOuySL2ghfjb0AM0eKZBAOVlLRKgVGOC4L1sLZiQtDs6i7S+1CymPuiGsMGiYOA
rwQAFDWyihmXXP5yYL4PYMfLCc+2Uhpy+likRnZ/DDlWyy9OZaXHiGjkP2qo015X
6oVjMgOSCsaUo9iL5ZQfOEqea0zNldFa6EkGAJD58QDtOmJImwgJ5DqV9X6hhqO8
QM6GzPo3agY9IEijyJSwHaTvfBQtZgsTtMUyM7bw/CHooG9THTBrYMviYp7CEGv2
BMGEL0ZoAmuCM0KFfiLZo12ISxRrJ0TtdTuehq3q8+Oe7Xk5IV2ATqgAfC7CT+Ce
LvReGm+Ca+lhcuUYCZdFm4dlosz0nGFv9YsJHGIAV1SqSNAeXVnnPpLc1lnVIaWJ
vrypT+uaA9TPN77ZahiQ91LtN5CALomHoSgbn1h87CNLzl+/YpLAxLICsUK0EA1T
HDOigbbpSJMyUE/NTSOZI+eZy+D80jEAOdkehJf5h27S+h+/bgLQrSmzZAUmUYzw
bSn3ppIVudahoCZlfp0l2YyuhEMa2dApdnZatcKApFx+05bxZOUzURTRHaC5cL+R
ONl9fzt/1OAXduWQf0Ra7oMzZS6zcDii6gLejIVXTNAlkhLmUWjqps+6SR0GO1K4
jsQZpVukkA9ovSdCoI1cLYv9kKfYeInAYPMntKKjcXpaoP3zDlwepBWLBF+0MMmQ
3f8MPXHjdCGl3Nc5mv1HkFIRKvuUpyoUQmITYTl4crmITfo9zzQrfE6f6b0tB9DV
x/M82w9QNGH9OQmG2HJM1dv35ITWWTmNMFoBqoMoEo3vG8Q6WBW68AdALF3oTMR0
Nmrqajls7Xp3RFgcjA/Ghy7NCfm7MLM+VgXJMQkz3ZQxCnBf5FpRn3KPDH2ske/o
ENPbirph3wiIJ7Z3bgjlKtxjtwP1e60XRbrcUNSM36OUo1wdPw9Tqz5G//OKHQL7
RihBHr9E43HvqNUMN5Hhpa+QwnnSmGJvncH0NPkAiskwlx/uoqkpEOiC2TRGIAFO
a07Lg0La0kGLV77zBRpayIZa9YKSZdST2K1teFZZFns3p7jalCNdJsoY2HIIMzBm
0ulrNA9ZhB+sk/SgI9nnbzkYlVXRpBPH/pVxR09zgBs63mgojaAXUlcRYUCijy7b
g4ZMw2rJE/U3nFM/Q2Ua0Y9DE88zVvjSFxq91n1vh1vqFNLCdGMI3GK6pfzNNPpo
jUWbgEcc8yoZ2Xwt9gpwbd8BOZFjupXnmDUKVwbuNw9jDJGizRhR2T7SDqAxX73E
I7afltjCrTbtnCfQnLQEdE8NN6eRf+zbSGoPjWLCB2ZcUOpxOMW/0xEi47fHy+p+
VSvX5aRC2k1Fa/Q6pytAzYg1pNx5kvKCEJ2hyWNcArWuF2g0SikFjrs/8BraTAvV
IHuiGeKQm7sAsOsmZp7J6XPoGjnMgOq2M/GUxHZTobT/HVDWVkTYGmGuX7dUfNwJ
BlnGMRJqlT906+1QgEEMI7fbqvePmnW9Hf9QnR9HdxxKx7Xcy3mx/yRzbc/o7H4g
6g+ZbsKEyDuYkJAhh4LjK6ILZswh9EghbE0rtk6WN/Ps2rlLJVwU5jbqCbGngZrZ
4aiFw1XPdfJAg+Ryz155+a0eTLCWYMAMps5iDAZf6pwymTO6h7BJJz90KGrpTqrv
QCi1ua+JGRWIhsFVq7HTswbSeVDE1J5F/SsY4IrOMJpKx3Poe0ZXZx+Rak6Oqej7
3JRvodlGGQKccD7hN84sXEC7olk4vLKOdsXJIyL/edT1GiZG3N0cm9W9eudTpebC
oVwDfK1AZIPgwkBrh7cqqfSYwwuc+QYhKQ5YOaUeLjdHsi8zWbU7wVsG+3f1DM7z
DIS9GErLiuJ14SdHY1B9v5cBweQdmwBA0gycICHCgDIkUUm8+VXkj7jOIKkg2dbw
oNvmTx7HpMCJzYFg8FANoELT6DRDX+2fgwCa3XIyZZPnfeowhmqSlRrp8DLb3EIS
6+zBMmC9UDCM+JrZgMeU28R+2MZVrxKPCA6XPBHhAlOhKQG83GvJAwfg8ZWgxwjG
jelTIdGM8x6aqiOAgn7gALP7cISEgLP3CQk5FJrLvfcvnfvUqSMn4YPOIaZBaMS7
dE+xzgmUMPeswNstatbWUaY8RfqIxGtIerIS+2Elcz1iG9Cr74XaJ9J0AOyf5RbB
rIMKV75sQstyhdCuisnDYWru1bo3ga8fIcWgTRW3tR34LY8ZcYmEc2ssm1xXan8o
vnsMDh63Ev0gsF5rQm3WhQgORRpoLzFfD3CPH4WCrv/C11/TticTmxZPdIyGsDem
3zhYptv2yFnWomR2T7uwcDMX/uvbiyiPZpH9Ty2SuKzgx/1l//A7CuapUcMajojP
FYBNUQhbdn+9+p5Js4+wqU4084dB+Xw/eej+MZXHrA3z6eY19K4JJImmYCNhht9d
IilMvyTNJ5RLOx/oLEjWjfguhIA2bFGtmDCf73rgDS0mf4J2a9Ff7YLnu6vTDahn
rIgljtcM5lI3wAVGQREcRcKSPPVLUBK77JmMd0jE3kdf3aVp+4pqDZOhw9gYrDt1
nQTzmTgm9k3G800oAUrlc128zKLP1A9rsmq0TZ9g2Sly/fqoTNCzaNU4ZuU6+vFB
jAR9YR3HYDbg6FjyCtA2NF0lwt84myWyYLDlh3wiPLTxSU/XVNp6HqK1Na5fxL10
rV1xAsbiwicFVN9oFvXQyRsD6jHx7W78CsmAWzycziSF3ZrHFSQLFjRgTZcOf2GG
AK6406v3ZR19pA8cEuqwU7bHtAKppEq6SRJ0pQnbWoY+BfwSC/u4s5b/vJX3SDnY
dvnBetYWGW1p5CO3HDqLI159CJXHjw04zpm5VO8keWAa7cR2HZXzvj1CwEAU8bPs
UrgF1uU3iTo9oSX60BFTQ3k7JLZ9vdfBOlkwU9TsAWzOD8FE8NYWL4zx4sL3OPGr
wb9ADosMfF4ZTHPFCsPHOUGKylswULj5zVET4fajZMYFvhw+1OCDcBnq1JHN4HfS
oCN4GyEwtVB5JctWxnNAw4ecWLHbFdq3Qaq7gm1NQd37bOdhO+d9sITXMAvhKY/0
S6E73Dx4cP/yYHScytqg+dGIm5iUbJYSO69XyC832pDAYsRf9uKZguIPsYtAAhxu
7BEbi88IxBZ0eP9pSoxFuNWbk3EikpxmdfYRVg/bQgdX4vSI3E/+gQa3X1TPvqyT
wcXuQr6UyGJdgOu1r5FQkDLOLx6I/N4to2XOlUzrydjhr2V+PgEU46ifgvgwqEto
jo7HmxZcvNelTAw2PghRBkIN5enbmXA+dy++wATOaPc8JZcHPMUGOePU3hW31ORf
m/WXBHy6yIcC6qrKMft98y+RUsDQ5CMSARa/rESunVDRZp3mE3FluDpqaVeECvm/
cVsP3oSsj6B2FltVHVoLeVY6zUbJLkiU1zZrqqIZMIOe+TRMsHUHVJFfkrBq7pM5
IvXHElebMMAbDJsPWhOEXmJtaOjIZ3gWwVkhs8/CHJh0RhKH1ZN/wq+agge6GEXK
Sys9WjHQlOkrvLrPKd/nmUL+kVA4WqGTF78RG/d50VR4VIk7Nt/EXLFpOBxtbw0K
x9UoDNQ5t8huvuzHIlD0mOLRV0LVBUG0s8FR818O0nKXvClZkaIrf/ePbuLe+vCt
LJs3BvxfG0fwPDpn2ivxuc15EEwfbJSdUJnQCKxATimB2TonLToi+Uff9drqAlWe
sK/huV5mklF+x8agvOBc/+G4l93bhk6D8XmWJ2oxubReWPcpZqSEP+mZ2cznh/ni
iUhln5PDCKxHtdYilio1CfYSzxRFcs3QAUraqdBwl6l+A61mg52VB1gs6RqoYyV4
F/BPYu0jR90M+Z2gy26frKea2jvOrvmR01nDbiQqsjdymJjUhRCnri4ljr8UErc6
f8C9q6asONK/wJgx+v/ZlSFlFNo1V3tzgwXA1BeYXFc+c77a3Bdd5OkDiuQBWljt
URx6N4SFs/UrUF20gxcrS2dRoqXAaTBIvDvkB6elQ82zudMGIfsuFjXHsWs/1I7F
AKcHzvSUA+2rYuCvRrUKyF2UocVwNJsf/qgTFR+tyAGVfhfZTXZrCc6xLzJi+mpY
306RMowEdMyaXlsm1Aa7LXEdw2ky92YKaS2zV4PJyLH1fFjB2T1BwNibAoCVWLS9
GfWFtAwuny7eZEo58Utp3HIZTlCy5j6eUBovg4pMLd0lej/yMFiiEhEVOH1+gi8x
8RT+fbgxHIV39F2vDw1guXSCJEG/2TIdtitzg3Kku24MSo+Yep8ZPDptklQxEd1p
1gm38NOHXnMQqxTwZ8sQKeNgRczNJc92sVskHETN4BVZY7AVDDXRFUi7htft3/qt
XkAOG76M8kgyFZ7/QP4WIQmeyCxf93PRvmX/77AJMrUC+bxl9T7FA0V+AeAvr+uA
xGxAd3DeZjLbVCjTLcQpj8DIquACQAEFZEWX5hHptDxsyIaip4RoKAnpse79APWx
hzwG7mY65w2QdgGo7FnqSO+jkVKpmqrIvlgLiFW/CMhHslEsNVhxeRRt9k7k3U98
PFC9LweK1G+7G3pAKah9vcxNInRuPZbdhijmUVBRoHww096CLic9LJm9nMwczs9D
dSBfDXWGzSukyIKh7cWeo49us8+ycQSxlDvcF9kruyad/ZMCHt9ZYPpxMt+eZSTH
UMB2B0dDIxy4byrOLtX57SiWfWHDba9ROCNy4RV12xXCCqISYYTfSTSrJ1qj+kCy
RxC/5ZhuEfkuoEP+aZiwnnmFFfeZNBXwuHGGiee80sdKZVjv81JXpc+QTXd2XNyd
AWIiwXJKWwR00zfEa776AP3eI17JGzlwpvMLYR8pJJuqluwJxqZ80q15ef+1Ov23
aGp+k26hNraEifREwI0pjaJYNGzsAWalUcUDjLhBUFYO1AF87yXuFStRD3v+AIbq
Saaj0bL5ktxKn8YtMgrA5rXisdQoQxIvXEotEBUjSyMarCxO2XFOvUCH/5lLHT9x
uT83SX77qHStwtZJuIWImfeRk/muRbxwBQsggAfAoD9v5G2oI7M/KpvFEDoyBmqj
q8VtaBgUNAlv+LLMWxfAAmuURVpjxT78PK0EgXDzveJpui6qguLggTXnTe3kXiZw
6fV9O595vFyE90cIjcvMFIqeh8FW6Tf09HlvUz4FVFuAczrygAPTn3bcJeWqrQX6
dIaUaDif0XguAg9He1+iSjxOq+eDUNEqGL8NzZJR8U9cw7yjBrfNe0qV7UTPAdP0
rn/fU+14bGQ0gt4YG8eAnyPkdAKfSn0pLa8itbpFPxWISIIdYL14YHsNH54B5uNZ
nBjVcP2Xf6vnV5p7UTyJahyopjMJaH6vWBguTuEXpAaNESSdYTXwCExBsR8S8y/n
sy6uM0Bjomk+n321hHBM6bXs3Uoh1ZfO+59rQT8n95nkcujbvbsMGKKdfyrg33yM
aHpKrlWV3OrFiKVxlQtctPdinQUjyfgiNVQ8cBbvYdB+M3gcJdTjx9yg/35HfAlB
G27TxPW2jndyyMn9haBsUQkLMCeoDdTW6VtIOgUqg9ox2Ty+IgKZ3M47Y1oGy44J
LY663p/YtXLfEZ+VuxVhsQS6IvTHmaAtYq1x2WCgtBbDzZQia4E6GsKH27MRqVua
3fLTBlSLVlEvR9PCyCkV0rlR59X3p+3Vpx6VWyw6X6OYpxTMupx2j0t9OfEINbRW
883pIAc0eXkfVCr1tu2CuEdsAl/xzwgrETLFntCgHk3h8XZdheVPkzHXL6TLRyaf
iQsGh08YsI9+pYka9I/BHYnneFAQ7tqOXAb+1UzdnTBAee3rBAZucoY2XTzp5s0W
bMmok9ftOjhIIpjjv9Rb4jab2syl8VKriMPSjimlXtET1FYHTsxaQ6ZUpC64qSXF
keXL8ncxPgVKgYlP0ofed60rvcYiF8dNnZPob/FRRv7mR+pGdYd8GvxvfFhpykDy
pI+cLSkQnGsEEG7oOaO18zn10pfyZtJU3W7yn/1Rh4Ul8GQpkaEDM53ICVqgShr4
E/iLXEZZpYiA/pIZuQGHn5/S+D5X+SDBNCqqCmkLz0Y2VHqxzW9tIKfiuFpx7mwh
NUK1GP9KOGJAV9AynTclkOMV3+kyaB3uohQUv0Otv+i9IEfSx1xggxnAzIa4pxZ8
GhmZG0iXScIYqr6cVnptOdAHx11Z3j2LZ30A3uC1ldPNv97potjBv+T2BsMYREi8
Tii0es1WL1h/m2sLSEVu5VlFtGN0Y/dmLkvdrxfM1qVNMu0xZ4YX/d535fZh8mAy
AC5WYooR6NPcO+rmjhwlcLKv7xsRYZY9AJzHeCxo1U4A8cw320dz8qVoCQMtULzq
BQeabB4WIOQ/Zx9AH4KSCdLxrgJOmo4Td/p1/qSLeHOyl0afVn8sZltXC0ahwSe6
rZ38Wmp1Ec7KarOetrzieGo+fO7N6A1j/S0Z0FGUKrJ8ww2/xo3uyQRsoK73jeY9
OtMEpEpHmHy1wovygJ2v7sLejQ6TULBMQNXTqn2JhnrSQohE3FFKR1AJa9XjjFjU
1jsFPIEw/xESktvt3bu55q4beNPeVUus478lQFidEUfaUgNnREOfdzdrrvpS3oQb
OsKBCbpSRI0onnteqEf96jiaEayaSZuPpaO/QNvjP++lAwNUbZFzmscfMzlOkHVH
aAtRat2aIxZYf+zo2ggR0+hbFcO8hSN9O8nWY9zNyntZIbgiqZf+bqyyRupEfI5O
bBLjL9e+JoSqpUDIayh2bn9iAvgCvPTYypYEmEX30Cp1K9pqc/i0V3VOWmaAe4c4
0x3WzJir8RMZOHBkYH8yzdM0KkIAc9kgDmhLC0uKjdT+AsCIYbAXH3qMiR5ch2is
qvXXtrOVjnxPI3u9uqo1n3zU7LMpiDkDjTIzpBqMJSfAl+YdySUOYLVhha/eEcfJ
bah72M4omXNlx90GReL12mHWwo+vlQDSel/CZb3s6My8sUKewAAXGihPQug3owyO
iLeEhwIi5dbdsvQbnwfrODQgZh4/wWzl8R/WET2CP6WaODVbFYnUJp5Tg8RYjZR0
2iDfpquRKjD6jwAtpkvFnhanlnWbqt3EzyJFI18V+uXsSiUbqTVItbwoK7I0FSWM
xeMZJutHOUc2hVXL45K8qBu6Iu0WoD99pN9DQqbj/PhFXnWMsoBQkGoWXur1ktIW
z5VfLIUCtmrPDBJVadJdm/3yawyp0m/aFkrfhlQ9EhI9+ge1qeT3PxCVmC+YX8r9
CXmZ11cdm17G4qMg9IG3L4TN7wKUgvxxjZH0SbTPKNwy8CtmYRbBdGMpRWrHnYbl
vKTRmIgN7t45ZVuyyNse3rbznkxmUV9bOZ8zy4nex/uSb4LMXYBT20em1Pfnleu3
u7VkljBUfwUVRG/fZbs4VynFkgrZLnqNE0QWIQ46was7/2elulPP3k6Mm+u+vn0J
c3+sKjeJzmAHWcQ5yA8X4I437iHfK8Xq8TbDgVqro7qO2gC2JF3dpyXKgPjiBcWV
VefrWHQG0EVoC3bwunDeZlsfN81YGhGX+d5A4WYSt5YfBjeqDbWU8BxjI6fte2cd
PNQFAHr0JXFsFDeWU0ZkMZ1EZ/RJtAAju2nzc4zSPkXc1Wo3IUgCPEVYFTkj1m5D
YRdsNbthqC1FJZ/4anyrz8o3kXFKLDZ0olhkC0i2IFtGWqMoQe81/C2TXmZG1OKF
wTK5Ttm7zIFQ+BjOWegXPS1JgOJC4HfCU4JNICiaPJJ6hnd3MeUemyAFFRgzXBiq
D9GrhRM/FHvdZTZ3OAO+KwI9xViOMBY32H6GcCUVEiEX0bGrSAyeiuxcj9WL+6pg
0zDEa74TV98DMyXEqaU46DWLsYbbLOk5wxt6mS/MwkhUzsnZzxBGqldOeOlF53d2
s47s5LfLGyYWAV5BfAY80OVP9ch2r3Y3K+Vpu9mz8hVYSSqEu4TOX2UdEE7j0f03
PwIn29iDei31/F+x1HGKo8O3tmLdsWdZp+mvWrDlg1OZUmO3thbHlvuEytDj29ZK
z5+pibKzKTDM9CJMxjS91tMl7LY8gkRZS6Dp3DdXRgVBz0mZTOyY650uwrsUyIAS
r3QjarS2Hu9xOv8puXfqNEZn86BVrn8vML0V2Q+7tZKMrhoOGZfOaOLAkwdc+LUo
IjkfafUyWFxhaceMr/9zudnoEBRIJWnuN0yFNnUdXfEarz8I79VVXiBebxuLglnJ
Lj0DTZLk/3lcl2Lvi2OIv4YebqzB/MhMi5rdcXDrElMAJXD6jO0+s5AE3G4T9qm0
tmql79srDC5fq+uMUfSfQI76Eyl6c6sfecgbCwgvuqEMlTighpr+KlD+1CQPjimj
Sn435HOrEr7XQYijzSaQ7OLuWcRnIe9hLA50GmZChZKZBDQwCkut/hOnB0vv4mJU
SqTY0g+ygrPZzUM9j4aiNra/492YmiHRKRsoafgr7Wxb4cKb1RzJt5RXyMgfQD6f
LQAr1Us+JGKr/10YdKLCQaD84z8OidnMKlJuIrXhG5c3alHas2gPFMKwELqGH8es
rMrRZF7v7e0Rex/amNJ5UiQ5glURZcKHWDkJnAmr6m14Et5LPhQ3qnDrkLOMA6oA
HoKfn9tiu6C5CxlxxmtUKMWA8jvaOWkIKl6ws3gpA/jlX+kbHT750QP48rddptPc
kDc0Z/qVEpBwl/VkHw9r2Djl2KA0sN3ExiOUM/8DMYkTaDgcJljdYilUUU5lF+u3
iEZRFwAjUIY9suY/FQsJi9HQQnhfU3r34TrCweWHxLSV4j0wLDYkJilvaBK39kcM
praMZTRNTEIDMzuJXxSCgJ90rTtN/3Vsr7g7YaZ21HlNCF4Tcm/lDYg0iolychWB
tUpatxgXhdRAsUMuiB37oux4vkYBLv2uqWQYn7qifNs7COp//Cowy0PATuSaI3UN
dCStzPH2q+TEOeGfs04RMK5FMqcu+leuVoC8gWsueOT0699LWM3MZ89UkD1rGqao
xKhaRN8hd/qggLsHjzICpktsOqcWC19m+O49IbRytARHkIc+0X6xXMlptA9yK0TN
XuTBMhsWICxP7q2e+nsiWaE1mj9s1RdaQMJR+SBVZRE6dPy+R93ZBZxta5uj+W9l
nMvDG6PYLSc7UorY2ODnFRaIMVMTKUxjir4duRoBLqDV6Pxw0R1mtz8InzaOhbb9
4G9rHOzo51JCWcCZHK2X/XL8BLuez65/GWQvihAHLbpkPiJMGatb7yITqY1w9bb/
tU4owp37JvX51V1DX/l4ebBZW5zfv+oI4ZiK5SP7+Ccqx47fhX3t/t9Dytg/IVZF
XjtoFFXKvtKyWg6PTSpODx7g2EQ/ZeG2Rv1yzMhMW/95l6PqXykVIpzQkT+25BAx
1QaV/1jg9e6hiexWpexlmy9QKYHdthdJ7Vh0rS3F37tFHvu/cvjLZxUL+xDrCgdv
A50g8EtMUkmCthO2q7CSWGrX1aYsN51Gw5PXP8OWszjUYpYN/Fz9seUSlJP3EgRG
N5LtSI2LhSK62arqFD021/y6texRIdf2Ry2JNLPjqiXdYJVXi3z9XRBR8mMZobmh
u02vCaJxANjjR3n4FMPvyCM/eGoIQreO5xdH3uwHCSyK/J3P1gQRxjg6yKZoMwOx
sPJW+bCbyOoSkOeH5NlKtuXJvDaXHhBHScqruiBzK8xzDRtFk4JCGG/Xy6HDFjkk
uaIdNaH7VsQUNS3lUx4z6MWYdK+xym55xAf02XVsBMJOFaaSZihp2nTd7OFFDmqL
TC9QYYAmQoQk3yYNUbcXKl5aIRfQ8ILLjirsTy4Imm9jLh9WBk2N/VU9joBgs5yL
hxWoJxLCqAc7NsGq542hOrv9kBWNqn9+vslK2JNC08fmHHjymZ0EiZCrHKdq2OAK
WA830fzzvb01ot0BBOo+4uQRqAHPAsTe/0EuqaGu7NOAxslwSpRUfM/aP8XO46zq
0pvPmOU6NS7WJxqP/ITesO1i4TmBfFB5pB4MqxxYnk9x1PzasvGlnUeiq/1o+ggA
YsGmX23WdEnuDL2FgMTJ3kXRDH2HTERgoaFDBebT4OJ2y6fu1dK3yVPUyXT1XluP
yfk3Uo56i75tKepZWp5OpwXPPGRycvRTKswyuV/Qwnif4xs7GTXlN0IMN8subMcM
lJi0mLQybukvO8FO6hdXvebAV0SoOgFYOAgrHPFcO+cjr9/1IMazCpnBYkuo/mOL
o44rniobZ+zKm23r7HGjeF/5dWsTTB/smq2/PuoMrKoQ8YdW+WatG2pVsg/VeLFo
jDr8wugizyIbNE1wZQdEsjtO5C337YXyX77rddzI3UMC1g2H7U2kok5d/1rFRNBX
kOqUcRi3VxhmFzfVJt2qpKpJRMJETdA5vuXX/MwVkAHrEiR7vuK77bG2I3ly6xeH
tCgjJ7UiXCA6uOAF444YGvmlLKEtbJqbRcdnYClE3hb5xty+6vufX+e847jQG4Xt
Y54hZ6JRRQxEq9id6Ww/rEGg1p6LP5IY9YNVYvUdNGuuAyfXJ4q/2jXZjzgNKHRu
ruP/UmvVeSesxurlcr/biC5/iCcTjYORHBvsgTfHENfJyl/JzsDSR8LT75bOlxkN
Yjs8ThRnlq3H7LiPofNX1fWxW4e3JnCalsDkQq+q9YGUWT3TbGiQYQp7PwIKhYRQ
N1/mR7lEIoHNKpSVrLQ+B2Qg3/tmy5qqALZFFhnRXmrgWs/xJVVqI+sKcV8VSDXH
hl0638kEJuDW6KsHJdEiy0D59EdGm03AGT5kFzgsezP1Cep00+VWqjiMx839ce9q
nHxKeWSDe3RCckFE41aSA6zkyY1W3EKbO3LmTtLU8+ErDfpRJK7h5ngGbrGDykA7
Gyu+ZqCIYJffefWjvwnqbvtjYRzWdBTwvw3KGxo57UE6b0YkOg0bbj6vHeNPhbSr
4kI6glVb6Q/1PxmfIyFIRaxyswNTW+5K66r9EpDiHHsBlmtr/8l01lr0dsiWjMip
EtMFW25lZm4bYSIkxCVyqw1BsWBNbhNZ+EyVSazJPJKdAo2hicMoIssVoYXg5gQV
Q7ycOI1H/q2xObZUtY/kir2olJ9S7Hl1mXY2RdBDBx4lgg2GCm8h7F2vqh8/FRIe
6LgvojDxhWe441lxGUUlRI2a7AY15BcXmdeNbKroO+xL8oDSAZ0qMuE2tFwIn5dH
PBQwOVrkPeLZRHgnYCpG1TeHz+H7qbSS5lNUWmBZmpcvZfNC+jiKeJyWQrEpHpkE
hP9Ol535oyFKY4H3E2jvRgNRXkoF8e5ERstaDnAIyRAinkPU/2m324vWPm/pGo+E
s7Oh5O9kEX5Eg3NXe6Iu2q4sWRd/5jOSZiig2e07dnK8pgqido9cGWiRJg0mvTAP
pIjcwld3iS1A4HsvPKd3hvi8Vf19p4hvAkIpQARrjEpkIKLekASlX1yfI/bKZxMD
G7yzNREYgbFkGZIcoazgYzPj5Ob3GrZYbvsUmf4P0TM/L0KMf2yK7y0jmZd3++Mt
0bguI1qQe4orMmC6FX3u1496raJUSmYC8L31babnnEmeZg3Xa68SFNGwrlCh5jrW
trswU0v4RNv0cqgFIGrh69nHB4axW43TSr2FJtfRVc8pTdIcG7w+eOJXfC7RPPal
RcpUsP5jS38AlCwEIQUWK+gbZP2fqelb+9Z/dKUAC73xQikZ74IDU7x4BnJTBiyz
lOV5PLEFUDQcWwH56Qd9Ij1ollTN7gW4LKXHxwcZQVid7E1jPdgrw9RMFFF1shtt
VdbREqwjFOt80xpXcuQFvPcEhorxt5NvVISG0eoVLysLsMYSnRlQI1kF341N9j6e
iNjbJCUtJdHMGc2yryH6bNuNZ9j3NHnKxMYdo5HRrTCHQfhcv+f83GjiE2fYdchp
3zIxmfvV3n36JgDVmqiuB2KMtpOKqVvPaW73O5FzR8fW3gBa68ILfb4VqaXeXank
P6VuCNv4dzBg1EhbbcPIkz1g6feuhT4L137M1udFWO6bcJJS7m7wUHJpB6Aj+9ql
UOWqPS6CvDKOSoogLfi9dyvD01TAFlvSkFzCiOR33IbA6aBoIvxHUISutFTaRcSB
P29i/veA8cUA83B2waPVl/bvhbBomT4Vb9PnlXwx4dFM5Ynd3jDPhitKPcgHXeA3
3wYBXjX/YLZpbtuXrs2kRrBoBOhXY9T4WWeAeOUfoFnLRjSjQ/+gqQ9IQHy/2BYy
dfoJmg3ZC/vBovqbDcwz2XPhxro8asO26PcjBVMiv7W+sC7W0NAt+epKnEktEZju
Fo44ox3UkjCdjEesZTSx5KHHGdN1xJtJAhfSDoztgUd3yFdGpE0SV82Pvd8qknTW
9yJ/G8UqBwtsW+OgnltifcZmWTodi6IM90KuphxVWHTP/RUNjOL35/FRSEsv1GLG
lBvIUqu4sHMcKjJnS4YnBkumq28rG6Ieqb3gpr7EZ06sxO2jGiMytJvzFrmMpJ8e
LjCPFyi5lJo3+k+x8iA50gtfSrokgb2qxnzVJYnBUFrlRzHWfeiOTmdZASL6A+ap
tiAcqItR09MRUcMq504wm3gMQAzIRa5y45iSoyuak0p/9+GXhryXY3m+RmB8fBmt
V1V+4RbGp/SKsKJEKqZAjAhoGsWec0MTr+EOiXznqqAFzJOIYharVCQ122VR91Ht
s8FsbsLbmTKmZ8IJQxjlpkKa3n90iGM+74377+39KDs4XwrtDxqTeavp4WhCExrP
vFEUFyDBEBMZ2iRgDvM03e6SXmWB4rNUHapQjabG6BoySwfZjBy5nXyrJ8ALvtJ5
3K2UZ2t2KA0frc6A6JsWLOcSXAfkT22+koE/bWtaf+BQF4ZvCgQI4fH9KX/IpwO8
qz4YFqFfUtvkuBvcbOOva0UFMSqrTQNPvH4D2k45Rtle58ONJPgZ6qVBKYPZsPoa
7ssGmnY5Aup/wAN6hLS4eakrn39+Une8u1CJModHoxyB8Sb9ZNy2Pjd/cEByRszd
odwkf2d2Qifs7THn8GYL/C4qyslDwqmaZOOX9jmCPOcerfDF5G4vptnuHatZX5Wc
wZDhmUR6OoH1Mvw2JwNEvzE1fLBhY8xMMdGS8bGo0lVlIQOKXqgjLO+4XtYWrhCg
95e47kIFjM9E4VTdkfv7kb7tpNnsirKu6Hk6vorhq0jEonet8bTV+cScG3Kep5Ue
nS7YnLKBd/oXRBL9/LZFMgpnY56nfP3sXHf8Okbv6Kx60QVS60ynblbj0dO6BTcL
ghCs5KzUp1056t1yviZCZz/bywDGQNpQy6K6egLLn3DsJVMZfyJfYGCMJsQLtIKu
rl6HI5DTfZPsl09YKd3AXNUd8uFrcl9mhW/PidL0TuoxFf1aU5942V3O84ZDEe2r
LvZFSazWSAM/x2xRvzWT4pCS9Im0h4RsP23IaqRl+ONcSjztSZgbJlT0Et1tCAtz
gZ8acE6Gbkqr+a3rsHRveGeg5elmvPkivstCjNUFBhL+psVJdQO2MxtP6Jpe0gCy
SCqTDcbmf+gGhNa6fKwoqF2OF4TF1IxK1gSUEHP3DMdssvwskPHXnJM7l3cBo4e5
cCf8lgipeM5IQJHOsds2OjeO3uthcZyb4U4kXqoVCfVr2SALzhyMNgf0WbbJ1Gjz
0PCba97YDwXGTHC/XXWLRRO+9MIlEXSgScMJmxHx0IqQyak9Fx2ukrN1028hmoXE
hjj9XMc+2/zS1tgDke0Sg3RvVkx2cmHcZe14iyHR8X/jNuWVbs0n45IyS32Es3gi
26koa7YYHTEGQyORpeJV2PR1NHJrWTQeiETyk8wLVeuSUFZq8WLVT2+5lw8E6YYs
Is86joEnavVU6LdWsUV243LB32/Iv5c3aaISx2aSx4/cAckLjqLyhTYMp7jmUcsh
31Vbr+Ikyu4+k1yEBCtn2LEPHo1eqaCtMKdXh+1CUAYhW9NBbn6he+avvRnNoj0S
er/R7wWyRQtnLjMCRcoZTbvElDUj1vOeUD8eMR201aLsnKXYUqgzLavmu6JDgW7Y
bQW73nQBZSK0NE2PF2J3SGqZAyyU05TqBeMeLiXlFNiGmj35Qp6B49LG90w/JJ3c
Unh52Pr1VXn2ROWB+9JzARxq0zytctsO8rZJxRKXtSY044V13sXqXL6gsTDhWcyd
A/mzd6I7N6yIB0gvn6zkjHUJXNcTOpcFYi9EqdUfFm25TA54z7bE7xEoi6zWqx1L
FBio26QfOnAWpLTEo4sYTMthb/V0f+TaeAicOPUi47a8fE+srUXu0IBl4Jj8oX3h
PTPzdjUp4APx/PrpVESYy46Glo0mQz7ipusVB6cFdKAICf+WjYbnBc34lg6vb5/v
WkTYB3oZc/QOCH0bWJuT/5+9RbPShksuzzsdK3r9GZk3DsODRNJmeSQZiKK+HP04
RbymAu7hCPWl2TS8jM1N18nr0MA5rxyfU/xWCw8xs5sm3UW7NF6eJ9Zyxgtmj3b7
6WOTUM8KENBNXh7uAinC/2+DF7+PovPs9P4k8LO5RCYjlBO/EJ/+uSncOGCQ7OdY
lvJPNNb9aepz7KajNOGTk3yd7cXszQ9uPS2ehFcqxW5Bf8xxJ6d6vEvVBqTj8Sl6
d7cePih9hz1aMtXBeDyfGO0JjmTWFPsYaMVkvHsIUcUFygh9o/g+waDCdoFXZcry
vXa64eofUuTXuUJQchvhS7CXPCvVF1HxGy9XAc1CGeB/HbsWymM2oTlKOYHfz2pY
oElG1yEHHpiUs0HdMUAlOecF4/awPV1YEvwhLwvCamnExoC4mLh3d1covyVzgn/7
iU8ZE/cPs7AamlejHu09bWHFracBlYj4ilwnJlk6sjLQOua0s5eMQUci3IRB3feL
ZtgP6uMsPmBH8sqIqqNjHpq9sVxaeZrqdd/hW35PBDjs74RJkoIFDmHqSn13Vyjy
083gg4dZR7YSyzx/TUb31yqeRT2UsM2yIvOfxiv5ydK1MpBvBcXmY/E5I4iEzPFr
vye8Ot9j+xICWc+QLeDLhXVnbTnPQ5ladV1XEZNBh1gWmxGNOJT52yjUZAmwK720
rHGFu+Nnk30/W2dSYZdFZl64EsCFo0Nv1FaInROWTXnfFnCjq8HvRZDSy31T5KQC
HvcaybVaKFOlRmN7+EX17NqM/jWWXRTBogS932V9dOuQfRiGK0Cwlesp/wnVjXpd
6a1ldyJlYHuUDrqLKSY1bQIFzmT4+HPbvJ0RwCuhwojfi/Ys3GTkTKQoLQsKJsKs
qTsWzB2EfRyN6q5oY4Qyl6NgIQXzTAX3IcjfrI0mo5GeQEjo1zmAz5pX4ndoy4Rb
WWgqe2k3ki3t6O5cbzXF6+xcU8uTSTF2h+CjZ5iFA/YkdbDp/3gR9A7p2aUNSAiv
dpfe40DV1MJFsImi/C1/CcZL/mJwb3+NmAMBCyJk21WTNDUpTI7T17Ib3vV85/nW
G4gX3cKMB5VzbzWZFFms2Zclihl5AMX9DBGvhhaqwcMRjfhSqrTY4YK4vfD/cr7A
svzi/1FormKAGvmk+w7LnZvp78XLEl9kEYcgiE8t/fRPY8YaexKs5MH8KtBLubXX
8aH+zOnkXPuug0pH/8pNXZb7QA9CqlUm1HrGlz5vcJII5QTsLtQeR4Qq9V5xJvpQ
nIyJwOogIMA5QY8Wp7V8U7VTsAOYWtrm2/80MzDOIg+GVIqH3wcsYrRwEChZPODN
jA3Hy5Sf2t7yV11yGt7mtCWYXv+Py6pe3IA7DBUgyaCMD+6Pb57JdILcHJG/WKPP
uK+dSQhDYKLd4Y8I/QwFOZJb/v1c2PFRQm4dd9mkKa+70QfBVekyuuDKWzO5IHwr
GGL1OVodrJERPiEGThUZPoQmtGuCro3nC2UUJ0NX1UAynczY0EExiByKvaSzwHQT
CMJTM7gjLJvtlEsm2u/1/MKtWlBfNbDJTQjVOfLNT/7iVQQD9CuA7afhx7aeCRQk
bnIFVdNbiDR4zB82BTzwqy0V91lhaLblOLlDD05MV6FQKtMa5PXKNg0t5S0IHyfv
eE+2KnWXqvSXQp0ZD9VwVg3C9ML7oxrKmSrfVmIJglP+EYKrH83pI7yPfOOrD/xM
jxKU3n1NLlUgwJwUxxNW6qd4C+xGs8xxJQ/tmeb2QpQmj7kwJm5veWXZu9fp8npL
a9C8kCrpBfNij5bVPvkTLdNDe6YyigkyvFay4sc+9QeOOAZEvtEwCRoG0OeYyuSu
WVP0ae4RItbtH1EOWDt4rDp9LkQuH2xlgdjPK1l5OWAh2O4m+x7iKf4GZBRGdOw+
73wCspzgxgyMMQegn/0NMuwAxQ0FNDYcgcoZ2u8NYb+8yMIzigezi/DssT2MPJGz
QMkMccNrRwsQDmekfkt+lJcgyQV3jwjnaYcV8h2gIAnEa63U8Gn4GNew2ZS1eVjW
jnWx9zN93Vtf0ptgN+RbdwFQvfvdPPXnBC6hve9Hv39ipzot0X4mLIzD8h4ivjyW
jvSC3XF+3TcjDJ6R/5TiPYGJE+VSlvrwsNHFZHTn0tqJFCUhqmlg69AeHDdordVt
aS7MiuhtECsCr8XOmi7Aq2X4UDXjQ1yV0qtXluNxNrXyfQueMYwV+L6azpjM8k9e
N25W62O3aKyGj98YR3biUoM/vj7VbXgWeSKrOo6uPuJaA+yRF4CoUK73kVe15xFf
0u58d4bUD3cb/CY95XFfIuKaqCh3OLeU1pA7Sd9oUTocvfFZreEX+L+/Pq0cxQKV
IxkbiGT/foh/MBCgHXVADAu1sm7O46i0LBYpoyHIK8WHhdKFk9Jzn1m+jNnGj8de
0gewGz8E85CNC9d9hLZPmaDnwsNMwDfsPXAvArUHGpKnsui0P+lpPHRZzruf0fdS
cne9fp4RmTFqKl5R0Aq4oNO+gSMd2wSb7Dep+6eX5WesVsU5yszTsTzJ4hCBupGr
soMtTntrGYNwO2sGtvSwPClnrhTHglk+3T7UQnWoK77iTsFTQrjPhn+pB9UpRVqi
0Io9tf9Wkrb5zbifiVIqu3JeYRAhlXmqaXhQh0MfSW1hcMuChoXx6ME7RljgIXig
WiFQwdA01JPNdT1VFHIxZRIs5mHj4BqObbRFmw+DGmHACGtnJUcXYgs1v67LAOEw
stePw7kaGQlcf8x1crppk6nCvRBa7eqNbfvSnai2KmB/nVsnSRwf1RohDTdVQdxo
l6jH7GOWRX/vxU8Fa/mJ9a0T73jwT//ASzEpTxpt3bo5LDT7hljMF6M/XxTCHkn2
Bzs6WKCnlgn+euK3mmH1Vz9BWqdFPYLDXmnuotBGIDQCfDEN764ycpE6J/vM0XK6
DIgpsEtD8s9IuanR1j40Qa1gNSF750FICyssjY1QnMZ4Rfn4LjP5YdpFZRQuvJU0
FiqkzwUMxZ2rwf2jyam5LlfP84BwAqnhlTpumXIG19MnhHRIw+3fFoQLPeZrCVlS
2vSphp4BMNMBzvJGa3ln6RcyaHrBNraEVKq2SaDMoTCt/HX9DM2P1JSwp1kPyHAy
82/h0IwoAJGuyaCSGB58ZUzX9g6wzDml4yAYrf5Un+8gvEkWdIwOJyQ2741FqqLw
1u4+pbRl/33sk08PhAp09dq3b7m2uV1+w6Snh0FUNB5lmbl03ErykbVaKCAeGvH8
IR1x2E4uTVgyNML9JMMLGk6n87X0PisICaa5fOBn7fT8bh2XERnkhWGJ0sntDkrh
1636F+k50QH6lPcH98RQTCmbn7Dbm7cLShaJBjYld+up/V3TAYSl1TxR9U1j9S6H
1uQBeoi9dSLL3hoLZlof5tDGHAhKasv3fBnL3+pfGg2coOGUqKR1B5nZFWaHFt57
9RIVf5p7oz6sckpvaQiZ9L2BOVVjTMayNKdNKLxHAb6Z715Ry2FJ+iNDLClt4fmX
dd+lawtHPzYhlZkHi1MjGYFgnxrr+utA0KtR8E3fXmZIM81HJYssLAqpZ6HGSynY
Prf/akFqRIjeEocJeS3m0w3m5KZAoKSfqc9FXXR3zOtJU2tM4SuC728g+kTGDcD/
/Qxg9BdNQBDplqWIMobw7Odto7sYPaVscxfFkNyIhX4915X5OT1ciQ+CCoDnx4Dl
IVsjepdHddVvgQ4qwH5/t82c12vXOpgcjBUvulbUFvdoS2ILlZyQ0qGssDPjLG9N
zWDcIA3Qkj2whQHV1OBw3n9ma7b590Gek+JpdFPKckfaaXhxiFZ7G3PIj4vPYEAT
GDPCsXYy7ia1SybcdwdkhO4lj5CsxiMJzAe/12YfNU/Sdu7YfohozF9ggNhSI7pX
0k9RQTYYam02atjbjQLSXFJwTp7akEHsqCJBo4fuhSJ+BlaK8NI+Myt0Iq7vxJXz
I5VxXiEQDZwwqdUVbH/a35vjMpyem4mtDUW4zEibcE9Eqd3IRf3lbsveMp+HP+Mq
ChPETrM/PkKXjQ8Kc7b1IuXAmzuQ5Ku16NFRTaiOo7lyO52GgMLSJh1an+YgcQxF
8jZ8nQHfQoz6GlAhMAPXTCtrBETzFmtBmt9r3bPL1lj/dSfHpHnxAxq5Y4O8XijE
7qf0EOniy+jJW45TT3lUQc61hkG1QUBKyJuMh2HmoeU/m5hYnI1FVVmuHMvdZ36a
2tgVGdivWIfkZx2TSjrWyOCQVhBShKdnt7gLpTjpbMMU44rWMs2XEaP9Tw3qZskf
KAgMVnW+qqmy7/urHIAbzoRddIjuHtbT4w6a68SlWJfjZGfrr3A2EkrupUAitL/p
oShFGDm7VgoGfkhypONF1aZjYQse6HF9/jL9YBRnp6DbDEJGv2n/aA00uWA21/eG
2YULDNYzU+AdIFrl5FXa8Idb6jxs90A3B9YCZqp1KWI9kJnlUCA3tdjhIlWgNAk8
mcgvQ9BVa6doNhUIjhx90h+vaa8ITmfJPlZ7QGfAZ5BdoEkR/7NEbVXZBsU4XJPQ
VaU57eZ5XoUsG5nGMO4rTHCI+7IJB5OjkkAcqlz9itWVdspMdn01CXaUT9VIaeQ/
Wy3nCoRt305j+OKqJUxdVs6e9XBBx/yyvQDYBBU9uqYhiytvXaA3GSmriMXMnit/
QbSucUHXxlKoCLlG0ZOAZHdtOYiLXBKB2WRxsZQOxc386EQf6pmJ3XXtPAOq0kt1
wW+lM9HNijg3dkT7Ne9q4JjaUyn7y+mDTvMP/ZMCTCiITr35C2dpkgki2O/wJBAG
ekOhp1eA5/wzyWCOlMSKrLhTaNhS2gADjeIAxqugiYbU2tYFRMTGPQQ8+WqEz67C
pSKk/vah8vd5IQzsPPX5pHB+wUNxVlF9YZ+se9TN9fGg8g62SFsFwW0IJAeJEibl
F1ihqgUxymoWgJ+qXeiuNQTVQl2eqfjnk1xF4uiRga7LQOtd3/RD/fhfF3cUWRFu
JXExhC275Ad+fM98N4aLtV1wFW6rAp5lonLaKYRdsiG9faS4Y3UmxNHEippvTdhN
xneExA7gelSbBna8dqDfmFTUO7p2J44Le50pKSUogi3R8mesT6Awc+bC3F689TIC
rhjA55uImfTw8H5b1B2MkD51y323gRgVT+xC53OnIY8fWR3aJUqyy5yorwFrfYUM
Byd7aieMMHb3aiNAWU5CsZWcvjjkIgaLrQlLK4JpK+qdtz84UlyGzcB36YqMI0s3
rzeKW9mjLgGeTFmRKSU/LEozU4Lx1mhCQefbXJI7tC6hhtZD6qYrqTOL4C9raTo/
e3IiiwquPXy90mPztiS0+XEM3NBDyoo2H8RHGDC7Rs8WBA5V9aFRSh+WgaMwXe/R
CKb0um4BT2FyXvYiK4oEaV+J3guuA2mc5sw7HuCtlxF/XahDnUWLKgcZ+a8ipodV
451t1In8nTCJqPAVL4h8oqvTOKyVAc7RwO1dT0GM+65eZ4OZsskRSbJE48X7Ts/D
6P3pDSb7WWpSq64JghTG36eCdt48G4drG6dTXmYRUQHcookya/wHv0F/YDqGAfk2
Jm10TpLxxYne1KkZvtzrIWvjcNYFdhPHiUgPknyxvJ5KI0ksx3Y49DxxpD7d4wqe
QlMNTSmeWGF3TwZUyBub8BwCguMQPrvFYsaGYwaxjECL8jrDFf8F6M71l9fhv5KD
tl8YFIQvL35W5TPvv9QH5CCL0rC3j15ZkXFX5B7pxbNadAjvtPRndslhbCYdZeDp
JAm8uchHkFJccsOOdSfevV8IEbBsDQ78TlRON9dC083dUnRUBMxm/monm8sVvXjJ
pCHXw8M2QKQwslLyTLHaMdfaRwXuXb2x/X4aSPlcgKxtfE+SxPhgZpYjThognOPn
CqFuhsYg2yRHt1Zee+2JiRjQRzOiAqkjM3FH37cGgm3vb32rE5dv1NdeyRq1HoWa
SxV2020s6j9JisNWiSEeM6i0Lymzycsj+hMnMMes1Bh0fX9E9kVR4V1ow56+3/yY
bO2Bz6ZWGDPSURchyT6Q+AVrF/vUvsWH2g8O23NpqOXvbnaGaxP0W7u1KDIk521e
if1+hI2XKqF7Qp4XmbRow+n7lbRmGjlRaA+sMK9U+lWbdmWhxqHNCGRR4KK9b8co
FFbR0HXFnuDgf8a6yOjB6ybSWQKggaG9OP/V/78WPG+7QrkgJYSc9yN7gkpcVSdD
+2md5rtiFLNPHgd4rbpLmrzZZfMkIUuP7mieXtG/tYfzbLXQ66FVFSe+Y7hHnjCu
FD+2/noxGwhCfLVWHNntvhaqoGAeQY6hq7faJuiEUgxwwy/dAv+MnfdgqJUl3zkX
6Cu0WcfEQrP4ITvyuCC27pVWhCoPL0efyt3iIm7vFYjb3Mpsgh+4rQrznPih1pFj
rPsfASQ2JOzJNB023khQwYAycNm/S2qZmyoRLJfs5+mzI3gNKXiqqlx/m/7b+tez
S2/fahX66GLl0wv1q8gVindxDiAysYBwqU4jH2CrqXnuLDrkto8gnLuvT0qLyXyj
AQb2tAFhEwzj4MelYt/c3FoDVVxR8VtRaex7G55ucTAaK9xeG7HWguAKdJzAaXWz
wjcJE7w41qq3cR5EQDBIP710hqT75vlS9kDOwQwvq5JJZpcgj5rj0T5rH0GwRw/j
vBxyP4HFFnNzC5M0A8xAxUPd/CBy5Qx6oe6qeURzwP4zCM1WKtzByNuLRcCZiYxR
8eyx3FigG91ooccpsUObElt07yY5v8Tiwgvrhfbi5eWM5HwXKg892HOkBVLSPyoE
+s1FPcw0jpnOYv6bAyF3VeWkqw4V8dJ2UIatCIMeuaZGW/4nKf8HdKllVc3/JRiY
KCtIl9k78bKv8FFY/offhf4eOXSeurTSycssPb+dgBK3OvS3UCYNXFK6E42z99Gk
Ps0XyyC3Ln1EPMKuDJlyQ5FdW6v8By99SLN2NcLBDDav9bEgF6OhofB9V8c6XG0H
CmdYDDaaZDNiApiQ01kbdKK8ErKitUNqzrVtDIQ6M1HaLeg9KkpSQvtb2WBcgNUJ
McxBSEN9Iwlqn6AaRr+BhvbLuJzlDH0x0woGT+R0dpov4xB+g2ZQEJXIy2Z5t0sc
iEfwk49P1zmLpR2iHh85XF7tF9WhUYL/1o9SMVvkgOdDjfKb9BNZIVIVWAUGc0QE
eG0aJqpekCxJwDLUQG7hy2ogTJ/Amg4Ithm3cZSH242yf8WvwotViPG6NFJC7tph
j71vXUBmLljnEJ1N7RXIgcG90aJdbapH/wn7QolWL/wvUcyy3msPTwgnujEq7EyF
fp5vaXnwKVSdwWcWXek4iwUWQ97qByBDtMgkhAbn91wJjgYTleJKhlnhay+pudV6
Km8cya1n2rDCKnZ/FbDm76MykAFf5fNpzSws9NrC//YI9vSUJ5GVIAxn+fGXpyNE
2b8lt0nSJKUiIf9oEJblyJTdHyDtPcC1myTg6JGZrJbx7sumzDHD/cpk5XNHGwWt
BGJ+HD60iShros2+QnXDqHWZ6kU8+vDMUCMLWKi/zzFbmHEZqN+/nhYEDZKiqLJD
NCgDi48MYVHgzsYr2LRfkcv/QlVmgY6mm0uBFkCRVdotCHXrH97pheX8bk8XUlPx
yjQxd8wPYK8zDAI2DljaUJ1hpLvq9N/ED7U6fwXsP/moJI/3oS3ncLYZgnPIXO4Y
eJRXEkHMakpSlSIsuv09sN3ufpDiSYH6qtGEEylm5mfBz2W42P3D9PT81wm9OpcD
R2YWZ2w7fwYI7moGxLIi57RkWP2aQg6p7F7omoJ7czcafj/oJ9hMZyioVVpqGFhw
qeYzc7nuDndR6XyfLhV52wqdwE1bUdZovdsskpBHDryW7IiK8bHh+MnYK4YBCJ0D
1Nl1SGXjCtjnyKpu0y5G89ARhqJfjNwoaxExSZ1Nr6X8ktjVTVvn3cbNh8igutg0
lA7I8qkY2IxncRxY9WW4j3l6A6+2ChWPNu7nGL7/GdeysMrEGgh2bWOPZYUapvRo
FHV7oo7V5JvVOaC1uH7CdnzBMhBWllPBbJOwiAJJx+POeqY+GoFceUG/Y/aIGtjH
7lquTdu5h4owKm4D2y4YPqJ+IYWc2b3SfhTHg4qz7QxCA1iWwPHRvlHdlhZy9g5v
2ZJSJJdlNLcmjsw8qvt+3cUbgtXQ7o0cbOFkKjXtig5y6E2vBc6WI0wN/R4VJO7S
Mdslmr2PA8ubk00roDKpL+gId4Cv3U/b2KrMTW/N12TQWMmRgw3Yjz9pP89NRIxj
e954KHZEs0LqCV8B2HclENQeP9KyqnaTEeh58+PwsWtiCu+u2s0oj1trPEgLw+pQ
7yRwgFHY3Mgmin7eg9ZSpGfGDcq7iuEKD9n07RXFjxxEs4YdscxrfnuYPh2BA4H5
myqVMFkfesXrKAcQKsjoImNpdp7q4KD8PWTVnqWYybDGyvHay8C40TGqP/NdP9HA
w1vkKnqcDR32QZAe5txYYsnRY6uizTrlAPkm1G3BGcDoL1BcEnhS/NvCcpr4J6G5
XtbLtstJKQywTkvKO4KHG/P0SSfd+6myU/C/mXKG5O3rmf7AfazO2j/Hh8LfErif
9EZQUT1Ovfdbe78NnW+qqYIyFCq7GhnpsPF7s+A7nGgTfd0CEYb5ccpxsrAZtf6t
uQhAf9RbINtYOnb+vspMZptRW0uzkbbFm3eHm/uyCb2tALeDXg4LTYs8huKBsyBN
7fxgFGW/iEbl3ThFz6+GCoMg6VetLgcRTh80Yd5B4ODPTMekm6pbumUHmpCS9XRL
2xJS56Iu1DEJaW8CZClYIPHSCCQimzmcHIGAN133GRG7Rtp6oe1ER4a/wOc3AF70
3Yxfc7LrU06n7JMfsj0LCoIhQpY48MD6/Ne+hGYTvfCBTTu0KsGFwgu60AMLPbqI
WWEcHKcwudQmax7KsU5TFp8ysxyR5GGUc/FVkLMeJkzL1+YK189YP/phnuCfbpZ8
bflZmTrCrlTeNk+vetq8FmE49Rg+OyoO7oPOoY6zcAXhMfZp7qUpfle83/GYHzga
2q9uFiaxhsc1yaszRL90ot2+olU2iSuH1l0ZnEimIh/VXSAaCaofzXPSSBD4agaX
lpQVLGGEHRLWNYUJwkmVTDzXlKHvNJ5e3X+nUSptFk7dyel1MYtSFAYWZT8B9ZXV
FzzVCJ2+Xf0SpfYg0+QgJideYUlrK5dsUXmZEzGpC2X2U56/hfgbuaKn4EDUcp8i
Us+Seh5QeP/3IJd5Zc+YiUF5bDvb3RbsK+FZsD4sP+CyBNkaO45CTuL1Up0yJYdb
huzISKexSPRm2K/P3Qtn0ZCTroCsErlULVmtN8k5Sj6EvEgni+pjUua9bSpDLH8w
jXIffwuLH58vnjY9Aj62CPsU75DgYGkNwRxQ7R0Xrnj0t0+tUL9LS/fBST1zvzy4
j2qZamHo/NyFcYs62CnEPABl9zdIFl2Ib7fN117G/qHmxLabKhEI7bpLEfaqYEsS
mVHm3cww1XkVYch0y2tR10iUTnl8BVtXPGDBFfW1ucYFh0s95hC0l4sWpW19r/VU
wS/QlZ7fTg54dXPapldyhYQUQk7pCJ4BEUz2Aii5Y0ihRxUJJh2xkvWVtxQo30/1
H4xx7HQI5p0VOtCzikQ2Yb1Pj48G2dUVFexD1Hxflz5RjGVC62yisGfo3aNo4xnp
jRV/tmy67eIWMBIDxWMfVDbfMOFQUYKVlVJRZpM5Tdqu1RDf2xwJCr3sF4fjTeE7
kVy6C2+ka6AaeM5Rg17NO1BreEQa/ml2qWvZKwvZJ8lq3Dv3rUinBctnNXvhKSWc
lVc7e+XTlnAn4ZpZzmReV8V/SbedZUQdnU9awCzBPLm7SkrBKraiIr8SCO+vyN8f
l0rLsQls4/iFMitBrwoC6VjFjL3Td+Y3gTyPz3Da5DnFka96QlSTMB+Dv5TbcGYB
QNFz2kJxDbA4EE372YlLs5+yReS52IRIl4Wo3pNKMGJ6DrplllBAUi23/+fbXUXp
76E1e7iCYoX/Y1GOvPOG81otZ02/6HZSnlMUiVrSMI2oq36aEFbd/Q9wj3FBw7tu
1Gj85xPdTEWiKzghFwEDd0Mstw4ydkpz2b8ZYcuSsNhlIK8/dVomen4PXF5x/clb
RMOcc2vOK4bAcFZ3tkTbuQNfUhMMd4tV5lwnTPOrSg/x8hmVjFg2c65dXG5Iiypx
FR0TgpUzT2PQnUu8L7F9/fNH2KUdAl32PDLHzYqmLJAsVHjYpnRYCSFYxmamhYqP
aD8SmE+aZ33TStqLATkNhnHVApD5ZjxVZbNiayhbrpP3sBd96LOm81t4XnPXiYN0
vPOY5kYnliIK7lNhZElO21YPWGjuKn/XoZM9U1ObeTf3FhLYfhYuayqzX3owj7iT
O6faWu+rnfMUYIvNJwHM1at3gWEgak88lAeUt10/e8VCoi0Y2qzMry6qLAY1Rov2
9P8YpyQYtQO4dJOetGbv+UPivx74Ag5W0kMjlzlE/wSdc0c2ecMOD2U/uuK1atct
W3UO0+d59iOqcguM8Sko13V8/RMZtvtEPhqnXqPQEsr8pS/55AAMPhaqXFCqGHOb
NbapC/MbGUYxRgqpPloSd4ff28u7lh9RtMlz4FwToXHiTur0m7RYFsEjw6V45hUM
XiSOe14McrgrWF69l5W+c0Z1fgrcK8nKwBnQacQ59cxD6sX4V2Q+KkERCBGipq8V
n/tNsWRsDmtmvnXbrscV+addOB2PKqgSPeSjd/1m7Y8PqLyFfOmhaPQIPj0O0hCd
fMm5O4c5FbGhHMSvp9fKmYrICk/CnYeoCHasKJOHmQZ6wMWGBne8BwAymBR3SNBf
U6OVJP+6YXO2roANPOzN5PLAMXZCpZibYxI8JSulLSPpwNUuW4BKBoKV3Mme2Lpk
hdX7RbsPojKXzqQSLAYCB4D0MVj+8Nphe4nnuQRYgluiQT/zV1b0oslWnWIhFJR7
iM5Ij8gmMjAq+9QkLZNSUDOKFkErW2EUs895VcTce/oSuNfmVYBP/vD1l/AYuLGm
MFTjr577Ppryay2p0qyUcUgT7ahaxhTjcJuClQ7R6LlOVLXQzXQEyyTxgWtGKsC/
HoVm6qU4tmFpt6AeNlLlNWjjAiDkMfHG3befWiQSyeYJsb5XW7bShCSzFYxEGunY
1ACpswBB4pmkW3cdluhSzt/oOSNG7OJ5wtK+aYZCT1RK9HeA90oOTAyMB8+HcIA4
IyLxs7NAWJnaLhgldmOmv/391DDkPChLqPOWuJpqk793mjuwO6FpFgw1oCvi87Qe
f76lWnGearc4mO9wGgYXrXnoptc1tElKVFBXh2r1wCyd0aikZbppz5mCjKKjgPip
QAWctDm6xagjBbvJj3Hx2higgI9hq/VfuRskTQcpw8+LfJEeKpNvSUSxQKbW+Ry4
PtMeFVy6Qq0+mF7Uuf/mIelxhCpz0YqpXHmKQdhnhl+2o+kSrodudp76hftfRt4R
X72awUBYR/TuTlFk3Y61La73BVz9lKIOA8ofunXQet7P8h9ORT4ejTMW/rIvHA5t
QP+XYXMDTwk+749X8A4ZFEy/PC4TSZJoTKGXW6jYeHBBUOJGrc2odBJq5/9/WbC3
nO4bbMaVeGl96l/uPJPYRRLUlsGMZufMeBVtMeqEBTm92iH/PHkien8cXLForivN
UFMhwGxK5yVOTiMSbsc7b8lysrfejlwMA6im0dHsUdY09aOKRTw3MoO21RAIU0gU
nP5XDwoPCghbZH/10x9waUXhNZvg7o6JWc5PHPdIuLOWyXgTTwEaxtvSaoVYeSx4
jhWXsSyFPcPecClzRJ0GDH9m4t5sRzO1NrzwyhGK9zbw95zLA3SNMLF6ixAL5jm0
9yO388kUT4tpwtEGFH+Iq4dhfXe2YT5gaf2sattXYJZg+ZruCeBpCWLRviluComL
iWzH7wtOLi2GQE+rsHFwJizLWdI7+s8YzYF4/EkcPiHv3goAl6BSakjIyjcC2IWv
oS81sIWpn0R9VDgb+EtvtI1ENVLEx09dyooqJ3/CUXvg44emKGplyS2kyONiAENo
aUl4H2t0M/fSpWldTQ0Xm3AK5AoTKqj+dCrZnsZGM9iCoGLZ8BzJEKAZOyGJbWwO
d6lhBa7jqXwruWD2CRrqUSwRUV6UrO3AMue0SufrmvKCDKaiIPwSYdoFD7AzUfJh
urs3RaOHVc4vxx6pFfC0f6q/d+WKY0l9P4IIe90Ud5B15+lcvPlgQ2q6dEbWPIo2
p9V3/TP4mRkUQzhaRezxdXH9jzZJMZ42S1IZBmmsiLR2gaUOFCPicGGn8uQ7vmn7
laUdyEBo3u6ewH2v+t8hrE6gHYMorHjrRHR9T7ZranB4DHyVxrT2QaSUjbMgozDD
0yMcBOk/fhIFfGWL75vSdfU4IniUPoLv8Bhxjrv0zXSRHYVtHwNeVRQORrGCWEg6
ze/jtMCRl65/4jAQ257MnNcAfhc8qXwudp1FB20P6eQn7R9oyreoZlUs6hltTtlC
sVZ3Fdf/gETlg9Ubx0dizCgXLKRyoIKQhxE5kyb1AJjxwz/8xaNLEAvFVC6ccFmE
fLWflaYQDgyKXoCXs6dcVqXCjo3N8XgIrUeX7pRLEPqiG5FulbB4uBgchtR28s3w
zkdf8E/Rlknr4Iq6Aq05uVM6lA1/VQ5fkuEuu0+jtG7WKI3w/KPhGWnNrsIB5dEX
3L1KAoCcsfiULgkTRdgCfZRvfZ2z9bJUtm12wzTNie2sD3X5BiJPwdVUCOrT9TBu
x2oP/BgSV/u5bC0HZ+EXkain5OJA7e5rMHjldaSQbiuexsrEkmrDcNsL3t45MhD6
IAn04hG8BdL0kcd0Sbqf/Ul7lgXlAwBRT0+yvFwdOvh2TPQtLCGs+PmzRP/8/2C5
VAf0juxLZj6VXJHb8USQNZKKLtzLtgleLRe2eDibVbVsPDASH08vptRtoHdzXI3j
QiZHFpxHikn7by4bFwUddJi1cqA40HEXUgty1uejI5E12iiu8SBmv0U8Wm/4Zeh/
9cFvrJVBF8A6dSw2MQZCGdPCSsWw/IHOeJNXy8cMcti4JZZqxpk0MOeFpG+Fxt6r
1enIBVL27wch2hkayOZXkzv5MjrLsHWRRgEDKU0WmzXKG8kClplak7oBMSRrIMqd
EfBDJlKo5Jd/uE066psD8YUCzEMGMbPIwK1fw0LsAaerBuq3lAjkuN+bob0DcDkn
iam/ia12WJPeSC1nowa+5kEZHkdiLD6ifvDFiRL2MQOJqAImjjdg3rtKV6sIX4d0
xlwCdEWhnzLFEnysuA8Lsv6jgJdyNpRsnu7Zvb98e4cSGw4NCOkBzei3HGpX6KzI
WkcXUPNaMTo+IwuGITNnOA/zxrh6np6EBw3sCCeU5tWrKU0bTnH/FQ/7KlMEFHxm
wx2vD1FGcYOS/u3iZmJDTwhqF4QCtVNzgTsv98epsNfg+nUrDTraro7KVcymOohf
T3eLz6Xx5FUiI9GEIZt6rSmAcLyhfnRA8y+6sdPMVPNdy0icKX59MuZhpvjiJSXn
tsBGuNRNe1xoIq83CHc/9lQXFP649kcCKrOiR0aSY44uuGuLD5gotaAioYOHk/mJ
9K9furO1VkM/wrrXGnRY/oKQmg+ZtDdi8UqWSCEeyvuCqnudmxuodh3ZnXgGlfHA
Y0F5zq/y510MfgjGN1gw2Azy/idUeyFiXwz77pwkvK/tOsguNNSTvmdClxh8/Yuy
6bvBjfcBZj6CKa9Yu/UbZxz+7BQXCx8pJuEowQ1ncn+TQORd/kxWOBoyS0HgumrK
uSk+jrFRYaERWAGqkJpOW6DIm9EKnz7dFVyYtD/wkKpIGUUXZM3sitc1gN4NDir4
QXWYeMY6mwo3wY8yeELjGOa3QLXjOhpE4Ev3R4jJetdFc4VA4IyzfpOK1O2kzC4X
78uXg23AzkyyrSUDAMwna/3uRt31nPOzOoh5MdrMeE25Nv0BdJEOWf55mT5mKjre
q2kbpkLR0/tgtCxxWQAutcKzXGOsoMPieDQI3NWvZcGIZvyOXVqKtTWWlhtI7tyx
n2zjKRZT/0Zf8EwHDK+z6BYvYIa7oxKyPXKmUZWiCwbI7Om7I1j0QMYCw4qRZSGo
mtGG9Mdzf6dM6D97RsLaU17yIdSJmrvJcC2M/f7yHDrs/mFSKedMkR6brPSFocBx
+CKlAOXHfH/LvB0hGSriv6/4FcIOLqkSBZaoiDExYYhERPu5+NwEC8hhs490AC1L
ZLrFb7TkqXhCIOKG8DZQr17d9Ok8Srl0BnydKXjlN28cIQ6SNx/AeZlxaN5LUkGj
L6Cl4lDz1RQ3AZKSBAK21ocELTDipzKqCbU0/XCxRlQ8gDggYy/WmoQmfa52YF1w
bZOWMqqjrSq01EZhBBV7J5T9JesXPPt4UKbl2Zdm+vhr3deJVasptoim4E/B6dnX
6v83X83slulwxPYHowyMIfK74o/Mu7K3koEN1d0UGYw2+GaUUo8INwOEJ5YiCDtZ
DFJncgxG8h6BPaDvshvJgdX7tAM52InFcp3jyA6rOr1sMZfFMmAZOn/B0M4LKhBM
TS/K/h4JFWuYw3BiOyU18st+iypGEBAIFobvpF+GTSrcuq/sGeiocsY1+8a3hMD+
GSONjX2l1iRolkEvpJuwHbyPusJ7H2aG6oH1r7/kBMwQRMTWZqrCDvnecZzVEeJJ
j1gfuZC1Nq8tnvRuzvtegCsDpmtV0fu1dWiDYkHTrQC1nW+ak1wHaSALuUSs17pQ
EvvvSrxdabOJOep1RlC+6093SRJ461HE03E4s9ulrRX4HH5vIw3fMpW7JYD6EcSe
XTvBqwvzCoiHN8YMojPO1S3SXFiIGn5zm9c1aDAX0HqBPkQgI4bjF1T3HGt3Ocb6
IR/ZPQzV1AteDIhmzIiYQz+0Pb9ItBhEH+UYnDPxZRqQHCbzkS5Vdo3P6xlFm7LT
/hY3kUYQYSr0YkHyD7Nclszr6+mU0YYohm+XUq1D4xu98iL4XKJoCeH6xl4W94HH
kvRj8sSLASnglUFRd2/lD2pKSpMcLMz+/tFK9rry03LxyfdfF8XZFbUfvZwoD0UQ
tgjyJ/bENHy/D9KHP0Sx1QgnzcFAK8qPlhcOiw/p3gFoWKgJjZiftGvY6y6q1Iqm
dCTwXBLPaXzPE7ADLziqgJQ47oM874WzInzoarZsoEtRrxRypl7+0EqV1wfpC+ed
mE4mCBqx4msTzkByGxtcOum6B1gaT+MY0xL2+YpbpqcXQR23sheOjh3j/MKdWXyG
50eKSeMpcAGx81cflFFg2fOBC0z3wdxiI99PgxdjwAgmixGP+p9SyvwcD9yAEWE4
wCrp0NWozgpi32ETjyLQak+7cZrRj3QExhtBoCP5/+nrIywlsHq7g4uRZ21deskJ
uK7vfsPfsbiMysvWEzKYTHK89LbFWJ7Ee1gHBW7Gr3bXc5eFfjSSKoQZCck1K/g5
xPywDdqRvOPIMvdMEWDBdh8CAgOkDv5A05wVGXU6stEz9VA9D9PJS3J2EVYfmbwX
5ckU0jdekoFg1jsR8jT5jqFG9ilxGm05KcSnUCvZU9ljle3vV+xpcgtvoM5DrtxN
wOe4atqdCys5V1YQiFK1egBOVBN3lOlfEFYU0IBy7jJDFtyJl9IZFRGe0J5qc28Y
MEOjlBMfA/JRiCM2pB40Q3VosmI7rRr6EzTC7of0CSwBNdwqtAHoh6VPbomW3sbN
pHLA8maUynIs+3LZh0lSpeF7/E+UAHwh6yxwFSTYwkTo3K7UBeNW4Adnmzh4kNqD
SUJ4HMNkJeuDoTD6VSFbEsULcFokjnn9B7zTc1XgIvKr9EM30N0sCHiNMm1ljQmJ
91mXWJnzNmUuCAFdd1RH5aVnS+Y2gZGCefJURmOj/birTob0T7JA3t79rqz+Azz6
CEe0y3eT4SXsqTPyaogvAMWUorLRR/Cx6MjGrO3XSsWwcgy7pJfViQ3TTZ+kyIWd
FHUZbPFxo4JuPFCvIjgpxC6+k59bTf8hB11jpJShdp3UiGrsZ27LPMVaINUy7u/u
bdep1SKnX3S3Ddt1bPZ+oULX44ObNqhJxV7HP52lB84MxJ1+8SMv+1Iz5Az0XrKc
vupvGkVfz0AKhIoZk5OA0jF7kDQlzSESBBYWQuNZ9jVifZNnhWHHQyN2XEao/FuU
FIreoreGURxbbBkSpn7GSk8NlUNmCI+GiMqGTOBuxu8oaL22mRoT1Rz2j4BQDDtx
z7+KsBEC9ZqHWzuhewqAvjVBvwl22+BDcbvjkALYsWPdnYJQ+6Dy5oEeifT/YBlc
TQ95Vtv7F8LTkJCzzMqSRQ1roVJ/K9+ccAm8rHI63tZfWDDSHoYAGx5+ld6C2kik
ocUB1c+mL9DaONjXtEckfxfTfx4KDAY1ZiFub9bcE6Jrkc2RkwcOXdx5hzxdaRvy
CNHr704+NIVgG9eJrhl23L38NqzVUBTzudLpbGEu5US+eYLF8zny5Chk+KMfyS3n
mcVv6Igg7djQJr+PdgELj+lQY2zEZTEWbJCemfOgDiD8LD1KNaSjfOG41AG+gH1B
mPpNrpCQ1H7pUL5hQGO8t5xn9O4tQ4ztIeetsNyQ/WL2LiVFaocew+mqI/9qCbxO
WL8zVsTVdkMoA5G1xr5QeGK8ld2bMMeJCnHOISn/4KGNfY1QH23TNj1ItJDtu3UB
fjO0y8gcoX4zddihtwUJAhupEQWyQD//kZ/e7D0vTuLr+vauLnmTfk+ogiYLL0Z7
sFZm3/UENR/DPS5UTsueuCSsXamVEYWDLFyakphuju1q102Jr+oilL/aoNos0ESP
BymhbhJKrvturRCtXWtn04m3Qc1v5DgEGjtKVo5ObMg+8ykLSf3H3++Ny2EGgPde
atRMBdxxSpnXMFkkKzSRs3jQQXqBg3Ep62Fb4L02SI3FIFiMCTbINLmWR6bHTiEp
6/Bv3FFGafKqY5YOH7ImFGX76U0UKWGFJQ9DA2dRTDvp3AkPN6yxeHTZy7kqdVtH
i+hT6AJfrDjKvKQSVKJHSdpYjlFWvEL00h9zk4VDgLr+KHW3ZfiCMY9jrz9xhCIA
JVZqCNO8XfiYKxUccEp2uOTz6Xn3E7T1bZY8MZVJid8clkuT6ES8yeiwSxiFo8WP
u6evTmNkM7jBjDxByT+eWq4hiKoB1aWswNmT1BTh74X6M0ynzBj7lOlSFiSwRPfj
0hEiVhHEJtZ25wxqbt8fGd7HV4unNcY88ZP7y+jNtrCFMzTzQGGTTiTyp1sG8QB1
qNK8T1BFDQUiclmUnCvvU7Liej1eRbQy1/MS4v/qWxlNpygTbpxHtoI4qvSDhAcx
lbmemtyDIvC5TAK9c6OpWrpIIeFBg23+3/Q4/CDmfWK/vRjWDvlXcW7jRaA0R0Av
BLYzzl+UvuJeMBK/PzcW6yxesH9jfoD0dBy0l1F5gvymkRTECiE+1BJKtm53d+Rp
t6HSjLtlHEeHLCZ572XGQNkMPXF17FxsECWI1CHNTdYx7BJ+7DBvaVcgUyt9rrtv
oD2QhYJBqENeQaw+wyUbsM6nl2/uBhLlK/zvwXe4sEh6oYLHYXpbxC5zmrZXoBxY
45z7eYWbhSrgFKlbAHhlz9yOO4nY8yAb9kUKbLt+W4CkEUJc+L7YfDL+FVArket/
pqb5QUbRYBS2SPQsKU8twXIPqsF/LSPQJC1NWFabBf5mMyR2oyYHRqNmbflSMqFX
0iLhCn+pi9LrIiUjHoX1ZgljnI3jmxoKb/To7CEPZ2Ji+/bcYLi2Om8hWnLM+Ugk
Co084zjqKWGMAY88VT8Bnjf/OFRRrWxOyFrYNTnJI8XRLpuJE7Wo8ewdBTLKAHOg
OD2EQ3skmYsVkN5zUm1Wl2wv7eKBPDdnskalMkRd/Kf/pS7g27K28k0oGCxKbZvW
Q8uaGUF8gNK//fiAkvaEY0fTD4BOl2SYnz7zcWRm83JpFDvCwWl+WXSypOAvJOlk
t6QXFp9k/2emzWeLItaqk6fzhlOemOPuPCfRgaXkoK+x0uW7oTB7UlFlfYTCgEYj
XCJk4ymV39chaD3snC/4Eae/eK2ji/oDj0RpoXghi9RJOpBcxLMAoO99HS2xQHuD
cK6RDhzLTkGiC7zMoZciar/TynCJxsUD/ekTk4MU5sR0Rlz0ukQes4tbGNIc4aNz
HPGu3t7qKSCFao5g7F2G64sKcXWsUHQhg+8VzVIS9YtlGr1tdngcQHwQV6IK/nYy
1hOcxdCUR4BPT7/cvP2C6tkjYV6xbG+kLVJYDGbx05xMDUughaErnYeLN2Tv+bQX
HR/ONj84diPfnS7udgNjj8MJ9P8jDTHCzEXi0tQvu8IxY3HNF71fUxvpkCuKe4Kv
pndauSjLHcferPXMFHr8y/uw4pqey3G8cEr9QAREKbh5wUSRSKxj0C/bWAI/ZMcg
d4JoO9KFwy/HHG+Ms/3A0QrC3Cw8Uyue+CJkbH67n1IORpWsiW4xqG0vxtmXnwbL
QjeIg/+SEviSyQTN+6tc1xXuIlwSO31JES8lhN1t7PO/2jqtbDCboq7ALMc9raDm
lxYl2+SJ5MXDXwhBc9DHuwWDFFpS5qkAWYfa4VW7aRGaFa5A3VLL7SzFBk6F+One
5lnUNlv8Tz9VPnXVbrEuImyztk5fL97wdhSMusQzFNC1BnNBmJbYQPmWaJwZyKoy
7M5DNgpeOhom0VEW8hIsWC7Iq3zqu8wEt4ziwc7PJItP6OUPEUaAESn57erZbpjb
Mi95KT1m+o62aeBSw6jFb03/BbWCGbbk4r31sSmNSbp5xlAtJXfSpRCEDRrwoGYD
5mYPqrA7/wE3RYuK4YfBnni/wR+Qe38QdHwa07qzvMTnrwhDcKfm2QGktH7e053e
TYu8LnCzq55GMQNhq/xvlHee5K+vzchD+lnA/mSJeA8Jc3BSoS+eMZm6Q03wmMNn
3Bn6iLE9GEDFS+p6anCr8pO4uCpb5IQG/EkO9rctM5h6WdgAlSivMECHNHbGkF/M
F3vlJbF6RMmzCSlX+usdC4oH3dWTq1EVkG/e/QQC4RurNibicV+mfbTApFugDfnX
0E5nwwNTpZwsN7YV5wYHGmJZh+KOp6eOFoh3x/o8hDaMTKWwDQlvI+WfzqyHZVAm
1HtTJb1dnX192jYaC8yxX3LzpnJDMUrd7q0QK5aiMzubjV/AaGEAyPtCaXpBvTy7
KqrRzvTpXgQ5h00DoHQNqwLhfQp5v6hS3CfIyPpVWjcMvRLkNMMrrLYy+lkNueAs
z7dYTqmcBsMFI82kskoiVkqpMKj+USR+1vPyzinzgJVd0qAfaHiRCKXvWuwicIAq
NKxBXyrOHM5V+DG4sXELoDIsvB9MqXTCp5Jffm2Ub+Qd5tOM5kAQyEhr/rIYvMel
eeXlD8fsHFaapR0VtF2k+fILDYXPeE8x7mj2XXB+JO2SREkHwRHIfZ2hQD3m0h6P
DyD2bDcLj5bRokjhgwl1g6Khza50wLX4DWd+ftANVcrPHOm+FkBewVrEy+dpmhzq
qLnp83x7alzm0QgMbh4+GhIOzH+PfnfjJeaQomUjEnitaat+6Pzl2Aa7AgV6T4Is
85evY1dasVXdxQmcvy+3s+tjF65dxg3la+WSbw4B2J7fg1E+jMXMxIsvh3C0b7W1
sv/MwZxFjMIbQDxIyLvOVInfdM9+znE56RE5whjNPAlpbr3VPpkXckYpmcjdJtjX
aMvkXzTfjtVXe5nIRpvDFAamHdhhdKmz4exz40+U/SzYpoa0KFa9LQtotRiLW4Fj
+gMYKPAl2R3oKcH6NQSZdmgrKw2jdsTbYzwgk2qBKqWo6xfiZDJ2bAmXb+o+G+sD
c2sUHJQLH2SV5sj1IXUhrVjUBZq0zjz9L7l3odDXOMxRAfM/LBWNRub1B6r/y/ga
T38lvjtMcTPcmLmis/2nYgHhGVNPcsG3K4Q+gBvWqkAXSn95uxjJC4lPns2TsdWF
VavSlOM/e8rp2VuT0OjA61Qwl8lCnSBwVq7Nasd7LIPCYFQjH/sYHN9YpJFZ6iU3
4qYDo8j68iyHpLn7Yyz8UyEBDrY/NzrQkW1g92u0CbzYJAvuloRAnI4MBMQNLOte
qw7VuljmKoVixxxWv9U8DkirlBo9my8ZPCk9DOtnM3l53rGcJDEz/moqhQa5ikKT
SbyRw3O3VxxpcGQ8aXtYPYgHuRUZnCt1en3FGQpcwh+xKZW3aNtSZXkvLcHJEiaG
yBhsvrq30CTpr359YPp2/mGI/yWzDt6TJs0OhjYLgn/zIAWtgxKsaaqQlmEqcwrt
hLaSIfH0Xf+UVcTLlW6Un+i8XUmpEdebwBN0Jd2WBUcFCaCn69zUBgf0uNMWRWtL
Nz2lTEFe1OIuc02XzVikJ3FpvZG1CLsoeEM10yI4M7DPN161ZP0wfttM/cvHM1D4
9W8NBsPcVyaLcHbBw3+Z9CGRFwG4EhG+IPsKtX2oIYlkweI2XeG4ZDC/BO/lcN8H
a8AUYBeZDZ9nTt7dMR2FFKkovA8aheqQ2cDwlvj88o25IrFRrt/+9aNsjtmyhpHM
SYSjSsAWEo8lDKkh7EWdBGdyveBThYSX0TenSmGRlh+bwzdfgLlbSBODsVXPnEBD
WEuY2fDR9H2bxl4lO0FaqnMcUf7UVoVLhGGcRrLyCDfTwmaxWFHmD6jGyrl8f7Wu
BrDn9LiDHG7ibOd02X01V4CwthfqoL7Yzqxax4hppV38lk8tv9y74oMcxYjT/THP
B1IQ2x3bJLsbyvVp9JEGaZNuHA+91+ZTCHbcC/GQXMp5k06APUwedBxS+ZoUbhNi
mYe+A681UN2d+3MO0eWxIlYlyQjrSqOl04El0MJ5GpChR+4QymCC6B5Rik1VBqRw
pcTECS4NpykBn0iuFmoCoF3AnokGgitBCge8rJAELK3ponm9bnkiHCYF90iVmMhZ
kamOhQfUUjz/UB+e0gHpMNL4TUWGz60drl7NgyA2jjava9o0jHOysQrdlUwBGdic
SEiJhWZudPrq9d9kkNQw+l6etiVcX1HUAMHwwbY3H9Jt16ed4HCE6zJ6jW6OAoSi
CSvPVoJoClHmJMgNU2qCJ7U23QrMgPLz/gOfEYGl/knAuUFcp2wypFN4HXiGLIlU
1FOPgxIQv+436Y4XW417/WMsSqMoMlg6vImLbtpzBOsI13vUOFJSWgZXymbf2Xb/
pZ45uCb63Gij3ut6YkgaS5hLPTKnZLz05+HWtTBw8Z1aMQI7i5hjBQnARo4D6KWl
GASoei6NHjzg6/QubuV63ktmGuKxROO3Udco3IuwheZcseDTleqjnl18lKMmQHWO
Zae+XldYUGIE5sfLQ/sLFBQn68AMF/vDldfqZ+yCJuHUOr0i4hQG/WNlBfjqi8ZG
i/DDoQ79zqI/rwWm44e5zpaamC2cKOTDSYTruTzaIgroFAEXuEZCdPpJCo6jtHPa
tGR+GeZBlzlJgV+jT5FjtzJSgGeuJSaIZctN4I+yKWZYPhwqkgE6q2A5G4ifSwe1
gBCvNjJaej2+rVFvYWzvMDksJhMK4X7Q9RYL9D5RHaFeSJ+6ftSAqe7xf1VEyp/v
RVliBmJ60LPUe7exUnAA+SihgxYHsU2rFM9zPuqRPmN2CoIgby/lRgDd19/qKAFc
jOE6uFFSAXotKsCHihrdtzqjrzfYlt38OcSz9btoevH4PSkERkX06e3E6SQzE+zZ
Y0p7ZIyuSFsRD9jIbXSZyEShf7owR/ZYCTAT56Y3TLmlPp2Ua9XSXC3mEd35ZlrC
wjuHExxAw/oelvcdyj+q1+fOrJos/wMqwjoEyzNugo6bLmaHMy0FqsMRICjiRa2U
ea6TXJIwMMTAT636eDVR/8hwdAN6G6F3KcmxZjhY5MeA8KKodH6fFsfgt3p4DrYB
TH2kyYYjajGg0B/otI5sP6qgWsPkXpqL3SaKpN98N7WjTc8SEOZW3SJu2fmE5c29
I37X2wbkJ1GC+x7qIwXucIcGmL2dvnbAD3qupfN6bt4yh9oSWjNnKUw+LSGegbYL
4d7EQFUaIp1X6cQdlA6MiLi/YJ0hDSzvttcNuV4DzvPYhEttKE14v7qN83SBqi5p
f8uS7LJdMFcYDBw1kP42rlydzJCb+yCUgN0SijW5ZWZGn5zl2ciZ9Fd8KdnPtg68
zqMQ8GCi8ds+sHsR4Eo2LqdWe5y+61g34nk1LaxOmLqwBqPnWA/2drVghLLlG8TU
iHXhL7+evWeElfm8CrKIbx6wdrf4qZbn+2KxLo2Opg6y216QNzrtcdNIQgQ05Nyy
A77+gMqmEDmTXyWqCozixa0cYk5qBwmC4XwwiKUNIYeigVzew1ivUms66y2t2i4/
GxsaYdW6OBMKawpvOv7rVb5XwVpCtkruz2ZvO1U4527LpkyIdE2uT8cetUNoJevC
sxG4MwKRlv5GGQIz/bu22dbGAgMC+sJ7omz0QCg7N5x6KlYwNYT+kDrq5tBPOO/+
290HFviiPs5CF8GLbMQV/9hhjZenXA1GWTtTh+ejgFSml/HrD533ljt8VJIs42Kl
HzLM8au88+yGN8VLIMVsCUvWi+P+jb9LMqBK2bY+XTBcC9oEMf2gurvFZK2hUvqz
TlSTINqb9FOxkzDOSdedbuqkBR5IZonPyIkbYlUsk5F0KWuI9EwpxdTalRyrWoRH
HF1lpACwy5jXPPiIirbnPC/d9prU2p1g7BtuEDgZr1MI+8gZpb/1NbjLd3uJtiLg
7mg0UF8gEdzJhzIXgbxLI3HnYAk293KBJBdhKhAqfs50EMh70GXy9y48T5s4AkaV
foOBs/5eKwZOzmAHYi5JvpKAJgBUscbqvm3+SaNG9VuXQKms1FsRzJjFqrmn04wc
hgfNVjycU89imyYvBsdFGe/emdS4ONBwDfEo5+cze65sdtgD52M5CYxnjmFh00MV
NoqZPg9KJ8fVZX48M98nXJCDpNTosXD0nfy+x5lR6uDL7J8lggmjGSsbI4dhlvBX
JzfVDSArJf+BsbqaWUPCaTigQjfPJMnrPHYwR7OMVLLT3pfLTEWttRTs12ny3VUT
bg/YicFO6c6Y6RCWc4CUaMm1v2LSaCZLsSmdngOCGxzicH+Bv61KtDwi3Iqv9a/f
AOU+8JcWOQUXsY/fYo5vakd6xUyNXo5z6HisWmdyht82Bzm3A3mt9mTlIEyvwCjH
YYkOrJ4Yn3L45FmDhPislK4tv+0OAPpyUmAINcT+Vh3iViK2ktzeivOEQCr5X//L
sac6xSoIgCrXmKpxnZJWcBKBXW/7OLlp9Ik/45FhLVeGxYYWYb2u24HcA2vF8L4O
mtqRYAZYi8SBv3Le/4fyVKpNJN6tLHe7wQ9VCWkRlRZdGb7QqLlmNy/xT0cQm6WC
m25RM2oTewi/EXyiTeog0iCwFFIBq/8ToK/ZPaj+qI7T9HLWxtv746BK26OLwSQP
6zhf4LXXJxM9QwB3mgOPHTBb6p3GbGiFTIKJMNk6fhADN/ynzklZhT/8LfrL4y6X
OVLz6KCCITXFUQwElDmsz48fqfzhMHMaVpucjYSS3XIkvBDyVMbRainyp20uTKEt
nhY0aHu0q/5CnGMcFoaY7U6fhEteUujDuitR0Kk8YG+EiYx3RrL8BJMkQaWn2Et3
YfoXl6Qie/oRkkNjliUjW2O3RQcOHxtWQFqDYg/ICz7A9nP7OLWo8OZv1Dz8fao3
w1u8A4smth0be+6bO8OhP3Yni/flkS1G96l69S6cRdoW8zlhgcn9krdVPKUzk9ra
NDMbYS9YxVlDlA0mnfCeMUj5ptpF0eZKKQOQGDwZkvkJuALehFsH6UBTn+/uTBPC
mXmgqAn/0Ze12EuwUsb2AqgUBImk7YRC/iIEihPiuVysL2QMxsayAa517ppnLfLj
+stDjfnfqzqa1kXpG8cNWA1il9EFbRBNw991BwNTSzL1yGpRLPJtf5t6x8EwWBoe
dD3TxBUKdPaeS6D4qaZwBf4EbIoZXN93PQs6n5OdyJFG78NLuE++MzKqinHkj7eG
ld1zQqPUgRbW4QJxrAaIhmlJY+7+dRwLYGZLZJXM3tDVWj07MMf52C2llEX5VoO+
yMQV26enMWtUgblPKVWlpnFweyevrDxWLysnG2yqXXqn7qASxeVrZPou6vPvoOuS
GS6n1Wp6oLvpdWvqF7X9YXHvYc4ow0nFLdygB83e1Gz3q0BDqe0hRf+2hN2C7hMj
lkKJGe1EquZZsfgFz3ImgvWfYIJsPr4MaeqP1X4g8I91nzMApOYqfmqytSrKXrgY
c9Zb+6BQIlz0wO4xy7/pPnUXKZctzxYJ188aPqjoc0XwwU+N3vESX2M1Pj/o8POe
E0R1cgQr7ukfGpOQD2S8Q7uH7k7UKQirZ7l5eRqMKezzBRL+RU6XhfxWd68XOZak
sb2wLTsj43xO/FkXjxI5sxVkoB3JPYzMN80t7kXK8roGCF2PBnhYA4PUM81Lba4S
d23JvQvi/UJAg/cG2sa6/p1to7I36MIFv2rJJAphnHcUzgbMcFuPrjO8ZYSsIIGS
MM54lb2ZaWwqQ4nXaeeL9jZjjZLSEetr9NU6oufpgm6ed3gss5t6OHXZwQGww9Xb
fOf0rUt+GLpcoXgzzqfvxiJY1PFHH+6ZwLyCB0tEgPNd8JxJ52qT7aBiRRMB0NU5
AeeuluLTMRyiURplBvDP2ZNxNMlRwNmSYntnuR0WREbNHiLc9Zz7twsNyCIIW2BN
xtkF2/Khj4oqRyU3DL2qympp386gR5zaLoVpMoLpE8KZQvpa5wMncnqnPbXlu3eo
EZQhUxI85Uhb/EBWd2oq+XDmWeOeBPoDzUS2ziDFxf4uWTqIOf79B0BV2irSeVWo
mU4Da3A2XHWKKe0+DsPeX7VxqpxrX/akbSMskOKh0stZNC4YFYGUGXAIwlPlbHri
xZKzws//OpCXoooPNw5gPzguNgCPvRbY8gqWy2BALs5pTzhtFlhCnfSo1Q4U8mDi
5qYOFNHeVN+vy1TspIIbpVI6+uvVP5qlP6/EBk2ajRVRkAwafaZJ2VGKs/5Ti0YN
P2X2FnLtZ6Vx3iLzdrAgM+nfXaxMpWLulIu1sZxpJLWAlQpCsQkt5h1BkBuShKuO
guIvEdzo+xBTjxcLdHzhbjL7ykpyej5x8pUhjRZJWRaQ/SHSKValV/CxkR64KFcO
ie+BaNZyQpLNmIg6TXD2J3poa0qWZ/o2eUawwmKN2bco20b3g13VfhkPanyi0BZl
v7subB5vLg868TwMg4IPdLOF7K68ThTSMLtc94GK4I+ICFsIADoAXApowtIYcPcr
G0mrMiRqw1/EW3L8g77udLIjatdwWr+Q1M+U2yIwOX7UU2eZ4ZmGc6h3ZkdtbG1Y
sC59S16GeZqqAx1Zitc9nIfNA7Ze0oNvhJApUX1jpt9JlcZKsVaVcFIwOdNmid4P
ZQUUa5AQjcmeUPUyruz0BqEzdTgx0gCY6Fe8o+WBOjWtIkkaZ3J7QPvY2jQ3m1IP
7ThviHnE7GyLfCpUza7rSBRgOecSt9ErGL8QO+TvK4dcGvzJgdRVNR61ypCoQX1I
ZvONr3dXiVR/W8tBjf33T88hzYWUfE6fSo8q6kvytwQVlqceuxMHvcOEnAt159FI
xZZRetV4D0XyONBJ4ky2iAWvGvHt6vsZXYyIAqfWRE9Gt+6U0/YkZ/cUyc9IHGQD
mAeoclojEXnqY7Y6Y6hRcaSWeucG3oxK8Ew+4zQsbfY02URzCzIEfBhkTzbohtDb
lwPpJDeXJOAoy7kyghekxEyQ0VofDWxxztrrIt0zNl3m3kbkHcQDAwnOZmpWKj9/
18OooX/TBl1po8fpQKwq92GA3vSdtdwL8SGdgFm0BnUOKJOmiY1Gy/A5haMCUsdB
KWYAaXEUmve91yILAnosXGIq7IkO9PR6D/djfyyEs1eljRNYT0NnAoEvapEWSXW8
+v4t4QIFkprQ1CE46Ilm4qCADR7PbsG7FYpB4C63y2lEfiFZKc2gUcsAmt6VIyl8
jmMiD20E95RP4Q/LTHS28d0czO0nj+SA5mWrgO8inNJXETiCsfEpuHZt84CulUtt
NSwiRsbpQ6b5BCAu7V3vht/9IGf9ycGbX0Re1AhDRNMc8W1eoijgmLWN5f51cqSL
cWeOY7UZxWBWOljYuVIVg4m3Mhp7tnDRlIW2KW7UazlF1oo2bW147N7vPoJrvyM8
7A+KsX8DDCBPiVxdYBF8SqCBSWmetF3zviMTo6WFGrmNCpmR6inIosj4OuDQGXkB
VUUkFT4V5RA0gUSei2mRA92EW2PN4gQt0TONiC9LbMbgarE08ibrlyxtAKLGNy+C
LWKAV5sObVmV/ERIjXZ6Z1ZX3THKK2NAnC29wmchcNZ2H4u4pFC4mFvgQVqwrlvN
rAzI6meI9LK6GBmfbGM9ETJvx1af/kr+Tgdw2X2bUpJn1ugcnpe3pU2g65N+8R3f
T2pGhsq19Uy39UgmjD9+oWSM97w2RWrP77J9cn68RmbInEEDODGKA+iYyjtXzZN8
CPI5LCGmJRDjyUnkEjzP8m8c1had22cdH7WpmyN3HgpnamXwgs61GvGEprQTnIE+
Y9CwhEtBJrBr9zR9fLLFUm6x3nDOmwvD4uUdGBW5sXMoGWHKPKQ9Kv5lSoR7UtDf
w5ProqQwwhXyWpqcC86w5skY5r6SPixx53/5fOc28/46Vyzori+lOvTgJdXt7UlS
ZdXeHKKbDXE8Wtwj0uMIulNCtU8tQADwbxuoMr7pyj7aad88bn+I02RKPT5PJnzT
sdXkdgCHhRSm+x9Am6N27cDVzokKxwB/Bq+nMU9rIVMHbEpsIxgeeCdt4uo5jcyk
hHNI1ICFRJoQHaoNX8sO8YJmSRCa5cZNlxyEhNEJJI02482VnzMbqkzq9zaz3NCp
gZxmmEWZ9Er+afLVvUVsFxGoL4YyEmwjgazOin+ZiRGREtL0iXYxnLIqh7dNQqxe
nHm5uk9NPIDWM/SOpCZLdKUSXqt4tCzPijlfGB15hFqOPAQWEjCYZ0Dz9UM4edEa
QW8se2pjHBVFbVrKVy694cisati+tlnIU/+hei4n78f+FgaOhc+OJLxg7bNF4M0S
zqdeq/2hUKBg3Vy5LJBofJDgJyoyWQkVToTGNVdPpvWaBUGrjXvszrKKjFD3k9Hq
p7SYM7IN8TUCcj71OvMNaYCPjM3msBgdSNEZKi3N/wJi+zZSqtQBpbklaRw/JrZV
JvskYWcdTq1IPFSmKvOhzo+XKXY4AZR1kbkyQVKFokh2ERp3Dj+hC0d8SKJXWMJt
JV03UE9RwQTvcxIcnds3j+ESoimnP/rHCzdx5syp4qSbV+Klvegcmhn5vLucSCxP
qTOXqHRjWHLW7THV2N1if2sZVMjEl28QxtCd/qQOszMUhIzUGfONqz7rm4ZqLUmV
M2CjwzdtIsKPvRw19KmVlrjQjg2to75hwYGmbeqeUF1iPQDegiVsRKamlqOOGUIM
39tBqRr6wtydfCqgI5NTiiZSLtZmKkx4ArArQtRa+v1YnMw16aJnb+OBBMRROrmC
VZni/iv8uEnODEzvjBHzlTgIUnB82TN8GQ9XWMXKjHMcXoXxyJtBGCPdfY3rqflt
6g6OxvQDNN22EGVwBWpLd92ifXVQFZ/Po/fj1+Ua6AwacWPfFCzaXfnZtD/kCRMB
sOqQ7eit4+6CaL2S10YLE/V9+22kOQMzIAvZdZ7Rj1M7aqQwgmZ+YT3V2czKk42z
Iu5qB68d4SKRN++MVsjvdhvtacNJb9X+necjrAcgn+aTbk3jjB5yz5Lbt6LCFN78
Hmh8eJXtXnF1oUuozbs36Wh18fmqPYzOHLFy4pSh1egY/JirVWBVHGisiy+QUbNz
4HNBWIYK3GbAQ8QErspuymcjoQsC56LbPtIN2DP5byENHN0iwbhk7s19RYCDHh2I
nBNIHeZJnN2JmFY0TVRQlvNqCQaw/LRbdY81I7tzpw1t0f6tIytXnR8RfsH7Muli
CmCLvz/WHc/HCpa/TBr8LAShzDBLhfgvlp3CNYGKWlDn1mE2fXlMP4AgKnQEV58w
BamWH4ii4uCHskotlnYowSf/Lim1hvG3ukBxzg6hVu/RxZhd1oDdYvV6LLC88Wsf
zIRzzpDRZBkerOhY5XOAzxMPlC/3BJFDNttV2222VINBv1U9FlrUzDRALS7MGMnf
tRYb0KtjbZgTPySwpNOOMtSJcSvVGNYn1R9WHlOidBM8PGZQrJL5vZhFsATcNeg2
MEzmopsz3HdNwrPHVUMkmxCT5pqSLFmW8R+gAHpt7zNVM6dZV9fQ9s+swPVmDtad
9zhEE7e05/iPYGnFKv+LAC8StVLZkELk2U6NQsiBCR7da1F6QVPjz3eeSR/2FSJl
ey6cnXWop9RwUIuUzoyirZDfekDG3bQ0CrQtQXCstPMN4JNS3dyocUt6+Rc5lyz6
c/3fmbfOSYcUjoIOkzCXFYmtNxwP/WnOODqJeIbwe01q9/XMnfVv6i8JUHTWa1m/
yDPK5RVt61v7i40T/wGFwEK1vscvzjzhRWYiKS8Iu2NOe8q9hkka2/4L0/w36y6h
CzQF41w+FuwxeebDFbdHT6fZdqskG9WrKYmT8W1j98/g557NAanfUybu1YCMEJKt
WpZLf2+9TfocBGo0fSh7r+wOI4OIgOvx2jZyhXWfLA6stfa6hVkSze1ch+COneDX
rJj6ONdHI4vY3K//tW5hk6kVlUSeKoXSS9Om41xcdZ+thNfJIY6s9H247FWulOsW
FX7mQ+nlNqcGZeU7ePAmcx/RvqceTG17Vh+guo5VDB/9l6hHP7U7751cxKC7rfB/
0mp/b/lyeO1sK3RWZVm7ma3XzCAU6BAX1bEYrd1LgLlwGKnn5U+5pChWY2eMZ7hg
OcV1Lgz2DBTQFoc9l7pShMhC0j1jFuMk6GUQ7xXNEfpw1+Rx2Bf3VNBWt+5dzUfV
yHpp3ut5zecGV2ALMITGugN5e2Wn7ijW0v/ysnouupWgX7RTfg3iNUmV1j03fRjB
tAJ8P+3ovTGeWb6WpoSw+/4E/M4KE+x93V0g0jJggpKMjcdPEVApv9z7RQ2128nx
cLXxAzTWb9tLt8lWFASVq+kpCqD9gkXn74T4+8TrEkWysPPg38qG73mHHQpfOC6l
7CHM0rAn8nnKx7ZlntyWU4cP3R3sX5ebgtPqUCMkQf+WNnG3XHjna4raGoadGDW9
FN0WyV2MPgDkquwppV8J3BkmkDZjhnTvEtGxnLPBi+9RHsuYY49avN1uTZYLmxTe
5Jz13Z0M2TXo2muARRqSc0dEqrtuEF7pbZGibBRgU503BwUhL4wZ4zo8B1oGmqhc
yOzNC6/9vLkfnpzMEapB5D2+X2ly7la7GINMthGpOM7br46O5lpw2eQ5m7v266Mx
/31wa+cSO+rQmAeKM85/EX4M+rGhz8gkL6QMMn7tGGJgzEf+ZgsxH+I38eBpWngd
WrIR/yq76F7Yn3CmPa04KQCkjaB8g4nKqJ5AC/OmFzxmhkv4gKrgc2ug/i0ymjJr
sZiJU/0fVf0KU7cRwfApfdX+eIC2hWsJdsiBc/r67f94NSJTH5H3Oi0kAMXchykL
lzFqkOit0UKTpJjdweMDytOcbCYppv+NH4wAnRoI9174yRCJKkFZS1xWBv5y7v6f
1VkD1zErngIXEr49dxOSyv2g4Ltim0GnLZ5mQ+z2GfFFsYiP4uB2H9cNr3VIU+Qw
VvlixezbiDuMwPo692eh485WhSsgFI5Y3HtKz26lQgjyx7esiLrDie9gJAui4W8g
JFfHVx8MLfKcbKnsiPplZrdJYDXIBEmlCtB5wmf/SHH9gn9r+xzeNIrKrNldaphW
xTt46xHwz29IRVNF8WOOh4sLIM5uj1TpjO4WO1osOOzVef+0d4dAa7bFKtIz+nkp
dbiGWPEe3fKKE1QSVE2sr/m5YSHAMBSaoa3rGSbKl92gUwMM503BOGH7YNTQhAaF
p0MuT+NAIjpCvOmubarmJAwW/nrqgpLWoukpFe+RO99YQtVxbj6LbNsevscjWH7L
trQ0sSuCH9w06oUwl0Mh8iZSr4aSxb9NPiNiXFCnHpZkUkDnpzuFB+A3ZRmXLjGX
s1RlmsS2Aunr+uCG3o9dvTMtCi7ndZYSjqLckB75IAYTdKtK38i9R+GcKahjnmVP
dA3M2Tw/t2QGedJpyA1VLdcRbsHaU20OSyEBH3Fm9hrHc3SLMGAOvJxGAMtKIE/L
NXoxtAA6Gxi0pyOowX/ymlVwNa4cVi1pRa6NSkw+XkTnIcdRW9hA54HpdqT5Vg2t
9ZHtrJXWy0cjywB4439ycpJJbbRz4Mu+V0tl+oscH6ZM6wEmkYp1AXcsQW0ysma4
5k5LeLHFvS3XcrG4ZNGUw9TyvzjTIITbIBdx0YTOcV1pdW+rp4mtHEgCUYG1HTvi
9M176ajzI7gPSlttHgABoVKhduKlqr85+LQ4LSaKBBlEh7PXB7J1CQJMvYVnCBJo
Bfa3zidmAa3On6AypoRtJLFLIXlJiYM0D7ay7ir92u7lAzMwMraOV2Kd3FG4XHUe
GrE5jn0AZlcrS12Tabh5pyQp51i+sKh0ypvXWMgvAU9R/kjCC/JQxPZZhrNwLQLT
WIDAT7Ixn8ewRwzmOqreQYisl94ZFh5SUi1btFV+h2JXQR5hXN8JiYbu99TRKNSU
odV6dMzuDrrq7m6xE+lYaSATPpUE7Adg+lfbxOQBUqmwLA6Ne+fsCfFye+vJVvyH
eN3QjyqqGVIxKHuogGhtR8BcpttjS5Jo2B5UqeMaOewKI4DRWxvBx+4GXHv6JR1z
ZZ/mESL9a2jBVG49DXaU3SZ/WWvwsZT9Fq5xIfXNfH+7aukxMKqjEUoHDYFgMqB/
gVvC5DcI6pgMLuZhSko+5+le42xrrMChRhsyRLlF7so1yPMqpLF3T3T+WJXjENsQ
t6Rzyn73lXh8YjM0XcqcKBsIEmTefq4DY00bJkP8eoD8lNRdJ3f8/ydgn3to8wNA
9EwaP3Wy7rI40HWplv9hXMV7Nfbvk9y6urjTduU12289TAUTS0eiOiECywP3Eqfg
uAGfY7Im8ZiXPsLXWcq1+ZQyhHsUsJPizumBnjH1rzWPX2QUKjpNiNLqoWKrJNrd
osavA/Q0P9Cy7VwyNqXjHIwXE6wqOB/jSu5J30Wyoh89Dv0U/wHwqi2BWWmE+5Ys
75gpwUoLSCkpdne9nskQoKhJes0EFhUwlKLPhyvlPQGmlVAxTE/P9zDPp2pEHXvD
/sY6pvNNLC2bt1fs8A45mOcmn4vS22TsbZiPeS4aVAFwrYYAmkztiihghASe7KfC
YeSRePYroWIb3ym8PVEk2CMlYUgDtotl3/eX89ul5q64SjVeAUbsoB8NmqLfRAf9
ry1mObgT/HYiNl0UX4JCcYb6SUwSfG23LSxkyza/xPZOoZbLmsOn+1utiUzqeG9F
pqlM5sm60cOZ0ZfD27nsP5thW/RMQlpHmbBZu5sEdOg9cE3t63FT/oA0sxBpeKp3
o8Px9ckXx0+Bdm4JhkgAJexaj4TqgMILvxezNNzVPTMUd7zdozoXxofQ0xz90omk
mmfY5ZHSYo7yvR4WWq26Q7I8ay6xZ+WLB5QBau8NXTWMygNCM9CeMK8E/WoS3FYm
QnWP5m84G/SRXIJz/dzuVy/HBOI+iuvX4E9LtB0DICgn0D8mJesHVGF8gnMH79d9
AlRgF97Ag1JBKS1G/7GR/pyAAfqtJxAaWqnSRb4VLS9CtOUKlszVuzDsLBNjdL1p
p2zArerkwjwlPZ6LvbuPE0PEA0sLd463rvM9TVAMtY5C7X4HRWLCocV+aGyLuNGT
p/covc4Pn+GX6bByGCp/Wh21SdBnkLzDa6SEOcCvHQj9v3X46+OhMAOya1tqT2Gp
Xr9yHyygWLI/vZWiKLqC2efgIAE0j3RZsYtOQSV3Uci6e20L87E1AmUe7M6VwaYs
CEKLpamW8W+REoQKObtaTZxBZJ1w7Bc5aoR14mn2oc7MOxZhTTWOtc090utmf6d9
/YvcKExJ+io9JqiwzZB0snm6RUi7ye5DmIn0oM3B2TIbz8H9w6qdvktigBJ/I854
41RL1FL8J0qn7j7cDq7/hV+b9xBC18b455FN9NkUR/EMkB3HKeIDqJeWh5erF7e1
SHuGty1c9KKY/QfVezCHQVztyV7q2REYxvFGxBlVpcLwvWnfhmo6TlOMdxS+tpN5
1k7cZRHcdaJkbe8Oy1vMGMfKMsY6moX5OOyxX1JVttjyzZabwDQTxFyvJEOQ++P/
lGQ8NObCNvGnaBkP4GIYoYMIhJBkKDEffEPpvnJShvBh33yewUjrB3s2q2+gpJQP
WyKUu/LKHXh9XK6tOArGjOp3zR9BOB7yd0vRe/1F8XoTGH8FW9r/7ycjXh5dFZcH
3FfJxUPyUDgwHIwf6htvy5TK+MxT0PXOZ7gqn3m9cYuJNp1ClJLYBPbSBDgVoO8M
1LRGoiPl8z0rFhDf/5pWans1IEYUCx0f1wX8RzJ/92lCsUSCBMHpt0ZNxTod1RzO
FWoImzsf84EwqEugA17Dc0F+uxtLixwVpwHU0ou9mz9pExlKaiihMwIYVe6C+qiE
C2+n7eIi/IWwI7Fj021XiwkEwEwO84WEqqdl9JYazmHsRHyimonvwbeffBpLGhKk
fA/VpBASTZkh4KFVX0fPPJOsUgUoJCBymlC+rL9AZYiz4XzrjHfTHcQJA/8Jnmt3
ZX8rMHEwJ+iuzYWaJ+ellZHCVHLydRXLAuHDk6EP+3VaESoIoPrejLatxz6MDFn/
uzaiy6Ko24BWDr8pe7e/Bw3EdIsP+VEdAEAMUgbBSS83nbXL2gpefbZC/hzSTMva
3zpUVRkTzI3J2kBP5rAip+rp3dRyPeM15q7iQbiIVJhOaG2DKqNeKX+bg1xtaRAg
nNSZ+RW/CbJlN8rEuGfYOwPBc3ARo1Va2nEURS0Kdh2EfXUvZIkz0BfvSom8MA7R
zAQZv/9dYVOUGKVEdGq3Ebom+/9gx1Gb828huUxOImctiOLc+2mBeiim6gEjJaxV
Dt/FtxY8wgfRwyXWjMbxiGUdUgoGCz99QtPRBQ72GigV6grd/tcC6ayIbGbDXssU
FWtu00zvTiy3qBGPy5z6m6rfqK5o5LgPAKwAU2l2CRoPl7fWjP2a+gJ3Av9xx8Pg
DgfVU/dPh7hOOSUQjz2injQYMFT/L9rulaN5f1TD2Kq3gkiaFA0YueSngBFTD0T3
s++5ghtaGbbNGe22EKQIw24uNQPFRQKXFkLjQMTflX2+qH1cPf859m+UzB0gcg4y
+ZsfsWPxP8LNGuFhMe2A0moPOqJmPop+6mLArMGgTU+IPeqg8iwmhFsQZK+aQuCr
t86ShT+sfIwxDL9/UoEV8lSncZVe2fPyeWZbt85fwQzI+N/X6TTOsP0AHqJluOga
EWd4dxGVN/2ixRsS+SwJ8gwGS64zMzS5tzXDP6BPD+7XEOkPQrnq1N6WVHfQLGOv
BAPq5sbADEmT6iYrdTuxIsiRlibjuAZyEEhzgnXKcuYf5IpXbIIukef0Or6HBioN
vDOSrmGcH7+AiNbm26KOAGBXOc3+kloIhRXibaayleCcgh3+/gR5/P7lZn0AcCwZ
da9HB86sqbYHT2v/z3oNdxEbcumnc4+Zfyy9buya5cdLvd93DbIHmFEZw7BPsU/p
/Jsm8D9OfR/HarATmmdtkRvNdzvbm9/3TksOOCALJjU17x+AeGreYANkxlQLv6dx
AqJbWs9Iog6fQJdwilRNS6amCKqMqGkkVMlkxUTZgW846yptOUUGYteu23TsQaEJ
dRfBuCk6GW60+1s4zRB4RELGx9WCzkgJw1m4fFu3xaEN+9eor5UAqA+I2JzmIWNI
+pS+adclzXKuzzxI8FWcbJ2TzOY3GjfI2D+NK4KptPUdeqqzXqhaA8fX1hEZD77p
FCGMO5uXv7iR19NAvpTl84ooRCstM2MXOwebwax4IJpOKzNw+Q+erDpy7ZGp13U1
x79tk4beriD+3g1cyR1mXlKJISucpRt+PvUw3985s9GBYMBKEY1ahD0Reb9Aavf8
1318siGr0FWLPA2D+s8QUGvVkUxzRrqCKG9+0pn9xKeSlXl9v7lx1md7uDFfyEae
teC3JWCXDNZRIxV7MydlfhmFQmW9RwX+K/ab0wr/cT1O/L1d9B/HGB7MRt4fK9+v
/uIZfhC5EJFf2+rPXQ1fco+WIOR5KH6b/biYXN4gkuMkRu9YlCXrjSREl+hASqdS
IeIsOIU4JIH2Fx10YZcgc12eyVdSnspBDFTUVYVleXbdyJFg1Ch2wdoWuJ7cwUi3
Vy/NTc+YeozWKys3j5tm6AyJ4vMGMx4n7L7DWIfaYQloiSNrK+/r393PhYhqkYmU
Dxp4ZhBGdtqwYW6pGUMqtjkJ6JlkBK/Xm91WqvFWWnolugrMS9wFJH3nntxHQor7
HF3O0o3TMjULA7FkIskg50dSYUBb63pveVcWdiPfrlrtDQaHHWXsjRczjtjQrPzF
rycaTMJX/3X+Oc3jGq++P+6H3o64TxAJSDYEd89Jsx5aXJnDAjxATEA4u51R2bf6
mjxLv4pJnwKGA17gHf7oPFWxbI3BuFP3cCsQ2pPnaZl1RVCLHvWIUa5TRhEVvan1
0sJoHrpYSflN8tZCRbB29ws5bglVBTWKHbC9kjT2+Iys5SUzoEtqXJhxBQOxRh7t
9QcGiANeSbK7afIvJO4kv1C+kMjDR6FTx3t36KXr6cxMTAi7KporXa6bGARj38q3
0ZCX/R2fo8050KOeQnPGPJzF1qBgldShWk7GwJxv+koeb3KWUFfH6pzZrCmzERDF
XC56u0AOodkYLetLvedhVW4xZbiRm3gxI5IkHtuyuEaF7kHUJrEdL6zs51LyMm2n
ZVdub/0QeFGk5XG29hFKekeTtBgFLi87jTGXrN15i1eWHfBYD00ZOK7tMBI5/MBD
myGCmUPvfCzH/WpDUemqk2VtmUaMl3+mZIrAM94dszd7xu3LE8v9L3co3er+tB5C
3OnV9J7h/o8fEaZu/5isoFFye5zt1yjgU73d1yRLAnT0GaEaVcdoDS58r24ZBUdu
BKRLCDv4naKF/hq/wN9SWBgUYj8NZQRWOoJdg+S66+HFv7DMXy/m9jHyrSdjCVNW
8T+RQz8giDwj4PzIcZNxJIpZGHxJH93M1ovn7QLc31Pfulpx+W6KQaj79IMUKmWp
tIoqhQ2yb4r8yxyoVtDFarzjnd/AGOXN85sipCWQK+TWxFTQg5dts5q6TlXuXiv+
q5Ku2hJvuJp7QDyiOm2aRpaaTJJyy/Vln4B7Lyyyt6bGHzrnpDgPYEp7Sg2EA4xA
P24I8j3UbsmZvBaQdNmKcDUJ4yW5X7D9VVWmbjPdvytlzytSIOaHxnwkUfgQ6hzv
YcLH9sZvxR9Y83QFOqZlvbfmcj3ZsQ+6MqzaCzfIblgeyOj+ntVJw2c/nDpuAiPT
0+8teNfPezwjmjWaRGXhRYeXN4BWwA2VolxuYfhdSxooQJOpouyrpAYyAsCTOQb/
h8/LJ66XgEsprWbhucoGfdoMijCOFKPyJT9/EBcpaB1mKaaAMpzussoSDqpkIUSx
Yyl6kWIxVQ7sMO/aO/mgw/pnzhxaCqDmtQkenB2P7oTMGqnbpO3EOJcP2PbsJaEq
xt/XmxmWPffhxcYgez1RViHbxNnNb4xUmNUIvbjMbLNIgV9FJZzX8U1h8v4Sjrte
/fFhOt/IM19wi6/CtNPUnjD2V8me+8dC3Oy6w+in7Sj9In1+ctVZgM7c7xP6cbEd
n6JkEj5h5LyrclWjPsTLeJ7AXDIuU4wcCxKUOWgHRIEMpJgGaQwnTLAiK4OmG9cs
M7ChGHgY46e1EVm3EWgoXbI7kLdULtQzaB+RBHXumGwtyI7zJX6ETPVvl3WMd5sn
6zzEY1+FtZzMOgEHcPYZnUoGD3qNxxJRMuvHwRUNUcItb+JUMW4ebDer4Ohhy0TX
Td/pvnWzQVlwg9tE5sIiFcOl0/hk3AXYiWa+MoDw+8mcZbQ2LqBml4mctfk6Vd5c
wBMHAd7dLRVrLIBFWEpz/VG6sancJHuHE4K3qamC67ZRcv8oZtwX/O/vC+7EtZUx
Zr91VrUQkD3I/N1Ul8NVclAPZTEaueqMH7F04enN+YxM5AGdFvuBYBwGAAH4gSPM
kVfeB6OMp3Rk7s9Xyj2a6KKOJEOt22Mu4FtRLIcJk8THWze45L1HKcaUOR0GldAi
iCh3Yzy3sCrh/tUDe7DyFLFAE3tbjUuJVUzuejGJ/POptVNP413DX0lnp8QImkpO
r7p1zmuLDSLB1bklosQFMDefaHY465XrT5Kvrb2orrpChoGaax4ZyGJ1iCJHk6/j
zF0hbRvDZDPl5NmzCZece9rc0wwLKQ8qyF11JI9x2kqJK4ojgK2904daBz8pIinK
DNHFdtiDpwV+AMQidg/Pal0Vsbn/fzegVEFpdAEPSDb6CT+xkjdXcTAx7r8ZphXb
sX+lBh250NEBxjxNW5UeR/ADU/fQfk408L8jB+d8oigyriw3tOnSFRMG9tVemWt6
qg3uJ9mwrqJHay69+AS9Iz2eLfXODYJGJVSUcPuBNvyrpna72EHqHkiON8TD+QXb
HPC58mPZ7XvB3Z+BC3Z3VPKhRXsQLyoBn5L3+iGH9ENhf/H7Kx3b4m4vgJ7pj3fP
JpQpe6VGuMXnZeYIPqodgEI9XlUQ68EfyBI6QwxWDlnCd2ZXpuW/8RIKg58Ya8oE
77k6pv9EuRv6rgKWaGT56VHDqrEsC3+CEuBXc5OdUS2tDgweOJvIrwQtLBD8A4lS
I1JhrxylxHLzcib5rnWOfBWXXiBal9346lfjL32OtabDrySBytY9IY3qEhibwJKW
75YAh8HUoRFwLU0FufmgXsHgMtfWF/lCMxiuTw/LiSzjr3DBAveK2ncWOMsUwFw3
FUYxv97ctUBMUUF1u0muoQbhSHPnlXjKAGnYP1k//s9nDMQwOSxWTUDl21I+Byx6
ud7EGe8KwTqTcxImZiBSYodCIrz+jR/kHqEyxfT3E4dVS7Bi7tFC7iC2tfGiZBhH
gRkmrub30O45Tc4EsAWHqbOuf5MGY0Ln4f9S2OfeaKIFRnRWBAvgTkd40136uiHO
0Wr8UaMNBebWrGvUhuFGJJ3OCnKX5ZZVqNo+hp6osXefzMlCCcToEJpCWRN8ilwp
XB4HViAll4W+omsQpTwPXJ9s3O9rbPCSgwJED55EsCU1RzrWbmAld6DEmqeCNviv
74pd7GK6xNTi9BdTSrUFE1TevnZaSYPKXvkcVUNoTmPMZOzj3r4KfN0qjipwmoiT
rQj8qt0XCmMfyYJZBb0UDQO2B+8HIGCuJ4+fgnSyEfhyxICSUMFL5kID6QSnUwhE
lFK+7x1b51Mn8dOPDcB6V9bf/cfGwU/KE6+SHKlhPpFCf3SdVEL5PrsAe4p78tdQ
SAtNtRxgSkjtLPU2pIGPr3WTnsseZkivsDUm+GNYbFBIlwuiStlZQAEEbB16sgJ7
eXhnr2T7ZcIcm0kEgtPYVSEOK7xC67mWna+XcLKslVpPKh/TfpaWSNQ3aFE8GwCq
qjgxemz77TCBzuYbvHSqtXUCRpM1BPtc8Q0T7lc2rb062fPZO48FkhjrxMpwL27c
/6RG8LKpvuNraEuJ78FgXqmixlYNbQWGL/9zu6zCrD5+QJNXNhvidawiJG/b/9Yj
SgcC4WsJ4JR8QyRyrtXj4zbA7dfhvsi0vF885+Ve5Jmt1OZ70wghG7SaZ7ybZke2
ehgRQ3O7iJlRC7B5I46IN2JAdrmfzwWQZpj07SW5e7RrqS5J0bwrG2Wnk7f5BDeT
T5Rpsn0XuEaf/iLwhRMYogBJJhN5mkY7czY9M/bN1n1h+XEWA4XZNbOR5u1HvRRq
gXvs/VUePR8Sdg1tsGaRxP66Wqt71lgHbOE9datus4mIrT2HpYSapPfxTt4d/01m
lNXEcmHxEZNNa5tbpS0eXs5anwOnrJC7xGUpzkK8Rfj/fY73JlTv5o/Gq0xGvwbr
fNefykxsISMRb7Ou9JUMYIhVXIwtHG9VsksZMlsN0n5AZ2HxpFkUVdZoQtINtAwe
PVFdugKe41T3OFJEwE/5XEPJPy/gStQ2BF4Iz4M9QH4V2+NnwbSmsTV5bJtDdQdW
k7C/ZHGKhKP7kShaiYX4Nc/k/SHZ1lCsDwzL3H+1Upo9TqJ5rTmps/2JtZjZ95Sv
EIAG11DV3/eTrkodWvr4QT2RHRL/gBAkVpzWYE/WjcygyB6mofhg8ovDwyul1pb7
VA6wWH3/bSDDsyVAsz3fob8sZrQwTdoSneo+O+30lNlsMgx3POf5hOjDeOzmluia
ipt7y+DLYSADs26DOKUR7HzjHPgqnb+bReLN1ihD0wBHtpcm6Wziu4CvfaCEjWAh
mlJE9li8Mmk2b1Bzd31W7Dwfx/XZlaPqsYvy6xQJw4ufZjjXtIqyfCl+BIvQed62
24Hez6RPlmFVAOoJJ+NQPNAUcpC2riH7GuY1CmyC2qjPO9d+DOtKCjiupH3pgcyK
eTStRpE+xLL0w7zhqg6oxW2iQJfyHFE0opI2WBqdsBzGI6lM1vT0+tdELN4x5a7W
XcqnWNn9qkTJfJ3lMuPYXMzKl+g1XIWEy+t2ikljtVirijILvc1roAcqlV1sHXkj
vDtBXFdSrRH/+SnaNckRCF9zLVUqSFfpcfCXlozv9rDESoCRR9F1ad6PEaxbWG6i
3TMdT3Kv8G/QX+4kNO3GRG/coJmWRLBJx0UsNHFyGnE/en0pMADS/5OPIrRbi76G
De4WSjztKxQs6WH/fIsO3XCd4pKnTF5WesTa6USnT9R6eI8EmR8Xu+nRvYDZL7lg
nYWFCMA3EMpj1jJm3mXrshCA5RSC3EmKMjx4W+vG8rL1posA+n7gGObWkENvpMcm
vppnbqsgGcoC4fVblM0T0xp4p1aShP9vugyGa4rIn+3FQSiSwQBDekL3ybByRrfm
MHfPy4D/vQ4iiExz5WUlOtVQKb04YcXztRQw++/tWwx3S4a6FjSmsnxAXOKEO3Lm
/AD20o0D9wX0bKPFAHqbUVA11LwIMn/lqDqEzTKxLjpVvbOY/Se6Chs+vQf/I9cj
rYbLi/ll8qxadBQTEf5T9nQIlw2aIoZHqbk6GOnxXSm54Ue5DM2TP1CsWscKVtFd
VmL5z7xo8cLLodMLKfVXZAP4PtMk3wBb8uGDyRCKbJLS9hTT1yO63dEYPM75x50q
AR+BXb6xucV9S+zp2RGnFvUwDF1i97tbVV7zRCqQgPdzSYYXoQlpOX0zyqVyO3xk
ogeuv5ZE32qtMEoeYnRfzRIjooDiLUZ/o3exgKnE1ntcXRCWG6CyAJFYC9GxKiWF
eGXs+7gWKil1Y/RsL0a2ePWLYqBlideXwCtKJPg+fcBx3qTBKGB5c7rvTMQWC/Qj
aQtCdfD8X5GMZexqOUg4/0YiPgb+jkPpT8PjsYtxgJcBuPKBIO86NDjT1fKoGKOq
EaIn/GdVQbyMJqYLeB7vLstz66L03pzfmpA5p9P9JN8a21zECbSEHbPXJ3rl4hHI
WmbALpb/sdHO9gGZ/rOk19sKAizOjCsdJM4W+AG7fQClVM1GgqACsLKE9jfBAqEl
4AKn08pjLkG6coIG7XDsRu8yo81tyq+dSETwjWHLNzPYH7w/iEuLE/rAW9RFUjmu
xOvOYxHqh2RI3RL7NqKmJYMHHOSM1LuPNSOBTn3cUSQ49imXlMd7pkFifJ16nNiF
+Zkp/E5MHO6rbf0PYt8fy/2xxAr51z2Iqv3LiAMeNr4U4G0SBc2GmrkQgLYWSc5E
C/r5FzkJEvZGBy2a3d34PelObyhc8zbvGh0nfNL64CultOITFnEj3vf32Ri6/Aan
oLHc4pS29uWNBpnwGGP9hUT7nIlXV9pHufUpjBvZ8FXtEqQ3LpXg2f2nYHWo+4Zn
ECFBlhdwD+nRW4TWZkSnqWb2BuPXeIh9j2S5chIvt/fnqIFUHrdC7m/KCjoMQmxv
yNbrbdsr4dyq80GqUJlgh5/RNj+Hdk8wF72CW7duGxMKcDPM5XPfIAoJmL0SMKKk
OhsvQbjInSQcksisBf9p49SO/T9rYeGLj7f906RBfgGI4r85cV3HEzgz+SDuAiWr
n6oaliyrlq+Q2Irs/DqOr0l1Iv/RjFwUErWCsqnvTVyHKpcIAX2kpsizpgE0oRRp
SmkSyVOG97nzxIpu86/6FOphefGj+pBbjQdkkf2gggXb1pEJfoQLU8cP3hPk7tlI
v5cWHf6ChUKdwaWqtY9r2+VaHFFAn69J+FrBAysaaEerIYHrDXes/1KyxwnZJdye
3UHObbk/OBrUCJzryUAvraAOWtHSvS5T+mo1ScQK8q9w9X9N97zT0OpNI01CsRwG
qKj35NX70WYUZlTIrET+yXKtUwO9KGvdStchsI4yqTRHXg+aIT4uSb51Sj3AyHVk
ilMldsiTprep5XAWhvlcuAcuietGOpZSs11eDAjKMiW1pu4FQZwJPF6bovGlSkWE
fcXZ47nB26Ytf0OK5ZL+SRh0UkomyY7y7fSg+vbXo+MDY2Kt7Q0MGeWtIlM5fSS4
U/V51wlTtUChqHGXzoBbzLhXRGH64ODCCeJnggwEWU1y+MD6chVPeyvp6yejaoAC
GhwC9mwvH8jmGQb1bN8ZgYpPQd6HBoIY73iGeA35L3KgnHoT4rZ73x5DrEFk87jc
RMRqgBAyXNF0kqkqdoK/eGPuehyH2OFdyJ5S2y8UuV3U0CuT2RhAPhxMFrZPaN67
wSnss7oIZ3jtfVhNVIqgiAOIUM5ZDrnQDDiTSnlKZHe1B1bkNGvdA9zRKEkKmGYm
FwV15bUD0MM3JGK96lwp4fknbcnDkNDFsptjEcwIoruBXfdOscPvYWWWFyQ15IsE
bQJ3JvCWtMTkdNpZnmUwM5DHDDf+wK6U4JONgmLf3LFCO7DqmhmPwDLEpWQs6nRY
ViE2nAi4cpYLYy/z8o1qB88laKzbaw4h1iJvlK2yHm028zM9NImJzwd5x+kJdYlU
KYXi2i/VF5AKHPIWSqOvYk4uRlN61jRYtlsI0cyfP1pXrShuWOgl5qH7N3eB0UC5
tSJtGTaG5+llvNrw/8YpkT1mkogi8FYmuLTxyqE8opv6FP6jAUGPNxAqdBYs2Jgk
TS8caSUnnU4UKIPcAdezQTbnamuvJa8y5YWlgSWGCpMfALY8ELYG17iLOzoEJzGf
Z1iL/m9WR1M3BgTUd9kdW//mI2PgPoBAb5rNEQ5EB+PS/kiXtxxJdmvNo2NFCx0q
gZqqrBqWHoAanhjalDq+KhxOA/WXWa13ppKc1TXE0UNfvVhQStUfXJhXvPF+FPY0
hQzuSnnhNPn3Bwn4XoOqod+e4g677FRA+AfVtgQdet0Xm0Ip8PKw+zUXdQrdexrb
bqmrzz1FP5FZRL0xY+sb5YEJN6SLC0y7WYwhS/uRMP4pNt4anjDiDhEToFpKOmhf
+90/3nOFA+r/tLYJbJb90EURtY3FyHzjUmt64DVXfYmqm9QHOH7DBiFpgOiq6tvk
rU+VPt0XZxKzTTbM8liEvYD6+1NPA19TFf4rmH5sfLdrrgxH5ns+OYghnghi0q+t
KlS8KXClL4QOSy3ZqLcKFppAIO/yZfFWAYZWTGFTc6u0vTOPyqRJsG/z1iIGf9Hw
pWFZUqq6sF/FOtFfLA3LGTk5lee/9TFB7d9ilGy1FgIncC61lZtI5UZUtKzGT4FR
tGHL6HWrB1dNY0RfM3/nJ1u9DtrIizG9oS+nXKEeFFiNHG7Pfc4q2d8WaiYh1wFR
j5IjMOyaME0/B1YQT8myxrsV9KmaqrN/Mz2YrJcyt9jhgnGrv3/ECAaCwQWpB92z
tFWLdBhoEnTtaug16Jpi6cB09u6dQZ8A6jlBu8go/6zf/uN7MFwLcO85yCDQs9PM
/HNZXH7jLFC8j7lEg5f83J+ytUXkPCBOJ4QmsQz6JN5kSfeb6nuKjjM7gU4m9KR4
+g4r9nufL4CcPZlkBza3HCvoJlbn9ortLZGPM1jinzpBGMVGGwi3Kipi8bG6cUQU
5ZWsZ4/lKb5UaLsGQ+6gMAwdQg625t5m2kZE2DG6+wONaVAF+pmtvwiHE7xF7Se6
wNLqb/UCarm+S7jkK3h5myEoR9hkfcQCQOmmkNtYgDDbz3qUyOqXG8M1RjFTo7H1
M+5g9VF0MYaE/TQ5QP4XVQVTln1h+uItgmmYGwkjkHeaJFDQ2hOYTZjw5AH1CYwi
jRVhweSindsYvnPrZ0hVLz5s0hHaQ13q2dxgXKKVj5jQdAja4peSMwjX84ttwvwz
m22eYS5T422+MMRQtRrVYA9MN3SR4W5D2n+n9RlT6WICN7cx09sk2HxByvsS513Z
HEni7AG6aNuZAEfMW6ANO+Tn/mKpL3/NGjMrxGnJPk3lMbkjSfnsWsxmEEpqK2pc
McY3WxWR6SVU8qh/UIzot8q89m+je7u4P85arXVSPXB4oAu3JPPavEp2UekGJbFv
VSGHrc9GjlwEeLpgcX58etzAloMJmFPZXtE8WUGT01V8+QArOeBvqJPS61PtJp3e
+DENmorpDbDpJ11PwgLuHBDq/WE5E90AKN89BqtVhONox42uzEDr6DaQQDAv4+gU
YOITLsvO/2Y9aUTUc3AYFO0PPmKIfjZggwJz9iECK4mdZ5iVSpu8upqVyt7nvSIs
qF7s0YEiqbTl4p8EGvIbI6WbXTc5HunyLjqF8cQIOA0d/wLkUbUg75E4bLnTlHYh
b6hegkCPlgPPLWEy71X3imx2mvtKLJ1DoZAyuz3Q6nzYqH1RncCWIbHshld0UjnX
buM3zJ8+XJPwtxjzKhBZcZKulGO67FGyh5EGIeEtwQa+xD4qSYjBFM6NGgeO3lBf
izJHHNR88h/UQ31x77Rvrz4iQyjeHRk9n77FoLJgbARtboJaR6J+EQHbizA9Cs9+
wTwxaIT7hqS1R+TBRPHkJPorGb2/+K4bdu+F+sPMmH7V+goFDFc0Xaaf7iGsvkrF
h4cVXt02birnTm8bq7VI1bCi9/9H7NNaxDXUmJ72wDfeUJI+6jf6Oezr5v+AVZHL
cJTFAQazr3EJIw2U5MM8nS2nGQhtOHI4EjK6k31JHgLjoimDLvlEatc9BaSm9yeo
3A5knkPec9bFwifWyOi1WUZRv6eGvkLL97qw6ZiH2uAdREWAYvWQZzmL/XGN8U3n
W8v3QB2zKCtTXviNJgnOhS2rc5E6E6DGWJmZ3A2Z3w9ebmuF+K61TniqfJWAZq5H
9iB1eZYtTkiMkuDIMEh4rKTTB4W/6eIoNOjF6y43SnMdqDRa5waAZvyjWozwycDr
ZPa89JU1ZTKfBruHybUhYOlk87PJjUflWR7HRrakunSjnC8TOou5wzahSQJI33J0
Rr7qcVRFXwCtAoXlevTjFGlBcNLs5S8uOPDeYJNoml3Uj9XzRnafn+f1y5H3LdN/
1/8sffVFenD3OqqGkU1qDKAtBA5GckV5FT/mr7BbfG6YnEQbhcUvFES1gpUTA6fl
JqzpOQTKsptiuAv/9UlTIdvStBEF1Y46tbCvctuLQNLXF+7ZLZUpDVaiKgJ1Rjek
PSz7gQq1i78czuuLUpqCSkoCFJCnjp0u6q7BvHn5MV2dpSix5JS8ebxXpeMKtY0S
007UEjkhodSQ5A7AeakhhnTwaw2WHBAhodD9iKGxL0EJ8nW9VBWmnWhouewIYrPV
xwxrbUv3dacLXGnT5AdtnjzLsVF9zupXUejqeWvjoSmZSWq374IgTbEmqH/SvAka
g2Xgj+FNrkxh6xTerZrsBNX8jUryPKuat5b8HZYS6krMv4LCtXvcyy8g2ItjCAgD
K0OT+56X3MlOxDAFw0lp480Tusf4GCAhSYOcFehYdiW+hkSpu4mVdhHOLV665eGo
ez5xXcd0rsLHOA6oPX91aIN8u5LsdGkT+vOlZgTnuwu4fquIo5Meaf0Zbe6WAZIJ
1XfxEbJpV3ymK/xEzo7+cvrPGkkwAuVm3odUMxoZn8GBTLRcHE6EL0QJRTIoC3Rs
7fSPNPMh7m3eBOJkNF/e74SCokPSW7RoR5B3iOKSGB0hwAFZ6Qf55Op9JITh6c+q
t5isqNu9KOUh+EgQW//c/B0dIrhKLicvwwytYdPx2J2KNWDIe6jVxF7qqz3OyB5I
gwfIB/vR2dsBPkNumsksMUSm/m1IM8uXQ7E1CKjEQFvgclKUxRcWJVu3iVjiNTXG
FiO7IRgHj4NmwftWr7Yizx/QJkGPF5sIBml/KPgv90goxwhlCcouqHlbv5DYFXFF
YDLUnvgvThjWv8Vkv3YM2Cxf8qwLuFme/r49UFnBn/SzVy0bVFqB8PHo+vCkNlVV
AZ/msef5wM6A+JGP00HjugpjkHgUZurOlyJ7ta5O2AqPC6HhhDeDmz4mVDiapyiu
b3lKFENJ9R22AnJxrTkYB/jHfGeTEmZhEV54Szo1q2M/xm7Q6N1eclhm8OW0jyzO
mRZN1bt64bEt3Fb9KP+kRQd8edfF+l+kJJXrfHHrPAXAoJ+Gs+lsJdsmhGc42O3x
Fsl/cWWt6TPTmKcHup1JzRynO+spgydmAMsQxvAoVBdubkMzG66Xc0IIdnR61lnj
vdNdmOvNRbGH1wDv6DeD50isflYlOJ9VFBti4G3ON7ZpBQ9HSISfKsTB7GGPkK7w
WRAGmGmLgBIchYnG6VeP6wkOjyBMXamBXHzZoAgiXHVwH3kqBkAW129VdTlmtAZC
us34pjVyHq4l9UuXPk6lDovZVl5qwVpwZGbQ1ddbalFvA3mTgya2RUozaS9vCbTK
WMD/AvedfGW+eDoHS/7GgQHpQLhEkqkDymIgZILEgwf4Bgt0WiyTv2kCQ/nKTiXX
kmnh02/4U2NHyU5yjkvDR0eTRSw5bg5w7KyBXCClP8XGw37Ck2tjiXXBuoHmQ/KI
dYBh+rpsC+5uZq0SCvnmgf5DUSqdE+Qt0NW9CdvPezqSC9pG/CdT7ivKm62FWJ2I
+zdI7HoqRuorOww9VyBTFmih8BzcbmdAQVYFDUbttfgPgtMmlU5MM9IAVc9F80NN
CZIO1gnfDGfBAEt0EH7Qj7F78feqDayqHnsUjVXuLiHCTN0Kk2CuWsxX2kU3s060
j/888ROCLyIrCrUlYV920SqeDnUwofSL/cso4GOOGan9NcKVGr54tSoEB/6UdxSK
vzpWxs21LuxUzBux6IVY2QbdPMCsmbZJi1IPuxFUDW8pvf5WRoVF/vjgpIuVvQzq
HpF/ewSIB6Yhl63cYIU+yfmmGpv8DNhG0sT4oUoaK+yk/DnK8w7jPhPLyQXtgNZW
pfLn6VCwe6SaIO81WjGVe1WpuimzskkWd6czMikxp7dvwCEGqMavzq+jQYRj/fHW
mLQaCDJEsTF/FU+y3dpc3Q8hahJb/8koe93fn5uJiCR2xk84LDzCmjxiK9IXT50X
s4Lp3Wgz7gYKTpnHXf9PWh6je866H9MnDSx9o6Bzr2QWU9siYrBMgVkVS8nNTeJ4
l9v1Bjy/Potusl7v20tG05dZ0qS/bgizP+08dFAmi+KJ7iMGdrq/9LhHcoVig4oh
Qz0ECx0i6iLKv8aQKNf1p0B3eIY56F3V9VJSqa+OHV7JV/sbEW/AJRfofedtakBk
zZbYqeE+W4YySWpeLsEFyEWWlEuUwkOnd4gxtW5rdaL5kIuD2HSTf0YpoOSj5wwZ
hf5EPpXqPiW4CqrpvcxhH7LJQw5z9bO355hHdgPxIiO2CfD7Viyx7z/DxOKuHqft
+p62EUfq5/TFgccobIPrOWrj1Mt018f0p+Dgju2U43pqnZYF4G81NCPBHDuEwEkI
xK9svBoRhPZsI7DkA5z7bl3PKt7j00Q+eOFJUd20BkYRE4z5AwIB6VnvKR4LWAPQ
g6fucMNEcj2RAHLa18DdQTpzCtoCvJAWLLQntGyDEYiD2zGd7UaGF0EUeHjjQlXl
yLDmGm4JVWo5VTiFkFe1hQOpCUH/h0AeO0GLLs2eY4T8Q1wTP8X6a/DaLWop6DbT
8mlI0QFRfQmzprE867Se2L3/u3QSEuMgnKihYAbd2AIysbLebvWnOKKTUAJa76Ui
euhPzoU/wAIR5GtacK24VXF8k7xG3LjAMFl9Lz+qaoIudCTegy/Qt39x7YcEeCpD
Hr4a6mbLiE24pJdt8p4HDMZWOYs2/DwEeHiCTfQrpSXHcr2I92TMdpZW1PAz9/qS
+feUYXlUHJkWo7TEnoNrYwaq3i7+DI7NxgP1aMAgvJebdYPx5fiSyhNdx0ULlmol
bj4XJa3BOhQfSd8Jv4OoW+vsyuV6j9+td3ldAT9/I3zVAgh+oXIjas2zsy5KTrtM
QNB8e+crbNNB9s3+gKkFYSB8Y/1QexBJvgHEPif8UfR7XKlueBCVW3pUwJq/N5PK
WJSXx5ya5wCdsOoTXph8XR6s1pm0+wK8AO+a6ELyCLSMF6P4g9caCqptzU/mzAsT
tI3eVEiYC1IkuR2pntxUeg2i/Xjg0hvT4Q6+BdEzafs0FXwZf3ONJyJVbkPuvYfk
sF4Npf1M9jQPJqN+iLlRnmoPdvFonOBpHgiE1nqOrEPIDYkBOsijGs9yCtZvAZUx
noxkPxQAbi9zPYzfNXF82VNdhdtZuwdNFO8dv+hUISN+lURwWQ8qE+WOJA7RNvev
zPjlOcKzE6Y4nwNmMdPcTO+h8WZxGfkQQ3fH/oHrGz5RCO0f8jSgVmifUVidPzOA
ARIScsWDJiehhBCxUj1YrPw8lj8mtP8ktrJwnyEdBbLiESyoIzPHh+MpzcJCJXX7
VKPtwNrPqqUQPy27GpBVt8HeodZYrikZccvcWr/+xJRnRDeDHpzhSQim0pwjszb9
mLH6TUKBjiprC/IwZzpLn1AMymU6S1FeBcBJ5S50TmDWtwQxomzP0QUo8GgfLkVj
E4ag/MreZ5Wx4mRWMnRW+f4Z+SEAu6DrEo5KIasgewqHTTxZNC1dK4rOihpnzJ+r
Tphcoxgr4JWo2Pmx/UmNrlAWQ5f1p1i8tZ6IGteIr0uxHg2S1v3ojYnS2XKHnM1R
5RZLI59v1vIxs1UvehqFIy+lErKtP+045DZWQMiGIXnAA419C+ISLp6WeVn1deaf
tdClDE9YyCqaNGiRy4AwvTl8OriK+45rKTZbpkiypoJkYHGWHZEWCElqi/gX0mPO
14MswFERM7cSelNNN5qTPqzm2kP3sOsLdr3qkf+M+n0OGm42RUG2O9N247081gQ8
YhR0wc1g7U9tf/DkHhUbFJ9eOpYcur+NlX4NOYc7aG8y0N04yibJNF00QBAnBcBf
u5mdrqWSBdkiPmDb+lcVowE7lCVIPmnJMhtvyJTPaP5xJudQi5R8Z0lz8w651Q/s
pqkHY+BFRIxpwJWya1wFyApCgUYGXv8r5FGEXFDqnCyLBTxJhtu1AyKaBAEd6rSZ
YllBqyxs381q1w6Pt0bCNbfk/kJdrOsx38+V4A1hh5b8vWFSZEBJpLNtEhI41N8v
1+dtkQ5Wr8b+yqN6dn7nqGM/cP9akGbjcJgbyZIuS1R9WGy/lWDbNKDW2Y7h/st4
hRE2UoIiSh+rLAMwDKve0sZ1RaElmJeCGhIl2/R5tegUVJCznUnVlqeP7rFBWQlY
txcjhHFskUuZrPcXhp4YTJb+XWqUDl4cZV6YSjuhg1/D729N2Hj7UlfgbNKqNtab
kqqy6d1nfaaY8No/KHpjSEDFnCXPQFmWDOI8TzyP3tV/7Bhaoh8s4sZIVHOIHfyA
rd7JTmZc3fCiCPqIr1TJhI/kps/lVuV/iCNPhhPZ+GuZnpEmpcTM+9Mu9Jqpw5Fc
v6bfE9iSMegxC5zPWu5cdzByLa2iwvr+dyYlpTHEjC47xa70zIi1Ez4xvOoaDPU/
3GDs7/2QAVIhfi9OoAbt60YfCNJYiUVvbID9m6UDrBvGvsTyTBIy4yi3RUHWsFHE
4dHF6UwrnrPfXcFL2FFNaW6UiHLphsOorXxhrxBh7Z+8RsNxg5c38FPgqcvBWsQh
haZCCCwTRfTRiX+Yw0CszFBo/15AUfW0pPfbKExf5KnhcPdlssjowE1l69wTnWNH
CEy0GrBpdl/zR+rmeNJgit4ZxdKB4ocFrCVjTXDkiYQHYmX0BLCrdvJhr2y1QJWe
rV6KWqzgr/WP5o/uRzaTbO8KMRtc6Fdbpl/+4f/eltsftDko0mN/H+92pYWM6nYX
/52otbbqsPTFbUay42L8sy6c4aFBSDtPhuqGcBy74mFqqT7LFqoDGVU5geoS4l2h
fnLsViNkGZ7Hr/77W+GOlmGbCtG3NGdPBQIQ6HKATNEotsDSfjPyu7HhI4KtvSXF
10mCLFmQvxl0+22AstuKLzM9PixRXMBVf8QdjMJrsq4XFRh3n1g8p+JMstqEpYJ5
oeILB12C3mIiuBkxCMA4Uz2v618E8M/kdqLwFR20uUGPPTSGWtWeLeAecw0nsRQy
rcvRtyMpp5IOQEdOs8x+YrXM26WlaVEwWtNpuRsKUNxuAV836cNMGwh8+QSgT3yd
9mEROq4WFHQ3lXftitZY6XjMDKpV2hpci+ee7iN6e/rwYiIeh3Pcikw3db8eVqrR
jUeXq7lfa/qJKAidpmYIhzH2tTvOklFHVTialy4bWxFqspIAAEM8j2/wOrcXenVV
NdFveAxta9/ofZ/oS1EToKzHzQTsVtj/CB8W2TpXh97MZMCl2ZW9M+DeNwEjLSNY
5mxiCAr49A0+RpxM9ESn+sUfmKfaIO07fWCpBq1sXhTp1muJzqfoffcZA4lBrjBH
ouOS3BjldjxNT+LXeHjIbEUM0J484IfvPCcEdzyuKiFhhUPlAAJPWWRUu4ctED59
5u/MflSf1Nojbso8b62/vCf1IFA4w/8kaYzRgDapveyFqz/yEr63P9Zd0/Psbu1K
PmyoHa10GVKY9ZsFvLYAmGYAsrakBPSiYwkuhgR0Iwu7KDdleWetZHVOu/7sOYf1
r9hP0VOjIuK0VC8MfKmS7IuI+rK3tr4o7faJat+IcZem8M72xZyrGYh4Jy6njSIu
LwRIqmjsnKEkWj0hLs+h0c4t27pfe0TQS1DjQl8/PpgvwukXHn1ZoqryAdgFmn4R
QUE8gLbTeRzk794KwKoSTC6bq809zWnCN+dTcrgI8fEwuDSqkZPIlTq7OV1Km7px
bW6CMAFX1DofNajBPNXhP6ldRdTRNPCBBqhL8ygmEnh1yRaFuY+uAQ2Z5hGIc6hv
GiDZDnyRcWObtCunV/tMZo9C7rqtJglR0ZGmbCuuJjOTo0mihf9omAD8NY2F5z8L
gb8dx3BwIkJxIQIRB7BHb+4pnVX/itoh91quF864EIoX5peodXza26JgPetgkNcx
cLOdhWO8a6RpgXkkFkCyczoNv7G8MYV02ptjmadEcVEwBo0+UANOF/51NT8W9hfE
cd6x+LTwB860iaDe58J7J3acNBagTHjLWbpTX7fuicyrELCqiXyFal5nKXpHFBza
SjnhRHGJfORzDnTVykXnW+FH5DdoMoOQlHTDfPmcOkyRWQGqR3OAsk33GLHemTVj
noX90HgR7YfquXzPhWIeGA19eT/Uy9q+14Dxmt38ONLygytmAFOZVX++82JJOd3D
DRxGPnEONvWb/tCKylsLFoF8pey7lk9BBNxerYsfEXxhkJCqYAhYcyxn05nLSdtq
KqacYJv/vT1mdU/TgYdPNRrXxRHYWrqucQpMkwpcXwyxekBrCoon07pHANSrJrvQ
LuDOFo4PLUaM7SOrcPRfaB/WAm3JTnLm7ANpSnXqD/2TwkpcHV0u8m5vm5hkXhI5
jewMDjLwT0EIfZ42ju2TJnMP1uorGkysTzN+PeKJl5lguOhZi71nPXN7ayupzoDo
wYm8SJw8PtHs3laJCyunqN8FQ7ZoZxByBDkSPhBdtfIFYpdVFCP8EtNGtILPJFPJ
B2iikKFREbIC20fctINHexQWybVOMYv578a+YxVfxxpLK4elTTQ8rb7+Bay6I9/4
eS/8dtc4wLzLQY0nByzCoxrByzBj7nsdkQUg2jchSPUcCzUL4wbRU509ocGQzbDX
1ajn+Rd8yO+kAiMfD6w1zg24lHOmO/XWuc6wCATmJ3fJU7xS68LIsK6AnMRxUM8r
IW/omKDsJK/No+2r63HAqJI++gkHAlWoVbyPlT/gF75joG3j5GQdSxplv9DVznea
g1Sv2zDIkkpPuFnmeVM2DAn1ifFsWqPefeZfVl+UGyPUn2qe0StFepfvaH5xf5LS
VwiHnRsYP5t6bHQFvfcLd0CwLV9ofHNM55pyXXEHGD4uHHffb2q6x/qzVAQKTA2u
ME3MVtf/HXLEcDDh2Qs8tzgdz3p94k1vynnAfCIM0z+2SlIUKKf5tRWIEsCINLzU
F+7SoWpCtsiAGuKOTTVMRuIc1DL3CzfHZ2QZjmF911Va403excyoKkUmb1tdMnbg
J/QK+pmyYsGFLNFd0Uy7IyMcDGiMgNLHD8OTydIK+rUCS6uv0sdkBc13la6hNIPR
06qVW9wIkeTY8cU11uXIinoqgiG4bJ6JtDRVLBZZ7zXbZc7Uln3+fW6b2Wtyv9Oj
1vJnyTzy4ZH/hgsUpk/2+OPS2kX8uYRzhXo+OfeaHsfExIO3jAXVTeuJigUqnefp
XhWnyUosSkmyCpJaPfzwAi6jtG/VD9/HICsEwIwDq1gqxpWDzm92vf3u8KtgOm4l
mENbp2qGC0LNB6RPR6HotfQ2YeiGcPhpT3Rw52SoqvVmhhPwYkL5Fotp3quqkmUK
3QVHqbFncw7GEw2m9C8Tmbe9tZa51uBErMyQpybbto9W5t8sXLdhsezApirlaY3L
+Dn9n5Da4GxrivIw86wjwMSVeSmHAHeudMQC1XWZXSj25PWFtbE58kh/2tR8R38q
NHQrhetp3JyFmXOcaFJ/38wq7tWzTg5ZTSJkImiKtk+UZ+YwcegOnin8AYn3d4Pp
Q9pLtTpzzTA8NpTw/4JqMU3Zfcighdy/aBDgnx+qEasuP93wsYwNUdtpE418VCzP
kADBtnlyDwBWF+Q98eqHMIrY8CB9ooeC7w8pJr+biltfTbarsagVsPRJUdzwiLPn
aiWZtIXoNk8ihSNvUPJodlop/7d9pQXN9aEtNUj7hCQ+zxajnTEURP8U/GI2Gk/k
PsEG1gJxVmrd/drtP5rWQZ+c9+/fL96fZhQVz3MkN5IOdzDyZiOD+RkAmS2h4rrr
aa+c2nR5WUQ2drh0+mFvD9MJYmx1i7O5DWDcvAS+y+6SmkF7BikZb0AZd1UekXms
UtycQgbkvUSXrNZswhTHT4Q8lEZiF1M/48FJ5X5uR54IFWqQJw5n12ZDERHCw+hI
iP69ZuuX6vIqYQ/E+eInyzkV9vin2neOKPdvIZ5DKAmOwg8Z31Yb8yrTz1GwaSIJ
gridzV2AcipIcj8XdICTnQ0oG+ZscAe1QHO+9tgrnxeE/sn64GfNwbXg6v3Klo9j
ET9SEh3sIVodRAeryvN6BNqxAyLEf7WpyPIcQHtjkiUA9BYRPLJq0388Zj8QSCL4
7h5+tsWpnuagBOPUaVeivBFmiMiOM5xz5Kksu/n8RZ8HR5Y5XTRZyO+w9cItn9k5
2DXrYPwZi2NNIUTgRn4RNWgCdWmk18GkAUC1CkaLc7V7FA7XE8Ch/P4M/ziYYENk
w3FVbBFx1M7qGs80CX/bsIp3rlEtg8NGHo1uxjyyNZU/czzPv2UvRRhVRCjK83kh
8R1xG8I8COIR38y4dPNIYiznzJ6Td8YXAmnOC5abuTxTawQffqYozQBUI03kEy8G
khk51LK5T1+oHZzo/Rx2zUWMuMZhZBAEwX0ebXIoTg4WpTwu5t8a/j3TSda2lggN
lXytz1pnsflFb+PThGEuXiNtecaA2XxP/nDRu1wBSB6VdTMXADwlu/RDsRT/8LTU
HtUA0hxlQwheK+vXwXRkr/Y5MloRIV72l/tLcQXCWJaR2na9AVaa2VxVSio0sEWs
NApWuAhIso2p1pZ8S0Pe55Wse9M9SRMpZwS12HcfPGF0U59qur+NCvPswnDOZBui
GtDCRqYEylZ5xO7IRQ5XfvwrLOJBEsfuXjiFVz8WWM7Cia0M+sk+Mro78XeEemZk
rKV9Rk642g1MR+FbgvAB92jKF6zqTdk41mK4wNvFGQpMm3vABbr2DMb+j/3kiHB6
7bat9D9tzfFQ9yWcTLGOtKQpRd3FuuyO1uy6nYwCUwL+ExICQoyw4l92Dq1E1mVY
6foKttvzkcuwAYvVpn/jklqDotqO8IVVqPGGopWg5UZyVE8aDKK0tuZoUN6CMlEH
xP52BCTlUuxbA6EA7PC2YVfuJn9foOBipA3/88PYIFKFyLFmu8JrqRNcYIGO86zC
YhijE8MqUXlG4ucMKfagSyBYUzpGskPnKbEgZayvTF5DFZ8z6UesFvIttzmSffed
iIMqa8+imiSs5M4WcOIbxYM3HXanhbMTkDIVGxDkzZqwdHfQZgz0ruTwUTlsrrlV
4OwWIvZcYPfi0qOztMFXP8eby1IoNjP032kp7x3WXqf6+LHOTjwGxpA8VJitl5rx
XiuEjz54Mm37Z9JGmwuD6hw4NR3y3B5wirsZcbxVAsytfz4ztKdRfW6tdqVzXNNU
pcwUJM9QJC1PZnMuGTp52fJqGQDRcpAf7uqWvu1NZJejtZrdFpbrXY8xnL58KzJE
fXlWgyynNAcmbUUOzj0wBa+zpBs9w1ZHeHTztRooyAP4nk64yPiMpRBPj5y2SQsB
nXMLMu56kAZFzpug/qczuWhcClK/Cj3h5SrHV8gex24PsIGPLpmxfwOIMEoXaPm8
cvfP0iy8DSnhF0RaoslYc5ZNisGcw/QYtq5H/t+KyKXfgOToiQdxHXoLkDTyBlwd
nGWY+ee1pTHQB2sblHUzE4wfSNsYgCVhZ6XsaO/PEEtK7IU1fkznHY4DeyUtHVpM
+V37JDixVwvwlujP3jFiocT6soQrEGb6MVEWNWIzZnfYC62265jCKJtI3Y6E2OZ7
gCBDLpJQqHzWh8vknmE6vsm+2xAygCsT5h8lJOdGXcwEg0hLK47uFM1AHaq62xma
BHJy4qD38SrczdmFZ2s29Pf1VPJktYwLtShpgF5J3l8BNIcNbq98VQ5nJatP1Ck2
HD7UE+7boN5JD3IdSIBrnw7bGYbk56q90rAFOZfOk3q626RMBlksQLwOEnOLA0ky
E4blHdMeo7prDYwX8AulcYtXVCJ0KB3WMglgE8Aa2ww96YpDbVPWDhDgvqzxLWlX
O8/zqC7031puCDe7+JTsqLBGwqkpSFWRKeFAkvArrO+qMFOwWmg55ekiQPasdT5+
ZtaVvgyaj/92dZHXV6J19hqpLl+8ikHGkPoAerslocd2WfYtRrGTaeodQPD54hF+
6mAVaW9jS+UkNJn6sQXzw3jRwPHUoYBSyyLAaateLeOvjn4A0kbkcHKiPCF9TjZS
9sCnZAbPBPNaove0eDCY0n27l9J65aLR0JrSwPMfvLqUKiaYpH5MH/A+Jo+g9wmY
OrDtbLN3Ntt6Bf9VgCPjn3oLjG+WSNBvGa4SVywenQUgmd2J6x99GGdCSUAu515Z
1BLoFeqrxIFvt3PBbQ7yWuAcvoTxg88rI1GMZA/QVfCaoHlW3WzBNoMaXWhuUvuZ
vxnLu/SfS59miDqEUFumewWvH4aerspbaEbwQR8ewsn8lbX+N+uUwiglRKQRoBJ/
mH3zJ/HEFx0xMQHgAenR00uOZ1MNww2NFnPfpXuWRnJ2xiEgyyyhTLlb7IfoiEf6
Z8eTj3y8HG9JmbHzJCNhWsyIDVC/MrxR24PzFxWlWlAvmQXgUEtcJ93gBDZ1/Htw
oHaW4VppJlHX1pjWqcFE26XpuqZpLYTcsJqBK6pqOmc41GZqk5e/JfHp+XopwA3s
KqU/dnmHNs8ED64cAh+xeF4WEBWxc+DEau4126FbT47LHRjxkav9Xx/PHj0U6kV1
7TyArnZG43PL/GZdDiZN2vTIsnxN9l+HnGdW8jX/iSM3VdgdS9Ok4gifd9SzIEXD
2Mpe3eU9Pfphfmt7yBotBt7/fNVACtLRo/19C31WSzmq+LmesVlbQNloIKWg5TTI
LojDqYUJ6eBmG2D0/tmG/i9MeNapCkYZH654jYYdl4eTEqwnPOgceuu5q1VqnYq3
JdSvMy1at7igruPkq3UAGhQmWw6BdB+46un1ML0Nh4U0uw8KdogjcTwZmBXjr6IF
V3GfwJ2E4RXgNQIqQ9aTQHlnqMINSpBTGe4GJ8G41uC7OE63sJCJZD9tz/mmsEuv
77RRaZkdzxuzDvUmFgovPy66PO7OL5X9ImXnBQp/QNEWlS7SHPfRbDP2J4XS6v4k
/ncvjcZmI/XzjRM7PfzTeEGeDpAGlxXVUxNDGSYzXCfy1ToMsn5cuMl8/046l/O3
MrIRsmekD90HNeLnmgf/b9UhxMxMnbmB3Hfkyc1j2BhMwhBSJlJtP91SoRt3qrIv
CgjaRy++iXvZzkl3L81mtao2z9G6eakcmfTybdFbKYNOFnaYvythCQaDUmtYHpFK
pITBqStxZ4nUfmMCR0Pxj8OmF/vXDYdTa6g0yUF7xkw+Gmks+0A85uIcrW+jI9z1
3b8g8IAVgXwN58jm8TvVI4r4GQFKNAFestOlF6S/AB5rOm7G/Ipr5KTewHuj3SpC
iWYnMZ5bugru8OYq3V6lBbhSUr8MKH/zVtakbqq9RXdXp1q8QPXg02MXR+2jQQz4
mihZQlRwN0EdsWXsv/2XfwP3nz3ZiSFNhUr4AlLxlA9307lmwBMmH0bwh67BimGn
B7iHtPre6qHAp7GXZTGq8A2Ux7jvca/McGudSVxA3ELbaV1ZtuRCZmkL/EwnyBmH
fUgA9pELin1dGyQ9Kz2z5lRg/dSoBhEr1uvkdyGD2y1lRjRxsVPT+3Pqu3P3aWQW
+aPnHTp1w+Ro/l8NvIqH5k+vBQCf/sinUW+c+kBjm7pIn6u5O1Uyc7cb80kaBjI1
OOf5VDjGo/NblMqqjgynxoT8EQMq22AQ7/25Igjh43VM1lObJbABm6ADFlHxY/dG
fcUCrPx7na2MLSHNqcOplwglXhrq5i14J45r2ryUbJ+HuKTpuywen88T2StDq2Sw
/UvvA4f1/g9AD7Iz5U8y2FJR9svk1/AhQHL2flasZau5dTofHsKIGP/UXhInoXU2
BloZUtzlPoYR9og3XBaky2uXXTQ9MXLFvJV5w6hVmSBbZ8Gwi9fceUghC73YvHDl
8tqWmlRv8T7/rr5xkBT+7E0zNyknA10m3FD2c6KbKku1XZCR/uDH1Dr2RuCjaD0i
Xj/KqYvRslWm7B7qk6TdSdNkWCrwNtafGfVdAKCXx+VADniQFN+RuMRsvr5xVst9
W34ed29pceHtCiuk3qOEqFgkAea2xHwAaS7sKMZIfmaQPLQhH+0DJts5a1f3x3bk
vbjE0/nMYrc4Dbavqqy5p5xzCtk+FXC4WTUslOIqfvTDSoH3Je7Y7rgN8lc10P/M
flqavgQyIvGu7RSRaHucSNTKcCpce6LwciwxnkFJUtnIdleznm9L5Fu9Y6Ek5Sq/
xxt9n4cQNGeolBuB3/AKjOFaFCMjJd/afo2ZgpttlTjF/M2bRmwmbu/6FIRosbRu
8CTZ81yXc/NgPGZSJI0qqSzvOm6G5ox9XNdU5nutOf744dsW0QecvXd00pusMG16
IgXVab84Wjr1aB39Z32KwJ6IWdn80ULT9UHX4O4/loDkP+PSMFR18TLbQmFys+L0
yK3/8SR1O9lm7nnCjTD9YYpuJ1aIo5jlgbcJDwZDsWV4YTmLbjCDPwptX6BeJ9pe
813tXPupvcKBugYfBieOi3rFPEp4/+7alAaeW39LAhzAWe7LgXOyGGzJt5QeshAD
2UwljYt8q8K4Ha2woRBugTICGA5/wdAiol5M+7oUKZ85HleQSxL07yKTEbYR1ets
VFk8m5RDfPpJNUGFVoFIKc67MWxymCBAAEOWTsLszzF34gx0bYPWCAxTRGg35k+8
v8yrEs4W/COGNGMb5M7k5JkCVkoVr2fw67xwzyf2SkmpDsc4RllibGGsKjGPa+V6
CRMUghtr1cffUBqUUfkpYCO6U48MrHDoK3nzalDvXWuZ6Vvmls8XBOMNYQ+bOFgj
7ojhRzKSc7oGK6UQSkkckxUoK9Kv7HTWMFUnJkibDaEktLxk1PlqpfunVPJIYbgv
jwqTMooHQsJeLCGK97ySWNi9ArgK2XHMm5As9x9V20HKil+++sUwdt/bLgFZ5gou
rONXox4NolBATt5fZcqrHLtm4S/ne1OfYQoIOXBe1dTDmlPtM8fUBH2/CkztdSdC
0ZpvJSJdKXnGSSzIn3hb6ly180iIIg8i3gEvtoud4xm2pCZrquYsSZa+2y5XbVdb
PE5ktZaiG+g4Fa3o5SGPCGYTfhHa3iJSDxxL3SueDUvGWWijvNrJnmdRK2S3b9XU
QVJ3B+UsdoucZRlA9Ox+kpta4DJ4L56vPjkyRWKjPuPgEgADJkvD46Acvdt/IB33
loCmPPytWsIPXL5orZwHf1ku33VwC29Fc0qN727CC872qIRPgRoH1+KYq2GSOLWO
szQSMmLcBz8Y3LfgcjWh9kMDMD5nLT8mWkfupSsUwE+SP4sguArJnxZo66tGCxIi
/ykm0gQz5nsze9zLG53tAskvoDwt0WMFEmrU18UM+OAfimqo0i6Fq+U68m2TLLOO
l8Gm+UkKbipRF7IThZulEa7nl5djU/6U3/88dDBWwIiUbo9CballizvGrr4V8lAZ
vMLsoVZwQ0XGqBB2juns2C1jYi7dTQnTPNj8GQ2oINrFTlZR/lbhHpp8AaWLB0Wq
gly/IBgWkpdZLGruPhwksH+mD+ivrd6OOznDXwDkqs1rPeRoyXwYEaSWRCFd1UVo
qfu3KK2lJivUkwlZSzL0lHrE495pLlx+fQH2F8irHiDJ60VMcMhgqz69oNY9nCUp
WnOzkTc8lldpvN0dyiGxeTgF9gSFwDwaQ6cVbofBHmY0bNn40tyj469rLzCdIzoS
mHN9R5E834ItsH8ho+YDLWtxiqWAJq0RfofldvfDVTdOujOYJaEGO4wn0It/Aifr
pJIEH48x86XgYPYzhyzdY6OTV0FRrUvOLY6CKa2pJhBsf63G5FCG0elGTXUWmET9
1SQuspgCcb4hIiWC6j2xefuoxzgNfwfduc3uIBRbPzWij6qry+eD+kMTJgR1TdtG
Vqf+E4Dtup/g1r7AgFYT3i3maunER8r1IRZNbiFKstCjCABDWRvHwwu7z5HRrZC7
zxPxFsv7SIuwI8wrzFw9Omh03GkK3Nd7OW5sKpKvwSo+2IEC794kT7W3+Dm2XSk0
4dpIzKiZp1VGm5KXkbzX5Nb6iCsr7+wUKmhMG27q6YvHdpH8t960mYQEs20EQahk
OissRslgDg0SLBx8SJrz0nEKoV+2cMyE0VwYKqOYhH0rKIr1HhWRscDkQMlOhXD2
6mK0XsnPoTd9UtCMkA/vUcsVhxHmd0xGGqb0juBrC42SAsdxpz9cx2hdeN1uukmP
doxTQae7OdJQzyukGwR2k5voNR3K9SS2xZD7P2kyQosJahXaZq0DxE6uEx0N5Thq
8IRq+zkmGHU2GstscB+QLvfCOUPvM8X/juplwdGvanBUZJPjxtwDjgDvMjTrSaSi
bi6p6wrYhPyodPuBgnlXxPFiUVK1swYndd9tY+KseO9DUplSg/PWLQZquHY9fHsV
7rauJxRiefztnstUKq/TL88R1/TI5WmMW+1ozOtycAz5FrrXmkEkCCrUWfbDrFgd
BI9Rhs2kMXNYnet0oDbNBGiFrziYOZ01UbUTGO0DcJVPefpMcZDJ392rOHO4EMwV
6daBTmTvAdqD1FAzpsfFMNPNbt4WB9kxs/PU/oACwitUhoxY8ERQgZ6K7NjzKKUG
5rBYDe4DwsJ5rHezxGsflkcOeR3sWNHpi/+ehWCdD/eONOwNmdIQ3RBeQoqxWBe4
V5yEliIv+HfmHjxy1//9rrvPYPsz2RFdw2j8p38QqEUZTLCuU/fIkaocH3lASE8C
AnA94qVWYuGM0Yy2YWBZKzqQb8OH1bwiGuY5NpdiQd79ixS0e9hJHnCm7BLKf+cE
rW43iJBVVkjlSmvMy1z4rMPcpusbjDqNCzl6hFCnbvivhQCAFW5dYX2IPAjEy9Fv
y6HZSviUlurynNQexOx7ldKl7I18rIGGuT63e+HrocOA6OLFNdZV6r7gxbA2wJsn
VsA577vlMa4Xtr+7JADQTYr/B50ZaL+SQ68kV9iZEwfGxmWtkiik9ruzkLBswVo7
hbYqa6mIOCZ1J5dU8PRqAuId6mRva9yA3YfY/3hmq95qGa1rxBEONnyQbd+mHNKr
2d6EnmR25K6OcmZFEKxB13ycWfq7+UT1wewq0mjvbwKRdWe+TLAYbYzy8Jdo1TCq
TnPWi2eX/zB0vD5hAwjk9T3dhdyBB5THy8PTafadCByYj70nMEMuzoFsUYk0qfKi
He2wOk1Ho1ozXNhRsjZyI+H4J9JEGn9JQ0IX0vaDhY/G43OkygBEiyeIpg3eWAke
bMes0rs/XSp+1OS9rjIuZJpr7bfYt6k6+orz+J5o5z0UqssrUaYvfL0uuFkrSB/s
BUKlo3vAjZ0Zxyat7GaTFCaF29sn2BnAVWvdPDXs+xq2mAgbm59djzxOFvBHrG+E
06QWujbDsrIWNwQpKsA7Y6PbjQe0zDDjxAirfh7DfWiAyy7BmgNMapRBCk49xIHI
0fMEXGDYph2C8iwPMQefcc3iv37Y6CqLHjsP++txnQtnF/6k7BdLeYDu1pmcqIkK
sgbyqh1NJYKbI7S0aAJjFdcB2KjjVQX1+gOtHmowb06nBsFDMPW4r32ehRwkADnm
n9tU/FReh33MHoLiDz7zaCVt5FzhfxQLfFbWP+5mS6n5LVg4Fr80mJsNQCJD3Ury
37kPv9zATwEigmQESVlFf0qIWcfcrg4rB6J0wBqIjieORFZMUhHfCQWzfcFajsRe
Dg5ogAMy0ysfN1lAZerS8C97hkkgbJqkwwwV3y1Q6+87Zw/HCfMsktvjnkA3M8Nk
AIDtC23+V68mvDSZjHYl1iFM/5Mte5YCrXrn7udLyBrhI5a9xUvMjXI19wPfirFT
oY/4HdMgP7qwJ4OH1og3XBlHgy2vw9wonwAsL1Go0RqLetPJNywGQCmTgsfNrST5
wrRz3T+INRiwBdsVfRwrtHEtZwo0M9AL9ztPNNcP65tGHYv3gEPRuyPSQq8260Sr
BIZQhZAutG7HC2gt8dNg0acRMqpXKfIQzNWuUshr8Pma0OMEU+2YqYdG8fpOn28v
4s9uusKo05lerHQ4atezFmjlboLeVDbFXwm46NCBqFsec8U3Da5bNX8TGC7pz3M3
tx0EA24iu7Uc+Gg2dUE1zLBwBMvfIxUI+DLuDvXuY6BzlB50ZNCILyEXWaALN0wt
NXHvUrt7aK/cYCIacsfVD6NU+owAT7YS4zFTsnYcxSCzbcJqniBJm9twOSrwIq/A
SFRihUEDT8qCn/FOW+S0ktB4twRl0CkeHKHWXzKjhxBPiF7390Vgh+g+1j7SWD1Y
bYG04liDAEmwD85ZUGwwO5QowR/9Jl9x/mh0XpXO11dcgQg6DGm2ZcDZ4PDz7nov
BuBxFPm1eysMX/q28tLoelex+6gHMVfW8ZAJGowMInYBzaLaibXfbPLfWpkc+Sd6
Uo3Hbwnn+sOCqOXKCGNS4K9Zibrrzl0ukeRQneTVXj+1wvn8/io0dEekttrNja0h
jJ0exwCBDiHYWoJAxys+n13iZtB7E4s0UyDq3btQsChny/Hu6pguU4kR4COJ8+Z1
fqdlIdxo6SIVzO3km9j3/8K68LXn77NxnRhnVXk4j0oTz+ZfiRMC0x4kjgsB+GKK
lU1kM5KX28P6+mzMZvKaOf9NFzTFiNDE4KN4+IuS39qljsS94s9rGESxS0THY7zt
/NG+EfQX4pVzbxEjHmai9wzbXGAiv3ZjooDRxpTrVA12u0LlM0uQ0Blcovaw3kiD
hk55Ars2g1aUpgnieHO+kYCMBKPFAl4oPNGv1JAyOLysDA2ryF2yTvAx2Brgoucs
vwGgfkMWFYuNiB+KY/keA74sXoNkTp+mw6tVJ3twRelKpk9ndMjyfWmIszhPBBjk
UA0eVsqkvUq3idpYJJbGvSGfnFpjisd34TaZxUrHcSuCroPxft2PoF0rnR4vRei2
r4BYb1mB5E+O59a9hRtDLj4s+qhvUPcpgVv7oQjYh7BV9OE4OucRyPRjhqA5MqSJ
4CiJOPvkvVZD76DX99ExuOEwf7LJvcSXa+ZdjDaP2KQ3TvYh+RQNfH1aywcJFBvn
ErngN0hW6YlQ194X+sdDRbom5+r9JHhI4omKvjoR/3yOhsDfkCRDck4DgxVO4Ws8
qwitYOmJd/aTWpJAytG0heoZTCMLLRoN2GHbck5O6XB/EFthnbrrVC9TDj7z6cFZ
eIiFUIC1rNyof9CR593QIm4XmPqJ065aaP3KUbFs9KnL2D4p8bd5znZSPbRVBN64
RtPWdOJNvJpRcg7V2Hj5elNmDt3LvpEZooD8hMekqbFm9NjBhT4aNdEA1WqmHp+e
Bk1MKYfAEjyhwRKCHXXc2msNzFTXrOWmy6SIarmvBuvEDzcknydzHFBZvp+hDa5s
grO1TI0AphC2wmRfJPkqmGiyvdgIojgBH/VCkzO37fxazE86uGJK+uGfKTHATfHL
dKUhq7jWaZJU4bB/GWY+arVwx21Q08dizYPzWbPqdL9a/gO7nqqsGB10F4kyb5Fh
k8W7bJjJdWI0uMmTCNM+m/EwMjG1B2iyAU9sKDGoj5kMfUHXClAo0bSHFLPWUKSq
uFKvT3s0vIwgPGYqNtql/iNp3q/YrY+51qIOT3lP7RmoIrl9JRGZniQkubBT+aCx
lFC/kmoUYNKkI8ACBs9kMc6/3R6iSOOYSSD2nUd3LhSvs4ZNwRgaq32CSIYwqUip
XvhOJ05lWWD7tD+UJtYeZKhnQ4o22z3RvTupCMPZWgOMyk5ZvlgpP0jzs66rHaKv
vt/OtMxL09Wykjal2OUxSxMvd981c0KYF55vHjwtJALLql3nlpAEPgbc/wvdiCD/
uhBOt8OEENr7LW9YAmCZxgL8cehrYrEHrwDd7/hMcovHxrdN4s1aA4PSM+YKyoID
Zn9mZWtUC8VQSTDtdlIlyednmZhWQoOSoZn861HrvLf/K3UYMq28aYZ/4x9AmCgR
+pNhyJGHX5sVN7OWCpE3YiIo49EgbmbnWYu2Az1+G84dEUwob/Wy+wbAQkrJ3nrd
SwtyZHcH4iMyg1R3rsxVkOkJ7iu2yl1kBPMkb4YzkpPiZL0jlJV3uXHNe/p0OFBn
gpA/0MvKYzDb/QMgQXO+6byn9UDjF55IlzhOaU+g4ah+kGaBtmE76/rWit/x8Rwn
J2jcwt/lSwQnUAMMxdaDnFEPPafpWa+dq79G2rk+ejNBj1Mq/ldO7mVTjVoDHr9X
ryfGmsyOQ0+3vWL4EYBjX8/HqVIKEe7fRBLKiA4fkyKr88m2hXMianTFXf/10OkD
/QwIFpzulOU5UfHfNF0zHgGO9h7GRxi20NwFdrDc0djrlo9BXEC2HdfYPOJfmSn0
0MPhYDVmrlVs7+8s4wdn0Zou+cbX5qSniAgl6PRlMbpdugasxRLRK7AIf+7Yo5EQ
obLanabG8XJKFrv7yQ7yufR1oWM9Bef6fN2SHSMum6dchP72T64SmD6vWjgu1+qU
mBrlStGQHv5AQFJm8S8WwiGFHSK8IIZG6YZ5t668L5vpR9B7NzjpRAgek0j0XayQ
VOMPzMIxjUABt0ovaydzt4/uKN4h/m+JBtHAVRD6RbpTYY1Khi5z8V7OTfP2wDpu
Iorh7jA8RKenXbHgi3TO4I5hPgZ+1ylCEguhsxiiTvZNhct33SXsQno3GSxdspll
BhltJ5F+n8y4wcCVAfvLM4cemd49VqujGJ+Z/sZtJAxi9y6HPd1alHmRXqqMrpiT
+W1yCaA+2EdQBNnrVmoTM0DZAc4z2VwfiI2k+OGg8DZa97u29EH2xhvRqHgYN5cW
YhMiAL907rZSm15OQpF/a8QXd3tIDW7PitswsweW1dfSG5jDD/vj3FtAz0LLC3+n
Y62Vge9MWddBFe7SPZQKN4h/Xr36Hu/IH2XPiN0WjGdU3xUWqJyqS4DSQG1zQTA2
Hxx9/JDrYATQqGuQbO7N0uC6FytezQUA7qK+z1ONBqY4odIP7cETb1wgh+9gTk4J
m8ITjKqqxopxT1HFozttFtXtUZmsrs192wMf8ZYAJDlMRMOhHops8lOCvP0jY5Nq
ahMV7s91C5CmOzzmUTki0nqPbg4fSgEmEZby2+HcQDNK/cv2VGVOV2Q4UAihu8Zf
iD8rKbx/LyNagdGFYedyNlv7IyewoCrrCELXXwPCnXLv8FfYcZwSAeHIwJ0u9reO
9MMauW4+59u8axJLnBHl7g84JffUVCP3heQB1I+o8RUTMF5xxzxWjhLJ+XAbDdPY
AtP/AcIB7UpwFQiOCkx9wwPiEZSB8BYcA/My/zbH3uJL0Yc0zY7By5Ds3yjyw90y
iQdDZTAaOSFawIh/zJXSb4kP6j7dms2WTLV+mM/6iv9V4DlxRp0jD171vheP62kV
CtLmOnlwo5qibosZdE09PqRnIvQfu8SEtIYhFPUcQa0zdN2C8buqS6GTWxXzX3H0
aFTzFxgY0xkpcNODrH6qF4tzQwKDqU2YraV9HDzlARNOb6FGyh1hU0SuIZ9oibXm
Qj6YfOCsv1JKcKbztJM8yAmCb3n11cT0LbSaRiA4cE9H753lbY5pA+RNaOrizF5K
8gz4q40DFckYthnDL3w9/5zbvH3kwkAlyUBGbxKGXNAAVlQ8wC3K0Skus4+nMwjZ
TRY2jd1xh1EQSTwCYmmbi5QSoJ20nDwaDi6ol8kcBIc4ajbVJF44hTeUMnf0YBSB
vY4r6DfL6sMEP9R36cAPO99jNTSnAObfjQDkZC8FeJSBVVcq6vc3WBhUEh32/N4R
nsCLWJE/W3nDC6p9gwy1cicbfynkPEZ63x3LwAPhIG5mF/gTRdTw2i52+KiNhcwi
mQoliYV0Tm0UdQ8VxeJm842v453wAobMpGnbyPu4e/yDTisU165nTxLGi6MnryFL
TcI1S/NUrjeQF01IgCfgXpVxvGy9T2YeK4HXJQKqI/GmTuln03O4Jgrq00E+2a7K
Uz5LIUxhvwmbBGSAPyOag6ha/IsEVH2mu4P9HwT/BenriTeM1EgGIg1Qxfu7VGOV
hZlwGXhZTP2h+Z6gT74tGMfGN24+8UOBJsqPRgbGFtJQK6kiCmO+0FIhs8fJBH2i
etFebCnvp7xv90fFfJbMLDqntKKy0Sgf8o4ABPdSTgUQfpw9Y3yaFL1e5vyGj9du
/MRxdnTdNXvrJN08jk5zEWYp2yY75IooLTAY2ZbSDhkLGi2xoHdUW26I71U3LuU5
rQybqhEPhqlSzI3SD/5SisPwNswPKNs5C/TB5D+Fd2VkBvlI+gUKOsXcQjwu6N4q
3jBEQ2cRfFOQXJ0u5LRi8lkDjD4c+HX5aj/cXleR0ty9/ExzGgZh/TJjPwBvJ6gH
gPmmKUtMC+TYk3bap01myj8kGto8a7ykiPlzm8Zq8kz5SAayFsJMydlHISfAP/fE
7H/dWonL9c56H8ChK9qVo/DVsrjPNh+FBHtDen2P+Fqy9cr9BQ7urh9igwU1FRc5
UfawmsaOAQk2eySSe0bZwZrlFyX0fzudJK/9FneqwlWsCuMJcVY0/xudyWg64Uss
M+Xh2FlJVnbhdzsHKwRdtHS6u+4h25akwhnjgIkt73sIXMMEACekOElTQIf7GqwU
DSEGFM9SB+nJ3xj/cDGtx0x5N4hTqlWSDYuNx5qW0lwqvxsefJ6FBsFiemiAIj4d
OUgn9VpelvNrTG7GYEoSf36xXe0bTFgJz7w8hUtFYondkkme+WVKOKv4pTLIjh2o
a6cVd9+WXs6bU1WAyZdhxV5Kd/kCyzZ+24w5UzbrvkY0Q/QPps3XmNsNPKqDpf5L
lsse2Eibm+e4vNpx7NDc+nL27RbKB1h2zTmP4um2WxTvDw/MqT1PUoHlpHLUXgAZ
eHU32sd2rhxJYDALFSSmfh4IwsrAr6g0MdIQaK3il0NGlGIFikENqhxi4ZtnVp2o
i/rhZkRei2Eafe13afwnKVu8lnbmM1gJaXYYI1hZVgOj0HHV9R+H1g2rqLm9puK8
2f7W4lyrd7F+1hXf+6QLc/tCuuaT45aJeohYIf1muFYP7JCUiqhdraLe7OIJji/C
KHTkYS1DTLmatfHFwoPE2QRaH8C+40B3b9YO2sWG59jDG4d/y2rXVUTlyt3+Q38/
vgz9p/IVWRwFhNS9JZ+bRSq5dAfHV8YJxBcmAUcmtqJY6jWBsmBqi5bkv1DgDuvl
0vRvqE6bj0PrINZdgeav2XjiSNe1Pf57BTfOILgo8Pr7oAPAevCvnD/diIfjAKyA
raTCG2CEnkez56xQQ0MvZDY0EgRxPGmJ+HOmRbzJBkSMzFb9hIwcZnO9QPdVHi5k
O4rf14206lkF5HnBsI2zys7+jKVOnwCEm+uRB83YNzCF4kfBZ2hBYeDta/c71HFo
AyJPPvmsffn91auvwofvTToY/Olu/vQ9emd6HurlN6SgDZ/oeiZPvXQ5S5YE2GTO
BXbEisYN2UfbYmoFVcUk6qC0r8CODqmgBId+m5TehFmT+y2ghuBuFA4NjATArPZI
79NJ7DFwOHUQPTEH4cLT4MfdjAjdrGvdH0fr31vGXy+JrS+1Ate69QNOJZqiAyNe
xLXDOvHav5e5c/y6aW59Mi16mKn6F73BMTmSpJRbFvGcTtti82gmgow79I8XgNDM
3k0af0FhravY+dJgMgS69jiYVDxQAB6mcCzxUqjt5i7hUm6yKGkP5ytBNeYKUlvX
ve3zUQk8vLCNxzp5ziZ9qxpLtbQS1EvRu2HKlIDTHYOUifVEwQFckK7sFGKvYQtG
SPx9ys7gz2idq4mi9iGckUqUB5vaueORlWRS2emZMYc+r58wBOqFxwpipeJ/lTQm
L1f6CN5drZT22NovMj2TooNEZb9Kdwlo77eMu1xE+OLZIYMU+7XPplIuK/wjbayW
H83IstAJXMoAE0qbCyZWEY6Lmds0inWG4YBhEF197Vxh1qSXKxfVhE8B6ftpBwL+
kCZq3NUIWs8LmeA+Bwkj8b5OKRXmIRImPPQ5+rr7rEgtXFLmIspLPqMSCBYy8gI1
/KX3Y2mlxxHwePJ5O7DpoTCSAnZlr+sKy7mxCezvi7MdTuYNSRufekJbBXt+sVLY
TPTCE6W3U2b85lkc0P4wYFdJ1Gp68bPppO369zxZYJBu1pp3NpwafCVynsMGEGFD
BYrCRzm7/DPnEdSkLrMUfr2seUam1+q1lSmiyVC/vfvNzWMaC/yQBk3gWns5dhG9
eprFGMqZaXPmCm8edLDbRMU1RYFG0bZKnrTwpFpcOEQJQZCju1kU2yKmH4BqCo60
GmDlKZPzeiwQVXtvjxMbwcEdu0KBfMOkfHunDhm64/ojPK9ROy+sd3TICTBe7tcb
uq2LeXLASRa2IFru7BZ3AzUITqi9BJfUid7Cj5HAtB73GzSa64pcXf+bGtgASugs
lYnTJp82AGAhmj7YR/GMqEaC+HjBnwEkxf+dsL2mIAl1g09Ys1xemVy6jGdmFh+9
Gs1s6Qe79V08YG06p42bpqXVEX7GDQfteQdAybTvJSpICJ+2yiazSIx8PpkaqRgb
B0/K/WApokzuBN1F49zHpVeZHvSbS+wdua325WsJXnmECIxh6lHocpCPyQ1OSqWb
XodyQj9L4RzBoOZ1pDEc9cuKp0G+Jw72z7Ediw0NWihKaTVEIrZrVoG9pYZnfGvV
dwknZRTOVIY8nsukO/Y81uTJ3j4OYAL9/7+hFBs+1tbNy4JgsBgm8uH6Y2iXDU8X
hiW/OH6t1cW34YymQLijkCEmv3moT6s0zbivswLrirpwwudYRDaimHizXwbUxGOS
eS0c6diWWcBGMAcrPw27tIXcA7IFBWLsegmzzSYAcXpTbX0FR8vjRvfujSDlc1ZR
nEfqi0fXv9R0LGF3WHE+gg0tRGILvuDoaBlR987cOb5dbAUiC2p70YvIEvC7YhIu
Cr/lJZXSEx+zNJEY74JprWb0QLiBhf+i5/PmuzkTxd1beD5/lXvU+ihsuwxL/nUx
849PEQ3UOAmUAxZNwnYFp6iF4c70KZB8dHeSjJgoK0bCjjvRtanFn4AlF1kQMTtC
LzxVyujvBFHBOXfWGzsP+zL/K3xU9tX8UaCqoiCKzilFQJw10E1tBrOkb3zCtpXg
q9qeIdxEecrU4Vbz+d8VggfbZ/S5ZinH1oZ2dIR0cX+/e2KtQcvJo/3/H0P3VDaG
3/8hidtv48qS4Z9AzIptuJowVf0QjeVbyIO5pSj+nwvqMmBXsQ5pyjdJYGC/S4vL
Bpsm1QKBVVcPyCnzV3Pe8uIzpq7dpwNpRifYpTczgUREuH6Jd+13GubOjJfNfny+
FosCiNYI2/kKW32O3U/oncxHV4pSW9K8BRjabQiB/g/eH4F8HfNzhLj+khjNTc/I
hhlM9TyIMPNMdEUI5RiRqA+8rWZNsQMKAyf0Skk706wBUubBi8xdpWTrrKhxi1gs
lFrOu8RPEKrshepJuE7oWhQOrdSposP2340g+skB5aP46FUrxo4Qo0ZVhBHAZo8V
2toERwgH69k5n0NAxODh9xRUOUGjjCGz1ZRH3DJy1/2/os4xOLjmhKGpzNs8Y3nt
tUMsWe/PRYBo+XAuFpPX8K65/l3iAEIKvUWjgwZ+ubIA187ggFLvg0s1QSsUA+TR
b8ZHWYiDylw+/Lucxdha7fg0Jrg8vDbfghqNmnGbXBm/AfGGkZA4YodHaDyciYmZ
w6wDJbNqVx8Ca56pJUGrkQoZo4SDFSmGIvu6VjaFyXxcEpAXkeZBQWtAOqsP9wZC
Ga0tQX+demkvxYeLwTGa7fx7g4CZSvT/l1L8GH4DtpVgj06KksrsV9fsjjX39ObY
W99t8rnHvPsyHLePtFKfJ1vGnkwzfWLYbqjIfMq/wc1js6E3ynILsKTsKDSa1oHc
B9XIN/hJzmvNXjsnlpGudcDlDZHyTw7EubLu6fG8wfUcKcBk1Zao+XCL6QT9LkZC
SjCROQpmEFxtzmWiqlTziDMdKchJtACe62T1Frf5TzEr7Fok41ZZfOy0zOUx9u7v
k0HPCozAXaTv1t4tsdxuLKIkkBVmlpLICovXgKFqfT6RwNLnIAxRXOEXeHaTA5Md
2/2/3ZsB6wSAWwuXffOgLuiOu/j+VhgbzgE5DWB40uaaJ/gXHaaranoUoOyQoF6S
yFsBBc6yxraZ2ovvYXLQvq08Psm7YggYieAPyie5kLwh30Ed/ffh96PMlC602ez3
amoB/HiK1X7h0ghp5XpTIx00BEyitaC1fRP265B3jMJVVIXy5YxGCnfgAB50VkCv
O1NjdxLKZ/BM9IlTkt+bvxljpiqTuVK49nJfmLZOnpgD3nMaoQPWFKXjfjikiv6V
xKZ3ylD2aliRf5lmuVJk3ptt1Gtr8zCWCW4dq3zpLmMvzi6unwVPrvpBjQ2SQGjL
f2ryTrKsANsfP9w1iXbvjILKSbNJylJ3IkWZ70hv1+FQpIsg2Z/GGMmbAafjzZkf
eGQGSEAIP9JCUDLEdt+vQOI8UFJKv3KaeNVTYu1fVGeHaYm6b51qCqJx0aiCVlac
2HAcZz9Pgq9LvnjFWnnOFMzgGtYJ7MTFSyyZ+tkdSrWWaEPdDqa6OcTXhIfcex6T
25GGDcetiz96mELqeQ88zBTIDJmA+AN3V/sc+ISKX3vbOcXY6+ERCC0QJ22tgkWf
lDBVBDL4V5rvuj/0seLNSd5Hb0yFIY0utvU5+hDqYV3tcUUDndWZ7rwd63rv537Y
HyaeBIG0IKSC6eeiVNyWrw/2leSltNouirPcUgzjDbFFaAKYYzJnGdw7VqImBEmE
if79hu0ja+rxaL4X053ZUyza0a+s0kgXS4KOw3csK4SkBXKAA6a24G3tundt3kdg
/vkzRY3YfSwonF2kixdcAgQi5ebRzkMehxjDEQW7Hd9Qw1xt1dbTa/bmPG09O151
sXsr+ZOIo+0E95yKxrrQX8oRl1M51+yIDe5pcy9h52wM0C8Vg/lh5eLTjf/zm8GQ
Y0zRaZn17P01s6W4PT3rbnfX2A/mdrXxf488B83tAVg3gkD53fhhwrSUjyc5Lw2m
Ntxm9D4aKr4vkJbGurlECbTJQYwqtuV6lY6d2FmPseI3+JFiE3pIXalitSnUs+j7
VyUP9Ew+fpwalB28qC7FZAP8MMt99L8q+2VxLXsdKtPwz3qJKRgeBVNca1n1pGLi
RvWwgfgbLk0KYC61c0N0Bc2QWXSIjkpGlRN9rnqODhj6qUpU4y9bHIBwROMBYFFP
46sAsldtu0mCsT16iHd1j1rqLHDQeGxb2MsyA8yoXBahxScpUD1kFyi6jKpc7uw2
+N3xfuIM62dHqSYoCpG7nvwrHWrkPChB1rT8/yFfRsP3mPEWwYvzZh7+WWKRgm5e
pCXUQy5rnxcOgC6+bT1+aqenOQRvVS56ZOKtuv728c+XtbPS2MbikmbFKDSIUuGl
kOqX5ljBHpMUUEL9UXthCkq0y04ts0IPdPtL+eAKX5widQB6/nE0j2NFH+7zOfKK
UVi+39WzPZ9UCO0jobWnOvZbO9RgnzALSgt97euA3Zh12upz9zkQvqkn+YPvzRfr
dAXs8Ik46/wI+gqweSBVaxyvs4gtwdskjPVhLGX3imE2CDRt7r8H8h+Yb7D+RdKv
tw6YdFaSBk43AFXUIgPSgHzWskiCo61DVV9D8g+SlXZIxI5ZRlmm+MKMVQmAgNJd
BmT1SiwBG62tv9pmfYcnb+kd/quVNoUNpBcuci6Q5oF0eZLfn3sU8enkLIfVx9Ws
gxGafGCt/wys8CbWJuhG3+z/FgVMXPRmYwIpYjoqxnv/CuDoAcplfpHWco0MCSE+
NOxLR5ZQuYO9ZIuOFDlMxRjn8okVDJrT2OV+9MpwcSrok+60Ck4vNSRJ7bJshaNg
syb/Yp159OrAVATHVhRf2wbyJd7nZSyQQoV3L2YjABr7BULaI+jY8xkUSwr+IXcN
cmXnvyYqSfxVHYq/M6nZQvDwVaH/+R5YVLbajK7mpPzqd2nEqlPkGNzMqUQq3ood
Hd26acsv52jBs8+tC+ikSJkpAJ/EI3venY/CpcrWFY3+mnp+aNs/oyVyaRg5+mtt
q87ytA7DkSHVaYHwPpYb7ddgeXvDErAQEBlU+3+yQnBi8f+b4Q4amuAz3q/MJEJ0
asndG0iqUUkuULRvfl0IBdpeDRpSMi4VDNn/3qCnM8deUqHoiLKI8w5NKJDuNW7g
knNE7My+zDl9sI8+Ipb3cpl89gNw5nUqagiETXkx9VRssnCqY1CKs2IgOYiBo0dC
IVbEp8tdxDAU6fKp60H1REK+nSRm54MOXwhXw8rQmjKHoe7AGWKjVB/3KuXsePF5
M2t8YebR1tqLSiNvKeeHdTO25bb4y78A9+UPz+IOgskc02mbnPVFiFW6Y0AA11ID
J6cpNqYQMAxeu6HMdEq8pYWf0rH7yl8ALwtRi5/9RtGkUhuvC3jcRrlnM/PJJSfw
ZIbJ/yqkySjLw73hn8KvZHBQIcM9tLwOHgoCWFNpRn25nyTbGE++xiLfSpbblpSK
J6ng+C/YVivujUPskK6303FYUsA9p0qc33VmriNWQUCVCv9gjBpsn68Yy3Z3Q/xN
6SKowoM6TURy70+LLPjF2jncq/fyP/PZWp3CZ3qCu0dL9E1mtDCGfmE9uay2qXKK
tDPQXVxtnmzncmsfbyBbESEQ8mqfDavPZ26OLhlPu8HpfPT0h2MPAGMq1kcVYo+L
SGbxLyUtk6Q0aRk/SFRMNiQQQkNV8R/HWw6OrKgCnpaQRr6aQLYZH9az2gH+5Wgg
HwZ+vOg0W1Gozwj0R49C+fHu8aNXlIEOD2GUz7ygu4qixO7dmEQNCX5kvWnvFD6i
SpTOhhyf33gpTIzmOwmq4hgUCIYiADedQUF4bMhGoKfw+oVxwGt0Twy6GAm0m8zw
eFN19v2mNMHghK1sRzukmzBNM2hak5YFyz3DgSwGNnL5jfNS8Ic3jtmQZHyMLrSy
1pz5FhztdyDnJYGBU5EI7GVPA9N+p4d6qFLRu9Gj5hrYsFN0M7Cmlu4N6fdIXKaR
Q3r9dxj2YF4GXzLipnwk7HolI8e/vrri/RgFRAUVOTtYp5tkAVsq9K4K8cJHuTRm
ZEyIdwstDZEPC8t0jx+rMy8qM+o96JYEvltsPaWZQ3x/oICgzXghgQRLgh4yj/SM
6BIAMLlrFyd2Ij6Ld2CDeJgXvFW3Fw6vBGDeftImBC9Q0+CSQmRNd/UQ/RBVsHjq
xHhM1AEf7yo1W6HBDOzo7YXITKkStKZ81bHZ/dp63Ho32wMiMwvprpEubY/LZMb4
QZQ2Lh1Zv5tq8pdmRKgWLpR8PXgMSYuCSVVARU7fdOhJPaF1vZtdGyreGchZTuD2
5R+82uCYoAJ3lvS5mE5BwHxuBh9Ovy5HJcUsoYcrZ8iwUKnVg5tmOrO9HS91dhRD
11A4V2jnn7ECO99la4MwWYlTA0ImAeaJoqdsMRnnuGLcc20k6oo9txi7WVrJfrgP
6RGtTMJ9Vn0pFe5Lnf9fSqbOXaGFsELwYUUezI9AR+r431zigB0Uk5IiLyTPcXlX
G1oRWv/GRz+gawdNt7TX14/D6+zqj1sywhuhB9maiNproJVj03hU4kHHHeKLrmW5
DTG8m+YE3Vzp3rK/RAhnxuFTtiW2CYV7dcPpijscBGGprQ6JiXVnmknKW1uPyEB1
4myKzepBOZJxeDCtmER47qC9bCo3NJqbtJ1X/TSNpOvwGu55+z11+5uX0g5oY5vg
5n9Oc8ZIFgEsvSDSWENs1p+Ak4QiGXnmaGloVD+d0yu2rrrk8Z/WuUWAVZr/S7Au
HU81fW7WEFrbb14/+ZdWo8zwDs8BaVhkRbfawesIZ6DkCz4DT+wr8ukXSdu679Km
bvVZVhbChXqIpTv7OWGFemRflYoDP9Hzyto+Lc/tJoD3RgFHb2ymHyOduxd0lR7Q
sGkx9Ma8NgSkA8SOZe0rT3YycemQFbcqYwc41Ym5C5/B/YfyYY+GVnnxlZ+OSryG
wNn2ZhjjzV3VZ3hniqd7S62IcAyUSIPwDT+7JF5tgyidL7Fphbrn601afzL2t7HF
jnXGkUdC0u7HQWK3VVoB6a2raL6tZ+8Kr7oiFw2si1mcxjMAjmn/z+OYIGr0Zlp8
NPCjVSeZsLBuFOXYnlxRk49WGqsG8ItjP4qmIEJdgAXjOdihGAnG+lcQ4RvLp3a1
MvJuXMf51XMMiry0nww6EZvWloaMsg9u/VRFjHWQhUL2xes2E4f6xLJJkSOYZWX6
zwB0frMyVoHb0tgm+DOWKMB5pWklp6sUZqUpw3mHMYAuOvnW9j+D1FFDjZ33wwDG
XHCbcIN9I5CtTSz/iSRYx940hfHtbHxCjFi36hYgeG+llnOnmxN8Ec7fqXM/s+WJ
iSs5OoX1xmJ+MDdLx4nVYYp3+6IhbbaSIB184FopEpGs16mwwo9m9xWtGeqIZoM+
NFA++Vfgmro1x4ESiYSeDwbKSezbZ68Cm17yvcbtrquRsoSEAOrxMXOQNfcSJku4
ZdD30yWqx0Lqkn8xYnslBLClCJplwxfUnajcKlxjrPuSGyEqaR+K2Ww2LOmXR/ED
tX62dOBRIQdWQl7offfQqeRdA5tCyzzyopH2pQ/eeZp0m9ZWQoUsHRRLi6qk5R46
TdU+GuKLFwJ2MVK7UH7ehwoAmEOi9M3qUqrwgv4FQpOt99med5iaiNoWsmOWPrkA
PGxBhhAyeP2/mFPbfI/IR+W3lhgjJLMMIhTmo1VOhRIYjCZu79vcwk2Lr7KTC+G7
aP2rH5oSM+lpbhCPu1tkybyo9BiO0vIQpW5i/ZOCZaV6GCVw52EEMAn939qh9Go6
ZpCKRpKanI4Z3aUwjNaUZyh7tjlw8VgP57HLthpKOmY7tQXOUTI/zrQPCN7edKnw
xwV9JDWJs4WnMpIgFV5TaQGxb+VPkyy/5rlsU206k1Km6JelUegzRj/68XNKHQNX
Ag55uV9wNb/y7e4h81cGju3ycw2So0I8I12IFTcZXklvh1hivrSdyrcI/mpxL0Cg
3s+XH7c1pPV5ET75VRQpfLhLXXDHFp8/hnH9OhdNNgJDZOwiIC7XHqXjGZBJUig7
Q8cu+Q6cWC/tpLCuu6nbkexd2DyKwipjlLdGy7e17bLmURAs71j8e/MOnaYltNO6
MuQBIqK5IqVRIQTLmu2nNADFih5qhQCIVUBG4DTfZ6xz2PJra5u9i8vEiE84ipB/
g+v01Z8BjkfzFOmsIvcEupCq5t/b/f2KYwCj4lQfp/ZWMlZFDRC0DZL5sKp6HCq+
zYs+R1gg/+y58XYgcLNje+ODb7PeKa5OADMAh+r7Jb1oirdeIPFnwlSZl/Emxiew
J1N128K4ajF4iq2hEiniMDa30rBkavtPKslkqL4+8oyOozcbTPaKIC42jKi6BwsZ
Xi1ItoRQ0GGqGUXLW2Rh58sscKssMEyqTC09bf7Q4uzqcWo2S6pO8CuoEqneDPMa
lNCVPwropmlzEwU1V2DUWwg1rD3K69DuFzmDUYM1FrCw9rCBm30u8M1SQ4d0cdvo
8QKT00jgICZmYuLCH0FE9LE1mzSOccUobD4znSaaZLUIlHwAC2bCMLDYpaKiOFDQ
End59ejnhT2UELF+891UJFgAmG15HnPK3L/Jdty7prho4cTCeraBIyLV3KMEzh3/
SC8H8u7OfyQdPzQLgrcDekKZmwiM44JHaDuVrEvqpbWVC5pUrgGJBYRhTMlTBNmI
4dZHPr3+EjMTeKLMjh9k1C3FgQ9UzLDN8Y3DodMe6+XtFHV+3sTfSrhZ+8WWHGxj
pSphvoj9bHAsfDppLZ2vrCXxsGRJUKQYGmqYnM5OMYgmei9qxJWMl8i9pF8WIlmr
LBotyP6KOUe6JJkMSrq5q78AUkdd/AjC/crDFMBTJw4ZtqQFQ1NfJD7fW66mFDIm
FLixlA1uNJ9r1psrUVwc8X5feTHBwZf70wn6aXgvZzOQLnsHvHoyfUlkK6dQzL3O
mw+tjyrDhbQfqHJG4YMsOYRwJjx+pcZZDwrZC1W7BcaLSCfvXNQ5pKSbPRrDR5z4
c8J0TxSemwuQoAwEjykZQvD69Ynnrz4QHsFormPOsFMoLiJZuTvunkFr0hqobx2G
mb4b8mx4ocz/PF/UD9iL5T2erwiwtRq8A6THu0xynQN9iB/0qINGdCO/DeVOD6r3
xBhX3gZVM1OI+RaQn5xxJYQEzN27HhEALvBxjv/bSFJ9gAb0XvJcErKP3rSCuTWS
5lopeDnkhJjIR45u8idMzolqDMUSmHakHQ0leEejkSRhIo3ltSNgoAKt3ccqK3ii
Ku0hPOxYnf3GlMMOjznenpohMAJn2Rn1woKhCTvMQq/0W5kL1aSpw3lBI0+Uy2tX
DtYCR1RnEInW0pmKjOzX77Oy0ngDI6hl3D2YENjvOgG72BTJleJzc2n2LeE3kYmE
v8m6j/vEuoDIbAkt7V5jrglBdOou0tRvM61pJ+VLSBMEXRKsRr6q7cRhR3ijYD5t
hDORud900oi3/0qKp+65GbH3yDt/b81y2wbkT2i+WFd49J+IuzXBdXqvujRZ2ch7
u4GciJhCi31yDN3JqqCKBF8pGeu7JIu7/MuN5cxE/6GLh13XDKnA9tJFiEQngVrb
J/nRuIWZCD5BB8JgzV3nnzY5Wz7VJMVg7HWKfvVRSpiznObmn6DLQlpnIJDWlSHd
MdmiLv5iN5lyGq+f/NlvuNNICQ/Zvz8WhTorArzPtc0/bAADWI90SsmT4u/Fvhi6
DwE3cGXORObBMEeYQ4N+wZsitL7HXfvR01oJW86dri45pnvKKKoJwF388DWd06PI
Nouz0SL0WOCQt+exzo+ofem4noE6AtRZXotuQjzyfaxv3TN1VZvM36C55Ttp1uPS
uP77OpHEWpn/nCHkkXYEMbNMFnZv3VQ4ZO46o+gAzYRFsXxdBaioQ7EimnP6lWJd
8/dX6vPsPGRbrJLMOlRxBv0Pnuv2g5dXLkNRsUoeuRavh5nmu9RkVp/uLjW0c3uS
azVZTUerEl8OrAES6mbj+USu84OXyPmPAZ7CPakX1WKGGTu5i3xJr+OtBj2IjGrX
DPI8gtJbMf/YgwMUTvLv2UHpceUf19tZJDkQVH41OAhkV+1cKlUjNatgLFWjhRlC
ffwB4uGirn2aYIx856dhv02auchZosiKBShYiksoLGgZqBB74VwJeBIOcL/PNVYf
sTz6xb+HNAhI2ta8Lk/OIydR7KAhIJHTq02twaGMk5DtEuwWREui+k6u8tFlt3aj
FQNTv9Kci7P2TPm88n6v9+ZjIG7dzNvuBRiRF0SAeMgA78esxj/2daXcy1FPT1tc
04I9IPR6eD5+EdIyavNeFmbZg5tC1U3E1/l9mPwJP6WnN54CjDaSzGh+qSlAo+KC
xefpO1rcIK3WPqQIst9s43hDXeE31YWcecXVmeRRPMWiAJhHY6L3w4YvBEiLjm0Y
F4L3FQ6VPnLsyMG/IGxnLQJk6noAApRUDtg8ZfYQf6c1tSh2tFjGzseljaOm4W20
TUnJo6I6bghA+IPNug4zXuyxHJI/SBwTK3ywE8Rr0mrzXD9FiPzCZthbpl0rAwa9
m6kH68zwUGE5ixvuTus9vgXmm4LHeU+9g4hOXUis7LAl821zRnB/YauRPvspoEbE
X5b7El59CrSnNSApq7NmFO8Fdp0zB20cyTxp36FcQcwK7PhytIq2PUBjH9dedNCV
pQ7JRjIHMXu2JCdiifERzVBlY/51FkDbPUfcnWIKbOOVgdjCnSmK5QokBO63TkZt
67+Ro77v6kuCA7dMnID+Kf3t82YWeVJnG0Bo7JExVf5OpwdDP/JApWxfEk68e4rN
yJob7lRqLJZdzPiWHZyVESZHmuFm8zPDn/52XlMFJjVXYpG1uu2QekoCmKdXLvs8
E7HCwOv+veViev1U3u3fpxMt1lErO9lVCP0z5Wq/gYiHqg3xScMcv6v/kNRq8NNB
RKy+nH8BT2Q4Nghi0qUh/NfZ9lmujWPORUJXR1OzP5Hg4mSIpSj2l3OzVU2IcAg0
uK9IfC0dwUyi2I4X4CKHXcICSCkGR/rKOKkLeGmWA9nY9liQvSlc4QLSUFTGLFcz
fU41Md/vUwVy/0bv3z5W5l5qsW71sQIUgZMeJWcIqBj4MlV30zC/riIRveKeCGPo
/k5lFp+zS/fFJdL3+AhlLf/1TvKjkhAqlJ12KGo1T0kgl8CuZLH8fMTE6ViTIjw8
UMqmEo1ANYUWb+zMATT1XjkasVYcul7yQxF7GhN2DHZcZjkOpW307gy3kNQ/wZzS
53vWkKwL/jAoaj8JQuw49i+vMoRnbBNjl1Qio4qn2gcDn+X/4TgWlmWeQLAdUVgn
BLhuXz+u4oxRqb8+kkCSWVjyIUNXvtnaxXkxoIAuP71x6xoxKqwV+HITMBJIcEzA
ekirhyRkYf9svyXvuNu9i4izKIJwyZ6JF9leyI3VfTuX9GiEEQK46mr+ayH2mlw/
OyMrgBLqbcOdsnHKIRQQZCdooarbVHklBiBIVShPd/t897H6RSKHAztLQnxKUaA2
jsCeyTrRphfvD7e20kYvCfD38cGY0h7XpSaJDXPibiW5+lRbkWDyUTwnSwFgHIwf
vFgW6F74X42kwN82ajiHujVzuT/DK6pT7gI4b0IIQR25gUUMIVm8EGkVx3aw/p+1
ichBrLISXeYeVMUGzD7L9NlOadkSh6rex02/ZTrIZMyMXWsiPaP06H7HWVPRrCeb
bu+Y76bxVR2JaLRqCEjDY1CANTofP564DajfQ0o9trSR8v4mMlbntWrwG492D2Re
bHWFwC0RkoVRBEUKBxNPL+mNySs+uFfOHcg2nSPEwbIRgcENW4DgbF3Oxxeo+ac6
UHwFj0IR+alWluCQHCwbDNsTEWYwtN+Yk3rh5q8c4NeZrZH4BWhIAXa4h55GIytj
uNdcAgsGg3s9MehyarWJm97e0VLzq2Zqi/5w6pVLfkncTXaCM4/2yABq8KfnXAaf
38JNTCSSqCohrk3KgSNC8Fu4/FxPTEr/JsU+8skTEl7H3f+Ufc303ty0xnfvtiC+
UI7BhUQa4izRgQlR/0LgVYExa7a38+4jV7LjHuu91cdkNtinBDkBIEcEWZGU0vPJ
CNHxJ96OUnMQMK9fBp4r0whnBBlH7+qKjNFhe6VTedYgQ3efcfgO+l45eUE1Vred
MQK0pi+yC1ZR97aVQ1/x2/INMVMMWZk9jXnPbuD9lGUe32zRi/8fFKg9sFOchwfo
ABvsNL4m7KHWBPBYgG2FNcrrHcjWvO9hwBR+Z2ggm/PELkGIYL6rD3dijk3c+644
FYsJlvdCGTN8n8x5vS5j91q2JtOYgoA3DzeJq2AlR6+cItZ5ptcEI1fbtiqZiuzK
Peq5JV9lOy7faLCx3MHm1h0VbcNXIqbLMZN3Nwny3NBN27+w9McY9rswuYN9P5VE
pYFP6Gg6VEGHb47ZGjtNonkCNkb+8Fy3SyE0OW8hyn8NBNKRNCd4wZ1MHL71QUDn
JSMePEUM+yrrHeOkE4mzIDYkknXmeAzqV6CERl2w7u6kuE6OswpP3j5+9moaF57Y
uBMA4fadOMoukdu29SyzKv5lKShLPnWHIMsBPo6hmfzpe5jeNJitNu8fYKdA9zlM
1W0LFLhl34egEKIwhK/50N3bvBHXVrR6wXhJVPJ/MjZZWsuYo7tV4rrhVzUMKKT7
eyVzts6ZfS9qsb0bbnMXSSHgFIs38HIZom2+PUiW0ZBYMhD9DNZIxWnSNsmxxycb
JGG86qOzDk5UURDJc2UPVtuGegGkshL637/uZAKJ3nKNyC1cvUrdTfu+6akozCDn
Fn7KTKal0jEg+8BnSm8vI2waDfl1KZhttQYArMMeQIeH/xNp1a5bYmaRQMeAZ8bZ
zgYIwC4d6FRt2PfY31HqK9jkQcZbYtJ3RbXlLRJwY9G/cT3I/ZjkZct/+RFV/+Er
qR4a/ADaVJcotWzvrnuolWjT0vTCgZA7mF5TbJg/XHXQClTDhbK/YnlUaujUG51P
mZGC1hkN5LI+/9V2u5F2P+fmZjN0JJU+JaXg1ESYxO+fpSR5HleyGFWBk7s6MEo9
eQ2nqhjv1NS6tuAtFQjmiYlbqt4fgChP8lPcBZ+GjZXIN2tG/AvED9F3ao3sf1dV
DMQFkOUPNZRm27uUrE8oJGsdHAiEX38TMN4gO6G4smf0hbp9XU4fd7Qw+g5SCL8N
DWIp8gdKL2kg3t3GswHiM0FABj1FsTrZ6mhym3N+ydig9c61MbUFSKp4vfWY3VMj
BU2gbToBHdLQWZhE0y9RbOtrgabB89OwK6oyJiYMN4hAabuhfCWLtkNFcxGMLZ2F
n+sHK1095+U7jbGgQO0uYEuRYMjRjW0AAtIQFu2ToQ/M8qPjggxQ+Bkfxo7nMs3b
RGAIIc9U1wQuISegvnrMLGPEYdoeomhdRQ2C1XV/U70Ercpfzkb0y4x8vrK58p6f
Sr4ut5CrW8rArImpNZwCo3vOeC7tBRpH8e8JdmomaE/3pELqiLdYYBlZHxBOwiSs
n3NLg0Pimy3pB/CGBLUY0z+NAX77ChwK24CJ8S7UcmpaY6EFC/9wqEiS4zgZBCv2
YW4S+sDsxpJsQkS1eeYPuovoM8rrk6YNyWJYaRyPshsIQyoH+T9gP5dx+8LvYqzz
KUk4AgSUbP4ub/mLmV+py+xtaTSNzLdrf+KbFTXOPaXmXCK11vnRXw+qOtdAP2Ww
Syt2jVze8Pi33yocy+kovYAyNVs7fX2/LWH9tKd2pGOT5SdrF+Yvdf87gFWfdnBB
qnZaJEfKowzWLwpOGi9JoTUM95iU9iQ4Evd8iLef4wVrIhWMuZB+LEwRP5cnepBw
Yn1cw9bYfGmrrcTO3KFa/sdat+f8pWwVAh6RP8zJOJFjNlAWQU4lZpifa1plJ5c9
u80O59Ycrbr9IHwjBaj4o3m5F5OZklI3mFIpd7AEtMgGp+blXkJntadi74d3EVAe
npyLQlEiwKr+mg364GpDJKGICTDlb7P7lWnnO8pSGB3z9gwHTVxrxntSFji5Toi/
xlmjgWMqp3ZclcoFyY1z8jsnXOOW6tD7LVWb1yS6d/IMUXmESW7LOOxhxgt4z8EK
YoVEhVpBP8Ox+fKHTOS9O9DzF6GpMsvDBkiZSt+ghvDwQ9gLZi1H42T4OwsOKFne
2mj0pFVPZ8dher91dk+nn829AYUYsipEMyAaIh/MXa54ClZ17eIJ3tZTo2c2KnQT
nGSBhmkG+kEUrGGLwQGEfiGbBXIaR10H9adKzvu/FpPYawVd4GVFMQkOf12YdZfR
jmzJ53LRA2shaeIf32JhIl/T1SnQboA/gs/Ck15B3LnpBfvrDPuzhkJd7mvNvX8m
VvS/0d7J2cG7mjM+HEgkiJs29EkdG9AK/dOgeKF68Mx4IIU2eP9akIhJljpfJgwq
t6NwKxgQI20Yi/cf3NPYBD1z48oV6rw9p+pdsa0HLJACK5qn+EDx1axIWDrneXO6
TYt/rAZTsg7G/zADWImb/NkK+A8WyCl4+Mkhfz/dJd/VsOLFz0wwUDcb3ZNxVc1U
6NX4gArklryQUFMGKuM3eUfkG+NvzvMKhnXjiGEt/Hmr9GsV+yIi8k6DcvLU0mR9
jbM1ZWbIVWp9gI6txsnvWZHZgOqouCui4OtSo0wVHY+r5y6Uujt9fvNP63I9cBX1
WXLmN2f4GYXFtxH5skbcx7D5fwXeX07u853ZNsU9FDqCLaSDepzyb8swgD1jr5ki
HVWeOFOY8X+cQbu7WsP61RTrhGPHioqyejwCe0LAVVFphPrOFhJ8z6h9QY2mwL4v
Ohv7zFPi0TKbGG3Kg87HYKFktw8062LA6JWGVXJ1Fvnmcj9E5r5QEKIbYb92uTa8
MEl2hQt6uOyH2vI2n7rDaxY60wADRQ+cFrrI2YWP5LRA/k7RwD4k7KKZ5TNZm/jC
jXSbbOB6Tb79cJwUefn0LFmO2dzS8KWAXeT0w2CmDoFNjzUS/kHnXFNusVcbTWJu
01+2YhNVFhqJwc+0DZel1iz0/WvNredOSGUwoAF0RaiksEO3vbnYZVSQ/nEdu8Q5
+tBcoGayI2zlVmWCARDqwesKvI+smXQ8JpEyF5IfKiw8CDUcQ8YZI9KzSVJd8Udf
TromNEKZUJzX8AnBlJWZeHxNasaYOz8gACIBT6Ubl/TId43tMEh29LCL19wtPh3G
FbBjOf3RCoWx8JKQWveUWPjVXcgjnR31NezDQRFpLeGWKEgtTntjbR1fIpIrt4zH
sQtB85MtkA9C8KDGfD9MVW3duvJ8nCFtMxcm8svJ3zdJMpRIxP+9HdWIhT3XsNd1
NOWK5cZlxMTsSLhe1eZ98OQFzxEgFaCy4DMXcVS5eFyeM2MeVvkgIxXkvoMwq3Pc
ctMs2khcUGSrH7y1e1WF3sm57XZON2APgbhgNwIoE9xQVH/5We1YR6xKwj5QBsS/
vptq9+kYId1xjAbRUXlC8QM66Srzy2IjFQeXEUAXOaAjBbNS9Ot3oSD3ypD13rdS
/bQzmA7ecxQPRx9WAFemzkZYdQlJoDIh0nqMspPwaHFE+qSaiZHtjNjm1iNBFkkF
YOr8wnngIOwnNxeOJEvPq+YPpOaMbxkvv0dcDKGWHSRIj+vxpT4Ctj0C+VkZrbZC
QV0IZC3GKqlmuewMe4eqOSfK5kVX1C2yT7ojITSmmi7nh90aYPGmV5KW0+piS1q7
QUNzFcPRGCLOsqbdGhamzoJdyYy9KqdCj6p+MDaz003kI6GfjimpakRLjr3ke/oz
vg9hsOvTguvOS1TeimuKdXWBEYzdtc/ylzkTuYWctDySny1Wn6uguYmXXuLau1oU
uKlO1P85IFxhcijGEiOpKLQGhWfIKkgT3mXcCx/5IzRAXtihpwIPPbqiQxa6tY44
JxQSMVLQHn+POiyc/eeCvNYecin7+akOGuTe02DzTCRTaQkn3w38sPTO/fxqJHvw
dkSfgeg/3gjHfKeBMa4ldC6JYaYRvnf6KHsHXDjgMpyYEGLkxfT3bcFokIFgj4k2
fWv8Bw920pbIz3edPrLi1EMmC5V8KBigiHvM7dhi3lHPr1NjaiaAI35TccYAPSEx
hQuidPb31gFI1kmKtRLzGDxtkAoKAGFLVYDNEb5FhLDTK/mmX7qhpriB6MyZDB+i
Gcd4ZvqAGuIPEVHk/Plo4Mt2O3nEfKNfElFd4ScPt/hna4QgIaq80xJXeY0pcYj7
16Fs9rhhXP7Xr36G5iVNnKr2LKM6CR9HGd8pozDkJUqBCAZd/Kyf6ZleDL2rT8xl
walYW5FVPdojeGmQ4R7aTHDED/un7+6mBIJk4J29HpacLTwc8p4GBQgTMWhtLNqA
1w36axLBVzKYWVQjLJDejarYn6hSsjLgF9FGr5X3OpAaTEN4TJBGZUfqIsukymbo
PfNtGPyupH1IDOWhlf3M9dUuz/iipfN/4ZtvoZGg9PzT4z5F4lqGRznR8GhO3aG9
e3j7TODbBUBZr1Sj6aqvQg1hpNIzanEHXkYdTkZBgeQocW84DEMPRtVcIChhmYW7
v14drawf6Jtw/WsBt+AUd4p6gluPdKfhARCnb4RDes6ykSKdA9hsiAf3HlJ5Dsl5
NPtivCzbety81s/mBPHhQgo5GvtJrR2iDNmcqsBQEvGuu+fynmwVd8cyPz+PBsPg
YRwW3VeEXNhsQtDXa2i7en7ZKTWST7+C1VciTxYPUWl+Z/oLMc+R5DzA2uCrG2bq
keBSYu4nXUuohmU9rEw2orgHpnFQLkJQ7EPTlIEczDxtB1ccX6WYOFWP/5F2sijC
Qtjho4FrmMVkmul+SozO0usanZvDBcXWz6dZgHE6NNU6SPWSTMeR+nHsYJ01zsQA
9EMBlLXWIOnao/oXhnrVRzU/KX74tQWEu257Pu4/+nndCdiBUiGG4plNyPnKg7rQ
447cbQGMhIcKKOGfA/JImNIun6KkP21iG4JQL8OPD6MpBWKbSj1XPI1HJzEOCV0l
hYIJOHEzx+p/728dUJKSt3EtFXCgpdVkiSMYFgw6rZHSzz1qv4tXnBPGI8RqLQIa
Q//f8zqrgdjeiYadhb+Mxv5q+Wc5IQK0Y7d+j/nvhCkoNlET/10M3T4DoK+kbu/l
nxwvof5mKnR5gK/F9oOyqcr5Mq0bTmlpTGaNVQD0KcFyY9rDQwvJqI6kA8iSnImr
Yk9L8O2V4m3sM1nqh7suHljQomo1ljhnc9x4R5RcOyw/RfZT6BHOpY8Sjs4Wv0rf
x2TGpm3TuEY+BJ2eywj8hvB96FQx+/ixtd3y4Y9cG1nT2MYF5wdBVtgXNN45c5+4
U1ncRVdpT//5m4QbzL0fIgoUimgbHy3coZFTcjR7o6c4x7trVv6Td5WSEDa8FO84
Y5ZibtrhLsGtU4fKBwM+UpfQabZMypTq58O/+kJgU2tmz7TvSyPJXqU8P8s/6EnG
3QobxydhgieZ1h7p2xXbkYQSNcrNdzuGv6hcM7fo/lXxMyDULI1yVDyBc5gPc85S
+A9NQMwGMsZj1tCOOzU6YcclXfsetJQ/morlcDTFzdLGoymjLRQ9X44OjVzMhPht
iKOdz5G2fevJnNPTWlZBhOxPLSqX+jsNVLHfVELDn7nzRzm6zlu4V5jm8aiJf/vV
vmixX5Fdp7NRle5i4st5ptwr1SlYVZrcfPIbX54a8zp5zX1nFrcAKcI5pKY1pL0V
Ar2J3E0onobGUyGXfjMz103zOY5U0D32/SfqZEoSkc7e9M7PgPq5Ax7n8ISBxSUM
TAHcmhFwtSN+7z6UwhxyDM1/25eSuWVxCglakwOLl2c4jtE8s9ia8Hsic4qxFp67
NnJ+25F4P/7UVqeAbEg6b7t3BX1PdEN8i0MEHXCNvqYlXueLjkWZWXw9f2lAiF9R
Q8Qgd2292wRZdY7HQ8bUc3/svi/7Sa2LGSrGKCOJbMHrsaKfAfK/+/KUDLXI0wRm
Bo/kVzHFjExm4D46gLh7wEMFaK/ZABBNDkJpGIeHtg0nPPtRLcq8jYw48OR2DK68
adTucRVIEXR4hISfxA97GIVhKIDuhxqflh/38IVPojp/OMp2EkIqF3MUs4Zcg7xZ
+kLHPbeikbG1Z1Rk+DRxDm148xet/TWlON4uyhpNtABYGXkaFmWFJlUbPHM5SpuV
duItBI0Fh2plKmFUYpLmV4HcS2Ta+zT4zW5rE57Tt7AuUAQBniSYk7Rz5LlnUuZ7
5Ls1X/keiy886jbfZ3tJphLeIsR56C8DeE4njsGvMrfZ7y3aKKWP8ctZvMNDnh/0
GKwogOGqfbWEgnfnaNfZ+8j/+E9ICoecZpuT5Nxkwl01Yt0dga3qcgCWDekeJumG
LNxxuypCSGEPO4y6y/3JWrdbdBcZbdsUS3ZkVg3h+huSoREMl1Gxuq364pZLtLA5
JX4vkQpvhbwtwU30kDGd6D9WNuQTOqnbIckHk8RvPKzwSjTdXfD08FBgK22mH0zD
7eOqEMrgBz+FDHTFoR8ggoZK+S8gThxkWyraU+s0FBcKaAITFcWNspheut+YVezF
sToa7TI/LH/C3O0n1XFLL0TFtpqS7XZevQRnbFXfxWO7HYH0pMcPRrl3a9ZLQ1Ne
tScW4S3aGGpg1Lcogje7kZyAW7GcCOpesKWftjT3U9TUPNPoDHkTLi9b+e+RL0fA
VhwRm9+wgNrzMgcaVboND5x/wKL8SvHgCNKL7zRYWASxiuV9aaid+sHmWEtfxPh2
5j/fxn30KIyoffulASxNMtxhObhcZnQKkexvVo9UaG8lucZJgfC7GE0Y+fRzuvXK
WxA3OLBZOIV2saDsS1qlRdg22sa2ksKPCxMk9G9i9jCnaSlO7nhxS2sxyBO8LxB2
FTkuCIYctwv1lMqbtfR0gnzKUhXA+lQavbZGfbm3qs1NBf9MuLP7cXj8c48aA+8p
AL0BBg4SpWnUNiTMiAOrBbMXPfw3ZJSYT4m8KJRs1bCNUK1m4GT0LgX3Vq0UR0kq
lfuB/+CvEj8eNgi1kx64VomocN1c8yEiRPajzyIsKMtK0XmhH6Bq8kcFg7kEWcs1
ZPK+0gMzGCFcnNJQLst2Q11bjitbsmXa7t+evwJ/n5m4sD90mH92IO9DnTDUWL45
ZVHLZSsaM/0qlHyXtboMTon4g210XW1dYzr86939gKMR5cGelXZKJ10Gwc2u+Mym
YKEGvCGZvpINdu7Ka15XHILmvlPuQlEKy4uJ4u4vbQS4cA0gEXd6CvpNwo5PmtjU
ui8lRllqzbK0i/3t/B+mEhHUQ64730rBI5uOeUSS/GX26XzqMvYtIivPQVOfCTkx
4AVLDZwyLPAb+g6HnPEfBYc1XVOgFs3WTthYWuEyLIzEm+MiQDRUhfXubmC1Nfp7
YEuLE3vYhXi86SABO9adAcbGqbrMIozuWcvOSf5zvpuNej44hLKkANrK1kyOHXZD
/C/2ngPjg4DnYd4XqlghXWjpPWzYIyDBWDDzKuOEgVux84ewhgZSgGP0mCqWgy3g
csoQNC5LZuLV9VFP9W1ooRiLDMaACE7DB93inl1jtbx3yw3rZDh/l6tbvWZr8vhf
k778mZTFuGsn8f5IVNVOr8IoG6xwk/Khzr+5lXqdiBKAnapboKnC15dQrZm1tJz0
yAz3OxIN43HHCOVu99bMYZ7ssdzPAhfP9hFiPbEBvCq0iTB4zLfcap9FnNcoADJ6
Bwz496waFqAM0KR0Rw/uJ7KPJLcKYNGAJzLc6tErkQ51TjxYcxgUJm+//e15yX1T
fJghtxHmpsDTUJxHN5TEYjVXnLLZ7JHAhz2nfoHpDpac+JXgHmTdkye+f/JM/bti
4dbI+15gTHA+Nq1/0Tu/Gl/8CyKLYRpShm36IrOmAYkASPR/Y74k532oQZ2WziRV
lBiTDVPsKSXmqnp/9mPt5xRHOyWqR0XTrKWWZeqSYmSTI4X8K/smRi5YVWVfOvT3
ZxzbrYqiAoVsMTiKjNMxprGnafj6r3YgN8Pq+YKyJlJtQmuxp1BhtL1USTk+6SdX
cNTyy62IYYt+goLuY9RUXIBvYxQpv1Q2Ab3tVQ3l57x5h2v8nRQsCQmwz0tiR9b6
1or2hEQ7LIZlljwJ4nSZT4AeKZS5Ow5bekZvbv6L9/hN5dt5t4TuQK79CnzwZ9PV
H/7306GzC60yR3z7DyemPDJL28HyN+NLcyySYe09pFUXs6x2lC/Ly+eZrzDVLy6i
2e2dOo2bfw5OyhljRgTiy4NKScZd0dLQv5OlLDHWu0QDElqCUWqYCdu80T2XfUST
eDbY0DcEnT3B0tQeYTvb1nCEh7nzXFsfTwzI8HAMvD99m0y5kIuw+9VkLPhhWqay
bxnklijOZGau4be0ID5c5rLeAGi+NBRAsAIPlAUM1QXDaDMHDTFz2hIYvg9iqbE6
B/qMPK7wo9Vckm6wrJj0LbbVEEDdWwEo3rV+5GdZp1OqQOWrAlsq1im4oaZhbNPX
Dgp45fbcxR4c92cLRx9rpcROaVqRHAJqJq045d+WRiaPLbMSES2uX7+5GutMj/TP
jggqoQ6eZt+Uma84zER1t8lanTiqNwSTI6yiEl1UlhHe4Z5tbDLf9S3wjUkzAEM2
1aNiFUmWW8V9NCD0sYLcDxTZDee2mYmU9W0rmPnf9mRX0Fq9Xxgb1/QK2UZOBAEg
BqBFNP7s7ivJzvzoCbZnIpzN4+vwQTeJ3CVQCIMKlQxPAEQlHtDPO/RuD0PXcEFb
yXz5/JqetXy77GW5FhwkfviLQ6nO1Hgq6x25vUamQ940lSQJk3KQLSX8YtSsh3Wh
+ZvCKOIN4DVI7x3cgCBAHdNKnMymBD0qdfBjSjkdWEfHF5Y0/rW8ZMEfYW1m7ECf
RT672T21AhDKVyD5qZN6TulYJFsAy2TclZPEJANl33Y7IaLM165wZtZjl4ZbiLki
vt/92SsJWSJ1Hm3EPyG6svX2rQW+NNRjvsVuQCxNXG3LTfmt1diY9/+7p4+4yw5v
fkALCjCQ1Ceii/y4vrLfYR660H7lqRqL6O/2uY3+HayYpz4cRhMbQFMS8FzowmV8
8Bxu5pRnYnw/Jwz4U49QsUf543foxNtVQg/ANCLWXf7AEqM54ogfFLxWPuUQFmc7
DYvnlmmheUJBOCHjXF/u2XXlGP6ZYn6YrEdD3487iGmAML0DB2CiaJ5SLLlnwGPg
GOfSL7Q5BEIg594weFA9BxKJEebtPa4LH/BgHTqA5IAdanWSJOz4idh9GS506U/u
QNRqEus+HrhTalNtVTZ0XFNMXoVt7yJznt54sKpY09a1giv8DVwP82gQDI4FYG76
owELw29fFfDgvaMcX2LYNj3N9T0Fv/TVJEPQRFWhA84SuIo+3Z08yJ7xPvJPlwGf
Rmlfl6XvqSQEJne/I1teK0sSehYjwGsrnw8kw4a1nyLQYR++Ib1+IvfL3WXo/4mF
QbpTt4Nod3QsZGvZnIIyKhgUNKonycEqgET11ivbM8ex507OrX15OTa8WwfwWm/l
bjWmlOQ4qwwQcNBIn6v23j1l05O5NjA0W7hwo7Mfh0GRFx7dnQ2+F6Ln7Z6MD9gB
afoZMEDbOR0IVnHIrPYo52c6wWU8+3DP4/fiFRHloBIVXQwz2d7k771sZRhz4S5b
ygLqUSENsMN/ugRbeSulyP6QQ36e73bq1p+KjeFdZklbWbNk3yYZF3UWejRWtlTG
t8ldPAgc7yDtkdQWeOEBxmUq8iSP3Bw/85qVErTbJxy0jKJPNuF8O1nb+3TBxxPb
Ma8FR1sm9w1SQhERjtSEjC+FyopwmJyCCtAG5xiK7NZI7eYYyTEDCXGReqm5rEQW
XGHk4gv39TEg5s/H8K7AKhoZwOAeALYkgiQYHNyG9vKA49ByBomwbNIf+uNAIcti
V4t+dQ1W1/ZXXZyudAzaf6l+/CLig0dGxa8Ctnkn/kM1vswZ2hPpPEiTg0feclLz
H3YFrZS78RBbsv3vWDZb+YMsYTc1/GpVYc/dkA1epMlJYnogM3P0XgX9+VyQzKmb
5zFIoSk15Xa3+f5wVqadyOTgerV5GEOyco2FMkfUA6CJaPRtBq249TrBo6xoZ0Hy
pSrC/Z/3dxn9s3+PDxGk5Pljz9LF1LtanNTqwfKMAoWMo9hYLbvDrglt98T0IgEe
aPdX4x8G/IDfWW6JuUb79CUThwNVM3Jwvxi5iXZygCCpEui5ophFa2ZBPH8yuyr4
fuUb8ubidUPaKO73BIxxSf0GwCebTut9SUHQY1opkR33tbqNnRE27f6H+ylzcRnz
ASQfYwhP0ZIeKDrL8y1GE7jWJKOCEOLq92hURU8avFNydPT8D/7l6JChVn28n+MB
dQlAvG8c6163eKQrc+eKftkk2spNd1emrh0Qfu0q9elhg6eoVnoz8gK8XQs5xYLJ
aXc0o0NrVXKp5q73MXItp6Z4dS019G9nzGCJuX+wIP7Tm8OkWWdf5pdIpcIsdplm
K7f9KniX23EVmUmSwzF5cSWhDexTMzxfjknTGU2QyG15NyzZBIGhy/oEUCIth+by
x6kji+LD+rL8uG5+WkYku4ducW75BEW1mZHQ8H/gfl9P6dFcpekicm0PJKwVooAb
Ro2oBZ+SV6bigsR9/X39jg+btnAoE/h1NqmnK2p42pFhQTPUVn3VbC5S0IY36Izq
AryVFYTxWaPX5aF2s51AW67+U195T7YxzaioDdM96oz85R5NU1xheI+SJg0aR1Fw
LD1DSOYPDRttRT46bS12BB3psZ9eJWHvIA/acw76Me+fKF45amYNmOxU0Ib2suDt
CRMPXllTaTtpo0uey+a/Ir7QRoU+0g0yIWvLATvjrgXQBY5i+aMx8PoQ60GcBTY5
8mn+c56MUjBhzuIaNYloymfLT6R5vN5d7A3LnwnD6L7zqrmsaC4IfEXgTeRNHis9
S+zNcOgAwLkk1aNvJCyc5XLBq8UKC1dIz/pMyRNfk6QDjtnAmW1Q1EKj3DwoHTMa
RhOw9dusS6FO6tZP95zEZy5JavTjMWWszvYojE3YzxhuTbtm0JFW5j/qgEWtR5tf
ktiV2T4JFy9w2BtPnMgFhdy2XqU9IvhORlp2exwMJ4HDLDAp1g5KTQWxQo3ex9X5
jNLecwMIPpv9dio35uFouVpvbneAgeyytVSxvTgVWhR39F/0T7C+lkLnfYTyM4rJ
f8Jf9B8aXlH90zJh/yLh8Xqy+TQ8OCpAS/QWS2l2AQK/5tyBWOsV4ZLWYA/BTf77
1PFwV9f+KU0lBDNRQ9SufXHiZZx4N+xFso49FgHS0kcDPMWS22Ep3g19uBAD5KoA
l3rQ41SDgR4Z+wD7WrkfB4UrSqgDUPBR6kNkpbR8QoMgNPFvFjY7+jXI+09YSFn9
pR4zxH1qDsfcdEM0Pl9tyzIw+yWiD8nby4g2bt0UAU62uN2rSImGcZRycpjZV4xe
1v9sWu+AvpLdbZ480hzmjutbdJr5Cprgat2jaeBrCfbePIZy7MFsRZHyz8JfMuC2
lX8mGIYd5QGBO0RBxsGELPrgtBd633um1DUEC0wJ+la4hvdpv+RI18F8guKrGR9L
hp/q4KgfYNwdbEGZcronmgteiaQH+nSU6eXx5rnC673VzhjEVM2mx3BzDkuKER98
2n4ZjYPflo5hSsvFUPsftz2h8uXxlWUpPwWrG+cAhJOqsnUEBaDl21s0h2NYhbhb
cCqgBHNKjSLxiCS4+kPYSDtE47pF/IaUtFSG18kMG8zyETH8WxEErgTp75T0WS8y
vHSWCCT4EJXvQ6j0VAIrfcA0UFNG54KuZq1T5iDoEZNxUIXGEgiTxDvjnBrCXgLT
cvGPPdzTLC1KFb6flYm2wt+lIIjOpWIfyA0lnNTYfhcCeFHzoDI66u7TUSXpQfMY
UdJyv4ZMRbWnO58wjd+sdL00eKNpFV7gKAGHvbIzisMotsqfug7NFbgjyHgvY1B2
N+OD1ZHE7bMgAK2UYHhNP/EXUUOyiY8x69cAwtXkhHd1IMZs/7Im7jgAwt58J00b
z0QfZ8fMn8J6a1/Eo0Hp2UBeGr6O+cdGdfyOTr8CSiE0Y2VmJX6H1kFt7hT4Mop2
2MSUNQGNJBWvFpu17NBjjhKVms1bnmX4nVZ3p17fVzo677xSA8QLiFizyJpD90q+
Un2qvgs4EtnmsEI2eZ41nENf8wC7RM+Y2Q28Zsh1mdgSJqIRK6N6+DShTChHYrRO
UnYF4CA3IqcMQd/7VJOIZytuoD/PPGaHheFhjyFDxP3p/7S2WakwLz/7lUkkDUIj
dlkUV0Yn9e6caCsJKHChu2BqNOSM936+anu2hW1fyAXYVYg60EnmI/TagSHNvS5w
VQQ4oMfJiAoHbJoO8Ylm+bGnTUu5A8CY4lEC1UW+FNs8FyYzhzUp2LcwezE0sqm1
+BBD6y8AZGhETJV9e/aTY1vqY4css7Ssl00QcQYCJJVTVQfB4RHNJdt7D5oZVBDj
scFTxjasniVajgIztXyuZUUYcH7DilVRvULb3l5SVb0+Bm+Kiv9tlnffsY76wwqg
dH8z29ujpaFgOkWsMIbFHMCpUaPfKXw0XyMAGS9wXkYfZyQh8UqmpxaddRAaGEOO
0UlDRrjdhly02GZvY7MYtBTCKO+5B2sNiXeQ9WAhyZdLJwPqEytyzdJKbO7yVl+H
pX6GhXDEYpvIZELMsupYqEORs8hAIImsHNKQJVYIVOTvMzBhy1+oMoXmQzmnAMIT
GVjUJT5yCWpvyLenU6XEEsFz1TN8Gpy/ZBsd8ROG5JLufo1U++iG0qlM9BxoE5rx
QqdfojGZZ1gn1XORKVKJ/0vMWFeqiLUp76XtePLleuvT/MXpVk8UhmwhDnd8cgxe
ratcx0RKmulB/mdN9dFLMPl+TMXpLqTTT3C+5t4wtUIZD/yzqu3qAubNYESn4c83
xVP0ceWrldD4eHKSIHVfScuQA9z7110WzM4nPJDo44UFzHVByOpcX5ROic3BvtFB
EYPlnsmANN25tYlIxMEqwaYCEqpjpCpRWd20pz6jhWwjLZAPUYi7y8k6pSLt0vQU
JhuQrxWMkLt0vvGcXXEoSah4dY5wZqTvrYXUzDAv0H4L37p/lPj/7iUL7RKN3f6V
y0RAUlzCDGCPhcyq6wsv7D0t+Ib7OuEv6s1c8uso8M7NWWRBaDn253DDWxPYdu8v
eQiSzdBT3ezHBUpIGhcr4tDIU7f4GLws6XgCutJ7q1J1y3UpVFdn00q3TDgctOBs
pOwacIRxba67KGCv6az0/p1xz7Xcbteys8fpCpOZ1xQXeaKBlpdUI/jD9y/iCuLd
4YHs/DylreKWkd9VK/1FF4lzbMYll4uv/foFCmQLcCFBRvOGhQu7VSBhyvl8nMEf
95/4yiDsFmBl4X3iM3uvm6Q/i+MElV/lRdWRVsdEGWD73wbR503MqBWFP+fMyIU5
ntvXFUlZvwNgg8FN7hcwzTtRJW6IKXNTvrN0zc+dvfPnGb7KUn7ddsNFnb5o0VTk
EDeTrNGrbGCmjJ7Jd181XqyBSqxZ9pio4Q/H9QX4031ymQVs7YJAFFWoAxennenM
egYqpBqURU9gYCNA0hnyXDpEY/i2ridU/pihF6dVO2u1fp+X1GxsFbCUNhLVk9+F
0BjnciZyXhUbUTlD4HpfglIGvRYSpZQ3daLvSP/TUJjGm76BpN7IJO00fljwrObF
hlseg3svg8X2wNasZBVJF2ovWLAKS0m+yMkkSGQwrGtuNvTeFD30RotYR2MbqeCA
5I6g2uKAboE4yh2SqhW7ET3KVhQXe8n/cPUJiM9RjXiXPB6zwA3XxOvfklvRYJlb
PP7Bx3N9oErKFRpmHfPApIqWhpisGLQYC12DZJwiCOTOC2SDxowOZao6vIRx21OI
9dcp2V5Gd8sCRmr5Bj8QkXXo/8UNhX+dcp1TIJM38vTJvyWKRyXHFaOnMCG+FltO
ASWJB0qBpwdKah4v5jro71Q88pDyRvQBPWcdoc3yso1gI4gQRSTDQAyvgUfDZCwG
sADa41LuXDQYv5m15W0N0BTNBxDAjAt+oAW2GagTKhojLJeLWeA2aGj/n2DhF89C
PvlxFwFtUPvNQNaKPs96UuTHbFeiyFNe8Ewy0UhcYMRlnuSx4xGg7fbA2PLHzcvn
K36s7U6KzDa7Ay13bzmZ3hOP/O71zZFR4eV1zKx1gIbrXcOx+nx3HlofH9EgGdLi
YUakmDHs8dNLQ+qULaX4D3FZ8cetyEtUjwaKFm98nW9270IKcrJrdAwSiACVHKMy
0FaT9vbQ/J7q0KKhwuT/wd0OhHTzQaq8ZYpQy1z618jdX3SoRwQtBHGgAXT43jOY
JPuJe51dq6OGgLyXzdNSGacWtD1hJQmyTEPx+L2BqDbyMfNHV7++yBFq8AgOmSYU
4TwihHClXsGA06NoWRR7+9lSYCVFml5u0Y+GDnpACZx38JDyM9pmFORtLXaFvE/K
B84q221jmk5zB4Uvo4wR5S/tAuYva3F8bcKDiGiuXAspQRsmR8OKyRyLmB5FxXyg
fbktwrYKxemfqNlPEkMt+eKVw7PlxlFvzAZghCsfNuKo64GPdHQkMkglTrnONQWW
pADbRzK0n9b/13DOyqxG9WgRrHem1rdmv7EM0RN2781QEWAIq11JR3LgUiJ4nNz9
ANfkRAAVpYQzVe1UMs0rsABpvuifwlcdRLqbrT3k3ht5zlkCjIVZxHI3DlPr90Uo
xq/E8KrP/W6qP9VPAn1Xyd1jgM9BXQC2sWI8UNZ5Zh7zqkQlKJE4WeYprj55QaVZ
gjwaocKAiojBM3UbcSz+Q5ASqsfO3rVj6z+8maZ9JZHhd0Zxx5H5kCD4GHfHogeQ
zevzkHPIx1yNL1ih5Omg6hdbGaKniXD6ZrVui/FrXwfryBIArKJPGRUA2BlwpPr8
6dW2u35FMSp1aQBt6P2UQCGzAEz0AM+FOtVhiTyRQUGotdFaFkxoISrgbXQKuW2w
Cr0WPCrhIbXnjNn+EYcaT64+LWz6r6l6sg0ceJ0XLLeVMvS4fRUcViBrBDhQqg3j
1+oTk6vFP61cz8gmtSNKRuFwFO2yYM9lJSelu244eVbuwu3qC0I4ts4BJZjxPPHu
398BUItn6UMmhCuuKeUBvEHFbJGaodQuRFIt8qWdRI0Z6iaF2N+VTbnU3c9qDkBI
9lwxUEslCCfKuVRmAG2NSJEuPntQGRKKrBOtlMB57YEtqhab221TXv8DZAmobtQx
E9dFHuMKlv0lxPLBa48qY0kcFWxUXHU9CAKAqPZA/v+RvYZ6GIzyTorFIkWxI+En
O+0GIVL0+P7/fkYsUEb5h4onKjPx84IwePxDWVamgRBFRizObmeEhAGcY+KbfKlq
DORiWLT29iZW7dwL91p1/6Lb4OHQoUWgYEAx6LhAD1nhxgJ/8E+1G0+kNB4BkyG6
84OJIRul0CO/Jst0A1IgZJrDt8GebgrmAI3cvr1Qrs0X5TXJ9gVhVr9ts3BFtjwG
aFSyEAxP9ybx2G4hFXNSz4DOZARaVIXxBJlTgi15dTOTvWfe/neHSb21kQ2f1aAE
Lo7iJPShFqioM7gc6XIOfvMAUYAQWpnDbJTqC13U3JI+e/q6sJwxO6IodJaHgAvL
yCN98IBYJf0kLzRCX129Kmx+4pYGnRn2hK7nEC6COwnHWoHpUVZ4GYNV/G5e8FO5
HL0MgHKeIhrSHKYdbU/GjR2eOUWvnqII6wafHerulfQCNvCAZSA1luENgaQZzI1V
fYBj9iVuAnx0Upj5gkaEISGERp/Wxsi88E3bnbgtCC22z/DcXPg+Gm6DRXxOBhXZ
LNntJdIst6WwvoQcARtLATUrnEWa/grV/Ji7i82+MMH9HoGBcsmg9hsPZ1eiJF6J
17hx5jlWcVOOZk4WHsv0xUq0UcHbp+q13f0E7XJNzT+4JQVAsnPTvJUFb5YYIxj5
ZJxmYTPnPn/33q9Iw1kK2t3ojodALOJK6BOjMfvVLj3CqqbJEE8v+D6H7J6Y4Vpo
zVJvm2CUQozrfRSBm08RgpoNMPLI0ah+9iW0UUsHc6+ODgywgMSwSOgSPHckFsHR
x8EEjTn3voY2Ds4cxNIz/IlHNaWj0pIAr5yOqScYgQK/NQj770TrYYt8UIaPwX+Q
nIc3kOz3+v4xF3RjBysmnL3rMjyYvpSIyeKk/vFeAa8BmDG3rmy0Aw+aiDpPn7uh
fAbQ5/icXeUXmprqyu1WIiOvZa0NowernCL1lqEP5M7jaGhFHE2/Y+8dgvmwerhw
qynY2HI6i6HHfOFs7otPDJpzPOVPEMqErvGwnr/hATY86mGKoLpJTahs1/AfZonZ
Kde2LIkDHbo6X/thCXbFKvKFenbo/v0ZeeKTQ617UGxYiori9Kd5vpcjiTnGVQML
kJNax8SmDn5Q3xER02YGJB0gFNVdvJg9e3kpPIGrXxD62znzbSqgT6FgvrB0AUHT
zxEMjnevIGNeDIoaLWV3tR3RH5C8lkTJKM5m0TWD+NY6vWQZpiGAoN6t5hgNv2jk
E9opXKG3NsAWbHuxJ/xRU6azEcoyldsVBUnHwN1ZbCaCnBCglFeDtO08jQDFQDu1
2jDvS+CZDiPvzxEwoBhOSDo2iENeMzDMK9FPjJa1Q1aeb4gO5lA+M1UK0H8w4Hsj
DROv65hIXye4TjjK0TezNFf8o4649aP23Vn+BsoBq4XgnKLC0dFq3o5u4TeOF0J4
cTq/IxRxaZwlTdJOxSnnmJ4rzmLhWK3CG5k06z8TOQ/psZkERJrm4M6JCWPMVsI4
OwnDuwcyvvNo2NkOk7Dmx7jzeFflP1dlHLxzEupG5JTbQLlwOZ0QRoLXJHi5S1ME
yNzgVUtVikAM04yjMwT+8c0saB5725vTFcbvY8i0YBtCsKD9TFfgICgpSAszNbAU
309JiAvDbZ5BaWQvnM5wX5NlgwSf2VViEEXVR21IfXXENTZwyzGaRuNeWJOd9hFo
iohCVUMpVNXF3qVxT28LTM98Ze7Lspgpfde3pMTUq5fPr1wz0glWJWwTbHbEY2+i
PJbjCF+32Semt2gaoOqQyL/IhK1YVpwtP1p5lzHTPZ9uLsd/0vazVY/VR4pp1Jvf
+XS+xC0IalKHYePUg6gnD87ih1b/oqhTvJGn2v0VX4uwKLPNKFE58ixrhdpciMVX
+MLZySHiJKxvnQvN6PRoqk2Ufppy5eZXidYoQMKins9oDcPkLevpKze0NgKypPov
mBylUyKO2Av9vQC+xjCLQjb0RX/0ChjDzraWwiAvx1QS/k3Xvgkp5Fe5A6BTzOuJ
GDMmGZdF/WxJqqQ45wEXNdUODFOupxNq3Qnm4Ih//tuP/WzH7dwyzlorZeFH571I
ZzwFH0xMWs6VcOf+KGTmORPPbTh7WiQ7l8HkxAerZjgaQTS72jdEYFmynWi0krTW
+quJ7jg7L0imBj5ycYAUpjJdp7iV5g8ml6QsjN9ViIl/3ASuR0kdQBbcEK7Wl9Lq
qm7ZxPP3jDCP8GuxQPzEjtA0fwDwSVk1mmbw0Kf7O3C4Fe/9XXwnua9r/Pe9fM2d
2mlWaPfXYhBSB5xaH+iRG86obsLv/BJassidYA9366ysE1huPTzwrc9O9Rq8toOB
+gyUlfsNGfI2uSIQiQeGJ0AFjy/ITPIXg7EbLlWNhiVnaal/FEST3zdB/lkWZb2O
ECgWVpGYfP91AzXnO4szxAnrkpnf3nqp/KmmfejOnEIc7tffL5FPpz0mfeAUtYRl
sxi5DNAGOesY1rvqFxoGWDQS8xyOg8n8fkXAAht9Wp2XtUElUULs1JXDwCVXbk2S
09U+0D8Bnn+eZH3/jFHNi9hFC8ME979fuDwohq+boIpEJV5irYmAD0/fz13XO8qK
pvux4JhIdeNj7HDwSjduSujBJ2SUIdAcRQSXcx4p7IKFmtHr/uLCu5BTh9XVE2um
HM+cw6Xx3RaRH4ztodgLhbo4f3eyFkvIPvDSTizQm1nxIG5OGEMWZfb8tc7ksSZJ
qPBiiy8t5RYLBOpJp3jsXWUT95dFVZ9SSmFDuYJlKIHZsFz1vJV+FqrpB4oBzc09
cPirIBqObz74z+P2OC1OJqNiHEPD+QUnCgEBL/YU1FFBuCaFWEHP7E20Qq6RiLsV
NejXxQjXqqdqxtki/92NvnDExXHHJMPfMNuByqQH2MShNFv5/hUgY/czGwnBZlqm
kgqTI2Klj2ZryTewYistHpHffIqBRbQuJmXjJEro0egn87rfYxBBJYrYonJxuj0s
/I2Xq2CIAHgAeJkBv7Yni6C+jloC1WhclacI9jElSEdIdM9sFg1bE60mlDyrCLdM
WvGBassJKLcXh6NGwoEYzyt2dW1VUJC15OLgMXyJJdQ+iQEitu6EC3FvrdZbXT6Z
61I8P0y5FOTujMvFWiUiqLsQ/0rRjFx1wkefBB3BEqvN+HmjH4/pIzXyAu1vGK9t
67EsdvVFJ5NUzAypE2a+FPT42KJeyhrObjpH0l6L6xgZH5fh44Ns9j6PIbil2A37
YhGnvCMe46sZJt90bS9rGLsMmZh8U81yDZeEryoxyrDqwGtMyMujGoV7PzsQ30l3
nutws3/EhMyWwAD0jB/+7oiB3MbjFozXq7+c/8bmF239rn5s+sHkHmgWQAazYiNB
H2jDaLvZzl+eKrSgt7F4Sn4K4qYVGwjX/7z3nrRvP31cm5Vv+jr7SP6THLGHczcP
jkYchcZOyGw0/9cgBFwt2HR4f3mU5Eu7IOG7gyAkpIsLAqwcvIWW4Sgiu7zg1POX
XiHTgqY503v2w1n6/ZB7JHulCmbgpE3pQWAfQoL9xmH2wMJuguutWgBvgqtFKRaJ
HeTqoHiCIiweQkF+rrJibvFvdgitlmtCrgKio2QdCag5lbTsAbqKxGQ4ofwquiQx
vsncN5rK1d/Pu7d2kABs8QbGRzn53gjVwrZuZUlH86ybXhWlQ+/ednJXdfpLp+SO
/jv2jlZUmBrTy3HxKfHFZCkQzczYWQjzFGxvcRapgBFYhC9nvLBvM/71pGX8eexO
lficCi9wSqrbNZpI1DlXyQn4RI8ubeu40z7Vz5FUhrHP65QPWuL8kNA/XN3+DahJ
bT0H6ON3VDcrxyRkn93i2leicANGxFdK2PtyqpLykRIFj2TCcWFR/JAy/p4Dk7qZ
9UKa0J2M5yrGRPzEfgj6SoUyrgMLXQ/G6wv8bD26h99rorJiBzNOpuL2tv9M9zDS
qvtuLceVOy4ZCXGxdCQ1MzDCegXItbzbfeIniitOWX+vZ+zLV7BljjSKkpODYDIS
B0hjCp0aFayLHxjZ6oG4u1j45FkppC6xMOLXrwW/hbCJTgaTmubpQ7obxxmB3eNh
3BBV4hjAckHPuD1s9qRtez/Ye2XuzZ9dgiq5VhXZ5pIbaFKnDEiTDQTg9FYo/Ela
ry7xhIDxKYHJuIWlmcPCbMoL7DAxR3YpuU0UwYGhpjLgE/SWNw0qBmQLo1ozbPkL
fBo4k1MpSj6wQDK7X/rjMIf9y93DjGa0W1C5N0BFILxK4KaJObbPp/lNsRAZPf7T
D9oAerpZCBndiZjI2hk+b7M2RKfNY28jjXDh6HtG/hdxWtT6JUql81SvpRG7VOyj
DYsj6YmyU4UDIij/2FCvkdD5SZzEm+dvs+/XAi6JwcfZ/eNqUd1V2tBaQTbd4n3A
ERbiUM0RQkZFi0t1OKhssxaGCt/kKfGXxOmA2MvWHWMaOGdoJ8axndo5BtGFL6Zk
qZKbnCQNqK6zh0uVOCfZXQ32B+EVQ1HH/MWJxStkzYcwBymiUYeAcu/MCo2kXfAp
ZIfqiZeWtik9DHpXwvvGu7p8sGbrzaLhwVHSmdGCn7yHD7OS9zlGY+jXDNDOanZr
xI5yhbQk3buuFKn+AIyf646GT9WNpwyYLr0/PcpiWltoVkzQATPys5TNTg4MPEuK
3gj5LBRHukUTEavbtFt1jFlkzamWLjjsDrKkHMPeoKQdU2FSR8vi3HAKQmUSod5l
Ppkmd8xAxdtQNcY1mMdVYtydYSGM2ZV9tDMOIEZaF57KocVPGRpzCgYdovaOkKFs
C9hHagi9uJPPZEGQjzM6spgk3q3jIBfDGIuUOhBY5pDVri3cDjhfOlNS9ikmRCdu
jelF4uhiUcA9wZ2NUt/bGL/gJ0F8K7GjBzpcAbEi5F1K6UZKpqgNC4jP/ki3MaHu
dYFHHmFwC6i+ZDqgQFgW9FmET3spi1smjBbogFjvy8TX62jQ4EU5TMv0/TFnA8Bc
a9402mUMvlqAuJ84mVbNOkGoT6TbJs+NcNH/FWPPl4M+einAp8mqT3Qqt4PvVcFQ
itM3RXi6ZokfzoXOIXA138Swbmfq90Bn6TCXFL5vRjpnvui+ltdbww7Po7Dpcsol
5nvkABDCpfedT37Q6X2tT2OpWz6zRSOeJxHOQiO1Dbm0UmQuJf6LjjoqV9nRLQkV
dyA0vF4Q2i6lZ3jXwQxa1PlVAIsJ+8YjWyfwosOPmqkX+F6JIWfkk8U+xsF4Ud14
6mHm4pwBNcCxljWY0mMONxej/cP7Fl+LlVJjBRZB8XSE0PlBbyt0wH6uVzTVsg+E
zkJQgTjp89mhHLQo4eGdjHYzVNm4yWZw83EQXL2i4YXfLGuh7NwUaGGnBXqOzrC5
OXCvFMVjtH2v4kkuncyIfbB4ZT53Y7Z7PCZ9NWkZhPgIsDlsM5L+TjEOmY1Eg7dI
cWO6Tlll+o8obYAR9Mpq/SKEE1MN4QDZ2FHCHYZNkHAaSo1g5pSe60iXeGtbpBmE
O+fG5IvIMTVashXBy9kYMTMeycVqf0x9O5jpgH+G9m6ACizGFyuwSYcfrQuu4g7K
Npjqg+a/z0rsuITgHDbagy2HDgiBqc3Nb4OumdrBLSFd2v2W08ZRmHWtsNXegHP5
6jTQgHZ/I4FlV+Xm9II6Pi3RZj9Du9d2/5UxLaxx1xuBj5J+2vTbA/IDVuKxVXQ+
v9YuytEAnBxH75Ie0g8gHYRls2BTU7L9dETDBmGskpYpZYowxyTFgyG9U+qww1MX
4we1juIqytfpJxTWMniK+UmbK2cNgvhFXrBQDwIW/o9QyvjW3l+GNgT7r5ohPOlB
jEmniUGW0ZucU77O/gLvOA9qMij3Eu6xHYA4Mx+PXsHhyDn53sRlhXiCy163u+6T
7KwcogmDd7CCwpBistbQpA8oS4eYMrhMYZCvHoqBqqD+eG0GtTaSBg0ssc83rTYH
MEz5W08Z9E4ldBdD/V8U4MJYYQVIZWGWV6DS3WSI1Gr2Pli8sWWUaI7SD7PtKcxJ
Dz658NTpEYt2FzGq4kPPpcKnNr0qZge87a8cgxd5EY1U3W/jTL8FIJAirVjoQ/Th
poKa7ZDgJiK/WjbONt0Ddd7DIlbgXCGfNymTOhS7auJcPOXQHfOEa3ahXuLtmulD
9j7qjANcyqix50HnVH4KzHn3QuqMIg/vDL3AF0pKnJwUbFQ8vPSdCj+rojwMK8He
IjUEFFdO7RV9x1OIHA9RnEnqlsFc5cSRjRs9GyCtwGZPzWkOVbcX6KbCiQQdV77a
bKJ5U/FA34Uv3/ptZkZtqsXTDJ7ubVaLI1vIwnwDlSiKIuYRc6y5isDXnCiXRAXc
D47Vs94vqLpgqw1V20Cugzr9y4Utsc8yY/fpVtvTgvxb1o5otyRQRks1HS1C4nfx
ihJs2oWAY5NfMR5Wo7iSoi5uFvNTY7V1NgFlux5k+r3VmIb/RqqbN774naoyp0kX
Nob3DglpGw6BS6xtM7rZ5dJ5hBNcjHbVLNdrmU6//bVL9sXB6H6d4ZGk5vMd91gp
aei1lLFnAaz74H6e1jV1R0qEkHBlxV5FSibB6ruynROLteIHxTR4Zbahdam0qp7y
SyclEnqHxG9z7PT6syuUtdJfjWefs3TUH1viGwpcl4s5JMLFYYIsQwYI+zciNW3V
ZKlpkUElMHqRLR04BqnEplkmVm99NPtD/2xWl4f4AVtgsRj6OJBp+LUx6BlapFk+
E5s61yY+fw/E8EisqjZTn+xTZ63ckHSw7Y6RirrmZ2LlprWUFmP6bKd0KuE9CVi1
pxlyt/l+r9QX9bWlA3xiA68bmTLqS8pCByD8rzh2iRHR2PquTQwxuFerybcyUyEM
ECc9bAoJw3viJ0iQ/rC6bG4gAEQ/lsn81QFuMSO0dt5F4hUTCOdeT+dmVf+C7xGO
AR5qovqMfmX9imVEEoho8A+3hOuBin4eXGbApxpFDgiSIpZPjSDU5YyvSqK5yXmB
TZiRcVV1iZQfuiQnkiJI99/6Lqh3SRHPkYZMB1TqkHojG/CFGiJ4ySEgGiPYWbSh
6xU68qu4dKW/xBfZR4Kd0xu6xAHjagZcWRSeog/k7ypkV+M/HZwC0u7jm18oDnYN
G7a5MAghOKP9Dj4dcQrp0eoWlqbyZt8oNwHfw4jsYm9PsVLV9me319asvT7z6U7r
jPmu2GiCfg2FxYuI5PtpniInQptVsqNdu9ra0hEa8ON5ds9TkM36pHTXdMVOX+qc
PWV3e2x3Qo3xYZFEFNA9rkDXxm91/6l13Y8Jt26rrRBJWBLrHni2uE/a1vKuGyQH
UxJvt1mnmVd0KQBl3fBxq1rcLB8lqsUPw3oMWKdCCtUsjtQZtyr+G6+dB41j8/8E
XYAKQb00x99TSNdztposFn6ZfAJdzJjIEb95PW6Qyu95faMCT7uvu3N5WaXVcNjt
B1fS1fRwVAxE5baz310pQinJx7MEO0uZuSYefHxKkR9mbC1SeUXOfYkv3Xpud9BM
H4DHBFqOl1Ds7/sLDsXdCx/VWZruWdPaQ5XlmUvWPV1vS9h2bw/YVRrOylVZUflP
JEowvZCM28LEq3KXRt6Fu02lPvYXFIyr0tM56k1WHzHgBua9iWMfogR+SOIHiESG
9h6D1r9LS3CywwIGUjnCJ4IRlN6/zSq5RRt1lihbb0BB7uDljDr/YkCnYeu2tbmK
aym7ZN3VDHkshkF+hr+u9XzKfPWhNtamOPk6rLKLy4WH/XLVQa0Mt7IVxSe2tJoS
4i2MZlTlT61QJEkHwEhvOu/0FyHfknYbuFbwL9Dq1Xe/tUmf86JMDQx5XFQuSU34
JRYgJIcvDqI16Kmr3XUTmlbv+8rBUUF5Qt6UJ/aBRISWVIotKzSfe/7jYWAToMPR
R2EoSWcZddhRYTyFSSjXX/MRYd0Z4WLsyBGsJY6PHYc5HT7kpgCJSyjCCEubJhXp
/65jHPPttZLq0Um+fCkJwkNc+w9RyvXkTUP40cYCJH8CQ5t4mul8nOnRaYQJZrdj
8C6HLeREisKXVdY18KGDoaeK6AMJ7YAOb1oqyEIFskNXXthLO46yPUD4piTnwhGy
LYQQcxrvmLMmMAyvJhZLg+mXGE4YDta4LnHOyTUuM/UcZiLXCyJCpKWmP6LNwgM3
AYB2hOlt+bsyqbzUU5UmVaOWviDDRjLKyxO+aFXROZE3/0KpLY1qgejKMDYCKqpC
f0aB95DY32VEZntaDIUY4jJ8BZsazM6h0scQhqc5bgjwfNCWfAw8GLJTx3ExsOQ5
evxyUtic4vta3pva2F/jUlR4GPwDP+5aRjwjZ2bst7E6sDsbyu/G/1YjvI6NiE4x
TlkgvElsq+mpQAZla1uSkFbk8JpN9Bhg3LO0GQYbyWZy9GzpdApB8dLobsbQAtok
jCcjk6kBiDuUHGBlI1ycOpThEq3l4fpcJqUSti/YltrfJkWcM0oCrQT9/EEbFjhA
F0ZB4BScJhqB/0I20AdDT2HEyanyE4bXnoCQqTpx3JAedmhK1W3fV2sqI/w4Xo55
uFfLXUq3gV6s5UzI0wQWoxihZtW6qBnz2FGycwha+EtDEnDLbsD5GtnfH1129Lzs
0eTvwSVUIt+939QJhLgQJgN4bkTv2fjEGK5DB26hM1IX7TAwk6M2uNCK2xp3pvIQ
wdtDEK5qWGAjTiUDA0S3URkinPZ1bzDH8+o+SdYmcBufgcAn3LceP5A+SlTMsH0W
YFeWdXyHWXVhk5Y8DUCQN1ZxXwLEzy1cP60jZ4sLVe5YzS4iTGGM2GrW6B/PZ/fP
+4OWAlsjk266sA2fRysqM0v4K9rFF8W8fIQGuAo49mzajGvghv/x+smhC5KpJlKk
+KmsGdessAaARGZxsbs85Phk/xDiL9RJccgQiT8QQrfCVbdXA2CHHRG3q9L95ibc
lJuS2lFv1rEWbkc2VOc0i0L/aGeT6fCtcL39t24lCSdQdXhWZVJVtbI2zQYeM71i
/x4t2gb4OJk6SpC2QRV6m4gjM2c7dss6LREZn5CeMS9Sf/XmzBlkQphWBgt07Zu/
2BP2kETaNjR6lnpu4Bxa+hJbjPo2bzxnhnfq/l53bmsIZBO+Y/JkiOM2Xel9B7+O
q0y32Snt/Upd2C3CwDT9nthazfRf3wNoh+rFnxxwLrzHYunLFniisftbNCouBJh7
+Ub5d4bjOBJmJlaqugebr18ks41srVukBVgifCoxdohOxauGCJwI1xJiG8kvMfjo
eJkBe2q8A0srTHOQ8MUW3PPIivovF/D+a8YXsYdBrHOiw/tdy2EbJmhMGBAnhaXr
Rv8qwuDNz/7pnVmPShFb64ck5SCDJAdh+QWMH3gLW6rNET1FBz0GnYG+17BMCyP8
XOnDNez40TvLFn0aPg2BTf1fu+JPvUhmvxkvs/NH7+UxCrWHAg3Rf0iU3CfzYagC
AGHMV8yUB7lz5ORsKfU9HZmKGKn/O9GVUHDMQuVcziSVolZOS/7hY6wvZrP5Nb3G
ukBgd+YYwavAlPXVlAy32VZF9S7yYSbIo/wR/y38I0hs4H7FJoMyHB2XIW9ujOnr
asO+7m4INHpD1ZSROhzQ6dMlJRCZSZvPobKEjrSDbNOCPe4zxmyiOSV7ox2w5bBS
c/YHhiOxcfcMY38DLsf1B3rFnBu3mNq1yTXog1D235pA6psDBMJbUsh7G1KKuVsW
jVlgqjTSjjFDT+ffm5DzVKIMoYT5r1R/sC9ymBVKYfkFbqipZ45CIQdwjlTPvnGx
5YT5QnW9OPdXZS/t4V/7yMVjMTsoKCwO+bvi3QSUguyF9POLpUll7bz4VPA8Y2T5
0fr3uRmxdLgVAk6+FZgHLCe+qCtBChPjZuwK6aGrHPadY14UU34AbjOO9HanFdT9
RtSFoJDcwZsq08pbheJrki0fRq2Fis+sRAKipdgBlCGQ9TRjqmlEGznYXEBpwocz
CxqrlmnrtCY23JFMLkbx2mAK2vHZawJxWRsw7cYugZIpGstUnSGDOGc4Jd/CRPOf
rvyL5nEMfQ7/OgIkBYbM5pQqD+oKo4KA/qBSdL5lX01dLsY42DDKg88JoV+5EU//
9EOmtn0LiVrV8SNm9mYZovZ46tJ4fo6roPYA9/z1Lq2f4fltgOMgIVqYd6E6x3Yp
RK2DUeoknBVMf082NK5yeY5FrlZELU2RYImd1427+Sv9LFOs0/EEUeiurh2U1/N9
LrctJwkBU4zP0XFshFYdlOy02nNm8SON/0cwg6hICaZtPciu+PbonfF0IeBXfKr+
naD/VRhI6rUKKWJOIuTgIHQ/bsg8kYePWMJzerul7mL7QnWZCKgjqzs9lFLXPVf2
nQzACO5g1rQwV5ghBPvo8/bXQcr3EuLJGP3wr3cIlVmcCG+jVh3U1gJD/q5F3Cw4
1ETxD7jm/YqSKVM4SDTe1Pr2rQ3Ie6PgyLgtoLR2PHDJDTcH66t+pXPyKoj0XpmY
HZKYXNNkEkw13c1saNZkqpieRqakibrg3NXztuJYazd7ERKz3DAi9pZdlSYXUvRe
OBWCQC5GtZiXqicBq3Q+q4IaDQvdIAkZOQA8kC7mrKI9oA7gDl59/Q48vMD+8Nou
DcnDvZS2Da0TsJZpbpYxWz1tyEflcGAGEkgI/1G/XsYdlK15gfvLnfZ5o9rshvPo
JRni825LKlKzkQi3WYSwB8Z9/iANBR9CuZuFclWpXsdULjx1J04CjX6COqDoIync
gINuyz4NZ0QGMaUBvtXDZjrgzqLbCKhD/HnehgaynnsG4nozovwMRATt6bTEq27y
njZIaSiDm/u2lITqc0AqIht/kHtUvuUFjfZcsQzUv93UZ3W6iBCjUFyxlNkqAhSd
L3XSVGndt4WPczYNX0IVhUPFr+GjsGCTpnujXDNzn2ZkO/1nOvWLiVCj9GIyUBh9
CXZmLx0iRj/F8/4GVu80nZHh+ph9w8GERdld3xwsQPcnTOwTT4GPZ7PgYx0FfjNl
BGdX3RYGGiYC7QLIZ8FxCgdPajiMYdo2Y1zmm9t21LT3zSMREc/pNpapm1YXNXPy
bGEiGMUNrsgVVyTKGI4+hCY7Qwxknu5QaTOcYPgvc9TGakQ0PIKpXqWT59SJH1nN
3ntXYP2xo+s7/+3NIV91OJMFAX4flSGsZ7+YxBnEe3tlhYL6XV+/cXHHrS49uNyD
GQsJYi/6nnrYH5//9GpSA7FayaR2YmqCbA5TEaFxYivFF08oSZBzehuLy5mCo4o+
ep4wrPsDNNZ3LdiT3O2QbHMtKaIVPTlvIyapbRwE8IAbJgv4QvVU+svVIJvoFvu/
m7xbsUeA4VG6w/RqCvsZ/OPaex6hYfH5P6ONahZsTg+9bYQQfPn/H0Xx9G2/84oN
FJaecq/4pWorjReDU8ZoiHYzummdTJ4pQZ6sOkPoKChfDDP8j8DGczHT5kHPizPt
ObL3FZ8vfycRswVR3M39HqnfXyS03hTbJfTVZGQ3+gNokPNecrgvl8QV0Hfapom6
0k8mHH7TF7MkPJoh0VL9YPeudQlcre7l+biWPcAscNQ4ZoM6jiKO0gsI3V1dGc2U
SjAjf2GAW8ceFca73LkNzUu/sf+undrj5IJt+KmOKXOFXAb2xeMbNtv+hompxxgm
36vXozIJibN0/TLicyy7cAv63weukAh2hc19tVCYxXryfNmFVo/dDtmRvZUHp/Yk
bfHAdTHN5JHmWiCoDuGSFZr2kZHnikrwg/jU903pIgXfFHia1WvXovBWbRXnNFLf
PrilzCOxm1IWmiPoq6C2iy7MrZ1BxBiuOiG0WXhD/Rbo70iuew9DvzrDNP/AXxSR
xcgUmQ9O/Q3K+zQk1IiohjSnoJ0EaEtjyXzgnJWhy4VLJICPsrRWGUDdF3pW7I2I
INcg7JlB/3zfemXPbcVs4dD2MQ+lGng1L6cUy/RfUTixTL9my1d7LEw0R3WzuW0Y
WLcmqc382LSGZ753ztomDK9vabdG2HpQKPmDk1aEbAow00oPHGAcdSBFnUnDEVK5
pljq+RFNQUuqRUhSZjOGXRiNSkbDqIvn2CuUOomJqGgAO8rPjPLJL7qpGcFK2HOu
zUSXrtOjg9iiwajQGw0ZgLPF2fTHPIgZJ/sizOi/leukFyZlNXM8KhEsoTdGBwNG
L7+oujCa8UfTXvyMFgORy8bWtQ5QL7DSn4k8/sIO5hx+khrp/ipZdfp6vBy/E0Bq
9ET6UmT1zXAcctAvgT8jPwTeo8+sIN3qIYQuy6aQDwDD83tdAWILPeyKOa82L6/t
FbxcFCb+VwCDxAyv1STs6SFBiYXiLs8S0Qys900qjhNAaeMfEJslDulqC/wp8WmF
goZo8D2qLOh4M7k2RAIENrhECBCr9/76wq2494yx1hVttUVs4jp0Z9zqDQyocF1p
fpXbmyGny6XJLxmUYwSWZdR+M4Tn7N/9fSBXYk7SLmrDJHMdODDv3pPIrHBBVo40
wGm8O9Ll2ruQcqOK/7IMK12ka/sKr2xs0HcHdqbEMfFZJDGhDlQ6ILb/9zYFnoFJ
WUSZv8F07y2WDsrstGU02rqPl261PtITjkCkKb+FtAWP/hXk5ra9FoDfXRkMowoI
9afXWvavHQ42gmZMMlcI0/xnIE4KJWJg+1kauN6FhEb6RUX0g/HzDenWM9AMQ73E
seoNfnC5QzqgctI9mhOCI8zZ/ZR4LAxOD0GERffCucouizjr0QnMss+Kpp76zxOj
tNETK6hI0eIEPIX5GoEqiu+8jkqEd/3YuqZXFsBatrFBF41Iw7d6lfsuOLxNa4H4
Gb6Jdg6ZbK1pGT22Kp4O4a10fEz0LcQEi8MGzsiSqvJOPFtKorhsmflILsk34FW6
gf4sZrVBIu7hWs2PwoWEtAb1iGRACdef2T2+6PGeXzmKFeyMoFsQpM19v7bv74vB
llt2Zlc2b/3LuboC+XEusigVDa0W5lkGLpjtkofpLC4VBM4vzuSCSLjhbOK0H3jU
NgaNksouFwt/dxgfQ3aV3VyobUQ5XTB81U+eArbnojfkxnP8O8l5l+IummJcb2lu
xChOaMb70qd54PZoXO9aKQqwnTJEuljP+FSV9GGrYBD6hM3mBdjonn7XcohW4KG1
tHQVHDm2P5yvmBTm6X5kQC89x797F9U1sY9WrFYFAI0XZwt9aXXdLYk0N6EQCbNh
SZO2jlLSxAuI5fmHS8uX3pA7morWKia7aAZN3YBj3S7FAlZltRd12EZaWbBYStrU
pX+B2ZXauWs/08xXuArC5jgXMgr016NZ73yJtRy9TCuxHrUjiK1fc3cbHDEEyNMV
/jbtRKnC5H9r/DvfVz7j/lWc1UsZGNTENmCcR5hmfvepVStnXWh6FgKWcMRghMtg
ekHgTtH3+dQztz9jlTCPNpmKxT0KhAWGrdPWGwMhuGJxUzCTSxD69FPSgibQ/Fpz
O5UTH9wCyedhV8XILuka57k0b0kIlMOX7l0zz7wKK0YEeHdej/mA8wAmxR8zA+an
yrh/sfIAnQ9y4NUFmQra0lL732BLq1sjqgotmSoodTX+D5rBjKwJHMGOlS5EUyx/
NFttT+veUewyxBCD+MP8VfJ70H8zBndfpV1iLCvAGSt01oJWw8P6WozBBrgtYStO
hoEpZkAot5Kz6rn9G2sOKrqCewWNatpGdiAwKCZ3vJNPUvPOI2A/GLkSjSuqN9dS
Cb21ZWK5dFdSqme3BfKSXsOlKmwPT6F51H8kP905nmgbL1+mT97OSWCga3SVNp08
UzCfpmY+nbyq1eQUdJb97otugLhEe4bBEjAvrmZWg+X6rn6j8sE3Bapofncj41k5
mW8zpkoODGpWP6ZZ/O4R1Kv04UKNjBAKfXWX3neeo3mdMMXn7z32zY2zjGjFZNCM
oeDNuzG6nvjixi1+eS4zWCRfrW9+pHgaaiw06jONYx+W5oboDRVX05rKJ3f901pT
1xiXyVcJW0PBn5W9yZkc126HUKc40/qEzdH2LymwXN6UMMF7ebh1XClor8t8ameo
0DJ0zRG121Aw3vzqvuzmLempa3b5bBP3XphO5NGfg7Dtx9AIvrGFhDZQEs/dDwEG
9HHyWmYpAvgYh9fV2sYDnZLA89VOvW3MJB/slqc5PnR2UfzGpStNZkxiVHQZyWVV
gCuYzdQFzXAaMic+7mwIqLp9Nomw+n97q8cdERJGC7APCEG7tBVmm2WSRbvsMjDF
U5ZV+RMZ1EqxzJLdGwks1aNpq/dQ+ItjcvdYhKzXv82WjJ29onv7jE7KHnHB5rCD
uu1V2jY3ySQyRoSNOu6sxe8ViiIncHNjJlx+xIHI8EnPzAVaL1A7EESoW44lPMBU
8FvLqyKqkPuNzY0Onk1WnhEpDvnD/GnSvQRCxvbs2cODu12o2IXyazz3C99P6VmC
/X5bogvM6RGckaDEAb30jyc50Berpx5FIx8HBKM8jhsxiFHJF7uV8ZIXmzxe0f9S
S3YvjUOVzRNcVtX5nO60FHF53bEW/P2VfSsjxBccbJPOMjvCzM/dZkr/FHIGHX//
AxAAyU7org+6hmmpOMb57+D3PQBbDHTicb4Dd3049LgpKIjgd/Slelr4Rz2wkFt2
WbW5o7QCFyHE9lcmfG68Ryf9MG9xRGmXW4wUzCKAZFcCObFoW3UZXj6KpIzoOEuw
Knv+9BTcev19QSxP2dUN5WZ0B9K6WXMabxaOe4C620hvFdIbwn9oAistqNY+FydY
0r/uDx/MI0dJEXMvtNlMFTS/AMzNcgVcRtMb1pATffuuQ8ot5hylrL3hAg3FwIMS
/HofWpDyMHb83k7UhV3bhXxwxBmGI1cgK0d54zRztwiqkhYX25hh/fDiq2Pwl2y5
YOVb78iqB2c3chvybEiNXK7IM4noP+clPnozl6g7KH66hGm7FLTsIKhaaIIzUbuE
Jjqpa2ZwJ8l9jm54PBv30l+8iZRh4g08Vm1+zgeF8nOIOAvjvY5p1S5dowDq+CcT
rri77NXuuARbrs9g04cy/sLbpqtsuq0/Go13f7C7cfEQhAmehKIyILeao+HaNBaP
Y7qYKWXYRrSTIydIxAKIRu7ggFY3OSCNAkNQgYZ3QuTTGTOrXQPTofIhzf3VYDvt
8rX9vwhJw4qFwJlss8Xe45J8ZMISI7jrGZaiP9EJ5FBvu4FkHJhrnt/IP9xW+o3b
bRl4td3WIQGdBKML7F7PgHcdJ4vwaC2j32eUX+EUeZl7g+VZ+mBYnYzpToejVJz3
r9jgsOhLl6RxS3pSom5Qk02nOIx8XYl7chkXP/cyPMz+t2xGQlfaaYqV3lvlfydc
r3O4pY0qSYantdlCoMPrMAlZ/qeYQILxGJ6VD31/MvrfQ8/oV/8umUhY/BKoltWq
b1FRrbIW/FtZEwT5Q81vp548BJ1DW6r7nlZsDCioRY3PqJO93YGuQAA2sl6LlPgE
0rHBVtM3+bcZ/rEeCRwUs2vbAaTa5uavM2SJDwpKA8lPVgXOmDSSlzuZAX3uOV9M
iDDYtNL/jdjPvUK+VSlS77iVpulHXMSB0zhK0vj72wTZOEMKuytguNK0XXndoCvv
LoLib5qzzZGG8tKbPWHPdrCuAZ5A8bGfiQQMsrFnWI19TV+sVPlbszGqK/CRHYvo
7+42YMwRsTAL9C9i5Txdg0MziWd8fxlKNkc4SduHznrPjLDm4tYoXoDJ0ev+sM6u
fHElN88sY3jrC7Y4S6JX/9p0NiaT0tzq1DX1RBqBWu7MxWV6ghcwYn5qS8EbBJ7U
8OMFqzo8oq6/xURTnE1BCQO2ognJVkW8QLy2/moHR+I9BGCVH1tUPjfUETMDOu+z
AfiR2srAjr9UYb233B6gv8u4+efxYhAvtLIbcp0sKxt/kbcD+t/hzV2wenUkjnQU
N1uhHDT28KKMD8eOo5uVibKCMkAsS8vmQ2uKIiDVW8ZiOzUQLXBskFKH+IB9Oe4I
uWVufbPoQi93WqOi+3EjlCkEINfCrH6ie95SGkEfXoxIiQt/zZktHEm12VEcHeoq
MFPU7RtsZf3Tvvu+S2VVW72cDiKRTrYAu78QRhrmSwaMBen3b4eJwxuN6hB4EOsR
Hg4ab7Lcj8GzERA8wHHDlLoTPX/J6pXvhCXZ+tDXhh+a2I2TUYKRYKFZUAKCLGRv
36QBLi3kvqEGJUGtRRio4VE2mgin15ANjTVrn/r3Bv+npmDiGq1joT7bkJUsNqqa
/2dTfEkVsY1nl05OYEbAc5FprYlMkaOEuy41XYkslEzhWPeonvAIk6877ow6XwOE
STarsSPKQnml740MjeUF/w==
`pragma protect end_protected
