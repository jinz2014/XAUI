// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:32 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ajka/2XROSFeUxMpmXlZzBKhDRn8IrQM+rt08Fy772ZuM9Cfd+txF3q799dGDZJM
BbwSglqq81Ed8ofEqn+qzoT8TdAtAuvba0yuvX4MG3fMVBp6CO/JrAdDjRNahFrT
yzVwIIj+zYwCQ5rUvneW6ha8fK/7tgbTLQkcVoT2Fug=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2448)
mS8Lts1FnBImnT9Qy7CHXkFWOQ9o2bFtdvBUtb0rQQUprLDqQssp5BYvW9RN2n/W
PTjVWkljDjaWe6UoGOo4VKi0dedEFhdi3QmgLxRtGEB4Xkx2zogZ1VRmxVeB/uav
MVLGslx+/6CjmhmuYgaDpJr20IW4J9hEPFM0IMv/Ka0b9bjYd8OLfqzRL12Fom+H
4m+xfcsvyPt075xG7S63eXeckdg8/B4p4G9u4c1Vu1qpj0ny6KoFPlUVd1Q13By8
EA3f4Y9ciX43PI3BbaFueg8biOmQ891DIXlidqOGvX4g8OtkSxja5ZE9ASi+AuOg
Stuz80jXqBkQMVQd2YTX6DIYEteiQPy68A+FbiBq6/gyYvyf7eCNZUyrz/o6UsIt
bep76R5tvqMBZR9vw9uW53F+zkDaP+xMfaaKGqkiFNp9UBh4SeXeIDFApilttZgT
ufZXWVg1mE5FBow0PcvK4XIPbPIuUmpag2jdPht2rzJCOM4dyT4MkzmPeK6LEUNm
IkBA7mBkeGnBrvbINCeF3AxYPV/SIaFVr9tgvb10ENMnu2Y7+axaxd+RZhVBfB6D
shuvMaBS8fytwb6mjp1fKOvIBpqBJ8xgppe5vYvQLbD7mYKmgvAXWNfrLhna9c/t
v/NWXWSBiHSN21qAwLomNjAam7zL4Ggt7d0bVtbQmFikvziJMDniI1jNuBZmxWTc
mCeq1sEAtt4FSPXKdOYqSkGcua0r8YruHO7fWcS8NJTL64X+83tRP7laA2irvIAK
07xIZNO/qbv3rUq2z87B5w+hrMdo+8U4U9ShiOnAMHQtwxjETWaMaaB9KX6836Js
hxK5rHda0HK+xGfTQhS+WLpaBpYOxNh9+VR1bnLNuoA2ZSdb40lBz7AQNSW2bL+S
N6smrfXvoOtg38nhQuPk6s9dJfgtgIr2yTTmFAsn1yFdKZWDUTCbL6HDtoirz4VD
lGQQtOJ+kUPJ+XDBjpr0WZ48/huWcgkTUe/xdy5bht9gbTP3VYtZspfZ8KEMi3w/
IVQwLXeWgmQIRwrU5J79MoVwdQMsM6ZI+bjR6gYEpLIX/T6NdMhIcZsxjCBgpD2R
6P0Cs2sPx6Itxd51BSRRuj6xT4ltQ5UXY+RSla0CrPoQsHVp7AEJBM9Y5NsuZFUw
bJfTcI4zYYes/ncxAuVy1/ITnS0LtWUfRi6PS6fPvfmdXebMPoE7RSWyfIGfoPTV
TD4Ied7GRPsmwB1mSFBsrf0PmbKqWNkLNtZ652XNFa71vUutetPOU7X4rwpUC9jj
V9cFYX/bLiK6X5BRvUuToc4lNuhLvjZ7v5wmzPoPKRhAE1Msw8AI0Jn/yKuYTbfe
GXnTZ+gDRWfVNHYx2qQm4xt56o+BEZe//J3BA5wr+tIleQPkVPax6H43hh+cv6Ep
b/ZkKqrj8m0hu6jiyAQpq1/wrNa+48FUdObxRvkZPI9VpkJMM9OvCsfWPBMjn9zS
Q4aLzJPkN4VDIypgztSH24ZTlAhVdjMc4lYSDX1ebDOgPe2xylooS/452DDqWaen
rhQhVOVvkMabGGVfS4CDLwjWojt8cJH/GaVlXgZ4q9rjub6B9o6TQmU2RK23VAXY
SHkWB6qDzOaUuM5HRRrmtZnl/A/NPr9bSlBBPUYLYk9S0Z5H/zH3RKxQE0GfJMkD
EndkGaa2Qk6HtbJPX+lt+5nfhTVOaGqUmjlja/GZCG6a2jsDdt4ya/dnVtL92SG3
vMvHmCOmm8TNruA8PMpwwBEbjg7pbpNl+pwZ7V4I3ODu8Da0Unu2ifX0pLJT3Vv5
JQeBrLEdt2SJHZw7r9cDxt+06CuW9F4czPTCFCoBneYg6SJFBuX8M6X+zIHHrK/M
cawovUJ7PVUyi+vxoxa+6h2RKhcvauVmqis968X4XFzljoXwgvDJ9iliWTtN5bm8
TI8i3nMdW8z48CcrsZutmgRAETuZiMV3QZh5K9anHkCBepricpmCl0geaw17toUl
RrdniL72auVwceF1HYyrMVB75oRrL+KxE+OMqp5C5l0CvA+E8U1dQ410yCHSnBdP
Pr4G76IK46onPNLv5S4Qyxdk0t6NWwHdXRrI8GKSkvcm42MRf+9o+gsO/Ztp7J9O
nbwMfQ45l19sW1z3To/n4qfVFxsDEzZ8JeA6R4/PYTKp5ymQiMjbFF46ie+o/CsQ
V8a3gCA7H5LmLywhLVhRw8H8eVmHJqnPK8zDTeDqpWemXVGEjaaU0VmW///7xQsz
ld7575jvvmfHKHcXg7Mv8xTmHPgXOMGVnHONm7kwBxodNUah1mNv0McRMx04GUpT
MJUfnnV19rq1eJcGQjf+W8D1c7gb8wSW5VBb2t3sLEeBeB0w1/cVih++fFUVvCFJ
04Rrz5uJ2b+h/bC8LjbGDcFFt05Mz/6KE/NOIBXe7VJIznKLY441hDpXcHruP3gU
bNE1NpnoGKR60dEofkewEXSNvikDZ0DLcuJcUz0bnt1+hutwND/dE/WZDcln3rVg
crizkhN/lPo7hcZrUJ7IAyRZiY4E9wZh8hYcsYYvad4BZ8I12btdzF0+VkH2xfnD
i7trK5t3CLPnlzXslj0mnB7xoKkCEhco/4yBayAleOeSTEwQBKUjY/fcWSaI0JDY
NAofQtiyx37evsjz4gpRIdl6lsMXyaOpFdC7IBaykDzUiXUKS9626CfWpYCTUABW
6X0bDaW2J7JxrzEg3visBeEOdFfFpRqz99sKoQF8zKkXGmd61vitqQdGZNo51fyA
DeewK9q+VEbXva7QaeV7fHwKEd38y3mote4gCsiS6uXQXsI7byl/x9Ji0VpVpttB
vA0kXrKh6qnj77I+jflgIjz88pSYek8SUqNaBD9mOkoXC6+q7tANTCUdoIWrlxrF
sP650XpFzeSGYaotnSVJ6NnSiwZujDOkdXqTStNtjXCqOtMvRyMbcveWMcakbONe
ha/qymCSVDaTWb7F4DCoOCeFrxhEa6VaQb4cKw1y0FQulfkulOzXB/3Bz4KwCFQp
3IM4lyFjol2j5rMkVzP1r3vFWktY4IVxOXDObdyFlCakELNohJ5pcVAeCauP7xqD
NSZ24QnCFFkF90v5COsvAjA3zDi7xeMyF46/Fxguzq5Gj5hIApwLdARLQW+HcZPn
oE/Qr2N9/HiXIEafi2zOvic0eMv3bLAhUCvy6cqivHqXt5g7kUl2iLtEXmJOxkh4
BdTaTeBPl9eKXBdC92d9nUm8kDfw5+sRt1to34UMuf/1BeH3pD97YvS+VsjhDQJo
`pragma protect end_protected
