// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C15DuamX82iNkshQvQPXnH4T7ON2W6eugywl2mwSIiGlDX05C5INGOYtpuKrYqFa
JZzHQLPZvGWm8UYzADp0lXs4jcMw5VjvH37kvMpa5Jg4jodh6c+c2nZLEIg3j8Um
qMAoFd90yiMz4do+wIdBGG5lXopRZ5m+mnj5DPZcza8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11184)
o5pn/je3bB6G8+MfhChVKZ+uKInQ8Wz0w23F8ar4oO/kosEZ70486edhwA3l/4PC
BAXnuzHgJOw6wBjRg00mBhmMbZaz5+C6aGFctH+8L1JjfPY0MHe5m7rExPZXvMjD
c2H7uvos52N1doSIz18nGDxICdSycFAYudxvu+n7vv9a9ukE+Ppv6PjlruZjPfMK
QTZte+WCS+uvXukgvKB8RS/u7L4Yu5KZ1A/Nn6lXsu3Us71ikAFRwKLKPLa/oK73
Hk277gLcJS10nUltmqcObWz87SyedsP1e55x99gbcaqms1+asoiTZPD6hzqhzkbp
yx2Bad3DwLJhroHceRiQmheRb+d5s1XDSvxy9Xq4zf18Cbiw2XOWx1hqmlD2FFQ+
sAjYOkiYZQHCKGDk7KXvBlXqJBIs2gs6iWMJfsTeah+s7o0vovFkjItUW7wXWPyh
wfCXmSK5q+crExE3keUPPn0gNz3YwsLvJdONXG7AH5prI0NaWuoWczd/xLanzABs
l+HpCEU/G3iIcVd7j6S/6nTo1snLkKLhLCxFWReUPe9VqDFRJHi4BadWrECB6r+a
PmMqwIVN6pDAx1FDuW2jevrvTRmaUdBDHZgOpFHNYjesd1iq7yC82PQE9b+1LvFN
FZVd2GN+QSWSEuFx/mIkDambZdmeV++SYV6Su6qwq+nffQfHXtvKItvzd/+7Es7V
rq3AypU/RMEXEr1HZTBe/K5tbn84D1x52t16+bulUO5HylJG40wvhRdW1xbozfcF
nZkoyx7p9Es2XkC9cfxfpllSF1rJT9CELuNL6rBBhGdToQcugE75A8zKjEgoykB1
gwLtXUGJmFN6jr0jR9LNZgIvDSvbgtkwNmZhmkhudS/inCg+zu12sU69qeqqoKmg
OhaQMjKjGYWUQjw580HB7wOZaUwj8UJ/S1YG6HIeyzci2CEWqG34DDWjObMK5P0h
jc0bRMfppOwksoaxcLzTLaBWeg+NCWcp6XdU+RAwxnsUgCbbg8vd7yE2/sfi3Tno
H0OJELb26D8Bx35Ac8cnAhnWVshJ6+LGLamsUV/tVYOR3vmjWwQcD3IH9iq+3uEz
QH/UMv/oLhYMLI0ZNgVDmQW4RxdQoDW69QmVup+5xBBlh3xZP5IFJHe/YFINfMxD
cC9HJ1YzLJQJ1NzY+GhlERG7xfeRRKuhAI7jhO+0uYydPcSZp+e/1uSytP3Kz03y
i3m0NXpo4KCrsfH9NacKzd+2zqFpz4qNg3dW2LK6kywiXeBmyP/4wnlLLLc+BRNu
YQmGm3dfMX4+xiGBI/QnzpU5x/zfQIY9faDA/83v2g6iiuNXZlmoCNlHgh/QvWQX
/V1SbnyodwYODuoli+uVcJm7ukpaQFASriYkuITn8xBdbw01ZtB9q5nnfdLp8ebU
MblgjjWW8uXdrDHujADtmVy5TxFHK9s/6FABHA2Swv9WZuoEk1R5/punDCGbX08Y
w42H14fhIeqVkOxZjEuX2EhlXGj5jwybFIV+XbHVDZlKQWRBy+WSibp4dMKWGRGE
hzjjJWnTWzfkyD64Hv8PIrC6jcW3npGeAouOOT/Ojw+c55WdGx9Kgd/UFv7gR49x
bMZMbV9vFPnyBfxFOlpgTE8oJmf3YhGF53964ik1MbEmCArOQpwJBBZXjJMDi1lh
LJzag0XwT5ZW1e+NU5pqGedXWJean83AiRkrS3dJLjY/W1cJghyB9h4gJLLfNQ9+
1/uJD5RvcWZ36SRTP+pwgKJUc/26CPmcRQEhyPSKucbCYm267b/PqpB063oVtS3T
iME24yURpRiTA21EQ+c+b8Wx3nnLy1iEuXiktuIPS/EmC4M7MPJWXadxlE7WQ9Q/
eLl7u/b6vA2dLZGKFB6dSwX2iQlcuSjPNA5Fi+6OYe+8k4drSuQ7AHEyzLARe/Hy
KmjlrFrKPqy4psF21ulWz1ly9PF+OhrQVoz4FS4Vv88SrBW0hVS+J6cV+n1B5/OA
qdfQmVX3/stgkdZiAfOdJIR10CdviEi/LfKOaixqwe+fRZ0GXqY/7TDosdLxOV7O
JqKJEnFuaF05ED4+b+2sE0cpD0w5enj2KAqLknparxRIflou8IiJ/LvXtGsAfKCy
CRHEz6EYOfoRs25r5zDGj015VpV7Mx40pEoKEEw5+phC2DwcifYTT4RIoFduO+q4
+jI+9fWBXzt2NgAAcWYpoQeccIHTw7nxcko8E7zFKZna0QH4AyVKRJfhUd6heUdH
yk3ZnjIF0UBhIqTYmbuNeNwZfK/S97hTMY82C/SyhSRiWRUU11yD8oL6+kr1dOAE
sgu5BnVFusul2goKAuFXi7SpT/a930QSlHlsR8KSpzoEu3ZSDXhcEuLF+uZkjpU0
/1Dh01nyzb3VqcZy0GrUHzyu9vhtumiaCZ3iGgphoDRWvmRg0piCpOmKRohBI++9
7psV2Ides4k4pUsORKypzd9FnkEZFqtJ7HevtydR+nio1ZX4G4EQ+eW1HLknZjgW
potlYdbWm9Y1PFlVveUP6+Il0nyXEj/NYHpkbHAWYTeSyzd1guCoimgPYVpYpc3R
tKHcsW8lbrfGiM9QdhTga392r1R9TFaPhiAItdCtauFC79zmb64HfT8e/qvLa7z3
HvR9A0rpDZBgvbxWBhFY1XZ15MHr0qMdnvGKaupe/8LBmq2fZyUJVkOqPevzsqGt
+ZVsEJF148hrV3KaDmsSnQP13pMcaIO/nm3H4xkt0yFY/zztwxRF83isyOrbyYN8
uCN05bHiNaynhMliveqR5ivTi6XZEl6tB+btxpW0I6AFfJSGQzW3l3830qDqAuSk
T3F1aOgPdTeFJtqAlMfs/VdEU0ORF6jZ7ZeXeBP/F3/Iml/sEMR2iE/0k1Yt2fj9
RYZw/IzgUZNZHwMrhVzRoPXFIePmn5dSKY8jM9cBX7VSBcbPJ1xOoGQtWtlE8vSv
htBN/KRjA98vc+9pkOpeO1gevWrJqGGeb0mdMt/02N1/CRMlrnSio4kV8cSXPuEO
+cWc42NkRN4WV7CfhdHysTjsSPdq6DbTN0U6ABZkewfNG4wBQyXqM1tGRKnaDEVA
IrZvQdRBRcRdMwnaPwvisBIvDB72CqyKNgnZJKKFgFhbUmFbuy+OrlPtG0QO7sNE
/duDDM5PFobdYkwVlo/icxmJSHIt8SiS6GL3li1xZ2mMtKSQPa73eT/Peg20gNIo
+UosRXf3v8A3Gat8UKSoNe7uDTDQqf992/9XkPzT719cmuTbNewF3NUgsZRLLcDF
6x2bmC4ek7j2FLVbrpkS0AEZ6jVcMuBfEVp71m6pL8KmSCqMsb5COQhYvHRON3dm
SYWlpBitm1ISYH0xEuseI9TyHZfloj2CypVlYvy5+z6+6NMF83szkiGODaOvMOkI
YSMkuXLVmKD7HEpk3TDEvPfljJz4cNCxuasv0C/0VIpTtuyVE4iGUcHEitT2YCTz
C9VpI1lSZnX1WcUP2xMgWNtRPePDtqhkP6USebSuEH3baBuNxChQ6aMNy+AepIx+
ny7kILFtSecBVfuojNbAywjaGjTrKILMhlp/9OwVxX9AaN14BO4w44OgAuri/xyK
P05aFTk14r0YBw8I+aEtVMjXRQxN/WSfyRy3Uel+LCFlWVl0vZV4mfatUU4VUGAA
I2jBmlcSTdvvkUtekk9ZbPlh/kOTxmH0KlhNl1giLwCDOOQLFHAsOW0ZGaLqO6MA
3NnrwyRV313X4fPfN6J72Z+12k0GeWXpX5PMjyGUPkAxo8bPPh3ZYc305gc7peqS
ORxQSFB1IGyV/oj6JO1+tnfh3jYUAdIZo6ZDV5L4fnZ098v89rHQxYFVbELVnZ35
nqzRkM3/WZPUmhmhFkIyv1YojV7X/r5q/wQNV1xPp6Ra7Bou9ddosT67TdNlvIbN
Kp4y+IOGMn9o1IbNboFNahmutjNbWStYhaehggX8vKZBAY7UW7PlFzFPPdzSgV4N
ycMQjO/vns9PCxEC6E7S2gX42bsuYL0zXzs+dFL8Sl3133hdU1lazOU7TBnZDSCh
V/Be2dUjJaeuhR1jOh8nbKGZb/xu8NARJ+aL2Xl1TVtUCTjNj5UAvWJNKZDeEqn+
PkML8eBwV25+qhsG4g1/8SV6Ud96KQhNsu44XbcFkx3N8+NbfNf3TjCNsaqpblRJ
z+4/MtxB2j2ifmi6cuiM9zRhKTNep7jTkaME01RGr24L9+8EAfRpaN1EjT68oBLF
tWISfLhh1id6Zakp1FrRodhObKWc+I61eIiVR1GVQsWc24idDj+TdkF33XzLI4ta
ubeGH3nVbXe3FEQtPC07dLPUTxhWuuQKcGfBQl/L0UCDQjWIxB8aHeZkwRlHMudF
Y6z0xLSkNXT6q1Pq6K4zYRwCnD1d8SS9xLxHdvO8c9gdR1D0tOLAS2Gd2kwFSmPh
jWbA2WlRDYaC0qU7TCMaPEG3yYjdu8gCxAZe3ApjK/LsWLKNPUqXn6BiZI76bGcn
Ny0RmeXIM6dyzhXnrLZUCJ3R0yDmXupSFEBIxwKG+m9uZfWq8gL14SkB7NQBMRY8
cjRtmRqL9KzWMfTaQp9sVVqE9GF+QE3/6cPZY9gmRAx0b118ndPxd5J4vHacebS7
2l7iB2OANDy8jzQczPfouPkou9l6xHZiqmWgjsn/wOYYpHXFHjNQReZyjGz0HvAB
2O8rTFkvy15HspsZTp8imDbPa7SbqzDTut3C4ZFFZCWBA8Fx+qSYLzdcW3evZulA
a/MJNJdGI/Gzoq9y1Uvw0udHvc+V6sJAgkzEKrxryA3M+yBFeZsY+Tchx6XhcZpo
ti2pnCF5EYdw9kLSVpADRmwlct7VXI1ZlFhWo7H0kwQpeKgGKbn9NaR7OQQXLbn1
4UpaJ7cutonrou9vHdmwqs+I/q0uNimflnkXoqr1Cs+IriO0viavkfUsy6C2IHkf
xd9WB0Fd44nX2BXshZPqQAhjOBZx4TXU+weOoR02P1s/+V6kcSPHG9YZ+W+8zcEl
XMySS9jBxd0inBf+aRREy6nRinDBRe9Q2eLFRjJ1OQCm0MOlWP7HSv87J3QA7hs8
nUXb3zvu5+TTF7f02+cCeVmr/LJloufqv8fULehKAh1tOYPH6C0azRtDV8IQXzk5
g7i1jVA3ar+f9s8Z0++VyRWqjpWxq8E/d4KxwajHrYWTC9lmbv3+8/i9oh/IT+Zu
93uq4IkTSDD1Afot3e3e/O6ynLmBx9D9QAciKIAOAOSK3xQB6um2Lge5DJcqy7uW
hTfJjT4lGN/EYHbehkptSQiQPTu+abfgl80tDrUegCoeAU4vFA3sAYjByCU7KuAv
5zGz975ikEXTsFI6VoTnS3zxQ3qxF1kBJlcv3VKcqMdhtqhw3DebYa4Jtw/AWi6c
ubqKYNCOdGpiBbPhQxBQmph42AM8JP6HuvAMvIlrzeO7uGJDdbu7goPMr2pSbLtJ
Eiy0ktDvQhqmKiDj9RcA46Syvr93/RPEXctEouLUU/xUGof6/AkdiqGFeMYfzxxC
bnniHQ8mmaA+QaUltSALpYLH0w5m30EAdwm7AiSBLvKVLtm8k0flhug8NYiXklhf
5TwPcunqzm2boVi/7XKhlcyL6WqSkNeXxJ5ZK5LJoqk9OG6CwocoyX1e4pnCRkO8
2c9to+PiuzHrOijwIroSVqal8jebrJTAFWCGNBEyCrs/dLVEe2OX1OL1vlmTATdV
co17tCTbxR7ndTRDHMPXMnMU6TFuSeGIBbImJ9lxSIV/EYeoVNpVwWvER84nD20t
uD3+48HqhC1YVVNoC+5jNfgAnj7aNIAzW4ZmJtp0ROqNhz/VemaVDU7a2TWozuob
ZblqqXy6l9GkbEX6ZM2kGlwV/87HymZUBGKqkADdctvkOlijUJmL03oWLzEPZCfj
oV7nvAas7D01B0/ipQ8XGJSrL/RNi0e8FBKogVo8LVaRhbxmlw39YsBHSn+roStj
rDpMlugu5CqA4cCmU6kn7EltMKTON15zYuQDzzaLMxWJwaOQ84Ks3KrHCz4YMrtb
F3/nQEURK50Rk/ErbCCjRE79I90iS3uYnDr8w1hhxKKWwn7NO0wXHg8aDVIrhX58
cF3Kb6rfpDvZxWOCXfE6mjPm5lfclsbE9ms3ZSawrRJOV3fDF689aj6oYWnlnRxH
dEkBEEwXjHvuiY+kQji2X6YFMmVec3QV231KxVce9k2G41MF9vEe3tgThyWUYlXN
VrkEgpqGs/LsITGzweXdeBOg0ncBCDQIpbI54vSc+bXbAEU3zeCTVIvJuKSSZkLX
zpKJrPOLHnVQfd/KzUfrnx4X6yZbQmORc5SMauRt0lBq0Zsig8X4uO6H6yUyDKt2
DsutuUbYrtWEEFQvIKihqdiOJmMjk5zkrh8rXMpPvfQ8ZeqGE9DQevZ8GauSO942
bSuNwbA18bGCLsxTyXHU4ViVz8pDnTnuqaAserSXeaeU5jya/ne4+eOwKO1RPfV1
8llu7+MXrqP49fIr9rwUqJsqTFKFHMvZcHy3RUaOlQP5EXSH7XbEPPp5wB+PSknK
k3+ooWqb9s2fZ8j8nCj2Fb/LHbANJ7A3z8ILCaxnvnoNSg3zdH2Bx4d4eBp+au1A
W/tP/led7ST7eTuJqyA1m5D26Kq7KrKWnWDbUyHw48wvjqyJOCal0/Wuems/ZN5X
ITlP4SgZLcMivhZrUFOvkfsLrRSOiRRO8jvM8Au8J4ytQSaFalYYrjPdSml2DS7q
XjAOgxgncgnKHyb50RSu49u5W+q26Eee859HrVLmwFoWFkDtuhtOrzqlshaifBuK
Do1H+Ay6mzw6NZxzoAaJCs/5+Sr2kLnsqwdgtE3Rawuf1kfyVyC+p+rrnvF83cGM
FqqMblTBSZK2jkMY5VL+p09MdXbbyKD2OkPhH/mzZg9KCkQPW3NLvEHBe5eWGUMc
F+F3irUNs1Rtc2yjakb9SKB8YFnwTE1HboicxOCBk7vQFBpkrTGnb9onx9VdDoyE
sjI7K8ugbSA3wERs0ki/OUpG2ZjMj8xop5WkvIPmDlg8A7KFo4ACcP7lE01GA5j8
ltfk344jOrpI0d7gaXsX65Ypn630bSI7iA6Au3SD+MDjnqyytHPVibcCCI2nQR0j
NWsNqhd/pSzeMNcPG+8Z7YvsJOePsN0VKFcF/8i8ImaQEqYthGq8hbmn2lK05EQN
V/ffXGCMqXJ9YlbOMA2YH2AqLXhG8F3j7WywV9p5/gPLbmcPzrgxAFHEeM4jnKnu
EbJ3GKbRK6QIpsL01Kwdly7zH3cXGopu5MscQS1oGJqFSDt/BRQNRgw+h9Alf++S
0Bha0b8SbWSRk3DEP3krmZz9tXKJzsOFltOYmDhVB73zzIuOMFybYGfDuoCr/xYK
4eVa4eORR9hDkkkQAQ0CSbFW/63+InqRjPNTeKOuMBqZjnuHNKPI3FJ0amwnT4Y+
SEcnM+lNgMGrdChzNfJEaxqfsG+bIzOGp6puSI2q92SjREBtXvkTJjd+V9CQf/pQ
/farhFAZn3CuyJ4Hl9bXCI6ADNRk1fcHofa6x1AAMPPUgKutiwjLf/ZfClQTMVkD
7IwOf2g7ClMp6hVvT+7IepaursCXZ4ZIOGPwYDm2ifRPr4rotcOwWeSlfgaimTQF
2W0ASEpLNdl6HqrPRuVCw3Z+Ta9ViVeFTSWtT6ZQValpNlGPzlaKz+YxoU2nfc9G
a1kMl1QtvXeqDBIQ6AG+IQHd9U7S6WCXxp6MfgldN+smojAuNNxRcnaH9FnD4fh8
IYHwnLXe/s//2enpPhwk1eRHlueog+0B2LKeT3buab4uCTDIGpBJIYxk+sVaISX1
nblnOCeh2ZxR+7X+N0cCy+YLLOKtqtXfAyk9C+yIXB2FHRSgW7YDE5js9cumg/P/
xZuEbk+HgPn4CpfbBTJtIhvbyxpqbgnBt9W7RQeXoKZd3dTuUg4swCZXD1DjqaDB
kYDwVfIA6h+yJEh4WXgPyW4E+ZZjs7mt2Kw/WA73cawsCrWAA+/p3TbfC5i4MbcF
qWgpLIl08A+ToYS9Al892HsWfRPZXB7OTXHHJQH6YvBc+l09pI1dkxGoFf9Janaj
riKaxwu05DJInjU49vhL0LKmK56o8L+h8e6Z7v6T43Gtf9pORY7v53PETTU4mCGN
1Uiy970/vNwJpG6Ua2hMSJU813CB28XBnTq7NFZPurrGVPs38XkkH5+377wEi+sD
3tDctzukaBUOTPLF4hLwCgbHBkUEuI5CujaemxxgBKe3/6qGcXhRXxLW4Ou8ixbf
L6VphFnGm/V0WYv6mGwcVlIOMm7rhbPzJq0FTJ06y3LmBNw0/lT+vDSTbvrMa/UR
S6pbZxLvPsdP6Yr34SoRgA57JUwzc00/4Jhrlbti4rbBJ8kzin59pO3eUZ7BdmAm
3BOVoFr+/gQ94fVgv61Bu7NGoRdUqkLJ2AM0HUs0NRc2WLxFlCFTe+n3KVvspWX/
O3C8y/pbMMQ8GdxYB++x0oHy6cNi8OIXFejUQ7lrUMLq1FUJ0VNTSB4h1UtvhpHj
AFdMva9gWYkzKSIR8CeFNEDT59p3GbT/bBUNWH0PNx5gIXVR+fOXGfQOvoL49cRp
h21Go8lwex0V+EybLFV0szOM/+n2mGAxYUBhPunWitL/FMVLZG2MsT7Lr1Hfp7jy
8VTPNHEdqGIQlO55k4taePcFaFBdExQIKVAosF2pBETlUZolpcbxQ3V0FR5prR2E
jAY3UC4D1kFSY7x2f4VJsAD8UshYV8fLMs4FCsszngnDduPRWtnVcRYh4pINTUFt
TuTu7ZFgmyXJRtMny6RaLENtP5XJEtScSw13LLKtQ+s8XpPn4gIYZbQG3hbnrJVu
jkmuYAkBpGOpeNssQ578nSQg5nbDKpdkCXuYTTbbgL56kYKX0arFimS5fT3c4ZJ9
yTBlI+JKQKLVgLYSxG0eeTk+tDmA+YxbOtq6QyNwqBcHwnlpIw7ZR6bssmqlCWRj
1MGIocSa9apx7ctVelnj4kogGfm0+n6/O3pN8/6mLTgCflw5cTo6sG6UJx9A/5OH
lC52jHgBESfkkFxGLMy4c39EUWeq6X/lAZbXR0v9YnL2flgubKPpfteI0qnOHf2s
e8HAdf+WwKOSVZ7AiTCAA9gWbNAbKO4/YJTvLMgepnQkp7Ed4aPDnjfooqp6PGRJ
mYPGUMVf4L7LiigDoELfXirTcBwAaCcahD0wvMVTm/DOh8zHh0lawhyOGsi7jcrK
baG18zIXenP8ItBFgpw3C1wsCzAf5U8kcgWDxFvkFPCvHi0eo/RRWtIeriLz/qn0
UMbX/+YTyRjbe/kfxuw8sUHsto1oQH7qN1z62RgGgQUl71EP6+OTiMA6zkOHUyMR
SjVt7SXM2gP6cEiH4Lnz6mNqeejWbsqLiU1fq0Z8b1J5Y9s10abu2rKXlO24BUSL
U4keD3u7sJezYYJvj2A3y9LXcrk0J3RKF4dmFVeYDG89lESDsJAk2Z+38LU/sdvU
GLvoUMv8ur9XZDrAxraYql8bCiLNrMBEZ9OBmtr4tVpD046ZQ5CjQlo07PB75xsj
6c/mcP5R8N447Py43dB58aqE6KZf9eaCeiMu0r4IjB4i5UjxzGY2dFnsHgD7gBa+
2FNmGN6SfXOUsOWmntNcNLIWF4i6Yoo5wIBp1Hp2X271lZDWkWpht3FhOFZt4JYe
hcn7HwKxvAb7A+i3jmKZPnGBdZYA/FlR8CBIiJwb4Jt/aeBSPkVz3JIlRGRCpB8I
PctEG23TVchAHBvICeRGZp+R+beI7xu/T7tVCjmC9FbMwDPNCdHklUA3cUVlT6G/
saxw6IHszAf6krnAGKhCEGCEmvcMghNymEEnNxOsQ6q1rNnT6NjquSYeqxtTADhG
bEEefYi5CRzbuCe3o6C5GqkAIyamR+WrozmIfacYQwIS1ZfwRryCY+IHQqbH5rsC
zmdbZ2buJcY/IduHkmNFcDN3TObLNZ0IXq3DM7+l93i6PnBIFqidlNrKpezSeSNJ
itbOwrPrM4v8osUtoMgaPIh3GKTdHtsUBe7/Vkw70o59H1T9EE+q1wmYG29qQoJX
Pmw8QJA/Q8SQ+QNepFQl96SSZeONHIMMBzKs0Zn/z4RurMuuYuOLfMmAhJRhyHr7
4AZ+iawcpK3c7IjvWP1FJxlXdczx3N1dJ41UKZPj2PVeWEp41EXZZZpkB6ggh9u5
rjbkfgBXYfU058fZn5DDRexVrghA8n264e3+bc90hpIcCc5cmsUYszbT2eWg3V8Q
WQSwTI52EZFwXrmN5XZ6wNfxi0cXSdziHEPpMJJAR6lX4u1ex+cG7EdrAtxiLK42
dEOv6MfAHmrvZlZOXkoWleTs8XcAyROS5d6s7WEO61dXnBd4vCiCxZPWvuv3W5Xu
/nCQ4hNCnlIex0Ki+f86K5cg20aUU8o1xDjvDpnYyiNJvENwWVGLCuTqPu9SueH8
+2DHLSdoooGhnxTgr5YNcSbwe3iIH+29qaLm8OHnzp/jFAQycKy1a1VV2GcANEl3
o9pfT+gMyKGyWw3Z5hVA6cC1y2iUJSVKXfA6O0/DcLQm6VfWAUvH91F1zSpeKepR
DCPQTBfEj+KJ+xWVAP2gwsUgjAYpPN6c8Ks9zlWuEy101TQVsT2qhlUOK9FFR0VM
nyEVnQS/FBU91og4u+ph+6IxVJ1fTxzcQ9sUuIG9BUpm6vTrURRRSixwry/GE2To
cXRrEFEVs0i95yU8we+JpghrZushi9LKlSoXCvvC5jEh56kOzh8u+DSiMrZ8lDn8
uKEflx55IllSGxaVw+T3rgOoVkq6dpegT4PeiEFwgcn1SD1GzuDEmcnD3dE02RFJ
E8OFIyZf7m+QDJenyFsnc+4YXlU/1NpMeRpHZyy6wXzDEQ7nSHGUMzlW//7fOG6i
vPZumQ6Vr0+vBMNmb9d8VpWCqoAdyDrnIuoE03uFli+t0UXHTXlgwm3xNpiHJTFN
PH0xHxxW4//gu+2ubKuQbfVSL73/9yx0D0Fn8UCP2nBsuJGLB0VlBNCUJZVzV0+J
X/vQl9l0qme0MEv7gulUUkgxlfrRvp3aHlUD0E3aN4NYnhpTjQ0ldAJsXG6JfaC7
wBGp4axNW74r7r6615O9x9JRyimof7btlOQL525stVjPQ8ZZ8FATu++8qg/7Eskx
2bkq4k+go78WGKxuVhKkxKRd/VIkG4cBLN9FT537zt1BOgYTz9JOpC2gPk/lqVlW
uoIgVFtjdLNh7rlt8Ahz4uAGP2nRZb7ldc1Oq3RCs3xUF6rQ0iLOMVw+HPIqjglc
NY3lAzOUGI4RpGtRpryGQm62SxE3QkbP8GaprVKx3nqcTVAXjn3M/3FWZANUQvYZ
ZA7tY/uX0PpxnZi6Lk7zGVm1xP0kVK6ay7PoQ+Y0y2kujbDtLIGKAW6cufSk5sPU
QIkZ7AI40QYokquGpMwPcqRy7raL8r5hvmdYF57tbLFRfoSvCr44pgpOcXa90GTb
C6CpIvwhTcBuEApDAzlA+Bsnqg5y4azlfv5bdEdJiQB0+OsiuRM9PSPJDt5rnVnE
Co9vVtQhBcatunHbDb5Lf+S5RWntmaFeYNXK8CrKJ82gfdnJKWifmbIp05pkCTqU
ClUStB7WskFD5R93vMIGBmx1YbLUuwZ6cEGl1Ag2LVf3iLAHkTUCulWoJ3GfFkEt
z23zhPtHrABLI/dx491n1QEuTLJ+0v9xnoqoLA/vylaMxHkEvwxUxOd9E68hxfCs
7qDUiGN6BPXkv73kEto8bQjiHcrqef7S1XAcrh84w4TO5nRR/5owe7/ngBv3V96s
j1VeFr7IcrFkeK7BXVEtDSrCKEMlCgJf2G5GLsU8dcMSXjDf19eqEEZ5kas2H6Bh
JAmCoo3mMyikiZvAvqr7+zbG1hw5pz2UwYXFkabhOGUW7r0y4g29d/S2VuaxQZoG
cWrVyOmH7rFcOjUcYaEe7saTRP1kOudEx6YGOt9StQsyGXjbDm+XDQOBbJ7Tm2KH
ztGhXz2OBokXFW39L0oa7DW/WIgIF/DpIiturxk8Suq1/pmMyqdqu3Q6SdvApeN+
iicRayg4iUUQoy4mNbZNkpodCQWTrO6QNDM07n6DoBv/1/Es21FZou+Ba2UrD9UF
3HHti+WmMu+QAQtuM8gXltS6i7YyTbm8AeTaDChjI6ZwHiCR3XFz0oqrjpHl6f+8
y5b39AM3MYI3j7/vEEVdhpgi0upiUl7N8OanpW+ICC8byoNMTDq5zXP3rbTPR8l2
UStFNeXtkPmQkT7uSGCmNM7HFvhoq9YKhEMLodugseS4Vej5CYDgw86Btio+Nugt
V29ZQVLbkNVoqbc6O4Ui68s9s7FO8keJn6Y0fEDfEEWYgzbE2br5uFKomQ/VvJAc
ZpXQVw1EGfOSNWsfsFKyoafchHlFDpLhVADTa1QUOx7Oa9O0v90lq91k0t37lOAW
3mr6RB595eRVhbugeUTg+M+vmZYx6A5lZqM/8CQFvQEbsO6rC94EcYvAFw+Kb+sA
dY+gIlnrbd8ImFjAqNU3OTHDknyb5Qo5j9Kjl1CTtvBBsxlQB9w0T+libeHSum+K
Huad6xUFEgoZ5quHvPPg47hMPFps/Wabhbke6mMI9U0W4k4J4JDGgaANyBs0Sjug
QCOMFmxAkX+bmMMKryoSRfLGPglaLvQgfUb5m6y6YEK2DQ2Am11aZpnB+Yp+32kJ
ycX3nIOMu9GxJbZrSU4+qUNTppUINqMQpdcHY+3U0JYiQOGxzSYTIQ7LXQCTWe9+
S7b8FaTuKTLUarE4hAQwQ8bx+AoADTrN021Q3KA4W1xdbSA1IUlAAqR4vV5EQs/B
cIOspzzNWfXlKwunas7UE7BV/xhWIzpvWjP+KnThOstFF2LTgaIshiSrlJ3xsCQr
LJlScCxfECC90MZb2bAi39rRp5jufNKBJWdq7MihHzZ3cZJRShpHWa68uoT8cXS+
q64Hic0fSytj+rjPgbfyns+pIDStY1PuDG9IvIMnpw9xa48KtBIi+X/vdMSk02iL
vVJ+hKFRKfxl7xRbU8WIu0CeTvl/pBTbFUDl6utr70etsaUORo3ZsKmw263fhk0o
FzBLsPykHVxFa+0NFzzJAD23M8yA2rln0CTMzG1H4DTotOWxvuSFCaIGdul6Rtc3
JnqkGaoOYe5l8yzuS/i/R9Qx3i77vq7z/686vIlg1yVRhXA6JqlITZYQTpN0eDG/
KwhfJdVhi4Z2+5l8fYrmmedN0ALJkFH4dSID8whNEgVvoFn6aRiP3mJ9my7Mqr/5
Gn4xwrHyvZD4PAD5oXlwNf21lgTIU9Zz6FKRrIjJ4CQllmQHxoLTUZ2sDNZ2aAWT
yIkKZgFytOxvTmCXExuN8qQdyuzTl+zP4W78ESesEwWhsEt8cPk6jkuNXV/0dKJ7
U5VGRn6hzD9NfXEpZ2+7CbCxRARq46+soApxQ2r+3plI9kdPvJxmV9j8sym6+8eo
PIbxvxzo8ISfi0nlSuJFA2y77QjiErWzz6cg3Ab4f+0JozjHZRYjWAiwIGDECuEM
R5GFVAczG+CWAp6KlhNnmersyPXloZGXNTR26WmBR8o/2H916bVR1es0w4MWF/dO
Y1vyx0RAPDioxKGFjvEUawhZ2c4MPgAKuI8AXbtFPBiq0gBJpSYX7StKNdpW1KzH
gwrrTFrYKGZ76XsNL7GqitownCUXyQZNh7LjhSx0KCSXTXh4yW6qM5PxY5EHzuJC
+gK5BUW8M2wAOC7GyVB3Hjs/iGFNPIVuld3m/YGRL8WjlCruIwGPGrYbZp3EcDll
xFqzbacZ8bDxDvwJgqvRhNwcaTQ/Hy+QHLszyRzkGlKN+QrPoSgxAT0b/J5UVa6p
aBoqpdeV6wGOsQDyM6OszzUA/tLGyRboDq/lxEtjAtZk5hzQ+QI+uNyeuI7nD5bI
dGBf5lwgFYIZ3I+Bl4NIfIovZgzteltE6xDLfeYM42XnzHQMtI/IBv2GNHkDP+Vc
yd+foQG41xjavm7BKNbynd3IzgGpjPotdc0c9yPmu2YxrBmKu6fQTvBjPKC0pU3l
liX1g6xo2HWnbjCuKG33EkBXHHG8X0x/rUhsFB6QFDuvx/GQfl+9iGe7IURzA1VX
/er5g28f5uriWBUKlygoBQO/Yph5wcsZnUsbdRgZ+2KynJCwpdDc3vpO9Gg4FQ3i
zG163RP/uoLHGrUv4IMxkTqzDO3zUmlfhiCiq+GTiZhzbWiHgfqNVVR84UEdyGXl
ustpAiicME1csKgxTk6l8INH4p/ZwlJ+Y4P57/fe5bnjhkJqXc+ioNvUMA1nckFz
T3XcY6jvR6Mqo30+R3v32OESEm+jrmYqF9y39DJo2Fp8HMINN2AImC+CD0PJiixV
BWPw/urBrqMz2nATJE4ExUZYw2PdHKCGDa21ybyqu8lozdUa8zB4Bcd8G7ED5TEW
hyxCrisjz/SXDnWCLorb2n1xs0r1ypMfVbZakZBByePuHOGZnnwgO5mqmiIXv+rx
lznrYHBhDjYpXQGe1qPNlxOZ5OzuIbH/fox99T44RHpaLrfVcODrkPwpyFmHGR2t
6WbfpdpeftdDIF+cV9jbX+2r6CZCvJy2YYWJsQcp6a3emwv67hGYs469O4TNL6cy
zgEaUyI4m2MrrEROiDarFbYRAsDCidv/g7qeW8UsRKsa5UuahtnAqkO/pKvbeZv3
AI7CG6TK8arzi0sGzkXuONIHShE6xHPvyyjCQoRANHZ+yOyS2otvgOITK+1j6aTe
0Q8cJcKsJ61X9Gf0h+VZipVRlmuT/MOeRnbzLmtINBcw7SEou7ZCbfPEkrEhICuq
4xE/onlHoyIdwqpUVrol8MflX9z4tLOqzOD04DCIJgv6oG7MR/MdXlWF/r3cNEI1
pLHpBveKHTE9rQbSWs4+L2Ro/wlv2ykn3I38l3T3Lwdo/ABrRChr9+klY+dtBIKP
`pragma protect end_protected
