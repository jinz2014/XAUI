// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aiBREc/8OK6OLPkmBv2sEBTq6BHr7cY2eMp5lcgKlpD7N04/tdwzjes6x+oH/pdH
r7iyeaNvGQS+dUMX4MCVGJt8a9z/jtLThnJtd2UGLJae0EIus997NR0t22SbiO2m
HGN9DADY3qpeBf3i2/XZKknQmtnRTVFenltvhePBmGs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 319968)
FKHRNOm0elxZq0/TD7HG9U86ZrnT+T72s47661JM7Xp1q+GUbWQ4u9JRWH6pVTF9
A9y+OKGhvtoDNhWAXimlwtnSfsDwKqT19e0aIMxQ4/m8NrKZ0WKEAn1p6qsLSYCQ
TgZtdLQ2P5GNXfubqd+xUISqvz+QQkO5cH6x+xa52H9IY7kIt4M6eBkbRwY33Ey6
0Gpbb92Zi7FUGPD3e6KfG89vkLZk3JGyg+SUQj+mB2KzXsUQ0ir38ttzAVSsuwlQ
pT+JomaMCfwRTTjyy6S26rSRPhihwm5TPSPKTQu2ZTTw6ILQBl09svTh6QEHsM63
IcZ1mLdpkmS2QQ+MPG0/S7fT2Wre25GNRr3YR4QxNRS92y6bF1oIRTDMisTXq4ie
5MRiXJMfTu4g7KNa8DW2TKutqzzZown+1QLwnDVjBtF5Y9Oi3pVkhJFpmVz07V8R
eKds753YPJ4GVQuOYISHNWvMWyRs4zqliLYYbWKJceoT9H9rK9ju4Z2ZPbVmiavQ
LgQwcBs30QlCDRUnbDJyBCBCteZrlsaNuN0BUQKMhg7G6iCzNEdrFz70Nh7t4SZU
Es5uqS8e9lU0tIEQMMd85sgH+eVqMhUAlfz2sjchVxvBUrKf4dKpvlMeOP8E5QSH
1EXmNgU7ec9KW0OaK3hAkXJGNtQdJCIsN6o2XT5rVTCGZr09ZgHZyl2o/7edtabk
qzB64f9UFLvyEmMKuEJLq/9mkO8bLxsHm5guluuJno+vcHGTKKbTaKR5inuAMjGh
7oWa+YjGt8sfeCHFhqUjqEDqwOjl7AAW8YcF+srXDzPeh4e4xsJMgwMRm1bBrRRq
WfdearKoxd7cUftAIuQOegEVsOpOQKMvtAyKfsSJ5VcAFDC0vBMol7TSjP1DNa2R
iNA+GOpgglw4WCz2NAVprcs3Kty510IEkpkgZjUoyIavyTQ2FNvRFZwXzsWw/1qp
vf92bYSF04ATNK3fdL07T+kdwOaEhXO72/bm1y8tbq16eALZiLvSDzKbPLo3ittS
YlIZOtYzvF5CN709iPpfam0GbfqP3I7oqa53WKzwFJZFV6Fvp++aadSb+TrxurM/
89qVJ6G4mU8sBc16rQLparPEP/0FRbHExJI/gHq8QroZNOPn/uAFRJbCCXszCqzr
hH8pa05gjEvcjJrN2GxO9XJqnTExYLXssLx0s4Qm5BMXAglGlmIqVkt2t87m7Gwz
RejKB7W7vMyeUybMu83QCAou9DhtGdvWs3PJ59cWPxAWJG3sfqXoYfiHPE3OATbq
p7ZlTthxkBhVhntlfuIZIZ9Z9T1Pwx/ttOSbQCB8emxOhgdfDsJGrSk3k3GW42g+
YqCG+CSn11dCtugbfHILqtYLal5ujC5dAcoYbNCP4VvSbJd3UoAEG0Levma4+oEi
JiKiue5/ZZLmoxltSkr4IAZSSJ+7PEjpU1xShZcVjzgMujm68ISvdHiK8XfYqD7P
AoOvOLLYrqAEH/VeErm4A6PfHD1xycmUvY7AyJFVecMc9G8ZPt/5VS6RTD/D/3p4
nqXz1L4L7bjw1bfCtgbUX01wa27xvK9krq313DM/wXgzsKw7kMj/yR733Kj/8bqJ
nQozvFiszKORosG6BH3akVw28YITyCITeplXMjCL1oz4INOhM9ap75iUx1lBEEpx
ZL5MNOC+TgT3nIfFdQE+Yppk18Cdx370ShZzpDbcmXo5g7kJ8QeTdWFGXnrT7IbX
NVHx9X3m5DRDY4N7o1WB+oEYaXfH8A4uYtcXP0CQfbRi4Hcf7hKgczFo9nR1nNZZ
IRB5QgVRW2c/sO05LvgNjXWohejve93P0tHkSVaYRxscnaeEJs40qpCaOOJ+DzNy
fNn1V+uE+anFJ9/PpIzoIKkews9quUviTFCx2Ayz53S3BkPsU29YQ1XlK9iJNydV
jyy+KxTl5prg2wmdSimRi1rrvRMfhohj0wcA5q4C6Bw70XcdjzcCPtevOQ4PI7mC
ZgaMpF73hGTcIPLd+otsgz6lFYHKLZRP6ngIKWbmxauxe8fcJHBz/wZ2/0ZDYF0z
wxstskP4y+QVChs9xImOeucCgESZ4V7+3J1x/r+E4JXAyyLSJNMAYrqdb8gCil41
C43ify4V4nFPwp8s0Boh1mvdxqnuzXQRzAyley7QN24qGCFM7+T/3n2U1i2oWHyK
BX1UibrVd2YPyrCN37vmyktU3w4yKToYdaLx7r9qQsGeDwH+PuX3AIiwYNejGetz
wSC8e7X66FMJFB9uOGTZE8M+u46+DxrrdUgG1mNAvuq3gSycK0wmKFaq9/62WoY0
UPvgscob4vuIIbmbl0swfOnbQR6zXq1b4cpPxUtxpn7WYc1ZH4xpjDJu+4GydvXV
PnKhSE1lDLbdqFEdtWFFAr4Cg+fVtcdpUbpEcp+EUyFbv0H7X3J1RwZ2sS5qDXNk
uQ3nKSGiEdbcoaSI4Jah7bwhUIUWnd/rUyS9+91j2TZI8dx4H7d0oLBeklj0h+C0
5jhjJXwE8jSUxDRIOeX+x9QFAPQ1OMiBcXyVxunHkiohPpcrppVhX2iwz9dLEDht
7p/ZGH0xSUL8p13q6X+GLROJb6o5Ok34QwJyxhWtfhByiQrYtcC1ui02l/bPhlUs
Gk7C149ONCB1DEkAz4RM4vsGdqPdLPPV2xTFya9PlURNPuOu7r6by6oBsFXSo7U2
M26eB/vb6peiP4tbu5+evZFJ3j72+MRKROECeeXv5ZMfEyA8VKgGhXoWB4MOLDfl
ld3ExuRPq40G2IFw34wHfHLqo2hwWxgnqPVCkcd17TuWDLdT50LYGCJ5aW6iIEw4
SVNDR0G/ZOVaZtPM0K6Die+ZLEuJvNmSVj09gld61THTtduGl7L5lgZkQdl3DfVV
Cihxa9GeId1764klFFhw2fzZJ57mAtmpsaajvktf+etNcdEVUmRd5qWJLeGxZt7x
9OewW+/t7upFsZiTw39cCA62l44gdk1Nn3V+8sLG2kDSmwJWLD4biynmw9dIcmER
ZCcve766AlzzYuyoNBsjKGQiSI9P8Clxj42EfYrUA5LMW9D21ka49XMqKcUZE5e2
C+qNdiCLEeJ/BOj5iPZC3lUpi3Qjc4/TsvjxDBwADISuqu+w1k1NH/Rm8FqFgvLC
JAijZ3043zjPj4iMCtCMx61YC5LRsK9SpdLJCyMegVfEcZc48DzxbFuXo5lwbGbd
ZYSTNPzfF43RHB2uwEfYcJuDRw47fzlMteTjcEH0CxGSUcUjiniXj3ISAy3fhpzE
twilyDKUwc9YH9oI3q66idwz9xGa/o2ShpfPUx7ICSORKeHjV5/d+VW+9nRE66fU
RI4/1vEkkC0ZHlHfoP61jZL2lspy5TOhJgFhYqVmNV8bTGBiSj2hoeiXZhXU/Kg/
RqemOvbQDICI11SaboQLQ3EB3MTGmKnNGAEHgT/OSZ4qZ6nQYdK1STzniZrv/dYG
4tcQM6wIfLa4vd+AvMUWJ9umWLEs6vLKC8FUial4tHyR3v+JXCuJdbL6y+lp3nne
cYo4XWsoIW7Q/ReSFQUNxk3PTHCWEbPx6PSHNXwXWfQPXBVzsUIUuFVHLtgpLWdx
d/oYbFlHpHUCNAr/2CzCkOIJJxJqeLDao3y5fH4gpIT32LVnoy1OgIGs+3UgE9qp
zys+V/QT0JayIZWo/EYfyY+xvf6Nz/YJd1qvKumXoKSbfdRA8PpupuN3XRTfnU8i
vivZkmyiUWouomnAJdTypDj1CPAK556L/IIbmoRCPPvVCOWIEqUPaRolqtGunNeo
lSm4iV7GtMA+ioS8r5dVc0szdkkGfZLy7kMnqO+hxt5g/Pas7oRmRpWoU2JUbYGt
EzEgRWw5I6/skQ5oCDvlXzsI4K7NVmDS20fl7lXzcC7l2pIA566Pr4Lw6qpi0Z7A
8y1yelxejQOsGVDtIdEEofNMqQgjtKpjoxDAf+vjYElFfzcG70SFU8CKhLuU2KXw
YrGlkyCGOnALnDMTeX/ecJTsx07Lbs+BOvAYF/Mhveq527VFOki1RBptt2sMKdXU
G+62VaZkaMYmqFNWvwUvVFIJqiQjK841/NdQNjLLokOjsOvgXXCrMlowhLp/S2Y1
Us0NiJ/vRzdErI2V8SuygIxDS2WG2VRgOYkUXlnqIezoPcqu2sHraBHa7OzNMSdd
pjqecseW5ASKe/YTEMnLBlVS+QLRlv4/9xqyfiV+jscD+dszbbXXoJlkVZiolpzX
JOjsnt2gMxdvhjPD2MhjNpOJbcB/DSDCiI/+HREbVnMxVYk+E2H8Rww37REeX1Wf
IT0UHnYVOmCLN02cmiP2XOpajaeT9HbVZHM5yhV1njdTtpdrVi84otu/M9CAgJ3+
obowIQOKwI+d8Nepjty7tHABrTG3m2XkxJDGsLo9+dvXiMz0CH5HMJCbOIjk6vEl
n5bxmOaydgYy5YVHPdJqmScXlRsPFC4YgQ+F10XBObmyE/z8lBYZH+ZzfLFfKWAE
nMRqWwHGb9gHHhzwIu3cdTDB3//NldAFKGagRZo6X5a7WvWEYShRuayo0mfNY4v2
SZhwmBhXkh2H9EkE6fhYCyp6CJBpzKPXzfckSxQBJOze90o+DKskV8oh1F1o1XX4
zSxt0F3x6fVA3fVX7Thq8xtCcdr20rFWSJUIfAp3/U68nWBfcCbK3vUm4zCUpcwZ
v+nTmp59ohJFOrKkNGP0qh42no5Wa1g2e7Lv9PtIZefRNUeVxnW4o/kpl2i1mRNx
BazpvbmXvAj1i+U9Iq4doNk/e8BBAD6fk0Aq4XI1UTWq6WA8gTMUcPambaLGL2vL
5Cz3tjqbD2I4l7WlWpJyOfPoGgzXOTuXS4GOz15uxLVOGbExPPhMc9KXj1d5CUQj
UWp5qn78t8suRhspJq8j+PGOePvoTghvbYlYtk1SGqdpZbB1jFTmP5InDHKTA8ob
mlCsusBkzjgv77L/E0RFGJ1OXiwuB+NPh9DRewjDa1h8Ob4dOP2JqkJhVQ3LdKqB
BZYvr2+FnV16WCYU7bJE3YxWZZ3TrHGKO6L85t4yKYc5L6vVWXMpowQ/TvxY7Q9V
Uqyc3ixO+mG7zcjbWbHc5r/7QMUBoNT6oCprBmhk2knl9ihLhGJKx0qsFK4csvpZ
YhywuW4YbIGWuhlVPaHxNZkypFFgsuxtaT+d8PORdwjDaRkUqyROUzsJZqJI8aED
IBA5KZXBF6/ICUvN1iE0zJvHdtgfkUmwD8zLCJkxRfZ0uMlyT5yokG21s/Dmf59l
35+v/CI0BR0XoqteSxagtWwdawgnKtTMKaJmg0IQHZiV+wWfaS/QiQ6blJSDkJov
LLXDDAqTTwzmck18Q3gtmr+eOtsI6B49BuVSLupWqr5sJEEDbfJaP0TpVzUhV0JG
mfeBNgmkgQ4Qjix3qIpFv/VOzsiyLU5pgZ6Fvsk03J69lGcCJoIxWVbmPiCb/En2
46v5vPcth6ChDonhpYKHAtnM7sNs5Z2BDoSTenrsu/9pB7N5KaaEzc5bKEC1Bavu
BrynYaVcb875h6z7U1osh/+ZXT6gdKvhb889xZLu8lfi4hTS7UZ+lz81dg7lBqhi
bzLHlE2fA5Wzi7jEywmIioKnKkBBINKKsu7AEvOaGYmrqk4lYAKEBoIqZb6hKcz/
jQ5lATlCuI1vCnAS6yBJDhWCz+MPXKvunYHl4OTLbkYFeO/H+ESnrjEJX0ptfhUU
lj62EhFwqjOZzLNGHdXmGnO6SG0zaeb7o87zbpiTyOR3dor7DBoE3zqtqJOrAuB7
jpoebnQZyDOQdq4NElHj1Dr+h5hDNacrRpp6f8B1veO9TvyBfbtlYusTQaN8l++T
4+JGgt+02mCeT9Y0vOJ1I84ev2iBw0iRU0VSSu1t3vByHzQAn5Ho0vEWDOV2WXfE
6dodcD6uPVPD3Ffpu4RBwwplgOCRlMNTjzsHY1kNpE+Oe6g/+5VIR+5FjTdOCBGm
rdPhvGCeT1vxlBQ4bx6pBnJ/Q22bSVlhS3p841ftmKJyZCdKFcRKmnhaaXhuhtbZ
BG8YoBXA1iT+UUdtR/9FYk7Bk2cnSfbmMkJmKlwQdx8VVxYexKIAFwKIz/5dG+gK
mk9dlNcDWSueDl+T1lm0UVVfHmIU5MQBGUzN+IaLhSo6EVeiro1rx+jemhYqNIiU
Kt53+eWCpX0WriA/AMcSOJkEfA9PlViLkFcc1/aTFcL3X2Tn2+OUtmVHYNTXLJjZ
elnmLfwvIyZOiv5A6dyDgFNedLDDem+Ev8XqTChMojyciwMpvasX4mKDNztYgYvV
jypHzfhZPVht8NDN2HD1URkl94dlwdB6zwgxHu81FAWih78Zgd0JmiVrSpBhXF1v
JgBTnylUp4xaksYQGmoaeWlbrbmV4Nz9BA4UCUYIMzpe2zUa/tO8PrHNytWkMD2b
znEU0nKeY5CLeofD5+FvkRVMpaxRUoHkKWbHDi68W7bzC5ZJpAsxTgBDwUNgyudv
dSr6UyhDfmpfydbTZDTtpQY4o+58y+EtQas7J+uFVSDU+4wkfit5MohYafXKKIKQ
IB+kgaHMjA5jByFb4DP+G7DdCJRfcnz0LbBe0iI7HXaUJ3UC20vNBWXlzvPpu+lt
dvbBeE14XjmkegtsNc1NNzfqAcklu8Esi7kHBvzRuOHu7Ud4c560pCDuBNFk+wPz
OujE0rDq2NpNamIw2fjREkOdnFPre9AGcLtDN1yJr78hU/w7t+hnJuJsiYHScRk9
lOERyV8pBjk7Lm+YfXNF4Q6dzgl8gxT7b5PmzOg9SvCbn71iZ2oPoX2C0b1MRN21
s3rzUm6XypSbhaRbbr6TgpQpIH1nwRrw62bWt7nTsOB20t0dfZ2k6yxhjpNxVwjw
76UjY/zbMss+S/NKZy47uQipmRBNopMe+51wAozkiasRcWJa2YQxjnmLuvhLq7rJ
ydJ74UPNuKEEdb6i2g5z4+5lgJcXgsyOngMNRh9Mbene/ZkV1PvMLv9ILSMR+j4g
a/u5YTSDUf/pen2TuK3BJy9TuDTXJCBdoOqMeVTW4Mc+pr8aPB3LpIKTpbx1v3Mh
P3adIiQ8vqlBZQe1LmVbkZqF6UPeUdzk/SVITw8MNJOjKPQLkbrMClkYCH/H0Pof
D9I924pt943jpbd6x2i7nPvQNavq+DVJFxGNkclwMLKTYdeuNUx3PU4UNOy0sFOy
XhmnNDnmlGnkttV/HrW4LO3jpEjSwOJ3kq0CtK8D+Ly5p9Bpkj3kXamTIXKFtJAS
VIkuARoguEFaPUKmCQYgjbqX4Tg+uWMDH+I1Lq01W8Hey7fnnA3ladj9OusMwCVP
Pe0B6l4zzLt1B7p9MCnAlNii9A9uSRK4P87bPN6+O1qy48Ke8+DypixAGNwyQtAh
bv/asxXaR9tWyjZpd6g4OMSvTl5riWf6W44OIvIO2u6yzLNGLroo52SC3Z6hPyqs
gZyjSxAcCh9z5dFSfFgoBQgWsa84pRUz5fST7Eum40vjxgY/N9H5CTxlfKxeNpBX
w9g1imiAZoX77xMYmY3FKqHixcyBQcb7cLUWdXxsSYgihQr6NV8aZq/sx5nCkP1o
RMUscdb16yYIxTlPpZP/rxRHf+G3ofkgUat1OHNF/wOUcHi3Bmv08RbQg3rfy8Zs
usFonVTpW4e0Fdwv3l6H1Ad58MHDAftQmjkh/lYPhQhP/6QtOd/wh0H1F+RB4964
8zZxNgAgnnsq0S86F6AZCji6mftTmKnn5u1WSLOztQv8AK1JyJ7h7BDA4cJQ4uYf
2anMplsxo0WHl9ExqJ8rcYPQTDE9nuu35Yh/70ZAakir9T93VsNeCxretIvh++yU
ZzwH+9BfiKhcAocomvKMTsxHK4002BSNgtq0CZJVwkf/RDMVoymumiRY6WE8dbpS
m0cJWDB+E8paV1DJndAKycRivXpWnUrFbnw7hC+wQqRXo19qMh6KBdDjuCwMSzGC
RfKTiMfMyFM6lzLGo3yov+OAl0LBsubluiDgp7GHsXKdIgET4sbHUz+7sSnjIg6t
XHpQPer8iNo8iyIWMWxFjlnSKA3/cI+y2gKVc92rBEwH6i6xkOkQCKNZp1MZTvNK
7TXSWCchWCouddTWL/2qcZ0He/JKvoLKc7pUk6a6X3glr2LTnhiLxyqH8MV1bSz4
O2zKggqnjQZfRBhCkUjjIZXOkhLFa6ssK1Ujjtd08ITn58Sll0uBGfzPCuQbLWS6
CUvz3h8aWvjBIrWAw6UXPPdXzXgRe733V91kvIlW9ybiYTQEjbE8FHIQ12EJSsP+
1/8kUvE3DHBVvsQEEaoRMEXY07PSlG1v2Fw88bg5IenpeSqxQk51d9QufV97pjZk
s/TTW52bgtASso339/t91APzGcwN2REQL53+5iAMqv9w2GzXmZVRu00v31V4Zp/u
+AkTgBsH1DsLQMiCtEFkNHxTXqC47ukVrDkp/PD+SUP5cMCwoOUXOmnerSb7G2Ob
oEDbYl6XF36tK+CDXvKR35pYApbwGIOZVxQDUQ0ULEZNlEx2ZkgKvwBHDbHLSgP8
w6D0zfVByDc6Sim3VIkSV6+pUC4xp9aZWzHM4XyCrmOfZ3TXrpmJi75wW4t1QMuj
tBrEb9O4aoQyUViQLOozkyY9HVsdkKm8Q26ugXCgHumpAjoUtw9ffwx8HLkILpwl
+FViXKNJLQAMTIurxKDm3XlkPO2hyxqNbOFEnME9mF+fKh7S71IZpMwfQmiwYRPq
JgQGAg+mkmlN/yaVoOiRcs4J+pCFlDwTsDSW2aSxkgoZWxfjBZRHmffgidIDzRGm
O3MjvYnRfqR0pyQE3tCjOBbSXNGY9x3wt/+kG2sMd4ixI/mrPbRDotiBsSWZx7A1
lRkgUYbn3RHck4Jc6vVQOFq3XYrZxrXm3buWurW/KanfzWaBnPNbqp9icebujN/e
+oOwFXbDc6M2WZk1AhaVbCDMLjIWX/YNE9GldsUcqb4qjajYaFTeoDqZhLvQW0j/
143DnLUtWovGRKEpd2CnB21GRHXxQc0jdTx9aIYWu/+S6wQQBtB/UCLX/agaywVl
4HMetO/eMKKfKIAcjjbLZOSFSWbcuvjasCp9mzKW5q25l5n9udNUoQA2SyElDbH4
XvmH79jg5biQ5D0U/YyaRas6qDZ4aWiApsDNMg4nwbiz7QlvZU0mx6Mie8rST4IB
Kcl9dXdevOSkowLcwpwTulpM3fLRkjIY6aERPqEHADGMBs0ud6scQtFIYL3gFQw0
+3DHCYI9+gYgKXsnnGLrPIyVgpV/kFKI10npUAiQ1zVw2tfFuzsoZO03rO8VH1mP
gNM/CNV6tIAWxPpU0iKidEOYe8Y6R0zskQ4K4pSLY3EFOVMoXu6DzC/8gwGSXBdv
HdbeNeFs27DGNbqmNADjrYx45X7tO9h8IpvSEO+Cu5o4bHQlyN6mWEWO0CBGT84u
vbbrrf2FxRkJrvwBHr6r8GligfyxW83etoX8MXJN4PCtzMgTVgkxUQtS1cG4CFAR
Gwuf1gAJh9l7uK866CYudtkgMcUFAod9J48Be51r6TIZJDjh66EDIL8JcmPwVUhZ
+W0YO7D8LwMtrGRkmpypwIc3k5TcIw2jAEqLnShnuliYAQWsk2kf4CxsmmKwzKZ9
lxAuo8vmyl0ypzCfR8R4lvmij0vtc13uc6xasByriocwRVXCI2C1MTqTC4GbVwiU
NEFlVcE0HjD4KL+udyxZkeAtxx5m91PSQGYyB57ZYLLSQ5K0AaN+cJ65Hpip//YH
xyYfeQFtSoq1lMwabE5c/3u1mp/ZltOIqzMwKYdsJeGFEN9D7y3CqWgUtAEEvHEz
vDEF61s+pR/IY/TktMkw8hFHk4/llGW0JCYruUdvefWceEP25bz3o0ncb9omaAPr
I86Lbfh51AMoBNXQ8tqVReCOY4p62vZxi78+kwkeK6POJ5df4JEnSQnwY9jBLb8r
6XnT4PTviHkdlKEPTl7PmM1AouqRAGX4YZAsnWHwIHWCKlJsOnFgJxVNrP3ON2P9
HDyotzl8dnJegjE2BBZKU0CxjapmxNlwPg2RMABWx1ltbYTIGfM9+xa53Mr4q1u6
iyNaPFeAeLgh00ABlYa8yyPFHfScJhUEDYINyFt0i6FAvKNsjoU1vf/cEomjB623
be+A+fy+0NmWIjAhBoGxo1j38512XTqOQfg3VSmSmoHSDLbCzlEJ3TmKbDrhAolK
AbOGIvvA2gzkd5vFDOmFo9hFKu5UQ2hiXafeg/dTVt8FLT9tJ1IfK6iZUdGdw1e3
3aSJcBiAcGCHBIEhT6RwWC6hRFO10tqgnqrlhOEI5p0zk/GzViJLyTDt7L5zVgkP
PN9inieJjuzD6zfrhbKG5JZvA+Kgau5QSYnIKvDnaTAeeMQ+T+Xx//2MZQmWikvK
n+XuYj/hpoBTyS0dhQMe1isCMsySkuvlqdcECffstbbNEeWS4GR11zw2yLPLKW2N
SxIa/orvQxsRVE9dSNHLZ4LCK5JLZ9IlHs2gzPlaI3zNc9E2rK6SnvaOlv899uCh
/8QxzZZdoIb++vVn1FPqFIGZLN63tvyzAqzLn/zvROLve0Vg0VinkNyfqzxdDyfK
19jyptOtawtz2R7mLqW3O7NZOUnxkBuMkhEWxnhwLA7kROtzqfT75oIufZBaxVij
R4YHFKejSch3DqY0pTo1GKa9LWNaP4bTIghLZ6dkO6wQqDuhfqIKE3pWBgmIzrY4
srKX9yZvJWG2dpGjUD/RDv6F4KI0l8HrIGfAZb9Cq9oHnFU020FHUEIFd6pvnRxA
+HFfzJCge8x9c9n+Ue/oUNAf/rlQsgKge+5ueHE3lFFslLYbOYznXulVWJ3MWjly
BEKttr9ow92PXlfYBnGr7iPz4pot/ckHOHRbkm5Y849sPEOb2dJR7xMFsiz4vDMS
uUOJtcmOEAcY1oofuLW4uZDDV4Yx+hgLFrGLrvoTET7yREE1U2fmKil9ECjKIkqg
1Cp/N/LpEGJborw1JpPQrQMfXlAKtAjPasa1+xVQz/CTUvyZ/FRmMJc8TY624Ult
ABT98HEdil+roSUGmy8pOpGsNVlho4p/uUUzUqrk6Ank8zgzLzL4aGt4ualVjw9T
n0jQ+oQ8FsPdH2sAcejgGTgRiYqVjbFGMCJnDzvN6ePgRLBdBV7rxzFbXrHsncwZ
s5/WZeNxPAaq2xQ93RBV4b/wzkx6bbo5kZ3OP/r6ucjOsBzJU691K0B99cjSg4ig
ZepngbgUA4RoHlmyQezSc6Eg+2cz+Uyjs4mcv4uuMVRlAPii51h8XxJ14SCcg5FV
iTEjqeSaHWSxs8BWadWe0k0Pm86Er3Jj95VO7FyL+fouUtVge8uCBVOch0S4Pedq
/7DUbCH3zVfDDlkJchy6rGx26FAxxKM7RJUYaGdrpqNyaTy6WGFFB+SCx0SHiDVO
FtRwPImMbpj1jyjxEcsAMkKEQLgK/RAlTQqfqIxuNtPgYhH5K1vL76CGtZVoy/vL
/AyRaf5ZP8Mok+/tH8N2o87rnOnTw+X9jH6l7zlOmp7pEO08U4xRbWl8aMNHiOId
mZbXuHjDoyXHuynfMBYpx8rHuDCbFmlb7E83hYor1JVPhkX48S1Y2vlwrzEogKYD
J2FZkuCbL5bxH2qZJTJ9RmPyW13/ZHyMzl4wsmXD/a5CxHYkrql0iKlMgYe4HG2E
a2mD8MQg33MmBmbIwFp786ypud5Es8PqMMRyu2nr8Nrtdp+cpur57+6PVyjnx9F4
3I9xSLWOthQb1t5IeinITDhv6teFTsEsUYi4H2bVyWWn1hOI39NW8Sop2v28d8FZ
YEAp/dZ+vucllDOOrtutDyn3Xm5qpB7EN3YDYwDXgE1wUGVWs56MmkJRxXx/95Rz
BCAQ8izZ/dGcW9MaB/s4hcnljKwNGompnlJNPBCj52GSsIynw71j3DQWg1wub1Hs
LSzUD47+B0/jKBmDCyfIKvK9rR0ZPChlxpnsf9fOONdpKlK/bGBvDliR//Lb20Lc
/e8lN62kUqdjF5WINTmlxfI+O8xFZdPE6u8KjZWYY/cSj+jjR+u63v6o/1qwkk75
GDZ51XT/oNXH6cDbfbEXrbrE/qGd67/RQ/cK3D24S3+RrFKoxhm9V1pdl11yh/3v
SibBUj9dLrYgZOopNceg+IesN5W4+u2uP636uqLd9LZh1WCKsFBcNAbaoVZuEk/q
HoSokLw+E4C0fgH7BiB3CcXc2ur5dL6IIH+bpGRd88vDFh4HT6QhRT7TfXztxYSG
2G/1Vq8xbTqxfzrlzmupeHNpujrIw9qsIfw2Pamn2oFx63KZgAoDcyfiRkthH8Xy
YdVF3xNtkiGX7oS16w20hzmnkYimFkYSsCg188WtajESzc35DQFdX6odqB45jenF
7DxjwPoZmBJfBFiJrMQQS+qBGixxcQ9hEKBjGN920p2WnSKWJcpZ6efareH09xez
hkg6mVi6lMbT83qxYRGTKjbyZkAkuxxSkJa47d3re70Cpzn9d1C6FK3ZZuwa2F3M
0Hkr452vYGkCPNSp7RCJUWRUMNGhF5ksyz4KEkiQORd76pNc1dSD0EF4DtZ9IKk2
lxCrOnXGvGQ4SzOk0aE5z6eayGWzYM0Z4SxmfBs3GrHVKXlUt0tdSdNFFRZNX8Vh
owI++TSLON04P7ZMbyo4La+U8P2SLvT75cbd6fbChu0b6pk9Xss91m2uKuu7t/kJ
aaiHoIyM+PnzTDZ7T2AImkF78nK07vvmw7JOe4Mfw2HRUNSO517yP4QVRbOCIMop
9Kt4+XjR/zHFAvE2IeENVqy52r60Nms6Tu4IE4j40WVRjtD7Hzs60WHautwYQPFX
De9uwDyQxMg3O9kGS//J4GInm+mzqfHlFGnhHn97I7mqYWny3yMueiAmgU48YG3A
vxS6pdIlAHBuszkE0N8IOTblUNLI8xa8jpsQGBf+JkbkCinRoUA0FlmDv3GlqXZy
QRTjZ262fhOTb/xcH14ydZhJGh1idQEne2X1YpLdZkO9T+KU358x/2ajRSmvZHG6
8Ehxik4HOpI54gho3oiOU70zDJi43sNvoQJF6Cq4Xzp0bsWR/E5m6zMwPozQdKKq
NB72eCHvsMStf3n1KEVZYTqzYBB3BAHitOj175BmRsfDZHGfY3Y+NYwv47uxCpgN
2Us9XHMr8WUmOnvJSIE26PSNEr1zAcYEujr1gp5yDMB/dbL51Hyx/SaHy2u/YROl
e6IOscOZV/mp5Y7izFT8NZsht00BTcnwVnakSZJTOaV/D4gB4cR0bHSw9Hr1BoiS
wwbTuQrqVVhuX0otQ3L8WQFV9xlXCNARezncIWHiH14LVejx1c0wkmWtTL1iJ7H3
jgt658n4DLxjG9qR7NXSSt9RU2eTAq2phn3GZPQi/NkRhSeWPy1UAL20XZdwSX5e
qERLXFFCsC4XBye5EzsrJuBCbJq0G2hgpKIzbVFXupCLNROWFSLyW1NemMod+HUw
SD7kK4DFgf//9xYlghEe2EOWAxrEcBFgj/6iBCjylXvMc0mFwhttS18Uzy/N8yja
TxMohAPG/7/0babseO+yI1OpI5Zu2sM6ZA5tQgkZNxixIpbuHix8oqoXOhII967S
rFAF4HKPMsWru4I9ncwFrQSMt3fH3WjOFpsRjPGEprpSBdGB5sfPwNz05/buy92m
jcUiCoorIKeSX+IkRbjRKy7gEuokH7myvY9i75+6euSV3nVnYOoV0iA45n471Ish
ZdA64UGjNsFtTbATmo7CbTws900xKbBy5EF4xBh/ljchAQK2dSMHVIoGsdOXZsEL
7vqGzq2DplX0nM0jRbqWZDle+V+LoqtBT6I62BcmdSNbsCDehmMj8WHuKrdAc23W
DIklTv8wPaNtSFUR5gzsuFJhdkWjmxXzeCynU8KqB288SM1zxeYs4x1i43oMGbDM
aPgalaXQUD7MHsdx3bRimTBQGZtHnTN/DbSdTqw6lYGikRdC+w355lCGwW3JYhwp
S1cm1/vAMeLEeEx5m3Hj6IFUcTNI88AsW73Umk5ecKeQKePKsyOqKaDSSup/DKWt
MZWlxPX/3xIq7qkFytY/e/36e05bPL5p+UAZTDEKRwnqeuwIycnKg9hJS4TmKzyN
836mNzHZlHGYergtQPk7/MH2MuqrCsyKIdYasPd9jk57/04mS7Fx2YIXDbvSYAc6
/Z/QoJGZoC/+TdiSxKWV3PQgQoobpYWGwqFyLYIOSPZpfB2JpovGDfyIHi9utlQF
K/kQYrybvjL9wBOklsja8qDmNBuxnx2DrxZfDcXolsRezwd+jyxkotTRceQOeV/S
OsFrJszrDDw20sBfWxo9C9wIW39dRCw2eDEM67JoPywkflI13uQagYWUyawTY4AJ
TpJra27sRR8O0ct/KvZgdpQkJS0MqXWGyjDYhcxH7C8aBTxeqJag5/j1bMxvVa0M
c2jJuHP3Nt1fy62Vl/hQ8IpbMXl/CwjGDCCv4uAJyVtkSSaSgL7dNMajdqtEuW5K
LKm2hWhGcAvXDzyypQhgpqOfIeZHQa/vkWQip2bSQv7ldRU79d5GNwHSiUzkc6/g
7fxzxbf1xJZKdcKrgzXCIB8XZ7iJOsnUrJ7eB6QfHl4MWKg4lrwSu5kRz/f7a4Xb
HoZE1QRtHpb/zYlIx7CiCclBCdDkEjLslcYpbuclV22lzlrsBN1oDDSVn+C6IJQI
BanXDGD8VN4jfvQ5Rt2SNSgWtXpTZYUvzWOmvdE12kNt0Vwl59rt5yC5O1wD/ju6
8yxC9R8LQ12ZW/2F9K1I6bZYKHMI5qhZt7grxDZPUrtmfG+CAJcgmP4DK+4YXwBM
7wpuKGFGUKpctt8suD1/NfMkGOEfL8d9BqUuol3tkt3VaZeGvfG3QlpGsdD17Lgl
ide60JORfMT3s9hqaSRF4m0FqLkIU/llaaZ/NCg4blONESJH/FEmd/8/dsb7ylbE
TzVdrsEl3jA+8fSP1GvY0qWw3B5NwymvijCr0XQ4tzKD9pjptc1+5fc+MptVLrv1
IUXwCB4o7d9a4dl0JsOnD/lh0RsyHDftZSijYC7hy4jljtaPVv5Q1EJVtRbODCdy
243zlQhkBvtDgBbozw+T8MMdRdk6KEM3YRPxPxZfWgfbDR0pMYOyEosD6oEFMiyo
vdWUdQbke7jnsHFzSEKGSGU6CN0MOldm3JXoKIi2f6/GhwxLY/sBuqnyKRXkOYWd
QgwwrX/xcKim5AYGBtUp562+5JLWieWl9Gi4pUs+DZlbUPKRYk10TlTg0KinOJm5
2bfgNzQKb9KGWJ3IZAlD2TOzVZ7x06HFHbr5U+gndZykT5TBhBEjX/qWMofJwbvZ
hEf4HssxYF9REmob6okxhWK2jyvi+PC5qPUcQA8Jj1I8vDmYly4XtP+mAtgWKGAE
EBX7nWQ6A6D6QwD0xW5/XhNOIc8/mlg46q5tgM8Hn/9GxA4aPGVmw3xlJwhkpFs7
RM/zxTJv3RxRdKyubOS4cgITEB5r/gHVoDeC5chUUgNaL+3MCGTIpP5rOq0dSD8g
/OZeRzNXRZ0zqYCP2OAE5h/N5lyxAEnwXgO4pePdjhVKtGwutgwQ2QHE8TQHHrnd
Xha4DryEbHPp0O+xNfB+E27V+MnXNuShI7EhKv8ryRhJZUSxyZ8eUwgXoxsO1Kkh
vP0UoKdqMwrVCl49V8kpBKvA3YNDTm4kI1nFPR5JdB3FrQHE3ARF+aYu/+G0MU8+
OieI4EnnucmffkjF9bFgtXIkyIURdm/G4q8FEma0bftQg0PVHQjfHo+wXqMZgs6k
JLicAO93V9mzspWrRdlMXuJtkeK8wT35Csem6q0fwUNneQ5pNHG2Fzh50CA7Eh3m
KvtZamGQp//8SmgliuwSt7PKgexO4e3hiECYLHAV5h4VdG40QufC7pDZZ49qHZiV
jPGurRhpxzGrbfjW0uDRl9oKnQZbrfb0ECh1gbqGrnsrOM2mL1U80wd/NlkleiPO
u5R8cdnHWUJmPpUGYDEG1NlQzXwuhC0eRuoMSxA8xgvbxvUSAufsxJXm6IzKWj55
rW4Lv2zI6AyYtT4BRfuHTEjENc+QT154V3TEe91xj9unuRAAXYdeuC4sMFMbwYkb
jE8tjGBKymuExnw4Mir40BCDmPbbCe8+RPQCjUQKX14PuO2xoSniqLb/0B9zi986
RGswBOXUo1Gg70Seaj0urnrnOxS8QI33/ZG9YkfoOP1FGt4h9OIG+0wET5igdF4w
igKvb1C96kN65mHl/IFSZ9hDvVbCxshZbdUlcagyunKBA/uCrtQlVNZud4NfLE/y
ECrHZgdQ2GQ+e5M7BqvZ3ZMr8YB+F5XeLmxG/6XMT0WkblN6Kc9rjSmiJB56EFuA
kmft+FiYIBePNAWVQAcvkBhxBAlE9E23Es0UJDZj8ehP5ZanyzvPyLc1itrSwh7R
x2riy4N6mwuyDDQwnnbX64x9Xf6M90Lf95L7HCDNtUvOW4qosnBUARZj8BJBBQuy
k/UE9XEtrbTPkFaPVqJduRhMRRRJhszJLk9WX3bzNOCSUNsFIL+9T+kHrW5jVfcH
YXN/64GAdNysl6FvX/Ga4u70iG2+O8H+fcrw0uCrZE3ej55IF87JZ7TAReFar9/A
QdPu5m3QSAmJ5VNfjABhZtg/HmDIXRdl3i9NXRnQYxwMsBjS09L+DBEcFDKFbPox
OgaEM7ErzbSAp/bLcx01nxOqIXX7b9PoBCsP2Z4rpegBu8k8qvrMJSKmVzh38aPx
Yuud5aEZTar8uSiofCiNcDOdKCdmYnNwS0jLx9xm02KF4Y8YnqiiIpQJYm+lG5Vn
liWTtoPLK0oH8kTGEaqgZxY/JrmhPNIicP9udkOUwD5IqOKvqs4FoJISEX/IoDdj
DM9SBueAExGJx++Sy/MjjDxC4wrPHx0eoLt2dcghyhuCi+s96UUQGEm6YJswQ6WN
4G6Vl8M3XAcybEgfwYoQ6/oUc6AjR8R78gah1dvGI9jX7ilSeitzKN5wxLBarAx7
MBbjKl9qR1oVSIHtoYxCkB4AQkw4LBToy+MySpb7US0JVlWrvwOUyONJXbxQyVdk
6SQ95bFZU6JFjMUEaZCnq5xF/nkIk4HAna6gTmn34WPjUQURV3lGVdsGt2abPmvG
abZg+PQlWm2CxeqwXMJ8WRHHcWRS1fHsd/jdIH13yp2V5r8mmeaqgQbRZnrHippA
VKC5l0n8n68JgLoQSCNAPxP1wTk8kVKHLWUEjvx2iGLbBquNFS89Qyx1mCSO/6IX
YeV/BCBsMYejy9z8PNlD3FRgrJdxXtna0QmzzMSNblkFMUGZmwKLx8lR5UpJC8YI
lE/ZeuT8T+W/1IVD60UFe2mgho9j9BjmfEffGBrWHrgXSRTnFxQm9aBRxddQfxfp
lL7O5FJQUHHiXSkYFd2PsEwBoK63P+1ony95m8XTNPhMKijvfxLy7ePD2WLjHBq9
1lCe1dDTKk8Qo45zE+pRTqouwO6vThXjx5XiqpUyrsQIZY/T9RlUKtjb10N3jc/P
dvpBqlz0XcTo6mX/uR4+YWuK+Qq3leDmue/xyqbI4FMqD5pwVFHo5r71DKrKCyJo
kZx8YQiqIEWlrSeL4gEjjqJeBMZEa0Htm8IB1wM2I7a3vg8ig29dE/DLhjtYHxdd
4cK8Lr2ftDM28+FVPt1Zg7to++JtR+30m52WS18JyX+4tOoIN4SbDupXudHc3eqU
ONh9FRXSwJRfn4uYw7KysHiD1l22pFQN9fzi2CkxHaAMLGIVJDPP4JWqtJjeZQRw
3Q22EjSU90/0EfQu/mqrTrcSy6OwVkvTY2zk1QwXyB3J0xq9Ava2ZT7xtmQTF5hk
BWMxmfr46NuzKSf5gi4Cc1FyskHokI4olw3WvTRKwAKQw7nB0Xj+mQNbIdepNGuA
9uo8iFm3egNDcpE5vOqtqPvnmZ8hFgz6TPEx/vRfO8yB3eCpNguHyK8+eMqZRizu
7VbpL+iMR6tqB5lqGB1spmmVJKYSB6zFOdoe5Vd/5SMcupvx3b3zMpjTEqAWFMPI
GxJjFh6y9dP30JED+pYeC6wQJMR3l7/JSpQQHps/x+KgjQQd9fG43/YfuH0iA0kn
c3RM/1/nDgOvhKmQlI8NVDUyokcsGGPvnAtgWV3KaFmT0nz0lD9a9Oz8uCTakRfi
2XlGhJS7qiEvDG1y8UIkN6ok0mWnZt4QS7HU+FWV2BbZGpyHl7b4b5lsUCMcV/KT
HEfz18bGZ5/FM+aQIwDgxXVTmcfFmrOQDeL/COE/Fuyx1SFIup8kgBsQQi2aZb/6
cornbnd6hQON3rk5jBJft+pAZuLe1UHuRU0KLgh8Gu6fEqXDTe/GvhZqD6Gr/sEc
lByC3VhRmGHnaM8fEhGNt+L0Ugk4ph2Y1X1X84AADgAmXwhyPOFjUPFU7rvFFo3U
ACUf51xc335bi76jnuCt20xCgGSGyK6eX0pZmkYDUs9wfjo48NLZlBbY7FmXVPnc
ccq99d7w5dZh6LgPDxejDOY66BgsPR5GdhkHbKf4KEsQwfGjCcHWqZTw7xsRhpM1
kVp7zEc2PWJz83uBa9af4CxBp5ja/VES3WFm0O0uYIdHFcOCNRxlc8Sk6rGbatyj
FRwcJdmxyu1cV6CqFOlnXZlxwOmo9FtzmjUiLucq2hXTgJl6vlY0NPY5XVCySlsc
HqN4wOQvzt6HxjH7weGLsmHe5WfKsqMXqKW0KWbY0PqH+aQeyX5k+NFqMUJDVqF9
QmDcBMsqB6ISvwZ/JEm+3E6AACwai2sDu3qv6jXZJc0jm2csI1obB3k2hccyAgz2
4sPSFOgWjrGUYDQDmE1AjHsAV4lTz/HQ+VS4RENXX1MPqyD7l73mHIBE/FFnWUkY
7WSY8X04lCqmZIBs4l04+vLeDAryM9TQfLC28hgXJ1SBHuRZDSdLFX6o0nmYkhB9
Pep9jQTu5uJClWvz6UN9F44Ydrmuh9MAsNBgJUZ4Qk7N01JnAL8pGrxWGY4wXspH
DSl88JODnuTmhgyX+iqqHXtluWoHvL79epga+rbxBTxRetddLW4QNfOcxA2Axln6
OIlqTUaa03P7XaU81OjXzi71nhxQx10DAz3PD9RLfBdPo3qWLHBCftM9A+gpOQAz
sfWUnq30N61ZYC7NEKrhSFT/BkYa0V49tBtNZmoJshwATlOXwWoKomvhWIApgqgi
/uxMN8Ry5w3rEaLFIS941BJji7cAmaYuO770kuV2/wlM400lXvLKdGEzaDsKs8HU
6msBHWqyH1TgaOuuOldpBRVeQrVakhavlBh3wiWw2Od5LDwWnAdUxKKtCP5pLjam
O9+VUi8/X2n5Cy4xDsODL/7VLFMmwJ7dydVkYd6XtHGUx6P3cyCgx3mb9lFNg0Vw
iLFYsIfwiIypT0g1QQQV7yHsulG1SCcd/zNJhM3RS352VU9TBd6bF54fPv1ey1Y6
Jn8NYJ1/Zmt5gK0Z6bzPQXNJpk4th2byzurwPev3F6weojXG4c0mYAtLR9zrJsUl
q9377QHqMOE8ZzNu7KKB+Trgb/r3sB9u6tXgK8yEgPxIEKu9Sk7bHyvg4LQAMDA9
MeSefyoQ2TFX+FekEkSP8GYh/kDQaADytJ+2QGyKL9k3RIAIQGjIiPCuheezTOVV
2K4dnZeSvZoTIYOK2nTPQGRiVVc+qjY44M4l2f9WeCwPrSHip3YF8RYe1FJTumah
FzHJc9yBAS5+qyUbdqd4H2WqnkwEAyW55+WSWftoVLnj5LN5xvedfLK6rKWsa96D
dZZ138172Q1wiXqUo7iPs9he6JzCIXNfYCf38xiu9kfzpoOEK9l304bk2ISLAB7G
FTXe2IusyYnqpulPOxW3LGOue5sVdy4kKZfo6fxDqruMzhQgs73ymzmS49owR3SC
tD58V/etTGOxew4SpLiwSrVUTXusokPilky8mpLUNqehtvtSaquMWiRQXuOjWwaQ
5a7BS3lZ/yv6T2tCmMsH0P1bgEy/hHHu7mLV2ASU8WF6r305dm8whI0Q30kbr/Py
9/1K4uIkZ8HVLlkqQqOrjEUP1ezPssCxFJLa8XB+G5AJ6VsJEDIBBHbD8iLSHJqT
NWhkLhTZ49f20AcePWSKaVt3zU9lfxA5H9P7j+qah2sWymW/bHQLN0L47eYBle54
LPtssm39Ax4Wg+g+/FWGtwzQStsUkDhDATTVhEFBniZKnfYfUL8cV0CTpWA/htb6
ezMDnMDKunnw+bh9GxBuxBo6BCrAQ+Vmn05xTGLlXx995Hl1OBAI2w4TQNBf98Jx
c2EqhhQ4x1zllb51v8Tx1Zg+p/KkILD/usypEWQpKngxa7gj7l0W4EQmPA0+evnN
5+FlDpJ2I+X4R/Tbka/UpbfwihrnD0zyamMsrI4bNhSMB+4gIZZfNlFz7GzPpPe3
+qqEtFR/3ttG7L42hzn7ir6GZsmo0y2PyrMVJ0I83HArrE7v50elb5RR/XAiQ5pe
VKIiu4PFvE08Dy5mWVZyHpUiG0YfcXfsW2ENIzrkkdsRjAiG3u+z+yUjAc39zbDA
WDwpW+D0kENK7VcAJEPOcs/PyALl5MXgp0HpAnb77bZ7d3cA57w8GNKZgaRFed/1
3fjOZEb37BHbM59Lib+vX+FIbLgcSJJjou0oPEUtxXgAF8yJhEWWxJ8yktYElNSv
j1+Zo1iYatsyDME2NDbPpwM8or+Lib2p9iY0+a2CcJCV1T9dQVTqXuyruFutjcJz
SKGt33jhGaPzAOMd48kaR/fALwrGsALTY5bnFi/d8C67FYzmob3V2gOMpx5Zwrva
EO/2fvgo3qR1CjgNINFZfjS/v0N76xl6tGdpKkWyWFIoQqBAm/i1R9EpTpUuZxaT
mNp3eeyZ3PovbfZSRgJBQumJ7ZG5n+mC/17t8jmEEm+4qHbM/IM1yvGfg8CSSqcW
h+q2UBdFY+WxrexThLIHiQ4byDXcTAQ3PUDcJCD1hqpC+QW+oWfjMtfJeQExXo04
rdenHyAT+w7OlHkHZ8XSfvySS4XKDS9xnUxpl6/nIddUHvmP748Z7DFozzAbIFg2
b3vFRIFL+HPEyLYpCTeYGak/NkK64VFhwAQhdjnfgy1bdK36g8VOg0GMNaf2k5F8
AK71ZYxF2G5OFXdAhW3FNSYPsWALDtr5ulP3oGoQCifMyEt1D/WbFdFxmvaAA+rY
9PP34bIz5/bGPmnoXcLq6yhSoHkTPVtjB0OYK7/pg2/7rGg+Gx0mjqhBHv9CLexH
70o8MjCIJZUv8e8ArgqFcaraIPc79HuHECGTxWJ4bFH/NtBaOCJ6bXxDdfP1MMS0
Yryb3wiswoHN/AozNLT2QKGjkbscGimVsWFg96gnGzpoBgon3C/NHlHLOB6WCSer
C14tegYK7tNEoOCtVFsDYmG7seqS8jahMmtzIVnKq8dCrkBZAfeYDu5r8GbAcCnJ
FNFVf7d+EN/0d+4yD3dbWw/O3/Xefi7wGtG+Z/aPcD1C4uEfQ9Akt8oE/3Q6fTE2
on5TAuUTBabgAEyK6Kexya3cEWvo1ZbmM5uvXHq5f1bxwog24H1Ok7c9arRL/Wk/
oZ8zkcAJtG9OfQZ8p20cJj9rz9XqTSPAzcfDri6fd4qw0WIi05j3ctmqTMXb2+F/
Gp6CVORw114PeaGNs+xreNNG8Rm4CxltkSoSKM9OR/rb8C//eZUOopr8YfdETAQ8
yuqaumJBQDHdotNF7JlqoNTSBLnLlay1LNecC1InTtskqHUdJtVlMejNsG8KMFHN
gHgE49roJlQtH7RFWI67RFeQjvdNTLB+NGo2hp2FlgX1Jnc4yFMcvhsaJNb2emaG
ycgSqtSD61G25WZuDZfchp9x+O2JW7AFim899rCNbipMoFxftGjqvS7OifdxK7lH
hVNAKXZAcKBfbRiqa2+GvsBmj5hz4toJuDxPSM0kjWSDNSGaUDzMVjnxBHyx3bZ7
8j7occM8escZmUxZJnreozD3aKwBnD3AsuLhfyWDyRiwOi6o687GRxkbK/OI7XZB
4odVEvVuKWDlETlm73Xv14JeAVMV/0bPFUwSWqecnfQoqPjhFjKZ0+culI+tqCb3
dXT3xNbxN6zwkUpdlgXCkJ91o1GA2DmZfLq/9suamvp/kUjOrxsRqmmuPybZR4sL
YbZacs/wNknU84K2BUUrJMUnxDJ9t8nkL6vH5xJ6eeeQ0q1VuriCAt7Y7qyKJTKP
WjO+i5G+aiOSWqYSUm7Ei/4p/PvTkEDH+QEqUV/bwahSlRUWrr4MIy9bff/EOJIs
gZ0svXg4vuBkZpzamyeKhoiWNZBdUBHxS6PmtLBwM/udcmBVT+m7M8xCS+BWepWf
z+oZrCB5/juJ0WuRG23drLhj59ECre8ZOfJnejl5NMAL8x4ac2aDyx0m8YApzWA0
+HMYhtW11sTJvj9VmTnLl4/YfRFT8g28GB7ReWJHDqTg8qTXp1b9Ua4LTDjo2sL3
s2U4yWXeQd1EGhqeoL5w9XGg5QcBeEzoFTJh48DtLHgs3+Lk80oubKYuUqinbOuy
GlfPkTiKSneeV8uOFXOWE0nMcK+uaDQym31yOhqvMBSwReUWUW4xkb9Dy9MNllPO
9UWcA7sIzcQYmhEcKgY0W0lQJOcjQZcndzYwzpMsm2R4Q8nh6fXcRvvfelgH0tSV
AZCrCxYjxeVDBeirM8c6/XoR0FOLHXt4+cqTpWzEVmBR1JC6yyBe8+6O+10zFr8q
+S0eQT4XTb/BX/GT5lKYDglUdaD8JNT8jUZn+xY68I2YfGbVq9piJBnTx9TbDK/6
aycq6o91cUSVZJ6mC+ghzdzq2bFPnU2L5RZGPWmDDlqgwwNZmSkHxVXFXhgf3SI+
9kOaxy1ePbRTQmcGjzTlnQIX51VGl16anZSB4F9vC2XJ40NNMgbrCOq5NyF3WPq6
mHtCZozyGORyaxYSl20Vvo5gWReqGci2QPcKJC1g2RycqQJ1Yza42O9/FrTYr+Mc
1DzfInSvbd4xFDpuHvLC8JJtIhQB23q61AGDsloFxuumQFJ8DhRJxtR+q5GZ2teD
tnYkmKlWPVkZkCJwGXExU/CJiuU1N6APdlQxNuZJZWRoSB+To/ZBSVJqsnY63/ja
H6rlkS0diYCuAKBZ2PwyU/XZwQn0UgIq3wIDSpuhaTjuk/6sfexaUvkgssis5KNc
EIV3bHiiiY4dUeFDs51NPhT5VIBQLa76B/tbsvZu2NqTtoJhUodOmp8NoPgpYdtn
B3C3P7t361LtXS+DmHyXWlKa+1bLLXDRCjtltd9XOmxvQycllz10VxefyP6hSAeR
OtPc81WswRcUYbEp21KaUwrsEK4oJYu6+Ya6T+NYpv42u8I0mIaNARk6tFHsZTg5
fubks8O98nQtGYOuC88fzH/lpZcELNPsnl26k85GKyUywhHjY/wBraVys7HFovqr
QENcrqLXwBM9sj5FlRept6edH1+rsVYmKHImdpsgewK+UFkE6o7X7SXXkT2sLmAF
qk9EJw9PggYthf+rliWhMvm02H9moZv/EGILN87shF7hlZhGcw8Zghcq/nJtb3sg
zKWduBMd5uJzgjammxATY/RF93iNyv1r8COA1x2dm6X2OyFz8E3BzsTukrmOw5wl
SBexW7+rIoga2Yefw7PFwozBA+i5Kv8vtycLU14L5YFlJf5+JqIuzqbJG3aR15EP
MY6X6PDCKVhiKhSiiDVe7fEGSeEmfQPY48+IzdIkO1LUJy3mTpxZvHwqGor7rTTr
6eaBwPbABodylEH2a+NbeOyKaeJPxoJR2yH5tlOc7+RVx6I1rEokAH4He2hBhydq
qn4y83xypej2PTfEFiV+Ag144y8xsm2p9UmooaLYbyOI7NDrxYjFWXpicGSabh22
VUPlCkcsSN96XTUW4UOvJaIeBBxoOcVi2leVPUGS/mP7cgEV/5Xs4crqk3EBz0Dx
WT3H/Pc3uR30Zu5vyiGEW7WRWsr0sdWs//MclwWLt2/hYQwkvU+x2uY/l3kOZ6AI
/IAiUg1buhz3GsX5U+Lpn58L2Cz3P++pbY14bj//zxNBTDiLJ0NU9cUb1OYSso4r
m3X87s15RbuBKlbJ76PFtHO3lv1nDTBnWUhgrUUbTRJcLt8MgNTU1/AibwSxaD61
X2jDVkKsdYjR32dLbrzc414hWmdqQtapd8+wUhTvSTFGNZCRnNAFdESzRUmpSBYK
4sHTKjkH3/fvk6Tm6g+RvrDH4DXFwxSkhZV2IoTbcSeqUV8/HU2fwT5KODePi/MU
kOZorZA16Uu8ui+5yI10SPMdSSkjgRfUQ1o/Wwkb4SjK2d1LtRWI0ml5uACMnda7
CVs6fOj1KX+PDtvMgDJW//wyiUGE2fwjh5qdcgc3vePhMIxh5tTXDAYrYk8C4rYT
jlu5PIQahPTSWEAdo7obxV5gTFz9VQBuojvF4l04EmuLFuQYMC2srRfKzwNvQMJU
xdkvBY+dKZgZpCgLWzeEqZyWEv6VEdxb+B6C8vg6y7mHJ6RUb10ll1LZuTSkFWYg
fQwwPmhoT8BJlaeLvPy458NCD/3WjPkIoScDRviyqd+G6eDH0DmOYqG2fiRLFfKF
t2NhP8rc0G4k+V3zfosM+3h7cc2Yxe0UJioFa9a+IcipUoerpiyZQvlejJxCXqhx
UHPFd81Dt9VL+B/ENZPj7FsKEhVf2yJPWCzGRdwLPl6v1l31SRVAml4qZsyrr1rb
Mrh3tQRKaHZJV+01LYqgVh7xnxflv41blnxzSCuRum59JGHxbhnE0OVXfZCdxOxC
lEIy8xl9i/NbQ2JrOiiicatPEy7NAwdMIzRcRrq5f9iuKoXmjukLE4wkLShT9BXR
lSB6pXxtstmXjJ7L4gfdAWNkLJU9+KJuxv+NlaBlw7XY/DEtnCd1UTjvG4+hS661
wecXl4QnVE1JIqj2WUhOTef/0r+R8UAo+vyzFX3VCMEV/lWdTgzjplxYlgyITZFs
3Gg3UAe/AS6cjbHt1NJ1rPt6zzYowJUi3GFPMg/pfLMBlql0zMS7Y05FfSj0DidP
2fw8WL6IAetbzM8w0iIyDgpzC7A8W9koPmGm2QUZpVBI+3CN+IrFhG7ZMo5Ui0Hm
vLo9Lh+Z+U8maGMTAX+Pe66RtzIVbgF37icAeDjiSzRIm+zidob4jLfGW7Aljtzq
JWFGJSRPVDslvnlX9WYw21x1rk9iXEGt+tb13ChFeGhVROxd64sbzQ6aIny4MWf0
VOWnzgmOtt3U3IiJObepNdxDSDRvc+JACQi70UhKnOdC6m+PssnZ7AcEHWeHJ+zV
1gSX/RhmqJLGN9WC0wy0TClfjb5ZFGHbW8nwWEHr5+7CcA+Js7BnEYBEDNqGmpTY
ASdQ9kO5u/IRIW4bl3SE9du0KvgT1Pn6QTiXTNVzf7Xt0oL5K0BHpDsIa26LHwrf
bC0VSd53LpVTKaIPhq2ozhpIJhK8cBJsYhpiQrHUU2PapGSD6DDRUmgMDXI/pXR2
cNRMxQhg41NWIbclGSv4WRjGjkQxX6Nt3TkCwn0rDZq9/Zd1rNdIOAFxFt80HDYe
r7/hXDZaQxXcPOT1lW1nzhHiNbNuuJGn38n89MgrpX5UnYwAjVUN8ptNnZaQTRM8
/dV4I2BAImqicIkFBJlt/xGztfk2qVjhAfiO56wFYrwEQBO4xGUg7OuS1gwZnyC3
mJQz6CYlCr/jkVKNIcKZSvmGl5YubcVcGeVlce5dOYtXRMIeMwIkUTJSqov9wIqD
qoSV6emsjeNO/qVK1hU2K9Xu/8nYhH74QnQlPYSmPEyxF1iRyUnx7snD5jOkhzet
vgFlknKuWGqHLcw4znWhTtZUCLGt6UnsVRRfr1oYbP2hyPsaN4Bz0oyPMo7y+wXz
PXJ+dODh8htLsDVXShgcOhWHL+kGRbjjokl5efWymVxAjEfAXom+bNWKdTtOebld
T3+GRODzAcL2lbkA5RIvlqal0ahX3l5J3XbYZhlBQwZ9INhOjy1RoD0h0j6M9OpZ
tICUS5JUvElOsmtvXYuFVmeHj2mu3mWJQ3PcjAFaSnJbZ+3lY+rVs9mXCD8IGsTT
lvRBBsx4KhmLkTgdYdQw+xzt6FRTL2XNncyOroD1RlUa66BHJyBgGgx3Jz26VmEW
k9WovZlxwcRV+i0/Bf/64SolADIkm/QYE1O4/t8PLGbNPyN9n9wTBDh9TOKUJLdJ
zgx55Sjrm7LcJKBB3juWudxi6FWiDE29Oi3UNW1Tbvvk+DaqagxYiDfAUMR89Oyk
dJZhf+4jGksc47Fjt4HUtEdL+G94e0mTIaUGRyatJgTXIFG0qeaeFoNdCSnos1C3
PC1MTHD5mHi7znNXmge6wV/vSlL/UnK8PQTKWrlV1H0Hc3mIfJ8HuvUt7BN2ArSH
Zo9aA5gLGJrtuZzKAM8E78PYfdJ9zTqFnJD9xFfEnTZ8oAxSeEhEmdfyL8Aqrtty
1ee6JOLTjEJXuSs4CfWwDG0GTUaD86ZU1XcdHf5NyccpUlHbJUFBXjcMfCBQexGG
2dtXFz6lrscydOfKZS/IiWP6hsx83gHfrRDdHNIehbTCfemZX8vmtRa3qhQxEU+l
UUyBUUzPvduQy/eOQawJHY2IvilRFlgi9hG0XjwBRpUvvBVDElRkUHaUA4nisR7F
sEmNhJAC5JLhOokrY0stsSFkRfWAeayfUgk6DaOES10sADUWVtqFOqmKNaSxxoJu
rgnFqpVVPsNy9CjE5rqRO7utG8XTNtVP8T6j2aNJbNY/BT7I6ieYk9h8RyKfla0l
36hb6nRjToY/M8iFvjKwm4jzg5SfGBPqADW7ds/P5dxuSL81tbbQ71MV7ANJBbzp
PZKjbX6RAEo1BS9QDbbjV4rak3YuHBBmbqJ34B/dyfDRbAM4C+mzHjYiZc21loFf
UYVJm4v8ZJzLiY4VWZMCdOk0vE5fGejlxCo+GzEN7Kbs34qFJV8AxcPhApbPQAh/
Ybunf/FbxFCt03BZgZtAYh4OcIkJlZKkyHzrLGpwrwYdq08oXjMBmXsonJBrlbGL
WAge4+Sg1WGt+nBiUtq73FuYXNMBNSrBtqQj8cOu55/bSKSrEwQaQq1ovKLaRcu8
Xc4oRmaxqXso054j2rZHro/KWYWE/4W+qaEEq1EZaocJZA0pdW783bh4EnZ3gh2h
60vo0+i1W8So6xrh+oJ81KY/SRJqYgKsUcCvFZYIf3xZQh36U87nfEzWZYTZ6bVx
yeLPdQb5YmX2ws3/WSdQD6BL24gR8r07z4e143yZOyMp8M+MzpBgeujNY3y0OaR+
l5y5zh3GGZXFUki9FQFEkJ0Kqjsw7LBI2E1nJRNbQgtdHdcdnUFA9b+NvCi6VZIp
ndHq7m+1+C+zhHwmrByVGXkmC+plJoq72M+bOb7OzS2DNWpxcMlMYDfo8QtCsXup
JVka5IqKVE2LWoZdfPAcIisoNqwuIsUBnVImUAQ//CR4dR6M6nbWIdbhnIfgJ3Fu
dyLkawxWB4DzEwCKucHjDNMeO2hZ5hnpWSxxIZOovJKvilHjIjH+sE7uKZDsFHUt
h5DvGbCm2VfGfqDpUAE8wx7wH0IpoOzd4Mce8npA8WG3JZqgH9HUzkBS00o163ah
4pPr7JwfVdVRZtGHE8sAAuT8/0ADISNpfEcz7FDGeIMUDHMS4c+u5Jso4/ipLF38
hatDylKC5INXxpNljRipCh1syGmzV1G2xBtSHjtPclBqLaU66snJ+iJDmBLVRHRc
I/eHJLh8AVGjNCUA2G9usH+OlZTiZn5WII9e5CpfYrkIdhyv822VE4I0T7rZZMnO
XnMOghmQUXwdJX+OWBJYzr5BH8dqWsrMqVDXoJ07gAblaky5sVpdGSix23Rb/ATl
svmA4Yl8s131GnNuSWOeu7Gan075pv+vzYMhL23QwZdY1RL1NnwTUKNVd+z5VxN7
1+Ex2fu2uxK2QhsJrq5o6hrKI4Ei7/16X9lXJQjkhvNUyZ4piPahBQhZqx3NJpfX
wQWf+FmC7DCU/JKBfk2Ga6QS4Xgyfso9gjXs96VeKV+jvMXTrPnzBfSjTju6fqP1
hNLEvelu3sFoCs/C0qfQWEGdeNeW3EROz83uI+tRcuHOXgQuOKnY7q7gMIuUpDFn
lULMT5TGvZY0fiu2Q3UEcar+TlLAHGSLu08cVr/WMsq9lX7TDp0gIIArxLkYxPoo
Jvt7ae07JHvfePWkJDIZq8BmBHL5bD/dwXV8bAJ9RStmubVcDnZD0cADXL9tpX7J
kbJUPO1PGQ5ZQPNq/6F4zmuiEyOccVB3DLdC9VG3YzG25lEqJeK5IHsCOGdpfI/Q
OrI8+t/YGjZ/BtuIhYjzT0VIqQOZLd4Ii8Td97wBWQmvnssieqEVhxkbaxnxN43f
0N3Qds3cvVmHaaxn8MRikQB+MC0WUH5MeOPwPG/Ev/0rO1zEfYRufNsYh/5eaLaY
BNWvzPq6jepgzsZPhzJ26eFsTW1H7UvxW7pTmOZdH2WztDcpuEMH+2jGZCAQ9vmp
SJvamjTLUHuQxW+syajR+LsUqZxBAz1cvyfxoEcmPIxSqWsoqwP5Gs3VSt6PXiJB
6E7KFjrPSgJMUvKogleX/+rM8eKn2a2BDrPIsVAFHbNaENlouSHBD59pVKPf4ua6
XeRj6P0TJhRkILtliicEm6FFAz4j4fLasNXLeHchV2Q9eu9IAy9kwdL6AMpT9Qhp
MmTmug4AtJNMXocI+GOdZdkCyfzJaa2SZtcYSnTGXteSfFID91JBgnQElt+eswxE
yaGWEXk0OJzpjr/S1pUczpwz0o3R1luuaQOhwXpaZPwIlczTxsaxMjFJjH+AhxcP
xnf09058l+G0toGMMFAF28+q/aloMv1wPqH91jJo0H6HsvhgqFC5Zq1qaWPMHWHe
Xmdxe1fmtulamfgBdXqUoPIm6E0wP7w3mkURGYVpDiIWJ99DagLWnrHGM1vjfSvc
YPqwxyLmKAK6zub9luhc7BfzejrwFXWLeUlDz2zWAFJWKkIMcoaonQPX13X7qloc
DCpqWvWtGxMtGN3CjLv72g+nrw7I8NHXDDchu84FF5Bxt+NR1fRMP6WAYxUDbnyz
89OshUQgznRP1KLEE05whecO6MLnfJ662/ZXUvZZztNROFnstpwkSyLVbaGblrT7
VXs+mNjbih7xN84uC09qix/eloTE8Hua3TZdTda9w85Hg2my7hnic8v463I38sB2
HpxsBaTuQsRBcuLrVbBfUdKja8wdBT2C1x5G7bQmEQJbd9NoiUOav6kFj4nwvR5g
CvCyAKH8zGj0cX3BWbJ6Y1iyMxqTAzIMVFVPa8XddyQBZXPCgVmLm2wtj3QkeD4g
OdhtdTFLDFuKNCFMHu79EmMtw9r6fBI1llm1JKOCBNRyx5Mi+zCXOzFAfwWUBgQm
AEQH/4mrkEo3H5hy4XHYqOkS2PXzisKTkoPl2NEo5GNMb6bRikFfrUVSh6aCYUW8
SMQT4SifSClWrO27F/aw75F3nTQ4LtA5Gpa9ntVCVNuu5bl8NVBXA7vKfh5Og8Fe
jsl3h5Kn3uCa1Fb03kQ1lzUzJLEhSmiyw+ilczwlZvDDBN25zK4mm3IWtPuFoC14
5yg5bHzvij13CAFwHWCqQuchvcz15D86eDWOg06UYYo3BXbouG0YNaJbTEZtSgFi
oZ9Sz2oRhKqp+DDzKJqvYMHhY3RNU269gj+/jZAYsAQDj+0kIW7K61vUPCPDSJaN
0GTreIo9IDvihaoTwjfXI/JmUQ+27HIahoPI8luF8yD3mJOa02bmPVWAmZ35O/Nn
5MFk2Ek2Av0qbHzrwXTCwMzhP833ZrydG5wM5RY8idg8vj8lkeVSKPdKiSupA2ki
+gP+9eSvLKS5VT5gOf3P5XBgkYWE7h+2YkJWX8Y/PHWBwggN361sdbnQmEzxPIjc
35tUauRtHGsW0wWAruxkc49krFE3ZE1UQ7xPs5C0QPD4KaIA0m8MrN0WEpkgMQMC
B75MpkMXqUyjCBTyoATuWKr6un6WTmu0APE22z2g9WfVZVrJP6QRySw8r/hjGrYB
gSudJ0NZXvVTMAONO+KIPcnepCxc/xrgUJWmSVommyDIhZKPjKTEtPHOPoCsgXO+
OwiPMy8NIRxUI5phFiGMFSsUro9Rchpk2Bx6pu1lVdfRjpn9tUbFKkg5uBW2j2H5
E2p18I+Qa7Ucy1UHfyiucgGPJSof+TUXYNzu8+WUf8oGhyy/ISaVsOIh6VE7plYW
869Hs9eu2d0bphHviMv6JJL27VVaJXXkvNH3hwtso3jTJOrV6B40BmSAeV2X4J+7
bibdhpIpSq72Xj8LfiZ0U5ewF3SaFz2DKuQ2m5qboSMelVh/fWIblUUGueqxH/RZ
ntn71rnldAzqvm7TI2+MCpaWYj70i+MI59NtNUXk+M49vOTD+NCpb70b7suN4+On
HHypreWpIgX52XJPYN7B7fnjmeknImvyKfNSIfUyMPAjzRr/gP90fnsqtwFUI8CE
23oeC1ESu5RKhH2V6Xdg31u5jWXFn+xabFq+XtXOj79M+ilSAHdGKCeHJkd11yF4
G/V/GLcwemMWZqR5RR/+986WUhmFYYZobxDgHZ/UYvTCwGOl78vvQfV3ANTAcmfa
Al3CsEcyi9/2JEdwH6ZbUr0CpJMRMvp8ZE0mA7J8V2Og/3GJqnDQW/vdxzhUbrPB
iuKBrSVRfv74BQz9/FBZlBr+n+AUyxlpbTJcqmcDKLX9RyuGXQYHcPn9mm4Ln/uN
JZAGrus+k9sZ6aWM15PhKRQVEIAlYap/CVOZwgmGLcb+Lav9Tc0i02c4jGZOhE2z
+Vmm4AT7jpZw7ITe2XrzLOgbLRMMiLoopVQVD4JFQb9bAfNgcK1UX/kRx3W+44jH
ZjhLtXONIPrfjk5hBh7oJmOE+pbKjHQVI+zFnWAt2SfZvwoWY3vROAhR8skJxT3h
gRSx+fJFKp6dDe/8MqFOBrKAMsSIEWELQPe9qRv74kunToj4kFkpVthpB7yvOURY
N1NrQTCY0G+wjpnwkwQVuviJjSqvLagZuNWulN1hExtoLkJvS6TbPl0TDn3lipKx
GQscP4lMZkgLIaHqBr4ep72pvQA4a0OMs4iheLUCei+Qwr7TKQ/dtdP2bu4z0LfP
8lyuYFzL9SteJqTK65nwhoc1IQJU/X8G3hnAnK9jG/X0cKAV1o9Di+VFNKHrkzdj
a6s+RkIcRF3KwqZ0P2H3FeUOMZfog3b8gVSLFcZ2WdLvD0UlfIhoJNElHd8IYOg5
ACa7KkPUHgylpj4OrtWRtuc2sjbCafjASFTxTwYaXWav/giOlRsXk42KwLGMSJW7
FTx0fJ8gruHmJ1A3DgJ47VBJoyCpOhb/pRFP42wf/cXDieMa3/u4gCswMWIJMWPf
b3CfXvUWVLdAl95p4JjOfku3uwdqyMo2angm4d71gsDfgVZfw2L1PEENchf18/o+
C/rt+2zMVfK1srO91x/XRT/MS0c7Xor8vBHtuEsuqSD8SEfF/XhnOcA4M1Ge0k5E
IlkIgxvr1nDaiAu/HyYUdnOUtGg3B/2Y6MFfWB8gFncLYvrVORTmPKb0en5KTqQf
m621WcHsPzenGJCma0Jj0BbeToMPFyT8aXTKoe1VQVzBwx9RmpyKyPI6ySmQEVbo
QP8tH7QqjCwFORCBruQL7M8VZBPsLPxSrC9TrCG/3/7VKxXBfzjDbg4zDNNAsbmD
dKM+8++P/Zz02pO3ChWHol//6LgJw7EnvZogSENltuFezbaOLmJ1MRgIB36/29x/
TXxtlI1eoi7/vWOPCcfVZmKGmp/satJZcK5Z+3tFInz3qQN+W9xQiVs2TcDy6mw4
B6W3TeMzzxTP8yPnhX1RIZ5oZO+qXcwbdNj6cFlv5IjK2Jj52i/lFY9kvxP50nYa
43Ij9TZ7bkxvadKVWnyTatI9OBY35dWBcy68inqAxQx9rzS91bqNOZYhEWzOtFc1
2I6GLtjyapWPd7t/PKRftWCT9ARxrkq/XIBEIUW+yafmLc/AL42xEGRNVhiUzpWg
SIZfMHXq/MPHo3/qp4GELIAngke4WFtCs6Pg3brp9BYVjeyMiuiFlQjw9tuXjzBK
r1AuobpLNamrphWvngqz24cXafyovkXeNHnuMwxf1OXMPuo9FfdsXYK+jl8iwjvN
KBdyGLQ7cfTN2vnHLSXOMOzw+aC9wFK3ouKBStils9Neo2WjG9L4xpDUrsh0YRKF
ZTCKuVCEnNv+BB6P7LSG4zauwniWEyux/IP6ZtTwQCR+ZQgjEBQOW9B1FjMG8BQm
l28mwx/hRCEvw97aKJCTelINGWiOtdldAqm+hxDIO4DgHGuM3sj2h/nCdX0Kebag
FHotDvpiCXVVjjvI6h3C8itF0gxnsxVLQTWwT8yIOPxWwyMH1IrPG8cRen4ZXs5b
7+kNCHQcRukWohcKOue//c452OFfuzAfF4Wbj/1P5su4XciotykOOIhFRZjEfU7C
lKqqPCOZ5loo8UcMoL5Z1vq/R2wlZIrR3Y6MtucuYeHu6CHfWYDDZxAoEdxBAbBK
OmA04X5SsqYTcLEOcztyj9/WtX+LBw8vBwdKkq7RXLnM04O33a92pg+Ajs3AVnX7
ZKN1Sx71yfgUHgtNugSOSmNgkbNTki5QGvijjMIPR9BXAzxmxMRaQW56QOzCvUTu
qLBWvrfKr97QjN54vNYgXF+zRFCd+BSG23oYzJXdG40IbKtDg0VjcvhyhADbF9lj
Q1nkC9y4y17sU5VugnTcnzAd2v8jyoUbB2qVVO0iisYS9awUvSS0eAK4g2ljNvRI
8UIR8ur0s5ibNdxVCmbNidmsO1LxlmcC9vGcxL+9g+yI5g16OlPuzUyJVzjsI8Me
jOouefglgItcYsICTwfp0P2a1iK7ha5JWotgMA+DKIDJlFD5HhJsMIsOIZ6vs3qL
exPY3+svNlV0YwDU0HNtw0lIp6APGESXI3KOh0Wpqk1/pTsno4PnxZhhD11cZ9e5
0MBGflnG92m8qg9Q06ji4KzbxqyNDWwiZMDKs5kpd3NdsvmK8aFHyM+9UifcdrT0
RZb8GkKk0iGMpAghLcTj2uos0/iKhwd/b9+JAeHNiqhXidqARDcn2EP0SmrBhqao
B37fhkdXuARVv7H4IDO19LCrPMDDtSgxhOJTDoVuOmHf96E29P6f49fNNxIjGbRY
5O4j0uHDs3JzPhSz20W4SnEwBKKFe1/Ptq/OkgqR9m1x00baAedYY/KBV8xk8ql6
mdeFod5xoytmafZJsQAIOldft1j9vHxScvkF5x9FHKaJlC0lPzGB9b80YdZfDvNy
m9PmfSDaStVz3nDrqwR5dJcEOWdpPV874X95xZHAOWh/vXKC2GHxoW3vES2vNUez
rXENzpZfeRLsxzDmzdq7eiX39he7O4+ZoCaDcFJZmTcf2u0kSzz11OANy60UNcmT
5nYKWch7oYNu3mw1l38tGZx9oLI8LmxBaXOYQfeEq3wHJSLYrmvWxTYVx86p4UZr
jBMRu1NQJRbKhrKbzrTTD31CcziRV+T8s0WiAmjqlhhvokhEqKANypw2tIm8FgNW
i/udBfpSFMZEhn/54n9AZP2xrdANsoYP6r6LKus90uvoLsveb/YaiT4SSdmkCGMm
8t5a2hxFM9KhWsiFVzfwZlfHoe0n3D4BDBTUPxHdako8+9g9KenFGwPwl3TrxhXC
GgaXJg82uu7AqjJH3qiWkHVyg2FbUUyoGwtwvfQCgbo2uYjryouxhQmBRGwnGbPS
0EbN7Y1oYOcZ4ew0L+NMKyMcV+aqaI7uw0LdX659Fz/O1GOZHF71yfIpwfAnPuqT
DAg3RwLsu7spWPfGarztsm+vqa3YwJJeLZiWXpc6/seM1QTFtxIBtxmn+T4MBAB7
g++JfjzygDKdGLEgykFsq2MNr5WQoefzqLTSDoXpuIUeNQs7WEYhFfMZebzV8Ptj
tHF6zfk0wJHufNWzyt463ydaYNbFrhWFdFCnkeh76Rds2RSEocGjc+MFm0vF6qR7
TWSbwb7DB6sptjW+6iYus1TTMbVGuL0eGhW0uHlgess44ueLzpV56CxOmkWyhU0M
gX1zSCZOH105vXz8F4pJFjBC1s2NwqWZwDCFaq7icQVVxXsxof3WzZ24+WXA4gwz
9pHSfpIi2gR9dghzzkDs3TPLTA1MSNyFAO5RyDYLRwBOVyvfvHRsFfMS/YhVkaxU
BsjrnBrgt03yoKnwzD2XB+7zSM0rlX0uVN5nrlMnSFZ3WgHKbcAY3wRsVEj/25NK
ooU/v5TkZ+PcR9ng+ARL4+U6SWpGXznkVF/ff2H84H9W22X/Qp9lXGNKIOp5xmUt
NsbzNf6qKbitLA0Jzw/aH/rRJu/5012qfwt8ZVRWvoOb0oANYqpy3Z88efCqKDH8
AFqRMn9D30Z6n6kB5xg83eMcDn4hsOpe9TFioP3vT6Iafmcrl56ZxIaSqLx+B9mF
GMhTH1IYFUuwKDqjP3g2VQMiSROm5tdS7E5iesje0P4h3BKJGaA6M2JCUeFgwurZ
0VsJjTCkpAZwRp1PDousFGrRLwS0VgRsBgGTQzlfqVfMjHbxSlRZyZpDjRUKYYM2
5gejfTBjYT5/iNgXPoqSfACvhOHP16PghrAfIhPvQSwDfwPOfJnIc/McWhsoSG25
z5zNQzK6dH7EkVgtKx9pchF2jTNArHG8oYy0WnFldUjXi39PiSn+fAQF98zsoXxi
wqYlgSEnnm9rvqd61kIXcSGcNRvmYe3AO9Fq8ItrqyZPUOlcSQ1QNuX7yEbZd+gQ
pzDH+yIqwhWIIQGwaEZLkxXjSei3GA7sbe9qqSsbdkZQ5Bo5LE9BUnAMr2ye2WsB
3mc/nDU9T89UGO+hs91YjBjeF95U413ieqX+AW6rK51qeVTJx1FJ6RSL8ASs5gfF
19kDO/mpJnwDfycPuPZ4BrqXW2d6OjaKbM/3vsdjTOjQsD5YU8IV1JDAUNBkO5cV
1koSyOPpTcZoDBcCE73WfUYafNKIaz28tor9BBg5Kwbs16BSbRKl2wRzCqva1XWk
TF2Sl5aV6Durdv+sF9sKpiRlYl5hVE5/A5OCmgBah6lY3wJ3/a5+pqRQJ3+qf9fw
OrjUPfKT87fllNywePasDtJ1yYbc8Wh41KPBHdlv64i6QbJkFtVfektPgKbyzHbK
VRckkkO4UiFMxo7EQxQfy1p+GFo8CTalLzdRfrQq4KK+5S9h/H/um48i/kIbqClq
Ej8qORE7aEAFT/urIQs9Q4tBjlFvm2Ox+YD/hdPT4WjdeZasHSGI3u0Oej8HFVgE
eL77h6tfADYoVtBO1+hz/NkMVB1QRe7ta5NCpb+vZzFLF5NkfhiD4NldhQIsVBdR
lKlaPMUzGLZQZncypbaLpM9qe220zPy3p2PFDtxw2/5ynZ87/b4aJ32Bnnf1oKvb
kw7poyA7o1Cf1MFBSYI0Sf/MQXmAbGK8fgkhLS7FcCfljJDcOartO9Kaw2IAcfBK
Ou8XaeX2S1+CD4YPHFByZmsxhN8oZBr4KiF/02cjq2UBZ/2ABRBvJmVL2/QuW/T+
cOMKVmHzSGnvq8DGZpp1erhmWWwE7Iw1j5brwWOm3+O/qRQRHnIkRvd8L143ImNb
uW29n3I6vBQ2lB+R75ZFbt3Ommomloj1Tk0jYlojb08NxPMKBK73234rljnSbh3S
OBVyw20ldlr+xe5b6vE5ypXZctfl33Bh6HJrHa2ICYbbXK3H+LKejQjh0hjY343b
oLEKZtV723EYX7MaD1aOQzExykORmR/2EUg6JMEFUDBWzCDgEyzWnEC6seIgvTp/
3YEZrrqnrXYCzK/DW9aENoJGrC7dGJhokHOdcnyBVVXA2W507DN9GQ4QhntgCWZk
4LVrkuRCDCF4SK++ip7BKZ1o7oaHMhoqML19lbBFAVh/eGZJPs812fVECDZlnwPo
ano33//CWfcE5tVxpbjUv5GihS1h6O3TUyYX5gsPBQ2NEOd0+GH8YFAGG+bKJsR/
brY1piezDWATsWZsHIqPDsPco3GD8ikMsbQZFgooFbu+AnXRA30TShzkucnKt33H
i0TvKmXRESJ0n8dl0tGscewL1ryN3YstOGRGFJ5K9aTfAJwNj09FwCUcYGV0dCqU
pU3JbSGCNQS+wOerhFPOLNyZdpHQj9VnE0e2y5pPHswCT4IQufKWRZYB69kqwqMn
6ZsXacCGqaLK3s8fNYGaoReMpnNnHBKnAdj42ltKH/sQI0H7CbfcohJmo7pCMSOT
LIOuErej7iaR4BhtLJGKl8hRba+63WPBDQM1wMf2f8RTkES9URjKIDP+MOs6ZUSK
eLd65o9/kcCYc6BJ3qd27CsrA88Yo9C2COZQoKr4n8GUambsofuswMbs+v9oqhy5
BlFezBPOSTXfHSv3nodgPYl5m6UBhAfZGJpWDeiawXZcUYnvWPob8ZdUV92rFKuJ
aOMxXZy7+rNtxjSMZnR7CvXGqTmawS4sPJtg9w2o+xPOkVqyGqzNhx9qhB7P8upt
el2YGPN56UsG15pxKiozFcuT0/T8VJuBfe6r+z4TVeTV1gXrrwr2Gvqloh0rkAFr
C4AabKFb8gcLsOHgzNzuJ8r/kYn7RGGJJvGmA3yiy+UEhdAUrjiiPzjwPKJYCisI
7Cv6Qex6IKwxbfzevP2k3FVAQYmKrGIG0FZxNv39F6+MITRJg96UtjNjL8HvTalg
huVUs58K3hiP+O3WkLJjDvpqRgqPd/jnSQI3k+Z5fOcn/IWkxT6JyjkhaUs7rqz6
g616sp8s5lFpDpozfK+QmlJmUgAIt9uDlssXq8JTfE00KSVMnHf0foTqffzyBQCW
HMxqDxgQxfObUE09DcfU1LPf920lbEuTi/4gz5/azC/7i0XdGtWLyDDh5XlRRwV7
7AsHa5sPCwv/Kqh+69Us2Z70RFgXYZqD4taVzr2HDNrI2zqBk+PBoHZFrnjx4UKt
Ga3+Fyr0XGwIzC6Oq5lAlX49+lItxvxAkG4dly+epLQcYWrwe0kOR0VXfqUP2Tle
h7i66gsmx9dtiOozBOuvJq+/le36gXWzl5dlwrr2zdkbmWvjcgTKNVM2jlzG5vq5
wDhp0v8GQqFt03ExI9ilQTVSoiz1KfZetLJHjtDO5p7ei9tUptP9345Z0rO54vOf
ipDXF3g3GzpIiknpKMjMqauts9I+Wtxh4ghBJ8M/PzWG2la0llQsj1cjE/uGyt9t
gB6kHWgVb2E492ym6Kfp3D/mszhMHBvcZowwhUueYl8lSvsAv9IQFdvr1hFH/boe
cWT/JrF2GRF7gpzEf+L2M9MTCQuuN8jf3ij5YSBjhNRDaowGjgcH1d1cpMl60vM9
3dqCfUrQgMBcWK2eCQoNrs2bOl44hc4VDpcz1+Mi+/BbKRtwifPl15D2bryx68wO
hO91P/sCOMI51dx3f3esEcUKqJcj/9gb8TtbtWolvMpoEGIbcVlXz7K+/RI64or5
mpWTwYWt5PLMza2Gu4bcfHs5pyt7IXd/hhITKirytjZuewqQ/69eSiejh9yqG9by
LgUlCZz/KAwBdgI4jRiYTYVqprsnjgELDGblGHrm2Eljnkh9TYt9et/mezV1BalR
e6XfPX4nhXVssGWvmo4AcpNmfxAkD7TzbChEYHQWkuZX9tj3nUDX5levoXd+P0Bo
9ZoahOjOa19oUikASc9JjQEKfl6v+uc+1eWhhKAwlBYOnQPbNnkx6mF8merork4Y
VFCOnWMq5yjgmxpRsa2j698H7tAAKZVYUz16s+ZM9mYcoF/wEAbAJ6BOgQkqPyu+
t/J9AmKJlL0waZXZS4jOFR0Thq3Sd5GxQYK81c3FZ8Rua8nNI7kkq/GwTisItSWA
Zb+zC5qcvrTHok4aCD4y/drZvcBlVyUdLCjPbzb1VIgTtTZnrwNUNof62nkkkkBw
ozlJF7jsLdiSRGXbyRAbr3yXxQUtWybUa2RjdLYCmTABNJR6xw1uMFiOwQIP44Hr
UXutIQpIdoTK7E5jUBwWBTl5yIsrcHU0K43IULMbs0DwMHFt8gYGb8GsKmQIG+yt
/3xvNUlXy/FJbcN7duLnKCleksOq1OmetgTBlvFJg8Ki9ZxbQ9B/xHL22z0TUKSa
vXSqVo3GwGftQNe2pTU2mEhSLEjLh6FkE2K3YIqnpaxoko08w3OYOt0qbqYGXdIR
kZhzQbuvsqQs8r6jW6iQ7daaPaaD7IlBSMcHa+qI7yM6CtHA8ElENyrjvnYw1M5D
VQ3Pgitgcg6MS57vyjskMoC0rCsKBY/uv65SfvgSFVQPPhibkYXerQbPvHMa2qZz
T3KzAsU1gCpoz2nEqwUqRt1vZ0h6UgS0Vs95noKBN1o3Ss36LWXOzT9SznRd6Lkl
/0j2ZSicO/3IRjdNmFZmAlsATQsJzp5RrRmoNFt1dOqnjI2EBuiKKZ6RNfVab9pe
UUesZ/ixaREy2BHvjhAT0RPJqTmEP5UpMCENeVq0zQvMrmYxx4UALWr18rN3cRyf
UnGXbHmayiU6xi18aDSgw8RO4eDjxZRU14Ju7WN+6P2MOyYg8JicexjzBFfRpgOB
AqghM4MrJ9wP5lKiDGQdjLGu7+NCd6eXucxxBrqE7oA7GiiNq3Pq0wY8kCgVrCYJ
VL3GARbFWG3mRLFH/2W4HldCNkPpKSfsDSGOiPp4NRL9Yv2bwcRijctKhQA/AcBT
4n0YfmjnuWsU+yEvNGCLPvWYFWkIxEz5QBglTIkqk+DGxePfCUSp0SeUdOUErXct
sc/TC0QQV3O+Mzab6z3z5LuZf51ZvtrTuLg8OIGYf7XppbMMv9+/waPLDiXC4qZf
9bHSMzc+VUoXHhQ7ecaHVztYzOuFJlLY9cVdHrivXJ+5TgjEwujhvagVqfnzcg6c
cSdKrBGnRNtIdVd+zn2UTU57yydFp6vYBjZF2sCXl12gXsTRBawRCDeOWRPFsq0h
PJ40D0UB73Zwh5HeyLj/TcFfW5+Tm2A6hW9anJU7LW1MOngYsMbwNNxx4RjDDii4
hocxJMwZombJvTbNLy/AREWIF0n6MlC3exetHJ9mFj5qE9vSueGs6n4dZcr8gJEb
b8wCFnyHR6hIbPkfKY0PbPhjQqja/6NXTaqX4qRiiN9ai6viJmn4/CeGfHEsPRvS
dS2LNQyzTiswoQI9pIGK4NoRaKH6FXExxOQMCjVIacTkQ0xSj7ciCKD3BOcLJbIe
wBrqxrhY8JEUYUsLVoHB0af7vhsfrWMhEK5eaSvB4vR1Lol5lAoICY61HT6v6pDh
p5cXH0zfKY34E28hyNfQWydyFZACD7txP4KxI3W141ryeltb7MHXVkkxgnIcenpI
dXP1wsAwXTjp8W4zW1peuMcZRgRlpTvtS9KX/XMny2pwQYyWB9MdiGlKfRYmD7eI
M+sAqwPBzh22L7HbQ7zrSObhY85fakrsvXLNAoWw6rdMQ4SplxNXSB+jLFlQw84Z
bKn0brbQnxzPiqgE1uvz0JgxW5wueacijtJmxibIvNvZ1LGq0WMkVFLyO4Ehn2/A
Y/iYUsGyMfjAVHxW94mFsd1k7gAVEJpcexq+O4V5dpTDuVGbQwcQn1W0MwD4LZHh
ogywDwjUspxjEo7k9zkQ0iF+N5nWBSywmmsMx1VxO9z0/YCfVJY/7J2Cg00nNrFX
b1hYFZEhvEAki2i3GMYNLA6OjXZczKB9BbRbl42MPEuoir50511ZGlMUGzz/SIM6
2MXtjIxfAldADOb0ttVNe9f7R6QrK98oPXRfYILQbTpCKABuUoTKnauD0LZQnCRL
NB+2WxjZAMHlgzlBHZsKafkJ5SS5cqSneZILkx/3YMJXXDVHRK5Ep9hzCcrgJFQh
4/Xai0ZJq5+x1663Gw0QmKRNFgJNjC1V2hKibtNMJSJCVe3xLtQFiyLjVXlWlhi5
pSXyq2AT+hin3k1AYiqfE3QwdI+fzUm+6XF0BBgEfAusjLFaWNXPoZKt+9JwlmjB
FLCMk+blWj09ptRmk5JwBAbK3f4E/3bfS0a42M7bMhjcoSuGTnErm8HSkndVnPre
l/IDSbn6a8Q3rNjtFZXBMe85F0PDWPP600dQFzJhl1KcPfhN1eMJN4uSrmrxAqC0
lpwh98aw8j+dLhftM3IueZRwdIMJv4zv+1FqByi8XHAszfgDx1Z6rjbhwL1YjG2u
4VJAjZRPNHG28zKpaLst5T4OxuHQoLRGQxq//URv5zuzPRHrut1pPXHa3lyrvRND
LeVcXfJX3B4/bc4ENRgYd+rWvUpi4d8KroMpQ6hzEWfa1xw673pY7raFoODGwSx+
NcBMkXPEFjR6cBbRgFzwTE109ydKaEeLObWDLMqdCltASqB4k4ntPWpKxjAS8wBX
b1akRhM5JUnsKYokeMxrOph1J7ZplotWOYl2N8yXd1ncPmHutezs/0GOGHDCEczT
eLa4Di5mX67XeZih4aDwbqr/28/Y3vRbW9DMh8OI97XTFS6zCRw+Ksfcg76sl7zO
ghu3tJnWQ5g6W1O2P8qEHUlY/V5yLiRSvJ1uZfK/ELx85woCOO1NuMAF6s9snGac
OAi38ZZGr/ZYFCc9dZgyiimNrrL9x9lemXXkRAY3oIkLDvZam6ApO8YAGBRTzIaG
aU5KY2dke8y0NuxtKGEq4ukF/o9hHjDwgNY/Mc8w+hxeONuiqFQi2tUUBJO7KB3c
l/UIDdrJwtBFhorKFrAiyQzSEQJUJf0O7AJsqxpFsf8VuFSI0s22npsTkQiLyECF
v2s4+28Jx+UE1uGqGEItY5pWClXnaZ9WzOoQ5UfwcKjvwzbI3Vlz7V3sJwBEvI+y
kTZpZQ7z5khhYCbZ2pbTehAV6LijO0eTVf8xL9ra3i1NrGfEjREmDT7EmZtfzcn2
6SBzCAboqzqXzsfhyU17x/hPhMg0VQ5Z1+VlZAkJDvBN6TNT4Ve1dZceGVo7L6i5
8jaMyOWGhxFKhRVLNFRjtCCOHQifPx5NdU3Mry1WqFvZIIxVTihtGrBKsdaQvpvK
t9I1fikYN6DV5ZB8dUn13GzvKMnosCRbsOT7l9kCcd46Pn8q9gbYX3d/4SF2Hliu
94goEOSZDcXqFMvVKm2lidW2SxdzDh4bl2ocfte9VSd6buB5AD9nLAJ/LL2gChl7
IF/WjC+XTYuawAxHHoeJgX9ar/IFasAHW4Z3VM8BzttocA04xi5PWTgVhFOblh7C
rvrH2rfB9kE06z5R1HmgjqB4VTzqvfHIYwrJLADifOXONpfSo+IWekemTEZZYIO+
9lvPWtD/ihm0Jgn+XeS0g+tburWGVbo0HB2gitjVJpKuC9dCHMMe/e9pRYxlYz26
tAKiKjjeQMNNcXtWxUq4NwZKREq5dkaWCPpdGtJtYKXnGbJyVJnbONGmNrb3mNB+
9Ju6BPFxdXYy35Zq1AD1FxwUBygkrnbmfSL2H6fR4pR2HJtqimIFqBm9KFswBk+p
foxVeWSGX3koxHOaTVatRpmH8z8b+bNNvtXpA5CvN6sumXRK2pOTy95UpurrCPZy
HpTmVAdmScJFrDxDWgd7IhKl772Ao9pIXHPCoe//i4hv5foFQHOIU9C6saFFeeHV
bUSHQ3u4R9l8BU/4ILFTIgkZpXPlcIQlljMJDUTIe4y65Wkl2wJviQyWt3ja3rRV
KWAy3taeEuBuQ5AFeJFWsx2OGpv0wgN6ioqTmyYTVHdZmbw6F/nQLP1f29KRlpGz
rExc2J4zvvlNXCMXuoi6qiGwa2yguM+XM5FxgzqwIjFvj/bJX35mfn7+GYU1qNA8
iugSyQqb3CHviY1SWScMINyihgxu36doTJiMW8/fwfpDb5EJRxQ3SXyarSkJOyfM
i/PTFp+GYYDTQCTYwOCme6aCk2liFQxYuO/4q3zhlnYaif7pLKHzRI5Orq0BJFTh
n9qS7h1IWk6g384FApV8LsGbKEG/YYRI8CaDpTKUDBGVX396OvwgZT8E6hY8MIwr
D+GJyF0gtvHd+7bzKM3OZaHNuQCVj1+ARAkIqTSHGrOE27/QdTXnV4iNqPs4I9e0
qu/9LHmHxPIerWBFBbtRNmilV3v5yo7xPLOhufAeOyA7le2ULmMp73WH0fTeYatA
OKzvXfzPCSLh6nnxCnq2ClquhGqMF7d0QotyRNgtqtWvArRc/oAGqplLzKXkuG1N
tXanEd7ANz5f2rXcFfULb11pcgIPqKO5OZf5P6ch5JUlM7r4ny+UgDRNaWBwdQFb
9jEsF5hA3xaaPZzVnOmL6PvoLxER65gerNvP9wcrHKHKjljXT9vG8z97ABkH23NI
Iu/3nsm3gCgqUoD1K3kQnR1PZ4b6GcRPbZkimm/Rm0lwvc+XUbigPjlIDIvAukND
c+z4vUpiGdsBnNJmnS9fZPvshvMEBPrRTMpZ1zm11gQ6XlGe+SOBiPx0YMMq5mP5
SIHb08eVNEyRYWZvpkeWHLW4Abu8pTH3x6XDKrJO+0z8vVELeLaTXSY9ysrH9vLF
LaQTdW8LAfiMH0HUqeI6eCJjzMOmYrN3NwOdX9vq3PzU3JsAuaWiITsP0M3iQy0U
rXGjPW3m/f5Nz8LDXguFVVXlC4PKmtUP4Gm2CDUeHP2SQhNXkkj60QoauxMVounR
hK2WmMTod6gw9UO6AYNsK0E0PFUmt5NIJvdr108bzmlJV1m5VcJdyTYW9DnC5Wt4
eEt78W+wzy6kWENaKqsG7+cnnvlJvNJ4QzM8C5vpGndrk+T42hCRF+rwL13a+RN+
hngSZtAA4FktnHuJjYwIGFwABhadAfsjCJC97qKy7eicTvWsoV7UhSYU2U5TmwvP
dkQMnluZnIiMRvUYmYkiAkyj4CIv2qAXooOs0WQlKBKrxWQJwqZvBpK/xJ52jQSx
cIk1ty+zbExGq+HzuZk3V2Gema6O2xi1l7tIRjzmBaoazxY8U/DfB/O7uGxy4Hsy
KzyTogKCZGk6uW6IvLkOgpm8HUYQx3kPBG49I7ESPJq62A/F2Q+guXXq1+GUtukc
5306OcqLnG2D2xdXlvqTVSdhZgR72JuRbS1mIYWeIppH0C911AdMS81LeRaLsrxI
YQJfWCD3ojw4aIKn/LVVSARCacIYSSHL7kZpp74HYyUePOudZURECtdvmHbFaR7B
w8gh+S6v1HiB/tWXWCku+9G7D0Wbdhgl5CXelIfSzJohKlIGi1V4aysMrMsX6Hig
Gge1Jb2NBn7P5vFxZANVZF5dwNCaxS+EonXqn8IPffptYrvwoFCRJXuMO2xbooIM
j8KjtSZFLMbRecp2paCnRCvBufj5kRTYV6zWwlkrtzSv1W3bXfj5pNe2P6bmQr2Q
n+3itvvBuWkrxJYfOeGH7uA+PM9+ObnlJryo+U+MC7Te5bbhEEe1T79LXmbAUezI
bWRGtY86EJ6rSZ2FRT4vRtpNPEuE+epr42fBIkjMcioOKBOOjwsPnYF7AkPMtR+r
smrsvX0yy6PpBQZN0RjI9K1nIP1CMUSB0dx0V8Mo5u6MptirGNI6LDWNRvngA1sD
yfAAOZ5MCmlmuDC6W9bQXav+vCL78jC7THUb54Hwgbf1nMeWWnEIolSsQ8ngdm41
7X+ijMkeOGhCrsh8Hd2ENgStQxAEW2tlsCvAzRArR2bxdy4jYY6G0Um+nQUfNIaL
zhAMlMQAhoZhFInCr9gZp2JxiTw4cHpQhxKs5SvewPHG71TYp+aR8RE4lics/KCA
PtdkIOZQXD7LD+ZEeCCYF/PWRe6MtJxWCDCcQ8pp846vbdD58fFHlqRUiqBwdPeE
OgBa8ureYNL78GJl0UJpajniFWGGy0IajJ13vSlbFsBDEOxentKvt2Ht836cOTfq
GTPBW7Go/yNxnFse94aM+TMpB6RZ+qIVvss6UrKBuo8W0KnLudDxAimotMPi4ILM
D0zZeRJFOusjRHiVTmgik2vjtVnnkR7/pDMQZgLJQtGMQI3DbgXhlLHUBLZOxXSH
yCSPISqFpSyS1VUYOcZUUST9Qn2HUm7moCb6Cp+ww/1wnNEFb5rsSYFEdXXMcvjf
auanGWB1DVrGxQgDLH56MNs01s4TtyXcy70Ecdz4Z2TFtbFp2I3nkHW/RHEIyQxC
BvjshDkBQGAcvA5PSfNK05IvtXHB5azmTioEm0NRsjW4bAWSt6TFbe636H7BqaYO
4xJH/8ueG6bgWLGg7+k6kQCLWdqHS5REtu8/OPz2LPiXnkJcHi+uhpNzNsAjS8j+
e3d9EMEleain3WQXqDzcJSAPfHLqNYestHgmZr1VA3DcaKthAUzDNlNUtKrLD7GQ
06oH82/lDygz/YXl7blcz6/c4E69J4+9fXSqLVvGEPPzKD+c4Tgusp2gnHSBt4M9
r5kMJ+13HcgNuIkObZ35vQg6L/Jg3oovaNnTZFpt22IVTPeJsmz+ebeeX71PUPXS
vc7JVd+1NOZ5Sm3i5lvgGqXyBGV2HaC3T7svlzUSbQ47swk4E4+hf1lJ2CKi3cCZ
oiaJRNlJWM0P753bza1Dd6wlj53533SCUyoUrO4wSBb7TRP/v9+TY0LGH9TI686t
yM6jqE0EDl4q3sSRI3r0iCPuHtEK47TZQRNbJy5HPioeZ9yF06CxpvhO6xJ6R+hn
d7D2uieAQHS/quiPSxsyv5FDjroXkHN7Pgcu8kfc6Q7fIRMBu4Kpb0G9+5qwawST
p8BgQTLCXKi4zoYbrQbhSneTs8uRj59ugDUcRarqf78Z65ffJP0YzcZNHPdiRyy8
CHrazhgkKGVMBr6X7m6YYDfA4hTH3mFNSCEbqIaIGcp3FYyYKvHmieZp9WKcNqGF
RsbebhZ9dJhy0NP0cKZS7qFIqpv7v+IdfKpX4Q9e0rZjbiO+o/ql+r/xUmuBCvEA
A0ivlHy62QSFhgrJFivfyNU0rkCi9QlkOJ4YYLHNjQDU6/qM1zp4nh3MIyQ7HwXy
xGA0WvVQGlR1WhXlf1sZdixR+IL66vtJSVlmvu2q9I3JAAu4eCuP947TAO4OymZT
kNFvFC2Z0nTiVv57HfwiK2Tqmt9ULoL9vsTioQqS1o2/8mqt9j3yNFRpXo4Op1NL
qOwNTQtKb4tDx1kTHUyp6P9ADsnNeoHxp+yBoeEQyMyhaP3D16SXJmr6ufp4Zpq3
tCaKP1lhg1FZrPv/+Nf8BU6NNHacc9EEHYYsoWSomuu2vIVp1qioarnbVuNHpMC9
G3/TZFrUq7UionGv5b4qplMzX1MG+QLXIJb4mbU9zrUoe0gVIwMO4vCSUdkNjwdF
dMOsGXRKTEapzlyI6Ap5hhpWv9tdpfUl127LroXwCgfMUWFvlJPCjOn/FYWB4jgh
tlJwluCqs/e4FwR3UaGJDcCjJhkRwXmPCOoNu+5JMwLjLzWMHz0YUji6kuc1vOpl
SsMGKa6WjQZYq4aB8Xq40PVHBK4hKoEH5f42fhLSp7Mcewww41WVGCZiVjuzhE68
twf8qDdT+ZOguFYgroaXzxTAw/RLYMo77OqaxtQ5aw7Cac7gijryb5WoB9XrNtuj
esrSn4DT6XruxPS8cdokXxfskkvQFkJkCUPNR6jW9qNfzKQSQOj3bdwN89eEJJ9s
rQyFtexC5ytBniBMhiza99UcMmmzUU3SHzc6SdCeIAG51OKzJxfUlztbPJqx+hX0
aDqBwqzD/Zpkvu3sEoi5jnI9vZoTmQanE3+ZSuPQVWa0GQ0hwSDe/H9AXlBKOZFJ
NOxNl8dkUHLpj1vOms8AF3UIz5QiRvtLb2FfHj2Gxc6ukUf0BocRKPbk9yoWuBsW
p1qEJ+ljOMOXP/ak9kTPUBS/qWooiQrFwVHjUkgkgzYhJUycm/zwuBPkOaErmAAK
SqE5/xahXOb6pJpsj6IebqCvy2N9A5nZ4JKf4/Exv9Zu87QiX8pMH3u50s9prY9O
03GPCfG/zB7yYhR6Xl6ydqGg7s2k0sgRzH8EYr1OgswcFzt6Q9m1HX9jdLtOIAgx
qt1yOewGhqM5hTN+rDIjp33+fvLAtVv6AM079+fBbxsAC+Xvvf07zoOtWhBU4uBP
EASjJVqtLOpMCLoiD4+je8rtaOMbhoLj2koOV7JuLUbpCPpGWNKHHmSWMcPU6KLB
Ej2wjKmQJy+4Z24uPU5to4OlnLULaAHWHJJKX9tZCLYzoiN76D3RzoyOpttGzv0y
YUVz1hox+DAuN6AxSF0kyQOOoe//95dO7CrLAMTIYFymJS3EC7iqER8ky2l1sjGb
u+E1JduZZ0CA0r/iZpJDUpK8m7qpobAVFGByZCk3kVzSNeWAGOkwarTQQdMhBWkO
xAtsx0EcPQMTXZEbSr+V0mSXGCXBIMQI8wrTQIZCyMtdd5hj5Qp0GO7i/4keLqb7
s0ycu4lMQoSvSX6AjluBmnZWlKH6HxrHG/ymdyaRpSZeuURoZktvsSCKgZ0z5UpE
98Ln6jrIIheZzVuDik4sYZdyimCcvzJjK2B9zy4y6+ID+5z3cdh+0ncjpH/LFFLi
AtNoJIW7bMpVneAg3AE1h1mB9VQFpSpljkdXQ1soZUVVAjYspzhVymYB5mNvY9hq
7PajamCxkyQBGd2mJsazbTXy5J/F85Slqu1Z9SBYPWsXhTEUuaLZocXRxBPVN1uI
DU4wZyMRSPoHKwltiXFvrkFvINq1FKaswE12t5IbxsKF4k9onXjY21SxUwLZp7Q1
AXxJmH/QaZc1aUJ2Net4c/uOIYfPJIUXrKH8GAlrIdet+Z2ZVoc0Sfd+2orLaAe9
24OVvPp7CH8M96hkASqY2YR3POvJftbeeLlujFDgwTkAdZIzA/alPnb7hcgbD9T7
ueMrdVwgmw4eyGljv645ZZGOS5L0xob6BjVAvvpQQH+e7TtuNzyPJ5Fz9OJ9v0Cf
L93nezus1heop6DaPBZSVy6Es8FL224jdN+YN+LUTj4nH4w+oQfoQjctdhu9v7Hy
UMcq14+opI/9eBLaLaeJXqxo2AndvI5mbUQHSqMlqUwV/QhZQIRPleqAbwSbL/Es
84t9J0PXAB9EEwrBwgOa2qfti/F07mOQIU3VWoXHtkbnOQOBhcgOreBCUdVBYtOg
tRqjGpov1fF+jatPRUmenBrLFQpV/yX5RfLXYmtKkfdTewN5XxYYb3bv8ZiNvrKx
fCWUmUKStOXojCgPkqlSpXi7a/dMof7qhjqaYGJXbhuZ1eAZd07Vat7pwhSn4GZI
IdQlM6tH1cZn3Z4iznAydbbd5p594n1d89xNjvdLb6ggMhc/WwiIdbeFBXIYH9tg
/RwPBgpYedyrEOSdyUiqLpa37DXI9MkL3YpEwWbdLSiWEX38KoQKjwyPXwq6Hdnz
Z/BfGVGQY9jAUQk+3f0oIkQxmLj5y+kAPEjJhZVVxpML4/5fXnqSR5y9uN/X8sb0
PsENfwPdOmwXNa4idI/jsQY3CTllBwXcRSo5zUmfQgU9y97Dv7bEKFvwiw42+a5B
oMIXFBPX9HV3kmg/BWVD9h1wzP6R76+aqLDscl74U6od/KpYi3u/Opwlo0nl2KzO
qPLLKEnFCoH6nxzhw43V4SyJ5ZRm0fveLyk2PfPkcygA7tAdtYHSN0mh/x9I4uE+
rQ4vh0VpGNfpIp+u1V0GJhIDFLRFpG93ED/cNjbHbd9wmK0x2h1xjLkg0NGjLqVX
ZPmhO2ZXSNKi61OWtcy4qEwod3MH52UAGDrkUEg+Z6X96DRbOIQEXrEteHG05MvH
yuLCR9GTWVQCuWwqxZ2fUHK31z4m21H2OpgkEhZRBWJd3oY/IoWvPZ0sO3MlvukM
kgwnl8ownSwjI8yO8dmecZKt6PsQ2XuIfXyh22qNVqyDPUPo8cihnwDl4KeiWKP6
yIDvDnKgTs7g4nwEcux2a35sFZkQUzKMcCoj70OuSCYTBKEZwsQAM+6YFfiCUvv0
TyU+VKD80Ik0EfV0+ZAManSvF9U/Kc5vwhZsg7rUIEN/hbWYuVtjApdbzsHOqzXi
r4IcC9iPbaQPf6db9/upZANwgCPNzxLXJ6ks5WhPs3mXpUyFcvioKJlL7ZnE4EnY
EY1vTpARc35ok+nIB9+i62zrCeVL7QmMSgHwu0RJ0n6Ie2AIPdNrUbWNnb283vmX
rx5hlaFf1Hg912wR8te/9zN3+gwbKpl5TT4JeAoTN58+V3G1cE5sO9Hz7Ur9cFpk
hMt/4KP+ja+etBhlm4RHuilx29kYu8HK7JOrHQ84euP5FcfdrXgbJ2rfRP0/2PPy
ofTmUh7AMk80LlAaML94+om6jWtpZTmOkytBVRMq7BjiW/X3fkOE+CA+px/GKLsS
J1GQllXgcrk/QihxG7AKGQi44okD5y9w003PowVRTDi/3j81RjlmR+6PjpA1OYQb
uUQi1+d6BWxgs31V69odndC6zn9oBaBbPQrRra7amPCD7YlbIzurM/T4gyXYJDdx
nMZ7V9jXCoaNgI7xl6uHWCQBxp+/NGFuAvZRdlM+6pIViflr0sG/esfqK3PTrMxd
UAxEI+0AycKscmZh9PyzeeWIFZTti6/7qbc/1EC8drVodduE3Ea0H7w/R0GSi915
BQVgrpVTHbKA1qb/aVeIyvfsMCVhDqShUSqHqcNP6rjraS/cp+GgLZ2CIjg+H1om
BfGtoIf+WLBL8WcxeMGUbNMrHSMkmCpKSdV0xuRvQOTLETayIo+o02j3C1cj8Cu+
hdNFdUzFf2f3tbLidx3fzBxlpDXaQk9egJsNnCwW3HOaTDQ+uCH2sR6fysJH92KD
xxK+vC5yyqplw9T2CQP2bncHIqPRNDCWk3hBrcOvB1fsWxilhQkK/zRJtvhUQivV
6RWmgSJCtBh1SQJ4B+IGSLxVBUKOoxy2ChJd2F6GlmHFl6QkwKQ62JpSy77UxLCS
RNWNFex5gTId7Az8UFKLm9JJAC3DytAFCIwRW9L2sKjuusIxDa8tKxNhJcZFKztQ
jyh9zUP63XcRTa7jjdHC81lyneVJ2vzqMMCRklcGRJjz15QcMgeaU29q+Hygrv6k
inkTQrCQQ01cMJodlUk7ZvmM9lgXuB6NvFk9pC609R7RNeXPTN/zTEcCC0XcYwff
rnhGR82y/zuwgRvij22zKVeK01YmWR75EJo/Lh32eXry7k4+zSNyX+saQ51/vB2K
UlKHQSjWCYYOaahGtuGz8rBwajOCOoMjBflV4dYn7hLFxvjeyYsxShVtfLRs7amm
6xso8xJUkPjrcciyg0BQIDwZPUAlSxXPyJQ4sa3xPjTfI4MVxsVYKtGyKgM8MvYX
C5JUnzsSVznV/Ku4MLcfov5hVLNSCyPeaLLwNTUbbSEJB9Fy34QwhMl6VVebU9BC
uymq76V1O+aJ1S+DtDpqtAQ9CFzTCiO2Pv8riUwxKu1enl2cvzzeW59HYJ4ikRAq
+q7wzoAGJMBvxAQ0q3DEhpLDPV3VeB/+y2XV35K/Tto4PKhRjiMbjbN9CM28NGjZ
+tLn0FN2yDwpZ+To5WTJ736IqSCzfB/COB/fRlVVM3ignmrsNq59m0mP1vmS7Cbz
RoozaKJuN+LTnZsfIBZkV9nlN/ogEuvk+Rzk6x45TetLHsedlW6OkVWD5y7/6JJv
WiGBNetCN7WQ1cVKJjTaErl28Fnl68aLiLAMrG1jsrujIwOmoCiMBqgrLY27BnXv
zEklG2561NnKgFXkJ8rGR1Oy3tmZN0H5lZvYEkBNgGWT+NwSYiTmHORCp17DBREk
wVCmRGllmn6+mE5UjlrmMfs++QYn6RI5vD7utl2HdPV2wNyyFamMOkLvERXYXkxT
QwCAjPVDgzHAynGdJz023zx500ShYOQ1khH78bhBG82rARTy1hbw/CP76I4+T96u
msjbmqBT0+hcT+7AR4ZoOxRzXCIZSbLoXhq/pLKi+eFb8TKxjZQZbKWgitmfFPUi
QH20OUAhFge886RMJuU/nYbr245oeL+uR5IBCmwe6q3iEcoEbkVj5wFOD06EWcba
p+htLo3lfZ9A2IEbO2dxtgmeTeJpgriVmdgY8H2OC+veHnxYwrNVU5HInBiHKkEG
qjzJjL+/rAf4UJBKLoKplfZhUCjX85ekGDJN7vv9jNQA/TfN/Tzm67kd1/3nmwLP
RDN1CKQnV5TWDMbDLkxXhy5Lo0VWcNkkIGJ50fG6TvJDpJIOUTr5nbvp/jsc0vr4
NiQQ6UCPP8VSvU3B0FdrzVgLEGGAa+v2bRvKHiOw9plBUCipL8s5EQIZqRMCeK05
BCnp/cuEiaV6bND7SRLmJBqfgKoPE9/HFsTBW4TLLESK6mLk4BnuTaTu/Z9XrgmT
K1zAUBTViD2Zi9PIsLfCun8iDUo40XY/pidgS6AcR/T/UuT8Ic3dpjS83IHW8YCW
brMexmFsJBZumBJ4rOwYU2yPJ8pGfiqlgWqz0NJmtlRE0mnhkeLq9t/HxmuBTPVf
voo7shJDcPJBrmL0Nu/jGgQMJtjhsv92y0MSACQl7iA/rXz6Y0brUmcElHe8OQJP
obGnsFz8FxYhoRmhydjJcmIKKdq2Xl0f9ImPE/bQb12wHP/37A912Ih+e+M4k/+k
TcN6bKeHNTAS0V2rA0n2vuikuMS8oOaKNUL3Gh/+0ZR1k/SaDrdo/f6VAyeQOwio
DdtFsKKA0P5r+SKIJleLaEZ8SOYRvLQqirW4h5ImdoWRNFMCYbzhvIXa/XWMwUbH
zBngscmITIA612iJSgeNlXmcA47cdMx7L7TvD4gKAROOneonz1wYBCvQEvzThsDC
75iDQLlodLs1OBXCcXR1U7UusZ/5jekvkYayYZ4FP8dRNPC9av1tAlAC2GSbiYdi
FYBxJQwXwJYBbikDTBlMQJ5cP8Yk/ojRRANcoGbjIWmErPWDiFtxu6TB6yyqRNXg
W0GNUAPOl+bt3deBTQ6TATd1DTWVdUp7fhPXEzOo8zHQonw7lLDGV4boKQFLnfgQ
Y7/H+hw3OBnx8RghndHsqejZKoUKqiNSBA1ZjcZ87D20IiGl0l96w8tAyhXhrdNL
FNbosJW82MYuNxuYQCIbqacWZJ5iBfmxdDcFJwgFstE7itCl8MDPHX22FoAqpnU1
kTVaNgkUpk+nIngT7jOpWUHD4BP8GAbbfuS1N9Id4Qz9u9IhxoltODVtPiHdeA9W
tynCrtOBPIxtvkrYx5KEtBCUXGlk+S6BUKG1SukWL4kNNIBjgvBkYLQiOimF6SBK
dqt7nnvsvgDn6VMQVfB7Qfaqt9TLDbnwAZR8LcJJg/mw1VUZ/kM2Q/dtwwlwe5uc
mH+lr5O3Tfd2e5YTSsDAxchIj00pDzg6oVCSkNDXeRZf9XkmkvJqq2/UBJxKflSF
els6xI2u4DqMCqfsShxSh7mcsJWuIGuccwcugTj/4P+TZr6zPUJIJ6wtCeiVpQ3I
dBC1npQmsJ7S301UKRHngdwEL0u7Ab8fBN12A4lS2RoN84PUiTsTh5i4e4fV7HZM
2lt2rcfDxMrdUFsXU9Psc47lFzxGVhMi5RGPTc/3YrWIaAM7jqTBD6RkmR6pEFdz
DRJEehjLi0aUe/KS0fhwsd/BECL7XAbDoYs4DthAnymBT92yydmTHSVwjkT6qA39
tRu4wiRyAMUTNzFO8pLmD0l8vdMzeBm+3zJzqgYblPV9af+9/IypuJ3lQfWbS8e/
N51cVyOlQtBvzld+x5/NmwrTHG/LQyJJmz4gvVXQ8CMnv0meg1U7p+Oh/eTjP9WV
O7ZI3ZSKHRLFBhGYhUMUTEf1hQUOxWUf6ikZ37i9oLr0FM6ctALlBhNs3vzDpfzl
CzZP7I+UNiooSij8JzqlrBwKpP0QCqhXEDtQ2Fuv2sRqwpBZ0WbPR87jlbtM9lck
5kUGU5pGIEhMpXD2E/KO4twNx+aEEs6Jr2lzVM5LsCJbbQL26gXBkKCpeRXQQ/2d
u7kqNQx/pq0bULiJNunGEIJZ+b8QyAn+wHbHZcs+dpdn74H1px31Q0WZbRtOdWHi
AcOXBTNomTweMsPX6jJ/1V6Sm0/KJc0adk53OYWpXPYZrymuVJsEj//2Bu+IwKWZ
WHehpayG6rLd1086HlfHrQ3uJZBgwKuGx8Fy8SEJuMPPH7pJVjML+Q5W60UkA1SS
kWSxoOMP/WgBshdDjZ5kDclHCSVbljPS5onPh9c0cPlZfTb7nZ1NVqyajkEnXeuX
BBnrt4T0uBVZcADQElDaauy8ee+OYT9n52Tmzimz0IVUCbLgcV8PztiLc5deFVNC
Z60wg8uB/Ijuwa4XwdP3YVgpPvqQkAeQD4xAX1awd6LYRnRY2eMCt9lLTiMPOSiK
6Q2ZM9+oicIDva66KzRVfZjP6qjpvEUt1pbJqwI4P0ypLVN4rOreaBDJZ24k932o
JDePVUFISE+rBaxcP33X1MAcSkzHBozh73ofdo9HZ2dxhoeoX3IkYQvllHF2tgLQ
iDjZICf79ytJVKeHJ7qrzvD2F6EpG9OmhVFrBHVjqLqGUXTvEAHcKDcj/PILpnCD
h8dwHfz+b64TZiyQO2zhlegc30Er8VdK0hfem2h9aZqM3mMQgKC7FPf5zKdCPOW/
ql2Uvqi3rJVUiTXD66P4Ef08mEP72IupOHLa0Sd8MdHVmRAjzRnb7snanTfCKAwv
xQ65oYsry0SzkinkQcmXnC5WKnWbVxn9Zg0STFrhIlerTiIGg5fBjVT6Q273/7sf
jqtUGnYyCFPBA+kIP/FHe6qtbitVQvqOZFKum3jLmBS7Y1H8z/MXjof1PCixAGDi
v+FYaqA+CryHG+4abt9Do1rY0FR7pu5HCnu8cdRLM0dhHaR+6Pt+UyWJiO09YBuf
F2VMS5V704dSS3P1ldPq61AHGS0lOgrIHnu5ZbNiElfUVMcrd49EvhSknwgy+u8F
ILCwggvzstGqFfFQzdCTizrO4gZJIu8sIsfWQvmJLIXca03MxSk+WgxxDPBIzEwY
obVxgM+0++sSXyqPpqqYT/f+uq5eIMko2j0BO6evSOczbO9bWTmT665ys4oSzeBD
prmjZHZqJhN3SYenyk6jxLCMjU4wXCzDl+xvyv1dAwGEy5HKikBuTSepWgSMZcLh
oPXRZ0j88Z49uyAONDb07P2IqFXlgpK72kmYqtqSWPyjz+fDHroIiubh7ZMSTgry
4sK4R/noBU3HS8pjePJY4HUo11FHhfBLxJD/2N7QM/1l9+9/hehRTAU//+BP342N
x3PWMD1uefm1dlW9aFuSKH7f8jm46ENR/jm77MqnaUdl8W4XY1L6XWia2AdpU9o9
9aBz401ruNQN2OsLiYoB5LWQB3WEoNrBoYG11mddQduBlSOuA/SyBUh9DiVA5UZY
1qe+L5SU1SZdCH9WyxyTaiP1Ke0VQaKUU3cszPsUs3+BqE0db1y5c5PXqSc7Y6hv
Vhj2q6RjkfuwEs0+TQq8TicrwIYz8GbY6kDJoa81iaVZ9mHYO23Fe84nZ8ziAMtC
ZaXnqxoaZ0yuzxuqp0jT1S7Fi+iXfH+8mSOo4G7CupGR6mxjszWRFQp1AufivHfJ
P4O1z4BBvCvp6grDTR8TqBOhZ5+ippLiM0ePgDES28t3iUMBXNBgKtD0Zu52fLcu
XqNOZ0T6bNvGFg0y/wwK2PPCDGT2yZGE3mWPc19tiAHOjgF4SSwfYBPuuVOcZXha
qg3o7jRvHt99YiU5nDgZec1Bvd2XMRDx7Gk6WT33oNRfivp5I7SK7xXM2sKod1Xb
HrnQos+LcQyL+z8Otq7bB76eaQw/GqKEBLBN1lp5zZbEIIhmxTFp0Qy4/FmoXwRV
HOwNwaJKCIoEIkp8bJJPPLTBQZBGxKgfCY34dfkuwGI60Cq+p8N/odUU9YSWlfBj
k6mIZWo6oZ9lc0Dj960p2REWh6PpsVT6URseb/eRaZyT7egRi50rA3pAagcuVFEm
RYC9B4VRX7Zzx61fPpUm+/ePPxIIpWuduR+rckyprwGV1TJ4vIKovozaMsnfe7qo
gRmaU6ojq1YQmCODuSG3Pk7dTvgIno194zmnMqt6LMag76xklO7I4f4nyK1hlZy6
+RcCtajb3a2vIQ/WMtyui1ABo+5ZUeEBvOAocYFZw0s5YYZdtIJbtsuL8dNUkEjW
P4m5Rwj8c3hCcmXxVks3NLAe9jgNMvyKFiUQmPKEzqe9wFCUhgDCsDLT0t4dd6IB
b08Olqe1VixsyWoKfGlSVqPnzwOJkZO/4uau/58LUwX6/LQ187mMrLZfmbDw2eb+
hZea0VRHMrauhp+xNkGG28mUKZIzHKuM0h01LojPV715XDVVciXeQzc7XigKbzRI
6r4TYf6pwYttDhSl7Bj4YqcQHuI396+iyerhR4ni1IYR59V2WpVeRdmVuenQUDyn
laCBJOPFXSOnUd75QkJgi/WmcFUkRWjJXOeblHDFXHsUlHAA3wFcii1QWMV8c5s4
cWc5u2tVeOQw5zf85d/ezKGWBn+1DlyN0ekjNJnbNyslM4BlWqwT0oMDnQkimDbW
bHpi7eFIQTVDPrErja5sOLUev+l7DNONFR2ki3hxjl/qPxXpcktUwVgll6uKtAVr
+xqSHYQDlh6Q7eOn2N1uYFL2nsIoA96BEIv0x6cTqmI9hFU4YO8djOwwICvlJfdz
V9FPoMRyB1pU/18P3cuN2o4E+AAZiJNV1yybbna+fnRwgVpEQ8B47jlEDaUfFmVY
zULiOctLcA2jVnYRwTYbcJQbrlbgsBPwCmONjEOXjRimi/wHqq9p2TYSpPzCDCNl
41vU6Yynz3HzUvBz1+mEMJNN0hM+VDcxp5uucSl9NL0IiU0lkyaDj8069gLhr93y
9banoq7ZCSlonAmwphvV9DLRzV53TRSBaoASR+N0vWDEp8pPsA1paYUe2nUwIAZm
CtxnR6qXOi4auAqnSLjmTTlOdCXZ7q4uiWve+RyHTGdXh1nLTJAU64EUYhlrCa3Y
eX1z+X7bqOAHrh+4L/PSOoUy8/of6jOSd0MTOERw9E4D8ztr9nE98i5Uwgf3Yi//
3ylL5wtwiqcMm8koPsYOdjl9DusreepmC3UsMrTZ11upXMAyJkKQFlDewgeJJMPa
peDRbKq+qLS06ud91GtnCnbThXIauo1SW2pYcs/C55rl8ygXKwb7gBSkDMYfkgH8
NGzs0UdQyOlfURgsSV4ItWXmqm2l7tP3tEGHuwkOkRHcC7o57tS0lBthxEmMVYtz
zbSw3/0/IpWXZWMxcAUy5ecqeuWbkB/vTfX6PIg70J9xxgwbDTbpfULrKZZPMVLa
l9pqcTFjt+RryNFpujzdfIRGi4pNd1M4VxBbxLNcdv+cPvHeWZp51diUCN196EMJ
v96Ifl+BfGpg/wa+ozKWn91UhJoZiu3dNUD9Vl6J2F9RCd+xyfsfH2/JQ1UMCxxM
oqMXibu077PoCkzktd8Yx/mA6C+Aqn4xm7S8zE8I/E92LoC1uiGHTWX2sT9CgTvE
ZpTwaqG+qz14J3cT77ULtBVuAwUOhu91Sa0rn9EsUKNe7pe/fHuucFEtnS80Dfvh
N3TuY1TWLVjZL9WBPUGZFU1ZNKJzqiCYJxhnNInfKZqgA12+g1PQC4rcelhzP9Ds
ttBRzRm2t/FTL7ZV5h9eYe1k4JO7FxuGmf337MIU7XevMZronNJ6o3Ulym+/ghR9
Bzi48U3XJNJmoeRmEkwOjUhPsFSliJ9Hh95Ywcx7iTa1ZToPIZHejVBJcQvFBIyS
I0o2W95oJUFagQ4DX0VmRj73BqAo00FdG0VqW+fIJXtgJ3btcdA4vfGRZSZWnfjR
y1xrrq5B4TBtyD+8Hzqkvncz9XXmWqeblkCu+VXCaIsNl0WM7ZqkHeHKsW9DR/Hx
Wq3mBoHeEBujOmmxppVz6+GW96DExICGC0G1IQayyFBWhSvs49zb7pvlScjR33Ec
8vAQz/GKsV9I/KSs2h5HPYETXiVgKCdD3TMwMZyJW759kdCPFD/COhfASZ8jn0/3
39KXUPJuGTJ9aMIZSigAYSnLb0rvgLekOK0i0QjQFSzjqe/J9oKmXSM3XJcqQQxF
VsdpNmqLLNSlGd4XLaxLBhCGnIqK1d2iPXaET7RzTk4ukZ+PRDqK7ZDOjZNP0Nwm
HlGgyjNbuSHODE0m3Yz8vIJYFwlYCJegRLuQ9/lLW48GhvKPzAfzMIC65G5HvgNw
/n53shqBRhq2YsQfD7PmA775mxh+iOTrND6Sstww18Gye1UOeeCrvENq5Zn1HpkO
RDHRwhxEENmg0V4inZp/irBIwjWwVl6tm1TBZXNFUvYBaw743ov0nGYsqM+1TehR
5RyGEHXj0wXcdrEIpeazwmVJZccoNkvJN2Ip1tMw1NBWZn5wHozWkdWnAsjFofBN
Nxv9VqjWh4J8Lr9vqFd7H5NSNhavqqHs/CQ/xuTuxdOWRYafHlwRhlfxGhiFY8Bw
zlua7i+8QdRMWcwJn+N6AYmQzJcozHA+giugxqGAfMsBSruyv7qNdnxuBgM7fBRZ
TzUrj9U6L120M0829aekIZNCp6Mcv4gFKTZfrVBWq73jADX6zR2bMfAB56RJOM0o
fWPDZW/UeZuCVwObcEcG0dFqLV3its4vnb47TWy/4KlkWlZOAET2fmik06usPs52
g2GKl9EgRa7p0CK9kTmrZhBjlR4qvKsPdilH1zmAGCCmuImlvO1sQY0tcGS/gLaq
dfipzp+xEiiAeArwJlV3FhGEQQ94MKnup0/gY4yfHi/Q06eZPH6scAk8Fe7XFoh5
1nOXQxGWQb9oRcvU2iYv/9oblaMiFwlLLanXalKP/tFhYYelOFLxmfDWvAjm6jFp
7CltmRuNTOBY0q/nJY9PqNch/HGPY5FKhr85svZoF53uAwCYT3zdJqPoIcHK6qPy
v2rfzzj6DUboKP5Mh6wtJKOiReDKsACXC4xKlelmdns/TsMeD7E8vDzYiFael7jK
/XLsCm26cShfDdEIiWavQmT7YrcQlF1h/aIVbqrT6UYIOjqQ4QgoKEh8rK5oLxgi
VCmzPRKW+n9O0D+R5PrN97LTBTTQeiyHUtU6W/8x03uFSP1t2TMmzqJflQ+/PTME
SYYCeTem/uHHdQvG4s4Zn8DzEaUQ9qSSJ6SrhHj9hUfvBkCNczXRbdNaIYRUAxR6
G2J6yCc4eo5aE9wIrQwjmfSbI+eIuhrolk4hALpanFDUSQr4Lt36UsmyJnWaty2n
bTTRcbmrRyIxWd8JhJ+i4RIrHMj5VRgRdx9CHP3OzLAncD5jFFmbFam/BLcgbBbb
dCR92B2axwpiKLx0SjnaKBy4hIMNCTDm4FnPDGe+YUVhJjdcjMpwTN3Qrmv/QpWn
GXLQgvjpLyTtSpNyKuR+11pEm/XBsucPrkjuLvEB/9X9o/ARr/10NdU7WQC96HS9
3mhiXpaW6AjI/N3Z4bM8gH/ilulLyq4NrOnDolQaSjznLyputaGKvH8x+QGY/rhc
ET6zVJK/K4Ehk3tAZzH2DOm3iU5DaiULyVYqcKhEXITtGE5Re5rX85fp+mB+nK0H
2Gpg87DlZqM3GelTLII+bcF96BV0ts2olUkwum6hDpAC1Yyr+m8rTzp/Nv9OPJvN
HmU8JG+Vy2TbalCP/gxcum9DwgUldNFfGm0fM9kn4VlRW5IgHlJ5mb2w66tc/mrx
ED1UP9W+K2MFUxv9JxOsnCwH/b7F8pD3Xywlc8vOMiuPWn0tcG9pr6pKTXQNyt5S
70o2bzV8fc+hMtKmpLDPZwe+qOFMSXXpfbWXPspHLmUsfTtXv9JYqIzp2j1NrBT9
vuQy5t4Fij8iYjEA3wRcVtEAoj4YL7yy7UPLWJillHl2PVxT8AcMVi0AFbw67kYf
vPKSdbIfB7v5GQJrFgHJiMe7yOZhPV4RJixaaStiYiiboD/BGrnpMpa52Lh6QTUO
kEpdCu+bpV8HsnwfmA62bARKck39h/ZHFCb3GbIOTVCAN6l2EmPRHwOLWOz/IrVY
qhpwZb9ICDAJrAy4i7E2aA826uIS2yRRy0xc4UyCgcLrWCRWPsmQGXrhPay7ik11
PWYl56ALQNsuPd4AMfHiarRlWRe7QTrfyDFFq5WUa9svinpmUsVLKt3J4umhCskP
/z8a/7bOMUatFv82iuQ4tX5QPscjlEIhU1rrM6IXCAmNMN+rGM2wbmt43U1/MuN1
Ks7/Sf56Sk/IE86ntWOl+JqZoC0oqQ0OM7dis8lrZ1u9dgDwHtumReHPj7CpHi5h
gZSF4bJb/Q6ypKt+kKu26pQv7BOPjRws1osFVDtCv7UFZbBy2Yw7ix9BIkWo/w0G
bcG70JB6UBeJlgIc6hWCkaBwB4xEUdnMAi+Pmoy4Jfji/xzhnImusbHoppnu2UUn
gl1JrFRQBDlAYVv8gnd8U8XbvhpY8/EHEOUIU5WU0zc1nSzye8/vOxqYdxWvdEge
xwIHRnysDh+JpY0c6nOnapOZomu7Af4WODSz0Sj5yepLyaN5Xoi7f/TB6puga2By
kwbuJv5C6wgLlB2IASkX+JExjbzy+RF0dlMfif1chvv+l+NorCqI4odRA/dEtNPP
9IWC7wzYaVZ7WXezjZQM4eP+FMzsTNfMA6lgs5WEig3dF9jj5wkmakIbZvS/gZ7u
gNJDUTEQ86uagk9QeXGAAzxkT1Cg0O7Fgi5uP8buIzN7GBZFmJAN2R/Bj+wRU+Iq
8e95JtPV6sBjaJvcCVWXw24hiny5Qyj5YAezn7KhFFNuEqg1c/faUuJ0iUNb/Qot
g4VMbAxiQlO5erpQp+YmcrVlaTyilTehTKuspZSBdolRP7N1C0vJhUARtWjVxdUC
BtUl773JcpU4x/BVfaVYRuUI+pab7SdhN8K9Ww4qx34QfkJcxsClBvDA2J9oAzgp
ZB8av8+bbIuJIb1w+D7Dojo/ZjMYfP1uPr6V9mTGBFponLv5mP7T+BsUEWkLz/ak
tIxMTH6nKe+8J5JLdrlHYNKMjwfFVm3pDHxTTt4W7aVJ+OGGDDyolFaPsjhLQH/p
s+qlYllv4tmpcbKaZRvBJBIdTax4DyOg1CLE+c0jPHyVJa+bavqINb/l0zqfzaVx
VgajJM8bvIxHYn+N1AvzscUsQaNIPMsF9zkXcWKY4WcgtvkHZXsCDI34CHX1D5ai
vKYO4Lelwefi2YBmgaZqbF8fKEWk7laP0DLjw/2khAhlpnk1AkxxSG22cTk2LV9z
PYTZunXE/g3tMQ95mmQSW4tZkkRoPownUKbaI+PyUlG/2waeh7Elw1tQ0L4zv9ml
G16ddcClZC7wmqzS9f4EP3Ej638HVDRbCs3W1s1b20TZOTS9z7rLU2OWy5T4TdF7
tPQKMiyI2JYETLrwwA+pn5n0teiAsmiiVEu9KfT5tgTe7QMxYyxzC4iO5X26NyAI
gtoaPnCN6isgKXVygJYtSBM8s1LcLeTuSW0ptDCUNbCuyb6fSBPl3mjHrDxhiMPW
3jyiRtiMtRFjJZtvlFTABhAXGdR4Of6JuMKP6eMEW6WXcXvnrF4Im8LXR5kRjsAR
0IJDU/3H/9lihvNb2l/+aPDuF3vH8lqZGulOXzM2X3lrBTvPLXELjVdHenD77M04
qLkR8nOyXsqcub7PIzzzaJHXiBw6RsbfQ2ErIh7sV0/FG+66/R6LYAoSECigPaPC
XM+Y+XdZ9wKHBmAmtV7GRlAPAfE/AoIfF++JGNbGfHnkqsgLxmo55tfcwG6yo0Sq
Q3OCUQ+BD5WBsr+4b+AC2nwsWigpyHLUnDFT6exeWsuuYjCwq5hk/lMBkFVb3Xc1
+tK0o98ZXU9nK14NujOanVFeeTqISX7je9hkiHofsqVZD3vBhnMxjynpfT1iSk2E
DjBJ3YXJTayxdewKlDvWbIs3eCa0+P77wmFbVIeImN6elfp8Qgep16fCgJ9sw072
QOw5ldPW9TAz7hpDxNP6KtZ3YYuPXZVv597r4FfKujBnOamqvWNyqAuONjdKnVme
MP+TfICtJwnDxvdyOgCPc0HPkJi+qImmSYbW9IxLUFjuuGKGJ7JevFqJICzmSNTW
vRhZMlDY00kM1xjryrg12pE09xfHh3ctR0LsIf4s4+rzgv3IJn/6MXp4g5sf6zVs
iQ2z+CdwayHGeHShrVrfHiEUQ20FhqFG7NP/sH8oHoYpc6WWTcUmlDBnXfy8f5Rd
zCfroWEXJlR0JATORpn7xnMU1wYSfu441isjl8CCI9MOJOlVk32c6zGTROX5Ko0b
/GZUWZTopAVVAT2crTo/XARXOXqYzAkCRGlxU9mPEYC5mngyhZCKLHpXBEr56ADf
Xb+m5V+lOC5+L7wDImjV/ihrAGAaK9nLUIvNkfDbI/btRObjCkXCKagac/0OtHpS
FonLFb1RUZAwaEkoslPBElx924adssArK/5yvIQ07QupxbofVkvzeKb7028mEiVv
oz5g/itxcNsrwOmOxsXUc60S0WXc4tX4ZCTO2RAc4wuZ3ZJfKcWU3TWjVxbIxf44
rfe8H+XWpSGCzLOFxQaYQMci9FnR6AZwnCn/lDKCM9Ao53q/9w1Tbe62zjO5MxXD
jNmUselxgtJgmXEqN1YTrUigf0WHKVJLyasudoO4D9Cob1tYv/algPwPDacr1m86
7aXOL2WWpHAMLs+xJGBewLy7HeAReFmmiNharhaC6JHjcHm74AaTFyvBnsWbWrcm
e26yShBcb2X/vqZA3iMsbqvq1wSgHqDxXqgs/OSONtpNvPNB8hSq/iWs4nZXsjgp
y3DeL/xErEDfA4yfB4fiahgWyVAj14vj8902BKc5YJ9MlYAwFuMSULHbzb6kWbcU
zvW7TsGC1sImmLProFXDem5AK/b6XpyXtqBcyf4YZaV9P/Z6q6RQezgIrTWH2LdZ
zBpdiDK35MHfkq2xUR4KUwDDQrDAzR6hD9k1nMP6RSFfJhRbTJk2+mL7uHWpyQkj
bQ/5Rl4PbTBNiNT3kYzb4/9laCu7E8ykpgkm1k3i8uFcXBK0O/ocF09KFM29Nb5m
1RDN1F5dfcz7JNJyVUgHvrk8xhMxyQkVVSGEJTI3spoFmrHcqbKB+iFuRK8lTZqe
6nlLVxjrVB+AEoFUTDODs0BAM/uvUooYkn+f+xAS745pwaXb6NkoSymyj/ve5s4g
pZMTfXzFWpk65sHN4BgEaZhLLI7mOV3kld9WwGZwkOMdu2vB/0KJkIU1D/JqCYYS
kH73MfZOO41L0VOab1oLsgTFys/V1BBCCSDE6PvY4FR1FrR9nZAUkJ5Zawc8mnnk
uJ1x7sGNQJSYhzHBOnOljfS2CmV21/+Rg5fs93cQMC30YXhFuuEBQsnBfE3SFBP5
LjSAoiQF5ULC6Huf3Egpm5dkrWbBf0/tCasEmwFmhG4pXdYS15EmKPCjwyO9RnV8
gB9hGvtVvf2hcOc3qCYijMqJnDV5nb/ex9aEnviaRyz+dBzQ3RAT1s2dSfurxJaL
lTtKKkwhjr0WTxBopXpOJCZgJRBgxnUdFubDv5d1UzQqB7IKY79ef0KXXD08mW4W
ZNFpRf2jKaNyCbGM52v0GSPDyARiRlfafxytRtEQO2km+Ph45GhD1yOJNVlvV1rr
l6j5w13hpXjenEKpBAyeOM6cDt3Ya4Gj+34xSipqLyY82zYs7GY8un2S7r3P6pe3
RDVPIMcHFZ5b8XvWUro5jBNmpiVYlTgDYHMShTxa+pRXum0qvsqVg6dSumo/T+7u
oiNo1BgkjWhn5/o/cFXR6ZT7r2nXImuYoyygHwT4ZBwSEI+nVgeE9QkRi38vKE1E
ceZRRQasH2toAWZ9ZVe2D28BYJOuPZ7r4utz9c6jQfl2PVPBBKq4CYfSELXXzvp7
8xGoomQNL42n0IhqgvNhun3Y3ruwYlbWNFJvr3F35kNB3V9Gf3eCQvYH1w12kL2t
2mKoCbJgwaZTs1QSIAqljzaeIOWBc1QMrfpItvye3tn2ULOwxYw78VaPDyvIRozO
Fq+hnb3zQh14MP5P12NgTCYR9+IvNmmu8I9dEzIBpyLlTmHKkN7M3yVTOr20Ajbm
RxxSzDop4QWSQMrzqg5MgdjJ9nuBI6e7cwvQ57p3+HwkJFlB/+k+vA5zghFqjcaM
je2ouoZhVoohLDc6CqEBg5UzMZBaHphyPZ5vO++r/nL4dd3HaDx+IHwQXL85Dumt
WQtgVPGXSTJFjNjhxaQ6Q5Tdno0EM533PN+/cgEcV3nsfjZ2/FjmXpTDg5hGkSd5
Eaot6wJpiSpSYjmiFXWZhAg98Ib179YL+RQtwT1fatJfPr4g3bvRAWmOhiVWR0ep
O6gr8knplHoIE4nO/7eqG5h5e2jDEVCwPNKTPjmMvVkR741/s7gsJ9HFVMrXfviF
uxR7ZZaXV9YyVxk7FS1NKkAkeFuYH3DwZJb/lGeNlDT0Ogf+xQaVXwbUeds6XUSF
iHRq1C1Visfjb/D9bD8gpR+8K7mrLh8lqlOz4MTuKdLhsUEUpDDfCNja56OhzvT3
BtTXXB6C9ZiC+P7VQnFub4l8eLdIiSxW2OjJGvrimEy7N2AOUNtq+itz/t+2KzpA
bvkllRyEg9QD277QtkQpaQ0tPbxw6XXqSERoftHh58/sGJUrKyS6K3FrabQltFfZ
7rxb7RwQqrYf0mmKcisEnwY+ypbBNyrvTRc+e5shHQOBhNK7aBOXhgY/FvoQV6Wj
7QMkifuOmc0DunMcXqGN+HNR43YZJwaZ20kyzXZJZcBjrGQKr/DumUyvoguCWBmO
Vp68LLW8m+3AFe/riaZJgRjtvfUtmRT7DlXtX+3q0PLiYLMuWvjyyn/dLNq2ufwE
PnIYmIXyePm8saE23u1YAAaddvMSXCXTvt0z1KDYiUFqQohkxMq9NW4JR9f0mgyG
SNo7wJLidWXtCSw9YAgFPuLWqQZIg0JsUhhX0+LoprAE7QLrHjbmlH4rx5xobEWG
R4hpJSODKiOlUccY8WzQJ0egBiEmilR/OeqRCiP5Pcc/Wd6/iNKkzqoaSBBi+MHM
fXfsGXBkzT9r1P8KUzssAlYsJOQOFOxov0ceNrTN8iu+DyKZleQVeZ3JRZ5uyhRt
/Dg392P3B60O6CWWK0abOLipmSoJy8Z0XVRVjuaHPj0NSgq5KWE1M4R2a3NghbTj
tA+AUpo1F8h/QEeDwxZHzOQ4H2n24Iz12/A18dAm10wee379z3K0lG3VIipMwYdD
8zrGaWY7zGWqmdaLWdjUYN7jwH7YbpyeVTCqk6Ry9mTd/N5kU7JCp7lLft4FZ3hB
zVHooJxStt9nhctbcyBeV0wxuEdrQzwmrBFhMgXLagimLF59+ddw53k1PpKwvVtz
QRiC3K16NJnqrno1F13i1uSLvctIr3lgJq61yG5Qf98w5py8McW4WcW3O2PAFawe
noR5UykwfY5sXv63z83fPP31Mdkul+whFbQAR15fLtYvNeYnFyoTXudJDcg6DkDu
XUsBBb6xxDni+fqrLeLtP18aVyik41mqmB1qKJJa+bivxDVCPeP9cw/bd7WvpvOw
+RM7jaTNztayCmrfWtzCVRM6Is9XXnlle/Cp24zuer9aj7kTj9CQCyRm9kRPc4Ql
ZIoZH54ty7a9thGgiArfEG7ISo482GOWUFi+KpglpG/OhqcNf6PQ+bqZi5shD47z
pxb5qPWNJ7926UmJLohhdLI1R5RsHn2qb0SoCDwfiZa2N+r/Q71IuKbcSV9B+uuQ
90JjnD1HqXIscXtsuF6z2pqrhM1BpZnhueO4fdSANgZwFG2ZrPZ4ktElIj6jptxL
5fHeJj5EMxkQJqbaHYwRO4Gf/xLDN2Fv/gUIRzFPtaosazofzHmvC8ve2kTu0Scx
GkShMJW3bB3TDUvRpmJrWcLaZ3gADsPCJdJG5k7e5hHJiANzKqyqA+flXNQvDA/b
HPQd8VReQbDkm2nKQbPanShd/kI0sEiHcA5JzB3hAl6dzDEVaWeOhekFx/tIf9/u
NUCEh0AXS0Y8HWWNEU81OBkVf+KGCnIPxfRLOrW8Rkyhv3p9VvuGPTBvjMR4FepP
/AKPLoAfwSeTbmTrPV5SkOmozYLLUHbFBLNkNSAFFuS1s9LYml0fG+PqGndaC4re
WaHEbB7EKDeNSVE+9SccR/X6NdcJ3HrexUK2rmynd0y53kF478cBnPzu2UY+rj4s
15G5BMFMxKnCf6xx7sBIc24WjbX1D4ynMezjHGKnQn3z8grQalB52pKpQmVt7mS8
d7/1i8+Y6A+Ej989QWB/MRKDXeViw3u+yC29RpObVwVf3JfW2up8i63svllryjpU
UMLKMT/r8k+dgn1OIzGSfNYRfmS9ZQnu3tjNLXLbLDhTyJg28lkpyD3Vc6ju+2UA
1scYQFZWpc+fvq88BmK4bq1Wj0SmnXIxCzxCIka0hznuRkJ36/6nxI4yy3apUEpy
HwSGtOJZfVthIOplb0CzCLggoTqa6uSmP+NdChza0Ufi1WhgGHa/WGCxQmayCehj
83lC3Ryj2KGsesInyCOdEhqTRVUE+x8mYkkHWU0kPiofDOa3F5EdGWmeQo1dPbkK
oFY067/LgupYoCnQwNY7solYFEgd81FfT61iXqyt5XvUShXk3TDlGIsZjoKyR9Ph
am9f2vx0OmsWGJpbezzs148fWKHF09gxAODvFOlhS+38BW0iXDD/7iZAQgJeVs1w
lLy9QeN/lgKRtnhNFkclmI+4XDVaZnSligxyb7U0jBV5ldJzzXRSrAdwlo0YnWMA
ZRM4mhlThbmS9cr3SjYv30ObZKDWMvj89va+DnalQLSKpUkEuDHYv2TXli7WPWKB
/UzYd+IiYU9vnytjzit6+qaEI5vZHWJPdFicmP5tUwaJYkXTIgazKynEZB1uy4H6
j5REXKe5H+ePRuRBRiN1rCMlKpCez6t9P/rTb93rAm86VyLOYyqFQhs8MyfTY7uN
OeATYrlXDFYkDZqSt/mtR35gKDVY+0XmOqoF5L12peRI/vWVyKH848vZQD+QS7T5
3GeT4W9sTF3YNPAq0FB0G9FHbp5H0Pe0FRJEAifYKibiVnvcLVrssS+CUo14EB5q
jO+6gmC5gG3z/QwElDXWk9DpprlpKBBsd1nhpbWrbziShxD+0zvZCCTBAUry+STv
52gQ+jUZPRM0rL0j0caV8MV8qTZIU0R4T/mO2lfFhz0gR9Xbt3LVbT4KOtXcyGr8
TAhJwtv2t4ARYT0rhavRn5Ny78u1eVse+iN6IPg8ApMSQEPZLS6uVKWmiv2A6aoZ
Kpxl4u8Up5i0LLsHvhvki1goCHsjD59Ye6AMNsGNNIW2WKT8JpnpkZtfsMaiENs4
7pOklexUEj33Lkd9nAk9LLv6GHgHzRup/xy5TTL9iTnmD1DorF1EK/EIkF1whnXN
q55ozK/rXAKwjFD2MEs6THUOINqJZiOY7COSQEZvIwYdG2Lf+ZPz1OlpA20JbO7t
KI+5kQjqISxnTlILK/AtVL1U3aOjcCAbyvXUQi5OZnnc5+yBiSmvI4a7Dh3ns3ZO
sjb+boJmB2vdz8wXHm47GkGgxnUyXVzge1/fVlDGjdeG2AGFNV+fFAjDwfcfrbLi
HiE7pdcbwVe+CnOanwIT5OesS8rWhYNIXLS/vE67h7nf9lRgC03WlcWtD+ku1/KE
Xj4Wo5NGM//q6jRv7NB4oQg4ui7r03hw+FI4iFy60Fd2SD3Jdw1UJQf5g6xdvAiJ
jSukvozUrYvjvK/UfIb+XZf5s4721vqY6dCeIEorr/39piyJNhZ3qV+jDUR5fHLU
GPiCiVhw7Tqd7U094HbeEma/stABCrwwnZLeMkRDcFrBoAJd0bIGBnWTv8rMvorm
zsdzfAA8qOgluKbAuWYfXGikT/aW/RoY4s3X+ByqqZP9bJHOGG2ECpWleCQTgBLO
bBa6iEqHToCZgOFqzVcAv4RoiTccmCrW1gMidXnbO+Ne3O6RETAm83YKRuuQ3ycV
fC6juLQ5ls9c+ab0VuKvJpnGbwp0+R9iFdHTkvZHZKFYVLEdDYxQYwMH9+N9DDwU
bo42JIr8F29KLJ7fxJ9iP9XHceb1zUkSGxEiUbxYk5+yfuuCoYTPIxYeb4px2lWt
fvmE6k4fYNi+Y8JJG5+KiwciCFUvsK/2xyowDKzRwFIVrK6mMTPf4j5UFaXnOL7R
g76AB66hiI+FrLta/FKyBKykHQ+hhRzw6oVAoos4hDrcpUcvzcS78QhNe5q6TnUX
SBE1f0bTOMFKPhljw1vElONs1JkkG+jK4GOWyJf1In/Fth/iACDwVkwwP+PDKanK
kbUWC5i9ZUwukK41t1MVCeEeloSBRk/zkC62yINnHbg9TuE06Es9rh1GUMaav5vz
9O9lp1nh+kj5uzVoilNX5DpWJOuCI2nTliQggRzC66tPlf8IwsguKzKyEPlerxNW
s5JgdnysqlnnicPgq+MLlDpjl8SD4Z3QidDwEdTmijGk9sJt9muymnHruMgClkkm
WoOT8q3rwKcnF1yvZ9uoHZ/xedYKZFsLBPBfZ9P9ZsE4okzjUwTF20ep8/xtygA2
33HIOJ2/q0hBpBzXIoE8ktRebOAqeewq2vYU+S4K+tllju8RzAtrQNUDZwnuIWXf
EgSmBgT8ic2JjFd37d+1iMBmLbsu8kg69yc+HqXbFqvemtv2Xyx9UR4c0vDClrVE
S14i2hrwbr9fAuTjyQ6lyPHQcNHmu8n7z9GYdLtrFC5cld8me03ippnR/iy3+pBo
S3dIaEnWZdV3+orOQcQPJNO1Ji3MhzZw2aldZeDlYpl6WYs5AHb4Pz7zikvZt5R2
g8sTikPsqMvUmxghGYzFfSOCe6H3bK0wWH8P68USBzh2773MC3NTpJpAOlrXstCd
po705+FS3mCbAbXuVGOBzOzj2spR6TH0qmelEe1Fxh6Fgt9IhvW+oczp/ZShNEP8
Wwf4meu3owbdrFrNm5G4OteEkRl0SDEeTUxrAhj3EzJnHP8KMmeoLTV7mGOSvOWr
2JlZ4cp0jaI24+WE1xXwZvLcSWyPpkJV05WWK20S+y1SZ9icS/OaG3rHwKEB9DcD
rgwlrJ1lT+ME5TPCxUDLKhv/BSo27+yrLISldXxBukvhLMkqUFWHfMcCYmzad1A9
AuI218nP7gErAAmhbq/XfLtTGPPLMdlzxABbi06qXkpaevYUx1UAYCGmM8sQFpeu
dPkue7IThm91ZQjze/tFQJvbJpHmTc0xfg9aphlvcUM4F7Q42vfP5a9/uqtctiYJ
dndneVxvAsFSJGc2rx6KkJx2R6/z1Q7R7eGemevSZq+B8Osv4dPZOUyeydjDUEOZ
PH0/sD7ZWXLOu30GD8heTT6jQ5TWczJ7sv6DaJu7GGnZ5LWJEdVg8HjtbqCzI/DF
CnodA8wHYOQkq6SsqLa14I+uM3eMoQ4hleD/kEa2XqG4t1D7bDDbsCqg9OoUAK1s
kvow+gjvLl+aBM+GCw9jJd5dUL1EBUT1hw3ZjXGH0URjP4iTRpJEMXAwvbI55cCe
gcw3irji4tvZ3YPyyYFmN6OYQ4/ySs3nkJT3LjBAJbSywDp3pr8uXY8expg2Jl5Y
A2wVks65nTGk08dsqNaZzHGocrFLw81IfJ950kpXB7ej7dZD6G06EcL5jFVmeEDt
PDLZsEVW4VCZOH7OHN4A6j/7dKbkaCXQGh3UDmn9MNx7FfS0Kq+4ehfN+X11PKLs
uUbu6fzDrB8wlgj6ftnVkF4Qbv/5NSARqf4EoIQ5kVZ3RDsAIElK0R3oj8KhDvNj
V02aa90DvjkQBzVP8uvVazbXBXs5Ch9Kpdva5ciuiw+vRulpTh0u8bMXI+dIVwdI
AfAOJd6cIATrHkTMCg/yJeVwb9uVo5McfCPrl2W4dADfcUyX9JcPjx+w91aDTkZd
wrwC9CZ4ttv/fhBXlQACWb8+R/PnQhmKvLzymlHN6ZwXpVd6prVYcisHpZwaF/eH
WHRXsDNp92YGGb+3yYbXY2mGEOE7FQBHcA2wVG23U2B86fzaTSQDGo4CsuiL3zxz
yZ9Jl1jGIsysd7XVcEVMxOZNLB6gwtnpugOJEEEJzbS2AAhGRFMxZ/XZyD+z6dYr
Q06zUftrL6Gnrp8J4g/sY9k30EBqchngm9uQKCs0IqGWSj05o4n2eef2BJ3an4L1
dkXBxxMYWbuIcLogxpXDl3kqPD9fMN5z6pU/AQNYakZy9hoZDuBvK4TU2eJMAC6L
XZYWI44YuxZLulr/z0+ylJvGHczKjxs5h+0nlcspr0GA5bheQHZkzmw7vQe4bpDd
kc/wU+1zwVAJjnPRbtyl3hI2q7SnhTxzL2HusP7Pna/9B+FfWt8/ywVebKX5gFr2
IhYKwpgPe5NWkFwhmZPa8ulQG0tKrYnilSQ3LPvguiaBit19rwwhK9wtRvsmN3I3
Livcz6U62G/jeM2B+xcT1uocc6pIziu6wLD7fj5HMa5yIBKyeG7Vhzk98ywZgq00
eq1RXGfqT6NVa/waSaC38IRpJqXfQdQM9ea35egMjozEOV7vsXHEZYVVdVHQYA7C
6JW9fzx1lDSFA50kdduLWMK3L1SMgkVpIxE9bQJGg3pybqhesNR1EvyyS0iMcDzu
yb8GQwTJQwigLC2hXVDYf1YZz9/VFp6nlCRdSaoiRV6KAWDQoa4Uh5+6AtCMlX5g
OwRrYBN6jXDq+Ino/nyvU5F4JYv7ZdjOn6CMFdHCd0bHJXM/3s7sWBcJvXFqMms0
mCRp5Li2X842RexIJhqye+y8ZjtRXqj2n769lbFM+mqLHIXSFOpycd5+T1+N9s9X
vD4DzPLccvbCqxnRg8qCKApmHNRus20PP9FZJtU8aMPKkilhpilNevJgJ3jqfrz0
41+8+p1Dc+llPMWK7CEFDzFJKjMAy9A5jG3ZpqkREOOR7oVVqFQpwvbSSB5sJIpU
7oUFvgXpRB5JxVOqVwBrRapvXU6brtAbDIqbL5jtjQKSFobghcL/NQFHzsxIsmCO
6SSClk1sby1x7PM/xRfzhfYs85L0PIhcCZhfcXo4f8Q/JqQSDLgx7pWgtdHWFxih
ObQD7/ewIjYAgSMRSBTaUj6T6HSxNC+H/yVdHegwENT0p8xaucRhclwsaaUj5nT7
2LI8aWGxOiaq/LCK1HraByubTEUwyogc0tfteX5sSZIUPYG9zQxnZ5a73O0vGHc0
72/AavAnorGfxxGkzDe+/VYTkzu9++TuTDlg3Ur3MnbZ64e8Fp6CjXrVsShrY0km
VePgaYNdHIr3n7Fa5VCyHY2Wh3bHq4W3YIjG/pBSRCFcPYucAtxPuNJN7w2Yg0ZE
KHXSv1JxOlOOcdABexqjoH56+3JVN6O///quIOwHRD5Wfd5X8IsphHbsZNh1PKWU
QM49VRXnPuDicVcDnA29lR1O7v5SznWPyhEMdjUsX0xWVAHdr6AEXghAaDCdE87D
y3lFBk/mHU4Q+qZMFJJJeg5Y60UAvKieMViNZxHp488BShGRxE6zmRKbXlTJc8o6
Dy06KxSEZbSamqESZqc4fOfbFCssTT5rD/E1Irx8zCQL0Bgz6J8ICc5pcGhmBuVr
P/AhLnHXXfayy84hxLaco3G0EKOyb52KBTfL2/FfW7qVgPUgGfUKIWEGINFC1aBv
KqSIispOmYqSHzGzSuGREg95xKxQaCtwdtw0coByxzRgTij4gudPWp6qu6Sv1h30
Y0dymZ1sMY23TcW1fYRmr3tXHt/Swf/zjzVBEKFqTfZ6j5CFUXp7E6EyI6yZLgz4
47YzZvkTu8RrIx1Aa7IrhRfCD/D/1GCqQdZ/2Zrq3V1TF8fO+WS0j1iz+W5jQtk6
Zp3suOQfvCCgq2rUqDeGS0kZiEF8PtllZ3aAO/UGgaRbAvFsZe8Bihkcz1YNoDaa
TvsGQWDwSRZamF9eLmUUuTA0VDOG75iBLGm3FeanPSNfwr9tekpzuLA2AyTr0wvX
36lPtTUFy4czVq1sgYeqw83vm3ajIenGrR+mXARCg/fv8zycDxSmpzZFLlljtk43
V0DC/Z412hD2XZV+w1P6RWRiz2a3Jb40K9cPviHxvJOchVX907M2NXw+p8ATcQQE
Wc5BUeu+/GTsyiWLbR7pppg1f7acjSmlun4iLNAVe9YAePI49usqUckj0EPFQFsD
gkXfj9MyZslKwfdH2LbKCf+9e6+3IEdDnMVRVYWgxI9Tj1Sz82qeI/L3mdjvz10g
C5HAWxN/+rjJqYOjpRam/XjDex384bt0Lz/Jz9IGobsS0diW4zLNw/GxYAlV1tpy
/R0j/5lc1yvaT/aMJq/y2J/gxzNTJKlup95nHiwqEhIgLnadey8qZpuhecvEQBvJ
Q+B6nMhvtNVlXsY3Bm3BYAESyNhW+4svW8x+xESQqQGUEpnK3mZ5t60UJ6pj+zlE
y80+nHbHvIhevWmgc2beVvekzSIXa3bGiblh9TRz4ofiLHe47YbEKuwAEyCNkbCL
ml0BU5NRXAug9fCxa5K/VB4frJurJSGJYB2v8hHhgBjj7O0QdMPd/C/xKIFSPC24
h5924cn1MaFanRAbKJvW9gFvLTp+oukKxxedrerIkC9Ga8IVdELhwOx3ptMN1W4v
gJ2sLCYyonCLKORLZurjr5DTkigcT3M834EKrJmoTZ4UfHS7az6fXFpaik2Ha4nH
cbGbXGaoYSx1E8k/V5jtFl+Ndki+jVqCrBHa/vCSzd0lOAev3K4+DIV8s66ZkBlp
9TRmgLVtsNuV4Jl5YY/XkbncTy0rDFL4oAnuoeakp8PShgU3WxerdxvSN3FGqRHX
6765zDSe5sOod14+qBRMRNHV4MmwA5+BBgBDTIg6tmwynAS68n/nOzzjOZiNISB3
3QDiORegJWbPvgrC8eU83Bqp+cZDUJSuKsW2pv45b+GC9OCpN8ec1zMiS6WFya3v
mMHzvl30Gx0TcGN7NhR0HGiMGrdDPhVIVbRktddZFWaMUML+peQgxfSjjKFhvUc2
fWITT9jmhVwCqlSpN8YRifsYXYu24ow2dJbleMXetYONuaFZd4l6j8MlbpHJCdja
TOlG9TSGhWTpC1HEKbatuoNLZPgvS0LQ1WUTCBteSIpfLRFAdiVNSSLW1u9s3adO
mRPElU/IaHlUM89ENRhukSd3+nUckBlsrX97KujS8O78KTgJKdbQoMMkhuTboXKs
L9vfbjrElGEE/fxuH3oIvg/IncSF/jXpT+lDavLgpBdmtD+whTjPmU0mQnJagbZM
K7PcFTutDMg1jItX/Tqm6vipqwEb/a23RmPnhjk9RU28cgO3/P/EUu9lTPd2Kmue
6O2mwF656u6LHmUJ3jp7Wf0u1l8fPUvv4kftWnB3/q1b7JspwB8SGR+26HOIe3In
u0xD1aEZ3SXS0mNBsCVORgXxdEqfWTifLgcmv/Y/SiyZt0jSXPDZ96qFbsS7ya3V
DirtiKJKwUWU2owMThsTabrDpLY5S9H+sv4EWASitML4ruHi2jwPeGWEcRzcYD6u
ZgPa8XbyISfe0cPoXFwpGNc2IZTjB/B3Sn4NDGpsq1elRSUkWQfc/SZ5pf9TCuh6
kK1bmBjeP9YLhjipOhhI47JPZ8btV5EXGi9vpk6ltyvLE1I7L5zueyvKhE81MHI/
T6rf9UryOC6fWVmDTmTBvzcWkE9F87KSI8mcdm9pE7rPbDPILhyzEbI23iHZz8QW
paynZaYYeaD/EOiWnSVuRuiBil9caQht2auSN5FnmsSbRASUTFkhhS0SiiZVsy49
nnu6fDy51j032OA8Z5eN3jHlWtGLDD3Q2iPAie91NPF4SbT5R+4BVqvjWlt06kcs
iiRH7cnwMoqk/Je7qz+8lsJ6fTsL55yYpISuarAjy9b7Sf9MGLfbK5i4hPwZMNsO
vpRNZ0x/FFP04diW3g+7xV/WlFU+8tbjW1jlw8hW4clCBL1nta6GkVuZfp2mpUbM
g4OWRfLBarpkQGdO030hCW86mVNCCGd+Ur99s9c5Uuv20X6u1tPhnLiCEkbVi1c3
UxeS1CN1tBkPfv9KARMYSkoK79WsNvS9ATsJX7cbl/Sw8AnKT0W7YUHb0L435pYP
UGOD8e60bmX+f+yKd/e4NppYnPG4wx7ZyfNfpiKUsEjdf9rbTdpG2LzdATZ4KNIL
+1xe3RqhgEDOhpRdDszCkmo2n1l54RD2zTOJceBNeZn23W71kPN03uaQ2FofGYXq
IH51IO5ZvkGIvqyO7TDkF1oxGT1Eu6KWUbIYGkZSl63HrvNaoUuHm8NVR6Fpo6mv
ENcXB4WSLNO9L6On6IO8J8eSj6rY0u1cgAkMCSL0rMdiIjWkPryOMj3OlGLID0HX
tEpNtqPo/RrbaZGxQa3EUvAR4RIL4jASRnYeR1ADgA047VNQ50atD2XfZKiors1+
Lpq5YJNDAi9AYBHyH4YXz6Fi6j3LLh8Cwh5G8nUxu3csd6bjnRHR1oURl/CuubjD
+cmJYRixkJySSJLbTSrQ0MMgaFuSOZ8colTaAasxG6Mt9Z7b/PeyHSvzCK22nyPu
H7tnzneSLSbyt4uZVfjJ4Qs2FkgQkGrhb3ab3AbvllTfQfSbznpgwYHIL41Hvc43
puZ4c8pb1IEGxDQQ+Q880mi/AjVXIRmaxYRaspXfIqI11dNhZXBJSkKYXnu4WnKw
PSegqEz5lipHXFHJwwtDCOwxuwc5Pwchblw3RsWsXurpygBR7nycq5BuCy7GVQBd
8mjFbO2rwsFdFZY6ZseYVTMwOoZaOyAa2xjN6Fwxgxm18+IowSce8gybaPbbRffn
m4xALc25a2skjtN8LkkdiL/nzrSGnUWJ3gj3NtYHkOPMeCIZ/bK0vfWcnCGCYXI4
d3jCOlEju2VBd65do6XbUrfMjqPHYkaAsP1+9JNR7pPDRlqWZ1Px6/6i6SsrertD
HogbA8IuYzL1CvSLhDsxQW6UPF8QEzAWlMfJOI5jwfZ3xMdehU9+yN1E5YH37lLe
TfEfj2TtgX1sZdEh98cYcKwU5VHo+h+ZgYaJbq8uzBOOAnqf1n0n+uiRMp4yc0KN
jDuNRwrI6guUbee8G50xq10lKaYbFMx4/ynCB0guvyPDlQvzdM96EmMWOPzVdIqi
4rDf6RmkS6/w/RDtuBkG/qu4/1T+Hp9MBn+802zj4nksLPKhB2Alxvm6PAyOZCOG
qWhHo+Q1UPzoI1aQaDKZvC6SkSvljTkMT04W/NCrlYKAyRsWA53DA77xEzpsWvsu
rnUHc/B9lLQHdALJKNQ9dQNL7RDp1pa3XU6wGrmx6WimLqd3DFqKwVF3hHFz8IAH
Z5HoWqaZixhTvlrgytBVs3wDzm0tPHGpGUcQ4KUX1yqm+QIFP/EWpcft21L4o1m9
o8Ml42umho3EmkC71xqHvZl2nGcix09OKMJqKWg4ZMjipZFkpmBAsCZfvs4Kagi0
7z8Nj4jtvoBiyL1sYfU3j+u5+sUTsVx/g4ND2OJhHky0IYxnPxcvGSct79vye060
r5tnBMuWz1XtGLngAri4XNnQDqDXbz0Wp3rXXC7POEduPhLekpsWxI6fCi+51OZd
t75YnsbV8p4dI0abyAF+/qgTxood47eEJih2Yphfl/U2qUaiqG8Ep8JsrphELKIK
7O9/kWstQZv5Np3tuXlzkL9zAduU13roBtik3FpuMrDD6CQq1vcCT6JCfxyaHe4p
M3lVZyBACl2LKG7ILahnUMqG1fsXbR0FT2vZ7EMJAUqihBsYNtee0MW/3nn3WPJP
TcfJ1JNcQq5k8P7TJfPUf7XSHV6JeiyrqINbnNyPosNf8HXGHWyrH8KT5JGG8JRz
ExC/U0y52FtLpFCn+g3aTouHSRefAMbaY+luSm4suCnJ6tlXcp1dWSemn23GZOoJ
ebRfiP9hqDAqz86pTOjl59QjahPbSj1iwFMyLWA+VVXWwxwoI2salGAHmh/acwFQ
6YjM8q/QmG37biX3P6WSy0kMsMgKIhR1+pgmSUAKXVf4BBopYyoCLlvsWjAv7BpJ
dzXQKaY9wMxfXl4GvZnPsk1i3WaPtkXsS6BACAMk0dSeZ5ykEobVvbZbXcaml2f0
iwsOfEuCx7g5wQomtM+r9RSic0UlUprcRA8zU0o4AtFBortr/T12ZZi2xTJHaiDW
OUslZBGgrg45AiKNeerWIAz1z1VPmSHjLM/hcQMFlowfy3m5STCNYIEitPkLoatZ
+WbLiezlDlGreP7v2aLahwVjicA2Qbsubg/Le9HP+eFd9X3NnnKBfuhDtF9dVnM1
qyKrkrh6pa9UUcvf1lRqCWTte1yuFddZQGFTwh8H6hGuMRGDP2laeKdiN+XnH3gk
eR9t1+v+kAkIvPFqVqTj3ZPlQxOKj1tJTAU4g0/ULWyuciR3ifwRQh73YOtn+a/N
z+aK2NhmqTgPcjoqi0b1b+ByHvQphYyJE5maH+ib4NnsU3aEMqRssjD0TLELMtEx
tKqmRSlmpIwDV2uHdH9Wx6d/XtKtCCqljyEfcq7KisolhhnENA42PRUJTsxwfD53
1CYyRHd25eur6pbSEWXTXNdEHeiJgLUY1JaHppqY9FL+gLB/1GaAHDw0NSHdIBF8
Nq1m488e48N3W9Ja2GeuIoV0DsfRHCt+4uDVUW165YFKBoxxj34UcAratDZuMdgf
9gKbyxsJatc7P3taBwI+Iy8ewTcQ4Bpl2zBq16rnSzrMDVsoWrlX2OLVbvH6lgWm
VbDAQyArizIjl/+usqvodF3x2WBAgMqdmsj5s3qU9FNJrSlDagEQ55V4VfTiho/n
3ewZR4xZ7yjy2iCxm7aW7MM4/EJp9smGr5+g/t1Uq6ye9qm5PzcSO51ZFS78dpd+
E4UmR60g/IBbArW7EjZznaIaP/S4ExA6NTt4axcORat7SwXumrtAiYGSRmB7VpNn
Ass1GHT6PvjP6wA2kxdRW6Da2dKPgr3Kvw3ajwuF+W/Avl8a6IzCICT1mZQlRzBx
5LuMEWymSvWg6gcyhVj/LN4MkUc/t9J+nvzZYaoioYow75+mIbsfTPLJqC/DOcHx
z/JQRkSfbB+nldUXedCtlYoJCTkv5+XmXTJDKuk2ctcZYVdvxZx4ZQoV/imvj9r3
n8PlorMO4/aeUfAQjPSnAmCap6FGgx+FtM/nKdfzyF5TB9RbyH5obHSBBW6hCO0e
sGpd8ODdgRUUw9pU8cd9e4fF2uDo7fbUEAkRCAJja9jplnpjHrLrKsKAhIYM8e2F
nZ4xJrCisgRewamOH1AYlliU9XPgWFd83Yz2b7tciLrwrYe8/pTwu+l/2uCZikAj
HmiXaB9A+qfsrVcvzCYAV5n3Lh45jzkx+7FF81y6CmwhjN7hs4TsPSBVROYemnfQ
aU9BvReDrVh+b+X/JTKkmRw5LJBsEQ8mJJS0+Zg6hwfoFG7OByj+K2ctNmWaKMxq
G6ikHD5vRPdblfwFDDoaD2AByD69Ex0QaklXB+8Fapu9N8ODo+yqV7XLEUG8B3HC
UFrVPzspcgnnAV2ENyl87kZHxZBEastUlq4RZZIsGnFsq+2uOS60ebAtd1k5YHW6
fDGIVxvBi/bJI1KvCYyLDKUi2VHxTBA1dhlcFxAauoEajMksKVKOPnQeWBVJ09LD
/Hb3hFhIe3tei09LYg8qTxeIMkjkLQ0r95jzj9kCbbLV5dONnB9Vjh0jpF54jOu4
FHsiYajYU6QNo8Pe7NwpkGckCG5U+gBTuar74nPvbFl51JW8+JnXSH+mE0d6drxf
wsHhzeSiDerf/3clYtTxfRrMC0gNOCMYOSytU+taNxxCJKo5lSlalnTP06MGfGcx
OJ0bY51B4sNqEFhu9Cm9w1zlokdsx1Q6HDh/R185FVcCUHRkZ+pDel9nWRiIZ5hD
jLN4520J6vtmBvbfdK+XAQJrh4zAxUIvoMiArQ2pehDPWe3h54dMz5FWmx/Lkz3G
O7avH1M5S7MltjnJjUnfIRYVZyyt52cWefLFa4w6Ze1NQo+ZHp4XquT2tQcMaHBW
+Q1DfjFufGG6jprCogkyv7X/9WN3EPOmc19vSty0SQO9R/e1jVzr5OzyNWSLgsko
syAn8DPul8QiVtYywAJheW0gUXRWcM6D2o3BV4Xk5WXLqIpRcYZkFSaBPrZFgjGO
LirGDg8m3JfRqUp6M9m20Lqc3hy3RTtqycOHiN2ZiC5Y/l+VzPUORPNPKD+uW4Ov
K4DWGzXvZp5lzhkc4jl6fOoQy7owOgkFvz1Q1RrHWoVbDRYHRTXxxqCsTj5FT8QL
UNdWFcKaY8NiLOw+J1ZbZT02BNccZU1uKKdYbwBbMiDpBblVpLm5txHCAnvEm2KX
sb7elsMULYM/I55dMa1+0oIXAwiqc1IYhvK132pttRvweN7fXryg9FWNdyUD2U/F
EHM/rU6a3ApNnZ4Zu0sVxIte68epRRrBp3kNQDPUkhB3iB0ud8FKGBnGYkT2eLhj
iCdBKOLnfdRk0HpMhfehFE5hFF8ycQrje8TrdfXCvG+RNGkT4w+bsG4KyxA3jKZT
xORD4kqj4nCwnF8XwivnU5hv5XfDjVQ1mZkZS3CjJPFEK+JQOlxTjKTCVH4dHIKP
Zn42BsfHpt7CtwqieZHE0fPA42QXlM0FWidriKsKcran3wjcETu/T55LMkzRCTiv
Hv3B4/WxsT2U/5Jk90MmvulaUAcV2YYkrIkwCeNq7kK0AQh2dRIGypaU4JexXABL
tXs+BYTKhEMRsfInLoN9JqqSfdv8oCzfaNdYGXbYqW/A7yTE562EEZv2BLuHLytj
Spo8iMjTaJXG4Ti+gnwMsP1PHRy9yqUpOOHSDZyARtCjxDlV4mtGWJrbAw81eB7M
getI0zAuV3/G/aPasBzGFikWpAlSuIg9EG/RrbfbxsfKA7dp0eNwhI0r8pJXwQZA
VtYgbmGPNq60KQbZ2agIlO0atYO74FcVNSWK2+tmA4WgSF0IlvsbqhIT22C6thlw
sHIbrI84D4Rk8MgN4niBqMf9Sac2BTBHhO9YgsSrHgkPrfpV4U2JTix8CwsOjjKt
BeXuozg4WuKMfCdEGp/Tlptz2xcBdsLqycXYW2FEW9gID1RlC0rnzMCGN9HxKyyO
Nn0i0wsQDZJEpcJWk2RPrsf2gZNWAgMvqNiGO1qgjyijtrf9Dkdraso0ZV5rKXHj
IvL0KPdd7fHvClocTXieSqPqlSGiAdIYqByQd338DFFOxJNg0GPVRR9JZXQmgE+d
lsI6wYFasfBzlpzXceoxqeUUVVtlJjVQzX7/19+IIU1d+3ZXKexTVKQ6qkk8hXYX
I0oMWlkBD4oIb9u08eBclCCoAaFS6ii0VVZ2rKRAQ1VFNgRTXNQnWkmgVDHJlR/m
dfLKZ/mX2qifb0uIqGftBbnfDXasZT3EjR4ECO25lfOx6mzvZD6VK/fX6qhRTQrZ
rhS7WB5cBIs9zNkz1N5hl8xibZtVwtS2Q5tf0D9AS1UEC/8epwvjnJg5cV3jPQ+Y
kagIDpWXi4cjs2jcPULfCycb/X3zg0Iips6UlfQHYUs8tmN174a30dLkWyjsdAUO
Q+Zxn3XLz5517cX54oKTAJ+u+tg17llI1mM+Rt8W2W1ajJ/jnkiwAiK78b9rv1J1
erIAnWom7Ev13A41rUsAQXjaF/Pxu7RleIxL72kHMXN8WZ1p2w3pJEYwiljqd7s7
HsiB2BT9JGcwXODeukFbNMObb3NSbvMsYxGDJNl0VX96j4rZtBl2gK0RXcQZ+8id
e9Uvnxj85vCce6filFyAuyOrtqIf82qHuWoP+wgt0GHgoIu0n50UnQYxRVWLpFU1
kZ6f0x2LSGvm+vZHGitGfdN3pISLGpC2XdnA8zcAUU+cX531KheK2KA7cgozGGkd
SdIDaaoxMoszMeA4uHjtvpE3Pr4JL8mw/bNHQcpPhhNk2orrJy53SxA+WiMlaLSF
igatCuDFHi8zbqXluLfViXWqzPci6qCrauYyk5MgQj7A4itdSslblSHAWCqGCAwE
/oRxquomAckN4CJ6ZXw4AsR9AooPnI4ANj1BBV8k5tZ78SJyJcgiSQhBBj50KslO
FuLMIaTm+fO2HO1peC3NU+KSNXmH8QXKTKNCwp11Dfm7e7dSDrNe3Nnn4PdM6QKX
a0POwaraVzyX61tKAsyGg49b7TRKoPZIpFZNCPQTBZOiOYEd6fz8gmCet0PoUYIp
TqFIG3Ak3HME4vyEHrwaI/JaYzkgjhvcu+OlXGVIhHBBlHY8opBdpwTSPxCH2gVE
uzXLJsvzVT3mwrJfQ2xmanf8PfMz+SbC2ID2+FdN7p5AHLhtRMTDl0S34hu+HBKJ
uXm0xpNcP62eX4BeMrs0w6jcres4GiSdEfiLa3VmXmCWzEfv98JF9V7Av+EXXwty
IzOtp2g/gfZh2Xw/FnOs3qQhQZB99zdFqA5XPCWKQHv2Wuu1yqCxiidelCWgnu+2
80MzCyWIF483i9J2fx5dDGwLAC6xB6jEswtt+SS1qReYmTgp0opm8Is8PbcpPD1s
FwX+cQFYlluJOsZIJrIgSguA9dTMc3P0La531JJAFT44F8wiPD/tcIGLM4hHvGh4
FM0ZFAnH7dah5lRFfoT1BRpGo2C1/py4PrghS6aNR2CnY7OcGNwypFJtivdex7Re
WTTvTIRz/7at/l1tzdWAEAKqO+18U0sTu29aBTp8lOT/Bhp1jrQrcfUgCDAO2FR8
MdE/wkAArL7OT6vDt6TgCLTD0AiXdFq68STcef5uc1f/y1RBZQP0FteQATgE624K
2dmFMstolHFSjaKhhIsZCBFECY6WjzGtI2+cBDhpjz3A5w3FidwagkGvPREEFklq
2VeyWscjD5YUsBZSVVGzDoWA/glD409Nd8usf6pbsP3sjsBPX3scy1EmcLQ5mH9t
1z2Yq/Ts0RHJZoXp9Wqd3MrOCUBIkf8EFCVeHEUMK62o8sdZPvjQreCZL1o0rrLr
F7pyr1u8K0J5wyGTTeSbGVbZhryyLi54kVME4etBgU9BuYtnMQZQjFQYHqFHl72w
AGdpb+h2wHJGcIJ8dlVl+620TGvIAL89+hn9upZVpbLNuvhS8T8SFKkImEl1wPbb
UAVc72B83WjVCoNqm37LCmzmd1/ZrCVq8QeMaevlXgGoDExtudyE8jjJ6Sh8SNhW
VLo1fgbfhcU1QZjkgGm4bKhyOsG5AnRDUojOIofhyrj2erXGKYAG/LK1Ktd36rDo
iLPXp4lz2dax5Lsyke5HoFz72xefcv6uNnTpswxe55p65+JWKPzQREy2P6/zEK1R
K57v6QtMDrvHPUSpxdUARL1TP0pdxTdqlgrgOwV2FNS+p3bDD7fL8NPB3To+5MAW
bendR63yWB0g8bpwjjmL0/gpSEELc8R9SR3NK4NBYmxlmLH+fNwY5Xzl4GjQwuvw
wDXslESU/SHM3Eg4UA8A/0f4z1RzgVeF2eQ3cnKETP2lmWaiZQktavUhoRvtHp95
7dvbk+CQTJi5QE5V+vYFi8S/0j5gSBZbt/zyVlNR1ypf7+2idTD21KSXHY2bePUo
bzzYJqf+u7tGmYIDX4FDO+GpmiB0afv14Lw2fDOl8EvtLoEXGh378PcSwQAPQvZA
OJDneswPQUzClcbIJHSwwxa79Eu2vzIs3TbjpvrM2jyAvcT5QDxz/wF26FyeODrX
HUmwWpwSNB0TfLzUR7sbEvyl0RPACbeyBgZPkn+ZWXhpW5gghCZ/jnMLLUFmvqAz
iJ3e+q8T1ex4XvpwLnGCWp8YDd43JxHiIjGoFZWlLO4twr7ROrwbw3u95k1TLG2r
dO1/U2E/qpwgpoOK3ca1J8ig4hnppghCW5AZzCZ9a6zfDFJ4zBT/TJe5zHoKao3L
GILy0mYjnIqNNYO+HouR46VgFmJar6wFqOdMxRdC54WysWn7XILtD/xk4EXXXZRK
/g0/zaGkyrwu+M8USttRU0B0+3qMbXyk3RzZ1oAkJimuNNhX+N34yjtIKFoWnnTf
4GFii4bKoBL/Msc3PhbQSVceycRYXjOr/N+CiZjAXzgH9m74VKA8zuAQkDX+wDI9
OsE1SmP0cMVLZOa/bMHo8fjfYs91gmK8QQyJVyZEWIlkIzP2Ov6b8vKFidkTnP6S
vN7qmdcxS1vFmW4w6ducTZ40YprLx6RN4kN6AXqZfWsmaUkC0eBbKXBeT9SNqOvv
wQNZllSZfPLeWVG5mZgu2ILPZ749eoYLUChwAFuHXH2ThFWcmrT6G2x5BcYAa8KO
p/7WeSi192iU/O1Xt/bT9Syb0j2+A/Fu4FxycVd2AbhjPqJlD344UPq5/wRWkbO7
JwgN//6UU9hDCeGbAsn2DTGg3+wEIPhFIdDbkmJSGp0XLs/nSUjlv0W0mz1o9zYb
N5oS7ZjVPpmAl5tp2kO1Q8Thn8meWI3Cm76SbLhNcGemLprHJqOOy+1EApishQa+
wKLpMHyXBdgogf4kJnHKP6QbcL2l/Htp7jJXYTPJGX57xDYlLBLwu4Wupt/SqRqL
7PnmX5+GmSpFJ82gn8j8zq9IlKKaHy0dthbw1NUlLc80FSW5b58u+hyVbhAEBDcc
lf88giNu8k5SJdgYgR3+ughPxgoy7NcXWvoAVu1o+JITLqQqD62zeCPEgV1GZlDV
0UDO/8WyO5U/feK9/z3kuXJTMoHMY7q9d+dMp0J4sRrO3c6uPgNHftV61I5aB9N1
O55ly+RF+Z4kpUXgWIPwbjJl1xIYgE87UV+HUPOiNZJaNb2OL0Pbxpzky9/fNlqv
GIUxZqEaPb28w6ux2Ap865tTbtL2/Xx3HhZS/Jw61c8ySdXJ+xqYUqzDAABZzHCy
VWimtedFrckvXMY3UIkfJgYJIdbnZzO1ojIPSUgEdSVvQWMy5+l7IjVbr/ws64lg
ONvQZ80DfRb33N72kiN0vgj/10FdqVwWCo9826KJSsHHz7yMSGAsesJaLsLLqnOh
H2+cc36EM71oxWT5OhZ6EO4XF1dw9hRLvXz4+GNIu+R1PBwoEgX0c2KH0lkNONWG
n5NPJj6VKAXeDRCKr2GAWDRouxrxGGy+Jt1MQuCwPHJL9C6IvF1asoB0hM0zAG34
TK/waGiSGUqsQL2ufgrmjC7x2HmrRUKAyIbWEo/laxYo7LMKpebydKyDBwE0/mxD
Kl/lVSG1p3Gq65VtjnoJRjLBLR+3kckF2RY/3q+2vp/95kYxYmXmJkz+6bY8buPf
hGGvFyJ86ABl2bj9TBP9zuv/Z+R8JChrHF6OQeVGmvqxMKTwCbhPo1N8M41UXrDo
uC1eqxbyLs8UxcVRzZp+6FeXHY97zVTZHXlFp8VTGFsL2pK/AaLzCRT3Qcu6RRKi
efTL6xMya/pxgW3hGZzJdKUqt5hbtlUW+Oq5pMWyoNsvm8HFP5Wds6sRIek26w4n
439ZrLvV9kZR/loRBboF3/ExScqNoBCAGGgikGYe18k49ivC9pwiQX/eIxnAX+/H
QW1GVPLrz6/eFJPYNLloKWWfPqMb1P+0ajbXO7JPI9BRDYhOJX1Re1WiHawyCUb8
xry8ohNcNdzAk5G1auqIyaxtiXOYkX/sDJoA5ktdFoHbfsjoVlwyiwAYl5CM+QNy
WlLqTc42f/j2t+lNg/zDSRzIYDSFULvvvJDCDzMMKnqIqnI7aogoB6rWZLsnH6a6
d3mJgZOWfN/qNQDS2zcF8AhmeVyE/mj6LERvcpQ9/oeqIy/j+AEfArod2zHwzZVQ
YM8im6O89dtC+NjCJtVULyoBC/dv3ErzvtxVdtzjfT70V8idEPlA7H//NHmaSiA5
xPXJCXRPakEB790gTJdf+Vsoe3FPJJTNKmcR7pOMhDpSXR9Z1Mwc5Qde+XPIZ4ci
flDy5CkZWTC7116jmOSupn8KNPgEJWBDk6Mj59sgDpDh+/ERJVkqJL6xUzQKAlrI
DjMIsY3ELo/QrgVS4OgLf6KBZvMvVuF44lhJiS5KCUgDZIM56fqqEhW7fn2hewie
9YX91mKZeLIOGYnzO9kcCzIvTlBriFflF1Q/gof0x6MxM8BQv0fSAR0BwmBm+VO/
S0UqG2tzcCxAUlAcFUgK38LDZfGzA4yij/8WAYqd1hkj9xrp+FJJWfVXTvt0Ryf7
79lPgU874a6RUAJeQ+p2NHwj1fpeMVlKIgnFH9JEwy/AHvmNaFx3OgxMnmV5PWY/
W1fz7vUYPmgUBOjkb/F7R7exxNdmPPDdxeR38Q0BC90+p9dOLy17naLcCk6z1N3g
J5Zx06SswixFR+pM09LeJcSI4/NOyJ3acj2C4AZ2mkpeT+lLmncYPz6JtFtomduX
J1XewXZJMiRyJjA8+/tIw3qz/+ieGkjAURCnUlykUGFo6IEDoD6MuQ/8K11CQt0d
fiWjJzf4RvfMkE7YGCgehpKTkjiPO0ENw/KBTSli5Mlq381bwBjiRQG34CBHnJz1
PkrfWADaosM/CJ1rezpMvGZ0wlLky+pzjWhW5vA3xNLNdlDpSA3jS4szYEUBjnpf
ZsXbXCsDv5hvkehHaKVimPI+0m8EfXg1RdGver9yI+5tE8AECUp8BKKrzdJll0dR
SBLc0PgqGME4cK9MWAuJfDdlupEzLr3eKViHe3VDsvM8nqp06EAUtbswjVdAqKo6
vk8rv4bHoDoaZTZOOMuI51j7uxX79t7DHNW+UJSFT3Y/igvcuE26iVeS/i93nUtr
7vKyQ5d2B1g1da4yKzlc73mvJnrOTnkm3DfyWQmBlki2ujFSglYuDCBygiD1rpJb
IBfgn6AagalJAeJicAE7z2O4idRohtHu8iznGBDSNdqOt5vGyAjLfsTh3l6xfCfH
7A3azh0rUHMTOy7XiwAY/TFp8VhidQG/DdGNB6ZOgIq8w5h2M+9ZOgRI5WU9v9Vl
NZ6Gia2Fh1gnEkP99+o9llzLniBrjWETbAwgBfL3CALafiNRZ3//bFqYVHiEtfdO
BUfvmHaScKv34uLNyhreNcVRtnawk8B8z3V4qjVhDnurF4EA6snCGMJwVrOgjDYI
TLDz9ayqQQLofi0Xn8if2PUCzqKPJdarxGiBQ6I1MVhYsOqS2Oz7wc7uoGGizePE
t4m2iyiyBwtxkIsp6dzJ0ZEtM7s6VqkOJu2A9AXHNg8gu3xXK+hiu91Y8DI7rA1t
YJP6kcmyravxrXNuY93ytRXo+3HgRntVHZHVKCHVbLU6omHhKfAMGLv9t6RRUGsq
dwPg5ZYtEZicOfvquGSaBJmEZ5kU2rRSK4/+OytMsyszvZdMgYPBpu3L00S0PhqK
eOb6xiIk2Ql7mHTae2aTNvv2ZFuijeBIP0lAKLSzV84Bo7f67LZFeDQJp1iqRi/Q
71fYO/uHKKBGTyT5/5g8k1JFALgq6We9MFbnBcL6aCizdEIRwkviiip3frSAeD82
WNgeB+PY/JvL1YykIsMoAqyXpQ6wvE4pI23688tKGHf3cH/HwynCoPtT7GPe8kUf
ANslbzT6Fh2x3WaCIlIdJwTEbciVCELgQSL6iV7QY7Z+p0bZiMomeuOmvVSbWkfX
4JQgXHJCie0CX++hig+vSUjljozHTgliJN4e/DhpcCOY6H0XZ+bTWq2sIp3K9fpg
Qlp3MgkxvUEx5DZHH/49C7lFocHMh5XsP2hRoAz46+vGzDHJKRORKfcUDwFMBX4I
Txiu0DabjXahbERYOOhWENGPrQATc+af6TNGc1uQcOpT3KDJCEmP5xgY+k08MGLh
n00+0YqoYmX92N02dBgx6EJlqz7TP8v6wIMw/GhqkqY13OZg96IEWM5yAlMGlfPR
aUehNJqm49YUgHmZZ83KDLnkx/ic7yrpJ3qof/GXMG3lC3bZN8U0bitSkbuPZxm8
o/hl+CCWggbsRsqaEEnE7LWyker1l/ml7KW4w7Z+pfn8Xg2T7yAqOsd9HiL1eeKL
40rw3EQ1Gd8KADk0BQmLVEQ7HhUflJq0DyscmI7CvspW/j2ofEJ/4mBkRnzJJ6K0
bihVDGkOliNwMfnmXYPAm2JoV7xG0nksv45D2Zn+CU13OAUYMhgfBRv+FHaGf4yl
XFSDOzlJ/6vLeqgKk3dYbT/jH1OGKhzBBV/BUdBRmDcMGFyE1eu4/mCsE3bvxI6g
9ypyvibZ0rAGLP+Sp96q8z46zAKgGLBYAgWRd1QOJaE0xmcLWrZ5VQpspQD8Ujqm
Crk2W2nsvClLhBHUjeWHNN3TAL6QKKT+66UpMYhhC0RZbsz3AE2GEpV/j9A+zoiw
vefncmWunYZ1NdkG4SLux7o+pdClJ8yDmuH+hw5fmvzLl+gSK+xdb8VSdB/GxhL8
e7nTrGrCWVOSJW2/JZ0aCDnbuc8UJlHi1ojM8BJ7LAVr07NfDefgvjmiBbCnP6og
cwGVJNROUIEZJQfgiscJEQSIPCjf92fkmZFXH91qlXZPqKsRuGhCV2Wu/tgt3qPB
0QbmLEZaj7EWCUyWfMWtaoCk5ah1xv/V/Pz9A0gMpAMnsw5l7Fb5JdNBtr79YDTw
i6Ol3dCCazXvwB0tWB23/cIV8IHcNFdDxMF/lwf7Hy3kJHF+qrUQyRfFIxkXBcW8
/VKbTfg7uVpftZyCyINMknUhwdwMqGSqjY3kqUpvTwHimhFoHmfKwD+Hrx9XuFZr
6t8hF2VfEEpnEDZrFYvbfjv0aKIDV8LIsc3MIV6XbiBxAEWvHb9rDllhVrKXEqLG
pgbbhI3IlVvQmJx+XlyT53M9DR7GPXIJ5jsl6K31LAoFuM+LerZ+sWoHD/hbleIN
HVmsTf79sa4aGz3sP8CPFJZceSLOWyWm0gbRLsiNIB4B+gNuA/qmFIpB9hwf6g7h
2bzW4uW1Rea2WCDiQXAnVjsOiGBWthIjwkonMXFmgJ5OEY9E2US9DCSQXtn4IU4q
mtXVMmntu4Kv6i9THDL1XtV8AcORjRUURerOenSfM2uLbIGGqkjBs1Hmp/lysKPy
X7uWCjpzI4Q4+kzqiYPrJNxiCjoA071jAs9SRRMvsASKwbnwcNzt8Uk7i3csF3mT
CGsJuARqu+HflFf2VxUeaX//AKdndQIOSMl0uAG1BWtzHjC+7Qr89mbe0yzGBI49
2PcFa5h8JQLL+lSMSOUXSMWl9YQW6fp1a9iZn7RxwKEBoU5F8iqEPCiv04nfSgY2
TBY7EBEhLMz0imzOYlfrd8HPoZsUhWgrvBPHb5pbjcDJSQmLrDqKQoctAGg0rBoy
/z+YhAUK/D2KkAs6vY4riCndRnX3psZSPTpTwGx7YnRagflpuQOhoA0tTPvzGT6K
vlUhFJIFYBWa9bBwbARPQ0CCGDwxvvJX8p77UbbmOd0K7HSZX7ET0bpJhBNexNVl
YNL7PQVHzMN05MJW+kJajAkwoA0YGIL/sFd7Q3/c5bQQp4Y3JFFIBSZiB9nd7evz
j2SB6jAD50hll+OCvMZarlNNOEcbb3dp9+JEv7Fhvrfref7boUOYw5pq0tqi1k0F
mJVFlm0KHveYhjkmwiQcgRdZB+p/dqpWg9vYSoWk4JC5E4Zi9m6lWVFvypDcYvXm
e0uj+T1e01gCWzfw8jqG3ArwPg54J7t70qXUyEnaoyH28RRbu2XTZmRIqYwNtG82
06KBEcUi4RlOr8oNzIkZzPkUyoeXTwVoKz8AVvdgP3iKh1LTH4igRo5d9X6KIgvE
Pqt+urdiEOujEd4v/y4wul7bGYFQEB1Z4P5SMoBi5NZUYHcCA8JPQtRSG3F8adQp
5QFTBbjcDaRsrIdm9AjZj7s9qcKfxC7gp4S3FUoe40UbW/XphJZ6A8co3vdqY/nl
LUobIZjlyLq+d+BgutkZM+XnV3oImABeSQWcQFWUYelzLGc6Qxo+I+PhrmbDVNQ4
8Wd34XiAhIlhSpEMQfU2PIbVp0e1R9s7I9qJCmVRZqyr75RIcY9xChU1zJpyY41l
g2fGZdsadp2pgk6J2c+x28tmUS1T4l3nMKFDoB82omQ4gwF+v47O+4YbghwP+rRD
gPjxsSELNPEcZR8ftZoK3dxcOrH9kCTa9Md/7/v7xmNiiX1S0rJVtI/IKxAkkbpT
vvbeX4P5IzxCoaMR1KCf88+1OhutsYRg1UGRF3DD4GjnQ9nsXoIAhABI4a4bME8w
5Mc+RnSDqWkIXI64Feh/EpvuTS/05/VgWggnAIA416ijQKCiUcXNNYH676K00xrR
3FOsNPho1vVqlKznI7IhQH9F7EGvrqesZeB2m22sprhd8cMCyh2R/BiPdx0q8apx
mhI8Z9imFKMUyG7kfvz6y0Q4qevTY02HYEtI8xPx5rSNHeIQd4o3h4plmzWanoxB
JjPbPy7d49zzAuu8H9imsCTmikaTi26XPlmpO+tPNOhVBbVmz3Pe3YAKoYHs9pX+
vDCudopoi23P9LSqFY7FOfy32GsHIPqVgbPHYFx4dLjkIgIlT22Eu45/fu+9HOBB
MvpBN94CnyfSg8aEo9I5OhyH1bU+DEnDhWvO5kSPcbabu3+aKkTYSjXcQG5eXGmW
/RjKspAMOdRFTaJB2YuV9MSEX+9FSaW4Zy7q9KFOsLVuoofAwrJ8El0XcakmmwYb
7qCRwI9+VmAXLfawJyLet4dh6yKHrU7kYsKcwJh/sUN/QHXcKbp5zFUgpSPdGamI
H/fCuCzr7LSisQU5G1SQLCCKRwPWNDxxwmRuo5M8IHipohx/R5gDXhG70enCh7Xj
kEyRmJvqAoy3sDAHcCYHUk5mXKhjOzAWSTZ7jjUWgVsPZhP0DHrZCqWlWjMgcUVR
EfqzI6rwZZvZ2WXEw4el+C3/+TYsV5SNc4C0GPXMtrqgN5rzE2zLwFEAauUynpjl
jGIOUjAoJ/aTgwCyq3G6mr0WaI1Qn/1gvfbQZuHlxdJLrr4oaOmnEwwFrZUUbC/v
wQeOu/rc2nPzSqsV8298LIPQdG9OKZLNy5B82XHt7AAQ/2r40KJ8744n7KNeNiM4
6zcjYwNtzxKNqPRm5GCxt50JiamF6C//tfVBblzrcNIj4Igmbrsjx5/o/x+43kXv
IJhMbh0CnytFf6dvL94OvMnD25tIf6+r+zPzXRv6LuojLViQotkxm/S/M+NxJa5A
KxvJTloufZDxhprBjWdX3y54BqA5MRSbQnvdTgZJqDRoPEFFHgRmZiM5vwp9DF58
ijtNglgJflWPSY2cxiyjdQvBdlqGy9BSs7QmHbTegikJFXV2yWvuky/F2w2z25TK
63JsakacXDjpiDzCwCk/H+fMhjNra95jpERhVrCtyE6lQvEB0xSiJU7XHWF0nZ4I
xbKUH4CyLdvApSuvXpW835a6GufISISKm55KvxOGXQkpEIAkpQQxiE/t2cbgrBxD
RwYJJpFrs2VHyyJzeKVvMy3sMTqsPwYwUq/4b8wi7emIZrVjmMnJZ6zeQBnBOvXp
R5/b+vPd4FU6+eXfgMMbeEmWKoMq2uHLL4pFYhNwwPc81yxMZ8cmziHkylVzPb3u
nClcwD9TStnDABK7UXBcACjhM4UJHXlWGGK239Wi19YPiwFQ/m0mlWt0kTxRSzEF
FQO6MmrPSTDlPdMYoF1Fdilc+kJ72gI+3p7PUKzZph2tnr41s+VXwmXfdJrFVkC5
Osj8NR7lQbfdu/mAeaX3mvng0MGyxMzXByDAWKFkVp3h3WQG1l/TSzGMn9cjLh5Y
cBxRSGefFTrJPoYjaUlMEHgi16rWIqDNVxmiVBWZjkRqXonq0KMVa3Seah1G0Brp
/vAhxoY8YVf0FRrLXgXHGifh9ODYuSUNR9yMwJ6ZaWt+j1qdvIhZ9xWbi4TrlXL5
KF/fTevJ02+SYS5UC/U9NfpZKeLM6LBNNoL+AI4+XBTzhfHLt3zPur6CVuohzFjs
IdsDcZftaX1M52oBwaJpkbq5m0QSw6WHbZbm688x71GSL+FLN/K58G/M84xJRGDw
qCHukNmVC4m8uabLTvbS6LB+OvVAP23q/9mOmH/dC5MiEJgLChFHWDB6Fgqkxcve
nlipmavCMDB3XlpaD6zZqh5N2jApEVI97j+8v11/V5XgQCPOFJQRthd92XiOTLg/
OIjvBAONM4209VsTOFj9SRXrWsY4I0UtMQjFRjS2E4+D6a9f34PmjHnuT/PhTMYv
QkUOC2L2lH2dac8UafI3GQ7XkKcDkC7Meu4mpNJH3PhCqqqf49KZDg0pP1HFW9hb
BLPem13h0eVq3m7qNxQjfIxXbJn0KP3qpjgtmPO+XQxW06zdg76DNEOMbbwil8i9
TMeLyQY6i8FiRwLv5rhh7v+ntfZ/oVDVpJBAk8hmhj2TfADvLNVOYWOybsXH03+n
Vw+mSUnebv682CCyHfkLKl4e6W5mEPbmF5lCcczDEf2iHKlpqvJmQ8B1dPbgQY+J
FP7sRYWPwyhZOB4h0eUoRNTz9hYaY3wFCEZ1X2FWFgoVgkwhaCpfREPafZlNkDaP
Fv1ULWCkeWBIFTkI73h3ugdtj4egIdLmv1h7PlFmxoshueBbj33j1n4k5PDfPGZ8
NBs9pqsdVs2Y4/+/Vt4u1YeL+CefWN9i1ewKwgypt+l0rDmetWMSvvlOdy5Nw+V8
yqrLi6SafdIZgIgJe7+JKowt/KC5BKfvq9H/IdGv+iccXT3bJbcxpXJl+i/VCyzp
jpJWARrLq+xBVq2MS6DrsEd0QcWRg6yqasYMdBhCRtKeCqxZzzM8EAfC8bkDMK5x
zv8frd13T3H6KnRyfYQ07FJlitFB4o0XeQ0RaiLzqGs6myF80mhXQpkMZWU6k+39
a7GzHjHVyf/qRB+dnY4Te57nTYs7msTMGqhGYQs3mnh71bKeB2X6NRteFYIAhXTm
xKaEwvbbGHofSrCbUy7JYY/3rOWaYbD9NcBCGdDjTAzRBnop3Fz9x6K6Yk7odpx8
d94OaeGlHq5Mw+07yl6Mz7BHQG9/iEGodazCAQGhgBTzJaxrGVOOFho19ZcAqrCR
UDjt9JKSPjqW10SdGo5VqX4kIH8qR7oBKoaqDyq+8T2TbP0a8sZ5/Az9b0wqfTCe
XkGCuR34vwRaxwakdGHsdOPgmf9VBxac/5YWDtfZyop0aIJxohwF/7lOqBF/qJM4
SbLI/EWLpbcnQvpgqDAa2OP6NBjM47i7RDqZfSLLhsqXqUorwGWyVvinDppJGb6z
otAf8MWcwZs/fdZE6rGuEeNQu/BU8Jelkw3I9p63VZGjCTthjcw96H4O2lEa/ozj
JPaIMYqTNIfiSj6MrDbtM3x/rbH1MtiabGRAYizfemCru30VdC4DnvyEYBZlsntg
abgOOQPnBN2lWAe1/qy2nExfGWIvIENZ6aZscpAoYnrfoTBO0t5dP2YY3UF8CjKE
CuXKPMTLWR5d9vAlZsidPhiqDJeNO9yRL+0lJzMY+0Rps1EchPnzL6Mw+9WhB0fu
rlEarig1I6EPRHmT1DRTwTw5CCSKTMNRSTT89F3xNJnp+vrCZkN/0xcYwMMHuqDB
O75Dw0x2dHStj9NqBRiZ5s2G1nyGczn9rZIMH4MoSs9q2ILYXdUmGJKfikksarTE
6PYIp+YXzAGk0FrVtDeys7T26YKDouvsknSPp3qCbMN82Qsk1KwGvqqFK1LByj6Y
dz6b2mVVifHFqF8hYZY0B1rWIS5TkVZF45uiodsvaaLwPa2bVMGgJVmjCDOjH3xq
Df8xjFVszzpvzI6fgcPV/AdpxyjO2rnCMHM8QMKb5zw+fsu6imiNwRuWJ9ebzUD0
7wRTpo2LYfEaiOs0oghUM2hljbTcTuf+xZJbjg3mMJoBwoy4Mvtot4doXPuBHPxn
0ssmY/lQnch8qT5+DgaEv4xXZAl9S6b/zg269vOPPxYUnbETc0+9ppiVB5Se49Ni
Rf+WR67scR1loDoVEpLrkwdlZn0rG+EMYhy+kIKW8jl20oGE0vtSmiUHtNOGvi0i
YgyjwgFJtfWJdwaoYp2nKdwlmky0r66u8E+J+ImA55Uf+sM4VEg6kQLU2k+V5enY
r1H9BtRju6SuPoBld5KXHQqoxY0zJoLG1URkhLORuJv3ntCCGV8xc0VUnhBrwsOP
IyOzHf11kZtR/ZsNF5hzrw3mKAVtbN6sIMVC+vLwvZzgVqsS9NhD2/ZpcEYcnmb/
SYj6OmQfiZWZ9rZIzexIfDE9YqHhoTKM1X/GIUX15mX6LEicuB4Y0BMHy0tNPSfm
Jl/dMwaSwlQ5ImOK0NEmXEX2/MFXc+yGSXc1sJBsfalD9ct/XxeYaWYZTPdF4iut
3ZoEwiM0bHSXyq2wL203VWcQX06v96xG0jyR7kCZr9is5GibmUhE4iU6vxxyh7lk
Iymfxa+5I8qJDgMuP1AzICjBiQODrrkTrxw1sW/vXHQgX+iGkayTB32QjHxY0OM6
HgkR2NUW2jIUwAjrxTxig5Id567MeKyoU2rLzYcGQvcaL81kgy8GPcYulq0jHxtp
NKdZ5yr1bXlVQHs4IfASrNC8AfWebtiJIDy/HN1g89z6cXIZJJXYD16aHPWlFrd+
qBHMlVe1kU/50qD3qhie61KuesiZjicWeN+qOoEia5QBHBh6FVNArllty7vnK0L+
ZsQIQ4mhrwmKD+YLkSA2APLUIJL0+/4rgFBxitpqbBTZ5IfehdzwQiojatZTWMos
TDBorYCTPUmnk/xahglDVq6ijQfJvs6DiRyRuB6s0ChLvNXAF2GG4i1SCy1UfBWF
99JDIyWAoS+bq+theqky+Z8s/uk50fZKLGw2fp8Pg6xPdrdVjE+Q1ib2qs//Qzur
2OzJI8wM8BbIRAZg8xt+dsHPGMwh5mJTv/yJzp7g3vWTGb+Z3ZhKvP3gwiw7i4lq
2ofWbaBxh2Vua1kJyFfYN/iEjWG85LOFJEmQWfVmf+W50IlCgBqSNi3oX9XforY5
krR8S5jlQhir0fAuJIW+nkycthT1h129cskZBYSg95P/gGz5MGbFDPs9nN561Ssl
qH5RVzAM9k5E/v//V0n/DK7Jiid1w6GH/yVnBcLDQAn5ArOAECD8LVqpk0CA06WH
S2rSIAMmG2WX38+teXYxvP4GIGfX/bLplLegIXAbhXyEi7SdD4Yde6CvvD3X4WkK
U9e77IOMyY294NINH7s79ccrIsVN/f7gttSzRfV5nPkhnTopHlpxq9eXifDgqBoK
GOO0msDL4+GBjJaMKu6Vy7CO8/jgYOAMxU6jqV9+qxxKzbdV67ot3YUXHDUBQoOH
M3RZhx5CAwil4JX2bcLZ39/9mAe3odvPnQ0m7t3Ts6Vb/V+meD8/YqlwCNqkdeBs
hugBDoYThU3/k0ws0Q1sc3wz2Cb8a/Lzy2HkjqIoiNSTp8yNeYXmmw/pPs/Noj92
J5gX9+UDu+zlN1ZifQd7htKq3EJoqS554tXgPvhRbjLgL03905wOgj+m9RhtjidD
8jFH9K4LThse8/85zcGStH108H/9eX04+DNGpdSk+R1MOK52PYjDSlvuRrfvbrFF
T7x3XFhzNOP2TmprLO/idroETHsa9UfmQ6+d6HzITTMNs921pU/J5MIsDIKiY/AX
b3pfEyvkWfWm5tsEbtHaBElyicO2vWYEGIyCdP+8Y80Hhu8QzxnqOV0tu1RM7bL+
fh1SbBA6osgZwo8eeUcKDFvHhTs67o5HakbYF08hCGck8uP6bSG53jb0O0x85bdA
ioSEQcz2yLhY2TouUwGCKjHBS3Je9QJ16CvklfsQr/Set3w6c6A7OB/cmuK/xkev
sztv5RpdN3Tqlhsz9jzFPU6LPc6qbGJ2BG7MddjpqhXz1nqiSzUbpgVKdNrbE7ny
VPA+0itGacc/dWJ3Sz/DU9BKDrQC5M3hDgeSb1c+UhdvaM/nwZvAQS8ZVpMulcdk
FsKFIcZ8DQE7AaeaHV5JKRoMeSItSbfv3dvvERv3lxRFBCipLFGe4nY2ogAAygEa
Qyu2bN2gt/OPddqB7PG5OjFm6oYrtp3d/8XE34UWhPuC3HVFk+WbJALqxZLFXomi
09Dw1Fve49n8byqAQE+xZD1MD3bJlsocsyaHUhjq9tGerrLzSAu6Gerwe8i8/HPM
yWLXjDzgsp9oK88qqMT/+jSSyg5tsZdcFPFMGeSIGvJfQKXewzMIxdveSIcNY4QL
cy57eS0E2aEPUePcOL5xXaNnzgUkO8pRqcBUYIdf0j4nDp+zqYcDZTOAU7dmclVg
+lqFeg/2MyeJsgdzRN+qdXVsS/SxkxDghTquodV3VlRXZvj4pg/moVOCSXT6dl6u
hvA9HN+HSQJ/K5fLOHzky3jOZ7CLIU2AMq1wZah/ixXZ/xcsCcxHSEsFpVPNvC33
UrBfJJQIihxPEsfEhl+lxpxLgsHqS8I9YILYHPtEYtMEcFQTXOvOklw+s+eu6xEy
srRvAz2Pxw4D34eYMa5KA/7cKDv4odzNXx87FbAbSmPy0f4F5zmHVGlZCHuVNuuq
uqirDlYHjD1AwrObnW96cpemRcC685om8ATuf95TvPLUO7WwTB8uMSEIxxEsk7QX
Rdhy2l/mhD9+s/I3AYqAl7BQMxp2wbhrKj/et0iJmmYgc3SJPb62+yRjNZt5DKEs
hrEhUIcRRFYVUmx1ycMKEJkFmZwga0+xrwfV5uiAnpgvROCvhG+61yMFy4n2Dt17
Ii8Sh7QGdUh0CjrtoxdvZrFJHKGSktG9McB1FKqz+pHWfu54DBxucg7pT6bARW7M
YiyCRmrYz0sk7R7H/XU63LTNW78CDFbNPbLmVFjrUQcQx+21j/p9ActgqnrGDMJ5
bMxpKTQQxo6imZECizOcfPsqMFQ1tZ3sA4DfQaSywabN54pVAQTkh0QcXH0sKvYD
/wEBZjEqYIhnLgNrSEQiCGSwDA15XqFbSnqJX+cdpk87caNYNzO8IvVKjWYFRIpT
RjnzzIOpWxDExEnuONjPEmIPvmRbOW0ZiEXwBKt0S9JDDWtMExIiSA/2lCa71Rb2
2sXZYLNQXhJNBBOzWDDLFcirKY1Gl0LoxVE7+OLGRT2INoJa067BkRGfOQUOMUms
qLqCivJ8H8wu0DucbjgQSvwzCJU1vPE8SDygBRap1ZRR/zwuCazbkT5TzJnNu6sA
SPEXlHimh3HWEf6u18DNjeZqJtC9GyvdwXb7k/v3JN/InMQ4imfpr3CruWGc4oyp
+m/aGl7UhcAE5UqZf1cnTQTl5sI3oqLVJjOn4LfPxFUy/kR+ZUurt19z2Oo8B01a
ZLDX+M5ua/LSchaTTZmGSUaOWc3IQNx7RY1TjzWsUHd2d+lbMDKhxBj3rWujyhnX
9AwEdbY+rZC7dxX6J7zeiHp/JG3YfKjCm0ovMj+K1x2xdVxSTgkjsOHWM8wE2P+H
6zpnWByPvOHQmi1NRPrMG9KPZIxzgfqSXFCmodFwKB75dMxpbIhg2OL2wP34vu0l
twhPtCrq0vUmWaXckdBA30y0WYI4wBjvW6my2AhRCnQ/AlJrE1QBd5a4Ghxdad3X
8od0VcazggawI6VtzPx4cIa9TefyFO9Orlm6J4a9iDdejUsxXyBEXThfTPlvioH0
6b4NRBkYgCmMW/oVgdr0h4iIf71SSLshZlzzYJUsSR+q5MkB6gzvAAs4+D5DAiAV
uWPTQ06ltJok/+zlbJJPEiVoDU6LAzX8zoa2xp5UaRxWQpyITuN7aq+KcRMXcdxh
cLW4Q+wgUSym5HqsTUMi2GKnuYAJR4Bnp1cRXVcw5uQN5K8mnSxs7TIK8WONOHcw
54rTTJR5LOC+Du37hVfWTqWEr0t1oKcwJ8dRhsi3rMPxxyNzfeWxDPyXmza3fcDx
vCQbvQJs02o1+2gy79JLWMKzi6f2dcjHXbaDUYxAEavlCtjZs7l04OE+6AtgR6JK
MdcNRR5B2bt/L1og9xf4HT4p2cHiKfDqcAiTVo1/PDr9py8o1gBuLYgSsbW4B4Wq
z97ASFt1LQkGHnf2t3MYN9YADKqM4aB+LV1JKlLRXhq7ZUhBOVn0lv2n5Waso6nc
maXu7MWMkV/CF12sWCdE81ITM7igMjH4jhqTr3wstAozUAmE+pU+fgDvQFi1h0Rl
ho2sxmxFwQoIpE2+lYCDnL3fGg9MWGObKl/YdtUiPKuKqtCqHYAZ92lZwF9X6XFl
xQT2OlDx2jNosLnDrwr0s8ZdSTikwbeFOqMJW5fDU0FnUQ9uv6eTmgL+JmiJP6wq
6iyGdpKDbjZp0tvCRghA6xarf/D7sdonOuBBKY97+/wgX/ZIHU7H1kun8dZ/PBJZ
jGU1lPcK/3n2MvWtoSBQ8AQuzZi8afAF3fdMZF7ess3xI6QfAzHlO0U7BnGwSrnB
kAw6/YfLX79FJ+OQW7qgEe49kIaNAsDG6SJeaSEHdJXt+zT4k1liZoJCVe1Ly449
TaQ6ZGP9JYY76IG+hQ0UoyLo+0wd8rSrWllWMF+Dc43GFD9Nm+n35UbwAgqreGOP
p0hyTK6/OkfYhNJJHBD5NqAtwncS9YOcHhEBgSUsSVf2Bjkkg81FOuj/R1eUfYog
v5UfVU5mOxPbRmNHXDZyJECkvtCh+fmjhl/bYfdqyhsBMAm7AmMuQB4N2Imryjee
BS0GLFpaRgFs5KpntSVUA0JX7+YnCc+G8jxmtyLVwIne+5QMIUrvdcirgMY/jqvE
KE6YvSImKajn+ffRWWAfwe0amTQpo1fl6MDjtU4lnD7+KWx1TJsrCdeyijWlR98g
5G/K4U44b35mI+JHN8c4ubpj5VbtdEA8JbwJGxEQQwTrkRajNCX6FuSDVKJs+f50
3prP0sisbqzYfKuJqxzL4xvtr0dmizVs9oFWy9JE8mBDfKjvvQTgLQE1s8nmHHvc
9yQOT/sqNsmNaFiwRk1wURVH0ZvXvFQPMqhFlicFrKS5ZYZ8dbxDuvSwHlFIbO4k
d5tqRtf/49S7Nfe8oqCHJ4gx19qEXBF1Xo5L6rpKXpnvOr4yeFhrUDqe6RHzz88m
fFfvCtjA7IPoQhy0XKszWKIJRbvGoh41TEEXgSxUQ3NeE5/2tEW+cMGXyVbRoYf1
OjCRpuLWXc1ZjTFITjDngPUpfxgRQ2HPp6y1J8FGT76Z98cU+Yehl7rZtDYvUo7L
LRohG6q9hAx+ZAyE/RePh4QVBWDcBQhToDN/wVeI6uFHGsxHixtJQZpaD6lbnoLW
t9eB5AxHBQhx+h1EwORBSuaTDmrgt1to/Yx12kSwZmZ2RED/W0XyU1IDGg3saZ8s
DplOjRkkmPP0nq4U6smQGKV16lay67hNNHFNqVjFb7GbtpWxmdEZ/YINd6q2Jozr
qRZXRaee9j60OrUHWtcTjksoK1K8ae1qzRP7qdsKMUllypoafNIKWGOTME4iPyZ+
8dgguE740sJc4kfvMZcI8ntg0YhvZiAuMd3ZS/V4m28kNqn3Qxr4Umo6/LC1cMFz
ebJOhOnRUSIdebssUl6nD5jHbabNOd5GwlsNcsOr2Bltw1DvTQxZ7IjZZUQMtZji
a+Jm9Yq3+US6/CVBOuKF8QMOaNjdcLAvliJq8M5XVA6iYD2DgWYA8ZwFKfeTxZW1
woJCJra3vc1HfjHrCWxG29ft84aUdT54PUvJaz2cedIO+dV3d/AkN3ZS1Mej1ka6
E66RkyxcM0kWn+NAvYWRsX2Vk/qgBr2bWv0Wo0BrHf/EJzltodMhu8aYJEc/6MUA
80Dfpqs/besADl34Tptw+GLu96dcVxJAEj+z8nA6YgFC1JHgmMYsWEz9QRzTiub1
b9zYas/fm3xY+EaCnPktR7iR8m3BP3FmbV5EP18pXf314LV+7M+/q3aJgmTZ+N+a
xjE2yIixne1VLOt2STOc0zsfNtzvHv/HxyGSKuq+yJxiWvxmGsFtJYo6XjV3nP5l
N0CtcABamvSRx5BhciGJwIHqD3Ot/U93rE7xnvFJL4dMDK1q6wes1og4SvVg8KdJ
/2ROm6gHqkQb/NMY5ur3rElmVJbg9qY/7Rek9pBu0wJML+uszJxgwbVUsbC/RC7P
tAou48M6mdBoyIpHNuP2E94ibjhc/1dXTtqo6jjQO7zDMFa5ldT7c7kq1GJYjm6M
tTHjR7tM6rHlt50Ye1wTFOKwCGfw88NJ7M1pJlySWhXEtifwaOtgJwMbmE2xeWUU
WZZ4+mg37vSjNDB5+gfuLSy8ThNwaD+DMGTorENj6Ckalx7Jogu7cnuDOw7wVE79
Of/LWJWt0D3C9EkkngaTfHGNBYKm5DRXbPfLfzNlMPRlsabn5YWTyuNleM7ZDxXK
Sz9oQvFoFELWJ/Nlpzy0GPOwPEz6Dq67YHZ1a6PiVnAq+i67YdlsVyNzE+Wjc6LS
CDDkXVGd+fgh49BfQ3YYZk1mHUVK0tapD2jNa1PUJbFJ9hhUoYPOLNtAjRVzM7sl
VyQ2HRgGvaN/EHR3GhYBTBrVzIde3pMqenQ+ttY4Llr9E32vD9QCzsvORbonJv0n
DEQAZ1lA+J+kUy2zKPB+68gihMOJN+M2LwGwGCPXpIY7Rx7YrzeIZblFdzSYjl1D
q3KdYFvTq2DWDPj3i7393Xreg1YFfCGb4Nf2SlsdEtUnP5S85g8ny67n+62hp/sQ
LRnSApohAggB8PiIjv358w/kJfRs7vLU567YQ7x1sj/pDGYDcRPd3L/R/NGjojkv
Jo2fqX4LUXy9UL6ne2czmC1oSmaOIEpFWOvH+oWTYg1KGUonBsTZiLH3SvvkJTHN
sbqVzHgeQre+vyrRoXu+43jxrh8ehMOVsYFXFQ9YkZ/RBKVe1b0t41Fs4RrR4yCG
fldu3w0ZSj1j+poomgyrR/LDXCqlQOjOVPybGyx8q5/Dqf7vMnLvgnHA9MBIrCKl
6KC0I03EM/8xW4oZ7beFQ+g0UaZCqtGmPdvWGoAGVXVsawchhDINK+B1PoKM7WYL
ssfm+AY72mnk/3ku/zvimovdBpNyCmN4b4aOpAvlZuZKp2ACoK69N2rlBhdJ25t7
7Fl36U140PAvLXf0vQrqyFh0imLTW3nKvyTOKAwwkeBwmiYP6r3A9BeUNtYH1ACN
XJ0GSCXClLYLlVdSoO/ZNjRI3jmeY765DEDVg/TgVra8kiYSdGGbwzY5DlJoZcW9
kOWt6X2lEtKZ12nHwWCMPjIqSMyNTxgR2aKYMKnWsru4zzAVkgx0MDFslDlID31T
KgSvD4sjT3vJNdBYU+VA0AqojwE15Z/+0t5pKmIq+oVYQtH365zSDf1RjiguHoxv
f4FWJokl/wm9UMcFZ/77SvfD+wM8HI6NrD1OQEovhqvFp3WHN1jyub28AnNTPlF9
Or78ilBVyvUqpxGvBy2p/lTlYuLnd5hBfDVvCqGPWdDfjbH9KgQulRypwBhN6Bfu
x+6VyGMADz3kZQ/Q8KoMN8bqrs8/7/5frzWVrfZbmUCp1cBwjc0sprOPAr9XklB6
WnJmxcbKAVSFlQ2n7LO3u6xR1tZZigmIQicsbN/YSIQiB0JKlSLN0LoeXMM+3m68
GoOFwmCgIaKyFQCl1GqI7LjSGwoaBODcXDhxt9CoXKIfA/EKSAiTl72u97Up5Sfl
DYbZI85p/icM7XiIgcO/bvjncVDBAvXYm+sMVnohYLedIfP/fDhm8/7nI8vJnZW3
ewQVSF6nehf+J6PeThLuuPu+vE4gn3mY7XC/+sPcLIPR7BJmjMW0Is8wljq8LXel
dVluJjDHGgbZMSqeFgihiGkpoOGuuz0X1IyQOr2OXFe/pbJsngnGwbEOKb19M5yM
CpdCaD0R2pC3d0yrHZWe+KAxaxsNePXFgibGYu4WHTasMTIveMWY4bJT9pOBgJcu
Hjfk/i0wCgW0dMBVMyaBSrYF+iSavfgSVmP8YfC0jfcAoYxJsizIxVQ0KispmoMc
Xtx8YVHqpF5GmpxHd24MU/SVyLNkt+muI4SZgRIKlH2nVafYo/tKazE4Ypwm+DSN
xL2+26w+KxA7igPe9ZBw86FgFze5xspIczYC6P0mznhvtQ3l0GMpDn7fAgv6ALrU
ddEGy0f3s84OOtrbwLDORBroeXcSnIyxIDpNKRZC77R5UJA8ZbSiTCgzyyGDq2jY
tN1nxEqCweTtmh9X9cVljKyeQS/vO/YR6R6oUlRFZfr82aN83xi7xung+/ATjK75
MuTRLB7x9i6Ndn5L44teHTiKwS2C5hHkyvcGplIIo1qeMTekMJLAnD3MSC1Ngsaw
AytGq+gINhBPRLUSQGZxbvn9rd4l3Yz9Eo549CsiyCDfGNRVOa3ZWxxvR7AX2Zc0
I6KjzwyNktQy9v4fG/DexR4nAfDtuSMxFeURPQmAeXy0sGW6JrFvBYHsEGzFydmD
VK/XkfxabMS0d2zKssc9FQPAObUG1FBMjbn4gl2dj60LgHzsLAVfclJ/fIoyVSVU
Ok5JpSFy8k9xF/MuW/1QZBAM0e8Vo3yy4RfqoMiZSmt0I6LS/jdW1reG6muDPuVt
a0nuNvBZzVcnwQTSDq6so3D0c+LIFp5aYCAYfAhZozA2o9v+K6LnDdV6JymQHNcY
jixa1axo70nFSc+2CkHPLoLGarkEwTnh+N6LICMGZW1ospxLwv/lwgg/9EEEzJky
zw1Zz8UnC4bNrEB/Xhf/RbJ19M6O03uzZcQjOLpFBitz5nJTfriS/e7H21vv4O9p
gyfUWvLaS2tXiaBUgAsCFbJKrZCkXwcJOBgdAPc2DiVPkvZVydGLl4bqFSKCooNa
18mnymUwfgJxNOAzU6+XFzlx6/fRxetDpobdQCK4B/ymz95H3OYhqrUhwgS4zwVo
1E07PVdgKQyHXn2opyRYp37QTRLxWailxP+0N6BfXUfaW7eZilSPsOxyUECJas03
gyVfnLWSd0vpR5/vh0Hrw2fAGvVjgJA/4nu2hoDPaLwJg+EiJI3wNAjGX/O2DvKv
EpMEms0JuD8pboKIQHCqBsSCZUW+WBEBakeRMQxM3boKWt23ARRvRsmJe4oR2uGf
euTMIQyuA/cx4jkYlcgsKC8KNOObU384FS3LbQIdA+5/Gn7uCMt8fHPTdJWMaD7L
Xc14arhRk+QzqXzJLdeHbw4D86c84ncr5xt17ylDjvWrlOrluPZQLu4/tdxeC8Ys
ZOGFwUm7/Axj9u+fbVye+6qf6/618b4UGOhxVEFX22CvW4I7dGo2+g6uDKmossAG
K/VVZ4oNfuYeA8ZACjEVCIiZSD0+3KNotMkeeRlhLie8N1wU8Utu4YU/PawB7K0A
hQSYErq1HtveUBy/XXlUaVjqT79xLmRgVLWgz4OLd5axF0JN40fvtzdElcD4+7o3
ZwzqrluJRf/tfeyoXNQOX9XkDJD62cPYuLV1ZE7Tdk0Rld2xQzCjGQ/Xd/aLLjvE
oPUptVdvDBsPdeJ7ThADiS2J2JTH81scP9l5igAQ91Mlos//RTBRDfucKwpTc0Hv
EPGjgv90M2pPgPJVru7NhGYDKAx6AR7JYKnPLnRm0yexMtykkv4GtiqfMRN8rE0a
zaJYybCcvNRyQK+e78Ns7TeX/jDBpZAMB3HiDAAqqIcMVZuzXqrn7a4CBFU9Km2c
cpNZPJkfUXKaK/HJAlwy2GNI0Av8vjy23SczPbK6JShOMvi8skOCJZiiy7ly/+dY
dKZHrQPFXVt1VLNq8FB75ltgmQ87uLpAthG3PEo6aZf+J3aNUWQMLjURvr8Z0ZmT
mTwwReulxPh0nvjyIgTKzS/Q/uzIuSDvoGwLI7P6KjrHEpXseNNR3VXKw9rUdQzF
aWSeKjJShkTk2ebkpakSGuzxuaUzwTMXZxG+DRNF9HIiV93iq8WuyjQ0fFiPpFw+
eEowk9xpJ6ynFx6loyTi0IhSJ5brlLMifW8W1jal7ksVMKIvNxRW9c8f/9dulDUC
0PGuf1LUt7NgitQPQ7lZCVREztUtHohSrQHA7DyD7zhoRTF0a3I19WzALW4K+PcK
h7z4rRox/LCaySUHQzIOe15LkNxTgtRDJDPZ/F2cFRqBRRz9JPMctsOrhhAkt5UX
WdWIpejJF8dr+HVTbN/XoqjR8QSja69r7ItDb4oNi0jyaTrSMTNEqpNhq1ny8v5E
fGWxLOQoYn/N3j8cN+IgmaQsJKo026M2MCXfRVzK7JAqRWenCtQz+EANXgYm/LJW
SFeGEvIxmiaTs2jOx/r57DK5qubpXzWv0tVfg2HcgyfCK+SS2l/XiM1ucDSQcyvq
Uqzwej6DoPjALBEyvPlkBe5HPNnrTH5sIW/SE92jRJhpLBgY3ugYt5UTB0IIQdAf
Qhv6EXbAHYfodO72oJQDyRmnkbHEiEnjD4/P59vhbjMP0oMQtVGu2AC97Hz1eIXZ
rqSiK4ybwBZW27/Hykffp3t6iAydzqN1j5p5WeJigUq5atOLzbOgrIJ/pQadRPv0
QFpqona0REzbxLTQeEfmGMtAGm2y5xEqXZu/KeyXDkHXY+2zhSq42M0U2r/xfh2n
TtkLidUUijaqussyDLT3oZ1TTTVe4sk3uzomrgf/EnUCpirunUgJpz95EHwfSDX0
Ofa6y7GDX5lKzQ8/10xXMWDgj1wXq/CB3fXCEBWRXzdZ3pVKOlQZTWIHRf+RFJth
aB+ibusXaFzT7aakW7F82a8yZ5M3gcOuWfaU5BqFwzmLlH6Kjd37JbV/5+n+OFjK
oLAcD7HMV0yJFNjrbIM/4afn9RdPT1DGHlZ2+kKj9gP1SNnPzoBn6gHKLnC8mEHC
uoIaP6WKTU2/kSokWspRG1bG+8+lG0sYy4agH/GuPYCOi8NOYYVUXwCyHphUtCMk
mMMTe874jhqf8r3ZI11axNp92dSWas6u/Se5gIjjgvBBwBjavJpmh3ipIIcCjHlL
2DTd7uMobTmHEEjnyuhvUrwwPZqUWO1rikTddvRNX1iH/LO9OEvPCECJKe4lFoCx
/nHH9Nd0jix9dFbuirGJSWGu5LokQTAe1OHKdwZVTowa7zHjfq4s58m1u8GgAA9C
QIlIsPV2w1w6+Mwz3vv5BOJ3NTOjE24e/bphGLPzIKya7Zi9DesiIoDqqBPqb+tG
/kleAgMvJiGEd7Q6y3OVDgBUdWIkmtBKlNPeTinOI5925pg2fvT7C0HUVa9e6Ol1
AsxZFRkhuPTiGDadIXu0nS6d3/T+KVNzXRnD2EPAb8Dg1bgcbQSHQN22rttqVW78
13H2YTbv84CE/IxASF8l6csPmCfY4rXqfPe4DX1FW804ySUCFnUH8xr26q5Ih4GB
lAEduWWvvyqzZzlACdR4JnkqmZ/stN8tDNOYYs88VGxpskS+82331ksVpIe52FsQ
h4Js74TzasZ8Zfyn5IDYm6BwEDZWYEN2b3CoRACRrbxJaC8y7oFnZRg+aS17i1P6
BQxucCefYdrmwpdTJWUROJcwMqCepf84RFbTOLEeCqGTFUJJsbqYRr9jUogEi8ir
/+FDS6R9OsQmEUi5IRF8FNhyTrsFQjEKjiI/6bSWAUdjSEeqMonTR9ZIa422VJFG
NDu7VPhc7dmLWIP7MUyzLmer7afbL99T8CCzbVTNgD212USI7MgN5wFGqCSPKaYn
wlQEfzDCdKIfvMaPWw9FZZiGC+mYPuYhtkOuip4vtqo0jR9VQbsUOsAETNdJVt6s
FPLxXGr4ocxBUOWpEXZmwc6vfUMmTdJ0ehn6+rIJhh8kzZzFFU809rCgqDeat6Mc
U2VfHclmhZe9HD2Ey3xvc0yBDUVttjPIrBvp2vidYO2Y18wD3QbjbauVluBYwVzY
HKMao4+PlK5q7xzrluwnCFu0t/i6BZ6D9jgtBvaCkHKAJ8s6bTsJoMzjSwY6GUke
mIsN4p9rBRnw3i5zp/cqQZeCNkHVWAU30L0NQp7ilPzw4+/nsHeuIU5g5ShuSXVP
gZSHwp2wjjsMJOJOcj9KSfQaUtiMLYTD+u9mH0bdCDvw1SNwDwLm906LJfeMy7Sz
ZQBUX3SW9lp14Rb1cBvF7m1b7lNNnU3elC0+2/+06sy76s75rOngJPBjBz5uS8OZ
epRUVxJUj/96X05k+otYDb6V2iX2jNfj3Akvon0vxxI85FN0fZTnWGeFjQWKz5En
GxBufiMqy5F1T8+zjf4BHABmvDHJUew0yqZGVGpmTpf4kL0vRJJtrE9N1Bshz7PO
4piiCm6pYE/DLKCayOJDpKIhn9MLWD6DDH4ITdzyX4I4tFjsJ3BuMBt0Sif0yQZv
+dUrqyDUQWo+3T0vD9XCS5Rbt5tgy4xE9UzdG5DDzNCylbHFqc5buUpZhMziym7j
kWnzTUnWNfO71Qsawn03yyUXFumBRRZBrJIour25mLtdvzPzYSJJnTl80/2IlPE4
QWnA0DeCI99qzKoOVu/NZRedr4Tyke7vr0fHzKhSgXigogyCVcxExLzJDfj3LdFL
Xvyf4AnLVSWUc5j6laVLtUQKl77D1iA1TUp7AtZaPTM4izWqAM90AlF1f6W0w4Dt
ZF9TBX7GZG+R/7WxhEKAwtk3ONVc6/1E6NzZXfAGyX41r/Wo4pZ4Rnrr0PwGkab7
ydzimQhFk+yy4X66B6SeoDQ1NCKKtvBrtJEfFdng7F8yLCsvTBZTM9IzAUq7i6PT
kMLgEZJvIvTiPvIYDSlJ+ktxy/KM89wg9GHH7kbTcu7HuA4/80Yhw6YllQpBBkvh
hnS8IxdgWh85xqrtgl9EfCWJez8IpspXl/Agky9BlHj+LMZCyObjMv/slFKi6P0e
6DR5R2vX3WhN50qEWacA9jJoITb6GkSUVdjfQC7fdO9pfStqM8diLAss7EM3PkFc
sO/ya/jcz7jd2Zln28u9zGgmD6Q8IDYACzHCxN18eXnzkBnnBh2GEvohBpatDKI2
Q1naCRxcMfUaeZXgrTCYyMOrTvvMkccK6qQsBWisxf9oHunTiZG2TA+y5gVQFW3s
Q2kwfrbiWhXyfcpuGOrnqSUVXDkMItuYA/ik1WFK5ASMOEfnDPSKavjCbpjUilDC
JSjDaZjXdW1IEXeZH93CRbxIJ6nE5atuoryCG2eXb6sWBDpZ+qMGVISpyUGSlCq8
tsJpqDPUz/zXRlhjc5Phh59fUuxjoS+wg60GRerwrZv+0KPFqe8lp+S9R/B+uCEy
n5m7oxw+E36DWBT991hvBCUWNsYzvcioy+Pt6CFhNzYunmXh3ijxsZgFi+sItaYS
tMxdWmZmc2CJ+UtPfwB/nU6CvTqQjLOuYvrCcACtwCe4+Y1vqoAEgKTb+NHo6HYy
Eo6qyqDuNxR3/l26FiAM9mQdh6lIUbwbF9IXBspBlujjyn9qtdkBV1riwyjpUol8
b3qvqc2UexqnpiWg81PaKlec2bPXSCTwc9PAetpUMcPTxozf6Qs98RcTiLk5kGkM
S5tIjAItK44p4ozMzGzyZP6rt1mPHbnq66XLrJvFeUsLF+clPvlUMaL8gaxVm1pC
88HN0T7k1wp3rsURbT8GIrX1RWwtDr25cfw7ijG4KjyVTv4RFoutTw+x6flwpwMJ
Rk4LWmPTPZ6YA/CxQE8kKYXKtnVzUH+RH5QFzPmomem4IkG6QIKB73zm5W3XRsvg
sc4eKPY3EPKWSf4f9mtNFR7RHjTd/1o2rCqpsdheCW5hFHJtHgiAlFpxzeodfgrq
gHMk1y7uvkS/dWwbLnRCqTb9ZRcSRPcKtpG2Nldl/qrq4vcPETCnlVYgivGLMzzg
SClzOTOvfcRjvfp2YyK6VCnQzW9JESjkt9hiK83+Mv+1eL2SqICetgJAcYS4qLbk
52/eB0Tzxd1Nsx6H/OuTgrTD6nqTcEC2JfStalx3n/B416Hcjw6Gcdah81ZEWaey
Dux24YP1QfKTtm19qSVyVPJ1rJ9BcFxQR8peR3KwOls1ByTE0zfBr+Pu2ftcehz8
rLTb3KA62yXlk28Hvd+lclqcFT/glhTJjVr4u9pwOevqDMo71gwi4dqVtfcP/LQt
WEiB3n5rKLCbyU8a+UTXUaIsiU5zG3fKRQmm89uLK50ShGJyWM5gSUF6l2uMxaq+
vOfhwCd9U3F4MD8KsEXyxTY/XTd/DEmXtwhJUwGdnmfIGv4FqoeN4YGfwB9LD7eW
K4HBVNccJFwV/SLqb093PKqmWnYVL2X8jIod9125Yj4npNP7uOVswKafnmDkUMy6
eygT5YLPRjoISTZbTp/JPKlApBpczhXLSws9oNEMF6dvItavEUeo8j/vazLy4ujJ
3oKf74VZ0W+NxWNMt4XUxeHeNH8AKeTKyR12f7V6zcd4zwflvKiUU7aKuq3THQM1
DHJ/HLXRE/AQFeD7Tn9eVNo/V9Izlemo2JyXoTBZEByD8/kFjWx3KkSSu2Vbp8oB
MBOJjAjsCnJzlHqoXF+QIpvuh9fJ3c8xu3Kf5LBD8ARIvGAaHw4yGrfa1aBtbyQl
bZ7Ds2mOS9+TGGY7rxKvp50DzMAA7ERHSZkw/Ok0sDP4CxPItqD3b6Zm+F6JGdtr
uMklN2nBFPPBK4Gmgqv04gJWEsgf0q/qwouu8xJkK25Du6/13vGCBt84ES5qozVq
L5FnfeRZzcoQudmO3bOnLOOHAzIVOkBJD4HcayKkC5MthTcqHzirPtGeRc7X5bqV
UAddT7xhbDlMU7Gvu8uiVqd5pUvpte0y/VyJBQc+ZlQ4p2ElEsfAtU/5Xu+3nmaS
HBV7RJil5fpIKtM+0qm67KQ41+pu+UMs/2IgfHEbEqemAG58hPlQM89doEzl8z7u
YvUi7sjqXnIvChfZmHXzTEySQqg8dF/E6pE7X+0nMYo95DbMvWWK9X5zA56plzFx
OgLPW6L3QFtujVhaSNBoGB6bW3TS/YPV2SBkezoytOLvpfPK8HhmQCz68PdAslwA
zXB+i6r0x1Yy+387KDeDEVLuuc5fUadwD3MQBO0n8fLoVc7GKq/qUI3AUsvVx+kP
57z6nitzMrH1M7JGleaejfKXezjMvOH5quOuDdjUxXASZf3w4lrP9WO1sNRGPi9b
SUggWjtc3fsi+VD4NqPuz2VAp0XRNW9eZdT+9CXpqTPGpWkRqQFfzqClHWhS6xFG
GU9jNosgJX9PhI/mSZrgjGvIPVogm7SrDzuDICdgorXnkoqmWHRmb+udCprmJAAI
IBvnd79HKvtYz5k1FdTU70DC7t84bGdL1o742HIKtQj3z2F+qgdzWHpFuLMgF1NV
Egw/eYq6L+iC/ut2QTZqiJqj7LhoR690qCBgVT9OwJfylGBAZBNRU+EFnyVCjaB9
lc5h+vsiG4fdlw7bkfM7DM9eHHFAHNM/zX6U0nz+cWnGIYZW2k8bfGfyQ+bZuAw8
eh/YcHg3E7frM1kTRkVwGs93Z1Rn2ndIiP7NRt93e4MZM5x74CSVs80l+BpA335V
+g9WhTdZz43RSdl/Xg9C1ntnK2pgJaF8M+OOdv6tMsJhczdcQ5XLEqyTZyAKlrju
XNc0Hg4tOIlMchAfOxJeJToH6p7S5Epa6kieU6/2A9cOSEoo6E6+EFX9d8gyFMLi
jjX5pJjBPXcJZwj5owkTQule5mz0Uq5JoNW4f/0eUK7QR8n5GcrpIeSA37W/V2I6
35ws5hLopPPH3UfmlNPmm6JFtC2SosFnCptH/1P023OKDeKu1zpNAmOjBfQUJzJH
UHCtso2XmsLlqyhw6AzTcR2jNMul+e786yhR4/QECZY0/aOhvSN3x57KwA5MaBpY
dZBNrKIDe7MpqBOTvHiuO+Fq9pid9adO07If65Rbr72CL49apaM6aFymeoMraSV4
ZQJUyEhyI7eYnyOfGF3M0A0SlZnut8j4RUH3pqybos0NJJF/N6G2WuHfmhW18z7v
9pp9w8qCj9fIBl+WJ0KbvZdu63GDx9yBYK8NBsYZ2pV74lzQijDAI+MxejE5sqop
sn+VFB1LAVfkcfmImNW34V64Bo/DO49syv9Pc+LtksECZCJCv7VzW9JOVIFw4QRQ
GFcfCTz/7k2WfkP4EVlRgYqW22dkucOOFQQDr05AFyrZa4cR0ijIzB4xxfS6/QHC
TgfEUf+jI2I9aBXCT2cDV2oZKpE3zPIb/wpVWClltRpzLpIfGmXPNOfTtg0taVI3
GeUnyt4c71djKDISCeGSyUCrk8ihXj20TSeXV847a7pmn4dzNE+LrutyciVPjXBo
yvFBqoFRNCuWteT8hM1EEYD3CZ4xdQpNzvzX2Z10+cNlk5hkZ0hUfpKgb8N7KMgH
HsjDv5Y3XSfi+O77/OQ3KGOT4Sc/SOOAPDdAnvrwIs++l8H9U/qCNleP5xHlRvv3
JOV+2ROfjYuQ2Q6jUrZBqTv/vBeR0qv5i1h39YoEIbahaSXFZfL8p88HQZbMXDrL
io4YxtqDCgjytPANuoh33uGDCR1sV72/eZGBLNCMXasbAGII1wLMRvu/pA31AoHO
tbDsdFpkwwvVFpctN9lT6oYm+VTlC8Flur23LW2WGrdI00Jn/gWyQwfhLeHnOQij
//+YFk1QsayuLDRv4QdIJE5QkOSx1Ph6aJsuoJeowBJfz0YWZx3GSw8kjucq/cdV
gaemuihmAwiXqQp+knkKJZ65i7k8bai06FqxA+FHA3DYLSiQeVjBqjzAhg7quHro
hElirrbdVcupURov3FR5bqNyVL6EDXVwlOYml5g3TP+P5lAbS+vCjhSm5Mhk+GOu
X2SrCURdxPFXiziUh5vk2DEKVFNZY8lSDxAiBsv8abgk9oUiFLExgKb9AkkHdQ9a
aNYZmk7fBhQqkFmuoHAFLi5ETX41jeSTLv29Ojry4mvAC43gouGJsQlNyLc6qZFP
uc7DtLZ8Cuvg/sGIM4k/INdJNwM5Ic7zqBYDN1R0sb/u5wKOBqXaxi19C+sLpziP
Eb9nFZyhdv7t2Nib2jR+gjAD05XNecK82UikAMlspC2nMHCVnFBBxwmARjC7/ASk
WCDW4WnRzu46mJHRdyjivTEd/HgdbXIIWIVFiGyTdwk5TPHdod53qfei3ARhbrxc
2ImmMWg+JRekkEdYJI2TUb5p0Q6g/HpPi7lLM27T6970gc1XERvqDBNEAu1hjBDm
3MefzXI5gH43ebBEdI3vVZVxLmGJZE1b9mqjJPJ3wJc3kfh2zFOaIT/SqvgWgZDJ
U+swY3mlyV1T8FGplMSsrfIy+wNnmwyK5EAC+dM6+d2zor5Ymrj7SZvOp4W2c+b4
VBCQ+MQX8km/f7pdeDOPQhjINBhDo/M9/21b38GfySDDezfGkSDhiBYGB2iztQAF
H44JXr3UqAvosoHIxGAI3ZQmsBS+D4Bdtw8aP1OoDcM0M8zNT39AivFFk06QtYGv
TewUWwsf6J2Ok7rEIzN5f0u/GrfaSdRoSCEv+EILu7qH9ctA4MO4GT4hAt5yzI7/
5+DPIB0hpMBN16uGTYsumhw5uFtzp10DSjnp4QU3/ypX/aQzbrQYkZIJRYFmGAkj
L9e7ul2weEt2yd7OL4D/5hPPyDTy634Yiix4QZeJS9dHaxZbD3/Fgb4AmkIt8tzp
2myoI6SMp7hgb5DsVCYYNzW2PZvqzhjhUZyjliHf5pjyQr+ucvveCoNjlZnTmNw9
B7W8u7TXieW4j++YpKGsspbAHTS1fu9YhvQ7WjjrS1FSCq9gxHtZ6B4KtJf1+REG
DOwak3O7SE3E61TbZemaWGNexsyBmPOS3FECJItKO05/HLtG/Csu4vGMiLOK8vsR
y37wzapxqr15TOiVIiAODVrHJ6QrMmrHlm0oseR+e+0/3xius2ZpXqHpnowFBkjE
3tu3CKNgdaKzB7TxBBjX69EAShWXfpcb4wmLZpKZRC1qkKcUL/qp2JYMZHJgU3/u
6hGde3Ib6YhkFOXkR+J3nUoONK09+TqbMZFUD0j3ukoAw1h3CkhFegZhX66rqkMm
0602kIe5XD6Cu78sfb74Kk9a7WwWuPdA5iPJfukb0c9EyqXPJZdgaPaAEMuMyYFq
ND+xorC3p2gWO9zvaqfXzfvSD4r75WZS3WYdZar4HfynJb/ExASvfBI/EGm8HKgw
ArIbKAd1anyaFx1rfiUO5aB2DI86rJXaLd+oxtgQq0l/Z4rkFNLZygZ1EsSQdqoJ
syXrcF84IAGs4hltyWQe2hu5e/hLYW2kv5AI3pHEpawq2RSbdhRGkLxsMlx3ybXN
hBMLTRhl95OCdDuXut4P97yJEXTB0jEGF13Ith4KVptvd7XKhcikF0hAL/A7J1p5
O6t8g9vGdGG6BpjpROfMDI3IpVxs53PHhEZdMH9LCvM9KbKCNMusmPdD/1bJmy4l
wUGjDhJHFPc9FrBlcEnvTr5AHUPmVWptqDXiOwvRTfU4WVTh7cqcQQ+YKio2CDVD
xtWHjcxMhVgIgbwuTmQhevESCXOkqjMr9eP9gd/0pRKusTumX9nxlglgYV93e6wy
hTcpvQAa7D58A0MyqIpVfa7aX4ZlYQGuHarMe5q09ZJi/nxY8B7S9/YulLEaUp7q
YKlhh+iLgjUkeMpT9TuicAemPeJh2wjlMIAWuMorevBtjhWGDeDsd5ZlbgbOcE+T
dogaPUzRysFi3jQ2QLaQbT3VkIDPgh8rNL732E40R+JjhoT5D0L4wJEvBoks+M7N
qytDyly+tjPNxOUXQKxN8JsQDzZL8tbQKCaqJPh0NNSRfKEDEQYEbecyTsl9OroO
WZFl9LSpq0aF3FIW2JKE6YtRRUxFqrdPVoqlxsJRQYRGPMKz5zmfOKZ8/Fkr3jAq
PzmJxtIx48PfjHCQotYxsf7blJajBzLsUYmKVAibF0YCiGgwFFCeUC6xRsMTJLcM
WEP0V+mCD3aYgQPzBEJwSVDRo5AWu4fjVKvKxC8BuK+5cv0sKEg8tUq3RTtW2bv+
Kl9m6Z8ssxD1OKvJJ0FBUcyK7qI8Hs02iv+R5NshtjBJTX3clEJhzKe85H+S03XU
oHLS86zHR3CPk4gKQGy9dUN4pEx+kUWsRkq6LZoajwWDKhHNcvFaX3bX4fqw9Eg+
SO/B1Xt51gyTolkdst4Yw6zZsh6j8kQzlNtapMqCxfYDwJef6+h11MmMl+uLGglW
TWl1Zp4/9RxznRmg9N0jJB0crjzGB/jyLGURXhbuZQ3/tcTFPn9oqTr4GrmkRPNN
ZdVb2/WP2CL1DDUH+BsV4TZIP1ETk3C8YQvjgQqgr5oVFJzoiYDD3khL7BOy4A0k
72gAiqqO6zwYzDqb3h0UOnxfftZ4VWmIVVRHhT29g1Qwpb3HMHwTJtI0xlYxVtxo
FuzZhIyKHbqJTUAVXUxfPmfi2R5lZF70KjP7t7s46oq53KFR6GveSVUs5/YGhZF+
qDdebHCxpg+QteK4fPas/aVulHxvTF6CjIQvZaMj2bF1w/CVCtbiIKjIQGn6QaGs
HrgHmCUKE47GWwVSERFCW+vdK6+COZXjQSvie4W3i1bICQRsWUDVRRHJFmAV0Ccv
r17TDfKYcUYqSfSB2tM0bZT3kaPgK+xBU2m9dile9B5Xx3GzLqvYZbCelxiNF6Z6
TGwwPA/oPlxu1MVcnTIIRGp2fNu4vIrGSEFQat/kpoo7+EILlwyAQnM2nmTq3eqd
PBD4/xPfziBV8HsYg1KVaE/dd3eW5ygooSwn8JolterOtc2kDMi37BaEqxBSJxcE
XoOedx6P2FgdAWHYSr/Zs2FDAYoHywGTLdlD6LlBMXdGoigNXjegO66SLh6yQAZe
+benqWfeDz76tftlXPHmHZDGJ4DIAgXkbQsG0XbSoqWYrx21+elKO2Lj+a+StPnr
GcWNnX+s6f6qhZLFQjbrXFOkdB5iZcmVkeflqG+1yShy23WPKGULy+xD0b4PBswe
U5vkTibW26JyBsyDPCCMkDO1wan3IzY0VnTUP28EdtP2nm2pbDj5pq/otVfFHI8e
VabOSMWls3l3ATefZ1G8Wxj/Lo3gDBDhJiNSZc82WiBpDN8hUL4+p0Wj1j4VBc6+
8hN49KPN/2UQ8/VxhRIzn0gCDo4OQeShTPbUnziwU4wDwqmD/f1gwcEbRXe+FWQn
/WLAiN9977zrxfB2XxqrsldCy67a2B8Ij0MOs+kOqvUyfCHbTHjM2fJAmYeYKvY1
bUUxNpyQ/bFiP1P6OWT9ZF7WOn9Zx8buYCvoJY8Ntc0rVvl8oR7YTQjYyZFHIxO4
YtmFroNj6G9hdUq63iDHu9lIZsefJdMaU1mAPJ4beNvXaADm1eF6Hm14+IsH9cMb
s8Lvgee+e5LCjs0H/HaVRb27MCJ6pX8RNz66OEd1RHT3GuhiDeNmxK8XCv6J0dtm
nVI6AJqDh+mtJFYw1V4mcB0oNfEKxF5LnP9mA1g4Ff/9RFI9CFHVci75vocv0K7C
nJEcESGodZ7PUMBy31Q6PVNP7dZQB2Uc7gUNzTJSR2cWLtOOr4pSeM12j9rsNwif
+hdAm/uk0mxUkE6BfYKxemYJgBYhT1fyv0zLp3KywyeegCX1+86nh7UVGRLoQd4m
MjyLYxOG+5nK3sCDNhf4fw9fD+zp3Wnz3F3WH7Q548tBpVS3BUeegjGeVSopu5hC
lxo/ZiPJuAuJS/YfAmDLci8jc84IXzsYWG7kWaQezydrVUJCGb5fJMpWrt1vCXhD
r4egpV7Q6LamXmQAqL3A+FruLcmfMd++50Va8HNzYnpMtHDfGzfaShOBButh7hqq
0waZptcdh4BRUN15UhAlPs4Z2SIVKnE1ZINFvfx44eIt89ej2DQ8ckMbSbA6IM2F
Hbaes8RgvThIs9U+WfqGIczxMEumyScl6HC9RnJ/IjeAvPDViTPxdnEjJvD2A2xw
sdkV5rQvdI8wICaDozSgEr/iuq5g5TrXIn/98Wbaq+CnuMUnaeyu2nckvknb/zCD
N5gGHTBB1Z40uCad2RR1w7WRJFzbZleUommOeOBYuct7aX+JVnAlJpF8bYuhLFN6
uGRvoc8c85z4J/gYoB6npRCyBzOw5w+p+HCNw4MRrvkVw/vJdD1KoDqlHohO+jhC
X3Sfiwsv5fTYKqyCleyVF8m31QHZyoN40SjzT3+s+pGtpwacGyKYAIplOTDUW6pZ
23iRcDG5rg7V6sjHDOYLCcdhJtyuCZX6sWXKBRJw1/IbfZBu4QHw/DeRAIJZ1PjO
1nuUSqUfuTJirt/XkQfwlZT4LtEHz9QawjLjj9XVjKUu1DkrQHrCKd6V4KxXelyy
uagu+lgFr/UuLlcqO2M6kWvAc/mmJW6c6MNdDbT+HrExQqil23i69CSTjOrrBHJM
PLXRO+4HGvpZjsdusCa5Grkv8VqKSuPygtYrZCymTvQEY3M0JnOtB0/0kl8fqRMm
OI1hqXLCEYa3ap6/2/NPyxeGle0iyF0UNq6CadVycBSPu2IC2sg+2Z7CJrFUyRai
Cno6b2u55rCeUa8W9r/gVibWK1/f33YK9s3rWhsTcL9c5blfiY/9S6ustT8AmsPw
0zCA+vPzFmup3iprjn+2jNkcTTlDCMaz44x9HoPm33gQoMThP1SxIm6ZVOsqfJel
UYCtq2vjvksEutjDX2B6XhbSIEm9s09BlefVHkE2xm5jRKOuSO8txLHQpu56RZle
zCn6P5OBDMzebYDYtbRMvk9lJxYd5azHKa4HFoedax1b1FE2FonkpPJJSTQS7DUZ
jZutZ4krNBdeEAAgZ+yO7JsmWGWwCy8ZTKUmxS0AXWyPk4xaAj/68dBlSFEcBiIW
QV/sUme0iAyBdHfcCQzPTJFjjvv7sdJe04faq6S71CE7ScACYh/vKIukt0wrczuG
6nmhH50ZvS6tgbwvEKb1Xr4IXXPakUC6zCbZT+r/cHBra+qBUlgEG9XvOSao1amB
QdJcsN/1JZRejv1vw/e8ngPyrczNcn8gVwWRJKpImE94NZvS7ByWeWtPiuaClfZF
1ZNdVh/Qh8kGN73cJ9MAn5cdQKIFf/sC58lPVYLjNjo/f7M4mkl3IcE89smZ1puV
MyhSnV6LOpy/YbkF6Smq/h+3XO9AG9W59P3QD4XAm/QjRSBH51RIn2ei2T1+dD5I
idxFkU3MDPUQTyxShpjgCosuPJ9m/6jMIpB8TSlT7umKm08viyfM8PFS9rB69XnC
tFhScKGk+ub92AIeSCnEPZGB+VJ0NCrrbdizuFc+rOUEbMxE9C5PoTXt6cMbXIRz
a8TLhTpZhMDCOuc5yChdr0kNIpivIUa6E/e6zP+WDUJSC9Df9Phtm7XmfOHdZeh4
clDWynVYEUK50vLXNiCaiJlWFbIVaxSYbkkQCVE0hYxbefYAL1EzUJp6L1XZ8NQj
qKiNBlQpewAcp/GcxZz0+Z5fFbSTEKU9zqv70ZivWJMTUW94c4yqK7D67+njjcbr
yTmYZE2pto4jg+OnIholCy/uHCpDIei+QUzit7JeukjWa25w8hXAnIv/7AWqGvgK
Lba5Szie0odE6wrn2S99hYOQ8tPvfCh51M+oNTnfDc6FuXZgVrTXpYxYHPpTMRtF
tSQlULG23wSScGuL6TxDgewHsAmfzPI9s9+OgvsfRyLNVvK0RpskLwDdYL7c5eNZ
6F87MssdSTETU1P34Soe/A7Begt0dYWmKkPPN6w149rSezTsoCOD2lQwR71V5VqU
zKE9R8Mw0eP6T2zKyD/sBr9Kuo4pT/kZDHq4lcETee5l6Thvi35OBvBlw86pPQYw
MsTMXZovYQSr5+V7uSK0EF6z7SfORDbCxhpyp5dnAmQGzngC1uPmbs/U51qG87PT
b030CP4PY/HZnA5bmh+2JvCxoCucsBxodb2Yw8xSevqGym1IP8Adsccv+v9wNG0x
+iAyKmMfdPEUXoH6xCPvmbYZXgFP7BzdmZyhf2VfyFESOsqPKiLdzYok4UXtC+vJ
iR+pbrZlAVD8dm+jI0tJMwxkk9rQnXrnK5KP+/qIK3wUR3NlwOLVWO0pBeVy3uix
LJ7jXc6BvqnD9VyG00jiKyUv0xycpD7G3tLzqANhizN9oWtYhnpCKYwjojbtbEHU
wZkLvIadgZKxFhAQyzTOeSewWSzkiNn1aq7PX+F2VR2jC37eONxCrGUJvDljgEWp
/Ik+BdxzXOvlHj34pPFGAhjsMhs4c9o/LmdgRlcWsCHRW7jiEZO+lgJCCJUxCTQg
ZaPw5DJQJP3ZAKud0PPtOHwCRDGD9Lp4DB4CaX7Pb8WDjIr1ngm8LlYqxe1OdZvQ
hKviaGZOg1uS75eVNOnhy+Z/TG8mqZidHw98jS6qb1Wo4WRIw//3akR1vptZ2x6M
wdiX6tlp3pPX9nLvIChmIWKun51651MB27y29xrJCfwcRVEr+enoyC1NCxwowY/M
fwl+UJ6aKYfM2KRxroT/cg7sA60vcK5G8lDDf1f37RJMX0pIape5a59Kk7XoLUWU
CfuX3hiw/oVXYrQdqLbywoB0Xf/geq0QWInArxR9WMpM0BympyzPZFk/ReUYfYvY
Hk+uR9f4Buh9Crp8CkY5dItTc0NJODp+2YhfOAxU+mjNbmQ8tWmK/DAxNE6d5wmN
4QoBkv1oGucFSC+fZ1FNaoMH+d5FulT8GHvrZyLh/47MOkAXTXAFXPyDy5VYwV9M
k5wN/sDcjQl1/Kar35XEvFYtiAw+QcjDfWE9oCImnAREREsO3nGK952ik9jI7xWp
Kou2wYjI6htWeqfGpAA/6wDcMe3h/bFP/y9f9Ir8ise1W6iRLtu5nCH1HFLWCNtl
blXCyBFWxosiNPlls/ZrpeKffwZK0l/Z65HIRwyz7LFPQdNaWJmdji7Cet331AHk
j0X5ZPqQMsx9rywe67FtgRh+snCTfzjkuRidQYMIGsB1/UldR+MQHZ0wXV0v0svy
5yjtwPmhkSizqpFWUHsW8gkDEWYVmeMCQyqSCu+LrXj+6c1vi/QV71oIRxxroKPw
qNBu8T+4TyOYPmyXnyPaVNA7/I5axnaBxecoezoE0tb4rKB78Yk16dfWz1VHyiZy
N4anmh9YLtxXSRYF6lQo/5nhdfYQ2TvPUbP3ea9S5/ioqIC+MWF0l4sW0E9xOQby
F5G5QUbO/lRMa0FxP4ybc2Ycqn+ZcOG4B6CB2VcLWXRQc3P+7EQcu/ARWvZm8Dlx
BJ6acJhtgiNz7bVZAjxqXNGYgf3AyC+G2xPHnISZpu2jAEvsGvJQdIhISFV8Nqc7
veXfiPRQOFH+DgPZwbAyr96/QgEb3OgTkl1+wbye/7vCXD7+crg5nc3RWQi2+RHU
QRgcl+M0xWLtcoBWk24hCx8ZJGjgG5TA/iVORKrMVFeP8aoiglLSHFzIBNFp+Wr0
jTXF+fBQdqd0mLJw97jNasq8z3u7s+KWvxM+7G2kPAcB5cgKYc+ZRdOP20YpCx3n
XOZ9SpLrFqqpgw5MiMyHS3bVofaojbrIPZ2BPAhAuZ3hSS6Q4eJ/nlt5IR3gBVSu
cUEcSxZSDPMUoni1wfovaaEBtRpCvp5C2jX0YCdMFqhGAfK6E+lMObjlnNljqhGz
4xqDXlvOKl8+XKSbB5AOtV+s96LZsGVnDTNsxaEn7dSShGMQfDgGjjvONqqi+Ktk
4Z31d0JByrxQTxkJvX8XwjMTyFBEfuRACwW+a5Ky8NwZ9M8g1jpiO4I5dlm8h9rt
W7/W1ddy5r2jo6YPV3DOUA01tPTEscEYufCC+3WFy8JXby+6uQN57JbftRKmU73M
JX4eSzQJVuxAoAI1Ocw1+6tx9i2QabKyVaNAINLBMK1Z9BQvgEabhbBWmil4ezAu
3Ax0MNwrAjJlRdrrgNShuI/TL194tSRS7wgNiNXrWokw0/0cL7KIBPRBdMiH4ImR
dJwbJ4OIEJCryjEYOoUQv1ZqLFbU+NwTIu/UBEVMFMjMn/vYYmkSl24Jpy+HL1cT
z8/OehxY2K2ObrbUELj7o2eGEUXmF+pZmJK+tCJQ78KBctvdQpAB6wbjA7ciwc9f
OWhtW7Sut4ftL3ZxbskjBDYQyojJXpDm0fnpBbgzhqNPaILKP3m38DUSQiEzXK+B
8KjYEhudBRsd+0LKaGcTOpxcGhy5YiCICGawDR7RBxHmo60hXDNsMe4U452bnnm3
iwcPJ2D3YWyX3r782Tx0kCQQv8erk3Kh6XbSudMoniQy4UWEMlruG3mosjw5Bhv+
95+1t8VwvKNz3n67kVOy5oHpb70U1OkO8qXHbUWq3EOuHkBOpQpkOQ5KY0wglGuO
Ql2gNyKR4ImvuAMoiGrt+ppc+myiHt6U4WUBG5axYjDYSbjmuCG/qA0uQvFwY05e
iHPcKewrA3Bh2c808066DcVdnnLPB9o+VwFxI3hBLcls1vJoHdV1A81sH6geMyv8
/GimhXEChvoElTXDYFdM4fE36rZaxloAiekCg2KoKhF07U4n4MCI+hCiAWtGbbbH
fGKqOTLgBHlAtQzFEABF5Y7jARkjwOBpcDd7j8civ7Fpbe6mk5WnbmTKI/OnuSdF
PLMIq+WVUiNeWNrkxJe00OaskW49I35vhGrwMzJv2JkrlDlPGxMtQUYRIEZy4Il8
0wPm3y19b17wehykAVYcqP5vcv/uUdfI4EfD7q6aF3lkHSGI5n+3jIX3SQttZk52
2y4HpeRxs5GOqpbzk+9GGkY2loxcuuNbbhxv3ioW0BwJbYc4mvA8Y0olhgdJ9yBr
VyEvjqOSsLgm1WHCFLlZZE4//b1NpGJSctH1M8dBvTJyqloFOAY6XZ9IvQSo3S/s
/3Q31TrZwhcMJk6yIiJ3TVx7Jmm6LLARdaov8+CRQeJE2T4QEtbLB3YEDVZjvp1n
1xLmIQUiZWACNR0eDswM22c92FbHwFVZd0IZ3FnzsxVT66fwBFjSZ6uvk03mXhJc
37I0GItRglW58wfo7GPhnFJH6+fbzTeinjIff97LUNLCo6K/TfE70d57HNnuqLRi
pkBGUy5XJJIo4C6VsxQm0HZ01MUjnMA9+7sFIEI1c4uOEVkE6R1BXHizBO2IdOyr
RRLx4U+NT3tQH3/kh86xmqxV8IocqAeZEjMv+vklGbunE0lPLuXYNf1TTSq7aMGX
1QJN4bOZ3pXczGzQaaOLeE5Lj4y88WRRORnQSReW6Fbg/jtAxhqINC212H/ROtLc
D8mK+S2tiWtfzHlEd0g2TqrGNtGy+bXF0VvjLMBIpykozPoTsoQp2c/TNEyANsBH
agTKN/9fq3NjBHAiazcChScIsor8MuyxUge6yg04WLK9rleOWyF8dd2J/5vnorAK
mbu/Gzc94DDMF8K8JYSvYBJF8K1SbUvKgW9QeunKqDhCOg/YszP5/kDzyXBEmYtt
laqUPF4YQxtaHi78UECwjZclzUY4kH3aLQVztscabsly+7pqjp8y6uG9vX1aRC3L
ee7et99SHBJO7i5VM2UM0T2oVSTP2eGS5xvSllSeIuXUIiC0mN1XD+Ni3yZUoaJ6
RDcrS93bQ0pVGOmcwh/3RPIyvClvDqCXNQfSFVcszqwntSi49O86ByULUD5w4zcK
EPi059YievkAPnUxomU9M+DQ52wfIP/ZTz3qw+VIjdCiuXbrCMirxaSKKjP5SFWk
MOrVhU515SdBSqA8P9jpwmsshBvkiTTzIXvE0a0AEpkFAWQkHoz3L3TyDZ73bdEi
c8dh0X+Nkp3XFiV+0KycdO+zMFMPKsR9VSxKjMqGP3Ii8nvyffz9ACo5rZzU6eS6
5/xH7Hix/74KJ48W8NlPMyIpQ6/63k1/F6I2ISsCqdPPo5TjxJ8rpK7Q+gOtQRgF
fAxBQf6c7AM+JKSBlDIJGh1ADFWa+U4TgHpwBd48QhXfjzQV1R1mrJTsi1iPf91/
f4wOs7LfPPJ9dy9z5RGBxt/pwEMGmenuIJaah+7em/GOcs8oyciKtL1UR2drWuFK
dRRLiRaUonDY6MQZUU/5OgsYCWJG4uSToKern/V0Nm3AXShcbiPcSR4aAqX3RO+a
CNs6o0ALPIatWdEnb3UTqTzpndDt2MjHk65fygjOkyygj+y5vyj2Jagh3UroA3Bw
4s0I0r67W4z00KKQ7bQZK+I3GnD+9jXLVJ+fmBbxUe74g69eeUEw4G0Xgw9tOfGr
jhuQoCDbiM3TESABdLClAnnlxSZ2H7ryEG5Xj0O6A+I7xRwJZRYcCLmY9GCfDzyc
KiGNMkLP7+9Bu/Tj9WZBx0eqKVDdtQxPVT+OO8dghMo/nRLYukQcXb1+31GTaFuK
GtxJFyNNv1GewSm9KBb9eOTpewXhtTraWkaZ6fX4VgMNThmmIFDAHXxlgboasWoO
nNOGcmXyFk808Fn87wCWaWYdcZOKGT9L8xfdBBGnLPg+O3qKVdjDjrrVblBcqhts
ox5Aeap8gUGhkOzrEY1TuBxXI1Z+AqkL/hbPl4SSs/QvOSP7xj8ZAzbu9SD3Ws5I
TPY0nx5U8pS94NT5QAnEQ9vXXNtwAME7cD9teqzvFfQRC1MWQHnkbmJBARt7hsOo
2d6sV/7Ao4T/MtNrm9Cl2HpvZ0zhIqP+bVIhKq/022ukd1bZIyHzfniFs8Tk7ELm
jqLusUekrB9N/6t5JsScXcjH4ODO9LLAL6JI+opaYS36kfuHXc0nmzU8e0zDrFF8
n+8zBH7OGtIqjlrk23LgL9vKepblPi4PClPk78vF6Wexjv/BmtUZMi2P5kwpBpOG
PSuC+oEabocLMsaEk8TP/JB4YcwiC9n//Yuq6Fwj9q7RCzhXFG3jU2AzSfUZId84
4N9O4KZaHg8hORJaTZ9tPibK/k0WgEfN5o+io+A9oiP6T6OduRzzbRrc2hGrYRAy
iX74JeG1/RsICWEu6+IJU0fmgv/DU68taIvOYOj2zSXlUHSUVDnSpjeOyyKTcEuW
Uublu0VzHzjyu1jlcjFlSj750bRCiLydQzSMif92OyKmAmlS7UsZxXP4JqTQRUxw
6Yqk+koNWYtuGEqlEeK8dzDT+dYDSEdQDq8+il7IpCnNf+Z9tyOVJnfgwNV6AH0J
q+OClkaTq9MHMEj1d9i/IrCH7NDn5k0jkUijnnK2IbrCwWofaHEyRTk5DRfvk5Yx
+yv958xX72JHpNjsLsf7wKHiYg6oSK5PBFj9fqIj/poQulwU6eP9+WzO4yYnj/gI
gqUa4rL5Gk3btplcS5QIeUGcvCXfKWnQ6aRolDxWw5utZ5GBM2xE3orsiNVQJ9ty
aD85oohZfCiBX/b46jmtEjXHsCKU1hyavWBvnaL/jfu9Q2/cn0BTqZvJDdmpCwdp
THemzt8hs1PU6KRCgFPTvVYYB9Vtu7axCFbzAVEu7f90xhamR5da8aNiDm/PIcoQ
ErvsWKOlPJWWq7DnyX992Du/AaAmrTMVMHn1NtkX0DSAlYU9vonynfHW0WgWBXvO
j47YiVQjvnG5Dr/0R1H0UNSqjso1CYsF/XXUmDqASH6PkOuc0kJ8eLr5Lo5qMLaG
ndNgmmVOfQD/emNrDKsbpiOkvQERc/QRjAOnGfkS2kb1xKtBa8Zzj9p5QoU4hMQS
1htV5RABRJqCv9GxQMwHSYemF07QHc/Bq3lWGO66IZvN4lJYsR+v3JlGR7dy51DU
1L6bR1qyvDpurEhljnq26XcVblMQH38aEfOdQdU7HriXtcnQszyBFqNuPMX6pzrX
h421Lezb7teXjKD7GGHobN2qQiwqpQXOvwD1fcbHQxIKGFaGq9q9EAZJhczdcCqx
8WUSvjTt7OjDsiAXQFXe86YY5Cvu66Xzxzw6NspLLGTakAk3/z0+AKDlVd3dGWWF
+EsEmbHfFxQyJtxByez98QnOafj21flXB7lbpl5W8bDKkOZq/abqktgHnmUoFTfD
fRS+z6iwOaqpqeEd5p3Nsn3R0+Oru0gRSb0uODhhe7CsOwLsyuzFwu4mGz0MPOFG
qvlXTMGs5CsT7u795mFAK84izGivgcfLWijmqQqoZtJo3BIe1yn7rmGvnAWvYv0T
E+69Q2oT7s3mWjlwVplchHnkOVQsg/Bl6Kx+BijJELzAeenS5yk/B29ZmTfhSgUF
OM/lmzB6sF/RChUm4YCc4mhVug0IvyulDDtaFwCPy3Utn9PKbAEXQw5yGv3hP+tY
WFlBXFXnW0b7K3/pnLzf1jz4A5u6y+jcCAm2tifZr6lxab3bqYg7QYvRhNl9v70r
pAXzzHSGacX0uX/QA9P5LFE0+gOfPzvyr/uSfLT9mBSGwFLns6tKQlxIlc8H5Nid
KHd0IDfPu2efaz0CN3oDwh0KOArWi+BT2OqMQXTp1AIDm9iuFj3nkuCgDiwYZI8C
6/bh9LU5NxE/u7KpHmgllIawtGyWa1GCk7HDp6feOQvmCUNx/9rXr2knzqYd9s5j
gIuR/lz/2Vtfjn1Q1yTbnk4JzNp7AlOyyoQcZjvJN6KXxoSJ3W6fNzupwVzyktMW
UkNB4rPYg2NpEk84QGvOiOU2KbQVsi4oDnlPCe7/UmF3QC8+ULewt8vmQTWVIDdA
ptdh7jC30fd2rhXKjd/iVg54rngZAEkUty/AteU2dl2WIIK2RKssKBgMouVeOdw9
zk6SsP28ibnEId88zc2FuHYivblSF95SyHQoJGH3qp9I9ZPQJw9J6KObhuj2+KQ0
aXpkRv0sfd+5Ab1qKB7Wn/NJaTpJhdoNRuTJLUyWuPI5k0lnlfQ7CDrMbqT4Hhbi
UnLCsZwsXuKD78Qly54hGfr/b9ofhd0GL8sJZylV2ncrqWrY8jDg024Zm5VP+wZ4
pCMtOgxGNh92TdNd6mLSjNsSsTStJ5KqiObDWu1WnW95T+bN1sTDK2x+gWgnsjYn
SUNeWLyQ/+8KsMG5NSjyf+CI4BpHkG+e0jM7xg5cF40hFYXhwofsXd2fYr8pwwPL
HXjwjzTvca++YtYcyUt+cEcA85EipUaLtY0hV2XO1QOmu/PD4bjz+sYq5yYlIVnW
6aWuej90HDEd/WTtlj1mA/ZZrRyHN1IrqBXJJqfb0XWVa9OBCPBqJqJN0MeTHukE
5gdfwCO0r94oWmjE+VYE+zwbjT3ojpjiUiDCkchjGfl7h/DfPgDSqiwYD6AKLiAJ
pPa3aXaLfxskB8rW+ztcocaGow31+6jyewLAQ/WtZnUsGMsGhTE2AuzKorncDQMR
tfcwOd4TTuNogki7aoM6NYPdukIeKVpAQdu8Nq0C5mmR2lfJEnjRoeWC+z0WTQVo
GFn3/F2yvtQ+UJgNnl3GWZ+nqS4Vt4/cGBxTLaDpHfRxrDYfQXZz/imIrlDaGEBR
nyZX2P8/V6xSmvvA70aM9lyj/aF+bPEhL363bzR3DMgXoOacU9pia1MZ8OLRSnYR
66YEdVHKA1Dv6UBi8SvUTuBulf/jCm5J+8ANw7LkoRkL0FymDVTZvYBrxJaY3Ido
S520T1pT9ttQnWuKFnxf7hI/bIOxsfuhVRGW+9o/PUrmkdf9iQSziMOQ8uqV5lvo
BeEMZTctDFWxs4kEJPTd6Brha3WPwVV3XLZCuocZJ50nL/D71nDoCftcD+dOACSA
4DXIzMUscc5V9MHRUal26n0q2quWv+T+/bGGHADXbGxKhNzKyi4wGSt5pvk1oeFN
vf/vaf3yGnJrTVJ004Z89V0xBOglkOIu3qxQhF8zu1VU2vhAYWkoHc3oeMYjg7X/
tUqXgET4r2HGSpdnTDj+kEl3cRCHh6uH+vXhglzkxd3Mw5IbUVW4iz0jUzkKh+7X
54TveFzZKqZcUlKoWH1VHkTDotLDkoMtHknlQl3ky0+2PDjD5NiN7pintj6jBkm3
Uej31A/SjXvG2uHo1BLFS+kktkiu6eoeJsOFmKKTdOGI4unHE56tnJOdAKp8+I7J
WzpEBWHEQw2b6bHFeEJ9hx34L1TSNb2RURsgNF1Y4mrJ19yyU1irXVJ6bIiT3J9m
jxLGOI7HmnpY7yt7yueVCr70XqOw9UrKTeZoqgng9cwF/jJ8GdNrAbl1pDafourN
p5DkLp6rBmsVgfYwtG7HgLSGUP1wrYNLRC8beBQLsljCVPp9pB8D0VFxQJyJ3TzK
Hx0WpPw+7Jy0cgNQ/nMg0z9Sheo1XBdcwwdW5QXZvBFxOqmz0Vn7CAJs5xpM7JHd
PNBAch+JiWTgsIAIF8fZpzSgC7cMkVfrGkoFjoJMrBFOESjHSQiy6Zci/Iaav6Lm
dxPpuDeWuUkIa6vQ+eh+Gle4wUAg96/OfRPpDMAxQa/qldGoclQ9e8bkjpzD3/fj
J33tku2qpmKlSH+GMk5axM8hbT96gjQW2pwMujnTpgsXriPRCRPT2yzX42TzLriz
urYNwrrGNXZmQD2Gum2vgbPLDc4T8e6c8YEeC4Ce7lfhS9vsycVpsdkWkd2NBHtJ
Ao8cEQuz5FygNY4/wCYX9d7+Uo4NqobnWb7jc4ypxHtn7xjo4N8SBVW1eRcmmCPH
fe9tjHHoPB1PRCjN0hJyT4nj5hBQDPlXZtNgr43W7OS3mBj7aO1r9hbxO0oT4nz+
2OS8dSPAV1YLfQ56Lef4dsG8ps7DXH3UTSg3KAOB8gtFq/4YQ0oqtvbGVKkaQtai
Gmibp4X4+NwwKd1nffcoIKe0F4pcFkrsZODmA/9eCCYcjcg0r5kYKM3o0gXZFi2Q
BnS7vffh5c16a2+rUnoq/wTRNgNwGMjXUUYTDaliNgLFBdlj+FZE0ay0kuc5l3+X
Vv7n9X4eDxHjAbt3q+UMcp+82lHCvJ0+P5Tg7caNTkqECvTBDqsA5PbhpJ6mOdR3
pNzUvPaKQurnlqoTl8gHbtygvRI9E4NyHvLOxAYOFU+nJeo86GIbsIBOn93md2RQ
/WQPMntvL2STYcc3G+QMfqtXjNVftc15AOzViwZ9fXC3/+FyX+nAUM2N8QIpJWSq
9aO2jcvwIvN8Sr5Bgi8HdlU+3av0mfPLOXigxNoDqI8DeUNa+jso330ZgzeRyPV5
2tz2jy55Aze46OadmoUD/omXyRfOih6Dgvs1QvbeHze0L0w2pXLPa22HhMww0X4h
tOMMzS6DpAxeLrhtAZ6WG6BLiPgPTeu8AOqj/1nY3etO1u7/a+7VbJzMAh2KokNQ
eOYn6INGWVW2fsgUL1lsclvl9JTq337dm3JUxLiY5YpjV0ClwklA2PgEYSnk5a1n
Vkb/u0z8LhMiqEexlfqFAYad4f0LjmqfoF9ztSFkrEhFi0fGbzMGlsql7YGX5Xbi
ltbnlsYHee/M5ePGNl3VP9s5T6KUkwPSFRFhDbPmaIuELIFCnLi067tTrPYwujbH
qhnBJ7J8EVujE1Ygk7vRuJb9kY9RNUblmvLqBqyyIPYAnS/FmKMNSiCjqBD44KIU
dgaQ2ti29iYPYsZV/qaEJexz1xwFFgFQE1AVSLjFKio78X2WgO4RRh4iKHAoG/o/
TcBtBFiRd5eJB/9LEYG8iam0JxxhsBkqhEBQPs1Dxxm2pWd+MMO1WdYnZoFYSXWg
kvgzdhgNb1uqcCSjV64sbe/xbJ7v6PMruvoL+75J5QR4EpAy8PT3co5gX6iVsXdq
qmTem0Rs4bqPCDH2EvhrfZBCaMjIHRC7cqYn9qQWIYO64KFU4c6nSsXx3CgEIPwn
3ExPuncoxywkGcy97QWbPtLMAP0u9z/9KMZhu8WYHOonKnVMst3XyFBuEn796FB+
b134gms3NCXtvdYcJ6InAoovZiDq1xTkhoZ+eKsTD7Pc5ZqY/+82h6tjHUxfpgs/
zojefiIBpcPmmGvcXAA010ft+DmqndvW2V0gabqvG2fW8w8/nAktgGvmFS0+hAHN
9+uAUcUrd9ctYnaTVCgVzb6BuoD+qt7mX8pIdBAW79Iry1nQ3IILdf6lKYHHm9TM
jpuVzlx5tZL7tyEkMXI5QzuvJqd9YfNMCAAGQikoEqmteDunR2KiDzibqvyMCQZT
2nibnYSqqPqQNQ6Hsl0Tlu6R1A9LYzack/R5sMTFZ/omrSBUNSzgbKac2D2d9oK1
8ZUiwae7JGxZYdHV8r+3bIspMuiK/TmnIcFtFeAQzeKVrBHL18LHdnxnUaml0Uro
EHLd6UR5aDcWVEzkZLQU7Ci4aswwOmcQHYgDT02OEfF6lYW21vdAwyeZq0W4kOqu
k4+BStcL0+SucAJ0In2jt06pYk/8bJyEnLIkgDBzeP16Ctqmkanpb5XW1c5TxOYc
3WQonbxv+rLqmImQ35w7muk53UTV1Oq8I/MWCyW6aA0zN80n+GO67vE56xqIeHP2
OOuzkIbruIsHqIGIfzposZF6aLyXeAKC6sdU4uu20fhey2GS3PtMXClBwoWL0XUZ
rMd/8Y3urIAgFHGc9c+A7D7RntxYJlMCGZXIEHsE/dYEL2CcF2mFR19baAK215LN
zFsHY+93dMyNwG0MhpcxoYMPSamfuw4ai6IhwRp+YtykruejW1wPkje+fOZ9IUoP
XEwanM85k7UNzQhYM3tE8M1Mj7Nt6nIYCjWumO16ofh931RLotzU7I9z6jwJSwKD
CP+26m2tRktfGy+v4v1jmKWvZzYEZkevipJGhsA/F0OPUVU+h+fGUwOOisx4M7jL
zaezJJD4AhWvhA8AKmRV++L2AdhZRyrOHAbPRG/Q/XybJ80o9+ESluvZgeX8NEgR
HD07Bf5OEhERTVLPAItlmz+WSXhizV08M6xbY5uxuTBPDaZniTEm0Kw0P3bzNOOS
9kwnFaoFzivl2oh918VHlmQ15yZ9JdeoQUKPJ8D6RpBixVE9vBUE4782GEXgYhmG
c+F3iO/ch26PuQfaxpfyaOFmM5eLTqRF8lN0E+Nyiy6SqUhJO21bXrzcBp/JoFaY
zcY/BvDmrGdJidWHODrsSqj8eJ6eLqLyXyPsuqT2BsDsHxZcGlI+Bh7izI7FV0UU
ZE1wIldxJ3dc6O1D9CoAed2RnpsBRKUQCfDMP0EpFyBn2xEbbQUh8oQ6wF0kOKe2
a8Z4+2HtjmBtJpSv3arpTWPlgmeTNEMf8lEqV8Nl4/wH7GkOu7UJ+tUKzAfZA101
ZA8hlVX0DqVfMGol8Mgs87xmOqFHDER2OjvOclPb+PWPiXbPS2836drnyb7D2tzg
jG505ZSZppYp5WKVlxL4wLMUxic+WlZw+ucxGU1ktXgCzYj3d+/nNtQ9LrchZ4oO
gaEaj0MuviSB66z6Tl3VOrsCAyWcHOrKP1+jdaVB53RoAR1cKHWUm5y+qTXH07tI
Q9392Drm3kKCZPwDKFPiDWiqzyo4zUO0DkfSQ1md8wveZnIPc5iEyAF37sbInoVP
3MCVKSI+Y++OAtzgn13cqJ/EQjWKmUJljjW4Kon3p/POonKKIpgxeKpHzzfnpeX3
L3yT8LDrDjZzRECQ4xPw1R3NB/QlSWsY90rGJhQLxcUy6XcZH3ENwyK+e6KCxcPy
kDJqOpWA0EWiEUJkPmRU8xW5KmvXhfJsgKfHqv0Mon1xCwj4BWngPGy8PbLvuKIq
yDetX5pgE+PsoeJYjxc97Fbu4tyEoNCzAKu2pOm8jWlihzaobtmN3L0cPbnQ24Kr
/tLstRfcIgR0z/P+MfRqZU1xa5V8LMapvKqd3akJBAftqdNavUK/2cW2CJNGbHNM
Zl0RE03g/tpiNeeAEICMiejGMs1iNdt1nSMMv/iNt0T47uFt3Be2VP2DNsWoeKxu
bLy2R45VLDkFE8oKfvUcfTcpRxZwPUFhgPvH/IKXyy+6j4wWobhom4XErvzN2Zm7
jh72zwVDfRu0MzZI5lbLq+Rh3D/PG1G5P97mc37s8b3o6rjLOFT32sI9L2coqvjx
igrrjNqVycx+IZIMhv/Ks9lMRgJJGvdHqHL+sfWc2IJLVZFjoPiUTqiTNYijKhG7
F8ZA43Z5nlVJLMkS9fd7U6f9d0sS1LT4/TN+/FepSD3G9AxY6YHXVevHYhJRlMvz
AIKn1gbwDkjbXpW2XkovaHcl/EDxnhldr7XHuY6yaFr2uRiBZ6uGTAoP81WQ/RsY
kws2vIkIAgj4zlJc1paizVJ9EXB1CprbN8p6SX+6HGKtxGhJ69PbZDAIpHv/7USW
FFlK0Yy4mvumyaRqZxt5ob/VfbMDJPdZ+F8OSoN6v5CD3n1SsvNcY5raE99eVBZB
FwGVsM9ZwmZGaTSgLnosBqbqVVZBrqyx4GfENQgRH5rOk2zYG9vFQuGiNC6zXJYU
XlqcIrIcS5+HBaI1yv1OscvzF3BoQwWgvAFq2NVdXkTwlKuBu7SO273Q+RU1MqKE
DzcaOzqcOwbTpgcduN0Q2nOLVWrSXTf16Ea6vNE+Jomf57gA25tvV9+coaT/pMoz
jDyS2yBf4qx9iUvdngq0QmD//FzhxiPPersvEzZ6I0Jc+17qX2hAEzd2au1x/YH1
Xi73tO3Jqd8l5tXJc+5bkms970XQRaDbTHTMRgjgCfoHNu4D3uJIJh+/ijlUwsb2
QBUEQK6rEs5SGxM/6i6daMP+0srWoYfHn7TJgv29nEKtKGwY9mGz7pbT7qWXCqIA
xGvKPVctzwZqPH7cjP46IYqyaPjuN4orR4qkSabwf9ECVG/sAsljWoKO7s2REM4K
OEHjuRKsZ/mO5YXs7bUufzcZdCzs/tOBeyEQa4yKC0mh5EP20+Y3pXqN7oX/TcQ0
yhE4pb7wwoodHokOeHwPYFx2lBMnZVgfhzwCj1gMSEJ6pg8W3scz3c4ncwKR4Huc
nyA+4MPLa7lUkF3ETveaKcfigZ3CKbDE+VuLMWITjeybVF4QYPz0jL0dTW3Me8uI
QDbXyIV1LLNbv3bKamOYZRX8w9sH1tcOEOZijeHU+yZ+VQCe4qJZ9ZFJJqMjSREB
cuPFccmdal9EwxXekQ5QAP7Jk5UU3P4YKQa93ThEOtl2MDr+9jGhBvUUV2i4mhuk
ydX0k65UALTjDAV8tOmw3cxtUqW1O4QceSYkNnPXGwlheT5Ry8lG797Dol39BT5v
jxNsfQ22qgpRtkAldKaZBS32bqc3aeM7kVSrMyMzrXT5EBxg6Ukt7f3bLHZUTL7l
JQLYImS7rdnA6zMa9RxhF6/DehMxx6m2LpWMRvtu6SqZ67nEek99fJu6am6waIbL
qIvWtJR8xTvDP6PfXc9oNkmlXXThbTARkkk2EjYr/lRh0mK8/hLrN5xivayFPP8z
QXbOm0r+RWaC7kAoxcdNsxprzXplBQi50heAbxY3j1bzb3vCD3wXzo1icCEymg4C
tUAMV3cCtSg+7AUlljiZnUCSFuQ1WO4xXuX3gJ7qUADahmd+azu/4XP6l8lgqR93
GXGGNj1vDUOVcsuE7QmdsDOkvFK+b7qFVQTUgeEFgHyZ9CAzEqBNckPT5I63jedN
QaNpMHAw1pgI17TpJ5y1VN4h9ACXiuwsEPwY0qHn2Ba+Hz8YEzUyKfiaYOfoW6Rx
/yet2LGXLmDAjkOjaZ9fmkIX9Rj1TM8WF10CJy3gdQXhOiT6/KhMXOtgG6MbhuOL
JtNsdD/RExDNSpzfkrsc4S/GxfwhebfBFH+ugbBj+jyEYbA4uzc7fW6/KN+7DEOz
Q2T6Mye8CcwQJFGim5wFdd6P32bLMPTaYz/H68ePpDKN5cEQ8fgj25hodU63NYds
HxI0PwZkSxM8EcjCF0yDi2zH3ij4uqYsIpx7UytiG3v0uSWINndr0YZyylaQ2NQB
1VPAFv2lkJqaqpMPJia6U9wVfgjKureJOwxU5I7WBTOpERgXOPU+0rSjTsl4eBRt
ZvyZ2V7Qmwm85xDkVkBoiDjr4Ym8MVkrxXtFrKXC9IuiqtT9L+MXaOlIMeWb1Z8T
9w77QVxNE2wdxgaPqO/ZPTjcUhA9VlTqz1mcde1Al8gFyP2a1K4us9Qz4HpAvsUB
yz+Vvkz9IPsLB1hq7NgHm3pEIGsGora4J6eUinOQDivkCUUh2dG2a9fP8l8dwyIu
CgFAYLg5LK9btrPKfFy6QF4WyN8w4vPU5GK7EU1AVxo9dIhWImxRO/n8wJNsRU6q
dSx3MwlRs+nfxsQmFnd/bZmha46xnh3M36Ag5EWttXUJwc56+iQOqaPKcD7K1Yn0
iMnSOJE0LSrk9ck8yB6E03pp2l/URth/Swf5gy41+7kJ3L9uEMfWgGOgtDo9C+X5
QPuIlxrC15inM3YJ9DtJEHnYraogi2zEiVVxAFycm0CsDbATuZLa4o2m4Uy5ntcF
TxY0ACn32SjJtQDWb48o7MzdWGmfCoucB2aYpa634hcC2WZDh3CQAGs8pVYU1F1+
4miU9b7e8P+W1V/v5PD3DDMTaldGUQyaGL3QevvX37fgPACNyECktpASFqCoY7UB
+uw88Fx1AAiv4Utr8NyzLk+GJe8BXJ2hU55xwC067Zv/j8HshXMCqsYIh8uHiWEM
wvbZIDlRHvfSrjiCnTFuR55xEe6QvGgb8M5WCaq2zBz3FSml40x8KHP4nhriWnRa
NIhPiYJtSXnX3bv7EtTfCydRYc8LBfEs3qXp3ZqgLXBEh5aIm4dzJSU6JB4t8saU
YEhCjxerAxlL5PMJ+SJWAtqh+opIK/Vp1KrbG/ys12Ryh4BWZ5r5e433v5afXACg
7wd01h/CO69qVPiOg2AZq7ZHVzFbDm/jGWqAcPdaMRV9nASLbicOt8Ujc7j0Pfvv
WHL0W/tboB4k/E6n16bcwuc8QF6iEhbhPqsYq2rGn2gz1bBE/kdCPv1J1bxSIQED
VISq8uDd241HeU5FtpNxYKOS/E8zygbuEa9wm7T1KEJWoisL2Y8/hPC/H9QB7HWC
CLcy9afE6L7N+cibxK4oXNlrSGnaYZSjr1OhQgL1Mpn5D/NMF77bN7/25WgWQQ8k
hSXY/3dD2kTN5MfcxM2p2Qmkq+wnZxr+jk+bDpsQQB28c1YFeQo2YoDbOey8Ilbl
WXuH/lK+DcD6Tuo1ox6QQbH5A1i1hTAIlZVFBP7KH+HNUODh/2Vy+SOOmltMN7yS
8rD7J4WJ3hI8SU2TvPK9PFVFY4MIE2h2rgYDQTNO2fYkJoq5GTrhCYC3oyWIpKZi
iQlFn03VGRBZkJUDByZLdMYMkDd0nltSBTcL5wQMFA/8VOtLBRjGQ6+qmZuJ4GpS
My32eKL+eAjX0nVGuCFbUdxJG6DheyYAdbxY2ebL9Oq27uLDd7dXmoxlrQhBwcni
5yP/QRqiLo6GFwXaQzZIGyKMxGmJ33mpQJ9n7YNWWiyH5O+Gcb9RBzGH2vEXEPwG
lV+2f0pCk836xf81FzmPMPkXSeDrswcsOwPHmjkc2Yc3oARNxIBD6s33FqNTjlU8
UVLjFlueO8Q9t8BciEzRSlzyiKdDhekv2iv8KzUfFy/B3nWvLRagq1NcOqe31GHK
ykfatct7kCBTmdcMuQ2dfXZxSZctO/8MXDT4DSa2tmRd+0KdjjxdCvuNSqPCnJKf
2r0WFE93x6FxmTAdeCE3xNxOiUckyC7HukDMrVBKpKrqcSwrIE+7c2GF8L019Esq
lRpeQMd2H++xyc3oMD2jCYm+tcVxSbXLM6Rzc1gUVKKR/EZiaYLOhXbdwohjyW3m
Kr87Mc5LfnQ09y0WiiXAgpK6mI65jd6DLFB7VgnFe5CnqwjXVBpLEcwy9vRLbTea
9wX64+7cCdXCZl90BHmqXp33qSOz9GIMmUhcnTPFEwlFeFbI2gtsMWGM3qOJFGTM
e2Qs4lQ5UJ6e1YuUqDIOWzKIBbvdl0DnrGNJY3/uynzibF8kjL4WwLanzDRqTcWF
3sNg+05Qo79ukuCBQ+09Fqq+Vx1RkLjbmt+Gf3xlVm8sZTvJW8b6Mhj04AjSerCx
BT6gIHZklSdQtKkD3k7dM6zeQCq7GAsQhDICxQhwWIIKXpRhfN5iqoYKboeWIfzT
hefFFl8J0LNszZqW9hjarPmeo/uXuqhot7JEu+aObZ2Teg6EEziCg4BibYl1GtHV
RYKG2Zq1TXsKL+RZMs5a3eCGt01RMO4FSEIlGhT1zV3HlRXYGcpD5h4J6g4lkbGy
2LA1Kso+50BCq3D0ny9vnQI+uEYTujtjd31EkQJQ+LrwN5qcLK0EyH56U2PZG09+
8xhaF5wSix8EciwVkGAcLZBAXeM1HcyfenUSh8TebWx9KdB86bl1vSPGkI5dPdDR
ZrpkwHEC4zBAKLXlgX7CokelmVbNGNCe4ZFNfgtJoe9+EEUntidIEIsXBotfMtKj
mNc9lxip6Rg9wS0YGl8lWLQiTcetZRPjd6Q3ZxE66DWvwNlJANFqWeqyGEU00LJA
PKy100kwhDP7Vrls4PbV5NEdBm7HBp3tCVt15wHSWch5Cf1CQH6qJBVtZevuSWu/
GqAKO0jkzNnMbVuSRCCgxKzXbBSJgcoaxgR+8NJMRlU6uGkJNhy7ckpH0qF2aCrs
/BTJ3GcxOvfNV790YsCccWDSLHoSvkGDHH5PhF+lr+529Qb1Zn78kh5w2fSa8Dko
E1UMO7QTXXa2vGqqaQF0u7yMX0OEFL+9G934fJx0UMiLdb8UnazUxDW15+0rOV8s
XoE0j5QePSI7cnpTiC4HNU/TAAiAV+cFSOC+ovzvdc1G2i8rQ9T5WLoib4KHUguF
YYJ7SEnFsy4PQceD17y3OJOXSwLuzov3mXm4J2U6B6FjpLiPjkhou1X44VfH0/ue
+wjZUFKx5JAnbkBkBFBBP2mFatJUZPuQyAmh1LDfUnksOIb4r+7exLWKU0WjHXTK
eyJdvLCsGjX5hginkn1KqrHcoYEA7v27RDNT7k1WDos+rF2rw/rRXmZiWtgHwWBW
6/bLdt/Agz8nGNZq7hGSf+16+mZ3Ux5c+d44OvTI+GzrdqMfPI28xGXsSMEInfe+
IUlE4D8Ud7EQ94xhFaxzUSQdHUFp9tOC9feoOIO1YzZkj0sq5DmceXWANUYHxR4s
jIklrmrSfxdPHAXF4PxTNlwQGDlJat8FqFYCgRWYSpAWIkS56JzZ4RToa9Ckmagm
uOWncr2UqFKb8/s2WikkiozKHsWZG2jyJFTGggz4PZf1Ruwi1CSCRWILrBvXbFDt
ox9hS3jx87mLI0FH+w3POzr8fBC8pFa3XpvTzU6q8+oR0BlxHM52ma73CWA2Mir2
iODgocmggJp8rlntA4vRoWSlXCe0YPVR1pJEfmeJXRkrOs0N6KsRUMajFrrff+S1
Spd4H3f6JZycnXO/XhR23lE0e7UHRikg/TyG30CfzcfEJv5WCJIwaWKYArc0aLgx
eDbkQEm9uHwFRJP6B1y7hUVZ03pZ1KAh7BfkT074KyEheWA/EtBj21HAf8XeT5kK
OLswFBGvoUtF1uXwv5JCnE6bFPfkHvrpdC6BfgxhE91fWq/Nd3iG0jJza5LvkSdz
BTpPOOZCw3uiFf4kBNPefR3PA9yED6awcLbNyo/InC27rSNRvtnT2jL1AfXkXlZj
trEFY/fX8qUSURq/phMv5S46m6zfWrq47G6LbVJ0leHLe5xRlyWbartA/TjLZZ7K
rFPJoUG8Sq/pI7McWJOGmKBhf11iiOE5qDFxEeHTkr5IhzlHhV5+VkW4VUnKX8T9
oWoQguAOJdcPBVjMfb2kT11tFQjfnDMocDsAgDve6OBsRW6Slesk6VyXku875TbI
fdjRjpDSvC6f6catT2F7FqsaI1kyG2oxSF/kfq8ow5hvcMuf9YFpDOU40CNalmsG
qf9dRgNtGHtj29+0Uqj8RqT7pAmEdzZMeJ1ee+ctA8Ajjs7nE1efUu9Qcb21w+yG
WZbKB/2G8XmsGO2ilL6fmaWH9vfCrxHvfuAxCFHQ9GVjWacD88NK90LinpLoUaN5
CGLYX9lEiHlFK6U8VELtmeZh1NRx2k9C6PzJ6PSW3qXqVamn5wdkKa+riQPllKHG
vcPhZZVcorN28pIooOjkN0PtmPCdSiPsV9KG6q8Hq3NjJBHfqE+wn+LJBtcGFFcs
YmuxRQM+A2LcY3MiuqdvYEOJbLnM9RUog7/q1wY5ubkCvjb8lrHZIjYuCp3khuIM
etqWvCmBKvkI2PVroCtiMVtU9NxCiBjkWY4u8pGeJLKz+PgH0zTfDz6QvTX2L0FK
EjHXDr2EypsHW40vnYxzeAfCIwwn07NfGCJ3Q38shKdLBA4K8k5PXFnhBuxiJx/g
bAb1Y9bLNakU8U4kFNwQtUysUV00/sfTggC7wYTP2/FCMKnkVOIFxchCqdxC3CTH
c2ip+eDAB/Aq2jWKIi359zDdzBOtw6RP4HNdqWBlNPRbg+rVPXrbNt6rzjzUpsGV
mXPFfVzoxk8ioT4ujhRrfr00f74bMj91iKGxBtxojm+tNX41NB0q+zEERUe/2zAD
GNlsjld+92At/y3FE+nf+qddpjUnMDWqMhZSdMCfd8UDSspznfShwTaxw59roVIP
RFGpvuNeM6lNJHPXTWWrADp42YCRavDykgJhJRO/aagglG6+V3pdUxKXDPOteTFJ
ULnIKnIdLxhi6FYJFJwOkK95AdNOM2Mi7poBu1exikh6EcL6Uy25J409fEIh47VJ
V6pz5YUOlCVWaWsnq6d2k5637BB7NmU8qSoI0spsXLHcXpfj59XEi6DzC5NOdNyH
1Q6hPxIXaBbe4LP+Y/FVG9y/KOwuH3ei8x0QltasVKNocs6EBt0EHjwmrq/4d9H2
hdpG3dLRT3WcpkIEMp1NqscJPV8IGMcJx8SUvxbcDt9vyaF08mdvhk2b3NXFze03
QaCBAh3m78KfxMLj5/gDEywCpqSC+J+WE3vUiVYIM9T1c4+lclxpMmXliTHLkBWo
JsQFA7eQ1NpcfT2dOPX9LFkGBjAgWYS4aSKSwaZYrY8GMHSpy/T/i/8ozhF0WyGR
pJgRyPV7j+seHvm333xPnJhj8N4DbzTJekrWHbj+iMZcNcdORtU0USiFKGLvpMzZ
MNMpmGZrUesIfiAxvZxFW65l0nS5fI/aLAkyys4Lcl3jbRDI49fJHOju6TABGQmm
1I8sr65+gOU+HrWQCi9hrRpHF64L6H++vXztoXpCj9VwcDYIwF9cGE9hCmtVCHid
eTxoXw2+PllRF2kSbgxE6HTv3QgIkQTeNAJQ60iyfR5TTumwsZNGdKL7nCngoque
n2chwB8cpzyAYZzaKmcmVmFudmEwzX7E0Ot2MVZouqpGqpAVSIzEDmOhXjTKhfIG
fodS6+0qQOaqoFW/L403DheYDwMnb0cCphtZOkN3glvOb6LZOA2XNc+2k9co64dt
HnxktvQrSFeFmWWPiQ5815wX1/O9619WJbI0EdYh9+LipHqrGk1R6EmmtcTgXznb
PiUkzlplHzUjDVpVII7NS70WfdVl2J4KIlNkRnwNZRLM1iC1sQ4bfUk32B6WXKsP
fTl1roVjgyeMl00bzjjswWEbgWlKjZMC7NA7cjRbZt94lWkbfE5T6xZyhGQ91ob6
waC7xiVJ0aH/SFCANu0R8q3b/6ZrJYC8Rj+K7aiUliHRpnoapjfMWXFYJwICq9AT
f6HE1r1sMuH2QjVdCWE8InC8zZ2lhcVxR4LRc5BEQrbueD7fNxekXpMoALH4MtY+
wJsWDl4M1lLznrcDxidPiPcJH6BSSuYta1tDmNzjuSt2BgxPsVqUd/QGTkuH1fuX
IgZFeZTcqGlbvMIXyZrrT/DzVoVfxnAU9cLK/d655epmnrwrLhQzXf7sK0NP6jIk
M3a3KrERx+2jUKBZD6w7jJxaqdjZgaXU4gUrVYKsjGb8fvm/frW21eCXsPulba1D
n4/rXHMwpEvVBekwWwPtWJPtoCI0BRo5QpKn9IzwUJBUMdg+IXoXVjIQ5VPtCzHA
CKySy/ohxUdwnn6yZYL11rafChsgY73nJHRdCpwHM2UiwaIwpvwKolFE1OBexmWt
AL2H7czV+K6yucsQ1WZU4Rb1qLnq7oofTkLvEu4fo+b53VxFfvN0YQo9xh1h/bQo
0AF3jo1FtZPH5EZg0mNr34bVwByUg+PFH1dNb2g6VP3fxy6xHAmLUUmSMmY5Xd/6
akEdTMOE4A/w1YTNDhGz2LTNxNA4zxe/z0OPbYd60GAbcIgzYHkql44fPBdCJav5
L3N1cCAnJ45OC2YdKGyqgv4WGzM50DIYHGN78txjkVhnRirMiZA8elst2qUxnlHU
VGRLlofanlhNmvhoxhG42gDBOvHaEIxtfo0aAqglxTSwm01oEDsxavzOD/p4TYTC
yxI2fS61uuHirus26Mu7hfnC1rV13/TtJY2KJEmWugyxf+m7XggNo8drLdlTBqAa
NzbAQiySLUCUP3Wwwa8lYywjz314xp1cIQNjy4G9PZCtqorz46qYm5Q0p/Rs1x6/
Rx66hmbEfLuG7uvZaxDaRk/Jj+P19eR6WO/uAl6dppreonLPKwH6ordwm8EwkYeF
/XiXDzEqOfo3hCmwb4mPPJM1ljJZAJkKFd/KZ9DRPn1lj76xZ0dV4NqdS63bOqKX
I0JwjaaWgnL6kfj1xf1YBvSwtO7q5JBh5YRpz8+uAnYZ+k/ZljFrv2UaxkRedElQ
akOJsWYdkuzLKoGIt+iWFZV4kiMq82TArIXEIGZsX7waay2na4AZSPSO8uc5szF6
t44Fnwm9PZwVTmEYuJf5KtJmUne828D0XTdFSp+FpxxHWpGtCHe2NRhS6kTzhfkH
5CacWgAtVxA+jbE1O63egYx+1rkvY9zKf+Zhnts4gBHyeekB1f5eW0IosEOmYKfH
M62dHXPoOlzdZyKfb8rwHTIvIgYWhvAxPE80Laf9eGk7o9RcCjK6ZWj+OCNzkbwJ
J/2DLcrC7EQuvVAc8G8EqpdxcgSoFu76QiSU0CEAAQ44+rwn7dvOaPd2jNpaYfpC
7XmL8RwuMJiMDnapruJiknVoTvEjQUY7fXezaZE60tU5qXJyv6ERa4G76RCCH/iQ
GTXKF4hWLAc1ltx/9LhjcJw1HhSpphaptm23qvB5qyNfVyLMM6H2wqqKWbapAcsd
7OtPbgO/Y2oQkypY8VMGgiINg8aJhHM8uZAJkTsgnHGRmps9+JKXcelF7NWviQs/
qQoH/Xoj9G0nHXNUg1TER6ifDb17pNmRTcAbJbMEfv3aWU7oh6yhcIUgKkY2z+Ha
bASoEvPyIr/tQx+vCzUflukR5lEdf6H6wtMWGm25hlp/yQgF+6uFqsv56USZzZIY
HcZjJBYFttTF0hB23BiWm797DP7FURzXZtvD/WSWaUUdhIm3G/8w7dh67q7eI7Ff
a9bl4VcG8yoxgoFn7NTdTn+BIlWyG2wVnDuEAlYZUhbTQqSoFB/jaTi12molr2XQ
y+kWv2+gTY7VzYgr7zWCpKCd51KkZcRMjZDQ0NVnZMO1dx+/WiBANp8jeN7foJyy
A9vfii1kJ3t64pkGmNtcqi3yZJfDxtkRn4znEVUTGwWUbcvxoyomP6glWI24/Zjw
Fq5unHviOWr+3fJL+YVNLJlWGh1drSbqpanMYykJ5Xsnqkz5bgQQ+iNQZJUT2Hsp
vOz4GpAfD/IEh5l44OUIv4LJ5+J8Z7sGUzCGyKZPlPUjO+jPCiBDxMsAnUqcfI2L
BxqjeeH55Qsf4DqJMgdLODtWjLcIx6cWRdSaomRmEU9OILzfqhTZr51ksHXyWtLQ
baFIkrzg/vaaq+GO3gH7hQP01cV6G0m8b5gOtY2AIpMKmtLG8O3T4xxnrA+pPQW3
FH8rFg5Wld0VLn17PtUSFZc9aayMjb3nuhgXtmHpKkYyr6X4hF9+abnht1enl81q
G1O5crz/jVZj9vugxYLBC9qWs4kIGOXyw0VWaG8wJy6sma2bJcur+TNwa1nQpawX
HPscPSWnYgIMoDjYSFRaKX1YovD/DIJKttdqN6q42ne2a25lKHwxFi4lORhqvJpQ
vfsPNjZe1z8fPF4chDYBJzdPj6eP5QUKnYZMO5J5iSM01f3Vd6+s2c5hN+yeTU6R
Uhf+smx2qMDpZDNYBPPMNQQtZyJhrzP/8oIWFc9rpEWwepHoM2xAIuXn/PcED2kY
8uNha3T5TcfU4A+vCCUKp4f+j6bTyYDmqrrbLYRsNlSxlFVZPT2RJu3cLASPFaae
QHY/HlyhHb4/6dzvAQrJ3a8+hVP5VlMMFlIumO/xWVWlZxYYaQUYYMU/qZov5NLa
QOE5WFDyDkl7MJc29EGaU8VAzd/xmgquVFqo5UHdQp1zdeIHUrRrDMh/4UiDgeOc
x+sV3gdVwReKxtDShORHs3BSp1B9Wi/H5HjtWcTswdumlJe2i19rI3BUFl7wwypR
wgRmuTd+qjMcGIQ+seAZ7REijdHLafENA1A284m0q69+o0dc0VSnRFkp7Gyw+WId
MpYw2D+4P3Np3+CPpmIAkKZSOngzw4b3+5EZjspQRvnimmj3S1mqDbkIS48ZZDC3
rvxhWBkLHQ1469eho2B9pSuyhuF+Tod2oFHYr04qVj1dEhs4PVZvIY8GqvtZyvA+
bh+DT7v/XYANmhq3xiGrLIRAYNPI6xyolIgOc/CxDgvTE1KT6Wmv9OGOrxLv7Gu3
FDHG/ldS6/bkWINWwTvuhsRPQtcc3MVe9MpAqpmkUAZ+TD7buMKwYGL2U2rGNRjh
FGdp+SrseA772LnXzAaGOAzUM+87IO485KERLEywh2EZJO/ZAU1KxQaP+kBtMj2Q
Zw6h4kyf6G++P4VZNS24bkQmTWgBXs8kRJJvNet4Hc9QxQvZrSJfg9+ZzNkEYwyx
opNPOan8Q43sTOLYTCtAP9IJRZF+TMydxBjVcwh7UtAeHpJPTYLUWEC9hq5sjaxV
sUwltqKDSxPU0zINti9f3h0n7gQR1O0P8n6+AZ01G414hKgaAgbm6JP5z8oCwv6Y
WfX+rvi62gxwBWI92PBQ0iw5wreAm4OsJijD/2O5LVebVNHrqYujYwWkvu/oYDny
sD28aJXjUmMee1193iKdgRhDIWR0XkdMf9vjOvOpdNE1zOnJoqaqQ7K9uzuVqHff
W2DebFJb4VBYY7pmSoMhjrfdqpxVcy3uj4WHPZXJKCn03EGv121VnNKEDYfaNDJi
jUWGLhjcNFnLXM4hKKJ9jcsxQNEdhdF5FxYw/TQadGwq2sb4yWzs5d8F1MDRXPNB
nVzF307k9VYPrCR+gzmL5i15KhPAGQAQT8VINuFm60+ZxbmPpzRy9W9pF9PAUTrD
0ub3zeSeNQzHAZUsf4hwSXketJAIBmvynvfRBxS92+qRs98V8P5tkCJk1imt5c0J
QeK3Yng44vjSXFG58GQze+ZC69MpzloQp2hyzWKpPJPMY4DCmMpAf7ImumH9LhTa
tN0TY5+Mhd5nvrP9rJsZmWj3HKaqRl57vDuNCZcB2JoJvL6eO34OFfiBEcgNLPFy
6DqW3e44F5yr4QlI65vRsapLlo4mTWE9tF3HxXMBWUhX/6XhEDqx4LRIJ4uNVBdY
w0Mvdx8ISGDM4kXgMLVWGlPTdetz6wFOu5+O9e2Xa6czUbd4WlybEjF2rnxSnlQP
pLGQTKUdR7dORG5UOM+I/VzJZlBW7i7CXkLBryAHs8iTqNsHk+oPqKqGqs/qld8/
sSnf7idxvmqp5oEqu9/Ed3eD6WlFJHhvuyI3YrVshAnXgSmEoVElUEtNJJTmv01w
y5mDSs6sO4hlJsc6yYfrz4ub2y6+Y8x+WD1GSmW4bmKEyBahbngB62j7asRTO1f9
C45rCaxfendmrXYjvclbn9ua1fCGEtZztYtxyhtzg9zvJbXV/NGA94Braaz5ib3z
edmdis2uz2Q5/Xj1dPHjeP79jOCHnahGZuwmvH7R46otjVQPKFDXbo43uk+k1CRg
yS0SPIo/neZoJ49TADsj3YrRLjP11KR28iyCCFcvsIc5ex4eNe9Ycf/7C4/h+XFj
MLUmquXjfayCIWMm/tDLEOwZaIESa82TL7cFvJF0vu/9LABiUdMqzPHaJX4bOEaO
kDHMBwWgeuZuwEgtvqyYko5+azwM6UgJIT8KmzQcLyuiDQh1uUJhiq1HTMhZbsU8
4/jRLfJKNovqM630wjE5rURgDp5rqoZr+/HqH92wcL85DNwkmJqumfnDZRkWMyQf
jNQcBty75tfAEgM5A5x+MWJssvTYCvjan+k2d2Zq0eRpoIQfIMm9/QF38dO2E+Xn
heE5Ph4Se+fObKqzaPQbOqtmHxfgjO+Ys6BX/tgF41Kjl4G/9qoMmocenJ2oNZtL
TdvJHnAUbKnjFDcD55HpMtax6OO0F4PSTAUjIBcvhDaqk4hq7oDTnpRVKNiFyodd
DqtxAMFCy5jbA73IIelN8RjNmTGHKJ0vCHXpJ2fYJHKg1ndEQqZs9MX6s/GpOdfI
udtDjkiKBIMqkew6jiJjjOoimRPc8di8P8+oeJvsjPUQkAuhqjal679W3l2jnxvN
/iGyoY6UFpP2ajZMfWI6C5QV1YdtqM2yyksZvr/GcYACrmUC4N1P9+eH7fRdd93k
cvvu3+LwdIR6UVG0u2Dcb/TTtBDHDVTxusTwS2WZ06f39ruQ50cl6iKw4BYvpBaa
87kfpKOMNI2NYM0gL4ElyNOsr9glT39ENskwFkVtk+xLwCJevCsjI/hhwsk0nUSD
iWvfB6uyr+Be+0mgRbI/EZu8QkXeNg0btx2NcnyXRHSs9ZAhkgSSe+1NpD+l3v5e
815uEPwiTRC1DaEmE//wSdy6UypNjenngzkc5WU89+jxkuJC9Tb3We1y3Xwp24M5
F7fyBWbP0OWKXxoe43oKab+Gv56RmQit4OG2aFV77Ma5v0khVhQ/YQ7efLKu1RcI
G6ErFXdgVaotoaKDFLOVgAAY/7t7RPDf4NXVf94u6teAgJ9Felrx914HEU2MZVJ4
6OLQFiGFNK1mME1P0GNGutwl2qVlXTQHk1G0IbMORtTbOJOlP+G8g7QxgTeprG4b
GTUR5L0DelRN4JYImfeduwWLlpM7kNcY/kQrJINWdjcE5kmXIgKyq61C95srS3XT
uzvg7I//y162GgmZUTIENJ9x1yePhEDCsxz6XikACtjCY/J04cn5x9Kq5utlr6uU
EPsyBvpCMvcUTRwMTTnf1D/y7rM4t9kBWpmG/AYClMfnAIhit76uEdjNpb20EBpT
Lqb0KoPO8IbwRltSfwy4GJplQCfXDY+TWMHO+oiPswM8tAvFzFW6nXXd9rGPSImL
YjEI1Nfrez85ktsa3c3VbtqtxpQsbf+9+G/IrY3vbuIp0wrJt/bhINKWd1EIFi5g
sx5PBQIcaDn0m8alvCTr7tRkvOf+tFjcVf2lOnOwQeLDVGB62nID6OaOXYFlY/D3
cFMrasPRk047P/SySvkEPnNRK3GvEEClKrTdJYFwwMCq9E0KM9jdkHcaq14gN2sl
CwfcFWetwMZwx6ytJ4pZnW2xKjJm1+qOfoJB50sPLViEwbf+tfcSdJc5rDAcH3PW
gIpcXhVcH/OI6pM8TwStuhMV+tvJtRBA8ofGAcDrJ3zLCe7L8zP3jHsCl3QrcGr+
hXA5PvjMak6+UEixXr/KcwyDhZKnLL6IBFmrjhLvEBxy1yqeI1CfBQ5lHpPbLv6I
iGtP0m1DOmgmer1IavHadQYBQm7LVim0DfYalg9EhbzZVRLawVqpJzXjlPResvEL
Z4SzJqwLw0NYUKEiSUzpoNIWFvzp/ulwF7ac4k4Flpu6lyugvpdnDx8pbrLlA5SD
Q1LF3dmSuWA9khec92E45n0+lQOUlfYZdbSubcZ5xnBRRaWT3GiU+hA18rW0xM3K
VHEV+EuyWv66kpwlgp5quiJVuJtlV4GVkqv8wB/gLeG5lWDpLe4DHMcyrFE1vsNA
CIIQUVd27NZrrFk9TFVTtjOEcIkPLlNWUcl5Aej/6oqGM89Kbvmd+R/1pKH8BGGb
JuMBQbvw7T3lPocZTX4h+6FwrMmMTIbqkBGdfJkx1Orc3DFEYIuZT8MRWyKv3H0T
wKdgImx9Iw/gvaxN3cNZPr/i3w59YrHJMMFs9dQxTBQM1hY/DWjiImNhcaxR59pG
IMJZu1Cfg/gWHccokxE1mjVRh3ldWwFCYYdz34mI3QPAXEy30Nk9pbNgTRWTcTPL
406X6j3kDVcVt4bSYNvZeusIA6dOAhcyB7rMwN+k7NA1WDLXfueqRQv7EWPt9E76
UlIN+2AmVsap9XMHLKqj9pgZRITe+4MrD/Rf5Tj5ENb2lPkBGgOtALP+KhfrgzpP
r98zzLNVLxP8XliTGetkfIXIkZgVHVXbDOOYEkq2Zbdv6HWi8Tnin49dl1w2BHCR
Lo4t5UMMQ/et70OcNY9j0rD8BvflT0z0MYYoYM0HrsqFgQYwM0/yPcOXWf5m6Zwy
IjPK6jBRJxoCpRG4MtYTuSksLXBfdQ/xKlOAAgoZ9kzTxFux0e/oQ07oiW1/h1iW
PR7dBsR9t7BSV4ybzFkhJoWdJ2dcO5tVHwOxCEsCeIB5Ac1AszrQ/ORVkYDFBPeu
nIJ/JFZsR8zHZIP3tqK0weBLq8h71uNisHy4QhDBiOAQz8kdmgvGGNzJQZFL2u6c
Hp24EGdCuBNegFl/QJAda3G/bhJLtDFwz0UInnLTFRQ6OfXUj3MNoEWvtT0QxNFK
ozmzJMjMIU0w8tttKYf/BTE/M7cObmnJXFcq8fs6LEbYGoV3bDhvjxkvPA4dtyJd
0GGbJUteJwzIwWVioZSiNoDplmSFuKjEdRboZrTFjAIJvijl9y1qpkDIx+JX66V7
vPhvKSgDsPJwyIESPhIVSVCe26KN+UUMbiowwxhEs94/ohocU3bAdScn/4LdY6+f
JzELQkkvh80qyuE85yPkmeMk17xyYyQWrwGllsvmFXlP5tJoSAlP4svzpSDUsWJ9
+rz7+qSH+SFvs71nxGJCIUkQYyy1tH7Fyy0MbsdxVLEK8v8x5BLGnjCxtl6aRbnC
RDKKBof/aQ7t1nTnXqyGnmpXbz+Z+pxK8Gr9i+xbQuaFH4T6izC9mlmZ9AE5W1gk
HQX/Hp3YBuaswN07ofVNjyRZdZrKMSjiEAZCBVeFx5zoDYznkpia2IgGi1GcD2Wl
a9q1G0soIzCIZpyEm8JsIY3rl92AnEkigu8C1hWFkMoty4nqX0QdnLHwpTq8G8Sc
R6/1SFjchDclcH1yXmlfejAkwwpi/j73d+/zI+gjmB3X8I4KKieShAuZRShdni0k
Oxbak/vsqp9jXgRbqvLonQeSFNt6UzqBbc96xcbZr5hvXRZENepu6r45qOQXPmun
uXpTSAfupYtE62VgUz50ltbYUOwTyr2t5U78779YWzCqJzDTabhVHR/9Suxka16G
ViUPkv28RmhcXdEs8EyjbMMoGI1Q8RXclf8MlfKEJqU1iwyrZwPZGlXraUJlNRP3
qoig0KcEv+enBsYzOjPlGPt40PUzqW+th5ORmnKVxCAw76AciO99gW3X37OalNbf
kwZkqOQI9ogiCU5iGKUvMsuz77AaViXKmjRI8rFAbp79iUcWUr3EOwAcG4TyotJu
NkHLu6KakAGLDbAdwwBrSv9Ws6tJV/VUupAo+TG2THnveHQ2Hlwsa6qGpqoPPp6C
bDbiuXXnXeD4G+yxyXSvguLPZ10YkuAkBAQxlC96QHdhdXBn60MLjclABATW9Lhw
wAYWe4lFFBabLbqaCkSiCqGdDSZ5BriUORBOItFRJDDeYD6nARCMDPkcJn/JnMpl
JJoscCA/JtnXQRgRoMadOlRFc4u42Iy95rBOv5n0rZda11pf35/zpGlpWM5D7u4U
risnqH8+0qV9QDy8Bw9PAF7RQ2V99pOGvpieUItXtrHXuAiLLqhom977n+a/oGmM
htCs7kyiXSmdpQAgJPpr3XEwz91NltQyJnl4ZV/rbY7W1Woyi3BT9+nvMnUf80QD
FrXMvWpAsnlvAVC520I71y2xnhwtSMIlz+BH1Ak6mzfenHKDrYdxg5egwH0d2Q6X
ova5TWbf1K+NW84NKLr0y7XVJ6HZKtI43vZ0GUxRzFjwXFM1uO0Zq/homN/GCC6z
FwbLGb05EYqHbbd1dWYm7JewmEZyEBNReUgIh4LVczWVpDkoApgoWSDrV2TPZufA
R8yMmoZ8afw89t82hhW5+3do1PY7oIf8RST6TfymAP2Jx+nxkpM5p1jBa+1ceyJS
aqhIT4UI1nEOBdSWTW+e3Ve5NGdkt/Uoy2P/jZvWslBROgEj1T9BycqkkE1uua61
j/maPHhoO44Hhcg7/PMuFkssszgvUjMS2o6OlAufq4m7tWLBTqNAciW3ZJzBL1Z/
enHjBRTJncNKPf/7lq9iWMg+r9GvLPkqLu6TaGuuatVIlTzxiazvo0JT4FmSZJtq
s98S20MdB+nBuDe0SvIjw1+qUZoE9DOGkpPwM6v652x6hDIuMOeDT7Mjnu68doca
tegZYbfTr9yVwAcDFzjzs9ZC5zMsMUlHl23JBA0sC1/fTOcdx1DvDZh6fVI7YAsL
I6kPpqvsWrChQV0lbVUJEGVy0U9ZvzdHvaghxzcHaWY5raPEhB7cZ9YlfR4FmSdB
MRKXe7sOqRYwx1LeddhBsebyjPwvYCthUGg49ErAFgcT+SQEI7vtmxhj+Qyjd4c7
Qo3uxf4L3N8paydbAXfASpvbB/YTJ/LTrgnKWYx7qrowYyLTUs5MUgriVQM+igLp
YMpmzZb09C8Nt3PFXkANmlXQ683dsL7I4Xano0nO6YcVmxRRecvuvANI7HucyOBY
AyxAdj+hD1H98AgoZIu2nVIPv49AZ1UQWRZJAmXTKjbiDx8ZTMg74vQEqroFLUv/
LSmKo+6aehkmajJFl+GuJiZoa0Iq9pXfOOFGbdPjeCpp2C2ehSKdSoa25UAP2+61
uK4FxyVwk55xY+DqDpUqUkgV0zPafTcGBh8Goh/Qkw1R0VKcnVmG/B688ksmyP+i
zOGqO/Hg7Bb65/7rzCYQ4MMCm7oSrZL5SBCRL90CkgbcTD01Zo+zRidKbHI8B9WN
K/NPL3ejdLSdSATwHABhfIly/Vk0eeC1I5N7XB0aPV7m19a4ywoOD+NphTnewiMv
LBX5uj8IVgz3IHHxMA3jXMObsHeRuN/UcsTufAljKp+xHVX+M5yaAysaEOh/VSBm
Lom2fk9P5sn0HAKdUT57BOJgZGsJtgx7GkzZHYZ3UAp5/1TUS9Ee9AsksBpGALZi
05fE1Ijcgq4N1p0zYbFNT2j3vWirSFlpBYu2JECgk+Nd89gqmzGVDk2yvR5OCH6v
9FY+8m6Q9MNIHEZtH6JuBH55JU1EhM5jIET/iQ7lsSsrLiN9+dN/nTiOGyxS+uzC
/GXmz8RgwXkEj5whmcoJyWNhVnN6iHAial8j27uozs94Pf1rTKqINXR+yhhrBKDZ
MfEG/b3B8qZbZ6pFJPAWzAFCChVsnmTarG+8VQafuQlO2C/zmIz3b5Bf6Q6KyYai
YTYwEhWE/vjd23V2nCsaFqtCk5+QsOp6V78tYS9aryg4CjD2lTnAT9U7v/fwMGgS
YxXp8KyOWx8wQUMuI6AA60etgPdjJP8ZFvUe7IFmr5oP5mZ1UP5XopHDiNFurHIO
lARVe/4Uh4qa/vHePB26JI4scOpfVNHjOPI53oEEreMWjRktkukY/Y4i1Sj5MMMm
M4TQFRE5pep+00TKZM9XuPh9Io55SwFZiXgzU64HgZ9hot2031ns2MMHdlH1qXsH
UUiAHZz9cUUxCUjGTpH3fHA/wOzD5uYdKpLgaoNLRqv+e1KWe0G3iOq5zTWANmPk
nZuFMoT3EpLkBzHFGWman8SaTXf2KfiP5C8wmM8t+kRgNcQD/R3mPmcE/Rzl9D4x
bo7UYzlkrWLV1u4IeJK2icPGYbi/XMRhS+iTA5k78cNFZgymjxjMxEyBLoLRDyln
Lo8ruyZW1+S4LO6JDZmAR3kjF1TxP+KtNgjei2DGY8i07POehXJ3Vxwfpy3hy4KC
XoRbgBrYtIDa2WWg3kUCTLRt6B7rnrbIA50CuRcJgo5Pg/Bykv0lIUvL5kj2eQp/
2GRwppYJA041VkBoP5S4q6WLJsSeUejkqvDWQxwrV09zZqir48OnJknZqI4bRkUi
7nSQgfGhqZkcecd01UmOpa78/91cm+lNJqgmqvufQz6+QknGk0SFZ4XrxJbBk19b
RVf7eZyZbWDK4o+nGlZo8oYrmUz4magPNwSZHoey/76oY0FvFB7R1+6DZFA0KUdg
xQgf641OyfmEWVRtfJZ3s/aSWPMak5OiItHQjWuvpFyTg1Y70eaNYQwenSYBjx5q
GHXuqk3YOAHyolFmQJ1d5qHsPSqdLCAtL8zzgF8HTUwFt7ffzp71tSYq+4+ngUcI
ligTpwlyD6tz99KskHlBhSJRr0KQzQgqEIuoNU9QsrEE5aoudLpG0WVQjkEMlUWs
ER8Aaaz+5SAMbepPPGnQjwqmZ5FF4EHb6a7KUxEiEvuHE1ccpV8DDHnRJIKYmlxg
w4XaiTjGO05jW3QvYJVCwYOWV73MPSggXNQFnYDnvLlep5oq3TJLzZ2ESrGO3sU/
Cctvhd0od9B2wNsT0k4kYvOERjwoyeVoeLtCAmfXbrKYYTIk1Z9RbwQxBf/+an21
/40Tq5KU0rmzlJph0B4gybM3qfspGdpDmh2PwrB51r5wHrRqo+sBuNTcFR/zKUFn
NlUEV5pPVNsB8u2ZJODSug13eoHvRhrnuuNtnR4FARtZJ2apFo65iSC4xqcjN9ss
XdekqthF5Yi/cQG6VRCZh/RlaCX0IIcGWdFEDRWfDC4dkprTqb39dt/+nDaY3oRw
NVdNGKWnBIItjo3yoJzcIStQ8frfmJYiozSH6g31VIEZogc9K5yORfPTHwtO6G/j
a6mL3WW2QLVZuGlbh5phFLOZZ8ydVBu7CMj1uC2D127K5j2u2PjIyOqtseeZrYsO
d0QDho35sbu5ZB5x4R+R9dl8an5lywyEaO9Jy1fWZnKqDUdo9kCrTzv9VV/9vF3z
OO+tPMLAALyiTxozsU56y2LA/U8polZGYQdKwy/nsnUYWuuzO2dNUNe1zJonkJ60
vRbFFRKomj7guZ4zhEqKpqr4hdyx7CWtfUPl3MaAHUpgjuQ2kEMh3cnAV1vpq4nW
97f3eNUTGcW014fMC/lZNO+XTgosshZ0ynHp1M5SuTDv8TWqfsSOjRjEhVAFJ4PQ
R3OiH9cNy+eXfArd4OEEwW52aW9KwpaeAV5rHwDLqOEy4yvrapQlyvSgBOE+Or3l
HTt7NKIpTClpDoYwV98+9oNJkVk85RxTHhklizuuzoZgUN5xb8moHwvfPVjYv3ft
RdQ76RLTA+YzJy3bfjT7n3xTqWr+ijOkqv/93C0j3Wb2HFw14CMgV2TuodM6joSl
v8X/MaHjNe95mfR6D6ZMPyzVYl85HYw5B1+mAJV86kgL2yzy2Zo/srqblTqwCU9A
r2DJjADoXpjWpRpfD9GB+Lf0LhrfW08Yji+Isajn4tJ5ASzrthHAt5HCY7AR2PSn
Eb7hZi7MeFM3T42fDxnypW+E5Ll6VPE2+CJHxLCrbqeW1ZSqBD8olLIBh9us59Si
VXTamFZfD2MjF8O6TYFsxzmSWMFgri3gyQ1YZEhOzfJW592tnCbuYhDfw2uw9CaD
xZTxcM1uCtcZtXRQFu2UJqFZXIy5Z7kWgK/4StgzuAXvL786sTuthH4MFhbGKyPS
2f1uKO+SygcQu0pNVIi3ZFzT6t9xMaxV934M8b5rKBQrlvu2hQ70KLRihBYw5z/0
QzetY3/g6SfF+/IRNH4xtIXULflTb7jAkeJqRKXVYzxRvCq+v5gY9R1HKnIWTBaj
pgRioGwblLouwVKErXMD+M60W7BXHUgugWJZ8MaxKQphistF1E/IiPHhsSguc4or
ggwTjJ7zWQJPzWFLILaytlwo8ma8AbIOEWfAlkwYrw5NZlFyJ24l2p1KBWJT14aN
KUm6krBjhzIBya2edQK+e8T7woVFgEs5Be1lf9PNojO4OTnGcQNAFXq2f4F7pThT
sQcRP3XXZr8/+aWofMwxnC7UoZ1Es64Kp9phrhB3TewosBejzWm4R2yo1Q6wWU3E
k34Jq3WY2hBFlUUixOEhtXK4PkE0WxPXt0VZ8BSlJFbq3s5nXPuHu587+rkOCYoc
+dMO3YvEfHE/JnfBWayFb9TSdzD8hARaCIoXDcPLAt+dNQVuO4N97nsEzNAZKGCR
GI3ufani/KYyFyISJf5GxHIih1RyyoGN/o6XZ95DrGtvBkck19AAzpm6McdfGaac
21aAKlMeOuDJ6TWt4XMT/dApyPeC/UGvOr8zHxza6PVoHj81Hi+V9EqwIj6svgaR
lOaJXvWm/ONspkcv0T5Cqsik+jsH31t32aQIwADibjFjs6P8cJrSJE06R8LxV58R
Pj/EzMPNmzrWMzK5vleJ00Na/DDcmFIhu8/Nef//IC2uFXwChYtoNCEHNzCWfhyg
jKI7o7JbyefwycSUcG5Vdz62Sak+2sSkO+Rw+ZzFjaHtO8LqSaKXYr3hTWlpiyqX
NNFp7GStpIYTDS3clikIal3iKeBZO9JDJqsWAmz2IzOdEvdzplaQaKCEpepl0FDA
Z7KqM7eWCytOULOV3aAHtERKN4iFmxdEyrWhuDiKhhKi0B+AHqEdBx1P5+qKDC2S
ZKSIfDRhpiOMPfg2YEHrKGlj1z4U2v8uiNmKqQxbP8JC6dSvZTLvj+RpSXBgpn5V
o75CCKzvQE8I1jnJsdsCqSV9rTLPVLUnIDVf7wiG20XdHTq+zFsy63sjR52Um/VX
Y4C+66ru7FI6+D1AbS9hsIb+RsHux2d9qnvJpP9knd1ZpXKlXcxAL7SNXeY2yAij
K73u4rqTgr+8c8I0kq66jFxNtalwLenMPwA7EHRtMGorAf6/EMW/Ovf/ebBfG+7T
RigSJpX9Demry3em/ysM/ksFd4hl5h9BjIE9g0C7kyX7hSUjYZy7+TLhND8Qz/Ec
zsVWxikO9AncVbra7DUJMp+7ge2Bjp5lLpIrpu7SIfF7TgWtXZfkAySOIg5eyWN8
dqoFfL4FKu6WilNnAjU+yN+eFwaXGfjYwEJ5IPIWY0xwTFqg1scogyNVJbbTSQz7
UYiWSaq6b5ZNnrc9LzuvmsP4pKLqfevKCqJsOQeNchCKLoGKKYOdv1IbdAZs4X+R
/DEa5IloKx+TMarrwRDKv+IpE5EmtJoGfFEIzf5ltEZxUkP4MSg7dOMBKYrJwYtD
EjZTuIRIww24JFr6CYY1kvLQMgzaBSAODfSICep1SHFn/LhVxuvFI+p8+/MQ6B53
+mUI0fvkE7bHgBYbN2Mf5w60ElJjbjYCDNlIsjWCns5zPMB5p9v2U+p6gZxwEmaS
+UAIZM452dqHwClcpgldDkgd0c/j9+/r/OXQAXJ+3fsTEAcF4tlkhsLEqb6sv6F2
CHcXhg9mSC0oJQRCtQy66Vp2tRwnM8hR7Qzm0eGIBcfg5j9KBOSlv0+mwZF2FLqR
mHyBT4R9SW5lNxoAfXHQxUy4I33pfijDj7dbRuIa4o09opDp2kQfkc3xFmQqgWtO
02UtUsIh7WpLgahpvFFfy+raXkC1H//ijBNDcVGeTO57GQX5AkHRjTlOUVoaVLmo
8rOn1T8rxDf25gcLioEnXmi5oM2dXJP3sHOO044OS2LnHSLKSoGNKKLeW+yyD5uH
xzh4e6atKQjnh7bZKAmHwR5Rs5X5C9sK8Jhy597Hw7dGaykuMxXZ+BCSjVS2mNH+
CnPlVTXS7mybk/ofcCunGHKHRH28RZu4c4J+hm+j4U+tbQNZQjjWFm8rSUU704Zf
48Tym0RvzhrT1O6xsuUdP3S+EaYRe6neFxtXGQhYwt8Ta0V/hUO9od/OG1Fg+EDk
nC1xhqIdFcbr09GWWqUTDhUwzqT6cE0ca1ahn1/NXSGbKlRhRgApuLikoqJQmxS9
saSOjHeGq7QG82PSaYNbyLPnwO/gGkBu6h9d5qZCzKqxjAywbwXacPEd505LZ3FR
HFioMjK4zFys7u45YQLXYYazGThDQJt+b00jX634UcRPR9WcQgCC64WKOJEPeOVO
WruDiydPO/45Sg5+455+ZCWFJE212JrJG5CMh+mn6GLdpASBg7bo6E1OqIbwn2Zu
I2uFb6cfvit9WDMEUcVMfQSbx/QU8BIZJuMqKKOtLdxG7uFwP+o/4dzWsPlSp6R+
Ey7tllyEBV+nMXguijsDtj/9XQoai0cR3jG0Ox2cArrluQqzvHKs3AYUmECiArAJ
CFbzt//iPU6jMr02w4mq2UOFp8+Avmg3T2DVe2ZOL8xSYcDFSVbYHWEHbChGfsZu
WoBsmbxYr5GLmSw2Lk1MoBiOcphFxsTj9k6GGxzKmB41GxlFgG2TVn89ozUmdJAb
NP/wmu1auG93LqUjqbUja8sOUQPR0qALAZAcvJ+HIZH2UBycmt3BRSkwR6FiuDhC
DuLEiWKvTW70b9KCyET0Iavuvghip8X+f2CVFBz1bkcYlxdJASj6AwQId6D8VnVN
Cix0hSAvTt8D9ZvWFbC/jwi+9cbqtZGXjrrmZacCeONy6+hlKbsSRBwqIW8ZNduq
ByXL/Vb5PdLhAQL+bM2Dz+enFrWu9m1RI4cuYONGrtnBJVW6Y46IaY8yFtTeVCiC
HUcw6zAnFyNKAVGdCew+5A1pNk5whBhVFJgx8Qa71Lmi7SYLyZ8GoykqqnogGnvL
WLF6GQyHiu5W4dn5FQ+tvs/rQR4GFwOc3bqXrIHKRr/ACpKlvQg9cUvOr0nCpDik
Wv0PpWy/AtrBZVgZIYMHxsd2nWJoPT+XxKhAyhHS1b4zqnEcucJY+H8OdKMMuPk8
nfEfuEEcvD2eRi9KY0XfMjBlziQrnnKhpXijRtlKuBMgNU61mw/wtePPpNu3TAwU
G8oiT/RErCYCII3B51SBSRXeh/aFyspWqrMY7oBF+PN8mkgfWPjGJwtDR3AOdahi
jTrnTzBFq76gQlF+hQTW4486v9cnesBV8N6Gz9SUKLVGiMY50fz5Y7A2SOjXk5IN
pon2rd2+eIfYk4ZdLtYoyUIcvku3vY6qlpTRl0cbEz46Ea1dbfZxFuynxZe6Wsbz
ZbferMSm6Uw1BRy3lTDehdCgg5H4+Nh4Cqo1tjSRH2SqtuyTBUyhA5B76nQqxseA
NWodEL2jPcEwRtC0WeMrrbpGCzny6TDJjD3ohuDNPp9D0nAabb3zAxM40JsPtKU2
yKHCuoObOzyG+FMXkq3zaoNmLYNkzaNQPzpPbu7jJMR9qB1qxWCDBehqW9V83fEg
ikIwo9kE64UY+y22chsVhEJTG+2mhPXEEJ1AfCnVw3wlGWKkiXDONQDirwbW5QA3
za4UxrRmZj0NSF8wE1+ysjGMcb8sW9GifkTCl1L+VzFj8/tB6ItxECRSq/t1YhXB
HznZPmiXOvRi1Ratjgy0ZMK/0aVZKvcn1ba+RHadvpFtw4VkCWuEhDOH9Lo28P7o
Ga8T/w5d+PSMqhIsl07JZ2qU1xcrTB7ztk7fdd10xZnFZJJuKEHXEdCi1mREgYtz
+Urk43NbVjy/Txj8N/IFBvdmldCQgC0UG2qUc7HkTwflI17f4mzl5TFeYvG7B2KL
ug2pUFfoOE9cK/RC4qQaJi4OlOZ8zH1yqo17T/XxR0pgzlkAqXVO5/LgTXsrkXqH
Zt+j0oQrSK7nHBNGNWmtTHcpN8W9VfaDRQTpMHwjHKrI5miTkc7R6R0Vb3Sf5toe
7MK9hJW7QB7wsF5idZnEnDXOLojoa4I6eVs7Ns0zuLIoB9gBEvE0PL2L+pmIT3Ef
8MiViNsoMbhuUw6D8d7YZ9mtOf0A/Pg13dGhXlThfwhmrSInqaSUpS4K63TudzV4
+5QXKjBJFSStER9FOvS9l+1zBH+iQnDhCed8b9SKjrp0xnWIlStkfM+0X1ZAEr4G
tvJ4VdEXuzUbUYeFu41TBynKi541hbi51B+FAoajZWJXyWwv5DKj/r6/3Pus4+wD
PMcGbRPoUOr91YoEG2v85FChn5g8+Ti0K2Du4Np+9e4R2EjBWTSuK2SfSMsbEpyB
YRaXP5gkT35rrYnP70otinPuULDuV/FTQQJklydZ5XyoiItCxFceySSsCLJWxf7D
RCq9XpO0iEm2ByF2xMS9tZSLcY7Z+tffqb9uUVobHXteilQ2d4x/TMkm9WN3Yywe
C80vM5jHD13TVp4Ca6F2cwJLdfy0vi0yAKD0dG/2S9oWeoCi1zk2u/1Y7PjV5hFk
LLrX+L3njWakZTTeGNOpM6KtIa6AH9GZ14KDZDv9jOA/g4Rd6XdPPulTW+7PlKTe
/uE9UUYm5jGV5hiuOJrB1WV/3yJ0hIiXv1x5vcBRLFTJ+q856V0+bXyOgB83GW/D
PDypSEygueFd6n0VOVdoWG0UYHUDPdPmqbyfkqhZJdKCblLDsQvyaucDxhzgyVxf
x9k3o+nFfy+IYkiMP/UOosIUBqklm+uGu1veW4SLy/iVGpJqvSBfRkCGgqcSIXu1
sSEg6Jy5hwMvhdeGByZ+Bj9VkAASpRcU43EY5m+sx018QFXmgeId09EpxATKQjml
9F3MNKU+f2dJFabgwLA/dBCF5sn2zBUy5NKR69+YTGOvYNJIZSfdGHfroGaKCAi1
NCpCaot9pynMOOn1loAPzi3lbmAkqt9ikZLVm29iYj8NniW5UaIx3MB2OFhKRRP0
6m+mCffYWQP6WlOj1sb76a61N4skYAXCJMkdX1jos58MPj6MGB1OLX/xsb4NnsD0
5wYee4kT/exIXoQyNiuLerlyyGWv5N8VpNIMmddUYU9F4igz01SZfSs1y+4sg3pg
gtpf8kM+TrAkkn1q7DtzjBfLjxxqQ0AADJqsaWQONuHPak5GydO4B/k58df6vnK4
GLYJnMpyDF2KYv9B8Sa9hzf/HtVJXXpCpGcJ/dVqx94KTq4Zyga+RTGYJdbIfwuu
KFSIslHyjJWPmNTFt445thiF3sZcgzavAHwDvqadh2KvXtnn3wDgkmSoRLzuil1F
nApvY/+zylIoF1wGOd9MTZ0agh9NTMZIsu+qoZnyaLqIT6dKK1z/P5TUuS3iuGuN
e9wJiudzUM9wsHr2EoyK+IgsrLEdA3qNgWG9QRxHTUxnZaYya869uYKPO3KLlztx
wwVEbRyyoSLfYo5JUSdrnLKuzgnKLY8yBKsjrUNjXmT0e0gJXnQifR3+Df1ij8Ic
q3RqYqoTPlwokABwy4xBAGc2KCoWF42LaF9nMLkTOP2dyleLMOeRrBRETccmGC2f
5Z/uowMvccRW+Tj4jL7Ifv3fldke5dl5A/Bkk8bUEVQ588BOsu17lfQJwqlXsJPH
U6VZGLdC4ug/sm/fvaYsFkY5DW4+CddVCkKEEbjIAk5kFMgj9DM5pKFdxEB7+W+w
hvFgj2rIgnPIy4k9JTOIKV1L/fCDlMvi7DJ+oCwh1Jrx+2AM8FT+7PUUL7nM5dpl
5jefbOb+tSiw7CmuPL6bkju+roSX/e2ZDumAFihwXoaWjlYma7ebSSk+SCwvLHtO
FYNymqxbaN2TyGPpuwtRB86LG7mByP2SaXstGfjBmP1BNPVDmt6RyMlm/GXT9SYj
CYx4PZqCt9lYEfJV8mgTTG4irnN83f589vDH6uqhxGTdy0IGf3PBnSzzK/D/WG6g
2fOQ+NXkmcDUwb9SbMg8jkzQpIEnfXeR345yw8jUYqQwvvrBZjO7pwOoP43OO+FS
+OYGExQ5CucIdVttsZ0SUNVnl+r9QUgpDD3z340cbfqTVNgRgHqQunos7BSMH1cC
CHhyZ0/MdD2N8+FPGqOhKf4eNLtay7fw/Ph4tRJYt2XrULXT+b9rQgNOn+VJCn4N
nYIbqg1XdGAybzRFVGW+4xTCZeaAdrxFCBkVGXnhmnKZoAIyOUmjrFaSZfU0CH9q
LFxhBhTYF4mrU3DiftSLk+s/77yJeIsQzvmXY1m4imO8TAyFifWaL8GikBbZ8mBb
1gRLI/hyPEDV9HDkfiMyvHTYPrMnILL5mhFOG74ex/YZEZaQ+eiDzBYJidzrmvAq
/9ePVPNXY3AZQUyjOMZazbHY06j4uLGHL6ohptzvMtch9vxzzuXBhZG8qpdrA0vl
IT+Auf5KRn+ZniWhxJAJqPNPNWGxsc7XOXhUDKdYfUlZ10NYXZTi37ld+s2lrSKJ
O4x0mBs0q69DCyzT83KbUUc2QNEH7Fw5aZpeea7BuV8Az3tVTNJfbaqX3yuFJiXs
j9/OhFuYnKQkUQFGWtss6JrK8H5VJ++d6oNaHvIUSMgmiiVxsr9dyo7hmYb3EIOY
lyeFJoIO145UN3JsHHLjJUNGaoYSfrnGwvNGZKRA7uMfuGKB7cP0E0RSApvslVmS
NjG6hvknOVnFd9hyRPMlfY7uV35K2ZDBLPQuQ63tZ7/MYO39Pgx+yr8mLVjdMoET
Ff8iSV2YbIfOL6kacn/3WBBQ2rg5cmQjtAB6qR8J4Zas/9peWD9OrBaLBVCVM0dg
yBN/h9rHgZgX0dbWyaVRTkJ6tfjz28at7hN1MC7lde/oodbB8cLi1EG8LChY+yEC
lZSJneMXXR0x/HfbUFFcC2O9HfgVvCQRR5E06YsHJme7AIm5Nbl8+5DYTLiH0lbZ
Qexahky7kRPPVv3LbHiOloBwPqtnidzmg067xjESl7oNq8JkmhKJVmb6Gdb5A/eT
lnPdCfKrIygwo2MCISst0wZUbftN/JAd3eHmHCihD9n96EV1vhnDkJsWk+xOEBni
IssKT1zM1TYUQCLUjQeFiWjQ+l9UwksBN2LNB3TQ4n77QpsrMd2dApi7nExCMm8I
e+Rxti0/I6Cb5+WJIQD3FufDmRlx8pn69yvB/c6tseMGYxiKRAkQjJSBASQi6RTS
4AyMCFW2bfE9SsIHQFLX392BYZ8P447dQpzbeve68zoAYKhzk43VlFYx8SDcWur4
U/wl4ZXy/GSjnqeMWdmUREKtZUnfAUqYCFpI8a014r2Z/TQvdD1TZZ/h8WPVRQ16
+o8d4cGa8seDupIop9z6wZeqEJrj3VaBWljgLL8dFbKuicqO82JDpmmybtEN0AJD
x0D1g5Zn4EBScwEv+j4HORVj3GK+R7CvkGzczSL9EA9cYHHWxIw77O/+I3UwOE8Y
SuZdQ8BH44fAaP21sJCVM8GcNl0uYeacBdHlOZg6F+bdcAhhbqU1LmmL+eSkbac1
h0iy5WEM7fTrwSsV4uo0ETsaVSOou51JYkd8DtSQ/TPwHHek6oldPGgi0UDxZ5yF
NEJzrQ8PIzX0QvsOp06glFo8CfEhTTD0MPym/r7DX5YnLh0KJj68rQsfqN56S9sr
wprFeWCMgREYt/epfx4OnyR6JNYhccBapNo74uPG3yrcc0agdr/ATWLqy5YKrHwN
xbPAhbe8Vp1VuN/XzP0O+cEfKpERwRneMwvqmDRdEpYPcXxMiY/N2OE498Ek2PaP
fsXYuxPagGCFvLJmmcxMWOomASWJiZIZOv8qQ6n+uOKvkOB7eMzwu9k1H216pg7j
Q3r7S5EuZSRNFlmdp2W4g8W+TDSM4MV51ISm5zBTTUUICpiN5uvvuu/KKV5s9rvr
pQJsbY2zt1GejZZrKbqUmhq7mqNsussCX6lAMeQoPaVb7/hnJLn9q2VUplNJvDaA
GaA7oQwzjiaFd4Zv+vwJ/2qFnDARCqOP5hr9AX2YLg+N2S25hCDshi1k7LLflsOM
iMAuxXCMia7tS7CjRR+xcimtYXrq3n+m4NYlg0u1rjQYDpyktwxXQBNe6HFmov31
f3BEXN0Np8wSpavvbkuInORFt3oQduIqdwhlVYcy9jOWkd+eqA0nLKFcIfhaD0oP
xyfwNHVmM816kWFU+r14Rgf6RZiGoFBOmo0soL0ULKqpvQ6wiROCRuFdUXnX2HMD
nzj1HwTAQ2sQguXVtW6qJVZ8gVnjb3zljxZxk8VT5Mch+IUmi7NmtS64w6+akaIY
qfmIO1n6tJaXLLMP4VGWE57VyeyxA2unpGz4C2SFEauLI58tgDAD1kGwwPY6dEjV
O4+jOWs170i+KWPOpo37HQxmkzGvkKQDEnROBRcQwVTJkCMA0FX8bkdvMJv5brZH
OBpPR9QqgI7lIxvbaWG97rKaOVxz2uwNWeYWTSP8aJ5V9MycGRWmD2eG1v9H1dOV
KDwfoj5hcmKr6IiC3MsIdoTMbetC+WLVvSOoIAURMz2sLfwHJiS6IljN5EUBnoXJ
IJvtP3ZoaPyNADnTA9cLKzzYsB3P4ST1mccaEkpg9dFdYRxQhbYR1+drJfRxQR0o
7OA7AF16jMwhkR9toYq6TAIImoJb7Vv1PK4NiAruoTI88hnhLn+PBbLPqTKzrr4N
6ihiMHhewjoDBsLUfNiIuOrfFIAZ95q/Rrs02pS3QISqhW7nCAiYmBOV5p+OKmk/
KbvDrYOCVuo5Ykwn1ZfVmtU6daiaPZ8+IaxQVXbDPl4Mi9X3jw03FOts9s0H+Aq9
i+d4p/cW6fFE2rwIAqqZpkJFYpt/SRaLDClil5WfgD3SNlNOQi/uVYDDaBhQN3Df
rZvD77bCKKZYaY4QPGeJIIFoQvIL9QZD1WPeihk0zwfsP7tdzD19nPtAeSj/s9/8
CLsI9FwTKrPH/rJfqo/qzMAn3b2bD9rx+sIGECDP0ctG2dfN7GaRmf9Ye0vmhWEM
mhSLoFx/1s9LjBgLjhLFW9imtLMaQ1m9QT+oKCf37hpwECFbv+4pIpcxOsVSgw+y
EWbctHASZwnOfdl6IrGCDmAbvHxhNcfJFPAdl7sBsfa0O16WjU8P7tymH5p57SQZ
7hw9ZTwmXnjNb8SEJdtIIKxnQlVBobICyGoovRl+FjPL5ooawYBFM9nyikUph8iU
gqVBuLSuMhEFlt1FR8wFZl0eNMtcFiSCrEnySAUbSyKytyC2o9XP9J95+pNyu5j7
0heKoXo01GqeDQC1Nx9Jheie1rIO1iinnq97hHw9ajrwJs/qXFRIG9bkHsRZ07Ic
roWbgO0IGPvRwZTh2zyJuWhzJw1EZaeRn7xQhFFMV1MLyQz9AoBJTOMZgJJGeOTo
80xjD6c/rWsEUjMkAhvyyJBtT1MA7QSv92jWss/pbwyWPHe05/zWLKFO7vUzgc9k
cqyKQW+kxzBVLICQJi0OWMTyEbiNbmTfumx4pHcbczj/GztDyS5rSLKMGO1BVBT4
TGBOHX2IMn6tZv/u0J/N7NicsMJhsAICtiLgLkb+9U/jOqDJlKtIG54STN1CwLdb
yV0+AkxpuuNfLRNyFDzABNRpq0ojaCd0X1/4gQdtlwLzwHbQotaZfOIfqwR8Q4T6
Pw+w+MUVD0wP4i/l9qQ1gFgoYjM4/6RAN91Np4m9u7NBYuYNr+Hfum+iflb+jMoS
E63Pxr9eBwjGlCOzb6uBWlC15zEGWsHiLMzl3YCHJVZY44vKCYgKOorNzLQ4fKYM
DsRTA/dd93b92lvxFvBOq2BqmGS2MCuFDLSp4NN9neE6THpkoN1CHvk11ppIcpgD
XR9T66t8oqumWE9r1HQ2NeWuVYeHK5m8+Qy18fY6Y5nhDCaxvT3ka16easLZGIBD
XS4JNjZQFAQvTQYnZCKSNOAZG5kvJYD0MY/xxTaHPAfWaqdlllJLli5XOPwkcSEG
wXT/BbQfzJSj2ZUpE+UQcMhMUQrJKplbXEQSXtQ3SjylwgMMsiBLdkMTcUOpwHp4
ovT6lUQrr3xk4YLBglgYoybxNRDH54nXhnPjnXEOqWorH64Ssv649kKmBM+SN+Ul
wiVFf8YB+mypkuIADjvnn07uN3rrr2l6ACftWNvVBQ5I9FvCRnykqO5rns7mS91f
jCH2C80YK121b1vCV7KrR9c2X1eVcBCTDihNenuogsRuxrYXVdrA4igZVnM7e5dz
hCU988hwZfszVNb8GJhGPl0/pPDNclvG6w/kgRhgvFvbYqCPtYvxoqZshAyCOq0N
VzhDysJwBWIBG4rLDpfv6XC+8B03u3Nm4wglYU1BfBoDG63RBAltlyzPJ/bbosMQ
ZJJGSURlxGCfOGbmyH3IU75OW38CdTAdJB77332uue9rwFgssYqfOtmAv4ahrXwF
Kl9Dqr2hEpkcqiFzhPRPsRxS3x3wl2pDgq4UasXC8gCS0G4T34+M7aFbbfOFXR9Z
YEHeu/nzC5+l0hSYNdKpwBMxKTqr1SEg8ISwdoJZHdbvl/1W6em2C9wr6u28lKqJ
EWb14E6P3PzbkGJuOHn0iIDllJOFmnTVTw3xlNKiDlJEcaOKapxHsyhy2ogqf8Rh
WQ/GPabK5M590EEqcODU/jWS0SjNSUVmilG33p/gwtlNW2FvwmfTaBzx/plmGfvG
vaJhC/TZaCOqB1j3wnKQx7sgxmTdXWqnaMbVG2sm9j94tjdZhjL3NsrljDmZ01qE
UDkHIc4G+d4qsNkHNK0yIOZN9APVCvk3mmdo/z/69dGvkxmyb5tm7ICumxtmJ4XM
E6QcSue8Au1KGIdL6me/vIYvLG4SQ1Ih0ksbclZt7uozdDrxP9rriLBxHp2p4gsz
KPQ15zeVrborVIu5N5INxo6o1QRPJzziJ7viLbMRohIMPOL6hvvriq3MF4oKBt1Y
L83RwbHw/kcPFAyIhd+Uhqo7izS1KualQjHmTLxMKjQpmvYjyHNNkfzkHwN+Aetv
e4SZFU/04cBucLIPttB/jTIvxqh/mOKFcb+mNAAQJDjYpBnIExmQ7XH967IsXDyi
R4c1Elc78LAzJbiYYnHYyMFsvv5C2KMfXY5Df/RuC0eMDCjPKvTg6HdOVhipWy3N
Yf59dFCFlHfHdvwLFngDT7eMwJBscnBCXI+QrYtZC6CP4PS774a/tR45zw6ePr7Y
scfINI8Vdh50ui3g6x/nJx4OY9zyjsivXPl0UWe9QPXZNJ5Er3xTaCpOAOeitLmf
pBpYRz3T71FZIVKPkY9MGgC3ODRXKM+UrPO+xE5R4Fn2O3p+Lhr4YNDmx/i5XsFl
q5BpkFxsvNoFy+XGcPzcxWj/PoneNbtQkTvAz7F1PAxsCWRzEzzjXzLVF3b+ycrA
8Y/83jEquHQnqCx56uh6MImnfwfg65ehLO8BhcJDlvniH8s3rq0rxP6v2OQWf5q0
DEcuIn4I9AS2v2lyK+H66Lp2P5aXulYe6O3QTfn+oNixjDtXKhfDS1gbGR/h9LsZ
jnsJrdQFjKibl2OiTHU2WdVfiWrqFLWtffZwGKEZrBNQ5jaTDFGnOdLrcno2SEvi
/OMJ20kq6PH6TTGrWwlcvwnYpYFCdhmlVvTl3QuXFNkO9B2DAlGKEBgPat9Y3SAe
JoBniQSP3lW2TydIVsOxkKruxWOrWM87cMYfyBxH7rs8TFqWyBM794gBp5qw8bWA
J5jXTfkYPo7WSkCgiFMKUdrmk7kAyjzX3SD8in/Xl0HYeco3XMPt9xbaNNwechF+
3ZgZMg16qBoHqQWKCOccR2FdMRNjUM60P9daGCBTP2Z2WkhLwP7UuS2wNWHu/Mzy
z0s88o82iJy30GP97g+DgwyujspePJjAthb/e6/QN7Cfavo5G+SRsnAe+C3LAmjj
unKFB53GwrgO+J3mLSb5WbhLzWkrV16i19pjTbdbVuivnY/6e6rzWmjtxw5ecUXm
ifjCWJsCXkPT70yVmMy2EIoKzT86PJGeFbrsZXauSiMdUSKUebKtx07zgPEfeW6l
m4qNSJoh6iJLW+nkga003Z9ECV9CDSMIFhdtE3LLTwmefIUUeWBl9EFcHWv69LWo
vv5KqmB4nX673L6BsHZFWo2DY+h4qZDNCGb9o9LE+8sSbWaLUkeKeuXAqWm7Ko8w
PqvOwdisYbJXVMDDa5kfrgdd82u7/eqfOMThql+Vx8c3+drdknjPuy4riAAO6sbe
/JX+UiQvNYWps8UvTnOSmDG/B7CQr6Q3GREj8MCYXf7uLm9TMvi7zIF9E9uJPexm
LzPHNLNsHP0cQtspLBACmJs9h8xvqiFGrIWCB3Ji8c1+xgOfq+ctKHjpWpK1MmMt
XWxAkb7MZwW6rvggx5G3S/0bBu3JvF/0dYYxkHgoqO6tkuiMg0ooTYGGViuXNyaK
3/x5p4/7QDnjRrJHiK15x7nhL3oxNI/7InTJ4O3+YDejqS27KA6+v2KMbIHw45P/
I7AX5KkAweW6IJVtBo2ziDoBZkaRcDeQhVuPUs7rvn6YOpcNhyxxoJr7t4aoNp86
WXEpBtk3H8tznO7sor5DPlxn7WGdq6tPY4bK+rzrty/LFOkov37lVP1kzhjSDpnk
ZCcx5ihH6ZSVt222KwuKFDKMkeoxfttaMAVwoWZAnfg0Hl2i45zzKp18UKFMOVFZ
8DtYTfhgK8Y2uI2g9xn7vN6hosY2D220eHsWk6ZeCzS9FfPdbXfIPb62Ho5WyKqc
LmLuVOdjbHPmznNza0n93CkB+5f95pTPwXJSZLanqmmMHI7MUOsHaFdSQGFFgesp
bprRLYIR07ELagkx3aiN20bPYMFqTwZSPwCTe7kxYR5aXwgs9q3l2WOgpEF+dzUH
N5ipRuJOGjjUV6Kzxu82v4YTpPIoQB882D5MlbQZAxRQrJ5zzTvfkyua5SwHkSHD
xUcmj21XDqTzHWKON5C6vFCFv93WZN0PfbR6Gm1yuX9qR6dmmN7W6bfD2dckr3KJ
pLM03HF/qfeN296QJRZFChNmxt1tFqxJwxK4Z1MtPQ0r326jawEA0F9cRPcfOuo2
okRtnSPsWszrOLJ5YSAFUJS641wGFkcq4g/hmg9AgtX200HRD2tLcZdiKSEH/btH
uR6OFLRvTc0SdjPzkfL2AJWXS4Kxfd5xp/IQ3DDu0qaDvPanVFSxsseDUr3Mm4vz
ljKrwL61pmgmiQoGw1NGwAiIBZMPvw9Ua1hNsgnbb8yudh4eosdeDreT7hk4FmVR
REPzotfYKIUmLaZAlgPM2QKD72LmS0WpOSdT3W0x0DRIyqW/LzFbPys4jaOzWaLS
Gg3rtdj5OkPCPQ1khhnpCZQK8p+iQcBPqF13sqzd/RS4I6sXt8x6bElwDAsv2p3I
Hxl3X9BGf8+giT4QHpzGVJeWDMMyiH6Y0i7vUzlx5c6VjFsn1QMWGWGA+/uPGnW6
6wr2Etx4ZE7OnvaUzc+ABhVjJ76E9o8xVnxROFomugqv/62zY+Ve7OW4yLGEA1AL
RJSwGZeyys/5vjvM9WCqNUq6PiicspY4DsfB86JjOywHzTtEcfepOBs/z+vZFePm
gAv32UUVXY5NitSxu3qd+iy4GmykQRm9LtylDUReMAiwTaRJVPRtXMGzYOKttpwm
4k2yF5dBWu+bdqB1LwHC8JLpzinHyh8NAa6NRVzVIZY3gvjVGkewMVlN1MFYkSrq
+MprdEGRIZV3T6UosFD8x7eyGxxV+QRhPFAvx1ToBiSWHRcTLgvIDBJDv7Zg1TYJ
R87T8riZcjiVpZT5WijW0X8QNO5P3MTzSDRAjYmmMKNdsUwXWf9X/WpXr940ZXh7
Lu7e0g1ewbCWE8I+xDLs4KAmqKyZocACUEjRfMtcUp0+2ClqrA3C2HiI6vd1pzYF
rIamcrKoZgOyu4QUEc6xoX/EHjdhdsgSikh1nrRkcIL+u2kqXKZNj7Ma1x/zFsC+
zQknKr5FK0gVYaiZS2Jn3W88toThf2c4fdYoLEr8fYdBU1zVylUc/SI6rw4WoWb/
aSd19RyETFFXAiAyMxJkSN1YCXvnvBxwNHhaP9SLB/k6S4gbJJcnVo7z/P5edy6s
rAWANvSTAPi/xKfeEmq6nnSm7OSGRHZ00QqJ9QBbhslvJNTRQmim69KdY+w2AKtS
J3LeO4+Tix5P2hQQF3X8YqFhU2oKAmFRyyQNwWV52lUOl43AC/ZaKkqnvFaBOpTM
kC9O+rf46+QUjrO1wk7TeNIpdOoAV6mKTt2kNh6qds2/feE86fiNNuZOMd1XPz+o
6LGXm+iZqZ6Agqn6IKdiH6bQYkNckgzIiX4aFxW6Fbop+2QOa51ux6ljT0dwXzz4
Gfl8mzKPSsNJlkX9tyoRrxuU5DVtmyJebGIoS8mbBHc4ZRh7vVdezjOAzNuKcaM4
VKLEfcJqqIvCcXSyqT0qcO24Xe+y/Ip8RdrCEpafyIZwaJQVmDRDSpy5bSUGYyEc
6niRMUYrBse8dksPQek4EZ4/I5SNIsYhraZ9ruUFMHu6Ly1XZbTyZQxj5liBPEr+
lXpJ6+4f72itKBJ4eUK8ClpbVTWkd8XcWS5Jp0UKr1AtH/Fo5BQg7xg59KUuAZeV
tMA1/pH9FIgHACyyxTo/6Bfxru4a5SNzJwdfcCYSNcgp9bBawaYFLY0gbKgmQkK9
pBvy4c7zE+9NuWuXcRgDGL+KfM23ncSugCzx71cNLteIFCG/VCi9oa562cFBOjp5
pHvgOIVkkr7faIRSt1epSNmBupg1veRghv7fxZUTZTOLkLkjCihrP5DNMC06xuQj
HAFag6Huu2cqcYN3pJ8WLPhcfby1gh+q+LgiFIWFvLWL8JWIVYYBEiwKGdeWZhbP
RBuhRmJMZzM2gq0Lsx+qMkhQ+yZqTbv4l5ntdB7pWkFaGRu57u1PVri9vynb37oX
epRa7831HTS5UZzEP77xOkVZ1YnQ/5D4y9QVa92jX6StLrGhduDTo7PozRpx1sbs
BT/EIcVHlHVl9XSdXOUfkNwFw5ZLeGvgfpQ6fp7bBVhlv01W78bPZ9DIgj5p1ta9
qXiML/vwW21m/+i0L5vgrw21KIyKJ1OADm5zAd8sX84nGKl1466YkaNOyO87/POv
w5/ml8JZmwsE6/70yfvbjJGgWjQIRrm/f5VLvXNQxQ97jnCRw/+Z3qRRK1t27Q+n
F/wqxBRbgPm539eX0f0XIyfmJLzkXj6rHr9ikQ1EScyXDRfk5nZteu6VZDTu0ZnO
T02ZDa3uHr1sxfY/rfufT8umDX8yB43+VunyeiZTVc5hPmoVbrQFragFfyYYLRdM
sDnsQ7aPgJw1W59UDbRpxUOeCc7vlL4ztn8o7DVlTy/jZAvXuNMKit57DOvo7pZj
eSZH/thzs6Scf62euB+WPapaVYZZseh+eQMz7mw2101wQmHwN5bd9uESH6cfuZcA
/7bvPYwhDMgLPY8xd5DugBDcArN+muXY2q0n2u2zG+VVLyshWe5o4/3XF63I6SKC
QIAE/YT/mnN6/XrYMsl8sJBbnr18+sTPJq1d9fXdBYyX4rlGNm6GfevhgDa5N7nc
+K9ZM0RgbZjF28CJgRPD1KafZyDotPyOknN0ousCPd0VsK6fs5UjPgmBmdL83/cp
NSOj3cXPsxTLNK+kkqfG5W2HqydOSRUYSot9BsLFMLvboWWRX64EPcaeEf0AKQ+N
y3p+sDN49yF1VFHmdmIV8eehpaAGX1BQXYZemNwnyJoyjZ/G51bHFrejkJjL3WTB
ZA6yDfwK9a1Qvxr6lltqvvmLBWIBMyKrMuZEnTBUMMo86O2ZDBnpsyE8sddfCPtn
3eze4aBDNf45E5xSgNMRu2uLjNLRLe21zGooF08jjBH5NkE6N4aAbOiWqvpNIv0U
lhpS47S3yFxPkH4CFNjvPzp+arWu/PETWdk46gzxiAO+TwB86nKB7KwgtHE35K4y
rP+Tp+gHa2ddXWx4DJMPxFIXRkBl/71N2Zgoy/beZUBbGmiegqo1Bm0zGZ83pIGz
x5WjtjypRKdOOMEbD6vKxbJykk1PYLnzvreRrI6fHNEd7Vxz+PXqhqyw1E7ruo+P
gfLahQPB8wTnU9o7FKZ630+cqBYoe9l08VccA7YL+P0LeYoDARUcDeB7L0qk9xyp
ua1DMBUX7HWS5p/NzzaNpg2U0eWzAkhLxTssSINKf0VpyuWyl5+CFO+AOjoxKYXA
ngeVy5230CnLIIFSQhupK/acoaw8BWwuw4DYBxuMrylQpEeJ7TpbzUQMBSQ2ALep
rVYTnOAVHonkgXL/ZfybpWI/8HbncUFczf3FS9omXjfnzV/D5h0B04SyBGPIgeWT
hU1LiXcRikHeDjfbi76ZgSFtVbv0ejTVEAlaIXHaUINSCuwdIoDwq73HhgQ0Uy4B
fiqjHcY4krade5xxG8aCnlya1b8mPziF+Zab1loahQR8i+qf+Ik7d2GmWXg3zTMI
wNXlsC5o8mp7Zdu6V6eYfAeH6vou7i7bZA922CovTTjbLKb9t0rKTTQAfrdfyKRy
CCJUA5Zo7s5lxNu4+KdRNr+Up8FJtWuAk0BbsHqsHMBY+RdA0/yMptg/VMrsZZ7e
Zo0vl+hJdFQWIyYfFs+snKMnVUTmAvhEkTY7RQjCmYctpx90nYmo1/TaLRcAHzKL
0kPrTiPzBzfqxolmaXqCMIzpbgQXR3poRxNBEsHtDH1cKAkr+ox1yuRLE29Or/Gs
/Np5vZgo6N5to9MpREEZjkaDcUm849cIO40fXz7BNp2wZjy7e8OYqdFCqk6nr5xl
UVADQ1IJVFb+Jy4wHlE12ccutbZq7R8USOl8jVlPVKChGxCEMn7uN2ifzvZJGaJr
y7+TNGNZTZF36bMvwLjdJo/csyBytGqt/8wBW8nQsPUFtPW+GgDqIIZyHKCwgkn0
s7auBCjfV9yylBJTw7eq3uydAYO9RiEr1Hcbg19++znnUPIPlUu6uM2984fySaBH
4jY+O+pZFdTazPM+w5NQtkyj/DVKyjIkeBthWFPB5DR3pr/KJ8ScF9vArBNJpIqx
pN9xTiNQMYibJ/3B8R8D5IPJ672V/aaKkpfasInMzdi9fqu3MOOtMNEAG9Jk5s6/
eTOMRQJ+YjfU0e4pwVMAZg65xTnmGDyLR9Dd1oXFItVeXBQtwLbREW0aL45OhdTO
eHnCDTr4DYXTBL6pL1aCsoUMJMv96Ou4ia9UtsOoX1cLVoU/8SptrXj+97AXR6Ck
NWdsHKoD1mzN9bd4XD2142QjMmVTAZEAMu4ki3hF3VdV+oJjEsKkOQMwJVUt4aFZ
GFlAm/C9QTC4mMNOlwXEBrN3zJfb9Boa6EPixMluLRNBEQhhah+UiP8ebognaS0j
4e45wa8LCbtSMc0dulnP97UhifxbouI74uMt/9QhXke/hjAbt+ZVCQXoAmpkPBvi
8Xin3FP4SjKxy/9LahmzjWPZM4oMh68Rq/muPXg1Hy4o7sekQv1llRSk0eHoC8q9
WieiUdUxxZ/QcgUIAzLVwboGySZlDzdmlMVMEfV0ck5pZwJmYIFK4GMmaXCsd+Wj
M3RKD6zeoXKm4XwuOsKM0lP0jSnswef57w8g0M06vJNW5Bf9J+Y1FRCrpD6kVBI5
gwWqQzXzXpqyzaopRhgBXNH+M2JSXoS6HxvfussSvJpx1oRCKm+8w6r3puaZtWQ4
Z0MQ5BG1s2BpR+5eTnYL0C5fm1tQ7OYEcMSL7DQaX9p8iUQFeYdJ3+MTibHb4j9o
5xKbDr/lb0eY/li6zwc5pXVKfCGYbkiwb5AxK0Sn2CaKjWPn9l/4A7Vjx0CrxyuD
NMAUU9h68GbktkS6177cQP+dZVERZMhLE6s99gCDlY7wc4E8MmnnE3PACRKqWz4I
jv+HJfnykKUZNxRU41wo6f+BRwTANL5JhdHIVPTQ5m61BnC8sUNywvXqFvG9KPqQ
p3oKYctgQEKI/NRNrm3qHFeGcAogtTQ7anYtptG9JmEcfwjbQ0GcU1rpqC343/9c
cD+f68H71WaWZpcZ3JgGdAwRNVMgqGu3J+sT21p+zWyF5Gp0jDcxsbYzNKjulMnP
khashdNzcHO/hoXWIlHXcQ7uqSBKZwB/mTpnhR07I3VGaWph5fZm1r7tUiNOXdAx
Z/lIDIOITuj3MXcBXLCgmCwS9T3hVN55MnLVrAhhvxc8Ma1Ellp52effA7zOK8ll
2FR1wLF/Zz8oHx/LDJfSbRVCPTgtP3bhudgqxQFDvq5Qwp3JtS62LlEC11qZYxtb
zlr59DSZctSL5hkaEQZOhm88/5Qa/Nlfd1pv12jqfM4zJfyFAmAdi5S1/QwzWUTB
bX3+Z3e5wLFkzlTLFGjAENOPL4jkoPTQaeppBJJPr79BCc62GGZIk7OYh6XZ3yGK
IbRaua6NsB6T3mx2JR9Mb/f8qxBYe9gvwVsu0uqX5InOWytle4D9ZkjAvWUSZi2R
AT0ewIHunLD1vj+Uhep4TnsubVXe+LOrBPBoolJp0ijJF9pQoNVmKY4JBfO7//XD
cNvYgGqGklCs0oUG6tPvahwx9evtLNwB+92tAqUp5BULRaRLZDUUeioKO37RjS19
eYrG0nasA/CDLtDJnlTu+/0nTVRmION1Pot+AF1kApQKfpQS5zSWbGbvx9lk627B
vfLTe8ku3v7AJ3HS8j2J8kwrbkjgUlEdQbwuk1TLG5vkw1CyFoUmJltsBGjet6JE
sSJQIse2e4ZaKiL0umAYk8b6fPLkaGo+AfXcbQ6qWsPQFJ2csJx92yb/0urMKj0l
uZh2TZa07d71abCFLUEjaLMzDSGO6GDofcjZQcqECmGRNX0/YV+vh8wvRiKTDJHt
lrHZyirI0yt3bQxDDIu8bPT5CwLmYfcVjV40zaiHVdD8i7gU4q9bR3rD7VnSuPIT
KG0/z3SbWwcLEqPIdMEggw6bMGciUhZ9TqKMINLlYgqeKYb/FHw8yocRbO2ggJpv
DNQPOOez9KNt07GjwmMykp0sAeEZOuT5vBaxuhrrkW9nkdyevp3S91xK7jVuv3bv
em+0qfz4MGpV0gU4LL2B6DAblcb9iHJ+iQQorQa0HF0Gx75JXTolu0w8slMp18pF
rZmx40r04QYh/lPjOl5fqznTlXdF4iH1GpO2P9thHnfpWnmRiathIFmrCF6nEFi4
xpLg1pIYXhoCxeRE1e4h+s9izcnxnPkpmkrcwVDwXaYx40OI6MHJtz6Dz2ZHEMP0
eXJA6P2P69oQ7/S0I0LQPc2kHQ3ii8cY1fqy//1Q+2Vp5Fg+oTJFXNdEv6B1iID3
m4c5Vyz4ycUZwSF+f9O8ZyfLE1f7o75jAQE8O44v2DeMopaUTh0IRYXgaM2V+e9P
/3AwfiY2K4v5NO+NmpexmNktbSfo1TsQQu4Jfo/UYK0sHTW4eJaUzpu7Dll6Yu26
bA+6fW0NF00londfX2Da6/fFGgcT6rWeDhdy6rWwBTCw5RJAeIew2eMCmxv8jXah
ecN7ommYRoR433pmFN91i1zlPahoPZr5iaFxb7G0D1eAVTdiNuuZEQ7FJxLc1EWj
05lA+7RUhiJPxs4RcuFp1IExsBJrW+RdGDCcxXvecqecvYBBu7DCeOAz5hWlALHB
bRhXIwlRQCfKocLxiqjucW5uZZ+LrXbfpVe7oNZyo6LU/BQ5ZJ+QUoeTlxhctqNu
JZfq7ewuMmQF2gujA/YmJaZmnYOTM3MwgZpLL0sMAaZvWu5oe1pocKW7VhBbkNiX
ffsqlZW827nsSy3CJ7o9JIjsYSPh5L+fVR1bQunWsxSk+YpCYJBumHftlhZywXl6
CaiTwPsXpiFkINPti7MiAOo166sOhTeGy4WZfU4Sk5gBegzIE05xn90bYyMhaNNt
25PhoHj+t+ytLzIsri6njVZV/O4jZtXkVCIH/KXocF3F2gpIgUcbEdXSyrvxTVHV
Xfy4ZuA47XWNJZ2M7xsUPvOf7BnS9EhoIpAe48ece7wlny4/nZYbI9OzGXea95Zp
YdTwJ7+W7yXZ2ArtdVQz8MBppssmuDlKcDb99FR7eQ0tVbCQ3dW6gMh4ZuryHgz2
Wu1jIlQYqmwjOt9CAolBtUR58sb3kktHp5jBb91sZ+fM2tAWOfF2vwKW2qiLQAlS
qCXHLW77LQZolme8yztkfH2OpE8vTEQHVmm2/CcwATEpd2ntrQyggF76Y9RROxTK
lbkSCr2XjNQfzLFb36p6gITb52L1ezn68nGYJAwbuCOdJkDMefH6yGoHGu6ddt6F
66s1yKEpgADz+G1xOjnT1n294vcFw5FMjQ5QwETvuH4aEtbPrPoDYiSTzgToUzop
XsCG+Dj02KEUOn0bSk35uN7aXS2FR/uBG18FArKyygnz3/eL+bR7qmaD0uOzpHFh
PcPqUC1tlQDr5pieKbbSR2RKdlkJm8cRN94lub671bM5RCOHlVKnW9OeCIWj5pS2
v7DuDWQz89wzFUor9Ut2diNUamIIFcv6ynrItafuvL6NpIDgirw0A+7q8DFu+VXu
eFzG69hKUWg85YCGvXX1sQ3tYCkm4mM0E85odXYGeHrBG40DNFak6/m9rCxG3g9z
nx+0NTd3UuWmS74XvWzY/lcJY7+G7iPEsJajLIorhgKX1IckRh9gPmUjNCSoZUse
pR50k2qOtnnypNDOSIZ22j14kuRaoV/qdsRR7/WyQN1Hw0oGACT/W57iQAfd47gd
bVTXe8iQKCVfIa2AMo7ugYmnpb1/rV3ti/fws6m2Sndi/7SLnXZbOhT5JmF5SGjf
JBsGR/VIyKnS2BAIUXlycV0sUAQL4UjtrHMj/z/22GqM2zY8Ho78czTueilNgPX4
SgeXQVgCJpp5AFvgZ7EL8ycKG5qP7QQ6saa3YL5qi7rQms7Di+RFXfrlfxTUBVej
aR2ScTP+grgo7bRobBQ5mk6DFMsRzv6N+Dd8MSJBqYrCou7h5o9VtvEddOLXxFBc
5NnAYy+N9NQTjnpNvcvQHvSkwNGWOYMeLqDcak78NIv3LBATtmwsxdAGTRWEfwc6
4GKjhLMvX+tTPc+djv6VrqxiZInt6rF4rpYJQIOHxiPxbuUiva99XYFeQl5AQR/Q
Eg0V8MM7Bc4iQJ0tPM7dhfmvobhF+fMZ5ZhYOSPwcJNxWfnRmhsyEz1hVHCefqvA
QOSJh+8t0uIPGpQrICWmc8dqZT7yhjOJT8/lz6LUR5f5qZJXdsqaQw//zSz/gljE
nX+Jf/n4SLJ8Ico8c6ecQch0E5FdyYIP26re2XVhfiwLkXVJEw3ph1HQ5ytACTVC
6AoC7HNnfzCj3xcw83kpr8kuxTAxOf3xktk9TTKAow9r+kQeibszhJceeB7b35di
84OgChJA1lx1d6XVrEZt7xON0RgnzrnX4EogP4zru2QtQZRa/K9s2lxVNAMj3d7E
bfK5ry+ERq6pIi4fzSCd23JQHjDgITkyN0gC5GoYvYX+Qa2bNC/gzsnlaBp67KSb
Hwo6rp5aekMNXhxf4tcmn6/MTtUXbdX+oC1Hz7VcLQ1nBRSNF+Kz5PnxfPFTn0yw
wi0IeVnCFDunzKK4c8vBTS9reINUYI8OFgC4PC8rq3shNrlgTl7ouEpUqu76zzsk
FF89Q4leh4xA3Z3ZmA3Es0RngRZ6Sx0n3nClBsFONN5FZzSnd25yisWUyis3qzNn
D70jVUvXnEwMdhzGugmB+7Tq9StjwGmpXJRr4QJUOIvAFbNVwVohIyEflSXwka8l
BsZnTktcOT8ynAZBcRKOBgXLyBN5wv2wXRaB0n/1M1vH35aLlzcBS2UjQz6OOhF3
aB2wWh5xM+muibHADD2c0McPVp6e77+0wvQ4fjsPSdbpkhL3cQheScZO5vYYHiez
yprbx2HZ4qgcBx7kKXcBNHMV4vFwhx+9b5coAczj66qPNktpXUPvKSVoVyVN5RAR
aZzbTk+Egp7dRD8OqAJofdh5R//wU1HXgrvSCepgKBebU3UV5WLHzDcvSFmltisQ
ZqgGqjLDpmtbz4Ifv2do3QqdF/l/mwD5i2+nnAxWUEYhsUIUEw9OH0/UUGQjBXX0
BHAT2hhDNuBvinIPeAHL4C1I3L5XXrS4KY9lyH034hjH9E6kaw2n+37zuQwAjGLn
/TKOuSesZgJ/9iZGqdOPS5owmOT0ZsENTpfYM6u4ly/6Q3C9kOzUSn5/8t28UpN0
a45x9p9leduCKJ1OX95CCj7H/gHSvdJRQSPQboJuH7mUEMFPFby0yrFFOLKHQPKG
bcIH0pqWRi28yo0QGjatEFMW617gCMsmaeaiNUGZYh2jFcNKA4A1VjAaxGFcprY+
Tt6GNnFgJ8korGvENS7QNvhSvHHYf54R5QVRwhmbgNrs5u+P6cxnIP2Gy6h5dT5W
v0Cfvc2vUN5oQ9qGT4q6kbmsfhyXrDyFhZWFqRBBYRUYN+sr08VCfEarlKCeAg8v
EYehCUSr84rcmuDERBPRjFfSYaHnOTzolS4oIEPWa5K43lPdKfDr/FucwtODC1GQ
E9aqDeLtUV+MiurBUMnSqoDLe3WGTKcGTQ9bvuelq1GOvFzvzpRnT2mwEYr9DT3l
HCtx35XOho/YQgZuafdyYKTeTjDHwvYykGoX6bRLnz9k9szDzRB3nNPogL34M+fB
Dz06C2FCDwpbZJIsgbMqvda14l2MHjFM2rs2k33iPk8W6r1zAuPgLdEWzQAWqbvz
znUZVnQLf8M2n44z6m8/Wu6J/lKk3JyRBdPHCRAWRH+XcFpAprUaaIklGUzsGyQW
5NvDfKFH0Yww7qSyK6jsUO7Oqed6QLs5w6J12BvglINZkRys0O5SvqfhP9ME+XZY
FMm4oTxFC3n1HPakfhmHTgAdBcWXyNDjggjKTW2M+SdnZeeIPde4Yfgrt8B8LOf+
SLecKEg37GRPZ95d/Op6USNNWOhLogOIfJUT/Ak6Gv14eM/H21QTG8ZJX/NDNq5Q
p+j62dk/Hx5TQI0oyN3+UYZ8Pv42uL/fAdXBWQsJwJ5y8QgZEPtk1P61g2yLWnE/
C9o+1NOCZ0Wg5V5ifmQlWb6rrhkir78a6j3dMDqy2UBjBAdLq7qhxh+QqiLNG+3j
wn08AAPBWBzE7mRevcR0YqOucL/dmfvulNOMfPIY3Atgkq+zSYsD7QMbQ+vyjh9c
xarubcimvXyxvMKJ0IVscQlnFpKIlsUoG/pTVL6yFOWycxRCQ9mqWek/0/xKyBc1
HAK5E0X8zEpwXK/Q4Ox4JQh05dRKQZIwomOWdHPO23aB+88A+iKLj1s+2g1TmJt8
UcQTaypUDRRjD3gGh/PW0BrO6hJ21bskVAiN4vM1mcJS1dsMQ7MvkxMdVUMefnwd
VU0fIeur+gnQelYjJEdwInqcLA5TdZN/+1q794iB47wOTF8lMyMp5PeIDkCGUofS
5hV2ZHDj7+KFRePI9HSnpZ2P9HXvu0HjFLGFk5nz77JDWbMA+gHY2zel51Y0P334
3/jAVNeJJ2SBZwA0+kSnoNM3u5AUSdv+KReA4wHOml+HGVR5fBHAxqkRwFdzKdQZ
OAZx/NhCfa9n+aS9AI47xn4R6DpjVPRPTQCKrCCFb7HbpqSbe4dHNgEt4xDF2lPd
CVZD/DzNh3RLRGJz/1tKcCkPwWxEOpBGT9eDrUDjX/N04VWi3MwmyF4elzxu/sM8
/UbSZDgnXUmzkgvN0SeWpKICf9GaWhVbM2iOzQUu2EjAVigVJM/yNfwvEJmr9UoB
u8oUdMxlApplUGC6d1qgJFL90chbj+AD5o4jkD2G0QT3FplexJkpHUlcrtOyHIuN
i4JssuxMNJP7gioFIdndvC3cO059qPS4XcQ6JT9lZ/fixBg9wwnEk9NG5qHT4Vvf
m7rI3nrJA32VAjMAYoDbikRoAsb+whZvGqFoY9VALTUfoMW87zfcBvyllA2jVOXE
T8HMkBtCQDoRRmrfBWV6yc5Y42njb8cl+jcxiGT3CXL41NOC9LlYhSIKWR1pfpqP
kozmc5LzON9fGVPubVa6dcqa+dx9IETiCDiIhZiEblWDEihQl/T6cdadwS6Qbd8U
Vb/1SATU6lGnXS2KO7xJ6P0bhfA0Bl2sIxTozybCIMFJYpmdCLrGEINUV0CoV/9H
uUi+X9yD9YhuTTkiK8M/qDYF8CEk0QDh3in9Ze0QrzQNmc3uGZa+K1RCp1/Dxc/T
CHCA5YKBwiKGAIn44nlALYQSVDIH50Bhmc/ONVBJFUYGTm3jEQHDkFETYm/InXhA
Gn5q1kE3093c6Xu5lQUwV83bvmDBikZFk4yXIv9J+Ur2Ooq2izyxfi9Q4RMJ5L4X
lTspJ0P5wK4WUcEnNrVcABS/uYTS+B4pe+8u4dLU88HbsnRqD2DghsJfwWW0H563
ssHC4DZ5a3DfJr7bo54dehIff7uIVw2gVPGCCWAleRGuJrUOBsRLrNAQHM3v0qgX
LU/iJpLoxSU1AwLqmRzXzVZi0Fhj78sAbksV9qJuf9jSzn4wAl3mU7Nnhwb9bYN1
HyA13SjYXH3H1L0SpeAJ/m1s1l67DX2ba5Kh/8H/yp604iXDY+d2BF7oDDWewWgu
n3BoMLiHiGhNJGNdNXV1EcX2GNdy4+72CgUz8YgcklUc5ESC0bsXfRp16RPjx9pL
kjaOiu201lTBnfMayk28pioqFffkmxaO6WoIFpm16DasgRp5EaADQE6z7XlfBYOI
BId/flbK2rCTEdVW2pY3jzFlYpm1A8aw6ap99LNiH1ROuGqzyzGn9akRcmgwyQTZ
fBS3yjqthTew0q4Ig/bSPX0RI81jAHmxR7UD2C17+ptVpdXd64zWZfg8nPZIE7SJ
Lj0iu3MqSbDFlsbRTrLuz4EZWYf7zTMLz1k3vbg2JJUgDSFBiNEHVP+xqf42xAUo
kVYIoNIIrhAcnIY9FBC92f9pIdpOfzPBN0TTz6W+19nGI7gF+1uuRGzjbr5fVEqh
MRqagxY7QwbcNJa6bpnIvSP1xz1ukLL/9/kWtABDEgKiXtgT/HRaeVmG2Wy9CrDZ
SD7g53mN06aTugnSoaqAdvEGLJNH3ck2BVL0IdtNPln4AC+d4N/Pg19WfVhT/fds
gEPl+YowvFA8a+tMbh4VHig80VneoDNml5Va1zsk1CEr1yc7axrjlpUKZBSrddM+
3zVLP9+2v4FABk+RGX7gRolE+jTM53BfutLK6GPrOPUt4vCmnfTPJP09l6JrSRYU
6j9yJRj2sz+Wh3uNuArCNMMHY97qo8dC4O+L2+ndTPF1vyhouU+8WHPeE7RPDEa+
bG6hUSk6O2hHp0v8BxHeSZqcilMCs3n0enTNae3tGpfQ0lHigh3YWouo+rMrRdYJ
YNgTGiuTaJqD8uIlfXPbQo29Ozh7c6KEuEIS4Lvizl0EHlOKEk64yw9UZKb1qyCV
9s5u0US+N0AioKD6jMpqNTKT2CqEDuRZzQar9xz1a5FjZ6y4PAtHyVqAfT5Mpk9P
Qnzf1pb+8lhbQztPPM9Lu3xVfdwjDZOOkzl+5k8SbQlMbG8OnRJQbom+FZZ3m7+L
x5kbYOHKBykFZEfB6sixiFIlmF9r52se83eMk7yN0R6sGvgbu+dnd9sGBeETyQ7d
tDhdPRJ1ToBJhelEIvTP2OrYl3N9nkPOn4ieJw53IDNH7WE/oUVJMBYZVtey9bSI
aPf2LJh8K6BPhctRKfXuk2j/hkcv+dy4DdOv/hPYjcUXQMZLJMhv9AL6RIViNXu0
YhNbwSaL8FKY+gng6EuZcRgXHtmL2a5Sk6PBkXQkThEuKWnOop7gHU6E5K30IWnp
krtuh+m+t1No8H8olDbYvmaLJmKoQRks+Qt+Tsj9uoqLBeogakp/9AEd7f1cpnji
fhz0JFZ7xnEZP51PeNzxNM/Ecsad7MNb+0GqkwZt0hC/1ov1kNLWgIjT4yg+mggY
cz80+Z/dl9zcZG81OphgutUfEWFS7sIFo7y2wmTInvLZ+BvVXk0WMvQqAoHTzR3H
0jwXfJL/SusIt0vFWB3+0E6crMHzOKT/7YAMHutuTNPVZPUt4tmxc1L6RNsOpMIr
aPC3CB3KeGSR4SaLB+G4TWSyJbrEMYv0gi2XpEuIlJaoQrNmRZr7qOi//GkHCN+M
aBMdkJJngq5VeIjMQKiBydYD0clT3GMbhoBSqUzz42+1SVSrqWDGH9O/1duoYxSa
JP/z9yKW832VDmkQ9kohv+KQJOGesKGN9C8msGzRAJcmahDTTsHcGC4kNGaxNx5y
on0Tt/V2fY6X9aPmU+TSsalmUxg3AsKiOCZCKEqRvVPAsnMG/vPpD9ZYz1Y9uuws
Qgbh2Zp/zxBFI95Reo0FXc+JVgXHkEzwXgUeroF00eArSoQ3d3Efoo2KEGIYj/HH
YJxH5ajmoWfjXpHG34QNz2P9n+/sX8+GOttvGu0+PYRQR09AE5yQNFsVzth11XZE
ikE8Kaahh8Ftj4cfgvyXiOwFWksglBCEHzGW45ex1s2hJImsjmhFQY9PPTfvyn4C
szKCQYCX1N1iGoO62hBCwY0pmHR6EbsJ60Mq/sGMjT6Pi7TeNRqMCpjgKMfORcN5
r0ukwQNjXoVhY6D64FLyuwKiOOsABJ2naAB+4QNy2KlCqLF1Cb4xmwGSZ1UIJy38
sbv/2zSRKnoIiBJbsLTEaHskHnuzdEC0zH7/Z/JaqbOJK4u9G59BEO1EvwmBEiBR
9blqtkJa5WK3zjkfBP1OJaBKk+U/vBFObPXmVQ4cmeG/VAXzRKoDtrOsNfVGyqvu
YU7WV4Wo1YMp18B5ZlmCS9n5F0ojkYDCXX9Gra52bi5cmvDDufs94aueaesAj+19
fCJ07zAV6b9fn83RGgnBaF/Hs6MNixMFmZ/TlAjcWj1g0ETyQWqAWKNHjVfwh2FO
WtvdD3RYovdQhJxg2JwDxphj+fFXrlVrurxE4C4Voll7qE76qnf/1fFxDYDVNQbf
/KUZBG20+9ZeTR0jSCAklYIsOfIGwlpAbSJ6FhNI4BaEO1VfT8i7PxYpTC+SYTXP
EaVeAN/rFtBOs04n2MwFbx+wFi6N4RMjtsrMgUJpLNAF/iOtpqEqTlYKQXw8QIXq
sKVqLxpsnyYqBIkotrNp5ulIpPtjDV5unVwRhiNGZ03Btq5SkFKkFCnj+OirPMLm
z2hHrGvrqMIsBl572Q/VRvKVZxsNfqO8xzFj7e1kIqpul3Qb/rnXA5F2sst3qVEu
xrvJ5oqyFiTlKY5VxYUJUb3rcn8zW2tz7X5uYaLnZuEJuXuXj2LwXfT4poiepjrD
f7ULqZBwtUJV66KNASlU359yoxTP2dKGv1Pl311ySur+m4E4mdreDYQBeZrWM/6p
kn8WUeoigKG6VRBAaAqTZ9Mjn/lBDWsuRgxbiguvZjZdQ+FJaIQwtozGR6X+/YX6
ylups+uEZZs5R49YrsRIMihUPonXEni6J8cnujexJgEzhgN24PkfqVl5l0z1BJ/c
QA7LM7LIT9f0yiYK8wjWqb500ALpYESIuICDCob6P9JvJOkgjTzz+otrIt5eAi6X
Ag8edRPrHuXdGmM/9mFeTDWJwFb/CoV5PHhNeKHRgjofgPSG6C2eqwY2bzJ8KCA0
fm5wbXwO3izgrI1dOnVegXpPcrFIk8I3AdKaRgyEGCeKBQcuxtpfcZ2+EEHT2cRg
yGUKpMVB4pgo5eKmAlEIGhUcKgJ4et2Clb3XnpPFy6UkL7C9P9DQXo+7mwGhL5+U
8veKqFS5yQdH6Cs6S8CLqZqbDFjvQhaAiMtPPhQlvqQNN5gCNSy7b6wyhae7GnPM
pYjL/QAwGAM+1pB7u5M6yTZCz1RS6HndmWwZdicAB2NXF8tFYlD42ayoVBrwG6Fs
2JzJv2tngs7N9pmzWHnb7BceNF2c4/pJkkfSyycTSEyHi9uL3zqXdh4Q2msvjdeS
1Jc/ozz9FXugeRB/F4QsUHukmW2Sm1ut2teeD4h/w7tvLwGaZspMWS/DExTrkQMo
lIpSX7gJn5mcUSXROZwV6+ZkW7rcZ+XhbZkU0BwkWBzR+orzpKmfSw704v86Cd0J
AVQII14OgWidK6fvi3ewCCP0TvIbkPyBOYWA7f+yFOUA+4mRvCIi3mK18OKFQ9VC
QhsE3WJplY9E0FrN2rRMwr6vNL7e44oOdHSjkOYK5d3qrbwTSbhv0MwcgMkR2t5c
anopdzQChgsOkjNU8RM0oZAowZp7b4PoBkgy8yf+dIH2tACKwE1HfkFe2aIACxG4
LM8zs/6O6aAiPTElQEKkPSUJPoJ8SV5PzSo2D4MRSxJS4tkh6QveTyFYIXBklr4u
uAdhSg++Wv6ppaF/WGUDBkBWQJFO8BlfFfQcGJyQICqcAO5o7oF9f5iLQbpHP13W
RvH/VPnV1i58kWePw41t61W/dz97fUwXfAzqSbcBN+OEq65m+ZsZZGFdQXrocdla
ww0AJg++Bfp5C7gVFI77Qp+3+ktVwgQ1zgn/oegfGOEevrI0xaIxPpc0+l1astiH
BqIbwmZabVTL8Unw9gNbLfYNjpJqdaYEsiOsWBaFUPXTtxpzIXPuEXJ30Xd5MOhr
7yM6/nElINfuHRYeGjwT3bNvhxH8i/Zfz/IvsoPR1vrKQIFntPTgGYlQxj5Zf37q
t+XXKjKw9u8e9pDFyqODdCFINrMljzzYu2QBsowrl2B0jeORM+5xz/f28PCIN0tN
PJikt3IDszARh8zHC7n9eLOtZGiB4RzwlE2GEgb5KAKqs6n00OR+8kMZqtXPRWWz
7MYpR0qLPaz22l7jIc2O13fHrjWxPzsVpVgYtNiysCG7xpU+wLRs8lY75cvLR8ic
F7e8IP2uQCOajH8tCWX9sh8CiwPlewuWet7CZZqNlUFC6dWHR99DnZBahVQ5pXFT
JQBIXaqmvtJ35dMJUFfv6Fwp+AngYdUCfr8WSNwSF5K6HS9/d18hXZ4Q/FNMEFrm
wQpNgRT7kSwQvVTeEBLgyI1+QVwUd7ZBkDOrZGS9vTYeIMxZVuImXrlMPGfF4vP4
93vWdSNmGryAHYqlhccCwFO+6OOA70YWCvTwQlkIedynWVeD2aaZzpqBxrVyMDKq
1n8mqVtG02nf+InmXkzTezOV/F341y7x0JH6zpd0KveMfVFVqnZc33QJalpD2QcT
xYUQ71Afs91FY1BWXaH6XBaIMAErPBu3sNabeIcwJSzQSpEquauQSASXSI5VMaw8
NABBwawUr36+Dl3dY7wOE6aw6aP71xsZy/UjyR8SpTWC5chq02vhtHRO8FKa8SFt
EChU4EXNhraF6Og7qrmY7Nbcg0ubvlGvBQ9TWb0JFuRmZ5zIBbzBct7n1pOTDQR7
lJebiX8iIVvFVFsVJS9RhsMtywhKXPzfG8yddZGvlQID/yPM0sDZ6Qa7u6eIH4+u
bCjIKs5wOoh2eBy5neGceJxNSUy/BdYfhKHzjfRyzboBpn8ZDM/+YNJXcy3dkGts
ksAR5SMJsPzkqqookZWXn/dIKaF+fzXr2HpyvT6O048jUfXmJo/v8wU/Hpu7dcAc
rr0rz9h8mdNXOudp2d+U8WXG+KZ2YVBy6txtCsMvAlpNB2We/Uy/Fzvh6uCNQHoZ
IA8RNEz2/A68gm/Ds8fgSFYwx7/JYI8bS0w5mIo+6n1bkWYJrxb/ldUfwf2Z6j69
VaUy4rojZ4ASFd5xIpQMndK06Ek5g5sn4br0eZFBEFanTRQtrNrbnXwzkRMc9nXZ
KzHkKOnSSnhZY2cy8hUFNF7h9WDaEm8IVt5azwBLsChx0dwf3p0pZAIrsuUckJkp
BufsaaqtKunRvaC6gl35mOAb8PyBrrKPTmEuVGshqPbbbVTDNsjt118VZrTk1iOj
1Fek3oNZkgMbea77y8++OrdAbttM0W9GEQaLJIRDoTTt03TFC8ffFpQo0XwW7PZA
065HFRGMNSXGQimnMM2NveaViqDfnz4uAH3bidBsLFEPdNMAH0075GwmcMtpgaft
7ozm72P6LFJVKpj5pRda6jXYA125QnVu+39Prf7vo1XXQtTd3dU+A45Vp3yJvLbS
krGkxcLnXriabxKsUQVKLlEFDVY/QddRUWJgGk5kRhsTlA2q9abfqeZjmhmjz2eP
Bf1T3+DizJyTbzTgBQTTPuAZkTCtkgBQHWEEYMhOBpSNrGrIajl4HZVehDbpC3o5
92zo9i5AmbsFq0NzXuj2KRhEfaolLFgOcDY3F3q1HhTfQ1b6D1C2JNSvzaz+rNEY
UVc8qSsuf1AX/36roq4ZnzOKZL/XKGyKzUc8fAnS4prKQaeAHeLZsW5kjli4U66f
ie7YZslM1KWmBYhnb4EZVAvG6g+rAOxPBns4bALHw4rfu+v+1/cRWFnOJfFO0r83
iz20pDCAJ96gUgcYMTAHmoh6vCeygDxrglo5ElJ5wiFzd73Wfuw+bbvGxKZiIq2O
CRiB1xFG6j5lV3dN3ij+CQ2TZ/HjR49MZWpEOTrycgeuCkTP1nTvbhhfoKPAHRZH
f+st2mbXjOAt1zqTUKSQIefwEbFTz3AOhNrow1YMGZ1Dm+HpLlB7ERNlufTWNi64
FweRaoY8BvMgCUgjC0fd7ey8MQkCQnPHgfhDOj8dhEsKS+iGTnWz7R3hRTQK7G64
qHOoc+k4kuA5YXcDZZN/HeAl+wqVMb7ujuo2RTQsbu8H5jLYH1emo2c52a+B9l4w
dF6CU7ZHmz3ZQShZvHxn6meD8j/jCOp6SRGEWoHhcuu0y1+xkXdAtBpzty1lcqsS
yL8xPr7AINA6ZJkYQZsxLQj6nSiO/JeviFDMIG5Q68DSkjYqQnYZVGN/OI7UDpOJ
RMaAr2aUhmfbZyQaZLvSsTSzM4NnHI5jApO3meMqmZ1JZEpjgFwZ9CkJdyRweGCT
T4W98eV3yFBlZVhCEhtLj7iOA33ABl5n/NS10a3xE2Hczq1NjPMXN3qq9K/hJ2QK
usjPiSP7fNloB5cSKjOuPke6jmgEmIkbVlgUNez58mFfiv/03Nd8mFBc2ZySRMbe
C6n8mpKIiVcgC4VU9mBcfUk2Y9liJCDNizmN6kC0kMbnoXlLJrUIuZT6hf6rCn8t
oiq7GloKYb8SbN0xcrOsDM8FCAHadOGrmdMIFlukaWkaAJ8FN5aXTI0hq2R+aoLa
W3/TblxogLt4UQ5w5YZ0g7rz+YLvD8bvwUkAgy86/U4sKxBSD5/QxfQsmCatBXDd
JbwmsFAlf0VXYfKl0bXS3xYXnIVCqiT75cBVEKRNlfbIZeGFW6TLjWJFTLGIklzb
QmsePtdnuU01YdSMDfUZv0EXTrYZ/DtE/CcfqT6MwrOHAGMJcJWSRaww238SY3S8
YJXM9pn4KE/2Vu1VC9TCj8enqYNX+fymSyVxQi0a2D0O3WTDRRnQ1ZzoqvHzemMi
7pjxaz7Tn0kWDV1+ahf0crD+5RuLz7V7+n0cq36Gcm+cxTwukNZrut8r90zLmsP6
M6eIwCC0slvbtWh5Ay5YLg3SokO1ojxxJRoVHW4+PcGCmPt7uo+bNjIu4c7/wjDY
IS31YR2lay5wc94zbCVcZU7G6CBQtROgm/HuWEqIDC0jL5mKavk7NTgHhcPQmE3d
01pVzaeuJijVAc2hVXgSfGKh/2Kp2o3BkvHd3stjYIr7D7gzzxjAZKDcr9zq+os1
wp0BhFVLU9bunsIWuq1ihyF9vbMy93l4zgLLIMzEUqUrXsq0Nj7RAOLvyY6nfIa/
vakztPf+L42ZLcHGqZXLE1BCxfiufLe74d7N+DiQC5vGzowgJ+sAFA98ocxoLjLI
IjYsjB9X34ZGDQZF1DR0YZjajBvXy6HyNpPuyJ094uFhMv+KWqTDe60e7nBj/MrR
vIUKMyCJpk21pXPp+heMIr4kltuKuEJnr873WNsTmT7D/Ms9hckzWGW2JqsIk0hl
u13sMmwcVAyGCBX5W3TjhwX76siREOrLPqyFHsMUeYHC2gIHl/2cLeocz7JA5pTF
8miKY+DHcWU/vEQbYZZEluGm/aD3SZNIJ6zvna0tADn7yCFNvEf+AUXIvxUMRUt+
t3zbfM5faibaKkCkaBmUQ5fvyCPbwpWQoj0IiIF7fNjP03SJBldnZ/im7YNey1to
hs9mZ/o6h9suwJC4ghzYhsFWc4bPPtWfkg7CP95/zz9HYKkoF7FJMKfRXdDsfTpI
sl05fkyAt9GRGNY5wh3G83ewtt/mlRh2HepqmQr1t/Kc+OeVVlaW94Q7XlFt3o7o
mfJl5tO6qvIEd0hQ/SXSJRbONksxD6a/kMBDyY/AjB19Mb4sZZhoZZLZyC7UUyuL
sOswy5Wu0jV3wNTVrt+RXu9JNrFq7VWItpkABSWLUX25tk5y23Jt9i3ZA7KmiGdA
dKXk2iQlU2Adr4ulgzOxFVdzUa06kwkbIla+WK4ANDpLxhESyfTMrpIAyRw2ftMH
9PglFcc6Dp/Wy+K7G944fBVM5TPklRuhwVHlbva21liAf3ucBEeVenKbcUZNqn3p
tqjKPP+KPp4SZD5e4jXmM1n7xGdMAluw49hTISM5dkusaAMbGN9pXpxr6dcPtjbx
jf3iWVayQeVeiu9RGZBlf5NoBGLqG5aU0EHgy6BkXYlA9qJFIToc6/vcVTkGUlKI
2TUnYub5HQ6n/2jw5/pSQEFvptbgdwHkIwL+6HvNZsw4ZAfVqjYZ/BSSZxA4Lix7
/U063HIWyVlStRIY0pvBP+beqEbVEWTxOZhldfTRwo3Or8alT8iuD1Y7lTt/IvSo
FrTBiObyWD81q73sewzLTrHpkgdVn+jp8KcN4z9o9Sa7OKuZsjhX8VofjcM59dnJ
m3o2red+u+egsDb22e07Ag3A9gmXyXo7LOhPpKmfYAMNOcEosXWepso40tEcD0VF
o00bL0FHFZetsSW9iQrWBIMXzsHS1ulFa7tGKNdrUd5vhwFqKh+gJer3BsWbO3eE
uztVGSMFnq7yHFMyZj89vxKl0pwQYYNMnIIlt0ykuJljxkFgFP0TI7VcDvhGwF1r
hjkCrWQ5UoDkdV+jU5N8sOa6F/zchGsXrW5nTyGTll4G3lLRxYoVGfpx1D+gQBZ5
2jCMrOyujOGFysWeeegXOivAOslIb8qoOknB9NohH50/SEwLbxzfbIlOe1RiDuuC
3ZrGvn/mAG9SJUNKNTwbZh9jelDFPxVBK8+L1l/VU71aFCptQAxPSxhLRWnEsccK
EZP8vhJ9FRJ4rtuCjf4UELOtl6/D5+Z7dgF/jkIeG5wBXCnDSEhh5WujTjuZNp+o
YQzjdm39PSXvoEtHHWK/jkkD/+43L0axlZ6QqrAocdsX07fHMrc4yyTCBG1O/UtJ
NydnlZhovYwzeckKUre+EcTsj7vZGKUzui4iMwCxglZ7ht/rf1KulMUr0dFgjxkZ
M6Ece+TIqRU0AuPyWKtvVnqZslnaEJByvVJCKHG7TPz81PzGTaeOb2hMaouToF7w
ZfE5624sxQiJASo+whdbhSL+QJaR0zRsIrMqYdRFnflKm3CiY/LwSfueTbZNhWF8
zUoIQX3zAA8SAhiBAQcwDuNCw4Ow2tbKxLhVs4/5QSa/1gif3dR0STlbUbLgdGjt
MB9EKnpoyJJxLYgRXqixuZL8H7ENPJoYA8BKLJCd2IPE0OelhCWnZMdSw2lWlph2
cAxZiRbTQb5R6EbK0a5hF58sSASazJ2dE0dvNJIbyAdSGKAHiIa4vOcY4ZQE+xsT
YWvbtbQQsviW8vV/ETdVipvzBdXho89OT8YdU9iEIuairO9+olrc6o6iiypXBvhf
u9jB1Ypq54e5aFb6E/UNgKlnUywXzx48RUNuhWkprwqmuKmFjcR142QrM9pDH94C
QnPVSgoj2RxNDDptEWEZzaadcN0H/GSyrnJsIau8Dy1s381j2mrLcreQyy7ilIDb
A4e+RfwG/92BhnX9EPhTjv7vH6Xmq9rQjntklsYtqXMpDgq2YOsQd6hVnIcj8acj
J4/hUvHuoKslXLcMGViHqlsymA189Adovyw4IZWtBR3lQpV2rrkgdi3LTZJdmMcu
LjS6tai7qrap3m5sg0lk/Dr7bEWGkJmjymdmOOKnfOx+Zi33gUtgASAljcYbkN9j
rCkIb4cYF4JWD4SsLDSYwg96Rq1XEZEmoprQqB2nNzgCorpbPtB3HtXlx4AnFaMp
Q5LnMqn4FCIzaIEZsn0m3YvYXyHpDx8ag3WrADnGl9xmUTFK8Myze/SmN2/yDVMM
f2ZJPReDX9cdCg3vBL/I2qFBU64ef3ajOm8fjK9GghaO+M6prj/zg+VvZFtZaK45
ypRWkdTKB3Vk2fmN9NfczRc0JMt95dI8oI8u2PgDZpG4Ligu4/fkU09IxqBJGvpH
Esys6eET3yydcXwNeCoGr9vYN63Rb1xXcoUvUXIHZWaeWaDAaHzUMk6AIgvF1YFb
irl6T9oY1SYrGF9Glo4MvDYCzJFWbZyPGnMnej6TVSk7dSBetUfOOGtfBJF7q+pp
eEt8vycy8pkxHH1rn6uL3jtfGNZgBWCUIh3t6wEpEuFwwmLi5DsfamhAzlkaYina
wX9PMvE15JydPvNZKymEjf8PhDi7OMzJ0SPuwBmTNMKXPN5xMuDPNfLlrdbPdTOL
RCNkQKUOTz4EN8553e8qwHKvsMp7GVJZu9YDLKUUjyTfddOFjBT1mX/7eWcUYvIg
uYaekCv8XSMMuey1BrnYxUy64ODi6vuPIsmTlXaQXq1SFvqMKYjRCopAr2XMe7jd
YhLMs6JGshi0PXlBhOlwLQOR/OJmLN/bxc+kmzwoIbGSEnVPgNUVbGUKmwfCRCoS
WWcxeOdhSGuuCMYKHLHVBdQo+Kj77HWC8IIsZt8VEoIDhHDxOUTyPn0wrSkhDYs/
uD57jijIgnU3Fq8FBomQWtsqs/IIavdGT5TMqJDTcc97hmZdE1KtSIPyiZkm5Sly
9QgxPUWgYUMiNWsUFV5Uyn30pFX7UjUAEOWZnaXjFryUfJ6WA4AR6efi0cQtL9PE
prgW9rO0U5zXmuP+LdBkvUmuOZ4aWVbIB3L2+PAp9O37oDCwuRAwDnHuyM8ESU0n
JMlwKKjkeByy9QHO090fb40qc6fIwzXWn3g3gfY7xUwdp7oSK9IbTTQiav7JG7jk
2Ci7/tShppUbS/85kfAAn5wsIzSqKnWlsYt1ww9jkrcmbQ8UkoPf2hurSTkuPtOG
eL4eg2XzSQ5Jd961iDseVn7vJpDM7hZ1pZWju7QoWZ0+255o6nn68u27HUY0yaqr
7LYXcmlPA2F+K7B9B/ISwkwNETbIoq5Tu1X4/e5EnV371ZRCY0LwugGVPqt4bXLk
Pqp6cNhD7pSOI6yDWBYE5m6j1t8lCPehsn4hlUk+imIPa8EFjsFDrb/9BpqLhbxg
UDPvPnYOtxemd7okwl4458/bOMnfiULzddxdtVgUg3asfSnHFLhE87SO4et5usVP
/HkhbMK/lnFU8BTvTqppKwufpDabEax1vank/qzkhDxa+/qFCmrelyUy2gJvFpmm
sUzXz7UNFwT9JdfA/vaCyaXImSzx1PM4upw3YdKCtQrpcHRX8tb1oxZc/wOo/DSV
FE1o2MGhEetVTZsyeksb9j+1PFID1afuo16BiWHqv8Kj3JwFvmCrtFnrPpyH5dKH
/Z86tMNe9F8uf8XCHlBfOQfANDenKlalDZAxfhiVk9fp5PQOch6+pf82L4rAWiG4
cnKDnh1tAbZpvBbO9evW4AAL+DJuUSb66HtAcWQdYgw47p7RZnRvdPWr0DlG3+54
TO0xbkmLZmRm6eyniBKF6mJPDHp2KBvhcMs3tkTOh32V/5r+eYMmN/ehnD0xUti4
QMDtezR+q56QJn/JjIjoELznwpJKvqFP5dAgjJzddtZGXRqzevUcNZBwVD8Yi8+3
MuxuHiU+V/BaL4cawIPs+XTHpalXWrxTEbTYhFW84KYuEM0RwKvxN6GnPM5fORA3
cmQJIvQi3NdwjBYysCtdnKI8aTZD1njImEvtn8NDgUf6eRlfpI7hLTH05VMJEFlE
9k1UecaRRUhQ01dcYIlB7V0qamM3DlnbBFRxycUrHgaWXb/eH0GrmQ5jq7xxoJqU
wNKUrqTvbeFPlJ2dt7gzzwPIpb65XiQQxFrNM+P8tVo8ujqe5Sdp/LVGeUwzPBeD
PvQKmm45qjZh/vl4sjyzGmrpfwnWQFJig4DSm23E78Bc6e1LJb0vz/u3XBIwFDpN
fuzbisrkeH1pJQYu99P/A+1qXGJy4k5hGXbbsK7wCFUn/JmuFzFYLDld2Sg5O6AD
vySLG6VlLRJFsWcO2lWidbX1DRNyDlncTFco0hrONPtgr9CxrzgjxjdnEew25S77
vREgZldT26Uo3QOpJIlk9FZF/+3w6LFi5RHN4JyvRzP6EegDcKKlX/AhIKRoKBUd
7xxScuisV5uJ2rkdahMp6+GIZ2Pdb5jg5EK8X4owXj/TxSjESbfWvrS6KpeBKcuz
uVTwtZIFDo73JQAYtwOsOQ1Te/6lWnfSudODNXtlLM+CXPDKtOz25cIOuWJlx5BV
YruCrQLa2Y9Uq9PJinbBPmo5T8fMyB+pATB6R/KEPKbFU9ZCp798TNI/GBn3/IQH
9uI8v+JkxwooL9aNNj8L4HBP2Ah6fGDXYe/E+chWFFBkvRpBM/SL9t8svpAeZMt8
kXLeg7jkEX3ipvVhhwNUqd8HoNNAT/Klwdh8pTJTFzyUbqxDU61R/zDu7B8WnAz4
HKsb8fwPnCvjBjY7MS1F8q/ig/TCFrB9LuIMXLfHW6QiqPyg7f3G1EqArIwOajsl
I4M9Tch53XoUQFz6Zts+20fRBYCTeGRRfFQugn+ObUK8Bwkj0hkFtzIAWbnv3/oa
0vaPR09gHnwtmf0Fs6jbB8OTDenXdauS3DdulNcyDH5KFendCSYK4xA5F/o9/OAK
O9MBVONt3dwWEDKRqmNcpDW545sTv/eQoh+fPZbTL0EdgVPGM7KMoXXIzeyLTrFN
dQndtDOv7y37ASkN3G2U9TPYVgNuB7ruG+D0iGxKaYbXkdqhuSdx2s1sBgyI5x5g
5LKqbPxIqAxSUQjs/JDdZQpFWXo+th6tVNTRVrmc2JRQt7eEbh7k1YHaKVo5JNeU
Fb1HjL4XxM25b2ysjI8nvbCMoPDYCoRI8ZetEL/0PTKe7q4W1amT0091YQFXJC4/
vuf0y39VNRzqgmSwg4SvzwyoH+NYs0CtVXguIbHYqzYhL3wy4JWobHPe4Bh7yA69
9fGJseap++P2a7qYb7LuoSGM1qj85kB6A0ik8KGMh3Mpn573hItqkEfWWF5YNKtn
uMdLk8cwWyWzNb8Bg6aUCYtawe2zLo+NYLG6+UMdzV246krY7RmxK7XFqP3ORza7
6xu8+O4+nVIG8H8kFhwK+RP4ScGkIii0M+WtHiARg52RkwXRyzA6G7y7hGwxwWHx
TKCYPcpOuOkHNHfSUNBmrmsZCHwKsh4uHYVubu+mfz1yoX78Owlpe3rg+q216/Xp
t7iQ0sHe1vdPPppSaQpBtVcSbxeYKbnmEAAp3KmE8pvXHozTPiy25VpbdX2tR46Y
bqdAexZag6xMP43HH1EZ1LL177yy3MXDyaoUbrJ6CLv2KAslSAJIKE7xFzOeO15H
E/Zp4vT6LQhiTrjUBxDvDYXudcUJItMx/b1xMS9fnat602HyRYuucfzuNBPMIZL6
Yl77Pje0iUoT0hESWMIsJHusoKD++BbPCVc8k7w1Dn6PlM/OwPNzJkoifHBV2FcB
e1jV6yg8C8zaq5JIg8UuSZzwg/29j5dbKsLK9/iYBamboIZhm9N3mQUKcBwfmu3F
/J/DwQprFOkdmjTg43s6RheMwBRQy7h0OvpLa4xKMYO2UqO3RsHv24NeWlx9GPEy
fYok0C+hQRPc7fT8xhL4DDV2cp5Rc1HJvGQfs5g0mqO+C1AoNL2pRdrgFutTfwft
Bf9yrqapwnTIGmNvoE02cZttieNv0bkQA7qyjtEf43M6bTrwevA2vq7/BJqGLG3q
UI/LqWH1e8zmGZorBTlaOkMUyFKC+peQ9siBp6RCly/67unCtLOQt3bQbmRotkTM
HeSUh/5LUJ0hXm+fQf4QiNq8nNkiJVFvQgMqAP3YQiDCTcwmefUjnnPf/lzhRlr0
5kpOCnDWC2OzeoAsc/tjhdSHjJqSoY0e6IXqXJX39sWsqect4HvveWhuJ1NxOJhj
DGSARgH//FO8nkq/UKTVPKe2y4Chz4V3RJzcSNfA3W90BHE7Gf0ZOgFAPq3z8pWH
+HTKaRfcPvuIf1fF5VUXAOW4vshHPvnz3rbANb+g38trrxd7u9ZKXwIVcc/nGegW
I1j2yu1CYMgmSGBXLus8fFZsWyVysAjlxRJ7r971EuGZhPtS0Co5KhouypOF3T2W
mQv8v49pHj3XjOZzRmBa0bWNSti71fPmVpnjuQ73g5hRJEJUYNC3UVR5vzSExwtY
lDbE96EAyA1Kc8UvzN8atEXcrXNnBhK/FVrGlGL3QijqZWJl4RfogqAdHf1PZYjY
mtRlcAnUrU64847nBxUUDJJl/T76SpWJ8zuxOT4D+bYLEkuO9qMiKOGbB5ndYGZx
2B7B7CnKWeuyValGkdUYRuK3E+1KlhDB5XIAckpqoOThcNBzp4kb2xbtMRCi/ipO
kZYIHjnis3xQYKRR30RFszhFfucBJi9pcuS0G50KgiVO77qm1XdBIVDy6z+0iR7g
SRs/wQrPz0ailAqt87mg/mg/rylCewXMDEm4ACyg6klkevAiAZqRBir1hQXfj41W
qX51wyFZNfvz7j7COK70NGcOY1yF7xMt3b/nc1taxMnkpnGfx+9/AbUJ4+XqU+l4
7rHmRQMbKxJJBHJTViOZUbLY9iOBXtITzl0AFCMSw0V9MQ7dRCmtR6Q2zo5fAiWa
bjoO8zCz+vbsl5Tb5npGYXjqHXzC4sAkaD3ivAqd0xCvgMSx5QOj6whWX7MIUMEx
obxcNV4nva102pVWJJJRLcVsWMHTMa4N6qBLV4FZVs4afJeSDAYm7I6xopn8mm+t
CC5FH9PmxXU3pYFxoMt1uQySDJeixxwzGPJ8crr+EWwUnD/roXInBOE+V0+MM1U+
Id5MIpiBZTk613IU7HzLcLTaXdFpGeMFEpTdC0Wq4WLxynqEoImPKbS4Gh0oTaql
y/H5EJKPu4PaR7HrHu8I1a90oM7HLpeNfQUDEsXZKe8kflsD3uYOXmAx6lIQcBBT
uP580nnSLYYEQJT7+dNc+TLppLNd8kUSey0SJI2ka0glvPlOc6I9PR0S3kidBkEs
OmBF4jF+ipCTBVAvltQzlx+jAayF0H5P2IUkBRx24d0OPrWIBmgKJubfeKVjlxFb
GvkAaHW8swcIBoJhODuv+S9bXPyLS+yUk2xth92ve8SXE/uZJ6/rH8GJDq88mM3B
HD/+Vp4GaUrW8SXcRB4Z2Le8TuVcqgZ5/Ya+i3VjGU3rMsWf1SY1tKihwy+0aNjK
8iKjpZoZusmaW2ADmhIURM2VsTPcusSfnF1PYNhqmau+yg0Ho6eBsEEG/AWYhvvJ
dRTxYhSJ7mO8czgDpZbNAkQa9coCqT1C+QijcdoXQgv2E6snUOX0FO3/4fH7T6Zc
f2ZsA/hvYYYfSDeV8vVmxrq/0NwhIbelzVQWMoA8dJO4csYhQSu/67THOpI6WNDZ
mJQnh9JNpdEpOdOP3YzhLPbS6PpLII2KeAknBc8CMrn/TT2wkjsOL8YNa3XnmZbl
GtgB6liEkGM0G1W7hh9MWYHudygZXxKyPqkeQBnrmosKrq1Anmz31/UYvj/wIGJU
0B0YT2d2eFjuoTC4158UoX9b3S4BUsbVmLuVTKVad8d7rdIKKU0BJ2pfBrcXLlLT
ei5Zq0r7S1iH6JJ1g498NDNT5US2iuYHVDpTwhRmeptsrnGVr7VJwgLZioII7SGE
GczJJMoIyus92xOyAs7bFlihosWjZlLv25/RVZrWJJT2xN34Qax+xe56+mI/cxfe
7tD9ysOzpnarlh7mNpNrHyA60Bn+bRmq7BXo6V7bUwLYJNMykaEzSbIwk4ILpqP8
4U3P0AaUCyPjvSDvkPqFa+Ia6w5QC5nEh5bqRxrTjFlDWiL/79gWJDuH8xUqb5sf
/e2Blaai/0kiOWUpQni1xb9UwEtN2n7SkZ7cDgGTpewTIipt/OVgod7vbeSFvWRI
PTmFQMSy42GXvqW8m0EMdiN148R9OOJLICxPevIkbvWn+fab0huZAgJg9iL48FE7
eJyPdDQjoaUP0SR2NolqRP0a/0nEFzwWQjQhvzWGg8m/08aaPlfPcrX0t1uKkUYs
wybfaRfW6zzNZFIzQzFNEKamQGmvydyJ9sL6GxkRsGyxgxWBHQ86klx0xhlBCMzl
NC2rlK4wl9mJNmbsqFKldKAPsO5AC9CNEKmLs9pPHbKaecUI0vKS7u8w6Uoc8mZu
EHSBHiNgSFdwBgY3vYxnipx5kao2F3m2/hAi+I0oFUCr2MufdDb/vUBbyX7WtcZd
6qsEKghH5ZdTgvwV8FM5oSkZ84YYhUKXHTWQDDc04mlZxEB/HLQb7nQ1OHFXWUym
lyjcHGNEcTMiETvQOo69JUlKIeC5KWH/+VG8eqwhclOUbDVgwpAD/6ULvPhuUN2N
eHzlGYDdurW2d7X/l7XpNc0vKFOj/Jes2VBmdDd79VmlvhSv2AJ00CcbF1O6sxnB
Ma+nxdGcPuWrUEjo46ztJmaEzrO6UcLaH4X4QK0sxxTgInyVpd3qM42bjLtbj+hZ
6MoXWRkp7jprCoP8Yd5wAYW/cU0/8WgdmavV6kpDCyzuYU36WfdeYeNgjZjp6xzy
sQ67O6aS1g7ME/SDoYTDitupkNBCl2JhiNlW06MPXCZ2/xhbQlQkPPejJsjXadCo
DBvhxJZBFlDA9jaigp20N2bRwaKb91Ws/k5vv6sGM7+RKoaoqrUsRGJYZ2qtenGk
fhNQLUESEbSo87BrSVnqWpjnXlX2Q8F8X295RiPS3zmons7+nBQ5k0QlBwwpkbvF
hP9fHUk1x2mc7SlVELpfWcurRdvp7RHxhX8E135rQfB+ia51KFM7F/JV3H+8gYTA
XplEXPLvK1Pj+gn+f+ukogmo/q0bEBtVzSse9C452Rloc5HXpzrAFxHwH+awGTpB
lHSXs0Ylad+nJLohqI3BXvJiJCsry0Guh0mKU5vh+k1HY9r3gOBJvGa6UsptXehq
FJOCVOidkF6uR7qJgs4NYAYC1iad6xCCa9q2u11WlCH46SjSKH+94L3I+6rxXUJb
ZZrSCSa2hq4+eSBOBdALJJI6KJxneszUvwwFBYjlnErAP8pLBR/zsJev6TVdJyYm
zjBYv9BPMqGm2FHL6WT8WATb/rboG46E455xrOCNgXNqamW2Eoo03cqzvmZNGrfe
xfxA/vYEeFaL20dBNzW6feAvnoZWeDM2xNf+kZcAFTHRcXjeo5/tMKZVTb3qnxKe
pQsuuVEjX8oljsrL3zYBxk2ZVJuI0HAxOtyoupejh0EqHhA9dIg5yWSkjNopvMwW
7hPixR1dHkL0CUfx3e5DyhmT8CvIpZYxIVlCqYtx5794VRQRpwZsPc5S8qnoRg5l
rO+XgBAQZ0z5vBdfyqlvCvoTzv+iORenDd8XvH8MmW32jyb+zBPV/XG+smL2Nr6G
3sWv9+D5PK3oLE4kxhVUyTYPhgeF0qV+px0gHvtHP2VfuBEikUX24hAENATQ2i3o
riGQwLyQGf9kJ2TO6XZorzvyqLfWwKX2+2if//hqB2DOnRDGL+3xdG3k2ORuVwDb
5Ts/m6D6znTmIU9ZImZns9ovKPpIL/OQayju+iUNu8+TFsCrYTJ5eyQW3aiS9alU
HtC73tF4gAhrD1904SLIemtUuQa+6qd8b+m4vrolooseuAmOr948McKTa/Suaa/x
rYIyt1Pc9w/F1yNEyAuT8wKKe9HBpQVr4X21KDBINq/rkRx/WvtbqjuXRI1Au7fA
sM5aj5EN6o/yJWtykhVoQ/csMWp5PbHW/aJoty+o1BNUxQqEl0TPzwLvkx76fCSB
bE733pMCSbBKzOlHX9FM9EUQsyouUrYX/2Ruhrru8RGHcte1ZjRXPK0vXTbJdknL
T/tJRMJnYfoAh47I4jLsDh2Qj4bQUd5A0lTnh316C/GHe16iVKlEl20iB3qX6oMI
RFfSy5hwQjW/17YfLQJIwsrLbyMfKuZUKUTU/qqg5RoFKU6V+zRHPnniDwxaIgcO
UrgKQtK3o7xPenLNgkS6xH/xvvmcEZVrqV3CgY1aTfo3jws8VXo4h2v7vnCNcEFx
RHkOH4Ks4eutt1B0yw1j/IFt/0UtmYke2yvLQoz/zvEvAzNJheQtblpBwOhjnjw5
oiy2BeSzxrCHFmlPzhC9Dns4pBZe0/9+Q28y5WNRnsqPL6iIacQLvxO1phYEgxKU
3wCeAhg0NCQsAI7Pqmj2BmS8qQ2duRS5lte1Fi4ApQzS8ptYXRrFEapY5Ihrw8ia
LDLP4CCLXwJGHbW4dcHQhKIiwgpFMS8nf6p2I5AjTzETuE4tltogXnKKy7O0/9xk
HtobWlSXPgizNJcZWPMOARCoaSZRE1yUoGUi0s1SoGUpO8nDgwZkw3T2Uc991dRx
ynxW+WAjYgQnom/v9FEB/YPzCQIq+GqdJUAEdnbtqr46dw1P6LIm23Zrx/SWK176
/MDb3KZeXTzoFM25IhqvywaRU48EQg9r2fMtgqx0ObC+b62+fq8hF+OUFkvu17ig
W5UymVP52WUlu+rlEIXgYfiecSsXwEqjaOCtnHSp2IxyAZVpmQQXbIqkwYBTO0qI
B6QKr2MncAZCrW0+X1GnskkPNZz3Iz7m30ZfM1vwqnY5+ja0R2qHmf+rPY3YwTCP
OEBCs3jUyWvo9/1io8WALTQ8Xc5nO90W+ZH09UWU+2X5BuVgeZq8mEXUDD61d+mB
98pRWgEgoUoNBGSe29xHiA7st6GEzI8NMJnVGEKdeoAIRIlQyTGGeX2FxG6lsxQz
p3/ep18zx4dHllLHT2IEhL3SzSQ6n/5XfHfZVaP5xMh9gzwsQZQaI193+ae21v/d
xn6IdDHjoD1RHut+jqTaeZAOf0PzePVElJsU0uqTO91NboUYUxEazHEcQnzGcdRX
bokBtl6vv7qgJN3rVpD38CjCI7IU8fqIHM/XWbA+dIOdRzGJSdAsil7MluKM4Yyw
5xbZ5gk9n1R+jUoe5FOmUrPOLIKWfq5ExJtVA+7nqtoV6ckrYZjcR0f/gT1g0ZQV
Iere1aSXAUjvLtiB/QLTzCd6YDsjDnVNE4+FsgCXOVEWC+NvjA3DEl26hf1GoUtw
pXm/LGshNMO/aAC5W6dBBXTxqTEDHT8oZ5BLkmQqVf1hsXLseJb1QWW7x28n/KWI
9giV3VV8KLc00eWNyBrsRahIcj8igpIfpqt81bgTxq3435wshqo7UCp0i/8Yibhh
UTAjDFblPYs/0boE3BlSNQJav3ERW4LDXvpDy6dzD0qQ2/dNUCB1kTxvYPlcDxdr
oIAXwLFVAOzUwtTBni52W+7q6ld4ZWPvEGxuvqFC/MCVlhQGmFLOzhxQYsOq+PoH
QWgqfp2dWpugk8MkYoApkv8PDPbXuJ9/ucpRv/76cLO8WHddLhGFnDQOerKoqFe3
7dj4Zg3chNqa/izh5hHNlU3osK7vm1mDzGsfGy/dZIfXhJ0WYmYeBSPpDHsvjZ4V
54gLXvq9HyQxHittOAdSSxjBtc/YZ/MAN1xwVG335dX3chB0+pU6ropcfQTxi8iP
Qpc40JmsbdOAiijajANDTZOXUg2/pSJ9ML7GucA4NrUgJi8R1H+bTc39S1WUajoO
9SfpkojnFmkz64oM0380g5p3DANczgZ7dvNGb1DdQ/KE7J1npHi6rn1JdGAGCDTp
Ssj2AJfBn4FTbK0x05MaqAnYQLozo6InGAtaV2EUnbt2nnsHzuAoHjFriogrxzse
pgY+Q3md5/35Z15VO3aLOiobXegIViHw7hO+fvcNr2ZcDqYABRh+QFpW2IgFwGOf
IbCjdBn6QnFuyuznjFcoD5Bz+3HthtzAxbayrkw66Ivh/TlZ2iRcXMFjlq1omsZ/
c+83x09GiuCJu+esNaOyARcG/IgQ3pE1zitYP9K3CNY2HjlCmfX4JuU1DxV+XOiS
jh5Z1Fy2ih/kIKF3dzLycPYMjEB3c6Kv6kIKx0YSJLl7/sILb7wUFdS6zjeGZkR3
1hCqzg7DQm+FylbiVzZ7EC3M8yIDLYaE+DEC61+Ids3BVGpj1eZpUM178VukSHLq
Pou4dr3Hhkl/SiCFVeri3Um/bjHF8T54vlocJAGxwoLgYju5ZaEUErKr5zECZTT0
kWQrukjMe3e4QADefcBCGrFMYIHMjYb1V1Mz3AGW/+0pM5Nmpb0Cd7gfX96hWW6o
RhzBw48OGKeEMIuKY2SQC3MalaXe7156tmZEIHjofeOvZ+pg1+n+YI+TiW1I0+yn
8EaPhnnNWbv8Eg8OJSzg/WgesznoNF6eWHzNbEA4itpzdM5a7mMix2FXs2XwSEkb
dapBml9KL0i90OvJOYGOTowRmTsaW2tJgwUd0eJAVD5NA+vQJ15vSdWIZMNPUXaf
VZUb1t5owy2YpXMjDpUVdli9bYPAGDaYpxi76Af8vK3WcH+szEiMqBDvb3cKV3GP
alW+f0OzCOT6ZF2bHOsvmzj7mceHxa1LMcQ4RybCGtgw6/Rl9w1osvDlQda36VWb
Iz8lV2EegLSrsuhC95rXY9J9dpg7MLa2ND2ByHVUXRx44N4/Y3zKRIEBUBi50zLn
VYkdoODnGgllCaPUb2+0pmZNvdhoxt665w4wnr62Av8k31oGg/FakYJPp6P1vtfL
pvaiU44oH6Jor7hmZHf94cAzHek+StIhKnodOWV8E+v9kAonvgcIGH9DMgX/xVy9
2h6Aov7IOHvcXEHxG9fW2BrD9g4u/VdFJIDrV9vLSPsxZ1CZ8HvbHYnycZhGrmtS
j3hLXF62hNPWQV+QdctoeUsEDFPHIZBx7ZvGSTabrfOH8weYCb8KXvod8IqxQ7VV
1/V1/YCFKkHxWP0YMvircx/mRV3FTMI7bSxtQzAu6wGpxuVe/eySNL/dHgtWU6fq
TQQjLZAskfLu8mKLa9n7Qukw0ullzyebYsg2yi5/NHXYHOqqZnf9aY8qa/rP5Gwb
UsxmaTzJuSfhdTBxFa1jVIvO92RiOZ0t+P2xAnTI9EDlQK1rGOxkLn/0noxIBJGL
YQ2AKv85XNQ4vT40Nu3XW6B33t1WaJriAMqWv7C+JhFed11nSUjaCmjrkgOm/oNn
Hs1Nx7+AhdKorZmC2G6aVLCWajo9y89lMJI9MEsqe05hpMUMG9s0xhOUYSMvFd5W
0AYuwSkl9peTJVTGQMbsaGrCXaQgQkIe3QuinvMEANrME/VeLQC03xe6kp0OeaMn
LRZL13/VFDntKbw+8HD3nCUTYDwr+fS3SJmQt0fdkGJzubSCKrB7FLLn25lSLr/7
aeeHg06y9lgDtAdpHIG4BAx6NSGUEas0Ac7ozdoK1QrHk8pkFTE5O7zjufpoF7Uc
PE3h6OodLv0O9ttGXRRCrTbz9f9hten8fFO7m2edjkwSy0QPm1VPrAxwWq5Pr1LS
2rcmB9TQZf4t/eUkLNBLZgUaPz8JuxcFaSHcKHuyGQfduwp5Um7KmacqVIgFuZez
3H6MDOpyhaSVA1SF0EGlESZPWySdUefh15AUgq3kileJb6EtLIhiILWLs9XO6A/N
B0w3fPWfppxb/ECQ3HeSZll1M68+6v4SEkgsJyNFT0I+g5a10/DkdYwgI2OnovmN
WaWNfID1vCLLc2/s3JMKrze37rsUBv2aNdYtVNA9N4o09Q5bPjXUfpHBE6DS7C6r
OJHmYl9EhS0CdBX6N3hBIA3c8suWmhLubO5aUpUOIKbd6PnEz9EcP09khVGlEa58
hJJclYrD9D8VgLQe53OchKdI1ft/ou+bLJGV14UBxF0CwqW+vJA8lBkh9YdhkmvG
L53WxH7lPoulb1WPiW2VAL6ncYv3CX+ATGNYOxDsew9WJ100C7JB1ff5o1++ZJj/
zvIDJphYlazNYPWli+fxkzjawn6ygnQhkmMDwQpAJ7K4+b7aMRyizKllnNs8eCne
fLE2peebPVoBhlYqhDAVS1NM0t6xmvYavKytL7EZhLThAtORMuHtz8LEjPIeOcmJ
64icqSJ2AB95lGYhdRrA2j6quRNsGlpe+oW4/Hbsw1E1APk48SXLwBH/JeAUJYXQ
RAtJ2NhUqd7uv191xf9+eo5c7a1pZqDWA2iCl2P3wi7f0jByGOHTnGGEhhnaWNDv
HpviIzcIet1LvYNN1JYcb3Fho7r4ETa6z2jSoM85EikN9A/qcrhQUg9DqiqouM+b
O6NqbHa3okBP2Nrp25X5KHLIOqA7PgPqAugJEFNPpLodapWshODrhq72N2KQOhET
OQ6jhOWUF5bZklocKp+wEahn+3ikhzxbm/tWCM0osLEDEZ+u5zdVr4q9h+1jBoUJ
WN+JJEgzh3JG6uYDdqVflj/DgsRuZhAvbiA/OCJF2hNjtKxpRo2T/iWB44ugM1nV
RN4smCs6gCa6Q6BQQ4NSJEsdzEEc8A8WvkJrPGqwgapnlLvKTH2TBYhW1gF7oX3J
CGnGJbAABQrrLRX6WMyqfUTTW2KeyZLL8s/ZNmmpz9jvnb0GNAeTXQB1vR4Y/xzQ
JeSY5P+t/TS2g67iIK5mfAj+R+tHcdBxMDFzuTstgoig3ZztgKfjPL1KVuh3C369
ApYGlvcI33CVkC9RtOM8ZZ8Ek4gkdynCf9pD0f3Z3vnptOYbPxUWLjuLZTQZuqP8
2NbSBzDLlEfHBzZZdrHKU2hnPrvKZsQ0XFjd9PQBH1vbqPzDXh4ubKc3EMOWJKt2
Bpp4pff0UAQfF8+YBMJeUMKtSEmHwAZy511RZRleFDeGoh1CYbIcIekzRKCtAUEA
VKjoiIztEo2uoqSrcaQ+ZygtH3ofLCGOecYeMeSmIGkLe5s9IHHldMaGhRGWL9zQ
DMmvaLerwpCK+sSi9wkE1zRMsFl/Sro4tN31K5/mL01gk8meuJL8Y4y0UA4sB2BU
cclxNM9Qmtsja3tiop6GHVapq7jWnKD1+U+V5CM6RDywVMqif80s7LA9hx2CnizI
CcgRrNhKsC5Rqjw/BCwzhZsYTvcabR5itfHuctSBGj1NHdd40hdsh7srO8PCLyVM
dJv0qU2A//Dbqa5VJFkX40iZuBkMvPR6f5dAT3CsiraF0M6BkvVivl8JYQnCMuJX
KsG0ptByScE737+P04/3pxYvgfRa4JvIqcaD8r7TKOzfVpLjpK/lFsXHpxeQ2j4Q
SxmQncv7GxwK7KaT++LfY2IGxfBtpa8Gkxn/4jX6nq4xYglPB4Fzy4zegd/T/O7H
pip/H6yheBMS8JnHL95OrWWzMd9g5+5KnAcZfZRxlyKgxtsnGUoFeoORXpqFim3x
QiZNCO5o4BN7OMskaAby5nP3LZNxFGvAUPetBeWx9mEbFieTRqea37IGE5q+ZMW9
5Dxoa7FD8m9iWcZQBAbDsWn8U4boRpMLx1KIQcfu5RiwH5mZd/r5E3C1MXqWgFUI
h71B+5Esfe9oC1IfgHfsgYQUsPzAtp6DqAgAKYI6GToIP23W6209LeDyarGTyDzO
FRwZGZ2m+3xDQ09Erm8MWPQbLLj482OU/GAm3POyvEZSWQ2PGiNtQrNjiCe98jmL
Bt4/cN0BQiDtJXR1syF5eYencXxXvXZMdVIW+Ft+xDZpWdx1uEpr80at61QXaoLU
2fL+GRGWXXyFu41gwDj7u23MATNGtjY45l+yKSrsm3f/nX8Yd6VwF/u9H77MHTXQ
a/sgMd69SRm6xXeBqXin1TqUv49GPd2DmanMXPyCoPNRwUrs09Th3IPoq3jQ2thM
CKIkvTssFo1rFfSJ/7NLNbZaEmeQSMzNaBrAYa+ERVShZ3w7csOGOja1fcmVNKOu
SLpab4U1+U9qqfuyOcf1bZ/f2A8OodiQ/lBV+dMWqvHN45uVsqlNq3oD/6qUSmTv
z6vRPkLFm2v3kMkAFP9p+cc9qbW9p0zrlXLjx1Hrbvk+TjzQUbQRfkq0EYp/sRIM
LxsVHDVMHXSw8xI4h0qRXqkkCYRz6X0/XYD16M0Cn9ob5q88PTrV6RD19eP44kkA
6ywestnw3AknY5iWIzddropB6AFU8/3AfEIS3EXr9QPDgPe5lxtCKiSbe4dpoETs
8e1poJsECkvOmxJEcG3/atfUb6Wjyax6w4ujF+tjBjeRvvdSxkR5hkcWIOD3BRpi
CytpzTB5k8xsnfzSYI1Q1N6vGxEaju7UlBKk23HBzTN/7cZWbl6IJ3cUgxtjSBi9
Gg1SL9m3VIiG2WeeJZIyYM0gWuXrFpBLNaHmQW8OBZBzQBshAKcdH7tzAp/ZkfKp
+azuMfiTxTztW/oQc9VMvrFaiMEONN4samymRQlf723OFoZcFY/cQMLPRBxnYs2+
FxfyuAcEiUDxD9+VN1+7ygfDxgihOsYws4xaqmz5cY8FaNd1ookhQqYWwUKiS1AE
zk2haDjmghptZNNAeONGh5ih8X7pXsN60YBtvSNiP71qDAmETAU+ws+wn8NJNN7o
SaXsF+3kjgYzTESoir3U271IT5e0xu/8S2Jk/7ZvmRL5N1M+9jz0acc8T/IMoajy
jgylZ3dn+mzDQQ6ZIKQqjtq/OTNsk8wgtepw6IixgAUJjSL8q3lex6G44zbShppx
eoRRQD2Ua0h4VR25gCfUR29a+dVT0atECBv+WbbUA/pCQGxWs6OvWfpSrrcrj2N5
IYxnqEPywouKiSY0EkYQbtcT3dK7kLDiVdG+rXEFuiwsfhXG7p7r5B7AzsLkCk11
n4KzYFqQ5RsKwZOXnfYWMMw8dtCLD2BlkJ9WZP88teuVjU3iHLxQmGoIyoMGD+JA
wNK5FPML6031syQsAN8HIIA8EXvpCS5c2CjBeQCQIAMMPQzRZKIgq4kNLrHTegUM
u34WCLIKExkbCZllKFX9UVCaRoD91iCdLhKzHDwoMbpdI0MjCUeOKeNpOIgTA+GX
5FBBkS1aa0HnblkkrFhvL7UyDudsTGkA9EP4pR1kgdk9Zpk0M6tdeVfRd8cucB14
U1JemCYHCRLZlfti2/GTjQMT2ILGwKEJ/Ps78ZJE2mdrrMQ67TlAI4j+bwqZvVb7
/N1wmVrkDYug+bBnnykHSJabh60Jw8LdDwBVysxjA7/2VeSDF5DFB+MpCgcuR1fL
YNOUdCsNwYySDIdLKykxINcPsQZFrBsqzpRLEPwwmUbdlGUeju0Q3O0Eqswr02Qc
8O8WxIJi0MDu29XJOnn94Y/wg+QW3LaBOFRJU4AngyGL/X2ZZWZUjgSFAt7VFJEf
wdoOBtZz0EIW//LHM5YOu5ugEOQ5naXM6VxlGGJizCqznCI3Ta0Lj0m3PHbKOIlU
AstcwTNQgsGqWStBQddDcBkz8Gv9a3P15KMYo6wKSa6jiKfJRmIaogANoKb6nC9R
Oczkzvf2dYF1jJ4I6V+LaXrY956BMizbZusv1aDCob1+dtcFKVYYrv8x+RrPY73l
lPJBVPhKE/GEoZ+tw0N0rjvVoraRNAJlcY0lnJDnEOWM5iUFV7ilORj6dGZCky5k
Rjdjdy+b5opV8oHphRUnl/zwGjn6FAT10tQglc00zTIOutkQLpVhyCoCD4Ahu/Yw
rf5LLTAKCYi8Ih8HLm78bUbz/iw/T681lttd7Ai/5nI0EHbIY9TOSVRFa0ef7l1T
q9Lks6NWnOPogmy46dbRa+VB/vhBNRuApp2aq3x1XaDPLHv9wmAfnTZzUTDfc2QZ
+9WPhUFVBf5CRjttcPteotbW1hXQfy5ZFSgiefQlR7paM+36s0codRYMUzaDOXMF
HVcI8AvEmBuopTjs5GHBoPouiHCGAmDsuNpUrt5mRZOZkdjiEq08Oo5r7wFGthk8
XdLg6wuZHLEJ31j343OU+GtDtXZlL8TrVPW0Np70dhfKLMGWyYHa6tNjOpyriTBJ
zrrzf1pXE9XH9J5HF8KXhWgi1/Qj1WSQhbH8aFMTB9ur6WHZnMM4Hxx/tUDdAxnP
/kwaXVxOzZWJGe2YfBM5Nnd5LspnjPsKWcIUAUHFbb24R9ujs/9Dg9x9nnQVAk/a
CkhlsHa2aOwwHqnzdyFX5IAX2u9RTxTnjBVg3XP5cZWPac5kr27bHww6dYsxIV25
Ll5KDdWV07TAU62GkR5pm087AASu7GJtMVDnhJeZ2+C7hr2psKfO4qtfe1fcm+dq
mCVP/5rfibc0x3mpJzIzgpuFzHMzAX115s/uGg7VFkfN3PNczdSjct7RyiWo2ryM
adyuoBiCCxLwrgY1pHGmv8WhcS9SyDCOwT7Pk3NtPxK9xydCY9Q3CvhUhxplZ2mF
nTnj5zmXoOGTbHyGuDvIqzAg01PcX0vefzw5KZqoi5Auhj44g3C0jJwxRxoMAHZH
CSaDwdwQEYMMx5NNTPto7rksDPplZoZmkEvGpyVdjS29cK8NzXI8MdC26lJXCboX
Qs9R84yd9QR0QRO0ZiwJbgMbBd1n99wiY2GuAbHu6PXGsSRjU3zglFTibtnDWsQ3
Zvf7alNJNBt4NwNpqSj3tZ+1DLacjStEngLdXOtuNJ4bpO57Nj6o7YpI+h7KkAaI
iqtdYNlo6OteYoq058T5PHmJXYRs+T/U6bfIT10sY2qf7pW/yo5iMA8LZzZtvP3i
073PQCgdIQq/wjGhQRcRexkKOARctJcTtA/pAV/QvWQJYAUc6shTRD0xKzEWgHh8
GjizhqfvBJYnEtkoRdALe1CpOPD3vd7Qvs+h3ga76nibJsrROUFXLQwE19vBCKEB
oMamYwLSRac8IUQyM9iRx3H8bXG+60XUUBvv0xSyCmBLBLlPWCIEBFxHmq6/u/pd
SXNSfG8f+CvmKqNMqEOS63cvvUDp4aqoa2E9pspT8z65jFtrgI31mWhV4jIJmag/
n0rLXatvYwcQsHo1KP7vWS3R44Vz6I/cFzgaNuTiooSF/5VqG/D5cbIuBXAKVAEF
KtSAPW2rsU9VFLQ8vxfw9bhWTkhSpYV0+vtR5qjkV8+EqHXGbq7eOZzPo48XeMKZ
BImJl84BuzbU+0zBlKPSwsd+dp27BhjujxtnMvkl4R4NuLP9vE8Lva+2OlE5dIKH
yoSWSHq2+mA6YO+KlKbNzLIi++n9oGBn38x4sB4K/A+xwvDfXF3H/z4yAYb+kvwG
n12R4TB3NSk2BzCA9vo1+EAmuikxbipqcjfcTwhjN31fsv2c0NJE97Q0FJd9O1zh
ea5FASUwcd18RI5ZVdP83Q1TwPHbpBItar2fkLaMv6Y7GiXHHasck90o3CStFJWK
+btfdk6P0op6JxahsPQu9qo3qXuuZwJiszwKHNQCoOcPwaUOAe3secg8LyAmK45b
VSW4QkoSusLfNhihHp4dmHwgJnhXFU0fqftmgFYkrxmxCNdi2QJGYyBNRX2VjP9K
deNm7MaX850NfLFXkyr1MpFn4kkLpSZVbQSPgQTgsBtmQpDjTT7g1tRfvdpaNaGx
QslpmKm/2Ze+8Xe3OFgWaBlVL4uUEHW5CFy3DbQzEwQjwtIIp0loY7qKYFtqjoET
cN3WpmZA9+ZTCGEvQQx19LLxYgWYbi0zhupwcemYODXp4a4gX1Jmu9x0KndWnUrR
4lKy7XlicjaEw988HON/QIPkzkdZp8Rm866ArwIKE+IVZ9OP24vnPB3JJPeZY0nz
dlBSyWNqYRUXiaXi7EWAumCplLmUFL7C5Sp09Q/6rJNroW9/sDiejziHf5XYc+1Q
PaHU8LoQ/F4VFTEhARsvf7m0wnyYQd4JwcGIQ0wDj7N/KK+ERHPEFvNImAZOtwmZ
opXnxVsCqDM77pZh3ulwV1cK3FGKu1d4ZcmHvhdU5ugmv8duRkyteclDi7tGyNxN
vNxA7x0YkQaYoXi62O+98A+IXhF/Ig2ETRfAwQptEAohEhwXBbvfa15+0T4U+jp7
IgHfHVfKppzaNe6Bw/K5CYaDswoBVWfaTx7t6iUFI0PQ5QrvPfhn/0jH+qMsxvtz
TQHvdDKo9ZxMgePDmM3PwrNR6YwAFkC1MrkWVXxeg4d8Ww+FzPOdhVAKaOuGcJI/
6qE0v/cT7xJOjClKqplJmyIClgLwNLeKqmCKJCFPG8VG7O6NpV5ugWC9ft9SUlwZ
eeaQCRtmxCzxiEjuCFAxKBLMJDQMD2DAsryFQN/U7OPo3jfYhuo+Adupb7YUBnaE
Stx44U2pUvTSM2ExKeiO6dZhEYVoPqg2t8AO3mTrSGkoxmQF31DebqwqTkvr4l0y
ENh30XJnAsGZGN87aqr4iU6dVGX9VGfR/Cym8h7fI4csBNjhdDX1/E7DF1w0RAfx
3qMOxHIbkTezmNimN1lIbORlGxXSb2ARJBscfjnmuet5m2zxwj1ZOvcYx6Q7LcFS
VdXbTp6FqzCDyI/m1/aBNCuyM4DgNV+uY7oJrqo2SfSwJ9+a0WXkpZpqfhklzdRD
0JfHjWPS39E4+Dny/G8FGXPrVfJ6aXuGwJF3N/dXJZQXu7gVHmiNNI8GwnzdfBg7
aPuOeYO8zs6FJNgzyrVvKto9y1AvabOcbd8e27Q//FZcIK0LUS9MN94csFYns/T/
xGCZ2b9vqGbYf6eoFYrYbSiygh2SesZ1D3G44n/r/oeEUnfPBYWvGfQCx8bCMpr3
oo6AL+Bmjng5xzVm48CAGDktVUbTgXeeb/B0L3k91Rfpd8Og8UL5K1FMe/H2jCFF
qr3P8mWHj8jAy0oD+JNWD0Y/jl9zVxkhjsWS4G+QevuYaIiFeNdJYYBmO4gW6kHF
qd4y9reGOuBy2peIHm+5oiOggAUaniEAPfIYBbTY+I9MJtspaZkp65WEL/AQxJr+
PcDH6PlvkJWI9BFmfIbWrGK6zK8YFqmt7GYRwRXx1VEhNw1Iq9hStCofQMnxh01L
uTYx/2gR8Ijt16+VvcJ7vKMi8OpuPcIttTKuDgcEdvFin91qQ9T5TTvmJPDRw2rm
dIR/P0W5OZjXXQvUyE0HnKFKl25S3v39hWdq0TrANixYBRI/IYRe3y99vAEnJ4Bk
3dPyhX50gUwAskJOgTF6gJU4iTmf1u6bWIf1kovgu/mimE+YJx/b1cWW40ojluPb
VwOj05PKIOiF9wzAcmxPRUOTy3I5jqey2ko9lCj2TBgrRhKBbSa9TbCPuIgv1gng
tLS5SjBJH+CH9n6HoZvcRSFMRFPed/LspFvFepHR8qRO9gf8IQpffcBKOxzc5iw3
fwvmpdLsV1fxqRpF0nE3j9OyesCG7KQAC6aE8GpWpputSxsdOElPOlY9qW+z9PBK
OXb8gsWG03l5WvMsODkvTrigNiguH9ti6J8HYg5A37sN4KJIBkOsECTLSsh8wCce
frs7M9tDq3G/gojpzwKqPU7TGHubSFdZCB0iMnXEuLyeescQKfVurQXr+2dGG4S+
HUWx4U/rTDKJ1NVqo1VgiVHKlGl4PVFIx8snn3FzS8cAGRCsIGl1/sW7qpIul/+n
x27ZGDZP7gCIhf25GCydhIatGT78P6JpWFApzsWIOKLq3IDXFfYNCV2yPWLi5zlj
0EidIvFDGdIHBOPtytYqNIyi3IacaqyNGs6M5ElFN9EHD+cdand69XgaHZzUHIw3
pm5dRUaltiDrko/OhDKl0PvKYhEEBhBsDwsSZlEBjvnD8KASiayVGVpEf72isX62
pzRU5FXVnHaWoDi8xen/fzq7xKf706Y4DTtDJC8Z/byOBvRD+VlW6rfrhkSFJauW
+Qk1Snr+tQSoh3WEwAESA6wH28rEQy9c1xg9WqHEFBXSkCyhFqpKTwpL18Pu75tB
53nQuBnDhvP6FYkOtolZdUoefw/Eze9jlvuc4NEtxe2nObtZHCMX3xvT0yJOAvc3
ACPfbCHWpFpYjVtAKnjLjlk2nc3PSfHWWTCf1mz05Hn5dgKyzkRcIfQ/OQdvnVPm
oVShVRFDMoCoHUEJJtxGu9zwwKpVsx0zaqEGAEOr1Z8O+UOqMm0bsBIiBjP3RFRO
/ATZh4SCCDWdkXfd5fkgWEjRL0i93O5X/z6P4POPUrrRcfiojA17cBFW9AvzaRhW
Nl87b9YXISGWCuVZBrwjWbdAY0wNu9xxYDIiFjC9JXNYvcjSqNYIB0BwvC7+Hv0T
ZWlV+/2uWauRx1evVNau2rQS/rttN9m7vjonMj+7tJ4YP6FvmyHXz4O3xpNZnn7c
wt9qEVMHfW4rz+9FKsUX2gqY993e9qCWT8Gv1vooMEUIswR0WFxjiGoPhcWROs4j
KCS+yyXKUk7PCJ+gbrPCegXTRdwHgfn+cdg3YeqpRCMKfyeOwy7saSgOeaoPv+01
ytLmCjU2KA031EIeztc/QNflt0WAeftM6wIbXUTkC8BdyA6CDIfMMaR78pS2JGpE
epjs72pEL1vsNb8F0CxRV8iXOGkb7W1WKc9OtDkr6DLHuWrU+x+hoCfcOyE1zBIg
Tgldt3H6rSlKL+ktqzT1fmCB1xUHQ9oIjIu0Tu/JJezYrX/eTz7hbb/DMR7h0195
PkU6jRjnKjczqJFLtM9qdTbc0k+Y1fUvc0SiUZm9U6bUquFHoGMQYuck+DnfQt6+
IILnVWgQQrNI/gSL9oia6qQg3nkgfWtZk57Oia4zwRyUR/Dx/W7x8jJrvC1gr6YV
HeUBgsoX+RKhbecnqWbRwB8ZievlTg+J45jHnGNsJjbuWkzHKTiSD7+SRh5+JBtg
spTN/TizjRaV/lZ29x44fNklA6bIdS3BLasDbBpWrBA/saQVnZimjowhP2mlYB4s
1w+jjY3lFRpm0hUJQjZhmEQMOxZ9T0BZ2uRK4u/+oEfOznJLjVBImOjQ3lHlzYba
SW38AOGgmrr3f3z6n9rIZT+CO6i5sIiHJNLNU42aKac3XWps/pCpERVmyXqoV/54
lIC8cqfiRhvTqbg0yoHqr118220eRqnkGRZDEqtYcCcqF13zBRQAvJRr2rQ+F1a7
iA3Z6NxPV9bqK22n+waqYwDjg1kbZYOSB+KUDaNtWzisHe6a7F8c6dIsTG/6qeLS
8Vs9uoycxh0RW6FwyR7ltZQUWRiwVNhSJxhciLSzemcsedHzE2ln1c8kwOinQJ9G
PiEwf4JaPsQ6OAdOqQrZU2mxUdP5fWUv33Mx4jsN2H7xnMr8769/ddj7PoQulgmK
KKRsdIsTGOW3dEs3zbLJx+o6KprU6vQxenkIJnKlUzXPA5vOQGKxeq7Vf2H2pSDt
IKSyN21D7icBTg0Vs2hWaOS+6GXJ6mfIuOwy1LHAm/kW+AUxxQeBdQ7BW2pSlZhA
kIsedEggnj6sxWffZrhp9ZKuUVNRrpJUWN56iPeZwQzv926f1OlcJalmJjpZVUs0
B7FlLKfT/EA2EtCjHASdOzdIUCnx+nhlkvyGoJTLXYivCgFZJXQ/ZZlcMPvKFoRr
215iMeQU+3jvT0mokOFNR/ubDYXgwWihRMDrxeNYiv1wS7LhIfewo2RfxX2JqKSa
SlEslN3FyCrjt9JiCZsl9ejs+G00N0ucOxVgF2u/bOQT6YP3AC1PvG+HfuFlikgl
HL7wQH7zK41x8XJRGMZnqrQjxGClUICSxS9WaSDZ7VPqrn9croEixRmWSm1Cskcs
QC/kEkiDp3gYsC8fmrcPXsce4M6W2MP/2rWuR6+ep+D9vbEpueco3hhLCBEyufFt
X/cB5aNMx3+cjkQWJfucTOh+jQTSgeWcuoaDxakbXJKYKkJMxKn+KszT4oiuNa/Y
L3UGnhpW/6tiJgXMxE1lq7pZwuz+7fPRfakakZQcb3CDO6hqVTZ4NKdSsvXXNQfZ
Gwvbl3VQuKmXRaekHjoB2DpX19Xe+GSX2ueDZ9uozDXR2fw73RMKWk18iraiNwCI
nCeavWeVKH5EjFtWNBsplzneSPyuNUE51fHe6VOswQQ8k1p/PCF07SWSXNkWpjVZ
uSsSLS2MM4hfZdLNFasqGq/wshilvEP1lqzpw4kRZf7sN1jZWV2NOh3gz2Hd8sD/
/GJGZjRr0dbP3zMc4kFzd3pWOB67KU4XfsIEIMwQY1bneeVM3++8nlcfFiy8TDgf
SlOxmE8p22HAJzowxSap5yf/vuh+fhIs6HmNc3lSb/59mrGjiTG7D3VXJfZauc27
4uFOBFoRIJugNQ6SIUH4So5qYH+G35qG6K8U0xJXVhoKvkcsclIj1D+chOfYQ0eZ
dKHNWFHRemQoauTCjJyNEmSU/uJe57VT6IA5Y5rTpbt8AoXXKjamTgpkMhIdQwHw
HaR5zE8TNSeDco1iy+44p7yj2vJcG7NskskrxdqgGpUbhSgdylmpHBTFHI/PLkOc
IBRlqrMz+OCNjm/SyGLYmT/qOq/Tu23M3V3Q+DEPQMeZAqpKMIF+hCZlCC+lP9gW
MymuUwF6ldCc9Zo/2wVMqkVwxSxDQUgq3n0fy/wPvOUYlSZLSsvK6RIph5SdWgfC
FzDydfIfzT0FxI9Dz4orJSycSrSkxrN2HWkkXac4C0VDVe1w75lWKYsEP+LfuT0N
m0MXyhZCWm1VHN5R+Sz5dEZLTnfL17RheOBS0wIpd5d7kaSI5GBS1phYfKezQE15
RBDaJckMBATAcv6NiDgxKa1wluFaJDAGKt9iOJOto16yP3UjjEFMOpHZBjR8AP0o
VmRz16cz0HCWC7bPzvRzgbKsj80Ff6fzqNw1FRHVU62TSxCtkXlGizX3xTB5L/n8
+aTGScSWk0xtnDCDUGz2W1z58bEMqkRVPHX9Kyrc/Rn1MoF6awq9rAIamyqpKQVs
jzMPkqJHd6v4aSvGBOK6Bq5BPYlanq6OjOjc78B7Y6U2WqiXxHcyKjp4y9PK3y9x
x1zwObW/+lBHdbhygV9JniFpRh4UzPXZvoCmb5TcUhpRp2w+LQ93o1cNzUtJxO9S
hCktId9eHupxANb5XbhDoE78+cKzSEpuR0H/Uht0b/STwVHpC37pwzGx1FGgLiy9
kl1mW1jmVgdHX0D3l/vnJ68sDXm504KYqN+s571oM/C1Yt0z5H+X55V9II6PyEUT
0cnk8tKfgHVDNus4TPAl1dzNJN7qpbwokkGEAZyBf4V+uN0VFXpr9seG8ZIHm8pg
byAA8GBHtrsoxL4AAYHxFxv0ZSth8Arspyn5FoaqV8o2q0CZwrTGncWvba9GkH4P
gcsTWfAwxKpxRVsNh2M+hoV8IzxSKa/xSvaENT/tvlj4H+KOeGCCbqpRp9GJDsw0
G620JleNgftP024KcDMKzYBPxgjYGvbW2wTRBr9AHIvezYePiWU0YreE9EWzCkqr
DeaG1iuoGcJAVV1hrtWeL5JvQEtyn04VNsiKD2unODtGS3xDPHCqQRWD8ERbD199
oNDM1tu4uGuYaYH/KsNQC3pnJYN22RykBFNMNdzeVa/dNmooNWLzdBiemQBjvmlh
udvbIr9DA5wv2p9VkIX6Yv8A2jfNLnZCoHSv06hUxg8Es9yU84vkXu5+01y0l6QY
ZGT06+w4eVWtjnM71mMZzfLdmcSwcdwetSuEYprOhg242VS7m7IZVzwVVyGPevIS
U/5t1PTlU3r8HtiYJ2Wp0IRCBJlqYTHBiuIuZ4r94E/vSD3yAX1Et438vLuBi/PT
Fv6DMGX3BS6JzsjgAh+szSC+Ppm2MDIFcEZ3nCRMovuh0BO9FymYakk5BPHGqDd2
hdCNWoWSrwHpobE2ofcbP/wbne46fTgABgFFP0h9Bkyo/oJ7Efl24I4tFVHIOuon
59nmX6Ev+aqg6sPWX+gzSve5N9lyKHMVkDE9TaOOsNeM6FqYpVUXI/lAw2fkMUIU
j/Lt1RlJxxiwncOWNedgvUFIiBs4NkMrcyhCksmBWp0SnduWxvDJu4CRsqVbrNNi
hwmGFdBKQeRayWYLlLXOXLHCFcmvdmo39g88mAlaqGI0YsjV8p9GizWKUyu0S13r
Io3oaba5zjD7ZFZwRX/1lBgAFeoSxOYP/9+PaGlyfDdPEq814tsEAdeOLnIxqLJf
FM2l5KM6v8Udn3rOIyqLWMyyaZbXgu8WmgVUB+JRUtwg5IY48Jr8xr0bSngk5ezC
VOmEwOqKLcGG0YWsK0OuF4d1Kww56TjCe5Bhj6gHgi3RtnGqykXWuS4SD60uFtMT
ffHeFAroIvcFm/K7jxO+25sFU6GUEq99HFknd+aqsSRJYkZ8ebwg/vcA/8Xr3QlC
yPEK+5tfcip1slLce9wZOKTikjx0hZa4A4O4WagrLuiCXjzD9rIiagZMGgSnGKoQ
92OepM2IUmwtzS2f9wUZASkYfsWOfAdN7Hx+WGX4+jhVDKQHHFN85PZ8+RHTTJ+e
MlVBakErm1UHs6VqDDWgOP8DkC+LdQtQbVaAb10bomjD55IOqejrawhekN9CjwMT
E4UyNot2Dk+8xn8CIIAApoh+53aLD8T7ClYrfSrJ3nTVi6zx44mD7wKMVMB5fZWX
WQ784KVuj/0P1YGSBYsN2S8mlMR5FArPauS7y9HjPWEZ2k1U35/XPzIGt0SPLTtT
TFE4QbpG0ViuSjTwQALqOlYVOBV0nzwjxefCffkC+ly60jP6riuORIV6OsCwc9wY
4Ihde3B+FOqkm4mslhQ6Bp/BwmYOC8sYYCySYoGwtTe2m5m9CwiXiOQcZ2T34v0I
LcZCRNUC0xu1rXSr5lIU+PDltXkMwvK5SaY44QCXjaJiYErT0+J1+si4Lbae1mpm
EnlTYFD7503OTzsxDzQdj5n84xYSfqGUctYYwXr4zfj12w+naskJmcu1fH+y8uHq
o2HgwaeofgXyI3/7C1E97Bs3SEW1OzCJQKhCg8JoFDmmIOOqhHwt+d5XO84q6Ebn
dc92RsHapIbRLTu1wYzBAWP5xAU/752Yk/dbuJQH96UR3W28sUvCkjhLh93scD3y
M6Hp93ZzypXqmuw3S6JskQPYU71bpY5IyFCvm9qpe5xZ3onCqWS6Eny0b8h9kC5q
AAc8x/x/pULt2CCq3mITQWE66RWn3ISQoBwGPoyBScG+E2fBjcFbggeR5/HipKuz
a6wPfStJX1wUjrft+cd7U66/u9YHguGxZ6Wmih/T3eLPKyssTl4GchTtrxdHqsOa
tVg47TJ/OOh44ECZVnIz2BVWJI/hQ+6ZzpowROaPptTgAfA4TrYenRIV1TXJeOQZ
+nis8/72568V8wldZ8+Y+hp7Ha7RgVG7rkIRbvVgi981xjg6utTheMvIOJg6zALS
JvZu+bOftPPqsyoWS/txUhKzInQMnmKh6+tTzbxrZEsgeukv/hQGm5ADe4O1hnjM
LF7nhBIMArLiBJH7fSySXBVEo4Vnwt9YwNEO6FJy+NrSqF5kXeLYzCnOkfOtsqjy
9MhoMzTOLalzbkZ29MRudtRGx3K3BEnwYb0QyLPgP0Lr0V7rtvlphuB0MiT5ToLe
uzBPUUGdhsezOgMPGIBUOzj20f5DBTQIUU94v/8ypLi72nNOuxcuTSLC2d4H1O95
icigLYe3Iqi9yvg6ld3UXez/pX87dY0Q5ZD2UTJFtBWwljCBpRoRypMX07KFMP3R
nfwdjtE5hvTpP1BkxRrJPY6IsK/ZcuAIztf6mfuZcKe+3hPskb++dlF4iVZn3OQd
gu/NzhITbsJrqNCHMAUKmD8WJc1FZ1PIeP9BqvruQz5ZC+MvkYoXL9AD4AVJN69P
tCil8f6OIL/WVZYuYJojEY+zGw6XJ9Zdrg5i+pc6x4OivaNtbIvVa4TWwni5buJk
Vi+mP7Oysad2gqrLhAtQ+VMBwGCWjcgXn9oV7O5XwXe+x4VrDy462pXX05i4NdTb
W6k1kBdCidGaw1f9czwcxi6Ymp4M/x9zeWMPmwrmWIFIeU/DPNZM2CGIvk5/yOxr
U+9v3dNIVm7c34bQ+YNrs//fNSSaopEcc+rzK0f/Mi0PcE7NSkaFp49QySmIUmXV
+puFPf0gWzebxeCfn+88xPpYRjXIeJFSK5L1XAPCgyjdzmtDxsjuic73+kPz5oD4
jyHqjwUn51SyMwue4nE44KzDBI/x9M5Tx+1WrpdHXsdemKp6f2lYt8ymjlWlrPi6
ySzXbi69swXjh8QxdGg8U6EDrZbexPEZAa2IMTnvW1kK6OrBekqEB4GiEPOJfqB/
+SYeyRqjW2UCx4WTiFfAfSWOGS+yayP4NM4oyZLNAtIGMkdpoWvLHy2RR+pCXguH
v4JaH2WQUvjq4dpIu8l2c2EXoYHWr76+euECt095lTVxaqPDd8to6S8BxGkpG0m5
BOKA01cvZWqHMmsj26dvAThLd47CvacVEm7q2ZMb4ppW4Cde3I+HP7MY9lK5Pb4f
OTJazRxLYo+qDJ7BPCxjP6eo1/M1ZHuj7/WAOiJLKqG6MfrIbbH9aRq9KWYVGXjz
2ppffzXhKBh/EBXZoFH38aiKytUZd+ICQNF65FK2mcVChNeRLDCVLqSomu5shdrA
ydnbmeq53Cz9+Bs0KV+c8RTKTR2AJyV3FxW1ooPqWN0meBbRGxIFlBXLzXnGXl/j
tXuh8eo+LG/ZfJi/VejpNePNr62S7NwjyQ6paUzcVIKaqWzC2uNPHrCAZXPseFv7
LgTSihRkwUv9PRD2stfw9B4ILbxqwlArXJ+dh7PlyInRV30847E2MsL2/LoKs+ZX
s6rtz5L5B+9/3IeOfS1D4tCiUuxNbp9fD8xIqLdy3jLabel7maU3Rl60d1wyq0fl
gtDUW2ZkhN18OAMOHA9Cv8obZ8+oEhqFZvxlMt7E2MO0Qc56feXsVLsEu1Ax2DGa
2JpUMmmT5SyKz5Hy651cnuKvcSlJEeEff0+iXAj7du7N8ttq8XEVkOqBis60QCn8
j4epfCL5LmQzcR+45qbr6mAFVvmOlHSObuR7E4mfS0Ti8Coz419RQPQUVpArJPGp
A0F3I9jguzNu1SRru12SRgaJ0uQ0p/gF502nn625PRx3uDjEHUsWe27fOaTAMMd8
uj405hazwTg5vurJy029ezMuW86uL+Bzhm64rg+KmfXZouJTw6Bz5BJCZovpJUdB
KMrNwK6tNZYyZRodGyVK/KEYS6wj77GOxXawO0ROHen3HQjqxwCHSp4/PlL7J3is
YK3kgECW7SAGsssbxGRgj4fFm16t499y5cNYXL3zZ9uJHTUHLSifkUDn7oyvMEs6
FHlvUyXDdF/W6Imlf2qRyuTkqU6b3JHHpN49A7caRX/iX+rdHflLclVjFlbtvpvn
B5J5NVINJOlve2rScNaAaYWCtpeWk8jx38rQXpy+3TE4kIf+5H5YStkK4bZ1BPkv
c2vmnRT+naNlDLXHKs0DpRAK+Mh+1u8A3gps7S5PxTB3Zy8b4qAdJLKp2GwuL0Ks
wl8DqUInmIA7i5qviV6c0w0ebInA8jnZaiIOc29ftCnlvIAz71Zrd3CpkDXBo+JK
7dgxxggAqEDVSv7rQOmBZZfN32wLSqcPMNd4cAJGFv5HsI+MK7rFPIJv0ZRria7Z
IEbu4OsasOdoZYYEoEbD5wOeWyi0zx/uANc6Lx5DVOn+KMN4GA1KDKGNxWBy1muH
+6KTxFszi46lQYYX73+hIY54nrJbyoG3/GbF96hfZcw7AwM3Tyacn2OwOiyUi1qh
uU6xgLVsq6aIpwrHf+o/eZXWyGTA1DysDn+Ly8oJs5q/VOsWJMafHxNr+XkxCp1x
lj89HeG4hRqDzNvQ/SmcwGoV1kCQDk6WtqRB+WA4q7m4pLoQ2rCJ5GsNZXRjxwbi
/qnEq5jAOhbE8CCUthQ/d9lqHxI0x/wTVEGNCAXHqV8YtkEggvEmZWUCP2M+gYT6
VGfepN26UmMd+ZawlVmeaWw9cUoBLOeg1hgTQ2c4J5tGaLq5y6SU86gDR8GZu8f7
c8A9C6aOQNHlxmEKMaOJ+8nDRm4Mt1CtgWP9ZKpkLfh7/PGCFV2wbk/0k5/RPFAP
4deiWj0RiyHF7PtABHBq/cxfuY8UC2x1mYCRhvR/q5Hq79YQPedlvQW/CKwlQAsf
TouLBH3CmCnJfJDjMg7PlJUGvz4uPTReUFe5jlwtsGMXCY0H4WzeBU88fMAgbTMl
OJNeEM423Pyo88U6Zhqf6xjzTQfGJFAM/kChheFXbN+htwjS8SISuhUyk7Q1NK0h
TBuOFA1iYtzcX3MRjSPYDHp7nWqrxWZQ4K7PiXDWE39aEITvq79FeKfoAGFfAdt8
VkhlRK6XoAqATffLWh30FcjjWX7x/+75+qJjCBxGX/IVDM0662/gcMQRmHEyk4xH
7S+QAF7bWQjt8OxeMRw2xwJICLUHGcC5vjT8y6NtDFL/gMXUollJUkwSrTJ2/UpX
QSuIClmC1wGLczQACnqkw7G7SJ7zWWaLBZWCmjOrZY79zEJVJBmT2kbMQXcV941M
75rwx3Js+5eRXAUn7x1JzlmgGkcFZ63h24iIzriZlSyprpVmynj6Tnhe13dDqBRU
SBHGL57oE2TS/6+TdpasgDSmC+k2G8lgEK6L+/fXgG2f0CG+UXWWDuZChl02vkwm
Ful9T2e8gLfvH8kwiDP/GGF+GRMf7hqnYgLhzuj7yxOX6bF05+lEM8ron3LyoF0w
qvgRdYp2SgSbluF7R1c+VHAtGorPqW3/oQbvZ+/B64EhFoaOcMswTPSiEgPdaXqQ
CCzpt9/LjdcQQuziO3F8ketWyNSUQuxPCrDsJYnoMfPIwFBNQ8N9LNbksNraYMIF
RsY8uPsvbpNGuXxDyAX2ovRER3733/JWME6Z8xvXc2H7dwO4fOvyA0ihztwKQRcU
6i1EYBkSTqGdC4UgIhRYZak6ZxR5cfjV15pU789OQSvizJHSScDrzkh1CuI0GF/Q
hUhhMrLHSviFNG3Ezld+dTpqD0+bEyL6BkKithu9Rrgfyo+ysM3h07Od+xAd56ru
V619szeERaE+cxZU16fc7Jym3T0o6astlU2WI60T/rKKQwPelRWrBDr2Gp0/wRgQ
tXgCvxFnVQOZHVFCphZU764nYbNkNV8vE/HlVr/DU03av/NgORX/c7DKdyuwJub5
W6BP73sc0ZXRH7qdn3zWNLDT31jmL6XW1g90uyevzZKno2RelTXKs8XN6hYxflOe
1Gbd7B/QH8kFzWsf9DY9owMTleokporNkvWMav+oybwtYaXoWBAMifJ+kPmVfziZ
cEDeyuqoZGMIKyNaRv3D+qfwemsIZW7FF9YLSYTIIscZAw7aVRn2EQ9x1HfnAkZz
kiQqu4NJNyb0O0OUYMk+vaZB6d4hmeA0prH5njyobMRvPcVFG0t9ZmPBPTI5oItd
fmCnLyKCMXVcdsf+W1gD8jzK02SaAWv+83GTV/B6Z6rUUl18gP0dNS4mzWzemdF9
QJrn03chxfJ0lf944E10rOy8NbxJtwYq0TlTLrwy97cRBLeW5Y+iehOzq3I/aR1m
UZ5Qqs1md3e4jtdZBzM2W3ln9oLs6YWNH4hNrPpwkPprpJwEHTKEdi8/bLR62SE/
olA6y9EUGIkXXuSF+uDCHv61zD68avDVhdVuJU1YHGGbhn/Tw7LktmlL3I7tXqv2
6I44l2Hu9iFCHdHynCyluDtww4p3xIo1eSVRcUpm5mSUiUUWuLuj148BzLSA/RK2
N0wgH+VO7h9L3UF35La4q9/s40yCm8ONEugyJyIn2uUiW/sPnoG3Fzub4XY2MgL2
LZN1dpULtuDSJJVRj/Qdn0R5/dZo9y5zdHyIX/La8GAsyHBzPx00WSZ6ZrGB6zjD
bUT43M7IyYlFIfwYm7qtR4cYbb/DqUDbEy75lnD7+Cqpwo1z0RfAleIr3rSXPtE1
IyU7P1fBJ+tRzgTGdgAkWHmwJFmza+zrLEyYQYfQjDCIazyOdyWifq7rUwh2reZt
EX+MQxIu1XAfSrCr7kc6rjT/pPrvDkvz6d62n3d5dEZE38sud5Yv7VFQm6BDbKTS
rlnNcB1a0zQUVCqK0CyKb17bq2Hkl3BmGmwzAQdJpSrMLC+9LdBD/VkWt2a/Jy82
cumU9WP5PBVyVKJpwMRLlVhSQ4F8AGI7J+jlPakok4MjYKcp42EIsiMoQjUBVHG+
N+uNdx1lX/yEjJx67DqC+DzZiiwY4Q2pAKOmV1SO678FrMKCVqL2Xh8PUIl9aw6j
vPj558P6M10WwwV2nGDvccm5lXXvdj07k+uXVeJ7kgPn6RPcpfg2YVhquB/1cc2h
Ojhy9BtyNcIHHS2hLOY2WXBe5lUSnatzRuTHd23aChODOc/w4oRuhpbi6N/djK8S
5iOugstbfK9e0FnDyzY9TxTW4eRfRCb9S5ldFGdOFfP8MnogNCX18GxMT2vmPnwT
pW1Jwl13AMTrljP/9SB9skpoZEkPxJjZy4j+Mc45ZOLrFo+wZ+Dtp1Jrp/WPqWJ7
d9nh6eCLzi40+9TMYXuIBvTOXAR9aHv6x6HCrLKdQpdgSM2OJigDMR8GvOzY9Sj4
McSznAlAzDFJSFKXmwzShP1TzSlonC/v1l36t15uuQC130IJlH+Lgg8YoQfuHhel
2abxidd+hEDbM2vlc5KO9Plqa0eV0P+D9JtBWmqIlrww314TDLiO13AZBiObBfVl
Cv6BuESGkxLwAJ7b6t1jc34ereBgU/MkzQBOvF73tLIukUb4sexHZwJsFCDz57cN
sL+8FKUoYcuQCSEaunGl4j9agtV8KzN1808SwYSRsGe9PjTXgRCMGPTlq+50jomh
DUtQ+yJbywkywvvYymvvMy1o2gu6iHYYvF2il6mSOekelWrE2fQWFw1SbNVYE0Fz
4AxZD59UnHbGGzN8YBV9VDBejzFREPj2qCP9ERfVKNgE8hu9JRU35Fmm9GFNVPzk
/ef9kwKZ690nF/QUL1EWKQYEtBrxMUnMChp7TYeBThTGgYy3CnTyuVvOj4FD39aT
wPzJGEZlTFk66ECRDQVnxlIL90aO/qlKKDOaK9Gg62Tljc5MkZjAOD2ueVP1YLPM
ws2pqUSd/NDKj4KbgphQy5sPHIYo5+L04AqKULoTQrbeZeMl1cq714VoF4xpq/kw
W/tumgq/hpJYuJn2mm3+tPM50dgKuDmrAlymNKG3UhounhWKQXZPyF/L1GjD4yrL
iSAklcP7vS02B+LqzIkAanX7kBzQ48v403QAN7s7BBxzMX8eEgwQ2DCFdz9MzSey
se4Mq1o73MKq8JgkSmkQ++2lwzN+yFlLHVzMxeLA4b/EwWVakaiSDwUgsourn2i9
HtArMurprarglBLhuOADumqbC2KkkSW7oMbPTOFYOG8b44ndF8FqcQ5VSdSeaSeu
3EPZWEwLrNMsriWKhKwCzLr+3CmqTukZuuEr3OTrd1Hp4lKZeuteFTDCEzbQQxC1
2V8sQGA+GqRoOdaih6fWgfqWgNSU3wDqOGFmF+XmS6t64srNtB0He85LDgAh+G8+
xlw26YgI9cO6JI7Wh0zDzH7TsA7xBMebmlNs6WW8wEbJJMidVNQLxxMBQ5PVQcHl
UhDammw/G3wsyKfQgiLnhCHiKe3ftu8BISMjTAWSq4eVMZ3nxg0JRiG7dOpZzjM+
n7ppcJu4xLzVrvylPZSbf2nDTXWJGgKrd+LX4+y2udfOoinC0dyUeIRovKID5twm
vjtAAZipvU5u4RX3dNdBKabsY8rtP+N84KeM32l9FPAaTzlUO8Gq1Z7tmONnTucX
zNzNbtmCwIe1Kda5QVP3v9p3s2tDCe0eI5ez8eLqEE62Azqro2qtY99/avS71Zdu
Ze8wFqb5DNR5pLLfuVDaEGKdne6bgEzEAzx50IAqWC9pLTBvIidJUVcD2Fug79WJ
NNu9bM4b3KxJ5Ll3CcHzx2LLsBQwQE1MZlL5YdPyEKKTY5vDo3IbnOBVDz+Zkig9
/UJS4aWkCvxs9bxF7gR/6Pb9FT9mUAgqNoPAsC7+Z/Nj5M5ekTHEGivb8aJQiYJM
8/mH3zcoTxurWyQgykRON4gZyptIHRN5cMwfwr7cQ0mPouIZnBRg3hPXiArlg/mz
YgGVsvTd+Hv/GYUMPVtWYgTn6eE+vISg7K+OS1++xMnwdubyIxHeUbOZi748syoO
ztw/eZ36Q32dEBvkfJopjjBiZ2+kVjlih6uJ1V63gTLZH5E/iyPm/BmSL0eBP9dm
Q6JhHZacRehetHcLFI76DdQq0myzd2ibTwAsDrleJWk9Bz76PgvF/kBhRPjjP/tg
fBBphyxI0fK/p790wMW/V/9uzOF5GBYyjMvpyomsRbDgJn9Abxy/epvwoMNl0Iqt
DbzIJYKly/NW1I7P8lRikESQ+7BhRFjjeLCucMXBG70oewZ1Qe15S8OIfUHspR3n
QRoA+qAdIk2zq1yvKRQIasULGaNoNDK77k7O/kubSW8e0wXezLOkxIn8oCj7rxH2
GyuVDjH88pdkIvJPaRzEYUWIKb2Ak9nD4BzVUPR35HReNbu7o/7NRGBE9QoVu050
8PkUyDy+TxA9ajwWvbhwWhnMJDP1EHk1x9WadfpDzv2RjvLD5/tuKJwtScAlCF3w
I1uwip/98VE7J9rHjL33WvaprfBep0n7OdYwks2k/ra2qnhKxoo9Av0vE4n/bCj9
Smifw5HThvMPHpTYagc+uPb2Vih+rFygukkNHjdcK2b4DeJ69raAGD+7bl/GcBiO
9ZemE7cD+M73pbaFovRYnsXMyLDgCg6Fnz4PONrVeEu/eigbHHK8Fs3JDTi6r5md
JqcFEgrJtqkL1x8oWkbqf8P90frjyi1z/hAuKoBhbUM5jMGtVSv5ZtrcPOtoaPXz
XXK2OOgqFmu1DcCRaRn7UfquXo+ZeDePUJEMoYPPJHnXVrGPoZpXAo3LV+NFMehF
wlOxxDbGR3/WXAoPrAKHB5lsw8NNPdUV33U6Jj9iOt7NJzBmk165J4RrRxeBV7Hp
LpicILCKyaz0YYjrq98rxquw/akXzhszSJ/b7IosqYujdjn2xOYb95+eIHlKzpE3
LFHc8d6QrXFi61UI5l5lodK7sPjFIhcDgjNIUdz6HgpzsHmjDr5ha+Ubmvrz9bMZ
d1TF122MAbIXfxDAJfx366DTvRVptCkuzFTlVB88fUlYClDMsXBHibeEAVzV78VR
FVwydy2gczhCKeRB12hUbCillMh9muBjfvEP1X0Kiejknx1ySSJj1JVq+BrFU1Xd
uVXKarGdHmH1vmtCx4RY1lE1xqvlE+/0dREoO7mVWROQ8JetWq0Nq/l14wGZExgP
qYO/xIzyTZcsQJUDU4i3Kgm1NMxYNvlv2/56dy45YeFmonOMQmrW+L5z51C8aeqh
rTQOM6TZcLdlLOIzkhIfzk4EiQLGbPoHhU2w39i9kF6YRILfZmIgZPjTHUnWraDK
pRvbWrO4KTsyNCd9JdZ7mElTGOltB28mffPednGtuaTm5fMRcpFT4k20SlLQHzn3
OzTXHa8kuELTARvt4nIXbgipy04D2fWleZcfxsHua2Im3qd8+MvGjkJA5HJ9La2V
t2n5pIJm/1a2NrK1bhbP4DDzOfuX8iysUFF/Aufsyx7LiAOUxZpKS7lkttMPikO4
1PbRac6hF/pCVOGI7RDiFPXxo5fqfdLJsltYx+1VXdW0/Ja7tEMplsU783kUebTR
6R1QSKwNSo3Mzjq5ZbW9og0WTVbr5wa5oT4iexmDlYPI6ApzsY0ZNQkZK0Hd7fFT
l8YvQ+12X10jq+iezzsYzNRQx+PQhesCCxEYdcchukYZb+Jh0DEOzwGw1eJDIjyu
GpG1LfmfCQ4FQZhzWT4lqjlyOxKzDzIo785LYQI6153wEQzSZfawy0wFYFtOpcl9
9rmfgmRaBCM3qdz4rxF+x/+eX7kEX9SfqPs3glGyaPPDCQI5Atz5Z3AZc3wmwapw
gwPgGwnqKm9EAqd1uUrKfpRlkqgGAtV3OFYMVzYtBqZ43QVWmpMFsitAEaBqkWFg
icBFc+pm6Io/5qtKbTiudQbl4FidvJ7ZTYzbsMtL6bm7nWMwFKG1kE6V0nZ/YQMO
GpZP7OjB7soHpTxE4WTmqPqIYZEy4x6P9ef6K3eMXSuF9kXw62CQPTqgOsqlPkJT
lsB5Gle+LMbL79bq1iaQKINxvrWuk59UpBCxG6y9FxYLYfFLs8HXZSV6RIJx8CWh
zxm8hHGSl9w4rfh6viHOqrpa2Vwk8LRI6mzyOa9JpGmIWDvEO8fcai0y7SiZ5pnN
Y5LVm6S49sfyc0VXXGCxT4nVBJFdC2/xm70sXCDWPxZa+kbh8mIYcdSN7i0CDA2o
kiMEB3absvBrLpJZ/md2ZfR2G8JZigr9e4nt4dPkyUafaHcVD1uQ4cJgYrkjCD3Q
AGeMFCkHgEoiM77ONocrvvLbthu2ceeBZAX6Ew62jNWV0XyyPZ2z7+6sje7Goth3
7QwpkgWkxG2HOdIQGg0uRrXJHqsV2P8xf9UUjnJewnjjrTnaDUFVs10BNlVEDwPK
t4069iVxnDPtgerR5rrzefALhcoa6bv372NJfkZjXmw+cjCOP9GceUdvbam+tEPF
iLo6TFHmiinv2iyUFTt5HC9JCB1mbT593yvprWcL7VlkkJNmJphMYmSH1gYQg6u6
WwRYuFi814wdNa+wrYljaQKOlqGQDOjTcAeYUqYtSNFeGquFyWeTVyxiazwCMEji
84RbSHoi0ajWwpyWgELFt4MoqLtl3Oee+dFhEut+zctETamHg/6uhV+nQOS8cgPH
c9tL4Eh8GwMzuwIpce8k7p9udvaSidzM1+gbJH6Lbz/J+XeJuJHTDZywCBCo3pEQ
5BYzToopGHqFoWV7HtL0z+rSyrqv/uniSAvUFqJfdTSi15KW2XqKeJygzddnQQoZ
PX2smJpwO74ze44jOEfzP93GxdxXsqtr1JPq6vumDMkHXsLJsU+zahPQPgi35Jlh
yZO9iR4+BiNy92wW0ZdCxCHjBQqTeWZRwxtImVYJKbwPH+OO2fpwFeZpTKP0O9Ob
B0d2OPhs4Oyrcq/gWC6OKiSv9D/uY3JN9CdjwlJiAeAu2zxz4XQ+RuY0vQga3R52
Q4OohGmSzK/ecdgWSOB5TOxKgP4KdRtZjs+DOWa+xN/q4kSKHQ0iWnJz6vrtP9Yl
FkCYbK8oYfRdoQX6k7v37FhmHsVLKultT0e2O4/N7oZBVLaJH0sEN24vNivkLyql
GiVKguez4h9D62zs/J7gp5EebQrqRdkbjU7sVtTf+VGw0Ih1whpkKhIqV0e7kykA
LPJbPkrb9jVaVdohU+ZUr01f9T4uKFDUO7lCmYjOolvZatVORJzxbEaH97gZO9cu
Eof+72xqNJ2DGe7OpeIfPvr9MFj1wvPjm9MzkzZvvWIxEZOU5+Y6HY5AQIk5a6Hh
xecx6X8LqEwCThDyKTVktLDrUNERneUqbE2vo2WI7oyd3zudbwFqPLmBojGJ1Qdw
l/UOKEa6RwvsLB6LAf7Zr9wxoIqZL9ouA333fJPAyY+w5iggVXP6aOTYD77OeucM
udNJ9WR3SvVJJfaxdC94QWKgTYuHgtrZyCWyzCICmGGRM35DGUZ1nMxnUyglgdQs
kb7RKWkAwVIwrlcqrICQ0EYuPb4imYhGTJzBr+SycrKlxvCWyRL9aUjSe+8myo0T
acwFSgYeKWgQ42A/EvBlRcNNxqHbJ/pdBXg6PVe5ogMAjItX2aJucfZP/+Bl1Db+
/71EOZF/fCxqdMK0YGmL3eu3ArjHntFEtY1nfLyBoSkhSm0NnVlBDxpYPSWNQKi/
1FtWiFgdndd0ODCnYsxV0q8BHONAiEaLZihyRw1f2xSbIu68cdbJpKJtGcRqdlhj
4a1Nu/6bgwIEC1OXlCr2XHdScDV8LZGtP1b5+gXOeMd01rdfEijTMi6FCbV2J6Kl
Qzc9U/UA5aIWkR3322uBh2y9U+8H/BbDU2ZlWh0ilaezL+2oBtvqWw000zIKYr4k
XX34I1dnFHwBJOazZ9PjCE04I93w6uqPxjM+fVXAChTigznhI8a8aBpW26KH0qpo
eA1TBMkqd9AQWxnZ+fQ+/rpjsrcsh6P1wCIXBa03RtkuDW12+Ww9wdGhJSdJWrKm
X6mqFj8ojGtbDFyJk8qQrJJSBb8fWnxWp9ojtjDFa4g0TOpn1mXsLlOZRhMRlvLH
AHJKx/xbuLmvHjm4lnzweQ0oTKvZGME+YIrHYApkMDboPddlHTID9Yb0aEQAX0ci
ERpAJZ3Soo/hLMytFNhR058rbRDc9tby+uoBmRvCYEUKaKQVnanKxmxR4xYnTEZb
SWhooJVOIkQkObLapRzP1RzwA7PONrFPEMKNqE4bzvsupXjBC7S/lxARerQ0WwtL
8CjvZ994GLqDj0tqW1awXdE4ycobpKNPklTGNrigxPoIeQfiea6jStOwQadd5TTx
nuzQkHk+zDNfDKhA8d6Zm3BZw6YEqGAacWC730s8jGDX5voKHHPzs+oQuR3+bh6K
xAUwR1Cg8pmeyOUFa6QjnTe9ziEmWB1RkeTj7atc0nJNSkvvou2tBJOLfyapOWMH
G8XS4XvyBtA3/uEhIJw4HhZsqjDjLmQavcLfkcWEve1VEsyLA8TePdgIpgL+cxsy
bQWz6fGYoIJyH3g1f4ATYiMEXGZAw4ZvTkuiF1GUdxUgiBQgs6tqRM8l+EyGxEVL
c877sw3X37jYaulz8eekNxCUD4v9dPxIuRXcDebftFY5hRLEDWen/9OM/hugx3hd
kjZ5A6h3oxtUlv4elrVH9I+E+kmGvYgfAYVrKycwBfqFN27Ki5U0gYjgOKVSWDcY
QYgHFFGu11pUTCaQdavpkT81G6OL3ZrG32zJvPsDUzobPUhAmZPiMM9yoQfuqsPy
jL7A3PLKNA99+Sa4G9QRv2xJ/siH11qb4FmL4A6y5dOWX9tEW6pPZiqBAHPXSNOn
iKHa4wPRCSjo4PO1JKOihgBj0SfqPCi/SaUcYmJCvVCm+KFZhpKXyfDY8KjhPHdE
GX4mY4vXLZ2xGGRTAe42is4t7Aiw2LvtJfWHVeVRpL6BS+usuuyTaQL9FK3AIcgr
owP+mPpzNaQKp6GTZUyDsvAbN1JDF2QefwAWEhHQg+ZYem+TE7O6uPGRsnjQnWLq
MJmxHqV4MZpUYTCWBfamc/btAyaZF7RCow67iLQnQdGm9Ct4tAa5DgLKvq0yRinV
PdQohWBAUtmbJrDVzxvJWvm1RGHRsHCk4LFO9cz50C7OsOKNgjDp9DnTc01scTNd
Lpywom0OfBzRGiKAZeBBVC18rWbx588MHQ3KZ7EAUepKKyzpGu2AhjXlybcRzd4t
8ylLgGmScBliJFSWD9LS6CDzkJdj8vesDO1gw/h99dM8WggG05rrpKRfZ8DcAWa2
1JgF8gc4pK6/u8S4iH+mpMcS5Jj8Ls+pVpoj0Y/GIVSk4vdFjAtubljpm5czir3m
sW3NDEuik2g10amr5726cg+Ovz8nCn92HkjOmlNOP47pHRVUpswi8SW0glDSwJxJ
vJY2y8mluOtTmvDRopbzpRrU0gZ7kJA+sKt+OVnX1W82hhEr9hgmu9Pldsp462SH
kKT/rN/Uk7zBTOz3z2lGxf+OZil/+buy65PiL5ZiQ6leE/Y1nhlREnjzcOGmJHdw
K0ngnoGiLiDE/2ADZy6lWDjwucghw5sbtNQOTEOhpmliiUWGNkb0RWPqeZ5FPL11
2D3lJXOD6rPqtMGiQ+3rOxw7pESEb8ciPC8yHR30QpY+Q9OeaBOgNc1YeAD0LDNP
ROzNvhZkbaxQIJwPT86witrXt7VCpx9DVqtC1/mLtIi8AWgUP1aM/6T6f9EI17CV
jJyY8s7fc754PSUCcllVZDDYRKAlhbz1E4/MJQ3P/zT3EAh/zEqxzx7X4drAnVpr
tYs231AWMKrM0XcP/6mDXynDXX2a3bijROrrwr9rjl46RMf5VDByxHI0qY9PQNqD
fBUaPKzJaz+gbyg9yz2WMhgJ55Bi1M6OehaK5cc6QHaKvQp7In/VT5M6jhFgcltM
WEU8GDn/c1YGsw/1PHY+GzyRT7NUNYBtkFTawrHTIgHjgvracgCjWkrQlIiU3eOT
WV15GD1gTmr8tQSqEX5QYB7dGzPoueFMkl3q0sqBOO95vL2y26ZD372b+AJ79+Kl
7wS7ay/8Y+PZaEKBqshI8meTcSZdtqWDd+yI+ZfYgnWnGFRTRaglDiEa9wgh1jcc
7Hny+b4aE9qsWmwcHfUT32SGzfJ3zwbD3ZXBx5ziZxAJi7Ml8ZmyS9GcKvrZl6FN
ygD55YRHPihHj1NqS7uhZc1cYExbdI/n5KAZ3oQXngZw/BFeb9br3/wHOqRtW7jP
CUvlALII0x3GlEgWNteB/2K7+uj+BZv23W5phyZOsGi6gIilafsk2bb1t8G75Wth
6nMtrtTcr0g7Amnu7pCsPwRNfGnPri/1b/LQkWDyqMhpeTMLcv09DQ/lMqNYP/3t
TQnsYenMbesJsjSilbb6gfdKavkYfT4Ie182jWbpPDshaRnYN4Xo+ilOK5Z0oLmQ
EkvAKFT4FkVKJsdQA02GPOnlVK3wgYIfFbj+xhIRi8Wau1/WMxtWurC6UgW1BEWp
Deo2mybSWwQFktneB8EiPqQ9tSz6MBfq0+Xdb6n/zJdNnzGk+IQk9NoSHp3qU2bf
UW2p9e2yNTJrMNf9UeSP3ayA+3wzoYpfdQUea3NDJ0SHe7dPRjui7nKFk2nsoL+f
YTYO0Lp9BmucaYzY78TWm+fzkjJ8fcrrTSyebZZqt4mxn4dZb6UxsFBE1DUMKw5V
Y1t/6B5BJ/sdhAtF04Jy8jldLRJWjaRzC3yGACz22UBdNgArrqGdnpURwnvaroHZ
Phua9+aCrm8k/fGGenviJ+NMXRxkv0B7or9zI1+TAf9yvhOeRvsFwf1H3MyVqc6N
1Meu4daghlvboc6V6hF+KMRfhhjdJ/YzwlevpycugvatG5LiO5piiU6bR2gy+QDi
4wEAn7DswXbYMgYb2pX+hl8G22XphtxbLh2kAkis8iYDkkOBDvL6sU3Y7PQ9/9sF
biAeF/XvMMCKGmhUeJT5wJxLjWg0KetSAuzOodU/TN8ju+cQPSO+s2Dj6b3Z/T2H
DNGIFaWNTkJAIdUN8ry6awuvmyjTi5pvb1WOYsa39ts6i9AkVkk6pZUh0uDGZnxY
Sx10K6bKlxZBbAbHAFqXcGXsvUPNlhykzWPV/YV8BOUqwVG56OVt/rabnwcb7sbK
YhwmREY+pL+Uc/zg9DUd89yOhM8AYKKOQMMW0UQDg4aLWiWvDBOgUGBn8ZWplDcF
C/EAoTfliof86+l2PsKcbJxtcPpycvBiKFv7qC98aNIvwCD/iTlm1ZlzDRq55LRE
0mvEzhcRRsBo9fXpj9PH9quR2Vw8Xm61i5vUPuuhOpAazzcpWAJIORBNJbBPE2aX
k25TcC8zRLNj8UgOIj7ahfaU72/wUa84zmVd1hegJJYYbg+3DAjmY1JPzamb4vvJ
ndreO3fmTSsLfdgYJ5elzEAMCdCe4w3JdKEfsuNaw0ktaje6fos5MMyJcVMl9BSj
/bOhYlS4auKC+5hh/+Fk7vqNpgNx0g+ue9XUl3skyYzCXBSdwLyvVQO0MfGPhkJW
v7j0qvuKdQOybgHwQpuex+Jy9A2OT/JnMiGdogX541tuf/Apm0iCdRNrJLyzCdOV
VN86n1SFEw3ZmPoGIYfyapUolKzGFKayhztldBbPLHsfAxRNkLl/f3QY42hUf4EM
v0JJe/Kf1H7AblyX/YyfDTXyvneIijDecJV6iTlyleMmzj8HxBcclo1nUDmZjxCd
5bOfwANCINmrYU8o+UPqEFtWt/SmfOXCQtXaqQhmftI68XktPmDHSx9xLZHA4v8w
IXt2VZ/S/AWA+/5V6YDSKNiLHb++C0AN6HiYDjMqDc6XOGNVvwOezricne2uSGIo
CHJ+9ETUAVYNGyLYcDkm+QWw0UbdkxZ0NlbxTvaPhTZ975yg4SYGHqE2uhkMAnL7
9k4i2ql4cqG6wLbcTN8+sl/11iTt2tCfa7aS58RTNxOYeEDRpOsKpuOGZ3aQkL+v
PT7Iga94V86qNSNDB0nUpDi2XJIBGvF36OIH1Mz5IXak86wavhoSYOVuhjcU86rx
FE9zUbBtzXO0r6AqpnWmd1PUjbpyPCXb5o14BrYUtvxRxRmd4/5dfw8QzX6VltEr
mQV+C869IYOTng3H7/au4DX2OHopmjiROn90nRTRwQpsbGxnxqsiU15apPv1qTyj
OoprtI/zlZJzd0IiYWZzkn6CRyCU8qcmNwShu4x4z2eyftf5LZxtJcrvuhLgjSfv
WDp2D+Wh2jP6zEd2QdfUObjICeauLrhzy42Mi/yhv8VGXHqPcNIWiwK5bPnD9sI4
0PFHUUgN+/ZKOr3z5uG7jO/qeBLVnmKB29D8AiDFHW1ogIVRZLj1y2ZZDeHUsITr
oXXRLSZos8/MaPTF37c/92g6K7qLB5/bYSUMIHSmjVYW86iEjNdv+yQQfdf/M2Tl
XU+qn4WF2JNzbJc225oPoE1qdcUUQgadzQ4EMV1ktUPD7srpBZxUxjgfjBvrU2CX
7I6HT8T9C/UNfJ80LZxaZT8vUQSwHMThBLKL9QDgSn9TiHc9dHbLZSAJ1s1ULVh3
HYKsxfXbZEyPfE0GUkou7yf3fM4yETvqB/gyPj1NJ9C2ZGCI1Dm6YyRxmOkuX3Mj
v1jwkUosd789yqm0HSRbIZ2MerfWg71xmoGSbkJoP70L8jI0btBNOjXJ+QaiRpB0
yHz/KCDGUJYfB+TTLAIUvXNViZq18dYukl8ERH2sH7ft89cnr5kO7ee/rpyM7yrb
s0+IiTbj0PHeTCKX69Fb5yMfAQJxZ5lS12RgUzz0S0YC2oaeoVFY8emV/Jj9N5uC
q4t/mm1Ot5GWExyMdiTZaosvwTD8ud+TpAT6WJaU/I9pQG1A91jS9wIzN46RIY6U
wEFDu3t2h0Kpur3ETR19ZvtG3F0qoQt7PkrHklk5IyAr97pVAw5mgf857f7+Y+oB
oIMYa0j3mOiYutYARzd9gtaybfcU06YeM+g3G9srGP3rgPtLNjoLxtlc4PdisLj0
hgky8p4Z2Nch27nB7iI6akxxcvUJiR81/yRj5F1RtmL+d29CUHSD2+evLX03eVek
mAqnPsEdplgIHrnfRDpkiRVDBsjlEX16GDR4Plps9oSzhOhhSWT1CWyFxJDHrZZL
e2BS5TXBhaTrd00eRyz8YEWJyF4w/bH9BWISCOWQlu158Kut8E5uHBv8TKE0sGo0
ElwZvloeibbK11GJmXlQRGmwu+WUibjZaYtZNV+5CTdvIzpwfbVFAKjmbdQ+aLH3
qu38UlQyJml6/3uhQ1xRljfAiX89W6Rb73i9xg8hNtLLeF8M96wzLHAJjxzmA9gp
lDYbzyXfpOC/Q9ejqjjxWO02O8L3oR1yX54nQsyGf3D+v3Sj/ZbEtYtKReTz89IA
xOqo4CtYyeXbQewIJmOezxyjf1BGMnRvJFrVHQTO7a3K+zsNeVqJVqhakIimeCjc
f4rWD/x66VQT5MkCdNlMrW2e6JRsZjA7vpR/ZLipz9C1G5ZedGf1KRlcT2h6FPVx
QRX05wJtOYfTMScp84XfbAPt+jfaV5wocWK5h0vEvzwCMve4T7u3Jaec7N24hU+e
w6kZIzcYrmUY8qaECksTRys4iDgb7GeHUX12LT7TFj1QZU3xEYauU3/twa/ZUktX
pSiRRz+zRrkDEm3A5mdycqfoe5Z2Fj2nABoDmH5aMJKcEj+xbg+In99zZVIT0hiB
3zzMBeYZaOjAixnCH+dFQQGSN0erC9qfoYBki/JMpY2kA9APU+EnK4lz5lcj9Bmg
TBWvpkZZ3msLFKiZYFe3CEsArV5iGEv0CTJ8bE/E0k4MB7sBg7NRH9e2yQWSmC4e
fBcgBAMmn9lBBeoEEQMoekf/ql5+7wmniAOVexrdR45xqxty8dFJOq/RaUvkhXQ/
AD0dyicOHsDtD30Znex4ar1NR+b2yvsG4BWnxsTemQIqABaNjvb2XtuKQc4SHhgi
V1Jao1Ve6NeSIqZDy5DLtbqJ4JNDP4M182lyYGmiGhkagMvwr8GhzZPc48EgXLsH
8MUGD+ajGkrBiTF+HgzCeyK/JpTlLcfBtk8w7Y56LYjRaeiRySvPGFjiD7xm3RbI
Qnk8CTbGMA0lGovDBCN185kLfEE51T0JICZs/naQbWfdNqMtzvBYBZTFpBmc7qqF
SADy1puvx/zEnGmBsFkxbnvwUMf7eiWLOYoLTYyFqSmLOMEl0OyHAKv/Dj6DsO5n
1OwJBDb+dVjC3Jpb8OnT05WrQ/yTncU9rH9EWg7+CJ9rt5KsJ2JLNpuXO+Dc63SO
dSzFUO9rrTXZlEXTQq5+7w0oNVwKUGhtWxPiRt4/3PqgSRqtpO+Qojd9XnMQKd1q
7P0miI6LJn95QRUnMbEnbjVck2anv6+sOFslLXws7Ue1EG2iuZEdnWaevZ6qLmAT
CBzD675kQlyIaMW188zJQZtB25mFEbv17fqgYluoCECEmMqwpaPs/jUtTnfEwzoW
XKug8LJk3fiHNZ6C1T2eovpHX15A465Zsq56mB3lMEx7H5AzEI8LHcce1TfVNUgq
MA5z8oUnkc7k/8rkpWIBgv3WwvdMKoZ033Qjs2BhmDOgNojU2xZ4Z+UHOVaf1c+N
xHA5Z+TFnwlSaPdiQuypgr3lLtwx0ig69vPPVcgymDObON8w5WG1SxjKrJdR0Vnm
V8efb38MX7Oz3l8VGE3vN7egvTVMv7/juNtsoi4B+XhpHitM2thZ7A5sGcBjBeh5
KN5gvwfrv/aQMjvQDrp9Y8qRLfWDrwIld4S6XIFrhkRP1zy70E/rjlxw+313MbkT
aXPa7MhMPDH+KjrZrd2mFvoyZBqJZa1Ahlbk8RkvMYty6vYPWhOyLkIasuHl7Jwy
r8spZXxcydbI+OIDs2TUWmg6V91LKVsrBpPMGPD/OUBf2XBkiBaN1vmsFZPPUwI/
fj/bm4UyuYE5yJqfzH+rrnL8lxIi+rWbakS7LEvcRwpWwJcXODdHFM6udWfcJ6Oa
fcw0kBaIAiiOQNmo9zVr0cGb1MRlcufE9OJBqg55qDQ6zeBBJpe1wI/sNbHYpu/z
rPL3iGEGKYK+LNrEcK7qfDT03+dIQjIpeZS6LtUDph90amL9OtNATsxgj6+aP3p3
lVmvMeaCzK56vDz3A5Di/czzaDqyEMp8Tuf73jPFNGvDlFYmOUF4qNtAKIZ/NaJ5
9AYnwv3ODhKrK9GDnycETculGteUJXwBfNKLeNPbuVxxli9TcT3MBI1jh69MTrCT
R7gEaU8MJYY8CTPl1MP2UYMNRYDJMyeoYyTdpP2EhyFu/hJgK5lFDjaNWIAGGCnA
jfqFU13ebX0CMzw1yQ2qLwec5zLnxN8Ne7LZRidRmp/KOULE8csfVuEYCV/CYYQs
qJzLbemCr6Xh2z5wr2sbql2JUB7xqij7LG4Zkeck649SgEk5h0Oiuns0WL0rpPbi
OG3qJH76X1EMmbtdR7LjxW1io2eDRUGa20yLj0nYfgqJa4JIxBtOUCtAtosQ/Hjo
6/31FMpDYnPxzvw6YeLrYHk3N38DuMUtQU/KUhNWsXHM2kzY2lNtS2s7PCwdGApl
w3FWAq85QgoVkSO2JXutFL0bczb5hw7do5AilGZak74cx5rXHNpjw5X5kkRHJECZ
HHS7qD5N1zn39drzDVLQU3++cdhSkZH/L6BpVl6zbDJKjUT+DZqUZjrAUOadeFdE
hcXsnpLx27/rPwpLIN7fS0JOvKGQWi+tMTRkVzPksgEP71hwxXPuu5DyFoLMsCAD
b2NLyT4ou7ku750vgei/kq70Az6hJLSktAno3hlSeaA720+fnEmUNIOPH79l5cUK
kjpGTFl33/J27ed3B72K9tY+uwYzImpC5fjRwpAqP33StUIL9a77dqUozeiLaLk5
1+wlflpMBdIombBLYawDCEdeMj0f/NqnI+OpUy5jDxuPf6y5sn0QE55o2r+W1dAD
laNHfSMvhPCv5dSdteWp11cNWgb+hN34NFMtM7bC3tB57Ae8RjPCFtSAStuPO4rK
Oa/lSNSvRzprta/y1l+cUouEnkY4OV4hHX+D6zqwssenljvZpXbR1BCqVUa4jjgu
T2RGDGKiqqF7gtNln7yHo0MdJBNtgYy7xrMDngt479s33knuDA5wLxExPNSlWo3+
bDGgqLbqeWGDoggw2Gmy/RgImWrX8lE5xPRmCKthp7mzljjhmHE0Wq2UOrQEYtlI
4MPZ8h0HYpWu8LJlnybH56uzkeCQFan0t3zV+MQtJ0R9Bq+ciGPHUODyXC75sq6t
6fETksx+xtJEEkhRo9CR2hDXsIFDENEXDKuk1S1bA9dL5xSdg+wpBr795C2eFB6U
Ygcrt/RLOwE5fy17Njx07R9qY7PnVKwqSXMM53Bq699nmbx6nnB/jyxZuseiin9P
LJ9v6BTwGAcuVPubeFIKsnwTD+otPDlPWRDcPAQ7SBuRAQw1dT9RIqEIV0mCdOYN
AkVoTmo3B2aqVAgP3EZZL4aM3PLqDX+frPbtrsQ117sUXwFN2RO26q9Bb805kupp
D3rCsGX436BLw2gPPN40v6vU6RG/DtzSg0ko9ychEnlrfDUXiaYvrHQLR186FwF2
9zGFePHGUWYUL4DylAipcWiUBqNQlheBU0RyQwN0p0C0bp6/bdsBOEC+TcL450IW
5A75/xP3HANwc+5b8F8m1oJMkXSF9ZmOyR0zYGA8uk499SRptOFHB2CdOWszBk85
nJlpchWEbk/ic6/dQorV4FC1a4BOPjE7CWawIOrquBIpVWPR419TUN3ejzOEivFJ
dxg2Dw/VPgE3t1X0MXNPralUA11+IWKWdu/lDuzLcK0ADl4x4GgYMlo5pMmsP+Wn
1VEgrJ2bXA1WTZc7If8NpdGzoAu3gVTF7aTA//TOhTtb/yASiyHeWvO9ZljM8Ykc
uXXYYYB/jk0daQPlt7YWlqnnTNKTysIT7B3GFcisvcT2kUl8EDnxtG/1dhT/zUwg
PfqDUaxHknEextyjeRGEF2tYpIXG9LGL6kleuf+vjO75UDfzqXV8lp/yjxzJEIMD
piBKgVqAd0gaANVBKSPbTXzVTIL/1ZCmCt4IIhq4NS8SFFy5iqDZZc9n4xSKxnFj
Hx32Qa7Veng9d3+kJb2LEXmTwbmR/cIlAC8fVC6PSM5QqsijMIuFMexoC4AKcx4U
gTMIUqRvPWw4qPbWM73+MYdfX/v1+FJom0jTTSXQjrQ5HVuI7DTYdY74YJqlnMV4
YQUoUDxDn/8MdVNpJnaVssDzSWGYzFkD5TIWteuN5eLyrVvUDPWDo8VPKTzP+EGp
tQXYwQJ//RWy/Dbjg6sOJeDsVC3rGwTofnM/wCE4/9yvvNlGZi1x+AVd9MyodRU9
0GS6c7oKdNYbHqYcgiD5IiaNrvgr8OskN9YsVpGmxlIEHC50eIwK2cwhIYJSeVjI
9dfYmKRDt3xBxt1Y5SKBIHB4x1edxs8LRclyg33U4JriDWREW5IzemfQoUKcNRhj
TyaUiXYgKnA/gOIjQrnK61wm1KDxYwp6JMLZ8FgFYhYzj5qIXmIH2IuB5r0r68eB
WPAY0EdSIBADvUQDMXzpDxLJreWblgorggs3Wp72ZZVp5F5wi+R5TlVFlcJcZ55S
Mun+xCWKaAiuZ2DfpwcuIHzFTUPCjPg+XVeqOV1/3MXeS1dbKvP3vDBmVBixDTgC
/AWvbNG/kKlD9eFYYu2CxPPhZg+Ijph4CGEMqP4sYD5KDT/sNOFgiYJtBSsBcvns
SODwXdl6UF/6iuarwUU2+B6u1UJKOXs+wYF55ZWWLnLcOh3m2Oau6KXFbeu/9xo1
PMifhaAAolYWMsDTr+0vA/P/i0QP9abrV6I+lTaiVB4aAxpU1tIOkT8E71uR6+hy
rGiYV+6rXm4MZS5qR2daCBTjmkQWpbFbVyoypDGpc8RjE3lzZLZX2Ah1Odn1/Ogn
9obcKwR7W1+NCIVO8wrb2dV+6bpeiXDYkghGNjjjkX2w0Y4dmI0c2lDVViiungrB
8stcjKFgE9PRY4TBPMux4Q1op0NSkKex6Xtp5uLAdrAQP0klvNz5Jc8Evs5kbPvK
9yTVEhDjgHFTonhWo/hWPNvMjX7u2jniAU7zPVE3Mh+YvWQIiK6pfmGVZE5UhMVO
aROmNY9m7Nkg4P+UL6EKugGi1U0Lwo8lHI1+/4INhTU9XjxlaYcr0dNbPYvObseA
KwmHspx0n98isL7s7VAltj3YMpbvWq/9VI6JUo3sVtsN4KCXUOLTJJc9T8eQimX+
nSkKeMZZ+bqyPShVnRnUqf4Yfet8MIwQT6/9oA4GwwXIyoLU7QOt+/GEKaQuI/Vu
cR5ANIBHSaVknZ3buk9dthLMLO1A3Ku/s2VELV/Xpu9kWuWf/8+jaogKpWuTHM4W
nw/NuLbCoJuKFAEPua74HIsx6hLcuajAHUL6NNBESQqjV9839LNUM03b+WnALF5s
wydGy112Z7RWcYpS2Hpx3cdjL8unRZdCAqWUf64PjkxL+W0OTl2bVmw08wGG2qjD
QIwue3RRKuJIUHsuiIDahpj2Nhd931OIaY8FdlAkMIGap1iqpl6fuZpXehvdaSwB
Ju1w73aTG/fta5f3z/gWhBICuwdNuB6uXZZ6lyTsLsY7y+oTqFbCYvpV4FWivWPV
MtWc0oD1jcKwXWpe3e16KSk01EgiEzqu6ZOkxYWMzcmlkYwQo1YypdLKX94Rwhlr
MgoAKt87md66MMz9QHYTRcWHECW++qha2gquSULmog4TZM08103kVG7HxRcmbo2e
XAFLWL+9cwBPcn3Ss/Cza3zFEmqmTwfZZkVduin5unKdhFRYLPXbhysLPZpYWz8k
MbCoPDPzTVtIbqi0mUXHzCBmk0CBH0+LjWhKOu41oRgjiBwdlp72mugbEP/jsRXn
dgV4cLWXwKLydhs8XmrlMCXCezveDqrFlRwvu1mmy7rXKziLuF7+B5imuRatjefM
2yDhaC9VehqP9zZxIqa+SBYd1EEn2l8xOZ/BrOZKTkmLZfqrxYrV+BJi2p02muqQ
ZSdBPDbPzH5DW5Z7Xv+CS6WRKJJuTQFTMZBVa5wzab32hDjRj3exMRTLnQLPXUM4
RjYHKkQA0S0uchzMEy3jwNKA/geuX8rLf7rTCZSQsXAbqgo2Zid9KyeONxyseZeQ
ndvy+rpiOmzD/kBIv1EAQ6tVIw58NvgkQnk17fOQupqwqqL4l4jkAm6K2DZqfUYf
dNGdvvbIIZNeIuJ65SByO2geChuF62vw6R2BP7545HLcyMEHLPqPtXFZmgZCWAOB
KBs4jqlh2VcHR4oIZpe5mvo/5exf2zLPpe8kNHvd4vBspsc6b1NUPsgmZN5CpFtW
EtjSP+SSop1+jZ6yL6N/JUnkWlv51Pj05J5svIVWncFKT7yz1rbEJLxk9EkmGQln
hJjZfNRnLZHPyuRThNme7Z3o/qfIfcSjQYLc8VM+NWQl+7ZduvEr+GacHkRKvQoi
gV4BIC7emXc77g4yRM9MBD0Ez6f7/95uV4rv9nALvUt/w608kZMu0XNq2B0uYwoK
YjPgptWXw2sNTeECKRkc/Mwxf3ZsGWRdIlNAUE+yQNxEhewLPXnOcsk10w8u3sHN
ZT6UXMPPQh6ft1UzziwtlNeOl6SHsZ7vYpI1zlj/Q745LTrfWxFFP5QnrjyKX/7w
EYdW5kPcVB5Cwrn4pw3W56Ia/xfH0SQ6j2IWY+yDG4L5l8I2dd9y0sHcJ1T2wFmz
hZ/on8XEDKyX29PElOfikczrctcowgEBQOADizriHPThfylV1GKTvDWS1AxVG+06
rX536KKNTiIuIAr4ElyMysqke8DbDdx0Hq5wPDIVtyrbu9XzIAFeKhqxgvIjhBcA
ipeaXnXalQwgOfX4KEFadFOTESrRm8nDreyw8vIY+CRlRKKYM+wgLXD7zjojUthb
3M6Lyoso2uNapWTLNI2LkIFpXwWXT5FPBkQuTxNuVLhZKwyBXbCQpourNQ1MnASX
Gra6aXt8B+WbRlihUwR158Utwwt2v166s5FvtAv+Nkko+0GxcU4BX/AZ0KUZxfLY
q6ZlN3jX3fMPQttTnUV0Wye7aS/kJEqk8CBywcuI95Ee6KH8Vsk1ZZoczCf8dUGa
Qfn26s/p8Dzlz0oUJNRl4WAZdFU3C1FnFnsTDcA8N3jjf9cY4RvHcHSpcNA0HQaT
kQ/CY6+xfpCqYkH/7TaNdh6fQge3QJQWLlOQzZU9pkEo5Dm7Fi4Qrf/qfdPDZRJx
AE6Ar+opj3e4+xFXy1+4yjx+0tHEscrT6VdEc7L5U/V/1Rm1HngA2U8xf7OFBkks
R0HDV6EOd/I4ZszVdjIOHWYK2UiPfuyk6LGM/YdAQPHH9D6TnqHtB9DR8C6VFTZj
eOz0vNyNxvlABfYH9dEj8S7QeYjjR7ShJmGl/YIjsE6MvYr3/jCUfrE4ddokZhzw
uXuyS4KolDAttVfOjv03d1F6iuJS5GDs8yds4PrCmlhdDOjpt+IeFzycFnxHKpDl
DOEHxLEk8AKQKQeNZFFL6U2PLIvzGDBoYIPXI7xnSTICXag351aX2DM4Q8zVjaWj
0ZT7hhlfkH2E9Y6l7XZ5eHN3+Lp5tgEtrl+tJDVDXU2S6OBSoA3XM3cHykBGHclC
8KHwz4UHP+Cx6VehIDsr4b9F61+d7x9JjrYeVbY/dBVUXZfqMmDK/lKWM1DR++FJ
M24sgZvbpcq/a9+YStWzI9f3Z84UEDpVxmwHx8NqaUpAMykRpcdH/E7r+82Ex2Qu
YT7brFRzErNFLOkZ7lzRRbQRlU3TmOF+s/44HrsUUQioRE3+jG0Ob55s4CdiRCCJ
pYWNAAU6zUlaPfwZq7UcSIdCVwtjwKPnTAkXbd0U70Iwo7X8cJNzCxlm0mb9Pyqn
sOmJ8sPoH6KtnQ7/UWBpnQJVlXM99aAxuU6/HsVyKC5NBm4iZE34JN8KYEur/jt6
fQ3QRWp+tMHh7+NorqhtF633RC1en9PziiJ2XwxkvHQjEEdl7kDNP52kz6s4ZGy7
d/5b2sH7CMfJ5jAFFrsTaTmEf2ce3Xi5ll3TTTOTzdjCSf2sQfukS9tYbo07S+ch
8eFZrVhOPdxKYBh3UHCPuPJF0K//HmC+siSRprModkQjHBTReHEj40dD0Q3IsMNz
yaRBldJY/YCo59xAaurzvU/rh6tsSdxbkD5/2dUE5AFfndVSbrhmO4fBM8bfNxlr
G3oPif8uUhrn/Xmu7bTDNIunKa5Uxrc1BRNVHpb5Rx2f8WloyaME9gV9yzpJtzP8
jq6YlIHNuaJ9glDkHXjxfCqdmFF+itd8U51AlzWIVqGOu4ehwGa76bxZLQ8VtOId
iFW9nOX3RR6q7BVI8KS4lh5Io5arJdNw+mGxNQc9YnEJFjxkXIsUWqA7ciUeYDra
gbvukCUfDlSB0kTdRk5OIhe/XL61sEsJGHSfvJOP4+zMyMr91976hOFkPSrQtuI5
HHFxt5/sW+53ypYRNKtH0VGIyj3an7WKhdsQS2ZbufAGILHPndqXNukmTEc/EkEO
s6NFUOOTO/GauYyib0QfEC3akcSkhSCyBODkjrkZCGwBcDg3VORzvj0dPlsbAk0V
Y1J+kfDJh794sDsaTG6zWXY/1T5qAq4uvIRE0otIz3Kpd67H4pNPVeQuWRO5tnZi
lyg+N7BRy/wTsVQtEVgVHGvrhnQzpNj15phWJMBi26e4o5YHchdayiETJ7KigctC
/1bOg+3iHsTXavS/WWJew4pSpR2bmAEwDd3VacQVFHfWRNumaTHXZwiMjeHLnHDW
Vl9DnDzYHMA4UsusD1SAA3FBqGFaZ0LIqdyp7Vu8PI+OqqmjwavdBP3s321vJ5rh
+6XMrfKjzNWd+5inXfToCR3k/ucrLYkHnCMLh7c6Z3w/toU51XrFdayeftNB730o
f3zRCzZdAv4/TiAly/3VnaNxRHo7O4sP5i46edLtTvVgv9rfN8bHhgtXR4AdJ2Ls
5dQrTDeyAizqi6uRrgxe3ZmLIrnaShqBJL5azSFYvdIbo7t+vALOsM2ZEwLTMGM9
Tn6xVd5YKpaqxSWEQLv39O/QC04LHx6XOki87cRJNq9LY3QTAnIvnjvlQ72L3xNf
IppW6eSUHkgEWfH65+73py6ejxJw5ti2JEPwQK12arDWs9x41/mrVfMMYmBskvSi
hYl/jpC/HzXjK5J81IlJ5BAtVGH2WwFFDEcczZ7rWdXaZjYn1OlnBYvtBIVEEeA4
GinFqxc+y7xuSe+VtXB17StI2+OJM8sImKw7OL9VlFNWGCHkmjg3g5BhirkD+GxU
O4wsJjEX1ZpT8O/FLS492CL3xhsFVuqsZEAoSneMClT/Ts3iWV1qDgUO+xSzoz0t
eTiyGcpoKwD+xdTUP2NQv7klDKk0veObD5G7AuKXRSU4YdwXUIGYd6WC8bYRJiYK
qyMux/cWmUIxoWuPjZji+oZeHGHk1NPiXfj6vPzSnKY39pYpN11juZFigbmmS5ak
rG6BE1ZgD7kc34497ca/Oi+8g/KqmfrIcdwO+eRzRAHuou0Awe8oyBf+OeccbGKV
QoKqn38l3AfnOcA96+SeLWXTZ4/Qo1IOQksKpbtV0HeGcp/gLB4RebHJ/j8F3bTQ
tNuvGpj47gfbyGQCSb3K7rAyZUNTqAtKZjgckCJHILYw9s3NIBnfQXPAWq9gUQ4e
dNp2TpbifH4iDK58BHE9JZLtOosW8GyYitwV0pYycPlR/73JQ6YT0Guq7mWZpeFs
kYnpcfiQmP/P8PIdqcoD+bU4a3frm/OeNHi8oOySNvKh1n/3X7nZCAxl5bY1QWOG
DLfQGjguSKWI3dn2VAIcqVzP37VVwoO+nQ63TZuQGDHZgGUTIFmLGgeaTaU7xLd2
1ZTJmrjarEfKt23avpPpgfCGePiSXjLuqK0czKDj7d+OzFwBSRUUv/8ROIzPAQow
LdipwFNpFS42mE1RGmeMWlsEOhNHHm1jP4wClKcmnbPs/diRrS7h7TjXcYyT4SEc
Q5ZdxFTyRizsD2l8Rw4vf1l+Uf6h9ANibsR2eJRJoqyzdSGwvZnOCKROO+5QYwHj
WGABjtZpVSO3Jrn0PUpSYe1Q3a7ku5aFSLAsp4yWNnzl3exb26h5eernjNdX4WCV
oFj7ikf/Mg7c6QMKI/HgZ3km4XA1Dsbyeqpp4rPG9cF7UYS90zlKoH71RDvzo6cC
62z0unePBOKxx+WqmRoKQ5CfzV2ytY/Rq9Dgpa9yEnp2tbUOkbguX+8nN3mS2TW5
0MTbVke4rgfbDbNYEwe2/7dF3IS5LShCK1yNbiCWe4W8mPfGQpKcUPlW9OIlDiKF
fE9oWFSM+wZxcegXDTwAa6exMIDeZC1XZdkSQm1MQM/5m2j377Kx48mPLhtMEXNi
snH9RuUkIHBhLuKzybxPNGCQNu2r93od6kTir4GKDqykHtlcVDvmkWia79nmyXE8
t/OndnpAVP+QMRPDFOjFoUJ7nelzE/8zXBC684gEB1tGoo5vVubs21XZB1M8zHhx
1TyzGVnyEivmR8PZkAQx/Bg+zU8drBfKCXexzVtVwMzOmCgcNWtUiz5Wx443lbSP
zBQ+VK+lt+a1lwyG8bQwpn5x0t39oAVMqjuwHNVJT+S7YO/+X3w12zl2d/7nqVKu
10NHCUCM7qnPLdeQy1ez4213lOCLro65Gv0XI2dseDYMbP3G7LRJ4kAr3/PbXE0O
w/0VRcQ3JRuC5B/I1BF3KXgFOoQgTpB8lROE9NlPNTJDB1eNjOIdDvfPowjWl32F
aVYbGdFrVg4wlbDkWgBD+vV7o2i46pesL6oprWB/CSHCaWw/5zQ8XQiv2Pw8PIEX
D6IA0bZRj1dPH39k/+TrM45iv4foyGTF+FByC5CFKKMREjVFSS2SPx2gak1SFk/P
KLINcFtmt4yyf0z22RfCFzJGkRaO0IlSbW4ZoCBWagpoDfXVhIWsYONj/A/L8dNo
rfMz7mkGhkNouCoAHyOlGsTCpsWfeqJNbfTcmaCVHXp+tT/6tOS9NTedgXEu1ycD
qKCgASrhkTWqudoa9uMwgTe9nOcK1+vPFWIaY6lCvoYhPXLZlJoMQlnPP9ZyKf+1
Cu1lMUafVlrcTrlI3FUikJcJYnrhke/xbbfvZg5/HcH2xJgnnFY0bdq9wTywwhk2
Vl0gagfdbzK83clEvlzWfmFlzwVlrEqyJkrgmnLn3jg0W5lm+bCJ8lEIiEIF+6kA
t3Li8N97oYmDzEKK63J3dxgd6OQ5zUQ57INRBHFBkFrNyI9yV0F/IlTv71qrwWVp
kHL9y3tKyjYEqeNBwwCIYMUiD6zrxkauISZpqub5cMW5cC4UuoeI6vfLPvBIst7u
1QRhmImd+Fuk+clr8NieMjK5zTD7STKcVNhkGtRSEoV3v8NXuhnjdDVh5g6SMb7F
4Kwirh4qaWDJjZjF0zUmM+dcNsTi7tmc6sZIX4LloIO7gHSz4gjj9tbH7lvmNeLP
TU2Htn7mq52mLCr9ex+VtkRUrooxZ0BQPIUrdOu1nZGYlupi2QykMZKgb9/qkEPb
qHLN4ZUPOUOxZmKb6D578dsVwNUKU82BrM1S/kaYLEWukb7lqvK3AqeoliDBYqMr
630EhvBe0MlmCAsnoHqMbYn7a9m176hdLN6TiwNC4Va/n+QGhZjH9CDA11Lr9az7
VQClCdS6FdutxoJCPZWAY8Hi7uS23SJ8W4xrvPFzodgzy5NF0jAOByPqUp9z86E2
N77CTHYEPEHlfFP3b4cclBDZ1TxjLiHLnXD1dqI9l0hAzF69/UOXQydAVcWr9e3e
uo8J5geSML+DjW8TKGPhmWaHd34mKjeEd5YTRod5mcvcdwGWuzdRLhxV5ex00ocY
bGpqz7JnMiJoGs9nnR4EPTEgyxJtwZFrbrYlQK+c9PLG314cyHFXw+BY7hfZoG5u
gpdpoIuoOUcEqgvYmubFrKLqp3/zbzTRzTeLpXaAPOqFIyi6L1sYEg+J00XQo51R
iqG5/1KmmO1iNlgguK4slUS2Ww/9VtPnPH1LCZXmN+HjFHGUsVwSTzZQoxz4Gf3F
4WRF5I+6o2foJIHO/K0bm1puQkS0KwksdEl7EfTyLzUYZYJiHhU3+nsa5GA0YRAA
g/SXikt7Xsk2YYuoAaC+PVR3Lk4gl0WfjADyz+DsYFqRtEqXeW4xvMJS2qinf8Ql
n6Ym+fWGdS0h079AAkfVrf2dLCuQLnOP8WMpTCqAvUeLapZ35qBVUWIsZmeYKkQf
u60fY6RPijRb+rU+B6HSQ7LsTKk2nf+tKcMr6FjxDfehif1VTu8EMfYOFPjTiyzD
I4yKtj2wRsOS+FhSq40lHUW1LVcd1o2Cr/jp/13Ie4cyVZ8zdDuCNh46BdadSmxU
j3fyEbU8JDFYfSeorxYSN0bYt1HtZtswmaEKgrwVYNaGVuIJvINAb2bK3RSoBXtZ
EJ8vHWxP7dDGuLuqkkkzPShgKCUNuwMBnC6ObbNtqGCa0+qy+Lo8FCxpzo6gBvGq
Omq0LJNgvN2h+OBK5Snj3Fav+q1aE15ui1xR9SI7aBqIzeEKTnB5vaTxrlSS6w5d
0PQzmYlfQ4VAL1rFdWMJqekYyaJZptJJOCqlUa8x2LFgGQIKErHqzXaLx4HeOWVU
dmr2XIfCFquhDVSgt5lvr4APDuueAKCDrBWodoKsSPu174DssPqK8YyDXemjUfns
N3k+/8Wgu7+7nHrC0hoG6GC3clYYFtHkDpJ8KyEsSQ42NoMGGzDKECMbNyBCCOyO
B8t/eWny6DUI597DAYHNvHS+M0kl8KGRWvxoYMuEDd8eTheBmsTOZWUdjA3Zillb
ArzrknYRim7plvPsAJNmQ6RUtmvzqDuLnsrX4PcXuRUiVxMfEELu4R8sZvcvElz+
Qqumy6n3rq1y0KuigKoFAFlBOp5wCi/9xlVYOqENqiZeyGOSZLtFJ/B8/0T6obdt
QiLqThpyDWgfC6eANQhb/1EfIupa9qaKykKTFu2IaZy0AD9eVYaWiJMg4gJuca4O
m+5dBVrFmsXj7/xHjEJLRGKNzjJAA7Xlm/FH3i/VtkayeSp16fitmECdYHHm/M2n
25FoQuh1+YgUgtZihnoQeRCtCjQNzIXaMLECfTSdQvDKwO7BiDvD+VcphX8+FssM
Vn4Gyf/miORPribD9YtpksPrDoU0X9ebO7Ox78GOgZEFcrjGgIUdfdZF6uKI5xf1
op8CjTL1jz0iykvvO+GsxpdT8joKANLnCqBvrgoeKnw1wL/zcPkPSFKU7VRxcbMe
SgKyZ38RGtUAhGE4VEwlJU5/ljZweKqss82fSW6Bjq/EDSWXV/WasUaWm6yqiOGe
sGyoZvXZuH/3Co8u1PIDSpq0HWx/gJZEnK99TWcJwm5rj2iCIOYhUiSKIPBe8DB5
yDRiZi+DSR38iK886pfSmjHS7VTXt4S/M8kY6k8CRTAl8eOFJzsBMdDF8z6UU0dg
xk9NeozbHhf4EBNdQY5Wh9bHt6gLI4wMDy9FXwPRbjM596rBnl3ks3DMz/pbWClM
q/CGC5aOA7zLJ7VJxs3t9tKKmC6vDsc6CUphNmzDE7ma0iDv0PTL2fA+mCwyBuUs
p5eAfTigjvHifGtCQr9yzfL7EEq46MzyGa8wgCa21oKZpKDoGa/uDeDYpxUcLhYw
cOd5DZ65AukikrXQQ0nG4cdG9wxaL8WFkz3WBLUVh9bdaxd+0evcURweTuy7T9x/
5tKN9i9+ArnIr0hkwH4fipNnCWXItz+hiV/K7f340RIzxr6Hcf7FEL9mFfPoncio
46IdjEMv0HA44cwCDz5JMMHWlqWbX2asRJQ2zSMmSBNzfLEvG/gSyengGI27FaRY
OggXCZVzvlv+zBLRDOJ8nFNZAEIGBIHsKJCryx/F/50227w1rGBusdwC5X6GF4/p
nn0o012ONYBrkpDYyGzpHS/Rg1vtK5a/dtOm6WmSrSBq8ctXdn0qVQRD7d6YYvok
O6B+yANOTc3RvxcQIc1zim+9YNNEW8BeaB8DsuPL6JHDHUKUhLXZgih87RY69IcL
//9tPrFUn6euJVfaz87PD+WabTD9kEzyhLbgo6EtO/O1q4lg2kmtlTsAjv3DjFOA
9Up+yd27LX6w5FnW1C9iMZFJtbbrkfBkOI06HW7+gvpE6w9T71EhJRQKzxHIVUj2
0pFOb8wVSEuhUFcdwFR5eFN1sMlWyTrlpcMvcvJMtO/2isUfcDna7h8sVwW/5vM7
bzADYSZnoMqjFBJcoOheL8DMwW9jwBShm9gES1eVYro79mLcF7Dhd4myF4poFGXj
lr7XnlE3OMFJJQbZvYPlrBTqFWFQQLgS4LBmp0DA43STxkzD5iBbiqXFw0tJlpBi
yLtuziaqxgXEflchkY2L15zwAKhDl67OcDDqi5mrXd5phqs2V3h6dZy6jYjVfIS9
YSwxxNi+JEm6DkMWfn01g5YpdfFqZoJQ1BS0kHQLCuaJdYAawRzTO4oR72gGe+YZ
1BSV64H5I46m2tju1L2qiT5Vd3tB1w8cB4/rS67MUtaxaPa1dATui95oxQB5CiOL
DFa3p0xSRGOmPqdHCd4PD9W/8s5EQElWKPXCYuyyjDZ+O4rmml6mPQaKOhpgQrtQ
EyURFyIx/XYesphE/ZZBklBXTdQbb4EPwGuqsSV8akN0l2uNPuiuNxDRn7NL4yeb
80zTPddS0P+ICmM3cpxrOrf4FoT04VXl7AK9yGEi7pwyCVyHwFlJwwDwXE7h0Fi/
s1tseKnvw52EqrzEWFMQQFUqYo4aEjw/nk9WwxwvjxYDVxFKZ88sPJjgubeEGDSm
+kdfwDiL7hUA9Urt/6tgPIGgcBScONQ0R/4goXe3KTTDaN0c6UzFeIIXT0007rK5
Sf9b8eyc3fUXeL4Ah3UTGZkOe8ranxf1JhyW9v9h6p7eiR9xaCQd6GbWxP+/43/d
cmJyg+QBzIT1oALYbGpH4LRcXLzoU/fVfcMl65wOCC8dIpsVZdi8vphU9YG/AFJm
mSrkRmTNJiMO67mhV/4Avh79Kzq8iJDUGUz9euVD+3DG1RxTKmAAGcNxVxlMuQZm
T1FY2NCxVCYtX3extj2+/E9iwz1qq6zMyR4A5PoJU9eCDf+J7D7jPFMsIr9iU3iA
b1RMn3/tcIaktSTTMRawc34iraZu0TS1InvTk89TsZjzhz9etPe1djZ93grHHpuj
vkOr9FUFOUUgeRdG1athCOgRRFvuekne4KD0bmNXPnlQhj73f5sdBaWO0/90Xhh9
gv4nYEMXpMMEZOUZ31caAGDzKvlKz9CH2owCEtNYsepfZHEjd3/fFqdHDhZ6WAD5
yecAQqRBke9zNlbuwfZDwzyh3TE4oGd0Fe6sGu6yg7dVA3UVAu8ErQ1pnvKhiDDw
lckPMqwerk+h8zw5S+BYeXIuBqFR2fXrvBLSpDlXKv3/ZDOLnPyeLwiwQqMXvEmm
Dj6HwruOGbpK4PL06R+nCnu1zgaR3QHG2P64DpmPZNWZDmJ4glElQgHXaJD1geGR
qxOm+DL4YCS6SrjWZI+XpiiKEWWGyLPpKW5pU/VhcbESa3Z5Dwn0rRbjxVwHyOSS
KaX/1ujbZK28YQ+x3+2WxGUi2v3hMyUKY8mgKvzgCBM5pmmww0htwD7ZH3A6TYas
z0LIOJGZqKVXe6ZKgLacwKc9Gc6yCWS7+MMdSR8095xN5JXBryW03jro+m4UC/se
N1clGiuXC2QYA3rMCC6pvysD1ocu8yFJpndDS2M3V27rF4Blddc8hx0O/p+l7Pdx
LMtbdv5KpFFoWnZd4uQBo4pHR20bda5oyDELT/eKjiv4okyXtmJq5SFtjO8QdMvE
RsWkCy5mFLUmC+mvGU4LCT+JQ2VNCnn2mQYNqoE2m7955+GXzdDZl/Zkce0OU+9G
BB1UwHs+/5O8HuXWyt7Dqxyt03/Rs1n8stz40Ah7e7CTqi4mrE+qNZQQFfy4OTC4
zDossh5n3I8Kc52gHYqolV3DgLIxiFcDX7YwIhjeyuPPORfkdJYA5RMNMPqn5gjc
HiGdJKfBXTW3NPz/i0s7F0gpPwx9CG2x80YZtqDuJYg20iTPAsu1U59QDWzGtntC
f0C4c1YipHN+I2VGxBFo+BlLdYg99NDZH9a87+qTGIxoTbydrzRdsalHH7VzZrQ5
6ydS9JZOEnoHxcYsCDOz37y7qRZxL4iaQfQA06yKx4Yv1v5NxwpHK370j7IIXlXD
RNLKsZLHed+yleYM2HENHqvaFMLBQn7x2DkPeiOku8Ewvidc+UyoHHR4pPyNbaB8
kDBvvjQ1GWwaKFLmK/xt0DPAkaL/4EG6XeFyWUtaugucbbutUCnBUUO05m3dgbRO
qDzG/5WtDB7c4XAtmBDYqetmrd3YlBn+1n9jwhJh9yuL3eAHWA7D8hUukSUHOd+8
m7IDOLcH+jzY3MoRfJrv7E+/kq8D/h1KbFTJicPBZ0dOqo3IuAyWcSKH8EjtjY7q
iofJH8BTgrxGVhzQhf7HRHk4X1siB6nZi7nyiTc80bRK0IoibK1Q9pNtm7CbF76R
P9MTtca8LZ8koxbNEpINvJr3CopSvSO9pDeSowlVSTr0/UvDAyWArQddHZ35p9g8
YZg0SIezY+/Xh6baWzoTT4hK3Ob7fEl+PcSTXnAKGpceay+KdcANc0xn6L8IFcO3
EzHhNbNttPAmwAzJ5lVYFpKUFffDySAU0r26EWIJhF9XCQ95Ds8GiWwO6TGi0dSk
NLIjunTsAq+YJvRyxZa7FAbpKLAYT93yjGjwq7PZH20gOPSOvfG5fIHHyC3YYtGv
S1D6bpndT9eqzjJCfPezndS1BtEvvaotYX11zBYYYJLHeZMLT+JdxQuIf/z9yq00
jePAAzGPDz22woLPW2SJFz2kWtmWJdAx5WsNezhTmscFmaelJLo8cfBe6kpUEi1T
bjaX1dpp6sAjUTRaRFVjC8B3Yo0NgNqB8HSd1hm0hLQW5PS+uk2bHRs51ullhX39
/Y0Me9McYvy/lhgag5Pd1s9q85A41eN/raz6VaSPBjeD+BD2k6saXZu6xm5VKIKW
sU9Y1VPWY/NYc1UBMr9Xv46099Umn+jLFFg5ObcogfB7OU3n1iTdgD/ueZkOJ8+c
4Ipp6FB4UoVT5qvdVrwZIb1SPGm0m4kd9q5SRTCXF2nnHl//lmhOwU0zgS/fw/aZ
I5ItfVFfua1wsWBN8fQHjxZC3qgffEzjnTsYiQ9RXswrD6tDd4Wqgy4Br3d5yu/f
poJBqzG20yCZ2DsyJOF1WUHHcu5RBkm0aW2QX5R5JTVn1EvaNwQFu1dcENkvCvbZ
Im8ROeWh+7DGvZhJlkM+YE8i31vdl3/oQOFyjrQ7L4FzacUrHw86xz9NVsXL7Rdf
lBLwJYaWy5jDZkeNFWV1THIoaiko0WZPuXDmSOFMhRSOMbhA/x3bHiJqV9zC5KMI
VH2ujHXY85F9q82bIa2lDvfY9xTeoX5JKy0OGHPM6/r+kbx0TZwOeAMT3MVg2FsQ
2ZoJhsFm6XumhltfrYh07cbt1MVu5QCMTbdQnTJ+Iu0f1MRNLS/Z8ShEuMOoJT+D
54cj7dNfC5LA3WSun6NjgLjlrMQmBeghiZtJs0QvBQAaWlYYSI3lOYvwYXQL/4IQ
ke531fIgH6cSm7H2U5eg7rr+MpHWnXQ2Z6pKqjtWJyKpMOnvMTqiGTYCDFmoU+n5
ACW1hAGNewGNkD3JOZLZbO9vGxsdxgQpoJZwfk1e1bNrerIvbSnfh+UZbZlkIAbp
XpWka/tB3EkIMvrnnB5FO0EwwcMTeKr0htbPYN1cLvV4n1N2ZiBX7vHWkas0vmZI
lYpVXZcAISU+x8by9tCy2ZMpzNbddw9IP+haNEzd+Lptc5X4FcPFAJriXJoTL9gd
Ajs7E+zXGoA8jaDcjGkoqQMHkZN0xyFtIlYvP0xSLm0XC7csSM8y7nDVsjeMkW+Z
dKlrpi0WtnU/OVdEb5duK5D2wzSMFHDTGdpGh5jUUsgsW3W78O6xluW8l9Fn+NvU
wL+xH3EgEQm2cs/3fWcva+XhUx/GkLRaBlUMG5oQdVYmZb/PjICHSVgrdn4luWRw
/QdXG6iZpIx4VG4JifdoOLUgW2wn931w4Eu551p0ttT0rEPUht6Q6TBu34tVLNcf
hk9qMzrh9axLUjgKWcYK6sCvctSC/NyjAXXLgBpXbpaItpw3TAEKSZBgRWvWvGVA
eXcEpkww0PV5Y0VCctXUjrsWMlmpwmh+691PgNmAXZEhXNkdLd34LeUKfo4h2Gyg
YHmIwqYDAimS3V3wUnV4vTysPOg3nNAC6SIJOkOSfo6AK9iinMxrC4cLmXuyCphW
qQaQ2zhMy0ZySdS4zXuxoBVAv3u8pgdXJy5N+MkpqRBVTr9HVg1zubDldRosylUZ
63hR7rXOwp59a3+2plAAvExDzGkYnaEPmOxMhxuYH8wRJyUVeXxd8Zt0a/4YSEjo
U2xW6y4n2nMBV4dgxqv+nD62fMEh4K3o5TL1JeBdVen2nZBl1NVHm1Z0pRJ1iR23
qvqaiQ8iaDbqouMV8sjtNvTT4V6YvlWTfMIuUGGT9xZIBplwbUONv2THJ70C1pwB
Ya2mHwn0ibVaICEdpq6wuSpOlD+6VfvIlP2TOpvDVrJMT8Nhta+6wknVER0SXywe
LfCOEmJZkRo+SNnceKL7O9FBzLBckvKoTw7Iifj+p13RPanKUrhPopDrwqSRCr2T
UmiV6bTrX14E6qZakr98Rpkm9ILeBaqn5176pbik93/cegsPO1p88zrVECmvStDC
yZFn+Cel/ql38ZCRFSu/iMx7YgHNDxbXj9/meZBqP1Pggfq1D1VEFyABN6SNYho3
+PHthcE2Qo78Am8HfqqaxULw7HExZA0Tziy760GEazfgq98V+kS4fbB+GHIfVZ1j
LDOZ5ntCoDviVKd6n/+bR1It/x23Jb+/oy4z3/uriqiuEZ9mJ1fNuaxDrHdFo128
LY8QA0aqgS5l3fIfOVh0QsykinVMrfVE59P3XlIq070dH8jz2c7uz7sHNJRl4w7r
KigQm0bkcmm4K6jGiyWgBpD+bHMAYvbX6J6FsldEHVvoJDCDAZaGcnGYQv4jygKf
49b7EwonCCtXLzoaKkn5qeSsNJYhM+yKLWIrsLeYKhASDLdRQPJMPNiBssENmGEF
JH9MXx4xJnM6l3lePE51bHneQllImuBq2Gm0ABy4Cq7lP/4fMD9MM9vRh6ENigTm
HisHNHfhH0L/5ZAUfymNf35vnqRMqcMf/7/UsBxqatjgnpMnEGt2h+F49DV0pn+j
gG0FZKyjAt+f/fJp58TWz6+z7bVPIvcggTueZ4rHjId+0wygY/ge4pMyRBGxzsXl
smt7KCDvOoqdkNRLeFD9HV0YJmL/qbxSEyEp9o9UoxFCQOqqPdefnZDzFLjoITJp
BrLMosFnkDev5aYEqpZG/jzBTrhxloUi2FjUd24asFWAK3JVVbxqC+wipAMVGAv6
UeqHog90CWYXLLCUB7cUrX5uqGN6wuNUB4pdzJ1zwwrnp6PyOTvqxvrby1QA7Kfj
o4zcBT6+RtxQTLQgd19Jcfiq3gTCwCJYZZQp6JYhwsvodNy7O4rLOngjdhRK5onS
TuI66eG45v5HL7CbgrzTnOLLRpgiizMYRtzAqJOUgh/p9l0BbTZ5HYL0elSh28D7
N4CKQMhXaqj47CDfrQiPA41C+VKnFXDCSMhrbz5Ur9LCWpwbzgPCZbficfNmamwu
XSIJhyuSDH8xDEr3MiixQrJUiXV6fBs/LPrkFSbFip7B1ODMbcQOL8AcxByXqVCn
Fp5eBUkq8DNWa7aTp14dqTNjiV3OY/jjE4aiUafmonLmcoZWfMdv8Aha9na4DxDa
7DENkJ6nCjkMl/riDBmpylXfBzrr13CSao03ugmJvxxDN+6lI6j1cKV4dbe8oCHm
Wmnf4mHhQb8gBEazfNejMqDBDYiq9XA1ualekOtWypgCb8tPJeUW8vl6mG0wyEww
owRhhNLZEMWjB1Hzsq9T6UvhrbwvcPz5dJqHXtUVLXJHMtM1SKPdb+efyc2jzMrE
fBZncq5VZ3iGDPNFAFDB+w/SznXJHETkfHXeiXBl7rXBJsqx6qyaL0WEuvFOHIZy
qzsw4yUQTBhfnNVkKKDb38v/54qPeOWMQ3Idz3f+HkP+mDt+dOE9uUS8KddYMthw
CKi2B/VdsP5XAUU13btZG70MQsHbCkUY6o+WrVPPLV+rOK8ERxB3/yhROGmbVuHy
/ZpuNg+ihHCzrG3jwh45fdurrBO8CK9EipGNnaEsevo/5FcqjqIA2RJ7fjfSX2QA
nVdRo+Ezx/ZceQpZjm1VpUP5yIFjzSClc83vLi8c8vDEtJNRSGAiVxweOlawnLxF
4mSlf643JqSEfuVf0aJvMMMSU/bzb8XJgzMB0tW3BF7bhaa3oPGMBVAkB+Bdi5Wc
STduQ5OQZ4+UxHCNsX0KjQgJfFZYL769xg2khYNCA8M/pOHGSUIOlw+jJyBJCw1R
uMNPcgUlrDH0XaUhgGMmRSDzCFFFr35NzVJrlizTLgvtZhhnzSVrnU/ig5F9Gjye
fnanI2W2pL3EJsHpAcUeiGJC5ioJRdyIpNOsgdJJ/d0Gkefx4js3kKkyoIpWY38B
OH5a5pyFa6/CVQMfh4Qpe0vlPnfzr7TffHxur1lAmgYrd3c/vvI+WBJ6wy0bLbST
f/WazuuaN6OGmYfHr+Q+CfflFjXQBTYHp048E1I2YinpYLTLNofiEKiaClszMB4T
JjwBDQWckGXd+inH4U6l+Jd9Dh71OkYioBvGzb0bxINOXmM1llU1RVJGSn+1NMtI
2TcVQJwnJDwbwUkqVplE/oqQ2oesvXzB6nq79dtJW0OscEVIKcbkrw8mi0v7COCS
SAWxPlZ1kR5atRwUiwmG1CpLVD5ioPYmaZXqo+wZHcJpilDTkL1vNsrMzo3pM7oA
UsKKgMmZkKTkoLwkhq/RrgCPUSkbP1v9vOs5J9QCx3EHk34daIN3C03fSX1SxhkM
FOMjahGCdaJyLLqdC2ZW1tTvb6DWf6DPcBKB8g0vrK8m0EE6jDuyGLCSV7uFx4+F
2Zmpdi0dflS0UslYlQcL2J224HsauS8rVWrd0RUME9jUqY94rDa4jhyfup6NRvVS
INnC7aMkt9EpHhmH2l3hOv65sjL6mW/o9q3A8Z86s1lM1aIRrwFl8+fvQvpZM0hu
zPb/SuQMcRx1bO/LJdj5/0EEANkMqJInXrXLC0bnnWvwW9AF6VWbvmWC5PrBsKWo
EOWbYlF9wKct1G2FpxOt1xfBVCVjr0BKjWQB64SWLIDWaLLxNXASu/kKIRck2fBM
Qo0Z1SCRCJDbo0hO0SiVYptegRY8F0LYsRy89A8E94yIjfc9kGve8HlnXGZNs8yQ
EfN2a+oICV/fnrS2X8+KLCs3usNIIhUHj7Pc27l6KGtakE5vPQYICZ6rZ0iGJYBe
um/TSbxqXaVyh2TWRAWRlSJV4H8Jg63GFZOrs4NwxjX77MQAYMaAZ1cqvj28qlnm
zIj6vUHhZenYjrdJXH10V2VhgPuABOcpg9Ofd3ej8pUYUi/yQnHtbCvEefr5hnOJ
BQ/BCusfBTyss3ouACd3OGjwD5Ty/SqrgNeHaGTMP/kHhpHvD/p5NjXla3xxBesy
8xkHu3SA3gz8wIT3CzvG6nX5QCVYOBBMY+mOEBXfVwpU8yVy6KxCxUjPYUl9CaLu
9D0x2ev1q3sPwMnqln/mByMdPCzBmzJ3h6A0cjmOWKLRiaB7LMWRlBWPmjgI+BzJ
EGw5BKZnAaXqCL61/9p0Zvw7yIYdhfX079BfZSZedc01VpF1Ie4XIEhZ1eOH4CjH
jYelvh5Hn5/j+eTXOyfMuXK0GWo4oGvjAEO6DYZOtU+cR92XpeEtqQvcT/JU//Pk
IKQDUtRzTBZRxc30Ags1Cx7GPGEIJsDLqvRXz5KPr8WagtSPOc8C+i3vS16RSBtn
eju4builraiKVO9dWu3jOipt39WESZ2o4lDkPi69Ahjf7WVx2lkdMgqxyZCp96Yw
WIP+Gmii6cidtUAti8qYlG7fZxPDLScNa9WyYXkQ0UerOElGlpOMKB+vGao1p8z9
I21tMNR/W6DRkh9iNI9BqbE2woh+eyPvpYXmISD1k6onBaKqaVJLGIDdAKgVt/H7
XuS8OAHg0OA/VByixkvSqrPYbUYxNk5qG6/HBv/QOth3BH+J/8TslePV4uamGLsY
ibdo3I3HxpAIhXww06yE/WU82Tb3a6friwcj2kq/E60xV1td2bWKnmVCN5ELQ26l
4Bv8ocE9AaNWONNqQ9k2OkI92KBsOJv7h1G4lRqkIgAYw1cYTtjYWeANTLdJ0XQv
Fo1TNJxo+Ro9wbJceUsAKHA67h3EngVWlNdWaVNuN/PXII3KAWNDNVl/7K0pGuAL
Ly9+9pdKc0WcY/82Bu8EhpPWpJeN9ZrnaVsUR9GxfM0WcTZmPhF+yoEUduyWNycy
8eqB4cyIpmAYGachL+5n4osrXlIybKh7bWN1f8WEo/Nm1j3IgHMUGTxUK+I4ENnH
+aUc/DBSUdR4ER1GzhQrWFVv0MdVgIOtFBQQf+UgqYjKPNtnVhKAkRTtEdHRrXgr
banlSwVvYE9UtZnkqwj7ySjhSNd7JbdtWIFxq0yI6+KrGDwmFiJQB/KpLamsdFcf
6zAhNwJiFVhKM0Tu18SpM4J4bkhe0tnONxOMaGrXu/EPtedlM4f30hD1+ZR0/7UJ
oP7rK9WFRFcanddkQHCxpd2d7nNZvwzaiZtUqH9htpTL5S2rZ8p5hk+7Vfv1PJBM
7zhM+YMIr+piKnAh1LxMY8aDvcBiKSWK4e6H2tYsFJDip92/ER4lRTQd6rlPvVOB
7FDDHY8yMQYeqg8y8dVtjErbW0JTGa1GyJ6vHPjfS0xAmmIsjOSHiS3As2HZ+1Pf
EqNH6xeME9hgfunTxVZMBZJ/rTNwFprzH2WLRyjkSpKaxBdZ6wXnURW82ZG/KnXg
0UfkNeUu4t1LA3QQPeTsruQ7qRHa/bn3rZDBcXAJJvK5syL8dMaudc2F3BmEnTwx
2N2sYh4ZpfYMdXiBC1tlsmNjHF6IikYVL0OFvTjKyqbGfBzbVZnxHZ9EtnLBjH3Y
kwnfWWIPhiYt9V1AUmMzrae77U4omF0i+9VMXehPgvt0FqQHlXt/PHyIJDJHHjsP
Y53WNAxGJleacjboRzV9d70QwzyCdHBIazNGXwLdhWWZgxnnVwLmBAfdLWF+P/ma
NVRu7eDEB2O3Vl6RbV4/uuIgbKP9IRHXLP90ZOkoT+jyHVlJSiSJLxx362xRrmJ4
DITFbN3m5+30OHCxHYYGGLYwF5WK9maSZFFuujfEnAHvE3bLZad2IJS1RtwjmsoZ
d6EHJTAGN54PQ6b2ViweR4CvldJUH/yQZwxskGs6m7bVmLpwP+ZBzio2jesG8Gid
Ipt2quJ/Mx3tyTNTiPUU5ms/DypIaEN4IG3Yr69OBYMdNwp0XDKxAVro4ImI5RAh
7j8xbfsHkK5II3DmjwQo/PidvN3LAZa30YAdVSO1ctmqqOKT8UZLYU76jomtmQpB
QBLLvNShhD8K/rZn7+b7CqOcPDu95Y7CbM6ulX0fUorqcXyCWIbSapn8Waf02LbN
mO553Q8SlvznbUWhhWKDJO/nK9QtdWfIwSHJrYmHtL6IV9kwlktQuQ30HNjzqG6/
GQmaQ2X4N6hQ+ofimrX1r/wYYQXkT+V087EgTD+ai9oqE4nJjP6xT1WkSgQwQgGU
uRJFgR2K1PaS379TKzkccleNXwKFAjis9wgxe3Q0OY1aNAOnnPb1aG7f3DiG/Lxv
tv/ZkRVcs2JTiv0R2VtZgmHjLdJiEH26hrELkzyLvzlbJ4Y+kMlKKZawRhSu+9/S
BRKkgAY2Fm43/8QP9G3QiG5mo0HOdGLijQkO/4ZxDRYYqwR67VFuOUFcjnkiWGEf
W8Xad5155MxXf9buhUNDAUHtOunTfX/m6/we5PzgAQubaLJkGAzCBgwflEJq6ZKn
pVguWt9/z4rQ0D0/WHIAZVHQaeIJUdO+UpdKLm+J5AfuNWegRF5nYXqOot5mjyAn
SfzL1H0UItWQyffK1TR0BgMExlgXU02/FTY+nGHT8HECzbaC+FqqBR5nY7Zxg4JY
ajyhhmi5isi8+hchJdkvaWK4YgcKKs9znHkbWphqaF7kvLnM8bTUoVFqs0XUwXGN
x/R//nLda2Z6fSQf9Hzgj1ai1Q3SdKMtTzRId340u1OCcjqD1p/e3H4xEa6tOK6O
cHT3EYlggBonGlU8aIZNYW1HOsRvw4SPEWr0lqmG/oXt4cI9Anu85cIqAihqy2l+
CZEGRqeBetz2z6qTTBgF+7Ha4KZbN7O/FMY7DMkNslgBLRKq6/4gHrw8y6qxO7ze
hxbNGgYU0AEd5SuYRzJNfeCxbOcOrcFq5KsohTtX5vu9DsW/JJe6Bp8fpbtX1COR
eesrONbSUJzpq4UbWjksUMDOr1EHvVOtj+MCkzFqRC+oh4OQb+57x7V/JaeS8hU1
BFxEMdpX0ExtHsCIBql5YXT5xRYcX32jA/ZgkVpIXgLlZAm1fZH3ursS6W6j8nj6
PsuR/Kex1PO6VsaMXLVra8FP53ZntElreVQAAKsskuBxUwZcJ0xHwm5HN0rJRVnY
VPCGEJQa5W5P4OHtv3G8tozGXOpJmBBH0aupC3QSMWwxb6newGEvV8TUXyVFtKBz
OOWeaPunmV3OQ1apbcRT+8fy8egOlS01QCpdddpVgktsLhMRW9e+jc34Yd0quIJl
B9BttluMzlSrKAw8kvXbkg41oW+sIf+mWjzIoko80cunRnM5UqmfSfg/zpsMdMGm
XlMYEdKRWmIZdLy8FuRdGPrdXqOg9C03oI7GDZD0kpKVM0g6ZRawfFuAf10x3Saj
SENJDPGUCMyfRfd3p4u7SYwD4gUG3qk/FAxEd1YYmFyNnpQ9LHHlfL7IVHd7VRHN
uR55ZvyPlSSKdEM1kes0q/nvoZOamfiUHDHWSFU2z4PbhW4hPqbzp7bwKkUJvB97
HjHhsID36gFSEuASVIMopI9BrYUUcD5oa4usKkhdaMBG+PMr69LoAjG9/1zWZIfq
KKVSaBmmW30GNUIiLXc2N4xCXaX2pb3fx5yKqiQgaaHSzDWYh4dFfND6Yrguz5ul
Zob0NkPWgtBbvX8Hxv86hF+3dxONpjgqDxJbZb7i+0tnuY30XETfHcaTkBgz1zjd
B6u3JMrXIFU9e6o30X84XO1Ix9ZrKd1CcahsSo30K/LESUPOBgSR/5HVbUcnMEqs
KqDbzynVVUiMGzG9Uy4buijzpblLfVQWIA70e9u8z6SIsP4YDAZ40z9FE7cV6F/4
/7SqXBYDnMvdTdh4gwpWUDpRannI5VqxfV+OAI7wx8DbHkoXPoUe44l4zkK8PbFi
ZBN3VhUoopvcsslCFa/wVvghenQDF00p7XLGHL3A5mwdylC2TboWFa/YS/iNbmbl
VNbE0zp60eR+pl2NCEzk4I9Aen8pHlp9bJkm+fLwqDmJ46yYJB88n37C97VeMpg9
u09euG9seixLKV52AAoaaZdwDHPIsMMqID3hmY/HN1SVqK1LsAsnGhnQiEfGoxW/
P6ZtCvu3f1up+yfnfumwx8h6bNe9aBKUSqlU+IHH+Oo6FGnvalVHNGHjQG2hEMMA
CuGQcjOlOfKpQf4Wto38JUMgREK0j8Onqp5VWSer+R+2dM1T1Ty6RLuuKl5/OHJV
qR38DO9O29XSgRKBj2HtZOBxcEuYDnB3qjWUrfaF3V17Pd55DCh1eBQCmXKXocig
yEOXJLF2ni2MHGxQiCTqsoqeg+dc7JfMeocXxnauK2qSaX0w8POvjBYFLXMEvbw6
XNJ6Thpyy3aHb9RC8JVFzj1+QxQHlZCI6sfaCT15fpKMuSepmmlsi/4Nerpo9PT/
9+tDFEmTtQJL8vmNAi+TyQ0gbeV2gSOHAWnV5Xb2YxttfmCmUu+qg336fQTXQ6F+
ltIMVAzXxmwHGzeA6R8sBZixxtTT4rxRRKvEYxlaQwY4uSc5q4+NXtTx3NhyaJQT
N18T1J+/o6YZWjwWNkaZyosRx/iTmfFIaCFuXEtmLEL6rYw5I6Ri3MNEnzXM6TFc
zmWdMgpw3ZoQymKr+TnNK3LjJavFLFoBH6xVAjEsVOcxm0VaL/8OotR6iQkNNFjv
FhRDtUxng2AqFnzBsdZ3WHmgxmozEevLLfnLt8tyx1BNpI6BlrV6neWAYFkV6Uk2
/tX6xO7pKbRmzB3I4Ger0PK5ebrDD58tLd54eOtljFL+ML6wlGjD3RI5LY4JSpJb
e2CZj5BX2MYjJS1i0g3Y7OWjKPWdVxJ4GulSY08ENl7hYLRZAPHbHLCwLLVL+wPI
eGb7mqun0lCyB61XxjQEsecOZ9M4Rm+BPM0VfE0Tf2dM+9zyH+K1EGt2uqtKpIDh
vROBmL6bu1FLqp9RmwtbpFF1H1t7sqNRaXWBvwJ7aw5qocRZmhJ5QysVwgQ9Wbe0
kL6g1ZTumgf1S//+B76I7+mmwMpFjbZPdBAbM2UBAVxZYsXG8TYLbJtMzReZy37B
tlHQaTZZIlQ9SL0Uxwr+fSGFjIci8E/cM2CD5iq9DZy9rgSowA35iR8lcEDNSQ+B
pDexABFvPIaB88saea/P9FDn9GbU44XBMVKDFnW/3zclDFmlWMztAUPgd/qxyD40
1Kj28SyxNqOAftdhSpZMETO38CiOhdUZB1dsm32F73JcTEuMs935lNaHglqdZ+Qu
Q7V2zl89rIL37d2du8iS+1JtXl3JSL1wom8/r5dOt4SMIMUeAXf6dSpKPCo0CCeX
mLnMH5mkkexp3n3IfnjpnabvMSCjY9c8Y1oZQw3tcAGu/P7HzXckRhgUvhxrA94n
H7rOLftQirTWrRxkXOrLJzKOII5SHmLU8y4L6SsdXVsC8KhAUo5g6pPA38HTdA/h
v4NVB9nsWKMIgrdaEgFw7Yx9Jctaa0OvWj/ISSIUcYnvRP8GdQ9WtWCl03PdNy9p
4eFWQpm7Z80B2ubSvtF81T5gRI+WVOTQtUzOKv6zYchhnpzsobeRD+5tgvxc1Zl/
7mtFrsKUplO3g80l8TqzlFSIELgCLryC6mw9tNRrJOe3Xrwv4WX3aAm9jzWHCidJ
4zJilm+qT4bWGTu8gTAt84mnk0aU8KwVvHlcnCTjNWkJ3MG2MoupxFhKdDa9NCof
122gv307ATkMHztmZBWmVMqaytfEPn6yOfDCeF+FW1plCXPqXbF29iuOdnwrJSTJ
qWEme7zf8M2gl9cpYZ8uw/XGBCi9y8Fzre6TjVH/L+aGZnnBOifUBkj53Iye3m++
0zcl3HNLUMkxozjiqRkoNnDen7A7gQKZJAQ3+m8/N+jo4MpULJFVva3Pwksy8aaJ
wG69vMio2k08STwHnBvU3YBCsgME7mhyyoqKuc7JO+PBuSI+fADiQyLX47xqvZhE
zMh/M8yJe58oP5aDgyEXlrGwf3VfnTrS286kfGHbUFfZKyGpNKAaGafSV86PANKu
qZXNpE6v7lrn99ptihF4r+cDDFqd4N+YtDPLdD97KGDXsIoVzzVEI3ERmoXwi+34
WorzFX7HFRkFbhWiZFna3co2ErnDvoUMs0G1b4ULaNuj8Pia/kTkTJCoKSf8RuX6
/Kq7cALcwFpPhaUoNWLjvEsy1xs8SWMOSYUxwT80flNJ2HCHz3aHZRsInp9jVIFR
MmULwx2GU110Jfl49wICpxltA7mu6tNNpEw8uM14kpaZyihdSPpRcqugMbayEaC3
8xwNRqz9zrloDp5d2QxoAT4GRhELPTITMOXXjKiwfgzIQ4f85yfYYgOusZdS1A+7
PTevkpH6EGwrWgRDV6JAD85kYSiSK8dILb3V9DdGQu9keJ5xT9t6kOmPLFUYcZOn
g0ftSrdu6zSTt8z2R7mpC2rBKNJx81QhfnkV6idr1GCSTqN7VTXmaCelPTGAgTks
nNrdA0p56rytWkvr5yO6630JK34RP3YWPphHsMAp22C0XpstR5JTurjmf1jy9sKh
mSjJNezoY4/pvOg97n+FG2UY0AuPPwsUmTBkUSWeLD4vJrWnM2cU9gVlzdGXqswx
WCMW/+ar2IR5mduFj5X76A4Ntbi5lS3vNqd/Gj/8k5WsUOMCMp1HaSeDNOnkSoDS
dz5ELBwsZwrEhDOmObC+E2ua8Tz8FNx639cc8CvVpyRaAARK5EKHqtFsP15ZmnIa
stdxzdRCF8oZjVqkTCyXmpuywKwyXflxfCFE5zlLtKOpilocaeq4/JhfOsdIUNsX
JsOvb+pOUmrRSbID5UtoL1zmcJyav4u5u3kDbTGkQ9Me/z5QJ3H6r50C3tneJGbp
uct+tAh1K+GUxYQ2NkrhDo9a5Fx+8UcAuIMOuqA985NwxpBbcKqySI9U4W2EPMCn
+T7AUZ6aOAEiHH7fd+e99FgP71MLqdt8NeBHbN0EELTxO5Qey6orGhPhVU1np9eU
CDlc8VVCjrxr1T9eSIDuEvY/f0nTPMRyVAFgQkyvbKZalrFjHWB1ABJfF/jUUbSi
RrfYRJZ83hpZ4NbfXPQMGqxJl1agtNXs8x3zK9w3P/hB4eKRNN9rj1A8oo+LFwad
U3o+3MC7D4YtbjbF7O9hOZ3IR0NGGZDu5U8o3IqEYxBWlvgCBXKTXiNzYdxZaKHa
0zNtiOhIzNlQE5+ryMnFPxyLxC47yLTIxU/phjzXoRkpkfSLiftYB8ZvFDJLXmZb
kCRFkphBMzCnBqULwj82scFCA4K5O/RjvVtB7Y0LehYneA9ceFggGgGdsIbDnMkF
ksJIZRYus0v1sEhmQDlQFoWWoMP0UmY5OqSzR6MTVy3ThFwJUM359JC0qbqcoppY
5lvCt2cpbM2wBfxpB+Fkfs7dYZ/xnNqmkqe64P/HropHO/8/Q5T4wUcmSjhaB3fk
UVT1s4r0UcVecEQm1nxafJefHZXndG36tAEiRfXfeiCp8ceY1wm6Iq4ce1Fdgan4
O977ypXxFFxVSdYvtb3LG8wmCar7+WhEqULpFO9xkzbsm/7nFWOt8sullAcMsqcG
LVRd/9J8SGRdMPdGgNfVNI5PizQT1cCcQKZjrqvYTHLxhFpNS/4RgJSE+TGJ1Rl/
oy2rGeBO+EDNx9nOy+4uhRaWFE02ofYlkKniMVTGdVSKStLZkAbTzJ772+hESkf0
ueNA6LWDj1SfMmTUOTIGPapWY006NiiG98+ps6CqKUXPwzVdLG7ibUfMDk3Abt+X
CH4AIBBYDL5CeMV/rU1YSA/JOptCxDeBrp95eve72iNpMQTuPpUeb8cKLCoFBqNB
H3sBLWiE6j3Ll5hE4jnPspvhbr5pJIpeC2s14Juij+ROO6ku9LGsetdAd9nvps+Z
cAiUBOAYGFTJ1hm0We3w6LphU+4Jrd8Wz7qsAPcKl0f4NW8HuUjo3CLbwFre4JCD
5Hov+vaAmnvEsYSFweZG/GmHVN04ghyJN8pFPsijyBCO/nBmJbMuhTPawSacxPfx
NFW61J1zkzmuNDt+BsYDIex4gczxEZZNxdyVOI1bIMmifpFkJOjXAhKheT91WdJH
sl/BID3/2IKPjfs/wpLupr8xw3lvenc9YeY7Mj788KXr5bJMyMTzMtmOmzVdJbWw
D9UN6qSCyMoqAqzOfV4gBJ8kguHDyUsYJS/76WLn4M8zzZEx9JJ2Aw+jtbrXUkDu
RnmCvnq/J7XDb/k4bYd43JLCmedV2yQRmjp5OYKg8ct2wNINyJCWmGiimHPYyUWp
J52Oq9edEJo39c/1rFsAN2DIisf3NhmL5m5lAr8Yu9RRtGxr24zog5abTS1WB4Mc
OEaeb08Tn39cTpF+ws3zQWCYzAKVfItMcVDmPxLVAGJJYSuQ7mCmuXSgPiSqIYq4
qGXDAZz3BJul824dp1hIkGghqtceJc4eMFEUrq+b/jRg3PElqy3GG6DlIJjOchi4
zfJ4dXjC7l/sl72Gy6VCPPY8AtO09gZaf/LAOAkBBYL6mos2BOV1h7pCMNsuxQlj
EzV1D22dnDKE/wHixlrz1XNoFsEmGreXk3tHEUFXnP0ui+DqTaLyyQxGqSk6fCzA
zr6EGY1kOcNX6fXi/sOJfpqGYTnhY2BGtop7dxY5LYns9z3P5ZIfHbsviqnwipsE
all+8c+ESrodhJiGL1z/1ERD5Z/mq+7FyeEdg55YBCZ8s25Z+QY4VoL1HH7oxLZc
qYTgiD2PQAazvMFWwn895c1YUDNmRQ/Yxgrarfiyw0ss28LBMrcEq/Iw+kKTJi2e
/6jkz+7yfaOvQB6+W7e0/OOM2nj4qZXE6+JvErDA9cv6Jrv6UeXEjdMr/V8a51fn
5b2yFzqE6Dlfmafp82RVAEtgMCRGyaL4Dk6ZsczeuckM7QF9x0PCdzMJPaf6ipys
9SdVjWpFWwhTVCs7cC4soJBHr32leVNIDaKGybBfNksdFluplEpLAm8hjPWzksRy
lKd3l+Z7Baa2ZNA/3ara+uAZfjm9pSdi1eRWlvIdCfxTFN5lAkC05G7Os1Lz60y4
+GtifSW5T4k8By7kuRgDetB/U5ldURfK/XdyIw5tr2UyFrmnIZI8PaYwcjPbQDoq
dzP9fIU9JOwm0B8c92FtilrCl4twGFn0zktLQi922L0Y4QNFoMtNx9LcYOjypkop
YeGGe/nkffJ/IHv8Z8IYZFZuUvlT81Jt5hXRobp2iS0XmVJgCYqNioMYiha0Y8+1
av0tKVWNvJbuVNw0N803PcrAu6ZO3ow6E/aT9YjFyd65O5lggm3BWTFm9nmSyJLG
KuJSuAP3tS6w0ttYZ/uR8eiTrs3oxURkxK8UKmKKFdJOCIub4mwPPJ1eHAbpEynL
P3IUx9awLKXZc1xl5FGx0A7NLqDuvvl3llNrNr4MYqyD3b82vFWa5wvlH815rRcs
QfgHmXtUyFURwsAnNiRSAdwjT0rlMX26rnj3o72s8MrxYdZeBPy6P0qpZU7eGy6G
A/MPDyq1SNrnMM/Cse6WqA361IwHrYud8+rWCl5mvC6x6hTX6Sno4BQ9iSCXV6JN
RtAYgbebwKH+tWrtqitfQrUhnVHikjWEF2f5QgMum3srMRoSPUk0RRrCtyDn9QNl
goQNo+t+4/OO659q5HnqBeq0Xiq8SSp5ydUmxANohPcf6yeO4NTijfm2ZIuI7AFx
xyYAfTofZ8WlCEyHKenV1HTj3xZYZtiQJ2+eO2avAIbUS0urfJCV/aNdqGPUhYcf
KHWQbQ6XApCin950AU/9ne48mcFeNxOgGXftEOGRvnPaLw3qCndqz1HXGd+9To69
seTK6OpYjIa1ttS711GxtU59wLq//QbM62gz0Ze3XuKXil4+USGD3Oc4XGHPLE/d
Z/JebaHVDQo7wU3Xvvj3CEpOVJru1NMGesNcbD9+RV+q/PjTgb3/viFczzZGW2U0
m0tJjt2z7T7MwxRR6AcXeGZo7njUpnJiTJKOLvaM+rLFD2HJ2Lrwd+Lbzgdsno8v
6kB/vgakxy6Gzqhv/oEmokFgs/knieYAirT8WsjIIbG7BlsT92A6OK3IA9bW+W3R
7CPs29hr/ykIVxKO3h6NrQIpS7sr/D8qmr4Nt7Y8P7wYtdQ5wXUP27PHSbwJNC5V
T+MXUEau10QZM9C5FXacTLkktJ+K/fhOkkP99i6yjHIFi4Z+z0rCxxu3LfJ5bwpS
V2t63gDSeuQCyS/Spv7dPTk/oGBZI2STVnTmr8b1jSt3TCYH5kDypFze5Rs7bAHb
TDP/NixOO7KiG1heehX8voTUa6ElftVQsw6Y46wIQ2u9cj8CqCmL0i7h1ubvmu/W
4PnEG7ovwo+1qmn0woHmYlait7oYtfgrzOYcSLftoUGAPuYSPySQKATlhPqdV37x
lmroC2HDlku8sQwo/aNOFw42gzvbkayvktVosxYUY7fqxLJBHobJvT1gDmlwiRmi
HePROJIVn48nT59DWFo19+eNQHRSp/j7raWz+VZwQKu1diNxusDsLLAGjrKAk1dE
MTzOsVU17OuQQ4sSSQ9j5+/uTJRGgK/N9dtNfjfRhMyf4sVefkUqnuQnWgwjUvmW
TuFtXlGZEksNPl5azrKDnzncSqiN8Px3QsvnxiAprOTtLC0Qfq7AF2A9fFle1o/2
mx+Brsflz0wiv/+2b2rBPg5uY7t2IHHdQYoXPB05Gszo7J/Se3QC6X/O8hphtrr7
xBZXUJnWWNXE1TP2D2qtPlktkd0qV9xY4433wbVEAsZnfZQgt8WTnXB/d6yEHDIa
SbJIEIieZMN15jnvNwLnz+w2Uai/5TMKJ0O9fMyp2hTSIykLB0eyi2HW+fht0fWJ
dy6+6O8f3t3t9vWPPNCoyQE6sPD7SOCQTcODWQPJGdZY+zhkXfiUQKMg29aanF73
qg/nj2LTvP5S17e6JYS4a1eZ+uSEgHDe01dXMlg6/LcO73KrJn2GaH1IgIrmRIDn
5Ap6tkPOyXQ98tEqva/jYVdSVm5HwqbgqQBbLAhtZQ7bJSu1CvUfylqafD2xX/Gc
zaf5TS46TNqBCKfL3ElUWHfTuqttLsOfXwzsOeYn0JCkQtdHc7wfaegSqDCHMtlG
wKTGFjNHMgRqs0cxVKyzVZUzTL0T9xHg80yWpX+BV1RwS8yMVJuKGda9I4S1CrT9
Ghzz0g6Wz7PgcXSpDA6RFPsLaF8bpCeQSrZPVC/B/aFuQayfO2y/QATKU69daMkV
Q4GcKeplPu1423ApktMCDAiMoQ4Gp0L/2GIr2XYsLClwFYC57V0dPj3pN+oQumcA
Ui0KuCouDd2ToJrQFUXYS6IGt0B4mXaFBJt6W77rPTvMgsVmv39h0IfqE1WEPtxN
WvgJqKG0/Bg5CN9Q6f36gAIWzBiz9nya7VNP6Be8zLS9+bcGohMoLfC2cVRkPLYS
fVwluq30JqpWppUeDTW6jq8bln1Q/L2rZl2prKkZwUyaPqcu1FOBRYjRRrWf+8MH
h8OlTkAX0VkhxMgiOVmZQIyEOiEM7PoJh8SafdlcK+iDkk5euit4i81/awceofWc
bvdui8U0+UZdOcBXD+wvZf7ZWmQ/k3WLFwI+lMfeDKaJeGCbhGi1sajATQ722xEq
fHvpLdjZrQNf0n5d2OzxN1ka1mpfNjSOKah8BqgG2PlFyqbXk1DHfwNr0oV++y74
/tjs9Qf+Kt24HGwcTI5uZ9SucZkn3YcXmx2hSzVY/mQixlCOIuhbjVByyuwWgE+E
RiJba+Pdc4AFDAdOKFM9rPecFdlKfPT2Kqt5beLNiYW4dDAvDzyMFEiVOpA5DKGR
T32toDfrlD+c0GRfPih1Rjhf4Sk10GzvTZo4K++abbd8gQLcWE706TuNfgVPNCWp
YbSqT/dcD/7N6MzWNXQIUOlm2G2SMkjaa6RylLfiyF5O8OgirnQAo/Exekmq8yoF
O2BOpJUuDXJkg3j9IQo3rl4heJ28mZJ7sDdVde4EskfuQUDgyD89CgNqGpBzRwDx
WGtBX3/MyomSZOXPo4V3ouCHluIWEmRMzLN0lsHgJ4EltqcojFJbRIHMmr84fHog
5+7VaMemTYrHRy28J98XyB9FBJ5rV/arZILp8jKbuHbFZac2sBE80yvUvTBfR54u
7wgxrsqrQVRf4d/ZrEgaV59CilW6njV2JLKz1E6z1dwUJbxG1n+5+/H9y05sK9Pl
0VqPQVAJkWJETSd/n+Gcv/BDJG0O8eBeo54UOQVsa9VEnz2CRM1fMyij0KM5HTut
4hh8BQG+LqYQbRPwApXIAV+Kx8MvWMrtAqGWtO/XsNGKp+4bz3hCvUpvLsI0Lbgq
2wT15JT4s/qiEKWyTuajXa3KefxDxF3055j1kEeOXpchoA7lywj5K5akg7l3YeHP
oVa9x/vujYASFmH7Q3HkHG1xTphde1E/3PF0HRN8Hr1uUlBgqRPb/xluvbJmdyA1
4YKfcVQb6jRFWUBVblbvukWCXs/PvSs6UIwEZNd2+A7Z6qDm0zs24sUmTKuXNUrq
AI2PznAEIKkc0H56AAd3mRTsy43G4XwcsBmQSxeVFssELwOSj/3hN5bD0hUOq4DU
6hK/YXyEKSea7ZV8wMGAGDJEQUxPwoym7EViz3S5UMbJNYquHDfdnBMcDw8XoBGb
QkmMNYDNoALdfcmIP55LpWYlDwyqszJ5vmgrdLQGLhbne/+BUNnpN79/+sKNksy6
TwfDO3+//4Hh1GlcQJEr8IqGmb+RIc48SwygCkf2AdHzc88OcBX+bVWwgS7DUJUp
xn6cRieTkaWjvtYE5S4ylRwqPBbyihToXI2Rria01IX/MZLEjNuSQhVqbgKde8z+
HCAfU6DjQRLCvPi+WzkSGa5U/NmtJNMJtxh8KDAJfVf/Oghd1kcAKBgRsfOT+YKA
//f5P+LdFwmr+VEpiwEyUc9zjbQp7fUKQl18o5jV550PbysR7MrNiRtoqdLIcwwT
WUWVaqoxfkxTKeHHwXyX3yu8Ofepxt+KbIkI6Y6jlMgJ+VT5DrcDlaXeV8r8tWGu
CDrbbvzlApmYGF5f3fj8+HOTQ6azbY1dCjfNOdfWltfYLONGLALXyopJLaTuD6P8
j867GLGAcgmANs0oqwVavDJ4r92PqiNtqoRQU0pKYkrHlvUknk0TyFvfgzkfeF9U
EnCoofeh//wx15DS0P9CFgoxvpBuHRU8RGhr6s3PUwbxSMkKmJJA03cdDTyWgv6M
E/SjjzRnR5qv06yYK1fQJCgDTnQn6t9XYBngy7tnnGJk2dUospn1Zv3psveDa4PN
S/OsG1flIP0moczIjN/c32F3QyVl564ADdkQYUO4EsQxUitFj86gph0K5FB6rnhe
vN3rf/uYuhX6AAgFS0tByH0KVZS0l0XSAEwnrz/rvVF4PpFsqL0em7uxNMjzlPtV
dSY3esenXcfo5ObjjQd3ieAGql8dYb2/oM0esJF+1W94lYTdPwJ2SevDlQtHXPq1
N+2X6U85tEQIVPQFJ/c8LpbjXhAhays9w+0QDdnHlUzxa6I+/7v/PoLB4ysxpQYy
hhcsgebEF6+uGFziOhgUnnMCg0vNHODxmZ6uXfCX0IP/gvIPC5dwNAcVdK8s5g19
6HFqTasWSqU6F6GG4qKJoItJ2sn0VK5W7sCfU5APsYJd3wuY3ukquwUpwd7mFago
n0jxOubWD2G7ShRklp2xBqKZEQKnj/VtnE7MzRlcEGlz0jfvbyl+CAouyZHnWmUi
+Uqhc/9QUKJ/3TrF0J6HmZ8fWXWFrdW0lXjjtWM2QpOyMgsANs+k/uGcmZTGxHEx
VupJYO1tXs9WM+8+gbWRG17ZmVmonvGMs8qmiLyEpGcIHzvuu/rMLVZhqA0GM3UO
pNa+cF2zbTQGIR1z7kWewVL4W9dXBrTE8Cna4MZlDexWEr5OwIZASzJTZEfd8soc
CMepcI1gKSvzfN5PFedYDiHdHMkwdPNBvR+N7lCerhfWy0hiAk7JDaaRgu9fHC9r
oMLAiIhKviZq9La/Vbco+GmTfCCSpDQa24xRO6pWQaP/NLYFmuowac+nD+XDHGTD
lK9ER2SRaPULrLXHaDpvLhItmpqov2Yf6vvqUe0khRqOL4FLLgl73kJ8G7KnkPIN
BgYJAVWgig6RAoXTpeKboTgz56oQv4FMmYH3/3tD9trvc8Y0QSO45gB028zrguBq
o4k6rW9khHtICEHkw0q7oV2eHKr2BNNI3TQ0ertIAcOi2U3TIWJixVxKxxSHOenM
+QhwlFzpuDDGi7Fe74PcNhv8ye/ytQI8CxrxTUffaB71c1DiBA5P7L+GsBZ0ZcOD
PRhzVnjDgxtebrhT/vxV/e9Xh6QmfTTjIZYs41Xdcs28yHnOL3y3pbPvl493LPUe
5zhp8b/apQdqYYTAV9gFStaKAhPELtHblFmXpxzDj13NTQAfJt0mXDBPGbJkWiaV
xP3s2/QzJFgErLZkzKNZxNM3yZq49xrTSFxA+04oKLSTkUaJhqt8efEN7SB/E6og
0Xw5swIWQeM1/HHsU1EV5t/gTVlr1kwJJmAGwEJc56JysDHAWavXafiS10XSI9CR
FW95uTKNckfHN/HGmuZaKErjWL0j873ubIwM/ulg7JcUWVLgOg9P6KrFTTkYrO5+
pAD1vKBLUmpIJrAePGu4KLcQgVEMrvzluSi0+xaMNIU/wURiEnV82VkF/i+50enU
Yy4N4oY6MJlKOkN+R4GZ+5koRzvNnuaRMe3wvlxh8YI+OUjGG4AbA9GZbNcdISwK
m6st80LnEWfeH7xGd5wM/9W4pkcb0Ohfti4DyVyDYT8duCzLurRZQvLgp87JEscm
PsHmRSx/tM7ceOs0KXnLW1MpFx45cimPgqps3Hm7/5Ld0NGc0IXb4p7uS2IDrLa3
1izX+B8w5P94TjPdxDfHEch14T2hoHNcTX16VgSVK763y+a7wi3c/rFY8QI+TYRj
qXT9MTzeai51xc+BEHKGn8n3HTi3eU/J1yRln1PmZ7qDJPVYom0Nu1BEC34/RgfW
olIKf/g6zc2mezZOwGCNsyISVIi3lFNIu3WSH+qvaWcjLiL0k7hmKdv9MGgckxkW
MgYxTrNUhDT//IAf9nZ5BcP6xbjo2OW0S4QMy8uQ5nGhL4Zgw/sz0O/qkkPPDuQv
qM/KhAWJ95k3XS0LSxpVnHhlldHoiWBKFGZ2HoRgcKrhTTeqwo5uJMhDnRNY2bDG
B0vug959LMPIcu+NtFx996P3kpMYnl1BymDk8ROJuUt5b/E0VV8XhvFr2zrQCezB
GPvkBpwebJ6lQU3rPIlx/JSOowgtP4AlwA4PySmsObu9llJdEeSAEgkEurztfUk4
rBfi7EZxNeNyG604k5xQKy+Ba9Ll5RYueG86i9UrUXncJGQNcFNpQNTbGuiAtA9b
VwOUA7psuBrlKyvZUqAj3B15271jI1XbpbKzmig1S3wyKB6XI66E4vndhtdLCsog
AtpI27g4lZFfpvgGC3jBUGXB6SrW1Wi+Oo0epZ8KF/od/xuG8+o8CaaUk5surrr0
g74qtXJ0V97rr6dgRQfX2mVrw5hpEaz+tX48eQ5YpcpFfgO7FC0gGTrXblETZdOS
9xJXT/gVZw66JViwBnnLsLMYndNvzRd9F03vLpWk975Q0ariua9pM1UZy7Q8LYg0
sSS9eChJOxT46BCQpgvRMoWgyo7pYROBaSiLvxUVMhvs1cCaWXVXx3EWxFQ14zXa
Z9mTVbSoioL1kwGQtWJFDzVVPri/t3r8JL6OiM8iT+OHadUFrtWwGPgiC9Rxj+14
hpVV/FN18zut6GIFOK1jl4wZXs4QO2u8C12VfBnuvDQlkbJdWUFAjIVWAd2bodgP
mzc5Lc77xQoWWbcOiNmC3xhzwikfT6GZjmVFt5OF+uttsHpXk97QE8Okkdlu/cEp
gG+9jAHwN0HJXqlhv5J9t9Xhl2V8y59lHBbFJrVQlvdwclRofIdKaeQgTOdBW3Jw
XpOJnTRNDCWFyttTmMeFGmqEQlpkMG3AU/jC9Md0IgliO6HJIbp9bbQY7ofx7+em
VroxRYdrMoLO1v3jcO0wIVzNzS1zuFablkFefjQT1TP/xQ3vq6/TW7mh/xVqRa0b
AP25/2J4NEkZgvqVEAQDamI10yXDfpFjr+zASS0dA3oGF/xb3wXXIbpo/Vupd2Zp
blcoq/2EyURjCktu0CIhtcttU8o9UoKxp+cSce3kXGyvvr0NPk3U91UjW1XCrHGD
o7iL4PjG0/DgLpPghhGDlyV6n1tM0HK+Fw2fo19f/b3RoklvvFgSfcGvzW/tRlwF
WQeM9WvRlYmhsBj/puDFeB/VmVJ1qlfgLQLmbBouvwhaL29UrUcLMKrrzvitKsr8
p/IAv3Bb5P89RFG2LnPeIUjyNX7dzkM2VAlBj+9azJQ5F8UNckaQw1AVpt55qS/s
5mqzg/tq7Mg4UyjUA2/ttxzGV2OxTqUxj/DD4Rp2YZfTSh5+YkbU1ttSBCnMgfug
2ZeBokvksPApbLF5ky+zhgOVxywDnWSaKX3hWtvs23fue5hkGqw4TtdY3+Hy8GXy
xDP4xMAsZtEHZ2qrbdQrMtZUAY9dgSULP27+ZrFBaP9car4BNBvpi/3CLtrm07IE
Is3BpOU9mZuaG5yFJS6ZF8X7bAmAw3pCQDqhAn7hQjV0/O70689H+qkivVHL98vy
p7uqhncgMQGeHlaKXxWaGcUn/+lcMM+ohDPxd6e/z4safHeqVF75znh8qldRhnTL
GsVMNuZmiKPvTF5kNCvqmo/ymxuugzcpGvPsr2Bin9S6iQg7CN5FyvBVyaXvm2FY
RMhv5z6WO3fB7udrSz4HaHUxIFP6jAuV9+bd5TOMm38q48pn0vu7Z/rBcnlnyMRN
tBV9Jwvx7YrrATSgslPppw5yVr5begud+1/xd3Aabz/l3nZdYn+qobqgRbfR0Q+L
WP1sYKT5LRu90zAqLxfug5Zng4Sg4M3bV7vhTS1gfmGtt2sFu38jiwJSwJeQuVnv
FEUCE/LAPzz+kcPAHWDbdJcPtrvtVlaLEh9rdcqbKKWlfY9OO9c4gIwlH/G49BsQ
hpH+Ltm3NeKoozAZHjzhS/tHMfLcj7/FlhA7yGySjtQiLrVWBsdxYY/VWWxCgoiW
X0Q9HCrmlfBKz/CZjDa+Jp4q1REVdNarHFS0wwNHq4s4jjYtx63d7UzyrFgqYk/4
E+2O5e7W1utjqiQmvhW2xmA5BittNhuVPax0wt7HmwJzXL0fy+XWfeULRvjgKbHc
6ZBa/MOW1tdzn4t1Q24owXSsvffxizHsp+PLjzBrTG/nUh38AbPkT+lx4vHNEGE8
jNaTeyMsDXeNrJRK7ot9GVWCK4Y1hZ0UKPJk0IsiyhpTAPn33ZMGIGOIAocDYE4i
Gzm/F2VjOjnZ33PACr0QUspqbHeaKQvccUuIZWaFrirwh1ip0WSgbXUTf7xnTa2L
jf486/g7YiDLEiFrU/5eOLoaR64c2oiKdRZfi0hqKN6wM0YiSnLFe6GzpDv5kbFi
8mqmgKXmYLV4+WCRWCe5bDIlWiWasdnK/Wugn40BIOwcPH9JEsh85HFO/kvIS3ZR
ker/YiKc2IWCpsscafWjvpEKhJICQe5O8tPS41tvZtNyJpMZuSUDPJG/hFVobIhH
uOTGWwR3SWq2/q5HlO1uDGzuIuLfe2T1Z4xrELKre0zq5/cB6wMrBaqSflFARSJq
WnVVQnEHjeQ5xPcSA810mU2TgJHssbHS/yqFHZZuUoE2ZGK9ltPp6hlZ1I6uL6dP
6gVKpG0epVo86Gz2Vz4APU7fQHXj944TYNppE3E14yb6oyiEVQpJTx/nMSIDG4Ly
+huZ6SdCdhmb+V+t6ZleAAW5w2gD46xtP9JaQovhoYkIjlzF0U2ZVqfMRLejPF04
S3LPS7WPxXa9395QAltIqOz7xOo7cNvYpBic/f1Od0wWJ38179rPWJ0Leh0/7waS
9RGcxGIyXu6zNR6WaGHN6HASAtMuG1SBfYDlasNW05nO6UxbwKi8s6MPfjZOYFI3
d6Q4JS9JTnq4+ILEd3pagDwju3wgcXSRN2mHFxeJ8G49qN4TDu23Iv8PbUGiJaHj
nZ8tvRWuj3P1eKYewrjSVrDooH05vEdcCn7oLxEsNJG35RtZbsMrv6+NDyfuTkCG
M7pQYRdvs+bc5oZQFJNSZVq0cqmNAigarN6LvP44ysNSEiZjOAUiMwvZn6Re9lyI
/Ri438v5tRAjjWxX2bpYWOcu2uVNpmqKCQnqypIHEm4aGFzw8uVcJ0IjJ2LMZ2k6
fZrMb+Hq8lVWM8Eh2U4GP8NF3nVh69iexOTltifSenTolFxx6bFJV6FxffvtUnoa
pOjSJ+UPC/A1RyWH/ATSC1hk+LO1j3gzLYa66o1WURJ8Zmr8o7/6afiFOq41393V
a1LXbuHaxU/w1IsopQNs0VwguWa5sY+mLnY08iiBWTNBieMLE7rQeb/TwbJiKjpE
DG6HXsEkidSOM1jVKtLS5ITYWbEI0KgjMe6nOgVLC0MNpK9a/oQEx+64EMuO/D18
hoVmiG9mk6CbAQS3pHJzVFkwaMDaGEvbAJsHNqeVfRGNw99JMDQXZSIoJiB1PD79
KvFDbScZpom9jK1OlGdtTA9dt0S+GOKRKk7x0zmejtKBAkHmxSp9vw5vCb0t6NpD
LXM6Qqd5kHwjCfA9+KxroyXcUs3tTsViZgMHPuQ9X1v2PdZkAhLeXAQ80ob/gOR2
E9j8jHyeDgYjCvmLGtVsTjbwcJtSPpHerU2WDm+JCBM+JCkJvLU3ljQNjOxg4DFo
zixSrR6YTO+NWy4bmlTSHVX9E/KjHERZHbq3RfwnPvSdtuG0V7T1HS9m3jBu6WeP
4Osrg/Jnv7uKQLc/LqJLlmxjbbmREvwmIibmKUM/5wDyagsZdzm4bLJD4Qlyxs16
34WuHj18SlPIP5xD9OCMX7tyKB8Iogzkdf0hl35BMRHksHHNu6Aa4lrSVx+iBv3e
Ki9FtIe0KcnTyIGhEwMKorg/vR5Cw+5RV6E7y/rWSVTep2xCmb2hjx8zm4e0TnlJ
JsNMgF6xOOEG+dYf6TFggG8qVBZQWpLBBP//IfZg7MWpzn3ZCfqajFJ9Qiy0H0Il
hMmGA77QHmpM2bVfQIfINmvGgF6/OZynIkbmmHk/5UVLkc3HaEWu9/B1raLe6ZTO
S6/gKEoHOW7UvY6c7iusfAizjTBGoYDlgd+b8CFYckZg+AEdiE+yOb3e8DR1URxc
mDXlQ9OIivXUmjYYS51fQY92lclzaxY+ITcHPbiLslUZZ+0UPxiIMCAEWqrDOPTl
oRNCk7clqrorLMYetjmb1HhAXMM3qRo7k6DggkGpIMoAyiydIJRUiqYsCPAaBtBZ
HNVpGjjGC6zM4dJj/XlhVQWcjlE/US/D5BmvWSRO08SSkior/fdBdq6vN4NCKLbg
57YQ5w4KN/cjOc05J1bx6A2Vu+lGunxF4UzPGXKY6driqDgfF6vH6/TOloNgxmbP
zTp4VIDBqmh3g8XI0Fhy9djSFajeLoZWSrxb2e0HmkkILKIYsbeOU5FHz2ZeEiPI
PcO0UXtphTbWrkOqtFquCPKoAkNyp9lsV0WnbT/fXZ5FVxecPijuWJD72JlGXo9U
bxyEotxPBrq0XS8jVLa9noR86sq37knYGtK0WTREd8WSYy3hxs7iXUMfaLKWkymm
IhM8sPUT4SdMvwYQjvwBh+/8xR0GP9WjbGmNBA/L26NOvmUT8CuH6VC3TfxX+RQq
fZDQEueecN60i5diPvfTfRj4ThSxi8jN58tfXUGYxmqU6hd2Qi2PQwW9XK+XLTZM
1TIrYCb4xsvEsitgCCyoGPqn3I3aRfhQLk6rksZC7wMNkiEIminZTL01cAfg07hJ
QFpdfs3c3bC1ef8+eJ/ylQsUxLjYaPlCT36J5ISqWF41uJW3eZiZAfSWx5NimCIg
9e3rcVF4rXexoSZZ6Jr9QvSQ299uVucVwKLzFFX1+WIOQ2tFXJpFsy47LBw19flt
BFjG+vdXIJCZsjqc2eStDmjbfERZdhUm48TVofW4pEeqpeKJVVkZnGuQpS7oYXWe
sVFIkS0UPIAn+3YJTzKR1qX5zV/jEGJ9LSmTgMXSMaRYgwmRQbzJ6UjJslLRaJab
AvNlU5tPY5MxPSjxslD3KvEQUfSK9Bvee02eMuz/TuHUEuJ+pUDRnUB0hCmlfadg
fXIBwbz1nCGRMLUiw7yTmtRaQgvtO9xr1BT0+fusl/bE3dhvSvDLzSqpOtwNGRR4
YwkibeL4C+Dhu2XNaTg0jCwId14ld+9H27srcU2rycAC61pLpbuchuc3qPNNb8aq
RMtd+akvPWJtnAsYCTfuSNW/kMdLUWZJSsFQMksaIMniu2QIchRcAuwSzbId1Z1g
bZxoGI1tYexTRE5CGnWvT+DBZQRK9yHdoSlk6R4VfE2eigKr2r7xAWDVbOIq3svh
te5ZzVfN7cJyAn6rpKNPIYlm26x2sS/h62mxVgqR8Xw4jDpAfJtoGDEHMp4Hkqs8
vuAYzlATJR7PH/tFucfwIV/jKfccB4fdNWjDjE+Jq9S9Dp19X8VATSIS4cLBTeF+
T5acGQ37xrVHBLpN88I05ayGMuxOaBRY6D+7ZCp2aNNOQfg++1IP80ZwYHi+6wrF
cOKINqKgLT8G8AaIeyUZv63+PPyoOdz1AKCmtlioLzfsOPGhSaOKwxu9PYGcA56i
/pMs6dqQIO+buABs98CQ/wgam84hV9zg5A793AB5jx8IYBO8NRHfyGeFQBqt01Fo
u8CMHrzvkjsgv2dz9y2hDoRmE2s/lKjL6M7zOzX2bFuidOsh/oe5f8nhoHVab6UJ
kg8szeTgJXPD1Gq1CWpeo0+Tfx3bgBODjmjhBpXu1zJLTjjErDp77e0Ibx8oX2gr
YH7yaWyrviJK5oEDKOEXlu0u9NPmqn60mW/i/nKe7Clq7rijX6N5e/7TJqRhkZb4
k6NTFq7Efm6eLf7sMmBiD6FH0tVShaKb7kKe+iL4pmu2THKTHuybfcTG+qZp/LOC
8+5Z9B2ZE/JfdZIoQO/FzY/DVcjaUB3reYU6y7A24Qa10GXQew+9vHwVTxIOnld+
hpWeHquyJiCwJVRam1VN1OTw7fq467sgFZVCvG1zIaQrxqrqnov9wv/zbCl3Cjqr
RZNyGxiPobWoPgeufG2MB+xjTPovFJLMVcEelDijcIMq5zJPqdzNlGthZLQC/aF0
nPTq0RzkOu0VdsSgHfwAXscGKFjDT7MmALBOkHqJLm1pZ9fEZB+KlXHHJIDt8/jZ
/n3fjzvhstM5fnbQDKzoe+TyRp5W8LafvjmOTLTHIJ6tvahebzSQvGUae8f73FH0
103f3w1me7xsjg+YVsENthMIXnyP02e3OHuCa+FKwG5mGfHDpAUjYDAzTXTK7d8k
dmRBey09+zQKGWYKKCcJd3hqocYVviEOBu9M/4X2tcVrD1lk1xTc51LJmcVwSTf1
BHbUAmeEJcUYz7PMn0na1yOtTFsqbEaOAhyv/JB6JWCkAbff8P5+uie0jKMkljja
E7d90aIHRjgO4k0mkQ76yZ7Uhaf8kDB3YHq0nGFbHP8f2qK2x1Wh9vIN5M2YxaDu
pjroLMkw3b81GHI7TRpVxe28cf8ZkBmO+3JBz/fZDt99/NcqBHLAhwTG1QxL99Rg
eoy0d/RH9pV3lIsxiqWTDLPnq5kWo1hHz3IcImO++Kmbs+9JIOQW7dCnjVsqLAFK
w5lHJcyfv4QMzl6qpgTWABiRragTJ0xMEfY+pANENQFbwH4AU1mz+VCzhL922Hwx
k9jPCy609f/DeutsLqEz6hZb8tjKq9ZJonHvermTngbjuqvaiZadr1xXcFBLdC6S
KAXePOODb7tiqqZ1PAYOpkG5HQCvwm6ZknboGJ0U/1IgXYpRme6BNy5Z3TO+eizQ
VzNQ0qXKV06nbTSUuW/WW+nljKgFuJXvj0b40Cucs1v9Zu60aa1hRv1cgTBn+KN+
i7jOFAKUYrAL5PJQV95ZZZ3dMlZs6EvijIQ7xYyUNJKSPAONbuYHasQ/zQul1PMO
g+tjJP/NqfBTjz3j4OZBR4sNi2vX1RXFm0NS031xDDbM92iM3+ASYEF9uxmPc2GA
LtCAEe+CWzlOKDwc0cUSziQi+onyvQt4luSxkvCVD9P1rEcUf+rg+Qq2Es+Mvz39
1xdU1iT0i1Or7TRG+vQvHMjG/l8aKBQ+Ljp1QKZ279t1hu+j3H+922dkMn43lZsS
COYvPPuQESkSY6kG2TEhnIQdJYANRGIQgD+O3BlCyC1S06ICOdlBnwdxNbCWjA4V
t1zcn150fwbS1PVBAv/NAJi3/PnJQIuh0DvLBWS9+bhK6vc2YIwU6CcvpYOqFQAC
8ZHD/1mCrfhSV7t2EdFc/pyRSoqo+XUijFYXjDfEJ1w0DnFJeUZKGYxSIrppnOom
4flvMEfLdTrfjgBV9UowDCA7CvgLpQOGxQUx9Bg6+Hw72SJsoAFXlKq1mw3k1Mp5
0dUoJulqN0v4wjp+shuakC6LlxXFuExuvj0BTVgsWMxarMb4ey70XD6SFv2fNQX+
XONgSjhXS428oyCYuyxOJ1IyoM70d/iwGAiJThjFq5QYE7orlwCx6lhKD7NrrQdQ
sYgq9aEz6f2oqHckV7KcAb6N02zEW8n8SwP/FnE2G957l0NLGNkIzKIMbNpPvfSW
mzYuytxu6wsf9jx3mhSwk2UKlXsXaxz1l2HGuluClI31ipCDf4d6bWzUlMM1Yadz
9qIMhI2AxoAVwRLNPrxsk1vNYFEfcBwGkWBicnR+Azx4GOpR/1QSVCGzbV5wxkpm
nF7Xq2F7oaMvL0xGSKH7IZbI1MEi2mD0S0Q+Xdo4K/ATTjuaTz8pZGL0mDa9viN5
Z7Rm+WEMXnhZ0hR9mYJ+k+1v+TRURcNtWC3YMVzDay6XM+yitvIamo/NaT5l4hXR
R4pFZkMCOUPCsXNDP1GhWiJjAaJusIWSjuzC/r9s+WYbJdVMR43HljmqP8eFiXkg
yiNfGKjhzfVK0vaCV8AxNsmLTj8TI2smb/i1svUN20qGDERnSLXTasb56DTdAXGK
aV8OyVQ2EhlpOmqIxQDH4E+viCiYqGMiMWJR+Qm7wDC4n8muMCGpfhmKOSORkwQr
LYY+ayH0iY0Mp4Ubm9clk7all+IAzvCJjutXndm8rWproPbqxBVZqhT359N34duI
/z4edtOE8xSdD+wjPT3z66nSJotIf1Jh/Raa50G49QM8qug6rd0xciF9gLP03JDO
7cxqSXYNHS/GfJyIG8QSV/WRB549pa8kFSy0t5fEvbAhQholeiSm8hGE07g6bvgz
haKq/TWMIlAkjRCwK15qrDFNha/ujlBWhtiKVebczBqxqGWsx+s7TSA+dgwTqY4Z
LLETYiANKsMElYQvDuMwVVVXqqx1zkLmc/BJmPBiMzj7hbj9Kf6Tk+7wIZ2WU+xa
RSvgWhlKT+IRWJljImAKI56FFEq4nYpzkpgaNGEJK6B4RS+0c+zWWT723ndGH3lb
0LQ6k1JJvlR4fC5zrxIpl09Te4OxdlOd9kIfoBKo/71lKaDTJgAv7IbRJ1XEWKzH
Bm8gfCdoTLaak1DmsnpNxjf+09RivomPnOPb9xtMQqpD03NHLEbaBBS0mPVt+pdm
mNizt5wSkqURoAJoQUvdRY4+d3EmOaoQp53wA9i1AbZESHFUHqe+ceGa6HNocEbR
RQoUV2k8qBYEVR1yDWTd2wqtdwanoP44NbX7jdKv1MNW7RVRiPP8Oo3xgdT17eEf
vGdp88UGE7yPEN/F1agcU8EnuYTwdVpPCYsOtAoaC6rdolkJWa3joCicDn4n3w1a
vEHs8QcuwqidL211gxq64mh1Gw6cIUSeJWv5Ikh71ASTvt0OB4/ZOiPgcvukdttz
KviUh0Ie5fMZ1FlNk0EjT+8QowmFB4Ug+y/3GK4iJHM2OBqy+v5otRZKHHJxob+8
S4Q9cZ85EthYQTGKX9ES41tyGrld8a3LlaWWyTX3UrbNVJRHpNdiqVklBxdqBMh7
sQiwkVYgxjjU9J6h+0qfC1uKiU7sqYu1gYJeFpxlzXpO8EvWrcmk5nE/x/27mKIZ
JcBFYxaT8A1w0XNo3CJlI0TzGnJVaJ2kkqCumr08eKZ7PfD1tI0wHtakz8aZB0aH
XAUGWPkiJpQ1qL84IpgnPd1vPTY+HHf4pF8OUgQkh4wChG7Oyycz7gxw9QNidYME
Jf5V/KnaszQTLib9QtPwiNQiKe2N7IdldLFLBXiwDHcxEYSuA5wCjXl73kS/RaXv
Mj2gamS6z6ZuXlAIMaD6TlGfwOPMVup4XOBqMs4SyKQkCzrphen63oM+kpy1VDf5
S4vO4dJTk/HvEfDpG8DlSqVAJpbQsCjP9BWRKO5KqTooumdPHZnxDpxi2cj6nYy+
tEsY4Hf8jIOiNPyKf8Naj+ttlUzpKizSgZPr//VjiBO4/wnCaiMpDHBjqu/hDaad
qEIo1l6Zit8nl9/Fr85oyVS+w/14UB90yDASdd+H12N+G1NaYVVjCxAAlfvXPeKc
uABAnCWJS1E/lK36FTIxsLIOZZSdKN53B8e83oaAvZQrkI3iSeWa3Gt3w8CFtZDw
Sc69z0ahN2wvdZFfmuYBV5n+Ut83H8h4ADqpyWUHlM42qciUp2/JXFAAlinkeMt+
WbVgX/OZn+L7TDEpzwJ4HI4mM30+4RpifRnkQK8RrXOeKsMNAq9Qq610HQdHnHaj
z3B1jJvYbwy98bcsH0ZMxVybORC8s1wJhYbDqwqeTmTw/Ysnh8OdK2DemCR47m7z
2T/4xBILVPVBeievb9SHu1KzmH4tHRLrCIp4GWIS/Y3ZyDKkC9o1j3YM8z3fVifu
CrTbSZIPNzoEQkXfKEGVl3W6FpPDJM30aBVBBt445G6qznPa7rjrbC86tnFw+86q
hyhVA+9i1ta4Qr+iF5/wBi7mvcB8GF5WjbVqHuujSWZunArUkyMot+VziDNTqDI0
9pI0FwvTLWyw/UFl69049RrPDmaluAG3xVEMdXdHNgGTLuLPp0LFdCr5yAK4xG4X
QO61tUfTltpSYw94FHPwDfSpj87tFTxIWanrTVUGnhuoQKLas+MysBezq8w+kG3m
fi5y9lYYwaZvghcZiebo+uu2lG/8s5uprqBWfl9aNQN+k/2RGQ5XLn6EfEoZVTOr
Y1AcU8UsVg3KitskuuMlQl45xIIE8YykU5GoxbtfCP6u0L+9S9kdgPh9yLpvpZT1
RLKpdtmHPziPcZB+QEuufEJIYphStTQ+vBePzeNC0lc93AW6GOrRGrmbRf1BlVXD
4PQWfIslpRbaLn40bQEwvx5YaT96k5q62WpUtQrdYdpto7Ds04j2tTJw0S+FLYMA
sgxVqzJi2iCRE5Yu39U0imXud1G4XFKm96MjDbpK/MsG4SniWfL5xG6IAHDIjCmX
MpI7w92UdGH00jGvUJ/MB871HVY2biU+vHWJYFzqyYeOi1uq//MRfeJG8YNKAUNR
ZzRt4RshF71+Cdop04luY5uus0zH6iC6TaF8ALsNwZxXbhjM/pAOc0wuPRzFjtwC
8sz78YfC2vgfVnc9Dgnu7ntdzQY1j4zk0J1ZsP23cCYpo4/YncKZPQcdbP4Gesg+
s/1quaIhMnd/ynFrWEYrrK+Vs3+wh7wnNhXjEAvxRzg2dfEdCGNBYGnrmE2LWqYA
8Y7bJ4Qn2+r5G4s173cBp1ntDsYxNezk9eZuMENUZQ/BDS7ZRIUNORHFl5ArpKrf
koV1/BJzxAVjExNIHMLRrOgC85x/Ru5GHtPFXSZSvSmo5vBDvQiSXuqldKL1zmmD
Fk9ui4dtyd30c2EMRalgNTm52x5rIMqt7VKZJrGMsuom8w2mJnXpEUi4BKb9/DJV
+Z14hdi0jVDyF5Kj5tq4JBP/0vz6Umtr8gHrl8I0ZLrQDcq1HQVoG9udoa1CtQpU
X3vdEvgO6WiYPl3/lkh+QxqPyeDVi45zGqCvZaX0xeL1e+DnKoWM1dg2i6GMfywO
YULhHXSdPdoPJUOIKJEvv5IQHdHPHglepHJoD5CHlUjW8MzYQGS29D/is/4IMcFi
fT8DNFHeXjurSqmOpuQ7WtxRwGh2fDdPuhhWSDvGo2cb24IApdT0+PLWYm2BfXOT
3bG1lBSF4xMN+z7qq8HOBS1+H1dbBgI4VGx+KfUysyjfeKHkjMVgq0j9eb0JBUr5
T3nMEU82Osg5itpYmqOp6uE+aCEoh8WQTU05ceiEwqqmM8rw0jkKpyoa3Ix7vbqH
DdjIGWr6/5a4kXMhMCzYMHSpa5EgmTAs63ckwPU8WSSCdq9B/kU78Z3zHX/ZLHrn
s9k61k2fMYdGsmIfoaUkXfMIDP/ZMRum/Z26CvZiSSzcVnQ9gPFKvPG0NTQm33ME
UJ6WDAfoP1ZZVy4DrlPqUgwTF893Q/MIK8/04XEn7fgashvfVHyVEQ9Enjq2lyR5
tbUxbzF6rFXVz6J6gwTCscxfCqqXHLcRdrBEsYSqU4wVyiUF0IfhGFf3ARtJFqsq
fDyjwbIecyOuzkF5tHa+GRrPtcyqwwrzbWWPLHX8h/D5cbE44V6qxamoDRnocBVo
4MxT/xtHblkG3iMIeyUKVaWQXIhO4Suh1f0Fm5i6QUoQdj0SQPZbicUrWZFtNzfT
XzDC01+KO6KDcF8pKTdszbh9mpIJcvQFcHZghnYP/oKAD9NIY/NEqwDYWZ6Rh8WA
EtzG1497PWT5ckNJmL+oS1jqgNU+tNu87AplFP6oVjeTlNkOxhk/vy8RKyE8SSMS
hUYqXCqFqQOpxp3RA2lsKjcyBYtG33/b++L5R7qyRzGL33uB5w/VbzchonJqEQ+7
oNeQOV7RYPEctYD+Yg928vJUO5yUIXxk7yaUDE6KYiXyOb1+P3XCNcsE7UqcMTOK
/ZGkGAiwHwpt4hQijFp3k6QnQkSTFQjkSNCWpD4vvlPQ4DfG/nhcQjDKfhOP6xcW
gJoM/1tIJou9RwKaG3/zDpRUWMdvYxGi3k3JT+/3aSxPFMC8fkrnW77Qxloi7iB4
6IZyPGNNwXyU9oWBYIDJ8HjnKiu6BJVmM4LEaB2qPHgO029E5m30UkTAh+Kql7qr
d6K3NcNNczgHXDUCbs6xBGvgzVBDiMTs8H7dHOAULPgbKboqEOBkIIm1FPBd4v3g
5/d8vJsR5qUQPtG7UcEMlXLURBuun30CuBNZmvpyJouOrvu7ladWZXkAI12BQ1Hu
SNKxKJOj/ybbcXqvNQSMAOfV8C3wwclcrTMlcyRj0QizV+XVwto8OYgkarRz2sAz
WUpL4ky3gdEaP55A8GyQQXPndAQsLF1dm/fKcN4z6+E2IaUtkqzFbI27t8UJJrAL
Nj9xyCBNUgc6ZLFnbg0TBSsLspxOy9Cx4v7YVh5HnJ7gG4X/xU01s0WeUqeZAlJC
4sLTjwxt9lnO0k8WU5Ahtw52r9dWOBbTHdeWjbBTFIFEjOxjn5MNSmnzduWGN1u1
USiQGfdwuoPgwZ2YXJ+QCmxKQMi388Xs4QWZ4pSc+P/1+t+pXYk0V1iXmi5YLT8y
ZRg+gpNX19m6aihl+GRJS7hd/U9vs7UQpw4nFPtZKTeUY6UGf1bBBiozq3w4IRw8
TiXBKLqStJaKGtRlWyiQBxNcbZlOMl4qBb+NVPaYwucXmBwW0DsfIDf6duKsPTWu
NR3wxpf/dZHGfWw+WkEDHrG48ZypXH9+6ltCPLNktOsqgPjnrqFb6904m6g6nOPH
LGOmt6vnTLP8DBR+DAoO2Eihvzf7vLB5VXZh+Ivl6gi2tus8WEqzA0hdJclx4zt0
Wwjg8IJeEhUJf0qtL1U+y11WTHHDdffKa4TzWCKfoLCR2vb05hGUoB948eZS2N8k
6RNW06tlmTxOtNZckV6jkdX8LrlEZrqsL1wOwGgd8v93cVFsVjrL7xZjnz7nLUJT
uHMhN/HM7B1BXanfsHTJY28XGOvzBlp2kubHoCEilPiFR3zVo5Nig/72NOsZG+Jq
p4EyXWkf138Sjz/T2ZbDBuqql/+OiVHHxBNoLzKZFyiEYF3tgC7DKFB0uK62zqQl
CcoXGm1oGk+PIOI1DBCAnzZM+lrqRlOiVLNDdWfw9rE7PMNPILxCFAJAtoEw9vg9
EmRH22XMUv/dePWxHMk8XPgSGRNOcb6cYpZJFM7cbPwBDGPH4b59gCJ6AJU9l0Sk
SWfO6Wd6ZVH/81BLGlpm5ARnO6sMhU3f+c7XN97Lb6OrTRx+QZAb4NxtLB7hpzsQ
a75yFYs5nxMQRVEz59pFlg6fY0U3DBXerv0E51Pn9v9IUMwJlxJcqbD8yHSZsaSJ
LBsLUUucdrKmNqJ8sOSeroIm9Ac1XAR6edsu6TrybRkyX6vz3QoTprlCGN3wR38D
URShQnBRIasbKVSDCU3J1GzUb/pMpGesN6s0j6Sp/PBde7c9/PGvDu/iRiBNrlxU
bqQK8dRcLRq8e1zOccCOpO+26Evv8W2u6OR92uOcz18zJ6E/Aq12/d0LHPGZG+uR
L8t5yWOeAgFRObF2wxuzoLzebH7aLlhCbpgGhJsaFH6hiAN0umhOZ+MmIg/G3f6/
HQ666tqK3Vb9vE0m7YmLRLGrfUtRHtfxLzgdp6oBwVzhiSfU48c1DATBy6FPSa+/
WwVHXxiYthDVE8lqJpBvvcQdHmU7l/9GlM8hqo4xM36oopUDayW+O9xTsWml0J4m
f4zNRjUf09hzHwyKsuTDwBwFxD++f6q4XvhXYOooP1vsBLi/qE88CHXJyiydvFkg
vUbg4va+FZapz3XxVB9xb2K4yl/ad/+pCpWv8EYypV7lvefQd2aJfIZh6ODQkCSb
pKU9FKqBUCFNShmJoopAmADLhmvCrSXKyFXmPq/eYfazolpnmH1C4qkFpv4dkwbw
GNTu1uKFv1zh/kHX2+rXpuoj7hrgdLFit262SpRIA30TGGQRoyEy0sIo6csfOcAS
1SjObT/3gi+AJi4Rpnpqrw2VPNfTa44ssB7tmvrkZAdf4FFGfW1XjG0tUxS7jGAs
oSbJKeZ7bycO1tPbX1EaGyFLE3bwYJxa0pHNaVAVuL96vxefOp0DjSJR8xf58Maa
Fm00vgAvpOYsFZURKTX+BfLm2xKhWeVnsoAYpqzt6f+Q+/dDiubNLeYr2mHu9gB7
AQapQ32v10sBrYQfgQ35+IkbtHfLJQtFrFNqJxl20J0umEbC2SqazjMQsWe8bUCl
EgwhJsJ5hRDEL7t6XB/VUYhUm5PzHPP5l3OfFxWkPssEHCJ2xDWvSsF+wKUiF0JP
UmviuxGFyWVsDTvAb7lmM5NcmYdfF8ISzTZVXgpAFMMZpk3ysy0PBpOF2z0kdY/W
OqTj828fh3xy72aT5QZkPYwGrxYdMksGLUy9psrXMOCHdf/URUEHulrK40jtVXIc
3M/GthFCW/q5hQXOxmdMOKlecehr90g7Z+ugTeLXQnjuYzZyZw1Ivp9tz7DtL2Qo
+fyiZo0JkPJzVthFsq1myLV/E1b4yxLOl2T5NyoPe0J/LjtmPYWHWxHLu9wPa5nY
X2mHUJTgIRMti0HfgPv/dlOFVrOYTcoD1C9njY3eHsOU2diY4msES8hmh7aNFEQ7
c9zGxosooHCmca+7NO4tv+xP9raWmdQrFHU8hyouFEYgkD+xWG009DPzO2nh1Ieb
DES9gAkYLA3mrrO71SZ3bszHfWQiDRpdhl6g4bPXLZESYd7YnspBDJ3NnXxdjxPC
GaDePoaBBc7UjoIVxZgMCZIMQGaTTXTmuW4KjP9OMSQmGB7GIb6ZeX8QK/DaPuNu
8KmjXg0UtZtU1J58oOWSFhheKnMqTVgu8z6+tEzJrQ+2L7l+21ze9vDxgbM5W3p8
Udc+E9TjSpASBwXx7FwZIzLVDFnP9CrJvXM/bjZtijFtIoulpZMgqhmHBi5igmOn
tGW3a/3OdZqBuYa64OGdVdqeXjlHL++AFmR1zeIyrPfNrG/LiqrvIugx+jA6Kl8p
9gj4DifC4Y8++6NWOyYOmpyJaKJ6RFAYTA0/+9aaSwfeV8YnaaNqQLdbKC97BSBn
Y86g7OddwbBsn8Yl5BgOq3ERamnmJbKR8Z711L/lobXAlAkXAHod0xJtdLCeFdLM
HK/jhS019JifGhhlDU0P0crhg78AQ1qZpYvBzHE1YEHDPkRT7h1jW/RN/+cu10A/
X5fTlh/OYmGzr35UMxuRmewuVq0fNDcW6zfbjr4KIISt72r0mAVelHeAZSor+3mQ
OfrgTut7mvgjhQMMMmy4Xua8rV1w2dsUCqsVTwShVfSHJ002iD1MKD4+mDhOUunJ
PkOszRNvw2KFitd0bk3L1xMPaDrugDeVLGcQuM9xTSHZ9BW62O8khi1gnVWUzrT9
IY+YZHf4DeYSYt38jyGq6ZoUiAM8tC5KTU7hd5oGFxR/KPykdpEJ1pWjBPX77v6t
jKYOzmGJvn/nGd6Z77aHBRHJ0NECEkOHrog+oKZh9VdONQZslhPLJCEsHK8HFhuJ
gZaU482/rP2WFMATLKfJi2T7mFbYj/GHzsI04720y9gykgoM0f5WTUXjX7si/+NL
kuPMrraxCIi8KSJX2w2V/BtmoMzlqT+L79ZRN0w+0Mjd3kylsZXZdrgenUizQURg
c2t1AA7dDfEHTkBGIQheKeXcQgHWVOHDMdkz2MzfiRFd9DxeeZQXuZ8JDf1JF/5b
NThr33km0eHeLONL7lktvnNKBSa3IKSGBSAnaLJxXthk2pG7hYoOVKUDFdz+Iwdj
aXOCkEGkTKFXkNz77+n00kA1GU6hzDH0TuVm7lKLQadYM3p3asUCNICfFl4ZE8gO
gQk0gw6EImzltkVwxt8lJF6iHCsw4x8gR00zxY/pT7QtB2WzEIF6rp9zDI2R5YDQ
Y65Vox3o/a6bESEYlhoFa5TVbHXB3e5iIEKttKv2Amx86vlJz30zupS5Ly32SuAC
ZdryALHkm7fJG/4bQXSxkgM8mSNOtmPKnlBRe84FdLeY57TbdpH4+KOeOHDuEmlh
QA17VY92UyJ7UkUbnXCxQfRdnUyqOYCPb2/y2o+ZJUu3WEPqUgmfgdgb1tWfjW4n
tTNvvDbuUOUGJiGxGI4SYIc/VzmJScXg2DnyZAwFOc2tNlyO9pk1x6r8nX8Hb2wH
OVE9L7qCzqtLR6M43mQsnycsy1akxvc9uKloAttgn4ppHUZz8+mIklu3sEgNC3BM
zr5ILf14zdWZ3D+fcofoXMoV82qZTAiO+9q37/GkgR5TwIJzqEvWt7KNoOCy2QZK
hFF7TEHFcyEn3R0dGlUnxhWmlaXD1XRYL1+XweEtMnIgDfrTbJ+/a+6DJt0Vraeb
aZWe6eQeG/x0I9XljjjyoQ/NMX9cr5xPBGhmk+hsXTyG7W4sV/j1y8PyQvsAtUjt
7vl9N58aT0zZHQk4FxHk6zzFc7LYANGhYtxGC6cdJQlnyjtdRMKYuyf2bk/1JYDe
C313B0PCsDqIws5lDH+TavGrVnXDHOP7eWPRknojSGpyvmcvfnfUZJfMQEVsY0LR
6n/zdy+0yiT/KAA4/kWPpVh5DBO9lxnGOHDqdoJnC1acgHFVK1WgmqOexnsyjVAk
p/BD6duMTA74GHXTGh/eQe7LF6AO4HMK2ZpitQSVBkqEJJ/RrqMNs6V5yiK/cU/Y
ajDIrX55i75GPDCfwhcljqDo2scb5Ue+3zAZjdqy9Mw+dIK63dDx9xM4PjiWnY/x
/LMtObl19QwI0j0ZlaqpTrZxQhiKr4Y753INsaKKkBSn2YXnN0mg2wU7mYjdaHyT
3VoDcLQrUtMIEdstYPPI2igYsClFP/956jSCQbblCQ84iJndRt5mkmePLEgqUfac
6biiP1DmIz2j3cJjY6/E8J+IzCzFC9xRX0IxWnMJr6j6cX4ib1Tl4ApXrXe7ZPTJ
0HfqouQ8AMLGX20/goKWHaP2j/xxCLcrro8VIe0H0WL0MI+CTIaLjpw5BqWNmFy6
GQHr5ZhQGA0Df5Fzd7fLnM6nMJE+Y7DUjb4cFmUiOFSonW/iFH1AaXSDCkeNpC8n
lmHWiWne/X5tWDI4dKwguGd8bpITV9fvCaXKa/+7WbRyCBxs1pYPFAtL3M4iCLcJ
U/jxtM8JgNMuQxrx+mxq2ZHvFNh5Eod6Hl9uInyXGIDKRYxjQ4PVr/IHiWDBAHuC
Dv2xWM5B7ZAuw5R7XozStQJTfWmyM5zRoi24mZ0Qt2/Glp27fqn7Fu6fxFLkN6zI
ELQFY6tBojkAAFNqzk7GAPPXAd85I8klg6PBk0DpblZr+koaAo1/jmXVMJtWqyPb
7QsMCV8AIbK3cankSzVjm1qt2xh/Nx+oDMuq4JOTINJl2KtQbdfoOIIJxhQB6gqf
xFK6hP7q1XUSHodxMVWWDVDKQvCax2XsbXIyyOW5s1KGPhOUaG0gnF7Z/kvUFdYq
WKFnH5678WBnSlsa6rmlIp8RktjMVhiCHPzN8vrFl+FqQO360E6jAIGF/FQB9cPK
NMLWR+/Dk/b5j2/F8SfgO9rcmZD4xrJHM3z23klGo6ytrCMFi1cQc+W50VqIPxQS
3Q9ezI3wfDTo+B+D0j5qTZs7F9cBevk9A0lEmlKgV6z6KHyFCbJej3L7BbLszKPI
c476ObWMxbhFkfAT8qSNKvavi+yRAlsq5C7lrEg303v9xzHMT7T4FVdMKBVfGS81
5x1zZF8MZb0G5hmtQ01AKsAnSNA+O3pMl71IYbDbLj9qhsMfh3vNZVhgMStGjTGE
FMVPQ4HGfd2hA4Sxjo9zNlpfxBmsi2wUv6nzLMgiRj9VU/vRAREWHGKHpj9guZfS
7pwdtxgw0hpw31vIt4kOJDabW3jdKwCDHMCM+mnoNZ12Tl7GY8SWLYpNHvBaPy8G
qRcPzuwjyLNCYgWfgHkFLBcf2vh3mFy5Co+YOEamMRiUiCGzfNkDV1JW58lXhRml
4Mp2W2hGjSFDsUhkmE2ID9Mo8gJrOx+I20qqrqlgGEI86D7CYc/pv9AgmWi1Xdu+
MCgfLzb+bygYvwRxwcpGYQ5L/Kp99Ksf5/Xa3AGvhkrTcE+bgE7r48Iu/0TI/s+Z
CspurG2bMgQleTHiylwW8/zIGfRxjChUL5iQg3j0HAMwRQmPfZPNM40hIS8zJvlr
zkwK9ivrRrHH/KCTG2kpVip4eSYUsPc+R0qzdzDGaDSJVj8cGv0mm0Pgl5Mjjqqw
rWeUbG06M8aGN5vnCLtcxDOOOxOdyccoOn+xzBmRZGun1EGqfsQYPcCpxB8TDTfS
Qke3z4TxEUF6suqkU8SAeAsSvpeQArEj3bFBAL+rm289l1gtUgP68SXruBymMGIQ
xhhDayYAc/HdXls1fV02YlBsrh1fHmzlSJqgbXa/VZ6zwNDo+u9qcvHChTha2jJY
TqvtdXEjio1nTnQwuw7wpVtl8kZ9PRX6yxQJKuth1mOdP4jSyvAxxRGTRLKdDS20
PrgNxq0nh6yRLGQGIJo27Ka7lB8VfEA6FXCWgqA0nhdV9ouE91lIMmNaqRkRvVaB
EpDZJiNaB4jeKKulLV9fI16NJIRCidTJrN4t6k9cubnidy8VrWo6J1co4P+o+rFs
cJkV1/aYYcpxEO1mxmydWnsDcJMCfayaT0LVNoRaDP9xUnLBW3wOJnR7UsPI+Vyy
XVm+1CoPysJGuVm6W6HTZ2IMRfDmVkDKwzwSyN8eAzwfWmzZgukFgnbMJpzbMSo9
Vz8iVrdkMjG13y1lW+RHmkbv7tKFV60BGrLCIbvwbOVkTh1E01tldHcv82SoTekN
ck4T/0+c4tX3eLEKHnj0KXEsF0jiVVoAUlrp89lRK8ZdCGDl26wOyamv+DUWOOyu
bem6lRYQciRV/7o340ZvdL5Zy6wRT5PVi6c+OmQU42G0xsdkpsRizAYfJPS/Cfds
WEQBHxoAOAu/qAJievrD8hdOdaY414dDV13Nb8KrZV8Io1vWwkuqc1c4VEw/jGKA
5YX6ZeAGKgV2fK5PKxI/Me42uPBvPyaAmgwxQRsAUsIet7dKSRvPPwXxnejhMNVo
UqqytCZgx8pCMVnPor55wr2mqdgsNnrH3ToRJalB4FmD7BC+wSlZcReqqzYh/fFf
5ZvjXC5FB42GyCeNRSG9CvQEpFDpHX34sP2bnvLiCB3BzjXGvunLmIqxgHa60/q/
ljIYjMlL6LLmv4QB/eycUxM1k6br+QyFKM2ebHMBN3KarY5mJMS7IrbVhwJYtZuh
5UVBZBHtO/tzo/p0Or0SHscTOC2USdqsc0STEbM0QlJEe1EphPMkq/w5514RnMAf
xHSWPdzsLh6vrWzsizmVclC2yktV/UvxK5ypyzV1u4zR7Szdl6twotvOpJ6YdnhA
zuhTDrWDTky4VbxNtmAqWKosIcfgbahoxJRq1eN1JV+LJIBfOUwq73nlOxzrUv97
l0x4UjuRRGu4wS88QtJtS9+gRS9xtYAhXzxjdTo6ICV0e7PtpDeDKBaQCFmopu0o
WQcSw7W+i0ovz6jHF+StSwAt1KX7slwvPoINcSlT4SheBrNVJPdybNAuIQIWMKJy
fZgNPaP5/74e3+5YODBdncUwT4Ogw7PWDk9js3NO5UdUcNre+IpKYFkjU3kOSHxe
9hnjugGtj4kcVF14f55ELdW1k9zpu/Qs775qbaHjR1pFsq7lMhz6Jm+1Dwq1Q+qe
DL+QybH9RDNgjjg1WM8TWoytxiWH5GdG2zKvPzryDj8DF9hL0N1lwmPE8/nFs2eK
61lYIoF385y06vxCsvF7B5exvuPnPyKXDRccf5aHJmT9WdSujD1Bryz/jEJZ33rv
4kfY1N1vEr/HVCUSFR55pQCvSSjCnksLVygCvKfIQEMfNu6b1n/fPHgyXpUmja52
qaEq8cWqUALgkZna29NJT0mEXacajo/RkdzkFdhxOxg9XjdhR8531Eih2Mfuh9WC
sZZEVcsU27EK66Dm9NwFGlBSV86DZLJfvrBPfgGRzz2dskCnB6XKknHaaUkODcla
xWATaoqteKY1mHSjFhTrIY/IH+JwABXyps9KIaPzeZvlSrYb8aVcDUahFimPI6LD
ZQhf9wroR3Eh5kX2NYwWnyIE6OjZlV10mCuw0Qa0RUeYKVfE1daWTmkJBEL1OYSd
B0ipw09iVRpY8EcALwsLHBrUIO6+rFq4CXojeVZnlR7dp9IdhpgsFz7Vf57Tx6yW
ROCNtiTrMfiAuKgRpFU5oH2UiT8YpD9aQ7szG0qCJGHnvHMgpGgqVRSs8EggBR+M
Ebi9EF0SrnSOjB0zP8f3V4dztkA5imxzWxrV904ZQx99YvemV9LrquYGuCwWNWwL
NPDAmoN8CaVCDHyxUhM31k/K7rmJrylBhp2+GeYl2tat+zvBknG1LIbDraGpjwDh
vy2U03IvZvRymJMNASZL0KwZslIpNb09vHq2cznQ+IvXjwtZY9g+cLg50jDQ5A14
VSz1X96Q55329q+FTYQ7L5S0U0L/GUB3QxYMM6mvD477qFT4zerPAu1uk11VlBzb
9bC6QXZ9iJ0UzKm8pLs1bRXdYg9Alt2rjIKMl3WgGH8wIAZPyrDvoYAKTxSlpnC8
bQszRPSfOJZYJDG5fzArU5rC0tbcTH6BaXR3qNKS4nZDT/+CzyityXdyJu5WncWB
uHzC2y2lLjKK91up9WfzgxBz7KUQVibzMat8kDw2nDQAKZlFe6p2nJLHGNtWMNxL
+46zu4eA1fJY931Kr2Lgw1G2SMiv3Kxb4H/Vgmj7YzVlOc52xaipHefAg8qs9W7g
gwG3UqhSRu6bWXQ70zdEuyPpbaFVCIsl04oeuvapBgP4kJF791/zAXAYbU9l8uto
5OQILsrX/a1K9BbOyObS3L0wVnInGx61jQ82MqP8M034dfF35M9g8K1CDWp5cd51
RorpIcw4gpvXg6yuHDbaNBErGvHT7gy/WOSeB/KS4V7zbqp+tbEHtxhdum4Th70A
v9h0L6LcDDWeVZDLNJi6wz4iS6qeLyBRbK+tMg6La0uuif8okzgJOk9tSDs0bD4S
7xyx4u43QNfrl+meQM0V7LaeCJQcPKviGrmuS5+9rNm3hK9qSAgkQFyfiwxUjZpM
CHRfcTD3dg1qrhl9mUCLTg+7qgRNgk0bwGd+SuULWT0s6zq2OXjly94BDZ0tDkrI
gbDoEAavKaR7YCtyXi43QLKnONKJUtdsF8YJ8xh1NpmcuTy7vQwvkOhxf0LmFjmf
DfrkO8EvVlrylpZFZfzrzNKoKyXiGn+LhiS8VQ64mxOpXsdIe/nxv5rH3dNeGgIy
vFEI8e5mpoIJ3bC/7xtJhMg4ZCg/rD1+kGbGOkfyDNKkktzCMgsyEnjp0ZG25WO6
+injPdlMWRQFow/qj18Fav4jiLK8BLfAqT6WtXkk1+7mJMMXmRXzoAvjt2Ueb4Lv
hwYaENniAQaVFe5Bv9AwSoRgtKHDFn0dcd35Wkf9GVUfD2eYuJGeB2mln3BLDoF+
bG50Juj60oJv0h5KbmDcqYsL2ZxijO+vpVoVZJTH7uwGwLVG/Mh4BOhyFVJY1ZwY
PiV7i45i4QYD4s7QiWXfmIvSIFTjiwEUjzXUpBxfUEM7+j4datr9BREGLmZo+sSG
HgPO+m4A/uaoooqqslux/qx2W62icLZ+cvq0IeAUPgGxQazK2wwSqyUBoAqFZcV5
SgEQ9+LfBoXGcHZ70p8akZPJ7/BKSlflElK8uWQgzD1nlfvArdZ5fD6ZqOlJiQPj
SpPfilbYcb4bvUwQeneyO/mev4NW8mG46KjXFw/3GBvTE9O7c2TeNPypQZ6gdGAX
dfQ49JvZv/BwzuvnqmjMicW6ZST+vdbeaWSnS/zjKTr9tNE0M4dka4RhQj+swYiu
+o/X+d7K3MLn8ezxkMGtcC4m/ko4uJt05RSW6DCWCxH9fPc2xMXUAxgRNDsqm1Fv
AE+b1hbIRNNeOw8J9Fqu/yRz8NJ3rfNzYER0hGFysBf+ZcWaJCUIVtAvUQU0OP+y
CZx/tC5jT8fwfCMffox95gnzlexFPEppzH6uG+bhBzwHEiKSk9qJ2h3c9YnGLdri
MwMGea4EVoxTz1MoNvt4dW3obS467wOOVABgkFgE0Fry90GmUTxMIgpIQvkJsgUq
V42TDaF1E/7MxYf4K0gcuvWbK+h0ba0C6InITNLTY71wTCyTZYYhMYFQuZLOBXMi
9fNtEWj9womHZPLIfr5VitnLKLHwhE/tLY/7mNgDEwzZZyczkC1Na9UD7FmVpnFz
V+GZZqrsizu10kVHdSDnhjtP8v0CkLL7XTbzoVzrmPGy7wfFObTnOBhLj3esql3j
xspgRG9PqIZAsniRAFHlvcHNYNIo7wOAYuWd/C2xe4gvU4qA3On/67G9XujCLVLV
SfcZH5n0N3lAmzlTT5GaAxp1dhnra31nTq7lzsC2gMlmJBrD5udr189XgbGOqE9R
utx7PfwGRN1cY5gEN/qHDzpLWfNYytgsrCvJpC7lCYB3Sa2FqV7/zcvOfnJTf3Jz
RDPKcmKoWByS8Q3Z0zqRsHazv5+N2gAC9nsnreJkOYgr0GL/pwp0t96m5S7P3AcR
MRemMJCK/XeUIW1xS6stX+S4SjHCMkyRuqQ0vMTB0ZIX6desBUCrSH6ep9Y5+iAc
ZCmPjPUiZ6GvSQWDWv/9Ly2zC5BvHP+f3XUJmnYGOpjnSjLqN9Iu31LR0sZd4OQ/
0SLHY19Bs6Dzm40XCKCj8UtN9mt/lYMMDgjbKJDVgHwA+Nq2SyRauAwEr52tSJZQ
Eb2IcIWLkvrSdHSn4tGNP4tjpsa3mi5Xa2ONjDGMaOxAqBzz9ieOPdQ+TG9+8RBo
yhfDKJSHWdyKjJLKmDka4Kj3rTENnPDZr3zOFNITIFDh2+O9LnTUzY1pw5iKR0Ju
InDRz1AnPrhajt60qXWXobrK/GkuWBHhQ6hy+bEFqojcGNtTUbkhRJceR+QaZ8Gz
vayFGl6MFYGF+x6CFE7RwNRBRGqkTM8BxVG4NllC6FEkpChzZ8M8PT/84xoUfh5/
vp7PiuZGJK8bZCFwcMG+MkYIRFEocuoJy/p2tbcfsVk1fmQPT584VGIfvDiSFwOm
kS35u5ZSNR+jzIFq7VrWahrofRWdiGKAiRC9UvOxYjulB/uf1ZPgkSrBDVsRJYSJ
+BUTrPSzQ6ZpO2ziTUWrt6XoG/slOShYBunGf8IaAc1Da1Oy46sSyUfNkq5wufhp
WMf91vXqgypATv502fSSYEvQSOnziYf0LQS6LAsZoVHJUQm+7CGoeYCELlQmdDfI
/IDN2xbsuzIuEFQmrSUlPaqF3GEtZRtQaIUi9OafcCTHDkafzeravst+QI3nWT2a
w9RpAAT4GAysv/pYLi7PDnTz3ahqYR4av1QDF5M6taFEGmGynmXaeFGMz4RGxSNA
z3jBcEzSbm28uXcwSv2FMomfbnZT9RLvJtM08tBtPoI+nrb6qp3zgxBLfEGoF4eV
mjj5jHSXUekJ2Xi5QcwUSSuOxL6PK0Po0zEeXGdVCSkcYH71VpqjsnGsUCFJ7UZn
8YWinYHzIi/iX16T97wiyuDI6ghk0WHnnZY6/xCtJvONhNaWN5ENU/NX5xr6QVfb
39SSDjYWvQYgvJVOn/DiE9S8LcBHFE3Zswqwpt0jDHCQN0raweoH1qXclXFzqJem
x7Gf/Ykct0RtrQTq+ENQOrCRhoEgoAjD6PB0LQcYbktiOIWfWl4qKce4FeGKCejb
nVwvggBQ35hpXn7ngoivL85rRfadV3jSaRw4q38fnhvIYytbPrOKhB9Fvw2Uqgv7
NN1OsP5HjYWFozjOFt/2o1RM08q33cGFjyu6LOl4GxgVRaY3mE1YOHFQ4Mk5RU8D
77sGT4F7Hh6sAHkbWU2p6YCPrbmw2RG1BSMd9kYcREqeohigfvDOjsL23+5R6MDR
j0BCZWZwH4caFU5cdYsc/Sj18fYRqT2tgN5sJTHIqWOH+rSe/yIvz5QkmK7nV6op
anP/Dtv/rzyd4oWsaiL0m/8X+4CSZjVR0wUatFHVzxU5c4+Ti2l30eQ8KX35N4Db
M+UiED/j8MjNmNa4s1O4G9Y70mG81inHn0+KmJ4dbYVEUmmHfL8j/zc1E2lSrFHk
ffBxxxoBXtEGtNZuc+8C+usE02Ygz6NPNZXPqW/2oWpgVJcDeOvgp+U6rMnJ5r80
5g64KNqXKz8ORBBER3UjgrTAn4On/hCK90MQozfQz4rYHQ4emaRxzouS3APlEQXP
SVC8tja2dGsPPPpfOPabbbg6BSmXYaATT6l41sVU7t3SEWCwGfyFIl0uwOgqQ/Az
lCtjGBc85g8aWnWmoSZzJDi33lPrLX3+VSMz94JIqp1BIUiYV3dBxZd7BoyWkBo7
1fd2Dwj3oCb6Zpgak9aZO1HRhcdlS8sOpPQl9D3SyZyAppQJaO8X8bP0hp6IWreG
jIJDz3/mGeH8A1I4w5KsTCz/lGvUewdECuA/5YZnVsXalnYl2yzadxQC52mRx78x
cDM0IVR394aJOLXDhbEfzmt3Al3VsbUKuMA+OIwt3xCBJ313PRGELahxEFr3OCUN
lE0jKdhZmYvTU1uuTEIn0YheQqUXaQUVoZBmFbVOoTb46VjoPb5dumrpHqdeLOwB
p8QDEXMb0mvSgVBNwy2jbtZoQPaS3gKK8dPQnlISivOyWj/LFuD1DPGI/AMY2CYt
fwDdIF5ifThGrgfv7/1iej/92O9EU+kdQdvlc/551ntS4E/lrLCba6YUUqKsrHb0
wj6FQaZS5WAbLWtJX2jJXeBieHwHSNMYW14rI2wyal1q5kG+V1Ip1sGMGdRShd0x
DHO6uMezEE16DkaKHGORti27SOgY0EVjyZDVcZX3sqsjc5gxAXlt2w9Sj36f7lTH
vzx40nE9mNrrUUjp3/Le0ShI16n+hlXixCOmNT3NcCm6UAHa0hxN6xGMEiEaWkRq
gYDszt9y8rh5UEbNNSF014zaA8VUu8BQGBIsv67p7Ct/nB9OfB0iMzEnH//F74vl
ZVs4i54kdOypG1QpzzUKJonfgYwODjKC3Jn4YzR9DnOaU1iRJF68QvaFzA0t9hB/
1IpsdXi3Fz8nivW2YjotcihC6O7JGqBSmSbmEJ+72UBDPN3gVj5ZbvBNsQ0Mzfyu
z2Vj08tvHbOlxvGWFd77S7iG4ALuVQqtSs2V5jimVN0FLFq3CtF8dqMeaGTvTyso
MNmyLYrLVRaWN7/Cw+Gx4NUkbNmuF2Q4/nh/9Jv/rGAT7pBANywCv0cU+vVRPhtn
MywUxJW/iDUQeakh/HSnCoemNI3tB7vrPcvpaeyM8F13wmLM3aV6HZsqsqgOavc5
iGIDXp9MMsxu0ZXPufxpD1oMaMD3i7djnH+6AVTQop3sfeDxXPpvkT2+3nsqdeBk
qhS53cAxmG+Z2f8TaNuggnsgMFX36Ij7rBhwr4LMr6SEuxwCgiNSe4JuRtDhMVBk
BP4MvgqgTSax3RpzpTUBXAmckJA9J4rBOFTx4zp9YchBXitruF85k7xekRDI7Y8j
OKHibQiRPS2OSAu0e1whyJkCdVevTI+k58kxEJMIhPqs23rWeUv0drjZ2mhrGTv9
o1AbKw/NdPpM5XwGWORhzawVoNmwrb+B2Mtipwiku8UiSy76ssukFfkef1Ochn+G
j2sCiSjAH9/GOKuP98g36mGF2x/J1jo/P8sZJtgjbfQpdCrhoOQADBFtyj6i+fQ9
Gcz2pW02v11uLjXAzWmb7bqrARXxnEVkZC+Fv0bHoZhLlP+fuendbVJMi78QAuiJ
McckdQgXu5jtt/ZcEbjAuFncJIY69aIZlUe4gNUA4GIfA3YnagGUNJoR6AH1UcA4
Sb1elFnVBqevA8FFgINYUwrWzvO9M6TFbwlc2/rCDAvMCTUfg9GJLvIOMPR0osvu
zuDElCjDk+nX+7v1iTLKBhnrN6Vqg8f84JKmrcsaqxUK6biFatOqU7xLA2LgH7uD
LDdALXxr7AmH5HDeevOl8kx0gom8B4vs+l9akTHLmtmqac3azXhWr61G8Cbxj7Cd
kR/+Vzy+izrCspig8ekmbHgC4Wzbx3MMb5KlaxE3LNwkQoFE9UZnhT+ku8iCcyCO
RMd2mqpMVX38n/8Y4EQt/IcQA5ix0QudBLad5X1B0rA1+9miL6FTO3hZYUn+1jcc
X/746E23TmbFtjeIopGgfBhFEDBCaYVYs1aI7ilTIEB0bKoFaQe/xeTsqcB0m7Gn
BXXqAAQqSjCIghuRNHILtGfY0M71m/Cf1z1VAuHWFcv/BY4Gy0QOaPy0m11OOLHJ
ZjVUSeuu4M2/Nkwg1HvDrF6HhNJVYNVBFFIp/WpZpBwQndwE8eO6nfFax/UkQqBG
yylsA8HP3hmMzKTC+I+JiPD2kKNAlKtdoLIy5nEKYXy+LV62mqb755EVlzc+H55R
Ed+5a0fg/TiWgxGS+ALdQM2UKdqSiyWM3Y19053gGPOorZoYUTsEpH1zJh3JJ3PA
81mtXVL5sl2YXmGTbyvEkI76x0giF2clqFaK1eLu12qhA6e20oHlk7DDsbWMyCGs
WJxcMON1Brhlu3tkFgoL98ly0Sb2yOrkX0wwcueGUs7LyIXQX8hX34WhIT9t2LGG
dhtdyDln+S52pPuxGABEf2yptvs85ZpemaCRH6Ofewi8OkL3/3LAQE0upPckgi83
MHbOJEm6g5R9jonJ3n+DPm9TqoIo1r8F+sTCoUA+epHThonG1zw+L24kNLf38E8G
Y2JlYkP58b4B5Cx9Ay57wq8zMDZRoFS2XjnNe7An7nqeKXW3fRHrP1xpXSlaW6Ws
FuYcJlKJOV4ae9iVzQC8RsVu4tpiEsTkTHVccbNslAdke3t1695E2EwXjidZaKpD
TzPuZQZXcwK7Z1icgVmoQ39wvt5p9R+E/5RcX/O3wrRqi0y5cua0Rgd+qGST6ZaI
ho6wBxR8bvvmH/NHxLz7pV6ds7h/SKuacpafjt/T1uazmRqNo46uMpPVhcn6xvqm
T8T9L7H5TPOi0xjS3570bjm2yBqZ6ucyMh5KokBcBc47IZAuPhGyMuWibB8JNT9o
4FNy/Yhj0mT5+nmRnJgsIdUZUAK7U6M+F5Ffm4UFfM+Aa3e2l/qGrVAH7UtndUqB
pjTt0fmJ41EkJQmJpcYbieqyON5/Sab4dlcr6RU/e0IYNPzlROdnY6BzOnB9ezGp
OIraeaf9QqoyYYV974UTbMnSukLIFj3xp3bM5VJoMj486EVhL2vNrrTdVGyEdijV
dY7lpb+C48gmr3BuOPLePavKQ69QLQHaZ50G9REVI/VxmUJcrhMv6meBQgd9nbNF
ojJgT7Dj0IUYOY8FmGZ0eefYGaERYjDubryEf4rMQ3eZQs+xwQgWUQJQp5yuTIh2
y8wI1FzlhpuftGZrYFgQoM15eRw6YmJhKjUFY6EFV5U+kvcJt/ljT8TQY2TTZPfn
c1ropgHC8RigT9LTfGmR7ziLeovAAm0vrP8ou575s+tz5VXdLhk2FvEtoFkw9oNV
0XxXwiXuQUdNQbkP3ndyeCNNe7bunnJdSB+9YOCEtptlwgObkMEoOFJB5BscFQaP
f2jl+n03lFZP2WA36oIiCuH7kfSmfg4U6GMzHT4pd4RT8Li3vWNJfVdbO//o0yQD
IJ+yt1hIRx0oCa8xThuX0y81NjlWA/QTgFTcOe0S2a8wS+D9b2HOEafmWl+/WzHh
jMGNQt+y3Es4QnS8gzCSXDCMI/M114DThcYoQYRNt6whWTVLBtKULkcNLHgATKTM
p8z3VRnEpcqBPKwz/ofjHp/Z1owE8gJU2YuNgRY/4L1iVxIL+aLX5DpkX0Kn5EM8
7mg2Zv0TljePQJU5OmgE0pWyw99fzkVdHrD/3dPhGL2/LtYSvd1ZOifoe9wyM69y
BJVYGIOYJtDLIKJQ2jZSu22bdkMkqo+H3I1ToH/Mw2RCW8V1pVIPffHwi3WzIetJ
o3u4SdGkkGY0sU9vlbXZyqfwQOuC4IPVQlVzQClaJWnKTp/xVzWuo3Qsf6WxVbzr
dF5Bhl0oiOyqLAUieqvlgcMoldtWi94CdEomOqId1cN8PClnBsEFNnnSijvmueYv
GIsErj9FtlEdnfjhU6JPRb4wdzWoc26NX6tPoDIcq3ktdR1pis4+QFe8UsUCwTQF
3KuXQk157TdB9dBDutNZe/i874DxjbyI260FWPlM3/e1CGEUfM7AV2F0LVHBEoME
lXksNLyMA6y1LMQxJHEMH4VM686ed/BTQkQatY8uZq9MpUdfrfh0pUEWFd+Nm7bl
mBdJVloZI1waUQ2obCQPvY1eXmpLiAQMy92lwPHZaxs7IUNsBNWetZJGYlYsnbpC
Ezb9RiLzAIvNVP/mXnY6t+VYd3YfET22cqmNZJTgYHBPbYAdunoKH4gF9swwkWbV
s0I3XaK6YBIJb3XdZvoeyhA+gsMiaNh9mtbzwK91dSFuen1vd7VnfclFU/AydJkz
GBfvosSl3s6WueBkHUpXDC6Chj+N2pIq6CZu54sO9MguwH6c0fxbMWdQoC/h9jNT
o1nZn7UU9c3/aoDbHWawIwsbNOgsohX48TYGRG4yRBPY7+AT3bj7MdjAUqnq6p+7
4POAgLVYIMEDPphjbxl1foj2w3EDIftCEk2lDf5dX+TzVKnHlxxi2ZtqGleCV5va
neff0QNp3qqVEY3We+gbmGAvYUjHwxxqiRkpqpV9R2TNpRQIvPVa0cFGl668axVQ
qwD4TlV0avhm7SYQpszIB0YsvtXR0+gUYhh0GHh8Vie890V58h6+2mpR6Oh8m7tD
tTZISCHZ1n0idbMrPurWst8h6VkmTaScy+V4Tf1lysjn9WDTO/FNWDz13WKW/B/b
CRYg509QP+lxf4tuyy0NmOfWItE91WEryIUa5dv0KPglilnzZ4CuAZkIvhfyIAvk
TJqblESIwW8FPOIx0jrjMxEhaml1PNlHkNRcFkzXSkV/ia2MftO433unCfZYxVBw
AubNccHJAXtUN7LfNECBa9g0tTm7givo5CCObHqV1Ks156DzI7onT+aDyy/OUNIN
CRkItGSd6exZduWgqhdjyXRpQhwWSrPM4DoyGJ/qr8d2HW+zwkyIumQbJb6iaKsx
5QwjLMja5CKtdC3jFg4LhtU9ss9Se5KvIoxWRcGJ9ciYz1oOBQk7i3p+WpkFZ30P
izoZLG420XHree61j7QsMaXqagu3HPotdROVzp8UhWTO5QFdW5mt5ZKwRhf8jOAF
WedRBiVwDUwxnscGkWiAr5KKEf1HQRlk8MzhbKOBTD0vBAaqRuo3SOLhpbOdtc0t
2atdeVg8zblc9CdwrrR80YrKOC6L7glY9+SHX7xjiGQW6C2Iva6eSHJokhBT6Tyg
kAYoi8uN+NJbM2aSwyRHo73CdXqNPB/9/n3TqARuwueXio7p6F5tQFeV52VU62pf
SXL3cXXmbOnrhzvNmvYHGrbo/afPLAQwHKKKfdhMhyWGv8+fm6vGGbJqckYfL38W
mc7PcFysR45UhnVVRFICFCsb4Av6KjiFOZU8OkSmJ7ZKwO8FxdIivAD6f0BKW7MW
bjNRFvnF138msCYVzzkiJAQiqd8ABhupIXavmq8FZN9OHeljl5YCaVSV4vIBK+zk
4WRGSd519KVvY9EFbMeXPui38l+T2LROFAI36TwUjKIQegpnRcY6Dk3sm36XwTPY
Gfi3eFSTdeZEGcDxHVu3cTLNH5wGn7sIXYo1o0nsN1xqGvOn7bSY83GgUQH25pTT
LLcIsFG+hw7Uta+vSATwkT+YOrD6Jqvu3nA1fNBYFFlNEVlJYs1Cu+87Rq8gYuQ8
VK2HYLNFDEZrH3J9wZKlA+EoS40KzAtauEunzoBqd/e3eXqP7SC+fAfGfTDA6tFT
UvOCNWNDgw4VOwqsKxuxlYXMbGGcySmDIsSz6ZHRmfoXSeRetHp7qoke66g4qQHu
UXIAdGw4hGiX1FomuhdSAO3mIQ23/+sA3mZkP5NjWgHy47gdwpoYsBB+mqLWvKG3
WCq4kDCeuDvfLY+y98ez5GBM9O+tGDQ8HJKQvYkCT1GRwiQoDZOBeR1cTe0wcvAu
ylNNvl17cefDt5Wg4dWF/HCANnok3d1OWrdoy1gWcXNbtTfFFTUkZAzGPzgdEcAJ
JyXdmrognqVoX6gOqHkl1iKYrOmHNVMwpsvHGmsDUCvrsOcZt1EBCrDJieLyd647
kWQc2FREkeKx52ODuYIRiyaqzmkRHKCUzFkUBozJZXty9MIUhFXK9txHYOyaSdaw
9Kyyw4ckyr2TlKXXhBbgAAGwL3HWoyJ6lpRf7XCTTq+5zUJOZam3jxftlfnKUuZb
lLXnvwjkr9mVDbD+4Hlg+HJWanytK49J77/WqkCQ7HXjLgZbsGQ84MSFBKtdRUIj
eESqfWfTVFX0e2HcsrbPvVOSRRk4qUee1eJnE0b6qNTMe54+e90JyqDZIGH1WV34
wNiHGhRmmZz/zxwwdBWSHAbBuEgguojKxOUAlKJCj8g+KXRhxdCxlGJeT5cHpZ2y
I+5zmTsYdQeOnxCQnl4m84bCMXDYY5LRbLzXiAbEMVBsOGd6IaLsKyQ+kawsRnn6
MgHYnirQie6kgCoD9gK6UT8IH3OCq0NNzbvUhsIG4ICfbLTIGxnS0PuF+e57xQHP
FxMNwXxu8HCxSpKiagZJLSTEPwQc0HC5DvCmkc4LQC8qeEWNukpCN+SQaWzcZfEJ
G8vxCyDdMOQdfhgXraYAWp1YlLBZCK3XOJ1PqpC805RImHqHjl3WURid1+Uj82Di
BOrNCSHMnvYx534ysPxFlwMjZSNHdYsF5geIeefW9bsAKL1tOIhgpAb1NHG1YZRy
WzW/nmJs+QAVok+XErTlmh3tezTPLE46OJydbPZPAtMon0ydqowBVadR34uCiPeo
/1gvjUP+UpevxLRzmIa0+xy6bCQqB0aUTCYkYaPwf7U+dhKjKcC20K8peaqtVf5r
dA8SrwUUzuEfrs/wyV+HehIx8nEDKYju2o9XNQ2qH9MIx75my2+GoCzcxnfXr7qK
ZMtP8TayH+h0WG7ypW71bDdkdgB3w47eV1YBICFEYEydBTZC3THS/d8Hx+WJaOrN
GI2hfujxB+r9C1XVliVAoYxwh1ceAe+Wodks9zhpkJTjBqLbTi26KJIVSUo6RqWD
B7OyihkZ1ix+op8JJojxrHGj3HjOGeW8L4DggH+6CNt2BJEOcZ/UyBVMtvRFO4NB
LCYlyCeJKRPlmAV1InbkcmZF+BFCceCf3gIKLXSPfkKD9q/bartQbjXah+ZRO/x/
sj+ttIaNcwpOMRduQV+iPCcq+M1CVrHINoeTw/ZtryEnSMGt5aJ/uYvG/g4CGnXo
edSzjdPSFH6ywI7ETpUo9OuZ07yXFs3Erprxg0oxCe4Pehuo530Z7BeHdKnFJbGf
UqCCADgrHJUxQ7OOkmLI5IeGNUfCIKQ9F/vHtmM4vMaClUf0Zhu0C27GpWnxmubQ
4TrM07vzayOQkSLNQXRp/Xe3fCUY2zXwVcI/Ss0JEYVSnu2uDwl75rfQZkpg3PMr
qKu72XgISi6DAlk0TtYRvONLNzOx4AHJaMTG3WRiKlk1lUU7oqX8NH6kF6CLp+PH
ZG/0s3ve9A9VKdSY6jwzCjzzHchovRn+M4PfOuHaVETTqyI1dggkb6/4A01V0fUE
5Wcj0Jk1XC52D4kcLR6r1otSikztIK84MuJnw0td2qyKHnzZcdp/EsurZzHsoxUE
SK+goPV1RUl6FolaPI4u9K0+zzKc3SyVlpq/FupmlMql4Ka/RHr0NZ/zWadYHHuJ
gWp6aLskJ+ln4xYVlx/B/HiReIGU3Ib3xqCju2IANpKh0aywFSCKXQL/ej3pLsd9
H507cpHc3CdPuApoV8qwcB4GjPSuVs4UuYlm6DA6ihHuJdOQYVGevsJqlgPF0NaT
FgmYjbjZOSoMC0oOwOkeBDdKs2Rty0/T/DYLKdUnjOEGgrgV+3pJXLJ2TIWsXxfE
+tFzAbDhT/oeRE42xgsLimaNJ7FqEfZdtJr60IhXWRL+4DxdYJssb3pEB8QXBhSD
IMGmDKHIHw9U+EfYu5qqAj1cz9TcgKnYwRyb1JkGC9X+G5TxFLt/d5w7oqaM4cms
HW52NdZK1MKKLTcbON86ovM+V93QiTBphmtA6JLGxv3HLHLxhinDludcRE3uAxYF
XZOtJm0PWw0yejCV8zLHSmVR7rILo6gCTxBMOBNQ0qHqdwGAuqrnc/oPbgsZtz6V
biI3Ug2pdy8HaRzNz4GDHDAXnby+fQlW/RMdcRQD8GQxIRIRqsIt8wm7T9X/Incv
0Y8GUg0iLvbywzxY8IW8w+4dBobEbmtO55qt7aqcRolbWi2LxFONs4WLK17V9z1G
4AMuSDLdzBu0dBTaOV7PNt5F+psmcfYGQmW7Hr68uflaQVRQRh0/omSTBQkVp728
oehdQNu18dKRfy2VNOlXVqowYShG/vHJZC6lK4DmfYgKnKsNddd5KwfcYKwg1qaV
qrHo+GHXepGfvNYatCLt38ZhGcbjS2fq1p9uaEjD08ySOuFZol8Uy+gu3sFEB3r/
Ypn51gfwtUu0AsXlX4TdiEmcszxmlnXZuRqbddQrYVIsaRgc3zrSbxFbUrXbkyrU
+G3W2QSakmFMGNW4CzFRRqywRMWkkhCOhF8irdgN+yyLXlI957wl40qawnKCiLm5
fSGe8NTGsqKH/iTZuqE2IGVETTXGOWswfoFHpmta7lmmoEpVUYZHz8BE/hjw5vHw
6N9m6zo1li0Sz0njFdflChJoSB53grPrvptTF0kVaR1szaZQXrNWJScH5xR5DYRX
MB0Lf77eiS2IhXScNdsYPQDa+LiAObmWBVbHNDZYhHHydwCeJsDYOl4VmzXKBD0f
aFzJtFqIyp1bFAYG/H0tQ/UJNcbexhQKdYl8TPhit3IPidbB4GrI3esSB1Su51bI
ktaEniRrwvMciL4JZv2arqyTNSOkYmqtmCyMSpmYISkXK1Mh+DWXs4IaHvKqerZ0
tFQohWKpnKZKV4wYHKPtreYmiOhXlu7v9S4B5VkpVsBIjCUOUIwinMerZaKMtVlq
9FpwnR5f2pXOnwRmMEejG10WUqOcnvCBv6mR7QZu5DaOw6U/NHsrC4WiW8BHEZgr
/K9A7FlM69D8BIk/ESH4EIgbUVQLueN/ozzfXzt8L4RozVOQ9aOzA2hGDZb7oUbt
siOZs29BbQyFZmdZ35mf75fXnCgiraITnSDedMWUfiDqT83yCTrNu3qTTLTZKpJm
43YHT3IxyW4ij5c+3mNQt8Q9V/R5rDgyh93erXWGefXwczqjHujCGzWbn1JAmIVE
zx0SmeqMLl6IR84l5gyacTEVCxxYeQ2RC5fZ0ZUOyWnYQ+p3ovBFuWhTQGN2MRFt
2lhoyTgyjDXUL1hord8dFBxjLB8zqW51G996qfsuNtCIDp0/ozU6Rdwt1OUtbp0Q
axcKUJajoIj08HPOA+mE23s8nS/zRiJh7jg1N3RAoikV86A5WSEoDvE4FrtE8u96
Pglj729EeCl1TCgNizqb0jL8fy49FSyDBucP88MOtxkNJPY+BLVKef8EpKzh0QDK
cabQe5bQr54UFybvGGmq2dBse3XzeVj4QQBRCQ5MMXs4oM1gcAc2nSvOP6Q2Odij
K2yCCoUwbBV1dkGJqy4f9d8CNbOO13K3uRJ1K/qDeVfMvkg65ToXcx7zNFzFxcO7
n12wduQweH/jaSGgzErNVVodcRbodI8XB5fRzy+k1LamTNPChiHC8oXMlACYlIfq
PfeBrRf5NwVDgkBARgClupWmRA4TVmoGMNZYPC3OSr4Mg1o2lUIf+PiOdyRkqxPg
7iOFu+2wQ3sWGFtHrgZ+9aAR5eQjEBEAGz/hKq+bFn1xhkAGuO+hkPz6LkeMbGeZ
SlAwIQE+C7ZQAD7/PFfM5hrye+0vq/ZjmRkj8T7sExhG0XDgxnQl6Fhf6YmLxsE/
MH8p7V9BMImnb/aq7wtOD/OSUx5w9Wswua8ijo7q9ceSI6S0Qdx4M4ey4jx5H7xF
nTwflrGuqZG7taqcVvlPNPq2R8YcIi8X7SdL20Vt3lecWPJtZM3SerOBmI25th3t
Vi1mfDhD0hDtYXSsd+wAF7i/D2mNzTbvFHhRLWlzl3n2UFAkVNEVQ4Q+qVklhREO
g7TORGN2tNLlVIjeUdIYhJhvTHe9n9qsaX/aPyVBhTKNk7Kcjt8ByTVuAGBvea87
3bw1kitJzDqmSFTuWRLPwa/e4+BW8O28FajiYy7YDNq01VawX2NASirFehugj/T2
OaitYcr1C6x1FjDvArO6dz8YUpXOikSrcza5D3+pZEY1ea99lQAIcymL0qfxIzvt
SFBm8aMrh4JjT45nvMTI5UeiTA/InNacWhpcsSTOo7luXJLQgLHz+vb6yy102FPj
UyqeaPiKX+5l8ZGgM9Ac7gtplNsPlzarLc1KIffrpedAM7Z05dgk9ePobDnwjt53
k9f7/fF6BmU6STQln/VOBTG43/2+ThcevkAvBPxaRM4ggmbOYFF+wQlQvOqNJVHE
CE2fXrBUWWULoVYFg8AYlYODb84BhPw6WInLswJAAe49Bv+4cRw71CT/0f+hWbTY
ZKqKVFjKMgmqP3dh9ao6LbA7bX6aWTC7OqqOm8bv484iBk/m0OO4iRmTVc7nyDSz
PakX6GgAjnhYlwV5MPHprnOUxqozHFwQQ5nC06RMTty4WXiGTOHL1oySI5ESFA4r
SUlv6cZwNvinPBkfS/7vMqOIgAI0ca6uLKS6YqM6LeW/Edo7dD/gRL1tW8K57CCh
nygcU0LoEzfKsIvJhPtPWWAfNvjEGsCyKVrEZpG5rt7XjqEM60/pe1fpYmGsKkb5
d5kZPg5KvigqozBxJ/q/SiVdZVaaMoGskioOjVAGtttbS9KQgdtS/ySKeoLeEUdW
St1sz66Eu0vvyYXcoGpTmBxQr/2gw+PKx8txaUSV/YelGokoLKixh6Vj03edUeqQ
tfejJMDnOOZLUdutlVZZHVH36jdem/XvHW4RIHpk3QqN0NnSyeBW5f1QDeq4P9sY
ZtCSdbw5xLvQ4U03TfuWYDT3BrHEORpZM8zJXFsAEzimEeRTXNLm1zx0uLjmKjlT
1Du2pxp9g1Q5Oby05Ee9O7tYXbkPgMr9hRF3NRiuSyI/e4u6ajtErBQev2Y/U2mT
ILeFBHOe+gfc031I5FWgOI1/WjCq85dbKOL/aIl07MC5Jw6pWE9cF4qEYN3ys4O4
ygDz3nRysbQhr4QNy7WfUrSjipBoNJA2IFXB/bWt1bT2mNE00Fp7dUFaxgfUaJWK
cqY9ZBdvnAKAEBx9WeGVRDcfBzXBWAdXOIOkiDMqQ9JFBvZx7ZGl6mOHFuZqJcIK
7tjhnQGT9SHLXdrvvpTZUAGZHi7XIBizMQ3vWAmjmuozrPBFmRVM/TUrbccsjqll
OMhDJtb8psVcyCjsUhGOv4fEv4ohPYPmbwbygtCsX/8t2zO5hTD7b421WAfT6ktW
HTteVd1ZzhMIWnAJKM93FtsqnQOftW0w2fG7Kvhx8QECvRbf/ryY8yK5NTWRZqe7
3/8IbOr8RpmG+Xm5LTL8u37fnppORyoVkGGUkkt504Bo/P0cYB/iMNbDIQ6uYPiR
i3MoPE+BExrDfMYTfdxWHTECbKIcyXBywmeSmw2RxCh+EgBRvORDL2LzLeAMczn8
Q4f0IOTE8FsNi5tXm6JiQDRDuQXzFzJCAO+rg+A4qpMgU7U7/2S5eq4nwWRAwrzS
h/rk+6XvaFlKb0wUPLTj2XzxhUlr4J/tGPSgtAL6kM+bcRIfSlKLCHPHNKGkFKYY
c8lVaQ6J1JK2VTTfNZso1sJOJrM1xERPrCdKaW3GMmBQxti9XLEuf/aX65MjKlhx
Cks6ykaI9zSESHHeN2Pm4O+ZsyA0p3OjBn3p3EFMmUB5lJWlLcip/njFfsbEJTnA
pBeymBINhgvA4dFYu29I/AnMCH4TX+2lUWW847zxP883cRZ6P4pKQDVvJVAmHJvZ
YfR6JpXQMOD57WLb5d5c6QM1GWz8oSi4v2mG+xCAoLNnFJWxJ/tFBvW/BsO2xwvA
EBjgb2RPjH+cii8tpEHG0+cuKOm8Q2ebJhISdnxwqEj6t2cy4YAkZyO6NmQTGWv+
1wrlPqJBlFwjfATO4sCsFGc8IYb1fyfixRYC18HI77S2snQJyol4HzY/7l5XhR2L
/+wJ1o+SD6TcDefJA/NZ51qZScklgtd9jmjDMINah79LW+7WjxaHAjPvjKibkH4h
GT0fiumqki9RhFALP1B5aflLWk6cHEjIlXo8ocHC+U+xGAAStaLJPjR9m55jZG1j
MBDLa1L8mQCRqMttBJ63yI8VEhN/0NJz3Ow2bsC5YVfnqxUz0Qcku75/hC540Ot7
Y3evRzLmKWnnrN7FkFEX033kO6+JVihJ+Hzl4m+C5l2Rn/pmOEhDkPPOv8R4Ms/O
udZN2FScIGqptm00u2oYfiRnmWo1qgm7LC1Ai6BZb3LAwioth02lezGMfQECESEh
MXqJ+IBPmBeOStblzkeRSbvlr3Jj49mrdHpGDx+8U60EBbvnU2ITVQrRnOK6pXha
D7qiz4TwkLlnc3NKPzwdCG5FnpbvNUODHHHm+ZwQZSPNiDoemREbfaqjGH1NWgMD
5Ez9FQs109f8ZTnPYzf1tSCZ9AsftvWZ2I8snruPIXfxxg9oMrRWeT2hnjIcnio1
1qCT29Y+kpssuIEbTM8zEruWELb0UcPdPfwkcCkS4DQyjI+A1dbZnIfRXtdqs+Fd
1d/ujqfU8en01t9aq1AEfTogXazWnP9JVXDfKbyu0CGBUaxnFxtF2IKqPp45Dc47
t+NnV/mbWQT3DjZ+Rd1qc+EU8bREY2bFIqVJRw53HXmqWuiOugCUlm4ORbTF7ATa
TNfL/0Xw6bOt4m2aQJ7dp+wj+kidb6wwaUg3LrIZsMB9is/1F6fdfxiXOu1K9v2w
oUdpuUL8asE072zPjcF3xHShzS+1AXaFHNlZb3QUzHBd9VS2RA/D7JIckUS+4p4Y
mMFNPy+dpOt6ozOUHCUggkBqCeaVzk4LSHjmv2lNuSysxxeZCs9uvDey1QzCoIm4
9OWr4J9g8AfNvaf5i2B72mrc9r+W4QcT303Pie6/WpJ3ypItoICZb7EjRxv9KvVw
sv1mNLgT1w4msFRAq+ngvlv35EEvA40s2yfeYlAwtUhaBBWOtnGEILxc1lElE0D3
Q34MhzzUnCFI9uE20GTLzpaUWmyLxmzsz1hkpnCuCFAJ11pmG+PK/Iis5wACw+7y
BV48e+QfZtMiO88kWsYlgF8OQ4qXbpilbaiGVgEoz4E23q0fHD08YZpt4/EOfZNz
/3JQdjarMVKOXk57OrzhrQV9ZoCAK280FmnXVsB1XbPE6dKsrRa5AgVN3nkamNAW
NRPDcIvvAL6/ysP078VZgnZio9vZweCSkjqosVDektr5OMtkuqyCsO4BTgYSlJkf
lszRU23/FWPYnbZQmM5PIiIujN6/HlQL16ylCCiAKVMW1TkgqF6chKDrHtgVj+3x
ealrn0PMbHvNsp1qfmw3Lfrmm/8WL8aWz5bWyE9a2tadg2oVvHnXHgDHOxWtWjX7
4XxHvu+YC1/bs5SE/bM5ywIvZeamvQPq4/AjA7hqlLI0y+TYhn92PDnMoy32pn0N
v8AtslKQQbLCew6TLIoOe6do9yzPvgvPluNcu4s0I6VdTlvEGmq+ZX59fauDNPCE
eIkemwMPRV9LOtAcB36UsLwgosg8WxCJ8yN/lyrPRtVoUqYyGVIFl3ZRr6Ev/BCo
MFardPsOqu9Mdr9ntHJIdZiYVNG/fFSIG9tAZqPt9960+qW18uXFi59LeGkztrM7
ck/HjUojYqbE3//GprjOHPExGe8634W/xMdFNBfpLSTAFPFvXrOWB1eKrtGlbkda
coGSotxHnWlBsZCJPci/+fqsGRsHUgyLXorGQTN8k1nLvHClVFLHr52xOhGwVmnG
FVuIqkYI16G2gjHH6o+a44NxbCi9WtYdXJ7oROzKOSLNErV746NXqPs9N0N1Oo0t
KYgKG91vUiKzlYYcWc/JkHnscVv5PRe0w39nwgPgAQGPwJ9Pn4khz9v7CbBS5/96
aSsEJwpajgba54ost48Sz5Of0tx2yOl7l0B0AfvKCA4ykn/KwphN9CuUSG/hTdw6
RNt+H5MmVDr9sDGpt3BFoCaPMWK4O756gNfDUuYYBkg6MYM49ixWMKFJVGw/Dz5B
p5FkVOBidwUIO/Ci74U3iKY/HSpYZQgBtxVsxcz+uznGb+fdJ+wFmLcONDlFEgrT
X7Q0A45a+e14TfOK3aJzec9GJR2bh+hxqvfZ3YKJe/Wvx2BTmnZ3Bew/PHZJ7Adx
nJHXiV/c8+Mtaw9QTCumUoSWbmAEB9XBJ9ajN4UuMExfTojFEVHKFgZZv5qrLrDQ
a2JuxwPTdhzYSO3EBgMWjj+AD3zLxSWPPIhHxm/B5EvEjB7hLcCwJBZOXW4sMEoC
ruMSovBjVbmQX8IwJdLO1OR+dIJSNgw5KohBMfs3Asb1eJRXe/6Kit2N/gWhVaFS
NbH4YaI1ZLYD1F8aQ9mVT0r511ioMBfUL9E96QBvVwmp1+xwzB2x546+Z1AUs5lp
Wj98rKSRb5X3HWFebMyNY6D5fEjVZGe6faEfQCmEcs5eHT0hOmLWSxg/Od9hy4jG
HD/CYtOKjrp3nWjTjQe3SWF42QDWhyJsHOk79xYlYG7nb6SzFVDbPT4ezYiYYEEA
3a3Bx9FfV4bgKTWliYS7y7QJLhIuVtj5lVm5S2RV8ro2vgZKcawc7lXiUV0TspE6
GQg6fzaev2EzNiLMNunf+SGxYj83KXYRQ1c2suyYTXbpfGMpad2gfteb0q4kLCgW
0wh+dNHkXbtz33iDQ2mTcGFvV+3+YOhvIguLgSwCVfERjiyq9oxuhrJXK+nMum/t
fifYuYg2FpbFa20PmNoR8RQNJLcvKZMh0lL/iFJM7rHoABpBWbM46doYh74dIJVs
abH968Tl8qDpI4lr/HxznWGCwNbQo+2wr1v9BJRetHJE40rKQJi32T5HLXhEhefp
K3IgH1Rlm6BjjB8Yz3cA/GPdB8MXHjiZvp4NXW4zLLh3HMAAuU57akyr8ZmYk39S
svEB0k5Bha8IdJxdSYzSKd4iagrdTSDDCI3Q8Sne2Dp4WqVQD8ZcIRoqfHepqjXx
kKb7k2jq8BXxs5OfioW7I7Sx7q4k3cP81jxY+awI4QJq9UMFzP8hDT0cOyXtZIs3
n0OZhTKvk5rTazL2RjZbZeGcOGZ48gjjIpg8ZpROj7/GQrf/n5vDMetxnPnJbS+1
L2jTKIGQeW8XPdYPOihXtSFWqcjUEGiAhRKgG7yxjB/h1d1rf8MqYVd9VuKxuBe6
tSmfRehXfYtvp4WGB1CwYVrdBWJQtjhhGtXiVWeAjjmaBWhTnix1S8Keb5FBVZ9y
zqj0GI6xN9/QQv+IvGMTXSpNcCt7MsYeXu6ua+DWwmMDGAnIbEt+dFgNBNgzjZZJ
jMBWBNG5+hGdxjj9AMSoXP9PL/jco8hjnoYi2T1kEmaZDALy2wUP+RYkQXvf2YQc
JVoMyGQjvRD8TvsvVhXFi9rIS5wvY6R2ELL+aCQVttafQK4dxYMbZBJfWTK7AE8t
CPP+75omfdkiY9F1Ir159ui8C/+EN65zhioUfOdDM3BRx6UybFW5qGOi2zUTX+d8
hBSQ6Tkvj+58KCZ+l6SQ/mOyPJbkmD/UXaxptHIyQ0uHuHx3JrYyUDuBo7FyRxp9
pYgswf6PdRv/Vh9lNNbzwAiqEJ/YicrITYkMtmn6wlovdpnLkInhv/bylhbUJIqs
tTQ+lritCJJ6K89NjOvZLwaNCHhQEKQeJuTJBIneGNTuH50YtrFGD00MdvJx1Wnn
GwXn9ePmPODakCZu3maL0Dc5SwmvhC+jpgqGk66srzHYu5N95/zTy1b3R59YnG0a
aBqkLk+V7JQ9Ci8Scb/bIHLLwLdGt7WJsBhY93OpTuCntv3+EDRtTk09BeyQ3PRU
HqL9vbIgxfPELhYKHKAlgZr8iw2UVNvt4pyAmWv87C0j0+4kq4Zxhb8C6z/nt4wz
gqbuCk7R8LPseU92FQPTD9OYlZp1bp3DMCv4gaiz4zrfrIsxv0dY0I+cWeP3Yldy
BTUTraOdtPR1L3jsP+wkMDKmHp8R2UzI/9ghZPJTz8ReIA7avOR8kAGsreFfPp2S
HXa/5nA1VX5B3uUtgo1+MoL1ZRt8V2l298ZXl+UgkTu5zYM4dTOtm2tBamBJoJgL
Ooq7xSY0GqTk6T2AIY6czpQN54+0OElOaZj+dw8y427YzDkKDbY77bcLwMpRMbWk
3FPaEYhG9ZfT/TyRtF6OsVZDeghUIWnLIbN8AI/ngARDOViUFJJmzGb+ln1dsDD3
nB/tFQdsY76RxHOeT7DsFAF+Adz18WcL5KD2H0+hbDyHDNMWmAlEaih1Rz0U1/bM
3RAOnVdrdJiSZSIeCbEPHkdI2qy9daH1F66as+kUk10OyWQz2Z0y9tKiFso74ozQ
4F9ryxWSkeT0s5rzycO6Knyz6b0irIHsHS/P5rt68DPGVMU45hhFr4cRtmraRINA
W5+Vz5G/5P3CJFNw0TUnBVicFDFeOozoZ9mf/XZuxJ2Aq8PCUZiLT/pcjK3iVLzb
W9YdYrSAvm9hvgqqCSQccrI6e2R3cgqvYvpL0FoVI3MeRJOHH/Ase1IG7nmGCoXX
QnRFOmpZE+fF6H+MUK5zT5FYKFe4UHVg8KzzVPNwcnorF+yMlQcpug9X7ouS9vfk
BVlpljvQl9HkgqBSeDS2tdqLZS7PUyn4cmjCBNRZglWSeHr+AUWEIZlekPIPjFs8
Z6syKKdaLBw/CTSXKZ2Rws8ULzMHX+OjGqKQRKdIJCPeexClzSd5FnFcCj0vk/YT
OImAqnJtOl8EGaVxo2HyXefvWsPdNADN2QZ6bKHX2+xai6nnq5EPrbtgXPQgZHgI
Mc7jXv3QY82TcPGwgSA5PXEgJ6z29wJe8/uP4Wv+V/0UO26wzJJjPwpKp7KhIj+q
MhQkqsXJkuFDNK+Zq1rO1SGKyaMGrERWVOOIVXU0o0ew9ZhOZxcyWYmELcrMMh9L
DGXtr4zF8YhM6hhxXTkNPP3q5Ven1nN321PNlyUq58gz03m0E9szHeZxaD3XWXbv
eLR/UZwTF6/+53UkEpU1aX/TefafHoWY9MqZG+iUIyvB5SeRRI03y+aD6HLp85SA
Fe0OlP41WC5JmZCmsfADgxavNZfY141IOIB2+LFmoYMsfqe+VUs9YOL3G+10623w
8hMkRZgkySQ7b9gdwXf4zACa4XQYwfgWk8JHUXaG6Eo7veYLBtSQJf6gEN6m3IMw
ZD31ZR0yM5gB3VwOFTiNfyswLkNPvbJCeYdViuCMQQ2T5YXkXH2o1slxe8wQ/ozK
8h/FTDvC/rt8dO5eEhsD89K6bjZrYgARGHrUjBXFfs4zCBtCBQjaPQb2moq/Bg6x
0M7MMsNpzKL7//mHkbRDMzOqOcQI5RnoDeq05hEMkVAY6TqmaE+iHqVB4V2SSdtG
Y89YZqJHrYX1CGXb1ITvnLIzuo9dlaH3E2P4m35G5VKmfCMA9DK2pK1nnFpYbm5U
ITs66RKSvbmMK/RUvPNgUyDvIz5sUzjV8orD5EDkSvYxRDMNm5ZFzIDJjnpQHhwX
uRl2WM2yjofvh+8n1K2wnavZ925QlmMcWDrDKyWM76iXH1dyjjOtayJH0rV7cNnW
BMK/1ofGcPXEJQxHbHwIfLLU1T0USuR7mTHjv1N0F9g6NZlAt01BIr1bD5zIf3Bz
vHPKBj6ZFrFHTjjm9jZTIySs6v5FxcdQuJ9QIrXX4rzmVG1t0HaAW6osDH0KNOm+
GpkbTMbJGR6XH1t8bNXX/6fJAFUH2cVzMOQmK1ywK7SA0u9kZjPscl87Ce3Orspn
amiufcvd9p/9E5q5pQRajgPLZHpzyhMZEmaJSoWV7JUIHUvwfzhKdVdXBUutHQHH
yBF/lmee3sFZvCPA3+Ama4Uz6DIPsLNSLg7hO/Nkol7Ay7qTUTh2A3HceNV9y0DK
jn199068w1CNj+Q1N2Z5U3mUT39bBIrndIuIj7EmrxE8gFVVnk/QFW76UQj3wxNX
E5DcOEx4ExEA0uJeLfQoHZ99qrzMuU1fBiyY99r+b9oy4DAind9fp9vJe6KgXPci
LZWPP9NJys1PIizTqjj+TWmS7K/kYlg9jJVnYX0XV8YO3P8QnspyebssmKpfDGFg
ALfqnHOKHi/izyUBxnBEkumvQ2GVP2eyc8zQ9SgHXnbmy+G43+cham04UBkWA/pt
F0y/2lpyBELVduQRKKF8wOelLJLMGhOyH0Nw+qyWip3A4yn2pDsmDq+N60aO8/l4
y5meLPMA/s9/+9CA+JWkDGNMCxWTr8+EwyDLNbkHMnR2+5V9VgkStxD5Zw3KSwo3
rzfNxeNi4zv3jah2PoQbar/ulUL2kARBHhLidM1yFVdrZGJrEv3neCpNd6in9+nk
Yw2BHE/nrLzNgcymohktipUNkf0+7m/4Xu42+4QUu6UujpF2+cNN4hl6SlDmyzGV
NVUhDnn80TQBUOOguKtJ07v/KGuiDxSur9jjF1J2iyaHFutkrvCuIcG5MmyE2vO2
vXsu+wojgOrmEOirs0d2dEKE53DDHWMQqJlb7B3DAhT34mixxhTUWpVDb0/6yrGZ
m5hug9vI2/F/rYfo+SMMDP9QpF42brEn/zvoZTPeouw/dpgnJKiMN3rk4iEwA8tc
WDu1SK8JRY/ci44Ef4HjRLbws+j7ZpygxmJH6l/NZ6+/Lhk6e+lWd8MWkQXe7rGu
9jlaLdFl2gYOneuhG9FdLKWSzldWFTNRvyt5W2wHRcUtToLwtKaGmBbPzfY926IG
VDgG1/JjkpSNowo6LtWOqLRSQcOu+tFAoUTNwrgiwZt57gS1qx/XD+CMV5b6i5MM
rgGI68upJ8BMzcFXyTcR48gmB99/qayQ0+f39FLuM/NHZfPLMvUDB9qkXo8bUYHe
thDtr7aVf8QU6FiU9FhIQDepEGXWMw69dnH0irU272A5ryH5I4QChKpIVF95C1IV
YvUDVzbwMZRAKy/oAoQBBe8/lJUWIfJTqw4LdWvExaC45M28tINwcVZho9/V9kTg
lDK29XckSnfXqB/nnUHeor/2VWvFitGqws5HVkpy+B7z81mbQibGbQMythlvDO/1
EThdfrU2ks9Y8BljUKtMmWvc2NO+hjpdH7Ou8n70Z09Xk2QOu9PWSlPAahYEtruI
n/ZQtosptPQcl0ZdZeqTJb2c2M0nyoC/QrKLaTy0NVO2UjANvb7sqXWoaLgMgqTB
ckpjaarf4H0pWwkwnQCNHXb4BfIR2fwGoV6nzXV/iQceDjlKnyctmnZx17g1C5ne
9VyxZG5/S2UUQhGlpqeMyfYPjwIsvr1u5bt3D4imV8YEQarqjw5oSDmXxOMYCwaI
OoYLAgCWNkZNpzSDtjOVkSkLmSjqfTu+yQMC/ZLIk4b1A+YOijWZ1wPWlnc3WL7r
DnUunsb2axJBJCovcc/lJSyFCC/HEPQZ/jWn2e5qQoIC757ZOlej/ypjARpwZGpd
ElfvhjA7Zrr1VFe+PyASMgfXFgSBwBaDKgz2Cd3iG/J6Tk+fT5ajkIYj3eEMkPZI
MjEwO3lmhjKtk1IAfTN1EF1NbAV9TwMeFYp3izvGOyi56QLX0gvAfov4/AAePz9Y
BLv8uRu9AOBqbatm8fVAx0TbdcZNiK9Rje5NeBFkZBaX3WF7AGoasZyNVVQVxlXk
j1f0W0w+HIJaLf5RpNWmFR7A0esLof8ahjil5z12EDu6k3iRQQzSxY2Si6sd3KGD
FhJHB3ERHO3G0sE4ItWaJBbSGU5KpHgZ0suO1i3s9Wih8z0s6fSIAgcyyTpIl23H
hnY7E+EZgBG5DxQYw7bwgr+Be0L+CBPUogVkQnc0HmH6jNFLFFMHUUv6H0hkPgQ/
VSdIclrWgTNiNka48Vi4Q3tjgkxsilE3MPjZeWCoH414Ts6FOoSFCzkExjIXHeQE
cOkPvCaQE5EsGCL6Kp9bc5Yt/AMXxV0mQmjbphPyjTTJOHUYNbW7eO2NX3DpFzGO
E5x1iJO2p+ufewyE3U4aHehFa8vgjcnXC7PuWpShH1nIq/ZGewZpZw4pn41GDJcN
XJaiwy/lej05mcI5SnkgBsC4Uu57ShiUCzjfX8B7Rqsx1QYPPgtBiFi+snB5R9+L
XxwNaGBTetjRHM5p7uu2Vy8EtLdZnV1P+TE65aJPXKYhl5SNVAEUfb00zdpsbxHF
f4X2WiG+IYutTTdRAF1WG+zP/t2Dcz+AHl1TfwvWwIqywIJ0fZH33adbSvuraR3v
0ZLGvv6yUM7nSxa3bZxbZ1WQsJTWcJy6XNByynzg4Y738jz0+ow8dP2raLI7HDek
7nu87uMwLxuJljRcI9zh835gOyCxo/kp54jcHiWSPMEzTTCukQcKGWJsHsr5jTPq
6rqXo5A1NG5gRS48z5VjgYtI6mguAbn0g817ZER26jJ+S7A1lBohrppC7/8E6OGD
Z1+nuRKuS1oGGh9AZ/Y9Rmqr2VVP/eYT5IBhUa2NO5LL7v7i5D7PYcaAu3P2p2RP
YMo6kdzbdv8BeoacJPixNxFrMQODUe1cL/xJtz8hZZRHXu+43VM/HX+/lX134KcX
9s5P54gqsXYkqlb2Xfr30N4sGvcl0eA/+NjIk8E1E1YeOSVGciYHA0X6HU9qCy7C
MhJO43iofoFamF4Bd5zT1gxK+DGQ1nAAQ69bSpCklQB0/RY1ezAES4/yk1EgODgV
MI4ZyI/S3N5XNGWr5tT9gUl8zBxIcvMvhFJkLBCNKjBxvJD8T+FmaADTm4kx4Lja
FXlHubayILdXLeqL5VLjYD0H+1g0sAl/Uq9BqTB1zF5CUXnxVmKkRwOkK9G+r/bZ
sPDOUfJPEYM7cMIYBtfClejwsz8PwoANHYsKmZ2bALmbfpe+HrVigE5gtjZZf0G9
RlwR05RLoweTEAapb2KreKdLF+X6+Nal2bFTbMuAm8Mlq6Einfa6cdoSNxBfns+P
j28OxMNqp8HpfhmGI92Sc7jhrdkQsDXAtewaR2Urln82vUcjAsbwtEJRC5KUJg3o
rmu0e4QJchpXuPYqH6eqpMCokDI7M1qyoTDpClKvzrDTnYOSbBUIUTMJiQM+Vp4u
fYY+/yP+E6r6yn+++oX9T48ACgNHXyoBQw+cot67GDH8mXCQ3Tl1n4soETDsLjgW
XkYyXmtjDc6Iq5XuU/dCNUBOiRtWPIJeCHrl20anINBOiiUSCLQBH4ZKjjAfmHtY
twgT06F/2c8i5E+0PQHt07h1uZY+N7IKXmL82GjDTVNC+4qk3LuRm3IuKYJ6aD/k
k9IccKd4SD9V1T+c6T4LA1ixPoi3Sb96AcNBKwck+fEuMOGiJyIkrLwgbNoawdQI
EAV5Es9l1SeDw6GGFjtQhuzoL9b/BgkuySEhaLTQHs+SMhBMzTm+RqvlsoSZrHTb
+JUZW0iyUfB5BnprqYAP/nNxTkOY9+zbiD4q4y8Fz7Yhu9SmucjXrExX2R5W8D4b
dtZ2smc3CWk8M6FdNZwKtGGmwa6ywnHaMjqX8JyoUVZX3+lMgijUdSUtHvzCKxio
Lw0bA2wMrGw0nGjcGGEy+MGsCzgO8fEkeQGp7KHxtuRNPjIxPY620q1Alz6aTBrt
FrCRZhVGyD7ihI74LE24r5HXnWcuxSOJTsiOQk0GbO8dv/2cKHuF7adhyW/bNOmB
Fr93Yd1+rhQ4uB+Rt6mBkyD0Z8dTgIJ4MFoilfcgbybI84EvAiopyQqsRPhhpLp6
imE3HGzXIyGGRjObyaQAUDUCp+D+jyhqkVtaLxfKh2Tt/WAKliKt85WX23FdyNf6
SZJAmdVe341j3uVXG3Lo4/9BRw9e4AP0KqkEJHd5Pg5EX6dgdvHQ7iUlQuP5kEhk
dACyupHOgBpaIuYu5+/KyBGpL9bWXOH1TSqNnH06SQ8/PWU3Lj8b/XM7m4uHxUei
/3xx7udby4WXawSREBktDCVZM0HORefFsE3DzWhHXGNTA2liUgB8KJ3IJLiowdo3
XM5+iupjmimY3AVQSEMDnaGu6XnxVXVspslLH6tOuJOMq4Ce+18ZPCjOGGLxmZlR
VJMPq+YQMF5F3wC0c29R7cBI5KORz9TvGah5IUEZzE6Zg4XWYq86ljpLtbObLnKF
YMKu10eAkCulRgrDN9big8apIWFlF+2+Dm7GMNyQtueOBKya+4DJRWaZA5afh+wJ
iWUaSNzZAn6CjetpMwpaPW/f9N3zkvKhGE4R39Tkm/BKaUZ5yjPPZ1XxNSPTHc3B
4Fx98Z8DPHdTNpLFDfzKAsG7jfKvVy7kzUBJxUCjsfukL2So+a/5fsdkO1A+eTMe
6fFcyEdKhIobIByfrGZC48wI9XBex2K9wpbGSK4sYxzEPtKQXkpouv8YJHAezDVh
JjMsovPaddOP+S98r4pcA/hLPGdpopgik3d8FJJOMJwEEku9SVsR9EtjJ5gAL6GE
M01tEANcNYtukg6txzoaH+awlI6f0eaUUsd9hnyEBCqRYl1stGUm2ygz1JU0e2ft
qcCcP1/6oV4aM1tJVmLFGqqyIX9KViq1fpFo+IhbdcOP8WVFEJqLAQqRbxcohxhm
geZYssGzGjIZZOTGmbW/0GlOYPHeiUt7A5wjvBcjw5D0sb7kq+B1Q9bnLGOSmdby
x28S0JEo0WpBXhMewkZBF2zYvbYy5zkiTFINtjeW/kpz6gldLPBdA2jw6E5OIqyT
wFfkHTy5LRwJc/ToXTLVbyw2T4+Y8zFJ7i3gMEJb9TAvxYQCgESLe9MC1qnETJSN
zCYV08CbOkoxCezJ8rc9riN4kXQVfE7TOseHrrc8ZDVO1fSK5urCVWhDbFFaFE/v
Mfr+9CMPJhbvfRi36WcQSLP3zTja0vJpOktsbt+fRKm9VIeIivyNesrPFGex6PVP
Ldyv5coEy9C0rmvO7FEr7Q+Hr7xoqHRIajUeq+I9UH+SyDm5n1QRc2J/SyhCcIZH
vgOsl83IbXzyJVkxVJu+tkCRKWitE/BFBix595QC97yvgcpaz5ey9PRJhTy/tsP+
TmdPAqwLTlHcyYprT9f7cnEkE0zdKjduVAFbiyPmvj/Ohv6TVOK4udROmLX8Cdmi
/LAwIzDyj0ovEq6l+PChR8J4m/s3MJPIyKPudaLN6rDGcWCSVemYLiPFU6SXbWdH
Co/oCRi7zZqmgBLhmZvMZ8yUxwhjw/5CAUZbMgWzn3d5h48xH7IVTcur+Zq8XTxU
3GFp4e4QgmJAtRB+yudj7UFCJ/d4dVW24R5rij58QB+omj7Doi6qs7bLsCJ8Ubn/
Musdg0+xJn1Y6/FTL6gOqqw6D20nOTfcgm6kJAgawfRmE+3adYnobscop668Ontm
FDH0PURojLdhHJi4f/HEGz9Gkxpve+MbYmk22yY+AJtmB6ehpTuPucAW7I9P6hI6
SZwX6WL0uANFpa+Y9dLgkhFfniAlDv6F//Tu7dabd++uDB605tyJVmharVeWtvA0
s/8zvJwghhd6nIE9ordo17wPNSFgnxgqsNwig9agyS/gb1dg41ODFemEXtN6W+c3
VyiQWmHBeeix1ZJT0721aozp7WqbPBynw/+IiLqfpsm9u0L0ZuLTuzIRvkNb0i1D
MZI3aNGakrTmUMMZbxmtwBY3Q9bFNqNUhizKONmd0H/Lqaf9J1LULOqo4gYfTJ3O
/mRNWBfJPzP1PQLv/yfRNs1ficlQLr+awDg0TV8AiJdd2Mx743gzMsTSAfBSn54C
G/Sw+WqsSiKXmzLXMSEeegkdlx8BXQKozwCAhBG5ycTErcvU4Bh8SjW6AbZGGeQe
o4awpA0o//+sOfIvYDvhmBE2+3yR4bXbP9vvDmMqNuV5mjBclvP6gx+0qW4xZJof
0pvMC9pIYTaVcPxTzUR4LhO724nHxe0ldsHw1Pcki3A80icHszETMF/678ez7OUk
iTb7Pvvn6Uv+fsoCwEzV2y86a0lX9vMrq2uUTjr63m3ZJ4BIwNy16oivlpVmoBpu
PiVBjQalKWv6VekI+ibM+ViXJLd/Jz2xwzsOU0ShFKn7s0RLDzxZQiFk7Yi5ZEPP
cc+P3wj5cef1M5DvMwArvBDmTbqW3xPYHBUhOHzLVTAUhAjVCuTEB7bhq5GUH7A5
QhINYh4bgHpsRHppwz3SZnI67KdVUtg8TW599ICmjnuSfyvTXGrMi4hrBxV/Y4bf
ElpFl55y1xBbToi7k/V3ySZJMmFzHtt+DXcxG3f5H1eZzjyDdo0SKpvidABGIql4
ks7Rzw8UNaj8sDXD3kstRB6TFk92A189btDSHWNHxx9dntAkyAahkykDpdLWINkp
YUqRCoCcAQsMXmlzPQEQHWyqQC1xyO/HxvrQr/Oouv9iwqk8NcC43NLtSuei3pJG
a++qxSMBeJz/nb/1sQhchx8Es5AKqlOlX0aOZvI6b3e4HiXZbuz8l6IyPwToyrQR
BtpiY1yFW7EtK83VdcR9VveKX3rdWlwTbX4H52yBbSzUvCB0xf4S9tyP6eiQkPj4
ydb9GkSmtOhcilp5RTfMq9y98G1Ww3p0NdjQdCbkAtidetvaQ40P90rWK2xONyUc
nZplzCvUxZoD1DV5v9GhzRxUV//SALM8kBjZglKR+ntKJ31yuHHiWSpE8V2zshT1
/FDXLYRJUBQN2TDIiYRuAo/ELFqp+gDT7XsRKDdISi7F9wWoKUQEAM7rcrFmdVzn
Frg2xgr0K9KafJlkDXR3etJfbQaj+yp/7iKNbuCFUT82pdbzqdXTP/pvaCYPbdYH
GWZBNfwbmB7dIn4FSbX6dPImO2E4wHczhRm6uHOATeAq0hlWVsj0ZQ8NWWV63dsy
4eecgMs8hChaKXHAtPLQ2FBe28Z9u0vHMboIRFMjN5zj4n0QxfxAzrdFy+kZpBJy
gOVHam49kH039ybkks0xCdhn+kGOpXeJuXMn/uU47JPckQhTo53kTBS34aIfTzbt
Z/cJMmzVNgB20oblsWpHZyhtJRASIS60GHWumSspvzeauDj2j4ZNjwxwkUyjVt0F
pGin/AXzQoQaA/yL5HAqyInhuNtEcVKdyN6qtL83tCa+Yz446Sh8gsFKBcdo8avx
5gL6lI+HK7GoVKLozsU/JzjmQbJNPriCyVIjtmNxhBcIxmJOYe3PHgJqB/Fape2s
lzpt/wDV9CzH8AhaFf5xJCK0vT8pp1yz104ZZ3DvBxdWMYmVvnBXaydu7kA+Db3l
1/ui+fT5DwSAW/OXagQSaBdBYCiWo1lbfW7khiCi+R5Zplt45Pqn+LBUAH0ECqsb
Vp2BOECGnwGxGl9SWK8bWTS+OJRmwzvlX2BqlO52R1iLW5ZWDxnRZD+GhbNo3fXV
B6KcNqS5/xRRCSI88OPcFJ1VCo1vPKQ0zK6fJIxJye50YxQXjQ0S6H7IEKsOau3m
fJgIpj+4qIcUEmJqyw+FpxgWrHP1cEtG1p22JgCq/FvTmP2quNpQoIkcjc5GvVZc
ShhpGhtDVlyAl0+zG4DO+JXArY2cRycZP8XlOhoe6noaWnJelmuTjM+Vcg37LxqV
qAcyrLhBcuC4/wUV+b9kBtn6n31yf72PGB6WZDytx9M650eAopJwm4YNKP+1IVfK
8K8bYATzg1IC03jF2Ff06YIdmttXOCGZN9jUEYT2DGSmJwIZ3Bk3XvcwmOvdMoRo
I+dRS0r2TmFfuv7vlaP1xRSWOgIuqH6LNU143bSVNdaushd2IzxUKgaljN2xZAc2
gn2waBKJrhh8MHsgFxoJsfIE0twwpsPGsDmPAGRiWvM6Iy/61qAuYyPwGjhxLVbz
WpsKE+owRqgOy1ApA04KXA0LZ/Llg+dq0ibYm6D+5Y2gjK4MRcBysog+83C5aadu
TWdj8MmVJmdk1YwnDnD7+H4DR4J3H/vCvq2rzbj4PsGd07+DfIZJzoxXjjGLJrt3
HGDSInmxd6Yt8rp5ojbTmBImJKg944Rc6PyNh6rLTgw0/igjAep+G1d88IpmPjqD
yg4fseWiNFNAMjd3ah1KVkzrdiFcgZiXPBCwotKr5JOPLkFKc0mKcc/AJGT/ZbWR
chC2A95IPa/equEjPj94RFi4LGJ+whPaMJdvJpYBeohxD+MonwvYVwq6Z3F643nH
p+cMQTARdWZkdSUNbaLadg1rqhXF4JDn3FwYJRAk84soCkqbDSIgDiGVc+cFu+At
vEYhErI9IRV5CAPXt/481S941OaypfuTH++LyxdPqAHTMWM7mhn8S2BtZ1AeHGUh
SRSipmhlZWLxH55ULBKGD7PQxEIUOp+bKBeaD5WCCTmmju50jXGA00ski8G/o7z5
MFHSHfgDhCCnjGSaAJrxYFK40EXfgywH24uKpSyM28zwtwxkSC50bmwCs9JGxWzW
IDd7QBJPL5U28CvL4UKzVNriAnommI92ApA8niirrxd/Kaar7NPSzvNdZwEb0S17
pEI2GCWLsZxUazHTrPe1YvE+Qt5GQHo+mGBw7LIbN61O7k50pa0vQIjmPwyJYT1J
Ge4vC8GmuzacMAJRm6mZVbUdzNdUJ3jEhzmhUt/oe5ALsdC+r7OdiRd92aglCfdr
diNK35tE5bJ2kz6vi/ypWdMAY8eE6lkN6D9T+LONOTVVCDtwrTYtR1K4tLtIVBTQ
nTcEeOx+iaGq9wmmjoheUhzsH3PbMbQ6JTmkeY1wvAg1Stby2npkA97SCbWNrwBs
cw577qI5adqAtEvkT8RrEAm4jhDAXCM4qt81Jf0vmnZgdBGOPHNiezKdiedMQJZR
tXNIA0dS+2zalo5alfZP+XX7VbQblYq14621nbxbs8UsfPUzMBb0rnlIGK7wLktV
ZyuEcrFcQYLW/qAjr+CxjnjokpIcrVKnmYY4kaAsSacIboS3OjaOAtfmj6WtClqU
/sL3dT3BhBBMdrqGHiG0FL3RJfe51R4JxT4eONwxwWuoV3IyZ2ZMEti70oc/GTR6
Dmnua+Fy21bU5NgSAcE0G0yB8tBTrakhTJ0Oory9bLWGjTvOFZOVKOSfaGAACM91
4BncRCHkpAfqYVfOIuZzBvWU38D3zcQw/T1fjt6q3z5fFEREb3zvJWJ09444xx9Z
EM1XTSPJm5i3cbeL2uYi4SCD8TvKVwQ2/LGBoTF0jp60Cl6Aj4Rj8UquvpUzfDlQ
40WADoBkqajZeoE4xP+zLwMaDTFZG7H1q+kM8MNfynumkxUsGvF02/muJyERcTQg
+KRaozuIZjKBuo1KFamlAZZMw2Cneus7edne4SDdWDwLF7LJgR3f6UgG3Cru6nA0
WNdAZSyXcPHTRcq89yemv6M9ZDhdOGD6g+6qo8u3IEfIA3hpjXVQapM97xRgD7V/
r1mxUhwRDa0IrLGxyKIM47PQ0Uf8LO4a2Njhm0uQo0EwXmGNbxG/cQxHn97HswLk
juFlZvM+X0a4xzdFQIQJvfyOjEVyzIMCEjuGeq4qM424L+wZTZxJGXSXCq6siz5C
hIpN2PWo6DMflCkzfxrcSxZ3QjfUPW+w619Se5Gvm51F1shon00SJfz25hGC+3Jf
/dUQ9pm1mlFzThgjMsJ26SHGsRJoz5OHav5CsbAwfw7SpjMttn/irvhVv9RxtcBR
GrI6x1YA2oaOH3Tp6THBy4xgrP2hB4GDByOmsPAydMKhVmrEZYk8F/5E/akmuLiH
IPu/w8Ogv9VkG1lGN9jZND773f81V9IgFeDRiJ8aW8CDMeGnEQBChZm22j/wURF7
SNB9JmG1wXl0C+VRROfxOAcQ7XsJ82khkiahYm8ZZEzNHHpa+6w1QIIPDRMLWnP1
LYMtTKFf16Tq8M95pR6z+hQAYHcpShhmE3gCIJh2WmSwenOKnpqgrIY+QMdoMmtQ
6HsrFbZCoVYCoLO1AHHHUramXFBqZzpeyUkya7Q0hbLqS2EcjBpBwirMVudqKSuO
Tl9Pc6+l66Mk6biGclAlhKqckTT9dWzAu8VGWdZaoMmVVLZUdo0quLbMAdjm3Ozl
yY3Ct5WzAmnhQc6wZfwi+4WHO9azlUiFbKGvDNUaF9pGBOpx4Lgl/mbCB06ZOvg9
D1qHaccgMERyVC2Y9JosBVutF9QwloWRff+fta2BfGbzBcff/8wxtMemI2orAmqc
jeg09z4c6uQrWi9ID8KxyO8xlTV5ACwqe6zX3W8gtoD40nITAXriwGz2T1olKE1m
XK0hptOYEAI1XyQLqYca9bNd7EJMSS87sJJjY8jD5jlWuMtXL9l+scBVG6/cuFq1
cs9l+51Z7o0dAnpN5rj4HoniWYmRyCpyOb39+mbekJ++auYWOVKYJrvfVc1TNkGV
E9T9YxnHYRZp+Qz0dvq8kyWvtFfOfPlGSE0NoiqnR4OhKB1F3yTF9eIEAjFVOEUq
EStLPeoPZR9t2VAZWj44Dgqg7Eng8EhM7+GnsF9P2hCb6SkAcyGBGDp7lCcyjl2M
98698GHVx1yz2ac6JW+vj4kA6kU+CT+GeT5VMRDmT4fP8qPp5TWw1i4MBwFRRl52
YqJsniPCqZf2AO/gry5mcHKr18uvmHGWo9VB/BqS4e6EPscqEq4D0yIq6LuK4Y+r
aoB7ZMU4YI/22r1iyup42Q6JLUE9mdUKFS5nfLs07PzY4806BtDAheb6JxQXadYn
KDHuWiJYfKSzT9Sy8Dt7ZC4p6fJ3KhMntmtsBywIK5oh8IBd86vg6Q5CXkxN14wM
P89hoZB7VRsP3o9ba2bQomQoimLGFEec+MV22sMtM35AdJZ7uvhVEleZ+C5VUXwp
PLSS59Wd81JsJNZ1n0x77tHJ4tPG0lfi6COnBJAK7VO1GPZBEDWEKy0OfOfTzCOM
Yr5M4cqCFtb7gwt6cTdtjW3Y2UGAPwg09hdUdaCdX76M8ScRTMBusd3wBvuR4sU/
qwkr4r1oQWdHMP5XiDq2CWwVW3mcjJuTnB9CzvLJniZSPQnBnaBBasixVC9WNeUW
ImbDrb7DTj2MqmQeuihG7HdoLA+Cr5a9JJ45ujK3kFkBFWYKUQDuyCmRx11mNvUt
YJe9XgJ8MS8+n1SAxQgYOvcHoL5c7BlxJjA1ZI69qjut/PetwDW6jVtVS8Dias6Z
XDbmeSrkAJW1VWHZv5zrwqxSq5g8FJsk6E/BbJNpakTijiTodaYIAWZQQBv4MxrX
IYJHMAHMkuGiC/iLWaRxKwBFCS0RGrVjadNNqygqWd282KubGnXhwWHai9XrJhFu
iovbzW6JeO+jLMfXnBANPRZ9nAQTyTVT3n8PtnyDql/2IxDBcqj0zYT+IyhoXHe4
cA3waHVYzhxDg0l6v5BQOLJS8VmD6U8SbkoTT3FzS/jVDRkAE5Pk2P+0aHSc8aOu
Y0qaMqiIPMdDPepkpQM20pZjIvSaZXXaQLo4bs5Ca9NvTBkfAAMhWzRISbEFLaV4
jZ7AsuIf5QVawrAmUd0Jpq3nBPFsFBqe59tqPktxOf/YzrbLh0gDn6Dpk1iQGKig
a93llMoulngevlbTktZqgqrJg2BBzLUJyAgR0nsSv9AfJ/N69AprM0KwljwAsgQQ
rU7AKFZ4fFoToJf86bE7qhk9zbV+wBSSXUe8k4M1tY0R5GbrfMorTpvO9s5HHLfe
IDP9u1mwQzR/ZRgoIs5i+6x4GT7OSdxQAWpdpdn192sV4Y3SuLF3WcHt7Y9WLz3K
ZSa8741zpKpVuBuxxd6w9qGjnBLkRsdBn2IKqtEawUEfzMJe6sJWS5aVKr+J3AXa
LqCZM6GO0z0jeGogIClpReI5WciKdq7f78kK7J42I1JrxG2vb6Pdc6KYDQdPuUHV
OiFulAjs+dH242D/OUP00BXPs3BJxZOSZDcH7uVdZLWj03586sWwnJhWw8k6FLTQ
C5zHu66O10pj2R6oJdl8CQ8n/PD/s0AUj0uDTDKHRIVXL6pp6SHRr/wPniRhtez7
GlaDJwEkSdW4B4b67lGFtSo/1r32vgNTywfR+aJbYepPm27WJawjaV+2hKESKbGL
3EuQkE0bn3oMux/4djbTl25k9NJjBbDvKfIrC+HtNb6z63f3zQvty7cmaP9NrwiZ
v3BYPXgDZIxy+e4ewdGvsloWmL03dk/cWA5dEE183MSlrepVhCmyyaBBMRq9lMcH
zdyi3vRTUyfMNHv4t3Hxzi12r7U9M0sR68/lqfDVPQfJCJx7RkuH89nbgMGYwHBS
UPcwrBoUsTNf/7MWfA1l9t+nt/SE1GuPuY81tO7439ma6k/KGJea1leqN47sHB/6
cFNw37nMc4cNvU2sgOYJAdVVOhIJmzS/YAjquNlC9WhBSRDLf7MQFNL7SVQvO9TY
i6fCE2WnemfdseS75gYHt9Gn9LZOSybNcCPcM/AJpzQM983eDiYjVUTMcUJDDE1S
HKzzBlTwkccPKT3maRdIxmbMeRyMMNV+MvXjXjc0oGm5/Zh5mdOsRsrxdzN4CMBD
BMEAM0auJjT8cr5dwXbLyj6pun2gW8NizB1gAioRATd8F+NM7Af4lnoXh/AJIpvj
ruD0xlWOiow/Dy22WStGfamh4ci/74rcWNdRFDsCSlx19Q8F3K58eSXqwok77r2D
PE/c0QkO5X4Sd+78840zkPZvQIF+vuDoEjV1lwYp3rdNEMSd4PEGm9m1fkEvKlED
N/KnOScfTeFc++8XbJprTzYIKFCwBk2ffR3KUjbOO6hA6kwVzUtmehd2A7Hr+ZMy
5JJjIQiTwoaW8h4xzWvv1s0nZnVWLOYfi5Vy7sPdlqkdpMldfBAJXmbrzQ8RKyAO
KYe8f5/Arvplt0yVKQaNbCjQ1NbZQ+ug2nCtqKTGgji5PgWli9GGqaRGigE0g69q
zXwl2dDlNJBMB2J+i4P1G36hUQ4wB7k1qbAA4QawLjRO8JnoIzsFAHdaAixiK/Lr
bOyG6bWMxDEtQfN2W5dLbdLxzFhWD+HVeqvGhAtpggttMdgv55fd1iGZj5vv6cps
GcKQ2T705gx+Rz1nWKAK/C1wZLTuEdzrr9WoK1Kto9GIX9ilHCUC7t7ZDfJIiB4U
Gcjj1G3kK59WYe9XohRxsk9O4xRfk8ZxlSq5M7vZzrMavMHgiYhLTnZfj6H9HQ+Y
ETC2Oa0O32ha7ztC0YQCskNtQjPYjD1x3+20qXdj5BG1E9AHtt4WSbZ63ICiqwPF
L/N+XKkovcYpntLwF6/YXjO+bNeLkUdSCNepcE5VudR4dcliKDzRDo4+uIoLybm3
lp2Jfo0wgnpRSefcV/eCD7lfQusQoz1ir+A8tNbQieLT63lXn73/0vTPYBhuD8Kv
i8KdLABrcJhUchxpf+jnqvplSS3bzCSxXbd6uxCenCq+60QbBchHgn7fA32hyWsc
DNKNMVpkfzPkUJpYXU0V6QMIqpNgQAcoVRRmI+Gq7CymWGds+xCDG4f9A9O0inoq
06MkDF9CgO0Tx5usxG4mM+TUMZwrvLwx4ZeaAUsCSUfOoPldp8emlAKpXcdhg49Q
WPdWSZm9nM3Sg6dX8VSS2LEw8OObGM7egWpL6kT3KmjTSYu8nXWUZfN9lte9nbIV
96iThGIYvyoOL/BhjXnIGUnXX9BqF9u7EXK3zf8ez/Hn8dubDlADLait86kwTS6u
I9qMO0JPs4Wwzz1uvhiimJ3GrYpo9QgAr69wlf/U6zpQeFOzU38TVwgRPFDJP8ds
MUP9i/VCWWHxsQ3W581Avp+WUxZvF19F9tboPqbb08zhrQpR/7borK4/njzi8M40
8bmLAWAgjSQ+HOuQa7OqeS5hQtav7JNmdpa+eHtPSquEizifmQ3W82xHxgBKrCXB
HYr5nXnLN/pyTjgcGglnsxewoFE8P2KCE256Qs83xT2lsEsaMG+gERf1nMa1fuDC
qLoBwrh7M6HtvRHfbKse9RA8gRR6jYh0Ue8cHqw1g59HGZ+UCzttYwwkpr6hrqbN
f7ITlhbmUv30SfPJ4r5chN4SZ3sEehSVPeldah7CbyBsh8UmC3FOmrqydIp6pGD1
NRCKvCmXU/1iIC4oT49J2XkAZmyPAZnLnHZ9+ZlNwCUuuZjfkgm84JHdui+E+Mfa
uo6ZuL0xgVybaWJgz6ammwYqHnkWdRjDkzOYMFvZKCCDlExiCB5VIhLBb1mcyGfK
BET/fLkBGmSpqvJbvxs/Sq5Lofd8J8CCAJX0KuXgpC/O8dUVJVAwOMZKV8enDeOD
5pedQrjeDLDFDlupaQCSG8/gLZrZYn+nj0RgyLK/lxdQIDXUsc9DB7PTiRQ8f+sV
2k/kn1QVm0zhKLlnE1TtPHuIJbwY3uTrtlDcZME21z+Eo/tLeY/z2rta4n0JOWkW
RKbfxf8fQxDpZxzQIpfxYo8fZBaEI/kB2G3pWP2PeoFoJ9skhmMnMP1AaQM1LEvM
xf9DGAn5w9ehffbBMjL4QcIMi1oQz0wtjP7aTVKLlX6J1bBTiIE/vpdexgMoGql/
DbsiYiK5HifVHuvZuYkTuzy6ShzusPK5o5wwyJwANI6ANuSphibPFLluz3YVQIVN
inFD5jC8ANDIhyxbn7Oy9F1EDGDbfuAvOpmcZEUeYNSoBiKlE4L3MNeXEa6ygDXu
FJnuZZAQRPO+mFlW/tny7YOQV3Ggv+lLexAkYMC6VTsxvWoxW+4wCdaEKdsR2Kgo
Ukr0ZfrPucRGJvzhj681ZxP9XAHHAwYBMgFU1dq4rcY01Zlpk25+R6KMIOH6+yZw
gbq/uoQkL18Y93y68I7W3b6gWEPH3boTvR/o3D1bRQ5X5uNYvUykSUWORrH3WoKX
XF+U6ecFcgoQ3/8JDrcQVkOwJ9uUlLTb+ePvg2r/ZRBh7d+nlDlhpKwJoqqyy5J+
W8fxogbWImn5wG05NYrlUt2IwEMkc0b0J+gdvCrj9Ez2hdT/DPPyTnsYYk0Pc7DD
N9bqzdf4pFbs0TA68vm6Agg+9H5TrjgR3Xoloyi4pujCNe/C7l4IYRTvE+F1jWJt
7nY9WzJ6allwPrmX/hLWZbUUXrJ9WCpX4r1d2ljB3BpN9C8weGGRIA8fdVY0eNjy
7fyqjEKIU75wIPleY23eAR6TAlaSI+eNwEAP6XwbP12QC6siQwkfFXVVjsAzYqr0
JNOaShi/WL/gNSv32cwzl8MXKNLaExP5OwVjn9fB2wR5JyCgEHawS//Y9bqTT9Vm
aaoGNTQ7hP8GTwGCejX8sPReJrRtJSQurMWV3jcWpPnEOrtbxN5gjAjcL9cHQppM
d0LG3NyAfJChCXwR3c1QeGyVpZmatIktg/diJUd/6eR3CJpRBv/F94yEctgR2dU7
0p8H+7Op7LfJD4HcKB9WvjdvgEsut9eU47ap1b0cFPhSYtAOkXt6JUdb9JVEzBA3
na9QP/Thtlq3kFIKA3G/YMIlFrwy8SBLRSat7zztT58HrZYkWSPDEC28swqto+Ol
bTtgg2/E/5r1CBYvy2/O7lQv63mb9+PozO2T1jWNi4kiycs8zDXzVZtYRc633joD
lONV/y7oQmTiGeLhySX/3EDx7Xs5lp3x6+u2pHk/rCCbnOb3gNhOUTIUUbbgDuu4
O5iaQH8qsmiIbjOyAY0ce0MBrzyafpQtFRpsdotpty5vGzVEqptjx+XPxAwY3q8N
8Sy0rO78adHgZS3miuNFxkj8CocPOreZkgIpK2wpzRu4AzfbjsrIUHptKVo7hEuJ
fJ1VoNyIflgM4GljCrVW8aTEwBmo863CObXeTavu4UfCKyPGyaXegZBP78ek57nO
hfG77DtwQzFKeOGIH+SwWs2UjOFWIXEnvElyWoOk4k0T0ZrMUD6YKdNOr2YULTYL
nnX1Qw0hRR3hqGcd7faV+XE8wx6PCvjWhELccfDXmqM7GG7AzQbH74fLjSDq6RxM
uFP9jQMbG56VzQ6igrVSOignHJPtTXlICch4J0f6gBpQttYDRhrR+n/vxexj27U/
k7YcBeF345y0cmedH4rLwEp8ndqUYDsPz3SsBONigiSwp4pFtilhAM0iGRBLANGW
y6j7sx6z5wG/t7X/VRxgdcjBGdnb0iaU0vtXgE5NGI8ffrWtPFvV68o1o7s1mGp/
DjlBj8P49FSwsyTw3+PuWJhBbuaug5KJptvf0hL7gehFI3ZiV/ve5e6a+vadt/ps
UTXr5scchC7gbB9mnesYwAnS0kN21sNoX3FefvV/9lRNjfytTcd3H0cO3TwTAtIw
2LWu+zy1GkY6/JPYa8KaZLmTj479oP0LwdGC1iAdWA/KubnqLkgWMThnk50s+YvW
1wfgqN/LPJrIo14TL4CWJm+bVFfo+LigRBkzMHfodS7fKsyKSjO//FyV12IETjbs
ybNOfrET7+nMfh0jvWnCpaE8hhvaxwdFqSpCwtnkbH+GSyGL9bIW0TQLfsp/v9CJ
+Q66Zu8Bzknn5vqDuRHWsO60Kf937c9JTgdjlN24jUSpRZCiG3lAqOKHm9ei+hkh
ab4RJq9rhVDS9TKtEDCEykYpfbipLp4ZHpRuhkux2YhGCCQkS0ddabggKU5Ytw3V
QR5bEn4OdPkabmsY7LJGc1z+IiewXo2bkxPOoL4CDRcOgOtXP6/a/WEYdgC4lzN5
42pZRKoMfE6+Q235G3I21kP8P4nAN/hioNXvhQSpYgSOO+aCckFtPsr5DAA8wJgd
7hSXYywFSDZU2lstv9hfgLIA0TaGILKJ7okJM2zOhNzxh3LUisEKFKCgyr6RwEP2
5a2R2lukUmNkIqSxo5r+/8jqWbWCA8ILZJKItC0l4I8kJTs6/PjlwZDF9Q6O2vXt
c0++dSicQVdobrb3R3Tb93bGVEglKgkxPojYl5eJmNQjCwAGW3KnDEL84HwE3gMp
Zz8bCTR2td2sA8V16RMhuAU2uuQiNn5P1MjScqwKJbJbANrrKt3+YW89DPYY4INB
kyg1ZJ7R1CwidFAJbqM2o3guaD8YwB84wydl6Wpuq0lFDgs0h/Upfj0Z2wUwAwt5
5Y3n2YgGwW2d2UTngEONQHu3HFQAG86k5C1615jckunZlqTeyMqQk7OhGRB6H75K
qp+GPBSTEBIe4gPW2EKX2eLQdynDbMIYgaKSFj2jHOwSAhY8DTEpmQb2473olfzE
4CLlbmhVOKhhuuZAUkzVdV/+XUXqJaxtJIoYwxql9dJORBb0HeGyaB3fF06Q1Nb9
bHCssW/nAA29ptDS5dam1isgXni1xdzA8r0loVLs5PjTAWqaTwa212YJtTlbuRvf
Qm0H9cEaHbkksVOsrMO7Lsgep9/auC3v8i5dp6DzuxncqxvhYuqtdejrK4J0BGAM
gCh9guO8cCk7TqiwDtkQaPtQ01HMlF705VnjS4bNQKe2oW1tlwAwU2+g3CezD/kh
LawYZm1DU3rbGe3QmV9SXrozKB2B/PtuSnAizlCk5sWsxJHaYcWedQoYj+ijqUt+
+0iPyIQn+WtrZOPozqgJ2EiFJPtWaGnvQp9kSC3Jo1bIoJgH11S5N30HSozv3drT
dLnCMPMhtLHPcUs3A1wuUeFQ3B4N+ySkv4pstnRbQbexa3HPJ/M7NXOmg3Yf9ivp
Gx3/TaYO9o++Pi/JQvk2IyP2CBiRs0Kt1i6L/Pkuez7ozsQMvfixdIh4VDJTwrw5
GTxDYnKLWW6zOBxSmuYAbsE6VrcGKF0jK96Z2NkFOHaqN94bSAfjOdfQHN9c7ool
h8od0swlJkHuPC12pUcd994qBuUqVgrkv7ijnGcqgkE3rN1xhn+6wjcjQyCMz6ql
06Ziyw/sDf9IIy4N4J7MhDuX4KYvtFOVQJnDA/JOITnaSqF855cZ9a8yPIfiWLHy
5HokWKL7Z+5hsYIoUJgTgTyWJNdclMoxEnc/H4CUxHkGaNtGy6DSciWj7MnoDzLN
xLrINAOJcpAnsFkcoRsmOp043K1rrTKDArajYeNNLFSYEX4cD8zfqZH8S1gaEski
AVltt9tRzs9ErY9tv1Vp8OPIQle9IEcJnwGBEG2Wm1Lb29mec3dhNI3eaJQWPE6S
GXDo1DUPe7UEkLUw/73FhDhf3crav6MsWXzazPrVg1Rkx3YnoDO04u84+v1FMyNu
uu/g1HdbD6npNIHdyqdx9awtOaoa0+OlY34CKqQivNjk63LP1FDGTmRx4OehSpiq
eMcYUJbvpZlHDkCH64yfbmN6xBvxF1psfzkmLjt+MFQjbXktVexNW89K13P4XQjH
KuX/7HCxdP6F4KVdnbPP8KYravJGL0nKiiQK6uLYUx+ROMQ/DRQNSO3m1rsAtMNN
t+rq2gkqFxhV4H4l91wT2u+qEO7OO+rkFhMiSX84QSQASUvzxNP2gwizJ+UwIHF6
EVUTG8L/Jz5kK+ymJ+KXWE1o+zHAA/cyI7W9h+yyDJ6IvkjGX2WWXlilR6e8d7mM
UY9Y4d1O2BqdLtIvVObHEP+/Ez7IZaWDjsayiSj8ubbjGhySzqwYpqCM9j3l3apQ
67iaTdtMVx9ZioDPnE0rOfmtNqtB4hHxF5GvI1glHwjF2hiQIWDAgmDddyB9GKkV
LybsvCii6Zry+xPBZrwU4UG9kI6yo6kpXCqi6U2zLeZgoVTGJWp+dnPaYmedkc1S
3k4/q1RubSLMMyDXQniKdH+hyP2SN2ED1AATvIx5EFXbdUnx4gEt+L0qECOetyxz
EgxsFGINbBGMXxmEOpL1gClQhXB6vntEvgvJFHld3Vqr1PULcFEFiOaCZvzbH7lY
cLWfefX8nrkNET9hH9AMjxNjTVd8qhOagWXDpgFoO8eX9CprzpTsuQwiRddoFsyD
NdF2KGDWpEwa3gUcievvtYrWSniYaYvOD2NFpCoWa31AWxPBPxeHkpsPgfmcPjNl
IUUjcABQcg8S4DXnm7gXfz2vkesdGEdYNwgl1PR6Z79xi/BzlIg8+IiYWco7vOSL
d2Ip9SFsvK3yw+Ebrb0+6TeomtkgZfHWYtAUyS4JvA2Els2XwaOObyzjb0Q6/UWL
AeV/noV+E43jMGYWqJeoDk9WMfeCO4zuX4IizqpfMQZcbT3DBj6dZyFVvgrDqrTm
Ohn7d+m9PwGpPot/izLg5gaYmMAgfUGUiYcOkJkuKymaznYdjhVSeKZB+yPHyoLq
oumvCAL9BQ553mF03IJAFAZMv6A1qmvQV9mhkfccOCgsayrcLnlWPNl5pGKT0MIU
YScoZMZ83phtH6rrKDOxknMIwvQRHeoictobKM/GmxFcGF2NzE3QyODMZGaQoIUi
U1G0BOPpuJFVdWDaEk7LO7RydPoV8Vm5e1Ap34b84QwnIxIbC5PoA/Ir0vmZcho7
rn9gVXwmEXlb6oplBjxtzlHRcVSSwmgNz3ycuEu8egzYbzEg8EyDXFT8+gxkaVIt
axFqboFZK/CJdkbqabhYh2aRhi2NN2cV9fr295SBqWvG2vSVxb4F5Y+Fy6r4438J
dNG5/rAfCn4tiEJxsbYVKSvTE25Fc6M49/TISHduLC7331kBbD5QN7uK6g2ejka2
dW0YatDbe1pvTTgchnI6L8WfS9eXDYjj1Xu3gX4ykpRqx65IES5B9XWuY05dLNIv
ZEMGvTt6FshcRsvZg1RDf22CZMLxYsZE6sKYNKyIX0h5PgUzf9LcqpDZ1NMLjE4O
4SBbMiGPeTIocDLBapSoOL4e3P9gYBeF/1mJacBh6TBf20L5DDRrC8AzMTqPp2Sr
AyzBpnXq4mzsifQAjXgG2G9rtQqScVRPX8sfHMhjBMimyOfGDBIxIXnCOqtl7K5H
Lo5dUq0BoEIFVCp7d81DJJ92B/ryg/feOPFqQCGO9tcS7WsuWOGi6YJ8fjYUpy7J
Xz96OPMsrf0eJGF+TeCkNRE4pYXIPzp325NZf+YPiNFIK0XUByQZe4hJKl3tdVzD
UllhYTZ9PBsPpHGUA1K7gFVu2807uX/Ph3uQo+sYGf2pQ7/cwfbj0ekDcDbqSr9U
B9HXUwuZwK3UQ2gInjcf4pNVD33+LStP/S3ELYBspBsnLN8ZQl+sVqOeVqgPaIBv
ncmzTTrSPZ5u5ilVOA5ogfP7ilx2pl1Tdz9fgmAlsXY8Fbf3Yv3csaGD3dcS32sN
rukTxJwo6to7sTvsQzrVyepS0lSScL6vxW672TVjIAEAWAqkBlCmTutLac7r8x5P
oEznVswfAX4Q3uZxT2/AX1Fh94eAZRRMQo7y+2brAVfOPaK3Oh7BuYoIygfsVb0B
0VUVZGv80uynyy1tqlR4HyOLLTUAO/N/yEkYgWucEEscfImkB6lU3s+1bidwbI2S
PmYGXk6UvxrsbMKTCKfdeNZKSCQ7d0xZX0tMSIWYjqdSO1Z/DxSPdsU8hdP2GDun
MMesIaDgLGi11Uqg6MOiofWLbkQw+VuG0o54+cvPfdwhll52fyItRAvjZRdmV56y
anTHLsN0R5RaGdBzT8DIfVO/s8sc7Pys/IyocTRuxeOvGpfe0v5MdWL1cITF5g+k
NiAkwU8x1o6l0gCDxVqfKMtiIjdhEKHeoOSoqtklEUVahGRJgnem3azgfd9yAGJh
ac0vI2cc0pK/GYs6FkCFMe00a0ICs57dr7icjvYyjY73YMHiigDsMgmN7Wm7m+Df
hGdX0Ru3yQgnnbDcroC90axN/AlFmiUtfaB8TLzt68Y2F9lUexlWK12MdcpqtrZJ
h1PRcJta2czjtDuYwL5ik/e9pxBdgFkVgoAXBN7yn+BQj5ax/CWzG5T0ho1XYMt0
GBRRTRkWK9Icn965o5PWl8WOwYAN2prA1OQOnxqNdswJtmImhQT9u0oRlUqi6dW2
gObC3sFRL3RA8r/9STtuWELqXFLB1ZKlXHuU11DBAYZGtuRMNcCIo6MkuhqEprjt
aovj5F0uPFiTVjFfwKthOMzdUZ36/EVHTMYzqusoGMh1+xCnhTgGgEeci2jCorlH
viLJxuhFvMlLwKnuqaRGRzBEfNDYofxMQxX4nPcCELndWsMz8+bnOiACdQd/c9nK
Rf8F/5xeMYvFOwz7thSRY2q1J1rI/KW//5pmqZXKHLL+u6dWZqhZKaefR3qzCOSD
vbFAYrCBm3wNN7Dryy/NcIB6ZPev/JvQSdlXic/ltQt26sKlm7y/dRLI+Pl4qjIH
hzGed3eIa74mYN8jPhhDIFs96vT5LrjtKFLbterPLF2IIgnnz8bD61QGjdWuYI2B
9JYBAzLaQbUh7CKJUvHFhGwZ/Rqk/JkShbwDq9vk4jY1K94mEQVr/jSWddGmSsBh
W5uRGCFXMKVnF16ubQ/QDD3nzYtaUfatu34kZFSDdppeanXupH4XCPvLYNB8X+ga
EK7ub+8AaWJx2VR12Xlzdtc+2v7mZdk5QIk6/saKX+9v6vmGYnPi+z6s8oCv1IZP
v3yIe1Do9yL/poDVDrbPPCqm4pHGA4GRFriIbL+lJpQaPuzBV4KAz75V2zraJo4k
o1Rtyh4EcCjJKgedp56mCrBPG1FvlgMBiXnktmsDe/gc4AsqOYAk5vk2rIUQQp2I
GH/BDoDkXQp970dwzpsgQJqKIx8bZD2qgVCFpHQ/fumum1eiIFep1nUpKWkZQjSz
XaQachDh8O/qIZ4eA4cnfrFd9RHCmqHId+GzrJ5/CbIWjCpZxkdfsvenulw8T9lw
NSciQfxpiAZ6DiYbyEK8JPseRF0voikBga/qa79MijhcIX0ypeSlgsmhX1UC9a+A
5ucsBV23KToT7CpsOKuDDXEZmItXmJHDK89lcSbhTtjobRYbvVKHgN49/UjI2irs
ysvqOBS6eYog2jGTjF0iCoGSegUnCs55oAuP/NtSNpoa1eRaRyH16aXW36Pv+VA6
87YMaJlElEis9GDpzGk6Ji6TSFlH98Yywly65CBhZNTYy5p2F2pPLABkl0JuIsuj
myRrd/uB6ospBJQVhkV8ffaz9YQkAwsTbiyYEFBO3uYaI52aemHDGQ5qDLlqZj6Y
oZHBbAWFL241Ag2qwhMUTPSWfDngSOIPiIUSOyIIq6xXAq7BOUcYGuX8yxI2C/o/
+kXU7QndcYHQtY+4xKDbkE/cmlBQBlo8CIeynbz7WrGFrzR2LksGTVJQJAluhvjs
oHKeC6zuGGHn1NXczAP2x+Vdwtl4XeW+nZzGbIKpsf090nqcCG/i4+BjuAQuRqGG
Otx+7YR0ygFFi/ceayk3M/hCuQvkyUDs8vsclwiDw/xbWcZsy0iUmT4Z9iLUTDL3
Sypp4C98rqLmrLqhcKcG5uGwnTwjatYUDXvFydMQEA6haqVEIsc4NvljaFLZhhsa
XOquvzWDhYg8+arAxHYQ6dcZJRdWigo00NDl6J1zRmAVvzAScbFkW+z8kGGjXVq3
lpAKYoFi7s9B5t2yVB7+aIT7Of/vL9z/YmSBOU0nVs8XWB5xK0aslvb2b2S+X1dB
KzzK8hHKDo/ec5YGq5SSw7TLAZ6VmqC0fiDuVZBUX86KhN4OtkywzzPhs2ZmsGoJ
efC0C/bsUIdPOAaE3eczTDiHodaGR2NIZz5H7s11Z2XhjUxjqhzMPM+NI0VvsAiG
aM8/+lBRZ5WRaVVvxQuN7pg4H6AN78QVhyx216N82Wa/44eZEzm+GrIX0UW1tiGF
nLRStDj4glwV36FG191GMz4jZU9xF2XQHOK/Z3Pm6T8L97F7VHNxycocaBDueuPJ
C4Id4+Lf1TbRs06mU9RzSoY5ayd1XucdOm4xGfxudl4e+dbMmGytOG2fAyhCEZ5i
tCin64jt4Gq8CLrsXfVNMwWXr0n0Q1JjIdLEUJAFNRGYFzn02hdjvrzcTszOf26t
JtApCRV3giRPgWJ5OKo13YcQQCvlt7DOL5qV4kKXt67dbPlKcQXqWQ9Hu5BlYpH0
MCk8i7IYn08/XE/GqkJezFd8O4XPKw/f3bPO8MNjNV+mTAtmWc+d3pI44HKyRyr8
uZ5WfwW4TcAS+Q9yg3gKerCtOhav9rZ/JwXSaRQuwEkGQs7WvVycX7dOt0U/yDWb
ngxxKxA1e4t3ZVllDN81Rzv/YduEjOw0zut9t73sKcrQbVhOxq/47uX+CErszJgp
+36w1119TVkyqYCUEmZnCuWeENODxf9DoImTaWSJkaMk4WpGdX2f+EeWHV90glfx
j20UvvHdiEcMaGbYvoVTKV54haKQ7Qq5wFfat/e1p5Ze/7WOGjAh4URgMG+E+Xno
D2H1j+qibwMAj7/x0kuwJm7Gje/AlbgQ3W1lXTMi8m42D9L188bzmTNwCUbKnC/W
/aGuoQ26Nc1mAXm0uW0jqdJ/DVlpF35UdSXR2xvwgPAEeMKlzY/hOmgqRnOwT52X
F7pjU8XAU6gxoApXd+/u7RcmuxD/8r9rFKMRYoL14T0hSivlCneqEcjlI2nKna/o
VUaNyBAhQVIjudONMDcYX3FX7skKwBq14PO2nRMrBLE0v8Op9YZKnswfkVotYhGT
NctCZYVzErC34jVBn8J1xVThoylHjEotpz7mEWSFzVeQ4eAioJ61cIQ5v7RgH90e
wh8LudwKaErq98nmUiwerbLVnMJNGx0APH8tv7t11ohQ5j72a8VxsG9AB33yL03I
HWXgt3JayFFdkcW31GHcDjxz3o1accW3k+DpgTaFraxE5NsohMySdTrdNaAISwgS
/tMr2Qx2Uiz2pagfjvpWSzLu8qQpoHBS1QjT6rgtx2ETT5as1iVdcNHGcczeW+OS
Y06T5lXvjfQIKB7FaEE6E30re2Rjni7Tvlq/LeUOo41km5XQoBG8ESLK0Uq3onWa
8JtT0REpSt696QGOOSHPKzd5zA+Hw5WQ8k3QzCTMAnEM/4x1FkJyLFIljJRUhc4q
qebgCu3F5rd2Zq19H+wQGvSiCV9ZGkrrgQvWXHBORZpgT9RDUMPaL2NYqpgXI+ra
u77/+LkYQ5xt/RvlbjFE1pB1GC6ZKrtaxyqHvv2+3KIeLFPe+lhgzq734qBXqECi
HbWt8mQktHtv51VyIIG1v05iGV9NhB4MWIg0LEyRRU88AUwZSY+GMr7FelKsMo50
W9Y7tNCp7YLJvZ41puX0uYg9b52MqsB9FvhLIDwMgG+0plzodzhtAVV/ObJPNnF8
pgfbSc26Z5BhtAyfMduWBPNAaUiMF+oDY9WE8dVzDxYfbiag0v7EiGyYJT1JLvvV
uu2qca0oltNs9+GbWrhQLL0irFv4lieWQo9d/mrCTCdm+w2gN6ya87DjIRHi4Ctd
4yWogNrgcWkAXvwdyIXoEdjh5N3AoQXWzvBk3OeOEo/keODqJtPtR+TRP+ilSKP8
JiPZh7Dbl4+aLgyxlxAnHYYaufGD6sgrklB98brDykPZWkNr3YIrD4hutxgoXEsl
p8t+VnSkMKiLQsWcvGTAK/g5ljkO64cFva99BZd/kxBPqPekZ1+9TXF26PKRtSpG
Ax/VCQp2w0JZsOVyOIoppnsByUW5WEqt9kgUDxWOEq7HAy3QmcU5oMgGpJGCjMT5
d/Py+RVQ05/wuFUBu/pwmlJZGGkL0RffE1vs03aBdEyyog9w4Z3MTlw+ox1wx3oW
w3xee50GZP98aIBimZTHDhiBlV0j1zkRKxKqHEe0G61so2JHcoW207hj2nNqag9F
pIMR0Wq43U3jH6nJ8Y6O1ZxJKo7pnHhPJJK9+VbKy9s9OydSg/hSBt+R03OInwVZ
ulcBQFL6g+yJlkjkbS5al534pMIiEH/2yTkTslZNgfF/19R9qB6cN5RMHFXCGzpP
xwW5eR4aO5B0kC7uinoLSxOumypAG+GLzMk0GptgGoX8ZYMOIf6wP24Zhnu+eqZo
tmEO50SXNtbxHvlq/l9V5562okMa7zKGenpNRbc1pe+zTj+ojJHtoKysd7f2vrhc
LzXQJVUkEUXfGn+Gh9nmUs86EBu5Oa39Zk3Ca0OOuLyHr93UbAXTHuPb1YldNZOC
n8/Ik1FowR0lHEGB7usmsqXcepw5SkSeTQ/KCLrEriDja+gQSo0qUaNGRXD/E5qS
hLagQwltCDRT1M+pK9MA9iFkjyAzBtwmAabHjimKMreR1ouiyU0pt4jTFVJoZAC1
wJmNek62dfBMONfwpz/p9xotACWOaDPln6Yjq1KyXv0V/Q4i2Xq5DLPGycxtYPlb
mUvUAqJpE5LSiJ7zXfYeBAiAXsRUFubVzZhQ5CTQuELhKXgAXxqwlgyt6zCpGKjq
q8DW92LNI1mDHyj0+pKW4BsvU3k7oBtzlejiKbxjm9SjRZhmYEh1aXZapjtUN+sz
D3cN4HKRW0Zpe7oyzRKPu4X6EkogLuskQnpdyLObVet24rbQVGoVcXX0DE4Np9C6
MBV6S4Py6F4pt7lvnKWhsfJrjPHzMYdnUHlkNVc2ZHQOYLUPxzosxKlNC6DNJozP
Zh49875szeptkMw5+4+2JZtG3VS5gEJRMPQRikVim/9DnE8JxDGkH5G/zsWmdwCF
904M7P5Zn7s0cPRDwGR32dWmPjC2YZaNccob48wn8sLVCd9l30tM28+My5NCbZ3a
E/FkF2rzfqcx37uwywCMOt82QCczGsz7UHT5M7cRPypJAYjzwGOKeiFRRj7IKi50
QNvuqnelzJUkRdSd/RG+0X8uqyh1zl/BuJ2addGj4cPJlURajRhiTQd9+Th0WwKx
t1N74+VO4YpK8mAIb7bWHMfUabXfOyKX5O1Ww5Al7oDEIQat6I2z7Zh0kfrq1jh9
Bc48CjBePZ6I63m7Ab6ot+h9VdXxehfnhlvSLY8BFNDArqYSH9MevruDoFjCOZU8
SL2nIoS+PGFTfV/tPbloV6I/SX042C2/GLjvFVqPaMktVJxXPfL/D2TiXN7sbaHS
rOsi3XUtvnydXQFit9rHaylUk+m1dB4RmLqhN+mvFhvpwzAOtGIHiDjq2JHnF3bm
t9B2MXCeQXJ36frkSvOjDEuzLCx1+2elghFcURf8WohJJOSBLq94FBayIwNtCf3Z
aLxJn2N+c9+esk7lW2Nk4PMAEMBeC2sZPs0xhctr3wW1wPnXCmjyZbeQIZ2Ecs0V
qCibIHNdi+AUJ7EMSM+AoC83m4NSIY1ZKLZhR+FcAwm/Ljhx438/yhPCq4bnUrjs
LhnLVfm92mxwkNEL/JrpdpJYMjyhO0Fr+RTjywXOIbCTD/9hsoM6qU8tBGfd/mfX
KQXwUOvWzX/UJpaGhqncz2j7gRQY385blMy+i8AT8iw9DsGTKeXQTMYu2u5q0VUR
Wjl6m/CS4vZWhNQFQibOIFUKMZstZbwOQAEJHhYo8Ri6HzmszWcMITSW4IkGtvd0
XiFUImfJ51DLuexioNHPAd61GEVX7vuy6hnlGX4hGdP0Q57hIA4Ad2nq/8qbO2zT
Ct9WK3PTJ9onS/qbz5cR3kBZsxJ+2jplnHOfwHTRTj4jdJXgE4ZhbD+cOtHIgHMO
Gj3WfAYAUjVfFSNSuQACKAlV7Z5gkW6XvRKoLJWwZOmI6GUp9DEYpp1jV/9x9Akv
abziwmnNTWBWnyA5jZ1QOLs37F/c2nXTPziXjbrPm7t7mje1frqekUSwig2u4h38
poA+7WFFcF3D0HPt31YaNpFmpFR1fPdmrVlZkF/HK5loDW5BzZDeR10/O87um4t8
rKMb0+CX9GVEQ3TdhDYrSXlMGnsiRIkxQUg5/P1hjgF/+MpZU/MpOQS+SvCqRlp8
mZhs2paHeYemL0HCj8leYOldwF5z+jcQhnafqkp1bZKkGAVAB1ka0daX4c2qXtOX
ZfLsMzlYGfcP1CUWGkB1wtm13xMNC2GT22sBV7gCFpeOaRyEFqx88hPEVT+8l/fG
d3fwZ20IPlzVXz6T7XG1Ri9V5a+kL2XydimsL4R3BtbwnypvCR52F3q2j9gqFTO8
DHaq3b+bRtnpJr3i/0Ex3Zt0Yw9le6GtA/bQW1UknjqdGim7C8MvQ/u7Siyh7eQn
Jn2CWeNNMGk4/MKFo3yOkaKmObUFiygWwcwD7edLwpu6dMTh54ZcwAKT0e8Wn60v
fOTmbpoOx4WJXt5WwzbWimJhQ0rkiVsRg3GxGO7Ui0DdUIvYNUtTtW2/KtIAXRqk
Oq98vPvlJyiB3oJR9LUmWnuZY1XqmIUSRMLmmzvZ27giFtLMfBK7LeM3MfcooAyj
TH+tn1MLkebXwclGTKEU59XgEX1UeZIWTOuzIMcIN8ZQIBeQUDQjYNgY7aP9GLyc
fXrSldQyobF9ZwvN9KFpnV98VACPKiwSF2pNU0yi7OesS6IvV0gKBPYuC6KYMh9+
27B09PWzOXuamCC0WGoVj2H9QP0CqnLOWZS53QdXeoNkWs0tdVFsFNq5VFE1crri
3DL8Y2DxIHWEKeT3Oq6mN+NJu7RWjsi57xHPH221En8RPDbfNzPrPdHTT9QBBHVQ
dtDcm8b1hcq6axIRVp7FQqwcIL4cfEepNUAoxZTf63sBd6Ccm4MiOAlccUgN4/96
rUSPOEOFTFCjZUnQcBFEq7AbbU5gE5PXtmGQ9gSTqPXzq5CtpvHpCLA8VPcG30Q+
nHfI8detULeov9JwIwXhSZk//xPtv3/lTkd6wXxteTaVl9T/xaeCAUbqX6wPLW/F
T9H4GiHMZcxjCaRxgd3xkkSutRpbBCVjOEXEUSsA+GD9NZw6NJcXVjsLU1EyKJ6W
5ZDimwyoFYibMneP2xREX+yWytZNQt0od2mA3sI58xwgv2GO9fWH0qovWKZgmm2A
SemxaQTsLLli9jySTM9DIs5fupPhBEjHOsKtGuY6QKBfLso0pQq4hkwEeqNeJ226
Uzsn8nlvQgSXLvSewNednmSS0FzPiQjusGfBM+GC07vhpsJOqccMQ0C1KFVhgIs6
xagqIR5TD773gjcGR+yj9g6h4qNbFRFI2ZdwexIdNIhdM7Jcb3y0xnmdCn1O174T
OMTD0vr7HgFo3sPa+oXIChNfHMcU2oytNFMjwvvJp1jxu3n0dmQiQYmdWvvmXrdB
D+fUzAPSI9COJkUh50mXm5jx3aw96Mj6PSt237mXvvjUdP8iVpju+45p5mpRH8rq
FBCEqzuWKIC7TF1RK5kdXMdmOUzc5OHZ0vSTNKp3aecbabPmwl2a8IQ35kSZYAj2
AgsrYWlk6L5Gv+syBxdxm2vv3YCdsKcbhCvYE3lXhPqdn2EEixcstr+GWWErXt8k
OsDUZUYCsxuyG/wxxY4kj0O3Ag+w+tUykVCWfbBxH5CsxzZbk0iZmL3WwrN7MnOV
6iepCqbq7kiYKXAhJVBsdyiGfTHfzVBiDEmvXOCXpUpnXW2Rlsjb3Z0TMzj2OpeL
E6Gv8ZA3cNVgoXsL2CCvpBe4iK9/j0nkKJat2v+quSaH8NCy1Pi5jSOxxRhyo22s
LjOjIqLYnbW1f3O/ffas4lz6zDerqIVQI8R79nfJXpCf4oY5ZhXe6Bj1/tke0iqo
kAraokms7kjlxrqcd9IjPzNaAvagP4Wtq/QvpnVGTyZ5Z/V+Mdp4ZeU9QSrgI32M
IpimsreoAFE+VJZsRxZHnwY3mMhrd7XD2+O9NsmUo8SXr+Ch4y8QJcNt7k0j3+9W
OidTFg6e4q9N/nnqCI5g7vcW9yWqQuVaC5p4XG33TOiv+XeuCjViRf+w3ZJQD+nu
sEDpMGB+Zbla4E8G4LJYjdASlO8JrgvEBu7k01nVcSLQc10w6zxi1BFZmhKmp81C
jhYTbefXFXkldzjeRgRxZ6OTEWZpZZrN2qs9UkfbX7BHZcjhG8w3J0BOZV3rT8hQ
d0mD2LoMfYeDGp4yEOGX9eulHFjqn4+PTRKSCvAdQvM0dU1nbmpHfRPGlOjNdjQ2
OK72bdRhinJZBljXB4GG41Vv3vE3dPoO1dENVR2tfjBxAhoWiVyNgMNYF0Ao9sVA
IF4F3qrA1677yDYDgkXzHsmNZPVkgJba7HjUQI4Omf4tB14Mghq/xS673/dZOmbt
BhkyVkjZ+haZoYLS2UcCjG08DOilc2uFQ6gV/TMVvoJ+2O6rN5zyLgowFjSKSn5l
SMzG/lAlPXZaJV6giOjOsiN7mgFer9mhKKG+wZPqsnUGl06JNSjjs1GOs2L8p7RC
JFO1eDxPoBViblLqOtnYCOYFe89P934VeeXaVWYyPT2egtex3XqocBxw9I0WJ/Rk
bccvlmdPRwkMCcvuF/Zx6vGS9vN7K6Ai1ioNK/5BAGqGZ9tzF7eoeaFOSvJXiaHY
xcV+Xs5IiuIKNoEf24phRD9lVwx/ZbPxfRBrJj/gXUK8of9tb1O1qyBuvP4tSh/8
WQMdq3tRewR3L3TSso3f0ANY/4VuxUG4Q7j406cHtLflyZ+4h5+VTHzFY+FCNDDo
7oExiGukKBK9p1tX0eCN0dsZyqbiKzw3q93M4BFg7UMwB0yRLp6dfKvide0SNGMU
YvPQeV0faErODwkYt28otSyuoB/jQ+l+iiTByKyo5wtpwakTVquSa4kkPw7yABWW
1d0/0BqrXPYWXJ34hpfpWqOiYmRRIsXDw0QqxQsWty/srTQwMDjMptpmDcBRBl++
Z1Yn70ZreBd3aBCxSGazO7tfGo2PWMAouW5N2euhXCdgTXBJWlhrd0u1Yf2t93+A
y+4m2A23c8FnuNeXv4lgHKEFWXoRB5ld275TTJ8GAYYjkfxYPCDucgZeDybjDZk+
j6P3CSU6Sl8gKScFEgirRpgbu+zq3k1m07lk2EPjVP/h8rzDN5HiKYhQK1JlSOnV
EXxsh7daoN9A+ODEkrAYa0nbsSx0kuhSKbNGU0DXiw3Gk2NJZHjs9XhDdq5xPV5E
kwlnQ46c1GTQA6tEG/SDQleSY4f8fpU34lACklESoFedkbDFzDZsVaNENY2CjFHf
SpYswTTT1VYha4C6ZcWfitbMzISKOS/vlgrEN66Q5FEkIRJawTQyeuj5CoNHuGNb
NhO6OKqDaZEQWdDwEiR3xndXURMvEazhjCmUdFGmiuiuO7qHnahk4alG3JjUKh9i
yNW5wdFB6QYKqTy+1etl6qqveZIn+LM+gTaE+833kkNBAasxwxl7NPGo7HJ7Mh14
wP2OLcVEVFL5KW5RNMc+NYyP8iYp2nT6imW1n+DUVNcsCCW1QeOU9EQqyQwt8Fel
qtssLfbLlefEKbONXlDWnJOLlZGS8cj03q8tgeQAOuwu5YcqyynTTVuupLf/7yfV
RyQAIKMJoL/Pj2vAShhZVRKvCd236ITCGcRj6wovFzcmjYEmejl6CL92SiXmoa4X
gJKk0LJ2G06vWZILlJuk10UjqJ/mXQkSxykXsDl4HVkqEJM7RLMJ6UTdxIdulZnx
4OC+49m7GcgxqZcXOGDSRxM0fKkqOzfDe1l+zUabdutwad+r0DbGadfux3YGdncC
UAamvAPpglZ6r5Un9X8WnIFLZg56QkRGofRol6l3qXtjCwBXQaHXjquCyvDQrTXw
iC3rdLJKYnKPALaubpZohmBKG03k+OeczOzBtAH11VOuH756MPTTy/EhNwWcnBe9
XukO26JHQtmGSt09RI028Heqq337vrGzTW6voYaaW/aIaebPEgNnWj2z0mXh4Fjz
6veKj6FaIbsPR9CihZ4tb/mLKkFOI5esw4weel/POSOv4bNz9tUiNULf2LKMsZvt
CDvc4yul9yTBBv07g/q5qhH7yVgnYo5wbkUuJZkI9asjEyBree/AieOdraZ5IUGi
R9sOd9cRvW85ttGilzmVaUexVx4awLJ0RIhYeryM8TXQHMWwODVaVD6uRTAsnhAl
0ynX06ZTqqslwnusT1EloldGT/4zfoZlMiOljsbX1Hbq9lJ43nkctih+ie2CndtS
UWHA9vldQH+RvNjvpibbGgC0AsPkAeprCza5wRK52qLeaUM/vjiDy68PXz4SPtpu
rD0cyK1BBTNheQrGO58fyqZIXchpgSksCElnSoKKJrTSrAthBFsdMNI7sMsn6JLh
XNX/qbDRV2MmbL+hGwlwei2i1+KcEd0+cAShIyWVHSZ8SiQPw9wlCaXUofuj2CWi
zI4NnkzIwEEQwR8dUICFJRoZb+r5ouInzsxAcmmYtJFwfx8+2hkedyIxUmO+RxGx
g8NGq6RqIpnSFoY2Kt3cxxT4abBb7ulhHX9E5bj+ZQ8q0zKXnLn2ztJ1k1osS4II
hUE1wwAaoP0rUIyKTZmuzLuro2Lb2cIADvTzo5t/u23BZdtrjHyHH367pmevCQQx
AnXMlnDeH+6O+xK0N1hOG9PFgCtDTIrXMRQQeSP+AGLEmCrMWG8NxmgoHnjPW39l
DMoauo66Nw1mqlzLNrdnGx+6f/SqgE6IovfAfZ+VfjuVBu7KMqhS+ezH9IdqCQ+b
Xm/VxbUrgOXmrYiIuUZNQzhSrfeo7rM6aASX/VwkzS5n2Nl+kWvkVavW2pHrwxga
6KSg2P+izpyUmm0X08CMjv1iFOqIGivtSH5kcIl4BdbQbrqzmO4Mo/QeY/njPGAB
SI2FzeiS3vnca1ApnWSH0vg1vW6S/blzuRlxVjQA347AP3zAr690ZxB9JXGFWVv5
aQs/uvlBanX2BmGXM9HT1tBkW10FusNA+PJCnLYYgeS0ntbdswmvNvnCvNZZOB6K
TdKyYzE8yV9s2hhUJjYY84eXSWEhKsW8IF6D4UcYqDda3BbG+xxD8tKwN00BrHbk
LbXZiTdxcAcapC/vfoXdFqt8I+/uaYi4gnaAezrEdtbNYn/WTJ0JN1UN5zTEJZp8
Q2LVAp5aG8QQFn0GJmfmIYSSb0alfkHgt3y57RdWiBcKhTXUriEshY0Ykv/A197J
I3oanAjBHPllGH78AOiKqhV0gVqg4lrWYa30Bh47vGs1/2AK31k+Lqlu/T2LoubD
N/Pm39vSWNa2GBGN/TwdLWR7j96B7M32wZXWct7/I+U0sWTc8I8Ravn3e4HZPgum
rnW7qrE54z02mpDOOo7TfU27Ughw0WKusFSFgqSb5cq8+4PSzCQ+twXKDMnSCXCH
S4nkEpQAJcqAOwS/R2PpRwltt6kK+mzIwITYf579/OqSNHXO7s8pJcLeI6hOT+UA
9SuNAn4OOm8KKal2xGAl21m6Xta/C7HrItXIzLgXL1ixfdx8ODCw26XekgaaqmbS
kiCF4NE6f1s7SOfddWThuTqmSEkQ74YDc/u1TX3nbqlynbehwCLrK2sfpSMsomUp
ysxJ/nkgVskpNN7EB4iJ2rl5FxCz1nvmo7gIbbzgnx4K5xZg2wCXzaD4XJ/s6mHu
Wte6qmxRhwSxQdXjgH1gk+YDXrCLEv1iNr+kySNRk55jZFz/eUYMgM/eZnJlHCSK
Ex3lBt0nLM7YNsG8FHegsjiCz5bHEsUTv9rhIYplo6QtNfByyHH6Ery2QJ84FDjY
vnL0Fk0VJXTXZ1irUGElYhOy2WnsHNbIoA0+Nzh8OSgpTvQVwqofy53tQizFmoHS
2BqeDSuo23UzwsM2t5s/5/kSJK8jVvKod8XP1xn6zgfRvzGG8Zr24DP0zm2MYq6l
gcqkzsD8sL/cb1W/Br/fE7sfv2yW3Bl2mUnzoRN65F+mVQqDJLUpGFctdpo1K5fu
6td/lls4NGE6DNWHFVdjdf1xqwoezViFvPWA21ZuFYRjHdS8ofq9HeLfu6d9Is5a
HQCVHttHJkdRc0ZsqsLBDE+GfAFnTGyV74cCenH3kGbxUMylzE3xqRhixWY++Hwu
h9Ru1E8wbgWwsvKkWMx7zrimxiYjefOCHZ0TWdExEqFuC0KnAkttFLu1r8v63sI7
VeOL+DOcH01mc4y5UddLBv/9ICsmQoNuRBooZKuq5vxoqT7pLzQHwD4JcFJbRrUA
yAlsUS490ofJNoxw0SSs/q5H2hZKrT9Bt3Uss3mriZ4XjOSNw/Yxo02yWr5Xl3nV
oU9MQXy3OALI/Vo2VvED07/479COQ0ofEv3cSDz4jyxO2b0r5h4mZPeKtk1twYZc
u+IvfrUdKeYmy1LDP830ABc6bPl5pyIfik5/wa/9GuXczFilyhI2ZwuvtlviKiIo
4mRWox6A+kYr6b1f+Nh3qcJjAqU0cc871vx0NVbbM8lQQEOFi7XVTLI9S93mxcjF
GnPkaYav0tSNL4Q26QqOVfmURAFQeS6HhFWTAI/xUfKA7I7xapbbURkO419bnXzD
s3SHpSraEH8p8aI/mWaYj+63J9YC59JTMHjtBJMqWlcEfXSoODzRJuTSo+qmda3C
yK2OYxje5lZZSrFCzEc79cZKXE6Nuw47YtF0Pls8LC/exBQ7MxGNrTHAI8PoO2wj
1+BDW2iQ1eiRMumX3+NTD27I4tlxfmf/I0FQVmNKXIJjaQmur68SLsd1kXZxvqpO
7q0f7AOoG1CWt0h9mI8gjTjUFCj3j2TxoWJWi7r9Vp3qR31UGnVHqSASOUnth00E
GY0vrXqmtq7qZ08zXRPBfZ7wB/K7+t+biu4Rwncko3EdNUGiuituNMEV/EpO5fGI
Fntc3TKjcJV9bsax5XUn+rUOgsoOWQl0KemDzU2bS6I5EByDB9uwuKqw5wZ660nh
MzzzJsWuKUXIb7gEUFMgJVl6sVJCOZXgmPNIKjdrocpuIl8KbmsCP2tPhaONt8Mp
80ZdROsXE8xzqQv9Vwk9QskO7//PKfAI4yKt+AaHwsZym9pD582VyEuzEc/iiwn0
UasnC4CNhiB7Gyhyald5XJibUnSIXI/kcjU5dtfJlkYzUlrUGxq+ghhVz/9uvnPJ
6g9Y1DIsZMMDs0iry9yR9WVodfKRjK49PVaGWBH5aYAPTXAMAiGH1P7tngGqMP09
znvEaCJcVvzIwI/Z1k/whWYJs1p+z77i0QRP/1xRPUwPbV3PEvm0V+uNQ1blPN73
ucpLVP+JVHhBacoCN4WMSzlI5Cl4QYuFNjuErSQ6q+g68olJKsV5vc5425EL4v7b
vDWH1Ck4dPfXOTXsv6/prrMRbcMjVeEzV7gnqAvYl3N4DG6YF/U5rB72A+h+vy76
R16uZ3cOf0KlbeOvWoUfDve8FRXAA1KRYQsSiB+FhOUqpbxfI/fiKUOLxPPFTyI+
JObuH5eSUPdaFuNiINVi+KHcMccogFkXEeg7Np8LIxMU9ZCsx6rASo/kQgx6GMZl
1I9LvFWNGYsm8TEwlgfvfSfkECynwfycXBBorvCD74fRzY91Gt1Or3u4XIRWZoWK
mASC4Uq4iyS0BlUsi4E1JLfqsKZbjdZYXgCqJ4wHR3iquR3Jqk2UZri0qRRNq0QJ
RYp2ngEjmbYiinOoMzpEMZRF8rd3obCfSOl93rKUw3XyrCCgenkf7xyFnIV7SGFC
EQnh5KbWuOwYoKL22IdbDcFNP546cTnadtgV0vYj2+YbSmabpDXhUX4BDTGIaKCT
cejc2wbi0Mwxbo3RnukvKNqooyhkBAWxoxSC3xItgp4eKA959q51f9hyuzXJwmqx
gQDzIfLItfAWDzYTfPLzMyhNSORh652wJ8yjdU/T99eWwnz6oyUjpHr11e70K9kS
H46+rISM6SalwykpGJJPOpPSOxmhDNixzohHZHJem/VEFVJ1f+YLRAM5JYQ1apGf
5QVbJwMKt6tSZ29jM08RplkxUYG9f1NEnuSy/yszCpx8abJuxXUEcJeuNmXLdOwI
OfjoYVOgqghiY/M2g6+b6htvGtSIbl2rJqC2OCcjZsWWozBpWhe3jFRNjFnFHQ6C
jwkCTbgTJn5or9lysCkGnEouF9UuoxUHp5afAxbd0eC1jdmvyv1GtrF3Xcyg4eAT
3JdBOtX+EwkCKXrNA3q4CUbbVa7JaY0YdEXIuphNT3VAOC64LFAZeig692wPrYTL
kYhPa/VYEDHn2Jgff8MnIszreb7PVkkImjdUc3wMfP+0PSwa2EgyM0Pt34GAkAq6
dlWT0QGABRfvwDokdpBelZkTSGEmR4Pj9fFwD6qV/xBbYsBYXG9FogvTmHpSEurZ
W+YJBkLooQiLFbrkCR4BulIW285P3ByIqQqt0HgCz6HcoLW8vslM6m9kCtOs3h2R
Bz0G+FI7mVpUVXE0CJggnpPEberLiyOiz3LB9Fzb/VkrDQ8hPp52jH/PZx94ZVDF
VVBxhR9zP4SEIfyx26lezJ1MUXqW1MtShyznp0cp9JndLGwnPS8TBK3EVhaCCWFz
iyuvhRbj8aNp+FIWlWAJMQBmQ/npVXpyNuw1WFOsjdwgnMS4n9uXRgLJIaOWS3Li
EEKvqMpzMX6QdwkTm7Ah0SIFDv62KqM3ShvCUCMFXcUbz13Vk5qfJxVgl4Xxp9F+
IT7a1jCTfxWY/gdiko2Ou0fAFKBklw+BDUekuHB8O2Q7vL345VHVtUOWLGqrE3qH
no/JiI9fAkRwtYaFKXDAKd9e59CkXi0CVwijUp3NnKEmytf0HgV7c2wYXupYx9bq
hGuvk2vxvPTwMEV+/D3TapFVyGscB2LxNDlH4Nk1SK568RBD/exaIjw+7V46pnDI
kBPRUiNAyEVA4hin6NkcIi7tm6myIl7yY0vMp72Zp4bsv7txVMqKP/vZAdclbbWp
sYvqbqquLpNFDRGXfxRj4Un1LdcBy9lDkMmUreLSrmy69/e7M8uRSRHV9NP4cfC1
TVLONaQodVxSxfbIC3pIkqH+a360W6/lDyrZl+ZasR5WB6SxGVgCz50DyTmcNoO5
pNYnFMOhmyx10KhyhBEROeZI+jbop0asoL9qjy1eDD8SwHQbIM/VclmKOfNAvUns
9y/viFfMkE6s8mBUS4akcm1TiHEC+RsQzetBInUoj+TMu2EZUMrIOfYxjHRQ7Un3
6tchGbjP0WJ02pqPt/rKPaU50OvteYWC0QTcWtjTuyJHS4yE8hvwOAin+U1kFAE9
Ixa/ok/mOm8WAoV+RyPjZ6mZER6gB07zHJ4oBdsop/v+YyWy0sGYohMRooCa4md7
5u6akFvEnROozvbPadwFJrYGDEUu42MP9bM2lmrTUpzfgOzvDwGvREnSEN57c/dh
zzwKQXzj9gpTke3YQw1AwdKK1bAMmkutEOrSlnTvoy0SWW72MJehL7rDXWOK3KiY
O3suubZSu9zsS1iUydVeq61V2E6tLoeQP237pLpnAAYGQTNF/rACeodNgWHsO5og
X11gaLxRsuN1yJvjQPbadBGIFiNlvsPehmDR4edeqqh7SzUQ8ZlaKrrXS2vk4LSj
FvQeG7O7M1dhgLNfvuSVYg/jPqMr80Mvl1Z7b2o11XODGb2LwEwAu/buE65MNUTu
utF2k0r3kd3B/5X4EWc+3YVR8Wm2ECr7gd8yCg05dswqPzMIj5k6SXbqNm2ggr0a
7AOLAII6A41w9cWMVI8qQoSDkT0cch4URLWHTQVt+YnhF3/2AmNkESwmVjHyC2bh
2TN6+OT7txreH1lNfxLpmLcch9Ywj5LXzKWLLeCLQraqjiocgtBOIFI9Ck1sf26X
2+hwiuhQ5VHU+jK4zaQr/XDk44f1rkVcb243NzkndLHarPr/NPugoeu8UWWT3O3U
+zdZ1LYVc6vcwwLv7Q/njJbOZCn/jWAhC4WdM3etkatrqAxx0ZixdecUaDxsYFuZ
Jv6mx6HUAHGpbnQ+0Liu2fWq6vtRjmzLOErXObYEQFJ2C0ETCEert+1KdulcN+2V
Na0z1lIPdqobtlG/XGqRnjFLtmj9dDoNQ24XdQbMlLPM7ydDK9RqEwdEuZWrzJmg
zhSuTpHBtjvzUJyiborp7ZSBJusO90IFJMn+EVaJKEBwSIEC5xu/YcWdSimTQRU1
uW+es/qHfhWV8BwQ6OxlcM2T/oK5F85WXjfweAb9S/zSjcrRpGyhD0jXwHsM/zM/
lvrLKDhce+aAfsNEKvW6QXN2KullHv4xqju4q/tEFzSEYG4r9aW4p/Xv2hUhIT08
j97mNN51wzOe+gd3eMu0dK+WD3dCvubFY9klxQDYtOeDgy/8t/4I3WWPgniHNxds
G/pqckx1HqR6Ic1vs1dXj1wUfhnpo1VOTDzaJTf67Ec+YnIRTEBbZP9jpowhSm4G
kLp1FVSYiS3gZULl5HPHuhzIS1m4/uGbBpQgf7lWgaByNwKmrejjwINkpMvM/m1p
d0F+jfzxWbRFtuFZq6dWkPBB6DRRKf2q5HVtGQ6bh+uBQWovj398HD62IZBhaZqS
ktvw6LLeaHJ6aov0tuuN7saXBJ3kB1YI/utyMyeIWX4ZuYMy/lm1PjB3cTALr2FE
iS/VTO9EbYpHVyCxtH4mZUbc9Z0GLRXOZFDySxzgxrjvy0SKB3Ed0cyCjgirsfre
vNeliyQqg1Lvb4Ai9TsVE/GsoH2jAN1bz1tJ6JIQ9E3yDDh06rDngeneMtSyI07v
BPBY+bdswLXM8FGANNzKQWxej6pG2bDY4ux51NPydhu4UIrjNz7LlVv3tYs5PsKY
FGfD9iuZJVCL3EGuMcKpiTWeBxzYRAeTogoqiKK6xx2ctPBmaRbkQ18cQVMGq2/+
1bMd/e9kh8tb2+7KV6hsnqXqPau9+AF/8pukoAiSMSyjmuWK32rcM7IsNZcWk2DU
wJe3Vp7aXWM53Bk7uwGe29cI4PIH2QqTnianaGS3PzRtl7lqnXgKlTeyIemwYlC5
AtburA0sERfRfjvyaW4/YmhGag7CLu8y/sl7CdUJyh8wEdtAbMOBOillDdCAzo5e
Kcat14ZUxoA8U22uI5SkaxHyChY8sVWVTRAcWmnwJ+RSws4TgnLG/vyRxlSvcUHh
yhd0Py7OjOiTPXFxc9S1luheAETHMYFSIZasOmY+Jc2ZY2Z5o+3m9z4QS1vM7ozj
2fC5QYl+kbwmhLIYGeAQmLobsDoQTNyTuJNPuy0M8vOFd8hIndaDYZiC7tD/E9Fm
6zNBlfnwlqgq9TZOq6W1icEgTb4isSwQ7zv23SEa2hiGTg/p4KnccrJQEzcy/DOx
OhJQ7CawXq4qQDfOzXXCCp9Jh9rwLtO4irEqmZMOJhR/wKKkn65PNSOYcFkNV5/l
4BJzYBU77ak/GtU2o2YbyL3J6dUW+cfAxA2CAMgBRriJR+O4ZvthZ1oumBjwUEht
nQf9HiJYDSfBRdBdno1RgO+PaJJ8TJGc9lZvnXcTFgIeXMSZyq8wvtFsJfhrBtj2
7mEiAGRjXiMzutYCF0G3GveyWQ3tkFCaa0K3BFIO99IhuglMsWH58mL3g8n/mxGm
fTMjjuP/nKJRZyt9pdbxrHjdf3JR/h7AoBP/wEIIwOQqo98hKBLJgqclgpeX+1Z6
n+IJcyfPkJSM2RMjlzCzCJ4GA4J4u9PANa05E/qLrO/tGYPbVhetJX+oie1USNHB
cjWifhxQ9DnMdLBymivFUGbQJqPioEhD60PsC+sSh2f+iPxyP+VN0HyM9HxvRU6J
MYcGbj+HKP1yfE+FkJk+1yyQa/6m1DHydGnotz8ssbWjQt9freM7sQRTazGZlkqD
Oav2ngc7wM2U3YWTrDoOh+7iGiaCWdQIpmOXz7xH4eQl8JNc/LFxfjxbNgPoTV8Z
UZ9CuJ497O4LSbHnoFMDcu3c8F3XTPEAg9ApjA/zOTIYAYBPCQbggMp1Alc04Hfw
5YGSy5jH0/3txCdkNj1oTF2CTgpG6eYaovOl++6MdUGpU6xJ1BMUTzBsvaf4mXX5
4s/I3OqwsWZpQsg9YFKOsl6dZZQX03pquucIeE1MY03+fgi3Ub6q4bOoHLu14Phz
n1Lx8/95Dalk66pWGlBteAv7io6VYABg3s0XFwy5ggX0ckzZuWsxAH0NDyG1AESp
8tnoVTslAqBrroP94h0bH+hruZIPwLA4XbuIUC3q1Gxg4fCHBOzvBG2xXbnniS4F
jdKbF6W9IrZ8Ne38/JGsEoksoDSXwJuMH3beqcmu0eS3m0Vo+A1Jey4SpRao+Gpz
9B1kvWL67ds7AAr7270sztZCNzdvtUKDkVH0TomyqE4HGdoTJgKqsKKHOjMY5HD7
qRhGqpjiwA48aXY/dyEMV2FqQK8pXo2bJiBEAShWK93ZxjidNr4HKpR0z0hzCbQE
tuulczTQG4Ox4y5zIUtMj0CbwqtHbFlSYsU0N53uFkgpggKmFg4KJot+0Hflky+B
JF3scb1FrvCRZCpU4p5SDF8vanbF717KrBm+v7e8I840WinkdvWDG+FkwniBsVjl
S9L5pdvD+qOdwUBtqlk/MjzZhq41vV+t8RHXxn1855Fcm8RWaMu1BreEDu52OWX9
WQBqdOS0KuowQcZENqA/BbMZSjGtMH5SExlq535M1zYE+wlOhyLCkWLisZJLvs82
JXxAHbrSsMhKlCK2su9jjkputeYogOKtxXjYRnBX68wgIOJwGcNqnd27S1r9fx7D
JJxgkf1CjGM79CV6mJ9OuVBYTrk7YD71WYmxxwMZGo9yziaA6HrZRvKf5l78Kbe2
k7PMCCU6LAKA2panflcqdl5G1Yhmm2+dYFl90BgaKsI6mV9wNTGtMcPfSUZm3V2l
0FOp+V3Yb7urZ/LYgMY6k+DpPIycuzpKHlYW7OqK9oA9pb0kZmXScbhxram7qAQx
u5K1UtF8sD6rKm65HWerKAKTwrfVaK/aESZR1vHIn9oHsgNp6zgCYCdcrIqBhnbZ
SIg0YaHTAAhscosGErB8C/4BGga+V7soxoBocxuXPJWF8TYbap9kVv5FTzcCOQUe
VE9oEE0RcubQPXJ9NqvWe2XvTKiehNtbZj1nTvUrWTfwGXtc7DRjmROStEFj+njg
0XuUl7CIcuRr0Hzc2WCLFrJQqDWfUOhr9nmDOvupo9arKrXhsisJddkC0AwpHvpQ
M3hGjgVc1fob56C4Wo9TR8rlgBHYE0Cq4SnMlk+xisE4gWipId1gyMi8zAoSTg3F
kTma+Cde9yZle00lej7CRSeSN50K5QnONb+7ito4lCcYaqgeJSzYJIr44zVxohOB
57JkM1QZEI5qafKcwmERYN/BpSDQ8cNAVkpBrizJPnfUxPWxTqcict4z3vTYLSqF
fEKgEH3GVfNRTambU5M48O6z/xHr0c5VoWfbtcn6IP+cNbjKKvic4MMzawQSbC1V
v+jOtwkj4Wt0aJwZTV90cjzjZX2y2nWIV/Aey5UZhWrRtYpk9ZprNgAloRjYeAYt
jXBQqgpIMPxTol/zXIv5H6aJHz/09oqw3PBRSrFmInybTBHYOBQ7SRf5f+m5imim
Cx2YuDUhQwOTsgUNN+lmIeRFCciNoJiMnDCSxuXvh/GnYClN/eK2gm1ZmtlVbSQ4
z8yBBL/mGzC2wwtRnOYo2wHFBE0Uakjii4MeqTOhViGyk3ARWjvk700XJl0VE534
00IpNDCXUuX4rFFR0KL8m2mxIK692Kh/jLyse1rbsCVfkPXh2zlC1oyxRK91P8re
w9gqPbDiv1SrG/yDwPdI7XjJ50JbHJPKGzi8yti4ev4UjgmgRF7XfJ6BVd7z5RLS
9ApuYpC8xfHX5Fc9aLgLh+EXOc4GfT/KUJXnvR3uaHxyfDjGTsGBaHduLfzeJDfm
1zJvSVnj5RJyA+5bt5i3Se899S+1lUbBnQt0CMQe1WZ4HGFhPDe04OFS9A3BEwWY
NnM0EPb7TNaEMqoZL7XopYuf6wH3emL7O5y/v8imYtt/8g3qy3rEU4BTT0aO6Zei
b3EkXM3CvGYjnFQ+n+t76STpex1I1xB+0ywDWnSAYtZXcaZAvKC9mlJUD9RWDPd2
sIx0N7L90mu0z3sROnXyPaZ2TGBnXQK3FxsabftXkgu5R2pUxc9lmoCMd7zvHK/1
i/TL7vnClI+mu7AqnxpdnlJV8coPqC3mj9o0T8oA/5i0L6BKUlId6z+vW0psenX9
sVsDXICA8IiuRBIbl9dHgYxFEXWXjrRJ2460XGMu3kfaGmjola35G1Kqnr7z6UPY
NPPuf9cylozKjmWakdh1uirBJZwOUgnHxrHdgZx0pquYFXi4Z1kZenbcARsZV1ng
2Ul+mP52vKVPWIGqNdRb1Kc8Psf5nX6yDfOG789fhH74G2tJ4TWn8ET6oLNNVR7B
wIdfq+7JJSKQPp2Z2Oa4eDCg24Xj311Es+AwaeIMxeFsBBcoTHd1Ye7Ly3+bSSvz
++LccDZCafCwuafkh7QlEe99wQXzf8Dlo65pX6n86NoHSXl25VSrWKSvATqEXA0z
OZBFcjwUhQnNx4pl2vlNXthXbAh5R38KzNdjsWftxYlaxiUFdnUzUJ1hvk/BsRLx
WXXM5N0YPmPQlbgQ7w2++PrVR9ee8e/LFjxKuthbOo6wNHmVLE1rHOV4ORuJdan4
hPBrIGqZap+3dM5/H3xICzQo21XQxnl1I5F6OqEDy7gjdm6dkc1Ipcxuptg9xGn1
xyH51s5t8G9KRbapxMkuS9IzHf9Khc0gUHr5hFpw4vzd5NEjwg6dKxlAbFoI2/lV
9RRABiw8+6dFpI+BJUUleX0I76WCvt34M9wm3XW7fGMHHXqSnlKfPDqrubr7jQ5C
03PrheJfzfZcGYdUXk1uOJv2XxP5juHIKOJCg+C0mTYVelWPKIergqDEnZs2wOcw
xju2COiFfz1jn0sgFvvbJWccQYZV3PQXyoPP3bYiPaOjxlHo7Gsr1988x6fggmsF
3FuABLCR3uG6zEaekUw9kKZU3CMIhJ/5mWAL5myOBbAV17rrlSILD17STD6R0xrt
JsGjEDM5CQQz3nkkS7XArWaU6d5zrFT84t8u8Jywh1aCt1CLf+QLGuHK63cfDQJm
CfWNRAJFpabytWsh97aEBthPLhe/0zZ+3VPmBSx5OHUfGAyiTg+4h6bi6IDublFS
7rBWi8oyVVOfV56aZnvxZM83tmAuBjSxSgtIznQHpKcdxBnA8SflAD1DqbH71V0l
a661YQjGMraEWOG9nhI7d7Ue8ObMGNYxoyB5yndMVGtn/MIVZQJjiL/2B1dpVvnk
WlwVwYdBuWoVDbaEAXUjd4lEmreOT/Q23ZHM75ffs39kdG2bobLZTWPFiNdM3Qjz
iRo+UmYERnnKKigxFqS5maU9DYQEs4vjtRdJKGqgwnUOyHCB2g8EjxWWtt+4eZBP
/BIOHZ9nrC8T3Lss49WSjmpDBFM/tmCrjvQOIWvO/KzXnw36dGgtGu00naO9pC5K
cJgVpE+YcGUOu7iXuBf4Y33ro7W8OmT+seJ1R/h6bTpph41TnNgcY/k2BcLF2khb
SG6b+73Q1gOxnUWNIc/siWKJg4KWUogWhyCrcl9MQfhhDg1C/iKjPT6/SKJoNr7b
3BZXkwy/B5D4iUm3QHv9LXJn45pMfJ0GzBT77sz3+AWmPvUgsAxRA1rhOxynOg9v
ZWrZZyY5QRXaavLH1GGHV8367hIwPsT6RdQ8w70dmfhBw5jYoVsv6F/bPlHT+sOq
yMDNZR/Cc1Ra/QnwPFKIpYtwM+xUjX/BBDb3oeQWjCYgQGFjG8R1KQOcwLPJq05s
7g3Ke2qGzehk+V3ouRtW5dUIZ7N9CxHBDtxK7gskDb8+97Ng0l1EC0bL49iRr7KC
PhyrWs6eyicAaLpt4sgSqk8J2Ae4NOHdcgtiitw389BENpPL5QHFtQ+sY4R4Xy8M
xjk/wNOrsbn+fqyIoRgppfFN1Xhu7kCHu2lowufdZvT5aVPW4NOu2P2RYKDCjbi/
935xyOdcBs4r74h5gVPdDWvpj7gk96w6xuebz4l8uwzEN6pj/SKRazWiUT9NeFok
wZTa/NT1O0L6cY/ID2+oVJ62ahJ6dmF//njegt7q3XVWtlqlfCRHu91wjo1f8Rsf
5SDWM8L5PcZDGDiz8GEy3LyTPlPK7tx3nKM6iKhKkPOGkwzdkRQ2Nta0b6xMDdTL
G62gPiC7VGYg5KMDZUZoHW0H/AH1b8j8Kgv4lQC765z9vofZB2ILi0WWN18D0a0Z
Vl/Nyj291gzr/0FK9T2uk87+5qbOTvkKHxbkF0+djrpdjgszgltrNX7llzFy7ISA
f/GNv0qzvVwIkX/AcswJvk1dsHiUFYANH1Zkiwv5MrLmjra8q1kTcIzHhbGrid+Q
6I+iB8YKinTDXanBXT5m2iLS5dVkMcYV4wZ9IN45b8gQd3gkMcPwniw6KZkZRiUv
B6S4B6w5grG+uEylZo9cykgXuaREWrvjYKU6DvtZ2LrDHbG1R9k9TkXFOWZKVEJh
BibWgEwPnuUwQ2zMr1i60M4quV+C2mX1vuWEw9RWYgwd2qGSXRdBZsUfQZT8RKXW
4jenndgTw1tCoweVBFrVyRtcBzIFQN5Tj6boPc2/DGyUu7U8+VIislar0XkSOD3e
2zNPQR37C63FwyfEhRU+1APAr8JQc2swWANt7zwYq54ormmRDD7A/c1ZyRPLI9jP
p+isfAOIAATqYnWPva/Xsbwb5WIPN/8De+wgJ+UVPUneQujaDJr6pFydvSJJXEh3
IXXvPTRXO8Oh/dH8CUsUv1glgbee/r3lhEmX3uKeRpRqjYUMc2G+fTOpk4QMn7NG
IFeUX4V+s+J/DwcC4JFuvslequ7cjs0BUobYfgcgmtzjHxlxlpU/xAyAUaV1GZBv
npeis0qCOdbjzupjnSruNCx57ENTqfPgUsyGjVoRRCoRDW6NSLHgq0VSCnTJPWLP
NEO5UxX9SRF4/yXZ0TqEDeNt1SD3LNw01lnXSq5sfy0Of3+nqh3NpmAxFYJVDiq5
UMiIPTap2ff/B4viziwx3efyunaO7x+WVqY15c+Bb9toeki9aCf3onnf50x38uFI
xIZfbznMTBM2q1Mozhyo+AAkgjul7PxEZst2WPlxjVpdX5Uz2wZ27iWXSb84k3up
U8DvlFF91Agjdu5q/lyniktG0J8+NuoGc/MNOuVBOr2g8UcAX3tIXxSrm1FUN/oV
1XrxfAnRMAC9RcyItBwOHbn8hi5Yrooeu0njOFrF3XAkfZMqhhEXz+0sYpCpwyov
mu5VbzmpiAVhVGD4xZ11+qBPdjFqE0xmT4YREH/DmDRLQu+sk3XbWnbqypsc734U
BE6eAd2loux2EeLbXJi1ygU2D+myS2xh8CVjCkRQm/zos2gQ2eB7pCv8LDKRGkIh
0Zd+841JBALMVs9XPFY4y3x8IwnnUwddDb++NwteyaIlr5hHprzfaPHFQ1hqNCp7
hrs2HWshmzXkpRfISq38angoyLJim5FHsrFkwpnnJ27OyZQPo+Xd6ezG6TvXC4T5
pnEb+h9yU8b6ptkNXMKPMr1zF9iIg8a38JZ+c41U317nmJwFO1PSKkJsHap2Lso0
2ydJYZ7m/2401YnccnHkV07zKLZcWUiw1NqcK8xF6hNNtoYaaCCkGApXWBj+UuQQ
JeLOBgYjDccGiU6QC0Fzk1ICzUAd+oBKsWaJfQ8OnXNfWzOLgqiAA/FjDn4x3gFt
xZoMMaH5X14CGL2AN/z0Z+oYNS5Nprv4skXpQqTzGSttSsWLjGaxPODzBJscnBGo
/VgXjPFWcewnZZ/f/R/rfogHsjftJ9B9DFZLC//iKlqQCiThzNsnhpBlitiFpjYO
R9NXnuidZR7yHbgyjjrlbntvm9XeZcsbaPjC/P4Gb4uHVCs9K48TVyYXHWitYRO3
DMDkmbamSr/p0vgokIBzs3z/2M1kxWWts7Zqu0Hci2Gs/yesZlSnoPWLPXAqwuZO
7XbQ0v/LWTrSpuFcU3tyuvvhxc5/8z403yGPRx+Vd0afJU1+tTcg1m8BAnN64KNu
GEVLVa9yOE2PaqHtvC4BbmC4pGePrwQTGhPe1wSdruXtQeafGC3j27dTbQ22jbJ2
In63++B7lqCaT+LXeL1q7uh2Hgg9vjm30slD8vpZmwqVRKHUTVkJ/MVguuriv5JG
cQNYJP3I78vxYfivXMM/gu4WffGl76kFkDcOJHDCjimdXH0FSztC2WG7cZGGMESh
+bhoGEOSEL7/ZgunZw2nMgZs04TaX0fww13jdsU1utSbzB0KSPaw5RdBFnyzDotE
FU1wX5dJB1gMxnszdHw3s3IGjLcb2oy7bRq7fvTw6Zam9m5aGdKY9R4EkqqqnfRS
j42D+aGbaO8ohrD/NS43XXUoAIorKVPdPaxjBTZP7jM9BFw4lCYjDHZJ0pAunAbd
oXpiTVWnEsH5CVMEtqx44e9SciU+I+xt/6GUF59wmNBXYXFK1VP72kT8OtKthW8u
Fy2AnBk7AUPUoc7gtDEEFeUceTgh/7zI3lWXY2ov/bE2IcsuzHo8v/aoR/hgq0zX
L3dXY9IyuoM2wqmRNeXW3R7fSkrMUG1PBVFsvWynu/OMf7W/9I3JyFUZ5tzC7Pbp
4Y0t+MgzfuLKyn6I7HdJJ9FN9ob/PPcNsDb9CY3AH3l2wPpGmdKvdPrDJ9Fq4uSQ
0Ehsr66fGMeOWub8W6byg50Pv/sU5uXnyzXbvWYILThifIyapaYQeOrWOTJQgr4Q
cypMIo2PVyBnw14a3zVFwv1P8DOCir5b5rZnQdVdjdoYDh6y1+2iy6ITCD2fFtiF
XZZ4zV4m/6UK0iSjgdhXu0V3WXP3j3goElpePdCl059h7DcA7HZgRz4m5uW2Ctl6
Z0cfL/m7+XdvBq/G0v93IDfzPcnBLHEbPvAk/HbuzCl9knwlWm3STpKmkfruqZJQ
b/ePs5D6/bKQNMLlyFeZ/DnVrWoqf4hBbzlIYdpB4WvYpp3s0FyMsghszykdPn3g
fp/eO2hmxU3nQwzVKuwN85GKXdGCmBy5lOjndsZHQVhDLrYQw3Qlwupf0pHDIURm
+yjEmF9vdsBZepDIOcH0GsXD72r7EbhRuqykepT23CWfQoStiESVkFor4u4mG/72
PsbLdKmwydpi+LNXcEcTLj/5nV9vCqi0nWMfLJiA1KWVET+8XXk4qWKW7u17GaFk
y/1OSRBUPFA2hHblmJyPAQCOYzB6X0gumje4bFiATMQ26+vOGe8WYrS4fPJSpjpW
BQsTJg3n6x1VfvgA4jiakZUOtqlgJ6un/vmEKqlTHEI+CxIhz5J1iKBaCmmpbgae
gtznmmEz54KfZHpG6WcV6sucevo2HLXcm0Mlxr6vzld67bTryGf+D9g9o4sFDiVf
E4nw3yEuGY1w3CAIk6qBu6eV5abVVtKrFeN+pqS7U6rXIDFzc/P+5jcAk20jXHrA
Wz6gQsVEy70RNyazvZMJfxDXT7mbTDa19h1kF5qqqg/0eX64ojH/Zr0SeZiKJoj/
/z2NHKICOnhvbQWMdV69J2s7/Jyl/hkq24DqUllxRDezMlCGVXp7lzWoie1M2Rzv
UBhdnrClPJ9upEDfjf4tpvti/c9SD5WUj4m0zh/b62FZoX4KmLNbwQ9qGEU+/GnG
+G5BCuhTt4AbmiuBHF3i76UrCaYX7mYb9Ho3hZy1DouKomOuUf20PY3+/iUAiE90
/3nDbXVB1TduiF7uFZngMZ6r7fn4aFnseuiNkHvsC57unMqitT6EXENwbRg7X+1u
wbpM3vgXEtzymvZvtBZ1T/1pmWMmvzF75C0x97SAiH4iLMuZBXq9ADaBS+8sainm
twNdoLQ2bCvEzEw9Iyd8sIG9U/snpWs1yLyv3wwCjG0RApwxFbwoWc1KXbbArva4
t02gh9/KcPaDcY+8nl0M3lL87gv5R2Uupb4y+OPWq0Fm7eSRCAJ3vHRHny7oXzFv
EE0Vrr60ov+40kw/NIbfiMW49zqOXKePPSCckuOOJzYSdJr4I/Zw+XCWYQ/RezJu
nn/LWONe2g95bQvcP1+2RuilhrNLM4f5Xpn0YRLVIC+jJ+SdeGfGRmOgL4B7GFVN
VLAz7SNj+u7YhRUqeBbdlgun1nEWM1fe0zwtGxLnLoy9PsNcG5W0OFX6Kh8VUANy
R+obfzizzYj8lRW/W2pvb+fF/P8ZztxGSRHHJppK8oOytEGTGKN43dmcD+QdruZL
HLopcit2mH2shPSOhIiZ27cONaBV5R/ar4KYhXpVdOgmul6fnbQlp2jopRcRxNul
Ah0KoonFq4ite3cnwZ70hRsEXw7OaSu6YP4RWO5d8FxQZrJLX1UfOTOVV+AJ0r79
v+nBahkEaozMqXr5boTGDwrRu3YJFWXjwlfvXlLgwi8PwxnuIRXHR7ls0q9bfiz0
cegQ6cXvHH6UuZtMRAcoxSBxKWP0bxiRTVOoUlQAKghj0V4/xUZtqGy3lQs/Nzxt
tMZFfmCeGbvJnSoiUVa/W05QebPh6Byq2jj16ERpkJMXxEoZ0odK3dVAAjSjP0Pb
ma3hedkqb8rSQgLp9geXKnQY9HFqwYiBxoab2osDRny/sW55fCtjODnyIxUWe3BX
JNq0dnHRQgPsihJs/Uqlaqr4NWtSJWzfTlb+WsxtkdxaY9LdQi2irAfLp9yTf5Q7
wrVnVe2KtffeJwlRoWTcK9ArdCX1JBRdpPgTGiygAxJYPoF7nrhpG1sp+dB3gMJ+
lOmbxkf+7rDJG9PfdjbM/8liFRVd5snrjkQ2nRdUzLvKXKM/VlYVVmn6q/ISQ9F3
V9dl1zYINNxXdXA7Rt71FrKKDmqxn8zluxHWyge+41vFW+k5J6u6t27QvIn/+BtP
5WOnAYHY/KkOS9CtSOXUhqosDfUxs4t+t/9Ul4vZdGF6qrYNleYbZx3cFqfbZfV2
1T2B3QCTuX9HJ5mQ1ymSxby4HO1jplz3ptO9JvpeeUOewCRois8PshA9qyBISdhV
NYcjH49wG+CszVpb0JchC7BbtGoKNXYsm+RsVgYjKnTc3ulP4omR6LEr+kW+8b0A
edRTg6bP3OIeF5QsCFfzmvxaCOPi/lJ1Q0HXPvf8AtYRkagzVLhyC0/v2n2LlOMh
xAxOKPffH73lG4PQEyclQMgu1yFD1I80kw9YX4G9h3oGhneygeuIkQl0AtFiSjBt
BnB/RGuObu2LwU1e0we4hMOaeQk5abVFqJVuuZ/cK/xAthYaOGU8dGrbAxJlDVYm
APP9I79FMYmYoTG06wwAJIrv69DPlUoNFBomfmnBBr6fc0X6xdHwkMoFAafBeOtx
wAU34Uh7uSfE0W5r8crnctEG4aRll38Bg23sSr2xHYN3+Lt9sT+QjIJ/OhqQfkhL
mSekPbuePmaxYkzKXU/bUuHqPChCmNE45EjH6Z1ok/nw86pEZWUQOxFWDcn4vKES
W5QBcmOSAEIMbjunIV4xeSgS9R6L65tD3tDQdNe9I9E27DcMXv4J54pQdvAhTaRL
YNPcZmgksSEH8EQAOOrE1+3t0GwbnewlBy3ziVSjPwZ7iecLDdagofUoCEMOip8W
6GGAfldQurOKjwD8JKuaWrM/0VXGs8VY1crvivZyobxMPfYyRGQq4cQvyrYKqvH0
EaeqBQld3egE/i2ijzJD6UzCCRhtyJTEGFcydPEFTfJzqIP752p4JAKd5sZp7e0H
nlIgpThWoNBvxaWr3wwvCT6n56lLRWzkXDC3F0K3VucKwSFnwap1oY23iO4JjaVt
RAkiyFwL+sFC6LPftGvlDuBSTmyOByKb0+lbxz5H0IK1Kwe2fdZSkah3Q4Ii+BlQ
ZPSB8aMX0dNczEqEU5jYGBd7b7OdaiogL+AxTssUGjmOucS5/Jznq8oWwbXvF8Zg
GP3nbKf604qc/P3xcTyvG0lPG8ZJPkBdYJbCYbxYSYJEZdOaT/rRlXL7FxzmQiz+
TBjDmswONEhfyz7Uofnkn1fyL6v9u7V9syqt4AOgr6Z6UjpzIQ+xF8b5mpWvSUjx
sVc2yufo4i2nH0vqv9L7UVy75PLfyT8jrMLoTG23AscBPsEoJGQqYR99UdC2t/lH
8bsMKf1HkRbWie2+VxOBWn1iECKNfeOj5mvdZGqxOsCYQhOdpGSDg+Pq9uB6u0CX
dxme2Qmq8Nk8+tubomMZwMRfF4xQE+uNMAiyt4fsXBOUAoU/MkMYhJtVi1Cx4o5T
etHayPZU7Y7+0TTU91F1v8q3p2P9e/BXSzIQpR3lzwz4g3BMPyeadgoqxR4+wfEa
dwfcXNHvDFVUON2klJiu3/lMGwRbNwgArQeBn9X+Mn4v5eA9vXYMx3me8KBKVvQi
dnnouPoN+cSwjxfSkLu++B3ci1DFEjPQnSk0pUr/Y42izXYK53zeTNHsL/Vqh6Fh
cHByWPVMkj5fWljClP1IrMVdQv/K76sWLEW/BmH8SkGQDZS3fGEA9WOkn9qRrlIf
P1MuJ2XO9PvA9Xa0Mrizfo5jGoHGiOA72zrG2KuhjCstDXwQcR2yCYBloSkybgCR
jnNfYlc13OoAHUdeW7qtZFJZfV/65S5ARv3GgB93fZDXGIVQWd1WgZTTrDXZ/ngC
UyI3QZTLmchWDQeJypXA5MXVeUV2dcCCPIErjspXgVtCFEcd6q2pjOAm5rmRN3cW
hdZ9aldLfAu9uscNedWpX6HrNxU+n5FXcVjwRR5Lj3teF0rMw1TcmVmCq6xZXgr5
01arwFJXN2bzOcOAnymsIr5RDwgURoU5KnoxDt2V3Irc95DbF+zUYNaZWeYkG1c7
NInGfLxztqOsje3cwjg/jjSBAl++3iS/0bKVDDjwYI0FNeXigCXjjFM1zHG6+YtI
HMz54agBx3MeiCdB2K3/PgkGD3IBRTOPZCUGV/EIgYLbHZX0070qXxhtynNYI6z6
l3DVWLe+0Yn2GjtZi/CMUCEHba/fdQ9Qo1MMZcyjKVQoJU3ao266o8GBuTdOVbLM
TpsL0RZNYArZWV3c/6iX17Pa2uTcx/lwZVUKdHIxBGQOUz4qX4hlp4rCONGVkyuF
SzAlytkwBKshRhk9Y0UEvXBOCFUejsBIzrr4HwVRoPajLxoptHGQZ8/SL14gLJvo
s/AEWxnJkKA1bAhMwQy61Ps3O1Pix/9HxpLTupd/hzWOmx4BQ+BG2vOz3bMItZYE
H+NdllzoocG+6O0XsGIkELb1QgapNI1juL9iC+XYdmIXPi8J6F0E22Yfp69e6wax
R/ROKT+Pu4Z4IKe8VnXteSr+jQMmJupnolYXKo3xmtvlxVZMKwmrpfH6f18jjdHP
YCc2FLhP72jxClITnvwGJ4dFXZ3S52UENAYq60VB5LvoiX2eCy2hgy6aSTgWMqxw
xWI7NMEdCCHE3MMjIRmtPjN9NeDpeVp83SLtLnO+2kMXksKFPnHpd+MUuAMArpNh
AXJUt37vVoNon0U2gLXJWrnNguumeeYj4tvZL909LTjThuAGEPfgA4WI1K65xiMM
MhFwuXG26yqqsJkg6pMhEsN9kyz35jUVh+ihpX/i/rITL0RzP9Km155NVWIGzuQB
rF+hNSMrxEyMYRV1sesru1jrfr4S+FepbxaOXWlH78yScMqwhorWuU6zWnaXUy+M
tPhew6tIlm+RBwJC10kgq2x7atSN8kvnNkGbZIAmiNlQiHEtpS/P7mR3qteTcwvs
7GN7b7+vqiUz+/dD2i9oD0bsfAhB1HLkdoEXWg/yoIGvgbGIqbYlUKNkS8J+SMnl
M5AA/TdHku871bh2vQaBvZtISEf7Xm0Q+KJGjUj9+bdUy2zmY9qZCJXrGzisQXMu
NErryMFMtsJhdVhNXbl5Yfg4K9ufTPNJ4hReXoZHCC6uui+R/14jrPemVI8DAxGk
qacV4orVQw2hHqAcyqt104TaaNBrYmOIkFxXLF1+APz1kBaJMVA8FE73Sw/8qb95
NJ6/ske2W11sFjXV6PQZE2pT92UM9sRCPzdVycws8QvkNAb1b5M1fPwYSu+NaCaN
IltmHHIy88S/zeXZOO3h8OTUNFIzh2TkTUo1OGqEDaxFEpiPHzz5GnHfF+wxWAcq
CXryIZxTo4pSwVAxtCRA4BQYxdPcRwzom+ciSyvWcJ1ObpVo3qiIHNYr71SXgI1C
9MjXro/5LI4Qq3ESssU9owWrAS866sXz6vZGp0ICQB+javYSc7Ux7ynIiN+8jygh
5vyTmwUxJsQP+9nglFVMvgnsfZDuavbFMYNT8+t62BCv2cHEXldxNWQFn4q5JfsW
er+yPqeiUAgCaZZBf4mZo8RUKSsxmtZk94YbdHeMjvoqF3cpjlNDp0sXJNBiffRa
d0k3zShERNAe/GZHvMDOJY5CnD8r7KKd86F+b7elxYflVfvlfprdQP7Y1V9ZEeDu
Bp5u68R89poHt9K49EkjOIc/f8sUG5meep2pWXi0c8cGLdL2rN4j17s8Vti0Jkjr
eCAbrWM/QCYzbFGJakGFqtawLC0HVD+GI9CRcdx3ZtiUz363YdcD1FzFde14v2mn
BWBieegqO9i99CiPgLyWL3IxTU5MvvkxKVuSifUWSVqbuemgTtSB/ZfR1RKHSw+f
8e+4KVPHkUCFTAtRa220T5e7UzuJr1q/B5mGjx4+Pq4TmD1h5XTLs9qz4kLD2UIp
rbRC/MFMQWID7WJqXuAbMxpqyOGMiupWv203NlPuKCyLYhiHe6hpBWc1z2PGNcJ7
lZ/JF+BZ9k/Uh/2uENXBFMY5kfPywIY1O0c0XpojPMADxxVAVbu4IYari7ne+IDP
e1zZatJtPkx9MFKqpOBjqFbFoAeSjcylurc0v291dNzQDUj5AtXohDQ4WR0yHbPD
Fx9PW8V47lCZneY6AuUDRSVMiGeV+Q6AG5OIuxGzyfOQOJ2WKhot9c0cwnZR0GWe
KCzA4N2FSreAsv8CuN+QowkPcvsTpqXdQ4Xo+NqKbCIRDF/ccWpNV73P7sALqnKz
qmDM3VWs2PFK+nxEISQ53LVNDvfenU0Tfg/xqUWUmIj22Wkr0qQ+yVMD73b0w8Cs
el79lg7j/fiM0knr+mKQftnYcrnd+q6zIf8LBS62VSMxib+etOZUsa44HF923Vc4
fx6rY57IuovRZbFaDywPzSgiV9BVRwFOHMzcQgHUH7O9iIQ4gGFvn1JP9/D9SWKu
hNc73xwWGd+aAbVrcXrPH6KiqK6itap3t2GPKSRumwisY99oeEFgIcvpK9eknTI5
ieKw8c+6rY5mwvfTTuJyKmbVoeQ2CpEC9lAmzESfUlcCaGnPFkENDOU5tgNHHDKy
WTRAwX04VHfauJK5wX7M9Z4NMBoWpXaV89hW1s1cwkwaj401Jw8Jy/SMrJlW12DI
ndUfnUC0xuvaney/O8p4BngGCBX+3op+g+UpFXPZ+a88+bDGwdNhqk5IIonzvwqz
LqdhOfSQIC1MAxy/PXEPFlTfTDkHaUj9lSYQyfitj2ZW7R3zMouLauKb0KyLOnUZ
s7nCKIVAt1dJWGcuvKPTWiI4tSjiRAF7YMtsrL3CuiyxkYvmz8Gs8St+VQdnQpHX
CoJ6YTZQjZ5xHurJlTcF8KHqT6ca18YgnTyaOCc/jNtEqv3ROk36yysD5BuAwtB5
e/NjkeuXIafbGl+dxHjcXuGIH9CaCwtpJYl4LPBm3l1YOew6swIWoxltXqEK/Mjn
1L0W/IPUTrrjz/xTWfgVtrabLCnANWbmGQKlVivXa7c1AykQvN6og+mQ07QcJzbt
tKyFAXkSR6pnfrSoEaNmnczs5YSmK93gBG/hDvedLByTgJBuaxcetxzpFN9Yiq/a
9P/jPzyyN+YT7C/sdz4uNVI2xPqmbj17bwRSw8lMt8KCDzR8GAddmzxwK4sV1xRW
YvkJZPBLeud3Vilm39XWwPDhQ5HjTfTVwGZPa8rK8QwRNcwdRR8RFhKlfqVDcav2
XDOeI+hMSoIt+dUEO71Sb0yRr2VuHnAX4NBmPHqWig0H90VDeKEmQqJqmq3POa07
RUz3KysnAUS7UVsOPhLrUN+L/1dOMUZwveLnRwZw07wZyjpPJASjXt+nYeptDN7O
VRXDXOpoejOYbskfOpiujnyeVQWOojB9dtySV6Z0oyNIcXnGTzGcUVQ9ydD0LjnB
3YFoMpHCbgZAfMRKWYdNZj95UMcKI/hhpMeumBSoEnpbL+5IKswzctf8AC9ytR6v
08DhYmoQEBlC7SbgIMk0m8LahTQBJxrcQ8qVW5pJd/7a8Q02Q+nkz4EroTzCRRXC
moIhcGBypVHhijtKcdJdIj2F5tMcHp74dD+VAgXAE9jF0r7QR4hIB5yw4jGKPPbB
+oczrfiqiG4IFkp31AgBBt/SsjQj3J7NSd2r37e1Nm3tWC9qLRISEeVUABTNpts4
S9+WbOmBBUrwPSGvG3rvM0v0ECq06IRwFQWpVtsqR6YCGVQKSk97PTpmXL/tcFLC
q1+xewNAsyEqFGPJM9MBnN2hf3GNEazyr2j4/mb4q4wCOBckyr3GAx691npF5S90
HI89JiwWCuBb4jln89l5MoH2Ib8aYb3NZD+Tu+0b6HN0pdE3aPhFxPYxI9/3oqKS
rCJWaHXHWpxcINKq/YI+ltTDe8fNi8j1uMUOaUVlXECKcMhsxgB1+rAixMXS86ue
I+Z6Ty2/MJMS7EVgY+1h1dLCsyT2n81SLNeXI45AdNMO1P8/BWZwLcrA5H3wqg7d
1VCX1KsUf+2L9HEi7FrHZQTfB185tV7tHYe4BuQYR3e47aF1KnRo60QC6V8pIBXx
R1FkNEbAUd+az03XVB1fyQaJTHnW8i7wLliaXTjopVSVmsBSguJCUwByK5mI232f
W5hqcArw6bY4tPfq80H4MMME5UlmgA9DaBgcstJdhtJalGI4rR/UgtFYNJOcYWjB
RWT2v5sFnYfsSy7KOWSERsWqBr7yeR4rng0p3DwQkkrCH4HD9fLpoKSYd2Vbq4NP
pjL55dpsLGqbnV0cWafMHDzIIns+P74QIfPA6tiUOFGzTDrIYPPXppJxmzrjd7bG
ttxnMvK47ANUKpGuFBX5p0bdCuzfpVXW1EL6G5suQ/Jo10VhdDfbKRdn66pxLbN9
JBlMgutphdn15QyWS7kFAgrKWpARiXNu2Y3hCVwWvY4o41mDaCT07r4UMIW5WtwV
5FwjYDrK8X1JT0+PjXMhQMXYFykzR6DhcwoLw53aiYRIgsN8+K+TcLrs8pOibFfG
5gugZDL9ogpG//I95/06vaZcWBNQ1q1QKYSCvh2YrNFsRD1vBKbMfmCWkiAuFwYu
to2iGK/OrLKiysTbujo2K8XsceqaoNwnppTX0U2cKSj8pDfJrLcv1rAsEWh6g94O
83ZzXuol+NdmIlvcjsd/RUE0EpKLuoiQmO3Wz33ooG9zzdT+gEyRatK7BOafLWsn
LzCJPGxl/KchxCLxUdpUMCsVMiHvbj0cxOpLVHhsZaE5K7h/OUV9OPd91a3TPOhR
7cEkjhan+04s8Ukgi+O3rgfjCUaXI9TiMTy9FwYDNsSzMUTavsTMToNlF3PRsbQm
jnKvjr/co/jEAtFR7XTWbzTFXXh2nukWL/UNkvumm7ZTWpmm/h4BHLEudSKGcWeR
M57Zq34vAWjSKiHiI2C98i+oG4gus305pmgLs9sUOvmMqXj2rmblPNo372gsz5fs
ebxEQYxKYyeNGXUS0EKbO1VWv3LE0uH2/KcITQ6/fSDCICbwelGdGMwdY0klNgBJ
f2mjiiIQYalBfRjOX4P07Fr8aBq5aRLtfJTUfv1gNXpnJUduhxj42M2obXEPxrDo
ZDbzLRRR7PpKVLeGUlLiYmscdmSJyKQBMsKl0VecPVq+0lSU8pZ9rq0esq7nWuyR
/pITPhWpA+7UsWd92/O/gH/jYcP3TKMN/w2GbN4xt6H/dfzyac7yhyDCJRsu5sSe
ikPFSR6tmo6sfllz/EdZ+KDLrr9VUNcSU4MhEW6lX8IPTcW/gVKqbXgillVAutZk
4lPIA5T2EkaXnzhjoseg49IpMdHFTYVzq0sUbbzCHBC9edREBhxW2Bu5TNT6kANG
Db3OHOnTrD+bGkqaRpd0X0K/o+TA/Er3fqFhgVPoFzZiIp7GXKgoQc0GNfQCO//r
B2O56qS1g18GnXQVAaVazZHhB+0Ezcl97KgghikrfUpNGWDb2iz5MceZb6gX98H1
1R+a7RDLlv7Ok+BG1DzLwHg5hsMYkS+ssFPbvPsgBap1YEc3OmGbKSGgPSpEnMKG
tYJhojyDa5pEwjEEVDzkdxAn664bXbGwoASE+DHys+PHHdKOokoaacJiduU25EI/
aeqjdU3iZmMpMzHFGYGcx5W74Snk/UDLYoL6pOCH3CS65rAFXbQsALvEPXAYJ5jH
9AVEcJ1VkuE2vvj8lAaeOIOIQPOLj3QXLZzStuomFlHMe1c6/eX6msacaQm03h90
XrrxLW4EKwNIXKlOPK6oq+rXXBm5MeRXRXKDgagQThgwfL+dPWWHzP7FhybRFPkv
qhcKFjpKSAHXYm1IeRoMu+BuhCF2r0oW9gMzZ8MFwzsKxwgnbP7B1Xvuc3Lgia9u
NrBFAxEYz326X9SkX/Goio0UxVxRxbtGeJ+/YDORNhO4M63m7gr2bc77SPiEwIKe
42+cvQL2AxqCT/IvZOXOfOS20jJjkrNi5GtHmuYBeyzWtG6JE+SoBnPOGR++PZOk
JL1mAj7MIjT1j+ePowpEElr7Xsnu9gx2BymJZVePlbwL/aHFHjPXXre8b0BvGeZf
RVXGwYh6Oa4O2Nww8LvLcPTWUqQFZSfd50x4IQN/v82rfRqeWIJKt4PZyPr1xTKp
cSDQEpItzjeBoR5NT/TW3udQH1MXnWeV+F3uuCUN8DIPYzdcXPxo4LeRefG26jYu
W26f6iBf7SQsuA5rxgCoiSx+cIoNXHS+9/UNJ/H58I23nktHMmgzpLUgdc2XfCIy
/C7FlBzwKls4Qh06xE95mKk/Ag6anwca8PQO7gVhZHB3dbbWb9++AmaX/EFeULPD
QPHY77c0KQLICyZ8FZ6IWGS/Dvq2L5f+TdktxBuJokxfwR7mCd9BqmLuw71hX07A
MMnkTLECeh3UT9bkUpaQniN0n82HGfwfiHrwphCq0zxZr8w72sI3M9MCxER1+IWQ
mId1bpPjcQb+koHFqMH4hXKMNh9DwUlckP433uZOOnwigQZK02T6NHpbyQLGXZhz
FP36CXWmBjRPCAgfqaPLgI6AcrdYOQQbvBAkrqscU+BT2y4CxzJp8dBUAP3uKBGl
uOAv6AAVFEMth+wu6FAjqZjqH/taUpHP8MI+ncsyEoQAytUAyGA7EALQvhvtL6+l
PV1eCJVidYiMrj2trdupkllGEDDjfnLtLFvrWUGKeQcapGPFLl89QIq+XYidoGch
VmK50iRqV6mBNYRCvatsdEQ2DZk6n/5dguRdnILVCotcuDcxj2QblqY+G77db9tB
Ws+IIivYsltMYAoVVdPtZSM0XfXie4FBAkxweuPXAm9KFFfO+0vFmKTPukni+cQ+
5nr3CHXV4HWRhMV4H5Q6VCqn08DLtC29VUIp/lRslrUXTrrwOzLhddnrV5VowK7X
rke4x6x/OJiZZE1IvpWZPqD/cJLw3a9aLouyNMixgzm7QBisjKZclpcRxnbOZbd/
5f35V9H/KyCrXQxw5Cm0QEWkCyYtJ1vA6ofdh0vJFcaIuLdswbsJw+Gvmf8UB1j1
HXL3+ZkAyz5K0lCrksifmiIGpRRqRG9YpzieGNMj7V33tOZoj5+m/cIkGESUh537
pt7KRUNCGO/QS6817ev8pBLERiXcJjT0vBb2IYNgw9g4flNAdjcFWCF+Xc5BaQpI
QiH7O3c8tqJKy0YIvLMCoUcKFxixueW+tcpZNWf5H+KUebtSTuufSrMPX5q4uklg
PFeG8SUWWUv0AIKoo/0uhLNmhtqvepJL54NZms/K9S0Vf3J0ic3LQPDvvE5nRf++
aGoMkv+2FGvMTbO02HbQShfYF1se+AGrzBMWlHlY4Cen0tb3xRi4LHV7shEVHML/
6tTSufRV9jom9ZudP1N30q53gH0b+hnxUZxzFWoJZKe7bi3bM4vuPkwn9/WIJikr
kr5sXA2LqU75aWazf7/SFwGg8YmNZoxAcXG+Di2+ep3JrfnpjhKCxm+fOxF3LBxE
uXoEdXcTrEORuUf8rK3Pqkkmbq/kBRF4FmwCHUJdZtmJVBh7aLeHwv9hpQF0JV1v
Nx4cE3srDkttmVyUaCOfWYAR1Q1L3+V1reRY3QB7cMm3h3RakrZYfqVfOEN0JRg2
xBIvxabr4Owc3ia/lXN5t7ZAkQA2WL3Runl2AbF3/iFRq+FmeIJyJfe2gxkhRyXo
sVQ6ajUulv2OLKTSICJDmH0t64emJP/Xb3LXJHIFTw990WX1VOxAJ/CmoUPdeyYy
iC1wi/Z9qyxNiVvM1lk1yiUlSY196ULkR2eyg0ePiM50HcP6WD1vkuTrXeeV7uW2
4nRedD2+IPWRHwIiilVezJfVw4sqjqTCHw8dc4tBMs2bcKh6XF/SvL+UvP+FOyBb
PUmxFmXmxQcUxWM6sNqa6pHsnREPiRmQr7lMfH+KU5iMnBKGKWIKb1pq4UjSgRGR
s5FHTYZNCEmTE+AVz5ZxKD4ceiitOnzF0zMnnMNqqj0RQjvKQFZEkVlzHFfSnDyR
B5LMyeDNvRJdl8scwEFoiPfaycn4OFSm2F6YPYJi6s2vfvt0aI76//gVkwAXEhpC
kBPeJtwxyKlFhivpX3As8oYtAL0+HfrC3t85YakTzUcK0qVzvxJ1MWT8NxDck6eZ
UzeoeAsOCLuJWuSiD8xS8m9mD7Z7SDas9SdJMi5tn3SUyPdAn+sUTPrRxO4JX2x7
KjbhRgBvryx8QdfJj5GRxiDy7ITEYlGCNGJoOkxVBwbthVS59ZSrjOPy3maeWF0w
5P/uqkjo9WlSVUMkyl/j1vYcWONnoKuUZ8yBDOdz/u89xAqjtmTayXIglO8yYbbL
v+jyoe1XuftvpzuseX9AqjOZOcutdBdKu5vWMD2VqCf7jTc2UzVWP3xzZf93QRvR
8BLq9RY38zVP5NHfRrbDdVhJ1qh8dd5EUwjBBy7l0DiNWoe0lVgDfPXTvBNxpB5T
1NZgycKpEHNOZrdc0ouVdT2NH/PIAHEEoVBMLUv9LDbPNIem1hjiyO2H7Yaltus/
dM+5pIoZM2cE8q28ygspQndbPc094VobNaqV9QSFMgBcvmNe65nHPGA1+rfl16Bw
IUpF1Z/5bJBF+KBGsI6HEOTEDUiGQ/08cQzMCP8h4WVtLd988XCYgElOF3WKw6+g
Nxf+VUex3WMJwFwyZ+qz98i7ndYi/IH6S2q3zVYf7VfAJB3IfvEYTj1MlbtWU0bv
NdJgwTSYbDoLwM7JSLwM3eIcp7NTd1dKFFaYhq5m3lbQIUSZAQ+/s8YwOhzSs3Rn
nDxVaxCumQInKbl9n9iVLLGntSW9+wNiR8QYNevkxKJqqEaD0zQsxYYhlrogNd3F
mkSSeWyPZPjt32byOE9adHIUDngDl9OG/5AV8VjqTx2OaQHCj3s174NAskr0+lTb
40FZS4hPUa4ZlQJh181mtfyNeF1vxUqaq0JiknqS785ImvsMDm/I+328Q91eu7Qs
OqJHN6NVRDZYKOCUOquG10CDoQUJ4HNlR14pjEOHrWR9J+QmOyXxwcCOr/ecl8P0
+2NGYrg4e5jQGHClegDbV01ujfKLK4uOM/cnZBaSoeNpE0arSxQ1gEL4JaSEEsfR
S5W7taKhh7ds9q0DGYpTqcZ+ZfU9pzy7FuE/1eBiud1JpX9BdRQuoJTduuPA4Hyq
sdRwt3/9bdb4nPqGPNfRbeLNHdsH0TFr+uq2Fr31gSjujl4EMtMOe/Gjl+W6PfXR
m2Aa/jkZnHKj1mUFGnn0oVXqLYaMB+XbgKnxpRYzlQ3aw4hB82oEoP0aopLToghO
i/YivAKrX3HGlcFwTiMSDXgok8zX8w/++DbpLkGJN9gS5qfAu+n0goWt0tFJVP8n
ax+PMfp/5VmLzVzPlDbwalWMw3GheHiAwiCIj9wa+AqhyOqeWXUAklPtXRLjHjH2
aK+xRd5g/yyz5TiasXkPZUAMxgiVU+mNFSoCCjMw09jynLvaXea9M2Xfpdtd9Lav
D8viX2f1Y0CrnNURAVuYisQ8+ZQZJkUgSPUv+gYpPHP19lQnPQ7L3qgAUpQoezT7
J7vxUOkbRjXlUiTbehoCr3qfqfD200IkZ1dDRExpXjPhJtd8c/AyDqR23lPYN5K+
cvMpSsafSsaxP57M/Mfw3SbytGPuvy9iwNXCKQoAVPg35yrl0OTTpiklMtWDXeJF
YqNB3KmZO2FnMKIlJY7TEGUlkDJcrMdENNhkYIDHBIxx8ZqVQsQYqW8pnawsbOjY
Y6QEvgZULU6VHORbYqNzNvOQ6UCW3XcOmpKoLcjPrelUlNAKPX5anjM8sN53CSLN
sHHk98/gdAWpPR95d7k/rwJiLcqGsV68WkxVy35jxVHlbsd3bL9NqT2mIsGV95U4
QbJputj3OzSBhYzCWvkNrlNP/RTDRVDlFrDSm1v1HF8/QDBs8u0KHx/5BY/M+z/S
x2q6J2LewL2eLKjhJcqs9b9r/qhrw4H7wKawX7csF/6x5NIfhkpaV5slCK6bMp4j
L1/iEBf3f1/ufydy8uLVlYrcwM/SOQ3+o68vqWPVzrShcA+oBJj8ij/7rUHAxiGd
RW90wByHaui6t9L4NIBklxMPwRlunyGIVuh/dT6xefAQlYzWk4jTn258DUva+Nqz
xrBkjmObL0OBezMddjFYaDJaa2NMig83pfFoLEzX0+ABy5o8yHEdUthX17OOTimW
WLoMQMUpVvc4xl0efB+i9eBF5RovfLiItvWCQwUSu0Tu0GLLNC2BGLcbPtyCBuQb
cM1sEwUFM7u3IKvprOjNV+RYy4WrLjejeTMQoNe4fvad8FbyKWMdLQtdfoVBU1jp
hqN+0OTpG5Q9WRGeO4H1VIj1v8LA3ULXKriTFksvZ+4LTbO1imCMYiAGT+p5Ez/U
UeJfmqyRABT3GJpMis2qIl/Tw3TT0IfhyT6JQNvp+DqZClmDPncYknlmxZFgmFgv
1Dnu0L1RloyVvjz5mCsAQFCo+udLEGZ/z/jhcs883ZxJf9m1uC/scFWHPv1qMx75
qGNy+o3gHux2oonnmDC0mXv7vNJ473onN6t7o0+yWatsa838HGAJ9a0xMfuzArJB
v3JL3ZSwMV30XAKGQUqQzvTARQayFHXO9L1wVDiIZgxZ53iEn28FFZZN1erUPo8d
MbqLzS+i/MhKwB9HZgN6P9K2ciowt64uWqeY8ET9WO3Imh3BD2v3rU7kVFHy42Ju
4zjgtAstL+21B+JxNxBvFGA3lfRDuTNwIduOsRnVG/dgw9YpNCiBPsIgCl/Eo2/g
apHD2L1qmr8k6ziN0rBGrzQdKop191kr1Jx8kAf0kLHgCW9Zq3omUSCe+h9aSMtI
ACwT7b2laJtalFROot9DV6Gvzz92Zb0q7a1P1HJmnNvZOErEcC4JG/O9qsR8tsqJ
8qiqMZnkXuptjY5lgejqaTMvY+yUlipCf4C9WrbXNt1bF9FYZiZwLZ98NUsSgDde
baaEC3v4YWY5Amd6o8aDQ5OBg4rz/fJa510ikFEH/vtj6ggxhb7vPcgWm3e2LLkT
48EahTXF6mcg/SoxgkMQT1A0EnJKfYHoIeVRKoNNpyhO4b8X7fK1WHP1fLCr07jb
I3FHCG4i0pRWwWDs6sZjDl8zCFFer4YilbFcGxM6cHxoiFngF1K97Z08zMuAO4tn
FocME6B3/x3l6EFZwZdHXbb9pKbz+nxVbhwnkD7zU+fJpaJsfw930fJu+joRQWCE
sqAYtLF2EYzwHOa3fIfMnobQ2P3hF+yX1Xk2p9SHEYYbFr/dzUhFgr2JHfJuKMMN
fzYZHULYZIkLqMxd5g1PELtpctLvDFb139XmMaOOjqM73jU5b99o7Y2rG/VsNWB0
cSK0Vbr0/NL8EF6aL1jakwo3Bd1rjgri0LXLktmBRxsXfI4/jZQF64VqSUcgw/u/
op3OPyboqeREnkrFECqcN/dnMuyfs9UZcHmH6pY5/W1vbak5BlE9FSgysFmMNSC2
N2hQg5NFywGb5WZ9E98sCRs4sswgUUlq/DpWK3Ndyi6IPNUuzkP2/+Y5gznevhgM
z//N521b0NDdPulz6Y32zjih6PYO+9w2nJ4cmIx/S7Shxb4BNGitu+vYWDRxOy9l
TBl0xxRJnKJ+PUux5+pD5QwvRxGH5gRAuvSDoXpCfQsPmvv8qu2JXyHCJvqChXlp
mFoOq733Zwq8YdgVgp9HhWYGAML6Hkmzt7Q2cymTGHqO+59zXEL5KmFcXBklkbaW
YQl2FIWeyXBJ0RQCc3LWqnJIhm6G12cwqiXDbnUOALIvtsxrXjrjuPYLkN5OmqaV
e1CILN93QgizLAIStYEjXuvjIku7Ga4hd21RLMq3xqv0b/jepA38OoSX7/FhwuLk
XP7x4YUkT/lx6fP6KJV6Kat3laQZGaZ9fu7Q501OAb+EjuI88pgMWZRv6z22sdfP
0HoQ6engkkg99d9JTteNCfVd1Y80SfRsvRMGMJC7qlgxSRMI8zDfq8bWuukFQngK
oT1OzO0RI8FUlXgsRnnKBx6UsycEcIsn2sFxI3/xgPSFs7XBFYFrY0a+qJdV3vA6
OA9i8urLgb1rLmJfy+LA4xpMSWSb98jbJxNjHi70C/k0mBfUYWMitb3GEwLzM7Tg
v1kpCXgf7nf/z3XA/oICOmItWU2liDR6niED9N908JDkcUBpXcZZQ9BgSbuEb12q
8y9QLkTqEE8g/KfjwCaOxtWlQvBdTfQyRlCn8ISmpiaD2OPpHUtSIQTFXat3ezAO
28TfvhW4xqVULdp93L1dVa3i8CfGjEA8HD4QgActEtCzWYPcay/4nj3PnQS/19Rq
C8xcJmSRxwrA1fhRFJ3Yff4poKioTtDLuMpLMbitT9Tai5TMH0yX1IEjTjwQhvTd
s7aPK/kzLyklTcYzu0RZ/uMX9otTBKrTtcGz0gTfwpX63BgdQ9wj9E4O0Tg0Kydu
ozL/jbNEkaLMw/3nX3XJDOj1r47j11l+rYDJxIjuhIEMe2Wq3foCWagRnKyKRs2R
93ZKwxF0UYUrA05y0ihoT+m12Q/CVr5EbfXnWhUhySmftPl87s3KCLv57/rnCBmL
kX0t2ggYbjx/y4KlkCjGFSlopn5QWBgh3tq4VMnsXfaysv/mZq03C7QSB/QqMVo+
NwS/O8ZLcJ70zCI+xr2KB3SqVWZHc0ly4wH5RX6TtDlyntWRsGRIu+bdln+XrLzr
gfLXsiltYCBKAW1CeT+iV+Tv9DRx+S/7j04A1n+9zRKlfgD3Xwpd/lW0PBcLTd4S
U35bnilaZgTIc+VJENmYlm0gG/1sa3bD0HvgqLZzj+EvPyXLZXOakQBlSeyNXWxj
IPg9FmboPq7WvXeXNeZVw1bnnGCPuGZvBld1dkMTNY0nzSJCBXa1alOuQkMTEVGz
SA+doIpaDHMo43Krp5M4I1XA3cbjuIZXE0JWu5aaQgVyZ4RrbuSBE+aNtdJD2VcR
mR9UNORaUkIrh/87181uIuc82A5mi7iv4vW62xUKC4i2uU1D/raSStrLyN8U+4ek
1vug+GUN1cGH7G1ZmTwPYczCxEhtSkvCZPUcjmIRr9IDX/RSkdCdZ0pAz4IlpNYI
m7qSEv4FB918aZKme/lw+w12NaXxBeYLgJer7m6+Czn58MVhVytwugY2NSG0dUXu
nLtjb+YMzCbLSnDeNr1V9msXwTc2id7CIa7Raf2qzuXCN6bC/w7brXnS+GbuPBUA
s99mhxtVrqgZOLQA4YKNSiy+h+54TBrH92HeKi3f/iwlT2RjJ66iY8lkh1VEKEgN
7+/rhYUKG1jkn12YpmVrKCDsQ1hf/Se7NzGshsJYvoO2cgGLBTn2IEybKQjk8XBB
Pc8KlQ6rlVrIB6dF/SOdxYXXL6A3mosS9TcUmr6fHzBu89w9rznHOIb1oC+eYO/i
YP4dKpHgmnAdIDdl+SUlCEJ2wDkNS8v1lJd6Yv/S2uCctP6DcZ++DqPlGu4iT/Lh
YpWzPWzQZNbU0rmON7n/Ts/Lo4W/kTWBOCykfaSr5UYnLweX0mHF4XfMq+p1F/AJ
78AFjQ2m49ZKJB/qTxofjTFMS0AZ8HmZ2qbIGibI9r4rXauyfwzTwyDqfGYISyJ2
pQqX+Z+er+igTUeP/2XuAXcI9sDEd6GpRbUlLqo450ECIHGJy8p46KL+f25QXrty
2o0cAsYa20OFUAxE4d6rgDO0K/f9uFysy8HIUoh3OTZNqdkBj8sP9XI2ukipkfsJ
jhN4o/d0zcAo9ITWwDcSMoQq+9/FLiLCD3MqMn3SuXU3ftGFRxZXkZRxrwqrNoov
XCQ45S/PQzlVt0u7P+3mPTz/Hq9nMwJHCVdhUkAadQfS/7AZc9IdS9fFrqUcTO9+
9El+VjwDP4MkHP1oMa7EAh0GX1JJBnEzpkA7+9iQ/38XKSc9sxB4xIl7Lup4KT7m
W/jUgG7BDVGxAqE1PzX6IKWRsusvxMqvGH8I2ed8q75ElK7dHC0TMxHvrVyBOI7f
StIPMLsTfBQ6VZGMMFIFYzHpiL1eZL9OdcVzBScO/KQtSaVlybcjB1/0b71ASqKv
cVWIW19P0tPVThmaFh8fjInu2S1XQcN074NLNapl1K7KnjLZm8/Zfpy9z8pifvQe
cmQKbul1/uqAvaQ5wnq7FjH4Y6zioMyP6YS9M+8J81b7wnPrWH4vCrR3mtsgj70Q
fI8Jl/+hYsg9wv7Gb53aJWYWLf7EOIOY0WpC2ylym6gK5nATyyCAHbxK7dDle0uR
IULQEzVDX1fHaQW5V6dMcuSF9bL1Lx3IwIxVBqWiReOoG33eSLsUStqZdna3Wjtg
jCpULZAdTcQ9N6j3qyrIdaBXjPtNFO9RX/OWoKxK5FchlpJU741ewWQ+ubZtgEFG
UmxaO47XwkoDsiwVA9yq6wHQyEQ1LCXX4iF7e7GKIDcVLsm4WOccs15gBkPV/AKC
BKff9k8n5KfXgGZChbul56VggT47gRGfIK3XYACwf0tnBzMgg6gSy74ka9BL//HZ
+Aq/nLCpqztLUwBVi0qZtJo093pMiNKjvng7F+p0rqcYs0/uUOF/tjfI8iausKab
P7JVBYjMJ2qnd5FrtZs0p1lfdCslGi15LoJYsP5JPRTKPkxclCOfpyfUezW1/ICh
yD/OVjCeSoHjrbQDh6dMkLTDeNRAVjl9qJdqb0ooNUjBtcacXpj7gN586hmWjEdR
p3Vm0XrMpNAHyNaKf725llefg/SmZtZ5ShUC6GCjtlX4vzYb3PnaaRktAuu/IL9V
K2CmgqzBDGnQHZIaZ7q7Dho9jaJNXmpCoPcdsD1iO7vV6XC/GHQ+bZuOM6Nb7Mvr
GM/ULLd8CWyHc452kRZ5ktmQPoZLu0Rd1wEQHp98ZVQMiG6+jfZDl0BPs0vCONmP
08oHzrRYZ+AAg4QwCDe6FgXrI6cIT7BaykItxzj7BG1xbuDoWxSklC0UyW8JwCcz
KKGdq9gB3E994fsDeYsQfCWMk0dK2gJlx5Ib5QTiu0kD77EnmKHIHsoYF+gXNmnf
JcMlN1Baqo+wdydfgum1DSEZ0Ss2qVxfZ0yAJBLTJrDekH+/+wS+NOPBhBN3BiE8
RgCyAUUbiVFVP8H3VJRJ+j2W06HfjXcB2ax1LSUx9GQvJo3vPC71xpbYrZZ1r9As
EeKRh2arDHX020XZhaT/MQ7AHiJv8CLsqnIVOLkAC/YaSQBzqYDOrBCFLN+EvyOp
gAuxV1EFYnbis8qUdEYODoBRz9NAKIZdrww3j9WMKagaLB7v9Ud0zaUWyXMA3TPb
lXjwmxi06ZqeFLwDWWgBJMQxYHYqLEs9CUXeGBpcrpl7PoJD4DyXHny1lBVRqfEv
EYYjbNZ21RTcLHR06M+V+rzgKBVnUhOpfWCKmJZCqRQ9JZPCrFUjN4UN20au7Sqj
R9fxmIwedaNUOmPCJBdsLPa6AWE6FenFoj9XOiYiiSW2uhm1NkimSJdC9D9vu1oN
8ohbzZscWYAo6bj/xhJ3A1mjpKowogNZiI7Jv4SSiXaneVirqNektJ2o7ias7VS9
AqLxw6OKPvC4ktvyAdQYWPmtRrgvy21Pfly8bUMYjf3hwqHUCzymBotlNpHOtz01
FB3vlOwTnEtcRxUAZivN71Y4Cgq+MQOivcboFJ5tUzRLBSru75KvVb7lKKkw4vjW
hTf9pZF97ZH39loef8/oX6Uy/j+lDQQ4TF64nyjbUP35DgQxiEuRlMk5CPvCyNHl
yy16hu3URtMgGLsFbGWRLcK4dna6nXg+dM2Z/za37GZ1zboPBPFx4EMLAeKlFlfx
eR+3CadU2bVta5OKejkVc8Ou3m2F38yCHCURFuny2jUkeP8eVpuI0XdjAy8zQJJo
UeCbjGGRUBnUoNWb4jbThGgcMOZoD4eeUmAEuuLRO6omtbP+Y7uZROGEPS/wBPpD
hqcovUZdWI6p5MBjpiiminc0mHJMvpJ6WPxsTMqLPbvWyjiqGKqHc/zGSYVoRbdu
5luTIRIbGcZFUt9pJSeRn/IoSdyEd54jmjZhCKV9VX/7bLt2xrA6PQOGO5Cg1N96
ZUiJmttTjVwlWbDNtTTG0TwbCBQr3PI/e2FVXm5QdOpk71RU8cUfVq8k4ReNytd1
vL4JI+VHvgB6HeFLAO6JwCqDHTqiP+m3AqrCzWYf8uUxRGXddSo12q3HV/dFlhtP
Dy6aC+Q+mXJzCHyT+1ISSW8XjHr/aBbhdyvWWr4limvpP2KD2CNtyGVbyDlSwKSQ
Ad6x+ox2er2KvmaCxpti4hU6jaqNTTyqcOgIkd18DEh8njGyvNSJvq6pO+BIBvlf
pi3eajRTIZJ1APWk1MDkw6ZDDvantLbeIrqtYDyK/c91C4X48mpY86k0EAQWuz8l
zXLx7wqhwZyu8Z7H/05xXWsfSZEW8nbRnrgUMex8i1v0P1gUwfRW8D8btEDapNyY
YosnuV+S5Kd+4h//Htzr9mv0QTmY8/dCmxEXstKCHmNc+eqJPHff/yQdL0azojdb
V/ulTwNvD9uVs6UfEJpyFHef9lFEzrGcrRnRRvBlY3iIaACHG8wq0XQJoH4neZvQ
5t2Tq4KfS77rjNYS31I1iurt9t+69ClIvOh8/iP38n3OSKxc1wr3QwPQi+mxo1Bs
dkq6g2FLpOojnoLVn7d0yhbZ6e0eXhBVqKZ5cj3T/pBMah26xAt1EepYfC4HKnbP
h2OndFscV8MKicU8RTzfd/ks2U6gWag234KWCKn0IXz6KmQeMp+R6duqqLXed/KN
oTK5KV+WigXUW/AlA4+0vcyuB6sKOAcCQ5ca2SW7P/BWyQ5TwCVO1VSvCPYFM8Fy
OJ7mwdiHFcCwzVKK6G/uZqH/OuVteHAf94VhGj+3oEFWlfoea7S88+wMPRGRSe43
jV+pEFxhQ1nFlcCvc5FIIboG7RvpwtCUUbyO2Y71WeTb5OdQ2i6Fn8SIkHpoLd7F
MEfZm+Fu2tBGgRYO67/65rOkBdtrMf9citeMG7dXhpGG34qwHDHD0huWtwYLOblR
IHzzRiP1oGG03acbtgISJiS5I3zbx83TTrbUXWQZPIeb727jom3KZ59Vy6JF8F24
I4OMhHRUZCDYC1dz+Vy8a+TucNCVi922ABT433IQhfCqSHMxX9S85fH4Ti+utKjq
Cmiq3elHZmDn4GJTho+dgJAa/Jb7uizcaeDbgf+wDNKZSPc6oUZBuMb+yLTd8bJr
Fw8vXgN92WaQY91uF4L+sCwssTFgU3Puj04N4b4RQhdaj/4L386kNjhllqtRGHfZ
PiNR6vbK9sGalLRXiH8tE/gJaB95E0xACJ3wcinMeJwICA9rbZW9xenGFCO61tdB
DWGR50+fEf9Hpuwte5PX0za+nwgcEhvbu9r0zGwCkeemgiQUqaHLl+FhEhLDrxX2
7m3tkEStaHuBhbgHbjMc1bY46EaW4lEbchelk5LHMfh9nTYvkUPvjJnLgm0dCnsq
KlnB2+iBD14MaDy67f5HNIlAn4flLW+lr4X9hemYpsn3oyFfIk9nPPF3tPyTJXER
Tjp/T61+mcqztzwux8Ogewzg1V6XkAd89LzxDZ3WGDGR8sTr+RhKr4+PmExqpOrN
BoUvXnizuzlDo0Etu5DsQ8n1Pyjwn3ZqN8V0RF7YZR9oHjScDMfF7SIZuHdeR0pN
KpRfmLHlM3RJ5N0e4XXNY4j6pQGsz9TsgoqXPPJEE8uhPCl7Z0nzsMYu3I2zAVUU
ysEZ5tV6TgwOgpVTQLDlM1sQ7Mc2W05d8vCjUE9AiNvlsikG0jLESanDuMyDA4Vb
wUQIL6M30IkwcsyRgT3Dp6+NlLDjK2ckOlzW/9YvQGWyhOfwalhJu5Ja5nt8roCU
+uFiljXwo78xMX2+1Akr8PZHdDr8g2HIa9eGPewL0u28xJr546HecJyDqML31YjN
w6R/TikBYkpgy8KKayZwqi3ilAHSdK5OaEQynBYVhDoQLgsLc1NdCTf73Rt/lkix
4hFYmWjsKfz5V/0dmg5oXVdiCpMYCAPqyYiGbanNo5A7MD7tUxzGSD+6cqP+H7/e
IyGsiihRzLXSuNCZv5IzOPs6jrEWAjesXcUYvYF6aezDrQVXD1ohYGP/6JkNsVWm
X3Xn6iT92cDjImuS2fJjOJ6EozwnSG0Q4sXG1P3fgNhZE/Q/3aLxXv+NYhKX2o51
bLuIPJF0aiAkMPW6I5R6JYcDglIju8IAobCawwWRLYq9xasIlfMAUoftCvLzM9oR
lYN6LaaBu3K2VhOK9bDST3GmqdPBHkUh/vL2uV0tNId3qOduloOR9D8S59c4htJw
84ktTnADtNI9yC+qyUe0AiD7DHma19Q4Vqwm20uyNoRqgZ55PLa+N/6zzSYFt3Tt
gOwLGl0ut4fKbiIxKg3S5GDQj8IWd/k3x/MYYAx2XI9pGJaohDREc2K/h35c/I2n
WEeF752TC7cQb4iS/7RoqnP7PrHmI5gzDS4DzjdHLdXZM9Jsh26Vslj8s0AI16UT
D27DT/kti1rH8UgkCEbNHgGp06mvVsWy9gvd5uQ9IHX2R4TqjmqPV+WNZUI3plK3
EOg4LwW3Afw4sLbB9crYbAb5DErNHkDGPtbSw5/Bm59LSvDZEAVDiJMeOnSsB0Vj
KjdPUgdUqy0oGMwReBbWuKtOFCvB1+kxBb9OO8f4uYcFTUZ6xAKkqCsNInlOcdib
AsV9rpQyCzQ1tyk/+QsylD4K39iZc6jej5UYWPsfqgWAst3aaTdyYD3xMDe2CaoS
5Inc8KqJanXMCvacwHf1lOXbtu9TFAkHxZugfQWg4U1t1C8HQimiWr7Mh27apX3G
NcJicI9nMIywu/HkCHJxfNsvr39dVsJy6OHs3PFgHQxltApYp73XoFCUA3VDTzoX
ifiaVjx51DE+f4Wj86EgmLFnjSlxvjybH82GsjifNja3VU0XvUjeoLBr6fJcu6pO
p+HP6W3gRGRhMaIiie86StuQLm3ynXQvwBlToKWqctMx7e1cOIHcabCZhuU/kqka
a0DFY+PnMWT+zpxjln5KAjgQjAbydUmOK8bp6H7Gl4hChnxYk/LVRG/YEfNP+Vp/
SvZ3CCNuNAFqyPoX47Nl/k716wZ/HbbLvJm2Hlt1ct8BsPi31wqvkRA3zNPb8U3t
5DYrACRP1uF+f58tZR5a3dBZhPUMCLbCkUepJ7vHigv1NQE6V75kCILMb1AvS+0c
zpBIhp7dMP9JQ7lDKewzRNUH+EOqGTcdGiG24Ia0vA39HPMrcEAVWMft/JKHbUEK
oUgaOEwVOx3Yo+ovieX6q9jisoOBJ/lTk5707LnyXN1U3M4H/lAtYNWI8Ymx/luf
jIhGl6exEoaGAdojOJBHgNA+IoWBxf4/pAFpdrcvuFjskT9QoCYeV3kvrAY8uVkG
JL3fivWrw1hXACp+4Iq3AxLr1x3HMeIY6B33gJTeVVxk3iYQ5mqfcmyWQDYDmOWq
oFy4unow7DwV/OlDRFnXbKxZsHgEK+VfDbrvx8QmsncmMTlTq1R4uKLBZHt4R0TR
Nu3sXiLotRmAjbUYvZEJq3wXE6TtA2f4rN+aiFQsVkcMZ2AU6+iP3QYOHCqL3xSm
Xitm5d6hQiwix12tA2avA+U9RMIyzfRwcUaM2hhASAwyH4RYb+fMvbYp/x6kbDHL
LOpR4by1KyrdPW42nTyWLc6edQSxuROWV20KbS3EiV7HKNKOFKRi94f6VcYsNabg
2m+rbTZKjRpFbDZySRovleHJyjBC0sATe/ry3Ig3eKtjZDh8T8mZ2Ve712tm7jSB
nAJfmQA0fhYvddIHvKV4CgTLgFOCkKQ0sGFyxFTLmZ9K8c0KZmsjs3kiIgMAHcyW
3LVCAOQDC8FuN7MhMQBPTSg3vrHzIs8gB2WY9KYO1pt4MuLsJfqQQs+01h+Usbyx
4IR6OtmUecNn0f1Pxrhwhm9qQqkx6lK7glboKDbEC9Z0SKZWGabz1B9kJZHTZ68Z
+atgrExCmq9lPH9GZVwL5c9B+znUEDoZuIY2wfTGXARhajD5KNgyUpLScEnvmDVj
7l5B5RIDg7OXtqs/nSwuQBbaLDszcjIJ2WEEzWuGwlEX08tbzgn4cR8+KSLHkZRQ
Tx0VPkheZ3tq3TBPEE8fLBIT2lEcpMRb1MU+zr9x2cBW0uPBhfSlddAxCtbKV8F2
qkyvK0ZsXtZWFGS3NXCvVzFUAsyGuNQg5G/VTi09eyGmQTDIAa3BiCginUq7QAqC
Z3eb78mgb3b7bLf7gGBWn8dNNUuMZmOeJKeEV50/KaPUSWt2zHPatPe39aZlwNPq
zipxFNy1aYsyI5NFy6jbyEKGL9r1xD7nidEAJ/9jAuUHx+WLf2lEUzy/6U72o51l
Fd/bHSOg/gbTSCEZVD+ft+zvbTt7nMBbc91dYBrL9hZKdu2SwuEzsNQRdU67uZOv
J6+sQouBoHbHZCgaAySYUMLkCLNTdUPRDoyCKtYBuUHPFGUgWu7sRWepw4OrtZQ8
k0nkuO4O8gS/azDHsYlA2/rd6kt08qAfWagLeihvYf5oRGNc5e5P7C8gUm2NCq22
2VukR9/E2uW4Vc0LVVZyGeCFDnJLBSDSO+n+Fu6Cxf5UD+mrh/tFfTZFOU7+crFK
TkIF1eouR/vB0BMoTm+/+aFMQOvGBxyxx8f56hYBJNo4DO9icDZPjmC+KcVNMxDs
dDeOzVs2agMJ0/4vhWk2I5xTfZv3gjFGFehTq6TNiyhhEAuBiNaTzVvRYuFEyc5j
YK3//rTMKSs+WVl4K4ouQfoZoN2YZ7PYm7fZK0jhgr4HcRWjBekrmTXp2jUdVXNe
yqNvnVM8X2Ah57PgUo+jVkhMkk6KNWBO5yr+GELcKMgAMUuFr80YXsvQT2H4Z6vH
mYToHuQhq4RImql7XzwZ0zuAFhOLwXNlp1Ua52yzilQgYUP4lW/ccRBB6utLJntf
eicYmgIQifbQ+px4v9D/tYRK5oo6s8qMfpGJ7XIupdyXV5JyIqzq2Oc4orglyD8t
RvRqpDdYoDFsiq8FmYitk7Mkjhs/eww4cfRPGkkSz2rS5hW/N4ycT/jMPkWS0SD0
UgCYslsGR5lKWr0Mz/eke4ONIGOk2FeCi59szURYK8CelaqdymvMcLU4RcArHQSm
7g1BvnV/2JEHSSlry/MG2oJpyxta5cw+fkE5BmiDafMfusK1EuXLZXOlN7jV+u6/
q08VKlb2nLHmCDlzNA8tvCrGEghaBZfoUrhGBSjDVGHi2koLK+RMNYktPICpr6X5
XsRd/rMYzvmFmsWEkn5GIkPuPxgDqPuqIgzE+dW9oQerTQHz5ltALunhDJKLEbTS
jwmCWdrkWEpbr6RxbMglwOvLaiMrJFpaDfn+JX3Iv+h0lTqauQpQHHEKJ3v1H5p7
SoX8m7+phQAHEqq+GqmvkZBomtpz9fDb7I0FpINb7PRYT+qEyzHI/tG/rjW+bfpV
ORdvmyhltUzw8lwxG4LYnbdg2bBEd6HEdJhQmJbWamXZupPajvA4BXkFZ9YNNoVU
+5Jrfa4Pjq+2ji3bdLEYeDCwnULfA6CMK2LwvENjG+dASFm69DUaexr350uw3Vyu
HIGP+FZYj6sPushAKxlPT4auG4o/aCD6HIhE0ZxDdhNxjpG+19pdV4FKLnSspv7y
Q+AipUMySqdno6AWZc4NzxhCdf1WdU3qkHKjwPgXZBmZ4oPPqOxgyE4HxTL/3MSC
/gubiCnA5mnkRtGTVUvs/xUv2K7JafQcI9BRrGTTid+gc+UjhqCiK4i4AfKIYNgz
Ux5zl1Enk0ej2b7ZKOEj4rPkCkqAxRcZM9YoO7Z3V7R9Hid1efYv+VsDyMfXW6CY
byMLPhXDkt041tk5VFEz0PI+I+rA1IgrpvG2rE9bVvIpKeqKOVL6EeX7UC5OAqAr
m1qhyh4o3tJFSyaKMizXizEhrc/iSQZh5S2MYhJ6AFJ8nk9N+em8qu49/aIxLFFa
GA6zjNCnr6X124UFxOLYQNS85PXvSzZ5RahUowsw0sGdlE9vQW0tEaJHSifnhc9K
ySO4RBAKK417sB3qH6uh591JoINFHJ2g8dbZMq5TMQnuxOtFpxszPqMQGxim+uTT
uU2JD6PKu4vkj/9SUfZj/FCB6lHYu6VBh2CsQf3j7KTfepcUvOd7nWelGM4SrlrB
oIY3O0PJyj7VwIFo2wxslSj6SHa8HJpHSURCU4cq+TIH7Nfch/2GzH+GyamwVBq+
satBZJ1ezT3YFu8LtzaDtDhsdTrmnCpKZvWDttcs4QRseGpVKimHQpqz+4DFxx5I
tDk616y5A5m0rJO/2r1Lkq2xBsRX3nSsx3vPrw4gROZ7B/6nACUBydkCtjxb2ggv
bD0qLiY6pouLiFmVBAI/nFQjIdYmuouqeo5b0gNravsF0M0Q3NyCvmn6gBBtoxaU
8wkyyyITJ7iq8AqGJuleWUIqZxh5ug1UL8ST8jXNnA3eHl/5/Wn9YLU5RS+Q+pPW
IV0j0kYfz2ivSazHMDx107MNqd2LaQOlOhcKiL9zivCB/Pb2jLWCLurS1ZcISXSZ
IwIUT41plOFZNgbrhA9irK8PYtaZRIntL+o4Ju1azgoDojWfbye0CJoR5rGBQCTr
HhTMkpYPiWWD3XpghJNSHeTmuy8fMOn9CsCYgvt1SbA0N6P5Z62/Au2y7n06S5+6
eKqA83N7kbq0f+fphYDXG2DvUofcJ5JaX9T7kZWaBNjlXOIekbXo4HQWtmJybZpE
+nhQ8rtqP6ZMhTUtjo45PNrUGyWgGgFoN7c8DhnVFVUoKyVLpxUfLR1LHXPATdBN
0/sSr6XbmakcVEZ5pw6v4FdHx1sRbSfG6O/AxIbYT0E174zndsBhZvV9IL+G61k9
5q4Sahqky9f31gVilrd2/51V0pOG93C/gfbbDhkFHQmQNG/sHaPqpDe+hC/jUy9W
OFEngle+ZctoHcQDWuH7Lgo4tXRWfypR37bJB/aglAMFKnLiYcJ8R4iFNsQ0kdxw
CxiBMWhynqCSR2g0OQByI271q/zqM5o7mJrVz2S81lCUrKWKaCjBr2TDNPFT/22X
9xNqrMA/2Upl5mFKpR+kw9nGLncezJ6otdClymDtlIxEbGi7wTLRA0POBQUZ2yPW
KQtsGfpueY2H+yjr4moug4gc2ZfknQujKuZLU5Z0PyqE5V8N7Hk4BQmgQTWpLQzA
Ug29f9wqyyT2ltfd6Da6jvzoZo0XKHGWrQ64XbO7ng4/lWMh5QW+UB0PdKBpfs9J
c0xLys3rRDv98Vg6yNCu2jAk8hxRvjYpZSgznDQvB5vczFdxYcp/NP0R5T4tSYT1
EqCl24ks+mK1Den5HcRBaYMTR+OdzOF9dBXY2by6BA9p2ahNrMUKnfSnq86wRiGI
hOt3BgZSXCq4+b7TJnFzu7mOPfRHwTnlbC06cOLNtJO+UmV4e07s1DiiYUqFVWFB
aiJx0bQjcyi65jqtPOLIdFl4Tc9u/ykg7SVcXXmf7szsVyQS5eNjEUPGonPvlsBr
Rxq3Zfki0rK4/e6QacCwgSDNR8VvQqieAOvjHQJDzvFBnIT6hKlOQRO5BcMFbxop
YkmwVCVtnLOs+Dz7skWg5z6KXKwLGkUClGZ5Z5FX/9abe/awAm4fWq8XYASewmkJ
zab89U3b0Fjy70dp8APPysvoOcGAuWZ9C5zxsJAvVGtlKeJW6WxxtZU1lzgi3jFn
GdYOSBVU+mzQZRZEx+wGZviho6TpQOlHqLgE1n1aqY1VmjXoQ6lLzk/+augzDTOx
t/AySFO4DyWx+iSFe7tG9nrmcBsRWhsZaOQFfCZo9wwW/ZhUJArso6rncRJ3Z7qq
X2VIyvdVAdl8T1iKRMMS8uISmYTBCv6pTyQeXLA1k0y/lsDrojV60o/USca7VZlV
6fJO6pGCc5HckWK9hVcoxekWelT7y2l2dCB0n0/h5f3fv59EX1RMVODUONMPmcQr
uKLzlqPpUeQadZZP20rpj/kXknZTMEfAsfKT6uo/onFWggc+3rIF1KNAqydfd1nq
gw6FQcMHPSSb8EG7niwUYodjtxECFdD6kuv2uSA5ZWO3LX6E1ZyD0Z3CyvVZD9DA
FboEimJgqGelou1nGfv+sioFBRQkUjBnUhg3jW0LHdxyESnKAr3ifISSlrpTDp+P
DkYilr0Ecr+1iPV1+rGbawP5GoaVysqqsnPDQ8ka785RntjrQUfgT6dWhcp3jqrz
K8uAQV2HowP9V4c5ck6NBUtTf1NwR9YDaL9wR7jskRN14U9K54EwQpxuWv9g70L9
aMf6/9pZhdLIRudZ59Wcv916GhMJ5HJLPoIBD3TSykLI/ovNssAFdKrC3wXfhPxo
XSvLwdJ0WyrqDP1K86NVRA0q7DcgJUHmSVmlF536zkWyVc9B0GQk4p1KXDIrHQpz
J5ifyAPPinIBfHWwUtBZLgEt11b3pMkkgVLovl57Ajt1bLlmHeXqIRZatYSP0IwS
jN6f6Yx9g0GLh3eBlAJfjbvzKm0YUXrfNIXhKv0rGP3ewKDTQ165Os/YymVSFmQm
0SZX6n50vhE+lXrM8p76aN/HE3M8sm2ONAxFpJeI6KZcW+1236Ccb6mhn9ya2Dpi
AbHs5DL79IWSOt7ypcqC8qQkkFm19LZKCpQrQfYn/AeN5JA7K3hMbH58J+OqY44E
E3R4YwAC5s2U3yFZhjfpl2yEclWAyOzxk5GTMfPcWoG7yF0JxsDP5MvSftX/719a
bXJ6Nutjb45kJ1qt3Ai09sGFhGFDQFkt6ZqviE+djc45f/1ekR4eoZWBhnms8VCB
tFAq5Ww121R94eg6DN6vxok2kxiU5GPlZWGlWjBeBMABX6B0EEYJCk9SaZBbWvUY
4RxIsqK33X5GAdUZ/enZahqS35IPob1IemLz209SNnzsAP1jRA0R3seJuR3iPk1a
R0ZlSIb469Vyo4QxSa7x0JTdtQV3l0QhMxKpWJlJwaE+5Q6LyiMGPt4s4TC7hQJL
UapoKFhrQGGMfwwDVRGQYYc0xsOb5T1UOT7f2J0081d1Wiq9nPaGnXUMHvEaZZ7X
2/X983YDw+hMzBsPWMSjQ3birg4m1qy5RkBh4k1UK6Wm5kc7SEn7tk169efIRsNI
4qAx7zkW3CJqIuW+JxfVF18ziQdomdYCYqRrz6dBiOVv1IhAcyKYH1tQKuZRFP79
gSs+qbOiwfSckss8RqC86DZC5wK62Ije9hrvzPloosMhYpOS9kIZOdWAosxarYjt
YuipfR9pQqpc31f6tY9R0MzHI6WRZB7Io0MspQ5mdVy/EL+Rnyn1L5hXZoSmZJze
V7dCNh5Y1dclRTQq5neH7rgQOUu2w+pqKXH2/le3fEx+tto731XhDVCk+ANReLyi
YhYWGTEuYalaDOrVdI9ztEhtvmFdadHqSMCALiVbab5ZIphikVWe/rFIhqjulfBN
kFozFR7y2nxzEIeQHB+rHAvTKBdIumquSHg53jB9jq1/dRc6ZmDPEyT/y1NLMS3m
TkCa284GygUerJVnSr1JDV802yHUA4lgbhbJkeygQg50R22udKhEdOL3WZFrX+q0
F8YDzV4WLjtsaVDScqIuMTf71AA1o1shPWpUaTea2rq5N9IUKKlLOsKXnkgfR155
3o3dBZ01H9oggYU2DvDvN+oWGOgxYWxqdv5mHMzz4MxxQowRaHBVyYFupuKYogvM
M/VLsr6+t8PV1cnjIsULODwk+KkOMvwvmr4K7PVqWgPQC7Z6ySyXkvaGDsfZN8W/
l478yaR8tS2oSpB8C8Xkqi7aodcWYgTz7zP7k4kf6IEPYe9ZsiSvhuFQ4iQpX10M
PlhEt/EZVXQabB9ambujO/Z+sSrLSF+zIHNOBP9LnP0b3v3mpKt3QDU0zn3+m5Kj
nHhlgsM9Ye4Cn6+wQRGr13eSJeKBa2IdVylnJu3tVX6FGKwd/UvSTyKu7j02NMot
tZ39FC7zdynSmCVH8XDZHUOHp1VSZ/XWQmpjJok/bg/IxR4aa6BWkZYPwFnzmOr4
2KDDJIjUXMXMWT1rOEHXb723uGXtQmPLCsMpDnQ9dylPUtvt14O5g9CB0r2AyjZG
V5w2rAqOJ3Fs9/7tBc7/gQy967th5hp4MNdYmnku573cR2GERBbAzNl/q6n/TmJu
7ITE8B2ecX9Csw88YPDPyqdh7Ok4eLnA9jFVd6M9rK2MmpEHBHNTY5VlGmVktgrQ
EI+A91KTArTaveiprQrBpLZ4YC8oDxUVfVSlk9TKom1waQJaUZ56STSVS5g5H5Dt
wHr07uU4WGuFi9nqVWkUoNqWOxvH3dnw18axl36WO1+GnBsOKx4F7npXicUe0Wre
DvD7tyzv4rKJUykMnjjKXJV4oEInoHBg6v3LoW6KYICGAuDHBtDzxT29Xv0PT/F0
GKXDyMXd4Ew2ODhovYBrGLlcB6KY4/PpHO9aCCr2n54eCVVs7JrM4TUWvOKSZIVJ
AEZfS3wrl/eh0s0mMwd5GwPUbwB1GNKFF6JP5bqG1YrkLAQIf/rCIeESl5wDMR9+
DjirVFeNYUimaCIzI7G+juJA2qbiyD10h6FrRLVGzZ0cPiz1kLwqZqBX0zMPUYFz
PrDgdoW0V4jY8DWPGguxRkIYpS0eSTKlyuLlbLEcm547ehfSaDicWC5F8VvdZqSp
bd+fCD7RqKyN/EDB3OuDLrQgvYEyZqShf2JtiGh+wcvuThdThU4K41lGdV/BK7d1
ektX8gC4KtXZrcrofKqNW4Vh8BBc7Kqxq92xBu+A0Nt2I7GIE9qZ4YpK11SEGqen
OZhVpHekThkRu1TTlhC3O3pbrcbEIt8hkHGyVJmeyVJH0H2ftrzYMR+mRcsr3rsD
z+aad1/EWPBq1MLfCJPjRqqKys9eOIKntixC9BEkLd3aFmqQSw86k2llmzUSclY0
XStwzO3H00+3Z8tpmR5xmFuAvfrDgoaHnP+PXvnIm/nfLzK9AxFbkiZ+w1xcLBgZ
Dcy6gaQbPHY81vEPfPQWGwUk4pIqnW6J1+92wn0z1bSYCk6CiUpcbFLlsvtoazLh
8Lq0pd0zve7YWgDREh9xPEq1WMGDPx7LrhCSlUfw61snMfMl2GJgp9VIf1MF+ciB
BXE7edKuDo86lY2FdulzxAkOzodWy1y7y8VLpByzFWqaZ+MpWzJbt8sVCaWX4iYH
F4Qst8TGdT9a3g9MXgrdEZ8b30lUuzmfi/4upW9iQmifDcP0DV6fpeaZvgEb3T/N
4UvQmDGsgbthOUyq+I07EsJFupDDxk4et1Uhj4TQMZXSNYy7FhAmZnBytoXP8Lo+
vV/tv3Bdvo7HxbDKs83sm+z/ph5dnshvO8CKgTKkywK4DQ9xNX2ysnR1eD4cd0mP
V8JEPOoNcz/udPBojk/w2JOfWttZgKhChuElxlhws3lPScuK/Zy4nLz6lqmt4KXL
FE3dzBgcDN01DFLzsBTb8fAOhjOsc7aXbHC1JwQvkiWJmIchTkZU0OdNgpe3Oglk
df60LZYskZxWm+bePoLSOJrFTiG1tnZ2I6jCg1HB/n9BkVeuGS3rxfBVjLaYDSVB
ETcQT9fmHvF0gaPdltjFb9S1gYTjoDaPw183D5tIWIkVQ9Nu9ufMBIfomcNgywX9
BeU4Br24OnAWuwGhnev1CWgrFi0QJsPcQTx4h5Fm1sHNXIHKNH3uRCRwRI7LuMSR
i79ROiCUakVLqrVhyVbCTWpF64LEvy7/wiStnKFgcnwKmhxPOp/erfI1O+Vzvf3f
UhErppFSunJ9AiPlJCsWlPFsUKfogsg0unALHQUSe2YdnV1TD8TJWqzNp8gcB2ii
CL9YRlVzU1kILgI/zfbajdMMtx8VAzF4kWVKiV/YgPwynewlhy3BYVJ1f/9AN/NL
yemUY9jQV8+iz5QdG2fpcXrb30R59+PksaiMRzVW3vmaMZZbMyh5jImLtwMsDtp0
R1GgW/3VcDjByXUlp20+i+MkYXP0U66rGKsnaXqH6JA+C/CMqIQ+Gsn3plAWsfrU
Sepn2Ek9+Oi0dHPRdnZeP+0kjwUdtht+YG1w1EF+KHdw3hw0RgVDYWjzvTyNpe/D
etPrwzZ3kJ36EapsYbiNE+x7HJ2aHCljYRuTiYmB7+ZstS2Mzyu2sdP+Ksj9iVJn
jBerQikE5PhxUPwMHMznzXtePZa1OihNoMsu6cxfRKILzTUeYTiC9unwaS7PqJ45
1MEslYUF43iAdFo5cvXdzctHZ7TAVc0cD14SUSq88bw3FONJZYavDQKXa51aHOnL
JSBfOk0NvwCcho7bWK9Qq+x0Ry5Ba1M/i4tCuIxj+EIrOdJd8g/MUy0C8IsdHHQG
vIuSiHpgqRUmyKXb9etgzOSVT54mxJYUwouP1YrixAdnq6U1GGK0UJxa4Fd7LEhU
t2SK2V0go3iMCJM38MS24WtmNwZG0xgaHARN7puT3Nm0kCCqrJVG/SQF2tztBshd
SsEcVPSmLfCwkbduJpA24IKKOvcmMPLTLXt3gIZ2QOoEqyA/PrqdfTREBJgg1K/3
11sGG7+/8rRDs3zL5IyjwdY+wfqoNPf21YSVS/KgdtL9eB+L4ETlQsH+XtI3OBq+
kl2wiOrTEV9YBM1lA5BhopjRFQVTldVNUEqw/0rkIvR+xJ9kZuQOKvMUig/frKgx
sKM5FR7KrYbsttsl1pWE6FMutpRBMb1med3Txl+fT221QMoJCrQ2vnVXmkU4RAVv
NI85nQv7sn4WuC2wH1EpZrTVYNbWv6nXCrBJxdR/vkj7kJL9YAilX2iSL4bUPlM8
IAkLwWlkE6F96kL90y3+gKUwF6IbqA5M64Tr+eHOM6QTWujTJHAe9RL5at0+uJUl
JOvUgzbkQm8lxnJAFYjm0+7tNGoUKygGnT6Pz7/xrscgujSTNzYmb4EZoStqIcy/
RKDqcI+SmQGn6niBYgdQKM2PCp5s0gFtTIAiV+SlU/xQdnkVR1y49UQzYcyGxR3Q
r2AMC49fJkMDzT9F19lfhgOfXLsfSg5T0dAjzdFyYrq1F5QiYvmfQAwNsZGJ0y2F
7hlK8POWHgDBF7i8/e6MkZ7ewlj+pFnQhrUTPaRXSByKyBPG1QdJ57x6O2cmQa5s
meWRnwupNNi+uCqKnFxCXOCgnGY5JvhM0ZeWMAJpMiH4Tzzg/D5JwmRAOSncAEPk
3i59/omE5U27DT8S6+XKP0H72RWZbVaONFfXxVAlb91MkR3Vcjr3+pJ/Qoss84q3
Cpc2hOwlfrkvDOXoIKe2aGzbKs4ONrQNiQ9wRIcV+bCUGE2j7PSSzEye7/+Wmx1T
VLABlH2VnWWknXHoSSQgxQymWg4CbU34PzKd0Njt6Uuuh9555BZobJ+CvXzr8e5M
P1tbmcKjBeOO7Ci1ovrxRjw1nQfVOJz3WLJSW3EpN5D0GNfU8VIZehwL1AERGI3C
DejNItyHsMX0ZvJmvHYQa14NIAyIT9D4EJFJMh2KapInLqg2lI0A7UTGXHChCvXB
eIbLPQxTz1WVG8OEg5rr4Lu0NRw/uX0Vwtbipn/K54WDuyiuh8VMHvZJm6B3/oT4
1R2NqsznuXcm4ZRM43oMlJ+Q6EQ34tALXGbt8hRhU5IuS/vOqP42Rd2iAsJGHy+v
sYyFAlLHppaanYjX19P5NuzDMjtcG0WIO3p6MQhyS6cjqYXy0cvuZaDZ7mjGJspV
JY+WlckbUAYtu+nXu/pGw2e6TB1MArw68F7LNHuUMJYvjyjP6QFJZnYD+SAWeoTz
6CJxN/BR1P7CQgqsiEypa5PV5Q4BTY/MkfSv/GCY/F14Wqs27dinx4jTeStZc7Ed
Tjrd5sDplqzDjOL/Ch1PZrudC+stPotUybkxC59Lbc/5B3uY0bNPhR+M1vY56ZRm
dd+rMyLa2hD4upQUxI8V7/vogua2QY7N3dpzSrDiy6W3/N3s5gCkBXsI8JsymAAu
swEbi5H4v1Qf+WO4qW+AX7ZFJ/22P5Hdx8tEzbKyVJYQWZPqSTAIoW16M8VHplPJ
iTDEmotvYVjHLmx9syoUKL3FxlbI/B5N8htoAs8j6oL+IUGgQdzkWOGHxorq77Hi
z+BVDtLmsaEdkv6yIEbV9GJgKeAaslJBkYbkSz7MvbqnEmbmKZRLi+9zmt3jR+IM
NrfEze1CY9WqyefkhiM/z1ZaXmtkuLEiBKKXB2ySCckwHpgp4uiRXu8P/dzyMYGt
HGyMZ7hIUo4ZKhKqDjwQVzFrhi7ncxS8rb/iItHDolvyqeQEVPAr6yNa8sFwSt9M
cQPRyxibUoqTz/iehzfzRIKSsTIQl6jVGxpVBiKUeUPTbs0afSIztctmPUmvCuos
mBhBJdM2wELXJjozbUNe4D14EQC+jc8Qn7bzd2qkmAZjzuugPnKWLMiUSJ87sxA4
rnnSk2P4G/+bez1aK2EBSqG9E62o0lwQkGLpixfXfONDdWhxXL1+6hraVHwy0A5F
CQf6YfpH2FiezTqfjHUVNt3QjYj19VhGru9gJrvCvbpl3KIIKZQoDHgy41l2BhYE
eCMy0Xj9OLObyWzHxfsazz0Oeq1z6e11BOXgH6nGl+TiS7r4p1ggRrCaKsgdDbM5
rWNSoi8BuZQu58rRW2+Zs6yavtOB3vTmaIFTrJr+M9OwCcQNKBgv0NbHAnjFfFbC
y0IyNPWv1TJOtf74kXggpuXlm4n7TVLetPHfXe9f65YdeMsk9opmirN6Qy3H18Gc
fZ9KoI+TDAVelM3usEyhPRTHHvo/XmCODXVvJBlMCTiodS5OhE/XTnUfjm8YxSnI
qKZk/D4KJFVQjlf12tcfjogGucxySBlGZg73Dg3fCl5AabNYhlCN0wnMn1C44+UD
JfeGshulvEbBzjhW7LIP0U8/6wDR93ZIqAaNy4uo+MSkdDtnmuUEZZxpulDYtUKT
Dq5kb3n4cUUS1a58QA9bVkF5jFySlGObBA/xcHjnLRNkWQRfXxQhTh539/FW+cGX
9uxiiuhMi53GPahjI3QOw1o1oGVHMZofY2ZWo7x8gf2vGFWucNHm5o6zUN5h3NGr
0O+0ge79e8iwDvWp8AKHBhc86cpNcgM9O1MFzBoYgpTIq1QGEcTRuPDYUm2JGTEP
LVzHMuWIaDMITJTfOPjygWkSBYwvRJ45LoCM5N283/aUbsQqnohGNMSJw4r4nV7s
prRtP7Hk4XW1l9I21p3LugFVjYg/cxTFZ6TtkbgMb2adtAReVNqmQgs1pdFE1vWq
tQgh3ySwP6M5etKBRoplqYRzQ5sU2+R93kAPOxLgnCP5nc0nJvrw7OAzKK7x3Xpm
KTnymFypmPo0JddxHrSXI/K3Bo7iQifSp//OtSZRJZn3ygLCXoYjY1nEMReGIiRP
exEwxqM+TahXzkaOh22XS0s+aFxFRphUMs2a7jg4A8M2Me9K8hjUNYlj69E12pEn
ZiCGWiKrOqYNf2HlOe8sbmEUJbC7yTce4slxOnkWxvK8O7cLRzqZlBoJMHYNSSkg
EdAcRthfFnTqtBy0bx4jQKWingHH3YziP22V+wU8+BqLwfT6kgLNHg7BbRtYXGrr
vFiLWK54GKfrzLhwYXzKXbFCBxJtOzFMy3AS7qD9NdySy97z21Uwl7V+0b4cLCrN
ds5LAMx6iUSrawdXctvx6HWiGXUWzWwwedRuSM7yMZdfEqHEUpsWXDrMonaVDCNq
H+srAZlBvjJg+2urkUsDL27cL5+zVO/B0fyyfOEsE7sDmW2mST7sn79OCanjK1Le
vyY7Or1/ES66YSEOSfILbZvdhWjpLZ5lt9NVa0EgnPualnJEty5cKzkr6RT+eNO7
Q99I43hgDZD6kxguEiUfZHGNvIASkfOhzIHI/uCcjNnFAg9I7/NY+Yazy9Y4z/P+
Rmy8rrdPMAJwW2hTho+2QC53vXQrotKCM349CllM5U+pcr57vUigOrStCVnIhCDp
KFx8/hhws356f62tGhZAcfjeK3/iMEwkAAVL7FZfNeS6zMPZ1rDkCM5xSGmtRbhZ
8/5Fb8vJdfk8/iObJoLusDz9N2xlmIEmXKTPT5vmVk8vRwe0x0AA66SnjQmotc3h
H1H7lqVYB36cR/uT9QIqkoD63vMdt6iBGBdHdVSXDSVHy92PyGce8LDlWMR/pF30
/6FPfRPSVZT+W5y4AnVrfUBtTmD5v8ZylHDDmT1PtbAOrBJbw7Sq8VSFHk12+4zN
mJMHUjZOr84ABxLWidn5oJoquIJLJux0YdK2yoX/8JCH5+dTTzsKWq/WX+lYp76K
B4UBd5ld8UkeNgFTwjG12Y99REkeG9L2c8yUqbiDHpC1mjLhlZpQhV9b8/qTjLU1
DOufPiN4U7bUyQPbpbXzMkFvzMA1LwR2/8bQUaXqgjAjL8uhljc0P2zXNFyi/Dz4
2/Mzb30W72sFW0/KZCnhYj8rf9jGhTdo8qlPDfvZxzim1dNpxXwf/EySCGxXdD00
Fe+9iojA3j1mmQYotSYy+uneOzioy7g9BWYtO9y4bdES+lPB7oeD6cacBz6yLlXX
/YQF4xXsdUA49ihnHCPgROesaTk3vgXlOUdVvVELdal6wKDapWN/FxUztWGOI9pX
2c8Ot5kNErOMWWCBytqmgl39uAN0NXWstGQmtz5SyUUtX8xId5It2DPJvxDiTzHm
mjOICn8rXtAk0hzBTJSofij4eGz5suuHu0vOGpAEkoiRVQ5UCByqLQSM6j8GCiz7
AbwFlUFYHPVNxVo06aoVINis67hN+DdD4hFRp/9pWIdNkUl7IrpsD9TfMzdemKLG
9D3ekuST6kAC5Z/XGZCRWbKmWMYK5GTcPHahSvjIc/f1Ry6UALsGoDGc440D0uPg
sJMVYyN9cPyCNZOarAtmqeo2wr6WTDtz8BJxHFxJyLMe3XqU8Gkgq4DiGXNa3QGf
0iujNVrjZDCgV+j+y/K8bxbjMkz8P5CuQjd7kHa0kU93q+VJuNfHW5ZkR+9R79xn
l/KBBtyJ8QEaFMu0dQz8pYtl4H3mMpBVSyyP4AMp+84/A+8Pf6a/CydpFgPRVuzE
Ngg97IjLQ0FwGdtTxnd4Uwm8VkW2DwbPnCxQq+h9oYmZ1/RVHGpt1Y6V2d+ZdDYo
JfGmxBNyyfxIaZxORvwY7yl5wbngiDZC2Y5VsCkdjtw6vj1bEmaOeoIYKSe6tQ36
3/KWq7aT2CDeXIB+03eAdgcXMolmYLRxZaClNE4B6KDAXfgeSezQmYXHnNXkeLm7
0500TMZ2lNIR96PJgMyqyGXoYB3B3E4HrcykNCVrDfY4YbDYPvWUsnpK7H+dQuA7
x9/lIgDX9alBSEe3tkDTgEw3HGagqx+ogWkby723mlyZr9xz1IpnmrMNsxA9Ylix
ssPTMLcHW3AR296AID6Qjp171VePaZ5NRJfCkAZsuY1CMb9plwOEb9cQ/yTPVNux
ePLg5Dm0po07q1HBtZMYIM4ZcAso76ZRIgAJ4EmAyb2pssKGwpvEwaXeLKdltwy9
8Hrg0b0Mr6kzW2MoEZy86Hph1bFk4yc24D764/Q2CiQMFU0hzcLBxOlozOq/5ynr
jtVsPpx3y/HFt/xthHfIdRFLFwwnSIDR6d2pHevsvDfFTcCR0EdEYCfE5xNl9HhP
gxYMVPrEkqQiq0FxVU7dVVQpL43ILdz0Ce5rYmmDaJEOIq2sQJSmsVRQ4ChGzysh
bauT6bZfEDRKm6nWlWegDCfLW/ceYhv8uwUTtrLT+n8D3Ava9m7JgMJrSiBVWIzo
Bud4NXUsMURAEPyHysWrPd4jH5fVMnI1dzsu8M52IfSFknNTidAtNNOIfljZ7LGY
wbTQnyI7PFD6JnNaRVhWbCFAo24R80ic10z1p934RxyQx/o/WC5JTE7oi887jOsX
a8EJ7O+/XIGKGrghw6x0JTV28MHiPqwt+xtThFoDJbpdZ3dcrOWKSxFnwQ5qSRuB
nNDRLImQnWNQhhSQO1EZnouwfB2OnqR0Z9tQ7k6yj+sFZQAuYZhV/XeL+YIrZkQX
YjGRkNqq8ALdDYhVhGdMo6ODf2T/6z/FXyS0+zvBJhMo0aeBOnRz9k2orYIhtKAB
5hgE4+oW1UoVF6sgGNO44BDVFB/rASlrLY3ZkMGkpFbjJ8VWfFfcoAGvaq7FqihN
scdeg9bWXKjTBcXD+lExzetX1vbEvJvfXXzg1++Dx/LyldKg7XtIzQiv4/AcOyZw
eXv257g9325wXQWepJpHQk1uLX+0D4UOTMfpHD84KKHsxe8CsFDoWFocubECrYy0
GdINKxsu/IR27Kprp+SB2hOxhL+8Z0Yd5T1ZMwV23Z4StNmXEzEFLtWlzqVpjUeK
btVFZvK3laMGaXHw53NQ4TGqEJf3uIwqhhMRpklkiLYr8QwUjrAP+1dATC567p1r
fO5d8InjCCnO0ABtmTyGtsOdbIzoq7DoS51qq42be+YHS1TImbNR7oSWek4RE3bS
/JMfedxB6fcdyVHlzU/06Y/+JoVTSGDMwIxYtGpqqmK7nXnjlHTtivgzoaD/spnq
kbZgoCadQyqKq5WFFL4DCFaDhxw7558paREboJOq7EIprkMSlBOEpj0Drc315TTX
aZavAZbWRmwJ8OvbbFnjJwFJiv2vsLMb4srhN3IM2LYoM62TAWOVpFmN2SLRSNe6
Dnj3wCJ04QYPCTSXhBKTqkvaF/ZWFXRJ39XgJMYL2O34FA8FA6iWi6QKh+eE+mhZ
LqnPy49G/vpZc290eU8DFuLvEzeNJz/FQGqognTQ3X2PVWO7a8CSryOi3luGlLSt
XmZRUggkpOALfhwpn5cfAtwLI2ppmz5qChY38HKJjOYRD0fGbnSsOmjeZQEtxuzF
2PRgG8t/EDb/c1EyRzfWejrEgjCqrezRUIaR/llrvrAXR2/fuI+XYZRPuBEkDkf8
kJMhJL3lO6+PBVwciANbw7e3GuhmYc2y/l0wt2q3chl0kLZXvsU+DttbHOsSuA1H
aml6YEsIox9bJ+HVHE8I0EchGgLHfEJEHK+S+3dKI9aTAjR3yH9afVikxi/hySD6
aw+y2AK5bPn2EjGEkyBroXdDFuenWDa0Rzk1sVv77mHWTeBbQeo5ieh02jtnBQfY
560VaZOWtWhWcPSY79Jcg68OJ6DfihEpCVMM+7xpIKOn4S2gPP8p2dAFXdle/EEv
xXe5ntAm1wgWPM7mKLyJkcFcUiHeTn/JGeY4YJFeT8Wu63w07ni+/IXXuGViFYhL
C9KV92aICVPrCRxG4eV6ureRNNT9kg8frMOnRDA+NWMu7jyH0tZJ53VPH44BPvs8
qK9DpcTA5DmPXQuhAUHHyR7s+A5vGbS+R8LXM+W7uSbU+8VHESTFxM2b8qLVJ2PT
Rmb15sV61nO0geNp92zbYHlThX2Jfobkr53B7+v0kQVAr74xAQ3Za+DS7FNP3MD9
lV/Lt4rNHeEAeZq4tWHBf4hnt1CjoORNu2BVLwn8EOcPMJF2URma5DojMiXGGgG/
6XGAiK1YEoDoXj3fL4E0g1X7zq3gzKtMDU07t6luBLcCa8rS44d+wLqqQ5T6IAhj
rpc0s9JSf4pziWT9r3j9VZeVc2voIEBG05eU6xlyMI08ptRw3wqRU2u86/fSHBy1
qBCnvZkjOxW8EWJPYWYPFwkFPv7JqNO7eltB1tL8MP71Y/pF+ZuNUkqOLi0S940f
H4TMCEhd3OcpKIVeOLNkC3WLYSKg4gapvwCtSKMbSROzIrhvS3iuFXA/3vn+MXnj
bmmTTtl9TyoNN/ifyh9WBNrLnnBGOous8YT9RJBiRhNOYNl+zpWEJBHsQ0kX2e2r
J3gRD4Ds4FtDYKxDjxf0RpkWBzYM3b1pFce3STRJPURVisaPB+BBEqiFYBTKMr7d
OotbyGd+FxLzKwRxlXnGEkC4D2QiqdwqPl7L0drSFgMwF2MokmGnotf/j2l9//5u
pTNDvX1rKnQAZ5M0jYuNBFA5RsCRNHTto3pxVfxogCkjFFqbqXU/DIXTbU/5Avje
QRrEWU6qaGZYqxP959xP4xiv0KXYrzt5XG+4OkLhO/HyhZL3C5/544NxCUvG2bfT
Or3ZhQd8g/0BQi9meXLUNE3PARLk1MrS2XgjexxBAJ4WLhPFNFc4ZR9XlJBwq1Xl
0NG6r6D9/w6vmPDSD9BIAB1OtMBDH5l92njlfMSQ+/m0CHHMVbRztuf6O1Q0Y3w2
7GxM5hO4bVz+x3Qdbvwr2pvVaKsN3422GUh6/bX8hdowFZzqg2tsMdZj9aNSQ5bO
AKcFc0cea/krUH/aBhH1TZ41td4JH5dgTaeJ3c995YAYtp4njAJqSWSfMAfWbgxB
fIGKkoYWqZ6i4uoy0pS2sbSbngi9HLalRJMfaSQeXsRbd02tVavqNItMV2AlUixL
mE9DE+BF1jv277+Pycx81PufNX5LS1kXEJaoIUTYblkfIJN1MKeUug2QnxR1xB+J
S6r7EGH7ta/k1cikXYnNNffQ2Xy4giGKfwe0WSyRV9gbRt5D9LG0S7Amt3H2h7G0
tQ/NS8c9Ak62qvK1AqobL8FwuaXJG+IasnHKYGfYcxFd7eisr2OajXMYbdKhyagc
7brQBihceYdWqidicwF6Br30ZuCtN8lTxo5GjF64bd99Hfp52M6WIMZUob6l1H3S
6QSqPgwNfHiEsfjKtibqDoiVV4gKwyVo7nOM+5dwk9NKak5r9gjfADYTUCnDi2V8
+h98+Ib1pHRUuSINiWNiwp8Tb/8YeW1rDSxHNxjwwNYl1llFSaxUkFzn9Sd8IJwP
Tta/3ybRrSPvwj+eDUvbLFNh6PByeFnwZlzK37Hl8iT87SZUrTH3jK70Xn/po7fI
nWgh6oCt0e6FQ7eEBPOpynkXjPEVaExJ0ovdAnd2UE95RKuKyfn6x/a1o4C629+U
C7eVpxm3/EgoO7nyIh4sR7hmIZ8wthf2iA5lCexy3x9GIPu2Klar8t8zF6Q9GphY
pv2f6v0+OVxskF2zj3G7a3l3qKRkhSJAE4f4lTiV5IH9mJRRm5GejoyByLR1uHoh
gcUu04baWhqBfkLNFukT0gO2wjJdQNtEQ3/YK5J4yD8y2IPwQ8VzNlBSnj7rwp4g
c+6Gz3SOKV3Mmxe+J5DtVTl5WPlGTLN9dwhJIv7D6ALl5sG7JKlzvbY+QVd1EZW3
f+w6zti3loHD2sxQZ/hXVBO5O84XIr4M0GbxAbWMsJcYBzuPT/qjtiZ4mLjtwMzI
6v/2gFLTB1rd01bBRb1ozw26/nPbEEIRiD3EsfwHFjzaDzokpCN9SMymPkcb7UNF
0wp7wrmagkAT/etddUdEioPF9CCJm8kfdWlZOY1CQfXc0RjRY2gYXQywx6V1wFMZ
jFeS22Aw/BW+d2iOCKIQEmI/zH1odSKpDt2VRLKksaugLUSP2Y3ZEsaAeh8TYqR2
YUbWRw+Z6zqvO/E7kaRUyYzzyXf8VgSqdiQl5NHaXiTYNih0gWTcdH2l+mC0bH7K
64dO89Qo99L8GMYdfJzcsq0IbKnhumPXTlFYDIODefdnNc0v0s1WJ1WCKPU2R9PO
ZoWi5KzdCDFgjAjGjonR0g4lzU3ur61yUQVQnH2ny87Rz+GLUeprIRwnbZZpHQ5R
VrX7xnaLZu1PdFh4XOBzYVY5ec0lKeTxpQp79ehNIA17phADQPgqIzV/dvqec4UJ
2YONi9J1mWZj6++0/5cYggmyHrN879W0yNQu0OjRUx83STimM7fzcjrbtitYOWby
VvTIRbDetN8S79inAfjAXUpF6K/OAeHsqiHejSxO2o0wL43fjhlTGldp5QCF/eLP
oEKjXMM2cw1TSk7Iw8+xFH1dvv/gf7h3/NdYERECQ6J7cJZUiToEGVp+MXvmtbZZ
FQpDSzs1G3aOF7io1+VijfgVZVpOcaP5fN4uK+rwsBNKTzjhcBDk05Z0KNzWF6d9
eRs1GgFdN+7RI8tO8kP8wsxSqCDz4Nsakc+K3gmVPqpBLVqsO/HG6QM/25fX8N1M
DxWvh3BfuIZ2nrI7A75l95A+IHi/Jiq+DXQ9i67DiiQntLO2Ttnc2qihwprTAWaW
CKlIXyBzZs9jfbM8qkMWW9l9RjUVKgr4s/dvrgXx+62+irP1JInlZB4BJ8VG03Qg
gCRvUBEEU2HLv/99gFatdPQEzZdYb13uLfXxZS8VDcyHCmYEkuk7XOeczh5TRSrX
wXyWudMD4W45m39Qv+kEXwvJ2USIyNuUowB3rj6uCz6n7lJ4OtbY7mdUU9DorvQ1
ENt9O0p++y09TtgenGoekoZnvYXJ0EH5I8lZ4AWTz36WrvfWCJBNNAhIOz9Pm2wZ
AMF8PA/duli1ho8fdfDHVzUWfu8zh3aP9AhkJFe+Pbr6CW6uqqCj7rEjDw/qoB9d
+E4Ndn4+rbiJNHAC22p/X1RPVXMNb2zggKkUui8x7UVj5i/8+7mzhLqIGc8wwXJI
vozdram20L8StZD+TfYBBU8H7bAfo0TvSZ3egWD5lj3FdnUtfpUi/b6gdOsYmMHd
vXYRm/T40IYVCqzOUpCbwVknTbXp0GsGyLFC/NWb3ja8mrZb7KzJEtiQ2mF6cWQd
/rKcRfoJuVZEi5BQ8gQ2YNkDHt8iY9n2uhdFHX2dK4kKgmg9e02jzotrd4iSnR4f
PAhouJfKb4LKgzb5VZ0YXxmT2XdKYL9IKGPxisPmLvqMnz2jay2Tw4xDGQZI5Blu
km7JMhv3UbMXuipQM827CBuNSu2XJc88uzON73he5Jx1+ykyzDeIZ1EmD3l+rYif
zgZtG3n/QyZxIfV954uCh/ZcV1rBDYthyPp9Gw/L5/nys/ppcNy42CX0VmQ5bbNT
kMKC1UnaL0RaY7Ty1Tzb7dRInFsLAp+xMRK5rO8cGknAcScRl4CgVVAnKDKW+w4A
c+KZW2LDu+W420Ru9iL+0c+EwUlfhxmnm5HRVuvrEHf/E/tG37M89sgMQ+ofIPMS
5N2gyluD7SIRdAYgYIxAMCWdNuUjOz/3bz1FvEARWsoacrQJQnWu3jSji7AK/SSV
yUZ+xVbQDFnTry3xf6tlVlGMwGSs7q4zKGuS9mieLyTrovVnv1omu5kXJNJdaEA9
pxC/iJtw5zyABCPFaLOD4cXtQXnlGor8obzg1Xo87G5I+/09h+/GQeTuVA73EOOX
5lQ2BKddW3/KxHAlQlq81BpTZ2yMkeYI97Dz4xFmdRvqPoCXkM8yPxFnpkBzC6IN
VoMNnZU41nNnfBj5I9XJ0ZSBMy5d7Ie+bwqZpbqKh/88Onwo4IHT3c78r21UvE33
Q4CzEBL3GyujLfwsYM5VorxHXg3zI0GG+6p2onBklLmNGCD6AMtuucV9BRCrcfuc
IpyqdFpHhmbhrvvzya2DRwuyH+ak8WIAcAHX47AH9ATSUudFVKiMN/SwWh8b+PZ6
GbjP1XzU5YJlzsgDRGn4MA2YFKh+/6RpuAYzseHz7OBymDeVQ+7hWDq/+3z4DsMe
JyJl4TwcrCK/tNegbMKa/iZljH1lVfv027XcjuWDGIPHJgZyN+A9BpOfi2+x9KdF
x+5bmoLFZZ85V27XIghaKNB2BvLN1fJ9VRhimQZ0S0kb8d11L96RxmVW3H0DOxUS
dPA3ocqmpylaxjQAbVFduJdEae5i3iGrIqIlWS2thnNWtAOfmONOSak3Fl0yMHgw
3Xy6RhnFcjcCw4YA/oiRWaJifk1OnNm4khLeFTf6P+s+NniudflXwtgsp3XlWfAI
pJv3nOLdmsPRdNLhvOw2ZP9+3pbcO1P+BQq8h1q+s+13mIiwN4LZmmYHeEmTka+L
NKtXuNCtx6YlWaOw6S60t5m9Ugq+wf15l9+tqRO1oW1K/XSfzEczILhOzZ5UaygL
1dawRaG9ERSUzipNMwkLsRzlvwvZN5nLYhW2+iy5UXaYVEAblKWWR7HR8IJ7tiH2
yS2q1+uLyGqBdzAEInULCQ0pXlCBLgGX9bcdsMiJUiaz+VbOf0CfvV2+Hm6mOaKO
pkjRB7n1DMJ38N5WI2dyLCm5PM7FuIgQEbEV58jss7BeJjbfYBA0BZFiQTApXgBM
w24fT8Y2xeYH+aDjWp9CAHirb4wacH+BP1wftDx8+9P1Fr35Lz7UqTsc5BzOrWiq
FHKmfCyOxBt5qySuB+pqLhY0fwMLYqP19xsj9q+MaI7LPjSt98BFZiX57DQtByFH
aPxesJh1SgMxO/56RhdMBOTEgrDYS7fQJLr8JlwE7btjQFWlHy5QC/I2ZBOixWOk
r0hEBwgbI0qx5QmILY0ekTYXlT7PsUgl/FyU6FE8DqvtDB3CEEtsnpE02ansVr5X
FS4tpqltnXnTMQ4OvBonBW+05x80wzlQkdrARFJDE57yOLAHq8y288VnK8kdk+uL
3leELKnVPlsS3opE9AxZGeJG0vjRqUbx+elIG5yG2k1lP8U5BRIf7F8pMD3Ys+yQ
P7KqK/7F4OzPjN2RoHd1drZaEJ96PumOLEPVgHyxKxNpXs3r+9TzO3mIlIaP9WKx
6pcB/dMRIMD9Yvxa3z5kFKGo3aEEM/exWWhUvuebwW2R07yVhJEisBe+r/SidZ7M
DfrZYSkgcezuxNzwpTbsWXKwh1QkTC07ONSAwP5Vzvbb1UexA5SgH28CFlJGPu/l
0FrjGVA+UAKwMuXdO7kXJO28Vha+Q3gqHgzVScZWYzI70schPIWuoJjBvJYEZ87g
urMxHgCdanQsCQs8YJywB9sut+LbsXKxR2Jjg8rr7PypuXPCRlOt/Ikr/CdX1ISj
1dwkew/9t3/AkFkAoqgvZ7+RFtdHFuUZRwfsdT8eZsEDlgUDDEswNWrbrOaAOah9
fM8FXXCXSUSy6cuH6n+pw1XzDSuRP3BaIzlBFjfA1v8j8cQ+6j5MLQVuhUaWfBw/
dUFN+FJ2sED5UcLheK0tbjoTVkVbhI0w5w+C9zg/0e4JfbRQ8qU2zpO0rJk140n9
hXWRy8noOSUModuPduSdkF48cldfX/DMeDKcxAbPGP2I8f43oYsy7tD0SR1T9FPS
TzTbqmu6mZXNf4ru1SVZl/3lf++lRS1oLZH273gM8Qf5zJODthYl8WlrGJSv40LF
tTPxUKDV7UsAqchwRZdFAydwBlwm2mZCTKuCq/QVOmukcledVSDWghsTBu+8jFW+
zRd1ILLkS2ZRGIbTG8wiXURDQH3PxEokOclmIk2C7ASibs/EhWM461GadQdrQqzk
dstiREgzBWr0MkTIAYAqsc4ul6GBrErfRr6Skm24eVNaROr3QVEzzBPfDkFLpfZo
bJK1kjBu1ixN95j+3dZwvhngJdRh1QasMsgBvz0OwRxyAHpIb6gGcBHOxyKMOawP
zLqqQxOVbDhLb2fz2M+rhGz1DjhtpNm7TcPBu+1WheMSKfhf0xYTu8zjt/2O0Tdj
klrmU1SwWeVVsTduUz5Nl3ZFMSN+A+I3XB/cLv4SmGw3P+0nh86v2TvXttKzG8Xh
gom3LHWHhtnd1vwdksiXtc//1i7TBKybvjjWlQ1yzwzKa+Bj5T1kGuaIyDSPChOk
IABUXkNqJarjIT5JNDjz8Bcm3bartBvNGQAdbGR7jr8c6o7To6tDmSNdVMi7Dpeq
bcl+Mcz+pmzVTpY9psBGsswyYSDXUJem6Q+WUsvK52o81HcCN/FnHr/GnYnyeO99
S54rZgMCxAnndVJypCpeQZmCz5br7BsBqSkOOE++rKX6Mo8CMNC0OrntzzYQgmoL
1017E0G4o4VjSuPKA//VraFj+OwOXbokeBJQiCOb3OiMMZ/0dqpnLTRhOW+F5xpq
98PeG8tbPtuaLs0qSXDxlH1pd9IKbFG8ZHj82kWuhL3r3fcEWErF+hG6140GS9h+
SGKtgPxOo+iMnGFCCg4akLcxqovcFUdRXt/2YIJCeCYZgRLQoDRfMZ6To/s7++3j
xBPFq8iEqfLmu6Lvi4uhXFG9sdimtoyal1UydK8z60DdtfY9AtK7k5u+cy9tkqcs
RAQ197HDZWK8a5WosX2nldDr1reEEOLhtChx/sOd2t8APQ8ynYiTg+NaDOx3DMcY
RLIliDdPI0zsvhyBdYX3fv+5D2R8Ahoo6UYKYfYJhppHqqOohr+EA2bnddwaAbtd
x6CVKPsd9gM1KQ5Jmykks6ryGpHOVgRy7p1ISokf7xPnOe6AarUbRaNDZD7+m+Cu
GZYxF/SVw2tIhPLkDxc7jkHj4Rv/aeY+c39CJyANcK3rv+Vn7unpUTAousUJihfC
dXXVek2RztnK1GxZaw4DgpwUs+TFWX2ydEmRn23uswVjZbd4GLB3z/77r1wtMiH7
4jgjJyYrkM0t1DqHNDMDJkQuNGBsOpOHBPKbge0Sfu7A7xMLB6KdUyEE7ON20cqM
iTQgcv2NSEbt8FxOdWSWk+Knuqn2TE2BKRgKkhyQeVhuAgrzhCS73Eo1sbBygwhD
JR/zYxg/E82XRpQshcFvWUAojUf5ZBXhgnM/QkgYbjrKlFXTdDzNp36S+kYGvGhk
fO5Nj4SgYCbgywGpMiiBBgHmDS5dM0HfWDmiZ4MWGTgoD3V2z0z0eyPiVYK3I1Xu
M1UiFiQLbE1QLwByYXb4OFlPduzItHV6H1Pcm7T+l5Gqqj3jzonvQnbEr/rqnVrC
/tdeNBvPQ1hvB0195rksMWVZ3l7jaWx01+MN4XC+WrPDzSNVKcoZ7a6Ti6aG1+nU
gQ/XaHI2fFaQ/jP0ZnRgKSKqFD9l4Y4U0DQYDTIftZnPP36npCEJ9WVg1rwO8zYr
v0omw1IX8ld3BMZBG+JtEjUV47yIXRsI3lxlgJ5Bit1rFqUgGatDOAx6JpUKJBSQ
n7I1oFJOLA+viWx6RM5NN1voXhjVAWMOg9ooZhAtLMRrXnY4Aq6LTaxnAyr+Ajf9
qujnCbNk8ZapqDQn5jjhMF1ukmeF2k+vqf5X4+Tpcu6Sb4/jzscERKYe9kSuDuta
l4ugmakxf1WxNiusYWzcUsl59MyRkzD149lhd6dug5uRejms6FUeeECzQDrdiGyL
ppADId+siOazMw5jKs8U1Pna5YMbZNCzFRTF4gx52llH5abDPamWj6AuorwnPNcR
lzCOnqOkMAImRfYK3HUJGhYim5WwF+F8n2pSSwQR3lZ9risWZDjwhINptucxvuZC
vIhUhAp4bAEPmAziibMzODZx+8YUWUYIb8AQrucbbCFsQF8wfhdFmr+T2WoV1wmn
HOVP/Rk7Na9ePCvy5R6qPjFwb011ahyD910J+h5opKxIg7LEK/9NeLEobGScovTb
4rVPoNglURZzQh4EhJcntv7YQj+jEBQirsdkJb94yWpcZ8eIh4hdBlP0YYkowlWL
vukgbEOZW49NDkeqqNOoo+PJ8FMTu/IaTSdrgtRaTOTqyYTniaHfWCjJErxeZPwz
yIf/1d72iowgwXoByWZLgqoaftuAiqYpM/040ySUW/M9c2468SVTqloVCQaOQ1om
aSjgbp4x9EZjJ8/jubee6YuFAG7PJKXTORO0ijl4v7S2Z1XEAtOI82wE5rjJxxYy
4BnT6zytL4vzWzqIjzIFMe43vwqYftiifPUIK8IFbsjas8sV0qR+H6s+uH82eXoy
K2uTe4QIUGqbp2IL1P5dN0SelPlpIqz5+XpsHgX4AJHoC98X98RAEohv8z98s8Ld
92xOwWKH9YkeCoojpY17WxOBDHUb7MXowjh9KlGYMzsIFJxScUveArs3Unp/NVYJ
M6qbBYvfbjHwtBslbpMKcJiLa07oOYFaxwl9CURwWlVTZkWejRD7LHDL8EgER4/J
giON6ap+1aBWcarz+TTToTAyEGVWj7/dHvCGTGxLuCj9c+IOajmeDS/0jQMcmXH8
bcR/ebCGYixswMAsU0J2frwuJVpJoPdf/tgAkutnXu0N/E56AVq23rq3dt3psum7
I+RtBGKJHkhME7hRzen9+zX5hQ/+9BSDt00j6czeIiGXo+ESPdrC8HpD0tYamuWA
x8L9R3YnISa6YlgIE14nM9KTSIgRnvQVGJ6VKbtLbcC5kHL/Macdnv8ZE+ZrUErR
E7gpAeCZ9na0AyW0/8ZLXpfVxhohO2wQQH1kSUyI1jCTfQC/ZAVc/aDCq2YXIQqP
LZez0mChYtsgm/SZ5KRAvPbqivKpC7ISCNB0eHJOF3tFGhUbSnKpBOGlrmSiG4id
MDIpkuZkWO1lvxp2w7EGxb17pF2vpBrt/0tB4/3WoH3ldKVxPheZqIo5vZKb4EmQ
EB5yS1ds3DTGjKYrUBqZAs3o/1vqaCo0c9FyXDkBCiAi/oEmR/dD/W9gqi/RylWb
gFMcKRce0TDzKrVCNGgPdKzJDVmEKWfn8lhel4L8AJYaH7JN9FDAOAJZw10R7gZx
OLubVRa1O6YgTiGi+UnRdqow+r3/QTyz6FEOpfKge0e9ngL3p1MbmcVVeYgUsIeI
K3fSywvSL1NbbsXaIXaWajVzugTYvbPYwb1XgxIWOpcTumUnNJv4eG8BZYXu7Z5H
m7nlr7w6l4oK/x/W4hpRwaoypOtQll3ylGZV4nVPTXH5aaiZqxvPxGSf8aiyb2AZ
91BwAk4ohg4yw8Es8fgHW7usjymxJ/mmC7yomD0T0DDD4Py6hX71G0Oyk4xzF+JT
vsd+rHvE1vSAbGs/ua9gCmJTeJVvN6HHv+lMVuqEeYEcrBQUKaDXGlISA4wGEuB7
aKJpAJmFwOIxBAC1Qhrkp09caCz4dqKYtNRWvKeOyY8ENdr4K4NJQZxGYH/rDVtc
sjcGlKO+u/mFEDVuz0nwVriPC0QtqC0ALwhCEZLgZGmhjpvP8AQN9aNqHB2K4/4s
VSEQpvdo3bRmM5eINXFvywpapH5veP8QYY5O0q/65SpDHHJD9tVGiOB0oQhMMD9l
03NyHqAoPnJZNQsYg6p3NUfXor0YtL3QP+YkjQ8MBldeYj4MkPa2bmPHk1/KFtPy
1euo469CuNpc1AYZxMUOfHbPkhWH7f+zY28NFJn6Bx4e3WHS6sq2NAiFJH04mDn4
3c9v5TmDrknFPXSxApVHSUDKa97daqnjdyhC8MfZwUvjsJ/YrCox8qo5Yx38UJgk
sps0x/1ZZgaOFT1Wkmkx3npt38AUjjbv1kfSZSHA/xQPdelVYf/FpcxQ1n8MWNPF
rx0fwzYxD2ehrdDE4FKA2KciO7dLVxDkIESV33xsdctDa38UGRYizk3O++zpc0CP
wRtSD8BtFKU6XA1Oqx/sl844wonT9P1pdT4UjzCIRNV+5DFJ86AARAnXQpUPGr0t
JmQ9gX2NgDFS8LTyxaPrUV0rdL8zQ981POCwAB+LaOrKB/JWu+lpP/1ORj2tVc/k
1LhbiT574vKcFzlfu4Unab66gsdaFWNSDV9DSymewnbap7X5g4H1OlpbQMnwMW/8
0Z84CJO/UllfEsfKwyskwSQSsJ2O+ju5aUp+ROJqxaecZhhaDU2nk5YEqTBByw4S
F9/lJYKeK0QHkI/aWZMT6Qf/bIJf32CgkbC0BZ3gCacfqI9z4epr7oXk3Bf5EZSx
Ee6Lo7GyDdZHzNnJxGbh/5c3RJ5h74k74kFiZC9QlPNjnXZK7dwef5UCVRBH4k2h
ZV/Zc9clkT1oJFZMt6wf2DK4BKshet62we1dq9lt2x2f3an3EoSamqitmWgylGxB
oedgK41uSfgXxoDISG7+H5owl2HsLjEWKgg+GBpVfuxUBSDjc0zVeIFF5juro1MR
ReonM8zhBfKb6Y3C4SxRxKErFJmtAuVd3bIQWc0fGqVDgSTTBfzXpcZdHatrBTTq
RNRZOLigfOVK+9SmsduqM2zum1T8KiWTzyESHkijK0C5x/MSo3P+M2cdj9Al5kiK
q7RWAo+k5fbj84/l9hL7mFDj4bgpnPPI3tLvf3P2+W1OIK3TTaFi7hVLLjkMmC3P
hgpg33cihyyWMw1FYWbk8q2FNnqAU6UjXxVbYOiJyw8aN5WSsvsLCC/6nlAqxMQ/
FkWV/aPKJDxbiGqakbtRxtyDbIUVHqSSsqVQBrFLkUTyqrYzlxOLP14xyK8XTOoE
UwJIrwRxADMWOFKcH7VKZPE5URLDoiqyh4uD7gDjBvtxBagypQk9fJuEQ+S6zTJP
SDfBlrmpL3cgWmn/xFDG0XCad4GRRlLGgJiF+LdV0kSevoAkNfY/vkbaDdvXo1cl
tyBaYseZe9hEg6v4i1ZtHg6ISv5YyrHkAvVhsr4SopkBMwcbz44EKnPe/oARPbT0
qhwlURedymM2lKxXLG0wV35IEUoMqOVf/Bd1BlIkQlJQT3PnUTV1qUnNDG8incFy
WdUe41WajaGc2SIk3qF8T3NOXMt3iAl3HVUo7gGD2RTYYZyUMdgcYy134zk2Mry0
N+7zxNSkj1N4CPHtp9n1D02OOl3nViY+/VgNB+1LMJl8SDlPw1P/ZZF6IiCHin4T
8Le4y/mpsgB64w6LGbiRWOn+QUZdM9+ove7+aTSnPnf1qRYxRApLjks8jvO9zcEA
HhRSjQvQjODFHgMUU1/jvq5UUXeSOZUdmA8zXufc+cYqvgCYiGdP0QGcASIisn7k
rIDO0kjEdf5YH+Lw9GhM1a2qUh2zW2G0PecCfKLGQ99S646zT1hQy7kXfJyObDVD
JsT4uCQsRAIEvDI4jRw13KYWY0Kg5Bexrr2WlQ7/47zqbLUwgQTPtvSmMOEuWAq9
yiNnL0qzmveXDW8bQKqsbtOSrwdyYfTDCklpBgGUa73yevx/Qcqh8dacSmxL0Yf0
iM9yfjZjZTldsTl09lzqOIgNBF2PzY1v5Fbg9aLcoGsyWnYLnPseoxyovF3s2KUn
qAPU7RkHfQgr2CugrG2Vdxjmf6w0PawrzLZRG5VGrvGAcDB+4kLAfOxA5pntB/rA
4iJR01YLFcxhzOAnhDWWv5j1dfEwiU31Oww7xBNr1WpYs3PlkFIMuXeIM+dgNvZ2
sR4L0lJRpBv31hG1c9dbP6V9pHLoN2Pnt9Js2oeyqKBsbAp3xBIJUgVVGb6d7MKT
8VF7rLxfsfdvHBDllTl8brk7UEqvGoUh6ut23KT3TsCnheO+gPvXN2MIN8U2WzJH
5kT59aatcYkTNj2nzDy812oX8QoDXBuEr9+uMAdtIzXXttM9xzAPLEpBONgDxPWy
L/S1pDeeDZe41NVQvDKwPLJNny5/a2fxm6K46QsAWmTJAPFGRT9x2Q6QTfo51Zg/
WrjTfRdVUgB60OA069H0c0LqPrbnC/ng0LnISS+U3S0nR0WCRxtCAKhrUt+4I4PC
OaHy8zEyGPxznyIfoba6GtKn1qMhoMFTNY8kcj7GDbgKuUDu21JZLp2CtDt9WW/r
oA3vaTbWfmg+i39FdXg3ftyrnCCPmIQXp2xlx9np+8+K3hNhXDpeOdlXdVc/ho4g
bPP/qdVcqIsZdlNwBgAYNxN3QZlZCzfkHoPPQaqal/CtR+dUOC4/46p1PnVjON8M
9b75K/yynfxA2MsfYZCCBFJ+TZPD521buJLskczVj3qrQaTan/HscJgkcnB4Z91U
3JotN/hdtlLDJ89Cq1ScO3H+E44lW+WEPtwPbfiGgF3tb/Xzz4JuD/0tK/zH5HuB
AT870R5LJwbo0sbtuxKPrbQEvoUSzgCz5J6Izi/u+u5Kh/TOakpgmBxPCOKvqG1s
GHHOSATc6+O4nTf5G7rw6z+1lBx/noy2maMr3tQqWyLexezZqbCiMiQsBYTU4XBk
k9noQV2ZuUJooJ8ZKyuaHbhxLy2rkNPjd2ADeRogSZ7wrNPiQO/yW7LhvrULHIFT
jT6w/Pdx4VGeUv9wovmQ8XtlP03wcVEz5SzqGms6xhpfz6/Qf7zxh8onBVKvobpm
nWoODgF/g9qOx7IY+ZI9+h1UzK9j4un9vnkqjaH7iQ7FoA+qT5eVsV+Wcirwunli
umPVLF7SXf759cOlNVFh417WLLiXVipmw0DZVoqMUD1SsyxCS//m/VcZUkY4Srd1
GS4HWJ6b3afNCXO6zjl0ZkjiDifduA/0N9ihKUuncNPdtgYMMhlJReGp9NnhezG7
FPZQO2YQrwXCh7TsTQBsqVk0uNgDThIYWHOMUc3HAWT1gQ8e70+RFB2dJCrCPY2w
uCL2j7J9hw75KnFSJfw2O4wLpw/f2c3p3JiQMiscTizKcfhHLRcrUakJA0k02ixk
6Ke8W9tvE8fe7N6AZg8wP/hJJonyB6zuANatbOodMQCGjO1bMeqiSOAaz3Mxymc/
Ui+Q7s0+45AeCdbynko4qOdI75EFhByVplDNKa1NofZZrSvyl8Da7q2q4EXJ+LZE
9RTrUhZ+2rt5MjKaqjzILPE5p5BkNZilw14PM1MrtmhqVU0Kc7yrfOzVNIost6bn
dcRrxb5Fw/SOFc8rIaGhq4qDVGNdt5vlXhFDTK6oe0qQy9Zgiu+qR9a6CH3XKFc/
XCKRnIhlKD+lo4kgZl3tU4LbG8dPj9KUQ8BpEYhm4FK6w2x/15D7X5Q+HcTTxrqd
CuH2MaOw/Uyq5cdLw+RLMIeh8Zo/XdI6iZJiJTZyR3Ytt1gqYqogWoF0mRZ5dFHn
gcQhQORNFUsGkNO2RJqhSvaF1Tl8wSpeIjJwqBVlnk55SfdzDGCsnCIdVJX/cHLP
OmtWmaB1qcTuScYV49FjU8t9m4zQYgfz4qwR8lM+2uiAP7v9by1n31Wkg7UCHYFu
AA1BmpRqvGdONnt0KW+oo53R/xzz0hN8Quaoq1XM2Qws/JFLV9uaCGyaHwlMXg2h
e6RW2tf4OUC3pTnGEObll2ZspO+M8UUhM+l+nJ44TiVAxQlVZQrB3jzK3Gx3aTUd
ZlUCTT6kEurxrbukwzeR/38A/zxgXielAKMEoZHfpn1UTKwwT+rmvNij8Jm+zl6s
jx1EZRPMxYO/noeTTeRMA6/2+NW4T0cpfG+I/NagxTMIHW1ms4AGKP1VUKRt8e+k
PNOCLMDA526iDMF8tlkE8Y8HaErJH3vR4+BrAgVqENj52zHbxxGeQE64K7mh5X5c
/RrK4LELgreL161VhAPSQ4HL01RzAMnKZHisx2L1SUq0EqyrKKLNvp08N40CY68L
sFyLyIFVWtmhs0rqgHNoMo3HOsEuiKpMjnHNKsbRCnHfXujTkGNR0IYgjdHG5t9+
VgmGB/bwLEJT2ZNjGbDdvMsui77Quh+1oLyHxr83cZddyUGCnx6Ersf0uGsc8WQf
RRVov9ahXwx0xciTrK2s9xi2zVTVHCrmwV+AgrSOIblFJb0L0zTPG0U1ALlXjl3f
47UqSZX9Uk52em0Vqclo6k847UTqsjz5nLit//9Pl6U1Uo3XfA0GwHoEXMc5L5K9
zQWMG5hsZIy1Hpk8sIWnKEoV0YnHERn9ild0BvfVRyMP02vQqf0x7vuOFExR4t/t
V8aOlpLCyd5Rrsoy4bOB7v6i90ZA5k9CKDIp5Dtc7o7eGsK/+w9WS6BKq1Ef9InK
UAuNp/hnlIwzNLZWL5GtFSx5tDoBQdyBCyi7xPq9pKTyQc1c/SazssftjENNruMH
liSMHWLPNE/X1gSwQMaFWptcWmKIiI25IH4wKo8qoFWwCBMo6luTbhZ7E7zYq9El
R8ecixLh1eFufJLggvzJsj/QbZtMqnBQ4xAliueZubK7YfSqFnj9yY54INXoSdps
dZjRo4E40qRcjbxDdE9Q48EIsk8Dm6dbyIjdHqYnJ3bmkuVggs3K6Q62AcSr/4b6
wnokDwFcKvz34HAPLuom4VPQNiu0Iul7fwBUkfS8Cf8NKgdmi/I6SvT1e0H1VFas
5bY2ZEUG+deV3RUlu5pKEg/MRZq6IwUdYlyWw3/Aoyg0kIOOReDiLsVt+V59EgPS
ql2Ivrw/J3BROLZoywKdKnBMSb4uh0bCgSFJI4XtviKJlGfvdjV4KvrjGN0L6mqw
AMAdbC1G7Ch7NmmF32vvvdX0tG6CHnB6NMonxRJiElmO7Qw4AY1rjUFgr8wUlGDx
89WJKXO3uiOd/0tU5784qF8WYm3wR0Oo9C09jbM25U4wryZneFAc9ZHRDtkku5AU
MiyT1AQi768y0lBFZL/ixce0OmROwuiFizwGSdu56VZwGQ/y2T82fGmt8eM15Cg2
9XN1CGdvnR1q+o3tlK7YkNSiLlKcR02ux2v5Gm569VwBRtWnAphmtCMFamUTxF8c
lqyHUiHKcMY9o6BK9hCPRee2Hh+8ypE4KwxA97ns1VZrmfi7cRyD4zDmTfpMYJ+D
5KveSFIgAU8CHIk17IdwyOhYbD9ZqQcoApHQVSR0CSMnM2ZVZUfWOfxCQa/lyXJE
0vBjXo8bVm5/5LAw9oMxjX0kOQFvJV/I+ar+mJo6Qt7AK0vJxEbfT6B7jwfOtIyx
wSxbV9uy2JkWY30KsbrbL+xe9yw1s4Ar6F5d9quf9O4BB5F1OJyzgH4aaPHq1rP2
gUU59QZ98JpU7iq8eaiDpAeiHMFULPVdcYZA8Xl0C4Q60DgV+g40C60+Gu/iiuGd
l10bjjcldJ9VM869FoLn1K4wehR2OR7fxpFVEm3Re2Nf6kB1J/8OGFrGfECM/iKQ
X1XgdjykB2eD/E5ws5SUVXE/aKiZUiKT8YajnKzIK+irZsn6AcvUbP/PeRh5UwB9
BQ+DRsY8E4BOBV3zNS4Hhl0weIlE3iq8R7x/4rm4j2awIRtJaQwWllsgo3uJYMUC
TGU4PiNaU6ZrNP4gkTU3JfgVYOq8RtyMgsITWhga/xjPJhlHzzZwY0U7oxtHju5E
wTV8bUY5GiBD/Esrurqlwf12maahs1f7BA3usbkuk8YlH0aTWPN+KDQ0FnK+5wS/
16cEUHhwJrhMub0/V2yUnp6aah9OsavgV/auk2reyk8TCXEQG3w5LqnggQej43Kv
y9mKCqDA9rC/obieQxxBwPQ6+GQkSLjVHgnhYTVb0R78UzwHErTfOOgP/5BSeaxR
HKf5hjX3sHC9aimOd+iKO16xX5iAl15z7kjZLl7RpkpHFgJQWZQVvy6fYKUPhHEF
L/giiEIVuArc/Q76vHtHvl6FUiV4qgA9DD0X2F6EvOUnS4jlI/pdEg4Xd7iiHIaP
gq/CFjiH4EPx8aO/OphQDPvWiDU6zXhbMvc+sKeK1SdzT7SoTbCsbd5PDB6f2a/c
5sZbWtPRp9gXGyOn1hxDYtmsFS9/gjgcAk+DhFxqHF4gPNCmGAma1kx+J2B+h5jP
YrqmqiRezSNgiDDY5CcQ1lQmRro78gXmBYBdrnwaIUapja1ynSDAX349Hy6cCb9L
SiboVhVuL8X/JDNQ+fabf6Mqp40dBXP7bELUfXJHTW2yF2MgpGnYkb+jm0CUCOEI
fWBl31qroG3wWkor/DZRxYnaZ1AR1WMIFiPig7Rj7XQ0CkorVIngaxfwNYqe3sF4
4wO5gptenT5d3pJZPBEzPR3+9hLUJHl2G8bVl7wTdud2r3NMoHSK2ka0wZCMEJAO
7wfxpvIkKnIBffw8dHZhgXydAoovq/3BfIsXuWCWnwyRRrtLi79s2zzayqpR4e9v
lIeLfV6ErF6PnwWgcyv34QVprZLUOtsuaAuMwmKj8T/Ng58i+6pgswIQG+OTmHho
gtu7h3RZXQMD+NdPP8JBsV9WVs0Eo0v7A+12ighlQjWO8nkUmvTELDi2t7MiBHcu
QZQ9JVmxDL7jj1X6Jq0ebjLOnarIKSiOepuqD5aICj1GwJhLg+5ygEjR434ABo1U
eFm1ozrgxKXbFZFhRKWdi8qaN5yftdbsW/OPX9pWI0WOQ+FFu+CCxbLL/GCWNKzd
Csqf9LST2hanQCUfxjOZMqlehRXPEhXfsaLkTJiDno5sP2ERWVCqzLKTQWI3IuDO
+v8VNFdx/KbZvFs806+MzaLoA/KsB0+ZvewWLVchYIfP+eF6BhRNDPX4a+F/sOpj
huo189Kwv6AMetvRU7RYUGAASByXZPX5WEGggz2dqSW2/XvprttXMPEMq/H/2qFh
VWCxsSvxCiR3b9TZ+Gzow+F98H9VWkm38Z/OkYNI/DndGmx9dK7xZC/oOcglT39I
PcSoX/WB0KHhyzUSaazddczeF50RO+826cXK4j8bhUkmdQxDK9ZKokOIvABs35Rg
f09ZzSsHClcR6mZPIR5pZDB1P4qnRjVH1sE7NQt4x/jAq1qrTSHWcgOvUOVgjapv
iiaMT6WXHE/ZfxmXnx9XZoIiSHsB/2KR77qvOSgx+B8dF9w+f9j0Qoejy/LqUMtZ
+pgx4IZZY2WHad+H5GwabIg4UjknKYg2DO8fWeKWRaPUn9IDc0OC5AmsAipRQu6h
DHg6n6Mmj1iMS7J6bivwWym5TW9B3V9VPbrRCz67Xzy3zCPbZSjXT4YQgrFvzKt4
j/zwcns1GarH7Q3j+5msQQ8S03IsI0y9r8B2D1MqefPCa20Vdn+EHGlidqsnaCDo
yqKgQu4B7vgbolFBaRld3atbhlKUIN80MhZXkZqQViZGnzA9PklQz+VnQO5YwW4H
H+MumTACXXIJCmgRZo5L7VMKM+muKh0JVjGg8eqSAR0GyeLvXiAZPYex9xhznKd/
ISGemeSQJQPb2R+fSOU3q0HA/aOspErMrYEY9CBkSM810gLNi8uvGB423XCVL6Zc
/sINrUvL/WyoEchvB5i+G7b6TLi3O+Qy6DPZtFowf+4yj9zF0x7Qzkx6ZMa35pmB
FpoUNO5jbgAawQ9EqNOrM2mX/xYAE7axr0EmAo/MSVZyFZiPujOKvfZ4j38ygQIr
kPrRHnwHegt8zgPWSMaVlGNJNu1VSKSG4WWNGrynX9fV2Sp5bywI106ZNUNm3QI3
Zo7Qfsn8msiLXjCKB13IoqwCgsB08cebtr/08w6jZ5BLPN1Tb/V/aVTT37ElTDkt
Xw2mHuZ4ZAjaRuydS64gFtaTbYpCaOY8vLYB+ufchc/jsCjwSyR9lWnkXIN+1D9D
D7Xs3/Gaz2DWgncmhtxQxmcv2g7P+QEaTOttvqlqNy58piAeDytsPsfxMWhQZgvj
v8qlH7KhboHSVPk7qDdA8wpxNzOAxlymWpsa5UETXa/D2XL2C1pAcCMd+WPaf/I9
zf8v5SU+DW+sSskFQOKHNHXexwmNREzCglNipdzJqFQWU1Xt38zcTh/N+09cIzal
gyZeuZUFvFMzRC+1YexGSKXDvZu6ZlY29RJAhW9CrAtveq04sGT2IzdUky4r059D
zfYxom0mSku6prISke6FA6qNGBnNNCKhVQ4I20zhstaUvNNxorUlfeDAsayYXwY6
NP77Bs7kvOQesaypI4blRLH7GJ50bZ71EqLVObGQKynQLEO77nN9WPgq53GYzKEs
3ieVwnOqYQ4VCo6ta5xClrkcfXkNfyydrylD+3rdmZwiwZa9kz4adfYNWPt3gLIm
B2uBn+43e7FuXS6donBolGP7aRltW2hduHjFc4U2PMwDY0GWeuPAFPf3/X2NF40m
ItIH778tFhQSTKOzYZCol8e253vQEfy4UNbOjj06/KbhEC93hRIqRtcMVvcpX2tn
/Uaa+cGkiw7Npdyjbmy8Lk/Dh5GBZf9mfDTxUFe2ZMVRIRTp2QOenN5UO8RKd/Q6
jU2Y+vhVW6oaJqr5r6QYyke/Nk9v3ncQDaPVCEgxLlliRaULmiznMLfrph+snbOn
ml8DMDS6pnS0QUMej29h/lIZTGXFiMjB0OAjWlEVWBxR0Q90g69mQgdBUeClKnGw
MwGAysyvWmnOUPwQPdLMoEPw49yVltrr7BfIfYk0hKlBHW4+Zi3RnqAtBMXcuMwD
C4Zu6kelsH2GdqixHKSLm+lRQHC7MrxBqqkU0JK2vBU8IcZ+05uMmynTQsTxaklh
LMz0iqdn6mkG1TxgBklWNOrdRr0h2PRkZU+VHhdSs02XhkQvF+4R0MxjkR90UhO5
HgbtzustaYb2cHqDl6tLijrViExIeoABonCK/D1J2dyvNy5iIyYDrMk6uQlL2x6A
opr5B/tgqcWKi0EScbFBM/kA7i6TJBqrRLlpT+zC5w94G/Ckmu1QutLdATk1Y8Qm
kmfLVTUkLJVAlPzKjizdEBCfl1arfMOijsSF6wgCB9Il+TMrlVXLKwx3osukZQX3
kk3j7a4Frhp5T88l8Jgn+XVYnQmBhY+9b6heT89Xo/OalxGv2ux2oMRclEvMl/9Y
uveXCwxg3Qyyyb57FKRSoobXSs2tDHClVKt5Wx7oIekkJgmfqIQDcvqfM14xbjuH
BgVnAQg3Z1YT47pulFn6smUpznLGR+WKwHMfUcUF8bOY+d+tb/VKh5iLIM0u6/EL
AEpGfBCaWIgpBizS0GTosnZcXM/Bfgsuz0OTAKj3Ig9YV+Iwl3a0SonRaZDZ0bh+
JusfoAZh/rD09+iYW+uMPFbNQUiRr8fZwZzSzpClTa4uKLFyoGxk/OZT4L/tHACW
a75AQ9VDhlrBF3edFG1ihjwjWNiDSHORgjHw+c90qhiFRStKJAfl9R00bkPjKAyp
ZUW/pKwWQfgxRLXwjVHF/aR5ctkcRISPb2vQlxUN75j4YlDSvatZuXj1U+fmYLpX
ufCebmxIAEN3F1ai3kj284bLABy7bBZhyyzKaLY4VsY+JOrsdNuPgoBp1od71hrI
p67ky88ZJyIL5A+ElQLgUNqMPOBwIi8MotRWMfNTJUaTuhtrNt27C0clb7QZm6Lm
5cRvezGpUrkw2l4/kezxMRYL+AkEXcu19tSJU351eVPdqgr9ZCYaUPNoVExXs1xz
/2Il+82lfZWfApcodRNmj57kq+RGNXl5RUqebf4yHbINmzuiNyofyXxq/c3HMIjJ
vivGxM3g8j979yORIqYG3vMZyvFVAey5J7FgTi/TwIr+QlK1iFLSeE4OWTJTen0V
evIgNH7A0IrhX3JT6UQ/l9HJk6xwgURowOZAFSPBQ4ZyJ1ktyJGoqPiFJ9eLXGwI
mpJd/bajb5z1EZZMSLLAmJhaks0ycT4mQ/IuUsQiMMzDgcpiQWGIYH1u3KZxSShe
bDyzl6l2w4K/pQZ8jIawdJ9HxWfdDEPx2AsFK3AQXQbrSNSzCAHMm0gKltsousQa
WZUlmxFx4ASRrt+Sy/agaVLxQA4kD6h0wbnD2WcU7xfBS5iqsCX8VqH7Bj0HMzN3
gFlG6Mkk0Lat5vtQHj/3l391F2AsLCVcBCy/qbpwMmxTZozuCJcxezUvlRbgvegx
Gl8aSF2mVBC/0khTQbtu2ySX9talrPGXqPw6N4k6rIW+rVZP9EfnJ3lN0r6gZH56
XVjrRFgWoF7dJBE6ry0u7EOIgaGQtnS4F8r6KqS7GNvLbvf1SEzac2tlT/mjaemJ
yojI4IK39fRBQ9+Dc5jkqjHaK6CQ2oZm1BovGP25+0vC1/QClPTJ/mYxppwjPnWD
ybJ4oOdZt/g5jGYyTvBzk3UjsnHvdKqhSvSjaYDX3my3yJIgDgBLCjtw3oBVRcd6
iwQIGYmwdatJH4FphNQ7B6GVceFja2VMnbd1Kww3ri4DRe1mV0LBhcxwd20s46s2
0F6Zew6bz/ExpZBp2jXK3BVjXZj7gxlWX0O0sAecXgmYhcb5hSJG2U7uJPgYr8X8
yh0oyHFFrCKxAyXLWAdm9FDweMnBDYOLwasyp5r4oWjE8zRfQqzOpI8lZMwdJDn/
s2MVEUxb7J6CEZWSgiDaVasPxgOtrG2+Ab/JxJrhcI+4mkPc7KQceQ25NpWfPZaN
yjVWBC+EkhnaFufS6ZHQC9AyeTYOsLpVNFlna5M8d/H++dRJvl9j5glBY+nu2nwD
qE4ThdH65BshGwq1KOFP8kb54MGrnFvGrWRhlMuNFYu0BbXq4KmugSVPojqfHS5o
ezhS5tFBRkbw7eaXyKxYFr2tbQI+4QZ5LvzqQK9QPStBArHQ1ndTA5ezQ4+9nH24
p15awKLSBf3zIl+p1GOcq2W/ZtWlH30Suz4AMn49I9BsYTo3xNuDFrLRLT+Mjdh4
VHZE+AmtMBz1TS7920BLHsJWSmIsc1cdq47ePaCRsB5RnXvd6Ul37hemDR4o5hVK
2g6tRv+enKz5o4p3MgpaNC6a0YfIpDTLjHbFfCCUZrHCRYeOKBSNAywz7zdBWSsg
h1RKCOBjNgJKkdLgIh5HfnE0ankp4qN0TryDBa6YBV8hTJKgmH2R1MvDjJIBq7+s
mfc84cgJdbJKPr7T7Ujn2bWH2Y5hbebHoOwd1UiLMiiTpHbMQQLxGj94BRq9MbMB
B8s4Ztho+b0QCklbAFB11MU07q0R/Rm6LvwF8J3tZH4FBpWxGZ4U6XxElGmWg/jI
DDKr/bdkHvdEE8qpszwuI9yjce8Od6tfLb08Im2kE9NU2TTA3PWSTMD7FAShBWRL
1YhCXh8Wwqid24pawEYqQiRZhY4CFVlHTE3qZsWulMLNdqj5D1wLFi9Pwrv2cNdR
jn2Wkr4BbgaOFcU+MhopZfeb4KgN36s36373BmrJ+v0DB8wTBRin1z+r8x7g9Kfj
YQc18jHOgx1v+A/804aCv1I9wNJMD2lgAKBOTA47iSesQ2vERSw7cVHIAWgAni6c
NPeu7F7qr2HqQI1Tpr+aU6QgAlxLeUjF3pTAKNf7e7tiTJAGP4F8MGlFStt6TStQ
Dx3jAWa2ZuIAbu8txfNJ/EhTvBmmF0ZLDPNw+iX2mReatLey0jqX06YYrQnVdFwK
XeT/HsC3lqk+ViWJYuWlwDAT3fj4DapQVr2nXpwr5lL4/RTnH1UM9dszHrogji7Y
JQvgI1kKzvckkgDWEJXuXTE5noWwbDyvJu+gjWAzvoAtYfSHaFJZ6fdB6iq1K8i8
ETJOeDsfwoZKyZaG3+xzxFWScH0SK2Ae/OX2lQEI1PC9fc+xDkx5gEjcWJxvMoVO
NQAWj+S8SDir7Tfnu0rznrKYo0UbHxQAyPicHtRYPKYtzsQjsuu0L3LJ0NW3uAR8
DT3y4GvtMO6eSZWnHvaVXw3gd/hlS2ZHoV/pECB9Z7ib3KkS4k0mY3Oh628ShS0C
B5MaZ44y6R0jJR0N0EdebpdwfSItEf3cBmNCtRaZK7hND1nABkcAM9wejSJzG69h
5YOS4Jz0xl4c/sdP8MZYacfRp4AJAOJhloRX7WBMUyc5vrsFMNjiDR9DpvJLxmYw
fGgVKIsnEmIFxJcL2FWUM3kDx41jT9vcfjexpOd9fEOYBXuLeZGavIqSY+90KVIr
f/jdnq5PWDmEQawwZemQDYSYE6mkMmrLWep0uXFqHKaj/INucB9zIp/Z1c0yRARx
uMf+xCcrleNTuYQmzzpEPQ8HZjJxUn9E9ZyGPgPnvZzVQJzULCelY855Qbn6mRYW
usYakWpId+2fvgSYI2BpOdwj7DaRNsscvqVeyesDCraZxX0zoWtjEQZrMMw7FyGn
PFJp1cVd7dUyrdJsk+T38KxWnAUV9vbIlS+zvvMbA1ByDFJg0ULPJAjgoJaUNNst
95BjExFt1IeXIbAoFnSJvdx4/TvQiQ/BTbO5gvyb+AUkZ1HeXtmon9E0C78+0b0L
RpTiDhbxXXI+u8ywQCpMHt8YSFOUBjk1ytH27Y/ug+fk/1FrbcieekhSyma+SW94
z58WXNionmpUriYu6Phe05Zp96qhaE3fcI88Pg8j7VClvDb8Hgo+wVT0JFVJ3GFh
QPeVBNqOJBTkCcfp6noy7/Iz0HNl10s0XzargS+gQHTqT20B4aUdwingdXXfpGRW
QvR5U4jracQ6PbW/9S/U50UkMvy8ccRgALsTFY+BTkBy57TnzXRNKIvnVFFu9G8A
g6KaPfoSCwWaImwhGaekIvX7qgoApiNJw1Oprf5M6UEjaHjXLySt1box0W5ArODU
X06BiwQLofKUxNltn0nBjhuWUlm/DJWBUoBhrHDLQDkYh9+VE7TH6bs/HzuDExH9
2fcojXf6GZIpICD4LknJ5cEjPWeHxycIFwIVDx7ql13xqugaPwZVnLA0woF5gEve
zB45Q7vwVJ3zq14FTFwrMmEl0L910M63vufBj3fMATQFeqzT4mdjE4xUvbQ6MVss
m16jgijceemRnO5fEz1vBu0IUCD+x7444PDJOIK+29rH/gfapezij2AIYFrjTWZ7
K+TQhb9zFvf9E7XfZnyxSCtON3W20QVHoV0y0kJirC5NdmTkZMb1chevydKwc24H
l5GFQHV2uiLxtmkEL9b25my2LSv7YA74MKEyKkNe+yWTLTwsHiEJy1yBNTY2sjcE
AnG9oI7xFDiDoFs/D+A4+1O/eIqvnijTP4+LclDKkcikV4NZP7s32nmP/m7KjVPa
EMznj78ZU5TkoYfF57OIc+4HHVnisYL2QJDppPzPGA9cjOoNgeR9b6/kGlkvFi3V
YXSqAVAmnUzgaggIqnNrqHguxiJHNliVaOluwtTqbjET3NtyQc6zZL8MWwRVrHIH
NIb69Q1eL9ssCvzlqhDp+VLp2OVyr51c0vUWMsGKzC25FQZzSByC9H68pucorTUR
PtJFulTPfLUF5rYSYiyLaOuwE8Dqn2XvhcO6CvNmOTsEqXEd3/I5HUTJniYSEOvK
ptj7ohmXxpajKnMqHWgEC3RHzJC1LMnjuzGTlaJdYy78a0e49XDBrqvngMugFqO+
xj9s5ZmgeKVTUwg60Kn4IUKLvAL7URcfHTkG97gqct8TZXhvx7xZ0vY3t6v9Meoc
3bmkKmOt09BMm/heDeywaTrACC3h0drJflwchSaYNMVwMzLdRCWqfrmoDOgKdD8z
SuRGIsMKaYB6o+zRo064Na02hczDSUAoqz1xB/sv6sjxHQqVB2081o0uMSXqfTMT
1c9nzlTtOrqLMBAxZKu2cVMWHpds4o3s195t5PgjBuXGlItcZNGImxSA5R9IzFq+
zNw4GKcnlOqebV8tcAgQWvsgDJ2jEhtGPfz+ZrcCaavbyxAwVdGQYH215pcFyfg4
u6XmoR00LkX8862eyLxmZBrMBADHZSk1IJttKmATFT4JPDF6IW7/u4sqpwzlhKEM
x1An/F1YVRSez4JK4nKIgMmdrfxd9TaiWwCc1ZU0nTBk2GMAP5gUMx4oDiBDml3+
UQyUYSKdpaK+eA64pgsXgQwUT12/ZnpLmJs99DujGNNtOXcEDMQNXWP6/Wb7CH8Z
mSNHCrsV9G/vyqBBNsOT+57AY/X2t5Z8qyuJ1002Y3/uWYsME7COzK0LiH/e8ca6
R9ATShl34wp9Y47+ipInNLApe8aW7w9RwRq7C1N4Q8aHlLZctj64BqSirg/f1vqE
5vy/Mj08UpITlnwrYWsr9iy90hPLHmj6SMP5nSdWhTvWhnYfYHEdCeiUgYSLNhD4
zsU2+Ul/PiYwN6etEEq9Af6+aEHHXUrQKVUr8lRL4CTzSr/wi8BQbpNT+wsIHv7Q
2NSZ6ruzvgpaBHYfjtSyi9al3fwIVcD7vMwg+n+IcSS83UfUqYSb0x4DSIO77y6t
lEN+MOdPymf+2MIvu5xmsx2tDkL1Z1xAevx8ZunMuWu/hWsjWPa9E92LBrmSzac0
3rKgqjlyR6bayTT/ABaHfqRXkRP7cdMvIO1p4TkpBJA9FptA1Dy3KxnQf/vrBe4L
cTKwjeKQN3Kdsr1+URSnkRM0cEXKhzoUZM1a1pZ0Mal5xzhVOHHvCOJvg8IYgMCN
F78+AK4KlHV134GY2kYhU406Q+TJ4q4IIQKx24QEMiO8Aa+6HFva7wO9XvFa0GH2
q5oMZb0kGRQWk/PwpiuAugdDM4fhh8DVRUrShAmJ/9EG7EmgTYwiwLFXZvtHImgC
4deHc161M/OqnzBigGSAwSGqI1MMpxHwmd7jhuuWU6p5kjtvf8bjecKek3lpmADA
44J/yOubH3q5SZikdgqxQG8ajhBnlD7ZScnVq30QlQ8RfjIjg66HEi3974ieI+Pk
eB+dFoOv4MmqJGNoSP7DRzednMJApL0FC9y7F77Zu/ue7yujp0AD8IIxzxvVtXz9
kXQJWQRidQixJHIikJvNCPh3b32JcLWF14rJ6Nr3fDpvVTsm5XgzwSAmDKX34IHw
XWW9ch+v+RPRP3VgPv/2fXju1htFMIWDhVVaGHHUTPAGV85KNpYSTgsHpTK/IorU
tY8ZGw1Fmvsb7PqEcuoV891kpGwUfBekLDxybwszx2zVAFH+xHGJlrgRsiqxAECs
JH2SYf1YfaISdpraulRfFHpg1uKadrlC05p6ZJTXsl3oOKI2nhxn+I9TMJ6zkuMv
WY2xfuP81ddlqDhGJS4+hhibY4JETL+uYNlZctswSjE03nHkYv9BmbhYqWfkW05Y
S886fdvZTI7OrzEnGF0Vq3KElZ9lbseCxB8yCG2/CV7yT+NrsRknEWe/tPHjFRRj
kozaLN7lYnd8/0QFSXMtP32MD8uL/JZMsEHZs7uafPYxlnns8qXsTKtq80vjVNdp
cvqU+4XpNToqlDxSBmoBdir80b1uW2xeeeIcKsDUw843MTUWNw3/2hU9u6IjkJMM
keoZHMsR80LeftWPvPhY3vwDiT9RRHwx0VQ5f4g+pU424I02L+6eOIje4edtmC7X
0nD+NoQCxee23oAevGdGk6N6db1nCg3cSOYyFH65eHPeJWwPnmVbh1RYiQcLpJ7R
VFE1GyDSiDggWDIGKZuffl/7dN7Wt2L4PYvUuy7lAO9YlWvJMNKy0vqZKtzYt5Sp
6cLysHb4JSrnlB4NsBXr2l1/QJvmBeJR8zPkRRrZDVLwNi/PHz20BgSVhr0uGVCg
cAzp1WH4awSe7h4Aac1OXByS+ipZLIMr9RyMOmKAScdf4t3BPO1dLEOWzm3RD3R/
1ruMzrFlt5ykyrBPe5WttI6m6muk95V9i7XVSzCvuVb7pXqUyMCFiixlj3EpmoSh
TvWYMazVzebYgIXf4QLvBRiDGhhVcCgH0/c+rLrMO3o1TWu3euVjdzVejzmMk+1f
pCcK1Byst6KYkkobLiWTd9txVGe0DS7r9PFuWDwcdF3gE6BTtKZDRldHI4q6L+BF
z8UK9ywMoKtL/J/4ajE6G31nywovCMMbhX3ksu8YIo1x8/G23od/4Ks0uRTeVj9q
KAnzBgV4z4IYZlOSq4NDGtF4vKrz0BOpe7FDigcZpwsV0DvwHHordS/gPHOm8o9G
2N7OVgyLO7Jh9voZqa4VNPNpWp2DvomgLGTU1f8i/fW7/sBd5yu0vHUblwpRXi5q
WViP5F++fd8yJMLtEEF8g2exT5MeV5iQq+Zs+ck8gWjImCPZaQURZIZuqotZpI7F
w3qPMzNXLZuWdvhpS/WyFfhIHoDSVihxT42ouFs2kkA1SAxTUci9l2X0kf828t+z
Xr40JIPjbzACEtEkcXMdwx7Ob5EwdStaJR9bgXbSb3RVRIKjYbOBb23QLBqlzYfP
/jGpy7tuCmHiys9ofweQpkiy2wDzCulHkd3C4Urce8WUfwTtYZXtQiRhMklLt0b7
KyVNwwyl3AnwKZmtC31PVKqIztRg6S2O+w/oKX2gxReTApGqNAyq15mIR3ZPNGG+
lPRKtpGT1SUnYexcYAEoFsL6pTgltdeYtOdiYNOvxKsouZIFp3hCz/gzCoZM278S
K45erIy5w7kQa84LWEVOhB67l1yZ8kUfy2IIqyzU6RW77XNpvD4Z45XR20CgauV8
dRqzGDHk9GHpu6Het4JcPCFbGmWxSmqYlDVxd6FH6YmrNiDUqN1ssbTbTMEHV1rG
Z9g5rTCyXsa+7az6+G09UNF5e3rxptu0HfS8+IIqVRI42o/HWQidyls3ClFY/msT
Og0Sqw/IxcWLIrAfM0w4u/B4PhLvO+lb6hYtuvlyYV2R/rsbBlxyLDkz5POh4PcZ
iuiSqTaqty2V1n0iPNAnayMHcLCaLQF8hFmyptGmHpen0eOZurXlBCeCbRXYHIVJ
elcNicdpuIrmoOhnUvf005adHgqXrfSTFAXAXVIdDaBozj7bVbXyqwU1L2qFDXVy
5B2/EO+EldT0wxSGX8iy/4d+Z7ilg9XcalYffeDNDyRhExjUDiBbzezcSUGABTBY
XwhmpjoFc1rc3ZLP6MSqazmJNmnf/L6S4ebNWjhAcTibCxqxtFSXcDndjl0u+hl3
XbJVtLqGZiz+raUMBdakjUwmjHLWFOs2gGw4sZbmQE0bb5eUkurpUizFEK1Vtefw
ipDZga66nSOIjgjPEeRx6hyTij2b0BmSRCD4VtDa/eT3N+tJMxEChHST//WLb9aS
XI/zG11gMQc46ISRxWeyxEaXZyScl2dQDOEItclqFQe86Z6aj+is+58lZMJ3hch4
jvEjpIL6R8O+RFlgPUOYp1iyxLtgpHGkakPceEYNKgQ5zEuqh+kl52hs7gugs97/
EBbgpF0yQuOWfCgggkR5csjj2Mw0gRnAnR8Qf9rNwI8G2qhTntrfT0oWUh0sJVAa
jyhW0pFgKOcQ+qoW9bjhhrKWgvN9zqs5kEFrMottgJLnDsnbWjt0Q2aeqN3lb310
jaaUr43mwSxsz8cEOX7asbIZFywvLhxF5ZNQ6LcJJhUKARGoTOYrmihstPkJsLS5
lOYON13W4QbIxuLxdUn+yfQarzUurPjrvIan4HFUl3keB1Z+poilhGd2OaONDGkP
PqKs88Yx4UYTelaY5gb70eKvJGV+pvK/SzRtQh+EjC1i5Ii42HyYLqyDKAXnzmcb
UL7ZDtodtGjI9xy2IWXE46gtlyFQOZw35Pflkv2FMVy2f2OCkNbGlF+nBwMpAv5X
8O0ahBxGG7WOiiJyZyvxp+SDkDHyXjgABaP0kJli5fEoCB1ioKB929pkRddKrJZB
lEFgOn1vyxxjmV2Aa+PPCm+dxjGzBLzXxqBy5BEuu3sbscLINK9GdGIlU3vvZsHu
oj33tCe0buMbvIwOeYVR1EKJ0DR2EJHq5GyBTdm0810yTymntOmqo8A2z1oI89GL
Vjl041K+JkeKIgNZXONNmvMXAvDb/3fD2PrRsfSn7dRZnUXKHjL4a2keP+JOTDqX
4QEDFAzPw4RNzmY7gPYEDxI/Ec4+/ct46l9CbsvzMySWnmVzsvgra/jwLm9AJiJG
cSNjxCugWN2XbqLHGt4kpzeTsvCChLx8px7+pYFxyVMOAvxwhLHOfaRm0lgLT0e6
pyNMN04TOmUSPz7SkKwWlvwYb3+eUYojsvxywc9G7WCJvY7Q2aoeX2rlKJr/A1lB
PPybDc+0AleLUaekuGb1anPPETFngmd/wtiuBEGYC446Pd5gZo8fOPK7quVy2v41
imcwDR0gSOpQTMFZci7NdcfhwUnn59LunN1KkLdg2U1/HovwP5UeB2yTVJtZdzKH
wFvUxjDQXDZs6/O2I1nnpEvhTOqI8lXgXskrMlmA1RxJJutDgHllvANfe/LyES8l
BEOu5509HFTv8VifRXsHx81XHOMmhk9p8FG0zvWUU81fpJDdpKW0T+mrfEyyz/yJ
qE4GCxBvIsdJ2JG2TziLflEsq3za+8+1d7pfL3OH1UvCys0QS/1PWcBacGBnU/eD
waIFFpDSAS4f47jGNqfrOCzj8TRfw29XtYnxswH3v1dbGwdRYsfJAyX9E//qcCFE
LoS32oz4U/5pFSDtLb+iAgFQFcdFtl3XS4mFp2dokFyXi57/7rr3nHTaFsQp7DQr
2N3l2P0QHispa7kb9FMXhA2Pl94gxaKclxwowfihYCe3NyOFXWIpXyEWWOu13aMG
QBQxc6LJQUVanIbSJzKTK/B5GHjohk/8EoBWsbK1bS8VknNne4cVbJaHK7M6oFED
yTNrgof3qZBVUKlcOL5I2oa3FnzCG3EIT14zsCJYxVbwVlnCi8cPu/ehWtGUl+KH
EQJMQRR2uCB5f2qyklXE9aVpWZqV9kC/H+UBTgrqxfbkH4iwnOEKvt1aAfyqJp5p
bEVeQjEUpm3tXq2RC5BDhkiYyUNbolHHi9qFpgzDrn9iHmGhm6jotEi6WeYyH0Z3
UCLGK4fcZb8rtrkNayYxyJ1nH+3tOUhNZ0fsSnlaImdeg+cY+ObwgVBKyGYMgIxK
qKMdUX27hV+1UrEOYXVD/9gCUBsM8DSDsORs9J8ov8XXq+Uitiap4PF4GjSnAkCH
J6Tz6iluJYVeqI7JYhPwSCs1X3zWrnBJnQGsZLOxY07XGxewMCKxw8Y00eFR52eG
QAYB9CCmruXz9414rrXNYA92pGN47r8cCsPVIXNYyP4ZlwfwCU/JDPQ1/q7dDSIy
iWybDyAkrYP2Moe5jyh1QqPbEtR+mAj7JdyBqnE0qMOYKcReYNjPlHtx27KdFxlu
FNcEF/UwqJM+AhDc9h7N/VoUzTHlsfwJYG+C5XLPfyu/AuriT52Yf3cvvq91hoHJ
WcDUKn27Rh9g5IhzKrEm76owKzKjHR2UaF8MQmHbC1ZodW2apF8QEQYIK2Rm++2e
DjGiRG7BtZYKrFlfHV5ikNW2ZrVTBlNFHRVGXzgzSRmjz9m+RILIRc8RgG7Ovo8R
6JaZQlDFLhDdaSWsPja645OAvIVLIgcI9Mxvc0bMVJH7Cv/ezjRfc9g+T51xqEJL
oBC6dR17+Eipr+lSLh/IY0pCpp/aHE2eVPkF4b9WWd8SJBvT0QqB6xLZpl3SrRW1
o3hW9V/GwLaSxtfH9YxqVtgM6Q3mOI1hJJpczHoCU0YALbySF8riCTEA7QeaFW9J
CNzPoeuY87X/nTI3tcTOA33sANII0MVeyaFKd+LCaPOvvtQYsTdOFa+wCrV0MvKa
ZyDEt+xAk8t9lgwaejvEz6drP2tR8kUJfHd+lNz6hr2tNy9x6SEJQ1vChMwngMxV
8cmVfrEiQcXurzxz6AJEIzDFr8S+pScJUAtMjoWOVcNTBotEHefAI+dBPli2niqP
uOiGmPtDVJymdTvv8KNwsj2akf1zDfqh70hurYo92PK1XUHIEktYgblB9oSawAUP
atmM5ELZEpnNgZA2DRCAe8bpkHGdomduu6W+AE3aoICi08LYWtWcyFv6aehaqUNq
beLC0SFsMhg3XlBkrYW5BRSuoN0p9m2HpPOSkZCqVffFj8je6XatiVN5DDqOxSWN
kA9bJrXabtfaUswCGRxa1wHsJAjHybiDOxlRSUrRvqJ+S28j5i5lucF2TCqvB6/h
oFP+I2+kycjPX4LmcFkba3Qz9HhufUJ9ju97DSpdSzjHWj2UlYCGd5T7audredBD
nH0SYf83BmSTRNZb4rZA48rSe/S/XKX3EBP7znaAJlQ+YMx+ftky2ipPzYfpB/6l
77dMcHoNU+tELO44JJY3tPsgrC5iiSn7G/ZF5lUA5vhDGxDm30Zwg976TiNNd6CK
l6hQ7pAMYXo3PoKCm5NSKBmhisFdXm5A9wj9zMg5eiMH/meOnI/6aN2wKlTdAg5j
zahJ107L2ii6Aepf4D+HJmEKBUuFiU59wT80QBSdg3o3pB34hm3Hc8K22wgjotNF
wjLMXqylakVHfijD1up7YGM07cbF8rZYqt99u4nOvFijfN8/J1otL3fhrYPBvjuC
H9I/R4tcjHqdoP20zUmcXrG8Zjw32zjPJ94+qghSfxE3STI1mVzpbDJTM28drzin
/lf6QkAi1UsVmfTM4e4dTbB+2DHzVZaMpMA8TSsl7+/XpzvBt9Yfe4ULLWQnwPCn
3OoU+Q29FK8wF7AkxkkhgEgLGO4tPQoHgcGIRN2plSajE8GbxQUBxSpv260Ydj/b
FTXXd2ccweg62K71D8vYyVnTa2m22FMTW7TMQUQ/Hu8lwkBbmzfLBKl3ORxwDuzE
TPzgyLDSbqHHSZYk/Wkv3q+VsxnoDF9KCkLAaOdRRkFUm5uk5CUudt+5tPj+WLGO
G953+4q5ecHJGwRkzOAUyVD0uf3kDxTZuNl1u3ec/RhbtnpfQ/+539jSepLhX+8j
pBg70PkJjH8FFZyCBGmns6D/kBPy1zWu4Q/HHfUKAoKPlFw6q9hqcr71POm5kCr3
Ga9LEwIgoIe99EfxpAnyz9ULptLpiyfLSRM16l7oLXv+J1+R1RaghYNQgOKX39/k
yRNGsgou58yz/NM4/nV4pGNzaoX9AT0f4WJdwwfDOD0FM9RBUT9tFwB6L1NeWFjQ
MPpolzcQSRYVdUOqh/5Vb6fasMSIV8AUBXhORUTteOpi8T1BYZieDge/ijKYjlDo
/AOxQvOZC1afrXccMCuy7uyiQQEYKg1qWp4/97znuA1GbtVxhDMfbHQMdnXMhZx7
GL6NdDCizBXqkIF5o+VMqrID2tueOZs1pCU0ZF4vh2S/c7b1JJD6bZ4oO8k/jPTy
+Vum5ZOFCmEO/jcznSK61jFadBepWRyX/3e27/nbYvkDCHy6Mxef5MMuMdcmZw8A
mkxl+7Jh71mCx4oagepf3/P8M0tG6JM8DuKB8jyZdrr/4CrGxTwuMuDbcKqVxJrC
uNQqTDifLTkx105tM6lADzTACpOu/OKCgC3fQV1gjEY04ckqDHMXXPB7xlkkVX8e
2wOgNA698Jmlj+unKeE8JNhk0uEkOX5pmqiciw7I5QDjvH4FKyEmvkusNGl5S6Ke
T9kQ+ZUBgz4Dwm15UnQg9yNXWsaxueHXLpbu1zooUnLpzr/xF2JeCh6kJ0++4oyp
DITPt2sO3oQUOrnnqgHPjF/PY5lQRsbQzAGLMjnmKjkzU6ZG9ZPfY+Q9St4t6/Jw
yLBbbcnjIJhhSbhT0r7QapcOmbTTK7Gc0T49nfLBTAboJ3R9J3Ip4hLjQ1Q8Pujj
MJGN4c+/9y6xY+eYLCuMyQNGwnlP8/3CPbuZ93vSdFrG6F8Ei/AqIyWA5oXmKSu3
caZz0NSca+xHs6rdAA8Y58wv2AwsmEpAdSosj8R6jJl1HueLGAl0HflzGLbuNzCo
bp4RVOzd2In3kfaFdZ4baJ6lnJ/M1+J8JdGcKUkGFF9BEj5PZS5UM00j8ip6L9VH
UbgfZeEVYGs7YMowoVyQxiz9V0jSXNQUqxh/Ba2mZKLPvpXC6KEyQMCsawdKQoHm
L5GMQeeHRvm8NqGiCggG0guwBhQo1k5eNsag+wdHrxN+CsdO2+rgYCfMuwNvRf1C
l/7Xhyfdff3m+wsDOieSeJEe4Np9cdhQeS1jU0mb30ag9V6FH9m8GkTG5TarmDUN
zEMi73vy7kIWg3vS1md5jPXFnn/TcNQemHmiVz30FXN+6XMOEe/9dKlZn2T49evt
eG/xvYLhKEKNe9mlVYmzsfIbXHgz0xMuVXJCThaVZ1w/9Kps6Uwd6aSaLDhxaBLK
vyZcUYrjukn/FZGxCa5wjIkj1ZMHoZ7cUkPiz8Y2lWxRXMXF0DggvUkZ5ZvXPwqp
0dQDyiyCQn35KC42gPmkCD20T7KOALysy44fEBdL2jEL497w2Q27W51FGGJwXGaS
VbZHAUzgTSILySQcSrOVXxpbikefHRU7x7xjica9Irang8/1HFSdhcd+IbL0QoHS
vz7WltAvRh9t6IAuXwIBh/yYAGA5dz1kpKSN/Zwwd7LbFzp8jBPXmQs79ckYpYde
vybo269MtjRnj1eS+4FUGWjGy+ijnK1e/vA+pfpO3Jm1J7QxhvbnMriyOfczbATC
HlttKHfA9+hE7SIdkzstTYIuyRj2TUk70xbSuzdsZM0ft0hTKcfw37r0PoNph4pc
W3P3xOHDfN33CNNJPGRgWhl2wh08g1g/ebt8dFytX3hww6SfBwJi51DcQfoY8Imc
IMEH8a3C8Or2S7ctFoh4cNNH6zUTLFs8erGcya+5I9jHWbWVui6zIwf5KIELHaeJ
GCJG7bkDN9QJeDBmoHGoUAT42/T3WtQXbP9eG3QXb0N/JSAOG/Mgl53KTjATY5EM
5QGItpPr6wwpZYKSC4QfDVM4/NRWmYi4/QOIBzQW5mDJCtUcBHp9vuzlYLWDE3j0
sWtBTRbdFzEXUBa6MvudDf9vux9mQYJLKILRnnlJyBRr9W9dG5EiCFiT6dAqCv1q
hDqWqFXA2C53rXQhbvPjOYavBQeR0SzSaC670LUWcZ9La8A7zw8vq8HJCXJbtScT
4GM+zT8lv3zYFoPDQpafOP8i0cCZAIrOidOg9b/WHrExcN6gTpauJ3A+3GJtPZ4M
vYKZr05CMHup/nKbaLV9nzh0JWgiDkVInYKhfISKvRNO2FOxy9do1DHfMYnvxusO
hd7NQ44UldTffCNddAbmEqlTPIdFEQO4RrcFpY/EEb/hqGcHGAa/7x1g646ow7So
evS/zvxm08M20dQqJFSNGJ4O0NAWqz7SwEDs71iFhXmujY5mcpFBYunLixB/BIk1
4+qZT/C+mq0GCFLhLd/s/6fOOhC75wWFpVmFevVJMKgXa3FumJl37qoYcVGSrXEO
tEG5DRQOK3uR8mRmEC81PoscwrKpkyg4EL6qJFKnXp1Js7jAA6Nz+YHJqiRwE3xD
Wz+XfSq+8KfZSphlsZ6k4NUftCoJnT/WH1IqCR7j9tRA1AXy/+1LP6ug45fzQ2nd
v4MEy7kKjTj9Sk0PBJRYm4WpeUYOo+mRShMUKwRwtNe02rxinTyFQVYfZsMla3wS
vmogXYPlir46hH7vuJGQqZOyMuclhSeZqECxxr60dOCtZGE9FYkrxuHRk4Ny2raz
lj5sMwWKm14OutHr8+0vG2Op/+qh2mGhyK2JUVnCdGLqQe9BEIdgYJyS2IWO4JDB
IUaW3GL9w67IVe09OUKArZCrDaOQlv0baGkm8dHHNlcve0ig4+H8iMaiM7/Ixs+i
V3C9d7ZGs8DMEG3wYSP/F8p8s5zYtMRar6BTuAkNTPoewGSdA/Y7SS0x/gr9mGiw
lYzaOWJzM33nXMqSjy69hNtr3/hmfX7+Sm60Xs+ObSXtAoGELRjBzYztrHyGYpAb
K9OvOO4DRDyNCObc2sjaFQ9Kovlq114OfTgdGVkn09juyZPwPjZLbRH8FrOrwovU
vKydfhWKfsN1F924hzBP8RvhsjJTBV58Dgpn9G4okrhZWbIYYl1Hf4t9NA4Vdhxl
cpgHlckom0zxpDagF9QHjP3Xknb4HKOaVy2hD05cXN0F3OvYA5EFOKcPxhC+YwaM
CoGNhXhYe8lWgIgUwGgdJG9rzQjOU0zM84LmMnGd0jAMk1FHkWAoX7JteJI28Qiu
jrYSWsqCHue306YFo4ksfKuBcYaYSQohd90YDIPQp54Yq8KGyAqMpp6rIpO2amsu
aH7NGeaP1AGyyi48/3xMA8Z1vEASXpo4p3x1Ryn4OMj1pG/diz43LwIGWqA1iaAd
tudS9r3pe/IBQpHNYOkrBb/WTvBHqYMxyZpx9Yaaojhi6X5rpcCpkLzsYreB3Zuv
+LoaMYZ2olbU6giNgjNQuPoF1hHuvKWqZWGtanhjBuuRlFIXNgheFqPxKoVlGipg
EofB7lmOTR/pMRYEZRqg1qrrkWlYPy1iQe3PlRe5krF7iqeF6fcNMoDQUxhB6UtR
v0PkEQUd3SN1kKrBWwK1DCUWTwHk0L1NEhi/GTbScEO/t9tjehPvj8xR9fkp2g+b
s7+/AwFUXGeHQGrzRCJ9YWCPyswCMnQvP47hEBmEEjvWRcN1Yh2YsE8oL4Gn+Zk6
+Y8IIAtPejPngopsquJ4WJYsmWha3B7V4jFXsPRGSH70EWvQwbBCNF+X03L0BmQo
H6GAYdvCaM1ScLZ8U7imJPLf/ZuUVUaJt5uoCJ1MOPYs5LMGfX2xThY/DCml6lz9
q88cspggGI16eEzSQeMr3eVhQKRZdZ6tX41+DT413lQ30USTFMeXGZYFQdO5vdt0
XUP/YJ3Yp6eKaVIxk0wvPWh1FAunUuDYcYU+Wgue74q0+/NwQRoft4HTwk1hZixm
DqeirkO+P4dAh3Uk0eymJK85YPqTlxNf8myM1emrYJX7UGx8V9U+GoCagotfaXQb
9TLOzGowiTN57vd+WlLsWd/DzO1ajkzVJtbll7cChIfcb23lR5z3tKXTExWZdAFo
HlIWYjda1tNIZ9TvQKuge+/Lhfc17BBFlSCkzweMywkwJDdjb7mi2V4hSRr63K6m
islZhPzmrzh0+b3uWDJ3BeoDH5YLh+OuUdVJkEr/BDm5LjA9Q80o+XK1/K7WTNi8
8jDwVErQgTUvvQnL8fi1RTP/r3UZ4Ulhjt/C2/IlucukzDwbf4rl8Ke4Xq4uv5p6
3yhSBL+sL6fQPLO4WvwnWk2o8dqfBudBqo8qYTann2/WcBgozQUSWJS3DZpxVM08
006zYJQZnH2y1FQwsgVnJrVMQfFnsVOhhyyEt0onyuMteNZ3FAQ2s3AR4iORQ3va
LXpxZSwBhpo3onGymJOJkACy3tgFGCCoDorfaHQQMfv5a0CI0RX0y9Azj1DD/LDt
Vio7eW3ZruWJQDEP3qZNZHSY7atFLPNPMjIwctDJi/p5kPecDLO/FphvfPaP6+sO
6cIq3tSIyLlfLkQuj4MH912rUT7AQLStETMHM1kGvClBxFGATSVfQdj37CKdAsJi
BBZw76ksZ35ve+ANsdvDmmh4NxtlivdbVfDs0Uuc7bTBHOzcyos3hOsCmhWrCIs3
kwKCFy07dGO/kogQeJyefNYKnJ49w8DVTMC2xLrTstAus3fTV5P8K7/HXI0p4WBa
CrOr8d3YTN4FzDLt1ToqLzCINexg7or7NMDXfHuJ7OceBPKbHlFUO0FkYjqVJjPW
YOKfttvck7PYYSrfEkKMezwZxBYuevGuQVYicov6fWJIDOq+E1q+9TFct7nFLYxM
osJYQvIWHCTtXYWle0q0CAkRt5LAVo8pTvWr2St7N30Wccgx+mKb+RxB657PSIFo
fK/iq2Att7T4y1NF09d0tXWIntYx1F74KK9oazQFhPt7KQxWWqvHoAKHmdOYNRfV
sbo/xqNsV/Lw0gNp4w2oehX7Ij+rvbSRfnOOG9GN7aHA5xv11vRgpBEIeqSrUDx0
S16xDIgH1QYkalk6UD5PiVj2Tnc+dx6GSXG/wWKnBRTj5jSm1KsvzeTpJfZB7F3d
fcBkSPvLWBOAOaUP+fHqX+Hqi/AQ38/pihtcGCyTFZIidg9lpwGXIlbGyC049ZTf
HMaTrIYnWedm+rDLCALzOIbpRnjpaxx2ux8HOWpySjB5TrbATFXJ3KMPpvs7VEbG
pGegoDHOAwWNWREGvRrp2FM28jzFGSkqDGRuMzrbi5UN7nMxpV1+qptapos6GWEI
COMFEV6CFe+F1SMk1QAHkixs0qT7C7OE6jpgmfgQlekOyO9BX7t/qozWrT+4RXPH
Qw3tmAzyGHo9kOK/f7c0qt45xo8J+mGWOWKjmcgQaxPEfN2KD9l669Bx5X35tu+b
469YQdRxiAdAxJosX013sGOiFbNt5uncOJDAOqKJdOK6Yg3lwpXxR1XjgS2IyrBv
LslMk9gNXsJYncoYqBo+8ZSwTanM+AtVqgeaSkIUgTc7mVBHuUeMdNj2xRd1Hw/c
+1ba4pUYL/9WJvzM62RF9u2qc4yGHLCMDrNPSbCuAemM0hkCCwKdDneQRUnDcpnB
7MNnvUGoPLiSEI4WWHtN/BhfLGnSOtcKO/ftrkOOG0VLfDoWIFKh4G8w3R9XHAHB
jIjqu6d8Tn4DTfMIy4LqIHQIGjFCzXul/+6jZT6e3XEF7Pey74kdQTPAzpp8uU0C
YhMFUajc6JcTmadfwRWXq6SAgBeR84Inw9y4k4phZKNn/MMF9pPhvS17CW+0NQjB
t3YtQ+uBpBFThwCnfvKVorjXkFXajFBZI1DRhOWYigR3v8NTGpU827S3k7yp55Uz
CBiETNGka/V33XfzwMQ+Ily6V60EwYFN7KkQAGXwBFpNe3bpwWz1lCCbO1bG2pVj
jWjAkByX3VJyzdFkv6INoWyRQVboMohe4s5sKad/iWMdzV24oVis0eOodg+CklAY
PhJ90tm7Gu78WXQXd6cX6kCA/NHYlpenC8JEc1ayj4xWz2vUr5qMyQR6CiwNZf6Q
OObZRQvjPlGGB/q4PAAF8/pBVee4cTg1KJduywy1DEM9cE3J2Ar68bF1FJiCk2dM
MMnfvfKPNDE4PzsIAQrO/S9lk+jISL8pKOgklRjrMiJeS1X4YiEB31tG6fvXAc3R
JgbphLl3QLUrhpsH8g6YPfH6nFFhZRIn2auS7q4VepCKk1k9v7ntEa84KY2Y2gxf
kQq+Pyn1GmK5X0IS3lzCvyYH/pe8pzj/PXxXQ7VL2G2UQisSkX/5/3WfXdRpmu+r
Aaxdu8H27ZfMjg5kX8v2xoxU4V5NeWAs3cq9mx0kfc7hb+dyYBsT1MRM8M4GLBBK
dggrb9mkvTGr2DMKMzO4Ge45NPGEuACpF/KuJJPd8On+dypK/RmeiVbrxScxnDmd
TEkld3E89Mo8pwNakD4VxgI5mOo+uv69ei47SogJAwFQrwKp8L6ZTuiT1KKmKJ/C
CuDaVpiZjz6BTkRxtkTcxIqZJTRgeFqcFbVJD0t7Ugm9fbPpC/HqzKK2iLrjHHhO
HVyFSxVIFDX8EOWFpajz9jP+SM5gCspBm4DXarS+iQnJlmQRBDb8Q2LeZm4Re9RC
RPwYABS0cHLZFDZQ7p+REZpuMZ2IVRvBIuRHAvrP4zKr/iywArIcJPXZUggdc7vG
Bt7sAmvMUcoqLeOBLVPQzib8fLRNzZCA7FG4hfEEyvb2cXXRhVSrFZQwVPkQbODy
KQRTVAKlbfXnzjh3GfctlUPSN/FO7vBdXIxGPuMP95zeTzqw4oSa1XPNxb/Z8WrN
FzjRX5jj1v6rvMjzsfNrID3hCu4zOuclX/rNbYk5zF3WK0MsmK1TxwB6tMiGcstq
qKjrkJuyr5HzDFdr7eAVC4fgy6nNsU7/0YtQtaUMeZ3bboeqqdhqq7Jn3Mx7g6PZ
lf6E7YwbPHgsb+uyTGWsHtnfO0qSTyU+J44PDSHGp6lUElxGmkYDb9+jRr4lNl0w
h1yO53tDjJxL6Jze9NPJyTTX8qVaVX9B50U5h5gP01sKk8kYRT1v9miEpk707uWv
eE8GL4Tz4KeNqhAJGDFJ6nXmggX4KhkDmrPrAm0EHRo1jSBaagWe4Q5LWCQ0eW6V
ghaoCtaQ2x+fLknKlKlXJsMXiPTEcI3bcPnFg7Z564hfHScVv6kj1Q6WXF1teK9g
Wkry0r4WE+lXhzX/W2lUhxShliAeFlwx5OiTJOUxSjbKCLftwJZ15gRFMbsid6WT
ASGMsVuXzmOm1WV3+1mj4XKuKn6RQNsIaIjdkajqTj/Tf7WxJ7HqisQj1GpxSDja
nZGtxTTk4eLda3nmLX8L3fAQ/Ajp2pSdPtEe+V1pYuR4HNvxYYBKuRkQcxmUJYzP
qyeBKvPAjG+fAcRnVj2VOzzDfHvLapMN5He8YpV9MMrQVF+yWY9H+7TiMoSWQAjs
9H6vgbA3ElrzN5mhX+XZ1OBKXDiMptoIUrA3DQK4lAhRX/4rW+fELPN69BTlHPmX
7X15IQhUHVcEdxvKPq9lhbTl5PKUfVcKszlsnnMX0sXNufaAwVSG2bAoDvRwhhbE
NzhPYmDYiZqOFESqSDjN6Oi4WTtiigG+2yASXqIAMdVgq381A2xmPmYJW/8Sci8a
A6vq9Ph0Q+Jeo6wSCpX3IHa3fOolJfWQD5Dp1mYKeWMxSPgjwYGwkCyGIroBvZaH
hCzTcBRbukJdmiFK6UiUwB3uG4UzDWw486W+QLa6TCHMvm2kGfCJavsn8QZF3NKd
+rsgFQsCMtiqLp1R05WcBbvIShDAEledAvizxE6eCBiT5utyRjYnn71dXBLR5YDY
dU2aJqdKeYzGy3TokyJoKCvoTKno/cGWWND5h3rwDUkJLGl3yNNXzDBPgRp93eLf
tJlcgQXTQCxXX30oj4eIg7tjmHwFNevFD9iM1w1RUHjf/wi15GkZvM7YOcIQgzXH
thhb1AA2F15gAmYfYKDncOzMSgTeE8H7jVQ2FnI4W5lb4WUphhAuNfojT1bOoDmn
YzeJBZU3uu9ZAyUGHRe44urZYTC1+KEODcRMswdlfIjJRWN9y1393Ng5aD7YMTcZ
p3CS2TVdhYNeq6Jj/vW5iJEg9rFgthnvA1WCMx/wz8G90DDLPz+IHIYbmxph1UXi
CtWYDTAR7OLUybQep678hyS+DnrmrgAcBInmQ2HL0guHleuKrhI+YdYgSjg7KZq4
5h0jkjpmBt6KUIrc+puHWCxLTZMw/Aa6C0eojHavkRONT+V4gnODrDBi7KlYKflE
KCF1RYu13QkLleX23rTvm+Kc7KNfuR3KixFCyFMkU4HqWX4RNiFH/lvRpOW/l3Aj
aAWlibxteF9uAKcR4rfk2TD1P+1PEWWJskT5708X/NQ8xOtUkSLvl+fFO1jv+7nk
3bWRWGqRxggyGdTTLtt8wavlPe1IYXLBVrb+L0vVLqekGCrBhMmPWxVGfjRDaXxA
kuxTcToWkTL6FBQqM6ii/fj6WBsd+F53NLOPH8cCbHG5NexmNOkngqsMyUllN2E8
h2Fhi6tHvi4iffIA6tFInGPcSQkiCSgCbpM0kRaHvIWT8IQdjFoq8Nvezd0zNy1h
meO0XRG8wkXeOqziKGdUR5ceoBrxIr99dCvLXFdI4KikWRs4ojccJstQBv9gO7/I
55UxN3ulIkISWXuK+uuZyRxWCbtCbSr5dcHeyncsIedPE/koWn59Qwh0h4spm5po
iCafVS6zqSLGFcy4+NALI6IanPiXwpl6GFhB7lysWkgw9OGM6mvPWfEK5v3H4CV0
136N/a9zFK8ZmbjrcHbaLQb0edPTFbhdb2S2Jkwg0YFzdDQHoxUmIG+JZpc8IV9b
JYMrGASWc61oj/njEfoOQ3E6L6PxPjX31renATLRMTvAb1WCD6s184pjaLLqngR1
22W6WxezwmJeVWqyERO8tnx89SS9Sa+XlI2J7nTO6yTZQBQuQAFHW0e3ZRcTBtae
LeDpHyF68Gegt+evudhYY35cTvmeV1bgbnRvasY85hteAQR/IubNpFodM0TNXYcU
xVVjxgzl2puyyVhSkaXkND+saVkkrKp88ONIqd/RD5wSoeiqh1Rajf45AsRuBMPG
KsnEk48J5eHRJaYnIZp6sJlL6Pr/VaxkBzN3cGPIGbRkKRFObVpyN/x0+dqakOzb
K2x6jxwUQmw8AijJcQHq0V8HTt8s2kK8bxRZwORYPp1VDg9XkvoQ4Ca7+aqbMdLE
LTP8QTeLmBzZIc+iTvkot7Av9h1AA81oX88tSiWM5j4F/VMjcAnJrp2/NI01C3e0
S7Dqy5fcR2Jv4zd9rFrCfyJeiMfP6QKy8wAAqP6t3CIRq7Ap3gPq1wtGamYd4/4D
5qe2IwplcQM1qoUXhdjYsR+gKhPDvtex6u9GXPlEHRzEYZ5EUSQTXMFk0qdfs464
0K7NAkcgHuwCeTF0lE46ykXfaHJcEwaE56D7ILqr8Rhl4Gp/ufzvtoCToz8gD8yC
3XZzGN5tav9OalFJVpp7SVuZyPG9igSwE7wJYAXznozKJBrK4hC9DxcOXRmF0Nov
cBsRSUhY36Rh6gQUwtyP7/yNQFHb5YX6fMMa5MaeuiiRMvma9WnNzp+I0bac33k5
kFjmCBoyxIo4h3ejbq6FaYby5eC6KpvbhzwBIDi7fx59SmNAXaiq9dMtt/KUzTLL
fOWdNWYBeRpV7U4gLL3ElRu75FK4fBvKhH0DFqxx7a03+WL+Mz+1dzBYaVHYOrsu
LzARHulLrt7cKZ+f3M4nR875uxky3OpMUl+3kEB22QVUcZzSLLHhgbyzcJ3VsInc
u2sJi7o/l4crMIF5dql9ndl1AcX2WnCLTnYJM5nRV6xkgPoFW+/hHqxr7zHdhE9c
9gBQEZ99GCjOXkZ+fQ3ti04oBXnUf8+ytGO1GQNdG2ro92vV4Zsgvqot/mkhcTwR
K1ZcoDLVmk0CijQD8gvINlOtJxfo71Rfa5kd3imXeZPw8ZAit7y1xvbS454j0RgF
JyWj7KVuPVSpulXzmAkaP6gsmbPRnomtPYwvl2QFWuELAlUMb98g5grHEj+5r2C6
GU5z3Cw4lp2cz5hRsblofe0aJCULcea3fjfOK9Chwi9UpUmCoAYzyVGModguL7r4
QC6zevwDE4giY+YnVVm0ueFjXdhUoqz6prBOFweFXMzy3Q3YRRU1g6LsbKMDccbs
soxH2ZwP2GHcS6JbiusKwNaiNV5pi5gg2X6PlLb1rHKMUoELa2SqYRxYKNg6nxIR
N4m7Dr7tF9x69hIHy0I1ovTbLJf4ZRT7g+7vIJAjKxvpemqHnZQXYcTqD8HOKM9W
RlNhe4XyqXYt509HM0I8GacBTLzSp+n5M5RlP5UNB1oSJ0G+nQnsp6Ce7qr6tO1u
rrbNNMe9GZukfORQCnl899NQVWdcvHRkwlj1HxYi25tPTlRp6pw9VqhJqdkbwKGS
2f7c9QfIpNTO/vOw9urZzyFPgA9Zcr17Y0xIqCuDchWwvuluC8sH1ePbdT6N45wn
CYfdEQXgIgOY36j5EXW+ygvNFIo6dJKwU0AbEOnzzPLf48We3FZ5x+4BhG3Szrl/
synObsjo8mCN9M0wBfqEXG6rOPnKYRa59/Ubm0Td58HkkkW7I0XG25x6HPQLtsPk
m4/FrLIyknOJdGDo4hFLCz4z871jsmnMF3DQPOX45GUEIqyjeixPO4wNIHYEWwqT
eXkz/c6kdTALFRruwwFvdye2Hkg3mHXuhKvr6CEpqgeZrQ0R+eoG3v7gOL+G3FLf
Kyi8JHmQKJ8ebI8IjGZM4iw8uSs+/jACzTP9xqen5PVmWb/qtJ4ebgb1huwriUl5
Uu0htTDDqhdhrJYTAvLxxkcxhsSQUovb26Xl4FKvD8nzQ6JgyjgFUc3oB0pLXdIs
qgh9LkE1cO8sNhbznIXUUEM4fRZ8UgY2Mb4aSppFqGj7DzIIg8rd773OEgw1WOFb
22215VrWO9961tTRFlOVpkhOhgZqYc6f1LC1zkcupMjnqbb6zNyuQ3DMogLmabhD
uHDxStQyEMz2vYlPqG1mEHJjSlB+lODTfLaYCehTEPLN+L7vJ0LUZQRWlB328PMa
7quVxrVaHlNMP/0LXof4ORDfWpA6+nuRWvcA6ljFJ+8udjsg2kmqaY82Bxidq27h
fS6jXNNONSQSO3LzaPtcwawvMCbODb1Jpw/0710hamZ8Z2c6hyxz00oFwtYfeGI2
jaImxxV+iP8D8mWPgdly5A5Ktr35nBAN3tqzNtPThgWwitUIkOJgIlqyk8r0CbkH
cL1srtV+kiguw/CmC7IB9nUkSh5Hlg+rCLjktz1Ivs2jO0YwWyiF3jT4XYt1ozY6
ax3Frn2KmznAngGxd35ZMxWUxCIKfd1+HwaThDuU0pDFKF0XPtPi25VxuLBuvhQA
hYKbZ71fis29v8RHNOejVeAT4WXjKSoKXtI83C0fKVErRxyHH/7KVqfG7tJjmr37
a4P5H8Wvijo/jorEcvCaMiZDJ5nG2+A9VmYj8IzVuRX6stu+4O3qyT3szeclrLcx
Tuu9IfVbwxEeVXB/+9lznfIVwAhxkcVsVNQdoYNXaYKCl6EisUw3UZ74Ej8D+aSQ
Vwm63l+0UfA2gZTtLQp+b5hdiTtTnZg3C08rblguqjP+CQSOLYheNz7fw6IXoy6W
7rW3pwy4fUth61P2DUzdSW9zhtdT1FCFNh9jA2JD4f/GpatZ9TaOPo4DlwS80GA+
cBXGJwSAS9Sa6Q3oWzY0axmmlDdYF+EhbEWBidnxBPsMLZ5oWlqKSUDgscKXWwZq
zO2uhg0A+cVF3xGmBK2LnBX8dshf2rlcXKNirXu90N1V52wtnynbUZGcSV4tNX17
UuNINSMwm45w8C5nDH+OUrKH4HbOL+IAnvPvUUwU3rXC6iaK9NN2dN6SUu1u/+ij
08wM5l5Br8AjaqB7NaaIgFdqFrZmHWJf6PJvMobzO/NwIB083+mnD9oSbmJ14cmW
LZw/Wbel9npyK/HEC+TK/0MUndlIY+oSCCcqZYzZGGa4izOnvBFebVli8U52XMnk
tT30940yMLT1MUOHMTU6x2w6x+DsMhDd34qU4dAYKg+YvDKAjbdGQbmaTLEuQLXp
bbFOMsl8Uwe0GOJFfyTb0NHRPHCeF9cfWCF4gYtQf2mJZGCmRI7ZO+bZsesdL19k
Y5oei49rE1S9UyIfuhad1op92NUwGU7ElX22UXhQC+WaFVjqcq0onAO3/68gdaa6
UE/+uDh4lFVj/0jFQGd8SHHcDlNqIj/MhEFJvvq5g3r+Zou9PAgn5a+js5djHwLb
d66ZDDIwrrUO/Lp829eYERaLDwDhm80LKrwB9x0zBXxI9UqNBpk0ELDHthTcZcll
o52MtAyKIK5xTGUZi1JJt6pIyLiWM6nXGAfiBDTlwuhE93ITahlO6nh+BpYO/jhY
wm7GtwwmJA9k7XhiHgQgXWrj46YnWULweKqd5aBfnmT8535Gl5cN8uYhEew4Z1j9
Z9rQbmsTYkgKi4uwHRV2ZdvXgfISC2zkYN+GEs4SMoxJCPqvww98ERinvSWMZTHC
WnfD9PAcSgIJ/IzDpEOwESt1trvZhsyg5PpWx+DLSJua8HW6R5v6GbtAKM52a2Yl
2WfCknUu8+vZai/q28ZRXWI3pmD7CBgkz5DE8jJV9mgRUPSqbUjdfOyYM2JMYqYf
KeZeYUhbLTnh/+UaCMf78ukC/6bPEi3WZUHyWmnmPGsTr66ADe0ELyOk5ZUGYZvj
uLybzCnd5r7xf87B1l+B/9ML8mAPJ/ocitYbZDe3OuLIVT7XDvgtFlNoY0ADT6sQ
KtMEg4bMRw6Qtn+kA5qz6pvEC2saFw7tYWtmWw2FEMZ/9AtFCvH+veH3TyTMah71
ApOFLQOxhL1MPTlEEtdc6fC8cNLfvtS2ZXrSfGGXRKr0maoFAEEYNkVIy6X5Gl9S
675v9KlUp5b9CWEdj5Kd+32/g/Zn69jiHY6whLQXiA206M5JFQn9wUzpbLOxnJ7I
efOx7nxmq/k+hESFmeKNtK7yQ5oxKLS/fjzQJcnFC6XKheV90LzE96EsZ9PMPZpR
GVSYTv1qMEL7gTJnjhQNSxUr1QP/TCLmKA1oO5EfRu4lKUbZ+/yWjPcwj8USWddg
fF10AnLnVl/nme4/hs9EeEEIcZQMnkjQQoLeeKOEV9dNYopJTXsidIFM7H5d7Z5Z
vLPpaLj0H7q2jshxjqu/dEp+9GMkF5TIBNVrbA9fK3yxPVNekuYt9Kd3B7grS+dm
DJx4TN/tTLr+uxqqSCVap//H0az9K+OeeZ4z7YIPliMljCL/EY6IZeflgPizi41h
UYAargcYXvQPQ9VHSWsnK50dvxMux92JDeH0UE3OwInw8khHkWgo27QdryAuHscY
Mj/sUhl/TFy6NNnGlU9onx/6eOR88ZFGpBARESWL0Uz0DfpKihooFHImAoTphTtY
bg266NTkAdCuyLFjR3d+2Kygz4lf8CMx+j4f+FYB5gsRbJ5iyY1+UME1WfO1Y70p
BA2rkVR2oE6IujFVXtUZNwmlnM+Kg4vbKdq36moREtcwLh5Ct83PM1au7rHtxWn0
N4ZTCSAToR857+l09b5/BV/4g3XhL16sMn85zdX2tPqNPLSA/ErEGSLTiX1q8gS/
ac8GH637bXUCh2GS0TYj7QTdUV6vj2HIDIhEbbbYO8zZ2HfIyCrxpPWO63FCGZN5
LM7URtA2N+S1/VBjhfAWk71hxZqwrNnaZ51zXU7teFBSoPcvbmByOkT8beHDsR3h
AckkEosqq+zsgufNmhdskpvPuZ21GattStsk+sncwSCttzR0WClicD3REFkvjNUy
ED0UHrGXaNQcHq1horCf/Vzh6HxAeoAqc2pi1i95qFveTnAu4F7oh4UNl13es5Ll
5HFPuP1j3K533mF9rd1HrgjeZexzihcwlpGQtNQdgfuKd14trXeuiTJ4Nxa22B8u
03w8styxBWIwTbxLDCaLKyZloOwhHc0UIT+cT6Oa0R+mE1trCct9HehZwwEyKba7
WO8+7ysT7X1UEcsLbhjxsqUIPT37ZNWsQKWubEKE7tiCFxwRmf5JEudEwko5Rtl2
mgl8lzkSU9ZLZKYYqXj8lkMnwgNuLpFWwjZq/O9OZVyCIXNlnnP5d4I4Du6zYyak
sN9Zgl+q2iKKEvZSXOcf9NkC1RmMeu2odkZ9rWat/oi1ACp4WblzSHb7rKkM7THK
tOlQqBjhR/twXGf/EACiwXH/vHfOWJc3dH7Hz9Zv5uF67MSdcmf2UnysCB05zUMW
B3MpHkSqRb9IqsjoBEpVvibfijqjSJaXk4v9QE2kSmMuCto59c5MmH/1BQcr/dNO
D+wN7GLXvHSMOuzFN4eQSQD2oDxdK+zucc7kQ+n0I2rUeDWao3C5tdITg94yXXy/
exqyLO0eAdPySuwPLienmqgVeS1WE9uTYTz1fLtkEexGfL+oDYhCQmYP+ldvs1Pj
PWh0MUaFdRxsyR2kCQXjXMmJcmWP971vTJI/56bBPI1adO6gXek+A2eoFf0T/LT3
rLQGZaPOXfvMbnCQFPypnLeeD5Ry58rK0NmrSegUCUNDJ5b58DbDwDdcgmR8P3jY
r2DO04zYEesDe8LnAUjPO/s27N6/1Ts5Q+RvX24hlUeDbC+yi2GYwGqW04FggMnR
4bSroj+GWU1EmwJ/7MDvLaroYJb6POF27t2RbMxJfpTzOyATBGdL9G5r4jY93Gh+
pW46z5N+ORtqq3N3FVrEFjEX2YCDmJpBnZLtFLiSYYGCVdz3ujGon3bJsR8B/XSr
SV/+/fTsh9dgFkhwL+fFXZn1wIixWrpu2JYQiv62+XTDBh283jauJMgEM0WlTauu
GSbdxha26H33yYZepaOkc+m4F5szavhsy9LHyRIduICyd+Q4RVtRUZ0LXLYN4nec
iHzajulOMtv08fNYY6f7JpqJZCyR2wAeHiAsTeGnfxDWHPiPmXH56OV1CIrQJZvv
fAuD1SY/WArc3DSycpxG02emacNmDl5djz2QJHzxes/LO4fpPQxGHLVqTswnbOM9
i3I5704/o9BANPBk2d5lZU5Qxddz1GZQZ4Kdo5TzLkAcg3xVApaqwWEdhloVq3gl
`pragma protect end_protected
