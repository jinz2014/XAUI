// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jweDjNwHMOYum2rN8L+9n4VT0HtFBq7fyioajHSjep1gClnSATzzudMARpxOPJsB
ZtnqPtSvLvLBpqH4D1HA2iAwvxNGIcLLP3nYFFYE6RjZYGOZhUX9Y9jysHcuFfh7
7MKtYXR15twxSuTUqtH9TzGeB/IkNeYy9ZUqGEkTElM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 45808)
zrBcqpEP6l3TgEt6uaEthnX1W5Du9bEcO02NiT1ypRUwDrC/nhpM5zDtfy3v9Pmr
BFrPHGPR3yhLK/458EFfFagktlR3QEpwI3zQVAC4inFxkfGkdHWwFOJ+4Zk3J7Ua
CqYjHV90ryzoQSgiv8RdqWidZhy+dS/hf63iDpBJjVZxqZDubAUyIEBkzg98Gcpe
/dTkBn9Vzn4xYJMb3872B2+erxs3VIrfbNo5W78OxDxJpxEUNBJzyXj5ihKDJIRu
Q89BK5o2RaeJXbTq747Lm8hk7jLJaaSiEQjiA1N9KE/cidiZIjcyhADPYr/yrxbv
YqXFSesJY6xJ8Y/Z/POjSENTdsjcHenU9AlPc7Nx0a/LQiS/SUbkHwHEga3P3bzE
gq2LooWQKsEjlm+J3IGlTYbrLp2sajolTp5ks1QaRzVpBuuGK5oZj/jreVewQfk+
aPg2wohvKhjHQI4a0qlR2MX6TAk+ONCr93nep8iMj5BQLSAHHT9WiIYRLH9x0fM4
rKBWI3AdAvmpLIKWzCjtHnEcFnLamrSEN27lHfAuD4+WN1jTErU7OpFLWZaXDspx
LBlZgIp6hHW+5/gRkrYkn7oUWTZZ0CVHpPKLZ6T9cbP0k2ge2X0DhYBZivodsav0
qVfZmnIgV1Y2CumK0mH+Vnuykr0inC+Xa7cJ6wbEnCxiNaUxsfY/PfsH0JHDkd8F
dinswEco9kB6sI1sCC0wNJC8wg4I0pWDNM4Hr4n3tyCJEgAc1XNjE541h1agR80P
kfovw5fX4J6HrssYFV0+TlHzXugUi/J72d30OnEe0phARAGcvphEmOp4E1H3Y6Cn
5Rv4MV8jWXdiHu78zPtF8Aw8KpR/jHSgTig+p8SmEd0U8/bt1vB2EpMT9aO+M6FD
NbPiVMB+02tPi5uoiMWchivNRUxaDl5FMofd0kEHWO8sDFmo0GM56Ad+hHsi738T
vbGdK0mCXt0Zn/XpeUxcNBOs0q2COYPV3lGhRhNEYm1lTWnyaJdvd7PO2SJBI/qJ
/JO2s4lAvoXpcGbxlvh8ylhh4SPXEKFz8mzvsaL7pGDiOfc31/SelSIEhbrVC8oz
kXJx+PnjBsdIu/bJUKpAlF0aztSD/mzgk613gyWXz7hWKieXJbg+jhSowZ63F30J
+q3R0iX03zygoVOwW8KNrO9vX2lORBL0LMky8Un4ot/oqprep8mcqqRyGF8zSM0Y
wzmR4VTX/r2hiZTORrgMRaxEt5wgghKiS8Vj+KXzHTeHM/IRQmgSR5OVTF0z7BEh
k2CUXLJmoI2nllQeFl3md73X3zCFoBER4aaKdMpID0dOFZIYZTPiZT333YUMfg7r
1EGhuosBMQ6qWPLrsFtUTKduy0wUfLKKQB9ZUzsm4kEQ66qzGS/CDHCfFBjPiDG8
O+GNVMXzeV3bnfyFhcWg37LdpiN9idym8hIpBiO7ePWxLqZShJEISKiU7EV+bSHF
8HDczdyKtu20/hYMeWbfCA89V1B7+l3rciq5oH7/t6j7exdhCY9tiYk5c1i8Mbsa
DTJxsFadFnXasCVqAu3XHz6GuR+FcDIV3sdqJsKar3bTZn6L3X931Uhy/DuoA1gS
oUFd6sXVgXC2HE5jkgRL8ni/b2xk7L8As7ljrMrYrRE+j8Unz+vWslMmLt+V1ocV
ER0warRrnuMZlpHgKtUeXkDe5zMFG/fkIOglmcOwykmoIdSxkvnYNYwQVlPNYE7Q
Ql93lKTGk2ygYD6FAo9Ib1VdYWuddGWPjzRqA1W8sd72EQPqIBes2hn+DT91Kd0+
wpdtmYsxFvRdo379/Q4BmZI0h724fnr/sNl37ZM+qf+JvNKvNibBKf3ude0k1p1v
rvaQd7ku0R32vrP80ssonL954d70hDt/3UBEdrb+5qSLWEXqaWql897YG+3dwraf
oyDe1pbbJuPtkC3JfLeMbX1NNy1eAbGpL0wzrbWi7NVn/IjRa5Nav52KZFLcTeQK
t8A7JzWQ2Zvgw9kXhekjrrklYPqkahw5RkYacLaQSXZszCZcqBn+e+X2SA2psD8f
2OwmCTxmkmwCfPZ39gYGxT89hrV3k356dsSave6aQskYUUxvR14eZXPwOZCNxX+e
m/zKlc1USJsssVKMxVQ7PyqbYuabPSqmTSXNDKNYMdXvGpV6He1jVUJ1EBy6gKHo
SsGLeHaPnRUDmGw3H58bXXJsHxgtVIBV1hAlyGhHPl956b1XJgUWT8N1lHlEp5ln
T4twn4Jl7GQGDGO3C/5Tt2RZSd8DzeTFdTaQMqtR+sThwdcdug/XfZWv9BzD9yWN
zTlB63ygKI4xpxSfkCAGgiUzLcBV/+y7B+CY3Yo49gDaIhnuLuALDzRh6Tpymn5H
fKJP4zwSKhc+FnRH0+0bidt3Plz7roGTLZWUX92QCNaZ+JVCkeE5HSfBjm97CId3
Z+IkodXeZK30JSHmKGkYVtLRUaabghM8ZCVUYDKuRWA9heFGUgX78p1pKSstD3c1
eJ1ljyre2M86ReBz/OtYRiYUBtUD88wYCKdiLdlTwk/zIeVni8ipLqQ6rw/O926+
6aKH5krL5KvVIS7TO6NXApp4e7vJyUGM2BfY+QcUTLjrQM62SCpV9cXeQXjM6xOS
YLz+RASv3bk0L8hDHe6/PwyAt8hd9VsYgRnRv2Wq7Kftb7nYzUNArarA04uM9Q1E
ZwNJLVSXhoObLCMD6JBMqeqbBsN0Rukm4rzFGg1q0R7PlJvqOS6UTgKmkJA2NlN7
VOjTKvr0fZP+IFIc2qQdcy9j1NeYk4cuxcatoYNkokrbO4G6bHcpeUV6GsfXegJG
/tKildySGrK8e3ypY+RYhc4ZabOUiUQZYGtGA8cqJM5Yuj0ZTZjQ3s8kkNB61m9i
RVApsjq+XpoGT9uUsAQLMjFdAs10hfwGPoKTui+gBtAztGuWdMZWYxT8LIrBkuq1
9T9QZdWdj1Rk0O6yuNVeawvO+wB0Zz+sM+P/oppdCpGJBCZRMebRRlWplzO9IOHL
vFKmFyblHIuEbzFus1X9JxEgAq+5t4QpXNVD+V07rE5OBfCTSm9htm8CnMG2yr5q
x9JMsIfMI6F28pprCfaxSYK2oBYVR5iD5pW+tncMPA81/t2kdxDQsG3WEddLNT2q
07vSz+L3a8zehqUkq8vgUCfWxhDGcCDlifQTgx8nlEimhJKpw0p03jKDbcisekpm
UVgCd/E9W65qJa5RO92Vc/jU0sYkyvCtphAufw6mJp0+TBJBKf8lcRbjljB8i7ds
OZmi9mDdKAeSyaWIkeXe5UgAyzuwjsNAByWHd1myO52//CiOCrlNm3RVyfv5GGFT
+0M/K+DD5ihbBWS0Pl4holUgeVD3CptZhzJsQYc1YqjCtKxI7NoR98dvKMleGRT/
AmTApFNhhV6sTqBSNSfGJCiSu/u5UwjvRxn//mv4Xsd2zcuxqWlBQtQJTyHgn2Oq
amig/opySIKccG9lxg1TGOf+2Zx5wqabk0H9UMSv5VeIgJzA02bfZ2afCW0Iw1vZ
u8Byj12/Qx8Zv4nFKFELY9p3CYBMp/kcGzkepIIvsR6HTNPHvkO72T6tKv3n049R
Q9bpUrYTfegleilN99IqPcHShDsCYU/Ph6ek6yOy1KAQhQrcqF8+Ep6+yY7/YYvx
ic+ek7TiJYhNRh+QjuZFE5Yddh+CdpzXo7YbDfJAbG7hxrMIcuiypQAQ8yUvDqwI
880xgWSvz3B4MBwqBqv3LcgxnPeJ4c4q+XgHtIx5mLgJKx+iekSv1Gz2HQvHfxy2
SlIyD+9D1i8VTkkynZeSYfucYnt+50znsTznyIlxxt2ttJgfaeH/CY6Bj1dEHQ35
3Zh7Nm8PZ0KO60S6xZo+ehO3KksxvmniS6jihcUi8NFsZuJl0IrEqEp3hTN6B5s8
CFfQyOaoMZtXXrREdIUOyOWATC3RL7HjfUjOTkDf3EBHyg8ASFbd5+QdIPPGrngA
vrnHHhsJ2ePtOhInd1x+JrZHjQWscF+16tDoDTAo1wp1OKyP9YtEbAWRRBtO38Jp
W/DIGZQi/lnAOyBfhpcpjrMTCUfN4jVzRnXb/xzd0QenwKGDvxzXW1nc1LyVaoO1
hxsZ/Ectd0Mp2C88reT7zx4MRcW4eyGDDooV32uXB5tGHc+d65qwfJf0fvopO4zW
0cWzOrj7TzMBN+yiV2kI47Q9BCB7+V1nvo3hRHKBXLgLgJl9zv+ujD3He7ZvJCsS
ATeQwkX9hj2mIApTuK5mgz61gTOdbwTXxQhL+0h7zkk52Pd3zV96R2ozYP1eNKKm
1h5D18uSJ6EMbP5gm4q84u51zYMOaV4dHHIhQ+XSp09yfINoKmeD+V+PMVsqyiBq
vlFVpt5qXSDdBeRDX1whqh1Nh+V+J87hR7jve+GT4P69D1WIcOyN1uT3XiTVIvQA
VF+pSNWhRDrh+v6QVBDPZcYSIHKBoFztXZIRRVc0E5O/fdsf890N5imdmC2otVzp
/gTTMKuGtaI5kFyPWipenjZEjZODzddHth97GomA0qaor2zTInTSxaQgwaByMvd6
cXhPHtYdDsnpjOnWndXaa7G050A7NrB02Q52BORb8fLSrHJCZEmDtbpKUSjzqwWB
nhWOTqsb5Ad77fM8gcTD1w8CmOIpdf2yAeF8sfXPrPCHw2AycpstQrwMBb1euJTz
80aKNt4AbV+2LR/zfzXMLSWNwh3Qiqy23J83kgLqebI70gbHfCYxf1UOc96r8wFm
dn6p+9Rr/o3twivSuvC0uK3Bqh4a7ZWvVk9TUIgdDDu6n6UZQdt5PLtVw2DFge4y
gHmCDqKq10frqMnTNbz3Lsc5jQPXjqpfr/eTl2sM2HSKpIseelzHtQZ113nYi8Tx
QYE+E2zpIvoebRpdljkatdxG0yM0Rm/IDoC9BlGuQ8znQYQFpenZlhQxEs16OThd
rTbQObc9kbTnaxTbDr9QrtqLBPcDyjcBjg/0wGerT/Uj8rtCpkQEZ2/ytkrqelIN
fLccKZMqEIQi6GA7/c28+gwEaEHSib6+PVJaPWtolHZijCXOZaqWcTiqk5NU8vsd
vUTwQCM8DR6Gk1Syzlro/8eOS26myP6ec0aPL6MEA6CNUDvAumrEIuIhbJbf9SBP
4mchXYloNTcGrkElKU7JHslXpI863vAZNG6ffKC7PFmrxh5QNX5UXguc75gH/5tP
ZSYm9bt59k55CVUkrerlK+MsYh+6/5t/fSGY0kiRUUmOFr4yjX419J0nZvByEh3h
xu4C/HzSXBKI9LDrl73/y4GjSiPqjnHOtLjOtI1wRsJnXz7tk0TerGlpfFBX7IX+
fUqSnIavG2kdJ/cZxVWMqESX7MoKC0KrvHRb+4Rj/J2WxuITS9zwGOSjkRHs/ht6
Rzs4n9i2vF1mtnAyIjtjQlkZveYSpdsgJQX4kzXvu/p5N60UxQ3hl6DEEAAGKRCx
3XPgD5IrWo9LU90dwrYjg1Clg0a/Mf1UkUHq0/9TOrJyIq+QEU4PyV0EskVyC3ZZ
UAGakDCFx7UPTjqgp36s+e/gHvBfp6E9nMitSSdCGWFkmH0gWvtP5B9OBgE0bqky
+UAQPSoJtql18gfda9HRGbHh31+5u4kPukqD9JnBiXK0oUUd+q6X/eoI5UdZtDaa
6b4LU5WXm9RPovDIK7F6nEkpNzhsBohlNoyqLG2/JcF4ly8uMpYlbzRR/UBjxZZf
EKRmpSCDHK4XFO3NK29AtFy3/TJiUeDvp9V6JzdbnmM9HYaALHoWUEI25qt/d9hX
yTTlaEn6/5C16EOjJSW/i00mor3db9PEwytH3SW2ZFgCil7emWhdVC+DPe3BJ+f8
g7g5OVf57j+ZkMZbM/2kKLprm7Xe5xvoX9BiCJrwESaAQrmQsDsqinyTT8IuhEXM
3FLU11n3d54JZt5kZQAEoFsCs8b0PdCYsSFsV8/f8hVR5yo80KJ0rIHYNI03P838
DjRwsrZalPGzwIEUXv2Loz2NDaHy19xMW8XKBq2/6jA0IcpWj43U+EBF34lOxdnQ
p4c9pTSiPkqpF6e6UqOq95VfQCeUIjzP5aNQu2Tdoyi9LtpINc7v1K2NAqihcaNa
Boa74K+v6lorv7B0VIboaTNq96gYcG5TXVB8/dHo7UC4Ir6oog3YZ4ZxZM5KWRmf
GNNDuQQ1lq62uv9fkF+CX1UyTi85+iy60uwXb1jjsrw7FJqrEo/uYkO+gRfb9zW/
fgC37t+VKPwNGHEqAm5ZlH+HhcHz8SZMHpbGZx+ondcxFv6FIRsPZ9cTB7iZIcp2
tjd3TRlQXPGd5S/N0hEhlykT9qvEctwKyMdpBumTpdh0fPkKelb/65CEc1EtPQkA
6t4PXbK/hzD4SOYFCphIWdqqENQMTWBbdJmHBnQ8gBQ2KlVEiBvgMO3EcxbNH2GN
jaWe7VyH53dsRls3s5iv53SCbfTSgfqyB3PVFiMpbqF93lXB55TGPIty+b15qTxk
ZGBLdhyeVDhbIyUjinyCILgB9Iv577cXCtVadqjLW6U3ZyE5zuy/q2Z1ppnj6PPY
p0tkQh1ilGbLFAGXRO/LSTvVRNDDJNwf7glPaUFOY5EwYQaRfMNvGXKmfY77ABgb
GodEjLSfgC6s/9oNifZv5yoyGwW1BXpn+X5Mey/evAfqsUwO+q9AOBzSFjO0sY1K
S1ZfDbfv6I/orG3ur4RqGrTMv28eXACLq/x4vN5HvJmZGrHhFOlw3Aehgzn6+KE1
6VmKiBaf85DjY/8SAXrtafk65smi5Fyn8jgySX5WCzBFYcZ5hfgv19L4jLpWtaAJ
hsQt6IabBIW4hbYsVGMjMGZe4YoS14kaERKqXDeiqk4JNsS+MGQbX8m69012EPqN
ssbp72xkvyYF2FRy5UvJB4Bpvm1K8HtdwrP0JPXoKgZj7TDAwHzlz8T75O05ggyB
fXhKlzhJfOax5I7K/ZweHzKFF8sUg52AFXXwHJ3Kg3tHSVYbL5Yh2HqjbULecsYx
O8cREyfxCdKURmRbSN/7XvepNr6pbQfWUfmjgUWffR4XwgdaLL4iqNBEi8mldf7R
hAc4o555M+S0Q0qh8ROQ302W+DTvv4APR0DjK1SLEZ4ufDHQoPb2QNeFwyRTLxjf
V2XsT0cCY6WkC4o1RDwvFH4DsLIfRNhXA5A7YkzWyEaBEOa8s8qhK150XFEDPstZ
NUzaq3/svj+XzObfi7YK/GxP8yREnG530FLZnODVDXxDjvBwcwJQJdeNgUc0Srg7
FaK8XC0/E8bDwJ67UjB+JA3YyXe152dASgGZ0Y/KYcU6vt4VIh5/fgQ48Dq5P0Jq
6o8xf0GCRhSShxdKMGnkVG7N6PaoxfQHHAirWcvpGn+2emdDYupTc3ms5IpC01uQ
+NQi8N8N4al4gX+fsHrbbA/b27on0tJM+htXOu+/3YRjKOXaMd26vQ+T8Zhya3Ob
uL39pre4ftNmt5TN/1lfjLQL2p6eLIDr+KbtHTuRYwAn2XLEzpHX3iT9vzi44a5a
Brn8H6x4fqDeSQ3DwhJGEnIc7VDIYD1pf5lu3c/MiZGqfRDZj6knYOX2NiBOsM8t
MVp5ZCkjDoExQ7+uNqdF7z/xGylkLwSOLXKnH4vMQ5PzMeHVriYlSMn2gqigexve
Q5gR0N99L+LgaJEuG7PXHd/x2usF/S3tcvD6ZAiz9NqVabN+ZJ6GFqf++N04cqRD
eYiNPuFqD0u8equRh2LwnuJCFzgl2tWZhr39qHtmabiujZ2Jv8WR8XFWtoJPmcNW
290ArnixpzETDia1ONsMVDYqJYRvepl3NbYS+L5jjGB/yrb+tZohGIrgPbDTx23l
A8zmHC9GpM3unZBVs4etTaAubQAMNtCk2lpjJB+s8mZD2c5egSRYLaqTKVvdqltO
H9x1kRTHf2+ETLdsr797WLFuY1dUyOwe1NPe9NhVhPDexJzTXQfxWLGzq0bB9Y0l
H7bwj7FFBH9OCoPKpSfedrdtabDs7lYB5uxRYy8JRZLmRz9h058AbT19A9sgo+1b
u+VrOR1+hXjMIVp1cC9jkrs8QRps9HX3kXTKApkHqCf7rGwxd3fMmTL49PWOXDmh
fgEuAR++K4K7lp77iVzRvBdy6o+c4toOd+12KeqgTdcuwNjWIl83n3v7JcvJfD7T
/RGKy1NT1CKyOv9P71zhNYSUc60+wdmiMxONRUTDBQnyvIIpqp3w6OZPx6JiIeXs
vtfAV9xTisvzE4uHKsTfy+Rf/b/Ju5G2fBmMPKM9cYp5yvnfNOr1pEacZaXVP4sC
DfCB6HlTUix7dHURj2M17s5uGaV3MEfbx436KOj524jNEGPIFJ1wXMjn5VhN9ev5
lLGBbCti6mKA+UmkZbj1KDW92xEhXZhKczBpA7bWahkIVBclVyCwtX5+Em4L7mNg
DQS9sUcPukW6ojI5Ng1s3cmWit8pWO3M+GZPBPwRUtCj9hnD3De3GhLSf13zQ0pP
zMpfjfF440eyA9C7k80uPisQUStHyg4nVizPvGFuGPQvvRpkEdM/QGnRt3bVMLgO
18GYtS0ClH9yNpFj8iQBHJSU6UJS3Cui9tGzVU7wuNLVW06C0w2FImyNm0hGks/K
SvmK+2P8LOyH6gJctRa5Y26iMNlVQEntB6HjdpQB+Us+pKJLfJkpvPK3E0zdSvGr
PfSgbF8+ISEKgJFEFdj8pTPBKSz/pFqvb8usRM/3CapGOv5DXDnlv49M3MTwf66+
9HtFyXO4+ODDdLaheFOcAluDGTwz0Sii05BflJfYC7UuBeNFTMjDCKIwvOiB8Q9g
antoWgdd5CK2+Pa5wTAYkldwQpP5drzkKpCXz+WK2913hmqIWYhrqr9xGUujGMH6
OBnqV8Iic5/xhk6edijWYspRpgGojD/mBL+raPpM4s0VaglVktcd5fEGIhDltAyT
2MpMyAb5uTF/odF6THLwgE5UPO7myjnCIoqkYwf/cdZTe26B0bYUC5BtGoMWVxCc
UQWn9BTulfFHmK4BOzJyNnwlYu44+6+f7hPOBzAMHj/uCIWp67gA2oPjsF2otp4d
gB7EHZ4aiaJc+MaRUsJO9layLrjODmTGcgAxFuL/VMzvDiGOPvsGIQD4+oeZjlZ8
gluA/Sl6jZ4hFwhYXlZaiwi5LnBlUGGDhz9qNC2TQj5rIINyd9hUTICwnguHyv76
tEJ1vjiSct7RW/ohxgVwnvnxYilW952KxpUd7y2dlSYzbp7N0tl904UvL9WjZxTC
zAm2r0Lbzcr+gD1CF/p7FV3ybzA50oapwIHR7CgBKdljqM3Bj4V3uDXwkyICggTA
hkdoRa8QS2EHy4zRXtSK3qoZgLMbD/skD6IZ+tbNJVL6y6uzHuWOCsEQCjOMmsco
CsvwNYMwvJ62RgIJja0mo5mCyzkoMbH2YTKEtC2kN2520lRcB7YeS7PCArQsqkCJ
IKJ1TYuuMtBzZxyVrppXpjvnmjmdowVutrC0+Ud8iz7gdfDVmAzCYadkAgl094cP
tQgekJUx3AV6DO3y46YL1HV8Qw0nIdicyalqaySaXdfxhwi5HDQxbiWl/tjCAScl
nrYGCghkZe6qF/pMJZxrxg1KkuTdCIfIm3GNxqX8nc58AOUfF+KxhurdcXaPOX7S
Ob3m6i13xaxZuB1Xo1g1Jysfdy7qoaj3BMp1YfLIpOZ+CpOrfauDY6LIgG77BOUX
/5hlT3dHHHzIV3ONEpHW6gTvMuiHsiRu2lYTcA8n+IlQoLQXTcaS4gjLR1PCQZrb
jakcpiQaPnpLPy7I61L86I//Vpb13UkLJZC5xlPJLETgF6bAFcR+oGzvBpuByAfZ
9htLZFhxfy4wCGDAq2uBE5gAAIw7tmDSJSugb2+omGL9pLZBRrkmh9yi5FfBAXPF
/r1hPbdVcZ5EoO0f5dL3WHoVwSsN+Dtkyu2fNiIqoN7Ok7rR/XxbQHZfmQIaqKVG
dBhqsG97M7Rl1AV37yZXmxQy/nM/QrxpHkX8DUQlKnEqX3+1GBggsB3d04mArosw
GUT8UB6lfOmUeYXP1OF/TSoUVXPdEBdIHtrr+28Y4pnARR4jpetIayMJeqs4J3zH
ymHjXpXQmOR3Q2L06ZLFD3wpXR7UqzhLcR1zFKarNrMCvoQmj2SYjGBya6zWjZEs
fpZS//bcZUr2mwclYmU5UyQdmeWEczP1cAq42GrLuGCu8M2ao7/AKhQ6P0eY5V5x
M+nVRcSL69Vk28SNZ6x4ixt9oRd1VSvYO0WIzqGr/rHe3/dJ48TuOqrfGPLUbygG
/kFvsbukVT/tVWwGLHEJ+ESEIZNV9cHkSCw6SgaV2nYaKDQOFEc8241NkNX4cCwz
yfpvWkTn5ZAQ6pkodVsUybp8L45Z3UVY+gUez4KYOqMxDdbz4R+Sjyp2pgygc957
YCNW553XHct0Sr1cEa/04GtXN/QLBH5eVbXbPf4lRXQ/FQwGg9CezDnaD+BF6+dv
gIUAo25et+Gp/4uQBHUhAfZPMgMlPIzLHxM9cbM0EyCV4MhIY7LNSFhW/lEKtf48
AVEQMIpYkKhedpZmpUEq7nFbxo4qkcTmbGIhMqyAU+5H6jVXshLysN6Nm3pkOpDf
iJ9+4XrZjHccl0+YnmztwGKMp3vxr9Sp5lHQwtqjZI85qiGxp0KRup0yTkEWe8l4
1XO8nP3kWi0/D0u7UNEb7brCzwUb4rpMYPc33WAt5098stf9oReyMd1lTSU4m9LZ
WNGM59AKkmDZ13Uu4DPWWz77e9eVXjtuzc4hfKNicHaG5IbSgpqUR2RVE+GZdEzJ
vZQrRrWdWCBwHw1eN356wRceL3fmiZUXlYnAdkpszsGIlC9XGQ2MqGFrWfAdGTfq
3lb4y8wo/AVu5R/RXdrCtB5X9QfOPw7fVGKHCBAiXeQ+o1PgDgC+N0+hbUqIvmFt
Kzm5dLkCUW73CehY4bNzVrDN0AQkJ88O8eJg/JKH3QYblpcV3Re3W2PXh4vlcGET
I88NM/IKIs4zwoSKITRYosGeyw3jvICGoTNE/ux/fuefAG2DDJ+Qbg7ovha9oNvU
c6BkSQrgephLZYQ/R2F6JlI2b1NKBXunMs55oKqQggQT42Rdg8HWDDNjDREepxN/
+Rua1lT3HXRxOnEw0mc3LfLYO3DVlVwJOTgG0HYE/hRxANfloARKPRN8eGXsDQ4O
FTxrOId4TofnmgKqvqsm4XfuPOYcNPgMdT1Cjtt6XwQlJtiYjGHvvNvaHHjyUGPF
3B91Vn3bmZlrK323JeBlaWTqDj5lNTkdn3N9F1G5WZ6IsURS/4Dits6DWyXYPgpf
nDzSu8Ilh2O0tnnyP4m2QVyAAc2iklN5ek+9L3p0cXFOLoDjvPDrxfYLFdXtHhI6
TmwKY+ekHXeuvg11xy2jfKaCKQ8Hc3KOINJ0o9BDUCx2tfC/g+l73WCGLMd1BPdA
pH9lQUzjGx8+wgFdssrnxZPyTPBy2ymf1Umr3wVfpVulSu0EHNAixfHIbNOVMxCs
On06OMDDqteGFn1FZCLXdird+zh1v6jLSuX2oa3WSU5IFnji4Lcmf0gTCo2tNhCF
Pv061KRuYxoUMNoXHecTHcPjS7HZJRHJbhgPzkkRlwDxEnGqGn+XgKNqXzehGWDq
uMXbeN7xv+dhphuWB49DSy/J81LNwE09OhwopNyV35/WIneZ6NafVvv7dEj8Ur2e
v5Z7XmlqlF3vAaNygGxweHoA7LwUB89ES/LYbfZv2WHfzGNheTg0bQ/HpdEvO0Yp
Vi89d8CPr9A+rstSAF2gS5YmmQBCk1ufyLOyaqedbZv1P/8UqTwUCBRSO0jTXBgW
2dLZA8pTUdCc/MMlGf/dUjFQQlMXrax/feGjyv8eSpqX5LBAodMD4VKR+n4uH4k0
20OEzK9Vdw7661ocyPkEhuE1nMTrDN8b9gcDiOMRuMLSdv31ydin4E9Nx9H8j/R/
l0Drx1I1lBy1Kms+BWhRc2lEt3aBo8URxi4zS4WBX54WabS8QSsyr0u94OjiwxLe
HKVHN2blzunFLEJdCa8/26Dy+CbR4jmoWNND3GdP/XL2kac2e2KahZzj8eNY2cDu
/rpxkEEDlAo79ceHJhCiIndJcUmFBbLiGOOc88E8tytVqdTlI+/nMbdKGjHEyXId
Oqj05yqvgxNh2Zgh4+maIVFE1iA6op28gTDpAurfhWcvz+Kh5y37vEn9ivYKRblM
rtEms8rT9V1THXqwQN4UKzz8q7NKHU4fAXCHkBL6LlCYMVwee3bDVP7KFshEZfV9
vEGzS0L+lhnHXJzOq9GOTHAZhGB+qve5NvmcewcWpbYb32c9+2gMRCjzvsQNzfE2
rZiioxU+m4OIPd4e5QLWb6lLzGOIX1yREylp5ENZlV0KRTxNZVfz/9Qcm4tkgwnz
2CG37Xna6+j0K1CwQbKbd/Y8P39Y4KdZrzEgEBRwwZt3KZcRE0MkbGSxUZFSPbWn
G5iKdHCztPve6AoBWE2I2/mjpn97XOQxRgqs9b/vuGWprbM9dPjmb8UHvYPhqiay
G/QM9O7K4Qrp6W3kFGlqDYtwzKF7hVtKWepOK5RZNNiMNv2QsydxtJAMBJazRyPL
DXmP4CjY7/jd8rHdUSweRedITE7CCqxsCf+yrLTMh0nQSfmrnfUeJttW1eoeMpwU
CYNUNx80sDdDNYGaihEIOvN8gvXm7dx5X82cPzIhe94u9sZ3VkfZIqpCWaw7TgkR
lOWSkVh8T/mrocHrU+jaM0Zu2sJcLAPC0gOZRRnlvUFqy9jQCKbjuYiKigc/14pD
PdKJz6LLOf/fcQ+S1uqniQ+5lAvpANcf2fSg24lH5qVqWh1YQ5sS34d4BXhCzaVY
ZrByV8S1p83iKs/Pb8pSnBlNG5wET5sMwViabTJHYDarNVa8FXvaiOsU8rKoXEUZ
Z6zSJDFinKy8CsfTzlv6BHKSbyiXKq5ir7VGqxGIE1Tp3MOTMClw2aXqKx+d0Pd7
wmxC87HjqnFNPEzvq3wFkCk0lRLNbdCGHWq1zG+KM3TxSPFMEE2xNKHveiy8t4Ui
brR2Iq/dm3LCmQNPrwE0v9idrcZp6wDklchyedjVVkCGv+dETRdaORKuV1C1MJd6
a/0BL0XPKmb20pUpc16LOoqz+iZYUAbcFSJlUjjNMDi0uxm+MfxmS5afjdB9CbsI
K6limB4hKygA8ex+gHfG0ofV5RidvVmIiz3NBSnqq/aN+Ld/YquWJnM09tfr42eM
r6BzBpWjQyg0hyX5ZHBVrALBuSFB0NhosH0eOZJO7Fk7yp/7iOLFUY4GRwSnj1gq
mQDJiAIhp06Tf1qgCfmrkufk7mCcnpxlUS6VjGGR0kf1Pz8mjjXFijL5ZrDBsdZY
IQEPOhiEtQMcYXyHyO3vM4IcivR3xVvq5pxurHY0xnWSbewtA1FpvOoAO4gynBw4
lgAIPwyMqI2O8FP/WUn1kcXsttFr2TUAGUqVQRhxCNVxniaGjGJiY7nVc+59z7W1
H3gkw4oCT3VwXd0PBd33PWQHgDa+WSSFGGfXfXnqNzBRhf1iMLSE2kh2kN3QQpjj
dEzlhO54mWKAAayHUYOuTZyLOPvnPAjWanzCMjN4oyLO+rJ1jRmr+DbnK8ieHJPV
RuAA+KlVbJ192en6V2chvgwE8zR5hU6MRodj4PZMsvCnDCxYzfSiez+RDoLWVvyj
Q3B0qddReZESiYjDLjXCLbFZkznMyh00STdXdic8IPnwB2xBrsN55RBd10M7EKUn
cDykZke9j2YUZ+ffm+8l5tqS43hFfhtGvV/nVAmeMW2Uz3ewANzrM2KFq5IfhkIB
zSBOrZWggJMqUbJI8JoXNBvJxcZWF44Q8SF9yQpkOb9kS4fpGHdjui4uT+43slb8
EH6DAnSdY4bifOSJiYalHCeR7wnPnMHscIGG8pCQhv+CPiR5GeSMLRUOB3omWNow
IVfYt/SsdpdNGAn/lbvHvcHYLQhmJz1CtWkFdxPa9cMsIlasfbMKWVHFCNQ/D9Ta
iPy173lq4y/+nGS1lKwGVowFElQYnHcI7RUNVOZy1shjSN80FQ+eMgI0GYUoadxc
XgWxLQ9h4i+V9L6+sLoXML1jK15nidXVKFe0RCAoDaSfalzZdlB2ADEoJAsaAAxp
70h4hATd6bqgGq2otZdIR2YzE1brJh4Bj1s+vC7MikpNe8cQzbgal7cMHHrGrXD8
Z5kRgiaB7vUVi8k9WHdXa/ZhhTGkVhaAbEk+Bllb5TfU0hf4lvzJu7aSvewAV50n
wBdGEWgEn9hHOguLuKCr+sxaUkqIFD34CzZNa7Yu+5Gw+nY2m4rXx0pQfqA/fH5X
akI5zhFhcn1OONY8O5rNO2IJVoPE7MCKJ87yeiNUtAMBxk4X8ct8RD5gCKy2Zc+V
cvn/dCRgKzWfFZIfhpgpJMPo2d6O7cW2cbBdWjnfz3larE2tLbHbqDSjR/ZgvRBS
ObwizFrGM+wgtvBkhCNG6ngHhiaF92kBrZBr9ZWATEDS+4TarH6OSEjCHjHFJVDv
keXk+zzhGol7rLLzvpNjWd0ftmPGIntQ2Vp5mWnEIfBEkSUqBkX1Zw0LSPciU/Vf
wolRPcK/NN9BtgMYuFmLb2YTNjsATmqfFksbxLSNeVdAl+lOO+XLqEY7KCN91JR1
zxCEmtdsOciIjdBth1H4obo7MuQwzskAE0Etw6sDgjpTkotjILE0twtKIT7QmboY
rghAVA878mJyKxOYM2hLYAxO4VtRItgdHJyUHFyjEd76s54S2ixRfvx4HtCA/yR7
wDdKZN61Nr3i8SnHZTy50LqJTBtuxWU3cQqyEfqUFJHdz4IP6Lln5/ZywgIeOY9x
33t8P6mrf+EAPrnJwSGI36R+cQr9hVshXxz48+xgVfyRjU/0a+bpG3vQEU10kqfl
ytwLhMXil9REHjdLql6JNWX6bAt745YEqsN44cacb2grjK4QSoBASH53/vZQ78jb
sMBRAjkiwtEvZpPfApRfiwb7fDk0aF49mZBWo9qDO+mC6uybewzJ2bHmneZkD+og
Z6BxrpFykZqhMPtkb7gYhZj4UGz7ptqXddTDyMLNi1exGV/smQZuOor2nMaumKSO
q5luyGFCUp8DjEnMABtZzZWThZYB75ctur9XIYu8Bm7V1suUJTjDZ8uRqq58tgWV
4zJw4+sTd4ChoeDaV2bQbsfv16/Ez+rN7mL83tlvx0lVPIodNd8RicSayk898Sgu
w+hcfkljTrUz0b+R/vXPj+9ERPbBHFrieWjvMak3m4BdDng461LUhsPQ1lNp33Kg
In12NysEIh3ZJFm84jwHCQWorgQhKm/8wCVp7bgq6qcAcoPNpb3ETFYY6GmxJl47
0SaJ8FPvIJu9sSlVof7ZMLfjqLM7DHNT5PbAic5ucdyF8GiPnZNJtlpkHTnt1Tp/
UbUxXxj6sTDMidzJtoqKWY1ljmDpjGVG8m/r53boQaZ1CV2N+0aeV8Fm/VCBJWw0
pw1k5kSavtsgPkZZhyHj6z6dDRgqiq4wjZEjN3X6JBOVU1lF5splex9cn1LhyU3x
0rww/RNkv4u0QjDd5oaaIAOWu7MkQNDlwGOML1IV9Bw3paa4eZ80+C/DEdQmMETi
ZJM3xZugmW4h5gWPzBLXu6AnXJP4YOtQuy+z0JCOMCkxsSvaKRCoU3Sn+q6YqtZA
0RiCEqMyIgbMBQ2Yp8B4yqoE48Y0mS6z94Gi5EPuP3vdMfRZsdVHDq2AUB3ktTfj
+ptyGqshJQ6TvdU1iXtoki3i/4M6dfe3lLLg7chYrWbeYkw3n8F4mXfwMYLZnrrT
F295WNF9aho9yUGF/+Gg7KTenD7+Hpy6gjyXv3WfdFT0HZsToOjnJk/vFFZDkpJp
lNRMsZUPgpH2rSP4Y9NCH6vT5p4IGbY1LhvLLpSdAJ/s4ZDauM1JM8dTzAlVQfHv
7WZC0QlnZWl+1p44HHYRn12PEL4JFMsYvjISQx49hj9I9voMfnGCM1UMAHFQ4Mti
F3Uxs1kcfBucguYbjMSwxWDp/BA6qCewCG+blh7FSduN2IMeUVmxUlek+WeJGTO5
5odZ6qOEqVYV3iLjQCtCTmRq48r9uKpz+/FELcmruIVT2hKcL55J6ojxoJCp23pO
zj+KRkGSC+/tPiEBwqVe3BY7+nao4dAk9PSFgBymfOoZTUQTphMzMry8oOyGfgX8
4ia9Wu+atXGb7ms3rTpDK2JFewSMmEjZYmDMiMUl3t9nXsL5i9qMYxpL3oEu57UA
HTCHJeBOl0nGVn69KnH2aTDZIQokdlYeJXMfYPeRYWKt7wby/ha9Gp6BuXeYL4jI
eVA5tO0kNnbl6mcJbPM1xwK3vgsDEBMN/w8AmlHG+ZZ64TCzufCzjQorttGbWgXu
JOXMoORIif0EeTFdmG9/mZE4aW+EagBgkWvsyjGS0FBW0S957E09rUkYGCEU2M7D
lwfwHvtUa75yo5k+I8SE1/dRm7+ck6EXPW/cXT8WUwC/AEYYtQ/tOqWZKWWs/PQj
7+nKRO2nugZteseb8HbyQRJVQ+RMTr8rm1W7Qkd2Y8VHHiw9gNo0zUCK90+rzhYU
ub8B9Wo412N/fa+2aCwCxnMg3VSn5xalwwlQel6PcRlhWV3k5e0MRvH5fzZ8hjSG
7GcKrL/HqgsH5MuQ1O/o+VaBdWf2vt6LUNhNrTJkqQSm5LYEsLD3Lje3UV2eRetk
4AoTrqLTTRile8p2+1QIChixQp+aVRuzD+cwWCw9h0ph4vd+Zxrv4pcPkQX/SG6c
9aS9923J611pCr6eLW3o1nufkKY5G1kIrlsV/dg/R0cmZ7bKurqjCiZcQR3IVene
X/XXmYi4ay5rpTsjAlB5lFFgR8SbloiVMdcghYDd5bNsZmhdZHcsv2vQpkGL9m+Q
EWzbNmb3jnUPwyBOSacObskzmX0DOq7mbFJ6OYh0ucLb8tBlfPRvBdSb3feZSOna
Zfl3Vh3PQ+hvHG3DZ8wB3Hn2bNbyiCWLDhPXA7fh/W/GSC6B7eyE0SzxH9Sf1RPO
KvTt5v04KHZjpVNb7G2bQx4jXPMxBLpEzCh/LdtSdpKSs/i9pmRZX61LSB30LmMb
GyUjWC8L5Lj25wlbUup+Qq3MxqifpmROSMQVmixOFC38YNGDObjNlG7mcUVPq5v/
IA2iP7+uuNABirJDj1eCBUtafYM7gVuwE54rsxFh/4ivFkCFKEWaVNFOzSPhYmfR
zK0LocZhM65rfNJwMC6pyR1Q0lCGr3d4u/F6jfScPkLFF4BNPeTQ7zqlSWbJksOs
zq3d5hXtXWdptaXfoeMVQrRKVKIeanml822OBM99jq+e0FX61/3kXYHkjY9Fh0Uo
LRVT7idAXAFDrD2vc0IguzWyDbmXLJAG1S6GZhDBLDcaWoiBZe5rM86r27tMz4YT
lp0M66alCjcqBOPU/4KtpB9VDn84SdeEajYWDVHwrtUkxUH4NfJnDA2Q3rDBBlwc
dAWGGhnjtOOENPpPX3TKBgauZUrd4YeszniqzARUlvm0rt+NZCZe4+7rK+SKcKfi
o84tqNZW2psyjjnEEPlHhFzBY16OcWTttTV/iCqDzUVgHRADrFjpB9At137uq0tw
tcACy/U68QYEI4d96+YkkUgn6p2IouLO8lvNqLP17TWCCKgocJHdbsxkVgrzt6z8
C02HYXEmasGxKnLF84+x6u4j5sRE8b3kip20Dgt9vfPJxxLPirsOFt5Fsfkn8f2Q
so8V4acB7pfDvLho/IMrARi5Aj5LF2TAYe3ISsKNjVNKb2awyahnsHtZ30ygaGfm
ternFj4EGyGaut19Vx4wcP4N44eM+raW0lUnsHKoN8i3N2nAJ0QKdmTmy466b0wj
myAx1VdpBv7nUwgfwOKUccbjk/ButARfHmuNlgNZ6fJ8EwyA86+2TioRAdatjRJC
5gZD+9J8kDz5JqRL4VmD2uOSlRpLCtKoTwZnVASovINb7yUluckN8K70aA3MPLkN
74qY2pgasHQi7LtS6Tv6Wl/aS5o4ot2Q9KQTy2Qp1H2wXrZaS2MCgyWpwJtdRM2u
hGFndKXpLBvGHSSFMZ1ex3j4/ArLHI8fZ9cCLG1cWCxq8oEzF43wB01ZJNlExqFR
y28sSJUbvZALXc+2d05/+7n9vLdXfsenAoVLZjwq/z9D3n4tNjWZFcLSm3k51V3u
WQjGmDp5DfJf0aAqtDl0zbAHDTXxk/W9aYRt3A5ZxsepnuVy6WRkwhIJBCAl522E
Wsvd7DdmlfRkQXuif/4ynuqwdc709wHAndnnYDV23PjFgFgYi5YeCmCSefBWw00w
sx2nOfob5YqkWzKtNhOvbcx5IK+OZJ66AetKMpiF62xXPhyvuDjflvTrsE6057bB
/AcebnL3pIAj55JoWP/0CTq1DJB15BWzOVpiZJ3oUMc0l3jNnb9iVpEepq9dJAC4
PbSgXVP8FWC65e2uQRanx1M1Oa1KfdvXokWm7SoLdWZEfuxPKrbHZnJWvYMorunH
KpCeAllSfR1+EGfr5/HBJvvk5F4i7z4dDQolANtfOeTVHeCyWtRYPS7jPoEV3Ixv
s4aKgWgc24b6+353RJcovlp39W8umjKjbm8oCgBDbP994GVu7f+smk4ws+12Rfq3
r4gf+7gnTvTWfV/DHO2nKU1EVW6vTd+OUXuT/tY2vZGO56koUGhEz2wlj06mVrPM
nluwKkAkNk16V/rYax4FbqMpokud+eJsidXrznIIQhRCgJTJTQsSCuybMNu9sZRs
asfiT+kWSnh2bW41IfW/o0Y1UCGJEiQH5AB4BqgiVImZA/l7mwsotVfC84pRp4vw
XEH0wbGhCkS8LqmvZBGCuBXCxa1hUz2L0HnL5DxnfBLTt/SPVicLwVBv4mbQ4lL3
iUbA1BfSDYEAaPGMuL5V0JYU3VsUku879sN/7J1OUnDyJhJR+GxlaBdC/arKJeLs
8JcDruFyEGjNZxgXmJvbnwVlzhis9MeGBWrd7ju2SxYC/F4ToU2IxzN+3jQQ8bN9
Pz7TAE895zZLz89uw7HsEm7HuPVOcnhTix37MU1Mm3Bl4Oj4G2KslWunR/XB4Jsx
b4+8AZHOmMreY0aYH+bO2djwhlSPIWXbQes1EVK0Ky38gAdFYlo/ZohSZb5Az395
SM+IRdPxB6l4dDaxm7iK3y10sN/K74pUAZ0/S1/msFTplqsTvSokUWWTYebGRRly
IExKY2gPpiJtBPZZRxjGPrsag1d/EqH2u+NVg4LRz5eXVm2JbK/SKXcUA6UCi6To
sijp5+1K/ehKTVgXCXK5B0w4akRjvwfqHBmFdl7klyk3UbZvuULEPuHx+UCm0PPa
Z0GOPByqpFcIc4HYPlJghx9DlVOIbatqdePChzLrUpSpcptJEEkIgUfL3l3cxPSi
bGkz28gG9tMBgFEQDzXBDmI/xYBlPOqgPB/SKQTs9k8jgPeq27YwWLaR2k40sp4C
RySrHiZ0xiImChnDTkv3fkq3ICn0JxUFX1BeFbGp38fQf61iAXDv7gycO9K04mmb
BxdA/ikYMVcUR5X/JK4PhkhTJlf+a0+BiZ31tZ7INytM/9T3BvgB56xSfaftN82I
hcssJuSKQU5IptLpQT4tuqRsIl1WjniqX8objHUxai+9ObkJC6+rOVNb42VlvLC5
PQyH8iofvco8VBgfMxaE0dpa2EbkIoZdze1Z7rQjoUfCSWJyeFxvLS/xaNiOx8lL
pwH7axQORKiZYYC1qdU5AGwObRSzcVtmGHEei3nHz+CoJ+Rz+BmemZ2qSBfNaCjP
SU3ZIxOCZ74boLiP1MyTCk8ADzWJeNug3x6vin2bUCem3QT1W6XJ3KXkswYPUIKp
2Fc+J0f81kpSvOG/izyGpqOFDx3e9qd18qy4YXYSlp9OfW48RpA87t3vlVVYgyEu
W6c5wukIRmCwwQvkqliCHQyii+Qjg93PpXnIcHBHHnjqv0osyWacUt2KJxWSB4rn
Tei6rVTEeFE7R9jezwrcKv+W4qAPs4pfX4zRLzQmTC/pvsj+IJPY3y6YuL81ahVK
R+Ut3jB+5Qtso6i6e6Q5bUV8Gds1tscXN7AdPYMfnQmoxp94/5Udcmqn+/+wx9h4
zwI1os4awqsM0STduGeaCfGpDzbDZODnLjaSQBZEp8mgAtuzGVE7OsQLQ/zDLGZZ
+Vl0Z6QQmkpLoTp5jVIFw2Tft9V7QT5slkhxS+DdLqTGpRsVrL6YnY/ySK5q9eti
3HxPUw2abLfWLnCcROV3XNlvq3LkqQOwRVcbxAv009roGpnM7tsFx2XJsGHUp2/i
QPNqQ0gTUXFCiPdIBP7Vm0ROr4HGzFTbyROQLNuYS6cCiJ2M4hPT9MebAkQvm5Mw
Krq0NHF+0t4o+cv3jckEIojUKIL7zjz7dGkWauWg4CKKWCJTJFquG18BmOjyDru6
UdRHNCJK+g0QReuM+oSFY9zKR2C0BwLBbghe7Y6mhF4iXgI5eaK/8sYBLeBphwNy
9xl6wVgg5Mj7ibgffRfOzK9xvTmcX5K4KMuKmhM+2UddKXioMC/B4q3GhiuPCpLI
jqoqS08XMP96U+BNeBIkpiApEfs+JLY9ZrS3zlIlpQ1GOpuSQX37tJMglZcrE9OQ
oGBFQ+iQNUiT1kmTJwkedgeR8McFifZH1EKnCchdBLBrcuHsuc8o7iiwMzECzilr
K+mSgyZ+tj0PMfNZevHxx2qwRlb1McE8O4FmogPVl9Fg+38+o2YdeFjGThpdKzCd
zdffRkqY8PhsRKuIbSH9cfP5IP9UPq5V1H9LOsfogDN6jjMYDoH1yHMcqgbHtzCg
c6GkOR0YHkhEsBCVUFYuhWohl1ijvgxehS5pUCkXOxAJwszVb+XoAxTNQI61WKDs
wIJgXnQmyaVAYzd2fi6POAVWJkKGzfztSu3mNGsfvW37Z9I/4GipfSZW0jEOmjR1
V4BT1tPtqvSEPdhWDGetvh8qSwi/Yy4iUEWr0BXF0YanyydOP7lACOfXkJUMx4Fm
X7dPdyT9a4A0oWaMTqFtrQtoeAtNtLned7FqftNjlI/I2NyhbhbexMB/6wzIvUGt
B+Wwa18duvAJU/UBNl5sE8iHcVipImH/J+Br8X9HNI2UaU2IDrWpzY6qr7sked/I
tcen8DHIro4XtKjU1Ax7jOJBl9hLcshE3YpL71qjAsjMlV0JjgeAe9A+8Wvy2k8t
gLcTWXm5/pSM4OiD1BuUAqlb8hbIhvko3OaiKPNCcT9KfSkZIvK3AkkKQyQa/W9z
XFlI2EQZZMNB5bABcks3A5XGpNtC2nvWsmUS/qPw59Sg90tJgVzqD/lUZvk4cX+C
CyU+YMKk6iGqpZfxdEoBs/cyBQgA3K01ICkyl4N0IwWGqJ6bKXVeXkknUQj6uVpr
hHNmGwUhmENhFzlRBM78mqX9MbIozjx7RebrU6sWOaFCfPGR5PvUVYcG2tv5wE92
Gs/Yu9Zxq6Lyq5iMQNl24jKJVRZdBf43lM6QioChnLQbg/oxroRGrqJWq9lr/hfP
eY9lsRxRWsCdC5NLH6jc76fAUT7Naj11jYZFEww15auDMAA6G5VwbNM5vnah9AIO
Pdis41qFDmJjN8+B5hD76UcLYvR8J4YiBdTcJZcwEmbblPEb5PsaRY509FueuYmN
QBQWDpV19zf9UHfda/szChGqmV/VKCBehnwildxaowHMtJjKp0b1GJsijF14C+QM
s5UiCDzl1Ku/8wTaLZlHmN/dX9AyzZ7UIRK4noRMi4KWNToZg3ufszTK7tC9aD9U
Q8iIlWFifEwY2xd5nh4oXY19wdHhcPybB6bOjWxC3FOaFaO4J80P8vKorPEdX7l0
778FrrpU6w1pExlhrzaQvyW/cHw3f7AjcFLjBi/SfeOSOSf4DFWQZJv74Qmur1Ns
kVtl5swELdwjNYoJ21pfVH6Ga+HVxiuIMLLXjv3quzgBxhuz8MArfr6SB8DtUto5
hRydJ8QDPH3RyjJc9FDB/3Wkqz6SLdKdrERRevIzae4MKiQYmMil3XIdws2ureRS
wFxfB7Akr4OFJKtPsgulHnk5cPolfQPl+IBWpnjNQqwoQzsg1FaAUOkztogVaLGj
yTi7C5V87WND4IMJyb9FNdL/HJSKKqGXcAfA/F+BZQFuuvRxZBhM1ky/ywlg/3h+
ex02LKQATlL2SAQ4i6hIPo34IykiOCfGDSXCj4M3Qdo5DOn79Ca7ejazAZE1dXSG
qftr9UywardBihx4Qw2g0TOEymTOvE8/S7ElqAJkPXAY45Z13jMMCNRU3hDyMw50
06MPNWJ4f0y64fshs1/VPStJg7M4PZefpCdkLDTVL1xxEYtjfaaWZCVxJASe4+fW
7Kj80GcK+CxHqhW+y1tWwGw/pudTO0d+DRpujM6enlG8m/gRnSY26UCMep3mFA39
prXiKBESZrddCyZnFxyiW1z8l2wsa+PEwOjv3oXLZR4KiH6sCjzsTOLIagOKamOd
6pNPjJlKy20SQl/gda7tuDp+JIXnWJKaSKwFGsxOGTPyif0D3v9YHujw7xliCY+5
uSWRHXdQ/sEaMOgH3CGuR7HylA7uD919s17uxSDqOHfp4AsNwQHHOOU8uGmgvs1G
7VlI+rK/wObDgmzmwVI1apD8Bcmx6KchiMwN/Kwkdcao+Nk1iWuy7qGPSArd8xOZ
NAZcXgXF+ApchhHkLrBX75Ubv083+lg4b7ulmM/Fqb5CxnHg9VxkVN61aIzhDIoE
mx0Q/j9hKncb4CGYMjxb4j3mkEwPJ7VGtelNuPiIYxyKtJlyWJQWB9V9TY+zAZmP
HFDQdlC1ieg/X+pGGxlhdjhh424i8MFkIhwYVMemta8Mq1vEd0EDyHfwfCOZGu7C
x1pPNaXVTG4+L6D/s6Hyn5tGs9Zn/2xiaQwuQLZ/dCGe17NJrNFaYu4t1aOyIfgZ
NWcjfHu+kAkv2lW91Yr9T0RkdfKTFSnbxeF8m9auKWK5S4ie1Y3OXZWkaykcVsTs
R1BwgWjXhmkjx9UeH/+LpW/Y3Z/dYGNc+F+uB07n0H8tpUaGaaYhGuzcYw6YxLsx
7eE7RexoqeJED1PPV7PZFRawQQ3shJ2XMd4EhcH4PJiFDKg9zaMyyrEA4I38+uPY
wV4Fz3XgAvjud5zwY4swKm0y+pDR3VbYZm4WsKRr0X/SKkFMKe+zKHZDGDDGhFaw
keTbjtNqUK8/pTMtTCKSNalgyfLOgywy5EVIqIGJeYtioODcoEzbVRxAUwqtNWev
pkjjvAcFTHxWsYiLK8M0IJgE9qS8wsBiLDDCBy8VVm2DrMhA3iK6Th5LY4/xl7tq
jZl6p7tWMRvPu+NOOoc2S8vNvKN4kOhZd/VjLuANAhAlBl7q4Dahap/li9s2KuxN
+Sld6EJ4Fw6BUUyUwCjqp/9uN6Web8uYwCByoSeS0CL63ey0MUAtU16narNDl+RB
NcC+THeTG9EEAal5xCD7o2I2kIiDVjo68l9gfIhwbyxsSdlsH7Jxl6pxrcT88dOG
YncEnlGF2bnRDhE+fLjr7ZgJCJz+Qri0sAmYz9NYrK+oY+eVGnl31OaqvBli4cZH
AeorqixDmWYPrbODssJg9yoOQESdtFYdbzMPxL8FMsY/JyPkGGJLFhnpVAi5UD+o
8fi1K2dZNG1ewE2AAGsdfXzGPuZwYXG3ooLJENOBsbaWRFdo0b8K62GS5oV0muF0
HkUgPT9Ak2hc9WURDl/oJXX8UrkgrOleillou6EBEocntk5L+FRFxWIcZ/q7wt0W
pBNQFHWL3z363R0z0YpMAYHDS4Wl9wtor6KyZdhg64JhTVMUlMg4SfW/mLg9UfEE
t9h+4m3u9+NcIdG4nUpjSvXjUPmhGUq+x9PRaAeHJuwLQUZLhIXaTR8GnTRMM+tD
2TLIjTcz10usJMdV2hGdyowwWWLLbpbXyJUwsIESTxXi6Ypxi9oIzz9tLPvovzKn
R8OcdRc2hJWvNwXFKsQSKxnmLSM0W7YK3cQuWVjgOl1xgm67b5+gcvVZj4PORSlP
H7uXD685BGMpk05fNNbD6AdPPkJAru7rD5c5fLz8G5gn/HZoyIKZdqe6YvD+hOH4
YCym6NUULA104FJgJogdWK+vuf3xjPgunYv3yJfkIRctQR7ATxJfjUudo9varGX5
k1cfaIZVahRY6MFBiPupD6b2WVL+XiuF+jUla1cRkkTf27mftdEOKKLwt4B7uOSf
a3e4EKJo3MMeXSg0obE7ZbXl2IbbghlMEHfZn2v/OqjD7pP/r7Zj7sXck/D3DYxU
Va2dHDngU+1/vKHnfxcbbvCtPDxw7b/2fDx+44hpIC7i/OfbaqVFN3PK4PkaCx9y
ggbQJ2a02Z7zmN1REdrS3Yt1cwYRsCu4dTK5kOD8wQCcou5+uOMm0Gol9NTrK2j7
TYsqMOuXHaJW5+LW/dGdmP/nd0HLX1I4vPE2jcpod+eVCvI32J87b7591GkI9k5V
KYMvSwKhYb0+GerFO9lHvYhoEUKW3W2uoS2iV0NHRcx6eWDlyCF8pV6HY0U2vU1E
SHAg5wQJBdFTmsPVHSy0LVlRhjtNI+TTHpuNZGcgt80mT3nih2wIhrdKWUKKECCp
Eo1rgDId1K70sUOTLQZp17gBhyYXBnoCVmdCFofUP9DIkLc5Maf/pEOPkZpVw1lv
G1ewANaHyYl+NNXKEsk30y4/k24rY9PduNTxQZIzA9unFSuYp9+TAEAOhXmYCGBR
IN5Qhr2QD/JqPoYQdXihWsNiH07WdE8kc7s47m1kZ12oAsAlY2Bq/3QDJcIIF1Q3
H2nUK8ZIjxy9ukJ6MoiJT4q4JOvCASOXRxKG8xb/nKkn0BPybal5SYxwUj9PtrPu
KsqRrvXYS8BgW9OWsfKMh0O3wrKwUFIPJUIieMEbSJjq0H81wv31DSK/aG4rv1kw
YvEBbGKo9niF9qsfMpZziPPO0hxTD8//4UVFcsCoH1sfnp63olH72PhwUgte5eXl
A0ZsJTgPA0oC+xBusPnceXkbJvd91+HkneogW+gQN5FK7S5qP/6tT2lIkzea2FpL
feaqxvmUj6Hhf85P4mIVKWjt9uqC6PLfWx7zSzAy1xiotZ/FLFVAbkxpsYzM/62w
n76+Nq/xXiRsCGpK86fRs3CWX+6lEFEm1hikI9jT9Kiu8X+YLQDaDKkrZtmZI/71
XTkSj5PtyaYtjF5aM8f9q/qUFTfQRjquJWDuzHKIa1cazJ+/uPwVSVMbP3ZvOd/r
oVDVb7F2W9O9F3oaZjpr7McRUextij7VSEH9GdwLKqvAmQ+GzCIR7zCd0aAN680X
4ZHmfoTsnKRyf5Uddfi6lQU0TVg06LHneOm11CViJUX4WE2hl6T3KkxK9iH5rrRZ
EnrUF3j1lvFMs0lqYOFCbw2HOEjOptplOCZ7eqO7tRjpJ9pa742yV8yzO5mqbBte
uP/bv4NNiz7IeezkWTXy5PonyCP5TIgHkQ+LS7k7Ro0EtPrkq/QdSfFulKqUWEiY
1s4pCBMkkancIIxbzcLJtMxs08N+trywKKThKN3r78fqacUGUPiGxNzkP3e9Jyrp
o7KGsnTAozYAWOa3nGuyvbqcpT/ZNs3qQ3WaRFE92dxJiASvN/jpO3rXsde1rWUh
JJzSn75OT/HKXAqFmpS47py2FzgAW8vuQUWhBJyEVKIonLNIU5DqSYMWjjKwR2zr
DXhnyKtU1P7ScVX4dz8T+qaoIwDcXibPSw0/umVtqGhkFkpKeFNgkZ+RxX8jx8DL
QYsh1zXR15iuuMKaGNMS/JKl6TzgYguNk+zlnoYT/INPTU2GKk5OOnoSfg7qmQXr
6TBmsGfV5o41wEdUuJKN71wmpIRbI49srOHIoAM5o0azVlvLCoEauZE5IMWtiIaZ
Dnlc2O5UxqFi2hFktdqu4s/4AWyt4tiqMMAh32mVK+NMGERlCLN1J6NGpizxqSiG
Mpa+ekydlj8aoY8/JyNNc/faIPjFK5TjFIKlYa58yfWcswZeeWJNg5fdGHL2ybg4
2MwV/2yO2ngSFlpk+EWMWriCw+mducb1O/uTWPL846uJshUa9m2F8L+syTIDjc+C
RdyrC79I3KJgZIRzwFL5cWudqdTM8zZsZqZq21YOzuclgOFF5s4lPKMk73QdLtbd
1EW71LIUMdz09NVk9RvWU0uCjrE2f8V4ZFAWC3Z3reY/FsXPDqQDODJJeK6XKTKS
de4FIb70Mebf7XntkUfsrrWNEBAhWAJP8sZuiVPqc0NaBnnqJZ3OBFLlTi9mQQHi
Lq/Y3wy3ftXoiGCwYCWrUHwHCxNysbQ86tDcExDkVghXbtxO/JQMEqx3Wn50aW3+
HdeHQuBPEJQ6300EA7tcKPo8FQrEK+c4Pvr8JlBU4Jrx6kOhbFwsWHFo108tIyLn
ohqNpPjpUvxDoEUkcbMMVhVKr+J7QmCSl3mfNRq5RHf1dnKHcS/c8lJSMUVWC2n+
Rtw0KpoP+YCU8NoLilNtGGudZfGaSpaFmx8GJ5DfJ2wygJeO8YVPab93J96s0VCJ
/L6ZP7OVg2dxY7p0iumqr6KWduqda1aUtN3lPRWKN2CuJqq1B152Hahq2dHfYRKK
/WDY+tOpFzyZoBHe9TzplSazcfKHRCnuJ3V63XmKSASNpH8/C2kUtv3kHUZhcuGT
OZ79B8BAp38+p33g8lns8NgLpviMlhq94mnlgUzfOn97GnEgaZJvb8SGHqDsvosH
B61ko34IZfcH8196tihL0cYyCwTuExnnpzu/r4F9+5EZZy/kJcPCKZcIZ3NWUDSp
kkF8aOqEy08U9Md8mb0+GbuOn3DU6FmbSTNEp9ZrDTdgW8stDbIGaoyJKTlam8NM
d0pG+g+1nlXB7KzjSPMy3Er+WZZ4L0kdZDpMhLJJ9EXO/yLrUc+UI7NRQZq929TR
vypwcaXUJlhagMSsd8R8JxL7s7zCIgJ+F1POm/mw7d4DJgk2l6CDzrZnnuCdlnEd
dWXWgQKGp4qWYILNV0QkhlcNRIN1w46JRWsUiABqzg8JvRC43SB7uQY5x0RWmbmL
HKD/o4T50ccVbguntEcOGMXxRKKF56e+6KgwcowTjiy8v28VUEjHp9tF6iClescd
oE8YrwzVTkUqg3gmkMKbI9w71ONF8vfPhcELrgdHyCetzzCKjydyOSJNe8FcaWDx
aN0qdFTsHm8D0F0XtFmioF0MptqaxH2d/3/2Lr8yZiyVgnROkTdxRGDzdfMBaxX1
38YxpMMF8ZIA6b3jjMCtZHYeXC3sHycFbdVBzWZd4TzCe2n10VdosLp4zJK8lFik
3DUMSqIJNkF23EuQuHlYHdS44VqxGwn/7H1NqiGevfJEfIpyau1rSHsN72ee3Nre
GSnDPIpdNDcCz3wSKEYoj8tI2ZXUyTzwFv+loBQb6yHQNSvo24V9VJoi5IuMjN1N
Dl25w45TZjerv7YEvIxTqjT0QZMSD4RSeCuXyBIz/dedAxHcKrQPaR5U3xt3FLrI
wza/7CU9gEe4T9dWMbTxoTW7GQSJOvmMvtZBqC/i2GVGzmjfe8O3jPioDfHxWh0t
/ji2axhoSI/0Y7evyI5iDZSZGfu7UB8SQmdwC2gANw27YD7LkEFCjRh+BuDZ2FNy
zR44iThsK02XW3C4U67MHng4snVz/O822ojKktF3cHfJHrGl9ANPJW2V6D5ERShj
XhjS0hYalPGxkN3YFsIWuZsrZjsDO2DL1NOZmAkHkc4YCCSXFfN/LwpA8NX1ZIxQ
7M1A8l3LMJskVs0Gxjj7VpexInmwD+TTEPO9fIZQ9Uk/BYBjlkly9lZi2tiUSgde
b47ZPcgZNrO7q72zDkWNitHg/bXZPlvPu2hIrEA9fc482tw+7SC7F1fdRBJHKzwm
V2DO8KT8aARPcN1SDS8gQceupvW9TnJ+0p9Tp9bJZ89X/I6j/QSefG/jhqVYXwnI
UIjdnd2yf4K6Juw9tgwd4beQKUWJkukQGIiy7aiKuWZmY1KG3xyNbAQWitUun90a
2XdSRDqidAYgP+5yNYcDsM1Xh8HTpj5+PUyFdVL6FbvoJd3YZjAh0WVvWs3x41fx
IBZ0HWDX5/YPDDXost5rWgWTAk/mcW+x5hPH6tUnSu9K9QyJ/3Y5a76wwBEgvDnc
x/o5/gMPr25sZQAIFU0SR7o7rAGz7pbKztvDvoeV+w+wxtfv3rYQeI95ffPe0iTX
zDuLDLVljIa8ofTl5UzrkZpJsyzXiysL9xlHNHibFy+4Tf3/QOFZEr1k3tiWFy51
lnlkyHznc8AjQo29qTGj6MshyL/dE2YJ8JpYjWSBiCRr0IXGaRzJ/w5EtdmEqfOc
RJH0LsXsSMpbrp4w9jZ8moXe1zXDXv815an1mlJLYtnTDgKcWV8En5WeMHXzwPC0
6mQFw7aAJ0cl0kNKw/Q/ih6TbT3JmX3Qgg39Pu8kKqFMATYcNANyfci0kRPt1BSh
HlwczUUAK9TpYaGVZBiVL2N1xAHb08wbudcywcepJZPf2LZTZ/FWzWTasYo23ZMr
bX9Q5m2Hx3Yyt/AkmcD2FsnhvIk60cFf1Yozno5oC7FIrK7fvxMwZyYcLtFlbFmh
SccxQrMssMMq0DdH0622FTT7NrVv9EOJTn5x5mURIfcLGN/f6Df1N0ptdVjbOYCL
WtHNAnCOAm2pGOWhqZ/SEXxxGa/WbxZiSSvZnXxQgxpZjuMbc9N/fWfhfyJDATu7
rXePqQPlLp9oflzaeTevEobBHnrF4spyrRcDnz1ifiGcI2WNU63YMr+vYT43HFpv
/nUVB4QnUhFCwVNvDv72YurcMqV0UrfVrrldFM01gdV7CPQWbnplD79wt98f6c6r
/rPOYGlvumi3svTT2ZDl5bguRNmcEsBPj3yoJypo/DQ7yZqECJeUQwLdj/Mdl8EW
gIhQG8rurVxi3wBhi1UOlz409f8BnqJ940Q1seh7z2RK6ENXbDbWSo/ZBuNzyMys
jpAofx8ja5rs2kFwLKfC1WHkfalS0bCGQFgYDRBVhUrXYYPJ1gloqbPJ5AeS+fM/
KKRAHDQpXIgAlaLHi80bXFkTHz21mcomftP4KyTjIJLPUWULuYP852kAxgWBT2nr
SgJiAm1L5R4zr2vE8IBkdy3VCL0zzIuoXQhCJOhOh4lTy8sOMmbqx5gjxcz3auFo
gD3WNqL3XtDBFzWKvAxXj/ipvfGwa+X5TuuAMZMJy/MMH3U43yp95DsZzfo/LOLn
wxGn95BbiZY+U8gZdSkioL77abGYs6apMurjlwC1cAIbU/hOEjGGNxQixcAapCXm
WDKaguQJCHDJFK3YAXjZBHSkURkLlkwrt+3fh/f7BHM8zjap2BIUXqa7mw1sC5Bx
78bdyJIH6uLv9t3AFg5H8B45HmDGelEDhKsxzetcaJJHJo3UzT8uTxvrI4kyhrS8
EkCUILdHU2jSvYqyfPdlcJk5iovlqi2W1c3arsKTXtsm3n6XfGqezCCrAqTgA8ku
97vngUM/99X64D9diRLMwcU+907fZ/VcD4vYCfA/RXh6qqzUXhf/dl+uc0mBCICS
9r6VBrgUghr1ILmwW91Gt0IvPswi7kwYxJiHIOHXmS6qz2JAV6y+SJryeitw1JOq
bJvczDePL0w22MgjGMLnJxa9dLcU4uPfsQKL0JGWl7e6E4gpgMOiO+q9WB5Mx435
hpf41BAk97fb+/tN6LOQNWMmC7Gob4MvVNZYs1sPlpgW/8cFC4s/v0oaIOrK6Vm4
tdXUEtG/AVVM7/PdvCPFQoRqOiHYeyhWlnINfeIVDY1QHrz8I60c7wkm7bQqfh/z
CRP44US9nndRwYp49Sssb6KY0cxOt1WnLNPMlnkFjwRcuWhx38yHWT6GO5feskuh
ZqpgxHp/ngdbiJ4n7vlF460rQwiLpzPG4CuGC9Xcj/kZK+JgyTE+vS23ZOZyDQvO
8ohk/obuFgDfkCO6tNPbEmRhfQq7wVpzpFvsbm+8i104D19XT3/4ymLkZs3JiiG3
6DEpW5+isryhYbF0r1al/7wuULbCLx4+eFMxkRSfEZTyFAU0qYykS0MyDm4+i/M8
BMUjs+p+xdS18qxw2Lw/YdNsEXdLt2KYTHUZMEClMU72Zk+fFHqkoxLIrSAfWKJ2
6qIMNE0tu0sfmnOg0rolXaE5Y6DAP/bl7klxA52YevJx1bSKdjmJK+rZHo9zC9C1
MG/ljwF1VfKyaM6uiQB7UnEIp+H9YOh4Nyq+7FUxt8mN5Limpmq5sR8zO8keJDhf
xoBVbH75so/OuzATQWli3v8AXnGhtN19ZcAKunsRYBjl6guzYeQEjnUYtdtCyhRZ
f3tzHJ4Cc/lQNNhbhLX1C118BVpmzsdNE3j684TUOcLsRPdhNj/ld90xHphrDJ/C
75QEg+hw/Y3CCiQGni3VNJzsJQ6+MhtpO78FezoWULeQUOi8oRiIX4w6/2ABsNt7
76VCHkXlNdCWyfSsa2OPSzt5X87atNxFqqDEOiesuheRgOxVvgpduYNlJEzaWIWi
TssGrOk21aVd+B+ddgewTPqzVsPQ8ZKrFX8Qf51n+APxOy7s37/2snmWIpgIejok
MVd830ApbRAk1QGaK9Ydak11PI5S6h9Bjm/uf+gx5Uir4afRyqlFQBvJiuFVvfZ6
9y2Phsi2AD8zqZzRQcvOb6Kw5JCNHhWqM95kViqlpLAxT8L7zMVYmmV9VU6R8OFZ
olY1BDFRRJP4rhV23N8vTKknN2Ibd/bPr2U4jTlt4UZbeiE7QB4T0yb1jjozBdwL
gS89ESG60Nr1Yk7Pv81VHh7DFZ3GaPVP84yirsqBVtpOVrqt5QO6AZ6EE5jsU2nk
w9j/Pnc0p3YnAEdnJF76iCn61+MvtvnCHJRls5alqpUXaPN6A8j4OHwrza7WHhb7
uWNDgVEusopbgz4ZcOqBWQTrMKJ8PddSoXqUVlxkFsOadjm8HuQrQTpdfwlFesLV
tSGM/tSkKi17QwG1JYM2+UA/Hs/+9JQqpsskMyobIkDeBdAod3dePd3yIfm3Zxzf
SjTD4V5wm/My3bteZAnpezO1DXYm9uQxh+HicXAdKdjBjIY7FvyixKnaJA+NPudZ
cntbkxC/2UGG3UtOVskcLUBE+qhgKtu15bYxpPgdb+pFVNDMjphN2lnGFjgPilkH
Fo6r/5qZEBAF0sr/i3q00bX7+JbnRYAhksmREWeTHuXg18DITy86Zd4S/bXQtCW1
KXC9QO/T5ysX0Fj7SdSfz6f/8xyYTYRdzaBekVbZlKcJ7gUtuE0Y8zFXiuOkRqql
U7D3n5Ae3wYDTjbccX2/3jUhFBb232EqFmW+932cAalzr0mJIirzNUygsJFwMwt4
jzHc6gW3xeBEKSM1d13OHJvdMHw78hd0SWFh7X6xII3lqAGIMQC9L4d93qSPxiSu
E4SRTNQhqX/MMdEEjegWD8+8KQ8neIald3t4D4GdlTw2bmWRhfQJ/QaeZVkQZis2
x4Eyk2zrrjDCJGAblEglN5ZRX660dgzQe8MA3zb78YaL0mYqU5TcB47OdbJ0VnAB
ILKGfRAS69oF7SnyPmOx4QOGBJZOCu4mUi29kg9pk6UFRMcxE+SDcnD05d/WWzW6
qfFeb7PIEiiNPE/kRqTE5swPm3FvjQ4ACiAU6/nPvGebZOtq1eqTX84ae6kdrKty
pfDWRjOmKJu1YKU7R0V9LW39FmC5yxbH5ACuKYavi1LgMLo0bc50usCtbox0TktI
KIgCojnfJsMFXeLuJ4RHStq6bG/yc4tz4lS1m8NcPiUhVdQVg6Z8KGt5fiZoVhEN
A7PW7wa+qLFojx7Bo3XSftnNj1fv5/JoDKU07NUDcKN+h4RnUtCI8BXXJ4PwevbA
BrNM+QzNyozvAQH0ChM3FHmZp5kOjjufHzkGWHcuaw4gGKjTeV0FzvQsFRDSiQVZ
sABfBzUdCVXWhb8p0XCheQNXdzP5HdcUHh2QnpQEggbmbvYQv6QpjxEL1UTYsoD7
JoFT8W/OSL1wLL7ovz3T/RdHv/f0LbtWB/IgChrarzQ5ozNIq41BpLDkniYZOrtG
s4AmQzgG1z5d+svMwA5cptJm8OMiVOxCTxB+zv41EeHqoXZBs1f7L3SRjo35I3mz
tOOVad2QFTLon8SGpr5z90tTshKkoKdVm0oUb3p/AjrL5WvdHrKGnNTHZdzvPJJ7
G9sMsnETdHTNvR1MIjdXuq8KpZagIfF5YrhqVFSZ9xeGU1TpAz9zZ07/L+tVo0Mk
SC7bg4lDvsgSMVpdq9sIM/+jxVREFRJU7S4CP1WdBIwNg99vD3Pzw2MDvYCbmltn
SUn9TGv1ABSUkNSpRtwhV9YNDXkbAYy7gLeg38Hh1ZlJutWnbncoQbLNRP2JaybM
yZZZu0w8YkFc50My+Iz0R9QccemqdPN3Cbd7A4+2e0PTjJfRHUl1KgW6AkSd8o1F
2eFY9rFsgrWTkIXioneLyvJ6CbZ02Tn7eH7pikO8IDwez1vMW5ZxiEzm2OghITFd
9HFXDd3OXn5S/m7nUcE7xz4/Xqu9Ch9zelAwYpWQgD7BobQJqGo53+/H8dnEOLZK
jEMDAzKSkBBWsJo3XEqU+PKfmm4mI/JTJyjHjtZllbUoCMH53P+NRhM9oTiPouzr
N+AOAzvLiowhousKSWKAIMN0PvIJsyt+Ec4IJIqlE2wvvFRwkaZSgoMj4Hjozjx6
9s67LKs1uHH4Q1jSW1o8WueGaaw+T2JtfVi+bZx4cEyX+rFIUoHJcxKNBllyhEe5
e7YbyO4AoLpv3pekcz2yoZ2gMnLHTEM0WSa2ld5bYhX1t2uNRV4Y+HBLVRSy5JNO
4SX/FwLhnsfXXmoNCNHEhQSCZxbVGu6rwnZoeDus5aNybYmTxGv8uQohewZWK2uv
ECCfHQw1ClZCDxzks4xmCOy/FF7nigCk9xuyMRHoa85lY3RtI4Ib8OPiNRu27vET
HYZvQQ8WYVVjU6VToVlHBB3FBgsvnZnlZYbhCEkAxmiDMg0Xxo7DL077wPN+nvog
EEr64wvPlpLrueiF4XHjNfc0xysMd+9+m/zdl9814hh5Lot4bJrBJ+7+L0vT1Lmr
CMEdzhUA1B/kRi4CC76YGjWpxMq/35YisGLu3oui00Ii/n9aLnnMD+a3Xkl3syDB
qlsnoLk90uYolL/bIKOdxzK4Bz2NffmxpGkfyKHghg0Lvl53r9Nck5oqeE8Vxq0q
4jbZkQEBG3RztydNIs6EYR4qErMRJyEHTk0nbteZ/uNYLsTEnosNmqQ5G+F1LUUR
42odEWsAbZMYk0LRZ7EhbKnKUfuNfC5sC3ffExI3LSyXKGgqj2wDOi+QsVHHmC+d
funnkfTTfx4OAcsMUeoP54abfD7S5cnDH9is6QNeqsMBNtpCSmDJUcoqek8H5hdz
u+RXT0CjAq/zGuuhfPiu6E+8Pp1W7roHpF7VqpYe9LLZxflnq0eNWrPzfV8s+r9/
FV5R32AlO6nrxKmkE0UvnjNNibA5w3BHWC7hLW41LF4VzM6ryCKzTfhZbR3onF+w
9jTxyBQK7YxzsOdGOsCPd8LjZvSzvW57WLWpwHoyJi2CdR1qvb/J5M9y0aVOMOzx
/iQT2j3lLpJB4Y/z9jSCe+0jai2785l3e+U57lGDar29QeZrLcSp0mCdiRn4UhuH
CfxhUnIdrq4D+g8xLLoNOMdzpIcR4zW3zSzNmCyfRZV7XlJew/ZKTSSgtASnWCCo
kClLwN11axkh52a6neUuq7EHkFYjyDbb1cFYtyJ+IrORSnC2bx09IQ3vZY7upIbl
Wjr+eocQfoQRvPJIOv5IGwOX/nyD4HyqsBLWO3MC6Ffp20j1buCAyva6h/Mdgoqo
dWA2XSGM1D0Yf4+qxFiJu3q5AYQO6p8/nG749Q5+9KOZkbAxBkjHhDSQ1Hfkx98E
raWwAydf+Zolxg8eAUsYCbOkN7QHdramcko4TzauSKu1/+IgUjmaKl91aB8cJuzK
euXRavwuBPOwDl7ijxCSpTjhbYEkNgMoUG1x/lO21TTINCywL5ZR6OpEAiPBfNLY
rJUGGzf8FiAMllcyXpCatl0B+cWwwTgix9VNBl2cQ7f0Frwqnyl8F+tSU0Dee+WZ
F8uz/4CWpbaIuRasBXQkVRHhqOGVJ7wROiVwavBdrr21Dsr4UemdyQneURY7HEXv
nvi9YlX1brGqGKx9jqFAzeSNQBgBktMhIjlfsKuyTMPbhLDjNkPcmpR4TJYRqYj6
EzaJN1R9u7VAL0w0CEAzb6wNPrn75SO8cKRjWCtDAxT6iePpkMt9LbxbaXUWEwC1
RbT3zhwG4O0zzd/lTRp2ITOWIBp9vkOh/+qHVwcflmYbAh+0D1Pwyoqu+GKXMy3v
kcuwj8yCLikzNySnAF32FhXBTkGX1plb+Axj74MHtjXU6p3PGR1K5xNcvCNmGl3E
gtaBxdLUYwaTIl1+SHs+Sd/08UVXRGlvIuvv0lrDzAypKr/Ho7gIG6QuNAd5S2xf
9bYzp75OpuN/x/rxnvVqrBn0AusEyr0pPUIjvouWDmwSvgMjz53i+SEMT2+W8gH5
ry1s7KqRaBdRk/Mvekd2LGyWoiv7F8KVcXcO1KDUsTpPyupP6f7cbMEuXaqvG9EF
HdMMGpLcIBs1uaWPkgQuzSnzfnf8NDZSp0P03CCP8inCtyHeDVPn0bSRzGYUORJ7
SdxI4EvJA2cE7y2cK9MDw/YpRGrIv2xTl0Iftfk8Mx7GOOMqtakoHuG9BDDXy6kz
/zPh7ltv9LT2tpDNXZU/ZX7woPewtW/Fmt0ubn1Th2bCiSnDocyAdP16GKztV6D7
prNAz7HClT6zvssa8O1/fw3QLLrkT7GCP73Bje/MTRrYDT10UmhtE80u7GUkqFoy
zMve+xtVSRVl34oEJ18DOpt/7/FaQdKJoH2FBZQMXgVExNqS4viLOoGYq7f347kC
I9qIFD6myzlWldXF311clZkgEb4gBWCPj5hXtEC1/9j1o7FPGl/SaheQZCi3A4BC
40GmyE0jUn5/KG8NBJ4k/yUH9WKOORFDNa7dO8y2jEqeLS4RyaEi2aXwPPbWq+fu
FyAkRV947xQwdBTxt6svPFQQYjavhs9Pcu2lZponE/NY9ouwxywB8/awjJaI7EtA
uqrEKJifPj5+bs6W0RqCIrxBP6nyy+AoWN8nl3LzjGOHM1f8luJRBMn/lVLocX4U
MTXd0r0nVXeV7cFW0e2X+CBsbPhvwYJQNd6aUZGV/gXAdc4GelYVBOvAjI/ufjQJ
NOTySXygA+J0EGSWFN1Mcamxt4cSEY1nxW7u7AENSi4EdW50Tmt3VEmbB/EZSSXq
i0FS7eXAcTAaCuDIMStowzTtv7o9o79fLuqT6ugWmFmiVL8zJ3hJ67RLWqykzSh0
sZxZWVWkBTYm1V/Gdd43kxUOOW657+m9JHWycVTN+d5jGgaCQ1DAhNUNBIpsxKKy
B+BBtrHzJDFx9CtAGcGC5vqCgImuaPCeLN4og3dPMVxWFOQCNbPUTYhAYd3dx6aW
q4/PUjJxs59bgJCCVxUZ4qyTYxEN5yu6c2YMxw1VkvzzWMivReMD+BKM7OOcbxTH
pnNWo1ydC8JHWn77GFa7d+2EmspcDXTJr7GxPT/faQxrXqpo/mD0nPA8TAxx0i35
ZdBhbUfzMSVMgHoQDCXPAZtYVFlLCJPQzQA3DaiPwY2otSepGnH0nuKxOFh12mie
wcqRc186VigErFVYrWOEZcFbSfZr3Xk1SNf1V9Yvo8VwqBmOIj8JP4gOepu0NWCC
4bjZXSX52qcw8+q2McRLiwlfub9YZ9JhUKs8x9WTIP0mQafiJgEhnnaTlMQLsdik
XtZ9AOwncjl5SDn68AxqdWXgP30hcmuw+p6lOynfWIbz2c/P3hS0PgVw26Ojln8E
EVFXURl50JDuhLnlrPquVdYk9hEswhCvQ6VJD3Xpx7RdfVeZHIbN60lW0HLyg6dr
rupQKZim6EnA1IkzQVVz+Ejb95sX6TIZZfNz+dEeDF9Yb/hvxNEs88+B3Wx3IGBp
V68MmMBgO7/fFOE7di8EIQj78DV64gCBnd2wncV+4I697BShLdAz7uxVYiyf/nJu
EekEoAKT4kbh0Ld+DXDodi9pIp7zgv8+sbdglYdxa4E0TKgPhLeQkI2AXD7PEgGU
AgYozM9XzYpcqDThsGbdIU8dr71TcjnTvifpgpRRAUUGxoxSR4pshH2afDq1mflq
Rzh0WGygRmAxaRlf+lZ8+NoPSf2YsKMfY1K/F9xkrTATuolxQHWfY08H4JQu7XaP
XJ7ClHbIoP+ia9T/3lhug5fXPHhUZI/2xvGEQaGMcGWIvG1NCkSuF+iC13Mp1r/J
NV5p6idRKhxwUAWwXS6GIwUKToT2ehdtMIowO4bFIY/dEnBtZsZo9le2BGeZlCD5
6B+e9t65VUhqc1hs/bOmEtzCSrnj3WjpbYVYBMTReBWp1/F6iy2JkPi0U03hkVF1
PbmBba/IwSwtkvFX6WuFOtkI9LGKvNjpMjrgwjClKBzauP/zlMD31f2qWjxsgTf0
QKsSlpnD0ZkpN0SoWID92928YrzfvpOM6Fvr/e61Z7P0uCBvwFk5TmKd94cvYMx6
Ker58cnVLfe/bzG0MJuOBP8uXFFR4CdLsQv5D86ASsnrA3yPTkTNKJhvVx2VAX/0
5KWH6IRQ+OY+45/aO/iVXs2Ys9ExWRz+y9VGvPcEsuhoDOkm0581k99vOji0iQ0t
8CL1SLCIhv+r8Aa4nb5nDLGgOn9t4yxJvizFi2fZndl8eg75MBJUV2Vdx76H1gOK
yDsWO6gg/WlOdwpqmCzCPv5yVbx9I7SCQhwRS6Wfkxd+5b/3PdP2q9+wba1MYJr8
2Vo/R1HF3hR+Is8KHfP9M0i6iFSNauzD16YaQQhUcO2oFL/3pwECiRj6xXwSq4/s
6jRQexaR+kfjsmny1C/Idgj83kYaccKw4bRypA7vJU39kxSHqb7elYnraNxlFeam
LOCwSVJwf8yBYOTC/ijHDFwt1n9Nz319fGLBWWj9IqDzBJ9cNsQ3NlZX//ZOd0V9
gfeZ/S5wAGLjGluXXPhe3XfSdvfYmXMofrltksdb2AU4J8UV91Z7IHy79H9gs/fX
K40ottymwYSadmM/Sx5wcEwB4R9wF2ETgwyJb6xfgnVl4iahRFWvNoB5DC4nHPte
PEXPfDeH2yOmoySjLcipG5nHbVBGWtYWsBPzFIuIQZp5kMIDmtwpeKsqc749W/Mr
0tNYYwhEzowShKYIVBLwqkXobMcjxHuPkx23eRqX+xfO7tBID0P/so3IF0TXyWTB
uo2w2GeiR2NeCfeYfjAy5jiJNktH9v/o5f8pgr6YaapeCGlZnRElQY5Ffqr4sgeS
S9GF4oJ+cTCh+VjkR+g2ZFbVzmpntXaD2dHk6yBFLQb78aR2iw4oVi+n3qB1ru2j
4nsx1k9bsz3G55jHl7YnZ/RhSScZw6A9IuWcZv2bSPbHOxwrBdQUTcB+G1pfnDoc
v9bU12sAhoexBgXpO4IED+MACehHAsjnxtAWsqWSBv3VBRzRd1cLN5bxGJcI+nA6
Wt5u/3BSNNfWswrbdQQf93xCETTb5FgJX/cpixvYV7Z4CTvdUFT3T2+25+2nTMe9
17A/3wkeTLMe+EUa0nS2s0HzqXucFnJdbuueR/E3qSIIp6TWpZ+t4NKgYr19jfzw
JUs478A7bdDCyaGu8JFfocoSffgFpiL0DgJ1Jh0B3Z1MwaI/sHYjm87YfCLbWY/R
3au+X8Yx9EM+vM9q84+oFKnw/wBCBjwmWT4eSPSsDAlCKTi1st+gZK8TrBGVLZyC
dQ+zQD8cRJUZyff7VZ6EVlwWj6guBNsgd0BtEjd+eWWLJplZKVDblMJvAbkG8Ct1
+LPCsk/f/0E5NBstrpOQg8NQLnBAMOWbYgOqu3UCP6YIIpFe2IrYROH67b7Y11FQ
HXJFDiSs9TBsJszV1jjBrNNLoK+ueRdXKHz8ASW41iPjBHMdqI00JigCPshyFrVU
+B3DAc7dWYFa9sbTBwowQU9CcNDK/9/GVUSo1HWdxPycai0ymvPLoV2lmqJBznuU
K0ABuy7jU7ifdCStFzyX3uMON2TJZpKejCO4FpfKNzkuM1BW0LruK9Tts7RI+GO2
VG9RCoBvr1yhDj+KpcRgfdkM4wo0faO3TLIfleDH9PUTBsalvT9q8hn/2k3y9doO
B8lkZ1O0ndMuW69ZmJ4QWuBOwQH24pONffNs7by4EKTJNPPAIfjTwmAYzwgi5DI3
Xe1ZmX4sa4lhkL3foGsinRCYvwb3aLDIGeajaG1E6jD0a9HLageboi2gfezyeQd1
K/K422wYeWouIad0YLWQYNC71YQ1ejHIHB2YyoFAKziGzalG5XOPcJjeta/NGSfa
XN+7lkbkIxBBYNPyAaqOtU8DguHCJPb/ZGSuhLwCNH8O7y8gbfiLUBvTLBLr6WIo
l44AUxOWb95vML8SXfR991imPBLRyDw7H8ktRkTefXJZeSacdPwTN6pIZZpF/p2x
NSYQS9rxkb2fVvC3lr5o45UK70jaetxsarpTeGmONOIssDYxLMOFArLHST+dDbX1
oS1PXNzOaH/KE2lfhcFMLkb8t7YSvsg5koUxS/8pIBojJipOcOLLLHCBgC9oHgy9
1S9cJENOBBwnfbh6PEMEjKu40rCFAgQ+YU53LuSs+MEyDdHo7yMxZfg87xSx7qhT
gNWD+MW2xwAMJTm9D6zBNNNQFJDsAXG+oOV1iBgWZ+LzUCP/EIMr660Yjsnbsm2j
pgfv7dhPrP918ab2MOCrIh4lt/R+sVOGkkl/42AHFMawf5ZO8DoHLGM+CsW5OteC
lrlxKnkX0tKzJengSrARc4lnBq3vHari4ks8b9q0P/pJqGl56yyfKK9lCgYYIVY6
IBVci8yfb8dgLp/rHSO6mphwBnazF0D4e+ELO6w4Fk2LsjUqWJbC7m1IzXQT6ndR
oL5ZZIx0mHSYsUjT2uvrNPTJUOfbhwV96kW4Z76wFlS/Rp+6N3U5WesJN642MD6V
uOUNCBuKygZ0055zsZdbY3P40o6UBNmP5P2hdUwehRjUebaTh9pEcsP2NxggS7XQ
Y9NpMa7vN64AUtYA4ur/FIn/Cki0ZGIkuH4UJj8bYFLSv+vJ8/wnRqdEwN8OzPf4
NGM0DydTAG1BBzVmLng4W3tVJ1aQ0SYSTyU9SGWOpav2kIWWxW+yEXF8yYtbKIkE
3JMzUALOdRRnLbEmy7fA+xAEZICWlH/nRCMk9NTU8IoGT+X/qM+/dw3DKKfUkb9h
xbj/EWyqjN+aLFuuzQU6BsGvGCbb9V71sJXj6ZGrWQ6SB8gYcDEzPh+tDcXR/S8Y
Msu0M6SDNpXEQge6SsYeISLMPmfbiGC6fYFStYNUNI5T9mSaxkTeOA1iRIXaVyAz
+PZDSHWUhwJdbULy3ND2y9FFJ1vCUlA+iM31YuPXS481uLFrtcKZtY5pMbR27GsF
j+H31FLbkZDep+vEogrmYtxdNfA8hL+ZRUW4MbW4RK0h9RS0PzTbq1CzwBjqHGgI
qDBvf0suaUFTJp4UNqxa9lq60SmBIYE8Hpj5Zlgs5Rbglh6v6dnIt0mMQ0tNd61a
b6xifFungTj3WLbM7zFQWQAZsBhCVH1ALyoK/Bq82h+gKhUigVGoQ9JJVl4awYww
10KvL+jk+cMaYAs+X8pfSqrZdPcouTZwoCBc0370BQXs2VPg8kJYSDlUSfkmzAgk
Y+q4BYym7J3N9kFY9LIhiaYL4tlhB8ozIfQR4uzhHAEXhOiiaMizkgxXcySCIr/1
OT3srz0feXhNDISf3GldpscqRW8AEeFiOGJOqKIpW0JODiHgPpToInsbzAvqn/Jt
6L9ee37q0s8tUoq05ETbaUR1hul6Sl7HLJYlddYaC8ncOF8Iecn8PwSMkyovTcy9
brLA6W7AuY1gLic/gzyL/OP2eiJSS1OZ7nF2QSPMyvJ079vy0MZnh/luzK7yDR3r
g19Fo1hW5Mw1XIPQwFbkIC9/O9bGqnHDq12aKys6Nt9k4fN5IO0ZvvGfKgkG1OVp
993eym9iTjtb6W6IJ3n9fgU8SJ9B3gInjYgB7HFjsUjxNuC4haYqeI+vsFywBRP4
r4wvffQ01sZtrI3Y9kqnfUvzAvmEX0iSQpMM1zA9CU8DQjP2hysLaHx6Of3xv3TQ
LUx7VjVXIApjOSJmcAVBTzYi18v8+mzE+vza3Wagv0/w4fy58S6hSfopLLySyoPs
B58EVwIDe0Gvd32mOu2n6D+/v7ZkEMNGhrvdY7pECMNOSxdYCaPyQrJXhW9ypXTh
6/TndWI0SQA1/1qVFJW8YwnfhSoNVFJrFAPsglh+7SlAq9hOgNQeTihVmaDqdw7q
/+ABrobMY46kZgf91u0L25gL6qxvc1i0il8O/UL3Q2asZoju2KmBUd50qHPqLwmh
lJNfSL6Hy50KDdcIok+ZGKVwXVjkyJpMBG9Y8fcvhu8eKHrH7Ik1UgtiUKq2EnuQ
TgWmBxp470WREpK+DeODvnjt9KrcdntQb8eEMVWtHE49zgYUzwlEPFPep9oDuK4o
uNS5+dtZvNEoIDps09IbWXzpd+7H7JPQwG4zHqZK6/uI/xALgJRFZhRdHigZ7ZW8
UObA+Vmtdx7kNH7NA2nF1B5BF2ccMOIvy9hlX5G8TeWk78ZSxqV71KIenyo8Xdm3
V6D3/tQYGuePz8CjlFjCIYf1+MhQ4VUtsxojGwKsj2nA7zpmEFA83zcyGAkkdbSB
ZhJQ+oY77Iy7s8LvQYO4tLdYPGNCkbOYC8WJWTmGwL1b3jnpKy3LKLYkkFNe7Pq+
TyjzWqrSNesZnmAvvUxoM0XzaME8PoDgT/Y+5/L5Eovk3Ej/5dBdTPvndmec0H39
dgb1zLadItlNxV0qlmQhP3y9iD4ETAoKrA22E0SxP9WroYLKn/9TIBlb/yrQeUE/
+AGUmeACh3/5oWmjRA9YO0bIpnq3rAhulyzUT8ZpITRzZQL/zFkFZEdq1VHy7kru
r3klwVaabHbTWWclEYwThSPJrehRPX1j5pV2Nc/RnxLeFUsjfYxzZymT6GWTe4Cw
9K7favawcRSOe7BMW22TnOnOfKTwA+o0COIN2JLxScbKUbxXieRNhA0b16MnStod
iZWyNEAO74/nLxESupDU5SzCDmc9qS1APJmh64I6LqD/qdTZy4ThqFPl+RhN2PfY
eROMnCldBouWo7y2qi62+U5jGkLoTi9vlLEBIx4JKw7Ps7gN9higVSpUGjzWaHyQ
9HeC4dq9cehCxfWrmpON1VQqhSPemGlu8vw8syk/frInfUI4QfrJ0vCM34wFhqhl
lT5QHc2jjFcSU5O4JpcUbUYFakiLeks/R90LheHCXXOxjJlKBuzZWqbCLXQHnUB9
6Yas48TOWCQW4K3w0ZfQ6pR+ko4jaWMESsDV3teyrlA8SP6B+7TRxEsrIvN7WIMv
wxmIkhht1W0G3/2EChd2DmcQ15T6gk8zwK/BIJ6kd1MMkd7rfQXxlyjmDwSz+x2S
2ACcEtLpKDqoY+NuFzhpZE+bLDRcRSJhIpmwNVRNsqxD1WY8dJmbt4rHS2kca5nA
Pg3JItqf7N1gV3/f/WYmT7tCqOr2bvhJvwOfUwcV9gLWpZt4sZmpXQFTMtGoC92l
dumLvnWtNq+ttJhgMrq7/ceI/e4x3XwRv4e0OGKEf+xHQQ6VtzACJOF2nrzxogOA
C0kdB3onT5GdArGGXLI7UYa3uICVQpIAh9XixRWoE2GPf9HKJWY8zvlySk/jxlXc
RunvIkiYh4yAg10MxCdnzQt+o8RI64bCa6+taFwcniT2jWb+jNjnn/vAUF9OH976
JK2fl3XcvE5GD4/jWtXslZES7ORIORr5Q2M2c5f+03QJaWAppZ6KkmmG8/IDcbPc
Foxad7UXM1X/UFaoRH+00RqVX+dvnvpfKhqbGBB7GqxW7IDDOdeZnqgAEyyfyXYo
t9ID4zo30k9CnTs8+Dz51ZwA5Y+t0lh1/JxEg3qmkbVciN0eOcBplVZZBx8A0lmK
vtrlUwEpRapYtfp+Gp+sDC94zsisYEAPqThCFUP49XYr1KKmAZgbYutK3NxNXfhb
OFi05FaZy552drRjNnDViSvb7oKbyamQu4TXtzmpFiOjBHhNw4KGw1xJYABucEWM
OSDFLIXdTSA4w1OUEMuh9J+q1UnLuQbOa6CLvqjr5qhdhFQ8nB651KnLuadOLi5X
HXv6J9qiT4oRzI6gCgM4sxaKktBZW+v3mjl+sYMOIzJsiuhXutOi9UXcvXnDwxmH
+knVdmezRVZJKT4oz+DsV0jbzP4TICimiWICjJFaVgedNa6m4loLxfma//OKoqS3
Yzq0nCB37+SLyMtsIxMDFUOCzVFWe1SNUaHEzppjGMir/O9+jjars0/+76wCBSGz
0PFHMzOZ+mff15pHOwAONIPepcDgb5itUFl6MS0UwKQ5O10ihIPDZD+JQGszlp2h
ndHjmSLlAA3H2ZZuzpWdzEAnXsnZ8+6hUg7ZPVkxSiRrwexxeaLiu/KY6JPTfFnS
swNcQK5LBjHgGNI/J0r3MiRjdvXeNxdMW1nNBFVGbxbF0N8PIhYmoyjD5auVnaU1
Or9auUG+5npMDnHRB5hZZDTVWeX+5X0v+7zD9ELPpID7lGPosUDR7zotslRPCeOi
WN7n19SC+zCTzDNOJRL0JQLMdnyFYmtQsiZYEjzLI6JafJd1k9rgidAOlHb7Mkc1
dcu3JcV31R++RZqgKxirupNbEEB0RU9c/o7SZNJbE2OktAHcqP//ZmVuy6sQZUhB
ghYM3hB44OoVd4V+uTpi3DWkDEwUIg5ExBZTN/qHIN23LOPcXhVpRyMxqB96cISX
eW1xvAhohJbbLvmyAt/7QpiYDM5WmswwUsusYWNOD7DaTvXoNL+EPCktst5/p8Dj
ur1ozDHqsYuHgql360ji2OnsuGY2TejDtI8Kt1ySMex5bvo6VBcIfJXm+g7gCnDA
6kw3S0Ebw7lp7O9noKdILPj2fMxHmarZyTD2V5CIpXyH+CF+wyhmx0ncQ/hSZfPg
IlHTV9hYJpHpHcNad2+1DT1sJALqdj9dEH3GCR3WsRZQ13KHPWADO3RHPgnzVyhY
de7RikGSX8ZGv1y7EVJ87xxfAvdKTPFNNLfswNuHQ2Edwc9bla+R7/nhgdMdg/8z
zkgCikIT1jBFoP1cU78WDIUfPdyVNF0IHcwYX+X8WvhCTAxfZ0ZN2+I0rPN6aZYC
CbUZln5HWVKVvsNanvEHogXQl7w7aJf9llIPivMhGITUFv0Zjvk+A4FidDiwTMON
rPTrZM6WaISdYD4v0N28PA6UtHM38xW0jSA+6yvOysKF+6Tglqqnbzui4ndgXEM8
GxqM3NBmDVJEitoMX/jRlBy98RH/xvSFos7pn8t8s9BY4xKOC5z3/28TRFZx6e9x
TTHGSFBEKVrr1Rv1s2a2IGwQRQ4yRzpwvDN+mWk8wRlYq5Ds7cPbGumX9pR2eyAA
SU0X+l3cuhpilUPWvz5m9RRSfYx514UEIq8Mb/FaTj6WU4gr4SOWE37WIZgz14MH
r3QH7yxcxBHrUW11iMVwaYxZus/xcWAPnEy7UsIzm4P6GDYWr9pLYg/1S7hw5y3v
jHqHxd3jNalOqcReX5d1PTyzdG5Y3PSLjO5LUy95qTUWl+tfwQ2wTZc2C5QHXi59
NQiF8mrs8DDIr5PvQeFmq43eYSqVeDQo+xRCtcCDMd5/0L0XA5oW6PCbg1SZYdYn
SvgHK+Ng/aXYrOVKxagjlaUxehVUwjLWgyZJuo0UWmVBPXCiI/0hprX6ejus61fK
AM1hiqyQU2IPL5hdUs1Y9jtQwEBHUtuXIOD1x1iCnhb4n829wPhg1+E22+kt7s1s
lsOjcNAKPAgl4p6ilSVMBgRDLDer6d/83jHBmr/7gNUuq+lQWSmTPkJsaoAeTI64
HhynTZTOS7DiVuUoixJrxmLrWHWYTXStSgKcSQcPlipG062pHANuUmz5taSBbojr
UyDhK0JgzBYVKKFXg5TudZLIh9uzKRLhnBIEjws5F8itYMPfrgYwvVaxwF/a5iDy
qltIwIuMwnaf5eBH8Ordu8UVqyx1b4aMDfLTXM7DtcFYlbGDExVsYIaGaacWMvI9
YVEqdHsTQxFz4Q7Vm+icLp91wDS5cn1GdL5MahshCkZGG96as/p+DfyYQ4VB7+HL
aRFpOLYD3EQ2tDox3U6nupwKsvV8U2+7Gw1Kuu712nR6utaLgeB7dCQm7xLC60SZ
m8p4qpVZCitFKqLh0zK6KupQS3MAQOOvrD8ydoUTfqsFP/yY47t26b6VEU2leT4T
V8OoJzyNwkuAixCZFdRZ2+BdhWM8YDQlkq8PNadRa+SMUZ0qxZkKqBbyCrTeANyO
btiPWc0q03oEz7HJd6S5VsWHZZB70QOkhSVtG2JHajs2eXDtc8zzMyNbR8WDWF2e
ImlM5FVp9ydt1R1TZ0Ozy/VBsMe4F800s0JOxbPPIi5uGNprQquuDgLzW7n68QgF
WdNgJpxZUxCcj7xylHGvxY2bzvDApyjHr+aJsSUNUdNyJtueNwf3lFUQZHwIU7de
hqmVBpvSzoFXQtXFTklsobxGo9nL6PqyWEixrkLvWumkTyHUe1pXy26/Hj+o97fW
J4wvu2QD6cgpe5xlNq54Z9yP4fcxfLItZSkj7Kl5jnS37hViqVctEshFigkhNdnq
SS4+HZYjVDzLGdiII22H+ATPdAEeG5p1CDT4S1kEWe0RoABmNtMvX/GcZ6BFKAkT
jkCiiKo2qa3uwNysKXeA41anJhI/gVeuh+2TVVWY3P//5r+1bVGyEowKt9M+QXcM
bsF5fgxfzIbcCiIwVgAJk3xbICEH+W4oHBsR99BGpqAk5M77uS5cLiCGEhytcaA4
qSXdBZF/bccEMvg65ahQoJnu8P6A0m2F2wrtoR1Haf+n/Z8jfmr1X9F/8rhytZLv
sVCUeo6Khd2xg6Xr5aVjp/Vt6OzFfajaLPpAZ1Aa5YKWsHHLKFJuwz8Ctmz2o8mU
C2IFit6kgKcxfz57O3ZgtHi7QmobS+JL7hSDfmmxocjp8NF7WCoOiSYiap36Cgag
85j2vQrfbaSpCrMtId7/WiYVEZnhBZrS4VqprSHVDgLOsIPlNjfu/aGqkaJVDZrH
3tFmUYmngKl8DdbEMxrseopZJdO/PonqJatgTWRKo82WPG5aRo4BQmU3DIEpbz9l
VcuHxJlWjd17Zc6VO0hsdNP6u4SzZX8IHQya3oduyJvr+XnXj9eryP7hc7rMEzOB
ylNjvVIMCbr5IW7OzWpii6Uyth+Mg9VgZKvavl/CXzzzMj9nq4RxUP58OVFfOgRm
fbOLP0Dz8tPI7t1gsNji9BM0e9Ha19Q4mXcrxWcYBTH1/1t6RQ3KgrF9GUty4MkD
+cMfhDmfN2HPkJCBQTEtAiB0hu+xn6EeD0Mo07dgRCvg3ZzHi7FDrlisFd2KkClo
nC8c3fnLXfAtlHLJyONy65KwxJ3C5uS7HTzROEkfASkxIU1JLe75TthUBTFKuwIZ
+jSI9crlvzoqKu+7jTSNqlBgTqCguzoH81KNpwC6J/f3ULao13fV16VbgaV2HGeD
v9vKYIzTTXfhiAwJe2EeEkH59sokAtWKQAxLjPhmkfDH3pJ9HhaZ1DVisY4C30Wp
p/R2RpPJyQJYhXYSq9MliRf8xwH/hNBcXElQe80/pq3hBybctf3i97G0W2oiZlBS
Z2bI8vkOz8DMmG8eMNqCeTy5YzmUTEBL1xD9HMX9DK9FJIw9HEgBfANp7Xp1KR/V
ifJVfqwfj7N5P2j9iuFTz0QpsTPI6lFsk6Y73EZ0vdY6nE0nay7/teLjjGyajO4a
ViO1p7rrTl9yUheIOGvaPtHVxrAc9V+BMF641YkpS79K1zwEvxB3bh1GuYAeEkJW
jfacE0+N1VXx0WB1PypeBazY8KcCEBCGFkf4l5u8nlM2wrLrCVNmkvJtRixEEWOz
RjQqLhMIh1Q1PP4bWADumQ3URWydrIut4j3NbtrWXXmRmSBJO+1XuLyYQ9sy/bmy
KPgz6+J/XMtV5l0h+ttgxWCFNwxOi/bW7Lp/Burlr3wH47bbSVapUPMeqSVn0KtK
gaiSuzCiJEtvV14cUcZd5UJDHG+S2HuMYayfUI4DluEUD/wKY3kbps4fqDx5p4qK
l6cKR2d6bfL+Zz2DMWH3rRKtQCh0TcsfasLxo234yWPQbxne+95drpEchL/XydvY
Rv5KeyRaTQM4fH6f4tzBRg6Hl3UMqLNwengusIJi+sciuFXk4OWFhYsvHfC7KaqX
ew+nWMy63FS2eEPEAU2ZEUg2+bhcxH40wOw2cTJxOQPsH15ECWNHbCtaXB2Z1/Nx
Aq1xSweWNy9ZPsPwqvKXyTORhnlsPK8hlCZh+y7KREWKEREFdJeX2ZJZLwNgYVrh
pTIPPTmwDIkV28wyWzwL400QgF0MQLu67HP1dni3vB2pE1SMkvO4YOIfhTp1Dygo
YJqp3CZc4fYtKEix6u3CfRwboytMYu515nkTxxRjg1h3sGm3zFtjcOTjhvhj/f23
fYVydipHyRq3QtiZ8VlvmJdTC4hy1t2Y1wPXDj6iKW4PpF1zWbXa7eNVXN/IHQt5
DJ7lL9ZAi654exB0ljarqOGOib/SPhNV8jsFOy2Ss9I87qO6pUe6ey4mcECZBcDf
ib+gaEm6aGrvh3nLa7mnVC0L3xYfpKTnc0825eC6XYRg4sqKhWQWPD6ZxPrWQUw4
WUIhlEl3laHyXmhWus9K3DIwl1aCu8W2xdn0D+tVlYqQonD3eZsjX48Gmfjb0iy5
EksZjU+W4k/r1dcqYqfhJjv7yodOFe10v6VKG4WRwpY4IJnijaSh8OYb2T4N1GUj
Aag1fprn4u4ttZPOPkloAEuwzvJ3V6TY7oTwG7Bfbt+aSxCUH5w+BvnYIlZ2DV6O
Gtn00Qu9RdkoGJGoU5/zJLQIODPpmmR3IksmiLLnj2s8SLl2ItylgEDYmZPZd7X5
cbVFfGt3kHSffRt4yaxeAtKIGubYYuv/lP+eWQa2xNY4rYGvZbgRzo5TW5aWISlJ
qK4P2cUrORuAqT6lNcSQc6/ZiiMD45uzPtkEM7cC2M8gmS63cpXN1TcuhkvLNj7y
BeEtn5kTMHOqPV8bVojGUtpE34UvHNnhhumk0Nj5MtOS6MYeooc9ffxNqb2v0nq/
006fur1wKfGMltYlBMbhHeply3ZakhRAUkoN99sf9XTYjmz64yLh3mXvyVz5IO01
ZD8HHlKjBRduyJMHXSg+BkIrHYAespLYkq11wyRKIaRdECdLhDgFXo++qlresyn2
zHgZz2zox6uAGiX+oimA9DnxM+koMQl9kHh0ED3oLidIi/ClQppGBrWkfhWFtZsw
Ja3W3yYGQE37M2oOyc/f0IQKnVWOrrNlTa0ypFFuOLL18crrXkSBRgtZlRS/oe5P
ixsKKatYZyGYiVwhSjfsxKVum2sAVDL1HrX7saMiOjQwTi38oAlW+BuLD8W94NRo
kQAihRGOmcC8H6d3di8zwK9E1R6Ed2PF3P9+1OewMza7P4syJxhv1yI2d6yyHAXl
X9qvgJ9/ftEzl/efT7rMmXh+sUpXuo3ZmcgR1S6gM/FO8OITxfk1BEthxPpuCE+7
Ehbi5GAuZsdxyhqLwKDiGbio10bQ4fSWYo53jRFf1qqnEWV8dce3+tfeowlv4Ubl
Pd4LXgmSUHjl8KjI5pT18vRlmnlt2tHYyFio8qTGfa6NFM01o9XOE/yq0W0aP3NL
wdV1cQ0pF7PmUacplG+HWysfsTccyb97C5AkF/Y498iVO9wp/aUBst0VH3nX+XZ+
pDoEzK6uWPx/1n5h3lcFwNqVy9/GY8duS2UDeQUxSxj/mYouUiapLgJcgZwxlzS/
VeDsi0zjwI8qtaKp5+RnBPQfIhtv7Sy0BgTzXt6cWgbHb2B6sNbtOBLUfI/6ntaG
PFG85JUw7sHCLSV4jdjhYcMiUj8dppUEBL4nHcRgcugx5otvkjmLQT3GUdrzY3MZ
qxRy0XJ7auxVcP3X8w6NQwWGOn2OZXwy9JkMiyyjjgi5E/j3lAidl3brH07iaHS/
U/ZeeOuOF2BhH+GkUVW0sAzhkXYmZszV6HIUU+iTWEqxVry1woq0ZERtem6om3Il
mH6LbpTLste6AbSJgomy1abbGzQnK01qMbLUHH0E36VLC50hyhTgy7tLTjrSFY5e
/7736pZUctanfAsMCGWCPMAzDhr3Sb75Roc6T30KwpYMceZHb3F5BWPCQg2v14mv
773R1AtFI9kISuMz82NnDiCmItGKjId5kL/c+5WgowiL7rmFv3hqsjUC+mGjUX4k
VWwD4bFOgKDkOkRCGDPyA+PBl5ug/6/a/ankd/4rKju59I+93PpXWSnw1vudI1es
v4hDfeUDkUPJAQAzeHYny6Vm7QoTXAGj2V4gWqHK/yOkFShZWAR69Wkxiihuy+1U
pxPoR9T5FnciEtPMYXmm/WjPDNGOulxaHFMGl4NgZqbSEuM8rBjitalirWNdB7N7
Y0RY3eSO2f6S4Qhh7CkmjV30i3O4bRruq4qAnwZ6rtI/oQuh+vp3BjJefjDit4aF
LOmHIN9SWhLRliDDUoD6db2HpRNasiZlCJaCLNAUvsOtafb8LktgxEPYmPi5rfc6
SEpTGgjnszkX1vogU8DzCJaQjXP3H/oIMz+ePqfiXhlfpUvH3eBYOY+ozDyyKk5z
ioyLzxngkuv2miTssNXvTLsxR0H7c/l3GQ60B3RLAV1DSCOKs9bH+WWRUBgHpI5G
2R8KD9LDymO3GwosuNg1pVKbUliJySF4t4mEcqROv7y+QXtsS7L+nqa7BkqjmFti
T2CQrQ280K33Y0Q3e3N9RTnrwfARbPzide9h4c8anHwe2/hwnXTBoNVdZmQLXP8x
AUvndmD6E/ltXC3KaXCsEvmpdwNxqW3Tohwb30z9ca12FCDG+o+w3/UjID4bOOY7
xf46fooSucbBaKI3qTdqwjzppp/IRiiRCJzybsERpZL7N5z6QJDbQCMy6Nd5tzYo
SHeAXeURqXepkpOWTbyZ4t11V/Gr3aFjV15Wqno+MO2kuqGN2BudHKum5sSU+daW
UkHuLj2v+8ITmIESUXhHmUxpJUA2uQncd5gLdNbwMsHeSRIMQcbeacycfK/NgoWS
4+mlcFIw3x+iF23J6IGqxzWVn9zkpR9631iyNeaC1BuA1njxrFPkTU+Ymt0+XyQX
Pg/cDFCsv+eEJHEBomgoA0Q9JwxrdfKc15LmOxqvNOMw9SfldagY8rkcwof02bWg
DjTimlK10Vutak84ixmxpC5tvxTahFE67e/TMvljDwvmhoHQmI0ksQufR6VowSMx
/7Clx7fGzt/xcB8q96z6HX3lCUlbbsN5HYQeilM/PKo8VdqSwttaeE6q1AiP5Rl9
V3RTAdvo7R+UAmgB0giY8HpV1KkDBAeS8VFTKVhki8HJ52xzz4OgZmDP9jl2KliG
DTFEseRAny2D5cxi6ZfWAmns31Uz9ve8zHSpsBsDQRsG18w1KjfJcE9QN8uUQQZt
sWLIe2rueqBMLT0EcuqSsEwwyDalcAyTPyNf4o+B1TUqlirgh7RG+sL/4zZgeUV3
mMv9ZJ9uib1k5RJa0LKbwSUBjoY7fVxVPiWKhzFzzrOvOQ0o2qVuAwE0R1ffvjz/
IFozl4RcFGBfAn2JT5CMt1Xle9vgYHLcwkbo3oEfvuehsgj/+Hz2ZkfFEGYQwpy0
Hz3Obx8ybBhaGEfjMgcbXN4kKu6Eyenrt5/HPXPD/FA3fI56iaHkbhS05BdyFUO0
k87o7SqXVR6INIE8TSL/lg2TPBc1waaShuq29zVljsMuoW83wrlznttNrcuI5Fqm
ZnxVp4seVmtcViqrnP9yadB6ezaeUTtPCKe3VikZS5VR7a5eNyR7eFRjaah7DxJC
KrreBuK4TBcJpqkFX47qGtawiJUUSr2JX5DI4/fAQZWeq9kThBIBy9m8SZvSbeh/
ahd+iYhviFW5G+jTEIFSco/WjuOe4LTGq7gQ55HPWw0okuE8uENuBydc0C0yCOSO
B1OIqUfRHfuNdHYSGA57Q7GMuFDNlx7Na+HdPkMKvvepnfQk60q3+YDsJg4+f6u7
9kIN+ZNaIJSuV/8cJvWq4+bz9xVRKV02g4xqcyYYkvbWqvJf8fG1pidr8Rbxdte8
rQwwRqis5Q1G+tYieBE41Hlk6ZsQ4SwYiRGC8czBtfeHa/pTkkRJmdjsscCYh31M
iNfy3QWgSrCz+4piTwK3iDKVRU0Ft86Gc7fWYdoofoowRBuGU6BoryKHemVRVMdd
wRZXz4dgv92t4t9E5Qu8LsYqvwX8K2qaARQFlTLQ5jA9tBWMdJ/lTA9z54m3rvqu
XOVRDvrOwm7F9mMhJ+ZHWh8Q8fMu+zVrAEi888kjzWfwKl8m00Sr/e09Yb6v5fRa
hCYj3tVB9NIjfPqibt+Z1NelfeD7uE6mK9qZpWMZVuvJDP13dv6fNG48M8VjaoJX
4dDZQS+KYuZuPyaiYfjxY3D1/jjeL9IwR7HK1UDOqmuyk1GlRlWDCaRvaA/aeX5W
s49Lc+2d5lxeL4n4pIf6mMSIY8xMgZ8W7+dhCgzfi0LRvm3GmwtvsHOxpYOQMJZT
NruUdJw5EPC1akt89GDkgx0kHBKMfTgMceHdn+evq8fASQojex4GoASSF+PdMUNh
oF6MawrPT+HPAHRafQvcm34OTXL2uV2A+677x6EI3J3nePcsl85YlXm2/CWWx0jU
mu0gXIkDJCWLEnydyZUhZqU8MaDAHTNdckaRucb5SwztUvJ7LOmnD4o4mpK1Q8At
e6PeejvsQxWEZx0rytfigefkNwKFXuUdzB5V4jn7cECvRm0+lbFHW/U8o81aiG/d
oMkqqCQNyZ5xxCLb6TYeMVkI2060KHeptOzPJdmNvB7QLs5Rl8ZotnW+/x71+9sz
LTnGKq2n9/7uQqaZ+RUb2G5tgwJekiQRj5+z+QKUAyKnuJbRNEtpnxHSUFKwobvU
d6nk3KmFBUWzZFAre7LKBppNb0NeqhGUTy61NmGMyHqSompzE9p88Cs7fdVO7o6k
4yD4F9CImaXEqd8XUoKUe5cOi6dzTCsgdxoqbi3Rrn316M/UrZqQkV4XFnn/8l5w
W27ZlGeYDZo81ONlRNxUI6+qiDnHEjVmDjNOpyOJBVB2wWOq/vVVUAiWUKTAsxlC
Jnv2WSVdYXTb/vXj5enYx8oWrB7Pw2j5MMlfJJ++iUkUs2rV6ZKLDTvHN+G2GjbZ
lJLAcv/9p2rU8m1/yVmtpdjYifiqYbX/ReKvxn1N02L+GO/bI0LTGqsmZSc6KCe/
hLN48LkKwtVS/fzRyInGABTA6bSE45AvdHOb8wNGbgh2b7Oc5M5/Y2gYpfwOn+sk
iFaEZ2aQQ8Sk4M0xxL3oMiUDlwNJlnybGAOBBSuLi87GsnxWvIvUrpfehQCjl2Tf
NzIqpYrCPM+0e+yhbRsBIgFStZ+K0UPIW3fCcVfhN5ihRuHuSNWQILHNEDkIZh2X
mPrRXbSBmXpNuV2NwEkErQFS3XXbUjvK7xqn1GSyTx9kLjmqqn4RjAJ3kFZspolD
sDjiVouPXrPONOs4VyvaoU95Tw+JHdHHDx0jJYcZuKyCd+3b4fYM0dP2GwdW5EOV
WyZpJvjOf3QpbCB5SqS5/wuk0+NE+D3zhQij147lXLOSCxw1qTLVd4e3/Sqn/3t+
9mceCfRykJXU/9l+MZFdCu3XgHQw4PDSQ11lxd8bj/iGQeIPQmhQren9vu4I5dVs
eRy/fhkHxhmM5rtmrPb/Qnbyr1B9krAOOmIurh11AiNOYNByLedtB1ruoWqYNmDA
GHLy1hngUuv+zrFbOGeIXqIfxdtf0r+vJ+8TNE7mF4wZZI3sPIyYpIUGhfXO3+d6
UugKZvCS3bF2OWl/5om5y7/WJIV6uRYJfxuA089E+dXW/BVyUdqfhgnUgVqnXHrG
7jQG0GQUOUMSyaAMcOsSuLe//5rPbGfzm3qebjkTnmdos+bwqrtO3t4PVie4OMFi
gQ+sm+uqJP9asuNogYdSZC8wJvuruW45hB3oIEx0EiLeLHEPbt7SMryX77A3jaRo
9RJMYYFm3V1VTmeE9hDCumEgcNezsoC69Q8JMbkF/uhgQX14g37S6aJ9PHDaAiha
kgSOBLUqtt+yZgQLeyQ6y8JH2tm8tbx6na2i8ncIgZa7PgND8lWIerd8kzfJct9s
eAAnDaF/qCyk/2q6UkUYcIQy/PjSZmdHLS2FmXHzjD6ilycoapE+udmDKvY+lIyf
Ezku5zNWVm5bnibm/sEArv9i7uOU67A0MzMhDrrEjGb55j7FpXmL/tCBayfH80Q2
Zrvh5cQGlT9Iu5Ts694yW6GR+jUnS3qrs6Av1cBQN3NTUqMLEc4Y5veOvFTHLGAy
ieIJzDgC6skDX50cXhN9p472Azj1yq27TX7uylbxD+gqfZcwyUd8UxkIAo/C2YBy
XV5rYrcphinCO2sKXcI1Jq1A5F5WJTAaVsk3nhlJ8Q0l60GhfjIHlzIWyZcw2cSo
3V2Q9Wgf375UkMXu6nSvVKKUjBEpmzf0FYndVh70XkBE7vkCvZ9gkWR7auBKHiTJ
UE+gtEQ8SyqEy1ERih0z5Mlu9NJxh3u6Lg3XMeY8bTeBG3ArmWed5yGSyfp3MTJb
TQOOZnrPm6ErKYVJj3cguH6xMPpGJqFWN+NXaErKRo2PUPm5UjJN/hqBy3oie9LQ
vRo/Yxaid3gDYuPoI0KZXj7LgrER7bee1gfARpztiiHnmffwjDQU1zRNpsvo8hUe
qI6t5el3HDNqvlIbFOwcViEoxHB5VVmQkeUVevrLyQXIQsFowAQfReWCYP5yQNt8
B9UmRBoBJEZgB0W9cci4GN6LVDjYK7yJPClIto4WpJW/LRkzuQP1XLHnPPpkfLoe
TSJw76Pvk+s/ihj5imkRn2L8iibW9EkNgme2JlcYLx1WxFyIdSx0iZxAiQx2U/QS
DxJ6UUUDVZcGhIJ2zn21Dy8cX8sl6IRQxLmpLX0q/LZirJ0ap6NTjBgC7qTmAqXR
RaHQdArYW3sgkFspflVtaxIi6q+5GHjWV8Yl7/1jR7Vtf5OWPCqbOaJ6TGyeG8vT
wpYuKwqfc7JgLmiuI4G785DMDfk1c693Kc+K/oiFOPq2tCklwNnGMXPhNlJkOgYa
5c2mewMypx6SDtmzofFesxQwbCPkB28TVWbQNmWLhc+UPRKMxETm9OC/ArxM3oVI
zHSQHXhuh3QNqewLeev26jpviwwU538QnmPOvFyO9sgDKQMw6xU1BZdkxcAyvBko
wLBTfKmNXVkXyZ88H+mTK9HlV+bXhsZbGKPEsL8FcMfDG2zuuDYZUVfByPyvsT3L
HVJEY/bqBkPCzTwAIU2hDhWZ76M19GHRsP/jJC52B4qOHFs9KR4+aVG06y+4jaoQ
n+Nt4ePbN3iXUMncY7+HyuCEBi7MrXIV1kRmAmYp7JYR1OpO5g3n17Y/UvZ+AFtD
3iDURDAk3wcnKeJJwfn9nQsvSrhaVnPkQOseTJJox05NHD2eW4SsbaxdIbAnkRy7
cg8691FjS85AEn4TFOVyE3lllTeVaGnMH9YvVDBoerCu/F8+MFlEDUva1bZhWjwu
wqrzqgO486skDZv370EQpcGfhRM96xewm603v/XDL09LkuCoBO7XXxCFsrgYNbyB
Av4S3lAanCMEC2eqQLi1TYfILWtLexbNWFwwXk4sWZJFALC+4CmghBmqJ5MkKrrV
cFPQo3xB/2AdEj/2BmIcbiix/7pOmXg8KBRJ+NIgjefyHxxhb5GgqfaHbwFN9h0B
QtzOhEqmf9xMs6Z1JLG0fnZAyyHdM4720YnDX9H141lHGLCHXLhvnu94Slabmggb
b6zwVxVwOYxfp+hixXPyA6Cyzx2lYIAgZejSmujBaekaHG3bjY/w7HsDA5R6SxzX
NmFuxfuyi6PoOzOxrlHy9/I0JG02RxVFrNzVbjxDjjWAZMVFG9hVRv5zv+S3QBmg
Pr550yh3s2AnQCn7yHOh0J1qsLi+7WhHzxDxWBgzXam9HqMib+uErDONK/f1pFP9
miVCZRj99E2Pn5wNY26miicPCAl+fdeMkHSWpe+RaIA86bq2ldRK2UVOVI7e2McG
hjSlkM7zhM4qIZqZ3ueMukM6f3bscMnlrnw9E5JtmX+stas9vmsveGOHPGlKa8s8
pVKC8lvnr3gzVCjxCT1s34UKHT/siCTRvc/BJGAWUXeLnVcoz1ieWD4oDWZMktPw
AbsWhCprdNlgVj8hXG88Gd9UDr/DsENp/KbNmoPgwpFzpUZ1ZIZBAvEbyCNyTg86
KgcNkwn3Bn2Ei3XrHX9H0+dkzAZBmg4BYZeZvIoILVk52oUTE7Lqr0y0eYya81Fs
alTeTGLvBoIA6+L6IgbsqOvfFapKYki4VgxpD5WSDw2zLQ0YjhxHSy1YvYbfxoWc
bepVo/v8jp9NmkxiCv8+jyv/4SpdElxK7nlI4Weleq5RYq2cWIoKy/Oawmb7ISC3
kxsjZP2fKzIcC6mECjBx3fHIbuc6XWeVMkbDyHIVmOzSb/L2HORW/9JK+1YIi2Nk
GgWDZdT2K44vlv7/sIJhdvrYDYImCJpf0py0IfmtLoQ+RjAU81i7flVlRKvYgwHH
I/BLyVPvvyRonOTHS6mEJzY8f1Z3OZ44PwWEiYmzEautLnpIaJtyz8f3yTCZ9Ux/
6lSRK0LtW5SPoyJlKtBlPHTVESE1Td4mS8U2LYW2DEHSNiUCK5Y2hRw8/1y2Mo8R
l1IpCmiXi6DxGyKKhrsnxzz4usC5vgPAGsSb0Djn4FGgXpPLY38V5st6wtxKIGR2
BzdY+9W15xl17tD21HhFqFbTYEai38Wm3G+OGoYGPLu70Jdth86qaFXaoMz4Tnia
CuGdR4O1CzdZAiUWk9u5v34dPujFwthZdR7M8tvlMDyEqEFCqSPDU1PWN3MERBjq
BkMT5UCRvuGQSSxArU7uCCV4znR6ANnWUpx6hgnITvFonu/uTnZON80SBXorNSym
yySbNxez5uKvzVuiAew4YXve/sHmQTmW94N+kvKEG2SdeheGbrbkgPI4qJN2FEph
14trwayJ0fzt71mqLZNyYIV3OM5UxmILjHq/jMmVX8Q9dYiq2b+cbOuUMC0oWPOi
JRiKCW5aPFanHy9lErjvPrRuw/by10+mCcwagAFBriEGiYxt6LMxxnsZMRQG8tQK
7Jii57lMrMO1MZl81LvaVOOhI53zLZfrtp+svpau6Z1sVGbAsHQB9aA8sU23RBjc
lwR/FAKtNF9e56SfpNmOq0Yj6a7V1hf6BeLeSH5iSFfio0euNejBH+ufVUifbJC2
tXtfxFndp4KsJfLB+9O6T1EUB3PCUb+3sMmXt57k1Q1+tcGf3B/uY7tfX4Ojwc3z
ErVxNPiRD55ZwndjpJDGW4qCNYn0PMkU47JvfnqYXqpCNk7///zqwGDUvrum2S3Z
0a3cR6HX7/RdVg0MIfnFkJ0yqw75ICLZBpDPtX6QRpiSXMCRAIpJNnWkAP3HB2SW
q7qFv8W83e9IJDIHIOX8NfdRRzUvQz13R1NtLIh0aDMEABFUtsoITKmX3wm9auBi
5Ws7zVAPOx1gKcj0+ROjFZ/gVmbiOZeWycGuTDaexCHAbz4GiPhIuSE4MwoZKrzT
l/C84h7qhze/mhM84wyMFwqq7VUrNL3VmDxO55RvGcjh7nGgdXgMfgg5I/lS4Ddg
asTSn9aoJhjbeYYC2/RObF1YJaMu3DyXaa8G15rxl58M2ahAwVBHh4vYjh00h/1x
Amhh5d12A2dE1UHGqOGRdPr1U/vmKbM4bsdWTRL9GDoBjQVjL1ND9OoupUr0t/5m
i4O2rcIUFIO/ymPJUP6qYGL8MknDtVKwecheY2XtJ5XlsReGxXYC1HyDtm6Zn8Jk
ViMJY5neold655Vo1CGG7KlwsLhMl3rmHHyi/Pl+am8XeoFQWfPpOJHAbFXYQr42
Pt+KZpeu6kjr0xaV+QvrJFFVMXZlv9my3+1D9Mj20fBSkT1Fam/b3Nwf/47r/v0z
zl9SVeG6UZ3x7Wh98+p1YIVizjqm0w1d4r/GKSyvFxh/400yIwHODQksmpgK54KE
IJov4UXK1Cs/lM8VMIbjgocOPujt1lWkiDjp7Oit+8Ir2QVMVwIbYIn4j2QpAQD5
NMbhdu5eRUkpijYcwzpLakd6Uhplx/RfWLfTA+q35dTyRLXnLNxjaYJ3c6NN45UO
jGJt8K1C4zHOZmvSN5tRgCqmsOOQIqNEKeXRlXTTOR5G39zkMQc+P+2nQB9hBVq9
TYdVjAWly+fdPDL0JCFTKygIbgs4INwRp8llpV1640gcmUhsR2evCovB+Lc3z4Wa
T4pW+AW0f5T08nMsKNRDn56s5J1I4/9l3QX0iPiF1qWqceQ+wTuZZWWhI0gSF3Uk
yXgw1jk7lUOZ8Mr39my7vdL6k/VEbSthV6E94OtkqRNJft/DfbX/KIIbTPb9x9ct
AvcWqSmJ4ReU43pZ4jzcLI0+ZMTmiYzA5AOHvhUVku5fNuDCmm9os1TkcJ+vV8TO
NfFFg8KS+CUpgihv3cBqSM2tAsa8UDCurPMTVPS2lAMTc7EGd2P6PSaW4c2Z0yl2
gHV2ZeXUEQYpBsvR2o9HqypOWKoP+bRRujXPtOUuKSPmvYB47ZoN0r7x5fdJuyVX
P+snI6ABlbFFXFu5m2TW5uiI447AJqORWpzv9+JghEyL3r2zE+GW2ynVpXTNhPxT
jTRZxUrb5LWY2vYvz/4QmVNG1xOHU1VGn7MVTn+7633kkZl0D/VSz9lGT75Z1yPP
kJlQTMnNnvT9B+grxPtEO03aIjUeW7kOhg/YrOeNQma9QI3x01HzPqxGJ0g1j8WR
t+JdpjerAeq7NakMqLcJPanylAFDHL4n0J5XOqqNMoT5hxgN6pgq1gmFIwmrqYWV
ee4PTLGk3CKMbrmQXHNb34+P9mQuqiGU9msc4wRme9tNV9wBH+ta9/1jt7gvEJu4
FWRiTxBrilHrdqqBIKhjHldeHh4eUXmvJUQ0VlFbD8a7nmc6P4tjvIl2DZxsyF0e
2xXkVUd0St662jdO/kn9N9pThOPxTNNbg+tU4hrOSX34mS4kyWdv5wJxTpS+MyTW
ySW9aSl1ZGI5WuOoFLRgbxEJELy9ztrDT4XkiNaNs6X51xJMCv5xFiSLeDg3xDWl
bVo4wmFMi3cjBhQx+G8tmSxNMzKUmL47gpKc+iuEcmYSTl86GEfUPQfrtvulSHgp
4JDLDUp2HxbSEggwkwY78TO5qGiCU4a9Yro9zwdCIY4P3g06sLdpXN/PQ42/2kyU
AFVSnY4KUZ3j6Vqty9etpBl8oaYRP+NiQDT2lNiyQHhmTUpwnPjUrY7B1mssBfUz
rkhBRSj3IebCwnmdkVJihAo0uc5Il8YfwdpPXX4iTJZdwqesLYzrcVPxZtoesfuC
zbX9h3qf82XjFrPV6xn/TqgKBiEo8QaPIY6b9Tyz1iBpMDG1kibVjroRt+12cRbC
0w2anMoMDWVViZP0NYTMLeFVzp41KpE7QvcnYvXdejU55PTrtmsB/2fd4HZXb+y6
jeed/HMPbXxiVm/Hh9x++kJ+oJ77G0MDuzVzL1dHr2AgBY3KR5Yg2NAAFQEXT0N0
MlqEnKOwS7mQvlqC3iko7CY3dAY8SAWoo+j1Q0YOyCF9Iyqp6nX0BMSiLwSsF35P
16tNhW7J88qmpZ4Zh6ntFj1qpt08EZJPXteUEm7sohB8Cuq6ccxToyLSohSY8Eog
0n51NoL08G/9TpEkd6/9cKbB/qnih/KGFGakC+YVrU3GdKffkeN6mmNDyhxbeitN
0hGbMQBNlU92mnSVNY9b6/Cy8XywmipCXuCCoobJF1G2cxmbyw5elUccWXovZoAa
1XgoSmqPpkyfiEpvXgSeXQaPuZ/SwZXwTLJmUAAg4bQEpwuVe8kXbhTPo7F3fPuB
geFv7OBovhRf37xW5Rkrmq2GEZvLsgLdvnAK81Udx6vitAUZ3/c4w0gh4mVew5EE
D5jkcT7MQ9Rn9dImujAFsmKykiCQvXBrQ83AvywGPnKGfoOKzTPRLl8xvqRpW+kn
98184G1br/06fnrSTQ/RlHaGngkPsOlHcOmMZ+mqh7prAwa4Hg8+JNK8iL3D3yrK
1j5D62tPBN2dhX6QvFoVc93cVuCsO6AhbFkDGnhM3gErh1F2N4OoxZ4dgWTUBNCO
jH64vRbfSiQsZImNJy7FQMyWQo893GSDbPgVl38vgTtp4MJ3H8IXrqjPuzP9dfpr
2mTWfJpS9pZtswT7RNf2A0p4g+VuzxjeuxB3XtmXBbg+Rgc/YO+vEtk/cKcpWaZu
FarTQYU2KZF3ukBY5VnZWAvKG/j3+e179EGUY6AHvgp7WHHxFbzIuaUuNbEGuRj8
bkqtf/8qSYE1zoCAopzA+RL252Zw+tREkGE0dN6VxvINcU7DVUwM2IRPKnr7HOft
P8YSx4wnX1y53ojsAsb57V3KB9xZgU0wrW3JkoxVi7rlbB6abF57Ghu56IXUxgO3
vy7Z4wRC2TwFzdy/T6+XRKkhq0cEsxKhWXa38Qfjq5S2L8kv8e15UzO1obDvnsGn
FSrt+hSkzD5p12lu9u40/sT6ELf9xuCnawDbR3gUE5TOzSAyhIC8WCLjbIC/O09l
GWs7M0IoyQQjuNXx7ZD+0od9kdO0TtWOfdCAjO9ogLyboWJQgKDG6tQRyDNb4q8M
sLtrdnb1rEe6C4C1xuJyF6F+dcaKtS4TqEe50rPo32tIAx9JSM96joUCGDNZDDVj
3GWWoX2z1wQgWoCucOXb1LWV3KZcBTFOZAA7ycc6w3BnFwelEdTCe/MiSG6DoJK0
N+DBOo0L6XwMj1UD4BBWR9TehhU8zFtw05k9vJ8Fxx8k5BCsXiZgMNTn4rrptoMM
JDMMSGuGSOUbJ+aNtFVD/RhIYC3yqM6sIUQQX3C0fNFqdcNhon5jIT2rcVKGQHAI
bUS/xCgU1ch6INvbZKi+HAjJlslpfQK8bh8+kGqe5mnkMN96TVPFICXzDKab8qUA
zvFS5whClftlz/BR6cc4Z2Am+gH8Q6uji6oUqR+JkvBGXVPm7TDQB6EZT/ygqbPM
3h0k3PHXRYMbTTng4CqmtpqsMybe2H4Tx/EPT2cgby+0xJ08KiogKfbBuLWoMJIO
0k0eTEAEbScY5qmFkgNLEvA9FGHX3CCGhrRUnW7QwmZ0aIBmXl48yw1mfV/J4vDY
L+hcmbLB61Qx6OiwjDs84Kl/YwD4oMln9coyrJTMto9TLqoHi5Tj24b7xYYTa7Ji
vJG7cbH9Js671IUW/kJJwkw6LByDudXPJHNnLAlnDYNBlIJP94Q3XxgLW3zBR0HH
80i13l7nUlBynlnMutjajygdcoidhUWQfN8Vw24/lvsUqYkgR8VXn2S5OzpgfhYO
Hc+6nttYq0WgEjl7AEmPHqegZUUNvP2lHRolNt/YcnrkRMd70FvhnLnT/Zapzeyb
3WCIks+cRbmfqhG/Yy4GOjmqZNOu6c/E1pWspirijeJQRnKob+dNXHdg2PXMmrwM
9ej0JZXx3/5eZOSXBBuUd7WS6ElbsF6FG+OyMr98wU69+HJavvnUU1HSFeVReVKq
3OHCXNT8oykGGZ2lwrLt54/YMilGpwjQI0I2VmZwd57CbssakI8hFmBpa5cQkriK
8S9F6i9vLd4o26Ho9V4+QQEpQoib9UpYTIYfu1o3qt7JcR9aFTQIn9vYtTcyxQIA
7FkIFNvd1YKDoNdKRHfnHp+pl4BvTZEY3CxQbi9mAFNEPQMjPAvFOZ/sNsDvhPSN
+DDQ/r3dArdOiSz2XSTvuoXfM5wTQI3QQqdK68pDJtkItbRSffEf6quE1i/JiFBH
rxje1mUCdTukLWO9i9lCPrz7O7GbvIKJjC/T8Bf27euRH/auwhEezHmOwCEACUZr
+yYv8I8JeVxxmrCboeV+xdUa6LV9nG41epfsCi4BwT88h/TixLT0B9u1G2Da7oqU
F4UXDrZEKlVTiJ+UZ/lZYVaA1dbt6W+4wNwHSxMTzBXLDa+HB8QzFSW3bi149DHt
emhTUItbtNeLuXO/9EGNz8tcsGGCu4ysi6QHaQccigNFdyyMsqpqkFuhSGXMOHYZ
URiqnzGSYKwYAmn9AOrOYWwyvjS7TkxKWy6MnS1Xb5snRW2usFA+cogQaxnd5HE+
KaWCL9f+qlIuKztICY2gBie00TqVct8+Jrx/XbV3iKRquR0dhkuJxxNBU4lcYWnR
Z/WjKYdAvsHeuV+YvRc6n1wcVflfmbM6JO0F0Cfa3uAShf4OIu7moqHpEEJiCDef
Yit4RDGWePQqnOzsV0eBTDOWf5Y7up40CSzsMIvlYqzGt8QAcmMStrAtlC5P+bXQ
0mm3g9x1mV6JEj+9i4fi/Lfrpnine7Riw59AJWYzi4QLQtphoP7MJSFAdca4gvbm
CaWdUPGJTaUrSi09iO0AVmwkvuPCOsGO70mA+azXghqiNQGNvV/YIPRQXs9dyjIq
HoPK9l6YSPEersnyHIFApCzmF4QsvhWWp7kaPuxLzpVFcFL4J1OACiUXMiI1Sr4E
pruODDxODDZ6wl8vido7Nmddr4AHEcCZqBEtI067WHZDE0VP/rnvrtFmCLxuMVHx
7p6f738d0EJaB97iygQkY4MapBr1tPVWeze7/nBokPR9Jpi0aunu/RPTIim5UhLQ
ZMZSS1fSzatC3IlIS8GNZ6OZeOH7U52cg2GDhifrqAi8C9M+uB/LF1n4+qalP7e/
pWp9ShlOTv7a1BqWyeLaN6MAfe5/UEGphV7yqbp3k5ZDzilj1+SutxlG/WKg6WC4
Kx94KdNYZD4lWEsymIH2zpE+QUqxBsFOD59iZS1wLYeKe4+racXvMuSlq6PGfkmK
1NJ20KDj/i1BEQ3fNlKNBBtYoxiQApZ6WT2pMVka5frshMu1xOJVUlEGOW0dgoTW
AvYridwIj6pibWBSOwqyN7Bh+DfNcqbImizt6zAV6bJUnNzRk4bwn9j3FFs2DOXO
1NpKgBzJTATsdbHD424efDvUzDFThQAWsiG0NW9PwpHndJEasti/yaBTSyY9MYXW
oSNJojz8tmowe81Ia59YTQ==
`pragma protect end_protected
