// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Q1YdDLhwK7WoWNw9UkzhxspAxsDscftP9Jav/LvV8BaIhfE4F3sEkU3BrsgL3O5r
0DOwxLOLQtKUC21+RAlm69YjrvG4B7Ecr4NDlGc46jZbn9FHlydlUsih3Mn08Fwj
MjY3C244l7uPFFmkTdXYR+yPtSzHYKbydCmGQaQ5fgc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8288)
da1INOg/s+yfbXPew+JLCLNBaORFuKvDSUPVI2zfRU5E/uxLQC/88plVZIBEYGsr
NnOgXfgFKF+auYe1tOSeDPhHQU2Tr0YZXYUY5V54UWNEJ5QH8/3vd1B1BonH+uef
byjFG6p9pCsK29c/8IoIsRjVSeMoUboSAldMDgSpkyzxo3017OULV/DYaBKsUbm/
C9wsZPaxhpklKWqmy3uwE4DHWxDBBprvPYWKS3szOdwNe2Bi8FXMbcvWQ0rgRpSK
JjgbEFs9kBGsRZ+PFyahFOgDrIE/DlKj7+PncUT8ppJZmLuPjLFYgAkmYsBT9p9L
bmvwGCoWzCzJFVQ+6ylAiVSbdwxC85Qf6FzesSmZgi9deV9gvQJwsuPvGzI+Hgfn
2kdh3aY+aEpuIkbEY6KEeiQVr47In+nPkN6QRWZgDuOBh//WCYV+mP8eKVXyZYMA
haZRWgSMDopLvHzxSW856OzVe7DDlf6QFOhWLZsatsMcxqccikusQAQ6nZcs4fnU
1ZFnqJp69r1pUNRm5bxPkP49WkpGATUZcoCMzFmCtcvlbPIxFIu6bxBIPFfOGyVK
gmFm5hxFVZhXsqD6yb42KsD9+N8Rs99reiHx+rAwZYreHHoVG0tn+sqv8FBvcnIx
LhOipZ2sqwL6lQhsn0ko0eZtUprHs3QGZLwc5SwWD6Sf5O/SSZNGdmBp7Qkbj5ys
FmHbZ/siov/pR+UezJFA/5SBLd+uQWjaxQHP88Tcl5Q1YXr1uQ+wPyzK52dvru/b
LTZEq3J2ZQtF6EIX4MhE9Xe3w6B8flItLVKDI1JiSsjDUqS3/XsS5+d758mrOV0l
yZmrCxDoHeM8NCsFSap3sCA/5sC3MGI79TbmbsGbzuYG72ShiZJGh1dUzznokBAg
REbLubNUlwU21EG4Kat95XZ1uIa0E1R4kLRTWy9oxKKpmTKga3EwZrAgAR9p4zDj
QaFnUwykIOW0YG14knLVMKZIXMcSJD86ic42otoIIwo42VHwPE/thtTaHwX5Ornf
IRWcFIWbPe8w6z01GIEjM65Fb0iev/f+X36voBEAW6XlXgB/Lgs1njdtPSXPJxtZ
e/6CJ0Y6elFcCg+/AC02AWWxrMwMPW4Fxrd0xMOYzr54Zdy2dLvrZ1bls6BYzlNn
fTRgqwtpJsMLcUXVTyXwy24lM/hNuhx3ObpED99Q3Q7Y9ixCTk+Q9PFmTAUkN8aE
j6OOS26JMnf9RWauWA/LskTv8jxcoPGzLt73pz64+Nr97kVv62HZL1YLkBtsbwLP
ck029YKhyOnYlP7I/HH5Ztezj8XIoSDlBGcWp4QhmM+GgzR/wHE0xNEIb1n6pHyN
So4ByqXfGohsO0UfdeHcCZ67TthAaexBxhacUQBnEksi1G+mOW8vknmau0YjxGGP
T2XYal3wY93kFIKXBKP3pb3IJIFNC6AY4A8HE/BrhBftEV8brQ1/1s/RHpErWG5Y
gCzRWU2osVQNSM+ni9ETKZEAJdg0RygAdQkUonK+jOm4iodqpcsr9zFq3XmghAYa
1p4/ajYdascENVX50PxkfvEjsLC8XjoKIkdqITb10yRhI0Aimc63eh/2SKlr3ph0
HjCyt9rVMqnfIh2o4IqmO869kaBorr9AehlpUqn4AT5Ad1TOBqgq5W3gLq5ECr8A
sZvvrlWgwepesBt/av4eem2UgDijvJ+49FCb2FG/9wwtTmT69MdpSV1JrTuPZK13
nPPBYoJJwRPVvfkbdSevgulS4PWIpr4BIXq6vdtV8QaL+3rSJYnAUjGP/pV3Fd8I
UK/tUmcXHqyGsQ37mNuXgzLc1hJZEv9lcRswnhLuUzrIDdDR9iYu1J/l8YkTefUe
ZGtfBX8Irsw1xPMnkD0Ww8Zt4ur90nIhR7euPbRFWFMyNSLau+SE4cxmJ9aLxgFt
Zw7x6hFna84IARjzwFWvsLo37jkLOOvBx7hrz/LOkre7TAqxExSfKIJyLESvkPpL
dKvjI476jRdXkD9JftdTiSyl0eX/vS4xOSrU8Da1hx9CdPnCrB8iFWu69KSIrJ15
G/1Ox9okNTyZOQa5rz9q1tGa2WzWgNiuo+Xcoa/EMn+c116jJyMCM5vkACiwWULy
SwXHibqWmHaBV33xlnDsNIuoh4sJQnlN4f5NO38E7CMN1gYACpQmr0NKJcuyfD5z
IL3/jjEUzuoviZfuXSx0/igxJ1HMKuHvYJQXEeAIHdMiMpO3ejHB8H13Sv5A17m+
k8ILlVHgbYTWDnnm2DJpq0/Nop2y0FlbIn4kOJqx4NQZv1R5ZqD/GNsVG9puL22X
Xre36IUDJod+ZtztpmmldROnuPjDjRDXkrLP1deJ0/QywoPq417XLNy+dnB0w1rL
HT7VjgeAigM8tK95dFdJPV9toyBjvusYIvyR3QGqU/ktiGXY8qOi5kTcusKGOZbh
ohP9+doCm/+YGstAfSDBh1VJPxgFWllnKxS/G0u1fPFGZrF76gIrbdmrBcBfLF3A
Dg4dXYN/CNOg99f8pQ62kdtdBCc4W4Gw1QozoBarDLGUdWVD26LMF4aac2OAswix
tkbah6czxNLwiJCQlDUu+IumMgnu+HmVZ/c0GaNJCIT+J5DdQk18Zsz4u0hWrPbC
a9gZZW7cdVeMoqyCzufkST9tIUUTGoSPNh4wNxO0ZbZnvvWQcIDWxYG1bTukqJbc
HweidlgIbeLdFy6TipA924IwpRFJyvYgM5YYVyvS2iJ/ZWKCa7D3WUSuGB6fUxJV
HNU/MAzf93YdTHPNo+SRMPQj+/h+3o5N+3XdcUJr3nOWjg5PlL3IMyP+5rI9Lzav
6ec3Ux3gSPZj3AHBHc9hzMKV4d1NfaPrEFxM/pYhe82rWi5YPl7Hc+Zt8BrAHxfR
HZgknFhgsF54+EG9qNckLIwFzqOySNImWSjIldbzsStfw96QDUBE0ktsvIOD6GRJ
X/Bjl4xaVE4CttQDI3Gw61U6VtnOVWIn36qNRPDY0cLwEAcksm7AzDZVqoIiANFc
DwdLtHfYvJeh++W3XBHs1GqKJjdATG1PO+YIerA1JAwHa6hrVkIniHqqXNT36bdi
nGL5CiLKpNX6nyTviayzm26TwYlYHVoGhJb0Hv6/GWmrHWqjv5P4b5o+tpQS5bAR
6BTogE6Qy6QVdPVWDZqXX/jjQhyZ97dZ6W0TuRPEi750rOrgOow4EY5mE3XWSXO0
s090lDymFlbnTe+hLiL3TiR21OvhTB6/AUJpplZ+FhA+SrWKezRC3ckkPW0adBYP
AfaqIJwHZ/sXs2FtcCxpRfm2RXdtgbuy7yL6626Msb6FnVm0tt696RkvCtW1Fbfw
KeQZz3kcHOeurd9LCc1C6XmV5ja/lhYaLiHLKg8gkhNmFCkCRDHsqYCbXVuJy+JH
0Hz4V8q4YoZMKUWfgkG0ciY/WdCF9P3oTqe7gm+lyeDEKAfMmV5Ox/ykzIlDV5Ye
tZx6R82X5mn79iLCBCg+YZLUOBMi/Po1124jh09eBKZJC5lfw8YQ6D4/kTM94Obm
//MDlDfYP111TVKTG6WsPbuxOirfkFNyhJrNqUk+BbS7+CzPqTuKuJeKd+O283wE
oUhHypwv1O/Ac9AXwrNzyFwgIbx/opjGIYHR8PsS/98TCpM/PfXNVFy9odr5ecPE
/6x1OXc5b7p6Lb52uDVHeChm5jHMyf9oKwHJ+aHt1pCxwkan/5KNScWk/4F2TPng
R4w+Glw1IQKxMiEEaT/YL8V/8lH7n64ccwSDl8pUhV3vgQrtd0mURit0Y/6oZls4
mKKLsarmKI5OHV/IMHrpLsYPaT90CrY9ftqH/k3qHtLJwA94k0EDGopWXcYUit1E
9pQa9Q2y1VGlP7iI7LkQC/t0CmHNI7+qEWRQtLqBrQoXCyUrtXHWwmd1sctj5W2i
merXKU+pb3caMKvDU6V1S6oLTJmstniGJqvxWGduhQk5jP4zLPeMc1j1DnWhNt9K
D+m2FThe2B+4OwmaoH0JXHYwrsXz7Kxv2e1dKCwrdTo5UzjDDBEPzH5k2Rk819ez
qvZNK8HEgpUCUM7yIKpTRbVaZDoodghcaP2J3QJRMVrKYd1f/zm5se2LVBzIp0qv
a37Z7YTnxsgYXAdoV/+QeUMoZaKnT64qqAWhV33WtwgvMF58Ttv4rUe+x75YVEdx
S9qEvKq9e0e8BHaaEJL/ABopMIP6n2DEt5OUeBzDfJllv5EvnIJSoBFKrsH772J2
zeuziLee95ty4cgd6s3ozYdaqgxwSkrF9yhokKYfYiFKzgjW2VfD2KLSQ9ruFQQ4
uUUD+ssKCLg9ojscWbFHuS1NdE214miFXN2TXO2ES3ZJ9aeDLq1jI5YemadzigTI
azCGaSVyZXDJ+K/NgjywQscTBBS9jMxkUnGqrQ+h3dxIROoCUqH9/nZivSoMtvBG
QgiItNbFWfF/UkSzM7i8PFh42FaCTS7HlbUzGsHX29AN82it7jt7yO1nwhvRyLrn
8ngDhQAP2bFcELXTlX4yAeydZKZ+wqbotC+6AEeYtZM9xCt2kNKYA9FJGgdbVmQN
BbJGxpq7Hdb7jbFZvzIv7JhIDW9z1GHOi2PeiRw9OzUfbhoyGaSwVqLUDi06eEgJ
tOy8n4ij8tzQ5LjI8Q8DWsUyD82KrIAY+nCOzhjN1ZYquccJB3S6JUF+iVOYn2ne
8O50SM0Iseq+wR61Gaho7GNcs5CWZRSyeYpHV1IK3/L30jr5YOdgdsRKOyF7lpTU
dokRIv+dShIvLgJ9H9cN0IrOo/6yUd0qRPiJ8yGLIxh9W6FcU23E9eXpXIIcjwn9
NUVuN9qt6KP3XMTIENAPKoATFKZg7KQmJVRA+ZSQ4nQOK1eu8ZnDDaI7dwWWD8Vx
Uv3Pdqq6UXVkZLn2Rcw7TtCkYwoqkVtoBWWS/VCDaFjdJpER8CAQa2F0JR8AysEr
/g1/e4MCry8yQYUwWh5fZVAcV3t7fi7qfXAKDAO1mbcwFtgiw8Zoq9if2/SJ9obD
Wmx7kZqW3HBGF+6pPGkfIic2EVuHqkF5/7i4v+XA2PDyIYN6JWGz4hGZQZUcOxFf
dcr/R8JsD+4xLR98VHBg2GBguzOG8o9i6uPHNRJXSTPL1zhQ0qDjWcJ/Bw+dZ5Qz
m18CCyJsOEwIyittwdj+TTwzEo/7pdvZSYlX/90kCvx8tdm3RgPmxVRgq4TzeMmC
mswn1iwoHpFrW4xNvPTBE9X/FbU2cVvwJ0DfmiWCiMiUxtQI6kgsBndY21cEJsp7
z0YsZ3/g1P1C4UkvN5XZ5Y2TwiHoG/5NZySP/67goNK06I6bCOZwmj3qx3NgeCjj
K1hvwm4TAPOsSsFKEq8AyVAemfbF7hBtJ8kH6tDUeLjx6SKYDZTGGw1UFx9+dL/R
Gj79OT1xC0+XWmSkIoqKSrQiT8t3VB6VVT0oOWOOtDYNIqrnsuGg68S2q1HwkhIN
oMGts5bZiOnzB4kaZ/RpEuY0ubGEseUDk265xVC3TnT3wJz3//dNK76wx2rZz5qK
eBfiAdi0Lex0uTKswkuqlvdIIs+GlhG/5hsCG6EoUKrC2vwPPT8ZHbBuBtoGKhZc
F885D2uX+7pvV+qploStlEUIPyPSeMyUpIqDGte3wyg4SvN3RYeId6cEYETV25Dp
T4t+hpSvey7FIehHLzX7ol3Ar/1YkaarMJSQ39SRHl+xWwDEx0aKyRiTIdp4R4kj
kaH4k+DS3Njc+FbMZvupucB1xinN4eqyjQGP/NkvyMlFSK4aS/xemEd8dot0V0dR
gF9MBR7XwRYaL1qTHWFejr+HfggfskEAUe9gwR0UeKVX2ULw08zwQJ88HKKQoiif
Xb8m7UCO3G535KHjjSqXIZbz1HAS3ykC7jCoOiNTXopLEohkKCKHhXINphuVKuEU
I+P9jTaKoTkLs8moveAvPuoY47nfStLpvJcuEzoqBG2O41Od/uwC+ok7crx3Y8I0
JrDMfwrMogf/l4So8csnCPKaDc7UEpS5p/fijr5fYuyDZ1pEcYm6GjiIxXfoYm2w
9Xwe840Am1Y15XiRcCC8QmNXJP5AspRWAAKCMWefKfFRZR+2nlpHKMS6dC975mx8
5xruCtCvilMc178mZXIZf0xgZNjDao7JUiumShHhw7mJ/t6uz+Af6hc22n9QS4z3
IGssOJL7B5aXAocPqxYUXdg9Wn4mKya06ZWkt4Ke3HZnVVO2skPKLLuTC1jUmfGq
QdPKV0TnjTAmFUWs442DLmtqm1pmK7A8rabkTcXi3ATPSU0hWKuPurFvRyNz/TN+
34aDwpgZsJxWoHGjWAE9qGnws2EBSzusl8fP6+G7mTngnt0yyq8CMADAi5jCbnJ0
ufDu1uSVypWSMOSTpRRe/947jccAnu03VUethvySb1s+38pfaJ0h2JZOdQt6jbSK
9XhlIs5iKLBMbO3dbqkz1JIjKPGfxeNjb9IusCMhGG4pcbeG1e8CnSptYouWZUNm
oqMcJxE/TlsFUBnMCcdYGFEScRx8cEMeiZfNVfsqV6kbWZFHiPpcjq0VBKzT7JF5
Jscm38rbgT7SqcPf32VOCfA51Zad2X5HlLqfadjuc5q8XoYJJYUekEuPY0C/UkS4
dPBW5e1ZBh8m3mrMv5odlKdDK0vgg7GyXKeyiN7fzSoR0Pq3kNBm2Y4WtOgj40YL
kN4e0lw//vjs60FZ/tuTLB5p7ovfoEBjBKnlV8WeERuSzkmdMLGiVCofu+mRE5PI
PgoAJnSJaj/A1L7Bd6JRSvJJ05EEtc9URWUogNWTZ/ido2mz3nQV955G5sYg6ntz
VL58woJdOK4AxnmB/MIGm6IVDh52BgrLKY85mf30rKyi1hQdGhgbvlzKVcUaVWkf
o5h5R6ocEm8wYj/vtFtqUP1Uajg/Rh1RM7uG5BJa9RkleOyix/wc+ORyGGZxARLk
pzeTxkHPHoiKtIey0Bn5ioAyoOx3T1A8c6Lz7KtfQ84/wEcMxYaJcOID9rsOG8gn
g2b1DtiWR9sR+S62gEYh4cnaFuaZCCff+izVkwqHw0u1Sjdfvl5TMuxOGX8khaaQ
LVGsWTlCn5iVobwCdOuQpY7rkIED6asGkzK3DPW0cg10MEVCZ4/XHc53qW2gp1dL
wIgh4S/Zn9x5TmrFX/0yzBWSfKA2gBsMIXL3fQe0Sv1a0MUwQy0BLI26h5mCQwTr
p1ZA9ZDG2RDBoabkghMn+WJ8bURyGq8KgLlFyrslIs39Uj6DYTzcp4bpw/7iTH/J
GliZVe33TKZZRWFMEg/8KfvH4WzrMAZRMvxEeFjxhOE1rqiLxI7qBHddsgseEx0u
iUdfPgQ8ujVFs3HFTIUGH4QNS7sdmIiipUr/uI5ezJZJa6Hbi68482MWfkaGICZX
DSB6cjGfvB4beoZ6DfRWlAAjGas8DBLQ83H3Ul5P04C+qnFbWpC5Cwz/Sc+u2i5F
xkS7PL08Nb217YSqVUAzSh4XSFbg6BT0/QrTiqLMBEO+slI65PrRQBkm44IjXY8c
f4hTWXuZ8OXuR/1r/dpE6QQMUGRT20a1NGwW6QzLUCC/cyekdqqF1M+t1QYpH4nf
6eVWQur9ORGyxUzt2hwNb85XV3jfjMuNlaYwBRBsov8vsnHepuniaoqVTx5ShhrI
FjEUAbBq+Aw9jiidE+KIZ7AzLJBBckYFlylILlgsFf85LYFPxHKdceKJYj+nr8Vk
UJiFTMiFgtJOVPhNd32cK98q1MJfEp4wVk51d8sr7OGX2CyXm2jlVZbnEIG5bLlJ
UY3dzDP72sI+rH7E0vOQu7yIg6ZYn74WJtHDk/S42nT+psqvvfV0j9EWUOsdAO09
exbdSjxRciZr2CY22GSgt0JPN1J5vR0GnBmHBR/oqVLtu/1HTVs0mKeCRbxrA9hw
FlN1BpWSsf+4U9JSkqWA1uwBoAYGdS8N2jVjPlZr3eYjmMM3HJgs39Exmbdv/8ow
Ap9S0fyS7aFiwOSdJG55W8w1P5b5SyH0BuePrcB1H5JwiRKZ7EnmkZq8DZA36iud
7J5+wo1kMKPQMymccGthBvmx5hCKNU67Vlfy/WLRDV1DoarZfMkasoVSkJ+Piad1
aYvepGASekBKXTfZmDUToh13QeMluXQa1PI3GqwNUyt0Ff+pJ8BKgFruP4Z9X7wP
gla4a0JnWhmP5u8PT3dYKmUam1zz56JYR4A53xwvWLWPci0oRqI6BLHn5LVNLgs9
kvnoRDyYKNK1QLiNpZKWtfCZK+6KLQ2uCD1ICRiPJrfitRes/Nb7ljyeBRQHuhaX
K8YNpvtAJLtAkvD4dwV10HaIEFbJdBtjSwcAUNZDDTKqUS6VMbZCfOqpPxxk+Lj/
kGXJyK207F9T9TK8leH/dlblYtqbQxYWVYUIRUAEMtX5BblX5JoeLq+wdKHj2i2L
h0ps6WyLpkcEA5kgTHbHjxDkDseJFQSWsB5JATaUu6a3Ic74InSZUxf4e6C+3XWJ
DVAO6ZjlxMgdUzJmVdRGvxqLbmisJ5vWVI/sWqoCHBk9eEd4o4MTsC45VUD2c+6N
TvcgitvhVkMQcByHfsiZEPSY260Tp1UNsUh2lxsFJlbU117UuFuyH6Q/6mZez6LO
02+teLzanCer5e0K6gTIXiw4nYWE1ubU1Ccdg4PaPa8hZ87pOAh+s+qy7keHKHRZ
uqhJxA6NEV1P4+Qw3Kby7BzYvduH2j4Kg+aE6dM6o3tjnmbEB7zGLhNo3cbHBXrj
/qeqFcwUA6N099u0zkKDG8ovJ5CLndaOGXNTBtaCEXhGzKpdQ/278mpzg3j7tr5w
UVCaaMoz+jjsQ5pDGGicYCyEwMRAOd6reBx+gdETZSPt+9mSi/6hXeiWDh99hyq6
1oCDnmVThJTQu3HmPypgxuzo5kxVMEkSo7AHlbQwZPfOSTBaGxdGV0y0NZ7JZFE/
kdIbZLHp5WmZnNSK8xP7fiN2wIAI/uda1/iwSMDxTm3rzkKXfRdFHosnM0AJjAgE
vOvHRHUhmTMVw7QrSDdjazYkH6P5PmATZz7B+GJbkvHmRe6N99ExXWkqXH+w08xO
Q5Xjc7P/EU0URv5HhB9WzvY99aTNGpenQ5sL/JvvXLDyuhn75sgtZi8IvjX0MEPL
8f/4jTh9azl7qgo1MeSJqwwU/daK8a95kn07LJRsb3D+ejVcEnYUV4j12Ihgx6x2
Gv26QbqEu1LQRi0+OiD49/zppodiWSmSu6oNOBlO0w/o3Mjz9MzRN4bk7Fe1kAIS
sYjmTu0hue5pwoeA5ktBXJXF0N/Eyf8zILs02o24FgT/tAQA3wOBLvYtkan5+1R7
4emFEbvJmi4SY2Gcddunb1bjGBNcKgIjY2bwjNzBs6cGTzN9KuMFDqEHxuh5GYz/
ghiF42O1XUqe+5viLHOTUHGbhhKGqeLN1bDh+d0U1L2ouyS03tBDQKjfB2ZEtS0S
TqzC6aH0IslXxHMIN9ANl29d75C6eX3EaBfnuKzAY8FfYo17jR6mNvCIvB3KuZjJ
pCslCGfFBQ9uep8ohqma2nxGpuRhXzXZy2fI3J4thbs3b3IlC0C1UM8Npd5Kvrth
QKM2cGIo5d6PK2zDXNTAbGiC7ksKfxw6PmnlxE+q9STXfXj4hlTErVbxA6BrbmeU
3lPShsvFpSPk2JS7Xk+LkhH7eSJwwtRaRw51pXaneYUvAP8T4uhRMBF7U3S5uA4C
KV8DO2q8k/70wg1lQi4CglSizf60Y9rMw0aKCQhY9+ApKB/jXAhA89Fbk+9IXwno
BtZ/iuX13fzPjVoxM9kokmIAYJ/Hr3C3C2cIpb8I2Dp1JTLjH9PQ6cz3s5s70XLY
lpGfE31eSuzq+8lTMjLClpaN6s/tf0ccGphv/Hw56pdyYCMhou8wrc69isvPkj2k
yr+4D5KbuRzodBjT3av8wrru1UHzL8K/Q/XmK1duCVK8SbgBlNqIdPwjSfnRUsw+
XqF59NrlRrykuhpZo6cVE1nRskdsXRN0P8fc2L3dynTRPA0IwIigMMb8C+ZLGi1d
vLazoPQ2OOQDqb80skZtbD2iHEnGnaXi6MVwgkwKT+e9I0iJ8sqIas6+N/bg4Hiv
m+81BGy4Vd9SmAYh7zt3iF3Yyp0jJHqv1BJrTtSQzogNJS1V1c2pPvdO9QpafRcp
yqhxqJjWUW8AIm5isUnaNgCbbgUaVtC3wRjFl6EhxGJw23lX7zoFtkz8wldFyVXc
bHIl01D4zgXo2h+VAiCeHxeLtecARioEg2sT984JLrFNTPG2JJ+4IDdllRZBcChz
CUET+g3zv73xO7Uno+sCYTu9GN3P2itKZ7VPXT9dVn+2JIAXOJpFWEvDRNjo1nAV
nOiJLOMGfPbtiC92/YniNh/YCw520I8NekhiNyIBxvFxHYnXGY65cU5CoeUUoQ3Y
BMb/mwSCMD2JuHhw+fDw6YA74T7RXf0h8R1BlFYxjLGWuWFF7lbiTauzOldp0YbT
PoyVF+mi+eF1PC0WH8f3CWlUHgNwq4Mtv/gJXHYYV1kCvvJhdHJ5TY1NQdJ1PwpG
/Ei88lTRtJgQcAwb8nNwg7qftaAJ6Hy8+RFRSTU481Oh5/ZQNT9WR4u3tkBKoCHk
reXRoF5/Dds33ZlfRbUv8mEGlNX6PVmdYzfqQMcPmURh8jkqUDJHrSlaO6TPwyKM
JtcuDbWG+R1Ec11CB7Qk0GjHrGqqsOk7H62srm1q4HhZvISBtB05iLT9Phy952JE
gW8njQ3rQT/CTZAE8ZgxcVf812ymoM7aLMMyKJ5KprAFVEScZHf816kLMARBb/cl
0MDsWlLljzuZ0FrlBUFe8nthSUsZFobHtthDrWIQkgQ6pwq+IRMJPLApLZYF1lcY
dXn2lbruHDfH/sKczfAwvDxpJID+RIaIWwIYdLC5dAwNQ4k46MPzUajbWO/CpbpF
z8RRtbVh/jktnbmJ6ctXmeOtcvxdEfVAWGqHcE3oH29xGJDTAUn0X95xTkIQQ2MD
zO92Yg1Ja5eX83ZCmopQJw2lemmD+zyrz2oxUSPY+3wA/S8dOGYuBtuhnk6ye8AM
gXs/ORPa/F/YcSkyCgM4dWDtajtmOscYaAOwSXijWgs=
`pragma protect end_protected
