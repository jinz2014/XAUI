// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cByGC2rXZKZk7lWuOLEFlVHqTyKSgkbnDyZf7UYpQt7ozphCbwPtlIPxssxQIijG
n8BcCIN0vMy3tHR+kzWFS5w9JLF2VdOxAmfnuYuMganIQYIjy0H8SeoTZfUkSjKV
HFkamLDuJAOeM9mXX2iuXuB/iHp3I/JCIWDi4imy7d4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3328)
G5ryAAUZTaBO8R9gKqHQcpzvSdRf2X03v7KPIYHlA0bP6TzsRFN3Hs1+AwhcRWfW
TobZmx3Zw14N4q+G6EdpHZmHgYNwLsyHA7WUIUisRml0yubWW3wOeTi2bTwpxS5Q
cgqqsPov8WBaWqOKlpQLKemjNptM1znbCMuhdopepu+NIJRqSA6GQSDPdG+zKxOY
+nJkstRI/VIWLdQcywmuC/zX5rguNpmN1bqlzXh30KZgXjw6GCBAdlvXp06T2f6J
cEiVtMRYcg4Gi6KwhqamiVzA3kBy1aTMewEXGPiOifdtIWJPc4wmgUs3/FUxZYhk
Znj//NGAbYTyh8zIcNnWYzLX+Io33eCTvlCSDoISm1Ex33BHbyLRr+zJpmw6Wcc+
XFadeCUoTkmQ3AZ/jLOYDjY04w+0xTBkeyHmATE26x19F8CDv9euF7ib/QLdy2ux
1FJD/1bAMuZi09brIIUdUhJq6fLFgFFVfifx7VLt38PWsCfXFkHLmFM5E0JjA7FT
tM7NpYaY2fMkDxqSsmkLRn9U23mrFCieIvCRytduUU1KHBex17M88jd1gvFTJGUM
tTCd67bW6zZgl1isror7L+fh+wigv8+hEnuRx6hCFH1NhFID2l2ErkuqIMbG+iFA
lbwtWvf1/rg9euk+DfDY/g6L17Z3VHev7VlJilpSjeK4tq4RlFBZ4DiknQaF1Ta8
Dl5Z9Y8R1u/Qei99Yz3urZ/jw0iE9PRRKUavVaCaHpvTcai3k2HiRE4TtY2tzgMC
5T1Hkoej8zkIn5oOCSvObNBj4nB8mwXJFJqpvDKpmv4K53RFt71Jdu+Fjc308wNj
Ap8St13G3cQabrViGyF/aN73AoanND/Irg4r1RA4rHvUppnqXRg84A9xMkCKxHUS
H6/VaVDO7r+95EPGjf5j+hOm9x+ARvmGyGtI8VA5g4CVU9KAyxv/jRuCRMXLVmCU
tlCWq+Bte/6dkL6WEyWVAzyanLLrN3wohSZikLNyJ5l4/OMfs/rHK2tapfqLGkG1
jMtavsG7jGnHatPTavF6H8boq5ZHk3GOa0YWtW0gs1x/Z3f2+vRZ2SkW3FSg/kLC
CEWaHOSTkDjLp8dJ6N55CeQplYPgI+7QmB/l/PjoWa/8u8myzZIIDo+jBlZlLOmp
1PXvPpmX5VZneCOBculOnjqemflLlt/oyivqOiVqohYQWfEMTK77NObakYQASKH3
yfQyeJU39NjZ/uizwwwmEWWCZUg+2mExYYDObJbKINhpVaN3F3OK+F7ufTrUWCZQ
DoCu2tWL5m96efjEopAzJbsuu1HY/eTl4FmXUrPPEjIhKd9LH/5+QVvrFVFXEaV+
mFvblWuFpDgZ2vCFjB5w1x9idQ2yWh+hhvijQHdjD2PI+tZlrU/ckYRWySeVKNEK
6HsltIrGnLhJNSsTdcyJx2ErjRRtcIyhCw5XhnarfPuzShOYfR720PEZleki3b3X
nXa1lMLjWZE0jnBJvfllZKnupN9gHJZ2CBlvhNctjVuZS+306BFxsVo/nqfrk3Oc
SvZxK2ZAIGN/TywBP/RVd6gQpNAbpeR+7PlV9Nuw7CjI9DO9ZIGyLzRxq9CKUDvo
tHe1T+3nj8Q4cJEaoEcGYUuus/zSTiB/FmK/4sepWhci3FgXmD1Pg8dGasiycPci
Er8UJ0f1Xl8FwRLKjhdk1FNt/gFcrmvzNyrCYWO6zWMwGAwWC7luxQ1fbNJ8WfeS
CbXEd428W+Va/zL91E8l1fgWXK7K+7WXXucYL6N2PuuzUrx2TxfIB9zhX3zBI2KG
7eT0ypaWmEA5mNJMRKfcHcTMSqIcYKBXutk+m9N9R8TOvtJ50HhrB/a5b7ekBWqJ
gE3QIkGls6Dxaz7cNqZLZ38gVjpOgId9G+WxjjXXfDWll9YKUcKChZ+Strac2isY
5hL/AQl9660F0yGXNIClpize3QzoWuMk+dv4h7OMx7sivzY1ygkYjCH4DvzVftyb
mNVIeGe83ZJ7tTJ58tha1hC8lJjTxjLgf30L96EhRck3BgYGuqzFxgIeTb32gNHW
Pi/sKlrNUpb/IbZzeUqsV+PHjL7Rg5d97TXXqt7+8vGvk1mcO+cd0wEZJVzU6JW1
d7A9Er6EWOoTIXNBo63nS57U3pQvrtBfeKhpHSVVytnxE/tWLuOxORLiAjA5ybKg
2FVPgB0UmINO5NNU6WajLJeaNperX5jKoX2mX43xQ/C2TSDDO368/K0PmnXbDWVo
sUbfdl75TTR/ZXw6mnY9hm5nmmiRD0ulmArnn/oYNhASnqpZCTaZK9bJnoDY+JOC
JMxFgRPx1gKYbvbfC92UBn6qWYY8eRvbu5FMmwNMEUhz2f1qv7FTw6aoUCoOUCQK
oTM4gNM0GygaeHcMvhtxBf28IjhjDcR4pz/+4G0EJ3PaAzSRcWSNKidBYxN1/bct
VkYY/wisaTXqjwbZkZcOkweUJolZLYJZ6F3W9SD6tXPpIo+dwfwvPxCwjWRfOHQS
5kcS7rL8lIIGvxf3Ph5KfhEKp7FUwqL4TASkMUhB/p/QUcsbhLF12jq5HxcwQDkg
tiu6iCMcYNNHqU4kDf2OUESPAV8LCtPjLZG5Sao+p37RKGoS2oL8s+LMYyS0IpMB
lZRclEYVSKZwp8j6qsaSIJ+ThAr78UqJb7aZ1ZW2qsmgJcAeZrfcQqLSZGD0ApRY
y8PAtBpAxvoqyHmMxdnAaKnS1kefew8FM25sp7/AX7N3facmcJNNo5jisJpxUHqN
H/ulVS5Mk4nfy5mLXwsjWa/TC2Yhq2YI3GSz4Z/+RyPpY7QnK/qrA2A3XhSprsGj
t9Yo06UKuoefo3/LaCJckKYuSbnSfymbVLLU7EbbrPA6r7hW1rO/kLdpO9I9FXn7
6BAQ2LDjB02Mnt6GNLHB/AtMXvOZWoousmDSTWI+/fyVJOVuDe6nl8AtkTdlZHsQ
2w/DW+9W9DZZd1Eq67/F+B8L54pYaMMGGuiwlGXRcj/p5Y01Ws8UGsehVms211dg
nfiWkas24bx5mB7k0qAz25UFTuxkPwlv/kg4p7aig1Hhj02+NgJk6HGRdGXrXOVn
9zpW+dpJolwIDAIL4L/Kq38QNnCFL/XO+j4LxBqnfEOL/onOutS+wI48bwLN4BMb
sKB9Kl3gP6fUuhfGqeYMxtX1kad1ttyQ+TsUvwYQrsrprrj4g8g7s5qyFnvcm5IQ
ybQJ1lGxs4lb0/iZ9llq3Qybw/QpprlofEEeFe+BzaqdRfgQDTVqfQKF4P9Dlnsn
f9cu1O0odxdgewEL/jOjKm66aosXzliB6Zitf+tbRiLA/mFeNWH3v9Z4d1Eiwx/J
951GXOflPdrt08xGQNo8X2yWyes/RE4IoQDWDl6wsU0b6fqo27Z9EXAhuID/UnWA
tdohbe2pVglYRF6aZzAonj03tzhn9VMZaQmwBLlbHUEx2wfEXYJH9B4CzCzp6wP6
aZJGQxGe4QYEkTOVB8kTt70PE5E/tArp8guaZ57vi9IRs+rwKHUnvGs3ADPNTqLM
iE2I8Lzl222V1S7TUiNOFnnjzMafxRn39Apo9WY7oc1DH1XaDg3IwvDCGj/MrTKw
a6mjvZcECCAhYfz0dqvpK9Xre/hEVWOS/LULIX6taq64g4g8yLxDisbSmdK/gPa5
We9FVyTF4VUni6Xzlqh6wPVmT+jzYiMljvysJSvoabn8FLUOfHuEKCxTNmucAFlQ
T2mTH6Sz2DEpuyZZlkcfLEBPgZOyCYfGRY5iAd5S51zjba/Xd+PHVcrjPtBpXXPe
56ofIAidnqnjxtkZ4BpGTPgY6IA9lpa0/4LeoPmHQfSzMFrS+0Ae7Fz5OkTbQJgr
n2qidJi2lvYcz7cB+DkSg6PDcku9Chi7VR5MoHBpfdf82GCypW7uCK02RL2rHij2
2GW6cHPii0sgdS/+qQC3y5tKFV7KdQmBHRCY3o9lU80G3qZivBzxg3HNvs60tTE7
qIKKeqJMdNLEnSWlHSYUrgRE3zNgd52QkWqkjTG7+LKUhSvdHi6RqtESt+BV+Koq
GxdNj3LutqlR1DHOvzjrXWYeHVn5ZfW24rIIY/1YFLsT/f6qEWofCo/JKTp6w40o
hezy2n2iBmZdc/PdRCf90M+/kRdbHRenCr4HWoZhbNXJbjt2U7l5XifYc8KhdRYV
P4OHzNFHiZRC78j/UQE7ZmFJjXrnNPtWyZzI7O3bXqqRwkrri0/CHLSLbgwp1Euf
XayHfYEChArJDL9OUGomdwthj6TN/snlj7Du55LXDnZLNuYAqwCGi6w0CLRBVuPc
gEMEBiU66Fq4LgzhJnwrbhuI4NGUoHh6wd0wJr5r6lYtk9z0v0JVClzSpwfAHgDO
i+J8jT9wlCOjYiYCInLU9sJPHd9vYzZRVBgioTw4mWtD6m+/6+P6C9uoky6vq5XP
5afJLHE8kbg3K9vW6wDmiw==
`pragma protect end_protected
