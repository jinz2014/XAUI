// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FU6CFR0phQ/xdHWIvjuwt6SCmNRDJ5vgU55hxnn8R5lZ0ct3n/yiV/hl89/Cnf0S
POC1520mZeXAXSkDN2xwKpBO0sK7q61bSLrLswyhw308iC8OwokyRFB8ogpck+67
nIREsL8FOawiIYNjgRjHAt6ZQ0dVJS6pXBK93E5yZzs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
653KjRTLldWSUu/Nwz2XgGB4Px0tm9xgERHy564R9VLWtKclNQc38xX6zteS0ea+
hxD064CUArt8Bb6yXc5hCOM6kZ3NASOmsObiU6xJ0F784889Fgw3xdm4JjTBoWy0
5vFtySmrxBa6uGvxo4ebx9SHyUfcC4BQX5t27VyozhmScov6kM84HnMFMqtM2wNA
ogg2H9hjLh+SoTNPesko8ZDcOlTzwNgwR8DPAAdNsX076wAAbHWwcf4FF7AEmYrT
rLLgSnaoEYj7scEfrgyEX45WsSNdDzz5lHn1y0+dgIX6q3nCSKLZj+V8DzdEdfFX
Wi766K0pJTeDhmzNxnO1x70sYAsG1ZsgpjGfHfhUzgaIK/MfI6Hy5nQZPdBv/ALD
Wmgzb/SXfkIPzirSLNJ0ddf2b7jHdJIFILramekhZwPgfARiuXA8fbJzVJz0mMal
lVCyuyewSX6KMM/6i6HW2q2cKW/tc7V49EdgzVaX4LyZgYlBvDkLVzMI2kuQRGz5
r8ruz7PzAYkTvTXJkPG+XbZA1DgK5EpevVWSVhyitDPW35Qk9h+SwUbI2lV2cw34
evA0o1fluzbIqC03IH5VqgTqfsgEsEo4BcW0ZaDaYV1mErp6QWkvSysG23OFZG+R
MsYSjI03euQHkdKJQof4ktNPxP6+sfxJ9wraPD+Uclim6OTTNmNz03vqephWUQKk
BsAowCfmAunSpkhye2t8GwU7G/yBh/0ImcedczH3OQkhiB/nylK9affNd9p9v16d
Ptgns/Y5t9OIPexm+4yDPHt4j4JPP8iL9lB8E2pMRIMlors2Lua1e3Aenr7p1TXQ
e+SuF3praTKvq7kUPctncrvAU9qZ0NsU5fDKW7zv5SY8FoV1cAMEf+Og6o5Hu2Ek
hPsa9VmJaUYYpJhSpf4empclQmjZB95Wc0D2MAVLlebTVj38S1bJN0kvGMhkyMGw
Ol0zksfHt0qEMOGtH9MyoLQIFYIm8FQ7kI+dm7vygF0dvvmAHgT+lsgB7rQq8KXc
cz+v4IQLYj0BHKVSbcxZvbVLfBdqBIIPB97ofnw2+fE/D30GFoHAjnpb5UOAfTgZ
Sx16JcAn9/SOPTBa2Y14ct/QRc1UXqj+K6/CG6i2/irPgaRc+eO7veRa9JMnauNA
7tbGj32Z4f9AO2Bk/C5Y0tNAZJYDtR/u3r8nZqZnr5xSQuCRxKlZU4/8HS8T2O+T
omWSa5FBrPPTzwnLBh9d5BfOmHNyyiiLrZH9eCXGcoI+5s2UWtX8v3megYKRPL4h
ld2/C6d6DyYa+XGbuC3JwRaDh7l4+mOZATk5rtDrSHRDSRANeqZoz2K25/iQVEPI
jmjUcUNhHhF442RXzFdc7ZY6EXur3URtDQGhcttZ8B4r86rLrK5A3RX3GFBf0lG+
scjqEjyQlZeLYuNyWwv1NR93Jua2r+y7a8/G+zpdJkP5Re+5DyTt9oqriL57IkJR
FTY48pGz7vNnr4rR6tXqImItHqs1gkS6WdBsLT+lwTUjgRUf5Rm+mZQgqKLh4DWk
aMnaJmoZtNQg8PLnDh3Z5pA4dWJufiQaILbcif217hBo5Y9hyEHsOVa1aHhtJEyf
vVEZAtYbmyrYLbzyBISBJmJIOta6nUaqFUNwoigqSlOcktzlTvKsKKoYoIrnAJQo
AoC0pnLCtxc6wrT3VvtJVqbyYxDwcOeyJItyTjv9/GbRQuxZP+pgNPW/ME6ue6G/
N6JSr7Brdpl34cIF5ksLqVsGFjo73zqwQBYDIi9SbA873GtwYgQ0wJmXljDJyuxv
ZG+ORTWaz8Cr1SNiOjqndvlqBRU9juM+3Squvrxv+bUpgHhffpMUt/8sSol4ZiSv
ycjN9sj+fC5S0laF3nATGt1cEuJdAK/JN0jjiCEahuchYOZ9aGp+tc8IEFF8qiaL
4s8nU881Ytibp3hD3CLq9LvbP39t5mrQIwCKdjnyLQSiX6eJ9xm6ZublEE4rQ6BS
7WSx7n2kH5KuUcNYaH/wBRSv9YKs6A/HtMl8xMBlHUu13UHRHRMDGsEbfVp9tYL1
Q6PSteDz2NgQT/U8TiI0zUIqT4OImjPjXewXCKQ/ZpIZ32qagPUn6U85BDbab6nj
q6ehVShfpTLigam22jNDJjs0DbMC4AiJGYJ92N+obmeSGnFCOn6LXnXLL2wPhJmp
BY7QW7PIf1EcfDfDlhs/JpX6weanxSB7ihqNcc7mGDNrHkqb25ucONotaM/98Z+8
19CaisFdXhW/1d0dcKGuNkIReF9AV6utaEC0jlEGOZneyEkYFPv+6Q24NwlGzvKl
q6UPM8FpOnE9ZNSRTYKaXrCGvbj0eDe4ThUD89W/7dkGcLS83C2oSdDeCs1j1gaC
XpaL0vhMHkqTlcCvyEkD+llvDckwl0H/ZAgBsQfbMKcuhWH96w5bWpagmMolV4rw
UP6DDDpddOsMbHDKHsYzyTYoD/ajhbnkfOHQaMsYiuDxTMILrnwuxCpg3pTxJF+N
qiIOCSe7NiJ2QOyrtfDSlYRDCF+JrfYOAD6mxczXZfvq/6QjX54i7JfU7uxwWRQM
vn+edOmx7qJlVuVuqTsAVaWqHLMdKkipfqOBQy2hUV76D3Oh1aWSGJtTFgkPv+8W
sYwa1NaoMvKB69M1GosiE/EPzAg78E+aLKLryR6Ly5tD+/2qkjMQoBUrR92gAByL
pwO2xnh53QC1HQ9Ow9j4KlMEcp+a8NiLrsBYcioOdAuZoMGaPzmYeMkGDdO6xUqu
x9V4XfW4cL1EgA4IBX8RdMtZ/DA/R4LlAyRQL98u23fJF7mml22tuzo6I64QB2lU
7SqewKbvArJndk5JceBxnqkGLCDeMblmfAlXiBvDv0AomcRPo+6QB+WcMPuvypdT
LkSjzUQ3s0E2M+p9gRZgLKBUURR14mCFWG/iDEcJgWXDvm6fys7Z3vTGTx2Vo7I5
cLIThQrEtBhdjbIi6qjUl//oJqmsrY3RE2hiWq5Rmbxdmj5hkQkZ+2Es1HDU5pZn
GSaHOWKDVNRE9n+/pydZzS8rNlLN/yQFt/IAUViieORyvP01shnBQpgPjRxPDO7o
yQvfCCqD8pXCyIp9+Hg42S3TJUS0ZyD4OCCNbidbDe6CFNTkswPBTHpGMqjnZrwm
5zyBnxqKAFvuHUHNDu6Zc3LXZn4+6QEZEWXY39pE2TsIbE8W4g8w+izQy67NqUja
mtuIjJ9Ax3CWDAf0l92N65lgiUPH6thpZf+LkOWKk62d0mHEdkTtiiVLFOs62oz7
wpn2fNx+GtwtUnQaF9yy3GIX9CfyMqA4bLJICG0XXBKnlYJ1gKIGl8XTj4U4V13f
NheViaAZ9Yhi0tWck0c3vLtyRm6TALL+PUC6W1eg/HZaxpES0qGAxeQ3PerJ9Pv6
3tTc1SBsttgMmDpFPlvPQLzZEYqWqy8lV1l85KxZJJ0Ix0A8ZicE3MrdhBqzdmGz
yiFUCXRnRhUYA45K0VAM1Fn34vzXMG47zDzagqlHhSsLXcGcnBFPSNKmnAbsDnAU
W04J9J5/XqZvJ9onQ7sTmUS5y80HTF6rx18lemRzTwOlmFlyzq+wY43VPILj9e3F
yDxEhYHFLyDhHrUFVYELsbF2rOMn738fOrugBdKB2gD1/4gTY8pE7TT/ntzDDbK8
kl/pX5TUGjjDePPkIsDgUcZB9J4w6jdJV011eXuVmbF8TtfSVXsUMzcML9sEVhwN
rmU0lEjDmIAhDU2vKIh+L98wnuiCXp/xdHWcZitDOd3zjfBqh8scyCO8sxqcKNKm
0/Wx+9T62wJ1BMGJUBayYADdaerL1wd7WPgUCVdzyr6/tEUl0RhcXHVHKWUYkyjZ
2QSaBPGqn0jP5rAApTJ6vMZLxh7SS3/idlLEF4SX4Ot0dWRZyuTL9gk8PcjEexef
BoyW+WakQSMqtLMMHX7rnG1zezrHEZvIy2MvZnR/ti6HFxD/tL3ZR+ZUGXY0OMKG
vyPY9wyUtytBYLTd3aWi8hP7qTW26Mcix9BAYXqyhmaCUsX2i7T2hMsP9Nclrq4i
iYESX66e8i3s1YM0s/ulow==
`pragma protect end_protected
