// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MeEluPulL9n+YW1Jxxl1x2XEOXsXDE2KSyVB8uiuuFBZpySqCJH4qB3z/yIigsYn
9lHWNeow8Zuu51yTDnFXFFf2RwGwXfVTQq23+aueiOmAwJeMZrurB8uO8/RC8RgI
V640LwtaBHiEZWjV0yZMlEPgHDdLU/h7YhAjaw1N4vA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6480)
dpEXDPP7e90fFw6EyX/iyDjTG15D31LRk1DuHv+3aFEKBTkNhEJSGvI79NUROL/s
CbvRjia/B2LCeF7AfIA9vLI1pIclthiFpUytVvJbw4yKBnlTyv1g/28Hz5dxwI7m
FwX6nGPKfr0TezsJtogDPF8HxJazns1Ve5L5VhzP0MBwZJ+bsM/+PTN8m+htLtwn
JJQ2FVf50/IlUUUNnds95iWckPOtMvWu4nlC7cQvR6b1bJLA/FcH+RwlVZ3bYipG
NaWiiLJie1Ybgg4nN5e+D1qIEcF17wsUb9jJXvepiNlXsXWKLLN+Mgi7CMwdp2ex
LUpSGra4BAnAbLzpRrvms1qTGaRUvaxe+B4xpiDBsa5Oir6doE7+czRmo474ngDs
RhNTweBasQTZzfZvzXO8HLeK9QThqOzVqRWGOS278ZEQbz5z9RtLcbaEwSK3YMuG
8/J0H8JwhKQ/wvIa1SKG1uTcqQM3vIJSJDNJM+k7IMoFDfFK+2k8DIQUGqhUBK7n
oYStPqnDMp+gOX7SzFFd7sxnB2N6z/ySgaf5yIETYbq4GC70b9Q7B3vMuX1QqknO
7ET0iourMh6ua2m5qqJjrjJGW9IhFODzU0aEHj9fCEVzjskJn7YZPq8h2xEW4Pb2
2zTyNSi9ECQxvQhPwN+kDI5DiUsPEwGFijANiMz+woYzApGA2CZXjPUfpWcJSMK3
E/6T5CdIGVct4RWSydAN4TE6rQBIAC095V/LQW7ID5CL3z7QoMM5QiaRq2RQBpgI
mabrLG50qwt50sFTl4ZlPsq7n23ha+UkBPHA88rmOYcLKNtMdDuAp/CqIblaY/c5
xspz0szYA4B5cJINeug4wbIi/uueeFmmpMcVby7XJQ1xh6YpgiQZdlYA8RsxQEMd
HZYxewuw4wicwJ7CJIFUAcsZqsLMUtzeij4BVy1LaUpSFTp6HPexuZXtYFZIBsaQ
1T3L2986uJdoyW1PSrsao0y5ipNO2Y6WwL0q2S34gCA2NetRr76phQcR8ORvqcEW
QTOUXcMV6M8X4GQHiXuKknuST0VbL/JRzN1CBdwx1lF1PbzlJmKSoAOtlMe3aHCu
JGGEvtM0tEFu+479eC18MTy2AT78H9tOa1EzybhwwoFzXxjQKdEJGCmbgA6yjozT
9IxCZoP6ak+QMiJl8AEsYJ/osOLV44k/Vm8uP6T028a2zsaFeUW6G4kfoCbgtYex
PcgLAotCPI0EofnVvtAqfVSH8Fg6xstmCOukaTSF6/P8F/eXQrx2JkFlZFzo5aT2
AoFjrI5AZO6TTkfIM8PHWRSIjOwnUivwLwLtJpvlBLk2xBPnuiqVExLJQND9LxJq
Z8ewwj1pHZuXmLFlyAzL68/nDIRWhnIA16rpe9WJDxP+EFKovnMlm9Vfljcl7W8D
iO4d++/VMlcixkDkt9+kAwfzZHhPZTdSRwi51hshiG0oXyEUXLBJd3IaJ8flfkzl
rBQtNNCCEhbHGNNO7Eg1Hnk/l1r45awEpoA+ahGJV63kS9xtiSL685BM2Y5rVdRG
ZKzDCzGMIdiog/k0qSW2tb9f3S7ostKMNNXcL0/CiLoK/NqbuoIaIwddgGYpoCZY
XcODYUOfw5yhuAJJR6rsFBR+py3UQCXvF8WKAqR0ZodTmn9+5Bn4vpixZKIiav00
/iSDAyKM5h5LqxJsstzJpP0WQ0FXCc2SEvB5lm+7ta11xVkBM4Pkit5fvszU7mM6
xQFowTlImQ6LsA7FMnxGNYA+rz2JY88lhcBOjfKGzN5tZM0mEiRyEC2DPQM8iWtg
fJtEe/rFd2cvUrvAFFmFMPZ3a5VLtcGTeCGiMsiBZETzpTM2+nZK3Mbd7QCT7Wv0
+T+nsfXyjXDBTGvdjGKSD5kKtJBY5jPmdmLp4XJ4BOIeFJ9Cy6M1onfU8up+hztZ
pJbvuaFvDfesqkxnbEcLIWkgnLOa84F8LJUfIx7Szxyy5KV8ufT80vp2Tm4C0T+P
XpeGq4XDGjbECJ0CwHSDwdKqwUp0zfIN7lipWDvWHeZ7aQ9gBN8sAcld0Fc4wvq8
QpFIQQ/rIKX3ukOZQ8y5R03cl6yD13VNuALqtFbozIvMN+gZslJkmSwfUw2EeDp9
Q6BNAAEhyNS1a7KOisK2Vg2u3AOJ4Gm2xxhP8xIqLQhGAVfEUfWvRhYuA95IifDI
eYTmjt3L547jZztcdF0RRKRiDh1KfY+O5vkqgezDM8YWyFAv8nP5GA4CJNHMKNlB
zkUdEXbiBCn4p4Uo8xyarBQUXMLk1cxCdELi8nfOsAIW3tTGnRPGErucI+nhwiGs
XVkFZDh0AoKblWN0LXlhryvdSGBFdrCTDdzwROAwkGPjgBRymyMDxF1HOrE1ip+X
0++umI+TDdGpfu4HVb8kby3XGWZNfgamlu/7OTevCvDnT9au3HaZYlvRh5OAUqAt
KfZ7iEOgfi+RJOsyORHiMPDyF5HE3roodhcRTZ82S5xykksixI04/9uf/ej52bo5
NC4W4fIbDpYSKqVPE4aSsBsaR6VTB/3IpKFbP5oJWNu3T1aEVQI6Uxskl+EBP/ms
oPUJbeyLwe3uNJs8nx5sENfAiAhYzOJnZvtzLXA2wQ9XqUaUZnijxrrNnC7/krdn
7OA4L0lFnjXNulpxvvfezbEUTOXiJG1FvMoXy9I+1mpjiZor4vidPMi/7BuwEGqo
HdrAjpHtYB0bCpU3Zs1CdbkQMFmJCKoJsNMlw5j+sxI2zI4I+PvYN8kwFRRYsJO1
uwyXLymLOBLFYBFGjPhETOWZHJleBC48Fcr8HMXrrgXn6XxrHBDmdqDXwWoeL4JC
r+Xm67szjR8uz5/7OUfB2kK/s6+8yXbgMVPTtp9qYQXyYTXyj9EXEmYG3jE11M0R
O57D8nDgDVSWu5gfkEQdCg2lMmIvy5JJjjntJYnn1UTQTDez3nEUDVzTP3RMODqO
931Ay46oBeiJB8m+5XY/O5FRNaRBi21DPFA8NF3Bhm86IimGKJ6avLjFvfr/qVkR
cGyvwwDydCzXvQa2oZme1by6voH781nCnKU5wbv6xoLTBdctcwRbLZT2HE2JiG4Q
YPFcVuGq/ogTKTmZtB/35UIx6Csad+zXCdbmCb+Zo+q2JPDXJTwZzkJreyqkF9Ws
VAUIP84OMRNLQIHjQXVdEbJSBO1VygJLfnvGQ0HOUZomkMI/GJoc5MJfSrAPG1E/
YKalXBti+lKxzApavb/yBnbBTmXKo2tjm2Q0pCEfNTnwaAF97RGoeLocopc0v1vB
SpHbjDnXSnnGgNsXRQeslOANBXkT5ng2sWaN//UY3X6HZj8I9GYveF47T3TKU+h5
oipw1p8PMPOfdHP2E5sNavPhaVIhGFE1WyQIfxvp5zVdLwmcdwe49L+6mCo8xHOh
t8rrJBuJkD8EiqcjQQGNMrheQ0KDH2nL2JHx6M122ei9L3I6DxL/yNWEOdAJic18
5l4Q60J1Wy5mIYSAM/QcLd1aybqThhwOC/Rum/3/i4O2e+eKyaJvbVQYnZWmIkeE
SGSbXBoHTCeNpv1CgLQRpWxW0ZyXOqUE4fQRiRFCFpKRjf9GhSncDy+7Ejq7mkmu
hYV/IMn87XAkiPW6tLn5y+F62F+t+59aDA8KmwM9IRQTtEKnfev/1LFxl04Ydy3K
raQ7G1WI9/FBCAWD9ALX0vLfmY2sxGZ4HG897Oil/0N72yy7XBKp8A119UJQgKZn
BEvBtBDfZ24fvIBJZvZVMf5whNga4BMkBLDlPWJJScgrOWkd1m/AktChUcjSNS6i
irMb1zK0vKgbQigbsj76XxFwOSnqBqZ/Kx7RcuZsHpLoR9xJuTOiIYBXEhUW9l44
j+EcM09Ke/l6K2lZ1Oe5RShr/OlLwKBzT1Lvyv0Oyy18bBpmkLf75y+jBeJAHapq
dA69N3mXS9tHnS9hA0sxv7yNQHUs7IhCopup85bnjs+yMVI2O20R35ZKZ3hJIy0t
MCF3AQOr8bbtfNog/QBKSImyFjTL0Ub/rlDoVSifagjTE81mMnPjGQxS0fziyi7y
gBfARJEnOMYY2k3k+o1ip9QeyOkTuDC98SsBfOJYz5OIdgDfRdvsg6b2lzg6LSss
qxr6oN6xzVtvDXPx0Ct/QXlUTRt8WaYDT1L612pbo7tcWWWa6BUH8v6ybfCkvHfa
85As676xCR6LKxsJlBsmsuiRCHY+FsUPoRoV4WNy0M8HHFKxQTzB3zEFN3I3YlcI
1G1tSh5wlW8HI2NrU7Cef9nGkPSAulqW8VAARcXYce0WdLrkLxNizfDeKRkPlIH2
/D5W5pQlPoloKcB9tkCuzeGQ/Xoj9x1HYVeje/Pd4tj2Um2HZrrqNO74wicWZE4S
pUK2cISp7snrWP7xROM0qldgMKxwNEoMlSSodjrn9k0KvfW6SCOrDFiFyq4cIolB
jvhLjHWFeOXIh4H5FPykQJ2i5VNCT86D3iKArYrj1oqHq280Trt7Gpi6jFHzZmNj
cXeNCANHD7WkHzTWwiEFEAHpo7+rtBDjDEfkpmDiO04wTdUsveA0DKWSVngRxjPZ
xOek4NNN++vCwplL7UdW5ESqHxRqd83cmeoSKkcm/I/vM4tpckiqHj0vJurNF0gP
9nezWWkBhbv/DT+901V2nc0cYZ9Bp9nrrfT1/2qOhWhk43NER6946bNWVP99BOl8
PWLRcmino6X3WC4ySKV8GxhP1mwxz2U8b7/rqWZ+l2g2PsvV2nehaZn9DizlfGUl
xViA1yI4bWNLxCZnWRVDpau3WVHQcYoZ3xB63utj+phgC+h+VYnYxgeMHzInMqcS
ry0BJ2dFWjTTk2tx1dm3fWccZWETSTgdJV0saKDyHcJ63KSFvjuuF8eilSLMjN1i
qNKtRTHw4pVaTpR0b1RB+RPEff2z26ISIZoUlT9U1/KUbNawFoP7UqBt/lKTzouR
bi5hTjde0kbq6ApVRA8LiZa8eqMdUfD4XoEyZu/T6+aYCzfot6fiMNFYneiF8rco
5VeHbrF/BWR/bZngNeJo/puBoQaimdSgppSjCMSqHX1fdYptXcP7Mvdwl/9cupP7
T9f5YtFyQYM33UbcUzI6HLZS+Y5GzsmCzH4sk8aY8XhZxIxkmqJ8k61dCFoVhMoX
YbNxtPNpPJ/mZ9bl7YflNWTHLYfxVRiMrM630iY2ImPzOtWBu5TorK5JeNVTqS3m
NrgSHqEB5LOIlQRbESRHqoKS1bb5oxlaNqV6q+6mo/wwc/hXBfcvF4/6f7h+CSIg
wEx026vbGF4QoLxVxnZzsrs9/dx4wSDGyB6p8TVseSidIERvRv4nNOB3qFWf7zup
RqxW/vzbjf+uADkYLhS6EV54D3rrgj/1od0tWKxyljR3coOWKxbECb4QgEybAuA6
valVJyIjeErSZV8s11Lgt6dxhZ8mIPlzDZyJupEroczBwqowGHF+LuKnF7VTpGxO
AfDl/w2mWhIFKSgARnavaMFLO5l0oiZwPdCYl6F5klvKSBlTNTMaTzvYvQ2axj/J
Teoyi0w0rFsyAkOfNKuSZA9iCc8XR1Qldl+x4jRB/aM7hKxPqIBTF0BiP6dKzSIb
/aF9533M+Yp9LeY7mtGoS2EYZVyNo5cAvPORtetls9ygSuMgsvm/vfepaixdYyG/
cl2oWV6b+aIlUEE62xsTAoRJrehk3kGtMnAJs6poRuTSnmzcjmcDwiiw2w3J3lqD
5t+7yHG8AJka0hQLJTq6klay0+JqGyCOXFc9HXGylt9pQB2hunbo1ZVMT0cEZyny
VQdW2lQH8y/YfoPe06GhUkQGK1B+U9eFmMe4RDLCIojvfIAEc1BDdzjWn6O7US/i
6oNcrZrQuWDAINpg9l2adqsyl6+liqII7wBt9sIL8qM1Zowh/1b5TajRE/TFpish
boprVRAVWOrzyct/OyE+3sK6aeebJRhSZTVTTHz6ksDT6yaRRb20XBo+PPn8K+mo
aaJ8XyuqLqEPdwYii8R5aE24pJ3PyL2DCGx3y3Nj7YMyveieatqIvXD+FCLFrkW9
5jMZgtn4YKjW/LKeR1U6/8zoi1/5HEbxIhxdSYqbN5ki79NBRrquhTF9xLyamIWL
0qn8z38H45u2iamCWqbKXs5/SyhMCj3pdLzCWy9aRh22BmgcYnRJa6tuuUgooLYa
3g0IjVSDawN8k+qQ12PVYhNcHYGA/41Lqbmpbf3nGuiQDfcDXvevZJRFsPaA4Qe9
A+aCtAA3ZE1jTSwiJQQKVDNcpeKHvea6/5l+fMh23h8+PdpOFms7gHhzgUupnQb4
yZbIgk9+YOp+u5tGA9aT/7/JiC4YA6blOOl+Ta06DLuueLKshc/HJTEx7QxsXNsq
asKViPe+oN+VRzTZ1APFS+EQvNFq8zeDgrF8Mwau8M575t/km+Jo1AYomWAkIUvu
Lzm+HPktjKx5b+grEKqepil+/vlj3WawnzZO6iAxEsjMo1zt/REqLl2BGZsMrzFF
BVHQd5slnLohZt+CfaUltcw0AX5Y1m5QTJhXU2Dwex6TRkDImo29NuZgVdpWIpm+
RKiLEwDqpJtoNHUnZ+1zUh58tUDCdDkUDDKEN5AvV1wx3omg9nbtjWFwJF4YTNQJ
dBFPZ5vKXPCD31HY4sxfG0G//TNBgTYf21e38VoODbbc3gH7tOAGZsVrkVhL6WYC
PcEOmburne4OFbBMumQp6hlouGcr3rytLBwMwY3E4yX+I8txAS0yFLDxdmzSrRRG
TUGH/rIjIEbBKPaKNQ9/WLgZpZufPU3pD4VgmZXvhmK2akH1/TwLeOzfF+0c+tmT
eh6nSyiBJatP4b5JyO1OqwndyL7tv375WiTCg+ZphcAGSMQ0+1LcllQnW6d4wONd
QDJzHAWrwjvWxBXuTRbY2EDGYYdBoLCCodFjwPYbOA+xRFKJKIcX+qsmynZ4gKX2
JSJ2jPe53MUrneFD8r8Km/2V7V82bqkurBSbVwNLp2U6MX8UEd+Qp6wmx0AaZ/cX
DBalG3h3rKIF3rqYedezIVuDaX23NhXrhqFustl87nFLiTuqjgCsL1jqZevHJPjl
65Cr0bcgr7/gVppk/kawUygqh0dqP48xOc40MSXZEo1QyRSzCdWcdHRgZEV40IAO
dC7IH+tYCP7jlzPpN0HTA6LrSoLcVWnKwQElrXjTP9T46v+ifKkF5WgsfmMP2gXN
QBOtwMDyJGRSa6i8qqdtFRytD2PJgfSN1aQPQPpuAnYHPZVphMHCEvQGqrOpjUs9
SeuJrFNKWu3ImjIeLtgesyguLmc/I4ikGK3qn/MHLVb43VwHlaM7snGG84I9ibL3
8+PHG6uoVSJNwl3GAFza0dSsVlWvcSiHrQSzFlvS1oX+ukE04bZL4oeIoyHLMIfM
9Zc1eWEEZ1deJlBFwnxC18IQk6oZPu7Cr2zFdJX+62Fahx5nXydILB51coztHswe
J/Lt6Hj0QeMFR4HcWPOmr+/Iho2WSYYGmPdLRDPEdqA5N0WlcOlR/XT1LiJWPAmm
kDRlSGmcCNB7lwSLBQF+on6dLBKwZ08M3c7qj+fTWvZSCqvpKIMH0lo/Cuc2Al6d
q9Za5mhzG/iPAsAsOEvlKh8q6l38CC5FQHRoWjAndlhxpFbLuTRuawBFxxYR5RPh
0//R9Pxv5fWy0UzGXBS7eozsfk2QGBz+NdqbB6DXRcIlc6Ea/Co8UlKVQbw/Zq+T
P4EoxqJKicoRT6vjeVc7s4w0J4aQ53Vn4neVPtFu/KT8JyAZ3WgGWVgwwDqj2gjW
CrUiRZ+LrNfYgxOLbl7jxSkJiNNjpwjpdAABS9FeZWFEXigRweSwmZ31vc1g/M8X
V9hf6Eai/7qEnDT1RaFLC1TYFMyfnJGRUkfRbPZCHqzMe+8+78YtsuSASMpSWbI7
R/4qXQ/w9OQWuOUoPpMwkXGyHeNChQx6tpPfgcv/NJM0BKsvka3Sohfi2J3NyYme
P646eIs3Js5K7agxTzqmiuChE2LoCDA20wQ7GFZtno6y5XKL4TkUHG8b+dPZ6oFd
i5mcGJOsXeZwP0ik3Zsjk4tqxqk3c+Gag2Y/1vSNeiJamSKssMMK+iWF9RyLkw78
jILg0kmU1+44+aw27q0Ov09eSW7uQZfq04RUemn3H62U2NwroiE8EG8xwOUVp/+4
iWi198/v3q+aB8c3+Ck6pvMvoIs7X9m2Lgs+xnwa4YYTIv8QkSe22SYAzRr6wb4H
Lct/QDhXl7x7L86tn6J16nZ58iXGge8XSJ23+Z6wEF50QaQ6/XxxCnKl4uFqBZj9
rnBmkV7quoIangQ7/XrHaTS52OyKrNt31BYQ+quWG02k8i9800wQYZbY/e4FKta3
+TIx92ku9epkU+Mlan4Dup/4wCZ7AMYFnlciqhsRE+MAGA0185/tegMNoWc7yUD5
1xB83gWUMN7U5lFegp6s/8+9cHrJjh/Rx9ukhRPwEaMIrykE87ngNjkD3MtkZ/WI
KzGWBTN9I6FEWVCTjxAzALSQWA9wqFW9UnHpd2Q1onNThDbFoVqMkag4gQq8AVxB
fR9n2hDKTHECJ8///Lj13mlxveillmkB4PqNbJBNU/46LW72P2oBrD3aiD7ViqPQ
/xAGUAkvPdX2bd7E4YLX5Bq5Jf7MWiNyS5dctNJK3/V6Ff/rzxU90WcL/5rPqg9C
`pragma protect end_protected
