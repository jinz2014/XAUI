// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:31 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IgQenmPxqFQk8pbJ/UQmfVHioFKstClQf5jI0zJvWAX0zCjd/O1njr8dZ3wEm1fH
dOynBPWPoYa/Oa0sojVta+2xAw0av4mHKnS/Anu5h3rdr7GnfKBn+vD8wRCz8ROf
ng+1m5KYcp264mXKdlW3a6/SaCVDDrkfWOdWa5huflo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42416)
lgaP3VdYzlRBCFPcYjlnulYsoxsGm0eZGRK1FvEgYczC62E+/MHLX6/Hel86AHaA
+ahT7mochyBNm2RN3bTXpwIqAjPS9k8DGA8/8SG0vTPPdR1RBqkY4L6NcgtXCMNF
Ur1ePmo9Ejc/Ir+HPlWNkK8OPmjZTOYvjBZQLnJSuDx6W+odooSvcUW6FUbfbzWX
cdH8W92yuCi/A1PV17mYw4t1p252U9FwODk+7caSuKbIHCoXOQnbMv7zUUmWv++Z
/M5SneDZ7msZikAweXwDb4DSru6rMBLlaVhrSYYBli6sDI/GEqlh0KQQ8M625V4E
2vORb83TFiV5ZN8DRi6vp9LG6dGhpfkxcZo2+o9UJg12Sv0yERuWoqDruIStjfXb
QbiRytyqUyUtUCS4M3oL+f18FJxoLOOMOI73x8PxYNpqyjccfACAxbVWpGs046Nd
N0wddr9itMES+9usxUBbciFgvOcNlIz5Eutk+T7GIo8h2kzA4gKQ2b9yphj++wOr
/QbyZln/LxICPkHJ6aDQjWz86PoM+EyZyUGhhMieKJlPEMhYwXj19HoOsrPN/mPY
6V0KsVCjFGNizvo62Dg/pk5z+QqaN/hhkoFXxQ7NYea8rGvtBdNroJe25zuvouku
Ysxbe9kzIWUSc2iVbDXljygaS1rxVVUNUXCc7xm8iAi5JXCKgt6enz02Aq/2q9SB
X6zcZ2NLTR3wdbGR+8gOVq3ahO8rfmLhqdTlaVHMMv+cXUGdjXc/ZsYibVDG0Ivh
OUI6B+3bm/+mxijpCCAAPOE2t9SBhh6hq/GyQ/Ztc5f7RG5ywirnESnii2/sW2b9
39kLI3q6FslHknZ/UC8N2HsJzGxWm7A4VtqGdZZdfQyqVD0VISTe2Ytjpyny5qeN
aH3VQrevsHpyGefn8O2nU6RNbrvGmbh+VDBbsGMgmEEVIVKztjOrd5Zlb3YGS1JQ
ORwaY7MvOqQtHGskElZpH4SeNd8saYvDYs1o88cJZ2gFwLk5Sheat0nQifHUaX4Z
aInyvn2ePrIk4T9BGpkcSD1iclFC+7Mi652Y6X/8lbs6Uv99+jzijdHc82GQ/xA1
5zwBVWKj0AcHMtiF6K2uvdUHoVoEiKnKorMtTEUQW5Qb/cfEenBTDdXrrLCW1ioI
i0Hp9yJykH43DsQTUA9pkOidpTilZS2ac6doDbs3f1O81DpEG6yoCmbrKpwfXcVT
hViOarh5UrSYVCXQf1MvxftpBDh4O6SniG7Xm7Jkc5tpiZVIhtaNplTDI2vXNzKe
p7lAi+f7KYiBaFUHE9rMCrHlf12J0Xxtj/fHjYrBoATxgnnzU9ImZH2W1U0CMMXy
7fSU0SctZlWfaMMUYkicXs4TeAQF3VjZ6qy0fPibvHNTF3HMuRz7eJGM/mD8mSdO
/Y892jpTQ1eHql/Aaxh0cSermiHy+FVjROSCrf1hjIiIOs3sE/08G6M5NofWx+Vh
UmU7lRoqmkRmRpJdXDRoPvyjfRP0Budr8iic3LuhYQlrRp2UF7u+iww8GLAcSX1I
zBzxsQZa6487EJzBA8GwgXu7vmNITd4Er15zzklcpoURYBrOzvSOUUdOR4sALr98
PiNzLcJffPaARFioyKvame3wTwn4uesd/3nfLP1zIo1rDj84HnU+3drJCe0aaLru
C4HIqVrS8Xvw5xDR14Rvo9DvSdWiqhNbrknWONlomXBi2Fq3B4Fh3b5ALvfbfriC
1sldSkzsFOD8Y1nJCFZdontW7KhnKiTftaLgWtVxkT8n085o5tpPfxLA37v+/Unj
evjwjZ3W+1frdDI5Bugsp8fUZYb/PE3i54VPCCFeYOp/94ooXI+B9dCkoPizEtvP
pNJ2iOzwwH4nH3emxBZKax6DGVBr8Z9G22lNzM16Li2zzVLyr/lDexoBQprLn6/p
DAgTUdAa8+9M961O5DIMK+xo/VCCa9MgE3NZpt0HioexrC9aWh3g9SM7oim3+WH/
ASAOlYPmB5M+O00PelD+CrtT1SWBwF21hcheos6dQVvoL1cYYrgotiECoS9g6gYd
xJwcnsgrZJmQthiaczn7wV+QvllLB/UnHoAbQNXuWyWvk3EUtfkNe/z2bjlejif8
JEL7jJCYq0f2DkJLUMQRdjawSnUU4uUDici5p4Q0xMSsgl5ayapEDNsvw/mjQPTH
I5hviG5HiWNrwFf//jNVkHIlxHNC4jaah9CEtZflWUAABrDUimWDKw73Jfq+2z7U
LeDT+3ZXYpPAw9TqktL2onLTEtn2d+1+0OsbedTkOfbfnXUZKpIwJqyS0J5JG+gN
Sz3ufoUUQ28dibhKzcPzht2vn5SK8RhlCVfq618cQmhQv3MPS/8ifiYyX1dV9hg1
I9uPCytXO8xDsW/AjNj6u357DRlDSaXCAYCU6V9hNsluXFaG3iXiYFGGmUwQvJP+
4feqKEGtLXt1NYS9D0Up4+dYJB/UW0PgW3iYhpQi7vqHvWyi7yRqh5YxCHA0LlgA
uWYDu9XVW7f/HmVOyzUpYjSXS/h+EEQ1+IPScsDDD12+deYHqNYqX9YmJX5pLDaf
1CegUKnUTvCNtJ8lFsC2v01wgwr0ZtjpAOkYmYLay6dEcBGrgllFzkqzU3otHXCb
JE6m53pgVJgmoLUNFXtNJWrM50CPXP4tTbPKNUmDz9TRI4GGdMPbdF+IWBJURu3H
M4yheGkMZ51nioobLyD42Ad9KS2sXMmtDOJ6zcYW4oy4RhYIV9252oTNQwe5cDJP
2rHUKy8UI8HjELoUkNDhxkagGkCQKPAtrefPWSvKfCkdYIO1hUjALKjfczRlEroL
shEDKN0+1xKjG2/r1Whx7VrY+mle0Ry+twLi+mbXETsf9ipDVz1D4dDNsS7lh8OL
0I/Jnxpv2YSSGN4a9ZehKmaJbZxU78dXC0+l8zK2BlXfoHdf4QCXE3/O4cclJhoz
RYQyTKtqeYcAVCj9CqU2VVKQx7vnPOt8gj1ByTApVA7EUiMvKhVBykndDUB/jTU8
zw3UU4cW0c/UOKyhD/QuCNbmPB3Ocq5rpzMqAwLlE3iUoeLILvdDbJ377eCtDW8n
5+Qget/vIXHwKvy8psvfVAaPIUOmqf7QNKQz6+sfyVB5Pnf3C1pqU+XSp4E3k7bO
r0yrE6oArVBRmUa2JzTsP42Ftx258WDbCDZyHm15Y63ssHBoyGTE2HdFbsbzoPOn
EsxZzppKpY93jdpHU3d728uXp7KbZnzkucOgUtk/Ua6Pn67NASLwSIDTj6gJAGlU
7M0HPwYKum7+WPUt2CZrjzlHNx6tGDXJw+fxoT83ErvtR82XA8tUPHGD0z0W9Bpm
pdVbUXFEWoZU8L0Dfiy02rFvGj0JQ4RhUrqJP8xhWiPSLU+Yl5/L4voM+yhdxZTF
kBdTO0lj2sM0dmwPkc49ped1qf9AqzWi1YCxDgnM7vSHNOoHE1z9ZZfT0fu111RP
MMUmr61OLy0S6ObO6unJAdgo329Dz1Enlhskjag6KhCIl4WJ+tNK89hKKnaMMR9d
RGmm/8T/xc6gDXqY7jwYriZ8CVqr4dHStxqXust7FjDRiIAH+tTQkWjZWqMztvL/
1Zr3Jg0Lx0yGCky5OM1CuYh6f5bdrVMX1NTnPki0sPS1Ej05/twf8Z9R2wqyG/X7
3XxXjSCp9DWAafBTYIcubRJxxgcR9XDTYCnWwVDSJ3HzhkxWSGWMNzaasXPI0UUU
0kWTtbl6y/mr/Ur/j1QSWdHyh9e9aJ0DrT+XpJ4f50zYD7QKakEa6ugQGt56AY/+
azTK+bBX5evTPan9GgEXchPEDOoEOT3zQNzg06WrINhh3BRgpEZlVJzDVMDg3P4T
1AFD5bvK32oq8QJsdjbVc37aDbQp1eK0dBE9MS2OwTQVyaHy2awqB5S8HkTV1/+y
m2GBLMdwn+ds8VJ10APyfwqv8Z8pxV+aZDrqO9ClzIsi9t91v7DAMR9MMRO7QzkM
PnNP4RgCAaLRfZE57DOUoe7cigUwHy5xzUbL5mLAnZHYdkum6KQpWQwgPx6MYUqD
qi9kKwAsqi1l0vY5mxYsU17tADitjcO17aO61N0hOEflznbcpvkZygeLRvLl2agX
7t0B/n2KuLj0cl8GaaWAVmU9SClKLP1Q5xAEx8tVVv3Z0Uu/J4tpiKD5qezP+azK
JLxrsAFo3zcwhMGVT+Dep6OUAaM3p2YLdiI4gC/BgM++Yd92qKg20hH4VcdhN8d2
+pBnI3AX+YCDF79LQkFoVLOaqLUvY6HCBoGu0wuf2HP0ozCBEH8XoGAUJ2XJkOjM
hfhkIdnE08vQkIgfIqTChWmxzpjz0Be5wrX8HFWWlsr4BsdzPzQQWFdnuE5OZVgR
YzwfnJyKSMubJ9Sfz2C2960sTRgpv98FRQLL9Uw5W1MD5b3QvSLTDYRRW2WWucM3
dRmSSs5J2cr//PXG6k5q6QZ+0LpynU3TToSWcxpU1vvDGRJVowKc9F4eP24u7/IU
/kXbvmXfXPBkjRxBM/dHoLefuU8GffZS+rx5R/lYJw42Eu2ZOJjjp5oCBDV3WykW
KrF6nULHFZIKtoZKsc6jjqoxtNSSeaeDJWJ+sEe3GfQNqJW03Wmg19kWGs+cVM/D
7X1kAC8OG75NHkoAxAxPTz+eydIBhopBWWzkBgz5DEN7lETOYV2lUxOiczabYw8A
ZmJdVvClwxdIjdltmnvJgdXF+kOPd7tBTpoTk4P9ab5sTL6BDEFu3oFwED2lRb7I
ppgrU/+w67c0sf4aKQ7GhHq5AVyxAMDtCYbSUVKr/PVaySfnljg57bltOLILntRV
qm5m0oG4BADnOZu78miu/VjEnb15aXM/1itknNbj1GStXv6UahgApeB5TGY5Neai
CXNkuH+IlaGA3Pgvm9lZuP8lS+/0g+t//cv/F49FctcMcnY7tc4TUveYbSVadXwe
GmoyRSgTq+ajRf/elRPTlBz7G2zGyWbUBz0pXQJ7reO9jjHbcChDkMte/yLRyFjk
EfMV3o8l+9b/m6XNwY84XdLUM2kytgx9mX8zld4CH1i4b7mTSMeuEON7pm3PQazG
yISM7ch/K0XlEaIfEBxrxTYE6mjrxx0f3F6p22gTEhw5TmcDhTPN5ircqGgSkPCT
0n0OrChSbW+7rFcpC2zU515Vm1X/a0pvstWrtEfYdajeKoW82+tHFKT4tm9tgmVJ
nyav61FCwFfNdHR2OEaBLBumOGcjr9Yu5Ct0WD+J1/i1bmfINKE0iNXgxmYzGBGs
FS5/ib9gyL3ya7NYSnlbo7BVQVgqPzT0rtuNR2ij0JDHVbC0qsaYRqdWDFW4op93
trxVv79RKITSjvhP9VXiSZONU+aLYiY6m/Jo3YlcbjCBbDGxaTSjTmlX8WHlV1hV
yiqXIZlRdeh03cN9o+ji7KiMfsPZMS4Y+aXYdZMvuZDSE1RzJbSjlYUhp9p1cThi
5F5jY81PDB3uzZvdd3Hao95er6b7bg5kWkMf5aTzfwcIPM5JmkVpR015i/bzb5H0
r47tLGFZFRWaDGBldNAHea7+s36GImHP0VThE3fbYHSAdj3zqY7MiQV7rj87VxPH
ZLRKuWN40oFW53OdO55UCQ0Itdki9dKbFx/oEXThpG41Eq2k2awmhaBar7YKsBfP
XtgqteeS6t4on+Y6RODu9NloK6lO9WP67cCwUqebV89/XnJf4yjR3EvmZEHCWwpS
HCUU56sNWzsQ18nSoo61IUSTXihCAslFdK8MWwhARNhBVVJx2XLkDQGagOfsoO0C
lByHmtZV1lWPtprrjmE3Urd1Xh1K7zY6QEEoO2WZZc22wCLbHzRWou76XkHUwguM
ayEhqRR54wjnP9DkuT4qjGaJWAIzxythL5mZ7eAYj8bV+n8Znpp2ocKgMqfetTzq
G07uve/oS5kwZXCAehuJtkK4jUpgRoMW6+KArCKcr46q8z3PWF8FOQgdePBbw7zt
2s8F3v31yBUirGnSnIBVR3o7uMAj64hsK+hlKYCNlwi7SAKU1vZeaY2ohTMk/+xZ
KtkWxzRpTp3pR73Y5P2TaEJbViKjnvWiKMpIuo0fUUa7WOfGFW4390jJ9WllzoAA
Cn3vwEuGNxvXlqKK/xpROP6PP/QYA7U1XSkKt3AYqu9IyKFZ23fMPOBGPeUBsExJ
btN72K1CZOM8+wwcsNRfgFwnySOPxl1AGHUHkXGZHIxF2pDih8MamqDEnk3F3Kdq
dTs9PBi+LxxehM30sdzzTYdT353Kn6vrJkVvA39Q+/wguJWz8DEjCT3BE24Ganuh
ULpilM3AwAk8eunOVGbtdAdvqk+CM5rd0M4a5nNY+DZsPfEyJKGPVgGLSJK45Y8k
Gb/p7mhhU7vTwWld8OtH3onx+7LLtqCVxZkketmmrIU/ft/gmcnlh+Anh/cPfHbc
7VXiYUQz84+KiAjDJu6/h86lV9a9vQGqLIizdRyhkvAhnyhnVebAkW7qZZK4pO/T
2uh7SEiC1b9mUB6B4/93ikzMrbCOo5iqVplqp2291bU6A0bJ9tVzsSGWs8TF1bRE
Sat3cE0gJZ1JLKJ4jGPAAqB7zmeSSL3GsI/43nRFVSQAMVkvYXF/hcSQogT5uRyx
Z5ecsqv+/spRwmiBiOAYh9D8ceNoJwogRDjgviXGiL/uWqvJQwUXL8HmR1w6YGSQ
CSnG8pe0gLf9NawdyOAb59qMKrlMKFHeVg5QGQ810nnXbvJ8aLoFuIAwBOFk3bjg
MGj8QYADSpaXXF8ykXofseFmj1+Drw8U2EytxuNqy3WBqayYIAXvaW0ylZFhHsXX
RiT9ytvoNX7v78r1lLbFOtddSx3D/YeEL7+uGuu/G6OjESm60LPx3B3WTgpcokY3
qbQxjnCfUclHPtES7jeg+kG+yki5hI0SgdxnMVaLhgYmRjur6B2/7zwquhzVHXZ/
PcvmEHcgXpCKS/AM9IdL9Vpw7mR38rirYpMeDMTMaNmnJfXZV0/MXhGxPt1xl+2+
C8YWG/lgDK+V/ZQf/55yNOv1vOEr71Y5Fl7paOhD+12lbpnFQvKGSyh4NU2XVlgq
LpVdpmufyvc8Mnw7Qbb2ok840sG/ObCMr8fatkVxwwb31k8i4um9PSV1M+VNiVgq
yGkNku0/wjT+t9mZ8O5Z91oJtILolH/q3/aeOb+7BQ8ZEYvl95Bl9hNLmf5Hb2j2
ORG4QbdVAFweGu3v36yCBAyfjzvE8dTzXVfv48kkc6m+RqowEW7v0k0DXpwosuvN
+B0595BSi8sTyvP3kqmmFXJ0ry+1QDM7Nt92RtoJqFTFlmgm/Qk5VkQ9H+yvdzRF
g5tB1OVCcF5TP6EyTy997cGSJnvOQyqJKx250vdrr+1PHOehyfJezJnZvqrtUS3y
lEwDBPgjAxJ+P0pgYuu8oaLrO4AqC+DfgEunm0ZsjNqchrHsxg/Xpp7q7dxntJvF
PnwexAd/7Iz5ZAqHszLblpKz5Z5osXPYGnPsMUB0S/1cxLVSzvgA0p3u8OhWkbWU
EBRCPTt6AbsKr1LVHYfi0giu82GLGjPvI9dR4Pk435enZKObX/0cg38AzL0e8Q38
MyUH+XfGEulFH3axwzcNelSRN7tpT/R4oM7CVLm665FguqlCAjQBPIlg6nyAlC2W
uT4KAgyg+Sa4XgoCegJvdIO0c3inRYLdFLdyz3A/rql5A+1x7LGCG2J37uzSfxhq
bQ+nKkBlj4IpAF5/yf7vcIjZslVunxyWC4VnrBSBNbjG1zzK/ADgq6H1pUv0nUU4
D/nnu3i3UWH/pwgj/RWpVKgVxlZ7p4YqFdJk93IF87fDWKra6NSXIL20rt1JYKDU
K/T2zwwpaMJ7/fCBSYn2MKq3zfzbhXawpm/5HwDUSOAZl28OARr9dTO8yXuiUm4Q
fAck1LxZcy/I3EW3QPsqFfZIGRkAaONA671ghLJ4GJkhWZf9LkX9VFb6bJ8qKS68
DB9U8T4EN8fxRit7OV8XqyXLQGZldMdWI3pnzXYb8uDYbx4ImSDlOUo/bixBF97i
MyQZWLg5WCbK3aArSLuyVKWwPlpAR8/eme8WH90QoIene+lkdqtwN+hTP0emqgd7
esRRBM9XucHv5Z5pKP6dVPnzwlHa/4s+jjaTtJSJ/WP1+HdnunheLE9WYa+pIPqR
7aRZpFEW5vm/NnAFBzw/Oe9Bal8H8kMD33NgClThMJ38lmkxdPD+ANP3TBr3Mqlw
b083LOicm/16fRN9Z2vuPqiO3X+uuhj2EYdcxAGAxzZerHQZyQ3LNgZ/yGGTrkbI
ImsGuK/HEHyZ7BnywzN2zaf1t3r8wv4igNWTij/HiqcOYL90wHgAcfhcFJt0gIgF
ot94RkTCLP0I4igmQQSHObCk2yQTnC6qvJybHyCbFCGXgJsGkDaRgzmxw1urws4k
KPveXaQtxowilUyfPRcECGleTWh1zLimmMztyE6in/lpDOaFNAUkgWjASMRC/RRT
u2Cte19llgcxxipFKTUOb8Iokl6ixAnm31Beog1qj/k5UuCdd7K4sNXGsmlCRGsH
jYq3bLYoIcBdh9zPTx1RE7Q54CmMZapyPwdphF4JRHM7S2ffeyOPp2trH1SxxTBt
jPTh/SJ0r3bn0tahetzFtf8ek9sfvDIAnyCjm+LxmoJ9qU21hClP9pziuixEJQa4
s3FrLBQMhGeibj75QzLqvjF63qE6ccKcycIVa9ILtyNi5HSJ5CYpI7gUfL5yVGcv
EixsNseSSOOCeYE2opqUPeMXVs6kn8honqVYh2XSoYMMoHFAB41+3CA2SIOdce8+
+2eocORz8f4PzLaDsZq6NQjTgmqplWvS15N3iZ6sAady2y3q1lgGAcikcsXsOiM1
QNg8mJP+6l1FutTg7TL1AWXgwLakCf5yKXJNG8jSsZWzrhbHzElG+MG4OOUsMRTM
TBbv4il4lniUe08OIWSw9ylEErq7JqwQ0jMyX4vCKWa/vSUjF1QfS0Tb21M5mxpV
fy1fqMnVlZF78sLqyewR0fGUMMCgrPGDbwBGubW3HyHX7z9uASy8LqRqguuv5Arh
3R0nc+XMhJgHtN0RS3wFdrKfIMGP6Ed/Nt9+4mdBOkA1emxevr18AdiOtsprcOtx
dbHlImtgJfX8CopV7NZOpXSZr8F6Ovthc+uE6eTVqeKe5LTeBBwB/fzmI82uNjGV
69o141HEKmoWHWP2r2z4NXSuDNRLfH6FY8zT7P/d/Ze+l86IuFzVi3eK9zbL56u2
FMoYvMt5FBGZw30dqaEuPsunZAImMWvwc4OdztH43zlcnU2b9RDU9WCgjXG37Xos
ffgqIdbW5eqzUK719AM4wEvb823FzW40/tfxfwpH8FYAdSwgi33hTPd5St5W4GqB
2FDpC9A2xMsZ2zF6g9VbxgxX5LTV1UXmoOUCO4mhqhEsaL/sCeEoR/lo4qyX6J1Q
n/NIGNOHvIO79rvm8mij5q7Zw1MeNsqHQO4/H1mI0q7qmz+/iQdFswxUabtv8EwX
6COkgk3wWglt0OnryIKCduoWCrkuzf0ThkSL/BH4AT0fklamQfCmJgCMPCMO7Ua7
xKzVOsqa0gL0YcReYfIt6iqDDSOq01npTFvia5M/SbdHFcnLKF6FbA/6WBP6x2lK
e4FKk6/mVRz0L6U8fL2Qmes1jWkHMaUZFcMgdW6/DycTXd/jHFCqJDFvgyJRsmS6
C7CBpGfeOsPbYuxbzQgfkHlcuwilxJziTBKVK3TTZSMjxCarJmBVeFdLOUFzxBTe
NQ/J862pqwNpf5A+dhblk/8+yiRpdmcs2Ks2KTbfZlcfggCoHyNR/Io9yx4SbcW7
GE3jCAxIURogs/nHwGdYP21XCncu7o/PRw5oEZtZ5AWevppjHfFkP+SmS/27v6W0
3j0sQCJkwzSRjc/VMjWRmTUYF1gBN5Tnoxio+jbBwfKHuSfI60DcxcNGjMbtWypr
peZw93WeXd1VtL2yCwBLhv+PkHyuYkIjGc0C3L2JK5cGaGVXGh0uCgcrDcvnrZuj
cGYl24PSD1rCmtqwpI1Gvcc2y6VysMuwULlATwQ3zRZsz1XDkaeZnJi9Jt/03amU
tpcnVu9ROQa49BtFsdrPjdonkq3L79HJy+HUig6BOWDh9ce7FELpsc1QBssSITyM
xkDFsy8z6QS0a3rnTH7/dfOglgBf2c08EmRKCXguPLQb42XWDOWkqqlCbVSznr2l
Wx/Spo9xGjphsLNnsyEK4aFxl08boxsR/YrKvQ5VoFBOTX8gTc81JaKn4VOwjSst
W8g+MTRDHO135pActq5X0Ynwp2AfgFS8D8m72KUZWVu4JXtK1kdxjpjISp/s8qPQ
oLjZ9SAIg6pxJoEuxSWA3vn8VvkdaRwNYLswsIBmvf8dwDaKZlPcNGtk8llFxJ6+
SWiphrPDhVLsJYR0Y42SltIIJlzKAIEdyMvoLq37ENgiuMyaGQUqHwqr7SgRPNc2
aAZDk69la6IbS/k9OwHAvGDVBalMGFRh+mIZRD08jeVAPvH6HiAOVg38JQwijjxr
eD9HjXZRT0JtjFRTFxTwnmhfdeWHaQ2nCUqUcAvSBz8uJOsUQb6MXANjC2C6Zs9I
z1pRPIAlklkx89M7qgiNM2yzOQv9r2CaxhWADnZ6v4ySwRMl8jqotYSDUMetV2Ev
Wup+IH2DKwG/RFZLWyQXBFRTnE3pb5QJo0SqciWsiLF0VnE9g3Z0C8w5pDJtTdj+
aA/eRCoNSD1c61vQPYra7vDfFJGMmiA4GuyUAXVgoDGKJHqMOe07RvlVbNEbU6GL
w915zH42jleoq55+Ct5sWbLv5X/kx980GMd5WPzzswwYq4JaFzeSMFQiO7C7WX0R
sTjISf6AECeOFdH+mPspJ5oOUuPCSwxfb+JZkqR3NV43Ox+Ln7xqBbpEgCRshfL+
aFgeoRWs3ac6gusYk/cHnli9xR+FCoZdQl3ooiNty0zWPfpkbpOsjjEQ1vAlrsr4
rSimeYNPwKVzhBc+cd6RccJjb+sEuBQV5yvsY5Jzrc7zIlk1/Hbky8avPZI3uZQE
2tEuL/n9ItJx1VfHpEkc0jLMSvBaLqWXHT5YnO1R1Ly1Z0I0IMbjW0f/2GC83Lp4
dl4cHTOHtDMpVhupA+b9173lfweu2RXokYiHNg9HiJC8kVwlA3RYizFsz+iPC9Un
awpR/6ZcYxfxcbcL47n1yJeU1F5lBm/cjdmQ+pXC6Yr1HPcM4WJYzNoymUYLCAod
h1uypVVu6dWniCPau1PAKMdmo7wYJToHtFCFgO1V2bVkmcdILhLIUht6Cy6CQPo1
Md3b/uRfS1VgFE7d14frC0kqcx3vN2S8tlvstrsjuTSLzmVtltXDuB1TC1TFFdJm
9l3nvGfYE06ONwpyRGHna+S6ZBJRKwYlauVLL0u96t21pD9gHdSfIO4UT1svw0tT
AtKVw6NoD46v6NI66oFw2IImejuPUfB8VNVrTY2EYkGg2zUMZ2VBhRqwn8vI0fyw
oYe7NlA/tPgOI00X1UhoZ46F2AWclRWICJLfqqGAEa98PSUH+EQbYf16atYcyqs9
O/qgY924AQBNXDnfg6fnymgDhmLAAGZBmFyCbCtGGNtzTRjP8x65TWppZpm2mX0m
9EwBmM2JDlt/4xhYX4zRAXVrElHaLMFjOFdq7Otb663VVLXUckT4Y8t+2j5htrtY
24r1IgrqxkyL1yLgM1U2SiMsiEU7ZmkOizzaqgLPgF5gP9odU41DvpcN8QMCdlwB
UgzpBHoAGgqtx9qsXD2Y796Q7O1pNCngwg82wAjhHRTJdSIpKyo99Vvmf1SGrrGk
ZsAtswjN/0pEx2gtPKzwdvTd5jXbOijiM81xkRQ2XC5i3ifzV/iwZznGLYHLf3qs
rRiOIpSOkb5rhLcs1dgpKU/QILsp19ox7IjpBnJCr6en70z3AD80Lg+1+uZQyoXT
UC/rEtAOwjiZXPgl7htqsb4QDwEV/tHLCzLxMfzaYdrNppttKBtlswj6mqqHhJxK
j8rRG8CBMcIDwFBDauv0MIHX0PZa2im/ykH1dr1APS4kvqT8kCGaC7D00PShFP/g
2nd59E0MPDEFj3CSyvJxXvMwEE5w4SWjhFjmvrttzTF77diCpiaGNPJ0o+/S/mKE
XnuWzoF3puzGCOtgTL11lA7Y/1JFkoN1ZH0/adjd/GcKAx1lDRgwEcWucNlpBSt8
HjSq3KdxsZ3LjqSq1nNrFObK0fBMr/md/H54SAOh5JxLwv8dp4f5ZtvanRVeyqJT
+sg0nE8u7NUSY0B/KJ2jOdp6VIL+WXTZLOuJ+j98CTSbf1XU+RT+znJhW2oCBiXI
BqM+1t5rZx4prBvt1i8ivEbPNxicJrR8+PXcvep4sAx1chlYE4oAAuIIs707kyWM
hdvYc2iQcRmphN6P5ghNpv+8vYJYWZMQcF3/bimj8ICdVoEBnvX4LlpTAQKb5GzZ
XMzjKfaZwltJy9lz0zt5ftGY2HGiDtDxAfsOhGkKhi4KxVfkGVpSVyzg/kZurzTz
9qpKfwvslOXWvfwQoWGTnL0OA0GShNXP1r0QjZufL9Pp/8A4DhaWrdcfTJqvUH0w
WKGc1dMFHoZaMeCPQzqK+IAcHg4dkIv/jrPHCkFyHzMA4nSMdFUjr0q2t+UsoHj/
9gUEE5lsltCsZMpVd8ZepzAeRckehI6elvX5Ogv4dIwRjibnW8Wz0FjkftB4Z6jW
H3fFlK2u5oH9f5c0yezU7OJuKSjstXalg5xB7fByL5wh4ny3wSgh4Wxb5Ft0mnXn
q9qWZiaGgdPTmwFKk9U/S9bYGoO9lde5aV1CH3cf2ZBVBAE7BvbdrX82tD9dsr88
ch3bfT02nAkB6g3vvcqE/EPFG0aHVvOFLstkkbvr9VblwGxkmz+p3ec+stjYgt/t
nRyj/s5YfTvb30aOKmMqsl6jS4cLz42XGfCRO+UNQrRSLJFhjyP6H7zubrpIzF6G
Pvh95+R9NpB9wLGaafiS68AOH+0A+NOeS6Rl9k6TKlR1C7cOBvd7uzZVWLO62K5Q
RX3sbfjQt3ZkwHd6OmVMWUxk2WUnXf3KWwp3UlGPTLhmodqbs0mve0Sog0LFc5s+
3qIOtwlifP2MQCBqdVdA7ZyzY3OvvzynktdPW7sjKduHBUV1POxkWy2saUQpcH3X
b3X52Aokm0yxjcQrcRXy942QlMrbO9HKptdoYkLwB4LWsNlhTL63PMy5DsrOCSWM
Dcnp3Ek7tzF2/NR3m19Pep8MGKoRClFPG+wBT4olqxJhdy7B1n415IIUVgkhaYiX
VjWxxkIuJ7qpqIJMj6VKpVrPnjaamHQEcTOSBmdPXD2VRdeLKWxBubI4o0XyrYfB
5L/bNPnahUQvB4jM5mFXnuCLq2pJ4VT6gVP/UUWxlkpOr8OUmphCbGSFJi9VVjgY
L9YyGtdTGqvlpgslGDANA6h+t8eH0FBMHPxmbLU7vz3rBEjFsEV5Pek0dqrXuCPC
9Nq+S/YeL7d4CkUHwxPfFSXU9t0rzKiPT+V/sE4f1icUsfGPiawUO0lNkmhBvaHI
Ur1tMwe/CA4lariAIyrhcZP3SZnk769NteQNDN+phkbdoaO1r0d2jvqR31Ty4Qyw
DOtKnZr9YF4pQZBl9s955XDHH33M5F8+456plLym6xdhE8t4ZTCgNn6VTLQcLtrJ
whSUV2LJ435TmjjDE2z/8ijXFs5DBvOA8SdXZ4CYmdVcs4PGqgMWfEvdxiFMEQA1
wdS8VXeKyvo1hiJBfyrDDTe8KurMzKw2EdmMo+KiBkEWib+kQjhYYCLvrrmqs803
98cwnZnZzzkKwh1GMocPzvnvkRz8NMPi76/DioODwhRiVSDXoy+LECxRsF+Q7yvK
1KTtGIrHrfNmMocCeAiV5KVReDVHlDx6dpvxBG+yWTtOQmf3PD4rhb4CSJM7SwpU
kFrpGFBD9a4XF2YMQPCSZ5dpRe3CAg362coLpT6w2NCPLZNi30Oyff6aF2c3mHBo
xe0esj0piZxc6dDJ4BeDKMFHb16H9dAJU90sfzwUlmjmGfaXqtTOttw80gAEDK/U
fLKK4JTaPWHQhOOtPbI52fIdkCuSLxPHU5BMNvcSAEHY0S4rK2mR3PygxBPPY1HJ
ffD2qGBAI+dZSLzC2qStY7VqG5qiYAQ5b1msifMwsiAaK6LaXSaPZGfpGFjHxhP7
1fPMHS4G5FFZ9kBPFaBWcVBxXHh+M4qSUZUCgZ+o134xj+FqidTzT7fwVnUOjdav
lNCo63QOk9Kc6OK9X2oAYn+56SEwNC0h2dBL4JbvmkKq5rGhKx/7QebGkw0rmSzn
rjY45E4tPa6LSqSH51u3QM4kEXrhS9pyM3byF2qRo/X5SV/2DVBY62HWj9tgoF+C
hb3oHWLeiOGW8KHHQvvSHR+dfg/zm6fTgKlHt7lU8HPFq0fQlTtHJHMQzkeCrfG2
8JsXiDfkAjlkS/vlFzb5ZND8fo9VQJxmAvT36TU2chfOAhMm2dMmV9P7fXILkvHR
J6ntwY1yd5aDEclkgT6cHKSPdCyyw1/VH/zpt2pgkzH9WgYt7D3qsgA3bYArAkkI
iR+QKCjz6o4aeKR5j/N7laOBE1JUnZt8sZPvzXvykxnVUDC8qSObl6dWprsQH1h2
i2861nfhCX5fygnUT2lyPAJ6wZB+zSh9mbb3SpV5WWJRyRhkK9vAwO+oIMOWRFGk
hStWJIiJdWLt/wa9+m0Ks/daDk1Byftz5/tIkuzUj2m/3yGBnzFrUP8JBZTAhdeq
SogppdC5zupP5VZsB0A4zgkYXCVt/Qjo/0zTbU4qSwB9IyZvp42gN5oNKHew1tye
dA1eB6tGsI+dUZmmxBZ/R2nNA776Leh0PB7qgKHg5ifLtD14yx7N/Zhj14kDyM22
nEhsaF6gM98ZgRNXOJU+vZLyVGPwmy0SvOfj1lXL4/l9uNy8ai7rkiRKlh22OeDL
lwz4T7Mue2AR8EfHOzDLgcpEFplGH+/Jfyd8phjkmopZfq8Ss5gSJBYkcxHESA4Y
5/GsZ3g0JcocRx/zsnE4Semw+eBMZAdxBepkIoTPg8SFbXkGb6hd2PfO2emyDvpj
QNCEs+ynj8n7UZdxPLLwz+87LDhm0o/TD1GY3ggGA94VVjb6YwBzkxCVMKwmA1K9
MzWNqQWpO35ujXzdvdi9kHOHQysrMfTyK3Of2ya6HsY2zCx24kF9a7gvux0cjUmV
zebNB8fqIerqyEpYUbpt+cUYL9CEWLa3mqu1GBiMMIkDhIYHdozAGQ94mPXxwkkm
Xr0G+xz/XDtLGg7SPO8+4ffU6AAfRVmwUaoKJ1n6qaInAZfMKC7fIO/yB2CVfnm3
4Kf/2ASQ5CkjHah4nlZHygarqOhQfv3SX4nr3mgDNeVmeSqlsJhdv6y+dnsUCAM8
QoL2W2sWYnXTakNfgeBUFROuNpW+t8SVDmaTJ6jkZCw/nxYi2iJEG58uqlELA2Tx
G40s3j2tzYcbIx37rQgTmC+1pY3P9X/c6+xQryRBpL0GY/4DHqz7FBv/rLBGI7nY
V2zShL+3L1IIFQXmqqddmCbc4F1Jno2x5SYO9c8fWpwRnp5G9BuJlOavJXknBqL2
xevY/1aS+Lh4cWmtZzdeiDlvPw2Eyxaxw1K1oU+9YAv7V2/saBb8MrbJDInzK8KR
Qgi3RGjHZePVRhZDpeseT/mzUVOSZ8DoThgknoGb9E/oChyceBL8UWtHYpLZlO1G
e2AjtOJOMtQ6xS49Y1mm7HvYgepGhGRy7/ZKViM8LDu3XPTfzqgH33cn6GENunLR
0v3cKBvbt9E+KrGyhXnImyHK6WHRo0CnsFa/gOtrbZhEK7hbZAgcYlpSgMa3VIj/
+KTG1dx81qPGminfs9UUrVDmMYKPSOkjoKiDriUzMQcJ9AbmBaDALPKJqrxNpGWm
uZuXKV8iItR6sDGpHdu7JIB9FQv2YoJDzE2tf5zOgV76uG82qbOGmZMG6WV8FJZX
sHNYrTzm1VQGM0rpd68YdSw1wamiF/yRQVY7RD8aJQ2BscIzserfInHjvF9AhZOW
NflFgkS5hl0w0Di3UeDMX3vgCnPuOFhci3kkrRW9wwbBw6MyCBja2W8m24VJF85V
MK+Mb1arNEAhBF97D7yxDVhKi/XoOEDOqhG6PWDshGOyYcNXi2sfK15uOQVmjEqV
ky027GvrWRSqVWnSKBezFpNYS2HIvOaxVX0BQivlNbjg0r+/W1kk852C2AB11Lbs
HshQm5SYW5dVhLsknJlCe+zJe+eRtHrpZpLvNqyn5D+0Qma6pjqrMsRlSIgDetsW
tfAX0IQ3A2lJwypIJUtWMTyGGQssFNyeZUVYZFACI6mK8F6/mY+8YAnMQN2tMCBa
hnaVdIIqrYQJxCTI48JyI7qrkK0B4Z3MIufnXfO/xB7J/e/y5q+qoiHXIprrZsIa
wvi4SS8qi32KEgLKiJeWZf4ff9DWduAayw4e9JjlyJY0kbGBIFWbt0hHdVc6CCLu
U/c0xZWthbClviCtHJBo713wlQR6eT74zgZFkrO9LC6WOCneNkYNHi5cimNZETXE
VZbQQSdkfGk3ChGksMw6BoMxc+ORdE1oIo8x3K1Ku1neOctGikGbpgib6j9qymbP
u2ZKBmE3lrrpgFBVn+9wiCNLlX1cNXnnj2mHnY9itJlZNq8tdFGqdhwO+qLlFmrB
HI0WVXrsibFYSgf9EWCaHNypLJJnvanIekarQBxqTauMcHkgsLqKZAFqIEZUQoPU
+o4X/1ygt1yMV17Ubizf2nH52x6uQe4kFPhDB7Ivme+KXzGGkt6hkAyUVMlpKpfU
IH2iSL+tbF+x/y/kJzqYUlssVyiNE7mkeDw2f1Jw1G7I8LjkDmxaLy8FcJJJR4Da
WeDaWyIOmcXqH4x22chH91zyCs4Vnz2lZvp/PaIWSN6eNUw1r9RMbl1Pw9pTO9Ie
gJNPCJXyt3Uy84kPXI2q7izbwdfcL737vUJe6gjOSnZCpvrw0OaJODgcWPyHT3q6
bP6UwBt47aGDoi/wm58i9m8frMa1IMzx2Bm3wAJa+/B/t3HJbVr8v8Q9AQqYU7Ov
yfcJ9wz1MrbIX3uqZz104XK5sQ0csxlvjOn7YQawT7Wl3RnRiJIU0TqpxKkRJLdg
iqS7qfItjXtzwF2BwzNShsc4+/bpJniGBfh6Bdynji3uGbfOHKv1MwxzMzDlVcln
luSdO44hpOPIvxy6E8Qgalg2KtAtzgj+aD2+wV8QbyVAfQ80lgJd9SiIwrzyMqJb
4QZ8up/XvBO4JecHwFzv9usvxoG52uz5k24bINi7NAq8fksMx0RdmPv+TGgpdOok
BLDjFGcrxyHirDgvMB8Bkt4VfNfy8OoOGL4Yf2g96bBF4KRAtVLENzq4tMBg7R6/
KFmvW+E39dJafImNpx32dTUidWeHc3Nk3XzNT7gwZfgtCQtLcg5eUrJjX8BVV4TL
qriV1nyzhP1dqaCJNAW3N9HkwJ1qiuc7+hfv58bm6ys1ICvhriM65p7lZV03n4ZD
4gmQlQnG7ko9lUjgXnA59MQJDfLv/wKjZ9V0xs8gfl9TU5Qaav0n0AMRk4U+v3lX
k6jqpbQPZNsmICKywPWjY4peJNljGmjhqDOG6ErQJYCmtu+G4hbmZuqF09t80T1t
kMMYWxzv1lzW617+og+oE3VVeFPYm/4yepCRSiQwKUV04B8a2Qf2g3gP7060YzqG
b3Rmdot3QtseeNHHYF6MUvJALLUDqfBGTi8/mEOIC40hf4bsTK9US4BFfyEmB86x
IppfD02hgfSplELKKk0RCVNMqt55LlANuCxzxHURcxPh7tA8u5mjUjiMjc6Xwvo8
pkjDBSoauAnsU47TY4hqiXzi8eXO/CsA4AkJageJSnUgsliZwo2W4KOys1AYlHez
iIj5YOCDk00k5fsQg8EBXjAP1ioSFo5tPi9GCMJarwJdj4rs6z3k1QR1PxkFlQtS
qPxknzWEi3wnCC5eIeeIPZ2xdhTQuG5KfhXFoZ4UREdZDOMoYLnRPDWgymlg5O3T
6sWJd3yuzsToRWETjHhPK752cueKaPdmfhyWEJEqvxFQ337TKcjv/xlvWBKLKumt
PwTJp/gDKYY8OB4oyTsa1JR/Mg5A82FQn8tDR/TBAPxq9G1bTmGhPu82nEv1heVO
6xUX8DCH7T88y+e6wAa0xADx1r005VfV2su7aCyQoXdljUMmywzwU8CBRkydLcDo
8Tnr4cv2OeQqUBr+d4Ls8pceQcp08To/0uQhVyuj/uInkOEWdoJacCvcw9xCcKL7
866r8NV38G1CRyG6jCwkrbBQBbBZH7W8jN9jE1WCRFdKcW02IDk+TlxSkfTPbr6+
Ny9UDnB/+GELhhY8IygQU5Pp2glbz/vwEiaI6PLPK6AQhWTxJ8R+pygqbAjcXvVC
hwtnXOy8QxsVHVUU8fKAwLHfP/+jNK3Tw5sMwCXUrdSdMQcvUsBHG3IjpNhbhcjG
YL/6820JhY3m0DEnkNthmw9pGFdnqgm/qY4lhLRLETlbRK/d8AfQR9E/l5Ab0xmx
/4fEBWt1LMX0gweTmu4tjQXoh2os1hURzvrVVMkZNwvz9wQPfCGfKkwclP/sVy5q
PwJiixYFCxLjz/OCQK4Cpg4PSG5mtL7xL+/Cjp0GldceG1uSKr2S7/qXeuVGnovS
YPQrz+9LzaMvcFEoZ8rorhMocFepLKomHqZ1D9GDfRGS6KtFHFZARpTZAcMbxAP+
8G64xpds6q4sZH9UG341RApkwKVPN2LvZmMyVs/3A51yvMxiyLwLzUVEa1f8OaTw
p6JUUVjgfSRA+o9p0HTEjrYdwzx99fvqzHg5MlwqZbsgKY9slxDblbsYF/LwBiGV
RRBwLJEPG+bPm5VLB4V0JtSorcYDLy1KRPYC4CETz3t+QFNUwQ3/tR0KN9G1DGgn
O6NI0gIBAefPb3ygw9bhdieQLzK8AyzFEmW5EKgVKZSrJMUnE0F2uEVkU+/bii9B
681l39UEvukbIP9oJa6GVWzmqGuWXj8p3mDyDDy4qpgn/eNBOKMIYZHGugtmI+Ba
SY9/t3dJk9OEgEfNLmcVTQpBWLKyUBdINP1erqb/GtC1VctiFWhmP0ClLcrXhRC4
CYEHhr74/fBmnN7UmyicqXtl9dMCD3L6pE/TOkyZjPfC1ZZh07m1HT/YEMBKXhiw
lLHtoPI8S8mVzmRBtI+yeOTQIyE5BVDYSJxZJKSTexa8ndbgvYwDkaCko+MY0LKc
3CfHafPfb+2DmniIRsKXQRUAAkByC1tZX0Utxa1/4M0HYK9TdY3ytFtB+TvjgndS
yf+HINKgh61Ut2G0UfJHyNa/nhohtxC9cxTRaBbIs2zg1HFvsE5Za0OO+AGfBVpB
VEZZYFoIK0bby9sWHkEMf41hO+2LrdIF3PjR0QoNVB6tSb8rUoSDZbIOWRcJVcCv
qAPZh4oyeGO5zaAVpqGuWpKG+mObPeH/vfuVT+1P2VIUejRdOrHbVuLXX820qTTO
4A1z2wavushr6zQuJSZS5cPOPlJbvqYLRWG4XVITNfeXEnL3xI6gHtiAhLilSzMn
XD1uw5lPhjsN51FKbLMdxIIEHV/uMNy6hiFZM3dgkG0Qw6OxxLZAWdokxFgDGBQo
kTETEUpJv5r/huxRTonqXWmGJXpqs/fNRmvhEjIusJ4H4QF44IUIAYGsEFKlMPDl
cygfxol6fSsFWertHas866GfkFohwDuk/SbwZJ1xCX4aPAZshlit39Qp1YGIreaR
r59Vf5l2zKmX9Ig7KjwonuK5ZEmRWdtgzDuHSf/isLfTFlcklqDwmDCUjP5jJT+j
VNfjEk3VYKnMtAdfNH9Pi6aJD3EyI7IK76h63cB0WRgmSNHyHwyiRc2sderxwbXf
OzwBh692OBMx4BA5LEodkGmIRO1kx4rJ63HHpjs6Uem0FpkkWipaT8CZpnezbKCZ
t5/fip70kVldrSSSm9nWImyICWzCeh3Ejzfgu75VRor5SProUzeLZ4tobJxtuCIx
rmElHme5gkSeeiqDGP23E4y/UDJaszdpb1yqM4XaLXUHZiMuxSBjYMGV/juUEFRf
ynmtUV1FbqUyXf29xwoPg5TZdmA4YhdBol4wm263vaGQSsv6qgVRftCa63dSYhBu
DpAyv3sS+ovUQhX0cg1teeGreoSKnSBvqtaOze/Or3U/Q78WyN8G7Cnbq5sZWWUk
4WTF426ujxPHyhQmgbz2bikMyk77JalE70RUpHpXq85MaKNNzrM/LukSkxfsED0l
Q/oaWvQ+UR/a6y5x5PVVYhTIWhuyvCd3G3XNq97zuIeYtI50RCWScoqhk1QketWC
RlBBFt45ee4ab7d+fZhQgGUMcVfQI9+0Sp5qCOZOBxJoKcCFa5ynvEwqmSyd1lQV
VScMQwjxH/LyBmmUDcYoqV+DL8H+gnba2POAVQSFEvfalorYXgpZzLogrpjZh7pT
N+KoHBl28BRNgL+HYpE0VJ8P+kTbiEnBk9Mvy8Xq65LmhoJL3ocdpOvmtKN8hvHS
DFqE1YitK3PBDsMArZudhTa7OMnPzqqMNEba6YD4EwqTeFHhUNq27uP4Bzarz6VE
3MjUP7zDJlwzglZWrj1lRW3AVMEcc2yFtWcK0CDkFq2cnr3ClI62/BQBZzJH2IVc
8lATbu/wMfzEo3JEr3fi2ooJr3ZZu/gejVqVAn1c8ASB06cpCANGDjDEIDxe3cGk
7MhToVhgCg/Qq1xRl9Qh+NtcOWefIsqH8x4/wasBa01+K3ykRT5TER2iW6J/H9G6
4jikLV12GEccRFSUINAR+aBZI6jdTQv2/+a2SyFfAGuAj2DRv1tq2DDQWzPolplZ
UAUfSI74zrHYwWhnhxNus+V6dNkAs0JvMGl6/p3QZycdM6Vf69ROV4d1le4wKvfH
4hCe/Ck902qA0ZSHMPUGYd9dnsmTV0f8dt/jsn+xDBMNlYrneHUVGdMhMpjCMb+s
mULb0uZ73DKPsXARwVtpG2HX5gTRmWOhn/Hu08CpXXsn6hPDTGKr3aje6BKBaHv1
uHVjk8Ogc82G6x7+BrBMt5ZR2tbpcikb6eUvz+zYCouuo/1/U8OWvAl9VR+YQ0nx
4VGeTfy15zt1vr5nfWAlST2H0/xrIneRAiZQJyO1h3oPNEzettJqB85IHnmI8nfK
GjH3JwW8ElACuAXQzW9owbf1NIh/xXHJkfAS2kM2Lf1yxqNimsbyCCXJqqXx1k7V
ItxB7+aYxMb3+idHJWcAF4V22pf7XVGfuDWDuO2njSqBDsNrGRff6nWXTsGX/0LI
wG+INejvP2nPt43PVFYmwQp+ZJUBGlYQ8HyUslf20SE+ovflNorlkIJQHVl037XS
sip5sJpUAOM3lmKAKwiUHGrVvqStP4yPvpgbGuIlM5ciavvRb8ka0XspK01hkrIu
DWID7sMAn65FhiYARcF4A6+QzTbAnsPHRH0Bi3pa2/rZIzHoQgPYS+EIJiaLLB68
JPlCpxW85VL1boIAEQZ7c7HDh3Rd1eievqVR8KoVA7RWHNadQg55rKzVMPZp2le1
t8In98wXOsjWcDfgpJpirDqkX+OwAen8P9MM8CJb+EAYq40X6WZY2s3eorLzmTRU
4I1nSzHSI7aa6Tz1oKACPG4WgKwpQcbw2NTIUL/xGToOIPNQ+jIk/Ix8576CIKl5
dCgOFGXFip5kwm8h6wLHy3fO8N+E+ZqCBE/aP+rsKH3Z/p//OKlEw5ompXdCO6eH
qCk+AMl9deyLT5H2Nfllp17eg03mLx30e0pYtGV7KK/JGN3wOsQhNFRKPgxNB1aP
G8QgQwhv95osVLyKiVm2nwkT4rKlk7zZw0DvsHcGAwOCO0yb9r86ILzTxvEj4rVJ
odEwXlBUZLVLB+lE8n/Pqa9KWmS/40SCaehpSwQqTKyCsPdteaQxEqCrJyiiOcbc
KAqKusqiwUIz2HNsPjSt+iQLdiRZA8IvchFkxpXjueTUDNs0lIhnaAk5cm58EKR8
HdfCwU+VKKZNbKmgI6OccYBY/8QCPc5derQEr6lfe9vndhAC7VxFuKvN/Ed8o58W
5lhIE5IwsfCmNottYoFcd/JZ/uBPAtLOzYOhbUG7YORU8x+PG+NywYDk/Hp+6owt
vqSj2/CMgVbIDipB4o2sjD6fr32lHsfch4NFXXIbDcPQwnlLb/7gW4qtPpcaXBzd
Sz0SY1qgbmauEcPhDyDWpVS1zt8KPoQAJX0FVy8202URA780PTZGVujV8VpEguZ0
PBvkQWIhrSEftFENxZvrDxbZb5H3jpaVNGDNRG1ak7Ytjs7sxu4gn7jsAO+K8CdV
4WBJ3r02E3L/JLklK+dnMu+JNAvCCv7ahKdalWjzJVa8/mz4jvUHcXaTy6lUWps0
Nqw7TTY2SRFKRTx0cfFp6LrfRLpWs6EnZbasZAJA9Zc6LCMIpkw6Mna8HauZf5Mo
Mm/hqq99QoWb0IHmQOXs9go/sZItGtUZkCDFlsJRAIls64SS/pfAnc34ILEYlf4Y
p+pf65e4pON2VYejYcd5nWqHfS6In1c5EJSWtV4oNIdVa9ZoDMyzROq06p/x5Vza
cNqtV24luFaB/DNUDwp+BQdp7L0I1jEjkFK3f+QwELc5xpLJVkxa8XqHi2Nr2USX
/u3cXWrnapTQNrQdRSt5xztX/LrTNvJc4ivpNb4elMu8F48hmB3nATG/2uoKXc5P
7S/e9v8hvRz/15ikY8d2rgS2lv/b2PW8xXnjiZBh86u7ETwZHib9Dr+cfXCvCiLN
skYJ40hpf6v1OaxvBvcJM0Nv+brCdM2plhaw/AqcRaFT5iR2CayOsji2m7yC0BK2
f6NcbMjk6WIsJrbDvQXaAeWdIRezvJZ7yU1meTTOCbg+r5xfI1YPHXowOo3pISyV
N3gWuR74bJcWN8Y0yGGySEV/zFpKUifIrPWpjIN6zn37m3AAvJV5V7XRAdoFYE6f
BavmjHCCgFqAQtDcxQMSRGjEcnRc8MQi/w5VnESNEu0diqhjsPv0GIPJFiPY1+W9
9F+1lp4VqOoxZOioqR1k3ik4wBABbesathHCzT2gW5q26ZaatNHlIH97RqsINnCX
T1ToZkZK9kHfhxp47XwoQzb4iRW2o7RJhLwTMHzc6B+C9DbeiE6av1zuV2RG/D6X
1qLfh15NRaQ1n8IcxLL69DH0rZ099zsqpAsostFP3ZgfN3BCoNL4D3m12sX2BHIu
l/0NN51AE+GTNBe5m7Mj/tUDokNd66cJRseL0tuLwhP9EzPwftpFVqbQGxQAdwVK
Nkihza327wN/3xWuBjZ9pKAoEmbMZ+UUkl1vlvMg3HGOuCFePLRuLh1aR9Mz/Rkr
SMvJ3MGHREgzUYhDsh4xtfmLB9z2Lm61p+L9BRKlq2QYY4KquUr9WwVi+W/H2t3R
n4zUZnoozfDF2GSCcpT7tAJQhcoSH1El0EMcJQtWjlPevdnvtFCJ2KlRSDxBRiNs
z+kiO7yjgw+UeSnCXkkdJTGbJcOh6fxzUfs9BIgCitBCxkbY/3HIo3Pk3Tm1Hkbv
zrVf3tFwPLKNObTNlYicO8cvD5bB0rMRACOTQgcgY96N9mbHOprSNPEEh2zCwcKO
KLx2PrdEgeL1fLGqMqipK2aurNTIDAV2uCq1tL5qy4zvtiVsAuILeRl704VdWBte
IjB/8TcKch/Ud4QaFT1oumHpebMD4/U3sR9v7U0ZbtLbkjx3tSZQa8EFNA3Rq6eS
9ao38NNjZ1uCb1J16pQmhRHsgqE6oSie5b+qvZU0P2N4yHOpAuXBPLQZMP7ZJuWC
ahMGH3mLf3X2fWARp3+VVmk5fxtXSHaduqnysZ19Uvliz6DPGWFTdrN72EKX7ZNc
/zE4CF6aa0kJ42vp4+/039JT8HXoU28fGOjnbHtlJJGXWoPicJKJ9WC9akpPtfxv
3PJ3sDfUaidCHHL92J33UzFA21O2lEp8+7PmjMg2MQudv6AtfdAoBKkmmFUQYPC4
ccqJe7zWsinQMxlMExZV78hmey7fEuKDcGmjyqfa807idkAqEBlXxomVFnZ2WOQp
4hXZWvDCHSBALjA5tVm1uz28TQrqURYOpg8IkLImz3flj/26s2qT594t3RAuEHow
F3NapPrhuyi452OAe1vtwKC8Pxrtz4k5qaHpaXIFSSKNgZTK4H7yEnLv22Zkw/cm
deAhArx9isdTs252SwxNJv/i+/fEDDvZyO136hnugXnMEJBCy8fsfepLKYOLOS1M
5SLD1fB8ZB9T5NptDq7yY1EJmJ0zalV5USiuy7KTKXjPKOvHe8Aa55KeWVsLSNkG
D2+PFtCPhVLCgshyiXQQ8FjUUh6EDA85i4CH3gDd+pcOYeniS7hz3fFyuM6YoSW4
NsU7AuUyP6zwJLxhOD3TdlEOlfza6WLfJDkjcPtY1Ras6zrjdyyhxFKP3uc5eKLN
KM4mNbWhXS9tfSN7VFnPGxWb8hD67FHfh0YGKfIoPl1QcU62Jt5+JxFMnjX05aZb
5ub8vrAqR5TFdDAWAeiAOE8gryf/oNVF8J0RThsNfGYhMeKy6yfaPWcNJ3G/OjF7
Ss5u497JG6qOX2MFT4CYy6Lsj3tuB/8JXmr2Y7rAKLX82uV1WV94MUn3/oKIlo/e
VIs1BGIp06xWrSeeFBzgVff9+LXI+1bvjdeisnEiAhycn5BOs0FFOma11uj1tKsG
8rxpOzL1wE/3ly1p+NtDCT8xmXOdx7hOKWM93IADqVDD9IfW3ITapBp0AJmOZp2N
jfCAgYwmscqqXFgvykwmhkFC4yi5EML//1Y4nY9vFkppRMJGiYpfmP2XsT8hiOtl
Kvs+jJzOrqOtTKN+I/B/4m6G7nqFNFq6R1O+h36Uob1+RHhwlT6pQ64O5ybm2akr
ix7xSmVISqbw98GNINTFjqOvDBOl8AaTykgZ/NRzGrUuNx9QpnMT8idr8fxg6p6v
vWARGDPoRmLMpcbJkNugu/3/EPuRRuSUVpIRipdoaMKkBs7edmiGos3+uuJpYnMU
1qtbwNb/D9zjHFYfzMNmr9qzgEOnVrDOkknRKvHatZDiSNs0SdwDAPAwmoyU5Nk9
s1STd+Bje+ySYOYaOwdmFtlmKAyDfzB+pKx6yeWUKlbQJalwlvLihVb0yFk9dt8J
tVDIiyGSbQk55CSvvsBUPzlqcB+GN2lcenRcuRGMcr2lEiZPR0/3IFuBfLobq7BZ
xpRfMxwkoFFRrp6t3u5cwBC4A5Ay8O6WnRYLNFGhlMx3FC93YKi+rqdBpPLc84nt
yUZmag8LrMus2PtEtIJ9WBWgezIl2FWH23z7s/YzXeV+zpZe6CKAfBFlEj/2LTkp
CNyTqzYTeVTwBdQmEnf9NOqFeFS5l/KrtG+mutzWvW+gbsYjq0NZWdWGP0luymDi
b7PHNvToH+s7mnmX/mNQSosXbQhB0/kUqnLTEWCzNThupeN+RweAMwoLfH48oUtr
NYZnmuOOPoWwGfv7R66/H9DpWXbk/05vz2doJqVSkTRiwY8UQDyUqiwkayvCMR8V
kt8XI3O4Wd0wj2FnPyinf9nFWxrn1oYOiKPpGDVPK8v465m0Y62DYF2cCUiBwICf
HpJMWIAIfEBX1cxIWiVLXySLMl2hck43wP/ZUq7j8q0uB1rOrvG1cxEMSt9jrOrh
Qi2GGuKdesbub64C6o6jw2b156uV7nDZi/lLoWVRa2G0G4GKMZbLB1vzsUy8LOqH
/k9cxCX6B4FQSiEb1be3IIh6ZhHcR4s+1JwJhKHbk6KEWq8lWozrEBiSL5VlYYei
9yB7WAiNy5DzK3L0pq48DgBuMKEDLrDuyGP7fFdgGoRVNI8ikABFhqSuSd8IwPXk
MmKjqYfk8/xd6CjAfvbXqxyUfdhKH68Gk870FD5JoIAWqPGvNo2n69IGhfnHqUV1
aHtpq4EiaSYn4NQGtFf12OM38T7BfPd2+dEUseyMH+9Y+gryjDgSOwIUnpDewJ66
LN8Da5WhSVRa7yNmTgYzO2MeP+YuIWGN4Jxj9UMflVpPZpNgGv2a/UtcbqKl1VKQ
B9CTTESaqyERF2oAzG2BUXe5hADsXT8ChP9La/vfWUTC8LFMlHi3ctI5l2CGNxnv
9KydALEWg+0a9s5M3Ze2u9zP/oTPVK7Jd6LYDTriIPkeRRoCEWGVkPgsQjW3XNNl
nOhgT32MBlItjY4t8f9i0gZc/yU2AHVUW7J6dx0IHUkkhvawKp3MuDTS134kizMV
QBzdWoDMVMLYYHSoIOCtJzZMkkYAwQlJ+JfyQJGZ6IzfajoXe3qzzrUVYl5tDD92
Cx/84C+jzVtGA3M7KPjQZ0NLN2FJxJaSZEsUN0e7jT4GxdmLhYarW/ebJn9xSzHU
P/66V+wqvQmOYDm4B+s/k2HA4aQOe+nLRuh7eoZ8EvkQ2ZNiSnao+0VGxv15QGEM
tMMQvI3tKWOp4eLsxLkUGDJhqhHJOez2XXD9tOiD1RdqW+ayAxVERFCbDOmKgJyq
v67NvflPDYYnBjr3rIL4KHiiax8XwNyHATnuEb8LXKAHSpnK2k/B1TCkVo77hTa/
RnqP7VAhj4hkQmpXyAeXbY8iBUPfAQAgaiY9si3ZVEVXnBx1OrrIeY0lfdVdfLgk
gtHB5psbNDR3P5dyrjXxcv9/hteGPfmHG0aP6xHOVBLG9zLWjwKPnm711iYtr3+a
Rbr0cXVZcckWKIh0hWOcpHRAKRDeKai9+WFu54dj7zQlDPDBuxt6+hT5KI8HZkMv
Nt8vTP6Hde71y7sdwXMeFQltMfqozoZqbc5MBPgpM0lDpX1+LXumZLaaWqBDjYrR
Dkh3ueWVGVeh1mMkx9G/72oKkgr4fHDkfCYNl9dseWOd/4FeMaNXu0Zfdzg1qyhd
OyHGnvDoezntnUqlI8pBFOTNl3wbVcevP9fkR7rJmroMW36+Pjv2vsPHdwmYQRGC
B6HAvxoBrEKbMs3k/0BwuhXCYnpeuflfTJzwsQ+VwFgNgRafXjnKHZVTDmLxOmb2
NSmF4mKKj1WPNLZxEaqo03nSsbtJGGszy5NNvaOSlxOh1feA0fl7Qu67NJMQ/m0v
VUPfMfj4eWCAKwWtqRCtz/yYc9Lf0Wxd9nJMTt7FzEtgt2beSDP9YxeBPu09CGkT
OUkD1T3qldY/sX+4FLxnJFzFnPcnZ9SJPuiXUVpwXL5kDJx7xmzE3KuhgnD0ui0q
tn4cxY51EmYlbWQzfuweDDifwLtoj8I1vpFGUkkim+NwK5FevffWKxJpK4EgvM7K
UwYTqOgyW16/VYkux8gUZn8vYuOiPPBh2LesR/HAxEtWBpwnyagwfdb2rih8uszV
/B1CYsM7zOURSBDdOh5h44uhZeGg/0XHMXLzR2ixNiO3sGc9334bZIUYyd6xH5jf
dp/bp2+TfO1k/k1wVqyKaTAl67RcqD6ONg7rjJ6PokA3xrZNMuL+olnC4mkO38Jk
3ZxsygYC9uehP//1xBehM7264vzLkMq1vMpo6+iCl7Gk/hA//jxrYgY1qwAapQv1
6UHM6T9+i7I90kY6KQCJqY2Qg7vw/gsxmU1nliGJUeoOQOXm19IN+6D5In5LNDC2
ZKNHueSlBP/xxKcWt0i+dziSTuYM4lmmsjplm//RhtSMh/HF0Pra5QYCaB6tZO7k
DRGsFpOrltnEIMnGU5l59+yV4VGdHWAJCWFd1eegclWsab3goPs4K6Z6Ur3Y7N5T
jsilkBwjXhemp2b5mmEmaMCfS910ELhgbcv7MzB1j0hhCcQ9giot3xGN30CBXRMC
IkigAqHJHomzxM9lHiFv0df23lEmN6FtjaxqA3CzpY8Zwc7gSwzoXwCVqGrbK41c
9PqYaBWIKogrFyFpyBrj1ZlmwoKs3ze/Dh3zahC1+BL0d/vaXZTVTFB4jDsTjMPe
ZPopFFxql/xjCm6dhCDgg3Qz9J99zV6a8LO+91K+sDNVSpUAScZO2ynkLodbx6tl
gt9jDHccJNLFGxnGl1S1fA4rr1qD16YnfqpRnbKNOMR36Z6jcA4+xkMOI7F5Qgw5
KzPRxwXLP2kQU4Mw3afnidKzCSc2HWqXWAkDcwu6qHFufAQHHy8ET3QPyMxGQfxq
mr6d7sYV1p5pqAywZtKvrYYBJjYVuEVS1aPf/XpCif04biAQadFCqhu7HYPrJBKH
RYPX3h4fwRjkDy6pOoYj9L7ajyk6sJG3qthCu2ae7s01u+paNFMzJIEkg1P98cxA
NsrfQykd+pbcCIeJ+Ru9NVW9UOPSNNVIlxpqSoNVJeS8U2euBn39tqr76cdwIFaH
4N7IG8oPA7BEi3nSXwoXj8S3u1qa9RoDs4JdFld17rqaq5etNaO74JWRVO1g7/G+
2Ufw4Mrq87j/r1dMhD6Q1YcMzPDZQQc21pLTmLm3dDtPYpzot64ZLFltT+4m9zAx
Y31wi8gxvxXy45RQsLs3JGDSO8H73Km6kh7XH9fidzmTdix8ffcGo92WwaVSOttU
CLzEt1hzI1sctxiA4fOYUjI1C2eR88gM3ZzhGvCQeYlsClZgwVZ2lJ2EPv6ugU/0
QpaXaqevLO7Y2L4SqS/FQs1cpicRikLHLlHiIB5pYRf5Jqf/j2IESx2LBjZR4KhW
qYVWpQ+NNBgNnH1tFl7vCNHIxhix03a4nL9gFuVhPgrxUDpKUCMVSP40XTWUwcY3
7ZkW06QrH87GFNRn6L9vDKpaAdSVA0obabvIUzkjVx7sdnPJSB7Yg5vm3OjlQkNt
IXmxQDPO0/dNnDn1G4Aoe0IsJlkQabsR/zmChwubM3G1Ff0JcLyAxgEW7nNsbqWA
wakeuLbwdlk0BPu+CJoNuWoUWc8cgAotiMEvZvE6WMSTG5FLM4PaMF4wiXeYNCju
2CHdqzdoi/IFRggErriKm+yvQCRwGY2NwGOh2vTabea3y46N0WVk/xSyunK/Appk
jzDyFGpkOOQjuiMwvTd83hhy0eoFoH6V+86cyVMkxHyiy9u/bZs9KYM68FXL1VJN
ZpoIz+MU1dxoizeOJv1cP83n30mMT99oEQ9P115hj+28mO//LBDthb+P8JIWO7ej
PnzACor7/ZeRx4ZBpLRJYMTqQauxxb6Wz1qGIprNsv0dOKa+QmsAH1sSKTomVDIT
8pnOngBCqZ+OfvcEyKVvKhwJ0NHBTDwmU1NhKocPUo0peqTQ0/Thg3ZZM+uUDiMj
1/984OakMHQh7+geJq2AaNLmWfdnnf3yl3rUY3S85pyisPdgAWc+gCcaZpkUrDET
AqjqCE6P0vpEFsujkmxtNvLeaOy9J4CMpnLbfA+Uo5dVP+hQftOfsQQWEYaxpfd2
YUfnORk8154zZ7Uv3drM4Pk0xuKIHnTpzOT8xo/YSSHTqtfxJami/pctUNZotdBo
u6Pmk27nPP0oz+WYQooSrXcIjYcLq8kqumHY5SMtu5UoO7pV1/eit6essCg4ZiIW
FGe5hRF6QMYlNKwc7nvRCfkFwnHmpDclDVlIVuUPKJHj05uPhuQJVoRmKzo+RKGl
ufJ7iYgXrGOrfiR2nKHs/50WLWvB/D+x1XLCIlIxmtcjxHQsSV52TI2GDVm0s6ES
qszb9JdDmaFw4VH/t/GZ+RaKuxuQZo4hqRwKbyI3uuJ2xPQji+qjX3gHnq85gkjP
K1Czd+lA7oI2Q68HbHLbdOzcAjVSOO2frtzRFMnR8XsdkRLm2ehYaXJg4EpDmyN2
lUgBqtc01gvddXQcbrJaK6FGVC8NPdUxHkb7pxDQwfU10/rjPyOkmqDSIdGM0haA
R6/FJl3k+R3yuCneR5xM/VlwnR5Zitqp1/6ReYkYEH8V6E8irCOGNciKNpKJA0oC
DkOzW8wYg94qisTOVetuGwDxNpz0N+fdxTunh9iKJfxhKNhZiYxlgevJcq7XTPCs
A2ZySV1IB2wcG/mptXMYcO4rJ1epGtyXLGrejBwbur8luN5QE1oG/Buf0DS6q2SI
RY/2Ym66QRswKceFqyrqT9Upsrybc1IyNB2o5lOlIc5Hr/Zg8CaXPoLgdOkpQfsP
8C1L3v51+/EY/1VJH3X9+cTO1E6Mx3215MmG7a1KeKNySVoSbh75LxUbevdY4iWj
SwQH6U/NA46TVvoq814U/nztzjcRkLhZ8GD4GtTOoYlV1ezf32HxVEuCnaHrCDBX
l7LGh0nKehbcszoqwr6HRqLj/j2lvsU0BJ7Ba3d/+hKSFlgz3QMxBj/wHB/FlD2N
RBZ+28Czf9klyYCL+gcKCmBkuk/T6vtsWAUqMTKYQxzy/sD5p/wpljFP3g9wA1y2
GakGe8ehZm7j2QSmvHCDozqaTZVM9BP/h4UQ8NDZlC0BKnl68tGDrR6U3SrehXAY
1j9+T0eyajjQB6NRgLh6tem/z/rO2+dHqSlGlFeP+9nLoX8diHj8ArHxWb4TGda1
ijiGkqJW2dekzIZ5LeP9ZrZ5+ZYB1LXizJ4hTdYPBqk5QJAqVHo30IFyc2reKGtZ
1xxQYL3cvc7nuV/3z+L8Odbh8u2Bi07YiQymG6r9s6WNyxB3uicxz//+dZqwm8R+
1kFUAH7ZohBxJ4bKsIVHUOT9sOMpqu6+4C7p8J9q7jMTYwsYNQ2tQvxFNQQJUUty
k1AwfQmPs0VtwFwob1AU3qTAFuc8Iz5XjlNTxm3E6CK8c6jkpR+i2wXKrHms3Sak
oHMage7EwECs/HIa++gDbKNriZ4NEuSDFT9U908vWNpmMFhovhhaqDp8LzJyPzsQ
htSo9tbhpqVrMj+ycemk3BcHqjwv1ypkUZ3rQKWX9pKXZGHs4zN51nEcptFarbon
trMMMLKMWl907Wi4kRkhFIMvJXwgPdtSaDAUCccxPQuvci17J63zCN0ncL7zY0zZ
bzPG4ovwwy3s9NHkNHLAlkYjt495EWOU8dMnyY2F3zxzqekOACZn1qQMXvNITdS4
zKekDwjdmaC3uoSBhufvntn7YMfOUUerPTYIsJ/Ni06gocRgqoo1j2OcvrZF0XPP
bAQoIiDYrWVt3pRSB+K6UiCTH7Tn1Rwab48vyzNvriXTjddhoYZdc1J3Kd0CGFGk
jWkg+7trcXoN95wWQHkjYzrUDLBgCAmayimPSzpxTrIYzvT61Trx+bOWXTQCDPr1
O/MyiUeVBYX7iwasmst3HAnLq/2cqHr9v3Dvug+kuhq3RyqVaJx69rLv4jeo5hkD
Cp8HBgbPqYLwKQ7iSvejOL2iymo8IZNJSOwU0nH9DvHn7vXuTA8DXbVMEtJ0F0z1
ddQHC7DBh+EyfCqcGME782FM+1VJSUMLkgEFGiSpudbt1mbh2yKUappuQoEgTf7G
hK9uhISDrwbWOEzMOBalmMlFLWBc80L9bPiwdGMfFl5PV4vqphuKS6ZOgVsgEwfS
lw6EsxXKWv4TCnIwKqwSCuXMq/7G5JJ+k26rp98B25hLIMMKb2Pxt6u9VIzqM3fg
/YBeX/+ooHPAqlj+rTaPf/n/4TTba/usE8ZD4WgjbLVNF6FRwbmJ/SU4aVx33dn5
2VyelggAhBsEn/LslWjhCLXhSqTsL8pbQBUTP5q3sqDJ2n+rYwo8XpXde1WgAmfq
Nga0mQZv/Yiz1jNr2zqkMK3yhEyn2LqZE4ig0hocRWMhYEcFgPxSTXv23oyANHgi
QJPr1Aj6FxE3R+YVT8A79fQO+V6OQH6r9577rkYa/8kc85kOGkHHoECALAac93w1
7FBc87ve2L6aqvJfhqh+iihi/njdHWzzlGmZfh1tJrC8pbtz+yH1/BQUjPr+Y9pq
poGaFy/aKpclW1kK2Czw54ISix/6lfbSgJ3dYaCeG1gvIFKOYr2/IWZ6cvYM/wFw
s+uJan6Yd75aKXj/lzviW0R1JUI4tP7PtzMxtyq70UUO7r1Zjlpx66nMK0nlwTc2
DoYW6NpVpAiY8GKh6JnAx32QoTwHVIME+1dj/nUAbcxBjpIwK2p3X4zCMDHXNwao
fnxyrWCALx9d8BSEztOMFI1XMunuWjjmrK1eGgAFOIKla25cHLmuhR4Nsxd8DqKm
Y/RS546RgS344mdQ8Q+SzrgqYsszOne5ahp3QGK2+AXN+akP0K88H3n9eK4GDWUR
X8gj7IkZsCO6FULswzePAgZf/1bW+24d87HGATf1DumrjflqOL1jrOedQC77vS+2
j6m99h8TtAAwJX6NH7Du95AxJPJxXi+p+drwEEGGuNSVXOQzSZWnA5ZRGJhYvOUI
UcqsyC1QNM4Lbd3MO9UkLsT2f7K4jo6jzsX686FRdq82grvUJHo0EprYg/YfFCLo
81ztys6kRfYZCl7839MGeG8TjZx1gaMFCEIbWKfvd1dUVvTUBxEXGJC78F2FDdKu
En1JQt/lF3A+XZNPgZzg+IYFMpGFBX32c5AT3+yeJihuKlG4tCvdT8yFfF1dKGLI
Wb8p0pRQuFobWB6QdhYuQgG1PH9Jy7Dw2ZrXoBvYqYucVokINSduqacWFdglhe91
pclD8bkCu1AdoWgxZG8EZCZsNFXfbphNukOUInDLUq0gpFKOQhbVrytzA4+d8PJe
B96xK0wlPtdwKmloOYYCbbK9wx78oCCgQu1GNuteQMlXzukFw3xoLDN2LROhS7Ue
1KYOObvw8cPiDfDfxb/Em5hywDjh16W0SjcQ9/jROLF1KbEzrYCjCLLLbcgq2PlJ
nwk4YRXErT8qFfOlnQ3l38RaOkf3jHRO5m6jls9qEBghod0tro5dcupaqNgKnEgg
KKW73vCggVWxMxRAaK+N79igmsNr/FC8Tx8ThfFOgaGKXbJsEV4cdphXfEu0h4fo
FBuQiHXYFG1qc2o4jfhlq1rBeHtNYnTU/ADJuNKKAkzP+BbMdE0yuKRC/zIAu3pq
s/4e2+OmhFJ/mco+m9wPU+49Iyk1VLzM4t+RMgenieJ7SWkYhi/qdFAQAC2/zr9M
Pe4LbfXh2qdTQgEMFNv/0j0PhOIWFQeb1eLuDWsN5kfgOAu9s5gfzvxuC65fGUNH
HVESk1fF6oEz4xDCJVvEdlA+CoRyTOCoq9bRxx/VVbZ9gzX0poYzdM44M2H0PsJN
GMkCheu75Z1fpRFrLXLvD3gdc/nVAQFuP/l4ykrrhdKWGC33lwVAxNDLRhL665mI
+b60w9B69yTmLSg6o5UXTUqKpN8Or2CJRihu9wOSfmEeBPjOR/lzPbo2TU2xRd5f
VZFTn8nkqnsE94xmJywSXdlA/2CNygnfiOXSD911ONCRERng+pM+x+T7U2iz8M1K
bsVD4/HKW990oRpwKwd7FeL51jxzkZCSIw8KzaUHtz4xeVRtC0ozMXIYT94flZQ4
Dnu6JNdAEHJMRg5F9Oj5r/Tho4z9M0WMuQj+SYi4SYp1XgZrWinlyA+ub1+wADyQ
XcD1kZY/bn+1OyZhMnE7N34tH94F4UIPeJogLMhEu2FSAqmXqZEitlx2t6gJ3IC0
dwUApw7gEYJ2bpRVhw7Wdv0ypybHISwRFDgpkM4OYVnkpKxdSA6V7vLv5y97kEiC
A/LV4dH7C1vP5251aDuyjdkUPxMt8zB3DCAtDUaN6G7f52Op/Ky12sKXAc57/QfE
7pobUMndZBDSCJTjM1Lf+Jgy7FEGnuXJrXzJe2nObIOCLBnXqa0YN/wwCi6Ysx97
izJ1NQsbaTCC++hvdArna5Fe3axSSVKNzncDCCywzkipDg6788HNBqR7yzVqs1vd
7bQSZwOAWWz1zlcYkcmohWLSY5KdNv64S07LxFJjuwWcpQBiNwzkG4GjKTOY9fQ8
w9XUkMvqPrX+sEBIZNW/yisVo8hXJxr9hFI8XBCZIlhFTidpkEI5+FsMP387Qb/P
YG1N5ZfV+mOBFSU48zHZWnVRuaAldQDwz4FLuFxdVtsMUsKMLkYkaF+cXsA8P8YB
CnEqNyciW4+WLZfeiRYGw3fyX3DR3sJhB6xO0XUsezlnO88KJf/ZYgG0ygV3CiBK
kdkD82d/9+pDh6DJAifg1tGB0kKN7+5zvDemNTstwkonz6dV29d1xxTSeGeXYv3U
qzvsLwCIu696JsUCkXzDfgB1OxU3M6C8Q4AzTa7Df4bFIJigriGyS5LPGNIlhXZ6
rISk4BH1CckKFJgH7nRuzzfpjc3UZHge7d/m7q1s1JfOGoT0MUHH9g7Lm+R0Ccl9
MQWnb3qhVr3vcLhSccz7u3IaIpIB/02nI5DrWNq5AZgWq0j5fcRcEgKieA5S4ss5
AO+CQxGc9dKlvMVfE/pN4x+f0WOo+GNZLHjYfESM9VJotEtPAW+dnwAYshKD3tku
qgnaIOon8asoEOycagnHPQjLlFUFG8efspsovmkntbOQefFIXCKbzTd+JkEZlv7Y
DzopXxiKNxQki8PzYh5PQ7y90YjxbmKZ4Xivfua+SsThtZSWOYhCXRQwgcTwuhdy
N9DbRsEZ4CnONTEvtMFCoTyt+gH9eL+weVBjbZMXKobz1l32rVt7K78KTc2pi64c
mmI0VRB7NEIVd4GvZlwakYrTS3aQhzvoNlwc/+pijI/Ejl5ZTR8Gu/NJv1mcc13r
xXRcHpA/6wZQ5Jn2xCgcgI2b9TJeCtHs5Ody4YN13egllVErN0Bx3t+E8O3LiIC6
sfY0rgSndN2oaHeuz++o5/WAgLxYTty257XwgVlnIuYCAxM6AMjH8cKixCHXyTMu
j1BZPQtR9iZw72JMu5pbeeEj7s/PsK3ZE1UaGf017Sg5M93jMOy6KCEyjdASODr0
Q6sRUTY/R5tFXjZm034haYKsUIbfNp0Az3AnMW1vVM9Wq7Ge018JCLpiNTOrpc0m
Fibf6QokcDt1TmZL1m7F8fXhI7R22YKNmuQ6AVQiem9JimPaCq0eKGmG4dc/N+Ge
70Dv6jB8dmcd24Lr2alPtj3HlYFELxFJ4KfrN6yVru8QDUuioXXdGOLieceMRuxZ
VFn+7deu52tb7rj/gw4fV2Qfr25mo2LpxZuWfV6aRTjYMYlUwyeQnOd5aQeZIyBO
Qp8yPRjAouPcBILbwF2B+UMgqlMRzcKWResUO3gRXBdRu+WOqmgHJnPEHUJ6b7YL
WWVvYkS9EX8pbdvJelaqOpbA302pE96Y2XX4OkEVKGGHMq3cNKfkGrW4jlSEIHx7
IRoAgCpnTp09wMqHQbR4ay6GLj+MhNGza36WJ+W2aWPQHOHbQ0fUt9I7X8Eo+JHo
N4Aiavc4oxNhgt8YLIFuOcEetYrETH6TkSCVSfKACHnp2AwpX5KObo5Cejdlxz09
2hPx1Eh8/Ym6qyNIrKXUHQcELCW7T5ZkMeAeHQ89fPAwGf9zob+5swCQmtrbZAkd
k+3NBjccn1l296wm2ZwoyqBzsgxlYhq2+Opz5XdkQtXmlDZ3HNaJpFtWQnb1z+kW
TnXekj8cbuzNs+iRTgNq3Ux5uqL+PK9MRQXgHNshllymHtBQ5oYdbbFltynwj0Tk
1pK59vQKdzmdT1XHXDVE3KrFhPB76fbg9qBSTl3xPCGhe+FrJtHE4O+SnzhTLDUB
6H3qlgLG5AoA819fQD6P5WU/Z2J9e9NcBEjleLUIdpxIGIYgfxiPcoA/+/0bG3Kc
9uLYaHp6Gbj1Kpt4wUZJGR7SVfbSpyfqpUTydvfEFaV8THaZP7Zsthl8FxPXaoCd
Oit3zp6cYP45f3cvNil66MCO7N511+2bFYTo9MyoTQ+JxGSoafc+Q98/8rerfIfx
0nLKAytJslpobZz+Edy5i1aS0eeVh4ZD7+Hc0dLeDSOm0s2xAtme/HyiZP9zDfxK
1vO21HBO69g/vEqZydmOjPyaQTtmBVoUzCCxP0IQPZbf1Wp9ZrQviOYEYrqqsXCD
Vn6AKjNeMlWnzq3EKGFDEhByanr6x6RmiURkx2etSlU58q+I7dEu5EjB5X4P6uHF
vVsbNkWFzl37zwKoU2z2Fz3xbOV7dJqCMSCOmTKtUOdoYF6NeyfT2anhxxIrZRr1
dQVzlGyGcp5i8bSkg6kqgALBSO3vBHnQr3J4WVDYIvmVxSlBZg/D9p8GDPAAGp+d
g8YTIBRFWgnTfxW07B0zefvnX9LdCxP0PJ1NLMMjxUGOIArap8E0xOuhKwg44RYo
VX+3rTpv5odGWOqB+A5izvvna2bo8uDY8nX6M7JMp+8UFdatD3L11edkvmJbxpAI
GQ2nmR+iq/6dT09VJhJQGWDYYeW6nsiD4IvnoWRWSXP/BCgs9SSh2yPFPn2xZRz4
DFdi8OI70LsWOOwxf75V/0wObyf8Nj8RPOaT/bE1Vikg4NWsqYkY6CgEA99bH871
RQXbU7phWwjo5xzW0Yma5HXuPqTL26IcgVJCJG5PvJjxyIvHQ2yF0wI19zDsf1yY
3tQixCXi8jsp/3mQ0g+D2jV/ZtFjrNvL5U2fKGdyciDzjcP7nKlUdl0hES1xV0qU
qDUBFNXu2jTOlcaic2nKRR3ylSbd/fieyg5+8W+ntRpyGQ76q1d/4zyk1xBFuepO
+hcaHQ9qXQEZ12403Avtf7FUnKOKtzSmqEkslhzhMDlTCl8eNzP+L56cYYZYWz0Z
rAGUXdwUyGLLSiGMvPCRlMkxrNcr0gTWZuUhUwR6toPH4LGvcaLwx6a3a7ZSxK7q
8xYint3jhuoblR9M7WcYuXF/mPqZ/yYagytjySr6qAD9LhGpFR+wnackWvEB4s+K
6EG/vf2QQSm5IPLMczSD+3UGL/Mvw2IYdnRh+G7V6i6o2s7qvlFic81AxPSBIkpe
Kme6t/yevM03fhxps/DE/p08PYGmPYzByj+uhUZgDRmVkVd5cL61tGafwOHYkykn
2kfEiXdNVyfQyJ/Y6oCWRIh4Dwkm1kg/MhAeS/gdm4ZJN96yxhByP4V9jqKQrwgM
o7oXZWg693DT29rnwfc+Jzaimw6I3tR2o7HpdFlLBJfADT/6Z61nq2EEiZTFWhCh
JU/uND2K40hh8GZNuM8hA4SltjVHhGQx4Phj8BZmVGfbX7S49tFkw6CHGEdq6H/P
ZN3ynl2hUAuRLWJ2wGVa0fnM9daCZ6HnqNKBUHXsfTUdCDBhXDxcZXbBmtpe+Pxi
0ciGYn3GTCNfLepNDTCm+U6VQRv5IJHlQZ+HMdBR8AYDLdEYta5U6CQClhnbH+ao
kSus9th/A2uzbpFGAp77SPnLJxZw0pk0fog7VgVMQGtqRy22Fn8GFxYdKftQC1DC
YJ0L+5iv8EU16mFnsF7fb/uDgRBGA8yqNjSqs49l+2TSifz1wUMeeG5OQ3Xc7b+z
7+nMxSQjgAVIXgDEECp6zlicy84NNXRrpligoU5GWuxqZ5e4mP4lV0NPZNd0hjU9
jZ04BSZcU3oCkwnaM4GaWJ0j9FOPjiam+E1UnbGVEcN6pveOk9JnvXd3NqgCCNo6
u1YNm6cgrIrId1mnFflhJ2RdZ+6Xg2TzHFBEgf/ZZnr+wGPs5WdMUiInCskAUz/1
n+dbUok47TLZjQQ6RxFnQRr6pThJ7WZf2CzVz0nr1MSoOnGBLvOO3jG2zW5ePxJO
XB7MG5A2Z9Vo1NXy3KvR0mnsE9KGCVSAmCw1NkNXmJvqCnjzI/NtKylWKYOJpt54
E0W09VfbgWROWQBfI1OHptuoXpi+ZDOHZJQZnQqp2XXP0aLgYKjE/06Vu3zWD3EV
QLMhqW/AAI9zuF6m6+QKeVp6OON8wX6iJmPJe3vwaTpWQO+P4VoChx184iimHcD2
BBOsOKK0V655NrwZH/bLkNK3R8LoIRDaIQzWUWTxfKQCb8fCLT8VeWK7FXH5uhN3
Q9XbX9HsTHNDVKznYF3RpEc1Z9jCDAEDaRy7VwgQQztO5n4MaSc34coydTncMJs0
rF9QYIcfMSbQrQAEaqqqoj088g8HOK46hhXWE7QnPb8nRatUA/PzWM1BjCUqE8ee
YaMc1I+XsHsaJE9KUUS06OzYp9bAtRzOk36T2q3R8UUT62COxAy3EsZONtbsJmFF
2cHPw95d8sb1qLtnZ1ax9MvzNdIrKb2v7wBKGdJZ2gdB8rnJOKG0o/ybE9VCjOwM
2plo3lSsFue00Xu7CNQl3uqezuNVx+j3ncee42GCxO8XGYnouAMcrjzjNbUzycOq
B+bgbi28982qnwIWVy8OIszZaIDubHosTb4kIEHVEu60HXHNu2c19+notBj49J5Q
KNL11FMzCqZSjGEsUTE8PDVooHu93bkQ6RPcyFqo257dxDdxnpK72nt6x2Dovix7
2BucMNwP67NzH8hokThyELCF5n/p4P03BC5gV2ggOF1FJ2KFi7tttHA5iInXWiI/
iK/GRDmPkuYzHjZbAwdwAwFF5erpK4Ac9Y5Rgh/4gQckrmyxltLpwla/fR6tIxnZ
vFMgiGCqIubqF710FyLGzfTdHLeBym+eSEz1EU7/NpAaDgnxtp6nw0DcVYVavBQM
lzXHtnvK8Ec2zqc6jChPdjYkbGJMRcnMfvo8ga4bnZai2MOH9I4k6GTIBze8nKS7
3xWqp6AXib7UPHUz1Gjcfp5isFuiZpV8ikA5kpyIMfwWNRBxEsFCjCMqXc+m6EgC
1qSRh+TLwujBC79VKcY4f52s2nwAINxFyJ4w3Vjz5yN54gG7XTIdjyDnrVAbs+G9
MfdK+GcMTpx6Z88wXSAES8147dHbw4c28P3neDWsjFUE8WoGrvgmbeTbl5RpTak/
IIihOyMMS2iYP9dLO7d4N+hNrr9PCgtrbIUqcmp98//m8MKBLlJ/M/SnGLaCWaFR
HwxveqIF0SUnhKHe5Yg3IGGQ5kgifg5QXLy6EAXqusXSn1D1vow5lQyNWtupVokm
l38cKSdKF3lYJ9OAkihdwPvnnoFU7FR13Uu7dW23IHUyK55ACza4tHXb0JKmAIZu
Y/ZF/XctNUoChMZOYvW1Pg2O0foW1MMrW7Pa00wEMQUn41fEphLijlUMMW1CwwZS
Dlp09Y50PzA/ljPcWkNRIMnlw2n2JKSxkpb4dBMzWxoLxh2zwIMD1lLykL9hIX5D
31/ka1HI505/KPAx2oUII8W9oCj8/E8GVK1KF8Vre0EEB1c6tOtXGxsaMxGZiuU1
9k0gs3Cq494tQory7WyQlOgFseOjY7uYYXVfEtz4iagobgYmqs3cVxqLaLyc0s/t
9OMP72p+mJeDn17/JT6TFUYLPteMwy8Xt6/dEBS/F6ZoFtCR3AZHhQqP7nNj9KyO
NX28K+l2r2hXEd4O01YwNFw557foB0XXUh/WwbaPtelENs4p+lIKqQddTabWCx67
gEB/Mu6kNGeELXbLPs/QEhYTcD20/EDoQHggjhLNXJRMlWZrisON7IyhV35x6yw1
RpW76XPNr3KJMUmPeCeQyWEXznSvialslWwyQAeHpGzqQKjLKf/PufA50b2Y07bo
GRMvonh2qNzjl3758TLIZYb8Oa6l/9EWY2MBXSEborjaHduDdDpwmO52rPw+ZdHc
noMqWfTmE6KmGu2BXVqPEsqI0LVDI+b6bt2R+Jbm7aIOqQWgw7EPFsVG706VzGBu
NdoCECUi8DOUuGlsRvKyLif0h2wnU1D7zY4GvGQLUaa25RKB48OClzO5seX3kiXi
+tC3q0CRkJkPNN1Xq8j97blompfha6P5DEwMfefq4FPJpw1En98TXH0S4WKucyPW
MEB3fyyHOJ/AqOmXuhZ82quA2czzye2cnvvN3RTFRDkM5HNh0dG/nhSK+u6RGD9X
NKCschYBGV8Y5bP8EK5Rid5cSrgZNtmFpoPB6qW3krE0otkF/unipw51X1kdQTay
nFZ38Zr6aGJCdyvJ/u6HAniq7ytuMoNKNfjXWlQuOhD3KsxWGndvUwEPNRtcLME0
PQiNssZ41/yS0TeQH1noSeDFB4IduBJ+hn3HBRZ5dzO32oD9XdrKYQQVvXwWyF7K
q2fM4I73+e7mLs0VJ7RTXDm81DyKVM/UfcfW+FVDUEd2HmUF5h8GIbNg7/u8cRCz
66MqJVsyAOF4i2eGHmAclBHdjTkjMwCSHez5ALFPT6hg+3eqx0IAntN7exnKatnl
q9c6hyYE2fsGms8Shpqzqtqmf4zdcUt1W8og3hB/pU21TcqzvROANGRFRlSCtnGB
yi0jM7AQw7CqPyUwXIO85+1dXnm2HfRsmWogJXI0wUNwgVc33Xln6CqSW8fdhMR0
6cYrgW23UZxXPFSlENNU9DrAVjvtJvWdfDjXNj9ZRQGPMS5w/6AFeBy63pT2oI3g
pAHcBHvvibu/NDQcq0N2X0cMfoOU0KIE+6xhITy0gCbKqq/YegdeuL+wD+z5Nb7j
XqCnz9HL0c2bGeFDPDJcaSHK4Qz/Xanx+w7S1Wt53gj5dKEgvtDHzLmTbN9La++a
yLwNPOAVp2wCiCN8m9+0j2725mQ33p50fwnipxKW6fYo0RdKoguvYTBOEIg13d7G
XrG66DX7XjiNzdBEMQPGryaOkGxheD2KljQGhOV09oUxB6KoVh3SfZnfr1kDMduV
0YPEcqE0V6HgTAq8U+JmJFjPLxfVoOC9jJ9SXjz/54F89NbB5YROqWMRkyOJC5ml
M12x12KzJGnmYPx/whnWktKL2PaOQ+1CpzxmRhDEnSCclsy5Msgba8Na6bGAlJfK
rZX2HX0Gg66Lc9vkND0Zke7u93WKJDIcTJZPxFyf4CR9Ns8tjyYtnvn+q1DRekb5
F/nA7IhrNExL6e0FCtdBeaeVA+VD7t1FTYuqTwyg8lM9hIBSJY9NRgmxXo/yJ1+u
ekNpJekciTRMne7TEGXJja2b8C7mkhkTPxIE8gur9uu4QvzChSs8c2W9BoxJPZc4
1Q7/KnMzdOvDp2H8qOfzD+4IMOdYtUlUUBcrwfsV/pOgfJqvoqhoz6K4hCttW+sI
ytmAkAMIRp1+joWQfAp6Pg5Ti4D/C5axDfJ8e8GG9nQghCEz9l/j4SYb9mBrYulc
yfMZ/mopDUqzyBaheXIr2jXnh4IE2toeT+VsSlncHqQEYuLO58dfegUD/IZjs7iJ
73F76q2KXR6zTv8vUuAA6ZOHIRuPD3vvii4b4jnjX2mnE278E5Ul+k+7/ka4mq2+
dxgLXAnETjnDmN1w+9noWShV44+zgYo5t2n9EVHM2HCTY5PZ1561o0+Ms7qMUftQ
rCxYSC/EcHJcOHDw3HFdPunz19HicYuKty2RUQ7Hl2p3nHObQsVR9mkUDu9lho+o
QGwpuu4dfqbMOtR0RuZS0UkZPI9WIApXJ41badnWnBP4L0DdPK2oD5TmBcfCR5o8
e1YszOTSrxYEAMGSmXOa2DnHAQcx05vCD/1eVu1w0gqLum2zDxZFr+aUHQNJNbHG
hLUiDyMbo/KERSUlsKICHEBtzijoCIhXbfTpRpWDP9MN6cvV1X7dl1QqQaZnUk8u
VKxlUs5VtRfc3l4OOTiIDgoUo6EEd+3EhXCfapy59qTOIycJtTE1RH8YfsepRzdX
nDqStLYmzx5jdN12p8u8iW1TbkyR6ILfqO4cegR/OFTeATTlwu1mS/i3PWz+o5Z0
DnPNDFs6XavX2s6V9GgznlJkZhLHLljezxmcq+VVeN42fVcC4K4Jv3ibr8JtvR2d
uFGgvXd1SvynH4W62j0FsfG9cC1aQ3GVKFMQ2SLGncRmxIOO5tpsdymJzasm4/mz
pEn7IW/rNQiHK8r1H36lhTGy26moj8vNvx8LW1Rp8e1/Zx5pZB40KgoFH+WbWw21
LJLnzC2L8LBX8Lq4gEjVsg05yR9asOj2w5Cg62s+tVyECPsp/QCxmK4NXiVJFylj
srethVC+TjBV14rei0+4obxGd6AhBX6+9KWf5WbAJh8mwgPK7oGUVIk8tj1KzI8k
RMjZoIrhSLny80hk4fbWX4gd9RVho3G+aUtPk/l0lwuGpTcfxYRLg8CWPg0grZrs
BecPJANjwShDYMzrl0PAIMQZgCctVyVryVIvYE2Y5f7zHoVsFkRvUzfD0iQ4hxZv
bYqFLgAvdB72FuYM5NOBQCLao7x/GY53+Wb8MSOIkzGVx36/6PKMNqssfmHlbMmt
ppoVIdfo5kmt/W/gbnx0wnx8Km2Uaiz4hz5emDR245TRnfQYBFmV3HYaadyYvEdF
SeojPr9qndMMVqik9oCzxHG4J1YDQgX5bX/C+ySPLNevsF7S3OHr5MM3xDOxx4C6
JbNWy2AGoeZYw2HFDsdwYFkbAZ6HUk1B5H0oa80sQh9YbnXqVm6V9Zc9D3nB9u53
dyk7cuYtiGf4CnMC59hMnLTew5HZRCE1ch6+T5ssBl/r66VX0v094viWKmpPNKe1
iLO3E1+Ch/WhHi0EseWfsS7uWBI/DwvS4niGK4EWlAxLSWv693UW+O8/eO921jLs
ls2B8Pl3qbdhfRnvGH0RP+4lXeCMXtlifvEDAUrY4aMpR2s+S9k0yxIGNTd4V8a0
jOPaOEnf7qzmzyd918I0xciTwSNtTort850C2jR2PfirezvnNlS2ACs57irQgHdq
b/lNhQQfUddfCkVpuZfL7gAcAh2A4hvhz9e9e/sP27j+QWcjIU1j1tDoGkV0/1v7
eLowxOYCLDjyYMgisbjYNyKEP50npSUrP59yv8Z3nPHQfB9FsVkCRv5Ja2qasSvO
ERZDN5BBhSnRWUCXUaRIxrq1Y+OQs1Gc87ZNz4gBdLC4y2EiG7mhTGvkmb0/xuvt
iR1gO2cvBdU7BVK9x9w7QBmx3kIncC6PCSgE8UkU/QM/ZQEn06hOpIxonh98RwzN
ymhlnergzjqfYPQOaSGbfGlzXjA2cVyOyO9BlcjAf3OZWzFQngBIwPR1xxKZsfiq
hmPm3saWx5A0FtZ1v7jdZw2HNKbPomucAzaBHacn2wjjplM+tGYn0q9KVjoREhJ2
jZoMe1w3AsIk3jdQQGc2UfDf7SZ5IRXHXscCaEDgYbfANAxkElnNLoEXZZLW6I3w
ToRklE9pRwtbtxaqF0D/QYGqhcO1JaYA7AAf1nlOF8ERqYEsfh3k+JZBcnLJJEXv
tHXUIYF0soHS2eZBlAGTg0qtsUZpND0IoO5aQAyjwt9gRZ0boWTdXcoLw7AfPXC0
+2iBYd3QlmgOMFoCs6mjX35mzapYNLBwOGmpxuvssR1p6isL1g2LwV7D0mdJDDoC
EDuK9XQLUgFn027NQgkYL97L39DbwANF/yAb15iB4MFeDYGLhItJmoQ6fi1UJl+A
MCEGnoRCrh6dLWwHJp2NF49EV8W6M9E59izaLBncWdtPD32sZo+96gwL/8jEtUQU
xw3N2AHCBU+it34clq7tgP35s8fMBKm8yt2ahndwHjyaOVDVYSQaCg7myeUgvLRQ
a+61815B9GvKegOyzlB2Ev5hX8Ypc01xzoo70eueVy5N98GktrffE13vnVbOTOPy
0TZzFm42wPv70v8Tgm3Ki7dhBkyqGyMl6xbwCmE7yzYtHIuIgqFpgrR4MmHyNE0I
8Vum2WREQdXrSqcU+L0twJoPhKw84XSkErQYfMRu+EhyC5DKyor837r/967hVHOr
E9r5lKdIoXjJOThlQ4GW+6pHr5IhGgWkMpuOmFPHfjBxasIPNjjgVO33axSrbg2s
GDlivgr7X2fSjdbEZToZewiN9EE4FujrgeMe6s1Rnbp+SwyjXgxVjjFioG3m0TPQ
zukeDxDUX4TKg3mBgUzyOfIW2Bx0lAX1lKcWjMLBqqN2Q/6ugd68VK1gc5hhcF84
QcbAKBq8ZUE518Mi7yOwAPe+135o6Z2cDFa/s39Z6KOKW0SdU4W59GE3MtNAcY2Z
4EAP6z9vYifYKZqX4kYGDqAs1rTGc4itLpvL6pN1zlGS2OMKTafN+e55kTu2NC6B
SQet6SsA0fsXQIg4OT/y/pOWfqjtB5LerHny6JfV+gS30mGRa5OdDOJA7ZxkrnB2
77SMa0WOA2mKHtPDQcwvSvdDLcnol2T0uZj6g9UqIs2+7/IvObn7FD3ZWL1Ee618
VxPCUH3xne/S7nP+mHtiboNrX9yefqS//ayLW9gClMhArb6W+sCy/7LjJ/Yxor/7
oXMGU6iJQp3lNH+VYFlW1BgAwroShWcp+bnsr3yfu1AJQQZBZSdVCPKPVh0hB/dd
W0tiY9yfhytPwWlo3RKDmrO4ha8fw2fP45XGFP8e5tEX72DD7u2PSqkzI/3gXQbb
RU31yK6N8s3D+BBzO5Mmybds6CrBaW1zgoVnFChiNMBL/fCXam1yN/GHQvMDXowR
RmtPfrnyn0VL3z5IN7KR4MegTJKNhvcoEvC4cucYs9NYXxtiElLARdHkY1MnI2aZ
ysyA+mE70Ov5U//LMGiwxbMtP3R5Rx5KZhRCNIojKZiDB00ro0XWDNibVi3mECyZ
e4g4U1/p1c51BdCfJygp3wWNybt0IHG17vuM44Ohfl0pet0k2mLEyjvC5sehEfcy
16/M99L4uNxZpXMjHC95QvVk0phiHCGAwx382OgbgwOdEptHhTKbovXI96nx44sG
/0xD6Uvq5sg91TcPO2RNzX+VZSf7TctGqQ1sfT8NPAPLQ47RuOUZRZXGlAckSB92
bsYHBcly4l2050YY70Y/sSJIJXJFR6o1cRt+9FjmQgRKcr9FsXQAX96jm/fcLkQ2
YNQITSFV0Tt28mmw4dAcUAF6bOODoRfNS3Fyeb/9M8yNcunfJlKoeSCab9FffYbw
A+PSAH9hcpQDoJCTIv4PvcBzfvH2DikZyTUULHLbAK+MoXPEP2D5OIDPwdUxllso
lHjeGUr9sAAoDeSntbGdfQuKm3BFGIgNmrUWyRTaeHWjPDUDndmzkxs3B82xSLBl
Xpj077njQrQuAkkJJIx0OwemSNuoNN9wXdw87QumAAIdUGrs48+rgypdr9ecgyYN
3HW3kWyWxtoxxCKSL7o8vzM/3ntoycnRiogXuDjlPX/qlHR+rtpzlzRVIOrro3lM
qoyuoDmj3GuNlcFYQWSz9uCfIsEKq1j3jrAfICSHlXsyH7K7uWUyEQqbAo6lHUdQ
3njHAKjwses5LHYn5pUyBpg+0oL/F+8mig75SXUzOH9Y4+eABPH5L6+B7fjgESdf
5uK+hxKnE3CoVhyFbfEI01hhUZm2m/rCmFWqzWFKMowMlro6PYz3cvUVF4XMPu2R
t+n2jIbKcDhrS7xcgS9HoRjPxaXrE2t5R/+fiaYbP/n52luqECiUKjFrJw2uJJYa
7PZJc1g47f8hSbXJck8yOJW3h2Q8OEjqk3XeV0VXdDXQ74zYs1uhO5hDuBmH/hp6
7lYAGhhh7nBXgk3xCt0nQdeumEggg9i4jYVBHlNd95HVvEKGJ3EwfVBrwI8KJuUz
18XCy+12DZc/xh+9Ifi/6XXp1xWayYOzHIbJi1ny2lGFFZ4AxiXYoERO03GF9Bqp
CFMHyFTihSBhw6x1/1LIAOqZNEqiPON3uQ8rDw8P3LT1J4HZUunMYaoW948awdrk
Xl4newXbdHmZ0jlsiOSp8sFg0BS3rdhAvKl4MBBWXDesdt7YeEhKYOowZmv5gZtv
u2iceklvvZTYGxITBCI46g+tnZso2gSVhItU1+erPRSw30SotnQTBCle9tkgxl6J
mH9A8yR2Ea7Su3YyGHpMLOsvQpXTszKQ1NZQ2oraXw/K0b8aUWQO4mulkfN6G57b
6bMCDQNcwRns68PXXYMK1nb60h6mNcy2vo3qJZpPsc27SFMoLbsJtMxDgZRv5Wu1
AMPhhmYvMpM1TLR3x33duaVbnct7hkH2yjDWb/ZdxkNjb9Di16b7GYJjD+wovYsK
dB0+ubjnrLl1GwN/RWLkfy9SWW3b0YFIXcxxtnt9XN2PW2PYbboJDC2YI4q5afQ9
X/RZfYCn0w3rXqplR9mzYLATObUR2+6Jl2h2PUByfdKej8F72zBDJR0AbX3VvckI
Qcc2ms6sSoBF5RfByKBgarCxxvqy/jGmHgOCrTSiSwe6Z8sjtiCErs1vMWZH9wyb
vCa9Oj7nkIh8cGkUk/pRGXQ7HKAUtU8GYtMbgFtSyuAoDmKldBmHCiECuwAWLT0t
6MIIqpLlXUVJO4Ub3g7rRwEUZffvwSBPM0Dgu7TIXHbPoHwpmK5A+bxgzBIP9JdE
luKg4hgJGpBLDYlpa5lqNdaAINjuZiP5fzzmeady9UmmQ1joU+GgAbj/n5sXMZxU
MrhwsNiZ6hftyybSj7I9nnMtt9MYCESr1Y+5RJUXKHInFHEmFnM18QN2o0ZnFZe3
LrDmNS6Cir1cVbnNnfq1NM0y3o6DOHcaJkM1gvnpszLGW901ZXns/TM0rj7vIqDJ
6t3XKBYUe44vEW+nwOhcSPKJhfNlg69TF1zgYgKptyMU8uD/JFNX11bjhZKKH0Cb
oXOYk1WIPXDC4sNF8FPd0um4hiewEXC2vr7GsU2dexdOUb63kxLACT96m/t1D1ST
3/GRDxHc16LrIfHH227dvMvdz1wPj3mpl6KZbEDpgrr+44GRsxn2Y4R3vgv/xdGk
r+nwtaXUpgvUiXUt5QKD9LzoSpx8cQdyXhQtSol2a6F/Pc/HDTow/HptbLMFxSPH
1zOhk8+nzPDJ+2SBAo72E2JtA9SbDhZgPDQPCflwv5AKSt28xY98tTE69HcQk+Ed
oN9nfQrY+3+BcRWnZQCjEnNkxqlfnHHZM555ldm2aqvlz+8r8CZd1cOq4fjau6Sz
w5UkMqO1hmOrlLOflvWE7dcq8yNNgrbr+dQRW8VmKZP5SS46goTnyo19+vuCRme2
zE18vBqoPNz+tyVHnmsH2dgiqsI1uGGP45RvlYMeWzr+GjNeG6i/KmOLFxBQd39b
SvYs3RO2cg0qHhTHYeoW/NmhTzAqpfRbNFbEXUiJGhp7mzEDI3BbYzFTQ3mxERGj
piOptaDaWYsiMscSiX4ZRYVkegnwf0ZGG3TXOROLUu2UjQ5aEoCS18SF07y1efK9
NX2E0ndwiT7OoPIc9/kWx/wfn6wz/qABQ8Dves7QQAzmW5ZBsL2+Ovop5gsaYSvr
bQzDlJNMjEPLG5lflYm9LzOFiJZJ/tVn+eZfwRcyqjb1ujHM+qu57MVZLem2vSQG
fdJ9m782EqpEHYQICB42XrAbUP/YmrIRzTIK2fsca3v1h6oqZBKdhXdolQHGBQ1M
qVfE3bCieOWtL2irgwtlIwb0SL31oNtoNaMjue534hpm1INT/N5B0A7mX82xdd2V
BUq5CwhHeshJNw0oVKRQgt3HHxsBK1wr3IdP754sXZIcr5IcGCUBkh/jMXTWONYb
ajiyf95bmwJ0GtKipl3lkLDsUGc3ifyW/HegiCsYmyVdBW3o/mTyv72TVkooBp8Y
pApT4y7tFPwAaoyZ0kah7dYrrUeQsWox4fXmfg8QSa1iAD4wMWj9T2vGtSVH6F4Q
8w3yk8z2FV3bxymn/5B+LWOrD0lhu2xsNUMx//QQrQ8QaGn6eApFls/Vdugj0GxN
dCVTpPr1h2tuyYabrqO3P7Kmg2e6ooqUVDt2M1xxq11jRyGymdQK/sePqY7GbYkK
fvyLjIvE59FdtNpHEDAJPXSwAhj91ZIRJj/KNPN8PW6Fiok9MiuGTMNNJzDOMOEh
yfWkKMSBkpU+m0b/U92vgQtYReZk7dwtwWi6YyWP6MH7okqiV5eXvYwirl/PCmq/
soIEQ2K2V/rH+sSAM/kuhBrRaLdLo6iLD2ElSSrRM3OC1Ie0Waj9L8Igp2fV9Hpd
rHUF8wJC9HmRLiBIh1g9XQzsd5pfsvx/bjiKNIbjseJHqMGmFrQ6ATsxSCNvGlnm
uQq6BQywR8I4v05UyqYao4Jj3FAH2bww7j0Fw6mAfQgY7eckRZllGY8jgYrlWuSK
klmVSAE0JZvKmHtnTnj7vwLy5ZZTqpAeoDrmdMzc/IJM7VC3zaPhewxjMGK2euN3
D+HzPCyis24RUSmlnezOcq3ZWR2d5wXgcGl5rOwDGXWtz+wAKoI/i5InDd80DxmF
4HAyw55XbnALrIuif3IpyMA/G6LlqHblWrOkj53gvEk6esz7qG3VEPjvOyFy6+x8
dzsMnk30ZItbWi6tnkWtPoifD9+xGe1w3uBt3DpMsGkB5XRPHbGL+SMldzv3VC1R
ljq4tV8YKT7qtANyQCdAbcVbRk+8aVYOecN/Z5LBJ24l6VWtgUts5G9OYQWXzK/I
wN8E3ludRp8KMS04x7H83ZRAaevzk1hztJeRXp+1ulPW7/GiDYRbQ3DTrKEvuJ2s
wJXcZIVNIGjccETr7asJEFM0S3lZusYyhAmGtSDbowdvusVfLv61G3RssKEcQ5E/
zFO2GGbNYu4yFyMJ/71NxZ/pbIVtgNLOgOgcZBqN44eBTDZ2M3e7O/UBRoc4YA7K
lQxkgC27hzyOnVkXJpxwhE4rlCfnXybvVdq5XRwxMwjlLgpyczoc9vzKNNKCIkfJ
wkVhXR5w/ha9c2L8YKo9HvtncfBMBgcvpth1XDYZFmio5Kqbsp7qG1RaCJ3FUE+3
grGgW75n0EYDvcYomfFv7vIke1ElZqiiMilNTqd9Ar1HT8gVptN3yC25s8zU7qSS
aYbZNGOmCrgOMY030llbSh9WeXBRlh+knwSV9e3t0Ebqg8kYXnkNylqxfriHWeZD
oqd0Xv+q+SFJpg2gPMDDQ15Db9AQGDajpsgDUtg7IHtMasqDyDqTM5/8WTUJC64P
37vddit33DYFqyg1q+wbeWw+bYv/oZ2uixFKYH9g22H/0iPxPy19BNaoGR8wljGC
61FYAicnbAbzErc/e0k6r5d6Vh+qmKtdmHXRm8Jbkc9gPjOi+C5QEo0l7ngfBBLp
UOE9raIeFQCauFAwegpfZPzQdCVxHOkfrutcvykRBkAoZHElK5PRuXWEMOZyrW/p
DqcGVqfymNF648Rx0sw/GMAs7AQVCmY4PY/q8V4r4k36CMjNGyeISUpf0/cFDovl
uahz5sQAcr5gi96/LTyj59jsrF4u208LwpibYaYwrWzSppFCCFhKXtTDY4JfmD1I
A0Vnq90viegu4m73Wje/d5xxl/lftTmjJnF1wQdn4TYu7rYMHTcpfGeTsDxJcSt5
tPk4CpOukBoa4luu2mUcdfafirBo/eURQl7YMXa2urwc2+vjCVwtcqr8VMJqJRTG
rHX+in7+ggfQQ9Lv8f/ZZQewRotwjNXPiqqAC8F7EeE7V6ZFbkuHo+XJD/SBWyxk
aEYf74ODbKW5pqUiiuSek8gmkOwTn6Xyt4R6nFglbopurDWPNvAZXvrNhMfTBRPa
AspbWRtn6mNcYQcl39HOeqVuvQpTSmtUqZMQeun9qOYudXjqpHEgrRJivbVDODrA
eA0KDz7seczVhzhC+IYmLYOkFCbOajIxPGwaXPTPw0cRNAmfbC6ACNVXOCq/hprq
yDUqf+XafSELwJDXmwO4iZDOIMMDNZZr5rYYi3cTN2hy55fWdjCEpxi0JwLS5LfB
5EMAE26QoybNUgSbtQkwOF7PK1GV9owBybmL32SAsb3CSl1bF2J42KvunN/W1/ku
bz9fbHrnW/VVz576NDH5hmBjpPCCw0XU7kXEu6pPiwqKCwnAzFFn0KY1CZQytxq/
GlqOHHTokgUNGwjzs4iMvM9+TPxbcFSPxC543CRn+QRFSLO8e+9sLY8FxisTBR4w
wB1OyEQWI4YEXkWvUXA9Y3JKs9Lt2R5byvVdN1CZbGviJF6ZQbakQ26om20tyDad
3vaPDIkKTCQSp1AuRH3nNy8sNIpib+Bl1UhDl70aQxWiJVWQ2hvP0u/EpQE3reZt
PcP+LJYlWgrEmHOtrnS4nYUvduBcHTwYTKzUE8/E9tNfMHaRaN7ZK44UP1Ppj1tf
2oKDJXWDf0mhSgT7V7PfeE+ycqXWUEQcXF0dXok2XmCn5huqRP8pmbCtNBc5URzz
PEjf+mr8X9dN7Y5iMGKYIMfAMoZD915L8Wi2zv3JB+VYg9DprJhUvWNfsPDEmOK7
BCG29nuYOngimwAfUi/+jb7+nAhjPmds09cmpbucTWRMqrDLYaRDmla+uuD2AxP1
6QO+ia+sR7vVK7M8ff3hXmXYPcO1BBBqNZarM/ZFVWAOvdXwmPdg2TA85p3MYOQz
5wRoGxn1HvWFOycJiV9Zrb0zFoHVYgFxcT5cFNSvDLKv9VtnrqwzQNjK0cFhGNUq
E0NAK3e07sv27ozoIXIrYhMnQEQ0yrDWOW5xZgxMjEFNAimLpf9F9tveWM8yYyGN
9mgdLn53sGP6NZslSMKjwEsA+9/p5hUohc4vL+b2x2+u9hkMoFBSV9q3QUuFhdvD
Qr/ZzWR/u9ZeRb1bD6qH25W6NJSfogIsRJ3Y1Dwqz0+FLC6CIJP77GiZioePYh57
GwPXsLywsnLoXYzaqv2lFWC/dWQcusLMrWHeJRKNwzDMhq4c3Nx1xrGwdeicPWiE
jjlDTHmxiAzEIveDB6KX9Fk7k2TwSQVtg1dTB1EIuZUkE+3R1SxEw3PvygLuXPk8
aJ5ZF3TlWWqmMONUaeMJA5LyrWXL/dQ/bapc7GLsHRK6pliEAHCQYb9tJ4LGs5F1
VmHEtIPXeoAvOjHrGhOuv9CC4CgMqy6FwksqIK3Hvuj4J9ZHiczDwwx88kUzl1BQ
1whQloxoAavPBcqUf7rdKL+H2QY7joA7P73h6Nhs+dMont9UEyWkudp/hFW71/N8
B+q6oIHto+iVmKFVJywLOCjREaPB+KCQvaF9kL0JBUGcxuty64MW/iQG1bXv1Fzr
aeg7Whm5aVjph7DKIC7irOt+S/6wnpiR/ntRcL2IMwRQrHeLF7yZRZ68drE3TmCj
87CMY8hxMxgbOxc/Cnr+99+B5je6M4UTjUqzkKKehyEXbHv83FGKNtgxxFlyxXRm
ia2lGBBSiXTF0+x2xo9qAXDPyrLd27CQ4drGc+b/G8FvkvO5kFJjLqJDcpE6sbDi
Yu3iVVTqnJoQ5bGVzwD6SpJoTxy8oSYZmQbkGtRXMZ9VUbZLiMRLxWFwtAu78R+x
12Kv+KsFYYxgv0pMLSKgp9jqdPk327TlL6n+GiGiZjoRL3ELb80WwwEEMU1OgRgU
uy6G2MbEdiUNEV97aW0IbxEp1g5UnJX3RuETlcaLBp5ueLKrljRtdzdLg0/cSTJ0
58yqMZof2+FTpUG1tN4U6TlEB/mNbXILdnyi7bnaufDYaYcblCkQqzaarbL7hFiq
33Yna5Shm4hTguAazFIXGURYHnK4ZOW4kUjpdkAmpDgMo1IlBkap3lJf8cJ6RyI4
Q3vhHGAGKQajTxBJ/8pQC1O0TfS5eedbMvOuxG0M6Eu3l0k0yE0vJhciqGrzJw+Y
9bxosw4N3uxrY8clvJXrvMiECL9nnClyTT7hO+rkix0fWIWrJ+0S3ILEntLuCL3n
qIpvt6Y1F8jevUtxyu/FBlVrQudPZ0NLXlQ06yM/2HhowHGQ12caefsAUgDPBlAY
kL96rAA/OphQlKnY2mUKm1btjtz64k7xRHM7gdpAI1pL8K8zHuYQBMF28eT005Cs
tw3V/RvQ1PABxmAbD1dXJbKPhkG2uRHZr2hgjFVJQ8/hE+UoJw8KVdX4VGPEBTbp
ESCyPZp91WtVEJzaECRr2cPGHiGK81xfn+R+XtYuKix3aeOmMxOSSXytiy3W84A5
9sWqTynyNrLYTPSuMWJW1LPDQIrC9eEq7olN8e2JWZU7Oc9wheUXxo3bC3n1XaU7
/m5J74bNhIKgfoyaTe+6mnxTw4CzqHmu1MhUAP6YZgWtz9wF49OeB9EF7G2HK1jv
du7HA8rmDevBEzEHuH9y5c74A6u4GWribdKhuhbN4gPF5L68hA3zhBLDB2jDtMzO
BwiZRjPHYW5FEQSgHW/+w5ooeJKnHoyg35f/bMybmhTbb0xSglKdDOzr+ZnNgo39
kWIi3MzjWphdqC+G9qWOwMtb4WEXcsRPmbxrd7a/5mrJfPRBPQb/1RTIUqFZcxqa
hYjkirCgRQwdjZ71YW8MqZNk89mFFXkvXenx5BmhtwltaL33r0fW+26fZo7kVeAF
CH2XEN5D5iH6k0HM4P+nBgJJmHzE3iUpF9/VnQrRkhq5j3ooZbMCDxRGl4NXQqkU
7G+hAyRLTMNU+2EqTymzSkEY+jODnmX7l+1mWYTOa09RKd7p5kJr9A7APL8y67Aq
ump0wEEsfxDTn3HD6wpzRY86ka8weSfRbes25sGrTmGV4tr91znRZN3G0Foi0y8O
KdolJyy0IzqMPQr+yYdLeEnBLY8Ot28+fdysGA71Z1+wTgwMARmLEITMmxYOwkES
W7/x9GJq4wrbs2JecKj6X/+z81iHFtEzBgW1VpcBBqf9YyOnu3ABsDsd6qOh3oDl
WwdX2HEzDg3uFAKJqESVXtM5aNrKmu+yYW6cWi4RfJuGt5ZhUrzw/BilxcpkInQK
wgrRhMtYhKpHaKeTAxFtnYBgB3maj1QxG9ioTk3Eqa5e5BqTj7bBK+Z5S4u4xOQp
Mu5X526TFhVtawUUvrcrE2oCXKfR07jZghQzDq7mUfDMsli2N1yhe0bQMhfwGMg6
7IjbCLqYodGDd6o6ycSmDipDDhQwtie/Za8y6IONx02wye90/hxR1MJwdvwmb7FH
03ilhyoB7bnsSyCYI4EgEft8Y1IkWRTFb0gOaRsLxQEPHZhJFbym7P0Qr3As226F
O6rh3EgafMPVVyaAU1Opd9HzZ0dkyZZpVNkNo+79zJsBPOmNRoFETwh02vGOv6+w
hY6tY6sgf7s2p+Mmh41fKGTjjutFKCPZh9lkot740eF7fT3f9MaQ6bmBDZr79pZI
6F1InARZ1sLammnq8DSPoxuHkohHrmu1rM6DuUk9La4MmUhh7q3YuoffnlW4dxTZ
yFlj345bLTxRhdVenfeMoKAtyNW6X5OGt70F73q22cugYiBxuRuvGhGEjDi6NBze
iSg6d4CcvNzl3Eyhex1k+MLngZfcy1kvUNDt5uwa3iION3kHcD56zcihMYtDKpil
uQWtnCyuhrEmJmXmZu1Hi7tvztKYhPO6x3mY4WMgYjEm4/o9UF4msxBUZ6xryEby
LufP7ZK1wN8kQpBEZvgj6UetsWev6n5RrQ3iIfYUEK3HtqskUanEJ9TmP3ZWQqX9
f6tWXtLivHUqqGwbni+wyb+32njGqVpNhCmbhszpg0ZHDi35ZyE1MJQU2FhEnGGX
imtfP6UCfKBdUvEjo9ATYsRPV08jp0L+UM64HyKy/qvbZ5dsqh6iw8IGZCO+LrwU
YYHIZarLTiXcy9Y/pF5QV14qL3miglNN3cvRyvOR0RLC6IdfS9VEeh4kuYekZGxT
NLl+cIQAmBBvcotKtdyhsIrH2ESygiTYAGf5lHnl2dSLSefRtWn5dJWuxyNs6Bck
IhstKeCUzyc27anH0t8tUel5Lmd1fr+dCmKGXrV0ax0tcY/kIXfCrWuMzdBOMLcl
mZa/2u24tRnHG7UYgzo6f5tCNlO8N0Jss+N/vOLk7iWl3dWofdKHYZzWWSNJFGWy
b8B2jCxZXP5IlBMyHe0y3qgHgzN2vbdQi94T0vVdTxj48KcFzuS0NDPt7P6/HMdD
7SPPZWp3rP5kIgW8foeA3fS8H1XZsDgxWnowk1Jw04MvokjWUEZBQDdMCpgaTm4i
B4bfbs8O7d/rTXrg9UFu2OoT0O5wN3MfAoRmK4dWgZNKI7Xc6q9N5eoP7zd60rRd
SfvMcD425dCPgLIHVPh2WaTClo6s4gHK8jkelUiVEpOiQQW6Nc1TuWJ9qv7giQ+s
OXpnLXPta1Cn3rVQB6vhoiKLVpY7x1N7bDYf2NYP31y1diO05W40lfk20DWvwuBv
8YyI2+9ZnqiQ8Qppjsiehx/L/vqK6BCRptsDnHwfysf3j+vNQ0EbA90k1onvfRGO
3FpsPjajgFHmWqUyKqZF92TrwMvShrEq6dZ4U4vKCbep+71wVNvvyo5PwaUorPvU
I/5OUw1l6ih/cs8FIfMwVa+yn3vUDV/MI90fxX5O09UQctTvzOtfqp8F+2KtL/0S
3mQvd+aaMDAc85mEedOLQP7TGFjZTTKMwAOvn4WnpHyf4WINfRn7PSBRURFilxRM
VUaukLEhvPd4ySqMEoXYSJ/AZiUpF68UkIJdfeJeT7dEAg51fCvieI3bie3kZJKu
lRCfkVDe6Y2YPZO7L3mLZtxDyF8UcEGNhqx0RxYdUz7CfiPp6OQUZv5ZzrecbVLm
gmnNSbGBSV4LfQbZngjZ+v+ds6d+w8zkK1yEuDjaD8OKAVZTB/gXONLaY0TLbVsj
H6RLJEhf5XeedzM2JUOFO55KLw5N2/ETOp9C7Opwbb/lR+3GS+8GHUOWTmciYi8q
d1ySU0Awjqt9oEgk+gqjr6JHB3tGdZPOsk9owEKhtSGX9DFuDxHnmPVWc92Uk8c9
05s+2jc8B5CCiAEOX4644UryH17Z+HQqTmZn+EBN9w7VG9SqxmHa/ozUvnSJCoGd
qgDFAZyLM6H1ZvcbLiWE9jdyHvUE8svyOZFCgm6/xe90Oen4p5DAqCgszJlsVi8B
7gd/XEHfNjiM2XnjFgGzm9kVto6AZqR5fE1AWl/06pCY4XVyIPEN/MCFypJ+Im4A
x3T2FIEv1ZFc6GIsth3Dzl+fijdRnLEP7G8ldIFW82Zq4AAsh6FW+rxVv6ALQEJP
ybzf7n5v7Qzyj4UYWF4ePE35WEeiyBLpDL2EzHpXD3DNNZpDkAhaxKdogDpf35fa
EQSjemchuj2eDKpq/bxg6+sXEwpGN3vToiaGXN9i2shGMOjweNEKa44/4M5jDqef
hArMIWsW5oP6GzhHLtCNPY7tXTSadFaRGtm4k6Ef9KsMb6y9qoC3Oj2Z1YNYmW/r
WXup/8xkk7Qz5Q7SrkT4Iw6oSiDEx2rVlfYmeA3o28okjzsRVBS2KUeDu5QAL+FS
uCsOU04Cf7Q+A/CRDMdpgTHktnqFIC0J/xw2Ezp57+HVGqKHH2TCF61JvAA+MLD5
uWd1AC0ZQvSAlgauLsNCjUw2EXwmhiDOAsHt9RW+VFfHFiLww2C4Wiy5EOwpPhgR
Qq2wri/xcWgFpJbfUSs74cuyH8SLHzRYeQQjnpcTa7wMGB0beHm2Ang977UAz7EV
PaNecYGlJgb1mnL9W/gsHqjOXDrKJhbG/0FX2kE6jWlFJQXveajn/FGHldDFUnVK
2Alsda/EpY4TXllxloNrtJkRyoKTQ/yIjShddM71CbWSVLIZMfwKGbbfuf5A8K7b
shtaSauo5WT/+0kwqbtYbj/0OINnLOVilV7XHoSRXz1V4F0MkQAVigqbw91kU6nI
aCotewTsJ5rGzRrZOCDoGxIH/NBvbVYe+ZPemrQycDgtyn6f8myf3ZTdFSsSaXCc
XEmpiyVJYK3XTOq3UqS/CRTzS0u417+2a4Ud1CtLl0gAKw9FlXlfS4jGEJ5+J5Hq
Dk/oEJqPGek7fycjgmTzejpz4WgPhCL43O4L0Fg/cfQeHuVAbskWg2ATTpC03NqM
8We3WDapslDo18PbIOHnGMS6ar3MOMO8AxBWvzlSPbxzeMVb4n426KsxTbywOL2V
zcG6w4ZRcCKekD6RrKzkcn+FXRvQuOmIV7TmkqAWc4xJ0110rsQdMA82mqbOMSiU
u62aeAOSHWlqUP9c39RZrEyvNI8OkGPhnfsm8n8q5ic+In2Jm6GFPGics14olBi/
rgw4YOa+qXsd9M+59k851dTE55+0gFJhpms+81JEkvnWz272GsZYcoVhdqudOLac
4PrihBonnBjPWAtemuZuFKgJ5yiDXW/rzRuky/M24vXN8reJI7LT2pW7PCbKHANU
BQrLFPklUciV/NnoEyii7H6ClVouPznsvFsfoAv9jKYpRFAbioql34HclQOVgaw1
AloCZeKNc9CBvLMMzFQs566AbXYTbv9VrgNWSlFLoffrr8hdG+CkJbWRm2ghbGQS
Jyvhqsn6zsMMviTH7WfFqn0S46DRrfU2lmAh/DUupR/uTgjt39V1NH1cdYklyP1g
QBpeFEG5udQrYEYmKyalq80+iFQytMkJzCmR0UkscBr/sObXTyKvmGOQX/yfuxIy
hvT/9OEyfmeHeY54xXtTb8aPdk7ERbNVGLAE9eah766CdihYO8dRYGBHEIwVTOTA
2a8r2OV0+zKCzQAfLYPSdeQ7vBKTEneLmv61df2wDVY54H2jY181PVN+TLLK5n7v
kZYRoYju0cPheu7/1kCNi9lCGQu6TNr+WHuoeOY9TWJPjQBcEeIm0w03snv8tyVv
fQcXqXqXCm0atHfcL4THhinc4rwJJ9XWdiPdyKOnSVQO9jmy5ik/qtcXFwyJWph0
ITr0BKQd5V4ImVvoYmMfOu3nIk38yBZr51iKyw/uQ9tFuV5nL0qoA2L4aXZA1Isk
xB+JlKgWHthpGuSYH2fF7Z8U9JVOQEu+5uzQMZT49KOm30slSi349+i8uv+JY6UG
1xmrFp8f+hM1NCkxPebtbr8/9JmDm/XwQP7vdXz2IMNTp4L7yAZFmCggXCFrVz/F
kj4M1fW1qZ5h//QDMTlDh4pSoJQ8IA6loGcdTNMEve+xjmCWPPXWfUYhZVsMoCX5
aXe7i3VE27BBN+WNmCLmRmHUC3WJqwTaT8tmJFicfgBAme+6BaAWTD0snpF2+9cn
o9CDnwl+M4GVGjBVkPffrK2hOhoJZ4Nvx9ROJP91yJH4Vw2gnk1NBWDaxxEXH0so
++K/EYwLAyAd+4MUP0alKZjQuF1lZqrWR4yKGpAHziomLIJ05QrMdcXs8kJtEtd0
HxuUsOWdAns7eGf7VXr6BMvuejZ8pywDofWoqCUIUXU=
`pragma protect end_protected
