// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
O0JulkgvoK5Whg9T0eHR0kAiEPy2cCN8kafdhrawxCtuJKU2qb2iJ3uZnhnPolOe
9BvcD/KCiHr5R9RrDbPZLwhif43av9dPZLNgPTbMiwbEEGz73evne01MkPONarQ1
o7VsuphyqFIsyPHPQVjhDQuPqYPbPFikXcbji0kokO4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29584)
qmwpfWl/Oq3sCG4BhbiMvbtRd8qM/sqvOLjyIlf0+FQF+NEd1qbr/4Oc422/NTKU
WN4ln1fVf2GnBYXB823euoN7F+4/Yy89byXoFl+mEcpGl7K6JC0SSbh/SFwLU7gn
bEQBzQ41qwuRUKgYYgp51JM6fQFJcfzs0q9nKrjg969Wrt0Qdg16FP+x6KOPLKiU
0sJQ3olVL/+8Gt8CNg6DtXGu//KF2J3cPulVlWrIK06MRqFcKmLVImIYvW6KfFss
EwCUXqoGWTW683ngGQIHuZkxtTDozQ5JGANfLW5OPvztT22nf+AHTHUGBrYZCCW4
sdieHG5RqERJG4wf2cgNp240AWMtKAIIZYkhoKDNS+DoFprdemGaR5ShhfODusMw
y4HW7z0e0tq93gvswIb5ijqe93juI+fiO2FgAA62X+nx9Ir1VAkdqCMWD4FalGM8
5o4/6iEKMscKgGCtjgoAk6IlNTu3vuPnlKW+JpBjUSkSLHUTfGLVxzYiX6t/jPFV
kYphETDmyA2r1RKDfb5v83mn5LgM4ufK/rpp8N0TZlXvLEdmkfvqGRgnCF9svtyO
qMqFTWdTesUj0jvXdsUa/3hMbhmH08MH/Gu2rhIX8KWF+C8HBC0NKz95gmmZaPUx
8FXTlXAY8bT3QF2UIKVYO3fx7RQkpuEsNLao4ITDPHCjQizCHqzT6a3E4VAdVQNe
5xSy5Y242pS93nDN5jn6m8d4dwQenPRFRL9YqkfePrHhY87S2ExdAMCMtqAgKbw5
H7ksYPVOfO5zH8EfH14W1tX3uLmwIKvrIdhFiuseIPKwwAK89uMr0bjhbPzPaQZ6
VAOfIgt/LSyfnuz+D7fBYUdPBSTLeasD6q4pZ0k+kAWKzaCJq/6crQJNUtfn8qdD
qeswH5eaMj8Ygn8CKy8uwyl/F/cVGjRCW9IAUPGb8YCp+zLRiHNaKaN2k/jpBjln
guFld+9/HHZfChfNQwSGo8OxWotuWBLmZfZbR8KKpPjAdJtos38s6WDE3wNPjujs
WW7Zpq2M9JzPqWQc4rOI27p2xSiXeXIIuRYJfoBm2UawjKazShKv2c5HA3ERVw0g
SE9Zvnc1H1yNDbWiRbqvplJs+wJGuTwe0LzTimNEHzAcqASENsDPbJCF5j7qv4P4
fkNdxlcL2MhLGDbC3samt7o+bRVwe1tqbk6Oz4LXdtNszn4VZhJyGXK0EJxldVu+
JcPhZ3+w237xW7h0EXeVEjeRxIxjIqhm3HX784WmCtHrKb/7boz0990fUqtwJo1b
Pcp4By/f5NUMCSTm9QGPuo78INEiT18SovHu20kx0+jxN9HW6J9kwKzNdQ8GgvSI
7pFvW3yfAr8d7MnctxkQNiNMptVJSjHObW+cdGhM+rNtl97d9bRM2oGK6umM7h4l
VrTKvL2n5LnnCkYdMDcX0qXuTHlcEKz8WznEmR9CzPXYXj/I8vcUPH+d9Z43Q+5m
at6Sz+WUTFDB7Wmf+GuMEhNP+mHlqP2STrkHnflH5gyy4E+iV3jzht+yh/0FDFKv
md3+JsBRJkboPfzWHVAe3uNi8Br2tRWOE7eF9jHhY1TnvMel6IhtbAUk3Wlx32N/
5S5Ng8sjzEMB7ZmV67sbb5JucVpySvJz4TvrYObIX85CdQbBqkBdfSndbAVrAgVs
R3AYkVquBS/xSKsYu98Wu1x+n4zbnwrFW792QsPuXI7SuZXEvZ+a3HdPlaXMhCWl
NKJMYSwAye2fSBRMbJIpCZqXp/A0+eYlZmv/Grm5HSvk6WlMl9WSwWsxiF7CTGlq
CAOuCFXe7zw0vHZlEIqwQDC1DVJZ0tOpf6MS0qVABQmaIJTSJxVDhVKURpNgsaTG
i78YlyzXCgCyCQdfuHVl2njy1Vs/vdwpnJL01J0X79DQYwc61fnfB5zQwe+djgI/
dvTKwPrJHYuA477nKub5hoa1x7TjD5z+44P9uNML638ubpJ0b63n6gdVW9ANLPY5
c/OygkW9ZfEsNkcbp9TP+HWBG6VmvUEg4T+uohEIyVWM0UOFYZO0Vc+J2zUx86X/
EZJIdLCCH7ST+yJKSY+zvpaK1LQFsCWvq82zSTJk5hEhZZ8LE084Ff8I5qSKJc2j
0HW7LjKf60WGpklQfRCkrbbLfaDvuLNnAv5WSX33Seqrcp2qKoP/rpGxl+wFRoe/
SSRBYIw5ICdnKk07dmYnUstdWi9X4Nv68PFyrYe+8ySwbn58U/qfFeMqaPOryWFh
hN5qiiBbWQ3EwFYv0NnWmo1jRyGvEUxCFCw3OsXTDIMSHrcxVVLhf8bMOhAEFP+v
R0kg6Zi/jTjW8p3a2qSM1JDGpIh6Wv7hkuHxFV9NVsC1HcPfKJr2ICLMeNBo2/1f
B5R8oY6mKl5BmXDvQV8FxbuXgyRW/JZpKXLwnyLNrBsEpRzjXeP6S7A8RHHWFeV+
iggT70Z6Ukp68ksN79Jp9AI/RxElrsaTpIIhTuCT7SYn/Prqx8IPsRVm0fTwgfW0
38K5WgMfVSuNeXPCruzg2saUXGzZAKBDMie4ikFrdQ79xVOyijeGzxc/y5OW6QgR
MiZNva23wlRLCrWOgEIbNsnAxSHj84hZ3hTMz+u5X9MG/YK1boQnaVpT9jEiDV7L
JEWR/xm6Irk8VCckn/vSHl2X0Nfuh+3GhQJrIrSZDj7knvuyTlDqA5boaY06kFNc
BOSgqup7f+qeQxvCkjpcuHFCZ26Gz5aqIUXCMKf+vr+2eQjwFmfSfIgjem9uFa99
8CpI392JGdS1Hgmp7QDgZ3TQi2hgOjL12/XH0sg5x1DXPM1cdB8XsmV0PchEbNpb
010l1p1RXiNWb4MTwv8VikGGrZBO5NJzdJ2V70NdpnFuS4epBoTSHvcPJAlyshIG
wPz+wM5gFIRvxzvOnh2ttSKoq0o9Rq5ys8uPBCNhAMseYm0ZjqPq9wmBv7CngVhC
VAeGBApW+ExFhszs4d2gbm1Ak0U1D30aq280NM/oZ9iBwgU5lourvhacQrNPqD5h
UhW+kPCWIkhFyDigkDROiaI5fAoU6bhvgo6BKceQqNm0HYtkvMrIvRVUW1UH8lU/
i9d+20gACKmXSfDjHEQNQAHHvVcQ/twPU3oEbcfLkP8kl70YPiGBGphGHwXiA2WV
zUmUvWC+mQZaW9WPkelPV2u1Bjfp7vaZaV0MuhMgv0P+Zx9jKIIp5brZLUaHl6UW
aPEuROmFJq4HmxmTfXRZ8m/4qEiPPci9jui092kVYMk4Lfl54PT9QK/SHqqACUGq
Naw/SNQ3sqwLPGZPpw3NTp3HQBfHRffKAkvPU2aZt1N3CAr/t/VikehlKr2Fvs4F
+LiTJYRMosuxQWEWUdpRPBI6uXIZCYhzngBE5F4B63ykdLgUnInbAOVyem2PRssS
+0x6A+DJdpL8d74HycRkjTZr6thbtV+0QkwpxwH8KYVmVp2yWQwgZoW5Yz/IERDh
vuejKehjYOTosA9YQCxXQPSHhAWS1a9BaZrWvVTlF3PrONUXE3HnL1wzQHqdYdsc
D+DM7iIuMgW2mFkau6WQWSIzwi2Ijv2BZBnUaPjd3aEcJA5saKEhnL7/NctohFtU
LPf4pt6Ih68RABZuxfGSGxnN6u4LPj32cz+Sp6+BrtvjIZrhetowhEbw+UanCL0Y
WeSDOurtL9UCuazViqddGawFRD2qaOP6BhKuT7lQn9lokcB90eJ7mZnjoC913Gu1
IdvHf3ficcuXBN+mNhnKKTTEejaCnXOrckeBbN/a8tue5qoLTezYeYpDS+OFs2jg
nfX3n6l1q3ZqtdVzLD6saLL2dBY3HH1sasybb5QBxFXov4TEN6/ezJa+/mqYF7M5
7v+SXtwDINUCp75F6VToGdZ5hkX1nTWA5SAH/BiF/PSvgGYwRLe4mQVIqToWyGqp
LHwKC8f9OtF41sjEj6QN98+WJlvYQODgenhKRJU4A6TtIg/JF/pcnzvV9OaekMBu
B58NCp6jMtuBdnJXaJ62ARMzysOQU0++FERkLd1BbAZllP42rpEM1xkAFxVnqjaA
e2y2b9PxafnC4Mil0Z46jcJbbkw24dIPeI7mGRPZoBjPj8iEHz2DFa/emS0NP/Jw
JNsYV4nHEUAk4fBIFwTk84yyGJdf1ANTrzjfnE82U6BoeRwTIlcdyNCK0u8ezh+o
LiyCx4RyWqMAXOBLZdE4gNlwynY/q1dlEvFiiw2Z8ODifno7JXzU7D85Ur1i9zhF
BRnfH8uaYngtQyDS0rNSq1YozVZ7PgPy2Syg2H2xSyovkugDKWOZs4f6bhoxljgM
OHPi23Bu1mGU7xjD/kOP1J828T4T92Sxz6vjBZ6mBK9kj1KOcYfSNGdCMM8iJ8Uh
IhSQE9G15jN2QCB0CIRholIQF8LtqWd1awQTiuWQa4pXESWN8hdFkesw3bZh9a21
rg/4HKEISfBz6dREJvhTjjZ1WnMfxOyqImlVBvMMqEpHYMAWOJ1mlXj8Ht6tQfOf
1BorwSg6lyW8mCCr9OnlgqnZxe9chYMnr0FV7ai3fcgpIsnquz3A2qwe5cnwI9Hw
skN42+JJ06+q20Qj6csHKNfM6FC3rOBjjjNEcv/GvqWmjqDxxBmU2olukKyppDer
E865rLmgl0LBx/HhCVHZ7B/uSiVLD0ZB3BC74Z3n/KIEa06lIBGmjvWBrMAY54mr
UrDIGR0dtMMey8O3psdzzztZM9U+aGZ+dG5MHQn68FyMvzovpjRHnaeElyJ+a7QR
7G1OVxKzXO0as0/la0DzjEU1qM/r1INX0JNfqoqzU0vuwGJ2hv0vQu0KsTr+oXHk
HLPZoN7FrPt849KpBDbeeEap62ylVmzlkKN/mUkNA5b3t82puwm0u3ix6zEWXtk9
e46VlIAG93cVtzANmHvjtywf3PUZuwv3WIBFIVJRpvVNjyuPJOuQT/YJ8z7/i9Zt
NguTOS7ZmpABo92HnTMPZjrQ4Nfx+PGsY732eN4jCEGO9jI80rafZNpTodJeJJwN
aoch0BoEPAS7l4bQC5JJQbq5ga71LXwFPvOCa9ojSPlDJaZP9cAZppBEUPbLV27O
VADkskw9xaDITJRsJbVCQhMpQjwB2VqhHyVVLoIYGvxsm5w46Kea0gEh9bO+I/rT
3nE7I4MWaedaZCvKCn5FRKYwj1576Kf4nEp7AHamAXCTsBCuF0YdzoJrDEudhfnf
hbpvO6kMXIANaJWJS0jHP44Dk63xPr26+eSaPI5wPARICqiFlC0jVRKgNZf3wwjp
9b5+e/VjTzRMPwY4sPFg2RdeAkQQLF3VhYNly/BBqRPasRrzJhSSULwrEQle2d7q
DIdKgjrZXKj3ripd+FRf+ATFl2gobhHb+W9FybwxiJ7PZkPww0d1+A++qWJgiqk7
b/n5PML/XTnCQYHosBvUZlnOAFnTUrkUfDdvFFeXX7nPkc8q67MibZ/zPUAhWje4
Zuiaq6Kvu8a58vGV6z6JfdimBqL7Mw8gwUm1PWXWBM0EiuZD1mjPyKklXQjlcM8b
YZF1FTWeaIfd3k4SkwXXoDPFEz6IG1AgRUGGUYpKwZ8bC5Nnw+kXDiS9CUv7mF0/
ZpqmGovOxbV+5H/6Kv0Lr7M9g0u6PQyqxEksj00t+lMVFjPQKCItp7Syu4f+vs+x
bs+wNEZ3swPSyriunAHPyRsrCL/hZcl9nxcbMqGzTJtzVTm0gLkPVBwiI0s+I9/4
FEGqn99s5Nn22/2ewNnhczgGqYrcYSjQyx+1HdQk4uzD8NXkMvZTeA74fktvNBet
XAyLEcCHohkRO/78qwaveJ9XElu0VjUjn4ZpxraOAQZiFLX8ZnQnBHKTIXWwUyeA
ertJDN8h2u0UjS9H3e8y4N0JOwDKOM1pVu9CLpRVhMcChmgtrjnzObJuN10/xECo
7RZgTzBir65MLIsz3qXsYHqcOmVmV6qkew/jUF39XDnTqd/02lCKNWdTXhNGPIcP
ozg87r8oDTGBgEbzKHEFtAMGUNX8nYwYC2uEnSh7b9+wbZADao0LoTh0xhOLI7+G
DI5FnAJqrCEBAzJoLIjVyfH15MgBosquRHXh6djpSFay/2uv9YipzqwWR+/LLw5Z
vNJKNRVLYHoBjh/n5rSGTZNoFc4RyaXMl4fr2F16v/HMltUrZrwUbxb7lTJsZU2b
smFpMdtCPcuD5H4btObBMI3PyFb5fD4OZQHiUJn+Nbk4R8QmRV5VKoUTNrLFpdHu
ZNlyIeSThCR1bwIj74Kn9pMfbJ2bPuTORtCUGfW6WMlDJLgcNIKnKJYkDerU4AuF
FOoeWWF2fJGnyKCxBQ/h/tsKK0KXZm0p+K73dlyqKZ/Hx+OGf0jJAL8bAocXK8z6
1LrBs8BXGGrzJXE8zGTVuh/VgkXJXrDuKTOcBNvWQiFYeI528QdSGq5xRnObnIK+
aWpLOrXVOcpfJwYorErJ3s5A6c51kORVzysIlCO6hD8hNNi5fHO9P9keULCmP5PZ
u3KR1NbsS/LhxF7Eeia9vNJO9oYkdvgovuIE3ErVTnWWYbFkOAnHApevkH/tEaFo
PSExTVwEdnhXCDUt80qScDulS4ukfgD9bEm0ITVIvPRy4ItDgHUYhSGYCAmH13hG
0cR2nlNBX5yuExPI1kG/j+6ZT6gJUNDcEtciYmgb5Sw9AVvpQ3ZPwLLtwKNuJ6Uf
DjQh7VMyAuxaivY9kkSRXQbZPdweZyzaf4C96mDSa54oyI378n9WpzGmHR6/9T1T
lOtkFFIVIPjJ1vwaEcNMKi7CqQ3J2HuGCgvqgMNRYgjpoX+vrATTQbIsMEFano6p
Z2qPzCqFMwfSmq3U6eCboACuVV8FdAc9y014uHorR8+9Y+ugmAsrRNMaXeTe7oB3
IsQoeI3Co0nvio8QuX6kJHbfpxe3AZo6Q8THZFo8NnZtaHDQC/1Q9Wv4jo2LJ+/1
4f4oJHHAXzxiigXnpWz92Z0xrmiGS4QCB6oTo+KKv+5NkopFSMwp36snGEdSjvlY
eJHa525pMyHjYR19aqPbzbFt0cxFlrFc7QSOxRrFYHLBNurs/3lg3w5xVKUFD8cQ
kvNdW27IFDFRyIPMf4pgSSoDJhs2sbnh79q9so6vFdtIQ6R8lgHanM3X1KJUBIkj
xxSVQPX/xPCoSyQuxHYE31bpevzq5qMzEXzBKKnlmy9oSwmgxy8/67wqDLgKtMY6
l3zY5VZwdvnQSJb6P8B5BgI+QJVbK6xqF9rcexOWcVAUQUgIVgcXyhLvTexqAWhp
eS1ap7mTcNvYXxV6bjhbQEnbT1gXwxKUWIaJqcTej3Bqnr4JFl6ln1p4Ycoc9TXX
VcAofY+PcbbUHthVI1gcsUFEIntjb8dIXjT3LiR5W0Y40nZU6jDmWjfu+/3yz8DB
1n9mLqMl9CTYIApzkzW5vf6tw9ixsEQ4ZeOu79KdfVB53kvz8BEsS8GwF7GvyThh
/0R2PeW/hHxlvyHXvuymXaEvcz+fVJtqVWMCTyogEKJ9XLzf9mc7ixWCh59J1EvW
Qd1lGNS3eH7JjAx4pKHUm2vb7jN2Jqllc3BcKZMg7DTD5PUX8oIYmIELb9z4MU7u
waGi/yLJny88jZ0YUO57FrqXiKv0s32tYK2MTmM+rRuIpKJaX271x+bVvNfQiR9b
IW7iLXM6u6Y3UFVgVeqGcnp1pa1r30FbijYk/D/4giIA70Hn+59l95MM5va5aM0h
/V7emOo547ww8T14q+jTPTEJ8a8dGJoUPw3TlVL0bUaW5iQ8edmMr/D1x8HwTR53
ww08T0GYloTxaBkYMtC6V641xg4/p282f4SXW+0GGUAgvmztXVDb9ubeiDubUPmv
R4PCmR3m+tXweEcdDEAhB8aj/b17cfGvpqeti9bPuZvUqn+0wh1rqqY5roTtCCWf
eqFoXyP2HN481x/CJULD8Qibk5KSq4OXx5u7CRXC03ir6cylIla+lCWaYBw91LtQ
/JngLufShG1fTvNTVja03Z1JxKyQ2ZTiMAG+ybaBgkFf5hBNekH5OBRZc/+WuWTs
+7xNdor43U5A6prSKJ9szg7pfmBdm5kmutA2GoGbSx3wteybflTR2bFcTpoUJfAZ
zAm1mLSWCd9w4Cn9oAvESvJ1J/4/L+KRo8wfJ5ammNj+0AJanvD95ZsJMImsSkuA
uR4zhkQ69R537JElTsoLbBVfNz/fuOWUUl7cHHDvp8IJbHg3lW/mpQtIVAFbBHRN
tR+b3aonmGhBJ7X1Zco0Pb7qkyqOcSPqyiJ9k6kG1n7XfGXbQkmKtat4JsJSYO5L
cGXjI9YcI30jzaLiJhBZbvzopMZw2G8C1J5fW21nBMfM1/fRmEkmZqgLx7fxDxHC
M682PrfH1OMQaAID7sQlNIZe26gPdVbTD1nLAkLhhSYxyijHeCG4nYYL8zRExX82
HY7x/ZqQjRyXuwResSIFw7PM1eba1SgFxX4RcuyXm3s9ezs3dQp3adOFqZ63g+qf
brdEBtKwCk3fltWGq1xNhXl3Qz20TmVRJOVSMGMprcLd3mpCRj6i2o7aPwT+4kZc
1vtExNcd2J4fjvIQL6dIDavcEgoxigLp4+vxpa+qcOcZMoSzCqTv7flsFslhhLmo
vStJTi5aoxuRecF9jfiPI4ETerW4kwsKbrdeXJBSTBfHAT4FW+UO4k+vlTcnR/06
7IX64yVSo6fNXOf/kIbxwSyWRJfNveR/FqWzsgAM+BcGZdyDoFgK3D+wG8B/uZD/
eAtLHHsv/1lGeCYiLJwGvu66STZjEDLeQwVTZo+Wjzs/jcXWzCkBiqc2fdtIPAjN
rV3z6zvwgwxp5cVD4rnkSjbQ5Vk/A4cziDXuGMg3J3PYC4/Gd7oUGMGgEmN6dqfj
AVnymRAoOloCoiz7qRNEvy5Ljd1DrLDkao9L2SXU3SXOwISuK6nxNyOvXbbj2MAy
TqVXw4eYXBU7nt7WBxO4H3y/Ec60/S84n6P7chaaHlodDE5wwZvevQt4RaF5QAfY
g7QqkBCnu6rkKAm0IQUAbdFri7iqjB+2I6zN6fmYAQNF54xC3tdP36hYH0RNC5XC
uxpHCQmT1QKt827c82zAiYE5/l5bVg6Hlm7HJYBY6E5IdbdJbOgHOocJBYuDh0RD
NYqL2vloumUbByPVWu2Ao/QXFpmK9A7Nl86ulmRvqLV0HMP2F21WvztFUdn8vamL
Iglob3NjRWsWYb5eL4bxF0ZEMSU9Dax9WWxeij3dy5cHpzP0Lxp4pDM+jAHpsuQI
ylkx1C19kmDs9FuunnbRo+wNPbw0GslR0V2HEjlXD2aB4wBFwpKvm8edAs18Ki0X
TWeKUVvhSldeF8TUWU9Xp8w8P5qhCWQ1lTjgfAVWGySO7gJ2uaCXctMpM4hk7wDn
5iIAtCjEwpgQrA0vLUMgRErGTbyRoxzMT/M4D1/dlraxQK0kDZpor5aNzz6VX6mU
nv/vVVpuX66GDOc+dgzsZYJxXvvmozb1TxRQowftKJyxn7twk3T8/LRVlWT5RI2u
3C2QnM6kmlxD/Z0mKF+9f7wQ3ci8TgSfq8cp+i6PrhG9mYEDVqgjMTHYtkR1xA1f
DimzQpEtEhuMRhkTK2ksZ4jcAWfnrHm5mDwQtM1YE6Dkjnr0GdNgd3OTncYDjwlr
fXFwOdvBrH+/RaL+eLPJi4n7cHDnEM9UVjOmqRSWMvluobONC0utrYjwvE9b+OQ5
U8ey8pzrmrVKhQGNuEH4UXUWo3xKKXmBsox2Ea99pmOdigV+R4RpSy4I76UH9op/
v1NGvKHgc6jToVcUv+UWZrgrJFnHCl9+MiIVSB4+gzqBys9H0tOzufgRQB4wVSZm
wft+znjPadGX4qly831KsPtOQrOVr6+bcG0K9ZMMc4RaeuhKY90fLvlDX7MROvyX
hGrEpGl4nyu4quXIhYk3qUBLfFlx9TglftSVOuZH9vWgsKturcL1g/xXPBwVbsTk
Ito1ggxq+YPsow3ieoVesqCeV/qQWPlMv0p1J+F80+G3JBMzQ2PuLC1/NO+ylR5J
MYol7BceaK3tE7ldofMO33M1NzcD/qBEKDSj9uqmfWXemm7v1uHofrTJacC4wnjG
Qq0v3LOFeEAS/XhPGiafv4M2gCVi/cbWSQXvO2EXQ3wemGHwglNjlK92LJo4stqc
WYXLJD3PI7QkD/Xb2IpZ8mep3/g2fszkyNNUqtQb8YjRKf9rBiW1mUMq0woYeebm
HTY7FUutNqV6Zg6EYT/tthHvjRVTZRAMG4RZKvPEfsii2khqPEi7Yw38+ZJnCh7h
yd38eoxPw13uKRvEj2R7KFmK4vCzS4A5s4svDwH718wT3cE1kCoZSaEZF4vEW/zl
6JCpmYSSXAmBRsjQXM3jZWqy2fhIlhzDhJqi7+esZBm+in2vj5IP4Yts3QWUafMx
YHlxB6QlAh5ChP3w1B6ztyJeZRU5o7YWENIuDxNfiUFfiGx1w4etR3+CSAlCIFfZ
0VhwY3OfyErWHokIE97/WLDbtwDleU85j/Zqd9ADfhkP09dmVlJerI3Dy27xrrvS
u4dAxCDTcQy/li1ev2vm9Aps3E5WvOYVEsPG7pLddO4RNVYz+1MmkcpHuJQjYAFe
KUGps9Dc/bi9x7RLFvOwVRpX1rTatZ5PyseZQ8C5qz5gxnINB5JqZGWHclktSJDw
GTMtRwf/HMLafmJk3fb9uT2Ofv5RtAVtLUbXpCWj0sGazW3o6xhScnNZ/Lzxp7x/
qnQkbn2KmaGBj2mPQvtX7SyPicrh1Txcd+b3KvcOxW+Z8VaqIS4NEcOXTK38bjz6
JvryluYZdM+v8mu4jAAOUO7OAZbHA+NJp1fhwg4R3hWd+zeDpyFWmmqg8cJSCyLN
plczTK3eIcpDjB5GXzUw3npJkdAYzC8bbDDaGl2LSaDnOjwD8QrMVc5gMoanZgui
n8Br+NsyNzYcpbvX+SEoQg5PmhcS1n79dZ6NfUTbtZ9by37xIXPFedEUXx0bz0BD
Vmyn6lZZMIKlQp/6/oX/EU/+qtjnRUzxurY+8CiXJblYtgr6PIF3d+Tm/XFI0guk
uXlae+Ng9MjBML8DrtHXHZXrX/Volggzl2EDLBoOYIIy/WyVrSzb++YiumnPxBvO
6dTVcG1NOJuk1SezInwQpcbu3iLK/YrG1xPmcxq1/Oe4r+o3T3cDBDSuNtLFxPJa
KnnTwmmwneYOzQkTA2m4VNjgOtl5nE1f46WiKuZTkshsdt3blZj2scO0mJyFR+Mj
TSE0JIQs015Mmwvdg/1/h6B5j0aQRV6LnJUK4jndyobqIrx8EKpS+ijr8Sy7fCtf
7DDkAuJ3COrLdlayav+8t5AJyAmURTG/oL+CkdqYrEPhj/rOhHdWlr0XuaTqewny
12evvFvx3vANFbTeYbTrq/WLeBvYnnD8/1omfOl/iU3M8ecsGh+e6JWKz5lGiDBx
KuN3/AbwdDarvLqyPJem3JgMucDzSEDaAKZYsT+uazTwV0+ly/jlSJ77RLqZE6w1
RDz/t6EDb6oozFpaigNBKZIptFhryn9WQg6eHg8KE1nt9Uq7YKvnK32fSax4lGK/
zhNwSy6j28Gy/yajud8J5FN4PxDLlDTkuQpLVJMeWqlU1l6QlQMNumU/RKkap74+
CxIl9SfsbhGXzgNYk7q2JmjjpT9RTCNNQJBCNfZLZCEkzSzIzJW2tFkCZnnOhWR1
hwJlEUG45+ptyWzdYJcnO813bjET80TV9RanzdHaWviq3ZmzdqmSXKl/J9vEHwAa
CxQueJuUHaKzAs8Uw7EvJhE7zri1Nv8XtsruHn05o0cNuOScqkp+EolS6Y9jmSjn
2d1WvMxCWThOQT4ixzEC7QiMDx8Tn+jN0UbX/4F7RcUJZ0RpFiB4r4YcrsCCsVDB
z98TxsEdQYCFnPbYw/1qRhk1V3Aql+Lt1exiHphl/acDILQD4HUewObbDWWcQvaJ
qK6vs81/R5EAax8TDfD5/ymhHbQC7uA/CAw7O+9OCYnk/MlNu+V4Ig6P99ROmOcc
flOUaF7bjDv4M+01pkaC60bf+pg2qllqjSTUdhaULqXdb8HvrVo7/u99lnbkpz1X
HHaPXzACAwb6mwcono3jY2aJyGBLgxivQ2Siajfl2aiAZtRa6LmCuZIa1fUzLjMp
dvCrgkX1zD1qttAIJtZvWmfLYvg5vWSWq0JbGwBX74OICA5Cnd3sBzloVBodrUzg
OzkW0f4hTyfo3GNWzyk4fkgdSbLw8IEsokN5/rXsKfv9lGcP9yErV+vYCoGF+mG4
v1hKEZSK5IuFULQqbMRbZkiywV+eWc2uD+/IExHmKt8C20ll/AoxNBvD3Zhl7I58
3M5qKLO7nY6df1jIdIHCWaliRI8DqhVxLwKLJbEFKA8UFBAXO1BXv4JU8+dF9rl8
3yxUQbCP/P3GNAAGFjVBbqX2LZhv4wkvcyS4b5Y++f+Rzp+EEkEZ3/mKou20eOrG
e8l6HkAWsl5twN8DmYDYRRRiilfnbQITW0JFtv6ZdIk6RVw7cW9SdArsgVNbBizt
kXL6tN2q/fktGtoRwMeA19vU6gdG3G4pkYUiOwZYWVDbfyes44/BOTZ7kEB3HFgr
QH1lclMFF9TfNiuBWfhj2pE1HTJBFF6g3RUcaHV0GpSsyTMxesu8fLERN8iGfg2H
hsUolrr8fVrLewgMrBY5JMEQfn8HponiOyVzZ4G5nXR0yCVnf6xDI8P7liGarYR1
UOd6AUgnSZxNQoamg7O/tfGbRnTZKdykPzjXAXwmMJGRoAWur2QMEyeFpRCTjZn5
HOgiNe29j2eztfiMyLA9BZ1qa8Cj0gYF0ABG2N7dUxnnoRyeBoHD5ybSZZFQKgZI
X51WTcAp1Z27seyDcFInDgEHcj7qT3FaO5odBrnFYvGCLP1NYjtqK5T8m4EosSAc
Jb0JRlfOFDYV51yEh03mo0g6xRk6H0wGsh6kiELXqeK2HT0/PYQDSVS/+Nx/zx+G
FdP5bt2R9QER0dFeqw72xvPdZr6apGMfhEPg1vvKSaTLyp8kKe3uOPNLJWX9czv/
czHF+1pWW+hnwUYAFK967uLJioeENRV6vWWap5IRhTaXBMqfcEORPKakKmgwC2t3
db/9jb2mfGRYMJHnbCRiHjeQ7z53Bmc2ZTYbY+z40eK/F29lMVl36wtYQfoft50f
y3Gl2zpW8s9PvQYGTEvWGhtBmtmF4Pood2pNGNOYls/2xkotBpWJZUlSM6/03x2B
r/evMn4oBVDseaVhV/wKxgBWnBknOb2qthJ0WdgAdH0KnV4VfbOX5nAW81JOw6RA
m/a/vDIKQMSNCap6Y1Ne/Fp0MrpTS+OAJ6Szhao2lR9+zn4JIqmM0hSqfn7WoNpC
RXAATvDPtZsXHk3DPnLYcOUs3HsCdqcXI6XY4VQZ+j3jCMl6rtavxAYljJ2z15sE
HKcitQEO/qi2DKIG2Gn1jQPD3/cUDlCTPk8W0gHGWOCIOdzLaGNP7DeVdWwpCdGj
MfLf0m3sHcaEhrgRc+0aZ1igsaUmSogRDkoO5Z6hRfnyCXm/GpLbNHZmh3lcSyxR
iY2P2GnSgasctfErgoIw6rZnPTnhG0phBSjl19QhSVgPolzEZVH/xc4cNUUMJV87
ItSylAJR9tz3sQw1v0+ibe03aB3c+e3GxjJZSCVxoI3aoNChmQvXTMtrltrKLoBk
09XBiG9SHitrjz+X33dpstGcwYWcg5GvaKCkyudsO+eLbPdg7eqQCrn4k4//4tS/
c4hWmAyPcISpamwUif7nhGe/Gy7llYOY+p+MHGpZpanwypuTdqRTmbD88UgQl9pm
HQAVORyFhF5oM2g2yaOzgY9wox4zsdPfDieK9Gdr+qq/PG46eCGCmruERREXVJLW
A4Y0qeR0d38X1ZAMzuwIt4CVJIon3WF3OCV0IyxdWLptct01SUIz7ZlgXeg8QLeK
6Fldg+ktXfmWU8uIV0FhBzJctpQpyHK4XI0naK0FKK9tqfnSnbZN9Ick3dfskw+9
LACdG1zG+CAIATF5hXVF/VMS++t8nmDfc2ALH2jI4e9Z07BPmIclvADnnzu1F0EI
DdrzngKiV5veKKeXRoGxK+YTNGHQSMRiOVNwQ7GPhsuAbEKpNTuGpYNxBCgiON48
alQEJ/v+69DS8M0cJ7RFLoDrKq8Bxcsx/Z4YyAh2I5An14FpH9SNptceE/qvbuOE
4o2jq/9jcdXyWAzE1MG51kxJYJvBENguSrUJAWeFk8emYjRepbLZDzAq5rqyia0I
EN/CPZAGKrGEPpee4mElU8tOeSg+iDkDGTTaHhu11ewup70bCo6/sii8QDhnApwx
HCAcNzUYBh/Y5GapZET0QtAl27/k22lT48kaaH0AuW4FWKEHhgnwQhBb1DNaXRi/
c3Mogz1qah4UWUQZ35oAZqZ87zUDQWFUqScHrjeZPf44gngbembsOOGBe9tm9eNH
+SkITdRlFBCLaGPP6c45L0ouOaOhr2BZ+mMLn2ZEdH2LkKBmGcqe1bHBY1YDBua2
0Ml01Oy7cdgmoTPGu3UiSDbRABLGBZqqS+xkCjn0vYT6SYlQbvpiqVaNpxETlYNh
wQV0LFHw9E1snRLYPtnBPNoX7V34pjAvYigG0/FQS3ygd/jJTjnENCD4mQRT3+uZ
UrUqHKhFEfPZ5++SLcVFK2mE2kNmPmABzmskjmNre0fDWGKEberrX82lRnfHmOYn
vV3zYP2m9z14HSEYaCirF8jZcP1HPLP1kkJZTurf/wnaQHRv0ionpilgXHARFner
aMLybDf7VbyC0pVSRWWEEJHTqgW9Wz/wcdZiqvVPi0lGv6iTMrsi1d62LhaW/CIF
v4yOw3CXix7kckN4gA0MH0WgyfGPZTgn8PeXFuO3+i/Nreye2AxUFihzlP8wqCwt
r0Esean8A1yfywYfA1mnWQ7mtv9P9uEealGASpODbQoP4xWcDkkCK3/LC5LzZnZL
kx7IPsKUggWQFVYCtDG2cdUcYmns9smaBgu54pOSR2RJkEU58jB2VMDbgAnePxYF
SfhcwTV/MQXEMff4lmj+1SNrnt0ycG5l+qzP2iv5Blw+6U6E7P98dgc+IKEnvlPx
TR/1VVcTxVllPn+IqrRNGeDg+8sQkkGe6QFkIEqLzNXDljc/SCqMZYdj10OYVn4E
1XW3KeBRn2i7BS7REnkxx1+aC3FKk26xDBknGNsOutuV15tDtcpPtYAW8+0ubZjb
zEQHt4iDzcvQSpatFBu+B8zz5uKn7iiTR0ysRXIS7w6YYuaBNr7rM7q88o+N2deL
57SuQ9KLTvTMewavOEV4Tk/STmyACe4Gyn1FYxjbrauNNAZrKAWDxGlc2gbPsrEa
2G5bKKQxHs6k41biLGbGQPKWFw2tK8WMMwbinGqFTFYR1U2C7Xq7fkuyGnZjJ/5J
WVQgXH2LKRtfm5I3Ba/27M7X/AHFLDqS+tjnUZOkPSAkhotFqsskaQh9nXUN2yOP
lJF+mYcdiay7bmXLf7VX3EP3wAHptB+EUX2Yso8Ls969Vo4BwQ7fb5fbCnoTmT5f
Z+mgjq3vtqLw8XfScO0dhBpRdXl8CiwyLuqeeZVA33dUi/VjNriPA6pX17RLQOBL
92ARPAsiqHyYgbSkoBgBeaDb1jw2LPDUWA/ey440OLEnbW+4en7ZYCcIh+DasKw7
k0ljhDfoVWLEHnr6N4UL9oNDJn8oW3b9yXcizLQbuVimT740vGwgRN1MLToiWvyo
/rLGNIKi7T0Nyafgs3lONNrHNQM/EtDDBB0jcpDY1Y9o7YlQupCJiwZGfaH4sgBT
Xdh+TiDY77yfQBJpDY+gJcKLPvHjMDKdYiv1WxyQAGQvHGWjMd6kk9PZpeZDbjY1
DSDqxqEqXlMAIkoQEwLupQpE5hM7A6WDBw9ljNas75UUUnDdcYjZ2TCEBgIe629K
zRGYZEk0luQa2WjK71nNDNryKMvGuHUAq9A7AuUTXBimSpMvmBGDhXTyt/A8uRCR
2P0KeMbwz8JglfhkGnYT2KEVgKzRg0cOjx4RIvzDonOiDy0FBICHf8E5TgRUOUPO
F5HbwhWbP5Ng7rtINK4Fr5ofvdvOX+UQhZUTegvMOS/9mjPgY0WbvacPqbztHn9W
gxnPR8sQSvDbxO+Tj31gQ81LPKEsN7f3YZc9l0VDmM24AiOJcrpvRWekHFdeJFm9
kZGQlW9bclQera7D2iCpHRtk+SozRVNmZxySYdhtp9q5T6paarc0HKMdYplOb8jA
SCsAO8DPFM7DYN+R8xES9n+Yd9FKslrIuDIMHBBs4MEF6oncDoHoqULnlgmCXhNN
Rb1zianz2UZejwPVMA8KXRmeVZBWrL5ZuFXshMgx0wZNEeIiOC9uQ0eidBT8edSl
SgksitXrbg+o+ZF0BDfjny7RIjdnnH7VYtlO2wl/G57rUSY/pp1PFKF6Xjpo7VT3
WSAGX3Xr/q880Awc8j70FPFgRBH8DOK8uvwms1dGTYlj9qEhLyzLda6XVQTVV9Mr
9uA07XI0G15MhzA9imNuX1E5YnW9ckWMqAoprwdLItjNDaDW37+Cz7TW+Up1758w
JpTBi6xbqlCZG8zcIZIyFRugo2sG8Q8zFB/nnr8pkdSe8P32IzMhlSQkqLMOlHay
srDQR3gs+7xmohHJrdLsIMIR4SiFkaab687nYzXkzdKi+zSvlyS7JHi7ioFhGjDs
j/2EI6Q9d9kyXQKt8xvDPIf2tiqguOJtA4KIMy9YqORDkJjXVdbLKdW/uoi+XXTt
ZnWSdefkouLGZYX2bGPNVMNRCvNPjwr74b9gfWt0jWZtu88wQ+pKg6rDD0kmYSUV
jr3bp/HPWhsHg5QyJCMLg7ILm3GoXvGrd7MImOYycliQcXRZyLVNePsnpttpUwgC
tjQwMt8Ge2oJSYEyN9y/fEdVYBPz1YQGSqkpMLbnwkrx9KnefDeaQkRTUDsteORX
/hdZZPL/WzNQvak5hTxWr/tiweaMkfOZrSLWl82XIPnY+i83UOdkxaHOkZwsy2Qr
qxsLM3iotS4FUw2MqAvTRepVNIMssmoDOWw+TiUbj1s8JV0CIuMGAjwQ0/vWrtSp
UPbrcDoR9VR/5xcoWXgxOLhzzLc7Je/GxKceAA5Z48NMSzEmM3CfU/JiCYmM3CYN
xebL/FT7E3/yTOrsGPr0U71iC2dRlYl3hEYDlpUyK+UVuLwl91qLkeNiCiZXkcmX
1ph9YIS/R1cP1EM6kRcz5fMlelyMOj54QimZrKiknFw2hjdvWcnO/q0OGQmDzoP9
5WqaiO+4+/wbLGFZJck2+3yGhifZ71cq1WtBGyKk/TJ+1OaW5eDGVGK0sI6zS2JT
BsK+IaWgWdB1W+iI8oMks+M7vE6ILTGGVTmMu7vpQejGJKz+f2N+gu7bEcY9lNWi
DnZwY269SE3rMJBT9zBChSXKi3W419vNzJNhN1KfLje0f4wtVvGoprhQqq9rR9Oq
egfb1clAM9ylzRS/s+dOUGb1cvqjdJPY4qow2tHMKwfFZx2vmjSnA8fNDOAT0FkZ
3ofQXDR9AmrBeI/v5cZxZsUKFsbZjjzlbpUkAkfIPxzlqggMeAUHdMpaYUyviX/2
3bQFmJ8ziFYpLG97yjgb0PyvNHJoKPdkGl1RYuau+jhZ4CEydR8BIS3nQY42CAAd
mBekNX6C6q8001soMZSpW0yGLn+3k/+UjvTN7c+jglRUMFh3nSYRDSvjVixJBz4R
gutx2sMfQ2vHaJzYTQZgdIyrljDGjC5EfSX/I7uB1pNfHn5EcRuGMUIc191tSJ56
+ikmNvs/G+X7Eb00U7G/IUPPXk5BexSU/RPfGdwD96YvzpHZqKc4u15lTrJjHSxC
FmJKqUzAJ7fsVnK/u2LOj80eOBLLZMmwpGeak7kRJtk8zhRCW5Vv/2fzNzJhdj4z
17HY0f8i55eZEaAf8qV7q9tEJhS30F8iOphfvkhaWWuXRhD5QOXkzDp/QNkbpHLh
xgARxEmjLJ1wCVgAsTOwhJcOuLerA8+AAZiCKToOKUVIyj6ixnAO2Wya8OMd2OIT
UzlZEQgiefENhmoPEpkadHOdX0ug2kFCVmNBpsWLE7JSpMADJkWPPEFz0b96GdCq
M9kf9ITjFnIgxL6Ee4IKiVHFjqJVRP1FYmxo2BuQxo/2Uz6UhtyR7gq9bQnJKAtU
SLqe8AiGaODmCt5G8bIJ9E9yFmADgfAO3/+qdjaM1XIYYjySB7o5wB1yMHxRJGd8
uCbPG28PQL9BqDXma+7s2Z1Q8lg51C03VXzLWlK3CgYMqX+nG8NWnhAiC5pjubLW
Bo66fmmYjvCRaQ4NNEnM0c2LRFYcI6wB0GRiqYrHhuj6mf+J+E9UJMyzUQdzWlUY
EmjopJwImE57KW2lw1xtGMn3C5z9UOILQk0+oLmLqpfKN11kWMmFu9YhA75fbIhS
F4j59GsMbc+ijyQKfz9eCf1e55pmuX1R041+x7tQwVqnVT+oJwSFnx+QllHUYA/C
ENy9X/V8eAw1f42dyJJO7U6ZsO6SzMNemG2uNp5WuarUfG22Bom5/+lvjFQiqDxD
8PO27x1XNWUjOiHld9fjR3v7274iIAgaXkoOurLjX6DjZBBFBnZ/+wMxQqAEZzuS
zBi6dPt15lRhZ70wxjVbFxsuK+GgWp07+zin6tDzVy8Sep9VdTjnIlIO+dGwpg0i
YHsb9lHYgU93hEHZLavjUa5zjj5XLThxZiyHE3q1DDMv8E+HceEfOIP7v2CDykuD
NivA7TCrgWk5W8y/R96QTFbojWbMU0oisKKogf3XqYj8R/z5YTaLYtB+kV0Eh26E
g2g5ilmfmGdz3gxkT37/yLL25WHFHNX+pp0LB0cYS77PyuvR7MUwESaEjPY6NpL0
YHexlU5ij9g48OjU18mmRF9PX66zithQYQc1/mdAnFrITJ1q/8zwwp1he3cufqYB
ZDhxUgM7xVTYcOJPir1WP1vqia1UFbJTiZD+OhihKjOtr5Qidw29vNGee/4hghnz
E31pECuARo736IOjPqDiSYPc79nXi1eBeZ+G1oJX3R9jtZTap1tTT9z3GeWHfWHN
t8wZZbhbZMtiEk169bFX0toAdmMFEt9WbXjwFHlGhdFjzQ7dIP8IFXQkQEaeLpUR
GJyIkNvPsZKmSyxOVprevpqmfp9CTOPK78Xr3ULAZh6BxhTq83NgwcOeluI6BuL7
ZNzb+h10CrgRQ/xRv6UsKPi+kBZe5qSJb2xAS9T0UPYFtTLp7y4dqQcUeC/2OTdk
OmBF7rI19pO0Ls62AXb9cwWZBpk064821n8oAs9mCNnbo8wCjtw5yu81kXKagKp+
H5mgnMTtQRyGiJabJuPLkKiUxyZYQtCPQuizE01NZNPkgwtUskrZK3OHHviYFOBo
tPjQSAJN97IAzY5+x/AtI5mQytc85IiuSK2u1Yjl6s4xPGaWoBIZPeLyTP4nb0yD
ncSa6EUBGOrU373XxyjCGBTPvTl5ZaKocOsz+/j4Ly/jvqOifjgOFCx1mc6HWi7k
vU9zuqykyXaxnCLPuPnip04zXT3Frx4Y4p47ds6jPJhv/BjICiZ0eYJWsNo+QCyo
KNgDWxXp3a8DAQPGP0ict7tO5sVBKrqP8dvSIjv/G5i8Tqjggtq4X9q+97Qy/6im
mCl8EBlS3KAENpD1jI5cSpvkcsXXL2ZE+hAuxS43rWNqzIMz9KnetIJhzU51h/Yn
4Ox2AHWz/ngEKYwH8b1KkhzdcDvLgT5kaBFpAZbt0nCSttPkXoEi+UNTEAkDpwDq
rphhLDHz3QGIHS13oWURuzf9SDubWy9EY76huU8zxu57dDTdDHHChathiHMHshBa
rrTAhB6cgnqBYW8tKKYWQyfKteE7jXuGdsRQSwU/zqtbUtx2KntfGOI4fsUCiHPZ
LPFMNxwClXvV8bNbtMaO6TBUsDioB5uNptApIoMttON02m80nlHhO6werQUR/1TY
1nP5f8UcKtXwcyyrnfgvnbLweOEQplu2+ed1Fs3pSYnUbQooTwn0GzOj69whWitl
Q1y/Bl7EEJ0DH2iaOH1njf1aypfhL4cxbtzBW+S8LgEJ91wfoMXqUA2xlFJTCjjM
jV4QLf9n4cnZxndVZGOq4PSSHDHjhjy3m5Ps53LXaSixmaWo7BoZOsEUWspMRKiF
eM1BxXwvT75fNdy0mu3uOOBTTyhHv+iPmg9TY+HE5McStt5TAT0VG7vzISUhiSkR
UjPA801eYVGkS909dPWbtLoS7O09hYR5o3evXY2r/my+45rDi7MeoAHY5kndX4LB
OKdxJDjV9rQjEL6H2Lf/xQpkeLCOBkIVMPWpFTLgPaYdpNDgvq0BAoReYtrzmWs7
X0615VyfOnmDApfEE3ZKNDzSDru2JmSPPu2y8iL12EJf4Tb2sseAbTi1OghGotBo
Kxj+DI5gJZcLNK58c12SdXKu/H1YGMm3J1dLNEuJQufiwOyIMwozIRxYHMUmxAHJ
pW++1QoqEIQyg+jDR+KwtFg7LKeI5kNgs4FgFGp9dTlADmNAeaX/fjS1h2OCrPWT
HySQ0iyeNLrKTa4V4VwIm0lK2XayQrRJKhIXO+3MCE5ueH/ZOHG6JoDXJhrjM5xS
29KqZQEzV7zRcpgLIVE+26Wb6Ob/zrA/NkqrzmenikEPdNGa4HeRENVezbOfSH8g
WWAjRdmnoApu7Y+cztaltge/jpt197y3r9Q9cEpr059stiBj38WG9Wgn25BGdYQJ
EpsXpbDlGUrXlLTi5F9ft62rG3fBJdJ5TK7NJ7nOODfPvkwkTq8xHKTgP4kL9jkS
ML56DcZGWp4hspqgZ9OZATuElIsvU/hNjzWvwIbWfcPayGzKakKC/mj/1XnNZJ2p
R3aC/HDR7nBzfsQw4fqwn/NrvmfqNQCGgbAxSUUamT3vNE5IZfi3V32N5SuugZre
zzcSZxW8HsTFXiuxXBHGawLo6uX6krF7nlni24fgGtWLhpoiOw9IqtJJezkLQTBe
nCoFMQWEl+LTdzT5smRluEpWhaVw2lqfgY3C0g017mSJ+PkH/n6cxbOPJ90W5hbw
HP1Ujw4LjYwvMFZUUWzwzYXT4m7fffpTML97hsLNf+wnWv+L7NkIQrJHDL/wHWaj
2XxVtx70bvhdoOalGlYSI78MvpzJ8ooUJGtgelB4QHrjkKVt8rIMWDAi+64lFf36
uzEOO9lak/iZjlTZ/w0DR577ivMD2s5kqX73GXGZzBOBo3ph+tGTWWRLo5veWdP/
cKHeD932nXowB9CvA9+K4hWKhh3wWUocmQybxwUmT8DCzyzTrbTpwFeDLRYJNfq1
YsmrF/fDGSOl3NEJDN245wei5nZ3Z9AcPkV8QEqyJHBmVoGdtKbyR5QX3KmagsGE
juYLiEoYwxKyngr3jegNG9GbEtAPLpq1B2U9exERhrOopZPBJt7MaNJCCHkY8od1
j+f5CvhOEyo7G6Eb0p3H+enI9jUOXhh6r0zbPYl/aoD56vvo0clLOhk+TdQUQjmg
vikdQjlNjr9BQG8V3LMfU+AYYhbl1QuoJoS1tAQwQudQ7Mt49XQuyiKmUYby339O
kpOBKShBjaymc8UIW40lsLUjpLiml58SabTPCQNKPvsNXrAQ8Xf+cxo4Bgk4+raR
kq4zdgq/qWA6AF6nM6AmmEdYJ2eCPxmRwTuUSLJqHZKvZEX06lcSp9VvdPMYz8FT
itSrxxVu1y7MYK9PqqCN5mc7jwOhVAW0H3zwF1Q6H2a3S6H4iWFmF63xeZGORFEX
IlmdJwuEiom3ImPS1UpHgVU4o3OBaGXcLIEV3uQYPhFYDeNXiLi2by2hQZO1Uy/9
QfE/cdZkzoBY+7MbuuR914i8H8jrYQVfwimnxa2wfh5TkE50aHZwAAGk6cucVor6
uPMCadgkOscQm29G/1ZNzoJLfjTGt7o/rkXLctEbMHywBhrM/vdCP+M7+Dzg11mv
1b8jK0kkYZz31Jpo1k4MRgTtCqOYJPIxeJIRY9faxc59wj3WizSSK3FPCjzJfz9R
XuOTrprClOAg4ZiSEIUek22MOLt06YLjcnyNWBEjwxXKX9lDaSRGczrsHcspK626
zNQHmI56ENHCguxCBt9utZHgWNZ8mb5NoeUWi7K5izEUMZba6eeuXvF6J5UGxkH3
U1y8klYwR828lXxc3Isyw7Oav9KnnoExsraehsqLk/bdt3ZsEu4e00y1Zl2ckiPD
rHlyflslz9PDCM06wN5ijqilFaohdWlkA5DCBykxmI4PdAa341u5vPd3UNuDjvPd
GtzMHpV9WLmtP0tdN6WBe34Enu65niRpiPdKxfV/YK7w9i503SrrHucdKckqj5OH
BnVvb//Q1260QKd6ZGs+dzA6iiHBn4dakqXlPSoQDVIQ7EeqJcTWTtKiPAtqlTNb
zLKQdiuZsW0ll2VlKjFWSbVJQLpfHPcx+mfC6qYNTNmO/r4s1jhizHCmQCqTgHp+
TDDIS/RszyWa9Fx1QGvoxktPT2oFfkxuv09otGstyecyleJkL6giDAiCOYePEior
UDNFsNWs2DiHjNCdQwcVvZ2oacdhDf0BAW9v7iViMdLHg9rOhM8kby9CWolBqTrB
w4yKxRXsqZQ1rF6i9SFADzjPd7UlE7inSZvhnkjBg636hu+azax17VG2hRh544ry
AV4cBibByiNCxHFZVPGvNZXESw3rT1Q1mquzdmi3gRbVGtRPUCoFoLalq50mLP9k
0Sz+NEEZAm6+b7MHHV2DiQXbLLOTTDEjEa6hcTn2gxFll/bTIg+GoR8ZUk8wZ33O
go96i43yHcgO7ISTEhoJakqc1E0D2pBl2cG5zya8YwgFwQ0FbO24uzP7hGRWJOnM
g0HzLNYJdQPDkZ8ARtZ/z0uAeiA3AHXy6AePTZG0Vm5IaPQWPAyXpJ0MoJmPhG1l
2WYxhNCVA2WJjVxhavN+O3V51+/JMMBZOMf8+22/DDpv1W42i6ciFkbOKdXU8Ebd
g1HPoM7DuYZlWALbu+42QYdwOwCdTjOercldBmShko6pytsGpGF2ilJAuexARV7F
PPllE83CoThf0LK5mxlyE1xmPdCOj4WEdRRqFac6qsO7/It4ktHsfiiovsXkmuFU
VipSS2Tb5v6Wj0dbNcXgd7/hi4OJFaeKiAZWZTVU298Z22tH3SoNvI65cYnTTgb+
qqDbrC5lkrG3gT/RjOkbDcHAxwtQRpCJBeg6O8buXsg4kc3Om4H2eth2B0eqwFqb
GemvCqzzYN/HfiLwkKPqoHsDs1jH7Thk8n9HvwhUsA4mQXNGQ03lFI03mjxOtyKM
71LWRIa10Fe1jIOJEA7wnEB2RuMtv4ILkzgLYOGjmcfME4QDOY5uKPyxVfcTzcn0
s8EETgrqN2kYEwHFDTMlXEGQ84HrYZqUJRzQ7AI8Hq12X54PquBhnwt6pLM7O+8Q
RgJKmGqYrrN+RJ1njwZy47//ZKFtilRsb/VFfIaid7d+pCRboi1EgsrXRn5ISAb+
GB90NjK25hNhYFdEDtL4tEkx40UHdez8I1wpgZSxQX8g6Gkqh7yOmxU6nkAxkxET
oY+hqZ3/iC12CN2R3JkAa/DSiHEYZjAZEGUpsdWAT0R29gM7YP/Rtn1fy9GVZhdL
h2fY0gEcCufncTy4HknOzVYwTVlvOhAOTv0l5LmIkM8kt+8qofsMgyDMqsw/P2B7
f6SQSZBRUenmrJ0OWDAgfGbyPYdTyv6q29pcxCbhnLLtfXEpDvNPKcYi/EGl+cgM
DN4F3b9W7txLeaKl2RQrBi4hK87wYhkpvh7L8wokClbJ1XrflFGaPYNp0PIgqN8g
tfWaI6e7xyn26oP1QCQMc7uosGWhxMegrv8G/SDBKCRmlbOfuE5A71SKkDfrrbM9
CpyUw2hzJ0yatRONuwr18aAJF9IrJ2QUzwwrx+7Gm/zHgXsapoPFACu07mVpXNb6
LSpNnJkJ949wyEzg0ofTm/Co2+4SfiJrerslfmurPSYAyIDY93qjOsgnXrDJf6qS
29oygva8myOFcDUpFc7qQxYd2qTwljKgFD0pW+e0PDoITzyCHg5YNGSRnEaD1FtG
BrXsRApILLjCICOaJdr6Qds0Y53tr1xj2rQ3kex6fWr2zP93wdxztB7iU6vGVWcE
q8/GUHeXT7yCYDaERgm7TPREHsjt+69+ba4LUXT4wGMJyj03/PV8nFLaBhNix1w/
djQQ98W8c/omRHgKqJfOa0tw99RTv5dlP1isF1hjXY0jC2qjsaUy7i4MURXFs8MV
JXzJj9G+9KBEIpOm415yDmM0X8oYogNMtYp5UF9QUV7uBB0KbQfEDEQaJZ+OW1H6
e+nHNPuKCnMPKY57sE8F/QAdO4MRa+aQGS2HMuLVk+ZOaZ3Inv+psFebZxbFxIzD
/zP5YqPWGXToqHyTf3EhIIHFQ7XitpTx/OtJ++HNSXevI7vmjJS4abHY04r/3hNg
FsxNnfgbFD7BnExZaZsusVQissUUf7BUcLoMgZsOx7xRxi5WbrKSyyGvtDcxUwwc
o9WF3ZbKZrpS6vfldGfiFwA3HNYo+A06dObUNrtwBJg0bsggPkQBcU+JDPHYgl1a
Few1Llg3Aukr9UI9KBOA2jAy20XUZKTE9i3Crp1rJKAle2Q4u9XOxQgUa0Ett7vU
HYo0mLOPjw2Ob9gSBzjTHfj/eVRXMFTD3hrbtVdQRfwny6Ew3dWdQR+jblUvfXPd
ZZVxWQDldpwL31YPJrLokfaNBLfN0gdtAayr0CaqjJVf1wivnAhJL7aaxh2UP2cW
IErQxFVG8o1IlN/g4GKMCGfIM7+wvfCKeiKFxzXIBLEwuIGQaeNihWG8LMxsUdZA
a6fdLe0h+JiXL8LX87KK2lG7SSILp7FtTVjQkX71luTvBjiVJzSvdnAv0UcavFUL
EraxVEQ26Q1MKFZc/hQGGpghAzwrh7mXO5k/v+stBLuDGxiTEZEwGEK9scevdLnR
51xDdiNH0cbtcUcUMPSH2Pyrr9ScTf6TcV7BSSdZ1xTU2mqaSzQGLDx3v44QmABZ
Mnpivg8hxIs2dScgoRmtEOQ288O0uJ1se9yCULXISbIjh+kilXEpDbzkYVoW1MHq
1ZlCm0TlbhxuTj3iLIZx5gN8K0nFyv8Ho21N0/LUhSKdLlmSa3L2n77k0DaMO09J
X9CnlcO4HK64+AYA9wzBfH7ZMusAeh/sXdktOzP0FGb2a4uO7WtFz9j4MTTz+pPu
GGkPYiBUrQWIgxIPYZoLFpBaX9EHXcYWViD84+stQbbg1YG6ia/b1SELkpuwA4He
jVK+O+7sSUyjyqf1eA61fseLJVNL5Y245BRYKEUs2k1q1SPOcczalOzSoc8ZzheW
b9BgcvcgJe+mfowP/+F7+jZ/iIXwat6xdVNKvS2FtVKn2yV5ukkGbGzwJFnzgybf
J2lOXRuGJhJOnNj4FSVZb7nvI2n7i2Gdh2uD0l7kAm8A6npRNay93OiSMZf/J/nP
ZX+JUTzi0s5kffyojDDBOT0wpEAZMrtQd4Iq8gvH/sg/qrYK4mFM1F/oaie+9rCJ
05actNmhmRrKNCKgJXh9IUucwbVKzt760b0izewoAS7W1EpOAoRIeeH3odsU3Y3Y
Y/JZ5v3GN/vZhrL6rl3crWm8Qx4vpcdUkF5AmNCGxkjhxw0IExNEdXM7fz8em6N6
U1ijzwKGlOwlhqGrgADN4lQekwCtpxRr/OabIjKhmtpolbJxvy4OIF7uN5/4cA3m
Az4nKtbm7EWi39R10VJC5bmGlTHIeGjcoJOteZnlSNCjhXiWskJavXQ1duQGlmkM
2mNGO2GWD+UMtQlDPwXn6MMXBXOmHgDT1KHwbqv2dz8W0yFqSCzNWyUjSYZqU0da
6JrjecBkT4NVoWVm9h0z6noIM4Mu6geZSSgV7yKp8dFq49WGLzAXa7/FAxFHNPo+
jhU0vcAtYEs+gKcWhcFf5hNvzn3d1+ih8yhOOadJwRT5HdltHLCGQlp2swwid5W1
+BWfNWojwSEiGRjEmKPqWEb4xoDn1IO+Lx+ilmZAJxzWJvHM5l18Ba86ZGIkGbws
iScUngcQKvx+QL3e5cGwGjdaWvYVdQo5SnKKSyCeRtfLqthi/eQQ/DTa9ZcK6vDK
Z/UtHm+JXnCthwpQ+/EZdkIBuYltKL1xEVYcg4ILjlAA/j7PVQTVTZMEyL496KA+
lCLjgW7hm/eYhwdqr41MGAHfAUmL/g4vH0hh8AZ1Dq214P/W7zYyfI7oai+ALn/K
zMw9Zwh1OJwplXc8ty8zC9rN0G9mFuBXtwF6oxfLBoq6Nn2SBuZjvP7UW1/LbVxB
b6EY/MjfRc5rimlCtj2TTbKY2WzONtrjuqRaD0XtIP2pP7dW/BHizy3gHAVAgTyl
nNFjY1Pw3In68WjD3vCeiarSGYMu2W65mdWXn2TEH8s14G0t/2ZlmBPpyhGJMkZk
RZKsFWivbLnkvg7ImrF46bVWThoYmeLEaftiEIjm7UxB+W/GsBHLHxRozh6WyBe7
5MpnNjvxhTtQUfQER6v5tZa4D/1ERKmthIZeu1fnMXQ0GGFDMEynxabuz487ROa9
PE8d2VLZq35zs9QFCMu7vatFfCNEUaeoN2gNvAzeMmYWVn6zM/wx1Ko8xyis41Wz
Bw26nROwFrdt8WYFfRq2pQ1dI/3feCMNWYlBpeurLgxqij0zPQeijfPZLaN2qywl
oxw4xFavr9xeoG9Y5iyTazqYHVK/wEc0up6iZ4S1OTGbuRRtu5s5Gl+vcuPnX22I
ggY7pO8av+3O3TtqdUVMMkTYKE0EksSeB6tHp+9TkkFdLSWJR73Sy9aWxH0kM4SA
bNVGKDkAdNJSucyVuNWnwz8ytl0TIH2IffG6YSnw50ZTV+f3QyYgNMu+1PIi3dwR
1o1h9XCRbo5o+G6oLNY5ZvlHz9VeJrLnVGjhjRrdPlAi0ZoQu/jhGI9XwNSOKs8B
reDv3BCj4FdwPEQOTD4c/ms5BYNqYN34E9/vipbwiERYGBLulh2FwRhxj94kGOwI
ghtBUmZXTwvf00PNfEPEhopD2AWI2J+banr/f64xDWs7utOmliVAGGqueRuShqgs
Endn9UcQssKTjuiCbDk0aMsi/qh9SW3VKvzAxc2uajGA1jCBUgRT2wsxDLlCZgbQ
EHfOzgYkNupWKt8K3owtgMOoX7nGNJvk+XOfiRa6x9YCeb136cCz/0Shn3zV/gIC
KrSp+vL1WYGgKzYSGoyIYwr/9zbPR4hb1jRqnThNIT7qihDERZx51nOF3wxYWob1
nIq5VjEA382IMjRv7Q3+Pl8omClyYO3eK5jbMo7t/VvhTXs0vTxhhrOL3polV6jv
GURboMdxNnQ3k2wsxR9dsV4Cm/V7PX8dni9K2SWA1Z0M9F6DITJxuORA6V/BOJKv
lkxSxDw28uZnZjqn4UKIJXRoPX49qDozd+w+4hAN/iAVZhKHXiESVpSq5q06VCCx
rbGbCC+OSOs1DgphNMReAFwnSHmNsUs8clIQoff24PGfGqV+XqJJYH5qOW+n60FA
ziF64YB50iZNqTJDQ8EPZnlG/T660YiBuPS86el5Z34VrfnJUXAIy/gZ609cGZNd
30RODF64p0VDKA3bN37lT0/SItxeFrNUstoeaXNM6+NQuBl7G+7KztXelezFWo6c
aprYwvaGsp+frA15WNzCMQ3gFiZCkle43btIJQE4rFo3RyqXzMVvpzPIUls94cy1
8NClTLrR2wtFvm/8z91gFpTp8UloIC96q1w+9VJuoEsC7f6aEuXPQQ3HQKkL25a6
iZR5YtdF3qiIXkR8/rTcP8wnUikz/3i+xPN8CcSscpSKpCKFNmgKG7Htj58Vh2qG
o5BKqV9yG261ZpEStX8RyR2v6Lbd+L2p4f3wRUfJUfuRoAxOcqVQTqOfBlZyadz5
rKt/AtLTlI3JBLbgjeT6U/LRHTaXBxGm6qPs/Zo7H6xpSBG3AUve9F6cZf07FUm1
hd1MFyWslZu/x9T8B5Zeyz6Z3S/SE+XQwraLN9JN+ZH+Ec3aAwH3/VgbdS38/nsC
DaJ+bceu6tL1weBCDWk3LF18ywr16dlATPSeEBPqh2k0/i2BEJXE3bLVpSdMfU9o
jwr7oZt9kMnLKwPMtZWUmLfpc6ylKuqemVPvtWyLrw3RGhk/khlD115cVWmcFn7l
oGudvHkwueB86mgz6W39rc2X10ZtM+6j9Rk/Oa1xp3A5wS3DhDi8GlAc/S45gKBf
sbabmOY1Zo0V7Vg+YPcyy2cHrlrwQGCRjf3ujMbqketdBGf4mVWjtD9tUp5LY1nj
LLWb8SUpg1YvXHdw+lJbNcHaPsmmgZlUydk+ckfdY6lqUFpp26stl9N/AjV3vKwp
5qF6sq7MwoNT2oPmuYKo0Z+5+2zNjW+w+3ESJZEk6w3eVCADRTCKnBYmYuGG0r8T
/wKrf1obqS/HwPD1VH8RTPSXr+ugli3CQrjmvMIPjPlnmcS/neV/TCnfuHidqPlY
G2w5QFN96lZm0A014ya/XCX3ad+fiPB/xpX2J9Qf7W9uoYhEoWIHAi96x1uzXCp1
8CzM0rP5zVTrsMJOsJCLyks5TOTMe9PouAT9wFc16ZU/5/gT932chE3iMyYptzoc
BpsR3SvFbZ0Vuf9o7/NR493F25CrdRHEB4mRsfYxSEoJcjOLHdrEenWYrJB2IJAO
k+0rfGRsICcWL/0jNAAmzwItVGmDNpFfBFiU3TGXCDCIy2Z3/y+IE7VumbPNZpa7
Hezhg/0djFFyTPwjzlp2dThBOXMrIbePnnAji5a8egXCwUpkZR4xcag/MKT1SFhW
NeqR8rv/RFgJVhsB+XKNnq3mHY1ZQ1w9v81wiM+qMQPL/RxpiBoq767+zub3Uzox
q8q8hvHUtUEYJnLRT7IpCKJSHhG1nJB2aRzBZb2jhA2XEggNx3u0hYz6MvHGdyPj
bfAd10y7M3PzKlA4amhAetuaga4ODqJgSjFWPrSEzva8AtBs0RQmXIPPHWAlVIvs
/WeROCXXmajCxhmN/+/qDz20SHPhsrwk27P78fD8/pIMUBb4hr9pCLMAY0Y7LOaP
CPSS7cUQPqUgVg2TKPK9Maxq+gMoUeThMDuPt+DY6O+8XhThkEZWCTiwf+Q++M3r
rIWPst8WGxBk3u+Whw1ECYbi4KBCxC1YWBDhtTf+oeQOz5InCbYnuDgoYu18v9Ua
B9TElLAt/MkcJJ3SPe8ocbCYf+KeZiDj1a1hPt9KM+I0PbV97utZ/HpiUwnQHq9V
x7cIGtQUtGAPY+COAL0Ip36RvCFJBJQrKy6uMiufeFBD+oI5tyCen3ulT9i9YNcs
FBuSriDmvo4YBWSxzUmk2+Yqv1VhlA2vFXAbHSSqDXml8jhyaUa/bkWVG9laCupH
GcjNi5shnYZlL/7U5GL9U0MRU6YZPRTK6GEKg30j5FUXqflhLEXpfEHT7XmpXwtU
4oVZdfvrq6K5pTLAnrDr/aYye3QaKaObrOVv0aq4UOetO+eS+Ux/dNZieFzf2w51
qo0cgVeAkIxXK/ufHnOa/btaIE/qTUEuQC+oNxBQIQLffhUJabeF898fkHEtMHiB
Z6WBOHP7II0NPNse7gouTCUymJISZ9H5qeL955JkTpLMp9ifQsRSAyIzvdTSCAli
hhO8WmCU7+qL3AZ6qd4BYslL4au6w6VxscrzpKppIFUaQ9+GTl4k2XSAnW5QxTJJ
Fiofv1pWewCi2MLYJVCejS2g+6WSvz85cbqB3JimsmiAVsmVhYlNAyUTTB3pLkPK
Ako0TA3HT4eWBLosXMkGC9vA6GBZQVexEJ4h0An65gmYLTeYxitVaOXnvlnxgE3x
mZvGF8Q3/b4bdqE9Vjhznmb7TSrMiG2Td1F2dVwFrFIK+BnRtQqqAgNGk7rxd5cm
h7Fwb4vAsfSgqEGjAYwkiIslt+AXHrg7Fr2/wUo9HqxiqllxU776B7W5rqPYnZ0B
08nztov/UqTCbleq6Fz2s0EEjiQgB5qFWstsLCWSM/okoRJNaxTRBwBE/jDzUZQy
YAF4RJ8OOGn/KtXqpHpte1VHagAU+INd0crE0FHOUcHzmFPyY+uWC0x/rJDoTcpO
+PZW1jZoaOzn1odSc9rgsUS9h2TY66vJkm6H78SpnWYFkqlLLs610ifvJhu/zg/3
rzZna0k2RLQHh9aNf4/HRLKvqPZPwdwtQF/t0wMeVjKf7gJyAV35yyEQMvoIg6vS
jeMtDKqBGPomyCNx34UKfHwQB0SHWD0QB1SLUcfIkiIJqgiQxA9gvsZYQveWA+Ge
LlNvuHTBUhTA79UnnTQXe03vYMB0GzuE1tyOGQjIYGc0VnE/6x7MG2d5j646muiK
eBO7f3pTDTd/qXaAtJUCWEJae/lNSFSBPwTkyZiUTUTWxxDLEAlruEEpj8BaOqp3
+C+fBmEeEkkeT8Ce6ZcjHN8E9kk+HU0YI+hbp0qnpFd9WyBTMzMuWqITuiUylX3e
N00gWW64ieXvc6h3iSZO6AZFD8Ir2FZrXrsQINXkvEVhFhpwCc8rR6redtNtRPXR
DiOfkt+ieFtWjkv6rYxgNjbKh5OLnMBoDUmGPUrYGfon+AeMvpYNyHAGEHtW4pe8
OXgUCKz76YZVyFMOdr5JlDytnb28eFhp7jTWtLiFNZtZsShB/l1EiYIcuffGLdnK
yuVVXxDvHx7gB9VVeOo6r3OxUDFoMWvMCYZQmUqF3zBaBS/cXDEmM/N1QNX3rKBZ
Bb2lXs/K0yz2d3D2PsaY0mmGWaoP48dddx2zleIDOo1GdVCP20Sdyr8fUjKn/Ztt
bSiBGBuJuGKlHDm7+nyro90UsDEQH5mYrzjDaclDNbIWsnPsVu2zj3xhKkNFWoVz
q4MD4Um24YA9jxq+VOYAIyG6++cwf8n3H0jtMYgLPM0MZLbuKKFkFV/q6RVLlu27
42+GY7jTsKYB13w9nU7bPdD/4qGneL8nhFffuct5/GWxTex+P4w2xbMRqq0W8U/v
WRp0J/F53aGAHKtOPN8CcupHQtBOVvVH6onTaVgHWhAI3wFp8WsPwtBCeV3UvaS3
wRz9qsO5WdjF2HvDVHWW90mfF4vitApGwbwmdJId1T/XaoGTgh0AfyG/txnIm86i
J90d9XMFSTlOztDXtS6+lrag41fb1ZAfCj9sQqcCSASV4Sv29Hqp1QB4muyRG7eV
g4T0OqhKIUOLctWJDLQY9JOhbnUyaQ8SZ6uDWRIW1QTiYMOGRtrRADRpDh5C/zkc
pSXs2cDjjXvRH5x5jE5vcOmQCBQd5Gt26zCfX4wmGLzPHdB5UillJG7rC/hmZe9m
kElHG2YJLxADqdA/YyL1WLJP/tHeBdbwJujP+SWq3twCALyDfiEjuBSP2KemA6bE
aM+AZfxDLh2qwtNdRwVcQ1d/qA8J8jDopKjwDSDd18VnkBafwbaRP+a8KjV053cn
Oo8feTIu2YheqgDBSQ5waEeU8IggAR/No48bKC5qnvefcnWhoQB8+GJeIb31nbmu
a7Yp0oVRksHo1NhQye76hVMLIf5Y/QodFTWIG39uatHyNUnfw5LDko7D+2r1WYx/
8k5JBsWdjmcl8BtqEYu1XokQ1C+xgKmiE+mgkmo/+j0n9+C4gjF2QKQrkowVYSDK
azGF0Qv9nv/xVcWx+1+eUVcJMBk3z89Ibx2CHNltj/FYuCZeZFeIel5JZGYEk+8V
IKlzmnTaQX+ICFEiAjUxE1sGPq3qoshXxljQ3Ro22SoTADdYMjGPbRPpjehPNXo4
RWZBxI34vhtTOpz+d99Fw/wvEH0IkwxO3ZhgYz6GgJnPYGn8rDg9Pl0bpZUpkPu2
W7qozS4PiAWnx6TQ8BzL/Xqp5P9beXTqHaShNFamVJDVjSN8XzEc9umk+xUVow+8
b4w0I/NmSYaRaKpoLkaYIAEIIEMYt4FK0fCbAh0zkTo7qe+VQ2QEZxcA7XB/xcLe
t/bn2MxTnkZNB2xdJYbsFM5j3KKb7iZFLmD/qV+16FxQIobbgJL6R6FsWutEDn1L
CjrCCJKZSWFcTvxH+61JhfSD0IeNmUH3sMlbnTXB5dF0VKG7vUyj8xMMowWiUETN
6xMv7M7gxbS4Uy8+QUdYCEUsV22yExyb17sNTQr6NL1LeRzh20Ckk7lHDHvHFJ+P
lOUA7QnBnByJyDFe2oNDkB5EwFVf6siAcoXtxn8sY2mC8VjS/H9/ByPvahq4dY7i
yp1UNbXMSUKNdckbCcnwQmWf82ectn2FlX2chc+iP/7iKyXGKgVA+XjpO5WlD7hL
Ng9dEYozba+odD4snLClA6u+d7s+Z/g/nLD/ECSAqE2BSkGA8Ahujjd4VAsxjth8
8iJc2UQjDVcUywXdNAMdwXUleuA1Xu4nF9r+pZiKLq2j75umeoQ3JSTepCrL7eQe
SuPt4t1nrTIsP+cpfelPwmjwjiiJazS6avYWWSOphx48vD3ZHTL2OTZ0jwEBN4wL
eO2W2dmLNAx5jN4Zvyx9lpkFHQ45qCcMayoSLjeJmFzrhcZUxxdkTGJ6USGuDmxM
PfO3i5FlVvQRx5o4jQY8bI0WsceSEx2lSQoGUlzorgn6/3tB4tK/3y9khh2c/3rd
9x4AIsy/DwVt73EHeTZnMzk4cZOaoKet8PVwPmv1HEbzygKwsjOaq2F02yeZsNHY
pItHiMZx8g3CErAR5oRJLhYR8rTIfSBd477xvwCcOjbLaRXT1c0wD0CfIpKOSptw
BQgW/5TaZsMPC4yYjGpzarmK/kCPn42CdommKCRHI0PCLWro3X7ZI1o9QU5SyYpY
TedvOI281STnd/DGIP6jdhMqXNo48sO0HDEUECnbkmULq1Yrf5KjU1aRMbIkHsxk
jFJffGPMkcatkivmRzmJIc5+HhXKjw8Ylf+V9AZ3WAaag4XRejFb31gtsQ/Jv0+p
XXpcWytdo04ngAhQQGGlanOYdp4h31XHyejpKmpJjjTUcYG/Jj1Uutc9wRsGfujB
fYv78MGIKs8geaabi6xsdCQc2oCJ5K8Yvv/exUP7rgP7V8HbCC/FR3xoz+wmntpi
V43oQu6JAOa08b94wFPnnC7oBul3n4cA7UhaYjYv/uV/QrqfZhTLlTq+eqges16L
yOu9i6GUUEv9+XwrX809MzV+GAM5/G2w/DL51X+GoRnuVoeCGaoqAZd6cJhX2NH5
0u+btem3v1KHUthyC5jX5PD3AVAqGbPzCAe+84DoLlTxCr52/BHvBRNBHlHn2F79
f8Xq4fZ4KFclhuLWeQcp5albGcutD4XPHHdG/HeFuw6F1KpNwepocF41uykqvRfj
2+b8Z4X17EHeizlEp/idTmRHXQ0InL4kuqdcSFFHLMKWT3G+LfL24uQVcs9UgcWz
914gsXRcJ17xoPnbEXpvniXd0HvbZ4nbmL/xyPoSmv+GlsTL9if4pSrknkDANVnq
c9izUjJs/B/Y5m+X5znu46t8RrTRfK0v3QUYBvhSpIBv56symQDQ4AFNDDHgdYXK
dh3PTA515QzBamDG+iPEE46uh+AjkIho2gN5wZOMcl0o7ygCYWV0b72jbbQwRGxt
Et6zJa0eYJ3QhDCbahXgUkY0qT21HO7ZN+UTE7QOORUNAVrS5VXsmqo/Xul8xco7
vGPd2lvx3/snzvTMIUHu4q7snZLuX+zXbDYsLOhD3eO4OfPR+M1VKkfG862N2NNw
Q3sjbwdTOW+2HM0XyuiewDC0yEr6hEdf8d0EVhjDGNM/u3OxNehFim4gU5IERvGu
DYHg2YyBRSvVstxrna4yKShU+8H8b/dPxW9OmdC9tQS8OtoMTKIspy4vBwUbBBlN
eeZSdccD+hCOCr3fSl4+7JKmagWKD9vtaC/xC6Q+UuQvj3/8SM4/b1fV7Qvol/+v
yVFDOM0YTDyNl57zFqkdsq4reE094cEkS3S7FUkZCpFqXjMNLDspHv3A5lCKTe1S
N+xe2GEjR/gRnhHV0ZP3e/GyCWKB+XMSJ6uzzW9NSKi8MNja/pLO0RB3R/Lo5T29
x1qYSj9an09QG6DgLDG3G/MH0O6vk20Q2dgFz+foFVyxGr4he6LHG37ffCtIeyIs
cZOj0adJpYZY0fRZ+mMRpV1Y0U7ixGlvTxwPXTn/dASI8crumRKpx91+a/n2STOB
G66Or+X4cZ20ft6kaN3+anVgT3x9itYq70xtxq6S436Vw7Yie4ILZKS+R1U5tKcL
eZYPeYNdJAwFJ+0i4iv7TD1IgqqQcxyMkd1MJZ/ifx9PAckwIrXALc+A4/Vj3LY9
71iGfiGFAFgqFUa89gXj7gm2Nz58+6NbQ2XqyM56d/KATaa2mGp75Mtsvm/3w/Pw
5Y6v9+lQP3cF+2SXpp7vfAaM6z9q5CTt+2b+NDirMeBHIC6SRET16ySP7K4oJXtC
Tihzs7XKvhhMyw7h26wvlaE1oetSUsCY7qLk0AXuLv3vRx+YdeI+dxvQGjrQHgRB
Y82dvi5vz3GKxrDmiPaB2oOax3XifnPcXUYFei3Ms1NTniWip3UsI2AHQ+tBnIYD
QWvrHXGFjleq9jMO+/9Nof8MEzGj7K2MSb1ZWf4lDVq8BwiS0hpd7U23ea9fNm6o
1dpGMB6COtxRRVzFrwF8P8cUG4jGXvMFyk4u6E7bPBCiHLVjFIgYR56EpXXKeiO5
F1d4rsk4T9hZY4L4F0CC2EiWUcmOctdTME0x7HmzfdKzZYJC3XST60SFVxCkjc1q
TG7Yl48muZD+EmPZluiumfKOByR/myeAGDNtoKcEZEBb9PcPsUkzijiSH8Vtdj4c
YjxHsOFbMZRbNVT8Ge/YOt+9sx6y6aLvodB8MxyFjJH4gKg/vobPNBfcyUdYst9s
YB7rAT2ltumLnHpHXSI89eMnrMKsoxi8j7Wjn1yj0pg71MKLbQ61n44gB1GaRkcD
mr2f+lmky4R58BZqHfmx872WlSwcxyqg0IePXRpMI088zTzbDDkvhQPFxzwONYfQ
Ow0CBtSY4W9qRkI+j8QhrPz7379DANoPvPKFY2vNZapw06f72rk46DjvBVVZ0esv
tIar27MOFKSpKKKAzHmqXjxz92xifq+o2nQaQ8ezhMbRYUhKoAEDUTle2zsO4qfm
PoBhMm30sMFV/UkXd2OphKPdvUxhS8ZNzP28bNiA2JViSa1WmMRL7Y4gpIQx/4br
5dVyQxQmMvDoT+lUWvOsHhPTBysW/ipEE69YbxP5VwVXqo5xyMFJ0UW7A/ZVrUO2
+4EXdf963XiWdFoDOXvRvCk9bHssgqyiE2vs2S534nBjX87hVeikHDhr16S1/GFu
WjQNsXWt4VdWMHQRGmJyrv80dHVuVKSOC3JyuotBFiny2ShnqLN44ObJ4Sh2BlzH
+6fIpOhhx0I5WWhUJO+r4MqSsnDGshiBPTB42io2vJ1Cjfxr99zjwS4mY0DOr1q9
dnhCOEEtIaDLz8fg5gUlFRRLkhfNCBbn44EwmX2eOrNbzFRdr5CcUJyxhJ30vxaB
Ns9ErGZyft4q/t/WmnV6D/uuXzdpfQoZcKLOYyn1sdq3Up4aoWDeL/h4o5MXzs8+
66PoSLPTBS6bpPMoLKfCvQ65SRsHuvOTbUksuU9HQa/YmfOYiiCRvm9Px9i5QgJj
wnB83/ELspoKCaTs+2hm0zKh3pHlF7xCkTn0KQzvdZcOqbCmbGwA4yX26kqqoWOX
Mb3jJT/9vMDs7znWi3DrheEi0QicGwtjL2VQW4IOX3Z2KPsp9maafH2FRcYNQBJZ
Remsf0HFGqJoWLOen2Qo+xL3tPFe0fijlD7xPEh8pVOJuoGAtFm5QlTWV+nZS621
DW1BoxALxHGcaGfr2cLOy8zLp+QTMDBiXBo+9PuNcvjmAbx73rOTFZtAV0SKt79w
ey/GBLXlojvaye+EfDT2e3D1hAxgKh5yibcZpF4NT4eicc6LtbCYwAjv2ROTfWTi
03SLdsLTFuAMfNYW1/bQukOLERheFJJIKqQ7zJjkFtPnOTPV/ej1i+1oAgrsZo19
5QBgM3TDPkIoy6FxLJMfmBJZYumfFfLRYXgLEVlPGdaIZodw1Dp3uP4E0Qk8gy3a
vUjsnsho4LrYkEFBQBjErWWpaK6MTGxwR9+rDTQCpDVTF7xFhgJsxhBeeVfbUp37
5M8PcoNcIJaz2r+xYWtCIGIHPBLU7ncBKaqsyGdFoHMCj6Cywx34ym7kNP0hnZ+u
X5UyyryVkAl2aV1EawYFNIVXSpTPnH4xiWK1aup3MEcrCAHMWX3e0VF3tcvdQJwK
DbzHga5UxH719YtEt8iFcrN6MPxUejbTlbh7VTs5PSTf6OsbMVkXjmHBlj3uapPQ
u90jVvdvw2VrjGHArie/6dW2XIRroR8DajaN13JBT1yN3MKDbNeEGz6IJrGxl4ne
PDysiQjyy3F0LEJbtgOalRSjLK8NgUPHK8YdpTW9DKYBW08NQs1+fxkdyhk+s53Z
v9+ecGETO+G/fzVvkpJa/UpNYGktirncv3Kk5NSAgfoFCp/DFp7cGWeIK8C9kGPs
D3XwLnTFLQNFkjLPf+xN/xwJz6oiZJM9VU+cjoYZVZs3GaegLdUh2kGOHSUStdc/
lLxpzRQgzQpt17yYkBQuuJM//o3HbS5/cLMxCsS01NQu7Wt66TVYfDSjsus8s7ii
qArRgwEgnYQKzJFG9qhbWJHQoFuEeY3gyXrAysBEL8GjsfSTTP82OsDLpMlqCplj
ADYrEF6oDFfC12lFjuFiIgx25FfvHxUKeaSxoEcsYYuGULw115CL/uJyRw2WK8os
uAed0cbwN0cACSDmDneuPzWkjWZ9jnCROiwNV6lvBv76xgE1Mh0kwSHjBVHMP1go
IvXhuMONxC8t308fqdgkQq0diZQzrX7yx07Ubo+JtS8bLdvO2E2wSSlPOXQH5waO
wVRrj0GPgHeB4sMTppPC7VRUrCpoDIt7uqWNbRD7pyd9hNZbOO0Cn5jJ9jW6jamR
KPYLo+xLb3mnc6S//4xZJEKhilbHOg6vqQslLaa+4yFIuxs6383gi+fAqZAMT+4+
1Oe+sK5S+j8V5Vo3jFPnXaDCfC/qhJlZ5V3zIP7Il8n/gkISusla8AhRZ3IKEmtx
8w/JZnP4i5wh2/lSQ2cpnzK93+AHFOMQNhO9uRl5/o0jyclXisG61HkbMN+OISF9
CKBvUePaT9BWqapCSdSbT1WOoQaq1/DaA3KG58IYgftNdynxdNT8L3I400OTESLK
/PgOCf1eOfjrZO2KRat+txh6BiRVwT0UEXaRqcz9TyhgKS9Vv+WF64nIKhOAftLk
nmkHqdJo6k37E9GHo0XHurgtr/zUzlDOW8HrR09c7SHeUtlKhYIjvUwEW5xVfS0a
WtXMR8+IbrnL8HiINUiOvyPihxxqsTYeZigALg0RDwMeViKqTfFd4RHEAfNlvRpZ
cTnlHXD/OIwLdUk5afN8HWwTuUJ32l2LhFeTH4SMbA9N16KvtZkl7ON7mv8Weudh
32MA/DZK6qS43WYvjygyu6SlvqKnnI55oJ5VKX7ncz/OwbQn9qMbxiUSqq8MxMoM
gU3mjK6QD6gm0wjEgQTEyuaF4MFzWvq66ZBqQojagvW+vYO5IDLpy2amd7erw6eI
tz5DczWxpP/w69kyTi3RycjG57dsgFeFIlbZ2R7y4qoSq3wVA8jqZBZKAIyV7A5S
Q7/wdGorM9wPKarxb1o0xzR57WiLW4ZV+TEfH6L2XG0mkNR51sym67NdZWJLbigZ
gDNO3gQomakXTbdeyfO+VGhtuM8pn7j6bQV4eoH0+4KIFtbh8RyiTTB5EHt063XK
rPsnLfnp42bz/eSqHjmC7cxlD3P9VOBJahglN0D/U6Lb39Xmg9Tv3Hjuhxv9j+qR
vWvCoWlrhyYaU0eC3IaiD6pUzKIDSxvnUFSOXkH6a5nUo0noAy+WZVAsYcaEbaLH
TpLWGL2YkFdWXLUNw7Kt6AVGJC2En21OT5TYZfFsMcgxzNBxe9adxSZdDEagHAvw
F8KAOhrXPXEWLkOyu+XcaurcOabYm3DLghWWRnEvvF39hodwhhw3yzZzHj8wX59F
67muUfZJ+0Ns5t/XN669xb70eZcy1u42UpuHNc32maUB7dsaYCjxVoPSZyt6kGY0
FyGr9KQ+s8t+CUHXU1YNtNg7om5Iu5HepoNWO+PyyMDIPU/kAfnTXKT601atG75s
n0gnFcpA3FRFhcao7Bhod9GOoc2dB5X5TIdMA87cScRt6hxkiPDz6sKRfk7omsva
4QkhMVwzhw9dMnjTHicqZrIyckmXEjOc+VMWewPwp1uzalaLK5KBIcHCS4BlN8A8
d1jR6HimZfQDed9otEYkRXj9/Ks0NLbNYQRvDwQN13LLMkb6ANPvL65a2Mx+SB3+
6oujBjQEvFMTwPpxeunvlWuwTga8CTEY+Momveh0ac8yt0n6On2JQNsBbx4Nn8An
PTJWseY6OyGU60I9pTMyF3rLqdYZ2RZG61YqWGTTRfgA2hZTW+OMqyR+F1abwOnr
xxYdC4uCIFquAu06MsCEBsxEqmoSB5wF+psKOnI/hCvWixPj0KwXzJfkBNhSKBOE
45eLvkQqBZ2LdEB474g2O2C2/RDCWzprB2J1ji+6e/oLPD0OJhunVWbc0ycbHczW
wQis26X2jNnIJlACBOyg+M/mJYDqrX9JaDTB6VBoZlaWlU3leiDnlYEK/BxnqTiy
AKpBE2PfdELYg+xLKP6lH0yALsxnIcrJ/pnRtRBvomA0n7Lcc5V0LtEuuywjdRai
9/TLToKOC5/Knvoy4lttd6chgrIWHkj6VB0O+dnAegZyZvo1S2/ywKLv7k5YQZBl
l1SGMT8wyKW3G0UQJX8z50QB8Qb5DAYebwwsnIgQ/yFMeipA48sUDX40dTVk1aBS
eQUjdcvNj9AoeZgCLxo6yVefaHS+LSDn4n6PTddgr0jFZYhbs2YUZ6r6nGK7w2Is
Rm71N5/+doXVh4/R29AHYTb32HYj0vmfn334Y+JJYwUMraxz6s+g0WVVdoUG6xFR
LOmzXWvAKG0QKRWeTZF3SYzU0KXU/RUrC8cZ8MRJexYNTOE0t/EIGvFycQlGPGyr
0eE1tQMPYvmjQicQQvannig1BZOpwz1nkliYeUO7G/6mGCi8jT8A//zTZREozPEo
om3H0JoHgi0JvBcoYU9M5nRE97BxMXnUMcpn0/A1a0hIAJeDwd3lH2u2EcQCpg+v
YZpgU2cbGS6Ciq98ITshEgMF4o+IdcoRp5p+Jq5VujsfTS1ya0W1oHpKJLNvX0pB
cavhq3OM9qdRAZWPaspE2Jg1wJU8liQL7IVBmlzv588J8eoBCnR73IERswnpXgva
+T0ZN0ThqawTsYb1Kw4EW0MMVPqlYwViHdK+Zv7lW6XYsitS5u6VOanS1GVxtL9i
rvqTSIy6cC7xkvDGgbqfOghyi2UvlVT11xS4sg5QTL7cFmSBTZdMolhDK/UHmodY
nqt+mUpuq/WDdvPCX1TyV8V30eVvCavWJ0AyU/IbPWwwW7BEtosgqvDSpclCIWvj
D54Ov06mgB2nQK9v5ZRzHA==
`pragma protect end_protected
