// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SQZzsIukOoj3gqN0+sH7GK7Uh4w+Lu92aNHuTTojY+4QOeIHI+7QrcHT8u2t/P6f
4chbL8bj9LVt5yR0E7RUiSg804facJGXNUDyGNy2tCy8usuZTWTI/ZusuttHkK4l
sIx0/XE/N0B1q4D0W12y2LTOZ3O2+9UgiNneFMqTf0g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2784)
wI0JOksKXgh4luTX4XHWKKeK9dmso9igaPfrk79mLIR5hbnSZQ63tDGTxt4juU1Q
GyKTfqq1OYBf6f1ctwTvvXupZ94BDQF3jQ9L+/o8xKuohOWQhZQtnNRbWgNryDrE
HAriM7e7aYNIkc6iMKmMZ0SPpq8LPLe3dwWyii+S6RMxRBzkOL9y9v2e3rGFHgsG
C72pwdpF4nHqEk7a//zLZyhm7yN2JjkQnwtBCJYlg60Jje0y+UYVu47b8OpJjvDL
xWVzi6H4oTRSe+Uj+0Hf5yA4YAGYxdVYGK3aSOSjo3I1YBZeNnBWDnFJ/HbQ6Jkh
HtJtm2R5OU3GQwhxIY4xm2FMbyJWZbl6SxVC3xo8X6jdGvZn3UOS+C53utlfugHW
fPb7BueBiFZul39T+ubUpdNDuYtNAiIDefeoyrANwOAY7tkulSNzd4XMEHu1p5uN
u8hcy/UW3vYCiPIIr8DYW41K6mmFCHpIk9uxqz4DEyLOb+VAxs0vfP3qlGFxQE8C
zrEETT1Sl8j9Rmp5DI94A9HqzU+gImRAGECouQNh0/UWMpob183TF76WiqBi7sWX
0yQnDjKlN5+UsYTWPNPBUCem5sjXQ7nmB40l3dhUMLnxChdrOcQiLyKW4yfmBGB7
OonBr8pZiTTB0KDkoHp4WpvA6N/XWY+GduJy5eS5qczegsimUM0zaEIsPz8A9CjJ
dWPL/PrUAVJJ4NT/7cXj5wwQrWSxcUjHcCYZ2uhGrXqPozNd5iJifFXJ+/do0ocy
7vN6HKpVPruJvXPlccrMTi+IAIS070ki4Ll9OlCq3mATyxoPCCNb7fQcfp4JUBLU
Km2mMuAAuO/XB+QD3bnIzFffwEE5iZLUyGNEPdhdAyYSe9tuRFIuu4+cM5LbnDTy
i83jvTXNh8GH8yPveBn7VD//UHJewTZJdPlGalo6csv5ujuTpKTHlrmqf1swx9SZ
NnaPhKG8aC58FxvN8rEjDfSjpGHQ9/l+LpE5jNOTuYt1lnLyTEqKTt7pN9Dt3DPd
pGlwUKjpAfVp3LmzCtNhE6fldRvgZlyv/4qz1SCxpbx69uGTQInOV2irMv8x1ZCk
Mfl13oPwEB1SIjAUZp4/lU76I5mOFJ6O3+7CsqY5FpZrn2Hv+z+HHRA+RGBevP0O
6KJHF0nimBRfbp4Eg5ANqccIOTAp7bnMMGKpz3JNVdCUPoWhc1cxokLbldDAIlfv
TkUYsxDaKEIEVU8n8tsZ+NHaqdAGdl0bI5KAO6peVtDckm40Mbf/5RXfNIBSRm4Q
VLGq3Sf7XxTPsb1xyZ8VyEOISzIDu72aIo/61gx0ySeco9dAUU/RlWhlSLqlgBI1
h68aAL93/v++EoVhgpsQFJzJvsKr6pBvB+tFSTnf074kHIMF7xZLJ5tzfH7NOUfe
QBcPQ/sMoVV0VjTgUOnEvQRzIu2S7c4UpJQO2gKAlTm8rYMuRA23/0CTtIGDYy4J
RO4LIi/hJU5SmmR7qXfp3TUjVRrJOacb+QWz/e4figO2JQd/LbPRdGcmw3NB60jo
gJeQiRZUb9Fe6prfjEZmJbi/HmKX3nufirCMTmLrff9vehVCj11mQ7/tksLmZqS2
rrWOyh2OdX5oaLmnix3OZ48jBKilCL4gNY6EGjzepht7QaRJBzYCWVtw7dwh25Dm
Bsw71493GkoM0v1U+TL1DApiMsEDeuE9IyxwPi3+itHIxHV5NlUjFau/KyIyrJqp
89VFEgXXvMtCcHknSU7Y56tmDVSxIYSOspAl+3fJD/5LzpCC5feFZZ0vqJRW1BaQ
r2fQuewtU/Vi2krme4ABWWmenpm8O6ad25SuawMU6Ot8SA+CZfC2h2DMPsSikEG+
iHww8sn/E84MN0fkuuT4NGiL4aEl1a28jUZAb9CC1tIXajlNEedD02JmdlwWIAtH
BSjyxvoxWzkASipFdKOlTRtarvssIOxJOOU1IZlx0ZP8mchFliPg+gwtxONLQCYU
wZE0QXuElZ43dbj3bJR8vqOlyuAfFVjMj/tqHya7Ru6JVRsPabqojZRKIcBDSIov
NVFZiIn2ZwMG6qIqz9xGWdxRMohkEwfcM239Mas7lQ3TcNWWPyaNYUZElkLDCcxw
xtYnMBZR1dIaYOO3d2tKhG2zh/xu6xdTxMF8MnbL95xFEmi9JsxCgcTh0tkLUQgw
+avvqNmoogs2esc1kASIfEbX4L1mBlXrjVNsyZcAs93Qb/dcYDjJNVXtVWFfnKet
iomEwiUVLfgmW0DYwHFICwwey07TZeUUCNoR1hxkpUjp7GeuOc+35hKbipa3F3Ep
VjqosbDU3oPisaN4iHJqKfx8mfWgTxwO43NttorzlkAadJ8aoMWFXl8iKMjdJ2Z8
iGCZFiLfjqfsvXx3PXukMfrUPPZhQ3vjx/Kxoz3q4kW2kSAVvvRcSpBOZ42+RgtA
BhhUb3bjr2UPrn7KMubb/Zio7y77JaTuqjT7UNvimk4k48+tr8VN/P7fm2TYCIoa
b4aF4CdpNLf5oqeWFfalhiebqgAgpo80JKhBqjej536MeBOCACSfIQwAEY+V4CeF
msZShujgbI3XOji9x+ZXiQxSFCwcvgoNH/dIs0Va/hviE0DMmMQwmzmFHx9+np6a
V6GZut/ZP2MYMNSI0Sj0j7bYrde8L2kpgLhW9H36t8/5liEVJgeOnPhVME7J/X/c
q/IDerStPk11f+fW95Sh1ck0ePL6BYRxTeotKMBjYL3ms/SEutYdAb/UnBX+lBWY
15q4bHdDwaGe5CXBlBVREx0xE+4k4pb/FubBcKuwCYXGWwfbc/uKFCRa4bADRR9K
RoKTm6nG9Nd29LVnQGyss0svBcuu7M+i9kQz51hSJ3SDyEPP8YTRoo6HKMrl0ibN
9rKSBb5qxIxsQXUJoVhflEN0vQrsOmAsITlvBus6Qd6gpE0OUAslSEb7qIfrDTi7
jzYRYPS2l1YXWhVdfWrLhYbr+qcbDooWpKlpsFdKfncd3fh8FDScwtqDLTxf9lyP
sPzmcChZf0GR5oIqfqtIN3Ql03ilpnKV69VVsHHGevWDMyuJGOzCZgYnYTmXddRY
0mcZiw5kf8OK3vee1HExtmYblvtIjxLC2G/i7hUYYqsPNhyxSja7spdWKmImTCVk
R/ckTcpImMxuLks7YfEnSXCFzMIaYpkVnr9V8kAjDBKPteXG7h9PDNec+Yy3y69W
96Z8DBKZKlA9aea5cBHIgIfBspp9bC+HYPrCewleOFu0moJ2uZN04h1J+4AVOD0l
SbU1v02vDpKLVyd1ntvyweIzv5J6SmWKxp1XPZIA9x51kwbDoOzUXgR5T095ir0x
XFYGSKp5rw0z7UzUaCnF1hel/p43PWZAQYLPrZWCgjcUCZpLxk1qD86Zp5bTeAEK
QDMNNdYRybK010vJi4uBfcSRBwsrgENeU0ie+/ATT8cyKFJvZk/3P+1LtG9ANzUt
Ka5YZpG8R2OAtvyBDDua69qwZiSw446Dm8EfeVtzmw7Mt0AVuAdMSqppM1yisWeM
S09S6/6ZrnHJV+OIsjXf8H8dWJ7wyFJ7JXPmIje9A2+tomvn7e/wpcfXlyJipRsg
Qm2HgUNn5xCDztijuWF9TEwWnwgs6wV3zhIxj4Bvmyl7C0uXa8e4DXuNKOTCx8/u
mTrWPWfDJtdLuxb4cu8UaTMhpVEYSHl0xhO9wx5ZGUtmlj0FcDPvKOFkyyf3YzoK
`pragma protect end_protected
