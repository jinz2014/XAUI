// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FcKtVOOeNp6RFhbCS0/dAM1GUpxxeY74C9oJ5sa5kX22LvF1iVtlNrs03Mr5bXaq
6Fc+kARrTKR375ZQ3OsDSy3nUtO8YF6+KFmzxvqshVuUKt8GAChUS2UmnHYrGpi/
g7cTyMlFvLnxyNlGhu46HDeH44BHeXa3Ha7uyQmvwHw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58160)
wvPAo50nO2sDMl0Xba/JGAJuy1kydhskK+ztVuZc8ytVzffm3lIFu4VzmOoOQ+Bn
31qIEFRJBxvMMgCoGtrgxbKO1DCOKV2uQnJuSe94l5eQNUcC3GZi+whd46Tyl1dy
JHrVDpHNRFJ5pzR2J/kZnqq7a4s2LRcPI6BulD0dNMTk1brGbAcUgAk8DSa8tBVu
l509g27TM764j7M7JcxQGgorcIxUh9D7n9lpXhLbDPqHdYwzB1MoJg05ldcVskuI
p44yDwy4t4Jj/IUgr9Il0vrfOhWwC0emBg539XC6j0RXFLj7MRTkbOsiGJ25vjie
CrgyarsTHWPqyr86Qbt10Ilz07E+LeGWHmmx46HUPbCvxlx1I+yPM2JqoArbtSfF
GJQaqbWGOGBtQsUu9Sh5jZgraDgQi6VhIJrdV9KOqjyAzisQdL8eUtnmns19zmUM
4vwLQyXOazhUseR47/chogCUTrPHbNOqmU6ajZAskVX+e4UCWfVZVYsChbP+EG6L
AxbaT5HvEYP4TSzaSzTk6CvDirEyW9+HTOmP3ULqhRm4d1NWVE6ZH7gCjmnscVhO
PLPREg0FZepYeso8SlDp6QWcoJF//Sd4wV7FvgSdCzaSRwsfBhKqbpsSGAC0TdJv
VWsASd1sHhcNSsueI+s598Bw/qE4fvZ6sP1IcOxVjJFOx28UZDeIzVbT7+9jFGMC
OtX98ryO1ukeaOpziAxs5M3ALN+gQ/zHsWbzurnqL6ghlmnukshoSXFeenK3c9vU
pjh01Wcr8gPq2t98OEjfbo5efu9dlgVSCQ/giJooPNZsUJcQalQ2dPdk4JwnxsMM
FcG2bLG2W6sW6eFpO73SwUReZ5G/A24xoOCtB8U/uyI/BxKHs7mQ6FO56FX0kQ5S
9P8u4pV0Pe2EzKASHULoNwt8FV9qY8C1UqTXk/ayksBC9pkQpVVRI5n2lhAsZnaP
Y9O4ONRiNUAsKyVxpE2N2BhA/8fhMhzzSHQ0MKJdWqY6jIXI+EpwKtRbOlmkAIKC
zk4pajJVfVDvbVMFxHt8vy3FaMBea+gc+2h2U/kCW5uec83YFKrJ/utSy82/WT9T
FJs3dRWdZLY8QXvV8vKRvfBQI8lFA+076orxc+3NgiQfvXOhXLqSKtITdk/ly/Qe
cd3iWYyWET0pKXq74e/rQsc9Pkh9lxVRQAPk7d8L5b1XcboL+R9YXyFyD7iYmGOa
+/xUHLzJB38KEGZj5BLJXZrc5H5H3EhOhExypm2A/Xx37MCb69Q7jplnKlobxXfA
n7nenDtAMO3tuTOhho9SRvqnNlWcohlOl73Q4YzKrepTkiNjLwOH3GH4ENo1Gj/2
v187LGEeceLAnyY5ewpvMXWpcooH9bPRBgsoYwr6ErfoSXF7icmevSSGMQXayHwO
oQH3BKBFkQIhIK3Q5TT440OJtd60WkyTZVFC5taneCg6J/wvkh4LBtHvLdKwxJ/M
ESlHl6y5RpewW/QOOPG98xSqhtTkbYcB5/THJtxxkE+PACHxo87F/uZLuB5OkP55
4IxdIt6e8tBavPYixhoqMJDJz3gJDjKC4he9+uxmH965tmf0LDgX5hD72YEt9hHH
PSeUEMAhjgIbSeB3hrt4qUKL2FAbPSug79r/3dLPP4+MRuUgeE0yZ59JlzaRfcT6
MixNzBwrfeDrYCtWNxxFqXLJGqy9Qab5JF9Dc/DRChi5MbvsfJvZ3Vz/lwt9w7iT
4Cxpt6Nw3jP2JktHEmqxHn984PVYa6FcH9J7BGLN8tALbUJKPM3ON9ewD7B7NkSs
2Yg0i8HlxXoUxRQdXANNhhR81dimEKJp/mBnd3YWFX++vDa0xd33H/qg8ZZbTeXa
/Gg9Dwx4DVnbSMPHLZeR7Uqgf/RUNM0AOJhifg62X1nsF/ztgzKyoJPWL/OdZ7e3
LYqRVIc4lRVrIdjGlY8AhIWGN4e1usftbUmulG7/Rg2nxraCcbwjammWHhh4uSlt
eBrOVAyhNtTqZjBthsWObD8VXG2RqNNEQ0eF6H5wFNDecO+ZInPvzZUuYAl1WUVB
JGEpPJUhgPc8DBmQXivaIXUxHFQhup4WO8l+OcNtgsa7xOVOf+b3WmLoF4XQHOK1
/ickbxXP5+KqheV+lTSKeoDJFVfmwDP2BaXwHhw3AKaEWh+IdY4qyzTcLwwDK2Ii
MNpr47mIRaGM7SXgvBK4y4yJcr6H89LizzEHeM7bB85iHBHOCc+8pt9N+4jgP+A3
MnT+4wZAefA2Z0weqwY0LSAMu8LYjmAVKNDRfW154be7hC0/KJ0dCwmRAgQ1zwJZ
5zKfvYWYNFxpRfgP9f4KIoiwRXQSSYaZmKuH6W1qiBoGA0dRr0MyRyrzG1V2aAoQ
tSvJQDS96+t1hquFledpPsd/D7KsRe5ZLnJYBg7yf92Juqm0uurEKFOWj+X1qUGk
K9oo/evaYeGhzgRDht2fJvM51FWGBlErf7QdxjmyhGy63IHHWlaJ3K6F3AFPcKgj
q0HZLYuOmkCly4ji9iVDxKeeJJHyAkKTJ5a7QeNzaeN1JaKbSLdyTxZoztY3+AWQ
hfy3HTLenGolGkLds14CeJOPd+Cru1pHJ6K5Gpl5jnPaRtzxHoK+MGBBkHMgexZP
lDilkWoInC4cMjtIVBnp2Fx2Px3LjggsFT/8PN8VMPIaR+erNqOxvMmJyel8dQIK
ppFuIPVOarF2CAar4PBnSQAbvgC59+45/uRhiors4sIQxsLNPx0pX+Gwur3SK80l
SL8cSxFzEA/RFUp4WoW9ruOw3F7I1sItfkJCEw20fL/Dz1+rPNca2XYwXI5laOzV
a/CCGeMUjmsWrS8asWl3tp/Z7Fw6Bw8Or53xhVQK3mqL1gYWrnrhb0uEpTESv4sS
EZlRnqbHVdMY841FN938WjapmPoUI+bqDAuuiHoVfrqRdvbcCVYmhAEsoQnL0aLa
PLe1tvEaJZI5qZevG+A5qNudJkmT1o+3ZwL0lI0NlBux9wwnlDMV/uTTk6c6PveW
2il70iRXdjjom+7sqYkgsH8YHSd8ypjR47W1abk686OngorxhkdxorDog4kZAtEs
ZA6EJUKScAiocrpSR+aIxV/E1wO3v8clEylC5D93mK9GHyMcjEBPmJg/j99HWZci
on+8+h6zvULVvecb1ZpZgKolJyhUPJqRE+Arz1/y0/bJqYSfHkkmZJFkyucWpcEG
hrJJk85kNtT9HbtIP7xR6zCrSU/D4/HN68tvnoDHYfkQGo+zDrTljH+jskI2gpNy
WLvBk4y7LEinAovlx5nW4qphp1Ks8reYHRGoXK1zvqkOLD9Mle/a9yV/JS83xsZN
hxLsAPuk7Kfb4muOI2K9B+O1WNitrnKSeoPyRyKQHvCQTj7O+W+HMsQFGYq+nNBi
aw4m0ljgVJuB04YmE6pKsCxUl1I5HmlXoUDe4e8IQItGgHGREnJS4s2os+xCrWTo
h905gHpX/MkyjolLP05RFNhieBmKk3g85aLKD7slPjDZDOEh3r2Wo2yA5ZMEPP5/
/T26LGcb/T+nYInzX1E+XuZa7INtv260f0q1N4ntJlk/PlI/WmsngPP/GhsbMFrq
W9KkOcRedgSzWaumoz/RWnvYGCICKqN/EksQr67sBznILB++fvUjrQs2UlMg8SRO
8psUOoD6kMFSxqKysFmbrVUr5v2coU4UW3u1kvjZAcPn7AC8tbaYUauvOWsH8ktL
ZY9zDY2MzrWW4KqcNNGolO7S6OdVJlOirK3KvbwlPTuGNdK570tf1styv0QJrMJT
JU5V0n0FPoiym1ZMY93WXxHwkp39LWU8BNdrqGfC5pmahFCjeu664Rcm4LfN5tLZ
WDqLDGET5I8+j8OsyJzNMIp/nGvR8FdePV9aK8AXhHrpD4HLTD5fXfdT9t15DacN
9gDfeUAz7LHzQUyu0ZqBIlgR4YtbY02AC+/g7w7+lerz1h+Qb1E4ZYqLoRhz/Boy
eocTkBy2YY8Xlnw/fAb0eZ27a2O9/tUEquWAk9MDTGJpAUh0PzSNt8aQ0L7lCdMX
YCAEJC5AChTsk98vnX8EsDN2n6m0UswlpRNId4QnwJo4/Ts73Hnqv8qGaNplK7DR
kboHD+HNBSDCxVczonMJcXFlAhgKpdkFYsS3g/CPsUQU0tX8POEZ3a+3S9h/Yx2N
nHY2iaYlMpTBowTaGYkxq3uU0jCxiPaEtCyvEzTsqJNIhv6beDYp2sCn4p1WG2g5
X9md5x2acCYTSPTEkThY+NNXfsYsBo0Zj8tz5LbJSaFGqLBoFZeWLBKUvOFp/9Ku
y7DYCxix5v4QxIyp+JZdsnmAJ5UXmxdZmlIZKpcD5qkpuKjAnxDGyLST3h9wVZny
2ud0im378Ns4Ku5MxwHK2pqL2OehJGJvtJ4FBBQvT+w00cGP0/F/VWh97+Q4qV1J
xqo5xjrnujxhChSNGuZJgSykQGQkFd5zj/xwb06R8Z2N0RxJPwyC65ef0HEPRHon
ho1jSlI+oVIYHmLvS4HrlPmCHF+vKwwZ+CCoJ5CQUww7sb/s++LOJG4uea4mkrbk
nqpr0yDMhnmfM+YRL1LUOzuDyE6Tf4PhQ/RLjXNZvs9hF1WG8Vk5wYoh9THNtj20
n7UKXs4nDOwIGuyO2LV83ABo60Jr1gTKkrWD/4zCPo3k4ElCREn++IC5DW0yTv9B
Tv/8DWS321HxR+L4yqf6cbD/KSyfPqLa+rWKN4HGCr+J+iTqtx755zyRVDYN4L7d
/O2mdd0b5uQnp6J3k/v8mEt7gmNynR8trHp6jxkqeNolaoygf8hwsNOq7MQ5Z43w
9wVMnl8NileID5idjp1S1XktZPDtYw44psztzare7qn6nchFhbYPiqNw6Qcq6tfl
z3FQmRZ6U+yhfnl3ZbuJLQQM9zyk6LhwZFI769IXIfKSZm/2xyNGWvF82l6kiGAz
bNuST88OHtpNJFFnlPXgvt48HOr1+HlmQ19SVzkaMoCHMyKOkKYj2EEKh37wWPlk
/wu/Czn5mb9At/K5FXM5VGGweem0/uULuvrSehidJ3DOweUU1wbqTYtsN6vgEtzO
1K0FzevV8iot5CDxHfgtvK7RnY/paUIzoa3aKFyQ+O9a/9LkDRBFg82j3fwNHWNa
PBbdRvpndYN4TSu7baq5znlGV7USbvgSQtk9yoGEaByp2IERVK6aQSit3WpNyCFK
zDc6iNOt4BicBefbHgPwBvBiiLLIaNI0SweeFhQTu7HFN4quyGm5GO5x9xxBiW/0
knhNLxVqfcA3XpBn3OqMUvsMZ3a4er2fjQBVexs/SDQQ/FnZLdEko+G+dJaDMSZ4
JVxuCMlZ8GEFLF9C+ZTVP7nMPNiW4vsizBWger78NAXmUvj7jfGQQwYAOdw2CB6v
Y5hH3aDlU7PtqnWJERAY7l5C47U6zxI/1zvupgODjAzv8Lz4LOTJVbUit5N1SsXt
pK+FSAI4GCwhA0rGDGib2+hNjC0B05LYBq+kMqGBIRWRbptuYwY9JWM02w4NCQcu
3nJytaFHD2dpyg6zqGGJghbB1feuQ+00CrjjAF12Kp+adu4w2xmRQimxqRE1AevP
a6833+SWYny8Af5boOCftVKpktbBLmTm0h8Cu9fWfTSieM4//VxTNHhrzQLRaMsw
H0QfiuvTpKfzLE5cEOYKQXj1DE2G3GM5FcOwysw8CubZXRH+86hIe2tbGHKspvY5
I7hQ4kDkFmgdk2eZvxJl6kqHI7ZAp6cUOH9jicYOd6FToH3FK4+YzWy3WIBABKmd
wBMU8zH9Jv2eAs5EXHn5XJC7lMivQINGGMsY5cl6WjyiN+Kg3TdOuHFhX7aYa09f
jWFfkKSMiHys6PLmcoJQ0YGYEdVOPC534fKwXSFIxFhE5OphBfxV6+HtYUHjFS+r
Whnuj3tCNyABIM28MwkdCfdG+lZy9FxM9F5mkLSwReuHcw7u73SigDXMvp9bDcL7
8Si7C/1u5dkNPKqd0O/n733kqCbRfdTFSSiToj3N25uGLWnjKyWqxmJ1mmWiDufz
UMmvAPWaP6UekVOa9alX6vYYEIQ2kbi3SRM7sZELEk8CZn9XbATGJo4IZR4rSIok
qSDhh0yCG+n31C4rKtoXOauUlv5JHjKVjTrr+P24ve2yOaGgtMhZHrD6b14dA82x
CXh3xXmC4Rg0hG4KcpjEEfJm9LK64hiXXyKtyqPryK/XClwkUiNvS+T69i5n1kO8
0gPt2Fp4/TAw3qLDUM7nynTbww2ocQbEaGRIUpAEbAlUCNcw7BizqJB518j043Ur
tPcG8ApitbTehVVg3aqbp24gFmO2cik1o8gE0BZL6g7stnzhySkde+Z77T/lgWVo
T2MYkgjtxeGyJ+8cP+rG1gl7KcAKp9UMh8NIN9p8oUhP4y8jQEgiG5vW3TUSMPkq
l2N9mVgXS9G5PXivEup/NWIvKcjfpeckXtkrVPrKLgroycNg0kaKT9eZ/QKIJUVa
0qvWJlu5hIOkYRhFlauVh62rTaLGJFWW9Ix3aRgL8mgxfOtl22HMm9MebGOaj0Gu
CdJIKt99EwDyIVFIg6F6XW8fRsSI0MWEWN/d2pbozS99hdznn0a7/hpqpAD0t0tS
QXiBo01yGYIOaFycEjmGWQaAtJXgepfs6HC0qztxDvkS7xWN9CQ3P7QkUVx+PGBE
sgSzfzsHT3eRunprZjfZrpKWZuCiIAufd4vvRyHFnMxPRW0o3xfTnyeHZe0GAuEs
AEcsorKdJgZtTwYgdV5eqkhO4Sz3dFr6SydTF0cXDFf1fqecNK44odvV5Dotk50S
mAgEeJYXR+ux3HWqS3EKszEXo+wjDaxNgPo1X9nnvP445bo5qCEM5yvdEFJ0pa/S
Wf1jA57HM/wvpn1ktf5Thx84NOqBglLv2a1DIteivuqbLBaatBD9vZBoScm2KCLt
aG3E4mnEUiJRTVOZKWPDJat3RYvyEhVnwNjmb5TJn9OrhHCbKbvwcrsUO6vDEjIP
6Eyhj4WplYupCZ2SZhzWheH8nobu4EQZCogTXvIeeApcgPqd65lkmC+C5Cqlp272
g/sBih1GCSQP2YRU9cSYOlJ67IN15YzbWq2PqbJ0XZYcs4y7NoJAuL5ZW57m1Pqw
xdJJx2YaPVM1i8UfQxy/UU9iiXplRq8ggQMH/nL6PqkcrtdnCZX0QUJDzO3Gf6Ub
/V7Q/07F648agHajRpufmWXWKyFuuH1Rmwe+bYCGMCrJPwJcTjNpE64RdpU2culb
jlxbGYf7PuoIs4IAoCV83GLyRNzgRKe7/C6CiLA3CpweLMX6q0UdmNvKVhD8of6+
TjZhHi3LvanZVEo2wU5wNd0/qdySVwFF5WtsUyT36Gu7wCfd+7o2KfuhQPaMXO7u
QSSP4GMHE0vV8mo/2Xko4BuF/AhMObEJ+7rO87yw85+skGKjv8P8Kfw85kQMblZy
DWb6wQA91ewjeESOjxGJ3vPgUrP1bIQX+ovuXNb5gtEecKl3g0y0KwvtmBM7GR9J
Iq9uC3Q2eMtjwDeI1OFXFRV8uaEjkZT0fKN4c0341czaLG4RmfvgQxO87G6IXAtH
TCKp4rOpPawx9kOJq3rzfLIJUsIEGyNOGtr5IlEDIxNzHq1M3cv/8kX/d7hON+Oc
M0FK/Eu0TYPP/ugQ3WO0NQrF40ywyo1Oq2xbly0tU56L3sDYQOOqWJfk66bTYvHN
2VuTu2RP5XWNtBKHf6PfDTvBUT5lptzU6+v5V0TnT9uHlYYfH/HjmnkOM9p63aAm
w+s45pExxql9vNMZk2M7n4tj9/UgFX38KcFpMBS0qnBL1itUHyM+4BsYbVgCVnme
qb8enesYPAGV/b6A7xMRUMbCfcqJUJGHsN3pf5gdQGZNmkaJLUHyuMgwu4NbYare
1Y+hmUWyJewIHP9XKLc01U8WCsNMPDcD2ULKcPsx9E/OAfrpOAlX3Nja378AeV5i
aZd4l1fGQvK+bT98KMO1Exr7/6ZB+TVoKehM8gZIsV8vLiUjZsAxpOr8kX9j2viC
XUuGoCUqaFfhP3qAHY4k38GSPLK9ZNaBTqdOWdkQ++3tUkVdGcIWulM9pk/SK613
7CbwBoI9iLLW7ZkaZOv0nyNXVqc2kEfNqrKPsF3Hj6KQxNC0WzAkgUqu7zQwjATQ
6oihAgYP3lAXuSGhI0g26CJUxgYJDpxC7vYqobcuyzlKWFoEq3tHOiem6dY14/s6
WJ/niD4w9B9mou/7A52G406hMmMfwqyePD98+UQF8vcOW0JzNjGE5ZLe2bsTuNK3
M5TRuumgqoXn7V9JpcfTeWJLByXthYqbVFy4uOkLNS8vFg0cALyvlBBtO5RHapUS
7pN3PisI93OQ4tVXqlhAmIrabljba/LB7T6tkvxuUgNogxjED2AzZnSedV7yRh47
0g14HxeWuhOl8RUHf7/wgaa/j3DV9TK9EUBs2VX0gdEvniRCsAiKHiXPwWe4QarM
be5/gadDetYA4RyZlVGO6TK1Mrpnqbzhxr7Zu0kmBzZqxGg6m5lfXZxPgPFN5fKY
gsg+10Af137p+YfPvfOPsgMMei8pGL9X+P4fdm4VdglkLPu69S1LKYgSiiSWiusS
hEI7Wd9OqCNXOAyFbt/HnhfzDBuqKrEA/bsquPnhyzENB6t7oLJwOau3AWBtMLWm
UyGQkL9xHscT17oPtfQvUDr3qPWoosqJUMcyv/YH3GWIymcKGMNmd1vtEHx1+Ic4
QnflcJwKgBTfWl2plBkp2iSljgNNGhB40CKrfg4wcx0bvoT0S8kSxIe7mPPvMQhX
LF3aUC1y46tZXzWgvt9UnpAI1T44vdNjraLsHL9J9HDKH0wK28rO9DliqWiQHguk
wUhht8TAHYTuHpb8kUAk+Y6WgmxQ2Ep9zN5eDrz22xAKRGSjdXY/ohoIVXS8XrcB
LgSm+ljnjtG72aegyNN3ceOjMwC3gAIyYxrK37i/I3hGGcRnEsW8puy6gQ/d7NjB
c1372rA78yV67E9Wt1r/xy6smRItSNqp1Zr6BZj2FedraQjMV71tLeLQAQNvxhdc
aX3yKF0LCTiPxmlm0yy1W5uOsOIk6NHm0luS2FcfrBrp84J5LljT43x8IdELkRkW
BSsKik0E2OtEenhWafGr0t6Yq1VQie+jAOJ8imTEc/veIMXJGC3AM+rd/WOYq7/O
augZk3e3BpuXLlJcoL/UmsONUL8F7L6iVf5FvbQnuDiFDnFrE/hCu0aNTPnBANYn
55Kj0UYrzOS2TUK76YhuhFuOughr5GyvaHlVLr/i9rpdytXCD2JGmjR8uokSKOjd
SwBrTH+5KUewpcVB2PsC7EVsqfb+QWts4ssDkd7YvTpz71bVD/mCwAk7AGCFXuBS
rQbiLoDjq7cY65R0TC6kxrqhigX4KVB5tNMIV33c19+cyc+vlHdzRgvTaqsu8lmy
YUNRwbKr1g5Fzhz80LIRzTXEqWSBj01Z5DAXHAcClmGtpBf5S3J/3YFMQj5y81Qt
cf5qf5Rda1TbI6bDd5jJOIBxAr948yr/QB6qvEFkac9VvYpjxQwhdi4jgeUjhjiX
eRX72xtkW2xmvu7fcu/oe60Ub4vZuUmqdAeNrtXqfe12FpELlujHCVxhbYb9qDFI
LKO1de2qubdG0MjfCdlwIRASv4DDOcqoHs9G2Wn83dcjoq+mbIZTnWW4Hmu6xfZ9
+0EQFtWUbMnLe5KD0WczFqDfwuZ6EjpjjGbQqEl81+VXNnPm+s5I+JkSTzCywuDa
HNEwvfKvvARgkweqZEbcY1tCEDWxtigFJpYC6Zn/FQzvGy7Sciq/YOj26vxkS4v2
lWVVVMUge57txBPTHrOsxsOUQIz8h1fHayi+4JwmyRuq8BR0Buc0N4STqEPNKgWO
Rw4IZ7fOBSiPCvBT8DDfkpkiI/cMDsc26rhEXbfn8Dr2j8XXK5X+8sBXjr0p2CaV
O8z0fMI+ijKydE3DSF7L0C59jvVaK8T3YDcjRQtshxMCqgppp0y2ptJNIi/FNy56
S04JMN3tLbWUdzPnSkd+fNMCybYBVmd5CuseQZqBxgy8P/4QAgsZeIqjmyZYd2RH
NnKg3DpfmFBn5f/tkNy1Jpkh2aKB9bOdebaGx6x6X9Egf2QmPk6qjrgoL+1K1Dq4
JV4ydq1ZzPH16xhRCiGQXOfLIsXDxTKCnmSWLSHzcq5ZaCFA63RvdDtuCexF27aR
yom9DMC3B5ENZb3NlFeBpmrjKT+7GwfGehV+d4i3p6D7QSiZesPMU3oF+vMvWXp/
NQigIJXLz6qW0BDfF0PSKTmX4rhIEjjJk1jGMawMBMhPRI+RXgk2SIgDJhf+UmCC
m5fyX/dKsJtjaDn+Aqn8sfIF4RduHGHb8ClBSNWV1SY4lq4wGWXy6ShvkRENMuKy
3kIToTrbkakzS94ks3PADnAt+pEF5Lxh5VCMymxGdkrnb3uYt+m/CBJKU6KKYNUv
uCdNvPJfhMAzGkBzOeEhyyQ+g7yTiC+xuJbK06o8Gy9cgNKHQ4y+7XuqeJW4I7MR
hQ17DBKxWRSvgor/2yYf53/0QLvYiBLz/PYljEpNBsHB2aSpsESfF4tASrE+K3uL
0nJhtCwSjivZrxXDENLUiVmvUxAI0j/rIo0kDjNShqGivzY+ae2BwMC6+UEBr4XD
JT6zyRxYaryNAeZhFLhcHEbS7/xqZjLunkwrb4vzN8TO8+ETEdAk/GO8CpCCi1ZJ
id725QpQGEmaIx6Sv8b6JmbPT57t2hTYyK2DFxOp7tr820l2SbKXQDw3ERq+CbTG
T0nZRF28iEBETCH5aPVBakEakbg8k9ylCTQ4uO49mRCiQT826e9OqI9HEP9uhJhW
v3/z+Cp+VnsYH4mxqvn97BkT66VhHxqe42V5mtTJbD4KKRjPcBo3zb0qeXwWrj2n
KR5zedb4NZaVDz4nUM5eZCpFSHr9F3asxiIJ6OVNbBftywDY8VgkQXlcACujU5CL
r4kf9VOn3iI7+v2u8Nvw9KskWcHtUB9ktQI/p1bfNb8bmlkY9CJP7v4l9hv7sZI1
fZEm1UbDwkFUqq3oUrJbPuTlVTb0eAzM6D9L+eDIrxJLkXEVblz+W6JZ/7utkYlQ
EFW26e+jU3NuMT2ujW+FWFCzj8LHAJ6mKJN9Vh/Z/jduQgQYkoPnaCXUi4aqimGi
riJecJkEUkTxlUpKoQQCy7lqFYGQxI9r7/gAmj3DE8z7QZdO/lMsGQHOtkUHWHuG
tUyOisHaaNo24P0p2uA6anhDJFJ5Z7u/0uCjh5ykGM7p9+iEdVsGrSYJr3nNVbdJ
nlu2FmppuEpQCZCcmJGi2giJx7ZHrBzDABbwNQ1ea0GKf79KOTEigBrDzja4FGtW
qjyFo+8pUAzjFtvPUeAeDtjRBSUY2+1EnwtcEe9kiHxj0OTPlPDF1EKNPtWXJF/v
BKREUrp2b8n5aZmnTkA6VJznYC6AnvaS96ziUR6K7l2yeDVx48VWWkQ4r3wKfNXY
v4qDTvq4g5KtdnhFnu03se6fUiBexf5ImZKFjWfhwgzBqV/bWLRcYWLU078fb1m8
3pVCf1LEne0WRBlCF0uxo0uGr7Oz+ju400kcf/9Rnm9Ds+/n8gLM77fvmz8t6k3/
POLTNwmbOKsHvoa4wYawUTy4RZMyfDhOUyHqs51LO46NyAnoPHhf11786dFAuu9z
VDb4fD9ihKbGtiuSY9eFCcxMPPaaK2YDu1W+7w611zwQTz8Nr6p9ac4/ycQ81O7Z
QugRJCjDmFXPp7ojjTdGM0xRXuxr10kNTZUWSfq6nFwOvhGwcT91D8vx3N1yxRD6
QMtBR7xgF5mGOrUZ7WjBkeijQeARSEQt6U8IEF5ifpDBbVzeJEgEy2Vt7k1oesXZ
9btu2Rzlv9UywpxgOI5FD+HWY0gZwprerNJ8hTX08C/r3svkf2k8Q42wbghgC51l
auEWvkEoaOTPy2917O3PwXKAiTPVognCzCZTQ3CC+Bb7AgNqAtUMVmY9TCvWUMj5
YbbegXXrU1aRT/bCdLVSOvgTRG8a9CHLfzZl7pxQfDhFz94nBQSaneCUbMWzhHiU
K5UExIFXvP1HccwIPlXIE55OvzG9B05+KANSLDPUPLRdtV8tCfs9chOAfdU2DWDM
M2ZAYNkkifEo6kzqoGXGiygInxsHPgXNX1tOFSRFKjEAmhPVnWSst7hKFdOeCNpz
aoluTUoWZ/5As8aYLCpJtYoZjhCPmLq8Byyw+UBYEdBPppCNS4+vdZR+tETiz4Kd
2gQ/9ucG8xQTC+d9Zodjd9PgK8nj89BB4iLU0dem3hvYWyqqegUP/rs/E7Cpl5QR
CqZg6znib50MnLdiJAuYz1AV5PaYMJLC47Z+2XmWVARAT73H0FXgStHoIzbKjtpP
/3Sgv3MnxRb4eBRzIsScr+qnJljgKHCmTgc6XrHXTEwADx+1SZotbDF5deNclKiw
h6JsIJRqnMpZVGSSR/OenDjH98p/5eiQCG5SlzhJ7gr8mZC6Yv8cLqKMuaCtwvAp
7ikmTm46jBoMXJSVmH4tjLgExVfmpAjoc5NVGUYy+x5axy+CsL9+oy67x2tc4B1Q
UlHglwSTynUjyKAhrzJaQ1x7kOd4q8RXSGECitjZk8BIQHCpTKkpEcPVDD4j0sUk
0rXWeyxsliRusZUNKCt9TYhLuxNtvDwGC/jRbSOZYISGM+uKH8NeWOCCjfXxkDg7
QdP0S9/hzBBqNF8kJjDNyIcCOo68PWVDfPfJtx9sgfA4HNGABVtiZes2/29IZVEf
KXNC3DXZF7ZtL/tJ4J+dhfOiE+iOEDWCiVmyoUTkbPKW5j5KjFtKrNmZFPcTapQj
r/JKfCipigloJmVfCytlg+U4C9h60N4IAbu2VlcEzEHpIXUrQdQI8X+jcFr4PiU8
t9PBd7OAbqpMnj14sa3zYNcmNB40K5leZdJIZw0oKy11z3bFHxvgGuPfXBFsHJCu
Ii3oxmSXyjYpTuJ81rNop1NH6kgQgsMAxMkhjmRz0eSWjAZHpgJ3O4ji1V9+X3WD
OxMQ8tGwjDb+cSxongNO9HvuNS5GEpbhLKBri+tkqbsd5E3NVNjFUrC4kevnWzlE
b5yTpJbypBt65IHMWOlNNgmJcCK7u64V6z2TkYdX4m/2vblsUPrMumPaT3vSYqGn
VgJExRrb7PoJrdttU6Pn3bumzl5NLmqctTnin9W01gGbM1i5qqbP6h+bFJsDikGS
GXxOGtsG4wDuR2DKZ74R7LllU9EBIE0b0OSSZmHGp+fL4KR2M7zYhNQR0PgjuQn6
GpeI76SD4Lpi9iPoNQdjUQyZjvN5tWuCJqr5KoLGTmol5uhHYF0QNwzYmp6tlNFF
yqhUcDyvxnqLBDeMMVRMo1GMZUmnE5c2z69eZ9PHXHMhif+PksxQon9SLpRR47h1
74W48s/vEgv/U7aPgsNsewqt9BP+ERSLEH1rxttZViDFAvPRhYorb9lnbuOre5eC
dk9DXXMJob0tFA+w1+cwvsoHtxYiTllbRHbMfZbZeznwMoOaX+0VUU9fk6qkG0FZ
Udd0l1gvq3fRZBKBNm/JU0deU7o75XTWwSXxgt4+lxaM8xWjvhNA4dvdxG3igPGw
4BecYxN5jC49xyif9dBx7cPab8tYO/NkIQORDI0GdV3BYYRKkOqYZvTUEUrJgMqC
M9jIUOsTfV5xBUjRt3qKgId+3PKTJZcmWl5dDtZ4I+3xpC+fPxQsTqMZNhgKcZPH
76FXoHUAqcBaNpnu4kmEEuyo9Z4BAa7O+8j7LzIAe27rZ/pvcouFCalejAGwRqzG
15+4pi3BLtyr2ezY/ao+VqwxoC2ty5NG021NHHFfN0d/giHc7sdfuxdIez/ZFCH0
8iUyqdStDxsu+R8t97wZ444Arb39EZpeuyMin5fwL0+zZxm6hZPggz/RKXc4XrUu
hnPGwQZ9Q0OIwyAnARlCT+G/pz9e935FRQV6xfkAwUJjhZTiJ8zH5+aN86ikh0cW
/v2WO/z4v4LjmCByN0XBQhdTV+H5m6SW0Sr/MrDYhrlqS5ntIJ6S9AFwZlw6ecP8
yJWAPmNsbKshnLe5x4XC0WDtiymshB44NBawdXU2quiPuT/cRtU17yH+TfJiDnYb
5gwZUz036qJq33WYS44kk/kckc89vwCg47tgpNNylYCsIRCfLWNAsX6QAPBBkwzT
3sDTweefUxrfkNIdqJIQXy2rCHqfklZEV5OYPK2ZQC9ol3j1zzjzFJsZjrs96CL/
zvT8djKCwM4w5PFHA8eFInKX8NoJTahtqXmJXgZRq4ammnku+NrMrTvA1peggulD
UhjO8S4IaH2Z0uE2cs6Koa9nQ7YyHDboydNOzD4SZAcj8KAfu5cx2Nj4abOvYydf
m8tGgUKhMT7aAgdN2C7nHkUmdJBaA6PU2fF1IBqpso9na+hIrnhDxh64n0GFU2vk
ztjhNLnS40KskWz952yw/xSSeSHy4tBr3WcWy02NZuCrPyk4yp/+aWCb6U7Q2R97
R7ptv9JbVnF/1015qAZzSo44Okd6qAcYyWF7Rp9WAEe5dYHMF2Nqrby2lMHpAQdA
j0jnK+JvQOvsoS2EON2gMB1nISEOewvswcS1OmhpmRgiqhURZFdZ//k3RCrYb4fo
R8fOW4lrnel+Qs3CP9CFKvLZMg93gml1XxST+C7Uskm/HNP2YHVX1Tjd5+XVDndg
yKicvuzV+azHoTdgYYkZPiHhij/yHB0wORtslOBdWxp9LQOL4n92fnSb49st40qk
iD5Udb+J9KWG3qIGPiF8U6MWUcT+voACJR13DkOEn3uoeaopngJWjel1H+aDeD3t
TczdVB6mxVzpfxF9/ENr/2O7o1+yqMwji6sGMumb5U/P7ieO8w395pUgvjbjVRfT
ZxHqCGDwf7N4DfU9nrO2ZVyV7drgN5g+aS6vKO2ryAuaQKxliLJWEygntybxbL+3
PKhGDAR4+6DrwnLZIOtxUOc1OXEJMhz+uXqKwpNulvkKRs/WFbPMpMYiqAdKRTBU
VOcP7TwApIElLrp0BeEkoU6rS2beLxt8o7nZ6DefEH9es5LPOKp7jXgImFnCiNzq
kp9rx244CyDYZMxpTksBJ/0QAPsq+xzJiHQvej1vcr3PaCgfuVOcCzoXZF7WKy2R
v6IUhHj4MLpXbr6W52h/0Xhz6hV6nYdSHjsRJdICz4aS5ietaeeMEqhvYeU6o/pn
8kFkPzlN7L16wtp11g9lSQ8Jvva7EvFJslr+eOOBpMDZkq072x0h9seYHDSPnWtQ
pSP9oQKaaYENUBA8cEmhNcjluGWo2+N0aYdBKr76ujA2pGI+vmxoKhTaT4HKA491
PM9TcjpYpinIJgqkTpNh0mq7SVWjOK22Vp9ZhCe2MuZ3FF9GEHulSp3V9r83GN/Z
kg0zQ/rLQg44yQqrI5PtosGT3NSH8Fh+z5DlfUfr8RP4v8DEWZNDZEdgfMd7pzHJ
aV4TfQO3l6wYMDvXnEECgRB3pfq70IBavqGoTJtxOVB8yGfSrpSVl+W9srGAZlYF
vCI3Cvt7z8YJ5C1KmJiKFVvEA0JoXcFALfr7Pxws0zAfpkL2QJMJJamOp8mzpwlM
tbBrqn5D0L7KUW/dNfzSAzv8vRdpm3iL8PVZX1EmJYsqP79yEoTTA9q/sxqIv65G
DlK8cXkhSkxlFCE4lINxuCv7C8Ti3PUA2dvlZwn6DhSCZxOsnQ/IKZRvc9aKvcb6
5cH0YdMEMRFW7ZUI+krcLm7hSzTkPs4SQQA5wBog8Dh1KVnDUh1sPEHD6+44TpLk
n40Ceq4Jy4Pwd6pF8A08NszFspBlyhpP2a+yA96ukeFRbbLzDYxxoKSqhC+vt8/H
MNN4pLqZXZEvbZu909QbBZZTlGyM3KbiZm9s0+n2+uEkjSZMTkhfHwIeYhp3US27
XweY5LHamG2SXNZgMOSivxpbw0qkzHN8mT+gHYT052Ed/aDLLpqr7PLNxjjXWF2d
4Q/kpRVurGQHtzr42fMdNYgDAljRgVN2RKYrL9kVEAnaht2B/s1PuzS8v3G94mBd
KHRLuiEv5SCrXWa1FfuBJDNVLA5hf5WID5TFlQevBk11mZAENzNWwDj0YVoUZayU
BfAQMhjfncav1Hx7tycw1y6NBo5hG1JFWpTwit88R+Ilhr7ctBsJ68Os7tbPTpJ7
m02UHEvg9aO+2ZMpsp/hRhkgHyZyvl2BmGD18yJ8BL35kgh4diS5jdPIZ0W6nsKF
j7qno1XnvqKvJRhv67/Ge9FT1mM6CidQKtyKO+WzTzgnKOjWy64KIqlwyZAtPQjO
3+eUeyo/W8a9S2RVWM4yZ4moGPKGEsj0wrHX3diK/E3p6jU9LhangRBnyUC1aI4E
B+q1RFQJAZNdexI/fPqoQWL36ek1f90lCmG0Z3jJe6fZigyNpgXpc9g+X7utpjPk
8SmPUNAzvqEFLGdKnk6vzsI+7/P7GhGopwfMsgbLTqnhSYTaQ00w+noHjlrpjUzW
/hyNP0Xoc6R0E2oW6MfkTbTPe5zgZgUV26j9/Id6dNdUZTm1RMZG74R3JWGkpZYY
wC2uBnM9NTXDMstOEXeC5a2LUDyIHO/lgQwyvmT4XwA1Y9knJdhwa//Wn8uHXd44
+FfTg0ZJl1ePJi5yeG02/Etf1VLIR1B0P1PhkKNYLL+e7qXS+KH5yT3ZouS06Dh1
YLHe8vk5NmT1dtL4vabEq76BUNCSTliY+GbWf2Sg9H+WpxIYYlhVz2kA6dFELF5x
eO1xexfAFD0Fz3Jcsrlv9dMwah/ap/zO+yRRST28bjhTI7pwxl8/yHfUJy/V7d1i
jGt2XYnibL3yGISjz2bgjNeMY+U5sri7rH+uIUE8uUzRqi7nwXpNg1RxbBPmkeCy
Gy4JFlnj2jmOZzjcXxhqzZAwd07f3VpO+0XB8wJ+P8CnY2dmBsSwu877Q9q0ugT6
IxTrBLhXO67QCwJfvqM3XD2lYBR17Cpf29zBViPoMVP2USq9yFrgoHQiyKotj7fe
msz+orIo8oTOdXaAuo4YCw+EEjf2c1YkAMUqXpEt4vmG9PPXrRk8WkurEc9MV40E
RknrNU6xwv5eK+FWLn7cfnPu7SU+9SxE4vuJR1JHbRESw9N9wEoSJ7DXhKSScVGV
hkwG7+4j+XocKg7Mk13g311JkxZt76/+UkLwGfk6FCjfm4LVLjc73hpZJUrQPEvj
a4/k+8ZOaRbjThNQfqXkIqQKUd3R+MgBYB5PuV/kti0pkwuVe4Bf3H8QKIRndUB8
ZYQKEyueZyT4uHl5hK3o7yEGJqc800bz6jVg943mi4CpvrYT5uDQkni/QZ3Mo9pM
N1I7OZ+usjllQdiZbhgxe/wZ4bXBuAKN05V6faYGHVHUJIWk/2K+qeBAzHt32Sds
zG/2qwmU+eNe0TjsFVrNrT6fvWlrhrjbKLW7OWCz5WfYzwIol6t4Ko1+Y72BRqrg
3cEI5cGJzSkJaru54tWBXT5vOsNUGzd8aEvjmqgEleDIfWc7oA7vIqvuaam/t+m+
nbJ0WAojShZCY559IInqPTYNuYMSqbjl90eX2wObpZwcxz83m1KKmAW/vBzzpwa6
X/7FBvw59uZDk9s86+2CMlq/CMQ9DsPA7PqCW//7hzsse91lbx7Ma7IfAkL8i9Cy
Vt0snoCRQo3DUU8AEk1W59JqeKSNWfwTVaojiw0QPzPKgtvVriGNlnkz4LFehxkv
bF6TjxQks8daM+OPgU0YyZ8RKl46NOPNzR99GWWeb8syV3lSEHgoVXgYPPSvA7pw
BQgFlmP0Ipo8isYzt+NEgVvDyKmuJ7jVfqo8amEBOeL93+E4xVepkXrji0KYoF+Q
1P3P187PEBCEMGXfDDzEoBFu0zBDuMv6HkT3RKhQ3EO3vlElEVQfXo/BNz3zCi/I
Ohv94BZtEbaExikNC5iJTkSncIZODpbdUl2hH19rJ/lkEpRTdY6gHPeA4l/268OO
BMw/P2E97OyBbeLtIl6B83Y/Jizs+UGRE0SZ1U2Nxea5UQD8EqD6ubTXx+VJ3KrI
zHDqTWlcuUeM+RS25XroPo8JqCbG0KuSpB6c3pGiUfo5r4fBBD+xaDOv7/dGCprQ
dNisVc2KWCm2tQLD6nsxKEHTq0HJ9WuSSvdWuRIRTA7pZdj0yUZ6FXFGdnKswNgd
PhNPIEtrhp3hvfA/0KpeVR/0b1fyuO0CfEBZ5kiRF28chezAzqhxlLAMvgQ7VwfH
/cXsoitPB4WgHMfaaPreg7ZlStPTyiCT5IzoNV6upGTFGefLKzlJuqoglsnDm6+Y
6kOxaMlmi4lWn85U/RIBNQGdelQkQJQ1nr0CayWWs5zz3bsO3+logAQAdc/j04sr
ImMQkmBXQ41MrHdE93oZw4Q6K9D1L0031iHrixGY+H50zfbC9wRsr90qetip8Nzh
PB6QHeJbJY9Av+iOIjY77IWCcQ6YmmqJoL6fSJ5gKTOHjBRQpJQLRo/OLHXTf//I
8oDSVnxYSgfd96GarcLoPalW7IAPus+HNI0jA2so8iaH3bZVXeJv8krr918Y4XMa
mt+s7sNP0MsWjbX6AFjvccADOj/yhonKOHm0blRH40DjRg6iQaAZ8dT8kGfMLVXD
JiR4aA1GtDfnGzuEs/VNyWYLhLPE95goKfGANspcSWUREAZVXoXib8k9fk25TBix
rEGbMpK2XsIl53+9GuuAY6VrRi7piRej+2uRDNwO1IdMfXBqULvWs0bT+eu+rao5
E5WX/cOUQvf7W3uogVbK8mnZiWo2nVGi6DxlOu9nUutUM7QipD3KhTP6rZRiQ4y9
Hi2aWuKQuBylb6z0HpNYFrEzDRJMbWrCN1hTW634PdyAl007W/7Dmu/mZh8kLbv+
UKIBk9Np7I5T1IAL1fjEc9kebATMjvxP4auMWrKRwxaeyXn3OOB/0UQITnuPv4uZ
rmLGYzS7HnvJdFlfjPci0JKglS9vnvVHz7twisLg04yI7qMkIjDAfTOrvenrdH1W
nKeNi7e+rpl74g3zmtHaPQ79lkDU4KXtzv3t/ZXT/GL1V5lVLoC8t4zMggkIPzKy
mZySySgNyosBvQNrlvwhw7NaZaNE+Hn7N3ISiZHqhQmhHPCfO3hsoPNssSVbS0s5
bO3XDW8XN7XSW+VWQY3TEZ+4t3zM3vi8vRFrwzqeVQEQeazt3gtdZqAGUCZQ877X
fs8vJkkpNke37FSzVmUPA93xw1A77SS5hdzqW5PZvf2H7b1jFxQ6AEP/sNH2YIK+
9naLN5Bi3Utb9aRFzErCoe/Yhi4lFfk31d8xMIcsel1bamK/ROeL0CnbGTxW2Frb
MV7jCK9I8ZUulo55AyTNpFVrUXOQpRulRZE0Z8HTnlDGOmxP9qfTkf7zad4PeRUm
3JTegwFPkbHkPaojZqu/cqOq2mthfsoaWh9wbroP2NnKMq5YgAA4AWT8AhaPh5Py
VvklWRcqHOq920cZ7mKjwNTGh53hBjpJ/49bRX3Sr23O8MZtxH9Z3lYE8gBSrYxd
8g85OxHV+t4sbw96AFPdUYuZT9jnmj46oBrmyuzyBzCYhiPjnvoXCK5BZd4dxl4m
/Hr9j4DbeK2/2n4wRfjY9rJb6bpMHZjNSMk9bwT1dpDahpDFXrT/fgjcmLuj6sBf
muQGDMUG7x4SEBmJ8o9ACoImQs8ZG4YfUmqTemXoVn9PacHaRTjv+CGBtCbCPxud
lhywl54kicRbMoSLD/O0gwJw898Rs0PZhVf4ynsqEBlU3f977lLU2uY2Wk4d3eGR
CuVZWJLbOrMu12AIz+a/eoqpakrwY8HVXQ8BX0j27t658yTI+PW0jmXEmvbU8h1o
0E4ubDRugHv7WbU3tGgQb1JYC2EeyaH3G0b/bUVuX71XkZkE9DPkA9H/gowB4j0k
9X3k6JQFq4tkIQ2UOzliFkKJf8cwRXfc/1jLrCDaxohS+JXB0dIo4CrkguCosRw5
dPs219sLVi2Svr0ScuLbBok8zLh8lydlrN8eQZrTZUM52xPGRTVyC2RRqBto4JAs
wxCDZXyYqvC2BzU2KU2URZaSBgUdGAhVQOXZRIbuc4FUXIcpKKkwanqKl/DMcTQ/
txzCXW9XH1/K5okI6M/WwNppdiOlH6V97BjtyG175Y7JJvwqaPVcI6zJjcEDTKzd
yG309XAqhXgj7+Xs0dxdfx2QnCcvdtyluLDe+HrzdqVcfeScdMP68H50FqVegQn7
5q9jjCnrV/ccG3Bbd7k5glpvXkxPj8Q3KjBXlZSQJEvI8M1VqSLURNnVqrZgo15i
DQ2oUQoNyATwsNn99erGS7E/tSkoCojxAxp84lHiZAuam8WMYEHqow7sXmf9KtG1
RPDquIK7wJ9Imuu99DvDh3WFaz+xIyRwmsqpDAcOLdE4vaRMiprr9alNS3mk2LTC
4KYOvDKRuo6DopC7VpRs1OlQkkeVa5+TFzxVJ4Bd+/XjOA4DIifgtC2ZVEHIayQa
ac00tJx5CoXQHke9Q0Prs9+wJ5LuUUeFiAI43agUaq2zHBY7HJj1x1Z0KaTP7uRP
BmSX4Zi84yqxVkBNljIdycy43qW045vmr06w3qEiGJAHL/VTRsb6D98JqoiuQOt/
cZvrTs1pL0/3110F9GMcl9b1AhyTW82zCECCOvOYTEHgg95/HSnuaUTa5CTrAzo+
2QHKrDR9gj6Fdd0nuqu113nrQPWdRzUZpuWhMGWZaLKRxNfekrjjgYltIBmAvcOo
8dBBCmBdUBMIMslo6ecUAq8ltb/idXULsnc8HikmCD9Wg3XJunk9pZokYUlSe9K4
rRJW06J/Jlc8x6iyTNxOE0RgrVToz2sL0Z32ggA9r0aF8GLUutWl3h3Af+NoYp6R
U/ko83NDlHjBvCPgURVmPlyz3YQi8EhfvRYG6GxEgLFPF1PTlDVZrtIcdIm7e0Fw
smLKTFVam79la6jvlLglerVLIL0Sz3hgzuji4ZCrUfFOESWbFat+0kFftdnBo9NQ
ygFQV/EA9RNUNClsupmCkStxJo7HzpqpvNqMcgiXOsh3UruABcobzrAOyOQjIqmZ
LxMshTHC4H3MhDIdvU65tIQiryUbk71Cba8eaueXtijG6Xy+mlial//NqRRC3CQg
QWErTIrcp3cokiczU2092rx1vJFSHHvln8JVIeFw/hAPiTiNUuPW3zshN43iEyVH
0OmEywgcidP5Hf5q+SljS83LZqoRqIa4YcjMsRWgAHnQ26TPtoHYa7vsURD3jcAU
6EGdxvkBimtASl54U1VRf5hB+Rm+ECNGBphDAI3PYfSy4gft3t5CFe6dYb8rX7U6
GAV1dDofwl1OTBmHSk1DAu3ZO7Cpu5MGAonaIB1qzGkasibXY8Ov85VyPk0U0IOB
UAj0HqK2vv6KXT+L+dbSCO7BSn/bqtBeL54Zh22fM7/1ppySZniqGrD0IeYVmgqs
WsYoDOh9EAsjD/OfMohs9nju9cSK5AdNpIhEEsygdZl3QYR7aAxAKr0QcIyQm8Uf
7b9KnPPqo2pMkHt86AfTlRptwnt7YaGNNYQHQHe0EuvHyy2wEQGjaEaLjMafsGT2
m+cTcSC0IM9egzw+stqSdOqAS8rmVgcj1IeqfvYf2B1GJ9UBfPJyl1w1Rq5Dztvw
EPbaHoTIvkn4PuV6ba1l/PFF9qO/3GMhTlK2rCNf9Sk9iEBeld6QScz4RRJh2pfq
7g3HjJgsvgshcCrcAFXyPQNCToQsuu2LsYo8I5Vc1RDWxZWEuY7kc7yLqa6DI/EU
z1yqaJ+w9SAKSP8atwkGULILaE3YGUCuhUFGQft/J+YP+Zs6orinc4vvRKR5mvXB
F8K90MqUkreqH3ITqZvn4fXJBjl2E8qVGM4yBhKfgzzXXuPN+WTl13J4WGz8pl++
IRu4lcjOcX+Ks0RebNWZyGv8tIV4g/+27xe15mrgE+e5dt7Yy7Qg1pKA4GgAnukP
ekTIOEz8rmLMnjkqSPF0F/XARdtxQayYlLqnLp8VH+yIBbxCav1eKiTcSPK//bB4
1DcpfWQMzRhJpKih5VOQDJfBI05BZEJYAk1g7/wultC0W4E7tA8IudV4aCgL13D9
VwWM9lFGQR3AKGculBr9SLViY3gu2i0MeIK+NVefO5t+518/K1M2oezWel3DJTZ6
xiMrbPE0LthbNQjhsbpU519nUxW3HBKfDZLSxIYjmSFE9tFt55GFjZkV3+YfkI30
b1H/+6gevmcZTQskiOvrf1UxpNifEGi9/xrOY3bhcoVb33wqbZAo1sxpnH4NG/K1
lVbd1nnjoutYQgHgzqbulTBiWR1ielFrhxwKsY0E+3M3KMFRJlt25qUPf1o7KI4q
UlRe+8nCMJnY12DS2CkSkJAyIWsJGv2V0GICQELMz6k4u9HLqQwI8rokQRW/7NvJ
JHIHE66EwBJFA+a3hLD6ZThkp2xWGGio2XW9VEB27hGllKHqNsIGVYB/XUnNSbQ/
GSSIRVtv50X5NlEUWDpd8C5p3Tbupmk5bHSQaT/Kdbha3mKZoMa1ZAQIxb4VWK0b
X2SDHV3gh9Jm45Got6VYtFjHzSNfb/+JOCp4N1iSdNIB3UH1dJurxsI6OISJ6t5c
oVAFVzvtX3Na+sTGtKQKQl2qBz92RtSTpDQg6vOhsqj4ObM2bEGXFxNx9CBNyahW
sNSCtgthiAAJqvOtOVm6qTrqt6us4Wx/nv4/EMOnGueV4x3ar7oKHHbGZRAVZ3yO
8weqxlRra6c5+VhQUK/CPXHqUV5d6hJ8USifLlfeEtYHvnnHi2js7m3ZgFRD7ZIr
Zqd0QrUBlRO7wOxF25FXsjYwnLjvtPVzi7sQBDkRprNpn3HemhoOeh333ge6dq3n
9xAW7KReM0zEB+gKM6v4OK+8UHLLaiYP1uRn9laPdQfw5804Fn4+5Vvl14LtG5Pk
46oGJT53FeIfuUl0dvBRH43ipZ2zDxdnbkXRE7Sv44CvikCgrKCAdaDjDORIPOa1
gAKnpK/vC2ul4aNceMS+HzI2EzigvZJQL45IArROWuLMVA6wkYb860hBqrvzOZ2L
GdadZOkXg/by/aVCEgHWtXjDlcJzK3HuC9kw1JKWo3HPVhk3E9+GW43OatU8uwd9
+01QIfDKvc6oQjWiwI/G8Vii5L/quNiquOrgGUoht9kQhywe5/tbHV/+BwApJZ0f
Bq8UlWSLjgKpReb508zGpIW3GC2QW+G3+QCMVCV4gKmLVrsGOJwW2SMrxlkvDIk5
CEzL+9JVaxRC+XZwInZ4WyM00ox9Paxj0yYn6BKOeRHiirGAePm6QMjEJpxIFTe5
/LwetM6rtPgvHgNDtstlTCoPJclXqNLYRqxfTYqY5n1LEpcd+gezWdInpLjI/Am5
Wj6/4J09xB7ZZlnXygIRncVasvH7+VrhJ6ofuHc6Y0okICgmbHFNzTXZgu3OPbGn
r/yrLyq8N1vGiXrSjHdRjyJx/N4uWeyWTuIbuiTW9TufKzTkxO8sXG5Xyomur4QB
lKKrG95YJUmcaob1D/JWROhJKHz+SngX3FPnSqunxvZbqD1nvWTp2iD6MaT+Gevw
g8zD9SWzFBa00Vq6MVgxuEuTPQWEL9ebbl9PaJU/fy6naC1CIa5+D5Q0XEyR02qn
XouA/b9CzgU+In5/hjDQelbzg1Tuq7iUI1yFPqzGrxJLpU91V4uTJEM3e9Vbi4YO
qCa53aqzSVSPemenu/JejHzyHM69nQbAqO7kjl/CVl+phoxv/T7IMHAyNent7cq8
aK3AU1TcvHzU/ZzICOS+UZEKSAzJoRFQHl24AH8Nou4SuF19qCGrF5mYqCKuL4Hq
y8bbJQJULY4dVt3MFJFLgeXfhKg74Ew/W1QEpcpbS9ww/KCC3tZcFtf6Bct7T/A3
FLdUfqv2PHwXRj0daV/nskL/AEZSADqJs73SeTszYLOvr+OaGILgSoSpoDr/C28E
ULPYd8PRiFaI1CEn9KR25saAIPG0s4c6TOffQc+L0mxRcapqUpcKBxwlz1ftkKmB
GVVc4JmpvlC+jqUiCo3s9YQtWvxk9ku5FxNF/bdFAjAPzDHs0EK2lF3jPVB3cAMQ
lds0EwmAnzvnceP0SbIKwjUHOnI7kMXwIcvvEEgNDBFwGnXMstYtMh7EuoWzPIOc
vBTnY08wXmGYZG6CnyDS/aI7UxI35faUkrA3yRGn3lFtVLYflDFbJKreUdWKiEBH
Z+e/pZvFZBUsSdgwnhKgYgqBq8WMUgYqTXznHxjLML8YzLT/mamiY6OGifGqAfPH
tZo1pjKe0/miyOho9U9asDrxaBGtPClFm2y2eHFXSpE1gCLJZLGF4voQVIah7Zao
/v0wKM9wjyWnRHTyPWbKsqOUgR/mM9R+stH673kVhBctikQ+EoHIf1VgfHZsExVB
7OiV68qBnRgK+QZ3UJNCygw6BGx9vgHg4X5K6WB6lyA5pPKIcypo1dpUJby2g4Bn
+IzCIpbHK4b1T74MajOMxIbiAninNhTEUU+QT185RheGhUqIiCmz6CvPRS8TDTAh
IN1zlqtizTmMGVq1qppXbMUrjflhI1ZZjQY3JcgyTOw7yfoNYk/6qIvlcoUjil7p
HLg21aJglEB5i+iDaXT1Px6mnn1d4xC9gsY4w28UkN91AAc95ktCMH0vh7aHGV/4
6ULHrrl/YwWxHhqxK06H12jG2oY/Tcebhq5faHH8gjfqO2QOiaGpTHjDa8Bye/fp
v5+G6KEdnhDnLNkDMzxFidMBvcg6pKwInmnAGWIwqUYInOZce90+78AETfXTcEfS
JDA5G6MnekIIgeZVySO429hFfKIsd2UpjiLXq4mLLYwUkPXRL5yaVWi8sljOsXnt
9OEJlgJ+ql7vr4JTyd1KqgyCT0xQ19BTlycg1iSxwtnxtBCTRXmCeF4vWWpXVTEL
1xKDECJ9djB8z+QSQCgofA7gjrB9daQUZryfuh1GZwH3IHe7PGPndnC2f5a+PfrY
R4AyZCFdChMEA+/Vmgpi1lsGDDhE7uhWITT4d05g/sB8DkbNrNuFJZ3JrkG8QfQA
wFN8mZibkW/ETfROLrHgiNB13doSvVaDZeV5I0oNa2ZFR1OVXJKQXmYHf3gI2Grl
2+QPtuN7y0eSbMPIZPOuXyQVwhHO6JRokMHqI7cv+oSAN/GrcrqOo5eOapX9Hf2b
tAEte3Pc/WK/F98gToHu1hzvEARRxw8LJsweV0tpKs2FjGh7K1kXKa53F0XXCDd+
mDkH5qXZieTa9upjZhCmFWMSL8ZIme28QCfIE6V1rFzaYUphvBUG9GZ0nQ91TItE
WP3wjCmdLAk7YV0UUhH6yTD8bMtmgEn/nZ5m87GTEHpkdT1dIn4FL/36tJp7vqW9
jqBRaoSE8N3ngNj2XGnCPqRF+hrYjIZdygeFo3vabVDRdFqNHQitk+Z8Qt4+U4xR
NcSF1o9V2OLY9qMsln4Xtfy2Tm8oyGbThlGk9qAhgIFRxHFXsKstSHCdhlRWofmN
wwyw9/G+at+et5i9GA9gzMH4VNhu6ogPGWEhAN0PdmJ30+AZ9MVPM4CYzNR6+d30
EpdRRBeEOqioTK10EaK9ka4JQcgTYLhjXEdKuG/r00n4VzNpt1Y8H7CBIsuw4xs6
E2VBWoIfLxnf2zAJMQYucFWX+JIfsu7iwwcVmCHu9Lfnxjf3LRT7gjkRSc+ltB+Y
E0SkN5KLjR13vY+sdF4q+rBQ3LhbVcFm9l086976oAgAJGg02dpyf4KDXopkuoS/
Cv2eNVrTfbeMLEDokFjqGHSRBDmAFPw8JKFEg0nHxDFQkVmpPl6cAknKHrkpT91A
1KmKQKUDZTzdy9u0Gd8o95d9oR0cw3qzvpFiete1rUI91PFhVB9bop+9ingi176w
iY/QesyZAVdcnMWu20PsOkeGxFLhMZAI5Ec1/mzpgyF4+FHEMb9BpYD0PWQt48XT
SSzMxXyK7CexaXIunsfpt8ug9MuXNpTFH7jXsGblpSX/FR3o6axVOTx9shgdVQcU
XJhj5cuVjfshMGA2He9qC3gx7iBZtw1jJMgP3JaB31iphqdTzF3BiSICV43xePoH
RcDZhSKvBIzeaorYRiJOMVYQV5q8uq4a+1ymzZdT9eIGgvytQDCtZUEUr+heow0X
O5MpAAU+SzqR2g8SFFOuBVwCfbEuGAbWjnIkIY3gl7EGhLdHqC+tH3n+c3Ru4dw+
fXRXozqbPDcEVx6BVyH4lSx+P1X5fPmGJwluwzxwd5CJwBV3RYan7rg2uZCT/MGn
rKDKOZlJG7Ys/vzbDdsQVKZGVqIo0QZfGA82xjNaoRmrNn8tWzeuYhJdZ8fGL0wH
rNKwkDTz+AwAkf8lw4NDSknsLLFfHTbm225oVtaVHMEysBa/2/MFng50g2iMTApy
yUDTJJ0TJuQV3ppSZYlyvxGwvxijxU+iDl39baVjLTJr+n8q0Hxcf9GytutDodmT
JNO5ARoyVRuWivTLdoFG1yCTRyS9AdldX2k3Tn8AF3gs/H7XIXvCupRPYybtOx5u
So8vfhwj9jV4AHbRrnlTVqVWVnmkXh4F1FBPeg2/T2J3Mypa4hqjp+0KOtpfTatp
46Dhsy5awEyzUdDdzVhKw/MqCw/Te07h20KpI9HoFcSNUgQi0c+GnO1KEJ1IZvmh
iuW9emEP7u3BSx6T5LM1yQXyGUj847Z9wLY+3jBeGuUghXKMnkwCqU/cozUHko05
9MgWzeEPEodD1YzOUGU35kxvCxIPDI95GelG/lCh3gwGh34UanHsqVup6tFmtupD
NvnFmfDuXkfNFp5otSg6iygFVtCyYe0q25wwHxkA/zfc25WDHjVXNpNM0Hwnl79k
b/WkguptNkNB+btZBgnDZXXOcbOteAihXpJI1+egG9cGS7Tr0k8uj/xURZbDK4P9
DYw7g8nkimIIySA1Be0gvRVSsPpJnBJ251CTTRkZylgW20yWX0lxrq91Thnk5EhI
S2PQJmtK68aHOtXfTQRD2eilq8LYY/hKfsNcgDjFgEpe19tByuaSQBrDvwL8Plhr
GpdBBvbXaurm2W/HC4AzHsqxXWZc+klchWN9AgvNTKhgQzd3CTkS9bZ7qB0gOngM
g0GWD0qdpo8YO4vrVQobBIKApSqaULqL87xJR3/PlJu+AlBIEMI0d9tD2yQWdCxb
90lYPILM88oJH0gxr6pGYeU7qT/NTFX+gzpRPYepcSh7XHDwbGj+562N4ImrpL4E
xgbb1IV/VMPTv0PjnEx9A5dNKVwDPAbOR1JJASb9WvDfvgGzilo8o6wX9SjPEwmo
vkwiq7MXQLYZl8iV7oLRjNv+cxBFiy82LUYPhVE4VSwRS10iMvDHa+Z/B0aO6ukQ
LplqidYIX99uOGFntfnMmKgeSIvRC9wXEAWvHPa0wnJ4jH//kI9FZ+SDMdzUctUf
Lak29JbghyJTKdxajg4ctBeoFre3vVnujlPatU3WEETHxcnT3SujHyo/rdg4R9Ya
qlOvveeiXMU+oLJCo1VtaBhsMft39qBqv4TYNd5NHLytlmGAWbFRMHuC90Sovf0t
CprWhD2wMxT5U8CPx7qedaZreCQf6IuVQ57jCnAV0C66VYxQ2D4uxdL46kFBoY3R
bpX5cbZ8a9nmIUWmiuPHUjUM+bXq/cBt6JWoIk5t2qNo7h6lTXXqvxNqnX1RaDIl
ZnkLdQxb4uBJR5v2yK+PKhw/htvMgzJYRtUy8MgODX9Di+7W1OWbd58jIO+WIp+I
Y0IiL01l1DBt7SED36FvPRXdix+p5cgjZd9qEalIjyQT/jN5MKWwox9bmJM0xcvN
iABLn9pDyb2wnwl3ykjgludbo4RQM8k/USHpzgN+e98/2ChRI8UfLeWm1x8w9dIm
+mXAqVhw9ctVWtgPJTngBT3wLKGSF7fpDA/K1VXyV3+YGO+aTrfr89R+a8bmXwqX
n0km7DwVMVEMezX9GgCqwI+WhIlqBGynZ0aR9XxiVtbHGJQLhw6gfLsmKaAqylMF
Wzd+IK8kimcPps+mZY7QFvoeUQD2Rv/lLQsmHiUdCV3BOk8qn/bfdnHx5fgmaRF+
MF9dVZtFrbo+x55jJRaTryvKzGl9C076tnEUqZdhG46LdP2L0O48t3ZaIwovyoyp
HIcRnoiAd4tYwy7lUJ7K9YSGn9qOEXMc64PhXJ7kCL/9d+Z1Usy+E5tSzeqLkKF3
tJiA69h1CHI2yD58loVfMCAeCmt4/5eHxDCru2HaglMX6JqzIsg9hsvn5jUM81u2
+nfUazZ2dtHh5Iv0Yl/dAOlKmQtANGZ1cfzOFpK9kUoRtTxPSlTI60Jca0N+ho9b
ZHh9Rb4F+DckQyN/bznIWEsnlv4rOrD9bW9hfut6ufLGfJrWaVmJ2ovnmfJGmEVa
qtNRg6OamfZ/aY66jPqUm3XbIRmvQVkQQnOUioC0pVVd86xRodQ+8Thx1KadL2iW
YbCvF+vHptPegIRONMNY5nK/TmMNEEWQKUQqUKjlbHmC3GG2Qlez3Y2EGV2v96nY
00LEZWyU0CF9A6TtSiG0fk2sAeqRmm3ivkQVYWDxFWJtjIPvT07Q5wYepuHjJEKx
VzAp1ELX8lLXe+S078AmQs7rEYk8zbNJ8/LsQvEJmiP9vbL8NFDXqrBjhL7vfuyM
+7hY+h+IH1lSQlKc2aXvuzt1s1WqaO6+TOQp0D/hW3UupTfUqLpmXcotQr6nAXjr
Ne0AoLccXyKrnmCLzLrwhgoHRJlIGGLxnTxrqynlKXY5pp5d7/pAoBK5jnGhzdO5
Vf4igawIdE9Av47R3LA5tBFf45fYKGK0C1Nruojd5s3If8co+Mle5LnnAqY1DI0c
jMD5K8VtokIy/sYXKsqgF50mJoGOZDg8mdtsApPSQ+L+IZIDDtR9EFOYiISQfqRZ
FdwNlxFCxdKoK9VSYKRUkVoJ5qY/twLh2g/Y5PLlbNA4j4Vjpy3p7EVDPyPTYtF5
sA6rqwFhiVTqZ41S/ZmXKLquN5pdJAAB4HWnIs2Gz3+oq0llEWHT4WCba3lZfsW7
zC2TRDLU3JL1haqlXnLZZnnm9UFYjdb1EA1jW4sNU4HyVKGfAd3vIG6t4w16aCfX
Qo3W1zX4PHjFZ/Yh6rut+Tu3JY+pA5g5zqA6ZCoJceA+bSXH28T2RwUoDvHXsIqp
drLsPOJfnzzpj+4jJCUpb0QFuLKiJucVdbxblf9yfyWrZXBFrwxqI+EeOHTqLIjc
TYvrTpf26TmMEE4pUh1CUaDGfZwPlnzBsclct1EP4b2SD61MiLAhnYkmcsj7vjo1
znEnO04+kIC7OEa/jIMyW7DBFLs6NCNYAqmOXpn4QGq9hvorcsU+guRjHE79DUnJ
FPtf41+tO4tCZHNNxfUT7Edw6b3NpjWvk7H+wt0HX9SWAJ9Kq7P6px8CgIQQJnET
gosB6msBxw7S6SunxRKpm6cEYdfADuhTVTrmpFuJUL7ue9H6wFS5RvZMSxCq+j41
KnnUiAyXEVvwwANqcLZOyDTwCf6G4p/WRex/uX3LhAH3M8Ii6M8wBHG+KNcn1jU0
+EZO8wt6TlJtgqJACP0SDuiHypTgQdkYQ7QSzEbSnlgG3yP+AmA72hopqvva0zay
/t1a4+/cPHw0fk8j5zmmtJ5OCLk6BHypw2Ze1EThh83BT15ZzQ6cfPN7lVOSN4WW
9dcCMtFI1bYt+ZQB/VzambEypNXr8i/olyzGRW4pVloHrf8NAYcm0xJDiiH3tFG1
2u7N6uFYxD5sVG2nzOtXikTurWgsNoly4Jx8pAyjCKN182hP/FdGKd1QMGf6P3J9
V3VZzQdMeWaYSwVI7w7KZKrmUkV3qbKx+4d/BUaXDH7xAlMkhMUDsFKIN70pJpXV
6k6JmUveCKM3+16YQRYvsR0dwFJ8hs93OliQ36zLb413w5v6M0oQWtbvxA+ZnyrC
OZAG60yCB2WGo5+W8NTEo572N1AhYKj0Tm8eNj+xeb5pKi1GTRgTBLCDnIWZdTd7
fcqIKF/efF1QSkchxfDZL2uGvleYsGjCWEBQvr8vrXtPvn5lVh3yKB8ws2srxQfp
HEikwsyzh2jX7gqjg1WLpPUWdCYzOR76bVFWdQsotEQadUYs6E9rdLsoutgpHGAr
UBEvGm92voAPDjyH1Jy95h4PzEmMl9U401Ht0ISso6VB6M3lnGkQHVGNo7vT1Xah
cRAKFrYK1bAM1Y2ysHpxKcpjGGXn3FYDJYX3lszHiNAj7gxO44/ffNyKP2YCjbhK
zfQGPm+Q7chlVR40gpWlD+NINe/faT7vddJ/hvqx6jJvHi7AhTktxYif1I2UrjDY
IuLSmWtUldfI8lRc0A+f4otpxFMcJRmJ7upC1WC7JE2lTE512+BF4y6+CDWpnljv
1KWsc83FsGZBKVl4oXlqZdxtJYFzBgicLDqH0igtE9bnVrXsfiGCmHRk7o6BWznY
yHyfz5WxYV1/g7AyrPYeZF95f99bjqspsftyL04HBW2lpxtO3TTacDkb7aVdckw/
/HYggFgkud5FSJHpPIo+H7MM6Hq//shh80jwYL2U3QVoB+SlSh1MUJA+pC2M5BiJ
E18bXtuEVrikIbYMwhI0agGOxfdjeSQ5BWTTK0HQSNQHRRlm7vuKivBmYzW0DSoL
A8ZQI6sCWx09zOTK6bGa8xC/LA9ieG19Pj/yscTFx7uWz+NoEtSG/S6+kBNsY0do
NwcsPVd+C+zmBrMuFjfeZTxPA8h01RqprNC9Td2VW5ep0amsanjJkZUm7vQayzGU
HvfVFy/Qir+bql1Vbc7t9y4XwEeYSVFesr/tLj7ZQFv+VgMKKt5Z+q6M2YpK6v7n
P1ztAkAebtTW97Zu5eyxP0NouuJ7CU4YCi5x2NlUI6Np/LnLGbwkjvWxks6sq7Yb
jmSTd1x+6XMKt4IPlGzAMWxz7TeQX+LVz7Pfnqb6bobaORCrMQeVSm4Zbb/2/UMc
2nyTjzSk8As7PivhMNAAIL+MkcAsbRlrmjAeq4yj6VEAXqPHx1YBWsB84y9qC8pe
uT/Wmt9JqSRRbA7kzsGcV9QKT+WJR9/valaDTlVkxkxif2kFrLztPH1DBRXWHqw/
kQe82ldzisVRWdaZ3tPfag+kTkjBZmquOwQqXv31bS4kf3DzCrH3lgqaiUICqWc8
8wL8JUloaF+xNTI01/RUq3DlM5OYQ9qp0ne2mEQ8zvKp+KjOYo2hj7UKU1SXthIQ
KGvH+PMaU+unf+N/57ZJltRoR8XZDXo9SjZVMq6g7hb2hRcFTk4U2HqUtlS/2Ko3
MNUy1fRSVCM/5rMT5bpvDuA7FoOWPOVMs4RDtxmJAhR9SLu5yKGxIBAZzNlbKZol
hjVwxq4Z5b2FgmHo+vDWmMvuNMbFcXcDlWkcdvDpofZJ5jEKPC8Nls3frYJ4OcAO
KQGnA2P2GkLaOxMI/4RiQkDAtdml2dVhpjElixV2VBn27YwKHG2daWcQYfleeBs/
WmrBcxu20Q4ar0YE0ySqBJmmCJn3bAv7AP5/s5iQ1dtxVloOqtB8NuakR0VXzqVE
EfNIwbBdmld3QVSwfGB9XuO2tIg6l4oiHW8c7SXliRT+gk7CyybexDVcciWglKUv
zhIq+DoDMcaO0CSM5NSk/wZdbdbPMa4nNB0fKFDr2jXWNWFwSEVcx39uUE/763YW
DM6YpswpD1maiChgfVchNbXEkXmd1xkQIufhXPuYikrowUerEI6fJ+O1SHPoiZJr
yhlFWW4I7qdIv+fzJy8OC/0ugyrIuUqzjNyDBINa/+VMhuQlRlNlD51Cin9CkzCC
UVZhlZf8IulVKnR0PAwY9TcJojy+28RwyDctlSptjpb1KunRcQeqk3Gli/kuPm9+
a7e9sxKEpA4YcsgyD7DdqnnoA+jJClRzhNtTlL9pJTzZBOfdkANj579kOYNSXnw3
Y7iKRn0/JzymHHIxCrH2QGPovz40oBlQw+D/Vh0p98SqweI2pyRHwA/XKEWVz9ko
qKv8bRPvl83jlN3CJy4iQi/2luiq8V2lcg7q55zXYiizqfu/4gGyvXY+HCI1K4/z
Wpuqnge461HPrUyN1vlDwQvIovJwNpKNPB4CXe7FF79qJPb8CXf4y2wKTpKR2V3T
yrQ3IF54lToopdxp2T0SOkl+urVOzsFIcPzOwm17x9FZgy0kWeKrcr+SLFfEBteO
Dh+RWqsJfE26ljS10b0ggd5n3GPRcrzPlSRHYyg40U8ckvvYj5v7UAhrJwilMvzi
1oaeIje/w7zGRJ8VVM1tblT3iUWxWl3yEO8fXZf7FwBtHU51qjWIqbiCn+ot41CZ
i3EQgz4hwrcy/h0p6gBzVds7/AQzZ511V0+2nQTfnOTdwwMRWwVmGIafGsStzXl/
flrUMUbxHdaSS8l3xf44Jm2fpuZeG14Srwt5qtF2bT5lw/n7ZD3QclE2WG6WLUge
apA4Aej9tqnHuIEbNsjHHixOylwppVHe47IXkXhz9sLcqBpw3uPNZJOCeDFK9aRE
cdlqDyL2/kY8dJn2Q46/QuaPXWyd52Jka5NQRcUVrMQU3ZyeXEWWkEnH2hWedftB
sXJ5eaalojZVgunCAAjWd6uNYMU44OPjI0LNJOsaIM7X3Lr8cSnD+bVlQoUpFK1l
NnND5fU8m9M7/2iRWcP0uOSIcUjh65xZtRPDQBj4UnKjgAqmmw1wttyCELt93QeD
dmaIqB6FP2JRjZUyAcCOI6zUb5SQOG0ouhaWp/KRGxpyBrpT0E1oWQmH2oJln5e4
skEtI1eWIufbvhblm1NGPDPrMZhF/gsiiY+tepXYjFUtlfztrBqPnKt6MStd0bvZ
cFMmnXfLD2Db/HJjGbMdN86DGdrphkm+Y8cKIHxqtzKt/pFgO9rqa68bw+G5RPFj
/zwbezQesoGLPK0Xzx6WgrcBMCrB/t75WF3fv7fmP8MGcIJmtIQsWsUOKxzmOqSt
ZKPe2FpAbyqC0gANGIOxAJMBBExPWlN6BiyFO4KTilelZ/Eys0jQjgbWvpj4Bj34
71qY0bLGjruY+W0+Hd7p1F9UUdLbMQRGq3HFGdsbxrepZnUmOCpbNbtQzXwVLHKI
1QrlmEMZtUL381INFmG7yrhigJmWm8WwtjPms0A29K1DeKpfj9zCA/0TxlP04aNc
MS9XBmSaTYfEsm1ltMcLmf/5z3nNl/3xFiKICN8KL0FP6oldDPWy5TjsaqbrnHNt
4PG7bQ1GexPRq8IfFXoOvAYmtGN/QcARM5n3EFjnSawtQ5PnHOss+KNRlcoyQy1q
C/NkVZ8Z48WslsTD+hf36NgC3lTqP2z04B03JniFAOEJB91X0AGBsa7EKy9rOsuX
M57EejygPgSEZCBgttZ6mEoBomI0ph6s2aSa0uAB/dg2/7ulITNRdlQQEDVE1cPP
Q0Bfw2PWCuoBn0Ew3JcYSYWcktI/EMCtfLqSYiro4nNKGa8BiI5SMngTpy06qfZS
jZGaW7r1wnAKF1WkrYJ63XSZiWYuWgXn4jGbahPOkee+xPujJJPCytHyobNf/ZC6
BGIwGLlpM9oFYOZNbKY8zcsL0L7DFgV6RSaMFO4lXBW4HKUtGGz660hDQ5SBlJx9
tj+xluzaY9TO9wokBRTh3uoAHmGvH3Z7Qt75ck3EM56GiPMmYWV7jmUwIV/+ynro
Bws/iUFl0Glofl7fV8dfd+mQ7FIUCswBXhFZDMoMBsyrUzQ7nl8/frHIl16B2K4h
fl1Qnlit/otGr8V+5yjTTQ00fPAtX36UXuhawwM7B4k0vc4KMFGIF8OV+9YdG2lN
mtdPUUE9Wg3VngCiqsq66gO1Fvsn9yBTddqEQbac/jDfrzZhqaLGCXoCi/kOp7dM
6Dckcd/VscE/1ZSoYoK5HO3mz+1ZBS/TWG33ITCesceK4WzMcfzcrt+1zJPdoYAB
Lgnv5hBVGCmClDaApVuQyFVWL9dWjY/wYRcB4NdGP9svcVaw6/GApsH5icQjcif3
Or72sEcyxhBwtxlCnPC8LGO4ygYWftut2Zql3pVCUdlUGU5MNU07UY0EHh6j40uM
+EiuOq02qeaBFqOTwTGZTCQ00VrPR3pTo3Wfqik2TNyYMrlIayOy6tCMyYxjuaVL
UpaBjFWi077d5N6z4C58GKzuapaocFSnBW27sKQmJBZWgF0Y38FFYihQrcVADhQo
VyoV10vU9PAVfF7YTpeRN40jeZU/tDLZ/rH+5q7noZ00o0oajDFc/8fbeweZEUCn
rwebOlCrGMMX2HOvJlourDMSwrdm3qt9jXFFp3OhX1PKrUg8cg1HkvPduyWpLmC8
UTp7onEv4vhh7BCjK94wv6c75kRV2nDgJd9ib77nTalHNHH21M+qkUIskMImi/cr
qaseU+q7KptsXfykvb/WkZrCFAM8iN08FI0Cynlm13Z8lKDBiY+xAiNVcy2Hig3Q
xcbxHAUA0v+8v+1pey2LMilD8J4FjqKBHqtwDbi2PAzZ34ndNPanmJBjN9VCtEjt
oq2QJ4UFxpw6DKumfYP5d8f0RlDcOP11sXANOtCW8nKWJ7a7NzfjvoKZGtmfp8zM
y374KqBWufCQIFGcNCLcksbX9sioZ0Ou/h+kT69zBBvlas18zTcbIOQTmZd2Dqcw
8pz/m/zGEriJLTSuQE1Rr4/CwR1/2fXSj5TIqRe5JBzdBOuF6ghpT3b1F9103doD
X6NXpnnNF5Rktj3eyP9DLAb/BtpnJLvz+R4rBOgKP4GXQRB3tw24wRlQBBh+zKnx
MxiogJWq12CXa3EYVg4YiHxK3VeFEvUnTn5t8/a5EwIFrwIqLh+EUHkUpDUOM619
bbANLoA0TzU4/yD76CVBwwR5y+x6G5hQfCXofYCqhB0ZJ5zaxbgGIoJu88J3eTsZ
G9e42Ou1McWun162BAjgRNNbq2JuxtryifGpbd1sERHuGMSqHdLXytoQ+juwiisM
LUDSNfFo0DZVbOa7hb01ZTWxIcZKROi143HsOKNleL+uomEgfDEkfORKBEuzLPZU
JxKlp9u+WLF3zThNKKimfhvN3966/DfHS7DPAjlADgHyQQdBrLyFJfjPHdw+SK+W
gQcicgWbXYSmqQrUXJRWBmpsb0Nx8yvV9Pr72jhI1oDd9BUr+QyqqMS2iSQ3fitk
Kz5OcDNKIQcjNbRGECe2XXbsxN+nKFElQSG9BhUnDf3dW+fxFQ9x84tDqzj0soae
F4ptN9fbuQaiV7hwq7EHLGQIEaG1kDR3xJ2a7/PAUqgoQ2rTYbqWZUHMHhKesiQ7
WEbgt4uO9mjDL04rCAiy2GKm8IcedCwGNXxWbdvx4kVMz+GunXDbdyOb1F45h5JM
IswkGmjxlfckScxTC/H9u0eBnaCHGVLO6r/SBXUB+ULiUGrwoGR1JgaYYLFVgaQ7
3QRd8VL50xgK7DffKiaEmfuGRoHhx8Y2VDShej3V3EmtPF6vBPA1tmnPzcAlZH35
iZ0a4qZVh7s9uvyVMhUtXjFkuzqZSHS4+duV3uwE/pLpVb4i4ZbWyF4YkNsp1dWa
IXTWKHsOqNGgkBQ7PZzDhWlwGjHVnb0Xrh5mAPiDXB1XIsUulIpyhaudkh/v9JyE
kc9EDn7j4qyJ9DwW0DpZ/gqYMenY49PhwesB/ZpWldvRIm+9xQdMyirJtJtKhJRH
4EMVfUECJYEvqDnT8coTcCjiIp/Zx5B9lTgEynNn1xGGAr5JBKSpyxFGhNIC5qeF
33lslco3+PaPOP54Ijh+xwiGG+zOdvYaN2ezkqxLXmLoURnFXnamsbBmjGJKaq15
ODu06rGfwOIp5jj/chU7eqht4WRDOEa/qxbqsFadEbh59YFrE59DBoRQkLI4SjfZ
M/wGimo5Gi4jcMhI5vNqV5j8lcyAxGYx3Jr/RnJhQK0RnWvf/qUy3ttZghtVgHah
eTMcH62+y/hMZAJQQpl6cZz3EfO8tTa87PXLjw+FI0zYLjtcBCAXnUiRHzdE5bwy
VJpXFvuEKJIo7+d79HNSD+08syTlw2Nv5EVUibiSEy2O84tn+X96gMsl9YorJDuR
UQG5fGxzA5tThKutpxjx98jHT7+h8gj5RuPuxH94I1mKabMonXRjPQOcC5QKIPSd
xJLqyTPanP9GiNzP0nqK624ihmTr6QWugz7hQfHa0XRns4igRNtNDNPZprNilQjj
ExD3PYMVlGRWYcDtGnS94F0BwwihJB4G6fbWm3r+Cpc6IzrkXO0bSsU7lNUiddR3
JMc03RFMmyupNAefbvMPfmJ56JypoXdSacocEGt8SkLLJgkDfDh+WVystIO3hej0
TVme/eSIi7HXs4+cFfO6m2pnU9f8HwsLs7NDSVBtoxgYA/Rpo3mBX+PFyjhH0PS4
n2E1aJ/6drQFAK9S8hI8v0gbaRvz++z6ctcjiqJS4g31vznncTBeQuMhI6gTIJq9
JChHnM/qCErgzPFa5L7rD0Hw8Ifl7aaCPJ7KGefg9eOr9zCP7vNWwrvnW0kICH3I
/eBTbuhzXqBljzHs3D6peVZAyGRuOlclqiURsAM7B4jThuygEtQYCiyqp//1PzsG
/2dZCI1E6C2blnmAd8Lv5kEsNyeehbhXM25C8JBViC934enGaT0GoLkbtrausZ8O
HeHXEaHfMKx208UXDNC+ytnI2t2TIYN2HVEmY2D8HHlGl5iSMw7bufKsCTpm3/MC
GcYCToWHaMGOsgbm/jYF+3q0N61FnEtTEWMJ0+1a+PNi5UYSS+mNSXJmtUOTOT/q
lUwxghyYN7yUlI87kJoY1PIZ9NKrUGwFKtdl/ApHG9sQTiRbP7C8SSpWVdc86e/1
8tGHufmQUJekdUvRbXBurtkC8L4r4J42WoKJRECRBhhCbOoeOEAAQxNHP+/zP3tM
aLDm8j3qGyrZXcN+m8Hi71nhi2m340eFBEZ3dYaN2QEd6DAIuDz2SjYStCQP3PFt
m9pqAcYTlqtBtFfoK/t0NYAEAhup9UDElESJSMC3bEowN36hWF9rMyCMjo3bV3zN
qrG0NQBCkVDn8bw7wLmA2Fgp9ltasToQgToyBFVPAF8hsH16qR/KGU1WGuRamNmx
kNN1VN0D0rMqecQwrysM/SBZNIioXm2vlxdigSb1rVZSIoaI4RVAaFCbzZNmzKC2
mh/0Q21tjhZ5g47BGipM9QBz5PAuKE8UMJOB7BZTwKno6t8fr8nBuzXqdadzxeoF
oujnazflGHragTG+jEbLlMl9FKUN1rAJgfQF9ik8JConBffD54NJFe1XAkHDaCtE
mCezuXZEPrdkDhacmXG++Cbde3Wzqwmvass2GLHqXHC7KXR6I+mX0O+xGrG3zCMA
Dt1Ehq+c6fy8rJft6bGhuLEJDmF8eO77Q/o8REhxjNhpczaL50lJuYLs9kEhQC5u
JkGNagi0LdgP3FCmDS7lOJdRyzuDBCsfeYXgcI7nNIXZNY52Nx0udGDet3L1dK2v
xujHsCB4FXFO0InkV1FyGeuGVtT9/H/z9l8/np7EsPDTR4LW5wTVM5hXE+ESIpiY
kd7dQALy2OGfNmj7h6qLniQSAE+YHccK3e9/sN7YY/tJ1rSLDCjuoVZeTqs7WAxu
O7xSedF4nfAisK+DZztjQ8qmOnyi1vs2qybKpLrQf1f3x3ZDLyuueuogfGXk3PFB
UQlYFGQVtCvYPwPCUYIdEGmj10Hr5ltL6B9FjUpoodKtGHt/Fct4IdxvXe9Ghr3S
CubiD8GbAMBAQQsju0QNJ0kD3cy1hjkCia5rZgOfIaRotZ75eA5JeQRYYituoL2Y
OUI9WOKW15a0w2ezWjipABP3Y3T0ualf17Lx+a+yn2l2phtj6Ny+rVwOptHeiD5J
dPkbo+LGOxzus1xp1+rZ5ziPfRhG0eqymvpNvK57IE768pT4rhl6Jq8vGajtSKf6
cEmss8ek9MWu+KXO3aZH7yi05fMq+h/8xXbfiS1+fDQeT3xx48HiqfCcWq+sTmC8
HgN7AeYryyKm9IN9A3mksrxi6+KDMaNLOUQhHXzVfgphKeQEb8yNaig9vvHpmHDO
mX9FzMHMu76O2NUzQFZtbV6+7H6qzQn2gbKyLh523C3iLcgMQbbAYPo3LTbXwF6G
rbJ2hjEtTj0NE816nGbT7WpGW2sqK4+kJQ9jotgxZlL/zgF4zX+H2ppN5icaQ9Pg
2lvMFlt3+xbIPXY2fKHgpIO4K51vWHH+4TU0LNyo3Eb0nepB/YAPq2JzJ8wccqZI
mLxwCUjD9fMSqgPIMrW8U+U2Rlk7hkleQlqk7JZ5wO4H8zOPcWAySD+OV/GqeXMi
4LG+QsLKkc7mLSsEURuRabY+fitxrFRwFuAoAVlNPmXn/E7z5Z3WsE9Tf/ZWz+3p
2BrGYQGJnOrDqstxFt50CLOKBd5ImClodw+XUPvz1bJal/dVPWNXqenehryZuUGx
5lqovsbx5H4/LQZd3FjQO/2xq80jTzBPLGJO1OYHi9h3ymKYdoGHnDPxErtsS/GD
JTJnLr0xeFQZtmEfaOAPWor1H/PS5iiJM6bAmnJ7/GDGPRaaW/wRkoQ7UjUdpvO2
NiXdQJxYPe4sfzNValgw9vENR9K/qBHDv2fz/xbFig9WbC5thRr2vN3bVQEJUwvk
t5Ltg5bdQeAIsomPn2LcwwOwurCVkKVH7e/awBP1XslVBSb5vzV2NYjVOkKx27+j
6+k6pzCijRbiSk0dwocgyBJcv7iffSYBZ2A/w8aUFBOnKg1zzy7cmkpP5ceJff7Y
ouk2d93KPtK3p62LmIlXskOZl1CRnlKquzM++f6Wp7okMGxLRNVT8K20rHMiIyQ8
pU0uN31O/eBwKaXd3GFnPFoVwMV83LR86nNlmYQ0rAULLatV4PC3OpTR6KIEVElS
ttL2sygzSaZlVgwb0zhVWoIsCxqRNKqgFYWul46Sto1up0z3AI+dXIvX7I95jTrd
ejSO01yfZGYsX0VBKMd6cZhOwm65elolGCGPC97SvzFPJuSUmqHodtXZb6lv+GS4
poDxWi85TvMo+VmIGQ11XmVBiCGTppOfX3acDZ5O6euri0DjBDeCvTLYryazk5gU
hAwV1Z3COcyXttXrA5SKdJdxOd5gJqMvvIb19Y72HRv+/mhELg39+BTLTxHuUg73
piWWlXywOMOaKQhpbEalKcq0xubZUo88cKm0BEJVS4vq55JPGIVy88ktZygDYZ04
/fhC36d+qjXlkalSs2gvhRlW1Sy24QMS++lbj1zMBARkYFaS+nV/AAGLaAB/q5Bi
cF5efaKzsSWt4dEr2c+K/oUiL2s6+lWHUwC4bLfljjLZuTLUW8DlxjuY9JP65ycL
9fVBaTlqU+wJzZ72EYuALGCJbjUuP7Md/Xvzy5D8vaIml1B6uZnbvqhAXqeRASIC
6m34vQWx3DWjByYFtywjCSZfRW/qdEEKg3pKFsx91wk/khGvt8oFnElgEUtkHc+K
vYKOhlsl6AYhIZKQNa04HZ9bHaarTiek5bq4RSHFnsJAvvosKnYjznvDkG24dWtk
ZavO5rUG138RriGP9FH9hBa5o0I9EZ1qF0nqsmNpkpDsJn12edLfKjSMlumKFDp4
aFRT+vctFiXvggarY0F9sxbtxzOYeTnjry7vmnVO7AKda/TAq6Od2LQNE3ryvpqy
/azBXTN2BD4sM3QgHkhyKtpR3XETxCFaxS5GjRd5UG5FlMzKvbo5QHEFS6iynOcz
VMMHkJ2SgsS3s5fQE+DMwoX66mw4128QCISfFgv2Q+dZY3AefX+6KBGouq8paQwk
fVD8Uq89jRn0oSG7rcKzk38wbKtspDMKoknWzdxS66+Hpprw7TORiUw1NrdoBdGl
jXu1gGhCpaoQxQf7tWP+hT2FSbvJcqb0fkzxzZsHvahCVUij6Cn9BZt48h0RbGKm
6uPDQ7FKjLxKo0vnFLlXt7E430/aBkM6C58KSPFrPIqRFiGWP5NKpf8TQskoIH3c
R+zHze1Thi0++wvXoUn7eH8RecGNaUJDwMWR/uBHyG5KSHB/Y1nQCVFIp2s6dCC2
G0B/O5vu1FFmozHPvnI+f/RaDxtsdAd/gXegqhZKKN+LMky5hwHSpbGkZE6zwYmv
EtDVTB3xoTiVUUP9VSq+LoS0rIQtsrMnGVYAuGpMnK6wZNf0AJEfx5fmmRuvgIVs
Ruz/ypAxnJ9AADy6ultmlfYtjotfAEj/A+h1WQ8ZAhaKb+hiKUdGZrVbO3Ch5V1O
Fy1IYZCIHYzmpzut7RMjaABNjrlB0UiICRfMj+/BLVWsm5UCnPBMNQ5p3ETfl5sY
+uGpGEXYzd6mnTeVHJ4zkcxLwrHzDFpcC1yeji0Bsn/dN0sRTZeX0Asdb9nKx8ok
etsg80fbRvigjGPdS15/iBEgdiipHdeSMEdAFURcels6X5t6RmEXoQ50XpwkRg6H
o4ZPN8UghfaaSuw16jPlYYUxapG6NCuX60mNZfxbnYd9FMpocaAz0WViQJjfhkz8
1pQ+9wSmCyeDUhseYGGeZ/kLjaYMJoiPyFcgG9ph+xHnbVF02rqKZyfeyqO0Hjcv
wrEb9gvwqENSGpet5M8tUKp2Gp9lI0BUXlGgrQgm3+lplERLnSHjr4KhE/5hhljc
pVXEE9YR+UsSsiyolq0pi+lbkmkQDsBpZI4RmzVI8seKLbvqZ4kGmgz5yU6PTZcy
3k2kDrLavz4S8JbvdziouSDOxu7jVTWE2JHc7L4Iu4y+eOsxiYEPjGMTPxDZ0Wo6
AjIV4184LiinFVvLbwX541rdo7XJvT7HOvPbBKbHDvG06zeL5nCLdOFN5VZy2jk6
dGJqAsgc+/QkD5Vnq3UdcmvJmrbJP1zVjqC94fR5WNj20pSQlJEgoWleIrhz908U
B52X1AfEv6wxwxjeX02CtuGb7WxtzN9u0nPX4SzWGhhEBr37zEdyKGHDWnCOjlmd
WirJ9e8howsf32CQn8L0FH+uyvw/romLsFs2K6EwmiepfmawqFvl8f9fRcl32b1g
lYVew67kA8sRYQDPyE5qpAPvVnp1t8vToj2KyPdgqUax9DLV0ySZW6hJ25+xNrja
u+85kTox4z98kGvmN8yOHDThAdmvuBh9M+WfJ9RHNhJHNd/eFJa874MJZnmyBzvA
rQc5Pu47Biz038YR9YYXOSEa/03Op7iCxJVgaRLLC1n/3zv2737FmC629W8ckY+C
0lx9tvSFzeTtojwv9ATWpZGc8MImG4G6h8T0JBFg9UvjRJ2fFTKsNn7XlL9ckgvc
v/6O6+Wg1iNi258yVr+CGrE1O0nHyGF24R4m3EM2UaZ2YsioE88UkKF2CslYxSfR
VS/ftp0MiRae+/ryrYGMW4lt2QiGLIkrhFVgLfs/YQmEQCJXzbW8uuCdaKYEieHX
7nDKILdmaEXNc5Sv4bzf5TsXOfNDCC3FxRlHCU9VXe9yJYWR1Y9Hlx/roxXCHwbS
fU4HqVw9h30nRXKjvmIG1uF7Oe6Y+9PP4+DxWVs1n+W6AQn/esnbZZ7A4qU5iAIu
ZzWf0lSUHICgrVo7ZUvFJkzgzz594lhGBf6lgKhBe7GIzb/OZDtAnFlV50li4uPi
ZWq9zw72n83iVcDUdPW/Pl9lHA7AeyXV+GVKLR5wfPwBnJMad6PMmaLzcByttPWC
SBVwUWvimPxbhb7xs7ZRyY2lArLldCFT7RNlCK/RNlyU3wzWBlYCl0qUOEYYYBcB
Jr4Bf4yelzOvEq1GRqv7q+bq+i6gVLuPD2pzwXKvOGB3ByxsDzRxaKGkF4e6zNf6
oND405/SWy0PXhYILkDDQ/dNjbqrfr1W4ssikpi3fK2RgOAkJkMiS5GAg3vZs9zH
9/6zEZz7rilO9miBDJ5hCHNTspC2Y2FISSVM5SuxkxqQb4uPdE875rn9Ipv2no92
PEsU2ztzwPJ05m5PtK+4XHktJFle+yydyE2lxIGcB69QvNdUyc9/lhk8kmC34rp2
nrtVW8/Z3TvRh/zxOe1Wc/ERvdiRVxM765vhVk6N7KcPoUK071ePXcZ1OY3SidTp
y1RnaQLFVqF40UWsxSVPVdmKvQrhv4NKcUVBwsispSrs1++YkFPq9hntVBgOswi8
8WPjyfYtPNTybr/MOoAeA5WR0A70QhI3Ai5gxOBmZjOe/W12YOwwq9kDUzE2Ei90
hfhjswaJ8ik+FZCAaKdKc3uNtP//e2z/ZXzbRgmJWBbOiUryETArWBeREh6w/3OG
R2cETt7I7bMiGmyKheb5hslPNupBgq49Gh7emQ25aSJDxSSgO30ZBEarDQPvSGLK
UJjnL+oHuRbB/6GbWN8kQnbbB80JggV+RZwiNEvAlly6jDCLeR4yoAItpw3tdE6H
i9dmv8BF5j4TGJ/X8CHzVv2XyT6qfWLgeMZ5y30SHwZO9YzrZ3XzsYTjNXSxQQ/z
UvXi9hn7Nvb15aWiWmk6UeDHb6S4sWU8nEtmXQpDWdBYpzV8eTuEsNoPsB3VDjbc
LqkesCc/Vy9OcODA6yAVFAaqT8CPchm8srggkQZlBYfvt7s5WPMAdqRhWyjL/NP9
ni7620j37beLS1xKoKG50orX6yjWF55K801KKgjXMuiCliQgCCvEWdLFL9q65TMg
6nI4f5NVxWKKvhm2IRSU+s5tol22iA/RIbpc+yKwI4AaMQs3SJcFUPjQp1GaXCJZ
y1auSg8Zc7qr3zPOr6zrNRstLHC1IfsATJzuH5sExi+3xssSHAyOVToo/3Eel6yl
9TkyWG8xhs0emAhpYK9YRahJx3gQyv0+yRAZQFO+S56YrAX/owm3X1SxmCjPW6VY
aJ2joPEY+/eq8Dlmv0/3XnzV015i/qWJNuZJSUANQFkfQxTJqUi4C5nopZKifrfS
DeTOPyxmuQkTTXbqh8PXET64Yx1X22wqlYXSc8PNMe0FpmZzq6R+rHBMtSs/Hith
rtfGOV/aO+01xk+AM+smRCY6QrC6Sep+ci8BgQKcxMnqTqKaZqqK9s0EzIJFbqoL
9v/IJMCk8/U82ULGXhs9Q/x7S1H7d53fuM03XgSo5cQRG9UsSeCHCYSjQLOovotc
Iho9JJRVSd4oZG82Awhc992sHJ7uW+en8UGhO06kRys5TMnBqsSuOfubDkGcDR0O
IYJ4Je6YjgXRrW76cxJC8VACQlauVApsFE7y13YAydMCIQ22eJ9iW6Eji/4m9Q+9
GF+nyHb30M22Wo+UolCOWesq9buRCm7E2jvIjjPQR0XHJUqqvi5ijctjYQs2c+BC
Jio49V99s/sQ/lUVpTKfcka+qMZnIt97uuvcjYqtGV8eUoV8FBDFhuFinNRGLl3O
c6xjQmOzl7DZzrhpeaX2N7mlVJYh4dkL23NuFOckbTGnpj85QkE35gODMq5TFoFh
9qtK+2rcbZ/TNR2u478+ztOnDVjdUCDDnDrv9DP4la3qSPHmKP5tHbqZ4+8mcj4j
KBskxOIPV2xjnNAfsAVw2EiyXgafu6bPV+8Z0Sg6tyqAOIl7lva4wJx3Vh4dGbK7
mrZpbgJfGnRKukxDORJJZ7BgOSAAenGzVRaugVFFyiwSQXvYZ8O/UNF020a8d3bX
yZS6zXE6xEdo3mjq23Z8L7OUz0nxlmtHg/DDGoQJVanayQ0QhhejH7oOnMZdN8Q+
Wkxzt/zVRDpWNZVBuPFsm4hzPHV0ZPPrwbHGeGYRS6dVWLHNc2+a9ySQSfQpHSR/
hdIE8j7KeLuzpQYU9+sCoS8IkzeRj3nSObKndq2OxbATyl8z72uDG3CWWR33oA1W
CuQBqMK8qnpfIntQDGm7Ae5eR8Y/FXXhNq2Ioff0JQxcvU/p4xuX8gnFY+kOWmWp
sJ2iuTZGrWvncTTNdYB/KeDNwGlN6mrn9BMaqGbSwvVg07pUGcqT3WaSw/84o3nw
iguYIQb85yW4x8CBn5mMJqTwnJmTasBbiJaDsxWJpfzZzWKEpQIWuXI3W8ywWi8B
UIM+CMpHWtZCTsS0Kw1za66OKtX3kXostStpuhr4UA64KLfR2lrhZ/scftJm6ChT
9Ifc7+ZfE2J257IITmx7qyN57/3VHPmUHVvOQm1SlbVyYO1rLfnB8uptjur4yKRV
aCOe/t6+qQNw1Is5uLu8zuiprJD+xuKGvqF/SQPvChoNPAu3c3PmtZ5OHsltsdyD
XkhEhWT29xaUiZvx8RpbSCVvPOrunsIPLj0ozxMigqI5pzDBB3p6RC0TRChEtjeO
0aqkHFvOt/eDDaEkVqQF68fKs3BHG9rmDuYU6a1Ntd4dBWg2oayoDY1LPcVAtIX7
wdsOl4CIRgyUVOMHlA5F5nRT6dF1s7MGis39wzCbFVwSU16EkQ8oer6gq7ioo66C
g/Ruc/A7dNVWe7Y12viI/2YBrqK4mpK8iUjtNYn+LQmM/ATdwh2iSmaMuOVTZssk
JYX4gIuIlywTBd0S/52z5dosB/SMbdRDbZsjBRXuzzVivscuqw2mU6AmznblLbd7
eqn3CcA7aLWlDL1e5GleHgpvDgF2RYh2R3M5mf1gXqmeMkL2SHJxgzUEJ9fx24BX
Sl5P8NnbTzPv6BaPIHh2lVi4BAQqQkrXj3Dg+lf96BkFOgLQQoUM0/gxrguhJ1Q8
wAI8xq+eNo+0PP3yTpx1eaCp3137TfFLprDO8T7ksLYYH4DFwrXr27aXCjuo4xqb
mNjOWORHFi6XZbnUWYjVFTKEPxmxUEWKr5txmzRbgXVRxxPaWbsZIveucC0J64WL
ujUF8NIpAEF4uIdnRxOuraiXNwcDkGC8mOmnTxqRBIHpf1AgROcgLq+fZKRDOaFw
9BwKjixvdw9kyEP+3JXDVvzVa/dkeQnjH6DcknUV/Rq4zT6dl2qKGiPaj7LHDyuE
yQYMXPM9d2B5HgylA94cwCoIEuwGgzsbN+URvFM8H9UNS2q1TAoQdN+b3WR0ubmZ
c7xNL3cct1XbhKCCKdSH8JtC2+/OnQ/tTBB6ZpNZXHy+Y6nNiwhWwEAJvjZoD7Q6
m4R3cmK5TpwPjr2kgBcAbr1EamsnotTecwxhdwkJ6DvTUkQvobaGFSEvlgyYxAJG
Chzx2jkH8BUT+3uCSnosNAx9q9BXDsYXUM04syUdy0dcOHBXYJ4zAHAwbGXqKhiF
oAlDtOr0FfvXjZetJ88fsGj6xJqb6GUp9IMceB74UkqMXLinQbtgYysGbcZWdk6A
bDxGwkKwk0zZDpFAsKPEkokwddfZt36Xima1Crupr+sWBh73Jf/YMOOaYoGUa2++
8UXxvyIXm/T9wZ7sOd3S7eJf3bgrqFERHPdcBYWiYpj3GwxqI10eb78legteUgHE
VcZsNF9FhyOvNGXXGrd7UU/am+o3oO96xirv8Jl/mIRu0Q1FPUN1FFHp3Ov7kXfV
TsGWyz9AO+E7L8iat2Wcz9ohUOEw8wW5iq0xURsnKezgewlUpcNrbGpfrsR8OlBU
CgPWZI3cUbWJG3eViuOOXhG7CtezuX37PCWCDC/QNSqYJVPC5hJioRulUuECm3h3
VuNpl2hUZLwPDjXfSt1xd6G56SkvTftFM7oNLi5ZYp8r2IT2LE5eu0WC265+uivi
mzS+wHjb8AHibn9b2odkePD74rpBZWyqOidLYcGUf1AtBoYA3dIolmNST2/N6r+i
+j71ZKuay+E1rC+9eCQxmjGiaUV7/LkfzU1AVlC9BzQFofIUhmM8ImaeKAimVpuT
d8KvAi4XZjwjEtbwkUwm5lccXjCjNJ65LbCQ+GDqO5DmdFrIdlzQFBIRCwjILcGd
pjyLUWiyCwO1XEu9kXiq28/r07e8qDFe00v5r4juB5qkVWyvu7y5KeZUUJxPVSur
Rd/deZdZdvxI0yNoRbqR+jxnylRJpx/QskcUQpWulhV/KlAagC6eY8laJ3d0ec6C
ivjq873NxuFX8Mhs2XfWcOpQpytBuQgZ5nRdPvr3iSPA0JtYgfnb/ZxnZUxAeTwG
zZ4xjHL6TBFAiYcGMw/GaTlDJZ7gNJovpu5HgtM4XCtBor3Y1UpTU+gp/BK2OX4C
DYW+fjQv7t5Ha6zHCUpKnKr8wi/INm54sSfSg+lBxsgn+UuA+i8vXj/9ErGpUPR6
DqRQPmvpRz/Ap9jjsAhp5wDrCF+UbqLqCpa92oCZN03NKVwQgCTn1tTrBJ8rPK+w
DxLCuBDvVZ5bOUu6/ow5J4AcIXEO3989kVMQmWAPyLD4LE2RHbtxq7P8Vvefvc1a
jYPQgMnfZKQ5tkHSO55gAnZAUY9nhcLmJ08br4fVtfaaq/OTROpW69QZD5/B9SLl
SXBBEGBNRd8E8c5yyrRkiIUljGEVSvgHOdoiz6qLYYw+/qtFXYwdvP8tl7bbvEu6
CAWUNI9xNAiBxXGvnd3zzb63rGgL8zUZ5Cx/MONRsmkDuO9sIKNLVcAMrLGw5ySI
cRf+J2TIwccAEtJkRT+8zPbBUuRVijSTdSiJxonXlo1d0w+Kbhwz5r3gOBr+27W8
kDXPHUNYQDGfTk4WdxM7kjCkWz1oLYzVNKWg/NC/FmBkLWdzPA0RcAv2vGgcIUls
uY0Ajem+Tbr/zgs1bXhnnp00CxHpsxL85/Qm4QBBFElV9siDxLhwyKxE77aRHEYC
7vgAifdMlNqByHx0iUa+aeEmoJkzsvbQg/vWsIx55iXm0pHE8jk/pIjF4MEO4U4c
4bdNeV5/t6mfSO16sUgYd+FifXZTjSBREd804R9q6CBQ4Qlln+rAjUM5dRGcoATG
qnWf3KoOK/a7srtN5CGnKQ1V89DPeBPxnk+AGPcJhn+mZslWkQOSg22BkBGGo5M3
C9OGCdOr0qKxQtke0tw1xmM1FV+78n42UUQU5scPVMElgfkikM+WYruBe2+xgc1I
TObHxGE0DUq7qnrhLaDKbasAuyoBvB1aGhYRAVxlFjGsx7gyDQV7vb/MfjusnrtP
y6NLDLTJsOGOdtU8nBml3hDzQUuETc57CakIbAYoyJQOBkKG/El5tsmfgSuur+lH
3HpPI7wBaVC4M1FuiERaHX+n3yDgTZb7rxjbqk5hWAnvJeI2mJdnsWK5xYOzSyC2
xsmC9jhAXOWJ9jWAjxzdwDveDZsr7eIheDOMhJYjaWKzgTAn6MCvMkZwHUHUBOqh
FYLIbI8/Ufx3XMHBpm/VLso4kjvuR/1DP+u6Oi+a8I6W2EnS14hkIshfNVuby81O
sgrk0xuoUa9ozHv2zpObJPFiHnpd5Ma+Dof5+dEnYB3dp11hq/o50WEtlaW712aZ
9GUuEzXdW5I5syJxxdIS43LFrHK3IVLhfHdL1IJE2+wYEOxU6JphSWLOObyKiooJ
l8gXPgIW+00rloU30AXCc2uTRdSTF9E7n0OC/cHpfifNSgx15F68OiGHk93YYEyu
Cjiy/NYqESoQDiU+yRxddPqWrIkGWlNdzQ+oms1TlU5TemrUrvCMn8yd3OibRxuN
nrPLF/PVysUSOzHR6DBHTpnoWfdrwANqAzIa92eB15V/soJVusUtM6ea3wGMxk7c
H6wymB9aauW/+K9Z/onS29S0+mVO1ez4djKjfQ5dzsyJLfniT99VOqGyt/4xu0oX
sgt2nW84DzP5DwtsDgeOmGwqC1JPENlSYuqoAlDFLfrAQbGKmiD0ME5Mlb/UUmt/
x6csGEOlrXXAvS5WyUJacChBa1YvChmfLqrLhpkf7Dv+z/wpWfik3Wx35pWLaLgJ
dSA1kCBLJIUNZHgXGc9fQLxFzBePN7pl1GI+uiJJuga/40rc3HujmY77uBgmz8Cd
ZksTCPGmEVRadxbPb7EP3J2YMZjqrJ7yODu0KO9hYtXd19Ahl6XHPU/4I+GyXcg1
QXa2w4fpMRGddy4VEEcixDQBB53Dxwzi0g0+8Py8wob8Jo9onW9GiTscgVHoA4rU
PNUjiHJM0HIFjFoW1nhXgr9Y6BRLbg2NhL/dExPSjkTGsLLredBOtEJzYJjv4TYV
ff892FvmZfM+snhvV66vRr2OXGfRVpwYED0An2ddC3u4TFHfolCVeGQfMPpxlA1d
2oz26ZNt89R2iCFrjki8XmPNcA2N8jjcFhYwz7v6kbP36VJy7CeOYjBDkrfL219y
FC0ePjqYht/jOooUrqLlnlg44QuuKcqgzYBLtyiIkayfFtjmxU8Ufdzoyq9c4zXT
LzxxwlNDM6aRmou919LDMRulEOrs4/Z6Ttm8dErI0nCMUQDsa1b0fXd4ifqYLipz
Tc+TtYM/9TmqTG5xLurVaxHxh2aOh26jIKi0UqqRn9s7VoFNmGedUloAjQX7pLzY
VVFHsv5AQq1j7W/tttp1zOXRABWTg/5KcteMnTM8rpePDWn32m6PpMIejmgmNEJA
7ynfpXKKDQrEdpTQ3TbTBvwkZEyVaeUGlq8yg3hhU1e8tAJv5GkK+I3VeO2djw/g
0PXTIvoDlsHq2w1e1SbYxbW9WZOTUV2o7Y76sPQz6fmcP+YcxzKd6g0//U0BHC4+
iK5VbMR/S4pSKF+rj4+mUrCOgGlD/qipAGAAawolYBgBbcs+YFbct8tOaAXZS36z
lqiRWWudYZo4iZI1D2YwOnZ/xtm/az6LyucxJwz/S2xBDPE/3XjN5hBe6LcI4LAp
rxTYS7MCSUKmi5Vr1qI604ZTnZw8Fx86DfTUKunQWMQkAs3fRN5YTHtzaues86uY
I6nVQRyiIqSXwchOf3EPIwm1wpbglSuwhWu/oCpKDXB0M3CgPwia0YoP342x+NhW
5h+zGH5ExhMogrfRf/YiKXcLyewRpvPetjhkmqt4MVjput16GvGFiKX1BOygKW2k
MZlklJjbCNcgxVbOISGTqG/yjVKptPl0sFaaHwhwX5eDLS3xgsfrWuUBtuxvZfIj
UudEZ5eFT+hWwujnDB6ayMnMGlQbjWwl8luaPEY1c5WrAbQtJTLsmJQHdGt4Aj+Z
+tHHBQApESYECZQf5z5HRZFrsVfNQpidt+B7MaSeNg6hZSJw+mrA/gD3SO5c3zFx
D7VxsxM+vwjY5eCE/dBkMZGn4NOu1AnvZz+kGYrkCrjuZlZx2bzMQE2ncOWlUeo1
GEPzft+ZpebLAnTVE6PdPl7jmCSqYHtqHxMc3Yx3zNE4cc9sXoBxl5yttDfIr1Qz
p16tabZXCN0wjDymaiH+PNhlSD6d03wiKcYk4xr2iNHbtBOijcFKs6k9genUiEjD
gpmyn6RGR5zK0nZSHIyF290GL6TQLFhmtWDMS++usukeE3Jl/RV/mtVKhQcYysk/
sFvYin/83Q41V8Ybi9uK3MRWiYEUpDPcuCr2wtIxahWWw4LAcirn7V6Uss/1Weu9
eI/FWk/R0yp//7JpyQ5SHnXKKXA1wjZtzOTbckVWfbUrpqRiL21J+LH7Qx66vf6q
DROPVhRTW8pIFrdViDtYA6NL5e5iUDuQ/tRu4ihmmwhCk+nZ7EturcgNO2jnIsfz
xQJqJWtNH7WfHx4sVXV3svBSuQVAu56ESSIz8ph1ZDNJPCQgeA/LhXkBoUpv5FdN
sccD0w7fQjZZQ72MIag7Z9BaalrpsZkzOjVNBFG30vVzboOzm9gjsNu+1f71Dwl6
dnSzj9vp8LC3BEJGQuKt6C2ke5PxiLs6JNukyJRvy3T/L9tJNWXrufcmf8RpOIzN
KXCD+MAIV00F3l/1xqdVST4zUMB3X4SQmdNUYH8pSU+MmkKuqiX7cTUg3kF8bKF9
FwjZuAhmn53k9He9ltrEY8nCnmbPOIyxBYIemp1tWCqCnQquPk19uoDq3Y5cb525
JBaVZM8L/ZrO/kP2t7Ihq816TZqkKJvZZXeDIegm/70uFrJicHqqUgvWBNeWk/W8
NYG9lVuFms3PMBfEqxqoWe3/TPw3xOH51GBl7djcVcok4TJMBFYCfRUbQ/7KtnLW
nDX6w1PczBX0LTUFe4Zherl+OI/sS0t13Ylb1vYvTKFFlz9SUv7o/411A3oYIg5a
0sP8k7HjJBx4bI0UDdFZJvcC9GWnODRiLnoyywKysz4eD1zQoGMbIsPbdpPiqsO2
7inkneUYsFYcBEI0OjAh28NK1M2f9yLaH0Dn/U0O9VgNJv+iERh+tlIco8G8tn8R
uQ8yaELuhwoBFCAzCsHZsRPUBr1s0LlVXExeLcouZwtvd7vto5jyvwOgk0MyZyXW
NSVRa8gBPlB2MKOMW1GB2tADZ0X27KesOb558ipZIkDoQ41PcciroH/yWUebSatn
dYB0mehOUdTlMAzuSVTI9ODtYwvSkS1oANI2BLkO7GFxghZ4Tf8uVIXP+3jzFnH+
KW3ba9QcreRP5NgAI2aBqhTdY9Of+Ptpj2Zl4S6ghGnoKCMlNc4gKy8iJl+RB48K
g4FJThKcCMQV0rTi3za18zr4rtx+tLpEz6j6p8P2Crq8MD3uOECZ7Xm8SJkg5rIh
3ORyGkIw8m3O8tpvnaaZK8ghO1aMRFFw5MT6FZTp0mfMfDXPIraxlHJZBl/kMYvn
GQAiicLAFp6ur+D1qMixMUpacHyZ4NsnBwwFsq/LdgZFkfBg2+e3yR5EC6vKNXvL
8MSEkULsrIpQKXgp5Xg0fPfwEucMp1rTzTXfovBs4tNRlfuYUUXkDpTNlOQOGF92
K3num28IgJ7XCMcxN9iF50EfQPyojkQAUbraTVIwwHwI8i2tdqzfTvZ0UbqgErh5
/N7tlpIXY7tMXGky9JHfXNf85Tjn4A6HJlUEQENAm8daPO6lqWiSSheRRQa4Xj0r
dze+rUGFIaWh9uTaH//Hy9MyIU4fsyCHpHle5txY0ABT0+v7XYf/pHQTRRlxwVJH
XH0KZbRTYlQKWcdzUWKWyJCdWg8YWnM1P6yXf/cRWhqa229W0/+MQ68qU17Jgi3W
ZNqiANrd2FQANSTRlLJll3fRnQDDaNXOyqgUnapvAJvkrh8w8nD9amo1zyNMHTFG
78nJnomrNuuA9SUKGvAcabWfZeBHDRBhsTm8Urzgv2Wx0YNsFR6wRrMgaEXhkMDD
AFlVV4uPjRK6dsMYI17AnMzYCRpisRFbPJLKLZLqR6CYFHjJg0XxFSDmNh0XZe6I
WfpU4GsE4DTjYxtTV1nyv8ZEx8BzN6cXeVR3HpyxbvRD4iy1YG+e1FoLu/lWU3GN
U28KTWQxjd3QHbJoXXcRQg2xWu1GUi5F/2E8K5J2YnVH2H3EdccjzuRgP/RZHbn4
oWuq1DzdsAo4i9xUL/26F/1raMz3GzIxXnqkJvDc8Br2kN7UNLj+jR/OSaR8yJdw
yImBHTQnSoQT7yezMw14ZW+WFRwCAxno1wa75rrQgJ6A59+QKczT3A7f+w2a6nhu
MRHVqQJGXARKFeA8UyWGbYejrHOT6HLXF6Av8BdgTaI13GshDLCBtXs43kX10RbV
Sphfpw/A+lzDKbRslrNJWi3Idb4/aq4ReXyepVaO7bIwTvJsSINav1kw9qOLYVF4
Iq5FvVWaByOUUSaEkTR6pLoH4STsnKIGlP/ypkb+d6wGfF+3mZdyzkAwu+Ltb3+m
T2hL713R6zSVh8qNQQ9YBQeszdZVm+9xNRuLa3IRq14xHyc/1YXXaQ93Ab8sdmp2
3PScc0Pku9+v0mLpFqyeo2XNVP8bWH81ptCXWEtejyqkShl5MKUkgmbKPRaidF9B
9L0S4wAaWu90EM+XdfOFcwtrmhT3nVuOJr7hZAk3FSFuLt4/dP/PHAsEwAejGaS4
znovPRbfAWcFdCxk6FksDepjUk1vE/KMxNjj+T1Af3Vw0vsiAUl1Q5c6+jjg3ttf
nkfvymvUIIrEMUXVX3z08yG2MO+3ZFIwp0hG8KUY51xlTmljAkUQNGwJVmLhP/Re
8RN4FkPrIL1GkdiD3A9EIi7QSkQPH7Wjn+opHwRu8f0dmnfpf4cQNxr7Ch3NfnT+
S9/svXTTtwfOr1qEkqaOITxDqx4MJ1x2sKUbeCUZCIOoWsSd2xOGDiP0qleF9jkw
UR9qTQ0WPilwlDRjUZOVTldR5oZaFTIiNHC9E8Uk4YbmVsGxmBpnzkZF9HWElvTK
qtJrbTHIRj3/03NZ2FQoCi1eOHcrU0RJOq6ZzLwq+bey1TzNejhxk54rGJpiQm11
gAlVYvTggQX3Yr0Vsy5KYt88CcHqBRpHh4jZtaHeCZu3NWw3+1f+aHK/FGN4H1l5
+mdWcXHhsrT2YW5IwYRocGPtct8LaHLcqcqpaoBaVntDHD8yj4CN1EtIVfr7L2a+
TvEb3k30akv5qh4u4IrrXxoxY5sfhaskWb9Af4La/WhE6wggLYFvWeCwCpsMMm0P
u3HBCem8Ey/EhRNpEurRCtRAyXD48LLp/xEzTTw1qHVPkUS7NhS9zfnLcLEjOOMY
0xYoSOCwW3nOa31gk2MJ23ABNnBriS2QmyrJsAtbaJeYJ+J/5g2IP0A+T1rrMlo1
OlDMNDM3bxcQ5BHVkfHO19zEYYIfrJoGdnW+irMXHle7RKY6DZq8wukmaCVD7uLh
7g2xVBq911OIWrd2ME3u312Ba/VaNGoYWKnhqkKMVxNPvEFqDd9ukYCwt/oW0P+S
D3Y8df6+nG7DDi14ifLnRTWnODHiwiWRxcZPNmyoTi/AR/d+uGvHfalmru3GJSBR
1FcDUHlwhYgKX6jtmNhNRkgh0LCgCYQp4jsbHm2lVcBmW0TcHrL6h5D673gzSlHd
Rn0fbvyjfVpUuCytRrhgTq2RmyYf9nbeSvET0FwkkOICfVRgPh+xFPlDcrPcVCBM
eMzR2ntOBXeqf9SEKn/PN4yAXiBwShRx22NPN/c6ehC8Wft5cmIRnFGlk1ulYjfb
VrG9FH4NcwjJi1NQex4TVXR+a/XbTZeJ6UurAPSqFmBn7zs6LRiJLzjwNSF/hvKO
AG9sRoIQO+fqbHw9AdjXIp+O3JGoZRG4e58+5nneN8aSeJFXKciODt/vtNm8bbh7
obQfxQeQa5cMXUm9I68i/bWPdcZxd/pnjyulAfyDhkWtNcAZWXtxoWfRtKS2N7Nk
p88u7VLEbCZw/tYhW6Qr+g715pMTMtKiyq+gu47eJ7eETRFnmX5TAyo7OfgBJVEg
7zUINtKalA/Pa2Ki8DYUn+8kKE7Llsvd9dxEHWyMP8LI+1s6wustwdEj/2U3JEWS
LZMk3Ij2ORZV4AUZwYnLJgLnl02rtaWVpUx8PkCkf4Uo0iVSoW2OooA7NGCvQFoZ
CDuUtaT/JofVricHRC1i0aTZwAgkxIP86B56Lk2AwYd1LQTBtARuzuRXKwAG3EYp
EaJLARagnHAmbSRB6G7peei7mIgaHo5vHrqlizI7uAUWJlQtXrE7ItBtiWJTQXJ7
xnP792grZf/IbLZtqm/wa/BdUcXR3GXAME6Dn+E9QWyeMuWKy+t6xyfE0ISckfff
0xvya5+01Kjtse+Y6+6SZJDrDF/qNyGF17UdaUhTEJ4jRToN5hnW2tmk/SmAbssG
MEpYLIZBRlRoiTaFjC9pWqgWkOAbBgf7JOpXsWywoGMxQSehSumIyisKSHwlE54J
tg4t/JMytusQKVV6rtvSKmVMcNzaqUhOnVmdD3Y1uspZvMhIflViy3Xgt2QSCv74
8VWoQC0aY+OG7shV909sLJ556WMHRB8cwWtPOmFQRcEkZLy7tPCRu+yR7lfL0IMN
UNm4KVFjrdQ1NwyFM9Sd2L6IPQmOhBaL95oFITAd3TF26VOkKr0M2HIkDq2uLi7n
tz2LGHKHxTvp2Sr76zTHz0kc4r1EMNzmaQ8ZuedtzYTfXpp+h8qe/e0t6M/7GVnZ
vsVNmJQ9Y1fZkA01Tygzd7f1X6GXxDEfq1g/cfHnug2BabasaV9Fq+mRgsbnHEqw
A0RSlkQUl/MFKaUbmY9VpzjRX7CSpK+d48Xihnm/dWB5uekkZGy782NXP33WRUeF
QKTFMrLX7Xs5NcepfpZSbJZ0mDjSKa3HaUoFDaG4MUe+f1dmqa7pJakZAU2nNvcN
1g2UgOLd60py6ybC2AkzrC0+bmqWSpq+HbEocYf8lY+9zam2/hSZcPONzZdjRdOL
Ghqb59v486OqR0SFso3WDNtNCTfZtlop7KaEfdrGGVH2EWxCPLW08mbEMOdkiLCK
JMe6zi2lkNHAS1/eyDpXca5v3iHBmQpB527SdwfOk+JRpz9c6BxUqyH6TaNn05UB
QGb/6vektNS37ORBUvl3QjFeFspiRG68Q5v7JOe9UHBOjZ8eh7E+c55cVG3+qqtb
r81Ncq651Bn07iUCVblHe5V/zD6S5ryjQs0jU+WiMXqq4bIEzOcw2n5csGNnRM4P
4vxpcv0S75c4RBwOcgedo9ys2YefI4m/eJEewrFUTBSbeUF48XDN1n3CZm73t5Fw
oRKFxUxfMa+/asABFTAoeAAmeWfJxmZWaFchZpVRhiluYZ/KKvjcxByGN7esLrTf
C/gYRl3uzhgyxQegDJds2FlDDqEjg29Nl4gAx+L3HPj9T9l7kK1u5SbHeV2QHHFH
+jYaMTxGkzOKsA93FA2tuA2518oLTfoUa+9latthjSQBse/uyuJVOc1BH+F2UHLn
SmXoupJ6VRJElPqjgU1VBP2srpCoXApePYRUYFMb5/QgUTUJric0SkwM/eCcN07W
MU5L5tZwRpHUACBlukI9Qc6kHAe/rpye0XlE7NgmViTPVr0dmzvhWrAOBA/ycabM
rLFk0vNoAUmoKyAGIIniX/bMMXLfA3zmIc9viN103oL5UPac3Y+zmdbyCuHM2/Ls
5EIRWPlRvgW92PYYpdTeMgEm85wMSq2r4O6V99uZ4JyjgtQL94hmb2OMfdGv+YHw
O0GpTX+9RwAcJkg6bywWrtN9s4GgQJyo8Pw7BimWkQgZYitMMqsVymEnpD+BdrM8
EuBTa2uY6iZWrPrWVjjQT73wQaHRAFNmKsqO8zKTYFEjh61bX1KxMB+yhnZWZvQP
qy0ABWEb0wjoL+jSu8Gd9Qh3NGEatVrl5FMJfcCd8kzXv5sA8ofuC9Ag4x75/bqP
zXalbeVez6huMdlOVhBCwmU1eIZf8nccCFiSoFfRkGY4LYXCqUY2MhKsc01vNRWN
rNlrI4QzE8mDkTSwr7AzdYHQeJNe61I/w6JESu5soH8Sx1icet9fz97P3CDuLKZb
CfKdVLVj0GBo1H1yOB71RpIgCweFsmEnxQqfIhin3Fu0QHjCPu2OXSZEU4e2yUVD
+zaOAOPGA4DOn4g1OWBDCz6Rn/K7PgBXTn8IyPm/zaW/mYdLZIjijGTlP+y59+sh
qmxfGErtGD65/NsnVR3bnUJWcbdqm+i0+3rlHI9Um5IYeuGz6Os/s4cKYE8uIxCL
FS6EpcwCvSjMmlykyOv+PfO2GABL11V1QiV6x6xPRXjP1VqiQKnjVvWCbjE0YAkl
ViruY9/ztEd6ZnJF2JXuDda6KLnwV2bQVkXiISSIvapA4sE4U6x/feyuyMv9pXLV
Efo+d+XKGMuNfzU8/M2Luc2ZZTAVRvGMHvGreTRJFkuUfaAzJV6p0Iu++MOUISoX
tDO7TkDzk8aoN2WWJVfK8GWdE+tDB3T50q+0n+mGNwJ0w/OU3hZxub/J91OAwZ+g
YdX5B/HOJYreU5gNBskoC387JsZk1PjpM38B1WsR+68SgMW1G8fPzuDr6JOgw1Ov
1CzOMbymq/DSdog7+uvC3Oz2ze6/fu0HXsiH6rYXOFzQrqZm1lwbtTwMqQoGR6wE
KVhYTZaPnSwCBpKGgJ5myL/2Ypwh3EYJicPCFI1jx0viDDmdlfoRVu3hSi5KPc+m
M0WpxHDWBS8d0kXt/APZt8bePodk5h74+P4gEmdgxO6tv2J76+6dYEUFDd7gNAsO
RL70dRs1vgAN6xBgIEK3EQh2QpWzmUg4yIADzHApYE/U/u6FrCkpjp6ugxQMFcj2
W3nyh+f/RWIbfkz8DkrxQYpVB4eJDiy4ZcdO9VwfMV0dc3nThKFR0fpnKD4VJvXf
VDKnfoddHpwFZoTj1m7fNDbjpUtN+jFsfyeLkShGKMoeX7qi6i1mRX8EAXAva4Rj
/PGkCB1QjfYmxai6jPReSDbCUs9d5k+4ogOmMy4q3B3+gRrIQmpoABJTsSyloIha
n6h8EfSfolEVbYNU6JxbiIs2qDSronBw8OkFdiSb9OuZeEPKZQtXP5IkgeVsdelm
jSUTiro9Ph6p4jK9zmKeVyLQt/i0ybNWiK2Eoun0zOkG8KD3J+iObSWRCkcieqOJ
C/WZ8Ce/rSKSjqJZVXIGCLme8u1D6H3m0XE8C09XJ20BWLKPoopxbKZ7TeKGfRQF
+xyJzpaMrJe+WmhOhE5Kxl3bwrujlyWg2Vmx2Yueh9127a+WX6FGxQir/1k/K4dw
zj4lReDNN2f3dfurE/elxKaq+l+OJ6HEIsnSDkZXPqRM0Ui3AlI0Se+ju+X0vpHF
U1/FW4kBUr7xaoWOgIigexAbIesFbgnl8EV6N6ksIRmBLKerT4UJm1gSt33LMgZv
P9bHS1YTp+0q6V02ew1Ke1WzP1iR72v3D2pw9LeOYDHLho3blWL6oty8fkG0Bb88
MMdsSJDw5k7WFBGKOyKaMdvcWubgMRt/YjCXihNryVUJZGBFqlGj8Su/mCprf+FF
iaw4+cPdlzZAfBtN8FpuqlskYIO1APYuann7ksn/uQ6AwkXGcurdG4XwJcg0Ix/i
8qVVhPxaiRFZFP6tic7hqT4pQ7IGRNApxlKYS2uZ0hFm4s+zjDR0MCIaHe3iQ+ip
cq+LCBdsgILIZeNGDa5q0hYLyspKp8X1DLfxoqOUgiBELGj/q/CfMeoY3WDGFauZ
oMV59iGmbPzrHN1VbtlrhuPAHW09/YvxOw33ia+fQNLoF7LhYDEvaLxbCq1xuUiY
vqIQyWUJhtO80tSgrFL2nJKeT5CqUZZNJC/Es+4LTbXRoptSTHBZfGZ7746CYAKF
ttayXM0HTGB/DKVzch+dWBN2FE5hsOE0Esph8TAgB1GEzOoFNrPo15l9zqw0vHxa
EtFAu1fuvv3K/J1jAjkj6pAQdIAlQxes23Bc40cdHM7cMlNCkfpqB0yA0sD7gIr1
CDHc8oYeXkiPfuPwC+dEGXCv3VK2kvcuu3TXGoR6g96pIzskfV8wD3bOh9VU2tes
ojIIpJuC6dJ1dZ/9A+Xsmab2/YHzFbCiX+SQKWj+Tn9w6WOhtQPKTE8GLt5p23eb
p59/IReMjgPQWRPVCRxBE0lPDZ+x49LIyYa5lsZZDo1DKgoZdPlkGEGc6ivBCMBF
1rxOO3bN/GE9CcKiPXqvBrg0qwdTlKW01wRmk8cODxVG9Snf9re8pphlx3eCTfKI
xxDiBvneeLf0XzSNobzzjqGviCj73GJFFpQT17R2DiMAbi+TWNCjaPtJuUkdHB1d
d1htjbm9urNNRrx6ZQRICrtnJNPml0hAvVg4zcpe0II26e98msmPwptpp4KPi0Wr
Uoqal0nYssAjOX2sw26vtD692mqDIBtlijpqywyMEX/z54iKq3oqyHbWQ1LI0tDa
OJ8sIS/E0yFVeJc5L/eVZcE1cSoHn5faA5fj6x37pVJw6M/j3I5/ICBPc29l5RoA
oOXf107zRNv/RopE+sLkMzzoEhwDno6pB3tfWKHQRc8SzXpR+7RDGPpvpotIrzXp
P0d8vz6qBnZF0WN7PluerrDcvAAVx19QQg5NAs9c92WYbxI/X1VFrWlVLAjPifYj
fhlxRKOibD8R9VQWsa39oWV/YfvMK9kbTsOiFDw0OlBqx6CDP9yC4x6xpq3NG0dU
QQ+3YCBR4IjAWso5PLOx+QzK54f5iG058+8xaYalg5bgmn9bUtHeJjwxL4aPeeZR
oh27F+6ER4gGWQxti9AgC+dGbQQa2G/MbVM/ATClSG452bnOeBOCElsWGa5S+5Mr
meOCbMpByKsuk2UUu85T0M2lXjqXHQaSVoonvEslOUy9f/DoQZlYNm2JQUhTkI9M
PMXlcI4E8KJJQ/Np3BN2MvaXxDNPckC76gH++fIXgTvzsJMLGUtnD57jTPnNtgSH
5BRhNAWw0hWGkHIixgD7BZP/ONgXfxZqXfn5SDehcRjimHpJ/2wn98jBwq0ZpFxt
sXOajBM3XLeaxL0nQsuvSxwiVuy9fpc4OAB7HWQPvRZXeGb+3SZkh3yCGyEyg8t8
U9LADRF1bfpKPp5LuUG3ZIf20BHM071k0CZBBBzCC3Eedy/cOGQeYzyKeZwCskUd
Slvx8u1dhCGeLAsni10Tuw0RkOtQAPOP/RDLm0nBE03DDtDdMPfkMoy23sIf/Dxh
zJdSWJ6IVKpqeEYs1olhNbXskKVs1kQVebLvO63eSVqhOePlpLx79cmbmFNysqRr
M5s2Pk2V+ycy5JrZV/7VqcFX9OgwZK6xwEDI3XkESEIiyheLNc5gg2pks8NmNUjW
HxRJ7pZDYNrmRRLGfP2qlvfYMU+kIOfu4RPTYWj7enX3JzxVYEfogvqixwBYxo4X
3fQsNGWM3LuEGAxameKl2IqfX6MC0z5urAq5RhLHz8gC4B3aZae3H1koCz20oJDV
XhWwW7+YIIrOGZeodmeM4jIpkJsq17bohFpNnnoixTAhFLxp/hNF6l1sgdHtT/zk
k8s2aSQ5voujXP5EWzx7ewdYMXJdQ7BGAHhUbiCIUsvwjHysl1YczJrajx7F2rbU
Ep5UvtPdEBVMS1giXsN4TxRSNVv3rgdgy99/CxhSPC3Hw8FeZ72l+mYAUrtAEX2K
UFVtSnsQ6SXcsHhVtiiXY+csF3OKAakqX15iDAEMsTEfYoCEhQ9hU6dNV3x5vfG6
+PcE82YoiUaZrhiI7AHenXJknRRgncOnhjKolZL9heT0anBo5w+wVrKIxcuzYeFh
t6R9NbaHh0sC/eetqTN2m/dQh2jKvjoS1xWy7r2cD7G2pBg0i0YCmbR2vx1C5cB7
4dv9iNWc93DNDTHlBWwkzj/0qwWc1ZbMnNML8mfqSOBDDewWSQDhF2j/ydJWn0TA
6BkSJYabEFafUQgQQQ/OccohsWhZrhgtbUBHhKnLc0/mew5cvtyNGl7mLcRhVr5b
14L3sRWIVpXeq2r7y4GUgij+kGpLFnuOThLfqq8gMDfWEiL4DNsoBHWHW59yncqp
qemN7iFJ9yP7wUtN2CdO4bTG2TVkr42YGvCwngN9feKob4z377CRst0loYMtHL3u
IhJfv+DFtzXGf+hpHDLEdRdEKunCOnNmiGHyMXyAXAgYXAG/Pz7xnETGl4QIeILa
7I2ArZz36EGZh6ssnhmIIcXGaOOlrqdGpKiZka/SVr7oWhVBOBSdbXdLU4LnUtkF
csgvyfLQByeuruqojhjUJJ1zarc3yuf9O07VRU6P78v786ITVTIRD//BxJm29AM4
GF9Xz+XTEH4DZEHJNL8JN2WmbYqXaoRCY6XKBQ2eMo1qsclo+A4cotfEYjMfM/xw
zOeUGSgOiYo0U+sZpSOgISJHWFKInq9ekjZ3fbJQIxqDxdri/IbNWT2itiwORNOh
isxAlnSHPYwRgR+SHdtkGANBtSx9/+gmFgVuwP7b6ryGFlDTo4Lpr4AHZBal9lQb
eyATAwHdQb3e4ZyLCL/mlGkgGLUo2poLhafQSaA6Z+XJF0PfDfza1VJpvPlU80LU
rCx656rH9+ZNJI4TWcZXQ0bJjd7GMBW8QdQX91AD+/hlWwzW0IfDuKAbbzSRMZt5
D7WavXNNNUxpHwPGDF+iIbZEFvuU57wFZuu3HmkibHUDbdf1P0MgzRMDMUsU6SrS
xTnfFJjyL/M1xmCiIajgttoc8OVDLbDgsgQDEsnODxe5kZkCu1diLhIuv/M09vx4
F15kdXG2g87MYToHYcCdZqEAvO1ZrWv3/thcjzR8vecWli27pkh7cEZUAP2uzhgk
MhaXee2LMuV2VC9ZmoFMkPLUjxD1jHWyHEtniUTTE0zoJ8+JIWV+oCCG8dBOuWBF
CS8AdcsmmM2wGgMUQNOSm/jigvzdjuFFJw8fXP4vsuVfJPfB21h0E2+Cl+lA+kEg
mKZ8TOjGH2yXaDJmRn4eV6Q4CstUM/tgUcfz0UGDkkIblSQXBszLvNJK6SLXC1Ip
wX8YVs2p9vE0Wkcrjj3TiM3aymLg6Vpg09Hnw9ciCXsZVQ3QugLBoH3YU17f9MVv
W6rvkMtSzd5DYX9rouTsFhGP5ZdUKbfApfdwXdfRa1/WClYb9L4BKq4SzHmd57Iw
9Jaj2drHo7/HFAK/6DiqkLZjfOMAURTiejAU9t74sWSctUo3BdYgVVZRpi/JsSNN
VzainGdFfyLI6URxX4dILV5rlnsDYfFNbbTQD0raOtwYWdxIYmtWd3+XbxrKuvaw
xEuaGRagi9/7f5whpPqqCZrwSSgVhPwrNJi+HiRMOYeEnp6kMxDS+fExTXtM/Orn
OgnCgegxk7/aaH/tTkHTb7MM5KYuD7KxoAw7YzJBdVvhEbIZS9oLynsSkA+83OhQ
1+hTOsF7Yiyd+jdH2OzKf4d4SExwqs2HYPcgtCNBlPNmMtzCVIq8w3JdbD4sRyk+
djAkBryn4XNi3f8DUCUISIkk2tUgkerGDJcyFabAOYJH+5550j18JuNNtAMfaBk7
XqFEGcQ1gv0g141tvLp37XsaE2d+3fgeejPdZZb1ocP7UKx6j+cJjzi2yAxcYPEj
UIXkC6n+IvlFHzw902wf5iew8FM9oWGGCE9e87f59adLO3NbFEnk45sSII33HkLD
IVfYTU5P79lXJv1duAfL0xB7+FONGkIR522Ym9gizgx8P13YZBE3AUjLaZRv5C8F
iFzTH56gBAS+4mM2kZa8T9y278jdnWiXGfmNzRtdOfbjwBHA5cx4z/u1pW/Uxssf
xU/eJ7AbEbQV2XUuD0kFAcv39KUXy1l867MR4rciVIqhS0cHYfkCOU362jG3cQPT
V5Wzh0/ODVuc2LDlE3BAcTnzkwTM5v6AsPlIOCpwbQ1zKtjSLWKUXxIE0wFqwbpw
JR9gqw9/BSSt2+S/pTLQ1CFe3N+bhZpt6nBuDCpeTLB4RuEs9UuyenqeI9Idcwc8
nvEay9ycda01/GmxcB7Ahrj3C30AV+bHaI+9qXw9lQS1W5gb1wT2KwqUFgiyMwfk
7JpKERgdjxs2Mjil9T2fv59cWwGN5/OP7tbR6MHRTZxO//reJD9th/gunMw7y8IP
xCqdFPY2SvmeXR5yaNb2DOtrbGEGL75D1GPQ5vHAqFkcaV2nLAY1aNOHC3tHynAb
W3RIaOWxZfCfZKPdXqBZ/Y8VypNRV/ApS/rf5ZRNZ3wHkV/9rc8abE6eHT3ohiAj
KbKaYvlroYmXEdrgTXw9DfrXnrQcD0JS2TEIRdgUhSu4Pdp4JuzW8gXsRV4MhE0n
5GJtTMIRPGDhqtmFWqX7rL2vFaqMZLlXDEGUyVS3N/5fZnvFjT7P+py6OaBz9VTq
y1JxZwgjFdYp8aW9jBQrNn/G/7xX8wecfowY89fNUnqbFpJurn096K9fu1rYCX4O
XWZ4708I/fQHL9C7iLR958lQ820ZRMbDaaYpACc6iihJwSIFMrW/E9tC/t27FWIU
Y73N14E1KoXgHft+CeS7fuZnFAfehJOEAHP2N420A7fqEd5yi78Iuw+6i+lhsKB2
YWnlq4xw91Y7yGMWFwJFM3glUaSNj68VYfDFFzKDjzU8NyzJiN1wfRLNSO837Tw+
sIspuVSMAmNGbmYJVvfbOmoq9z80y6bcumkLGyfPCXnE3vhlLnMlLTD2OiJitI0+
RBetVE2ypdusvY+rXC1lGkxACy9trgWLfSRezUyDQDlHx/ZmOJS2mrHTD1PqAmhb
tYkqunr8jtnBHrwBzr3APWFPvaLwG/AE430rDgFgXrp6UDqga63JxkXV3rdtO1qr
Vj0CivT7T8UsUJIwTT28dAffzNptMe2naMLuqaaXpbhw6yKBKUATFvbaKmfaxwkK
cJCLUWWd54/evXizsOtUiMxquVcHdPUoL46BncF0+2anf7WzQY1oSCoe1363wK9A
t8HGpHRXAE3yCuxaSryX1PiWMcfNchIxVNrwf/TabF7izWBqzuSyROGh1vcdk1LA
EigIhjq6Ch3bWql72Ift4MX3rZj5PZV3x7lKq6wWhYmoFLUb0dhHj9OK8RhwhfR7
NzihFplzVRDAOW3gnWrMFs5lt7TYDA4exbiqkpbbp028Ia2o5TRve3UuVVC1DkTs
PcwWynA3/yzZpTdb5Rg276kmO3tCxqtTN9/isIJfWtg3oPvAnMbYpKytokv6bJpp
Q34gKly4WC2cc9Ts7qX+d3ykRfv63rBRHNn3nxD9L7YsFffQ3LKAPuIc9RWBG9IY
v1cYWQYT6k5xag33M5Tzn5y6DHv10nNHdERVyVIwsijfJRZFT6yL0ISWAz8npb+G
6Hd67huGTn1MoA7++/wdPq2UG1Qx7UKK4uFdjR4P1qL1SSV2gIZoP27bfWMBkOj1
a4qJ3sLhyYLSLN6ks/+JcW6uwFfmn0/Ov/FAsAvjMZ5NX0LhBjvErF54a5s0dwjs
TxVXTLIV7xhxpzvUxL9ZxyBiO+61L1yhI8t94wNuJCufscpp2x8SGDBysozRHQL+
N0+glwrJJ7Xcio7fFHoqMWYSBWu9iBZwxSRw36nEkvPMlhc+kdf6ITxfZy8VDeoI
SX/ElRFZ1UEWQo1nfSbmAh7odCAds/e4O3FyV6sj5vrMBELMty2rCciED7NDE6em
ApbIPutXnaJSDapElwM8qF1ZjfyW1Atdbg4jGc7Do5a/kR/CF2IyfGpNP92l1LNa
1UyJ3PKKlFImnFLiTQf9Q8u1X5fPCAULkIVPZ6Q1rHe340VL7zrR9USIXs450WOk
ZqtP+oaQSsjOLuIhY3kqW+9gkliqty0uaSHBo25J6Z084Pigb0RRVNaWJ0xtnvaw
rrczPJnY+9KVTp1th5NiEuQx4DN8VhK+3mRGGSw8zUu00bseCRDiBwHMEVRIhydF
K9CtrqzxtHd7LSktFGprtXab7xtFilDy2aP1ljYWuVI5l3EDNe9hJzpeMJZHdjPJ
m5cNVrrkkLQL3jesKY+/JxdiQLB68idUzdPPjuM4qmWhCqsVztmF8+mhB+ImfrOe
HQAU69vkGv6Q8cdA7PQwO4b6FxaTXZm26tk+IxlbvXnsEHz7Atf2n8y7krlNO/8Q
iwSO0jtCtMxMCqjZHNkarKxngcdn/5wtq3PySfiKxpgiBS1k6IpqpAX08gANeV6s
QQD7eNp8WUYvw9a1e/FiN2ZDFlVlkoc9QetPq/PcP/K3WRqWzsU5J0AIwJuaM/OB
oqR6MRcgvXZizTjP4k94qiysmOeG24Rq8H03hBv4b2XTrWhrZDTfXniv1EXGXx9Y
C683HBAYFDDEZg9/OiAErr+gFlBO26hBc9A3LFJlaHuPF9PKy4VotQwsuAJmfiKE
+7Gz0t/xT/mY/xGeIVO6CgSQGKtK8NJAAwrH3CxeQe1kMCIkeCJ9csberftdD79/
OsPygsSESiAP03fswuQJA4nqZm2IwheTI5Im68Pk2o8281jdMl3T++J1895qKMbV
1PxCVs6vYmrAE5ZY4qt+Bq84VDxh8Q1bgvstSd68EyEORe63sAfOhDhWu3WusucR
L3uCU64umAZtocsUyk1k5oTpGoguyqEKF2IhtrnkjBikTWj3Xvp8eRFaqm+Uo7Zx
gzBHaCVRa4/d2hlqXt/zCByUJK6j/1y7K5NKfIr09KYqTjUhy9weN02n1XZqMCQw
a63tMuPXPXRI5Oqw7+psagGGQEegg2XloxR30cir7MieqvQnZzETsrd78rb1A9g2
mQapFvozgSukWPqm9Qx7y2Em57KU9onJVb//UyBR/bgGBSKToN3JRhBfORZrq/Ec
jBg/tyBddvWk12PVnPFJ7bDTmMSXDPQKQ7CtVGlW6kk9nv8p33H75lvJEovtMudQ
1/SIc6tuibFRRecd3+oydBQFHdSkBKv2uwdjiBJVR31p55w0vh/py2hw0z8P0xcI
c51TLKxQNtkrNQtcFpiJF9GwV50uZpSt3P/XuHPgWdLCd7JLlDAs/MXM/zKGSORb
nj7UcwUgHFK7EET9k6KewuBIqJRs6RIRM2rNiA4btxcN6lyrUdfFfMD4hDYfX6kr
rApbZMCBnIDzQuT+nttK6A6JjiRbzcL9945cbte11xCsnWEomVkuJuL4xYme7Oac
icieXJkvtRzZuzxw1hSqumhqwQ8lm3m1EjnbkCSqUHhvmrSbQd2A3G+DOCSJRb71
1X9danPbnhBWuGEoKWRjHvGj9kB/XE9OEVLJuV5Jsww8Px62cCsiRJV/443+fuIS
2XCoABeOZ35YnO7QxkH+wJ92P/WCz1D2AVJLQCosxNGWdz9kM59pKX9Z0BOzsJxI
ImrCZiO+i0CSGejWK+SMlqxyK1MrZZ+3J8ihdDaRt/VxNP3uVE50KSI45jacxHSO
E6j6S/NKSacUx8raabU37H6iIgEOLGOUTCciwXsIY9Nt6SXZAo0lU5yX/ZgFRPYt
7bK9bUr6odHiinuBrC+JCQQd7mC4FrOs4csJf6GZKm6PZ5z59kp//0/hFGxYArBT
3a2KKruDUMfAM+T0saqPbDk9PyfZswh+GqhpcA03YpwuxVQ1Rnm/PBIsAWejm9ss
xXLu40teIy2DGryW1+bps6LyztftjmIWm51u/zwOhyBuZN79KTl/Fqbz2jxZD3EC
v1bsu5PSfDL1PICP00zKcwQxMzs662J+eutfgWMJQS3UbM+oXvmAZW8DlV8qKoQC
l80EYWpMwBgVUl5lp8ocdjCVAURgv+3hlog7PsnY9E/niQnEy76YeELNDkN/McKd
NMHV6RAMYcfZShD2dOmDaUVzcy8Jmwa0fDihI8sBA3V3cJW2nJM9QIZU92xEwuUg
APGknmVaagAKCs1+QPH+XTx/kTRNVFTc8VeN5sZ38Y8/0n0v0lGlEACTX90m9WS/
uA/4QwlMjXyw4ddxGbxBH/Lppvri6Q7STZ2kxnBxrEZkZnuafi4ycxf9OmQhpJI+
I1cjANQn4iFPl4W99UZ+krFW8FnX/+w7DzYm5Uzb0/EkcQF9dAMWmfl2YfcswIIh
GXxMc+98tDa45xQXu9lQg7vTWn/NRrDoFi5DIHA2+gBEQLCtpCemys0bdAvr5mtD
+Yxt0NWwHticp2hZs4dA/ehVFM4ky++w8okv9Nhr5mVqaidPcLv3tPszsuYWIg/z
8v7ziJ/dFYVIA8KAi+cgMpWGdmfxKHA8ULMMhCCsPDICOLK5ZW1cVDSIrpL9tGoq
X9XWQ5x/Htsc/drX23rXXioEc2x9GMwWJ6xIcIKX1JSN5I/CIuOwclDJAmZF3DLE
eFDfDPmJnarl0je4DD8UIM0TC72IWVe0JWIdBLtYv8vAkOHJabtLmk8tPBA4TeMx
7ZWxbiGmf3F31ox2cAGWlTjZ375X9y+ySjvWKGx/hPPHQJpNxcBkfBZuURoM+eB8
xGHHHoFH50+POOcjAAYezQNiC/6qSJTakc+NfrMt6CwfcX1BPsSZw/+oixyTFDHO
a9YFxKid6/yWRRrNnD/SEA7DLkejDNQYy8zzOEqipZCEx8VRF4dAnKrE6kpK8SLS
Glq6gTFVxMC5p1T7XO7XY6atXhBLxsRdWHy4wkazxLNoJyEaTBXi3gHuwzfI46xX
UW5k8svdqzKXu5CoMu7NyPAza8PcSqfv5D9onXKexcyYq6IMAju6iV2xeObRCBfg
0ae4VorLcxNkd/m3Kzedmspc+Huuupi7Yj2/257t4Etnq7UnyJY9XtD9VmkpCv5r
0aoH2giZzmLTHVGk55aOEp+TdBQe3qmdd2aeJhQ642PhmE+WX3iehrS2sJ8iV2lm
W6vwyw5fImKaZrh/RtcB7MsOjNAfVU4pgxa45NvlsPboJiBSjJayGmKb8qnDZpaP
MdiOzYV+VU6+wP+rXGYKnYe5jvYrcmsIqWjoz8QBED8aUdRhfit1eKU3vnNuvcbQ
SA0Ny90hT1Jf2QytmqbetRDG3L13CvAO6oBBALeVy0lAPdjJRkVPjxdV1I/f4Eht
GmhGZOYWYX6AtH7jviAlxMuSGkgrgKBdvIZnIlZBlZKeZRgVMX+hiUANk/tSYEGr
qPIVp7Li8KwPDQHUQNcGFvKlMMApnYfU9tNLYyr3LmGzP1ONO7QmeCf2xVSkrk8O
KraP+TWtPf1FRLPOXRp9ordkj3Lr9gMhD4njJFz8w5QTBD1cra5GVMf7FFC7Scf1
ZUvypmDaw8x5+LMqnm10cRkiYLDXBWnE+96wRgmUe2npiot219JU/63zFGl1ABfH
ByTb+gGIvwPZ/DemONSFeuzGgmLhrocvIcRev0DnioBxmTS+YFjYPg/pAt93YaRd
wPB7pnCOavIPOUGBx/SH/HTWI9bes09Jxx8oEOh4wEYT1JzXTgARFQXNa1lhdmjk
WZla5PMRLf/EXgPIWgaxVNLcErfo4EmYfNtXi1xmd8ZT8ZhoLJ9csRisQ0QwFY1E
njMO+bXVrcst+E+dkFHeAgjdSXWO9vN8tqzkuBooIVdP+TatVRC0un1uD4ZasPE7
mphYdeOVzMNllZS/Lrs+Rd0lKv2BEOOVnIeyAc/z+Rf2GKNrbRk3UagO0+JubnzN
O2wFrxqU+ivHyloipOShP4zSj0GXlOEgl7nNzFaR1Zz56YxZ4Lqqy5bQwpfWzYne
pD21eSYxig5Mo5Jz7rBdYR7Qc7cCQTYT6v7HFlbi00wek9p8Mfy6t9OxNVMd6wPR
pgMTMPDbCLLv4vdq5tXmYY4feNtXmehIEICF1f1FNNvTJzf9f2XeXruUeeTGCRuw
id1CNZhThUHf/hxoiJIUKddpux+5wpMokfkj9gA/XotyAySAYUUloin9nKH4ncMF
Ja+wT5nN1t6rxQdcbFOQ2pq+c0lgQ4aCEJMRVgdMmGGLevZmmN+V3yH5TEeZYjDT
+6k03TLoB484ur09sxbLCccVVq/L1nf8A1Cku8QuHcIVG8qkOdnNmLPagMZ/SHSC
mOUdv4mUGoyqzTcGePmBC7UCtdpdVOA2exICi4vhSDDzMGDwznMqwWNDh8pSX770
TUmiN21uVlF09G1lipCgF/hcbneczuaxNQ7nxOSvG62WcUw9ACuIvWomZyXr3O8z
tg8eGZK9E9+S2zYpXYx2xNFby+Funh4ExhX+6xgDUf7v1XAd4Z2EfAslC3f0yBAn
JGQprDh6a1ehP9jjhPPo5r/Hhpw+mhFYMDV+jtUUFNkrR7kR29fmVv1EARAPyu5/
wuFpZPhnbTzx86PD8UZUeNYwdiUcK1jLx8wgKfBfrUaHIPb/1+VLe0ZtPoCyUq6K
ksmqx/DyhibNIdOB5dPinb+ZkFEemuIJTyyacH67Itjt/qgQffDwrfYjB/5ULxxG
zJ6Xa/AafV53OSLU27udu4tSqXpL6ZHwKs55xpyqQAvQcwL36W93hS0ODXTSs3A4
LaCpv8yP+7ATnxVuqPYY4Y0arGqLHItY0yNvSZ33byzfelbKu1kj+RmNGX3bIrWm
deX8Z3TYgMwp2yuxGne3npwSFr9VcsIRPb84G5T2ySCP8slyYBvLBNNP/9iH6x6M
lfcgjmO0y/nQxC1q1Ia4WsObdOICPFeOovrP/vhIprQQa31/gTZTFX1Vh9xhWfou
LfxD1lkzp6iZ4q2VwPcDI43OdtGaVQMmj+qGbqX5FQz74CBa1S4KmOj48N2m+7t8
PNXGy5m2k+0JVx9g0ayX8DMjq+n3fdYjgap/BfeKtpZXEDhlIj68nzFHOTk3RTSP
R4bKUfAyCtCRDUSMExf4y+NuUrxyfB10ETjpeVWbtm2pFNMVZQEDsVePjXPC8tn8
oXY48OqHjlqWZgagY+Qls5UDjFsamZ4x6LersfoAfQaDk+0iCp2vpzok6rTxSP0Q
Qoj+kWoSwdMk59BM/SgzFacdQPfC4KfAWs79Y1mrejKDgWuaLthRsczxRzNlrEJB
fnk1KmERFB9X8jqFgEZovkuOfXE6z0GrwNueQhP79DwM2mwAK99I/x5CN1Gv/9UN
5aSj39zf4pjlWTtkZxpIq0G+Cxvxy6hk/9TNWnNaOzh+sg5hZKEDKEckp7e5r3gH
nS80K8h6fbTGxEABbsB262HDFu/HzBKUiSYFIgKBq60SGbF8hWU6xkwM5fXEFqdh
6YcBK7Q+2RTHylOs5cacn1nu4EDdAR7VCnK3OlQOdRHsrPT69/7jFqsgHj6s16iU
qAcjkNal55ocQClI5flX2CTc6oKnAWWGl61/9VILsFtQYrsE5mn2bMoBy8tCA9rK
v/Idn1zperHJ12LdXYVbVwtkR+bfl8PnBMxODMBCgBCWhmm6GcZE8kGZu/aLINCs
e2+g/hoyJlotwKsZIHDBvPbTQIG+aVi+3R35VoUHWzgKltM7zImW0uRC/FOJnNwf
Op3Z8QM8Uhi7+uvyyTF1T5u37Fk65f3ZMkKQQuad4XfkQRLkiLDDBdTC9uZAtoJd
T2P6hM0MlA4FebsPKz+7V72NtuF3WYSbqDEfw0hWECFPiIbgxEuiig7umOsBbt6H
mQq9n6UoP3VrZQj+umqNd6kjw9kdriySph9s8FQurf627QgTjUtHeVoBXg+MFB3E
Fsup3VXCf6FXsGucR44NsUU3XmzSC6WEtFm4wbu2z1JQOkT3yOMZ2XuDVr7RSIAP
TCc/7OiMvlL0ck4LgoHY3fuLS0KcreJJrS6HQFPvLbcDkX1XkTWVn61vEUuWkuul
YO87cP6ecymcuBgs0AIpH1VnfnyzZHADjg7DiDHYStgna67HbMiDw8OihlVzZgQN
IT2l3G0sT/UUgcBU9dOHNDCcsEL7TNDjCMzHfelNt37LVSAHwPsaXIC6pFnbwyh0
QZ0Afl5kdhLUDYvw3YMdyO1c4DRIIJoPKLMvpOaTyKxqeeI3bjl70LAwlbZpBjp9
YKoBGqodDH/htWjaRem6TSc5ux0U2uSP6TEC6Vsdm84T8RWztDbzUSRodRjZWReO
TkdvUGNE+2hmvbQSkiy2kXtLc8Dwg+/TSLrrob35zuzlvA+uMgapWCXsg3TZEil5
SaaAjvcw6wGsah+pckuSsNKqGVaZjbKw9xW63+2b6n5W5yzfBsp0mRkOgmbg28Ci
kAFVvguB/AzXvGGcbyApszptr9WEj/maEWFYfXef15SfhHUk4KK0K7q5/y0X+K7d
L8jKt+CjoHIUhcah4OnSclZpMcimbqxfgzsrngdUzYyOZuHcBePue1Vq27+Vu5j0
PikAew4+p37T9nU/y3BI7lZ0SMAoZGw7jL3puBaMVdq4sGApxYYAcZkJSuyOyabf
VRVkzBSp+3zArOvmZ7Ldnwi0gVxI2jSfmnkDwmwzki/htekfVvayeHWvZo74gcnf
oPB5VSCpQua4/StfxukJKW6epTM562CcN+EyaFXjBHOecIi/S0ld1AclZ61/wZJj
6hW27z/uE8/GXsE7YxZIE2eo7474gBmToLZpDWwmJV4As76gJVD2f2S5Z87VMnfa
etv0hYvrjo3Hyji1S+M2DpcYUd3C7iZGKavjiJktMcr/ZSmerE7f8mJ8Ye20uGrM
VQJ2U9L1myeaI6QpIUusax/weNpjwuJ62BZPwHfCof5tNtfAqdOKzZBuYku6z7Dh
CYIOcMHN5pX76nwetK4XhB+xtmYmjSvo8a9x1SxcD+BJ/W8zhGqdDGlptS/HTcOl
VNMZmdl6ku97rFdrpYrlOq+2nf953S2QNxF097gPiolnkGkkKHFNStfI29ESgwBW
mBnXytv8xG5UhuepuzrIAxv3odoXxgiYlaHzqaY+biLq2NprYVtRtx53m2plUB7x
lGuarIj9hOC1zB4HdPoLkKM/ymfV80ALiVXSBQ2WvjNXFom/f0msxtcfpBMdVdmj
VQLHZisxWmOS4QKhhe4ihzc8PDR25sNcGuDm/EjsF1h+iXkHQiItreMS2Ld70tDY
wcEJuy1LqQczRI/exWviHEf9gtzlLJ5llSyN16mqF+R/wtnDTpq90SLUvAsGf2kq
Kqq4TDauvFbI3us37uk7KEVL5LBEsUSHSgTWyoYnjCiiFybwoONz444z6Alm9u7y
FUia0JCj1oNNLZdfsxBwgjql5q9mhw/EMgrG6VXovdQjNeO9ZW9lrdIP4Ph++ZeZ
Nxw5mem6kGrwGgxOw3f5ERdH5QYBfOFoJ07Yq5ecVgiqX8GetXRvS2fOjPVzaHS6
yzgEBxX7vpbtUXvGh1ycPpOEfjlcsskWY+cQgNgVSRx++JddqqNEHQL2hlNh5qMf
zeW8R666b0JdkF98erAgH1AXThiezN8c79XW8ZUs5h+8LCEC9CARHv7akoF0McdF
7NnR8ZGUcZGqsC/2nnEmdSm7HlOs//V0wdWjvbeLycmUOnvUoOd+PedmfJhQ8l4s
Fo/Ma4ekEQ5abkWQtwmvfv71nplM8YqEIKNHisHB041lrfRjhd4gqJPqXJS2T6Tm
lPZO+uWZ3n6dFBHDlooE/wGZsu4OpjXUK844PnTnZJjBxSv1YLLIWuOBzSwJKJGs
p/079x1h3izSDpDHTkqdJ8MWoON8Sl6Ejuwqu42pujPqrn5QvxNlOIEve4vBN94F
DPEMqbn+BLUHAjtKr7Xc/M0+xa6/vNMicBKohIlf1glLD2X8d2BNvv8uKXp1UR76
69iOAPPIrfTMKCQyjhBKIVeRTGiqlTC098gkkZ9A3YHUu7bVYn9v6Uf34CRX38UE
iYuZnK3A6nWuSLjpKjkgIfFj3XmrqX3+52zYtAbhVVfJXKF+9U9+dc5CbNx+FJ6l
K+Bv3zdlmGUlaMPToZFx/HAx6bsNvRJxrS5NEWM7DWZy52NGS3yDPwFFOKoJgOpa
J1xi7siwuVVnKZlkqs5+vaq+oTxqy8HuSvye+cSCjB54bLrA653p9jzRPU03rGlK
DtNkOg10k7j17P1ygZfFpoYR7Pehs2tsey9WBX9+CkR+nXcI90tdjf7MGTSYfgaY
xsoffWbqIxN8ZY64ksAo5euIpjO4Rb9ZGYWKHhG6IShUXntnavp3FqfAxlJ1imBR
vIIPgoK4vb4zvb+5lJKTvNqP9FwvjqY/3SRdwZ1THSJTT0CunGc+EPRdZTAp10Nu
tdmUFGZUhkX3U6HRFMQJplxoUSjtGXpFlkFYcZ+JnzhOcFvjppyp7KNYz9bm6go7
gSH3De7VMY5ZJ9h2pbPE8KsYd7n1ZP/7KhxIMJEdJO/d1vnkoxEw6UQtN/4qV9Ek
2AcNZU5ieqhZkqVLN+pB3sdycUaChAKLIjRyAEeGOsMW6dSQuzOrWVHpnzORKTJd
6pTXe6enz5VGjwOm8uph8EX+jfCwZhbSK5vV2MNVIDkIwnUw7b5Jm0syaO7JK0ty
vXuUo+rJ+gXt0158gF5HU4cnry9NdJt4yHgbPjsZY4WtMD58I+i3nwfYORyxK+gH
fnc/bHRM4IxZcaSRs8eYDVLoktGTkoJSy19wNjQhO0+p6EtY6H2AjMU8muuRcmHJ
yWe6UZH6JPMb+4TVCM1Pwhuej2utTxQa8zy6ds2+kdblVKOn2Zr7902KmIdjCmqi
UnkePSZxFcQCCmvrHy28U1i3BLK2inCIdu6ZaQdhjOdb1auOyQO/ubuVD+8pFNyU
++qTO9mZwSNd4Q6U0VgSvTgkssu6yI6M55ho35ROmNZInsWoTupr4Ryb/Tyc0xiA
jJUVTZ8ss9caFnnZqfMv/AWQHia1YQBD5ldkdeARwuZucnUMOlmwN4TNrCtnovGG
PYb75HqI+plWULpkt2m9DY+u8BL1WLy8O2dyIj6jknq9jB0VKLglnta/8VeyyFIr
wG20Kw3svW8uUmP4Rq95RT8vMGK48dVouuYqVSZEsJuNw23NZU0WdJzirgisqay5
oEWlkD0bfK6k7h2kefwx+YFpBhY/iW9Q94g+00ZRFax3cCMHfwKm0ITbIcZsfDNh
6WSuSIgNzxsejN2o9nY4oS0YddL8tfEGEHoDRCRATc+LE5MLc0I10kx8AN1jzp5K
Udp2CyB2aEQtLVWo/TxBectJDb511X9ZHIW30qr62mkvQdqpZPmOJB90JD9DjAwH
y+K1GfM/4sQ7tsGoLUsecmJ+m/AmyBm4TMgWU7DbaWIMfV39Wku963voPidR8KNE
HPsWG5VVt8ar5HjLu6UpgrqqsAYmhmelKfjS5MQM6PZ4a/uU5vCP7BpiGxaCqWPn
wXKBxJ4fGEI/3EWPyqRn1ZcosEV0J0nMKbA+2rdmyOMuSN/zmUr5PH+kQBM5PzXj
UvL4sx+qZ5y08QF9ZMwOfP/Cqk2mn0V2lN0A65ffrTi+1fXMdyefFS2TxpRSos16
6P5HSFOsz2CJb9a2HriRBNQ2HIMyPsSQosHa6p+U1wVFKP2D1M0kbhyPILUmjJXq
CLG5oG3ZBHhy9xy4lNJFcPhdv9as+KWZCGPU0Qu3LT4R1AaJbJOyeuCvzAXI8bnX
EFV/xW/wTuu13E5jjWX9U+N/jZibb3LiM+yEhrjV563loCWbbShpjzFvxW86KtyW
yLFCXoazvATL9VMophCKqGkUBkPikY4XOM9MuhVy+ONsNY2mA2emNpYTeM1wPCad
+L+0ZcjzVZb+wk+IJ9Pb5QjOgNNutR1lBvtgIK2eYd6/sTk6/PhdnL3y44n/Fesg
HfLBqrROMBXdfgF+CmiRTEu3sc8t5VVlLnb/OynfYI5wEN60jrcnp4cI6TsKZRFS
tQ87Dh4egCkDopJkTgD4yg1ascghyXTtA2DJ6Y55gtTDIolvY8HipFp2Eele6aDg
nWySURjWnVftZxZ6GTmCOFDnOr5fOpTbxtT24ywEnMh97dpqI1vKvP7l94Z7AsIk
utN/EqazuPSpIm3hV1MSNuqv7W06qS8pbmJGJmrEidLo6X+IxDrsWu1z8zKmBajz
V6Cm9Oq72t36Gvybm1xuu1l/++aONGj6DotSlf4zVQ1m+L67CQObrcSBkC16Ygjb
LaaHAhecdKAoRmzjhONQI8Wnux7orAUObmEPZimA7IJ5uvMF0CAVuGapT3x6Ym9W
jL0X+v0AgHhcLrYjU+zFwnMxmbWVt66YhuGkRIdRlKnpw+Rf81Y1rHHJb5UiG97D
L++D9UQQC05vTeSKnQtb+vqscUEqhQVUYoMqY36BHKKMJoB7Mk9KfTuRI0Utcl7l
fdtqZmDxc6cvvpihCNKdTolZsyvauSQoyAdTVIGTvZKlMyV0xuNy6Ea5i7yWPN0W
wlsiamCcI5O4o2tNeR0pE7sRifxub0ZDINsJS0dAsLhWgYItIve+EMIYINIt4YDc
+iQpwXS+trBrUMKgEklsaNmW4elBe+ZXwvTuw402W91fKnTl8FEeWoWbXzhnsm0U
npPsAReOaD1LWT1oUy3dpHDqTLLP/k9j7CPBVy4QMyUt0/70I/6G08Ovgj1+mPKf
Ie06eirPev0kS5Fwh4JSQENslA8QlTH36unh4nuhSCBAZa+me+ju/6WeJxZLLBxd
Wy09zTt/q8+7pKI9f2YXdmuSn1dBWF87p41bh4HcA3InYW0gUhFODXjbc6FFf/DJ
wzB1D51NfkFUyrb/JXarT4eDU/iZn9qHHIqtwG6dsIvqkD2ONMlgRP8lrKKYgDMk
77sMUQR5YEkMJR16PhaI7QQ9b8q7ZntsPCvSDaTOrMwjfQ7/Lyn7aVT2AddcxOgZ
2WbANRrrXa5od0qyR4s+VA2fX0UUaioylTB/xZ7aN3/vXzo/cCSjAgavJdmUek0P
sxFZXd9/+V+vxQtdBKY8H7wRkDSucNTeiDLk+uD56pdY3/HVbLE78dtEqNQXGjZC
vKIQVpZOmMRKIlAbwDv/hrJb8y/2LPGz1y0fvncnfKKtjmWH5VBDPL3u18BsElc3
mXnYrsKFHpkVKr8JeQ7eg7yC6TUcZcaxYpZoh5kdi8vgnvI9ijlP+1V3CvObG6p7
+yAGVjhiOC1R4iKoGR6TYrtqt9+Ii82uairT2CV2c/8WYDXpS4lmnFoNsrYJOFUG
VA+A6nAwHIEwkqW1OJBRB6KK1N9N3JBx0VcX/gbexAl5Ukdxt810erEqjHad3rAn
6KD21+uf2ic7o85nCJ8nSM7e81A8zI7FC6JMIEZ6EnVjpnPbghYLP3cTrv5IANIH
cZ5Exk9y3AwrbICLFx5YQsuxUdRD8w35e+TN0MFArp7CpOQLKUuAaXtfzH3/1PCQ
I8AWNO8GuEvfznRh2tuavkK9Nh6MltT+XB6TF1SNBHnu5XAZnJHxhjJW/Ee/Kakx
u+VQVwVHf2tml9nYgijFYOSUsvscyuCsl0pwMRJQhC+hZjMRl5U0ErYIKlzOxin3
28b6wy40OjwNPdzAmThuFhTqpnIyVg7Pl1MnVHdF+OZ/j/Z3cLwd8HBuLmxRcT7y
AH9SJx4Fxg7bInaPFEIR+6hqki8RgpoeQzBzAp/yGUtT7XHgZW4hhG9T/UV/7DLE
qun0f2IXkur2mN7DVM1VdVQZq1xEi8n9t5GTGIAaj6inNK7+TPn13HeKY0mlf0Ei
ICRgBo7PI8zge1XZkzUhAA0J4NkMBTVXXblx8MXzfivsiUwBhw2xOk+nJSALSbtc
wXaRno6O4lUPJ5cwhZfDh+ngqzoMnjJKH+YiQ7KEpLyYXYHuYppIh2x8xml+HBXb
iYWWySuYA/Lc27/aNg62clOoJmInVmHTsdOPVp39dvEP3MeEhCSvb1+M8KAEuxjT
rm3a9GtRjIM0umZ15qJFBq4ARxMyUL1CflBlZhgkWCIxyVYyMgh3h3Vb7L7GUCpE
u3kJJaLhz/20SGuTBQO8vm5TydtaHChfoWDrIABhi99AtXzoKFG6uOSmHTz1jr0K
LQfdn2igUEaPxtvN4FXOcdwiwws9nmhrAmWFmn2bi7v4y3qrkiB+QW+ozZWvR3dP
5yhW2MHyGQMdZIYNrAcfASXOsgFuMeHO+n7yEhgyWR5CUF7RNcGR/oyyLdev/1nu
WzrRD7QjAVKu2/S66hQNaMBxmgS/t5H7f/3a3TeIrR2gVA/MNd14hoj1NdSJ0lXK
VTJ14mMH8xo0xdGMYRxK3Pzzvof3hRGU0HeGa82aPnEK/zsBCB7EMezatkx3ZbWE
lDMgJc5MSUcthXBcXq30GB6pDL8oaIqZ07yMT51VXvSnWbDHHwg62bKX6IMuWpQJ
V1/GclDMMJ2ahGeATxR+6+QK+5ldJ6AaOVPA89yvn2f2l+SDKo8rYk++3ngEgqPq
y1rFeVE+fvLI9O8cdTsHTlkwjOracjHQWMevl85LmmYgW3kBeKMPHZ5HZYEorUh8
6FED9SLFVR5FVx8vkOFW2PgB+tngQeYCtSakSGkWcBx01uKzzEfKsWUcsLO8VThM
SDiktwV/Rb1hXw6ZXVy4kdEiw7059wTEVIqisn6+gLZyie1d6aYS7eS0bbtPYYVc
mf/H+lZQeYaP/NDpSGSgwVOt14HYDIgmkIr98vh222UeSUIUAzv65884hl8Wtv6O
m8DjIMAsmxOXnmWzkcjaEVAnwcW/NufG12mhrLxxgm0CjoUuHiLiFR3pD7A4X1Fs
fhOgrlwbhFzFavwthSbi2b8Dlvh88lK39GIGq4Bbbm/+URQWlGpb24ZFTr4gQrte
NSs6VxmGgELwiGm74kiPxxTUmWKOBvVjx3KtoyFi/CgZPjYsX1KTHqvMDUIXkor1
nErPp48bLaJXekw6WEXXXLT4x/n+whTWq0jmmosWOssswBK2uEdWMNhYjRd36ZHk
DzbNL82IByJD0AcHxhPslvbkXoa2Ad4ey3J8fOzU0PYTx5ZGvr7GNRYWK0+g9zaC
9YhqDnsLPutaZvCJaJ7XLR2pu3MfhzRH6Qcg7sdfNyd+dQ3XXNSuT0Bua7xny5jw
5W7I6pNF/ZOJrOGOTHyd1VcoxHyNSYr1P/UK5xNgF2fDiVWMcPt8ZmoVwF0CN2OW
4amfAsZqlbWIupse3Hz2oqODbLZT9DwAcoiUWEQmyiMKrPr2WGPLB9vP87ldRpbX
iC1Ee7zXQ3xpPZX9cK9RIGOuNolQwjds5DT5n/7xBO0Bymvsl/I+nouu37b3/y09
qKzjxwqtweW+m40SEeP4L67xSRQAfe3BJPAZfuqPXrkFxL7t7sk9ORFkwjIDtAm0
nIYUjuwdLJenPDQnH9WeJAKP2FbbWeD/3XQLptsTNulw+0+CxzDy0sHcBZOAyabN
49gp0StW/L22QCIYMq3JhP3oteBskfMTKpO6rpqKUIG+zLwaiVdTuektfl/EzuC5
4CUaKBxeaMD9Zhaqhyib+7PyxvSGRxZEzBKs3wUnu1fS55RqeaNefBXCvVuRIUY5
KrpYRqPAATZGnpaEeK9FUXqT8QiILs94gEg2tZsXIoG7gX7VcKjEMxr9YmkrL61l
0GytXpBYjp4og7twNidMo+QhNb4Dsb1zhdWi0Z8MU53QlGcRZ/Eo8wOexdNlzn2q
XG9KCyiMrEMa7eIi9QK8nbVToJtkunkZeNooQt4WIEMAzsglP1D0leQUfTRwT/aT
ckHlctG5U5oi5KI1twFG+9A0n5Tgz0PfAAM1veQ/p2LvsmDbk7xhkaJCyq9kCx0G
F1H0vBJhwozIr/qvRbQQBNnP+FD4jYHd+DhZH9XM/Dj63hf8yToJi90DYi8JGdcC
1EcjZKJFTaFIlkyv6Yos185/vD+hMiKnYsdFSNtwOfC1GYR4lG/oLsYd5FOY1bQ6
S5vTdY0D+h0oNDBO+e1S/qTWfStAfu2n2/B1STgckzkGiL3Vv1+gt0sunw/Ai7ne
d8IkVqa1g5S/lacg+RrxWix/azDn0x/Xd4+TfIRxDWaW3XjEEmMMXjK3LN8FrSyj
aA6WznSYPrFji1g+lO55DVY3W0nazOb6R8YfjKJM2Df00KrHBVy8B7SZNg4miB2w
ZsTFSdXwFqiC3K1e2NUlVJZR6BEyJ4MXWhxgZoH1cJBUh0v2KANFHpknbi5UD9KE
D7XnRO0z44vlkakzr7qTRFJX3nuNvHHqDGddHJw1jxcKyObEEGZx5Mw4Wst7/Z8S
Xao3DKMyLAsoS6wR1rJnzUsEXHMhg9jdU+AocwF1o3qasjL/7CssXIbg7xsUKlgF
12HZXrqDrXVUBFFGSqM5B59FpWSUGefHOxWNbHN8LWEe8ggmnvqC7+SyR/MwDR5F
3e3VSyZrga1aXmnLhLJk8TUytaCRC1zGqym7ZUzXCdXZbT48hoobIn/j3yoBMT3i
SQyK12G5ZzKnUfe9Hnnm4Y0UStkfnrr+Km9J1HIauRhKFhXDm8sHiknZ2e8A8Sqj
FfYWb/CT/FeFCyo7KWc+BrNqrlbnpSZMUwlherb6j58xB5BOravWhd6fWNGuC3sN
NfhjhVoX3J/AkAiKPqd6Jv6zFww9bxj19BC9vrm3eTTSFGcxLa9eYStJG3TovIPl
GutcxNwTnL5iXaFATJpdnS+cBq+apaBxNug/I6QoKmtOA3vjbi0uTaqqemlVmg3e
pJf6ruOyj+Nk0LZDAvFNJMFeSoNX+z7FBc26MhdvMAjg0KMWIfHTD9xn/E542t4V
3xPFe50DQIK81ZCR9RkDillT0mWUHa7O45xJXgYx5+V/pxWVk7afwmtJFj7InMdD
QdJvja70op+PR7k/5EEe9AiGee2YYraJTGRkLFySTnHD3wL9FKB8UnMvsrPIgt1c
BSxZRGNIMyJwVaCCHuGqs9uOblx28LDF9doDIXfXnk08vDFx4syzgWOlhNTTXbfz
m5PuQNvZfvx2nvu5q2iErgmUtR4cJJXiEXC4okl/4gLsi7mNWzXWE983hkqbIfZO
dT0gRL4BqJX/k0sxWBSTDswdQQJ+eQbirOWjQ2SDfH1v4QjNLVIa+z0hacY81VjI
4BSnImjfDhLCDon9eUaP0etZSsAhNKOJrtKb7k7Z69I=
`pragma protect end_protected
