// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kL3BZasSFdsbeAZSuIZ9zpzgyZBbPMJvM7qgJv9ivmJwYR8Xt5F7vvp0jucjYV77
0A3zZ9zx7JQtlPzXjlyC6+97/F69M3QnSq/Kph8kNjfawKEDFnlmvlUmKgbvgn9H
q+WrYGAY460yNGczmRj8lNkCnrSlQNneSpNqWat7xAQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19712)
AgtHyoM6B9zoN3iYfYDTp2hvpv0tdTFDAvx0roK7RlQ6M9wmKegYmXiNEgUqeMed
LxinwccOhCQv4GpPPNxU2pEJ9jC4tnDU5bt2SwdaqglOYFxb+46aju81HddNvjH1
u7zs0kV6aTa4GGnElVWHCScyp0enFvygJGZGbRxoiTT9HLhnz1kI7CcQFJqCSLLH
HnFVArSwLszeJaUWA8b8CH1ER/kdi+3qdP3ZEpe2LbuXyBZYurwx5RMgutWzRjSJ
rGjpSBXnyYMh/XrA0e4LcfHuwdWxRYWzLdyhyqr+49JLUjbPg0fRUoVaTrOfNVRK
D/2JDHN7PsnqO9z3ioQnb091lKv4V0F2ARKnbP5OH1n5qEsOF9y2nCcz4x4DevpJ
AacnL+Y2K20lsYsqSplgOuT+L3msS/dvcGIAHq3Q3P3huuXzua1qRA+en6jC+sV6
pUkq2OHeRTveHN7nUOhITyQYV2rJflKXLxrQC3FfVCOTu8I0wT/ChrFNc1ohyAQD
b8gPrIf4FgCjDTfyxuc/4KSGZ0gEY4AE332T8S9FwjCyBJJjcdRJXfoiM0AylvWV
Za+zX474zYgwC+IU6CxHxl0kKYWlgfUZvXDa1wYEl9GvtPkMJckHm+RInEbqORep
6kv8PQ2Mt0zze4mWvARKq11U+6VsVlzkkIdGc/SIeeg4jAzhp5DWTBpejM7J+sfr
b9iAE6H7Pr7Iv/rHTfSJBnUJCWutdk8wg3tHBtduMWgJsRh+y4hxTMCAfkGNNDne
baPx04XBCDrLY6oUhptBerL91W0rzRPBUI53AZcCgZV23ldfX4ysvmLNtzOrNMH6
Uys9RBdLCWIvHS3KWJjJnxieide3FNqFVfG8jgijKXXkvhajAbb1gfb95PR/VI17
3dCSMKx9H67DW+k6pCAZhwQ/tVdoXudhnPz6Vkj6YkfyKrsS6T3s3gaNw2GQan3f
ghPBGbFlQJuDsdBYWajceZ4TUJeZseR9QXfGRcNc9/LGyEGvE9abHO51oAv/twuV
GZZFFsW5BrVwBx/JsTsxefaAJ0pe6kAnos9q2h9LCEMYuhScHy/APgRauVpIWQU+
zAgJMJo3VDOinmf6Ekxgb/BrxNjltfZ8m4VytU09M71zRi3FssoOZphpNSCZzXQF
dMW7rx3Nr0hs0UWYUxmZ0L3HHR0/4aKZcYYkuMyOjWtGLLHZF7ujx1YiIDfW7LHP
W+5WUqSwhQsWwRbHFRbL9eCWve06NFvFrMfhbXDgl2rm6wYsr0oP2VRPk/x+BJEP
tTrBBeBRpOqzV5cj4dSEgQhD+U+D4tUfp/dVPBT/uhHUlwslHfbvIPYB41uN+yMQ
ytYd20gUGYzpXTPCpgdH5jh0djWjxAbs1kpCoYsqaVtXgFffo6PDHU14MGL5OkIg
c/zVeQZ1ngh7yAHsaln8MR9B3KmEVURArxGoK1p6ocXc+veM65bskhvPYHtZ4Rq4
NzIkXMXyym7vioXiDqiOhzhs14FCmYhfDiFR01zWol7P5pfEwfaBI2wkscr6KHgO
R6ATLwWgkWo6+yM6VyCM/NFWwewWKeCQs/98pQsng7G0HeV0/z07m7Mjey1O1c5d
y88JS8Yql/kmh5hiVkzz2wT9BqaFxuI7a8cQ2cXoCdcNuFy4/5EtqZg2y4cm1D2M
p/pyuOM9L0C/YfVJSZJMOqlmHzljlNrRtE99eSq80A+ebXKVBVMieRjDtYZ6ro33
hWkK/sijqpin9S7+mP4rIF9VPSQVMa0za4yyhxwZea/gxB+YAZ/Hn6qidfstQa5C
gMnyYPKkBsOCkwjiww7V6Xgo6ZJDsLSGcDp1lpCH8GFIEqyZf/SIm9roDzV5plYh
qQ243eLxU5kFBJAIbcok5uzrCBAyyoVcZ+NxMLhBC1Q69Ydp8J65fWQa5TKDRAGp
B4NxjwN2L34TAvW/eMMnzl4qvchkZHlCyW58xhFTEwBPTnJZGTbgA0VPRbXWYP2a
w60aCzqeWE1guDUOy6ln+9wkr0HXZQChGNjaDPCjjv36z0T2bUhluR0tseMq9tnb
ukgSx0fOjUR7jfQOzPGvVrsG7HLtNk/XCQuFb6ZVkbpXFdilFcFj9vTTmS5BT84F
Q34QrnumVq6fY4xXQ2O8p0piZeaRixwb+SO7gqBx3fL3QYkcmQFqyGVkfB7IpAFX
cA5FFOu8bw3RdZAyaslqsAgasxIPJRNdsoJrAsDD0HrVizLd8E5OQjG4MsfG+GfT
j++lHq6So6NQ7Dhk2h/vzjThQwQZwxMbHtf47b8rmr+lwgmbrtmBZFZZqg5psLUI
kYU/TTFsYV3A5jtpjzQnmFWSfaIDWMte5pzeAOk2XlnyUoPFWNBNgy3dHRxCwA2T
nSsl1fN5is1g8fea5tIqQJOwBxD4ckWBawSX5fGIIKJ83UJj6tzcyR9IW97MiN2w
tPc5mWHyORsz0cqVH0MNJ4BiQj3rU4Ty+MYOAn5DYa6oVwU0PcYzsztXrjRXnXaT
Od2nTyiRPh0+DkpqbjIyJhPR7GmaIO9PfHQRRGZoUchNkL2goAnTkYROdU9mkEWY
hZPS+Fq1y6seO0JqXBSQLaghz3osrgDD8WUqM9oWFLLLs5b3x3TP9HgrJ9GsObEp
tWQGTVg7K1ko74wMD/g01VhckyvsZJgRzN4mGQp8iBTvT0XfrEr1qj5tBW23DOwF
s6R4T1/2+nketBfU1HCjdO7El6b+p27iL+zGhGSxOcXDv6DlkGyhPCH9kJcEsE1i
1rsIoPhNQC4g2aKKCkQ131DSJMWgn9CR7jzRu04FOgS6lC01X3vf4j6w4vNlaE7T
gNY35LWLHy6WRK9AiRe+AuGv4w1ZVv2xOnqnNljnFEpSpMDdGDm08eD7wuAxwGtl
8FDVYec+GgPRlzVgabvQ9WOPbbeNCv8czrLMLuHVwN3Ed1Hj/U3L6/VTDe78ptEK
AO0/7gsIGWI/NPTkstPlAcLA498T+GN++ikSCCSDT+OdYWPGTGXWtk4rlNSV6XiS
Q49TVycXwOvRoKrLX3zmyj3VEeRFoSFD+Cu4L5vJc7uy0txLLRyJxSrRS0DHlj4X
KatjjKzKrE2L7Wg0D0PR4NVQGnnKMW5nMWQmV9O/1PO2j0A/ZorVuSfxWffXw+mt
tWUD6fD+Lu8qhHxnvs248iyYqyIorMXXvVkLIuoiKYbn3iWkFYUqOFZNLnQtCusb
888tGXu8ZKSKrIMVlGbI9et/e30NqLuI95EMz0F5exbbeEwKmWqc2DCJa3m99mEP
c382WGEIEBbM8LrriPFLlJ000A2gF09aG1wOg1q2LFItIkt6CL90QyhbSB7Oz5ZQ
C14xMT7NBV8rJLoCk02G2YJumtYrWThU1L0oY+XBfE4bBKSo7O4wc8KVlVYiph8j
Fs5efcV8NV7hu5FUAEBrpAa5vc1nn/sPyXxgR6tvBj8yWqD/jx5mCCRUZ/q6gB/H
Pxn+MZhgPQbGoUlzXRfKHdyr9kRsPRePLquFYaXkZB2oX8/Hg6UsEHfaMTlV5wru
HgQOQ1y1TTFsvMrVKHcWd0c0czNesD3MJBzFE14qNqhtpA20WYZ87QblXFqwgdN7
SMO6LsZ0VzMPnVUKUmxtz5HKi93oiyou0zmAeewqznRgf75KcoCZ+23dQUmkZN9M
LUGu4017Rl7jL+eFu7bWwzGyRkKWt00TXKFQ4nsLVatrrAQ8nNMs+B2iWxJrPtw2
/ID5qLog+T+YDVKx6+Ac49y67dliQ7K67vJxuVSAh23m7u1HAfVFnWz0rCfYW98q
DW6hBx84iZ66BX75S1Be/TOHJGSO7WjwJX6gGC0eYc/WpTWVJDT6DZnMBydM5zE7
NOeffVeDfGoBMAG15NPcyBsQFPr0KfKhOfxTCRlWVhRRO2ltzdWqfzCajba5cwvq
ogtr6aw+247CAbF1EuhVJDfqW7wfIwjHaqolu7gGnnCdH5m4uW0eh2eXuGV6f71n
QzeG+2yH4BgCbwwMSWq38XcRkT+XdinfJKpzcQK3eezEz0bRjLmoHIOkY/pdn9X7
6mVZiEhU+JTJokkXNfHzwGyUeE8kBs7214NFYUevG0H5GI7mj6RREABGSk1At6oy
BH3tbAneHvGRrJlLXbM+csc77Uwlqeiuyt+cYElKWqdSeAs5FHtjD+KwpJiFYMYy
Q/RZkBlf/6WlLsvkZheDSVc3mWsw9fH/Phr7wvYYyDRnTy5kFwEaPrA3+QNBwxTf
dhSA+pKlauHtcnX8Xi7Sg0B8KAWvP2uxdaURSaEbjXw0wixMLPv9dZzyuOLbpDMp
0+KZOCHePs4U4NjMnK3XjhquDotyu4DNct0pajSHHoiZvcbtQRjry+X4/bcPgp/o
e8u7lL5pDR4ddvMP+Ymv75JnWxj1wWA2APTiRIMJLaoim1ICqnz+CIPhVZQ44aSn
41kl7Z0osJ1T/R2T/Pl+YvFv1tLK/fraLHfbs8bV2pUKvLkEaBvJ+w4L8ohk836c
Z1b6V2u5r+Eoqdn4kj6wHTWP84u5GCkCYOk4IVVnRpc9VOHjC7Lf+IopfpkL+o0N
s6j/JdH1odr1dGiE0NEb+VmbSe+63iNeBFefpg7VrZrmOCuN37SnSMVYYJPS3TKk
mzr9XOWkPWnVh3RHo6W0TkUlmEByEM2sZZSHv/wcjlOcx6thwcRxAAI39lm/1Gmi
sIvIV0qDlr9ra4gf8Um6RVuc7VzHZbz5EsqIwN14Lc+NCSmvPUKCZzffJuZEKZiy
iUWKFpu69VvJ7gQerdNHsdnHVU446KWxgiCFudEXXObai511Nas+Hg1E6/Gxihgy
enIg1lfP0bEWlXiAMVVbIZj92TnrNHx3FE6ZhHBGFB2t2jRGw+skAs+PuzbS66zO
PUizVmIksX/o44cpanHj5kPUotdyikLzaszHtrbvVabbDvjkYXeAaXOuB5RsJvkA
P2FLPi95HheKJtz3aGMybVVgRvFsRaeNGnjiR5TrcOiKN4UL7nnYiXmzRikpVvjq
MLv+IEQilDviojN+8MwMi94uFLGVUY0RizMTTC5kt/KOv985jqfY+4BUd23MO5xE
jFln/JFQCpnNgNxXQLnB9JVOhsRtOIievRe+JnQim51ToCCqRQsIScV/vl5EdXtz
y6ygIi65ye+rM6QUIDtK25tckO9ySimZPY0XP3iSXkv3FQE4r/cVaLwjNuK3oQIX
wqlBZpiUhgJiYPKyUXyffm4H+vAX8qANooaUz0th4dDOq5dZXMu4ZHQPYylchxln
Q/4yVlQUnP9ucegSFdWz0byFd1J4MXzeysoHlLgshDYeHnCsUrpacZfeOcaw7j5b
V8SQNMCPPhEq0O9l/evcw8ZZKrBuryAynw+bIa7i9Ws0rfG8sFWYRWiv7t3/zaez
LMox3ur97JU9m3iQDKBk5zIQP2NOZhIHt52faO0LnVQxelqX0PNy2K2tj+uywjoA
tw/5irXNCU3eVRbY2U4q21GIS9RaDJAA0/4TasR+a0zsgg/fwbkx+J3m7SXfmKzV
xCp+AkzlhBRWMOrUUhrTqgtp3hAiFxeQ/SzqrA0+ypUYVU/qvorqo4tnjKaD1OWK
1tk5+ZRR1h0Nx6sB1YJ+CxkNBkXc2nK/huf++jK6ZQnGn55C8RAaugc0a2Gq3/jq
v9+w7xuvMZ0787WP7xYK8D8kTTpHhkclFYwlgTYvY1jjgLEXpjX0DZt/a2zgt0g4
syrbQ9efWaWLiXp2Lq9SRAynunucY3NgE3zBJsv/2gE2FiojhibOYGMbjyfZIyS+
AFgPI0b+oDd3aaTdfYVkHxHbf+3o/Hu3FD3EPWoqJvjrZlf/Bq66Baw7QRYiOLO0
4cbpGz2aAVAjkhranL95iSJRU0842lu3NCv9fx8rJz//lPjjbTj+tbTlD1d2LBP9
RaprX8UjL1DHm5w1xmT2iAMWZTfvapNMj9EfFWj/z2raVbP3VClTImeGlE7ppIly
KTG119Sy4fNUcQJSz9tr5wbewex+w8L7Kj2WnTEMxj92d8n2lcOsHA7TOdZowFvD
imqzdOlrhZcIjbIru7WC0fs85/RutJhfydCYUD6uOiWwZD4C64obJysZYS3MhvIT
c9yN2DovlWaYMDLUMQL62eAhR494AojTkoOFH/lH8gM/wd+ohmaqswEmujYZOUTy
FQhazfe5CerPBvWaU7LkyGZuZnIcv1g6ib4PtmuX3Flu/uF3XkCwaM1g7aBSUCx/
FueYxPNXbwOTTqubjlnQLL8RgPNDZ+GKup3UgLy73AP4aoAChf45yEn70LRymZaA
ivNO9aPb+45FoMFbtvNx9iD15vsBeBQQzQPfrLagCx2sQeIuxqcU3fXqnE21lDrl
cSED2AA2u+WpUmQBr719/JFOM9OZcPs3GZjZJ7/1zPoejBJJmAs6DMO42Uh+y2EY
u5LoFfvedUa9CmeBE68ptPpGNumH1npvBkXyqM+xlgBdejUOnDSb4Cth1SWi+sup
unNd15+jgZfpprAWeEyR+lNvDvNgQRk+2rzeYjQiawmqWIpiRdOQE9/zo6Mh7ySF
v3ROURYwAkiqfB+Yjn+mPC16eDM853itNQ1CUqKY43OJ0qIrZAi/T7hW9ti3RR7Q
KDaJyBEHH1PrUUQlGDw3CDhwhGTRwO43Ed8ErrW+Qex2UtiuhW1sT+TNWnDB98eU
rI+LNgyrnUmNh4p6TtoysHWBUB8xpZ4vzxMpxNiwg04R5v8S0FAsURk7nE8hlUux
3tyfx/QBLQHgW/Q3Ps45iUl3msLvm0jP7frGOKmSPpryXCfo0KoR44MDBDeIP2aO
ykK/o/VYGJj2kARZO/ihz4Gi05zh7OS2JO5G8s/YbkXMpSfjolu9LdHhj3STmLyE
2tagrJs33ZaLOttOp0uMxLaze/0NGe0NgCHuIEnS7DVYWnNzlsffBvnqvngC+gKy
hILAFBLdqYyPN7VgCGxrjPyO3NTEGP8XLhf/tTpN5IqPIMA7OkLtjSyUMHcUBN4B
t8cElFkaQ1/dpaoRbs+8sPiJ5JBourUwuRVMj9u903NvdD/DQmUHSXJUjZUGQMQI
cqnljnh2V0zaaadNeE1HPjGOi6hkmHcAHLqa1TEU8lK1f5gX3mOsNJexYubnkf+b
8DSjKkgwcSAnZYuB+uFJDYyqhoPPbu2SSSOomWfvv5kAMoGHyKhMMDGEqSvOHPV5
RdaRQgFPwODdefsHXU/jLpTso2yArUk2z71el+vOuwUrb5ogOPb0+mCTzMDFzqUf
rgT3nWnA+klxDLjvRSVVM8rgf70Xk8/CK7cMhiufDkg/cUgUPD6/UP4Jqz6dPyC5
8r1sWEfwSDT14mvSJDy8KRx/D3jCySL2v3H2+2cUyByKgSZhfHrTUFbraczGzEXZ
ohnV8mPZSHJaAu4cRwvX3tOUVaFido62qW3FF/jD8eQ/gIXXSoppMpH6/qVFR8XX
fhHvclKig5e3bfJOiQyYh362serN0i1luwcWYJ+/Z4D7wOLstj1DcJoq52ubtPYV
R6jGw7pOXgzTB1yySmEM7iitgZU8w8CGafR3p4wfz0KOrPf8E1i/yel7dec8RmeQ
qlUYqs+Ihb1vX4IHu+CKr2TXJvP2zBwvAIPfF00GH3lbPOOkJWIDdgqKMPYB7YF6
7xEUDoqArl5zmpAmkQUlEpUeOP631CX26XCMXVZEwxJ0xX/Ds7Qpw/2tmOHta/IW
OMZmk78gvYu01su6hJY5srwheMLglqO9KNBmMUZgiGkft7AUuxk6Qu+MNAfOGI3w
FZW8iZtLkfDREFHQVhlrAJVr8t8dCZSC1KvBiW0cPZq30jPHfZeoO9SGva9hMd2B
KBO9vY/4rqGThRCQR2DQxVrs27APs7t6Yx40w17MVn5UldGfIi17cbd/sYST5PKP
OEs5J8ul6I2uIFDuf+9OvD3FoeFYq+HGaOhr5UCFsgTEwMGNZ/7If0ZRsK55xt3m
XBO/Xake+n2AjoPhUyR70jJ3Mte4YL5NhT45ZXZd6u5LEOAbU+qasHfoFDuoTfsS
S45qy+l83Mr8guDQtYuWTVcFpfhekhjIDsN3Idhf1AaNHPinSjdsuGbUTR3HOY+a
TX5lL1+U2wOWq9rwgKDi1X3n/zv/kYsrT20VdI73Vhn7FBsMcJzcbTXktly30Xwt
3JLTBuioqRezAvUkS5rmrAp+XmPbb8Wsb5879cKso1wtFiNTQ7feto73d0pqztJ3
QG/ZQTTt+IkMgi4uvdtKQJMUsI4wRQvRX26LIo61PoecPdb7C2FpaWZKs+xTyRVJ
Uc2ypiQQ4pHdREHf1W82uFdfmu/65Rf6qFBHu2MQcYxvgA2jtyxe1rApUDgaiUnJ
kfD4HlwGWg3YDBU5DelcgCHYFU2YnfFs6kd7g4e2U7LlRXdCI7FSFcOnPgIRgWrm
lsPXBPmRmYm0OhAfIKgp7yu12wIoZCqCJavUNiKp5K9Xo6qkiuh3SeCKZblPH5KV
4zTJonD3S45p1mV1Hds4KEzcEIjOXeY0sUK0sd5LsMHmv6OzqM58LUoZt4oyE88K
77DQoPqELHLdjAZIIH51r+IXANSoGlBpfDwJFNKO9z3yFYvpgjkX9kLeTRsqPqKV
Wqy9FQ7EfwLra0sujt/iW2mMvL8+urfXjT+TN4ArFnlNp3CRGtas6w4JXG2By4o6
ErRUwrsS56qZkDfsssy9c6xXHsZeLVbSqzDWxh52Shdu75ZQvv/qv955SS8YD8vV
2ZzKv1tDAvpMLPPkU5AvBpRYz/VM2FpjJdbX38ECkd1LpDe0n2VTx5ImQLfdXhjt
xaQ53FqPm3Y5geQ1gtSdNG/6Ycx2QrdK2eHhMRUntlZHmZ49niDsXvLiflpT8peD
qsqJwaIl+DVZg5dgcwCauqPtrW/B+cyQb9lgNVwbXW1bRORKKG6vH4DqY3gT5ZlF
ZV8V/6jta6YcKoflqeOlQPAIDjdkouSrrAoudwjgY1f6xnhJKF7rL4IaO/Gv9Ntn
O3UJovPi3hvGiLRTWqGUXDMZU5RXkRVyDb5NYjYZztIqw7gM0DPHUcO4dlpWnAmL
mTdX0v6o7Rpch21wQIa2duSwGvbEzM8WaPfGvxDiJ2Cdpz/0yuSlKbMcx6xPdfV7
beZdzuH/QD01kjUA8kaq/PlI5fFKaH0s9nydve/QikfOFWDJezxb78VTqlLphC0d
0rbtx2Kj9lchAGZeQf0ToqVobJt/QVsBTmjZZAjM2r08UIwR7xPo2F8/YK1F6+92
8A2Z/2LWxnyApeUlS4jCZXrs1B0CeYj3EHceTZ/jFfnG1MG4WVZ0O/wvSoa+OEpW
jUHXQlHfBXjNR0pr3AKxlFXvjgJ9JSvnAA4yGt/CpczJ/NNaI8TPuP2rSETMBfEr
fFYenLMcf8NNGwLihPE3HJ0StBhSbL9ppUYB0YdC4wZ3AP8CLSsEq8ORb+hvHyNP
WsTD7Fycj8PB4B8YZHooLCYs6PWzAbsR32C3nWBWoYRUNxza6MOLxOCVfMpGv+Yb
Ubez23pj7e4GerU0h1LyyyushrEtSsqmpvaWXj5/pO4qNXYoLlG1n1T0aFgqni0S
kFoj+2hVgC5EKF39De2VNK0tfNj7nscSgwtr8zaFUI4SVFxO0i80CxB5oKFqdqlu
n0KqGyMHPizeqesUPrIhs10/jO8Yvx9OkDQ9fSTlBDCrtu++AyjX0/lI/NpKpoxZ
qjuX8PBGkrqt4skxaGAMWmd01LVavP/fhYSeUE0aYxpHlaVgbUI5d51Yl4k9d1x1
v/m6nxROX9r7+RYma5PoCuN8OI41BUUQ9KGIHuu6X1by+MpC+kWhP95wpu0ia47b
OUR9K98Pfd00k6yBRUOeDr9xjy7nFB+sZ45WFE9p6PPewCJxlYKTAqiu32E1U/q4
rbadeIwgTydyRHqQ2Bqb6vn4A8BEG6oLLf+zg3t1ZN42kGavs9ezKJVYYsT9QrtW
+jF9BFZu6vJ7pFuV8fYRu8kVkbQMmeuCf6JH0G5okfzB4OdboFKlvAQk/5w6jc+u
cPAWEZbUsYVqRhUID4+S38V/3fjSyM21IxA1Y5kF/uM6ctGE7a0o/5IXmp6+0Ff/
6KCDL6biGYQPwAc40XeAqoY4RA1VhDmEh7Xfs0f3hU2G/yH0NqXj3HOObU6PTGhv
v0GG1tQZSjC9XOc6gpopMrXc8mWpxBgnhIE8j82fQtWiCVGwpGeYpVkwI4tIfCyL
qEYst1hMjpOs5bf7i/vzBlhPkhk6nhhTB9s1DCkUE/UAN/Zw56m8tmaAiwk+4fne
ckl6Gl6whOJX4iSCHwLURklwCo5evLeA7dIrEhdcST1IXu4EfJKnG6bwtSe8sxkB
m5d01tKyCqGZ2blpMhz3APgBh+vyADb2e1erTppRaVYcuEhqHkrBr98FikJeu2XW
ceKzGSBIIV2+Oa6cqUNcFK4yNAGGeClEeQ3AQ9hKaoqD98caMncYV8ngmSGsHurc
zfPdBDjIsj+GHm51So0bp0urX6KJ7sJHoo0wgMD7dwsmuRroklf1WiIiFkYDMR0h
LkN/FgFS3IT/UtfQHflbsYime8BhiBJYBah+pdZ5jky+/gfqvFwZl4GMXI6ac1Xk
xBAh5cPGMRK8H3mpD1VZtCM6vhBP0K7vVAxtMLOUoVzUa8GSBKJinTKJZHaPXwPp
OQKIKIo9Vbq1D0oJVkZ3fKDoA4niGGl7gIShOkBBeIPu1I0+c0vKChLTQfzZSPVr
Cjp3Ahsprw+LCH1ExPQVYBxr6n0EPGGZF4wJ0gsO5voo2Nc3xbsqvTNSWtXGdavt
lKNSYMaauF1qFKPZf0czZtw9YQ35G/FVqxjMZuJZ4kq8wa1Isac6jFL/pxRkIWa2
DvAUagcx6xT2bCcjqFOQZZflit6YLw8cr2bDyf3SzjNCtY51EM1Jd5ow4sv+Fx2B
8++7cMpLzM6KeG39bWoLd7C4cZLfGaaa9ahGjdMXuuz5x4RsU6LWKzS4DHV5INaJ
vGQ7zK+ZG46Q+TgvDuRjO3utFT4GYTKkU7kwHytk0dWe+PkJ/UAZvgSAJNWGNvRG
hQcoy2B/nNLp5ndznjEhMIiASReDKTGoT+kbRloycczg1F25uWngjivcUD1/pnI8
rJJnZHESTeX0O+R83OU0SOcO/1TzSk8V5BYWT3Io1A3a4IIByYgBKvOxbs4s3PeJ
JVkCI9CrKl45B+pg1zopOQwJW9srVYyy+TY74hK27pY7tODcWIyQ3Kuqw9bWw1nw
K8ENDnebeL2IbYf1+O38o5d9IaFpkv92R69j+5yUFosUFRqxbHZgBRTgt+iAgyFL
k0T9Aof1Kg8ytJAL4Yjxfy+j4jTIfkLshDIpb02g7OTbv5DgXUVAPUCL97LWwFF5
KeMp2VznfyquNC+DMm6khdaPLXPKiNmrUvR03qr+Z44MbQWAdNSEF2CqSroLIjZq
g3k0fvEP1SZ5Wdvs2BLTW1tJb104IbEUG9V8pzoNQUNFNy2WTdUisSKmsqRVtu7i
FhURm4+1e0K2sbkKxyYIZMf7pRFxZQuZyb3rLtXzzZar53xC1oeHhstgjoQ2nux2
Qb7WDVXrwja4pyyCuieSBKE8NraJtKMSQZDcNTCuQ/Vd2e7xWyPVLcZv8Imn6tKW
1v/zg+Wrr1YDvfIUF4yRrTtpQuDmv0vJopwHAGmEx8FMF1B73wokAnzCzJZKaNCn
vdGJ8hb8hpyVAQWedNBscOTnwUeX3t+4TihkuaocgMwwOECxEsjUKMzU+nbTKU0I
udHcAKlv7ubvV2WKDrTVKJj0G33AJxL0k+5d7RmUpCGKvTf8KuVTKh4+uRnVY4je
/DLj45B8ruNzGTQiHnhT/L4g2kVrtES2YLc9beCKG3j4l+CYhLZ5pP93gFFcOzgb
DbyF1ysrrRBy+d8FborR6mmGC0RVH4rEmKsN4gHx7B6XiP3G8Jdt9g2z4AMjeC+C
6EdpUEuNPhRvAVyjtmxpDhgG2Chf7wcJbMWkPg6wwmjJ6ThSv6bri2NWmQUDZ3Pg
9A8TA15L3jDSM+iyU2A+DhSolzHIR5dbZREOp9QgD82PB/iCvfYQq8CDEO3h9OdZ
GdvWhMPZRDaCGrFwOdKKbejPJw0AABLRocxwGiOCQ38Bo7QGoXHd01N6+8ULPMzb
PIWC9Iv0s4KEbnLEtDYM1hyujZV6o+wfFdzQhMO7Olvw7olDw6nO5mcyTCOPCgYd
huJi1H1Mjkr1RA617ZcYEm7IG+AJsZeu/178qhFVs2esJbp00iAq0TJ17Cw1jdeD
1Wz4KaWpNSKegtxazaSMO7XO4saF7I1mdOjul/XlzVRFJEtnEbEh3XVpGO6OX2zT
oNf9yfKaTpMiHeYI9vYoOlyhmFU9YaB7ERB+1iHN24f72dcrBemxAyNDIeucncb+
ZKgqNIHfm5j9tg2qE6/HvO3tBKO1fAtbQtKuzdf+kh/F6DU9P6L+4TF96WqDgSjL
DJZmjo+1OGMnP7AWbW0ESF8WCRbk5mvAF1IrmynYK7EAPv4qY1V6GP/U3dmfqQyL
TXJUU/AdwHH43aNbeppqZX92lAs+Ban54jxbcW2/So424prsNKvFVkzCdJST2yA3
w9U8lpDO2IoIkLheeMENfRKzrjvCqxSjnCEYXCLjICKvkelMHxp5Ul29z63WwIDh
zxKBp6LqL9mT84fzmm/1POvYPIFH6g9trYMer6nkzg0nyXHC7ViXlOUgbTeLANyn
Q/LrxW6uCOXlJw8uaOhYGx2KKAiqo+nhtZJWt7F2UqW5Tqt8mym+JnbnQlWRLnJk
ZFCSr5030ieWvkion4qZWAicx6PPMlmIi9Zc6R1xkd4rlOQO7FcRvdX2/mUa1ijc
VCYq3G6McNILd8+VSPrGc1S2j/3RXBGgEcFeLdvtFuL9CmcpFBtfhohU8H9cdztt
IXTENChMHIKM0WFJw1vc1CpIIShGZndsKGlpAfmtFt36NV+/uL7Jq+AC7YIiq4sY
V1vA/jkNOGshHiVMmGGrG8YbPEOpcXy20+giSilL9pcQ1CI25nH/A2vomBdiicLh
C2DOEBdfIjDrxjyKVITa5wvLFmX/UXEaZYqtg4xNeEfuRxav3ulPdiN8RTD2cANr
EQ9yFG7Cs3czNn/km+aJYGWBqNwOXyOlgVDlk2QH0wOrtYEJQSh6UR9LkE3FAo/h
5+pw86q3GrOgTfgOS++yfs+jyRBjbbFr+jkYSlE1kqmSd9YhXj8cHXlARNQA7li3
6sEQ82n69YdqIXgNWp5/ssgtkptUg9n/uLyYWVT+EdpW2uB4JjFZj9jvS8GeZkfJ
rUkDXzzs6usUNc1cNAFDI1xYWEMTFLL96AO1rfAyLLmd1Lck9HeDSYMYCHunWI9e
CAlbvQ2JCiOHTzYSFHHiKt7x3xC5mRyInXjcWUkN+bfZYvIoboc+bd4xLI3s4g0/
eo53Zcl8xbiyeKkkyJnXn14sHifUgnGLzIaNY4Zef6Kstscs70Nyq2WpTyTiT3Cx
aOEAzfELMoo+zHpYsskV5XFYDJDjBSaObWqgSWXKOilc1NGS7/IIKwbxUmWj4UFV
W96TvFC0yeMrz59tNchs9YXwTpALxkLdVijCkhuNprND40cBhN1Md6TwYhPH3EqN
En+cWrBLy8HkOb36N+WjbIhd8Gq/B2JbhOhj2/thuCi+C5xEFUIBxDXberVq4UPJ
BHsehwsJmSn8wW3SToUztzdpYinCZjMOoxrhnQcQHk2VKBrTkCsbp3k0IRfchGta
rzaZMW1O2mVp7CSE5B5eWqAhxHGNU+iPCA+qA3QLjdJOqMYto+pv2lOvNpNIzSx9
MJDdl22vWT7ssXPG1QDNXLnO3tKXemk+GEucaa+YlHhrYfakJJjVa2XNgem7s3k4
XJFOzAh6+JNgPD5IXAy0ZEzeyG+I1Faz+LCTP1IE1L67ynYK6mw3lhhIli1mRSTf
XyEKlOr//qryMvkUfjWr/4g/4Lqdi6MGqyUekgsglMKYPU4ygEAbLjI3NAociggq
bg2CsVfjwclPpUitykQqTDptp6/4i/ptEmfXnmPCKMSgi94byx5ZNpKS7LC0UBvB
aIV3Xk/heInkFsOx0Lqsz06VxUxUKAWX2QyUy7he+yrkylqRxfa74fpHY2HN4O7/
SQIu2OhMfin5iXcbrn6kgE6EFoU/ZMBJ9hsckMw4VG3XyhXpA69UYDNBuNVsH9mo
o0V2lbB+xEeiO7xBEwDgxxmDaAKA/9fBeBHXpBlwz2ss+ZfPM5Ma9p5R12RjKKup
RQw9+oDXpJyA71DzeiEFe0hWDqzRBWZy+uTAVwX4dhSXwgUKfpi6Yk0t8sKUHsy1
2JIOQGGRh5Wv6KY5aBuzLEBnXibDzJ0uMPa2ysPkvWDO3COZJ0T8DCzXDO/3mdWa
8HVnu+3gH3UuqPApbkSYkpV3W0xy9mbtMmlOEF9Pd7qpdvo3Y+QrbP185uajuLqR
7q05QR+TqnrC0YGc26bUTPDvtmLAhXkESfJ1ue0gwNz3TlYmV6dppgikw3zUonEh
QEzB9BEW3nUjYK74erW7DL0g914eCokBiOVWJOM6XlxAdbAQfX8FNKKP46nhpm1P
AAzVUVRb1qKS0TW3QU0zP3+W/czi0LX0Oo/OvxFwJ7TLwPopIWfwxG6/iJEyY16J
g9aTefpKAF+4NadzVflbi2zstLxX7iLsixsiQTbqjpWYI7nQy9Dikz+F+pb91q/T
Ck1sngfaBcRUA+2qEhjZrlci+CPkwmMxd5gElF32gRpvWWqduHXtXrmyzw2Gj3FK
NhFSsp3/a5kVn4ZwLgDQgpPWS7vG571pqL+CLWVk8ED/uQKOuWx9WKvYrj8CMHKE
XXAAyoUoR7HOYuyExL+krbqAk5XIDt+MnMhPcpQ9mfuOLpnJdkF0AYHeBELxgPs0
UmMmBlfPPbCiCSXhd4pnbOOStQ9HkpSNwax4CqiWBK8P0YfZGGlOJw30siZ1PQJV
DOTbiZoYvsmIVivZfKNlic8H8JBNZ8RbNu9E3z6sGa42+MCWTwFoGFpnznYBY9tZ
XW2odtXdCcEPKbF102JKRdiZL7Idq+ARuGY5Hs0IJXqjFh4xj+6hA/oi8+dmece9
uSm5JEbP3iglkeIPCeux9azQorBmUc82X8Oafh3pzINCj3nRZ/NQPYnSljzaaMCj
gwt1GDzdmJHPGjAgLU6P/EW3X66ohgeJAAn0eDE6jCx5aUE/2lf/wE9K8C5jMujj
hI5/6S2fbYZi8l0Ewz2D6SgLp1yFJQ2sy6Osrp7Wx/KUpRHq+94fa88O7AXI8P/4
DI66WAqHbYpU9u8/7kOtSLWDTv66VTPA9R26gvX2fN28HnDZq67dZ4ZmT/aL28F4
9UHLhs+stViTtOeZcMI3CB0btnzYTNAf/rmKDZe1q+69WKs3TtheWyCh13CuiVjN
cySDIh8UU7yPZBL4/opNISIBK0Pey11xSgqNat9bqJFZamKKLZtUEdeinrj9I9th
bvaNLVXq72ZAqP7W05RV6T4q5QO9uqG+pXso+Upm+KCICYh7EqX/ZbbcPhYbgAoG
TriVRworkPt1XgD6nQ27GK3PYMSPsbJuWwea9oPnxYtoxryqdFExGdzZ2T4riFa1
fJ0MRP5FI6SQonYKxGMv78f0O4bXD79nlb9iKpoVZf5gD3anKHFHK8KRLjYaTW6T
Ru7sntEgSSDwYo+5iLEp/pkLKrcXVg222+ESHwVXtQzsq8mhLPoZhllGyfiOuEeT
HnzytgIS6eyCna2DeLsrh1hfK+emPQBKm+G4fOyCRe6RITuSENy66t+1h64GX0o+
o7ojlwRch02FPqQ9sRL3b8ztkKSc3WrmlOAoU0M1x+AT9GfWXQ0KJXFF2ABgoqxj
rr/LzvGnN5UFOEFvuOqXRoa6daw19p8aRFbXjsPlZwM2QEOmarrSSphTknnmhagJ
bJZzBM3YvT3l0qIvqhBb7OrjTFlI5RGIxCPgim/429flyaRbtOnDMNApnXQ1pkIl
jl9d1UXHolDI0HqJSxjy+DUcj4+yIgH3qssGjuUQY1DtkUxoSMkZq8wg3YuQVvHg
xhzl6yUHFuF7bRxRSMj6uBpkhAzN0NRdqLq1ys+raTToGxblhdo8ZLQQPK5lKLRp
QLDi3RXnKvT03k/lkLaoxnEHp+X5Si06uAnWL10NeNTZGeai7b9fcTORuQDsn7AD
qtXFmM3iKGREqNh2GQNfpkqAPNTsqfxifJ09UgHAvlCbjMKd3Tq3iicaNud1f3zO
c6jmmcmUY+k2EZ3HrR6Om57FzAdpLaxHHHtFC9tPoou1+xshiDPn/LuXBaokYubQ
86x3316TfIfkMWzrvS/dZqoF9WhdxccrKgHQzrcP/JbHpr+q49ELnb4G2T1qPsOf
slEPDgXJNKkQ/Cqm82LOKGqKpg8v0mGic/Y3OWfSk5WRwcY4CUgyuS0j/rZ18V4+
phLn0atuSzvdc7eE1s5yi0DI/heCh/k5Y8jsArb9WqmFScHKBu+II890O8wdm604
4YXNESIpTJjNoiD3bSlkLMCt2Ml55sdQ9kdKqn5OUbjNIyfAzJ1trky/Ix2uMJFf
+FnCB4k6ZWDyInK1drB0cDJa+asrXD5ciJ5iZysgGkzTGDsPuPCLEzm+7AGhb0tk
5anB5hJtqHVfrthFaddg4NepCguchJmQJVwrFOI1/brO8mN7j/d7dVhPBVaLgREJ
bz6LvsZKapcIRPB/UuGr33nJFG9EFdMuOl18j8WqbDyBuyrEVk8JeQ6c/7YZo81h
ZwDcrfVUf8NO6I3G2C1qhsmPGiwGHT67Msw80e0bnOY9neT6PSSUk+wYFDnk53wH
+sTA+mZzfj1Ly1x8DcorCtny9C7LUQr+fMEuZ9V3TzEhYFC8BMTkIVlpqWlI7nB2
W+GnVTbakSKEjOuTkoh6IkcGQP0C9ZzEGms5a1xPjJ6lSzd3YYPLPxO5+TaoGWEt
+qhTx6ahOG3nq+vPJ+4KzYlka4QXibomIzW9ga3JXEj94svwcrO4Kxu2j7Iv/adX
DsWQhFals0Ly2nRaIYwcjne6tQweIeGGKfzcB16c+jpVFq7wltKHSZ05hAA1AKpK
7VDjTN79G74NmZr1NbWlUtcSLDrrtGCbiC3pHI6BH8qUALO4TqAxzfUheWEWMd8t
iTK5RA4FyWdwLatp2ASmTYdSjznoLlieBbbCwgnC/qlTPOnAilrEDv2OYntODKo2
8a2C5Z5Ts7INHMnwqYW+7tdH7q8rdvCqmZAsIBwtu45T58tDHTrL6nb7KqfL+zUp
bR4IxRtn8sQZeCZs/PQR3oAE/b+E3xOaOxxCXM7OhyEomki3o299HNKIB41BI3pN
EniWxOzSa6HyuHkkFyAXHvSX/9Zjz5fjwVVizQHXF1ti/ZlJwyH5hKHcIMEc0fPM
0cR5cuPldsLCdNq0YfAb1mqp/IL8nYHGG58mxCNb4u/E3750Et0MIe29W6KcDIXt
CdPynxOBp7XBtYtIRay/oMk/ZsqXfO5JgFOe8LTxcTcifHPHj/1hI3ZnpOU5y1MS
UGgMvf05p+ZVsgXER8lCfd0vIhoptH5MAltd2JL5f/GUJ+jdsmlmn9dpVcAyH3Qi
JYARMxT+rpX4HiGsx8Igm6ExFygFM2Y53DWiFhHSZpGAqr6tdlsdl0s5npko9eAV
O2U9illTWsv+kwVwuDp5fnvPG1XrQq7xCg3T25AxV+tzrJybQx2NPnI7KjHYM95o
MWtt3mu+vRrzobBGx2RsHRImKdaDMHnopdciSWbIEJ3BBEC8eX3aSgnw74zeearF
yiW+sguojp+s8jg/5Aomuiqy2pktc8DCArKMb0cRJIFnXiE6LwEOBxnTxFmyoqRz
oO7les7Ikij38cG+41zYG7T5C6eEPOc9dNMS/FyULS39NfWMFwFX5fuu0ladKXA3
ZFmtKq3sDmXq7sG8gYBtVZ0Ddn3V3l7mAV8zubY0U5Dx5VwYTJaDaTuc2KqlilG0
dIXYBIodXpOY9lrzWjxu/WiDuwamPmA4Fl1h9MjI9duaBp48BCjnjgQT0+YmMR/4
RV8D1j0Gf1sDci4bKBK29ucNoGjmW9GFxVfBIqryjDedZEI28Ty7hIbcdF9rhwn1
jx3O2z+owNgD5MnwDcQ4gW1f/MrI0ZX0G8ivEmyIjmiUNnHOIS3pHuTwgh5CEoVU
vMBX0qMDkDY/bK6t566BkqSDodfgxcmDamUpEZHyWJg37nnnLc6IPW4wrX6QYgN2
Site+cB54oW0fqzLZNRFlKbXu+OwZ/8W0r6A5HM5F6NvRjeGcgb+4zxJwa8mH3BD
4+K2518ooCdczVfC4+ckwIRO1iRFKqskDGBjRd5IpuPC21Nj8mGJ4jN2k0wpiwih
RFIFc6c5LPauFJE33KAhin2IfYnp1mPG6AYV86lM+3Kw6PwI992M3E/ZLw2bAAHZ
Pu/af3DKG8raSXyYMnjy9hF3S4pmWVf6P1e2I2wxzbV5Wi/rGQeBQpCIznsB2Gp8
ek2wyOkcrRx+NnsGd57ETL9u9hAUtUh2Ryox2C963ADdNPzFUsoputYql6nHDSBo
pD4se6FlzcTi5N1Qs4+rPeIePBbyUkYrOb4qVkIhY1aVTPEA8hYO8SpxYw46ymm9
gK++beUjWA4QFE26c97EUisGSs2osa1GcIqOaWPH+a3RB77jPya9wuEGJ964qYPx
qznMW/v9m78xIJEaJKvcPzm+zgm8UkVdD8CRnO8d0dYKwQn03ozyjvvJj8xE3Ptf
C+nCb1WC3kSCHUI4bFC5gGgnLcAuK7CHkt/FPQcaygKVDmPCngWhUcFrW+BO8lHC
z0nCWX1YsKK6A76VjenJh50PwflzH1TxKVjvWpKFX2ToQRCz2e2HvMnj4GKItOze
JAzo00PDFBsdmgoZ/6KNPqkYDBgUxgNDiOsJPhrrLWiOnU8STIQCUm/c+YWcE2it
64rfRTSJNYIGu/kBc1rXTyzpwaC05NKJEl0TYgq7HwipZTuSzOuAfb/9JtRUkxgK
+f60ZV4NjhFHFitBQtxUAQVhfTHcdbSYYBMe65/su+7eu3INm4G9WFOoOrxlmScH
3XhWxhcyfUdEq6CPs3MxWOTGi4HqEnw/JUffs9VQ6MFCSUMKTOSAboo09ecFd7Pq
HQf2YN/crOWPYCK6jWL7yz1vFgofTCt22r79s0gzxw6iAud0mabqEtXEBgEKOlH3
OMNIoKtSN4j5gd8+ZtfAf8jfEhOt/RCaLc6YlsTobV4eznf+nYhYVa17HPJUR0er
3zfnM+xOVyuZbZrt4tY8V+usGh6Bbohoib41DH88T8S7/++or0CLq/0ZHEMe8Uo3
EuPwZLGJ5w1oFN9SCmaro1fOznOs+1LG9WYiGKOE2Hll5eJCSZkxQeXrVchu3Xpw
TZOfHRzTg02p9B6qP4qwawteXwqG3gNsG+iPdjA6DuHZg1n+tz/PfH78ZUtHlpzK
pkVwsmwKRUej1sewZ0b25RWHA8Lv8+Sip5I3ppzLk0o8GeT4MQUjJGfIAc0ku/Xy
+2n3awG7fsgoAlOa4L07voChjA9nXvRitMXHRZ0Hglk5CrMJyftMHjhZBf2dk3P1
0pVLmDY/YhOga1S+GL2VeJrYaMqUcVzlVhqp63EnabHmfEV3hqPjAyiYcHpKfdtJ
WWZoruKfqRaZVzEzy6kLda0rh7uY+JxaFe67gtPT+6l35xYY8FBzQqqdi8Nc8ZTr
xY/GiWazpspNuOhPxmh/277VZuVVPNIENxupycLo+GtUeb7aXIgDscWKnU8TyCgK
midhbWILiG7I5alwHD4sNn1A/pqC7de8mAa3s+24jK6BWdi9tkisRz8pdl4zrY5p
UD6Tho9HcCh4pPyICHkuJCL7KOF8WjUaetGzEx83RpS2+wt98ic7tDBPADQvfy78
MhjOLP2upXoV+JMNxc4jKPQo+PAuQDls7ElU61CulpHcSI34ZlfWTJIMTaJPC9tr
qo4Yc1ygPuxEJMCEVTPjEg0TgdgRcNYtRelifI0/CkISn1Yy9pT786I/RyjIpeWU
KRsHQhvntmU+qhTAud+Bjrno2qMEDjm8lV9y0m5FhjUSRmZXjULI8hb2iyGCbrR/
QQLgBlsh+P1lRFITe5jGh3oc66L2L/pDurICYkVAfVqAlIqgTXSXnLDU8bSCujgy
hxy+nQhtev+Nu35gf3SJoMyuzQhLLcEinCb1lBpimv4yYESv3yQtVzZgSL3uD1Xs
iqvnqo80buYPhXr7k1i704YJ1G8Y6kPPOCO+crMZiHa69k1PobvHGsjrjlHFsuPr
vF1HId/kzYeMv1OaSk9HHPJawtw9BO34hA5RNu6GytFUHCQbcZKDaGJHehU4QNyy
lK3fnRjNXO+x+4zw8y0EzkQz7pE084tq0cMt+MAkA3xYzqw7uMa4XrcLr3N3jhyM
b9iuoatGCEZ7k5SDbZ5aVRKS9dCw+4GTqFxJqw3qRC9jojNqhWHBI4mbjq+jXeIh
allAbfD2gqI3i88jmB8T3A+mX10lmIvLAgVB8C6iHimBh+w/ppxO0RTKkgYcpQ0D
Bh4u+WqFs7bN1fUttWsKU8bgXkyH1MElMlF4RMBDL2/uk2qDO614riKU0vchlxG1
ztBZ2Vx3TMHPYoCNNfb+kKUqP0msIktZqZdMq4UdrkTO0N2GeTEUBmCuB3Z7IZ4I
ymRyYB5hnTeGL66qYkrsiGzUG1KK+vGNq2YOCiRi6yN6n+yOk6MwZAmOY18f+9Xa
44O26DaUqUgJPU9dWgx9mV7PBkVm9Qhj+WfgqlUCWD+WACWlWT1xrajXizx4lVFJ
qY8ifDe08+8Kv644hTA0H9wjrWJrQggvPfyZdAg6I2rRlmWp/B+ot0GsGUkWby3p
cpaAGWzc/mDQ0u8X+H+yjxrYCl+hzmvUuGCwQgzf1UvgF4CQGYbysScTjzJzWrK7
vfOyQnnzE7sj4GBQt21I4cm+UB8KDtYOhXGytR0ypqML1SknebAFSwHZHyLArJh8
8jCiEZlDiO0BkB7l5X0gPJj04itEg/oaIcbOtsWhVi5NIKOF5LONLSnXZ6XmVLoQ
3G8FEJHseaQp006jh1Kpk+WCiHOuZkDjN1khGVVu2zD0hgyJmN/E9Cpn1ie7wM1N
KYkTtAK70cupprl0GSJFX4XFToIyVv6FeFMN1Gofqkpj4oCNHxKYdS7OilGeNdcA
lBHjeQ5MmjTOafyXZJfCnfouWFb8WqZouDiWoG2uPmfmnokYW8S3/+8JWuQNNWaA
nfetaVy1H+8XaZ9/UKAeMoPX/kzgZ1+SJUL4NEH7AIaW/Fb9Ka5YuW9uSGSWNxlt
l8vRn+zslXpdYTES3RFIQA+agc5B/OfaZ1/a3AIPpuB9HaNFXlN8rKof7WvkSWoK
teqaS5DqQ7fMH2tR2spV6VjSMvgSezMsag2mGoOSB9nFOPooyN8GUN1ma3G9bkZ1
enmo21BdhCsgQpAZL5NSrmytPw8F988kPuwLx7LvBoaSSPdDlDsvY7Js6G8+FedF
LbqMUcMCqFFBiCAkcACuJ5K1Kpz+KeWHjRiJEvWuCrwo69GSVtTUQhg62kRFjK8l
hTj+Io20VFnwd8AAlKyu6UT9ulKsmH1MBkY948Lq0aj+9rb6PNkM15sbAaRBdWvC
h+7VFHt3HD6QfDoazDq3OShUi5vmvNJVDDTPGGCPVsZDtMRcp4Pos1XOH66YK6YD
DQ4drQ1B2mKLGwRlK5XgAt8GI1HMISv8Yw3/ZoKPseppX2+jVw+9Xztsbr6Qf8UZ
Ddy/SSo9+idmKcyypSZ29McRtSJAn676nBeI25QoWOHoV/dWSmi043SQF9SKRcL1
Kk8RjD2L+znHhQgiQOz1Q1KHOb02s/jTQDvlq8tCl0bhMnW2lfmQy27/xcGPxbWH
Umndzy4J635YXCKluhSIlfcStgX5JziWv2nDMxgF0dhj0ZDtMYyvndBHHEvVoUNh
yWbIj6yHyscj09CQxCa/hvs7IOGJceFB3GbADwmgA5inYv9Er6h8mnewNMzT9+mg
2lceXAP/JafCRpGo7Ncn7AkPa5ZZj6Xz1sxnKYUwsgGYxVvWoOKSY13iTo/ds9Tu
bIJ9vgEGp1fSSqgmz65n+97E0p8R2sIi8J3wJwjhhVi9lvAc66hHKEhfLLjDaiCa
7Qo63RpCRGNyTAPdREI3G0aWHPY0UFrP7tKFBd3CtKknlRF0YKgCKnqifr9IA1vJ
dHtqmPxH71SqOod4N2uU1CzW/FnnSlkIJ2NuG8Fc3jAkM/zefvGr7Czbw/u6vpBe
DQyiQINmWEZUAvXkAEOuJB1TlEgHey2dxWJEbz8jqAXLTi332QXVzL3Ec4RsO0LL
GTqyRthfmp8HrrRhf13pFPliWTmnuhA3NUq4rVclu7sQcSQVKhkql1xZbnC6nOrT
FN0DAlYLIIyyNV2u3LtWYeBilu3iGH60kS14oSNoWdVzemR/MsGKvdGowGMfGyUt
wkpZL61jivdIfzY85TSdKzTqC+8bt25FkfnpSThjgXCMoUUWbvghwS/+htup8fcm
TPsAjJuLsPDZZfFnfc4tsiuBBBQOpRrKOVMPcsXdkd7qCiRWj59Vo9avmOvh9bHo
/bvbuaoVH0yDBtnGKM33P2sUSf67niMXcrCXsMVM6nHILmrSnT0IUr/7Aa6Ja6Qo
x4qTDfry3Az3ZKa/7P9a6xPMrpjp88sBl5GGh1orfJdW+6vDkxcuM8XhmYfAtLte
HxhJOlIxsG/q7u4aXEmAmraRttCreeyXbywmcLJixFqptlD2urLnbUsZLrujpfZd
fySXD186KmVNHdscoMLe7EjfNm2XLNSII5YSUSKPAwjXg0dR/iIUg+lOzfR3kNdy
bYbI7vwhpGrD58hPHImuJwS3WtiZUyHkW0fnT4tUJ5F03XmefDund0XBay+FfKOp
oJbHl3ajpUVJIUGbw7R9ym/93ZKH9DDKF4YyGcD6acbSTTuOztgz7GVLkqOHlE4M
HZ0Z5u8W+lsEfGJBYIWexpqboDSvLqst3LLc6PjfqJR27oDqUee6xLJifBLMQKQD
QIyGkonnXaN6ULskzF/CUPXg/0lK2uW51PZsOGBv3qAPZj8m44rQqOy4r9TIvzHX
kpfQFMvwwbz/FBn6nfMf3MxsA9it2Xh0Jx/1KQUgO/McOVq8GjbG5rkoK+DKjV/0
ZndADyB10kzSMZGrfRk6hC2OueO3mvfd/6LuEm4D+GS5tC0drALIYeLR3hiB9sJM
ftGO/GAY260Ft1NdG//HcnSr8pxR728W+NB0GYbX0Smgoz91qBQT22Z+1vtsI+zf
2GeF9znCB+g/P2ZmJgvEkfiPJ06ua571Th8AG4wEPVsF6NvamfcrAmniIKvm2XRJ
9CoHMUdthbt/lFej1F+VqF7A6rhlaMHfaOCO7dxlP7gA7wqyp0nQVd9IdIwEjZEN
g9VO3lDgo6KFCBW394bzhAcZ5Eo95mPtwst1W1Q4n+HLOFpHxWqObitiwgrcSwaC
O2GKGRTr9hY5TLXBsLHR17uZnj0dQaUaxQsnubAvvYHvsBvrW38E4u1XcvhVP6A2
V1eJp8EM7VwpqdEwZVCMvaXp/UHj0yST/M2RuS6OJwr0M7UkFw5cuu4wP/RiXAdr
LFFNkoP/ZVmWgUC9wEwIpx6EXvZgnw/0awfGVzHdZsJ7n58wFA7tUjtWiHJy6Sw9
V9gEnLj7q/o1zhYZu2F3fwJ57xYi3mz1HFfqc20FIlff5x+9klVyUt3pQgJ5DrKX
QWICAo+pnzbBwPa9RkVVZM2E1wDSRR+jD/kZdC3LMhdclxE2OyqMuRMEhbdq2o0S
4noFmOPy6C/V5tEGyjhkEwkRu8I3yJiblPnIPlqM4lqG3N2zqm3NUSsbBLXwQS9p
77ddwSN1utlbB8zMvopv0ZE9WoF3CknBO7Jn7KXwmtZXT/UFhFrURsEZCmWujhke
mTWaiwYdCvWSpkjkKktyH/fNwqDhPWHOXG9FVAcWlhXOW8SlhfvaDGulKO9a7nM9
xKb5IzsZ/sU5LexfIei9TCoFc5rxQd4xfF2ZlPq2Mpax46jWuL3TYAydPxw/tExH
aZZwNUMePo8ltKxrqMwxm43McnFagZcp8traryuT2DuZl21y6WW9/t1Z68Z3DYVR
h7lCG0TlqzEm8HkjEX5Qc3fKiPFgZS5DLegSOTvYzIcCH4TMF6hBWgiFQYAn24Dw
RUfpfIU9ALeDkLcCFtuT/xR3a837O5jg/55nxs2yPN9EDRdZJuI3LybYN5+oE9Rl
xBrLlonxdDY4PK8VgK0nncqPQ7bG8GI1TTF7Tn4g3elD9tGYQ2PAJYH8OBBt7MSk
WnA7uMYU6VnBRnHSj4SBB4HJjlmESfE/xzmad/FhYqi1e1jEoNBZE4f6eRieZfpJ
6qNdvpJGiZhKx086SS8fKb/cjMvKsc0VE+k/uduRjeSP4t2+ICnjdDu2A4f1pye7
A19ae2vW34tCepfoEhB1JlomvesqK4kDfi5Ar+L2V44HXaFOvEMX1hBDa0NA7KJ7
pRDRWb4MJrozg1JA+ZSJhdyTmiLT/STQy1lyLeCLo7OYs97O6Bh4ySYNlW80WY0d
1Hb0XzTJdiOVz4BF/f5XuZLA5tdCtzSOLMA+uMWj5lcfCvAp/FDopFX9RJdUj9YL
005NCNOxylw8Bm4c8eHnUU33yFQ3DLj3KdB0UE9B8i8LKVYeMbWLMXBNU4wzdPXN
/M2F4Wo7x+6BSNNk9g4AoruBBsXWUqFhpFj7PlsU8LoYDX7kT3RwaOxdLoUWB3jA
sJ0E3GEgwFw+BLI4g7trh/Cgl7dJMCugqjq++l3nOP7jBXWUKHyd1EcEMy53XaSD
/Bc6Xme8N1UmVt0VdCtp61hvNF/Lc/C5uvX3jozmdmiE2h7W1JnZmukzaxi4+MPg
Lj6CrOBH0Wrsgl0XAavzeq6e8PZMnxg6T4TVCKrmFwnd1SVJimdWEKqEq//scaaK
cn22v9gIfTLzasM75rVgaq4dKIvQROt9799Soner8oiNSXsk9usQYuKWUuTciuEj
9UnXzubsnqPNhxcqmy4wPbHHsjePxXUFAYFxbwBOddQjug6dvnQ/rVlFh8jEW2yH
at7QtagT8C2pTy1axSfWwkQHB773fULMWRNC4u4hLu/CiznoVCAfx7/cO1tqWAs4
xlHYyX4TpuG4WjGu14dyD8gQV0q9qm5MbdCC3LJALGhrnvoSvv2+ackqPA1zK+Nl
0XmqgFkjG3lhcwcuGZrAlV9ryy4pWLCQ7AlE7/GWjupDMnKFLY4x3iTmHMZKP3RZ
abuT4jwKXmyWh/cJdyzzeHminlRQVY7bEwy9UHNoUSLGYn7ayQ2mYwfyz89aqfIT
2ucJ0xqO+Nc7bpkPFKN6uUcIWIin7xrGDH1+V/m5zAmJyxIM3aK90HKzF99ZBO0s
Nx8w9WyVSwnJYIJduPYqSvv11l7n1HjMTzD4WF/RKpLNbOYueCebnkKaFCK9gosH
5CXjHZgMxv7QkaulShm4iIZDMBg1OiA0sl/qjTqFlXdv3P5Zc9Zcvv3OQFfc6A6E
tOJYULBdBReH8QxUuunHS0fcr7PCfCdeYQmWNzbw9O4LHeqEx7BhniN+5CZDIGPK
N5pdc7f2Rw7gRSjqKw8OgRyH/Kl5Zlx0z69bvHslDCGUQENpU/yi3Est2fDODu1C
wMAfDIjNk5mnwNaguS5IYhFY/DyUNcN9vOCaTFMb5fm0bSUBj08x5e24/whBcnZ/
BGsr7ipUge6k8LgkMYN0/ISTYuWwRKN6oXutYJ/mgFq00Zn3LfqLYVg2MEeEQYQ/
KTdGxFq9qSZGpN8j8l8TyU0YOtrwAEG24xXkQwMFGeax8EbG4sOQmvsJ6Y8Vub5b
cbX3inpUwq9Oj6mW3fCz4ddf3u51JNez6Bi+t6snlPdeT38rdVrIZcWhMInjryUg
WDGKvBkQxloKEFlOQgTY2N587NENoAwpI1g685UGrgGnOgzxBnDcahdhmI+ei2cx
rY2tPwFLzuMSLS0UYyiNfwbLG8ajacVSZjzEQnmPkedYsuuGL8I4aC4RfJVA+6xQ
kAs6prreyPbr+smmQu09mAJM4TeEgWkehq3J8UmaMaIN2Yegky7Zf8EWcHpE0xKy
nJ9STn/v5t6VGHKJjaktw5RRdWh0KBvAOY1JTbCGpoqBzboyChtwxQRsJzXVFqiZ
VH6xo7icTXnUm7XTOrNOZtodF9jKPyy+OfyQMPJA+9SJD/ZL8k16Rv0TcTaQYyLK
hI2FSy23GlS7rHGqwyC8v5PLWuAL1kAMBlTbn4z00eWgTm/gE25NOT0PwBCgK0nz
2Wp+hW5KLYsUHURRW/O/iv8FwdBGX35J+aam8UmuAEw=
`pragma protect end_protected
