// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e9guBE7MweUsGk8QT2kGhxSLMNqmt5Cyj0okB72Q7Pa5cG27E0gwN4bS3qnwKEyD
A1MYiat8BLnkzEPePSL5pI0VkS1XMXLBjH79iizhtcS8Fzq47bhH9TAaWxVUsko0
Uf+aW8o8ntTjrZaPUt/GKVENCpwIiNH9vgFB1ZqME/0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23392)
2dCYEYgIqoK0aVNo53yi6+bbg+p/h2vbevL8GWlN3buCv5Q5unmM6pAssZ7fjDk/
nAn/0X4M8+p0okBZzsDaCSRAEdoJCWmUTDOCVVxWtjxmeMR2XnkKNtwkazk8Z0HB
M+YjlHJIwiYYgwA2oXga/1kDdAtp1+cgS7sUCicd4jmRlJ62kMv7daPIS0fNpPEs
VMeRElD3Hf1u440Rkchck86lGM5O2OWUFZWZc/Lvp8PvEMPifC4mamS65Hxd7GZb
oIpC3xa7RKMjvpmN+8+88TBcJ79SycRKEhEWfUCt1koLLyfHU7HX5jWpsDbueYR/
qAbEWgqzOuSr/noQLdlzxJlkjVjLO6cvu72erFJySUsP8JW3ag6I1cs9p0p9o2v8
ZjGgEG9BvGmRx+ZITv15PKM+fZiJADSaz98BrHf9rg3DNwhVd292UjYF/uqEDt2q
PrNk82sYyPi3QEk8e7l6SYsW1dLz7SfVUzk9HxcMqoG+hbrUla9ceNySzQwkozQN
I6k1jmDUWFe0J+9Kw9pIgyplv5XggtFy3xhmoxrzAchnnoMbPyfNHm/Kk0XOn1WP
V4IPT1C/wmw7XSY/IUro4GSa4OuPc6GZHYzh7B889TyUQBdip1cb4S1Bi75aqCY5
CpiTMWIzoXJWH1QNo4ZszKADlvZGf4ogRwlrIBWWtSlqPaCvAj2nBMQe1dqMcHFA
EigknaimKNO7CZbSK9dGvw1J5p3mozFB6GZlKPUHHdOqA8oH8QrV/izFoeOfZW4o
SKGC6HXLMkKlwy+zRjN7yynZw4NDmV4rvwyNlx0Phz8Y3tmJIVZvHm4jOuSsWZ9i
MrDMZwCG1mSTBnd+m+ww4Vu5I0oxxfbV5VUiZXzKbBlrxINDzc+oUXOyt9/3yL0h
WRqZNq2IFr+PK8Tqjs+8/25NXNHOpUk0JiFPuFo9KzIbDkc9tlHkyNBVuuALsd0M
Fi34BUJYKEjyZJP75mrQG40T8Yy1U0x9dtiSnfghPYcoGsALq0BUSyDJAY8VkrdK
VDEI4x1ZzNanpYRCqVdkElgzsMS1x5LDRX6XlB8HNFVClPpreRuwqmRUnzs83f8P
5cU+y72aMpHsZivaOAkHub3m7hdhXmXCQhRauKV+JuKcH/TKM/foxjcLWt2WCK0G
364MLbKtyUidW0KICsy7nO+vNJIYTW2Cu1fv3/Qat+6M2vIBkCHcWzhu8kRT9a/R
9iqEg55DkzMRRmIbavGjnvfDp/fw6or+tIhBI7KbQpDn8pFZ5MDJFGZSbPC6FMSr
gdefNb4JW0cgShgp+SDdZSYNgTGrxA4RtE8zSNpKZGPfklqMNsyjimPNxxWvVQqV
zhNx7ATr8B6DtGSgDA07FmEKnrrqIVSa5QF6353dO8uUHhMQFeH0I2Hwwm6Vpoz4
CKAmQOYrgKGIUtOYCuzXcECfonSftz84JK32YUOP1U2a2vxY4XRr0DGXFX1KZTdD
KIropGvww0uHv1QJD3nZ1pjZThdBsa5mAJy43jcSXrSoExPYbqNXQ4YoBRv7BCoQ
TJkVcv3juXXXNTHRY1xrHZwPAWOfdDg6QynfimSmztDchn5xF9Hxru1I9W2I8ZCN
gHX9ewjBtre40yGN7dsqEE/RslsgjmR694FfsfKnZLInaBGCv+0DrShqD7dq2j72
6fhj9NsPiXx9lLrAYf4L3Z3lTQNEimpgWijSzitEwa9jDzM0w5/exQgaO3v5mu/+
2kxLEgb/dnXW8UeWB/ZUdHHG8dy//Y4KH/xI+XuHOw2WwS0+Zjhv2zvSYzlu1aZa
Ge/L+ZWcBiTq9BjAE2fzdKelnOvCP2AhXJb6Mcta45+wla4TEUFG/HupYUGBU6Bn
KB0NlmsM6jKosizDv1Jo/NECcQJXEI+vscOiR6NG5/h3EC+e/zYhnZIxmLhuWJIB
UB12J0sy5nNjpmM3fFO4mhbaZFBu/1uWpXLACZtiJCvTxwS0Zddtc0eFKn9u3Fxa
Eah2tY9H9v8aC3AKZ0cZqg06AhitHcuxdtPFVp9BIVl2xbl7hYhEkq1NR0hYb4ia
4toE3Y10gB4mCd/nIL1Fox4gPwFPgubvUgusJMwkdauizXld9rNoy0ATR+cRTAbp
meoC2EcWvw/wVZUh62+OYXYqihBnwBM6GzCYjmQOfAJEs30u/hcGQ4IVKA7Rc3aG
xBQ78kbvSErFZog1JzKrutBj5sCtbj+DS+jkwAdknR8ebAJ5tCiBX8csc+osCgL/
wRPWjQU+pCXeH0nCg37anMjbz8cxmSX9kB4bVbS1Qh3fuOMlAQ3C4xNlpsLKIYEo
lmaYdiPe//mGKeWka8QT1dXTYMkm7YiAa/FO/J7/wj8hAFeDdBtFBdpt0rrre/NR
5C74Hop7t/j1l72c/xwWv2Q/FbGNhGPyDZgRS40q1hzO2QDTJKnJfSSf45QrmCk0
Jct4f87i5MKDU7gwcP4SPdjBHlGKXix2LDUo3sxVxASybBcMvsJdfgIIBVbNWvrL
hsYt9/3hwb9YuoneoJ5Z5vvu38uHlcG9iHvujQX65RnwsMwXu3BAzsBmimMRGLM2
EUWb2UXHAk9uNnjB9j17tXnCtzfjMMszStQ7+UECgUprWqL5hldXtXslPJ+Tv9ZB
9J/db2k79jLBtHPLcJY8w1WvcpDMQtpEaoJ01gAtEPVZ6swY0Pb48KfCoBV23/4P
qoDxklJYDNbPkh1QczdIfPzeyNmnHoFRV3BmmGTbSAumhsURz3cHI0FnPkm2gqAp
FWSgaASDJD3A2tVo5rqVCYv43gomzWBIJFHbtD1F+GaXYRGyTPNqY4SdCmnK/1F4
krzlOxhlnvI29G4PEd4KGrYhem27W0xDXB2P6FUH9QJ+VflrvXco0mBDsfOTUcL6
ehOqJjtCwJefNeB909pv5mCARqzjWEUo0E4OJPewRLkHuaBV7TN1bYhiTS1vLvd2
tS0cnKItjcwkU4lScYha5VvmDc+KITjbd7t9hSzUlSOWSj30FpiqnCLScXP34NZP
pfWnUWEYyUpzT4+n8NfJp/ktLiZo4ymT9StDb60r4+5r/E3ZsxCoDcvm5F64jB0v
320yto9HqT4mim4p5AdvfN+wx1NUP1W+8oyamdujVoy2HLwXaHWfxhPM+Oj1bNPE
j6W8bRo4CXm0e5IKiYeFaj/2L2FBfKSnVa/EXGwNdT6J1TbFhObYRr5qbfsuteEe
ikOMjiXZC+CJdG/P1w7fDnIl3TE4SbUQ8UNz39T/Tz/JwqkCAqORWtJ8KgDjfOf6
0R7JY7JSPTgyKnG4MXdZjh0A+HpS9ZEWlZb2W9WZXBhOHZRs0v31pTUmfnX6rNTD
Xjf7btpxO4JonjZRRH7aww2XaqxI+eBHTXsWgjKhmwWkQ55Jz2wE9LeRWvMH1AkZ
RtKzCFRPLraC88DzcoaW73sRuele2zfmzwC2vaLkSfOauGsiZAJusS+PzVNW0hYt
tHVEc5nt6MhPTdejsXUQzhKu35DZzneGxes3T0mdvBz3wM4E1vcVpSu8SzcoaBNM
CyNcBDbMKHrofQhy0hPQv0+hzqWINT0l5zOJm0v3lVrI6W+1iFdRuodkoL2Rhhjk
tyiVuVWXOcT6jI2DkI/wS8JptJVwHA+VXPq0Gq1UE9mGEEuxpGu3sd1DrtsAMPYx
S3zRsuMM8xOaZ8Ya6oJkIiArLhQJXpB5nwTgN8HEobvECBtuU6oq2XtPurEz5Wif
v5Od2NDFjym9Sixs2qlPlAbJy4NhJAQxeOhA8ikZPimGOlKJVF5eENXEr2FalNDD
8IotJNiGeLuq474s/UhA/AHDKhTlxxUx05Q/lZbsACUhQhU6wQhAEG/rpFe92kd/
PsYgAgfCW+FSQ0ZPuwD9NKSsKz2YmLUPEDYj9+hW9U99Lv3kZ3RBh2WrVOoPKWtu
f6ms7e/y2OVvK93xCTdi0qDjYcX3XQpTMOd9h5dgSP9VJSWw6otNBTZRI2IqhROO
RfjpCAtpPN6DhsjRZRssqLRki6/bO92T/lv1sJiazTL/1dO1dOcFzUMSnkutFXVq
pOpwikphB+CFbra+g9h7msGSlezMwDEZYGRF+uG1NNJkeeF8LsmboIdAQ0dfAxNy
uyATnA6LJedwX4U2a36Z1MN5w1RMlIcD7W3cqHhNcLdfXYsGqTaTJ0UA5Z0fBtgM
4UWyp5rRpV90qOlwPEjSesuWHGYlpNXc0JBvLLkt4rVryg9C2mhUg9bpEWJeOFRz
Sd0kAMl5ow7/YqYQLmWSXEt7VxLTOMUSCVhrNDGc4Y4JSSl5R2DriSfarECj/sFK
SVbSpYhMdJLqzizAXey1Bv6Xw0V0fdiLYw43LbInF/oIl9EGYtcZ/6lKHAZU4jAg
o9d1MjU1G56m7fPH+zAVIaRy6sHK9vr5B+CGhPCd4SIH3dVAAw6PFhbiqpdIygeT
k2Z+dGWJDDISme9Z9+xM4Eo5IH5ez9WPwn/Cc17FUS30blfVcAWm/ebMxVizCkNE
Yyxa5eOhGisk53iIjtYxufWKYOcihsz9eZXv9cLS5aO2zyf2MPSEblximS3p+DZC
wUeYR71OEtoleJTRHvfQ4+bTIjGLT0WOHVambaAkOMWN/aPD/QKk4anIeG2wkCos
fKZIlHJGDS+qthDJTane3I5S+EF/+D/3ajf1y0P9PoYp4ijMOsvfeS/sN3Iihrk0
27Ht7jqsTb3tmjQp/8oSv5drzdWBYIXWieWgbKxuySy9bsBd1ANec8F5NyFeFp6w
4WsvlTdxq3wK1FC1XH6SeObTBRoLRqJM3F/DhH7IYThQk+O5VTPg4EYDOQnvKort
a4wtiqNkwsUFs1YEPRbOHEcZbubx0suy0+8go8SzY+sfk+Q2IJCx7AxcTaEezsUR
nxVrNIGqC+Ws1CczX2QUVm8ORXIGG1E/ctbtdYL1spDmCrg/fyXsEjBwTx+8VkL3
fL0kL1NqJTBkqME0Lo7Cd8DmPVk13UWPSRnhkyuNHLni84wJNEujq17tCc7+QXrC
x4kZ+8YW2ylR3rnMP/uzEEm6Fq628bmuWZvkDFgsThh6fN0kP2q5KYSQDeVY4LYN
naHKJKQEKs1p/9aSZhc+cXnlpiluJbqgPM+umG1CHNZjhoE145oHEpXAXNCL9AEq
pTljZbBiKL8YiR3Rj3GTsf55HTYMi6Gw8UQz26/LPy7oM3cEbHc4MfMvRN74Bvg2
LRykTL+lKlYU7oaIfidRg1FePIr5ZKWDAbFkGjsKd+MjMRxhmAYyFI211aBd3h/T
ACd6C7hdwZRC8/N/n62VkGHJIJ1zFVZRQHrNVal1BUzxmT+pxukuMrBwGYdeL26l
sM+UN7hXqVwUlyLETv08hwamax56fezf3KmWt/Q8UToyxY2VaS8YqiDUyLEDrZuZ
YouutwLrGhCwurBI8Dnk6sli+hbQymfuwvuhzp5ciMJug/SvLaHAKppw6A68vCbo
MfFtTENwvbb392+oE2e4eyOoMFcsl2yqg9MiIMGY9B4vIXJYN0Ivl0sKDak0W8Xs
SDAPFmbK/1laBA9ZzzVI+jxKJBbHhOMYLeshRtcY8jOlv0BocCZNg0rN6CHxhNOo
fOYrF814v5ATgpwgiHFZAlbIPfGJp4GLSxCOkIe7Gvgc+1Gtwf8V115oyF7roBoq
PaxW2jmwcaxtFNcJrjv2p6xIo+OwRuEPEzKT3wTfjFPK9N5S32Z3qrbliqf+dNGR
LO+P+pi+yXDJZkLWiehRxy+vrR9pdiKo51ml3qr/OyCKlTo5F/zHjWezcl3LCKfz
NdBfdS8Iy4rJF2RFqG/V4ztQKfEFi3SqUQgvQFcT7u6lhZR8Tb1s8fhGxUljg5pj
5jEXiQjTjtsVTG/d9U5uQzQ+rUwb/Iws4/ASdWWYT5pIYzPco3r2BldBDo8k0qAs
jEEJ6Np+ndwVhec9W+cNnTEdg3ApNUlXLaGUKyrIC6oD1nE542rrgfotiKVjd72s
tbOv/WFp/LhJM2Z53tLailrjRKDBEAyLg1AEieR4kIXGQg95VAhfHq6soOuAWkub
2DODkNTTrg+Jfv///InKcXMPW40+MUFxZfrM7ZhNSOzhjTal6mEzOJr50V1xC7R8
wBeQBSl9PJ6YGVDjAEesuE9QqU2WRgl0l+zscAKmpL2rXgp5qVnu73XFlV7qINiy
8Z6UzTKwt2UfVynsMcpthTzkzpetuKOyKHycVVzZGbjKd5Fba3qAq3hGGIwqB1pn
iHwJxKXVS2IRVJkYD5DPiOOFs6iY7TO0LjOmZ5UPkoVqneDaT0o7n7rteS/G+tix
AFrK386mynZZX6QH+0jKSKL4bKqXYCMvUzoCutAUaqYBqwhKRElYxm7Kg7RNzin5
bmU7nvL0FjnlapIERmEPcjue9z4OX1rUHtpIC9m+ilMQBeXvI8QbsSlffBCg7RME
8Z6esEERt8FbjCK+CF1PR3zlQmGl11pl9qHYMR3PZZ+zlRrqJe9s0TvEyZaifcNB
jnt/zcBHzrnVr4VSm++5+XG1zizntDFHzDB5g0BzVyVpEEbwrqApOHdPCQCDXmkt
fv9vZ3ctugUpFnq7aUUmkFmdQBSc7BRNgEMjWQXlVWEhgy0Lm9xnpvfmuJxo5HuZ
wF+cRQTxXP518CIIJb00Sb2vb9LD3xTrKhGGY5Nj3uS32gGjBzZpiUgOcZP87nAD
zqnaBRVGeYjMppKzPWhM1jDCmVW2iV5mKzBxnH3sUu+a1lHBbzmxDjKcEDGv7Hih
sP0Hm/8er4iPHy0oGt7fHXZqUqU6/4sbQ6sWKXzFaJqvtUhXyDhMKvcYpDkQVcch
veVzZ0vT9mRP4hnqok3XcloLDZRy790NIQFG1ma+GAWdFz3mvsUcBOa5XJj2Uxxn
1Tbnoes6EePJHHKK67l+Iy6n+KdfnuI2zll7I0M2dBz1Exh0a/GYzmqD1mFpSspE
Uw/PljdtkrIWmvzGhDRr8/kQElAaY0ieSjT/k6IwD4pzcXDqJjojBaIhBWjvkBrM
fIQJxiClbx41ZEzojopGm0R2FxHNkjCA1+nMzTYa880NdjYlFyYhIiPrRpV+ppf6
4L3L+1+BnU76Nx6UMIvCT+eP0Y1NBnE7Oc9UB7vMhqSrme7sk/zdtlK2GM1WtLjD
hL9xGbPNwaChRKqwPeGtEyyd+ctoKlDs+y1aypaibsDHYiAPzgy31X0FgIv6+rfk
ajocpK+w2Q+NbqPL0SxOtNSU7fVWFf5wffdMcUcJ6Cl7jePsPHKIFuKtxAh6AXOS
xrqoI8GhgZA0tDvyMRqjm+9LyMAB6a2RnRfdVTBbkOSELEEF4Bq467nJup+01K2H
RsxLVMHBSx7Tr/vSMNH4YExlNfnNIFq5I77WZTihm9C1p/wN6msrGiZjVmWMR38e
qK+s+c5fMtmrT42GtksY44wA2NX4Y4X4HsDbcFXv56nTwOLRKQmkcAIKN3PmPWwK
iU2256SRP7jg1wuysUXEtjZD1xqS17LbZzaxKXyYb3vcN7XUaAbuXR4G1O0Y7VCS
2jZBELLypMxuj5nKn77wHcj/KoxeEM3x2IeOQ6YzzoCMN1e+SHF+bef9NrhTw2kn
4VgXMIWOfugiWRLbRyRa2zDYgcGcMMFoeJWzN5n5RfMogCAtDtJBQ2iehVpgnln+
L1FLUNEwHVqbdGeSB+WTmvF+yPeoomARSH1AVFDFQHYorembeo4t3HFZn2dMSq1H
jroeLMhpcSJsIMi5ZONNDjT4mH+JQdHKWOk11IefHI394Xr/i4l+eTifsRCRLZl7
3/FVl28NJdOEsLRYQNbAbHOJSEWyty7680RoZWiRcx47HJCeDaei/CT7qDBvyDTG
SZrs8Yh4MGi4IT8ZTz1AUBP/TbFS4EUZ4D0IHtdQwJDrVjhMPIFIw6L/LjpLwdzR
K9CAamjPzx4MAPYB7lYGv5fR9b/q6xlHLHdTQi6zVoZfI3y3WS5FH5Lf+a6gRSxR
v+1XQx/nbS150SgQ8O8R8RmC4y8WDUO1YUjKPmKq+O7kO9lTNY9nC4t2uOQyV0D0
TRNPEHe8tc0iiYWmsD5uMZP9T2tZfOXyQRqBLlLQDqAdh/I6s5cXNsAipEbYlEKf
8YABg+A15QBDiqRaDQFUKLRJYD6GE9mKrioBnXW7I4EyMNx5TUdLSPYw1nBUtyji
fZBUW0hsOBzQHKX0nnXRtlfmrVWxj4Gs4SmwvFsPoqvPYMjCq0TN2cF9hx6wM+hb
8GjyBUSwXQKlgHXuaWkoBKxyxNUBwczTr4ar0/pTZnn3urJVLHoFtER5AnSnQ6ll
ONA4P6emwkvXtCpc+awfaTdh0qQ39ShxwjqN15mMNmGi4g7gWiP7K7z52ir8KgK3
CkJui5MYpQzH/Roq0DaTkATwjV7qU5PDxmEY9PcRmtHE7Warr5/SLbySfzec/3ZY
hLEVd0EWBcb6GqcdqgsPwU5JVdKhem/pxcSS1jDEeHJxy/5mOSrKX1XXiGhY/pzi
XwvHvTcScPDQimQk3Cz6wRt1uv452sOzUGdV4c3usBX/HM8SdTrF2JdhkorLokix
fpA0QRtob53R585Hm6UBS8HiCUSAnK3tb3Dj+9yfQ7xdA3Xy5mn9CkrZuZLI53KU
2VUGklKrbCUfcWcl0w9C51sgqLMx+sQ6+T/xY4nqArw7tXRFlEtyA/niE5Ka7aXW
knLbuD/Nz+OFKDCK8SjOJ5WBBsZ5qXuiV8Vn3Fjl+M5BiKO2KDEWC+IzwQet9FFs
TtF16anXHFopTZ/tjIjG51rolKaDbudcOQzBWiY8XvRKMfVaYJFoweF4bboHzm2A
ruEaRFlvLmwfz9xtZXHAJv5o4Upx7x9lP3bJo/phfvHCDyjvcVmtby7Fe7Ksyor4
6aJXSYSrZFose1VOMAh0N++LzuCCHAdemVFY+00Tjd/owA4bFWS/CgO9QNmty/nj
/XNoQI2JaTu/byp/dcl9XP5fe6AA3xNz58VPIfTt6g0RBCu2PLeTW+bscM8ByOpd
bhSF6Vm2UjgTdvPD4oeV+wch92Z9FlSN/YuS1DGyfBOcLSLPOvbvfv3EisigAv/p
/hG4uUyjmjdMqEGfXvx8Aw4tXnCOmbs3Ig5p4EhUjqeS0a1F1IYnnfgafEtWNrv4
IR/ZbSgzzRp5TkjcBcwQyd6inA2KbT2QRbAT0SB9uZphbYH3nCWuK/z02w8XO4BI
DgzAYZF7VVa/eZHt5Q1VJkV3EJIui5T2/Iek3D6wLogr9bzwOoudfyWxxkOSDR8W
OZ7oSuEwqOXqL52fD95Xe2xJwT33PsdFU6d+oyx0+Kx57CNBbRzB87ItewRwbiNe
gIZO/1uJNYReiWJzpAQq60UGmLnIO8usi3bFqMbMSIGB9gYoiPbW9SsHbi7a1182
P6pvkwgnpXthmm2EuSw5rCNWaqHVic52IHUaLa8a+jIN8G7yS4lBuLZJnlaMpXrl
0TgR/dShdrP4TRbfuvL0GbYewwCMyXUtLtO/Y36e9d0V8QcWWhQQv+Ob7csSvLUW
Nzb/xl3O7WrxacEQ/nQeIZTF5ZYZ6vdpGg/pukPcCcKmUj6cuW4VWfpUjJkv6hnQ
ZGgs0JiWXliEm7hIAQ0tadf3tsrqfspAjBQLlADTZPwA1jANQxkW1xby1AAHzgWM
BWW0kBC4OTATyu7XtAfta/9FhsOVI2hyNaNmuLL94D/91QOYBGCa0wtwedgNhPB9
9eRhV8ayNumns68UFt43fZZAMZLFWx0wQ2jVNwCbtU7Q0JZ0I8G8rT9XvPFdbdco
0q3uB79A5X65lyn1Exw6HYo8cv1TeWkIgk+AYxUceziErQFnLCdmqx8Tl60UGKmN
KQw3dzLdUMdnhvako/aGiWnhcyU79J54Rwo10tg0Wsm4kiWGAnMV2l80xBtYu8/n
ye0g2z27Kv+wZ8EPq0JLzK08Pr+puwNR2yALNkhRB+v5Dq+dGDd0ZLxJsY8uauUI
PE/gnpoMfjdRZ10q+KiKfYJVviQWk8f0HfpDwjenSF+e5qy/FR7HLTQ2KH9/wKK3
4lOxRAYbS9gRSDPfzOVRvA/+0HVC6qROquFeAPMDZcjv91NGURYL9By8mflWyoim
OFngzJA2bcZkhqM5rn6VR8MmL7vv73MS5bMggKYq7h+kjYjls3hynO4etYzbj+6v
LWzd1thycB4wu25RgR6w6XydXDUfRoFO4gnWM+LmCuvWf5kPsGJF6iIM80/Qi4CI
Yt8WzH2UOCIIvygmdv1jnV6x+HBfpOgIF5r2zKTnp+kh+5q25LmVu/JK2Q/2KDUL
kWOjCaarPq9aTf/tkHs3PYkYZw5Dne3S/3CVf2nA1ntfZV06VS2epDSMZJNlMQO8
CJaSisGPbW3FMP1QrvUCbVxjTqhjW7EQBpgGLHpJcU3h5ofCoFgNyOvSJP/kGEGj
Rf9YNjiuV5OvfWA9fzEf/VBRmnuTQ5FbsfKqwKsP6onDruv2XKJ1ph9mlOJg/SQ3
pNuqXHj2sCe3oUhbocnzM1yfLP0PLeo1iKQs66wO68PKkCZSZ4dmuV1QQeaP+q8d
MLs01VE2lI4df0DXFuDyev5fOiTkUkspivIV7LC+06HoGrbv/2vMK4cVryfF3Z+1
C2QLNnx1EgUSjZdAuOHaEk1wLJ5AoKn2auB/xIR7388Hl1+Pj0IA3JKhv7eAEVOe
jVj2PKeH96jsOTRgh5xwX7T9eLMpg59iHUI7ny6rTwaNVaFkIjVNi7Bg0PaaDFyv
PivUWqfpA2TJnv+NyJDA7Nu36UFIpbA9cEmmGzesAkmF+ivMSk63Dk1HYCAsCFob
hm/R8F7A8Z+jBraVoSnvswe5h3d5brer9xJF3e5I8Fxy65lxUpTQRPpRrkuNw+Xp
Mt+0kcbVK5E4Q9soaoezhuy746I5FRGfifvs1K+IjZ/VNvCQSlRTro7ZwcQwPT16
84aKhduEpI+kgJbRKHmA1p5C1U4i+IpdN97aWKPN5yMx+EBS/a1hA9xGxkvG8RzX
GJaQu/auP4Ym3QaJeMw10yTiCN8Yi2RCXk19NuGgA6TlaH64wxfrk0z44sDIxFw8
Y/621Ri0lzgpHiP3/MsSocynOswcbP79+ddFTRfH5uwWtYZPzukpci4FI0fITeq8
n3eTBXWFvnT/IU1DysshC6ag6wawSs3q4jtuFJGXjvahDHBkmybl9WWlq1DWUX6h
r39RLSkgu3DRhMEnR53ao3ao5sWvvfyk/j2/cXCNYxKkIXyBHXyCQf1Q7lfqVwmH
Ir46uRbVfxJYVNF04Uwtpyc6VyYyFfdv6LrwvLUlcRkyGmqDkK5E8mMcXW1L9PVz
0y7HfmNndlRM2VmbNkeFIVqZTB7bptC3zxK/aK2QrDYahsX/10zJW2+DErm2vTN9
rNesRYKomAfn7YQXmMtp62gLYcI+zTobUT1OL62mbKXkIvMeBZ8UHiz6NhY1zsRH
mqo9JtzSlxgFVONu5YZL74KeF+wKHjPdej1vwBoW/0vp1LE/5tJnkbMAJpi3Vp0J
TIVFKfBQ/KLUqNN/LH2IZD+SkduTWCxjbNjxzp6uvGNvjmiZDm/WNz3veOluSqRp
BrpJZdJOcrMHj3rqMfYSroVggDxDbndXNQVQZ1afciJ3khhQzJIks9us6c1+btui
vlliAlkzrL5WIjFrjLCr+T2qVuvtVgFmmdw++u9TA8JXUFgDcfOdnWYvIjDXdDGJ
2ZFYkeFoV4tdjpJ/ynb9qe6vPFefnXtWERT0ywLaMJ/isrPHrUHxc97+Diab6OiJ
29A+UUbOA7Y8QeQ8zNn0Fgs/8MCzZR9cfNSs0TNimOgEm68h1X5dXK9eT1+3EIJL
9IguiwHjXTcnVncrZYwLz5EhHy77NDUJ/u4lQD5in8kFtYmX4mQQAfClK2GRZgHQ
FWtxd22cB/0hw1afckcbWj4UkJUggqi07YZMlJ8gUmxWI7QPtoQkMVaE7o+trqtB
iYVsyMUDp5YUpYILVphPPzmuqR6Z8zHRnrvsw7tNrXPB22hZIojQgDQXycjFNvyc
ypq/Wr54fSAks+qYzLZ/ojN4ExVP5ZLegCkvJbI8ALjE8o5YMMeIaAb18ncQwHHh
mstvK6+zfGxkcqvwyNYhVBD/OCleASejKrBdshFh68jCPutY0z9jQbkC1zDXoEkS
o9pLx1sdQ/7X8w0Y2JaFbjfRBHPQgPorX/p4jRkpwRgUejudwFKAIde4b/GG5Enf
Tk8w9DX226enJVmSO7I+FIYz66EekF5DFWbYjk5SgnTWKzppDkv+ejvu74ZFRQgN
tWjU00D2Nr+kjWeNzGeuzj0aifKLAww5QzHREKMD0pEJxHPOgYVVj7dvPJLUM6uq
kzlLJLRykjOkJJSHvgvjKIZWddIHlzhdn6LqIhX/pk+nT/RMKvnhYr7ry15Y9Cj0
cRMjVp+XR1KBrZZUGaFN0zVVAwqosBTxP4Zm0Gel//srlu/8FRcA3hspmL6iXgVz
kBHr4TCKJeg5InlGh51qw+wjScbZgGCCcBgZ0gZq1dm87USGMv6rqaJLDMhsh7LE
0buMPYkTgmMZKgEPAIvsJdr4KAgbPCh7mkhDDa10slmPiNGB/3kus5CEJXx1Fjvk
71nASTfOFoX6M+4V8lz8PqXJgXOBiZ1xxD/rgUEs0VrfuvwxEFffpsVXPVQmFedT
CUs7CSVz6LKRWHtLdDK6GzOOKVGPLXGOuvBwM3hkKGNk3n52+DnRhwkYwVhbNfgI
RBU+2z7pYp/Jv3yvZzoSAQhsvAP0VdCv3Qb3sKHufLV5QJWZ/HyLM5+B1okSihmd
DZeNXQkkrJbSn5tjsOO9ynPr1/JpaqaYFIOa312jye/y3pr+DrZdaFg3y9efw/Ee
MVKtgBvqHmKHJv3u9yTa3RJYh+ytCv2JZZPSdThZ57tErnCmskNKMbbF9dDoX6ET
RTr9b0bj97d0IQtgCkj7ElfssHq734YTfO8XxfH5PvH8ZFG4Lry2R5pGaG+ZeOvW
+BvVfNGMB9oLDAZnptRy/+Qv/+HK/28NstL6pvUtnXj9Tw9fllOcRn7pf0krPBjo
HCxbyD7xXQRpNYrUn2bMoUrkAo1jUjkFemsheMB5NeUTh4qPuU6wjRiJFkVi1AP7
PL/YCLSCfiRyBXlfpoTCcSQsZSlIfa4Fmvnj7g5+68jhDg1UYefq7Pvia7aEsUzI
Ffovysayn1/0FocnHqYX+ohv6+iDyPm0NgVJlUJdcC779iVKbvOVhzW08pljSmjb
2to7xxrlK+2xKKwqPeh7CD8QHSDKjvYFpAHWxIOAV0AVS/fj3jo2d/1aq0Kj9cRy
2U10AsLPeEQvvv9bc6ToexgsFOqpTCOrgPoTyqoDZV6d1EwDG86o4hV5hcCyl9SX
XUW/G1U69qjn0du7u3U91YOWbWqjdfbGYKfTc8SFUWngTXYiZJd6EValZW2ASCCc
VoLns87XWJRIC7EyiiT9pN7gGnpoeluQwCwHzQukpIaNDNbg4HKp9KLK2uV88dyT
eMUPPgn4BeNny0zNFZ19OHJN3pu2l7wmK/baVW/ZxLylyVejXMN6fOqpiOIi9aGz
uCKRMyjH+t7sue1D5Ccl7xZejiB4hp2sdI3WcXJ5XkZm0rQ4yjuqWdV4hzACGkAk
Ydfbx5b27oX/BQ7OxlSK3ASvgWFost/0kHXvudgWFCTfISTfPbjDwVEHBw9aNpmW
bLFqwQaowBcVmlc/q/wyg+5BFzo4ekgYbUg1LIfJAGxIxX0iqr8VTfCYwUGaGoNq
OjYP9Ope5UezkT5ryiJL+YNVWIjWnsd49t+pj+b1Qfsiy5Y9eKHcNSnJjkCnS3sI
zlc8VlRbW6/Roh9znouVQMAW4S6exGMxmiiI5M66Kt/v9BVypVA3OakcKBuK6kPD
z4WnzIn9y4sXP+DNBb7j2EA8U0zemKW2BrqiKa1NsPvKjQWxsTGQa3vfMBhryZ88
lgPlcCfsgyBF64hQy9rlQbF3CErGZ/UXnI8Sq8Iq3TtthTqFqlkSTrE6AwODDYY8
GF8TEevEyKqzbKtIxoBoMeDdt7+wO1HbsIDTWgU6+Ev9RP4CJRaAtmBG5liCDdpX
7EUGfmd3VZ3CoBeFMWvmvA3ZcL2dw186XgrFWfoeWJcH/9CDPyoqJFOvAGA1fJt3
8p6ddhUAFCsZ3+mOcqLGc3ZixpPSqxTojl+BYEDPleisI56RaaVuuRV5+geLRm0j
bj/1+Xyg++5SjNReTQvx4yYKL6euQ6XChmwsRCxd799ettCEcNK4POooLO2M1yex
uPPXTSfbdNS23zaN16YsTBXW1xJwoOes0tIBSHirfntBUp7aNBA67nNp8OG4GPao
4bzXZnNeWEw6ZkWdL23bEQ8kFmG9qf7m2mfzwYoojeL9QkqeMruvlqcke3Pce+9o
ArfrKaOlFpWo/OApIK5mhTcTqEfxC6K4T1MF6tpti6+mhnWtMu0I+mJQDGk3oUHy
qkV1TRrvp5DxYkEIkgdcCsPPbhhH/jsAOkJI/IZOEhHKVMkIMDuUou/roSseqxJd
tPb0OqfKZyb7ebSjnmDsLWqfuqB74AyJMPwWwusC6S5przqaGuLrbtgynFLujVL6
pwuGaOd599eUmI5a+WZvxpPhrIyWhQFlzotY9Z3a45qyHCKSufdtSaSUH8n4xrFZ
9eP95DdsCMf9Sj4iHIt09DFK16FdPFc/0b8bZc5YGKt9v2z4CMNLGkwOhsjQzTJw
WDnVgpIu1QeKougaAr5MCx5A+sKKYcpXuOQg8Gr+y04ZAweZmV3o9bBMlA47A2S9
eRtcbKSaAGvOZPlQL0HBah2rMgsCZd6hZ9wS/eLsJHRzBVGNeWTD/Kjdnx2mpTPC
4GUgN5AWXYJ/Y8uxNJlUTb4u5EqJwc+EX0G59SAg7QRRs2W8fzhuinklrhVFvzra
PsYz1wEx0mAa4wbA29gv09+VBWdKxqLB/Z7UN0KKD7GXp7B9gOcxPhCcenSnc4y3
I1OqWClLwIRe5iiWNYbMRO+4WIQQBox6FSnCtGt7v2cLCw6QHlbnIQauIDyjyq/C
Lb187Lox3VteeRBxtKWPtTLWzHSMK2d98L61y0///sIXNBbLDJYrluaZxgXWKMso
JSNnr4+IOQ5uj7r2J3NWK9Ii5JtxmAmVyWcZZlqad/PpTmdSph5PtDuPDkN05ht1
2ZLQP/4CGq/nJ8ClRWCKD14kNqVYDxUEUx/vLgI0dCbo9gg1x7o2gaJ+PaA4oRuC
Ueait9kgs5NbVBb4fvY6RHChiBpGE0Z9d51IhJBDaUUUeqiP1jHi0ecE6mVGKpm4
oCpCoLxcukFXhguyCpv+KjpB9YnEStOuUtfpGaximxOOkxly9srNScZOSFaL/lCA
rjezoE1Rnv7lGgGLtBV9W4MQP6HhkYaBj6O3DpmiQ2KuoWVDZRT2rQBxw6z9XIK6
25Csj8ZbRxRVBhdTGXbUMBy7VgVJs+MWHhKwFS7ZguAe4OMUI9lmwJtSSmtkxesY
0UiOVJLQHsge8i5BofRw1uroLaxZlydfDHxV2047fKmIda8i3RD6awBctFb6grcU
3nFE4ngx6KVDBn6R7WiCbd9lIpSLmlxFyNSLOgrT2ofynAEQVUOikI61lwXFlJAW
Nppcy2tKFnCvb2rmPGhns5piYgDNie/QlJyGbu6d2iFKZlG2aHW1DV4KTOtYa54m
s3ZDTEGf+oIukj1QtwsNpX+zQVOWAv/eaQNW+vOsMZwECrTQptwRv7NwC0QxnYgU
NFm017wPzMXSOwvLYKStR/R0tKc1xFO5gZO1GI+LZl7OrgFIZ170jSGA09jY6bo2
IcTg9vt4WwOz2TXmBMRK30uan/32vXbBcI/GTicnrx959AQVrVJ6Ua/Rkc4I2mbM
4RKYnrJfN37sJX4dExKCAXoO7GdtJCXChYXqyuKrrYzFhtQahsryPOM7sQ8ot8CV
P4HvcxIbXGaosQFFSu4c9Bavcnc7zUOyicdBM5t8PSB/7tnZKFOy8sqqR7B1vR/2
WCJ7epZ/vzZG5PBqIYVPLiWkkAhr6NQqASPl9J5+NqunK9ewAae/3Ditadn0gpEf
B88PAb24mtBFq/eBWiHyS4UxvWXyRJ/06mUsZiVYLunH83uuMOjbyLhNREhKS5/O
AB1B4zCQR7L3dZEDJfz3wRsYWcUkiD2RI9Ta0fjr/c/0ByZyeFFGr9FlgQe8waCi
TWgJEipgKNwZmi2WQ9SKT2frtuceIJSSmRaLyTVSDnSiQDbUmq4WqW/8w2uuZB0h
9OuloY0Hbf6y0BWBWzS0fDvQoeHmmnWaXw66Cmoy/bk7KocFRpWMuv9DktLK1L97
o9MSvMmk9M8gzbYBJbzvYjPYTzJuSbA+1KtW0KEG4YvgBc4GTdEV9B0s88mRgOMc
To75tfF/bSr9MbnCiWQ1Dk4micLWWRj1/AlqXVTkWKaaYSCQoaJkUOKLcoZE+yFE
crxD0duse/JRXFCrwnKQIAWDHgZv7lwqSWT1rv3I2drx6WGZ9OgnscG6IikqQrDg
W9cbscT6HO47RixvFcZBYuBTb/DOWK0vRVviNlENlh4yVbuChiBKUGwV1UIRE3GY
4XbEp4tGPEnF2LBrpriGM5AxtJFoPoO+pMBY7JKeCBJTKCQxHqXGHsf/TPdEls3t
mMp9TqYEYIbrdUSFNKrqIMglKZfuh89LlKTncG89ITZ7FQw+FGsPJTTJe0qZGMTh
denYrKfmgHJ8g08GzAOq6rI8UBsI2rkEzcWDbcUtZn7jrnMv5q5Fx8Ruk/UHmJCq
dt7N61YY4RdF4UKp2EXjsw6kmggGM9ch4gI2Nyb74cAFN/Z2BF+eY3fOhk8pJJio
xrcun1i0DXlblwt0rkrNy6nrPPbIo356J0a+0fURgO5UDj/zBVZWk0IuzrncuGQ8
jkLsDKGNHuZhOeCV9Y/OZGGWvmbRRPJvwpZUlRsK0gKJVhu7A3+49LZUxVN0fkkp
Xxb4GjQ/ClmeDfm1YnTryMVOUKvDvw2/lqG9W7Bgvo41MhSmKmK0HEhy0VcDcspW
Ca4bCmc+oXkrnzJI+A2BnC6TdetbmrafoVShAhBJntj4uxgXQaS54OLm96jJQD2i
mAtpZtozFxMG5aobwHIAs9UdhjoTVNBVnvzl8R0sO2FTQJsTfpQE1zwSdOdVyFrl
brjb3dg2P0TULwUG5MiYG1dd5Hftk8MNZEv76bsdlyBaRNw7iLhqB0ed6p3vxN6r
f6GNXd1P9JasEgaWgggpNFp9l0+9cerRGP34j/tnliwJb2t527OrFEDMvKHf48Sg
1eaRHR06MqOp6beJckuMGKHFb52xCzp/gjjdAxcZpPS1tzoIB0PlXD5iBKRwvZnw
qVjFqFnqtlhOLaPI2BqT75c4MVnWanDFUIFdpjibN+dZNPijE7RejI0txM4bPk44
+5QMfMPAU2yUb/gp5lw/tWlqbcyC+6GDmC5tp37zhZHj6o2LetbtCpPeimLzRFwB
Kp4mGr8EJlvOMrQ2KnwIKW1e7oPXxDoqwyPuvVIKlDeciV+Yw+iraeNMKcoLA1k3
/965HdoBSUfBEr5S6IDiVcvj4gx9lyr7XrCnKvPIp3ZPuDV+RlWXnFhhtZhhWTs7
xIlx1c/AKVHRGuMKOMnD+zXOu2IH2Z190i8ZzK9qb02uyvyIrzs/zE0AQYik61bT
3AoFdOSGtd04HiACnHsPdhCksLJ3ggFIDHbjlv6KyUCDbrmGgC5v5iQ6LGC5bori
7F4e+DMheHflUqagi+gQrt8/bQXCgw2yCP1eMVcnjcSf7FT9HleUWbRaAi9U6ICQ
5s8wAh1F/cuOexXVT+LE/+jKiNGDZIgjQzuHpUo28bUK3rDqKslpzQWB2px6cfLz
nCijWelInjAh6nqY4s3qIzAdtAkvycjBD6K9KXKOv7im2YWPPxLPaGmk4ghiEhdS
8OhsOYc+vN02e4rIpyNrjFUCYw2u7twVw3/yAtK2+PDzGzAM0SFOAbmUTnCcml9F
gqJJSJxRzL/Y+YnY+M+dNlZb2Jw2TVxDCfv/dAz7yjPP73/WbhRxlM3WvhaP/Eq2
PPC3vIIoqro3uR24ETwOixLK9ulqX4LXLDarJ5G/flwwxMLOFC1wm5RP9MnceqrD
gyULIZ5CoGrhbf32e0ndAERpZOvSlOzIUB22WObQdREWQc8ZHtZvPiDjRygx6sj7
yK0aZGYVIbhK5N8huwS5JyfEsSZhgqr+lGYypYSxtg444YNPWJDP8y+IstZjQ/rw
EUqu8OWXbFjl4+OrW0rj71tZcjg5hEUQesJ2NwGhEZJ0CvBAqJlLz5MYi86BVtHA
+EslJpmyI2A2YI1JckFD5u7Yp6W8WD8l5JS5yCQlNrPSN4WEy/9F4DfNQinp8yq6
4XXFqEsozFSh2uxZxZqLnFZmgSEFz+pukpuL/YL2s4Kc9RlcPCyb7ih1oKfCmySs
3vjoEA+dfI7lm5vRTYz7pJCpnihdg7HgmM5pP4KRfVHYM5aRQ4wQjlSf3LuCLkuf
U4XUzZHKVs4wTgeHqQ+RbgriW0KK8Ksxecy+AN3rrygZjkpOZCsRkUqvKxfOkNkr
Z3xFh6ito5kgSi4VivVdOZ0vgysMbhDJvWahowQrgiYJqFgjlmgQ/oNuPy7aNJoW
6MPUUURtLXPpRvjc0hfOKHTs2BXge179MVYsAKiBNlV3JjKC1iNv3y/Uafi7Zwq/
I42cyiJvhBNxXvcI6U6PNGn/5iwHxkTe/23nM2PDtCFedlVx40JUqvltjJqJIBTq
lL4WzZH10lahw58sX5+Q720YwEh/CahL1REA5iCyWvzV0f5PKhtsLp0/8W65Hy5l
89Ewmh+OyPyDfzNAFVRb6f3Gzrd4iwkaiD/kAZPp5oazWc9khUhnKRhIq/rljWEx
Etg65VYYKwCv8Y938USf0CZV1RNATQGW85bwjjnZBeNWzp7DdTqlYjJPZLVVuWuw
CRT++T5dY++SxSlw5TnxNBNR3ddl6LwLpN2D5rhjKwwXLlY4Rn1/4f9PiHMf3h5i
C6KKjKA8Z7isNaXB9OPdTzZ8vAv5q8pi5sLdSmjf0/pMiUeeILTlcORBCDHRt/Ui
jfCzoVRpXVMUM8JnbLo0Y/zhhGSYa26FavVtvjDc907R0kxC4CBqu/JkoeqFeW6l
OKf5C4sZx73geeDrDThi2G4wa0EpIphXodP0O2X9jOGSp/DGKN+WyQmebSis4qSI
LM6GAyT96ZzFAyK8BEOvZ964HSsaDKRn33mNuUlLlZ9RMXtwMvsEd94ESAVWy8t7
68heOM0SoI/RDJvm4bwGqQ5dLc37T42TX3OIMsu9gWtYqAwK5B7i49ukmKsJBGIm
6VmaVWaE4LsEZDthViLNQ3OnyIQoq7L+5QiZ6DZSJiJxoTv+hOoFXWkpc5Ak8Obl
jrX/VNwzqyx2ZsOB4YZ6ijY2E2EBCev5b7nxsLmft3bALkuX6tWZy8A7keLsr24F
zCRRiZ+5sl0EGQ3E8QDga2QoDJaYB3xKwDWvOHq8KAYdN7AuSbhv7/GbiEswfeUU
Zmit7mKq0TqUqNSAjki7LuwNjFqWpe9N4cMwZmRmEL+D3y2+b+ngYWITPXb+Pbsm
Yz+sIHETcNoZLBSfZXNgU31E/b4NWFTgEWiWn/mh9SGvdZc9vzJKJjuqUHxp24JJ
fXWlMRbiTJU0p4WoZNXpLRXGAoJGHJhMieDcj+AGXk6TM1GFCmhFb7S3tEDGJZCb
GsZcEEorR1wf5rZtBkU8tK9YRcyVMp806WJLBEc5vYMBMw3zQkti3b1Kqw6uQMez
jonAJrq+TZzRyeN5zsYwXoeOr0H6xVdTocoAIkFUEh3GWXdZd5L8H5xd0MoK50Lx
534Telv41dIE9iT8Ipclayd5KpMymIcSQ0SpZ5ZH9WEDjfmWUA8/CW9r+qREkUDO
QfzfQr4nxXgth0Fzf/W/93DiKvwKLbhv/hFisDsVERoB3j4/jG3co6sBmeuCH+mY
hRZU6RneTFfLgS/ikHPgF1zK74DPlVoFi1BQlHIY3Z2isZfH0kUv6Xwo/0xZf65O
a7h/GmM4/oyv4AvihJ7LeQY8x7RCcwjw/hyYiaDVIuogfpYlFX4gDMQO3cwus+OK
1yKpMsDJOrHB5CzCLU5ACsS74JdeLy6Uv0KpzkdhZXdB7qkhr39vU/m0fX2EnHX/
V2np6Uy4xgTDH8mKxMqUkLQIUIsmOCGOMUXC3CATwxsafN8+qW84+0gt3OpaWcwm
RzVuGQc5eAENav7iKLbRKRSIvZUX33D91ll2xIVZnMQgYbxP+/atQ38igKdusNYC
TxXL4KbcQmaImy6qNwKF4EctX4J1/XIcndTVgOLgD1wRr8G7OyTYjGOhyk0IrNrU
aUtXjxK3OmH7xte7+OiUIzwivBIY4G7LXSVs/zmImB3KSO9R4+DTEokzCQ+aX32B
AWpVq1YJyEh6g6HxW1eIl9a/frHMnElmDYpZs3L/m9XDBYhYXZ3kzY/UieLsplTl
M+CxUDy8+31Q7OqeKkZEp6wRmyexEP7YiLRx8FGiKoZNueglx5IarASFv1k+LRH3
l4imSV0zHTkISlClF/3fFAhL6edyJGzzb1yZDK9OY70tWoIhtKc6O16ocK0QUCLH
DAclxc3wmbWmsvrJJS5tdUk1sX2hvTkxSCTViwsxP/WPbbvsw+EMC/7FF9UYxhp9
zGJtmjMOdG5noKP3o+og0WstGXNuFSrBLHYc1geA17e1whwqk/CbiU0wAz5bRoG0
sya7S3gx7AVMwNU9ar7nWIyPjwrDGC8jKFN+R6Mc2w2uHVGx/oeFbsK4LnzkFJ8z
OTiqcSpYIJNN/5KtNgV9HflymAx1K70+kOqepEa+vc9ek1Sk3NwTvV+DO19O0lHX
zQ3/0Qw8jqHM8yE6B+y+WUUGGMe+D3wsJN0Z89mDSdskcNBsdALeHPnmxdgIQweF
01MRTz59daQqlqnpBp9jygGqg+scv790CjeaKdnMX6n0LkLNNwjc9a/wCv8IEb2C
D82h+pLrK7oOkqdBAvgXJZHCURR59Rv5XBkxU9gQuZhfaf8VN9CYS3jKr60Vj7nA
4R9D6VpvWnYbfgu7MRrFrjnLUemSHurj704ytywP8OI4uUhgCu3ev4Hny5y91jhj
2Zykw5I4OxMuuapbH/EL7nYTRWHQuphKDrAZ0msG8bCyPp5DWnBxdRaVAgeAkWK8
AX5gZphPPSVJ1CqfKjIYNKbt//hGL/u4i30fRcqjb3/QLeqRzeXjqAEBBAi8PugZ
OMLmmuzGosdZVL9XkjHOVqjXABwsF4fnWH2A5dkXbsk1CLls2/WYrnZHsl+gR9mz
FIQPhNJMdg91vLtHRzj+q3ufLYYSP8faHBnOjfpl3Xj3AKURui0OPOWMDLCJWs8A
5XIVUcfWG0WJeKVOkw3JxiOTA3hDTMTo8MFcJlQem5jsq9qf8imVuc6FSkw0ucdQ
YAg1V9TUkK9OpEFEIDFbcGXJewPEbVZjmuspQpTHZL25oGa0p27W71dVgHRQcfLU
uGEqA/lwAdt5Uv8pO/7OfoGMMqrkIWDffhNhF/bPkxASjw2KQrcYsTQysKuU43zi
pvg9bvcxYoopB8CEOuXU5UcxXxsz5kmTxY2Q+pzsWnBDAeeQjBGZtjm2Syk24LS+
C0zhzittZ3ysY1YaKgZdpYlJB5kVe9t071OnYj0NBkAHSv/H+2WR8x6sgprOIS4W
jCYp1nf1Co+dBJpVDIpecb+ZQyCRCqWIu3oKQ6M5cJ/08zbNg4vzehimPmN8aQ89
JvT0/AaDkgr4mszMSkS6Q1HRH0fpAzTEBS/HvepE0oqNooZOPHSISCudxB23JwQr
GKHQzAAzctPubWVRv3FLO8a2ehYoU9DqYGw6Pioqx+/XMld0t4rRQXhJR2DZDUGR
JkN/KPo62qsCP5dHf6GK1/jzso3adyuNZ+tOVVJzBCDi+kOAmCZpvbTPpwe/4r3j
D97Q3mPOe9TrnnfJwZ6kgkQ3d6VdMfmFSvn/0dPYnj9O2eZFVe8PEESH7nyUiSiI
VlAoYoWqc2vL9ttdsmNuuITMxlSY4Zx1lIFumUJN34TqNU0IFaOftbEzxjk2v1T4
HXlIolNhGqPZMoYUv+mpXu8XIzFp59xQSLQQFN6iFqKhG8dDkdFL2Zov+OicIdOh
czQG86bVagrCzzM29Zp6xO1vuMwnuaMI1LGza/NdRN8eWZ8/YcURuoMmowww3qCG
oyQFHLnAbjLvV9+XOxFplPdDXmS5a2mqb4FLmUYoWIz6p1G781zOPjNzVHtcgq/R
dZhdvtWOyyKnX3TQA1qdHldfgrpP6879ijFrpiAHdS4Spxte63aXpXBLDvdcgXPB
dE0xs0mhWB1wEN5lD9phcwL7r2VNY3a9ODSBiQ91G+GKT3hWm3HCom7DK10edjei
OBbUpxH2dACKhteJPTxFsFPR6lvW9YtHcW4sTHqsU7UO/3XS1Bv2tDBNfCMZ4Q7V
qSj5KC8cuZVyGiGW2kwYNroMQYGR2yo3c980Fl5+zfXEIvs/RRfouQ3IOZAP2Shl
N3WG5jiQsYf7k4kYA6b4M0ko3tbZwzEe2FBucBQrMXrK7eyQeSYK+JgLE+FuAzQ/
OqYjpNK5Dkz770n0rDhdU86saRRNxsj/PlZE8+y6CCIDNgE1oMX+x2dyZCotFAll
SUlT5jF9ZBIpvO016HA9AUBwqrL9G7I0yqCIWfIn/aQhF6tT6pr7JNvI1Xry1uzk
yVdHbDuhApE+3OkKYYsbNym9CukdElfGYGI/tCwW3umu6MK9VlVq5eDizx5GIseG
YSmj75Axz8cIW1uOs9d7bPsooUiNbYBrjbZP7Tz0M2X1SgxqQgIdNUGLV9kKpkKv
LzM7gNecPHXm3h2FyTBxKbk7P3VIkvRduy3+mRL8HD/xHI4VD6sA3Y+ipawq4S44
mJiALvD7g1s7ag07WxMJS96XNDth7jkwI2+sPcTSSMfDSwTbXeHSkG0IBQVE06MK
t6c3RIGxCyRdwda81OY22Bxu0/6QeaJKhx0KpUK30Ss1HaXK405F7TUVnX84NX95
P4mY8Z7s+XxWY8VfFDx0fz8xtMc4oTim4tFrBwd7TgvTYfx8iutPA3LDWNX6PuX3
cneLgKLGDcQ8JhRFGcePiVKGXO6D8OuLQthlTqljH3GbkmXhc3qzqgyIfzDvqbMN
GCufiJeh9vvUiQMiO1aPVS7pxTRBGOPamibfkXHSwTgzsuL1ia/Z1ku2Dlale2pV
FytoCH3k0bE+9yCcD/s3jQwHUSBibT6FbNw/jz+f7y8PKi/wAUkwbudNFICaargc
qsW3OlcCHG32VcYolRcep9cRcuv+C8ZmlZI7t609Q2Gmi+5HDx8LjZzLACmh9scD
20kkpH/RpFuxOpBJkFX0wM1TDljeUzQLPfj6B8+U3MRWpE/t/VA4iQJLRUQLap3b
yO+Rh7dPSXV6IC08m9PAVp4I5cI0Zle3oo6VgXV8Ye8n033RYZi6YQdHGFVaTiiF
Sh2hkD29ua8CI0B1ALYEPxqbc9z5B76WrIYlu8u6TIMgpvxYsGOsSVyb/+tWGQSF
iQZ3vUuN7fxUmKpAfb7bWgQaf7/iUVT0iwZj4Gnu20iNY1oQmeYU6W9lcgG3bV0h
BZR6vEIZyUBK9NQmguf+t0u3Fbs5oUO8hInEsNEktx1pAV4TbZjVvKTgB3r2T78N
NTJbCZFGPDYXOeF760KamogCRZWHPvmWbcnlTXI5Kz1ZLBw9+kGikWfwxsFnd90I
Hk7b+i42rYYB3e6h7N8KNyKlilwye7+yz1QPU1/ONgDh7J51pRsnuqEmMfiQtV7H
vuMG2f5LFCcjwcKmEc569OUCasHtpMz2WLgA12KTuI6j0RH9AFN3/uwIK9/qvU33
ABBs4ZgbwkkhmsuiPLgtATWQVfrY3O8EejktlHLlHg629A0EeAoCo3G2NYOGNsAK
0VyHlWSigM1ZI8L43Pmki72kWuoQ2aQz3MoietGCI5NAhC3Cm+0MIbrNUOaGTQqS
Y8ozErbJ02NJCQD08rcSLk7RhVzxTPmS5EgVKZhjFmTZD7suAjaBUt4/onFIA5am
xF4RFLmOdBLUvBRF6YmUSHBaHzYtnvPzZhN9jrKwVvoqnk2k7lw2N/vDmJs1FYMR
S/+7P8+PObx3y6E3sRioDVfcquXqeyqVuUCuMzflQXijJqY+jpgPPqUFoShh3bvd
HD/EwDYqi1uYxGPEQHw7Tq4EcDSBUX2ZT+gMyUnAZjvlhGWhXdF9g6vJuaQK7AVm
rEIZsktY1Gx8kIdgYc/GF/Dh0tZ87dSBdpNHodgj+PDkUsiVZpRelcRPMPt+dxxQ
YT+CRe1PDsanmgIMC819u++ywRoA7jmjN3FgqtO1PLrvmXA/5IamzW/fzm5Bb0V4
GRjBXqB2fIzdhkXB04VgnmBMprOuIEtxa1vPuOLw+Q3xYbhGM6hQU4usqm0Z5HyY
/T1HWbvbiYGp4msf67hdET642in+fiY17TekPkMqeN4gcxOKFHA0qywPwT/ONopd
bsojqac8hhwTaeBbtlVN6tglXrX0nPUQFBhHvFloU0LJyzzULnZak8yNiZI2h5N8
ZBhyDi6MB6GJeMIH/wQO2/fyCekuaG8k77GXrmgPa90NQnzPqDahgNRTcXuslwgJ
G00BkmI9xlHx8pU5xq4IJ2WB1xq0ZqsjwqRJ8NWBPg1J5eOpLx/YCLAOGn+Nh0QL
BZCcca9S53ybDpXRqf1cgjXkob5NkqHU84G+EhbEa0g9ENtXYzNxh5vFhzbnTeB5
kcPIrS8G9oXJFK0ckLoNTanbGOVquHm1R/18k4tuhLDuRcZLXhsSQHKjVDS3iG6t
0rsIdqAJueHbePWZKOVt1sqMuu8tJOTK3o52aHMckAqCQ2jJfa7xFZcxTv4L+OXy
S4QYt1aqK2c7TAW2TB1ibKLKjUj9wPs5sonkiuoovm8LUhM1AVJzhJ5IaCxJockY
HmqjlMUr601tdeCShbWf1wMM7f4hlnGaQ1PQITO8NwvcbzH0w3w8H2BE+fbpTSoc
HG12kzs11P/z9PNqOj4iRy9dYdYSyN9qpNp3dlywhcXiEVz9deZTrlRQUHqzyYOT
Yj7dQQ2KQwX6ovMSv9oDKRIy0mRACRpq10jrD1AuyiMYN8cWIsPsx2NbjYOsuhwN
Lv4jnUy1HCvLjh5fLkeDBugCt6ThBYf82Ds7sWlRpR/aXXfdvFkloVRWK8Ux4Iqk
k6zSevJQtvF9l+Im2COrUP71SFZGqeaI+Pu3Ct2yGKjAImDNt8nYFBh2pcoDcd2x
wbh3Vontm5HK8Njew85eCZPyBbv7s1+L5ww95ppuEscyUjBMCA5zOY/4rOdtOQ4m
mhMgRNHpXSmJ9hRzNxQ5HDgQhEdiS5Fw8d4stSQCI4b3Bo5M25XugsCmYeedloyh
iBv4Ky0xg0pfqzp/YVXpshJbzst+7K5QVhTMlHhAc5AWKnl6LrHzp5RX4W9jeAyh
5482YJhOsYYde3+CsxbaGxlf7pI4cHKIK3+FUBUmO3xEzLN4Aronsmg/TgFUnPv0
1qSfk6TCg2vjdjB2JHg5wZ+ZRRjjutTBmaQc1iy4vGKpDXueeX+Y09vXqMIlUzpN
Ps8OXlt1ZR01Ng059IRDUpB1m8GGS3wdrehRTCJlEZExxtQxqVj2lhBY9CURQBDR
OuvJVbNJjxkh8y4WugI9OjTIJ+YPVPQCMYjGrwRXQOjNaHx+jLWPnEF7zvmQcTNl
E0pWKxR/quKL4Vgool0lJMVhhNWGiPyDt5/tOYUH8s5UdHBlB0fLiHt9Z5sxVKUt
Ss8F4ovvjwIKVfc+aeZDIncvQDeZ3Vwt2x0JTWM5/4ybI6VuEZ3swtyWs6rQSxxw
gN31JXBt7rf+DsThGvqTwVLvg1RNUiwJBoz/roCgPuPnTCmfjxbB3sGNUszRJ20K
U0jIzAtngwWQRvAWqtIgkVHXu18A0LJAaxbE/g2NxH0caWMmhvXrDlhzvuni1CfO
tfBYfUTJoU0i8qBSypSLDjdA0I2VQmfajd6NrWOek/JKjYYJkGWUXZIIIAEuEUo4
7NO4FzJhyzDwY1ys6iXREuP2FKW34e+ctdyl7YfQhN/aUZe/TX58SLzWLEwK/o5z
HpXPAhdoPue9FFujnSoKXnxcoF75FyXwgS1OFggF2chFTl22OvcmtYdA/HCeTDCj
9uoxEPXaBE7EuNm1RC2ZWukV0CqbxFs2LHFJiQ8sznokBBmgU3+bL/tZIntDDiLl
hGKipZ4EmUCaGeFqYrAJCRj6JavhViCxpZNtTPSiafqfINCuHrsnkH0/MEo1LnGv
A0uA6jw5hGelLkQz5F6UAk6LpQrzlnsGblSdauA0NgqwjoSKiQB1UuwQYm0ufUwd
dgizahgJUU6/gERCnUCgICplibDt+rhApDFH3mHlv5W6MNqRc9DN27xZT+kBokoA
KbtCRBtUXlvcEfv+lnTQRCkwKYwvMo6WVOvlrzh8d04V/AbONpzc7Es/4eKIcNLx
rlHUVdIcKFpfFsk498xzOpzn7TfyxcT/22loD85teF8DwuTeXOUzHpqidOpIXqpU
U34gYAZ8lonB8jXiBc+lwotD2JOlQkzQJXugXLsynva138H/IeYLvjNQgc8u3yPD
uFMIbyb2JAjrCb4Kl+mHp5jSkqxD4/qEeYIh85TsThmdler7F+zRNSCEVSDRns3C
+tCWoFybreO8qtks4Djwelwd+ApoSGXZqmgqhSz9crNzwiWKUJlSP+xSFWn3nhdt
kVldN8brPahy7pPT7bYMFF894nxCOp0aSSCwsdAr+Txqb9AuhU//pV4qZFIM887d
hic97Rzn3SZWAay1rbnjcuZRRlEOfvsTdk88V2YtU0luBcik3MqdJ8Qwt88pyWkX
kE8+rI32+WvzCrKKRzNBQa2omof4PM+RufruTrdZMUyvK5VKLpACtqtqX3iyYnea
T3mQPqo/cfFiU0QLv83qnm9akRxZWOnzP1MuOkumZf2/4ZGxE0o35dR7MWE7zCwA
NN4BS2hTZcUzXSLqhLn1uvfGXakov6FRCUSpHr1OpkoFhVC8v4xGGMvH0A3Ytr1Y
oYthapetaU2254/veyvLfR7O+aYAHoM+i+1Hs3Z7xrptQzQdEvVUbcDJC3CbYTwE
9vDHpN0dt+4PESybBTIGosKw6tjyY5LgBZmwGNCF9arGRnCRiVupNGeL5kITjyak
ABvwy3MqJny3X4y+DTe35oRP0pY+dzFDojiWpTC1TbluYG98rvYi7e5YwfAFbhVu
7lBF4fC77gVrE+5qAHE33mdkdKlaux1f8Z7K8Rm6hu/rqICUCHF5oAo8jgkLd1aI
o28sWkW8+P0BbFnjrGy6KaV/XLzXeFBl0kAIspLeaHoBZQU+OTrz2j7NSxSUY9WH
UcIBxywd99oYpCGFw+IHQLh7i+t1BISUkAfM+7ExvGSRRU7n8I2zLfctkoBIg2/m
bz6w5LQwFp6YfC2BypFsKzQclvD+BIpjYxE4SJ8jkxlKAZrgk4g9CfdqJhTbSsQB
S/fCs9ZW71VPN1+1cSva+eeR3w+eSDW7KSK7GQXuKDIN68YxwjTPc+nhwl3GjKOz
rVO8WZcEuyrYVrMHYbhkSZ+kE1IRiNdT1Xicx+8+QrY/NK/F2asmxMVSEM0KAjtJ
7oIbnc+hTtk0pP8nK4bjr1NGFSzHy2692OXb3d2UoeCsBEBAWl2AH3keXmVITPhA
8e7ftYWZVg+nMQXmdPsJdCnQeeLYkoGWgLfg6KEGweEYkYZQ2QwPgBE/myAIHDwp
gXDS7SQVCTZWKmdat2JEeJ9tAeZ9Mnq9qmRcBfIQTYTn+FsNo3W2iEpUC3zz/xjB
TV/Gx+EpAQWPe983zXiqjwrNzlaPh20AjA9BfOVFpDvD+WLAT5+3WvBynS0nNlX9
gmSWJR5O+s31nrpJmKQsnc+qRO5EsDpLsHW9kajw4cBj3Gs01ONa/uBRVdNUKvl0
Efa2WsVu/2MQtOWEYbgnjwrBCbqBdi4QIemTb0rwsRFXsP/2tpwHwqqehrapnf6a
s7/CE56OUfkNEhVnObZF/biH8aOskkovFFbUP3LnLvccpZ5MBft/aTvUz3USizXm
1ghW8y3jHQwPUKkz16XW4j3Gk9HEfmtcCwiDS5PFR/qNTryW06M3sHLK1+qA7lqn
2sAkaYi6VsCIZg9Fa1lcsR8GsFYS/Y69rnK2aCxrLmLfAUz6mcp0esU7/EGMQaDD
Nas+4FK5ZhBga+KsPqnCBas9iOmDZ00vFP/nObPu718cIHyo/NJxKlS3NZE/6elZ
jJ4VyVVwQb4ov3A6442HRZYlLxcr0RDHoea+4Ku9s3vJr8HS4c+HcdJmj/xHzIHh
lF1ebGQdanA+lzZs0YujP9unBAuFNDkct6DFH9pslOo2F7vBp7WIsyKZEN7BApiC
pZODnkE5fbQeiqHmwAIfdpv48qEUvwGKy5+yHCfRIfBefziZpa9o7NR0RRJe+ofv
msq62Zi3IjA6aOt7OoS5r/JDdphNuB9oYbIj7trSHPIzBBm6zCbHrgpkr7Cde7eR
Xx7nuEXNpRzrl1ryBOYkRKdS/barR2q/68tSYoD3UsLQ/nZs4SQeVDQt21ytmq2i
+KL52Tf7w6YDGZVqM8C9UCW4rzJG5ffV+WP3hNYYSyWMMI2H81MqmzM/hLsGWWI7
inp7HzjL84DrV/KbOZ0Egr3D4XXt/qTQ8pd2QEb398bq/b6Knq949ELYxOxshqPC
kJAbcTZPwZMFcEZ7qPvCLtuxWQcBgY3h8puXK5HZBpWPxwZMVyg08lc+Ekq18PvX
2yUMV+gK1jJxB6Nrp+4Q3eYG3HMp3Nty0YCvFZtRow64V9qjWCnadtQTuP1Ggifw
ct+PW143l+WKGof10E/FvuUZo/jHhvVket83Cu1O0Nc4effFBwEm3+kJz0vMsKgt
Xt+7jUaDwtm/Q5OQ7G6gRmDLUKrt+q7YuZQnw0hPOrn+CbJv5s0AxIORrrbgh1DZ
yOgFNJoosU1FYDsw/440XfAeqHs+5KTmfvVrVuZ8bFEl+ysElNHdxUvmBRN4F0OQ
mAOm4rTPFZOvKqRARudKtCBU7fSK/mN9j2lXLUFgfdeGAkL4nPFV0IG1FdBzweIO
BKrPt4eKN15NhR5Npw0pel5elGhE+7MmTnesu5BuAPRNAi5XhrbprMq+hzDPdlhR
ZyhieRvlsGqD3JFgNTON7h0sN9m6zDyDWDHquQUSfZtxIR8U7NXXXLQFNQS+oF0N
jUDosbLs4fj4c8U36qjALAr0Vg4tfHziREISltgNnN9syGikZUyporJp1B10egVu
vJkxckyXTra4CLy/0QjB002AOzkq80MUyGcRtCHf4iGOtlmiOyKtalFaLszmRLZp
qWswuAXdVrSLtuwDWyf8gNjGQD9CyW+wF5oFbL+WhXopuNqijOjrenQlFXfe2Py1
zBT8FQ4ujXhY4LPeQBVfNoNefeED/4kCut5GZWfmF+oSrtl02Pj4UudLaEUP6gUy
25koHz9lTFZStNvrXC3CDiFrqqJpGq9mWtYjynbuS7LpGbmS26BDzpF7Tq4nhiGZ
Tkt/NhXSmD9TkIczLFb+MYXMApVMlePWtsbRQwZl3JEgJbljwRgiOdPJc1oUVhO1
LZVzuvxb/OaZ/wtLc6SBSmcnE0S/yin26Lu7jOO4nYwTrNAgM/dir6zt/+ZhyXKY
KeTsYaCTvNXB3MVxXmKAS3MCk6w42FMXXUnnqhHSrD6UiR8Tko7llmP4AXZGgCpq
6/vkR3MeLwdQSgxAklawZpT9cdBSIV4lGhD7ZvoJa+OI0OLhuHLUeEQ5Aiyhh6+y
/GdQTRfTi6u5CDcQ3XaRJT0Xjm4H3gQ5oCZs049gtZxZj8tc4D8o7SQxW42+rE8A
yQhgk2/z0ncA2OkKWnoZegv/sw5/+FtAEPWf1OcDslXu94pX+ijOxlVxnwxVN6+8
IagZ6Bq0wEU16dzKtX1hwgUZSlFJnC4iVPT3xhZElAQp1ICVKQYGE5tUHlD6B6wj
oHmmSeYOFFUm6dAK3s0Bd8WZW6CC1ipZ5zTlIZz3S7MYOFdb1Urx/aohBvOe8nPr
n6kZo1PRwPN3fcEy784KnD7hSYdiQMbCo8HqVJY3043IcekXbkL4cTvYz1hxAO9v
/Nbfkign9u2UV1r7oTK0XA+Gy+h/+1sLp5c+u2T4LjcEncrVDu600TbXoDikJShL
zFz+gALicnMe3vwCxrRHkCQcLWdPR6F2eKF/zT65mf6BypV5oW3Pq3UvUfiHi7Iq
KFjV+Fsre8E65aBc37XrxJ9Ik6BoBYSl9famQ0FqweEHUroQsWeqsNNWhBd/SwLy
nW1e4+KAi3UTZkhT1Lq9L+3O7yuByJxPJXEq+ph5gy0D08eSKh3PutoMiOK9m0Fy
Q1gxlGF0H2H02EJdstTD7f4ea6Xnh0EZCDP8WU+eIExxJGIplQ/rtoWt84gPF95/
nR7y/YzyxlcnQTGZloYsbagmcKx3eagZk9WwIPTPYtyhYV6m98sMziLBEMNFAe/7
pD9+ZQ8VCk5Yjp8CWvvOkqxbSoT7AqbGI95bSosUu24Vb5k/EznAPXPFOe9xAxG0
SXGrnuqSu2G84kY+LG4hLmuHglq2XpF02IKRscxpZz+mlxUUBXDhUUUVqowG0iPi
ZrzXs+gXKOk2SZtQA5DQ6HRLixd3gBJ8Cx8e0bI37I0UZvd7t8GiDcsXUNjxmHgM
59iVXrwzY5WMSDJv1IfHjlstwecCguJOaMBejJNrhqBk6ri0LF/SInm5nYtYXEMN
h9+VjqwRwCGna43zFDOEeaoDabmxe1S0kx7V7qrD2ArHshLY6PY5Xt2uWLhczxtG
S5IvP97742nbviHuO8l+VfAYXJTLxmpj+N9J0GEfqGBQY3Tp79W70//SOHYNJSJI
Byu2RxiEx8BBzKKJIRqpB05Ar6R1GtUlOhsJykRMKlWfCVR3JPhG3A5iYOmxOQbT
2zIdlqMIHo0M6mhwkPk5xm8BRhPi29ZHqkNHX6wNdfyDRl4IFKX5Z2Ofuq6QiD97
0IE8DXSS8pJF9O9Ghk5aQ5v4w1A+kirHWuzcRGGJRrcusX5ltD046g2D08c4ER9M
rbvy6bB9oH0+tRJ0NbQqo5EVPYXnm3dvp0AGQ1oYtd9V+sWU+Xp/USzK4rb0ZZ29
YFQFCyMU8f7N3leXMJTWFrjvu7ZWSpfKe+bztBQ4ar58J2+jS2czmI4voFf3NrLT
qT/MjM3nBPsbYrq2EJFc+g==
`pragma protect end_protected
