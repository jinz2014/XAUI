// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hGYLGZds7pcIMskWvU4U6Dq+87OBiptz0U/DjsrIkeeb8Bj6Vr+VeSJ/vMULY/MG
0RC3papFY8yk0ax9FLcHJQI5uKTtt3RAs1VQdoEhLaE+sP2MlD+pvihkWM77fS0n
fVBwDr+HeMOLAbN1I4znluvPnaP6pl0b2lWiC8C0TE8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5920)
fpKNLxTW7RX7jDvHRU8L/UZc9nWZCJ+j/QaGXJhuGY33B5vFQWYQJihqoWXjK5/Z
CHxQq7ADxBylA0bEYZve4IiLBEjzuVnGS+k4JNL9cCsqoihO6mlBP3vkrJHRJpWF
tWJZZ7IWKjpF8KmvgnwZbxnCtDeazrzyL9tzsElk9eoLz4q1hZ62GqUPsO8d97F4
6aA2wQaQMy5U1SPWFNVQdbB+MGXfYE+JzUSoOE8OMd0nWGt6mYJQIs2IztJnHfYJ
L2ZLaZN49W2Qu48Vuc7T/EDt97yyCuG1mBzzw9zC8SSkMwbpeEla4QP/d+U6kzMm
7u/0WhTRmaUjhgBWBuwvuZuaAZLmHMvWuKj+M5K9tUE5/PUxR5tuVJWs5s/thYXM
/OTZ89fpoUwFEHEEGFWi//f8UjV/pjk8Mq1qAa0Sehe6NdOOKWTgW8HnJGqMTsqZ
Y5v/yTOusdhs84Jae4147b0n+8xKaE5OCp3zbsryZSm0o/A3s43O6SC29snXwrPo
jlEGBnxeocu/lWqW7OfxivWRSCgduEoYifmMHojHktAd0rfdMiqeQ2kVPyUno7hD
8zhOtvTyYdeAYSzWhd+KtzfJ7u1DbEN5Mj3aLX62k92bE1TcUbWUjIqgyaIplKyh
obYJsazTT7BNFzOvOg0XnrcbRzIOl5LVJGyMg99mAWc4MRseyqwnOYZ4vGIAmwB+
z+f9ZmlmL4X5mjaEyuDKj+UXRUmKyHXdlf1K8Er5Ohr3KQG13h43y5jDPon0A+GR
KcvPwFT3LlNCbMgyxPhLECLPas/e/8Xh8vsmf/u9xAzY4kJfxApfw05jbUkbrjEx
5PhgOhv6wijd80rdhyZrsF6aLLVxpaWQrnrD5WQrStRxn02mYU5LC501H+Vpr657
3lSFcsI9fFObfNFk7LGtClmFx/SR26GnwYpH06UHKBpnvQLrk72pB8/kI1k31bA7
GZwUwA8SOGpWw8rh/rqcCIpe1DTVn6cykgzv19/+qZhHnvzajpcCU3UhpNZyjcip
YdD9aKlNel170SCfNAU+BMzkCfyId+GMpOuKmaRTQTuBgIzrPzqP9O10xtBVeoD3
V7LXTz6W4RL1m4Hq7TiDV52/d0n4XYv8pVq9gT163miw3kz2wDskrRioCe0iaENH
auFc2hG5GOKW50VJJ/32x9/sim/WY1aO30DnSDDpbcyPDTgvBjkfmVK/adlHWcMr
d9mqSSCG7wM2JMcCxNn6uDfmTkErlRbs2NsFAlwEGfQwx1UrytejnKjh0aityOC8
Kb06FlkdjNwTGozqINRwG44gwJOpXCa1tbtbNijWfPNDz9f483He73xnCLRU19e2
7qTvPD7zg6VpWfCpP8OZlaXwcP3YQyzQspd4uC0DImSKMhaAVsNHL8tePYN7hU7Q
eUY6UOxVg4Ao4qUZtam1E2VHX81qLFBvVF7VMCmAILL+JivRJGeZg+IkU2gkbZVO
KzPvy01aCQyw+BsUbglgRBRrWCoSgZuSlVoR+e6PTz3m0EnejKNOZVDWwQURkdLr
vJJSWo7xkHtRZ1icbsdclh8/u5a/jTi3VfusBFJiBM9uYGH0WCU9yPguHsT2cor1
FJBbJjk61HvlZuRT4g/10bFo76d77klUnBZ0AUcBnGmTQHuFII1AxAMMta7TGqkW
uZ1OUmIkFoTP3QUWqXosamL1Cp0dl2eNQ34sg0KDrRGP3SzrQvRF2iychES144jZ
bwPa0EG+ZaZIFw7UXMX0s1aOqjWxTKc8H2MNYUNjglHN2iKP5VdeLKVNuALD2ev1
ly/yIKJWINgPUn8K7kpm1vJH/PSo5LpHgCqcmwk76S2uoO1BcoP4oLdhwuhVMDDI
DOuDYrL5YKC7Qdq8lepFUyGNSeyuHiE3XhB36QM3rg+3q0QFv0w9FaHIGPY8xDvy
McrnYzw8fIZmOKqxW33W5arLElCz1Swmg7LbSmO4TaD9ZRwh68H5S87VKdEaHzG0
tFNCWgvLc3u9SBxo/Qyv5BKIqaEi95M/LmH5rnpjsvlG7kzJsmwJ7mDFDJ9c9OeG
JhDPnaWws3MV1ABZ0gtJyVUufjOrLkJOsfcr/IGF1UA1ds6Dhi02NJL/4HR52mss
Y205xD/DBhz61vQmT5lVUGa4XItFDSKrWtdxUa/ddTkVOqqUpP0WEjMHctLzYohr
JtqLmlsX+HqbMlNDrHCQyBG/W7fjSdYrwROOvU+toMmiJa2NNuzoC7ln4eTUmYO5
MaeH6IUi3PM71JFLZBXiVwmXp2UZgddyvvfbaEWk1Nl89YUMrrF8aZXcEPXXXHYp
avH4P7vn0qQ7aLYt2NunNPGKQ84ti3drXo3jTlsq4VFBDbjjTrysm8AIokLBYZhJ
UoY3nrWBNPOJU3iZSe31mWVdSQU+o9Ln0XpFd5uB5cHcUJwsKt226Bg5HZG9WrcS
FAYaYoU/IB4CuED8Adc4Tb5AhnnBPcVH8Kdjw4/M4CALvzZlncUg1T83tbycTUEC
fFUrBJvgsvjy3wvn9HnyzlL5i+IPs2+MfaVb4bH3+lxdn/FR/HIHakYZgqn5wBcr
6SoKFIsSwDJkGOYjqZljpu7Tcn9dbQ6moSbF2vbkvooIYxb1NF6BcAExnUD70XxY
nrkbyiCPKaQf5DsX1nlWH8KpxS52s/FIQPxG9TBTA8CGGGzv7KW/aPANBACXD7O0
vUV4p8IE3zkWCMOoHvkRWOk7T6YHNzk/bqGDDbTbOnyaZzN0OlDDk4ZygPcIv/ET
mGCRpZbP72nPpbKWWoT6qyapGxzVzdEco5t9UVgCxra1eNZTLYM0UH6Kaikkczmd
MvUyd/O9Wjan6PL/5G/y9HvUbJzgJhwN3B63G7SalLN3QB+GzKvVrCKyRKrFHS2H
e0CNGxeekAqVzoKhS8G7JYg7qE3daFRJmhXLuCrVCQzRWgfcFCWTtNkwpLTrg9TF
qhFHqpRsbmwesKZzn2MFKur6bA4Rz7QuK22pd1n6WbkB4fSygNitW7FUrR3hJtP0
oTRHA14H3WXLhlxplZ2ZGSTuSVv1Y21VEzwgNJdmA19q7VHWYdpX8i6R9gHnkVFY
TH7QvLFez1MwstYZvFcnuMqke1bcFzm8+grSOZrHVJdhbSLzaTc05a69UzoN8+WQ
cHL9Mn+vXzEzLmnn+XT/pzpFLrzMTZ+1LEkt0gNwFCO6t/un73yKpQQqvvgiEdbB
ssf+CuNDHbBJuizqoHID0TrfjibY3gnpPPItB/cgQ9qv5ApUV4gUZtdKbVhZCUDk
aQLlWBtfbzxxukDZrhZKsgx3ERcGweMLfjVyvyUyKFgicrY0/u5bwids/AtaftiN
mlM7WVDgdnmCYP673nsFkTjZPG1kt3kjP+rbUs4ItsNb9YzfAnY59d8exDOwwUKH
k3/zMzH8OFjCG0Rn2lQq6XTSgIyjKjNxZsR4JYNIvbo5t6EQB6qxH0/uLmdTwJ2W
eg69gBeIDQ0P4XT8uDNPBsvWKhADRUc+aDSb7dKvF6IDv7Ohu73xIqRJxCGgU3n9
lkR+LQv7CC1ULdxNiUUQA2pvj2gOQAm5q7+kh6sTi6KobWsz9V0nbNbcKsL+d513
XJtXlnO9HgK5xZMTcDYgh/EoPazAiDoa2aiEoMoejYN3gIvGShKw2D030C4O5pFr
u2NFb3R2YHn37ymuwvLfvcyJzMgVWwl0isFnBfQo1xc2ztlIr/YljjRyPxGVpbDx
i3hjkE+4dflUObKlKwRDKcYO2EO17Ospjsk9zFxqPKRma780LOjuf2+IO1MpG31/
t1QmivR+YENo8phnWWumHWtDyiH+lzcQy8neIj7xUitGn27WHS/C23Gx6ozkzF0N
4bfPe030/EEA1uua3m1oKXjzRpOrPKxpuG4k3cromNUajiyVVA/Xi0UJylBkn/N5
JqPw6YAFNsAZdQurc1OE/6OSa9jLAYSo6h1IClkLqL1ToDXvqcPJ4jeEi4UeHDfU
vFALBOHgFyfrG4a6XCQX2SUAcUKp/ezqhi567me43FanyIwA53NaKmWolFvDCY49
KhoDsI5GggJQMrpDpAzmICJVMIWaIfYwROUpXoKDiC8570s2S4cAoUGK42m3JVp6
mWvB7ywF2aEwlyeoXDJscWc3Snz+OZsYkVrvcc0FP6CKCe4ilzk5tw8sp566bPcj
lPn2BAxEqOuaW2O/xgijoR8AgMgClz8LND2GklnLMUPYoLk9Hz5anjGojpYNlT/N
EFt8lDlfmcxpEHpL2vWIVOCOzkO6lALin+sEsfoTUNEJrC45J8GdbakAq+l7zAIO
nPyeviCDZlFEacgcsC3dJ260V+z3GSEcKbGyAUrTRwwy9XTNpBEaGc7LBpvWv4At
IgsMK60+WicOdWuiNTza1uZaB+tFQAwAzP02SojfrWNe+hhxrvFU+E1im/uqkNk/
6zVFcVs4btx9NSbop2qHUXZe2byt85mjibQyL+0sbWxOQKKzD6M330BoF1X6Y56M
mMRj7wiyf9aZxWewHt5cWwc2C11PfWaoU4PvSFBMst5vtD7DNsFDgYO6WX3J7irX
0IkRD8EBrHD+7GXlz3H0aoEDr1FkKIJZeyEJ5ss9XtspN4XVNT4VDLnGX1HOstyj
e7eKmVuki9YtvgOJeFOtFz87qE03iZmAvqgBej/cN/mUONeG9qYKOb9aUL7fPmQv
OV2xBzxLyqME3qi5300ToNwZTd3IPZirbDmo0wSbLXIap4f+n4PIxZrNKUGr26t7
tCv3eFsmkctL/O1+u6dqPr0bHhDgkEBvNYqB7NxcsbBAR4UQbcc03cCqH0jOD2C4
WkGcUeVid7kzygvLQXh9W3JSyJGnUwhZEVF0u2Bsm9fgGylnwJUTV5n2Y9mdPMKz
5CqmlT9dz5odeqp8tKV9BBnbUikRl6wloWqAwlkXXGPBVaneU2pvYWpOm82XTgCx
ilmegLVfeoistGwygMRdpiVrX06hD3vef5iTuX5/+uyDhkpfcdAOd9pusIWjQNNx
1sE7B/hxB/GXzd3hfth8blpM9USL9eNjmhpuoO7W8xfx4Lx4RWpbKrr9VVCeZjia
+LKjKxEdO4xz7/sf+yc/cUdnE3MXOLysHM0C8ikftke+oDZSgN0dWFkWX5Jr5rn8
AUuvllavrKyWZjtk6IdhdM2w+1HakLetJZMT3n2sPXABLAQ9huHeZix0tsT3IR40
tRx3ZdIhR3Qbxrx7Y9xFckBr9UUtj8EesYNwlIDWyE8dC+Rrv3uHsutzGjteDSml
UFG+yE4yCySkgV8xnKYvsYG1WNh7LQp5E2wVkhdvalHcfoxiNZvc89QOSclzNpDH
PqlqW8hH4DrVxyTu6OuRzaaU1X0HTwl0V62rPcPF34DZw19QOCALNphmfcZvtvlH
sb8w8gmdu5IITJL7kParUX6E0QpC6OGq/dhbIBsKYUGihrKT+H7URiMucfVodxkF
CNV/ZgghH1ZNFX1SsHMURU1G5GLs5z34epPDYLyujTRRpG7fAX6yu2p36clUjseh
OmAggrqD6I5hfeUhTVMUTQGbRI9q2RVqyEi0wNwEoJIWIhcRIXXP7xwHsmHqqPXN
VWUPhRi9vX4WokceNbEsDOXQ4Zw3e4R+mL/pFFtPpSG7UbDbp78JjKb9Dm9y0+4s
X1m0ULah3AcFwnfqvh+aYC/Uc7JQBlz42STB2PKgIZpOWlaYttWogK3aDqe16jqk
p4QwR/FirtVdrgi7/PFFPGlLRPXBkKjf2PCdgsbYm3lHz4m3U3K6idQ0XUS+A1Yu
vbzZdwuVdXDoGxPODFPcPbWtUerxgCDwq/5Hr7giKOFQXxGTxvtgGmdRASINml9x
YEZtuS01J13/VIAPn7wvOACB0YA74Y39DPsz3NuvIUcJJjDdqPMwzdOeoE5mjcY0
wl9y/GvALez5CCD6lMEv2bKMnF9aLFkEfT1VANOaw92lMKEqlhrUNSjnSQ27DtFJ
K/OtIFwvCk1Fjy/6V461jFn1Ni3GJXSGlBJTu2vqP50+welGftxg6snQcejQa5uM
cu7lqsEZONVuhzj2rZhX0e2y8D/f47yKedAQaPoWUwtmQaQrcmQXRtpK4MkaICOD
b9x2xiijgXnRLP/dpuIZzPFLVB0r/ESSn2/2ihT4cGTqHfENUJB5KgpqyEwgHD5U
wHPkxscUSCBWTEuoXaeFmzAx/W+OrCbyI2qu0TrgIZhNV/soHXVzczaE905WHaJS
gnmsHg0bkgGvCiPn72prpiCmZtC1zwUlUh69JNIYFp249yf6HvynDUUk0r1M10be
jrmJcQJjg0oiILsINeDjpeRBZUoBXmYEX+4u+EKvA5KMZa2HWpKpRSacl8VX59Id
z/W8lnR8VesNoNGVBzpXaaqVMUORD2JB/2fuuP1rT3iAOyglvZEfJrb3Bc6UOMO3
H2JlGTYx0Vm5O8m9vamXleKrvzBCowcl5XnQsu5fyazIKen+u0Qor9keCEK8Ossj
TrEkHW3Fvx+Cgngyg4xCUM/57cmxSyVYyGx4RoxSvpAwcg4zOe6UwDpmiDEPp7rE
0OwwXp22inphDDo1BZsDHZ4buwW7ktVnFZLnAblrfGL1ZxW0qzwOte8hy+AS2DIN
idOpHtbvswmQwcZIf6h2ZCS7dLug/3OmgiscN7O6f4apMdIeOlvGRxkhDKqMU50v
DZmyfPd1o32MZhgYIxpR0gcDge1z5Pjo8FAPXHoNBYoiKvDMzaxrKi9lRWSZ6Y/O
2Ag7NQyQYCn3Qqi316GAwCoI+/gUBt8ej6FfHMa8zIAL5iJIBuRKRgSxt1qPWGVg
c3nwR+nQTYWOFjxGXBwp3wPqf2StTUOipP6a3bzydQAs5AHPUWosbbQjzo3276H4
tOS1YeuHk2fX2yFLqF0ij745/IHcXkhFEkcj7h7DsrnZ9iorqkHIfPP1bD6octrc
lxV255oOkjS2Ek+hgp7Q5VT6LpjPANjm93773ZYSxIu4Snz//nTeopzOFCjwPo1f
OdtIJmpWDGh9UpI9XGa69tQ4WW0NbYR4WcX4QPMsJhnZoLHA9sptKizJtKRik6kW
y0v5WAV4gH3BpA4xsBbQtXIp6S+h8I0sVhm6wy/AJ7nC8Qt8Bp5KENgPrlFEovPO
q6dG+uMumOUVuu2ycD5o/zyILlRzHoPrCB5pwX/0VK5uApecF806tXBdlGO4kMkV
AFImA9Oy3zViL44CtBSLH9xTdKgYGpOW1BR/kZAgWD+lViMt8mBe6c7/7dmrWeEs
svluSii494waiKlQUvdmX1oEo3w8rGlj+54ZYAbno8AbOpKX1SIlpMBokhHr8fyb
foknACroeB0x2cKjlf66wMbLxVbpSBYvc1ucnz+M5EnChRCg9o7lFqm0GHEUqO0v
JQZfK2Cw5KXP6ff+22gfPZeB6F8S9WRV4UjGkxCRXD2CL6QCt/Sqkzxww3F8NK2l
mQi1m/lnjlBF7g+pNZjEzg5ICqjUv1ib+wWUHtIcMpmkbtfQFD8gzu13u/3hHGFi
smRo8teAkR87mwjlKpdTpxbc/EZAu7y380TDXX9DBRwzS00pxnsjg/CMCerhbTzC
ZuPi1PrJ625nXXJFdFhQDBsXtZ9VmDHIgFwa1pAQL9HL8PdnuiZmeUSElF6tZZUc
xx8EmSegsHltRlHUezg59COfrWol8b7ptOS7X5xR8LzWREczw8Gnv4rZKgbiE3n/
57P4omnQr0olH8pq/aCHC4dcKLw2tFSEr9lfMgfCMWiZT8UelwzJKxmOu8t7lm1C
GOAAK9OiOjE0oHdh1z57x1v8uT9UuCnyiAA5YEyi87m+KU6XweR1rJjY6Z3u7Pfo
unmEGzadaifyPqhDL4dMHvdZOxclUgQ5gcC6/JDYLZ2Pw146Cy4NLLHJj62rQulk
hjdOj55C1CVw6zPjL42lSA==
`pragma protect end_protected
