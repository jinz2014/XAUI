// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YnTG4xz9r3WE8lXI8h7vlMgnjUIbo4fABGArCp5wqLbq7B6I28O6Gk8uEYRd38Ai
0JxB1HoEV9T3e2MJEBcAap1pgvZLay5yHNFmJciz9RMQxRqad6HIuncf9OwGH8Ct
fpxYLdIsqXEJlMKImDx/mG8Uvub2W5ZeEj7TfY9x3V4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21936)
FgH/DfkvPtM3IhFPgaAfSQay5CWEp/OqoXzfFhJKPAoL5M1iaf/+hp+JgymiBeRM
pmMr/9csyCHDqxJGjmJ5mY0Aauz+cnq6oj65QZWvgfbLNNO+k0X1CcEHRWtjDeOn
G3Nia+8P2OBsese9/IxpyL+0jinwRJ0ZVEAKft5cLv3LUlKcauEkESpQvtpTi8tE
v9iX1dyC2F1Q1Ji8m236L/IRAoR9W+epoOivsurjLzMEAiSvsWkXFbxyl1oG7rfr
/sRRsp0buVuEM22wZAE6hqex+g/eOe8ys5PJ43C+UQibivlfLUoCV2gy6jn1l+IY
d5KX+ogZGPoGwI73npTRpnR58phBHOfYXG6CNb0JoaqlIMKJAzozgtCJhrcYZkoU
+5i/qwYcSvaMUd4TN6Q2DN6PaFLvYZqfe9BYVB0m710uNZtWj/favqw9P7dFg9y1
Od7jElQ7XCDKryrbTH5GpHztbfxZymT1GwT/FO2FywL7JoCJ1W4oLpOI52FsnzkW
iBInpBgIqkYoMdGAtIbtAJSyzPBQMKq1M43Lw4AO8P5rZPj7HdLl8N3yWv/VgYgc
9p7Zk1UpH9q9KRXhSbTL65VS14i3DNzshck7UQzXBFeK5ck0iiwxR7XFp2kGtI9p
GGOLrRZMCsUnnw9EGjZdVYHdseqShnEu2Fm8zCh1HEvqRdDhVyUMUKE9t7JiKMso
+3RMltCpjsDhppb33zhtFgd/c+l94o1JdCjymEEHyKUXmE3jY2SpVzc9bis9BBr9
jhYcA32pC3x6uwm3GSbm1r32Fk27D9XOHzR5DeT/XrxJ8WNFpBXcnWkrHYtu71/V
Uf+tirAGYR82WhFr+KPtVkoc6csBgErCHP8FSqU4ys4A11P9sbRn/gNqYxCXZEIn
Kt7Z85m6sCqNGPCmIUqONi5J6UkkbuHKt7syUyRPHcVtK6aosLWa1VXL9zb2CjMt
MkntLeFp5AeADSscMoHuTB45Ybe4uJxeiQD3htHv2+qXpmwzNBW2BtyKqbW8xQel
YQcvHDdvv1m0z6HuN9aN1ilalFMXaFL8OklJm6l1cAxoNbK4o0qE3UVELGDZITPU
j5kVRaw1zw0BKWIFr8QcJPR5ElDwfsLGeXB9Npzus37ktC257mjpOHU1mCnrcwZC
KhwjPfgW02wfzrZhQbtvh9Nf5zcbnlxqu0BeA0d8AXtCTwLgKaixRCAfJnBagJUA
2tSPpk8rpgdgTjKpXZk49ZAgT4flKHmqHTbtg8zk5r1isuVZwCiOB863lOiv46xV
g/4A3KfVtYiMZDZUcK4NNV4iA4/npkXWnip30cr1E0RKW3UK1CBsUxD7GD7+axbD
zXPHZl2OdU0lEf6oiiJsqsgmid5mtGw2RXevcKGgyWfFMejDXAYJ2FjVievjTRZT
wYAltuQXhgjTYFE43gHbp6YGgnbOQnu03ofuR0MLmOtABJz+dsh4fRm3tl2Q7/BJ
Zq7CeLhQD4lDfwaTGxaO4kZG7Ik6JbBZW+mO3EcKqYUF8HtQD8wtoYYp12eTp7OI
QN1P5CyTE4RyKAraTuIoTlz/ENskENPTZ5AC3Ci6/iSpuTzCPtyiwVinckkxzm1S
SbW+DJmUcBA6O72jhM6PBvhkWVs3Dk0NVIpOqK1e+wFanONyaFfYEDSjs4lmCrxT
bV8j3p9imvg0ggsLGPopgmBa5bGXpGQn1dtxsYSK24/gTP5dc9u28EHPpHuVz65A
JsFUZ8VXqEvFGG1SDbiyyJeaP6oNhl+1qBL9xuyG9kTRuFIEImP2YNy/hcydlKtg
jRAtkQtGWj9xo7Z0dRctJsYqivTCKzS+GZp0mPEures9AbIUOaxCnxaxFTk1qqqq
2lKkSqKYFiXR3XkdxqhuuhIa5Nwhxwjlup5iEib0PGQovm/gOg36Bv+e7SwS5Oa8
XaIMaderONuLrlf1AS2jK9zDQx0yY4GPCXmSD0Phu6THp6dEoKijHPaaUGjHFfbf
Q2eWARnMr2zl7FEp84PXEBhBdiYuUaHhgdOpQFSRpQuXpIGRc5LVMrOx4v1rCA5d
kBHeUov4NfAOs5EuZrfGEDLaGjrw7DntUq4/KFbRgyOwv9z91Xi6Rmlq1kbwqnYe
eUsrycNuIjcoX70V3KB2fthRksjcKk5AUXa0w/w3S3+oFjtepwQAfK+5ErLTBI/3
jy/CFP3ztT14AkvTsotlg13lkS/EfNW6Gz+YHJjexzQuTYtcNVcXS6QpZyfJQnYf
ghdv8fhVbl/6g2SCbTMZjyzVxRLrf5tVOtkwmX4hsobnY6dryXziiHN9wNYY/UcQ
rABS0uCa+/nSCjMfeIIxi2kq9Si25vruclMm9kjCU0SDUHkmwrnm8oF5aYXu8YrX
LoaTcHJ0mIsgYMRKPe5lNT7L+l34yiZAsg7kmHLd7PBqbQSMaWU9WcH1p0+bfOkI
/I2vZgA7LiupLa7cOmBFoO1k1TuL9TGQ71I1UDFj1wxhDSMxa7RUy70pGFyHznKM
U9mD1NgUEpcYaCg5fjeedRRnvYOe0DYN6FCKJE/0Ac4OZDpfsbpcd7FV8cp8iJw8
2g7vKdMCYPHTbJEXBmKcR9Fui9c9/U/XHjDdDzrECs7eZWSNDifBWK0UHBVrwotg
EIffHOEX/naIEeFKfowKL8wA5N6vAn5+DTq77k6rW8xGtmJhuWoxyPXzYLMJWSfL
K+DkxsMTojkInIyM0hRndGvlw9+Dbw4fnysMeUPgO0tnQmJ/Nwtdk1JCuZ97chTU
eTUfUZQifXg0YUMRE42h4ECSoayDmHSRTHqRHipzFLs5mpg3zKogzG59oFgvMIkX
vIF8BO7cEhYqYPBtJGRGtyoW7d84m+J2fckt8Z88PExj8JPRVnSLpwuaYFxr2Qxw
4OrIdfR/E2DYezqyT08f8eMjZhuCl1mF89vjFqiZHuAP6TXQSoVtwRRiP/iJlnBq
wolKmWf6U5Y7IABeT2bOKw4iy9Xt6yEhz2kaRHaQlU0BhQMoP6TrrPqRk3UWpGul
X0Wsei7UAZoFwOuY2RyYdBFYQZuk6zv9fhTtxcwGnTYRK0/8MnjIXBbCmLw0eerN
d+xX/8/DEWXAhGMM0VO6XJLM3BRIrxc9oekVZf0ltq7qinLNyj5VghtIElzLnZTS
l0Z5dfCQbfSRSmEU+3mNel2OZ3iBpP93wJ9DMjKBkVSmdo02kexuGlzeV7fVTswW
7Iv09G6b4pDww9rbdEsOuCkqFRlY4p4u/5IdsX8c5ygR9kucEIW5CuyZ60E7V+ot
RkYSHX27Hx9NyrfHOaHujO+V+DIng6MYfprXFtlzZaa0eWGVSnj5kvKMiPRYJqqV
UkqRy1aWBL9v2TclZrVK5YrpPoh6SxOMnt3UoBKxmMltd0oQjarIrTydlE3yVzyi
OQPHB/hb69aaU9dkjKxi2hYcH+jgW2rf80py/mZ7WUVRKMjHP6k8mvr7hYpsUGG5
IfRm3sAIKsMZGPOnTfNop1cdXeg2jpTmCdtD5QkfNK0P04kvZ30sQPFjcK4/B7qF
+74wPXA1XRSWEKW7YgXc9DaxTQBOqenoRydGWbx8FZU4KMrUdR7tIq5xrgxkytub
Bc/mkDzX7x0XFjSzc/4mDt68cZvOf12Xsr4Qd8C90QCw8KK73ZylqKpKqDARF8x+
B0i/iZrI0dqfmFKL9Lvl4+NjinYj3P7CXmKNPlFUrLzfbrYAZyoYFicRyd5B0ldJ
r9X9Y8YFME8+nMYMxt9SqGXhmSitImJA7z8ryPqR8h5dnKfkrpSKs/PMXvaTOnJO
N3ch9N/ZvZMHXZgYUrf24RvdUoqoTzvU0Dn6OyWZZA2UB4IAD2Rml7w+NHwxBjUu
yyVrk1cdsQ4wMO4KmN44vyCJi6tqC6HO7pVXCZ/XBUdJZSSzzD1HKsxIkruDZ80s
wTaJf7SDv2HyYAkUD4eihdNNqRdEUeWNAFH/wQVFp735+Ko+5b+fSrP5QnJCSS0g
tSxnvP53oYOViHwBBgTXQKsZgTWfiv7EGgNs8w24GHdlpxiDYOMn5pj2TEUBYoa/
kFVVX1hAF0pM5/1Xs8IWaCxqCNrU69jwM5HLoscG4TGb+5v4t7CXIeCDSc08URta
DvEK/F92QpvJtt6VtTmd9JrN4lYVuMbljDOciAXJSG6SeDYjXWRN8ks1nYi1qbFP
F8IVZaKKc95Gu3mSkr3AN93iPUndoPrOavmCe9us0klDePSgPGEITAAhWGYdGV11
2A0dYKucSjbM70wtXCfaxn9VZMMRrgnIpotXF9WvWgPJAR1Rq5Sp5tAEeoNYqCJe
sXrGPYW9+ZVEZxDSk8xBebgVqdytKh2WJXNGnfNsEpD0p3NB4goEV0m/vEcovKWn
AXnFExcOx9M2y4lu0/ThqEFbiZfqjBl0DtfyDJmxEvC6xXq6tiKaBSaTz9CBIVZr
0ExJLk0F5BJ7BrB8BeBoYP3h/R+0GipO5Ylml26iAJlLCE6W/avWvYu1l0xXgqvR
xfBAmizLTt5eaXJDOJsESm9Aei1QaXGlY2KYBHAG2HJL2TSwMHeErwsCoXQxFaNL
Y7uUZ9teeSomuPz0YIiRESsePgCvADZBy2k1z3boXUMVW+WWN5ITWEY/mpwzdxSs
2dzsx5YpJnyMlZfdPN74LEF3S94xZijwa0lYLY1kMbTi0/t/l6coRNgz5jo9TP8m
BhGq834A3FDWdsazXqm83UDt02TDCEzSzZar9+eQBIaL4dRUEMmDefBfbCwtNrzw
0yoZv9hKnlgGqRmmnm5xPHEtTIOFCEFB/iRoZ2mMqAAJk4+D5yd2stdAQOqg6Sdj
jZwIWCuQp0EW0VwlhDJ6Mrw6CRcgUkwFr+oOOg7JInsiS8kW3O5hpWUNb4jEV9EM
RjqzdGT+Qb1hC1trkaAFkJIqzPBITW44oV8p2DWzAB9rWtl5srkIRDUtRR0/1C45
Xwcjm42VzrZLq/LIO2eatNfWknmD/fLVwntiIInk6eYpc8RcB3piGkmkFky1DkDC
NAIh6S3ipPU0Df5T3pokhENFLRUIvY8Bqiy9IhSOUsbMWhII2DOY9dlzzzdrbl5y
civaAPl6Qpw5+nHR/DgDl7KHU1/Cs14zTCPHdiIKQFK8lPMtHT96yP9pCn32a8A5
SNFwrJyvLCgOsDIB16yO2cQL8o+KI/NQYfxEmOzOuDb76F63xvg1f2ljr/8k1NXZ
0U8ss96v/Hc8cnmHAgn6cB0pMT3Eli8CprCpyfxz7HIRjOo3fxO1ggckzNskgeJ2
vD+9MwmH1wL4w/uKj/e1/UgAN4XbWkVquH2xUYkTV0lY7dnWnXczXqMiAlzoiYwF
SiZ0I10/WV3S9yasl/8SRFzbcRRacKli41tIBmP+hakBimhJdCPKwGqNlSUF5Nja
l555EbqIfRzDj7RZZB2K5ZMaxL3J1ZuzQdmv40J6bLspN9gX1E8KqYZfdSE9gGFZ
isWeMAmi3+nBqTSEfHDwH2xnkd1S4aorR0F5FPah6BEO/h7Sxv857+x+OEgHF/yl
r8bPtP+0jRUBolSwgxn4udB97aqZXPYNdJ9LmjJAJ4wEtedX9T5VVDiHYiAouLru
vBnL3CXlhKDLcUGoe20daBj8tsR7aL00Xz8CAmof/n11p/sCDpcRbARePFEiBZvX
Dw8tNwi8NmE887i15rwBsPu6bux9ehiZ0BXeoZrxcnFcjygtrxVCACnZR107blA6
N0mhBaBABlLeUeQuCTT0L9gDrbIkRUWZ82jMtURRQ3RXuTexjlf4FOKcS3EsZ6tD
SDiT76kDsOYNxNiKvk5E3X9o9yK5VwZdnEmw/zLKcPU2De1ap3Qu8Q1npoDATtFh
J1slFdjRZD5lDJHjmTq6ebE6r2AEOlBMxF66Kp90SP3KoDkACeg0A2gjKluVAoFc
fWZRmkuRhhlKLikGlNSbUn6iNph643i9/hVDx+qMvt6w/r2ksb2NKIUUpRVi+6JF
PmcjPc3fwo0okBWS0YAboIrOwl79HBR5JnuBTXsORp8AxVVP3eVOmDU8dH43NOWX
04RBeJfqokNkHd8hjdEXtON0vmSQmrY0ct/t6Qxh5jIfCMbrmsph5R6TojAZnbcO
2oVVRHsU2y9m1WYPivtZCZlrJDAwLwUy/YRSYqxnjAVzcIY1FYrzxgqFbquO3u+x
I81DBLUdNGMYkDmem5v7RTM8sPbBwJB26mXHKVDxFDOgfn5msQnfkfxvFeFlfEIg
/6jLCW1FPnnvR3ls2NSuaF3In3A+8PhSYJx4MVlIjuQKuhupFm5d2WShm1lwRmKp
YP6iSpwjC88PAN6doh/1VbTgfB+AnaKEW1IvGPTmPhEvpEAqwTtDayTKgeW95UV9
yi0i5/xyQiSzSY/z/N9+hMM+Og2fGGVZLLsgSl/+18Ji3FXBpN90W+21OuOJs5dV
tIZRAZmjjAF9uL1FAAmFym/LnvjHQXOXLgvDkulvuQDvWmzAICWpcyR4h+1DX236
Sji6I323tjboLo2LC6FTjvP0ZzbxnEHy8ssH51xIV5vqeMN/7XLwCOhit+759/AV
kmgNDCX7zKe+eXn4j6LL/2Zd97wscuF6kYit3kc7Npn9VoC9rfPD4wwrGGSIkDDI
ctSv59KMsvEzdKMLZH6iifauw+zRbYdF0XAKmkprcnPAqxlnhqjD7nhctKaurCcW
osZ96HEZWZfjOCpnUSq8sovuzxtFm90sx1z89h80/shLwHfzasAxQwNLs2dbngi+
zP75JfUyPmxpY1FoATvx1EvmUdJ9YpU/iMV4jJLPQDFZ4eiNVK0ixt1yagPBAtVJ
RGLThTYVwVjDwMM7/UQKtAWM2Ojb8oPSfBkP++L1dHEOtVyGEYQXzrIwVWOffij6
I9tHjmmDIjpTZJpRnqWWU4/QTO/j5g1d6bCaPq5GtBZ6YyVZVXiJUCCBkxsme7pF
m4w6rnTQywJ+gitxkvbt/Xe0BZ3QQ/U6YqQJDh6nd0VUfta0VosIMyeGaTsLgndN
YbHYV4g+k7s32X5wZJKyu/eDi95Ak3Gf58G/ucjjvXP0Wt8pc9uXeijyHPMpKvsT
TSgrZjGnvAKBVWax9tjNtpZikT9stemkjehjGS0YqiNHVcrDTXPxskE3nnoDwfJt
XeG43RjJ17jpGAGcrbqJUAyHBK6LXS9q2pFvGM8qXY5S1qFiyeZF0SXaPkgQA+0H
bYy2+MEjqKCpTvUM7l58/0D6WpdgXKh2IVlVicR2/QYRA8C/D0QzqKxDJQq1aTGH
5Oxn3Xl8BK+jAQCRPvXelNG+DNtF4FVLrVA8+cYHf0nxIhyG1MCGC3u4rtNok55C
WtnEAr0popmDeK3NMcpt9AVltjkBF0pHiU9cvDPEkHE+58sI8RQO4BpWwobIYj6j
ZRt3d9PlHcLRYMYtwA1RZkjhB/UeMDf81HuiinA//BoBK7awPbj708Gi/xKOMGJr
/r9woYdnvGKPhymAPuIqqZKJ17WJMPSxRqt54Ir11v2HhpMincYTLIoNOZEA6Eft
r3I90AnZl+dNcid+FI3Z8YQSo5pTYQe5/vQXaD34czrfHlmIeE43nDMOpqYRG/GJ
P0v5AgfvxZmpRAre8IIalHGK7+G46gbL76b3ESwTsPhV3E0AjretAwmGKYXhNi3y
4BwfsBglntYlmScD26/doIVhuYRQa0O4hERZv2/2cADwgMR/Tt5QqxspA/IhG1Ze
30d+rXFLHC/WoF/2HR0yR7thXIxRxGa/Ch8XFKoSLfLyJhqYSSLPRtti6alr7g9J
9TL6ei1bqv114vLH3VsHDeYaDilszNYvjR9HOImlu3sVay7gK0C90HFZJ2HkGWFJ
eagFCMPIBTq7s9EPHjx/CHlO6BcoLSzo+mpdFUn2t9zTeGZPHONYm/F2v+LuUwBK
g33fLujb/FMO3edTOtdeocQgouxwfyFb2NXGr9C3JzxWsxKW7LsiGo6wiWCByyDE
eBfF2F3aQhYpnP8qmOdhP5/UH6EVHiCbyCnVQi3/1PzpR+YHMGU0nf5PoY+QfZk1
Dvi8UvRp4tPbS+hbKrvlQ63OUXENOxrPCjzQMB81zU7z1Av0zl6f1ojGh+wuIcwD
IuBpBh2eJTCuyI13U1dv73Gl0UMoh5dfesFyE2UU0QbdZcXjincFfnKhVgTvEAg4
rsJ9eP2d7evCfznU6RxJ4X/Msw081YzGSlpmfiTe6f4SJtXI3P99Y6UP0QjSqdJF
UlH+Xq7jeqv0hC9JZj6BQr7Plc07Cz1th+bVNBxd6Hu0GxoG4/7dP9BsLknikHQ/
3ykjkne68Mg3eEaufE+/IBfBLay1Py6FlL/nwhbSvgflHpBBcYhLz+tbsws8SWgX
D48HJuNm2iEThokFyvJ3tPnZY4u8nhsz9btUBbV9UfB6KfGwYcnxRhp0ik7ybUtw
xoQ+nthCSHXlTHRPPMCTkAdF2aNIOTbCLOuQa9s5/Q/bqp2tzNwHRvieRusoX+PT
W4GG8Y8V6PBpAOtne7NtjmdET3axPFyAvLj8HcuQADrOr3/zjZd6OHTPODnqHGhP
w4vueq3QdTcK34bGV+ilSM8tvJfInpGrfiFZBg3px21N2J7LTo1nrLostc6FD2W5
w0lilNvOBV215GODs6VjBbscUO/rpnr6bMEFkeFzb/v18jmzZzX+pSrAouRtoHJ+
Wgv47UtrM6DrHeLwJX7OJmSNT+ZdO7Mnmx7FfH62gEoOTp+O/tuDgbLfuAtzHX7S
GbdUtpijf5s9xHGN5VbdgojI45KrrfbL6Dul+IcKZRsmG5cIG4BhpBe9hEl9B0+I
e4/UqOHMWX5UH72s2pvODZ8ErhtoN+VtQqJnG+nNmOC0YTpLEktE8Cqt4XdrYc8n
gCwo7ODUMHryM0o2GG1872HcJNRtiMp6zrSmOJEYA/g8VYJxT5wCxL8fyO2/auGl
YqpQAdBkcvzuMOBaGwBUo6jesnIUu0+ZdnHOJ04p2kjOhR5w20Twdr2QQ/GU885g
ZJrq1KIXFNYy58nRcYb3VqFCYQXXdLGRTe5bUsERi8/DE3ZPLmhluwQaRISW07zO
Vu8bXTpQVdCK3OEyYaLVTeprGKhZNGBHMMPV86TPWjcVrQJDr2pN0bEjsCOfAuNo
pltR7zfKR8AhAVZMj0BQvQcqX2dRU9QzeMlaEzaI49xEBUHnC6H5e80Uh1MLrZc7
KFHUpkZ3VXLkjrOt+mBmnly8dmhr3GmO7Zd5OgkKrl4DYJgKCONNnvNMYsYmNN3r
elVJ+qnNZ23DH9BoJyX0J/IFWU2e4KP5LxZueiQBGlWB28VRH98cZB5MgeHwLf5y
AV7bkBfRIg8xm+rnTcwDEFPL/mVHYeiDzzL4PPvpbFtWLVQ4J8J4JMjo/hvhWgt8
5b2xkDTJz87kmj3PJy4+0nVpTTn9v2DqX7Yulp9SkfWBhvATpa2Jn3qqjKUXQTAm
JyghVupEgQwSjc5O+KbRWQ2Sf4gPWTelHDiEtOQnq0Rh4FwsmfC2L1e8Dvs78xD1
AF0ApOwPK8ar4gUifg7YcmZk1N/dbSaOLgSGY7CnnxaePxVp9g1YK/jOKOiEYOMa
hPUprs8qOAJkxhjVtNGMjhW9+D/dNSayHODutdhQh0RuttzYIBVGUYp6z7Pqnzkw
sm5IZAAb+Lu77ZYyd0BV1LgRUUnI5Azonn1BPPSTCKvpkzZ5qE18NN+dHnEx3IgI
eqmnMObhjQBZN+FODlQL6kDxSMY1fuyIzEFdoqetHzqineh74OmTBQLvm3qc/xDX
cGEYpPKCqZLkQWi7v99WDQBt3bPPf9s2jOSdccpektvBziL5kZb6sbqmeD5JBCok
QwMZWVnA6PF4z0MIy6ivG6LxIjGQQm2jdgy5OGhrkoKs3BpLgZ3OAkvzJLd6NQbT
XQoN7pBpKnH+KuuuSJOPrbF3vBleswvNVQCKDH2SSoXvwLfIalSEK3sB1SCbbv2u
OOffRoF0vcx4z1xUp7j2hNBtw2cy4zbQKEVGoAfP8uULJlgV/KMs1JndAnd6wTTQ
876JVjLgfeXfOiypC0EHFWibq9AjTmOzi4OZiJeaQBTEgWuCFgvtnxkiwvqND+E2
Y5umnUU0wS1e4pr3rGf/bNg0nnImVnJbwY1eiSnWv/nQpn2LdVW4lmQHpfIlIBaN
PCXQ4H6qalMKx3l2HPnyOzVsPRovKhSCHjdMdJykHtialUTelGFLwjaix2VjCm+W
2inZzSa+Gr8G3/wg/n/ntoYmsuJjcKqUJtHr1t+L0n0BswX10oH0MD7nxEfQKmL+
xGGvyZx5jACQ/x78tE0BG3j48UeLNuEhPhEaTXCsMUs/moO1YOyxqqNbcC2dNKxP
9T+F9GgYdubNvVEIovUNaVnrbz3c444YqVwC002udsb3MACaZA6WC1GDaMd4djUl
yf17gsCAPl/PMOs04h8Yz1HzBzym+dPASjiqKOFiVnZuVwIA2gUMSFLrC/Wop/cc
0UfwE5Opmux2vop70dEK3NYGnVBgr4uDMd106D82f2gNSgm3mEsNNOE49AXvmmc+
KHT1NPbUOMuuwMS3h8TvZKgvE5Cn9CnynJv3n1qKibpiT/CxlhWY/ygNJ7U7vWT8
NGFGN+2De5wprnpfC6EAe4o9Wh9NcF4SdthoFLtwO5cbUzDGaDhkPR1bmeUr5YZ4
9KxVO2KfPI08HfqCF20MHQb3hu4LL/19vD023ZHhsHqtk9amK9JSpuWxm0/zlNIf
8UUpbqhp5sCwCNsoEVNqbKBIYcfXzdT3xq0OScri9nXG34sghwndbQXybqC9hEis
1o5mp2SGGKzEzVg5xYoYY/uN2lFWS7k/Z3oOLgYG5KyA/2JBuCoJSWyzXki6z4Ud
mXVGj31mfWxInUMAkvsdZR4KK5ISJlwM6+yLRPZqQuthif0SnYIiRPs66aEQ7VAk
V3hM4ncvoF2An0Wh1EYkZkSbCyWDktX+tqAnjGK291RNeTM4/RYV5xGjz1lmzt2z
dMUrbb/UxtP4MqaTp5MNpq7vTivEVbH21y7yP4tqrH+cyzNgAD1XYbnPMEX8ryAp
LQGii22Ys/w2zyHV6MqbuSNMPnvjNy7UZuKkevmfhR9UY360xOsFT/tvICHJMI+e
up51ZSoOSYbk2DVyoQ7KJQk3JcE0hDdCuqKkSkQGVIJ5Dw7ljzc8t1gNkLhJj1PN
V7O84LzcUba9Nm6wM30cXSq6fEVWppeyec1E7mJelM004W97KTg7CNKDX6EqLV2U
tz5QQB4i3zE0QchHKQ9vdm2QqJXHvU7fX6y4rcMy0dN+LXXO09qa5sNRFD0Ahpor
HyqJXikwEVnKFztfLS8EGU9eV2s8GxxeVUzKtWyTwxFbMaMisQB2eT52WR0gyiPL
jjpPH0ZynmGQyRzyo0dX7xD1Xxq85Q/jafaqe6kundJchNy6ouMpLZiDC1sZ3Yf3
9l4XT5Oxbn3RLtQkKCAFzj4nJ6DEZLR3QEwN21osuINvn/5gst6pYKE0ueN5snAu
RP/EoXbIYDc3iblCIejtYsdXqwHKes955sY3a6wMlJzbx7HD/PsYcBjx0QAnXFGq
BC8imQeOO/eKZCbLUqvn6ewQYr5JLkxb4HoJXkJx/9tmlzrHsD26W7q9eb7ntSH0
OW2KQITh8qCoDkIGUxEbDywOuGRnOJo1n7SAL2ooSxm0MMqzy5FjprDTdLtuxjLP
XPbpFsWyXw2LiXlp6r2OiYkYLEo3qdo2P9jVKDOPpY3ffPUeRRH6qe/3UIB7XPMk
gH5reTbAD7dL9fNgKf1U2WJtnvY9r9XJh99cZ1d9b1tBPrGAuETOHa6XnCGFE9Ie
ukULUHnkLkxDdD4ThXidTh8meWeZW867aW4xu2QQkXHCavgTteW6r4rrpZY2oWJk
sdAb3xm6V0/RsXdvf/rT+HTL1z7pnnTn4SzN0PFdl8TY1Jzv7PuhGdFki2wkzMAj
iaSDqBgaGZ7KPKWYg2I/iMFmwqVwDOocsODodzk3JPcX9e90394YyjID7RGKcXK2
O8N9H+p8uQVQ54S4RTBdhHcIyrp6kRMHlcxN3cjCgg2FU4wATU5Z2AVOxrxn5Hqv
VDo2bsPEd6qz85/ABK381SkI/tVqCqhiLAHEoMQxY0BFjwLkNgL4O4WERu9qsLat
7FOPOUBgMnlpOIwA9G3bNoZbwJi6Y38FzcmbtLQ+f7VKfeVBOWq8+DeDSH/g+cM6
YjHtIdxoV0AD9+ove+nwKUkk4ag+ALk344Xj5eThO1X84W1O8hV+jvnq/P1ifsdx
CrBaYU6eRU9FpzwDx1UW6Oed8iNRsk1fl5M9PMA/lfzegecJTlLgAwrolCcAyNiG
RWe3oQ71PwqYQ3g2M+4x4Cy4YhuI2ZoLz/+BblHeGV5AwJbJLOF5n+6td/6SrBxQ
J0gIdmRUDHO9d6Zex/dYrBrdv1TlTF1a/9t8FQaYdazo8nsvnRpE0K8cVQ020uIe
yxnZnLYdAXMS8b0QBpQZVb3tEOMJuY1U8Tvh6dOkdu2eLOaxIAKTdOwVv45++KJt
/i9SUU/iNV2urUbwnt77cGUSzOohrfWHLp/ST3lLmLxsuOHjLtiowtL2sYsmBlSj
OMUIMvOTd/AYhMYODxymZGQ7ooip+lVz7oQjkI0tLxNf+FrUv7n0e2rnvnVQpgVn
gTF+B6KUrBlXw+g0so9swoKVAwY+vGEt+x408tl8sNsjgAqpl5Yhjcjitj4eJ5Gm
hYi1560NVrIFCnaU1+kw0edb1lqDHvL+8T+Tb9XgvewKlATzDvAxYsaNHl0q8zXd
BgINCi4NKlpfAY/XKTpcEoeNkipMxm0QJ3CV0cQdZQ0I3bEiOJ1hHpwsB3LgNKht
etRRCn3iqXEcZ8x8jSUI4p3Rjger4ZLW+gsmmwbxPTY6olnW7kBGL5iEtJn6RAI4
+gEi8TbSoTXzBc0DjKsQ4SSE3U4YF3vjfEVEWxQeocBikb9SzaV2EcC+76derCsi
dUrPVALl0+6/HKCEQ5nKKOkJGO4Pn+8DXsWJC+KFDpIAzhsBoMq/Z5Ig9V5zQnFN
VDG2S0w8ehgODAlLu5ScThR0oX8QjXsXXN3QaekoA6Zu1PtbsbM3cgy8WdQ+Eavp
txGLjc3/DOoRqheqFIxYYmUQvdFUplh5xIhZfmlZZxoeyGLdM1MlejJ53yVhY9cZ
xfEu3ktkHrl9oqzTNUbTGC3ZaW0Yl9tleOeB6gvO2H6khCNrqIhGuLPsYm6P6mfB
Ic1tfQPFl087OxepkK7tcDMCMUxqZUzVCmsa8GRXXhG7YeEgRyEV8oQGe1hlTjxq
W6wvYQdaWr49IivhAWQeb0IxyE0jWgDN7pd22XmU1YFyIjc4iPatyL8B+RbSviC+
4MyBTg8FilVfBBAeXVvwECScgZumtVatT0MCg9Fl4EEMFKGM/nEwceX8Xy3Ixj5D
ird4iYTDt7K3QRjvZko6I4oWGNvmtayGdXfFDkB76g6VRQH3XQUIv+gxAUlbWZl3
nsxb6Z1c41DuRwvKv4VB9nTROb0p5Bful/E5MgemAa1x8POBuGFRo72h4hKU9yPz
2rDLKfcOTt66s0L/Wns925HUrjc4aQmMIOwyZfE9f/VAxBTSkSQmXxFeblvJJNOW
Ty85G7UOOW4q9dkMJU6hYikoT5I7ngiOWnAn5hkPPr8n7DoKZgmmyKSrH7IaqnJK
UMXxSv5McThHHSi7P/fUYkxyS3/7AtAQ8YOkyHDb02hDaQkBCNBC51DZZYjp7iAT
RIwLgycoJ2YuWa2ixgEifElcBPaSt4+R4H0oCD/kPFeZWEE+gXf0JDuJoQ8N2A/w
a7t9umnyfCBacgHfITtrTCxCQ8o06ZczREqnwitM8FSCSw0YqeyMCOUjDA3n8hUe
YoCBhpnmK3i8HJ4MDJYYjHWOJrdRIswKsCd0Q5Xi415LaZ3QZrvUql0y/zHvnc5M
v7D58rqcZUb7c3o7OCx3j+BeapJAK9laxCTblUm4i8JvSXFJAdRP9tB2oVAMXasT
cVAahIqV19FSfTxBNb5VVDJdgVhTBipmnkTmbcctZ2HrDenWhMLNB8hPYWhugVtm
i0pPAW4a9cid++jsXQbJ8v3yaocdPPoQ+NqoOA57YWO5HIREhPE1t3aLH3jYHQxq
flYVneZwdFlPuOLD7AXtphMAsAq8nqfT11hGxaRT5TmXiIjVCBEdMXwM/7JP+yoS
kbn+DHaWpyU2QWy57PYynx6nBar9kPqHCHQw0LL/2dU3XvpAlE8Lz8WyT8XSKOHm
tmUYuXF3zNb5BB5ifNW0/sk/41+5zFBQHyIesWLrLlA/xL5GbxVjvgKjDTWODw+p
0Zc9I5RjomD5fnyYNmO+k0LY3GSH/hYs4AirOlao/+MgNEstsel8Bz8sHfOjCTnF
miZVP45+WnFyUE5VwXhyO5Fzc7gFTVVqJsN4g3rIhGMSLYPCscIYfSfe/AWxLb9c
kzEyz/LEBpT+Pu7Yhqnahay3fzTmDQjCwAKc4CaN0pHL3I1wMsumzFB9bUWK3M4q
rsvQP0flsh94d+dn6yXfDmc3vThH4+azUEK6yWia5aYQaJ3fdq2SMuX5QA9IZMZM
jX70xH6NCEtdFo+RfC+9fzGBXRM2N3mhP64ekmfH5eniY7we47gp6creqF+I1C3+
UZdt9g0MhNe7jH5ZbtpPG/QqTNByUfHfEE3wddt0JKJAjmEVjAOkghQKKg9dkOE/
gzHcixthXhVYCziZTrADldRU91AvD9gIcYMNpPZ5c7HzVIZhwdDL118teXSONhxK
kdOoeGbaciP1w3cN2TB4oV5uAexeqrdfxbTPSpO6wQEenp75d0dG1UFMEnXVRems
NLDZOu9jZGuDVDuoLvl01xDkxGH8g2Uhr0NHEHj33s4nW0xPDniHtaKzZPJuwP00
+GIQxjBIfjDkwvnWz3y0GISnAhIOByBuyYxnj2S5cdygVlQCmD+g19XvALP0pUdn
FC6H2iIIni4Uy5Ba3bXpXYRRaBpQo+db0h9T7LGYddtBFgqMnG+zTizriPz2psyo
FAQPuiik8tVGTb25vZ3Lfq/AjHzTZ+BB/YDb3/ZYMYS5GEzi5hVTQDlyRB3Z2j4O
OZFXFCEN6IM7AgsYgmj7/cJgntyus07n4vMDlCJ9FqjbZ3kU6AaszRrIfkWUnEF1
EhT3kCOidwnmyzRKllz4fVFS8FFobKJxy8obV6qKZrypj2fU1IUWN60kI1MmQdG3
h830Tattbl7Mq1ExJdH4X06c2rhcj0KE4iw24Zd32p9CaiVms4Ib1ya4K7rJ+pfN
FtuFk9+kjYZy2JI0ISZYC5yzVN6+QR7MtTqtkMgCwr+tXysl1Tyj/yDBCgdhkwjq
w5m85H2AZDOVRQBvI5+dOyGweDqg8miCRrswixdCNZd+EBehWjvp0fSfBEJTVWnn
cdvbFbkyz4EHRAMIIy3b7t8DrubA8Q+Tv7P4JzsRqMyRLn5/AWQQ7yxOTwulAO1M
XXGWrNOak/ocbwfWM4TPz5rTt2PgTC/ibys5pvm1E5YciaU1dPeNhIUPlUcbdEAK
ii+Hegexyv/JHbjavO014AUpc/W1kg20Zzb8euryp/YLBGIu/ZgzXEF7CR3v+1gU
ffUXLScT/a8/fMgWSAqlDw+NsZVKPMROm8K540yi2keR1WH6bmZvLrcQEANF18rI
QZ9GWLye6KlKP8Qi1K6i7rHYbwGlfohzb3ldnUrdLaBPTbdbtQ3MAqDmBqCfoi17
7wbMTX8xqX6bC1/WOq6aLaQliywGj3rLwz4BE742WzQMrh/+P5RTcgbgM/Q7BDti
9IM8NeaZ6QLDJ9dhTpAbsrIi51e0Q0cyqvdC/ujQyLDFwnIA+wJrYdPgAEaXxQKj
+BAvRKzp/Qk/ZoLf5bcrM1B9aO0xsS+0VofzIU497Yl5M0o3pHfnF0wiSECM948g
BkRQY82+ft/vKGN8n/XkjxQM2ED+IlufRoqroBZEEcPhKdDdvJQymI/ptwZ0gGcG
8adSo+X3h9WbZjmRMfKSzMkSTsBGAS6V0ClSON+Seqwl6b+0LS13wa5MptfHPQRV
eE0iMx4Jpv/nCVjb/2tuPPLoEmhY9u7dpoyoSiwkreDFey83UeUdOuxieOxW1gDV
TjPVIEHJcw1BTS8W8fQICJi9CwavJJ2RFhLWq42AfjSWFtmQg78SG7xB+eQplYbG
eR83tJ+/exQbKsDx9exLXxvMXyYrAgzReuxwVyeFECGJidAxErTDxM7O8R/WJAtT
vmDl8yVsw4o2bvDvwhpIOKXRYK1gmsVfIOkT4J3gHqEUou/8Cjjd+2H4wZcv2Zn3
5EvZH6rczpVbq2LX0byzB32HNOhSE8kWGsITZgm433hWTf+4gMF41o3t0p0KgfuJ
H8k+qXgT+B+Q9FAnNmVQ8i+FbcemGpH5GJOAW+qqpskG8+kIjGEMPfFYBuQlE5+9
LhgTUCMGr6L0KMgIfCof4WJIAgRspgxvWBaWu0onGhBJtenqr8Kb2hAl8fOjuahs
4ItaNL75UlOhpA/mYHtnrDjKp3A5ovIQ09/GGESkuTW8rIAFQ+mRWT2ZcBmpWT/2
zZR9iOgAhzSvkgStzYhhK2e4Tu7ZQFQe80Ip9PfzKvBB+FrRKJVQg2uPsABTT3tl
8suHkF77wEeUW08fswGAPqIFTCy+sY1Gob7esq86WnOtp8Wg6D0XvbpVx7WN201K
azb6ZeFBbI6apCYugPT7/iB55lwXdoCGDt3Ujm8p4QMO7tlyGBDcmqqd0hyiBEMY
lZ16azdxXruLLZ6SvsLj9SgBNjU0uAbfJ6ngwRrsDn2Cwk732fpfufJXyJhcRYkv
ehFxMmYJ1JHlQ0czd1HOd3PWasLjDJKht5IoMMuDF5MYhgwFNcMMlysh7JSE03v+
l9dQa1CD3z75HcfRw+RltX0rfUFypSwW1PKAiVmtN9gqbW5VYVovK6YPbxCGCSNX
FrKiEiVrJQjMwnT/x+dp6nuEbfU0pUTxrb+zWj9JMo+UY8nvSXQX2lI1aMoFSXpO
4kzJ6P/l3sv+PPzFB4VdLpZJl97jxwG6MrVabrRqvSiCtY7VRjK+TiPAlCl+ISmA
zM/ovO2c/GqnZE1xHhqKcmOn+pLfizCN1Gn1Gwbd7RdxHznABazXjKUzcuA8ZOMo
hLcJKzkUmGErm1hU5LRPFtzSqxk815xyfq7F0ZfZ4/44uVKRC+zeG0hyPi070Xff
YG3LIc8JERoBsV353bgEPCH4lQcM2AwC2eNvX3RfGk/zyzxsmhTtT7p5Sy8Kjbfa
1S+O1tirs9C/4YAyl1ETH+SBdXpOoi9AUNwxvHT/8eMRB5a2m4YXRjjOK8fzV5u2
QuwbmXAHK2zadBKXfYzWFwOm7yya5PW1KiNpicdDtYYMdS7T83S1Ee1qdapVt3Wc
WTn+9pDVjf9uLBT9/LWyQGyelb0yfdiOfCYL0Gv5Gfmhx95bIYRQNvyCIKbhBMTr
lYZ2hOzjyVHAGFfeBuo3su+BLTwIugWdRLBJnAviRLzMJ0Me/R6zvQX2Fn+PuK65
vbFMtpqorV8VsYYFFf0cYednuOPSIpJ6s5FkU7MCvYjDOCjeWqC5QxGaHpqRqZt0
wNsYaDN4bvIzogYG3Y/m9EZcuVF4qMqJE95LN70SF0Utp1wWkpBOp9qtjZstZ9gz
jLe5vG9f9hGeI+AMxELNITp5JrAU0iidIAjmmvRARQaYeSABAb72n0u2vY5ejgz3
qmvN5Kt+/QFBecYrkbIG+enFFe4ML+YqWRFfMzn/Lj1ade+NaCEIBYN7Y4BiD26I
nfbm3xZ8Kh6fovkcRx2SAirbjoNAk4+3vBfgMKg5KrG2uo5op6x9tP+AaeOPdgHB
AmE76LlghhzAvLRVYFBGa4gAKK7iik82ac+XsFvsI2uzSTOUAeW6sX8cbNf60bNB
zdGas74BCDzpK9RSyB7YA/rSg9O2OlD6g0A1aDTCrBPU3HlxfmKpe9ACsvXsrKNn
1hAOgCGkffXmiUjYR9hLFuX5mdQzJHFX96oGS7PRS6R0RcRLDDIdc57tad90+BAB
SgNl1ec2yYJpGc4Q7/uEKxbLhfQKQK7ls3faoyGFyamt5uAe14oAFGOXJlZI2I71
YToFvecwmseUOFs8hy8ONmIsUdArvjlnp915nWzpm7fKq96+HldzR6NTV5iab6Xz
Ro7mfSEOmAOuvpDMHZBwjM4Y9Xew/ORMZM+M9RVUdKu+eMjaLD6Ni+mgX7jhjGri
Y9EJLFBs92oige4+YV3F54r1tWfjzhEko5Ze5s8evf54oHCbMw/Uo4z2bheYHvBP
JmZrZ7VBdAz+6oTwgsW7lkmwlMww7vxbLuwjXVqOxaysEcdiua4yWV66ef78lAjm
qUilHfrzp/R5nK4EiZ/HzIHBvcrVcdKaVwuoXpzdjdCDs5Lv+TxXGmOx+ALiSU5Q
OrVwlY9hrpkyx3F5iWpNIlDJ5dl8BNLNZyaE1L/pgG30PdkcR8W83HAYScgOe+vr
414qI3ELSnYnYhgBsOUuYmQV4GtxVSz+9AZFGCgHkbXue7dezyIqhO3duPdDSpzC
ygln8GnPq47ipex16FLvV9br2yNk9XcvlsUq8gkIganMB8xdDY9VQZCofXmcATl9
vnA0t3HwbXRv2kr1Gt4BdmIdQMDGqbABA9avph6OpeGKt1Al+MNnOY4UhkI76P7H
5y+VkckrfCn30m6CjFLT9DZLDkTvIl+1jDFGddYmXQgN6/6Ndrb2scTrAQ7EHlyS
uq1fBbr7EiUbisyFLfwnM2d8kR4z8bY4ns0bgeT4L7TNcNC8R25fRK4sD/8XHqaK
aXFut4Z0K3+zDvAKIlj9V49PT2SPQ6LmAhztTa3TkegzjdBm1PZgnxRpAhg4YnRs
Ai6uH7goMKPY9gB85RUbqV0QAQ/CeJv8TWLc8pnUWt0p11yo/Xbn1EHIlo5buIXA
8mK8BLsI/Nx5oMd0HSEX1KsgN/USMdwioG797jk8+88izQeUhdPTX1YQ91S58N5X
CBjiqD8AmjWMFgOuiCMdxLRKYZ1r21r9K4JA5k+y4hXKXpn0NPYufKglC3qOwMCq
aMhZBGQN9F9CZ7VQLzDsepy9AO9yJAQFawca0h2oYoWtKJF4tSMDFlnMfJu15iB9
nSn7wddt+us2R8Hku6iXUyp7vEsys8MAneE/ioATkzQz/qrj7/iAIZWurrJisI3C
5C05X+VxQ5/44KZ1b8bBpVyaI6XWbEqK88P+MOhPBzodxC+8Q7iUpzjYLRwWgkaR
m3FGFcQrmXP9l3GAtWxPryP7hZ0o8xeMVBeA1kLdr3QJr6BHjq2w6uCfKKdMODpD
Rqsgca3gD5xGRVU9/XOHBORRcNbgnON5YuHwQm3oT9N53O38CsnpZDHiYtAdd7OD
oxTQUP6rsH2rcf6U6rs/jNT68k4vG5vb8UGUDfuqaygSCUktfljlcY4bpwrMttm6
tHpEJFpkY4Nf0RenCuwSfK2fvHgCh0SyBCebnj/j1nPjI8AOFJi7uyFlmo9gMiyp
6WZ2PYfzX13zq0nfIQ8RDER9VI7U5XOwS4KvLa2NqKXvblYLndHgZMaXEga0luyW
d9NKqukbPNyCzPPuXbXdWo9z5aFuL48Texe26GyWhZglOmgSWpvuI+aJSeVa+HCk
0cHG3EFPrUDhVVqlWaDlixcv5fM4upS0uAtsO4GfKPM3hMpR2vaa34wq/w1uIYis
MD11BI88KaEqWDKPbk0MqWp9HACsuWxe+C7htruENihThmRTXs/ZhR29ZsVNuQ7z
sqB4foBobn1KsMzhyILKpukzxBPG9c467zRQDy1vJD32n+N4MLC+ObZBwlnlbnTP
RBnoS8W25O7MdS2SKe+0GLazBq3jw+T3cfrDnSo/HZLp+02dNrfwgFA2Qnx4fdPh
6FQmSEbj9eXyugPNA66ZldjKcjyBN+wRH5E3DBP5YcZY1nnu9U1qc3gZ+coISk4/
YehUzegOv/VIar2pwSeTr7QBvyZum4FsAKRzOTqKutFVwyAsIAtHqDQFC/2l1E0f
I0ulnYspigfnvu9ISXXLT97j2llJhNai+Gg6PbrgzqLN/f6uhIIy7w2b2Hjrrm3z
iUKxC6/qSTYjt3RO5IMhcjuOyB23IZe+ilW6K+d3X3vcXybDd1EmQm38YCU2jlDH
fLmpv8VK1ZC29HDxSF4OePECVfxHnKKlu1FgYkTbjzNLcdPHRPA6LasKuLw8llNZ
i5La8RPHmK28rupmJ2YSJOfiqdDcfj5qGKwG5kxHfd1K03PIPxgLHkMp4WPjd8m4
zv7vPe0RXDSEcicMzN1QcORzruwhDM2UJN84H4ciMYup/xR2VlKwqKZWK6zWHvQA
ja54WMRGL4ChV6ehPjJvHAnnmdl1Hrb0otIvmA/zMkRVcuqWFCsIB8SPxvW7z8NX
u8uiWtrz9OyCu+BT97EpaFHjmlM/cpUEzqLQ/p0FlzVGfrbZXZ2YKiJekBM4H3NI
TDNv4ybBIJYVWIVUBKBmLLIvabc59XuoyRezBz7WPsGmQf55tAkWZ7hfPa/rY0Jc
W87yWFaU3POe2puXS2/N6wU69b+/UgMZMJvjnG/es4/2/ARZ03/IA3pzW/UN7Pgy
Th1ZJ8CKezzWyTi3i8cftnQr2V/wSJoCrcqD+FfneRLh1mDvNHkGxAq4HO57GFpv
++aCmMHLzSnLYKootsEuoI5XgJnqPyYatVP349YrjnSYyCzX5zNWoazN0rW6WZJh
5mLs13RW50AW/AWHKKNaKRHl8OQmA9Vq6cGEsPGUtvdh8UFdM7eVnokkFvour6tv
v5Xes/9ujPnwZ98uLr+o+ZOI5B4YP6oI3KhuF9Vp7w/AR2MzaZtu6HBnVEb0ZgqU
FRnl1OwpXuOmZ/a3seiWy54yvaLCR+/SEUTb0wjqbaFcT2d+ma21/iBTEm13AUDK
TyOpv68Ne+DTqi8VFHazUz5jRazHFR3BZvLZEscrCCPfh1ztj+U8+TYPk65Z214u
+9wcF3pslFdyL/ILPqmkF2yJiji/jYC1IROp49phw6BPkHYqa/K2MwD/JF7E5Krz
FMQ6j2Na7Jjk5DNNh1sI3HM4tTKN9zbQuIZqd8l4XP/rAFMAZAOvOynP0amceh5F
Sj1Kio+aBR9MM6L3nByvyXEKSCvW5zk5XIMYXF0ylawGtOyUTx8B7w74y1z66lFL
JY+Nj2gvQTI6bKRoGIdHIIvgs28pHatBE+CUnOuRubHqPxrgQpXdcTsZgKGGVasE
3XzVdveATozOqXVWhZ5URAWXZ3uuL95ddOWukX8lBwysGmwkYWNQyamacfRDleY7
EZTvPvA/Xk/g3s4HzShDcNoeh4U6BPCZno9/ngLcD6TdiqW0NSftunXmaS3DidpX
agrIm3TmH4kUJZgic7m+FTlNk7StYehJ2f2q13h4yLCW6lkI+5Dek+R+5NFaXGGm
wdDs66CguGmR9vanOu21cMHuYUx9OZtbxn9DgPiBhecJJ3q5DCAYHD4vrElpFGTM
yFN+FNw+ouoHO8Kj5AcKbyxifVrwuN/ub1NX2hlzLyjZKzXYe2+7P4xeD4FRwJu2
HLVym1bDFVJo9uQXsUMl9HoOv+MI4UFyHxTFjX6wiI7PmniC6lL+Hz8QZELeEJAl
U4y0VqoLpxq9xketLa1UzZU6kXzZTT4NPxfOoFafVWa5t1QqH2S9+SW+j9WSjvMG
iC3OVo0/lGZtjU6yi9KzgezIcoWwdhBbT6zikPkp7q9dRbaFjrYUI0FjfZQfpcfK
LhiT9wtkBovw59qq7zx+1hoXT2/JTuTnqYpNh9s/fwsgKcqsqxO7721biRgjcGCP
dgHLsT0yKJC5LVwTHPwzuZsDGRkzIsgo60FXxQS6A4jlcegTsFLQoA1qkU0sEKFJ
+JUfyTT/l302pyt+ZcOwap9q4lYGIpZ9dhqbGmzamhGD2o2WYwDJ/7G/sqkB4zT+
P0s2lSwWrdcAgizqi+jvd6mDuI42m0ZhLqegkDgJ4XebPczVF5CqWYsF5kveXCXw
Xk4uT0v7nbfQ5hcfFJJ2RL/ELC3z6VWPHJMexs8fmjggdrjOGybqhbpwzf4LNCsL
vLyZVEeFwFdsnb3H9jLRR8oP/fgoDmkx/LNjSH7X2i22M6LfiABZIiu5C5ANO5ZH
qLgxEtISryPpNpjb7kyXboSBqy2HCkAOqqUxz5oTQhuDhMsAkfnCijoEdotX1xdM
GCgZmrhEeED400xpTT8tC4JXnhhCFcYFlFzKGJwxYA9DCuIr9a3qo/rLLVuLcywk
t2egpdrg0ImcyKNUG/orDXXChkEsudr+vGX3hMlQenxqz6wy+KHGr+5rhhOauNAC
Xi3C+lIfgKlrUASuHqnXlyjq7Hk5f+6GfIQiCWBTnMYlX9NJ8wItEE71m2Ks0RpR
VIZUQYnWgWGS1zE8857ONrJo4mkuYT3kzHBXIMtZ85AipgorBYyqrimF1UOjFx26
EoyitC/hyuR2uYVv5LbyN/GIGwR6jez3MMVkztX8odAafkml91sc93yKJ1owXPmo
ezbAz5i+41dtxjqY/PCRbPnfX0+2JydL/qFOOgkbdubT/MfEcNBTYSBJvdsnzkD/
oEahER3PddjXlzn3DLx3nHtqybHwAdgLnomZ3XbmIkFsMayEKOnsL0MnE5UTfQpW
x0EuXFrWZcgPng2kYLWn4lv1guvn34llGS32+FE2RCjmCB6jr6n4S+CTKrwi49vi
b5Jhtu2fy0+M7KhKRC0A1wdg2gsHANDJ2HhwV3DT13n9UnYG1PkVHxgIdWhcpYDD
5vq/ZlDHNeLQzT10NzyUcKsxeEOFvWESvvQIc4ixBGCV11s77ViHkvN6S09a+l8b
b6Jp9uDO3xJkcPUBIY0e80Ez9k2i+IkbdOHwrzjALxwTA8VHQLMOdkngrJ3FEKnd
s5YIfLeMUIwJ7Av5Bs89U8KWA5tOgCH+aWa2J45wBS5ozeAVT9X3OJArDGfWQwNC
de+MehQf+eOkLXoCdSOwCzAP9L8TYXAMZ/LgPe9vbr4BMb9LrowQW4LTfRCh2UMX
eBFd45FeMSWiJYCyteHPyW08gTXq8zMxQXvfFArc8Ra+QJpLFDoV25CEt6j/6rNz
ysraWwD9ewMY3G7PYKe1W3dSX6BdNJhr4El7OFD5w3rfK9uW02Dfl7SjkHAwTk8X
eK/9TK703T8x2K/R5BjS+jD92+S0o14Wx5W5zkyEc0iGxHQFkLaWuBcnJgorxIVV
ozys2nVPDsGcZSGb67zm6KsdNtyi1KfN7Hm5IB43t1oJ/5tiHQ0nYLxYCtgCKIbH
uP1831SMXUcDHEOOYdbERkinke9KvyWkndI5NXmk4AKTMJVkG34TQVPQaG7cbf2Y
raJ8B/YtIyHHnzZt8sSLHSMXmB8PG9GZQzxCJxutN6NozugOCfwbbWAQ4xPwkTko
7bLuUJT+p6hy2XjaV4TBjQACHU2zm1cp3MeucfglzzL5NXl0O1jPOZOIrbUFK3hX
vHkW/w6qH165P2uuSDR6GpVOacqFT1wPuYvuRKxZ28gHy0KkjMFENycYoXXHGRyy
x+hLaLp0YSOlFy6TGVCqf138Z3dweUxmPjMt86nagkAstDeOBRn9z08PHtLoassX
Pq0EJHLfLupidUd+tHgvbF0BKzDS75MS0jVyUEMHsokTz28V/TTuLiQ75IpRQXO0
rJuQo0gcYj5feOWphGZqbW0KPuNxpK2EAICLSaJEnc6LSZEv+Y5sYQQcOFt+oWhK
58SwNoaOD7FUHkPCia0kSNlOC2WCHkFHXE7lpv21APCFNF93uDD0CwsKI+iXav2Q
ZWnH4IyIh7fw1sDZcem4rdZHL74Q7euPeecxWiEHktEKbFvH5vqYJ9I4thAwLmno
RQspKQ0Jau2thxrAYRwYPd5N3KJH2CUZFtH8cy0iAx/2e/GbTKDo6WvOMw17BqMy
wmC7+TXQS47Aw0KCx5Guh5zlnc2RS5qj+vUNKPOlXtcHW+uGpzENO1+c1tRhOgH3
ztIMaXFFr+hwb7xPqiE7QofPRY/CJyHM+t5TmOfun3hIElLT4+MopTi9m8EB5Gh+
AOTxcQIcg2OayLgqzWGdPLOjLmjPg/mhOMThechQw93nNeESGCk6uM7F+UNhtoNo
u5mAyUnXdsJ1StoP0vTWfvnwcTe1RYS1kZ47vEcBYPfb0ofBtXNuAymvXNptLwD9
A9NQ9BYqrxbQI1WiRaxB2KqDlodlFFr85WPH5j0kP4E85I0FGRC0LwBLGw0/bkmP
C4fGx3xpxwix8rJlGU9I86GHkHfuZGaZVn+O4XpRaBwGwUEN0HkleW5+PDwVsYhE
IYv7xFO/RXgJotJZIgf39tYUHkvcebCqolBmbPiMEpNLRSCq3cACfsVhip/J5geb
ktLxboErJ/cHDAOJeRB1uz8aPwZ+KD8jPqLGXyNesRkvXCivheNj3FrHSECI+5/Z
qlk/H+r8w1x4Gj3YwErEWLVgZF79Z0QefXhf5buPoLUElirYC3qeMAM+XJ2BeNAp
19c5tb9EMOOV7CWhMDoeoRAuKXG4shV1r6/bHTbuYTO69o/qBYvzS7SdFlaDal0/
BFdlNKl3lLKHLyaDtW9OiUWJftFRay71zIBU0aAt9o/AMFZqeTQWiHy4XcAvGwrc
SAXdmFMff5a1o2cgJOQ54wMC0GZzLEzBbVjCOR5oQgna7ppu3vOj8i3wHSzoXiD2
eV/LCfSE/Vurvg1tUFJp/6xcFuV1uJ0E7+XBxHsJH/xabH5xxicKHURvrhEeNG3i
nwZOAVkX1WSddo9duyw4DJWC0l2FQgDwT0fFtRqPSutKPPa4r8/6waijMV/O3/qh
S0ATVAIqptWruyAZ+Bcn7h8l4d3OE8aoXuSA8vI5u2aXkSXaxJDeeLKDZnw17cRE
k0z9xkiNnXVTtvql+1tFlmr2WoS8hx/VggGUM6fGtmkEN7g8PLDJRHYhTMjavjrE
P/pjJdzut293TWVf0Iw3auj5OFE2fDHEMhYWESHJapeBWCB7qEmdPwd1M3Qimy2D
PVvjlVlaRWLet3D3qAwdjz+xmtSMqvW6DfFlJ3L6UXaITWEDrWN+rZ0RdCJ+/hq1
t6dpyTaCE0+IeSxwAz0jPltChzAlaBjK36w/RLlDPgKl6z0RxtNq8aGQ3OBzoyjj
zULc/0/3845Eu4npBq4guTHiYMYqBxB+8ycd6cGHbApENrnrrS+HjTvX0MImIm+8
jGnL1S7sSZ9DCEjhWOdOQskhcRDmaxnPfBWccllWtbmWB/1afD7HAEAbo7R5nyGe
rUFxLp5eAsr/gS+I8hX1oeyAol/+VNZC/p4e9U1bW+ASdZ4CtFOQMOFrTqmnp94X
IvJtWchc1lWGJEIURJSt9/zQ7gpWT/aBdbO7v3+m8LXPGYbBA961myf+cfpsWjPv
Gu7TEeJJFCeiNQYmPo/mJm4g123F0omfa60I8vHzOa881ffb2AckqxR9GQGrXygg
zl3fHN646KArxjhPKjRimsCRqcQ88Kzw9SVHZRAxWLJhsyd7wOQatxOY7UB5/SYf
+B4CcRMU6E1d91GoI6WsgOwsaRFd9RM9Z4I8P2CSOhMDqWXt0Du0SikDTbg7FRVL
CdKm63P0Q4/K9wWMGSaaQDGP4ey58YOSBbOVdkXU+cxTQyPg+0vHBcmsf2wgAuNY
PNkdx0iWmgTUOUUmPbY+5WKVJZs+8JlunfZzsX2o3lwvlACEM5XheKdQkfKat2nv
/451uIXAjiFWl38m4ePoQUK6B94LOnryP6YanlXc64BCXvAO0qJUaSJrdKKI7plc
eCIP/jOUcmTjpLkx9kR9UrQrDb2qM33sby1FxpAl2COHx8kD34eI/D3P+DgXWIem
JNQfV4e3ATrfy+TCavx0LCzS6CIYbpm52aCqNmDcj/31Vf6OXq3H3eN7td539vhZ
YTAZH/mDHzVRSHrzOWgG+1xyOGuFMMg0663dpIfTPzfIVurYOHH/XHbJOcFVyo1P
QtAH361/fkY+/+dpXTioQfuPSsFKwhB6y3Iik7WQ35/QpMJAP2OqCshlJE1KHAuz
K7Bd/ripvP2jahklVjArbqzUSTuGx9agXyZXaetYGg9dU+wDZ7Sb9FG0hGrFm0Dx
eWmfjKH3OvYppdQ4WC1Ltd3B0a6oyVaAThzWKhvb9EqnSg+bEvO+WmHfojagWqTo
nZEO7f94xKIr07yZSePi3h5usqpB0yGCvNBAlhaq0yZmy13VXCbu4N4qC1/ejlEG
zmNa3TZeZliTFuUhWCzpljVsGh6EAA3Fgkf4akrKLnNVKBD0iNqHMR6DT+0hh5B3
TL2tTXeqIqEtHp5BD1EX5eafMGzUEqC0c4FWVdns8/E7+HhhxHejbJ46p2U6kdlY
RM+aHoQJ3hs7NfLZKMwpjQ0RynQG9CEjfWHxCMIxSrnrHWWB+rzvrIu/TnAklJx7
c30hVEIbzYyBb/v9UQrMVomw9Z4FV+YWKKczpp9mQ7Wcc37pToR4FL4Rejkkics7
KpulFpfytcUz7Gko/fg02zxE0Oy4V4LjnV0bsH11X81YBHPch8vTN1UfGveTiID7
jVa8VjQ122kOstTQjcFmvxcaWq5sAGxsspn0gO63XsVaToPsxQFZNGTv6HO77/nY
cgsK+tXkCj0B8OO3xEjdSEXeWZV5566ECqTYcPcDlKv/PB800n3sU8njn8r8FYmS
0ZqnP/fLdCZAvu4650n8azVPdRgcVCi4gRsjUlt0ZmKwYFoWSa+f2z18r7y+GRRs
4fPATgj9tpLBA5gjp7JRBTVremBDUV0OvZhFBLeZAWY0D/KdmXTPR/Uquu0vIRV7
xLfifAo7kRfTqN+sYaFTcvs1oXkRu7yxgq6TUPh+pmA1+FgeiQ8J5pHgjohwjztT
FoKiELyPog2PhDa3qTDz3Z2G8azTiK11msrbu9sVdVCiuQrBlexMQFfF0P7Emu+L
1JotOWuFQBod7qsR+/h9//xsjmVQhQfyvzrnEZDYaEZ7DYRpRfHkldR9QQ4itqsL
+vWzOiHLEdn0Ahu5+fZDbtREJtP+ZXwktOzaG/nIO7NFC4cbO+5t2RU3+OxNUrID
Yk0rn9iOJX6ab4DUkgTtmYEtJorfFidg5i9WVPalxOiK93or/dQQIHxIoI6zQtms
v24UBNd2ggq2+JAt5Cv+mhhFngJxrqztchlHjIojD+KrsF4nwu7FMDu9fF4g1CqT
4Qf7d3uIxzvrtfODqlnoMiYxF4FzzDyLsO33gMJxki9nLASpoNgl0ChUUic5hlkT
ZfJVc9UeaPRVf+0gU29cYVOYv21/dyZRLg81JMnXWErEcj3ecy0ZZdpWD7YMa3F1
to0NkCarOFp8KUXejfLfJDebcTh4MAA1KbqKkmJrqivXCzD4TZv9v8evb2ev0ic6
YCvRRq/zZ5VIlOrrsNljrclFwN6/u3Ogf0EzfeEPJ0dAfMJ5FEjYN1whbkbVvMBS
f/Y3pHhGk7IO+bW8msTMX+GLXaO0hfWHTlJONHEErhygqa2j7sBUrE0h4kS0bhMJ
5qoUiZxE1BhBeRnbAj/qyxihoP4LOmeyUg/CvXC97hcxFUTlYlbvLo8W+0S5Hnzy
uYeXOsaB2KGmMQyZoFS/urPGc3uDxVJUJO5eMtCvEXC892oKUZmsutpo76DcKsST
VBMlj9ekH7ZNEnypekHBmjK+qpzRTPzbEg/12aowzEuFOBp/wKgHti8j+AC+SdP1
1ZZPmEAPbg35OGxm9kR2sYHBWNBL08HCEkH9Ac6kG9BZdF6C/YkRxY/tqw1ywp9t
90gfEOY5vSIVUi3MrAudLJvI/AMYxjvP8U6p0c06sho9rzXfXClwPjhObeWAL8ct
2maqvIJxjYfTRpO5uPyQq2dzb9Xd7K3gqQaMq+OWOYr4JYqvHrb9CnCwjMtzjd8U
sZO6y3rIXNsL0sEADPtaTLd5hN2kil0KkaD/nMBo8oq62l5vs1vb3JjnpZ4hf+BN
Ar8/mQo/Y76J5pW39gHTCv2GdELfIuQDn+YfrwCjxs0rmPIvbhNDs16tAjigjiyd
o8VN8TU++W8jbQ6iHz3LGuF0vaBqKGPC4O4T1WoSGvkhnfqDRRRsYwdmiubVo9JA
f5Y+Melt0xL3Z08cJkS2TMRQuNsHy56LKbTC80X8dwSVUO9rx0fil3xxZwbJncFa
kHDW0+F8JlZWq8bkOgNJz31p06tFBHGgFfJxfRkoBppMMHLp33JCyjXzQ/lIqLNL
AGIt7s2tDntns8+Z860D8UUAkKaJEKLT3dawFAzafKzGB9/jDvBu7S4J4QG81hxC
7wHjkglXRZ2n7vaHfjMxBz6uNi8LOf1nMhPHGyBUXlS26bM45rOcKZc4+hVaVP7e
n5JI+lsrcZIbjac4UaYPE4t03MdIw1DfEckH0WvSEjGsOjVSC1Pny4xytukQyQYH
i9LjiPU4gFVoEbusoRKbabeMcH8bmPtV/4JYTSuvWrGyepFSiljODFYY/NPh0B9m
lpuFJbt1rKYOa1iSK72MFWlaiV4Zpz6whfs7huUavdw63HjO8IHwzS+57Sr/b7KC
3/RSvCaMjofqGzml522PZ5OQZIk71HFqDCPEvNX4qdt/IJE5N9dDNxct9x4RPcqO
4tsqwsYADyh2VcNIniD8vz4VuqSNpgHiSGxTrUYMdXtu6X28r1L302v+0jYMIdNJ
qxtLUWpds7QAtf3Ronkvp4aB8tn0S0PeqwYMRTbrycFYap4PhFibJRfE6zkjG2rb
aFoivUmFjRQ5OxqFbQcf0pWR54bnKDvD2tV5b6Q+6tMv07OxuYzNJ2XIWq1imAdp
anJBCUEwe5QH60dNymKzi2CXdsdq7OAI35gVL1pe2lmVItSZJyFrotFGHmW7iA+p
uQfc4t4/hLGQtymAbkn5sa/TtvDa1bpdSFcpNbVXXTKjusqGdmpmDOa9ISgWI2zr
ucQQJ3YM4mGjAY389RP6qdnO9j6yRWBdfseaNWVHnnIt3hCRB5zzGcgEoCBL1ReA
XqfDGMjRy2AfUEfAYxxE5MixZAPI0wGzuqTm2FajzTZvMTL3gRYuoI1rIcmkldZL
QSZDONt8C2mF/sVWKPORtFVGxzY/k0qFUuWyEwEXTwf2L9qXhaazB0o06ZjP/1At
pgFpZVhcK0PcdBiZUcKrVeGwiem5PaaN3+039znpydhARUJJkfijr5QbT0pJACT/
wQNY8gfUfPyUgmzyzhiiGnKoi/GGZZq2Oe41pICOgfKevfJrqQEbVIr0lGPOPf10
kYhUczi+b/tyjS865iBkpUcYySzzfmUMv1lFUMpCwj/JgPi2pXzbKRPlcz8T14jg
`pragma protect end_protected
