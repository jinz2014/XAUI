// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ywoft6EqHXyOQFYU9pAnFMYRQSM8vMUVXth2BMCKbMCdT4Lxpsev0KQ4lNl6rVtJ
m8Z7VGlxZzgLWwIEXdOqP051MA7hn0olNfi0RSkkj8jAj9j1oT7FOgPg9cKSgYQw
C1cgIpNpEUA7xpXbyt9eAzEmfypmHF6hyxEcvgLsE04=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6400)
qnwHzW3ZP9jGsD2OjGuJIM7j9u7XYDILxnS0uOoVKHpoT9ujNhFZQ9owxN0xlmSW
q//tqkbb0+3/Cj7+h3WbRgl06En8gJy2gFToHEHJVKa56Ta/0mBG2bW9roBi4Exs
sNzSNpmJK4a6l8xFYB6CtlE69K9bFmiJq29BPdgOBFP3Q8EzbDCmCgEgIDkahjsU
wpVIOBwKr5kTmJ2X0Wqvqq3uGIZASHzwNq1X/zLq6wQMOGIMkL8EgAwO0HVVNf2o
qMga1oNs/rrodtUyAPJyZa2mKeWQC/f1WNgyZq9hs57QiUv9GBAupH5CDys7Tf1v
YmJoUWAYvMxZq+6je93mE0x5JlQfRC+8oNWUaMo1Js2qwo1NvqknUfWg98k4qi1n
GA4JtiejsaMxYtfSa2OJTwrwArM69AQSfzGw35kWDXWtEEGdYSAcu6ZXr+ILUuqc
TlJ4Cb3WRNjp9qkiLWt2gMRHGwch/ySuXmuuZarOU6UcDSo8/xPTNfk6rJd7x+yr
4SsBvTRYf0/kZYAwsJMIe9M4I11hHH/jrywzbLrO8oZ07zB1+XFM3F1bPMBYQeMH
28KqSY7+HHFM8to40ohMG9Jj/qfcQUQCBYS5hM/mZQtfZcZP/iJ694u4zolazF6z
l6+YCUFB9BDEnCDXvxhR/3ToxHVJ/MnUM4WZljnJu+G59IwF5+5FxIBIDHdtmL/e
vvbzfrXGaXkXey6aMHJSqQQLPsCMhfVmuYPKERZWJUPOazX8Yic3dvIhgIjKMeEE
6QLPzjhpr+8sRKY+eMk4V1kAaj2PUpLt3SkH99Rtn2qXeu+9TuwIH0kTc8wNPtJP
czp6qcIQKkrEMuJYTxaKg7nG0AjttwDhk0YFUH4EquRwwKj7YzuMXZfPDjzPo1s6
q2Rf9sp9buwVS2h95+DX778N+IplUKbDxq5cTpw2Ubw/reyHaIn60knkFIfuVPnE
5N2uBFfCd6Ju7q5ZtVb1wtLyxWgqM95psniBj1YTVmo8DrltJJQa4RqL+iVckt1+
4VFLqocwJ2oUxMa4Fg2CZtShthIpbAKgj4I2GYw9yGbfi4tUDX80h4t692EVSOG2
MkuI3llYM/b03SCeNBCGdvAannLhNcwxulnTkhp1xh5mNBjZ2aw1tOf7wjCjEivJ
DtB8F8OOV0WhLNrhBoJRUYtxfOUm2RgIwESf/vFDqyNjzVZFpQLxWhYb0SKwJnuF
qBMyTakGim928iCTwsF+mq5FVi/re6xPNZZi3Nn2go5MHdjCwwnC9mL/VIDo9X0c
IBbq1V/mJfaKBddN/VaqcAIjwFdrEXLHR30gB9UB7dF9SLiRCbJKs6Wwo6/FBzD+
JjCVjpNsyQUp9lhs0ILMOcIxxomcCLkTMxSmvmF5DnX/Jm6qQOYFWmJaMSxu+pxj
BrJzRGsBnmCMrhwIM2O2l7S9+zuTVLQCMPKB4KSKWma29DuyI784BC3sHVN/oXl/
HALhD+clFyxjZT/K3DVM38Np5DxPs5xsUZPiC5bbTxJ9YQv7si4uOgZ5vnJlTq6V
8FIG99oeFLX32EUF3KDEBmCihQ/BqlXloa1Ahx93x1yCekWfxb6wFyW6vxzriOGb
IK/z6yjecTzSQpoH5iUNOCoPLtZi0Ky+ohTgd5vUvAM7/ps9AP4Zz22reuzVTN3A
TUFAFdCFxWXUbLWHtndbYIl83bw1N7DeCFZxlA5HsewvieNUeN2bfwI9JwgYqOCu
9h2bynss5QXAi/bS4VhLI4KKTHp2Jf+n6iyyCHCBWVZ5cjvGMYJg6D2tOcuzffPt
sod16FdNWMR1d1KE0UWGk+NQivzUMshW3xHQLp99ow5netyk0Mtq4ea/IiJzDW6q
e92M9JZZMXoeRlDHudmSt9AoPkmgEMSwexmhZVHjw4SzDq/g6nF47xNWPugrfDYx
wgjvZsD8DdSwXAd3CGamEa/rSAgR+AC9KJxrs7kPy/+3hecJmsq3rDnfGXRhzDtr
avzZf+qvxtUGB9phlSzu0nbVUbYdnY7lHhByLYEXzizND0tMu6XEZR6f2qPxIVpf
Y9XaHERrtvzPyfETsTzP9tnYAuam+t4kl7si2pz8TIdHtkkGsWz+x/OpcFwdksR5
7fPQFYjsGbrWNKAXu3oplMYqx/E5xF1kIUMkU0sjiyR8rDhQk/DInqdllwhyxpqZ
Jv/xQrdq/yXA5X+9zDVdqHhEeP2d1ygU9ML1vG6C8JLclNMdl7iAcT87fTCmlFYQ
8lq8yXkq3Uyt0Gm9BFNxdXERwXNmYIeIsFKFe7hnMYlI73LkVIOGAxhL/xFaWgWv
QSuyAtax9UnSNpd5uNln/wfnuObnUOvOSJGXuPTTDmb9ZC+ud4stXttVhcZgOlnf
6Ac9i5pqJBildHh/HkADvBu1inxtwuJgUVBU3BvGGGV/C/KFHGP+rmRJvZfsOrG1
nwEwg0c49p+zesw2ozhTKK+3NbGnVueINHYk2Amp7BdMzQJJCa6tDGffhIVGPmBk
PzTQ0K7hvi5L6Io7c3f1BLAfqpdYreYSkMVHkNoIo7hWSLgZZjmoCfQVXd/hsLQZ
2Wv4eB438iXHGQv4lh575/kTIAMLyA9+YhERBAUuiN3067xs9nNy7k84sABhAj7r
aHlyhdX/U8DOe3pb5jprKF9iW8cglKub4hY3gS0X2HfVYLUV7yv2nwjj9hjIepgz
e4uhmX5SY4JxT+k+xAv89ySVlcr1XGgVg1v24eb8YJnx9EMbezXtrnOi+HJsD7AO
MEba0dxqLeYe2EiB6Fo1kQs55GpIokMQAp0iYHtkGDhFzesoEtvR3h+DekSva1Bv
3O4SJRrOXg4IJwsg7XFoQ9CHAbumsqK/36bw+M/PRB9iI3UwUAlnGd21IuSal5WB
rDBq6wh0dEGPPd3OvfmsePPcp6KyDyGfCiHxW7aNryVGavTzbNc+jo2U6PgfFAFF
q+3NFn4YN7jcYsmkETpr9yw6JQCGzD7EOtKezbpS5XxCnXiWLLkLiWT6ZPVeWfqx
QL5Kr5c60hjW8Im1I9m7oEwXTvJhCiq82L0gqr3ldFjmxpboIenRyIGpGp/qQxdD
l7w47uM6IkwfDpKa/0myq75mlt33UsIPor4yoJua3QWg+RnT0TM/xbrPgXuTu9PS
Yib+TCZJG8E+HT70KoKohXVOcbrrZldUpytUlytw/8PXMMAjUzMhynzSv+cVleTS
sMnAq0HiXJX+QXD6XfUxuJagVr/FHM/+2zR9HjjtOBcGajDfCl2Mx9igq5BOMaLw
zoSzib9L4+DJPIB6r8DpmLpBMDypGHvbp+mz+ddpOEQcM7QxXlGoct+J3BokhbMw
/XEyuyp+47rbGrqQgEphYX5gZyYGnYbkiJpyUu1k0ulLCyXtItw45CFS/E5Lmjwd
L3CwAzLI13UFf7iHRpsdWGLWbHEnnUH6kVMNVmWig2axJFajEOLHbW1csA2ZkH6j
YY8i0barMm9ymLP+N8JWw4G4A0OY8k+TvbQroMuFkV5gwcQbTapP2pvYcsriIkcR
FSntXC98hrquWtFzZDMG8nqV0oLRLAuYxpS4jFuvgu/+q014OhRbGzTFLOXeS7Pq
kpVOtWTXj5P2htogBF+SFU8wXrJTqjDt/7UyTdLfgMg08kSQO0jWf6pQRH0tE37R
L88M67hprDYs3J0xk8Gct0O+JOBK8PdN5WrEbVrmZK/OibkdYP8aMzVRHO+SZc9r
QJ+9gfDa8mw9XBp+vApn2f+l6oGOxviyCgQR5725kOL7woFNVchxVWguUYuu8j7M
dqtUxoRnq7L12FuDtgIKEqa5+UhXqsgHmPM6bb2f+7z0QKtrGLGFQLEwvv5ea3+Z
i+CqL2iOeMHA/8+wcfL3JjkegWZ7+NS2ziWWRKwu7C20hG3xmNiTbGfiaP2rx4MN
iMCYlMr6o2z9f3ca76FNJUTaSyzJ/3fOhyHNzRjyxOPjDqRu1FPQRUVZItj6t/RC
WIs/w1dO2isKy27ySxOiXIf0L9zV/QOhv3hr/WIZh4Ic9J4xbAz9J3NvrkCsy9Gb
IGewUZ5Tt+M858lvVSW+URjLkIX0mENRfDmS6tAC2LuY4PUQfNJGl13X5lfa7/QR
DCXuZ6GcTKl0+TmMcTdfr4XvUUjLUXQ3BkC72l5xsV5hW9Qu/DoLmFDQEfmPXAUd
HW+dN5yKWXZNpwst3e+RrD6phAAfnB4hY1caNKH7PMO8lNcnbIQZN93PIp61wVFJ
bXddaBTG6QvLKa91CijYR4/3KyDOpiJf98JZwqG0xN0Tq0/0BW/XtsEMTIcon9J2
c25s+PRpU404R8DdfO7aO/VWTjA8MA6F+bDSj9A3OqRTKw/aEIC0X8WU7AQsg3Gn
WOFIYrzDA+lhZyF9tz3/2+8ynwLpZyHptR1y+OnY1dgPrRvJMGHZfYNSkeco6nwu
PGtRm3jAjdVmTHiOGB6y9UEIcq+d3AmI5+lOUt0sP9FAjp57cPEXq7p9qtVIuLxZ
657nR48L2lmxslhrkxR+SNtywH/KGrDi/Xr60u1v5mAb6HitvnJNIZAbrTlUgMYO
az7EBbbj8MsGjuP91JvqwtslpcTRiulQX9FLj4p7GaYhDdGV3VkL2XmrHR/nWP8R
3tGNfLO2/VwTFMB/pOsYwDYW5qz2jQJkwIsPQbsByORoS5KZ+cZ/ArOD8lhHbmB5
2UVMcoUD/LpxxE1RmnxLfXJn3nUV2HaRHF/3JPABLjHhH1ekQPhQkr+HI95lNndt
d2CuQxE6O71bwCA6dOGl7D17QF8nVdym4G9wekz6vXH+8mcBuCeh/r/yTmlaRo2I
iwESLPppLUoR31aSblIL9+b19X00NLcFoY/ZRk5mLTlTW8uhmoaFDBvqT+YH9DRa
rG9mgnmaZXqzrAHx/jnWFwtLN2HUa31Tm0eOYvUgvobyy77UzmSKCTa0me9NgTLw
yXPN+6FD9TDO/DEUCCpWJh9gm0vaKel4S8fAhidSSxSzqpj1pnn3HsjPiGMZ1AOt
hgNbTSFs1UOuAe2/9BHIl2NkmevEAVaOOsNnrZcKqyKf8mS9l/4si553R49BceC8
2HRUtw6Oiud3tW9U49EhNkMaxLNpdCwjxayN03Ieqk6bCmsNUu3IkCHVzUxu7fpE
l4SZS7xxJItMDVQYi3RCFDwZl36Ba2G/sEVn6uRFgsoSWQrA50Sng4curn1E7D7L
5RGHjPwVa8E0U1SAuse6hg9hKdomxXzRkVmckCV3g2/cBRTdt0DrMxi/4BjYTB7c
SUHD90u1WLjMiJYpOTc3QIIaY7R0wu9zkWwX5W3HxOwGzsjm8Zzi3phm/j6u6XkY
O9DJ8TcAQdRPWiMK5rYmu3cbm6YINXWVokUsggVASFgNSb/UFCdA4iN/Nm2NcQYs
Bql62CbD4CKRStTuAR3BIT/ZYhe0PFQzk5+W+yVBh2I0jua2N10HuokKG81c/3PV
SUEhM4J/jYO6Jzn/kynaNAsU6MC8eRNkUK+xxBCW+RNF2GuupAMjI0NBkeJ1mQZw
vlGYpEhRwr7nC6OtPzEUzAJgbuXWfyPIOlw3yz4mRHSDS3T2HPdmXGnGeHhtgg9G
ZU+h4kMO0+tXSAsdBkyC0L3vd1uybyfqyYJTv/bQFQPjMWt9VoLL8lGyq2e2xtYz
GXSnEmPE1x2reFz2RGpcRwip4BJ3G+OD3ukBERyBfvmNDV/FqEUNQAjKD0ReGb3p
oU1SeZJJRj5TxTak4eGqC3LQC/xlIthdw23X42xowhAtnvRSPLev4C4GzkKO9/lz
MclqeOefxmJftiiKWZlVVHo86VD9U1nJquuS/fwAlb+aPM20l3yEvZ7XYmyMtoie
hoIZuN9ggeGvs8iJwEOCwk2dpvu3xRw3ub0WIPhNPluB6IkDRdyX95g/eGIjb66i
DVubYOb9rHV60AjEA8rdQLp+L7Guf2SPZHgx8pMqebwbLe8PkWScXiFLzkIwApSQ
4ObzM8mHayPX5nIbsOuSdTxFQnlI1Avv97zMPaiOz3k4qFKMzeKJanHlA7rK7dqb
Yg8r+qZqmGu2uju+gN/K9te4Mwaxj8E8rj1Wnnufu3PM2berQak8K4/vbwKtoES1
bj96YsCWmtSskD7/OF3w325xNGoRuVeMa+Cyo0eHWrkVbMRBCBjhZnpCtdC3wRVQ
+cr+lLW1gOUwn7iewstzZZ8pXvvkMtrp8/Yxbs2SyXPvWcf43A24FAO4O7CCnUsd
bAf+j1vbObxwpSpaghfpGBDP7ZivxXr12NSGdkUcINt06vQnAn7/0PoYbBz0eHuN
cflnWG7CRbNZOHA0t4yMR7vlHIRe0yPNVl8NTS0s+pt8yoJTT69vLKMQ4P7HZb36
gQNPZWz/2yxLKng/zkjf6k8ZN8NHHB4zKyYWLhlSRR2Enl9w67cTQF6q7fZJ+tUc
eqGfLPYAJBVBrFk+RTguXB7je8B2VqbFOh4bxjWcVpY/CGQm1f78Lfz0hF9sWHYf
9x0VSBJJaL4Y21BFIIHftdAcrhaAPcQwDAmPYsumFShoXxRDhtGRoGYlvDzxVaum
erZhg72wpbaxwWiW2bxDhX+X9opajqtcyX9Ljzpb/Nt0+KCbPNAMEAinfS+fWz/k
qnbSBHXN5JxrshumIb6/nZOqT5Z3BTOmCOg8Tkw/xo+gGKykATxBBEY5fojJndXQ
3xfCe9S/DobVT+i2KdkCRZmkTNa8uVbJKUTESpIPy4/by66JPB2EOMy80Cvl1qD3
dLakQZlOKnCrNdgpXQC6G4+VavUP55rWXEVg7RWk8BuEbxxr2p1b9nYrTh50YpER
adkTH9vWgeMennScmEPJ+Ucbuf6CW2MXLh8+Dzr/og4O9+cayYc7qv0u9deT/6D1
irC868yEcH5CzJIB5Iz7IlF5rH0WG8ZBogu7P8POMaS7M65+YncNq7/ewpvoWj7R
ijFJimx4KKicAkqMR46jbQqwc8fi/tLdr6IiTj5OoPxlh0Uz0F1BHFIGSp7+zEFL
GWVzzfGexJ2KbEJZSIWYnawr78VpjHRhiy9U7CLmflIpQ+2QyQ8DC8MOUVHZQo7D
Nap1gVholhpFeI7PLMq71Qotz24r1J7/Y/6nTE4yYNl0uTaLBo1JIbknsL3OyZY2
mQNFCecLxYgYqwawwMIRmzREdSADLNOoKuPiz/7ydnVCQFooqFg+PXNcbiI0O+Ij
0RkRI/xqnLfQAvkcPpOtXV1VXjrtmhsPenB9/qa6i2yrHqTE4MgvQ4KOJIoz95fN
us534nnH1k3EyFhko2imqzboOBu0Z6jmH7YLBo/ei83aUIRNib06W3iFEBgQRV1a
EVhwRI5CMAS76SUOBljCXz+8WixEpWA/IIyafJe3XV17VBOGYs569EKREWJHhL0r
8fBgVvsKlV/nmWJStWsf4FbkhCe3qWwhNxdrraF9KvD8J+ZZc6kB2QKZkTduyl7x
22Ata4EzkTFCraYlP/m+YMXKFQQKLjHWXVtQgWIAUfqxnWqSztIugfI4AxCJ735Q
AvdlGoo4UTIZCvIFDm+p2wpzmVBa4uNegL4arHgFOeWfkWphDspIsagCChb4JfqF
5TTap2OKqoMEeeJP9Fh6hMHAbz9F3Xdb5QBEKPvZlhDRc5H69GKQrTL6poy/Vbt7
MBi15f6uKztkct2CQz3FixWoLyaMTLpvJwoQ9f54+KwC/CPUzs7wihxeAR7i9L7B
jcUHagYOsrVLIQjF6t/9ZiTYQse0wghnvt6tBPr57fG4+0WOLUuzjxRZwzvcW7qX
/SG54Tl3l0AaKIbrEAfW4NKH0+gK/dfswCBEvV6xU0WzI+Y6Fs3dUviDQZEVONqB
MJOmkSVB4mReb9xd9/3KLMHh+5eRtXXAWc1hjWeBxryBbh8TJsnN1DSMum5J//Q0
OVAVv4VPK5SEkxH3ca4I85RAYZjU/inCz+3Lulg3yg6ilLQ9pqAZi7Qfuh+9xyqh
P8tSkHVf0VhEw3HWqzHrxcYOOi+vNObx+JFkrR4s2Aw8RAMx/uMWmtY8zm4+NOjY
L11WprdSg9iFIBv0MT8x8k3bO0OWDtGItEvClmdHS48bQ7vgi5DSGBehPcdC6oqZ
2s9rBKUGe3OrXyOf8PO5hoDLLZFFEKeD/IV4ZaIHdB0IdyJQF1VsxhEh4GN6O19L
3gxKvwGtbYtZzyjKi607lBG+xyHDQi5TdNdqtiqEwcUhFrY9k90VA4Pf821uFXV/
71sBjOI3agVOxyZUooIgtpTxoKwa7aP87B5JsYjj3UdFlVU/F7rWwHc69St3jbNv
jNgEuAQoOpGmWmgA4ynmFuYNrfyXtBpPeNga0STe7vA/kM856FfjC13Hq1dXSeCE
p9wKr/+gX73rQf85rqUcNr0L5OGK9lG/wRoswXT+JiQaqVfUIXEteidbiVgdUaAA
dY+N7Sorl9HnwH53q5FidS0duMNPO2HjSDzPtfolUuu20vlEIN7ctag7GfZUmJ+v
HTIg6wT9G9B66mAZB/R5Whfy3aIfmDITo3CLPwLHcFFrzOoVSTjpYu9R3QADJoY4
bgYOafM2HIGoecBzWR/AYw==
`pragma protect end_protected
