// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C66h92zA93C87kCLDHvgOUfvmmAT6T3RRuaTnoYwpKH1xnbrA20WSnbfaN3INzNN
KN9tlXEbmXAx5whnhJtW0D0VXjScRjyXHIJNpIl4lWwyeEpE1EkYF4VgICMIjgVW
jM2+xeORMlesxzs347UAwVgz8w9sfSEdddV179shCAw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5776)
/WLCFqtsWGfwdFhYwOr9VhhbnVe1g0huMRatT/Xf+pHQk8xx6PAtpDhKI06q7cXr
kZNVbS8SfsHC8Bupf5nm62b1/wldzK/oxW0aUu+rjBah4F/RlGyooDPoyRTCjv/g
s5Fq3ljQn+EhkPcK9gPAKUUkJH05rT4hyISpcJ3nhatpitti9Mud6IbwDyVOcy/P
aWuYUFGhA0sPB9GPwN55JWgKTL7ttn4oWefQrrwbOjLHIuK5CgCodp36qUIW704v
MCs5RRX9xDPlObL7Du5f5HHMaG6shhwxpEa+CY4hlJsa0FjqPOMWxy7DGqXWx3TN
EWf0SEB/VseJXbIy/KrfO070udgQOvtELZsVN8XRZBf17bpUHQnTPvd9A2xHh26k
UvGtT6h3O/5J6XxCHW/dW9KGyKeU1TCZ5ohGtpkmu4JSx6VsD/QKnFH7LcHqUB+O
lZWkcU+MWwQ95Wbu/FJhTgp4dKCocXg1fOJEE7Bmdg9ZDRtRFeOWUl8XDffJUbjl
A1WgQ2DJqTZHve1j1UV8dAylGBwEoIGxt8KZ32YFbSMQzunHm+6F4oi8ZEsyYi1M
hJcy6luHEKEcEY0TyT/gLaTGUOG0tMXm2qflKo8cQ6OlgoZaDn8AkjT7sKpZq75x
o0+nF3ONQ1+J0FvMmuMM/0cnNoiPLHEwsQYSWmu/xyuq0n/RVoA1JzvJWSr23R2w
wjNhhg4p7kpdk5hdj8ecPy7SRlfxsLOyBCsF+7ZynZ4Kr0KkjG+Ne9VrgxXYckLX
MqGgI0xkYFmThQMtxTbclvU8v9iEuRxod2BvxS3VkQt+9U2bFoeA5uyLt7BgP4Ym
drBIzUuXRqp4CFoglffCxDIKRHYHQyIpStan1WSrqu6dxhv7fbOpY+TqfzXFsJHq
fUnzzA1nJUN9Lt7PXMJcYK4ZL123u9e5X0Vml4MRN3SzeNGXv9G1lAbvPcfTJU6q
N8SjwLHyZTUGveonRFEzQv+HAZlMqebjSXd8PGxwql/gZ+7i/irsDP4TbsAz6z1n
3UqQ3WpjAm9/0TYdFiBbIChm3PS69voFB2uYDulAch/jxjqFsHfav37lUETC8ppO
/qzmqpjBu4WCbClZfHiOtSsEURN2OSrphHF/EESU9GSHKkNi8Q+anNYQFAslGEIx
/V36Tb8W0+Mn+r3Wv5ywYdEDlyiBIo5UBlFYMTLCItiXgRTffzwfX3CCmaxry5l9
RftlynlPlrr+acBZcYIDZAWos8GWK8VsdHO9kTEEvBiEeCy01ssVFOzF3SRdv/IW
nAdOnhCJvqGKrQoF6WgNqb2UsMKfJ6n2dyx3fLHRVyeK/bbFrzoCBkvA1xRAhlzR
EftSGG2VxgQVUqkZVnI4iEaSwvvccxarMNzecLt11W1bq7R52F8lH3q07tbX8TTy
c5WAWtni6p+tw1/O+gOH+ZnrA/H1DQEXFupxfMK+wJDe7U1jLHIvbKG5OAxW+uFM
Z7HHRrgnj5ix9EP4EBAH43YDHMY1bQolmKEsoUf3GQH5fihdgR1RIuGQXfZh/JK3
H0641k5oLiEcnOyBVhhUu/iUIrqo1yV74AWfR8Fl5bzeC79VuSsW6h+6f6lm+M3h
pXamYa2hyh/BKU/wdSO/+e3Ao3Nzv43MoAljmnIrEIC33NW5L5DwOwfvEALXmqG+
LT+7YIGbLhlm71AtvEEP9kzm+AU07sSKnsVdj8lyCBG23ZrvKdXGO1zGGvSjGPZo
hVMdTSVjNKOvdMbT2nDKYPRV8rhYuGmFflHh0KOV7xy15kKIAWoW5+d3LbZ+iBvA
oV6vWNYnUtQsvRDX+m0ALy0a1oHz7gEJFZWXvG/WfJABKRpsvCLqOa8dxx2JOZz2
tQqKzC7ezC8jjboX5klbldlltq3OsYm1TkcSRiAXd8KFcV+Hek6c1Aiq3NYe13uL
hmcefO+yghRYwmrVHMdRbvHhZMJspFFM4ulyv3rWrFRDoSjMgiAR8XG/n2XgZwXR
hYVWfX3jpEP7vAbPPMD5elfXehU5ds3wMm7jjR65cJMiZsHblRrGao1SDo8jjLru
HsDlaPE9nnqjwQp/P2MPEp9uBtqz2K/msSjuh49wON55A04QWpoXH/BIkBKOXeaJ
BXXJovLgwbwukvxad5fzkWj6JkcPqsnusDQ1UxWD6MvCcZj7m3qwCQu1/NIMK0FZ
ZGS3nUhuhViaj+MnJG3+a9kG472nCS2DWmfrx99VkrUPJRgsIFmHYoBKIodR04B7
XPty14boOd+KrrIPYOr+z3Wai8twHB2+Z10sPOFJvsg1ZQbBl6mZK/UjKBMpZbkO
c5hWoYWJWbYXaUGeXGQA641ExGM2cEJkUbny1eihZbhqI4ouXfxYLx3iKj36/Z8C
0o6jMfjNFUw0TIa6OiWMqQgDdy3KE0yfZFsppaqVcCtYBcT2QQd/Joo5/IP81Rq/
iqUkZpL+WlQT2z1RAAxjG/1uGXxIM4NRur0aJxETa6ZKCRPtPQFKyzwcxDhB3RfY
hXFwl5WOaw9eXP59Q58DDlB3s9XxrqveBdoQOCMzTfYoP6dPTuvlQMujLRHTX2jw
pRXaZ1wgcXP/5FD7GDOoLTwMaodPP97AbkRSxBHlqdGJHYlATZc1GT5yktr2BsyG
xWHTtA9OjxmZZJWvmDZZwLJIzmWFOP9/UszmfAL7gOphviV3Oa/DE0nVE9aYHeTI
9j70juCXMFNVY5RYzjZPwzJaLyLOhbrAhhAZ153hp0znV9Q996W30I8fdsoaQ1Qm
jUgnLq+5aKpgTinn/qsAoda1dHto8Li3NAl2LCTQKeZA0clsf84gSpKgc8ktH3kx
jDMOQHrFB/1FpPaPe/zr6q/ttDV4lFelUsVgE0GUA0nkU9QQVsFCikSy9s8ITnTJ
MDEifye5pNk99rDIv57Imm4WlITZgbJKS1qXH9M/UYbCEzHYtQXnS2/XQN5b6+W8
2qL45yKkpbB+mMqIUNmDW2SKcsn8HmVgzs2pdKOZqbBXmAQ8+DmIx8ZWKykhEyA4
yfBf9hbqrxZIN4Xt0qFUO01fgxC2Lde9EX/Jeu4hDFapOeibv6m9/EywiYyIFmz8
GVuW7wd4KrgljGQR6mFzHKYyjXIhwUYWam6IWWEUpjLc8aMRslCZ6dx5kdHJopO9
A2q3rFRFz4Nd3buF2gpmxhsXnCor8ty48hZTsvmr4eJYanZN1wg2ayLiwEi07zPg
7yGgFdSH4Dll+9hK/HAqSCyZsgBFSen3PexjIqzRQks4udQ/lJM66YaGHk51IPaU
ChfmNxmZdgh00hoqypmTPp4Leg2GvmelO1RtJw1XtK/rBrhTh4kQ1QQTRJ16xRrU
5RSecSMLqtHuZdOLaqnSgspow44Kd07JbqYJMRLg6wUkDTi/Hv1/yOOzIEDeeQzL
eL5JINxJ6osU27RSudiFfKlLBrgopjXZ3kBeejeZN1JWkvGfpufsNedWZ79i24aS
R/xcR/PzuJht4n0RhUa8/4UBd6SLWz+c4g7c9A8kEA9BluUQPB9EVBLTYR2X2AOj
0aZDzya7qGvuLgzg6kdzlpkJLuHtjJMDiNnAbI2YDYZZtKjF5QJWwgdkAMGnCP1N
BVl758h94ulymr2zhE+qA+C1SoxYGMjUp/TsSPhqJHo96AA1qo41FMPRTNfPA7v9
D1RTGn2ZnvFW9Qg1jNVO58zd089gFakUzVlfhw3qw49pmTkFSL9oGN8wvC4zpQwU
9di08UfLIU3kZDxMhKRKMcGjmuNy6x/4GghqcG9cjQ5wICMXqxvPDR00/u6X1fd5
kibee9MNMVuEemHLuAjy/TjY6CtotELJ8UjAoALfDytISLso+L/n1PC6XpDDYFUE
Ygt2mKCl4Q6gxfN4GoGln3X4m8zXKbvyQhi+hF5L560tZr/udC4QzO/QZ/gyszIK
iAgKxySt+XunxGUlSft5RAIN30atYd9SrMmgMdDrmhdLNOkZQ7TlazGyv14m+kVy
RB3lIYN340C74gZtZSYMvAW5WuM34+gnxPWVy3kh5rAzKZo9dnkhchcHmL9GvvM3
ee5ma4/FAX+sy2e3kyqqTt4y1wIZr4Cz0GIgA4f5plYeYw7nniEj38jXKfJw23DS
hosqy8W1MciyRTsJBRTnb2RZ18zcIQVYBapQ9lkyAA6OUeG1q/lNyZOb5vGUAMOr
vD+HqHAHtynBLTgRb7IrXr1cFNrLhD3EKioaLRR1lRdtalTaVLH94HlDNNTbJTdX
MNyTOjolJWNIqVMUbLXGlZsP7LF5UQE2HL8zVZCTrM9Txx8jZw+WU1ZVY2k1Xqph
ECVVquKYk0cGJr+crrk8cV7mkIuiKfmpBdqsNP3z+CoQLP6bCN/cL8upvkF18WOv
6V+xbvzeu02a03biP7/esxwuC4XJr+W8JKVy/98jnl1P/0F4v+9Or9wN4tu/D8+f
liOXoPBBbX6LMB1TQjDRSWY5ESq6OB59pLlJ4HO7962ls8SlLvzi4eBh+yVuOhb6
rIDLaeGi4syFp8ddl8DWYETFpSBVaP5QNdrdp2Vt9G+vJVVD4csk+kzKlizL1XPN
bt7f8045STC8KiBUwBi7cggwTIaFBIZP/2PQTSWO/wKBj9cg2eaEX+ohX3zQbNyO
g9niJdYzn60VSoH8xiKI1EEtpoBdDJk1Cz26hl3URtOD5i91OrMfz+wHLBgUNUYb
HjcSALe2j8IWnPDwBF6LsKB1/UGpneJCEEYq117tR3k/Ekr9O8DM2ZVY4xW+hz3r
Kvf9kc2jK1EU3dKztN+LE0TwhQh4bX7N0LqWyYW2LA66KLCd/Yr0WKOAEvo/8CwY
pA7vweIc3X+M8zPTCGKy5HwPDSs8PKttACbpc+1IqeQrDTDHz3VO2kdlrNYkcVay
x9Nv1uyFS9zACSXa7NHP+FqfcF7ko0HXI+UiHpOQL2Qx03VED4xaMjA53IZNpIUj
Wq7sHgP5F0+IMWBLZ4vmGx+iSwG5Y4TDuWgRlB7fm812TTEN7K7XrA0G4a1YekxS
HJkybd6Hi3YwvGhIGZEX1ZC0zIkRH/PrsTjOXGX0AcjnnCA3LwL7tGHSIb7A66QC
5S9eKUnDRi9fMR9FCjNeJUTgLycANumAKxMyngeQ4BANkNvgp/SFeITXTUQVXsrG
dGCF0bnYBG/MFpVMwZ4/KaM+207BKOqG2q+QPuPklkBDLT079LQ2g6xDT640Oi5o
RPRAtYlQgNf2q+1kg04ez+zHwMzXLqlfGIE29elHJO5LhzOzsZu1jvD7poBW60Vk
KzFZZ66o7vhKE3IjqDTlAq0RjsOrx2AlVEJBuPtu5gK14V/40pQttN6nvo/Riw5E
b2+4tXKlAK2Y4M0siy6WOxTFyj1mcM1Z04A3VcagPw1sf9qFiq5cd9BBDKWaiJRx
kVPihimAfgeTCGgLom5NbZovQ1Ltsu2wA/WHWWRTkZm/AK/LMlEko5XBJ2R8fs2T
WvW3tzMkL12D0dmQ3V3oTcr8W5dXjFM5cHP0YOGn01vVnFuooGwoMnDndSj0Sliw
EZlAkdcbWZ+Q3sEn4wXNBScx6lQ+SCEP2aQOUfZ8JiW40XR+36wD3w+uR2xi/Cl7
jlfgPPnbnZYVRG1LYtOGT2KFFgvCPk8G8zoyGflseoJ5ipub6kTtC3AfY6dRYnc6
+nbtvQFibVsoUqL3M7r4bzH6o8wzsfphblSoAQ3jIcKzCpUdHucsQZr6oDa+PkTG
yn+0EqVUp9CzJFdfiJ2SF2iV15yS92wTZPtUhL7y+I18OMMNOsx1JLVs9Zi1WzYk
GA0NN/MuDA0Dna0ssZoYIkxLa2dF41fnt4xKQYbVy0Zi03Tomr1hTFWaqR1yrihV
6nrrUn2OQRttiUrdtl1uHh+bPZhtHpnS3tbCAfI8oy6ic9kUUI9rtZGfTKH48FWJ
3S/Z8azZ4+QnsjcCnsVZ6YhkhT6uzOAzTBzA7NYbSdkNynZFiMOwqxlzkBIKov+I
JL3MO52rm7E6qTrG13OlJ3V/ENVfDCecsRaF47gMpvYTHxvJptOKfqMynbrN2JAN
1BhZ5odioSjnNbN9P7JVgOw4YZV76gkdkqjUblMZ+rIBKHg35yGrQMVY7f4+QFa9
XSVpxA4QwEMv4Prf5UOV4z5Bw4qZ55jdjBov6E84OVTEWKh091rJkqrKY7IQK3Qx
Xl3SHajZ7t1MQOYMTMGqJhmftZipxhcOGXO2NCzZQsVs2T4MYcstfy7SbNe51Q0f
5sY+VeA2cVkIhwdLAAK9yHBM+UkGS2X1Q5/Ar0kxVr3iYhvyZUAUx6TfdSyZWTXF
pM4zOFyQqM+Skc3SnMYLz3malK7IO8XJREfDjSTM65QZKvZbVjc977Dm1Mp1+25g
q9MWFkh1HnHVoyIvlZ3o4NLdLbxU+x9pq/n4nnpMmMFarBVD26u9JlnfVBsLyVST
0HzUbyI22x/Dmumpjna/Q5XyF/8g+IlohAyljjSAcJFR3PxPx5+2a5UgL1HSjGUo
4U02yLlmOtOBZ859z9oqinGSJPf8ijbP4nV9UP6zD3UgCHtOmPPFphASNt0egJ5g
goE1eDS5I0rM/M4D67IGvfcgdSvWhL8Q38fd4nYtULluJYRfeGUFT7xoi7o6XIlc
rYi/eJ61PYICLNWAOja1glK/WIPRjBQaKF51siYmBmpyeMczPMTvqUn8Q2lXUCKp
1bvNtAhNpJYCON9ZzkeeaB7x0Y3t1KB7JUYwqALxDj+CHeL6TuRIyOVFH9HEaAjd
5tWtd0eUkeNbRLmEkgHmwrrUTSt0npSLOg93TUH8+nbrcFxFynprZ1aiFiT9qRS/
nsUQjrnHFUFUP7VPEQKsfxQK2Qftq/DJ4Ism6vqo2jrCKWFJdVXbrETZWePnCDwT
QO8T4pDDa4SjXYXH0sWNgFFRp7dZIh9tXM42B3/1UKw611a2ewKKw/LRX1Z91L6y
HHjrpQZc+vzOQKom6/FXzNFyLxP04VwOlVfA0CPuEbhnml5ZMJY7ceGNzvoyq6jx
CNZQA+/3Q5ADlEa0McGBIFqAtogkFChE6Gtw3UlqLIK895gnfHJv1ZrgJEB8ArV4
H+Q6+QaQFLF/klXWCOYi8plpr7RWf+AbJwsP3xlTETDn9loJ5xvRu9vAV4n7mnnZ
xeZ/JpF0M8YHm/Le70nxAcGeqbyP4MfYcdBvlgErOLnYHfx0ArOH5ttOx0V7qtG6
L3SmUZmi/6BrP6gb6JmWLsj0wkY0+VEBF+Y2XiufiPoDP9Q7hcIy/ZgZ3jEmvMqT
v0ouNG7/1nfr3qKTSTfAnGWCCzJ9Xei/OnGmm2aUsgJvR5i3i1hTpCeMybKODQhG
iN25HAUn7xmblC/VZ4zRDnv8q0fLcITzJ5baOJEDw6Q/z5kkMN+fyPlfJ1RrRBs/
lw8/FghKhgwDDwQDsTBL6g/wLkB6eltSl+AufyP2JPU8/89r+psHl00AnvvcIpXh
xWFsNRWjZ6/YCMk2nl/lv0P2Y7cRvkDBun2DFbDIR1x/DYME486iamqmfJVaYbPB
XTqOnclmiyV1sNAgRyOzfVpxCdIiVg6kL84rHYtsJLUy4X7SbTUDkVUGeeo92p7V
fuz4i3h96QB8MraUVE53NWIZdEeUy6ACsyYZ+vHF7gkSDopTl3pHKKhl/Ef57kG1
Tt1WPvDR6oO7xNYneTvBZZPvVboH+NytPj56670WeQ2AVZRKp2Sq93qUTaVzPpMo
vEjb5Zcg2Rvz8jNaPlTtlw==
`pragma protect end_protected
