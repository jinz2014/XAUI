// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JWXf56CjpKWkoZKY6L0EIaDB3kc0a4J0S0z6pkxZOWT8zGL6Sc3rPz/WePvHdU32
VpUTwE+Qu6tPFwkBNUd2FqPYdIirb7dHPligRkqcXFoF6Cc2ooXQhDOnCiErO7N9
pHXCyHeJupTxqPdcdjcA0UBeCn07XcwhevsgSyeSY5w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12208)
n2/XFaM4j4UATCwOMQ3Acj55+HCYPapYzWIc2vvbqQYVdJifwv9jDrTgUTVUnH2l
MGyI9HwbsnzhxYO+mKmlobtHoPgcEasvRR+udOa6EF684QiZ01aELTh88sx1E+rJ
HM/xdZZ+Qi1QObGRBm+AMlyHzeZQ5613EjsehRFiDT3EYjqdv58SIULys5SylkgB
njTZiQI8g+4uy178I+H7Tm6C2cx3lvCYAFEV+YkDmBvQFIOw7kQ6syINQdUPsoc8
IDD2vtGZ3SvK21OvbT5TYmprsVODqXqyam5+Gu9NDw5SCy7Pt8poP71+sd8WRaE9
8K02UyJbtOrnAXiu6+BB+lR0v+Tgz3XDgZDH9K3Oe6gw/Gzbe8RvZpauBgE/LlMW
aCJ6emExzUGQJq9ZXKz7JbRO+FaZnf3235LvKylV2pUy8k4gOKXUoQBQt9alrZVb
s2qhaSM/l8+sfXOisjRgAy2XVHfQIJwiEEtdB3D5+4lviFCVwe/7fQU2MQsckttN
NwQBMkykQpuDNFYiu7/Jmv1Wb5AlUJMCn4M0QRzmQjJo+zjFCNQpmDbcWrtVyKPD
KQZjfyI9ei7yXcH5tgj/1+wAHTBDb0PE47EH74tC7YBMeqd4hcKxxUz6uRgv4kj6
vLdubp/Uwm09bQnYRHpZ/phXE9aVzz7SntYDS8pYnSpibLZhJ1xwn9Lihiop/6zc
zIQ+8etjYvxiRFpZwEvCcV5/3wJtRwgfZ3/uX4LatCoLivJbb0niH6DRCVOY9i0t
ef7exu7G/2Ua5CPUpgT0QQXA6t0sd2KoAF+snrWBpSBpJHkVAqtjc7yzrPyzu2OU
Bdpy3lUoU8FFrrK2TVH1KmO+1NIIzLGR1dQHQYI4FZ5QunzjtYbXGoeGE7jlWKC8
l2nkQzXV5HVxMDii6N67+u9ScNnUjlC2Ki2Wis/h+p4VGDwm8irUgddlhLJFbT2E
6QJ6UHIbTy4VP4pvLyjZeCpaeGQzOOhEv8rxLonii7t4k/T7LGAwzQv96c2WfA+f
4aYAnNKn1U+uHRSDC/4J4UqOGSRCqRV8pGp1xG1kjPFE1fFdNBIfg6yf9qClqMDH
DdPGc79xBHSxni7AVbW3PE/iWowDqUZd1BB4teU82/Cjr3b+VKT98ZjtoSrS+8Z9
OrUhY0To/q9oYTNo5BFTFnLyw2uDp+QAQywOm8IKD1SB3o+XGit+54ZaDuDb+ZN3
s1zom+ShCOOU0WPovOSa5GyUPilntgayQJX71ltd0laGNAdSw5LpwFwtmrU1PXwB
fXPsd2Ct2swPwRvVg8mL924f3XpdJidi4/ADBk1eUXeAF+ncfLZCtwKVEYnLzDX5
YUGJIdIjLWnIi3QFZ+xznaNPSEdVmrLXMh2S5ummf7BLkPyVMH23Ol7G1Sp1gDDa
Wm0nuax/QbTxy1Nx3LlCgBVsM/UEvr8zSZJAahPkRUBFealWQd6yvt31utJzcPPU
dg9ovC+tlNmmJxn2m80hOlFoa9BnE97S1wTA33fjehsums1/HIxmu1q3v8O2ULip
qiF1Dc+y5I1epGbcEqfp/EMoMMjR/k5XDBoZOYVf90vnF12mDuJP/+UijC6VTahh
lssBZu0/RFP1ZTaQUCHJBd/kGGITr/qzDjgGNJEOQehciYlp3ZO4hNHc8/tvw40F
fygkMP3ZbWrPOgDhYCEW1J+k6AGvGYtJx+2DPaVAqyK3qJuBHAXWKRk97glP1iTp
f1dNwQitpCwGMa7oydUMWTts8/VqkdfMPrjDpQm3sTe1XlkQ/bFuIV8fZD161dON
kDJkvzs0MJNXa+RYK2O4Mtrouhf8sP5XmPU0uOzXloC8eUYM7gdSNivr/hk5ppAM
YHCjIljlxOQtdUlgvYwSuSFXRfzQQRQKRkgGKXD+4Y71FOuIyLBeKf2NZgHVsIOu
Ow3FOEiD0r7X2Dqq92DyyjhiXZaduIKj7aUU+sHz+/5lf7CQM3sLmO/4Zkl6Cg87
YimT6BHcYNiGNLiaxUwlOp8zwqyVedKBUKp1FQkj3eKfTnANYEh+A+Z72A42iive
Le5EsaaUHSXkjARYLF2GgwAO/t2H0M2Ul+Rsiz86Y3JC3Gj1NPAl0TxQ2v/hxDBg
4hwCvtmOaTXohBV1+uTtUCV3JnRsWReOv+WPp+8qSJI3ov/c3k+BiW9/H7PfqD89
4wkt0nMUtVkzCt/2KJfZzJUjNLOLnFipnN/KzSRfNBWA1BBOFqyv3dEJqUSDPviI
1a+k3MB/kmrHtx+ROt8LMpnZ/iU69QWqycpfubpUq5dJO+kLDFol08Jh8JznPekB
gGPWXIHw19x5LrO6JN7YSn+VIIG//fjsl1Co8y9f8g8YaLmX65GTi5twhoX3XZ/E
Px+MNerEsq33fs0QTNkl+XQ8QTc+/C05zZprIbVwALM3j2UOxW4iLrOpd1izgZsf
tP4CAXNq9G1G0C66QUvwjK6oI+yOv2o+O4D4mTVJEeaJ8HxcJpTGkaefGqjuGbW/
HE8SSAJLtbJjoSKSnC58VsGO9A3UoAN7lyEPTiCRSpUnMnu55O6D28Wqv3N5BYX3
KekcJCn2MstaRnJDhws4KWK9z3XUWpWCHdZUCtdj/bx6Z+t6UZ5zVAUbTj3yJ1iW
+vLNjZTzjNpniIjLvWbXejlFaHNuD6xP1bMpQJ4ImNLOGeXFrDClNRzNhW6Slp0L
X0kU3ld0U14fGhZ/Ly8DSd+jtYQPn77HYD0honisLG+xvBwd90nWSwdvc5z/ARWn
nLL+yd2wWvrRZjDQ1y6PW+Ubuyy1K9gGdxlcLF2ODzWsqTb4QTVZrSn1G2gYH1yd
NFn4YZvmlG9DlP8YYWTm1ruAjIEBxtVPRL6rERxa7SPQXZphJ6U49L9dpCcp+gC8
4eb9bcsomcnqPuomo0XI3PHAY7hBM+7+srGgc4iLViFhTfUMajgl/X20hKJzwBOl
hxqwEvTRgAskaXS9o0Fl4F/R05/S2VwJ0TLJtZIyU4G37g9hFH0utNoONGhEzhLC
mGtk1UXwh3spL8PO4mUzL9VUhybz+bQDvmog2pnOl6SDo3vI4dla+TKkXawugkJD
NtHDaYk0ixemEkpM1ba56Jnqlowie9muG8n8BFa6AqhKzZ8sU9RP50e02jyEOOCK
2mUDqqVjN9zWkj495MfGdypR2ktitSn9I5tRQn1aUxGHG0JmOiS8VucgqEAJyl0E
HnLikX23yonhvFF5EPZvJjpis9TYPACklY99muhjGi0kn0o98SwirtmQnq0CcxcD
gPDff+XBkKOafIHjNY4EsMSoV7kuRLde5W2IkXjPZjkvold6spjYm0iwo526btZ3
6ddn36RtBqtFiMiblb4+u8ViyNMGcBcS2PgHdItQ9a6PQF1KPhAgaAtAXyn4ptH+
aE8ChL5TrOULXxrUTk1u+nNNq2MkUi2KSUbD+N/WLgWps6gBsGEilKG/W6NB96iY
KKd0rbk4OItYLt3tFW4Gp5S8JTKQNuFT3vGmpuiUnZnKcmF5qHakP1NKGscf4C/L
CLkWM+O44TCPnOh8wT4CLvOuvhvzQgeQ6UHUN0XGS9asLxeA9L3B6tTrhhRd0YWA
5WELuc4naR9k1eM7IdtV8LLDPdEtW+YQQC611KoBryRzdleLskbCfjv2UgesIdgz
ybVMa42kOVVN7QtbU1LwCIGP/prbyVzDqiVxJkIYT4Z6jLx1HbNqNcd0M42H7+SC
z0+4hi1//nOVuzaKOpeDQsyV6mOpEBUmW9r5SrbeKzVNHnY9/szgTHMUiFC2M4G4
hcbqrZExr24AK57EJbxM+MFpoOYR7mJOfswT5S4Cly12+ZljeSsdEBXd3FxSQOg5
I35VSxd0I6O+s2ctAsqz6uPqNtRkxYmo47TRFPpzRam4jbAETKGhLa0wva6vO3BQ
84FjcZIbZVSmu3gJzbgyhnQs2AYa5fXW2/m4jRTWBSWLRNK8yN13Z+43gHt0gyF0
F5hvftpbC17Cg0mQowNh8QImyik8f3GqwudBRRyU6Fm9GcFgDlZNQRt9DcyZX01m
RZSBo7eKEsq2wdwf83a0nrXJRP+PjPI8HJef06OCz5Sz5FMDFWO2SIx0ZkP5Xp3K
kmx2R4TodeM28mEsJDs1TxxpUPcYruvop3mRuN8JdYjt6PUKl8EzliSZulr6nlU4
zYDwdjBg0JTaf9nD5MNMloLAcqBta46uDe2e3hliBzwF2+W4+evi2TNFV6WHfuVH
7JcuDbN4utck24GRkcbOixfgxGFlY4qGcbN38cxqfCeF7Z8wwPcX+ZUpIclZNxai
rXaDJZAELAzRepvCkPRi1PDLTIiKJ+vH15aGAhzw1eoEhAWQurHUsBmA/Liwnkcl
ad4ys+P2BCmyyhu/XjB6aqYcK4ZME6rS5tnsBHh0zMdQt8czZld/VLkFQxJBNBNS
5la9/4Pw5e12kAmAOzKY9C8g+oeXfhl2N0hv8fXr2+yoTVbdH4httGTJ208bJitc
dm0igPdEhgzlXYMS9Y4rZgYDSJl1mFcruEL8sXcNqQxofK8AHYMd/H1fDVg/4zD1
IZIUNPFSKWCT2+jF3/OL2YA8GYdLBvtsqgmjJHXOnxBFfmxxvWhEZ6XMDumnpRP6
sW9oZB7dfQOTHneK/mwTQA3w28jQwWGRJ73iI4rQD1ELSzjOBO9cJdOGcuveTW0L
Seq6zTXsaPuzKiybeymXQJC7g+rJx+vkuUYIZ1DYrrirSropD9klTS+Wmzb5N18a
x+MUiEprcGhULzWdEELlfjd//zV/PuivxgLt71S2cO5g3IhB4TEv1B7dX9XcjiwU
u+5jWlFuLxVPf+frxYlJWIgj4KPflUOQ8pExl72l3Im32lwlkkIHG01fWGeLg9r8
AStL/RwaPUssz5XQq3+tedYKwFyr6gob8AGB07Bjl1uvHeNmdADQOuv1cHlhXH2O
blEO53TFWjgHuQBBS0PcFPKhM8EZ0VhRFYQBder0L+GjHwHBbvMTJHnfG/mXft2m
LgD8Hq2zxcwmW4Q2RgR87oEidng22UhANScRTWXB27sM1o3HWh+Z1Aah3zJk1kGA
uzPhp+aOWCrP8cO3E2twTeKlKlT/tbHUt1i8V7xtHPSES72z+YHwTWSi8JvT9Y/v
l8psyPTqcbhTtBFtuZUCRe7PW7fH6YVEWRFGWJ+T9El91DGyhVSf+ZLM+fKu//xi
V4ICIIlLuZrqsXaQF/u93MscNOvKauvUibE5jz3sozXvspvgqdWE1K3jOH3Edg4B
rqehsTViGdyW/+2vbyvLj/thT3OR+3nlcKN+4xtFVyfewCUjhmv4Ck8Fja3SNifX
Ypvl/1VssdDchww3uY1xKQmxLQERQvUfuTwmduDrP1jqfWCi20O3iPSK6VyUOoiI
X9SehrcpGU3x2BOLRDZeZ8tMD0nhACKjT/+axbc1bnLIu8zmIkkZiLDLNWnG8uev
kUvVs5bm0vUtK+pxkvHyR9BFOwWMd13m2KXV3iy1VtTmGKQcfJBAropddFKqB9ML
8RtLuLSIH6nSEPMBH+7PsSVJjbZhEkT1W/TD1QApxSIWYyaHmnmDEyq1BA5pVCR+
Ho7YwsjItoT0v/OPBSaV90Tm2TfEjENi+XS3MyLuvW2ytIDNk/CY3tAWOu8mOnlS
e9dN1Ql++CaDH6a6P61edW9XikV/dvJRelmkpjppBc+M27XAGJiGUeQ0G45ckp3V
B4R4nZbr5fKZ5mAOT+naywkwejXIu6U1pAVTnyfvxErdwj3mRPNi3beQiuMLORCZ
NaqoCliwt9i2UhtJiILfGm3eN8DG2C1x5mYoMgWB/RBuFSyTY/02M6ymhedGq1sI
TCMJfJu2dPXLAKH7jZz9EcWvVNWLbHzx9CFGkpI3d4PCj3150om4An/JAY3u++y1
8fXGwsa2Yytv+bo8sO1hl8rQKnRyQv6x6F9jZfrRDbX5SZhgY4w+JPUOU8tlItRA
BYlG84XgvnfzxvXelv47kRN+5Elh/6PhxgqW2BcLf6fJ1zHQacSoHLzwWKzf+297
E8ELY2Elu/ivqPal1RahY90wPNunx23qerDEc9mn8v7a4/51T++EPzXrXueYyFK5
HgDCX3hzHAHNE3v2jiq7myg3wsbT/34FG15B+XHst5l2PB5zT2c5bLF5qlqEt98n
YGeJm7nTXkcbHnIjhmeCUo+KwmdLTw51pAHAHGtOogOftADZx7W7fsG/SHEuBFsG
9IcYjT3LIvRwLl8OcFxaL3aUUppLLj/jTJpXDn6rm4+Cnbr8yYjkO34UmqWLgyQ1
t0YznROh+ojm5bkp/qn7+hFdgK1/fd4TuEw2BW2UISGM0D5bZr4VZHNTcoa/J//B
PdwhKI+/L6bFzyY+fX4rdutH1WjMHnBKnqk6LZ2cZ4rPc7jizt4Gyqh6YWSmQxtK
FadQpxTA7D4HiIBvsrnqqp3TR0pqaqCWWIuDzIdZnuamzSKe8L1GCjcEhFYiIqFi
ToV3uKW8urStZh/NLYcXMPTWL7tc4EOJQVS9k+zpfrNSaPc5kUSKFVci1P4P79BW
yvnh/3qvCiO5e0/+B2QJTVpsSEkTZ4eU8ygD+uahuD62vI+swNHI3/kQQOiWGPfS
73mgfb1Ds+5WKT3mWqZjmYYefLjMkmHP87RTxZEftKNgiOAfZ+nJPMXpiGZdIWpw
S/eFZ/DajgL42dOC8wsnHZ3BXlgj0PDEiNNklmcx/AF6eW2RBD2pwevTARquMSVT
FIuyvKtyOD0C/1tyZj0eCsLAkTJqk9iLbjNbpFzi2/AkbGhVbMmf4aGATB7j4ZoN
AwsgRudA+PwMEtQ/TM3RfxqGcYg+IKWMtjjAgoY/5Vs8TBxt6daaZhJYwz4buDi4
X70Jg4MZWY1FO4CjDEm4Xi1jHa1YIwppyP04liSxSLkncyC1HFRd2DEDXKse/5n5
qhX8uHqdhyG0Phu+/7GdbXwQthgiSb+es6bZmgo3M53UfrNcaGFMbp8jz7f26yRU
9TOCCpiZJwf/rD9Qmh1Uakhwmtf9nv77IyR/vnicgT4B6cNu/xX3PTB3iw6rwZ4c
wawPieuxPSwSr9wtasmUjnAZNRLH3ntBzBLullwoUskXwHAOp3o8VSE6RJsBkLSl
KQ6YMJh1FoC+83j0gNzVvqU9Anp2aSLVY+/+FMtLWaxzCydf4GZF5OpJzxL5hTfd
stheUwaRQAvMbVfplM9Em1BvebchOnFQ0Wu9WWdq3TxylVOSBPIGUXvrdfR0ki+P
XiXzVP5aiB0wXMo7VNLqFrRxu0uDt+6XHRS1lueVM7ajxmGR+bzC2xXAYEbTMB2n
+EQxho0aIVoXwGxhdW+Yza1DJqg1T1RI0QcGNRu4BqhJS17Ngkmwf+R4bySp/Jst
q3+i5wViUwTYC5xaFr+EmXDuuzm9Ns2cKvaItoeHDku92p0G2sOLaH+0wGRjhJcf
RgBLqpkyZXxEu2nyA9m5L53g60Do21GtBkTF2HZrQQxdRMR6v67IFttBH6KZe55n
mew7mqqR5r3zZGZfvOkWQka/QfVtn/40YjxdOhvJNuYTRCpsJHbzaFgUniPZPpyE
ijQEc1EdqwZlZ7HeaV4dI1ckTL7RIKrru5YHjUB84RCgpbR7u8XChGXBOH8jyyUB
OUdrFNIPnhCazZr8YxksjQUDG9T4bHbrKsGbFp9rSkknw834d/htqQU0CpP6geGp
dym5SRUDLY8H/mgXbQSYw3NKoMiI9jTYplxs0NB+wnMcfZP5koef/pj9dL+eEu5U
hwUuC8XRKt4XblUDkKSxx/ub4hD8KgY1JIWBwc7fdtkNkBnu8UGSuAI6kOr9bSz6
O02U0WOuTkXPmHeJMUwwwmXGHuxWjKL8ibHeHuv44OMsSmIzK3C/6BAITqPL9TT8
cS/8bsSQX5PyKZcaiWZ9SGM7KTTgJPmrbe0Mr+SrWKRe1AjvNgMJPYEbz9JUyPgg
QzasmC+vMxUfOELw7+HMka+m+u3kljdav6IMyXcCN17vLOzTwC6a/J1jH6q1MC5+
7wAc9jTohWV5Fhxkposqv4oomBTSE2Gu84/Fkw4ISePr9BblBIOn44zl8Soz4Gw3
f6pyDgGgK5+DYUtCwwImRmYJ/nBHy6eJd6pBotSbTVIrA5kWZo/SDOFUeslmvi4U
x1LzL43Es1bGBJc0/Id7GKW5U30sS0b2+GAn9xkpXO2dntMgsU9CZ+SHAIFGwFWG
o54hIz5vJlQQLEFOeo9zyOpXD+L1aciDFc9nISCsSALGt7FJEQz/HQvwVfu/bY7j
6iopUbELPXTZ6a0PuwXLp/+ehqoVWYCg+GtlWgZ/mdQYQ+lXg56tmrMCSs3gTKdW
GIGO/KdezAUhsELNMgUKDpBVfLxsInXnhqAc+amYbL2fRbH/QeJ7RS5H9A6MEXO7
U+92+bFtOK1Wq/rdyMQSExc3oWEBopMPcW3ngaOd7AUKcWkEqLbRzMVFpLGyeYNJ
8Dd3/4Hagt0yd00iOEkNDnrATVppFwvmjrBAIao3xt75YutNHuV64v7U5FK034Rl
OI6b2Msv42TKwLErYqGj0R8va/KCsjNPhsaPEJppcbDH1lXev6NL5zj8s0pPArgl
etisbcvyJyv8LvL2piu2hb6MQg7KhdiO4rip8ypu61AifINEKAddJkiZQk+yZ88S
CZGspCGg1fSB/aH4NYVuzpNzA1xuVWXQAQQgtEZLMkzG/ldq91bIWLVIxDtWXWYF
NsGfzHvu+U3v09pjXG7jtY7gx2+q8DnNnp3RTsxgn09r753o2BN1txCD9rZoPLSL
2fq8bmKAle4qb100+kvYzkm3Mb7VqoKVu8nJ4BxP8TH/ZHs+gOID9oLHR6vqSTr7
am/Hddj8m2FV/Q9rGwQ7pmOnb7enYgNUP9WePsR5sVzRBjIQw+xhwX/dLA17RcdE
HXmD3lOp5OrUk169+uAYCAYQc2IF43BSeNklOYnBkvxy8nSoHntsFhCDc8taXcLA
7YuVPgm2CzL/xeAe1I7hUbLIeawkA51DNHzRKGUTZoHz3mKrVrbIy0N2ceuCXOLU
THAq40chakXHvPAb6DMg3DknNKc+PSe3DzqPQ7yJ7PJFRWLdu5FfsJEFv7cC+sWk
LApT4aPR0b1DG4+ZjhO12izsL/HveWWPpqexwwEt+VOicAfINjZSgOww6YSMjEOO
GLzsWAWTvoIR9BR6op9G7pKkTOY3dRuwt+ceHiwPaPBqRixH9Dx39ohNbDVPqPMq
2OWyPaZJ2ejk/njGTCbBK9mfbttYVEMrhnSgP/n3+8KTq+yUbjmsvOT6KEKpsnMR
DYxeUD/lv1lfd1skHHWTjBKzSRG4LYKZg+xyTVnI9nvsEV0kYbUV3LeBqMnOuOa+
74j8DdB/l4pxwYAuFq8Snmck7FDJMFn6t9nHzLjPejV0e0/45A7wv31QoI75JHu3
cKbx9I1nMbcnCbXypj/sNddKQKVrfhYdkTJH02ZYIEZ64kAxuLvq3qR8kygyKUmS
rXwdv/7Q1RZ8HPPhZgiWwXr/hQk6gjxJCgWvwybTbuPypgfujurP5e41BaGsnGC7
7Y7mRuB8r+BFzngNdHToJgOqpgkeDNYnbT5BPgRcvS0efY2G5D7hmSsvQWm0tQ4l
5RbgIyd2k3gNCGuqB6oWYuistAPrlWsZ8ThlwyNwrrp00KxopXnZ0Jj4MOeNH2/5
mSa2/OqJOouzeuP8ra9vCIZXX1hSYpBVEq/V3uwD6WtOUCJf/N8x3pDd5jZuizLE
20+s270HdohPG5C6+XMBBtUj8/3TxZ96glyISEFBiqJokidLGgnLKnEIB3cX4hwa
3oXHNliIPKgSdzIrAD5xz+L4AgKwVftLhHVs5OUIH4f72DjSJm6zZ173OGEUEmWs
UMrGJ2Ozhy/wxe1UP6obTPza+vxiQGEl1kdqYFbGOOoKJOT2c4zas45VC6G2xzsi
rz7gZ9E8JujMEdpUucQ5g1ImpXBqOUA2H6z7Q543scG2Wj7OjVBgzVWwNhx0JG7A
/Q3Zl5xsNRlY0GtFiV38uWN6DssEXImzZgr1x9DI/hjpM3UT8lXXpIJ2jd1TBSVL
IEPKhmiO60ruZOJmNv4dWJOae3MkpU5MWzQ1FVz44Z9UdbalX8yiwy3VlVu4jXqH
bFaREb2QoNhgteAiWCdpiivhlHRzbA7wLpvOZVssi7pXNkHj1qw+IU/3EHOXTmDm
AWxjANjcDBRPYamkxNasLsZ0RvxqfIB6Y2H1r2BHA/vuQycZSYD5G//JQwIPecfm
VfIJ3kDUJZk537h3BYN43Y+/4oHRt8zvVf9dU7GN4ltmYd+M50T3VkZpE6VdvlhA
EHTYAQJYREW+10TQJj1XRz5bT6TnXgC5zpVLp0SZ3XP3ZcmCFwDNWld2sMdAnb2A
7jlZ/33FLh25IuI8O8/KP366aUrSNdc9RKjUzXLWco03S0xAeGuUb0zORZREwpLS
RhH49Kb0F7OAkqZFJF/1WTrUc0GG5DDo6oY0psyjRqpPvq2xYbVOIzN6TCeiovsW
HxSCV/ha8lEjYG7aZ/FoJ104uwEblRYRTtBUkpyxPz48YyqMOoK7gg4ZjCADBE1b
1fzXBiY6Ee8532gDxkDJuoB+U5s56IQDmFM9KKjfgTgLMELU4f1XUzfWl40k2XrQ
gO+GRu68Zb6F6Z/FssILACkB9dLAMdCUK8+VKpU8n6R2VkCv1D4Jt7x3rnwmhQ+A
JFEe6GSz7cwkRdF/83MdHI2rgBbJ0Hs9D7V7F9Y3u+zjCJVM5/efPuGeM3+eSiYq
BuPCI/ALr0LJdehQsaGKfrZHpPTJXdOxOyXo5QLnNVRy5JeLXuf52zkyAq2KkTLM
rLuZIDRsBx2CFvPpeKxlt58GQtYRdKKZmGUBRJDcTVVlnAjn2HxuI2bZ4H2/ZZmZ
glDfxVlg66UA3CMIo7o6TBNXzC346kIVmhpj1qP2EAsJAZ3grfD/uGqREJzTwCjd
bMi2vovviD+NxWY+kZWE15jzsUtNgo5mK2XrWb7LERRiz44/9ckrOTwJuAapDCsP
UlzpZ0cUFar8nvboYnrdwi4nQgpRO0cr7V03eS9VpRhWH38qmjNWL/Y3woH3k+Y9
n351nv2zBnanEaEgw0iwV8qlyC0iYBKr6A4Ok/0ytgRe1GChZTwcUcvLIygOZ7C7
dkdaKtfjpmpYZX5FqlXKwkDrqDLT/K5XGy+IosO5xaj7wxIZcPYA97e+07wCuR2V
ngUdWKu2jMOda0pfP3yJNeLcqxN6bxtl9hllg0ldA3bAmpfKfbuMr18TNr+mORRr
kjnfXlbSynohFdZecI/5LypR9lDKsfuANeku7dplmgY30aiZaEKJ7Akeqsm02fsA
s2ebBpmtV2kfyORZDfY3b7y/i9SjXrD73QGHgytv3xkzjHuk0omaOlN8CdpFP2bG
V34gODL4kV/+/1T2kx713t9QqI2fPpmynDRV+uwwOJqld+hLFQQ7HEjiCK3HX4XS
8+7OONK8ywVrpTZHz5ZGgTyyxjyWLkdGn5zKtfr2oYNaaPjJJcctGr6HFTcxem8B
3+JnuogUbLskhIDMVuzriPKCIJ9qVdYxZLncKmjPttBb0cTgTipkhtjcJiAiKTF+
222V1TvQvpqyXpI1CxHMivOKAbV+LSfhaMzmnh+9eTdAy1fdR698x4lTgNsSyhd0
uJ4F6b+EX/Jz8tEfohs2oC7vlqqnjgXhM5AYJ/QXAi1fLwFHy/ZgJO6VddbhIYbM
cuPIg1tWPfg4LmHMVZYo5/Yf6hpzleOBuyL/IDe1C2TQ7aZ1TmQ1vFH7GIWJOVhk
YIVrdzjQqbB8Ua9yErGocjJtvl/0Jr/i+BoqW68fUkuaBmjX0VSPhoImDlscxUvq
KLgnLQjt/4736jOmvXoWaE2TH3A2u0fh7UneeACF8io2fejDQpFzl9vLlURw+iXa
yBKCQw91mhvNt4lNbjy5lbF8n8AMMuQGjPvIvY8tP1ROYlozSv4a8eK/VQyTB1SB
cKrSFPlYXb0HsJRikBlVz9g7Xd2UH3M426DXSmLPKXhJU2UDFC3MGiIBvzDp+tdy
cqQIdeM7OrL3M8Nbmkt2Knp8tPbC4esBrP6bR6jD/uIDBnAJXptv/K60nJPDqzGV
9TRY60YRgpa2XzhNpc2znBF2zp09yoI+0iWPmoCkKPkcgaWl42MDxkvk+joJun7o
eXWPrG1D/PatV8Ior5ITtx5wVrTXxdgqows+Y0kdb1II2kjL9Il1sV+NciBKR5If
FBgZ5Zgh8Ufs/+sfF4Ye+6tFyYZ+iIuh3v8PoAm3KyzR8+OHKkaUiH6OUjWvMVWu
97HYk/2GyVWOs3PPfNUNstrwXFcZfzVo8mxL+GaZAojZdSoI2oXcR+FS2Rusu8w/
ZMp6o9Q1qGifQvG6EjWBVNidi54NbyFVYrJ23aFswSMcHVVAns1sPLZYK5++BBD1
Uth8+vp5Hc8Q0sZOVP89ggw7/9fw895HGizIbKqP9wU43PDrrzgaLWTt5pQ+4kcw
MLvXG2me+cL5Dng7nVztr5F8KRVPIWs4DeCJ91xIQa3Xr5yRtdqCLjJ4s8/hjfMK
S9ZoWQHNdq4In9eooiaWC0X/cxae919aGl6NWCNoNUA1ItgncvAEY9fa0bcrwc4H
hxlKuZvOFLuCnRc2bQGNwWvh9LwN4oVhbKEJ19soD89fk7WeAQUk1aYJnu35ZYuG
2iphWdimgiX32eELaG9b8QKcj6SCzwJmth5FT196Xnsu84lp50F9rsKb9kkfz7J3
xHTuVxCXXp88Z0shgKY4CvMLJZEGOlrfRdez+mRTiNoqLkt3t+ZdHyqu9NoCvlt2
I7jfQqNNeeMrGUrsZbTWPQ0QTEgWXP7FU89rZ+aGvKHhegPVhqo7z/43uWVDUoyc
e+E2+AOF7u+HK731F6recdQruujBqYiASdKHTv21Suwk7034dqOKZxFEYeBm2Jz3
PzlQI1388qx8o5s2lmQ+fXGySmAwamiOR10qsnpP2BqOi/JOs5yJp5MfTyim4v7+
fPOKbZEJPFGzLNetrLqD3+bI6IoRoNkKmFId0kOh+V8tTkb1O/t7dKhq4J3YKrOL
qBgLm6VD3egHdgRmj9uwfFScUKRAOjYNf3xbwAY6AWnIJEBliZNP/KQroluRZJt4
qFPEncLrCfVQY+3pvhukbpdRk7Cwd+io5awm4RQ3odqBzTGyVfCN3NNGP4FC9gxZ
t9y8j2WtzJWg3vJg+ELx2JEvDGh9JBiFmIFTvFuBFJpDLx2oDgW9t8CDkO6L1BjM
2NQCUulCXypDr+FSul7MXzaSTGuctMTvlH2VKiKsBlsU5Hb7shgAp0sFrOgCnJft
owWxuR3kJk7794bK/K7FJDC7M4x1Wk7vOvBKueL1cHzjJhEn5pLHyh3XQDVmiQOL
vZ1y++i/Ii8qWADl8b8A8CAcyEHbrR3a6gQaxvYnjb8dFUu80lJQbZ88YqUPd6uM
QSDqSlwUmrCXbwA/veT/EdnpB6ZQhYOCI/UNGI4Rs8MNxxsLpSqZYrFtIz3PTAYE
6iF2L+jo74+52XVOTXBhDkACuBXfFY3aeKc/tQCAxIlfKHrtiG6XQqooK8lpY4q0
BIg9ioBRfzOaDx7gJqKmpKJ6SLl62rK2tpSvNBdEva2VXbKs6KFNTN3HEPF6xY/h
DZUM9O/u8ROsjrtxHv/o+SFgVmWtAe2KJMiKYvM5vU/QzQI+a4vgrTm6A//VTRAx
EMnyRqgOn0qTnAoDeYt/zrATVSu2wYG+sgzlQS6Pl4rODXPxJ6N1tLvYGKCgWR9y
Fli52cRlFaH4knbC0eEpLL12NCRwz1J9iLTX0CchTCc2DzimRSmmlp1rdA4cV1IW
XiY5og6QF/lrv+/IUdCRVReEyGeE2164pdFDhBm7HBKXU+3+MSlPWzIbsDNjEUtR
iYQs6xIEInuCVPsXqknflhZC+jhQSqmJP5duemcHNsYPQpczIcFWXDmuXJrEoSmr
DoUM7ypGlZu20IlPAvMbah+FlN7yDypvdgb4upkEbHljc8BEgaRmNcb3hkE5fqRt
rJGCdkPtcTehKLHg0xiQrRMEwJHghvLVuiZzZjFjwaYHI52Xsaj1dNzHALyT88t2
q7eL6oKdcxryJ3bDirT0Xkzkbes5CM2JHtqwERMjMr3hDMUjQOZNV/77UghSruqu
jENXeD2Toe8jpdrg3ePtZPkYgIrRu8aO9By6AOIPHn2AkzZhXYVUgdlQkugKwTy3
UMyA9HoIKEseK/jfl4w+G1vdJUOzhJeUaxnH6gYK+I0IEK0AQZDbLdoHu8dLzubt
K0af4Wq6w5jo+qtxp7SUBihGggMekG9RSyvHQ5XWsJNQixcZzCSetstN1IkZSw6K
2Uy/c8z3KksgkCBg9OZjozDCkcXtmuSrLUBYriblTME3jT5ezcKI2tPqoRjaMWEQ
u2tLmcTi4rv+nVin2FkXu1HyAdMuhJW1PHm9q+6W7/qKchALd3x1fuZb4XjTJ2a2
Q1P0ERRQe9XuFQ+8IWPI1iiNxIKU2JuABcCDfVFW5u3U7Vi60jqDoXA4ujsmWRAM
KVcZvT/66M+jjLm4oKkflXAaTd6UCenIFRfk6FtBGKF/VLZthaDAYx7xXDWPvsK3
51R9pyUZYbYXqdylAXL5vI5m9bu+DW0cg9abjJa0xx8ju7bMkQ7VhmzDVHAik3vl
ypOZFJIVgSodKg2wbLzYEioJMBHsIbtGtKRIpigE+D4B/Wf5xPac9dzgJhvAs8Ik
9SgC4urIdwp6tY/mpsDM6vIuAI0T1DJhPdwm6x6Q0uitSTT099y/w7TkLNxKGT8x
XMYdOqh+/j4xp5BTSHW7YoLMDeg05akdqAOI7xF1pVzoNxdBgHIhb2oeMW7zs4i8
46Xu3usSKCph9g0BZvSo/lVBn3ygwzv1Kb+E4NtxCzFqeEX5n72D2Yn37VU1vCEc
MXCABhmfuX1Ap/qBZbSE4YwAGKcnbGL7E7LkylELmV3HGjWal2R0HbpLS10aaJFH
GBhTxeICgwFnOXSaBBULmoqKEm40+B+hThf+6pVrhVkJ5Fa/ls38JqtaniNo3NOC
tdKUO5ObPcDYQgnAr5z4F+cXWKHGkuwzsiLjvi4LuPBXu6fibo9Xq9QnLUzkKM59
uiRYpYXwykChgET/QU9Omhf/dp8DNgJOcMyWEMMI80VNvzoQ6yrklzljsRpUn5JR
c9yLwthXD1EAC6mNKs3T2ZJAnCDLYnQUFsvI+OU/yoXUyNZA1qUvAlG+wNGRWjbf
pAmi1ndGKpeq2ucbdN6C3oEuAtYVt8ZA6E9PwSj6zkg/mBhpS5gHtZijUXlEyjbq
dZrf1lmugK/E/RExzHp7lHueIJWI358uRGTEHE/zlPBAGi0UYAQTQ5oNBzN/YFlm
HzZmMeaf+kBRjQb8nAkgr6uNKOUCbGxBgGRLSeCAdb3uLjYdcuuQyLMYV//IYWSP
WQpUQksZKW4xvFIffoNdzYnbwGr14nsYCUjDpMyuf1dHa9gyPbIMKPbmvNxRAZ7O
Z0lg2rI/X+J/+2MAFnFMcsUY7Jo5VCRbs5JL9nFpdecetAJDUrDDXUZushpYybRu
TYq+ZXfEdix+OVothQzOAhPGRqNWlzMBklh0ZZIiZBTAwcCj4IgrCApHOCNy9nAO
+7fq5gRfZ2Vii8sBlOp06Yc5nQp6cWB8i7+EjMd1bEYfOrRjHuLu1RIDt/5oqSPF
WDDgQHq+HSBdZwisZI4exy35kzwMW8zUr2wX5bM8VWCFnx1RISzlyUWHuE72tc3d
4sjr2ZDrJQh4TCWc5LVD1jU3CC9yZLTtIOxBe7d0xfwJg7yXfGMMmPzfvFK2oc+c
WeHoKs+aAT2lIBb+/SwuyjwhwF2yTcKkLGWksGNq6txwm9yB1tcC8sIV3y+cjYd7
hOM2tGi3ouNbIlbdEjyGI6Iq/OYcdiTeb7vHTGRVlU7J+F3M0FQIFOZTOlUS7F8a
bwiT6pCr+7Akh3ytyrurY66LefFKfZSJX43U6q2ui7oYwbHECT3xwAFHYt7/RuUA
eiHAUj/HeDfNf6JLXKhmvps3WTnKlRnsJ2la+n/0PQ9sAwsHU21dU+3TtayshS4o
oyKODzyTVF2QCXiUa5jLcWkBsGgyAo10F3CAHpyQMUkuGdzgOtB6S4edRHoXxorC
nw/qU0KzbmqBKWhf8jLQhBeJ3u3NWrmdI4OryNPKfohJvgXHbUOfIXZrw8tQqUl8
zuBTtUu2F4ZvTNGI7WNRd9ER9bhvPUxVYEk/jYU4RQTfOYq06slCHUutnYEdu0r/
sIBkB7CRnUkiIN3/vvWxvA==
`pragma protect end_protected
