// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TyQy5Jx9H66qbuKDRwjfzx1el1Q31MNI35A9VTIeERmX1h+3mHmzK0Xe8kD0uMLT
uiosP7FiyP5nX56+P5pmEbgnVN3QcyR0Mso9quYNc9OhA59Lc8NOITVCrKkZCrMv
v+OBlETD4TlflWP5itNJU/Ffr6s+Y7y+x/Mp1bGFZB0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42880)
Kn94y9aVNc+FrxL4+Xi40V7Sqwxz8l4sOdOP7z0PXtHZX5SuGZtVTAgnqrhJIUeh
hSRrBTsL058Odl4/9sEiwVGTMbRKId+SPUZi/qaKLazpOYHBh10cD9aSEh90yKHf
M0nwv2CdMLcKCB36EIvsWpVun/FAFpAmtZnHB26SlzNJaMoeagN8xCzCNyx8gmHN
BIUuEycChxh2ohaipiy6qNMANHaGX96YRhw3QzD6if/VM9bhSgQBV6MLn8PCBGqn
3KonqcAWg7feI30BMeu9SGc3B+BZBPhPeJ7mCQouU4fN9C4CtYglEdRIau1AYY/Q
4l6bMNWIrg6/GDl0VCYbq28YI3iJou1rsaKotmZ7YoPnC5zcJXsbXgkLBRChYhc+
Um4XMGCSdknTUFYMXM/RbErEhMX7HBx37tfVSv7sXAdF9UWz4aMvZmfwF/5Q81ai
GbSdWWeylE9C/7MM6EaNmtAeb3PWSm2Oxx1VXT4RxZhQHA2IAty+RsOCI5pQgwe6
vR7+aF0lG3eN4zv3Ns6Oh2bKHOh+wittiTYKLcLnDj4NeNh+lO7OAdHGz/D7Apz5
0lT4UMnlX0TGQfg3NWaEPH9s6r9up7lvCQUZdqXHa2ZgoF3pYOXENAFdG/5CAoqs
rew7OcnUQLMWh7TpPkYfNOp5OhP9cbo1u8OOW3vMiaRYDT2r+KktfO8Ke9HQnIW1
d1p7B8yxDciphnIpr8GaYeR0qmJ9eUlbROZdhaDlSJfCI0QLz8Qm/xeGnYTePnpK
sp3N5nL39GAgYG9Ma3TTrsiWKtjbSl1FjZNcrwebu7o3mko4qDxJdd+lEbtSrhWY
JvBjHbUTEfEn5qpq8YUt4UtYa+TEz//8qW2CtYaei1JS8siUMeqA9AIV8su9IWkf
7ih65V/gLANBICUlK4M3lj/xVg/2w83NiXz/T9agxfkI0BiG3xYUybEF9hREhnwY
CchDdAONnbUYhIZbqRLxJpfmbje2bwWfReyWqaCBQWwraBTwrM7X6MD5Ok5PQ3fO
I+vc4ipPheLGdxt1aH1GrasPllstah7qnaWFJDO1f5/dE8jalmQfV+f6Eh6+zUmF
D0sA5g+5KueO3Ofej7T+Vr6mtGn2Gn3OohwJUwZI5bMjquwzNHsDqLm8jRhIv4Pb
oSyyd3xzpfeDQYrm4sNYENzECQg6At8MvozOiwSeab81wdeU3lLT93c4MKTmw/5B
1MmFSbAs77YtgvHkoMLigS/NVkrbPx/zrgyWLjP4VpxBFTg61/1yjUSjuFsCb6bb
oGA3RULwd+FGHbOR8G5NnMcMRS9hd5DcmgHVnXEia8/COvNhxquTJ77wtji4+a8h
eQzLMTsFxiH64VRGFtQs4WpL910NssnW8zVq+4KFMKWglQf4FSI/huCkEUx8iNn7
PklV4zNhk1ySxRnnXc/sUn5nP1x229I+ner3qqSvWxoXhnFItB92MyiI+4T8d6tu
mxdBXyRWtsDDBVG9LARY9rCk3Lln3LY9EZmTKHIcKmF6k06lciB3NRq0nDwR1L/d
Q2Z8MbZX0kILO26Y2RZfUkNstmgWEY/0FHwqGON8e2QELiApKxwXzb2sBaeTLSbd
X415XQmDC9HMgiZ/+SV3JB+CxH4RgG8fpuYZCenSYfzNxHWdmBG9T5Z735L0nEWJ
S/opUqxUcg9Av80KAHnRy1P/wcffOmAhlIapBNhNaISPRiPNlfk8hj6t8HVt7NjW
9fVmP7jb8C0Bug1kAMhLWhUuh8WONHkLJPr49wvRS1s5FePgXEW5Ifs6HCokLRMk
uV5/sZknBZC9g/O4BYgmAqOTiwPf/lLcXyppW5z2dvAHkdLKRbMrVg75SXemedfB
3CmlrU/W3mfbBOKKmQymLsx6+3q5r3CFOcdEc3pQ/RyXCxnJVFNLXHQf4HBVJSLk
bXI86w8DgcfG38fta+xjyf7G9804I3TFUyWGjn3WhBbYmChAxS/VA/1u/RhmWqrZ
nfduKjZIa3na8t09x8DjL61HcEbCOqvCE9OvF52AfBdgiyphkoMRnFifF/MJR4BV
wdOiS/BDRmN2VXQS+xITy+KFnCTYiGf3NkngElS5pCpBtmQGAbyDr+MQCeCGMIkZ
0Bj1Zou30uU0+msJ1gFiWxDPbfaNW58IgAgXhnDJFl3bJTevvXXL5lOCijBzIyKa
IToi/Jp69sNtH7DDY9QFZsvH54LbCc/zC7SxP9kM3z7c4TV4NZ63WLrMuVWd7Ia6
lOaRNp/ZvjHl+EGgWC6hV5dow8cXCJSK2VPsbh75RRqRM/uQREDVAzKUx9AJTa6a
zXFDYSzfLoRfvUwKbcJkGpSHRixSHUueGs60bBkovHsTTYVFG1yccLVperysjntr
T7cxqsmfTtvC269+c5IbsO871oYM1LtnTP/AXgMmNVt89Ml1mG3ppzb2vlsq5hLh
ENV9rgeXrCQZPvAshJrU/xikP/cJY+QU4aTUQquhfdwfuIJsKeU+STp3e7BNxlOD
5Bh33iP7KCgokxA5I53+Af5N6FRmGfWjvjhP8yXMWa5RH4s0etwnDuvi8eMwkldt
RpLAhqsKyjvXa9JN7Jr2gWPU1xdqG1cy8KKryA3UDr1cTag6QuFV+EOKvsRklCGd
1yasvfK8JjZhpaAFEqVF+oOD/76AOy4V+If5MKoGzGRen8c441MT1Q9fpymxn7dO
+9DxVzkGKrDClri42JcpQPyOjPp/BBypJGcsJdT7ZWoykbnLQwSLXGoXVxtQIxgq
wzfHDjI3LVdJUaZ6MAIEQV7/uIM7pzEUmGeU2u59B0ZAu7M6I/3xj021pHRmMDCP
hrvVrPDF3cEKGd8JJjh4KcxeYAmGM5FBWxwCAUYVEjENThosfjrnX6lOHH5IUbIk
GbIVjwiaz8rLOq1bZc7scxmmcod5Wkr3SYks3fcI3l+agqR7BERtYmKRjTzRON5e
gjPfuV+IJVgAUCUSS0amog0jTxptkR3vl4ZH/5xo/h890DQaxaEA3X6kha5eToq3
ei93IzQv9U4F7ycjkapsvdQucpPG2eajvjXoX5fjizvbMA0RmnP9hPHIfMxKJ5nj
BjXJGtPYgAB7ok0ZJiNZGcuxIJgdjOmLAsTSY32lzNBCOab4vk+B8CvwICmMI1NU
TsupQmjNbtKtTHxtooK8gGO2Ec1I1g9P4KNpqwheObRDovJlRtMByguyz5TjKYhL
eg77e/yMXLwN0gEdWtsRkV8BZCixlPvHhOroGhU5OfbURIlQxnAehrYADdYyzZS0
Kh/PVI0aW20Jb6magaRWBvot8GLLnBAii/yQl1+HuoWn2KbGeXLt/glwSOp6syUf
Jbj0X4DzqqLVDA90iU5y2faJrD/NU5u4ZPXu87JGMcpirL5kiKfvdJHaNqiOpR9i
+bGmXd9HsMVRy2MrpwfUbIOty6MQYP83phO4NW2HudN6bZU7CqFTvIqYRvuomKXy
Rnifmtf7m4X4x0Enui2h3IjfT99aq3hKrw95B4AagUj9JrXKh4ZgoCDzCtSO6/rU
6rgImmibKS/NXDO9DOi7eLfk27rX/Vfn1jn3Fh/pA1IOJ2O1hIABJGjy3tZxvCQn
8xRhfyhu5TyiBruPKnbKUiffIHWj2NtZ1NwNx0oZn0uesMFFL1DG6jvQFyiyDXay
BnRb9s+H2Qwv/72XGa05D1/oxCCrPAA72PiOhF23zT7DNhUCon7CqVRTFBuB2OOI
Xq4vgrA2LM5b+0yqzuQSHiaBZLLf5eCXiI/Yym0YBi68DOrwvCABcoVAzoYqIl8K
Kij6lRj/xUGmmuptabbZUwiqqRffbLpcApWw/jbFq68HZeSnC9gyw1aX05giod71
QzowKUSQnXMMQ+0sSNuqBiHhe00M2JO5cnKDqbC1EqxgkCMoAq9YywfxMlJ0vIaI
9mVHMSE+7iMfgFMtlDyQm/JHp48vdKa7zj+HoBZLeSqakFSY5d4qSKqqACxL5qyY
cyHLJ0viF+5wyEtQj/PU2ObgPGGxWlr9g+WV8Keml0vvteStKCoTD2TwZKUhxLk0
u5yF3FPnWuLsHyqMDSN+awlN2Pi6Mt4a7QnOLy+zsTaph61UQJ8JZM2vhfTO14wg
/0yjVazJNDy+XuneAnYBLXbMwtIffXakMMRlIhApF40Ackdg4Paz+7QacZShajEc
1Wl4L4SFLKJCcJPKoJgz+wntWNK08VpCb5hZhJWXw0AuZCwoJ9+acXZLozlyaPBq
sCm3J5BtcuCBq9Z4F69tXLOugif57WYdB0ocWlhUCW5kSW1mqjePq6LLvdE5DLIG
jbE/FLb11gpriJX/pi+gtidGbOmzH6hoSlnABMdh07l9nvKHriMlWfvnpVuH6fXs
Rp+iSF/Eq6QjMmzaEjVSkeBdZBQ4cjWZX/WTGGzVLjwtirhFDWV9Ovml6Iov05jI
BSsRS5OW3/IKx6ZXStxd9aI4boCOx8gabech7T0YMXqLB7IdVTn93cURoZtRsS2K
CcFzw43ZwCJjjX+Z9IDpYrXjCM8ECPFPfejwjCNhDrCgk98ESk1SWPOgIhGYalF0
Nq0don/IR9NDdkwkE+Go+fcJeUab3Tk9A95z+Wi3vgE5vG71tktGjk4cJYzhFp6E
GpV4MRIA6lhQq/65fceQa5KAagea9ioManVej7Cg+WSrEseZZx6MMg4IwIWIivBa
9Lqptpr5T5tzEXL9sWOydLomm8K/KDJQHQCFsErKwkbTGxWNJuWRqs2iO/aKItAO
fjwdi3V7r18YHgP4Ee7zO/GUNHrBJs96V4OUW5aCanpvu5TiW4Sea54Do34ExW7S
XAW+im7V9VCoPHw/SKZ0hltEhr0z87ztFZmSCYCzpJObsgOKXpMQqHANh09+INzn
GKI3x6eVqmVzNFw6/L5dwBXPHA/I54EqHdos5y5inoqOlabpCZsnhWfC6PgEw6pP
mr90EnF6W3eKgMakfkuLdscPNZivhVw1M93RJOKE4BmhZdFHj2jwSNCP572DRueC
eZwXpTmezRHEwXgfDD24E0ZuGT5TrN3gGb69JBAK9k4+T1hLjyfivdL5thRo/qz6
fgOwDkVYMC9HLyLsvVHriO/isF4vQ2g4lfO5Lit+/btGO9n9SaUejkKtIE1ZUAsR
T0vKXVgoWXNl6kWup/xYL8GILCA+xWCfo0jNy12FXAd6nkpdL0BIVoxTY6ORFZIs
7YtYwc/Egqa+jmtuKLPSzUh8uCq6Jxr4OKSNlhubPT+paDQ1kXMDcVew03CoJ8JX
FIdbrn7XJU1gS+VDgZNwG29EpIDBhPlDsSDDGhYWSsvtfiXNJbIREHjOKVrAFEaY
W3NPYz9pb5jAZAnXyzTYXzTiSX1MWwGIB6QC313ah363KCT1lYHfc1FIdgK9rJX4
SXubOlqGvPSjMPhrLu9JDw8emMZzfzTR5movtolgi7Qo1WFMTFnQFnJqKbw7yiaz
bgKDGDXr/T6xpXBnK+2jhmgLdjeRjpi8BbD6KM+RJTkq8t+6E+uU4UzLpDT4rqRH
W7MdOT+HhJfOkGM/drweIbw3b/FraXCipNSl7QleGJBljjERAcZPeun7I5p9fs25
S/lJqaNSEdfZhKwfn+ZtzGD3jk9wL+ehUFFRSw+RGU4MONLcsLx0w35CwONrJuhU
P6UBMAteawtvlQiwiAe1E4i3s/vk5eCYUWhm6Nnrpfvb0g9dxUGMxI/ydZGhuj5F
HVeo0iXPXTuBTX1Uye8SzFg3jSWOsKMF86xWp03N3dDAN4GBzkgOaZ7mhNN4Plca
e5kL4tbamhEfZh1VXtf1GYUi8BdtnbmRxnRIdINFZVPA+8zMhnWR9EjtUdF9/4uT
8NAQ760GQFoa6YthHb1er2mK3wlFQCeK2hW+26K6OP6GjixkfEVeeOX+2GEq9/9V
QM5NL30esmYjuEZiUuDKa4rRogB+O9X3bnszO+kjqirevdnlQ4eBJPQjMUpFkxQZ
Z5GMV3cKXh7Kywbp9rWEQErDbBTvn8QL88GtnRe0K4Vid/EVqx+Yp76zb1BDGSfb
Xd/Oq2/g1FtHj9DMyUooGShe1G6j6bXyYwEnWZ361HOY/pjl6gQ52Oc6wX1bzKVD
oxHhcCEfGm4RCjVc6mD6qn75K2KzDJUy0gxWgcUR3zZSnTFXh5fJyyeJnwsq6KRt
3lYC4+tm3LvxMFsoDkiPEF/Tsi2Kcbl42RH1ZDEWSIrORLq2O71JRb1v4pQ/vIKN
fEM7av9z6l8+Zq9kBLk47KTPHEvJElK9fqeXKwM8f/2sNIm3xcXDpPDK58ylQ9Uy
oHPi6d3r5Cjf4gFV6nUOTJqrGiH2Yr163lDaWpHHGga2bjoYqudndWI9hIS1PQVf
F/JDjpZBscgNyXO8kayfcQ8MEC9nMg816PenwVsYPD7z0uNtGSNQxiw/PQWnEHQw
jI1ptP+lvHORxPbk9N0SCDIlNcZmlYjUwNY3bpisZxYQYoylHR91W+Bsklc+hmC7
nsnubb2aRN4uSu+DyAINNLnq7wRZKD1qCMsWD/kqmDF5qVJ+0xgzw1ThvUsfIRLp
/2J3Kvy5sYR7q1wjE5e2jS2juJ115fcbv1pRmc6i7xvFPGVHySnZtJIZoOFP72FN
0G9pjzdA64/qiYx6lrAYovleuCnSt3xEsRw0u8tcBuVur2DXbcAJT5NF/u/bDqxt
jWRmkeMPufp7yRzGuCfPfszBMM2BDkux7xSLjW33fL3WXWk/upeae5YPIpL8Ddhg
eSA+c4TTN68FnEjGNmeI9xLo7HCiz10URq9rjR/T8QT8wam7SdnFlsYhRJ02BAIX
Tf8iOXmvNNmTvcZpuBYityL58D/3Vy4yDKRARu6bCj5lDDHDIALLRJUDpjLTHOvU
oLF/v2QcBB293Q5XE60YXpY7ko2Y6asRJJJ8h1lZ8q7SkmM2LChYo5AZwh55UQUg
2mGV5KxqNPkOsHnrTz7G0XC1dU7fMREiJ/MImG0aAWBZqjJJ93vcLizNCcK/r4v6
5eCbrnQ+rP9Ju/JzUmR7dUxl5zZnyConvCLLjtv0/wwuWaPbFDunaI+2rOxRqpre
z5//LRD8LXYqordfscXZ6HTdRuLPiGbzHQowwqrXvewF78NjBCSV7sOZdY+Ib7N1
hdu1DjAJOIY8yiEMEzBZJDKgEv62uVLpD/TIwHL1sVnl/dn+hfpqrAKqo7edm3Xi
wvNkUGlih3o16fgHkdoUuFCYMLt0RGMeIY+0+qTN8Y8NFjZbp956d2mh/WhjNJDH
+x89n7J18MkrntfhRZa7ZiiYQOuxm1FJ/38R2wbO2klCB1TwvjArxEwlfBmV+bvQ
sRvOnsnY3B9dDVpKudhXiaE9lRCN+EElFgaakCpePZyZB3vRZLUA19Z3sizk0ah+
QTwaPvaPPDkohWYbhp5+6/A7HMYzCXfkuk6HqVycfyabwu4R6iLbTal9mD+y6fdI
rHldCpZYvkBWPAMMjVk2jK/si2CoYOvNPvFcZuJcTkwaceWoeyMao9vamaRDw8SO
uXBHv5Y5JSYucin5pPoAr96nJn/elulpMm+K3wdtd6I+QZxXVJQRmx9Ba7knOdWw
fjNCYozCLgvQ7NAmCmOcRZCOM2RQDkf3UdBNflXProiG+xE0y8m2M/GbKjNot997
qrZYtJTZybiy1avJ6oJ6s1mTGs32jtyiTxR06C01CU+nkQqNfD9i1Jsv7hs5VJJx
72e3aJtzG+4HbA3vJxmBs1+Z6cSyvJcIpxHFrSxF9sdezCgnDCcQJ7ttw1ACwIXA
Jduf4m2M7x8Gq56DcPKeMZzgypdd968WeeTSIF4aT/sib1YXVzfL+pM9alyqHU0I
0Jjlk48rGmyfXd2FiV8l64ryuTcbircdPCtvOszWLOsCI/2TgDK+Gp6zt7cuTgSj
bjYQXEv5asPcplVtnwHCc+0gHslKXgrxzVSyHtyFwkyqsFU/ZyVzEw8fyHhMU30h
xdnWD6a1aCUNUTQQ2/5kRN1yU9ZIkYLaekjTzvRWU0yv3JMxPilMJamwxV8VSAgP
AOxc9/n4sPq5EE+0EWbFn/+j/B90cQSwp2ZDuzhNtjaYwRnwvYKCD4RmxdK/rvu2
5VeDhxgs1g2oZsGU0J3eWXXvH9LsVripQ+7xTZmWutXIhJmgZKSbx0jEIXXokABU
NZ2HWiHdEe5ZwerKgmpX9VbZnMtT9NvMLpcGtIeJaYLdGlbwxxwUWjsUyEA8ETmk
FIzsFNBfPHRO50y+iztqb2NWnvSqNlqfkwGFlUMEeb25FYxmhyL7E/qhOounEWDa
RAVWpnyMVJZh2ns7ZAC5jHsPFK0OerAzL00ltwaDNPb+X62/IHElis/4WHAV6YtM
yVWMARucN5dHJi6is7bDPArzMa/GKkQOb/Xq7CRPq98kn7SAzAwaOs/W3sXWmzjM
Y0PJ+T00STf6LnOU0d4uPUkkQE7ygmc74m79dQ+K+rao71AtT8z6DxAhUVTl6xPX
IMHKnV1KGF54OhVtidHMUiAQMIa7FL4t2/zc2hj3C1W5qHnd/SJi4sacn5bNfuFT
7fJLNEl2g5jBKpnTl8h4HQrg4OqP1d54bZgXeEytNetVDL6yv1xlAeV3pElFZaPD
sBy2Df/Ey0DxBVRUfUfSZBGduj5oGKcVuY6xKkdzjj4r17Hrpf5SpspE5CGXpegn
klVVAsQd7OvTlACYSgW4ccvS8Vkwct1XSgv8nq6hN8jUPtpjwy1o5K6qGIJsKFW/
RV+O2XZj2G6EPVdbaLGvXt1Nto9uch+hYFA7nVcshlwbrPYglWXsuu2EiYIZZrTO
moYzPAM0CDj+/mQe/CvvqCNuqy7DttPmm2PtBYe25XvIZRGC2HiovfT8n9Fxv+YT
7iCohzIVGoBygw56mpULF8ZUmRFZNL/gTvAk4EveDcun93VY2+z+7t4hdPAwE4NS
lvGCElOJjA26zQYWk7EU2MMGWroS5l9lwxlJNPE6G9fhBQThXG8DpHeX4sCkwd6t
85HKCb9ESeJrT3Al50xDE/dri+/nmaRvZk3ogNq+FWXA9R2/vQgff+v10SzmqEUU
hJjU4F/T5pfoDyHCCF/ywo+jZpPj7D3gyOquRU2MgBMZxnijhtnm50ZTdffjjjGw
ziEZn989lPw4QrMWwL5rhTr/t8Wa4LAd/tFCn9KA9ewKhm7XvYFKqH0L1Y0e4jd0
TlCoOKKIoJyFjSTMmVpW38HwwghEA6pP2JSOr5opW/NVNg1yU4nV8HvAJfi1yk7g
kQSWqOGMrrlMHGaqp8ttnjlp/xzBv68S9JzXOrAzbEqXirQTrCW3HgiH2RarMlX5
XLbjPoibqFu2qUiktFMbq4H2n5CmV17MrmKPi0V4D058lCQjFnXC5UqB/uBLeUND
+gyJcrAJY+Cezz1IMOVaeMdiKM9rd5XyxxfG2USjaIjVFV6TEdJMvupctJIJfusX
9oLzA6ZgE19Rh13gHPFpTNQzfRkSqOFiPSuSIe9cQ31Llk1fQRwMdjd7kXrv7p+6
Or/W2MJ2vtNkLoIzhGfnpPVa7KppNwu49aOhgNRRL06eaMqjUdGoss76r4vwA7Pr
cHwZPhuGY/d2D73ZER8Vw6Bleq03R6kT62cbCpWYRRgCpv6poB2vyg7UgqtE62uP
DKiX43RoiEwRXEUSiIihiOCwzA3Wi0dksZfsjrhXYCYfx+PEaqZWaCYQn5MSC9/c
Olf1B2ukvLufU5Pf4w95OEqPFt64rkqL2I99AoEKc10crG/PQwQOe33+a+b12Z/R
N/xbFSofXe2SiZmw24cxA+uin82SdLxU0Xx/sbEPwa5dBKSeyseuWgjvidtvvmUI
8gWTaP0rIz7173bTbwQx8mYMSmiABY4DFbn8Bd2kUEMwC+IDimGHHFhyqhzkH53G
zRQpJ5EHMRTeV3XjnfCAcm4ln5K+BIiufZZRk18dq3nD4s27BORCeBc0uWWq3ytf
NDT1uhqEdSI1PpQ3ZNXta7g3L0J6nqWOXoH6WFY9yQkYoHvv7Hm8AP8MIAPUyrCw
PAwsvnsqBrvYJTBdwHQgkweUFkiFuDmKQs6TnVULrmRqpjZuY6KD/q+kLl0GsTBh
GaSw6h42whp0C97eeXQctbWvqSNnGV22b7zVcofj2RUnp+ZFrFx4+yWqcXykc4In
qJuTeWgjTeVAJahht4X77MD2QBzoGUoZ2rLQ4k83TwIB0weTp3YnYabSR+7JToxY
eMPl20KgPsUbF0VLUJGr9Mg9wCSeUn1Sgh5B6851WHppfc0gDHpSxbvKFR2MSXTf
JfCSExSvPPoEb9z/Y5bBFc6R7veApLqf4sOt5+npSnaG5PIqRzaZ0tkJqbRS312l
uAkNVuK3bBJTUfrvGl5/KVNMoMLHqGyCZt11OxLx5aGUdsF7UkA0uuBK4dphCzQv
ECwjbsP/UPmJQEd8SzScqqiZNrgRgZhp7X4rWvlJElemrnbLRb4elL1qxFkSnF60
+whIB3cSdIBIARFNBOSY6x778dHOUI6QITn5GXYRwE7GoJqrRV6k8BW5W3MIfiWx
BKAHP1tEd/jAknb2g8tYuNl1C6tXlQL1C8j6u4o1n/02n0lSJWsvpjT82A6Vbn9/
DBfoyjemXJZb3g8u2k/YyWLsoFMbZklS/OOnTb0tkKPa0D0qxXacv6rBqCHbuMnn
+ym8atPZkwJcvGYMZY1jQU+4aS+HintyVv88mNTQlgJObHV7Sc/L83J6DfLo1c/q
deQfKmO2YYjRXX7gOnadhnbf1ejZW8wpo+WQYhCL4pSmFiGK6hLVbqzjztgpa1Lv
N8NuIWvi9gJBxsS2N00rX++qCE51v4G6/w71yteUid4MaVvGObGwcA27S2YgcXP0
ibpCAQwOPkG65QQcg+VrqiACz8rm5GramDsJqD4y2mdewdVQchl89VmqTIAuJlpR
EsAYg2hI/UFmnp7NNRR0LfLhC9GXC8B2m+IHiOQyBxtVt1QgLlP/FftASrCtLnGV
agjDy2G4p5pQTNhR+v7XFCrBxPoYTlm+alIZTx2/2PYELSenCCr1+7Vmx/kCCXNe
y5RWYvo98zEIX1key3IFMSyQE0YOOwF2lL4/zwl8iJf+ZSuicLZgXTJFH7TKVYZK
V8j/y9Dq4S+l63gWYfIJfeyd0d2MUlDC4aEmY8Rjj6fedBN6LZS5FYhax7gTGfC4
y8lZPd0Uc/uMO25rcInrSmRipWu0+EJv4aYJnRPgGf8vJYlgUG4jtlWD0GKoTORN
Z/9/QlpOypAwNOa5HHLWMn5/QgjxxJMlYd78ucqJvpABTVkA/EX3VcIf/pBCHj7c
WlOz3HjTF6rV3+Kp7B5l2l3fHDlyYmoZ1FjnsnNy4OtgzbhdDqmLz9A2ci4Jrh0y
6bw8bKBRCIMSGG+aNOkgmbhWmmeuRIh6blZhgeVwjhhA1COGgHRWuAwzUKRwMlGi
gb7b7EUoAAsynbaMfThCXW/Q77voWD9dOJnH//LdoWd39Wkmb++YY7qm3MTUnlmY
p5rHZL8ZZV7KOmQSWfGXYAgIQEze/iEBeidEX2tjEFf3KrpNAFwe6Y55RlCgptm9
ntZ7bK7xbj+rYSODrxgipIVeGS//etWixAR16D0ZsE5rEW/F47KOA35RT+KJKKx7
F+n4uUGAsPlHxLoZDiv6aZm8h19BDuW99JWxWU5TbQ5ymbJ153cP04TRXmeyoo6+
2jqmc/suC61honEL61t/5CjNUWUdCyJc4FPd4arw1lH+oxWMRZdUphrWjPdGylFV
jKK1AFzQxNj52aBOePBgLYfFwyKTG36hGSMVY7OQPNZwmmyeSX6VbD/Z4rpBqYPU
/uAMq69uDnIPp05SPJGEZuT5/apTzdPx3K/b+wk31WhIQJj6/JywKKexEE/z2bpX
qsQ+y4MWQ1EdAgA5qGohHBg0ZMkt6lWo0luoqVEWtMM27O1o3TggM0mVZ4uilZ12
6DuyRukRvKeCNLYfokz+ctVzSvg2hpR8siwz6zQs+9wv22puIJIDkQcg1k5NVI4o
IEOtnyFR5oaUtpB6zVrrROECjCepB6d+7H+TyTu5wLBa/Ri6zxTmbPqjBoMkvgNo
LbX1sZTkmE/OkL3IMSE2wg9QI1s9sdI3KLGR58MU+aKYuqZcJCUxanA5MUASz8L+
ZuQqQegPV35fwGUQjvnCaX3HUiCsFma3CdyJkSfzFBdYEFMC4VHdyEBiTHfbkMIE
3E73qgT3K5pLKrs2vlT1HcU4W+U8/hiUZ65Jv+ZhAZ1tECbtxUqkwvXm6dL74W4s
y8IXzES4JcR7So7go72UAZd5P+eLZiUz3quWPi/1KR9OrcLsFy//0R+zY+q6qItq
V/2n9mQqDqH1VPuCEV0hUiHdUHhUqP6gWlQqpDilUQtQ774rdz1n88aKfxsFjxdW
PFYEWzDUsHsI7adYRUaTqsgTO7yO4+tDcCNUrfEkPbMZ018HxGRBX4zeMf4cPIik
SP2nq7DVD4cyGZ6uRWobG2uSHl/gtP9JQ3GThtgBeeTc6TCobJ4s7vLSED1f/ZWE
EVypb27Xl8mQ9iRJ63oNOoxqOdjbT/WejfLUijnaWNyWfAOtbGef+P5cNMc4teyG
YfafnIeEw2PJ7C9VCCo9kHzmbwUuP9NOUaHxUQo8E+re6Md3zQPfDBIBTF8c7kFI
kdBfsJgFKWsmyjn3cZOobW4N1g60J4Vx8f7xzbvjZypXLgjsIKwQ0pqlsGQAoEsj
nhkQ7AXh4pHS5fajPOXXwnINxkl5KieDExw3zM4PnzfGbE427hJq01TVkppyPQS0
t/LFAP5zF1oErrsYLO79ZTaQPYkKeLu3k0NvaPQ9r0ny5IU/PvHK48Kc0jYrurwr
J2kbDp/lYE4XZDkRHlrZnwD11T71JY1hbYb1EpW5Cxpk4ka+i8fGctiC3l0wFYax
KaT3w5/JlR3dwUKTazHXLiSLIy1POVbiGVsYopewy17XYlTD/rapIrscgzWCbBoR
RbYfc6en5ULt9huX41MWVxVx6WsFmpMpvekVVmttcr4z3sxJzO/3zWF8WJnPvKIM
VzH84K6z0uKoA4EQyRgNkb03XcQzR6jGaMxQAP58woPOvMtU+ujFMcvFe2/PqZL+
el0dV/iBzqXm3Tn91PpnRcdPo5wEHxCAb+GIsXYpfqQZgQ9T5wE0nkiPOGcHd9oL
3f9E8KPa8QrIqzNl8gN2HMpvSviuptF8W/FMciUILgpqNHR/BadoNUN8tGONujIb
R1PY1m7ztoEp5bKp80ncuLahWPrqgN+wtIOyEvjVzFlbsmK6UpI87XAzgzOhrtR2
7wyZq0obzQtRsL1SLU6NpUWUBomS60hSEDNI5o1/6NLeCpqapdYs7FmGjqTdUx+t
D1COty404lz/GQF8h+HdjsLQ5/FzJGyg1S4/HH5z5Gq9I9jarJ0ZekNaTGludn7Y
vRlWGbyc6R9a0c4YBZrPl7TsKJr+f+tCqW87c+/gQWA75mqy6ptWg0bkB7bqEY9/
CdKqu8vbh/mDDaTljq93dJVN2WXlBEzFwKbVUqpyaVgm2fN+PWSxgzAUpJiDwizi
nQM1Sk4zcFBhP2RktkVhmHoExcrzp8r+8pPpZL48p+2p6cWfyjHeFHwjgDJMaRT9
1ElAXo4M/njpDgc0xj7biq4usIIGLI4DHybfIL64waICwT+Ece5zCoTFlCZrU/+8
GY6AcNioNqPGAhQpuXVmk3lO4+AkhuJA8p22bVLFl4455HRGFE5qVysECcQdZYqw
G26/03pj7sW4idC1MuaOv65FxcmyplOPnU4G9NM3qrdAh7br2QVb0mHvJ3BK8sgV
nJRst0r+ylLTINAX7jdqEoy7e8aE3Qgwp7keZCrdsVjgz/42etR7H+MV4+HoDhz5
J3omecHW1eBfxRo//7aeo+aS01S59Nl8ebR5i7snQ5YxJFFP+F7WPWkuNfNU7oDb
7UOSATN0Ih7+6kTxChRDrtqJbI0xr+Y0IG/UBH9+RhymrRFjvEkXe9pOgAGXZR6K
30WWWzHOEck47Firf/i9PGCxYDWfnev+thkHgu4DmKLSgTIM6Ry1UZypeWZYTxLU
uOD6I4KTPvzMOFPo6q3cCS6HggeR6m5R7azPmPIq0mXwbwt9vlM4MI8rtJB4IZRe
4pMCmRS0tXSVHEb/0uMtZO9ivzjsDMo88HfMvAyZfxVkIPEAhXtjGG0ztX6sDVIA
AL8LnKHf7/6txBxOacnlkxKNNr8wAdiuklhvIKnleIR4oVNDUZ97FECjFd99BPeB
0FF38kbQ0//JV5tmHUS9KegD4B/xdWXZRZUOsrAPRi5+8ZHmc1efbaYP+cajMXFU
9JMR9X5R+a10g58tonnvtYZq1bF39VVNN3/fRTWxaaRgVSNeN5bkcVbUGFleONVu
3SLtLhS4aWsx2UCYkKTAipz9l9vQxcVqbeW7uaXN+RNvz3ZZyMsSkcqyGYsM2UFa
vdJyUhwRZX3DQI0mR8uRTF4CtNZlvCM+uYGWUzTGCHbq+nhnwf6+Y1y+wWap2eob
cgr2DWN54IC8VFfpizdiphgyXxH2qw1mYpZUwoephNUyHc7kmK0CqzLsCWftkFJR
9NR1V9XbrMBEAi3p7R9DdG+EOT3CW3M1PdAQx6QgArGu7gIoNrZlXhxrpQJSXpgt
koY6L/PMG0tOFSCy9f5Jqf76iYJvyL37dK2MxTcvmJQALmskIOinDpZ/XUyTv03W
6U+r/fbfxGJQIK2kE0jtr3nb1E+BSm2JfjWqCvRjqG5XXi+c4WOHiIWb74BeOzEp
cuDUr2aWBb8rDu669ZgFnfuG90vS5tIhVLO6hCo9Tx0CfeIuDW9TDBvZQQaZ0/AG
8L2SAmYGtPZ2mtgbSPyyv7SbMEZvOJ7Ocq+/trAEUiKLFUlZ4noX3XpaQLwutoKt
eM2BbcSKSW0H0roiZFtQb81e3B3vJ6GqeF/JA0IHU2EzdH0D6yQIqB2Noje+LhnS
yde6p+xlvXnrHyi4rzL3IhPTdjcog8wmPxyXjWd31J7g1fjl+RrFIFAby/ZxiJL5
KfLLQQktZzT3NXoyertvm9QdvF1HLxEyvkx8AcB932XPTxDhJ+a60LUxCBcK7j1U
T5kjfp8K00aFoeJaBWeXIcKNqmUrXvuPXgRWWMvB7Qub9u0u5vyE0IhNyLlvA6/3
KvfxwBvX6aTdwHo9pxUQzYF0Ox3gX8IDVdYVTHhMW4PHPqzzEie880M9aIL1hgYF
dxG6bR9hJanWG8PbtBYkeDKLW/fn2DEtadF4fP7AWz55PxWpnMFKD9ti+/orBP9W
DsHJK1oVtUry3aoGSJj1wyQe4XEhUr5P+D4OpHurBp6WhgxJWjeMGsq2ggj0LZlG
FEG8bKiPj69l93C/rLTtzlh/L7lRt/2wEXrCSPuNwIz4koThRiWKv2863o9aGmgP
D4OJdzEttokOxJ/kD44QPYhijS2EMz6AdOUS2yQ51vpkzaFKueNSc0YA6d/SpNm0
br3rpg1ljAY2cwqVHQ7LdH11MXtE+0VWGsgDXQlEeA1ZZrN2/rr8YCZhQQ2iRmFJ
rSMyfiVB7/oqqr41ZeBgU8jTdfvQ+l1xFxclQb6dZUIOxeNWybXclh5pU6ZQYpAT
4hdOqrz3AjRv9AyGVN8jlhGHr1mAb6zKH4xN9Ec2FwO1yUoBmJHlI4uay3kBx5xR
tSFUSgQhLejRaS31G42ly3y9anlBuXsFrFAXUUUkuaDikHQWHGOb0o+f1s6XBSn6
zeA9mlIwRunoSfhRuHrxgVR5o482TTHNNn21zmgXfbd+f3tfqCUohPEnRg/qzj23
k+bnokF7vxz1+tcQfoXH08HngdJgUU5Ma/hgcfYryOhovtLBZB9hILJydYkEhFmh
x0odqEr/wUT/tPkJBZnW84KbnShhmxGOprMfMIL3wH04pGZJ1mZoN13BD5rrKvdE
IJAKNfnCOWmjQjEvfnTumwvrZKgOrtAAF5l02ZaWnfnVlpuZG8v8yVW8nEMxJkes
xNeZ+em319rdokBpT3Yz3GMuMP+kYpRkm2h3fjSSuUs+DrgJtZBCwX3FA+wnz70a
aX/zcdocyNbcswb4tVZzA2caQF96kAv+0Ai/tD0PuSV6N3vjndMhjFpTdcWS8Q33
AoZ1VD9nEyVOP5EHCtKaegq5+lYfz5Ira9M3NezQhaOCtNtfj9FYDmYJ1vn2DBMv
bpZlWWShyAfiRFOW4pzEGoutB3yzc+omuaXoAdDJkruLhXAsp/MADlrZ3dNcAfRj
mADXS4LljwXM7k8dQeuW3EPf+EJnJ6WYMotRJBwxHGNa1Rc3D69GMgxscJkvSzey
f/lQhgbWQZG6j2HPTDZXjPetW7Z4exaQGgYU2ZvNLx0IWsJvkBcACC05JTIe7vgT
PaC3EzhlsbOVvxwuWrXhqg34W8ZQZ7txsVZyA9Ap5rNXVNuxDoee+du24CFwr8x5
vaX1SSntIZa2LvQ7D7Dt8KG0ONkOfrTrlcGJN8GKq2+fvAdrHAyVg60geUFRRXTr
6Rm94uB/pCqRR8v8hO9jdx7fTMzlPI3IilFH3IVsbvBEIHXpFXr7hUgTxTcr1aiI
LloqQN/3D23xawpJMbwcX4DpXb1kc22uLYi5WllAM6LHFU3ATQM3+/Xk5NyGfGSH
ZVIaM2h9ItMkvOCAIMfcN5b8GLjgNl1RSSUafbGUZ3OGLeibeUF980WVOkVrZplb
OUoq5hQ6R7ZMtraYKXQsoO6qmr3aET7wzqRbYP40BA+582UQS03ns++OrnQ1wfhX
r1lg1uMaarcCGBs2+TTwGdF37OGfrB1i4TudgAlJgVKO/riOGH1pmPRN9kP5Kx/n
OZ/AYpkOznGFCMvEJoJ2lD9OG84sOd9gYsbEgaPkw7j0wVjgy/1BhUrfna97I4WX
VO+xwwtI/m2Pk0hsRsJkDd1kv+EvNdHhPNOIb2+XN0XWTUUSoMPpTlmYQFFqz1Ye
2deI2Ki9+BOVYwcQImM6Pl1XiqH0PxWcmc13nRXSUSKckqM65zBdnUlxlmngnCKt
mGorQo6qGN7/+kzHkpWBHTfB9HnQJ1aftpTQ6EQQTb3rl7rIIEneD8AYBbOf+kwP
j6CQuWhXbBsmN+h6suPk19t5OzJiu7074g+gLvHPi/kdt29jSjxXd0A9CAdMH6o5
WHj6hcsTzLkSV19yni6Sfmgx5Wzcg/oZQPXu07PdxPYghCe8fvlCSM/AR27o9svK
7bYhL16udY56lV+eSFW8C4ufwPwSfUAPcgJ3xlgfZka+h+9Jffds6+w8p/MTQ77K
EXb6uLd74wazUsTU4NF1fUDXYYjDSITsFsXw6XcUNjmyZq2a4B029ax4rYWYbz/L
8uzn3YPm5xSCOkNY14pGZL/Z+PZhl4eDj28ul+Q153nNMeReLHD9njVOMzDa/NIf
dti4pTltaDILNsqIj7L37JrQOxqqVuCLufDjfQtNIYZ+7XUsQdWCZGq78PfQFzWS
sUsjWKi8EaEtQ3WrWj42i0jjSHE1Z6+EbLpWcGaxarpoVnST7c/KV6i8AwuMION5
ySfxGzeP/EfBjBlpBt7D6lteCgaMheCwZbLdsVD46SOyXdv6jYowxhiskLA66lV4
CmGLIK3eE8+z7uORx2vS+el66Ws8eyz1V10dy8VafRpCEsyl7vnKc3xiNiXxzWf7
oYEMe4xYrbZcNw7XsgEzhDg7jD1FQ81vaPMZjnBYfZLgfzSR9sS+73olQo3fHSvh
L7OoS14CXJ52frrIvA8TiqxgATRzdTEkxaiBP1J7iT2H61XvMJmzg5eiguAjPOTl
q01W7NoGaC28cReLB8Nk2gctB1BFqB7dr7juRv14DcnHd1zJST4kBoVCoJSC4R+I
yZKTzU6fs3tRvBt46FmnqmqXZLNUDvEnKFV+qbtiMeYbMqt6uUb5vULCMUNrNogL
WDdoELr7+e+IEgKN9H3XngCp0Mp9cIQOj4v11m2kSJ1Gt3VJyOkO0OrMQa59M5r9
JhGNmEtGpCTlXqoSKvOaPwQBrifSX/MvrKaHjGTpg+uDYZK9KcVAQieneENX+t8+
jedtpvzGZC2s5MrQcU8keAXL7T1zJGdglQw1WxCp8sugBmS2ffl48qIFV5JhIYcx
y60v98SqOs2mqB0PYqjyylGQcRnOIlLY+GK0ZA0cKHHNSTUPSHc1z6DUzR4kHvpl
hl9QeE4A0dsYgN34W0LA6NppsA5FYCvTh8NYJ4yOvAzKuTU+WMCb6ks8CSUfS2HP
sLqKv0AS7QkNBwGlniE9Ub0Hwahm78ruXlJrH+/vup+aIb+Znp8POdCcNng4kKch
yisOAHe8FVzIlY/nOiEdfKeTf2JgGYiFLqkU/w4BshS909K2XMayjGAL8s0hXQec
/dkPPhOeiMGoyxxTJ3K4ykwYVFCSgjJKow2OPGztLgewmhjDGwAmVj2gsCCiPhhO
OXI+ZOzwXPMscI7U6I1STNfd7IRMqbHvHvoUlDi7I/Ba7+JNvPTt01iNOM0LnNCa
KrM3EPRMlGQ+voFOOyI0spA4pAu0oL8SIubAG1XYA9QbIwPO8hi3D2gVwGEw1zSn
pUyOAX0g7j64j0wJvBqrUchASzUmoa5QC8EexEmYvY+z84aj5lo6rqhVQ/hPKjVf
863bNgCM7o0bee5C3tayBem9MYJBCq6cYae/mMyMVXyyrJzkXDpp37as+aZqKXrK
jgpSs7ZtTXBj/RLhAWS0eaLWY2o/0V+2LWu7y1T+8Bf5WU6KzXIxUCja9t5O7Xzr
Rq07KSoK203+rsN3NbKSUWMsVg8I1DYy+RP56RixfbN9nF3SNX2mBLafOavfiPv6
6RIKpVzr35byR2mEYiTsyGxB0bGD6YJxC6URVQQc0PXreeBjkM55+8UXH6dIZIXX
c7N35g1JuPIW00c6bNArSdZXYJCBQSKr7zECi+27p+iYDmJaok4cHt5ZPNek3vmx
GvzBin+wVYtY4KgawhoKwHPfbR/tEYR7v9wpq9bSg0JZZ5fxongSaJwDBZTJaIrV
EpnBUwpbHqU84F/cbh8UFVix8ONfpLiMgjmtFjosrmHWjRleYSEDPaY2dkIxCtCn
LR1U1PnVkL6IOOYnI/LK6Rks76ses9EDWg9X97o2FlgcptI/jrY462ZGjjHk6TZ/
Y1uVPH8QzoNhnX2JoBm5Kp5ZiNSSzmZovOkoWwOPobANyHw8Rxd/f+KICy6BdThw
vbXIoybr92IsgCFA/BlSTdZGczBJPaMFDMPS4NwyVNznax1rrDv7xq7NQIjL2iC3
xJZTplWUGForejJuoBwt8HgXR5+ag90AgoA1e1QWe9c5P42ELA4cA45d+CF/XuRF
ueI1gzHfIf03KS8oir/5/QIr/a+XyGhpLnXSeZQwMG/P+dNtjrzZn1DZcWtseuG/
2wcNHmZM+Pc0uegKukSRmsnW+YeKhrarWuM6ux3sSfhx7Ni4A4BcXAEc+XYsHORy
yu7pC/6FPLpCSGLWpGZSiMo/I8L6nkRwE6+XOezqJRHAlbhs46SzU1lCh5KVy5WJ
MF3w+qrPtksMz/BevFI2K11a9XupKdXapNjPIk8q5Ql0wK1ovld/r52ZJNV57Q0E
Ym3uUX8KYnCZ2bwxa7HESc0UgOY7o12jvD5KSn0r2B2ptjxX1M7J9+99sh71Z+oU
qgc8ZlMYsdQDqr+fRIezAUNQzwlKAGbUw7BTd4wsoXM5NAOgkr3LF6TgLi7DkJdy
Sh6w3XrluQvCNdZ9XRa1WeodkIiJXcLRQoCJdtZ07AZvl1lXZ1WohM13p+ZWir4+
v0pOmroMl5YnR30Zq/SS5qlLl3Bhdw+u2AOT/zgcbCqnYQaO0eOeZH96ZH3+nQdq
ZrZQ5ZHJj9n+WCbfY2CghD0avG7eLtI5rKIKy0gb0sGvWruOY6hwvFq07tQNUCbJ
9s9RjO5kxk//kWvg6Kc/pX8A3NHacEXkoTPP+DquNOdWE65QaWdCDNFXO4oQF5dD
S+qwXJp6VQIRvi/ESVoWq9ED71P6ElAfa1suXCcZdhLkELzmtIjRp7tu0IVZTorD
yemYdXaiKIxETiqVaBHTBmuORQU3iWx3Wc+gs34B914HE5mKVq0pZcq00SpBmDoh
Pfsr9JEH6l+IxMdcV+9p/mrDIUkysXGySY/vlQw8Xn7qYF6Rdumgr3CQenqsdfwV
RYiynytpsCGylPveMTaJHFaJVAr2Ldi9TlMufDTLmaZ4FVSeaazXkYjWif7yI3W7
+KphfXU+bjigpszv+y12lbFgaVcjbiGefyl56wFbSkOl9DqinRqfukjDwDk3XmL5
4kV1zory4iu1KlVD5ZeFYiKQGaA0CxeFBF/9RVsGSJvyTgXAGKge7056ldVqfiBp
VG6svkpEDvmffN+GqY/SeQO0CJWDVZil6gFEZtLtTyaf701p+wDmM3+L3+Bi3NVU
HqCrURh6QNQAUPELBVA0z/Izze/Bw2U7Mcl+yto37abEBaPiOVxXXze3J9FEGr4V
uXjH0HrlqnftCV3bfy1k8ZxPNftnwjaqx6Kgb+zD7vwz2Z5YOVcSHfihZzTYxiB+
wtX4pZSW89vXfJ9IzVwdaTkq17CdQcTMyqxxXukFmBEpWv7W/Qidu2ENvyDdQ1rg
ssuCUoKpka1bFChtsykXdrQ2SjqQj4o6cwtN/ROE0opTFvjm7tq6SXxV5rtJrv6T
7u1JH0FylQ7vuXbw/qMSvzMkxklqH7SV32xMQSyyVHPFQoq4On4azVQJA303UzV8
HU3Zng0Cb/8IJuMilXUBOUarRwNMMr4AoOcq7Wc0MshSXOvxCA+9WIIADguWTGin
dSXyFR3TKafUVZqvdXpR5eVTLWLXF7pnoqrBmiv7WCvntJzL/kXjqpHZYxah2zkG
bFkDghwaKoaqA1NpczNoJWYaN00Uaa+vMIPp4YDhr8of4FzyH0XLmu4ikZmV4Ef2
YDCWzXBbRmHA6zxTWHyagWmblkHbUYIYr4ETaFsrp8KCyOQeWArWmCRMM9iskD0h
hKDw5awBavHJHA2Fknaa5vW0Tregk8BZqoVPVPLUD8P8OTH2uSYG1hUJKD2SkMKK
i43aDZOVG2E1fNW6jfrAg1Kc73Bs0o6+mT1t9eMi1lCPey1AGfHrdPa7oMuOeGYx
HMWpU6mNiwiVPHT5YBRHu2ptenQMKzPtyqr0qya0SFUSXjbiPXqPwOfmhENdpK/c
DufEkunoGuBCusOyiYnu+xnP37ODmUMb5a1kLrA7cWX/bV/Onj2b57Pie7/sdKIE
cN9j90HtarMDfijyn9tkkpOR69WwHrkONtaS8rBga7mLJBQ8KVc5BxkEz3qcD0+y
l0167bhe6xO2DX4ZNFprCKtZd+b6xTrL1PB3W+slhkJVqD1uv/TgqQsdYP67d6HD
nEs3shJXA9bF8yUbfJbkrOSBIfHUIhZgSOyVoHUPDQz+nigCd6UoRNulc/2rxE+5
kt1pk3KbdxMHifJ9Bl08n9iwQoB7FrmOAPO7Dz7jjEYZyKiJCcoLdHq5o22MFze8
HYKe7QL94nC96y2eS0+9RSZHoRLpnMK/QjWRFZs6ig8D5bmy+v5jQdNeohOp34gr
V8LKxSTP7aOzqkVL9hB4HiMPcq9YcKSqE5ZV+c1M2gzuNeJcJBVdBNHu8oLUSSd5
/sc4Pmnef7gw1BbONjIMLA7kFuDPnt96xttucWVO+nFaO8b1NS+5H+88oy+XoYo+
mZfYc5PIX77WKMKxIJvmcNhCvZJ+IgT3uJ5z1BjhOBtLZeC4fisuw0qNSmjzOxhq
1hNvRHMGx4CctsjxNA4AIqYQCkGnXGC3xw0/ZeZYODSbH4a/vo9TNFmwy936N+9x
vtT9DQGHksoEWDDow0sQu+aNPmcxrhuvC7AV1hF0uuZmxZXXZZ5PhJyhdtznPtYm
P8pnKXPk5axG03C4hTt+vy1CV8mK6jyNfmu9H2ZuMEYRIxH2VKy0uBlGqSWMfWeN
FK7cXjpJSj2Pidhk3rNfEf55VWQs7R2CfcUp2Q9+VW36ycP8BDYqOWilnzM2Pmp0
/0JT8AiT9M5rSK7zq76LgYu/7kvRv501l2kUNwbHhHk0M6M9/47fk+IkZJ9m/wez
gBm9Dv2I7xR8SBdP7krrhoHGPNNEoeOiyUlU6Q/0HD5tCfvtXJmn4SlJN/MmlxTQ
MmnuxXNiOHZObjJjAYE0LQAbJOcJyWdfcqeVLTzGZtqb0vEejy1KyA1J3iT/rlKq
bvkQF70Ko1SdqBmMPMPajItUBYmgccFC2IsevDqGfy4ZEPoDj2dp/OTVaghbkugM
q+h9TsNgEhr0FdCd46rCYvMMjapDUFA5WJ0U/9YcPkXl1tK6pVd88eEdV9+lyXo6
eAhcZRX0KXbE1tBesOB7bnz4MMY9rz1FainTo6w3XnDcH5NCOoOKJEc8JTbsDWk8
z5BCfZAu5Ky5BIWF65tOwkMqFivYihyx6PlWPKY7KoStHv1ub/YZxjp9x2fW69wC
eANCm3OnyexvUtrHkfk5FmPg1+vsnwXC82E8HmLRbPa4hSxK6euB9tfTY14JL5dG
ajk4pj6t+Bgx1+GjDnJKLnsGsngFM1EtlD7A5nhrtj1E3w1yJyjwUc78jwPgzJlT
0JdHIkGS9ZhnGjnUOx8fFWYH2LsdLWlQ2dyqkJ/qVyBJ42DiJHTiOuTtKeYBID40
NLAuG6uLijDK5K3oQzn2QXoe6WBm64oW/s11r/7zgoHCg+hENhMDka/C0rYvINf0
dZViUWMHKzWYWyrz3mLX/INbE/VJD2qIkPM4GShXY5/l7V52Eac3ukQjPJMksi/z
xabcqTpwT43rgJd1J0iiFKHlCgBcgRutIW2IHC1KLVZge6N9HFhfIGEqBsSzdHOj
LEQI2vGoIS2qg4lJ/iCKOmjR/RuNcwWXxCXEwAoupwvPPlGwp047iGJKokrNjfLl
46xKz8TvPDe5TNlwl9k9ZMqCShLlDS0J7jvM4KSRJHj2pdTyF+tdHpcSiEB4VO3t
ZuJkhHsiw8Gz8sRlthq15GLyhfKONcuc11xVB3+8R4xNfMyCgOGbe2mGYWlQv1Hb
y9cdb8+J3Mxfgp7LwVKIHpbXHS7PEF6ydoxfBcq+SchJ21WbNMSoQ/LYlPi3BKM1
DPHVBgwqsCZDSVQtDGCXP9NTJgBCDkiQoj4EWEd0srxkf7ObbfYsCvfrieHcLSax
y9L1wAR5FzOWTlyS0RQTh8oPu5yXtNLV/2ufK/aILF1FX9wvwjEFEH6ygkxFhX+6
xrCrIoxDbRLa5uI/ZMPVfcD2rt8Ljpdn0FVnPsuFmfcda+sBlUr2vX61170ynIg8
o46G6blIZ6diJK/5dfYbYgeotZvVbZDjl3rjAl87aoDL8M1BFfZ95RNq8QbNyjum
z+fuMgVsLRk43Nbc9dj4wtXHqhdQC1QVmCrs9ljwFgt6jGVYVyxRDumawNCW1cvh
5iQIyTZCWYsMVYE5u4XyUqUTV/cs1FjdkVBrxm7/suO0i3WAdHizdUB4cr0kOOvZ
FrLtgVzAjYFbPpIvQw0feqblbIycWn6NCnfpPde7PkMPlbikQlDFBliePG8tEUDN
VahrjKJQ/q6HdibxFSyRF7tUPpGDPKUbZa1MfS7UAOry1JBjFAWjdEhe8ozf7ZXZ
TSGhni9P/20HkG3PWYufLl59XXTvnHrWDf19ocZQpv43glqM0bmm93xT//1MdgYS
hEzl6MYUb3sVC0AuZ3wx9qNaEacRki2tbNfqFb/kVVF+PKbpJLlR3dK9prI9xoTX
ZcxUSiFHAUvrg22KvJ/jbZyOoYG1Tp5g+dSO+szM4IDYKNpQVqFdV8XRFH3hAdBl
fcJBvtRuyjtuqesMz/KuvC0iJgBCA9lYkvBhcA6pJj8ad3ZX6Li/U+Rv6yh0cvR2
sSVmasoc7lU8zqy3YPWpywAcfUKt0Jl33N7G8kkbkACQZz+2GLIwme29qGckkzqK
wYXKcQ9mHB9rejoAsofm4ecxO1DGQYR7c4QHBA1zzVXkS2eqWhdcF6x0xHpDYaXv
LcY1CqwbH1RUMuN7lwWeJdqUJ/+dKwqvLd85g7lK7q0TeOafRFWSXkAHgOH0dTZS
pkyrp+A734ovbk/pKeC80eH6vKzXmRnRtvomm06QYke+h81Gw9HECPMoMjR5eJw2
Ov2PxJTfhbzN++nerzFWxur6AhcZfhdvYEcDeH2sRA2+qv9sFOb7taKE/9wI/Dqc
o8P6yVoqimoLe4bcFCSIIjuQ5YHvuDmpvsdbw+F81w5KHm0OoCfDBLel4NPdKtV3
ka6tDovL/IFX90/iHnSUtY45cju9KmAOqms3aLeMx01G0m9NTvBdOE2XxrBoBWWQ
Z/M1imvMW5aR9o6aGSkwp6TtAsu1pYWUei5u2mPUMpQcKxKpuPTskSoRsvnKYRjx
CC8qpZZ6nH2MiBemRCl8T7MNnblcSvtlJOZ+pUq/YGokNpQxWZt4x7fYZa+p9Kvl
fQ/1LOmLbCW0KJz5MEJKsg9UB41njSDgLIt5zHbvVJjv2qvpuZZgbNamx3IEpdzu
WU8bEvlewCk0CmELsolYo1he/K+0d1MFs8fKBfeN98OW1JHBkUT+9aSaBKuwvOZd
5AaNvepKNrvzN3WKHY7qJ5W7tOJk20m/dLLdTQWJ+eHK2LhYguMMUWFdCx4EJYD7
I+qH2FT3+8n9Ng5kvWSpn0Npk/D90Le+DDVn377VPxUwTJEweWzy54VzxBfQtgGU
FA5o7pckSKs1dUKtW+cZfMU8czITvKvbiw3U5eG+Ncbxrl8eoDKbkser8tuZp3/f
Fmjdwt8w41yOpkcuiOOM+nZMHEN5C0v56e54VmqekP0PkwcBIgK8+MdSZU93fGyx
YfBC/bWlfpqwEhFezJHgPWbtlH9Op5dT5/2vULfCiETzPQsLa3Qhfd7S5YZt9Btb
8A1h6Z5zLay9DWb2H7NdNueTqnneSkbTDwZxyhXJTiU3asfUQJpoatKNhz+8tBPU
bU3WBicErVyKAnnZWVZ31vTqaLQEGcdL1u4lRMPypSba2xxmxIqsCcbVOGQM+ZuS
14a1eCRGsuOf4zAVFY9rhY5jA/fzqN+EHZXJomBx+ssqZzKk+9j2pQvEf8CQZ6+2
xK2Gu4Wa6eRxQREds7DhHn0NwavF8z7VPFIbqHJnkqz9/KrphUc7qhbo8Xew9ynb
S81dUAJ4rHECAWYULQs/A8z56lZTqQTVJA5yYNd0h7HF+D06m1T+kEcfS+AoG3PX
IG0PfWvBvXkRS1xIZOIb3xrbARdKp9r6HDoNMErWlT/zmqTZgh7QLDdF9kCeRhB4
/hBdgWzNCmTb5aC0YEaKJNfP/ZDxHkuaDsTRaZCyBz+Yd7SgJBO+9nIT+tPGcli+
RdVji/0v+HPAHyYTJHc2aZS7JcO5F0x4KzpAcgqDlmhW4WXYLsBwQ+7MSQQfvr6v
lSKKuiVF2UVPvBo+A9meuRIZ9yVbeVvB1ZC7GKxKw2KuRY67OpQof8r729jeSQIN
zyE+MRIn6En8HQtAYVZnPmjH/BOccBbjvVCFFGB7+5FCTMX55gHL4c7fQOVM6mie
9Wu/UmTDYrN+lRLhKP91qaijcprDr7lJpobidBuEv+xeYs/hGtOyolV272KRxUuq
tJDlwWafI/gprV/Nk/h9+ZMTnHM5Uff/ReudhT2e+mkDwt0QeixOqgBvn4Klm2zp
HawJcLvkyGgKJog1fNATS8LNht/YUzItadW0SBELRnFjg+cBEjzAVuVMxm2uq8ag
Nhwp46i35Sg8m1WOsE15tskBNRJl+2lzJa8YxLUxOd5yV/rJYgLGk5KrkRiSD+qU
7iBQ7zB785o/HKNnEKgGjbz/YGotEM0+a+5NpymVL8rLOqIj5YqEOT/HTV21/0Sb
fz2/Y+ucZ+rAkojz8/hI6UL8tUXHXmBGoJ0AfTtK1vTHxkdBf5qr6kWjWYevLgtk
NpbGO90MSsKPju8ZJO0mGI/a1u6ba31H1AGBYC1lWle+vh5riIlZZKb0O9r0vT0f
JukesVXBOLwp1M7fTREIeqGi7CuxRBK0qiLprEoKDRhITAd2HR7fNs7b7dXuGVXx
HvRHi3H1Yj683ra0fuJBEbMEZsNb6LJ679CqfQwAdPhKJawr1hMmOIhIO1lPrXXP
xfm4y40Sz6q4taYlRyRDRVZaIVBPBqqcXhT8Ph/LPdOSzk+fxqwekQ1JJGkVF/yP
WsEjt7hRIi5Yxw7FzMlsDXiMRqkBGQPd4kOu9ji9greLa2+vuQltTYPzDT5nMeW/
Q34L7DiC6SodNtL+l5DFkU3DBYo4VGZeqF+bklDneCdg7iOCZhSw3kvGmhjqB5/A
ipJJ2BcCKWroqLDWyKv/83d9exSJ4W6I5s15XBytg8mHB3ALhsKO85q/szlDCq5Q
D+Mihx8ZJeR2/yenr/PNqMVmFhTUe/LvFN3RA+vSXPU6HwY7E8bxUmGFJx4/R0PQ
WaGNuqrBteRdQxeummf9YlF+/WJHBOUbSJtmsK/WAfuGIu/AZgZqKgNRL54rEZwL
ffLyQjjgQ6zr5sZ6gsew/2ggiRc19WUYLYyswhez/GwDAwwRNYhsjvsN4cGNzVq1
tDyAZPI/bwQAeCk6sVD6Ax27x2UPplEPK4McpvpjjRD0E1mtHFYVDg6GoUTRwxDN
mfSq7aVZ6tJV2n9f8HT7O8PiWZCYqRNsYjDyX40xqnmAkzgMfOpmSgGtcSsghw8a
zquiga8kW3CDIFvEahsBnwaFC0eRoDB7wj0VmVaa+8XORou7byzFqcDBQ47EWPQn
Fee66L8E9+Cr3EwqIYzplRa1hsypzxz5+vw3syGsrWD4gJQNy2YottbD7Gyuvi6n
9P2xHcDAuDGCFuSWNJ7ks4NaW9WY5QvlsxVcbIPqAn4p8lX9VbVeJku90Dr5pAvh
J48b24iRr9ZNtjAhdzXAPSmfInbAKFkj17aw7EKzEUZU/licJB+OQtJpQ9Lev5v1
uLEoaKTx22RlwekIj5PGyxiSukI5YOvyPfwvWkjrfPmTKTcd29p94/59VlkNUkxl
byB347PTpnCMhhOISJjqmtUV/FJRTrlUoX+TbCeLQGTnKZIL+rtMigmLX3Dwk/Db
biAmRnfy+AEyOiUP7alZ9cH4UY0wVV6B6zFm4eEMlj3lNwNr+MpZ6bwuoT/rp3sL
7DaPs1NrCKnJizzhTY9YXBqIfYQIDh8L8Q51k1Uyrj83Aw/WfaU38G6yqvM8ebma
FrrFygHoxVny8f8eRuzOjoqWH/KFNbhr9fnhNuSirezxNarZW+fGmG0xpd30raRl
SOH4eJYhiaYbZpedjaCkPVCq6qklIDnWthjrsYJ7f66yJCrUPEkf0VSSRTf9BKO3
SvNfTNZygLkL258A1ZBCTqFR/os7p1jlzLe/wvjwaniV1HqTwN9qYQspuAFpMjLv
GR2YYRSSazIAFjQSI4HTi4yPxCunD+40BQfcIirWrHmDl5nGx4/GOWsv6es3lMl1
kCDIFmfOARxcu4N8x5jswIDCEHXMu8OqM7Zd2p3oylZu9ABgt1/1jFbfp30vEXus
EubZu2sRp96DUjIAF0eQofo0RrRdqG6/bEdjcrjreKqsXXNfDUjUZVxScvgRPahj
/l9MwV14qJI8/+P8jSk5REQ1l9+lBgSiXXUmIEScD/OMVHaFK5JCwNvhpWHuPpjL
kMIQ21UBylOJdVn4eZX1D7n/hrpqg0pX2DDJNA0qZG58llf2tQumNOSANF2uRL8W
ZfLuuQk3MjcKlK/98CYoDRNlKIgIFLoCIoF7A6GynWRqn1f9sYgUrXEI6jkZTRX9
u1qB4y7qpsWZaREy8XAqo6u8B6RNNtfYJzeHAKf/rLHSBEkOsI35PcyMCtMfjgYd
9SPrXAhpSltqV9D/zNKykW3w/X0RChDJJt4vwGfKkMg3MY9F1RzCChr2prDWUUkM
NaLN0M1F2pxuANmsod+PCBgjQMv1F/aZ5YwgEFa84cE9H7BbasFQH9UMXSIkCIjP
b9S4mZeHvWVYfpaYem/kRlYiHr+6kn35FsYG7lyGdTU035wyFUcnnn4cC/WGehFQ
ll20WblyuSNsGmrvrjRxUmdlkA/F7pDyJKUDJAv7lM7FzuD0CZjYdzOyjWe6pGRQ
rHH6T1FQ4+Rh+NpdMB9QR0TjkbuSylEtAkycCxMAxX9SfHBQfka/OChGQNXiBSMw
zDmirF476J+SyQaKHZc+f2fkomSNYxygM3UZFLgiRWZqUA8YPiFrmmQtweaLc+N7
UdT8bx0GBaoX+Zttg1YE5J4RykIe9SZqTNaI8y0mfomhHKe8FhsIBIw2fmrHAiGO
ZoMpAFxyjYzpl69QaY1h7MpAJEcZnSvQ032JqB+JPUz5x/AMcvJ+GoDa/zweEbMp
ZyPIh0SDs5Zqpp5MySJnUzTuHJT5sk980+zoTBlb6IOSV3dH+V+jsTIgrD5dZsKP
yLG5VR4j1+Da32OD8CV+1tE3crRMAJKfQ4NCyW9kBkBAhxmIxH0sLQjP/CyUxqVV
wI7oY3BmANMQWDZM9XYXTYFSzoZ5fom8dJod0sQ19NOE1EhyHV/mfBsNbN47M94j
7w42gSeWMDX9l/z3EvmCrBBuzqV9BA2ZoQQyYMXC+sgoC7VHI1zTtuHXJUSHYNXt
E2xSOVitX8Iylw6GFW3G5LzMQyU1tMOrBTkOnMHqbjriwduy/p1AniEilxxMvdNK
ug2CH0Q4KH+2322JZzjk6Auc+ZP62Bq/pvaT239+zlD6fsAGXBsagN6aM77VI78e
uFSQv17P4F4mRDZXCx5PAZG4qzgR+LdjCfSLTj1/R89Z2FMjjODnUzWkiYPK6Fvi
T+743Dpl07cIMwqzMxQxovXodWeqEufJxzYEiFw6fK6igDJq60+9P0EqmdohC46b
hzM6JfWznBZdIvvGmmT2QIhpIlfNEL4ksY3WL0wzaF4MaawtfdMElO0/EmbmPB6u
HuQGZX9dMqhmy7A35HI6M8+JbeA++1KcMfpnEWPuKyB2ICuVQTNq1QXBvh34H4el
AnFULkzCsftBg7aSZBy5fD5zYu2jK2fn4yQEWDlGju4A3UIW49aF7QzCzMcTMCBs
qIDtQfLy4jrzLkFDixtOBrE1EznQ3S/yt3N+HN/UeIe4dRtPkjCZUWIegH2VU9Lo
FSYiUHaNT0X16gZm6Z7yKWPmXhl/dsizNRezI/adX8IjVp2F2P24NJFZOZsSbiuL
Sdr1290lk5A8AMOSn1omyhajAuA11ZubWGZfd/T7IAEFdbL939Dy/e4/Xfcv4oC+
lEAeUoQGLtBrq2F+SYnRcGYfbiNLKSXusSSCKG5Ik6XFILwgQCFxd0SIzmkoUZVW
JQvrwG0v0vTz2SlV0x2PneWS7qrrC+iITNbA0AoKJ0ItxytlLgI2Nki9AN5Tdryt
yzd6d03s2wPGZOuEw8txy6d3cliKRJki5xn5/TODaB98ReImVCUQL7yzTr3+Se8+
BUJpZIcVqbbkawmu3i8T82B/zSD+CLInCgY+Tl0citgI0GmLoOqWF1iMS157Gl7b
S9JQKdWTW3nlG/H6QV327UOXkVfMFMkDcV3Fn7mcYCbPbTKfWy+magLynMF4rN1H
w1AbMi3Qx4pBhmOmUMHLHsxPL3FmWiZfUoLw81G2XYaAyzngNWsb71621qXUQdnM
UpXg1cLzG2cpEcl3nchWMS+JFggrldrwf7X5W/DFc/J6P8L7UujnDfIAFi+WGd+f
sdCjLYPo7SUDDq8EPvrH3l8iqwXiASzTamVFt0Lyd0KSoT5LmfRTpcpb6Sw0C7HN
R9kg0FYXetU4dlsLCKEwjQINeDgTwFauIQ0Y+fcv9tkszvshhhnuaHgbOm8xXAoB
dTUotmv1rN+VAFaLm2rP86qFvjqep0zdah8WllfTMSGaP4dV0xh6vj0CB17pJaJP
tW5NBf+LTvCBejAdvlYMtFWoBdM4LSsKNxDCDz5ChvL+ZJsDjztwe/+z9m0vLuyo
NURJ0LIWjcq1h1b5KB+oLxVXueTfBLZ0xlNMAvn8R8rKlQ8bz7BOgUYNMOKfYMNX
EmnSFIeK8/H4g29Npm+B7W4x8UX1Q515NCzQcFwmoVNg/1CMkHHOg2p8DvXvyb/q
NifRuBP1k6TsX39IBfzxPCWMyALT1AFalNAWEmA0qZoIbhAqPzXFjUrym7LsUbjo
i85NV2PIx+eypMDJVDMZhDpycIGae49A9dNEn8XGUmuQvN1PWOCZyhuIJOHqYplZ
7sba1W2wJJ7+bmXgoJ70zwMDTCGu3EyieZGdRjdoqIpsf0qbFLZrHSZFP8NZGkb/
lMBa7P1dNmWBuIl7BTTUVapXv1+STxQb0seSykXppyL3DucyjsSrncJ+9KGF0cnm
j/qgr1z4h2/GyEwENzaq2KwzwcwMcxZoqGMJs0l8s0EM2Q0hZ3q9oCYnmRN/bfqD
+gIWaCvICvstzsyIxLaY9WK2jYrQWOJv5AICWlqnqNRcrwE70UzKrRvn7tu1dJWF
SDV5ZQPuBkB68/3V5V76K4Qrmw1y/+l9ai0ysw7mM/naSt62S3GBRTABnowHakOd
3uuX1RLyblPAEKUwFuNLwEG1zf1E9HJfr/pCVskev52zDlhIC9IpSXZT0AGau0fa
Q9yhKM0/WA1jj9rrqC+X+XPm32omgAHbWTA42mOJ9jgb9EouwpIL6gPi90gjGN/l
HOC6CkxGZJ9fjQyjYJp/xpL5GjzYSjXn++0f/JL6n9oEWuNrjbeF4vEc6bssXv2R
Mcn1jQnMSOz2iSZpyNoix5TYBlt9c+K1z69xZpSns7Fz3Sk81d//alKOUXJZmlbA
1MJtNVEscjOrgQF4ZSB5gzpjgrTNmPU71ipwCFn6nDyCCjurEHEj/CTO37CmAj1J
N38qk6Ah3o4f4+z0veXlMQ+EvqzFh7CLjJ6m2yWJltYqgqTXCNT7lQzI1OrIaJx3
8WY6cA3I9/BfJuQ50eHZ4S3P/LTxo2AxEOJxJslb7UiybqVNpmiwsECMAuuao/uV
fxA5c/zcyvw2ggB0YABgRnxURlBrXSo9TLFz00FAWvo0t1Wf+lq3VXHoQJ45corl
oeY2FhD7Ba6rikjaA7r4so3B8LzfabDZGDWJisdD3KAe208L1YKjsMHZ+U0BWyzq
TS30gaiMDEBsKmZhGhO4fsVfCz3MbXb8u3xsNOX46skFjIRDlCcvwHy/xaCzr3O8
IqtlmN47QZeq1PfTP2AkUQgiovgIqcHUXx48HKneocaJIj+52v3eC2IeoAjsj9Ix
BMZjKAjHJkQhQZ6z+lev32Qk5scb6/D3quYNa8Owk6fBsMEQdDGtFHKsjMm8Gbv1
GOxeJtSOF/Pow6bb9As2DotiM0YDFSzS4acNCZMCGs3+vLRyxT4Fr7B2HOLeYbgQ
rYNV6schcct7Zi4bURMS4PdYijVAOk6zlsx3D2H215XbH6TknChr6e12FE3jdOpd
ZpD8e+JBNeZIiaVpCDraIBtsDjIb/XmweyhiQNGXVh3mqfHhkP3mnMKUpAvHsF8O
VJP4v/PmRVShv6EOratVEe4sIhxrOr1ZanCBcpg4ytQzd5tCMc5dYgyHqoVsTmMK
9A3lw5jXfNm74R9HONNMOhaZ6YvsBsJc+s1CDWpZjR9sPnQwLVnbKVWOIyus6m+f
ItMRm0+cG1cJVJs7rmoznBvtuQ6d4LGIEPnLxVKaK5pta0JHuquuINiVUjxKM6mD
/pBhKkzPCFoipGUIQ0mKI9kBfvhe0tS4BeMC8yCyNPgzzd0DSo0HwsqA6MmKxOFN
R+4HbZPN/0/OAh8ibnN71WMWRHEbDw8fcgnBznVQ9h68Dzv7fJWUeu+RvHXazKCg
Dxy4pDT80F2zgLO3yp8X2WRFl+lZGSbwbbZ6Xfm4TdyyAiI+7D3XTNaauzpYwCbF
Cf7tDivvaJzHJRWSIAGV4SVcyC32OcG7fSNjYJvvg27nBjEvn6rOwHmda0F5jG2C
utYluOOmQyVffNRb4txXozTd5PKl3LhfV+qy+jWLCimdEAWZGC4Q4CKDd+/ldLZ5
Zg4MtoOkSuFPOuAEKurIb5b5ePATHKsi8JbRutiCRQ9dW/LdNotuGdxl/zbcitxy
at73KGJ82Al0rtdrvfDIWuVZR+WJQRKrS8aIk7J74Y1y5edgTI5NlY9YLjVaSBD2
M8Hjr3KCRRsQ2l/3KIzzAOyMMOvA26ZxcQNtG+hhe0hYIBSDmxQwVukPKApJMWZw
Wof5VisK7jT/xXPAHFXOUgODTFVv8CGlYMHRMn7fxGWqF88/pehscZVCuiqHWABn
uSajtAG4tuT/5b6xMUJnQOG6Od58pIXKxvEqiikM1DApvdRMSkkjDVGiSqIeji2B
znfSLpBXZoHSNeaFMOG4PKWrBZ1Az6CGk/0C7XUntZ682B23S3AjbT6kyqgAP0dZ
hW14j9VklttGa1Jc5asa3VjNPSC3H8UeUgFykSLPUmCwxIJ8r/ksN4HrmVLAOZpD
TiYFtoquysED4t3ViCEx1V8wnpjuPVyjAdouOcP1zLYwIYSdOs7LLwlnGlJ3kc9d
qP9cANs4kaBaAs2cRnsJxOeecnWEakOu6aov76t93Bq6EgA4RFI3O7hzQiFfzL+F
x7tAUHk/irRjYNhkrC36+FzaFzLi3APyyn60BJfTUIMtl4wM4Lv6OV9fR2h/0yAN
t9hNe4PtSyiO3JpPhtbYR3RzwCy3lzgCtvjf7JL+PUxijygHPZfTgocdBn4zTzLR
E7pGFjuguWKYkY+8GdNhaSr7ZJrwvnJVbaPzlG2i9Q0Y76H6phHf94Kriu1HcG7c
aVNXStfacsTJibYTqtp6aoc8qUpXZSkkXs1gNcGs8gbeSh/ZoolLxJVSdmLlc/0l
4vB41qQVfCcwbaNacPaMw6zJ9zpooNUR8BD/RDV89KiAYTR08M36hc+QMIItwmFB
awM8Lz1oCrB06KSzwpXVzNB3Ha6rAoaAfpuJvgiZNnhlUFsRuqi85l4U2f5I0DwR
sB0aaC+cVraN1i/T86Y3NMEUTdtFVI/yrUtP2lZYehMAd6rTZNHIZhCBajjBdjCE
NwcBG4s9SrSOxnuBBlGMzmy8NfwSGqMWkHW1mmSsRQP2lA4DN/3Z2KIHyfCDJUWu
Dv8wlVyITWFNT7+r5+5WC7yHwKcUuIJ6J2rePtId18Zutqp7cAQn6Hawtghnj2/d
YhxjK8Yq4sxUiKyFHHIO8A9eMV3rVAdQ4ISDFElC3UwT3d+6yJDMwaRJTEE2TEV0
Gf7h7smUiQaSw/mIdSibSQNKQDoACBnZ/LJv4toce8fHyEdQAFeuTN+jZjGMie5G
NNxVJaDOdam/DJgfWCttHXiU3TpuQ7jUEt14m8V/AQ5KNfUqBYKf7b1igcuLg4IN
Koxy/jRUGrPWP/EqgItnfVrBy2gfQYPyILuhzWDGXDR9aMarieqHQxfOtuKR7Zi5
EluCu7iCkRcEW/UFsHp1os2hoM3xF2sZ5akR76SP3/9p9lnl+nqKtQnu516u/rsY
55kS1Zfkr/l0sXiqLSpXtVbPj6DOCQE7amb/aFtx0u1fPnFCiGXn6VMZws8r0l0a
+eAHcSUJSalMhN2vlicP+SqIGu+0qbOFjdlSvllv3VgfvGoVAS49GyYVKLGQ/F7A
cUCreog806IOWPZTT6Arb9Qurc1ItmGldBFxpYNIB6SE6DrXkQXl+kB8rhrpKeLX
D8cak26rnZI4fp5hEKQ+VN1q7TIfgO03I0rlimmsOLzAZNsKuyjcwrNPAGW5q8x4
nCKNDd8iwD7qYPyXzPlfPyOO9ztOBl2Q3gmYTtKWPxc3i5zWl6Ss+1VsqMQo6h01
HOYzj9chZ9ScR/qhMg7vHv6DuMF5X2GSHP1ZDTttWRvsAIDTj26QwO1ZeN23XHlD
LnUOftzZTp1UjJovyf3dLY29mD3hVtlnzd5hz4361myXWkA4MIAbF9iDmntj0R6J
hoZQY2moUgV2nCtUCSh2CDAsVt3KJ/GvIBKAqG8K0CuUUV1PDPGgBn5xXmdnmjHw
D5aWNe+UETFF3NPaJjq55yb2v/uhkIZLOS4Pc8RBE9WRmel6s499Kxqqbu+NFC0f
u8RpDoPHs4bFZcHQVNiKSdMB03rDDbiU0Am7tIHvGVGHBxUoEWsZesL2pnD5Pz4d
BuqfIVzdM3jc4DLuLzkpMCsjLpGY2rSrhL2RGZX0rgOi3oZIn8saEtOlIFZZ27ht
TxkQYyl+zIDU8h0t347trqlts4F0O8ug4W6eN6CZdZBmSvFbbrujE+Z24IdTTcTO
ea8LSIvvfnphPcRSw244S7ntz77lDSwd5FgZLodD7jZv3x0isia9pcoKa+yQNlkK
0U2r4CnN+5QPzDA0wLwq/HSAe/kijqyKP6GPebPRVqwpI9vSUjowFjAeIIUZ+G7H
SBX01LDjiVHwU9Z0OzXc3YTQ445EsP4La1bjT5ZcK6rKMuCurq6KApDHwZtPBcl5
YePrITuBynpahMOiTz/tEV3AOeHfIxl85GwqNKnjsr081/fmT62j8ZvhhjXtEIKd
VWGHCHpCDZpr63UkRZNj80/fNe2s3vxs98EfM/2YH0GN5bPtolSGf11Ly8yK/tYU
nQQWljW3P8FqYLoCn+BwwQbWhwnvx8xyEhRvdgoW48B8SA03ECAqz9sjiNKu7vhA
h7SLFqzoefZHa+8cuvmaJjCWcVYPU45RfAHmxCQ0hmKBpPPgCsYxJHyipeb2pqv+
T5oBGdz8BqlQoeMXH/MJv5s2D/GF6luD4yYd9Y+dDRoZjxDUUgnh1Xkv3IWvopc9
nXqvFrWLbmqe4RiwKgJrFrrIv/FA6u3XEPSwYzbhDzwQ946dNeDQ/OuxrbtL2wRw
VPM6Q+tn0nADYFeglgm7gurEqGaBE2x8e1dnk7N1iIyGEThyS1g2cqhVMnt8F1MA
sMUqzzbt4071Cg5LwgLecM8kSTs62AdjDWR/lSnvyGM3NhdVgi1bjE/a6XOaIYMJ
qgyR1wb3UK2iytSf0BKecxkPXnJzNU9SHfPE6GZ/Ip+mFGT41DCLcfRx026TQVAQ
VHbGFa4ashBg4ucuZHZxK1VFse+r99lU8UQNqIdpYsRtusIO9r9dbLMYbAJftqww
o68b27oAI2nc9YKaR9sD8dUoygVS3G14qanpKXMjx13ty4IFT7H9LGneu6T3CY5O
SCVuhF5qn/QYCdBuHudZ03AGdVS/2VTTIWVaHppDdjs9iux5BDHsHpZnlDvYcWqp
3dZdos7uH59wfMRirL5YvDHJ3nzflvAH6lAH1USc2wCJyAleAJk5qQb56NR5nYeQ
KBtION+fLs6BjUJlc72DvsL3RYtSVSbudpOqeipxKMgQ1haO49Xvmf+2amwYWX28
WKKpGONQ/GG1nVYBTaXzb2FDCSTV1O7iQnBObiLsHq3yUFA7GKVTxdbNEVc1UMXl
fyk1XUnaECiCc6dpzhTDaQ07sGSXRWRl+xAUWN/dGKoT4JWvPNE8bxx7zSLe+DIJ
tX4fW5sqykhLh4h++mhNtb+8b4SyjZHGOinLyIBVCG8DsFMrZo29sO0gIJjOVqgK
IhrX2OTXIYSeErDBFiUWJ1xNi+rZ/wUoJSCJFF/Dej5T5vFwtPmTRMaKuGKCPZkM
n68FwVkXpHGGeER7DKdB2Up40Okplhcmhj4yuiFUVJ0PtYahI+aYvqWg4RI/yfeb
aqShmjVUpJ1k+p6J/hEtGRpSNaeXR68nUoHvop58CxOlWIq8nt6FeYBrWJeaIv4N
o7RRrgJI6dJygxThf9y+MC12WWmdDyFqOrMKRDFFoBUgXQ394mNI0T23Z+41Xmh1
j9Mm1ZWGpPRlqXVVagBM9txehQ2A1W+envsmlyRyD7AeyZBfmS8S3wALs+IAD0Vm
TIhxBJbI++LtxNWgdFFihbwmpQt4IlL4S6lWcQMQ0oa2hoz/PaRiBzVsmvsH3/Lm
XuxbWeB4Olk12gEB8LpD2NF4fYZVuQ0FgRejkDZbUgO0HNKm6AT/iYieyARp9RzP
A/i/rip/jfvZAhBnkADcDzJyzGWeJQxwFSlXM9bUFGA+kLsJiKg1/1Yg8agsBK17
Mt6DzgEj5xiGzHFoRsYCmQWWQVbTBcYAsVKtr2o8RtBNeW4XaS82MiX6SmLhQRuZ
71t6h2QS0R6sd4kFAiz63dZRduTHULruWtA233dcJaA00ydPGKaB3PG5Njm8IgN6
gbVSjyKcuZRu9X5WNAQJfzKEk+LfojHztDq6EaHydvRtzZr87DrdfOrEDQsV3EBG
9fJ75wmfTDSgk5d0pl1JPuYfnZZoq+N4sLhYCzL/2zgtUKwCt+AE+7eXEkxxytxu
PCIcESRsCRkHoVNHWcx/PUCxhjmlXV2dmCkEfyHdwJs8jtrX495KjmRlUpONcxHd
ZwQ7nXwXy5G87k8gqL/zAt0firzifOZD3KgWNoafJWyT7P5PwuozutobhO8VMDf4
nTxpnGpW9SBTC9Cu+FamJzqAPg4BEAZOM0nZDYLj79rSyrNmr1RjrOtZtUdi3W8Q
FJRbSiIeXkQ8lA6m41eMKr5OLgyKLel3/bV/v3daZ6+hzWhYY0+RXLVKAGHp+dxd
/Wy/YmYbOyVj3T7eWXkrhqHO4YRgvpxKzRJJ+331+dSxlMybB3jATXR82sPI4uA5
Cbrgf9IE98T4poxs+bdEKLtkw5C/HbkDbVDn80dup7oKWhkIKjQDKbkoEhNSrTVS
DTb6Qn0EFbgZOt/De/COQOvlETaqc3H7HQ2Om009DtiPJpubNWTtVBDvRSMTLfGS
K8tC6a4vRkHvidokCZxYuTvxUmkASI0qP26z5ae/O0aO1heZMC0JY4Du8WN2emGA
NuM8iVAdmZT3+H1M1tOUB8hZwf+J6PtqaozrA5UkRkg/OYSxqPmPZjGyGCbiM2nG
ygek8e5gP2Zj9N4yuoTUGvcch/61tsVR/6cYlBTssbU8UcAp8mchRGkAZ846ZARD
WC0R8HRtqvSajfMF8pjUpTH/aDSTq7zHDeBT57bm9LI4aMyA3aZn0TRAcQwT4kVu
QqIBdS1Z/ODyAuUCYBShk2NkmOU8Q67QU3Cogiv7g1jvr4S1GHEb3gPJNOJoSVF7
hbWYJFsy3BGCBWDk1rfjxMypoX2cf6M6opxXIqf9ZpnHy83s/qe8L+zsQolJUvZx
UXg2hy7wIAKSvJpQYfKO7MtsjCCL9pH6oDU5u2n3N5tCBLu9ZIeUW1pJvtmyjyo4
JEYFvXMKrcw383NpWICixCygq6V5JhJfnSQctnRIubQRE/C2YT5N1/qH4CotXaOT
iNFOuZ+79TV2dJog4rUJnqVBHTslaAjD3fSL8++kQ4DnjF5vVo7+WLvxF3Ga5mne
932Ia3yK1mYYwFDW8gk8lK963zQPNVNKpkgP+5SxZkUkDIbgBcO1f00qLFP9TLIJ
DgsG2MrQh1kzduIep2hQFWzP8sWkbKO+1DL5Sk+qt+youjGlkVxWuwahGWG3pG9i
8pxaENY0Zyl0AmUQRyy/bmuiukoq6XNmWYAXEZ3fGN1YUSGKuoZz0+U0F0t+V5pf
8O66vEoirJ6fa5xNOx8SgPVL/xl785AcUWLANnmrprUyGmUV+nnG5iumQZfAiI+P
d+YGhQR6uIJalE2Fb8yadnEmR4XYeFmKjhMIHSITk4tnIK7nsrYfQgXpZApmh903
H4+cxtLi73n1DWxV03mIy16sGB1Rx451L7eJ0wOe21n+x8OvE9rNHCj8DAkEPNV2
b882BIfLuN4R7/x1ucF8ISRPLF9cXHG1oRsdwkzzEvJO4Rn8wZVgG2+lNLOvsQ5h
leuZZ+QQRJwbDLXz1HUxHsCEZxQbtHnunHrLgJFloTjoGz2+260mL8DdX86rR0hB
n7bpXa0fdT31CCRC5H4ixU3tmq0nZPB+Zk1pa0KpLQcG8c8VZpOtzR6XvBxjdPvQ
THKW9cB1nTpjKTd8MCLih2Mt3FJlx/2m0TOINet2XhGDOfQ2Pnjq2pC/pLMhBmbY
fdvZFOrSY7E7w+IUUBBuqt/rUpYMY8kCKvbTni3p5zcMlnL4yKN+7AHW9E+3RtpR
ncEdyV5hWxnOJ68QIThzubeZpAVla2+PFS7b1lZGlB1Vw+lO3s+hTiK1/uh4rRkW
iDkpeWEMXa1jNKxrZv6favNZnJMt4L9Aq6Uv64iIeH/RM0XLEA5cEbQ520TI/zHa
EH1K9xPmAls/H+83JATGB9O9fkPJ8nzJRFjkR2a+YA8foNIEoiSzHm73WJiH851I
DK5+gTmvaYJFV3OitxX+0gNeLwfmFU+MBjo1UHAuinipBFJV6PAAoq0TL5yr03r0
k11N8MZqppPaMQW0PF+hXNLChz9d2mpnf2d0k4LF7sbXKz3w9dY/HfMWWnXEnuQ3
wV6iGpRW79o+qghUTZbjxftCu4CeS+KzyT4gKLl4dcTKRyLHWG1cSHHXgMUuaY2Y
2xRzaHR0GGlUApzoyVzRiyCbr0olGTfj4xhrd0ooxjzjvqTbr30uvDg2VynaM/W9
l0bu8gkjNhkUoctKLz+ZLkzkb+HXepg+lupnJ5cRjWBwCMbAAjuKP+lCf37/uoam
R7LuNHvMxFa3nbO3eJ2AamIZdBcCz1klCXnHeZaNrT4CiJSW99YbGoznMfrSE1pr
ZKbRwCmIIDYTslArFHpFsmsJZjcruRc38rfmUC0Ibf8oaCYqUmoGo7lox4bSBE6j
JYLFRE7+mdXI2bnGwGvmJPmoj3+7rd6JsmJyE2ltO9/AN9O0wU0Jgm9KrGl6mD9p
6Dm90wzZSG/y8C7LmSRc4q2hjkxb62EkH+QPMPeyHdgKn1DH68S+49aUlSKkqERY
SKBe+/uuGsvV7bjStKMSFSzmsWxaH6LFZUHPoHoOd0DbfP0b21A/Jz+gW2Gl7/Gv
guPJYmgL4z9JZ+b/paN8D8d3I/h+jZKceq2sHSBneS1UzWF0zuVyWMN7Oqxvhl3p
VLReimhZvy3f9Z34MBgB72joYHIsqTdUuY0+hBjMtHOz+CfNq+19ajdDT2Rum+uA
yr96Ine/AuaWKinB44bUw7vjf/JTC2Nl084hjejFiz8tac4a9TfWSffRgpw+Ha7E
2uKfZV/y3bhDlhSK3xjz10f8Zcon0ANXKHbbyM+YpUg8gWQy3hDsK5Gh+15Ur/wc
wy+AIYMixSGblYCwf2flulR82/6shw1dgtukjDsuGK2f0s0Ztmlfu90b1wP8uak2
MwQVxlp2rmhV5pYCgkrbX01CVUn2dGHae2XBjdrvIfo0OvBHHK7AFhieU94jyvx7
38mlyh3IaAZ9yYpCKPkLoqerADSzrskaQGd+CjjcNB2hDZFW7LKPTW/YPTw7CRPj
GInBegnW5z/ywxcxKRNk364Y2zuk69fRMLEBgVYDbdcYEomXftpKr1hjeHmRsjZv
6MAjnEGqcYp+7ltc2P7Em2+x/cQaKKRheOWhQCMaP7hQAEq/jq1klVx+UPHQuKC/
xz3yQ8qtWx8O+7iY4SHMmDTXwaywe8NNxNW6lJwF8oWSLvAMml/czqwDhKsUD1mZ
ybzlZ2rad9xfW6hKjV4TJNDiNPAeIAEKUBwm0jrl8afFUR3xt4+G8Dcvx71zScYN
hWx9IrUAh4mdlt3G0fV+rXv8/r93u8njXf14+vRxybrGXQNLe0zKpcpXA2yuXOZx
btuYW4CEgXZDduwjGdN+gW+mnNgjO71VvSS6ClFxdKaBWRVOgxKDzLmJ3FXiKpCn
UtXYTugTyEcvZUfhFVRciwGXIokB4QSOR28zJjt+eaR/8I5hWbMkeQFfjjyWNnF4
/5vbJ7ROZ4z0BWc+ZuVmvtXYOX+SWZgAtz9zgTjsXJgX4+0car4GEumAndGZPuNy
zxDbo66p5duhgWI92U5+E1wG8hCEWxwm21iIbJoMDSb5Vd2zvKd0j65//D25EEM1
VFVnjH05SPTd6hBmlc9ikztHyj79nVsGxcPTYe4d86wAJfXRGCygw3UXy6d/iUUO
sZO1X3/ErspzYh4J/NtYra/P3TaXmpZpGZthAljb2/vmlyNekwBRFL+fV2BWcpBj
/TI9BT09tFxmaB5CeQdeaA5eD9c+oeMv6CuWPOdJIuJLMouGViEcApQKIm6gjMpK
UK1sBRBHQM6irroJGzOd97JHrdk3HnIeaENPVHA009Cd8TBqD9c7ddy8cAGkQjYT
qNK9pyzugsDM+sA5tcy+YzM9/t1VYpFAbvYnpS7NWkna0LlwhcBe92TWOBKxfOSm
VM3lsxwVLdWGHC+LqjWJNiJZLHbL/isgV/8yOCnHwsPfr9xpBdHLirBFku/hUQV7
XIj9E8FNA0PIFiAf71hqPQFz+MmEWzAxg7qGAwKkgURq4iHUgDYphyb4Yx1Svcf6
uC1H3IolQS13yWIG94Nx/8jLed7zCT5qGOC+0syaue9OYQdHeEj/al/fRnBC/vYC
xoFhXUzRYEdfLNROIVHpKj4WxpD8kceoF6T+kKt+QFQaQidRPF1II8LhAywrLCwx
8iwxXq/ULWv5NSAjx4uw3lndeQfxbkAMxorHaqiBIJWmdeeFBSIUF9DslDIirACF
fi+8stVW14clQsuSyARroei81oFsnG0OTp1Z3HfH0w8m+3GS7lPDN5nRx/F2jNmy
djqtv47UuFESE3Rp+YRdiSJamQai2y+egOLRCCN+12akWTNW/u1WNk2IrFKTW2Xy
L82pqSOlu249RGb5gTqJFjTfeGcTwZ6cDABq2gVElhfkowyAJcKknRaCaxhPqzGu
vHzgk4JRgAqyM2sl5U5f3tgJ+foyg88Nsn1RIcyf7SejAq6RhC2Yd/rfKnNraziP
UoRv8MdbKhkUzwjDmhlNkO20VbmVg5rxYqfOtnaEaiMNyVfCbUl59yHZeku6t1KS
lriUcD3mE9SHVChCn8ZgMDOnNkwD5BClLjk2N+CzIqhHyN4Mq1SQMxv0y3x4rpiA
pFIgfUmMRbmuQ2pOQqsFu1j0h5WLSCSzMn8obpq55kAvXba/iKmyBxf50iATCanP
m4JfgZmJ+lryXHorV1gUwRnCtIMTIxRLaIhC6QOJCETmsfwY/7+hUCHmDWpoGcaX
g+z+a3K7npH0JYEtupA+R3LlAPUqsElWPcjthm5Kf44cAnoC9WiHTtEbekBEWPKS
Mgasqm3qxeF3DP+ClkWND5X5jcjFTnecvBi17PBAwvOShXWZ/dVLECOWv4pZljwO
paeIBmS5mY5LlqLlY2x8FnjGq7H1m1KThx9E1uWrs9MovmKeRXl1fnPfhw2NuuLu
SWaNC3Bu+BtI8Agv4WqQj51H5Mnd9t7DXcXbuSU8qIZJpD0rzmoRs5pXN2iruBRM
qEEeJtBVtxZ1QWx9qiGsexxcRzSH+B+6C7BnlwZ5b0CFzHx0/tFVKcVikHlI6gTW
c4LNOUAwWxNfqVchwE77J5XX128KZPyb+7IaWfbz6qVemNe+uN3pqz7wR1fVySv0
HshN7CKx3x5TmU3JrFupUpik2PZ8TW50KhkaUFYbAiI7a5jdaKgpQAVegTQX8f6s
fm5DxW9qkjStJW9+XawVdq8Bq3kibotvD2eGszWVrqnfqr9/wc8zNtggsQeGPKZR
gpR8XzC/F2LM4c8saWPYo/0ZwNiQshrE9uyDSzyWMxvrUX871b+7Wd7tLroZvJY/
RswzacSsWiFES5hYvJRFiu4h1LSAhpiKWrUJEJk9LgdF7CSpQiKBBBQ7DBreswfH
Din0M7UZCNtLZXsi3G/1IEnt8PGBtilTBYai3dAfoZeM+JzmuN4NHim+f1PSBjqx
CcYkhyarAHKmkz/n2hL9dsNGD5Bhfzk20w/bM40O/QISGDXKvRvMwkseI9Oq9Wil
kmYuQ/mtutKie7DKMPKBGDxTm7xNd4rmncI7pLc3hAcV5jThsR4fpfpCyNoYp2vf
0LXqvDuz2hXct3An7XR9PIYOkq63iSoMx9mybInUxdWxMWnVGJNSUpfnKo4e7S0o
4O7/z44qInMdq0TNMh8ZECcAIDesL6pWulqKktkefJ5Ep8fu6hO3Phrp0UgHT1Vn
ZtVHD+RvwNfbmL9gqYX5sdfdBgt9ZRoNyLU4GZxUTcV3MUOiU6YAYKzX/mc+4PQ3
F3uBIIzOU2wspvt1IfPutWvNkBUPjwI8M8tpc4u0/FhvtLsT5TXPLhrKF30Mlqbj
gSHlzdo/9JropArLxyqb5jBVLepi0I0uI0mHaomQuljfhwrvfnfP1PiarKTMcP0x
PKNJBj1741Bkq/qWV2xVRUdipcEEkRZYsVKLZEjceQZ3ejPocRsJndKrZTdlRRqe
L9HpajMS2/knr5nXaQyc26uzezFAmS9+VJN7BHyG7V2fcT430UqKVrrS02CW1Jwl
olu1jy/x5BizwvEGkLfEhXilNTFZVVJ7nBNHF7l6/GUVJB4XZGxZqrVSvQVSmbVz
G7etguqWYM0aCZtETSMWkdJG0tlm9TFUVwYsdqsAznYx8glYuUyRscqSQSbuc9xB
KXhf3hYE/tnjtEb5L7YpRfVHSblsM4EKU35vyVYqILfK9S4KMFUEoG1tDm0Lkk2l
tQPsha5BN01Y723ykwBChN2Ra+FgueZpmNNNfcN6QFi6j62Lz0ULof/OcxQWBn1a
kpLFGomWGyfn+cBcSCoLBxklGTwuMW9zQgYR6OvoOKdu+gccdBpu92EnzBuCUUO6
+bLZ26Wr4zdo/ANUKxa0PPUHWtvxaTGfTdK8AZGwJC29+NMIlkoeRCww/yScx1Xl
mzWGL4DS9b7XPRm6uPWWSnebHhNI/Stn4gOxk4KvU9jyxQloNqPho4yFo0/WnrJQ
w+dBWIwdGV9x1TFMqTq7gRR79Hofd83Gl125Iaq8ulNhTbKgYWr7I9EbEHB2/QMn
5EAKcwhOcvtcxM1CxbzMEKzlOokwmoOBSKIWTlm10+w9YasWFzy4IetmEuwpVG2P
wOUUd2gWF4T8rHyldkBiQ87Kv+NeH4SyQnYX4F//peV06YMmD1hQeKvvSDsEKBGe
ZauyY3/Xe8jikG+uuVYnZl4YT+aDoDIbWtJAneN5qnvnkzBVWLtLFASvZgzSGSV8
j0CvHpCE/pjWk+KbJLG/j7sLDo1SXjNHYzOvm+iNPjx8HUCKXbReBnelIxBXBTSq
zxK6DGc6gA1ttE2w+Rjm5QMlq+gqU/kSQNNyLkd39Ijz6nyXAZ0rL55IuKnWXnkr
FTXZVPsDRVSkgeFYHg2gTFwEyzQ0uLkZrXeP/4Z7LAIOgPbDeXscKhvminQPSPkH
1j5BVtdcoWZZDtl9GRMZe47NXnWcqRS+cMcGclcG+aW4GuKajnkuvAG12pELFgts
JbUObK2U+eVxAQ4L8OzE5WXWA6Go7aTdXb68KJUjdW1khuou8eQCxvPxgY2iY/tg
URZXMwgLQDO8FKUwxW7RcCWJUo3FH62H0+z7HP7p7+vxzI6UoOUMDVxJD03jkoHk
/D9A+AoRz1qFYeMn2aVisfbSYbtsc6O1LApc+ElhkZSKofa+UorOWR2Fjq6YHBdw
QBpenHKpYXf8GVgfcwN6Mmf/uH2Q8QUQrfsVj4TEqeXG+FY6JkqDkaZ+ydvJkrwK
p+P8sTLjvFeRU9RatENudDx6ymgrC7CAYsoihdE5FW3KTV07dj9Vl79sMpEkRfhx
MZQe8LfXx9U2hMW5CHM+pBDZsCVir2eLH90mGc5M9SK7s1WkGGK37Rkdfw0ykvmX
FIhyFERpCBC+k2+y2bxlzje2aLbRTY8jJPNK5GPdp0bXv6yETld4OULAZ+IAwTym
3ILDCSHeNOK+y9t/GBZ/ZJ2iqiyNalICv13rVRGv/hy7wJMEELvZyiFOl1MybM1h
SYRQQpyrWCikUoYJcU4D1cYhBXC6+0eAiJqFseltpIHzRxiPnruXDuasc/CR4Dbw
KprWe/N65fEPE4gKzr9BLblgXS5lNifrXssunAj0c8BnQ/qQD1Xlq3r0Uwv37t9W
Uol5tAkQ6vjkIE7gpEmx0wyQ9BC4CjM7m4s9qRJFmPe9NOanTfsxDFy8IvZPRqqb
p8LJNXys7M/Ex0bdVbQv0+ho/w/RIia9u89Ny74mcm0A/cPaz3iHLWbORZSuChJ+
9QkShUu40sxquwJc8U5P0hKLxj6N/kDNe2RewGM5f4nvfuO0KAjYhuf3uZqepyi4
1MSaaQ8t7grdeu5XHVE8oYYT37/7FfmA0neLudzM3JLTJMvtofP/QD4GfFTcFSxF
fOoWpeajYrqjJ0jhr3BB6Z4kem6aYyuttMCvSpiwWHr40Lz8rzG5PKz2XHubbWUS
0DRokv1GiYN/UIkV1TKMMjk6uvRxWGxiNSOaO/hiKb05EwgIxpEpX8t1QHzys8x4
63SnleA/awGXnLAbVBTBDi2xBXkxFcqUnbYgIGFES1UgEESBJgdStxjmt2SPKbB2
BcUc1gCfcqNQygTQtExg83JUdDA1ILsgBeaGn8/g5K8EkgtwHoVgHD3dmoksCY5A
0YJXf0s47L1sOGDHzNsgwEm8voitDvBjCgQl3aAoWtLv9qfRoIqqG4WcflOXBQXl
EeWbePvtw/zOD15zffllW8OOCqLubZQcI++265naeCGpq0tY69iMx3g9o1rvKovp
Jrf6KWn6abjOLw+pkYT57BWiJ6O5FnPMwOerlqWKueI7EeWKSYD4pqNqF/yE4cGH
TUsbYfIogdgEZnRt06O9owQaR7/OnofnL01Mb987Qumo6gUiEYV1o7iNloZSkkYH
KGFLDZA2LZKVzJi2RA7BLmdha08OQs/N/6dqWbvFNn2NxlAvimmqk2gqJyqtFhoY
mVqSNeAip9z1U/f9FzAHkHevdy6qkBamKSS7jk2DOowK2LYlN119vN7G8aWQN26M
dmIDCFpE19Is3Ccc6KIOdFeQ3I8znPmTCIFkoBAfT6EFk0aLpCetWhPwvFGO6IzU
fJ6A8Vc7iKQQBkVJpb76nZ13mTyUObh4A6UYYFnd9tEf5apHiipW3M7u3KHsdSgC
uACCSE0MLnNPrVjm15vvSyCuygFNw6hmm9zHuLbYbUO9jU0ukpTOI93aGJT8uvGJ
C8w6Fj0SOy3e3Ehn5MfwV3wBhkbhcf1S6VPlXCKR5ogczLHgjTklL6yLwO6vYblX
L/4PKTo5WSj2fde1swjIlXwjydkAv8JONe7oUYWWGvra3ZCD4GCARZxC8JRDb8ya
jBS7XIl3y17cfnojfwhzwbFOMaR5k9Wkc8EBcNZZMQ5SZbs2khok8sybtiOlidc7
ro+NW81NhKZqV4EYzcfl5Q90ylK9jhm0meKJ/NmtWAsfZQREqcazfPcUR3xHfAlV
sbfXVlzFWBqPx0/ZaQhWQuAk6lKm5TwxpiOYwMx1ksflTeHF+iChg1sAHXQGYGuX
z3BO+tYRaIKzJx+IhrU4ga34dEnWl0VzUYAzql8W4sQoroitamekHya7EuDVApdG
reUE9HoO4v3znOSCFrQvz8YkEVhEdLVVdlLqKZKKA/d6S6HS5sMBhLLTGs+lMnhr
aXo0FWq84UphF+8u7sfF8sWZr0QTwS08rqHAm8xRGP8BI+ncTRd8AOeYSWsGthsm
gs8NqioP6mubhIxr5Azb6A5nDo00OMC2lUQf0suJLqKsQkeOlQM4NESy34r5U3c4
5+ZzUwWIFvhF4lSnhbgg4wHUoDzHAbQCBzw2VAbNHv1XzhbEXAbheLhMljzoa9/O
VzbvQvFqcadAz9WcN7n6ryZQKe3j9TP1n+VNjn+rzJNVLU0GvCcgok+bwrK08jBn
fvcjzzRZ7sj1R66u4CtmXEDaPnmNt+G/kn9cBhRSnmc58NI0IuFSRN9qoKYGvago
vBO6a6h+ADFLqvIH8otaa7CGSrNW4V6UNWYkoVYCsf2dAVbFDZ/Mtr6XCFfFVwJg
hHYyqef7tMBz4vYjzGkXeJtEaw74qmMB+PPcxArIlTKVf8OhDGkqLw3Mnr/lCFN7
5cvhaCd9hvDlFejouoyhzgwPNicSClxZwLLMUlOj7xhs0kgX0wOq+8Svoo66vV86
J/Qwh5kwedqTYiB0yAvn1JzJTeCVeL3QUy3wbWCtY+HSuHg6eqtIcd4LTKlj0Ph8
DmIf/NcjDRBKZH3OThcUWVrL0heywtg7BE64X9uWEfcu/pnfNTON1IMF2+KKsHob
9F8EIhvYQ+72VGyrNIrgnIh12kB4AfGqsJyZLZEPc3vrFJCkCMv4NX15eCQL2IT9
xPNddz8ZWNu4ZVdskUNQscw26rfJo9AyrJy+4dj0RwEL/usHxNbaw8MoXpkGflAK
lH3e8oLWEooiT9KkOYZ15+Slbr3j3jYRjOda0fK54K0pYu56iD59fNMowGlHGp63
Hmb3zYzK77tpKU0EpLO+7onUBNVc1+rbRr2ASIt0N5caAC5bMaZi3HgyUrLcVMxs
Q9/i+eDFQywKOy7WY/MBu3K2sSqUAidhDmfIp+BSPHbUKwPsrHVCu6qRuuFP+ONk
JvYLR51ox0WfhAedAJwffWU+zYXsBBQKsBh3ZyXDWxEEI21w1IlpURpJ0YbPg2/R
4xVV1xsyUBwq27jwIJBv3TB/pQOn4RGbVV7ZqOjaKQ+xmAO1/01D0bW7WEfaY3ax
KnAC9/HA9lKNl2dnBJIZ+WsPRb1oOwUM5n6/FfBJhEtAbl2PENiXEk8JwBGIOCau
pFtdOFbcJVyLb+nlSWSY5L4YklKqB2o9tIsSDWOx5XZp5yDB/wQE2UPegXe42i+J
s88W/cI62Cu8ftGp3KouhrAaS1C9tNx3fhDB3WXdK6FWdXysc+zYAXERzAl4y+Ua
Zkv+7Q9ZQHclLY3/4gIzhJUru/GfUm0u2DyzpHRj1IBOsucuea6waKqioJPAsJgB
6wQCCricdVL8FO32VMQAzqmXrer3+OwyPEVetXrh/Mx4PnedcqhmWhCAM7runEOZ
Ell85tdywEqOmTs5GzAWw9qSQNx9ceoCBH8no6eq4psWrHIz4wLn+gIXZIUccuNW
vAslySaBUDIHFaJeI4dgdEYw0myeVReARKnAf8saVpgyVTKR2QeF/H7ZdNomPcRk
0Gqzdj07aZH6IFiNii+cbZsGHeEh6soejkPGhLWup7CPOBJswv759OvIooKAALE8
FxAJ6fuvisLpmfL/Qdo0fnbFYpHr2SbiFM/Y+cUfpANs+ApeYjsoNGoz0tcEgsar
01U0rMv9Ei2DF1BwpMik3HBm9WU+pQ+xsW04/VfBglKsrHpYCRWfWB0e3BcoFKdV
EnvJFWkUgd7shswWz8DN6KvzP8h0kYbkptZsEdJpF+ZXjYSlSHRqnvG2gZBuoTbl
Wu7ej4s6l87dDUw/jVuDBRVq05IAE/35RWfqp19If5Fa/veiKTVrt/U3kzPyTsGk
xwFRnw4QagfnXBAAY3jOZJKyunyiev09p4tkwBstRw3i/ZgorLHttWF7SEy8qiaQ
BJxYCbgUCVszFUuTRC4TQcbYM4om87Xu4Mxgip3NhPvgSPx5O7jrkB+Pkhq8PonZ
zJic/zHF+FN7aLFe6z7m2zq9o09/59o1IZET7Hyt9NXL1ItrRqtahBbZ9HxOrAkZ
CNugOHqgcL1u88I00MCE4yTG0EmaYTQI/JWhukMOjgAQolAKsEPAUxgelVbYhH8T
N7k1nPqFJEv6gXEGAbxVvW84F4YpMr8mcFm/me4K5DshLfnHIFuvRGZSL7bUYz/1
gwVcY78/CEXsSgc+jzDk9tquYA9DbToKHB+CnvsZuDCzXPN1Kk5xWerPzQOwZZzN
RBZ0abIYWO6bdxAc2fQfHD1p4pJXO8ABAV4BSLu/+vdrmwC0nW/ppKuwShbotsx3
C2GVxZQqkpL/VBBDgMTUMjYIp++xAeNhaLQLa+JZ95bK895Beu0CSMdj66DK8V2+
Z+yCsjsCALYhmppPxsvNg9XWkm7I+rZtuHReoh6qkEC7JoVbvxcCCeukFI2VzQGL
MQsJj2cOUjQ/MvJU1rt66Nmh1uzTs0obqDlPH2Kh0w842L21GvoFyQWxwpSRPm/R
x/SNcCC9OFXXGg8b5mpm/J+/mItm3j4crjKOLGr3fdwLcBkP9W1rpX5t6/RCW9GP
a2RrW4oDdgUeEDRfUp3bm/gL2iD1jConK5wNdDfy1YgICzCRURWCovPPAaqyJjFz
I+VjM40QkBicUeRmF+IybALB4ZuncS+bO8SmIe82E1oPpUEiVQ9Z8v+nl4LNDWWm
vIA52kt9bPJ45iq/BqizO/x2GrzObdFRqGdJceXYe59/nn6PvL9fo2XXYO/AtPDY
SS/IkkB2U7lajqLQ9qWL/XzqpV0DD/oZ33RpXuJTTqwG7mmuTb3EGRAzWj/Bqzjr
ewxu1Z8Hr7EbWCrwjh05msNWUaFNVu+VEjvOKRf8RGiMpVJcL4hNZzbce8m0q5rI
ZcKL6YF7CKeJpBAFBkzpVruEml7lzeQ71SI9w/6Dm0GmFfeIOGRcBr3OT1hdaR3N
aR6UZAfHEe/ippAmQTp+wOTp5li785evsa/qROGZaeRrbp/h28fxZsGzJkCZ00Zq
KBtfjin/PVZllgXLFHsTA03/NX35X+zV4XxK4DZ9goUqcIMSUnwtB0NNO+liRsfC
MXRAAaLA7hRdngjqsAriIMCEkgLK0AdXFBGlwu2Ne216gP7x+8gFgoP4dgLtmTSf
NUSShar839dPrkz9scgawq/MdaLsX+zjes/KYeR5RZl7lrFH7vSh2XwaV5q4f9ap
3E/umHmOI2vbIZJcVxN6gFo6tHxrLOiq6WiSIbTU9o5bVpA65Zdr5fXz3tK3M3lx
Y3sgvKQu28TqDoTGMSndhqU1ml/DjzRS3CKNKyr4J5NFJAI1DcZX2tsuFQINExzW
1QLagY8anJDzprKSPxur1Ez3AtjIbEkoQbMFxbvhKe9luL7dFmVeAe351hFVJ0hx
Qd6wlCgD6rqgPS8edewbXLbq2IuRMMCoCkdd8b6TmBNgBDEL3TkmKC68EXB4o39s
6ZCfi6bzSdxOqX7Qc+Flx8JRnSB9s/nbcbbOXN2YKz8MwGwAS7fco250TfTHxvG/
lB89qKoM8LY7OH1uJt3Pijb8D7u1r+VIbWLPfD5AiTS96ONndzU9l9nKdJEZDcHF
/hmRwQPVgt3bUZ4KrRuOsLOMR4Dor2nfY9qGDDqiWMwbTM/Ouii9ZWTBRu+ntW4K
wpKSZhoHNLuTxzIndWEWXJlTnyvT8PiJOyoLcAjwhhc7kGIYDVuclk4rRhu6thzj
czmlXS/Oyd2k0tnJ8/s+I0Gd4ij2fgYSfS6KI6VkLlricE1TiPXGZ9U6TRVLvldT
3exMumCMiV2qFTgPOTiQjYCe3/zozihx6albJqY2MfOtU6/rBsAr4y+Fz9jvjf2k
r8LCJIMRY0HFkgx4iWuX59sLnybJ7jfJIj0wtz7GuDFJfulcImqJyILJRwwHCiq/
zG3fwwd158Bq8OqNMuDkgG3aOeTNaRjLOBMlepDfGVmCnWgjJ0l09pt9asSTk+es
H75MQFCG2o7VoDVXNlpoPJ7+dqtT27m25bvWddqO5aIvQgLTWhWsLSNf0szdjEYf
17/xqALXrngVFDRgY0WGT/cioBGI5h34B7h1R2/24Lh0PfyPGTDZj+DqVKneQTNA
skpS136ouT3ZMkyn9cow0OaazWO6AfT+0Qcg250pNZ+XdAMUyg1JEFHHFt1EVIzn
0OHx5RQ5lBJDHT8a0m2mG6y8kfHLDACbtv5Tx/Dl+hBTarwEi9zhH5es0pvvFpNV
jgXIVZ6SkmUEWTd8TATQ66gC6PBocjnxDpYjR9gBj1OpsQb5Ssn8k3thuPW8wXk8
24WYk2BuWjFgw6NzvKJyZLe1R2KMosuSfv65b8OiJuzXnXdiE4T5mOvul8ohcJo4
oCiJS0GMilL5/jHsxKqBvsruimfcTojHhhzwpUZNVgEyQMeKZyX1JRCmWjcb0ka7
DzVTcMBlJlnSkDGNcpkqIwEAtoUWnlWClLBlU3Q1vETewbBiGxu2kS7oDErROWj/
kbyzyyWCHKMn+BMuj8eRH3mrW/dOWXFjTKsWyTpCdZ3O74sNOQ6g51kxIgNO/k+m
86aD0LqQTl4JegBmJyN0ntQSQamqiXMIumd2uJkyhVR0FMNnC1NdNjXBKQt4h6tE
6e9B0RUH1EDMwTMfVPXVFytrYNF55MU/eZAtjCuszx8m2olG5YXRLfPxBP2649dG
LoB7voq46GKxAVfIK74K9qGJ8/pLItkhGNggGKuC8FwS1eI48uFZbcM+o+Clhw+1
LCCzD19t4k3sUYrj0oVWiJn9W6P0K6fvnDHB+2+txpFCw6H2zs7MKnzwLjYuNyjM
eT71Cvz4uxadR3NIIsAEocJsUlsk9RrUBqlcC13VvBquYe5sgkR9EEhBLjkWapJ9
1pD2PiANSHURuqirlxFuTId2UR5kYx+gF1ntnreGy2kLZzLjoZpzJfYKgskqtwEv
DH+oFXbJoyQoDVhMOFVkzI7HfooRBb2hPpDLgsf/YZW5jdNHFY0gKBqRDlY+NxQ2
t+CfM4R4Xg6Rl0HX3PmB9SswUL0qk6BW8oTH/HKFB9QVNecEAMpJxzB38i7nQIdy
qp5pPzIkGqx4MpEqtmX0gQ2odzf936gOGEdZFrsuf91ko2kLVSxnGC7g7uNgLyWc
2Ra9w5XRN6+3tM0QYDfCZ3647uU1KelSoyq5T0s3xQ7fjVhDhsQZ3SvID9KYYywa
7rvGzW7swNZmyidKNRt8GWhQFGv6MJGS2A/UVqxku31LXyGSEI8La11uEmEEg/7k
rsMRYc07F1O7z4DurTM8fVOxuH9SudfkpPTK/ddgH9FoXur95fnk2W0B5TYddG14
6X10WhY+BkKJvvilqIkJZXjK1ogvbZ15/Tyk0CcvAxnSofG3jffoxDIeF1Rgr21w
RGVh2U1UadQMr66f1jjFr4gLcQxgZSPPyY7bVMAX0+dnQ6nB0HHgM0BHPOIUOsvV
06OSVb2n0K8sLc6SSHW5w7Q8rDC4zBsFmktgdEoINYG8/Bmpkx9838tEQMRK7YJ8
rr95Z9XudeI68VRSMG/jlqfG6AM3WXY0re0imZXYJtqr1LOjYidD2FhKRcNyBoU1
jZ5yZpMF+xctjDJ5cqbyG3ns+52nO7A00DUYjYs+K33TonyUnz5frjvWhE1SKSL6
ubSZJTBSixaW8iDt7H9hKRVNYF9eLUhflHzCu87ANaBK2EHXYRGMaku5EvpjB8mM
cO4YWrMbrflWHxYGxSvRCoDTs7hh/PPwnys9uRXM9FbxMeYFqrFgoIz5mo4vk2D9
eeFTbfaufZlg6ZtstV24kEpl8LHR7slnuTsfwy4H3okY20yrC6juob1t8P7/YF2P
Aqli2DyreyfCcJUCKhcHFEgTUXNFRroiIMDdku6ls0HWG6XXWNI5iNWgvmE1jYbh
Rg+OjSL8Rufcc0A1KY2e62f9sSSmBL+sHk1n2APydxm38WQXkGLASNtnjDF/HrfC
nq7MhfeFuXnmlbxUBJ1zpCT3qrvDiPMvMY4/hSqch8DIcJnQySpI98rdZQ8X6HRX
NG7+tZ8j0jnpxO/wX/kt6cH9kIbNHXqtAEPT6DvNFvLP0L2ea+25n/FOMc6VtS94
yPK7ENGguCWWWO/zJcvlZlWqJBYMglTi6/0R7s+OFIJNq83beIivcTfRhIJUUuEO
FfNj1OOg8jKqIM/GWA/wWwMa3BMabD8UVwOoRQVCuBgwF9g9Nrg8l0YRI+9tSAvr
IuW9Pbjek9JlprOnIvlGEYcsL2H0HYqHol7dixjMtuh8Gimbpplg8fuOwj/PMkRc
7qzpcXub1f2I53Oda3O0cQGkRAhGqCN5aQxP3ZlSPlbuA70cO+sX7o28hIyOvJix
5Tb0chncv646bgtee8K8qvkti5Ew0qCByUnROBulWvKORJJ2JeSUo+LADVpTbFVP
ulfPKDiWItBdXlJ1fe+hkS7c0fpz3Q7ISWQfWqwx9AHFCh/5QPVS6h+y+fv2I6qJ
RR+fdLSvI2yK7xDwqUwmdR8naqZqKcNavV/f2VuSyVaCD/VSzVUvPYHt6kajiiN0
OWYUMzPO6jzs6KqJ4EfsZoXTk0u/PJoQGX/UCDAfj/7Ejcy+x9GYoOYlmrdvv6Ph
xKeXescuQI+Eldr3KRBiLURiFi76dsOKlS/GXz/MWKXXBT4dl+tlVHIBT51lB3jW
q4lOwBqEaYn8qWKS4B2rfxdbDiLcf7FolXhPG3HdlXlMvI5xMeXXUNjUnw4EGDTa
CEsoNbFO/53gkyVwn5gpJGrNwKtXKyuF0kGDMDF9sS0sDizmH2dTAUwQpT0i7z7M
1qTYPktxnOHqF6rOLVb9ewNN6rkvUcyfTCeoPvAeZmvG/NJfkaniF+G7CmUn/byQ
wb4UknpGNiXwu/v8cnkaOjIEgMzfYtDOSnt0+igznV2KpVrOEpNpgZx/UpPiLL/c
IzdHo3A6rLTJ3Fl4e443ZnQKj4JbR3f3gHkMASOH/cDG9sy2/3uHxzoFNnj8A/K7
SZ9IQ+99ww2FqzQw2O7+WGYPauif+/QELei3UmdiKu7XNxazeCUYoPc+keNl6I1j
U4oYWyiMe0Q/7KKPBl31AsaGXFHp7q3pgM1jxkbMO2l8IgUa9oUXIwAemZ/ZYWbg
F2oIDaN+glThPuANI8R2vs6WpWvLz13mpHbvh6ZTxOJ2lXoD+fC4TDW+0qda2/h3
RwJx1ZZXTYjjRWEuPpP/WQ1NqQb54wH2Yc2+qDKNT/COgBFiVhSs/fq2/ZztIcse
g1UPoYWELRm+aeaT5zh21Ne7IlP2yVKmrSFp/VvJ4az+AT8NowpIocV1OTUaMZ42
kuDsCt/p9Hnt6QooPOlWxMtRK8MxtD1EaHR+oHgaN1CDikGyD08UaNiM8vRroQI+
yXlYLz9chrfX/+fukMQZmHQegEmGUSnqymbWvRy6Tp8flttAFZjZHjY3f+x53OXw
46/dQ3RP3fAmri7N4sBEbCgcQNfPMMODfnGkDw9r67camgHjgmzrI8/mUqkgzKby
QFbcOgru7kpkzZBMH6iWwPEWv44/aCXIVoGjHa93GDrjrDj+Aei4LBHWyEyikNq+
IfOKdIIbf6T8lpTYtMOyz/OXqoh6/9jmVe8998Rrszw9ZpHU21gVnlpRZv11xV1L
60ZeE8VGxeDqge6/SzR+iqWKmYyeuCqyHDNtOphawXoQ6Szul2i11jTcJU37qm9L
epMUWMPSXWYdRGXYkAWQ8aufPxNJHlgOtYCHM0crQ+gxcnnhLlLAGuJmW/oaa0HL
3z5FpsVMUR18MJEimcaS1pH68hH+wfYkjWtV4IhOjSMEdjtylAjh/GvlsSIZ6Y9e
TEH6m1WcLtw14srv4+o321EFowfcV2kl0puLQpdqafJZXPopGjcQpVl0+be4ogJj
jloDu4XDPSr8FLdJKGRGwfY7Itd8GO7zZlbPppOktkTr1P4zYxXf+tfaJnqjelMH
8gXcuJJmD7fWF5RphJFky2LYqG17BWX8r4LKjkMEINNEQ50AsRhvyXWtArU99lq1
CF2JRk1qFrZjJ8Y7kyXTkHUIIWHx9+UhnuFziKdbCnqzMYqVadML/5RaTyfYmVPy
9wIfHHV7v19aqX8Hx9G+RWvimrILi7FOOcFaBfE3MpU54yR+FofULPF83D80HYc1
1UikTQhJnTLQhV/9fBNuiI4ZB3uE6bS//3iH/0vyJNPq/oulet3zM6B2ztNwXEup
lGO8PASd5LOiHsJ5H9bZNhiI3feb9uugMBvDzcxS80DikYYCdWQhavCERQ+hGgp/
DgYX4vfuV8Uc0tsrQdLXEv4CDahfU0ZjjXm5nBFhcTE8lgU/ntsti0YJxLThZmGe
YiBJa6HbuURUAK7+61nilC+3ViMfsL8xbgJI0kkaleFBK1bAzR6iaOu2eN77M8rQ
Hjn3BsQ1A6TQ3QunqO/obd1IjFLW3wglqeZ74G3tHaSqZpeyUyqvLXxbr9yG8prf
kkJpIs4hXWjKe4uiFrkcs+nPSIYOLTP/PJYD1tMOSLDmcwDbjF52OVd/q9UPIQVs
mDxDnvbcaLTBoqHZqfXfCGUzcNwAJeXHISD9X/f37ZlPTldCHjp4dJOMvsjvwMeA
uf/lJBlZ4rwe7pmTwl/ct4SKYk9YJpYFSAnPpRaoX0Qah5TQVGtXIi3dvheg8LNR
2bhyPb/bIBfd06/W0zQS8XWJN1cVlTpeslDe68bkb+XasyW4Hi1DhRMYMVjy11wc
aDy/bOWGEdBj1yZFHNyEQTBwXPy4P2CH55t+OGoCVmUQKdSDITHMzhMLE2VqH/8E
I5gxgGuNA3IBTJKsksYUSmX6f0pHFRtwNQYN/c9sMv1oOGji2cCL6sfAO9YqGnnK
iJqD11x8EU07WK5PkvsEIw8AflbtRAYZoV87pCglKf5BMLSlvbJLNQLfKUBCkvX6
V+R0WeKkJ+bl/kpB/JzYttPU16mH1i+tTxRERTBkWNQ6zAlwmhFjtIoXJo7yy3ho
51bdlbN8DBnn0SA2BKJTKtpWd1QqoNE5G1Da2TcR3jg6vbz1qZwHuXJxno98DcW0
oKeeBnfbEn6lZ7F0enGtPOV/d1tHNeiqcU69ZhKLbkKc+zIBfZpiJoXn/gOavofK
d743ksEZ6PKWMsgCkoZJkvHXaaA9szHg2GUv4nmeUuo+xF6g8XLrQjEY5C9V7lvI
zlAPELMp4EZDoTcgOIhqdk8MZqcj2Ia/xp1y7zVwqrCkyR1+BsDMSSgWeqCXBz+z
KyK+IhDoQN+3UmNYtd6BId72+G/1Yd7/RI437QV8zyaEMHiWi+AGGWtTV7vrOnhc
9Nb3ofQNpA6djmqmtNdB1vRLbu5BScC6emF1mwDIAqH1FH8y5CYTmq63j+14Ss0t
pWWc+16EPkb2FfA3dk+44P+m9/sZpdNwAbTcV6cWLVa6UahPk980eRx/sEca1Bia
s8QaEsbS3hcSLO4FNfbp6ynFJyuKMU4sJW0UfBxAIeVrWb1uSQGSgZIOdiSN7CLH
PtJa0WqSlLiX3QzjhP3Rui+I1sZeDia6Xw3buqhV9AK9RmdtYnz8xv4z61cGrywC
GgWMdrmGztr99q8g1c2ot23zjBinOQ1H+XbNLKb01bAV0TLOjrkO22eOg3R9CIf/
flDuoOuItF2hOnU+eMyhJk+b/gXj3a+a2mdAbYAm3nynqf4YgoMjVz4gJUzYTG7W
GyorqrEkcAiIed/M/SGXVzQJt35DmAODR3lCyXAtpMAhQqXN2wUTunVJ2mmwOh0l
hDPPssAWAkMApLpnMoeyDtvcAup7x6XT5F/Jkobn78SV0cByVOlsZERItr6MrgHC
RL2UNSUPOzQKj/T1sWVD1UfZdm1fNK8SCY1SPoYpF7kQDlkg7nQ0TgfBBB7bgQJ8
5XoTYmKk1a1w7Vjhl5CbqjOhSVegz89oXVRVf9XRoHU1imtvQ44QxAnYSp9boXTL
JBUjI6NYw2vP78dOPTRqPrpE2hGdGDiDk2eFf7f3j9GynJQDSAV0K+rWy3PWHMgh
EDh3h48jEEgtw6M0v9Z9PjNHkw/KZ5r2ARC2IQ5Er3gEwRDNrecUg8qkOs2GsulX
hZg3uV8aB5ss0j5N3nA2ynUV/vCadA5czAGpGCsI2dWEl4ezYZM2vhXTzoU8PzSY
aPM1zHbqJRy7Nod7luxlg3lVnZRQdck5SzNt2Tpj6CEY43qNTHizeISTsNOtTx5b
tuwCzO8RrNlcik/NeX4NbGHvajIl9mj4aHRXlYxJCxt8ImJecFMSLsR6uqRuuXfR
UyJkXGfobF+2cxEGf9VEiBD7AUe7UtWpAnPqlQK1DcJ1pPPh5TT8Av/GidQ++K7M
SMwBsizsnLPihslcI/7Ex6NPb3Lafy3iMm0nASzxsBsOiKobv1BsG1hIW4oCuJx7
/Z1d/fbcpLl+LYFsniqmgP4THIKw/To5XLdeT3X4UfDlhu7ByFZRsY7DubUZf02Y
PMp+qae2mzV8KNviUEsGHHw2rRMVsDsL3OqBNvw7Tt4umdTC6zMGSWh7cmmqnm6J
b9R4k7phzGs97vrODGL14R6ijqQxnbZg8pFtB7PNyDKuPe5lDlQTZE0eXhldnvlG
O8RaaqX9wezG7iVeykyfWSZrYK/ZkvwyajmI+4C07eh+KnhGG2TARtu/2vS+qOxk
cWAeWXQJyeJ2e6JUs7Pxw2JCfsIum8qtLakAqcwLyAr00Q1699b+2BdK1CKKTp5O
FXg+xFQuphUh0hlZASsSSU1Kcb3tfwFFQAblnB9W3ulpy3gC0wcZ3Od2CzuDHBlG
lBE8TlCrJ3WCvK+gBUYC6y78n4vQYsVd+0MWaCTWHhEbmBWb0MRtL7HI0bxIlMSn
RLtdVPM5rW0bxjunwdvPsTyBHNbsAs5mHum3POskMLLL5bp4YsY+ndYDxwKpOzvO
MOYDRRhVDJNj1bPXiKGMVjC85mmZNECN8yWwGvRoRPfmtdN5H5sPpgk3FnpBK+ij
PnrKZen50nbuzzJXZtY5R9BYwG1xzjySeHuzwq6jWtJc9QKKZuzYAVdz548JfkjS
WViX9+IT2DvNtENH99PjE4f72Pwiol9Fy2C7rxuVVInHfFn3xzUYnPtlELvpUF3A
vKvVBjaL/bb9tlFQXslT9Y02RZfvz3V3ZYJeiNqK9OR9cQvy+SCTncQ3mrtdjEcj
VJcPEzn9CXe3BweQZexy2cyK5iysb2BCpT2oufqN/nfgFixDh5WmdC48Rn7dI0Q8
dFvHip7fv5gtZvL368CBpvDtmlEzzdXS/atK3lIeh1v52SQHPjwbKZ4S+ip8gjkI
oCAvDwPsie/roGF2RbwN4lV0XOh1xD7qnzqM202Hqbu5J4jn6SoI9C1NawmREijY
amWSTWxKOSldj5+xUxxP1CPyXFhf8X5MeOpf3OmH53TbauUQKJWCkzLhHYvK2jXY
nCIX6RPzj0wxrb1de7ZrTPnZ/gWS6ik438iFkvwYlA4ti1JPbLIwv5SWwZpY0Kwy
iHDObWyJcgnonsoKUOGAzcGOFBPACsp9AmynRsX5HOlWNlH9E0UCtiNgKf9mvJpm
xa6AJARQFxRImpr9uWtNTBEluixW6XrLMuppuT8BBaLAS2iKH07EM0dMLCaxnB3m
ZcHG5GJuYIbkCRfevJYmiupcA9V+aj+k5YS8AZCdfetGTIVXnguohx1b63xNaGvd
BrbEhREiBYc0lYEcY0D6QFv4JQRfUUSFCU7zXrewOcZZzNFPdQ88MFOha4vAqFRv
jvGB/hKGYz9DgkpWbH6CZ7kiGdMXpzXwP0jTuiZLtVQ3ZG3SKzJOR1lpp3wcCx5N
Vw+g3QybUOX50qXdKRfvIw==
`pragma protect end_protected
