// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
M9pIPztXNc+yCRj+mnB0SoSco9FL9GALrcSCJwdit4z38EojVx4fOaKIIvn9P1Sy
JnAC2Tna00jaQne81F7hmCm4EQJd/6np3t3gdDkRTDRT6c4lgMIiiH+Yjr0+Y/kO
m+SGRUJD5917d+3U9wwK5kMXs4goWZXvi6jjqu6EtAQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3232)
AVYKgYmD6N4/mMsrlyna5bHLIqDTAAJXAMQtk4UaDStfrIhVQQEA0dT8YO+EyRlZ
Q+bpJ1oouz9eBVPM/ezb94+1aRS2PqXrtlwNhPINqP5d8FGK3lb48hR9A9eN7riF
VlazFO7jJWYKyEtAahWA0chPkTRffkTD5i1EX0MwLSTSBAJLETAOeCnESoKmsAqS
5w3fDPGRPJyjt7WMO8qNgcAvmNtaP1rAohkNuMCB1F9IlA8QAxhO4yXpQiRRTsjC
H4zJZtTGr4S6PIOGIcN1uLHLmgASUazZkSEqgrbfFGkbqH1gPELErNgYwsk1RXpJ
+10Mq8GT3euCZ4Jm65ycbuv5vyfmrjIxpbMKTjLCsyIL/lpctwwp6ahx6poRwZAo
rdoU5SpAt0hv3RWlZRfiWpw2w90yjlmCK/3Rti6X4oCeAHG5Bfyg17KRIACh7APx
w4b1re/wi/+mekEK9rhAeEGs0J1/SXfT2kx14+4w0Zn37MsznXGsgAVoZfcASR13
W+W9EzEuG+SNcsG1kOJGED3Wg91tOxgk5wQKj9BPI8j9oKsDeTaWvM01PRCSPieW
PoXvetQUZhYXnB7kDyfqUxALcjZF9zZkAnHkxf3pi1moqe4cbvbd1SNkV/SKabDW
C/KuTDm39FjfZCjIByTw28wENOYPnpK23/U/beYp3AS2oo4oRVMuTincYY4cuhlv
Cp5wm6mIAA9XlGrp4dGs53NGBf740FUc5l4cZts3CiCmZ//QKKNecADba+ODnlMo
pvfgyxFUmHvUF4hVlbhvi8sz80W+W8XoiVba0bb7HyW6H470HhAytEu81H+kmryC
a9VE/QRYcEQy5gKAND7oqDe1UvLyPkAcKeKOzEmA/JOOmZhMsukA0x9aT1pljBvU
s9r+fFCnj6AHlFnVgsXAPEMgyDpdC7zpB0CwEfC8Q+Q2EKijVDrU54W3MQtwOTp9
0K9/ksDuoTkMXPDYh0pr8UksFmx1Cpc2a81jlqeXFZTZzBjvu8zdaGUoLQ3awHBx
dKEYAg+J9wEtKCldb2mTCrbGzxBgQSupB92WXnATJIN+ScnfxY+ud33xMxHCcV/9
MM781A2fOxTlaQVQrh4yD1ZEYUro36SxdLU0EKnEWgKSSHmRxDqjYsLV1/DIkguO
ZjnhWCWGKC3cLsCBFNdilKZHy9w28eyR2w50GH1AgZ+IiN6cIituQl5Kfv1tl4cE
8//kdHyxfbPPfBQrssL521gYW1bCXyuUEkLQeDOfrnqt+vLq1FXZh5WM1XZAcAtb
Zq2yVesilnJvlqW0ZTb+XtC0TDuLM9gQtovN95SA4zA7TOCL3/CVpxJhGP+lH6S6
c0vZ9G5TVP2Vga6Lz6zqd3DzVLsr+GWznWFXhZanK0OdURcLiwxzfKrMY6zSDNaM
DLoKA0i3dp6d1Tp22xEL8iC5GuWz8FzyZJeqMLZybSsvxR5uyvhWdAubTKjRVYsb
tWO1qiqCt+qVMT7NyyWwl+HH1XPrNXJCDd8nyPfmTycXQVtWLJcxVddI0mKD8PHq
BCSvEBHUspEIbO+tpE6NCYJqZd4li6YWbfF9QLHx3fvNNTgaS3i0Uz4pyH7JcqGE
uBnZRlCYGmS1EokBIiAoIAGzvVgGqSz608fsWqmnmftOJ7N0TEPljn0j7lggkx7W
/XH04vjxVnihRENKO7yZRMGnllYX9Rwvj7VKLVV45X8q9IEy08ua5iv+sRR5s1G9
yLw6vBS87uI8Kn43VfSfU4M2SGdIYMwx2KH0PQqSvV/Z5xJDF2ZoaLq1uNKQrOSE
PWvo+gox3BFqhEEjj1qm5vvS5U55UaOYZ+OIUMmFT1FY2B7pjDHoAPXutgnq6aOi
vLvilpxTpLJ/oDJNnepKBwTcQIzcfr/8w3EtSpqhGs0Z6+ApbdP45KgVgXOBV2Kw
42Tq55DAw6GKUvS5GLv6SJH9wWcUvzxLAh1TAqeAysuToVxXzE1Ok0rJgMQcy/jg
RcpTtqBXu1txthJsmzeXwTO+yA6OZYT1FkN+oy4LKydDitdhVPaLYQmbBOlp1yUQ
dEaV0YIsIVSOvO7MI6EPU+/yUXcCRTGxWYhehY0jfpwX82BqpcTBMNtkzInjuZm1
1dQY3I6FAmjO+cj/Vcw3JCb/RFCW63/NmW6N/2HUIXtbUkYBP+6uScaVrdPDG7yk
0uXzdnHmL9x+3LuPVqKH1BUJllQj37y9WRbFojWiGNkjqIF8HYhXsCCowBVnG/yu
yns4n8RBy8uTRAi3YL0Zwld0B081cF3vInLdLP7no9nLbYorNEugcVnmhfJYYjNa
WYf5q/lD8DvUOhqTe2Ez/0XBEbbn0i8+0Iz4RbN5uQj7Bezx5DV/0E//++hl+GsA
MjMv2R381VSCDTxC0G8a9G1JybExQDIhRCYKly2a1/VwR4oBFVZfIGCSMooYppNF
VY/gR7GjaFs4obfWdbnvQx6FUWzVAzCnaGzqr5VB+0pub7fSnaCFxVZbdl2IBos4
zKMUKwp0h68EwakjbXg6RFmxln4Ai+jyuxBgvtsifciJTQDKzV2WKbu4NGjLhVm6
ZidDWztnbxd+K5aTSeeq4sfs8VX8GFvY9IWTQ2ikQe6Mep1I5lij+AKI8y9xbxkD
4aRpmmM8PYtrqFh7Zq/LGVVs7DBhOkvPM4TFePO58WAXPo8yk6W/cup9+GNXoLSZ
6N9+7kk6lAGNJ6l5ucSuUhY/zz921wOb2cnkHNdPWGnc6W5EodfG0IymE/L3b6QK
1i30NE0vlqlRYM0gadQ6YgpRFPe+RC/fM3RRUlRT0pagm5ayMCg5r19wAvGgbyse
jpZxLplvTDCrm3FGIm9hY6Pb3vF1HaZWJocpCJ4JhAFqkIMISrw6BpUNLBWlMOv1
nZUUBAY8plI4lmr79s9fFeG8aK5SGN3Wl5iDyUnVr0GSbTENm3VPUejm+aAdCmRf
2wTeXEML/X+6LWVCMvDYMgY2gcdoB8fTfr+z9J5Kv2Z9LQFlXPM+7dcNm+ZH+RKu
U6OGgbL4A9vmn7X93LTPJwSKwKFP55S/w2IeeOAddKkGj/iQIB6fc6Yb8Nv0sfnI
3jLDyMiy4UquKUEWjGNydBeRPsWWwBuRlcHM8mAYxwsx4mw5edPOnVjXeIRpaMJ4
MrBU6eBQ+bzo45eqNm3FSneSVXgOhAuCzHVE66KUov64eMriyV35G+/MjOHl8tKi
JuZqUNXwje6kuK2oq1KL4rhZySQYZHfF87U8Nmz/xBKtXA5F2d6vjMlgF6Vhuls7
GNPjV3jrBJNbqDFChce+8FYN4rZ/BVRXLNyOtsYPyu9Cg63xGMfzZ6beV5OFP0zy
WDvqNKHxNJt27vWGfs3w4G3ev+1YDTXA768aNf1aQbi9WDe9goSo48+Ok5noRkA7
eUmEAouCQ7Iz9Zf+hMJ1BQ+58OtVTFIldr+kdkDdAPCGYiHVTheKpn1rlA7ATtck
sgdn11LeKvKo1BbvXCoTXvAsT7d1gIHMdJapobGo9RFQgJrzKRU/VCDS/+JqOLED
vkNmliGAhtONjNnx/nX3oT+VWczMGxDtUQAvohnF+ebC/j+/LzNS0dcrJgytSE5B
+69CdFkPMYBk/0CTv+r+pblzYcN3UKtl/IG1NZ7aEPCXRoSvxoJEKziVOZX7+iWj
qccJlXqPnRyvNW1BeROwtihRt/CQ2AEMQtAyfXCmxBXHq5mgJuKahoB4eKhawG3Y
/SYnTHfnh7AUFkQOJdj+mHlXPsmH5MyW3jCUq/lwcvf7/9yJOwf1PZgHIFmZYUMI
+wOJ2bkzS1R3n9kzQsZtceHao79bV2SfMn1gERLuSX3DOOGEdd14v6fWtiYCoiAF
iCyFsQ/g75JItF2fiUljqWTJEYLT8mtQWlZspjzY88jMsiczQI9NTwKwzcJTLBSL
yJX2MkEZlbmi64eONedkLsIRlvK8012wGYXf8TBhdjcNnrhEDSF59UjB+cSJrLZc
ZPQBAp/tOn27g0PUUDgz6WsVfx5Bm1CrQRutNJFj2T98UBaGQvYrjT0ZddVx1iOh
EBVBv6CujXix+JDZ04mYQHWEsI6G+1U/Da2QTUMH5OPSSfpUPIUYTtifB1V75CFu
dK6hu/YW+u24m7xBP7KFigo+OeM7WHxzdhCLL1IviJ6HQi+Ht7Lxf283bj7OjmD7
NwOo0DVkhveNCyaP8uJy/5zppu4voRiicw4r51U8gWiKYPNbgDQQmpf/sgNaJhn/
pHSH0u/5ZqSphN531yUsB3DJ9AFEqrSVJyww14ev6+JMKNjkA4Re4jH5MTaN/GEQ
dDEZswB71hGCF9Xd2+DR4g==
`pragma protect end_protected
