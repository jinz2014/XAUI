// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jM18zpyywDsRCGX/XeSzYjRrirFnmSCIigCc+aXBeD+lpzYnzt75OWuv4TN3uWoq
pogRt2zmdMbqtLrNM6bvStYMP1wh19HG7rDGv/zS0Zg2pBC3hePqrb/vuWNULTzj
s89cyp9UUhrvoRiqE03uCBc7OttjTE3ecIjTQKz7l6I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31152)
Z4L78JuwUOTlUb5InQUFSxzzai7h40OQN2YjQiAf0Q27iJTVHO3vQ8K/J8qQcNi7
FPveIparBVnpz/nwR6lbvjS7EljtFDscSzQO8LVN4ESAA8ZOqsfpP89hAx/fa3AN
o7z2/xvaQ7xiLfcQ0zobhM0pVSP5GWmulYjN1oNcxOMc0oOvIPeN1fVgr5SvKt3q
Bv/xUsdf6f4cYrGqbRVeLDjy1XaTFSnKHBW+ZS1Q9CeldTHgGyISl3+HpAcB73PR
Ap3dDuVjR3XXJ5jengEM873HpGSLjI23D4TqYlSjpzFF52WOGEox/0imTsjlYa1D
Gt4i2Xa1e2dIkmvYha/Mhxkj2XlqAPmIYcQvV1X2Je4a0Y4zRh8YYVTb+MCo1g/h
yahssCQEQnlC4F+jCtuLDDcCpNt3nlqRCnx5GamkiXZiX4yEvRug0dELL2ekQwCa
/OHcE084t/MoStNGxsXhnHEeCuwHg7FB8F7TBKg5Yy/NqbE3teOiB2b1edL7GKix
2xOBaPot+ME3AmVYmoIMvyES2/dm9hmcCqKhgsQ6ZxBl3FhngU4jwDuzAJOVg6mm
sxfdzFQdLGN4PXF5s0ka2cYm2epvNGQC9moMLKzDf1zsq83q72+NKjcvGu7HGba4
ytZNi3qAaivHVewgZUCW/1LpjuEWu6SSP9c7EJEp0UIYQvaAPAI3u7wJgUkAwyai
pIxYikMieL3+8dE1chA/vamgADK+uZRFy111M04xsXSk8uKsOtAAEcHTBxmKYWoF
rTEe/8guefIlJw89jgaT5JdEGiTPRwoJe8NMfDXBVRrsD8oYuC9rG3JOsiwIMwea
3OlBgMIVnbcshCPw3EJ7TIdO+lgs4r+2IGdM6ze9StR2K5EMZ9G6h5g9v8B5AC9G
lfpn83a8BwcMVWsbV7nqQSiPr36gHuxfR2QAt8YsAI4nPR6D+L645Bxq96CCYfit
dOSp7DsNMdVY0J1ShBPuF6nUyRd1ZRBX6KD5+lxyLLOFtogCLM4TINnCQakQ6Xq3
SqiwijSm8CLnywspdzmuJ+zEiOctFjq0nNVqaoP3Qi2pfgUN0tevgrlHfyVB3Qhg
+84A8NK6cp1mXGd0+t6kx69q+EcnUwG/T2eAXHOhImJ9m+thwFJdItWp7yc6uvZt
kmUpL9K9mCB3XyJU1oyopCGpNe4O3yanftL++QvCxGro6Sw8WPoBYHKqPKptok63
N9ggg7z31OEHsTQWsdkk8l1MnM7rYThaPIe9bfrTkDX9TV2jNQ57RwlaciiHKatx
E3eP1aUoeDRa7t/g8DFa4yfMnIObnDNdbLFiZq/PF0KIHQDxNgNfgpO/52589fwC
JH8NbjLS1FngcCOLBtbiRDBPFNHNzBZsybCGUp8GvOBLXlLkbHfMRszD2ztbprhE
XdsXwm/ka/GFVhemjXl1efHdE3vfVtzQ+z21fflaMtiYrnUwThc63EO48W9KIuy+
DbF6wuTuLZS+d7Jsei9ymfxj5C9DiYHa23iosnHIG2C/Bn5z8XKyQVh0AmKCgarq
vRpCTJc8Pvk8NrbGOWQ/TJRCF7kiaWbUjZxdvoXMIOPATekDvzQcEzQBDw62SkYx
HZLrqQ7yTDrYkyCKbM6xPs6LUZK92mN5OkfX8uAF2D5rITaVmhV9nDxX+3aLhv35
ldkOqs/6kMq0juk0mR+DKdMwL0znEzyJ9XVf4JkjGY9VZgJlrpjgPIJASots82d5
pCMp3iSYOVEuyKu3YRCLdro/pM1qkMFxukyPK26n4uhfhCKOfJpeIs84fOsDc+On
8VEOF+5Va6fFGa5jPclXMSW9PEUocdoiVzVg8ljlK5ElyzvuRQYuPhDHndG4czsD
OTLM5qnHBrtCUYcUvdece1gpZXXBuQSpBO/ay2YOqTib7C5vtZb/nM44ahdHcwhI
0KfUIRzKsjxYcaWo2lInKshAeCKiwiTNxLaLeyGt8Q8stNjxhysXLCnca0eAZA/Z
Rhg2W6MAFExXzwPzrrqmDB9gSI2UOepB+wfIUKDlEwLlATC4wF9Bpri6eCg7VQVI
2AHWV1SuhrgLCTS6p5UU0hEOfaHRXEkRnv1e9Q4nzLV132jmIQNxHzB82N6ay66a
9l8pJitsqSwiOfDtOlg80hj3d1bQiftvnH30+9R1NjpajLj1vtCrHb32qvjksO3L
EC5V3EhRegY3J+JvClEGHiieDQU6qY9OSwYLktxmZYPDeSHkuPPz6LH1+jD8BlAx
1RUm0IdUsh7+2LIcgHcW5AVQURJX66osaiHDBu2lU0NdIWOGXgMtidYffBCWnICh
Qtfq+jJlDM2yavcBBfV6xgmF5mAzGDlPNPQpmAQ79GFIqPU+fqBeoV6qkHVeOeez
evtHzjMigc28alKTXLaKu0AHQm/RF0jJXOaVJZmjZkriV+AvmmggmxPEnyA1zLXl
AcYQ5I/2gZBvwOSz7pBRsA7HsR05KKCAzYR4ObFcUG50OIat+jDZpScaixSYT8r4
0KL6l09ck4VjQ5Q0zUTUS096zmVnsejAnRi/lxnwFbl2JD7jPaSffE7ZiZLnxC7a
VdbY1CqB/lvw6sf9lop/KRmU+9FGo899tTI1GgSsRwPB5bpbQX1I+eAVCARUMBHL
6+DqX+P9+QMFbTrj4ujUMW/iofYvbR3BRtw9jlrKlmrfFsKUHmTOywP7MLCUxo2t
ToRsyFnQtblm/7Obw2AtlSE4gZQseGawkc80pdjIbklraUJUWLwmUbD3vPu3r3jW
n9g2PTqIyOz9D+DVYa2o6jqXp2x1qwakESxxB1JvVZ+VOPhroB6BPqqoXaiX4HoJ
PuOmjkrv04qUM0zj9DCtqS6v5tKfQ2RfB1jt3zMnaPA1pCbPEAN5H1Ed+N5swUFx
5G/g2N3QfrU9g2c9wO7kUw259+NTOM2g4cBRS8fX9KUx52ixTb8zJCM6a4Bo3JhG
yeHDHL3FF8rYArAfyzWzGlyzOeEpBKKxwgtM3tXx7DmgREoQhwQFZEKzRw/xUW9a
lruReFyIOD0igoHoA9no6J7YElUzgNee1SHktrQpL9PFucOuvXtWzKtLadhIpOZF
CqSl+hxgcfDgnbTBrH8qYPtzN7zU9eHoLgJThjnhgnqB9X9xCcop7BnlPkTBz/S3
mDHjAMhpp1xn6va1f5eR1v4Zcb7PsXLf29zlrPXnZbPMfq55CobtwwEip9uov09N
OcicwDEXD9MIs3YYboTYbVnbnZieYmXZ+97b5Ghrr3tBGbRzd1klXAm+VEqOfsFz
dJPspMOOv+7TwEgjrYgSCrAQZVec56kdCMIYqjyJzTYzfNq49XsxOBdXuUn3wniG
Yis+gFx86afO3VV9PfVRtKmfMx2B0IqOZlzYu699g+4AHhVk+t/Y7hjfqbYzDJAl
jf3HA+A4BNOIrXdtAGk3kpkB0uMO17/+9EOdEJhgwguaDmnjOfiKRoYzTaXVmazq
06FrWq3lD5V+FGpH23guaR0Pe0mB8v5ByZbNnSBO+srNMCJZ43vUgJk//Vj5e7mL
iR/6tRB7tlGI5dJOdNZLhHeSoTvGn76cKYDWvq4qRwMoInjSzOCmtUvqBT4khFWC
+P3B87lidCDDNO1ZsbuCpsENyjTgPEaSEXSzA1DEcv7lhJvoQdwzXdEOs2DZScC6
BdF7kO75DH3MAjpgWCqTVeGcTXttjFxlqGGbNvRWSNfXIj9YSNmIC7H2MYvcEgYR
nby5v+XzHSvivLDiM26JKeeeDZtXtrftHqv0i3Lpfs8MM/8kSYBE4TUuB1Oh6Ii6
7+35MEyZvbfN20YNVje3ECLqcxNTTAGENwqyLjdXlgjWKcNXssJeUBHvQoBlBVEt
mJ31/FWyCbgXce9Nns+540OZYX4gKifPxHgqM6/L6Nb0vFsmIDUp+ndG1NDIO7y8
KkeKYVcubHUiizgrafzcM1W3j581Vrfh9nHvgQPcGn1euzkp14Cvzr3aBjXQxHTf
buD7qquWyGfIl+tiaJnz+VyuXhTPDo81Qe5SNTxVHYhgdbnYyXW8hy7JskU/VZ+3
VYEiLAH5nFz02WWGpCMlw/TN2PySSqy5bNPUPF9PGeSj0xhpyp7i6lu/Dgh63R3o
HP1owNF03lcK/oUFoB3tn3uAtyhjJNKQJy+p+/TFTjp0jtqijKmdwHnfYhu0DOD0
8nCKhlJeCLqvgBdeKWTwq/EBhSg3ONfo4KKdygkeDYjnWaeO5RiFg9ZqTwqhx3Gi
lUas7wcWvNc3z6ChTTGerLGnbJJLNygmG3neThN7UZd9Qb6tJh+d9A3neln8JT3L
Z5hBw/tgcVlwEr5M8yxsvYdJ3nYrqoF216OcJNdi0tffpNWhNf3QscxiUkGC4mta
p73m5erAA5OZAgXtdi9i15vqa9wxeC8VELZnowrv2p6PxY4OqHJCfbaqRiaMvw1d
WfSbrL8w7etgICblm3LNRivGRmtYKWhNVPfRPthVjKd5UAATV2jKbg5qjqHgI3Ul
BwTJ0hav6Fj5HOZGh9g3O+QmVGbsReHjk/V5uR/spWJxM7znxVnVGyiw9OeKE8Vc
FZsxDn2x1f7F45pAHoKuhUxv7YP5tKKRmArFjxgSI9ZZwu75/kiqUMcwwk3Gbbys
eJnKDPs27oluqrpab/G/JwkFyKaCN8MD/z4er0ZLfKQ29/Sg0YVe836G3Fh6P1iV
ChN+uuPXdktK5IeoiPs0w0D4+iSYnpX2/uhWPAO4VMpDnPOusdXOBwUGohCMpMKK
XF7sbFmVxOCW8HYIbv64qti9ZouHIVvbDS7us0lXJcFbVvKOzjrzDZRiysP7Tf52
1e1eIAAuJEWgIoqdI2cy8Z+RCA9f/iyOCWGIlP9f+XdJBJ3xSKcK5ctuzKlFhZTL
DK82MNMuS+Ujimmiwn4Tz9lXpujU0OM2jd2Rfpdzxn0A2+Z6/+rxRfnWkYTy5EHU
MXN/eebCJ3WeI1ELJIDLontBaH3cBw1CU4P0qCFvb8zRjBsKcMfl3NYdswXN+W0A
e+oCWhmhDnZddInPV+jHsQPLVDXhX8nCZ4flzz/WuyeUutefOseM2fIZcDR1EPCi
AzNypP79HWCd/6eZaMpEUxqfxPnzhYsiMXuTlgHz9ku8ldDF7MuTtNWz3ZyEUFQJ
YT+34S5VTLbhURyhAjixJ7mrTyVaIRy8tE6Tsnr+RcqW+/iCJ1298oYt16tB9pvV
mwam21v4GJPVzM7cLE3TbQOuXqA50FwWb4yLKXnumG3F14iJ5NLEhFYvscGJzn6l
b67GTADqJt9FWOgfsa9T1TpyzJHvO0Yedz/OZ+Ug4Mc/5Au3SUb/i4LklRkkeTaV
BIJavW+um9HMxHi59EmDVvaTjyFmrJkcs/fRytDweEVllIcZYse2/kt6CCf0LVUe
voWoXcriGJph/o6OrBbhRV8p2XSeW6OkcLaxkL6Tme7HJRlegV0oxQwDLaeMAtWp
x8w1sydeC/C1cmiFb54rXTSviANL9n2wfrxHowSaHr/sJxcjWnYqxl1NAKe+peu/
LHwZorF6j9L1hy4/Bu7eMIbzRuPVSW5a55EoMoaP3R9zfx1bV412rvAjYKdT4MK8
o13eDX8JiLhcjwKn7bTRhasGPOb1etCHenl2Xgqy4bb9/qLuknVqI2OiBV4M++0n
DVhQDh64o3Fo75jc4GMV+oCnCuUu/e61uoRdNXdVS0M7p2t2+ZZb5y2Q3K75ABnh
Tz+gxOcIRZ1Lbyx8DoBwVvAJLNVz+XFb+8x1rT6ngYf4iaIL/aKH2cvovWRY/0Ed
pLAUN7bYZoLGsyu7ysj6t+uL9QCEbTwTqI3RTsuowZlLsd5BAOZvXQOiHxT3AETz
ZNdEm9TT+hRHhO3R04S98Ya5/WbHSZFJAOJYxEjrRLmhErTi+AoXg75HdhvReI1Q
ux5ddnTbmNQC2r5JZ4IwfzBcuoQIn/DnYhuqW0vblKv/ZO50FZaelJKqQugFOnXA
jL1cicm0oGviewTaHz2mc3RSzxQPKBkYUhmUzKgGS+Vs+/OJTM5Gg5EKzWbZsJzk
beqQNP3sePaGw+CcdX0cb2p6oW8KmqUtyM021JT6EWKe+K2ThMGR2kJSPCECMZgl
qfbou+/wpR3ZSR+Ehp9RKtOc5hf5QFx1TpLW38CD5MgMYgJZ9TLfYjEHn6hOcUsV
nD0Hqi1m9rB0Sf+4tmCq7BiIkXLRcZ8LtHkozn/sSCsvSGFF07L+vJRU9/D0zmOD
79LNvQAMhESFyMK7ndSiva5Gwl13ASrv5PhHuGrpi/L4dcmpGvxs34F9OdavKg+d
jHbA831qb2la8ATqeiCJjc+ar7g2ioiod5r998P8mznUl53xZZqPN3xJP9lWKDQJ
H5AKn9Pyt3Cq8OGUpV8J28Nf41TtlNu1vzrdTg6fHyOuI94y6grhbKX52CjoAZGu
4WxezUosNGsroyNY6ESFU8rKUkqZzvDSEgTwWofnxsR9jxkvOd4TlvDdcCVeqkEz
QnNoayZ9ZrMdnHsGoR5GDAxI67br4rJKWL2G4D0M/x3N6WkSMIdSvldkQSN2RBii
hR9aOK/Otqcg6Rsnzt2NnYjNNhlxtKHuB2/gnsgh+5Ca6Jb2RRYLj+UfAQ4A5FtC
cWQ13HlzAlg9JSlPAo+/Ne+7kXWLegrUU8bwcOH6bn+B1Th3dG1oydgu/35jHxBL
aWvkxScQD/CPZ88Gr9Zq+Ikr68QfbZay8NtUCT1Wq8auMwLqhFgixQRo4N9McblF
1a56n8eou9xTiZYBhpSFKb2koYX56/E+KJDZC6YUGxu8LjmumeMbOtAdRzS4vw8T
ZaO29COqylNkD1UxZCVdQrndT+5gTMF+614l3ols9Hze7k1BnrJaW/f/cUNQSDL0
+kFOhtpJuxwBaLPggRCGhrKnzssW/DxQlwMTKumCScnvk3S27NAm78vyjo24zgRu
t8uP9zwOig6+vTKS46Irt3Ggwkm9PILaTE7olpw+QpD3V0q12x+6EOmp2LHzztI0
cNnbHPJWZMUdOp3ELMGolHS9yskAhU5EEMgGBoH3izKuT2KJ769pjMdyDlc+mv5S
RXkqwK7yd/w0smFVmRPJemuhwJ8QC/t9A/843DcziY12Zb20nmOuBnKs3bZpebKr
aGNFKgfdbjBBzjwty0F8QL/NNA7KlUqLaIAL/letro90dMnu9c69rdkIUbwPtbSO
Eqbeq0ay33xbHaEj7OK1E3kXw1NaZ1YzdqA+/iikzMO6DQcQ3v6oamFE6YCyBU0+
WGIt/Hi/yCsf2NHQdJFzeNVR8vhV4v8wWmJxqaDdZsys22ZUK30nE0fKWYIoc6SD
rnGPgx8qdLNOVqK90B3wtDT3sr+Vq/ZqD7Upjj0QIV6BjCi/IiCAGZDIz1EGHUbl
eG31V+w9BSnDRyCjBG7xfG/sABM2fw/sP3k57bYW6SX+TymuiYyAgG3PJ9JvscE5
gTfUC0bzyUc9y4I4jk3uQlOCkuiVvbbpvO3G1t5AQpRd/+yAy5WrmGNAn5VbHO/3
vId0MD2PHPOZMvgAVTJK78z54qStxtOUAtu/Gy98zhRNSUIlYYA8hEHH42kaAHuK
MLjbnZYo+NGKQ/vuWWbQKpeqoCqzhuvQbegPdJWPtyTWQrYoW5/1bViV3gVjfFfk
88JWszt3AYEHFUerSl0ngzWZyT+JoccVl2FzOThtscXTql3AYDrIr6iU7fh/9pTr
YyXf4Uhuw0CjFgGT8/3dc7sNphbIhJI8CLNfTOdz3i6asF4r25yNs9Sag+UDew2i
KlfbJK+XW2SfDI8BdYU1neVj7eWP15L6j28C+Tz4jRoY/XiRQmCM4bMkvjglR7ob
SetNowswyOmG2u3WRmrlvuOWqrmo+nUdiCHW5n//DN+EN/20VpZesqp0GhZAKOSY
ivmDwWxUY1nnmhhSTkZmr81cksKjheizFgSHHVjWKPpHJzHM+Jr6rKi2RdOcQI2D
ZTl/nn0YyO3OzmI8+mrAESRCRPFVeu512Wvwf4q7yOZqOrAigVMXjtKHaG7GeHw8
whwaWhK2gRfYmX3/kY2yXJQ+nS3FBM9fhUuJ4SgYkBAvmpnbopVi/PXn6BWBaZTY
Qd/kji+PXu+F1UO23M7DPvbFitrs5GPconAqeCukdqSUcHWyV3EvA/T/COWvFrc7
Z2kXhS0/P2xiaPKyOXwaOWvGm2CVayxEImyYiLqHEy0We4RTfdN+ppPUPn5sWLLY
A6IYhzaka78+sTVvHJSpx3PAJReGQRzXKuTf1HMWYtiq56oQrjY9Ok17kuNZQUf+
I3qRsyPRvmkJjSP828x5XLU9eKh4FFhLuCLh1XcoZ+lM9P3Ojt8ktGaKTKtDi5nR
yvad6ID6kdJNdbf3CKG/CD54q0C5RqNUS3brZtmI6opGQuj2xCDEXQ9A7dFprg76
uA3HVDy4oWqRK/ZMx1sApnSqtcaIKdhsi/Jf9mdNP0iCYIARjsC6eDlZbpJWhd1d
VvacC1HxOeXG4XQ0oGlJruiND7bWHehqhhlED3NIbBNuZVDZUFVFwZBBI9nrrkco
xO9q6AyVBPhMCehBBi5QY4AlKwHKqFvT/vEt3ZOfnqLGOeVCcBE4elMlS4ZILZ0v
x25xeNz3GZAG3U4vnr9mlyvLkfd57dttePWM2xKKdnUuKXM76KfcQidzAKsfrAWW
LtY1NokV5fbkkcBvDq8sS/Bt1lRwIK8X+AM4dWJubZE2X86xDM0UuRX6p4EKdt70
0gM7snCNGxJJldXQH2eu/Wkw3FBBM4ouNJpmkvBkwglIGRj8B/JPcAM8fCqDphIM
qfxlrZ56V70H8DDUtIYUDK5wNDqRMNCvgiINQCrXZoUzU4Sv7FGbS4GKpNOwDcC3
bWuXugVvdwZZSCI6Ru7+XiNlzUsP2gQwr3bcv4djQnPV68fzkcDagxwz/ABeDh6h
KSN0/xJWzms75nlPpwKWfK5hW1BPOIQdLjh+quit0wc+eLTx5a8nD/3D+zGAb14k
e7OyU7kysbFAic5aUNETw0BDZ3+hzQSp73NpnlkXav99qmpULEBvRrxJv+w5TK2t
ybJU9LWgprWIJEiJghPmWKbYfg886DdsKtrTCisUmjU0KuHFzoQRPrA/ScWhKYRM
R25kjzaHLv1HPWROCE8g5yQA53Q7P0lXOOra3ywDxDc7w7IOSPr4zej5qS30YXM0
+RwDSNZchKPAYeAofkqq49UsXJHOcDqmMiF6ZSDWLCIfLr5W0jscXazHLOaxLnAd
mVdy7baHj8WZ1oj1zI80/mVSNbwOBoP7U25OITd4cyecpKaGslpZakGh2YY6XJnV
6GC2070QrYgp+7gCXfGqG9YdUt0MRmSoVdQF9joHa542j4g7UfFvIDGZKpgJ8QSW
njqxKSbmI+NbkZeBJj6MdW9qEJ09Ugu/ZsIBxg7PYBe3VGjz1mYxBu+aL75LDWOW
szqdcC+Rrfqtfc7B70/iKDThNXAQHTwNb3b4YlLxgxtWB/WEUmCvS5akYUBtoFPA
LBtTW937WTQaCT24GXkyCxQBxFtXua1a2bDmIFNJVuyvtRNi+YALI2FcQU936pW1
Lz9a/Dk00ZIs6a2eWah+PQmHpOgNGGagv39kIGKe0SCXus/fLMFvm/IFPpkuayJr
Q7YwvDtocBFo8qyiaD1ORyBndcgPgZ9gMasHMVdHidH+h7klXTxT9AAJrAApP/8l
gcyDGCAESOus6p9qiv5lNrwPgMfe2md/QidtFE0i6942rx3Y94PRu/D9LWUZKlF1
bABQ0oGJOsnzDlpqcdRZZwschyeNlO2A/993aOTzVScnaS6R+PPNDWviKUcAXbhf
rtzvON1c8MRzQ1dXtcowm2JuxUxX7zwAiVZ1Qv9lsJ9vXNZ05k4Ec39lxXgqFl5R
4fIpA+uKCJqJHt387wB2qcct5BPbxzKpyXvxH8G1KxqvJ508fQTkZEQq5KbjYgkp
RUHjOZo9AQvQf1eX1AAudzZfwTiXMprEH9k5V6T9F1nKF7+gjRA087pO6A/2ewyl
C5vpdDKfKExAP14w15S8aR1ucJ+pZnZwnkt27HwSMcAROB2Qgk3CJdRt/E3CZ1b6
7VXtAzx/f3Rig1IDkLaEm9nzY6CRe1aKFNBapoTN926r3U2aMrwij346F+sF1eSR
CHZhIl8n3Hvdk+GsWHx7v14PQgETewlENFiXTmtQnx/sJ+21PyG5oiHzj28p11XL
iKW02e1GsK0OxiE56qRvthSzw0Zh9MY25Uhx5hpUbuqDGWAcIIP0c4sbcSQt0CNa
q3BmwAtZXyjCrfRmSS4jQtSUgo5lnmP4abJ3Vssh2KBH2OjgWk/ffj5dDeB01x2n
4v5ycozzkRoVudWqFIdU+lIs/ay6AYcEgy0i7AMCi5gV1Wi21ONgK7AAQQ27jquB
oEq71rPgwzSmtUD/Wl5rTlfP2ifT7WYk1T9vAk33YJ1QZaeghJpeAC6RUBCU7vuE
4azX4OVJxtBaG1paZ3nXZzZTMyA7LctnUKFB2h2Bbu/YGraHfuIK0H6JRU7rL8s4
MjiZ6alkRzlxSI3EyltBxerJVyUSvV8BUJK/787TrNzxFuKoobijinufFXMLkWdI
+stfBvbMl+vyo+7QwuEe/opOoAscR0tLB83kd1m1sdiqynnBtme9WRYLGUw33v78
6WS5KlX/8VUnup+2phheDtpm7DpC+jggPDTsRvb8wHlTam+QvHmLJ8dC7eM+U364
Lvv1Xwrx1jLfv79tprEiS6PE8Qxzx7EP4WVdNXU/e4m80AQ0HndcIC750GNIywfu
F3Tm1QlFbHxM3eiwXS+5HoNij2Ni1+jaazZOzuJeXxV5ff2azrTOFCYih0xFoo6J
KqWnCsk5ls6joPEOAee06aJhkTdGj2i83VsUBeEQ4Pfxf5OnpoYFbLDq0kHxs5jA
NRgpRedk81e6sdG8WcOlXLNJht05VG+jOWr6FqHWKepQeGOM0PodP/tIV9wCkg8k
QTyp0RW+OG60Yhf2DW7JgOnHajpfAcs9osM0KovJ6DlRRIRMRuaPoQmqm4T2faFw
LRT9h0yEhaeQYINEvIfAQjMVNUvfbfwkqkl1CxUc6IW/TgksLBKVzlo1MxhdhfwW
Rng7HGbmXdNcJ1kx76GmOCn4MVHVH1UnvwCmlq+rhiY5mbmIITX7QPud5CwJ2sxL
pmBDXYR4BfzlfHmUVrusKQe/c2waNrqXt7Rda2+uB+IEPOqnhMKNvYxn+ab/azdN
i4en27VeP9lSKlz2QrZPgW+fsSFZHNP4EgokQEnwwt/e4HpGLoH3ruh9b1X3zI0D
AGSt+YVuzVBllgq+S5FhiX6neM7MwJIxtV1K72HwYJ8Ig+q9lTzindmIsfI9bBd0
BFKVWb8tVwbX03S+wFk6Ovr6ij+zVBpjggRrFGnOXJlDkiHxp1xZA2SG+B+A/AXo
aGJ5JINa+5PSP+XIdaQXjNkF0m1YAV2OfHUDzmyzHqnon6gyY4ow96gI4WBOM4L5
GE9THzhAxWQACl0Olw2IR5FVdWQ4km1JVHrB4BqBaKmwQisX2nnyXaPD+/grwODI
/UMzcgsrzCM3HUSOVmCF4wG3UmvXP2GIif+aPxrWyyT3zZ8jHiCc6aPnaTU/X29+
L8dNrFFPkskGpEuL5oMw8uwJG+S1dTuUP2SyxjD1a5hH1HrV6lR6ROemKpWyS/vG
eYBQpVVZVnA1+kLNNYA9vXAHa/D7mdZ18fvfzM5SzMWpGNxfO6zZL2xBjXVO09g1
CZtFgzb1n2AVKuDBvhc2TSeDatn/ASHTft/KdVw31VDabgx6RoxuUHq/iY6dblw3
JX0sA9Bo6NiFZFWYOU4Vk9hUW0OQwSuVinsijTA+x+g2ZJRIYuDYEekxu6nnn6J5
/CXI4+PaGVAkg+SaASfNaO+1Q5VacTUGuvgfyeZHFlMX1HKonBpfYmCPHnSjKg1S
fWya8C1XDrkVDt41KrvNZFwe5fvOTcDF/2KVVlVi/CUNtmmX192Solbc23h0vjRf
ZLvup8Hi3xx7XivlS2bTPjHsk+s7xDilfNn2hdzYWKQw7M0vCTig7SncuPWB+mT3
R6G6CEJwJBb7fgAsZhZSsEESmcmlkohcEul4UZ6U7KjBnMBEMBQWOnS6JQGIujo4
CdOalTNd85LNRKjxie4TRQF9lN+Ju2OZ+7DduJEYBLZOZQ+LAwx7eRSLAREoIpg6
D60IdqqIsEYzkzwraXZ9D8srqg+xjlKp/Vlq04BG98e+hMlPTiFa4WIawAjdWWTO
sTVNkD/A44uU/hEVebcWX1oFUfXRDKhPCHHj4Zb0hfa7bPxBHofOzVnLWnuLnqsZ
OTPFa2EYTHo9jhg3qpKwxH4evfVidZNzA94ZFnQoZIyw52WNXZeknl4qnuJruevm
aLOaMYCmGZyf9OQ1JadKRZuSQngzj6c63mGfpCU/2t7k6DLkobrOnyOzinad0O+Z
ZOMhlKIkRNwR0KGy2kjFgaOy9CsWw58H+qnkwTQwgpZzUo/yhOrCWPMpQQOe2qu3
W5oELSFuRYLF5N7S0kfJHWnLFXCbmLwp1msaLHqiiGsuYu8h5YYiVqtycwpwp7c3
LHzhEjBw1DLqB133uWeIx0oqQFDAu/feV26fiSgdGdDDht96KjKk1p7P1sQe1Vk7
7s/kxltIe9APQ35F0XgDOxREAehdx4fyO03+F+qhFxfK59dCfahL7LoJ8PrDNosy
iVcW04iydrWH/neqDR/XDdYyNoupnSXWp4wyNSgI492+UlabPsXTNMxT7HPIDZA0
ekvmT7w7rX/iLxJsHaXXZzmLV8FRlsM57YrOX7+6rmxd6EY7GnAAQT/JgX14jo9V
mclEdbqdmLGKH/OmVU64esavAUdSsW/RW9Mt77yAwh9x4GN79SxFyoKAgoaB7xHz
GTxnp7cH4Q4pTbIOBARg/MubxQNOfyMviLGg/HF2UnuETX4kY/RXeR8EWQva8noE
BbhCGUr/s+rUJ/Ph/fx/kF9w/uA6rVaRIxzJoJhit1pF3TOQ+86rnS6dJZHL3UOO
i5Qid0+ThfFFkeEInXw4UiT6LYjhGiHrjIpYZPA1rB2vGUhpgjbQyatAFGIzfEJ0
yr38AdQcl01Qfx5wBwS6XhWfla3y5Gt9rGlzd9nVDeS7LdMKSSLTpWmj20e9p1R9
1/qU5sL11npVX1GTaC5vEqmcTs+hcMH7St9mQH64FFe1Aa6jsfiRerUsyT8MoseA
fOf6BlS84miuI7a4faqb1Wj6mHgz0ROn+9Tcl22Yq4wZtC+nAk6k6EfqtECYW8Ur
gpAaz2i6vVr5R0uvPD+IwuSgdesaYO9qWAq7hteYK5ezi61uR1MUkfdnHM0na8bm
n1acFWGvmPViJ0S6YFHlnA8oM8wPrOSpL39D+TpnCILv6cXZJ3W+NhKB9WEwed93
xQB3fUL7VKKehSaRaO+4jIjfFL6wMb8NqJGXBomec0JQYUUwEHI7VS4dC59MjuRn
wVSDdAuCHkEOP/WaFvCGGrbB2ZBQa9xQSioC+iyy6KT09pmBOyupXt3Ax+Aaqc53
dg/qANf0azob1UAwRUZ0DItgsXbADUGntQjPsDck7KkJ5IaUXZKnSgVc3Q9KCez2
7txXwWhCbpXt34VIS22Gijzvns5G3QaslmaveLWNIkg90oQ4mSA8vzW8un76PSQp
mgtG+K25YVM3W8I7ckadE19EEEL/rhP9J6TVRadAPlOJKDrVh3YsbpTchcSfH9He
dv+3wO26T5EmStwAjtbhin1s/9SuUsm2GXrrkIOB4WF/deuH9Cag18l+Sv9GsRZ4
XRMa3iTxi4OzKHBI5VovZyK8TIxDBeQMa1QuwQJYDCG1ajj9giwF4VZBCbU+qWQO
Q7JBAHDVmEgG+nTtr/fC/tibBhpiEWXTdMj7W2uxbx+XiiRXvrbAo31Ol/3CycKf
fACcs262CB2H91Bpkfqcs1sLiko1m+WCDVszbGnhmu/IwgSLk/YOzctSyTG0JUjD
6i57kHdKBV64v02u6vrd4K6mMhzjX+gGloVxCVzs8lTdcsFDuKUKwhO2hq2k6HFj
WyFMIlg0XFJmMZFvDg5Ks7ir3RWMBjHTkaBjviHA3it377s8f0iU/7S2kswrsNTa
EDYZHV9SzV9tPGeU0W6SVaxx/VQO/YcOtAtRTX9gs5jfwnMlheM4M8HZH4IR0tD/
W51XyuwPVoCp4XFCw9rMw6FQtpFk7ukwXuJqNSIhH9NoZJFWNumVR0yVtMWMYJPR
usebx/fGzla+dc53zHvtb6sCMzxY5sKNL0CBvcK9kEWo66I4oNPzLIBMPFZP/tTT
89RyYoV+pKa0D3AY6bt3mToZiOq9sF07bDCVq0CSQlU0v2vS95VeFp1VLgStZ0d+
nctc4El7CwVnJSuanhtQPGCYCmrQZqc1d9vYONPCZgEAVVQZet7OSYBQGopprAFI
Cfl1Vv+cx0MsE3nUC6JevSXBNC1leT0Iex7B0X+TSeOffDtoVDBjGTJPfhs2mrmV
GIJbh5SwZ3gx4EqpO+gLqdB8kD12MIJW4hlwxev6C0k+Np5rEiqXdL54DsGmS2oZ
LfTHbA+JgzItRpS3iriig0TR+ExEeAOrpf/BU/f5KVfvztNX6jg9mqR2ga5KKS5C
sob1imwaKxU+Nx0d9i0Bccggm1adCbGpRBiruxoltqoo/7sWsWap+xYyRmskj7TU
lbJq/2sXrnkEujq6Lfsf3p8XAU9UUnoSG2TTNlKjSrHF5D0JOVgCGsVp0KL0X1Gc
9n6V2YZT/mtkonK7uF+q9/ePE1Djd6VCMyRDnpfOeXhz/pSXkUOPVf7X3s13/O61
InxNI4Gpbt2clf0QIrpo2WYwGeLPqY/X/w/FwBzh6hwsDGRv4AaDvF36PrsiF1zc
enCXGsOSXYqUD7nvCOtr8amIIxS8x9KC2sUVCjWtugi7xA56c5/D4xUzJ3sHtiTd
nO4xi+8W9pza2t4d/2hizdUOI3lXTt1kX6QiioBS/qRb1yoeL5tKjOHfKYbdlZXM
36SEZoarvQae8gY4a8aV8ZjjTRm9tplNsRLtB2jWYpk4t7Z1s1nuwW3l9Nyr2hHC
g12VhP6/DJKpmPAYHdDuj4ZoODKTSO6iRUJ8SNDpX1mu7+f1AUSvM8PLcxiUDseb
Lo6/fKxssQJvtr34LZZkgQa1XS42cnAj9L+UHSimfWDPDA52QTLNjnVnjC7I1R+i
79wuoOCZDoVRO86DZOjdIahR81vjvtWlTqgZGlYjZh65nlxZ0AJ5Sv35jz8NG7+v
/MykD0jw4rb1lq2TMD9vw0OFwRtFQspmfxjvR6LIixxg2GTAIFP76TSJMm+PUeg5
54EInkry8gQIDkzYwSunxkv3+ZgD8N3SNxhYcEczAIwdRv3jcLTCPhrYAVK1AlS+
mNNkVo05omIp5fDkv9NeODHkrFjplaILmWRNy7PuoYL+4TYz7gPwg2W9P30RHbk2
cAaWcPd3an86DsSjKEHV0RtAfVmrTU51s8+o0NbvTAa3GkrerjhztyXs8dldSFpw
JZ9jAfjLJKasE5q3PAfnSMMnVj+E2VZm/9VyvDAFKuGrTPZMbExJwlVraVO0GYOS
KxywYlrT9gzUiXaUk8WrnZX6c5tD7XoFerx8RVKSinD/nbPcYhX89NA3XS6jUbZP
R9Fe+DyAm7i9pF6QGt+FyiUe9cHXQ0D4az3+UKCWKOVlrDTsALih3mj1SKh43Tc4
KC8AJ5qNUCXXqYaEHgoUzGumrb1+ZvdN7RVYEB+IISGz6WDd1Rt2CEa7J+iNenqZ
91kACO8Qp2Y3S+H9qvBT/5sUCVx4g0PhGfqPtI5W99kfWIqW+r5P2EDY9nODfFOR
NzpTAdsg7y0ZHQdXNwFVTI+3/Zx58OwYfj9C9n0UVVAIfvUwbctOwqO3bhLRwKnS
v9ozPfTn1Iz3Zi9qD8axakVNWOMzFqib3vMWPsoMUXHgOQ5kxsJ56cO5vPcQRTsY
dac50rWR27H7vz2WF2X5J6SJCjbaSfVl7o7+DJJ7IdM+9fDTlGyTWVNJGxwEKZUh
nCInvWyMEOZrw0+eE+cZJpfVwWliUOjVOxhx8RfB9JovjvemdjsGW6yDtGFxO1NT
gvo7bg1n402jcy+NP7BnXuWuslppAxmU3ITj2wS2GjXQ5Ugr8kOzqpngXQt0t/63
4hCM2G0vT+++iFpuIk08YZTRYseI9EGEO4Kv8xnH57CFEw1HYJAcSPGGBVKMgJ0S
Vr8Bu1eF5jHBrS8ueYaJGO2DOD9O2w82l2u2anjaYaZ/cAEG3FNSLOsDjWx7is7i
tzagka1YCm93ExlqIvyRuc6O5+7HsbHgK7LtY4rqbLQAH07eF31O3tlWsDIH2yXh
SfCHvjxRnYGr0EXiaPFBjKKvxl9g7rGwi05C5DVsygMjJiGv6wzd3/e6XbwZyPuF
caNf9fkzAw4Rfz/oP6iWgUMx8bo+L02CCT7yzb/H1XiVZmZJEeT+V9/AbnhLSFfS
VKD+PXM6tKmnWC5oMuzfGOzJbNVFyMTu+H3pfc2/AHEIfI/Kyz7DSPN6nweqIA3q
eLV0PbEQzTa0KkWvV7p6psGrzjb9mtdk9BvkvOCr7U1os20amAC/5ENR57ZYxxiI
/4VshOrgDVS56DL62syqak3ZoNE/Mz0ihU+1yG4sN7Z9QhP/RUWPWPdVRq6KAfDp
gD/qIFgpJnQt06CeohvZGuGpcYIpE/50LKnt5uX0cDnGQ02/rC/ak4rnUL+31O7x
eeG1XOc3Lsk2IMMjFOBZmhMQo24ChtlNzvm4lBazmpiq/4w6T3o+mUEaHDRyCa/V
X5JTbAWAhovRj5oJLMIm5mACygVdqi1RhiqzoF7KhszUgcD5GgfU1o8urm0JKs07
t8cltg4C15tvq5rmu7t4Rw0p2s2b5uXrz8xEropccXXxhKcxZIKAfxtBwZJ7HMT2
/0Nfgw+NZd3y3YPK11niX4ziDvZRykysTvfDPicWvvXr+hoT78TBc8IsYkg1F/d5
LQtvZwnDeW1Ey+CyubyDLhfmzAZsofCPcvHZnekJEN6aMe51DaAl8pgjwS9xaknu
qX8lO5qxnAwdqRUOmJpj5AtDFwJO+jRHOwyKc5760k0qZDpNqKs2BzMannLnqI6O
iNgl40W5NiKPYhLBrfG4NYVxDayEJApxj6IHC3RF/SYI3BfBrLf29iwQV9L8/WNC
KTvQvZ9XVNbfSvMa+8F5CN/LmMnJQCdjdH++8Z02ioTpNPB2toakv2owVom2jhuB
Ae5YYyS6NcdTRkEjG5NXW01DhPPeb83QVBIrfazKc8fxBQsfqHX88K48b2EDDow+
70waohbflqJvGASOXWEYnVjruwKOmZZ8iSuS9AVcEHZJPgUr5/5TYnMfqPEVy113
IaD1DFngekAkzPsRKmUDVhK2En3YoQGu/SDwnxr4lzmsy3vtWzghPtNvyj9Zw/CE
1xMauSVbCM6m5FKoQFElIk3XjCamHigPD6F3obz7CWpDfyZhXAsqE/2kEDYaajXg
a4hYPRUzEW0TYjevV2c9bOqHvM0fnxd2eUnnGY68MdDPY/c9lDSZR3X4JyUzRe1D
TQDhP+pLchIgkjnEN5S9B6TrD2t3noqlgJx1jzHYh25IHs7Xe8Zuo8BFW5FZ8bEu
IC5lRXA7NL/ppC2LE0OZKBe/NBTGIe81cH6XeLV5O9h+QtZ3DfoSWvCsgAtQmwbS
AMoPrjokMC657ttwHJ7YMeQzCsnRsfMg0SX/wqeJWCwtzXnwewJp2X1coCUo7d5/
pfjjpA6llOZajyY7jpfctLaSZ+5XKSSLKGskVgl4m58XYeqknLtEEMfnqYHdrPo5
Uhm9N/Z4bGn/YJevnC6VmNMoiB0VhEOpdFibpMbEW9f9xv1C0yg/FSCByKNEHgA+
Td8kYDJcBjIwvsvdAjKYjxK7l9kd3Mddu/O70l9M+gOGe7sjv+3P1qynKHpIRBM/
gDJ1K4N8oO3TPn7rnef5SZfq/6ylARe13LBZq0/fTa91DYHRcL79mpzm4Im7sl1s
2BWy+2K3pO1urQ9mZLsuTgaDRs4OTlKjpz2AOcHfOojtI4TA9cxsM4XjMH4brZa0
IHtWCmuNuICWkfysdXqr57stBT0hM3ORgPS8Iu7J5v89h9TEfbcFFtHSh8I2tMp7
8Wxwf24ZbhwyLxHD1UjPRhehsm2EgBFSuRXMyG8utqP4OGs/UMfNyEkwQ03p606i
NqkRRuDeC1Ww/W5BEtn0/9/X7i5FaknLsn6pVtBDlbBA4APPQKNxUBju9gSvvSiX
DE8+P+txjztltubFktbEIbnTlDaZe2J0LDGh6BCSv6utAsaFeuY/r8wlsyaE1ylb
36+hiDJm2QggYEDHLnyiqkui1qW13FKusMiHkirGqsl4ikfMmQgRauVTcx873kvf
1jYBPN+eyLYwIRsnxdfDF1/bYoh3uR5vAWceBkqqAxweGUJgDZqHzZNauCpBelE5
lhu4C2p2h9ZtLbR3XyL/PRwsCJJr7w9fSqh273GBMSkDIQhpp8eD3RKWPlom3zS8
PQ0MIBGZiy9tmtHQzEjoZH/0l/FBrpB/fnU9BD2irdxd3mHP2yOWdOvWTR/4jH3u
4QjWwqlp7F7gFocL+cHlGQoq/bv0iXh9FPsETc+v9rHQDw7wn46rbAShRX/Yi6hX
BUUBMDUInqrPLcLB3qSwLuF+i3hFVfYSyogut5alKtgEhci41IFl0FFLRfl3nKky
Rr5DDhZXQ7Nlk+C0HSt6nTjXUEQ9Z0YbjesTY19fOHDKiSbiYXrv58ORf03XNNI3
pDYxLaa+Y280eV7op3xnF8/1XcRR2+GCl+rkEmplOsPppF4XtsYrko0F2v9PT/vF
9GJsUo+1GNY/wv06v+/72/bw03wJW3C8zTonv6ImGRlivr+i9/HkRZXTNR754Qd7
2NP2PxgIvFwX6jSN0XCKyb6E9bLhNh6YSuRy0nCB0fl1IYqdPkRUPM/O2Rtt/1a9
m6Nxu8IOw5mDQvyC8m0pbyRFI6zOMc1lHjW39JXxa0tIzYYOJfjNXK6ndJiEqwMM
24Vm6gh/dsZt1djAM4IaJdVfQ1EbkGXSVhLTs6eMfVdSCHQDNnIWgOD1cSp/TQlB
uZN4bmPVYuqxmg8RoYADDm7AhBVLmhrDWR96ETSvBiG/k81rL+hw444kvhXp0Lh1
tAgvTbLye/ypU7rMAUvxiB3IunEaockDSkULyedx1F8Vu3UpVEPh5ApBjTmo09jx
aen4ZWaf19/jvVnvVYl9X7ylK4EcpnM+YByiaVuhh/JDx4+vWKh58W8L5gQHk5BQ
HV7scqRstHDSR/l8TWgrC7upU8jooUO5b9MizFvEZ8OzWKB0T6irljuIY0Sx2fdf
11FeFMP57jbDirv5zje10jvk2ve0u4oftOE/+tb+ytZkHGZaW3ZAYqSfg2f+Zfpp
8+XQqkaQ7sEBS6uCgDw/x8SkZlW+595CFQ357qEfY+20zxWrGW8JVF0z1OjE6qdD
BiU5fEUUWLYCKknKupVu7Z35vIBnRqhaX2tdqMLTlSwkSTKWWcdRUKURvXhFo1tD
UdJ3oboN6AsbjWZaDwq2y8gPqo6EJQ3E0u6ETxePboxskd52/dOZkVB4JLl2HaQK
mKGz4ZG7AwiBBEzYM3iqVspY7lccsK4aBFvQMvrvH0UZO4U6kvwh0H22ayOxo0r0
mFaWikWr6AnNSAVkcvk+bQjEKn41D664ifZDSu6T6j08idvv+la/SvkKZdMXHb6t
fDfsXXDUMUjP7ceMo13f8S0Y6fQCH3z82jkXQ/WvvwgB/gVHOKpN34A2dZ5TE1qX
yIxLepVYmtSjeBZSQB9UP31biGA/138eabG48T7CmiEJxj86P3eV9ESpRacE83Zj
ZMqK49bJq1EmBXDiKVRnsn2jWlQutkpjsG55EJC+inKtkpknVYY5nY2SwDyUSeOb
McYlQzf6q0202hfzmp1BmQTIzWL81t2G3/LQ63MDxE87oxBTSNGeJB9VYwCQJQRF
UN3tEzfWXmj4BSDMzTsgE6wVYwzdiNpJLY0FEIb2ZtL+bFMlZNWEghstJK0jVN85
18IUjrzLCyUag0GMmCFfZuz85iAgdkT6LzN6KEdn+gAv/1azOEZu3NB7ArcvKOqd
GJH5EluqQ9KOow4JvBTTmutkPhPx8ynMOfBUOv7ojXYUt/xr8XFs6gVqrOVA+Drf
N6r+2PrbGGH1p65YYNulRwxMLiJWR9puXjasafhOaId/VxPnSOWKTeEFHwJ9Pvu8
+f4sBmRlOpm+zwnRnPh26wrf7+THTYdIet7kSUoV0lBAdsZUI1v799Zj8F+LcUx+
kXKpgY+2+NOmdhItsFlokCHt3Px0yRo8D1etAKcEPgnNZWykV+4WlKxnBbQwf3LG
RIGnYRMZdWmy5hKRVQGoI9yRKuNjIFBqT4rerT6okFxpJvIlsrNVnpA0w+0NkoCM
tOyB9LvrzCoCDRka4zLRqqcMqg86PLYIoIT/clee4m46qnR2SrQIrXnixj4j63Z6
C3u7rsSMI4SvPijFAiRIJd8spIHSxEs0cteNx9Iv6MaDdcEqocfDbGoF/gLlugkU
757taJSco+0x8dhaNbMmWWjnhVXnCTCJQDs/jnKHocZhn6B5uideLvUhDF1+XvCY
3XFdAMgVFKO4yIAULYQzu+L1Hwklxfi2CAxaClRe/zW2hxl5oHUI4sFFgD7z0vck
PjviR+0rNxEcpN9a1QUWmD0pnTXEXwzZvKHHtXj8lwMXjDIwXTX9YrXyDUuVf6F/
hBFzwpIYjPiZIReRlQQxFqs8vXJ2ejclGaXnLcyv20ATPDX+rlpAR3L4vvcq75dA
/EEeKHIlhcg3g1ySSQG9KbfI3kONRnpkvbO9XNLfCLWZ5U/DUiNT+U037TMhZDAu
fuDsjVB+zFZoCTg3G85IHaHGtkzg9+EqusU+3+Mvu4hr5i2iDZizXMAebIoXh8ee
N32Pc+T+iTIDQs/BtZwsV18wcHocArsspZiiWUO95A9RhpVjcNOnfw8ey6mtfon3
OW7E8lcCjsIaj7yVwV4Ta6qIDD7DX6I+7WsH4FO+u2JPki3NxTiL05A72NkFFqb+
hPS9HWC9R4de35Su2aCKoatgQZMfL/A/DF6EPbRTqau9OLe8DUfEXcUv8kJFLI1s
Mf7wPs6PXn6A2DChD6tHxZXAF/Y3pgpAVXLhZYZPdr8gPCXwRHLqHzxhnto3gl0q
iV/7I1qZmaFc18I0CosbKFszXKUj9FsfmyTWw3uFt/sgC5z0h0EknR/b4FGKYiUY
z8s9FgBYGXDr491SigXD6XJOLlHorZMqYuqjh/qLR/1x0NU5+jNFIKb/r2CcsZt4
Th0Es4WbpOIVcFzphftwK6gX9I7+A5u/lt+ZpGsaAwRpohYEBmIjX98EpptYCJBa
soQa0LcVXpq6VfJ7hx99ayG1TjmcCKiuu+hwpjVAW6TE2p1fbpN4lJ3WQC0+bBT/
BvVtulXxdMIR4NtXaxwzJZH0vWLLvubNj5hXb1uRhZ4AgxIsS5WVrzeSE3/9r5Ot
mVdasGUMzoCdFfoYB67Pvf3dpw+mq/qIaQnf2qtK/lv6uPvVO3J5vK84jinNzCXM
BuObnb4nyMF2NuRsNKMXQ4viKwfFF5I/AH6lvF5MAtwUZwbM3ozxO45Dcb4a47LK
IwNKvIc3Wt175TX9oL4DgXSArsE0kBVZWEe1p+d7grR2WBg/i2ioGViNgnLDav4M
5XZg3YQJOOpTVke1MeRDQ8YMgyz36bmiEI1L/I2E22BArg6USu+duT9mnxQ69GnX
cYcAGDc9jpHgt+RIs76ZvqSr/qsq+NUmyuh2rqksDV8Yl8wXP4mJ5DBeqFnVAOZ2
7BB1VSV52pdfDX0AczdC9NPJ+o1LmjQIlKV2Osm4h94dfHhSlrPmFbe93LeJUzcx
9OkYicg8Gi3JNvqSh3ZfgQo0ysaxFI0JHIe+whNWDPH2FJEo6ilEjF/FlXeXfG23
AT2TjJI/Rue2FTYqc/CzV8rVeMyJmHoK3wULDmqHzAtwXIvswe114Yh5ulyYd+hk
QC3aHA1anq7zbnamlYZjg2Gh/1nZaJ6wWoMge89mbnkQicdZrSXr2tpBDasvvK42
ask9HBjHkDkppKbFRf+SnVmG/ge7wMRjorzNTvh6eor9p/76hhVZ62gE4YPWEuk9
EwrfpnI/E19KZfNFjRtLzwAZUycxO097S9wDMqNRdaCZo/n6+gQeUlybREQl736i
hYKz9tuQ/5I7qkqAZDwiQfXf0iaNta52xCg5Wn3rtT87E0WgS+vKOQXdIECMZYSV
6xYFMAK4HSytXMugv91VC3GuDgw3j/5cGoKP1wFpFuz3zwoADjp3Yl4nquMBWzDD
sZID92q3fzz5MPWqJJpMO+sM9t89L3ziYw4Xx5ZtBfsXII1qB5N+JvTU0Ndhb1WC
CH8aSJecrqWjvI0009zAnZLPttII8Ml+5VfZ61eP5Wazr0fK7loQko+VA6EdGrCf
G9gCQAdkgADPqfWnzJsorjwx7y00gQGG5iLWWbHffaJ2ncAA4q93B/qHDPnwDpJw
t/Kt51VLrkXPrNOuo9GEhwkGKUsHcIWNf24iTg2JD7YmXudFECLW58Ov40pnpv/y
k7ghr0a0Rp1J4fYSnJWZbFU2kzozvwBaag2MVQiwMLXtR996HedhV4iuX2z13f3+
iGsclRrYakNQzZospTws4PQW28ZrhZg0FF7/LliFFmIPKM3ELVvzI5LFhhzp3xRH
YyMpD8YlD9yL3y2vRA+JCA2yDnY6qV8v0WD5aF/WXc+YgrPM4+YcP2bY118Mz8+z
r0eSusqCmyagUSXKAiT5+ZnJjRCLcqToSLXjRhHUfkoHT/MVG0q1STIAT0xBPyhY
+AfAtQQQ72QH7PkJgPmopNHI3KVCfNER2ys6QNOaOcTM9EsTWiLRCxv7qMfXgOiD
i+bQmb05kfUoGJWwygxyfB0zQleC4b5+NGgs+gZQhyxByXUpEriDIMXZZwJXZDz3
5M1wpECK3OimsYyonTc97CGLK9k3O29JViit4J7SgeLKkWt8fuymxpCZWc2z8ezN
go96WwadsnXBte6DoirRPsFn1zk/5jhJbbEDsdxCbxcvLXu11k2X+/2SkJr7Wbx0
G4EszlZrtgMe5AfvHShBg2R0Pez9Y0+m70y8F//QrQjITozmcZtMgvlicHYePyUp
/nLPLGwOLRIpCybofIznV5aPutx1FuAtL4JVleM4lzuSUlWm0guhiYHVxJEGram8
E6xtH7evt7XyNvDmRMicgzLyZST3zQNyN85HSNW4SgZ3GtruJEvfQviMCllVMm4b
qN00p69L09Pi7ar1fIsTkfyB6RthUGU7xHVkUdWzdJtRe2LRsYCTsBLpouK2X8j8
Xoxq1TzA2O7PbaSDs0SGhddXUO5CEchdnZzq2wVRZ2oW/geEWNIDuA765jn//VrR
VRtH87yo7Vk4ycnLz18ab/P2gVU8ITiHNi/GhF8f8Kde+NGjfUVlSfLKRRqdutJ/
gXrIphwScQ4JkGGJx6jy+l6ew9lYucDmsFU53YTpogkuw9z2XN50FiD7r9l18MC3
mEi1EY0wZU9mIRG9TS/cJakn1EYASSgaSbori+lxtWYzaZTgkYkWlxxVl4hAD5Uo
pnAUVTFb3I3p//xayBu/kOw2GjcH7HgGg/YBjLV8mlGodcmNOvnr+ucwuWqxRLnx
CrgwCjcBadDNboZaQxYgj78xSB+nNqI1E6cskCw83gaxZBg8t8eW+wiyZk+QNdwp
ZnmRaGbO5CvWlwIJMYrZtLinnAEsoN/LBji7K84xs4aAHdSwkpwi/PvqupYGQqu1
GGBV+VO5kau3zBAncEDpiH3wfG4aT6FrYumzeUTZQvrnjP+W450JV9/CDMKYuHjJ
1lCfkjlU6iWAYszhtAFxe/fq0ZYoK6KWDpWYTznt8eZEnP6+x5VmGUVW6UpcjETf
qdtMLd/P7Kk98W5rN1FqpjWifdHcO4Z+YppCcGkCNnlHF7cO27vg5cBvBxSIkf1e
ziFo+5ARmjpcujbgs9VAx4gi3ZkPmO3D6pbzAU4esxpVmp265YhmlXUmoSPQeeTZ
uit1upjm3OiWExGNQwcoRvndBf8igJH5wwaAZJeY/RyKnbJ69fRPls04A+Vs4ALa
UbHXmguCuCih+zlIaZptn3wONnXrVmTiB7XGdhdaWNb+jiQmft/uMpeJhzK0Z92s
4eRr7XOfqDyZk1uyfkRtzcwNLoqgUbsOs0se59O3u96rLCiSivSWDNhzRHy8lcpb
s81hqoU46pV99zVE1EN15hNSUexXx+P69AEYmA8lvaDTDpiatfL1hYfCIgUC+bg5
G8Zm6lBkblNNu7PM/z02/FiSJoP5J9CAA6aw63p3N/V1F/ze3xKNPhrLCQ83lEo4
7HZ0zXoNY/0UYhI9C39zdHvZCinYB6Bl6XWkBwaawwHnCugEhKxgONfuIVSmp1Ko
URg67nTBGIo4iG1jEtAAZV4m3SHzlQVr1nKFjJwehBAcDisdtctBoUwyHS55esYa
rqpQp2APD17SAlnxMN1w9rsd9XBdlzRFFCD9Lj0471B5Mour5BYswys7F/OW1UiC
bMIj0+hmLmnGpGRq7GS0kgxmR4FL3PAq9Ri2D1qFBVYuMHd9gduR+ve9Sb33KG5L
o6q77ELhBfOdv1w2sTyugbN54E3SWm+63E64+TK2H4GdG25kjhgS2toxZevRlDJo
8Pz+csklgs3leGrU8AUY8uZSdRtFqTez+nhQe2MiIZk0sLtXuSSFD92BFXa2VGyc
QI5R2dTwx7ZPqDp/RTGfT/o5fJZieqMvY96d6RPxz5o4r9sa2umuP7Ni3xoYJLaG
ocAXAVGXcQOyKeAFSWqfQbaMNpZNu1m0Tvibperz/tkLJ1PB+FzMZcQdq19QhXlp
5Vb4E8wbpiuZgXKDwSDAYyMmovJfhafHZrx/xxyQcdjuQshqOWTBlyNjfxRQOXJr
q2fN9CiM6Ttwobqtmj/uPePPmGwVU9W7coW/HWXnyhJC72r2tumUTNUPqtuvtfof
jg7XpvEa5X7u+mE4cS89YSXmn5yYQt/HSzNJeI1gBvaOTGvPZGdDvIt5XKWDXsJk
qWuMKUc9OGveAsDLEZCtC5MkAoskormlIRehiiIrXO4LSwimg3TZXbbIem/umtF6
+l/maWHGWnS5slUggj7nHQYTP3o/5XrKJk+ytzzEymlh0pqzj1iv0OOVsX8hTmwf
jehCeJQnb4dDyBLBtVmokxy+QO2Fnej9KsIGjPIEXz9R86IW0N1YmqJyDmsHMXIl
PwqvG01NAM5KxZnPQfAcSjaIg7LEZJwLekLed+Ed/jQj+XCB2BhRCa3c4fZEZdS7
DkuH+S6d2aliuxqeZOynh2cv96M0BcAcfxJUQq1BddAkNkWGYzUqx0pBaIzT8p8d
3DJzB1cQFpBdgTNNIlkTtOf9A8Y68hEBQeCvDqJF3TfcEdsY3y7o0WmwORkPvXmq
bDgNvEXNbP76QFTMBMRC05Fry13n6WTKbXwsEnSjNRUVMyoVOUfgppIaYSsUoeYe
WGMc3yIGbK7VW6qMQDC8LmHlsEMvNXQcymuen1OnJ7/foo1X+PDlE1J6gAU22PHq
mm1b6TfCW+Bh+d/cn192tzkhz2Fgm0Q1x5hJhuB2ws+vB0vIqsr4BS3Hj0oDdKCP
irJhgPo4c4i1rYnNpNIBOkO94+Qjf9kSCsjpKSXYcPtKbI0YFYyz3jZLIa3k6DA3
oxLvuzlt5TdFhINQQt1k5v1ykDVGD+WKc4SZtUF64pCYukgx8PwEQ7ZEhYhkQdOr
9QpuCMrt7Bfm49lGT8N9Kz74uSeHumln7CFgOsg9lLt5jRk/98OZrOHuy7XUZBfy
rWRvnnFcGTeSemry3w1DRbBBDweaV/bxuNKsavDZ5J+QQO2TkIE63w/CEm2HMDMh
+neaYQEcyMQs3aG++nZrtmsSMg9m7mkxBaPXj70p24e8Sd55yBkL0OXzLCAw6AU8
+CYUqOaKuJ3meha9RYVKjzxbQajR2et2b7zlzR6U0ccfF3EJDZbOlYzRH1uXy0Lu
zHoMXL5JxXEMT65lbzRPsOKJAfnZl8LzqrNJEGo3jMOu3AyNbUsFIQxtWvuin+jb
+oKXtYeHN0h7UXI49Cu2TMr4k4zmXxnuSLq5DqUs9wfMryJX8w0mChn5CGRAgx3b
Xni7XrGp2UYXrxTj+VqcB8OG/L5LQijgehEFdOkLUPZucFqyp4o30mI0Oi874wMn
C7Sers4LwewINJBtinO2Xj8rCKuJDLCUxELV5j9H8IALb/2adJ5vELoRkHFqQnIj
BzNScXGp7F1SddnqF5BKAzOTMxReCncAbUngzuE5AjRdrIchzISYYiJmRQny0JnN
sY4GXKeGT4f/Jl9EAVma1JQYxNaMmM0LXd3dBj3TvpZwOE7IWH66Pr7D19XrZFFx
qBzc/AfiimG+LW3sl3DUlkTF9sa2gcNtBnk7MXIXF1/rnJyjPJr2artjLy+a+nxV
6U5pMlBgZATfQo4/5cIrhzizTnib3CsHq8xHJrD0IOl/oUOs0goOCOgngnxIxDkI
J/UOidV1kqNjnr/HjJ+E1TOd8JFPoSoV3GfaO+uCEgXQBipTvxAYT68Y2NgIZj4I
ERdsTDAF0rQwP6HM1o2b/K8GcR2sCmcKgVvqeQpQNhmC7B+taTS5PhT76C5w5Cm5
tgXLJlp9+adyG9wRISwWjCJJtivnFGRZSMxTQFbzB5VpYwNEIPxYQX/s6DJgD0rl
Ag0oKKy3bWpAlls2NuCeiDO9yD9QDllvx6U/LwK92vEcvBy1IGqHn5EqsZLFbokx
ZXlA9LcZezOXS+WcmiQybIlmtXFbquYxAVkzNkBtCSRs0jqbxOZOIG1FPLqIrKzw
EUu2SErF7C3PK/uSxmfMlfkEb6cfrnbp2TxAoAEC/egUburphwEtFLV4NDdBh9cf
j7TQjKB70xpY0ieFr00OcIxNUYnOSgSNQkhismIKxNcjhx7Rg2NI9Tl6FybK95uA
joC56QhfOOlbjzSJ3IL/x+i/HcWB/sLoCz+eg9dEy6NPzbvpPnYF78OcaDwH8Ksb
tObcWjIEmkXOj8RldbrgRkRZn1nar5atI64qCvWtx0q52pUD5pe1akBizmQ5GuQV
/g8C7KgOAoPjOwFfvI5ncZMr9uQc7t7dwdNamMydo8k+mMOBuZaYamvUQW0iIhSK
5ZkZvUqywbcViSQMRAgflMu1ebgEUUTlxviwCICQkkPWCpWoxyWnm+hnQA24qGXo
txdS7t12TFgRCRMDhIGhrgbX8za4pRrYnW4S/+dMTOdSHbyDx1B8XL9hRFEU+eGP
f14ZTrQdQTx8Jo+o0gPKZAZE2OKHI8CRbHL5aebnX7APDgfZpnMDAJzYtMeKX7pu
q7tF0g5t5m0A4KIEOpvEtJw42Ty+kpjBina7jxjsm39o93M7WEltptx5LyoVz4H8
+TtmPGeFF6yGyB6HUVgeLgA9IzE9SkZrpiulqJUsBFK6gwod0F1a1PqWUZgx2Ce5
T4s9p+qOkeyo2STxtCpd/IjG1TtbmeL9it3Wm4m3NdtUfi5ghjqRsLE+RWrAP+6L
1EUyQSieIZPZiOcacR9ZzqnTbii5um6jeqfnOE/ICF55iOGc61Kbwit1qoUDt8VA
TYtVzKc1thVKkgu9+B8iDRgnNpfRFSiDuFynBGF00N0uygIJQNYD/G7AjdD8RV/Z
3IoGx/gGREHAFK1dLt8x8tpF8h29jSJUJj+lCaOzreRrc8JLxjs3DJ0AnyqcsVaP
dvsl7uE2/AqysC4q+471UUQd1un5EOPTCpMhpimn+LNtwpXqhE89kJgBhri7gYhz
X15mpnplguU/IG9snjNvVx9P8hdxwM5rwLY5QLY3QBWGa+8FkVnxqWirBdi/ifYk
h6E35IBf77zqao35QeIMgEJtdbDgIm+8H8DISi7ekcMVkDaj86WSh+H9V6ZTebwA
8QdwjBh41NBDET3xYq4rgYYjJqrmwb6nxQacXHy6FfPoPt5ZgvkAAL0BcPLio5zA
1DrBBTjZWnmablxekaCLZeiCrv0Xdu0DtQ0S8jLJmyS8vZreefX/aThySQ0f5Eiu
jS1OQNR3fhP3F5ZLuwJxa4AL3tl86oLg5y8BJB8TGjU3w4mL/lsXv7t1Dx9r06g4
BTMsaEcUyhH8KljAWVEEIbcuEigqQZn+WZKFTt6TnGZI1/2Q2ae/IhZxlb3zb92x
RjC3g3T1eLsGUZhFC6SfRXz0UobSa3n91nWzGrNJuTv/Pm+jH+/vd3aJoLmaZzBt
MHoux9gUk4eQP9MkIwgk352QD2a8h3W6+6IbphanNACHYRmnZ691764RCoQkQ6jw
o7HqBJf7Ve8CN2TPzPcL+zGEIlNdDO8jN++LYk+f+ZkPqebgc9RgH8GRbos/gWfW
9cSlJEEw2pi804xrxjuWhUtPy2x7TZdOz6oaTS43ydMRIXGeUi1DFnE8UiIUcRRQ
QK6lVhORZCLbPKNU9GJfHvqzX8VR/Mo1HJaRaM9jV8vB8I2q9MiJArKi8ARSr/N+
V5ttNC6FMJYAmMCQfY9Ew9rmuUOzXM/2a+t/66iATrr6XtHHtiHYiV+R9pKiGSSE
f5xWyI9HlzrKnPq/1l4m/k5urDHtsCX7jRgsyJifgqKoUdVfYjO732Px10U1CLUe
QwUVGn1Z88TCPbUEapWrSKfcnPlHmp2ZUao0zMf3MVNsGHE0Z17xU6LUQT9EVOBY
QE2zn8IGHnJ4j4skiUd8eC0CLL+2g0eni9W9U4gXhGNpWTZcIfXEBGiMRznlcaTG
i4X9mSDj/Slf/mluv/8CO88PNHAkvex9937uveykuBAYBKy2VFlfLu65ObPadBEX
Nwie/Pd6z3AJxOAqRtPekE/KUH088siimk6D3WrGqqCb9MFRsxBKw3/AIbJ/rwCK
Sd7qHjbYeno8UZv4C5+ff9YbBv4m/TyAzIx35/2Uf2Vt/le3Ki/PCtn5jUF6Luov
7p+Z5CCpdF0QhimIbAGH/1otx7l7a2lchgZx7wZ3peiUzLqTpkoYrWVJxCbKN17q
ZQYptxIPD8RTMVJl4hwgHY0btiH97uynDSzuNzvg458Y6bA0BgrTiXJBJUfHGwsr
sLwwNk6ycIw/nrHiVfMHnRLernDuLZzVgzxSA6P+jPz6HyBzwTW+FRSi1GGZTcCl
sznE0ghcfkhPjbTOjKTL6TINGtTTWtDbVQx/MMoP6Ovunj00WO+6z5p3CVC+QedV
/0Z35RuXLH2wkelIzWF+mUasSU3wCo55g2jysjSDSP8oJAF0Ft0Wv2mW3z3gH3bo
9Kor/6IAQsnmuKsUDxdEANhV6ja0LGErhciRpVkgWYLpYOg5wlq3PBUV/CBjjO/d
rPMBwsV+YOLbk2mOBmvEwdUOAvpESY4wrs1MDP3CYSfVN03BSmoA7OiG4dyE6vdf
7RDZ4V+sh52u3udFfc1q+CRNzb8kRTAw1c10E1Ttdrdz0NK/dgbt2+OEFgUhh+xP
sLjP8qQe3Fd1vKJp+LoSzO27OK8fn6EgUIrQE55UVJC/skOCFaw59mPILg/oftSm
IHDY0Xtz5QKBFwebR96sFPYC0aOG3O2mG3NA/uSs+EUcOOwF63YCX4ZENKc/iZHL
9+sYtpKKQ5cB6QnP2MrnEBGs9VJJfqldNhAKCRJ1CP+LlWAKxHWvjCZOsZe6leoY
Uyw8+SN4+5vxcZf1vYelfLv5mAZw9T/e6NxaN8BJS5GxKFZxRqt92EZiLuym/8PS
HeJc1zf5FoT7ETG/bPxmO6M97I9wRGzulVIaJr6mdv/MQJJiiZFmoDFfZPZfkfA7
vY9h4GpBV+skEjqcVojJdLvt+WN7OcvDZBqvHjxEDYZHbxzAvbs+ckcVpiKiYPDA
FR/55EsSeqM1m8rCKbzOb1BBW0azhUeOkCrghriHJ7dYINH1GcYpe72+wyjnxoXU
PTVRGpLDno/9eBgCVz8tEnvlPpNUm/HzUsUTP05RvY0f2OX9U/aiOhqZ8W5ppFcu
b9OLqktmHy6FQf9vHJe5SkVtjO5AVk7owtbk1vBIma1R7BRNA9xquVHvv4H8H6PO
mlTnRBzarjsaGHaDWaWHzs8qP4Bqe7N6vXspr3BvzAi5SnRM3SKHHPDg3djf8gE5
8RrCSkI9ZW4jNz5lhTPLhiu+TvcDsKAZzJXDSgOq/c5ZJhMQY/DltzRXbuVLswI+
sHlabSpq0ikl309MxziJp1EN29hMSohrw/utGNFS5CeYVEThk7mpTAkWBHsSYsVs
60X0cHB74QQu9H/IrNWyCtOlCn9dDyLJkVXvzPFoIyAE5OkV4xMfGswAqWRinX13
uhXoDCWzk0tytlblvVYHG/Mpt6zFB7uk/57A3ejvWOgThcY/DpnOII1vj59fJYVA
+8vpTa21w2KdYYFH4hFL5Aq1yshUc8c2+jLErl8Zq2eYjXtN6fczeBqpz8a345jT
F2DBGwjq+9S0xxgxcOJ9V4HeP6+WtahO84GeOhxL2vEL4RGG3QQNy3HcKkufk8gp
jmFMzCT7iczkYxrPR5yILUnqz8otEf06mAYPdVMeveublAo8JeneCT0n6kyCPErM
qD3uAW+7ZqE6U3eNYNRwIQcpGXH+TsYfbeHDwlY6k2beBlr4kv5Jr0gt6hRSEI8u
XcbfPgs+3Rbmsis+kj+sDmvjc8dtbob29dp6PyJJZcS0gy5VzB4ufyo2Z32nSg70
JAnhHPl1yjsvk92ECetxsJcEJwKv3ET7t/nluEGeVV+gOh2NeSyXIljV1iXlLEQ4
8ptxUVkozY2CeqTWnAWWTvR+Yb/q/0Lh9OIp/rTkCs8zlol3ET+hnhymUegCKc2F
xyljs4IdrT5iB5dyForKCssogT5zX/rAZDKnpxygtad9jjMrP01wI5hB4Cnmr9yv
wjxLgNLmN9+XUfKZfIy1QRjq4TsdXYTq29QmexDMSa6tjUuiC2Qm/jMzGsOtiCQT
2uhyXhlQr2+UMCah+qNHHFtsckxb19NAlcsU0kZKhMLYMlQGNpYV8pOrikN1Q1ne
fqAJGiEyU7easTVtcku37D69APar7N6poT4tXd2HRoaAw3GGTYlHYawZ3Uqob5Zk
fUOIhSZqzej8xgAmv8C2IzQ013Kfe4Iu6o406KQ1p2m5cR5EuBLVUo74M+U7AUBy
mgNeFE21rY4HICebsTK6TEX5pRhQTPPzcdHE/xe+H+gFpancxdn8qwXsvZdCl8V4
BzUOIR2cBoNE/BcxCWVODPK6DsC/zujrfxxE8go/Cz0ZFNvWaA5LhT3DptxVzOBk
Wf3nG+6Cp7+lRXDIuLu7WH0M5WP4nlT+XL8m+n0bFDsgp9/JKVXE3D+74vvHD1dA
sBHohlezxUOS+tip0oDkdJPgwvFmLUt5EOVY0O2y4bo5Gj4cqnfcMcaTMPIlt1lx
edWF2sUWnB3qNoq4uvuXnRx6zEybR+hL2IwWaiOxobH/1zNvkWcio0HcJ2zQUzlm
/qvCSjmUr8hyJnIXBvQLmHBsKIjKLFw+1unnjx9ACy/DzPvCOSKWy8U/0IVSdMpO
L2q9k9J2C6nxbV4R1n/jlgEPVvHkAGvD+arKiPdP8SF0Xgq401TLAW8/HBf2II9M
y21oUOTmi7SUODnlaGM7bgQnGCmaKmIYWjLik5SQlf2dIpQp39bn7scRzFwC0Zkm
Fj5mwloFJNDuxqBr/uV/jwI6ZTDySib+CoHBXYAQttW/AsCL5uJPeyK9GtGzJHAD
1UYKgV6EvtnarjbYQu+1L6miV8+U39wUGUQUKIw88Q8Jp+ifFitCo/kq055K4aRN
OtgqkcUVh9BqIN5Ejb65nJkMIH1IfWyKBDip6NLMPKFe5yQZdq7oSHDmPhxbWnsW
kW28+AWa3Tkao+/qwEzyyMzPpagZeB7dgh97Lhmo31Srp5W8D/+ZHAWN8nQeojoN
xnER7oFnPTLPDKhfueKNmu4twQqx4+UI4J40kC6b4DwGfUZVqSZgO2Lf/Mot15Mm
23FWlz4HwG1CwxPEaT5YfK+RJlhFeLxydS16Lfd9m+SMTtXzeL7pqeYRJDgTS+It
vpmzpBDIJdBAbl1GA1/eClxP02mSECTi9YcZO+qKJ2cA7iQCr89VCbc68ow8QX4S
TPzqIwIsp1uw9fF/6I70yFvd2U7dEzO332hD54fm6XQF2S6OXLBaRGgo1miLsFvu
tFQDSLbZ5k7bCURvniaftrg2+yYHayFYAO/5uM/ZJhnsWUoWruHQJfpsnc4uSkhe
XJI1LkWv++rvI2wnIl3zNkXtH14Z0D98inO/Tg2L8WGMz3h1jNtQtyXNbCInRI+e
LY6v0HRUuI3GEODpsT3O6a0DMG3b20Vm2ZC6TQ0yWHvis7zCa9CRZbrvC596Ze9k
eFXt8Ah/ded7ck56/ieBju5P07Gzr6fNlKcMD+ZstLbsdLbnFqn5TYYrqG9aH4vq
OcErj0gG5CjWktzB0rH8oU1j2+1jeiOB2plUDsrI3olF+E8GKY9LXfGk3KkpCr8b
lFTy/FNbl2ZVeYDof2ZyGf3SJgzgWTS60JsuLzbt7n8PlPqlJB+gz6SvOZ7NOH8z
aA134THUvTmGfsIhOP7EwjzB/AEAJ1niEd1ZuuB4+eXB0BsVgIGGhza4DRySQLC9
VNcjPH22RvSFtY1Lr/lcHBnbSDfNEyu+2E8/q+DSRYxUPKU9+Euq0Es31qfq3JCA
mFcv/bO3jvv8iylQRJIflkFcvj1HoEyWVp52frtHfY3nVLFA67q+9bCkObKUZi21
LvYUAHq/lx4sKiYunxSXX2SVHn9XMG5X7UigmPYzGk17BlvwpZHaShLQHYaLF/Dm
lB7t3ETlTZTljpX6mCzb7c1h9dV8sfm8dCk3hdzWuu665SVITYuAQigiJJ+QKRM0
SP+dcNp+20TxXqDhcK9CZhltALbc4m7yl/pFymtaZogp2hu3sikpzPQ/4+/a7Z9v
EGg5zm4PI5mS0o2YzF07OprITmiBbbpp7xzJuBkV2eR9cdfIkolO12+X0Ujv2agU
eDn5Lj5xwolz+iYbjmEkAnL9rTWClsEuWAdFIeFfGuY7qtOP8bf5U5XGD3ZJlDP6
xWRRx4ozQDd/uaJtJ66vf9LYafRtTeOZOsNirO5hLF1NW6As7DqCO2roq3cETjLC
WE2GRhAlRHAjPreFMElf47PPApGp6xqUxuzZP+32PpahxzkvsmHTzjSUXXaF/9ye
Pzu5MmYXk7Cu8eth3zONglRY48F6qtK0IcYP9vSValS4JRf37NkNYWIkbGbH5oNz
FMb4Ua3mAAkJ5as4PaOiAzlSr8aglf0Nq9G2Vi1KgS7xxioUj1oxwYXERuB1JfAN
y17W3rzRmtv2x6NknI5zHgIZbOhHObh9lGAcLv2/U2GeK17AwvtzHkyXVjxpEt3+
aACusHRuDNibuiZyK+JwZUtcRtwJwpk6qR8aJMe0fs2J/r9heSI7jVdQuCixBTDF
KBxaIyJf8Z1o952kcLepMyFe/RKyUMDDKL/jow+etTfIE/v9cyFBq1IF83bKaT40
wEHC/EG/AVLRoLWyo2rG9SAVbY+mpdobJO+PK6oya22pprVIZSfvZrRz3vgsJ3mu
ema87SsQlqzWYr7+1J3+mpJHfyY2NE9eXlMHmdqGJWDfn1DrTBrJDiCP74eXIJAj
+qz+gpHW7mAR7Jqky+0W+PgTQPFvDnWin4yABy4CVy3zCjTQn8Fg0XngI3XnLb+s
QjWgsfVYSPjI5nAK5XIma160FWDFSsgAIEbr32w4hRGqwqpkDc65g9uuNFs/pwQi
PoQGsdHpivmXmhQSaH3zNtw3/mJ8hJ5OtjBkLswb2Nqu0sylZauQldH/Md6tJTlk
VeRaq0ZR4GBWvNUrIkviIwFT+eK9PagGGho6QpbuSe3aD6hUb8ydzK9Kv7QraFDA
dJRi+tgmCbhXfXM4/8JA94TlNTZICigKqNNVeBbR6NgrXa0g6T9NolrlcuQgn1yZ
5O9bU5p67fxqm3eXvFPYpOB2jbqRmq4m4SuMbdoWVDP9kyWEFGcCEScIEUV7DfNU
PD+SF0vYyJRZNLoa/7hiZV7WSCtJgB5zYVxDpyYD1LtVpPiI6IalQ0vp5X+4cv0Z
6mogxzYL8Q50yVvs8/qKbZEavd0fJO1dy1YR/tumHJSb9wlu6D2qS1IKccDoXps7
2cxKi8++S5OCTpXOOGPHJWS97fEvoiZCqg4mTgSqUvE9n1ybC8vFP8OqiFV8ac+F
wIRPe1rkxTtiLjdz8LnwMSPXcDA35PbLQRfx3RpkCi1UvePqAGynR3ALoMJomFgQ
/1QcThiS7gUqrc0bDbjOeffLr4732jCzNzwz0Hp69lJAetUYktXg+28pw2cPuJjP
FheCY7IUQHP1rLVvG/KPi0Pg50cjFK8nMVAj4zs1MKEKiBEKhO8Z9+l7lKaJksf8
xavqESwPU1o3MOSgi1d/C1vZuWUj3kuJMVaB28KWS+w5KFYSZdi44MZbkPTdUtbV
CJOv/p60ZK1zGW9yi80HGhLyP17Sp7TEAVuQmE52z8/tZAd7PWfkppDZqr4RUWzd
/5kfpnHRFTNxIGNV5fLPhSEVoiFvp9GXeL2hx8d0EAKkGYOPPnODZtGgN9vNuf6g
P4hWaXKSx3wzp/f9NidxuInl/rmBJIcuct1Or19gd2cOyaT2WYAw28gpvj/nWeG+
nqq4xNoiU//igb9WJeYR6y3ScryWN/I0ROaQetGRBMR3s6RYQxQCFdzBN4BLgd+H
0aNpW7KYs9dr9aCeHjtLhKagAegRsetyAicBsuI+me2NVV2EOSYz61pIEbO6BdiM
BjAvavx3gqPZtUub9MdAW+BO/0SaY0LEb7DBIKzHElXXxAbKRLFj3FBbcXnU5zUd
hLD0sQ1x4z/nSZ9YlAtjV1ZEUPpLVnphglEXTBOvZYC4Og0vn9P4zEzu3NwRUH9q
pBZ7Hgh06+oaB9MbFJHPNRA2Pa/3wRS6AT4CORvL6Em6Jt/j2SSwY7mKxoApQCTV
LafR99dR+2hE4hMQt53DIhWK2BoobrSXZv27ZziKNji/JlNukGshUkrsjKesk//v
K8BYc7TcFodURPo8vktsJz4SLbz4IpzOAJyvTvlJ+opS8OalmPr/yxvQaj+6qjr8
AoeI39fMRZQlb8FhqziPdN/6B8Kf2bdYB2y36/8sZvMM3RB8d2U0ih3frv/aRYvq
ny/QoJUxFtqvn78tw/PNt5bftHbCssUOx2kqO1wt697C0atzLCExKjvQxHgnDZsF
3cyok9sH5OdRMQ7n/8n0sFKGCawv+G7NAaFgWXMImAPxq4rmm8XAQuy39L4Al81g
ZW2yGCcaxw1Xr/Cuxh/Mi36mf3FyCfrEbQT18wwyFA9D/0uAeACcuEOVEd3YW1L0
eBrs6FX9Cb/FUqgUEVCSN7s7UriDRtF0AWH2gaCHqYn11a++q7uMxhiJAY9sbzvV
9E2SQQILDgRUa8Tlw5NA8JInqfKQRRBS/0I+6gi7oOC8O+IUzN4ZB5w1riVj2ePk
hamZJOjP0K6GLtGE8082BhGN9cCLK3Ks7hyKAihpxdoFX1orUQJLYo7dnEHw7ZaY
hGLJqVopaNyt0KGXJX5hU3R/ZqoyM3+jbuxZh/3X9Fos+RRhlA3hRBdnizZ6gDSb
zUXZ9rL9to1F41g8vsNH+OsquKVGzM1pTW/joj8nYZFgFwvDKC4nkkE5vf76zV4N
DnPagk7qM5EIq2ckwYepMPOzYrQR0UrH1AEyHcv8NC98Y4l+wj9Z1Q/E3eQ0GkBp
QTriXPjkvNYfeBpvVoPjfsC4zRkbB8E+irii44OP01AqvMn/h0xpWPkuifAwhlKt
jSfiZ8/IMK51+JqyxXfXX45C6Tu/rK4SAb+Uu9kEIDfBDXs1vBhRnGQsUPJ5EHlx
165jvLbbZb3oyYUznP6ElogEkdqoeInpCfn5HyytrqdqJRVFSzZ88cFTUj77xcpF
TOIJCLBnmF8aIvzx89de0SqtRJmsqI5qkV3Ycdn9Cnp29YNgm3kAaLy/LywpPSnR
x/U3UQtCw6VRs7s4nROTOCxemvAGNyACmccLbpoTT8HxcQkKOQH4LivtUke0e3Zl
Kd+EG7t9fo8vBwBONY9h4jHPrAaKNwnaGRga9LkRathKvo7y6KpL8IOk65bf41Rr
nTTIKxmzr6Eu3ylu2DRobBs+AbAzUYPHMH8JJyPdw7FOpTmfgeUEM6Z4z1Qfw3q0
0aRvAAE9IB0XLytCohzzphOMQxKRR53a4Iu9iPN/He9lan8cQJ75Gl0CysAc9VLD
Tu1ZvhUkYmIAtw6z3ERmhUxgcuYi7oLkSPs6/hNO3AUO6lv/NZBMxg9yo3zgaQcP
N3qjVbZwlw5iNawoRi7l1X+t/Lmx17fJ0uCw6h0au+vJ8LtoOoB+LuOU4XN+Rduf
kkq3X7jtGzUbRQVeZ/1fG5BUECQ7uW7lUGhNxzWJmWTRj8lBtzWR5pXKkw2faMtV
KD4e+wQhZqj6rBFi+9lJkk6TOkwQFi7jCnGw+muHprO+VfFZuDhtUlYSsdETCJSv
ad8kC0a43XNZRAP/GGIH+cXVmhBDMSdp2uzgMSnhR8JQQHu2SnmHzpFlk0uQHgae
9YOT/d1xZPoitxohPTgvfNs19I7nCQlCjVfvn4glY3IOyL9RwcxC6M6qbKXSCSR2
MCayaMGxYX/VFFIzswJWRGopTwCVlFuMah9pDjpf9uHMcvAWtu/4i79G2sSo8E24
X9WyJZlAmmmOhG5Sb9d2MfQwdAjE4dzQ+y5DqM0lTckzqBtkks/x0ca09A9ppfao
da/hY1gxV8iveRTu62iTVxJMW++Xu9fk5AKZfFREyeE2hsgpr6tfQ343vPySdP10
GiqjM9qi6Z1YkNkhn2T6Se6q44TMiD4vL6mwIoPxXGK9fadWL+sKKbQnxgMmGjz1
34f5yZQipx2GGMoLcBC/DhMzHSJf1JhQZfVmPXdd44NjMJZitYzoA6bTHV6sv6pm
mv4tU1kNmUb0VUe2LeYosMjcQJwip4fT52fNrEuytVUV9rZamagaW8rdZKLzQ/fl
TZf0C9L/J5ZQsc9CLqeHByEIHQQIXu4DbjSPw1BiwJR87bvDT3ZY2WK03iDoGg+2
2KEPVenFW2Q3IMxy6iZKahh8zR8lmxKWttkUf73uPHDrJh/KKQ4g7fy2NdAQBgWy
/G7sbWVFxOZjSXasB+iOkA0QHiPjTFuYZIr1OZmfxlXuhvl31jb8F58KglYdxFh/
ezv6UWjl8pSMyDBbxCNVA5M2BeGCWiBPb9ERoDaxbmuw00nFvnrD11MrQkBPhgRC
8lItH3AbOq4S8T3zni5Nl3fn2+OqUuT6f52f0Nko04ko9Ep/jLT0RBmnVU14jHrD
ugWxt9x6hZNITYC1nDNYR4qIyWRlPb5d1EJm3YPt1hnaXLMvbojTfrHZH5H8tK7k
yzuiH9pXwT3neyuOw7pkKwTiZ9rDz7V8dciIxUE95j0AtAVVzTVTrcoQBP+TkLQD
eKInCzFdGuXIC12fJgufiTMRSb+Un//relxfn24lKHPgOAYoHmv93cDl6D9ZBdiF
wyDHWkvxng/zcOI2qhbMe6ZU4n5t/MmMc3fhVVBwpePZumRYaGXYTu9XBKG+ulIv
Ky/hx8a7OxE6uWERFa35x1apXA4qwGspDHFloj3kUlf4tHGahQFx+N6A7YRHMdmm
Of/Ca2l6hFMtoE0o9hycG2IY7LPDviWfghmKeQ/LeVplHkT5f9NJpElPpGCPXIAp
3dwhBi/ZL0srSWcwLCJgjbGvNBrF0l2cpbXOaFjjHJ9Tcv89TrXvtVF1ayt1RHGt
HpKUm7J3fJAJk/f+pmJgY9ZbRSPk1JbbIhXtJ6u+Z47xS2JfH+OxOkBBXOa41r22
pp+1w3AeC8NQVB7r2xd6Rmz46co9ifnbV1p9kXr4y8HNhoZmeL77wVbRQRKhCScT
56J+S3b2NYPuLYxqhS9221C/vEaxKmyFKDyn2jMLsqpebQaOhLpklhJ+w5yLbrQb
j/IMUj5zf+Nv7tvrzAgHnzaEDI54jmQhm/52OXIJNZMxC9IivfRrG2VL/a9CJeiy
9duQKdvjyK6NuosHvUmlP+lvb/e/5I7lny+OVFfgpCrAhT+G0KbRCcNn4WO3E1JT
u0qOS5fJnkJRz9bURrhbX2Tope/mscx9XCc0YCEapeG2NqBZwes3/Yv5hAswmVZ9
gfYCDdgjqt6F6epzy/zQilXN2Eef0xipfxRqZ7uGuhOg5Tivz7Re9DxoQO56hAaO
J2oH4sNifRTIv/LjBvqWf6NpjLKt5iZDGgtSaFy8BLiNOfAoFvHTBKp/UMqVdVHc
abnBplRgt8zB9lDKuJJUuHTcKUjT3y605oFNDv8cpZFrR4QqeKPGPD/qDrCxdvEN
Z/WfBOQHumLc5xz/pAIVG0h+b4M5rjAlm6lO6zXJyAgMc5Ht7OmflFLIfxe26JbP
H+/NTorRpb+tIDMOhyG3ZXfPvYVy6HAeyJl3sOGSyUXi/0iayL7quD80wcSn0c5t
znvjvOds+lFfqacVILWYunGGjR1aOARyi8wssh07sFFf9xv4pN/GhbEkYyCPhYRS
0IRl6J2LCPAsO4mS8GxerqcP0GSPHwnaWE9uglZkQ9f7VRpApXEamKoV6rNEM2JV
998M8C/CAr6RIbe0RrGZxfi2vmZBgdITT1Z84zisO+tkawxTu7cerIMfbzfir4dU
FrZChbs/ojvmekFH/uBmrVgFJqyNfaZRM36zR59z2iZWOgrOWavuA39ejdv9D4W2
E0FIewYgaLJIzgMsNqMvNK/M3mAOzYjkFB6rJbeMV0KN52nOCC7AUnJu7j4iYVuJ
ek+snXZ6vJlZEOKl5UU0LqGieWyMWOSDwFeI0U5sqxTuUI/mJaoPKmBwE7KnJm5l
lwJ2XAT9RqTe+2nWC0KVJbUyhPfSALUdmX/hqL1XaTc/xKZvxjMqIqB+a6XWWCSK
xN+RFkxAbzXXSO3xaXuhoZ75QNMpWOheFrS1PaHLFUcZ/mc9X5UB3KOTf5D7CLlT
4DY2SpSZ64MKS1zBjbGnhZKk8GUatGikXdToj9LXLDY1F1sHxCbiAAMBhEuIy6U1
+yzBtpRPVEGBD29UuAvtyhe44TidX5chcekgVosnE2cKBL3BgdrzTLZcH4gOXwB/
n4FKshtCM9aqG1kHos1q2jPtYEIeXKSkLwu1djLjFak6S699zxIUsZbjxwspEZwI
XQoxds3y8lC8VbKwIMJB9BsMVD71w+t/uUia6zd+Hr9n6DbLwA83p3nAtQW+N/tQ
Fk6E+KY8y4gW4VlTPQ0W8aZwn2SNK9SQmfg+Oie1N/fhGZvOq3soEvpJyQuEqtLT
NR5aaec2ly07ABtdbPxIax4GmPqLL0JJX6hnmnd87csu7U9uszyxiOJ5T4nTUNmu
7gqH+3/j/bqajjKhCRlwp1SiwP35yyrqfLefK4pbHY6wuoFOfIEcuqlqY03ijDyw
+6hzwZZn0OEnEEcuHFultSklkm72F+QsBghtZy40y7FWG6j7+8oVuvxa1YjbDzw6
9IRfldzYCetDLlUOioeYvCO9lu/RdVQshXACogSsnSsu8+HbdN+/pYQAJJBlv7CN
sm8pqo1drz6Sy8E3ShrdTF9J+rn7zNZVIN8VnVE0BIWD3WiimY/qvVbG7/8ncnG0
yVhKpaH4AQHRq0GkMWqK6E33hX8wJ6zNfwFk5GIRQvK1pgmc776lAerkZgrrBa3r
3QN6ARFEiwRSERUCm45Sj/S6rUAfBEd1OmkvKCFL4jSBN52dm9Hl/DjXFuAuB3eE
FIysCEEoHBrHxOsVQjJQ+ZyXAcq7omjAkAAoCEL8pbCCt3PsuC6VLuB7THxqvboy
LmZbt9oaCYF5hjxSFk7Ra0kTkb1E5iDK7tMaxyVA3BRXwXUB5yPh8SasahphE1tu
GActgNPLeHG4xbdB4qnEKecaBDANJhsbCP1kfQYpCSrHLUsJnoBwiIpzNAF+D8re
t+Va4HpwoJsgjtfEbz64NpVnQIIOZrdA3CcDapxPjqR4HZKAyz2JIOKCAQG/A/wE
13M6ErsQdtLhZOUodeb6d7iN4mDMvVXmu1dtT3PuuwYZOsr6TZNxK06+bRC1bYRk
XqHA9lm5323GRBkWyIplqZZ5K5T7fAltAmbra3Yl0UceSNC1n1lqxi7mMgKb0f+j
eSKo/x1MUkS2kY0GQ05TxnpQUD3jg5xGAFGFFixFswyXeuz+YawH5Y1Ls7jSdn4/
TE+Z4oGz2hc4sqhprmHF5tJ9Ujj8OvODG/f8vMX1W6APr08livq+sGl7OIoSInoU
JUQjdV8A19CPacBnwD++8LC7TgpJ06bDsYZosCuxG2lA999SKLYHfxBj98MtQm0s
mGGgZgs8qbJd1X9PDwEEeo3lbJKeK7fvgBIRsDOCvnxeoYNHGQXE8oRp446frMT2
Ay33fACaxvoSZDWgmuILjfrvzwtmyy/+JpeP1/qhdSuVBQHFo/23nYBg4umYNIvP
aNj1Um6+0wUl/BEekH6OFgT0ilGxcQFsP2aYLQLqbXmK+f85jRrevMxVvh+FqP53
dA1snChWoVoBC/giwMb+m0a3SeXoLcdvnXdjHCFNycmYSlXrEx3/oiXZPlw+P1k1
15WeuSYlXwz5ET2ZE+W6LoB2NdpJpYHpFVMmpTopRvbUnmWzD5ukWQGIaPHxX3ts
tBGZQZNDeRGTLEuJHAxJNztRps5H37tGY8Hc8N/+hvcBaM1kJF2U0ARHgGZDABlA
Zzc1FfJKbMOItbPXHtZmKEFcSez7GwRDO0hNVoNYNQmO665KW550ZE8BV/56vss5
RJE+JlPgbBP5AIgQW67JaRJ5n4zc3LZ1wx9MBuWXXLlHGm9oGKsNnGGNPLf9FCeQ
eXIO0InEcrjuzMoPT5Ni/PIRps+h4/8ECaQJHC8Qx71ZEFEo7WR993Q4TOACdrjC
0DFZcvtafZMVJXYTvP1ANxh04w2a21Lm2v4pbauFeQkoJ2sL0vJnnsNFPzw3JpYF
nproWZL+Fi4bz2TW6UOvMXAYpdqn9+WQ8DiAktPLg+Dby2CjkY2nuFJrD80HS/iy
2tcep3g7SpcVnZY+s9+Z/mSaxZeXg3Q+U+89zT6gpSWF+GNWMHcEG2Q5I+reVmgy
aB4SmCW1oKTW1EOdlP5G4QF1NV7tj4cT9C7zazvMAygmaIypzeTf1lEfNVmGkSQc
hy9M4/ODC6qw2eD31j5GOYW6hGEij1/SM3KWGZJSmBzSfEgUmOGV2zhlbW4lKxgf
8bGK9yH+wj6L0LBSjiHzEDP/hPxFMZlsytT1PYqGJ2geQ0ItzUVUyJjnaU2Zchxe
GE3+dzIdBo+c4yCFXQKbxX//OTBvoPtHaon059S+nqQ4wPUojC8G373jIPOLoevV
39UtC6RPm0IbsMRi8JJzQ5pk9pMk7DCi/XsYz+bHb60Ek3hbzMS+V8qrXlH/ZgvB
jCUWMIqYPEeQ+JE/F0z0xhOS/oCVYUCxpxFHLADciK18HR7JFi/YVeiF8amwuKJ0
`pragma protect end_protected
