// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AGaXlftmutxKOULwpiPUZYphdCuhcplTF7fteNwynmFeNR389GttM6zvleQoY43W
t3uJvi3QIT3sIe9Oxd8VFemnEzuWv4ECI+ELu2MTVB2p4gpwZFoKA28r0vxsqg04
PJgrdodmfhhfA1VwLARihidg4GU1kQdMF20WoJjXbpM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3232)
tm94Vc+VjVVLq/MNf5sx/VZc43EJHVbn/LBlWA0/Vxu2ZZrrIrX/Q4m+E9ltsNeo
d0zbfV0WqWh0I/dAq5sDVpJaN4pOr8zsq3n2jKGUFtg1FoHhf9w0cft6WUFeli09
Vcz7FMaYwFsvF3cG2LD2FFKgQzt3r2IMB0rvgBnFmBK+W+Cf9+GTVvBmeMy2E7V0
h92z31gL8qv1mWa7H1HkGeOQ3X5Z0tLf0zNuWW9Zt/w06Kdf7l6h3NaiqfJZKxLN
QWJ3TX9m8sWC3FpidOoKh5DEjWcm0ynLT8f9ApHMAgO6eHL54jncT0Dne59j0wHn
n+bJ04XnMlLnaSGIkpQXvmTc393//FVHoqw4t7HlxwXEYktQKG/jW8DJmAOdVcDT
P31JBIKo9B8Bi96pbzSQCJOGS3jjmAQ16W2by89KNkqIPifpQu5cxiuMBIL+GRV4
h6jzRODxwjegQPqk2FTuSzhu/vjNj/AO3SPrRr6X1UOgpUZt3IpbMQcYs6GGipuO
FtwETjK4/5FB9QVtpSJ1RCN2y6jj8cM0THhjAUWH/BzCuS5bZRmxrGB7aatvcXkD
OyLFZEyhOiCeD8hNCjrrM+d2V2wIfseIYTjHbtestLK1iw8XK4awM/t66D48tK+E
IvGUtoweBkpU7lizssH3trbpfDsl/YGLvVYznXmTYHGR6c5DUyG0/ZB41spPBJ6g
BGas/ts8dja0rT68mqTmXHP9scOgcdOhxbhVp1wZpV8vdvtMSi1qxCwyFy/33mvC
TnroHh16ylZPMgCHeMu631z9CjJDAGH/TxbPm+hqrmR5PykweEvDh1ZhDdF5Qyxc
cWjUPILo5SRbM7D6kz4kCQEpHTQwpMR5vcUGxX9vAnp1XCyGDRcaRu5KPE5ak32d
uaIm+WXL9bIee1IGrYWDt0RcmOta9r4Blc/FdPlSmEhNryU7B6Z7H+D4XJLeEfEL
3t4lFxmFEEGfk62pnoUYkQPWwX++ZLzsqO0T9WrURV5HKkoOK20MVjcUNFLjRI0Y
PXJgooNI0MLbqH216VJ6acyBscuDcy8zWZMh36YmV6eVrOJlGNaar1qJ7VpClioJ
0ndUCg6/ia4wBMhQx/CEtWySY3uvN03L+unu4FOs+yFczReqpc+Frj8MkjO0UOB0
/KKt9gVJbe1msLrAb88sTHB8giTe7x6MiWsv/4Pa7iTqqgcy1ChkHdPvif/k0HgF
3hv4qyX62AIZ9yIDFV8+HKMU8XDYoLyDydj3HUZbdFoi4YeovEiekBOCbkQMMH83
s3zs7i2JWsbOebR4p50V9qG0pwknQgElTZ6ObQWsNhrANXdvEwFI1QiOUEGSgpHP
1k4GZ0T4a40/Pt7A1Y9o+RVn/dk7+Rv8ljgRG8fLJUuahxeSIwraugCXHax1GX+l
+KAnNNn1y0QCF5rUSfOuP0xXZ+xVdlTJpv+PtTw0E8xPeBxD8MebJz/csR1iOZ/0
1BmmZN5m377Xo0Pk12wbCPOAfcr3J/sVC/X6jtC8C7afSPWs9Kd77MGWLYBtk2q1
R8NG+0Ia/YwuTybVLP4iWY9bkVtlyAObn4ebhClwVoas+qw1nwpNhrsX9SOZRQ1t
MHL6WENId5vEv4ssd5TTdSWb5w9IdjWRr0az4Lc0IbXgTrB3TT8Zs3b50CgsIn61
+Wz/Qb3QhOXQOv0ymKrM20vY0ZI14b4x56tQ8BUpiaBar85IVS7z6EXZqbtyKT3L
qZE8miGL0zOWNxOBjWjdOG6DSG3HPIZYnXwgts/o6ZrYxokc2iz33sdprrNiY6X/
tzA8zVmwy0Wy6MYs/sqnSuVAVhK0Y8PKf2AKZiiI591mPR6vnSiJ90oA8Hd2FPWH
GaoxklKdoTZp4Mx+qnzLXTqdN7RmUW/eY1nhvgwPFeBBB8r7koN7FWLU+D/nrJEq
M1iqVcr/sgEvcgaRui9lGLx2yM99dfZjDwUDoMcCNTS4+XiG9hYq4dM3PNcDwsJ7
Mj6S9Kb8Q08CwQqFKXACmSrbD2jIR2Je78iCTUxjeVXIXQwvjAdCGW1JTPgIiGrT
Oeo6z2QlazCZ8sJVZTBUpsJ9viocy9NbtkmWo/Q0SjX0La8zH9Vb7oJlgHK1MV2F
XMFsSee+cBRtSFANYAwNIplNt5HH8AFsoXCInl69jMB1f5plA4pfIO2SKuPdJrtG
sBylx5cyHkhLVgC3dnmdHxOQQ5SegXLY9fqf5yvnrh++xKMcBrNzeh9LE1GMKNc1
UasSQhTFPJBlR9DsoJYCpnyL1Mdxr/mZIIXzKC1niZek0j2mbvqLeGOb4p3Coyo+
Fx3mKWEwuM1BzZpOFH1JlF00RebaTWBnfaCzeKwWSrCtMfSpFrUhHgOaEzM/vl7G
oaozFWCoSePmWzKPijzcZnRTgfcmzDf7NOji86sc8pbPFo+FBXRb6ZU6EY1AdYTJ
I1648Wy3zLLbpNH6417pPW9cQfkiTrUSLX3EYkkkJk9k5GGGfCnfavifXalIcJGH
GPh+w0c+YKU7FqY5FeBZl8+sFC05fBpa4GE461byaGq4mzhr0dQLJu6GH8JGyimS
cPIW7fs8WVc2o5TqG6ZuP7RunrDPhj7m1CGZtNxHxk+neUqjgJbTFpwmBWSKVPsw
Hh3rW0Z5/oB3JlDOQ7l7FzSZrjEnHfqeMdJc/6kXyxUtlfVSv0J00WR0+Bc/ukJe
oMPvTdrKNYbQvIlo2NHM7CBxBas2dLn/AcZmULcPLQjsW8ct7EOAoz5obpzNAWHz
T0yxYdnKfBjyEK321WS83746Z6rh122525WB9l/DfF4diRLp/PFHEwUZm8BP1gCM
JkPBvEra93VEN/stItadSD4g1B6wZgUCchabRz2rk04XHd7ZydPjSWgU4QCeK9E8
qmvv72Z5VOZUnWcJbVKSBLpNEpXXiXoMSYFAdh0PnzcYeXkuMOUwCHU64f7UPvwl
hV/eqDSyZVJB5lNKrfZEgmgJRMD6VEFYb0Brr05nNelPGWrHXcVf+lHb/qevbySS
0Cu3pfgp24sYAS77Qe/+4dHbT3Kkeu9L8p/8a8EI0/Rym/URE4T+ag7vMph/lcB7
NBKt9jZjF7ZfP8ZXeBiCQyDaMlHi0RKVsRLK5mfS/vJjo8XzO6ROvP4PTXW+acis
8Wk3sxGTD9eXexLUMNE1S3tzbCSHlHvlTkYuedB2hUcDCXegaG4XaP63hxOgfTYY
OQAToCxbvneWE1rIENk+TB8wjGmQ0A3ETBZMq69BrWTIXBbmEOf+KaSLaWMjz2Iq
2+Zhd+we7uW7h6PaEbflCizCXGSZjD4tLMJ2BL31biKHh7F1WQkWIjyh175ktrP7
90LYTvtTb/4Tc+qbV3iGUyw6Bo9DbFcYJ8uomfYj8emhmGVq6Sw+NFqfoow58Aro
qbztsGT6JjLbuzuHSwN83d/ab/oer3CZVT1SWiqSRl2pKyfHFtl+yydYuwyntYMP
W6HID5zH+5thOFkoTVMMoyr6MBwuKRJxdvbVjlcg5dscO/46fLYaY78OfRVIzvl8
jWm7VP3CEB8HVZ4nAq5wxGHVJ94AS6RwpDOOKVlbNYq6NaJJDJdxWMkGzHaZWp9r
q/l3VdW4BXG0MgVEynh3grGLPPaVS1Q1dfk4MNOzWIB898DfVNwViqZTkTENyHrp
DU/+Yu4vViGH2hXGwzp5ujybnQjUlSxkzhHvGzBTTlAXUJElcxXzEe4Hx+Sr4Qz/
HvCS7WUSbcQN3/e57n9HXjdEgxuQ9j2Onj40GauAg8IKQRqMYyPeM6F0Hn0M8q2+
tLdVxH4a1wy10u9cEtSah0uSJzqhRCzvhUmxGgeKqK5o6myHAb7cMn+msej6gIrp
XZBvTIp7An9JnhCU+ZNO5Lq8teavj+amKVklZNHvpUFSBDPLU28N1mkZOnSElqKm
hOzAiO/5J+7aD/S2MODeQTTv64oxZJsSHsbxyRpbKa9cRABGDo1mqF/gKt8UNJxP
giv8W/DvFBCuTtCeLNM5HW4oOlnFGd7GhS6qrJYaV4cv59dIC02jro0M6XPL41bJ
yfhenBRifPDuMcErau4m3N8Bw4TWVNMaBji+3N+0wu8syTadoDiNFJHfFUVY3qtB
05fzsLPtwL1XNDqdg1McdHowZCFSQoGbG8sPiEpROmTG1UlGRcjvpROXiW1Ek7PV
Ae+TR8Fdt/RG8h/Ui16Fc1fZPV8HqbQNFndC4QXE+QbV0fT5XQF+MSwrJfADYRUi
IVocTQyR2eMPuQeXoh9QUyJcN7PoRNlvGINtw+PicW5hhhp7/+VE0B+sLVtX8JDn
iHzMVJtlDkvO0v3GZwhdcw==
`pragma protect end_protected
