// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DQQQfzAshhwGOC/+nBoXhPppv0ElBQtIi1TBl7O4WQ8MFR9c6SORmmsbW8PxO2BT
QQoMxq2QWJQJgTn26kOARWD9drY/D8MXYIeBUEC5VR7F2vBC4xscKco9bqf5GBvb
DjkBXvFU81EBXEECej8L4nyI8HbC+hUPe9ehhgswk4Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3104)
9rCeUrPg3h7Ruqv5mKzVEYTA+iejIM8PDq6LEjYFpPU/NiRcSvqNsqUBJbJbLew4
zS71e4Ul8ZXQoc2L7ZWyHDzqSFyKQJRAGmELy5BHeFTZwytNZ2OClli5RmrMFTui
lDRG1MveBmW7m7bnu8+iwIIwIU7CsI+iGnhuwlRTdwVrhdmY9qwXGlrecj6PFXN+
FGHJCUoE43srN/kuPrchwFYOFWzO6W0jnXlRBvwGmJsRwJ5GNe/m+avYp9/3ZkgL
oeHNKamisf7EkjmA5Jau8CTahPzJQRAvm9VvKTUaCwo3EBmUYaTu8iVkHSdIKW4Q
3QUUZHLqpwnbV2an4BDVf67ppOfO8KyN+sNj8FnIsWFUC3swgyFfRYR4ooGETtkK
2vrKZWR/DItdMamm3Gu6cpiFYcXU5gawsPUPvPbjyX2rVxI12wimAKQn/TnKtRUv
nkuBm8EI3Tz2YmynHAapqXH5/ykFaR3+HBbDt4gkIsS+9mpvj7i8N0I0H4yIzhew
Ae7LwlwzkFr0L4oJyulKlHZMFLWQPp5JsS3+Vs1qHczuibKB+jlULHyhKfe7AL4r
qibKK8PcRZ4w1ujzPLkIW++65HMlgou360dMJxk3ESDOdqEhpA9dyYet/ZsvtZA3
Dbpw/ibSoxxxHdOf5/cJbm4swiQAjv42YBKa3diViGNqtmn0kjjJzbDLsAj9Qlnj
fn+W1Id0gKUFZaSRnPqkGUxEFB6cpkTxSb6Ycrtjg/I+i8AxT3LPR3WlqFDflsIo
1sJVh3LySAbooQ/DFE4bczEvHzDnAmjWoGgzoOrspR2RpmvvX4yn9fXRbg+n2/HZ
q/NzmfWxSR6us3IVKWrU1CkCwLocTVMBRiqDjYujCktioG1dzkFdpfQFVL4B3Z4A
v2HShruYkvKlu1No2NoclwTxB3ImAQDc9KB6X1d0DO/SGATW3Pc2kfLo1KRknHUN
S8JyLqU5YlF7A6NnYZI9KAa0D2BNSV+OZjW11JXft9JVNRp1Gj9kh1ngYCKYyuvR
ZmcXa5ur/zioO0goKZMvUpuby+XvBevLQTQEI8r+FY7fFyz9C5zCttTNOpCULBgX
BX4K8Bm110upF4AP7b+wkYDeUyjgX6/apNjIC+joqSy4kV8rnVWhOHvWD5Noh64y
zwvH7qSHsp1hSRKA7VijR3xQaNHFipN53yfDYc0xSZx891iVece+LcjrsMGhhct6
o75HjF9lyC7lpIfKGTBIiwj/lMemld1s2Q4QPwnwbbrmq7iPba7dG3gxewvvvcOb
sKStu33kyiRsOzGi1C79K+xS5ejOFTq0YK++JhCmYSjDxwJxiYpVAriGtgtdzD4A
G4g9asrqqG59pmQKg8ltf9Ch8X1h05+chGFfG2fi77kOgCqWfBYEkzzNBfQS2zsf
e1Ub8BBYfpBGHorhF44CM3/T+pJEfGUV766RcyJZB4pnfgoKSVumnNXlkaUaQued
MwL5Kzwcized9Zqn+ZnlT6XlNEfHvwNxnmtT3LeGWorflcuqDLzGRpNsQGKgz+sO
SNGZse0iiWAqxNIPSxP7Kqy8gRn93Bgq3lr/jVQJnwvdGduTdeC8tbBPRhWA4Dbb
rPrBX0TKTOYTU8CsV+n1sjfG2zU6C6ZBYERy379Zn2wq4hImhDlnY+yh+gWHjvGP
4ASa9PwRbduali8/nsuZWHZlTBvXVGr0xSktSmjyF1uwOsGT6HO3EEhRqxIjLOQv
5bKQrAqCBSD0ck7OwkMXCc5I5LgtJkrSihnIz92lmMv7RUCbRjilojWwYNz7YHp7
TLuhqiHhwjGLXkIjO7lpi/x8A9UvwDIzxbEWZnxF4pC1vkVFKYO/r1wOK4BYO4DP
pkgbDZjNCb1Uj0iL9SiJFmk/hwJOdpIwxCabwd9c9W8i3yL1a8czScjILJZC9yTS
9ZO58AuzxTRkM3Ui/vwkJHKVEsab9mW2fwWTGF6NW8ViGDmxf9FfT3D/cYLR5vid
guRn7HFhI+8+++WCFZpLYMXyFCLM/e5mNOsStIOJ00zs4h81QJH5FzC2Iw/aeP1O
dPgW1GCQPPKDSoyGf6QWaUPnVFshLd2mkzdL3fIfI84liybTEEAqZGEAlMDIZlgq
rcdXJowu1IMYvakpqbu0G3JbEYuFvcmTSn7cy7ZZeZiPOR/6srUG+l2JGQH4OAAG
ewNXs1RXwUGa78U03xJHmOnGoYFw/DsEJg4Hh2tg4cK3uuu7ffqQhFxH2vpy7BxA
5bu2yZSafgx5RWbfDbRrKdY3g3phrm6N5RlABqIMiPk4MV3N36ReHOmVRDBf0674
aD5+7pIxkgadkqSTP+ggegc5BPQaTl67aFJ1HaTi3duWnu7lENivNmuCiAh/g9i0
iOXsqAchZXl+/XqexSTCnnyN7aa9D46qtuBzL6Akd3qUyWGS0fQOM8aEBXP+xQQv
k2WE6fT8AtWqGeFGsmK5FDDQpyFHkeSlZMtDIcYJPEgDaRbEtfnhXxS4JroZwNF9
b4o5rAO1MwHMy7JMUw3JuNTgUYmYrFJ0clMg/5bR6vL+LtovJTZJ2khhjLvfiZFY
Y04x+IYd6vxK/AJFpyxlsaSgwhztivCW8IXACdI7nbyU05LQ3xJerRnmAoIKQrP9
pp45nemxldo0FH3xp2JF120xhs5lSiB52I8XedP00aJn96x4cl3eADYkJefZ2xpn
LyBG3w4xXOQQjUEeJQe3fCN2vTcb3ilU6ZgY8sDo38yNel5eaMLG/pmo7HzSHcUV
mOxGIqndoACndELi86wBtyktiEtiZtvC8SPOxVI/wdC2xe46c5shVmOf4NpaS3W8
goiq5j/qrllaAJGViyfEOWp190S6qT4cczTFm3du/hzgWCh7tUtjP1XCI6oJqwVc
2e3DV4FhkF9W0f+Rf+7UzHciUY3NgN/zUihkCuP0gm/gECO5CRjYGt/mUVnk3EVQ
t3tUFYFKJEE/jOzGBQNJnkU52ydG44Y66I8lkcP2HMMwkk0Phj9Kr2gDwgBAka7T
W/foqe8y9uLo4wFl/BRPEyB1qLhHM0jynubi9xtlR/cryNSceoZqEC1eSFjP6wqH
zVQQNCbCLqVxEwDInrh54XLLIsvE3cLWYlXStk0ggd98WBCq6qvAp6cBVnc6nzlH
Y3V00MMRNSQJJG0o1BqGQ0u2nhNcq2289yCy7TNIGAm4G+rXIl+h894KaREbHkJ7
s+7dhT/6jfSoyG/hdkbIH552bT/tKprQmscJ9XWyQCBVX/JrE3wUxsAVelsOUBfZ
JNmn8oPcLOZG9y+IfFAZKagjiaYJhh6phnlMUBTIumoTvqWM3vmiTHOUe+IiB76R
J/jZ6jq6ERoHrhrqKYNhjeXxFQI+HZEW+01N7W0oYPtnGfCEWYebV8kwNxp8h12M
cPFNRNnkhSMLAtNirnZSIk6+3/7XlYiveNJtL6tuL5q1kDd46sWbFpl+BDnXVOzr
LR2ME4o0EFkb9WnYPlUZkMwgJ2Wopwf5x4EVL5m/lGtS6IkQwEsbL5ozg5Cu+YHC
Z1p65jercEpeC0+s1Cyu2loRl2IBe1IyNxw6Y2ar3eP4v2b8FFZbGay+zVvb+XdF
QHoxmBi3t4Or75vN/8ii9S9CHhDRI4qdU44OxQHBr+FKJkh6+xsRtUHk1Jue80gr
B8dr7JVOi44mms2WIovFDHzTOIJFRt7Gawv34d6R1S1/M8M+MnUaFxAhLNPiYGN/
xYadNXUiUAUWMjVFtNSB/iU3nFsWGRXx22uPUUGKDQyDZasrJt1B6F2LZL9Yhxkq
w2ETqTxBSyI9B9g9SpAdGi2CvJtS9rhc96XZsFokmJV/+z1Bg/nsomGdCiwQUaCj
s8IULlAubDGxRJrQuU2Rk08hVtc2xQ8Wg2GrxJVC/K/x3jOYYiYkQ3ZET9Qgz1Y+
cz3otA2lH1vCtHflGg3iM7A0o56dA8zX8Q4rbdGAMvKiz/S6ilYmu5xXyaw0FM0P
JsCezYdLIsv6RdhNZBzhEzoIhR9fHailgA34CiP+XOLv+z8t3BeHj5gmgCRaWz9H
yN9pIXXpZB88QJR2qb9SHl08nyiMq42xEiV1trtAZW6yQF7E3PO+ZFxMML+e0OEA
lMFoUtjgI8uyiM1HYpH9751+Y5DJ4M0tDLtazMfh/kI=
`pragma protect end_protected
