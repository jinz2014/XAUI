// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GBwNdZtmr0p1/B0DSujsOFoJsS7QJ/8cy2H3FWWxVGJ8fM9L9Q3CPD9V/zUrhPkl
bT/UFYJ7i1oHFd/X5TEHUyMQe3dT4cwbkCj3pnrjTNfxp2jUNUd2w70lCJKO32gJ
GMBY1OqtPbZ4JbO6FO9s2BqX1VtoUx2ivbhgw3OkNg4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4240)
vxY+0ejAIMLHNDNMpcYK+hCFDa0LMPuA+gTJCnMiRE7qAV9l5moh6l0OrNPpuSRl
JShOUdHOohGoBHiGoaGcx8KQydzUmQMjqpB065j4TwV+NbkyR4Ro5kue7FGpNxt+
ExRgRLQ/aoOdgyj1nHilGHPHtBy+bFa844qvW0zHCg0hjBf3pJu4EkwRXrQ1N23g
18VtlvmuJWxoYUBph2YhjTyVb/w0GRK6I/izmxSlkrHzvjF7K8YTGdjoHMQf3a3i
OEvQkweOLTehneVcIsc+A3A+xXs9SUwqFRJIWVOoZMUX2b683vQk+xz9SV1c4ZxN
OHRtQtjTz+1fLdl1JSane+neuKjoMtJMfY7j4xvpSudVqZS1025OXdqlhzIQ2REG
qQ/gh3GZf99q3FoimIYLh0kbt5FOXv26O0wi5AZr1/2IhXK2F0yU7iIt03f6BCch
YefBL8CvIfrhR/eNJ69QEOaz100XG0erRKikI6EaogIKGpj0WOfKtH4C8/CKRyrh
XfS99KsyirhnJBnFx16KX3rF+M755s4Px+ogSNNChK3m44OvzI3eDT6333uESV0z
bmruNFsjFD7S+yM28EHQ2JtB1xMln3lBOkYXLZLcDHTAJBLpQCZcp+pNNRF+7PZ2
TQZg28sWIJKhQ0T7wHkCb9SooNgONiuW+jhG064BKtGkUGHtXEtaRrO6codq2VRW
mqIZPZmQkC6PeZrEHj/TENfm1BUSFHKsQ+u7+/erpI/OoK5ZmBrrYUJAXyFaRCav
ROEe/462Wti3c+aShdjz0mjyXtD1CR0qBa1XnKNUKA14YaN+sULMwIZyhXl3hGI9
mACFBQYTdVRFOGLqkgcUtkw7AKny/a5gJo0MMwg1Ysy8rAaOXPeDzr3yqJo13eCs
rjCEV8qbzqDAbGIbwKpvJUQkXNlgQoD3RcSqvIe2PSDejHSxjoemiucJXx7LdjLh
KdaiSOUlw33RQ19Z9JgrR+nF3w2epF94AahvrvlSn8XYz6euM7XNHIRIYJcfKSi9
iz9xL2a/67N7FtbpuskpOe6+kbHihbm6YDmknQ1vy4rA86S2hknnYBOTgSs42CAp
s6C0k/cpdZfIrYkc+EPbvFncrppt9TTKbRF2ewxgA8/mBsCWxRY1tbIkzUxM2/QG
uAh8AlHl7v5O9GnLMyG3De4285ymmuvDgW2f6d+rB5rLBzz7vqzKJBw+CCRKJvOn
RhDeeOSVb3NcMLl4ujIzaxdox+TIdnaYBwDkzbcLQijY0utysJYRkTcKnlboGp+r
JSWuz4yWLb4Yi35/TvV7DowC6Tvt9iamyF2lVc71jgMz5cQivB5eLIjzcIcVu0Xn
f7QLekddHwAnRRJq7wr0s/Oa05ujw9piReUg8nIYGhGUxKE0y2GRn280VD2ofeUL
if1TEdRv79RUB2dzPkfyWHuMvxzYa6P5VJZEoX+24hdVQYCLajvzWpiP0Qk0i6Tv
JnI2ogfRiBHswN2cBrK+SEDHRq9kcYVSO1omst/OlAwprxG7Zxz00iVIu/ugrb7s
aty+dxzp2c6Cc5qHszC2SBkjG+EiTVQQmWIE0czAS3GSAVIWLfRjvpGIhEwsb9Q4
T3wJQKCpCfAwYDKitkTEIy81nHVgMjLG4Zq253ZZbVyaecCrEvTWbGSbQvGu2Uwe
0uBLeuPy3npJFbGJ13/5iYvrfTiQ2bPNEWb1hBSOps/kO8fV8Y74t5LBOazQ4wk0
I/Zs9Se4jjuoZMUzx78mxPiLkLQvhQwpZbG8CcrgLQj06InwsGnSz7s4dOZBph7i
sofagsIvpJ08WT4TTbq36zXfgEYLRjK2S4kYbrzUzDhspssdh7IJjYnvh8ENwHEg
Se9KtvEkpo+hbf6Xwk8pqipThcpyC2Shox+tTI95A6KOyrZB6dRs6YeoDLjdlAM7
etanBl6o0M885s2NIZr5D34EJR4wVibG0Y8dVP6H2Uw/RoAc9RnPtMxlfrU6PYJW
YEuo4SyhUoNvoz/a/09T1De3qp5/CJ7A8aEAL/Ry9rXs6Epo4nE3g762LvU++v7N
c5iTtarfD1AhQdRsiGa1JkH0qcDd72limHVODFPoD0dIRfcO55SXHumKlQR25dnL
jRs9Tpw7UILnfnEWDkd8flfjCpYWaVc9RBs11RO0aJUlQGoTAtj+J8i1bpUvEJ0b
a27tlVqr9c6b1IBzQSQ0RKi1NYSFYQyMcMe3CEpZ0Cs87Hsq6kxNZJnDs71Gt9SI
cnja4bNvTEAvWw9C+vL//Ms9NPBvIorSOD+HdPMJruucJXxrG9UXTjgjl0uo8SA2
bqzkp69SL7AjFD6esAJ7BBM57fCfZN2zwWHuzUkDx97i4nHvkDBzPTy3Q7buarNx
b7xsYN2An30HDsP3IzazK0kxdv9ltjiqu6UHUqlRaERl/oc7Oj9ZwLXHpj4deBTX
MJplQqV1QKDfLemkXwemJTg+RfGdupBYWMd/v8dj79ADQc215/xBkxCyFGi0kNDo
tylcTexXxb3ta95lqva/S/E4ahKAym6pT9kkx8eU6lceiwpWg/gOF+rBaTqN1KJR
9rjSpJh6zlNc7bjNbSLfAVO5DVhNSpZY/TAX1apMsw/YQz4pBcywS4WGih+EXbWU
JmGGhtAJWrK+CSpYFeTrvIec9X0oOIiDqE7i1qgNJmUACA9QgmO2hYm7pnCfy1pr
LIzi6GkBjHbBUbzu/7Qj/V39Vwws4+YtcuG4fovmq0YQ9LmCYlpS6UrRocS9AHv/
QN1zU/u438nJvM4WBqi2RATMSD5wAvSiONgAZri47nPW1OgaT9xY6k6qu89Vkfys
y8u0xiLTNUS2qOrd06eQVF88x+QVRB831Y9cwq3YAyCEDO5UlV7XMDWPU6lV7Xwl
+Sjm1P5w1N758uinzyl+Juvx256F0nu4O4HL4R9HO/yELrnD74J4xJg/RiwW7oUq
oDEq2wCewCPY5q36AfjtTcXBWJ/H4K8mPhqRTba5ZdgLvJjayEiG9mnL1sxtE/C2
D4olnXewuSZit7ACEbnMYL/Ywc4Ud4U7Z/0/ZYbxQBRK7/WnLqRwc7VVdxWKjvSZ
iB32avA21xCXUwsxE5qeRxR7hmQPFta1ESXEwwuYzgEDhsgVU212VFy6RM9b1ioj
ulkz1qISdMkwVnqXxVQwDtDWhn/6cAwFjon9L5oYCrAIzRzDgg7hS/WlrE9fqbQ5
c5LjesJ8UWWLM/SmrwVALoVtuCV6wTONAbCORoyoIKalbNxs+hBn7L+Zs4WGzU3g
bQlFTbM+WY5SkpMw/Vn8bZa+W4w25DcbsP1rhpdUgAc4fMraJ8H41Wi3KbO9aM41
oS08nW/I4J+Bf9R7xpzi8VsHgGrcIwOD8sCEH2PGOIQjj0c7ENcXmj5wLRzG/Yjg
rWZcRe3MwdEY22zH4PzvJY8QY0QYuB+PwXnwVfWltjgcH/SZjh2XV2bqKKLeJB+1
fi2HDVZBg1UD622uEp/qWMZWpPN4nUi4dsjqXwi/Tc7VIxAc9sS2JG7bBf+ki/kN
EFMgRnROfJxqN5+xhcw76o67v/6RRMZ9eT8AzMlbGpxfDFYciNcf+F5nNcHEslD5
lcfiKtYDnSYZd/a+eAEsNbaXv00+TZtvdUo8uE3VRHZgbEPHIKcrBsPC08OIvFPj
XlpNgqvVew3pL37JyJZzSdPoDr2TD9eZcXTM5A8XxrOwosddgNf8TAFKfkgQv6MG
eOqRwc2u92jYgpMe0WecBbURcPv+PCdDasUvTR1EMaVvXvVqfq8MHxC2y3c5Kc3V
7gJkZX2aD/vFMhGdgiekf229DkdGG3E/uLwa0HCR/SYMx0nQviI9szXnGRY8/wXC
i8q1eTfP1ECAN6xmfHYK25BbWttekrGSEKIppktPkl+7w7XSOYLlcroys0InPv+f
MJf9PXtmpYbJByBDu/uUMdjqTp177O47lBlaxgi9lkmSBCKRGdlTWgyM3MJR1jZ/
9koTSX8E4yDw27ZvY96xluLs8cwosQP/5tiUwoOkBQvxYFNoGnKxDqbWLoeW0iro
adgfCEJggvA/nSoRDnog8xNtlASOKAYygmGVjk2A6D+7I+E2bovau9jhA95kVdS/
VsdE+sL0hBEEIC4UrXmUnjxAAD1ea4xLpsfny7KtVuRuQFLk+OVw5rdZIo6w53Q/
W0VEKD06x6A+m7CJaOsTFRGmuXq1zEWaNBw+Pg7vF/MAH6MUOE1z8FVGPSkVUDD9
93kbBDsKr4Rq0SIi1C+9VjKI+fyp55MQPsvcbQBsvXfwKF8maZQdIxBq/7AyPrXl
fBSiEg8Cqn4/L+ta0gv4TVzoaPX6noqBbH7gLXo2eWkDafl1pfMD+tmCem3JRPG3
+D1f60B24A5bcSEO3UQUzePdVjHRc2A59fooil8g6waj+1nJZLZnchYeCaBhDLYG
uCkgxLEhCowFPxYqAFxsmGBDEHdDNS8aYCxqKja17Qs7vnQD/xFn1LQnHJKCCO1R
8guC+DlTHkINiQBNFtskA8bSElhnj8fv2Nw+aEydpATz2iIos6fI++PgEz6TSvZq
GAj8pUuAGGnbZA/UUZZYKLilDuefHHuBWi/k0AgrhI3Hm3czM6ddWn/OZmpV+Unn
pUwpbF+NizOE9+2aswrtxnfagZ/uh6fSXAHbfRgaLziDnuh7dj+uw1sh/g5jhcGA
edW4kR2KCAFyiU+l6wYxc7BvXWV0TIXkC6W9cxMIOhHrIzgwAIyJ0GGrSHjSWApV
3Temk3wDnVXxymOnSnvdZiHHduTsRyiW/3S0CaGjD6wHYSxi6MlGwV9+Nz1idN8r
lFgUDseGdQXgkjFrag3Uxuinfoukm0KK5mO30DPxd+DpUX+AL5nCPi7CW8Jms4ds
1ffMdaMtu7W6HpxWfe7elGM2BqErB2kNbphgyrg9CpLykuj7f7Caot9vmcFfAgcA
XZEdE+sNGzDQqVyv0wLDyzPvgT+pK+7tIK/KVE15yLZoEYwT8ptVerCjU/4pDFSY
WQz0NA1D6qDTUzbRFGioB5FQRbOnEBG1QEnl2TYMVcYcKBKe8P8MBDyOUhg+5HhZ
cMQsxsd2hxPgPtANtmYGiLv24qcxTjHQQkWJHYLgFo3vc4+YIyT8k2Sd4Vafwd1a
W29Gq/7ngBVY7MQTFoiDvMwfvN60xzDHgCBqYLiH+p4idt6xM+qVsowOzOMp/BFP
TZxLRHMOss8DUmziaOedBWiT01Lvl7PPh0WW5ZS6EuNbDaEL6bQreYpTSwuAq70k
9nb2rwC58DyFOd31tb0WSy4/GYYAw1U8RugJNMOt9YB7uHO+sEeZDmEyhnGEwO41
7a2pIg8VWxcKTIvnpEjNs5c05RuLkDNW2VGu30FlwgMIktFpddQ9epfuvtAtic5S
Ol12rVv7DoHSMtwJQ3BMEeeoNXUxsV3bgzmOUVMw7nuY3zbTFFCAshBkvADmXcMu
HaHgSR1OJDXVpUc0GEX70ZAhxhd4CBYX4VJqYbo6wGnqxoS+esO3ZD3XZFH6sEfQ
fje5Ji3lS2J2le+Vq4rZ7Kaf2uMjNGNDxiETPJpjtjN4/wMgOjl0Qe+Qsey3QZM4
EMUfvR6ctXdlkH/dZIE/2Xim5gRNsQdMOTFEv0esog3fCjLkwXnMx1L+m1Kmn4T3
KPqCGPMtrSjvDASS+S1bww==
`pragma protect end_protected
