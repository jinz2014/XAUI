// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NT+1fFLt2IGwmq0Yb0yyCry3MmV6PT0Cii3r6jHvZYLAvzaA6FsZtSAFPLLqHDkQ
pK1ojl/IDZlIT5yPCUQwfiR82EErsUJ1XTmKrZoRW3ssQsXAISXolovN9MItc8FW
NVPhCSewDjVV4Nnw2Eqy3MehFCKAKjxH5DGlh7XQUAs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10128)
oOyz7XcJCNRw2rT6wju91MaKS5G8fuqSrKdbeIlgn5r9kYYe0ITbh/Kx+GtvEgEd
A8+O0fHZG6nRsCM0ugCkgKHe/uO2kB8MjOm5wjtvwS0af1TaW2zkpOgsFkVoQpsm
TqdGu+dLcVuCI/iEGcjeUN6C1oylUectEegABQiMGJkg0lvpqk5HQ91kyAiHiufM
99zpbgw+eL6JhrldXn3vyfKtndZJdEPbNvEfiazYQK2B3Dyr2Hi6dc+cP02jk/qo
j7HPJxJpd8i6YkuezSgO5j3b99izuoJkveJ/zCvTtM/Tw7GrskSAaQ9wK1kvcKm9
aPulgeYZLq9lqH9oUOX8wpMtvCQD1vGL0kf4N92QhEi+Rmb/BB7EfNif4QHKcqph
hNHDxfuNAdFPR3RcBZuekb1VT1inm0LiIIj/YgIo7cmoWRtWj0clusl91R60lWzc
T7NRqBrn9qK3CWuKmONTltJCHABLO0fBQNG7U/MY2WYpCBZGzta6IunvXlMrPWrN
8Onlzi4i53gJCcDp9dYSpEgEPwBkT/QRABEMbrWGuN+RrGeNdaY3QHLBcGpRgRWY
IZTy+8c2hpnO3db/VPDnQIJo3rhbw9h9Zo4c9Ni9yhymhRhOAmOrGec6JMnEwreW
bS4zNdT9MkpP0R239e02G7SSEX5gj4/Ts6sbUjDVfg0w5mDNITeWXdZMI2YowDIX
S1OmK+iNx7a9knjQkpJtxbwUsZwsT7gQtvlvbZKwFIg761qGwYK9saKEInURZCbf
jnY8a/Cm2ZoXNTCCysD4z/nCdM67eHQhVsFn/HgVGyu4rqTCBw0KdoErtZGlOhrS
rUYvF3j9UD9mJVZiLeq9dACjWYDJR5BtEGaNV5Ufy1mG8Ar40+9EZPlBEfk4VGop
v19DCp2IMmfIwsdGJrS+4ffFCcD2L9Zm0bbZFucLU1FoxEF4Lp3adqK3dvHUzGNb
hdwn0FQ3DCDQP0Rd6cClGcx/PRPdLG81Vl6lVi8YjD/BmAmkXpKPgAJ9qw3ONa68
tOalebefrZ7MJtLoNA0M4ZOsb14j7hjwe/SjLEidaYTj9diEELZ1MrCXCA5axR5S
m4TFo96C9raus3qqxblFAUZLXJ89xdhAq93jOo9I3DqNDfF3cBCGm3dZOe8DQ3tu
6lpEZnvh7T4qQNH6XS9JvU8lm6naRzMT9YtiElkte5nOcrnhaJXB2wbikDAuWCQ0
xnzmxy0yvjzaTx1naotByjYV9oIymv/xXGHS62/ce5/CPFPSiyyai6EuniqZ1cnB
U4ZxjAu2vFmlSimkL8TuhqIhGDk4z0sPHjf5NPZNtFnHTHHHpPH/mIrvNwi1HhDT
mIXRdLr2q7/3NC6bH8+zih9Rwo8QUt/ynOFutuCsRZwcjiuvZmKXmPFOVUxsIPnf
ZQ6AIJVTVeqeCkz0w0i+Dd+PKMlo68Lw5p4e46d02vGkyPf5S5mbcJsyaz0BGgZL
5s1UsV+foNWHeyHsZrlDfm1TM9cY1EVz+J6khLCgt3ZNER+BLzgXftrsB4LRJ9eE
z+nrp/b1LCByjLAHZ7mGDgnf6X+Sf5OqJi5seWZxyfjQ7yUpsh7Jt00SB0CLJ7RR
Ka0OYgRPtn3fj5bZ3YhDmlL9hLwlK9VSPbnm1PSJS61yi8UaDa4ZKKByDNPAL5DY
mD8Q8HHEZVUqv/epb/7NmRpj5Ov2iFceLzAMd+X7RK7HhujVMz6oovf2g7t06SP5
WUvR1bUAKEXODfBwreUac/oI2eSW0NFyzV46FhqnT3axtLfNTS9WeS6pRosnLMCB
RONkU2AAQpbUzPcOd0YCL1KS34dec4SHFQlHG3yTHr4fnOZALElvf+G0s5mlG214
NTY4xfZLJvgvPpWcngKgFwJTEkTfvRGhepIE+fi1va27OHY7YqyKhQL05NK4snkv
Hdc4wALsR0KjIfLSrhFSIipz0R4TkyeAS7zi1uV6f9ECegQqXodEx0qfSEzHmzbX
rqxPguIO3TPKDVjZnY7ldlN8mOw3UgpLWevUEkMrGCW0hJmRZdBfRQ2U3Qzk4XJp
XrZVK1Vebjgso08/C5Av3HG3Eza8kiZX2HYefUkRb4Jy3MniFNGxNhI9Y6RsqCJU
ukssR0smhlXm10LH5gxzFEdLB/2vR5PIiqZhKJymYga30EhSGe8sXDlamqkAdzIl
H+ULxXXX8klTQTKZg1nWcEc6U+fJLnyqjJesnbKjOKpf1O0KSclH4zioSlegK6A8
2U/fo6EzYniJ6YKnxK0TM2barckHnajlERCQFOjUiNStV0pKt9hFH6C/n9Z3cNyt
zvUZ4SgWfPFA93d1hSZgidN/g6WFRqSTVngznohb8ln0EXTcrZUWMo776DJR91T/
pt+oFA/o9Dldows6hNs3lV8S+m6Ul+S/Lnhyo5Gkmdt0JV9NUsaIpxLayPsHla/g
L1/tPdKC5jzZd0bhw0jowAT9QxUQEl14ixcTY6P2PfibhV59R2SrT6jBcyNMM93+
NjLsioVqbQy5Ow181kTTn4QFCjJrZEK9MY5kU6vYoCdsdXO5vk4Yn8p7xKAOmqkl
dKI/JUETsFULWBVkKP6R5DXYOs0IhbB6qwOZLxhIahvpKSLFVqruutt2kyYmUL1L
dcx89C+PlAHTDTeRJH+9aBXHsvQ7tgYIohKpeiefLOdOAPOGCKaqWqRL1lGj3Ur7
13JMHxY5dTQyOjFdFUWGpcuilKqXEhIe9s4Frt9dfpQozxo2HYrbLukAilPxhYKa
KaJ2yJuZQNXCkdh7WpP0Jei+Zmf6/HGg9kvzyVbMBDd3oWRc/rwQxDUHxPPjhUv7
HA3MxKvW4TtJKdbpogsocYlC/lr2+yHo5lG1Bq6STU5grE3wGzWEpfgPo0/2IO85
EGVgDEXC3dbe/4UvkvabXINv+/largAd1tFXmcERamzIEUc8EVCnm08ko354TobI
sN0DfDHCVkF1oGyBIePw5sZyfX2OwWQkf5IfMX6T5IaLoMST36LfTTsU7qX/DRby
Jj+jrB2iiHY02uYLe52+ZY2u7s1UB+UzCmi3BGDOD00Y2YQoj206juSwWw1Xm1SQ
+ahXSLQmtx25OTfZGymupLQHBtG/bcKsQAHmpZxWv2wsr4P9pB5+tKQUrzLvALgd
Ct+4x5nqshLFL/8dll6oyLN0RLm2gVMmyEjl9Wb/veoF/GVhtbsP+Ez1mkyle2Qx
/kJNR4UgqHLMX4UmJxQpaIv62pXxS4smLmJ3gpFjHDcFsw/1CUjbTf/yXAgWp6H/
WoE/aqMvUvl9bi+ID8p7m4RkZkF/ocethBDcGo3jA4o9zWsQvsFCfS0BxZdpugVj
WwERXCuRPDcf4ONq0N/YpJJx1CbLCS3crgpXMA/iAy0mYdgTVVBbkIMwA15etWbf
v2aZHSz+HnoSpw5dyLGRQo2lzxZjB1XiDv4gao2Frsiw1BGoPWAB2PDsfmXUZ3NQ
xEC65n2nXsQ0hXyDVL4NvmhbIHNHupM4sOy9pSYFsihMKSrCufwJHn9IDRiyGaOB
kZtb2vRE/rZW+SK/FW89b0nJZP2jx/QMarGxrHVkVNwOtjkLwI56hk85Mpm6IGZL
dmToLKD5jgNjlO2rG6BsCh8DHBJUPj0TXTDa4OZDx9CKaDuvy0n6GpwituSXlVkV
lwBSNJzioC8115t6HTMhaKRPxW4vR7/KGIpRxmPQ4Hx/LTDIfu7OyDd2I2kPuIOp
rKd8XiNypwFdLWV0AmUX4c5KLfqB6POZI21tGTiXy8z2iDCFOWEfYUuOIv/UH8B1
JHSzeqKWtU+lkR4ClTzC2C5jS5GBrgt44lpd3VaILBqFrbe8vi7CiT7mg90mpKvB
SSKEAhUk7EMWGNtn9mrGMncFaFxqH5jHowU83KS5MfbusfDcGhZKwrTCaDeCr43M
hjWr1x5+UXUCe3TLIx8lIJ2EwNPs7L6ewaD+Wom0qgFkjRaSo1MOYtrQdmVIYbqf
XlQzw1eq9BlYt3VYBtqO7U3RODuLlRG+x5s8Xd8x1zULcp//FpimLVu6s6U9IOb2
TDNAe4VYonOk5jlt1emYhkid126VEtI/va7X8D/j6Ob3+4RxS4QhZv/fAnpwE4dX
AyOck2Bui05rNDc2UjW9h+/Nv92BM/vA0zbrGeLz4Vtlyfbg3nas3aLnnDtzPslP
wwrt4q+2EODopj9e3aJwORyfvZ5doD1ktJByDGkqWYwcNqwU6qWw4+FiQIFwyjGC
u2wPJAAzB54RxhnBNjwfKrE0hTRGpZjzxGggHP1rJtmxQ7MnnJDmyeJjJ5QZr2Pe
7QnrcEN++hmffSeLep0iXQxfEIvU0O6PmrzB1Yxybdfymmp5sXgcJ7DrONs6F+Rh
VfcjGnNJDR8ga0NtcvrxVQwbYRtEp2u8OxWeq6y+HDPJcYZE+IdPqB2paaGgnoFH
w2T60jR/pk1+wpn61AZUzkEWntETzsIHANK/MLdx2uToKhoHQpuMIPPRIqPcU/Cj
vCr7RuSn94zxIbLVPqU0h9n00c1HJuoM/Cb3u5sbbQWjOw4T82tuslxzbZ4b4V3V
4dX8ZYRKcdVwBnGSQwJKDLY6wpBSw63W353pjSKcNcWI1bzxBYzpDV1kIJX8AFl/
LKTDyvgbTjrZkFl24M/inWok/9yEEsNpUbKz1GZD91OscbJgOwdMbcZ9M0AVnbb/
ZSmOmO0VVLa8btbyiT6+dDPQZwzcmVRfUH71fAn2ih8cyIW3ZJ7NnPSJhKHz9t5k
N6fCvw2zQtm6QsMRWue69QAoGgaTnZ2xWRtFYPRTMDHsiwxp1b1X6Raobg8EZu3x
NcxXY/9vrq1fhM0nPOr6ggZR/jdedsB44wCBs9ugJeBcUKX7HMVEoh0mD7eCphTd
Utn/CzYQCqgBNn+15ex+hJmgytmQHS7MxILCd38nJEWZIPIo6Mmhvn+rbMHdREUJ
gzujlzkJXEmSCWYmU1/v6n6kpMAkQQVnonOh2ahGDw6XcSe/VechnPTu2IPklBzq
z/lNNgzVxkXU7CeWoi6/KuNJIVtO7NmvvN+ZYwiYw4tXWSWxsQGqxT7ZG8SWN+fe
2boe485r/pFF43Hxn4rDNCXknQvK9OppyxPDy8c3Aa0Lo9obswtARf0HZYa0j4kE
1BiFyt7/GnSQ9eXgHFqrGOBvbohCDmLf1DmTPj9Mzh0E1MVOS4fqkJ2iTPvVmYTO
MlxrAhjj/hLu5SxJ1EDvZmvDksAd1bXtDgZm2QmsXl1DORLt3L15jMEIJQsrUht5
O4zSMpCx7QbeOhdj9SVtktSy1lZlWzX+BWagZ/rLS8hToubWNDYkxAiFn5T5hbPT
mQrWeM0idiaOuolzLoOasf0vq4fpYx8CTclDlYgBb/rSbL3vhc0HwSkhMUKYi28f
7mwfoOnKWIc9bpGyxpFWcrciFQfW6pL5/norkpUrNfFPdDKl0fAB+w4tcYi3rK7x
fmaF4rTaeQIPkvwEVkSoaXQ3UPT5vyc5wGVBuyFnJv0byV+KD+yBAjcdtxxUxuSo
VVuWBEwco5QeBZ6Eq0yWYUSAqAt/MHb1xXog3mJORnWyMnOrmWPXb7lZHfL9SwWw
oZwnSJE1891OYLOmqVEjyGt6KIOTUcQM75rA2V28icytOkmdAQxLVxqZbiertImG
Xgq/v2ydRLdfydFu3Uc6YQ4UfBcx7BI9N1Yxs8POlmD2JzaWK8YEERAsjpTHDWEQ
1oMvUH6WUJfqAEGsHsyrNf1wk0pMc+5pjvgYkiCyqOgFLVHht0NhzCohyMidRevW
nh+syLgPwEUbJAZ5Y49l55Mlavg1h+Iw3dJF+HVTD/if9/uIjzQUmWS4YYmGYZqq
bdPBdJCgNOwS2Z14qRtMYAT2TKUrXTPLkaiSMwMAmh1NKfBvx785GKBN04YbDIZZ
XIeU9g26dOX8HhvJrvrP8HQ5esexUHr03GjFWXXX8yhosSd1dxWEXCRpCUjzW2M6
XFKBwfD6tT8VSGe8fWGSLPpf0Sl5BrCrv5/F19SyVPk71jS/S9LVIC7wLmT4gr5s
iJdeTSdAXIl2PQXP0VWgbprRXG3/nSR/RNtVLGhCDQ9LrdEuAXHP7C+ggkJz4dqn
UL+Rtb+M4uuXITijojKHFjLakWLeP6QMj75pNQrCyT/iPPA9S0AtNdtrGdm4weAu
5R/mx4dWaCYfeITGUYu0b/BYOhyOriP7FTwckmxoGRQHf0ys4+80V/Wp0Fv+Ldk7
kuyQRixVOn578YrQKc1yGjFqPBfosZ2JnTQj/gZjfQJvYSQW8VathF8RHx5UV2Xl
gjfhnfLXIEUhNkqiC8+IayJlc5hTe17bLbNpBXRk+1qkEs/SkQiqW4+lZ/bHMl++
IxdJS4elbSK+RX+eZk85lw1yf7SsrOEeiKKtQt+/zB79EU1yJUqqUPC/K+GTWOdn
cohfzPhsMwYIKckEWiXsbJf1XRCStHK6Lo6E9KX7BH+kQZjnwoA4IloydyQ/JW4X
VlXjR7zKBkvnTVcGBNsuBqnpdMjt0wDw1N0b+AhPzMyPhDyuw/wPIB6jR/+iTCyS
KUJRu0iliqKoBTxYKw7vRt6c0kHTOZ5u+/WxvuxFgWSIv7zOVvz/K8mn0LkpojuF
z2b4mxzSefDyELM0M++QQ870vjZzRDNc5jaV5vgMumZx4TfhKG4E1sD4fcD2JnEO
tfP1+kKflii7D7JZOtIVK2q/oMQv0nDwVbQOupW4mf2tRNa6blBZBGfTkR8+QWXP
qnXWUlDdX63d1xRFoaD72AmI/uZ/vdj6Jt3zCiBLEIWEq3FXXoBBYb9Q/4/aYn7x
cltGI8zDhSBZzKiIcUNyVeLgnVvhg3MVo9RWBhTBYyx3ayjzFGNNnbTq2X2di2Cm
z9whPkv3hfCbns00IOGr8p7PiVUS1Zm7oUzqRRZkON/gZcoOZIHqiiMKGxMFa/ub
QmnW4VGRgKhcHNc9Wpaw8Z6gPCS6vTZfLofoWefgOTPBh5NKu+Zhj/vVOK8/oXbb
zmZaypI5TVwbGzDu//MboKWb/yo9RiDMRYOCa7jKh6Aukzcsl8ZDLokamdSlmhD9
/gcNbWDBNoTfAH7jtuEHs4Qgxl9B4mvDG28MJNwO+uAswJDdTtdWAP+RrGmWFJ6k
bL/4Ul7S5y2KOkJGYWXpp7O/61gyO2/TdaJ0R/GGOMfxupySKeccwsg0htaH3Q/p
sCLp2DsT1byx5bYw+LoFXjvhWmSBGWEfKomYbmsBAYiGiBD4RTioYKrmU7fES5Cn
slrliE2hgwCkP7FYzjW9g20HtwnyCJyLzpExKvbzI8LIoUOqZlj4kjAddVZeskmc
jTID2PcrsaYx1pDuoBm31wbU4B6m8ritluxm2D+VZ0EuJp29zMXXa17Vq5NELPaH
htptH0BnwARHkskFVjq0mAFv2+vqlSnbyGIolUYVD4bX/hBqDiPMHUX9SIRjmThE
DwSECgq6UChbnOuSh9bD5TqNfiwp3303+H4l2t+AOQOge5+YwV2N1vwEL5R64O1h
VPmX62odAQn2nmKHkxSVbGq85vfhguyWyjapE7KoLOPJ3UGYChjZvuBcdzpELzNy
C8o4dtlor+bmW6ku1A52olacS7qwO5d/YEDjO1qCgTNq8IFAGO8zUnYmgEnGtJFq
IJMvQvlTKMexiHOyhF56H4xjb01NmiTFKZSjakVkU7AsavLz0/2dzarQoRLi7MaR
dw2E/ciHBmU8Dm57jJdyy/s0gFjVZ+mQLgZc3TEey0a2auTRPltLZh0FiZ2EwwKF
YK/yZ2OD+5gmtQawN0nRaSXjh95T+TxVoK3GwtmLGdHEaegWt7BJcvEwyoHLcK7m
zh2xh7W/+YanHpUKXtIWMyJ8PIn8CadEEy3PGfWjuzlQB86+9mvxa1B2ltwgpvSs
DrhSc1JrwgWZEUaaVebi182A6IDTmBsm/0/0XD2ThlwVrRNUEeUGpeLQ2lC+QBsd
xgfq3UDm5dCwqXuaZ6g7ETmpXvh5yrTA6AaMsOO3boSabrGmRnAsJrkqfYCTc1le
4HSOWQStbK9n1LqF5f+eHUx1xCBkDZYls03M6CKOcmUBKntC13quKpyB2R/GsL3f
d1y9vvck5VH2DqYqo/Sp0Ul8tNdKF2VSkiUd0tOHlrTNakeaST0V81Q+fff8NGwF
E3Kq49pCMJyHMRTihFl+SpX6i4PDe1n+tr8nIP/EgPYcIb7Ktno09vWhTu49C8Rw
DL7lsqoPpkr7VJU6jAC8aKIIqK9BKF35ZrCtr+b2yJ/K670t98KM+EowLme+pttk
Yjas9DgGu5e7tiv4H7q1rLAmG25mzZeek/XEVv93FrPJ29eaMpwb/pAVUebXtWuZ
fVgYa9UPD0no3fvZmarwNxvkBSjPO7zXCLr4pHfZJT48SJc7AdOBDP0MsBFmtXlN
C6W8ctxJGfIaxLOFTzdDCUAeW68W3mRFc5IkopztiH7ojwj32PNnByP0tLFRxZpT
jcX8Yky2aFr8TsiXW6yXUWavmFu6hRCDtm/g4Az7m7tGag/sOu/EW6R1AhUO7pTP
x7cS6maK6U+5pZG5XfqyS+CCBLmKLuWqOrCHuvIkf1jcHfjUoBlFt1lCsrDioD4j
SiiGCn8PgB/JGVAxLrOJhRN5Q9C8iV9HKRCengAvwQIV81kOnO6qLHv37wOIfF1s
5uUHRcxZposVcekMqlzEQVoY22vFWW2YB82MyzarlFI+t4fL1ER038M86xMna/tR
fZ3mUUmx3M5YLhNuZjVnNEj3cJYdMa8vCTc+pruBzXWUx5LfME1i6F8UNpqg99EV
p2qL2KyfUVq2UgMD6gYxpKI4RF24PMPCKyGqzG9A5zURfoJMtGs23AdAafOJSxyZ
27KBRhwbXuLdSmTJyPwNeYQq0cVseoZJm4WAhWeaEo0H6MC6FfiRZ1z1REu11qek
4TUs19vnS2Z2mTVLDJaVdAxWwEvDlIAfSsjVLzpMlNEMZB57q9aGhCMvc/obUDu4
Cr4sqw7PF8nod1GDVWjMUnbiNCgPxIiX52YIm/B36YaoleSsgr7jg5O/QiBbGtMb
cfGhDXsLS/kSdYaSwgYL5kSdihcwa961m9nwJ+iKYlB05QoMSkAaEpsjEYH5yfgg
248bRS+3rH9Ub6ep+2676DCSXGFNkw0iPwcdNF0jagZaPMWVixwl9xJsdvHSrBrO
056iCp4s80DC4q+hDWfPh4fVDcD1Q5U//WLw5AjEJBlZEi/n5Edqm1zQnfxjTdM2
j5NHi+H2Vmun0hX8egpzTv0Ml8pGpsAh6Mf+cdGciZTR9iCzPxotxdmF+M0890dW
81hqzU/0jMVIigL2jktI4fMsqvDI+RMuK5Cy3qAtSUz+ScL+MO3W0NEN3AbOH2RK
vM7wAyEMIJf/1SDnVj4pMTN/0MAtSUvUuQK+HfUWqwtIeBET1keoKms2463ZoGI6
nanqQquwIxLXYxqQpf9sqzCHwXdbbG9mBlAkBRG71hl3CKQiiVOgRseSx5jO252Y
UN0SESphLJwzik1lAhTwiKiczl+BSQXib0Ki5jSO/W7xe+DrxKgUc54wuQf4x62x
34p93+tTgO2wOw35fkJ+IIfUWmPI6s0jgS+8SHFFF1iji8mQYtWhzIjWXjBgm96z
tHuUhqW1QwdkMlib0RK6Gj8mL1abk2odaPzELAcuDwSMi1xoTn6kzfl5DsozRqQa
QwdbfwDnCF9SYlof1+gdn7zAMRx0m7vGTnufT08S9eE4oVOWjJc38cc9UCV6TsXB
3D2SXeoB5U15bTT3jNZYQrvmLkw/4h68pL4IbeNzjN+/OGDs573+Hc1YgHvPg46V
FRlE7QkXkm0g4t80TgwG8QbJJtEiaHwqvpEDOJA6PkFZuoZs2myExSvD7BbyBewp
kvcdCYF/2Vl8b1+G0nz1+TNQY+onfpiZ3Jvo4UZzhwcyaKFSZmaXxub72gKnzIoL
cCIipammH6oNQW5xaxGLII2GJvUaClg3WZRhk403HR7NfmVjTtwNrKVtYFt/MwgU
zlfrkZhekr2iYig8hsnsqrfCyCZ8819ZH0c7rmZabUUiORPkzwmMEUhwCP7hjaJY
j/Dn36pnjIM9jLrXZxvBq+TZ7A2Hx/MeM3JHGDj/L2CGGzSwUfV8UXFecBsbF2TN
4rAQ5g62TbczOzdZu+P48iuvPiZ9z4x6lmdux3wvYefoNOzFVsSTmj+UP/bf0Aia
7aYCr8ZewT0dMXwTNLy0IQPPcnEd/v+KgkXGkLm8KStJrCc38iyWZGNbxvezc+c9
Vizj0gAhmQduy9eF+Gw4+Iy5SVjxsRWDpoDOjCRutMP2cTJ8DdY7Jx/80pZVc7Ti
LOBzMFT1gBw8ikX3xxVp1yyNTwiSiGZ3UDKxzdKkMWDbYz+2Hvpso89vVu3eJksh
+0lHqiVojulbvav0FzzckuyFqs036Non0ur8o9pbz7e4uGcpQI9HPgXAaqsIgs03
Mzuiv5Yfw5f1JJ93pGM0qCrAruP+JosISAhYnvo9Z7h6sFmsv8VIa1jbBO5lZFQi
IB5wNzslH/4iLTfICOlbYjRIjbA9QyCBDkraXsGNzqI9aZ3H/JJLrSrx3H/WUeLU
ys77YGV3YOQ6RzWf5LZbDW3FOJPgvGdGH9lQ0scVOTluRqP/eLfx30p1Kl09WQg7
Ax4VJ3rKVY4WJANahveIbpZM1XpnoVlYste96PvZdo39bmDQYvFiLn1Nw0MhV3A9
ySTUQctZQCI4vg/TH9Jx7xnvZRWM0ghjRvCo0CBeQT2g3hOlzeZ0RGBbtJMHeVo6
hyBALiqrVCWIBRN9PByw0BoYYHbZbYYrpvDgSLeWDLjq60etMSXMLBjEwqU/zFqL
EoM7zI8e2th12Yo/d3eusMR3olJVv3jri0xp+0+q1WYeBvPdst8+WLFxDRP9+4BL
8L5XZXr7JVHL417MjT73CPnUBbejYRiYw7vEcdy5E6wT8a0TiMEdmqg+VgVdJ5rh
h8siPsfctFv7UTc4lUg5P04tOb2A4y+Sultfty1b2UX3ni12CAW3cXJu11kfBXq9
/K4a0DdRZV2kSbuX0Y5JEVU4akOgo0FfG040Pctl5KQKzdTACl7Y4asKBAowTvbl
iK6X5UHbVQnSFg1Asob6oD4DbyBvViTka3DDH2e7i0R3dOkjP/bbVFHszrjLX0Z3
Q5ILCCy7zqD3Ly3T/s+IVYJGVIIopGX4xZqY9kwHvf6+8+oOhFD2JXuM68fPPzrw
WBAS9ZRwQGqkj1mZrfDbdl2hQPHGIxfpV+ychzXCycNCl7h1Sh2HM394QVP6W/88
cUspN47u2GoImgyAxf4dkhJ3o4RhGlJx6A/Tv6w67rZB8PgxMxtXf0oXT0eWt8DQ
g9RGL6y1LXKzZ07DBo+rzyvvLyujgDQibcrcDnf9d/KnBJNPgIsXuCTqFMXvHSaM
96NGhq90rnWCzxz0b8CGOTwkHumqMoUMl0e5RUbqhAl1lzTPio20F9k9xosfwHOv
QYdS7lE3FQ7rfLzRZlt+OFQZUiv1mce2zDytr0LAM/cQAvPZnhMNA8H6s7hezr1/
KfPTfqZCWtzT4/SIOfb4h7OQpPGLJkN0jknnjXY5nBzj6PB8PzScdv+ioBMUkZKI
Lc04TEd0xgHbgSO1d0TmOTSKwFNgXhT53DGMnUGnBk6JbbNZDJo7bUHQL54nE4k+
NhOCyQx+4dovbUApaxERn49K47p4SuZ+aTJNa+sey8aBF066fLjn4DDwbqFOAUEf
jS51k/qiK2Z2PPajXOZwDTHUdQjz9jkjUwHl9TE3ceMWJp0AB5hDpTMH/OvYU0u3
44eT4/U1OJLXK/l9/Lnux71sc8yzHwaXzUftRswLOCy4qfZ5FhBr09GucOLRL5LW
T9H7qPyKeowRzjVVHMrz+3mf0YdpZBesBxhnHPIgm3aZNXGbviXyTiuJREg14Aaz
1ThuVH1eqSBh3spdC3m0JBT2NTX293sZlcQat+ceyT+Ik8Hnoo1GE2yWXPEHgPVj
OjwG2Hky3u6BMnVrUtKuLUWjTmDVRJx/3YG/4o6CwYAbRv3fvwpEqjoy4Prj1hZs
XUkiv2ZpuxD6hLZXeeZEdkvFKsHw3Ne1sBb4EcFX4a+P9Fqg4JQXd7dZcZ44vCnK
ZvP8CrpVgiLowPNJz900nOTqEhLAjLfdkeAhZ0cQ8LNfXRN5yd2u4m9OX9Qka7jA
F3FM4eXHH+nFNuABE3zuHT8VfjwI9dy/Qf7llQbutRvuuI1TJEgdvQXAUiaVKNwW
aaiJEudQ7wd/+rnQqoXpsZ2u8B7qyXv1QJB01ENZNpaXsibAHjQfZvDcx0RUK9+5
rQoE9hK1tGdyrW3Epoe6A9AE+TXEwSX0Dr4xB6IGHdrOPzfWnZIIOC4kGJHyElJx
zDOCKWCeE6sSD0ioAFVBSWJCnkaFV3qbYy/nc/+pU3HW0FCE0yCyhfJibDAUWndo
m1o0zbBETNzSqOREN3L5U2mlT4IdsWxvWM6nzFiv0byBheqqf9Y/KtQJYvZMmUW/
ayDbu//HBZkdLpRVo/uK/n7t4J2OL8F/+u68Ld7I+AoEaTh8saTmz3wP41i1jXkN
ZG92UqFnHpDTcGQ+RW980yFeZs7bCKHFV6q0gMqkoOZgl21cy40LX6Si+kiVboiT
snjX+n6dwEc/8Hgkejhpt/hf6nPKC9iHyJuXFFAP+zwz02osu+mMSU7iBG09UJ87
pPIOZUpGCjJT8GWDkPsKuAxpd+ZDaV7sjDV5f6/8ZuBctI5954BtITaVl8KHqUmr
I7m19VHa0aG53oSBjHUXeVxR4yYrlIDOv6P1tSBN99zcHYjYim0sWmSLvULx67Un
JBsieRhL4uHXFkWTQhsorPTg6xF6hcLYozqyPhhy9wdkZ1RXU11lLMOljcd6xp9p
vWyynM8x1oT9N69i0XIa6xkMkvQC/n464QWNcAbl5Ia7tuOhh6u+B2eZGEDjkKoz
oCLo9ZiLxGjUwl4+qi4gEAkuRNxScPix5WzScs0V8ZJ4Up3JW+t5x8FQ+AZhUZ34
EiSBsFE8tLlgzJCoRYU/B/MXrxgcafILO4TwfkW8NnFAg80Yv6Jm1S1bzeSD1n3D
zAs2DeOvGj38ONWn7dWDMWASqJ+fR4hOfcDt/J9UXyQfxhfXIzvuQiTn0aueYLN/
3XrWzKV68hySRAuzdGr7RhykV+9zPsqAIU5zPKNJO41MI2i+qbs0Rq7D9cS7iu1B
aWvyoSVtI/5yAquWE2/DRUbKtbcLgJtWV6oKcaImVxYlX+Kmt0g1aWY1C7a+zPk6
i7IxouIoUzWXYf6Ta50dw83rMwigRHq3bJSa02bS2kBt8dtgyHThDwGYt7ih1AY3
13WSvLwFc2EXG89HUu220De1cdJkwZM/gQrkfftl9BGVu+W5dOaBEAROrx+YqZJg
JDyB3ctR5unMInOCDMMkgQ+7rGfx+EIcvUJ2cz7vSE5JNK0gd0hHuevZqyZb36Mt
AElpP8VRsP3QgNDEf9RI9fXFo7nKPCyCfv/wqAUT9+Ql4IXm+WL+UjEUQA8fVk4S
`pragma protect end_protected
