// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OSU7SXqXwzirDLe0qRTdEfxI/xBjreeYasev9oKwr8ln0NMdtbRnaTjJo3tG6qYH
WNuuX6bEZ2wZJ1NMso0NdVX9W8BQSsFC9UZSID+vvrFetKz+lTV4Jdn5vgkNxLlq
UOESq4k/yqgqJvjzDXuiDjIda9I2yxe2RUooOgwjZRU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5536)
2JpMVTck6akd8t9NUsj4FhyEnc80ubRqp0OJbLRVV1VCHDPVyipo0q7cmKA/+ywm
9F5HBaAJYzAVF7FjvWKMW+UvKhA5Zd/8kOzn315NqaAZTNkqSD4vDkyhc63tkNTF
digQUfFCwy9QFdXYLMDHHATDjZ4BLuz9xEEi8yP81j4+L57opK00Z229Rc/XcECH
khWapAwgODvJFUKagq6fUyWU1iofcYp1ITvZxg3pykbUCHwDwE7InFVLsX+W39pN
bB7vqkaadNfEXxAAaBxXL8dr/vfaG0Jsk/NYdTXPESriHU+p8deEhvGTfOJZqoIQ
1jxyYWPMYALLWF/H0Sgwj0takXwj2V8qFhz7HyLVFOJA+9Fu6G4XfYaOj+mGQ/Z8
4HxUjBo/UsNoqAcZ26hdsRZK7dermQGyHB5HS42u4gTniM8LCGGn19LltsqWwFJ0
uEqFBopNEsr23jKdMqCDqY2K9IXea3Z1warPIRfQrzw5djWjagC/G353vhbE8s32
Cxd9pvjZErTqgdO49WG9yEELNYI6d9gxcDFpFZCs9eXjrTPuVawF8jETuu7PxAog
/V8moqU2uk3bzUfV/QBM/SNSpWetHpThEYdrcCwLLM6GhaGe1pCAeA714IFu8TZx
bEuprwBr1m5fTwVZVFXiI5UqujQ5zL303uzvnee3FYoR53brBTDmROXdrkqkAB5t
tKer/NlN/DvJnn1NLOGKuHcIQ8iUmR7NpsJpqPHCrWZUSl0L3mL5TgRiEE5E/kIj
993oK77y3Oba6y4D4iVbtKxbijjA+Vrt3Bp/UqMomo/n44WEJnuzjjEPP2W6j20D
L4YPfWw3t6P86qf8F5FHKvSO1ulLHKYHWvKCbHIByyrZKCVIf6oIOQ0df2G+aVxT
AnAvYhfbW1a04vW20t9YI/qUH28wKbGzCCLWy4RdvfAzmwesXaqhbD0h93C0mQzi
ysSf9kX8ZYwQq235zXzNg5rR1m3VVCS/3aGBIew0GbyB9C/k5/aT9qbSSeOEcTl3
Oo8iD0JeYDo3GRx3e3KRzHgcAuiaVu8crz8vmGq1jXZeFsPAhcB4ALtq0zr/d/jj
vm6fy+B1JJhLBx/6uKZtDfyMgaeN/yQw6mX+umrRi33dbFg4LxPgSDPjb8oNGrer
oUYuxHVHfivBnYmTljVeR5XjAn2q5YSNe4l5CJ3NCihA1tqUHKukaSsT5CUi2NRZ
B+jMDCbEb+0zDj3YPIcgdLxd6+P7GxUy1FL4GmP+2Bt/Nh5sHnosxvwLT5l17cD0
R7KM1QkCZDq5qKQFI81+oaE+udFb6j4/9Tk2PXmUgCpbcaj0f2RlApX1ZN/kigiT
PfXzbHN7OsZ8jmw25LmadhtPkHfrUUKpyMC2rrsnnWQttY28ePeHyt+fbIeJ4VNv
NUujT4liEl2okYRVawk4ljcoHQYE+HBZ+G2Iuz9vxZ2Q2GYbb1uCEVMVIOgEsHuv
xXCC+W9wAoHeXw9wCDeu6fZ2Aui2hGr+H7ifYxL7OIZPm1kT//iKTEDMBtJQTuCs
egpSl2XjIXpH89Bc22J6OMiGgULtUYwUC+Ezc2ySCfPmwAKkVwoSlXboeSPkr2Um
umkhhB4t5mox8YM18QqE+IlSKDhaX1oQA8VQyoLib5wYtBY4EUcG8NfYbm4xgxyX
t52V0ZiA1PxUW4RNpxNcF1Pfy8LSLXpEkX31q43MvpG+fvVyn8YJKnsJkRODl5Jm
tftinkn7wOZ37HyPb1hQl3pc1R0/ArjWyqfJtIb7ZZnCVdgqhKlHMqPqqJEclnkE
ZXeCgow2MYhVUYvZmb3WqAbKJoum3dH01NTOrjwC4RpFipq9VUyUmPgfbbMdhelz
CqOEEfpXjo5JFi3+xtOFJxkFXA/dqJdEzhGK/9p/0jQTzsBsiTVWFz28Over3LPD
MT0PuUnt1jiiPMLKMb5KRGngMRdS4gMFhE0hXXxWHFA+ud0+Odit0qllwqeR7xPU
04JhlF3Bb0WBgRbc+V/EtzRdmpTQG+x2XBRTcqG6Y/XXhIU3Ph1Lp+EP5fua7tI7
wj4GoVbG/XFfGn29gV9KHc/75Occ2Za/xkF5Zn+tn+mcKtWmtou0eZgEtOvnwoOd
I1CIapJpdNzP0HaZ6jqbgoBJcEHY9TbuX7TbAb78bdOI6mqUS/xfnKfcH8jvw7RZ
JpNJTABeuCxZk3PqEAAih54xxtoDm5p3aBLxmw7mtkoqGHMhvA7twAhDoU0BGTNW
JzGfy+R+YiwTj2ki9n1n0dwKyNMorLlVGh/29d5hf4LlFAFJSDTi+TdbwQayLUqE
dcKJCqg9tqKua7Sc0RpPNfxIH7Uf4H2PhQGMFZKwCAoi6XxH2y5zYMlw/FaBJaEB
X8h6A8MOntEB8dHSqH3d8OVdtXsxc7WK4EhyD3BUqMXY/QwbCaUmMEY+MCqCU1Rs
W0OImsE9TgebI5ICtgxdDYnHMkE3h31WBnNO3kXKGhJlLGbd/jyLQfuVomjmA/HF
7vHwl3MdNRaQtu4FGA+uMZ7JimQw+8QPH7MN7grXSdsK038IpYLOxzMUuyHZypJk
2QdNl3hDHTz0GmxBQFpmZxul7V6uRHrD3tlen3/6/SRm0Fo00TZbY1RQr6wjLAAD
Kz34ELpj4y3Xw1Tiy/TkBrmQc/r5m5FOMaqhQGMByuI7f5hMszgsFnIPgxOWfQW9
0h7eOxoHPiOJ6mE1QQEe8/5I+HH0HVyjp+QTUn4QURuB7bFMU/IkC7j3jbTXn6aU
x4ow4oF0R57V+xWkYs/IzWCM/iM4du7wkH6OTX3BNZ8HnVEwsj0+0MpbQ0hnf0ww
ibXb3HAwUaxY093Qvd9ORQ/3uyDZxLqy8eyzN4nxiirymqkyS3sQ3D4HzpOzA+m2
Vr9g6al28poi3NboTqA3PnhcW5e114FPHDSGs7HwMMz9Dso9l74krkfab8aytW+M
LDTrvuR5EFVZupK+CkJ4eoLrrFSiU3a3+oA5XL20G5gQS3z9EjGB1STW4N0qR4zv
x6Haswo28WODMZibJ044ZOOcjmWDLp8gPFdf7hUSZUwG2rkgCuwHP8YLz9kEOZey
RUzW3WRDSatUGjew/W+bDO5IBkO9vjsrCd2bUw5jdA/1tLz2dweOY7a7lP65Xl8t
0lba0gmbviZl1T0XCGFijspP1b2HJpaHXMoo/FGjzYuGjaQ0vnbS4ic524NI6iGM
zdjbUEg8Sy2qgOtg/MjjB76Jww5YGrV76B90z2/GHG2WqpieQXlH5jCZxVSk5EDT
hd0oHhvg8b+0mkOGoXKw9vx0+Q1trkI++6nbKuKTlI6BR8qH1DaHWLhCdqUXPFok
g4tZ6K2Y0bokB/LfKKJN9hRy5IJ79pzFOUqZ2KqnZjmbf7pmxxLHQ4naldqLTIJq
Jo1Cnr0rhrAhVxHWTR+wkkQZDGfLriLaEZHjvgmDL3mZ6jOkSxG+2KkR9gAJrj5d
rTMDjdD4g1s3indeoC4mgDBxU7TRJ6+buNfZh5FZXa5Ostd9c6R/8RaAQ5V8jcT+
+ICWdAKGyQZ3OFg7AufWXmwdHePsA/vdnjEv1Mz65zOYLRMbRNx09DcjBZuMbbhS
9IcvS+UU2hqSvOjx7DCFivMP36STQL1ydikk4Eu7NqOvTX1ITRwpnzXWCdOzBV7f
wMcDkIOlWwSNN2TzTAdiT+OTDsB198lWEiADAxcQs4l6D8zrimHkwDzMOJPQrofg
O+Sq10LiGejG0pdQm91kHnESK71A+D/Ev/BXWyge6R7TcH6XDgfAjUAUyvCKg35X
fINRjtWJwNXrCvvi8KxoC0S6VZeVoIChGR8IWZGJY1CBpFxeSWbEfJghrY+7zUMy
wstGT2AQ/8jxbE8dmkeCHXQfk5RayNNxThVdvsG89+iE/iNp5Wt+8lm0+eKGS5l4
oxgykYJli/2pePtpP1nJqjwYqbIBH89XX8xyfUSyBZ6mkxOEC1q52jKNyw/xj3rf
CcRUGh1tQMVhCHu67vSSTOyHuClkXAg1GaxAYrWBtkIGSHetdpdzgyYTd/Z92AeV
emySN5vxZt+GzNfKqVFEppI5OyLTFa6EyWtiE+8Yvf2xTCe89y/c25KTnwyKVC49
P1hy2yliJ+kd5jOzJl/s7J72ezfpi73pHDdYh2JSAN7efio9FgQRmDhhDsEcWkUf
mFCWDQ0WtF6L56u9L5PQ3j5bMjJ3n6qmaw31ip1NZ1gk90PFgi43RqtUqURAGlK9
i7h6L6lpHYyd77rxaTSRnOb7jEtizBMJLs5Rlzp0AvHTjthL7Zr7Hu56cEzKY4u3
du5vNjRsEYRPQaNP/61IWR3/a/ddjfIxxq3R3VyiPd655c7FVzYUvM2JX8mDXqRM
DWWtD7ljYd+Nb2iQAbctRm7Yn2uSpOWAyUSyrcE8PejXvQtuOydP3mBNMDaHzPkk
qGEG8qA/x9cNN7qcw5dNsByqD9M0JB4FoqOkxkvnqWfFzDWP2qvCKwglhk7x5feN
cB4LQRH4m26lHeqZMbfC2zF3OzTNkTWloFH77VhnuxL5qGTAIA1u1hx91360io0q
jl1EBm3W2ENvOuKnTevift9U0ITbA8AFwz2yoJgVHXQSXi+H9ZoF+8Nm6ICCJcfs
gjN42YiX1RXRCFO5o8wASgFbuc8qVmpjY4dOHmvSl/m8sa8neV0fLLAJZ/ZEsqtd
ARe8DK1V9sLLkvUWHBkx1+36GICcuogTXQAbmyack+61fATLHu7oOfuzVq4keOpA
gjAvOizSHmSqxiPe6ZiZDuX2GjkVZMFtQuePR7951WW74NedcAXHJJqfMYtB6fQu
G335QYZ74mFktkNlL+T55xfqy0TXuJBQl5eBUaKtzslmJChXGZpT+IHgHJah2wbY
1OojF5dmhXWh5sw2ID0McKxirffHd/fYxHYaw2c4wLJBshPI4GdQqmJ4ko2Ws6S4
JSsLKu9ywoJJCbA8uk0lZ/xTtye+Q5edt0X2+M3jfsTWwMMWg6W6Tn/fZ0FyFzPD
JNOi0Yn/kGrHl0H0nVO8zBxRTj5HiXFQ4RchUnKZrLGuhHZlXLFUVWOBV1s1oof6
MjeCJhu1eaYtow1PJAgGHh1fLi/z8izLBeyy9GYj0F1SKhkmzeDgY7M7MWnPjZ15
2/E7M/rVrPFYQg1srrD2cfki9BIIzgdrxehDRWS6mBcMdJAxeZPNm4tXNPZmqdLc
tJVvn4uSr39FR75xDDgSM4aKhndNAEPJqIfTUiQfp56z1sV8i4CsyKzcalyG8i4f
9qhYjdwGvV+eeVjD4WxwBuXix0SjT8KpKL0ugJm5o5DlRMVXtP1382RZXuqGzBCc
Cden0aSdpeyo5P4jCWLlo/ypcd1JbLPhtd84+2nkCToeTMlmNBYU+A1kV8qvquNH
GZ0Z09H1EcnVHAEYdr64bLeNsxp4ZMYG8sJjIf5jZ7fbc6fgipYeG58YvD6ADQu6
5VN/uNBTTlXCA4u4E/2+sd1upaMVsGT8jC9ivmZYPRIX+ah4zacIU0ae1SnCVKFF
Ti+I6Q11XAYSx7p7hm7MMLVWv3Kpx32Jv0ZLErJKYmfwMFIb1ZBs8NpDguIGjAWC
NjnLNsBVMfwjRDpjax+DHcePiEmCxfA+R2ZkOo5z0PxC4EFGK+pYtz71qOVViWEA
g/g09LAy3q3ZAAnxmHANdd9kufRhZb6do2HStjFrCrrgUMZbU4/qXT74URvy20oe
vvGnCyQkSJ9IX4LkrSBfFPw20E5jeajsWeD/019KX+638Zjyc4cX5zLyGahWZAkB
5aQ7ZVS27SyyNufJpx1I6DS54VztBOESc7/VNaiIfYX9PKPUi94wNnJC4XtyFVoa
kWYKUULOaQpxDh/S+/gFVHKO6Ef5xPjYOATbPbruSuiXCUr0qfEZiFeAV4LODrQq
TwB66vxHgFwbbSxxJYGKT7uEyKN7BJKyIaNnVaYyB0Z6o8g6kluHU9vHOHAZ8FXF
KaELSFWW7VWouEyq6iKMcBK8j7jGJGJ8ryPkqLxUXQqKlbAJLo5ZnShay//4HlPN
h5+acFKVyq7Rx7aBSvOx0udBqA908Gd6u4SUVcdkXHOZ+7CIvjzKf5Sw3keOxrhe
rt9R6ftq1RmYjim7XA491pYbHFnYHXbTTQpS3pWr/MAKhnRxIyrg+eglyRcS8szZ
FWY+q678jqVWMRpt//4ynNxbcQr8WgyhMn8VgUFm9EqMcNIyNJBHfNiUxpWq4s8j
7QzBWkVukwHcHJM4tEwCk/tu0OlLXKYWmAyOP8PlpejN1FI/gWZ9Rz0u+jmN8Er2
XIBeOegTU7E1TOhZtGXiWjMGqCyaOO0ERgJQSYnLL3M76b8GPptuStCOj7GuusQ+
Icy1DUQ3JB62EVyMWXSt/ALbTwgbhlVu/73MrMWFmweJhERavJMsdXHd0/4vUFNc
oyOj8GkWvgCpC8Hk656w0bBI9ZBcC//FgDAn8bEexjPK4a1MA7kf3B+kUAuU6kej
F0s3UccI4JVO7TrnP+SaX/JBQAe5vjVbSVHhJG+cSw6RHCPiHWWl7MkZ2JzmJJE3
2pCtdOl09vZNyR5Je0EmxvGyhnA0zlovx2GwJcUOIzrYokd/2+XaLl4+BIZ7vREd
TI4dmwid7yo4k4ExIi8OfhXQp6gbHwrJfRjc7uDRqBY3ocb3HtzrImsZ9sI1PwvP
7nL/cVUKZ70qehlrZ+e2q6FxHD71PQs58Ldxp/y8bj6Fyay/HEpAmsY5SxqoAc9+
cNnzdDtFWntv3/g8H31zKCGlo1QcRJ5kUmzmNH9CZeeLgqC33KctFyVLrTF+bVp+
QHJRu4ubs5z+zFibBy/qiCgJFqzhjqo5qb41PTa1VlDnmseSwGMZ4QMf6uDEGLzF
XKmc2hVsoYsSGOFEXDxElW2j8FfZyklh0xuo1W6J4iId301H1Myg5u5rfdskLM86
VV9+hssQ9rFxNjg1JdaWCSOFSFmY5h3o3C4C+xE2IzwIw/SQDHxehFoIE2NKS+7N
hmJqeB56hwP9v5xxQcEnQ5KoDiT62qrLU4Clmek56Ne6beXR7G0ECnPEMnMdlgNV
TGTv9f4lE7QFRG0TJ7iqMKPlyutZ9p+WCF+upbvuW1Yjfc/wJf+cuZz/X4Hx6aIG
KbhEvshg62OjaWZxTM4LWyChVPtufHHBjiPJfc1yB3t6AmUenVQQNQrvKEmHDWrS
AMSZ69y3M57afcbD23m7nTlvCNZKfvxlZP/VhnUmt0EeQVk8fr7wLqhufO/mLJjj
uunceuHIipNtDcB4L2DbiDxxaA0me0kbzXwHDT2+CtV9b0b3M4iJhEwvbsvA96uc
wH84f8PJkozbEGigbY9p8ZynfUBlFhJrF+e0iprid7WEp+JdD0RGapU7zpr38e+r
8LiN2HmwwekXUB/rrgnyRg==
`pragma protect end_protected
