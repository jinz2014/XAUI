// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kYIxa9lrMuY5YzFFTmm5Ds579ZNU8kaIG+FHaXMr1lI90wyCr7x9o+/kqObkj2S3
mdT4TL/majdGNA7FTRc7twxg6XfUC1r2/BFFxWqoO7i+bjctX/KR0v9e4qYOZD4U
JdE6AB6ygxaClqIe8AW3XWIXIJr2R1DakejtAR6YmEY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 181040)
RYwcoq/G1hcujAL4oOcK/AzQRl4vx1dDpwCZJ1QiL5ncBaUA5uy+mTk5gXkoTocO
sSYaGhdyLWmBEAivlNC9kLt/KTAKDBSABMzjgNKtGj/K5wakVMmIvOrTeAq/x6SI
PEIqSiA9mlf542iFZ8Pe9QQ8GJICiHQJN+pj8Uxer8dxCWWUcOBYt2dz3+qBYqmh
27Y96iMY96UPKR+6mLhS2fjUdTfBE0T7YoG8Jpa/2eyLJDImkZwu7krMfeeF9x29
bTlqUcjbSk3IQA1/676jeC2sjwffjb6o7LgW/4xfE9fhd81Mxo+A7LyaYpqgi445
/rp+WjPctG6JO2lxQnnvPAyIyAuyJ6DkMx6zDLyrSbrKoVeOllLrULIi/mz5bXio
kuuhZX7DvAJVCSHCXQ3mjJM9lCLC31qiz96+D6MfuBCu/KIvEFflWpOO9TeRW9Cw
aRr94khX7sQvD93vRWbIRcZXWTwjSS2fdQKIjuvZ8yamQI7VT3SqauM4tprjSYX5
BIvPPgh+/h/+W4oqllIeADHZaj1/fP0Xl2IL5bINZwrfIPwYaGzEl5/blbFzuQ5t
JuSG64B775YFA7G6jooGHSZ0smumaZXPa1E0unakM6AAOqWQp3q4NQQTg7STqlek
KEVkPpbZLmAdn+RHcjKPyhVIstK48En5727P448+fdR317OtrIjUp8AoK05fktso
+FGiUOzhaWWPPalBkyRR8NsHKDXl1IRH+rwbtHhaZAeQtTdJpq4q1hjaQs1YsVDE
vzqJolPsSMO/Qwn3bEjfuaHLQsAN6EM93oGsCcma/ltZBvQbGFqHWQAQnq57DUd1
VprkxrFdipSKsevvQEHax7iwHssHRWNPlGgCJvQtoE9DPsPpnzKIiMW/E50iPBb4
yVE3HGkJ5DSrX5g74oagFowc3TP7nJ2Wry3L6XgwVioxrqgr71HA4NnPqAJ6J8gk
ekCVlPqLWGJwhsJDj5TOOlpeDkIBayT0E8R3cv14ef0wWlsVLtidE/z75P0fi50E
eqcX2RcmGI6uYXGUQqwRYSf9zmUap3b83d89Jj+t3Gq6cKVe2G3r/u9DVA+mkKyF
RkesNSXrYeTm/e6FomSwG72J9OnNbLdNWFqFg72K/crT+kL+NKPe9hITfYX0aUaV
c8CrUa9P143qCVKeaaIkvWIyUcTyUgPPykEGyCanZHYEojY7ZZBD+UBdrgy/ndu/
I68cmG/ODUGpaoNwLhZrfa7I+ePBpd8W878cwYAs3M3VFOLcqAtPS4kKiw4aPOU+
rtkmq48D/8L/GCHCNE/oD0Kocd2cD1D+sGxrXp19QZ7dKbFn/znY0De7lMr63S0j
CaCcBb4ugzTCnyQHkRMn6cokH3FDQoU6YcqzWJCur0zAb3A0AGg0Q7InHCwGFuc7
AL/vqOBJGEazWM67I+zIP8a0onEcpP29VwAQ6qpMsIUnFU5w9hQZTU17gtf4zWz+
m9VzA/9rprT+OIngcraeGv0nlHkBqCJsdXvnmiY7VzyYZZisVn/cJcorPsF/1RSQ
/OxsWYyc3t4PvTVQQ2//DtAL4CLRrCln94tfdCX+PjSHkq55VHh2w7o3jy2HlZ0F
ZVrKSaduM5eCJSSu1kEYqTuxHBAUEJAmfL3JV4KFP2OxSI43HnijaqysxIxtfPoT
d+B9Tahcb9PY7Hlg0BXlLW3pEdHHu7IKb2CARn/oXMETw57XxeBJSfJoymO8TLEl
y1b3awnKN8UrnpcnlnC1Bd1I2YJ8CudtxROaLonkqWG2Ij34VL2Ani001X9NHUv8
fYC/0UTnBm94X8SE0rNOD8BNW1BfZVrAavMQLJjkfJUNGVJJNHUKjrkMe1bgjRLo
aMzpH5eM1OifLS1SzcY0x05SFyHH4PhILovKg17s/CAl6LuODLySRHBHmkSs0sgj
E52r+pAsQTKI6IjmhZfcQ3EooaQjArPQu/TO4IWEFRgdUpmxy6Z89CkRTVLvc0Le
W8nPDSsTBPnefmF7YCAL2WvKwOwODYqkkj/l0PHN0eGkl7iIJgcD6kq4wRZYQxf2
SQNXE6HKAbUrhjn8ptqFvt/WdSD8Cw31WBMk1hko0YZOPCCPzG/e83NzF7HwTEsL
HLNpW4Sjs6Kf4JMbjXvugDK+V9EG3OS5l0L/x7NRWlkVsorJSzHvl1IRHy870lq9
w9yfS/axmxhz206TtKbhp0YZHLf3eNcZLG9qOIG8Az7JMqRnOr2jCI2RfJJPQBme
BfgBVkw/t6inymvWTU//ZaDWFptWvqpCRHmI65FJwsilqSuDjc5WSjPFBl4m98Cp
SMhwgcphAVxhGterYQmwC8a91LfGAWnW6tordHDkgv+BN35TNrgOJu1f/9k1paVD
C9dO/ISASXK6gac983UCFfhYdKA//NSwmOdR5s36Wd8r78dmSyRnFrfG4NDBqb2M
iCG9/H6ySGEmkH7e9sG4miBEDONQxJ6IE1xRg+yc3/1QJPzvcz/9LYd+CsdaZX3z
C1s44350gYxRmyzEmJfhN/65F/YEj21khnVUshc255ddml6DiZWIoXfMRldtSvwM
74rmZcJCcBBgLkP1nblM2HMt124Fcj+iKaEhEjbBn8vZ0jR7SdTdkTFr/E559mGi
oW94hpAA8ZJ0xL1UPltol8IY1+cT86/palPF2Xs7SRX3z67jkIav5H8Vah83fCm4
QaDwoQrHuAio/AUtl347M1hgu4KNQ9mGxiB33pgqS6NSgQkgdLEgwFRH/VWYKh+f
RtfT+3fxPb+qbJRAKpKabvaorDbdtRSGHOiv1hoRBeDA9vbU3zZhmwLbmlRRvyUK
xuMuAJTNzn8LhA5nDSIqoEJvOM81Ev9WsHztr0/1v4lLYHSFJ3BToRja/gXrmh6F
q/9R0OgxkbPhQDrElAADWNifKRPCuaKvMDaT+dcAMf6fEV7tT1ulik5vvY2frBD0
MMxz1lhsEpjc2IZDEOA9/HmyfESt5pJRQy5tPKoiXXlF0PWv+uUZr0Vc5Ly6yZ4B
PdfkViWvQm9NGY2BsBoEeivnFN1RuL+gnkjlajJyV/2uQ+QGh7OuOU9vp5o7Ap86
8/MQvkj+bqG2KiC65UBR4rLbh+ZiqQerU7Eet7AQhgfo9Kqe+EC2lL/q+EjSw1eF
MCXyuKgQkJHBG31Q4INq/oC3bMFRnMH9nZB9RDz9pO0Y0PyeHi3sMirxHs95wwFg
mn7gRfTi1y1BvP2t9lw0jn4DKkwuRBSfp7KxFgRhHFQ482tAHZ49whLfhtlqEn8W
NJ+YZIC75bJ2GLVnY4/r+HXms9jqfAP94AJTeDtCALHUme1J3cCWjP8xSCncTLzi
Pmro2jo6+ugoiVgRtxxTRyRUeIpsw7vNReFSegDiGNCdKB4j9bsbsmVq6QOu9Y5Z
IzGKyl5kpFDs1B1LEF29iWwZwZ8ctOFbnqqgZfsq/hPZ4bdbpWbfXn3U9sfvQ0Hj
ChVxwrDCx5Peu/sP7yIbDTbYiUAQ+5c2M6w0rrC6o+GqG+d8mU7qD9d2aH7PKB6i
0/PBIkPk0aI8HGE9ZUxLYjmHxmuRakgR2CyZ93QNoCPd7fOicIyJ8fLtJJjgglRC
sJkVy8tGLl8X/QKgnG3IxoojJv3KMcm5ACEPUtgaqZaN+MnyVbH4hzTe0CL0IJW8
9os5/3OW96RzOgHxFTopQpOufV/dTU39c47TYyWCscbOvlBAiesf7Al19sfhrzhx
vEjtT3RurQc1lqgMxdBNSHIY6yBHtd57ogjTQsng1FCIgxDUqknsbIOKndT0IK98
OXcUMG7TQP0OlEYDM3pfNP8qs8JCPQ8d9/bJR48rmUIeZLmBOiVm8QpP3F2Q7mi9
Op5EgwS+Dc7dSPLraHZNqxz9/jocreDfhLXv6GMfO6k3pH8eyNrvIiulQP2aSazi
2fOe2BwFxcwM+giQVgMBveqSZ4Z9fVrQu4232vd3J2swXNUhKTct3Nr/O4dfyal5
NMNCt/uOUU/PQM45lnKkFpAKHVivoEPbB52OWpBzE/JeVSpHRYi6tj+g3+P7wYK3
SccVGe3+6KivVjwtJqtGNPuiIr0ELev5F3i7LOmrRzCR2rhl5fnzZtb6hEYLmmMZ
zGbOoIAW6ZSaF9zduuROXQ7Jhl69bVfNcUWMCu+CuqOd1E8J4DoomuWKg4kvPcf0
bpe/xLYJ70Jwdiv8b0X6+z4OqG4ysL1Z6Mh1jky3vP11jpKhQse5jBE/vk4K4woh
kZUdJufDt5lSPCxr2tqplKJqd/U2xYxmtfP2DnSPT408aZT2IuvAUwL2jxzTAVVq
FBf9Hzp5gjFNK7rx2eoc2mjnxLaSUFRw/QidToltHOvCozWD9OZQ91026hH4c1Rb
xxMIs5ajHetHd9EoQ0XBPffrCAs8UdiSpmYZMlBSSFwylqBTdMUq44DsQBLCl7Nu
o2gf6HaSVWUkLa3CHQnkrq2G8qBq8tHyaBfn7VViN6vurRSHju6si48qSMXgdy0Q
LNi7ldkWSsEKrMNd/owue6nT7WqYZQD0RQ3CyPNX8u6D7G78e8X7LwWS1jagx8Zn
F6VoUV0Lff2vWBTYAQrqCak0T6e83tyFCyBfkXEzonyCsATs7HlSVlcRRFOzXJRc
IVkUHcTo514MrTLgHpXQT9D929gUGxrNjXZMisumQ0fV6CGL/vvYo5LIANFxTbMq
RNp6eN1AIOgd8RkQlePUN4lDQ/dCbZr34Q5QmTvkAqr9kv4zuYFGfytZ+3T6WOoi
FA5G0DZZfK0vnDNolxfHUbAGW06poBCGkfujiusXccbj2d8fY+lYS3bZSOjKZUra
batn6F2yIsLrWRDrJOb//7gDYy7jrsJx4GVreqlg4QObUx+gTRKUIOn/39UYYLbh
hOPrDCwJ5SYgQC4YdgziUraQ1l//tC1pbsJSITBkH/OgHGSnbB9EWI4f983KRKvY
4xjNIv4spYxU+8geBP8C+CSRbBycq8sB3zR4K//H/Bcpx+hjFmRj3tUY2HNozVfL
Sf/ZU3bfIZoZJGqautOmSEi5YmN310Bzb+uc4+BddC24a74qxgCDlFibi1yN1zsC
Irf0/Rb/m0ofqUk8WBCP6BGFjyMmDllh60qYpBIGl/ioOvdVLRMl8wtAMQfCFq9A
zS7O69vtDoDeF6QVKxuGB6TPhCIZVxvHZxNFOFomdgcjbQh8/nlZuCkmbPFZWUV8
G1x9goSdeKw8Z+GmZKB19FD+R0tzFmuDa9XG+2sbllMj35sH7Dx52P7WLskhJ1NS
4YLvch7OnxH6yXJkH83z+4tdkgJ5YIqCk3LrmfJGvTWSKsJagMLzqCjchbC5GVYR
wdAR5jY72aMzww9n7l3gyr/R4zGLr3oY+T7ledALG5VbjkbxkEt1hkHcOBQdP2S3
fFllIo6kCsZ8LgkiIAhSzJO401whk1mCeWcPpRyvtFGdYM6wRlhdtn726QK1ESr+
jZNZSrz/4T3/lsQgFS6NCGFK1e1ilRlhxRizYEEjt7d1272V7YX/H3kLPLvLRs6i
VZiSSN4/2h1SjmFp2/VJF6LvdYTetInbKqvkTSNTahrkee1WiwwPchOCOc43w32Y
OIHl5G7329wIBGVo89FOCeyGFutHfRYdhHdKo8TmXM2LSvk+lui+Psjt7IVba5Vr
9O8521+hnR2/uTG536ptIEFKRu3XK8Li3EbCZ2FMNF7wcfbvXrpppMCUuhE2QwBj
jpwg4qgUWTr9fed5KcVjX34QrIxDLT6vsKJTxlQOampFM7YCkzR7AW8O9IIZKsUK
ne+odQ7lCYJsuVLNGg1gf2EWt5rYtplPGkcVMwOEMhm33AA03q1t2PHr9kwCdhTT
V/npNzysgowhj5+ZuiIZFgtyu1frIRSLlA1GbCdAePGt2I0pZQ38OlDgi4WOeKH0
2QYDnu+RVfPrLTuFKfxZGX2ks2si3EB5GUiQm9z/b8aiqF9HXfL5UaHe5CM/KEGh
jcSggiZ9MRghO63vtQK2M7wkuzcQMecJbQdJvaMbRXVLvpB83OKUD69btoe0Oc67
mA06v9ltJCEQ6TCOTE9BZYzk/kUH0Hgq6ltXcRAGltLKd9giNjQ9WvweJuJC8CpV
ecn65kRhKqAGqDT3sWndpjjzdjvdAGOyiiixMrYynfpSAEkXY7EGUpq0GOAeSvVU
SvsPbRjzNprgS2+vjg9v2tNe8TFFqsZ20rdeAX5nYecB9KQ2vHiPr29zyC6vXNpS
5whXQ6/WXKAsQp2iqvGRD5qO/H05ACF5w4LgOIPJMjM46McH+zVCF8TAHmBNREWC
YQgiVKqJHhouO+G0dmW1HauDIbTORPOI2+04ygqJUOL8DrbGssaFGqk+jo/BeAYM
XXPHzHXuqRoZ6PStkotbw1yW/9H3jewIfj1lzO+ecjxp1v3UbQeNMdCdkBS8+hUN
UUlCFZS05UupIqo8lMNek4CYpRGPVEkPKgjEhWCLjzudSvP1E81PRTGJnHFfaS+8
bFcKlXtzEI38wu3uFYyTRopMlAWfOV74+JBgndzPuqW8RKXARas+F/CTH6ejWXNf
ryYIB2AJyXHwZf3pQD/oTQ0HtIgr+KGr87fTWB5XVxLbMJ9LQf6LXaRLxOwdsGfO
dUD05uapswn21OH/2LpUB2gFvxzv2iOAqT4zYMORREOUqxUZ+J6dWZ0mMxbQUSmK
Ij+theq4Nx2oF4VWEmPDfCl1v30IrQA6uWpAbLPYgPdVrkWYL68gyRDD9TL5osZp
NExCtD96nrOzovQba0TP7jk1nBYqCe7kI6YN/hivvcH3IFJdpYgssluVBc/yq8eo
gAXakVgtzUCEPLJemvVoLNGzKDZ/rHR43kq9osWgcSdsTSrJh2uGgz8/zBt5ULOA
/P0Tw4Xth7eLC37i4mJeLjtzYOSO9HI4FqHEQ7qe+PMcvJqfw8guTmL1g5Ttvtto
n4pgx7AoUdLw/OVLmyl89j9MZVrdH9NtoV7MxJri5Y4pezCMS6WxfqH95OB+IOrs
9WpgepeQ/B8ZgABGOnlx/ZpOPyReWIU15R0m6tOVx7oVtHTNovTd/H1Ei25DUr+d
9jkpzoNL7odlErwQzWWZNExtUuvVN9X+8Z7Q2o5XtzgaMFlq+Nyt0rqrlPoGn66g
ByOCcAzWrMkXPmrn+b37w1iuUxaaWsQvtIgqwFPA3SZ4Hc3KqbF99uMLYWupqLfm
Rdwyxe+SIijrOwlOOqu4pMrOVz82SA/IIpCJyeJ+ndWgpualQMGrIJs3fmzBa33X
yBAzUc1bGQUaLe2IJXvVtJgbgZFFDqBjRIW8xj4uJjlkwbIoYvvzEztL5DPpipIZ
Mw927r7btqFmmISodf6QECnbQo2/ohyZuuCE3rEXpbbSWSLDDdqGld5xBlWpv096
Fg2tnFBhtytdFCMk8w2N3QgmA61cnGzHqVA5u20aZvSdQ/XhodG9brKQnCA0Hylc
fGz0vQ2LRrJiVpcHdJyA2IqkrcfkyDd2QB6+gPnscMlY4SFFGSOrj43HuO8oTocj
uOMhePNItLaO9hGHidgF79fSgo9HyOKJ2ULtiQOYtQonuWYi3PPN4w1K3n7xiTXw
GZ50NyZ7f+SJUsIluFK6WZkfQeMthYVTI/TUdJuTsqmEWG2yw4daQRfINWT3thaP
u7H9BZka/EpChT2KZIUIL/XDIp+P/V48ITBaQrDPi3ZWbdYR+hdar6OFjfJOO/0w
hpik84sFCtrFx5hWmMRT6WaxxcbmzlC63Tv6AxtrDXYI+hjpoh2b+W1naMRUfPYs
MhXsheAbuUaemarKzSJSvb8pZmOJi8cmOvagTUHuCwTuoCwvDfxH+MaJ7fQ876W5
FGIp16ISK0ZHP4RlJd5C/mkmAnAvY0qoxLL0HUgf1Ppj9sMw3Ppgww1VjbC0RTfx
+yqHZDwZHVApECpRzpzrz61fzWExxSrc3IcCj/I7JOXo4EfLVTktN+jzUlW0gktX
ZicqSR4YNy8O1DsMJGYNyu2sc7uvrCbZLqM9zoiSqVoehAFTkJahQBuFcHuIvZWV
aIztUnEAP/+Oa5PxzxepXxS7NYjwZNGwYXjCE4MvomXlwjDV/H9vrIDbsMBdC80l
b76W/8LeI8TRCKDKxA+ibzYrmjcYegB5AOy3xmxbxIFVS+dl7ShJa5/exXPM0Xko
QXi1sTb6fNqpH9YkR1wOz4/J/ikvGguBA5v48q3ILqTY3pNK19ZNeHU5vKyf5bRd
bJRcqCNlAP8dNlyziyvOZDI+18wiTPRVby6ekELU5JsBNuvqHpxxTmGG7pBUVnFW
aiYuKGawV4SNUoCJQtv7h25QyTCsoXgetbOXhTo9SM/ryaNC2kSeR/13MiTH23CX
U9xJBumap6dTduLGJnDyoSGupf64KyO61z4dMgofevlgudl+KhC2A/91JGgtgfWe
6XbKH2RotkZWZWqsV4p9Jqyc0BGu+NvqEeJp3DcZxQYYI6Q9HdAUoec/j/N37dZz
P38l47uFfIAWvMYWRGOQkfJu2IWtAQxYd3222F/etmECEaWBfoWSF51kOV27UxDs
nb2C+qClxupivuh3IaM3QMoYVOPOvRRA4LsDbyz32saaE67v0fSjhstFTDT5qEbf
4jhKoNxnYwvCoLmEM1n+538zbyv/rrgEwsa4nLPKGLl5a/VckAcgXKvCsG1T/1xM
G5hx//WF4czuDUMYa6axALYmDt2eQ6WQ2zeiW4YiR7y5U1fK9Pmd/+B0FuXgKBwk
jjI1JmfsLQfuOVjwRZbdSczBlz1hr/munIUmsQ8DtFPFRXAWWeH1Ixkw3QHVJRax
5KKtrRYn4mOl53xHmZSBu2VE9WD7rAdYZ4xIzfuq/nxODEgGfsCBiDdPQ5cFetkL
qgRFcxdjDhuq9eX6thiVqyI86odu9mXH4B60PTj9jI/6hFkAwnTwIRMYnGdaGdqR
Bcm0YFEt3gXWiUtFygpd0qJuEzg/GGP4vKp8l9nhb2SOzYj8t7I5mzS8ZdP/8PYO
DbA+ojNkUGZDDLAWMrfHFax84UkbShGw5rndTlZNiKlevQNIEEVkLJOwFU4nJITw
wdlnUvfff/8qJrIjagTC68u/8kvtqeRpUn6JKs1RP4vyvp0uE4T9eF1qpEakBJwW
wiyUkirn8Tj0s89ySUbd9kJV0945SDyF3/a0k7qePQfVYSmtI4zXU2H41Sz5RK67
f1IZy9q42tQh0JTuAVfar5HdYIeU+Ot6hPRg4ZwXNw1L0dVJDSyT01ELuq2FSWqU
4XDXP710yjNLCXaqL1wUk5Bu0sthV8p3tI9kAl1kB3b+MDgF5PcnTLhwTcOWG+62
cBnD0ndIfTxz2s93293G5Zfi6N9Df9jcsE+OfX6YBpAbr4Mpk8M2babmKb5AUK+a
tUSycNej05rvBfBRb6IwaZkBffnh7hkJocGU6kcF/5beBGXr2shJErXLmoJJv5l0
Ubh95pWCzSJ/RtTrvycMIuvnni3irEvhW7MCyP/+KRqjm9uaWXR8doyIrq9i26+a
xcDLAePk+oBogR/SG/JoNY9Ew2uM+4G5h+bCngIWGz9suz5aIouGhX77ZXmpimAW
P+MwKG35faJH8zKG5kl+f7zSPqwKDISUh47wYRSg5Ye+kAOIEpTUN5mkM8UD/rlu
Kw5CdTi5RlmAtlfRLPnog74W+m023aVIejir/13RsTEkW1cOhR5pGCB/zsWFsDPZ
apKXOgYOVmeI6flN4cThzQG0rdZBnnIoxaisdquZ6y0PGt+6ahpZ34qSckKE8F4o
f6VH2h8xr2/Dz6tdYGgqyvYD5T7+fCgAj95UQSfoei9zBDXyHXocISNmtRULmziy
ye4hk7eMzGc49nHy0AkfSuxEImKuO5dC5HLTXneOZLfZ1/CztYph4DBPC4JbLHNG
VspGx0yX59H8pKNTPdMSk1q92pJnxtcSyepHiKgTtRihP37j/erJ4JvROLq3jfMG
FFT5OZ2Hf6OQUYdypfVxwnI4YQNAIXqCD5yaUeLvG1UqO92KSNYosag2wqoYIbVC
k7p6E7CkZHZffQ4gtZC/VZQ976YdSEz0hQYxzAUWAeD9/+oRjr5hAt+4R8P5X/DC
b+djTstKDSw+Gbr4XCnB+kZQJWxVDccNOHtvu8NhArG9fd5L+74RBqZ4RPxiV9Nn
a8+VW45UNVVhtfTzTi030/eroE7HIsJ1D4IMPbeMJso95tMmJs+SSUugfFjZZlGv
rKbHNXpo8SW/CybsCYmias4mDo0M7Sr8r+v9JH97TSlql/pfbtWerVbWAd+nOqxW
2cwVfii00rBEThHAjcTsTD083XFNJDHgm/J+NTUfc3EkUFnuS9ckCkrxdo6/0gqK
VcwiRA54SsJr+IU7QetcqxCq4NKxP5PvMawyk8kMsCSYc6ZBKjQxd4gds1aRkHx4
CblhasH7Zwa5DlN0L7nTmx3HQvnanC6u60GhD5ZtcfHSUSkgU7VM3GgubyIKGfFi
17h1rUBXY+B03txyU6/WBuW829GIB5dX+ksJWfWvfLV9yNj2MpeDMLP80OduOOrm
bJ2UqyS55v5FulnG5tqK/CzFxPBFGQHa1b+JcFbG4lgnIv/ALqCVSagjSjzX2z/9
Lw2EVEun7j5C1eF0st54ON6+ZLNW8DikUoVZZarowiBTFTlDdiY3PX9fdS+kNVgl
0MY6QvyrzK4GxW4ot5bd2IvoR4yCgKqDgUmbuMHWBqSWSbgFpQxsNC1gJMc5V1tk
D+DEaAKSI1SQnoMDoi3DpQjLXJM1PHVZBHyQ1zf0rrNOlo6+xHu+++5ld2/qjdQI
acFGNRF9gtSsLpdEa3ShQDvqhnnU4VKTWlDJed6gBm6Ocpz7kX78AExw8b2YCCAT
2CLmujxBMD9s5eN3CDNiUSjZ/HoEfKOIRHrKomNc+u59HS7Nt1pmrcnLvrN8I9Ve
GSBs4nmveshAcL03nxgORPktKe1vF3D3ivn6kUl8w1OJIaOVxsv5nZe3/fVoIc4C
pcWn2QXCPdlG39ihoNkbxowDDaaHctBmzDbkFTjQVPIO4KHprjgt1cRLxPkCsfRx
wcWJM4jLPyqVi7i3ZMTO1RBJLgFmHvau8/IksykCoTa0jNh1XmFk0+OejPIDun2n
hVzafCGAG6p21nf5retS7vbWRjP3n7NkjTeQuLPmQAO5//4RjX8AioL7wUz5rO3d
yZJFrl3LWN/hE2DpyqzKXO5x16eH2PXTysuE1ldpusWof6WksTEQNcW1oZuv44iZ
LzQT6pYEccJ09LoDKUosp27m+9aY/6lSsqB2zglTiSxlrw82THCcIR8lXKuvmhMA
BlZz6rYv+qmipFRcAbxFvNFfFsnp/AU6gdrDUmw3b+MLoFhU8Xb7+Bs0aE/jqtD6
ikdSC6iiQc6BEmTYuq/JC4Fo6gedL4qt9UwHm1ilVJ5rAr5zX2nt6eujgWKI3I+I
5xt0Awm7WDEmUp9ZyIvUKO2rgg0uZnycvzNsHx5kN58sBbWAlQIbdianYW06Y+gd
aNXwbjdSw8G5y+720UQAVwofAxKO9Ky/A44RE9Zt6kuhl+4AR7MbNCcoiQz/dZEf
/VC1EkUHhAaQ/iBeZZYaytN4o5w9BZqI3IIFLU0LC8DIagRtjVZqti9DGceMzcBK
4r3zOIegg0wIN/ys8ynW3ThAhGu0aEydYyLgKwwtDndxNXk255VHtyUK7RAZ1vHK
YwqkB+IpuAOsWTSAJQ1kfLl6BiZKXQ4so2E0QTyWXWApvrscK43WoSryPDOwbd7a
vRop0IvlKqwWZTKHq0McLWmt7xA1JC1crvWrrlsOgxXvUVq1eBojk+SwEjhz57hm
iY81xhMH7DWSUCfOp4kKjqCkxJrAFaLLyikVNzPY1tuvUfTuXpZy1oX2dbC7NIct
yd8hYUa6Jare7dvIVuwT/04TnBKiZR9hk15RynxXbBJWtB0HDFG3/sUIrGauLx5H
VxxFPUmJsHI1gRLxoS6e6EN+sGNg1+5dB33mtZWX/ModWBdwppzUoZhetJJcbcns
J1RnXK1Suv8c2RbHQCLk+wQ8thU4OEBMi65MvCkR5FFbUY7XNn3WXr5KUvz4Z22U
0+Wf6pSNuFLvfyvCIu2+SxlUIJMqWhqQA3fTtNO/NZsJgJ6fX+ZfVk0h3eks/Ibl
LdrRNhEmbvIxN2E1VlHH+qbzLLMtsxJfvd4ympHEwC7cniAfvVN4BhFTftMXXD5i
tySqqhdSVKGa8kTXsXVlRGQ8Xaatt82vS1gfi/WAul/04oR6sN3Q3wYQ3Q/F5VPi
b13bWsvXZpkitFGEFOIqMJDes32wbtKf6Lbksjdi98u9xRhbsSCpe4COtFJN5Kqp
ml7OForlGt+Gwia0IWCq+b38KzlrA4z73Pbm5xHhSGPz7y+gbnFtdM7oYGfvQjZ7
zRYGUxoWNA+tAO0kvA+Z2sQdTX8UhwJZm4ACXly+OdSNAFUgO3pXJV4bxKVGnjL0
wipzX0RPRRUhLLcucl/MtQ2fwMNLoImyD744h4YbXB6fbAjTc2W4g8+biuU3ZxgB
yAFM8lJLDO0tp1Wu64JZlBpeQiQMTkYbLf+H7IzFUISW2UQ7a3KT55bsC2QS+mPe
wgAKhlSk0sGLWVbzxf5tCdIRMHnpPF5XgPrXUUdXuHbwQ53bB1o8SSVxla6QE+P2
Urizu/8sH2NjnltOyVMZ12JKNMybVzXlU2ifdSP8RU00uANklAfsVBkiVNj/YdQS
8okNaRrM89KmKuG8o+76Hb8nJmogC3cGx7nbcw2gRYkAnckD2V4+HVbNT6A+rRXk
MpXTeEma2JK6Z4DuN+qQ8Px66cIr/qbkFWKvLxdw9+s+C0hddqi1MO0CzXW7C9wP
C8kU4dU/lGkBepIGzbpxEdth70/A+CWYk9kgofs2SSqsJ17Hu9TR9POFNbzRcTGh
6DMX1mITzsbw2ro/qTuqptQV2VbAwWZ3NviX1Zz+jQczqhKU3ufc67v96PBE3Mrr
wdK+HyO3j17r0tnslKMRop7h0nUdQndHY1pjVnQsz8Pe36pFCM44A2FY9MeAxdtP
F3HF5n1ssjU4eEPAEwelxxINxRDq45SynNfQl1aBnUxRpXllkerN2Wf6/TAb1lmq
NefUq+6TTvtejGWCkeFAiJiZYSSTsA8u/srlvBm6YAqb4nSQTsMG6mC/48Rc7aTw
t67X5ef4/9C1XGu0KLKKt+/RzbVYK0P7AQnm0yHQdLynumylG2/cFb4HByvd9oI6
x/L4NpXC+EfSEdiNepd4ro10QaCdeI3mb4erT88HzD/Khw2mC0SThIgLNWTkM+fd
9XuOL0KmTe6cW4o6zfqSojB2SxwZY1m98tDyfRUmD96ceCL7i0b58ihSyEft8cUv
QTimdqPkEdo9UOcEt7qMzfn0jzePcXlCefbxdDf+avbHbCYPwJB0U+9p+QJdHUjM
bRTSRQg7bhCX+vVWEhYKM2QJJUTQ652zl8tw7WhCnwkXEiMKEfByCVb1JimGPjwj
RKoOpBsvezbxgYe+VV3b7s+pXB+3465Ja7ZWYJMqmO5cQH3XRpOM4sU3RJr+70kk
5VkdK0hKVp2hyLvf6jKBE4qikOvC3fns3rMMvU2r/sXA5Tlv2UrI1jJhArNluEn3
yAxAueWc0S6GoB1lW65W+dRWTvwp4x3aJSolj9nAX6CMcln+YINulHZoj+RSu0AX
EUB9L4/LrgHEp9hl/HSjc8rcd9D6xPVZp7KSDNoRJ1Lf+LGWOccs9VnXY/6sdqwv
MzvysTCe+ZE9axnq92BCh8vbroZ/Gg8SDwQGlTTrzia0dsEncNOSiLkFPK334xhS
/gVn4piD43pFNoYOx/noywKILzEDWjZx1zjLDVmmWtOJaEMJCIbTymIr3Qt/8dBP
G8pF2VxCFaDjx3/40075rrO7tWeXd0NsUMXfXqJGU+w7whrcp4ZZNUxuZlxPi06M
IC2oHI7SMepngsooBANjysizogPr2VSuGTnCguTLxzNlzOH9+lr5QpFyc201jbEC
RHo+mLotTtU4HYAmrUiWO5zvPPD8/j6IgL1nBLKMctkAc4jaUsK8dSOpHkPWUvDL
Th4eBWpM22YjiHQkfh+ngnBVl/M48IiUy2/W8lxEtNPI5RyoPUZ9SqkNWwMfifYz
FjdfO7+yP3AKrdMd+zOjYwcovWUxs4PWqnO3c/O7STqSM0cUcZX8c9y7aYDnuLAl
RdUb4uRrzQey8YJ5GLyHLQ9xRADQgXPgeyt1XPgHyHd+ZAqdz6y++5d7ZF2zZ7oN
52TcOZ1blI7g5tDbbKVcXxf6Kn+jN0N2UvQucuh7L6kjv3PXrH8wuYAzdkhZq7Sy
noddvpX7OgqAF8+sxAZRYBdj9CpT0L6r5j9yrga93g9Be0ltyONBH6EKEFwYV2MX
b2vsn3LRhbLsyzKksYPI9FjbFcTvOyhf1ih2cxESuB2ZR0rqzbWXmQzDwSnRXQOB
gF6Pvmubs43GaosGwrtoGQqR2fR5BR6qMJ8WKthVOo7HkCEniCQ0sbwgotn0W5nM
MztPngeg9o13K1l9oISKZj00xIMxVZn+Jk+/hzmI3LWv9Whml5W9X1G6Oy0SxNYb
01vxXXG5H8fyvlbV/FBE6eCaZC8Q31dP94xI+cG4rIHSL+yPc3/iiRILm9BWaQaU
7MSGJgmtHgcuEDNmbEImrcsN8jUSnAYNMo2hRq1HUAeDfM0lhgr+bIaO1sxOBPqt
He6Hpg6Di1ZSsOn+akyeAocYxKe8Ur62KPEIEmGNGp7KchGQYuVw/ZFVrJFEtwQ9
jShaWQ6Z1cwlS6zs09yO8/K1yI7Bl4btu0uPzySQz1uBPy7+wgBRf9wVnoiq3f70
2Zs5ZjzlRBDeAkifWmsi8HZidyprscypK5BWGqJ/k3D6GgygQY02M/5RqH8ilSrW
8obP3W2/J0IUQdZbG7KybMJkH+G37tXVgtFOawJwLNUJC+SRLFC3QrjR/hbhgC4V
hpRUvsWebnpmzHt3WCaJWMDR9NcCWgTVBcCSD7xjF+0p7igGI27lzntjkiaWwkKw
Bj1977WeJ5iONLmgwZ9RyPeGRMY/KLzlpAsrkq9qV9MGVzF4mN3gv2/X17Pu4jeb
804UdcEkGRfVO0+KhrAWp3E495zysrcVo7Q9y9lw45OLo9+9ENmuHHUnCJBTGTuH
GnYA+rXJLhsXo+XQSbbTDT7RDMB2RIEdPweFHXnbHgnHg8uws30gH8wPaCIykSYX
xN8lBBc8MQ4WwAh3xEvo2PQl3q1A6CzfTjrWErcoDrphu2yxDejtAyJK6XuSMvRz
f3hRtIfZZY1ynQKhAR5Kw6oJZZyH7P5GIPeyqcGiENjKnUBR+41cZhH/sTW8YIt9
+3c7bjjs9QAdt2B17rkK4fJiNbZvx0kfTuBQfIbnlJhASWE/ON4nCFqjN9kE+Str
cmlEvk2589z1v+iua5K/mWpPTmWaZ8LIV4WrPF01OEOVzsDY8cKiwGmWG51reQVh
IDz++F82n8GjQsfsH9xqkvwIf8JTNR4X9A30gjXD6I/zH6uCD1DNVPjD0AADs0em
Fds8GJHk4Bx4ur7DO7hUK+n+ZHotpZQ+XeR75x0MkUNrlAdu840TdH1Zu4O98lTi
oZasJTl3iOjzfywTFQXAfeY8UBYcrtpNTMcEf1AhLnDprs2b8cMW0InrVq8rmXQt
+hqDV6pxzU95ElgFK2TgFMnMghI97fG0qRbzRPvTzrTKKRnXtADwbZ3KTX9HPe+O
wCpVBN0RjnZJDvxWKHK29wQwzgmz/DvvU8e8ZLd/FXshXRKEvjMt3FYv9KFi+lMT
TiwijDAfgCE7n6xV/zITj9zWfSG4PDAiZK1SCQ6stcPmxqSH1Bq78BheWToHTl6x
kM8PRWlk4zuTm0u9VB4cjFZh2t2GDsMttiVKg217HOHoXwc081iMc8UkPrEgXQ2Y
VJOW4cBekFRHiuYKlUiKdB2GBy7filkjQyKlD2u/n9v2vY3fwrdesDGVjvgM54Ls
7G+1Tv2h4MKym/OCv9KLm2jEzLgjeuluW4Ga4es+4rDVinAQiD1Chnrf3ApfaDxU
b8SWkQwYj3OF94sscoaWjJhh5NiKKts9WWhz79GQMN14Q5MufG0OPw23Y+et5Tlu
nGQM0kP5wopx7FbGauaz1noco6VKrXQf9gi1XpOnDuUi/AZeR+xM8PB9I+mbru/W
e0YKuh2s5X3UeyazTEpRh5kz8VJYihu2Fc98BydZx5BI9HFgcvRuOtJfETUWgsPF
Fn1Tnckcw5ADS8dOOf7tZJ5DuofEsdLIOSMhmO1zjgKBcleHJSCDp+T4+CL236kE
GE+c/moMdvfRybFF7AjEeOUudNfC33T+4ahtw0Cy5cOmAPj+QlNJI+T/nHpnh4yx
1fTAYVq7Zsgp4CJy1USpcMFmYB8mZRFeG6mrOssknKdKdDiKUHhYPGWuue47zawX
VZrCPbTipfChdxxnbwySJOOOm52N2WAxhhsoVT0XwlujT4rSy1f56mEhfIWLkRIG
RgQ4Y+0nRTymt6vEL9BS7nA5Pxs5kSIq4pIYtQ9RsAJro6cOqjpvAjTpYfmB+KYQ
naW6qyMYjuAkl3SLdugJavDN0L2VJ4RlkDT12N9LEEOkankiJ2S7SVYo+dbS9yc0
sfXJYJuFFrV5RSzg8TcyAPAlAFZnvGHgWlU4QvfNpmVs7P6d4oaInAZVRqGQJGOg
/FOvP6BVpqZK2FJTicGypBebMNgWa7f8vAJq4Rd8JndrdUE1HhxnwcGSL201B8VX
1S0dlAv6EPvW2ZdcCWiSoyhvZqEoT+vf0lrp0+OUD6dDqX2mlRdSp13E4NFhmygr
CgyeYHNgNwZDR0aSgCTodN8zwuabaOnZGPweHuJtKc1kcla+BBojerp5oMoxc6P+
Nk7UnbMpHWPjmEdC2422g0rQoRm37KSXIXQzMhmPIV5qlJDWRP4m6fvUM5Po6nEZ
AUIDrWLQgCZyd218HTDto6dK7jBRJN9fAssCW7J3i83s1RgemmlVHMd7bDdD5uJs
TPwVkAEHD/95up9akQZh8JhESAsdeV5XvYQmyH55tGTdX1b6g15hL5hpFGHI8upL
ZExbjk6rmT59SZlouw8sYY3hhHN3DbaAMjjCvpfsaFrlYETU6fxknZWWSvmDymRc
COw/A7BTrW2gv1lzjrMVFrdjGE/zOUtoC3Z1x8HCuYW2O4zGMgt1km9pTdxhslg7
E1No89SXbW4cSOcfhO3wc19PNxXG7p7XFh4KEPnqh0/LJ2/2YaG2gSSZGxS4M1AC
uGCzzDAVUQHPQAzjxzuqO6iS+h0lOXUf+uMIoMNaJOK7tOCTRA8VxDhi3V+CNdwU
aPJ/d1gCOLIzaUkci9LngcImCYQ2H2ZqcSc8x8sLmH2HXZ8jEEBKnHlRT8B9xdVl
jArycrlvjZ9hiTFyjUl8Mpb49jyRHt6If8QK2OSc+nvHahF9BPGnCTk2FAtjXzPU
4z9NMP7AqbwnXEVj5AtFCwTyyW6n8i7YHTr4c8h9uiKOpzRrjZn7m7PWCjM4NA/P
TJrr+etuaGSsbifbKvqeU6a2ocbgGgjmJRoOid0en8rNAvwjdN9BUf1mT15zUxFB
xQjEAq056Fq/IB8h8WZljUZNdesKAgPgM/KFGNomlRD88961WMF4C8C+ruWv6Xwr
rM9qbDQTaBuTufI8WpTMo180yInNpes1emsL4Uy0e6DKWxfiAoAXVgsXzuKCmsS+
73YKWPhuIyNDwNR2C6H5CEchMtm7Og3YzCbFym8lKRERujvrk7eYj6oXyR+3b00D
EyWdVduVEpeWQUDZoSmIgZ8WItZ+eOplLN3ifdnWW+UvVqNpmgBAs9pSOGB6f52V
oHSSRddGgh7DeKGb/Q9/7Q6Z+i5nOphgxkrK6Tz12xHMIEyUN0VaCyJBL8Ohl/Nx
NsOVuAqmXwtz1OUY040H6dF0odn6SdhdhwNsZHZ5IVFQZM7Yaow4yvdhk69J5AKl
HmqzNfvz9Kgzi0YXZg3VDJn4aFxHS40Ut9JmNhKbU+dFLmMkwQn4GdMhzcPRiHr8
4dPLzQgmsSkGDLQLrqepaiuLcFTtns5Hhp0aZCfGhCu3cBIvSjxec0ZTIFYuVWxJ
0LaJGsFINOuV8Vb9lkQ/qbglqW7ziob7N7RcZ4Jr9ORtLjOLqeiy7s1ejXDroZxo
kdXwGkISa7bl+tzKOmIcok47pLHdw6GdKlea3L3LYRHtyyBS40zrWaFQ6zNWlumz
R9eGlAJIzL1jHk8wg2n5trjw4VOmpCiBznOboFULJRhW3dcvnFsTav3wAbFdvqNH
t5eQPXmmGbYAO2cffP6XNYCs0eMUqD6AdSNkVRujvaa1us6P31o+MyEWd62dgYjR
SK5oO1e3GMX+1H7FPv8czwhcwSPlc+7DMDKcnh4Hju5YHINtXrwro1BwQfewS26+
boEZlkbE3qncgGX4uSN8ieS+6S27yu8d/WhtJnxsvjhKke3xqb9d7Hvaad5//ISq
QqFLKnkEoNXi5/JwbsDMDbK6JD+XQQcoaIfC/wLLMsOjzN5DTRTeML+VsI1sJ7q0
CHsPTP0IV8dfuHiparqIvT6LCIuxnynlj21706NcqUS91Nk5YYQUEy39VSJVVtwV
M1D+zT3Om8FnBLSaHMwyOuzxc8uTJX94m3XVzHNlUXPBNkPEFerI0gZfdVyB5pn5
iHlAxbR1e9CupPv51ijEfEX4Qzpt/vaf5ODjAWGLDCzuR1dDR86MQceijjT35RVC
HmfnOKQONsFKJY3/UGibiMnM8TmECbsyafDNA1Ji+li7Vb4xukutxLaE4Qo67mFT
YIr78tJ827R8B7pXqAyMMs4OMbu7bklQZLKMpF7o6IJhdaAm6EpvRPTzMGPR6epQ
NfGtmCrAV0Ji6KxeyBbSx2wWu2KLNplouIB5D0++276X4bwnhxvdkS8/DcmWKEd/
35TV2Q9thJ4HW8hBEG03C8fgLLBo5CuaPCBVqLXJC32Zu2UFlqnoZ8xAZCEzknZq
zszRPnnOOxOo4l5KN6hTminCCIXPYgYSjepel6pgWLDPK65KRJegzVbMV/m/D+Np
cvuidkMHH46LK1/TumaTo1k9jZQ7ZEZORkb8EtAk2nonRagtdEmju2fFqH+z8PVL
UeP72jLM+C0npxiTXx8qpviq3NyVBdRH6vZXi8BqtEoHYAQKYqXlHFLECAuuitdn
ydxFiYpOccZj2tX8IKVylqAPA8aO3bz0DOiXyrqh6kM8nVq2ngkDyAgWYydMybop
px0s8Zflf2V5KDalb0GGyD6wOGEsEtmTV89BaemJqHCcaX7quh+98lxdOf97LfU3
zp0Ka2rndnQw/9v6pfig6KX265Og32R65yhqlBfQiSSCWZBi6jyMW9MkZqLtDReZ
39ptKDc0kIcLLNXlBeuKArytDceWwbakvZ3R1q+nUCwhoy6KSP7XYWD9f+6d748f
xOQ56n9Bvt3157D0AVYq1KRGAiRC2MMTRTeDHut+YiZrmtfx9uOKwR7uoUo+Gcky
pjXbnGxFW2v62nhzGTyh/35aMODDgFu2dbo+Te4Rm7s+3w3M2btMdbe8zofkfon/
5d0OmahERcrj8HSjUEBVmN97JJ2q/mfr0RncVkrTNzvSKQ1HJd5GdP+BFP7mavFs
lfoDYCUD3dsbHxg1PrXlLbZOWBRNvZQ0QjVUxUDpz2qi9FqE0OTD31Jym0ehgPmJ
TyP4mNFuaj+6DbY3X1XQer5bUcwx23RxHXdOywdmbRjNuS7jqHqLm7uqqL1FC9/L
GFUc5MsVd+mq9JJL6raMZQA/44Zu+btZ6gEOentnmpTtYUE2rxWMqQ8i/1SaNWsO
1s2q2AX1SEcmyB0S9nhw37/hm2IPBLT3jMjTw9ZilM6XNWknxY14nQ3bTUantxKo
HrWlCd3x3vlQhtzl+jy1+Gio9gaXA1L4Kl9zQZKRXlVzDHKEwwS0BgFAQzjgOpKg
qbB8rU5cdz0sKONh8wYSY23ocD3cAzOFoI/Lky5DA2GUeZggAsAtJ6sd3eaE3yOz
sbE+hHdLtEmXAVwW2IDspVdo5bHsmAKxemnE5DHjc0RBdNbRxrqZawdhsk1HoXJe
a79MEyzZm6KuN6d54lHEKx3R7ZZ5n0MseT4o/JQCXwDYyNImfwvdk3UH3JPTYi/F
lN88b3oUNpSUSkjdfC63wRV7l42jBdytkqjOCCHJ8xOwjCvrDDNqDdPvebN9q3EA
c07TdBPae7Vf/khF9scrVDXKy8X81fhVFEx8g/xTD6HEJDSF1eleNBB+sYo43ayb
30GGrOYQWAwRiKSduXJDdz5eIlvU3kbUeW9kkLyGUpBQ1k66pJQ1ZX7bkifTHMon
joFPfHLpyQc6A6IpO4DAKQRQnXKwGlWHXZCEA7gSJ0QDWFL1H1GJMz2zKCMYH03e
OdWyXqXs6rl0Xj5KcgUXTTs3fRS3X8LGUFIAWFEKg34D9R16oF856yD9CSQGMudF
DXh/NFpGsS0q6BIrJJnGcDbqeabDbJ6LMkI3JH2HZta8xt1nuiv3ZEwPsEeqql4B
FJfzoOUy1DjUfieKLmwhh56YrLstlAtAzcI8QLO7vVKMl/T86exHdnQtdnU3KUcK
qfWHB9bi9rpRclvvVOfNuWN4FUJ2VUZGMbrHTbTAODOwHHH9egSM7VS1FPi2IS0w
Q3M0tkGi3vGDNWU4cfPErBgNkrvBS2kTeI3SxUaLW4avOF6s8VC1eBCgkqFjivOj
YtUR11DkSsKNjbblbom8ncHrIR/LX4Y2EvK/AR7MPv5+nMpL8J+y/OjQWJWJGi2J
2NjEmtpA79t8RAwtogaTSI/CorBOJ3kmKJ08T+2WDU6jlshW6N/lfr2hxzIZvM99
L3e3d2quVMKBdbF03pXa0FOaZNb3bXEVKV0WpTX1V93NsQc+3tYDkr9Ff7PKbq2w
M+NoW5Lznxsj9CV/p24nyEVwyce7lI7QUXzj4CZ8szy/iEGPvQoN+DGigAla3lEl
4tP2Xv4SCjUiE/KsX4x3wrXqccODfb1My3HCOCFC1bVVq0QprLtUk/wRIrAPovZf
K+MdfnjRkKRkcUXKfeKEyVDH8bl4g4AwaHb6lSaK0DDU3NhLBqF0f5USkHrwIpGr
XSUCsuIMZucpe6m1g0r+wcpONrj4LhrkwkKc1Ezw5DP2X84cqj/yWFUDEpksAGDD
j55wmno7diC/CDTOPn76gv9ogwuYIHDTIdDco6is0TR+nlKahU7I5vF/ryFrp2NA
Q4xwGacQ5BXcta01gndoCkF5mbmTkgSkqGfMqzXDLKS1f22o87fKPJFy1rwUfI//
10xjhoG7I7YVUnGqBVS0WEZvm5+6Y3deVHwKC8mMCP5K29f86/8pmZE1Qnxxoqqu
dTIt+b4kQkRfmx3QInRxV7WdPCXcqLKDVvglQDjCGLHgPudrq7K94AItVBOvRzQ2
XevnpnlPHTcw69PKkjLEuHJLaRvfYPWeRL8rCfcutIcewTOiMty53QvGZGko6++g
wkiOptFOi9TjQFg1/bG5MeCrrtym7VU19D7QYHhhevjZYLAQV25Ah2WVZlGXAq08
kMuvu01ICpHIQCmTC+biqv9avhZtaIjC0LY1T0Ok11361x9V3vmo0DMFKQiETm78
5jO/jwRYZc/G2/SgIntqxBYegIig8Z4Fm4KmcIb+TbiSn1485uBKczVDHYBJPdYZ
T2CNLTE+BAKspb2GDNGhfu+pwLLAA+7bipdatIwo0+djeBp4gp64pGdoTENjrhJ2
LiwHxHoryo4RrdrPTcNgQ1c6CsjNiaW6JFaIfc3uwPIvEj8lSGyrQbg8omrWErvJ
UqJ8A8tJ0BWFWy3RBAS9XWkjg4CSktZIOxTt8SAblk7rj89JD/BpM6i1e04lH7Ij
86dbeMgsQvfOlt3d1AuwTlSCu7oBbo+vLRwco4lt4AO3RnFfQ90oYmDAeohvk3PV
cXDvIkpV1ZjeOVASWbebIYN/CtgY6K9YhP4QmSpN9YvTq7IsFeYxMrK1t0KOZD+B
blYDtVoJpltj0xNw1A0OvhHKgN8d5LNFCxYuIlRXuLqZODPdkzzmIgLqqJeoa2+9
MNXcmI91ybspn+cJVDyGOtEKH2q0/9pl8bn4uOTowMNzZtq7Tad9mBzmbcE8M7Al
eMtV7Rs1WKWqzw+DPJftZYsyV13PlljKxXhxLnIMg35xB8IkUbYZNcaq1buXuS8v
93MVm/w16HhCc0tkhPTzrXWM6PXPwzBQh91Y4/IawszJ/7tITXAsXlzGPfCmMati
PLjj/qlE35oUG5fqEI8anYGwjs59qI9UEbiio3v4y75iJPHRQ/pguc7IPuC+XtDG
ZbURez6JjHtaKHmgkf1xIigt4JpNsYYlR2Gg5OShKHEICrZLbt/4P6AuV6y/Jq4w
rPO9hEt+AcavddJqRBgks2boYwZJudFwQBPu0E4r62kWzeQjt12RYfEwoc7MHoQ8
qW7U81zXef30+hIlHPSasZW6lKopQvUda6GzKXpPuteyT0EyrF5nd4EprohoxT7Q
7xaVSdbMq+AyYkxcQxXYHiqQChU8+1ECfIO5hY4aXlSxHnNaMbvwF10lJox7OBpl
cVMwj1w+FqV6LXrm3w0Gy9qLEX3IAMiBQ/KkzF2WtU/9UlfvVrSPbORWpRyL1YWm
ViCY9BTuMA9haR+8wysbf04mlyZPjjfM+siHIiCtPp8iyqWwVtt+EFGCFEEx0nsJ
g4MLWYprU81oaXggK8Jf2+IxP9ickDal8KXIKd0NMDFTWhVbDGviqed2cdD09Fr7
tKgPz0FkOBpwSh+giZP+mPdbklfsQIx1ZXxPIDgsCZ3MMfSAIPNjgd+7DDfJsHPS
d0HTYecFEyCnw+6/pdkSKTao1yL1FfMioT2EoUEX+jBIIvEWYu4BgaBYH0Jg3Zda
ePzYgHN5ygpwLBMKBLyH7+9izIJPmZDRxkD/vBR5RbGPJhHq2Ur2rWNYrNgwzvh2
Nhdoy+JQQhMM140NMqj7nEsm8cCi0OM/R3fNOgO/6EhXIQVaUrX6CZuYg47gAqFf
xSQzIaO/RZd8ML0jrWSQ775SIBKEvcQL3Nn5PgokWce/FLvnxiJTigChq4nx8cHz
wCKFYIG9ICyPY49tvfjbHKr7QsPY9MDZeR5m8pA1yD2nkKO8iURrohat8wT64YKe
1I2S1j6DXXXCtDFPmSBp2nLYr49yO1K76JCMtmaEzQgcFbgZm03ILnt6WMSJy87n
+jalR9WVOblTv/IUj4Pu8XposWmB2o8TzY7ZLoXKtIYtxqybhJpML/5LgZiZc+is
qUV1GhGui2P8buE1pHosUh0BAHsm9BQ8CyMuiqxrZ1fXsIVHBsiwy4ZlIyo3u/rA
RF+XoNZhSMR4/NI1PmftXiXgTd+ZoXz80FIwoDPj51Fn2NCBLJU1dASM8TA/TtyF
J2/giVXl4H9MXVswYGYtx3Vkz8ij9rzp/6ypLFDDB4fSFywQkOG439nOnXn7zAxM
GgPlrgqrlSufLCte4Zpq1ehKsJNYZh+IXx510Lwaj3vricA81xti4pqzLn3Xt1Io
WVwn5LAwbX6fB5Q/hiWuAe3o0fyX0FhkFSD6qXXOTtmyXL+NZHWSKAmoynJ6AYnd
4Qcp5F8sWxkBFgB5MTz2yXC5vVolHylBZqwvfaaG/JD0bthfzsrIOrafUyJKjFvy
/IkV8ZJnO7OJR+miXm7cR00sqeDA84woRkKYSuIm2yXNs+x4wbqge8YRkuBvWrnk
agyTSxfAO9L8AiWp/I9Qo5elID96fYT4R6cBcl8UqNI/JN9YbUhoEJs8zqk67rW+
l7rao20cRjdwtz7WLs8xfHgSFk1GUiBkK4CoJ4h8D/lUiq4PMRx9LAKScwZB4qG2
arlqsxCgkAsJuNDf31CIO/KCA6Nzo+E4ezbyofYlqNHdDncybpQVtMQdX35mUBug
DBojdRwLzShzdjblNddUgSvfKkWFgURAgI2O7S2h4TMRIExGaWY7drO8ee2JpfEw
OkdGlq+4JK2XzmrE81WdI2LLsICN5+XE7Udg32WbOvmQytrKfY6Yus4SY7/do82c
sz6iuI48hGwasfW6NtGB0FKrL8OPDB/OjRGCIy1F+8A+Gp5nk214rHeMONJ3G9n/
ZEtZGmS3Iqk5s8zD5DpzMn3QtaNBt+h+esuu5RMLS9rHwlq+rFExohPK/CvJzx8v
WOkrCygM3Kh/lfTvjrZ+fswev8xfAB3dt+gVLbibjY74wtjnbgatineB00J5iNtY
J2qZ3NY9sU4EcWnfZOMbJMyJC8bn39K7iONEVCYKaSGcVfLJqRIzZbTrq+OSwjZz
siJ2u3JSzSQT6q6cmzftKTaSKTZjMMP2RV0z3udlWxtODM3WmpXWGlWvqcjP2yfI
DwY/P3OjomddXlxGSft9Zy3/Cg09E6SDzLhvgB9YnbKnQr2njCIOwaQ5kwRMlw4/
jJcB4OXSCMHcaBi0ANL0GpXG+jmxRSEVj/g1J3tJPRM5z6I5kWbfkGjqRDsfolmB
XiMpE/h4hk0Bd9BRJpFGETCOFTgk64sIYtpcM0z/bHEJa/Pc3kxbkdn7fQRsM932
UxCIfSbsjPvWUX8UOKY8qK9dD2jdHjaGOruxmxBX/m3LzpDOHOMbp+qr3fD3nRaZ
3NGJbAybVTVWPUvG0sp9Vf04oM6A+ZGX8yRa3zF6NTrQtn1qh3+N3TjMkjTrZbQO
WVVl2r5cxZJ57mi+bPLRi+BOkDU6ohIxh4RGut+8OnvKgefVQlMteayPTInkv2eQ
jugE4An6WMyCHNAAYztKCps1Iet9kt8ZtZrWuUIrx3LdEzcfwftd0kJLE99vvVcK
VkwQGqesipQF+KJIvgPOHHcE1A1g57RsIP6ejNeu/Hr0mhQLLzz+ONQLTVn2O7mM
g31hYkrKE9bH4cAbjMYECJY/i4ykqZaxU0NnGu5W99WXqU+myms4ZzgVsiAAWTmx
n1jAX9bDjUPRW/VYw9sBxFHtrS8ZVLUlauHbSr/0XrG0DB/0ePcgz5AFcSBXSihT
egSq560NqIAwY9kx+1RXayqZQtp6ZBk2vJIGA805iG7diJiPcQZwOBto94Sat2Aw
X5druZezhQn/OyPqH0PFMVhAoOLFCZ51MqemV7Bjnxvt2J5mMuXgcupWJfC6TbAx
D6wfoKi1jIME/Vn5Pd5iQYFThT0KtRibYybE1/p9L1z2vu8amv0pD8nCBPvh1sdn
vNlYqDJOJRsslLJorkSPlAWSNpQS0M2O5eiwzY+X4D3Dms60hgkwDAZllxx8U3Mj
sJ2gT4qTMYKPToDm257jTGWm93uf4vuLdnSeX6VZeSZTPeRQtIh/pzYU4W5lAZNk
ZBA6iHkl59m26JOggecsIs6Xcb0TVwKrJ1gY00jKh3XR5nS+jtjTStqUfuCyKuNy
/RysAgneY2NwU+GZnLcalH9PPYxXK7BKJ+MMk0ild6uuwUnn3CkRul82ssjhOfB7
9C2u8TaCnIauN/3/TFM1DoVQYNbPjyf1fdhN7+rcorsITLdO+xHSHtyvwMCzgLSy
sXCpBy3eMiBARoK47xQxY6TGUC6g48U6i18qTdkR+zYTGF4utq4S1IXlp4Jm+KNu
kNe5JqqXD6YEgrnhSA6cK6RbiDr6Hb1u0DFi8OdYAbVc9MDW2iz8JyOWAZibMIpj
Dx+umf+TciSZaClEIc7JfAELeMfHjzX445Xi8rnyQ8BmQkxruJB7Nebfn2qBoUQX
ryBopiirQKCgU65kIVyTO0imFa/F8e/tmdnnd62QX8mPxkLX3HdmR67atdZVOmz+
r/gYQd2qH20lNJ0zkd4PzErA1wi9LsJRp+nLE/kWPdb3JdiEs+SNHZT1oyR0QwpW
6QQDZBZ1zgul47UQQH4CwdD78KkByuCbUz4v9eLKCdYDImnwoEj9vS+71Sn87tz0
wR0dM442VzIIVTSD46axnbLENo9bl5fMQMiRD5Sy1HYVd0yFse0g9PksfLYejq5V
1YzSwOk2JcHElKHM5FO0+L3XAe4WEqAE7n0Ah+rvnl596dS6CnQa42BShwb9H3cC
rthyWwBcIJtX1ezf/EDCOoKX3fvuIOfyTi58I1S7btqpWNi3PcbSAsbU9Xxx0FVy
FMazFuyLtgxP0rwsnXV30lWwe4golxBCM5Bf28QKUkTO6GeqBfQDtu5lmtckW5Dw
7BGJ+AqSaumBuP4lhqyqxjizlwjonM/YuF65bYwJlOFomrs/XNFsyrcb4iNO5APF
U5Ju3Ot3VDKeQ5hDHdhF/HUbsZAKmq6St2DVYxc5+OvP3mBswq+68JiMSszxsMQ7
Ia4hzFmmRGC6ZvMv4wbdFDHSFKo9JGsZPNWUmjevBfpaFZh8md4su8mAU0QRKdKf
zPqz7C+OgI4pF80M0lUwSsVLlyjvRwk2+FUAi0LSMasabVRtwZOyZJtGXpfGv9ZG
5aaoFZmFlEAsS0wEfwrrs22P3Sc/fWwmcHKle7iFzGT5LqRipg7EEcth0H37zsnM
96HYPyWV9g7S2tE3xJjOt8f+JiaDFSAsEy/fxgjEJntXOB6lqB6B2FHMOwPEeK0c
Zmjyvnx8N89Lc7qcU9Qj94Hhy6ui9dcmycrIlI8egA2dQ/S8sB+X2HWCzANXl4I5
rY7Z0SPr5NOHLqmQFbg3OhgdswpriWTIlliOP3PTvYvqNd9L8eh+uJZoelxE7ivs
vu2VR9YmPDaPbltmPRFNctoBzmovoHSE7DVGNVBk2iaByIN4/coJte/qjHS6fXHG
CtGcNezFTQJ8CuzSppYXujtoJy9YcUmHMoOQqB0yTuOmV05keJlZsD53udHgMtm+
HMqWhKK4YthGveDVFisSqTZRAHDuQq4jI5nNvqduaLGU9OG2hGABmoqxsgjy+HsM
UdV0X+zW+jHco4fardT1vPt/r8t1J2ewbTFR8Xt+jfITdzGtuh7/ePoF0B8riELf
BF4Zf4wRAnrRJrn5xDD8+vOQ8ez5WXvBCtP5xnM6cAsMXpP1m6DVj7D6SDGLV5Pb
0AvxfU8NLTzv52RsZxfladDdaBmLOF24N5uiD94OZgj+XcSGBY//T4/9342DyN83
5Ajprde7ktc2Igk+s8lcT+PdzRaonVr6f0RiSzlWK4TqAzmpE7rW2hc0EmKVcrFm
icL/O2mwNTuTmpRhX1CrIIKGFOOr+mYkAyOVWWEFNqitGvetbHkP+QoRlfM83/xg
reMZNOwAUB+ia1CWMK6an8gzSKdADodsWcUVHpV8ybn5IpuC1QNDdgIKMwxPUNTz
/SyICjw0V9TSWBWBC0R1gwydS1WgWrFlZBmuf9d992ttHL7RgZNpMNdg1CvS4m/y
B4uoICufo3ukXsDaWBu5Gag7rnOvV45JvN05ZtQ6ovLewfzAFnBd/qn/bvxcXMob
mGfhJXTdVIYXlEZ6BZAfX7mV2Fqe5Eyh4jNnNrD8adU7k4cSAgUUIyNRyF8UcoKP
G0RdTvwgdCblGP95Ee+grDNBPAa60PvdMc7Vv48ce3CwGd8psPrqHyz40C9MOImI
lwo/wMhUc3z81COu0Wkz6cWvM+fFKI0TfLoYISLbfu0zigLhf8Zr1Ga08rgTeG8D
m4ZY0lnsxYzIYT79KzjQbcaFL2pYwrRUSTPY4ts04e5l1e2GOLm99nBcXr2bA9ya
3NznEfqvUUs8DTlE12TMhLyg2ekvbl0v71Ry4jOKon7IjE4pvXj9XCxkBl83rGCd
xeXkpoFSBtKHMZa/zljO9Z2PWa8wDsl5u92faQ08eMtI5EjqaSipYAC1obHHDERo
jZ9nKakNacGXmuEJcJOY7sduzf2dJphrEmSc6Wwo6FvQ+o7wk8gw0Y/CkEbZNLy6
YYs11qewv+vO4YPjEjjHVX6h0tdMAvKs1Gn2Qt03u+mHN93derwF3fdifNqLwe6j
haeb2ab6UCuSt6QmL2S6aRzON+kMQnnMPeDzetYroxqPBdQ/FUUtfgdMV/rLfI15
yDjmtXfnUFnUUHEhUnSgbYkXtVNQzZFI0vqd41ErAISLIzJEqIs/UYNRHaKHyme5
HdRgHUDj8eT66rKZgJH17lRyp/JW91a9tPQVPlciHAfo0y6wK6Xc3Y8CQNk96d9t
pNG6uars76G5ikOS2GIH2HXLDczd4VI0dhA5mcchNwVFFAYLVMVUwPC3Wm0yLqAr
vsftQXSmdO3c7l17USoINKTURfvetj7LJisGwOTuhOdRs8+7heWKS2g6xfOtR+pX
e48W/k4Fc1iebZh82OcMAEwGMUCUZZdLNtbcZM2BHEmRjpH9EbCz26F0lFG3bJC9
eyFtPgzt9nhUbYqIV5mHcbGpKPhfjsTdSA5XJPTCyG1xqQJFkvnrNPANVSLfOQBg
mRJcPgUXco09cqkgteud64qfXuS3ufiJYWsybdSQ4zcVveWdo4u0YCr8ejMhUzMc
PfCmxDhJUZUWW9UQe8VV/KxM7CepPbNoQ+Kpl72SjQ+rLT0YSlYUzUg+8mCd9lCt
C8qah1qUDbvaCGPN98zmIRmdevRJBzSKPKfUZBwjV5OJe23DaaxcI/FQI+rG626g
tIReEssOCdc8AiZgzLCyuDcvkuUq09OiABpNFOD7Y/FTui4j15UvEZl5swLNAmBW
mzFzW2Zk0M4gFfIu2QVrsTpf32G6TzkicPNma90UqZEdmYqio5XqeCZ1SRNj7028
MAybTvk9xV1xSkOsctZdhmW5f0CQbQQNbQsUkVAOAYWWUDGqJqjuIH2rGaVf1/BE
VhSIkvaBxmdswXbeIuGtNX2xmexX7GQtobDCxioy9RgP9f87O04X1IG0aufD5i4z
xT/jvg/OkUZljB5nFE0jJnSMejdvmejG9EqBeasoSk4UtgF0R6RTpCb0KqTT8SOG
KR+3ceWYBvSEZPjlmkxSQ2M/d7+MdIhJbsqK2Pgnbisb0yF3Pw8dGZoBm2Gkkjeb
AAT4s04TFPQKQTXZ2FH5WXCseJKjh9lI/gHhvuzFSw95fBfof9obIHRTo5bnfu09
Dvscv8r7fX7DRGt1RT1XZr8KTXs3L0dBdmB8aHnkb6vDp2/6lM6OfFUqXLoemlfz
yM2z/qEb5prNC42tO3qafV3E5d4U0Jw0bz7+ehR7s69x60ESW7f/XakKML92P/D0
l3JGtvJiMRQoD0oFZCnKxE9uU7QKpXfuwuNiJod3afQSn22dJVV5M7+LCuZN0/x2
f5QLpKym7dbYHn6LxQDH5yttWLopHtBj7+Hzbj+LF6H+qBED0CpOo+LycC500wPf
0jd6iKt9uMei9sRC9gfxuJ3MOV0nHbPj02wPvF3DQ3HuCqHLB109h72UyVj9RSvP
KHqcmXtL/vd2jjhlf7RUoGnpXeftE+0HjhE7DJZE5vGKkJqzFB1c5WVDRXg9zBOq
+gt/uAMfTm/79eMiGZaXcyEEiwSt6+ew3s7iCoak9nLOFit8EPglcOrGUpifU1tZ
onFNL/jRhuUzOKTr1NEb6ISxG8354QBosw5eu0ZuWKU1YhqFJowMkQreMYeJo9wq
PA9HYWdez60kO+u8nSWJXGOjkCxt9nNXZDxTr2EdPhp0bz9izJYDT099CO+PEPrn
N5wT3OBJK5wfvirzFB3bHUeYhSEevDqC58Z08RacSJ30W+QxC5VwVK1K7Mzlnsde
SAlFPHaNfwSRCG2buvqSLANom2M+zC3bEiLqWc+Ra9nS/m0t+3mF0lUGyhaT90ou
rWcmuUTNV04va+WKoDDtEYoSnoQAduY7FqSRPfT3lImZaEui25XtGvdf0fruFcvv
po4F0RZJ+4czC4HIHrfMSfK01vgT/xxGaBTzknVCFht1zDGBGB6nd7CpqxMwA9Fh
bdeh/ZRnu+oZDSxadr1Wg5OYufJsWSabAvbZRblpRej96LDHgw5KlFU5qS3BeDtL
agB2Uw1Z/wn3jo29caabOQ6eCi99rpEtIM8IS5gADK/Nik0TEJr4d1agCyraXg1T
7knAIR1R91QIwYE4j6et8/HQOECgjcT4WNrhiXyaXOQT4AJ4deUrsEGFcKPNqx92
Uf8Z3nf6rOc0llkeKBKpob8SNCn3miRPFnNYCyIVbrZy91wyEtmkZJ0gLUuPWZFH
hIvUt6aVSaHPKP8KVGIhvKD4KYMDAQK1IeyTpbhe+uA02btuFLjy0ZpOwPhaQ25p
HMZWD6LGBvf+ASqnid4qUxGztO9fktwuVqbBYytsvSSjD5awmT0VFnF/l8IQB1n0
Zt9PbzFr3U0Y4eFosDfI+o/ViYqzrVJo6FSyBE7m2bFRh0q5v7dTYh7qsoh/iU1G
w9KlTr0BxuS2ICHMeUcGFDwD2v5jX/FrflYkJkQUGv8xcuLHH7dj0L/SRwc1PMik
8VfACv4SZvLDT7sX+jaDqm6KnwJjs7fA7hIA1Lbh0GTDs6lJlxKqN1tzVF0mueUr
BeXUlVeSNxkx2443EwhlZzc8ZWedBtpUTQaueqbjTSBK/QCaojmg1prbykVDcIIL
TNiEGtJTiIEeEOOFLo3kon1DhPaZvJem9G/pyNIVUa7op3iXH4ToVmwxdLW8ln/E
45WmHuiCcy63aRfDizAPQZkDsIOegkp4N3bqsg+qozuO+jYt/r75zWGlITA6YCFi
F4FtFHgudvPjtRI8Bm4dAxoUTIBRraLfhs/OQXzzdjM1cOfaJPFe815Uh7UN27aj
ir6UIXGlBZ80KBDgdhSOPpVjx9N77Wd7YoAi2d5paVHYgdEXnJ7GRvBtDLUvvXPq
2QpteN5/5lYrSire4Yv+gVHNvff2vkLXZEa+JzXA7mCVoZq0vF4R8wGqKW87snZa
9PoTzCtSNP9DDQIGPVQ4YAvZbmGACteKXXOlIcrlkd7rYCkrxZPh42cKG0+UZDJF
aUYxRj0SPm6rP9F8v6yBfxUcasuQnVivB6DVvaVRySWuqfUELrtUYUntON3gLEkz
DK5dhwy6XE6EoYHi7JTzpNxR+utlA8P+x2uMqllkFKiXZ+8VHFc5NyCnMm0diiwd
+2aA/P1PK+ROzCsnqd4t6JEJFw+gEOo99LV5x8Mvh6/A+j8grd8iSsI53aVwjefk
HNSM/ozKc2zkipPoohk1Vrgx08OCZ5WXmmXTXihKAyZHLhSD38PIBcT116ybn39A
PSq+TSQgkLnBi9YtcmOEZl9ucujkXouVCCVM/VtoiT+JD4gg407JMHdTXRxPeQB+
U7+prIpB7kYS+6XJOtW3TbjKvL0jo9/qDrzLKGxadgodQ0tZMZwBCeaax6xoie/4
vJp0wP1UgRxiMaYNLbFXY6vAfhM3OzIBHYAb3a1ytgnxwgBbWnwC87WGPBOZzQZz
9JWjTf/nq7LwhzVsZLW3cwz1eDJvxWmW6MwBz+cFvbR/1kutDO3tQFQw7aR8NZmP
d55krS+l0lNyraXqaVaC1CHMGOK7IqQ2UOaDgu4jL+fs2o094jOgBYjqAa8i/mc+
RbV+o9hhPugA78ynX60u4gtxojD7Vv/T+tI1zZ+rlR0soRtXOLA/PChFhBuHHW/Z
RA/FUlXqXJ0rXMFN0owp2bZOiwYjhg/3620oXMyNxY2G2mMh5uCUqx6/q3Kowd8a
KO74x8wajzUrpX/oc+qY/TlzMsVO2sB6uq1P8H+LeCjaVWuFzUilFgV5dFqj45PF
X3n4UXEr/XLHe7vMElQzMx1fETSLFZ5gfgvZk+zURodoYQptarL+Q+LUT+4JyXr9
qnnlnJUwn1EwRImmWJ6r8qyfQlL3JkHl2Jc6wFGM+Fl504ffMJ62VCp4JrJsbAU8
yJ2uablJm/Y6+D86UX6T8U7mpiIyYdDogdStNM4cxTETDxNW88tSHpwbYn2/I0Qw
0sS2E3LkwyP0kWSU9mcdBF7UDDXYgavQZr1pl52Kc2yhzJ9e2O/MbxoTNJxsJFmx
PkQmbuC4bpBPSkhJnphtpz31xHyX2Lak/+GjjSyjG/x/7GiklG5srmNV9PgwSUHT
f8Ou3OQpV6ZB2vk8PQIFhJvsaNtv3TAhDUVr0o5XwxLe+cLE89QSW7e4P9/AOS1M
pcyp/cG/Xxkwjo5dqJmvjfrQg+2F3ex3cTCeRJ2Hi/YlN/NAOnFcdISGN34jqsKm
LMVHKqW0EKu9mv+wrBTx/KhUCdVaxQ7M9AO/XbftUkWmJSMZ58QEK58PrWp28yni
1ZalCgt3UA7gBuBA/5sLT3DcwMHiicfhr47RmrSxwH5dVYcYyEV/G90dX2BkUrq5
9bq63r0tyehDB3x33nlw58H+rTJ3lwv6WvyGmdp6BQm2sR2byQfy4Ugo9fAmB3JE
+typ9l1WMQ+rKRSRFnMJhlrWTjAuDPRdZESupKY9HUOt66eLld2lueGi9dsASTCP
Ed4rjV5ws+M/XI2qBWgT6nSIwS3aDga+ItBZ2OASPmeV7VkEhPspoKx4TzLEpLJy
9VkDzlVCfwM9+9P9sRP5jJIzYVpGjHtzkbX2bzjzaCchggxhYcNVUS9OBj1cwX/f
qZgrauks5s3wCFJGJ398oD2SoJwtmAepExpZoodbrPwuioZpYHxSD9esOQSNdIU5
3yP9wAmfJr0VLJ4ljoAeVHFKKg10pahylAp7HsJHoRcZ1SFfYBp8stEeLRJYOjHq
d76NB2kGrmaMPU3hm+Vhub27muH+ByIncj4et+duc6vQU9tF3hlPyhcjYVuZMb/h
9j6zvsekkDjdrbCVnFWCamumR1K32qM6J26hmsSRTs7np1bOZRTGNLiba9siURUM
e70nYwcTSbCJR1vv2BJ6ifK3Oh/wYa+rf+i2yT8M7oztJUFU/2WAKTTg28x/OiUA
cW2QZlXrxx5s3dYKdGKH9dEiP9xOI7+2TmSuO9D2itPZcaZFlLbspxQT0iYZdJkE
93NIB4PWFHJhUiovjGu1vwp1R/ja9r2ud+tr4O9c/heq6Pmi7e3WUJCF4F63wPuD
IMpDQgi8U2nCibr/dDijH6WNJxrdCjwbZzWIXj/yd0ikdcXQy39sTimOTl7VeAg8
RPocAK9STW9mu5h1r2YM2oBgONgvfBAk2c/WTftmVFnAO6MtSZ+b9rOHuOeLeQYO
EKir3hF4LDd6NZxPOTTpfRgXUDJ3d9vDxv+ekrAXOhWBb1jV/JCohOC3k9FzIVBE
WnYBTYoBLbXFMsTHElzzDkRKeNPBe5xekKdmLIQoqM0LRFkNAfqcaHjWkL2LJ2yS
n7xbtZV+R9khhfX/mWDyLlVechvLDNc5wg/7QcySVG2HWDN4yMWYi9J5R/vFETK/
QfBZNMgyoWp78EbKyP39EWFRVV6jugw98hA2jkgNvb55J22leL9qbMlbztSmsSJu
dv/TBpIBqWLdQjqqi/m6siR+pgKZH2IiiftYAWxQ03xvkJqQdKvWfwhsoaaUx6Up
PIrDi1Os764EHKYX/DfnPffRHH3I2t4rpUIai6VGBKo9n5RTmstPeGwrFrIwceEn
rVNHPFw2uZMBl1De4JpISdD+yRMkGigiNtOspsFDBWVYhLKH1LYvxce9LcBzBpzb
Vq1SbSJMdXCnDnS8K5wJURK6jrb6OmPXaok0pG/f5VW2wLXh5u27NG4oed/NwZry
jQT7jXVxEJS6vOK8nfgZY1p2dSKnwi7m4jpNEavVvpl1unfUuWvhATZeudkFGK5d
kxdUsn3T2BtZBiMpdjeAENhwO63t8oXQOLrSsHq1HXZVUViABsfCTUTDwhH/VNqp
DbJqDsrLRxgGOMAng8QNynydFbrp6tDATdagJuuN/OOocKYwTv+/LVVoP83Q8Ahk
GIqkHZ91jF7I5wfIHtKPsjLd6NIV8VfAXXbkz5bcmpy95f9R/nlnY8TIHx4/DQ70
RL9vxCwWQnPXTp4C91L6Ku1LXqaDWi3qshnzrK+m9EN8YxUc90C2B47nQkk+BFju
YDcVu/ADcPtEY+3F+2TXQKGa3Wyi32mOZLgCJLtS3wBVBltFkVGGWDvnjaG0V1gu
3buI5kNFowmudm1D7hSoK180wkoqPmZwdKNUVeE7jYcdZZgC8QiuFLW2z2ox3s0j
iS+JggEVr4wTOFjfMICUiEnsfI3k0KMo7WF/n7JYsExxUTff5E2EW5DOzp2yfcyR
5njyIN23O0kuNA59LVofAExLXhqCSvSDnw9g+mAN2PYFCqoag7ejKuITtN2dmM7k
59d1hBJpIJnF91jXWBzszt5+c95gavrPGCHDxl7M1uwHBG8xwewWlZTkQK7UW15J
SXlXXdLOQZePFwtyNe0uwwbN2njjKcWmzX+YKIBMvhTAjleXg+7SWSHj0ur7I7Zh
k2LnNyh0EWFqYQ9QqbOTAaM993h6PRq/6er/1oLckOlRAn2xJjY+GUKhuPLP4f8a
lJje9P/kEkrI5s18RhZhbrowbWZVnVPTFKSsGmWilKOVXOAlFk/N9hSGIdeu7fFN
ioVahiHAdC7NlblIChR0UE7QQHf2LXXZbVqZ3IAAt775YVzoN36UWWTohTw5CDhG
bD2M+XOPUn7gf7lFX2qYmHULB/mOB65VakGXKazS0heSN1X/2QcH2CauWMY/KKWB
Mmn/dCSNZU6Mow182JRpD8yA+yj0Ekeq3Q8qBBVjL3oqA27vCDozP67i9VuWOr0w
4bokZrNjA63AXTN/5gFT08UqMYw2mntBtUeGrxk5o3jbcycboqGeSGH/YYZ/w3tP
8BPHj+HMMyGRxrbPopnwpDBbe8N+AyzxNVNGllz+3hKgi+gVGfbO9EgwhAoP3GnH
dfdlLAVkoMfTx+v37u3m80dEEOgw4DqPGwullKW5jenDPxrsjxTyOOOTwGPNw7XU
59kQm3hg7u7CN2/229/DKctotqJlO91ZKuW5ZWa18dEyLHiXQVHHdZQiczMqVXYa
oypn4jRY//DuoTgxVYcSfm1gjQcrstMloPJHnQtJ056b4zsw4BZRFEv6Q3epcm0w
4eAIm1qUAx3LzWzXCatOIQbXjt/q+1A4D63HuQHTTTitOi7wGfpylfcXMT77qgW1
Bw6SnHAkHNxV5p+r8kkEbn6PfSEeU2V2MlrRGbpsIv6waH7HTyCMayR5fmBO+M/G
uv6P8Bo/bbqKu7d9O+mxecqoklrLfOpJA0sbu+oKunQf2PyDs+KAPtgKXY0Dqfja
vJe3XQ5jsPMcx7jmHIN65Cq5HJk0Ui+l8luSAjRjJXyfOo1i7nZvaz48JqYQxreG
IV/DLos0iNf66JLvFU6NryClaSf05nZWU76qiHOh2HgP1TgBvC6OMdWU9FlyxUiI
n68pNoCBqMzUsesvklW8ps/Mkf/fEVMc9iC5XcUkMUi0rqqoY86q/8xjzqHFwNjr
zuKRra+D4ZDv0Qe1h1bqU0olld2CAA/8KyPmC0mtn6YPGfjzhk06zj/yr2vT0pHK
yQuS6JGVypJD6lgmCG96dBaQ93hLAfq5jIlSzMK4zQDP7ObCSCEZ9ildVE1X+lOF
xNEOZUYv+FgwYLfhxeu6Inrd9r4mJfsWQoEkjHTKm5aafNv6OD1tHnz5ctRVsVDB
h4eG6F02YWhvAIFRCgKdwfgH5ObXCa02dvYKLzrDgIdb9oO8tcn5VTZIhLgoU7Pk
EhekDkpalfb+V4pkFT5CsuXBWv5tsr+IrpWourfWpD8OUea0qL/QIhkQobuoOm0+
IlX3e27QFkMnyuRA9TpUqlMM97SEZXeYmqO9kKKP9JDovi8TAkGaXyWr++3q+tss
t0AvNX4FxQQv0zu1c5kt1g2DT/yDFmUx9vX707FETaUUtvbnMIpe8vKmDwVgLYgA
wmY2uYyGFPGQf3OIVDrDmODH9Qc4V8oc2dFZ01SHftWU+upyWE1IpzWGrI/sMW/J
e22GdhZluVS31+8N9VKu85iJnlm7DW6sZi9sNSJ07oRbMwBoY6YbQPGNIrP/mzi4
Fuy1oiiOEhIWv57YqC0KmqVORVuVl8jkFkAsUUfkT1YZf618HMPTEQaOkqKZAo2a
MgvhqYHyuKKNg+R4O8I5UQnAVsj1Jlo1xC4kACWUWAdxlW6Jt2l50B0mt/b1BQmX
lQj+KgNW0ZN5DwrvSqUJGnN66+lGCOUEXGTJmRoCPirgumueAio6xxa6ysPSf+sJ
IT1n4JCxb7wDM3Jja6eD+e2Ry5HGJ0ILkdlsZ3MLkWPF84sWoP5XnqvPUuK1P6eQ
Gp+48fcSXbCAB+1n26ExWhV38ZE75qvrLGKRlv5Q6oThqTWDcV28L3XcjQOLik1x
K2zBxbde37xFLXxRIRcwkSQsG1gyc8VqzaoxBUpc0QhKiMeUxOEHekUXnuVO0fXG
Jz9P6Dod3g2oCI11P5yeCRxUFH9ThnK3fDmzWtimEpOCXxF1Uzlj+AuIL0k1xRaw
dqWBEO92uFhbaFMIHn9G55Cj2hMQCAp0qcQ8akTUWODlgQV5xX1Lz9NsKq2+xCO4
oGsIWTuVc8TLlQmJVQgmlylzYcEwfG+Bf0kEsqDg+JPSEOVd6mOhRV7thKGuc8TS
64N73Fb+rGl5KyP7ejikd490b1IvzCd3cw0o8EHkU9LVWw7LqMUO5cSkXwg4GR01
joRhWnqq7T3p6eAZMy6PxhjaQv2eFjsjkRox6gSKonEQ2jVFrvlFJAZ0gzsMY3Rx
YY9DXvA6ry+XOjHzRf3V2qtT+d3dSCqDp2g8cE7SC8XD7JvupaYI+W+kbHNGWbz1
7gNKONPULt0Fuj8/IoMmlaG/jV2IuNl7kra39N5yQtth8TfQCMpXYLDAvlW9VGB9
5T/iW3Xqkxlr/8Q2yJ+9SfxLfJHPkG95uWRoC+xmEsamXIPXpEtijVGavhOVJfAU
3f/w7VEPx484xNDvh0oQLQfi1WXqWO5Y0Y8bRqHYjj0Y6c2ek9Eo4s37Rvj1Gdal
lOBjDD5F8cKclFwNlZH7fcnBfq2kB8X0guvI5uaudg7AKmaJWjqOVAuPCsABBqXe
W35I3nxD5lmQMLPryIfY+L6wJwRTF12+mq/r1E9/Y6bmgZUreuqx0QNCKnKx6NlP
NfuR8OmBoILV8Arwb4Y93PcRtAD4S6MYTTYhEtITAqqnJl1AGMZcHGIHz7mTiN4Q
J2A8gs6gQzydNAU/5rPZAgefeClGCWpVpvgxzi75xAhXjI9kTpFgAsBkA09n1P9A
kTZnQ3N54Atpbyd+DVdhFY9mawgsLXFJ1kgsGeXQ88s3svnXux14c96M7MB20AfS
QcB7LB5pJTfTPEEisJKPv8N30XDnxl58Nuzigr4GUoPyV0t/6jLSRrblCguDfDvH
w9f8e6g/rJH+R6Jtu8mcELSWzC9enf+Mg7gdKYrZCQHCXqYauc4RiuhUCF3lUaqv
QPy1w139gv9ASoHvBHElWzLvMFjvblY3dA+QXTSxb+2EzMrmpEzwHRHHYLxj4S/n
s5rz7I9ZQTna6/Gkex9BffwvXsVcmD7YrtbNK0iiXNInSg8vm793eRy5pMeNr+0e
fwmvOfpB9uEwP7m4JVdtusiDrGu0EPmlLHOdvgmC5WegSOMW8RONhwjN/XM2PAuI
eg8yp24RKtqltD//+UyLPO8aP7RV5shxuJ96ImYIHPftvyxOZzb8pYC2UemC+/4U
KkPlScagptRWqE9skm2wJDJhkcOn/bjk9wUDgUaacwQd9aCnhIidmb+lPT8ELpmf
++PKyTe2IRiW7BDIryV6ACY38FLDy2PKtc/ND/qTopF8QRhY16V4BKQ+qXRwDxiT
hcGOkT3lLPBTECm6+KEMBHgNrIqHwC1DMx8tHuSwgok+FDBDxIWPwPoGTrEmQPEx
+y9YQMNwz4QSBIiRNBefSe8znDAfg0rUYIEoVeucYT8xZAvFx/Q54JzyDW6HlqSn
mcwdgVxjwAgqVqoD9Abq3kEn+AbMyY0DenRALSwDRac/xvrAA4BqBpulZ41Dum4K
SObdji+1eIXJxw4+4ZXGAhkQziYvyga93RKRTvVn0wK5H/FLAHLVdaFYHjnpeFwn
Jp17WWru4PwOfY8KaspKlubEFkBsqz07zI7DpRYQXJgs50AfCYo5jWrj0Fh8AEtT
/idzf3cMX3c+ulv9oUqldrovyOtCQBCUka3WwvnyaSJR5Wrf/20dvicOPBJzeL2v
+yKPSKC1j08pX1zrnIcuubIgo2D0hHVavkQYsuTJDud9ztLhpcJp9iUlyocG4il9
r2wyJPQgwfHi77rrxAFMcfrBUbxd1G0xFvjn88qoM24cQtAe71ZRs/AMMv0jNlKD
RSRCXIiwUwxFtnrLRHTFDC96AvnUVnSAoHcpkO/nO74rdVMIh5Ufplb4CkQ8T7TE
Mh6KgxvLGj23sXGn0HcrRIpAEOV4BZToWfFxe6chz0fDpHFWp1HjLZ86tvWAFug6
m7I+01ZkVJknd/vQk/VqyeEJq2kwWO5w18Ay1WSCtGoDqFvrwvz3OTn0y3Fxn59t
3ybvI03NFS8Z7t/bpEB5NYsLCyuj+LVY6Yp4Drn0BGopKwPJLZXHYpbUVPJY32E7
lcu7enAgYNNuHzq02KiVpWnBWdDyZftEPWFF6n/Epy1oKTm4wfG+ltcXzGSXLbYe
0EnGMABbkDrRY3QyRQWqm/x2SN6PJajvf3IaoqXczUMp+iE9+jwAlp3+sFOwikZz
V5Ut9NX7NqVR+PldTVTqsVsMjzkNydRl1SHxDIfVnMQSmV1G95Qu2mISgySiMOts
XcLniv3mySlRmezOkcKo/d9zoQ1IwEnnX1an5zpthDr3hfZQ2xUtrbNKwXCjUT26
D+7UksSEwzYTDegXrjgOs7r96XNtFkkB6P5gB98tOvWM/8p8azrDLPsZbrAvurXO
RJAqaZipxzbRPg35tyPY0+zWDcAFXUNKDl3QwNjxfunyLPBt+QcHqzZ2jPQ1PUU2
ERFDmm08BzGvRBJz1dDjYlGt2p/2UBaTaYE4Dfh8l088y4aaCu87Z4kWZpG42pSW
ulXR78survpI6B6iQRLgH8pVlXcXF4bH9CtWjYD1KVQjY08BQQndinslL3ru6ESx
t6YMGbqKiIsyUgLnBydf8eihg49H6uWg2W/orLwJAh4d+THMS9RFU+vb4AoY1gmN
JqbWmCGNSiufuY4y7wTl4K1eKBWl6vomxYUFWqEy5h+RlyimXUT8PXebJfeUcDlH
lH3gEoto9ehx36IKlo/Relh+d+leWGZJPAR5X3jJZaFMRXIhM6OnNBV8cGg2XSgR
RSoIoOMWW2Gq4NjwJ2m0x+6WKNDyx8+zIjcvwQzt+DfWH6L75eoMHvtHT+svDx3N
0Esk8O5AnBBqK0QfXMc/Esqa6fx69JY7JkVkFaTWt7AFnsXh4PLzy6HWUGn/Hj6W
ZhKDOAVcJV7oiduuDd6qvstm5ay0+mQrYDPJsYKi9cLmSf5JDBkCX5FU/xmfhEXF
W87nF4NpB6+ZljvDJyxXidR312blxjWZY17I4XMVEobA8eTJdwpUylyvFt0Xcijd
2eUVg+sKrq099dxy3zxwozo4Gmz/8M/xQu0u9fK/hcGcOe1ULkfqdt4AWTWV7tmc
C2CNmwdr/nk7D1wm3qhGz6dRiDvBWMimDm3PL0KWHFi95YQWvlLoVDwX+eWKb/i3
kKlK9G/BAsAiV1dUF1pc5igOdzCGXM41cHe7rJk49lvZ1eSquH275twYCmKm3DXm
sFdT6VT9yyJR4BPwZzFOaayFsP5l+BQsS77OgKuFmu7i6l79c6DuVlNXUu8dwTX+
4Zfyp2hkzN9Q+FDnZnoVCLxAS142p67GmxoaxdZoXVmoHbwUCBvXdvqMimS8AdBe
8sij+9WQFWR3VlzTE6BKHo1nxqScn6djS5wq0ueG8gEWWTmxBZa3scaUxwuZRfpn
M0CZkVYq0eMOA8zhsZDdyCD2J8Qfwdj3Ho3aLB2gEaRXNIgfGgzSPBPZoHdezuwt
RmREwOD1+s+bCDF98VlgV2Bbx/1YZd1k5KL6DQO2mxRBfzROyHIB9kO4syIdjj8r
leD5pyG3hQRJs+/w4nZHeRamGA6dePnKMRUyCgauib7ZwPY6a2FvrD/irSANemc7
yWueGBoq3T3jOfToPe76aLElcCKQwDygvkzEWasCTCd/jkqNK0y8mBsNiZBVK8jq
jpL5qV3heLlS2m3d0SWpT71fjRC1Hlu7PSKAVtcsBEFHPgJhu56HtsbAq+5HU/QN
+YGPvxZ0fWIxll/ufv2yFg0c5wD8ypF4f4Ccwk6/IokgJFzhaick68LyDlBZyDOS
DI+gYQuwnO7MnJVDrbK9eqZLVLpyV2OZT9thb9F0N3a250H7EJKV8Fk9Z0/V2XZ5
fV3Mdmr42AZPo87swmbVWmPJCkQwHfe+lfEwj40hlAgl8X4ZphvXBJz2vp0qgSlR
or/lxAJlivqnwo8xsfflPG8tcr2XMGibZWWJvdXEijBICYvAScsK7KugMSdfXGz5
XJUMWEtPie2VJ/Y1g78PGlB9+2igzM/9tNurH36gdlYHHkOmbFtYoOFnuvuSjsp/
LeKB9Hp6SGwblAc3+TMMB7OTog82fhevMTyn0TYHfrTpUi+99QLQOTTCuHhNXrkY
ZV0M1UmXd6YpErIi9JEQvFPLdRVieSAp+fZ1Jry7ZhFF2Nwi4wHesDls1Y3kt5io
uVcB7wuJr826Ke636lWlc4DuwyRL+d//0cmf/jHeAqbPu7rxsAnlnWdEtCyiXOAn
x9Gn7zPZEa9l8F2svedvd2AGdE9OUT7WTEI9MUII76Oo+X+u3GhopW0NbnunfEpC
YyBYpswffcjzg2A8+kr3otpkeMN97Od/hek6z+JKuiPtXWKmIG2rDtSyS6LC0itA
XuAwH9ZwgW26mZRycpGzXxMlshyl5LjawPM33Z82Im+qlWX3+aDLfx8DcrvHZIyc
kYJyB5appZ5eoj2e7JqZqGt6IJcNaIK/opc/dtLuEfClTAoKLIyDdb66TNp/5H3e
c9jqIUP8jS6y+LyWsyIxloldsUnfMDvIZmpSKWno5CCGloICGD200KNRT8cf7/pv
05iul/JnAo2+PA+UJYybwSnyNVzSr7uxg6dxx9rYv84vM4crGb9g5LfQ2Ypr//xA
zNLSX19YRyXki2Z7p7Hask22RnFmNPMdQLTplcMJsHN4oW+DadWhHSu67ZzGsORO
AoER38W6tqJZY9fXLo/Hh8em5ouVyvRwdsuehEHr4kARe3xnL7F/9KZfn52/vTas
E0p2Uq+nCprjx9BfQHl2qQVfBMjIgoFw++T92gDr3jonOdPD6YL2tyx8VqrjgJlY
5QEAwkXikE5NSybORynrIH1D6rOKPESoJHrBJr12NfNGyh+UbEqOluZ4WQp131nr
D37Il9nLk4gaqZ9IX16REiolXQKVt0lZeDpSPUNEZ6Teqmkt3IstNCS5OT/sjJ7f
POh2cFuMpQCSNxyTcqKcSx5vz9gAmaY8WnW6wC9nX28O7AXdNRL7NQ8EDz2IuTn2
Ov53p4XFMGMsuJiptBiDMdrgbUoU0xJuJO+zjjWb98rpIoA33TSDD29WG7k9muZL
I5TYsKgvwsmIgkAr7vvhVnSd0rn8bHB8eicCnu0Cq1r6Z6AJqE0u3uwz24xUDcTm
UKrFb8IVYf4SsDJY5tJD9q58SdLkHgsTaKyCOsbh50uBRvD8VLRC0ToirgIZAqyC
Ovx3GU5HFTszZ9AG8uxeQ8c/rX9nqtiE86dYg4V8UtAgAGKIPGIYJIQtLK0tHRYx
3+h2pEAH3Y+c9Vh+FGpicnlnqCcvQYqT3Z8eYH9SJRFNV2P6DJLBNAuX3Jw2TUBU
dPIYecGkkYkgglRtMfTAhUKmeBNrVUf0vMML6Te6/CaO/+Bmp/coTqfF66uzNl4W
bGyC2tD82BgHOgi6Yg9Z4gnNuHUS6tG81Pg/sGgVT2V1500UjCBFITh2NFeki96L
kqrRJP5KKIKb2C4qQNqQ7jnT+PGNQMtyomH3pv/X63LWy1Gr3Tj+hbbKpUwKySFH
Vjbn7TtmPGshdLT8s3L37MxTZaK9F9aa9bxtKn4GEHwrsSBmWEOvLWa8KTF3ntCd
mbxp351t3N4wrTZXE6jryVJQ+2GYGgepV3iyc5ELbeDq4NiLwpr6OmTi1M8qtp0r
euBH2PoMJ+GEoUpT6vbyyiryWxszGMAh2EEH5Ex270pWxQQ1BDxZCgP8M03jjFtD
T2499L2CMIByctdxL7/iGk+vkmkuSHU9skL5noYjKoJxASi7Y0Uc122W98buR7+w
of8pUQ6U2IDLbiRN6Q+gnYvhxV5VZ5iYzzMPhXR4v+P5ZJL+LzQW5iq9xDqAWOjO
3poGXvzLHIi23EYYdMKh7PrvfYX0pU9c/62KPJ9b4z8RBdiXA9GULNSx3aDG+sHH
09iLUeLu0Di59QMV6fGKV/kvABoJuHv/i1rTEVNWUGwpLZQBvLBX9zgHJIt04upp
bY8PhvbqPgv1yDEueeLNpZr1XLbgMIWjWGDEaYmuAZ4Esbb9+XrNKZNoJAAH3xbO
mlzUDXvNROotgnx6B7W0MVnec301m744HpmMnuNOUnAXzbtJ75YPB5GCZeNXs4Ep
Gg95/HzroMIjE/Fw5xQnIx65VTfN+yperzPR6EBr8Qp5QCaiRtjStIky44B2ZWe0
1LW519M+mASQtOpobpwTSjOhjOe/Hgi7OavvrGInXHCU3S9Z1kYdQQebIigUHMv4
YFO2bbKDzjt7dAiZ7Fdc8IEKT9RW7kDiW36hQx+Agu6zQ4tTbS50ZvL2fvEXESZF
TgsbEu5RFGMRIxHzdMGjYFSaqtOujKfxR0J802p5NQivOVGN2p9O2cg7cQ53a+Hj
dAHxBvHe3LTsTrqQqX9rsp/Bhd8XdB8wbc/ogDS62x82rXFmeM7WJFUrLkBUDqhQ
CMXZi/R7CvNvsrRnpFgtCAW1mEiZNZOPObU5RVrNjgEdm9Jk4xaRgNFkUzUbDnFb
K9TMowNpNcvKuHztr6CIfIAOO5RvUIBLp+Tua1DQYqZtpHQ7gnTnYgN0m4ZrlDyl
3pRF6n0d6QC2Z4zLTaqxwEjcV2rwqr2glkra7rmUVGmiU6X7T+JirCYiKWM/4vOe
tdSxExg+kxi5JIpbTUROoD5nBQWYCpsum39RnA2soe+1tBypDJ7rjAvh6pfWaS0u
R4Oq+5Dtss1oUsQzeyhOwnloAJ0+uoOYNxjTew4PAeJx9MboWQWujmvahU7DXgcB
FSmXDWVlITW+Q5cJZTzcXkNyJUEVAeGRvHQ1/W2Jse3Jjta03v4LkfE8qHizqEMB
jD+R9Jhm8NKs2bQrt6RFu5OGY6l/Sl6bGSrUfik1bBe+H/9i7F+x08va784E91vr
2z54Y9zPfYA3XpQnDzkCYSkzHY5KS94Z4BS1khdKA+OzF6fOeda8uFfwNsrKH2XL
cslDBu1w2HQtWpyjDts+dVBU/GxYn3hcrz4OUxy6R/LPjndaaThRueYZpGOxXnEa
ph8AU6oyHJd57g7pol1Yw2aRjX3q22tJ5OUdBcMgd+06CGK+Gk3xwVb4TGkcaoC1
JQ8XJWT9l8ocX70lTS4RkoWtOEN0v8GcWpcRHBpG2Led1NvJy5DdMNWy2peMRyN4
ACsi+frtQpuMSpvqCTNgLr6Htqabj+WVMs21gorGM1/u04vuDvDb+Z10RMYy2WtX
G5OgWK/FHuYJYS2CaEoMLxG/yPPPUKw1iF3XPXxBUGmgppfuuCAjlkQ6Kc8q2ZFE
BFh3VpT7OC67w3NXF8YDOMMMYPaNSpRA0briZNNepeEh9l1fL+4j0E1aNndrnJLp
KNbqJWTsc4DjUnkfv5WfRUz6egKG4IYQN0F7kBDw7YPaW9M7fDWH7jsGgyiSWcbO
XFnSgyrLte3MIuNgUfNUZrjC2mZuUE//VZeq067WXTh89ZJ29XeXQjua1m2RfBIZ
Ph1cBM0Ma6dfyfFcD73EPN3nfCs68V99w3Zy0QBb9M0EpAjSauEF1MMSIUDuJM5U
L8x5ZgISUNS0Dao29gcx6hF90c0DP/D+op3xil91hLJgYOh65zxK6LzDLg86Nbzk
QOzYkctdiDPbLcFFpE2l6lqi2uqMraxfm2tVxYFyDXA1Rz1JXiVLV3AcZ8AnYPTn
/r9aZw9VNDfCBl/YuiftzXYs/85PJpbmPxQcfPpl1qNeltYQQk+R1sE6GlxEufbr
AaA/9RWrc4CA8UISweA0gLRtCF3KxaX3sEJi9dRn9yy3tKiTTjn5M9fOfSkBUKmw
/5LrVjLGkiuW1yWojSe135GerN4vD8duHo6xjSxckIDJScZ02OEk3su6rjmH5bu8
iN9OItfrFS/SWwD19sF8SApcS8590dTXHXSzckFa9QGq9hhcFu8AMdXBEmHuVs41
VR+8Gc3EgzQ/IpqNTfHdlGHQvNO8BItqmozFhIQccu2fHJajmolk6s/GC9sxYufT
qOalTsaM/yHDqLb6qPAnbdYR+vyxwUcV8f3bUIBhSm5mjOSsel+fX+rf+ZS7kvqi
GvoBqI71EaaQcRp0k0pko/V/HE5tUQb7nWCdydsg/+Mpm5yltelsyCow7b9YpNTr
v0lJ6QJH7V3TuEXcNLVHW925aPG90MyUvLfXQX0sZUs3tj7XOpNBxp+mpQADEg5R
Yp3R/qovg9aD0cnSLNYwKY1EfQBU62RuYfsE9DoUYP6++ZweJsWMCqBaCh42BOGZ
BryABcgxKtDxpk0CEMTXJeyuoe/Xxh30MCiR1SIE7Fk9pmbBmve5hZiR3bJAtQZ+
1BI7LWufC2VaC9qtuvoxY96QlAznnsAi4oG5BRsInEDymZaimlzKBWXVuKhmubyT
8CC2P9rlnIQputMOJLPDbQDfWh4uXrxa1JiokFQ8h2e3kBhTvX74KnJXC5KnYcZD
Pe2OhPk7r/tX1dIsSvO3w3G7JcF0YEpBYkXTPL8YVZUSU5QT7xGRGsoM57C+KD16
gFCXQ/Hp1mEVQIMS/yUILVBPYg1Y9uEwYLXmmsz0sCxXmIs7uiSQzhPzHiHBP1gL
0gMrhSzStQE+hss5eDylr4KHNslmF8umvyFZPf58Usrxhjz069B4HTwf21UzmCUM
286ztPYhzOWPBGRA7/Jkr5Oozfi+UDzbv/fFQ2TFChMJj1bFyw+KdG7+Wo8gXnBb
vRw52ye7Gf4HF+RgqUOt7YUpMb0+mab4X/qM5X6CUluihn6Xt+iWvTTFTb/yC6Qr
yyfXhuIalyzL0YeSRu/cyIoi9syM/O6DdhfLc+Pb4ZWlLvmrbQw8JFDw4wyGvHQI
nYOau7zeDi0TJ/lOUau+ym6NiTLYWSoi0Hfk/iQ82/wuZXIqbkKgjzZvn4XsXJvl
yFU5X6Fycrf45ZyTa4MSES06BiuA6RouEE5UIwYXP9Op59z/7+laAYHLLaa+14BA
ifsfbu2QPMSrsq+ZoGVd+CvwrJdND10TAwCoZJ+rhjHWAHBK+q8eUFURz9CTA7M0
PRgR9Q2SP48gnEuk2HwljhEQlYlgBUZI/NSGAca1JFuDl8Tgpq9l+LNYXoBajVRR
WY/VJ9GknjnUeVEjRuU4cuggLQIcx/dmNOMOLS+6yjZg9hrj6Y07j0GaOQoqrgL4
9QYU/tiRsfHOD9u5kHIwDFlGt0XIqjyZPkC8ck5+JQ80Pc0te2wxL8pVwANlI5hr
BXNspWThRrYpxu5LIDyLSRL0+4HOvHeclJt67MjP0uL5CWIqQPMK44rW1bniUEvf
1PY4T56ah4t/gP9RMwxnAfBNIoIZtlmIGlhLnxyPdx6UZW1WnN4bQfDVKDKpOAw9
uJL7pJEg6h3ETBoRXqNuWgKU65eoRNBOgVjklkod/EjAzVm8uapsJNDp5CXa0nZv
+JA33v8PGPQyekTdePR1MqR2eWFxZDDN2DxYY7x3hAObxL+4A3UqkMTN3ktNmy3S
RzQKijA3EMB64NOzji0mm/jn6QvN70zWTDGcrHkasW+1YtS5XGxAATea0p0nlMcI
RZc8OIAxzRH2/3gebjXprNn6O/8BUQNnRzk8/OwWR5CFWz0FjvVW2NnCe2YNPerq
cnqhk2/3YSh8eHrc2NHsDxaS6bTy3LzcgqglPi+snWlS664zgTl2SZT/9NvyUM7O
3SXqrzWc+rXhRY93NsOA41wtcRlimBPq8djQAPznmD72spvVki69DE8Vzrd5SCyN
ioCGyf6aysuBr+N/UjefkHceeILEQmwn7mXAk0qyDbw3ARTY1fdYG51K+XeY3qzS
esY+HbZo1B1DlQ1jIN0+ncrYXEuKBzlrLlkx5ShKnp+EyH3BXfBmU9HZy58AuOAX
V8U409B5LH8Kmbpi079+puzNiQd/Q1Gh67Ff0vaq0DPrrpozapbVMt2LRse4YkPv
xrSQLP5mK3u2+ccVYtcehpzlxgElrc8svpeVjZoiZ+chO8L0dPINVrfq9gaLvHKS
LwEjZKGNKg1WviH0Bmc08LX/E8DIO2EIVBknCpsAS9xZ66suJDp/SY9CHfkfDYi2
T2YzkWn3Ys3FIPk+02Y8i9N7atXbPMVxlZ2dJCl2c3XXI212J6pfipPPcO2hrwyc
c9cuyFD5kXOVk/2rwiB1DdYG9DyfF3WI7H+j2obXaj8m9TguxuWb3Aivs0uDtCWF
JV6sMzstcje9ibCgRgFrEEcZZAdMmivB/1yJKekohxXfhg9Wq/Cd36cSVx5vLw8D
U9SBYHLRbqOJQ4b+S/KoFfGihom6QaDlI1LMQrjQalCur7bG9gboxQGTE4zPNOo8
Sv7cKGTbl6sHCixDY9NDb1Cm0ijpbD4ZEkYzjaMm6cBA+rfBW/fw3GDouMTmE/GT
Uk2aM29cECcJ2vyif57ulDcOZMN0RheW9houhIvnxWIIz93yOAritiuRP4+Id0IV
EENy98PXzp9OiIeJMnhu3Xs4eWgjBbAX5mbEU3f9Yc6RZOBVz8kh1ldxHKjMXfbf
GfAprHerhDPbnfAbLiWXgfPJs39IDRegdGx4T/VB2cYuy/oRWViXzy/G9PF/BAbd
jvt8trpxuZZ/ejbVeLfV40DChwV3iCvkVU44VA+SgsrUooXk3qUSiLEzdC2IqEp4
3eSNkyy2Jk65f7lHtrQ8q81rttPN41qx/EJVoEPpe4QV2JLi5nRAU1n2BkfhTK6A
vN+tirjZaOZ+mMX8hcD+sVI2L9do0GKpLECGPLjxGthYv+c7WtabLRpFg6T4TIox
fe0jbrB+bGpy+tlz69KYaUVPTeNlWjEimEOY9lgYRUFhnvSceYLE+9L7R4a3yRwB
S9qss3QtHiM7kmo5X5jjuZVXpxA0wNjjuLAkwmaFudMU3nTm75mmxWqMnRaJWPup
IdpwI5Ufr6yEQbgin65bxPA/Pnam4EGjzIbw/De7GL/bgESocvSnXBb5SpnH2U6C
m0G7qZHLYIcYj44qe4rNmL2bQkuPAEFm2WHlHtK7GgQG8C4OrQFwvb3sQtqPijfV
pcG62PYw1lmrZCNpq8CKIedxctecZOyHdgLqTz4qio1XaOm0lstuty+950yBZ5q8
QeoiUpq7xIrIweH8UYtmMpIg0ZYRaltcnVcyltdNZdCqaENkITell/HqQpOKMraE
xBOF4n91bySaLV3ushX2+DgGnkbt6Kn814on1BIMuFGDPJ0G4Yj/s4ao3RmsfiJD
vab6LCNOvilkTJy+wrUDik7Aloe2gBiS5tB4lhnLwYajbGNu4+NVBMyxgFY+BSCQ
FIDgL1uqWAxZg31QaYEQwcC3Lm8coJLMAqKsGiJMRXFBLibiOvhg8/mK5ej/tT6/
T+2YPUREyo3DMjBZ8xJASrGjQ+7DaQ6Nid23tCAuQ47IT1y9o1h4akEaW7JY4wWN
mfkEB8XgxCkQLVPvHPTZkOpgyAeNKNL6VmPE/WugnLP4zs5JFdCbGkK6wz2WMWz+
kCkwz4T1OltbCUxky74L4tEW1qdOcqCpujeiH+c7zhxYIdBzM3v6dDQQUZDUXEAe
vo5uo0IBAzY/7RGcyC6JV1U0i8Zv1LZR24miCkcW2x1cGFUg5JiCNKt+aArqRZKd
1XUUFv+KP+UVcwjpvVNkKUG7/R5LQmoV9Dlk78VLFt3Fmtd+TBEISjcuajNUlrSZ
IG1NfV9RWdEszB0x12M5RREfUPSYgENFELsnO1HLRamtLD3vzuq9QstzgiyAygBV
qDpl7zqySPql2STQpD0K7mRcyaDpDeMyTwnWKW8h5SSvnl7HnLsMLj6wL2DM4rCM
UHsQD7mCuktMxBK28uCnPL/YBahNpNvslsMXWbREvOPSUIAjsDETEQaljJUD8jrL
MWk0976yCMQVnv2MU8gWOQewZITqs/Kroknkvt8/GDPLzHVd9r1miA/n9c1sj/tO
ekVo0c8M+ngc7dHYc5Ab9N6kbipKlr/GqjLJL2RwstRIWDm/kEy0zt7XzPsmD8KN
CEzZu/LBDXK1YvJgJOagl8BTPzBRIWLbOtFl5wvpGtb2OPKRM0USQ1M4EBPdbYD0
J/JjCffvjoruyJlDfDwHReXE65uq5YUx/6T6m5cPHkS2gj3ifipDtivYJWSowE+m
Cfi1srhj/zxiNFMZa7uJmDIW1j1YrMAFDmaMaMayIQ10IvhUPYgq1HQR+s+VEhlS
H/2BDaRlzBM6s/+CK3fFYlFvSgPScdLjrHjix9VboPd4dD2eQW921HV/kJA1HeW0
mPFUwLfVG16k4qSvFCFv7hhrZUwufOhbYcrGkMIQIwIzz9IHy0oeYNiGP2P/m+/M
oFN10MhgIu1vcOns4V3gjE8UQsO9TaWvV/uPK4hvTuV9nZNKEcrwt2c7SxrL0Toe
wwVJe9F1B46dMkpO13FxnhBM+dP25lCQtOjDtwj/wqwHjm2fMfc3JoTPsQiSxZDT
mE7nrqFjjmucvUXHc3Ro18ytxPVJQ3cruE+fxlOznOJyv8KovcwPaPbd/Qept40d
X0cogYbYY6CMbTNkqI/Tr9z/7NaTb8L3aq+SZNnlwU0rEcm+tYIopb+5WTssOXiV
7bgMGw5kfKmIlqTAwYUH/6Gv0Bplgxz4QxJqroRPo1Pa4KQrXTd56ZXNvpBnX3u/
3cQkaIMDusM2SMMC1Ly4DGJYmppfULBRSD9vDxDuOtHwgW+hYYvpF4rY1E26xao9
wzOPKVwUQt9NtIN/L1ETkSMHypXlZ0Vzr9FcvOXbu8WQU5nuhZNefXStPL+g+AtQ
2hPaCBi3HKGj4sSiaV7YrlbdivLblvDaB3ArKYtA5q4PPcgr8dke3rC+/1TlkYaV
VOvRmI/GoR7l2X1eObY4QEF+QndKW0Zk16U2COPDHfbHTid4zMnhwwMO43A5kjpZ
AcmNJFalfZTzRdhYWVTFMkb9UgnvhwLkgYNb4ieD7EPxetJv3qsnQTVr/dewONNW
IjUj8spC0cb3KBRXPil41Q/9npC7bQkzBJsqRwkUfDBBl9Ljt3Wly6ST0imzD3Ss
f9NU05eEvTEfxJy7ebIghJRBrg1be0CmQ1XdbJGUOZbcmlYn7K104q5icXgDBzcp
35+1kdiiMXisuj5sQCV0r5BzEEd72NVMBSFQpfeM20H/4a3/FnWbpUmUxif438Yd
dfsV8Mki4iMf9ja8LWSr855A0nVGA9+plouaKkefZOIE0YubHgOFoG0geNFgnNpc
UG5tPzrhkYW8/itLFdHeZDOy2aNrziA0wQ9IzDdUFR9QxGs0l/dKbdmlGgXEZhXd
3cWz/ZuG9/7Nhgao+umaYNzllahFeILR13uReU+BPkZj2Xg5erYw8qc9ElJF5ksc
5nfuxbQwa35J1I3hHlUaZk02i3p9chZZznn13o6lQbtt6rWhGZgj6FK1/Ucb3osp
FJXRr4iJhV7cEniRTsyHNFP1PvmSM6uYZ/ixc9baQrTAupQ3BiDYwiUOTQy0tcjS
BbqUTToR2AaJoRv6IEdLzhIhJIfQX1POA4wlBgDp+W+kcLsYziIhbPdaJilYkwj8
VgLe2xs8QDVcgC7iF0PoxHl02WYf8nq4PpXkeYRuVUC7TcgelwzFcDSBnUuKtw+e
mhNGMgOnh81GcwqZCcAAFQfzy2/jhwrp17o33zMvL9tfKQkqZFTf9KTkb/pBBYu/
TLk6TN0EcIqwJ3rZAaHP3uQZNEyGrxLaXCXiK4+JaEY1/RCP4KmVc/AVvrJJYmFa
z0kf45aqhVFhTnfRNfHRy45RvReI7NVjEgCTSKa9y96VB57FH4Q3kjKr6yT+hh9y
glk/lenWemn5UMSav3/HcVUxnhAICQsF8XRH9WN82ZPtB/8s1gjPArMybcWKmRmZ
e4QW4DqpL0d5SZM0NuahqCQkulLpku6q06BgDTTrT6nEN4YusNW/HMykuWPpAs8d
FZGB5qpyWTTYW3PwbZfXIon9fwgv4bVUMb90TBqixTHJbTZRc3CQu9mPxv0oPayU
meJnnjtt3OWjX86eXioYuROloTxsGKWncIa+RZbEAAw9wLckMXX3n0yvo/EBRbKE
1ylwzd+bgAiQqDTgL8qzoTcMjOk2+G0+KaO9MT9gmmEQ/GdQ9MrHCgm0E/eLB0hu
noVZocq9FKhRxbGh5ELENUSL66GBmvwGxRsyun9pfa5Z+jM4JSRZx0aQZQdyVHnF
lprqGSL784xtuYP8BK8xYLdgBXXdy181h41S4FlI+qPbb1tZXFa5LYigrRKfAKsY
CxnaNmlsM9lVNwdApYh81jJRtd20ERTCKfBSKbgZaAsBtQ4y4/AHzyXyDwyMnp2V
DwCKcSbj+NenfM3vvGglO6yt63Rs6lqWSrueq13cU8gwv4ylpxy6QYNg1gqc/F5A
fjC2Uut/VEl7fqKRrQAnIfGvQf5TMOuedhbn/uhGT6tQVSEBzxqfYygmmTD1zAsK
hZadaYiCau8VayZQYMXUGwyb4CDwm4hlEW/FcnuUa25kZFigciuFIkYGJkt16LNZ
6P0iIMbHvHTPDL6SmwwlZXJq1W+v2V3eOWGzUPvYa2PN67Horn+7cgHNuzZxv/yY
EmGoYZ3fpr+SM+9qG7XQox5D7RD0N4ogFkmbYdAz7WI/cOvfU+N3hX+GHGiP5Mzn
zms7BB9K1E/2NiqCfQCn7J7xwM9leY0tMhIV2B7Ztq8JYsw7wdJcTsq1lNNn18vI
jq98LYa7hydH1fVB+60EHPnNToGhwkOG4YSAqs3ENbPYnN8iURlxVqQhEFER3rcX
bm59HZKjRtEvj8wPHvys53Ph+8u/DoRK853RiZS/85zVCNqd6FVMaTZbeVmOa/Ce
IAcLJWAT7WxQ/03VAW6wxJKKau25jys8Xb8fECtzFh1U0e/Sx9kCZX9q/iXDF9cL
rA+1gQTg5bm1xvzEloXi7reaeMASvSQDTmQakklX1YsRkG80BspdUalH7sVAnE7p
V0/qw8B0kaoA9UI29QEU84RD8/gVYLO7IsyeeHQKsrMDJ9SAML/o/48AnZO7KSnC
2rqF+6mRvyCvGNF99RNSHIS7EUfwkBzVXZdMpKbhbmoNerXKsi98wb5TkbACOKfa
6V3xcCyWWTEyrxX+JqF8wM3CaqjaqWCIiSR90ERLMl+03pQnpvKgtIERDEOSJ4tj
eqKyWXeBZp7rz/UJ8HFnp57DC/JRQuJBeZH1e0q2WfxVu9WeMP1dC1zNfcLGulqv
MCcBtzkER32enPXFJ7EhHl8Lm70VPdmyf5a8iX01ezaLhZYOuS4nYVNvdbmri6pS
jF1JkAH2a6rARxVdbuoCj5/wsbkS3uWTKGv9EbtEuah3WJkNoF00Y7zYm6e1Gic0
z6HesSMkYGq/yW1kkgiEqJI1d8WJfsrQM4I5Q4jUgRZ65IIZCB7lRB1Je7aNCHF8
f/r51t+pGuBR+ZtSP00Q09WpjIRr2QEpxIIO4jmPxA0rpcTaVC6eSaxkP55gZsyB
z4ROlb1b3tIaftUQTGUSqGCBE65zOz42SQctAdxEeCP90XD7OiSWauw/pEkwd9Kj
jfo0CaTmjqR+rybJal2BWbzqvUfCERscSMqW2qrqBy+q4cftU5P9uqSNtMnbJU7h
zijSjZeaxzAW75dCxqcWJwfSRTrMuPqMESJ8bAEe+IOLKY46lwzoTjOqcc3O/rJ2
7hAPoc7OTEwHUyWUuz8X5x/NBwGkwJ0X4cRVrGmwca7dju2kALQshr9YMKEeNHLc
f+iJgbOjtQ1IUME1Kw9g3+khPGet0AbzWJ85ygwqrR5xIdZHaBD9+eXxdL+QD2Zi
v+W0NVhhT1BuPAl3Dw6CtRDa4iF6/ck1H3ile2bB3knRc/8qY8RPPHvilSab9MI6
7mtDxKbJDDedAHxuO713t7ZTcA2ffbCiQegTJsC0OQ6I/0ybLsRgwRE9xiPK09Do
XverLz0NQuoAg6Q6SjBGsvpUSUoT3wyZQS2dC5DuqjoAXZo4nhwIKrjbXdlnX68D
GmmTz0CHJH2FpbJdpUt795llhYamFFNTChiad1MT2ClCwib0nS5NFzPyUz2ChhkD
Oy5xaJ0mToP7b1eHBrFRGXC/jaKy4zts2t7f/RgaRcMZlnyO23pFfXa9Ld28ZWxO
aFTL2rIJCYWvkZfFSXVMRLi41wtlW6OA8obfQFWph+xdCWZ/WRggyl9eeeOVbNgi
9NVOxrEQW+D8T5soob9OmnxYBIX6JYR4OW9ueFc6mgXzDd3DMyb0a+w1abvohC6T
JkJrh22SH6lgrEHIuTCrPqKD5Xas1N6QVn8G95IQLW+9at3IdrnBiX3PwqPahjqP
KBkh1lHF70P6GaR7v9QzNY0AC3CzgSDx9ap3GBCdSSIcojjkZyMIyaZaMgJpGILv
qLdyu5wTbdTt/NczT3ibS6hjOEIsmEZi6rEIU6l2Ropga5vBWNCn9fpxEQKn/XMK
wbfX7VMhch3I+nqPdUHktT2nw8hC7b/Eh/wQS7J+pkq7yAuZomMcVht3sKZNlGhP
wDzkbDuKIr6cqTpEOZaIKD0gTPgDG7VdOWd7B8MtKWGL5d6+Y3dnhoO1W+hO+veC
xl/vAKyMGbiGOEJ7SIOr2JtWu5Cu0diX9lDW2UtlPm36lpeVsaaxS/3xWcRpAYf9
bnfqbckMTQR5gJZMJeX1zvu6bJ/wQFB8aEMGMJHYsgFlZBfGoYDDaORug40OBkWE
oToiz0Q762HbVOl/RPqiyT4+CKi7X9wpJvVcrBD992jgTxZSXkDwXLaT+TwMgpyq
wwgygFB6TyZbAJGshn9hYjs3TamIIXnJp+XVFNMUzic07k2FUL6hlPfgLNhJiHk0
HEU7tx02get8+5lfUgcOrcjAOaBjRehlRLUCDAmqZTW75h26eDty+1ak1mdk6OOO
wJZSn+O8X3QU7GlKKmaNIJLpbxYMz58AHjOjmy4hthUY9JMbaJ4QiINqF90Xqrwc
r0Su+xh6k3rjOK2SSQFVAPgYsvCrWg3pHu2qok3ME4tSaFNIgpzItupBeQ9pCqJF
ZcuG8NeT8pAQ3JMWYLlaAI5aSkSN0aTqon5XxZ3o5RtOx7yLq4ZUtlj/QOFKyyB1
lwlCblpYXfGUcpwDWwuouWdHU+YP08CXGcOwCBETQ4syAQg8O+InW14O/+xi/b2P
n/YASmzn3algQDjhnSQz1LveVacnDQ1zKXlMhhu8Rhkckj91JUVMHJSz57cDzGVu
f+6/84JtZcXOhjCb6aYlE5n1U7Gt7sbcv/IpXBT3f6HulclwYG67ByEx0TUOoNES
6yKkFx/tV7PwY/I59CufCPDsdXjlEkKKykwBCf422DLe2O9CZpElvOTcA3cRyEsn
pMiLzgVRu5MQXAx6Uh5PjNL2kSW6jLFyzYJ4724KRAT2xUTQDohyeX1Jwy0rN15Z
IojxkwhcklP6PbdZEzZmh8MQApk4pyehVe8lx58eBfJGNWlRaPl2cS7Zc7Ttpgy3
khQdwu5JGL3a25RPGtEEOn9dixIgUs0ZuekQNUQYWWtm65e/9hNmcOWmoNGiDYcw
7sajImdRAYMgxS2M3AHvtaK+pY2LYyidAFyA6bnIPMRcKiYRagVRIQ7blfqlbz+T
fW80/uXXfvYOT9yADxN98EV1vcPuUMDDMTKmh63Jefei+eqeOwNusKuFI72cKuSM
YC4Fy4Sa5S3xYuS7WMjO+WsuqjNmGikDqjHvXbh0HQUbH0vVzj6badePQQRzqoeX
Wokx/lEZ9UURG4KNhtbODHUikeD7aFGtXp3OX25bKr4iGsqxUgX5JKDiqP6JA+eM
mc3e2jwzp5t2roKBh0/+8HKUlsdd1xRvc/niYtGPh90FFB3ifXEGUAndmkMCKZYq
yOmXhwF/UZwlxynv+rwtCFmDxotRjBurNReOG3n5/MTZfTEuqRvKWnK51lYKfFzE
qQObO89o4qKwM5BtpenHLU6dOVK3QRWsuRWLBMlUP+Mn4/h/hG416SNfuhW1Qykk
pm8C2VtOfCcVamc4fpiozHiUoJWQ9YtpQMkYZk8YCGyVwGEROSHfa12lW78+xKc8
RpyhO12vPRYbfJxlEUxjKVNFdDVKJNHQttyc7Hh5z6cFoIgXgBRUsibR4hnvT6TQ
tHF0TvgtW7JsdTALMXzbxCPujQg9x0Wk26328dgbkK+ltCtSn4Q/V1KuHYwQ9D/D
zOF19axAxfQGszDL5vAcKX4BKVZQF+5nomp5Z5TlaimNLwSwuVCFB2KvL3ZBWGmL
BDijpujDCRxQeytOysgw8empU19iDPhwWyeGccGxM4b+FEBLDTCAqD35NVgOenw6
yL4fM+zMxMSu89t/3XmkK+ax+I4Vvp4w89HnmrFnFwnI7N7FGTM2YY7Xt+PwyTez
UESlPBBBUZp2ZpguzakQNc4gkT4XABmrGLLVMTK4pdbg3JORkPKTYyN6/lP9Omgn
VHB/WgHqwGiTP0owmpcTOxOFzAfDWTCGCDMe9hWZ3gtKrAJNuH0Z2j7H/oHYwd/y
aOH4XIXfZp3Am+rPhMugRROab4q0eOZGCOw0yl8x3HmNKpca9VJounrW842pQh9U
UKyoxCWaEsiYKVZLQ2K1aInfN1qh+3ryqe7iMSZQSBpWCe9J4hgtdAikTRwqzxAx
ClWCqI/sLq6vSiE9m+n32IiHrxueGqgQPYdy8r6GauXyyDk9gZICyILVEpeooWwx
SOf9SEy3kd/a/qAieK714gaIRgYAhzIgyBv/CP3lO0hbbzq53LiZJqJkm+kUGSYC
dkj3buvIIvqpiWFqkpKq57vP1tRkBmdJuYIbGaNQDNhmniyP2duMdcmsQ1Zb1KWa
U85JfyeMSvgIBDgmsAmw0Ijq7R4Rpq0W71HZohIzpsJsDKWzEslprB352qvoU7uG
PlgGignv5WhdGQO/hRBaYLxinDyMEAmyWuGinCakrMjy3NbD17vkf+lRXZvAv7zM
UA6bp0HRMOhDIf4QL//9XD/+z0hQG1MyJzs8HPuf1W6OsXqCfkE0qiA4ss60JwjH
cWHU+AF3iMobz8egf4Xoc0JocD+ZB5IvocZiGV/MH5Q0q7+g2ZUIDpZpoBiFfdBr
UzsX40fWtIIRXHR8/3jfTcuxp/9jo2M35eM7kfyNdScFMJRY44TL7NsmyrMpVZss
BlmJHbWzVboXJxIxV5HO19uFZUfM0Z+eh5RKJuygk7W4+QL1HEznll7qegI8M6z5
z76eaYjXxPAKgd2WG6oaKoyqS75dMCT1eg0SLrjaK/zl5YXzz59jzypzZg5BmN96
+89VAdlXAIoCtFgEaW7F0f7alpOALE/iT7NUsPXdxSKMvMMPORUQy3jAh0m6s/6+
Qpoayry64HhOboT3klQAobjSpHtPVOY5HP7R+oqWqCukSY1oi1DRx7qdJSeeRB4Z
zEE8+wtmaOG+w7wRB09Xhg+RUKEZia/QiOBvHf77LbIjM7l16Z4fEkf8K1g2l80D
VdQWgIwAba7JnFoZJGW0vtpWWstt88k1vJ4A/47dos5aTm1MQG0o3rfjgwqhDZRW
TKEi5fkzwypz1FeCSBGIY7LaVsrfbAcaU8h3SQRo6sVFMssIV9ELvRNieZIMp2y6
Nwg3dFR1y/eZ/HoellwWNYdXS/XKi5KkWKdyp9BIw9TWgiqEBFmEd0S2yqRhACIp
S/8FHFdrU86I86mwoA/j8AN12Gv5uulVV67E3bKETF07zLmma1Ew1//4zSrg8G5j
wilK7rJ2ZApCK6Bled+tb3/VLKEDq1V5J0iRsFrYIgTq6X3Q5yd1itiYnWgUZh65
ws5fUsuNv7ldr2OHSdqfAiFIBHOUaRtdYWKMiUEI+4Ualtq7r9Y8+hajKZSlT3fT
zkMnwD/8YAXhtZBhZ6qtqmfV1ATCt6+bjZxxitTUlXnnogLuFG8PaOWgxiWmTmsu
FndvJ2kOYUjzW23tNbwcFxuEq5fiOKbw6VDYB4kNsSA+VI1LXBi4Q4YacNoCFEek
wgDFhmwyTkqkX8IgqpIDpC1zHwl1kgfaofGGTuX/rCnApFnfmV2fSHWGIvPeVwY8
Wf4zE0Br4j/qfbHWI3eybeaYdAcS1NSo9SQ+k1gC9MT/ML8jQ6DMt+qAMvDZ9r4H
QV0asp3UMmnSTc19T3v4ydQfHZkwD1kb4DVXU4NUEOCtAH29IDrhnrIw5aNgAOrX
HofH2l6vYSLL2BjQnqCDtfCTpJ0/+2aNRgRGdoQ5QdUgx+DHCcETPp4fjblRbLnZ
GFt6DXyfz3BIoOfv84aP7szdwoB/gTr4GzS8DTdTm0Rd3Pdwj1MYYmiR+CZ74qZH
Pp3Y6V6o8mDde3zd/svYUwCrTrT9C/RdKTAkZI6p1bVs5kDvTbX0lx6owOmKCewE
elZLwqAZBHh4OuTTshRxtc6aNE8Rnp0OuuzCnh04vsLHnUewIIpQ18r36dyKqSGE
e09le15ikTxrdnGPkaI3yZWSuLVTlqpjutz2HuaBBz82fgYTLFG6GEP9eKleHe68
OpFrEtN4yrml2wvtmCbI4SDwjhkIOup/oWGkDXQth9J3/n4Plg82hE6D7SUcn9zT
PGPhHUITPWBjWGZZhPQ37RWzaLAfsIWiYwkZgaqTFxPPN2KbK1XkYedDrNGhYyHS
xLuIDusSHFNThZpPVjWJhvaH6Drir+68rh0KyoHH9rm02wdVIsiTYA1MEi3sk9Q+
WoM0AuogPLhdS8198vMoXcU22n5A7MlN9aO9HX/3m1B1Qoxg6amVkjo1OUZ6U91b
ZzDW9wUQvBASKyFhHEbrvM+0cl3udWGNG1pFbXQjTzdWIneJzir4jvMwkxSy0jSD
lnFkzQt+Ee6ivzDR07QUUTrambu00sM8NUkFWuxpiy9902CrNnptHekJuFF1wQ6y
KEOYfHl3NMwXQ1Fl+xsdOtwe/sz7iBKEELJVgM3QDHvT4HNLQCpE0q4eAFoIDVWh
GTzdpK2SeN7suv7xzZf+VutdbGYd/zvzhjFMBBLGtZWiOJxeU9CpnRo0SNQVbGdZ
uOX1UYKVIPd1StzafJuKuJ8FQiCIOmQ/jyZAEx0SKRwlvkaz/jTKxO8oUt71dLWc
DTlRh8yNOE2VVS2zvh5cZiWkaBBg7r4/HmiVUeGBk613fLCoOwKbZMaXycM0r7WP
6+Z5X29oBfqkSEwNVxGgcELEaZfHy4Kgct5/s3Oj5hqv6unhB3XF64DmgfelYy6Q
RJ95Otv2fZG3uGWpT0wC0iYsKAc7u2JOEimiBZO1FTGprfsYrova2gHZLciS4oDK
IIp16zgacW+Tdf1Y+aqOiINTc7jYGwVU1VnTAsU/inXiv4ikqxlSsNVgX+5Wi4t8
TGL5SUZ7+BSaZaqo2s4p250bCVOQ8iRA6ch9sWlhYSlTiLCutai5A1ygVdIdLJ2D
+asq842yTQuxtdxE8sL5AXrcN6PPs2ZwxYvWeGuxdbWYDxAgfBX0enntvT02Uu3v
ZXTgNamYfdp8pNNCdLG0BBMt2KSt9Acv0uJsPbfP8gDUO2h7xxs3MMo9WyEXlxax
T7ctIgXoiGN18vO7B6Y0zRLti8+JnB3nLackCJKHW15ejbNY8CFecFL7f7gnwbAS
vnSEdfq9cWw+RuWNKigbcKv83X6PvaZd4Ry0aJo+Sl8DtG/HRFRgb+Mvp0Qz/D72
2vLUuvzE4D/PI4KU+1sQWYAc/sS43G+K6cT4cK6oWFl+Tk3WMVYHiY9RFV1St+6L
DV2NvhQ+4fODAbTlBJA54jvFw+u6mVOZ7TapUZE16BPK1EU1bc1ur6u2abLqMi/f
Bu+qvveHLulc3TtQ1AhOTblwzcaxlVgzzZcr1Uc8uW70dLpQPHmafHcFnNgCsBJ1
13SUcCUL0qvhY1Am1Y1GuDWWiPvZwKvnJK4+YZwvnZI2rnpE8d96RFuzCbHo9zzC
U4GBZkjmbk8CG/a4sj0bj6RL0ioWocmSwTjQG8sQBCGe+xCwD4ff/a0ZvJ+Fc/ek
MFtKeFvUNuZHCUIT7mEZaToK4S8cJg/koadM9zE3XMO8W7N8CaMwy3LuUc8YEcYb
1JlW6lrXlqAs893bbOu7CFNmC+syUnsKfXx6wlbqLqgr3GfgOcZ/PF4YYGU4mkoj
NhmRqUgbrlUeNSzyNBpqojmAOE7tAlG3nHQO//Ym65MfBXh/4kFxnUh92sw+8Mdx
4Lhey7AhL2Zns3U4GDzr90DLdB76MxBcMyRJ8nazjgbehdocSl4ZgiQZxIyD5Ghd
w5eY9fZCyQrcTuxmTPLibL1H2gD4k2YIRxm6P/ygBvhbHKmGvUUaCIyx61iR83p+
JeIJongcTwx2oHPcbsJb7mztDn5Cxu+0OJXHZ7IOaAASM4mRNr7vddGRyxqaCmQY
4BOyZwZgfjZaX+rOB3t1u9phvkQ6U71R+XjeiHeqoQb3vyUBZjKJRaGDb7twZyZ+
3QIvlPXewOFEcLe25+lZNLUIuAE1CK9wWbWKp1JvfqwqTqQs01I7WVE1XSSZ1hmp
e+HwpizmPg08ZxB6MeoH5P25npD5VEoRBTRITjsViaNPxeNO+BPyLd3yDBssMx5k
Q2Gi8Lf7OWTuJelssNVfJuzi49AUA3ASA4vDnxk5lmpXK3adm/aOFP/qCRvLhQAG
oLx/JqV5iY3CEdFOdRBn7lcB9PqtRLPuL3oulcz1JgXTXLr24dkxMz+rDwnMmPb1
biJ/iyz4bMiAsIjiWGdHhAm/LtPjzLAi5LFlkXXJnktfJv9ZAXvag9TXK7jf9Ng3
B5MO8Mkx7poBD+KDbGYjCVy/d+t/ATMCsHy9MB7NfbEGe91z0mHrR3eQLI/d7LwC
Y9VHe8qto7yg9II595/HKswO3cqTGKGIa1gKwzC1w6bbri/sh7amYUXPMkX3P2dA
11OeD/UC6Xv3wPCd41cXJB97gKzBUCpLNpGPIUoLiTjsRHKQEq7kokGqsPfhOwaj
hSpDLS/2YSW/WNWOx+ZchnsPc/oSAO+KjtmC4Haey5XOBbVk2PXJKdFGE0OPgmon
4EhPPP6gJ7Dq07OWy4V900QpVublTz+wt5oGdeyiotwfNZ4fwS1q2yiYUJtH5jTT
SJnAy5FyQVSRmx4gTHw8Va9j+k283xP2+rhza8hdd8i6ZmdaKSISxqc5ZeLxiEUZ
uCOaCtsnOQzqBFY2M2sWxcdVNr/qqAfbJRaFGI3VnDZYh9FRMMVT6sRqd8Sez2CX
HqMT84ujwoGBXnzCyLxbxBHdU9ZdGPTFf08yOXo6bVz+YJiuaNyN6LLw5bFTU4k8
FwDPEKbTrPFk0NcJFFUZ3YpmxbbInuGQ35xmtxma9bGDykBAGbPrLfMGuEtxs+SX
KSriR/eRHhwOxjpVC7QEiZMIhL7ROG6M6SGI5ONRIC4fXFnRCSHgEXRuipCu8PtD
D/qhJfL1ztJuRGFDxSvYdLLLUo08uY5o8+yhAyns4LV5hAeQhWIEWnpXf6xEuGP4
8fY1cCvtq+hGmF8WxGCw6nNv+m/5qcRKfNBTdocDF2lge0AP4Pghh8fOPZxtqMlq
gflmKTp3aJ164RLGFCm0Nq/jnSDT6GrFF6BAbZL/QGl16klJVfTxkSDY87vy1cSS
jZTSG84+j9mOyTwT1pRsW7VdQQ7J6DuaF/wLUOSqoUWPY7jNAB9i8iZPzX/fYkzl
w2CPiAQlRBs6plIYVa7k30Y09RrIeqIGpgd/4ch5pP1k9F3qo/jqCXgBbijZd8Vv
PeLDecHjTNuEamfUPtIDc2AaEMAmLIJO/cx7nFwEamTsJn5mwGrrZJB7TIECr0c8
8LntZ68h8vGE0zaM+W/2KZefZpOu2euk/+NX3psV5Gha2AcdKaMlg3zl0s4Vv/+9
oxHA3Q33tCoDyPNaFLzISbS+7+WLItQ5j0qf998YMdOaEUYEc+yxkQMrqSzcew3V
dazZTI5HVikrJuh68tVl7K8blM24LrisVpGsj5lNoXPVxUyeuLBdOMHJ5wuSiLBm
BBHUbAYVHOkBo2dqJxH0/1Oh7SPWerF5SslQv52d2YfCgFKJ5xoFSiXeP0bc+Abv
9MDJUntyMY5HxFpoc/IfpHMCaw+ILmSC+P/HJE20MvivRGgm/2pJHx/IzIs2Dyx5
cVVK9AGTLmO/jXXdfZxe9X3i7YwllJyjFpenf7DAlbDgNDiFea6HKvZeeYPO54+1
GsquehNgBw3X0QGw+xZhSJb6FNcRL1FrYJPiaN+ZsJOeCsAlFmLrWSIlu6Azgo8P
An8mura9WEcqqaM/hJSQT2Iv2q97G0Y6rdg4I3I5zbHQljBNCQutW4+ecq8COEnS
ePc4pxcrCCGr4VMft1F26OGIliNGkDM9H5TBdCjepIHRyskJMHlOsVIoPVvUJmMd
B7IF6W6QjQtXhyx8LnlDfDzNIc+3VcnsPLgDt240MmgZtOi04qNQ9PcParaZ2k4y
RT/ubrBJx2Z36zKsdHIRshWtyZNJfNl7Q2ip3fx/b8F+0tUz5gSsenueMq2pTGwb
zjb1OW8o8w1wPdyz11P2m3UABz+T3gU2BdGCMHXv5+G7yb9OJjlE59wryNLKQe92
yG3m8Gw9hvwWf3v+otfIlMdkNF9bWNfXR8DV1SZzQ1/tJ3KP7BCZ/zrjqwZZ5Pja
NDp7Vti3dNd/+Hd9zEuHLthiNXW9wmLuLJ6DN+OFyp8ykwt5lXxCKrrOBj14TCu+
tDxoc5X+W6qE6rV2cM0AGi5FwW/ewa0w9pNtHSs9U2ELTf8g9CbK1EMVGvz9sDdD
p4AfR4tFL9UZf7+bGOenW7M6NTz1tKJlNWa3r8xLCmzMpugkT3WjJC80gk+T7W8X
Seh5gDX3MzQAW0yOI2u8842BZJukDctCQw6deFAjbkYGScGnmmmFYdkPcJP3KqgN
8HhFMWLxHgoEpk2PDdRWkfjjlLuWxcfaAdXEjUQhYQYEjq9u2mqfPefX9QLyWXHW
/Fo6zCXnaKnosWX6gg+BoKSkp8Vwb/j2/7r7wXPr4glmndCTZCEcRf+HKcyONHJO
o2dKNoc07olM2nxHhT83DLJGvFuPhdbMKhh6y9r6runhbUGKboChWdtIuU0/2maj
gR0WDrzrArBWTm3IWrYypK8eXils2JbS+3U60bjHSgv5kYw/HkLF12nSGEGtSjwN
LTOJ/qe5v8SWocQa8dnV0KQEEZxmxJizdGsZoaSEEe6xPdgsvolWJKwuT+YgPJvJ
nmWB47Mj+X7rTbuKv6yFFrz7o40RJn/qUX19kv7DEL4Lh09xpTwCWwixO+tzHKnE
e4CqdEErUBmG5TC1ITRm9klnt/I2L8H5Jr46U/E9y037QYrY6dVjfjnjzgyXQGyj
VLFV7W2iUysamF/uG7IaIuf2WLjgG0gtx8PFosTkN9wLmXzTNgpaGj30OpvLShpR
66MOs2wEr1ybB7XibtI/xDChObBpeYhSQk3XjgDlCzoKCoMG+hsSE1rtnJvXUd+x
1AQ7g2E7Ll30Qq5cqP/YrpBwjPLI4n3zOeqAO18vcOH0jgAZNQfLjqSaGC8vT6IN
FBLLRMPdVnjP6VO3H1m5NkSnZdVd21zoM9Q1q5q5aDOmIaKzD4qXuJYrVPJebESU
3cHRatO/JYHLqT8AHnehL2/G3EEgL25PNU1MCYl5lJfDde7X24rmRedfGxPom01a
MQ7uaZ+ltp/0dI37pBwupvwi4cziFp03x5SSJcesDfVK5eDvzEGQKYO40CRqOe4U
MFWsiH/jwwVwBk+kDuVtmlKtEttI0aM6rvOLqDOCnkulmFGoz9a3XAvkwVtnAXvH
Yy8qLPtuI05qDooYak/nG6ogAY9DbwGQwuzgOJ2wM9fmzpGyVyQK0brf+aycAQFv
3ndRjZhqzVxJg889j0+wbDtmvoNL10xCGYG6cZpi34ROh/JcH48zqZE2xc98m0H7
t6bSV22EGo02Y16S0vyyix52CK83u+qfcG3A1fmsrYcF5y2jQes3h/mAh7hTEo2n
zpFy0XmUwd/3ei34/QJHhfrc08Btn/6HiEpdyzWul3YcQGgH9xwxgLqkjI0Iqjdp
Ej/mP2CyOK1fkcSqEP1sl6FoK364ImHYQsJ3SXreX5cAJ5eB6Fq2G2ROkGWKtr+8
nOQ9d/nIk6z6+i80dlrK75NL4ZCYOJvcqJtOEC/EAVN72dwgOxmYS18xE/TkWpYt
Y40KowUirEP6zJ/LR59ttYulBdUa5MaWiw7GgAMLUbth/J3bw0jskwy8xMkMu5eA
1T8xBwbcbBZp2jXonDwzQsAfl8BtvLkOHQ93ENaYpSNNUk4rq6SX8zk7mL4ANVNG
HD6nyI9oZW9WNhHbPzlHhDF4ogDQb0HZMKf/1l3LTShthfZloyFEfevP1HrzReYF
PB4TY82bdbGK0nJ9mug3FJxETFe2eOMNPhbo+toiNpqEyuCz82hKMhHj4ykEfXYg
pF4q6LXPOS8Y5xQ0wjtNl8t+G/rU7t/6y7d9k/Yx2nukfiMxl2GvDeiziOW77xMh
oiIUod7JM1NYz5Lbgx0UgMNCKe/8zXgGL2BwJbbwQIeD68/mNPgCIo87j0tZ+FOA
4DvBafKTqfGydY9gUlDl0X4VNkdWvWr5JTHRwIV8bL4ARk76WA8/jq5C3RVjitwC
QEJSRJpXznb4KrrPc6jlVdWtSFxHv03PjefzyaYsz0kHAJ05oPqBSxDCT3Rdm87j
riOUZfo5GISwlLFfjPWANjMGBPQq2YgY3+5wFe4E3t7YKounIR6PLdeLdRnJAJCH
DDpeX8AbqFr2DFWceQFXt+0OtPFvLhdGUYk0rvDNkO8Brbti727OqOdgE+/Lqt1g
/X7XdEuBCG0TuigGrKw2pwwD1gJmghvOIwEYKCLlc5qq/C13do8V2mjt46nquvh1
RQjbdLdjT4BhQOdjfD5HpY1v1y0Kv1/2Sy+gxq2K6SNks9JwNTeOGjREbZ+2sjeF
TK6TBAHksuCxwIIVPBE85znr7UM/39F6gsMvUAmrim5uhoYwhw+3Q78Kqz8Mjcwc
asmqoXYvfSBMUJxOwQFz4hFoqK0zTZS0D6SWERjxvkMm7esXVvYmWM0qumgo8CRg
uJmZqCJ2RqdPxR0m11Xqt9YvAsgyYYHtZCI+4fIXAii3sT6y2VWVUfWew2OnYGu+
8u7V3yoXY3pXtD01L/tj6w8dHuEOSQl6KBNKXsmX7Y/7k1hXKdDEFodMQ3rZhzXj
OflO+Xx7apcsJGQjfOBXN2R1O7kDOdy7/JHKnXqxlsRiKVc+kT7gHmYOkP7CI3i3
QvZ6tKQyglHFzacDfexylOVQxW06TYDHkmGPdsmVvTD6XZm/or1/qLnzOtPCnZul
lAskSbCpi92JSSNbYIEYtfITuG+rRj9gIZcEsDszLVKP5ConKC0n3b7ItSAElgKg
qoUOjjBjEAaQE/ZZzs1UyqYKuhTzIjRbae3tB/ckC1x2l3Y23Pt0D4T8lW5EFMoC
j1ysoenVTdApA0aDKItKI5thH7AhWHTsS8KKoNe3d1dup+5p6muYNKWGnnz4tLnf
aTqEMPRasRfF1uXEG98WunfV0VWPyJhMSZr1yR3gR0Tyw+2WnBUDcTrnXPgedNuU
c2JfP4nlXO8hyE4BpKrHrNpA+Yr8Nq3SeMa++EJ7VGlpp3pAZZoR1+XpN+ynMgtQ
LEfupigaPZ2iGwUvY5XoBRKRsRW/AO5ZtlMtZHce9gM7q3BDy8zQ0RcwBGRmQ/7R
wCJTXUcvY/vWPQrRB9ZcCH9GcNHtJTGk9JE4q+bwP8b/UT/nGaEfVvbDxFtwd0n2
Tr4BOp8dqBwEDGmPKI3ahbqPtoa0mBMMEPkMqdlR/hwwkj63lkLFLZy/m1qn8114
5NjX8oVGWxc8OAZhXaYpKvzZo3d1+N1hPuk7c63lvUBPiN5DNTFfodOKNSD9SKev
fcwdEFMRNoBWQxrXiEGTNnEAmtQ792ZPL8yDCpAnutTk6wxHjgttlkLu60dQcewL
kfvkUpDDxXUc04rJ5/m3y46ZBhp7lKPmZrbX+GPJ9M0l/SCUYRomsKCtsNanJXqR
iPMATE2B9tz3JHmeW0KF6lvIELZYxvljYqzMvlXqria2IMzTDy83CAz7jKSz6qEV
PnX0zyesY54LSwqtjJwAmxyiJdMcw/efUQAMlnm+TY1vS8hc+AEwyMvFGWviQWix
+ah9m4sYNjjPbVWB2MDOl6DJKFgHh9ms4wItK8To2pMSqAWw1vRtQkKDKvy2Azii
mU13iYhvVZh/DkstZY4rI75B/g4vGL6aeAh7Fh2wFV68UktTwHvgcA2y/W6a39TA
wKq8d2po6yLncvVZB95eYJ6TMDlO0UbOAIYyTO5/anc5OedqsnpxBSfRt1eMcBmQ
K5tYSa9mr4RB0OO2ICNma/oLpx3qJfTKu9TLm0kfYfSUGtWLFz/7/JQlywmYKLaL
jOMode49xx6AE6402gU4Sh/t0M4LHnfJ1GzNe2uVRNYtnBaYMwEXi6GLEONUSutm
YuR+hRhwZe3xFVxKynh8bAkVhKW/LT/MsxsA7pGI/iWrRW5eAjd94OwFMZPAjo6h
TSQDphnaQEtXWjVTIynPJpVF+M2MZAqzgRK90Vz/oDF7BFiKRV8Zrd3zDPJ9ZWkD
hFhzS9ZyPbsO/Ivjt8h8MP4CHtV3nfvLcY6Z5674s7dD5qZM7YtKjs9sbv0m4abM
B4UrYym6hQ/y7vmADYTmgOk9O3RbEVBGXoC2k8aDhcHFu+GY/9Zu07KMvYAvmb7V
IhUXd0VXNTfevTCAd5nnjFA6df2li6bEuYKm1fTVKuxOI2uuc7M7t6NqovQIeibK
kexPjUYrmjG8Xq34hOIBD3j/90UFRvD8oAaFwOzmx48SsMm9vtSZKhErIQptwRk8
HO0t3XVSxLrTKpuo4ZAZVs8NmvYsnh492kNQ5L4yJnhNhKUPg+JTQ8kwRIBonx2t
X6sqSQQlHDVm+9Uj3PIzCvgkBBUsL9sCHrIPP1tJyLHep3uo0D1ORirffQBpp0Sb
NvmSFrM7jd2F8kK+ODMwuk6z4QX621zq4q0QfxrVHKe3wGlPY3zE/txGKgiRSAVm
WpcITqnE8PzCSn5oiR5tWP/OkOZR7HNFIBlzq6gooeX7AY3GGSryl9Yz6dF/jBCi
wnpb3ecnYBo6zxDUj28Vcl+y3ib+vG0+v0SDaI5Iq0LYt0TZoYb8pijaigYss9Mf
HfDUD33agwAtRlKQ6yBR3p0ilxxXhwRXu2N5u7Qz2cZGxE1Wzcv3OFsL/7eWhXrm
KAkHXFEufU5993qZqAFNd7M+4WDIVENaLR9z07FxaOW0iSR4W5dIfq77AWBEDAre
Fqisha/ZR448C++iKbuJYwXZAi4GwwxNa2PyVq7noJRm/HFn9/8QWmzW9CAtM9Xj
5E2rwHOi/4NXyagZz1iEIxBrCmCYtQAfV45qKVIFAsonizJil5oPS7xcEUPfN7+t
M8xqGVmzod2vDVo+M8SixqE87VjMJhR6GLgiXO1jWzbB7uBu3afSSh2+rXE+jjiq
wh8HTB8/wyhxXbukPEARz9lAdUmsjnCsM0HhFedXQvFK3TLhYXSPQGiTlnPtxYNB
M4HNmea12F6zFT0zlvDawhDNydiME3Jec+k7RWjzHKoaZVuBW4gcMGhVD7AMg9ha
FZtZhR24PwISdAzDSDIUctFUw5bMo905NtxLn59aF6KW3mnUiH8QefLTzJjrskni
KzsyxHx6QoWaMn1WUPW0RFi3tUp1ZIYN+rGUS3JF/ZrUka/0SoSvJIp4O/zRpGui
qBtioie1++6i1fUmiTpYfw95X8gWk2wCWa9f4I0buzfl3eXJXM8zmiYA1KG6FzeE
o/GfVJ2H4MNL75Ju/6rIJHsZOsnYFackrtcj8xz2r8MNjQeqKJNnrWPP6p9ql2F7
M9XP1tQqOVqPS2L52zVQo3CuIuFMfup9cvYBSGFWhBLDX84P/KhvHEvXmMTihQbe
WxEuvlNgMNpGtVV2FbmJXT85SmAWQ2JkP4HXiksnUKO+mLRX0XZN3B0+Utiyw4K8
jLHCV9s4blCrFQsHK9wPWibx/1pY7yzY/paXI1JLXFPoc+ZgybA50vFRJ6gjQSy7
JW3jPhuMVkEIWmHvE6nOQr8VjHxJg+o47u6qNjxgr0PEb9KLRrebDD+SCUfWnhBO
0DGD0ubalIt14KFquahWXE56VNu1500/80SC2MrX3g5un4RPwerEg4xL+88lN7x0
1p045CochpG79dlkgq0cLewx5VDXp9U2D5IDkKVMiTD6WSxHDXGPpNgvDFrbMK/l
ds4h+7vWsSVkkKDjC7TIL+yiDM8QMt9gYfm2RU3vQWlbuaswp4QAc6StJE+I/IhX
8LcJYMkNF+TdjS1s0eNr8akZw6KGeaHOzmHfj+aKVyjoeUkK8G4ju1znDN0PvGgm
yZYWKtrYdTHxmpws4TF3cRz4Go61T/FAvP/D8IbAEbXsl+INDU+Tys+SvwShYI9r
7nTLRSXye0q+SFy/xMEoHOtecqOYO6oN3PQkiPb0inzl73pguQsVaGsIroOce7aL
Muo9ir4iGFn7Xn6tk0Oo4uDQCHiLBXPbbS4w+FDzwVZI2HnPdJEh69usQkJp9H+z
DYI3sfR0birWpPQCmyt2Wo8rtOD8N6Z4TsSHHqaMS1WydkIf7VdBooSHiSQUxA8o
A77oWS6lGNIKXtmFOoT7N0YPMlV1wbCG/cLSrYN5G6581fBxfJeKslGMlwCIcobu
kHtx8AXbmQqFxKtjyNJFr16W93FKK0q005WfH6yqposW4Z66XAVqxRXYhaFJP467
nHYF3mG14fB2cBauglfzo5DDyegwChNFMzi5zBmXOyWM98tHAATlXhmTaJdPU9f3
E6jVl6NNW7X2dF/wOBaMLIgl4jL8LzkPHJ3IRYmzp2NSKJ1MU0uDu6vJLvXrY/kW
1l6Nky9sOXLp392qd6ky6VNsOlQbxi5uYg7WmxksxbOMXqtWC41RwMaD0FOe0MsV
6vAkcY+p3Va84kQYze7KxV+iFkQe5K4Ja12P/lSVZzJhfaKBg3H7jG5ci4SHR8qw
5NfnPfxzGMP8D7igen48XkZt9HfSXmFvYHmP7pefSQ1J+NWJrfV2K3MnfFEOrcdt
hp7TfIiH7QKK5ph3n73QC0piOwNJYw2uOuPESQ5J+KQ+HZ9yd8l6oa9Gd5stTt5B
IGENVCwQKSxc5Qcrda0CnDLW/vRXKnXov4zjVPwD60pW46P9W3dGHapKr5lzQk37
YaAyF1fl2YKQd0T5BoTYo0TYMLLe0Ea+R1WWgkxfzw5ND6Hviea7dAa/JBJWhELC
ErX+IPQ8NFwkl2vVtNQO6vBxYlwJ5oyLcXcupX4I0IwH2LKuwfyPb/In0TKrzDtA
dHTNdT6U2iF1JbTxDspQReeosa80E+rZZsDmT1DJYz69Qy1JCuFy/0HgY3eLhx6N
JxMoX5KeW5MPJTCVKho2vSMlAS2MrFs8XoYuSWMUmN7R+Xk9SaHAzeHnHKdgmuyK
rhgQxOkZJCb5ckZztgkH+vIUsDEs0oDQijaJ6SxkJml9GSY8c7YFHrgwhjbaIF8p
5DHWJo1A8HEa87r/dHhAJJJqiR5VDzvNzyvAH7IrNvjAP1eI4pJF4/apBTm4mHND
azZYqY6kM7NuGQz44F2zsonlE/DcSRcrwVZsqPuxV0IdopXlCK2BaSqpPzK9lb5/
WaL7x5+Ld+DLtysydVyhQ+sEeCuARTG+acXlP1F/0MPzVLtjK53Cj1+64Nq0P1J7
+q1hLycMEnnkrZSBevcoFIbbzDbdXPNVatF7GB7fPSK8oe4PJs3AXkHstKOAHQ2C
jqKK6duUn+iMDPmJahsKiGZm1F76EK1pjWwAjO/aWIpElDVF0BBuAlk+4kOXiKHb
baS0mkQxoy5w8OvzuUHEXzfhnSeyz+XqihITE/6OMUsi3QIBSZQnjgVeNnXLlioA
e9wA83xxFKH7GyZKvnlt0upUnVP3TMZw5vU1hnOdwIBbtrJjT0s+1PEmGIJx4vg7
J+GOh2puvu5uNyOu22IN/3GCtAcO1R3UzDLIKhhdA1uHVkGsTea18HItEYWxillF
zrINFnslqHWtLthsAF3U+vr5/sqGgzzat5O9ke3EDW3GhhMzpe1bI2Mz6mOXnCyG
wLZGFdM+d6Frz7uiWneWeZq3r+OKEzvQ3dZHywLcKmnPp3c9ndBhCJOm4ChKLVvr
hxB9uVuoeWWnAO6lMLY4OWcTb4gBS6OxsNvo38bZAtPb+rfOdHqR07VwG7OZZNv8
GWqt4dQxx8NVcDCNFyKhh7Z1BuuGNBLCMtwDYWLsEeQcw80C8AQwIqFo4ueheA9P
SPw2/fbZv7z8vRuWG3cqv7Ixi0ZQ7aGu1Z2IZ71EFhvzJ10GALY3jHiON2+Jev7a
tJJmeB3lF5ADT8dvZ5L2hFm20DjWWKtNTmr3nseL0AB+EMmjXZerdtmq0hinLqU/
N621QkgansgC6kTyWYOihlsXY+p/6wKHiZ6sfSjhJNfmaKBcGdQMmeW1iVrGqngG
HzALBgFoomKunRqjVkkaq3r0L6JNkSB9Kz3NVSl8s6LL/Ydi0XgtuUNTzZAGeMwf
tkDR6p3CoTahSOSMa0+tnYCM6xC6+1TAFpYHG8AEqvowIz8EFW/SjzsDm1oUiU5H
gaP1yn2eRKkopvMVY/tMph/qn21IfE3hzAdCTXU5e1qrOYVfd59QBgixmXvR77tO
Lf4JsL837qXhUlqKKQgnuNf/H8dDlE7QiL178TBjxqCXWFWw/Dg3lsbmtrGaCRqz
LlZdMm5wmKZEm62DgBifcdBr/AjrYjX3x2fVL/xFIYbEC7oSpeuA8fc3MiQ54K6k
7tsRuGmZLni722TpDBVu2xE/lNd+w15CT87jbvntFarlQfaujV4gwHvSBstDA7Qf
4PMhoxO2lgvH7SQdbObUlaPl0gw9T4uIALw2h/jd5zQSUlr9THm1jEY3djr6Ngt0
nhINtz0qgLbNHyl2XiOWr1mzz2MiFI5xSHuwD3LsgNV4RKVbNb9rlsBU0NnBXTIM
Vtl+SleEBCuorxOUZUn7gCgMRZOpO7jcBy9qLQYaOYm9dtM4LSk4r220ik26oxW+
4yVyRzC0RymQobJMmomaGSgjaxfzJvhaq1lgBgq1gTGGRZsLR9Vk/KMwNviiz5H0
Yq+wr8+EpP+9u+L5S/3p1Kj+roiWjVXp5On4y/e7elHZqOY7x/JG3XYKYrRb/U8S
xTH+i6Xc1+UaoOkt1uZfxR9NoxANIQ8xg7SG9cQ8XOXCzlJ1Ok6kg0QIdmYqq8bG
aqaHBl95ohsrp1fztcvU2GcBZ8EhRu/Db9ASp6p3BFIDyukkyAEG3gbyv8TDvLQ3
RBMUXiNXyqmDg+ePFLjEHGH44rDlg6I3wJKWvj85wqVWVTwlDIrltKDa5zPm6Ht0
BrB9epCDpv4pfTce+IWhAaHbFkBi9bJa8BF2iKQKLONX4ITqQdF8WpmGFyheXHqH
Rx2bpUjG0CFqS9TSUQ1TClCx3NrNpGO3SzS87/Y/nsPZ0jne1Jx2wiCI7H33g4IA
bBSgs7IHyYUGq5QsQkJj9zsRUirXN1Efx4d/EY4R7ek743/bsky/p94jC/fAhLM/
fjvjQ9+kASs2XmsBXgfSslqix4PdU5lYyR6EpEyzMbSJApVEz9H15BDxJ7n0qhoS
Qij5+0Vp0R/BeroH8mFolDcvPKXOdAT8sV/s3EW3C7HXKp29DjL5UiT1LqLQz9x4
lbh3Ese+KdY9lE5jLRgB7Q5qwLKEBHcPyarw4/CZWNELjbq0CYsulrlMhFDHGC0S
8iCSkKNHLcd6mI3KqbtgHleD/8nAHC+Mt4pR2d0TrrXwNoe1wfAUeWHpI+8rnf5i
nQlw7sYTBbxFfORTyXQ058tp0wlfthyegTHNcEUmGUJ6qm4Y0lDckEjXIGN8/Ge6
AnYd8r6Mv690aAgO+0v+bQULSrM3qcpS7vo6aKPg259tMe1Fq1Ql20tt47kYjO1a
SXHWSfi/bnW6g4QdjQeLqamaiHsN930P3QKMa4jUHNSQSuJbxh3NgKR6AKgzhwPT
yOVT0dD0uHdra0lyRCOv/blez1fBOgedNe4HicG0noZUMLpxth3OZt9iiYff+Jr+
0l6IrEBe7oFUBd6DjKOsf261sHl7b18TKSigqbccOQEP493ASjanxtY8b+aRksVd
i8Nho4eFZRU0Vrlxsqp8RPkecn62yp3ieqEUdWoAKwyvpu8zdOpeyaxHGTb/f34K
nAQwN+uDstCY/dtI9hDoZOf5d/VgIbU7QJzKetoXY1AZw1Yud43XSMfPy3DL7XnP
vrOem1TDcLhkRaRDFVopY5QTf+g1NbVHSaqG1uUw67gJVU8SgEpYUw4BsKipuJJg
6ew+xwgW0B41D/ZBK2/XelZjQkG/SP7TQ+znyjE6zynXtzWpXDK1yhLCkvpOQpgp
KFv/ONG/dWYpc2omQpLzap84Qat0fjF+ubIq19o+D0mikA5QcLSYUi9RvQoXvZ1M
gDvabMTEx6wkZvPzWxKx5EFsK/E28kST3ldgu2nczN4eyG8j7AllFqEMis3eCkaw
1NzWCyYrHn0xKHhtB3aevUvIYnXLecv22M8FVSx2HShvrduzmJ/R86VVjs0dCA2a
BDbWeZQmN1GHKDVHbPSPIN/mEXzIXGq+QSYVIsoC12o5DLDJ7NbI7b+YWaGqP76Y
Uj6Q0j8MvqpNPVhuOUVvZ3Ri/l5Ms1Vsb4YrLcq+cYAyO4HINQOypMbZaDIVIt96
/RuuCFCxDHsl3kGtooNH8Ln2ewLt0AIdxLdTeZoq8U7BqdmRDJT5i++hTO2dBurx
ZxLjOko18FeLgbPq2X+DODF5NllJ9XZxPhppc4yCsKSLtYzQUv6s0utmxAnJfnh5
B0zantVOka5JjHV4xnsMFiBjYgNciocSeFjsXsDPNLob7sXTr+X3H9JgdZu3vLfE
nN3lwUIDRxgRjPt0xw0ZU+ewy62NkWgB9WHhAmCvquyqKJwzmPDyCxW/qIb5uE2u
QtXdJkyRwlNdcWi/SzrAGgklbP0rHYbgFhpVkTXn2cXua9e0+2shBJTKuHTKj2JV
d31NJIeH6CfSHM+/OlKJRsSEzIGWzEaHQCEqtrpfLhh4HeUH+eG+tZkq7rjf54Am
xK4ZRnbqO+WXMsgzSR62kOWpea02Lz7P9VfbaQ+J8hJnchlta2SAY8MQRG9y8Cz0
1bld93+PT8V7YiMiwi56OmdUl/DABVib16rxxHKAT0byhgPnK/3b8guDoxVaprE+
IwBjT1Ldp4NmKWVyDe0J9CsqFULyTtbGERHI4XeZyVJHqIvnKCb2bT3EJC7FuEI0
pi2NpBhgMdwouiS+7UZYVLfWUl32SHq4hacRyDSG57+fr4ov+xGmx7vFBKB/elgf
htyea4omcrzJmG/pPka/vmeaQDf35EnPxp4ItCvjaoU5rbj7z1b8tIA+vdTP/CKg
f2wwvZzwkmTSHLjuRX7II0/M3MfEe0/EJsYw7TmiX9QQir7ODilEopAQ8A/GWCNv
U4n0z5fnh89pV4DznMBxQluAu2SYJK4mPsqmTv1HRgMqfcjhCDu4eBHMrYfyeOFy
Akg4/GBjzeqd5aYLcq50OqHMb2zPxWtN0TRkvFzObnwxwk94lZY5fePTuiPk3ZQI
VDxyIUSYGgd1q10dGZXBo8EJ0ffm7dxjHLVCJHO5GBiewCvwHm0QGChbniiELoB2
AvgZw3yHBQKiaJxGzW/xUsYd+SVhaZHc6i7Ug/Ttlw8AaY10kTdnjCfwtSIOM9MH
lT/ETRwTx7nOghEIxUiLI4W4pQ7aMfobOiNcqDxwfY6cU6Uj6If+2ankjMH0zQV2
VBDI1MOhe4oAFxIneOXY5vItK+q/bznyxWi8cEFoO8czkSzpSHMQkIUX6HbLy6JP
fwk6PNCg4/Fbm5rDFw9dqeAhvLMNu6qCzeMvWSeZDrHlc8o34DsXNhf6LgYg1R/n
L0ldRiOc1zP29xC54Yhh455GRjhAWVZUSPlFm/cxYqhxzNXBPPA9w3ega8ChPXgm
KcTROCdLBmyxC/HrXo35GdfYyjMOfdjpoBIhVcgw4G/Ue5r8B5mmPtxzkQIfxG/G
I2NwY0pT6w4IXhOGvcFrpFohdSYQ/sn0GITAo+aT6zwZOHU1h35ZhfV/yjAXFDp3
yKmfv10Rrki9NOV1WtYgf19CRIe2N1GTXA3IL8Ac6npTHcvqSmhGt0g25mGCaFht
XGyLG3gNZI33N3wfIjqTS/Zj8yt5b/0WkneSkNPtBwY1FObWzI2LXaBWe4qCFmlS
MTN8vgRTlIVnSkENUTdQ8cfMpubwvu0wB61F8Vp8XSJim05N3Uk0L8XkLvL1depb
5IFt7NtRoBw27g75+pHC9P6LVcgU5D7/mVi6onX9Uw7UVp1H0tFHpM0HTB6nTOGS
6swz+VrqXH8tx4XMPDIC0hjNvCzoa7zwlQQbxB6LTBIu54RVAS3UkTfT42zDEAtN
9IB9I36n20xR9tmNMA2hMztAnrRuJcimnEzS9CuGu3lFB5MA8LkLc17ZuJo7/hTc
L65iRhGMVTAuJh3cuV5hRiUFff6O4FnKMo2A4DDAAB7Zq13m3Ka4QqOoYe2pgaYc
qrr4FrrUG85LzsgkVzZxgV6DnpisyiHJu54Y7x1ar/5SIDoKi8lAu5oLnxDrP2w0
zpYsQy2J0UqDlRXzLcbDqF6loG1xBw/M6SrJxqZtCsFkIAsIVzcgdoIqkgxI4DNa
XMgaNQLOA9KbXB8g6h2DJEg0U0AMd10BF6Hp+ZiqVm6i20jUSO0q2m+m8y+v6QFg
6gEU676VdDsP9qRpzfijCAgI30Z8urG5Ga5dE0dZdfxzZ+E1W5xL8g1D8eZUXg/b
ySYVTC2F/Q2nXxC5UBRLgUHywkvJx3Ls1+l6JZBQpDs2NYyol9aeQOWWN7xeyVEQ
TzIHTZp91+Q0UoOAqzD2CPqR5Xwhn093SHtZBknKyXk2sIlzBvPR/BfVfQaRdjYr
uijXa1EaUfWVdWi/g8AWm05iQy3rdQhq1U3KjzS5rWtrACYDrfZzPROC2Hg8KZ2m
rbyHM2tDka9v6PN7ZunTM1Z2prSyYvreiCdyRk22ocO5RTYsJQS2PobXaXuPinKv
zZdE6+9MHFCZA8V86r1DyyxAFsq+OAG0a+VjR9LRGzDXO43w7J8jX0ePVTBS3GXG
3/LikmEbIREo1qanTtuUQjherNqfcAk6rbklGvCPsGUhd05gDBob9Jd86F1fIZtq
82UdzoxC8mtYzFwdoMjnEMjoPUM8xlteEO3997hPTbom/h+j2o6AgPxPRSki+MMy
gvN0QX51RMHsq8+MsH5hhLtTcv1qEO2sFxjzJoZTwQ2quELCu7lEgswiPXXiS9Ni
hHgE+34KPSqU74MCf2G6yrV/KEUbhol//pjr3B/P86OOBqC9NedTdYggfKMO4Cpp
3+FQi+IyP9pbJcwRXbIgAzFGehrekzFjDWsP73tjazZveZOhoGa4QvVlLWCP8jcq
eXeTFX+VdHk0qW8dvuqpkD1ozxNApzlotTPjbiGuKqamURJz5qtGe+XncSLcbiIV
NgzkBlf1GfNobtgwD8iBhuYgmWi/qcuk9qAanMhHUYbfbFKqJ6nrSLHVcSU+XSBC
hDUZV/ozJADIxgqt0spi5yI0BwlwOSTn3Y0k+E4g8z9atjC8EgccpuCJpx0dQOIY
DE43oKxLveMLaA90tH2hWGvx2Msme26UcRfU02/0jSXG2e1/jO+b2BLTSYFFIi04
KfAWhyz3rnK/RK/0YVMuiWWvoEyL9QHMn7l/gH65jFAVauUyz09bFwfkiNGYUpzd
2MYDwzVDPuvRynUYM9oJ7rBJ+BYGv9DSr5kOdWWLlY+laL+miiau1ff9cptNeIwx
z6pM1vzCxtBwE2LUnkOP2MQap2y4faTCPBszryhhXc340TIeM0f9OiUi4A07ueLp
gjt69pvjYqr4A0+go9NIMn9Rl10ti5mBWTIYsRNrWZk+2FnLc40rbx7Dv5ysJFdc
ta8vYm14Ilz36DtBEP4z0UALHbW/BThIAfYDZYFwQ4XIWkeT2Z5nx31eBiC3uVc5
VNkHmGNJANGHhBH1pUk08hWhWGwpAJOePkaG2An9lTvVHmmxJPEcABYJVW50Ndg2
fT2gGg56uQ5218qiuYRTKK1fvP8e2VLUp6JER367gO146kjJb03UO8CuWjyEBPOo
cVMcp8WOsMjUxrermiFSJg263m9CGxtBi7VVHMmjwXN7TwR8VFmfKGBDlm7rfLOu
scm9dQDd56Hcx3v5rTf3m4BKrV8nBRIYg4+EgN8nYwjkoTv1sY0S0gC+8gtMICcw
OZsAeFbRJBEq6EfZ7yiZtFbcc4e2ISqR6xoK5HOwQMtNeGgnN82mkaOXI3+uo82K
QQ+HuB57ocLx41bO0UrZYoSOND2rQYunr6LtjQkAmpbxEb07TaZ+/Ojn4pEKYr/P
N/HSpLE63s5ud2exfkYC3KDg1MuTLVzMDRrjG4BTOpB5Mn71bOqciCnLe2fdZrsl
DX2ZBk0gvTRs1vK3wyUmfgXfN3HgF4bOw8PBJuKD7PYTkyMw/NfybAEK5eRaTur/
5jR+cceA7m+Hvo+zkE4+fXIPeKeKktqiqKJa+BsUCC04aDCq7/tfAnoiAdH5Nw6A
DYTpN2JrQk4lqfDoNzWNpGXHFZhID9XqHf4+NVUW/+nIQAMoCBmcju7M06SvbvUG
lAIsvuuLt24tzbRFta27s/tn6NL0iQsX0KOHm0v7/p8kFd4zojfINqdfhjw9O4dE
V0zMBrtFnZywIlic9nUOm/NF0TXlLk7YPwqbKi86Q1gzeJbFcqfz2N+nv6PntuU/
PSOIidCqC+lFhzirsCG49iCPUEgm8DquBAw+xpMrbFI1DzwUkfzCp3gonn6CdYKk
GfUKMXtZ/Dex2c9oH9KxeQaFJJ2MSyzqW07HTnP5WpFC6e8GciDfZ/onCFQnjI50
SnZpwxB2ToemI85EBHCNsbvwu71vIoVoiJb/tV4w7JxujRrEFtITfvWzxZI3UMeU
pFXQFfZYPm4VXBKsmH3MX0P/A80hcm79PkfGtHaFaleCFYteOl8QAYfF+BNApx6+
GtxTC/rKechlw2B9HroaCp4vffZ7CbMj0Ky0Uc1vkXucTVaWdbT1dk7Yi+gn4WO4
AfJ2UCxrJYP9EXv6boKs8MGOBefLw1hZ4wo27U+Qkf7CrxpX4BIBP28hMgTzXWYD
KDVF4RpM4GnXcaowNu3LLPwaIx+5nwpGPTW2pK9IQyRaYL+i8OiKeSWFu42JzKPQ
fg42TEMYMMtKxll1Lf95olzea9dlavDds5QqhPngG5ve7mcgjSeZ4gYsvT81iSf7
wETiqGjIvvzVwIkwmT7Vz6G0NM7KkGcaNeeDWbbt/jwbjKpQTXb7DVxs9pQhq2yA
SqUbIndiq+s0VMPBW7jCE/EC/kdKmtEQn9hrNZwlxcO2X6tWgl4N866ZGJq7l0LK
HijsrwQkDia5vrIMXz1x3uhg6bis+uiW54VQA/8z3mrm/1puaCFzr9wJvwo1E8Su
X/nVR+jnNGZ+KEhq9+8Jkot6W/Hqpj05ryS+cXCc9xN2ywgZtk38wBWW8JBsBDaM
N68eMfcuOtpmGrK9vkdLNia/4z3XzZVLaVWTn/NnCMCnnPQy1eTxYM/5teQhzdex
f0WyYTjdSr8qyfuzHgyDJEWNW0LkTnfTkomAt+Zvb3ia1Bv3rPXQg8I5Zv3+FxT+
EpFSmhZCbTnoYqOiRXLNfXmigm2UKrO+1BfOHH6Wq0WYOhF2Y6w4NOhfcCz8bzyD
6RTC7GVP0bqxOnw0st1ZGPzzOYvyq9DYeZDys7Yy6agikkd5wH8PjTIA0L9XBAJF
rBeMTJyYA03S+0sMrB9KpSvjXH1DaxzcYa+Zp9qVKwKDtAOSytAmfBldgeOITDXd
oUamQQGOkZizRlUtLJRnMl4KQCYEXwbTzNIfXex0N5l1lJSOIWO3a860/z8HWcb8
EKIcghxYdBxe8Wc6yMapCDHUmyNTN1SI1VOxWc/ocWMQVxXUFf+Vc8F7OEwzFjn0
VjSO7rxIdGDV4VrpQtgxWCjouF8pzTj9lDrMg6YikWML1Usj2VCMu/W3VMY2wbbv
lxX1hCPK8hzmv12nhzoZqYS+Z1Px9H/wRUeDJb8LvVF5L6qP1R3fg9VMzzNztPXS
ua4XpfnnaTXjrkjWu2wR6EVN6rWH9PdX8jV19sh+10vRqN5Zo36LVVZ5K/Fyfqwe
lqAi25Fz8UaZsBi8OMb3Dx2r9IP95p0OO8e/oBane9JG7yXCEptniUUEUgTbriah
jAyQIpTMzCisy0B11Wn3gn8H3AHG8cdJ2JIbsG9wNA6+kjw8Vdecx4W+BvMVMLbq
QiZHf/T5HEyEJJo8GlDgM7iocj8JmNfA7SocwJJvQHrH5Dp+JIV9m6egUWMpuFBi
z9d/RW+rDOf4q774H62xN9/P1XrcvZmGNvp/PDUWUJXSeijrQMp4kDP+qlKg+e1K
8eCB3YflZs9JGkBHqXSMtmue6IgA4KzfP31Hx2hhZC/LHwLybPMSgQbuCGMvDS5L
XBECaT7ZPg4UAT5OgMGbXcPkr6dD3eTcubmD9KbGNPhBatGEwIT1wozcPiPCxhY8
I6UdNB9haEf93wmKqaVao3TbtTz7uIJtqpJ4BrL6rIMK6iMZ0k0Yqy0QSWBd45z7
241CbqHjs6d8Pm/Wq1DNmc5lcx2pkrNbG/EvOS+Sg8D6+vZJ3FMd+1dOviyCFtc6
IMyT4r70nlrU7hgehMQy/yGWAAo5kbmwa9zxrsfwNmHYoFWD5pHFTVt+gNMs/D0P
5PW16Wa4wHj8b+KwxoRYringOVnY7o/IYvIPYP5nFcZeL5q1ygZn7kOxBKbWBSV0
hCN4AlsiNALzN9oSBAc/I5wcZSrQ8y7f0jMSjfjuD6cOP09Sza9RIzycB4XuVUii
YDdu8NPgGShaI45lBP1VUFztgJCfb/El5nh5z2RVgJhzY1O+2++UeZJPyonfTPDF
oEbPaF1io2S2IjjjIJTeBbr15s+fuJdJnxEGfFPNTz0vRkdMyYLpGSm9ogMCOqEq
JE1RSuVmk+PQ9Mo56GyUAl13ootM66Tzc6eYa15W6PNMY9WePRp7C//zleKELY0Y
j4EUYOJSodGZu6T9fbNZjTNjvn1sKaptmuaRGhhs3MRBsTh/HYJfQVAcRo5SCS7B
qTT7+mrhTaVn4PqEAXNVhW/ZscfJCLVYTGa6U/VAXwPsFa/m0yejuvJhkPJCMtdk
3tY0YZmpYySLNsDJiCJZ8Lstf9pZgEWvkSlXaHt9wVxBJggUZBdDeVGqiXFd50Nq
+7hKq/m4NRkrY1MKS1cRrRG19IUDJYs3HW6mYVmW+e3C0VRONma01M7Vo047inbk
U77T8OGQDxCwzQWFZWEwRomWGfzx994W88miD2a0lqbxgOO4aWx32GfA3hwcwGmQ
709oaAOrSpZmPJ268s4wdblCEcS1TH5EfNJVcOeSYHqKuHk9F5ijfbMD8Hdy9Hhs
09oq1E8XjSFaQaStIjy0dfTHATSk32B3LFW1AzpV4JqEZRH0ubUdmcT8N4wXxTFu
ErAAqck1zE+rwuRhXnF4flw2gaYn7qfYiPzzLGeC4wxO7Sq+wVGLVcMMfVH50rEy
2SimW7/u5V4mZfHgzakJ2XRsT6TO1yBqS037YoauMN12vYlgTRprjbLpHjB6fGw5
DgwbCHX2bK/Qy2jKMyvAGjvTztqrt5hlfYU4GRR0lTftNwwclOVvHM+vHfQADZO6
RHINGU+sZIM8Z8mF5TukVDj22KxjuS0DsxWk5T6Xvf5Xi1A3DaoD810ZTj+QOFQs
BccCQMtDvU90fomt8CYaThhhzCdWjTWdQ0EKYaTfXRrF+PbXqzL0+Olmhru9FAdS
+tL25yne6XD5fw+6R3jNYhluo0hZ1k3E0VwvcFsqsJX5X5MBMDvwV+Fn2Ejq7rb4
6VcgYvU/bu88IkH+oEpNEhWBrCfHijG5sNnvDNMoH7NP6/cYechA+XQA7IQ3b90+
jwAjNrarXXt5LpXu6pUItaWCdWU2x8+7wIDb/YR3OAqdi3vMwbJ8+lKYEOGzvGEQ
yh1u904fGhqbeeZlW0RCmO1WTxdKICY9uJAww5T1kKh0bsRTuYJODlwx8J+YAfQB
hay5m6zwWBjFhFraMV2eqDzNU/PM8TtL0gELizDS33GxvzDlibpjR3oswHcqFXON
y6QxoPx5P56V+R+vUNTZSI4tSV/sXdXc6IXiNPdz2JTRIVogaf63SUpKdkCcCHUp
34ZK5RMhMjEhLXSuvyKyJezabnofIpD78pvFCZzYHFG2R0f8dzHJ8B/KjK7f5Awf
qq+5QNnOAQqlXfq4WM7i7KkHmnRnxIh527Xi5D5Yt6gkMspzdf/qvrX+xUGIQ2zh
mGlId3deeJbLYVWI4fIjN4ufOrfJOBQHO83QzPquiE24H9secYot4N4STtjL2znp
0DrzfeHqb6frOT6CU24FMctIBg3QDkha/8+v33OgndXm7PCMhXSkkgcW/SRqXYx6
vx2A9Dh448JSpIst/cD3Eb4WXcetCAi7DSyWkbxaK1DLNun9W0YtO64d3B6DFlLW
Si7mru9ls1Z0GbTzmVoWwtmuoQloqCXtaMyIocGaC4qAIECjANK70l7XKg14Drz1
g77saiXrKAM0QSy/DIuhqf0adnTnmgig+7C50bjYJrBaP3LO59TtYwUD7qQaLUVB
Dx4Qnz5AcqWPX7ChqdHTyktB3JQT38GM9hAVu/gqBrU5GgdsSPp4M21JOR7X/O8L
Nn9+h8GZsKVawDlVFulQGKz6v6/sLEFKp4xYROTuiT6M/smYjZS4YNapbe1saea9
v/6CKHr9GFjfAxbfTx329Ws3f4NeAPCD7iQfv2hgRgRlHLSp3nyEqW+aPRPuhcYk
sMhBZJcEQNRqaQuW71PJEy0ZSTxwteuZZS9gJke0Svw+N69Y8ow7i8R4DKHtUJYy
VsW0v5Hg5Tp3crp1drt3Ax/J+AlS5gNj+rYkMoqRUmuCS8QBpXuHtCOhUowelJKd
ALslXqBYJllfKblWn4+1ZBHISZz/gjlF1ZEQ1l0i5VL/A54USJmrJ7vMRNrMLVau
OwFf7s6DZTxjRinkT0uBdz/QH53KJ26Kevcjm+Wgo1Ukt6UHFvHalZkCxQwk+4Xc
WeW5vUr8Yv2BHzOkI/UoI46LGwOPEHzwpDiUl7WkBwU8brJpijuWUfuphVL3JLI9
a5vmlwJ5fFl0YiuWPx0nW1pvWR8bFiCdrA7bzxOlOb6MyKI0Q40w7Vg4ch+8JyV/
ttdiz0DGxFdzoicWwaHoFtz+MzEfwVo53rODQZKl9InsL4jPPufzTpvSvWjZt0pQ
dhKEjYYSqsJ4FFQdkAc8m1tvTQM3ywY8yRgPO1y1exhs1FmRQEL6efWWLJ6FrYWV
4Aw17SVKUC/TGysiZtlQRunKMHhE0NETTzRur9aaR/XOJ4mxU9d/3XjQxA0F3leP
RCHyi7uYAI4n/CEa/x2o5N8ajFfi72uWJIjzGBIFt1kitjXu2Ur9VMbpWt3Pf6y5
6JRO4gKgRWieB/yEjNcF7qyM+aPmXmODd4y1DloPZmQnAE73G7fpl9d21aCrEM6K
6zWPM/snnRfWnmZWpi0RNSv4Uh/L62sW1L5uA+LiMZJvnSW/lz5t955yVOFUC5IJ
kh7n0PJQQ7npuiSGbwLrTVpqxRawgyiPg+OEpegheXAuczbxwljx+wGH48gGIuyw
LWMp8J7eFSaTQ3Mj2H2IVihSJ/1smUJlATHGKOIIzoZ8lv2dHyamRoj2psMmZCR0
rb1me8s0e3EEG8fl4k+dAzaMIkJhnpN8dvmde96VoIGwZ2/kjh5ftUIeRla6Kij1
w36B/TIoISbdzeFz3t1HVg0hTVy0mPz3XWBC4VQc1jww0AXEZvt6iG1DDniPNFSf
qyxdgaf9U8cPYx3/neO3Rf/hG5UnJivlox2OJXUs8oAhM5d60SAPLMcFLoYO8Ns6
EjyO0+ohHUkdU/hT8AeQx10+xl5xHtTR7sKH8ugP2ZawshFgOA90iiXQkESe+wJ0
Qr2TzjcbDUzPACq3SEvANF9Iiz8AmTYCy8FSDpo4DgIV4IOcMs2S9e4CvEoVGgJA
Ln9aAjV/LvBBoznNl//EB8oe/a9d2gW9zt3BKMNRh7EEoBFhd8QMZtFaPF7m39jB
QCuw6jtN3gLZURfJ0C0guqxJDN4sB8lbr+dvjh5Xup0lcZWrr++MlPxGEOuBqq5C
2AzYWwHgwUnpzPZXlKv5UP4mRnREMIvCnsfRydMDUM9Q4xM92HRH1L+gSLX0Y+uo
LkgDj3BeyFmmQD/DOfz7HYKHLdD//5kfaKy2ul5xt7Fwt8ZqjH+zDIszvzjOQ51+
flhBtHl10R9hat7dsvlK80w1xFYiU9gvbhXEHHnjD5t1b7h9hHooBd3xZtVt+JnF
wgdllhshZmcdMQtdPAF8noAIkIeO8Daq2S3pD52NDg69mCI+WJ6PNTJPApl20cAo
QirjAGVK5P1MGv/1PyLO77KTuJ8vEOMXXirHy5TEJov8VGSBzYMGa+V4prKJKaZ1
Eq2wPHzrSpyD2uhfx45RK9tVGSpuefgCh0jz5z+W4Pevf4G0daKYycQaHpJzom3w
Zy1CsOlcM7+0ZbEfUiVDUXvi/2ZrrpFtHfXVbWwL8WbytEBz/qk5JEfY+i0vohdb
3TLv/VnYtKIuSQVeVAIkdTrVq9FMQLbVrmTwDPgxcsqwCotdgF9GVuAOWtsNwqPp
YMzIGM0g1UQc265IWDpdyHqrLqy82F9EbHFH4oCyGHArwH2NgSeq32XPK95piGSZ
lTUy9nVt1F5ZoGsvY8drPPxeukqsR43Q0534YJCz5eXtUk/9DLkNRpuv4FnitZm0
Rc/z6khxq2ifxhBWT6QRatuSmQM/JxiyY10iicDxzbpOUjyirPjIO22pOjtX0dGg
dMLxGrqn+/JHcPS95Xwjw74+R2q9LnfL6eKohYHuaGOl9TLgLm6ImCv5SVBSnwsc
chEZqCiUD4YvlAby1mWA+gvm7OJS9zS7qcLW24pJjrhLhm8xVh4iKFz2Z7l8BwXU
XCD+LUBprzl11AuNaEcLZ3aV901qOJPJJfsbcNz5BdL1MLusPJNeM10EosBm5svi
UeJV8rxN+Y5ZwdA/sRsJwi7IC1d7Qr/znbUecuRxe6pWlqkxfkjR8h29mx9N7p8W
Dm9nnRgrtX+LOe5FJ2zqIHP2fu1RLIkcG4DNvY7/LAnOXFYaDcrPQ4wHj1AvAh0L
oeEg6D6IvEXkGBNGhzUQRq6kk2vmar9yzxu6EDvhNRC+gCPfHRBdvVKQ5Z13CtH2
m1VxoytkGFBhrXV88Xc344YO9pWKgMDjrOcoKWbKdufmuwsL+b36nS09EWdJMWYi
9kQj2gYcP0MMLLypVhOosARDg3y9bCMmhhzMCUjM7ZTCbcJdlpokuNlyntkIGzWV
h1/V9piq/KDtL51AJMO7J2CqxCHfyzAZtizEHf1MtTsaEFAhRU+zXfRSBPf6hp/Z
YgrcOm9gvVYIbAEmx1rBG0oeaOLnZSbLDeVhFlU5G2bYfFW71i9syvXB1jTn2P1+
fN9T0QX01Wa/wZ0Tvd9Fh4SK92QeXG60n9ItJrhJ2fKN7A5eU1dAvgiOD+W+w02h
GXYhH+D+mK/RcnbqEj022T0XHoMx97uCLVBZ/ZIU6k27NW3xDmrwfWn9N9Ahra9B
wLC4mhUJzMeZNWuEVBixI+2CEK9JceAQ8wJDD+nqatQjqZLHEjKBWMkp+XDgA3dB
o6rYYx5w9R2ZRr0HMStGfwYugHhknbeWYLuB9A8a3oXbOX7PRI4XXyJbguSNroHD
mmmFoXr8QCvq98DH24cx8DQAinYdDaILxEHSXJmfV1VXzCLFEibTlyRLRtEJoDML
d0w5EGlSGSMoDEcTYghjuLN0bhODOFS5GyOdyDG3bDLttQC/I8wakbT+NQSxaIot
T9wWfqqLfMWoivwCacdrpsqbK2Yx6XVeB1lDbp/+XXg/iwjypNqFGwTznje1YasN
8bMMhURYzPwDTCJE5rczxFUhE7Pb+5kHrKY0hBuQyjoT9fxyZD8C4V7St8z3bTwE
EbgSDhxlOmdsvOTYGMN6pUwUIwFzTMa89nKjxAawu2fnWogvZh5mVIwYX9MqKqih
we6lY0raY8g7w94mxLsveLDtmESjjb5rpPNT8of3qrosObfVBvxGJ3EM5amiETQJ
DdkXY73FguGY6Ew13AO3TIPKskHVRKuMxZHx8tnN1Vp4c13AFYkF18TpCBHSwWP3
VhJRkAMu+WE56XS8t3aOT0nD3RwxIfwMLyBFqRUDDZyZpQbit3e9zqO4J0m77hqo
v+tai1s0b4r3W6MgWFlaKIGp5siSr1FDeatAPd+W2jivOEYtEpp9sJ1wvRPd1A7K
xobZzlx6hU5p64MlnXjDCROPvxmfX73n59aJtc9CVq5+umO+4h760Kn6Vs7Z0cEo
bNRpuuf4yCl1DSqFTk9x3k+zKrdTTHy8aSBzkIRMKVSQDf4RpH2R5L7rsKj6r3Ua
ohKLIS9k84Q0LgzdJwhSBbuRq9LauKOW8uqECOe27BjEnP6Q6RbUKbdGFehT5Xkq
0lvkCbhWfwBq3KitKCLcPVkfxiMXIgsZYvGRRkOyqQ1vZ0oG71iO0+CiHvec5PWw
+4ljS5iW37/xtuP9el1tMoi4pBAADuQVvm1XO+nWnPhr76T9t2Aak4vogo4mfxDC
c6CFZr7DcSeJuboNjkATZ5Zwf2MoGNfIYsYt7o0YTbuwspbcSbmwcOAhfScGO9rR
6xzKavRiSpmnAzwEmefWjjwwu3D/PPE7G2ZHAocwJTu+pmXTEW+ufNwkeOPJZcNd
x+Ms14CPVdFmTa8kNGe0/EN7dr4RpLuPME3KfvH41tGqF8r71J/60SX1mawfrn/p
PnrMQqljKM8rZJdAzcPVnrWKCLiAkwjzisp35sB++Hpt3V1sa0OLLXXkUhRSgHOd
DDIhI0dBlLyMOtA8gbju8rrO/GP5CokdT4CjyZxfSk+sBWyOg+LpBonNDkTX+92A
0XmRPqj5S0tIez7vE0Nj6UZBla43m1WNJs3XSCk7uW0IbHCFJ0Q62wyS+G4OVQYo
NGjDRTOgdXP8hVo2pmtLTsBjx7Gz859+PeKa1fNCHMgnFc8INOZT2f4DcqmEQy4I
f6qguupX6CAK0iyDjQh4B5UX4hyPAaLzEHXdY7/DTGnL3KdXbzTbY0pNUttkAj4g
z2E2C4vSQXte7rvGK+IxIgwa6y4+bL5k+lDKBQz/eI5eJC9n7GzJDPJFxsMrUEKJ
ONkCd5QuLpuq2NNAkumRUGRbG1l/vEQcSKShS58wsqqxKHrYiNyFb3QKIrH4fYzI
Uk2V5HLMITYDXfwSlOhSYkSVJ/e7k0lU6vuWcNDpiZSilTTu8vJH9GI64VTBjA+Z
0J/6FtBqlkN4rP9IrUJQyAFxDHBj1Ga4VLjL9dPW/hlC3/q86T/XxztSqAkR7PWC
GNbCRZa5X8WipxAmzSNDjg60D8O+w3pZj6T4ozz4Hf3IF/uOHWSS5SsW5NNzfANt
FV/zc5Q5kxUw7e+ji+y9kQif5n4JdeB/9EXVmUwYv27gXTZMGP5IvGPk28LBrrVI
dDMRG6W0qgvTIym4MlK0CdV/eZVJ2xVPDZ64yJMwzsv+hNLqb/27eHqaV6kYIJ9q
cGw4/kjnlcdk/A6GorctgQM7UaWiHBG7w+FEDW79fLYJQu4QczubBUd/88z2PPJ/
TVW4YBEzmVHEtEQlAg0T8s9BLAhCcxQvrldLBhP7t3kSeR65LbyoidKe877fJS1Q
RgdWoes/imoPIwSD41WjaRsIiZ+5dMJPSs1DaqFy80ztRM2F3NEeNt5649YXMMgU
EzYdd6B4Is1JNtCI49oK8WVzi2AHW/ZkurKQJuS4n5Lsd3SypxAfMM3XFl2XulRt
lp7qB7WT8Jn3N89v2BN/KtMgxXdbbmn9oHbMEd3vTJ/6tLH8nh5KdIjz5zpcnfy9
6F9r5uCjrgx4DKJvJYwQuXobYOHZVHXoYG0Kh+QYVLoAC63IJ/sMV9DMn4xmlYY6
QgKXgLvs0pj9wBzd/XrR3VWQlPlivK8CStYisLXdFQ1xr6R5zxmuzIsaJleavWSW
JzOcd0vP0G9vzH6RtrJrhsgtn0CJj2KWieOdxNRpLYcw4wneAj3wRMSrouQerBaq
NxXfUakR6Uqn4mBdG/mXHqScbIygR8KyhlDn4I8o4Gg0L5OgixYKitGAInQj0uQg
srO+nopBn6AWNEI7ncE6dKKuJariHd/8DrQjMKp5VWHpg8tqmrMPcwNebEm55qNn
AdKmlSgIYkW3A/RKYfyUit1ztCJz8Dnp3feIH4PCGeANR+ahl8MyFBcWNwDr0MjL
ASGhpEOFyEKD8SAC8BBh/zTxgczgNW6kip3RSTyNrh562TEmG9gFizcYe3549gaZ
l8ecmCnm4C5mNkXCu6Srwkq4qZ4znnM1vQIn/F1Un8gd99zcbcWjP0SAuV8s7pOf
BCmjfcmWS047wREyETTBGNAgI6MdkQi6hRdkltYPV+R3G56vOIOvSH4LqoU1ehGw
LPj+O6D4Qo5VADOLfKPAk6bcgRLvAoNizkkFKaXhXjZdvUQA+waC6YQ2wJxjOK4S
thzYiIgOnz2JSs2f87GS9q13704NrxO8TP1ew1ub8X+PeIL5B+YVlC4RRXLjzNXy
UztsjKEoi29lPdkmDX3pgA65k9X6cI3873fnvWG0+QttS/MZAx9WUmakzSAWudgy
Pie3AGaxuvY3qYMRUNzGtDeHW0PtK2/7pKUWKocLYK8ZfV4u1lGPP6QTUDNyID0l
2YDOaGAPuXdN/3zS0a4jSv2FE5Do8GuAXEXI2XlsLiY7RJIbA0x26S3bMwhESU33
AWNUACfI4K44zETB7Iz5RDJdPrsd66B5N/o5pJEnIivuS/P8EfZLgXxlyxrluGVl
jtKz867/w2tjY5KyI/fRZdfKkpGheY7S+lPIMmuDgMJ/Y9dNR7AaoC8QQCcBvYw3
6Q5K7CEmKhtFulKu+8WbYe074aqr7jNCPCA+Lj3/c8P8e3/ZgVTVuWUzOKNBZA46
SMjbp7EMWyDSDPW2ZUT0QmkQd3dyue0pycM0QYom3vBK5IT1Q8V59UB+DBkkwVOs
aDVOjox57z6FnJ0XJvrZPXfHzzdF3eFQG6c58ph0waBwJK6CeF/rBToKuCFBEsSr
GYuFwZwFYgd2sLZ82QEPg3NJG3tVtrxvEDti07Mu2CvU1nas/JLoNXt6v60iWE0V
iFZ+j8FdCGg6A7946DYrvckYmONrXE//YxdNjD+Azb4PPF9/HQmakUolh9dafziH
hkjAuOejg0pulvxf1Uo8pylRj/kmhqPFK2tkLsIYKXv+zuNoOeZZUiy6WU6WRk0R
Mheqs7OQxaDcCfO+tY8Q7GXn0qI57gra1tCSEPUoefvWS0wY/WJY5laHIMU5T1TL
6NB1XN/1Kvmla6RGUX6xAk16psyYCjXpNf/llXo7tDPQZ/iljqmb+Cr5Ei0wNsOt
Dvy+A9Tf8xdVHYJDpXqSHn+F4IBHZNoAF94nUz2/mi8lGHHe7KeNucCOn7mGmqa5
EkjUggVmSdwNohfJzHuc5oGl7YxfAJJe9CBxxXSlnV9WMdjxr2gNmPDL1UShBTji
ycYkqP7m3acKO1lRFe4t82YrLjcg6D+ygXh59reQCm8n66izSbJlapwcN7Aidfvz
JgoPxY0+29PgeBlHYqz1vXbuZGG04SLRMjbmBRh0bsmdQAa3Q191u/guT4sesAyh
ynEOlxvtsAY0oeIvZ6DS+XHNJSDr8OkGhdvee2bYtPQmqkU0hPhJTV938rC2ROF7
0nKd5ze0e8eM87J+8+prBR6WyMlUVF6WwUgBcuSjlywUlCSKkll8RdcUUST6cBxm
3uOmTIr3zoxEbnP4/fN8rCN3TtClncyUaTGCrVXxkClKda4OV8cr4O5X66lYwNVt
1WoUufC9N2XukBdpaUnBrzNAI83UR4a//mjnaePLn9GG++9LEeWMfqSDVPnBw9v9
m97/9wLnOEeJqw0fJmL2vmQxoiYdqTUCt3iKqNMilx1nnKnnz2UCSJX9BEkGjxIL
WMbXNnFnbXk5xC5hrRAL4Fk5VzGTaxAlJwIc862aPJG7gGlmO4jWYSHHxYpWG//k
4CnPN0j/TGQ6N5oKioggsHI23YfgtP9WAvG/MGC3Mlc6V8QJWEvHo6BFspiC7cqa
ZHawIzHoepEaKAWbeEcMcxUyYUjO7jTjPPMXAloOxBkqm15n2513jKBC/VwzZnN0
byCXycrkCfWOweDz7Zy1lnQuMy8WOfpe7Dls8c/2D5o2JQJZ5Itx0kKnusptoW3x
vuA/PueNFvVo0YnFB7WJJx0LybEQ+SBxSccLNPHz5ZpC3WK+ojpnRpHd5tZZUgdB
8Rfo2YTB6R85znYYKPI4IBLQFIm9vKuZM2doHV7TgAYlABfh6qa3HHZjnhJDjsBi
iPQFmLmQl7+zYq76yL4jaB2ysgWHjtG5XXmTQf0nJwB78tF0jcgRCsvaPK0xrM9C
O3xdJe+VqlzwmGx2bZwAOITsSr/L0Kvz0DIDVPsVTn73pKZ4n/3fNP6DFAcGocm+
ZvSgfKYLu5QTNWCwDPlpUMqn4QfmTKUUj7eSQih50lpOednbm7cFtshrL0JyWO65
BgCmMHVPnb81pDq1jB3A5QIDVIvZ1joTgBARelF2G6Iz5lcAMMWaYnSb8WqJNYpc
kN2iQ4TM7/SrYibzww5Z+NKuDi7NDIuCEifimOkC0Gm8TQ30IKsVb2w/Dn0agc4a
sBayJ9raGytRppAQDXIxFu24TWEYGUFecwPsBcV07kUsP6omw8bA+EfheJRekvl3
rdqICYcWiE9xVQafL0TJKUyXT2sfCHRZMuFh4MG4BjZEBt9+xd8zO7xhe/ymrMrH
shpQqjSX2Fek2NdKX+TnWtH9vx0zrBM1JyRLcwEWIVoSjFvWyoSEvwqywM0wjDfx
RB6PCtwPtA/vBpir5L02HN2rrhKPa0yz/gV2NEaPT7CZxuojTmytVnNOyzsZuIjb
PEgHcHX9XNB7HipAG1bV1La8Lw/A8+FgZrdvWMfourb+uIaDUS9dGEMVftLb4+jv
jAtbsAk7G4rFTXeXmOJUZItoY7VbQOZqvFRRMwRW7Ljs+lCHI0LqOLm2cyBxgY7+
Ihz202b2FC49C+FXvuJPOihQ6a+qlOh6LZFGo69wXb2O3AOM67co4eunSSn8SoGZ
5R+RlOKpifymWkXdoj9JixxnU2lKtWo4/Stq/8XtangZCejJQHXY84uLCLZNPUht
S9J+5P5vbkll2cazB/UwSn6+UmOxROWZLEXXwJtuJgBrdDQsUW+H6bvjgjItoSgm
lBzvLP25zhRBbxCPuuD4QosPqETywvFaG0h5iXxakMhHO8w++9Eq4cEHxQcMkSAL
laYdRJh0a6+VyJknqtTZnVcsUAgyVn137y8k0MQ0tIcL67Dzluhnm3lR2Oa/VUYF
wpvQ8HI/EC6R9hMwIPNXqvulWoQllYvlH7Ng8OVHY7+2D7SmFO/77bp1N8/vPtQL
jgHu40hmf2mpJiZ+RxDD+UgPrlHIDxtagjxWEzsYWAgJOWIdOVaQWOKVPrpkHZPF
84cVEdf5fTkObv/Ff+Jbf1F0i0kjVg422URIyGaq/ivCdtv3yXKoilaEjuAkddMI
+9gJPyaC1dbfCKOZwiVumIpIk9pj9KD7ULRmsO6LG9QW7HkI/2BHGOI9TWpboDjW
XpsaFteHsupPMRc9nlb1Z0T04eXGOeyULOSQnVrmk3BJ1Xkddw05i/qdAep4KYob
bEdX7lod0r9Qt/5+UKxHXffJrwWlIgpfoTb6zU506q0maREuWb4Q0c0CsVxikWcn
xLUnsjLeznGIEZuiHUrhYx95Lnj0nE0mcBr71Lbv/DWgeo8Hl8Jz3lg7P+kh/Gqm
lNBJ52BSVEqoYZH73+onORJHD6AhfiDajQJDSH5MW+55sSbm3IhpPuVR18LICH4b
CMzMxNGNlztw3JjhPzRK6ClYfRTOgb4QMC59gYk+5g7FOqcZGBYl9xAmPsSXpvjY
u4nxXeBqXNMom/uISSS5IqnOfMfnsOPhT81ZNEmPq0TDfT4O0G9uMeTH0lsVBeIn
bhSD57j8iy/FBBcMr1ZEJ5LMzDLPgTpckFOj6qDrj1QpihSlhFdGx1GEv9BnBq1O
7PjTdaqDuHCiOSdvD6hjxxWVuNM3m0CJu88lRkbJksklOVKbKPeHQMfUVtlxjvXC
OZ1a0EqqoXx68EEXDpnRr69aQyC9NbHpJRzZlPwnS1O12ohist+iRMA5aV+yd7oC
2PhLuYst9fsq8PhrL+0z6id9i2Cv9U7PUoMA5tYCA2I1f8jvL743mv0YSSvhcV1b
0COFhQdQfV1kjiibIb1KqS3mU8+2Tzwh+HvA9pahs8fHkqQiV86tETvLvfe56nko
SuAuKcPJshDjaPTrKe2ubr6NOZSPPvYX3fLgYpFKmArvEVY1nhjgSDMt/jNOnNnV
rIOcacLH5LU85WKsxeb8Y4AKWJpiy6h3whHdv+eiTz19tBHOnijzzOx+2mF05fZz
rNXCdOdbI8V1CaxVVOSjSNmtJC6V8GibTloJTKhZRv44iCOw7v//E1P8D7BrMSuT
7Tqn1sJfWep8kcUr1WMlzpDh7MEcSn24jVxGrqdTnQ6sn6Mx0/F3dR6DQFc+dzGL
D8UYk62pSI6UBXSj2Cn6agy+mIB2volUpyBxfeIqQVA+WBgQt5H2+i8guBCdq6x2
0ijfXN+Be1Z8eIDKXipq5+PTWyUrmmZT4zPeoXrDG6D7eQ07ASR1cjWhxceTK0pf
7ldCywR5e0IezUurIPGvmvxYek3Y3EW9TOM60VmtffOlMwgjFoIkafN1BikVlzF4
ai7Yp1Vd7Gk0PP/aXd0520+XvcYbyglQIALiBiFD0aKfcJuWfKjRwJaCHa4TqbbN
zlREDIQsvU4JUqXE2bCAsXF8jM8DhXvskAoIfgBWpbR5GssAixpQ58/9pOydqdoX
67rJ2OkhDAq2SHsxHyPKlG/btZnMZQ6vKoDEQGwa0nWpg/qSgbpX4NzU0BaG/OQf
kSR36trxfaKGxYxmVtXyFbuZSfZ+G1777LR7Dchz5Fk41e7OuU/Si6iao7tN39b0
6nfs5eor6/H4acXONam80Mwg7pZWXvoQbur4x+2kGyrk/lbvf63VG5zL53oAK6EG
VBzhb2yAKIEU+ZA6avYooy4h820yjYp1M88y5MPvOnDDywP9Y9iXqBUOY5mdETC1
af7rZ2KScHHTjJJufdOpcwxQ0USuQhwVUxjXMiUXMYRIVqScgZtdjeomooyv1s9H
3vU2VbkBIHqUkXQyZelyC0flMeInQsqJIBbn4SJWaUiVcEYwPu5n8oBFCTu0RV3s
C62jNNNVECkkPSz+QEvd2Qfcsn3298porjLjfhitF/1QO7fINwckG7myvk8ZbhbQ
7w81QSh+F0skDXUiyu01dZgQ2uwOxhsrA0WnXxQ7puyRugZRidN0VpHKdSbRZGMd
pY+yTvwU9NeWfjEgFefRBxTY/vQovMemXNbtN9lDGOAQfiF9zQNgGLp/O769Mpwj
STzVFk9j2otNPSoiIN8PnUaIQ1vgLpzbRxiMBRQWahUOBZcnSsR9r8FYfzrfK6U4
gq9HO2c2HYEMvCxXEoHqydR4VuP6TiIRxwW0SJySPJOr7pkW8zDy7Dp1Xl6Dtecl
QDOoQ6BJ97neegi+7sOT40Lb876Tr3E/qw0mvBfOsu7b2P7GRNogjWS0bpQUCCaW
+jE40TX1UbKiTAmcOIeaY/dmSz6Qy/KLL50gIBBGlzq3x2vwshVcSqGLDggeO/gm
GFG5SXSiRQgQj6kQHvH/pi0S844FPAo+tLTK4ni+UKEWGTdLxu2d+YnMgzyalwUV
Ah2I8m6r3NHdmganC7XzOK2IQsKQpoFjNaswiy3Cw4dRGAGdlHcMRqwloBYCNpL7
wt/RF+VfsPmcNuSgY91vzqvdwtkHGcGoE1T9OP2wPQL5d7xg+WlEmwGUq9Ps2rqZ
wk/dY1wigvlaIzDmBCT6kI9Z8D8kM76Y13R5btl5KOSbd+EFs/w92P5zri/cDiyP
FUKdHTSuuqXl75YT3vDfGfm0Uwlq5R680pN4RerlFz7Ik48qND/oikgBPjjS5RWY
xTwDMpg0Kp826FhyIjV2EuH8KiKlRp3PaP4D0JQG9AZo8sZG+CGW7R0UAZiVMNco
SRG95POP3TuhIWFm+gyalueDyLm0aYopXqoR7H4cQ0WP73Ie/7M8R32eZnF8VJEy
uYeKGKMs6AhI7T7xEo9+U7p9xbZXbybYmiK46MNPrD4o3VzQsA7i3jtqVZ/3YsyL
i0rY4nSStKCnlbKEthX5/Sa5UjQmZXiawDOjgwY9ytqYa4p1I9qkumV3Z1Iwcc9D
PCKRhIojyNdkxI+ZxmgFvDO+UJM2a/J+8ZgKn8e49PbsxPK7FGyh+RiDDQntMRxV
Lo+UGDBSZ+9i81KMHzakkD8ApwsSN2voGZ+2EuhrVKxIbe4MAgd6t8gZ7YVx/Qr/
SoPhQRv5wE780vwW5VgoyxAetR6RLpnU8B+9O8SJSBI73pwc8CwEggmM9jP7fFrr
y2eq5Zki8/T21Q3lKQTB1WA5sNN/CGmPv4fJxv16bb7Aix4/Ft5pcu1K0/dzfWcZ
9OLARrB8c8ghIxNK5M0vMheqkNfkq8e6gfeGcaX2GCXIpqSO7cXquqqFNLX2CETG
to5r2ipwW6FaTRJRAlDnO8DCPYNqkfKmHPQESPIGThiUVkxud3aIDifhQA6thyZk
UeZ9aU1NCUqgKoctnak+u7f3gG4VCh6qa6EoMIHkVcyjx/MM7P8pvLwgcEa8wd4O
TdI4SuylNadh03lhRANy+4LTuYVCQmGnRv2bOND6D4oHs7s4OfVrlWuvgA8HUNQP
X+INhkbTPSnvVx4q8p0qVMCeGh3G5MHyzxs2Eza+YUQ6RuU96V601Cr2hwCKu/P0
oz0vJocbevDvQZkGtWY0vZUiSWQM6ONT+d7E4G9nlu+DF5epFdZBGv1+ezuxW9wh
v8GI1UVvxCy+NjI9pusfw4BBBLMqU+O6CbgyDES8UVknGeexPetYb2kAyXcm8c11
r5hMuBBWDGvWnQwP4YyopYoy9RWcDs4BssPPyBrO2ZdK9TBsuUJY8Mb9A7G0WwPd
eck3AdN/QpRIY6AH+2Jg+wyc9EGGp7lb+6CV/b3jI6oG1Oo3UnXODGztSxyBGY+T
8azOcq5uw6xZjPEFpa4jcVjGf5hkln1WQfnRhWzhpG1ajqNrHDUHyE3KXLnQocgB
eTm6FdClplooySHtBE7KS98P2BZHz1Kx2HMHh+Cvfi02NhW4vqgvu+081OL3ZLZG
1x9hFzVJwmuPAeWvhJcM7YJCUd0w2fqQjXKdziI4aVBMb4/OCWvjm8hHKEIkpDrD
+gPxav2fS91/b5fxP5gnAmdwqleXP+TaerEQid5JIgjRpDEn4VXm+ryWjzjB5kGO
b/voJ8+UqEhozpTHS+nv3JHVcwpBPL0gYpticByf+bhzvInvMQdNMomdxMMjBK4C
GRohz9nZmhc51q1tA++ZufHxvUZ6LTSNn+P/pKUEPf+I2MJNPiB7rR6PGB4xuehb
MHbATrK8HLNvFujbZln7Fd522bphXXN8ElvCvyUhCBa18vse6wFZrd9EqhKjXTTr
TRyFDMi/CIuH7+kSCQUF+nPx8M+RMBK5sq4aVqJWfUX84V345h4ooiEl82W4GfNh
N1odXEmRZ1YmFkdRv3XY1UyGyQxpeb2QxdYDTAwJCW5W3Q+rBONwvru9iwPT3CEj
DnksLjSDF30N70gIdEqm4NH/WOESR5xPl8Cn8pHgv8SPnxwdKQEEAfAFiFrvTjB5
cba2qwVEP6RFt2n2T0FmAa9nsmc7kbBx4W1ujTnNBBlqFdiJcjq9xydubH9AhB7k
+l7twpSO5G8Ta+9EupgUhOjmBSKrgkzjqptYbPHbznsCwTZoV3xsINV1gt86nUhN
NJyk/nJkx5vOYLhO3sb4z1MhnXA7bRbqsvVQedzxtmArzHUEIOHgm8C+l+Ia/5Bf
nRLef4pcREKfP1Xe9CdS4Pni1Emo9sGT6V3LNCrumazeoQmkKu1HM+Yx4UC8qMRO
dJP5YCJLjUG5PoNL4ZWyV4IX8naiB7LmhJ48Giq3a2sbiBE7kqB9u1Q0odNm8lwe
6b1B8dotrYKQ77yj4VbuGmzxQEuTdwl50rq+DO9urE5HifEFuGCOuHA3LoilrkOj
l8wdUnBsugFhOw1WX3wzH9APFqOc+FC4gSMBfC4FlzZ2ZrdSf8tLr4A66IDMg0u1
70W+Qru6XIMTtCESBuWjEmJ5ZRx816p83qivN6WVZGOfzh5pT9TmTYKRvGRx+svV
lzYNsM2nPioiGifLzHAE3vWV/xaSVAW8iBc6SKMdb6myKDixxUNCjGFd8Rbq2XMB
w5y/SqpPS4kK2os/mjS5f2Pvhb32cZjAbrnAw7QUsO+EabIjHshiu+0hyjoTrdU/
K6G02Awx0CgRXdDajEI2m0UXvxwLgMcLPdeSdUkF6cayq56NcIT+hUxJ0l/KJ3k+
+IlapqLyQZlpT8f6DpRuX4iJgaeSqXgVV4DAGg496JDBhdGDF1ZlFf2ICZsMuWek
sjFuCbkoAJFvfjNPuk84ToDAWOe3c4Y9x857ZSWg//Ecd0/0ANbqg3MNTI6Ko+yE
o+anMxRmrlKlyWxcEGGo3O8ZDh0XNk4Hr3e+akr1jYDQVSadSEV6alZcOx+6Kq1t
zxinMLgH2Y54APWGNGZO4MEXx8MTHoAa3ek1wq9SV2diFEPnRRSUJcPWhFxVO0fw
2XXU5tcQ4ACIlbhNuFapBOrHKJQ+ToyC3SQ7HvbBUDd7DXrd3xOvTDORSFxTThkg
sBfjs+TrWdPJza9TeBCvAI/MWZQS6lBZdqoDuQ7pwlfiBqROI6ku8Eu9jhAYs5Wi
QcNnRxvQNA1TDpWTiAuP1Q56OEKD4P4SF8UeA78YMSPOaZ6jez63tNI/aDCG690V
DLDoKYq9wCPtlmEnl2dKGNgPe8dmmr6BdHpslEMH1M3fxnKB7zemi1Bq2d8i4DTC
lQuQxPn4fLen/M2QkzkIDkvYs2BM2Ep3fOKK4qeYSG4d7+HLt9Y8xIyNOoGLHbPs
4ORfk8M/pUkWwa0dlNpIO+f5AJ6Yss2kbT9s9I5JZzUf4u1ikOT3w2+XhXZp3l8g
/J1XPALRdipkJU7aaxQ+ahIltC6nZpqpD/DS7gMT8YVCwdgPQBNaynnqmksfrdAH
L/aVd8goiPXULjpHWsEQgdA6zKWl6e4Jto2nCiAVk6FZ+V2ZPCkH6240NBDL57Sk
zeVOhzNuQM1jC4B6d5ocGd9R/L6Ql546dePbcFITm7Xd1NicKBXhjX77i6jd2BJ6
mOg9M9rkJQWEij9Mzf6JLuVp+eonY59ZPHizDMRiiQ13uRp1dJPNIklTpUy+yRgX
ijq2KQrcQzTpI3bRWUdUwNZcBcknJYCJfCkDUyJREGMI4FH52zRYOC0Wgh6k/9M4
+4vNUqJhAeqQZnh2IZ+raaH5SajEUHByCEuWLQOp3SHSYxHpKhIT48XkBp1MJ8C3
L0d8jt42sN2CRismIhSrfj7uGrrc6yrvuo6poF22BWUWZ2sGyFJP7Q3VQ/dedh3k
DvOxZVhhKt9u20XYgxaboaj/W+AuldgmZQfTk7bSgFXOULUjumqO9vJa4VrkNtkn
G2dNYRrK4bnHcwuwbLu6cLwIGpFskCL1e6skmRMwJyd1t3+cDec3VoDNQFUcIZNd
volN6C2OZN03Dp66IHxTrLV3T0lNYWnhZxhKGwLJx3Q5Mn8QWqD3jjA2Q+FmHqp1
KNL8V7KKWKZlSzvtKWfcfjyl3wCK+knRxhGoxpGmX26a242ZHKFKtf62GgFVrk28
WBks1Xe/3G53UaI19PZWaq9tm/rmdJT7uw2d4wFU7Dl513+qp2rCs5FsdjG5/siB
W5Xz2jAv4h9OhFB4Hdo+Z6mMTHGyXgbOoi98xFzOQdE+DHZrAstBxsX4/HJzE/qT
89VNQrzOkjquwzFgqWZQnGr/sCshTNenlc8RwZ6fYO1DIKAe84roKao3DLnK4Igg
4lGwBiyiKVX/5umpg41xB6t9oJHN11qXW3js4jiXDQODYhg0PAo+aSvltlGCBABP
ksT/OSdZWmZEbBFWotMgIhP6jhI8t+IK8OKzXp3KKv7/PDzVMfm3hxYnUV9lhzzJ
Dj6oOjLQXFq6/2pzQYjQUz7G1r1cXlWF1jpx18gdOy+pA9LYSl7IPNiqfLSHkkfk
22P5aOVEobGGhFaY3X1orq+PHN/nF9wKFeIi3lgMV3mNO63eOJds68gnXr+fq6Gi
z166VzQWHyWwixHmQ0NSFIujzDM8WOmQLy01kaOCLYl5ttpwDxoZFVPg7WwTRW6J
feePLZy2oydsSkTXEHo3SWS5Bcf/bVZ9C6xZXSAVldiTQcNC/2BvUAcdI8L/zCYA
1ErEMQJ+7jyF2Jc9FgTfgFBsOdcszTHihwAF4UqNngOqRq3UTRB0h6OwTPaJzHBd
XngShZdTwrDre/22eBLEoewSv4lDafHtIdKbDTuyxrs824/tKszIrh6cC/Jhr2+V
OjUG0Tzfv9t9U30uAHIY0jtkALjYYzv6Jd3pnjqlRRKeQBrolY63FiToZe6ZxBCn
K5qDeQIpLXop9BykMy2PnQOV1dbz/2OSkLi28DxQoEc+sRci+qqyaClrIlCh3qBQ
2s6RHXuCS4XtbZ1VsoQd5OqQxIAQJLmKYXfes46J2Ly4xge3wmFKyvypPS5pqhae
9JEFQgO1hZqPVBIQZXIvIkHAYVHsDHUZgx1DEPS81EETR01nGkd4mYkfVSk07rzE
PtV98KEU3j/baBIn/GTBi/ZCS+igbqetu3foROlhowJ3hBklCXmCaoaoNiTUlTZV
b7QUUQfG/YQ3OYGRBh2qDMLEq6w21vN47/ObuV9UfCx73io7FujJOQyk0cS35OO+
unAoMKfcoLsVcUpJ4es/nVoE1Ucs1w0eo6LMdhyN9MxXKMe5POII3weqwFQHOSwO
wrKCB+hUfTy5T4UVN8+YVdxep/RQJYY7KTkQ+tanljHPpA9fk4b4uAWCY/VtpVB3
RBmMliVPQmE4AsiNutcCWA2wRsLUcHCnj/MRPWi9pMcuAylZyiiVpkD1tY1JMlWa
C6zp2nGS5fbz6UC0VlJcLZ+CcCs7LpdsPxOcBmZsfeGk40hvVEGnKFl+6AFg01lP
fkR0gJJMzdiAITwTDyqktmE40jngXdZ43btj2mSuTyQNYtwjdNHtEWquPUt3s8d2
ym+gir75SLdmIuZspUN+rfpfJBdT7M+iLS/dVqDL3/fRdpotSJvF4wYxKoegbQ+i
trqkL7XfZcMWqdCdNGh06+EXmqv2VFT+syBDYjKZuF0IQ/3X/DjMHHdO0hQIZCnr
o+QPRplgQjBWdYDSAkeQ0eGWi4kF1qPeSU4PVYRCI07O+oBMrZ6fmE3HiGg7h4kJ
emGxc3gJKN+YAGwicHY+1nLxKunwSNMvILRYJJuUI0Dsk7LjCnBDbLghVJvV52DI
tZkeR0fIbZipkwVQR9hNsK3nCJEinrG3Oo6HADfz0/rDuapxFAidvlVGgpiXiJnI
xnzkbx58D5C6P3pQWhirXvbrHTPAT4L3XHojUB/oty6g/fCluOYmql/i8nCIl3hz
StpVG8OtfGx34IWgdwCRgQn3MkBOkVhfpAbOhkx/1mfZyGh+wh+xpxuH0M8tA1zD
kGCBe7paTddV5V7D4vQnagb5jLGSi4uHgodS6IHu4BgwG46gzp/p6FrAcuB/mJO5
LgjSaFLj78Nd3wJXW4TvvGK/6z1K8IDRD8t5KYyq6RzkfTOgBQoPbgX4tSBeusHJ
8DH6L3eYvilKrF8N7844Au9PNVRI0zfxxJqrs6vFzCK8IYCHD6qBIGzQt0JUQRKH
mX0JoRqFx56aftHI1q5XIAay4ygJHJX2KMlGDi9ruJgzLpnWnbFSMoBaZG3Iort7
GgdJON68bPOaZcj24JsUoBOld4ZYPB07LeF6OiaqV208FnW09MXpugjlRDG2wBnA
3nFECOph3DzpMYv1jfMW8+KB6u4tZrPczSE0SR9FhEO0lBrHFQaxOFVbTC82lKL4
2cc3mXmISYbSfVAh9W8JrAdWHIxtM3lNE9jFmuzt4+NPWD9Z7quOcJ1Mut65FUj7
jZlGKwc21I2gfkQn81Cqpp8Vc5HvFIPWo07h0Axm91HlAADg84w9UMUUo/I5xfvx
0kgelxxf7thLpySPJJviDO1ZGlsoRWy4X/Y3I5di1aajWfzG9cWvR6vhh05TcFSd
SnOxj9lLbMx+u9TwkOMJEJ9VgGcEdNMI64UeIzqesE0DGf0QP6KPZKzwmJpoM+5u
cMS7ceK5ltd04FSWtj/GABO0DTbrrRU0aaS+wAASwk9C+/EbMXVQy+K6ojlVOiXB
uPKBRqG5ZPj2uo32BttNU5qbDbS+FFmWZcvirl49vC20m76LHCBCF3vxkKe6wA98
qs79hxRl9E5hG0tCeT5EMC1Lku4IhSQpEQ2ar8bIXPYLZafWz0ETGMflVauPyZ6N
N6whBeG5V5GgAZdsUwJYevvMayVcCjkUetjLSUbd30joeXTFQjxUuDuRRnhA1+Ob
230EDNGSP26blYnDnXZ455qh1wtnOLOhsp9HUEa6XGa7OymAVB6Y95r20LEfQnwK
33TcSWKndGiMIDamrTeanQB0JZ/HIP6OmFR1tLGQ0+4Z1nrcaFLTGIqBG+cPAitJ
vgfH5LUL/w7aAyIed+UkDmqLpl88ubXrUYZtGt/N0RsOdZEdsnXzRVGeN0E4UNK2
gTN5KMzyPyFdIYWUQFqV4O+zrnic+GYVytPKANyGRNlU7auwHu0cn+PdD80Pb9AB
gOvmDckBd68tvH3Vrho671az5+5d3uxofwf1TwW9+P/q+p6A24qiEHzrLJIfaSMB
dLdCBwCfnHkP56rz8W+KQRFMnBItX8j4VCgI7/VARUZZob9csrygy7veQiEcAkun
xJdPHGj7wp5ui8mAmuF8J8nx34RIBGbDS5PJQv9yAoFBoO6T9ggJVWI3Oj9t5xpd
V40Vy5xkqdqiWEMIZIYT5x1t8Fv0JYYS/Z98ZBRx8XqdRkQaQP/AsqVrzEgdxc+Z
+VOrbJyPm83MgJhLxhIP71yak5ik24WZqf7IOuxiIxfnIvooIxykweDIZelg/GuY
FpcSw/nNhxcrnVUYBoitB+jjvqEliOdoaExX9CVmkodxmoY8JjaYZj3euo5ST+NG
Mj3fHwwFWm1lU2Suo81J++EOqlK99cPhSQfaR9+0czoflYgh8AZmLYaMuUfcQI5h
ql2Ocva44MH4eXIwRH/jvLXphDWKKeP97HoGcGxrEc9HvZjIPyE6Y+o1S0W0uQkU
crVLodsx99BCqKiUNgK0RFZzYldMoz7Z+20/pNGdUfPI19t80FqE7BKAab7I11QV
FO73mZoIAqqLTSArlgVUDIHwd8iKC74CRl3GGwZ+HlbaxaEpVZyW7Qq965mZmCjn
fHuoBQJPuZIxkswJfvi/kIDx6NGn13CBBjICpWf/zPIyhg0ScflsaWli/NLbdKDG
W56gf3Sji82xlNW3R++QZ/BmyKqfOVl3xB6eKo9TDBU00an0z32vJ3dSznT11eRZ
5wkCnCzGHdcVFLOw/XsI5PoLT7GYpDlFeGMKlLNE+mN/qO5OfiFHSU9OEO+Bt6fg
xlnxM9+2mE51KSXwZ1X9MFNdwIw0JX34Q35o2OO7Y3ueD8WiYjp0Mz/6q1T2KoTf
czdrZ3ib4dOVggqU4Bb6nmQVljw8Gaea84MQoM8YckQar5DN4FALO2AzEsempOiv
VUoXrBIX2g8cUXoCO8mlMjedzlBa+yor7goEYviZ/OyUmUd9BgKVJd6barJKWy65
ktnj0otIW7Csl95UNYGJE5wamK3/rQcxv59gUH6Zvj0DsbHdzwehbc/aKC35UIWI
Ke8lnDvzGB0ujIE0c4KNSfscgedgfWEby/EvPltNGHG+BAQTMxRbq11E60ijiete
WSczrmRyW5QOkoLlyFqejI96hfazDnegjcfUPcmlV7Fwv7SVH2peWb7I83NO+Agw
Z0ZCfLCRm0J8yl7SKG1LFN7m01NboOl89In9AuCpmxDmUdC7X75i3uUTA4hU6Z0E
dRXYcomtw/6mBskh05QCC2wTwbwz74U9p4GPwzRsh2M1ECqvoVaevSK4rJVi+xe0
UZwIS02Brsnz5TztdqjgZ6y1RVi4MA3KaPBd74GFED7Qa90Suo1p+R2Fc04gGytu
dI2zuSOASOce51IdQDbIyy0NAeY6swjrsM9TB807GG9Y4bC4tfkLPjZZBWNr+rdA
+VCCG+F6b7FWtN1hLsSqC/zs8Hvj4wlUtmdXtzHf3CTL65ZGuzlMR1oVb8uJPSC7
YKWLw9sBE4CRczQ7UNNdyBbUeiJdwt0UrEKC5sPrSu6StOq5R/mMMVXyX5bHTujw
sts8kxtWWOOR3YpY6J0nHPPEKOUOCHsZV2tTgmCArI8rK6EtyraQHX8iD3b2hWpm
A7mJ+IFwlv+sESMZ43/0NWbTIcCxwBHE9ttQfOruh0xuIRzbmyWdo0OtZkyn7sSz
ZM0MAcGywWahHF1xpmLN2kLtqaQ/6BgwA6R/ufFSiQJ4p31G1NFS5cWQH/Brgcz+
IoANp2moNkTNpsTQ6hoZ/CaeCeQ6PVSYi90Mu6qqmv9/EJjqnWmNk27flQEm9YYW
+gaR3bhxRRv0XJOESB2N0hUaposzpzyXuRJm2K6qT2G0nbPy9tRoqcEhte6xoWWw
tvrMMLPtWlgN7iwi48tmGulPii+Hn915JxM1Mvg7Btdh5SXln8Nigg3VU09ACEQD
o++rQ90aw9Mk2mDb/a9N4vir/OWS2dYCbdxJ/yt8d+5jQzeccVx7SVlBhmJNjcaT
VlAnSGDXfvqdSPuxpslsCEjg1oDbFHygskVU+q8ugMXQgKVGsbIHJZpFr/prpwsj
EurQFWCRfob8LivgmP3NQKY3eHKquI/o0FqlzqRVqluiVrSP+SBhOjWw0KDRvj6n
vxVfFmRohZ4mEA/hGTvlicoMpl6BqTcvp8F9Q1WyGhabqqzrtuRGv/VJWXw4bzrR
dNby9CDyOFeGxSKgFPXRFN2ja/lAWa3otn9tSbyIjCiNmzkK7zTNec9PZ8bXY5fU
RbzghZC16WbscnjkCkD+t2XfMpvMJagxduOAdVFz/oHiTXM/XMZfrtBY1FEY0sbv
dPaxRmsg7XW8gAvOvkt6qlG0tdnuOyxQSMOJJHEB7h2NloYSzXNr3QVJrzP4CQia
VFPWAWIl8O2fcWMiG48HIYMjKsuFxfnyV3EIuBn0gcR1s5B/uikaf6+dpke7QEji
U28q+gqo07qwiLP16KdNYxtCbLn9Tlk8472bo/8w4vnIu8H1FeHLXWrmqsZWQE41
Ke4ZmwWKEBEG6KaAhRTAIPQKjwFJOMJnBrvs7ew4WVRCz4Fqm9UenfzU2bbGGoZ6
DppLUx4MCiej5lLUWhgukLzLO5f0ZPv+v9AlESh1d9JtIvF3hb+6uA1VAkUa1nJ0
5zoV3SzEKUq+paC9NL5UfTo3m1BOgXITGQ1oIeEryhK80MTdmNLgM0+TpFLjtLT4
g6JJ9WV9LwRzUOibiQ00TtFKNs8mTCO+rziiCA+UzWPU/f8LXkg9KgB7kp+l/W/U
1s4fzfutj60TL/Fz9FpPGF5BNUVfNS84SsGuejr8ixChdF7CQC7i+jXK9x8peVGo
6c9paWT+TRNSspX6C1oHW43Pz5ML5SodQa0NiocQV/7G48QWBQuAJjPV87e1uCh2
BFKeelDOwmnThboMblG0UhZSGbmjdmPM2RkcgH/OQnpAU8VvNqbJxXQBvbR63LMB
yJd8/WHvDeiqmcsjgzu1TuWnuYGH5lQAgWYCH/qMpEiYKVcwcowyidcAnSxkU7T2
5KBPy0E8WxcNF/sSv5xoOXfGdVUiBNxbpT31IiDLn4R7FDpGGQWPTqw3spfLK1kw
2+4csS2dtiWBiNy1jYfkELNZ9iQ4CCYNz9iEEPkH1tgfUouIbU7phfMt1/2RRLAl
zkt0h+M50oIqN+X1wpwehdQJMYAufAUTLVjJR2gk9LkEEyZtSoLBy6CIqc+Ufa4q
Kp08mUSG+VeC8E05bE/b6+VoV9G+borAmWUlDfeK5BpfyebcR90V/dVpKpn8ph7T
xtwlwfBEAjz4UUJSr+yCch1tUzzYcNrKvjfpFOavv7MB0UfpQhi4TQ6YU5FcUpSx
60brqpxEx6w8m9OkMTmY8PmhJHc20g5rSwuWjFJGq2y/PSZo5FcukDmmtidpL5+Q
O++l7WsgEcBKQhrnFkw4eMVLGIvbz9Rn52JLfDvtMqlXeHytChE/w08ez8NP6jkL
P0ayn9SYC1Cu3sJTumwf4FLJxFJ7Pj6jBRylgs4kour3QXwWkDkGy1eRJSn2g3B6
4SUQ4p04uQK7NGpWAzTHN72aGUShCLWrPzl9PFkYzbPby44t6f78FyxZe1pSeZiy
K+pRpvLy+yLLKKZMvCiNpnORYsM2enSNiKppLgxz/QqUMTtdteEeymRbGKuCCmLk
ooEAx1oGUw59kBQ6Yp12H42a5xSXI+6FYKtgpy5OT3HvVun86HcxjyWGcGFbwv1a
11YCTCiZaeKTxh9Z8OduJH8dvgBPQywsZifBrLfzgJWzzBp1zvsoAezqChc7YVuE
nM+fzpfGwQWGBYwl6q/+xDZ1lN17WatOZSgNZNTO/JMHKAKVBRPbA3QcVS5vwPsc
NqkeJDsZivYOa40AL68pbmSp+3U9FeyXMZ66sgBDhvoPRDHSMPN1BwJuCVcVMQ1b
Q6BZNxocW74P4RuEUZebJGXlUPs6xwJDjeRD6Na8EeNIGawAVfzfqKYWZQspKpg5
77mM0x0HuBFEbIT2rGntyoih7qExSFfJL40W23v2xP2xH3kZ3bof/L/DkWiMNWzY
roMUykjKyZA2FGC2KS8/DO6nFnlBp0LrSBnmpNW06tnfhfzxaI+L/SkUudqbs4je
L0FHFv20zVulnnw056KhjevHm3aWqD5/amPZJKAYA3N4N9SOXJEQLKq9s2GzGZW4
UdkYs3l5sSprNSvjxuChhzChAMlQ+p1llldhfTBbVN/QkhWWcu8uF4h8cZbFICB3
wMsOBpVtKN38YZj71gcrbn6QS2qPMMeppfWTo4cei2NvtT7IRCbtGRHq1pwoG9nD
zBoV/YSFZv8DrMZv9gYlh8SpNGEUnUUROn/cEX/HF4oV/aMx37oRclQY8WIOUKe/
3CmcfUKrdt0CnVQxVKklGNOjrgEWUzHG3xb3D8hAWXXLixAD1VP7gj8w77KEbSl2
YUAE4PlxYzKkD9HREIleNeVcZ7ztbyLOuv56QJRo40Rnn44Hs3i5UXh5lkAr/flw
y3I6lorPeKZhD+ztdR494webx+ydPDb6b1+cmB4VQVIH1Ce3ng8X3PZQejwL3d77
FtRxYws/mtQTMW64dct3veYwIzF+7kiTYRBuyToY9OwwbU0WqTdE3iOA6ytmBQY5
PCwFI/UutS3CsfzPLfYvemU+7D/2K7f1bssIQIx7/Ap+a/YO0IfstSTKi13p9Hdl
tgTerI+FtxjdbT/XeauPTemkpRgZSu3TXoZyv5YgQWLLyVaNwJ+AdidBfcwtWqjt
q243PkGVzVCdTtgLIKifp+7uELMVjXr26mWYVPpLLhfP5dPItqUu5zLBgI2cXWhU
1didJV7Xx/0DEuaLBqURAh1sKfOLdqnry8xibD9XRniWa3KxcJmo1SmfIns06u0l
w71gJ/DcKRUD+ksA2qrohFrrwOEK6KnAVTaUJIFej4pn1NO0LE1ujGkbuiEA8lr3
9OjzYO/rDCJeAbu//wtBJuwRjyJZK7gE0yffBydvnCLu16rL0qmFWUWGEy6+IFT1
UiBznDcI7qPeKblm6xY4kjw/Tp9PIH1RiY/tQiJl2i3YoSAxd0jUGhmtWuVIX2CF
7edVWZnbnJvU2Zk4mvBBIljH+8SHc8xqD9WJ+vvuqQMFJRyPBieBvKyK9AihfbtZ
5Rxsb90EE71rDexyBqH8NUyUoWTz3NcSdUyknFCN3/2fYbtN2ZvLefftu/jfv1Ni
S/vf/GaHivAEcusu2iPl4gbA8+86jRiCJ55pIxiBzYbU5ytZ2u/kzc+mkeI51/bU
FRONKhmY4Z17fty9RBNl6njJZ9incXcf/Y/tAjWU9iArd61lZ/plTm0ITdh4h9dA
JPWv98xlgiZzVgvRyqxNQdAosZ45TbpZ/N8BVo9fWpYPX2ios0wqh2VcdnCGYmFc
4VwC3vM20sJfabHEEVtbq56M9JUW3A7+zWyjk8tC0rCYvGbgpK9vpQ7c2mbR4AaV
P3L4wZrG9RJt+ihuFdpYkIHT8gy18+QAvWz9AX+6oBqfJK44kKqzMU+kvGuhcOhm
e61+DIuPq4csho7MHs341U8qe2F9oT4nJ5IgCpAAoa7+mVRPcYUgW8H+603Enfq9
gIU5KDtgzM4ypGEYCUKqnexFIsGkwJWAr0+3LypUMohVilYnhhkubs4O/sysGMAj
8CyGt0cDAb4tUrRQONfPQgXRsdNIzMiicn/05aR2jID9hjqeRgacs4ZBUuemcAK+
6IABZbKYjYs4K5bP2UDItVXvbnRf9kV+JwrlWHsczMIAQmXoFBbxHVkUVOdLTdNz
wJRP6/tGzXrAGmpPdf6qtE/qbOQy7NwQwVwsJ9R5+3FQOA0sQ9Qd6UixWcN62tD1
hUf/5GlJGnqOqokAvp2zVv47Bj8MUIHX8UCiSGTRqPezs8Ce0zcnX+xfuF38h431
j90lb4jd8nWy3ES2IpCCS1LCvhI0v5X3oOjgDwmB8StwSHFWd5w4fcKLbgarl9LZ
WB9IsviZYq3u9ghB51g4QoYe3c7SF4kqCgTPrUi/x6oHmLnw+/RkFS6ujRPv0Fs+
Z3n2Jk7cqxL+0LvBYz8COGFU66LUCXplwxLrBTRcmb+k4HDFKqfsMtaCosFzU++w
FhUOZTXa9F8SVtM+P1+3unUIc27dkDYAwk+VBKPu5Bn5pg7cq+/3Rgw2iSVugQ64
XfuIlQnxCuVIlQ+ri7jRxEabSMABOaf4mMkW+Iwu77PlMVBg6clyBW1jYdMWJ9WN
LpmOHv9UL3rs7TjGwbEz719hzquDb4Dx7QEdXmsuZYMdQyDlFn5MGXuAbHFrWhB2
FCQP20JGK/2DEN5lRVsLT/PyOzJYga7j6pObnOEr+WdYEeVzm0167w1u44U1eCtt
Dz/fyDro8ECERF6ij90QRBa9FNPqQ72SZXbozCBgJoA+aqSSXgB4pBc1PXc6lx7C
SUOplXVUfwwExvTUArl7itAj35BCbhpbyvizsius4zghbKJo1tYMJlGdOv/asXuK
2eed7430vyXtvE455Xaf3hcpa4119SiVnMJVfwEuyX4bdE7F+jW4q1a/5uvWcQy2
1vBY31DLaLvx4gkNu3cJB3oEPhW9Vjp7oXi8RFaCpD1CB9a9HiFl14tlvTG+3iXF
CGe0hgMyKFWAAXKBY6AFNzlcZ94WLaxkXiB45xVGplB5qlHCwyN6ZWj21j+o2t9c
hAZ2SLaN7wCqHdU95/FWl1iOfq3go/oJaCTRPkJKHqYRb3h+CHuJIWrqjp6O3aWU
VkPwyBMLtoVmtH7Frc2j3+1jPFErQCmTbqOTypndmwLSoucoj0qrALtOaqgbua+h
UrHKDL0o1KLCv57m/ok2OM/QyMnNqMJ9OcAXU4JpPGE4l4SuTa/3Amsb8Qu1EXO2
oVuOAb4SQNiVZ5oJMnNNi2/3Yf8foZry7IvVFOk/mUJh4bMgbXvbi7JoEWDbE23U
Ml06nej5BrUxcs4Uwchp6/1sjwLwLEYxqfNHrF9RczGvH/exhYs/fj8V02B61Oxi
eBQZVrCtFKrXxxJv1sAZKr1R/4uwMs6ewOUBsuxaTkSgdDLstxRhlh1CdOVR4Y3I
smLPBepWX/hvgYXBzDQPhJ0VeIbREu2EiaeNM8OpSosxqhAg+B+Jll+2/8mGa2Gz
TcrIpQgDs3de/OKrP6vr4lBPgS5MAdWo5ECya7Dpuzp83ebN0eouimjLK5p3nbou
lb/Qmn6XCyoD8uBatRavvq14QvnqtfDSC3OBvdTwDW5CEfyK5Oqj0YfoAmoVgSCA
Rj33RGZ+cv9am9ImZsPmhlb2xMW+jtDT+cBQ0VdtYooGB6AxE7CbIpqX394CDly2
rk6dxOV0xz7y8zf+VH8sFmgvMsdJmLO/dW4/Q32RV8JcQxQQUyrur9p9idt34RNw
PHWhWgMrxVQqJQVa3oUrXa05kpPf3avIgOInjXd8ygmFzMWrYPKYaKYN9g54Y15X
waiOrw93MfBIfniBCDmIrEZ9tSzdwu7AegwKJXklMSoDBaSMnuWYXN9Pl5p/9h70
ikuPz4d2n8ofBTHLSCx9+ALjehuIasKAZyc086iSikAEaJXgXZd9RgC/WM3EngeH
N7pkSl2ly+3sVTobykFAHFH0vGWFjsabR+m3IfypHuu8l7r0jhUkdvJrt4aJ6aCM
3OIVvnCpr8naK9FZmswVjiXZHJk/RKL2hU0hmA1YppM/6udIr8JA2a/ttuYENXzy
wTCVOOegCStPNBIZqb1LXGh7rJobupCjhuKtqqhEh6y98K+fIt1QIQ0wKCxdpdxm
8geHzBQg/v/TG2Q3xn0y101SNIM1orFBTPgjrsxBKNWR5m2VPVxu8hQz/ymvxn0G
I2SqWxRZhiANCHXqik/PYT8jofS+rwEp0BPpybkMJhm2vI4D9xgLkiqaYEXIOEnG
bgBPlS+pGIqOr7kjOLI/BG+ezA4F1Oi5Q44ttc0yNoPrYzS8cEBg6em8UWqDTUQT
IldWJWIf/yEMYW1nbW+KcJDznAmzEefMM+0w011qIbntIyEMJ5qRHSHS6vQtNr2a
Hgl1bga6M8wtdvScjgKJHywt1kId3JfZRPPsuWsg9Bf30Ziqfyrig+wjIFWHdwed
pRfRBhl2l+yrBLf6Ntmru5zn4b3NKLRlhvuoXG8eEVpOW0t2PyTvFeEpdWgYYcGt
wi23s6OdspAJOO0ScWhofVvhKmGzu3q3u9AFl/kkKJVO6XktPvdOUHNf8IiGTBcJ
X6sAb4zMVyJA4PeUtXjO+/DK6piTrHJf9fmqQL7b57zDZs4Tl78D4keX6zoIQGGC
KIoIXTaj+QsBdINx1L4kmDCTrAUkkYpXya3V6hV4a+RAJzusGXZUV7viEz3m8yd3
LPootxicoJABpdfJCL2dgy/xEnhJn9vdoUNIx2oMP8FkUEJ4QQHpTu7X9aQaktDx
CJPrI2kN82VCRVZwGza1xXo1IGVVstKv4yym645deP0vAi+MK3TKYHKR9BWjhTj1
50485ryFYXi37v0kiGaFZL70ZyriVQJxU0I8fNX75NnJgPVNNFIfCpWiEoj3zWYA
UhrxGzotnN5go5Eipb+ulJFbvxzHPl8+ITO20D5Pz1I8Tl2iiBBMOuRAghr8DHxT
5qT4G1khugFxBhnr9Bf+jAFptGTWAVVrpsHyljuApfSwQPRItTe28/qp/OjIRKw3
OdO7X1NI6pBDBAWJAieg3q4gQIb/VSW7fOsATITtPQRkQydciv6fFfVEn3UbeMUF
BSrWahJC6NK/1XvsJOTrVRt+0VwJOr3NM26VwZ/lJ8epln8RCJZavx1g+75fnYVi
3hj6z5joHZnUKSNw6vVylkn9pTpjtBsGmSMPvahJczYDSiV+2YoQPFA2VxmjkeaD
jSbe6g5DwkyWP1ZgvGEkHr5gO6/sIsWFXDPCcJo0I1Yp1mfajoyn8d76xxZ/NWwS
q9PP3WGUz/IsuB1cbIOgRZGe4rzGLZAJlR2ofWgWz4PG/pRcI9jrerw1MlL5xCeI
ZrQsPVsFVRSdpePoR9ebbossUJxRkjib2RLLRFHGJn23znTWpS7Eterbw903Pn76
HKWb2aHNxZGfKgNQgtvg9nSkXaI9LBb+5KZZB5kbj2CA3m2xY3L9W+gj9WnXD5A8
VtrYP0BZPHbregLqMMjLU/K18iZxj7CJT5x3qxHpv0Y1BpPYmKh+jkjiHKL7dLE4
mAFJ7OtGFOBbjg8t/GcKyHtVoTHfZK1YqNlLew3triQonNaCc8exrSH1hDhPDW/I
Fb5BRA4OYB/NsNUnxFw04l2tE91fFreRZ5B2OAXEfV5LXoqxuLp4nHDVIfIWumR2
PWhE5d/4ACrk2lvrRsnQfxDzAHrfZkJHEjNaxipN2uATP6g7xT37g/yueKWIZQP0
TEwA3q1cr/Zf7ztcfNYo59B+jF38s/c5YNjwGBFuKKqDaXOYNkZ92lzQ2aypdVTR
Ob95FPJDWrYZq9jchC6z7w9vzOKCwI2xUni66jznBB8rAjvjxCMIeq6PRg6/sdy0
sIDExD1pLkMKdQiPjGNjZ09pal5RWPoXqiAXqv/zKmtUfsEvvxnWm3YYbv8DQd7e
i1xONaZbk7WhMkciZfrKrLkPwdgbbQ01xB93Xh4065uryCU9XLjP3WX40nCNgEeB
r53qFUWdUccR6EnbHxqPwBZsLmZsqX/PiGd36Fhp9h8f3RQNEpGfMRofQzkjSzac
cWrGxvStzDar/gz9p6p6bhSnAJ8BHSFko5VlB9QNMmXQui/nMu1kkQB6y5wXxbKP
oPGrDqqS2Ky+mpfhrm50eAskUDhNEvMNrukxAIUbBWSggnx3tFY7XwhG2TP8VlEr
2DlCCZ0Q4y+Ybefw5T5M8SNIhOJrE9fnbgjILcjTn6kybD2cijnsjsFtze4OSnAV
wFgKFdpCMBZIImAvDKYKPxOdfz/HiB0y8DQYiiYY4nUgH1RgNl1ovURXaj8vV2Tt
NBYTDccx/PIEXioT5SDIfEgfI6xnTBiyRT2RzGXhQJyNBDD9qXM+UGlPy9Dqad/c
Gwacur+DDLdUoqTF15cEl5+6G2huXy6EKVyHEMEi2ADlyuOk8pz0bH25h4M2OhTF
E1B4zKqsc3B6Hib73bqoRTr0+G2W3YWKQlQWItRmZQnY2XjfHcO2G3zpdNxfG6SD
6EzmrqwN+bOGTvOf9JwZx5H6G69L3LzwYG05x2qSDhswbyrI7Cne0una4uWG4m0N
UW1HB8p1vNcxgWZGxgH0RDx2+qkBu8M+XwOj0gxQPXX0LczlmMOBvgSXzzMwFdR4
IsvxrkXn2BFi1pYuq+wHMFPfes5EVGF91mn/Vz8tje3h2gdVsP2++Xi7yDX1EGGW
9xq8Ce83EOS3ZWR6qWFoZL+aRmv1Ia6sDoNGr4isCmmugAe+xmZQESCPq1G/ENJ9
B+2BPTJOWazi8KUxbgyBiLkLKs4xjTrhZL5W1JnqlFv+S2QNI/s1V19UIEuoV9K/
UoAjUNPo4CcMby8/RRH5kJHYPPvpG8eMEXaAz3W0r2k82gwmsR16lLrmmcUUyOxH
jDkFEjjTRrf5C0/1AgfixObTFMDmW10teUonrCySU4NGl6gWxKSweBdHtfSGacX8
NAO/GBBI9LkQ13+XjzjiBVnmZX9v+o4SRjfIGBtPNi7eHdLgQSe3s6EMXDG3qMqU
2zIoWEWgvr6Kh4FZCJdZvbolzuljOS97PgdnZH8GZOejpFA36P6WrDxjCL0FLdoS
Xn4ejqDQ4XgkgExRoC4yNuBqJeZgaZpuEJbpIhq8e2J9a4DDcVbiJ4fw7B8hMxWg
YPhfD0BffTmryb5Nnvoe2/xB762RsSboFH7Nyq08XsX4pUmtgDoH+4Af8kaHGIqt
gFonxwoa2SLzL3QgwZtFPYMM4VuEs2HgK0l5oP5nbGI6VTb5sNghrPvcqcKpzTOX
qENoC7AP+BlgTfCqTP1fZCIMkITP+hcido7/77iT/xxE6cBr4JCjApTSo7Z0IjfP
gdgZVXAqZDVBVcRQKZ3+GM+Q1Uz72PblZQs7Kp11fKJzL8Egv5AiNQ9NRGuR258w
W2M8FhJAk8STsS45J25y0V0a2PXDr3zkIejkDPiRZdbUKCdSwJKqaXx16jb2RG+M
QhCu3Fu3BdgB+YSaG76biRtLGKOlhVLmdHiC2kD16L3IDB2F3yw6Pq3iRGhTwgxz
0kgy9d5TyYT8ccxbyeTAt/05mLWH12dGfN4+SrxhE+gjWug/J+oww/lzVLtw6r/H
HafajwQxTQc/EST11BogV1ioghskeTA3cwcTa3B6AQVPvVpMwsenwtmnmNXuGAyx
PNcT7yp2oEwTr0HS7BYKcrklGdeMvRoRfLr7zrjcaHrY6g4W+vcXQvU4KqSvJzng
jN2d8SB15U13HD6Yufan1kTaWp2FArgLIgAD2ZRJXVy27W3j8QTLV4J9wjHoe5rS
7CGhGb9GJ5e1ZWKoNhlvRa+1gN4FkzF5M2ZlJs0397SVZEy8jomgvUIx5gkdgcsN
T3wEtG34rMSUc2X8VTsaS4AlhHEasBdiPvma4lWLQpgGD3GENCRcGJ6melr1Bqqz
dH//fnwFy29G6yCU+CvmWYxdNdYH8D99HdgtnLOf2zOZZ7UrMonLiF75V+oURSP8
wovaXygKI8NMi/q9T8QBnb3/xoFT4p2nuYlqzBGCOhi7QUCfwLQLIKee2+7Qxm1E
d6ShloBV8rVCRfBY4JkPiU+kzrSkr6d9W5su1jNEvh9CrcZzXGUcfijnuOO5EtKr
J2V8YGz2Z6ZgyPDXTrH0JRZ0m3q3vrsUGLq1G7NTgNYiJZ+hR3z0XG+x/goLpBV7
fYhn6bUbmrbhi+HiQb3KwsVMCmDSOH9IJNdhQoOvsXH4/IUgqgox6HmOwM9fzFC8
14i2y3aMtAnCBhjOF4h22dQu/rSnnCA/dQjp1tX3bWvWOxSzUvTBsZBqIQZ6I6dq
UZ5Ybed2G/FmbPrjB1oYU4IfMvCxTtlkXAC4sI1FTtbG6F/+lm5BSTblHpN7H/mO
/hYdER6kzAzIQa6g1oHOlOGC2i0XQo0owvGmSKBjvF7cpXwX9NyI18xsyoqH0nCR
u/xRlCFghdwoRotz88PPG0nK/b7i6lxbb0N9nxZbTnN1v25XOII441SRN0nGsAbu
G9bJpv9Ng8SpJ7DSVLl1guJBe8zTe/0jk/xlzAzx1/KkRHLIUdnyCQdEjpMsXiif
Vlvgf9WeUIQRqFRwskpqb5rBs1vjrNddEXb/4cTeK2hyL6bDx46ju4SsCm9ZkJQJ
Fz0I12j0hGedxqCI9ImpEz1G/S7lY1akh7F26x6uT0IktStgej+l1B1WmIASWwd/
hM3S8QkhcgGA7I0R3rEsFBp/a3sHABf09cf0HGc3e4qWtndGxHCP1k5HdB7OjYoG
EVM+0nHpMWEN+zmIHixmvjC85onHdC0ZHst9RbdCs9KHtXgINYy4WDtcuSyc/U4S
w0AkwlTry6kIjIZaLva1NxTvjs45NS4Gxq48LXBdYgh6MvdMvpy5nQhng11cnfK9
PS5HVNTy7UYy+yHbv1Naodg3UwapieydwYt9IJaIBcnQMoIwyOHUaPEHuET8VrYr
21+WmvR4Lghf814D7y6rl0MS+OrXxUkq4le2XIKPPBR1X26EYPS1AD/RbUibcZNF
pBZh7N/EJ8km/7TYJRwbkRWb1LFETt8AyyfjTilpK+6Zj7sQeS83sSiFLEtfhlv7
LR3s0NZIlyiqzDoD/vXbZQG8GJasAD/JJ6uF93W8TenDo470UguUsutUY+Oa3aDF
fHoXtvhMuRY+JEOFIdiiAPZp5isLW1OibMXlfcDA+E+tAR3gl1nIblGjmDL7E7Gc
gwwPEeK2BZKxJuTnrvBJKPZ8nw4EEZMVtZXU11LDH2RaLdpLMnM+74PLPEyaK9HC
qX5EVFCePptvANCD56/fy+psRBlb59Z4qY3hdQcY/FohUSL3RYOaZSUvrjTEdEHw
9SPItGfjYOumtYFMFH2DFAJZ2c2ScOw3scEs/KGGZQvU1NFOTTLIXMwTNYRrDtpj
mjf5U2vEemE3xWQZTtP65+Cko7xi0gWosFombMXEShljqVx72//XnP3aXf6WLMqX
2ZJXmzlhA/O2gZMVVJ0kEyst0t8lbYI06mt+GxdMiVDTAtPFfQcVlQvFLPIFKOT6
6sv/aBF7hyJ6QV9b0d05jIrkzMqpXyDUD36SX9fUjAifsuucxbNpqXcN87oHop4P
+DaZ2cV+B28x0ugCcSEsi6kC8+XAFOzwQiXDjNwfUkdlw69s/qwADtcJjD/I72g8
G9rlxepthV2OLunF1278dCAMZ2cn98SegvQ9bgSNyfSdbHliVlkTxqWzR5TbgwPd
nlRMesW31o14nuSd1pikwl9LxuAS9b1Ri2XK/GhXeQRmTIBRObPqb7VCMQpEDPdr
ToMTRRe8xARNDJB5qMupPu+iKd8DMLRfVHs5VU6Qg5NHPerCRMgSb25zCzcD0rEm
iUdkGR7DLGUPmyVyBBA9JOBZ6niu+Lq7xrDIcLPoAO6v6unxUzJZUpnX2kyLsBsx
nUGe5jY34PL9VDrlo9fehaIHoU6jcYS25zXbNevEYybskLciZJ3+31o9xlEGCAuT
+q42dW82XgEi+//wi4S8nKTxsEjoEBk8sg28iFlP8heGF8ee1bWp08JFjN4KwqLC
MSAAs/9f2wamBNlyecbqBZsZ5bHcKPKkVSRivivbt+qnqpvGTe8q2BppYKj8NPKH
vyj5xH0uBJdJtAxfM9mzsbKlODM0UD7CJEHM0mkIuSLdopBiM35C+0XX2gDHdLU4
aK8cswpQsFhhtammIUPugLq/jenQ9qO3hmqMERYq3EHloQMTbt3SuHuMX4tix567
+OZUHM+CDF6zhLZLnp7Z1YninUFYEBwgv0HTo6wsMr7e5RFvdEU4rBOKKGznZh1e
2asMEAD2eks5jj87Ig/rl9cIkAmONzX8+MDc4EO3RupNy6tu+ZqTWx7ucJWgISr9
+rFmJC8cXTiqaCcTen/1IsPJlxv/iKasekcIpHt9J+0INg+Rfy97Op81o/25ToQj
NkfKYV9/oe3q70HWKg3gfr0nwuvqOjZaPvn0XQ73n3S1iMIiSn6VwfJnjsAPqr7u
moKDY7HBHuXi2J0AUQ3nA2alWHoIu+iTreSQ6zN4dz5KlSsFviZ0A6bufqLeA1sR
Y++aOpOwJY/dDk2Zcp9WAmg1OnO1NQ8qRXINo6SbCUesyE5lxmNoafFdYDRI8TPv
s5JLBkFZNPuQnnGRjW2GzAleSlxIn/N3MvoKcYiFMurltH2mhvInUL5PcPQpG3BM
7EFEI8GJxuPspR+/M648szFvx55d5dHfIBNUx5uIDhMAw2HoooF9CKAz9BHA/13f
YRw6a2FmqXZbCjwhxGU4oSHLD3Kh4j95MzLsVUhjfoeC7d2Sdi3oH4DdsyjXgK8X
0svkYJCzzjGWuNVLtdpnhlLPlYW3HjP+7KVgzfkR/xkg9NOp0REg6xIsAJfa8M16
KYRpubUBpEbsYDVUt5hyi6OBmg0qsEuLEjh+nG7UukZuTnClMUoPzqYc26wRHLb/
VURH9gHlzEbSn7zfscTCYBCz+/Kdg8VxapX3VLHb2Nt1lAOktObxiW8T14PV9rw8
KILNEJpa7640DF+lZVkwbVrRInF7GAuwSKjzZC8ov7/L82KgWKlj8MDnN6PxcpRF
8E1n6DQmskxYHgbxNQ8laPfsYjAEGmRIMW/kmrto+bUbxkpSDscW4iD6xSpLwWTC
T3GdCeXGqZVF1BFHeecRElorj2POFxHhZ5fjhPJ/cykEEydB+3M6TtUA5Fkjlnyk
4ZZEzMqAV5rcLJE1PuST1jSBLO14OWJKNqU+7+nqdpkZmGPXyjVM5ItaB5eVzN0T
nslPATjb8mRiNK1HN/e8YQUBCCRt6S10/rIlguAv1ulk1x/FQluBXAY3DIpIERLz
tnWweqnXwetzbo163tdjcGY/ryfSXyb4z9vI4bhcttqBwtkgKPQ6RfwweLcmrYot
8sPzGK0XdXxx5wAu3QDMwEYKZ8Sy5BNKNRsg8YdCaXse51ekHYC4nWT/iL+3R7G/
/v0sHAjbmPxw/KpxjvzicCDoHxOFtt2Co+f2dQuwy2VPxPt/X1IRxeqsej8P+HSA
ZQrtwt+i5nPH5NYkJDJOmuv273m8Dj2JJeYHKwycOWxddZ6omnA85aUwM53/10ws
vS2gKR+ySCVDDLmndHvYc0TPTo0X1lP7k7KoPmeASwHfJi6PhCZ1BY0kJNb9ynkf
Ryzpw+ei1sR/0R5FVBgYJSs12KanX3gvp3LKbzamEYPCF3rZTbXR59rpZMZCW7mY
BcFlH8SrI4WO2d0jx88yPdlNVAVSEbtuunA3mDO2w+KrKmqQor78NvBdtVk5EAcv
HopCmRe/GSBG4YMLcrGw98tb5hG7lmqfBrd6TYTc9o3EfAbuEbz8S23KXERpfmHN
m0coQYw9DXAjt116wGpPFxeepKTLprLX5NIKxL16MyMawzOSjwyQGmhVU8aXVi4K
+wmcSVdVnmnedfRmpmmOy2s4qCdMLyecBxVz6AW9T815I7c6qYDN43D2O25w4Q0f
oUIq1Rrz63y99PEK1O9KrPkYGwDomH5kVcpm8rAsx5zH9wSblQO+NalkHJdAXy7L
j5C71OjQKnH0wI2ysTpxG9NVXs/jkFYBEk0NyTdanWDJL59DkHu958kOViEVaBo1
VW7XzduB3VF8ccPbMDJ0q71v18f/J/wFa0l1Y2+ohMMCPGnIvDJ5mm0cCOgKLem3
KYfcV8dhACPhlQd/krdm4PtrhwhIHv7iS8XBijnJDFV4LCeTK0oXuR/q1qqkuD+W
oxQWo6LInJtv3Lx+Hb4V2MNBGJ+6jiz5rWSkAFyaHwGcK12WhN77QDP8NP0u9qYo
QVgdcapsC56lI0L2kgyitg31Npf1deNZ/GF4HzHM0IgwriiQyJOsMCC2kKYGhSkV
CaYXVMfvrWBDxbD6UpJ4lmpKOZd2dWmFmnCVm0viAoFrPPMFJQC2tZRTeJLdW/Wt
Cly0WQxg0IQwY95eiXpegjGnhyMw4ZPitw4XDW7eRQsL0I66TzG8VCMY2dl4YYmw
CIjbs8Z7FHt2vO/dm2JsYhn6Q/Y/eF4gDWSlFdfa4lbhPj5OVD5ilzC30QzZX4FU
+T2Ouf/PQgVDV3PbRQhvRCVg0doeSV0Q6GtxRJZcUw4xME1SGhLjSU9obsS9kii1
3SE+Wv7D72g6ukQj4pjC+iu9SFPIifJDvo+kjepkZaVq1JgDh1xQhDmp01s6NVEB
jqytIPNbeRZX9RJVO7J+r2EZMHVNAECIHiGuDQO451iFHeGY93NG+t85Y0OzIQ+8
uTI7ge+XP7rz0t4ndFc2n+kBYu7JzQQJZBJR9+nYbekHWhdQyPfclZaV1BBqHzvh
Ghdg5f/IpXfeSogeWOyensJaL/aA6+6VbOzXsr0py5V1z+dQmNaP4eGAusur8wfA
vdOpG3NDBZap4zhn3zz3tNRume4cudUCZYXEJbTTwivuID7VFb3tY0xnJ+lTGASG
tLWvUpCN8544iLZVycFSPf7BO36p/SZEqqX2AqGbVNgaHuoa/9DO9eV0lXjO5yRn
6ra1L67YORdbqlw6JIqaObgiasYLBeYtROkDUZSw5kalcgH008XZCeNqYy7iMX4y
irsTEuenbsMLnp2x2/QFEITuW4zKKrP+5So5XYA5HnI0NSWab0UHnJY9Zxi26EkP
mZGOpdKFFG3/szXKvFHWF2pZqEEKKjTZQIpYjBKNd1tARdjmW17wU2+q8OeoWtW1
PjQY2Tde82+1YlhT9LpbHUyCtPgjOfIEiaXKdI9NwvaRolAOQSzX+5mH+vBhsDJ+
4rRIv+fk5nz7ikDBJvh/GqqxP4s8FlDrPoZsj0vzM6cfS+6NhtoEbwhjuV/1AF23
Os00EGopWCPo4lDNKs2CdLQEsnEDvzBF8TbvWkhTU8GIrEhRh75nbj+BVa6u+sTK
3xMSqDxK59QrgnP0zWhRZYaKPn9xqan1HuVYnVWccGQsz61KZOU+eu8O2/nkb1Pb
SA4FWSvKrUcspj/aYjMf1m0gFiYwZcBTBzqVxT94aB6QGyk0PNCJiY8UMVLkpQPW
1uFonimfp0TwrtUxcXoUSJqgJ59+O1H5jfuS/luqUsv/o27x5wQwMCJqWMx09lIN
MdqfIWx5bAEEzTems1mVHOGP5oLijc3qCVavyncldF5DqNbA7sy1OsGMK847dQ1E
X8n7GaRWQPY6zMgB23IrDpPQI7sKptwVmlEoWlDh3PSF3b4hoDP1YC4JnWGCI9Lh
9VZmEuq58hMoJMB+LA1Kx+fi6kLjOysxn/QxiwutfI8i7z7UCBsBxYJj56JAHmPX
q2dxlm869xSnlQ0hucXbI373hcJqQZwnC3FBWqd82/BXYDGB0x2+UCL4G6HO80v7
LUTHf0oLR9XakoIJPHxNah8TUCzi8SrDdq6qtwzznD0CJuABUQFDf+lM3ZviA7JD
UEcWmH+sVK31ICvk81fFfqE74j2BdKbOalndMFMS8PGXPGPuhh4krIxuKV/yc5ZN
bMGGH6/q5Tjite378a7zR9UQhXBzxEFPAUB+V9yMtz7526FLYkrNmYGqV5mGXHTo
9wqzTL2lmhAMKT2pScJ6W3wW3MjNucrnfHWozjy+u/GGS1b8ixiu0WEnNsVkWao1
6KUIE3qOoImKDyqUsJNTlZBLvyM3BmafMOg2zevLfllDR6k/oLSWvBi60M+jTIFh
Kx/06ZbCC8hiv2/h+qQ8jCEGNTFEsyjf1K4bjwykZjjICNtiQEOyD0CeSVdh6EV4
yjhtdzYj2Bx2myt5xn5Bk5JfFN8XcxpUwtWODy83Cvfa/Ij3Vpgjyw2NGavnhZcN
XUlkwKAlOxBC/eckZ4xKsoPAPi0iw9F3+vsUI5Pga52hht1MgF48FO/TTAOqU5a5
Tf98AnSJRy5giSri/zwHT5StMdkmLVSZ93hAXZt31vwEPuzUH3XXIjm5HSrybbsG
FnizvGP/JophlCCwjtGFgCY+vrVsWz/F9nbzDnY3loHm5xL2I/744JLq9mE7fUCz
yzm0iqzCMovYO9+Ckn6ztgCCoRpULhXR7/wTolAcOd0tE338ctFpoCRfiATmmdas
SjdAX7LoW3wluwmiczis24EGwMJ6/1QCn7SQTULpfKTqEJj7KgkznxNFKPy09peI
kGsYByNXJEPhDEXOIrifL9DHd2mRzje/gmEdI5NQBQiQ8Fv0ayzdGy67pHyjfYRA
1v/74krWoxWyM0bLTJ86kPx9z+zzOB2ZNjm+rtSVvavChKI6uCTMvnWzFu1J6k8h
w/Qm9ckS1RVy7N32Rrzb/Zlt10YUGjbJDAqZmkw7djy8uZGpkgqurP171gguj08K
dcRvYsuTGG/rJIkqYjhmgedYgxElpQuIToGfBDe7VTZCdS5TXhEjFmPXlGkFeb0D
NeTFUCWADzNqrQQ1WuGisfHjp0VsrVX7Ip4MVjsnWynrX1saCUdCW2JNuK15IQO9
MGviCN8Gzfx6rUbSQESC1NO5jMN4VbWpMjWdoXmRhn+9gBzrKvEN40zRRdypjNMh
JR+NN/8hrY7a3sukVJC0Zuha2a2D2gWKMPdJ9NIkQbY2357LwqlXt4DIo0uTQigH
W1Bj9gi/8HpV4LHlQ/b9YGj/Ppbw9zE7S7wgw0uy9XwsQUqO/M1y9ghwdP8/F6jL
T9rdOUmBcFA0NDjOOOjuSxJkgmFzFcNwtF8ohqBB4r7QTTR2dh30zqQgYnZJrPIU
oM/M8ekgSg5g2BBH5bZWQcjOALOV+XT18FHP6m9V14uNt6xm4PfMK8NlN3UPbDwR
NJqCcNeqWfzZHL3BPDRkfbvTvHb+oM50TNeV5M8y+Ze1dqD2fMjj1SuqluPlAgNr
OCL8wjb2dY7y4v1/JvHDo/0lAB7+fCEIM7fOwvgboinGQqIkDmRatUNrdjiPlpce
t11GEigEyRoSP+Wzq/f3lvHSYVmE5MBQOX4+zJRiWd8h32HkLzg/rQtfwBglwBdd
OijiNOWaQFoSQIusJUed2x0P4ZRNGshuGEqmxpm9kIcB1QzGhR4xFj44/NFUN1HH
53SNdxG/GTSjq8fyRtI6seC923ILmjnShAkkFQs8tgEh/EIfRKD1WBdMObznt7PS
AXJYVqj9JwXjKRkFKo0Y0O1kTWAUREBGC+MMqIeKMt19O0uZOCUZzSTKfD8/tlSz
aDzDsWLlr8L7e97EmBWnEQ/VyVxZJvSfg+mYolNlAhOSG65fo0UY/g8OpfojXMNE
FF2t+RvHxMGKOzORIjQTv5vj+TNc/tFtfoWiQnUJWiZsgdDYvv6OGEuJKHR0F9Tj
5SAwvVz3B61aTwGXHRykS2+zEPM/NVB297j8rQayqwHTsijB/wUFq0MftiYrLgdH
bW2ML1qq9O67m8IhyuynVkiM27G/C+OTSOFIVBy7o1t9VTUqB+FR5BuG6V/wwx7g
0GVyh+ubgT2PmEtglvmLOSV91rL/+H7cCgq1t7yfgowQ1uJ7AE8Qq/X2jMnPMa2+
huvHciN29GbsduD/9pMcSZzvp50Y3ZPOj+ih1UBQ/ravIt8+xZSH/VdMQvyiovZx
MURjk++S/5jkhYIZcvNW0TduOOrKKpeGVAO8Ej4k4N7rsLOKIz0Cg22Su7tfQRQD
TSslR92PY9nxRBJh1CCFBod96chNpNb0vgzhS+cOmPcPFqiFHlE+0VwGUd0K8wex
bp2Pcs5UsdlR/At+QcV4A8E42A5nB9p4/wLQd09Vp0IV+Zi9RQdxjYS1z03wPMLi
+5C8PF5WYcKP0UP3xQh0NjxeamEcuGxO70AzxLTomHsphiMM5d0AByqdEcobhs6V
UI2UBHUaLaYR0ICxCTt6q7Rlwbwlw4moa8dFaVs5obkDssFknqofi2MSPReWIRSx
5MoChGUKnTGfZX1hlSVfoWR3deXUwwzADyUnqzm04LAtrDtUyV3Jtyd6B7zAEyLH
udvB0QL0O5gLjws5hfPwRdnbXy0XeU6I02lB8g3Dp5RrGPPeW4baututzpKSzzwo
pJhyIFKS1r/T5/n61MIe6m5lFUg+wJJmTB5tw1pZmjBtRdpvPQiIjXLn51vrO1tX
rudnZyx8xjcK/PZ6NxSbSqqYKIpbOXDfXJhA2KFyx+j9y2drDNQ6ZywaEpXtuF4Z
aXpdOSW78P70YcuThl/7puyixmvzdDhIn9P1tAJWGorvMOf7r/hh439+AG0kTek/
jFnoMLw/cMxu68woaftntHJfaNhDPhccFY4UEfx0cUEfW4CeLT2VLbk/ARIgOpLw
UNvXhTE+t/AfRn+xDhsivC+9wmZva7Cdp0ukXMTLPq9dO/rWvEh72wemkiJRHzIl
7gJ/Ul6HNeHTSj9NB6Jj/U7Oj9d89i7zBDyIRLbcLdALrsbSK7Jfvufh/eBAB+aZ
v62CjJqEM3ypSE/bKXm5DxfdYxMxRpFBaIJLnPOQcpIOgwGuTHnEKa1KozwV3JtH
U/8hxRWSkDDg4LhlA65w8bEE6Crh8K5BHr7czpnuQ+XCOnCGFyQNXQd7ycfrt7cK
2FKxIyKs1GhcKcJTmzdPj7YyaaideFBGC+ahrsJ35WtAvRO9CMSkzGhVXccgOZPk
SlqOt6c3zkoqhcJXkfEiGikS4AzJ8Y2Pq+cA5JnOHD5Kwb+D3tyLhq8thxWXtnq4
zuJt/4sS0hZPbSDtIcCoj1MWPKQ5Txbxs+2ePSTxYdIJeMpFf8Sosgj9atk0Hdjb
QOKGmdPeP8wFwFGd9BMn1599v7zY9b5LvAO5OzxIUK3hjeEuE90ym7vvj1YAbBCL
3HpO1Nbvhok0ZEeOajfvu10iit+8lz7KYBhxIiPUnLrgH3/e5+lbaXotzANMYOhC
RZErtAlaUDOswO/xckt2lS9NAkgQgV4/dN1XRSmBGJ9dX6IFTSwnofo9oIR9h5YQ
4X+LLc+bC6gyUjN2zfGtldRvE4ZKet8B2xpJaRfEcNZZqnCA5bv64zT1HBFWOH60
OlSdMNve9rLzbo3m0mSKtE4paG8R1WObFXNNtrbOQveabrWiAYSJne2szVuuVTXz
1Fyc0G5khPEWgweXvx/LDKnxz6Nf5Utaq4O8P5Hhbr0vbZc7yH7RXJ351PXA4YgE
88iAyq1QRDY1PgVg55C8SLkLAr0LiBxNUVxUn46I3vLjuhgouLOup/kaA5JMBZr3
o03RNxs6w7qrmIOqWb+CNyxx341/FX0tUWkJO3E/UldU3C1Mx4k9c35e8UKKqPFZ
7Fly6mFQF1chf18P3aNjKCCU+k+wc5zKeRdxrP0Rp8wAOxhya7EghCyqJAAJnGmT
eZxuqDW/g7GrHKEyx1NYpirotFM8QOXViSKfswX5PWAfDcEr13Uu7aq1wBqHNOGc
VPTbyRg2ahAimgd5RmSc5eCJT5frGPFmIROgL10mg8YrhBZ5hK3cn976pqTsX4/+
kqPNKbKNFnsF9LnZBnWK3vP6RzPDdbqpOVRW1PgBSrRBQ15oEzbJniSMBEEEeZyD
B7BCtu7LmiRX3VL7ycd7/SE6ZbBcvJujz5sSSDxMDdoyldSp24Jwwb1mmmkpIkZS
5LdPSGlRypyuWx092zaPLopz0kNe9NBIp1HXifddsLj10JvlcXi9vOttrynnNp2S
0GozN+ipQgMcFPId/p8VeuyiDt+OLBzK2GxcxhXEezdlZFmkPeci3fakQaenqrK1
s5FYjJujMt4CkIHvoT6uaOfeUy2NaLtNg1FvJfcOXRDa0Bn0O/YcDWadeUCW2TS9
pxJPMf11dAO8kx0/BvoVGqyDxkzrPdcjvSZpIzGeobjC/r9U/a9c14mds1ZgnRys
UQvNr5zFc0+BO2y4LXEWY/J4MYeOIfvcFWnqUBXWmyQiORrIJxXNxDiXHgaV0Ynj
8TzsBWWoR6siqILj8naadXiONrA8xXaAV15chIw53xetTrArRllEG4pr0BO0gbTW
35byRZv6BHuU3XcVAD39cZK0ROYuvPBPZzs+vfMUqvNPfAOMO3RNTzo4fXPA/+X3
rntv83iveuvMfD1xv6P34YTHFvsxElmGce7kQ5UlWJgcoDRgkg90fWz4a8S44i/s
05+iTayn4S8g03TYNFz1B+W8s2jLKedO2FagXpp34NmRTR3Jqi6mBkTMpsOpKEqE
r+28koI4oouTSVlHB9kUxZsGxZRsCWMmqycJfTlaTT1xTuacOQ3SDVdiorypJTQm
XLdH3PeuBb+rEy9MYQ9743BkkGwne98j+yXHE7gJoZPJIRbqO75/0SZtY8pva9iu
kS+6dkfCMKT1neYep0brboYTiVMaT6VYPtFDd8mSUecZJOZAD9Ha7SgA3ZME+hLh
AtFduPY1YpRU6sCCRbTtu6bO6Tk5HoL73AJ0NcI8c1k3Pwim+XowbAUKWaGuiGX8
vd5K6kSnlL2ebQJaxuVq2uU+q1ZOuRgpZv5ACt+1J7Kv5DKEOhHRJte93093Zq+B
n2wATMiK/v+yv6ts6Qq0c0IloXGA3c5IiX+98tOrnbM7wPDkrrjWPC94sPY34dYV
bSpSOiSS+f5czhuBpr3rUUKVbt2dTbHcVxEiTdOZaBjxH63fcnCGUjL9cLYbkjB1
UFMmlqnY7SNe8N6CD76qKoKQnM4gkXQshpfDDP+9evcOWcIKdyh8eNt4nKvLEzKk
14Yzq69x83wXJdav61la7idkhDZf1yedmseo0gTbeyGk4OoyYb03l3XshKaBFV2p
/h283tnOElD5YIUkRwF/4ln/66ZCDKUrEL1cfhCqt2qdyBv1mob80Z5CNWZSMS9c
LiRa4Wiw5ohUjpkZ3Aki5KE2nNj9y5KNZ+ixF6eGOYHtJDas1mGfrHiW0SlW37a3
+vMH4+bR2E1hPzufO8uVJHzdBeiQhjq9dmvXX/gSIPG1Y/N3imdQnDdsjV/BucM+
IgVEFlQgHUiF7FOSy7frqezNzGxTDVJ38a/TsVUmMJldMIuToa0r5Gh4jVdo+Dv6
9WPT1vMZJvYQMsckVmxcizGmfC3eF5SveVFtQ5yp+0x4yULU5bJCZdK3chYNE5FH
YiBkKVhACsXmAnTziL1KxENntWjxz6XinRlSjFvWLRfqZ5gRvDuJVquiCXPwfGeO
B4N0JO5ElPy+YWC/crcZVu1JV6dEbIDnrHYi6mfxR01K4RNSGKU/xjRtNYMZYrMN
9qXSxOPawLSwoHRhBmwlJUtmtxySD+wIjjYp9e82wDBkcnWcjD6ZuXxVKgKxJbJr
s+BoGJUq5mIDgz5Kvq+3PTxqsezaMQpaxAdZNNWthqp2FK4TnLpWUIWen+6tC9Ht
yHwHrdyDIM/AxaNdggtI30qQM7exzTvJ8FkyMOBeDiYDyXnk/akbFDNXm6EljOwy
ACZccw+INURJyok0GJNVFaPV/YoEZSQLbymfyGBdtTh+xvZDPO1de9gluo2ml5S1
AcAFn8IbieCjM5emRIt6Lb+9KYOm7u2tmQckA7qaYnjhH/HSEL0fnqiw/sUR6cEv
csiApZT+UUCsNrdnVTenAPY91siVSpc7yby/K98u8c61jI/o5Zl2ijI2DVANePkk
jAh8K7yYN76wP3Iux2bsLxFv9ZeR7HZzJ14fdegd+pZZ0wcSFVbdR5e1YHglw2Ow
VchrVDZQgY1EekSRexwtxn0xGCoYN/czJAoUqSPCf+PB8sRIIhZmBfFemAR5gEwe
TC+V5dycr8259ih/J/k9hRE7E6bEAvE36CcGU7mYGQShvycuI70C21zqeLH/UDeF
37z6KufyCbWfhJRPHqp94qLaatj5SxIar+stTw4Br5utSBSJufdrrphCvmiO5CJm
QtsOYsoDJN/KRdVIl2nkvI5lYor4DFgg0j2BKQgMNlacFoI0QrKEvEZevJxl9+7N
NNcb23vMIdWCcneYN8n2EGDYDlPh7sAUdZltyhOU2egy111dcKiCnPkpSevPk5Yn
TlAO7/+Mxjiy0AtHUjninTx55gEHK1ylVzw2D7EoZzWe0htPWHguOPPFakjn4uR8
HMOT5vkBQPzHjkjquMr756z5b0HkwPrLNUHBpVAonsVg747pFmR5P5IxxGhlpoSF
UDcxhjkPBEfTjFh9EObuUvJY4fPHs3Wz9ZLxp6YrM0OAmo/wFA4DPKQuVJvQVrqS
YgTO7aUPDTlBI8AT8MP7CYen5JXRes9dKoVN/ARahPJ/MuX8k3y62c5pXqdsM0DL
OqfTzdJLD8RFog1gmQhqhGMRlEdR89c27IiPq8qdj6E7cWypF1Uud2ok+2lC5ytV
vju2LkoD+wvOGi2EJZ9W6wx2maFjAU9VdKf5WCTybbE2ayVOvPabf2aPVbREKZ/n
+oxD/hTZ2pEZSvpMOq34qfwnVuGkne3Ql6oIvSgG7GXoexUAnS4daMnsXtNaaYzx
FvS8uHvTIR6xmsSYTWsHDWTBE3Z0Fe0EUJXXFPcYMMQWkdyPsXb01BzMdo9vsbXO
W9X+G4hKxgYYuTtKJ+4M4hQ9DpJevIKAsQCSHjDGDCXdOSNfgK3eY80ooKkbXshg
it7lY3DzBx/5zeuHU9/lGsytKpxE69vwWiYdjxsfyidwD1owQEJQeE5Rb6zDDVma
3wDnzBRBYdUEpY0lvNkhTcHgbiaWBnQ4ZhTDmso1GyzdAn3R5hp+4l4Bqn90qQ+W
rS1eeOqCv1Alp08jju7yTvsSX6cr54EDo/Grx8hBArMR/O63kAvKPbJ9yhcDHWu7
nd4qUEau9fPZaGnloRasYKZDr481mKmuq+0PihzNLoR6Cvkc+Dql17p5fLsTsDxM
Rg9tCT9913Mb896/VT8oB4IVJJPNYuRqAjm3BK5Yb7+9au1d2/Zr5qmNZaBuIW2B
QyPcjZ26XgDfh6mKkLmizUF7WjuhcwpPW6IjUgEb89ACBG177Nh6HvgUXqhB22pE
hnq9u62yg95OGhnI1DG9AbqNxaQqti2C+d9ru9nqJRg/IOTzxhW0szc8GOPHh7Sz
bbOXGfLVbFsCISXZ+Gm9r7Lp/Czaq10KgLBhcz8T2ZiCoqvhvA9Ze6V8eA49GcSB
q8Ppf81KDIBXGgIBRvXxz3VUHbVcysmXDxTmnEpiMIMao6jnq5E6exjSdBbS+Gn1
yfTE8O+JtFBuGKJY9zktDkyIIrGYxWf0ZIgYonYyKUOqjiu6lFJlGNcqpyXPkJmi
g9rp7Xr0SNzCVem8fVNqJoMhI7m9A7Ozzo0q2a/y9H+QLC1HHT+ApSCgC12+uOB9
XpnlLoWdgrdcQAD7zYBZnt65dvFMIwUzzTt35C8GPlQn5Z2SIXUIsDx4L1sbDMQu
dLE9FP7NUobBwKYucwhq+E8Keo3mOYyomVoYbiTpYWn6L9rmr8Xk1jOI2i0wI7G8
wrTG7htXg2IVYrwhUYMa6nYCKMhEZhx9Dz2XpJG8xvrP+szy6eMKUMakoLnUG4/r
bcRJ1vvARJvslWIVtqg36tOHCuqlhDK17shJ0+CnPvyKSi4C8LENh5ZTrb0ozGL4
0UaK9VflxxclX4MnnGt5v5FQdo1u/DWAvgoUMb95GE5jDfqRB8QlbYzRKpVXNpyb
sNemQMEQ6mZQB/tOvHnOyWWx+nq0iIC+zXG+KMlGorDIP14it+kcQ5LXOF96tAZC
8Zouv3hyB7jSSji+tlMNxL8kwLD9KQYLhaqArpEvmw2Do6a6npRLp9uArqU9uHFA
XjdMQ2wEe8/hT6GN7awS9teSgW0n3a/DPv3k1YhsPiGGo/txJhaZCvgaonvCsoju
5vxApdwJmTcMGBBgZHkzENISFI/a7wxwIM7WMsrQMae74CqSengPoDBuB0VaDA6e
9iJ+uuei8E7hoYZoEiE24VbjWAbnpiP3BDyhwk/TYxIkyLJDCZQdu6abfjhj4pw8
hTUlqzEkb8yTIvrKlSK47MIZdgPsWpBEpMXRg6OhfJF+rv5cilzvqsfEiynSEFLH
flQkps1hnZnMPUu5YT+TEnGVJEcsPmTMLgFi8dMMynHeaQtyTIf0SsFZfDZJJ27o
ewGrfdYdXIhmw2eiLax5j1osxtX+SdsesRXFY8p3xoViByhA3zF6w6EJiAuXGYkc
D5A2yKA3roR8rcu8OtnXpJcASp0VlNRFhainSEZZPGTGFF2ILNxtNhLvn04JkCLw
llDxMpwIQEWz8NE3CJVhUTVDr+26eDhnlvYA0R9x2jRgTOK7hsJlKAgbOs9u18tB
2G+/zayQ+G84xqYrrdk2MpZXR364ONWcklkKSvCDrj+z+tuXbduaNNGBULLrzItz
OT2QRPKch754iAc/JJS39d8VXC/iW2tHRqLlXcjUCY4SDyxBlx6VQsCskqKY+mwu
XRDUpCavEUb6A2c21pMQFkfWXwxDrth95w8ic9zd1H5yFSPkwSXClu1X1X2GB7KO
0sF9GGdO3z8oq+tj8Z/1JyeTso3m/Eyg+NRZl4AlOGFwCwbe/vxqpAleOsxkVjlP
LF4b/3HCSTyioG5hdKTZRihwZwF+5jQUNU0OExJ2aWpdJ3Uv7cTKgxBtBTKKBQDv
3OgyvxD/rUzu+gKwfrRuPl5mNnMZry71t6SldvBKnMcm/vmsp20oGP+3Okokg+ih
S1uN5lhm60FHSWBkuEaSJqChBJjtN2cRKGGlbq2J/kJvTOg+2oZ62vSfa8At8swY
TJJoYoiiInX1LN1oSqxRvLumqFTneOKSA6BUfxEheK+AWEaTEQ6Mz+J5IMXyd2KQ
yGVyG8o11yHUUn4iaNDMOuigsjqlN+pbY6a+/mpfKJDW1Vg43gXM5ZipC9wBu72r
IshHNx7U1Hz7687+mnlv2HyrvcEQk+nG/lTRIyn2K+hCcFu62nUeeuK0awHdr3Te
p0ogLB/Scz66PGHbqV50y5DdahziEd+ojnF4LYkVAiAJTMGRqnqzy+Fw5BMpW5Tc
PY7zfYL6el+PrC6JySMIDAJUfCAnKqRqqlNn6tVNLwE3usDvASHkx7WeuH6ZKr1R
LIgqzrhKyKeteKg8oJFlgcYmPcl3xCgg2aERtaZOZVJSQIjbRP/7VUPtlo/hyApT
AqII7ui28eKZKr9DHYLnYHKiNK/vZcGF8jbE/BESHHRH+RaIiDrXcoZKLAItKNNv
VuOHmWmm9s6q7szeKrbNkGkTb20D1aVusD484gKCPl1lNVvV5/TtvwxOiBI8BZe1
MKMCEQ9VhT016RDr0PE3BOhe3tAZ6SuEKGClkQVdoUAPyCsPaiLSjEFDExJPH4zc
G4Akews3+mXL7spcFxdQ4yBYnzmYaO3adH+gHaFCKd0LkRD93f1Kv0UMGN1Oka3w
1vC+rGXQlcnyQ+Esv0tfMzsQTOGAoc3lMhtqFRF08bEgLMjNlzHNFNhe62ZfrPwO
KHPFt7/SUDnfZNcOppD+ECtNdhhLKOqMFq/IIkJpSYJ2cYFz02Tu6XDEPLdXIBqb
7Tg+RVE4b84o+PinCBfGoPmrGSPUUJXJ78TR7ivEQLp6CdDeDSBnSmjouom6A9Ly
NqgvIJE39SEmZoVGYqSOHXAu0WCsl1cZw6xTCr+ix9otvDBi2wL3TazTR0o/+ZsJ
kBfSO50D8Y/LM8mfn1eXQktuGd3ZNrITLAljY3IWU617UpM4bDGC24+VFH1ylYWJ
GtDGopEOXn/whioH8hvAArEMyloJgtO/uxCgPPwOTB0X/zx4kz3xOw1E6JraUoCP
kjBK9//LKUKfFSY6kovQdCR+Nq+4FLSnSTuhbJTYnurOXH3sSxXEcJZ+pLfxXD2O
ycolcT2X9RkhD5oWaB2YatFUdLilICVzqgiahiMRuFif42jHkwBrw93OfCWHvW6H
Tq/mXBFXTdFSRRl455JgGjDyriQ3Zdqi61XW5Fk2t9WlRLOwcd4OLeVgzuzcM9Gh
zP1fFgzk4yiFCTkJ+b2wIhT2og7LLJ4zuk6O/EiCI/GJwRK23MSQicujQgSbDKRr
kY/e1YbeB97wEAetpCAYFyQrk6B4aFdkr1J6QtSBZBewixj9eQ7k63vXyIAi8Z2Z
Z6qZLVZtANQMY34d81NYLqJl9qNcCBG/LWmYn48YOHGkBuV/Z1QHsH43yYjdVBhR
tl3YICw/LgeEnq63uVoM/PzOSv23Hjz6BPgbchDDIwMl87YdgGpakyxVN26OmO0r
a5teM73p0qKvsK48OmGpwMNY557xF5WJsl/EupyfsBu4KfaK79OHsktlL6DWgvki
nW1rxFeQBSIkPipOEOPFB0F3IH4ePMtGqaljLZ/P5UHTMCd00JTjN4WXIZasTcqk
1U+8T2dMeCZ2TSrgksHfAwlwC1mwMxK8X+X9Tscg6U/HRtBC6UiyNA443B/mFM9T
8GAdgjhx8SomiuCRwRq9aWi6abR5sevP+VXGtsu8ZcqxMHmsf2whoIQLvlvaTZWS
dIa4TIAinVk4OtdbscyaObg71HW2h9hOEbiNwjmuWRT+iPLR//2MzBIzbNNpf07H
wsWgCl3ytJEy6J9cIqBPN/GgtNDlkpfWGoz2AQ4TSVv9Si4d7OPd+gv5bBuM54lE
2jo25OMRrcfvMuJLiURqiTyIvZJr7f4am6eY3W3NKArpefc7OPxpxxKygyV1u0L9
2OlWQ3cIfUWBos8AVVilKXAZzPicT2vvcOCo3fmJpRoU9tMUA6UHlePavaaQLBQo
RwMrubfFrzWmRa7dhbIyDBUt2vjyw4dupMsokajTwEn2qQvQfD3lxOfCvEK6VCap
PxzzYQEUz9+ScFCBMxHqkQ8zzo+OeLaF/aGTAGG9NMqmb3V6nMnNzNsQkP16lwNC
KGRjuH38Gc/+X06v/LZleS1LYQgCOHvzKv8kmJQR3N/tUoIr866P/GQTQs/73/uF
P3YUiOeV9pJEUYrV5TdfF6Da/9kl46KzAjXpc5pbavqYrUjwJDXodyU7QyPCxv2f
x79shgVlJ2DMqQjTxe5RpfJwUMkXKkW48kRlNsDq/XLY6bTefZsqf4fwJffTEPJg
0vLT7OtUAsvjhaff3VoGaA2oJmeCwPk0Hu6gGhecuJOt+nnR7TANwm03k6EExhT5
TXvtqTOKADQ4RzRJUPUd4YzJzR2yCyXDLImp0sELRFRRsyluNV1fhuCNyQYFzdzf
qJMxzVhsiS1UHn5aW117bOUVFDTSiOr/LbA8d9Kccf+18jUyY5Zp9agnKqpaSGQo
lOLbFn212473/ZVq3A5EhM7268umgVjcwgia2Y401obU4ijpLYPa9PECnwJYbN4S
yNYerFPJFoqwU2OWntxijMpolX2O/ZIoVF0qowBbSqZhsN/0STuvHHksGBHeRsgv
NAqolVlqFJJLJ2vCgYkequg9/BeMV+glzSyddtv6MwPxbjjjqsbRl+VotmqePEG+
8kT5vUEp2L3WfIrmoVrkvdjKwqAJ1VbaxC1Na4SOixnwt8/fsRw5WFby+AB4gF/H
PAap6pcwBd+dNzTDc3NE7kirGWab0ZE0jR0EIkZbJRDV8cU3Eyut+Cy3tqszCtxM
7NeiW7sRb6mIP4sNtXgNZVDtnTo5v0TtvxmA6HGXf5M8gWp4vyrpCUUB+AL3fRs5
9FZrCbIBGUzNGkMTbMSnSSM0CpNVRwExCbgOBrMX1iVxjz1dRyLbK8fsqWVDWkKM
YqzmDF2tv4iEz8lG/HT/45TKPBhRHY+RqLvP+g4gbKaxCNcjtBLDK8IXvk0E20hs
Wl7vbe+tBJClf0OVf1VJQBCsWwtyRLgWeutEryty+rVGACclmXQ2j4P9d4/Ck357
yi0HSWL1ZqKLwzv0VoLPXeeACyaCBTTpfgeaPyCSqT9Ft/RQPzFZeDLF06h2V+pW
B0q4VuegkT4mtJafS3eARO58C+70ELwpj1q2Okx3CR3iT+h2VQ2+ay+ZTV7e8HHW
S0WL5BSETNxqlzoV7QRjuyLW99iUoiaaY8kOGnCxO4HR/UGmgfC2RRfWAuWgNtKs
VEpJkOaApLD2U0wU5Ux1sD7+uT6Nvdb8/DheHaH1xakBqAhk/WlD1KMvLvnjKs77
wY4qCeR8HY0Qkdxv0gpe6mQTlTHksYWTFeEWcHT0R2qLom7MUip3X9Pb7IIf6LGB
KewJOGDV2LZfnS7bE+ipRHegpXT2sU5PV4p753v0BURZkH4EUMC2dsaAGtQuhqjN
EfXkq05sHTR8s0xRCkQrxXmLMV4TZUjy9/2WqesKBhGZ3um4cmF3E10pnk0pcT/c
I9TrwY4WMTAecKaL9IOuROhMXeD4SeLs713JpaGHkhnj6BfacK+FiJYnuvU5nt2O
gb70WCmlDnzAxor3dnaD4l33bhyWkcOL2YcVUpiZuEBpn/8JyCtaaIDSONnmnrT9
fPvzqtsc6HMNJcGQm7e0Yq5q/ztJCmxeMEvOyGW9d4fSqgxX+ANY4r3WokA5DlTI
Rl9IOs64B4z/kjIycF5RmXpgP+DeKK08poOR9YBjapvNeDmYGLXfXk1uvaLfi8Me
TD4vyPVOsuHcmKZdkR2EkxEA1iFbghbvYcm116cm3rX8PGOyK7A9n0QNY8EALbYB
VAxILxFmiPP4698x/3gVzLlQvW4cnIKUQKoxb2AZzLbN6sCohzbPw6KX0Atw0uMF
f3j1lLIqKU2VEIZ5hT67NxIzPE+noncQ0BnJqLqMv1D4WT5ir/QZIiNCJt/AKXSa
IO1snOLrjWHtXS3sSGr3XudsNcGtDUETzDGJ9ywGJN7iSV8RHbYcwYUbT0KFhWg4
EXEIByDW1AMYCeGhoAHoZ8sj8AEsZwdx8aROn1APo/eWx8rF4UnhuTANg5BJ5lHO
4tNUAT2A9i2VynM1i8q1FEZYbCqsEGL6rXgZD+9MTCGqObdfgXlUAl+EQn/Uyn2w
zXSvZpUDK4so7j9hEps8Efm7UH5kAKzAFzOzuEuracDL7rTznwxNyZL7Ly0HYw9b
ebqYuFj/gPdNa9mlYjxZxGvkE4pDfmd4HDWk186WhICywItNfRpasjB0XFXIL2/b
N0K7HCaWfMO7jFf/kcMi0j0N+amBaO7hZodOFIElXWVCTV4eAy7mmEGfFoN5UUub
43986TFiJLy6dQ7gUgr+SS1esT5r8fKmvcUKYrk+ImVp/lJ7ojbksqGCxk6894KI
OHlvk8SeZpKfGKaofP0fMewP0KrOU/Si19lAe0OW/UUUZ4cVYCRQzK6Bl7LlbzcW
AJ9LH1FqkLTlSEh+VkqWitRNMlXkdV1HMW62EIA4q5q9cH2jWZguuzDerEWJViSa
SxmQBBqB6CoKH/bWyY8VSadkrdVO3SxE/vV7tdgGQw7EW7TQwdMArHooJYKHV44x
A752SA6FFHyD7HeLeeHYk88O2olnYdcfka6jGFVC1wgdKA5+c2B9LwlSDKFxQynn
dCQr4aakyd5prHDU29rMgQSYirQDM25OdcgkfZmXhSohcXn3nCLf4WOAyZkObM8v
V+XfZfrZouTMGBcbG5bYkiQ7SfrOgCKzg8AM5jbPmVo7hFkDjgvKmpJ8Cj4rl6gM
E11FsuJs2XU5uiAOFPk9nEugrVVG9JQqYQGRfCp+JHNtHKU1Gu/b4K+Bq4BSIK8q
X+c8IkBSffR59xZfP30NSEKo4LqN6cnFfo9sVkRavKeveaEc/rceRFRkiQYKt6SF
4ivvDt1o3xUM0rBuYFc4NiRFOKJiS/8LTgEasbfWz5GvUIxSNs7tJzKTEJQOxP9v
XqVTtNsUT8IUeR5mqhH3Yd2eVtUjjBUn0rLuqkB5R5ZXNWqjs5Ov+96YRG49cuyj
Ar2UytAUB3NOcLEgxR9F+dDdDyX4/OwJHx1sal7t5JN038sehMvor5JC03WXPpVl
dPdGcd9dsF6Y0jrVSvMGLiozv2XIX/QkdaoCi9RBGjrMFvg0CJh4rFgZsvg2uRYg
m88rNxWXd/APrpLlJTXHZq8JeNq9WAnnnLs5+/Zamj2r97QJzNdhH5MpHON9hhbT
yp/kRSstmtmAUxZpMGLLx4aZuR8eOaDxQAcearwzR3yqSXkVeKDz59WyrTFmK27n
+/RnseOk31IQGjNQF8Mmcu/1xptBoss6Cf0en3bFjdJ44hjEw/KhEz4gpVlgbTSd
UFVjYdrcBLCW2mERxfkf6+p5t9hCcenvkMbjIGu1oSCCyYFrEEi/M4WCPBb/Lf4U
ys1jEciDcmrq+18cnH4yGmsg2C5PKJb6+24dmbIqXr42Fyhz4LO0SbfQ/EAwcIUq
4N+qW+M03PvRzyN7J+Lmcu1rSo3KpVsBr3EtzJMJkRmINecHqRbSb2OOr6TMbzpY
0fExMjfiDu3EeQwBtpZTaWx2xuHw0OjHdzEC+h6mgP14y0aWksuOeNlxpZqW2QgN
UajRAwWE55r3Bon8hJmZdCGbxVkk/1tjp+wPOY66qiRHfqW3ZNsgAc17zSuD6djv
j/q3RNwtqxOSrJ0/wvittWl0waJ4CKlxLa1PK9dOoFPQFMEgqyyXzpz2C865JpxH
dsN0mmU9rwKd8Xqri/EcrXcOoz97SXLi+EP8jN1qGOahnjtjUnWkBKwSR4qcLYBo
EO6r7SCuA098+av4CB0DBT3+Zhfl6Wgh8zQ0L5D99dFcSEZoMzRkq5S1adKAh2Y7
zADxEytlfmCYgM/UmjsZySYT6nKXBE+eiT2K4aWQrObkRz7dyb3tWTU8+Cdvcy1U
/fHP2CgiArD2iZ4Z0zCEdccD/RfxCB2mX0fU4VQFU0tt305JDIgE4AmFKmaC+GBK
bVCqTP7wFr00cLDeNa8gLTmEjcepHhCh3mpztsQM/wvbtkxUvvMG4xiSL+fWebtC
n2HFEaWw0FN7NSjoU4gdwvhm5i9e8X7CzV0zpYSbt8OniFnL/xewjv/lZCiiSwYD
MOK++AcfP9I93LAjLWsg8E8jIDUVkBNYtczei5Y7bEKrOMHZusTUKWTbqnyph5l5
skEWpY8ldEbeRwuxfpovl/9oGNhViihlBJyflk32Js4bmIEuDCMfmHAm2yqkUnIU
wepxzO/E5BSZQT2n2JBgaV7dnTeINg28YBKTfnyMQuLBrhj7N/TNihNFyRybt7ns
t3AlpkS/ieY3VP8zXEyHGFt+ZUmo7/KntViP94pfJUdjYR6sOlZKCCbNT3hfRe85
8msN7mazjz2X/KJ4uzYW71bZvEAfCTAaSv+SGFPKU5xzohbAZN82fxErc+mrbsed
vKAy+R+8zW6hHw7ZYR2T8jnc3oWUQl8wPCatOpYIQ9WACl17fscBRmaJtj1sg1w8
WcxJllEz1Ke9JBOSLg4QBB32yxOiBT3Wjg4tRcYDiB/dvxPb7X4BCnCC+CfUkRQk
n+nNNe6Ju4ZXKFV1cfqHOnMdLNAi3lPXnUxx57TzEVyfdHqmo5JnH68e+5bl06Z5
54k2yuYsAJFH3KKotAHIGudUkXRkURBSti9/IAoZHlHlGmMSTNGA7CJOOXoRCQUR
uErCuDTjhezQ8/Z+VpC1I2/c1JJtFIQsNsvA3v5GXZkRPPJ+hzeU5bexDKxtWHTI
Dwnb0po+6SS1M5QaVB8ps4fHPxPXQuSaH0lpt9+iktbsuQgDjATJ5h8jIk/2EuBD
ieGNzGTmwxtCli6hZOEbVAMp0kSxJU41pPY3oIoTAfuiyYbBLd0IksDb2jRFWSZ1
RX6jSPmGY0/X7y7bzTFO8z1ONP1yjkK2FAkpuo+b7wyctdSAhBar/15LiegCrs4M
JndVB1xbywVAxyNMDbgHcJjIDi6t128GdogQjmDbEZlUEQuQmVHnOYF0hQ6XCx/W
eQFNqhpSjwB8eGtotjTOIBuXQ10YZozNKmXUFfcaNi9vBmugu40vjDKeiNJW/M+P
QG/gq1JNFH6xA3WKddFhhKyN2T41gy06kOveX8a6jt8C9f2ymfDnOYobrL4gTpmu
YCdYgH1IV2TjuSu/QzISUO4RUNFHT1opf5bafX8LAgKjKQ6h4P4OT+3VZSsOcI+X
G6BkrTGkKzl453fTmSbEEG5dXuSCGapP1+IMLkN1buLiUtCBbjzn8tpNtyn3U3JK
4MBRGALII0ms15fvVZ7GKh6pCnA0x77KCglA4ljWqX9+ezRV8MB29Ye6sheLT32e
zN3jPnEfnm/hgzVMXGEdfJMMMghLKUQK+i1cR5D6zrB0XP6vYA6FxN9BgT7S6qeF
lZf3glHGcR+1Rx+ayR66YhpZ4TjYX6/7V24jCdXN4bHs6P7axDrMjametTFjvxOi
mxXKnws38KqEujL0Ldr7V0A3N6U12HQdjSQ1yOpg8PfwGt8chqDogjktcnLzJfn+
hPIgNWftONtkTftN/BGMtZobP64rIuY6253r+p4syz/ZKiRhje9q4f/hZ06KccPj
evhq9i/Aljp4OW4gwK8Gk/LckdtlHSQYMgwy4Ncx+DBQ2MJ5ZmqwwjfazPr1U/Oj
JqCu8nPLNTTL/prWOjIvit87QYg1OfSWGvsdTkSviRJgvDWvTZ0LBVMzwKYLVYi1
oFCzlJoGfjQwmhx59WD27XLEAzOKuEptZTYU5JjWpFC+iKsj+WzGoXp/pvVyQeCZ
6jFYhtmzrtQH00opNDKiYAZv8Y9oJ7Ba2SIFpACLk+zcOZcgSXo2j8jvAljyZHgv
Hs77pu1NlHExHEl2iIFEULUauHXidSdGoabZFpT1xeo0qlkrQCAH5Uf2h87ic0eW
zCQ3cQpxjZwHjSDcwVpFwj3HL44Y+hBNCKEN5SlwXv3nxPP+COJlN07JqIX+RDYQ
C2rpKkD7U0XbBnkmr4oM5LFij7hmcGTE+6CG7pWsudSVuZIJwtT4ZfDIfwjrz6zq
dCwIP6mu5mLaEmxmYVQgzLKL7lWL0F6rc27Y5QZ5MVtlGYO2HiA4+R9oHFKuZ+jq
Rulr/pJg1CuIsnQa/lvBr7zhXeOtixZiRhdgnDx29n3ijs5gVGimAjpcPODWV01k
WiFCu5rNCPpk5BG/oo4SRnCtYKyWTvNQGyDlNxeFSFEVHAC6B1Rs7lTEX6Zu6oVf
0I4hn9LCwgrTm+742tH03nB7zBY94G4uMrd3rW0rbelMNZlZkoZepy8rcowQsLMt
eK1aFTW/7NzYsfh5RLe7cN6RL6a12fGv5LZDwsy/O7sccf3qlUVqLkWZkVF2zqk/
Z0obS2LNa9X5w5Nro+im/0np477MSNSXd1XAQ9T6MI29e5onCSyUFZ5YYdiZPy3Q
b/qT95L5WWJ494F7xbtvJWY76akE5cvv17mGDe887WnrcwNlF+94M5phJBuCloJ4
2Lnu2VM2HLCd1eW/tQkHV6OwNWvVdZTSIISe5M2z0pppzHSJAXe1VL4yXCsKwg+Y
vnWAhcnbWs/s9Q00xbdY6nfabYcIUIhhTxVG+T5GzxI/xGfpEJ/ulvlUP6d/t1Pk
ezZ14z4srcsgMahBMgLoPaoz50JgxkKbC8pFMnckS8kaY/kBWNPNNEc1wKUKbIk8
mV/cDC+rMQbaWEIof1Jmk1vRqntSgPiWPIH1AfoWRx2SygZrVT0BQgf8r+Xac3z6
0ovOwAmEEc4UlhcKj+884t1CHMQdiF0OnhmDbtX5wzqNLSmoKIqRkHrocpNC2im9
0AzWVg1fdU6tmk6sMLf0oZHM0zGKeNqyGuMLC1rB52Oc9lEMnqImbrly0ZtFKRYs
cnld6NEucnZVsVZGf42SaSQJqazMUFMBpFwshW2DYhLgVEVjyZO9W0Z1rBStSuf7
2fjM3QbCLPhWx97E3n+9iSmgRybWlLMjCAL1J05UB9Nu2C8qWPULRw5PvG4qX+6n
nAgHkb/PByhNsruNVqcWhtFY01FwmX9UrFqKDunxqBWDsVoST/zTDV5IrN+gBIJp
1lytQ5xuyexmrabNGokOasX664ijYaCjEprq14wiX5+HWH6KeOudZXJ7BLMFOz6l
yWw/6P4aft8MrFPyt0mcZcT5QgWNeJk9oebro/O+KzNGKNrffViO0T00D2FRJ9eU
gx2KhkdC/SBaZQZhmynRLyrlMa+igdbI1nqvANZh1QrYhsCR75EZ97Zg7ivXfSd5
igPUZ1fwN3657NYgk9EYeYLJCfSSgKafkcH+mje/54EwUdsEoFcKRDCCTpAqkoZS
0KEES0MACExgaCgaN9GMkKMAUI5KdjlU7lmz1OuzjP2KTbuDAtCuNsniWg+9obEa
CE0gMCxoSc1w9eVU7odcEuiovd8NfR+o0ZtK1WTYSYvvOA77XsqDYIxOFrZhFvr2
Q6TLTlm6clYpcupa2pkTjy9IROvTfJ0fAlb27YjVZtQDpma4obge6rZE1zG18w4/
rmLqPS/I7vjliuWxkP6t9tS22xJCTD26iYJ0SK1iUN+2o7S5asu2IrvUQ1pIW7LF
v6V9ThSpl4RpJXQLWKW5L8gUS7USLrKTmidxSdh7YsXaBy9H6IM1ntrCrm4iHGu+
IpXA6NnrwDnPHHLrTcNDiAK7/FoE3bZQyxYJmgxKiWb05SaazlXDayNPEM6Xs7wk
Sh3ss4y5nWA7KRVaiZ2o25FDDhF0YVLyEJ77WIRIjC0nNPBk/uKRb0rB/P+uXefX
lSLknO8gM1agQ/Z2J+n2S3+79K8Ys3EdG7rV/QdlAkJFK6+ilirhwIqxj+HlRLM/
6bIxbIayppqhT+xWrp+r4Zj64YEKbeovTW0twC63+oOkHpr1d57GNZXZ0HkL6wrJ
NeQObMEymBHgfCrZBVYkDws+APpUAXg7Y9N7nePq+Z9n+oblQSCk7GfIEyO9UpoK
9KF3A6OosxCMIf7yvCrqu8vEBnGpq2csWC0YcSvmXLCiinsj7ou8x13bBaiRhyYb
/XWqpPbS88AOOQoqqKg9r3ocKnGjgaW8DKXBsh8Ro6u65eb603tLyhCcSBFOT2z7
XQFtp8QDFMcvV5QuOegbqIij4G0aKB/wBtI11D4UVPmXaRUC3sqnbqsvY3aR6F9D
LgK16N6aUeJGW7CLghFZfYxgU4XYIlTywYMTsztMVQBzLKBzbWQ6nfMC1VW+QWo9
9M3yO0aZ0rXO4NEZGlGJAKx7rT/fqG7jWqWiUV0aSzzVtIqzOJyiHQGJFTW2I+AO
t2CTKxEMScDO392fVE04TxvQky0aDd+T9Ccezcb7epkbRW0I2rvN88DW5syvMYPG
1GOgs6eOGFWB+XIbvtO22adElDexvhkAeVjvu72+rlYxO4FyGl8WSnscW4CDJpdB
j8dX2HhZ8M+2CR2lR9vuA/uaBVZcqkHXI+HUuKvyjtkk3YqZq/1jY+ZgrhenByft
QnqTmQPrzd/f2pvpeZGZTths6DaXzZl2NAMkgZ5j11rxaCBVhfKDbka0ByGQBrl3
hrLeoHZPAbmouRIoYXmI8pLIg1/nAXmvspn92ghg6z0QPlylVdllDsNPQMRKIafc
aM3yCIS4k2KXKLWT+384lBHLzihPaDLqc/R0kbhMKkjH/YDADARxcBjHYIpM0syO
0Llhe0auc4lQzufZwX5/x/5+mSzdZT7AGmwM7eHlUkFz+yGVqqpHldYgZT1NxiHS
7KJYbfuYQzuFEbcaWnT9ESES0m/brksDH0Je7pF/mMhqp9Xo+NfzIYw8UjKWl7Hp
1nZaC1EaAAkLUThsRto1EtpgDxfsLDwhpTdp2Bjc0gLRvseZ1s0hSfpoLBNsCMg8
yOfUNhPj+n/x0npdz4uLXoUjHDk0HAstwyzhz/uLVJ2nMvlG/d784Q7SqSsajN2D
iyHNFx337xpqbTC/FhqR5rCjtNzavaVuxKS1DuIMox97gm3wELgcwDuC+hSPfJx2
8gxZZwhP/Qwu0v7n1hzahIHsV2AATwraOsasUyi7FxfGAPyUcaVu3pFeVsyQ/jyc
D5qvquoi9n/j0elTTc3bPpIgim2ecgXl+eAlo84PyowLICkQpiPQAV9rNs2225o6
Zle22SDgqnnqXjaKlCKFZZo8XNAFatgbMQIv1j1Rs6rXErsR6Rjb9bynq49YSiJW
7aZyJ3rKZuxlI0K9s1EWHSP0jdEXZpEnaicg/+8I7eoNKm87DSeZ191XjhI0+Znm
P2p0N0e7NVXFe05oPfkv4tOg22flzqTD7BJnFcrQQKagIsEvuv4q4OWQSbmFifTC
tfyEbKR0T6d2XHqWml+fQ/R4I8FCCnkMhF+p+OUif+daeAQyRAQP3U7h+Hg+54m4
kdexQR06y4H9cdR0frBm52/qw+Hh1BkFZngtIFjSF0vOeu6mMxH2GyBDQli1W5Cu
KwcCtcz2csNoTqpmpo8ckvBZsdhg/NYa/9vxSdwOMSEN6WB3PYUwNmjaXMLV8G7y
Po24M5Moqhj35gCII2dLxLSZvlZdAWCAAPSBMuPy2eDNz76J51g3lJCwbj2nA5l5
UY565BIKkAU5tjWtIB59S0FzS8Wka4EaDJGh5oasi93oDI+Qt8a/i/zFfKOuZYaL
fSMGmZVLsihLPJs+Xbe53DiTrZOEU3Fi15pIrCL4n2m7K9E0gp30WVPEh6bqXBny
xGZ0PC4TwqHTHBQvq1cgYcuDTNJnhkCexD+xb6PoJm9tXVkHJILQnH2O9w6R0sm3
a1YMbIf/JAK/yes9vLddLJ56ePP+pd8QDuBI14LIfC1poP9Y8ESD2Q26AUIhTM6k
ByFD2Zd+q2CczYhK4TLCaR95TwkSr+WrQhWZ+8q4rBiVzboihQxGhKOuE7xspygP
v7IO+EcLR5o/gzVOejIlbLXRMZzZBK5m0YvSQb5+ujOXER4S6qAnCcluRPtl0vRa
nFTDfd+Ix2W+vil2JOfIH6S5nPcwFIvoAI/wK/7ZpxvFpl38iLDER1SLcRlIxf8Q
389YC5Mb+ekGxBY4FL+nB3QEdGH7m5olhremYdjJ9S5EyapUTAeYk11REeiQfUfy
6arPbqyyXAr30X0ZX+q/HyttXNDVeI2nbgkhjCUa9AngEh4uzfHz3ZkAtl54XHCY
nzzjFKed+vFdZJ2vA3RWNoci5lgtcz5hYj28yH0NZSDt4ZG5J1hKt3iUPsauCEW2
EAAoNghtu1X/fzvc8D4IcSHU0E5IZwqspqPwHPpcvtdr/yKrRnCjEQDMwim6DCaw
qDknCFRtDKqc648ugUu7k4d7jW9s0+WCJM8fKoEaPbYVRAqrLytYnNLPlv9WLZNj
806S9NuIh15ZvG0bxAJhFWOKlxZmjX9pdXJ9m+/hI6d6mmbjG0+AcPmKPRW9dnj4
nGl4mTp9+LduZCPXJAOOP9HwV8i9tuZ5Hv3xOUpbTF1xG2qDIFY/Gr3X/EglgolO
A1rPkmxeZ3I04dujFrfVFmLOJL1LP9OG3DqvmeXEtDcTiwy8qrpSJ2w7WRAWdUye
qImBjQndcxCKk+Z96bQnJuiYhJPXNHrN6UhBidwnn9cALwpqEh5zUECXHGxTeTTf
KpVxWclTC5BVkPfPPoEZOflPClftIXowdloxpGD6SOUFc7ZhNaZeFsyrvfVcAz/A
KB0++TFiHlASmr0qhtAgUgfs7uhUYu8FwUgKcYRlXaUF0kzipgk9AshePA/Vgzcx
qyvE1E9zYGccPr7XXN/FYkuqXl+cIhKoQCIGPhcOx2NjRY5V8AOyM+z7/GZE2/Kl
c0MuUL4Vkjh1+nKYUm4wP/3AvDFZGBcCZPRo1Q9HAbkQ6WV9RNLkbkKQPrPgXYVv
M8LehPU3Q0wM7VNiXX7W6tUbJCbKE7fjgRaXreM0GVcyOtqkl5nfgac2bH+JWQXc
gJyW5wOd6cRpZm2a7ia/Bxp9ax0DLPTbm8IXkhSvhWeprOlayfDkZaCmU3YmqoWh
+CSYFiFkd3DXqkB6j+kKrE5X2G5LsDZMLZ62U0U+O5ZHAWnUGW7VvsuwRgyZXZOi
5ajCGGL48nYUQ2BUfBo4gmncwOcUAvgI/PD8ixTPubTdPQH6pIZ1CeVoUzv4QWRZ
WYGkoLOgsREOPr5tRqF8/i0ikm0nIXuuvcAmhjMSlFrr6UVLpVSHKyYk30P0zxOj
S+ozf23xNazt5F/k0QjDEf9X31Qn5SfQs1s15C3RJ+1Fst24od7ZuwLeD2NpN+w1
6pEL6GuV4A40rdJk30gqEnf/p7hIR3hfmUp5Qt98SLbrG1Rq1PBmneSoWmIk8B6k
ebPy3GEnH0lYuScLLj1qcF1iniJAyPZoJa94UfZ+eeas6t7VoJsD7bEKLmFtBDci
iKfJzNsd2tXFllxE4Uj0Zp09Lk0hQSt8oSOMqiT8NTm1JLuCCSz/sflr8lmV6Z3u
xbRhe7MNkZ613LYCCJ/q4mtWJaU+RqZG0xtyODKPvp/733hozwA8uMSg9Al4kHIp
mJ7fK4/RDaEWkBB9X8hxrgL1Y9g1Nlsjnxx/bmdc8+N5OzrKdK2dJSiCqf4jURYn
5Rv6J5/WiabgoNXdgGfA/b645E7FKgJvklQPKZ8TuXMKkjfVL1Dha+imyMKjo8xF
CIsx82rd+LsTM/7E2TfnRBAN70zigCFtaEacfjRMq0mjbey1tj1Su5KGYCPm2KYq
tN74UUc4+ZoOXB7j7sqeOdSXZFkP9wllMPiC/p3YJPtd/oHEAqps+FuhLexhxAMP
KWly7mysLVDg8MQNBb1SpaXLyrfUmJ+m9j1o04W3ZTUfe25kee47gvWTlZV1POsZ
O5/UtCmLRs12KPJcPs1ooeRKZ5vTkHnHjZ8tH3zarLOQPkgCJKxJY5eawAcsOxcO
ggfe9renHTRgGQj3xtJ7mleK7g5arlkgQ0X6MWL9yTB9lCUHb3aqQDd8zINJWxUc
bgjGsO0PxgF+FmAwfzFdv2KS+rFWY9DK9VpF9c3QLzwuUwjGL69YWoTsNdIHdR/y
KhP+bZaoH0wfVTKgqPa8NggsIMZOBQH5tJlyTlmg6iu0ClSPZWlZOtkedt/WoqP4
AnPf0Bre5w+KOtG0BShxOn7I46SFCc7RXDyiTxPUs1mkPPqPBz8W3BA7buqKHh9D
VSbXTfLJ/BGRIIEDd5MolygLquI0s8D5llZSYgPMYCluYpGkJXQsyuISgGGPZpX3
DSbbIetOa47i8PUtGkp/wIzOZoHqG4BSnS0y+/HmJ6+YN3uLyXZYV/fDCii6BcbD
Lvn3z7Prd0e/cTQgwTCLcaPdAT3MWsFnkNmZJpsGFiPrSpM2EF8MlyHeeQw32vgi
6jJoACfFm4VQZSZxogZzU0iy6FW4VLspiQXC9UAX2mKPvGu3s638A+fv4xZBOyNa
5Iobb573r+aT5eeAxVzSeJxK2WzUQEqSDNa5frm6qKaFLsG9FG6K4sz5Eda0JDCX
/1jt1k4ZHjtKqw46pSgRGSu30IjP50lOpiqBhJQfRS4ryGisvh28j2Y4Bew1P+Fh
pzal+Km8Ykw+ST/UVv1Pokp0BTjE5lEAvjib/x2v4l3y1oQj25I8QHYrSVXjU3SZ
BaD9SLGzmg8wv7slFRf2FNu/CezzCPiPtQSPUDMfhsj4yhrtzrkksaM3Ezz2Bnxi
uKgpY2/P1BQVrXVYPdH3kDmrKKzk3pBFrH9akx/loiK9xWv2cTr0VMycvSgUmUGO
vdHIAtbnNvR2tS9+4OJuht3sXiup7YAuQUyrUhs6eBUFXMYaslrd0hssCaDN3K4g
s9rIsj/0IHiDpXC3sRnbK227zhYZld5NvM9hC4rAnWw1+sGquqoeoljb0M5ZF0gZ
sAUpJsOf+i0u+rl4d2aBuSYpAfAiabpRnlrDLuwZjlwn8RS6qMKD1vV2s+Y/IAXZ
HizFLtlZUf9PKlMEWWXOihmrU+9phRUAADDXFHGXGK8Lqq38CeT+pH/awmXagbDX
4bybHqckHs8LZE7x//UDHoCz16nvVkteqMczdN1wqWSqZOP0R9TjCJRI0WPD4smM
avXanyStsQk32SEtGF6hkwntG8yeiN+PrHydrsBculg/bnP+Mva4XM++3mw6C88R
QtZH5CtFwJAMihjfPWkI7jKv1P1nJx4iWIvRtgwd/RkN3QZIsJaA2bAtxdKKmHaW
7TbP4UjmfII6t4hO9HnEVwKNHhnKlfVCYHguys4XbVOKqEAip6TiqHBReZ6StMkd
lbEuO9iwKemtl5uC0uVZz0l4SAcfvGMlV5coXfoaTSnJKrb1UvRgyEGM8H5TVQE4
oolEIZx3J6+QASkSvOxsciEYrsN/Ldpa5tee+cGfNs+Mn8xG5OhzRRPxuPQeRWI9
fVyEL1ibptt9SblPMjLwUMVLplkd/yM3fOnH10CCfcGTa6zbYv/tfNtXrN5v0hYz
UXxAdgJ/GPwsTroKXcLtCOKPt3tGJT/82ObWBw9MZomtMXpkEqg2ZFB/lcbnvWnJ
blTD37dCwBxeeXRrTUODx/Sb8lyUujR3zR60vtLYud7JH9WXv7DBcIYKqxNEENAX
TrcY2h2D0MA+Wiq1qfxElmPTgVeaEjP7ynLnVTS1b9ohZRRGgUTat3EnHuluW8UT
VEkxBdvvlMjzOjj7lk0ls7FpGMmOMg29hWWePCjAjPI4WTrenDSpj2FICfTkQpNH
7BHCSleoIy3UOOjNPSKKYbN0hcLg7Tf3idWzoWOOpl4eeMlcRC/D8+dwJxI/XZny
BX1mO4TRBiz8wi81GCfJ3PHOYcNqZfMdVdnAhzmIGcphmYaIjTvIO2knPpFSpjsN
KY7Li5+uiUL720GyQYMcjtoWAXGs03GLk4oiF04fVQwomaAGpa4S+RAm0/DCnjli
JBBEnSFyuzrqiFBk4xlKjbG8S3hWKzwwnqzmaFmcXYnE1hbDylaiWPY52o2TlhQB
CP9T+0gVYlDSPgvt+fdj+KPRYW8gh91Ljwo7VJ0kDAoG85kg5eblEPcTY3GAQ2ee
8LA+PLIHuSSdZW6wLEwlDA6QXHLdXY/akCEBC/DcvuC9uRdcV14vOconq9GPAw3V
9jpLgjIcH7vOck1EK2ajsB56BbpLne98jHgDtBsp8trVfs1LLYpzrvQ99a50mDmm
eiaO3idZNktMslkEfI0D2S0cqBVhHFc1mr0kowb5xaNtakGcLhQ7djyc7y9/GCC6
WfacI8Z01wTWShYgTF2lCiP5b+PvzGYXipe/Xv4uPmB/m/HTpw7+ki/h4vVEuT7o
7gv5ECaA35SmUOppnAZw0a21wJ6+fRxpXwgxZqQwDL/S3fKVh3c7n764dHvcvRC+
ycEukDP6SWeTt5RIuCdLOmXw18C1M8pXm/XhPQpNzs6afkmQ3FIUc89WKiKn3bJY
gAtq56kqrwWoeDIOsJ9OBPI/Rx+ykhhflB8C8JsUau0sGVDI6gCxJLxjIBsOBIRF
AWYd0oDgPjz5mtmaEZdPaAAF73YXXPc6oZDnnCNIGh3yo0IgHyMg+yK/e2iuA5ir
2CVs5xj71SGLdXuPNnr1kvfXPZYTzLI066Kr7QoHCL0FSeLnbsBwvwvnlFaM8JgR
55HZb1WWVk7fVbuU2gn+4wBfLU9gfwy4gG8bdey3rGp/yI20lUdB/IbFhAYmiAZW
MgUjyZ9CZXScCvG/adwawe5UChFzIXNOz6qg1EqZwg048NM4iWb5pEk1IbVbcrEK
QtMTiunHjl1d+h37/SFt+8D6GqX9C2EK8gvTRAcMxeKi+PqG2C/lalxogaSEmbf6
oNavUxbFp0xI4G9Tmv/Gs+nBJ7Ud9XvOcTGWKJYdMRXvfH0w4ZqSFd8FcJNXyldI
yaMZnbaeWW8/eKK3/Ei5gqW7+pTBr6nh03E+YwMgE5e82+5XB/mEpVeePVHKK4tm
xs35LcV8DnHQrHvOoxwyjBfDbVo0UUzaAKdXXUsp3EHTqKLvF0iMkO01i92/tsC6
dGovqSwGT8ZKeG9eDwRaJ9uC+kFJVq/k+JMav1OSGGxcECIO1fT05ytxGBgSXp/m
StYEjT4EAigU3TuHe2125mhcYRL/1uJEcTzuGeyBL1JZ3DDyHWjDtksucgciFQu4
pRZDWSYg78iQGYCcKNEqFtdv/aEgcTuoerLCety2wImsNUxSY1Ij01CMS0SQX9ZW
sMeelzAUUbv+IEjXGR8wbihEGxbSD6E5kHFgmHbJvHb88HHzN1HEHlntnVM3UURo
JHvu/cUvaACdcFF/W+3LUqXzbfKgQhrdFa27RiH/gWxKIJqrhcU6uWZdj2eeProA
qRddv7HNtkesp11qQbNNgsW698vNWiQeOCX1LAbKE1Y9j8xyN7EA8agZxqXAbUFq
5RczFGoP1rT9noC/vFVR4u5WLjrsjIi9C8Q3/S7w6BQxaRspPwEJ9FLuLp8JwEvU
AYu9CVOYmRBEAIuT5pt2aMW5n8tQi5pZQDhzyaCg21IAu47yWZjS/BTyRzF5zdpW
4O+bLZqS3iaendUN3eQ+TvGT6BCVe0s9mxfVU+IH3/8jVFEpuMcvEwTvNCfVwmxs
XrEUsWrjP5nKsCADOcvL5lpnUv7em9qHGujAOS3KqMCA/3J3yZp9VBvkWia4jaSI
am1YKeCNFkbyo9/T+iks2TkMenPB88GzI9+lQqSW/Knv/zkLfSGE7UDte8XlLinX
MwNDDr8wn1tg/B6rNGN65rFT+RY05Au9DC0kr3tWouvlgAKoz7Tf6KHpkZcE5M+e
il628pORHcMMeI+lWlSQa3bW/tD8Jhfz3ORWb2+o0ge95H72q36+WXXFi8ZuiXYd
pRdm6MwfXYvX/BVs2x0vNguz9UMLleT4XaWifkw9wL8zbN8DmkitApW/j7/AhkuB
kqyHEnXAzF7XOCRjjb3M7iIgKqFc67N+b75o0ft/vAKfLTjuxm9HgBBwqJOfZFDW
l5tMNGc1bE5CBJje5HmJG/j41fsFQs+dBtZfOXgGRYst3PkXUVfEuAYikc1H/+BV
nROXuMyG410MiZpfVJNgssOJxhJk91L3GpY/AkIO3jxMl980jgw25mIxTNMmzbCp
fyrpgeGpf/VC3qRfnavLGKwHfIDcpIJHqrAPSStigHdXYJdZ/TTZu0sfeKJnbEjV
nE7crk49l0zcdHd3sk/rI1qTcQsBc8tva7pDSUWUsYIHVK61kGfHVEUPpSN35Joo
5YMy7uk3VE1Ys9wg96yOnruovmFP5T+uPUdzrGlJxyjoGVCOuH00y2MO+cOJtIs1
O1cbI1t4H5+5dahRM9c6qk6KoLDn7NxMtWeEgEgRS4UOaBPBfQBU8BggZlIChQVT
jwUB/I21QUGTWnySFvX1WRwB9Wy3qj0jJlCN0kxaqA4cxH4YIQfu2JcEq1MqnGb0
MXLv1HJ3o5M8j7MLjTsREHDzw5SJv7X6TKedfVDr2dVMMmac4xU0XrWyZQAyVteV
RGO/Iy8pJ6svroGFPf2JVtpUCibaamiq8YoX/MmWAtp+I6UDom95qX++jPsvmsSK
ScMXnRVW+yd/phOkxBtlN1b6MjJogE4NZvsgcjhRVd7Kx/zLx3BSLqypvoUZ3oMU
QRLZilqrgN3O/RVRWO2aigE9D7pwF1Snq/YltyuPqhOQXwELPDKsMyOq2ELUh6yg
pxjUlx/PMcYduK0qlbC7JKoxvusk31siimVO5pozzPnhOOdY2duVzUIed40E1vOb
ns9PvM6JawDcIyMz8ieXPz8o51QcFah19TEWJB/oCdr1Y+KTIRKgklu8KQpBCk0m
T1U/+ck2qAIler6xaK7FllefKd72mhtBq9pAjfLUS90QGkUfGj5tYeO0QTtEdb78
eUYIRCZSkhuQso3yJGHGPBgY9UivnhpvfTgVWgyi5Gbp1G/jlp9sg6BLsEf0k1Qy
WhVGwFlPejdbpShkUkgWImKmCEywQuxaGxXKi2zacBjFFNzHlJwknUTzxq5/2Bs2
MXiy4LCLf/gZ2S9q2qlWqFFEr9ZXjQIOsB4ZDsZfI4HmkzxmmVdErqVQnQd2nT4I
LJ89PjyEOtBBY8CizWqdStXp38aqhskjgLB9edGAhlGtd5lpuNC0NWMHaVO2Bwnw
xiLbGYXJQh3//w0i7EKOQQus9SnIX0EvCEue/Otg92Hz3qOC+9Nlp57wVrR1m6rx
3aH6PGc063CaREhI0kGWrajSOWlnJZtFO0Qgjzg/xVoPesJ1QYqtpzse8C8iwANz
LJYwCrafYo2OUXonzpKP5b6qa3qShUNxN9WJxaWon7oo/dDy7c6NTY+MZPaC36+G
R19Za2xY8HKAYfUkEGN80prqMCwTQTB+DO72i4y7upwZ5Q9hXW3ax4V6Fwvo8QVG
f82YJaU27v6QW4CdjlH9DjkQFynVgNW+GplHSCDgJu/+r4NdPEo9ulcaMpS+MzgG
hBAbD+OzhTO3Xeqy/sQXXkBYsoDZpYpgTwRBWxaMF/zhFoFhR2Uh+qi7C1/csMMP
3WP0ApU94UQRO6gymHGVb2jw9QVKxcF0tYi6wO60oFN5VNF7tnvuqcyCOP40qo9S
i2xfLEXlZveyqWCXEsThmL6wKUvsmegOnv0RLBYvSJphorxI19z7VmCeuhVnjIQP
+NOJcCVOpg93QheopLsZo5pHUqxq1ABxsjQZFUIdHHT0KCxiB1oa4eDARlC/5LtO
TzO+EXVWwPxm1L9QOj+5OKgys6U0ndigMwUPgsHrppp0erXQyirrpynkHCdYRLVO
j0U93aluOKZCa3290x9buDTKuHPWxSM20QJqmegWb5T40p3Aktk+5rXOLiBxkC/8
qKJKupmu9RcR3wf1IiquAqasceSQtAAgX3UlIqFF3GSd1Fb9DufLRJEVY7spsSPB
AXEHc3IVTRdjfd+8MEcZCwXtMkHmLeQd25e5jK1QcTHml7HXPpyNCfoCf0lF7Rgy
EJH+LTsmjB8ui61jK1kokzIz57EuB4bXRuTZPTPAwvImHwUAUyMHIXW89KyLm7gN
ShJ9TxUYjaQawI+iMZmXkcHwG2ztlsaPPUhg2YWt1dTKHpEGMxCy1ZDC8WZ022SM
URWdaOcIcNEHBPaVgFtPZu/+Pa7d/k12m/uCSGYJC6hr4yBksKFQJRQdBguyxiRL
T4D0LMp5BPXUmV5yoebP1RjqEVqrf8WtDFp5q882aFMFah0+ohSq4KvIMk5LtoEb
mVsNvC5qhcrWRwwy3WNTGxBN6R6d5NRz359V5BYFgDqlKlyESymNFEzwm7NM6iQ8
wua9BhJD6tp3IKGrONFwgcv89dwnh+n8Y9bfIE2Jdxt0OAB6/jqfMfw3v+4oOc2L
M6KONVbIcJgFVbh6eGk+4Fia6mxqdLX+8ex83Nr4nqvow88hjJNrn0efAajk92xH
EThg8k9tq40Cg8jIZfHe6Sc0OzG1STau/xVXbPAz/01BxCV8u4hV+7gizO7PZoES
ZYBNPYwo7ycinM3IY5d1444td2Q5ckO2kR10JdyzWn7n7JqyGF9HzuFq02JMuokL
+U5A+66EDcdhzBzvesyYJ2Yeenn1hVcGEJOyr3ChxGei9o6PDSeqbdxwtTPOgYbe
6zu88U/YanB+6WSjQMcKYwax34I1gjSKN0GXysTFwB++NM0tHFgM26ZurU8FYUnZ
BPh5dO3I7CL6TU8FEmD76Gf9ehqZrgFZ6sIUo8orFLgI8AkeGmzkEnO57OVX+H4R
LWCC+XK5d0HREGpN2Ol9vTLSUTRkRGCOjPUXG9I9L65vmf9jTQS0uE9YtCWbFALA
9Z9VZn3nWXgy9TPzsROf0c5BT+5o7RzVWasiIAMUHO7HI+PLs55FI8wopkm0v/PA
Dmdg6aqJytCdKY+R68UXABGcAE7ivW4LFip3lPNj1zewOId3wOR7SMFqCqRK+Bt9
ERYbu8q6tUEf4jZ+Vmmc9aB1InyAKegYGmxDuJrruZoxvR3uzlelImKRokoQVdHP
nPdeYDrOdO5HRVuZ6s6bAomBd75SyNUDTBGiQhZ7YeE2r2gQc5MRjYpZev4AB7RP
E1PQarqAy/k3wXUD8fG/htBW8T2TJ6m/67jJWXVpSPMgJUeIkS+v1VftvaDcM7r1
Jrrj8CnZfZTr6Mx6pzJDVoTPOhfMm3bEpZNhM6+eSNxg8BMtz+5uHwpmG6RJBVb4
xzqPuvj/vJufn3ddYCvlSk8mnv8EKKa1bwFDMRsiCawhzLPTSuNNHtPODSmzM2sB
V26cMCSCK+83/FEr5pSqiblWntWwCWbX9ICL+6TIhtGaFba06RhUqJ/zhJ6tdGkE
ipOQgozX3El+zy79QRmRztjRsD0wtX4mp+sKUtRBdrSZmBmehp0zDf/d7Ot4UGvB
scjcHQ4FUnLh12wQnVCuoRJCmOgkNdO5qlR7flR7lOcO8i+submg+x10jLvDuFZG
vfgPmYTTeg51ybCwn4li6/0l+0AhJsQDxN9n2tEyAGv6dktFtKV9n//+447c8sHK
v8emVpw0/Bg2WaqDYdFYngBOFNQmHc+ssWS0GiXucHQ7jrHr1x38zauuKNnXwprS
MNa8WsMXFbocJvzKju8YW5tRKnn1OSWTyJ21Ulw4/wEjKqetfAirRwbKAcK8DOny
DS8jWnsVWX5qKeTJ/hmPJDwniASUyCSNvc2H1bYF9n69pJt0Ywwk14PgeZhXFTIb
6sSthJZ0yLlTchXnTJYi5PpZ/Xwzc4LVb/WGC3T/XRHeUETklxMI6lezwI/bVjd2
6xr8JmYlWGBHSs8lFfhMsAO1i7X2tEUCMMk4F+d8W1OKVQZHHtlDjw7IN+P47o22
c+DBZNscqcGOuCMAmuh/vZS1FIeEGxjaasBGhprnCncy65DpmUAEVf/PjHgr28PQ
4domgCnJJ+owfZRDmUPigT8dc46ie7Z/ntGONd0Wdha0NuHFB2NQQFFnFOlJQlmo
LlT33Old8+V9213YoTr0NVAWYHBQGty9+7S3jUBJo9N28AD/MwMzc2FmhNh2SufF
/nnVYr1Iv87z1DYfucbbGSuSsXfwsiehxN5igvUGVULPD39OfBoOl9qHlTLMx6O3
eLZUCmppSNx6mbai2r6VnQS3nXWaO2hnO57ngzm7V6NxQDPvbOTlM6l76rNHVOag
yGmowLDQA5YbbaJmdVplFdsGbHGLNRrutRdwZDeuE8NJZth8ZxizP32WHoAQtbOS
M85qGXC1WH/HtSCbc0BPlrEY4gy4UVKpsfkBTaw6i9nXl5msMuapXroHFmNlDAAQ
hOleB6lSeHujJ3dt4oih9bf0tBKa4J4MqCN/aIVRJJOwbY+vj5awL0RBxbDQTaSy
vjBLypHOg70MmDoICjBUyr0dkMdLuGunZnk64sNXXzuPYGHPDq+bqvov2EyulJ+r
jP0ovty/2XFXvtKRp1KucsH8GaZ2Q56+1DHhAMXyfCR6Ur7+9OCYjQS4RStM9qR2
ZwE2HJzDbHd3lWA9AnaI3kp9TBhPDooWqc6ZqbFShmpmvDtfegTRFmN9UUTheHHi
t4Q73/tdIqmnKIzFVin1D1w4O1qRHIzhKHj4YrGoNjrPVAivRqintURxtokfdxRl
CpClmPoRl8geWvkdWZKTqxz30VnDXRKOy2UnRyVwR0kD1D5jzCv6zcTVYuAp9Jpu
kC3UImvoDoPzk3m4jHYF7l2oKq9zh56JXWLPMRypXgCX/aamAdPDAGQY6cFyEqGv
aGa2iW7vNqMglyPojemnicGYBXBpyZrNm2QjHKuVF3NTLiNHy8MSDb5zLQcIijAR
M7dxdVDp1PfIyYeBMGZt0kk1VVp29LT7JDosUKNZ6DNFyyTctVN5NVwAjiaC8Pbh
IrIO9i28JYxkmEZh4p9QRh1VQqlE0ycKqCA9hG4OsI1BEw15h17qppw7FghPd3Ek
sB4gVAnhmhakT8XUlQeGCIN8KUxYe37Bo7HAVUj2JLIiQnkexdQ+Jx/rZux4i7r3
52NSM0yrL46S3LTIa0hsjY8E9Nh06dk/ktBcl8OOgwV3FaRwmE3XQ2V1/bSFIcrl
VdnRODGWsy+3zgL02utXnq2CuVb5GHxin322yMZfaTmzsU0S7JuWbjdVY2BXuKwr
NuoFMzXnSRhbCMYD4MIGDv73Js3goS2u/6FlsLwcj1rAqxAQz2S9MhW65x27cBSw
hMQi6E2kxA9BmQaZi8ESYHk2BdwbPtw00YdP3zDeeKUuQTV786xUk88c7puJTzrj
R2gBfoTVArvKOrXmp4mjimlb3DQKAOnW43iwXoyiSFbPiMF1MKUsP8IT9C76z7OY
uqvR58p0Euy1A73bbdPfJF/sQX8Ett8Mdvm/OSF2tgMLRBJnOvUmlCkeOXi8xrkX
9UScZQXTsqyQVKNkCqSduMrhxLZIw6vC5xZcRm6BNUh7J+lZ/qQM65vyIuCbM5WS
SDnv61+lysLNUAVHtssSc92uwHQF9m0HA60IhniG1q/m2ScmLx1iiABbhcVWr65T
YyKZc8rd8OhdzWx6liQPZrc3wV0ObRu44QlDXtsXyNCfSA8Xkn1fpNZmqjB+okhf
PVWolhZECc9d6PXHZ029pELdfRmh2BFhuclpmpo05g6tYSkP2nVQrcOb98HIUOTq
h4y38H6W30n2wBCLOIltal2zrMfQuOyNyOjcXHfEPt4sQcYoTmw6yZxf2/KqxKqR
TaW+6ROtlUGIBFbNzyhbmMUDInuElp+Fn4SA0q9wOs4e+1aa53zVbb7KnIlv4zRg
6wJyeq+RMVHJDGwGWiZsCQTxP4C4gqVV71q+L5cXTKJ6eVt2nfd1z7UURmke8ffb
6yQujJr7pBcs+3Ur+UYuOqtk3ZlUqEJ+vcru9qIXUdAndTHRTz6F8EUNfvYWwF59
ms36u2zeuKRj4WiGtClzml0/qGhNpDCCIFgcMSuANGkrO3j4c26eQGcirFGa6izX
/ykqYsPd0y2pqeI1l+rI90eOwPZMPkCLpQmssxGfLBi8g/0S6e5hizbP8JTZzL9t
zR+Y+u2MHe/ggEVdQnSQwZJyt07LSCVV5TyfueKi6OjmuAm8bBRpf6U72FRDFGXx
txhS3QCkBwUBSOBc1vhuqnolqAPEfTkSm1ogNwZSHkNVhz5OqcYIu5KNWMiS4CUU
XKdbJydkbktJ1eBt4kuoa9HL0+i9sK9A/wbsSQKRFjdDSVUbh7obNs/Qe33bqOAP
2gkRuawaKG+AVbOoOUdQq67FkX2RH+8ETHlTWC5cbYqaSP9X/8WOZ8IGPg7gzDig
tCKiPfneKcWb/KWcGtwfZbBnVIdCmopw0gsnL4MIM7UYLwy47XINaEhoc8RdL/7i
/OMHGzXsqUEenvFEUsep36v8FihuWE6EhwjaZ3FChee31vvthBJDr8JKhkPVtRbL
RTjD62eTzBfQxP79komCgdAAycg5oAZWd4Dg1A1DV+LmCrN51U2VB6n8axE57bMc
xTy5h6Ma8Wpi2StaCHwMeHVvsJLzkoUl2roA6CS6Ruk6JituKpVQBp7AsSFhi9e3
w/IR2q5EjhyfiDw4Sj6qlqDsZQSzkaDfmJEzFd7Xc6uj6JmryC7W3WgiTGqvbqr5
1SZ9euFrAKqL8+oQ0xF8aIIqBjnYcXwlMZX/qair3FtvA5/XcX8Yo+GrW0vWCvwg
6d9ZThgoTr4bnPXOUsQYpyQMFuyQi5IIprPnIjF3GuG0Y6oyX3w2wn1gxNy1AXDP
yPB1byJkIFREQ31iTcAxyzahRw7Xh3KQIj90pQE+KSEV1/zyS+jg2c1wEqoGiCvQ
gnQp3GSVfGdFPoTFVxe+X/37SwvTiFVKLhOZ9bq0+vBFQY25MNdERX27NtNyh/hn
ltckSmbhQloRRPBAybIme/NUhVBZjB8VBykokzEq+2rJoZ8O9EOjo/OcUiAeHvBz
ktq+PT9M373c48mPhr+m9jpkhBjkMBgKXpv05EdA61ScTkUqbiuipDS7EYDC6qf2
JmZ6QTcs2F92AJUxryNEq6YtazU+LgIbf72fRPu5PTJFJASwPj66hKxZtiWVbRXh
Mj7ADi+SIix2uKhvmI7rBSpVnuYgGVYlZ8uvkxKEUWkyViXHmfy/E2sAYIX/3m+7
BxtFxrflw1ITU5pj4IGuzSdjimk0XdX/ntJOGaEN6KKa8eqh7059uNsvVz9XpqA8
T3JTiIQx+1b/DVvW5pD0kCo7Bndld33vzu8PZz7G4xKzYHDxLoF0mB9OHI2DBgTi
QXDALVeAiVQXZFghvzv5nR5J5MMcPyi81oCnCGpyxFbfo+lwcF5kBITRDUj/vdKb
iDVp3YEDVBmVkCVodaMZqGVe/KihyXjpOuxYIsBlfc/Rz9QSNmia00bLb3eFTBUz
+0siFIUc7RSsCMpNOeH1BYrtf+66d751tCGNEXzUrHiWza/Wb6IpDWRJAdC6N/pj
7e8tPH1CkstFuOrUfw+bfl9rALhBWPPz8NhH8Vd2cuq7tZrzkZJW2GxlOOzvXIn9
JpIoXcoQYRsUtXObOdIv6ENc0tTq2M5Rx3RU7nu71rhiDGnk+SwEy6nUEp97gMgM
iHrCm8N0Gds7WUFHyXjEd6p1zb+LB6qfJ4NL3d1sGxTaXF4X6KSf3Rhk2lLz9mwB
qwpSN+mUmpJSFze/5ktGLHTF/X+5g7V+jWo6sY9PHLkw9pV+kXcht18luJTWUov0
G6bw0dLcKYjise5U+s1BAhV3FB+ofnA9VutKxh/IuuYXzVVm7VBHNuJBcSNo1g2y
PBzWKga8aXHZ566WRVcoSQPpWR6J6/P/x0D5FBGwYNRmZ6gdiHhMaIRncCKvLIg6
rCk/U6xrw3f16ipkrbOCiyXD5w217/OI0Znz4VaRt/zHqeubhwBBomX5ZFPmO2xF
U70MsgyZQteAWpjNZQU/nFQKk44voBCEkrTo7To8N8NvBhallYpkJu9INlngYBY8
I5NyMTeqiTFJWDSJZoqgg7sqW/V9Vzih4veg0eBJELS6GuopB/tf2XdvBmKSIxb8
OsrAMZc6PBwqCJsQz9Wk+S5dgAAb0ImRNLgSNE1tjuDowq28Ej/fV/octBr1lpUq
XhvjZeE60pCYOFvijwvyvWnFYDzD7pHi/5SHLyLswaASqAfZ1/cV0bRSjZYSf3ge
75+NT0FnZPwZshaRtNFuywbEdGkvP4sN9x8mI83lyr1DuynDeT4YXTJCsWbuefe+
SUnMmCzUHE+tkT0TRrIyXQp5VFHESrte84NVXORhF/BN3iK2JIgX4dauAYD1zn7k
tA4sRT60PYj9O6uM84KOkQmMAy9aEjSM03KN9+ebO/GBDL2nfCBhuqDJr4k+fUJ5
lOb6aNzwAPw7yHenK4hvHezcW9AnWknpiN1pqxtw+0BZKUi3bwMdYLhzDM8kPoxq
Y9RT6qba0ROVA5xy8N0U4d+j9e3oYbyiy/unGBEztFN7NlVrS0UFDp9PTt9Zvy7Y
pxoXuY415qfSVnhVPXMwusVU0JHerzMiKvaV/PKWxEOJlgxT2Jv5fzMPwCPj8uen
xmH4PAmo7POAfuXan6PsokIZRBvjx31I84RouDLUj2Z71ZLa4rHypTxdd+bi56ch
EieTjrE/XoRs5ID9Ie424BAox3yQkP9GuQHqOgsYbhbKhfJ+L2/wuNDw4CEkPNod
m+VJ0EpzundSEd/2ujky6CRISy5HOELUnHg5SZZpp4ZC2HTh93sLzMtcw6FMUZV+
eG8lfYAs5l6Uh2os2MqYfy6InIGwzd0UAeIkDFTlMkN0NoKAiK7QS0BrR4MmIYhP
5JcmAPsGtqfpz4VzUPaHjwVQQxysVwavHhYLoh2UP1e4/zsjv0wk+yOdP2GbrmZE
vLNRYVrwer+N99Rd7zPge5+S6kdVxal3638s3nI9dhY851MLWuy2I2p0KiwezBWX
XXyKr7677n/F3EkaIBuMnIg5iR1V9lZHR/uUHtTlMCwimMQS8BkTZh6ljUV2z2Sl
g2Vh4TxoZDZrjrIbc03O9Zxicz90MgMgSf+/1pkfQr/tYu2nHmmp49dlxt8wxy63
62SBjukyGgPuUg51xqN3YnLUZ5MmVCGbZE6mY0L32a0lN0mIGntftWBNBuvOz3uk
k99olKiipBI4oEzfOs246uVvFMwPhgh6iBNREPuyowBKZCq2Tz/Z1CJG+LfRXTbM
yI44bMucg61Y9SWHZVzvWyI5S7S0u/n7MUnuMbk8ZNY9VMhJ3FPFFW+9sOdb4t2i
sbjRrJmTKizYneNMK4CSm1eRxkL9nkKY/mCGjJD8LBMrCkk9ZM+uiedpcG1N9MPz
AEBfu5Vf9gQ81GeYJa8avuwzzVShqFo1OuzXBUSV2VFaixO6TLZhHb2GtRx/2yhR
oiO5tqzS8Y7/LF/eVtSVLgJ0UuPZpe4Ly98lac5+heIlBysrXObMtDsG8Fvcq/QP
ny2ABU6qI0tzXTIyODCQy+Zkd8cjyzp/J/sYjW6Kh33ztwQUja8kRGxgE+rQUk9L
NV7GhXUc0k3Xo4EHhQdKbb+yJM9zhFAe2xf6saPf7ws7/htXWGD9g5fFG6iI2LlL
mXy+ImfZWBiwnNclAbXUGXWrv28R3e8H2bKLVao+Ipxk/wQm2UiO4+BrdH//CyQX
h5S1K8yiLvl6bb2nF+fndJaTyEy/wjPqZ6n5PIqHUF6oaTTb2wnUuYrDzYHlP9qo
AyY9msl+gnTreAdYOcM503pF8PqyyxPS49hJmw21S8chnmbgwIoSiAOtvP8SgVjM
5DvvJHtG/oZ3JGqvETIhzzZHglmGWSLtb9oGJi6vRBtyE94IxjCl35Sv3lYWTfRR
XVK8V8Rw/RF5RoTIyzGv10Auwu6+SchV67xmk05z8OxvIPKUqhobTUHrqPG8Uk84
6Vr3jY262wJAd94xZGWK0uzOZoIyzT/uSpi6V0+daCqEWMp7TtzYeIECpdlv62Ia
E8QsuxcdVH/1sfHCT6FHGQ/sjxUhMI+J4DBdbCYTwTg1IjTQeft2vRkPrXmKCnku
Dk4F5cvd5JpjMGE2xfOCcQvIakNHoJ1hG5WA95b0dWF8+/BoZC9DY/VEgme+y3Dv
qigJmQevgwQ4u050QE7Y28VxtiHHU/Mw8XpueNsm4AreAoOaAoGL/bkbDUhE8fS1
kipgx1d1feG1jDmobMFMcEI9kK+dWxYmEKQDWeT0qa+dr5RJEi047IYbQv03Yt+g
8mmblrk5U2XNGTK8t8enTqegOZvhU5Ry6ziNCNdRf/XzJNKr0zDUuYXOJY/9oMtX
X3FRp5ae+pwOEgDPEfLCQHWokzpOwG62bE+IZr7UwUMUaGU/j6z3mrF1lKDnamDZ
W99aUQLzQUgALZko8Vp3bmHaYw4VAKmWua8NuKI0qh46N3dMHaUYuFf79c/lURsE
ZpsRLkg7W9dbJ5O0gwugqu80GjpUHLvCqkAdVXX3pKsIY6Adxn5h5w6uAw+1BJP7
Vsr5BIBkBMkWbBrC2IEKCIM82JpDNPYn81myk4DVlpZFHdn5uHg/f/DaeTsrKZh2
KYWVkhOZgvqk/b3fbnXOAcRyoIqnBh8sYdZjLsWH6k1wbl38QVqKrH78uP0m+oOa
JcO47w6A4tKGtuyu0vp+k0yH0q5zWlwQl7kKo1005lYbCQbMjUZbg4UK0dPfIA2o
pon791ZOsW37rvQQVjW+4wQyUKOBHvwIYQ6DU/B5Rg+eankx19xEvIDo7283ZK4N
Bp9+q8LSBzk4vtzjlj/IUfpoqwRVVrW0f203TXad031uH/ALR4ubGI5+loklj3E8
XTw2l/kXjGYCqSbSrCV/DP/zaSxRsMbGNoh+TMQFGc/owxBCI9LoDv8dr570xT0V
o1PEOswp/a35NoE0CW2jAbR8npIdJL9UKxW1+tf72zoxqOrRMPwRfocOlTI94evc
wP/Bi1H8fOi7hBuQDNqNcOWV2P7WVXUUBhq1l6c+4DhI530ULC7a9tNFFRMKkRXq
4stBuSLf3TmHY/RaCgAuAx3CBJ56DnSGJkLYz4c/cFH4llCYKcHDAowUSBIfccKv
Jya7SnEpeoDTiJtU2fwX+iWJoFYdpZ4NHGt5HP2rligW0U5+qcKFhAc1pKsp3Xwv
7UKJD8X6i4HSUrEREfJojIwbC5upZyBNDw6EEvxpRiHj0RCHS3ODzo1clY5LMwqW
Bg0SNoRaMYKkJDLS5oRWB03lHd2xYHfnr+F10K/xwXW9hCNK1z0Qu5QzLyVnBh/A
NdAqGNDzeW1cdsZPMYKEEbGNLHq/e2Rhh4RH0IF8o4fvJXOuG1v8Sh/KIw3/UHmi
RMF0wU8nCox7/0RKE8E2wvpGkUd88Zx1oK3/AAnq/l+19M8EZuhyPZx1IaTTHWla
BwZYn6SoUG6Isr5LlMYbv6PsWJ0ffwSNeonJ6KpcF2rI+RdRf+AIZqH709K0JoYH
oQhlYBab0davRnMhUiDTyxsWxAycOXEUZ/B/nsE4xDb/Bhxbg8QlahEXELEN2BTu
FPvepVB5rHKzAdScncQecpCVOonXpWjqttAPQK1bdyVkdmnecM9W2lQuMqX+JM5A
ghVJ5UJIa6Mw7Bm3owc2L0sPy0qv2WFvt1gGfqhPjx5sqd6BlpR2c1H6OcW1Rszr
HetXXEOVdMBCduKbbdXvwk5j8A2lBA8J9TeyPH5NYDinyFlU3uYiShqsPwg2Xr1C
jLGJQ3B6B963Hj6+Iz6xXiGmjw4wYRPg6Y8XnDY969gexjNcg5VOVrxgZgI40GkC
uBfKeRtqNBT2fYPFJRB+ph+EDLz1Svf22Vj7XbUdkVTlKeFaHGhIwHDlXET2cFXR
y2wtYjj4wpY9JbSFRuzFoi6XT2oVNRhGW/Zu1eWSszVFE0pn+T/S9pGI4IrTwpM6
TzGxnXUprSkd5IQg2hXvk+epW4wE0L0Yro0lqK5X028aJxdxeZ5eDyM7a/zXKI7D
vk6N+ktqEeb49lhQ1FsTzxmxI4eduHcP7pj4MIUZQmrlw7o4QfBf9cwE0oXEzQb/
RKRcyPLTX/vHi+KzVHLngjUkCYh7saO9AIXUcVmD7M1EpzR8iCDhSTLVGjx0lqad
p8rqw4lQ1cK/PED49Qhto/Y57LzH/7mcj//VN0ynqbaC/nz9mSxK6TQr8/wq3LPB
exjgezVbbiKi4he2nd6Kt0icHrjjlcL3spLXxxMTntfqmeoSKFpEkQWNNgVOdZPn
j6fCdhOgvFq5DDkFqIOYd8FYCWpaZM8RaPSc14AAc82BABZskuJz+LqNHIUr7QIP
S7aEuGvoDaZ4RfpA8tDGV12oP3CUXnpJifDaQ18TLzzHd/TwhA8EfVXRZ6n+OAw2
3WfdWpFmHtYRWFRDQq71KvIJF3te8evRcab+Ioxq6fhgqT7t6I8sRhok31YY4eAA
NdzOFTluk6IUYeseck58/NWQLSVRteRnRQv59t0vGYh09n6/S5nEN+RO1Ye480o5
V2lIEc51sKfct6v48oAxEuPgmONB3ihKQm2bgcHW+QNYLBpuZfPVXN8mBzZI5olC
ZfGKqW9oiT9vQyZE07AP2pGggjY1IIpMDUc0x8MOWqFYbrEF4l6gbk9dFn9+1zxm
xj0i0KfqnykVJ35yYbQYUFpXs/hMEWnlH56z0c2ACq59e9st64KFxEmOlwIkKEA0
XZ983DlFrYFR9SWpJ1jIvsaoXFUVZUaNx+QE38c7ka2jL/rm9Ba2dRo4aMLkBjrM
iYPFyZ9xeuUZ4NnjzBUzyZbWPFfl4OykEcLOezJmGXrlnQ4nt4dWXrvJgyajNNDP
VRSG102bZ60gTOh78jsmLBiJjGQAFyFXEC1FK6kTzBg7t97qraTvNteSndDFfEKb
HQ0UHwB5vxexaSvNw3xuBXJ8Ya+wsoxQerbNYZwABwEV0Oc7L4zzn17mmMjHDeIn
N6VvnLqHBRTr/2ckUfkbooIbjm+1o/eDw4dLQ2VFvi7HFCTRNoTWM1WOF6aDxDLB
2sIFjPrS1ZaSe/NSdrmJcJ8QG9WQ0usao+UuvupIlYPib/xnD7KRn7lXkxCc/10r
01IzeQIr6C5nkp4EQFsc3ZPJIsEup2wi+8a7g/69IonFz+atBLqdmg9EUe5ORUCi
oQRUaLKwJtv0L92Fb3pFKXcDMmsgA8ysoxHvfhA3ln0g47osRsZ7+ZtJI1I89MZC
lCoIVm2z2fJVOfeAlEV5ly/Cby8DC0BQEUGu17Yb5wPo8M8kVVqr+Oqyrb7u2gPd
MGxsnxuSsZqLpzJBcLQx2ecjcebDqqyX+5BiH8AGsHdILPTOfxqPsv2cQw3BfBDQ
oSlIm7nQqlgEPvG0X3ZO6kZPxMeXk66MbzVKiFpFU/ehN+5nw5QOra1F2QgPITi5
q3Duxf7A+FVGY7YE2L9TeoVy1lclkiASbM8/c2yo51uGPZViRIrbmwkzoMr5aZ+t
ZvnZqNGQDe9XrsFt0fnvENpD2RLzQnuJwmBC4iFJDY3bDRg1FB4LZdTW8PDecBT3
InFb0dXFnOJgpgwu2scdfH4QeN0sRlpp+sWissR+yjSqY9YWRDgXT8gFN8fNK/Ko
VLD8GocGRkmXIrO6hapt/8xSAOew73ejgSPWe74MItYer829Lup98v+20hAvIsXo
i2bPvrr4HzIt/0n1Kum4QadrBkG5w4ElzKM9SMYl6AqIHjXbwQrhjKm7rwpuR77P
XzaPuQi/W0xw2wIkIR5feyVnqCANPBtMAblwBUvBAV3pQbbJFQ2ukMrSKMEXvFB2
TiSrfQR6Fv0/k7HxG6CNw11HgyuZ9vBivcXnPfFHTv3MR0RtKhDV18cQ9tay9AYW
ThVDWJBydevZ7/rcw4k2AJE5kpAidDEiAQY1jzF7+nxIpuhjs7OeMGhpi2zZeD5C
MP+vGG2N9dpDbhwW2B76bg7EpbbQR0jsiFncX/4QKa0xNjVa8cRLkONlrVEeHbaO
DRejhVmLNl+VGySfuyxpQp7ec48wIAcurIyanDIPMo8sgB8DTTJh5TkInhh9qhb0
qD/qj6hz6SZZkJXfuEyb0F+G8A+ktrgonFoln1wQbpqgqumPPNxVyXNpNOg2e60y
ZVBHC5jeR5YjpPbPFEU1npQoIQBXHCd5mEW7c/qBtVjkMz6EWmXtlvzlwwDArf4t
0TUx2rU26dy+9QWH32OfRNAAZBJbDvFIz449KIKTAz2SkWAJBhK7Vvjj/HCZMZWB
RAdN4qfppZIp0O9kqxkiU332QDZBB3c9Az/yBebN0aVGnFURHO92xrc7R/AXHP/Q
35y3FNixzhlhsa2een7h1AWq1152JAlxu5vYk8cfykxFmn1s9iVujDeSDIDBxiqw
fxkGApypin5X0WqgWpoVCfvJU5alizlDPhiPGKUIDcLsmD1/4cjnDD911182oHNR
ZK2LEry9QSPLrckkHk3sOMFX3v8l/Bz9unrDvuoFz5kYMCztFCZ8uASkQ1sI1Fhw
MlQqJ8LRXBQ69KBpYGiPrxHSzbrcKrFD4IsPEYWYxc98Bz/YpBv2Ywsi1KOSWi3y
czAVhKZrE4lb4fetlWYCYbqn1vlLMUsC9kML055lx6BxrcpCgXsr4H0Lj3Eigzoy
1h92bvUFkK7P399GDZZb4j+fZOtwwihZWN3vckR8gpDVkC7BbfmYi7++FTFmGTZO
SI6o56TDU/C9OHcgrJt3UV31JMP0nqb6ihSCg+TaFHf+ug/OpACDgLAfZPxRTW3b
FZNhjm0yTwbfp92MuukgnAUE5IIzgMHIz5yP/FKfrjbOHLYcQ4yILunUUO8zzICr
r1PorX2lA2zIFqf1PLRJMrIIGVOk3FoGZDaJaxaMOd5scj3n5N76V/T/rYcX1qJW
qvEj+FclORnf6OEC8j9HbhRM1+WzBMQGe2vht7zwO1WOjbRgm5U1+/G0eqfwKalC
Xa/5U1b2tZl8fOLGUmO4hxXGkVZczCon7lQcgdtyBM5+C3s9/aXh4DKhO8smeQAt
RgVNMc9uThTbplbEcdI29k3cOsKIeKpvUHmi/ZWVul1HKr00L/yRFiIaVj4qfOkq
pLQjMCy5C3n9FFifXIs3Vq/pU1bq5SXvhoKJdud3HDDsX44q4T4JM5RUKm7m5nbn
xUw8pk0iMq1Q7pGlz7oDylvINcw7hzX/b718ys7zsy8ccEkEGKhSmvtyvB7BQPJc
XtjoaPeV943KoOTMl9mFER8MU+s3jHKN8hfmwQQe+7qmFp4n0UUSlQaY2ID162Cz
HeHnb7QgbpUfC7JWAIElUpRCSjUfb2q5JgBbWsffjiQlvC838jjHRwGnxLzedZ1d
egA1nmTSNbEg1Y01vY/y02UAbYrLvHwMME7U7KU0kiLLPawsGUJmJiCGMpCoKn+Q
Dyp1gTluB28UUxjSofJekHQAxhGruOKAigox5Z+nespAMBoqHpg/U8FobD9bdlL0
X+tOEgZEyyHvQU6FjN5j6IDawvXw8+mljJknZwsKEk/5c5aW9gTfvP8Kegoh/4Gr
SaSvJNigt/W0j05ieZDLX57ilHessXqYTUU0BOSekvCbaci+bpszTvLBV11wXmg9
7AAJGjDysci8+y4d4wyZWirhEZ8FEW0B8H/qL9Gps6vTdSaMCfOgh5KB1AdNwgdQ
hE+IOUsoQ7//3F8TQU1nvhBNJMoe1Zd/mKqjd5wF35eCNk5hB6KaRoOC/iYOUDXO
Uc0R/8i6MpB93lS5MPfx82b/1gQZinqZmdyRMpSO8y6dMF+AH0n4rwQPX7cLNufC
WRDtkSGDOWm4jP9J3FVT0Dqq7UNwMT24BxjYWQRBsyxLHIAm4l64nRrNTbgHO3k8
iJj1X8yi1rwQZxMhQ7oGFusB5vxwUEaAfW75eRAqEmOfYsW2J6H3m1UlZTrH9WwE
l6Z6SxxLU0EjBliuVsBzmuVF7w+PQtX08L/8YZ0vj8GgJLj8/elF0rvA8tp6z7et
iqBtWKRblmGnbWZldwsx1MUU1TxJdAaD13HHUbWCAxR0AxpbLNgAp7+udVNxyN4s
Ev1CjKgicBNGx5HFc58GSFhCxJjuLL4NM+sTsnoyuC8Lhwj3mTViEVUaSLf+ukHL
wJUo91gY2/ldP77r7mMLfFyBXfdYqVKlz2IHqGEdP7vwWfvL59SHhs4IXUdzQYsc
aEq2wJeKkgnOGdw75U7X5Pnh6agFXqwVZVnlq1D7mdkHDjd1UQTxI9UdqnLzVvJc
4zO5vZIZhUYgbv6olmNATREcz8lMTR1IGSGSH6HlmVbpow4I6CVC9i1mVdyByAQv
Sv0emqfUv70bKUPyrIxhIAr7lclsxLDYWyUQZlhE8bqnAUGVCdX3Z5Owvb2NSQCL
V3X6FjDix12KckdpbDaOa8avbIooGvB8gvVH/rPEu41rpKD4vc5v6y2Z0LCGcV5p
8RE18sJl6G5+tenA3AspJajIw0CORLUNZ11dn01xYGlTbNHJvHi8U+LoMnthSISy
NNXwiAXq+F7dVylvnX4YLpfOu2ROUAC6nvpER06xIGKbw4AzF3vZyN98bkLFuvDa
f+VJBXvLKqv+WrA2oPgZYC7PdDKHii1ulGz1fabROBiRSpi9nORTC+Plgrk5sg5H
zB5GGC54Xgn6ld88m2yTz92Y/vp4Mr15DpLTU9RGElPm7TUulwsJylebHlqAfFOz
ykxUxZyo0AozXqg884OhoFTZUZPyBMn5EIYKbC3yuUU9XgicgcJaszTl5/zMfWlf
ZNOY0wTmfr6CtNvK9kbJeZa/MjheI8d5zSfHrKn88QUUCpFfc8CDX7OSISt9CHfA
VCpvnD5IcT/fGvguzVG5JSYT5q6g66kyZm4lI5zSjc7meFdhsHFlcRsbPWb2+NEZ
9NjuVNR+ew+LIdQl6EG+v4SOg4+rzkFrZ7RimqvdSElu+3+XnY30cgzEW0iNCOCG
SSWVS3ehS1FPM1RfM1DjmsfZMeFgrKUO6Ir8+Nw52gKSGJc/2d/+2cqkLsQUKRE0
PsU8SaWuvOMt6MspjyZFRkY95sE70tH+iwXWs4lrmiuWli0WxzN2ajVpHuAFsWZE
fE2cccLRB0pifB9xkNktgWLeKy5bz3b8XPOuT4/ULUTSH6eBeHyWFQ4Eevn/S+48
Ksyaysc96Hx7D1Styt2vOEgalVLTDSTK3iGXzJRIBKc4Y+Zr9lA0IW2rU0PsPk1i
w8tNewwtR1iLVdwksuYxI2bN95cd/QclMPRbTFhIZ+kGdMe4maWcH/7vZsxjylgI
2j356iFTKeE7daxk88PMYXOMivn+6XvNk9KxY3YJyVU9nOiylV3v8bKkECScies6
QCG+7/j7U35MKIUSpY9w18Wdd+YTJ5WN1RupBBh89CO0EKXKMN3hMiURtUckVBMH
evSQz0cT26pFtgf3+uF4QsEd2fhkU3SNCuNgzWLvR44Qxjph3ERejZzl6DGeRPXY
xaSV9hxht7qXa+PKqyumemCVk6mX45uEui1Cb2/FQFR1Lbmwvnqk3MCvF71j52gc
uK9BMA8lxowBhl49ufBmSoLKd35LATmKszexwOfOJ88gFEyzwVuEODZhcwqX+fyH
9/WiIm6rEFKlotG29ita3xHH5wlBnw+kUomEalqp83AqnSeIN/Gn2VQQJHXEeHK2
8/p3hknc4q2vwVjLuSuDzf0d8QdgMHOwLaF0J9T6Q+2sTqvlyqj5kMAL5LiWU+O+
MsWUEtc9dfu7NDyCLK6mCiktagQ5ShkozsFSdzTgBbhepb1ldCbX/aoAEmbTPh9Z
3MvlW5cUulkXwff1AM/jyvBQl+XESLhVHskgNr8xmevWZ0tbc94w2nN00EB/NDQp
82YAnXUPYoURoXflbg9U8C713nDTdr6W0b7I7MWz9pGqAiZa1dQzSDIUFsO7Oq58
ojVEkBowvLgqKuT0e7tfc2uC4Jn9pZ6mpTtNqGhgMzTCP5CyVyi7GV86nMghUESE
dy7uxg3vzTZvL8puLE1PzhiPU8pAigSIjDWVqzI5l2/rAHCehFRG1eRuiOGT0OUY
k8ZhupGFfdlsNzevYgDMlsrIhCFzFs+mOjrJAGIC83GE7i6NV+/4G5q4edNrMXx3
qNdEoy+tUDOtIA4fh+IfhKObfFuVT4HWDdHF9l9Z6y23hnooUjU6v+RRfmpQQlVr
+WY+K178d0b6YaaFMs1u820DOkaLPaf/1730N5PhqAge1GoJGkQGLDd5jR7/DQUj
cTTwTSgWfulr6DvJ5U6EGOy2KBCcshKXasinsjURPdNq+gZEtMj2AxP5DGg2xN7L
i9WZyLUXSFErUOoHnBK+AbdOjvBhiptRZxlzH2/ZCqnMW5sSDIgEfphYhlZP5aVv
Avy0q0TCPtgEEkhLOlPlUyMQlizcnAv+kYx1OTU79WI83rzE/sdeAELMr7uvNzV9
KWgKczn2kfDhqzjz5JU+FoNtrd9Q2PU8imtK1Odsycbh/tzJ8ivbqZhpZ1tKiv7l
kPTsIzWB5Ekc6LoXKk54Agy0Qdk0fGRP1rIHxGg+eSq+tenMbZ+brj2fH1SZVXvM
7ruhEOl06/JGyuswl3J0fP8vMaEd2Hd0hvWFXV3mETffEj8GsceSW2tR1KtYdr77
mDkCmT6q9VdUDHLoSpRToYeIBBAoQfOzP3BzC4ToLfpy//lKdYuXlzyPzfRyLEr4
F4ZTZ4RfjZEEUtiJBd2ysSGnz7PCdnnXVOlZojYwFMU3GmFaGpEFLDR4NJCKlRbr
5AeF/six6QEj4RQPjAfoWKSlyGDR2RH0oFfmAQKD3Qph145wfkN58K1xrBDZlY5i
bpFKiLs43IIFtFzIGaOXwNWkHfHr8oFZz6ZwnvaPVquvM4bqGOO1zexY35vfcy5R
wtfnyQ6qljnuu77XU+FgeGKD9rsHvGAPEFY74usaT7SMB3afoQ6bndZo39sOBfuL
u8k4SmWQ0XzQhb0FewaNYctXexEllkSEzVqs0nKMbCpWnD3O/eYAzyAxzFQrmCO9
XDO9dRpsYkl4g7uJtTlRJpsZ5Yuhg25ya/U6dnjIZ737MuPQgDQf4mFqfi1zRYuv
tYE7PtJhpWEyO1AfQ8TwWkc1rLcbnwN4xS9Jliv8Zdz0ZYwXeN18TmFgfVW5y+GM
x4h7zstYpRB5yVu7ZOxynfNgWkfd9pTiLjNNfLLhP8WWgNIs3JNizdLjPN7HKLHL
IFcwxrL1jy3sNTHjjYNaAggIyQ7mLA7nILJSXSMDu0kBKYJd+5/dU4Tq1SdSHxGl
8fjtQe8L1EG7AuvjhUZ5Ye1ZzX3DMQwlBtWTFJy4xwiMdq88FCTBsKAqtlcdc/zG
m8pAe12fUld/kDdt9DD4EAMI6pI3ck1Fin0v2emky4hPJx4FHLW4QdjQngKnGCqF
Rr9sfjqlxxz27MP9trX8Pj8eNRumWa/qGnnEIOgovK9EcBrOvF3v4ZRWMTFYEKn9
QLSQ6rKrb1p94Wx9XccncJvLAmZzrG5nx6jc+40coui0QuWZxUHzTUr6PA/qe8o3
D/n61EKtKMS9Jo7RcpTaP/+yqWhGztjs524bLd8eJxx1Vo5EZ7DrQxwwPXLS0xx3
tYbvbtsQFaFjx8RdSG0x65lwJkSfuouvLEIuXAY7c5trJbbRbCKAPGGUcdaUoJvy
4hHExxmy9dQmf1n3vNuJqKukn2roinjUSIobFnALJCPkpkmWMwnl5btwCpUo+ql7
9ljw9B+RgV0MVzix16pf1yCrz30bHg3B+RzQNY+Oi0MOpQHUVE3fLZCHc77Oojg+
UKvEAY4REXuloElLnpH1SZSjsyGkZYzD6MFvsYLWwYXUAwjYvub90jQ3oIyh1N84
+72afsfqg7e7yx8otA2oMpnGz+5NvH/XhTMzgOCQdiC7hHBn8oRdM/6Getu4Ir/O
ddOrSY4inci+a3AfMIGPFOFo2Q4dA00JmrvW5p9ORL47qUXsFK/fPdXVsXJZ+Oqj
OvA0znfpr3s+tkpBfiyOgj/UtJRcgZ/sh2Y1NIQ6AjJ4sceHy+RfQOWTrgWPFxb2
62vA5Ie5aWRFt8JtKFfusUDukHnurt+29SgTNj2ssJyBnPxA8mWLCyJgWE94aAM0
pXHN3NX7VTGKoo6tPek2hHEgOA73t8LZNrVtYs0J5oPqDqG7QnLrZegt8XzaPpgE
5uRazY4gwnA4Jl34CFyZpnGuYwv3jDsXkNpOHsV2+TDJYqRObDkL4OtCmOxCB9lA
skTc5+2nYF5DGC9XMUz1BAoGVggM115i6OunC8RrMfYkDOQ/s823dHxtrImqyVNG
6rFFvaUNABA91mxXLaTdw/FDtciRxtz+8eU7RfS53ZHfOvFXRxovWuE0HKIqhwr7
i+ZgMmQ6AB6W+h/Uu92B66VCql+Sh6OV7BdU9oKuhTgjTr1S5Bl84tlKUCqZiok4
4JOScLxdFc48n7sQT2373NtoqKIaC39Nx74cHrpp9+Jsxey6JN+7xk1OdIXZ1N1q
NQ+O04JcVGj5OXtcgb3FfmK0l6Ms6ZfKmhxxS2nyakdMh6eNJLpcCIe9oMrvrjz6
ZoPAI2P846BA6m5A6oetlpUfUADxc95fqejdmdpST1AiKdt07oMvp66KY/CFc3IY
Q9sWXkYM6XFrkxYHJjm6TEcR/BvVqqMbxkFAa7z/c/CUahYWywUldQ63niKeOgb1
kuN2lG6h6jkGSNdytLJ/DfaKVZI+RXxT9wAwOAEzTrSEC0Q+oc7JuvnKHKYNWpx5
6Q08RmveV5TEj29seaRt/DYqjweMmsxGFSr05w00Tfm48A+8v9NU+7oMnPcluHmb
hJkWlRtP+fW5WJ/FvRwxv+b4Y0ckeskmExh/0PdCksOEaSj9u9oPEO/RPqRXV46N
NL8zH9a+YC0qWXuH9U8PKtmPnfpG0qxcYNZWgbbqgQymHQsSTPGDajoUYrYjgD8s
K4dNF+yMmm9ZuPjH+LnWoDETGk7NELdWI3JFQmGZ42GlA6BI/qyrM2n7CtxFBDor
tplapxoj9FmipIcBJ6YC32gLxn5dwebdWEcYSnRN4xRGJ+24OQk6b9+EDjZcO6Q2
8P3u1lW+TbDZSytmaaBBwcyQAwGdIzYxtnZwT3o+vSEZL4Ft6U4Gav4FyBjMzhNe
sYnNSJu1DLRl6XQgAceVWxyNrDUMdRtVUiCyLDNqt8zZ+iLd6BI/F30PamdDBLWI
eiQwRN7uh5ALokLbi6qkQsYp/NBKfNhNryOF5CIOG6ZbJByPWx1Pk/LSHIsPzO1h
TJGX7D5ay6o5443qFccVWojVJQkgT4/YZUjtu7CVD2HnvjxFiUZ0di+dLR6KrERv
ioeqV8Iq+SUWYAWn6gmQpbMe61V3OF37+KbELV3aHNLUeHDZVwWD4XsdO5xTPAEn
1gkqwYFaLT8rXozK0M9gV2HbZUJgORcEymczQLzYCCztI0H/YD16tJgxHuCnIddO
LkroDdNYv4DKbr/sT5ULWVMNx0fybuJSOK28CpIY1yU0neLtcJspKe+MJbhffyuK
wkEojqK8SIyb+xu1frYBssBoxwoMdTZWYvAu5zRz0NsWYBKw2GOHDcTdXA8R2R4W
8pJ18k7Bf2LX6kMbyYj43ExOyVuCsiIGT5HcgFHfpqMBRb6uwiFhGi9vPUDrhgi/
JA3mZoMlTD0bi5amfOC/wazQMV/MaY0/LhVxCQRkz7Vb0hLG4bh9N/YL4BTn8qKB
00BNy4TGueIyaNULR/RauEosj3SbhA+IwsMqQfwtaGGAHHy9kwKXY964ued8KvXC
4RigJymMaISGQTcwK3JyY2GKV3wqMXBljK2F1UqiF9tmYL0gJZLmURfouc3lTrOT
vC42xgjgpuiU4BhzS2PRQmdHYZTh0feftm21+p+g/mgWnlAPvRtag41Oh2YIyjU9
hXDyu/EW0xim8rv26AZXwJ8/FKmaJiRBEUh9Ehik0HCWvw/bLciRn1ghm1rtIXeK
lCS/gEkOBmgQv3F2C1gtu/uLqfHBQqbq4sXUcaZQ4xnNmhmLRYQirQRjT4udyNJj
N+oDkZHPWfZ4rqmt8Ws5u09PhQHbWNeObwKfQhaIsWTL0qkJfDi0vLlbuVq2WCnX
MfmglSda8Knt9Sr5iZ9JOv4Xchcga1W4XoLAzc5lGk/JMa84+Ti5Sv7Tx0VtMOPI
+H4HLDVDi3ZWjiLzsOldorQhgj56D4XmXaHNnl+Tou+6p5kYseB8O7mZpUvhvdsi
3tMOjt8qgJB4Ql+XC7NZQtp70OZTxb11YjrpXMkCAXZponnBAZHy6EGTZpmzDsMu
wnJR4OCI5uAOHRPACoJHoTKWGLqNAhFXh2EUPQCmzdoX+iwwVdZZVUu2kg9oDbY4
jOdWLRCAG5ob6gnNISokQ22O0FeIVKJshNBNIpZ/6gJ1BYyOApOOUED6kRVQUdxO
47qgC9VDKF48+TRDfgeGz4aXIzom9royEBpY+xo2m1ZliNOgxc7tOL/sdTWw1kMD
K8n5VkWiro6I/k6jkLD1wLpW2UeNnJ/AKWz3JvRsD0algCRHyiK02b+9U0fOKyCC
BmYMH0gHtYNUoR/asQ0JwOYivrIv2E7xu2xfXE2MpZO7Wgc+674CrudzTepoPbDn
JfuL6sZYYZ/R30r6VxLXRwMNqjT5YWgw+QYkeXJvyg9nymiHgbtqrvWAhV6kk0Po
qagd7wMo+meH3DT/9PVKbQ0Lpp+w9jennLzHHJged6L9obN+mdo0f8uBqy2vrAsD
F/TOWSJUW8zhA5+LXGYT4zU2t2ofW9jwZmapGnc8Tjvd4yLBFCmciDBw4zXgmm2j
kMxkfKGGrvkI2L4towuJJd5HPej+jryYJDB7OBnwGRDpNzTWVhr+NkftREo3jAVf
4WzpMr7jH9TmNYCWoabNW8OS+UHPIj6vGmtkqKytVQrSwvAUPPCiESwni4mSfrym
nLwxVZG2XgFdrj8lwQWZieIIw/SXWjVV0RZsdQIcoH3nxlg+TdlhK0KQUX1QvffA
gz4vtJETIBt4qRzJZkUGVnSehhdKZkuJ0ynpyjX/HxV9bjZFjeqP7YHYReD3GsLK
AMewwYEp0jo75uL6v984d2g//CjetaKe10ED1lEQX4vnhrvApgxVmWFotCqXFUXo
3sm7sAwEQ5eJd67iec6JkuIhKq3A6yfLL9baR/SiW+rNiOVxgw6GSKvxKUBE9Nq4
GrIHONTLTBq7VeQR8s4PbwtVpFZoOoVODKjoAfBbv6Re5ZLy8PX8x163fQNgn85G
JH5udergyI+4Ko8NplP/uqkO0VKNReM901cS+UGZZcXCZ0tcx91Uu4hGV+uG2x30
MMmDgMdHbb9r/j9B+7JuRBrIFunkyM3u75OLg59/6E3pA3b39ErFLMtSR/5GA1G7
Rcf5glwq2dNP055ojZMPgN5P1SOgeDmRlENtmdLAHcsyQaNwowcDB80dVlp8Hd24
euOETB9DS26u/NR9e02PEXG9wguR6iSeoV5D2mPnID0wkd0T5+HZc/I4GFNCaMwZ
I3mNgTbEIhcEvWLFgerVaiGrwty06R1Ts+diJPCtFwpBxkwcuLh+kDEnOetf4Wlt
rXUD+/PgSIH4BoLfAkTJI4kWUtzzDUkic5f8a15Nq43VOyZbzZwqkZUDjKjS7OBV
HTIsES1LOoFUV0YsX42QUt4Xk5ULJqUq8uTOcKYsbHBnJKd2bCSSilWvZ6godJAp
FPGMLyGA0PGPKjpXahgQSnh1Y3x9F37i6otP0tYd8zYulHa5Lsb6eNFUe/068Znx
noJXdN9YRthVxJ18NF4WGIlBA1DvcbUEQFYFR74gwyfJTFBlv/8SKPuR0f38G3aC
3xyrSIoOylQRQ9SzVtqPPcMT11rLaAiPLBrxhkiZKVTNhb6KiV9SbTyI3Cvr87J4
elpLZbcEpZejvbTOn3v6Ja0l1IeUxxmG9/mZORY/82IIW0OmuaoSZ/QjJv/4K7Qr
Otkg9Ys8nuSEX4OWDil+Y8o2zCEqBQDIEc5N5WHWq09v4WePMX3IpLaJ9Z+qijLw
+ruTwJzPlVS4oWEqh3yPETVOIuJbwI4WQFdYrNoY//uDMd1xxSErGsvgy5M+rNVg
RdTimTGvD7JkM7Zdr7N6JKqWV+jyQSk6HuJifUc/2354Rq+BKFR1KqH/+8cCIG1B
irbjJrg9O5NFTL20MIWv+f06mGUniXfcsRMEzmOvqDu+o3DO9dNJl007+JY/6JQa
A32OMl25WwsogYFSrTjQw9Mdl578EmuTAXLfxESQyLirYop9otiYqf+qgZiGDocQ
l12DBdEjnUmWzSdyS07irsRDZds8y3UJT6TNNEUT18S+ZmAW6uYK6fRYaHRXmGnO
m5r9jioI25XuU/m3ufieUzD930LyRghL0uZCWCMQ2ZCe9D9nwD/as/dLayQNEBHP
QW8TN9wZZkNzA6/H9h6KHZzh6bsr36Nk2A3P/EDMH3p8W/3eT4CIXLfJnx/XqEn8
P6ZiofI5KysjumNuUrJ9fpChv0QfFr5kQOBazPQxvTZcjEKqClMfNEcU75YXfe+6
WEi/yxgx9ad6IK+mfilNEp4tJgkHc0F6Uqu7oVhVxGepRoKuRelJyy/mKhs6a73p
re3ptGEPYdwWP+lycUK4/1HL0Ois9+ZuQvH2VWJLvDY+ddv64Ms/j3+Kw7qpiRP9
855u1MXpbGG+RqBmZFHR1xZD0TGUHbHpuV91brDcCzFiex6cTj3s0pR5Vrqncacx
d16NOxyTMYmHIrkmdZELirTD+1iWp8wZS+kdHqdiuxQhJpBY/EktwMxZ2c71qixx
SvTY6njnmFuv0HIFSrLoB1ZCAMBL0uoUwXMYkU6otNoLl0Am74xHhRx9NJmCmc0d
LOOqK6QaMLzQwTwX/iNPlx+zc9KmSIUJYdGKlqxKefmzIlHTVLZJkB7LiBxrQnoS
UIl+iLOKPM7okcUrY8rP7R6jo4nOEt+7BydsqDfhnIGd6Xfl6t0wOnZEL54qMvwR
UAnGQpXRq0occkR6lq8gZFEJb8cUcktXe3uG/hsJnW8moEckvU87KWPM/GDYOUeQ
NqYRfqsnRH/rHkvT/y9UCjQGtCXvevfNsrsfvUQSYD/5S0iS/DsidpIXZJ5TDyDL
6wS25zHKWvMm9QNBHyCajyxFooQs8hUkA0ru8xmJruEhGnY+Rca3cXd5VzLeq/88
OrTkC+8jUmWjTc48Vac1gjT39v9+VdcUVr6ByHwaMfhfF6JAEyngp2S9hLlCHNKd
Z52TWv/wocx7k9CdfhRfLB5yDY2B7Lw2ys6vLHjwDajZUvD6pW0/3ahT/1H3HLCj
2RUbjo6Q6Jw7/eaqQFB0SjJUZqO5aLb6UkLol9Ki/6JAWqWq8Uxw+W8J/o/kGCDz
zCiX0jIy1Qs1HygE2t2EMiU52IdXGT6ZebN+25Y3VeRaQSYWF3JO5AU4pcgCJAnR
kfMbUvNp7OZ6TY0lgfRvLF3BzjnmFoA07rsY3q+0G7E+IExU6MoZ4yar9VQgHJZM
Lgv2mp0Ix9Dtj7eurVHqwRwdyrDlSMa41+0fw2ZXi9tPmozpJUOpNr0rhD2WeoSX
Zx6x0mSpreldkqkAntE+xKLz7KyMN6hYj+MvvQAZE3LFRQrwNPTrN1Mrf8pEsnZt
PE9A5YkFQO2hLmjqmGi3/7wjG833T2XugKWBMUlC8vRIIES8oDS1RXonSNBVWNnp
ADyyyIfLvJj+P8DWSU6EuFFYF5w0TMFv1EEreALqrDkwAM4hhJfQgRxKHsGiwRri
oiCFAAzCWsRwPMPcC5iSKvJY9WUZTGROLbgO/kTbduBqRhFIPx+wG86p4aeAid9Q
q3FJOdjKPuMH1kMLfmkQVW9AGlQoQxxATc4AXjOl5j8BhRZMO3z9LF61+YZZq5Fh
RQKI786iblMMaek3aPw+h6llCLFyJULFAgg+eSA/W7dj7/7jEhFtwFMG7fhCCk38
c4h79yjtGLPi3RSZJLrdBoSc1WcLSgNbKJNIbbEhtmPBTreoLmIXxxVCVW4CWSTM
NnBqJiSsjf6Kk4+t8dXArmhNnI1IYeIK97x8M5BRtusobU+ntTwfkBzBnHd+q6pz
x5s56rpUED74Sp0DXvxkBqB36rSb1jQrXG5MsCKF46rA8EVlHGPodFpMOcJBCia3
0zdd115pu4I72LrBBwEle8xsr1PaLFyrvnk+gcrYDQXhh7i7gmUqoYGheukFEa3k
fOcoQ5K4IYTDvv9NcmZyz3WvywgZKuhfTXtEJqUDi/0/NHcv6FqxVKtG+skz1F/A
hJe05ZBmWk8xbT9NkjMVH1TX92BQZ1yzaR5GcT46ToqE9dwRFSTxhw4DQv6ARfgB
4n+ZWFF82w9HzJ+C3ROAur8zi0DeyyWd9q8YQu4g+LJmB+LnOyFaFz0xnd4XPwhH
7dSuI/YnBQkx7t1Feh0Xr2FEdYEtqwaB6Y4B5qT6LKyYXpbCp8oiwhrsfSGxVVS8
dxZR37yCYt06N2Rz74Cw+DenX4Puu1iezdhduquzrUOSPL3aMhoxxK5MGmEXke6q
c7WXuJSJ/bADaeouCac5ekPFA8emzuw8oUR+leglF85DS89s6xLe1w/G0Ou5iVu7
NVb6nJZOnmmSLTlztef33fv2z2cEjYCXl4hBegw3DJdYMajXELjZbO9HLAgvPvrx
oUNGt8BK5iT13Bk9O09HLHxHju3jSzGIZf/bLPzaW3G01n/4HAzAcDnVfJ+5kv+H
YKuij8TWSGnHzIdZ9pxVOvI72BKHKmY6+EegOClo9InRidhQFjlzka7Y4eNo50n+
nc3oO2GkuQhPcjN0ZCOzwu0+3k11lp2xi5zv6APaOhEIjPj0YWf8fxlMjkJMLXdX
1iykeixW3wGiSGFacPf5h0bIY17wCZmM//LRkUnC8goVhMeWsrAeX9Sw/gSjGeM7
r7jh6pcdvKNZUqCv8CmhZoDurtYxGF21eecqEhidCU3IJaSfi/if+CzMpzPfIbti
JAjMFTYGNmJk6s6nHgglTpaNBTEq6mUMSTsYLgCHOD/eQxWpXnpW/Jy4pFmVHWlj
jwbXO26zWPfyPMB6zjNOZEEX15auP9e4Fuak7Ca8q5gRcbEz6YfbwyDynYPJ/umg
zw1dVZ8kqPPCbPzKTwhSn8GTb7oaeGtY0MohkOoaCbS4MTd0mPUPvL+JkHmebU6h
AY3KKsaIdZzTbns04CletmBp9bTPaBzA3srJf7H/lWEuIwSRJFOoJYX6llrX5NLc
dh56HslnPCKMMmhYiHmqfr+qb97V1bRw26oznljsnfWCanIYYj/LAJoFMnIUw22p
xeqoXhYjU3KZVUrUQAyE30gXPZoX7OKm3BPVXJE6xMzTtTlZEawFeodKNb46XhW5
NJIsKkF4SRV3sGUcZJYwbsD6Qu5fYRZrsIj8RvYbMnES8/wtGwHgX17KK2cw6eDO
CNGkVlvWTim3PNEDACsDczuJRgrNHbZFdF8879/M5J3IcbfICE8fqrLe7IKU7M1t
rMLRvSW/WYqP0Hi6NpbD0wCxagtOPqTN+zQcfFzvbTwznFgX0whOnI98wDaTAJm5
DSGX3YiQguWTxHaoHj1osjDULbs1mtxgSUzYanO0y8UJNd6sfFc5kTGfLi+xLbXK
xfS95hc0FK8bHyBuPyt1Qh8VzwbSdlpa4n5XUT9tKXwhcqR3ooJw+ZjS5eKIIjVh
Ho16AJ2RpP5HosvWCZGY7zHeV9xxr5rRqCgJSldlPPYXmfYU+tljpkI7SUNUbpgd
ucKmXCG+sQ9twIxoawdcC7hdCHJJTNrDZRvlbWJpOS44+QJgsPyqXYEbKG3qx7QQ
BLQVRzzo5ga2AChsKwcbVqUQFcufvPe+yAkIEDI0fnMrMpRO7APkfFb98kgbDhWk
BBURO0Ik5AIwdhi1K2tTP8saf9s9fOa3djpT+DU72AFeCZBg1LF8b5ocYY+OYRdp
ES8MZDx8PopVLe+GZPZzqxEuzyXTAByOnRimQA0vtSS3wIcRIaNamql3fZN1zvn3
GIkYkSV3n6x/oD7YnSPyrfCudpo9hDoy8UZZ0ryZeX6nRCdA92zAw3ODJp+0gFZj
5oWkvbHNGRx0iZ54xmlAuMuLJNrJjVz39SdPY61xdd38aNW8aMz1AUgPxHGKkOPh
a0YGK0ODPnHMrxsz8txwclgn1f39qY5dl6ml1kptBVjTgVpuX9Wz39YlwVZE6Qrf
9dHc4xQY+F9teraDo7V4GFQOK0CzZDnZYkKF6UVIdLCvq0nSVpEsTjahIna4wPo2
rr6tstE5YZCFTDi8tk63IxtDDTkc97QAqzuIK1SgcPTq4wNedTNQp/RYtyxnlfKS
Y5ZPA6QuyT9UJlwKG1X4RVRwhUvzvwjfLBOREA7TE2v5t+2hWzMARPjKbUlz9gE7
VY33/akejgoRO1yi3tFmv5Tg8zVAOXmgpvxEtOIp7UvQ/dUxrE92jPHt9r/pA2PC
DdVHCeq/F+/M8/H6dR0ayNaF/f97atfwrFJGViqPMwtnZTcXTDeig4MyFCU2J2Xa
PqNsGL9NPFn9xZ+BhxaahlNCgEEkdLtexVSzjDnc4UtHmBKiyWKJABpXFvunlMX1
NAGiNjQOkx5SZDGUqEOEuB3PIZMS7tUKYL1/+e1QDlaa7bleEorYAjluBPRiuToz
I3OQCUgY6PrzS6hIx4lERuIXZb1gi5zTYoD/46Yl7UcXS3+DwZ/CK9MksoaskWOh
DMtwYxZuuJHB3sppVPMOCcmI4N24nl0lv9sE9zdiEq7Uzs31m/IGVL8IrLMuyIsW
Ihqh5brF7GftMgKFuKT/JOWsfWV1mU/c/gDkm2VkZuSgniVVBVP/WV2M+irqAdM1
cAPi+aviDcExhCOfzEDlcax9p5otcuUJvd2DwFiuE/uuM6DdpoGUJIbbfLwWA5k4
yRH+4S8FAP6VkQUUcJWsSDsIXSRp+teeyykpbPws9LEAg76u30JJtVi5FA2DThFB
KASF4UVC1M1sKn78GjaNVM0cIHOG+h7o0bo82THLd3HgPrWKEbbM8qrVmrqz+rnu
u3d6kzN6LmgAJno7MoVbzb9EhZp2spZ8rkmWHYsTOQ8wD7ddPkJNg38yv14e4AHo
NJaGtqXF5xvI7+lw9yzA9gi5YhmqEmRX40ijfKr+yFBzzmSwL1rLOrZzf+b3bvdp
0pHSRtdlv+ds//ZppwT1IOMIWGqVS7WXZ+zSWlqymDUkwkE3mOa5DDwaxt24XhzN
ssqAUT0i/t/2WuiYXOlyHzish7CGfZVy9prKaOG9C/ItnbZzQNeiTc93F7LLcBSt
sIuU5VTEoXXCzc8ePxfsWWevkXpT2tHBSgMzKIUMswAKhtXx6/AswRZwRjYV7PVs
UXCBZGCr+MPGcEU5oi1m45vf85wMLBe9hHS7q5W20xqbHsJrIm2LR5EtAHMbOxPn
2xxydlveRVBbMXXXikl407/CFwCy2ViMMGsQWOxJYIi9tAkjaVTfXSKWyEnhK8sT
NW+OOF5OMTVdhRfHN1VD8L+MgDFzr7lD2xCCFf4mRfo1H6XSES5tU3rMVAQpUNIr
Gr0O8OciBaxugIwFTUuvqJz8delnqGgIK1havYPL8DdAFi8orZo+8hqhvawhL+p0
mgeY6W9AinmP/ZL2Ze1HH5pl+ffnKaj2gAmgEPjDLyU6PB1vx5PVFSkb56jhpjLg
ZLIVUTcqdzpvn9WK65Vit10USaZmuE/YDRiMlrPXg0lEPOOdMAI88iasfpysAkDb
/JiL8n0yncipCSI7TmjYkmBftBEp/009CYjn5Mu8w0u0tvHIo97SMHZ1oPQTK2tB
7UurkmKs2yQ6TWMzQdgGkJoyNHIu4wVB8z8cv4AhqWDzlaHUC3KiOjhRAXYKdIpi
RpVpKodk3wE2R54/IBeNQoMXvhfj90xMZGL8GkaK9WIYAoyFOn7RwAKs/l4E8ky1
xLJRQtzz+s4XmFdyvbV1BYL84uNaFwNRmbu3G69Dv2IsEIiFVGtmKt0ou1rfy/gI
t8M8yqV5X6PJcTcI7G5slg1q7ObBbNogtMUwMo/qIXKOcJZkSsWxWE0lPDTjxc6Z
ue2JeIoOP9zg3asgu6k3Iz41qiGdZ3DJZ4ApyVCgCmbM7BjWKlG4N2tmMCTwANrf
3Yg6hzSj8Bqta+sqjuWxKbw2/ITqCgZHbIe3I8ObILAkxClCZxl+r35fUe0FKh6i
ETHyGkMht6cMCb87WVFEPF7Js94t4NLLvlzUofV/5FakJzdWSQfeY19c1qL57ZAy
QzEjw4KgebXY8gVTMRehBRURCHYc8loKGCNUkWjM40vU4yEsVV8p4IfvcI7FMhfe
DbzPG50LXahpgyUAmjwYEsQrs/dwSW9PJ/QmtQl/M0maTzYLZ9I+kjDXt4YCQTwX
K3wxE7KrZCq8eUovdmd+XYFrgI3wzCJXtGy4jjdB8E/iX96wjkuhxk7wSkuv6Yp6
joSv1WVNk08ZSE07skc29kj8HvwMZF2XO/Q/Kda8dDeN3vuXlZve/PRl+QmNUkdg
QB7RJj3lGoKwU3nXqvrysG2Kr5LcXXw3vWUda/XrlRDZ+zBDnQKwtIZnEzKcXYgN
ks8hMnaZenkQGHSQY7d3Hxb387rQHwHjGRlCHaegl+6AXJH2rMhySeuS3WyjTIrU
o9qJy/qWPUl6wEXFK1YbEeqs6Ubt+O4C36LoGNb+lMjxNWW+A6G0S8HQtFxH43ct
prijfwQJbFH184QhPcRsYKQAPS4yP3izGDbY3uSmkInpkoytrjovZEM8amePoU39
t4cKBvcpIOQnjqcaSgAR85MT4GiVMtL8aMvmpgTKPL52Mh2tSmEkkOVJGUNVxRjM
hyV2p2TDOSMfMG4DEKDqoM7HXvCN0E5a3L7kPa7lwKTFpLYAdZuHtlf3RZ009gUC
VvYXLHLgkHGEhuY09jhuTzSdBhSkp3Ta1m6mljUONmv5bk0TtrNl+YIcpnAUadYc
pzHlbSB/RZYaoANY+PDZH0PEDp99VpwvGrThFWeNeHFHZZ2cRxZ4U3ig17ZE73X+
f4pnV+sl9N1kvunW02O5VvcRvBoAeqTwVHaWehATKAj3ql41ABtFT2R/nIIK6eJW
swLu+EOEGIBAina5RZLQ/+5mbYC29WWrqqEjK5/0nUKPaP2ucgv4q2TYWc6or6py
HSa/zzqcBB5Mpp8oAAUXV1Z4rnUyd6Jm0/75rWo0B5UBg5AKZhd2/yTs3IbOnBVX
ZQXUfosvIbzHEen4tWzNWNhMVkdSGKa6tDX3woTXh6t/tz3aW13PoWcjatDmIwaP
2tyMtFfgjlBfX7QxhcLyrH/Ma08WZOPXAQd5tuy7vci1WKD/41SCNOKoUmpyAO/N
1YmYuyDuScIcf1SCm5Xz9+bHt4MsZfP5fzQfsf4ubRK14IA7WivJmGFbaHoYO0oV
Xlqy5Oq8VsglMAPCthG4ZLlYMaEWGNfMHZdjxMlSVENvwrZ5/517I4DrUGKG0GMG
PIiT7LRCdivVXi+a4B1xBXyvUyjgiWva1OlMev5rcFK9lX7T1JaTzU3nmycYXrGh
CQzc9nxKraj32z1v0h9WjFryeuSgKim440XNN8fzLjQ/iWGB6NkaxdGr/z4Wvuv4
j395/iiD0cfdziUTtEw8ECG6ZCfdJdJR++1ldJkmJ3sQi1HLawKltSQIKwwYHHL2
GUHIzzV7+L2dkhMHXbm9fuwGLjHL+TThBNeFinaSE95awOOB8jDmearlhRjkH9Vt
vGMhrNPhrt4f+vZBeKda60jthXvWsuvKpaSkfk1LHR7pX9VYR1j96+9ArOPtBGQ1
wHS7oAIEY4NxhKL2KBYEfDucnaDtbw/ns+zdulXwxBjHZQ16O8MyhiJxTkevMTBh
M3nKFJbNhX6Q6lg+Z8QHK3mLWLx4CS5CL5yJonCFWL8VulrzMpERljNbXj2S2mRW
MBJVhSTk6Rf30JwAgzSVIuWB0iDfKdBuBCuuqZE11IVPqLkAOvJkS6MaOC2wQE8w
bf6nL2WIeulAK1Q6rsLOl9EAYnxXm4mV1KOHMocK/4e1mmg4N8i/QeY/16X7Svm0
vN7+wvwUEB1zpWjdh0fpkQrdZQ9CAo9pexSsisMqieu707P9rGaNUuO3EDtrps2i
NrT5hvID69A/VXqY1QjV1ekXBHUqvoCgcGLyLRzuvxreNlYbD+Q5ve0lXpN6aVOl
tx7deWUfLEa4A1DU8wPgbwUNTlKno4F2MMzOO08XIWwZH1XtnXjMY8s1+h8wqXcV
GkBYPqZUcsQ+mNFf2IXgNmnUgZ2UkN4zkVuJrmlxauhD01bnbGSsxZWAkZnat3kI
Kba4NWJ4cmMZ/lbW45fGGOTHEKQRlLNxi9HB2wgYeyiBJ/CwHuWhZkNsOptv8Mvi
bA7P5bkB56g12XI+x9sad5A15FVAe5xHRg33Ec3vDBMre42Rv496MZjZ6Blhtal1
8r1NV4wWONxjH+pZb/CH+6Pd8oeE7ICPsV5kLq1zkCf5F7piNbUeKFinHZQ+3tUi
FYsW5BI3nKQ1UI2yujMSvvk5w9UOvXtKhYjLdLat8jA2Gi285dGEr+vM/zjiEDWy
CIvjxdGNQb7x21v56z/vl2LrfPs51+XZY19HnEFnJkXm6WktODyFpm4lYHVDd3PV
jOYJJanmKxOGQM6O/yuMgDNKtGPB1xNRa6TCaGuaDF0oc06e0NBcQKWvlhq2XLmH
ht4RGecDE1xR58clIYf7Emz+++7M47gneL67crISLXiLrP4KdvS8FxM8DXt0bas/
FBUvWH5ftI6S30uQPO8lpxumDS/9iQ82HHx6lkjeLhbVa/qYJcBzmMoLEmErm5js
ci7HB+EBpc3Ki1g55VJK5ZxTgE2LkgSx+iNc/3dAhwE9Dpp4WvCvhV20/SWrEeZR
AwRY0LI2SCVAFAGm8z6UTePWJCefxBnmwlXJ7TNBfMwOMgD8TfG3AhzNOjrBNb5q
L3BDPiTMNS72KhIUXookdF8UC+0cj8hKyZPSkbC0hlHxH8LcpGDbtY8I862+DyOK
CNj70nutxgib+dQXiUWSk7sQ3EhevldH4NEaqHgCOjyiUjL1MzK2x4OuOGyN16x3
RsnF27FXTsmZWFy1an2BleLIixCtyMNLTN2Nrx4+C7P1La5bllfzp8wJSopOH6t1
NXTwy7xxM8ZcHIZTBhH9U+8v/xLc6Cc9LUYAK3nvYQJq291OkfA6lhO1C4t1TTcD
+mSbJQo8/7PkCV8lq1gZH7LAjnmEzM9okChwb/yvLXr3kzYE9JBD+qd2lTFAo8TY
xP9CIgTEmbxC35P0P94B4/lHZ3eMfO8g36Qgj4TutLi0uwdjJJC1VVy/oFWMY7R+
3GsJ2fykarYkIaS45wKF0x8JKrMLIZGJtWRzcX4sYJILi1s/XlNOCZH4oH22bMAt
KkSCH8OEE2YNEzc+Axf4NaN0pAEGuv2HXZHTRHie8OQfUW6obaP9zJZKzR0ngQv1
3/wA7rZ2Ng0Jkhe2P6jg19BiNKWdz0a9V/NlOJu0wB8lXO0UZCdk+29PzR3KS/B9
bWfUvQWKLL1cpMfAyM5PFf5bmny+Ob3h04Q3ISltmLmuOyZ7iWG9X9FWCgFLR/+t
Gf/czG00Z4zqRhqeKqcb9JoYwaL4XK6OPYM8J+0U1TY1zWyMLWgwtoc01mkqqaa3
gAVJKVXShz8rySF0zgZ6lrtvTfwSj70ORCwVRnx6rlQ24l16FYktW/YcwyTm+kaW
fqjInk63oxJiu0AYUDGtqjB1hSv5BC9MVmBa9wJp4UUdGaQ3XjAO/atwYP3sLyEz
ArEXOnqabRCSLjBHViDyGgGFWldlJyV5Z2xhzRcm/Wmy54lMREydCfwS6QlMa2tC
nGfUX0UfKlC3+h0Ulba2pR7tZdG3G1Q+VNV6/8vOLKCWf4ZhJ2uQvyUtPu9p2Q6Y
Lun2NXhu1Wthx1U7Y5tn8k2kEGqzp7QdrDtBCNy+zP7sT6Q7x8hy4NzTT4ycDsMF
2fe4z059hNO0WjoZ9vqqoQ2gGpP8F6dpgBfHfhPIlZSEjRcwjWdBuFGoOo+ysYiF
Dof7sah1Jn/uQeCn0ZUtntpI2ZYzL7x4hne/gPjDWeESUjVDg7WnfKJC3INZf550
fmuja8r/x6tslqxx8V0DYxrkZUvvo1XsA5nJ350Dg1CLu3NOMdU04dBGs9QffviC
H/Rrc2Kc1BuCHgVCRLcEwPUKQ7twKwxcFeGq0ehRD0abz5loXKgna+o4swUzeLyq
mmN+PsrMR2KOMJTJWdK7dXMmZr6/LD81rmTuR9VeHdz4ngV/NesFKVHllKpWI8VS
Ojbn+ZFZrOmM3hbXkP6Iy0wnGhqjx1ZGN78SHWg3ve4owe5lXfSJLQSwI97+rYqC
09Jp3o9YTM/STw8PU7O1y8kUkxcVUELhBVbDAbxYoGsM88vrx/MFwKEQtJiu8Ltw
PCD7YTdtczAEUj+5jLtikL3IN1EcZnlY98twTp5Tkz5DSVbKt6E3bsJnZUo3rIee
H5Bj9Ck1L6vNPBaHsDsQlk/T5Kcc8MRDaFYqIq74sU5+uRC5U6YB8fJVYnKdWnNk
NOND4jV5aORD0CPF2svEkkH40F1sbAWULAVg/5p92GCAt//TnP/Zq1uvnChDdRcY
MM0nyIakOnEMXy12GEJWY7tLC7oBTWhZkk8ahixLSESbbSpggwYD6DkKXVpzeuyN
keRgvQ55jBVaku5PN7q9mZCxk25K2bBAkJrEKoKoXPAf62mI3qSRIm72eso6AjCv
+JX/QGqfYKdbmxMzlSW4+tGAJC6NYy5pd1boTVz7fwgLipTPpPafT3efWGHHR8oD
mUfLe4RVljgM85v8PiBxBc1FEWWSb0ZhAxcH0VIzwwfkwosQZxWxS46MzwW0q66P
H/U754hcvX7zkWcvP2nN8YJrzO8mjF/vfybCMxWSnzAgrrCsqv/RH0lZnsTFqmXC
d8kuJonzO+swj79nE0s1qnHMKkuOVv3VwC3BGZj2Pv/NqjKsl11CRoERNPo9Kq0o
iOzT0nFw/5CQSxVHv7cOZVvb2KZ7EkAkWxSLMiUnxlTy1lNwKrxB5atBmio8Q1IZ
ZNVaC0DSF6YRx9k6c0yEbsMC+smzVSqrQ/GhsqW1WB04uq7x7ByVacmXuT36U1+u
mFhoHopq63VVFTyTrrt4RzXmUYSUlauKKlzdUp62dhMzkrby3lpJRSBEuyT06ZsA
N9zKgLoL1V+DPLvqJ50OvnRwWV7i3GMiQG9NohmHBcFdNwE8srbKLxIYVvkFSnFY
+tonM5NOL9pa+cntO18iPt9DrzjdNslWBDbJVeOsJlykcuZprmFs7Lx2OQIBxUHb
XvRzyp1Lm8nkWyzhMtZmb3w0OEeoLHw5McUgJ+2aZjpzsBR0ytvUBR5ZbEY4cX2U
U4fnHFXFaM1dLaMVYCO9ibnqHoIaFf0pAW3tRfsNGaE+Fb960H2wOMDgPpeupWqZ
AnZfWiaJejQ1WDIEN2So4Qtod5GMQKna6Gv7rEJ8UbZAfbw//bkzhkbKp9MYChLJ
TgXzNhfrM3swPMHufCP318CWbuZvHgdO9cBk95a3QqiPddjnHlP/vQ+LuCGuRqp3
e+lONRVzXK9QvkScUFzYmcOUkWUaqL1K9TKXZ0jwNSgHo7ljJog8yXA8i/BpUa/h
wSGWzAKyZCvYkGjkIUIOPqUq/FV0bHahZAnB3mWDt2/0Lwy1wkcFQNFaUqLxzSzh
lMRYd54KEf0zBd7yXyK0noTAhh83x1BZzd/cjTOR+5c6repJ8T+Hn5VuXj9Kp5zq
s8GOjV5/+cYbC0csJH/tEl56bctFvDw45n4uDoyVqS7aBKYmAB34NdnQycQ1HmwL
4eCL/hLp8l41vTH7ZOCwHhkmKiWcyF/5Q/j7Ncb30tzcrpCQhB7OC4sJU01dR4jY
SIbN5KpW2Dte2phZUO7TiRW5j7ku6cWNZnKWn/R0LFYn2Tfss7g/RIC2Xa7r79D6
WocS3tHPkfQzcaxdZqcpPNFUBIhhBTRYcy+R355SRm+iqh0yR0DE7ln5tTVPL62i
AjoyWycifPHYYF8kUFdMueLWklGqKx1584qI0mTcY9bf7Tcw3hA8ix9dB/sWVfAv
vWbY31jLKm27Uv+8+LHOKpDuvnqX332EFfgW/Lx8Tgerxhknthl3gNliWCptVdbp
ekswJVVsTtPQkxj/H8ENZ6vbT+q4pMLd1asLLN4bqrt68tQkUX9hJ/+60+a2DqGl
PBkgiu1sGCAOfIAXz0K9L9TYg4bVstPpxtR1V6CvyeJMoc84s07kj/96ACTX/qu0
0TinBgDT+YFCuDc7qcwOiaLBdW0uvfyy5hKwy4ip4iycDSa5VsuSvvAlC3r5FtV+
RhlTHzwVX3rJq5+nXoEppd4qtbfBHFVPQJ7YTTIS69JDOa0CPwvPKB1AtgnfUon4
ugGoDmZdta3fvcqTCPY+mg8qqM3U4jqVtRF2Ed9SZO++NkaMLiwTvv88/jxtT1EN
f86B8l+d9ZC+dMeg+m3JVM8LaiNtSGAJk6L2CYi8lcZSHEUoeSRhRNntoXo9IBEN
uB3XHpO8tF67wHa82mTyyMPsuctuJtwS+hk9s2OBzS9A0/9RwDw4Fb40SxMH+JLN
96PoNLLpN17cakvg76+iir65Kj77ISYWsY5KWsgYJ8118rzUCZ0etJdVFUrkedxf
9X+W9ExnLyTqS9qKfU/0FeP36oyFCCKRRVJc1Js4QXYfDAJfj2HpPduIMMFMtH5d
3XUMlnpU6Wea+U9zQvStbA/EWR7IIJd2m/ISej146QgAMgQELMC5NU/xnzjnA3Zj
FV7tMFO3IUPhsVu8fi3Pq6vDSKZBOMYSHDyfhzmTd1koB5EppyD6hWImodZFQYrd
LWTft2vf26qRM1sVA/1WslEEo9+r7z/sgDI0EH/ktl8+pVBG9NO4YvjldD3shdFy
IFl9SXvLU2Is3milbBRzbjlRXgwZoH4UoY6kuPHU8dnJyt0qpXUaCDNXlxrb9+DK
jV/u5RMhDVaH7JZBfD6w97jg4mHkGJz7FSidRsrd5GbyqpqHj+/UQFXzGCoTTbOO
/27J8ieDCqApwMj+tzK1XNtS02vETpX7+Ulrvy0cwY316DD7a22szSApBYMk/o41
Nj4tGaYOznymiB39824VrHoNKpvL+vd9Oo1IX0lHHzhsFS2beBMLN+ueza8Kn2+s
AS3EO2y9I9KXk30RIWGdyfVCepJS1+YHwxF4h/xLXbJrF65eFjn5Z6kc72WO0hc1
T/E7HmGMk/AvqbcEC5ypzbNEi0qnh2cY4AHV9uZAipkmV9Hk/Nvy5Ucia00XFwJj
/2X41tZKc7QfAD032s0QGuM4yZZk1ocqnxmVpJXWb11/LuFqfLZhKCvQ0IMK2VIC
UqQ8HgVvR9O1Hok1nYcFM/YA5eG+ipN/WMcZkB3OjjqheabOu8RC4JMA3yukcHde
KBbcIfawlKrlQkOaXxJRr11qGrVDjc/53BywYwN9KqmkS44D69YD6DY8C9VeyWE6
oEzz1mnd1ALXJ3MgMBvwPMCMf78o9++bElG/jDIleU1uIyA0FuIAOogmGbtnHQE3
ftMJDj9jsvbuBX8RW/hTwT1DfM52I5KmMIfCR8Cf6VLezQuBmFadWlnAIq832yHC
DACbE0H45s0YF6w39aP1ySQ/3Jydo+OdyTn8lC9zxyvTt3J5bDXh949U37TwKB0E
c/jdN4N5bJdVTBOKvHZ7QxwDlDM/Xcl9n7VibCq/K3SgNUh54Wp7NfVkZ+TbmCHu
9I9uXNizQKp2caVgnIesPuUZroTYPyrbxhoLodY4B21zftmwWnTOjzAHlU6nlTVr
Xhiuo/w+ZRPszplakj1Se1tkKS3+dIJ6blY0i3zxMsbXEFP5ymvGEci6DO7RWS1z
/hFsqblskkQ4A5N0MYLOnVQt73vrZTUeesPD+nJK6ALlTThSMELSgYydEFYnbe2D
Qjvc7XSLeQWf5W025Rbc/RT5YXmtP0381Dg6zBozkKFzOnTLVA1YM+bv14F3xoSy
8My17O3kz1HYvd5BzTznDRemjXz3jVi4JsKDHDoJL6aEeV8QbccGbjjL3iw+2N7v
DMM8L5w9czfsRwFYINM/DSxcYOL0LWmYJUAIkRkiA0n/6NCct8VBn/TDqBMkB9uV
ZW4Jr6E71BK3F2qRMUbwXOUscjHyDuGAS0BWijsNgCpfUJYQwpnn8dIdGQW4uZCE
cSTbnWQt2lnXKO39qY7PNPAoALXwD/j0Snd8mPEJoKlqhuxzVWbKmb2qUx+fDJdG
W6B0aRFNSduE73WQLkiP0Asr8uDGcgxDAY4YQuea/G5MG+DhAKeGQeSsZDNS+E6j
a71r6mA8BCVFdimQ1LdLRwRVOA78KdWVun+vK6p03YzW3mJ7uD8fNaRu10dFPWk3
qvh8QlGGY8B3RAEyXcKaCWW7VoNRJtzcPXME5ITnfyCz5E0iJlEZj3RWl0vbEOVm
jM+YtGXwuUJlTStgGmGcA+8TC5HQ4s4U8Ie4vDULkMn7BW8k03GYtLIWn2y7AjPq
yKOb0PJ4tRepMXz2l2MzN+oY5ADSh/yE1xyJeMxdJ9LMjZzwZwrSSOGGBJwmWTVF
FyfCt8RQUZ4nJhOwe7hpFJvkh9FBaI4QmHV0Mm0CNEoIHR/i69xg5sXinJenGNel
0mcdnfIgF8OES/WeVAwwIz2AYbzUbC13XsYeP4JYMSXmCtcC9I4Wk3Ufu9xOIl9a
FRHLaxZuaR/TQ6QoQk5ZTJccJUzdrJkt6MYO6k8UAukJq9UDC9gS1Bw0Mvadl/pa
/XzI4j4jYhZuDclFQTwJZ9rS3kceNvxvit4iv0cRBZUt6Ft/NMGIoma/WjMYKdiO
iuPP9FFeGtYRodgSuccohltAwjSozquR7u3OjA80PV/iAQoBhNi/Br8Qh4xBMNi1
hj8IepKOfOVm2nZiiJKlqbUsGX7/bll+QrX57BOEBxVo1vbOcxwcONbHEitka3fB
h06UAKfz5ayLR7PyqJMP8DwzT4wbC3I6s4/buDACPKMes9en3b/tofsqu2HKV/kS
Do4Kukp5fS+z53uyRvWPqIksJmGs8gNznRVOvkXi6zav+XjvwK5twvLDi3Qm5eXh
50qBakD+K94ynWjqvJzRbmfxjUmfAgYvzegL60kDh7kLeVn/+f0Ny4lqdB7YG3Lp
Hw5R5BISVrUQjqQKd18nyqkk469NAmYhcEYQwAc2HoHicrokMdjxOEkDr1m9LjSQ
VE3I+FP8MDJDL1WpV4L98GN1WwYykOodMdzFqHcMai1ZGiXnaFHoG23skt3pFDjw
R41sshm4TpMWpuDWQ1/kT/nG8r7rbAm4pew7AjvTF3SZsM4/V0PArxxVKhlziUtb
6M60JNqjSCB/AgkWqbJnpDHGfUiDXFsOOdoTls+GUdAw6KEOdolgTPqG7dTx551E
CQY/rSQWhJyRsxHPW1IzoG6pR03vPpxVBWdPwzJ2zX01LA6pMNUmuy2xzG493p7K
/Co3NSYBFeIC7+E/ZcCBwZ4WXb6xpkUnrToIxtfoINDZUvhEHkWOO4GshVphOY3/
hReNcOY3/GBiRRJ5Mxhbb48tltonlYEbg/NQgMCD4fN/m2iZtB+1WWe83e89nvT8
DvhvUyIEtMmePxq7WgDFS9QZVHcXWIao5k4bd/abxnepUxxgum8DPA0qyRouH26P
2IHTpAkLC/2zjpm66gCRgkWorcwfKsh7nuddlfMIibfoyWMUVd5nnrTiO58SNNV0
8kXukK7MKkpR5QWdiSjVghQ42oJJDwi2EIF4xbUt2UQqDvrEEyD2pfiOucQGd2F8
gdW6Y6IBs9N1ndVauJ5kcs+fefYolmzd8fJ7kdkAA/9uzab/2rQPdHbAZRZ2X3/c
InNdS8oWDOiomxTmDG7W43R0MqRaFIz8LKvwznQjaPxwGcaPsbWQIBlUg2yOLYQD
xGpWMDZb1V+Kah9ID9YPISrbpf68EliFCoYs0cl4rNzsM0qaQwp2t3xuQyf8dM0j
qet5Mg+Z4S/eHHYK406DFkgSkFu96FgssPk8pcgasct+T8Ja7sVBDxKYy7/aX7Sb
1jZ00OKotUao1IJ4B8tFIIrjJ7O3UQtksJHaCNFGAOEaeuEd9K1bzXyR/JW99Ra+
bGk4ecbw/zV6ZllGufeBlx1myLS4ElRyQfLfsIJrTOqQJYwjiiXRWT4Xx4WDusCO
O27/PKIh2mLBQQ85xaOmQW3cK3G1jR5HT9unYy08lMFZa1RzDvrUD3IdApXOkoiB
tUsnH441Gg5+GcFUQLDaMlbkVdEPWv+sbqhN6keZluSZa7JuePDz0KxlKPSrB7aZ
CWNPxv6BxxEzEIdWUnAdnbX9QGhuL47+ycUY8ZPlrhY9AdTxenNvbt6GyzNuKqfb
vHHWmgTkjPloEXfHewQIVq9G2TZda/w6WCTnM+rdgm6lQ+KBJ9IMCMBLRnRnBGLA
8JGyxEWfUibg8fHiKQkZqFygVX/zwcSPVkVeEzhcadFcD1I0j87tv/PPRIabH+76
9ctwdh5gC62tWa70dqlSLMf3SKa54U94lDFXQFWuAo8OfO9m9DIYsCC9bp5Li/qZ
fSocn1DrPvdPxSsmfEdLecqCdqVE8OMtcd7rZ1dlOtwF7+uNMPPMRBGaLlJVczp5
Wne5QGSZvSfbLEQxL08dWPemjAgCuSZ+avsElADxW2cVUYrbiS8jvcsLh9d7Ed3W
W8blIuWJft5/pfbk4b5cy4LEVeHdZHgqlSjg+5ILGxs5z8XD3XTVU6He3lPupySG
C4tcWyismsN/cT57z0ieAFvu+EtJdGI3SI+K260XdKWxeYXzyG+5hN8c6bEE7H3G
21jzHkDcm9LX5izJ6+j7Wu56XlluFBCh6HvMBVNxkXtFekVKowyCT4dk1bH8zOAc
9dEWH2qfF20Hk8wT6TSM3tO3YZIIUe0djn7tvfLHr5lY4Qo1AhTGXVrVnlAy5uxw
t9PDEIauN3wRPw8sxG9qE0291M+FNp5ic5GMrTty5KhENPVw/RCTYaseJSpQSLgr
f7dBa1hRCnnTDAZVI/Mc3Aiq7yGX1yWFIZQybqA5oLL2p8fYIYYFinBx2VtGMu/R
+e2gp65mBE2Sq4+abQYbK1GwfE57zcIXwN4abnLeqWnGBZT6c4Jqv2EvuLrtrM9B
K5dWMpeJPYer6VybrPiYm+YQ4gpW1IF/y1Mz9KsTM0mnZkZR4S4v+O9Wx82eVz8y
JK2tWEe0wGUbxfA+69MsvSdG4+ocBrfktB9ESWUF25uhwiIH6mOEI6Qg84Zw2q2x
dwQzf7P6tAOAEpSoiehcLashOYWqkkI6627rqyWisFwFDwI/tvlaI8BHCB/Q23hX
5n+MvkN9ivFa4WJZ+zPg61Ttvh9X6gkbeEjzGaqrdZAGcjaIYYp6Gk+oY0vly5a2
X+MQ6RzVIuA+hMiqnMnMwHyuL+IQjC2rLtRAOh9xj11yTIVfGDM03IOxsDmVtu6f
KDazgcyNb6s+vpgYDG80MqpF3BJQIgxc+yAY+I3o/FMgOWUEfDazAVM51Z2uOeiw
noEYHqTID56llF5yaS29CMggJ8NJoIiNQIuZ1e53Z4ME3b+19HLKLqgS+guIi6Is
GKKS8or8j/H8BDI8/x+F/DVV58A+avsd2BOSc6iCW6nDcSVAZHgjf1JQMyYnCv83
Q5uupIRvLLkKLjoARgGnm74PX2R/sFINmq6HlCdw6YPQyW81DlFDNilTWE1AzQyO
29vuDWjVQG2Dj3BUHkxsUM0UzAs7aplX8RkJl6gIzUX0zbrRNsxp7CdmT4oTivGo
4hQp0C8+O0pAbcVuePA1qZouiJ74+dUIHXMhHnmKahATYw36L+y5firSeI2XAJ0r
qFGgf2105rPb7A6W+G7j8OVM1QuPNKNFPxDBc534xGm81d9OXKnoNexFkzMwDPpY
UUe3xvkMBYJoLXbobbyy9Ql3z9sa3O1osEucHPvQsCwjl/8s7IojkGa278pebiJM
8TrVongNhx6K8WeYcxVHXKGQRwcPBGm0VTQPFdv/eILB/7Ezchw89WaolzK0db+v
Vz5U6s3bSvwQhs2TOlX4CvCGFkYsVbszs/nEGBYKtNKkwUiYdqfGME5WGIggT1j3
TXc0G93TRkqAJwmQ4NlKQg3st2GJ2EOA0wOHHfu3bp2xrvYYYUhjLzRxHyH7LcwW
CWAtBMqxT4VehviZRgPRlQADS/E1NUlhJpjfc7lstWGLjB1PVQnw5OUECSkeryJu
7fvWIM4ES+jYkH2AwhjEoXJbOWA1/PdWQTBQGhozjtFSl2TbRNwuv9HDvYEl9vUc
cRko/XIOso3qUsQlLSm4admqrfefwVIYNdBbO2P3GLPMSwhAPKkh0V+QAoOWLfLx
Lie/whAEjHOAFU5MOeeJanoAKu05tAnDE97vS+wyyioFrFaPTCjTJuSv2r8odFC2
gFuY+p4Xmsv3f7WXPNpC59twGCaMgNwlPNuYbT/dYPqCzsOJvG391HSpCO3swDIX
5ZOlLpWOGOFTBrkAH45ChuIWW43r8ZqPF2AqxcVnKQ02ZYra4iO3DWilEewcgKht
qLvrBKqNxIFgaNR7AKCY+qJbLmTcCnDAt3W59QailH0qAXG91obqS0fSekoyGZib
xiZOVKqek1Q7CchXZKoqpTCKZbuB71CjpZvTWGvUcKaJJozj1IRecXy0RdS9al1g
0NH48aukKmyBW+OIL2uVA+OZL9wig/fYVaP/GzYhhVUEmQqyQJ3lSiNeOp77wiK/
VO7OTkuP1wRjBNUADKQ3GK/1NvDxsvZqzlHNyloYDDknMODpjiXHSQD9qk/w1Ay5
BvqZ5Q++N/aOtQHlN9sZpd4/HaIhPEStQYRqr4XlGbBPXvaJ+PxULh0cjABtyK88
AibrWRtTB9z9LuZgpfKvf+PxaciSf3jMf3+rXqcwovh6p3CkLp7U+Oel4ot9jiBH
9jd5HMTQmTANqWZq3UgsaqFJNP4j2nGSMp8BNJDBKzk28nHE6vUve84bbOmSB1Pg
wPfMo6241MxewbDGMcQWzdD/TroE5x454S3yZ46EZCUIxOPzyuLEl95+7ZSMLWsi
PZTRVDu/T7Qrxmp+sDJHoY2DIOSvIA+lVL8cuFBp1oSRlXgBs9ePQjrUPeiVKMLI
ZuQ+o9yqPUEWFiWZzik+Lc/TH7Q3Vx6QVfJhkcj0rsYNIODKCRbawjUeACsCVz5V
RD4TpW3uO8sRrEdEZAajaXNC+85CSGkWmT1aTHRClJmPmM1Q4gdt6fjKrMBUf+mH
q+Z3LL0laizvsaPFDfs2AlrULmuh2APzGNje4m2faYCc/Ih1sjWxOFuLt++ZrG+V
j9grJrXiSdsZBdhXED4p/iGj9ioyovsh0YbA87EWe9LizajNxttcn23hEkIymBfP
N4rLwa0MCBA0ayh3f9wmAXj6C51wzZs2lNwA0DpXLiZAJNNz/Qp2Qk7MP8R4oXmF
kjgZ+Lm+HvWd6xK+1qJY9Ar6+Cs3/0TZadRrH1jXJXXUEAnzqX9+MKbzs3OME1BC
JDLuNrxF6G9tUVEIgsSsXlqPRL12YeRd4jLOG9Upg6IXolZ9E6LiY2jiwyjUtTLY
/lhYObok3CDMNvXKakhhT9I+dlD+/N87YUxkS04BfLR5UXo6uxOPd+7fcUPjM6xq
TwtgYkaRquehLtuoEAoG0HfKW4dqXxTR8Ciz1+bFLL8E1DHGakVaNbWtoBhixGu/
LnUEyiCsuXS0Qnx11brZEdxh/0ziQf6rYn8HS0uhfvNNDYr9aj1DYb5DyyGW9Fhv
fhfMVxDI1rMn6Id5lxr9x2XvBfQG8lmiyh6RcMZE80KMcpkLjOuuArgLdkVbActK
v0fpVGbz21xgg0jNXRTDOublKY15Bb307PEkPpFnDZWlUEnwEEdDi6d6j1IpruRs
eeCpQP115j5Mlyb8v0xhkQaLuWHsyOOZvGzhdOphLREKbnG0LtVRfQMl8BccNzCv
kLbyfym7xlMrrJ4cvUsJV31rawnjpsIJo+JeNK3E/NaVTrGZYM+B5cAjisKIPkpD
/k125X4Y9ak1SZvC0wleVinD8wh93T4zVT1Q4nZIp6e9dH28Zc87lowf3K8aDB9U
JNnNWGo/iIWGRqsCYsFg62Dwvor9Q6iganAwTzKfWEECTbVFfhWEu+vIiGa0NUjc
GuljXBwIA0vQLmosYHKnlESfJo28S1sgZzv/YjtKEyeB1Eh6DQMZaPSJSt1Y3UMP
1YYcy2wFjOAwyxyxDEEOtxqQixtJ6eAOnT9xdyOXR2ffkG7DVYs1ywMlXbZhSh/0
ia6uw939HKA9Mw3zPJCKIBrczCGrIea+VrXI42MbEcpOPYnWxszIvG7t/sMt9j5m
h8qsPCpEOePUiBOAcHR8qC05MS57IH0JUglSoKd+wZihsoBSiv/RY1SloHu5d+YT
doq5brT5bU5D52lvGLkBuSvlQKjnaEV4bF8q48fHictOiWrEDzP4n1qJRl7xkiAg
/UTmjhHTgEyWkojt6JQyCx0B0jpt2VOvHqlG1ZUOgQzEyrzscLISm/4zgV5GCV4C
qVAVNFtdpZEYZwTKXmWgOXiuoYIKbFECn+THyspyOefuZvsJF2nDTI/R+pgpAKj3
zlgVsUrNtzoQ07cQcQdoWEIZ2OiJwQE4skXFxnVL5uRQq0BGj1hP2G9r4FyaMaNO
HqpI7DXTfXqtC0W01m6uYrQHZ+l58ume9anLZpuEZerBApYyPKaH80ZgD8sgQa73
JbdJUy/6tRPlIn3An9dB3yUtBLg5hOjvHkd9kcnrjqPNdANSD3LBLWdjtxoufJ8v
ZUqT8oY3tgYNrNiaRo+/WvOxcPJzt/5/x+M4ToTiFf9xND/EOa/CZAlBeFisu45P
qC1Oq2/2pq2EoTPh2uN5hvzmZSuiyiKAF1QhTrBvL3LjcY2aPHJ3qUY885ZMCWxF
SL3t2vzLkhnbOHUZVEx1Ggq6wPOYAparS9s2xVnAQCov3aJmLEPrNA3xqb7GuxkY
cJLkv8dwtCoadDULot6VASE8TMQszyYSPS8m0B+NBwNgKOm2ouQO9KcxNIkTDKmk
Z7RPt3MFfvLJwY5RMeHwKBRocvXrQNRVz2coMLoIvlAmYfYukdIDq+zIRqCjMhWc
SOjZMwPcv1u1R3mijHf9Gs26OZEpSL/OdWc7ndGkghJFpWFIxfrHXZdUGrl1zkmD
oJDYJVNHti/DuWygzExEOZq7vFb4nsiQVDiESCZGPA7ePhz/QSuA8HdCqHYCIcyX
EIbVG1dNSrPTP7rNakXPZBMVo9Oly/J1FTB4ibs+Sdw5HYX8WB7/+MKDI1SqOiCF
TWwC4lv/rAzhJEErhiJZiUlzTP4D3/i9a3rK5+jCAaquOjUcFc6oHskSoPSPr09F
VYAC1lrcESKqp0EwSjfBYNNkltu8e1tDk/v1etBGvY9rLaVfIE/e7MQdieQ2XxTU
UsARneZLXo5+bOb59lK76B4BW6DlrbPuAU0UXZJEreTi5XMJ/MgW+MFyB+7V4BWf
9rNWDE4Jvpwjuk2upE1XD+Mtn6jssTeGaG8TwrVCkylb8qcFburICnZkCVXqjJce
kpUtwDAD1S5vbVW6BU2JHfkd8vpM7Sdp4exvq9C7d+THyfN6bjvb74pmzXgxy8nX
vAuHG2D3XzxWbEMT0bsHlGkJHFhbuZqrwb1F4ev3a+JGBwbT22dKXUny2On/KL8z
SaAxm4kcac+1rGCFbJV+EH4O3uT6R6FF7gNp9j5Fr5Haq2ZHpU69/Eb9e4MZWETZ
rLWXeeLUrnWqnYLKAWdFW0h+jAx4a9klAOpXBYK36RqMkk2K5EYx0/uJjJ1TzlJz
R7Ex0sPd1HiCEtFSWjDG58pkNceBYXDQ87FoX8pdvUIon8hTZT8woL56jyJejKA/
qobnAqnByrgomTfGfkgc0XWY81Kn/nWkVabblOuFUdF+cY07ZfXCZ9cIKcNR32mg
RCwYBcoSLgg4Nd9Bxpy3VWW+WRVTtYBc5GXu6/KLx9WZCR4/MS5cRncVL3+cR79E
9PJbBwqKKXqi/XRe8elKYYJvC9JpD3KMx1BNr4VXjaVULcohHr6u6BVJwnadJZ3T
YSNZDtMWy9L2e/ZY50e50sLKgUKrwoRKKCkWFEUS64DnHMCBpCKkHXghWr28Iiwc
QnD0m4VvKxmkOjRk42Db9iLtfKPLHrL3aSECf4u4/IV+bpf1dd4OIGmFtI9w9IMz
p41hDz4RMjH9+gMhPsVDOeWyQGW95f3CvB2o9hexoOFSpdkEYMal1SDeWB+aNBLR
nWkjcuHsu6zcCJz1D3gSaF2ltTAX/VoNNAoqVX2m+ZWnuNgrfaxa/TlWdOF/CJGt
KiT5A314/E9bIvGm/tVNoK5Eus2Vd54GRMmFCY2HKDDKdQ1zLQAq3j45uIHUbRtb
Zru7prIP/rLxFj0NKxK4JP8hZDlTRWvo5sp+y15LBQh2tFy4tOjsIjGzXi9isT4f
//nwTyAvRpmhUQgRcb36J1/Q+gbhuxlwfRs1H6TZLma1PW2RkxvIyRKGcs/jLIwi
46NtU1LBfLVNjExn5dI4l70q+UwnPp+cO+DTPkkIMDIcGMe3XC4izFvab7adzCEO
FVFzt8s1dn+apoxpwzW+N9n/vhUmi6VMPbErWhYVnaG8vRUS7DX1TtvYjCtAh76q
G97obWsk5c3YMcPOd72W03u+oMoLkAdjKZE6TJCnWWyWKzUt/D6+1ibONHCdcwgg
hReK6selmvEL8IjXaDXm1lqa4n5DY8xeICrjTMHbtKpP03sxMLOrMPMRYIR9RKDC
B3Y3J8TQvqwHZ4wDHiZSEaBLRXn/AX2cg1AuTLIeERgqtgWlVj5yVtUKnE+mxzYr
OwJ4cSV9LY4U+AL9fmAS9WEQDPEIs528ceSQKJl2gqr7r/6Mx6ZvzIfjBKTqxSCP
/Z9YrJoWioRUAOym4LIVulk5AV64xhUSGmv6QUqh3ikuzIasmuIQiJuwhYlt9Ehx
Dl/uQSPMWRvj50coN5fS6+V+YuHRRvWCfJ7gosjPua0oXDD8zB6LFb9ojw7TRZCT
Ky/xDLikvdkxHGf0DSdjyI5S2R4GhjeDVgKy+ZxyZ1k0IzXGfCUg4qo111BUZIba
ps7tbYWEydP+XrqhxlLsE0j523HfEE9Rc37B2yUl4sqUqvD1BBn5r5T25vyE3/Ws
JjJ/+SRpxOTEhVuJprvn6oiGg0qBWwKZzMQc327ejW1hJ2IMR6yuZpH3QnTyGQG2
Quvb8HSpjQgQGJ2t1kjyvUAIeOCIM8Ho4mcZ6BwAXu/iIikgMCSnC3dSJx82eZdo
dIURzvKl8EoPG68+K2CK4LKYWzTgiWQiTW8exdPSLVtBdg2CpzUI5cikmTyEZPIl
BIkB8sOAEMuFbFZr8FFFPU51NS3tvAEKdV6ki/9ihjTua2R/sqmkAZPZOG1akiEI
YetzOLO0neZlfjCsRgMpt6Y9NYauRvIXASx6IcEWqHuKqG9qcjNEDJmPlh7572vl
hXGnfkXEQs+e7huxJQwdezlPWbPTeIAOvnFdSmfzu5KQt4NMjdyjJnD2ipKvMqSX
tT5nI0S/2QHWv2gt8INIOuYbESkDZZ7wjE+JTgKnRCV921NNwTz/ovnEaX232zt5
US96mBYH+GyTkw1Lw1NWgMjBNLg1ngEvbrl7sNP5lDpnsNr6gZ4lvvKWdvbwJ+TU
c1tMbRarZ2R9eZzuMI1HYfN+O+C9ULg9OqwI9DqvlN1ZtYEMWLgWVghBTGWjSzQd
94nhxcUYmneZoTfpwvrTmAv7EK5Q69Us5pw90QoYzxfim9f5JxAc2FTsJuSLm89u
dq7vgFd54ILEbqDtdOnWhXYGndjxQIhQExcF7rnllPQViMzamKHb9in8TYzoICnl
q4VbKy77CdSh9QY7BrE8gArir5WatSs68ReDu6ZaIL7AniUl9/s/V8unFQaHjWyu
XeHhoHr6mlLV8mOaM2Jl92Zwf+pIi4jf4er1O+FGGxmlqO6nXSXw+y5Q/PfAkpdF
jEROgCPSSCMT3yxXEac3BZubx1/MvZ/hHZp8GdjQEOLLTeT6ieQF0VLWM9u63+fe
fOFTDuccXxxWlV+y5S5oSu/QsL+A9rYeQ90BO3daZFumaSfEmD9a8/OtuQJOxtZc
diwAw9fc2DMwtocc2vjtjyLyFJGrBjwC9mBWnGjzdXBfE+CVSXntzyntz54/GqQ9
mxRPq4KcyO54PPdRXSp9Y3FDoOV3TfOQUjFDvsdesB7jV9wLzBCYAccVvBHsVcBy
Z0+x9jBWhFWQiXN7b3MwI4FnTzhOwo/Hc7T8BdAhnsMmg3Mc3uwBnitTX5/lJvQb
6/pFBkkXL4TQSGYgOJiv8diQBy4LHYG7I2UNDXfXxG8NLHTZv8afuBf+oLSN9aje
/hEqjF2kWFVyxG4+6h9zHZo5o42v8daqJKWkAB5xyot7aBeC2XbSi8BX3RBbViQs
ogGN6LbaDuQBiNnxyONulxOOq/TFb9/2qUYX0nwyz7g+X/VL7E/QdYIM2/GH5Uq8
tvWLwH7MydnleUTXnCGyfCKNVaXAWus+sXJQWoz/50y7LzgZs5WvKoIsq+FPBwKb
G2nyCBHVZwWNIJ8+vJZSL6X4QypA7ne59Lga/k5320VLkMhQ6HFDNsIwuJmQ4OM1
NPM/z9x6h185vxVGAu/VsF9iVDokvuMgmto2VTSfuovhM4tjuWYpEjWnAapyl5jX
g2yDjKxzI0bRZj1fEcgQoeSw3Omn6LB+enutd+v1hYD2ovzxSpGbpl/QjlZRLLQh
rKU1OzAKnf02670JV6CSSUtHTpEZdsPgFd7DGjbT1PzLIMfxOU/XmDGfPRWtdD5h
4om2GhKPNtbHZ5XG70ZK48US2nWykyBE0FU1I4YVVGMVEABvTTEyrNXLKVPWT1uW
MRATSGswom1nQlt/6gj/UfP7RsBUMk8vVxb1U/XtSKv0hGyA71hXEJGhYQDxC6ek
b9733yX1TVuj4Tbk5KOwxneZtsXDKriP19OaNVIe1MI7W669muk799NxqVPCdmoG
YrsVSib1MEWkMqqkHrcAlwzrtmB9dxwXBqxqr5dxudI69JzMq0jwZMEjL1wfx13/
a9uDm1F5RYLnJRex7yokcSk7zIRpO/xysrO6Bq15egJ21Lk61spFA/WiyXeiMcUQ
NVki7WJbbDGI9DxAMXXC+0PV0AQC9Mj+tQPqxz/rYNo5Qc1HNbAOqLwVxOIYcU4C
bLDSU09AlNe2ngj8IpJliDHox5/CbwB/z7wcA7nzPOHHHvNdBF0RND3uQSuqcTAl
sHrBNUFu5JFxOBlgodUswBR9twF6j1jboggI5e6zE9REWYmVuEskakLp82fvV/Sq
2YvtcbY0wiWt6gMEqoaRSOAApsqyxKwQeMWbciSywGbWEwivRCZy/7tOWZsLBZkc
/EMgMTpPSbCCm6D5VjNr5b6SHQZm3NdoguEeQeyMX9eDnr4fjm6Ynhxfih/dh349
hdJKEo31pQSudw8VdDsm2ijqUdvuobT9wB1XeLvhV97MexpZ6HEmCF/zunVIS94A
zg8V8L2WxLz0ci/BhWNg9juTu7i/hV0YtzlpZfpdcp47pxKuUmigmaCPLzQi3NdI
AYF16cXldezApvODn63SsVvOs5a26sF3V0xq2hfifEa4qHcLp8Ylz4oYukryE4Ye
69s3RK4VT+ClVam57qVe1Gc+HsKzsz3R/HtlZTA2ytF7jJk6TuOhZQ/xf/eoRBYv
xQ9dd4A851Gmdi7VC5h/wpjo7ICv23JaP8Wkcr3dterLD/76FED3UJo23tflBT+z
xFRDeceR58dujwTxh6VZeZo9wrrB3OORe4bRuk+5xfrLruzQYC/TzFImdRZjprZp
R50dYi2m4E9hXYcG/hpsKJNrubilkXWkNHTSTs8ez3ZQzlSBCvlD4sLzlRvBWm9N
T+hEmRCNL0Hh4ec3q9GSrnDRkZ+3kGP/gKIwFVQJeEoo+q4Eer4tytQB9z52kS5B
Tg1YrS0N9JcxA56KKYTu8vVF3heoP7zDhirs72n8uUumyKteHBL+a6z+raHfGtFU
97FitUs2urTBBWtxWO7DUoMIRduOjWTX7Xq9H7ru/MiIYeE+weXdPRxLRre+HRBq
PJhmtvRlo0xjUhCs0EtuZbSMajNHVSq3KuyWSANNeeBKuN8mKzbVp9Plef9c8wid
9GdQbGqfnWTU3zkeM8wN7sajWYtI6Psp9YfV9b1isz1I5cUvY71iIcglot5BjChg
1D8Qx0mKUN1grsmbSFdD1fOtBSypp38b9SXCsbB19/7EdFAJ9es3RBOlrjHFZJVV
VkproeuNmCiXlQhY6QWkfQFIiB+f8Xz5/NAMXDy5904e6UII1KStWR5D1TiN+uCd
ZkTsg5T1znBOopQYt18WYowd/fux+mEtD1e4azFzWW0aX2N1NKU72WXx6ewqCGcR
GjPaV+w7K7BmlvlYs07Ntm3hpndPMyFogcrWiOTUg94VFDNMxasHLJYE4i4AoeHA
CpGFasrYWxYFwraX4byZQ2DZSoIDtOzDzp/MpwhgayMWzWFBWGd0FrBhmz4Sao9m
JN6mlTcKNVl3K0aJJh/+rF+Q5hbkhancAGH3PwuhQ0uX8kWJWeE0BN+1fev6Ie1J
jEmQsrB7gUfx/8ik7bWnGxPZgqYorWTyEgFk3JzXRd06FXeGw9P0hGxMzhMgau9g
kvKYqz4uSaW49EcHbUN7VsuE4T8IRf8eJgcbZCEPms44Jyj3F0chelKZ+wdW9rqi
NBaPSNmuDVGM1ejXrzKOK5LU+h0ZNdJSwyP5UlJRvqwfpydnxCNLqPqsMhTVfl37
2tHqGxW9bO/NmW8PoN4KUEMi/q/acv7N0Ltna/gC9a2Ie0nK6isw+0S+M1t9pS/A
ZYTdoSvq0DUDE0qTetDyevVPxbMLn0lSBURhokKQ9DKHHnwJQQ8V9nfvoWWIyFea
UTKrM4r7lEuiKTKbbl6suY1TLbwlqj35zaZ+kIAb8GWNC3DMtgTA2reS2WZ3UR+/
v/H8fnVCqyNfZZkyJY9wIRxgWFj+uFiRYO89z1Z+aSAUm6GSWHF/lRR48GGCe+zP
N9lE91YGKbqLcqpViDQy1kpdDwzPEqdAXJgpyzfF3epNGOUKg+iJ2GMIOStLpQoM
zZyZoUjhrYPFy9i44cdB/GtUJrU4zuHWj9G4kW2dxKew5KG/2jfLcGtqY8YbOx46
mOS3kNZifWJj81N8Pf5NmXyMuPa+iBvhYs0yXzHSjvhTNitFP6g3KadV7yaUAVkm
vCb/91b2pc/TxXq7ZTExDT8OpHBprTEuSKoKCWJgn04a33KOTmxfsIThND4VfIqc
4smA69aB0oxuZ/bIqbUXc2jl0uPdSZxz1uNQ6/zTe5G0mKw16BhS0HZqsHTG5Koq
MvkqgmN8vS4qEl2HRp2AfPeBj48VvUhkf6rRyWRjou1A/Ys8p2a0pfKfus9YeNKa
mBlSg39OhKHbRSJR3NkXgQ8/es48xLlD4SnLumvsvQ/D5yO/alqrHg79ip4HB+gn
9AFTUHBPjPVA2YvzqVxca1s9F9bp/sBeEjnEdo+qQn/gOHjTuPEA+nGNiLL5pVtS
Y6lDeNo4Tz/2sGRf9NttOCGouV7/qOS/NsNHIopZrzi0fXkLa1wSYYRi2OTlAS1/
MySp0VJZwN8I/TihsSus9AeiBDJB8Oa3D0/std1ekPyg3WvX52dBPKm/5GrmB+/N
8AOzT+NFk115DVcZExCywxjNjops3EZoYKqRLudmVvruKCOzktURthvqZeUixO3H
0aiUsVeBIOi+wrxEeooqDujtRTiwGfH2IKgmTWXRD6q8WUpL0QHtKpGlJc9s5h7q
/tcRpgo9WTuERq0uLsUUylYQp4zdtPGSRXAIlFqZqBv0ecNKV4ZQtc3j/D5OnUnW
k7wj7BRgmVTW4jj5Vylfz1vdoIbLP4/j1Otm+xvXUiC9oqHVGUPTVO7myTHaRKsr
pNebbwb4XN562Zwm3nKmFVZpu13Aqasq4QpRv/MpJ44XfTzzk1+VjJG1JfVZxRrs
E5zFsIgvuKhzsaH5Au5r1IP4JbVLNyFhzA6nhMjZDGSxCxoa3I0gpWFRovo2bmAB
tClenvbqmNJLD+5P7isWlFJqBdHgmefzQ/KpaDo6nzjqsSAz1oYx19ODap6CpePo
ZVFo6zWFVdgE3pVmaGjIkFFIATHVO5ylQfd6f1gAXM483BMbcV2tmuo4VDwT09zN
QIM5qdsuiiRn5aWUsqSgPFlg8HyZAP45/ToJzwrcU7t+LY/mF4upNyctbRIQXQ9d
OD9Q4PyObDEJV4h6k6VpT0crJhCEhO0qPvVluAC8OVEZtY7aQLPtPOwpC5uqGwvO
/RaJE7Va0HzJfxxcKZWG8VmwS5vJOVu4E3nX2tpBThN8vqJqz4pAQAzKPSGKHXJe
Z2dVMh+GE+oXVtnLeNlm4wMPj7VO6c5cWOuOh884HaNqCUobjyUqlnOCqnT3rnwT
TduizJ2k7vWsHa28aseUTPDWbednvmlVOLZH3TR6/c0zqpmScyI7caGUm/k1892/
akf89D7AObsvoRWyu3RobvEeDutEyEZwbfhMJb2JggHi0aENQu0A2LitTef0RpEx
wW9qXDBNAHaiPeY5On4z9K+lx9UTcQVYQtQ8sT14oIgxPumB0WnRUauNZs6KiJzt
yAzmUWf3LsB7TW0ajbWQXkYyrmpexiWL2lRXl0TVvIj/I7/W8YS0+wSejlyiJwCU
HuTegygk9H6dPRtVlhzXphv+r11GhkajYn1ZXGU1f4+Scaez/aoYeaXgM4YiPlJb
CCdn1/wktD0af+Vfv4U0/0jS9WaB8Iy2duQTXpGwrtFWzBqw2jRa/Z/Sh7ZyaJRF
SUuEmDVJUDdzuIX+doHARUnyWAc301tyRYPjNFg9zbJIHbRsq/+rBnkr5orE9ex0
lzlasnsXwFMdwvV7HMdiqEpfz0m0XDvdjp0ztXyDMNEZPtNJshZCGVV8gluXyiHX
g/9mUKuDn0igJ6zi5R/UPLWcdAAHUfpNArL6M/B8Bbz6PYRXZ6vS6XNiQU4I8QMt
SQkIYoykHrFn28C+W64plKhhRc47XbZrcWcpx/76yYI4PYXLS86eCi8SCVfc+7/b
jZiM6TlNF/hEc73t3uVqoJmr+UIFL5j77clEVO34FC4QzhCyKEAFaOYtMLpLTpNh
qNOyLVLcBqzdvOAGM9NcfBgWlAQQzZF/ae+QU8knTKYOy6oogKVmvml7hVnkwZPk
cNp/nKY4jrcvRIZQvt77ET+1UP/Vs34urpxlF1eaLwu7kpdFros3gEtyN8TaDCK/
WDK6NzljV1KAJKgy7jzM+icScWiznIRmkQ+Uz8m4JCIWXpITDBB38PxVLRQ+HPT3
osGSGPbragq1L4dV2jfWzzosg5/oH/88Aj7gEKIJZOa/GeIXzgX/sSWuXR5viiEz
ioCDY0G8EflU8XXlUsilbygFoAR4ofPPMN7kEQLIcyROKMC0AwADjkkKoqbA1r6L
ldt1qMwip8+1bvHHhxbBQDKUh6OIlgTWLlWw8SER8VTemYHD3XfO2FN5DIbmGpaO
bAoGr3hvteOxa5eOJta4XVvyYM6DeNP+ZUAUZqeXZf9IrQi6z9VRWc9+vbp0NUjm
oeB6tKViqgtZ+zEpjWY7y/v0n/QPoui3t4n4AUamE6j/wEPu32mR9JVonDdIaqrD
QYG/F1+9TUEFVUw9TP+Pa8z14Wg1sQRmf2Y/qqKC9V37mV4OSVe1IRVG4BB78PC2
ZeKEmygcbsDpftujqMbaeAVwuMUmYSGshGiDgDiBxj2i/R+UE9y2OIGDbB0c+4bs
3WkZHt4gnNgSUKQSRr6Q0Xt4DOJvFHdfQVy+Pw5B7my4iGR7cGxW8RkNY+DqKKvn
D6Av4R+XSapXKrKiiZWTPdgvHNpGgPC5afOXTx1dN/pKISNZ/e7Z4Ajdkdy/XWiw
rk+WXGMuuIClEiyEuFrwHQbbwLDpBbhVhA9f3HlDvk0rlukdGQ3D5MKEDrzu261f
CpdGL0QDjtZ5YiyMQkilgtTAiejjxwNy9Omkre5hXHsGLt2x9zi2w+u4PkTG16sm
OO6uJTdYzjSH5mQ2x5IchIzG9UioXRYdzR4Fuk7pI2yWeoWbHDiQxS3dBRn/BOYK
wio9EVFG2ZsnHpjRiPG/nhTOWsQHdBGqSzW38C2QH+DQ6ukhgQeXQugnFFKq/ZkK
6Lu6ModRq82HEEtQnn+zutJeIR88UXbT5MFbSWpcOSbXtCMeBoJ3aTPlS70jDNDu
8SeE37fBMzYMS8LTVcs8iywx/yb9zapmrJZT0ODFLCbyDGHmJqO+k5ZdIomB280X
QcYERb+YmXohQjgCFWYT0elckY/ErubncF6V0wyOkw+McjGrjtn9oq+jdkhM0rx6
k1JXMrl+jwKtsFz2I8AIaQQW3W8Ur5VQlnPWEzwsf8QSXcQyc85rwSWAAk7nFBR2
y06W/Q3WmOOrG6CfAqy1I0JeUwoZK/Vu6egrBA6YtlXi+8YwCAAf8NnaQ4cm3p11
jX9uChbsd/v40xFtYck8zE1KCiwzG2zk/UcELyimzY36EXcrdbrujIuzCO3U3URQ
Jr4KtH+sZb/Yc3AdJZ3D6MOgeOmuY4pIlw8ZLJm3fPEf4S+mjtTSOT33BBql1ANK
7BZeVVKDghO61PafvS5Pk3JYY23RvdUc2J8reLkbvvVzaH6Kk2XqOKMqYE2f3dPe
068Sdk7/mZZ3IjxVTu15i3B1vkHzWjeCvNppFSxWd7lIHsIi6g8IpMtxD2V4eAYQ
SHwn9ARvoPzjniBQJUsXU2B793ODieXDwN/wiyQMmX7MzSlySngFFa+zJqCKQqUv
1YP4t+MuycDKziCiGbgYoQ0x5JIQmB7Wp0WsYTm2bnU2u3HKeS3XWcAN6F3zgkF9
uKcz4qgJQRSVCPJjZnaJmnBsB1FqiLGAdLjFwriSRDz+lPFrDGG4VwPjuqT7XOGC
vUsWo+BLxRgtRSvVCRtrauv6MrYsha/m5XuHKWGflPLJdwmnRHtoN+Lea0uHkMWu
HI7u/Asd9VzUufVgpZWTK2U5Eouz+d8ra9X/YZFxKO3s19BiQ9BDEX3yFIS1UXO2
VVY2dBrTArtIYjb01dQPNp0STPpOBY5grJMvPaZQEvdiyIsCj2ugy8Y2vDlEfWic
jDXckbwwTdrk6+CDTyBX+u1rXR+EpGGwrVffPlYrMSbYTKvNTxRdxRIFnMTHpcZP
DOIhtB8CsLxsieaBi+3wapWLDGpol1gNWpNWnflOdE2jvIvNRXDgEOULP1e3x6oL
SR2nU0d2GFraebxfQ8f2d1L1YU0emet5E3x0iNakIWY3bRo1kulCZ925nxwKpAsR
duCCX8SKp1sTzfz77y3hr0t3jWPNbO1OIGKNk9xVVCPnVEp8+BNQx9/Pnie/+1B7
4PqSCdph+3svgobD6m/OqfmVJkpkq/2YuQ/gQVjKRiHdyWSCrfDT8BIF7m/ctqte
gKvWgF1velsp15JTnWk+19dxwaZlwno2nmXEaj1uekcfALtRdeZWXPOSvnRDTDMk
ry8WpqVcM+tcVuEOQkZxNC8mawm0/p9znc4iaZQxkY4/0P8of8QRXDXnlnqr60Ls
OdRFiJVo4+NWGjHlvo39w9uZcZPx3Prr4Tv2v2p6SSLDhedEnoC+AgJM3gxVaz4X
iMxcN0SQqj0V36uCy86V7n8pSy9jZR6LUw/uT6lJEmi/Vag9kVcK3HbOpBVhvdCZ
AMJCBa0siKLC14rZd2tWR6k6Gh9wdXX0MJxT8uS+6BHEe42/guSR2/966ZmM+fyo
7YjzGnSiaQONvuQjhnFXMvd6BrwB4ol9oytkuFFe3C7+NztuwLvzlv51tprv0/lI
InhREhp+2zOWDQs6vGf86vkvKgzgBRNmSq9OFCMFwar9oFagSAsSrWHQ2jOpzG7s
u+gMT2g4Pe7ghFrb7fL5Z/IkgMGY08Q+KCzppmtefxeV2ROrcYI4TrrY6wpcdf8J
SIX3wpFLloRj6NIY8IlQNK4ZdKoWsN3qzj6riXFhMfip3BWLenvXEVR6bYh3gHV2
6pS7r8IhO5dou1ERnTz+Z6UjAGcfhmJu1NL/Tt8kwjed4Y4vwm+vrbhVfpZSJx1f
Tw2NBe9UUq3/Wv/EGIg4xcjkrNxvoLQ7UOWrr7QnrHx8ShBb+HQsMT+lecFzD9O+
bKQAO9NJfMOMpz0mejLBE2j+EX4U7ZBDzG9wufDd4JAqXQf109EYTDebgDMzdACe
YolpXshPMFgSy/e+x18FE1xLppkoqmUaYfWOcvf7XVbx8nHX93Oj5Q6pPqrwi9gT
hAK/JqxvUnUUjgKIVnHUZu3VS4vdXqBZk9wbC/qvOUb6yt42cCnJwsGcIZ10+NTq
u1sNsIfVBhj6qgfaZqG57d+vGbdaG30zIHHWmO6dKGtbAtBFESAE3Q43dL4kzefV
nLmYlm1WZZL5jR4L+qXb7LSeYBFEb8CnmK3wOZGJnVR4Zv0pyvn2bLgldAhwQcnZ
8tehuPKYe9virNPS5QTMquKe3w4vhmhOf+JnqlBAm2F6PNL7Iu854EJD2D5jX6aQ
xjVT28HiCayvQ9mXx/2WYdsF+i4qJ9YbxejPJ7wL3X1TPSF7+MwQxjBsF+1FQZnd
X799OH6I4b8/O8qHiZ2GTA6k+KrbcnG4s0k3lrLa6vCvaQvlhkaOpRj0CBZZmS3m
lYygcnArftPcUGiTR7TFtD3B22wF+6JUb5m84aCefZIo/c0CqPRCpU1V0Jm6lN3n
apwuDufeY7fUDPEOsk8slIkFn4uIUfydIlgcDo+fqWYDUZJKDPqCbnsnid2IShe8
pub1/PHgRCX3hNbPO+InwBhWqWEsE2v9Zp82LpsvBDv347NMUFZmTaHazBO/3zBg
EkhfR2R6uwaBpfSUfTgfHB8peCBG6lmXk4kMHUU87KDdHvfhhifkNHLXFG+RQrWJ
eyD6MHYqG2tPNuSIFmrYtuZmFWLizdNh4iQqZv3GcUfFaQ3NNWhe3vaWZPMHVpsO
U26C5HeU0IY5ZIDxZ7EnJiC/IS05VjVNfLruxIV1pxoJUd2YPgE/WtkYUkIwVhI8
uCJM0DFSLiHLh5H7xqI9HQHMrQV/erMDsK2ukik4AzGz84q0+Nj8LwRHZMU4JYHP
eKK4WnNh1jM4HdUyXNju3pPEtrN1Fa4UPtwPzThyGSFNutdl35Qun4+5k75UMDTH
4HYDYGhnyLHSWBOqdrDlX3HpnlTA9j2d5hwIHiVR7V06OmKL87hI7CzOdaHY6ijT
KSqp2Wxm1H9SuvgBjtHvK23aCVgKOSl7nc1N1KhgartmD4nj+QFhuFZt9lapzXAd
XpyP/GOSoU/9j6kToEzZ4xTow33VPHBr64iUatHyvDwm/mEL9wCulFajEzL839fO
HKOOdVBWNol2cTlgEXQ5Gp5jIjndoD54eJORYlLlEFgZjvet/Y7wZvv/7RoOtIKA
A7smEBht0X7Ki7KTZ+ta5DTe7Wr99n4HbdVPa+c8gant8VqzbkEcfWlojQxqHnrH
23f1DJf4+KRTQAM5N20970EFcsdJzcdd9ufpNIMuIm2yxFJ00Y/sr+80WVPTbw1t
qZoY3aThrwb8wDdopAqGNX3b2VliUF3V9Kh4HgkwCJQqkOmgId32PUE7XflNjobn
bETsdMhKQzUGhqZN2mtq8KXUbFAfeGIvDezj+orgmBI1UzoxlCs4avH1J5To9db5
SllG4+8LZCeqIQKjYyMpYmSrS8YnhzcIRuFN+BY4gtiD7INVCaBgVjLTNGYdqVJZ
t4nffUPmhMHeDCvdcNuBj+a3xzMynVEH4jQbsRkCOgyVKk6rqFgMNoA/aBN/6k96
byvpw4T/cZa2nRe/UiPrTHex3pbM89uD3lLkczSXjsrfzC3QQ9jI/71W+OUR809k
jFRMsVTtSZfIM4Zj7Lb4YNVxvA4GCduCu+uH03MECnL0QWv4/FJCj2SQNVLa2kux
ERe32u6NlAfi2v8fzuFK1z7x9qYjkFDm2Yl4ptRELZsdGjirdDM9EWlNUJzjy6GT
IDbb/o9tTrFX12uFtawvC/qnK8uFyvkMBOo3t7oZIw/0Ri/V4GWM4rfjFbGRZqGs
m2gX9b9z7vpZB7QQUSz44MY0n02wOeXVRh2/RyIwQqcB+/aAw9ex/xm/CkLYWpME
m7a0VOnearQP0vomGB7BHaX2LQ4dnW/cove2y6uZ+2Fwb5j8GQvzOL5MOqnmalpR
rfZe06Hbmtuqc4kOpKZCggldW5tXlm5zz1GeQzAZ0Z/nIKxKxp8iN+ZXf5cAqnAB
Gzj2gxnDquq8DoCYpIMX1EzYchFE0vgDrlsN7h+QnPtmx4eGw0Gd2mD0SVMhzSXH
9fKXp7da5kscEQIEE7gCfwDsV2lEyq26DaI62+tAoXhRNSlmb+ZVeEo2/Nzi+wtT
jihvY/Z3f9rLrFGfuoGlhBe2D1vlmLZyLrdkSxc725Y6JyF1wohuW3YwbQFEYP4v
GzLH0C2wZP/OXiKK0nKZH0h5mdi7Jx+MkFmY/nQIrGz94/8MHSE7h6HoAJX8Ma/F
jbiq3xsMg53KUFxMtC9Kebsgv4rQf8bKu0rthxzuaerOt9Eb6sOfXDwkjFFbEJgV
+ZgZ9DccHh5NgUPtlDDjAKD3CoW+227if3ihn7xk5j+w3xNN/ClJuQ62miSy+FI+
Kag2Hx2UHntm1vxS+DMUKWUgLB5MvxKqrRxq/HQKp1fvK/vpJxJR9sYb4J+9jtPf
zvY4ib5NhqQfQ3D5bouwFzazY5I2iFh9DXVvJBULWWwoFrs5+0sxsJTIgielUUat
zfCuzu0btsAQ448f8ofSOBPV6Ijnjm/Kk5GH9QdmYrSnOjBVwzisfvX5GYaDW29Q
thqTAKFZ6kAyp2k7GXlsFefKiz8yLz0dc9h1SRMpn6AtjrIs76okLpXeSanjMbAr
sxquDMqzv7VVywwe13Vh8UJSv5/sfWydON/lMsCMJ/WpC1vCgL1ay2mSrXbyaCr2
BA8/NzZATqNwLIHYT5aCJAEcplaxFHuIX+MyDZsBtYVdnSnhGEJeEWv9aXRxkg4C
HiGWtjqouhmYcFF5/WfnavwocnmQZjiggPvHdwfEOloPxv2WWLsUz3ConTHn7Wt+
qO+4LSJ3mPluj3B9zcpLhFMCeI52hoHKeR8GC/uLNoxWj/wTBGNfmb5hYKViMrO4
4oHcU3BjRb5CYxTfaJxtY+7i5Frfr6F7kmGl6FcsomiZyj0NNMVJPp2EK2qGH7V6
pn0lHhjyULZPkgohCvDJqzRncY2arNzsHbomvHjPk87wQn7STYy1LGekWvG7dltp
4+UJsbOQcqgVSb4Wn3KROWabVKqZjIdywe+0f7J4r7SdmUjXcYnLFOlM3xYwl0kJ
T3sNiWgvxoXm5GlNDz6zCpb2AlxVkMqnddbw9eUC7UL7Eog/BAwBmqhdyfEXaxy5
OjOWmA+0BE87M46B88qmNA8phPoQZO4GXubkGE/k4R/KkM2SeRfH6kLfk0wSZpt1
dpyGD8LelGWslucbJfQUKH+wzgc6mFHIPs3VW9QUhvcQGfg7MQzEXqctu2riUPy/
0RE3xeeMnZ3JrFKOnNYBRQBEc5muxReNszBHm6g6szm/Eslw7Luk/vBtz/wqXqTO
WMeEdCqeCA5GtuzKhPHmwAJbuYYqnTn9T8JeaXh6osvQUI0qxbmFy3uVLl55HXVG
/Hy4xQqI0Cw84NznLSySgnuShGOYLHe+LwFmSY7pq88pnGM7bMOy+W8TlFTe0or3
+MPfAUH3Nu79XWtWcXYHm3s/s7xmDOW58Yd1GylZQEZAGEl0P+Kd6Zvs5lhUPacK
SqGuS42BQkFk83rMkPs6BWiNUeJGOxloIY/L8bTQiEtqfISIoOLbgKseIE9iDB/W
douNY2DkGeIZyzXcrg9eWFyFAB46+WdI2GcTZf4WHE6wXbeI6JIevPvrZo9oogTe
oybvqDcIFJUj5Utd3XARPl3oP36RuoK+2s+Jo4qDd+XLr/3b6H/qfMipsIk9qCac
ALDLRQ2AR1UFkazDjWp5V0YMiE9gFaFnRJD4Lko56saXGaHI2k9aDq/R8VEmIuSm
tLauqyEJyZUrfUtGv/dCntnOkmgN0zkJpw30OIBNV+x2RJXeLPHUuQaSROk28Opl
QdY0cpqxM2IWFTKrjWzsrfOPTHnIXGAM1py18Ke4qVfSEyaByP7dAl9P46kUTKdQ
gDfy219Uop8nhgRmyNGeLisu41M3dwqswhSeM4c4T6JAWxReWI5u6Wq9K3afBsD+
jwImYf0El2+Ml/VE3m6fuGw5Z7lmokfrc8GE8/3LZNI59b19J5o0Cq4sOfutTjeI
AeMVErhXTW40RdBkAsovefvTY9ndDRhgXodsYleLIhF1eVfwHJckDI1+TgKQrDEH
zqTz3h+c9+6/5ClD726HrtWlHOdEZ9ASsaKrQl46xqRkMDwedGOyFTTIle/7xaKI
GMJGCX5fP8sQ3gL5HXOYpvRJr0q5k8exjBXesQiwqlEygJZLOhRPWvh0bViCyMgE
JFJhpX6GBeS+pLKrYR9LWeiFrMyNGYjVbNsxwIcciUsYXC67ImWyfU2XVIIDVNVk
twuBqMBBfcBFXdOybwttcXbH3Rc639X/Nk1vyxnZ/xRva32b3W086FS1vtBwsX2H
orfbWETderYb1cGBj6csW/KXvHEobG6PEjv0+jyr4F2oCR/GdwqyseMRGoWJRi9W
Q+76h6iDQwweZRW6UgRlH+ZGywNGTaXXIaKBcbAxCQvwYqEcTtOT/88+4phEh5PV
9gemc3wP4yAlbKThg4QXyXSwzr9+Wlu/qGN/wIvIhJwPUR6Ud4Wgd/7Kyo9uFQbB
he07DcheAsLeo1gVQLUHpaTwSAcqOHp6sxjR6bmP3KM2Ed7eI/9UKMYr9H+zvBib
kXkVxMRBa1LNxaQCfxFlV6NTqjUY6WpWt3Po1Xw3C0z6Kd3zjWPToH+GnE2c/P2V
Ne9o/047cJdGi8MqBP7XXShq1/5zZm/ZzEdlDDuifuzr3vOvJyyZ+RhPHgbEjgTR
GzB29eosx3h7oRTXziNEyFO7K4WMw80Uxe54DRfhAp5HYKpSF6oY5vOOOSWgxtMU
ugCGKteeNAlHVbDXGAvIL2x+eaTbUi3FBt0gdobzhzU2jQr4UUVNrbmR/I3xWgOb
hMZtNHRC1ZjQMASJIj98/nb+rM9clmLryiOY0NVkHuKochxUB1TfVO6FygIUUtMN
1wE2+ByHeKwkmbi8dTFDDqr71ufHFIWSKYIHGxUCL04PT7TmQ0qynyM+nm4+p3O3
Qb65bErfA7FXnRGbUaqd4AsGb+P0CkpE5etgs+4pinfyf/w2eSOgWpJ9esxwUgxa
oFjEIEVG4rgxqGFt4p1iombTEHXCuZsAUaXi7GKX/EgvL3q3G7LRvSPNUgQKcGMa
yHvtIXzD64UaNPZ9bGYG71g6tsiL952HLTF312QxTqXZC1FSfWzDMjHMX2CfshR/
42kPdZmefi6pySRQ9Y6MkFoqMU8dcikUM3D+2p5wGmvZZv54pwUEMF4s8NjMMtgH
Lc0gIXDyDqZjGJEg4RD2tUryQNgkxXyVzl96MIsWPf51VgA3ltaAA1i0k4w2y6JD
kLJf6Aq5Nvsj+pBZVx9jYugOtDt6ewnzkY8zqyM7xQPfSs8+PLk9c4vqy6/47QAY
6p6tibi6kTBtjBif1AZ63fl0h0MrXnYVa7FHBkJOU93FylgAMw/dev9kh/WO3aRn
nnMhSoXmm556qT928io3os+AFUw8BLi7dHkuwclkJjt2pbTEhgvk6BKb9llMlXQN
i3OwtCDMbjJVbrcs3hsx+WvNw1o6aFus0igddRZWYAAykokTvb18TS41RP+x1GL0
ArHqQlesI4MRbR+oTxBMXC+BHyhg2o/qgypDU+GpOkj92YRua/gXDXDzvH1fJHpL
s6y8dAt3dIbWLX8Nl12LBQIgFIh6Y6ebu67383QHW3c787fExyL0v+yFkEfEZtis
u3poV9Gh8Cjlg2SbHW/FhaRwvq0cqkviJFAiHD/6mVN1JEhZ+3UIB5+zaaH5jmb1
edYiKFV60OE8bNe3iNzbs/DCd7hq8G7FqmtwOWT0KSyJ2U4+R7n8XbGNS3FAj3Xo
5sCE/CXSNoX+Jy6hpofThMGCGdkVCtQUCygHGtneb/SBa8l1tGnupS+WklTQA4RL
niRFt/L3uZ2+DvWs5+Q+0q+kE6hdoO3co6wFxCGpe5FAXrqYD+0MMxw8g4iDiLLO
aRgWm0DY2IKtpNfZsqxA+DVZBm6PSH8R8ix9uGA7glfoabr7sWy2qduDtNwgcIhF
mrOBkgdtjNr5ZKFcpdIXZy5TvcEbCikHWSbaOqc7rtGt1vyJojez0GYt+vMzK5Tb
iG8Qty/lqMB7uY/X4GruHDVcZh1c1ApZAoso9RVh9ihzeBwOqhOZA4AXAhjq+hJT
sgd3v+p+kiwasgeT4iOX0yDLeTm3PbvqQASpeyqGucF71nwZwy/dfQmqHL/T6ieb
INgroxeK3sjLLDGNLAOBc08BxOKFl+74Hy9DcxY6lUHAYSQZ0SwozxNaHZqtPC2Q
ePoj+KjkgWtaavD/LXoSaAM/Y4PTfUSNcG64TuDJ0eiBBZXVzapimnXMgIo5Vta0
Iio580l9t7EvpTB81w2bM8jLLICd7pVqyaD/BJJilYD4/waSIJ1maPlyn83BpcPP
JAmv8xPiSrp8qSMY/lbSyxY3D/wYYegJhC34uqHveO/3AVO6anVHAGTH8q7yFQdY
t+B7f1/TwhSEe4E4Mhtx2qnVFtlWO6b+1YPLqfPPgDuhEj9f/7Oc1rXQ+CRydKV+
+nn6dDfl8I6M6uUusGyPVJZpmjKwMfpvFYdcugLJZzwZcfZWLl+HJK6ajG3L8Sxn
Hmd5TK17/UgCNv/h9bQwAu4RCGRL06bf8ZU/wz9KW2g+nZuuVgiUAyorpqhpLCpY
85krhohmCLCAtEoesBDtzExxOZHTSWNWEx/bFK6EXOoJ89rCLMF9XR4FU2sLybCw
cB6RFVdUyEPkdY8ZFlmKjzojKtV7ixJIBVTbZLbf1oX8K0Z/b4u8IcB8e/4tCFez
yTbHyknkgLKsyAt9h1Ptlx41sTHd/gWqhkHGgVUoI76ZnK0JhxvysHGpAlS4Ow7Y
FZCbaGVVdKSU/9+Wx1Z7S0GDfgUuhClV0v84QY0TGIiIjAW86AnJZcJ0chCZFmee
eNCqC2e3bfjplSM6kG2BrtCHHXsvVGDFlnz5uvwfU6NP+6+yNc9ortCYCQhDTIdQ
MGmLfMjVwCuaeJBy2fC8udYbB+ELyJ9BLNwSs8KtpXye6bxnkT+eKz9F4qKHpNdx
+Thz+sTLJY5DiHRoXCq7YmzUNH8YNMig3f9NkGuMB+OmZA8kLeaZoE5Aov70Qk0P
4fuVLEcSqBwVQw7ptXjZJzLwJmivHp1xee6rERCOf9qdFphyjYhzbf1xP4ffAL9t
lTaMVKASkyxr1GhK2HvsWoIzxRPrXZxNME34Ftr+W99lm5sCONiYBImw74sPy9Dv
Czr69D2uyqcG6gg0EPOyTXctATOahnx1JswhcLsBQV6Wj9eVovftKVuKX2/AH1jH
nZVSzbi0R7Vz5w6UL73QyRTfGzSD4/XRB/F++bZCOT7rZGQrlGzphHxt2madlt/2
O2YG7EWhVwptLamc+PyKdGexQhklDsypq4IL2O1SKY0MzJdsrZgZ9W6RgV6ud6g3
9qTDxBWrrIAQajdly7SLn3sWCiabYXOc5n5SvaP3N1tST+2Vvq7V7Xm8kNrWyf7o
L447XRY+thzU0typGTMQleWxLwvbiYJSN/6OrcnlSFbFuEYih/DteqIf8xT+HJed
fxwYh+wfKUPf8XaFr/tfrXr8/SCxssAcnbRQ15m0HuSFVpFwYyysm63AMoz51cQM
BS5PE1BN10xBgYF4fFRnE5zqxON/LGqjYIancCT0HJCg1ccFYjZYeT9x5Zj4GxvD
U1klf9SxRk9J0Ju5lbax7R6Gdl24Y4l+mqeSZOCHq0C1R2ua67CjLBruwqOSmJ3l
mOFnapMsomfri5Fase7/cifN2QmfqMO/BOOioBHPIZeGYpWz17iiiKcRSyfQljw6
o3R5mqY6ZEdMCV8+J/MhBvoWCSpK4QgqDdE7O3u9eg//CSa5wSe2JZZjlUq/Qo3S
oQsLcTSNesiZlwFTqWhyk7t4FUkD9NB+Y0P9BBh+p/9TqOVBBOivIpQQLoHOLZOw
5QHziMYylBSFZHSpvQZU7/hmZXl+tj738Eyiqlx7UkVDUpzOyHiIlWUcvceaXF7L
g9WUlzgqSwQY4TV6k2xkPuU9+Lufz1JV6L0Z0m1HYSW6dhGjT73iYXW1qsR2PSr9
gtgKi1v+tq/RqQVELwSQLG4Jf94VvY0rXCQ43EWEL1C5dw//2M+fXZxzqzbOHbWv
oE/ZjxRQqouMsJT4KAXbaw3PoE1BCeZr1c3bFmVGu64LsAcLRR6EnzcFzaBEqEfu
y0WcjMrpnxFganmu7D8E2yS4zIm1r+YNwqij1f1GfKmiPM4GMJz4tRHLC+fhh8RG
+Y6VnktXPSPJYOwd1T1AiJTwyxEefiu2zyBiB1/Yvl+jLgukMmuLJcpIg1jDxsWL
7HrxeHCpI5wG8lr39VSVQruPk8Zo4J7sBGafUu+qRZ81dhMdbGp11EAUSC9OhJje
/1rcy9DPCpL0UifMsUatjMMz8mkeUouwyTNeK4/w25dAZs56xH0o1tJs63gu+MTy
C1uKjOVNJzYXA1y4tsg56FVr+gCbFEHTsu0U7n7N2SGAhN0e13ajughb7uKrFoXS
BuulFEBAd6uUpwXDDQyJVy+e/k7sNeq5hRdXBcTkWv0AO9nOVnM62VCOi4OPwiGE
HrvcfY3vEnzCb3LruROhHluCQgEDDNUdvkb/48lFlqtPpmT9rZLst3YVK2d5lTw2
35rhDGowkqzPDvEdEm3uew2YD3UYDuo4E/VovJR3oBjxO3q5yo+a7QRjJaFhOfyh
Zu/7DbYpLPjYrfruF6vy701sf/oFJCAy3rk/FAowR9a9jThFcCTIjGSur45H2BxW
7MXpAzqYGXZ/5v3+9kbg4AQEc2SihEtuK9cFK/SuY5qdVKsUh8Y0vTwn+mkFLMC8
3YzMMgFLWPZgsDK9hPNkLCfSrVkHmR0gI86reQg/1A8Ev1ikT6uXyjnlgbse4Qd7
AinwIC6CODkZPmYU9eMuS1Lf6croOTVz9+cXNiQsIrJ9YVas22FKTYOGEejBYn3K
E9IKBLhf8deEDmrJrp7aGzylSu4I5okkGfYquoJOSNPls+BbZqxgDsCPlhI86Eym
wnnf+TT9Jq3cu9SxkRxXzgMshN0K+sggeHLaj8jmiDr36QJ2tOSBIqlfIV+92BK9
R3Q0ytUJcymIs4hFbS5R50/F3VD35ROZmTropmBQM27/GUZzjAanjyNVxgK1hDpN
0fQ5iFUzBOmyvVAXwtIHqsf2OR28UytOFR5V1AMAgAMXaa0k0WA4oNifRrJEiS02
bdRLvc3wmIBgEPqSV4O5nW6PNaVKIFJkinmN/C6KkyGaXkRyIewi/0bMRjnw9odu
KZeZdYuvSjK9BNb88yh/YpKLvyqfLaSDvGmfUNdtbikikhE833J1hSgw/fq0w14n
wMZCg/VCkrdsmsjw6zTrpTIdhbTvdwSEdY1Jg/XNk5V+N7u4NiA8ONlKpUPYlekJ
wjVbvuVJmhb3hf7C58gTWWCxm1FPBRDiSa54wK2qcRFHihLD9nLC5eioEuoQpxUA
18mA5BC4lwpeCznQe2gGnq28/xrsL7PO48rssJY2FWCGqOSRjlkPZAt90L1kZzg8
i+2JByclWtvX3xNAjkQ8b4Y34WkbUWzT1HbcCTBdV9ftv2kmcPjszoa7OX5BDkfd
teiRfOBZbpwyh5GGl27GRmac+r9fBD2RZhsBQky9ihTrIwuUhKRz3mNVG9/4uYgL
N0/9mPnv8lU4mPpfSgLmP1psGDPLz49O864Mq3zMRegU7Z78Rjx4IGPN85Yuc/rI
z6PWLj6C2SZcZQ/X5esCS8zd20XhA8GPRHesiBLH2HJqr4kDYRKK8882MO1u9p6q
4i8UlRdReKrqR68ZffDVJsL3ZeNTrS2pqFYWiGAFSFMD1YKudpPeWkdERJm1ZmQe
daZu6pxKa0/1eqFzTigmu3EDBoZs+kIO+jRJdtK/vqC3sk22EnZE2M4fJ3PDSL6s
9IrNFyoKqvZbe2rTGAbeTqZu6Arb6W5xpHcoBjmbn5ZCdiAIZbfebHwMZz/GU0OW
9tzc/sZbEZTFh6F6kD+jmzIT28/2awat/FFW2B/1cgijqDyxc8hXBCqMFb77X5+W
IvmXlPnTAqqCT2ZO0PIZxYNCBKEUg3JMpuxNPTwgUiXxOJhRjrw68SJCjjFuXCLD
E7/9Hi6MHjTWjPkH1ZQpxus5UHCLSusYM6EEBMJc6iRsleevHBE+eW9Bld6qy5u+
nxLDTF0CVZ3MGZCp65hakjNt87b4EwYKm0Kpn9KE7qellkgNnhP2kcIxZOSdbBQX
Y92b5XNib94PEjeuD0s1vYBlJ3X9I+Ou0ibBNXZQv4tATMPWtT4je8vx4im2nYbE
pxuo98KNNQA6eEJDFDByV8HoIHB02racE6LGYuD8ORQ2H3ZylwbcB2UFGVhlWaZj
g/gVp+F0d32QaUtUnqG8fWWHLfC5jxYBrhUSRPb3yj8goJOLuYXV5Tl85AmmW2Ej
RZaBQbSwY3DE7KIw4cQWrroPziXO190q+S7NuJhz+N2MMz671DVgWef8RMq7Jg/x
gP8fW4FQF/AqwZd94p5iWr+Qrh5JhTESnV8hqrvNJyZrIffxNcDd2o9E1D6vwW6S
ZqfpUsKp2vJ1svniL36exQOu70oZpTmTwDvbz+M55qXc/GW0/bxzGocVviHIYKrg
N/vlEXk9gM7VV2stlyXvlNrG0d+lOp/Id5VB1udp6wD9e+IyUO6nttCNdSTMl2wS
Bh3jVnMmO4yTHliI1Bn6g41r73tm2ALKKhYwJNlrYJMkXRHTnJ2bk4NW2KuLoQAX
URwgE7jqqrz8UXmmu4XQqNdB+4oo8IM6mkQvMDWZiKnZPqDeekHB2tYBqfNwkt//
5cZvfRwvrkcY1iFzsDmog3MOlhF1HAU7WL50ZCkXGzhSS2EetAIJkKb9uTqBvRdg
qo7cgK5r2/GpDQjO0hfwbMgB2X3sX3LXsBBoWeOTffBQfodd8sjSL0KNMNmkDbjK
UU1hpdCro5HJ6Pht9aazx/xDNlF//KsoBL1NCend7M1dwQxRn0lE3VBUQY0P1xli
Xky9Pn1ALbyz2rGx1I6kVBtQUSDv4Gv/CccZuxqdXyvXYpL8Tw8m8qw5ME2so73+
3hW06QZVfnTyJy/K9Vf198UFI0w2hJJVftY7vcbICcQ9hCNXxwAzJpM8Rp0VQDzV
OZA42QnKqbw8ZdlRLIu1g7vunOYvkDuYVS4BV3bA3u3duSkLBXKeTGkYsD0Ia+wE
i07/BSnqip1tLiPvCkUdHlFoJ/gUUo8xT7Rvnq65sPXq4mGlsJmggtzqHpPmGM1t
64M/eGSAMQNbcW1jTQ2FQrMbZIm547fOFhsnbbrN3wSZniV4RWbYoKWPk6xurGMr
OWW8iWBCYzlerMIUC10yEH+KB5rraeyaoXM4ekOlqwtnij8zq1jtX67ArXtSBXe7
l4BG6xIQUrAtn4X6cCNSYQhMliZQvk2vO51zAIJTblaXpymRCZipccV3yX8G+1m8
iO2Trgom0/sRXpW2wXzUUdonKnNn4UavEZkejpGC9VvVzfiu/S5f0N+WOq41oSPZ
eTqAaG2tWeqT4EcCw31IvkA7fcSSl3mGbfOWG3GdF68K3tiSeEFq0hGqO+9MyGCK
tlgFi4YI0qSEkRv9H5yW5fFTRcy6Mn6+R0V4TUI0LyUNPRPrh+SQRgmIiJebjhth
hB756N5h2zzSyi+HAnCMGZAlCdNx8JUvaklFiTfYktr5Dkf9IGqOiLR88UeeFA2g
spJcCR7HgPPgvffd+k78F9a8fT6bA5FlficBUgTIsLEIU1PHGnBb9KpIby8AtkQP
ZjgRzbNPYNVfsY9GLvEntZQkUgIjhva4UZ0eME6fZY2vA5xo4Nxz7OTn8JkOvRoN
yygGfEAUO7vjbfp7xzMSlT33PS2hJeoACE4fTp7a10JQZmalgDuJu91WZ68ncFkN
mEWMjQ5YXTFmPx5pXcSW5uPSB2IyqFefM877wLhywhEGQv6ZyJL7YeFfChyfh0hk
yMlG5bxtUCmH84Motuszaf+d7xDrRE/soa0ur9azke9MDSIe8XONE35XwOR+an3A
mll4DF28aX19D+YfjR0TUIcN8ESmol6QZGK7FYx2jES6KjY1gDAyDImXXrK4cZQj
vLzCIgKOmm6UKxdw/zBEDrosxTR4h/aSsMBxdHGkXWzZahW8mqwfQChLV8LYXiV3
Cn2USLEFyaD8c87wG0brjfDzXB5myMyKeMaKAUsFMMPXg9D7GuVXZACHcfS9r/zO
PVn40iqpPxumEQfDgeXAGN+zsP4pVHOwvV3BzIIlpBIquLEQistaBJ87T5Xi+IGy
/wKtz7IsEGKxjzi/PdyLDuVCP6/UN9MhRvqaBdu0M7F7zx7xHSLQqMbRuPNIzNr0
YdbfywwQ978QblUudhXnO0fZCl27SVXSASuuosy/75pgwssKWBwv6Y4ZBPxHWvUe
zSR+sIHJNzbLlb8ZycJcyBdii0AQ79Uvv43N/ZyK6g5Gi7odMkEuftHA/pwA/oK0
uVFnhYY4lp1OnhIRrJcYklVBvKSWZOFvxrgpj4aIhqFGN2NVw0HQ7u6SkHw8MoQq
hB3Siqhc+3LFfwpHoCQJtGjNlp6VILwRIqYfDYH5lXvveI8VKunYe2/P3bnu1ko3
luZlbTRVODh7WRvCwi585Ljp9cgboizHzYWRi+rvukk9auajPfXb/75B54ui1vp7
SNsAnzizuHWg3qyWy99M+HMY2pnkamktHUcPIlY5Np8E/+DcjqsTAaQKf30uIiUr
7bFL+HgwpqUF/Q5HkD/X7WOw083qPqT81S8s9FEVfNSHlsjRe9s2cEwxPkJqCQZs
7gnQH4XKHc7Rl+B/eOW2GeY6nqWl8aGOjUmj8h1xAkoQk8vTjCwgu9ZZYIuLWK05
cCqqbOTD4AhoNzLkKHRitqQPXQFJwxQR+cMCy7Hj6sFAfCiVhTV+vN8Q7AlXb6sc
w1JZxM5HRyYcLZYtGSPpgtJ+JlMqCTXPSUiKUExUO4qatzCGuZ8+cPYBN9m+S4Ig
m+AWvoOluOXTXHSyt1sGVd7c+pzlBUUhYJOeVI344sgjK7pOIDo7hKbjIDTHN9dv
eEfZB0kxT3Rl0QfWr4e6ND0dKkMoVZGehiEa7MXE6sgpYLY2UY1Jz0MjffhLWkHS
cS3xMEXXnz7yFqleCp0EF9fMhgBYRvfSwoZj4hG2J+w+Cz6ypGgpaiWh98se8KjI
PZYOmDZApxIxsPmHOiLB0woXpVLDFCQRy+TadbS6rr+AZlmkf7GcvyM10dKVUDYJ
tlWedPBAVaTfS3zmovwDePRK3/6FpdeoA6C9prYC9pjXz6VpELGVqHV7fnFXNMsg
rR2fYVR/8p/6zbshGAR1uiEReQxrTPqScfXlD5X3ve2y/rhUFwJnHfZc6JLEwcPz
ULjSe5H5KBOyo87L2tV11UT/0MGloTR2Z6DVnyG/WuBOa3pcAQGBYtovSrLLo0Wa
55GlUV4n20LBxdpqJhbT3nKjLZEjQc5WBxC21FIvXyLjdg66YqXJPteYBfqClQ/E
WqgTOceYi44bkuuwQmLJFO/LR0QZ00N/kLqvOdViA9+xsYkhVn4LEL7g8WaUyGBQ
n3eYZqC4ElGhWHr90gSKUwScSqq2cNjENYfXfb3sE8LlVnBby2U7JBiHIVzAZauP
uME3qnVQwJAA4UhFaF32U60Rs/syp4VLhntLvBC6MRM4bWv+vnyGG9KA3eCCPK5a
fpcmLBTRuHWoW7kjAxU/9M8MBhCIJFiicYsRKWIuZ7EAbOBGo/DQEGi8k3pCEwvh
0h+6XwVX+7NXZJxwisQvCVyf7av5EjKZt3LoBvykaRCAarFKAi67MwAmMm75UViF
Vts6OXtCLrcH9iLjncrKX78mCDnpvYJtZHvYOLqMd5qtb8uMu1CER+AZf+F4B0kN
HB1Nf1QW6wJHgmf++ZRlhWD3O6xCT2pdSqcKv9QdlFaQx7iGvqRy1GwMOQWIElM2
JG9JepGqrqJyb7xFvwQw+pLrGLELoOiOOXpEaYbf1FV546iHfu5bDt8quj0c2Z50
QJyRzcbF/zPfSHQlYTB85b7/lA10g6qNBfHIcKEmxVG3j7FeEhsOJphV0G9uQkO+
zsVRP9ijZ4ws/z7gyY/emN63cv1JqnUNggCf7Au8su7cTwHO4ljY+/ZcdcSuTEz2
V5OQ+SfVCicTQ7KzL0ZHgKeMgWoOvMfYhxTuOhj8lJdKwQ0YiqzcEOnVWesZCM1w
iHuPwn2FjQcnl73T+Rj3V0CoYmW7tGy3XspX7WkU+kdUdNqW09lFv6K1ByYEBy1x
IIILAbeoStSRip2H4oAxFO0CdGcyJcVyIOCRSbd8eNQ7+YzFBmdJlMK4KwlKncJi
amGohc+4zN57ARhQ93NMmG0PW0GjsF/fptY1d00YOqAN+blxFiiqJihpCoeaFKGX
oqmwPSAVxNlYYZPDfwa/21GcZEDSzG/ZXih/iHy3dRjaemhEONjv73Hime1D1icL
6nomSepdGE88x9vMotd42AbMdVljEXuAlzZtvUbFiTKu4wp4lDmamUYfS97+Zw2k
+ZOo0sUikgOAc+hbDmqA8TY97mKt2xJmFvTow/60YeqyziNRZ56pdtBg1KEjc7Bi
/QOUpww0QkAPkx2un8IrDb22W0nd5iqscyfFzZ3oyT53Da0NaW217tFt7YKnULRP
cYIwJaaeaSStseA8JXViyHEqCj3xAFARbaveMfCIusqOLK/37c2d603L5vGbsHxl
hNpRMGOX5Opk+d+gFFzDWmuz/2ASSsec+BWk5lB4tENRpKcqzut+kpEzcFFLklJ4
jXg/GqazBv+b6APYvTNpyNwQWfeYRwKEnhx1RDs8W9wCGeaj4RnthbG95ACFtNDZ
2KmnVI5NsXilrpswhFRY3Um4AvAs9Vz2A4iRXl5jnfLjVpu8zItmcS89c0K39fqK
R9WxDOc+MYdX+dInp5lyjAey7mMqFAMG3rxOAR0TTDuMxZSbPv3umZ/PKScc/QTl
rAZjpQJ2xsvxA9tG3Z9Y1Zk0QiQtQyVESm9ZcN2KucAmY6e/1bU0e6I6ZeohDsvl
kK+yZh9YNcy21VCqS4vpVcJGYI/QbAEWzQlxgExyxq0qw8B3WNsj6+QZyJQ6KYDn
uSPDVojTXxRtTyOCP4qVTaKPTzIvmoY1fs5f5AupHg7bL40e1rc0UaRnI0p8b1VG
YJAEky21w+I+mb65SkZcxwKWBLnGoo6FMZ4CQRlboNkT7IjuoszmZwp5HfGnHHI8
5UvD2SWtzDmEDABftrGldmnSqB151IhhmdivXP8Zgf5CEnOMS/vrdzzLFVyTa1Dq
N+ojcuBlahBRVBZg2bntLmiR5otXYtWT6KngCXdJApWXThdAOxHaDnddMupsGKfS
6uATvGZCaqWRJmWB6Vwl7ousrcD9n6xwjaCryxEggSFanmbnzORlwgF+ZrQtC/vb
htBWYJvfCfviMSzPVF/UYhd2HqxS0STW9Y/fbvh28b8JyT4I/4KKGqn40nLqD3jQ
w1pWMTfadIss0ga4s9jL9ZEvC+YRBbJ9Nj9OQVpi8UTeW68qhwglYy5iuHbIuy5f
GuScLVbE8Hte+IKZo8zvAU3FIoa4RvcpnEzXKKIWsRta2m29q0JHT1J0jt9ptiLC
gyVxXQBBYfuvGLMByXHInDN9/WiPf2FJz/WvxEh6+qUul/HWIf8tp22GA88SagZh
ZyskhoUAVh62A/bhm2hq7+DaYLl4rPIt2nbuHFqIN9sbIG5ijcMRYVblUTKDNHS0
xtBd63cWnzBzXhUFkGjfpz2b96KeR5C7m3maazRA5sWjYMMa4JnxjdbLR6lO8GlI
WJXDHiX5TfNKyG1NCCCG7L+Mz2aZ4fy2zJ0f5v0nS5bTPJRdfmJPHnFgGx4ZgBJ4
7XEnpGR9lfhRTfgh4xviopHNNUHvd8yy4pbeW7F/ANZ1/jEQ470kvDlT9ohY5H1a
jpAsNyFOqfMqG6wEPRqeS6WtUSvMXiSaa9HxoU5rtP1TFzZ2HJQs2mNIYV/IQhkH
4la4q/tkqy60ETjls/qhkN0sozPe3qzDWt9dMSX0Jjc6E+p3yeWjNAWm6/6VjMUG
rUeF2tVt6tyCc6YDMQV6CoMGkUIRsway5j9O7k+O16MIJ7G95NGfcF1gqbUThqvJ
WnCkFb/WAmy2h+9hBfZFjuxpf8202mDNLdFGZ+i70fO4MQPhmgp6DuI4WCjRLQjB
1+S4pd0zabUQmb1JG+PVwMamt3h3gxWa08HUocXVwNML7ZXSK0OAC/7YVv3GDez7
a5juYtJPLpyoBRqwZQboroLqKt45knbFRk3DHda3JhEXGP7MwhLa70BE0hPxiway
7TV5etDxaK3p0n5heB86hS62b3rd+c/Duv9ARp/rK+hitq/RufK+UVf5xvxIYmHa
kgqDk/n+MQXgZGlpW9QuPlSOlhBXPtBcpf1rsrf9Ndrqw8FxRTawYtrvwshqzwhY
A6CoKlS6QQLDC7wbISTGxOJL5hunB/atFN785vk7K82lIorJRHgttkz2jCWrlZ30
P58ahiSef1YMzEjklM1fjVMqUkiENX+aPK0HygIKJ6B0GIWfqosPs1miGHvkJoVO
Fe6v5TrHu0faDfrcTrH0HqUcmMKpiBjo+nn7F6hPLymysskzY9Ty+Ipss0SlXvld
JOFesCB0ZgOAe4IAP3PH6oa3I0QvFi7kjjA2J7mn56H8+oaWzu+ogr2AsNJxYIIv
jy5QaQ2sKdVC0uBui79TyUiNl7LbY1pXUuM5lwEFDIM7CTL856TkQVs7wi8i4ofn
cS8LqCCN8wFAXYurVJWWCnxeZ1VpJAEp2eSbvVPgkNiOfD4Wb2BVtOOQCHkhQpJN
6P8/38eAA7UigkBWvTr8jPUmqXn1oG7eyEIopI7ITgp9mGAH9zuE3BaiBkQb2DJL
dDgfcv/xMPQhkJn6yPt2LEDzGqLTdl2S2BIy7+pIvjN6JNKH+yoXKVDVrl89a5yt
zFVh2voMWcSbVg1tYBidFyQtDmOFiMiAspi3WXZfQAciOLXDE/li3E7Yq7NDs7uW
ZCCjeeD5X+LjqaXaJpoO5YMvfu+ivf6QPAQY4uwoT0Br9RsMxezGnL+bqVLkHBv+
3kJ4xdlOFntkVnJhNfNXYXD3ad/HxmpngtSDvHVPF2C/9IpgGRw6YXkrLqDB5bCM
ZtjjsKUYJ75p0DC2tTH08Zvp0yc2NNxrJ3qrHhVQ/ihxdEyotnKF118OpiNmoQaA
VlJViIMi5evvt9DYN07XkeRi0yLk48kY/tzWRxqvjh8J0hWEwk1LZ5R4+fky9tZK
s7IiWgzEeJi4M3xcOh5JUEb49rhIlyVxQNfgrQSlgqs9EKsYH1F9cK/TirDKcQJN
UEb9TiFb+IifJ5ZRseJuMu9XW6PCeJEHhl2C33lGxYAcQRrezfil2AHl+RK6Uius
pVDlrF9B3jjexniqYTH5ovCOmPTEVvTtdhgYc3m82z2Rr0qCC85wn4SMwLo8Rt1v
a4swWJFy1XR0NrnlwtIhI52wHwENvBiGWQgxoTDDfdbXlVYQE79+af5q/ZzXZeML
rb5D2X9KfQniPsvppXEXioIbAs8nyG8QFnWTkY5w6NE9ZuisEfviXSpUO/sTWQAJ
WBMvWIIN+13xPTkZMaSKwLf3uWdUQcN3BT3kvqaZCHRFiqtXXXh6vXW6FqBduWcL
dLhmNn0gyw9Y6DQi4sNIHbS2BG8qBeh6jECHw9KUHNifhri/P/EjX3DN+83/nIoC
a/U37xNiSt0b3t2aaiFXzUwhhsRk09kgyzId3XQW0dknW/R+6ll8OkgnLlkRFerI
ftdS4/4YLoDybSlxZYuyJE8ST6s6kzOE13O25YFMnvQEBAloKrtDZGeVx+5p6lLA
Fe1xcGNZTXZbIk7NaDlavJlihY08IxPP1o2m3qWfKi3LTgvPtxp683Gp61jlmOWM
LkOWQzRYCvxBklkpypRKY2yVccQ5AA5v20AAJpnb/Qn0UkccDx7yaip+0R+ro72u
hf5FkdrflrHJTG77fXfjV2jjoszrHg3PhbVuN///BOQUiE3PE1GiYjzzDfXDLgNN
FrQc2BnYooB8kNsxIc9P8bZ+WQqMIw8Kb1MikCdIfjwNpunnKSNIGcV0vngZ+/aL
ixWFTaUBrCObFKUaiXzUCog02OaVk4EUvhtr2uNVo/e9k5jBRJjAsnBHEAK798sM
K5FqW5DnSTetAzDcQnnnoIzBz37lVbX7Q/5AXeG4/6cDMl1XEvkIMXcZbjlf4hHT
YlLLdYdKKCAaL894uB9AEq6MB2IHY7B8mwGiUD6pS3wZhgiluQNl97K5uEdyJf5V
fA9FQnpoDyYoxo7rz4wg0ddQvZhx/McXgyZOzq3t11eblw6DoNsWAu1kBLojrEKj
0bPak+xny9Ne5avbE4E/5/0J4n8CsdeidQFohNBp9mnNWoj6LNArb6zQPdfx1UAE
ZUstYKieEn+AVb5ct9mz72ecIEQwZuXDbW9tBWqTQyiXO6GU8FxxmIG/6ZMwrF96
N3HPKCW6VOzeZaPDkJDT66AqvXI4nUM9n1YSjg6WMjGhbeQyABHugFHsX1xCAyWX
znNvcJ1ep1zPkuLgAycgUPX9p2OSVLF8hfzPjuX6ML7hhYxM0f9xpXklG77VP0o8
9i7riSLxY53HyvA55VbumMK9xoghNm7TzDkUlPAjCMvvo0gkdwehGBH9rOW3MupC
bpg+XarnxOo038SxyJ5KQ3UQthQUuihvL4hBrknI4Rk5QOQJZO4MrW15dYh4gi/F
z/sBH/z7a16sCztZXGOJ7k+OtU3jlSDLb5kMzY7GO18cf58kpdpR+tGXjoxreKyC
V1XzViCJ6R+R+9crsny5JaLpINL1DQsmVVSlRv/zds6ezGFFnWsQE8/XeS1FrBuO
L49xj+Nsv4pExGxE7Dr96HsCl0Gtc9a64deREUmVC+EnWFne9plvjWUFqa2XJg0f
R9GOT5zXESfJrynNjbYpYFLysK2Pozl0n4x3kSnVX4rZ1Xb/N8rU+FHVHZbmfh0M
ts+UZnDKUHOvk68AQh0TaucShg/WJllKBebt9W278nvqH/k0ucbvTJiSXqSD8Kya
zFUiRw5DPf3mYQLtzreSjRLycLribfi4yMIFdYAmw0Q3YdFsrk5UgxRvLuFHZcdY
ISAYGGpdZEIq77xbzKCy4VutadBAqCI53odP7U4mfAehtoEqpU44RV/dWL7n1z5Y
XbusxuOS0FZPJZ88jHZ5d1l7taGKbUfytz7Q9YVEMkna1mhHItQlsELgO8pGpsuE
1HnvOIJrcFO9mZTAns8x5a7nEWx/gv/CHfCbkyk3ksYqLrJW0KcBKC2mzlAV21ol
UNw0vlLlq5QYf21sUE1beBo+pMGTTCdi6zTH3sj7oPVIHFHaiVmg7ZoT+xQFChVK
ykXv8f3c75vm+x3KULBkvmo0eAavAnUDExm2fbS3OadBsWrDvrSfn1xEuZF4432H
Ax8OeYvOEaxfeX64ypv6YfH8J/nKJS70E1zAxg13cB9g2SDlmGnSwQ/V+RxoLpqJ
vk9RC7ABQPzMJHEYmW9v/FInFU3X+EhyC58mAJMwYxR5mWffCW7Hq/bdKIGXUpuM
dOWJnQaNMkSddYjy6KG5PkUHN2amFWolZaef4Rq+cu7YVz1m562dr/Jg8ORVwGRg
4FEQvzr9a85cjFaoZ6cIR8mXPgDiDWiriIZ899YdlzcRNXDJZ3w4uTxyzfrbo8cf
e7WcE0D/KuhHKiCWTu6pA/zCO0LzF3qkUl4OEZCmz5OeR2Mz+NkjOz603OnTtELe
D5EUvFRTZRD8bWRZKWFJeyGLfO8A+g71AHcpBQnT67AWOTtlEcnFcTtOrt3zPCym
VeP7O5DTyTNcoYEYAUwcTePm/lvSDeR4ta/pwaqAKY6sIP2gbHY1+x6PqcXX4ROo
5nT2YQBd7X8W5SUxhGLBB4LjtVxxhLVLWmq8GG5RZamgVnSMZcr0uYVEd0qAsOvQ
OxAwjuZv9IzutVwQEATXP6zM8IHuaFz0Hk39ea4ioGceD1WM6BxptsmTsbz1/IeT
hBV0PkQseBgPv1BuFE+iPXQv+rufYHPSBK+9qJxUXm/1e8bwCKtEqvsRkYh9m69d
n+z+aTHH9bdk1VeLDbETZAintymm0g+Mjj+++FCitOYaYru2/TfOgtsz9ql+qhUa
x4UiZMkxeBJcF1YpXyoFegu1gXCD27f0xbFT9NtVPKuu5PvBcbwjHhm5iENQVTep
ki9k53PY/j17GtoobABvdX6BqXSgfKuVkxuALfFk9JxwqbOoTcaE/n7ynAvK4JCG
ERRUKK8wpFrb4MrecYoz6ivUxc3NYa/XHBxHulLmhnBpaVLOOJONEIiGq9Z3dEWA
OD03C48PxEU22Fj3JzpqX8cXKC+xQ66kQ+ifrqQgydr+o5Nb1UD5f13bxtua05wU
na5KLkd/C8F0BQDmi0mbhhHcuwO03P2/fxMS8aSjIylNrNeboMBEZY4WxAWgWozy
mf5MFXfzO5sR9Xg8lMxUydhDBSKGuHCbSGtQXvnSfu7Kp6DHkzKW8aXbXkhUBcIL
unM/m/+lnx35PHn4TFDPTPxnSIAjIHQU2/y9QZtObFIjKIwB4xwtjuMhjAsbGT4y
FmUyFcXaE1R/GYXnnVR5JeQmQoqQbnXuVtDSEhyFHoed78LKm79otnTxKu7ru4DT
xLGpiFKQn5/X77MrHQS/ENETCJwtL9I7YIutTlSNFob6I0y1nW5nnaRLRAgAbOju
WDRPP7+tKBijkPOQ+H6mwGYRmAJ/yQEYNZZ26iP7e2+h/dWlH3QHijQGi1hWFRnS
fxVigictMG8ugaZvEiQvgBS/AlwQOqCpTjPzFGtXfy+jG4PlZBNu+iGHLh8cO0U4
2JCuB+K0uSmd05PVU6BbzTfPIrC0thrRcOxr9eg5CY7iPb4OZoTWoXCJ0hPQDKgw
nskCjml+O39UIOg69hpgPdntq50/oXuM/vog9UbQmjKq48/Ja64SVOQ3maWZ+Wf4
rvuTtFKnOfVIet0ckF3BfVSepjQJnvasBB0T13LJ6+DKvY2XiTBLUpARDbbfYmVK
gjiSoyulzstMUawFRhLrjlqp7QFUyxzCBBQiwwAee3UryskUK4gNAvRRm8/fikWP
LFqcJ6RSqANJvCdsGly5NH4hvo1yXEWAB5TZpnI0WUCt8oCfAMVrFnb1uoetcDwG
pgnlZDR8CYAFv1YU7O+IOjloTK9JZAi00MA+KCDHtmGIy54B3YeUB3z+gqNwA0OK
jGeTQBkQsVZydFGaL3tw5DoSxDucnMoxrkMR6OKxmaIEPLQpTyU8xTKR2ksOMxXd
PB8JBoJ5AqTZRjewHO0zKlc++JnQO89yF55hQ97TV1ZgtG2l9LNPdKXlvk5/qWsW
wkd+RNA/NSXlKqdVdaNwHmJWumrc8P+zkWx6i8o7zyCcddCsJbn+5TgeOEuHpErE
Qcnch2jgsSQPouTPA5o03x0JEN2Y9RFIdfD0lo5W/NjmGnYDXLlF7MMEGky/JLVd
xljxjwMaLGEtldsYkCXWPcDOe+2MQLFXzmK/mbnqChy0iNhBnh/OH0bUei2jT0CI
Ri527uxbh847Zyuy+oNxFNDixNE3aRVpHFJa2yxZeoKO1mdStBAEtIwM9FOR0kJL
l71K/o07ss3BS45sPT73N+oizlOBWTDaAWY9Bs8iHPxfuIPFgtZz6/pwapqOGq6b
1yEZ9POWvphW8he8IBYrAc5tiEg2WtZ7lpHLHQgz39QATMzA9u4MD0Ll00kWlpic
I3cULPp1jUjCQtdOiy2NVxqD3haiYb/hJ83BETDBOJksE+B1Jto2XPxoI4y5BzN0
Tr3CphIgEM/PyHopqg1p79AiXRVhQS4a10rHGV0gjmbI1Z+Sl/+CFAa1HLep2/eK
XLrUz48Q+O0ut8DHHOGKQJxWf7xoYsTZ8tUGyMSJw1ufX1371FyIw6D0WChNaGzP
EzpAgUwwEplmCp7gSKOfqMNFqEoFHwSbfgp4AKidsczKDbuNfgzdg0CY9aNLqcP6
45WzRC2jeK5w1bqOGxLgDZ7WJC/ZbTlPX3ASVWO8jn9dZQumIaf/iS/bSfXm3Al4
uCmaqm9XbZ2W640O2gSLnW92aQPypNipz/Wey1LB6lNaBBKk9Ppd0+46Z72uYxst
UpZFC935flf2aoW02u8O4gma4FaztSm4bZFVNeIGBTcHH45g7ePtM3vAWy2FnC5s
TykU0mLM0oyBZ9VuBPH22XDgAi28EdIZdyNLkhrb0rsO+W0nXPWOOsN9wbMfaZKb
gnNvMwHz2D+0KyYRQNFX1oWKNyPGW2wUilZ4jOuHbZfcyydgH9BMDzXBzPpNBVmb
DOh8Dh4HDojz6detodYyaPqSrGqMpzwNQE37PEnGWnyGly/szJow3nU4fwSMO92F
IETJUg6LF46UMaaxTFbLs5nRs7tAtJHICo87JtMDXS6FJM+lNVziAJRn9kT5XTaB
fLBrG/dcCzjIi7wM/l1NfxdmY4BJfsto6f70d/gb6bGoHnIEYNyCIA5bXqvUkEuJ
JYPHj40/7HiysFmq7L8KrJhWf/mCov1NxidDiHPOjdEmxVN+4jZFScyzMS+qFaPF
7Jws9zDxUg748t2gcSay2469NOsbSap8v5CHPb0Or53UHcGUiiD5nwkL7doralWl
TZXuzcqvVp+5ZDH3OJS7PSDmZCO+v8lcs4h5CAjE0DXhf5x90GztjIZGJrhI1Z6W
zvOkmQ8aOJbEm2YJ2HJhGkxEeJ3kEYYnfWNfeHhQlVeLYZkVqpPQMS715r210kGk
TXaJpC84SLih0jlBlTUhedZisnrCUwNx2CawRoBr5TmCNy/bgL0DZtKZBIdNNm9u
Gpd+XSofDRi/tpm7G1w+EdShFoyv9VZuJkZy0zr8mk7Ps56MnZn/oT3uKn25xOBt
zT4WqT6QkwAc/sL3mG2EagdcgWp97qcwbPuushpz4k88VZ8yjUicYRo9xE4yzECM
1a+SPlMomZ8CQAbZT97de/RyzoqIazVSKhoOChTWqBvsKP7mEXTePm2OUbrv6HsK
+RhumBqlDX+B7YTT8l0XpoCFeDSRuFXNwCxjdOxbjbkQIIcXiz9/0mngPk2LuW+T
Qx/nwCxpwafeDCIcUF8/hLLPAxfMKZjJYpwMr23sLXz3PB55FK5fE4zVRG/Gzj98
z2P2DcyWZwvUyWobJ6zyWNY2v1/+aMcrV7MKH+W7vpMtb732kiqbuDe72yj6z7Vw
1ki25mapsauMErDG/v9GRc88lzGieoHOMptwy5bqwNdOF0XFKSSnAs+Em5Vyjmx4
DIt3XiqRmlSlajDg486xJYMp8TSP5+GsId2WcrUTbSf+rEETs1r7wZtks1e/T2Hn
dPu2O7Z9RkmECqnfPcTuY42XlbrZa+W1BBiwvIKuEqfRCug3+4i5Tv+17lHjI7Ne
c6W91RhhvQAM8JRpvjW8JI58Yro7ramDEHf3YGWEWKdBnYyrJLKHQf+hPoQWeqNG
CR1x2QlJWpQYlHkQEO3v+MXe4M02tCxI9dvypIvLFCB3sLLxlqRduyracMx8vSDq
OtYZJR96su+wrtBRYVcZeRA/D5nK0wgdzBf6ENbvtL7FIzz4ux+UEINjFGQ7U7f5
9mqfb6fx9J7GVi5eekRY11242CfB501aYUvjSkNBguvlsaDDDbAaxVYhda4+Psv4
gyjOx/7DpyiM+1T+UD7T5ru/gWUOkPOBoA5Rhg5vYMbIPsutucn6+/KLY6dyKBEK
yABdQovz/8DdyoR02y2Pzv2whUfIkGEkaBhWJKHuMwXXSgrgnFiIqP4uLb+J20H9
cTh/FMwNLP2tqFyHqazRd37Ed4JlZKCoNf+uvDfkFCRzrLKuyd9rMCUb2MXG5s6j
PsPOx/B3zl3Y2W2LG2Pl8eQzI0k/jnCB9lcLgbTS24X/NbaAeEq35sMGttwHLd3w
xcsPhOXUGf3R20K+m9H6J+41YyI7OpC8v/MEKzZV3tFmVH0f4/5MTEehzRrPughb
GxEjIfu8y6LHnAfT6EI0N+yqXPhPU8eQJ09w3ps8SbhhHfftXmJC8OWArs+qxScu
v86VYzQ0gEWPrU/taeZ+LgznstiLDc07Humw+9xJXu8hIm9bDYeoSo6FBT0N5ipr
FXhmIWnY7HyULXegqhMyES4ka9hHq30LlYWja58KIGAgtxauJkUmzVWgguTa8cZ3
qOoV9rXRGgR30wCrFS7U95cideVUeG3ht3+mluWpuiK5XSofREY5ev5n6EFEUEUO
VKNGWrbo+rAvlQOwex9GSOKCQDzPNPS81V6R77Q+c/kvVXZdAF5EmoF0b8qR38pe
XcqGf+N7mne4crTkagu29OPDPZnEewAHJ0uN+8tBjMUq9fUdf7KyePQSNSrB6/FG
+MMv8WMx4vaI2Ppew9272Y0vkjVzOYy9Y66xqrRbHngnRhTurvZ56dJnOnDcx+gY
e0+KXi57vK++OaJt0hvu9x2gbfHrWc1qmTPb/BRtVNmQyIzp69qxTeP/qIwsCkXq
J2EY4M8yXvo20kCX33OfZecOhqgGQUcH0UQ/lNTON0JhOdiLCi3sXXGzKsU48Vpv
rofg3740AsUFv3LsCmfLAHfc7TuSEyrbYAe8SHj8KCIgWwynFSu+MbgVwdC/UnyK
O2Dy9jV1ScDR0QJSpfo0wp8/e+440IOtEs3WmXPCWmjJr7f2iiF83D8ia/F3djcp
ZzzGbZgoqCZ+k9Nyg8zW7HSVA5IUnj7hfMUmR8D7FL4UpMpeR2KiCnJlJD1zC88f
G380Ky7ZVUwdw/ILr4ZpDdVsBjVdh3l7any8Bfh/7be4q5sxgxMinYtG95HzHHYI
+M0NR9M32S1+J81jCy2WaxuuUOa/RXKZIcbjWzhkagcar5wiarlutl576Mjp59QJ
npmMetOGqbM893au5es4IwCNCHnGCZcavX3HefalLv1DdcwFkBvanElCiUBUsYSY
xUZnGlX6Oz7EQiyUy0SpEH6AugiNzMMA7jYyXitSwRchi0bznF6cg6nRyjsx/bos
UvxgqIxPZNsiQcFUdVIszuhYedbtpK0+S7QRrewQUOTYay9KcU+XuE1C+RVEqoBL
9FJoliv8ycHYX0TVB7QFDdUZbuC1KWOS82sGBamE8lio4OW2SY5/8O87fIu/bAuB
gkZXnI05pFIrFJuhBrpGc0GRrWwi9BjBgryIKMQbihMbR9+257zLIRiO/Q+5AR1R
BiaUVU77qQdhFYjRf0Q7Oga/uaB/+k374do5Y82739NUn6zqJ2EVVkOKmukuRQUx
sIvMLgBaBVjyY9a2CJKxHD8eDcd4A9ZlgNe/Xubslz1E6D8sZDR4W1g9XmuIYbzl
TS8CcDuKKh8Ya+4GJUdygUU6NCMuJilQtYPSJcIL7FN94Iy9pF5shwdIfE4cCAQz
InQUU32NXewY/ABqn28v1r1NrRkcaXHaF53kA0nAAUG6UwnSVLZknzPsFM4RN6lU
/4sY0KBQK0KH1CDXmJHac4+k0Gp5jGq/i2FRdpk12URIeqWXuPp4mxuRYnDOvNqe
+KT/D5LfSZWEiAUGTqd0t52MINnDpoGRIUT5x+a56Qm2Crs4RrjGYaJj5iXqw5l3
G+Ep28+G9cpMGPYMcqjWYQIH/7YYA8o7nx0f3YId38M9C+fA8ep/Q1GI4SqjJWvL
7U+1KugOYfImnogSmcnm3ba1IAfCTrg/2Kf4Z8vm8MWzVxQTJPar+Q/8CRcGZKIx
20beApnt9mZci/ajXGqOCifNFQCvBEbSQoo7ecB9HnX4KA5YzzNLehNNn3mXU6Dz
BRiZtnpYps1IdNGgjdfSfxfzrLkg3Ow5I2s7GNEkqzQ83GyQPJU5QYyMybECWCcM
KtPhV1obwhvZiqPMle80YvVzbV0QFd/bZlbPQI28IGPmA29UluyUi5jRZJJjMQgW
Y2CEtZhtGaWMZDklyGJMLedCqvzLLsQSpQcz306R/u3T0cSqP8KM3GrRFKqlVKcW
/eitmd1Gkd9WK696ZIp7OdoXTZOXUcYrLYm7FEo3H3MNYxEFbdCzU5YsGTQx1yd0
XflKyoCqzIRNOALEG7fN3SjOxIqy2njj2ULQXmsLseXIw0ANyUAUV6PrhVR0KaZN
hQGwfYkSoC2PHuXXo/TjoVoGzIfgh7E3v37K4NblHRWdw2+rw1htzBcspbgmNqxU
sqnBbFWNqYzUYbGkIZXZnbzGe9qhT9BmEOvvk4wV+kHKMjAGllFoHamKHfo1HfLv
0LV92CV4TDmqeZZXwWtVegf5UWNHHXgX7sRGtGPsdf0OZjMlg6GynBYnV+A1eV2f
nB3j5NiQ19uAI3IM4yrNDuMBBL7nNVWNJixESxy0ayCEQnjNYVKJXCDmroO5VbJI
+IPCNfdVYcyFLX/vQdklq5pAWNfN7q8TDNqIpFaHUdGWs4FpnDiPph6gWnQ3gZnL
TzbVO9iqCDR4Jjx8t7RbaxQr9qf5mUiYlvp1utda/DJGCnwoHw380Q1TNUnTX4EU
8aSGztDS0RR0yJgVKoY0bR70QSdTpIfetDDJczEz/TtT5feYEQj0eSiEV2/eApXJ
eutSPNCzZAPmFdSTx8BA5cpir2QziPWs+cq/WRZixLxAEtMNXY5ya/v6qWn8ezZ/
igtIe4ULfPuR8TiJ1cEYes58asqoy9r/9mmYztwgFU4km4k0FPFiGY7Jbbsi4qh6
BDsEd5lKs+4ZcjqJYAj/mxLxmn/SeurAY0n7T6UOto80SlOO6bLtZpJYxfoyCtq/
7tEWaSzC2fCIXgMIaweoYs/w9SZeNTXNHc3d6F2Em/deJ6RUaV40Ce+pxFXpkYKq
ZSUYeXQ/WjJV1M9qVQxzt6oVg1y3h7rfCGdpd422hiHHzdvjONw9kDOHFpgsL+v7
9rY8NO8s+9+ZxZt/g826WNa7g0wDBFpbVTFu2+sE4CueROclh8fR/XEc5Z/1aLGk
boHEBL+8JbMhMPBnfXS5rjsKzKoCEREDnzb4dMbjzh1eHphDCWVntLu/OOp88JWG
nPmFBxOfnVnvgaM+RyvklvAZCjwEBAzrc0s9HKpOxAb0Sp53MRkhpmuWw+ZFCv4q
QxcVJmr+1QUNn8Sozj/Vmi83YcHJI9HrzEBl6iAM0qsg4s29qhDWZ2iZ2LN8HbhC
sEL0lBP65qStB8YmkjN/AfrEiwJ6ooC6LfZipajtnbDkeC2HCwur95aZe1vwz5L2
FcFv9BvdGBHUulPU5ujctzQA3SKE3TIY8rfizO7rOeQdBCUjPD7UWdBMKT8tK9dM
LHxagDeQcLIaUn2XVE1Nm9ZL/Abp0sR4NzCpMuSBvcZZIcgwhaL9MBofqzgWSMHH
cSV8luMwAJR4LuTGapxs7EtSecdFLtNkt/s6ZxROvQrwlzyClWNpJ+4KiOheYBHF
dOFKFpdVtY8CoN6vScUoKc8xJOa1hcUhfPVRRfvF3mQAuJywGSumcAZJzeZXhXyl
cO/xBxa5KFauBnXdh5gt3vj+nYaYCu/VPIlV5vG2gq1sCVdz1YNYSaKp85JZini2
aUkiyi8PgTt9kJyKScgL/kAqDzUQmtsg+346zI6jfyjnM6Kp6uXKdWNlbDipZARU
sY6J4IeN8EFIY7gKCH2UDQgmI5scP+hFHVBFqTqHA3WPTFX6FAFDpSmh0icfjgYV
LuljEuRWdUMEXXQdWyuURzZMK2CnIUo2izd0mqVnYo0yQ26uNBfyyO2xGDwRtZ3m
WMZtgWwdipoQMHAAiOo/N+hc3UtCx3uLwzxCBDe97aEfEpMvMR4KR9Prm3QXtDBF
AeM0KGVOlyW4ogkbkNBOC4PTyKEaWhz3UvvRvMrYCV3MEZBGJSC4GmatwX7D9fBR
/ZDdStQYrFuA4tew+u9KQ25DhUj7X9aPH4hamt1/fNaAntMwUs6CgzY0cgvNnOY2
ubjS2hPwefisvYKADy/yix/R5Ah+4lDghBtuwXFry4S/g+x3hewIrsZ4WQBvV4kZ
VXD/fhpPlcrZJVbOxBG0a6WbKLkVB8RO2Us8+laC5E3dOf8e/1Ly3FIoqjTs+EU+
YqzC9BAhpfJIaj7Xvi1YpiMnmLD1iPgIdaWawhYbvRjlbK2sWmN/dQ/UUVsmxxID
locvSjZMmJHROYGvfYS+NEleYBLTBlM/jkyFHSXPQ5flz/XJ6JkZ1LreRg6SDRU7
twONo6Hc3V7fBJ468I1xoWH4KH5f5SrVE3qJ6eByg4NxzxC8gtSqYH6qzF41klNO
/PRwmTlsHYyRRGk1U5fRLaVYzhhkMdpnceEQ7IK4eP1pGw+ZUyPRo2S6g5b3Qtk6
QJ6RAP1hIJYjEUgNk5bQZfd2J8PtvqPpHp4NPklDE1krYeE7PaNf4uai4Pa+0GQ1
Kz4v/f3glPmadhc07A2jHW/ujUUt351p2S92AT/Ka4oo9e2i2MENuUPD9IWfoh8/
V2h1NaDwy94blmW6QzEADcSQyOfuTo91yAk5uA5sr4pDGpjvX4vXT5zvYOokEsVR
PeqvlJijrdwZGc9B/jE2Xon4BRolmL44ZnMCVEtOARmol8rRs1Hn7dbD6NfxkGX6
G7TIlwnLFbNXU3HjF63agvaXVrbWjQzPtNI5OJWEyGncLJ7FUemv+9KyPkrOxnAa
EZoTF/qHW2ijQ5qC4xJMgmU8rT38xI6pBwk0grlGnE5899JqDSmuxDJ/caPaRENT
l0o8j9Nd91xyVxVFxBRtwtqhpCrfXY58DfwsSlW+gqTDOxTYSPHjZgGBdcBzmKT8
6y9vn8wzNHUjHIzSGOsqBJb4wcfXCwwv/XftsmR8kxEI8MXBPVWUNo8/+AUFrRMN
nnqJiM/WGjRWKFsEkf0qQbfoRFb7UuHnKq+Ah/C/UzrJyMd2pLOAwFKWidf2iakV
lpMQcmIsOk4sQFMCHQeUVHVowKN/kf4cYV0ciucqq0wko7YQxa56r6bYxeezR7/7
WqofSQ97kLp103Wj9wVmjorrpRdATRanetYTE5ud22shZFY2JRWREVJlW+e/I1P0
omsTrv01MU1AESKkk9FYSG7b/w2PUDrI5TdmLl30kbM9UHXo5BMfA0w5xzVKQH80
81NZppyee0J9K9UuSYEhajcRPqDQEKRf0XVGUlJeEJk7NHh5JfvTg4gc+8fZjCQK
CYrnJwMWJ3B8k+EEDVt6ijFKCmT+mXkwWfx8TBojQUlqPXJItIhB/0UJ4SbJprpz
mDfaXBaxVDFBHtCEV932PhBijCAul3sE9w3MuYFVhDMJNBZvfdDmQMyb8bRw6K1j
H6sbjFlNqHYHpRj1vX8oUS2gNeTWIxYRGWePfR70F11fhOqQ6vi7XP1anHKDDtiJ
uBQuD0mxLnAMhj6zwfLdfd5FWGlj+RTi39fMCRYHqmyRCz6ROB+Ehr92itPqgFc4
NPWwjH6eb+9mGiPYb3/xH2rGSOC1Pp2IqxUPdBVijss/5G0dHS9BgQCgxjT6PM+f
pa0Okc8wKte+Ogr9/DDkVQwJ5TcYjgmqGH76Cu40eabCLIhhN9kBWJI2z1bqdN7Y
URXOduSZtBuh+2gYBdf8LScKfB5PE6wYAonDxN9BZrFelkvekvyyQ3HRFHjrOtYg
tVTAgjTINMppsepPN7WdppGndBkysrYrb0GnnWI9XXIel5gbb/ub9UlkmhzRFZ91
UbCokzOiEPrDWtTeldyPjyZ3Ru+neYTWX+O8esZZH3jkBaCjoMa22YYmDpwrfwSE
qxmqxxvEk8uWOs27fogsWXtksepgwUA3SI+zBX5tppYLNS6+KMv2ywHN+KDPFwqY
iM1xLc8Un4sr0EaMjcBkkc/rBez3E0rmvINYvFSqId9pS3mUr0OAR+zgZmAXmR4v
HKkYQXx2wSMDB4F/GDcuxWCyBK7beOcM2HOrDyN2ctTPoiJCP+ca5NfW9kdI92s3
VVuA8nKAMXnFnEME3yK9yw2YKdqd7nXryP+WBVIGiIujHghtgOsRcQLKFtVucwCT
wzNhFf10C+k5i12iEXq5f7cl/iMKXBQCKHe8seGfaQKiYfAgJR4TYdTWB5uKkye+
NMgqum/3aFV+pNVIkx4NSOprT5UhNwFPMOf0aGWlDcgw5skTyjJyI27SNaDezgAP
0zeIiigxASuVBpzdm9PuPbF6MWrTJaWKD7PWMZ/elTYvlDYy8ghimNekwrKAzJee
08I1S+MHQMQVOyJ3jopByXOfrcojwDIrmt4eX1bul1VQCFqnZboupNFfq0ChILMJ
7ifys+1TpnSO8c2NAKm4Jz/GvjR3T7p+JBvAKjU2jqZpuqiXdYsTqMClfsdtrtoo
tksynHDEVroW/BUEM0pDWc8YfVVPJZj95BoVZscnlFrWQbA4SQPf3KLTKQ79pCjb
rllNqi+xCEyU3yFjKU25Amq3RCfmyjb9dfhS4paslxxqbzdCGTJjHATV0TVXPetl
E9giaV74xGD4kuT/lFiqRT8feiB4QZoB+eeGEJzZ4lgLB7rLDNNkmLArm1pRJdrF
DlMTd8H90Vn6dLolEHuc9BCYRlp/1fIEJPbGepFpuPFJ2lVyPjDGU66xgpR3b7nC
WFlLQNYEarDghjIc4vJSudgCnt8uqKhpxWhDAzbIUTksabU6+BkXC8s4VblB4J3V
kx5PsnhMUJOWfVjGEpDQJp5e/UVGV44JJKzYAE5WeXMvC4YWUUAOpXWNyzW7JO07
dIIQ8Yecpy4X0HP7WWfcP3zhDKQFTS9f8KsYcl/R4/0Kq3OLrnZ8XkU2cvItetya
ww0o5U7OLM8+FTWXDv5J4OW1bLAtsTfSkFbbABv+SrSSGoBBdgMXG5aD4kVissW0
yoysx9OGr4WUEW5vRt1BFA2o1TlMyu3gZuo1YwkXmQVyJpfJA1r4vGfKGDRbb3Ar
vaHppi+81ot3BBc1ObxjLhj92rZXemHiu11VsfNa9EWroQW5Fx5mAEewUH2MjJv0
19BEXdd3fTtSWgY9+AykZgVuvUC4Qf8z4S44MpMbw4DMfCN34DZuj1nSpTEnx8Vn
UeAtWzmPEk+kQwmP6qBbDKc7f1mMfPWce8euF8CKEu0L8KMzvrP6kJhl3N2nwoAN
SMtFrhqBpRGzbPKb3BRI+cKeTXr0Vp6fzMBL2puXO0Xae02wDXj4RQBqk5D0aACI
EZJe0h06MtnjJWv83w6TLXD4G6XtrIN8kRd/jY+l6E6DNsBPmvz2GkjMUkfuK3ZV
R+gNvwtylPWkRU1lBDw+JvMQ5WX77isrVCkha6OK3fEYnHFqKhslP55rd6RoGa1c
L8CWKQgw7XvXAM/k4fJ3hWsq+wVxCoJnvP1jCZsCh7tOKfTJI4Gb+da3DLrXqwK8
WTMbyQ6IDBzATdHEe3t7EiBw6Z4ezTIlDIIFcXeL5hFrUAu6iSkRUa1un/UtJd9Q
Hg9FFTDTbkDzdH4ajbEh30eF2ZaiQKXJyuFWwU+rwb4fzK7+duxKsFZ3isvyXvEL
dguTdzPiKZj3JuryAo/dWK1PN/h90WFRvlQ4mzRATrUuOtRbQkGQCJQWiBCUo6kB
ET9zPyvlv34n/HcvOpygv8skG2iWo4nXrN5hzwqsCwBfP5pxKgY5RNw98HK5fCK5
9OdkH1AFGEpxBNyD224hLgbMFLbGl4rJIsF2jSyQPFYm3HkRbGzXdieDM/aFbAbQ
NAMw6YJ6Y2WBtMyvn3xvQqWBKF+Vgar6LJPMLDosIwSWFODtglzLCP5WqZlERYQ9
deROBiLmvVkZo1oXCojaK7w1DIBSx46l4Q54IINe5dcU7dmKrBCP41kBtRD91ZS9
DLk/haVf1AHrD3HVUz5WsvLsjyZQr9O3dc/fa7svRMMvzRZNYttrgQnCONsCxAsJ
aDhSZjWOsAdL3H7F6jr6pLIt/K9zTpM3oNWcDlZEgxl0Wou2A6N1MGNQqXF6U7so
pflK/AXCAkO5ZZA8hnd43wlFxX2TLb3Z4rVYtt99Sk97PC4JQ9Dh0gMe2KUfxcxd
ud4jIF0aIpDmh4FnH/2DAIOe2SKGl9sIhxtP2z6h6Bqaz+cTDfJCYj0SlGIN4/yQ
W+cDuijej2FXydHzF+v8yzsjOIP+RWvd6g5RwE6ivrJ0kVSssRgh1rKeC2XRznVc
O/QN2NmuEBGveYzegY8K2qi3mcgB+o/Q2gDmRHLMC/ZLvTz8Jpa5fuSH8xuXpATS
Z5jqfknI/EQTOxlOGhcYKylLdXz6IqRBIhtW2XbsIK5cAY7wdGtTd1js7e9Dd6Ar
Oo1gST1lZ2JGBNrVnv9yIRB5B9TW8PHBf5AuoKLv38ZfbP0UsrG3eVgrDZWn4jce
HDbx6BgWbmHg5L65EFQO/vXvhHWteYtE6h+V+yV7/DZCHSOMfpnHG0sbHdIGTeZr
lTyS0JwbfyIn/zO9CCFDvflMgMiDQj8cR0gxIJPDJ93CL4t4UDnyVFBNzzSeYxDV
SlkpwZ1CufLALZrXX+0KWzgTjsvNd10sH9WbeFCOCLlYkevD018Mm0kLA3cHAF1U
fpt8lGq6g8XZFV0DjKmokZ9Vbbnpi1GZmQeux3tW9vBm+iVatZuZaHn3Ai7lRQzu
LnLh8E26c7xIzQg7GnzUy0zHC21iTO3CMLMr8rXABPe8VKiml0oMtRoLzZVb3XLd
SmygzFsmaU4y88XYncVWx246dpWzI8Hu5xpaxvPIfsXEM7lPeJsDoRRMtPra/a++
PVkFzwwZFPhks5qmj497q2CR4LFTNYpDm1vXzwCY6XBCAG/lxoXPvimLGDezI5ds
4GX3oP0bhKwpQLRDo/EDz1EuSElbPwPLpKGGuuhaaCDnOUpbYNeiCvnwPrlVsTjB
wY4T+QvjvDP8dWde6hgltbfn1A0hlIfl7HCo12cZSyxMb3OmIUuxSPBefD87kO+1
KuD5f+HT4rO7Rox3TjVYA31U2rnB4HeA2895Ee4UE0UtubMHGNP2yMUv4GGVQj+l
lX10Ei25s51JSJEkI+dueMh9J6W5Vc/Pq8PThuhGeRgJ704SjCD22w3myWi6nLM6
ZRHdSb3fMN9E2+6DPYWuTJgPhQ6Pi30oMGv5k6LaBsXfFsvYrlcBw5XOIR/r3ko3
6t0j3jP9zPxWZaj0rcfsGJQwzWeShd3WGL3QMRyt5K0SgaO8kCch9cjR08pArnrC
GEBMhy+fU0BBqIUQMqBfSDkSD+DLzFiNuVMXf9D99/YUyd6cIli5mwYb3Y/yrgJx
0p3yG6tanePx+i5OZLzalzlXBqIcuSOUB1l1bUri2fEVXGufFPyBBP4wfzET2/yW
Dhr7+UG8KWd+i5gbTCZvoCWpHmvkepHQ1BHWC2sC8fSa+gwsJDK1kC3rgnl8HFH2
RVyuVZjTTCoL0zRWxadUvEv5KRMvh4qDZ7l93izbSbMnRWnrtLaejlKBQi/4aMOD
K+b1Ir57tjKa+7bZUDEm1XHXImhADv+8WzfqeO9kC7aEzzzmwA3mE1RmhAQyZZ9F
TtLu1Q7pFCDE9YGQGmlK9WR10nIVXvoSe1xXJ7Pjfw6eufUmqrsqkBUPE+mB1VsE
rsaG857c6vJU25CTDQUhJdk6w/PkDikaxZaxfQNm1VMWuuT93Exa6zyHyCZ49u+b
daqGYi1tkpBoUGlbae1yueefhGOOS4Knx/UgduhLB8s/3QlHFhfNkTpkFqyNQSjl
Dq+tmc2S0/q6zAN0WkLkm6eZWcWeMylN5i9S929hzKhGtsXpdmVbKly5hQSTOV+7
O4S+NPSaJ1zE6N6VeB8iaf9pZlcCDOTeYuBLnrgln47DNeiYtkcs5qC3TCqGep1F
TwJ71VtKPx2QuMo7tHAhLUJcE7HkRcj0s6GF4ILg3CM8Lj7q6BSoXj0zKmxH0lC/
bvPTApLoblCTtcPY4RzUhULU8OjAJ8/0ebv89FFqd+AqStAIpUa/SgL7nCUveDTl
PEbHzMHm6p1opxSYSLN5xdHR12bjBolWJfrgVDwhUFtLzuXMzf5IHJ+OkkNkXBo+
McwsJ3qzMxewjBG/utahtLTLrVCrznmXQf7pRQCqip2WvC0uTH8IrZOEQG4TdSDp
T0uSc4116oHC00bxp7fIS78uhWU/JKAy5hZ62lH1+wUhA1yEG2OMH4aN3loVUw4v
IBADt3n+iInpORFQOG54vGdeeqx0oAIQJsZSw+JnnVCj7zPoT0EOo+r9mzN4K4iS
hFHY07I46xKgfItIeCwe/ax6uNxnGBMOJgF8L12IrupOLMD31IcWpwoCrd78+bvH
LpMWn9UtlQNu+fjE7l/z9HyMcz/yCDOE81GjWWNY9z1VTNkVqV6hF/xvbeNkgSA7
PdGith/9/lZo70cDObUbBWdthnOCWEOv6Ge5QGRppjTMjtIjh6B2w3Hq3KXETjBN
mmkuIDJ2/8tHXOzmWSLW3S154vIV6KgaYmPWLKccOFjRpZVqRqFRoNoYN2OUOp+m
WnWKGmw8iJAZFGbQW1pkrDoFmsBsEGWbM9FfyoDClPx8xCP6PJqkMVLqLawdA8JS
0/xwHQC4pGEvUUDPzJm1yf+XRCfTT8cOJZzC5Zx883A0by4q7jwnYO8VZJ5ScFqB
8W5I2FN0XMhbfFxLfpM7/Tt1njrJ+MlpIH6nmxdHQTCL265wMksa22j+FqUK8cnm
nO6P6PNTb3Jqvisjd9ekESKMlzmQZI/SWILBNDKZnqukQ3o9mWfzhbFhrXitmd04
mk6+7LwcJr8NAC70jZM9Ecn7wucAhUd0g6PkZEoJaHN33bBafz5EUvmmaH0zabNl
AQUyrmT6fQKIx8f9DvAA0oLqH6XSy+GB82FH24G3rRD9vMWlaKZRS33SWCTiQ8mf
WjfIegN4J0ZKLWJMKPjq88bCh12dpcOZ6L7obBwyHrKl7Zx1EZpm9O4Hpx2XhHC1
/P/DhR4I8K2V/dhdpRKozy6ZezS27eNm5HvV4eiWQDBlYwd/KE4ItoFKGGFQhRib
NWPyCyUUvNhN0jsXoGLpdQX3GEtff23wxuRzVd60/sedwYnLnR2XNhos0PQqNZex
jmUPcW7FqO+msvVuwYsqMzm6eddFik6kgRourRNdrZnuYnSictqW0L1H0Ku2hQ+m
yv7SnbxHmpBG0ZL4giNuY5a3V7CXqjJi4iOH/u8Ox92LxAUJjuxvblFGzBXBK6Re
ucOlW28EaCYPyLDW01sAEDFVCkasW/rSawzf7mvVg3Bb1TzWUKhVIZ9mar86wedy
B7H5ut2OkpKcV2KVhRgQab+6f4Fu/iJvrWFcEYdh+U+1Jo49KMyRMbr3EckVvyFy
MNeO9M6ZVz1v9IqrLoZThx1OG4g3Ngc14fn9dZ/G3kWpu37Xz8zQ77v/xnSMCcfz
uKlWBFVDTkF9r8qcPenG9JbCpuWrR9QLKBpghaCzuYQeBrsStlNUxEi6BnPijRF2
l6oOTMoOfjWRcNlhKSX2ao9QWRkJBDRROU1Erq/1KuJrt4j2HpYDIXjbeayONtx2
rqZ/+0okKWl5gcenDiXtnnWC06izjTK55am6JiZ4mwieOdHi0KWEx7ZiKPM9sDLR
6KQ3FNdJuQweh7orWR5amPfKPjX/lFxrBPru6BIPCh3db8czpntGFwgloyOpud1Q
YVITJ2vYjOyJtSyLjeY1zoCUBPka4odO4ji8+lu8steCmV1MkXvT1GhFhIVfe2FJ
RUmb9GG6V9+SR4rUfWzKrfyDcyKoagw78ZnVehkPqox/k+yQI0b/1Azo57iAyAtY
ibypwtaSpVSnAvkvqEwlsq+RfA9WDwdBM31mUOcafEtRmXeRcRI1O21fBGNZGPNU
aBlowCcTteFEXCiK67Q6BngSnvE2g/XMDViyfbL826xRfYF+C0uVex3GmAoYvUAS
D2iWgWxufk2luDbkCewVqBe2/wuTiRLYCSUlrp5PO4LVitv9krBRBVcrC3WFe23u
tmtuo9lNiIShh+xrDtSn32k5eHhYdFZgvqQk2sIkc6b6E9OLkTZXaQ9KZ4y/QZPo
p7A9A4eXTG26O6l4O2kQ6eT7jGEscjUoSPjsIHET5hfP3ZuTkzYbd9xlJDNSV7wG
14BklBulAULAGxgcB9AsfqZ6CHqzLagG8NHASAZghMDdXFbAkDLY/D9oWgaBUvw6
H5+fRHCF9Q48/o+tiIn3VtJ57o+ZKeF5+TC7DVnAHAU23V+4IWUupujYnxoW5zon
E4ZUouoddJLyekmYuHKfZxAJXXXbyIGZJ4Z18IxBvWRYC3omtOjR/SD/qF2kXU05
v8oaW/8mqKyI1i925ndgH++b1vZnW6+X4cQMLSOqgibr8sdGqrPJii0jryRLaah2
Uj69/c7ChZyOAFDKjpYB04fpmki5dpBo6fLhuwe+FFQl/hwu5OHogTX/l4gPsHYI
WiUOcivRmfY7KkmQf13nFbFLpexG+MKcxVDIUzotnZxDuGhY1DnYLoXA01/rjRgA
nYJGIwJp2dKkzSOvitAmmB0t1i8n2tpCVZuf2yAFEsgEujoavBWPLVhEkAz3vR/Y
Q1NFgti0H8t4EiCeYPc8vRbZdDDy6LkKlPPSIjeWdjyyuQVXrGULXrdaw7+RH0O+
3jlw0G4D1m+bNactVQukvYKFK1BeIaByJaZrFLWRBcSmEoyryXColGFv6u2XhCFf
PWaVc2n8HuMf/B3nhelkuOgfeCTwAdrkoZjxQUw38nxGlC3O9QdHXJ4giYo70Zif
Tb9RKkH0DashO6ea0RUhltdVT6ignON1zgT4/bm5axAacrcGfda6eXZK5V77LoPg
Z4jeAN23zWiNNDrqCp2jhi/NUrqGtD+9Ub3AIyLcJxaqIFjGxQBcfUa1RGKr7YJJ
lohCUkJOnqHNhY0iQEbnyhQ3QJcVdOv/yz0MUoWpV/j9WRyz4OYZpaPQTSN1z3EY
amP14ZEurC20NbfW/KLn16KiYt0bIGz6Be9QiTr6rTnABAK71sHj91fsSDYL0LDd
qYoLfzpSjlIjr1z8CcXJj2eRdFHRZz8xnPam/2gciQSNlMzMIsJQ2v93+n6CiASz
IXXxpO7/LCEhUfkCj1um6Hg52akiuU4ZYPH8guP1Bv8PSl8yVeL4yosK3jslOL2v
3JFQWl3RqCiBbkfl16BSntmKW+HZG55M1zxjJK7P8SW1Euj0EqWTGRSHB9zn7FSI
LuL4xC1WJ71zcQr7U20Zu6RIR5FhBbys44ZTImMOhT+Au7mpz3vja2Q1f3kh3SKQ
61uBAxAORYzByNBgitLcyVSCTBLvsfaZMKmRVoSlxIovk1uvXeZLNTM7kMU/fUB/
gcc/7jK315Ks3xUU0uxn+Kml+TB/2bUr+I0eRiyt20R3Z/nvnRZt/RO8T7ROgMTr
bGo/Av1ynONQU7fUoX5bxZE1Vf3XEgJSdMQjdOaFIx59xLTm4PGv77bsIEF58Mwu
aFGs12Lgp4UZR3YJ/MSFBSpVryvvIT+QF4MfNgEIWbBiLMPSytnCkQQEeoPQoE8R
tjSKGYiQzjPvOxCR9lukcN/KjtoTAUA89s2aCRVRDFcai1JLOXa+6DyLiF+th/Ld
Pf8JsQwdjcDWrzneaucmBLnYEi5WL6g1vEFVAhK6MG/6Exd6QFkH7G+pWPPgmfnG
RjgytRmr9kSddLStKp9NSLegXWqdPL6XrcwEew//fulOU6VTRaOt3+L2z6sc4J8w
Dmi9KOGOilZjOGFMnSUQnFACrFklx3MHWgxR3p34vMtHQK857Q9rzGLVnJezg39y
6ym/TVMtCDA/d4dHQ1mzjpIcf3/18lXyCJ0HDDSZBJmKI9DQAQ7zevNDVuymXXhd
O+DakM/TkcvJ98HZj/btKFCY8EubZfpb30yuxQQ9kq4bXIltIuF1/En5WvJLLqoH
UWtLi2vC8gVLsEtwhd5HB/8qXb1D6799Wud0PmEOzLmtxPvkLNy6CyuIqLAmkdyn
TNs/bIUeFK4n89jqN3Aux9fI97dFhx2auUciRHKPlS6A8jwRxjcPQKpTvVVhY8vH
Zn6aUtcMFUszRbxweT9olREccmY2nS7dx9H2HKNUB5KDpbBX0vFpnCBRAAtTzlAE
U9tgmfjCzuPgMkECxuRFVr+0ZTawrjyzGDlFvKSpv+Cs3Dv13hB7khAyLz6d58ga
bq9oPm1gQLZDdeMIeFG8Rn4B2po2TxRUVoz0vGtQgK6KrfvIez0ZTNHJITlHufWS
h6ltDFaq4cErUS89tQmL4XfDjmLWJll9689RBofIv5L5mcyYBPKVITJ4qUEVvlpk
4pvj/lR2hGwgigpQrzAPDm5dG00gLW09CEl17ZrV3CKTnv6eEXMOgyYZOs3Ih4RI
aO0wTFI0vNA79BJpC7xkFl3dY8sQY3LBaUSC+G8knv2R/DxzQMik2Hrak5tSmYFd
csMKkYwp7C5ZLtcy0AYvPteqjhbOYMCZEm9aL0bE6WDBzLdfWAipmm41SC3LcbHy
ZHqDZqUkV0gdtiz6w/G8gK+EIu+OR+6KCFal6O+F3SYo27w4XV1dKvKkyfGelkwU
lrMxit/gyW/Jg7tpEGBBxou/q8N09CvZcdjOjT9FKB5d+cRAlDPHnruu833iImNN
ixeglpdwIWDjmq/LzuO4HbnpFE4hx6vVi1PfriXYNaBqCTsYiCKuep/JQwW+T463
vccqzySGX4z1Ag+ZAaRSmY756fMjc+GhDXl1HfMqtFIlAQZvl7DtDmE0fxA8eAQB
4EHcVrgVfZBEkLiAYjqmmkIZPaU7YRMcxz583pTApOAneDzMOuu3/1z39wpeYuLT
W30D1z123+BRmbfxWzZFHy9F611Ay4I/mZ7vdtTGnaKFhpUcZqOsE1D2/d1uPFSF
Axv99hLsgNZyxjST9SRvkZ9dti7CFv27JFdOZ4Y5j0BIEklCUfcrdEQHyhn3Gknm
Sg4bY8cRcUhTnXvHTs7fAxMQzow9uTTAMCitZ82PdC7egBmwsRIPwrPRmtqonZsn
7Mfsa8ZHuEPNGLtAWOS2z50ZY2jW81L/qQt9MZhcAflheDMkw4e/WgupVt1mbg7D
3i8ec/ALwRP9cYSGEIdw7EEiTgSKCtAER2ckGVh71vjBh2GVIhUH2rhwFQhsg9Jn
cEo8nfsgWWMlUiFMgl6jWRSTYN66urL7Avi3lnGL3q1Ul5I6GuHBamCJVBX0tMui
+UcO6Xri20wCEwcwLI/YHXyvmjKO8YAxCdLFDHk6sfsqm+w1bXC0GlQiNOlNIpaW
0rFnzzB5aA5VOaP75hnnPjOE1xEJgtoSfZARQxA42cXUI4Kz2Osyfkvqr2R3x4HC
y+v4Ep9fwJOpWc3Mb8qXcdqx64YwhryBoZFiUrFzrU9Kk96I1kPSl+2eVTqhKCrU
lfWUcJjQeWoBK2OJF/hhqr8gyfIv0vvJRZNTWdQ8Ez9tH4JPv9BqDJEO+2201hO8
x3PgB36Fd/IO/8lzOetQCyyHtpaRrZS/jjAJ1ac4gbrRJbKIcahGE11uHhDTZV1e
mafYxO3/s78TrOy8szqIpSqeqzLpD6dQekx4hO35PHSIvRmp77AnT8NheaHGVd2E
w8PiY9B8vQIzVNRv6tVlyVF9vaDl/wFnJzCBWSqxvSq4ixJSigiDLw5rhf9yteTV
MwItxmLDlQrvoBFtWEva9Gtl2xYYsHZg6mODafHdBNKlR93aCnwLDi0mfoQCVvJC
F3/d27QrLCW3EObZfXPpZRs28hgbgOiOFOEO+YZ4uJLvyP27XuLbWu/CzhHRLs7P
TXNKWTvwE+ult5E9MWbzBa3E09eZlWnPYJ6POZZk/dUC61L5W+hH0S4Ly3wKAHIu
VLzJEl3ZOI8L9Ghq1x3lrd51fg0kCrGRVVPx+6cAH/ptDwZ6i1c01LL5/G+WHzbP
v1s69DlWGp4xlRe8TW8wgwhVNaCtMiB8IevNluumYTurShRBScMOs6NdvsPhd/8g
YzMb2Z1hZbiW0kDSmZdauFYRMRz+hbT90ynrpLc2viQ6Ddxo1Qfs8/fMMfgKbMyD
KC8qLGEUYfHsAYPxROhGYPyVSxwtDPLAkAVZhmKIsJ3adjHNe2Vc9+9fXPRhjDQn
Q4qs6G9+krcVN62MZmBAWPf46LfnYs+5wdtYpFf0/Zy1pm76OPiYqplAlwurf6fD
oav4t74FTPe+Iy5FBVjvUtaD6pNAIYlIh1xbiYRA52iE4dICyjbQief7l2PGhY0O
BA7Su5oCV2fklthDzxitkfhZAT7Rr34zSyxYkNnA7Nmt6YltS7AvFmflM8QMDR+K
OBrIW0pMXyQQ28tJKlNhKRYBYakwGYbzRA2/I1iO/urra/BB33pPH/UvlX95bIKq
v5WkQfrmRm+qE3ms1CQOdLjcr3oaViFqNSR2zNQoh7gquo6znkL5ljI4VAsBWYGj
Vmh8TzVE6jMQv18s2+/NuYYrSUCZNdRL4foclHv4bAW68ZdSNb5/yScyJgMSqlLr
Sz+dWlcMPvjfNUULQ/szWNJrW9SNeQ6LFuCMbJQMlxh+zAhgj3llhRNVkPvfX79H
EIwveoLtc0DGcCBJ0NkS+KKqxp6Y4fCdrH3R9Kq7txIgTg/CY1nH894Wh3nf5hrr
Qzkar6xexFDFhePcbCMXF2cWI6RIIS+76J/W3eRVfk4kfdsVDSlFnyfVRS3UC2+w
urYhLw9xFkEi041dOaA1dJkoFz8SNXXrpUM27AViX+Ytz4pRQsnmsthW4MBt7Bhv
NF+Qn659tv8TGPt5AH3JfL0TjujlYlRZSECc5BI+9Bd1TNbr/U/C1QSo3wvZUPfv
8e65ynUXL1zzIyDXF+TqELkJSeFfYGWESAUwfGzr5pf+xUsz5ksXbPNVUo1VDLjF
ZzNW3mQZWmwFprehdP6S/lyklw2/asTyBvL3TBgVqbm1slN9P2qlc0KESqc3EeH+
UriVAwRvI+obtct4TxEZJvLOnSaGTnee0mpYTYNTOgWIk6n2hfcXnddS+cto5Nw/
v6Qv5Eye/ULmtvbByOvth0n2g9sBGyqIojgvDzRo5/pNdyM5v+QtQtzloz+J72K4
uH/eGxYQuJ6DvzL82V9Fb8karLzkSFQvncqHaa34/OwUl1uVlZAu65S77K1+kfrv
GtKWBgQ2dkyLcwMbiw1PphfBNPevXskiqy82PHyqXs4VD2jcbN1jUT0IOZInqgd1
UUjQ4hfbgWO8qz7ODugmGeETmICXRU19X6aLDG2YtEHq+js/UlVrzIrxICdjk7X6
Ef9tneVp6aIkFeGDZyfMIurbX9GSJXYACreJCriOG/Tbh3WGgnv/uBlWCjJVyLjF
b7J8bRVBcJv06qszL85JXUOhr7E9i3q77/0pjYyCQBlavFgU9JsLbsMkbJF3Yyay
/xI4kHHI1Crd69JgxAzdmCEd9doDVnk0BuI5JrA9aIJ/Y81wLdZ5d9qEf1qBc49Q
iNH9hUN/xS0Qag0ki6c4soC3FpKkjWpQQl7f/sDYYvcApU0t5+1uZzCLJ1zxL9Na
Jx/pfPf6B6Hbhezs2h2B7UbJubU6gDafUyg1Y+/XDfeUwCrApQP4qBeLM8Y1Kwrl
CHkFEFYiYsba6Qn2dbJwXSnrPQc5QiacGmqREyuIRT7dN2dTk/9hfn9RITqREMCf
7jqOhOmZW31da0W1meV70uxsBIdOG66XTge0S2CIYdhSFf4GcD0PoghXev8/GYtb
Cj6n3DUPzSKdmhGgHDkGLCUfpjjBKTsA2WU2AaTKz5KBIrVZT/VZbEp5aoa7+tbK
nuaNDdiXgbq6qPsYWppKHfVlOIqhOH9ALNxIgSfgXu9Ax1fgTI3Q8uXXmwchkZ2I
mR2R8XuO2XfNOx9TPkb2kZdoaC5wJ7P6r5zPlHi9fEY/5bQ4VY4nuVZhBiEKia+m
a9Zv/TlFMEH8TeZ/4Oh3v7aTrJUfmlLJWNHc7r40TRDr9OusKoNLFQfFo6iusOiZ
UqrcXQpvfSEqbYFVnydJk8mYWcFkRTAKQF8JU5Nx+Vof2DcycG2+hPP/W1qsOQx/
uyJt2ztevo09c4czspXQUDKmgtJVJHc+pKse/SszAppUQ+oRVCpruafYwo4VFKTM
4iQBUYaF1i0M5dDQhrMv+5Z/tRpWLXVIVts42ghma1pJXk2dnB52r5wYYZKx7uVp
gL9YSG/vIy2ZuCYtfSPw2eZ4hv1orTGrLe2vLUlqEUiqbyj4oLxxubgYBO0jfbKR
2OgUMOLWTYwDcwEM1NSrq1z36d6PV61p2ByL9sRvlhgfHuhj2S2FaVAVckUewz81
ZscuicGSpqQ4uPFd4XGlWVIHZ2IhB/4Yh/4v2fdFuybECKTuWcZMXDxbOVgbvFp8
Cw/P7TqmCFJlef3jIxh6FCOPsf+u635WVUBImalVUF49OWJ6zB0V668mDR38OaXS
57aF+9v7D6xiWxaU8Pm5ktm2qTL/7WTNoEuuA5iZc+gstyd8438rzB/byvgw46ik
bNuQ9JrUCdilXzaYRVihLC90KVmpa8OWR/3g61C+rqVE6qr8Fb89xmAogKkYxM+v
T0WYcW1gAAbw95IPlDuziTV/PHi+3LAl1Xno5p0T9Rm9BSEFdraVpffznoZmyYaG
oKpxACSArq7zNrcp77PZsH1/2iDiGKeGBmbgLPwolTMxHrSSz7SeF0FeqqhGqelt
p6hQuo6itTAarDtPKk4s+/IvKpQMkVbhjABQ2+yTLbQ7bsjjZNknvPfDeOUBuCkV
F//gx6ifOZZ63Uinrn3NU+xkpf/lurMp0SQF5rlzECDiL1/6wKOyxW/VQ5IKa9Om
7hd75j+uE5NNQDoVzpGH1Btbw4meBiLXlylT+a35zKskf+JDJnqqKFny9AbSop4E
6yxMTyWL9fQth2ucMZnlVQN/y65tfaDWn47p/mY/l7TJdyVw+vdz24Zc8Z5kJZUx
f+y6vTsx4AqDA9PhVaPS2/+wcYdf7suHyE3TCGF0R/PqDRiUpgPA6am3ZOS6aUTW
UyUO/ywTe9IZ9B0HXfyujsA/Rgvrvnu8cGNwezeohSq5sTJIcgF9tMljDayyg7yL
sFtlOdo7Kmh+dxsz3XenWn18TT+gwIdoXhw93c+Zv4l9qP5LdlyhR7QDVxMrDbST
fS0bjGcLvW7QEdLXIiddqd4ZXc9Sd3Ud/k1iAErAMSMPmw9HrYvT5CL8hsFmOwwq
jXr5QrPdJ4yGfbZKoCXr0hESRd1BfWhqIkhGHa59oDfT+JWkybmRpXKphvz02aWj
XRTsvQOH4MWnKkh8Gkz62NXRvgqCk83uUhkM9D19I7X0f0QaW/SC3FnLUSRd23kx
AnwH8qh6jJR+TMMvyDHsf8uJtOf7q+5cGkO/U9tkSLPbaMB1+40WJYiWitCS3Pmf
8H4M9MlZo1rDqAcCxmwe2VdKyjBC4967z/k7xc66WJLi/SElF+0X1S86lQFdu/dS
CDSC/ZH6CbD6dJW5o2SIXmVhtJW6n0NSbt2Eaqk/0rJ7zeTWvb7Wz7sepxPvvBQU
eHze3C+re929/lvFxlUCfEmS/91Wem0TyDSdaRcj55JFAwwcG18QmdGQ4D8tUvf1
2qXvwlt/N3Mn27KY8hRqsOLYZszFNKD3fuATsmaUfK4cKusbfxrLoX+rphRogHNG
AOsZ+P35olD9waJkkd+/tIbqEC/3eYR4yp7kgtPdpyo=
`pragma protect end_protected
