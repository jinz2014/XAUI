// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fBzlTJyVaJNYD3EGsFPZCtohbzuHhYMgd7pLFnnOS1mLfZrmfHe4BGqHAj6sttJb
lMbKYrNQXs30KGtMEh0GVxZ9mQC1HwoYXHQZprA4zYMBzTzWJGbsUz9ngcj5WdJn
wf85q3JKhMSMWHT9WhqmdDPSaXhLQX0M+BDcxYE0xD0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25536)
HhEPR1mszjuD4kYMPEThO0op7z0Xy1zIMfe4eUgKZUTyhxoRqY6K86yH/BvE2Men
MlqoukcLRCqcGUe/HJ3ZgHHR3+dizaTUz1pbclknCiwD+gfvLZlLOrDbC09KQ8XG
kPPnV+bU1Or4uH9zeohj3IR3oSHQnmpyjyNDr9b++qFhuLrket9I7sMaGAOe0xH5
scKSyl/3/FZuO9RVugARFd2zSYY/Vnvk7aRu2r5N6aX3ibLfdoOw26Hruaz/6uxz
50PqN06tELNCbCE9NB2qGsqX/5K9PHPLcOXK1www8PzQshNMdeY1j4gsdiuEt4WY
IApLH16MJD/Ya+I+iHv7HiJ1aYIlZVfA1+2xWjBX0ep0tuUwPfIUdaSjRkw4bMCV
y5DwAtPEBB6lGk+JNV5TdLzbDe3CX2PQGAWeavcfUM17ZFUWmuBlYxakYyyctzrR
YZJ/0PoSDx1WjvU23EQBXKoqvEsg18Yp56cGeKeA4HfPmnbO216yQCsGgSEOG+L0
uLXSy8ZJYFtec8RarptuLOw+pimFWVH+uf7hEVdWoaWBazWJyrYVLpiapai1Zx9D
A36UjDlZEmICBM1rGT1cg6SFNmSpOlW8jKmYvGiQke4nWG5UnovBjk/kG+xweBo6
hj7Bdtci9u3dL3qwHVCJwOAyP7VVPOZ7SSCb5P0Np/bzT3Cj8LgRZkh7/txKEzf/
Wly9EjzIvk0Vlbidc3pwwv/h77DkKbc9FdLwfmjIeFoBdBOWROUAtlNUb4JzUa1x
L4V7FYvLqe1daVxyF4IfXqyOz+Q6odxVQAkhxlfhtv+yeNuMy6Yl8v3KmLlJJtZ9
Zklv4BpBK3bn3gAv34hpRbpmiPpl9O0y5+RYAQ9UhGoNKpwu8hsGLIcIYx2U5RYV
qazWtIC3jpSgL5KSDLzq33gmJhNITLUg1OxgYUr3SCZ26D0y7mzKeOo0PDX6CI6C
5XyPoGlagrbl/A153k5F7qNXAOOpzphSY4VyjY0x7K4kiN2HxTbNHVtIn0KpRRRy
o1FL4sjE3wWGJPwwYfb7vGEeFZu5vyP06s+M8SZbrbXjw9yVfYNC65Oxnc17XJGY
k97J6SxnVi8QNwvmntRu8hn6N/fvrUpkakh/fNIQmjvWWu+CZJJpv2baPKGgmfXj
D2wfEMP4t0mItKQR77xIf3lMNGUEYxOIJXM4uIIwc0Uk98ZiOVVdjR8PvonT7//c
p38FlYzLTdmDo6jrQfFhsqM1ZKI74xRoMFsosQtC8eAGMSPTnmztOit4NjdqsFPb
8/UFEhDEHPRu9LiJKnkGZtm3VVdKsdJpxektjeJ88BOOReOy40bw07T+84VhIu2g
81n4rIJnLVQwuxmOlMkF43TgOAVMBUFyyl3+3go8qWU/6WDIDUzSnsMfNO1a2NKA
DninMQDKGYwcQUB2ByvMnVA7jjId8CCkwzGfsySc5+0EmdbHggU/UyWx8po+JQwu
LbS/DT9BSp22qXeHW1zwTU1yAl8I5fxw68prZ3PDBKODXlOXhAQjjBTVMVmNz9wg
KcEUJf7FD6eyzwzhejvZAfaALswvBndpQeGKX4tLXW4mZNAkYPwMYhO3sFlXyVFl
DVkSlp5FZwT5CzY3SM3a1ZK0ukfzmp/Jt8sxVORSNXyLX8Zlr4ZoPVDB7mByQiCZ
kf244ECALqGJ9iwXa+81LsNQtxI5naJzQSlbHLYVRH4SDDuLJ27/ZmZZC79kIx2I
NX9d/Ik7gFf76ifWahKFsaRNrRw8cUuqOl/xEK+GOc7VguIqr/pDdOVk2eCZmyHk
2Yaq73Zw+vON8zYO3BasDdKIwUUcJNePY8meCMyU2TqkqUz6in+VnuYuZA9XTkGz
P+k5+T90Y/LqEUfcx8gPTB1bdV+B2ez4z1dwLCXBE5KabmjmKHN2C70G4B4diFCi
KGXALVePKCHaDbFBBTu5CzNLBhVZ1kr9FnXTJS9K4QK9tshTwoTXWPprwZh48xvZ
aoiHC7RZVZYNwGD1XMbu94Y2stpBddPftX4FLsy3VBn0jz45g7qJmtmI+JwSyFgb
zXz2te862ixdCFyyuW9mXXwhmda7gJXy5Sw5NrqldKEsKFofJXZlmJBICCmGsGxb
JskW2edNPEtHAQO02TigOJ7fy8++xNEp3Ecacs/cENoqflf4c66H4h8DpCLAcEQH
mEPPWHn9TJ35OO/YZT6eM3WsVFaG9b8/DyfxeSSIi1iWtRUW5x6SiKgmy73rMdeR
jyaRc8y4yCL6zwgHnOT9+Ef9G+wpl2du8EEV/ObjX+wE59XVPEfuC2bqjxaUYPxc
j3uduYn2s37vWDf8DwlxkvLMYeK2qHwzU3P5ZeKnex07YvK4y7HglRKxBG5PCATb
26G1PYOFq4dh+KsHFmSFeqqbx8XOjI4EL1Q9vErxfj7jCKoBRpnMn0CfCffAd7qN
p8KCxe9mCa1XNhCUrs/Tb4nTaCmLtxIsXp8lvdGWt5fZOXc1QPOhtni1WtIg6kln
mP/uKa8A5qYqOrEBCgNMLYkT47aGGtxd38aBmB07TtFEYOcdV7aPQYAFBfYyfhRl
SunhzYx2AeLqHY4FzNtU3xpomxTrvzigRiHB0wQfI4dh/NXcKRH9VEGBv9ReVsXF
3x0kvB4qOwZNQPPmNmhfBLoKKu1J56p3NDEfaxomKXoVZAPpyy8FyW8/63dXHfVv
5wrq65D8ro1ZZ3zuk9kcBlatHgbPMGvZd2L3LvsGEAmblC+zzDP9OKHc1Q0HIups
mlbygolFDMhsau1RUuaAQYw2fq+fRJzlSyo/YTGzPsyJ3oKFFuoA9lzTO9rt90Gx
oA5y09A+0++Bz6mnr/9yQ4fmJIUS4XMgtS+g4xzDMZUii02VLhf86S0DkI+IG8+h
VI7Iy5QAuhI3PG5MiVswIOUEMrghTjeFYBVgqTEjSqj+ZL6JJ0wiJTutO6tJiEFR
Zlo3kGLiHTU0iddWU/zNtGW3wEzyiop3P/9HDPJW03v1IhTC50hl1KxnpkorlfoM
BXFHtgYLIn5QQUGJEEIIqQ9/eHntlGZEHEhh2aAXqbvKbc2ulo5j0/Swj7ftzPk/
oBCFdI8NKNfJYHVukcru7UjK6oUjkGtYNBJkA0TH8FnwoGGp6Gbd+gjJsYHws9j4
0MWIJp6f5wk6Vw1MgoCx9YyKCQu94d2Obgwi1UbjcTUQC64ikxnPJ5qvsZSW8vj6
gvYieRPKMez26tlfp3ZErW1EB58aSC8YKJ0njCHlDjve3kzvDnqE/Qx2NANkfWEa
ttadDpfjPTZOnpCHRJonQwv4yIVvUXXKdaWXMHyl+Pm/ym2HC5djMgD5OhbbjTym
mlUV+GWdf97SJxCuaDtH+Jl40XoKew+LShuVx7P2L7/X7EAYUDLvFu5PVHPVCSzD
dW79vqVftHDPKICQWEpWK8Zfp2Yw2vUhlAqOS8mqDYDyWL9KmQchvBpdKRjJQNSj
MNNi5+oyJQgQXagMIuxp2rt1axivJz9zf5ENwye14AJT8aRieBx1FFQV5YHantvh
6xYo4w3V7+NS4MG+h0gzcWaS1EaUqK6J2ng5aNDBGIA6ZNkbFXs9RC3PDuRfkt6r
4vd50dFNbN6ZErxD12vteI33xZTAuWSkybxuH9cHsmm3Hb1As7Ej6ePXy8Llvvcw
29mcTqFucqjpyRMLfjKrBTiGh/0b50ltqt0HAf5f5WBTlkU3HoDMvx4yl6W/+fXn
YPdFSyzHmETa6kWU3i80hBePBtbTaroa/MvJ6njz/Hs7+k/8caE7XrNF4OaRNgcd
Ts00/BVDQSJNIqUamVBHyQyUVowkGtbrUjFAQut7zzB7ip9nLYy5kkQzp86ugjgz
i7R0GrufEn4+vOJ+PMjTPL4dj3UixlSQZSqejr4QxOv5NRnuSlkSYgxFYcjNspUP
QmT32u6s7zf5+iJQkGFC3sW2RmEonnqAg9EOVnbkkuOPyD+c+3k28mCU6Q6sfSu2
GBnU8vWOJvSRZU2crR09FUifEj9sLi7Km3eBEzCGUHD4/XqIYnMnEq1YHdrg/9OC
phGS8cl4mGZ/S5OxLpDBukP4smj3IDk1cJG7MGyoWyqRzK5Eqyob4A9ZjOTHt8Cx
QGEAOjzrYbwrt/7m2jNl7ahks0u2lWsZTdugv6oMxsW3QVsM9XvlPSxgP6C8n6rr
WqqRlazRRuSfWUh9DLkXqxf1JIZKEQvf7cXi0u2BOuAAquKzBZzmHrV9hA9IwiCl
JqqCqDTs5wXglFNJHsNoUt1If/1TOK5EGntE8vVLBbFWJtgiPvYpYsPl0clx+ca5
10uElYbeCjwrcu60H6SGNSLWFvPFJEFz4yD7LtisjUBunGj53IbNirsNpUvl5goz
RR8ZOOaZ/7wdrPfMQKzvh7f/FsnA4zD7pINIKhLzJIlzY4Bkb/KuvvDzhqCVN4hD
0ugKRO5/yMmoPx2jBfwe2zN5KJ6PPZI4ZVBIbLhABAh0rmrKN5jrBnvDdkGd0sgy
XIRviCX0GhC3iFJNUsoh2ZnTvjsPR7xu/Pin3fiW6a7H//YWmKrTBhvRUNWaIAx+
ayskGtjxUvMQ0oD7YJ8Ai4SfT+I9Akje7n4DmoOUfUp611d7Vay5YMAacovYt5U7
hliw6Yq6AZcxYUQfTCnTBTTeK1DG56eTfx4d35bcrNLV/HYovpoK4zL6PUiDsau4
bhV/02/n/yfaVtPKGHZMFfwLIXAct55t+c69oOr9QrfLxswuUNWvlLSArY761N1G
UvkgiuJpyBOQWNND9Agr3lVWBQWVW0zbziG3JdDy1xzZpTRhzQ6biXblQDoKInip
NMzLz4Hi2Vay/Mh5s2YHPLK75ahKIU10JPyUs0TiVhUjrw9tB27hgoqMgFw2nQ0c
4BPcqMGBiqly1TVSf6ebYEHDGkPGfFqh3csvkU6Fc1h0XhJYLs1jL6z8h2rjz946
cOPwI8ZV2bVMfph4gy5p3Qrk2RzohKuYGS+SKqyuxg9j2NyJRnR5ShMawRT9xOJR
sjhLsUsVWZabh7iVCiT3Bn81VRm7vMxHVc/mv6ojktBlO4E9HgFboJQyj47F54kg
B4vbhDssiPQHI/L0Wyi8bzRU9YqMgNIeS+Lck3yG8AXHy0cLbRl4qb99HIZrhk0+
PnTYcUQL/7Bua9w8oKJXVZ2xOiG6Z/u9oYu/ZHIOGF1H/57UlWfYjISXxXhNy6zN
Re/n3T1Ekfv+DWAQMHHxxur2HILGH8JjnWWSU49LQWmOr4Rlg0irXce/BOq8MIB3
xWwubmLeBSdoMVvyjNkVgUiB+lnlqM2iTXns5X/XvIys9WfLIDF+3o8r3q3+1igm
XkM0QQB+BsiDTIJCtTv9NapAd9eZvW/dzfSEVKF9NKGlBgBWmGm/a7TWKFnhPU/u
aF26auTNZbKU5vBDB3GvOV3xw1nvduqJGDAFYHyauj8UoNFIBrsVc6tw1cOe82af
x52GGq4d7PePVs/GgY2Nto3FY5L7YD2eB3C8Y2TZeeaCjYUlKZF1drnTCdsWjmKc
jehZFJp/5e3ztdRUjpZkaBRq9+0xdTw1Bbt4XC2L+ushGCgSENFP0p86yW1u8Zth
hqQmWFhiCm5JjAcd/IFAhEWeVDQY6dF4lzFScygwgygS8JlP2gS+kiIvWsVJcbma
dzw+xKisbzQl5duzgYVxhXR3na/nKx3C3CNiwqdLYUb8NYX8GSQ/fU2R9sjXCcpN
usPcrTPoy0ov/axhx/yeBx/op9zN7tgBcEl1c9LsjrO6pF54YNWlZUjYcb3NyUsN
Dv0s9J3XD90S5krB11EK+hBBCMtDkQjwQ55Q2iBnK22Z0vmp5N8aBS3NGzranyJ2
ENqQc7/2I+OaqseOAjknfXNvvmSJt1NeQmSg0tls+zdbwkTrrLsyUDtDB6brtiHh
Q5sfLGDblUyZ+IHRaOGJpdreKUi92MVTGHgJiFblQCES3CWHQ1WRPK1DnDR6er5d
5JjcsS5IxqlVU394/9c5jmv1J7N1djVw8azjsYWX6YYeuCFZRDGr7SAfUZyVBvMB
OvtZWcDfqgIhM7OwxzfBGtxJOVDrvEV+wZKR73MBczPOZ7r/JtwpsVwmOtRGgYM0
OF7qZgOkG5VZcXW9sG4p14KMHiCva4Nh6A3j9X6dF1rHpSEcrAuO6mF8tFmVpkgW
PoOnYJFPG1C08v3nxD+Wlp85uWoxv1B5d9/wyIF74XaNHHw197ik+wryj6AYlTlL
QL5VNceU5jjhzEWFqAF9DpIWW4Xw4/Lot5NjAjPKtETqpukPIm8AprgYEl05arlY
Q65PzfyI/DkxEvJfBxlqssOvzMGLKdO2CuJJTOa8gzR5Bda65klt9PL5FK6QhAJN
OLaiLRJpzZv7yn3oFNGVZIudmkSCQR+Y7ufHBAuRBlrJ0iDvfgTGP4lah4759RR4
XjkjY+K0FoBs4vo4zTwHFg1klnCVNgfi3Hfm7bo0YEoBwspWLJiF4JLV0NJgaakP
h7VF5nAioRdCANaFzk3ir2Et8Qh1kZ0AvFWY0nZ+O54I4T2aVAfDoWTycz1BYRGc
j3dDgUfqQNcVJwJWeqj9s0drnDt2wRsPbWLWF4MypMlfho54PYbqgJhLwwYon1Jm
4aSvV3ownHukO6uf0KVOin1xmnYApaZGY6BwnHMrFx4nB3CW5z6BwN9DvClKgpaR
2pgqCWXvosKwyanzh/fVafm+LqccFrEYLlIqCArTSDBE5M4v0Ds06n/q9X4IxYOj
d0SV/MiKyH1gfxgovJVzKKbvvJQ9HimVQHG4XXVtvmizuXWgjsGwWj397hjfI3DB
uCnop0ghUiz+/2/3OgOI7PegILFJ9dxteH2VsiMIsb92mRCo/W7XYq5UCylRy8vP
pa2Y1Ii33tW6zI133y75Gsh3XHYjg4sj/fB3/mNOV5n/diLJbIjnnpfYM4JMjMux
7bzmOzmbZO0rdL0R9iHqWScIQnaldHKuReDGokeh9euUMCvXzfigaPbNg3d9uXXq
rcO3jFcST95pOnpUjm3o8kPLKZSUM3xNjkbeRGo15wiJ7fIqqoiz2HKBlYx+T1qr
JLQCWbb4JZO0HOgUN44cnyF/VwC96GN8GbfFhr9YFfA2uQ36fBzzVJbrYJUwpX+0
wB6qGDNUpAilKOiOxwKWJAOl5De1Qx84rAkoAY1GgVTQEeq97WzVhI/jYVefrChA
JNnlsylomOGf3KVwvjCk+VnUQ8Pcb5E8Da465Tz8Q7h/+aIP9A1ptBFpJM2qlwkm
Sr/ECYbC/M3NhQhe4IQl6lGeTNoqtfu5FzmQqPiHedakAY4Xb+0Quscsa8HMZbV+
YrziOZaAOPpc2t7HhDKrSWz82nUAkouXeATxOP2Ez7VaT/duVl7QF3S83GdQUE4j
wJlBXgLb137OZt5+k79tPWxk4DJKr2pqURP5fnTBGmzxExchJ+etdXChSlsdQ9mc
lIz/9IcOCv7d2FBmSOItrjH1xapGaPz4GLxENFQvncmFZOfibgIAkGNIOs8wzyOV
ZvD6DbXOVUY5F+7RTVk1yKRW776Arwf7lS61K9slJ+kqGEjznswsbFm4gih1HMP5
bzJSVjmhrQzwtu/eDWoOZsnGnrnkCM2zP8x8MhfKKX7sBqE0jngqQybTLRkzQrwu
YU6SCzZeuB/Hu1bJ460XJ2gkkJCueMmYGwit5InwX8+tVFk6bueV3Ph+XrHqsry7
wupQ2sxBv90J70uMkaXqUYFtLTkYItraZeV/Yz5moRDGpyeaZ3pq81obg7VTplu5
yCYKN81q7Ep39pijC56QiNXp5l5zpHOEw/shQn01B8bGHMwq0BQtM4Rns2pCH4Kx
v7b6MoMvCPRzPfmQCqre0vTsK7YATkPx7RiRG3LNb/YZrekwanEWZhcmnFMNzndu
9fqkCKqDMtO+fA+yJdDm8Ksl2hV9WAtqZd4HeaLffDCj5akGm3MjOuAJjmeuF3xc
3d2FFfavPYfh1gEL9PA/y/vOerTZTjCVuCsM0QpEz+S01AiXYcYqu6ZxMTZFx8+y
x3iTEJwm6XpraFuiOlzAuIpvbhXRz/inGzHrDCHLIWdn5EHPkxKP95YBPY+UmrB6
qiJF2ofnM1uzW/qzrgZ8UiTCZYNgqyQwHbUNDfkSMqQrAEasHEmuzMoBeIW2avnU
sqVwnFj1hoTn2KIQ8aYXRHcHuLmUFHJ838L2q9CdObTfaMjah1B27eJ0iJtBUos7
H5kS+9gFd+ldEH8rqe5X3mEIUjpzadqa/AWaGCF0OZ4xEGYJvg1Tkc35LDebfF6r
pU3Kr8F1Hopi2Q8XyEVPQDUEYUopTmxl/UWbYl+nFI/dRLc6C4lz3ABFUjka/uOC
mhFpA7ZND3xf94kM1EivfMEuHWEy/QP+JisQKeTqsO0ACvTysp7AplBKIZMdSd66
Kb3ixtzZsvaLegAG/Xj+ikMGZOitn+jwLD3/ySw3uBSgJdPDCK75Mg2o0SE8VDVw
+YCTkWKA57nm1G3mgofDKH+zdh8P1LvRVnIZHJds1uEajAm3pjJi1ed1YTn3Zwiz
gtVJFzu/eyXjQc8ASM6gxMl1xeBGfNAaCulna4Eui4KxkoEiaeOseKA+eR6oTKHi
o3Ljh4ba0JPK7gTnTKvySQ7KGtgrWk0mV5T8a+iOtAuqeJqs2FKLM8FWIDncxYIO
kmlquXSfPBsc9sfYZuOmckxa9FWQUV7uUamtxR4qTksaz68+rawCk2pxBwHAVsHV
5lugJ7Xs60Cna2m+N2FpFTBtT67U6/jkWQlUXC1i0e+W+e0rGUOtFDv37J2ZnDE+
BsTVUU5xXEGDN3vDVFAXwd6RaElVF7lESuaMC89vmhaqmVh3m6gHpWWkB71aUUd2
hqqbFI5AG7zORG8JCz20CcsBd1wmgNeagUCZiqRC5f9QWkU8njXMd1cw/+z17JE5
+ZdTqoAB2YeM3iXNgiRF9i6XIB2iuqlIDk5oAhWMO3rYxkQLBzYcOW4Ol0U6amjt
tLWg6tSdFOVD96nR3fo6/VlO5hQE4//w2Cbh9fidV7LeQnDjm713sOBLOleVm9kY
7/w2DI4vgzFtirHAZmIFO6JRa96CvRnLEs1nBtVZF/0o2rCKAqSxXUX37v9NDInS
L7xP3qmcBgWAb9NfaSRLZ3w/dYodQogSfnIBOC1trCXhaZ0dNiCgzb2AC+HzJwJH
r3Rc/BxbEfcmQyhph5OPVo8La2o9Vmef3OkJbLaIuCAtmmU0Kc0EUbxOWR3gZOd9
csYsq5NRTk8lVC7lq1OSUStLkcMA+wJbAHyX9llwDNiZMH9cwap73QpYumKjabBq
4yeJTVRIdEmhnhqGPiaPbGTIfrZr1fsO44a9AT4335OkrKNfmJyjO4blwmbjSvz0
0GAQz1RTyVQzkHUptNRR0SkDM4nvB3+llDSG/mdhHPsS9W29WPlKYGr3+ah/nO0W
V8nQEoMI9UC6Yc6DY5xFwtn9zK4hL8ws8rmlpwNc7BPSvAJmDlkXfcQe+AuaDxjG
ikO7n+S84va5vG5RyF4c7EcQbdOJKg85KxF6hEA5PHERrJrpULvzfmK4FOFIoFAy
Jo0uz07epWz8dtG0pIo50bzV93bKk3Khydg5KBHfbfZikhWiB/uqZcTKzM7Ssq0U
zId+sJusf92EwQtdYw2JdR4cQe9/96W8q1IBsmaChjoDBWWpHrrqGWws8UxRTqTr
czZQ3+k0Val/+ogcEk1kd9EF+JiISVbmL4DUjnAOX49HI1izs7HZAnVDWPGNRDam
qYq9k0lg5t8B13ZUF1ZuzNjNAiiWt+jFrFKeYKuVpYeZBqGyvZ4HPVln+fqMrg1S
vI7WJsR0fjyfAZv0y4SDg6WB3OfpDafO9M+3oAj/yWsJz41q2MaFBcOzyRP5JvOZ
7qZ2Z71sBr+Tzzte3jv/7TUq36qTH1NWhVEqOgCVXURCi9KteD7QHelMRNDYCY/G
3sgsZfJ3rAsaLTpllQODNeIH00Dfb4li7lzgo6ntqW/mrXwFR0dt9tIXt+vomiKr
VVv+NC0QtlYEO4ngDytYXWX2OHCmBqMWNoC0RoAIV2RsPlWp3OEehUEj8N2CBFam
8/9cPAT0i04DHY2BI2Myh/b1tLJHCxpoS6YVRCFXi6GDm6oXjKT+EBZYmvyXY6vX
d2lbw2wVKINVyFtPL3N8v7Ry8zaalJC9eo75npkH3OZjK9nA9pcthhhPGfyjoptg
5Q8jBRa2ipVrEeYkJ6Gm6LigaR6wDsjV+gAjgXf0fmoyAYgJVpzvWE8Yo2hHymw7
ZfIwNU9MmsBJNLzziEKQuKIdjRywCWB9azernW21KccZFaIeVJSfxv+RJf1+9uMn
Q+QNq+sjf4fVpY6xW2hRDjO59gR3YdFDMUAfw630G1tG+6rNEPTSyK5LyWx3NXpF
b3BUe5qb+WpV1ZJVSigDqXjof14gLUBPTrbBeqFME0VkXTO1+nAhOkh9TrSFbWfL
Vn0ssIWds7rzHvJSpuHCZN4E6duaxGB0GiX25CinmwQwlfnA6Br18gMdgeZc8kpP
ZkBvRj9wMnbLoR+XRqmiJbm37Wutd07tCpeyiQLNR6ftxnqiyXf7e5rIz+Hv+YZN
Y2hfQGnI17DFJTyDnqNdqI9idm32eK0BmA+bv7sFhEVhus2u7UFRSRm6F2W94Y6v
E9cJRT58Nr9MUq8PgzVXo6Mh0b/O+Zh3a/fyLUwkspkdecAfTIfQfwliQYc9csrT
d26RGC02vfs9qnCbt0lU6QcDaX5JmK4VpPVkQr57+TzHlW/pJav+FLfZxBt4SL0w
prrcr+mfy5om0uXMree832fa2kO93Gbz4b47OIfY8+UT/qHHyKqYUTyh3P8Cv3Kg
piivhPo6VHCbO/Xuz2OERDX7UIfeyrjY6tDTqtZqG06KUIoQADDpuztWPKLdlk8c
/M9o/P4TJ6hSvbyhXm9n0hYYk7dxrrI21obc5+zuOEahzl5x1a/r8r+vs/pMAd0b
1looacvjXhQ7CKBpnDeooYSzhaY/mK21iPD6v651+PZZZnC9brZUo1D/Rvcmarjs
P3ArSvTTcLIPQnx+cd2la8JYHDIVfpEaWKN/4+MJLXosHLSghE6x9oAjFkEzXfrv
RE3p5x8q6dtl0ZZs3L84/q8a00VHomipcYcAOmL3jwulV+yqPIawP1pZCOru1J+V
wmYeG1JrD/B+KyWaBqS//Gin7xwnfFTWhg7zDIyR5/JTeC8A76MhGmQvsofDY3Z/
lMMoFTPosBn1i1FI0OIoPT/IZwxeR14Q0e3Zt6xu5xp8o+Hv3IUR/Q2uIc8tJB4+
4TyB6N2MJ0GS6meEJHA/Xacyng3nJT0hxztFJXAl1vhVNJmOzXALG2jH1MinSnQn
mBGl1zQvbNW7XYDeJt8dzbACvd7WcklMDWP/6QvW1ViNOqdUhFGznCusXftPy5uZ
QWbhB00gQtW/WrjFyyfJL05gMr+ubGFx3+ucZ19PjTHQSpTEoz2J0zwBYKYnQw6D
TQnq0g5Q+v8JTmR0Dioe92BaOh7VuJAG7Ma8yXoYf9Cg+OV3kNMO6K7okjR4d4L7
yw3i91UtzuCEDexNZXDVFHNa1pw8dbfgD0x9/fhe/DRteNXozAdylgVvJulcvQ3F
C+CydvuoHkmNf+TpLF7gczk/QvM53JcxU6yYBcEB+ININX6CbiE4zm06sYcE2p5O
uM3dH0k/Xbxc1rkSrJqcSyAFjXh+ms+nl8FSYqsiuyZsgR29QbYjUAJUatAyiyx+
UHV+gkCxpu16JHKYr7WHq+tLE8UUG8mG0f721uPyB9AhzpU5pjaZtCaEEBY3SDST
qQsYDv52YoIShU150gh2v3IVvtWvWd9RfiwnmiAhswdqjzEp5jqRX+cMZTJ5qH5w
2v9l2wIsc3samI5KsFxMf9kggjN+GX5IpTnQHxUL585d/LV2xPttUjJYsCBCc95X
g47kYpzi+OktFA1SG0xe4+9cJxP40+SQMIQRLN+c4AtGXzs0Kjg424o9oUssG+tR
xacDbY1YGgS41S4wtxAU7d2xOchXqatn5hDfxxt/M5+/iWFRV8aLP5zts48du2m+
pbLGyO6D8OmEDjdrKtES5LdAMP7A8H/TUXNTjpOOYVljVSsEChJzjBnyWmxmrfu1
+O3hn69XXv2toMTdgfWAR0fU3HB8hkEW/AAD0FoSwqlHWAiFy7nvALanMR2iZlWV
XuSyNgJOkhnJyN3VIrnHLQ26Fdvoxh9IPQhzcbFUmDaJsi0NjuPC0zi6B7ogAcLd
1iHOrpNMJJL6Em06m1rJfXlPwv3aTppzYcH/n2ZEHSuPYmLA9fo2rTac2wSqiLry
0DpZ0TL10TYPw7QYHct4VSco85n7T0B4qdGJWRGFOspq9mX0juzumxRvPD9txGuR
alB9XW8r0SZSAF9B8mKxP3Itxy0/G4tQqU2MeMcx+LYq1OL1qeBYlLyE0ok3yrDE
23H4yTs/jBwUidq8SYkrb1kbYQwfh1HSbfNRFIP6G859IiXHyd7GN3CzUg504gRK
gL/AOVFLERSRlHJieb94VtlWI/QYNGAFysK7dfM0d/mNDuXH3aUpTcxttOyQGEvw
INmeSy29RSgRk3ht8177dVYDi1QFqqx9U+whrJSdh6lcSOgBP161U/IkxVNBOlV0
WTzxA9yuARto7OTTLbsvd6/LYl5mhOf+OEwMDK/Ga4Voko/j7c1OtCcXZdtFqj6Z
DAijhhVRgH5Vy6GcEnjTzONR3ARXBJoCAzghQJ44e5yW+jW4P5I0UuRzRhP+ssIs
E9Xh6w9ZkHJ3gTeiw8HzOFMmvgA5sgkGYUoCcIVePZrBT+MC84uxGbPsIjR41Xzw
KssRfq4+GGuq1tnE6tao77TXIFZDH/frdA1FYThu8ESbYWtaNZJfYD8zkfVUI1c7
0sw2ElunVpNndDBc+L2OkU4+yjK90dIq0f81AOwhdFTtLQolaadq9v4R1Uk3EPZr
q9aVNCOZJG/AJwybyS7BeS1n+Mqz8XM+P5GAkgseFB84NK9ZOIlyi/zp3zWDN8zp
EuLOsT0MZJN3SlYOcXFbM9F6NQMR/rSNVFpaMaB+YZgGqmHfp32DGmGkaSImSzYO
9yextZS7HpiWMf6cHC+q8ugSr/fs5PgCtXS1Gzs6uOdpUGKoKvKlMUHcunmUZQKz
QaL3PQeh3VY+Vg2fDO0oDnwyGBN29Zg83GRfRNMMN2Kze3eSf0QGPr08cMWN+CPz
O2oWjawbl1JKav7Cw6d4mu3gKhkgzwIvHvZQvGiazvc1lVeX7wgxqjycpmv3CWb/
EvfFZ/1f8a61Wt9oJMPEAqVxzjSeyLybNTeJcn7g7kdmlkUYsvmnzFQRhyAZqc4a
EqLnhx6OO/XgJc7iIkq4HCn+IfuMElOwb+cbVMhKnHFDuiX8Z+alxRkQG6jVChWV
/GEUpUFsA/BYOPSGF4HCO6CsvheuSO5Fq/OR/8s/R29fISkYttolkocjuwPUOt6g
j0IUgQyzQUKSqg3sG3DaLQ2OeSxJD9g+XSx9twwmUZvZjaZDdG3fg7YRzICEKgt3
L6o/5jX+4lhzUnoQsJrf6l30wbHXvsLEEQwYf/ZNz0AWvYHp2ZTFLoEIvhkGL1V/
O1PFzzpE5Q9mDQlmkzFZdF28IvmYoNIRUAW0hXcTZ1Z3lGhN4e1sW24zmWV0cVrn
5uTFW3N26at5RuUUELsd/cYq8+SOX/GdJ+LHd3cIZaJ1KVsvEcjNJ2suQ06DFHab
6RqYALWHp4cXpPk6acA4/LwUtP3ztf4hKtbjioflyYV1QAm4GXaeBHZ4HaKf/G0w
TZpzeA1MNehQRelCKtuN+dnflfB/oPih38phz2Uk6+Q9v+wuiGIkCBu2+1QdA0zk
Itzc047Iv5ADgWV56ikB8ijwxOTmZlf9UMms03sfOpcy+5NsxWjoecVUIsH0L6/v
qXVQjS0KPF0PS9OsgGB0wrA0+oB94D1ilp2dMrooOqRuc6FW/q4FXdRjop6N6lk1
C4Cr+rdAJOM9o00lPDxgRmw4cuaWvWMAHMPZRDNwXVkjDgWel5/4Ue2gj2hJjMf/
Q8E5XhW8Wvw76jaM9az+CxEGwJxaXN27PXzP1UlS3hnmzQwau8t+PJX1mwFb0rvw
F2gFal7bb0iRMUU+8Y9ei3DN5j9RzrqgEKbpCkgIdQIljck4jUQu6YbwyWoV5Hah
TvlYYRL2LSHb+Vdbs5iTFNU1pCt5A3LjLBxJqQEJ4QjE5jOyxg2irYVwAq90YCfv
atJTze5YjOSvC0wY+S7AKvpLXr/KyBhAbSbpjtIMVaDQDO3BRcmmLZ2T8AzOrLlH
KgAaHg71Rm3X/fTxGX5SyiMNO8sIJAvYdHO9TOZUNO6FL2c06E7k9/ujFcYcBH9r
tan6iSoRfxblM2nYyJSRO87Q/yZt1se+X8zzRVRnG9sqycfXFAc5cdfMNXbA/BZD
284eqLD5PWR2DqNGMxTyq0tfuDoDiakEesReJYApLKQ6pyJhU4MZOPcZ0Po61E2W
lPQu5aIrKzxYDBmK8Y+8SVcL7LBS9v0U5n7Tp2nL+4Ck2zDs88Ni2tEvDZF2yXJe
XsGpunANdJaGnFnAcWVlDTsBmTKfMlZJBOj++YL9zZY/IN27QysQMI3uIDisDFiN
C22fMCPKtBi2OBQM5pe4xF0SOlGD5XGRifFwkiSmibp+7l61lB4ccfIg9RENzY1v
FMY7VbfbXytJSAKfe2DbFuBYef0am4Ngl0wwyWPzelMpwo49ldF/MD5XBdQM2fL2
jIUfEzJvoshkVYnMJBDZ5Y9PYa52rDEEpaqwtKFEnc5ELkvWgOruQClVS57ocGNe
HxLSKZHJPsOV9vRBs+YAJTaJwDo74c2iCK658gfbkjk0qCsLN/5cqyXlthRPWHgN
ecvBhZAOyq9tIqgx+q09kTw5Ta0dggk7q4quvXJd3nKlMUTb/dGkEUTeURPDI7o7
x89mIRlsvQWeh+4M7rcHdJrYH5sRGfBv1xP9SzepL1L9L49fLQOIRQ2NckVToW3j
Lt2nuTYCN/dyr1nEPypcSNbUaWmHnFA0JD379pBa7qPIRBpzXc29W0qJ7NgbMYIs
Eqyc2bsaL45xqg2qErP6RAEIEM2a2shjbE/wz65kRuoPhCefpNyHUcTHTZ2ldtja
7SPGsyZJjbjDFfHzdJAIK+lx/IU7/2u1FA4S6EUww05uSaYbPOKaZXfOLvHcOXTW
/s5OrWmTjIbDIZ1V+B7M5JCNnCjp0eHlv2W/thA25ch4Dt692XHVQKuCNEn5/T1s
Fc0dDu9yq9MIND8PWnydS/41XcDQbX7fEmLNyfGdtmN1gp81CX50WPEBDF9DF55y
bfwaM8W7PBk9tlXuz+YcLsIhk2JJlIy+mQmYJ+TnHCs4k2UGRGbr1DH04hmFkiEH
ecq0Ok2kgd1OoP322opqGOb7qzZwC0QDIEDLNwVfUSNae851RgV10aZhxkX4UQ/4
+mO1sOVwqisfY/74HuZBp9stNwZ0xz61ZGCGccQLKACmx+alwcIEfOxR8s6rFJ0K
QYWIc2YakTi2wZMMNdK0d5ehXvbgYvkn2z+uO5T46//LuxGXXtKszvYk0WxW+q2B
qFKFfOf1gSS5wwz8otC1uPs8FrdIi5o6M5ZAxxXQtQol2a5WoIez2wqpN4cU4lNg
W2ocVzLFc3ZAtOm0Fueecf+twZPnG46GF4EIeFS4k9ZnK2qI9W7uYTO54zXx8JOi
lYBzWb9wf80HhQbiB5d8XNEtfVfMH08QfoMGTBtvmKvzSD119jLy9L2Rv6F3zZnA
n7e+ijMkVPNIa35OrypdxibC4DiOKaUxL+dSTDYooccIU4Mxb68nEHnlKl0LsLQo
2zIiRSiJ89WocFCKkxryX/e2OErRoQQ9uwD/2EO27rXYzVRr2rWxgaz/vp3XILXP
o9XNMtrrYV/SOK1nDEe70fkt/tocEDwpCMbV22HhNWEYPIBCKCUG51Wa1IQ/AN3T
fqAPeBuYjLtUoOgiODeUOUFz3ZtDKc0I6kcLTqGMzI3JG1Q9WNwmRcdpUxfTqkV4
gptfzeKAP3oF98TKA4yGiiLjB6x1LzSqd2dUFxD9ovq99BZ3L1y0IQXFeh5B50xb
Z2P9pIjEDYOIZE3+UTWpQYLorfj5355de+hf9dO4XyArDPAqOFkQ1GrOJwuY5L1l
h0EHNNi5q+YyPBKLtitt2a+SYrxAFVMGz2OnJNv50GtOUnn7KJDJ6YM6ezuFHFz6
ZWKOKnRXAygHErqaCTyD4p1medG1ktWP38B4KCYjhT9pmeuPWQY7DENHgL96lgYa
Hf+L8oC4IlporxHfT/fhxhDZ37AsaJ3u962zxvRC8oCX3SehQxlPfKnjXGjHGjSK
zfonIlAafMRG1HgUfRgY1mSogbQqZdrXJQccvfAs7SINl9k5DOlad5kmGRAy0+Ts
OAJaL9ynVQMzmARgmDtxa+wRJBRnmXkLDWWF19wHxWQubVCgYpWnw041wZRGmcVI
iThWxH3Re3KlACEvNYn0Hmu8GC75HQrBcOiqgunENv95VMjBlJdQAtWegL2/FeAw
8jhY3ct43MThS8dJsXZBYumDIGNA7VylvmTavB40DIUYFqQNpW5fpaGcQP2mmoO6
umkAowoLzJwdUFtrDud+zK/ToD1XfvCpZnCy7cfP+AnEpZGUMQWWVBTPaRj3zemD
mNlP9nB+NuhdNmj10H651wYBwaI8orpI1Fp1O/eaZt3SJ0rEcv3yYuyHd0RSZIxI
r9ZmaAmUIXKm/h3airk9HQW4TjO7bkfJK38B4djRakBHi+yz4NMnNmoaVsWP4IxO
860gJjAKEiRLBiJph4TsmhKvFvx5dvLWK0sMjNpIC/lQ2+nSIaCiXibyduMGVdf5
1zwdHHkkAxzZGx3o8Th7DAYwaEondGh+tyfOG5e5wl3Vz11hCalu5d2aUo4XsPRj
WNPFySAaOrGjlUEIXQrT5zkoN91AEV9pcUqRukCtaEZIl4xoQwQFuN09tIp/wxb/
GyDpJ2H3Td/1zXPaOm1IsHhOs3FsDkNHZL+p+HwA2cVXyh8FXTN2nHgdqKz7J0nX
KHtPZTCwo9addgNOudYocAbIvxCOiW/pD/2cZbwg2cKXkHa00sS01h3i2p4n3HmR
i0uwMjuS56vLrzv7zOhplsHumI5iQ/Q5THESPKV3KbWe3KlVfPuGq6T1m4aEHyKf
sqJzd6kr0KH6JO5WCkBt2NLklen3uDzjSojNpfy3A2qRQ1aHOqckdWvzie8CDtsh
h1H/ItA62Nt8JvGOhh7jTD4O0u4fLphFKDYgRbJ4ioSncZ9aycA5vaUU03rtMU/d
rqGw2XbpopRsL+PKweL5xg0bIqw3IMMrdQa+4dWtqFiKXHFFA9vEdBQf8xD/bJDs
mDQoarklDYMd4C0uDV85ednDhrAkE3iByiBKNSDhPRfANkCqCyb9sJMZpuS87dNJ
18GpcJbuhGdYj6oZWyqsPncyBy5YLjIEAkfj/1igK73bpt8XPzxUgMeaU9EVpfRl
vFcUJ0vLoAYnndRYgKVFUj8IeBepWUmSHHT90HHqbj0Ep4SFAhVOms+AYy4IBm7L
vaAuKqG2Ft87Yrsb9U4NmlDBSobgJjUA3zIDm6ygf5a0ZIHokLHi9Ldu31R6gHlz
jAavx5Qj0teQ3nIpr5ZILdyIvf2HO6CtAs8QOA73ClSxLG9KgZuw4XW5xxeECjT7
ssnMtSlOH13ZlHKYB4GqwYU2oUzOX/HSIiMDxVTyJ7d4puJTxHItRut+fU2zTLkI
ZH9WV81UB+ZIBtaM6NvBc+FP7k8SfAcxpnddmgItnLojOJdQUsEq2kdGjPJ+X7y+
DUW/WloFwMPo1omO4pGub958UH+rhHqFa7iIjJa2V/ORDJKSt6vh7MRakcbbnEpX
3uLMlKkGhhx85YWx2P2fOQ0yv21ZPI0wf5ogpn9QZpVggsAXqJ1drAPicmCr4W7R
L0PK7cD5ofiB2Nbc3Wxcd9llxahDq/IhgqYsBSyCaCChV12ObhpmqJmqHyjCbiZ4
E7ASc/xL70+ztgtyOSVHdM/LQp8KhzOiUsk5l3RFC1Fmjo3I1UAVTvyDJbAvV4wF
0Cl0kUwfK2PmFUKH7MmUsjE5XG8BfsBlBJtsKOcVgr9K6aMCmX4lZx0aJutYMOYk
MkfVtXSy1QrGDdLK5POl1Ux7eBlg2H8Ejp5TdeZMtLIWDgHfEcX42qO4pfdg7nNl
BAAy4R8BuV8hI3iB/1mAQ0WD7GTIAXMbX1jHU4KEnkMfWEwN+3O/+NuxdBR6uNqO
uJKiJTe6lVgH2DbJ3wzpr5/x0qK8y+NCR5UHHRuFAOTb9lCzB4wlYgt1uWUe9JFx
4LB9axSjmw0MUgPtM/bbZDbpA4ynsefgVGHJYi9EPHj5KxRJcRI6iGyQTJ/6uo1j
HYZDigVkBhBC8zg5N9I5j/RlB7jKoG+ftjOdU4P2sinDGsbcP5Uv368/ulw3DKFU
N9WG5Gnpxr8vHfACvhcONiTJgcrexxLUAKSXrA1CHrTvy+clIlFYxJqThtgyHhSv
ogAw2C2DG95AYy5+rrOR/2K8PScWT4yudWccAFoDLWefSmEBXKgSfga41SB3B8P2
sFDPOvwQOZVq75dem8/+opLQCJkwqUPTCvN1eIpzSviQko1Q4fj2oPFlCWFfjYsJ
EYxoJ+QLn7TJCsBBVbvQEjC4Hp9HHFwlS1L2Mh5erHlseJgzvU5qkz+qID37XFCx
vCtw0VW38acnSYub88pEajmdVkpCRnJLpRWYMQ9hWIjoGu/1ZY1aYR+ziH8wEqHg
rRk6EwpnxnPiJaNIG/mZHGzuEJ4LF4zTxOmIYgsdJSlVKcMWA1qA7OGILaHDh/5r
Kc2ybVkD0Tr9/eJTIrh3RkUCMhMSUqOkeNDNPxzyCEyAB/0afvgZur/kyoYtYS5K
vU4O+oCX9awcXc0z5LQN5GISJ0PH31F4xOsAVzVmTILkm22yMEDT6Cbk97kb2DZX
Y5/dyGG2f6V2L/45Q2S9xiyTaRgjOIewNt+VjhkkY6Qboc4ad7rhqAJg7quw/B7q
AUyQlNOGpO9H2IPSQcsKVc6p6PV7vIeEdT9difVhDUoK6VjnNFMYLzW/whUb7Vup
wC9jbWdeCP5RDVExiZBBFPm/jtya9oNwu/R2d/QtGEajrAxGJdQ4MNDscYLVMFiU
YOrUVOA3Kb8LVGfaWGQSPPJTq1UV8pUbmmrLjrVKBSc4KMj6m//xosFelhI2qib2
sQ5XLJG16ifgmCPep2mtQGUZGtO3ixQMhAComZlgbmlLpgLHAtMoaQrJQnZJ/PXc
N+nOZ8YTkQPpAlQRVzBmOjHXdZv4C1lj1W7D7gLoKNyObfMFolzMuj4oCjOLrcIK
dpSmgrBb1eTdGDwfB6lfCeGai8U9XvTZTHV3DPvn1jMh79fTtj5ROmXkbVEiD9Bh
x7OnRwhfJ2IgNgBI04WZZKEHvsEtSTQ4z8C3mmwGfFUWJiXfkJBeJXvbLYzr4OTd
M/a4Vn37B56gdyoX/F+GedVy7eqQjYIE4P3DuvBWJmUa68mt19JXR1Egzl/BvYpH
zMvFvfBb1VwcnkkEuQzXEWLV3fDq/hXoYO+02m5AXBm0nc/mSk/9euDnbNX9ka8a
J8LXxpE1UoDZ9QcL9OY7xromZfreZdfWBbzUTDQWwNH4qc1/nVJV5mb3piul7F2c
sIBlBA6Qx+g/P3eLI8kPX6hMH+x72anrm2vkJvRh4n3lknXHP8hP8K3WnBMMHt57
HALdLUHu9XokMSvr5rHX+bbLuPbmOhmyfY8WkpdkD3t61VU5xEXMQXJDhcdIMrCV
pM3sNJX6fJTaeUieuuYFiAsNX1DG8SBe5C0vsK9Ul7xIH7oTCXOvkbRXkxI7FRHf
kvVoa2DKX04PDlN67QhV8QDAsZPLumwSkum0OTBGPiUNOdqGiTj08n22Q0yINKn7
wJtPBNGB099xrfNGO8Isx15bnIvvDAK1203thOBniCXZ6RsE26lsCybAk2ZQp3lj
YZe48KlCZPpBpOArTGP4HDCmxNAHpkzucwMnIedRXcPQFZXZ4ykzGECIH4RnMOYN
BWF4blcFxy7uOdrAJeBYBn4V9QqJjh9CwXIwnHWIG/Ry+lqoPGrY1UY9YHoiSwea
pCDkHg49VReIaCwC06vt1cH8Yad1nymUDPxl7hFEwwxh9U6P8h/yqjmEyPlVhjB6
a7GdHIsBHYzPSwhHxo5oQbOdvfYR/3dRRSRfUh+p1fFyPnFuysSe/gRpJ+JwXNw4
hTtTbADnx18fX24fyPWdaRrtFVGyl33S5FT5Y7iHofbMtD9UM8c1ULIS1MYnnfgZ
FZ3bLv6uRnOvJ9ytDQTNPKyoIl4GA0axJd+b2H7hMDdB1Nd1rGdau8VgmpvSePJL
6GjtI7bc8jmAwFYM2A6YPyLUA2xyG/JtZsTUDwcw6Bipeivyt1+hvtXSIAbU/cUI
76WFkUcOscXd9ZdzHKMiO/eD8OxRKa4Hu/A6XPALyzH5beDkQLeZ4Xz1wV9FLC1X
XAYeqq+KY6sH6YbuS5J5Zmb8tBpEWD8vAsSFRzg+nTf0cAMMeQ9r0T+q/Ww1a+3O
rA8gn5Q9S+a7AzPMujMYfLI6wtsSasuXLeGISoMehLWsuCfPTEgsayTL1Ix4SqGT
zIQ43Vd5vV2An/hG7LcSHDposT7pFmDvbTKV913iQyxWrej2ftMlWwOtimWlxGvv
5Ji5akFeuuQMzPu0zUNlZCHCwkDPaP6kIyyNdws0vLFw8Az4BI+JLAetD0u4JgId
rP5yty4xHUKg6pWKgbxE/iQy/pLawrTYy/v/andPNUmIiqczxuMEvPyixZk/aVwm
MaGTKc2n1oIrwg+TY7ttjdqLZzxUNNLaw5pCNnsCGMmQKyJZchfJlvF574lDjgRq
LDnHsyACv00vWY/gll3iCj19m2wZ5l26bCYEMfHYuUo/Tb20Up+Xe3x4Ib/sSdNw
nT0VrY81Bs4JKh0B79/QbbDVfN5WWj3xXp4AhZ2IWAP6O49ngiq7gMZ6ly+TMqZ3
BJDk4n49P0zZIY1fXi93nUPBlrTKKigmMmLNSCTN2CIYmgGuNd3UhaEOucu2QYth
NZ0Ehg/DL6btoxhT0GFzC5yzR0V7hpSwmqlEuosaK2fEHJVcZBMSNcqNkKodnkHi
jVao1hFmZS1LvasbN1Z3WfLETv8sYaMxkfujQFa/3m8dYaJz/IWI/gO4gvFDYrGc
pm6zOoWAWUgw/Ehg/onUSFGdhZsFaJClsTHiEug1l9Y5p2M+6S7CHJw3PC6Mxt4K
UdBpOlkUaD2SvzyEBEbOfJHKPv4laGKWROfV9SK9zwu2yUxb3ChDHjYUyThj9Enc
gkK/jCdRtG0PBH8UwhPWe46mkEySZ34PJ5BrtJHpD4RmcTAOoyn0rXjmdQmMQA79
ryXA9jhYElXfRD9pmKQ3ac5E7d4x663eTUeRbSRLRaZVyD+l33t/1XugZX7kACpf
wIdulgW0UWpgl0m96HctIpg6eIjs/weAH+Tz+O+vUWsdUyqR4jlaThpl0SWg2bbs
PzTDOibFiZR3gadnujd+k3CMWEtfKyXAck+QFb8F4sNqHVpARIrkCJIvnpZ1StjP
g8RxVEf0/nwS4voSHTpAWMr6bUK62NkECcM1uDk9x5x1lXl8HnINyAsSjOLZuT1X
OwQr6cL7js16bwI66AVka+OrrIJa0f7COYa/XYYdFLOu5WFgxilkuSyeTCU/vVek
Wg1qrprjmL07wSjpPXECtkwsgitC+q5M2lK6oiKW0mW+EjjOjDclQfyGVHI5KIed
sZC6dQEdGjGv8bb2vJNk8P7jrRoY18UmiV+jusB2NOy23CXdqM15pJoOFk7btCwT
z0Wt8/g43/iXuJL5C+ked4HzeZOe8KYX0iR5fxCiEu6LsJT04eEcspeCBRqCQVvb
6A/tPx6X2cRKYscGG9gh1Z3IJKvC9uQ0thlIrZemWw6nsdnpx+FnNo4mEJdkFQEE
wcStKmXnbBxklEC2Ic/ySEGFC3juAQkAk/zUMzTytgsAouutex7snZPGMD257kuh
Qo6754nbHPatXnj4CYZIJugMKKrddfZ6csd0JFAdOyYH5LPZU4TmXhf2aj9f4fqP
ba/guoSUeGQ1d4PFV0touGt+wFhlCfeP7zBzJAq0brXsVkG1/C/j813P8LImbVpC
dvheXguJ1yyHMEkItrqf7fJCYtaSZONjr3q75OwD1lZvhGWXcyWtW/T97UkVvkRC
DsJpCvPZ/TS5DHi+IRGx3tSi0m7GvqGOpC77j5+QRRFqoW4VnvTH8jK8XbNk+szV
oVEjS6O3bvCVzpnZ3VbJSYJUAuzOh1n4rxFULWiTLPop+P3nfsmh43JHl8w4NJd1
1OykSmLVm9i2R0lyQgamcPcpYhAkDUlhH4hiGeCwzjKD7y1U/qN3tCxldRbgAPaK
Q9ORg/YBZ7MTcA+nOV6A/UtOPANc2AbnwVGPQYomE9DW250lMASAgWVWscqiVX07
wDSOUalgcDn1j65FtM5qvBq/rYNyvECtEB6bmwwkifPhtgA+MsSGtY5PHNOBQqPn
02zRnLUA5mkIAqzsh4/vHSBDTD/niqw3BksroXNG3I4q+t7bZYIGjbQcdT+f0a41
kjT6BQnOGV2V5Qiu4MhwqXl4OmQjxf78fgteQwvpds1ZO9cf28PAECfg4jcjEFNP
d/tIdUuqktc3pUWBqvzZYwJ76TwWMB2h3szyLSTipc46IqpymrJLMuVn1PaDFc4j
NwIHxlfZNsRSt5Ma81diqdwx4UvvJ/ofWmAUdNY141Xemp9hu4ErYZjxmJqDyThv
tnpxTxdkTS9z6dwaWeSU//cIZ1NUDDeOnnXuyspNIwNHK7KyKBZ0uuKTmdDco+Da
tMR5eQWne9xUe1cqXTSmGCJE5cuKjOTBANbfPf/xt60Rw+sbmtb04MV+CQ5Ni8kN
O9MfXMlIqIygr0i6EnRVS+EV1RPVriPyUuh54SUMnpFJc+pCQV9IIuv0h+wPTWEQ
V99UYCdcKYptmrRBu7IH7+4T8M4NRlZuIKKc9mgVudiBe0Fepo9h+jNXfzJyKFQS
QpAJDfg3NHi5Q23CpbdubcFtB1WRgnIO+m6AVphxfw7ZztdPY1UVibCcz1O6Q0od
mbEzW0TiNNYWtjSObpxiHZJaqhkshbSnMl0gLVGQ3jUYpf1CppfcbbY1zVqk/0GI
DohdO9Pgb6uHpiIlE/OkemoH/Y9JnOO8pPjGS5Jw/UZXmnDeeKrmCbprbmOXj5XQ
49MlCUEWQG9D3XUTQjq21P2tKwmkUJfroWLOo9tfALk6sFm8pXLWx5hn1ecHI2pt
9t6FuTQui8GR4q1QmNgGvmCjpm5LqwhKQsCa4p+mXakJf5Y5ESiBimXWbyVJhXb/
/0sUadQPVnGzOdsfxw0VoZ7oppJTvwxFPNDczbwmVMW38cveTeNi7x/riEWnaVuz
lHIudSn+dtiJj8FUHaswhg9cYQpZG4xjh3xXauU5QPAtLcsPuL/bmVs1/S3Rn6nk
m+7Za31Hn+Ubu10VkyBQfDcxac2dAr+i7VnnnTa4SkBoElLDHq4JsvCgIX8dd55k
A+36XpcnBVvcAf/li/RZGRIAwii48jXYtxZEGqmXl82gukRSs7dWCG1ljgN5QWa0
RZ2VwP7MDmYrBXd2CdHWyrwiemFNZ3llaX3sAQwKj8DVwHTndxTUmnOa8WfUDpz/
BhkX+nrobCO8vr9yu6A66RwMI83fhR1xLAkNfsXUfsuXCg/5kJrPzjjpDXnMPLOj
WNqxw0SXh5N4JwkWi2S41VV6avatEjBZy36qJulBOXmNxUoGhmJZb9Qx/vsUt0dD
FuH2zH3HTp6h8N29nn2ZWpxASuVhC+w8X4Z8H6leHeaeX6hi7n+XiFWWWnYojFDh
5lvMZrxkQyPooWZpcnmu8G26Z4W9bjCoTRwu0RoQCjZiGIQQZAvhqIBQNmk7BaTR
IhTAbBCbUKU1Hqo+g8WP0m0Nqomb89dxjXZZRDFabqc8QouUVOCzmcXTUCm99UXU
quhgpUSGIL0ltsgWLLwGq7blpTEui+hbyoYIA3wZDEaBOETXwPBWSjMtzOd8bTyy
GEr2qjwbvj/FkqJ0t8TZAd8ritEfNMIGuNglt7norBvk4/yEsOJLg0xCutasognu
gI5LEDGzxOIaIW93G+4eTe9mEb/Psa87eI8MEllApb1mpexlUVYUEZO4+cDeHWCG
e6fGu49Uf0rGx59sW0E1COUG44oO9oxVRdmw8nkWy4FJejcGJ1LC7FRzWjgaWx3o
vhTPzrzyjP52vEjnH72R4OzZcwlKCGK5FXBcWHopCLBN9kjX+L6JRnnFJS0n7d17
uM3bu4dxutckbOFUqzZNeTA5MmLalfP/wA+V7lsVPtjTKwp/EX3Du3yeGENeed5D
EyFn8ayMLaoYjP/DaU0n8pBalUB1D085o0VXAaZr1X0MxxFMWZnP/zndfCew4lgL
jICLkR4qLMdqJCe5SlEr2Sx7HD8ifjvLuVIBXGRlK9Hep5j7sNzkPaSSzYczEmMX
WcgBcngaxCvlq2lwtwUUH0bjvihvd0hCiLTxRygxOZaYF+lFanso6DQQNYJ/xGix
axOl8GWxYsILHwRyY+coyMWj2aygqTM2uNlHDpX5KVA/n5uPqJRmcRGznTYmiDFz
63v3TZQHEn+JA+0u1EITVWqo3iNnuKlUFiINLSm8Nv1gtO0z8J+ublf/e6rnb5n2
uARdEJu8jD15PvZV66JtXgMBGAIjpf+NFo8kdrbOvoOvYvjmYlhZ8KPzo4d31Nd7
Lw9wdcrUr+cJfuQt28Au7vezBVxpdU9LRN1K1gDZt2COaC5L3luJDcOaSck56BRc
H3ZOiG1dWqy3vKcue9NGPmShh1ARb5VQkl8exoSF3feJH1zE4TlWyQdNSb0Xv7IN
X0WWXIIfmbxW8Muc6gyo/AAQdGzOxs8HZ9jFVJ+HCPdPR4/hii4EdC4vNfgBN9xu
IE2aShoP3/25rLvIDkBDC/ehzb08HRv68CvJm372g21cH4O81S7C20DUT4MaSduX
Ov1TTyG6cHGpqSsosepeHN5qNAXjxC9N5SjvEnOS1OtMjiIHDiukMezrp2oZ6l+j
LF9/0ARK5CuYsF1YWg/kNwfrqht6v018HOW/2dbRfpl7kXTgCAG6KrmfByGNe4l3
lO7E95TVyZpSxGjkzIVIeyGbS7Xs+hrrVqHDsbxMR5+WKHMFbQbiqBAXngU6OSce
oh9n6FUDrpWn9lkLkkKTlEqD/VdFn8h1xQElamw/YuCjcCrl7N0szGeFoFip0+S6
LpmTOKSwXF/0mw7grc0OMCrDR0WxKuBi7yspYXsa9GGLCqP6Wsj2yPq7S/goMpiw
BVqCjAsMlvco9G9VRX4azHAWipg+ge3s2mS7DnCNUCxn69PuYAkt1I5xskzEikKA
UHy/fHn8VlpWMbICcs7dQ6pdVFCIhbjpi8VrjMs38drfoMclOpxgdHEc9uXdJbD5
WYGFP4GlUUnVjVPBR91c5KHbxii3nUNlQ41TXSnUe1jYg38eCv7SeCcFak4HZob5
jVa5egnISXIwoX7bqj/1IvxlK/Zn1XHhulAAvFwiljzK5NXpYYVo6H8XTOBeElHZ
mNQgDM6hixzeXiSH9hZ5gsG990M+Rr/yBGTh++Ay3Nmzfb0UlK6cGOYMkt0XcRwI
xJzeED9M3hr1gFFU8ULl/rUfRxckGHVY7SWpzU/jcaWim+5/5WCKM7Ay+mpwz3e8
V8Y7yS2xaCiGy3371umE8NJWc15jE5nycnT/ZRPxKhTFlbVAWAvgWYKvI8N22dgL
AjoQFZn6fTwZEXyHDRS4FwGh9NXLRt4JICUETGXEm38AKVTpOAxPY42PWeT9MpuD
I6sAb0oasuc+P7UZix5CdHBGDm4zkRnhXDvpvNo5Q7iXooAnVXoICt9+8urovR6h
aYd8FKP++oqgYHd8adFY+kRQFz7BpH+iW430bYEmDuTjhPQsKjApe6FzKAqyhE0o
h6p7BkPJv0GEqSvpU7uCZcvMkVTzrZ/F2kt5RqlcwzTl/DzCY5XhUt/xvwIDkGte
XyiK6s6YyntvbqB2FjH4YurfFmPAaOhtgQR1CwwITEUx/iUtIDeBVC4ZqG45nMNG
xi2YrDM9u1xMKyjNQDfwgIjVwrTnvfoyetGvznoDVICaVoz51m5mdJkrdwBnf1V8
W/303SUJtTX2lvzr/EmHmnquDVFz8ynJlFeIvPw2IYHKCaRc3HclkGGa9Sgwstl1
Ig3xUFOAQOKYtTBIkaOaSct6gVFGrVBcETbxZK0vAzGZAIexA3yaCw45lHEfn8yc
U49IcBLTUsBom6HiQek7TacXHCFFGGiVBfl+pCsCcj4dUHRyT2by22NUEDuy+N8D
+PaIS0NRJl4GbwJ0HZpemJTL+kDwcAtIKt2WVnmafQvV7csDvHUMhVnB2N5A4V5r
EGyFbOJppP7Vlb8oYBAatIH40yaI4M0T2Kti1N7xAGt4ipVg0D1Fc8bm8v7essKJ
nlI5fq8HnGQNgzj3KXegETZSuOkhgqR076qIHku8jP9ykqbPcQ2ZAUwbr94GAE9a
4AX6F2dKvKpPJtRD0ownaShUoOwkdD1Gx0RZtEA3SaU3qAPf5T65H17E/mXCZwau
KMaFSbZZR8ST2J0fmpURVdAkto40y9yAhbnA4YJFgzLxSsA320OxEE2E667N8Ia6
Vn3pJt9rpCDVNLl6z8ZljF0qBE4Q9rgEyNmvZzdFLxaWpt0IT17rnnElVBq88Y8A
QQpkZ6VMokxwxXzWyEfnQZM5fhCisBw9c2cAOdDfxuFAWhxsPgOa89DxYhT5kaEj
V3kbTSspngSjLHaTMMltOfKIGg4dR3mc0fBZUjDE16tvk6FxakB+0KAYyZmwNo2s
EWgRYmRXrG2FVJXciSTTqJMSvb5H3Wyi/2L31XRKhL1LwaX/LGN3RPV2jKnEBVbV
K01yGSozySt5+N8Qp5RlKWSrM8ytY0eBxvzcmNO+FOe9fUwey7D+7JIiqu+4Z3QT
dSQPE/yrArCdc1zzUI2XAHhufjIJ0zFqxZyDzUIHhB5p84mNEyGD4yWDYFeV8R7E
3OAeaj6ZxW6rBJz+Q9YA/6d21N42u6nsOwJMIsxN7Zi4eSEwPxYvMhME1KkfpztT
QWmrx60rCpFijlG89Hi6HDjNRXCw5A1ugr+xlIL5c0niKUmccQTJX7gbxJxHShnt
Ky7vo8ijZELeymhqRsxj6YVP4J+WfdczsyJBU+wydLrD1pZmHFumYvyJm6j/sKG8
iv/uNHpfCuRDXgSRk/rY/mKA5OqgXlvXKv6gDEbfYoCfbG849Tdb6ne9B5cKOJ07
Crw6gAVM9Pfpm7iOiiAw78aGdPMdxFAiQsk11J5t7+S+e2FWyp2viOwYl2ASeQkb
tL7pLrSn6q+vidLNWQICyUcYX++DB4C4JQGb5D2fd4YNeY8tjFuDDUG+hZ3a2hBa
eL9lTHJyTfZRFxTWoaGiEI/+MKEfaZ0dKPz3doxB5cW3g3t9OULE0gV9FBV/Nunz
pp7rDKdnlKjFCJZs3SPa5hffM/JcID88dm5oV55CNtZoN88QHDlAKu5V+NeLC8qf
4mw364NNLqt2ah6Z+VUOS1BORcxJhdZWp6f4QCognznMT1V5jVmD2xX5cIAxISGE
HuFIjuaHCA1UnF73768/jnaMFcAgKIBxUQlmmw3w0C2xarDieGpdVxqBYhx02/kS
C1Kj/DHko63lmu1psfZBL+DL9enH8X2EXZCRVHZwNDyLxrLeyIcoDRjFnnH4y9zY
3mjBkkCU4/DHd1J8322VpJxaMP2tvQWaPtua+akjibr4bwvye0M/f+D9uXB6S4Wx
lmXJOX+cIa1Pq5/MTHwtUmE/u8LBNvN8yOxLyfGm+QkbDMPkUIVSKVnQaNGSgYUc
5MTPhfbX+hXDCFOnnbDOdcS0VRXmEXA7BOKmBN82hpcKmUXi2G00Ev+ncmuj1085
y8Nofd0hAgDLd+XNyj4k+Tf4CXn1lDhhBa50R6Et+kwe5YCiAlAsZQBz4dHTtTJw
GAyHu01HhRSzahPDf5YQqB2W2F4pIx/pgzQf1aMW1xUWWjSkGIlHXOEImaUiDRht
K9E/CZEY7wG3hytjV0Y3tTaZRQ04wzHTP4lOrQSDzOlulBsxkec5ZYOWuKDE394B
LdnauK+x77NKVzOGe47P7nj8ISkkCv13jDpc9nxhU/dzSr+fT+vkI65td9Jy3o4l
AY1N8Kggbmac8SqIwQ80ZZYja9e5c6F5VUToOPYjcsTI1ovu+f2SxlBE5EXryRqW
llDloxCy3k6zSffrcJGxGnDIyEVxX4fnmqNSU/fILo1kDKMYuqJ5tyfNygfonq7m
N9npUmNCRh4drhUDjZzGjPjcQNJy82zcEOuLxPMu8wyW5mAiW2INFYxZ9sxMzUdN
dQz99P8ZdFdaZpI+Wbpj7/TVzlAqP+qSUhocfVUkovWvr0JxSfhbesKpuWBjRhQT
rlMtjpmCBZe9/a/hEUw85smdwmQV+htgudlgO05vKhxGNTBA+QQQCggXUidUGwsW
Z4NgKZ6Jk8Ipw3c2ST7usz36hEKQ1D1J+mUbWKyLagti3P27NhTgTDIcumlAuRKE
I9zOz3QXpAS3GRiJDdTKVR19zPVSDAKt/fuqEYHoSdnRjN/e9fTrzDE/kJqmVeDo
p2QVNXunwAXwu5LNk3W2nMCzIPRzgq34z56QaQQHD1Jwj6p51n6OhmHlYe2w/YkU
7gVI1czrMSLzIUXTn0K6gY+Wv2VdVNQ/JQSixrLO2w07tO55L4jDVuiOHTNXLL/0
xKWIZYhUM8yc7qRT/kdXggGiTuTKrzNwjCfesjcGp5WRSw4v9G3pQbZdXPEHY9Ar
V0LlfgYM9V/uMHsMYr1Y7XudVS3trTqlNdUJWmrqSjeS0mr5/1mtd2RWV2YEinx3
2W4hqFw2oewwq5UwiwLHB2h11+r6UPnwTvPT0X3Si1Yk008x++UhW5y1Fw+MFYQZ
5SO71yaYdApHynJ6zKMOoqhEYLyQFzdSNiP/sO3kekaeLQ8i/BrpXVJf1XUaMvJ+
PypfMaQCIMXxIKfClSFc+sRPzHHB6Xfh9DJ9KSp6SKH5xXo9rEM61LZaXBin9Gci
aMnZcmhuChKcEq0/rNwHER7ijnGYvG2nvi0ODuABIv/NriaIif4hJF/+itYy/d+m
HQP3MvkiLmuJwLFLX4PkvTLKpUVfWyq0wDoWg1cTtQdQSA/DOzHqs0UoQIi0i51H
u4Hgdgva995HXQlxkS0W3MKHmKQBABSvg3UdVGOHEOmyev8JiBhsqgVZdvAFL0wr
nW9hGr4JwLQBYw7vzB1s26rIILvfOF4wp2BqoPsC648VT1lnGVdK7O72fhTvjALs
dlnnl3598Cg1A6TuyFncCH2vONPlwjaXP1iCj7qeXt+ANC4WauBK9JxcC2J6DhTN
NmEZ3FTmEcE1Yh2SC1U0DJNXt69GWWMsV++5wrzgl+LoVuWrKpkUQhKEL7fdblS0
FZBNN5nViJ02fsjfWGydANMP462HY/ERWVIq3/4079HYJg062a7HmOzfr0ucpNOV
HL3JmFxBnWPYA/l8iGWPnfPgefi9z5sIXc+FpsanVLzrIpUlqZNH5KoycWJT9zBl
eNgHgSo6IfYyAM0afuh20JfVzau+kiNb7V82KsMDx0VAan+FCKk/pbSdTkcxCh4c
qWBsRd6YvG+1nHyU8+eWvfpRHZBvqWeQbMPwIs9fxWh71P/ggXRepmoeI7tcj4Yn
db44++3GFDmsCLWkzxWZRmN5lr5h99Oak9440ws36Vx7ukcTAP907aBk4vBmmDtM
f7I91PbLR1jsSb64/NcU88t4Dxt8auKZZvqCrZBimNcloIuGFS+BJ4cA4ZzSmrFa
KBqqjFhRpFsSj9rS0RDuuM6XSLLCe1NBCCzizLIncJQmtUvArQY7gso3I0kHKfU4
g3VxtCSrWMh6EfntKuCLGAbSACOkEpid3rqH0vVjNHUmMJy1QVPU9XhRyLfyWVq+
W4xQCzqJk9FRPzZxqGcRusvf/Tjft0hhf1elxgzeyY9bzGQU4cEeO88rFasV/x88
irCrv6/VtltC6jbpnS7JSQB9Q3brLOGkoUKEpK0B2HvnRFMr0gtN7pPgHK/M+k5O
n2RSzkzRAhCMLZCi1eRxYiH+T+Rs4DK0EMD5O6vt5JZoQjTgvAKRkVuipdUhC4rR
bZYLedk36YO/X8e0ymcjMaX3GADySOCH3HLT5lvOqQrOVvpjHVMZU2+NtFr48bkL
/K+ZzT76+tWhtphnvudg77WrzwNu9l9evohTf0QKqDVRBawY2Jp9+GYrXe4AOHfA
DBkjARbwOTjYMoL8MUw+ghX5vYlm6Jj10wo+7IGDXkqIJCrftUCLikpLfJVHDdJU
fJoRtnuq5Ar+/GfuLUKk3dMmy6affy1etWIHMzrqpFPT3ihYPfrZvKtsjzBbTLWG
Yd5P4AF+2lOC+ySXx28PTTVgaInE+8IXIs/C0iDd18aL8d8IleOuydzX0qvOiX6L
QA5myFWSDBIv3ttNs0PPqrxYI/oCj9SrJwv/xYtwZ9WrhmZaJze2DKw5wWfJdMhg
6wfSA+UbBIPiJYWPMYuVZjIKg3m3W2a4IsVM+bu7napVoU/aefAGPdWignsEQ2Qf
mzniIHJkOTimlDr/JSQXNnfYKo5+vrzeS4IPS/Xh3FVnXxbVTunNxf0OezHEFBiU
9fOkL+unFLNA7eNcIg8PdYHl8CrjMefiYsz3NoQzWCvXglTxZC7wWyuIvYlYqX29
kHKtFqHJWDpuYXtruaZspE9F+2t905ALs8hFA64blcoaFwaFc+UKff1erMMA23P3
VzsDWxBpXz1r1ElyStdO8kn/Qc8cZeorHMII6icUP6pQ1svyBmE3+Y5SUM1dWJNb
VlAxnp5tB2kBoPecPCN+ljg/Dk8qWTiDo7Nc03fr7WobpvoFAZhlm8EjNaPck9JO
0NrttW7xL2FVLbnww2rpw9q++3ghO/570Idy2+4kOe/xfaEXbr2KuZwszy7aO4FI
1ij8JWeQzj29ywHg2pEyidd4UInz18jq6oNOQLdBbCivrO7qz4BuSLQwb51Y6KgM
mT7Qa8hs1Sxk0Ud+FwhwJU1gDtoDosPLC1mY3THQhW/LzmZVo0FxMD9Tl6aeFKtm
JSKdr9CHHAzl2zDmABQn1FrkC19nMN2i/ZyW65CJcpdvlSq4eEBSf7p76R1RfNcl
6YhdcxJcvG1tJqPrFcv5h3B14NY4GXaifeQLEHwqsAhdFPOiiHNNHxH6vdJr+6S/
MaBOaXWreTJ9EwLlzmm+YKyflGnc927t27EHNvkVC1SXZ5yWH2+v6txdBuzdYM4+
8xoGsoErVTxCe8rrWOThnXCHd1XB4zGsZa0KoMiG+a87EN9bVwSk9gzIvRS8toQz
NSQWyBykzjTh4vRLTRjpcojrpRraAojqNw63J7Cwxk7ORTUzqVV/lPGUIkuBTJgX
+5mkSqf6cLgNdyX1sGvJ0c29pOkgNiPE7ynLVoVnbuKPeV1e/OA2p8QxrBmQF8ny
FtpbKxd3lca4YSnfAoXhmRXbbx7iW4e4kylCxYIxYhTN5nxat/YRMMBqhojV7kfO
h9jO2nAw+HRuDYITWJ1Sq8LrJ+XJjHtnFRvcTVP6dCko+NDh9kcOsnrek7z2FKx4
9ASbl9EUIlqistjIQzxAtl8wKqqz6E0Tot6isp/A+DTEtFigMN3gcFh+V+TQmxAJ
Hne7SjOrvx42nB4wMo8azvrpPapX5gnxZt23FfpTXaOOZIb+jvYR9aqYb+adg5XX
AuUnPeLEzViB0jLJ2UpUkA0JEfZ/vCwrctbXPWp9JGU1QtL3CjdGnQG4CR49QvwR
pIyko1V3IRKZRWE5hh7A5en0S4oIA0GqFs6l1MFjvsblC2j0Xnr3VnFqd6cAvQal
zdHCO68QAMMjDLKVOtceQ2c3YFmIuQneqMgOMmrqy1FPn3AWTT+T1EEaOHT7HCfV
2td6+dIgr6vntrXvNkU7YcqRJOM5XmzeMHUfw4bYcmmrPbxJZjbXJcLU/8DwL+xr
1Y2Z/W3TLHX3hUC59LUBwmToPx2NvSu8UXEbWv99cuy0eo26iXYUWrcB9Kkxr0Kk
7DksUftTWLkCIj1Zhea69P1vEylSqS0gWxsXgDfEW8/CQPyOWnKc/MJA8/wqk7WO
SqSb55vOTFbVOlEjDGPrAM0NQ+XCmDbny+gdNmtkjC0DVCAl375l50xuzAUjXEyi
P6x9sUyo1351wBHthC3UxErCodMbWc/YfAQFaS8+r+Jz+vtS7qX1W+kdIhwg8HKb
KNumbIM9vsJSWpz4K3kyBP48Y138FGUQ4bKqZ1AH4WvreCarrDuZw3mNTgWaNrmv
22FDJbjUdVSkFz5IatrQYKQ8qMKMn4/1ZVRuK/YU4I3mL276wvsCpLPNXDRSG1kx
YpPAw1ZLjmYBojx+rAqWUZ/jwY+FtqHAHXEy2uM32WdgDGkataTUH2RIAxbjW5zo
0CpkYRwO7yTp6uhRbqpcoP4z8m6IGzIdHC/Bu9guEINb/rU92+/0MSFBeFr3J5pw
xC3NKDv10fR0qA2eO3/NJilR4RjB2rp33OX56Pdtu+wkL+K9zbbQSfUOTtc6v5g6
tnJ6RfqOKIZzY2cnJwSqGHN9qvjrEm4EujcYtVUP7k/49ZeyZdV0hzbhAq1jhRPY
zev1msQyqtJE+wItyYJNpRYV6ideZy6RW0B99DSCpkxN2+iIpvUAvy9YQA+9hKKQ
Jtn1jz6GuZlVWaHl4VLx/WrW6jU0ORIc+tC6q/w2Jie+Q1ij7/FoYGKwEl8ebdBU
C8NMBOxCHSIwoxB0DCupLSvcQ+GI4msTYYHkYfoQGXC/woKfYKRrAaoMKS8y/cMo
evJZDy7PsqwgEwscTFcF8alR8n3cr/1spyfC6NEvs8OD6Ho8ol2ytmmyYyvJQuwh
ardJvLmMfzwSbtDA/YB1Ft8HM/Rn+wfMv5OCGSl8EswKa6caVYQOPgXDmMdX7nO2
v+MBF73R0885NAv8lJHTaWW3MCUeQX4x5GXeEDCmTlvrLu8jkPlXXSI+PDPq/QMI
L+teHUXRX814YCztYDQzsHom/5empPdjPjIdy8exlqpEahSKJ/WWJ8AqJyzePOaG
4QimmB0iA5UOFudPmcWYUOIm6/cgFlb9V6YKuxxhKUMIVCslNtddjvaHamfA2pKR
nKvn3i9E+lfOm5HDCFKQM8H4jNaM6Ziarv6SFkrNj318lCiVppUOiV+m8e4jQ9PV
0oZECbfF/GlyWXUoMoAoX6A3IvbzMK6oSclzwP+czr5ybgQJPdiNz2bGwSPYNpXv
Tu2957+qE4Y/gTKc/F1JU2A/q5HFfdBYEfNbjPE89SioupyPM0K54GOpyeo65CwY
iZhEqZkul2x9QNvum9g5MIWKRXp0Kg3TblvQH/N+dClCWsGeEY5P2WsgaPmPIDH4
wTy8VUxRIUVcbjCaxflHFt1Xsg95wajRp1F0XVBiwomzLwBnGepukg+mu9JCEGRp
iEDTYcakCO7Y8MBw39ORMvil2i6tJAnsLI5zmwW+FzHeROwjRUifeGXmVmy9ABG3
/xHuNVOP80WRwa5llNQqPHiYsvkG62zPgoXPNWpWdPWHl9DLwzSoaVc3zumgdPfq
MSALRgfoC5DMqkcZ7RcIlKAKULO3G8Zwkh566GjDIMQsnucagOZHNYhlD6M1VeTO
63C3DltHLlmoK/OzKO8nKVFCWLfL9F52EYVx0Hmqy6gLS4bEgDltPsDm037Onotl
kreeW/ZrCvEeE1OGFGbXz1ECSwdUQDKYhm1wHmaKV2kGtfTcrsyB0yv/Tyoa1sfG
abPMHu1YdePSRtT/rwhD4UK6ZZ+e5f7PQh8oErHOMwkVZsAUzVMIwb4bgG8wxojp
gjM7SL11Jbf0aCIu4L8izMwBZaeJxVIyVW2cGJXV7NkSBVf6xVW7CP/8fekeW4jj
1a5zsObc/53m26IxsVcGtQ6rL+IhPCIIPew50l6Pp+cgy57egdtEmueIzG/W2PgO
`pragma protect end_protected
