// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aUOMJp9/1VvDYffMAGIHCZuKgnYt4X9uu87GBfX9kjyI3akZmG3Cbg5ayPEYaWCZ
AVtOVtnq9DAUIv8e2aHoEmAOjC3bnR8v07f34rSMyuEEn2UYSUFti0ydz+RdlOhT
UeAq6KH1OeVCQC8RYu5JSDQ8A0Ka2sD0Xx/1bsWtuRI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 193872)
RX74L90YXyT4uktnxdjze9bxnFEbmMBGauvAXwCgXU/lkU2nnEWPgZ8bFPOFc1Sy
T53k158FdQ+1kWT1l9R3LhR3aoTCrCUdlbaMAFEuUNhzRxxPHd9On2KRRmRua/L1
4WVOVODYAltzwoIgdWSsahbK6A6GYJUZL3QETjbHj7hwKu4MOY2Uc+VMemXANM/w
cUJfcSmChiWmSBgRVtg4FeVB6twiQ2QUZmzxc/3xZJ1vkeTgKkoOPN/DaZ6xFQK+
JdsrBAaXDDXhzsj5wlDgvC9+YJDZsw2+J4UC8V+5eQER0mPP9Ols1WnrmSe1TGw4
5B3/8e7gozcPwl/ZRdVy8nA7HHELWVYKIU9tydA0HNASIZwxM7DKNiqAK2gA98Xr
6mkiA6jKHH2L4JrjF3x3EIQPKDjCmYWZZy2Sej8yrxI+8aACHkAVUIUPWH1QoD2Q
pDXJrvKW9wSpomV/tfRga8Gh2uZ2M4mLr/NKK30RlKHHGCjEzGf8uPOItcYN0Vxs
3/ty8yOBJkxn67IfU9NvUIbeEVZq1TQkfQ2Vzs9ieeK76Ym7qlbxYFkrpEpjq80c
mqgep3QDsxVa8JayJDuNGWJnCDkkwFzslZIXCkYdhkF/iLCXIxZ4L5uyjVM+KDHr
azGYVGCllekwwJzasy/QENWkPGAudDyXE4vhrXleVjnksuBj/nw9SE+p3RFgMqLi
4LOxn6146QD9wbuRCdzgD6x2S0rdeWWqd1VpddauisHrO3nOU807Yp5BDe+oNp20
7TqAtOFekDRhETJdHNoA5uHIRG8+n1yfZlrajE+lFfdwpR3GSAXOmNYUvHd152ba
k3hpwezis3RFp9Sb0azifvXlDofSvsV5gARocaYd9LVLrsT+wEU4utnom5yNFeqw
Ll+/x6qC+coLIiJiTvzc52SRKimQ/5eMYQ6Ak6fbnTc24XVELIrl9j2E3aN87AEW
p/uARN6DfJAq2XxonIaU4pnj6lnGtxbDHlYKOTcmF1c7wCRewrt0qbvXpK8aywRA
AWMI4IT7WsYDZJGy8f95vY3Pka0wlk2TCVcYkZ1vfhukSoS5f+3Lnd55vilw3hML
YOX8zYfRN0+5IgcPiEiPPqS3VSC85p1Q14MfMO+BEH+ZjnowMJeTFQnvwdT9FsQa
yrWC8N2ZbmgdmZrGbbeSUzhPNeqZlKQ/A8ho7Ahc54+gTTsVIYcuqzX0VtUHp3zy
yKUZoPJ5Z6dZSeoV0/3ZehHNZtshS52wRJB8micuQr97r8+hGie/207iL0z/bCF3
yPnK5bqGuBM5/qwcwXLJXwrIny5Mrt9ngS56imN6XDEZdbZ2sVfIUOmSQ/mLtWW2
6F/KMmzdqQh/iyaKNxz2HteIBtEDmGSSGFPcmoaS+waSimiYBcgdmV9IhF2nezgS
WwSuBqaJX21TM27jyXgJbvS5+lBbiI8JTEfjR9Goof8wWIx+xWMiNDSJnBBImxN6
399IGBX/Cwh9zlzuDvznhs9apiYJutjnhPY+tIfDdQAvKSKNKgjC3EqQ06/xxUQF
v4OLOZyFycm9LzH+EPjW8RDtTQ1/1P4WrarZp6xXyj55YMre5uCbSgmTVkzhBVh8
a7yEEsCPgXoYHn86lfg9lxNp5lN5H8vq43DGRqcFWl4R/yaVumxgQe29nORqmZhD
NMMPyw87ENfcpE9OpphJL9Fyc9SgQdT9JAqr3NK5Da0M4Djlxj65KqRbJVXZDBI4
o5dE15KTQbXalhxKwgtdom2wKNFSj5KpcqyEV2XLyxtV4x+trc81DGB19TAU9jKZ
efqohRIrZ38z/y2GcatWWHlQHENlvQkkR1wbPRcnFknIUpj4qFuizyR5yw3e/fBz
YbufaClJmrO2Irbdr7AbVswF2ql92Q9kLLoD3wT5ax5sW9j6kmDGqiSBo4RZS+qj
Y21tpDbXly8phCWOEGMB0Sc9Xv1xxDNB9mGuk9fxLVWAmtzVU4Y0vFquL9X1bcof
GD+uhWLqa7K4jqy5zLkxcUVnUQ8kadmBrPDqHGhupybpWrOid++pNDGIkP8TamA5
3en+S2PoEzQUb9kc7FD2uT4I+iFmrXrziKLPWtUd+q0fQiy0ROZzTl7ZPbChQDVa
N7P+yaQIrwVrTD5/IO96jYBZrxjmLo4+czcJiud8fWntC+XvsyZ0Cw3tvzL/Cewa
xKREH+Dz3ySB7tx6/QxkvaGQG0TnUdCChNEOJ7YUPIai1wslB5BoB0dQNl7NHvZI
O9gfxHNgIQ+9oj7I53JjcxLR3Uc9ltN/cKmFqNMnbv77D3jZ2a98O4xnuxahKtd8
Wen44etO7/lfi2UGXZ6o3orvSSwdwmIS7AUuQuxHkjdN83RGxc+K6THP2NNrTNRx
x/uxt3GiCUQKXb1FGD7j68uFbFtkTZeykI+i8vNQbtlPFzotfmAenKwzkVT+Wu1N
BqfcmZ2bGLz6o7smMlOOT41xox5D3yc7BvedQRD6i81ABGoXJZvy7MsI/uLXdCNY
DnZ9oTGw6UIFWYxG7hh2z1PilSZ19FlGsL5PnNRZ0s8w38jIkpYv4o6jY+xzrpIq
qHSMWkkhGyLQ3SkxA4EGUxN8+5DpTVPVU4ezojMg6so5H6I7ueRr2oL54lRK3C5z
KWYzsHf2hLTdf2DVERTQ8d7sB6MCm38phpZLAk7SK5pNd9xLpV5YCXOIyjiOnFNi
lc5QYC4+ge6Z5BTMD9qNRe/UvI138sjH8qT0Hocbi8a9V9G91obS2w9OjeDYGPQ8
alPL9VUrdBk6E4DW0rNVS8J+f47q2nilx2sSXj4BOUQKrRa/KCOZF+MNjU+gQQ+J
CX7wC6be4W56u8HKnumggDYb9eAexncezLFNnSDe2rb3CYXWL+pWvNIIJuhgEC0D
Ch02t85YYGxeZg1UDpriJ5/8i9gu42dHd4Nwi3J9eWHkSP0mQFD4Bi9Z1WjtBppJ
0d+aTNrBp35+jsT11mWrLPqmqkpqXjs3vZFBMLmoTg0GHmw/zB8wJuqSbNK0TPUQ
T0T/N2Ttep7sc/GEvVjHqCbtTQ1c6Bzhsax86qCdTUzjiiVEv2D/HOumHZsE3kBu
ISW65uGsUNk6Yq+My+2IwTFtHvoOcUCNT22rHuxbqBCjMBmchcRmR5PXzLGu2j8A
kZVdP8WmneXfezYVbSup1RYlutb9rlnKxfWykerumbnhmQ59I8xq8XZp9pmWGnCq
A+43lQroLU3JpTOM9C7lHozsoc4w65L3MhOcZAVh4p6s7tej4J84yiHUvNvbwM7j
WvjaikUMX8qW/XWcFFWGdVUo2w1Wn0zD4HjEQ4vz++4pzMLVapzS69EUF7Sl6gBk
g7HexBWMhZYt2zzqI1NQSnzP8+fgj7MkePlIS0xVvVkvvegSDVSZ4kP/onFhT8Pw
ueqj5FDueImtx71W8XGiaat3oQlwQKQI4sYq6+sgAUo0KXdKpTLb4FRg+le9vCjA
ubFCffgIZBFVV18Q9yrmf/9TDMqbZs2XjccjZaB+mj0zOmIKN8VGiiXFgK4luNKS
/1Dk3NbrTin2/hH+Z8ggRkmMTxrC2FCfjxM/MJeHPDM7WEzj61WJYIUShPh6zVrm
LY1GPTVwoIV85LHj/dSbJwPzPImxGH6AVf3weUF8mAHCMOeRHOYKjqtMpXnqBHEG
Y4NlXzEuo+bKHsw21YqaYKENLQmUMW6nCcckOJ7bVfVPdsbni73BPSbCIKWxZaxn
Ree2xmbQvw4axbQe5xORYdBL+UCfojfkBgC+DIcDW/i/JqDl3UGP6BYYBjPF/xjp
cirYm6MZZK+H+vogU2mQns+t3ulUEQX4o+qFeIkHp5ZR6Ve6xW6s0cCOTarn2eds
eLj5+Dp443zDtibZaDY4NmL5KAmTzQNttnfCwWA/nwBEQMEDPj1dDqfF9k9xZule
yc0iPcLkIhKV8zjOVRiDOLlEhkgIB5n0J6Clm/JD4ulkBAtx50gUgKGIBTXODbI5
hXgxSMdjmw6Y7Z/VF1hgqo5Hc59D0n9wXxv6DU9C474lsyr81j38iP23Ph+Sq+g+
YOli95Dbq1FAOTdzBlgTw16xzXKWNMIcyzZoUIj6pKZ1/QIlWRrtDUaCo243AdDN
yKF+DOTFLmckzWfLuWmNbUdK4GcxGP036vbW5FgCqPymFwKEAydjR2eYzzbCrOt3
XdMwckGcXgIifA8ueSfi994osdziTaWdJYMnoElLbNfIaCfraYQa6jJ7l9LEO9pl
mSol2wC7U8xsLigwmB1eJ6CwzAApOwX9BFJ3l7zgPiwOERKzf5tWwJcDdeuY9ckL
gK0Dq5id9pGX5uyF6u+Ql1KUN45bHDTDHyUW+3dN6YDQJF8EXun190y5O6Zy6Pee
Njqt+lJkyXL9hqxWwHwkCbGnmHPdIyHrh+g9oNHSh6wcjVyLOm3lcILVjVbkgXYJ
jatwxOvlByFN0oNLDVS31DiiQAs1zemn8/lD3Vwi9bvJncUi17zjVjw5W02IFgDu
gh8HzGXfqE+DGHp86ttbhcjLuzYyb8cd7rQNywZhVulRB+/MyCiKQ9mOS1PhJx8L
vJBexCBSKOIVgotX4hFWSGVGA1+l7sLIFkMhDhIs5c1wPOC8ZxjpHSBoVxj4O1Qj
hwMmdfTxoqtyMCnoeFo+XpzO4P7W69tZMg4JrHfZHzHLWYiDfrLzFVtvK14fEByg
Z5p46X8x1OpaD8WUyIbkZXvyN/GMnrf2mURIG10WPUaU6WA7D03ZSjCdSslOr8db
syHEiUG6Y6Sbs+MJAv7m6UUUghvByxIF/Zyb/Rl6ATaxp348jFiEzh6ZRXWTI5BE
z0D1jmFWp2HkJ5WLtE9KsoPXExI7IP40GZDLg9A6Xq0pv25WzPCtxogLCqF8INJ9
xc0VaWoc7s9bIZdKF1yDotLo1HHanWyqlWBqBtsWFep1g4wk0B1BugHuhFfafuZI
E9R/KTENacRN0Qc9vnm1oKjgXTCKt7BhNYo3QNg3c0V1FJ7FlQfE05BIt63FaIgf
Y6fhOcWy6K0BN+r6X0uSEZpMlbiIACqaPLf6LP/d+qJk0E6Qb6AfcwQVmuPn3vlj
u53E/I6a1kVcsf06ul859lxY8sVGSpTlulAZDfweqDvQYmzDu32qXDExxzM2bq2M
7F/ESB4NC/5s1m8+bIhVGRRTOxuPnNuBkvCrhmtggA2vub1igFoncf1FF4lrIwMl
/gNGOwup50G2f06vmnK07zrvE0nGkzolMtZ1axi0wjcWSpL4gKr3wOMDNOoXV6/s
+T/zdFn8gM4ABIwVrH9xLmQ+DljGVtGdoqXxQYz3ItSHPpZLNCjSxeNs/0d0DaFt
6Vq/MspRsbySGNhCjJYHiERwtZRbszw1X9lpy5qbZ5j4HFlJZCEw9i8KWlOeHQ3Z
qkH4Fs5pEOXj5rW2J2uMo7u0yxwNRK5kBA9w6UGWRSyEfWLQX7YG14Cdb1uiqZYs
4Ikq6N9St4vCM1q7ngHQbQ4MMNVdTNw4hzFnoxn4A0Qv3p0NF0rKTDqJrydmnz+/
rO/FGD1hUGJnaPTevN+QWnx41x6MLY6EwtUSoInsz12VlnkAmReWdNMrT63n1tW1
LWXL+Dxo29oRRTyubo9CW//kGYlqBQBKvSVs+MR1L0rGOb2pQaBsIzQ2X/GBhc+Q
c8YsZpX1QuiYPAjrMabZISxOp/RjvsA3pDCMAwQuBh4C0J83gzben6JKEQLpCbzt
KFdqQTPUAeFXoqbCKAWgxHTx7odPp5bJATWUfbC2GUAzAB0nTnfxEsMhya7V6xuo
7V2JAomHz64fG0qIEsFxbXctk4uduyUMaywibg4qe6LerIrX3QYo785mwq0K2qYD
BvDZ3LjbRwoMLox7UX3mxNv9DrbfkHBPEvt0pinfqmW1led37CRDNQnlnuGvTylZ
sZ4LIsrYWvyiW0J4OURcpIkIWy727CY1nG6ScXnEtFJhkSOESTlXQXZQcvLIRK5E
jHMiVDahco7RMVbr63IvU//ue2VA7rtKR8euswLH0OJ1pKbSMz6iOfDriMmx0jRR
HCt8REYDmbfdV/mpUHqWAANwkxaHxR5E60J61A/EPreD64zbTt+K57oLTYNzzd47
Qf0IBQgLRdvU/hFLht4OVdcZ0im09gebXaeg0yqpsV09DE0mbZCV3udhIYHB8jMj
Dh8jauAqWBDXad0XeJ1AYAhu3Ay4Ac4Rkjzv5IXkxQ+OaF2rv8IOr+l9LyXLvP0v
Kss+/8wDztpqX2hFuu/3FMGlNOkBJ4tCe9NX42RP/69pv+rSE+1D2JItaP0jOTvK
mx4q+dbUnCoWNqXm5YR4QnO4U1QiG0/jGWihcVdepWAHErqGqEPBx12QvtW4ZCG8
b3YwSFNj/TbLvOTn/rlaz7xJEyyIVUQxd5NRpTRmBY3E7xlE4fLbaylaG1kP5rkE
Ligp4ZozSa/l+GpLcqOHCqyT/KPz2v0Ab2HcuMqqXJ5Z23dg6477djN/3hN0MwBo
PY703t4W/BDo1gn086+hvY55w6DydasykEzEcrIyspSXdefBHFzldDPGnGC5pgM+
KL86BK8bvI3uTmgvob40tAwgFD8mXYCANR0jniX820lbRIJyrVcGfAQddJuIX8PY
a+B+BvU3FkugELqOdTUG1GhZ512q2POHWVlLmPtPyUM794mc8qjold9Bm5ch9OTB
4zyF6kbmVk7BjC23hW8lrt1PHyYO2HgqZnPWwwpmZsYPLCdRgZQHShzuiEve/q69
y21bj/wut3WqY4w4K6jadIASJXnE01P1XfiFPAUI8f6MC6JMM2gQAO2cxT9HAIRq
oxekjy1CWFJmTAush1Sy1+Aq1+3PDgKcQTjCjU0TmQilZPcPld/ilqGEVl6mNf2A
5FLr1GUfqv4wolo4O6sKjq5KRzWETeKPKLKY9pcqsZpNFdRSxhm7E2q8CN9NgBGJ
/WDdrhm7d/83ZyViX3LUt4vt4sBOf8Q5kOXLXIvWdABpWJfBV7MeS0y7ZOdEb4MM
PyGdCP1R+Pxti8b4Bfa7i/m1lvNbfwFrGGWHI4qCPBVh5EbrQAUbBpzWszMcstUw
ypQg3hGsWYj8BHv2Zg0Yn/aI+32lmdlZTp8w7CF6G42ox95Dwc+IxGhi2s3yGl83
Fe9XWTv7DbKxMmXiIF5OjM8VA2f+1e4uyFEoGOCVCtf1SsCkzKhTpLyNJvFtTxVg
rUR4DqhgocvYhQ2n7mClK4fgaDFvBpfmf9i+Xpq/STjTdXKTcAzi/HcztCf1aaT2
ouzX0WENPnVLJcuQR5i2tQDlsL2W6MhiYruIFuWwZOv8p/vXfGKUUwsv05C38Qt1
8Wb+fUNU/75SInha8b2OjOMjOeejuWnWXe0+iQiHSvPZeJA1HAIEHGPTtshLPcG7
spEQEFiPpiW5r9rR4ekXECyOGXIfD2KuJ3sgH9KUmWa71v86/HesYxheJdf49PQ6
H+HuXr+usOFOJFJbkoqbO39HSTOAh6gmurpERRSDBPmxRs0QT7jHgdaBHT1Y/PDC
9aKW2Z/mjvsiOHpYO2Ayol2Me4LaC9qKChX9PISJUqbXMjyOLNG0jaEoTN2fvxoS
MFkuz9KVNOIHvXkQQ2Ji/91mLRWq7SH72MwRYc7yIRlumlJmyo25e5S/ilD6mJZM
hKY+87bsx4jgvU+kLVOp4I7TPU56dtLHVBX4Y9L/B3E6VGB4QlEHHbGsaHfbqZ0R
Lp10sT3cvI1OdQRClgFkOHejyyPeS6jSH1G0ZEyKWExHI6eKrDLPKZwfBIkHRUmt
UKU/sF2Yqkq32v0UdSUN+fZTmbbA4QeeXb9HGu+5qvVB5dnx4ycJCiDfbOrzvrdc
xzMZ+rSPuptsFx7z4oAB1kYFApA6jNxHo+/uAarc66566ujomRgFqBmJE/QlJvO3
Kor7S0vdeErps4NdxdGd6hvflGrr43HMVwPzoRu3nMcLuhILo/ZysLI92JuQyXcI
yvNk4Qqu9VSApY5JVmDYLolEbPTjky9pj+G5yuPnG6tOoIcFnS8v9iFpHoq7mmP5
U8kaVlQipQ/9DHTuen+jmQYAIiXuXVfisJQZkk7WnQQZTnYI58p3pmwvxr3ID77t
E2tPEjb78B4dHUpqFcaTsXG909gNvEq0obp/Rwi09KLGYMbOj1i9dej4/uUe3i1e
lUBkfxvYHCH2argYV9ZI6Lo0MQaYiEsQtJuvYOUIgK5SpURxbcI9/xmpcuQNnypV
TpHhAan6PctcPjYvoghn0p5LSjAZ/K/TzZp/M+M/BZRfNSxz6DfzW40HYlUbuXP7
xpBfIdxtknVTojx8/PvAEY2b6Nf5pfOCWF/gIZ/CFiUUY04edvn4Lfjo/Qfa/4bM
xr3A5vQJh8dQVL3X8YsjHE05UOOE37sK4eqUI5USaOx+OW7VkKcLYmtfdKfxsgIm
7siM/rbTSibZUYdistHtMdJ7WinMGG/lJ4AeIdaZEy8E8PhZkSigscovhFBx/DwB
DFND2ofXmEUMmjNuGyeIc0uXwq3pmQv/MWFddhYel6uw6ilU2K8+7POSsOCCzo6/
YP9ShhgkN3W+Xf6WTucXrpg+TbDwlkPOfPaPjO1/XAM7GSYyEcsJDQQzWag998VF
8ejANF2vApnZJ39b+v5xVOIrj6LATQOuuwG5z2tSYIJTRvX9Mz0y/6+sjOlQ7mmQ
DoETq6P0zbSli6Z+mG3kwEeoGeCgfDaUzdGoQRDzzGjE7NQe2nFgDNlcFVg+9mUl
PniYyMaGwfmFnbcePAV6Y8qQDMD9YI5KwN9tdga/o4VPHKVMTQ2ggSAD0M0KnZ4g
CF2YNnjQaCtyawZ06th0MEdQa1rZ1sXbOKpLn1k3AJPi3gnhnAt5mOKz8PcgN4S8
BAevEZugXMIs33+4C33vi8AI5DawFW2SQEkCO9UFTq7Kkfbxa1xX7VWCAFQx1EkO
y7wXW3IxKrDGyWCkM/6vv1pLdTcB6pGA4EL0L/5BZHr1Fu09/qDCP1yXkAuhh/g+
Nph/Yx6JlZ/mlj28QYyNXVovoM7Tzmtlk71VT0lw9+lFzBPuQ8hllV1dENohJERD
AV7Bs7UVE6YU8GwBhCI4/8+1Zzi8j1d4bqrPoynwG+vlD1MEghcUZ1NJI5+0kbTv
+hC2IzUrT9DvnaAzMG0vFqbrc8NeqXwq5a7cOsomXV8hDo3yunYFMmN8rO15ByY3
pPLchTxjf/9rWuhimOKQGMhtX/aRXbBlWU6dov3g0HOMW0J26U681zn9vx+z3we3
8XKQu+P9iaa3X3g7pyJ5TIsL19AbpArqU2PKeayKhgoVZcNcyrE/jSNjZNIffhPv
u3WhtA0vMAIKGy9/3fIvH1Jpe/7koh3ZoWYLbr5rm/6hj9VFOw9c87hyHJSQUyFZ
68T/z4lArOwF1KMObEUMr+jzfIfz6il+TxhImB9bktXMB9jJOWWj2/Qmyh5MDgsq
YVChbShZY2YX2gMIBtznPmxNnyNuRKPK4GKVxWQpABPD2O8xpLiPyPCrYaAkP4xu
7MLLe79uEPh8yFmvp4FOkR+Sd1flclG3PYJWVVh69jsOzBqqWFvjdd/03/90YRfS
bi14GAM+nVJck8Fv0PHEmgk/zurjzjJFrzJekRRKH/vN7sky5O3UQEf+nri04+9J
he90nbbRXxouJWryMtCXKqCb6shR8YZaAAcFCYoHw2IHcJL10tSeuZMLsGM4pyR6
8Xy4S3qPxxVdx1UcYJIdGTmd1fRBDwxap5juu+52fWs3EMecSBthOqTVYnrYm/kc
Th9GAC/n3n+HXDC3AZ+2G1nuwk8aOBD2glBJP0u8Rh+WMSEWEidhT8QQw5Fn1JqW
/5juqXEJJU+CZzl2senCQnK2ziEMBHu9pOdTzCGKn184ijgoFKHZiMNCXfTcXldW
IAFaC1SBx4wrOZ2Vy/MuCgHF6v/ya4ykzEJCuCigJJGpkahiYgIP3EwolU4prT+1
PHO6BVl8blGk5vgKc7GlwLDsCbUoeA7zleq0UI5FmgSQImUrj/PFRbGL7PBlOquZ
3xJFYq5Ho1CcrICaikTcBpWc2itewN7O2Z5WXh0/iXACbHlA50D+h1EMUWi5tuZm
gIECc9L5OtGfyJX4WKk/HjjQwgqKqBs5D1JTIsj2razLFiKYPg/IadeoOl/Op6qS
eY4kJwsi7AiEEKeCv/NrmxF5vHGZn75vs/kF/qLJpA+E+uu6h6U0l8WzcI3zDzL/
OjNluGgtMA0Zbd3Zfd0srAidwVb5O/R/1dpdvZWiLNL4WWoi6XcZ/kqESv/BMX1P
8nW7BberScHSVXos+mCfz0fFK3RDFC3xTnevnj56TjeaA+XFq9NbYotkGvn4nm62
M1Dg3csVikdCKGvai5pDVE/NPn5joP/jOKhS12ca91bKBpTq0ohWyGHWBVMxDYzJ
m4J0gGpejdob0NIaQgeUbBH+nuzufUso5frA8pKxpSsqKDYj+XxYBAjDV7y10IRg
3z6eTzuPUtWst28xFZxnGGNCutxrXSUSagnVeLaOlkzTffo9dBtoVVotxa+yiWmn
xT+irppy2GnFWKYirK5wmfmbzzHmSoDmRbjisnhapljJbWQq+iYjiVIs6PnF5b8L
LcIWD7pDkHMVcmmD3HfgnGkVjEgZM7PvDkx9u3s5xjC6s9UmghNqGvc0L+pDK0gT
nfeObC2OdLFKKjQJxo7C5Wmr4tIBhqbCHf9BYxe6gVJdManAzLy9DoQmY5MWF9/N
QTx5OJ0wCv9ZUXCag6A6Q2NJrpNTVyKFfH9i/aHWFMFcQm5pB1StnXEWeI/kWN9d
k/a8+sBEiqKPgj32QZRcMiYh+yzK74eVpGBShm8FnuNoQ1YN/HJrjpqh++vq5TrN
QLyTq5OqDZI+92CgcpzGJgDrUI382jpKQ0P7xS5eQgZWTA8m7RgwMOsnEAqMvCOe
JZAPXFstges0gB5HDtRQ5HuhZmrZW5s04BXc/psFnF/3ufPxgVN7Hfl+GaxBe9Ch
yBayileT4Jau39dDwj+YmCvY+f6oTw7VXl/LzMa/ldYZT4yOsh/FQchp1+d+lgQX
7FSyqJy1smQ8djeAWUPJqYdZEdkJyTWKtbn4tbzHhrjQePhg/xHp+8sjWOCuusAd
VtlIl45W6KkXb87gfBuwnR6wG/kEi9FtCkcvGHiGdiegxD+CZ3bbQlDmB2gK2OFa
ahU2ctN9ImMTb2vdgWApWnKV1wZgjZGffWd1m+BdPLBbZlpcMNGC6JEAzbbJFx5q
eGqY4z+ePBZTduIAoGB0GEwg9yomV7Jqz2Uysw1yuSS48HYVMJYWJwbocNRQoo8q
8B24ovliY1tGzt5JeZuwMmaEkkSiOv7wTv3RHDdtm6/Rqg9nQpqIgDWXudyGfd9N
KvRgjodSN3liu9FuGLl2Mkd2TpIBdj4iUJntV3LSEXxDRPy+M9xvieC6bdUuxLRD
btgTCSS7sdtayWRyeLRrO3uBKr44ydFnXfDaHSJ2CpKi44+m4BgaXRpBBkuvXpho
ClxINjIqX6H5yHpVY5Bn7XxTzDSq+o1bGlO98WiI0dbSjiwSHP9PCaRvXiHYDsEx
p6UhUxNOTrN8G0JNtLG+Eg2OZ9VKVg15cQdromI7lA0ZUsFK6LSIycSyqbdNSFYJ
opOna3B2pK4mK5SF3JgEVCjsgwfEqMvffpEGJEu2+uBJLtsSet4R8iBjsq1zcnaQ
KfOw5HyXYg7zvzlysrl6IpK3A5Wmfk/tXk4t5mkv4BrJPKzq0gzStncdutI4boAt
ZUeQGAxWtlyobT4TPxc5yQG6wlQidaqWnUiYGy+fmxzgTqRFzrv8KELJccV0vpzf
BAure1aopncvg8PDGLNC1roUkC7IhDzWFc8OUkFM9LoMOS25geW/6BSDiDHYxo8L
/6UaZQBd6XNXJAdxfZjbyS05PMRLJT/V3Y//V3AHiwPJasS6lazuspalhe7TFENO
vse6lsOJ20RMYaN01zWatSQJBE008Jpu+5xlQihMHGZl7QDjTFvcVDXFkyUvqSqV
FefDryh4VT8w52MeMmLpQELjKiSL6vqnfmsoGa5JMsq9/ZPY/BueZLJJtkdHOPmj
L4BGpgJkWs4ywCOHBj3lPda35BGTnOcwvMFnp8E9tt8PQrppoKmmdiqlMYiAJ4U1
Agyl5uZlsP3O3g+1fnOVixIRm6Nb0UuZi6gSxYd5Q2aJ5s9Ve49voFYjMr4tt8Vw
mK+hD7ZOkL4bJvUXWMtTPkfIkS30MRYAaz/26k+aGKqXyy43iBUJuzDNmFnayYST
Zo0rlb7FFuEXVL3ss/NPmUfzDzshlEl0Ew06nWPCQb5EFNorB+8iy2d9KF/iHMoQ
mzW9G4nyP59DA2lxFHVGYLl0WjMmd6sd8MBvdnMQKsKauKywmTKW00VrqPwsf39Q
/ms2rf8UOOI4xfqRoLLPbjmv4fie2o7gjATKIQ/Gk9hG6tapIhiGKHfs495UCt61
p2CUn0rU0RNyqjBMU3aZSsDHpP1KSycRhkQNOdVZguYzHpSXa+mZIoD9xg2XSwoq
uI3CWvHx2d2W7o+iF0zRJlETk3MrrbrggtmgEnOgzdS2HSIDcgvSG+gyhvOUxxdZ
WrWKDN8/eHIIEYj/2peINTN/EGK0NGHf6Ff/3CeWEk69vh/y/o0Qeghgtu7yRU34
+LTGmNMFp3WAqHSSXoKis+HERis9DNVYlzuhQHlMRfuYw2wbJv7jFQQi6St7CUE5
6pLE3Br6EhWsNcqlclOsi2wSXq9fjreiXlcnxXpSo+DVyuk9fmiZv9DDh5bfemLq
dOaB9c8ooNbKMMhmLJVFnxQcV9ZTg6hNdfy0Kvp/9kwRtsr2z8JZI7FXfVGdqyOL
8xhlEvLkZZL3NSAwA0SOGK4De0J2mB7WaMPRPBLH1l5agtwONV9/x6Ke4A4c30Xn
eWSXJBsTfXVhK1yylY98iij4g5fJmH7/mxhDvqWHJeWzxDEfuejFYFhtmsSz0SM4
dGVOvMtQn/MBBEghEIgfhMBvlspPv1++IrjKnkhQXXnvPmqyZEzmk9+dDS+F1717
MTeEd3kCSXEHt0OT2ooOmap29f6Y5TAjKkUlKuAQzE6ojtVXwsFPLf60cN47m1fM
F3xZlNnP/Z1ytlyxHTMO0k7pX4sMhTjPmEYGcl0yr2RwcEkb+oBP2wRTNXnyPDGT
ZpAIVAb9QLk2sdA1b+GmyD6vQIFJ+Vur/X+tupXdCzWfDuX0m+Q8Ang5Efypy/Aq
ENBGA48XRq9ij+g6bI01gqSGuXZHku8TV+p6NKrZMrthY7VoSRd4ZSwLxpNOFyw/
rqnweZ038Z4mrU2KijFsThl/2o2EQBLJypj4YVTy3QNRv8Bnv+aBVV3aIe68/Vi8
fnJYe8tkr3kyjDtiexDlkN2kYI29I/aN1EkRBqYCxuhKrRuHXP7LpgHMQo1PwpAM
74CtmOfZBZgbKWbO7g6j+K7+wOc1pYWOP147JjKU1nZNKwuMsvDb690glMwfWC93
GFtKkgL6qurL50lipGzujxAbxce533Gm2Wtjg29h7wYmdbrCpkkz7qzRzE421oGB
LebLbFpoKDYx3AtyY1VPY8zaC6YqcvZjShuLIBzvdZELdHjajk6QPMBqpUkSX001
WtIDADWLFJQI43qZ2iUO+t7iQDJcCLEabB9TkKYJC1R7sZyeIyMx3wfzZDvjyPkj
HEz9QK2DJXBLHNGzAx8EqWBdvu/riG+sAu/F9K6DIriNw+qGOcsVLne6mWX2ELMw
OtFKV0T4UjMYi1KpyiZZLs9GKKH8BFnJbNyZHjKw1yAqpSDIJhu6l4j7W+UD7mDl
+/IXbj4yk3dQz9O5C/4ZNjO+Kou0FGGzb2pOUcsS+ac0uZjnwH9jaNUEu2V5lN1y
WJLCM+oJH+/S694F3DD26sJvkSyAdrlwtsP4CHErxcw/PYdkkQpuQsP1coGBOsap
n9s18WFgkJLmiV/ArJ2cJmLqx+UCblCRrwKyFo01gyO7ZIzqLpgK89BfkEfVmTvs
/AP9mCaPhWPiV8/hvwY6nqeu0Y8X7Uw0MC9DlI2eqYJoKINMAPGGXG1UWz0U6XJh
Jayg/lUIiqYx2JDNASAR85W74FAQg10Jsiw9ZE0Ck6OFwmKuoySBCnjcRh5HxA6K
9kISmaAhleF8hShOvPCkwGVsq+66DGzNfeaRXEQThCLLPRa58Weax1quNdEppOrU
n7pQ2X+Vbga280qZHk2zDz2LDD+CuJdNCCGP4QU9V9XvXvzRSrVuUBlobE3O5+jS
gpOZGtjvpjVK9hn5XtOpddRFo0ckl+Qvx780o7r8bmCNRRkWudwpCLrl0gtyafBO
va7EaZECNYojMDJMsb1lxPylNwoX1Lk8K1a5jURoeL9EAqz4QWwTB5SmGJHfb2BJ
rFiTqZcTR15/InJAaHwnpt1OGapYTp2lPpUke0Gpb/CaIicfeJDM5W9VQZLymXdL
xSEYFmE18N4UB9ft5jyZVkg1MWd5b8QbEkqerEi1Su6S3QZSsYO8YFX88zjMwE1V
7Rs/hmXDJTktU0UX6HTdZ4+tbDUWLCO5GzfCtnjVqsN5dxGWLYjN82pzA4ft9Yyz
ggNZ7v+TJfr2TFctcfU+EAVS8nu52q2ElEDQZXbA5DHZC12hwUMqe3a6z7ounk1Z
+ikNX4h5a785K8JtC9GiAcxBkWHTbwmAY4nkj4T9x8m5D6doyzwWO1bVpclnnFCi
1tlLMUWkZ1s5OM4c3WUqzVcxcCSzGfWPjE2pCvgLqphUyDZaVkZJzzAAvX1pt96c
4KprKXZSoPWNPjHZQnzAO5R0hBntBdyjMyGgeP0EgN9PEyKMa2/M4qaJhvJnIg6c
rUq6RdDpK8VU7Gpg4+wUS0hIyj5feOr8cQjLQBCNUNITDo+I/UMuzU3eR4V1QUUP
zXuivcm9knN6t70zZny0YInvBcS9jqtmJX33T7/UAUYzsdOsO2hTJnNgVPluzKT5
V893oXyhBsME7BU+HNXqrH2dpJEDMjiPx3C65qpXX+831u9jg5azLeuK0+4s4IF0
03BOzf2JiMcJlm0XlVlf7d3c0IPNuWzOZt/0zt9LU5vXfpzqwxsJC0VdpS9eUxQ0
qo3rWFowL24QLTIf2SXN8xZO0Dg0fe/A0NBZbay8z7hz6GUhhPyPatKUFWHn8WB4
1mLmG8BWwFLAxrrD2Jufttci1NUu0jVYLGEmBX+BZ6NXpOUlDWBh/mGVbp88K8Jz
8zsZiMuJ7jOijwaU839XEvbnKTPnSEVGhsxL3phGP+e6Cz4zIDQhEf8Q0vtQvOl9
pa+y7r4zsFQO9ODWYRzDE1TcsxJJWMMnZ2SYAAkw9Fdkm1cr6ZOdnoUuvri9WXN0
GiZbWaUSgmDCFHjqwbcC8mMpf3kjUcsIqSxmA1bu/WhkVLRPBLDC5flxITTfI75E
qOpBtwaXXTw3rtloKFkONJuINeqnunlewqmiUV/57/QQnfoWTVcKBWXcFbZ+tEm6
gcgZYG6PxzyK0XRfjUondn0ZURIpFz3zK1HjIz0bDzTVdt8yDI391KS0hpbIS5e8
wfHMND2CQ4xFwZ2P7Msyh7oVDR8ntnVWxveQKKybkIYDRy5J13eP616xaZm+8PJM
EvHgfbYbys91CDLJG8XeAPR6PJGMNw8lhW4X0QmKJroME2x0smaHAQXyOF5JsO+I
Bwe0BIaoHpoK5u1XhkxneqfXcOas3gWHPzo0q9PP797HNj1JXfqElK3otPa4SBYx
qinFu82LuRkxkG0v1cq10hPVFzUguuiwHp7Jxz6Q902bTBIXWZmlF6ZMVuafOoyq
/wWYuHCUNFhMP0dq1DDRUSrloeuddwf0q0uhhAFc7qKzwKSrn5RSuNV8ESEOvdQe
/2Eq81BVA4TWmUcrfAg9hQxJQVd0i/npJU++lmGyHMW2kmapIBHhcqHpSStZ7urg
F+iPjPIkWyBW4nP5V5vbpLYUNMg5OaI2F95Lr+HkQWibnypb93pAE0kCdQ6XUW3R
XkecAahDzNsKEbhJZ1czZYfU/jxbZgXwpJFvWXLZ5YsujE97F23KnvqCqSri9boK
LrtWNNwwsuASTC/Yu/gCbuTaXwqQbGuXyQ+zfynoZhOvbqDvAtLd1HQLRhpzxMnc
3EO1b6+mwOFeeJCkd3KWbjLMMbFrhqz/19H9NgS5EOcHvJWj/zJWQIb8+5xyP145
xTecqNghK6FD2Qa1LFAEtBmiFkk+mf++lSVq7IBVYMMmHSVR7Gzr8VdsoQWAFni+
UsxJcR1cMpCvjjVBdaonv1+5Vnwor0uNuvPtW0pcgLg8IQ9ikTft1n6O8kZbggpg
u5UvKRJA1ciP8UTYJpQLLplWPuBUX9fL/dbnf1S6jWktUqhLJpFpSKoRoYjOybxz
Cc2rC1qgQVImG5v9GYSpRc+R3v6zuE8/HkuhfiAokGnH9dUIe+WFHyPlrx2EcbhN
el1j1Q09lMEAda6a596N0YXMJzLwZsVeOOaI7zMgPn9iSDusqibaXLeX18KOK8oA
WUn7SBcIXS5IZqI1jwgmliB3DUFhxSLr0kZi29sVgC2t8pGtddQr8DKDh8OA8JR+
O3y7fAn/IL2y7qL9l/jV52z/+IOA0AZ2p+/lC4ME4fjum1W1IiVhugyw7UzkdhZf
rKjPbdu/mm/KN+lpLM8LJd38MMn6HjKCm7WLV3hT92hgemrmv3eMbXImynp8WGd4
JLLHGFv3dvjsbCWLCmtF4mGYTBET4YGBsgRV0IaHyte52mfXxHIz8h+5Qa6l4Pnm
nmhBPlGGGhKRzZNTx2rfNr9eu/Xg7qhZ4SyJ4q42Q1TPvPOMBFN1Dx0oxYbPrcrJ
eP0b4OWauncoLLfEm6qNJlh6iHuT9qsFSCRcJNDIp/eA8NNer+lvXX5JwLB7Bbmx
vUkNPbu3/76Q1TujKmoq5QqMRTRxAn2FXFpXLnoRA5x3J6rWXiHt85R/Sc2PBtwt
xRDxGr745pf6QQ0WYwlJ3HfOZOwbkoZLefvvFTsCPyTs+AuMv198CCppoNEA33SJ
xzFdoDJ8P0Q3zvNmO6Xl4htETWd0qwQ32u7qtX/cjqJs3GXGEWAANtnamDDRly9V
83PEHgpwV/wd0bf4Lxn8W821zAsUyxNOzJT7RzVz8skL/xc4zjbEqpokYgBaKbyk
84WaSIWqzTloVXYxmXNLR07LmI8KSbZXSxPnG1/HEnGr49lJmGOyxmVK1Vw0Bgly
EVAut6jQHSQjn6MMNDgrA8O60vlypmgAMIkuqCu0AKpaB3YDfYSxGlA2NrvElVw9
99f8ETsxbT2TedzrSTqn0ftXZrL3ZgpgsB57TMb4vfKgCbS2oky8I3bcIAPJx4bU
EOWT/wEcWb8y0qMDBlE7z6O636QEgr2E+VQAH+yxEpPdxtoeOSxxVNdUBWRWwZDG
/gNcTkFo/cajVWVBK8I1oMlY/JXk3L5jW2MFQM3p71XyEhyS3NTwc642XjOMKqG6
2EXj/VBw18gHhBm8XQoAYoG8hKUQ9Usgr56wolvirAn1bZug9pGyA4DtjbopDEYZ
L+PKSM1MBqZrkFLM9bZhJlVLZrmjEf29rvtZSdIJu9v2p0SijDfhyUEkJiko9JF1
+e51TFzuXIK6kBDie1XWpijwZZPdIRR+F/4J2XP4wBs9rsbbVjNhdaQFRoXI9VrR
KpuH09Fo+xZCBlJPm+3Byu+y/oGEnDIOq7+saVNR2Ky5Y28+kjZ4TXQiHKNLoPw0
Zt9UWbBorI4Fd6GRsmH7mjii25BpLNEvfJ4oCM/ePBrzJ3k5g9RqOTt4oVF1msJ8
S3aUz+n2vbAV6buEiK68/sTAcYPg67WGURy1GPp35cYud8XOo4AHthnqT0KKPbT5
LFLPvkDbAc83Bxvq6h057nQCbiad2/Y94lnkJEMlB+s58eSE68/Y5aeJsJsAHSMP
+ElXfVnOeoyTva2JGiirQNbrnCqzuyZAbAmIndCIY3WqRIeOWbg8MldLha2Z0fn+
3S15MY8o8uq6QK0avxcbQ+GBLG9CkxNy26UYC/JSWenrJG7NEgV3fNyIuVrzUibs
Wilm6Cq8Sp+ymmIYJa8jRtZQKUXR+oFW7Z5vXEEO2wO6jDgFLNqGqVtVs2I2/Xhp
o9iqY7L5tsKGIS4sVWWR9ssVQwgNPDGikRbvH12H+zWROcHI3n64d/tipytXgNvq
J4BmYsaBeEs+y7BSomBi9xC4HNGzrD7sVIYIscIeKNIc60j9od3ve5ipVewMMTg8
k1Ni0jiiTgJSjK5aacNmGtLx44NgsNME9bl5X3jO65lVOEBrm4VAlhkAK82eddbK
KlXxhT5eXy0TItG3kxPviR+XDemDS0Zgmwj/LMRtrFOhcAhrhJrJesMUENzHG8WL
HdIjPEEHd+TSP3taJdrPZB5IzupwPiOZcOjnS4MeEcjWxDWTETtbdJHo0xnj7Ny6
bwMPrqjmFoXSW+LlbWp1s9KTQoZ4FclTPr04jDm2q/fe2uaVBwbhkVjHDGFURndC
sK1e5JoNid4Lenr+uVeyx/70X3BOQPMS/2U2HdeV+nVAKxeuvJufIbi3aDK4WbUo
yLXRlmZN90/QBlz106qyb82Uv1Ak+FmGC/PX26IpJE5tHJ9s/m2qgHxGZBnSyLtl
xVICUVt1jChiFAYq2Yahyvja2JY//DpHTuewVLZotrOkpYujUQEHiYp2OBZ47vz3
i+aRjlcnzZfg9SV2JWjYm0K/qpLTgeKvNqWvUVgvlIqURYhGqgWltvrucoMuJ//7
sbkpJefYZa4XN0WDAhDkUJ79f320xqVpy/1IC06niWS6m8j22XAOd3vjv9VsW/00
5xXGcuuR0vjVF0dwxb7K5TXcSErvYS8EAFZ58Vy/Bv370bZvk2BffeXOQa/qXgOm
FWfEaEy5UD2ORidb7yNeAdzfoXfy/TsDGGC15APT5h9wMsW6cpZodSBSPjiWC2uU
6SPlq/WqaGEOLbCZuYt/ZqBPSWez6xzGZM3Jj5YTLZcO9jXbvPl8y3zpOKpBSSbA
yr3yNztVAvXJ0dZszmgJNzz5nei7RDew3zVTGqr3NG1JvzBGyXOtTBVEGcx5wHFU
g7DniUJyT4f4xuP5adGGGktzDPzYh3SWFWCu/MR/3isiG7B5SHcORLoar2gjdh6x
97tTIR//GDtQ3KkgWHUOMXspYEh6amkBGj13l5JF9SAVnHdOyrWMs3loz4i4cuEz
kShq/fai44rUczfG40FQSAwMv1Bu+ggJsGC6zwzJMa4YZBOzUqNUOqbepdUx4m6Q
SG6icusLsr5qFmj1W0lnB+HhZMpNSlv4alGicGVe0oAYmmYm6gjzVUiv6NukfJAQ
6/6vW0Y1vskqFW1IOjyJpjwbGrblJEUJGAQt4btGygas4UrEM/OMQFsP9Vb+szF/
MZSeZc0igod4v/H9kNz3A+0WKxkeiGQEIjs07DE9KkyeJo+pbacTrp2vjkKn4m26
qZNvXGdmE3+GKxLn/dNJH5fWSTLgCpVAVdYxUxasNBztkSWBgeD6ouvCl9zVUDeE
x4eEzHi1sglJ8JORLsDWIpMc/XC5eGjtH6/ItN/0tyHdEu2vAXT0cG3ZtCSbJIVy
09DMC0RPJCfDGv6dJKpDaZ8Fs1lVXtaECh2JlmVwXxe8kMwAEHFLbSq8yD6vNNCW
a6PIbpxYt4U6TE1OTQu++fSg/LtoJlHh6iot6lpQmT5QPkvxIs7mwEFPje7C/jhH
y3VXTamsi2Hd+M+cPVJcySyJ4oRoNU359iXOYWJHtYOl86W2mOa8ePNA3NTdqp/W
Jrxhh7H3ZJ9lYIXDLiRzS+1kraIdwIkwZ/FKEbZXWzOchhpul1eOQltBw4R51dBr
YEcavu95zKu3YPlaZBn4U67Nyx5/R4h5v2J9j6qRROtzSeptrX2CvQ38idpWdaq8
kPwQQm2eWm5R8G3f7jySZ6DEvdTxnJBbpFcKvEAGhglMsXFSknE8xFdOjRbK6Qgz
P5YblSEfTBVpxLDHFTzmkGKQf3q7gEqAtJNrj2rpoMCb2l61idy/8xR2i4lN9vef
AuIhTPVQAEJHLn2ZLsNP1pJwq9qgvW72SXTgzbvz+Y60rHIr6kJQqwkY2eP9tUNh
MyHUdx2uO5/fUGHj0VZXkdpwbwvv/9/DHcJyJ50myHGWPVgW6NdFzOdJbROSQLy8
IEy1NcwmfHBUU5Fw0Pjp1zRpTgJNAeNJyjmwLYMP8Evj/UySp5X7/itnkDYFoLnN
Kcewvkd/2BzAZhbULrnW9/yFi1uvsDZcO80o/GNDj4I2Ye/bp6wKvYroaZ1FWjLw
GeKVsGgIfr5xKKy0CvFNvf8eflnTHGJHuA0vYZYGX8MV4tqezWikFXLQGty67n4J
eysj/5IBoyneMa6zdlRuACtHT4YjuSoi5BuNSgaVmZGLiYYcdM34PtF9KkCAvxHQ
u7kIRS2xwLMHmjY9mxPMT19rNvZaqO8cuU9tn7r9QNIyY68CEQUEL/6GZmNh3jjQ
9Q2v2F0TkkOU0VzGhiselWkLw7FWbcf6iwaDJmX8DDcMiRNJ9ix2evVyyvqCNSA7
n6eJTORZ8B7Vyo0l+tFi9fewZ4Wn84ktT2M1SQEOdXmeNZ75t/NYiFUlQNXyKQ0C
AiRWGbot3n1Xb2yljc402blggQkIcFv8V2ygehcK5kpD3hTC40VZeGjgXmBcBAff
ROPM+sSae0vC2yK14gXTpd9OtTJM/FTIxz38eP+Xnacma8UyTFFvy6IN+on1QE9+
VoTRKc3BOYWR2SD4FHRP1hpL1O3t4BJsmIvKIxvreLDUX4Wj96JcQO7cpFTbrjPr
gNlsROM/6JsoxOd7zD47T7Vg+sF+ompVlJhtr2l2iOFQ0CFpYJgAx9tRwBgBYoNl
s1TM630K+9UQ3ILU3V9PHpIxtij1IxT2SOQis1MDr4Zve6SHfn7ZqK0da5NWr72Y
0yY33JLdTparh61fj8hH+02lv64VXUArJB08lvlg+iO3ULCZBoDlH3I+vTp+yo5o
Oei/E9JI/7JzWALijDnjiW2KyZ3yIrUatkrvvXHtjV5yNQWqIeNBNsuvst7B4tcF
7UYrNkF7ctxlW8tKXE7U/C+Cp+HwXGwxccZ3R1k1narw2gdGH4QWNT+YO4baEtb7
k22Exon20+E1+pZ64NoK5xfRqsg2ZBmjcsWQJTdwQg4CMavCc/PP9vlnWdYsP0Wo
0xAzKcTgnwZ8pknG13tG1XAe5euxMFCS+oQhiV6BV/wjsk7m0nLiRmUZ6bxiUTlJ
bNBNT5pynghA0AnqY13o10bOv/wLUu4uESjGYvNuW0dJOPz7gFvH7HOTYYEVnwTC
ZPjAbrvHteO5s/kk3VB8NZKo50hbxZgl6UOjoFTfdnSh6bYhcfFHNtVLXAqnZbGb
E3FLZxV+h0QoasZyZOQSIfkVxw3Dpf8k78Bmr0R8C2jsHHmY9Gca2Mtz84ZcP+2a
h8tN7HDYsBr4ArD8eAiaB/rnbCn2z/Qg1AQNFKXfjj+oJAYTJLd58+NE8rtPXsl9
G9ydiHtXN3xNsNVckGoSit0e0M0zmK8z+LcDxqt5RavS5rzlqZyKhndb8QCKMLdP
iTGMcpBPldphhMf2lMnDOf5elkioAZI+VHx3pSsBg/tGRMIfYRXfJHWsBve/ZZk4
NFXL6xbcuV5ZsSobp18QxNVRhF0t1R+TXh+4uui0vpFpDlwJ3qStcW3SspQAAu5T
pXfqaP+HcpHCQQP+JIU/ttMeLdYSVx9PZcXVM7yCtvz2FFzVen9X3g++RGNziPYq
0TZR02zVtCj5Cbk/FGFfcFY77Kx787pTmnLshajcrEywhh0Y08eMunbMhf40/jFt
08ydYWjvhSNrk6P4Io7ps582GRORAW5PFr1mJJwfSOrPUx0j/SvpAT+rTvSXiefg
d+GX3vWOOhHV+YNsIJyLlqER4X6+78Ir2rSPUW5G5YEclu8keNfz7NPkbvSQwEgC
+q/tvEFZSVGT3E32533319WpWAWWDjH/79NxTvR2Ph7VPu1h+MNaky2mIW9sxoV6
8NnQwMea6aRG4RAWDLLd/g5B+NPfAhKNrhJBhr/j8lTnTPz1xrN427Cq4XsYLYLy
Ehuc7cYkCid4W1KW1EVJNoBO3X3vzl0ll/vG6075gJfCL7CdZoaYi7KwGa9CDAOj
H8aq1KwKFoezcssG3YOtfiXEo57jiODN4/Nbk+uxhos5qwgIawxKyx7sL9Zz8Z/D
1s4ry1m4ypXlH+8XqiEhBGUn/v3a8VhcS+7WkjWgp0AebGAAi3cDPVq2zPK11fMy
figxOj2AKGi+chHRxUAdq6cyAu0vdRg/78qp58sVk06XkA/U3ye/1MshLJJiT8Uw
l8Ev0/M5tbN8iU8Mj27PfW9gsGR32mYYDP2M5XO7Xf1CB61tlz3vms3MSh7w6G86
qZfIiorc0pWcUblD2EGBS/t0txTwepjCYPcRo4aPH4AVF8OD/lyvW947oexZruUK
cdoazJDNevg9WORANOzbNbx4GnB8YAoXcvnfmWf/VClh04R1pRcbMPNKETaZsqzK
VNlqb1L5n4A3OTPQpgC1/GltQEI4hen1fiVasUp+tqsZufyJZ5f9bHVO2w5YhAcg
VpN+RAaU+7PdwQD3nhpdMRzyCW8/VB4HI1R79AtpRq4srTczMxZ4VH+fVQQv6GSB
QX3CV4KWkOtvPd0TQC9Od9Cua9mA1V8SsE4YFexoiMx7cKxVSi02iMveZHIYLCjl
hfSmii5pZ110LIux+ZgRQUdVKvca4Kx6yjTfj4Hw3QOqM1ikhPgOskuXC9AVORGR
wQARrVUkizLAZCuxER2wX4fSl45ioDoH5vnsuCDO1/RNKSXwpTq+1/0UN3L6Ieib
JI1HsjlGmA+9/rtNI847Ev2NEFhbE9D6wZ9/7JcEfxEm9Br+YHfe/nUPXUpKoIVi
sOnw3WT1uaDph1CqITBbs4W0VCYCRFS2a0686cLMepQO+xX9ZAzBquD9fzS0HJpq
0vtBGmEGbTFDfQccM4fToTR+AlzuJKZU4V9cqbT69fDbBI8qA97BQZzwi7fHgIhG
I+6JgEpzTWuUxxxUZF2lGNKN6AmmucA3dkWQNLK6UAthkhhml+gdxItswZiYNNYZ
XQKcNErZMS/pdVBoPS0OI+xeuD3D0dF3aYwFKMcHDy5zlea4vBaxyCDsXpzslzjo
aGCIbWj+Eb+JfqXtJlYqt66Of2c097ix4hIuX5Qh1PxelBfkU6TTuF2zJtKn+KZu
l7DtkAmEeCeINb9OuBi0w05vOXHSDTiRULgVFr5ukVpjXLwFaCuWfaaeBJtNt2kT
xmcg+jZMmbtPfc5ZMbCGJ5nzmppqhE4buSrAmD/CH54/YPurTp3c3wnNLSdccFei
CZ4tFX3tZyOObKCpFL0eqDeNUpnxZsxDjXYWngvsZraqetOTaa+SUdLTIQhLTH7S
BX8A+kDPuVRr11y2JdKt650g9eTwsC5JS4y2Zv/h7HDOB5xi6vb6DL7Vkfq39HBG
ojFXNMmEA+m+WY1cBevaIL1mva9PIybLTNhdn0xZx3FlG6i2VChRnH6j5HqkR+hw
cymFyHulFlJ4Xg6vU88ftGUiV19pIbmIxIWtKVswkOlA+Gxnkxq6gjOHPOHnyXY5
YnjHwuAaz8a3HrxE3Di2ZvKUFplpwLGqfanSJGKoNjwIxwYkv/DrFx9LkM3hKFDW
FDxkIW9z97GTvNZLxo7DTZNREZwQiwTX2fKCEnUl9ltYWFixS9Hw+5GcpAfA2JhM
mvScwEZwoV/feaYhgGxBXXzGtpT3N4P+LxtuVZIi/nM+6CkK33eTVFlDcPGvwyNM
vhXS3WkNRrSAR9JD7sw66DiTJ7qgaaNwZBe/vzLuVhc80IljDQf4AAtUaFHsZsXy
lBoqg23De14R8gjQPwJkd+w5qonVi+qzWCxBkKro//G3fY8SxZZgQ08oyCTcx0Xi
YRzax9/AuJr4EuUcaHZUOq4tFdoi74CcRnlO+4lJF2dST0SQXqWgDzmqVvrkt+3U
8/NMT4KaMyCr5cucV1Lfj7gxFtGrZb93PYMmpx8O7zzd0AqEyf/7z1iuRnr4SQxz
sNppvbTMRRo9HITFBrpftVQ1w69Ss7W/Q6BiOmvpL/7gW+7xVxplzDa4RM3pLH2X
ihJDawjIWRC9/Btjzh9Qm9B4MBGB9CQlNr09OppIufnKMc473PqBsGC1rWtlJ8fq
BF0Xz9AWyvqaKrEzsSQMg41kdb9FchxXVR8bH5S64xwNiKrthWws0Z93+7fXv5p/
OrgkOm8IrUVWHVdc7SHkVSouU94kHaXJgSlkawEGOUgP9AqNkUNT/GQ7IIs6G9Mt
AWaKPNXQ7RiwtzPCECO1PcphP85Oi5+CCz+NCN1ZcuZyWXZ1GUSKh7KAWEdT0EtM
0QbsYjffH1ePVhoXCvBLIYMfjRMT7QY8LdNIv2HceX2ykLevirAr8fjxx0iZDnsM
4lH3O82W/s8Vm0Iw5FaiGtE39crr5jos4K+2bdnYgqDedVkpdR2po3LCzoIt5O3O
tJO4jvJ2IErJmKQ9ZrgeclQ8mzbYpyjbIbZXHPyiP9wzW7rzcIFzcyT1CezygdpZ
jVTAziM2MfNa1qqXWBIjwtOjbbGM2Kq6ElEhFfbG3V+JkNwriTy84PsV3Tg5sEjG
1RzKNn9XRvrZ6Qx8g1tCpyi4DCZv1j8ioceF9sm7ZfkA27InVxOoblAa+aIlSur2
sOHUxFeHAbceI9FNhKRnamHsJrE3hLSIiyuKy8oEmPPdGxL+r+cyaW+5YJ6Skg/j
ooxj3t1JJbLWqBe0Hzh2+fE+97E2/jg0UDcgjoON0fBTN3d3g0ywkAirJVEboiEU
mPhbP9Bl56aTFbORWSbFkE+oaAmycr+pl5mpGeZKA+4xn5KGJWYw8S/FreVrj7c3
9tKGptf+9Zp/d56c/rgAODU4OQPVBuUQ2Lgrlh9r/igYOwE01YB7iP1uwXNrMgqt
IwQ0wTlbo9N43tzx0kfeVBTWVLTn68nTCY1Ns3yrRyitHe4Qu2g4tMik6ucxXBLe
2uJdVtoQWA05q1/vzEJjMneePNvzkK5Xvg9halyoDc4HS5EJgPpOlOEtcivZ5o/M
Fr+gweSXUo3gv2Cd+LNv6MwyRv5tPTQSGWRLjUoAgHkh09jZd6dIlbrunsnPve1E
wc1F/H/ksWN75+onpfng6nHUcOGc/Cbb1Se3Vn7SNxvjjRh9IYHY6ly27KZgn5mP
MOhBP9rF1spSX+Ownm11xAJBReJYqw59hQNVwRNqtHiVccMqn1Ro/O3yWqGfpXp+
LBnTY16G89yDQ9PHAdesvT0A1Rt7uIJNimOb9txm3cqPRWqgm2TY2dAlvDxc+kxD
UWRpHdRZMb8ydG2SSDlw/f0Zgfsxo8tfn1iLrN7MAPLw0M3n94bjt0R/ea4TYRrY
XLTymfDXMzHBOfwsaUkame6RQ1kmiTwZ27O6hNkf496Zdd0vhMFoY90GCOkwF3P+
QVrzWPtP8YetHNVVCqOfCyHijxsuwrkUXzzb8KZObtqRmmM+8YiE45stbtgQdpFX
MdamRSUwo3RdOND+aZkMTbSmSWYidfJ6wxMCfjTvZaEuypj783ALe28uC/n+VSIv
SF+Hpw9FLlnIUniFudtWmdrJjEILYAIcaFRgLXk2zylSK3g02GtPrSpJyyG2PbCs
oAr7FYQ8ACYGVOwd3txjaqDgGHHXxB4KIrWC7ClOIBueyLRV3qwgvKp2HWMZsHQm
75LEtR59uHMs2tDJbt8QhuXGOepeVZDqmIhLQs6/scgOkwzl/TJG28nkZfSfWocw
4MYwD/ylgaUhloSS4/SM4TKnmsoAOjgU2oSvj/RswOk863npttTa0qoNZYFcq/Z9
EtxnffJlQg5qjwf03FFiVDB5VrNWxMYRscaaPIgm9D8z5rDB4EMkx025W0HwUnEF
4Btv1wf848MTuP6SCu6nU4TlpK8uCTFTGg4rQqSDckhO9+bwgeNDGQ36bDGThSfx
67IMbT4+I4L/AcCLnRmNf3XMB83tw8n1O2z5yMRdlWq/9rN6Dyhk9O+9YHvJMfqV
qdSBlW7Wx8OQTiUAL9P1782dtvviqKkdFAS5NVM7XXjSDk3zgpZOWUig2NcfH0x1
yGFIHJQg67+RHly1DTizUz4o/VsrLrjGpXJlD0cILnD+NWfuM2KsPVzzPodAxwDI
lcKCsA7XPQUkSRMF05yOV58sFLTKWcexKXyV9GtlIebhz5DDjWSiM8+Qz/t0Iqcc
VKny9st6+DPym8RfEQN/TmcwVZMBYIpBLHpM66KhQlF3gB1UKiXAH5UyvhUMD8Uc
8UpM3hDkqWiNISbFIr6Qqz6dTdRc0KnGzGx/hjL4Os+CsNx6vzsFJ3ErQyfw3wAd
AxVv1DNqRK6a+luPpVM/yJeDBmaIG5d0Ewp665KQL7n8DkoW76+5p0pGUuYMKqX7
c75wYZsr8WyPNzekq62dQMOnotMXIub/EwOQ8JHL16RpwqaOnb/UjNOHquwTz0iK
AEuOna+CTKRIWoYykjaBAcK2GGmekqHzsV3BiEgY6KHO1P2fu8GoPijnV2uSXmnY
jHF/ZsDuO4OWyTWJC72X7AY1YDbLuibNtgI2iOKm7inEV300i9YWiMmaI4TAq3JG
6EaUZPKNhvSeqe5JHeMSTdJ8FGwswiupR9zp0pgL2MZsSOVM6uXdaP+WtGZobL+m
dVdzKFugX2MO40sU0o0VyuqN1bK6C+lwtM2JoIZ7rBgZLNEZfGWa3lbaTLbrd7Pm
Jj3Sz/F19P7Y4BluS98MeevRZqQEVE+leitCZcCr2SnskojI8jDIf1Q6Z/bkt1VQ
nJKPbBRB/Q/cqOVkjBfU4+OhTCOKwcnY20HqOXsEK2dNP6zY+jKrKExSS9xEt97/
l/fRgSp0e9jntCQmtjVlmXSf8If2mx3PkHR4gaFkPnnD9GfEYNUWOwOzpj+KQDqJ
bZUvrfdYkZjo/smNkLBvC3rpOXlR1nYtX4HeVGe6pbqF+s5Lm8Id9FFNvU96v6IM
qwEGEUQ+8TI3ayacr3MTznWvY82+LIo7QCY/zlhuZuLB0uj6CsjUjuxthJSacVS+
PeX5JvxpfnkM5Tjcw60qWM/MPQx/17xxE2dmFH+5P14TUCvXpc/hwX8uKkdN92l4
8knxzmYEYzR+TsqL0Oj5MJV8K2NHkOVvbk0PcJ2O3Gaw8yw+wuPTEPzyGlKts6rH
JrbRqNgr6HGahYCKkk8odOb22rWfQ8fJhl267VXmq31LgSgbsSH/r7TPdZJfqjdt
R7bChMt1wEnBybRlD8kFqKm/rxy3bYbZ2lZCZ3dS/ou/LHIa3ds+8+DiM8RGhf1/
B4BisTQyYNJWRDRjml1ayeNjNW/OtCf7DRIkCJtzUqoaEbIl6i7nZuFdySKpd9ZS
cl6VAdvACzJWLsXKoODMXdDuBPia12hD6qbjBu4vri6NXFcaciEZyoNehq2dm6nj
MaoaTiCSC1vE/8w9LBTZhAUw/MbORFM6OOMwhEOvr4TykKeACnEFu5MZxH5Ydvks
+cnVEGwRskcYRyP9G3lMrFH3CYlTYBAhmAgADcHMGKcpSOj5ZETBvYOkQQgujY8U
aLnmK1+BU5I6A3Zb0c9W7R1mBqG6Y97emZ0I2eIYtjEHcEB2C5vqzHZox7gW/P5J
kJh5rFYmBpYWRM2NaWbgoW5KOxM+GN8L418RjpTBflv8A0+CMxndLVG5eNlp1R6z
04oOVAAIe6Rf0bToMxP3iRVcmxyadiklDIPyvB1ZmK5GEia84WCTLg7WX5u+lJhV
44ToxfwTZaioi1/a84Y0OtXsgkbzssmusGsVYRHS9F5/dFIQi1dMfrk7Nl1d22Ro
wOoPJAcFnGctRui9CKRXkmZ60PphKDtPGjMVmZySZHl8uxQOoAxJKjXxVdqEvAcS
rNUDYiGIFYWZxBla7QHFwHT4RPUoHID57M7O3EYuDQwkbPzMuo4KgX+SEHi3qKLh
k/C4Oged4Yncd2raM1rIkaoq/JgN9PAtO5D2O/7tpjEriqAAxa0HCocHNh+bIYm9
eE7ALctVwmcAHVx8f6hAAsJtB7xwi9yZKp8mso2RqRkQXl4k+Kk5+Mzcn0H8ttia
66gO6qYZVWiwGtyWunRcb1Tv7COi8VgLtzOhGDBeUIiqXtjcezVr2u1Feka2pjRU
AfX/+AavKeafyxSaBiKC9q2EjZ0Gqid1/MNfGoazE97dnKchB5b2pLBRYzZjWl/A
pWOV1ZJw5b+JbsSenw4S4ajYZ4G2yRYq4jdY/aGK/Y5+bWe8NU7fgbyRxjzzY1XE
LIaU2CNCrZelNXAdUEHRdErN1mOKbfQ+r/RxmbLSei+N827MIsLbMaCb8CeYkPMw
ovAGtV4ZRNoMw9rn89hM0499aMB8p+er0Xbi6JWe4Nw8qCW5vudMMOVhGJ1T3BUO
8upStPOttCkuiY5nAR2wrmrYkJQwWAgSMEs9UR8zCfDG2WCaWDsguP6P2/oINnBU
25olN2f+XZTGD4ztfdbFDui/rdqIww4q95HtPgwb5rH57kkbSKO4DX3fLoNlfo9P
6Mxwx2trhhEBhHee09TvH6QRfilUu95bkbyZ0qz/OsLQ3WHkZIPURy3LcFxjUiRB
i4OywSWwE86AdCsNIii6k+RNrz+1SMHXbioR1lwhqIBugLSKl7fcB3KCthhB2M5c
ZGDs0hi4VR0jwVxsAxJXARMcCt43rcoAWtT+xiU8NhWlI4v/sBZc9Rj1Ng72RS3j
NkGcRj/8GkUkG/11oAUbmye8v0xRrn6UzNJE7yLpi+E2VTR9bsBMb3A50ocJVKOJ
cofKgslBT8vqZj89Zfp9ZKR3zByTw7d9RGmfuHPkg2zq7tJ82e12+dtPYkPTWmlG
0tibxYpR7y78q6FStXrwO8E2/F1mTafqLLEYT8NqBearvvA77xYyrDofafRF8lc2
eRth1wXP/zxCRBaj1Beb9OH3lhsqYbqs/9gIN7GfeNfHqKm9YY/RUJFQ8NZcKXI4
/k/YIQAXewq8hq4PNNiMV3JC+VU3SndqJZnNh9/Ia2qXCgwaAIicUI7DiPWjLWTS
Amh+iXGJFAjMiIJnN13ZdFsFd0NOWmxyfgWDJz2hItJqwNe8Fh8jcZK0fiH+kwz7
rYu48+l+2xZGFimdozh/c5nB3a1IPk79shkdeiSpb0Xi7XpXg/NHnSvhaVsJB47Q
DpAuDtgrimsUc2eAzIqqhbAYA+vPKEAmzeY+IxCrZ9q+DxQf6n1MhYqXv4UKJPZF
ySGadFHGRD+x2okSMZVp43kvcMYUHaFPTUOmkPFmDLxM9Ou48aa54Q7HZd3MA4Mp
ulCgHnEbo/JBhHtuI+P1sutseZpkWhdn64CYjNYwxxcjZK6D976fQAwRF483ua1V
Q91A+hU4V/gHdTukpiD2uIHNmFHRjRPd+qAy8c0b+yxFEZUZbRTWcT5bbbZ2RDsm
P2Oxch8XAVT5Z5yqsgveVezeQLqQBAPu1tP4+E6XqRV7YA+Zf7vCFuvvs2nvCQNU
ytPYWc3cDk4Q5ZL32rzkjLFoWc8i3iONWQiNx4WTYq6oSnecKqHt4vpP4HYdXBFR
skzDbJi7kbervbcx2Hgt/MxvpavwxNyy1kH9SXx+l3NSOSwmoQXUP4NJSyMX/Jj2
Kg8AlTvIjW+V3ozII07h4Rrp3UCnVo8lHSRHBd139xhAdbaa/rGj88+DdsQ1SeDK
Xdf47/atFa3jhzpXkJmDufT4nsEYsTsc4/ggzUFl1HIQR05bQISVfm+rk0tepe8+
Z0jjJj2NWbmTiswLR5j+xlKGLnu0MToULso/zXKsvF6DDiGJGuGo1ZT+F3rrA/kn
XmmqO3IibiNJd0fy8hQ7nhxibabqHzZJvgPm/xW/6LP3I2NAUryVQilk+Gen8Xo5
ixUjPYHP3GdjqTlse9jTgwYhRQx5cXyd5OO9NKl2EK1kIq7sPKFkYDoQOhNh8qXQ
7wdatjGVtnIB9hEFpUJ31sNbu4AzyHdVMatdTK+1Hd32aV/lVjTQLmmBbtRb10yg
33/prR2totW6ObFVDk2iVZAdIrGoEkMCsVy+id5Pw0vwHP2dDyk5ct4G20ODQSkO
lyBxZLW4nT8gqGioJ0hSaf6FX6qeWZcsTuKDGrF9cHtfT7jpaUNFKkpfYD91pHTh
4NJFcC6Bj+rPrJpQ9DJlYmfP91WFpJ9uJpTp06xK7O5XIASP7GZ8S5piFTqpYaYJ
SeVMzogPHcAnMx/wfBPcbSwPxDrxX7JZxFZl1cCqJITQl8e0HLSXf2vHsZipUxkR
pK7JmlE+CTnRwA7X7+ZUKgkCkK8XNk6HUhxN1xc/ONf+qqT+B5OKOkl3b/TYKPtI
+yK5TkPvP7K23HcHjWBf1sBTFsQQrXLzxuiCFMt+UTb1kYMACCzZqQLKBkfVy9Fn
kegEfXf1klqyPx6D7AcNXe4TmMr2bYG+SB6wo/TeA5D3qSUvaknj5dqCva6rIRx1
MV3/4hC8yOK0I+v+nOcKeAPHj+HRZRH9BmjEUzoZrdLcZHzKKfhf62UenIKexofJ
eJ7e3zSC0NOqqyM6hZNfL0l5tgyHc69NuNGzVbTXh3R34vo7bbUKOr5fDMnH10kn
Ez14Nbr18FCL3EAV8/gt0XrWpKdWxd4T/VS12hB+TazVNOqru9XOMkSJMl1TAI4V
zJdpL6jwXqXuWx3R+xz/jEyiqjYGM5eDhkE7IqYLocS2iP1X4kubnx0nRrc2oRCk
EwhUsaVFiQ77o0AWLpBfA9hiYmaRs+dDp/eCQ5kZbYKrOTMgGlHRabPzhUQ48FVn
8B5TJjGGabX71Lm0NJ6aGiZdjsJBmLIFlVaGCpM4ykJalCsjoanSUxL+rbUhmmhB
PPDHUcvjvMIgYmc+XuHDzv4NLjlKhn7pwqvqJZuXjdB+DHv7VQYj2bzDlEoLbHko
YCkQmZ2zBY5wxyrCsbz1yaFNtlXDBPAf1FxB3UlZIDe4P9JgaUwpFOe6EvB8IbQG
0b3uLXhXN7mPBB9XkAlhI/CSzjkYADHL6u6/2BNiEMj7H28JEX+bKmKXs75scc9e
F0UwPxgNmhJjc6TMgMY6OZFsbe7SnCR7SEEO9OmjF77xwwh7DXptonZSfgxGEx1U
71qWn++Ny9nrr52fjXPcRCnEG/6OoSHiQD37N2tF2ewX5hzXXslTVNKRIjBo/fBQ
sgOoMWHwmvrSt5HzAdQ2rfNvFE9JlvWhrNL1gqi2mOqWz23oMd7GpjB4JMz8QWyx
utD0cI83sKdfjlxAKlCaQViFqEpoZhw41rZgGUiS8LGU/kAFpzyMvYSIznn+9FiY
nicvripRPZwx6GE95ne7t/MxTECUamxlRWwzFTs761TyUTboOiqVCDb6FKN6i86X
mB08bB08taxFsW6QXHMkVTetONzM6HfkDp3yFjYyeTAdIOwIeEFY2M+E/zytEkE5
t1LCusGskNu10RWO3YbN+YeBtMrJsrGM2AvFMwfl63h6bieCt70Ziu4OMtcu2oQj
AfLivMUUOdXA5qHC5a/+7sVhp3rEwwQDSwEY/ePAg58yv2j3uZma6AsGg1ENhws9
99JjdNk7nSrZdnETmbiAwx+YeH87IJnoAPUNt5kTKV3HAJDY6OrZ+2Zl99tkdB6Z
9pWGJcIooBSjQnZWQtnQstYfseVODeYlv0GIXNN0/mDfMdYX9DMueT1Bt2STyTZa
jdFwyBsgsecF6VfKP2USbiLG2LqOGaz7zXPVmnYTUGFU+yC3s3z/Sx8yjcj9KgX2
pUbTvEg3+tK7a4QFguYOzO+CXykOZGtwMUjr9oT5am/MHSUlSg2m+h47UEHvqnEA
g+gIVo3vMFznRz/yY/+B/3AZs1gMg60tpS+jImBaTVzL/oEC0cnUcrhQeLtqW2Pk
BW9NtLfqx2AYmmH92DpBqMTHiDRmGHlwc3Lqjw5W7FdzQRYMZXUhXjZadfomiqpc
zxO68gVu04b6bLXBPMOenmuliNfg6+ckPsPLuEcxvYwudfmMDo8FqxcSphjM5faO
yuSEDt2zI3I3nJH23sDnChuOIFz9DRJIBg9qAPGxt1BM78GIPKOpRQJNg4BZ8rLt
TW8g+9iqxZDx/OViTncnQxZGvm5j5Iu7Ox+ZWjU8VAzHXRX30zp0AdBWPrccbHZ5
GOmLASxI5GdkhD5gWQHDerJ4VnORWoZw5f41Cp35oBRclP62y0Da3iUAxyS+05qh
AFPaaHRGtCe1nNfKMIt+++7vpJGrekpPQCGzlgBbm7OMcgrDrXKaf/5zYEYGLOwi
9eXIj0dNUuKIs1ExtaH9DMnt5lC77m1vloq4UZkOEosIVIM7p4O5w7XJMFTun2/g
KLntnvgrlGAVScwGEyCfsLVrj6dDUZdpqZszEI4xHjMuWfW6mREmn9YlNKVcSy+i
VyrM9AUuZsfxqJbcyuQzSIDCu1LaGvHQqyLXIW1h+o6iOuySmmnLbg1r9ThscBWE
K8epBf3USSkS2OvW5VnqFh6MIWqoy/QV4Qzox1phhwh30ru0qQcIKLk+Mf6PD1L2
oQBCEN3q96W+Rw7Vdbfwpm+lLOap77WyK6zuaG1mYTquv51+dQiAiPCwaGiVGkxZ
g3WJEm0yh0f2Qu8m8eFgPZH4Vb5orTvKXTITMhL4iVTr72mEag3Rra9MLmXqQteq
mio6nDU7FkXNtZ8IYhZjcFI5jIzMS1f5sBaj/f9srvzTYK9x1THbjXAqnkvLBqWy
pIZI3poux4jPqxnVkTpAUR5zZ4+9nXrRhtfzRU77n7lHwSs0Hanirl/ois4h0L+u
7SIgSPBiMOJLJXeNjU7I+y1a2OQfNnPpXDV1fMz93I46GD4Z//a7Kt2xClciV/Ib
c8XKoNgqcUPCFNAqpFAR/vOaiDA6i8gCOCqIc0kfv5KkNzUttlDI1pZooMo04I+Z
Hue/d5kt0GBGZipXnVc7OCNdfJeBBEcpXADeS5b04vjoYfI9nL/78w4NFfCTVFmy
wK5hG9RZgoFmZq4ogptkHl1EWYGbBDpw6FJEdJR2+Hl1rJob01C3jG07SgfeyF2I
a6+TNiGJ5bTzx8oan4ldOmexzHG4QstI0aF95viO27GlaWfvyeemIi+N0TZL8eC+
BZGjObcyOeo3v2HLjSjW6lp71vKPSDEkmxt50+kvCfcydk1n3VlrJN8K+S8idxw4
D5lGktiq3nyomdmkKdg2YZEYuSXc9lju20bSJc9+HacFogEQsRfqfZuTcI5kcmoB
8J15kov/IyjmL3XKJjERsLK3cbuohFpnhyU8XlrybYu+znHMomaA1xZDO3oHk1kc
GaV+GRyisisA9oEBY4Cl/7XgAVvT1brqqq3PxvC5d7Xjr15Rk0PZtphUKlgdSiUU
emaKzfiwY5irnAnhBfA35eqZUYpzbb4V1mUEMQ9gPDYVKS5IEN9v+hRyfS+uKxLC
n963gxzUtAqZBQzQVo0jbKIji+GF2oE7XyKDDFXZNU+8gKh/UVu6UCFX4DDZA0FF
hV0kNzUL8beWiJgqyVtvHQFn3QfTyN6z/1BNa1WnhGXgnB6aEV/IZfsJSoy8cnMq
SHGeUbgl9r9L4UUqBun6AZQDl9+AgDdigcmFREMgT9FIMk3DQ2CBnjXR1i4W2XVU
Z2emiUszkmcBLzgvzXKefxhoQXnSpSlFiRFGYPd9t07dokJRqeNn0WM8R2VGO9cp
xOF99McUo8gH1AdnwWh0Wwf9pAcnmopq5+kKslFCPcSbs/Kw9asXeg4Yb87N12Vq
ahT39sR0HBtJrKk7bNZWE7YrO3kbyh+sPs7hDu6bZssJNkELThCJYueX2QsTRG5P
rOJFk8oL2mxFtQVtz2Hif36n0n0OgSbZCMGbeTm8xaBofRFWA+uzB/OhyzRE7UsD
hmFIltKgARi5y7uGXQVc857o+c+m6SIguNtPhHj4FnY6HpipgPERRqd4CIPHYHvq
96OrQ0Ty5Tp1eKrxIKH/y8OYgOrLPqzoAuHDKEc/cj+PrngBXhLfaX/mLVcjStcp
o1Zb3EjoxEWAZrjPxALwZS5xJ6ssTgvodhqOKX9vhjhJ5qsOZfyCqFd9rKY7Cn7j
F+fj5SK++dp7KUyVY3fbGqcl5Ikua3hvLYclwt3/8dIsiZZo92T0QX73bjDA3eDF
GVHYgfqTubHMxwSYQjtf8yFjmxv3eEKh5gbaOOy5hC6aQEsF7dy16KWSRKCi+bXj
pqQ7EGfH1KmI+DU5G88wyZg9CY2KhOLrp+xCU0mJODti3xxdRDW02Z6MpY8+gktL
dRXDYZm+NNAUESDPtEB7DP/K6n1eIYb1zpiB3mPXOYCEli1R7Otf70ZDcZs5JzUB
9RPVJ9G8JLMkuZcSgQn5tiIT5ds9bLG4Qy6A7kDzTMMG781HPQcdDC2IDe4/7G/W
y1VuAHxwyOKAq4bmZzCDgHKIq9pbJF9sQN8M2hCqmxc2ejBZ7NWqv3XivtHiHtmj
aFVDvgPjHpwwfCpuE8WXv8ZbAJrLQEWWKBfGsJj7w9/QqjSmTj0Z8jlzrFDV/01Q
rFylW0UkxcvTjTlPQjTYEzH++yXauC6b76aFlzgk7dW/qOyIivGiIh0ufzFWQyqr
koDfVRXkPxCH2mXBtlssv4CfJBeYyhjnS6DK1SOkez0iic5X9JJABb6tMJhRsL7G
w2xBoOKyoxlE55qgkTRA/rOJzeW9iMwkIivT4YSJm+5ZqkP0X6yv7Qur7vwssJEi
goTEbtGZ2pgKPXlls82rMDIkywXe1B5vqAirkgPv/tqVxbhlGAciD+ZB1WDgIyn/
9p0dQ3Ay4B4fNZNi9aQjf8HdAO9Ts3iBYVeSvf6AT33hP2iIkZuXbZUPNQp7ebhl
aUlTjvxR5X8ta8QlB8/aUJMsg0vqnlfLN7QjXqukuqsAhT2IxXb5H1Xl9J9ovg3z
h2wpoPLrY7glMvu0tJgLdM9Xj7XavuCWUu+/Y1u6HaJX58XO7lfAPUSpYe9pdKdi
mBKSUqxna9NvW2wTA36SJPJIb8TlzWOgZi/8k/X3t/m1/sIqfQRG0GkVEgrmDByR
SgbK6hXE/QvENBq4cax/JDEVqeao5wklFaAFBvtEJhzyVsat33OaQiTkpNZiCv7J
mjNlYjNM8e/m1IGHvarNKydHYZERzx78KFoxTbJBRwb4uwN1PAy02OVHTSwly6Uk
LnaMTYotGNx9mdz/bOf/M2cqmamNGe7qav5uOb6p9iF72GfLHfoqQMoPsBIff028
jwCsI3gqxhSq42yZQSjKPncnqvQ1+xsAjYXGgIv2AG1o9ikecXLtwjvuTd0dyh2U
lOhyEclJkYrS3v/ij/vIaHLPhXxHnsKf3jsOJuEZmsmc7Qc1eyKhVAdBp0d+rsPX
MjJO7MojLwjrDn8eJ580sz2Ir5JWSw8nZX7i0QCiistptPgcb4kBoSf8iRTvec1I
ZVUMmaNSuZJlzrxeSyIUunad4wj0qhrHixlxxc+nzoS0YS4z8ThP0uUYvgUzl5ft
+bPQaNCpmAB+rSTrKq9BwYM5akYrZMcIRqpk0BbSgnUQlEaZqlXUnclNGBCb8Uuw
JBrxKUXYmiD9nEnx3qOaxiF2zNmKqDvr9uGjhwztYPk94zpO3wP34foLOtMjVWmq
FLSOlXljroj+uLn4THjYOCb7gG7tZqJZEWSSRdjs5GFJJOkYKKUdOqyLAfk5AwMN
++9JrzxTKsIE1FuQoQwfBfGoR5SycoJ+SQJltJQBAZNHarQ1iLApZjDw7cMLyDRI
0h5qwRS6oKj8ZxNx20s6CqFBvs0aIB8nTOAFrv9LkD2fUXxREzsTFTrIVXVBgu8p
AzyCS9KiAFu6wOBMDfSSVzXf9K3Z8Rocxe18DFhEFifG6I1ssEFvFbTmhrFSB8HP
yAJUy5A7itl1ezBGuDwfuaHQ3yu0RaXLVHAxseCNYx/V+kJMjEK0XueINSWJlzMB
ZXG5Iu5d9mMrB/Vss4e2EliS6qfjKNTMbsFNX0/Zef7eUyy41yaljNxDmuIa+ps2
St4IUHGW4pthfKU8SLTbaYRLryHk/JZtwiD7bJ3kFcyqCsvnjGpgxrPdHOkkP7UH
CfM480oBPaks5eWGl5icPb3swriWYXK3JjcyjAk8QK9kYGA/MIPbhU+LPzQW6lBs
kOb17VxC/YutQtQN1F8q6bSc+/gQggx5uTg1Qp4jyrfwCrNQTtDVDoJr1IfMPyyT
ZDtxkc51iHVSFOD79Fti+YvBEm7vRNA2OHZJoZ60JJEFmVcqRo+SEAMdtAHXcIIG
09fcgHULZu2OFDbkZlBu6FFlw60ICaw52LFoiaXb63fJhugQbemBRmuPZs/QPNEH
I32ixrIDd3jzEKmli4p+mHE9+62+gEmJT5x7QDBA2elWGlUV1xs7/FDwj33ZwHTd
7cenLCm4RLAz19HNQFkJaLkrNa/Ggjli0nnjoYTXEMW7izcZDUIVm4lhNjCxq59+
ovWeGfVcs+1sx2hwhYajRfvAsfdJApVB7eAVyy/jeqn30NTzwsUZR8eqw8e83zFn
OLN1fdzcrlwp2VTEihLKr6T0khY/l50l1tl9FUNeajpjgicockzRHHR8h2+qUv50
Z7X7LSiRLSgPe1HRT2GRTLQiveFrtcGVKgTjNyTIWOH3ei8uvU+gdhryTG5DdKU9
K8qLornWD8VQec9nk/nIUk5WLLvbdbQRBLhol75/QK3ue1lq3uYRxjbwLvsvJ5d3
uyThmRZ2vcZD5f3z6tq5h/GXYPTW36+1wprihZ5twyD+yu/htigi2k5vaXxG946F
TjI3L7xHKvuwPqIBnGBaRo5rD+3AA3Eb80nvsut4S0OQ2yVA2pO7TK2HDPoEk65D
6FdjufbquyWFTPt8whE5w0jPZjpycBfiR3CMOj9RYVmKMYO1HXM52r7bZ+zgu4BG
Nt0EjDCX12qdrRGUTsWs2KUHnvqFdP1Y9j668tEg/UpqDmBBOe43R0ufriUzjvqz
SBmkkw33zn0hL0osRKw+vIyY/b4jQYgY6n/+GiYZvS9y/pMaalPJT1FH0QQVArmQ
Fy/wYUkrERIvMmrspL/LxSQDEnwoyYUPoO4rIlc7rpOMP+GjsAMFM/v37ixlmNrz
+el9wGXCflo5+htK80Pb3Em0y1WXORXG/k7And7TIOsFiTQuMx0YEQ39WiE556/L
yZn3jQt0WhQffiIzNr184R+0igswrUzZV8DSgAWQ8YN9oNKCjeppdEdLoSVOPBME
GO3EWQM8B/fW/Qx6Xu0KZ58WCd9Jxe8tXtQjRVPQgs0wRoWQJiiWMncNshw6x8pv
RsImal7u/CyFOaypqoZo6UBXagdsBCTUPc5YKoMoT9IZSu1qPNlF9UcAmAXOkJlX
JW3E6gBiW3r9imqf9pJ70CwfLPocFLkKZbMf8tdlG1NdnNTNE7SKcEZQX+VhYNoP
d9MOPXJXdWww+MLnB97L6ssVE23xwbQdBwygLZFODK96jlOPtqYO+8OqsLIftKn4
rES10QJGP7MkWNs6RKGJFLp7ef1aa6J5IALphAlLtTi/o2cz0DPDkIrMOAYS22xX
/ddbbm0UkX4akteLalCLRGS+f2L1zcmdp84qFOBcyC2vZkSHndomPScYDyxP7OAC
VGSjnHTh2yqXLA3v9QPDpxJPQ2MH29EB9AkgYw27lNM4MVZw11jw3ykC6p7GpGbv
DA5udxRxRrhlZrz5YeIzs8D5pF+KMLAx4g0ptH0kV813pEvT0Y10OKkBTqIJQVce
zjUETVNt9PDBdRjBVld1Y9UeKDxkZ5dvfVhij77LUNd14AeDTLrM6Rnb712DA1aw
MM/ahaQrgKznO+MeTrloGOkF6Yi8fAVV8VbrGYzVLSQkA2QV+VWyBLajUc3hWRW1
7qpV+c67eip3x5MYlmV+9YPgNm1yk8tqfMwyBkQCpnABU1fDpr838jieEU7p0O5F
ksxPhAfrbw/NbeMGzh/q1tThN8uKmv7DMXRcDsiHCXrlC1goq00CtMPOL68fVKtW
7qLtPThObGwMmpGINIom6g9bQKQpiPSXxQK+xy/vDaQtolxedhxCsbfx7SnxNCBX
phg+jGFXs0rVVC4coZzy2vyQdCIXxjjxgJz8Ci6HkpAQ+mtVuELkSp/mmzaSmQMf
h0Ny5vVvO+mybcfmiysTzuwziaKqk7jZG4Q6jvsWtATnzKQbPOqpyEAhxM5+Clx7
als6Lvp4CUSZ2d47tinD+Gbja8DgnthzK89qOwqOzYsi1oKk+y0BAA7fxCGnP+7b
iEy/u50AX5jKHwRg6tZ7D90Pz3wAeW5qBVO+4G9VobO4wDKoT2cFEkH0dN85d8J9
Ppeu2pFwpXfFNiR2RF6xICoaaZTWUOcwRpeeS6UEKduJ2F7MZ3TPjd1qigJr84Pv
jmLTYi9ECzZghRfRXWSTtUkvIHUIQShgsLXCbUwqZy+CU6kwVDG7xM4QlKaADwqM
2C+xJbHXxYkKL6Nn8kyh63LzKisx6XIdYXjHSGjRRgAqG14atpdFngL2Uth+47d6
ArC1NtmRUJnEa2dZdOepqQJYyQMtWy0bYWaUPU4UEIKVER0UW5PW9olY0GJGenRb
ZAtOY/H2AvabelUNFr4jM274A8dY2l0hvH5q9EgHvKpfyLr1L5Sg5gOKq98IetLX
evSU8aJFQukn+PybbbZgsFzLKJ3d0QaTWv9qZM+O/bimCt3PI5ug9QYtGitoS01Z
OPL8G8rmIt90R5VswkoGTcrgHwxQP+TAhkYGcmVq/2OuwQYtJbj7xOlbiTe99Vy5
0ytkeWx30PR07tXga0xC2fVW4BNnUkvxGtUgebqHUdKcHpUadneGxtmvfa6hcT5o
9M1MsPxDtvkI6fPliU0ij1uEgDPGj4A8AcwZoWq/kZ3yuJ7HypHMMq6jlvj1FpeF
s8fjkfsSq4FvmlDYk0QrL/afPDA8EoGIVoyJRTwunHqXBxLHkSXlznrkULorpkv3
qjg9OIZ1wCxEsjWhYe1UhAfgi72NmvjASlI0dxKi8Pxsnw4opI9TyYhB9Ypgqokk
wYgtaFLP6lLj/8OOUxhheCV7scApWsndBOUu3RpLgj0FJ76FgKLt1/GBHWpccT1x
IKLKxtju5rHQIeAlB1js0tfEk1qyypYoSjf3uTIxD520/hLifCLhIPZZLtZJ59d+
8z0a6oDf20C2b9QdwyQrchgEgXs6FkSu9sctQp8/ypGzKjUfPlvEDrLB8ll3SJOc
MhhqrjVvOEp0vmmx+v2Uz7Mg10OhgvnkexkqVzCwWeQowGhEsJHI5aMDg8c5con1
cVdA4d1coaIS6iI4Ciamvv5R/kOqYZz8nCSnIMhgznikgZoBM2OKa9yAJJ4rp4LD
9UsugR0pwh9iH3LbLWhicBHVTsuoNFbfnsf0fhu64c2O5qcvHrxGQ0Npzywnvuvl
J3E5SgtfhPq1fGxK3OUeeBq51KEU6+WLHiCKjSSQbrQuK1S2zUDZ0aw22IlODgcT
fXNcPAWNqoLxNLMn6Z5kr/DJ3Ko8fm4xSP1clQqtHtc9KQQPeMr8x/+fEvIxki8R
gJMBohU6EQ1Hh5jIY/KgILjN98KW6Emnit6tmyWKiZPxIez/A1VdJGc5QCcFUxGN
ZSvfnGfd3XZi6ZsVkVfpE+km0Qk93IX2d0qaFXKdXisT858H57m+JebDxPJpE2iQ
qqqc5cHb7LTisWvJICxvC3qh+0KYO8IZV3yzSRRr+0I9eps4Hwj7vkLaGfPooEQo
WDHXlFSvUudTZSYoJScBwbdBxEtjzIqgIwMSR3chhAdSEyOWyYb2B57ZMDEjDVQp
4JQ2fHadZErFVBmAvLltN/AWRUqQpy3LfuuLqUvjT9MTY0U+ZKg2Ep/3luan5S6V
989U/6xLZ7jcW/8HMn7bw/SxMc7EnSC0vFvGCkcIvJx1e2gfaHoo1jEBy1oZqxcK
LZ0Eu+CdXJvGqn1rSejOIPztdgvB3QvJMFT1ThERgKPAiNohu/6DqZiWKQ9CRogk
OXBykZqDTBxEf/Q/jp6gPC03zOozht5T7gotzMIhSBqbIGGkCW/BxLnxjPQsuFTg
gcVHTHAA78EuSvdwCbMD+WcQVtJzy3rJpI13qpixeALEPyPOeJCG0oLuBcoWoQ4e
RhL3ZGTqAPIFGUwu/afwoRcoandVLkyrzDTbT2RtXRro3IUFJc1vh6NwlfK/A3Ya
Y+TfZgTMa1My0TGphHnGg0hu8qw4KeIOIEsiDjDaYakln28CfuWF8CohbxkQqNbD
x7j6q2cEny0dhDyh94OPEAI/yM+LhHYxt+P7n2IUDfvqgLWx1lKTAKgDqL0yf7tW
LVM4YvjKGYyTY9aJHgx6dE7VTpIo/a5JYuodhXmLOTgFqoxV+rIsDzkHxs9DRkz7
d82Wpq44n1FsKrE+XE14WfJw7upko5nW81TDoUpDBolLzXcOTAZ85dll2L9XT+ai
FDA5alBok+2tZ7DlkPCLF4eKIrfhqstFgGwwnvJqdGGh6clYqovsIwJqltZAyOrV
UHsjSM7JeEQmivpQAKJZ2tge9C9+Q/JhTFcsmvx792hHzKSTbJXmJgAdKKV7DcgA
idu2Q2kiWHvG7qCRtgokdIczzAW1i+XHQ2DoqiH40AnXCNFNkCZ0aWcbNi94h1o0
0qjesXq2GEmwEOk4l3zPO/B0MG0+5/SR9EXF/gBSK7KlnQBIB8K2nfbwzIgtvIVY
8W+U3dlA0U5Aw2QRwhHv3c4QUt+XZneqWS04NnMI9lkLMBJz6v/bHwuMeSLDcM3j
A54OQAgEEZobJA6ejs6iTLtOCTDh6agE4fsNttULJQ93OYRxesJPdiKU1B5lVCyB
SYXcXr2kgm6PC8sNqJbZGOKtKHSiBx8wjLTjJAnAg3FQQYSOjArCRavGkIJgQUI2
e41/gc9KLcLesbTURcsi4P1B68KKJLsveOANvnnsSDAH/TDc6Rb6bxvXpYptMeYz
LvKpm37Ula9Bm91x60HEwwDxkMQ/acTKW5RKU2icyYe9Nch/iKuHKdtyypYOVdJy
HSWpbRBKMYcyE47b0VwCgPzgAyoV2geDm0deiRFw9Qdtd/Ii7ZN6lW5mUtq+CzdD
+LTrv7fHKil1A/S/IHSIKAL0An8qfMAeBv/d4wqelsVj9L0b0sxHY8tr3DRSzkMo
TWkE+KsIm9DCmPqOlcqR6FIEwa5VuZABUdrDnd8fxwlKta+nf9Nd/uz4xVh4KIRM
LfCpK4M6c2bgpKZT+zt0fm4Z32II5/ooOmzRLiSU6DPi7IBdj8UlO7KFMfri+TVH
rIWYdDTCq2Zr21EVRWJbCND5/a3oO1SwMeZilcKQsKEgmPBGUa4gK+cF3m+zVfGl
Gie/reYJJmNxx7hD8N6YdXjLk6OFWhAJWIng1J726m6asnVDHePpi7U83DEq2lat
/Oog4y8Uhzacl6jSkveViyGQslsMzc4Fvafk1l48EzEQahsptZq2xpKCstI0QP44
eriuPSByGyDdOu/KtFQOukJxCLDg6nhSVBPqHhG1vYYZ96jxLVHnWo9tMyMk4+fS
NCkvXTexHD01RBRdVolKUljacoXqQZrbyMNltN7JVcig/Y5CCqjItqLtOFVx9dNG
PVCGXdZLgK+UP22CgfndfHAPWbG7QND2WWWItuuDyj8uaR7k0PQwhtTSkQptWGW2
xCyTsXKzG9FRea/qY4coQbZMC5vs94dpGExWN9bTgSjDEzvqkS/BuiWxmyODes6s
Kw0Wd4skSHk3J1YwRnzNwAvRPlqbQAS1OQZDwhTwSnNWTdgCVa/VJhxOjwfTFLyg
xB9qWQoZVeWBTgcxA1xrcm+Lk62XmmSJohRnTpk0rYdEaAkf8Eb3rafbTp+u8Tbv
0A5GTHv9t4T1RcW9ZCiOkshOsKjGxw+yKWXXW3PXc3vYzTfIT9beeZy3WOd+W4He
Lol+U891J3yzekdydKqFq74MIDx5wGAKSABKIV76GxRKf4MkDKRfKL0HF0hOxVtU
3GrPRO2bQmF0xGOJ/MQxFyu1v9JAtdUndmtOESjXwGRV5y7kdfkVhNhBwJaCccUY
O0EJ4bEdr+NjPNzWEvfziAlupPK+fDJeNcegpK/Y56V3FJdW41EvzEEaLhI9otFh
xxW0YUuk6Vj+BN1cuX67K2NfMGzXDe2/WZqfglMfPDel39XkRGpT4chwNaMPmoCA
Us7sALsuYQS3kO5AdocnZBjrxm6iglYrivBJY7ohf4vMCmrcXLWE29zjPTkPRMw5
sRoKyJTM5jTFgTwRDswkl//iHRMB60tiJ+U3rQ5cXu9N+vjakWkYpYKOL5t1v3/x
Dtn8KdDTKPAPCTxGR5IiNywuvI+jNXENjlM/UmWX46acREOBACoI/xw61nczS01Y
qs7kFfkTOtNuBj6SLEVaaidgUhR4x/00GTYKpqyRUZmXGcVK8Q+mdzQvjwPWVgne
VV31yCXV3+gnTOOytnIAl05EkGxp/JMREf3qtYl9WKn9VMHx/Vm8SfhgogKoAqsg
LZ9vguKnsGEs+US6ZbBIZX8sUI8c8hbsuUj6q+UYBADpTpktDTPd4F//GH/qD0Bx
mZFpZpfYog29A8mlxmOTgWKlPodO1KYXIh4qsLJO/8ASmddm8Dy6eUkZawXhfoYG
FoJy9ljiJ/LlzP1tN/ca+vZXahyOKV905KKIOzjx3CeFbRXnmDq1A/Ogu7yf5YGq
S1LejUsz5dhxieR6HPFvGjvbIFehbBGw3i1A7Nm72G96312xoXCTFZyT3NNO+Xcb
F9GMNw28kdT3EZnmLcCPi0GtHy/zK1nG/MiqSrQRDqrFSKDga/JKs3uFVatM0OLN
W4YMLpnFLU90uvmrMQMSzTKnvwlqtCKk4mL0R9wVarbyOQRlEOmDJlbwIpLdliHS
xmHlI1vPbfZ33EzpZRfuvw8IlIMBPtOmxhMTh50pY2Af8MieVbGtKK/1lqH8zAC5
wdDb6ee8sS3H3j58lIiezIczK1ANrT1g5WakERz/BjB2/vEpcNKrPVrpq4H2Be9G
UCjBIqzPZcnxOsncQNl8D2CL2DN1HQmV360anBibxEjeTMtVC+Er4jnrOB4vwhWC
4y7uDTyw9bStjWLg8YayWXM5O1/M5CLUtK0zNm+eT8oY2jCI5RDVfRZ0JXq0/99p
QFnTZjkpKIDXIqrsp9A2tG/wvyT7/t0jUufzZnKnaK0n8aNBNwAv01NFYjqRXpCQ
75VUcsoLc/1hPe6Cvzctok9qstVLMDl74CBkWz0g+KKjwH90aJ4rgaxFaE/w2Snm
muFgiAH0T/V/MF0z97Zw2w3c7e3QzDeq65/KNi28WfI+TLktH4mcddHbpMbvE6YU
OOeKwJNcLPm7e7/C+8JmzOoEqtjl4QJyh7EY6XcFP71i4ib1NxLwpSZ/MpvYOuXL
lC9mbBMxV1xhvvOdhOfuQ6br6muy88mVLrNiKcF1IZMP/7+dkbgVypg1Kyslcbvg
3E6Gn/xI+tP5YD9Nrr2puVGCR+5D4cds5fYfsVlbWePw7MlZLKxSbcFZ/z4FGjsK
XkSDOZ1agxbW1uFfC3j5l1OlVsuf5/XpV89MvaxRWHXxmVvfv8kDZyyZUkuGPMd+
I+oszFoPuPbGy9PnqmeohWQX7in0L/4AWvkBZ6uVmgwMB8OlnpT9JFsLleS00og2
98qKiNK0gpShExPYLAZQSIpspMlDtNqN6cICThhg+98ZJ87vARaXrX0v4xC4dB+8
Fm6Dx0P4XkMhCMCF8zRl6BcTdCc5Nq+2P7gWZQgHWElpTnnTBkyncwKmF74AX+cN
g+LKOE6AYo4N9/zuUd5RYgzqqLYiTI7lnoMmlgHZaYYtIPh5hTBZRqctZDqdBwTH
yIdeM4Bd08v8dfvF6ggZ0PrkbSM0cq4tLs4P8FgaFGXCfhRXCbN89kvqEdM0U+7A
URiycHlaEGDHwOqMW1kJo0+r9hYc7tEmmKbAXOIybAp0MaoGGRUHrBLAjTYOS1sB
oMnuUcVLiptf4wRfIGsNnH18urpp+CLsU2nv8+JzghasVEUYg/PZG+xAPISxAWaV
z0830sCiqDulqDmwNEIcmGUYz4+UXVWlxawxhYhZ9BR4TNybWosAI5oEixJl2fur
/GHAZuVogoWe3V6XbH6+ysq6Q0HnokfcTtyawvK3//mAZm3j+waixZYWpl9N9THh
6Lfn61yY2V2wlj01iTTOthbEBGew+gei9SR/Ned4bp6T2uKl2g4f2tPtyDUBvHHv
NVp0pL8zCWOxicxSk7lwWj3Ofv6ndIupCUWeiLxY2ujVF1FI0IJn6KyU1IjGPK4K
xCCyugXObn6Alktf9JYWCWnd7hGvMSIL7EGCPiHdDBXSCReLAvZWDwrL++1YFEa8
Ul2PpI+Xw/iTnrVayODxE2E/0fk+c5Tn1XSbRe36eDejc1PbLawuVzzOCLEJwFnk
R1NfGlRy2xt7DULvyBk6UKcM46h3cmJLLuvrYiN1cRUFtAV9vIyqlwrgby/gmYmw
/yA0vP0Q714qwa1o52h4m3s9vPQ58dV7OVjxIMwkwxjm+ou7Hu3y3vVYcFbrlqPE
UmOOjQZK4+dOCnAPwNl4vHOHobw4tXhsAhxFpYC0v93tQErlPCsh/gVuKbqT0bws
nNrrnw5Piji7HErFDhg8vPpdjMUzFP5TpenBsm4lMJ+xarVliWWItHj2AL1wpFhk
05xnldBrkdIcATYyseqXvGZFYfKNSvfFrsGzI6a9FyL4BwPk04c4CNif+g9sOsrp
oOIGnmsf7yFSzKZToh7iKvHpIEAl7ixA7YEfHaF1u/0+54gIlQa2V4GEk1ZfE1Pi
CQ8VbPBAYpR012JBem8tIt1UG6F7fPQlGnONf1JRJEUMGl9fYx3P5c4mfrw0HpZw
LIi1kY7CxB0K0PQa8UIePFbSW/QrSzqi5vU8ekBiFpJ8UzKUZrwCev2p8I2Gc6/7
42Rksdit3/exKnrLGqiOusaD0xvlNN2qxTyJnjjX9k1Xwp34VbcEsOP9ilkR6phZ
h0NR3U4gMJXn6Qp/vnTh2jbqQmLrF8xOtIdjy5GMh+LNLHHaosU2n2P33LkZQUQs
0ze27OtMDGqc64WgxrQrzOtgoBxDzG0ZTxFWt/1PVhGYabjoSar303PPd6EEHuLb
GS7JldATZWhQut6ITfVqHTplyjM0op0VyNAiBSvKLP0UhTDOwADrZWWAEEi9qy3B
mOrZU3iLdq6z3wIQBWAY5D9QdTlk4idF7dbCzO4St3vhpGMMiBLXK3eYVWMa80fw
Vi9p1XeFi0i22tev1Njj+G8tKX6KzeY5NVWRYcy/Rl5Wmugdqgn1iFQCs382/ILt
qc7y2+/vyz9Ck1oGYDTC9GUCpUWaf+dX6cSVDSBbj7Oe58vOA5MV/WFHKZTGK75m
fOCQiHGBr9A57s0l0JnJPPCpsHDvRoOEkMqc/5H/iL4m414WGa+LHpCdTZKy/nsK
tqLp1qwkDBsHA51Ir5QFfTGpWXd7woWuRm8bgcOLQbSXfx4gbeMpfQJmOwvdC56E
IE1dCyVbNNc/ZSlbJWGMo66wZT5ccI8l2XDRC3A5ettcPipswD+3INMBKE7qOoDQ
cL4MTqu2cr4rgpxDvicgxDZZD47xu70OlYdqHuGj4FidTnVkKGo5tKEe5UOu3KVN
FZs8llTQ/oC4VPsYhQQaBUxckxxRUVbHqMuUpMc4Q+U9bfa2SRqoPZasnrJjMb5u
EpUiHshsJRmGNjbRYr0gG7qEXa0C3PhqctDIodLK8xzLynmG7jOl4Fa3DCS8u4Gv
BQNwpJeuo5S5/eVYOKCJ/qLf+8RfMN6Fk1N/kdPwfoMXrlHYooFRZ/JyrpVtr54u
3nZLUQemY84KVWiVRlwI/Oa/BUjSgteuslWfaiu7ZDgugt8RydbIdIZETsueUYuK
fIDy1+lCJNJ4EOe/Vg1XNdjzEHPQ6h/EiTGcZp2ltde6VF3BMQ3tA5HR6pxNkvue
f+RQJ85+/Me59PlWRp6GYTV9dXYwJ643hd/NiIWWlK3P23a67tyup9ad9bF/vFPf
509kg88QqcOIylYfEzCHn9HwCDKpA1z+WnzFc855eB4APJBeLF8oe+biVfUQkUNN
3MK9idhiTvwzbwSciJECxq3VbHNerqD0Wluyaim+QX1lCAOGzuwE0GEWsCPpKpsF
lTCu7O4B5uUAiE8fVJ1qvY7jUGFYF0+xDorwxCD1cVAY60Bm0rdJfvIRQMZWzVAZ
Gb3R4gx9G0aF/x/us+JPRinpoI530DFwA1WCbe0xxh6c3lE7Bu2yxMgR1kLU7BT/
ex5GNiUAWNcCc/LLYL8JeqQZy9qFHaOD+844IOgUsnMHORTQGj4XSu4QC7PMN6fU
X8aUgKsB3h6XQHCGw466xw2UdUBQQG0KLXdf1j98HNNUlSWPnwaawm/K/wA3b+Or
L+XExcI8fLaEUgc9QivCid4EUIOEps/vH0m5iSNjC3eTZoK6bJGGP2FHG68lGv0H
LiLtZfCp7NHsWMHTRqAQv1ECDPfadINQCaNPAHWqf4YKnSPlcBLoKPQ3JheBQv3R
dL0lKlECWBgzoVUTgTqf3Sn2FmQuBFvMpEdosxxTI+5WdGTFJ+z88sn3zTpWxmDB
XhiQBevGtQWmCHmb06hYy/swoU30l+LCfwosKOliUhdaa6CVyxiTic7nEiRhtME4
FOW5U4iOG9o+A6Yf2c6eoDMCT0+CWpLiVNLp0LVz5YGzl7S9GcT6ruyZfvyh6YxM
50YtF57Ht/pXvJmFw1/dwUWmLxsOIuU59oXi2JjxMGvrB1veUVSQwRp4FFQbRVKu
lry96lFImwbYVxpVm8Z7SKy0F+k/SkTmRMQehCuDyemMvkINgq8eRbkePbdKaeZh
2/IEelnseRGSI5F/FUp0Wir9iFJ2TKKLe6nPuSb6brUMiJEar/G/9wT1EWSQ5qDb
ik23JRa56d2IMgnzpU4CrrKNXa3HjjrHWjJrEzXYXkUsECeO59IubuVfLhzdrKov
jkwSe9zDFnO3HEqhXRZAbZOu445CnZgk8HgnNXJTcWIrGand6oav0tT1NoSH2kk0
SKDziROFHxuJJrVfFGN3ApDEL2qT81u6By2Df80nnCDxkX1714bhMlQPTd1AOoH8
y6nHMh0STo/SNwYbk1oQGYLBruz+wNlhn9m2NeWt7NMrswUSFTf+0YNTEcmmz11I
Rmzfr8T0yUQcOHfekZToQxK3AR3KHoHqK2fSPV2mWXobZEEoRKXuft7N3JyDX2mp
3rLrzPk+xOKUs0W9N6Fg6ZfjLIg+WLINn1/BLBrPvW2GLVtcXQ+zAmUMNLhHEzxW
hQZ2yCWWqC+TlnBvy51SxXTfRtEnRK/7R+OlTlb3SdfHu2VYj6JfzUEfMnlaINQ2
Na4k3YRBKtwufOfCJRbZCu3gTzrTdauzKob7GlI9MsxCwxclLaNM1BS/BjwKZVmd
piceTI80OMgKbLW+sQ4GtEWExTNTopnwZUoO7cKHoBimTH7cY7KaS6YOaN+d5QZk
gIR7Z+YXkf7OC5Ju+Miofr/vKFR3kkgmcSITXpUCMBZibXXVsCHjkIX4jX83k97Y
CM8BXYO4ZyOzDBi3b1o2AqCd2mqQDgKu1YxC+ghufihfP8bo9RXh2IOdgAszglcg
HWY4J91yT38VVuOkhjFhHSZqGOPRdNvC3+QVrHIKDtukJUvI09OLrF5ZFInnmYxX
3yJau/2mHVsFOfM6KQ7no9C+ruAIpCsBcochGV8dd8Yt3VIx+0e6Xu2m7u4ulUho
ZrOhLnrtBY7PPzFP8SpJQbSb2U3P55D+GS9W38XIKFAlyF3szzbkWVOgsu8ijlTB
vK0NFGB3Y/yZliLWFgndEp6kTkg0mwkGkku+6WM64k1WWi6nqF+39t/5SX2fg7EJ
eKoZ8ypEO/t2Tvn/3/ufr/Q4WyiJphP56202btdTznn17amzMPdIxf9WVw6gb1Dt
8C6eMgH70hxQJhcefxewLwqna5fdxZfLYcGUBUpyb3CcZij/jicb3oKNl9ANNi2S
NwYtiZKrRqeKGjvbPc2S6tX7yKMYkI4NkAYI044Mw3q3qMSSYkJT2JXZAT31MKnY
iRCQ6WO7oU33GxC32E4/ZOE/TExtK8V2HC9ta/3Fr0hDuPawu8/kXtgbODQZDbhQ
C0F2cpQlD8jYxFDhp9bcHOR5qQWUG4aPcW3oH6I+hEpSpk5XrRmi/M0VNnX//UYy
H2rec++W8XhWpqx7fewh+qeNWsW6cfMbXl/KdofxRUIeXwmmcQmVkjZ4g9rw5BxS
Fq5at/zu8s0ptJQvOJNPtR0e753xNENOSI0x68LNCj5o0o5PgJIae9PZkvMKoWZk
H5Two1lNri/FhX7/XCl5tI2WR+PkK3fCNmZUW7Cp0sATainSwwSNDjIsVeoao72P
4xhT7b0+s2+sHUTbQdic488tyDGU91kLyk/5d+pFugFXDf1zklYFQ0NIbGZWZaYQ
3M50etKhd9IHpjRANWmn3WWNAqQtr47pXcw8Cp5ho3zojoTbxYU4/+GP5MOyNl/7
/U3LAUqegyVQ9u3QA02XjLxZK/CS2pOGmiG4n8bsG7eBo2kB6liTmPscOyZm6DjH
8Ra6xG4y9T0tInTEGYMvqbl8qZAbIicCXY6vSKiGyBaEaRq9k2sIZj8R6iLuZ5Gl
4m3wau6R/ieMQGo3S+cRU1vxA77RB5nQ/odpz5uqlZY8sJATtwhu+P75WdMf1hLe
B1AkArCwD2sODxebQRfJh++i6//rzsiibClMd0BT2lCoeLcfAnhApViT6NaHj6VN
yNYTNmvVU8cdy9sNvzwmOuiJ+GkSMDmvF94VD2/NfCJRv8mPFHxeuV18Ee8EKGeE
GbIzwPgZka8WDNmECV9JEMstjgIEG8b6ASMh9n9eAkNLYejOydsM8HDF6n/7xBKa
L+EUKMI2GByFQ1v+66HVafl+yd7ptstpjz+CzwGSXv4XpEqQArlVGikbuzjr4uka
qwwCjMgC8MbvvDthfofIWdSpgY4EJgHD0JTR0BodZcIlOG6mo9O+W6AbWsXRSBkr
zRlgyGnDAbpfwiVEw2+Esf0T/X9qW3JYa5N9vq7UcUdWbjDdA0hT4YxR02lVa573
IlV5Q3nEwfo9NsLck2B/qVaLwYWJ4PH4Z7+Kw/+xBtQBnrfX6ADpr+QgwbOe+Sp/
MkV9UG7u/fac0mOGLUruXjoGYCo3u4PirqQ1iq9/on1c1FhUimYsbFyDSo4gJDUt
6QAnyhE7yzEmhjr5EqDQinCZDcMmVLOzlzvvQabIlcD67ccXk/BYHq0ZVOeGHcHe
EDFvI9HMcOvFnryFNReHze/Q2fLLRjRw8Evzs44srpeGIcOEvc0fc0+yhB0VA1SX
A+IqgJ9GInBN0rZPS+YG5t7CUrNzd6QjfkT81RJK72wAmTrLTsOwqBXTq399BmjS
Ps1gQ7T4YTDk+FpdNufKirw6QntXWsZ2X09GPVb55tiEg2NBadXsyq2c3dKyyQOp
7QJJ5abWsRD3cl8VhBk9auElC61q4H0MLxXIzauvnam+MvU+q/DT6v0CGM0kUoYT
inqYcveLQo3nZKmmao6Cg0TxgnVNcmtIjtAp1sw70bYtsFi+161xrOfYNwMkOgSX
RZRu9GkeKHyvZvRfWkuKY3nsHepM5P7ltVuRTfjjw+sO0zM2WbIFIN35/NRRXU+5
rsKfSAx2Qto9DWiaAzZm7+8KC6jeW3rCDvnkgboMwaTnVcZEnxUlTJWMmviozqFH
c6l6+yafxpT3wIDlQJh3EPZ3Z/VDmB0uBTdIAQLk1NhBltqoe75DmSCq44oTJc1k
MPKGD0YrYKCY3P3P3rFcWojpurJiR9E1V5kijwhjYhkEJrLTUmTDMNbIXAz5CKAI
oeBHkocswFIkjstOv3iCo0oaBws1Izx0SYPWvnCNBVaFggeEPF4/XCIIQfdggrWn
e1fe0f6JbB7jn0yfGBPswhqBjp/ic4ci9+xavgdeAcSnVysA1gFy+do5bDkH46B1
5+3hMW+DSPKmroB9h6/racpKnAjLOg8/UIE0+g+N0ceVFhn2FXEMaKK9XWwKgIXu
EeiOgazgDtvN84ArYcSUpU7tqtMqecCikkwM/tmPcc0IoMszXM/wRpZLFzvI2Wjy
Cjtr4m2mxmXvLYROXP9q0ANm3i5OKDEUnyCUEnnRr6uzoYC9eeJaaWxahhA7QvaX
t9j97LFzAeokVeWYIELOZyYZSeEwY96JXOclKgLv0b6oOMLRE2s/eoGi3Iml37ZI
kLUNuodGjkCHdLhAsR+1TdWmHmIV/wNcugKOQ0nQPsJ0fb+lDbpvT9dBzvzqdROm
cIm+24+YlbPM7EJ0xg+SC3qVfSFLZLLAQUiXi+yH1CDv3LmTrwd5+SqbRDh586um
eEkC+HmWNUF2RGtIn6/4p0PVSjaFYdXF+q3/pH5s9nEOVJGok6RZPqY9VZ3wsBjk
19CGfmqv4DV5DgD/5aW7OAqAhPOCla0NVSK1MFtYYWnVLMNT44+rOG0M6LT5LXxq
BQ/1OMYZB4kgCnxuac+tWjowailwJTmXIdl9IgJ7j3J3Qp3g3SIkmpW6ObtMViv9
7wNem1LH4cRvFzNHqPUgHip8CU1ya+mS7vb81YIRagyflLnfKXk5yb7eJrnWAu/N
I6ST29sSll/4HFUcg1/aNR5tTv//Nd6n11xOOo35DEhH4ZEARnLRN/WTasLx8lXj
NYo0vxNFJWS3TOyg08etZoAYQaEBOXDKS+MYMJ2w3QTGgEcxFtMFb+Qe7Z78T8KT
qRZhAYQM19CelzaCBPCfUGqG0CeXzbXykW0CnF0hdnk6bb1ejTT5lbq9n0AiAAZw
lyqzvWgTIMBHmhxLEAQDX0mmhDjH2OjjonSMZMAAArn/Z8tm7CHr/jt3TTsXUA9d
K9cmuL3ZRPcTnnupKQMnLrHxWBNJAAGt8ZHiod/f/VoTabk1TwF5ObkAHOTItiEr
rAMYexfm3Yjj5lm68AnvdbwesC6R1MSAfSYykFvE6mGWGFfdY3xwN5Fk0YwdLphu
F696y/xsiuah7YS61OTjCj9qZ66cEqOL2UIsL9vRmAOa/nb22xrSmN/2YCvGbhVJ
rFRyz/d6lQIaIxxL1mLtCKNWm1k3QMbmKTac6jtplehsOHQRl0LAiXqQUxZpAbDH
TtCwxKtw6ehDlZLSBZ0h6r9bh9yP3kUbWZS2k7IPXZu7DsSO/4M1VQCer5kJkNsg
Ac3e8I1y4425TzjKbmc6mHsM64+5rccRkdd4/RlrMgXrkZy71Ewjvj81egKNbVAS
Cx8D8D0i+Lai4tk7D6Rwc7DlLAv4lhxcYligISLlV4w/zeQXk4dMHUkSU8kFA1v7
XPkGSUAbNAbFZ61OF+Tyz3FKxehqvZFRY2xZBzt5wutzFMm0b8yuJHRQOJcNstU4
qVW7JppulAyiAlBN3L75n7hViOs4kaImJPGpkNhycBOxCXR2GZbCmKdh6moGiqQM
o//3lnDJ0jef2SXwz+LWwqs5EboRn2gHMEsi6DOdL3CJmilfBGFrcBOL80Qb4EaZ
rmS5h9wJNgI3wuXWjnWzXpDYoybSGr7HgNm12zKnTyuk7XkTBS+HBl++NeVYeV3S
0eojIi56I4gyOtKEZSAcoshB+3eHovSnevV64n4p8iuV5i52vk3OZKCwk4kVovRd
BTwHtKRrQEL9lAD8lT3EXJf1jqhNKsrqXtTcXj8+1zwJ/iujTUzdIS+euQqJHfFn
njHcwKmgMR/AryTr+KPR/EFYa9PW2FQfH7HGSdgs/n7c+ntGs19hUBLdhL44p/an
KOoGJflEKC9Iy5LAu+YYRb/5gR3tuRRTS07pNs/dgbCLw7yzh4jibc4MqedUXbSx
q1au+gIW+vPzSInYhErn5hBryGVS8H4FocNv/C29QZYA8g5FxeQpz4mMUbAyPqf6
D/7ZWzBO6Pw9aqKxapRtBfG5mgDyMyNbCm3qb8ArNTsgTc5O/0UpL6TS6dK+0JQ9
vWrx1dSAnkZDifN7xgrk00vkPtZUAcWtRuAAbRqUFd+xfQdYhkq/eZ+vCqaVLMTJ
BHvPoht6xzO3cgCzpEq/DoLZjQngIwXV7g1uQX3fYFBBTMQ+aPTSLSUq3aCYpI+I
Yi0lnVfLerbQwVZkGkotDw1yZG7TaMY3aiA2oLw1n/ZO9k94up7lQircg3OLBDBm
QSy8PapFqonapEtGxC/InGhRqXOmI+6+RzipAwA/VBghsCalOAiX4kIbYXzJytfR
idnB4camxEa9OSM/uMq0bQTDLRMID6Xk9k51uyXdO/69eTjTwqo9h5e+n9/RcbnN
hKpsP9olz7BsrEMCadIo3M3kOGdBxtpIac/B9liElQKD4v4L1x8s/Ofp0O0bvY7b
cOaBGqA9kEyzwE5sGItNTiHyAYI98QcPtAqD9pnKtHcyE9QwTfq0fXWLFz4FbGHC
PTXR/759YSVeHmPLLCiFMo35UFsnIaBIrpGK5gKJYZLUMGLCqWBMBR3Sl/yQ+nmp
vX9U/7c5pIROIC/uU9BkO5p01S0fLoCzvwMmpGVgbYw2s3Fx3fhxtxEYL9G4ZDRz
HboudCjJrUBRVwCzaa9HULr3mwu+5L8sRDl0DimC/wv/Ov686j8TSuiZ5k9Iqf0u
uPt3VfIJT/GvqdTdNGKRdrlu6WUrWd9XJXYQk7qV5o+p5+OgeH1G9jrZW51Lfje1
pYep6AUghDB7FM828NQs5yoKLTlFcsOzJ9L1Bit+m+q69AypJBZUWKwQl+ISWeP2
uTQTteyuIm2g1DjOM/cXG7kjU7yJa8NU5xcimDum2hRUdk3QcnUqTGXLVb9w7Qd7
zKPX4Wf0HQo13eXFX9iR3hjKJsHTdVxZJLIMqBG/rv22Gc1VqUCmp5CLJ0O/WJDA
LFW4G3NzsqpzwfHFBxtBg6qkz+rJjR737nZQDcAQSHjeSXZkA+xt2dsi/7nxrbJF
bspV33hKus3y08O6KGUI5+AcLmTysrpLGkw2VsJp2lrsb4ve18VKbReS+UFL1Dn+
+PNJZolymcr2i07DW76Xt+hXLbgVRinsmh5DpBixf2nTkHVOldGhTIQNEoC1vnbB
dWGVLVkvtxp9Hk7+uc1NHYmNVEbAlhc2EQpWKRxdNZEqFXvc1S63GSNJH7sdMiJy
0X+24EXMYFXheytD2BU3lNIE1DwPTwxxSNjHyqBrkfAu4WCUHGWHA6GoX2jDQySW
nL0I3qZEpCnaStzX6Q8OAAvO6vCUpyW3IzHbXZqArJkVTXL5Q7yJPfU6H4Vnl1H/
kYbe9RN6aAObvPC6uYS8+2Q7pciulHe1M+3TcrT/ibYoetpJJtndPlbKDi4wbTrS
n8PfaZrZOHGy8nbyZNjSaC/lA54rTFllV+05Sola5/wZthbmp+WYKfqhMmiF2Lgt
CP3SOx95ng9aLuVbBbpW/F3nD3zv0CIzVgcDf6UptWzHbd+wDpm4XiSj2HDYIIBt
EhFogb88LliNa8dCCMKUY3DHElU5dQ0Hr6abWcSX5+lxZdCaLUuu1CYE79TCV2ki
OvgvwdHa1RaFIU/Yirqhn2p3vxKFokv0AHJYNiLtM3OJwiy3O80dYbGc2jrN1Ahu
TCrmG9A3pdIEwPcHWP7NLjM6G95UmND4ChhW7eCyXDmRTjmlqGbYufAveLV1ZiKU
wpBfo08j65hhRozKXhiqRN7+aC//JxwNGTO8k4B68zUhRa/ymd3rPGcm0mmj+RnV
ISs8xu7VtHAYZiSbnCRjDvO/e4lVIMjcuj20YNA/gTyOvNXx0blf5axnGzMeIM0j
XAG8T7XltHDenDrlczAWLD+ny/jDp4cbU3c9rVMu+wOsX9OwxJGRKc1Hp1GDcRe1
sV9/1UJXSlcv1zYuhg+uphGT6eaVLEpoK72wQV9tK66AsD/wZXEDru0QOY+KO9sS
e2qMxzvgE/o6s5CzjiuhP6nkLvdfKh03SVyYaSu2H4EP5jIfFERWLE0LQvZVlZZB
m3xnl3mKqdx6R4xZMHYAa3DefVPtn+OMRJzQnF7sIQA2Fwmr6+fQoDoFxvvGBA8B
W724PKkN2C6KHSgQETFwqCC+6sU2oCg4HUOe53cQZqo3xltHlvm2Jfg7sux9+z3s
7moMQqYoZw4Kf+VaE10kj+FVgD+7o66K9lapuqzOWSw303QL+49uukM8fKU+1PoE
sukXBwtUhADnfM8ReFisbt1vIaFm61/xgXrk0huByP8gmkq71PfRyIaQbxo5mQ5+
fdSX4IFDkadllk4qhK0wDd9mD8URkklWeLRCRnhieFfIyXv52+CwFq6oVdsKPZXE
Mn7o7TBukkYwwyr+fPYEnoi0rpNux2xtxhUthRwqDgVTtT1rBqP6nIh4VCvfjlaD
9+HVRhAcaK6x/LgMYZ/DdBcXRVk50AwyC0gNOx9SElCs/yMKPzwup0X9ijUCZwAX
a6qzZNtGKm34s5qjMHI1upQLKEIjThFFnGgnAzzQUwuDR9PjQ6syTIQIbG/RDcq7
cCcPmGHOE392xXi1lFG6g0qc2MG+Y/8ere7IkOaHYKPhq+VXUfmn0g3tAofN9GOS
nYcP6uUdSfPT2PDmNFMnmhgKvXBiQJ7YNyH5CPZSGexxVvIoVI+cOY8fveyav7s4
1YrVtno5cJ1+AD+fnTixdpFnF1yrM235Z0Nyj9r45baiBNre/pXRzCbszSk1AwfX
D0Iwfhyh2mL4p6pYbgO8EiXJtTUevPTBpMZrmBsw5ZUaPCYtluJBWp2mqgU1q2Kn
oqKCICOsgRvM25VLc3wtUNFmsRCFdcCONOoC3kMuHkzBgsuRjdQT7UNZGvUrynFz
zBJbpZ4EXPTbIaY9SbweG6PMJNxN9CkCi8FlcfmD/t9kkGbsQgNxuL4mMRMhZqEM
q8DzVvddq5H1ilLzzctCogkL15cH6TzI2AX2unr31+/C2MTp2cvJyiOwUjH830WX
DXjJSSvKlhJFuJNu945okgr0mn46Ncu38toe/yD2kgYI7rkX2jvehVPajUNvZeOa
9sZ5oj1+rps1A7a3azZJbqOZiT+C2h0PLMDFoDh7WRQrYMiiF7EOM5Uo61TyJeUd
TtN9Y9ioqBh58AzQYfJ5aVD3szAVI0iN5nI2O6KKOBlbrbN20ZoWMQ55CG6mkdpD
IeOLFrQ+2lH1BEY1AGgCdANsw7U5aChIRUNa3Y6GdM/mPT2hN0UG97WmTxGDCm3k
e5fHT/MhqNbp85hNcj6vOlE2xAioQ/7iXhtGVXxGDPxG6X45A4MoXMWuJwpKUQrq
kGkgLQxwlbbJIgucUEUUHL4VGdM3KqYZL3L2R0s5j8dBFyWtAiTSCVS8hPdHLQ9T
2hXcDX9cqoHrM0bPMRIAHcJvFqfEgmbPPmfZ+bvybDuMmU+OFpv6REitky0xfjZc
zdat9vIczIHcDc+VMl5MPodhTRGeduO62yGzjjcEOciwekJcfNL0l8iFebAemc71
QGO8woD1RBUHRd1Cqqg+5zG22MQumx14mUY1nWPF///gGm0Ml4K8j2VGKMZgkhwH
N0uSwGU9/hs1IEqgX7GA2pZlDbk72+75TOis7GdpnNM2nxmD3UTxCymWxCNTjs4U
6vbLgyJAr0iPzQEkxvKAWuxlS9WGWfczVK3v1g85rIQ/G66d+E9RyWiElv03d4Ns
aeGCC+ekVuuEPihIKSldJdMMSeGiAJSCfeuOhjQf6nuLJ/WzDdq+Qb4sW9ZC4Zqs
+xPtzrmieo0Fkuq/mY2+oE530vBpk31xWGD0Pjuh8CscukMA1nHv0DOdo+sAnugx
zY9plsPLc3yxcwTuysWoo4Uo4ZMj6OLrH+B9PcxWFDWYGOoK+xjrCF91UUD+L/a3
u3bxjOqrqFeynYI/e39yWtwittc5o73C8wHy/C9v/Uz9Tc7AaWCAbUNNLqGvgaPz
zcko2b+Ekxa8hl8/w6w1m20/oN98PhctoHG3PJTKdeHSgnHz2eVzO3nILg0RRwEh
esNslSz4IbGfgVmEKTvAzSa0djsmfCmTnXKUtiwkxyX1JpRjeODC9dAoeiLZOOy6
/KwK5z7Vg3nk14Z5hcols3T8mM73L7qsL5fe0U5Qs8gpUUMprpCai4gRF+TcKTOs
cqY7sE0yPXqirFJYBp6JA/9/9LWhWrTyUmm5uyq5BdCp3GBDeizQ5rBG1mmTfCVM
IxEdmEDx02mBJ5+gBsiW43VPo6gDeNJ8sba6voBSfSk6DgkfL7j+WkCA1FCvi8B+
5Swhrln0z7eDv7KRVd58HUuzzMJWOoQbteDfZz9M/877Y2XZeUk0PvWVBs3eo4fG
WH9+9XQfzkLL+KSNyhSHfjR8xlf7jD0V4V885ex0sq1zQ+HeF+e5DwXTPMfIezu+
Ry5ufafGd/tJDxKUKTeQq3fXdIrNuNWtRcdQKZZmsWmxebb2T7JKB/tosT8gtsYE
ee567WxNDB5Vx++ELhfkw6TyK8mY689xlcUWYapHkHpzHw33f/BhE4ycVr1RStCO
+9L2Q6Wv5qjryF+eoxWUSIcXCoPqjBYJQlNnHKAc98DJGJ7e2Z0cDNRauyRS6Cck
LQ5jBfWlMlM4xD++fDMpQ+89zg+YUDabhsm1EE7/TPmK9+9JTClATnHu3RdJLpUR
GhxQAQGmxwjk1GxiGDlcuxGs52nV4fcXkm5RN2kab17kMq+i3MiSnDmZDblJ3ubm
NGWjW+ifGwOntHHm2NRkVSXo4PZFz8A4P+nJ093KWmTnoo2woIa2jYOurF2PBQXq
LTCD8L3eQ6KqrdBw8LEJEZ47MuglbtOjkU7nzbz+f9qrBgTGNBtiogk5xwp4Mey2
OW0vRAFb/8+b/cjzgtr7/ZVR09cKyNN+0Q0X42UvcHmL1izkG6spxRq3rkUHxJKA
7WqhNXc7/SZ2O95TJ2oymSdWaZ760drjnsYLKlGPqcJK2dzOa6ieec3TXTwUH0lE
1xGIdOviXFRX0qA8utCYrPNBLNStXCCfIBZj4obpoERobyg6G5y4LS6U4lWXL+9o
mgu695G7dORRu6hy+OQn6S4dePfHchfp2cjCaugXpX+t9dL9/C/mHDvUXO/8yXub
AesG/EcoMhsbw+717hJIwZ04oPbWMgdAzvbvGpnYx30TWdEgSrJXJnn9JYrhJApi
RFgZl+OHlmNoencW645Gp7U0nMrUCAOB8sC9iLZ3pPQugEchYyug/JO0LxpCJEdz
SUZyh5q8pmVjzKPTZlHg3vm79uqfCcOfPmJr8THgzHPbOCLjjwy1ggygN0lmYdTt
khgTfH8tp0be+UOzXIVRliOnovcZMVZkyvYa8kLL4uy2z4ic8Jkzjq7hjiizuIYT
PusoMPl7aNjF84KFo6RGK2BzjKWkXUQRleNJHXRAr4qOSJ/SRW8XFgZtSNahe0id
1jzt30E9U7dpRjM+QBzcdmuEjrjh5WT1IVRRpGAiGAX3jp5zxLJ13Iwh7aH2ZGYi
R9AWUEJOS37XHjpRAAtjgaxWhXLs58rMQ50WVP+cxdaH2wRb0GvmTp8TnY3beNOX
bYBOODdFqHGauphjC+vWhHLARQ81FMDtLmiUHv0/WCottqo3oJHC7KBJyqyAYMWD
KIpO9VV/7OOqtiA8+sMDGEc9qdbKARaVsRKQNNvCu41NOXo8AeJqJrVm5ddwoU38
amRXt91bXW38Jlm9IRy9BxkDEGGRuvlUz0M3DAMPaDx/xcyTr6OvCc0dIyGgSGOV
zqpi2e3PPFZdndz6YFyERtf2pp9OwV4d/eqj3FahA2BDrZvyCUIaFyDyDcT/c6cR
S49VkfdtvL/huFefFdyIcthq9p5LHf0z080EeWpXyqoWKRAbb4zgLOla8JhKzQa3
AfXncj+Q6yObgH5ZmZWeN3GjuCEtRfIHpZKDkItOt2Jl2PbIDjLzE0c/nfDEPwtj
cQ7S3bIdyVYaJArZGAeTSPMcxMLI9p18VkAYYqszD7ndx2lplGUNTYLUst5XXZOg
NkNMc9uE7qAV55vuo9mRWc1Z9IC2yBoSvFF04/9jwjdwgQ0HGJP8k5IMtQbUxvdq
FfRUHraIsFpXOCd7iOF78t7Nzt0BEznpmLEJEcP7/0331ujWCvLW8KIck0mMFaJ/
uOG/Q1YyoXnoRsKpQGPx1oWHP4r5zMJOVx3nGjdHqpfmOECpbBgOp2bgEquJ4qaP
Oy4wkeAVgjtAv4pMP81n+AJa2R3RfSeWnQdtiWJVNB/AjANqjle6NpckVTCLmAE1
95rU4RmhYRTd4VIuXiNlLXJTESAlc3YsbfnrWA/KUnAsoZGTtjz8g9wixnbBKyny
qAck+Wl+Bde81aOGEPBUhOAEq4lykKsLWlWRU/pXydtVA0f+RzQK6YMX+55XaAM6
7hHS822Ms7F1JdQxEW8G8zRzwi7CFxbABhZt3x5Gf6nO6W6ksZDSdJBSfmtELBEC
2yYfatdix5ZJkfd1HmsK4Voqx2K3pW1NtCJ/8rdJ8v3j9xRwEBxRFEZqI4oJ43Z4
rRIyUrSEnvN5dVWbUMcygIHpinws2QVGPrVgfnQWBwOArMjuawMuO0811nTAu7AR
O6RL275fJIDkmrFP8D4QSy3GFYGYB7tX+JDdpK4MOhxbRqCbaxiKzZLL57PdwyDU
eBDz+mwUslcHW4E7DoEmCBN7so8CTDPfOkOc6AW+pO8zRvD2qtncTA1zA5PVI1OR
+fNhv2dXtOYCbvUyjc1v/51XaAUTelLWKR3WSFsTZTAwjR5PGVrFPtQIx8bm/PSB
1MM3ApoIGktGxGGPt8SXBWjpVtNjX4QvU26KSVNbSkwrAceez8mtcyDaaJZd9d++
Ni6EU4OZ0+Trh5Y8diH4T5rieUJLVbkUBxZCcFV55CSX6rc2+Fz1OrlVIozV8GCB
uogmhlSl7WPogkgtmeS6gRNssYLuS+uBNxRZooa4qwwQ7apvk0J2mhlo3sZceCmV
GCbjMV5fpe6oSOk+BKJYNMlcpVESRuMmn+tl3BsJpA8nXtd/Q59kakHxqjOG3ZcH
gp8ZI5XRmtlXCD1Ts1jn0oivoSiuUnS0p4wtT18zYh7aakTPtrr9dOiypy9dAu1e
/BmpMGIj+Uecu7Ssx9sjib1mPQJ4oniJ7JldgFKJ3YRHf4aFCiqT2e4vkloMv/4G
4ZO/0LdMXZxINca0TFGsfkdebfGG5RRR2TI4BSYMJ55uuDyHbYy8yzgjKbWe8p4K
cJx1wch8ok4OrwFTMgUTZUScFQuCayyBTCMINSCWwGdNW1GWPSMocy+cae6g+L0F
6Pr4Swdom0H/+xDFp1mz1nElb5gU8CDa46WeVZ99r73xHJxQd9kjmCbS1JcaqSyU
TYzNz2XDMwmi87QyH1hXxJjeiu8Hol9Ss7qaJ3JMnq6VyawNaIUoWbltuR5JpPRK
/DNaag0Gei9i//QUDFA0xYUjqUsNLgPtSam4IimSp0vHQIRfdL12osXUD3A3TX1E
EvNvxVxd9VS2Q++FA/7Xg7B5z4EH86AuLoJGxfr7Tq371zjcsJ6j9fLe2lFiD7Lw
76YG//xYbQxih4994OKDF20DRPG4/ruqn8RuqWWRVByJOYZkiMKfihG8rNrYqPCg
zHcrO23P0YJMojTDFP1TJOu19YA4puZdS7zm4/h97oRcOmGQZJIb4S8Oyx8vZevO
DS0KQwIZBnRgKryiacn2cqr2NCQGAJxdIyrl2mQwFQNyo22Sc9wOwrWUTeOExq/b
gGvFhMahvnU9NFhlcXmm0Sx/jlzSmagPSjdfjIQ5QeGaSjk3SpGqyYluH8Tmub1J
2nCpsZUhGMHcZ2YQKObKgtkGyYDvELV6qruiBvU9LBNStfcZZXwI4oWMpxi8Feur
x1cPJ6pugF88/m+FKAjZHQdgsV9otGjuPf/celPBBa9/n8MG4VmsGfMpc+13DFAZ
Dom95ykYcxgwtiTVopTJEHo3MfXqiRZH2qcbbN3e5R+CEAYNv0+mzX1RIJC7kFsO
hZep83Xm2pbzRLINO1zlZav8hW+xCj9Q8/32zU1ag/ZHBpcw52/xuM5VYIQ7xkvn
yAtMNykxzN0+DKKs/pa0SR0plxXkSyHOjVjO0NXJcslu2FCkrA/+/ur5hsNomkxq
AEG+Htt16pI8A8PQQIc5ODlp8E9d81TWjFB70KaOvr4GWz++WuTKrZzeoNO3uYC0
br2Y7ZR0TTS8ol08wmGpM5iJNdPNrQO1g59qsn9+ykw3dyCGUNd11Geg2r0QZO3+
oNz8m2LNdfAPRWpHDzMWBZe6O9FyvhHwPLzvzKbyS9iUOeHps1IzOM9Do20aY6vJ
HRxhzpE4L038hNnBIOKCEZBZRpP/SPDgb8uVBIwYslzgukEp3s2/JqXxZpyDvaXU
BZjuYiFQ5DNq6yX9seH9apc0kDlisAmH2D6iKvc02IT8LyWuZ4kJp13vCnBEN3rQ
GEKei5/MDbpValiFAwTglLg1/3PVkACXR3CvVDEPmifUPvBzDh7kem8rlj0vpJdq
tFsFXybIlgwBjiXdsLx5PBkgjiaR6GK3/JMtZ7V1RbTfSzX0yzsBDoaxTwlw6KL/
+8ywcIZF/wjaJhwQSp2vIIw9D9puMkfytxSoNqK4eqebUbXDMyTTOE6kOkcZJxhz
FTY0bLR3MnOE/exfEnx97VE+AA6V5ScQdDa9FwvQpO6UQJZcnXNcWqFAB2Lpn8v7
kXy4JfTMF0nOyHiurxxmH7w1lRjYp5XY4Xi6RXXX1cw8zwQcTuZSBin6wx7njzJl
9WWYUsDmwAaSG0d8NnVhhr22syp38FnBYkcgECAsnUp8xdkbB0tNHLWMvATLKcN2
AiH3bL59pIEtq74PlNE8/e9DZ/8e/jmOA2t2q0E8kzpaBNcnMqCg7QghDk1ubfM7
7d9S2AG2zIFhnXx5DumQHp5S3/M5tor+768KucmK2EGyBUdlIN4v+mQsXNNAh+lT
cIBa/p9zFwVrcPrRTq21PV88BriBqUMiMa6uQqh+XIDnCCPV9TqrK+XkDT5R6gZq
DuVA71wXu0Yh8POy9pjsSCSyTpEiHcuc6iFB0ivSfu4zjSGsVs0R9Q9R3x1+3UYo
wB2AjXMuqsJxWUdLguqtD/HfwSRmkDuDjZgeECm2EPZej29IqMj1cyPFCuvcap8i
/ILU7YZo62XUhQJWbjhb25Kk6TMks6E6QqMoljQqxiOTXwh8y1U6QH6XHx8TebFb
qSWUWTwoIkpYPs80MpDr/p5dkHeUGywcOMnxw+/aLWJqf4LeyxDk+vXyODqQEw+U
BQQwfMWC+03VC5syZi3AmWkP6V0HgzNJtYtGCcIvxwpI9vYh4KfEy+84AuJ+XXLg
hGDavbfFZGW1svqfFOvd+nmtCMwi+OeBDo24wm3zuqbbM1UJ55i839nmyFNEIiFX
J9OL32qCT6TAfiqiCwS29stnRmCgcEIudoE0N4FTIKUX9b8xXYz7Q5VA3S9Gnyho
jAC93OrL46Md1OWElftsalSWkAqrQhJVXOO4/97uoFP4l2qNrvFnt8EMA53X3o4C
ntheEPYgdjHuByDgeQSlMPcBlncHmDr2fJmUC4GaUDXJTwNyrVTwmW86WXCLU4Ye
DIKuWss8ktJ5eRxuhMNfuOSzb7IwqvDLxMZQRu+0F0c5rwp2FQmrX29PJHi0GOdw
DnGkn8ooqpzKhMrkHl1RM3tAzWODVEn6x/5vkRcK7asPpJzmQstDPKUYqmpbIyQV
/uwPVx45XbvL8ls6UUwc+PbfPdZupeVYhinMtyckqohtf5lIprZmiAxEwaqhKxBZ
uwtnKEvGPVi/JM6zAJpX4yxAc7rSsqEiDBeYzNKkYguKYQGT4iB5SiXdrOna/7rj
H56PcfV8R5Tkrv7nLIahLnOHtKmuJH7PwERebVIld7MWrUoKmOzxCuHZ4dk0/xld
grITj4WoPZeQPZVundVL2Ut2NnAGPxhdd2BQ62l6TW9lFoX6ilb4NAKziJTxNCXL
kf6FU37tQOIMo6Oh0dDx9sZUjYlOG8CBkHrmIrO/BKjFtvgg/kV+mBZhhc9SYehH
ezfDaKkb6QRHiAGczaEit7ylpi1u/vVuIaEHOGq/pz3zUP+QNWD3OuDbw/oxC8vJ
SosizL/5PBvdWvAvlr1a9t1S0CeNfoofteG1VYvaM/mWApdTJlLaGN7Krp6Rs1AB
NFhF5PDqyzpAGc6kxv2hIXkAjsgjmXWgYSpKgK+xS3r0YFdQvjox/jTd7lacI9yH
SIBP1bkCJfWy0MWYo9UnWvEyP1C3Cbkj+B7W/8tddDEsVoIdKRCe+jI4y2O49/dA
suJatE3VcTXqZl2SPnfgoR5RtrNlR0tLGwi6mChhp13HPYM45mOu9XEZ7cqqxRg8
+mGb3EHfacvmBp5Y8e0qtqkE95ptFW59W4L/T1A60xeje+WpkKUHrgFs6ZpvF29X
+OuJ/PtSe8XAQZoMrEGFVIi0yXwCgqaApzVlcSOixu7VGCeHaKzKs7K/opYmG83o
ku1MaNakRt3EhsIoQzUIZ5NCoioTXOi3m+QoQi+sv7+AGGxgei9Xh49eLDmUFK7y
1jSyLRk92bKXqyOM1jyPwtl11Bv8gdBPNsYLnogLOGIT7Q+ZKYfgJLsO1RUNyaLr
qCOo2x5YxkkrGBmYizTSML9ZcsVJYNPRpCKuchhciDfsmdtdkZZ5xPu7jV+kPLn4
W8UyEu8XAyJEiCLB9vgl71Mhn7M/QKU4rBzwWwHR3htAyHZ7Ez/YDW5no1/k3jQb
QTL4NG1GPyoX2v5c6P0jU6uGMW3fED7TEHSjk2z4cEvW0U97eyFSC9XTTQwPs84X
CD0QPQ6VDim0+JrK48oSYx/iKgmUWHr6PaZMM/JIwYuoW0QMNaejDaDNo5DpOBii
4F7vvOk6FyArmUySfeJgPX13kCc2GIFDK5XrOUZa2v6Mb27FGjZ6704Z5Vb/+n5N
oNFAyXssoGLC6+pk0ZTCR6J+Dv+vgfNqAsM7DT2FMCv36+AQcmurm8IwXR7Dxdn9
pDnbPoMznJykdVSOX8ZhKj0WLn/unxpUOIihtdP47cRErdnylt88VFsUGmLKpA1J
M1nz6qEAYAHnRkRLWPmsXWB/487h+cpns3WrxZ+7RX0XhfN4YzR8NNbKIRGTAElu
fjvMLfzCQ+ZzJiKBE77BLWHcu4h9FwUz1DjBxaBrpu28sGj7OLxTSntwRHfp76SE
58cPxexHVdGCoWYmVtMJpoDgnotmbYB+RXArB+leS6IIDIyYmpROUqxE2B9VGDQg
PPxL9KM90UWiyhdMomuyo0tP+jTT7h3POPxReboMF3NTCMgobZ+QZse2dCWAveg7
iok0E+1jkLN0hZQdDmQDiWyK+Ow2m9vl5poFcegloXSOHXVjO+rGG5jd0JvbE0AY
Ym0pnPAYL6WbjPVju1JMIXGkSKXvX1ke7S5CM02IPTlAYw8RFMB8WsPgnjfI37+E
eEzMwJBjLBiqho1jfl1bPvOsJkHVIMXUtlkq3EIR51/5Hq6WLWYeilfI1UpoVgvh
LRdbUvp4HAHGMKmlVqpLiLFOQ1pVCNcRjdDrdZOuBSb/OknRxLShS3Jp4grT4Aiu
IjVbGTwd7qNd5qFCCuqBnU+LYuSk4mYBwdFUYKSkS+b6toTlRv5ZGmdDfGJj3/We
rFki1EPYyUB9ND8Y5/s6lmLV3o3tb3YmHgZ7/7cfmZpI9fXbNv6NzGioiDKVv6qe
wYwtNLELm9ij8Edup2DKw8GllMSaCRV3hceGDBWvfVDH5lQuvZQOpY5Wpe5606W2
d8pHjzDdTBEYwvlXQL4HpV/yZBUAw25Ze7pdKYGf7wADLm3mPnxMD1+5eelSb8AU
vCt4qoSU1sBQS8DlFZvEoKwjstkyodAaLSD53Es777TtH7ZbEJ2CmVVTK68l+c/7
aqAEnGLD3tskKFUu8EYet6BM17GwJWS2L/L4TcCB6zrZMrrk1FLc/JyYqA3kwh+C
w4oUefuLn7dSy6ATqLyyjVoFjKAHp4A6K/FVY5s8duwkY3jVrkLyH3IXnqskHhaM
rmkMBZTgyLg+NBnIeGtZQ94ReE6Fb0IcLKO+8thtGdvBj7PUuooIw9lpL3MPhlaH
4tUw/odoeNIcXaB3SUHFsy+02+HSuGF+M95b+dVO4wfO70NOMJ21oW6k4bo8rZoQ
QSQQhsceSKeBxeEjczN/vX/oKEVN2zPShaOowq2e/NqhjM+YPmQR6oJBiwNs7+CD
WXTav3nHbehuaZCy65oevRnW/uoDsyTLB4XdzzCZltLjJMkZrTqabTRnPRIWIk4H
6z/Dof3kwkC1LSUZ70wHJyTuLXkbhPfKzam1WCemRW7fl0Y6PK+OZY1SNOCZz57t
/UDDl1TojJ/BJDq7Jl7XiL0EUYh4suRtypyIPBufNefybpwJOT2qrpq0Rn1zTr/s
cKyvrqtknuO5gIZVeZRdaEJgy7XAmxwwCza+dWRNWwXssy3FvgsMNMcQxePBYbmW
hIBOejRGqqyFY8s41lu2uYe+M+yycw5mNa3sVpFL5JkolGpYpRgzsu4YOnUHR7zF
IbYLdGifvHq/W/B9s9ikw6adRFRumTGrxaGHQF7IyJEGZao6AVjLdKx+ZOtM3Jru
qgviHkZTrbXE9IfqIcMs3GZzRmOoDgC7Q6ORF3BAemBnoaAwDnMlZRdh5jS5+xoE
teBEcvSSMTjHRP3BJREQ+p/TwbiaEio1FTHEovtRjJs89LQJ84QP/MoJxPwYvbEV
C6VHz3bX/WrU2eEoiwxYd1Smlx/wjzZswxm2cJr5DVLgQ03wIFKWoFz75N0Ko/eY
mPUxZIwaC1EFm2GhYkvkgYQTccBEGQ6zI2yq0suxfhEipu4tHeVUiFVoVVHiaUrE
92ATc9WK35LWBcwUmJuPEgfg+Jjpg7TcpOlRMgiNbtKaqOB+LIaOLyPLAvtkoeGb
pN9zSMQMcAm4cyo3VuzRu5u+4DTm/fpn8UD5GD1me3mO+XAV2noGbaEFqWynbro2
2yX8BQaDk+Pc/cazskU6CtyPSAYNgE7LUjL/YzzDBzRl/GhGSCj0FY+Su3jjH1UE
X81MSAQ1aLq6TLg2a031KsIidq6mx45EkV+f5YlyRAgSyKLmRbP0ddp/UxTkFsDg
6uuDPRrpfaXXfRzpBFp6/j4U8XCE5DnDGBEr43w99xe8wwpscazPcW6WoXIZAvIF
TWokEm1v/S97E8B5fCl5VlXVan3F2rVYNuRB6+SKtAsAb31jq1+OexUc7UNBKIEb
KpvBhHQpcV9iiwSTHRQ+U2nB2d32NpOT9KmizosaYL0YXXiIt2pnqaMSkLP8lvGK
GF4sUJuU7xp5dKZU6G2olUmBBaAGPPa4kkLTI7iO1Dg0VME8zhiy+c2e23o2VjbO
UBviVyBZ86IPeM9IF9v5nVJll5Mpej23i8fzOlpdDKBBkZ6I5k3jDqYPqinTIdAJ
WguRNTh5pYFKBwR4I/gq8eYA8G9QKxNa1eMI2iBemgC9s1phqGbOF/HVhTFoyI4n
igqHcW4N/HaFXfBNrOItIxJ9SbCCnOlpY4kSQOJY0DhI0ZvQhpxchIcD7VTP/Slo
z4W8pTip/XeUpRp8R+WEuMRCQHMjDBVnF4ppBqGpqOGvAyrs5SzsE9RjHz8+KsJI
/5ZDmrfX/st6L7Z5tULmyRLI4FO3wCkuqBHVWc0/mGO4ZtM61pFjkFMKbwJCb823
c/XfN3APvc0gYOhxkyWMjkXcHS9cAS/AvI4y2iD6CFBVVE5yLRNOvWynPuKWX3uR
ZehKzhbmcFGP0FDxryyvXmeWCQeLibyOYei5rXDIF2KtriRhJNxzo7AmnushMDRg
3bpTf3lgqQX+poXLwoDQxicZBcOKfnKsEBF5lpO6+XWZLQ/xNPy66UfXpwi9g2QK
hGA3HKWDLAD8+ITsg4z9D31G7S+c2znLMQ+EUrfXnzEBuPm2GglmFldDYpGAnL1+
9FR+f2++1eSyWhStBOdAyoETWFFuRaKbEmjc8lEAqv7XML+Bz5vqDbb5kyNtIXXw
BSqKab3WUTPnaL4bVOGmjAEDcomD26RFYEJmp0/AM7EXfixk5oxHSeWmBIe7OCtn
DPxcxYfmarRLw7i2xsHvLzRKpKHzMU+0eozZzEw1muPUopLwxjIT8E4FSPv/M7ew
Hy+btwVVl6hHr+oDAw4acpEf+ICDa4NesZEuiGeEo+F41+ujli0SRO+7RsPsVCdB
K6cLzzBR9PkIdHbcBB79DZwhh+FLUkw5Z4kVoGmdbdWEHzGyRYqiCJAruAQBGNDF
oeU/OkyWqO6KyjlZh7MPvuvJk91rZqZIf+3Lg8h4jWILHNxGeVnUQvz4p+9suNDS
DmfuyWKxcnIzTmNdroRzkWbYrGbirJGaRraCSdOA0I7ySV2tOC7YNxIhe+jSrLLH
gzOChW2ufn/xNEmSVyl2vfcW6StJ0AVokZfjREUaLUQX8DkWnz51v83w0ArK7INm
96ke0ImZTKsMWkOfnlD1uloNugeJJ9Gv2HmvBLC4Jwi48LvIqKjT6Fz3gqQUZT2R
ILHcQksgBCtrL6xFeQ83Jqi1EOYHKIXCzCNoA+ggr3yp+OhdYZMxULIrknulZxZD
vjHOpgTJNMXZsgDmpu6NyFG+D9/t8GhgWthfJXfiyPef+XvwsIOkw3CbuHsT21rC
woy68+3ROer727ycSbPaOTOs+M3+YdLSiyeyEnL3pbz+ZcjxRiQpZP3HOfqrkI83
g+Buv9X3gBNFEauEx/cwOdpIi5/zqW6EPuzlygfnLdm1yVU3kltsZeiAf8KhcJax
zesdO3ODn21F7d1kaz6prO7VxZup+6sj+gKQL453oOdg9JRWb3c23W7gwSNluYLE
Pj0otHp2avzlkJj78+pqLZRSTxaOlcdjaJLhBWiC6OJIUbw0O1qI0exMdRU3lIhd
L3USZ3t2Y8sCWHvZxNpn3VE3Tkkd04YURbd1p5mf2wT7Uz9a/NhLdQG/Zl3Fj0/l
8w8tILtpUFCeFzCfn1COlqm15KXSsGJ7rfaMwuLgeYJz+z3P6m0b6rjq8L4qiYex
8d/ymg/DiTKX0FO+FtnAe3mocHIo3x5a8TrsHW4Uv/Sbop7EQil0D/nJrs3RxFS4
haU2CMgHJyak02ytsdSparRmf1cmlnOjYXq9CLVLb8xudpWxfd7KmqcJp3Mkz6dX
HncfmDot+kjPjEYg4i4QShFgO6Cy9Wvc+F4RnQCU9EDcQI4z6VqmtiS59YN95OLq
Ghw3oibYyBqHsieCSy56U8wXpUwxSMxhsiLwrf2lmnHl8OXWaAH3jyfQvaGycn2Q
SIhhMUtPfEIAEwe5SzU7j6u5mD5i7DsEo8cOul9iu0n/aResqgwxC2hyjEIJKU4P
ML1CM3EN8XWOxaXqkRVpmQroX26eKLNUXAW5WOeYD2+HbuEhvO4rWnILG+q4icH4
o8iJTTJgslCP6spAKX+7zteOX03qNI75EQGGxRtJLga2IrZF3yTFPco0/AUJVH5Z
bhkAm3WDG2+hCCCsxXOhXy1uvFn5jD0vWaFn7jXX/dFYbEc3zHfqv4hk2rMv3TfF
70ftB7PFAvNJHa4ELZzmx44u98GIMK4OxSOplwVFUse9Nfoooga7mBEYitlK5wKu
ysos31MYkfaH5nS6BJyDrFh+IQ1I9J55Hd29Nea2xNTsWe76zDbcfha+UlfiPswd
jgAR2ng9kWc+8RRVmWp7fA9Js9ENyGY9bRaQ3YY0knKUTL7kwvaD1GNLoTCQMyH3
R23mnqCF1rXnsDCLdBBgPjdwp+OQrPJjwbfahEcrMEZmN3Ltz/ynAjBx6/BGip2Y
o+L5MoN/a6y1jmZaHuoWMp47QGnGl3B0xuoX6TkDlqu8dfqtpI4GbrIjdqp5IY8P
SsYgC4wjanMCBkxAopck88y+6Hi/aU2u7JD7/MGsba41O857p43fuCnx3ENOpOf9
e8Bv2wIijFVwR0NGFskelycw9JM0cvZUixkFIEWOW5VVIRft3XtePgx97vNwx5Bt
e6qcT7ZaohFzA5UzBTKta+zKzISjSOeoLLZdFFMnVkrr6/P+4cSayJfnHkFCgh5N
mtWo3SUzml07vf2tzDpsWLvlI70W7DVbD/s1brh2FMAoNx8S1Zq+H5Lv9fpPTA4G
DmdNlRg0FpmmAA2A8mrobSr4NnPeOhkt12Sm5XE/EXNeV/BoQbs8iUhZQ0OKNlm7
5onA3ykRVSddCQswX1w/VpBfXSIHjhMZ8igHr2cBcEbdEX2qhLFJssWsIryZUi0G
udlciICkNXLFO6sZJRe3WL2MUkkJS7BapTd6DR5op6FxVoahp0ay7YTzp0Gc3JPj
nMUJdOMx897GPbHQc4MpvhD+RpoQqh2dT3XRRUkn/fMKzxIVlXgMWogd85Y1EqNR
uj6JOvsT5A5hXxV4RRkeOdB5UjpRnZYBWloLmi5Qi2Bk00wCx7XByGmdMXLDAzXO
xiJ4hVq+2d+Fq/2ffwZZ7o4zk3O/MNzKPP+MqSnRqmGMDL9S4UQtCI/MGjrc6KIC
Q9IqWJ8vjnn8Rhp6RzUgf0jpn/0CEhpZuBKh1xn5MkNYBwaYP3oYqG0WNEhxsKgd
S0jVini9phu/n+/arWGv9rIOz9yZ630fwlqgJ9/3PGn7QS2BbLgmzQaOHEfaa90z
DfNMFTcWV04w08khD6/tGJfYeVu1Lt2H//iCvNK4Fkt8vQe5sdWmce3aNvGnv7Xf
9RYHpXbJjKS9GusX9TgzyVl3NjoER4Gzk5QYzRldQryZarOntz+zpDS/75HnANwZ
Sw4QttBSZ+9zH2ea/rYrfRjf4VEVErnmxKpofcJ/qJ73nqJZYsWgtl6c37C5sdte
APOn7tFrQl19jJj+KEM03NdE5vi3D4QR3LWd3OmDE67FEEpAQX+ae7Sz8xrChUus
tes1gvTmBcs1jvGvYmDAk5pjVG8JrTDvYqKVYXANCuZyW3D2c/JwOPapkKRXPe4A
EqD9cZKPFMBIvfYkEQ4G+m6HF910a5Bl5H2irJesTsbiYA/12ufAdfQuSqjExEGi
+5qBg0KImAUhHXOzCdaxIQJFP85ucS1IfUPDiLInkr4KlgN1sxjXcrMxgqSvdGQC
hEQBm57QgZaBcSjFK0YPP/UMplfHM4aNoSeGkaZHSnlIoQzW/bdx3lTzQqibtYcW
3iQ0BEo9Q4SOK5DeyFoz+P7wsm8nIpDcAebL5leOntT8vIX+KzV4TEkPsGEBJJkC
v6bKTMDfdxPgAPyMyHnxkMSn0b+2AcIy24xP9L6Izcqu4OiIWQakV5rr/AqOZZRw
wLsZ88nkgJqd07RUtmwlOCtxKlWUqLOkXvVkQfvIRsWZHp/5FZsvCFjPspLdtqcn
xcmmKA153iVCrpkD3w3BDpzdHGRt9vcRSBn1ZjQCY5OZ8CkW5EbQKOnfTqS+ShYQ
d0rDJwbh+HES5IclD8r0SXl/KfSYISaCaVLBQDpr1CDHr9FeVVIXScDB9Is8wxSk
jMnajccNsNk7CutuE50Qg/QjursqofwcKStmX8LhAXHLQILQ+3wcD8S/o5axxsDV
dIE4FzFQHuRMRdGL1lxzP86teNwY52i776dWx3aWkIsYAs8b6m6tV6SrFGhXDpCR
4ZP83WiCXmH57mrYh93lZFGglFJN8fvCR19Fst4MoYL3+8XxyfSvmydjYlEed9D3
cshes9qu+1j/fbXDIiq1y+dqoV3jkelnjmPgFSJcNJnqTlQ/E+j8/j0IXs9wyFQu
bw7YVk9FLedfL64bNDKeesWPeW6duGBTyMfCfHZUay+C0rekV/9otmzCpmcC8yVr
E7QxJWCJ1ECZVke4EHo+Rj/565wy0oUeyFB/06oMxOmmIrawiImY9SiTdS7YRjg6
6bT6R1oAHJyyuYvSW1nXdOejg932pUEeJ3xe6tcO5YU+c4CDH0pI/ylAr4AxJ1Gh
JM7uIt6fZAxXnpobjWblXvmapl7ALAi/hhpRrbvzlX8YcpkZ5XYXDGoOS9ikXEV2
AJAE5mpZgc82pN3H+Qip/ZY8vEvbXaxv5tjDEk19HzhwAi26/UsQSvMkSgqGGAGS
YFf+SVkpGL0fv1Xqj0d4PXdJkaOFFIivzM5Qj9lP248kTipxcPosLuDdjF5eL/Jh
Pf+c+0j4XAiLxeAFGA/cScqizOxNtYdBKIIRNirERi1vSql/klRjG4e4ntIZKd+8
8rw6vhfDZWIxDzkvC4dJnEVDJESKTPyy0lopazUCoa1hOYIM2qWTRwmoOUptKD93
184cuaG/Tq13eZXvl7ZHTjpKzooy0m7Zdk25YzzvLF1DxPS3QOV2k1TnbS7NvGJ8
RlqDEkFpUcPXDolZ2vjvlMCmMUXjWDUoAgfUwUYo2S/wFoq6wmI17sAZ0mpxfaAB
ArK9+UJzH/PwuHoFTr95bBZets6HatcFVIdgWpoG4Cd0QBEECpbwGksubiomi6ba
gV7nfU7czKVBtJa8tKuo7C7NcneLuJJGtTNjoTh4y8YULzfUGg+jkdaVv0+y7mJ5
8hRlglputoyCJIm/TU+QUTeFXVKATe409Z2s24ymtWVLKrluXJS2lz3PRahgxivh
dV5vxcRj2WUHuA4BDTEvxS0WA5THREbIv8/fFeBLXjpZHFCHBzyjGS/bHnODuYLs
lYqQzab48cttoatPgDmZWLOfY2SQxv7x2wrMGiESboEjYX94RoPscYYr0Qewbg2s
YFdoHmuqS+P+Tjfxmfm17641X+rdjME3+rYZr6q/vIg7Yj2FGIGSTnye2qtfGgig
3lLSPjRM09Pz+YzbVAsyueF+kgKQxYN6CmRFY2m7sek0CjBxsZn2+OirSuCXdbVL
8EgfAMGA7PAGNOAZwagJm6R1Vj9vUwNNFSg9exjwhSZfYv0Hy2PzqMzzRwugoDti
00UB5K3bAcAWJF7XHJLVUguGzjP0mTX7Yflagc2YZe5gS89CS4mZ4OrdLIwFRYB2
OOGpu8uSiJHliFRhAmLp63B63YuP3lR/MDXY0VUOgVbyrKtbCVhFJDixEHZEgQZ/
oNGsGg4/rM2OXUrrc+9L7qipJiL1iIV4HgGd/SB8Tn55qCqFovsggBu+TYRvb5AS
KSQuXt5XrnHgxUPJ8zybw7i07ETJsZC2mbu6Mljqf1kSzk1M7SKBNmnEgovrGwv2
aQG0Oh70y/gBw5pjCdANLIrDoaxun/CGI4IXQuCQr6cDWZZ+IH7gfi6DaMEuyN+H
WTCmbM5PlacBLlIpPjXDRV0I9KbqxZvMUqn+7aBWgaIzERXw9gJOvFjvTQpKUWCY
8Fk9Eo5vL2Wer6zjLmdCIoZSnxYDDcYTrc6OPdZmrcjn/kymEdSleQJiaBa7TzK7
QmKuKhmdVb3Yl348A2JFkkAx5+Sk4eMDnmtdgPVd09qs6zFTwOYZVhe03GX4pZrk
M/akdF68uswd4/qIUau1Dhu1goEQa9evtAwn5xsS3Z/FF7T/xrs57vGkd8mhrX2T
P+EPXg8c7pB/OsxxEacU8bjwa+r8tISqrmZmhKFLgOaquX8kdcA219G5vkDa0FHv
NUQBc0P2DczPw+0KBQ1HPGvQS31T1/T1taQTq1sMdXDsyBdTcEb0fiSdy+jhndtj
/+BL0/gTt4seElc6PP445l7V4jBuU07kEBgJUlyGREmoipdFdmn6m/CAExpuEG91
J4S+rkj1pSv1wn+9eqvRUY752MLQcQMX6+Ekcmm9QMIK+DOZ4VJZBqprKO3grePP
gXE1L9Ni8jfUxv0twVnMKTfddM9+r3IZ9cXnOe3ZO+TZen05K6ol8+VeXWO0cmUG
i81UgxobnzctKueO3XmnDcBjvFT1beVKqTIxyroG3RLUqf/3ULuQGclJKMV/VZJn
0SpwYefxgpuh5FnOAufKqZvMqFwdmWUNUx+gL0qu/Xg9PT6fMownmCqw/yGNIvyF
IV2127cqIqit+FUwhf68tyyXEuHEm/GWolAP3BVoONztMzZDZPMVmvW4O/RfweHo
uvVAT+RGVuYtMQ041c24HI2/jZlZS3WSWLbH35plT0mWtQ2mZLhv3d0YhHhkz82v
wVStrvqKx2vvsFIwRmQUbHoZPDd39q2IuwShEz3fSwNSZhlSFf0hizTSGHfq17u9
qX50hvAgvN0nyssbt2lgJ1ZOSjzHs2nvTFLpJlKBOHWf8h4RRYnLk4mzimWyHRXP
BmxBsPQnMQ3Ca5EKs1dTghcJm3FGp6Jj1xwAT7ZFW1Hs46HPAu4uLiGMTsPdjAKe
o+L1djgiZTTOeQlBtDKLwvxh2s3ZFBUvq6GZRfUuB/FZKzGVHqn7LxcpwUm5l0gN
Aewuot1h3d5w53IAp8X1DQIJArARVAW2M4RXhscdVoXL/Zhycot1ZzXwuWhrhnw2
T8KP03OauEVwgmBfKXNQ0x9y/08wjdWA84n9zokeifqNiASQmGL/v2B4k7XFInCU
cgc1z2rSVFaJhZIJOjvFTYV7SfBgHxsk8SBvYbG9NZBmPfjTPtSbDMJWZjIeZeu5
+aYl2epnOt2GKV8Miayj74Q0sFFSIJ7BWeSsElaP1rv0ab3S8cgQEEYSLJyxHv/n
9W5y+mbXK0tQf/uM1nhkgeYQXsS52oSKWQgMnA5F+03o1XIpVEcW7WjaSjGm48bD
hK24IO77IXAHKjAoFTnFNHlq7LbMEflsaQefmDCFSY8yhTAI6Mg33UG7qfETKTUd
/VlOZ7Bc35GCuaLB1+S6/uUqic2GWXiExB9jx5uMrRiLvPSibaleFl+lX8ZOysPk
eiW4/sCijN501G/BqBEqyOrXtrBOmPaxN4jVa9gyRH2Sd+nFFgJXS65q8ZdN0tZw
L4ygyZ/fBGFDOeJ0rii8zi2VlDwxRuoCDZudPernxgd689MQefhghL6zYFh3jqnp
rqCXsERkinXBukUbklJmVGLQ0XYCfpZhF7w7xFYxqae5pnGMCQFcx3lLZuhhnNyz
/w6DeVlzPydFQwe1fNVVLm8MoVP9irfB+LU16Fo9kMA0HGQ5aSMFJJ5/ehUlrJnk
GLe/q9+ODNCpgrOfA9OEtcEIriI3V7AA+MZMCsVkITZaJudroQvKQyqBQ94GAvdo
+mznUYKLWvXo5el/Fj0KFVxeWKVBwE081Vex+EfwonndyXaUzeSRG2H2YtgKFdmm
UGaD6FIR/jY068sdZJRHODBcKWvqBBhWPvxc6QKOISEDqnTlNH4tDeKxbiVVTkqr
bT3hcIcUJN+8FLn/V5UqP0VyXYw2Z3tPL4j2GtWu9T9YnRY+IV1nwj/YFvbVHj8U
MA6cAiXAHDNbFfDuweroqcQXNIXudQfWFP4pNjWpOYJ5zpfCQR+cU3RkbQ+9VbNg
AVrkyOkDz1pA3kPPb2+91JHqfbM5WRoI4xY+x0od2NRTBeOTzh9rZjQA9Ujl7C/g
HfAew22ZVRtQoW4XbvgS7L94ot8j9AikvC9OePQzhoELK8pStck3qWSnkjmFz3iE
BIyKyNYJHTAeNUr3oC9aqaKUEsvqzISOmZ4vUPGX13jXse3wiYJ5S+AvNXba+ZKE
g2KuIGbTPPI9ghauoFLzV8vPPUAHu6e0994OE2d7QO5oWdmd+kLyjm9+Cw/TheK8
vBJNR2KJH554LT6boKFSPfQW0iEtKJefXOOskZKfXFyHVMTrxt43db6VySzCI+rV
GnXG36BoD5PYrZWYKtq0vMtSXmauwrV2kM+V6GsjRMJWs5lS4IrhYFgG4QLnFv8m
qmAJxw3xQNcKKDkKrqkcjLsMdxG5jhicSuYjdw2MQqmlfclz+sw/uYIqw4NGTwS7
wvayWxSNdJjxNa0NlKCDeZYJvXRoiRvgQ1za0ZEx2ihNH5q/tDAWcdHMR+C30cED
wS0gk5xmUVf+gXRUm7OHxF7MlSGZe/y5vcvzGr92u6Dt31EOeyzxhiifZIXcTkYt
i9NO6JqAcCvT38ZcrNB0RAGkN49ADmuEvflAF2PcHUsmqZQvuhbr8hDW1I2PvOVB
v2tIFmgnJjKchTY8awkhTwN+JvA2+Na/HC419RBh1jJfp/c1ObkBwKmtO3D0rpXt
3XtQhJFmF/3mwCmJjRVtIdixgp0dyOfCLiXXEnAyhGuugeTA7FQ0pwarA2DUbPxy
fr62O6Jovh+dxPoFtzgAqm4wwQ7cjzCvIuJJezD6sGdZllgqfO/q+GE8B7DXH59w
z7X3YW91ucfsM0YWV6j7ehaLSjEg+JjNmmCY6EHBh+dHEOYtBFtdEVJnrdNNacQi
B78xzcR+dfBJQwKapYnMUIO1YZlr4kdTlx1bIRAIT2TSUpjoJiJesx5MIJEegE+x
Eqq0p80/lltji3ayb83Ros6URcrkUm02RmuGLEQHk/yLGTnJ+dG4VZHjsLauN8eo
34fWyOX+G648sy6n8ybN3X/bpdbPjnLSY2xkTMAZ+7y3Tj+Pl/s/3AXCW0tLLJ+o
hR5wtrNSRP/ry7dUfawxnfLnnIhvSicCIKC4yOOWXxZMWaL1tKd+oSNj2kuZv0IM
D1jH2V4IdDrZ+l1immHWcyOeOrZYNCOcPz+GFsTase3HtLlDY7Ut4+p/5pP/TScI
43dSwlkfEJW7ivR6hiUORcVx2YumsClua0rMvBVMYmfR6NyI9xE4IVbKRebGpN4J
1d4VRfgFe2y+6LkqWntmAajE/sliu7OK4+7t0pgmB2h0MJvaUsx982zIdGI1C8Gf
rKX8w5XMyH8L8yPlFegtSw8k3NM8bLDBg+20Bvjox6hddl4xeNGK7TxZRaLKOxEN
hfoZpneMH3VmQ752+qw0KLJ0XIK5ZfmhsK2vbC/3M+jOTBTymGB9gS8HM3gk8LNd
VIyx+yP76b6OMPUwdvBOauK2/FrK5Rp5Sted0uatlMe4n1XmD/KjtSogAVdJKLKz
TKucDHKTOFUq7OCYZ1g1a5DyZ5otUKj1KjJn0Vptd9BmJcuoIOKVShgVdS8txi+P
R7MsjF9YeFBZBJtSGINaMnQktdHZeiCbOhwVZwyyZAahotIlx3KpItatRat8Xm31
2d0peQCH/RNBPY8BtTrwDOMNT1U7ifDBGz7AiYJRvcyBLRYzibYL3X35oB5bSxby
THh4RBFeDMUfJmFynpQovrKFDE0LxLlFQy7+gj7Bw5tYDy9P/xVDlA6jFm9C8Mk/
dKDjmyZPXTiiAnKNz/ug1M1hfwJOBe5CtwqI1oHy9teFMNr08E0HH4YKbUWwJrMq
PanXnhWLCQfTHhTfNEw+cPnfMACZ1Mt62oMWqahaQKRrtBm1Cu5lZ0VXvujGe6C0
IM8QP2nddZl5qpXJpngaRJI/mKwgnJWDnXMXSzsBWvC3dpUWrMNkaZEh/TzsXUHG
Yw9/E3GloC5CkrgcBUWopQ2DJKNyT+h5dEPJV3zU0Se1gfEHNCFSUFZRh2wWse8Y
2/uCWpG6SG9Xi01bWyM1lC0ZrVjtRJH+EIS1qIXtEyHlVNlIPUzNCpWfh02Wlw3h
20Gqe764jsIJYxlwHrvJRdEMe6zxvYqMyCEty+bgKONGbLA9iQt1apvV8Ke0EI79
FME52AOuav6TLcyVc39wvu+IFaaestBQLx0IjBqRcqdCl/dcexdq+Cl9wX0sk9qc
66qclJVdecuztitIdvUi4oJ40aBEUJVuF6kC7w3vZIrbT3dlXtRR1jYeSsOzzB0l
qUXrGMx2ty3U1D91dFheRkaZgFmSYZDhUutB1SYyJC+ME8kV9e3OpJiA5HUMGTfD
aGLe7/9Jc/aXRl6cisrDi8ChcWncU9K+XTZksh3WjXTo84FE5pF2oVyc5CM42dRk
34hbKV1WB10gN/y1Sx3Jo25/ISfTl8f8+5f2cavMIybWF4BB8pJdkR1Xh4Yn0w5n
uw3pBBbXURIrwkmbT8CQ8JTuYd6LbmBIicNyNgN3clA/vV77WYpkbX+QZY6tu6m8
ffqZDi832AmoEHYiaXVEtB3xV06OCzFaTUkydBe4yc1VMldY37a/wOYklAiocvQw
djZ/DKyoBs25XEccpPI3ixphrZEHy+rajkT07gKbZRL50K4HJOiq4TsUnu1VDDxZ
bvpCMEYlBjsbzdizZJGKGvRX2fs0+KLCFe9r34A5LVhdXDZosn5BCaquhyKJrwrO
Co8A7rcM26r9ulm1ig9NdaUzMKyhhulWRvEaSD9t2KA+5PF7M269oN9ag7nxwtJ4
ZS9CKIGeNV1l1oHw9fK9BV8qqZ6O77unJyb2fS9GiYv/clQnEBSoT+2l3we0zgDU
/JdEVC8JQkMEYtOqAhBlXXES6Sc8l1YrIZfHHUm2rIRWuFnxkI2HjGxKVf3enfzA
LZOvcxLcucrnQOW38EYkKifef9vStCd+uOGo/nHysgWdgxLcJgCYFveeVGJ5n5R2
bRC+6sgIGXqH9Pxu6VTHIK5Qvp72oyctXocfl2ZghfNs90hCVDsnYjt5/VUxKY9s
NWJGsFdjwOpkfghEDj8+keMuBm/3FXTH3MbSlzfbpPKDZAkKmWEb40M2Ka5tAVpX
cpsSq0TCM2UQR5g/oG5m+TVk57JunIYFHi6cHbTL0w3dLTdRk0936kpTvYUlv5eG
hWTb7IO4kPWhR2vfG6JShXehNR7QyzrNbWJxqOqOov+3q9cNVJALgr3rWLfWbOl7
KLVpsgBzS6tl7TeklbQW/H/eluqeXn28eiG722kBVjshDrVmq0dkD/AtUIHzFA5n
nNn7Qzc2cpja3exjzsbJtaqPIUFu+oMYd1skqobWHaqmsBFu3KZDi8gRYScA2CnQ
Evm4CjaSvnBrrWMma8kW5Ko9pZwnk3QDtrJzfTs0Pg/t+RAOD9hUgPqcv2AkGfCX
HmFGqjUw2cTpPYvQTD7AlVOT4VVnNBC1POXQ7ZwbEq33ajubbMk1WvgOvrhvkvw/
yHpQGPfPWSXC/HnoqC/gMUzzhQLBgGRivSF5m46Hr6F1oAMkBQcmS5SdVrg3CvMu
LAG6pg7UNWI8ZOCMJRn7YaCpUEge0HhPTOv80lG0tLYL4FhXsfXX67CdIwztZ1ED
jpIqSKiUaasd8j0XJ3GYbH9dSJ1Hblg2gTzrivv57214LSEcwPNDCU/n2FYHKzWD
Yxh+c3oWBgvyTct4V4bjFkDOzW4Ry9YhI3sjCpBtUFDnu3PJj11u9tEngm+wsfc5
MzJidY9WTGKff29LA/yW12JZko8Ul80+bgH27B11OgRz1SEIdVxOt2U4T4ToNfRU
ELO7lsNWbtbWB2SkZTgDjrZbZmgL/BdHUoqMbxnktCVtZzTpXJXBIhgz5TQcDdf9
5Yw3zXKYVcsA4h4DqKyDZBdDyhel1c6C8aV/k4bZNFzaGv7wRjf6wWTscEO8e67Y
Z07q+BnD9roBZu0iTGr1MHTCiZbUo90EdY9ZDw2oEGgpnUFnp6aLxwAOjijJ/CVX
ppL+oiAxc3NAWxpsW2vmmgkDNF4kSk4p0/6x7xrnbOmTe1dCxsrx1cI7npQM9lDR
Gf3oi4UlHGAs5zpc/MvSpwLnGPo3dZ1k06sG7VodzdtkVVi4Yjt4SITS9tMCLri3
X14e2Dpl/inBYzlKw0Zp91Rw41aI+7CRn4c8ph9CQWc1LL/hqOQGhp2qhtK5GG1u
hU3BA9T4m/ChKn/EHrzd0gRhLPyxtZpqSysE+3R3ObErkgUEWFQJgV35auqmsnJF
N3jCDTwRZls+W2a+XVlmEN8HfxF5FbTf79w3zf50etb84o68B/KGF/uP/DMCLB7E
k9A6ktg8Kz9hluMiIx3I/lTSCt0dSkvzSrIzDO0FEvfk8LCDQsRzF0F3mc8h4BYa
0ZcxqWcTdQqTWOg/l+SM0hOf7rCUfC9MHOPQJdX89S0uk66HZjHM3OTT62pu+f01
TLbuP/LEQmVUvuIGo6TOD24i4IwJR074MSb2/mYo/EeI5DGnfKbL8Me+d7GzO0dg
maPpO7UE2Z7IrqtkLDeVV6pIqY4B+1QyPRoMK9WHs8qbDJpiQ/qU4OGdTwMP0jM2
DRVTrGWIZS8xJqOulhkpvpqKW6iAGAgiUrMbnlvuDoT1nNxB8a57fa9I30dUZAOD
oBd/45RUeYAwNzrCd18mnpjDIigiPN6y1148yh9g/i84sWeQ+o36qbYZy1XV7tCV
5ab1Bu5HPrSeycKqCDEJ+ugohfDipqyN2ZlSLwwW5OZfobDbYbhZVFExL8unt47x
CzksN66YOSUbz8yMrggT8ptQuW2CDjUtEqtgSXxDThyO5tn2AA9B6R5mDDtCIRj1
xz4RL0nZpqEQUryw0pLURxH4ZsPYoTMOGNzE2yA9AIt8esaKYsBU9WSphMIT+sD/
Yz2C9Q6mDjdLjWpAF/E4LZ4/9stDyO8AtChvIGcQgKLlMGL1cZYEyxJ6sXK/B37G
6KjwcNKpLv9WFx/XqNd5YjMy8jrfw1u80vE7CHmXiW7/JESsB+YSS45Hu8WyS7CB
DTw+/NzHxRTeZ5WeDZiO77t2mn9YKREpeEL1Y26HS0jfU6CdaXUxIbsTHvsvEK+B
V1N7W30aBEbQSLbaKTNB8tXgUS0MCajvE+qKyscZVzTjTlanGzLA4CATP46qRofU
62wbpjIRQEDweFUW48GQus5bEJoGf+K4YYnkmLDoWbnumEK6gBuxf8VEfNJZd1HH
W+ArUTWnB81HQadP/7vhGBY3aznSV2RuUkjv6CVQxJNqGKTSjyk3wDITo+hrM7VK
vQfkZfthr0yLHme5GYU+5Dar55dNQ3PU9ib5hE4CmhtNeMGl2AvxE0VhHkiz2F0Z
4q8gBbPklfPiTeYfqDVuNuMClOh51lGS8mR/SENtuLjoEaZV/FivqyxK5f2snczd
L6eGCEs2HliFIRHazMTLxMQ3S6eVK1GtPqBhR7adxVpEtgUZyx9VspTIbQiB2bZF
R25kFsPgTYeoklUACNBSTevOkCXBaOXy6AuswyedsfeHESlWSE6K6oTDD1g0sRFW
64petuW7fIYQj8VNa6lmPBthdBZe5Bhmza/xWRe354uUb8I2UGZ+fK16UCLHDe8r
3XouK1scH480CTj9+Bj8huUiodRLiWhggsbGm9f4whhbghecDfGM+K0jYI7TxyOz
8OdyjrZCMECsHO1sTImg8MfM2v9uDuCvRwPNjXn5SnzuoR2mpp+DPnWDHNJyqQV+
bURvgV/ryMbVt/a3E8eaAdASQ+PyX01l4creUeBZr4TJ+a6lfZbHXfIKSPZ49qYr
9c2J4lecoT3GDg8aqEw3ByuUSQiMUtu3DdCqDWKRnbG1Rz6ND57ZWTqZmpzF0HzC
CBaQTbs5d5EqBogDIrGxD578tl/T4jGWr90i4FyXov+AXprZdLUcxrl9siwiNjiq
xV2azAL8SSX1HdPAtHdLiMgzBI+KIAnhuMLn/oNCrhAuybFQAG3EMO21UYsjZ4Ke
1SVNdsfqKiHLhPlNBqoqo1jyTb3a97ufqw99e6YtQEQ3wcnfMGnAuZGJXnajb34+
9csSPxh9fDiYqPyO0C2HWgdlgtYgnH4ziFoPw2cUX9y/7xbNXX4zWuWB8a3GR6ZB
wxgLocGCFb4k1XSOG9WoSs+gRVIItrU+n0iR4nEb32OVj28dO66FlmA8rJiP7//c
LuqjBKaZjEqFML+FHajx05TsdwZKtZC08OhGYAnrpay6QhInsfaPj37CYHI00olh
8yWLD0IeWoVUImQMsfJ128/2zR832oFc/5Zff7GYRf1a1ye5sJXG5QoULx41QNhb
/BEL9IGmKGhY9Bo7KVsgUDKl4mGHlBr+3jg4lr7EJgutKlk0/yEJyHVRKWHyq4R8
WQOd6C8XQNUb6MNClvDyVd6nFln0b1t9JrKwdOkbkSgQ9CF4LhFWGlAbk2p5deb+
KI2qn10C9sETCaOukTUfyxuFCmXnjfOf+4rnuxgK/buNR2bPpfOV6bV2OLbzYDQo
LwPwdYyMkCzckXNyv6zNoJkuhbE9l6Jns07novcWDZa2LkFvv6EDZ96eMpeDtH4G
yk4yz4Ix14WijO1tX+y+DYmvh2uhMzdJuaX0v6lTrLXEIOaUwiZjnL33t59TOPh2
fsbD64tqM3Zu4rCGcJqIhUEsR3LWP8WlEG4iQweypqGamirK6SPpEcm+gN+D630O
Y7uGWHHHQOGQEGR7POC7kcyQd7uUGBkXNeSqCwbR729CYibwTud3k2inzHBoLTap
jUUhYWJhiFYc0+s/RTsNWWyiPe+YhWzUO3reCoSJXWYPsWegj9iu7kibrN7/LgpP
s5taZPfjcKjc8PKTr7yX0fePsK2UGBZw56dOvVM0xA6JTKDLtSdFqW5lLBeb0ORx
YVOVIx/oyMbhds06bTY/70Ul5iwTTXUuydBF08bQVmD18U/Ma+xcfFrEHW09MIgo
gdOt6090BFTuvG0ZDUOE/KZE9WFl1SkHMJ/XZvoH4WH/BQWaipzh4GY4wT6GVniO
Mtvi86PaI5hosgBA2+KK/zetvhjZSQpbO4eVZDSsWqdBdC1R0JIPvyNKKNfIHijF
/D3f6LbEWuAY8QpPYyxyBfPcpJGjCvYzIGDM9lUAVmbxWCbea+Dxntu3gZNupsms
GlAX/IeyEWkcMOebZy52aBnZVpM/Y0Nuyev4Urex5LkRPjBV452T+dEEl1yILVFe
VxAauAknmhuKnEGsoemxAlKZgNLg+uGghuHwug75FLXmSUTV9cSpT8RL/UnUY/b4
4o3xixpJ3Hg7fxVRQ5mnCg2GnaIjhq7SLwZ9MNX/R9ixdY0QEAecxNFrZ1xjrJ0D
TGCjwrl7MXXPAjm+XpqQQBkP8hyQB4eGAN5uS+qw03dRrgvKyG66/TLrhYMhqZ6o
iedFWcj8mwRRCyVxDaV5NnzH46cJZ9HchqexEFpcEhX2ymLY3SJdjChZMbmE1khR
/BxC0jUpz4bjp3HjIPba9W+PhUaDJUZD6XphRjGOAllUPabcoOuA8MQ0GFd3iTmK
J3kqanceQuqknqcAiKZD24Xe76iSxxsKhvWmfTqn63+kuRbfDK46x09mlnXDNSMo
y/Z1ixpK44jVPl9jjUZTqoCjaEK0Bo/DoIQ5GmBsr59lCN6UiZQzKNMBwTnLaO87
34UZ6WuN7qUUW259XmLHS2UnX6PA2xT9th4PeTzVXC3/U/BmIL22bVDDy8sNvGsB
F7ivaZtR+WUlFuHKVNRc5H6DGxDN4MUZAsF/OdpNIfpzHEI2AqCKvtU9voo35Qpw
4tpYsW7U3lCfIcVVj/yhV8y6rVtQUHkD5UOT3zhotVBq3+1cHDemZlGfkk2+Swou
zHIM+PDwuWz5PhmXLdAFzOo8n7QF/fwidf2WgSGO/Z//8NRcrhC39mt3VSJVJoCB
kUNNY4ZQWHOMXH1COYduktJy4cMIP7pAj//pMc03G+3PleIzQyK5wLEYx9UGorrA
3hKc5t3hs9h1Ep1/1uZ3vbJhKUzSf4fEDFzWwuNdPGneP6q6gQGILZhebRb8zF7l
AL00MeACEGGM4xqkeoqyzjAycoIqD1EvPFAHfHHPDD26JUjAMjDIWoGXuRHDxXte
8sWnIcoeILtcopoTMO/nSBJV31HkftvsY5MALMpIHTvJXjoSMRJYd+PqpO10xhBe
NZ2Nk9KpDe9crlctvwSGvZsZ8yZWM8sdYL7xNDbShliOQT1HwE/uCwfbMGXlNP8B
k7NDOheGhpAFIaZBVFD9vqnrwiHr2P+7et0Q1eUAHGa5i0eVm4KKvXCoET3a7Kpc
dZWLK86A3vTPR3WB5pru0C1RossIWYX+eBe3ThOkqwt3Rxd6xr21St73OAxLbb+d
8dCfdU21uygI/6p/YKXJIosz9PiUgvIDMVt2r6f6PHO9A8uxRptyPP15VTinRb+i
X3pcLE+NX31QGrToczkc6ksyXpIqrvMd3KL6CbCUyCHG8OT6a14yfefK+8SHHeav
XLdzxsk1WNHZTCNtDkULNTNxFJPGNtjQUgq2PpI1EyzBMdfI+4IlLBpYdyEzP/un
eVnRJGJwwR9TDe59bhqB27aYRhLBXXOCuHnQBEA7nX4fsqwfSoR6R6KBPUdfRyHD
NME0+j9xQFrm/yUIivUySOyJgTWo3v88hDoNNbcq0sDCZrPqbdvDxkim4FWVI1lQ
hChZff9hUtandyYE8B8GFFmMexiHeEgfWEjCblsWMIeYMEFtGtf4l6FPu0d/cZa5
WwEAeMZ5qm7SAsXfBhDwgaud4QJnmgY4KFSRyP5L5iQ+27IkTMIlTd2ifdDm/IWJ
O2ncV+KLH+Q69xkoGQn2m99rMPJq52eKb42uQSeAtuOdZlkNM0iVqCDVhOEEU+gT
S2vU7eUM39T0fXHFjuPKt4xnzTJOCPG3GKzfudEjjOidF/ItbrsxI6r8/u5mjaCL
e5iEB3/N86Kbv3u/X+rNgF8NkJSSZE4GXarqcUIF3R2TcgyWR6FNYN07acRgoEwg
tpx6k6gXbb1vwPNQDw+Up/tJy6jH5J9Gf7AwY7xX2WVrHxuosSiDZX9WXAj0jVis
fNu3KK0FCQ9oHCnqVW7IdzVnoXp2bGo1QKLJuPcQKlRGqYPuwZWh3lYMInfGcC2Q
UQuMMCBi/XuO+cN5lXpgEmio3TWdS23Fu2tX06T2Bo0p08IveXzq9G/qDwhwrano
gZVczFBP/zvKCqLkEpkTpG5X8+AE9/Tr6MLqQB+xG3iV8uzl3gBEj9qIhOU7WZWR
4B9AbR3ZY9WvM4J2PlF+1+4E7kxASKKJiOit99sMoRP5hyrE1YF4ljMoDFlsip8t
QiwuXg/PIQldQ7DiXDaA/x5qj1k1WhkwSVgTh+pwK/niv8kU50ndCQZZWVCodJDI
W04z1bQaXgybXYQz7g9tTGn8vPFbk9SS7qCpteb0T1Wm0eEPq+WlGqsxht5deUwi
03Jh8p7xjY1AYmISpm7hQGasY1dJSt+HC708a0CIeqgGlCEeoCO8CZabD3L06liv
EicpqSGJT9JjTEV2/rJe/bNgu9SSOLcfOaqQI4BhP4ARu7+j1129nx+SPw+VyIQt
V/2yyYgVoPYlIWq78bFJyJmEpcv4dVTD6Dgp5rHPiD0NAuEXaBffLKHP+GpYRSxs
WO+1sj1JmhghVayeETSagfYjB+koUbg3tegiSgm/4Lcm/7zjaggMFAXADiMwJCYo
nROclEWraIlws5GJYJB1uLBfSU/+Ys6n3FpDG9E37gVyJTzA6u5FK+27dYli3zAt
d0zPROy0fT4ZdADRUd7oXE40byW/27/1m622nvceQAhJyz5mgsdeB+MiovZxn/XJ
9rQttWDcT0hFCrX9yUwqNSLB+ZFyLYhmsAY1rQBjzjq5M1mX3x4mugwiU2ILRxAp
UzKxYfDR8uhH0EtD/xLg8+k2KWMvjMakQA5Ui4OiWn00yvNJScSwVySFrW6UfqYT
jHuZU1Iv0/V5U9Lldt5FJfymku6AF/GpRbq+0NrPzZd+MPhCYzoy3qxScqO7TJTX
qOgj3wV0e1/OxDLxTROXd4NVv5KUl4/GshabWA5XC/rZFEybQIwHqKb7PFNd4pKA
HGnP9vGTQshx19CWVJSseDrJoTRPZo1e160QdjMPamLJYdfP7bRiicIAhKt8ZDsc
0fGQybY9y4UjE5/r/7JtC4e5D3UJoO8trY13sKfI3ax4/df2/aCzI49enQmunqdy
FxVTrCHHPkmDGCKBr4pgHJV3KF0SlV0s24VKdUHvQ15cupc/8u/NaZKJoJBd7wOS
Z/FICjDQcwNWtEFqVp1IijcwGxxNm7XlrhGfmHKH/vfL2erdZ7k7tAqEksUVtgys
kLFy63s/x+jS5QDuhB0HAm86GZ9l7IfUJ4gUyq2V/T50HYDTklDHbBWfzApp9Lrv
5exgRGPdX4SEkm+g5CvuKQ3x8oeJOVgMIUdiou03zRHDo7dp0ErFC6ndk6zQz5L9
+5NpeBdeWwOgTbyv83efEHYspU7JcKIZBVS2yYnJLxAJvkEq+Sa9vPx4yu4vkeVb
otUDpmS2a/cammLC5kMkKr79sxT65bAUUffh/ZLlVTOBniEAGpNk5vGTnD6zdjyJ
8DnOdSlHeHZkibM6YBnLxBaB2DhfWhf/J2zNpRkZ4CWsFITiqs1uxn8UgX4Q+HPN
tjjUkdbjx3U24lnA9/JWPy9SUPbfACokKA6Lg1kYqp1gyNuWbjpzmSCZ6chknEix
1MCXDpKAeMIN6x14yZrDD9q/wQ3SHs/k1th38Zbv4w0Qu936RUUxwAa1U+R+hzSd
oVVqrmzXM6jBf2s2AZlGwqts5gzgVXWsU3HS21nZKzVP5tiadqID3piBMd7SZfAu
NgbNA0DUqaBgC+YsH4ZZyt/gXGtHOqimchGd9v7gEEhnhWK2pp+TbaWn9P6RHAx2
RxrzcCPKAsqcSR42CtkEK7Pb4JmAny9Qnlsr/psSmgy9caoF8zWD5pIGa0v/BlOI
SLvHuo0bhsOvr1FWFxO/lIV/7BKYbE01SYKW5A3CBTEY0s+ys+FWclLRlpq4piQB
Ppx3Qsk201q9iSl+54tRm8k7K3crI8dps0wAhAcJr9glemPpLgveoSJaonah+uhT
40cC22o3A9g9cQy/4q4/oJeCr0TBpTOMRJzRNz3LwtWr/doFDM2vaxq5Ye/0Drw2
olIiGikLgxxY3w74mhpVN0QRI1YbdZjtFuPMPmhpGQ6bEd/tcz9uUuhBl8kTeMRF
tw35bhI1XpHOMKnhmgkpqyf8L1fOzVRpjEZP15CuNhOmzb+yH4Wxz0JIhMdABWq5
nhnt30K0MegfmhdTQ5vbLXf8jki39xUNg1YNihbaJz9SU5Pty24ls5LFQ3QPbRJv
3iD0DH7Iy8dPqcvkaWvst2MjY+7AGHdpweYDuuM5ca/lbczLFIetJRq16I8JmukZ
bdppbicI5Tf1o6eYkqrxfnz+hIAjjd6teNIu04g1fN5lLPsh/p4c2H/S0811IogE
7WOQytcNWV2DHkl11QumU69mjGYRtsV6tGbqYGOu6GPbAcx59a4VGILSsq5VeJ83
8JlCfPZ1ZXujLz1QAw/7ueeX2TOLTVOXTNLAvhUyjReyZptaMKjzva9ItNhAjO+9
F/M5yR0VQvSISBaiVaKK4YrjUbHulbGXR2gPxpyD5NW224UnPx3KvAwbtyFK9J+f
WMQSXUz1Hto2VvJD6urG75dV/V05zJ7dg8BX2v1eECaGHi7B481WQx8O9rrFrFxd
TYGM4uoEQiPf4L+B5tX+BxQuw7SD0MB04mxi4xe1LBV+CGBan1NrZZerl2BE+ThU
vfZVRTeROenKiUlDjm1XpTQ3kk0mdsAabiqE14MZWhNLXfhM7yzfthXz8Yv2onoQ
ckdbMCdjjaN6g2RW8mgNCaSZmS9ZwpMWZ9tUun92qSZs7yOnBai9cAqcFF3TmA6z
Cp9alW1tPzVLHbWzsM01KKz1wariuG4EAg+GxDg0kuHtkN1JXr3ODGGuUB87rDIx
cu1TNa7DQhcq8ZetfWGple6/0/wI6uMwqZVrF+b0yzCLVtOa+nEsFou0KDOQ1Uve
2Y9VQJ2VYpUJ5/Ein1cBEkRzKdyCzUADBxK0YSrayWRF1QMZghzHBSYxvwteUmaV
n/8j086A1KPtY0ASvFh0HFX6TVLkdQQ8GhyZrmlRUdNBYHv3iYkTOuxMg0tge00D
HwZklsZ5cgQWys6yjGH3ptrHDKNMlbcAhrtZk3+LZ2k6Te8qF+lAVhCDzAYQ9nPg
VEtX5juux11aC5jiw+axG2GG9PLusawX7nZ8zM9FPNiGmaXG98JHnIdpfBwCfIxU
z4wOAOoC0t4hWlHjsh4uQsRm3V+2bBcXW7N53c5sm1c7mxnQnj1yRuvitlvMA8Ab
ti0W7s6XSbvDSJP7OBoXLY4AX+lXQjzZMsaq9wFROcgmYo6w//ZUzoRXbPmwmX91
oJb+ZjxHmhx2XPJ57dlmBoybQEjNLy5kuIyWpL44xOZJr1ZwE0nR+inN03X8WD3Z
HOOdpVW1yUCAVzKmmcDoVptlP06alv57KU9FHCuuswpMvBjLDoL/zXqFD/9XjEeJ
4EM7WLrq6GfP5m+4GTcbD9VfNMZ1Wh8rzldHsmtOP8jjt0Bb7nDJc1+sGv9Nr6wd
f8RCZvIZW2eLh/n9TSOjWeVchQrEcaP9cj4IyTrtAU3yN0f9bc6Ig4EwyI5pHcFE
ukjYjXA9Skpi6m0QQXNHS+6E5TxuHlN4iBoteNR1jDyXXXYQ93WZV3ZFIZYuaJaS
jZ047KuyGFDuDpUJI5WJ92mWoQvn7oOZ6szt6yh8X3y9sgTB+m+qVDZ4jtqAxmlS
OJEeWdmK+nqqJN3eVcbqetnTjlvr7SLhDVPVVsPInpoZK7h33FvqgQXidKcQRexx
nWmM4qcFfppSVU+NenUNOk4qk3IOgQT3cPPqOQIeZYmxeiW3WyFuXMTSrdVk40Fl
yDFyPhIZsiRC5E5LVmkFroIEIN23HHKoXSuSZ/k9qyeOmMtKOncUV9+bFBRBsmFE
YA0DUDa/0foM6NXMIyV2HhZ682HgCapt1o75trfJfCmNXPDYUFkAYSwdYrpCj2kD
UGTP1A+vAL0XjMjBrJqshgFnCSxB6nZXulcD2IpRVT9a/S/zJwKWqolpXe1dZNOv
SADdR87zSFHp549E9T1nRi4WXrUJMCvzjPzRz0HEGai3F5wpEWGI5dB34PELWWIo
glwBoI7o5cSmi8b1IzIvqsp2oaPXBS9Nh8i2cHI5Oz6CBfVLOhZzTPu+E7VGLraG
+8l5PG6kiZAuiyocc3f1Rj6jeLreuWEk91LxX7uhdjGoPzyD0Yy7lVijRgr4t+pe
v7ukj3tpn/laLqXsJUWDCfo6/RGxhHqjHwJedSQ5VOXDhANP6xqN+vVW16pjrzg1
h/hrHdf7guyWJYbkAoz/r91t0h0IMs71uHl31bMJZPySe0cXVmPrhsDrqYIOABB4
gKzF5N1yXetlm4XzcWH3iIq/r/GFhTROtJVE+AnkwZTRxbcUyjr2i22BQvrRKKU/
jcP4If5tp1NkTvD+mNJD9kM7drARSHIZR0x15RRa1niCFZnsqzAWPlR7bxZD9Dv1
nhJW4Oh4/LxYotGhtoDwB2Ms/m234RCcIo7J+6fgDm8NYDzJ3cy8161sQpBcXYu8
WyVY1vppUsi8vKgaRpSJ4jgt1cEHcRDxdgUDtVqRJvAy0KVvDb2/dDKteNTAnf9l
L0zJBQKA/aY8drCUCoMAVnAlbASm4N2FQsLXx3WGOlIUjS+tKn3RMKflEV4KB5Ip
Gdk7Zbn0WQE1bp+KUTxEGxkdJzDVLA5ZaVUMbcCgjnLBDp0mdA8IK2vg9yUasXjj
93wdzlyLiMoxEiQRZAPvR8TELfLxn4NBko0JCFuNcU5c3P/F1S2IyFrp9AOf9Kmn
ieWuIoy6QVEI/e1KrfCuCLVN9qed1T4jz8nDz6gsiHVuA3kq0ZPRZXeAzKAAj93z
DDYodal06N821dNlXLiGoOcY6LkMsURANUEJMRgvEz2jMARGNMeco7jtIhNEBPBa
wyTCFHmTXo1kwdt1gTPj4X1aYH8w6L8J8zdA8oHhITRMiSFf/ATpkvPPZIFAO3Aa
jLQ0q70D+prRA5Q0gioDdGdN7Iuyoe099qk+JjYG4aZETtLrdO1dol9G2Ztk01Za
gvc6ssAC6oG8yfs0VAVr97J5Ff+g9LOZwnzeCel+jEFgT1uiaqcjRA6LqwgvvGHJ
FY2ldHy0uKmRDlP+GycJCcuumSfiLf8fw7j8G3oalMZQT5KcpTpcM7nHB5BmvJXs
ddqDgpvGZ034IxY2ftTJRHWKcvbwmZ16MW+Cf1QLJZJgk1nX/g+C4lLh7Bg3wG32
uzcOhxjKyCPShQQ0DUhBU8atlnWrhDwtUY5622zYHCKFW5Bo+tMmPt7njnmjGqkg
Nw+i27fN2X6ZAbpelAqPNzrdq91m513cvonfra/5hOWmaV5n9wwnenAyyp2CGjad
xQ+MMxX6jV8bmHXqvbfPYOFGHotIEsbUTpi1eJHSH/9axMmQM3hhQjhUmxKwTi9o
kGL28RrEYFMxMMrogpd+RwX2lGveVuNaIl5vbDsExnYWYo06wwr1YBJXfGcukrNp
AVjA5aD1qrNGs1u9V/LasJoURHlPX8PJocXTrWfjcbLx3r+eoKPBp0IGEYGzdA6s
Iq6roFddgATcsHpEwClyATRhBGEZFg2GZePQS+Ug+rOAuuhg2oWHL06wtOpTdHWn
jZ9T23IRMC5sq/c6TOFxZCbfiARZ5oecFZzhvFcKYXM19/Z3uNwXNB0wjcCrfnhO
DLzZoIc6wmF8zMwqqHf/UxLw/Oku2iBcPVHP79GgUy/yFnqu/0BbO8FaZAAJk4aY
/Vmzepw3wQ9fDx9hwpgLxwCm+i+aweSJp+YItx/0PybWsAOkr4PwZqpxcMTdgnx/
Nx65UucayrsJTlAfx4d4crMWP88Lue6NInu8bWxQ5pIzo1hX3PaTS7uprLS04jfD
QuSD0fwrzhgfu2nFIWkS/7cAM9Tq5dbAXJdqUBn2T1I+WEUvBCAQ5Q6MdIF8LyoW
ZVJV+c+mXjSn3t5jp0Oa1kzPJLExhc6VdOYkkt30rQEy+7cqBqLtYoS7BIhAxBVH
e4uGJ3zkGRj045f7zOVYNk5ATN0mtGeaumeV0PDxSGukIZpX2EABzAm1+BWDDcOe
Hsai8dJFKdDjA9Bg8XAqDvc6GNJimd5CtSIrz+VbcBGe1Q12r7itULMLYDncLeMx
8qpJ7hvivSlUXc4WDKEGHHoxJ+M6IncNZHw7hwA6gA2LIW0jHo6xOcy6Z+ygj83j
d8FYtF5tRU98oqWTg5YmupHm+d8IS/0BQnWUxJMnYJ+Kodf4fHdiUjENel81YQ8O
vyJJZ8AwYjIkZ5A/uYP9MZ+7lnxdYte7bYHzPqykVidJwzvWdjjbfMziMl/dp2SS
Jpb3FOfEyGNPO2fTxY7VwW5NsjTqborD9y7Jb/QqV/bRxVkGKM0SFfvTtenL2nUC
krPynkr+x5I6GgSFxPtGq48AWzR7IfkxJd/WcJb6uvFU22j8KYgjfERAYw9X3ozT
98ZcXW8uAFiXLnXj1GJqdA5upzFtV5Krz0Zg6BISw+eBcuA5Nw1apy9+a3Efwm7l
k18UaDSrz29UUU9TvyNpabEzJXjMeCgX2fipPfvU+ky3x0s2h+0Pkz4K6WC6c9Rl
4in70a5i8ixXK8k73xf1MrJkP+xaDWyQXKZN8vjRc85+t/HXO3U7oBPWCrb3wg0D
2vVSAibJX3Uc9AgVYX+XZmm1UasECyr+CBvysteUrQEIES/E9cGq5wzMYUa+g+4q
BRYOBH4nFQcQ+nZ/mqNnacEsrJZLhyK8rTJ4a8D9Vbmmts5YnnUbKLYstgobaO5Q
Jxn4Y2vXYBc+sk2GZOyDdy0atBEwfXrB9OOFeXyb8I8kigTRScw8PWu/dUa9lcIp
O081tJv1Ma9eMk2cNETRjRxuKNO/yJ0yKqMEXDK671CaSF5CKXADZWz4IZrVb+dc
K3GCuZ7nl191tAA6PRZkNglWBd5I0IXpWRmVb7CEHi09CQhrrhrjcw6IWq5qvpCy
uPtHx9uVb3T8Ly0UGpu/WMj4wWR7Yq6O2H0d6KQx4Pr1Om7WVJV8tQs2m7qmCB8I
Z9tEH2UCWrzYevuh4/wxrSg0ZCzfMFVUQ5gfL91VpCog3RzfyfFTi3bJVeh0sSAf
yhgMrjvP0SuWXu8b6KB3t3vM6rqAoFZYfKrs28yAyJs6x6sNAoNoA3x7mJm9GiLl
gZ7p/8Xg/xMGA2QwsxhLYzUVEPYFmB9TyuSXuzEOO3SG6MESYgj3SUQfp3iiNHE2
TASiRLdZbpQk4UVkK2ger6Ij5Bi88p5zka+/0lzN8j08KGRP2GJAkd8imw0DFj1b
psf+XIO7rKjzSNp4S/ar83ukSto+T+Hi/4OpzLnjbTEA48kwqOts0r/dbQzJ4col
t1AZsXNE45nn/fUdZjU4eNhHmHWGg87zrvHi9x0ef8yZnS9t2LOJfxQ+ZxN8hNI5
mF5Y3gjDykOhmRVUSQ1ebEvkB2vOSeF08mZBMhRp9YkHR1OsOYCL1ngM0VD7wsbO
P0AAvsJkoXwDeDL0nfVr1qPzrDMOFAp9XT/8/fLP304wX2J07rnE6GzfrPDajNO4
gu5kzUFHWJUtMiIUGnGOXXy76zyA9W/hZRHvCCEqG9RiT3vt2vxJ5wQquJTvxpB6
JAEP9uN6VAU1GGHX3RTcd8hSVQdwp9mLCOwuuooUxXM3j0n8vho6m13d+DN1wDUA
sP114N1xoxzixsGI82Q1GHXjyQ9xztCrKZiTZUJaInaCAf2ln54Sa6flIAwUyxEI
ho8+DjJrcHYa8PyXbvPMfXI/oP/QM3r2/FB9Jf4QmCbOdw/rT1qXfpxsAEWcxPX1
AvuKdX33KYQBcNoDh+AYSvqd+StzTUkC3vgiZ2tEmvkwKW8i4659PO0oNRc7ause
sFJZtlXJGW8R63dUbaOYjtOf83XfCxeKGvuI29yDEsKLDGNCt1daMKaOP7eTY9D/
v4wYbz5L4m+hHStgOMQK0YENHA/tdXyizKJXyLGmnnaAAGEFwR93IyP0vuphRU+s
fRiqUvBgHt0IPZhHs+19N4FJlvJ1aqsdu7gzeAcJz8W/ytm18i5JOjednRr39IhC
GFdfEJikWpVJhUmpBuXy3dmaEjTb5WbUMvKF8GA1C6vXdhIFHwxq7VcQMhtarJ25
GObWdBe3ePNNrFexkQghrwEHC8Xuk8WuHAybGyBHZI5ZkGv/IowpqKAlcMC19QiQ
P0l8ZS2G7ZDDSulaz0mS3RiW3uQv/4LQrP7/HgLnse+/QXxYGfrz9Z4BUJ+7Vg42
2UG9EtMrQtjyRvYvtdKL8NJg5gY5VDd1ucxcNWGhJ5kYcHaK3ydNg0eoBffBF7sE
dYta742N/C5I1BltwZPz+mbyqTfLwEgXoVEMKiigCpSNM/gtwt3BXheU0LQD6U0M
Tr5Xmo320NZAE7SIDe8SxqiVwZOjkHxQpK5LuYpPJU7w1Tm+Yq1GDBIBTjWBJqWv
NYJIUddv/bOm3QeYxhHwdHLR4sKIKk6Fgw8Sadt8F/qRPD/KIfEphiG+GbAbdHYp
7i5nczZ3wVs/vwWCSzNoL+DlqhbZIlc6E9u+W6m/erFmFvAfwShHXbsMhUa5+swf
tQ/jh6Iuz9gLMuMMR3Ahlj2LCZ+Kl1DocHOK83taSCMPzJzPUK9DiOkqGoN9k8cO
vNHLEN7XS8M/qKelvazhjQpzioaXIPC43ro4mFoR6tTSaU68eHam7d/gAvAjKR6t
8/sB+qOQ0r5a+Wgz3SqLqmDyhx5rZ+aEjhMXbxURn90esLVkQHDox9HGjpYTmBXI
/tJsnaF1QNjT2j9wnljVG+u/38dvnrvykXzTd6R76DH92Ulb1xkLFrZzLYouJgFd
yCmOXrBYhMS5kSovAljGogFOzunUfJ1f4u+xMsN1QFtil0/ZKd+7bEkFEg4DXa8J
YuyWzwrVNiEjgzJmj+V0W/udrAuvPFX/lOShj6kutUNP1fl1FOh5odkGdevWXKxq
ccrq2JEMcCUmB3+jtMXGDQ26OHfOX0HQqbj8enSKmuZsYnBPg8spZnQhFYNsbOH2
ZCpwb1eK5K1hp/P9cu2XUjvGfXM+sVUSs5tQWydY/ukg+ClDucQf73Jkhls360/G
eJcqBa08vUFwjGoBOPY7c/QOCjDbTWmxdCkVfBesuAIzPyp/ArMfeuy4JUsPzFwG
pny2ZimR7nUPJs1RrwNT23oXyqzHcf5/rqYlVMnBRFsYpadv0nyxJxfnFxUoKB9t
0WLvChWSvMyejCO/ncZKpW92NJnkmV2n/qL9gg5KY2Ro4UT7mOIcxOezcklOXwpq
16emC9KDA+ZyXbn6k7uDjpQLGZvjwKdPYqUInUyqWVZHfkGZw0SYZoXLawInQB2J
7VM3CY1u41QzupFh/b0cZFlvZGwtQCy8oC1sBQmRVrdC7IVVaw1QJMdkCObOeUFO
sOWXGlPYSGPsQ7gaOxZxDIS65JtH6PeCYAm9LX7Z4pnLSSA67KTk2fkfkvfmKQ6r
5k16po4zkyOsoVanVZOpOSDLxqp8K+8LvMrOo99conejqoEpo9+ARLNxyPw94aZz
9sbxd4wzXOR7FFSeF8EyTjL8uROEAFYtUkde5Z3QgSXyyrBOBnypf2rDiya99asd
NHsRYLZi0nm7z8u91g1cxZRefr82fjNQjzjpgABpjnfcZsfe5qNTqz0onmrpgc1V
1pDE32EELJuPyLk/sWsdWtR1z26gdEmcTAnkrDZn7vKmFmR+Bylvze1LbZSIbP9e
jIGczFFdt8nXruJNi5d4HSO9f8iKlVwlLa6eCYGH9PbdVJGUwTwlwWEy7gpJRvRy
GWoLj0077OjoTHhNWPu9QS1MomO/NPCA30vl+bOlUf3QDz+3Q9lMTPqEfZJQlHf/
suvnkM24f6HI55UQ4hxxFTsWV9n6PcRH+CjRCySCEf487m9zivHRo0RWWI80ryJn
6WycHw9at1MqVkWSOFLGV5U526k4Re85cx1wfAiYwM2SUw81vF0dGdlI+Vj3X9VB
x/lJ4dhFwWOmPaUChpicPcT8bus2Fdz0kT5Q+Hem/yTaj/sBUCM5nxvOePNgaeOA
5V1OpHjxbS7nrXw0gezTf/1kMuus7Q8NLOxz+gj54gx+0zOhyvgm02esN9vcdvP3
8+YOmLOs276P/SfXuaYgcBtG56KI3DhGT++UVAcjNroHj88C6Slfow1hbvtgY3T8
6qZluq1ki+0cVontV9DsSRlj6g/f7lIzqTLatAXoe37GB5WU3RWBt6SEgf3Ubs/U
kG7KtGoDjh3YAPWNESLbs7Mnshy+m/Mb+wBLofoGMDQ8Q/eRdGdFA6HeF3fx70F2
TbKx5RyRDKm5lxgBmlnVlu6BBjCpJqTSM0ldmqueQzk9Y7FP5O42idk3fMMgvXic
EOmca0QbGfsXMVQrh37hAWwnVfqP4L6rFZ7CbN2FDoxYYwjOWKci/fR7RJ8axZHu
6Yjdn3WEB/xH9bTYku+PUUBr8sNKjVS0kcYanhvuCtnviiKyLfh/yRLM1PRlInzW
JxbRdjPgMcjARnK0NlgwAVtIBJI1HjsJZ+3Pc1tEpxnoQUz//sQJjvpE4AhUarEm
fjlUjTvyO635+hfBD2L8+AmQCCX/pGdU3fYokC6iICJAsSz6gVNcdnlPJmpvhQoA
Jp1Hfuz6fTa9zmUoSHcZucMtl3crmVdcVUWZHuMOpo6YA/bZaQ3VXnKvZhJ3gFd5
bP5/PeoDNh8+V4SCa8lPowkLuiR8Zdd4oFo5hxK8sjfWzCn3yUaQ2s9xwvAU4iwO
NWkS/7NNqJkGjUuFfgTzSn6xANuNvxP/gz5E5vfPjqsl8w1ppoAaCi6VwBIjBZLA
AoiGx5kBUA5sj7sAc5WqiEZznD60YJd7PG2xS1zZsRcZlEETS4LtnWeTG+EDj76d
RCMrKigQf0/k2NmuC0fjDo26hNwj7iaWkqoxJsvc6anxr5lLJYhHFIyYf+JssgDF
nZcZZL6W1XhqG6ri+FyvcEQUT1VIjP+DCAdrok8x98p7CVbt6tao2q9TgSbQhtjQ
45u8vWxQk5h0VINpcn5pmAL7Xrt07DviY3Sa8NxN+Z/voO9FdgOciPkyuZGvhnFv
NJveD2I7+w8wIgShh6w+cl7/Nh4N9NBUV423S0+ae84Tuy4XJYx18JdiXzpnglYr
SdEhnUctVLJvj9oqe74mRuZP8p/pzoglnWFnZU12DmXuKBJwvUoVRbnJvfvGMJiG
7/4ctUiaiSW/XTB7H5FX1SXJ0kiZvFWFFQ6PlNvdfuBMmTBgloIbaFrjsEaoG4co
EneRuOZVOGu4gPcollIkyo+CuY+kN59EcIbZHQJdcGJxwRxo0lxPDcDrhKkO0CPY
TkaFW3P6hRO4VNAiUr01z9w8XVR8S3BpCMn/zGyIyibcy9WODOQVUeuTGpXOuxLR
2fcEPTHdDiiOlf7k3NwREHx6RoTM6/09+Q5dVQS1L7j969Oi8rTZsqba+DrNQoOt
SPHovL5mJS8kpSJ7lu+ou+CHCNgo6QvkjyHj73hRqpgpHS35hBIJfJTEnQ9swTZB
pKPmyC8fn+fc1rxFWbMPYeBvNPxCrlcZOwIMa3lHDP/V90ek4tBvQ3l3f//U+Ubo
wyt16yLxb0HiJ8OkJzoEvpu0IVoS/7XnINCoqljXLv37DZAdI8kSXZWbexHpl0qo
8cH3k7YdiO5Exjyk8ZhcCJFf+h+cF8Hd47G+lvZIOqSLImGOat/yaVvozJ3VK0w2
qjKue+HcjFhZrV5V6Ez/iyHHpMGEOWZ/j7YpHsVP5wC46VJtHelwnw3xXf3WfbVs
S5fnKiehJsVI9AXRR7WM8LurJyKbgFpi+wtMUvXQ438+4xsnK6uAUs3pe5P+3gaW
ymYG9xxQIQWOsNuTmKeL4jOWBP73LzoW1aB5Bkkzc83p+x2pQ4F8HKJxZ2AxoczI
lFhUJgPySLqmTxbuwVVvupCDQet1GKg9bb+uGSqeVSrJxPxTTxusP93NE2iokF3L
ntKS5pp+unzAB4XCw6IX7lEePU1Np2cpNYRlVIA4sOOeToDYCq10dz8PUaPRLRIQ
bRY3HwsVw4Ayos+0jZ+IeCCR+xxl3ywTQd2LvXLC+TiL5TJqWRMs79818CuklokP
kzdjiWTesgX3h8lRvmfXlpG86tOPsKOpTE7uE3xhvcGtgslaPdoEdgOCaw66RMSh
7Pk4wOYX8AyOj6mrtRvHy061a2hUnWLkY3SpmbrTkx60wJt0Yw7pdGL6dwlON/oX
qjWdKUkT8fJIEQjje4aCejsEOVI7QWQ+dVB/noDkkLWh+jR5hKesTyodGmCla3ux
okYhmwG37DQNxwQbWMiX493QT7u1ALOO/rFpG/xIAosyF1ml90SgDx70FO6mbH9m
Zt44HaUiVH12OXAvQFDIqzHlyMnvdsbwbhlR3bTRdC54jm5/JecT5dg/mO1/cJVp
Sm6rfVJasswcY1+9eW+S1NO3m8lJNztA5/FW4MLYtgb/Ekxi6GdocsYjLmefCc2y
qbLtyV5+5quDbYhI3WVYHX9T+JC9ehbk/rTtykEkuphnxoTw5ZhFG7R+s5KPPZd0
p9MXt8hqPBcq5UGXOFiDXju3cZ4oOBIfl9Rdz93Ka2JWMhHmLpjFFWXkKqLXxvdy
ocV66dkZS4WRZb0nVHUSXnEmPoqOsqlJOyFVuuzgw4T6156Nmjb1p4ozsSO0vSN2
tlXF3SwDo+a/lYsz2FrpatG/Pt4JdmeL4/K2CEWhAH7M/v2DwrmZFrhnLHhZGkF5
6d60+kueS6c3/NxU04bzbnrrXX6PPlfIv0V3dOup24V2G7g8zyvDiztfmp3t+KWG
2bHvG6XLlLlNumorbLP/GeaC/Ch7G7EuYSgRNvPxGnffMtuZ099hq8zKbQjqoN9n
1K67B3A4PPzXw2AOzTB5TASx5BUZFklBmORlw3ctoqlluDMNnL/k2ltDAhuZF+UD
g0tZkhsu9YslO9wqJ9pp3DRWq4CIjHl2/RtwTQ+F9wdnFjwAgwIoypccswZIQWb3
fprOsk+Jv/w2brDc2lzf8Pw6oenjGSNvba6UO7G9WVFTuQTZFV1w90CF6d2ARn4n
Klp9pt8p+nDeKDt/Ng12TM6jl411jlW/5D1OE7ncLjSJvg94m3JbS/+ZbZHun3qL
mUrgbhDWgc8UELpgZ1K3M7FYjzzUqeHmLXkQX5yuvfSlAL/5R5QqnnT5w003RXFH
N4N7r/as4d8INqhlGD4i9rV6AvyltrivEwSJhNIA3TE46yp9kexv9XTIQ+NFcEMr
0KMBo5Mjkcpt/xhk12a3kj0J7msPhY3fFMSLnVP7tmD0cmE8imF4C8GzEbgUTlZ1
B9vSaGKFm/Fprk5xUbAxnCnYt080ly7BJf7D9uQOvGeGKlxVDhUoOlqvKQo2Gk/s
wd99zfBiUOfqR+jJIL2uUwH10W7pLcZgX3cgUoS95xbaOU2yL1ZsV/qFB5Dtjzsa
IMWQN42cStXDr86osXp8cmfBhIDr5myCUa0m+eNJs3ylWEPY3zbM/UjjfukT0chk
3G2GnPM71Kx+tsW4q7pOalezybGScYdie1JrsvpEZ8Tqgr22oP2nujBTefZoUgma
xkKtGwKH/WXyFLduI39xxjWrbg6xDbM1uqYAprhMwBjooQy4LF4eSBBGc0nFIKmH
KpSs+3NVdzzmzT+DBRX3WbEYjc+lxbZluMJP1w7ytom/nDeaxh0A74oftYkUVwMk
egGM5zKFueO+IJ6JmP52rrdCoS19PGSxCI1r3mbJGf1XGCkIQK7tzOpXe47bVeNB
yLejlOrXW+F908rKq6BOqcM4LBNor98Qf0Ls3Lbz0a5Z/IXR5/2G5/ZmTJ6ppGKQ
z4euQwwsMlPMkBilS/GwVk2hQwp2IgqlRDPLHEl19n0RnD/7GpomaWnShfLK35fX
jwwCQE0HuZ6WEsQwMZCMMO9bPzFKAcNpY5UCA6YuY6naKy9quK1bg+zfvqovA5Ol
m4KOdpw3SCQdteuo/9jBZGooQfNNB1obs4vtF0XvliYipe/fham41+gii76ytY2B
/O+ZjGsudLCRdseDqhOjHEbRSojpSi+ijP7d5cJQhCvcyVVUTjsHFAf5qbn8dE61
hRnsQdBlML4fALW3ELMw+C9VNbbXxAKE1+7jVE+H60JhxPWdx5oVtYEg6S8Zx2uo
SKpQYV/A8D4+t/38N5r8ucphVaCyf5dqfzhmV5fSm/ibrvSz3I/UVrso66pyMnTb
4fX/8FTn83xl1AIpgUPXfSHLu520RUikDmcivJ7jbxAqJ8M1/wHt5idq1RXTjfmP
nQQB5hqLp4VN0k60F9UPKVh5n7Oii8WjnPcWa/dmQQUtZ+KhEvQmBUh0B/ORGypV
ud4C5mnoEmNeOMmNx12Lhc+5gFE9VlTg07qXbewgen6HSJypJBHziEU3cbD3vpnb
jRUBTDxuo2V0wXLfxGvzu2JLmeREbd9KWZ5V5sArpfH0l3boPINY9bBnzhMMwOwK
0KJ6E7avTH5l0nkTIvU80+Pb1JQ/VJv2oQQS7vEZPg/ptXaiakBm4TDUA4SXJvYK
q5Ry2hroIxgPbA3GW20jO4TPLskdvSyZA9HJGPQ50ghq+uvqKrNGRCXNZvgybyVK
tEBoWwL1ExxO5gfJnTkuLMKC6Zkm+Z58fqU34dx18AuAW0kUDbHvzMHYcTaKSMeT
dreujKXdiFSz4+unN0A+y7GjbcyhLukoLlrZzzaAh2bbQ/xkFBP19h3IdyNXsw2X
10KXz52noZGT4tZPz1a2APBcFK1rajWNiWy4PEVpVAG7ZLTQzIMnzgUWh/HJX0a5
Ole6t07QC2udYGWpC9QusYmEQYJQnUqC7Fnm7iZHVebfnMPNFcKvzRFGv4iOi97p
P6KmIO9AN6nMoAEm6cnSEjrLOz9ihW4YgC8w/qoxXAtZSuVJVm6z/RybByHknA8D
Kq4uwW1/e74oi5KOD77zCf6m3swwaGtCw8cNxZbMBUBNyZX+qX48aFKkE76d8p4w
TCRFVskMKU95fO2zzuId0n37Kc9Satm6h/qkwgv+/uNeA/ZXfQ/biWXGl7P4PJOU
rMl76MFiB080pqkBrqEN29trrB3L/srmavyITJE1tl7QhAuXQTWDVmUEO15i5VV/
xWgOSFZyvo3eDtB7DThOGkbK4cZMgGnaY2ZOZWlYQfspAPcYhWk71R/kvFhoC8Qo
bmxBxQX0pI5KkRZdOdjhlJ5J9tgULRxGnS5VEbM3Bxd52pgXMNzTvFdxZYvoBDo0
G6RBlwtmnDOlouZA51j0vA6zzTQD5kL5Uz2mAugl/cE/yMCZZzsxj9igA/13SQSC
6JzssAWiS/UnYQcFKmwK6uhL/H6wVjFyXawqg0T7bNlA2szqJRuekrlyRv+bFk/Y
uCESJGD7HY5jZYFC6VfZEQOrCOCtKn++Gdz4pN7Xqyf3VPL51yNWfaePz7qddSGf
3lxwHm56WHrcmORAtrlJDGiZ0JRcdRVCbiFX/CHTZ164wt9SM4vQ58PwrITzxlai
RzNVp+2uK9ht4guPquYhROfQDMjzVucvAgmPWK7s/99LE4h6eOAPC+wlHvq94RPT
CUSSllaR3aSQlPxdODNARV0xviNXMAIpPe0JpTl9pbHuykfHiuqTM9kdHnrFeudc
OEsuU3qYhNiFYIT2RtnwX1B8kav3XgZTE/NAKrOpAbp0ncbnR3fFy3MOVGPtbdlD
SH9e8MHwZYvHoTLv3ZE7hIKg/2PPnbOxyzzjscAzEyCK3PfAC057Wf42lPkkPEl6
gUdtseim9lK9B1fwAPNvTT8QFWo3OLBXwjnOzcdhDs78FHvccxoBed5Zmtczi47e
fJVoxWsCgl2YJ+3r+F5aeGoHAJvxt+URWGba8P87SsnY1XsS2+Uemd21BHDsP0Po
OgBtc6S54AmXsBUipE5170V2uTezLB/bEC27nSLhGg1XZR6BworVDUWsib+scH2m
xKKdfY4KB/ZAd8avuGa70MkRL7JqKkg/QiHyTWxH2SGQeu1Shu4ibGYdENpG2W3o
jSs9RsNPZVGXbEn9Y1zZXHX2eklYkKsbo8y8mMsVR+2/Bvn+IxHpHNgdcvLkEzKN
v9mMqGBCpevk4SbziUh1lTmsS9QjFhLzV60Sj0Byyioij6nKjc/VrYsm1T0eExWP
jX94zEUcOA1Ec/y7Zey4suj2ujXFqv+JPCpl+/SS4RoMEc8McgzMucfInLFjp0LB
Ol5xsVvIr5T18T3RLPLRTFoL9U8/GDuCk6ExB0JEgk/D0Mlg1ZY9P0W0bRoY5odu
SRMzqQHglNkOkyveQZtovW7OXJexEEf8pLTgEU9yUBtmNaA5v7UBrzziBPXvxsjA
8g01xnUbeKpyggDrqzt7A5JxrQLow2d7pCYD9rHCnVVacRhpzBxrAlCNw9bcWOA1
3xmIKmiPkhsZrfB+mE2S4NyqVhNF9wxNq9jjWVpFRIlA7JkpBFa9fAMxVyEvWzP3
VcCpW4oA5xVeaQsn1qBuls6qT9Xc/gFv8Z3CoaqzlxoQFJCjv4M+SnEBoPyWhFZp
9ey6lWLOQ3iu2lG2+ae03OqZxFJkK2X9lnLRrsrFpkJgls5/i/w8IY01wQufNj/9
IlQV3aDyTucEv+HHh8J9ZbT8TiMS/u2i79RAMAPa98P4SXVhTpT+4JqW38TJZYwm
1nxXzmhVayllK1PTsey+VkrJ0pzhYl66GGL0k00tergnM4M6JodvrHZerG2mAJOZ
KaFD5j8y0fAp47gTvfJbWvZNvCxPDAl8MXStUH7ThYKHi7+q1grqwIFusd2rSZTC
vuVSu9pPNJzg2aOlI4UuDbIrMbxK6zgt2Im0+OyNRhLBnxxgSw0RuP0lwFHV6NoR
6AWN3HDtCJV9aa1ZC9R/acVd7nnqSjbDPgV0OLDBK3yvuEXRIGvTliWlXnH0Qm1I
unWR/MUSTDkxHoq6/CRtmwRofbO9c6xxPsto42SUMVhgs7hoj4FSx2kVEc2lF/mY
17tjgxHPa2eWA+e64l7hKg34YqPFnikNhnhDDWtpoHlgooLai/Auc+vSOV/rYQsO
iNZTy9adFe5TsjPZPZBcu+JCbfoX0n6nXw5xFiOMqCEzwH6b+5oe6jhFgXIeNnN8
DE7PogY+WCaylwUuaVnBwlyddZk1fCRvGbyDJ9yIDD+cfBtsgW7I6E9X60jw6uhL
1j/8ffu1xtZBQkCc4Iv+yrb1iJChdqGGPjwhC1gBXf8hjpYxcfTOVnGY8HLWU5XV
WBHnMuHQjBUtapwUPlO6zYuZFEMlMijikrrxIUHmQEzX1yKQL/z4JYvXWi8pYdLa
eXHO7bPAzWXEAa1AVSebYU2JHZ4B4QwSFhNjheFFk48fauQu91RCGfgPiImPsixq
KJ5wotpAhxlqq7fajpOdKa+RsU9Ia5mZbW2usuZ45Fb2yATBJQ0J+g0t+qIjgtR/
fASmnP2S5InxD/Wb90a+GjRVlK/g4RFqyhzRHv9GFdtSOsU33hxET2foZZKhInpQ
LH7v80TroUnGbSmOkb7LdUNBCpil+RCPsQWsTO0owV65xQxgK1ZYop0GJL/HZyL6
3d1V8XTwkxuB2vHoFAPptFpbxZuNv2bqqdqQSBKZ+6fZdsXZ+RXJnjTOFn613DjF
9gtdbAJXq4aHDDkW7Z623iR+b8qMlViB9GKPPPIxBsswyZ7AJa68oX7fww/qmMcH
ZMgmgqcezO4xn7PISmPxHLM9FNOJcp2hqZP816VBB201qap24Lqxh1TIAfc5Bz1M
fhmIJOEgli+yMru5SO+KM4PLgXOiCwC0VtEMltgMFIeG+u7kLwNGlACXOyFfSIIC
GlgfrEEKIJgze4NNLRUn4FQ7AJ4UwZCzAb+3DT7KGJh972J2FzPskmh82oywuoE4
f3L4hR02jjbmL6BanF0SaBc0Xy3O10XkGHNMgWZ3TWQLIxexbtZJMb2HAF/TjfsR
ex/PALs37Q+zVIBIUg+5WFCH3Oa5m4pB7PaNWU2dLlD8cGo7smRI/NRtANCTsqAF
YCQaI2VhEGPWI4WD49OkzEqDodyDP1z/MMxL/3VDzlJ98bqPD7kvR61JQFVknWUB
BNFQHbWIgC+rVyhzrINMIDFDoSE+mZmPvxXE06pdWcxVYia2figNIN9ifU7ZJoVx
GL8Dwg2vNp/RHIpd+Tva4egvLrZEmRAlQagD36CNJKMOsg13gUq66VkcJynLtNe+
pclVU1VRnjzdXvrm/H0RRmckofyu94Cz/EEpFvrl/LghxfjhPebfczjlXdjnRtFe
JZPPhB0Z+8Wu55C03JYcNzYJjj5KvccbBMMK7MiUpXaIL20gei+gr41jR9XeUlTm
cLfpHFISKoPHV7m8DQfzCHuWSx1OG+zjvqqrT5REb7ZYUYdE1J2+7xUhabFxY+N+
eUw5PDM+36XK3U3zK31p7VJlUNVLH1mITBkjhpnTu4PKkRirlRJhafBEEWuJSnKr
yrfjVsuxS8dOITVjvzagWmSMz9iqhU2peggkHI9PmEva50f0XdUXFJKmk2U+vcHv
QLlY8HrY5Ppst/JvpDryUvOYgksV+XjRKXvqbByZ1cpag8IN87mO4lTWliUJdzup
ei+eBLamwuuefuBsad2ELhNo2Mp7RLxYAjPp3u45u4l+Es2sTtiVL+cP6F7o/SaI
Ip96yRxkJJ/7/6RpSmcRIAkLH+p7TyzyGYRl9kO80zT+8n47AIzW+AzEaVz9j6Or
y3GCAGYiO4ZVtsZRJm5X+eW0pr3/NnMkksVBY+OWLhsGWnr5M71HxzWpevZJpMov
c9zalyE8ZblwhHiMeQmZ5G3PFUdIXGh2n1L0dEE9K149vCnj4BADGiNBIDwW1meh
VNdve2tQa89YNAP64PsJ3kFUIl+mxQ4SjrKOOFYXqPpx1A0s87QKjhcpSnfPhwq2
znXObmMTwBRcclE/qsQpSeja0PFCI8OQr9EA/im/y0L5WIRGA+MZMcxcacZhXVJe
OTrOlATpWkLPZaXsAvMz3gq8Lo9h6YEG6tONidXR4CnmbhjAkvZY5aqJt4DLVPyh
UMHMuMErCEIP1Vb+k/BqwqPj+5KgR+tvVZMxdTkrF+ndOAsAuaSYWgfVD59k5ECL
Zig9m6qBj4CwaJ4nnnAdml7SWOWKSPZkqvL5FlJt9BZYaQ2G6Dtz+R+T8Xj0bSR7
yiLOFfyZSes6MGBuFP8LShq28weto2s1O5e9wEDCc75du69ltjHKd4tzbgiEig9C
icK0/wxN8PjP/kKD241auJVHlRYCZJdBgfcfu+c5nZsdMQR9F6Vf/GCDB4elWogX
gfPOTMRmg0/2C/sxrtQdjrm6LnidcO7BcctHu9rVlMdTIKmuQHfcWDHOpaNABLq+
uvN6SWaY4FhT0TmliucxF+A3Cw28asH1+0aOMPzZPyI8IaIbFnxDFKEj21DILIlm
8yuVneWZ5rsEMzSXeSWXCKbQwyKxEbHSLSfN4QDKKZETbxBT7KIF9hNfiBvopHiJ
/gM3GbVzs+4WlZ2uqxINthanGvjuvPHF5kVhSQbEwcvUz7ayCKdad9lfDlz2OCpP
7rgpx7BI6uUZMXaSAuymzeZp56z9Sf8rQ1pgtD0zLZUZWsPs+Hj5+jc3xOXneJ2l
H43ikrdTfSgYpHnnXfd3z6YlrDAgk3nJKhRKfSoywVOjfdr+NrMVnpc6z07cqbIf
Lod26zy85oL8AWhAMPu8YknKsy2SfSE6+6yNgWvIdZoCp2So/WmsDqXIV/ndJ0vj
xvz1Jf/0bRedgjn94C/MqR+8LvXKpzay/qllzQMeHBNyqdictrFvSz6pGnp+LFxr
iQ/WBkxmcljRCNSeu/I77bGXyD9bnLND4+22z0yYi+LCOPGsWbP4EpHJvlrhJNKJ
K9DdPTdxY9KTAQgnyxGN35t7lzHhIWs+lNEVgwI3t0E0zyH7S4EORMJz48XTPXj7
rsRoQJmrgQILpBcUayzuv5YbMjQyEP7WdJfoz7NFV3LPmwG9H6VMfbQuHxhReVbc
qeeArZMULmOowxVga4ROePv5Syn6Q+d2Nxh1cMP947RxRQiARkxUh14eKrUB3FLF
IlJE/mkgf936+6KKdutdfwb2oMpOkOyYFAmB0vZUgbZeFMWg/RvTV7awnZwD9r2y
XfBHZaxdGJ7VngHxA42SXk2BjUE0XgIDCubn5YinoV0v0x2EDfEyfAldfo9RAyi4
dfHMPGe5Go5JzPtYsCvyAEYWl+emLaCEips2lfqaZ0w2nWXKQJlq9vslzQqbgVxa
nBZruDRcn6sVqc3a6F4HqV2pbg4ABBVUv3PZ49avsKg8oguwFGrIAc/CMLqRYGv2
PFBIzixZppme0KQkxxgCNtjBpRhDpiWUeD+w107JISgKQ9Ulavmc9DyQh50rv2PT
cnzmpmOMNTTaGZWA758MsceCyuofGeD9B0Wfe+3uTK4WqqEWe2pQnbPvMGZezJt+
HGF0tBCkeqWE3yIv0g3OeqwYyTjtNSk0MFZQX/DMSAwAG8k/FPl2f5lF7SF91Jjc
z2H892mlHxJ9bZehqUPHI70I2fxIzq+ICXj8UJGG9ocWfeQxhShOtxkaentEKLEd
gqyBcMakcBZKWnouhEBOU7yF8M9BmHwrHIKkMDjbC1if2jNPFjAptVBLRC6Hw2we
kthiLq1h0o2j5eTTkqhDfAyNmf/aWImHN9v2rzOwAA9keN9A4EYDc21lJGLlHwF+
vpjyoo033HCANJFmUx1+9pARtzN9VJAieW9/NnfLNNwiveHA3R/kIgJ/x30q4gdq
Mq0gQVPpP3vClObOWFhwe1zaSyn1E8J5yz46cklnsYh2ptYdkVBElkrvfNzes75k
pQ7mN3dJ/RCCg0UDpso4uFXmz6gxEfkRi1VQvHnh+qWO5Td17mpTVFIyBPGIFyR2
Wnza1EcWyHMow3BTH6Os4ujLlbdx4YCQUQR6qE7wcrR4QkcQKufu8sWB+zvgmzG2
WzQdOQMSqKIvoG2Lo93pW5ujHlKHeSk1wx3XGQLR1FSOM/SCecmoEmDbuE/azEDw
fkZQnVqjDen3L0KZ+OO0wVKQyEa2Gt8Xfg+UoYdgCXrryjZrANa9cXy6TFhXI6w2
rSfjuzOS8rhYg28jSQg5PwoSw9D27FDJnuh7Uh4QZ+2BQQudFJjrMoI+jBux575u
oFyXw4Ub+3IvbkUYHh18ZPvgHf+43zwVqEWSkMBN3hwkDksXsN/15inBE/eD8CYU
GqFadziO3bzncuU6sK7huUY9/4kNZNoo0KBYJTW8YVIy57xny5JEniIQgpbswmXH
RxC4XCCl1gn6EFYPgfdlTAuy8/a037Xtluf6gmgKZqsPLoTYiqo+6piRIz9+8F0G
WlAFiI0btUE+43UNPDuMp7SFevLlyBUHNHbmM8/Zwe+6dHD6hOL0zJ7tsa/pfyt9
binkYiLcszvPaRaI043oX6AGzeRHlCMPFVUMGqSivuDPmX2hTBppiLACceu3o4oO
8iucWMfWJQDVxi9Hj6zKSCNUc39mx2mMj1Gf+2xZCWjj6glwBX+/AukIUDv0Y9gv
MO5/Wa4hmOHydU56hwLjYTt5PVPEiQYjCuBsdYRrhwIitBZVKTSvnbLxrszUn6gt
YJGkULSf/jLsFcJOtdBBpgiNJ0YACSM8XBfWe2crFCvpTNHA4SqV6zCNSlspAQlG
puHAgNylWvKEZd1a59OaNxD8VogorZ6ppP+2a9qGu1XF9DHbK9uCWBIzL0uDJDfz
3dHt7e23Wc+nimNZEV5HSNul+X9BD1fSGXXIGh4ZCgL98/mN6/0Bd9M0CRv7zLPg
3oKY8qKpTNj3YS4FdBUDxeacHZDKv+ChjVTBoknFtgo+RpuL5P0rr777C8Ao14gS
hFp78IaeJVjTPfzd8TRJ5/4uTRckqyCl/Ts/EESMRJ9UvQHHW6VKbMeIJ7dbtyy9
LXL8bs89dd8DDzgFRnFCCOkaCSRdtVIPEB3F0HJDmH5I4ySabley0cdQvZ1fXfiw
ODMueEpkYqfz5bXNddutwuu32M+GmtGlwY/O8zeBVy61b6tiBPzBET7uQjLLdTpQ
uQYuoddGhqAOt66yY+o4epRZGBnXUdqQfVQmslGuSkCspFiF9JH2LpwF/SZ5L2t4
MUTvyA1aiVYT1UJjStUsAPg8kRV2zSk/bCjqNcA1z3/wXnfBOWd7q1u5I9GAJQRF
uoQ/B+lNZJ6GBCo4FbILsxTS715RNGfZ6U+BOSN28l19UhgTX0t0jXVSCL0botdK
dt5lsD742Gs0RdS2+b7RRZBQpdNheogmMYxRi4YVOsKRnVpvkTrysY5hPTf2n4X5
S7ZMvSDpW/xVBGxa89fpiAKqhZDGy7EROr+KUFGt3WmJmAwq19C110jNUCX30NpH
eEdXYF55jsvLNF81KX15fFDYy2cqGH5gK2oN1rLsuO9/k00U+047i/qrZ4M7h2CS
C6OyEs2TsuW7K/65JdxiV/gufRNsJPEYsh3QMN/5xx4Y1eBfVglJplzInf/FfKmf
hTbS1giPNOXs4sEJERAe/qE7ZzpaA2zr4dykd0EWc2akp7pbXjc+cj3xGoA7/9tl
sKiNKpiDLWRCEiwfXstuksOnGhwtmJCjvWld8LbUME0piH44KH2l4eRAUpEAp/2Y
g4V5M7ljNy31RaZnAjvI3CmjOi/ulDAOZXxtXTPLaZLXMP1h6GV0F4OJjYgOyeLc
7Jb8belpiLhks+YVpCCeYG99UYw7XdnuDKaW8jPPb6iQx8PIjzVaTcMHE8+ntEMe
qEd3NVnlmkTuqC9/e5ZdhKiqZjv27CjmHNbPCyebT3nnCY6qs8sffO63NOH1Y9dx
st1a1APjvZzgUpAwvpL/sT3f2TZFYE6y4izPc4wAoOhez5eWDysntJZhqb6ndTHk
abR0i4QVDG9jG1W0uB3EEEPiXUSiWBopsBQHfF9ugrTG1Bp91o2ESkY0g4b2Ddxq
GuffeMYrIiXmtRrf86vn/kddrztrKsQ9fUs4teKCmN4PQEoznX0fIABv5WT71XqD
7VAzgRFRFKcjEu7aVFn64zavzwmH5iID3y07py+AwOqEhM5wIFb483jaXSUfLvTF
ur/ydjit8sJGeDJ+6b9uqgI1kZqM749Oy6FoDq3loW5ts7v87Yq+ZGRl8wFnki9x
zxmm4J3DxtQKSKurPdJSFP0RnZmv32chAbkNWBFnYJmc7/dm9xp/Lf7qvKX5YjON
Wyfy/KfWRmUgzHxTQ34mxh+LOgUSeFAhH98KA2WstyA4cJdpanMYCyQ5ZHPngkFS
x9KwxnX3FYEDsWq0jDEpIIxN4fFZtzUB96mviGjCc/ngz1pvOOUK7VlexVzIJI1Z
RIqndigArzHnkZJKqWDIf8G3UTT+ve2VlvozuKWAxd1I5J/IgbNA25wGxAwN6wgh
eCFzPujyeqdjLYwt7/vVsHzHL/Js3WjsYoXmAEgI0c6oldHEUP8fVe+9QeOKUKcM
spzKtB8u/6a2H/qSP8zQUWe3dso4xmbFcXo+N+L9WUKr676qqcwEMuqZ0wz1rpdV
J+jHuiKGH6HjmCDrLiVW11v/4mGsZEstONMjDBpBHv+JMXnXVKcAL3HXg0VjlZAH
xMAK9MCEQL25kObOeiEA3HDmSJ+AY+d/k5P6ZnXIV9LGgOPFqu8+ilXpRgdekfww
DiTDdKIJQkPC9pqLP8Oc7GqohaTUGMNMmCqNrpZHKV/DiuhY0Zes/f79ttk/UQsb
be3RjROTEshCjrVd8ZAv+sdjfNJ6JJGaefU3TM+lgn4C6o+yTpkZGQQXfYlE/WSz
f645mqt5GddbJ7sBQ6DJIVDqXRngccdD7UrkguhBj/ABrulu+ICWu62BzKNuED4u
1YagqZKeR6jBNHnHzIPayJEjFBcDJC70L6XHvdObMMk68dRe4LjJRd/Sfsd4g3d4
T3UlaKOYZADtbPAjrvltbNxKC0KEpo3ul/CQNsF3ro1UQxJrQRqWPe4NnNhnnetO
la+3lJeafIfZ0n62xI34EVLHWevg5CWk/h2nOwcZYnr7VAZSZ9LQksg6hVG5lhA8
gOJ1rY2SRpoKZujtq9JDFmR2UEk70Iz6BIc/0TwmCjqph22ZyG7fDs0NRStpfDKm
fWy6FGhcRomW9nAapTgTHP8wq/d8fccirh6Tw1/ps6fipjDOqQbD7PYKQ9jnLSTh
Z05jqo5Y4hcnFrcMtf+81Im7b7pRtRjJsrEOXqWPht23uiMlDUGDgmgtJGF6mtsc
Ffph7hs0klPt3ohT0XFD6BiiJCPf6/gyMtpevgn07eY+SlMjruAqRScbEC4RglI8
CRwNw0PQ7Aou8DvC6TDI+kXE9qjaVlp9IBfH+X56XrTac1g+nsJK3Ud2MW4cYz3Q
311hWKYhj09wrvEDPA6vpZCJ51GOkWHObalX9nSTYNF+IcUAnG1sTwAbUtQT+4rg
tcZlp0jyT7V9wMUfhqO/RV/MWoXZz9/4Ht3mAEgLdW9Zb7/fR/fQkWpRXWhmXJbi
EpO1zzj5G+uEPZ0wbl4qBnQ6qkMMVyn4naLnHctsRfc0a/ERg/onIJVZpKPXEFkJ
n92iq4551/jiTgy+OGJUHRjRPrJfqCqs1deTCC5kHmoc2tAMmqBGJwawQWKDTKAl
EljGORpxg+J+87P5MQQM7nC7Cw6i+BcgeT7yNODfoitiTsP9ClxP/a4vpSaeAxGw
mINHxj4+r2n2LHKtB9TjvPJh85rrSlMEjIagdQIImyYfGT88m+c9hMviPqOAc6Pi
eIh1jzhBQDknAiG0a2MN77Cb+LTOMykc+8LxTsX1h3eFE+qwQr+RdUU9LPEdW+8z
Usjv9hnZWwNDNCr35PaqS+IyuoyN+1pmC0tpJecwsAeNnQBTjL+8Ih4blkqPSmWF
txsT3qLkqNnxeeWBjeLsrYwVIfEdktwXOw+iVgdXXvFkblxRMfvmH+4amPdel0qk
j5KRF3ijQoxoUlh81R9ICHrYBCCYyALnoHkGZhyS/Rx03E9izP0wSMTD+TFVMwqi
Fu/qe+PZa08vgD57bO4PQdEpl7ECpwZa+f/yjvGDUm+7UX1eCsEW4TOsj3Z+6OpL
XYHVpIkt3liQeYp2Xmsy/03GmBpBxmKV/OnJGQYAyuRhaYXymEE4UjIv4hhmQHgE
yQiR5UEHkE2ufr8Zoq+HKE0TN7dhNpMnf6YaA0e6D4RPky8Kpu9A6IJhwBb5LQ0b
ut4Uo6wnsrZ1itaG3vU6tvsDJ9b7Io+xl+OQwN6M/YW3FWNN+A7zSFWbQlYtjL44
CT0cLGcVanEiqr5pFw7tWxy3upR46cpnmnuj1HxitnRHfuG71SiNNkHpYUUyYvVh
+D3Vo+d7jiluZhFRtAlBHSAKiIkRs5UH/zd+g5VMjk08uZQIo7Zb6OMTW5ikHZzF
rSUOJGazMeQ7lsm6v3D8kk+F5qxfVczwu4K8aHhADiUxTfc0EzebHEt9nUUjaFvV
Hi/Q7Qox9EKl0kvFZT0QgLTdEDfu9CtM3BFLvXGOZ51dr5AXABU2gCXqaqjEzRbb
Q7xk+fvt5TAJ8r7Ml6lRZ5kMJap6eIBgLZv7sg4laCErV55ZxO7W1gmguV2jugR2
D7fO2vNu98DEkcp1o7S/ADpdcPwZfaPqrACs8nWxZT+oY7ybUkyf331alAsIg8yU
v1ZqoxSoFDTtkc2Ck4D5ESmAiKLtyLoBoPs5OixaiAWGo+rNxztQkK5aoJEDOw3X
kgLtd/WHmLfc/oj/5O2OB8fgeL89UuZhUYiZUe3gNzvTfn7F56vGpGpen67akFvt
XkYLAiLp7FKlf8fNgWboHQqa52jis9aq83Y/i90iJvjABv9qsLxlVt1ifc23+Do5
P/lsPDozwEDFrFBCFyWpcY4Mxo1ln0pmrGdsHaOuf9WqitT7pk8AbEy5P0p2lMRt
1bBG6zDAT6DIqFVtA1n7f9rIniOEqO9jqZHorZSb9+A5uPiKu7d3uua7WyG38mSz
y2t3Rm8AQ3ilbRyf29/xDiM8/2Nc/ypbOXsciRX6FfZH/jHIspNGzV8g49tBjcf9
1M+NK6db8JAX/s0FVKQKpJBaFftzcCSqGE8P6er76ejWFUHqsTA81MtAOmb6r1oZ
IAcHesqpMxzX/PFIfuRmjpLkNNJVIBgvudW/MokfYyYuybSTM7R5os16wd3b+tpX
N+fbfBKH0/TnzTH8SL1XDkALS+Vn/Qj2amtyRFWV8tOhOakqtnR4lRyNwRd0gK4P
qgM1UJK9WdXsB8BmoPQrDvZ/R/Gyhuxecg3tzgJrDpwdCR06zSr8jYIjVTyOlJJk
htm+lNkfFi6iRo4klIBJ2MRlxYt3noJU2IgADECEjagoRywetQ6W4A7/3d22AQMo
MyozwMdul4DhW3ggopaOfuG1fHzgCVnJJUaYV9vj4UorfBZEmFHtrXPs9d+msl2C
eXv0d7cn4MyLWzv9CQBNqhYf8YoDoSAwdZ2lLN/foteULbuNKAYLY86lMzCMUn/Q
xBI9hxxbO9UodaqOxRkpDePR09gjBptoJdKRCDb0XHZiksJM25AQCtR6TnMXp9B6
uwd0Mgrp77VhByirTDajjkamwzWGRpBi6JpQUdDgmaxUmvvlfVCtdDTQ0YVc4GX5
Gi7gNbg+UDybpmYmnpqMtixowmGYwZ68t/6KPoU/wazMQ9/WeVd8R98apwzLUZpA
5OEWah3M4Ehn8RmWw0Pf4wrTjU1h8+qExWmEek7b50UFkO5YwrgNhApBh/ACCPUQ
E42YpgMGbeyhS3COIcPBasI2QaX5//+Xrna6gFjkvfCA3neMUPBl+xXZ90lr1D+e
gkI2znx4xghbvOWCOAnuK7w3kW9S7O6ye6SBkaTeojz0/madNN7aXXo/S4b6L8kc
eF+0kpLeveRJXc84KlrJMcSjIQcc7kTqL1PS2Yhwwyj7L51LPKD10OK3hak2SMXa
XYAOnZNOx5N2CsoowdpczSzuLmXwn8ed09se2qS3qQGifQwbaFhH3kXuHUpXtFdX
8XfizfOJ7MDH9pU2eGifAR9+imhi4t6ARSIuuSfcb3YkWPWCbM+ITTvcmh+YtQEE
MTkZ6x2BkTrcS+u4y1LmlhRji+2tLhaTDqXTnnuuE4mXBG3x+RJOXv9/NSIzwdmD
9sGF+BBVMOV3uh+Rrv2skiZdJVCi3kDcFUbv3OLyfurLRfp2E985YV1z9gx3o79x
pkjg3iQXJD+IUzSH4dUGzsBXQFxMlLENgIQwNSVrYzvkycuimFo0wPbslEHZDm3h
DbRcrYv0JhJ/YT+WmlhYPRYRCtNFf4LlWR/V//wVl+F2rqLCrSeLv1QkLsJM/i8k
7+2rrav7D/VzI6rhey7q1a+SMu1Kh/d6jpyab13Ysox/cpkJ/YQ7WuyI4NgICA4V
YBokjgZ1TPwEmBshHa4QEQ7O5galT/nDifOCg52lXhtbsv7FCaEl/v8l42d4MGJu
h1q5Iz8MCpxmXrWBwWRuoOTqvVmb2a9+F2yzKKHjOtALn3nVOPI0yhN9q6gP1PVF
yRjbksP1W2CvSkNvuRktZ6GX0E38qEYMGDTU0Q5etcjDV7OzJlJT4yZPQAESoQXd
L1RM8W8XPSgVipLPZIm1+ml554GEOry1HhdqiDPIaH9rqYgjCC14mubmpw2HKPqp
9aBAIVt0IXeG9DCcowr7zmYraHfAEdls6lDz/1S7+dee4kdX/oPXYYQ88UkqxysJ
EZFCC6ZQhHUoW6BcCIyi2JwS2w/OCwbuUx7AJ+On16v02ZPrToKqV35SJkkiOy/R
HvqyE3zJQi4iaWVHesGUA3CVjlnJydvO0UcweUxHILKyYda3eTRaRqmiSZw1LAMF
Sv0b8xUTA58h8xDdA106peG/MBKU04QIBbTTW+2FlZrrVAsC4xy4uu6T8JAJoG7+
IBViAHiUVkIIebbLdbNhl4lJuqJ8x2/AodIe/iCAAfRZ39KgdL7ouwDArVBecxSM
at7DpDnoyX2pEGnStDYz53AuIBalmyT/6uTx9vT/p3iuOhgjRFT7YtnbaYndjfq+
Tf89iJVxwhefujpVZq2RUE/IfuEypWC90a1l1O4NoHAaqL0IJQSLQmvmTo3wRKMQ
7PBc4CCQCrghRlg/kXHhp6hqa0R/2SuuYk3qg1GRl0f2vU3Lwd3lzOMuxxmCC9Dp
VWBNutFWT/FlOnujcrF1fKawG+v3puogXQsXILihh2/rY4EMSgt2WSz0wRx67p+1
v0P/EKZOkAWJmLGzAZ1MyjawOuuA1W02DbFbukM0efs78awyDIZx8Ve+z/XGjYLM
X5PyAlV6BaHEgX4W3zUZeDybpMjcfCafILphgScUgk3QBNNvdykoXyPwXAGzaqZt
491QQ/4mHm25LwWLIFwnnCAsFN3P0gHQsZXMIKFR0eO7QLBDTHZ/j4fH8U43svu+
0gRorwrYgzdmHP0lRiWEG1c2g1E8hoEVe24osiev3F3nnhvs14yhG/PzGbavb2f6
oz5ZBtkY9lEm98zR+L39c5PIFOfAa1OsRom/j0ucXnh4ztRPrPQQJ2aoxKpdvC8G
j3xVJ7lhT/1NNaorKF8XRqu5EO3nepz2FruiT+jarkUFN/5uLiXigmgVLvuDp73b
fu1qVgCr9ykmXgwB6zc3htVA6AGJjmRh0P5O7VzOgIEBnS+pXRDn8Xh6/d5v1rDd
qHIwerNM64ZoemRcB0x9BmVB9au8bkMV92IL+Utyu6FvthjwUiXJdj96lM5Xd4jg
wowrYG1kp1LOafniJQOWmThv1OW5wGBAN2io8mPot5JMDIhW7mo4xHRyrTbbVFiU
FWtrZDzRwiNUyvbghdS1zQwUd9jP72ljMGdCTVevLGI4FZk3o4SuE6JdV0Xske3Z
KsG65c46thtoy45e9AyJ7ZwfSjjkh6Q/isX3+EFzYgxvHvBTuZTCQiH/el3+gZob
JMBj2/B/EiuklB7NMmVu3ai/b8pslozbTEB26nkz/DKKoY+RwhUIUrCSn3lEbR3t
IMoB3RCmZqIRguYWlejde6y9f6iMjZKrqeb3D3zNbdOnSY84lpg8uvXqbSOfaGY6
XuNDFD/4zaVUtE9CFNEF2B4EFjsEVG2apvAeTLJpj/emVCAtWXtDvvg5tpIM5mGI
MDtT0TWhBkbpzy2ppxkBXg6cbDXxhvu42/reLFdnYKrxCtncQVTWJEDoQtTrTP69
pHThGA68Wv/qN1h+jcYq+1G6ZBV6vQYMSB6+UqCWQzaJdMQaT7YrrNLGZbf4NAxr
3hFpR429drsTdYaXaepM1J1ex4FFyCvO4bpvtFwkcnSASjfMrqBwWgeRVXr4pkp9
16KngHX2SOtcIaw4xZC0+Qe/Pb7kDc7h7UQ0kYBdkgmBML9kdXFHDGmJoBlTIUxx
fCOjnhsobJYAjMGjP1fW7o1YbAveuGs/AxtyFCr397casHq58oX5OQWHStXOvbo2
DvkPliSnZWnW2HvS5W2WZtK4u7QQkhDUBjp+FKaha3BeJazIMZ/xXWGwSN9FAFle
LiHIKGkXmAidKFQpucooLnvo3dATqSGMZH/myr3VeYZBCbwUdjzLu6uxFqLEKQCW
SWuDQUSpFe8CZzSSlilUQ7p8wRUghFzcZaPrPHvsiubdfjwQPzeh9cNiZ2+h1i26
gYEWwJyvV+k5Yr1aXOtXOqSB8E/nWE15QSEDVEzwhj12mEoJyf1/p5E8xKgVjhmo
b0cmLmhuJ7F7k1/0UtKxRa6jBMv4W0e9JDozJ/WLdvgvPqrFpG0ivN7xdwZDMg8R
JCwT4st56Ha0K5uik9/1Nj11uCa0Cdi4FqkueeH2tWZyKdihpeLSSYAIoFlce49g
ncWJovoa6kvof9L4Xvdak7FGnRJ2XHAVEjVNZSfZjTCMThbs2rN4w8qmhpIGhI1w
xrpFK8/K6KCHyKYsB7xObwJS0CrEDm+25vAatvZpTGOXEU/tllWrHuLnkAC0iWbO
e1VNdkT9vdX7CrFkKqBRq9imOGe5lRarzG6NEsdL4hFIVGmiH6qhzcMH7VaDe++A
NrQSc/Mkses5GFsYGnkrQ30VWVFx0ul+HmKuNUP1bzBQGiyIcO9EgppWNqhp66JJ
GvqcJ6TlBH8HozpOei/TewMzgJY43b68UqjBANQ9jYd6mVAiJAnWfZS00MMFS8Jj
XzAz1HbJVgHKsE2xPESk7sKe90Q91AMbuJrQQKdSpEh7HUCL1rPS3jfSGsglI03C
jTPRh/GP/N+M1VciSjWPtc5M7TFk7NSkjRDs0aLYU0FW7rgwKD4fzvPeMFv3oy7Z
J23MeSa6anlH/vMUb9XQchHxqHmVWCweaDok0Oegj4xk/WJqXB1r4jjrclN/81gj
bo15ms8LdM4q0xvyUD2VOv6AinTXa1cjOGWqQDyyFlQA7xiTUcTTmRdunP9OBfpt
koStjE+2K96dzkcYhNDhTM1fW1n4bAL/ovqQiqqdFV7iWR2bffKQmAnmTDTDKZn1
ZVPkrKSSh/aWm9bMzJGe6a/ZDZ/NzRItfHG9NZ6WWSvFvvcuwwhQPZkzK/jE2Q0B
xLa993XhDT30G1VNomViIUGR2LgSTRAhZR4l90emzgiTsiH23bFGar2ileSr4DNS
LvS0IaFyG3cM0cONEhPXDD04yUIsvmB16MuPRJ6K6Ey7eugMhAhbso2ou6kaJpL3
k/3Uyj+pWg4vLPe+c3mpf8zcoTn3UGpswducAO82CxY1xGJH2ZSDvZ8EYhgl6tOC
vTClguXGwAxKHKv65GbiQLv0FHp9wvvc9XQ0t1Ba3bskZUZ8db4IaeEa2TYTIWM0
KAcWnhwoODxSJFApxxwK0NiAtL5/mKW0oHzkXFBe1ysQGtzBQJTUwGiIP8+X9LKp
eUC9ymgXTy43It6DDz8s1B19ZE89/3P0EPiOyQLy4wSzAinmdspga5rK4wuh16dp
fjGaTc0pq1bNuw3G0VzpYIw0heplmZLl3eMzDxSuhhP2I0pubednLSdn+/RoGjgd
vEZEhpmA0A7UTXpeN1JmGp2yS4jNXUfy7kcqzCnkw74tHRdwtyMyvwvIebBYJvxB
C4KTV9ijZgoth9M0Pyl+AQBZr9xN+ym4jumjxV2ikz1R5X8zYdrF9+Ky7MS1CqRs
Au9NwzJXAwBBy0e5eTt99hx8F6/7orgHtNcJZ4cWXDqV3UvGE99y0hlVshw+I6rz
TG+XsTSuzer+5Syb0+zNXVpNeeu4NXwbAgbkrQF1nF1dJAYXbzBOpg8MOe81dkk+
uIVSqwCq8cMwvorYJtjl7gqSAi5U0c5yq/1MV+OHiG/HNfjihVM/c6UYT3VY93Au
n4m4uYjHJEaYgX0YE+2/j3EBB0MbSn8qH5XRXDQ4kVg969rpQgRx2faDdmR6E59K
/je5TeyFcb+N3yUtGAPkYRs453jYLe6X+95aQDqCXGB6Ph0+CZpEoUEEor5cVy6j
eXFJjkla9psXRbva8TohJ56ZBezRHtUwi8m0s5QPjMdyAgwGDNZjG1CFjfYQAYvH
W10vDF0d/RLMUHY2BYeHSNVQ7t7Axr1ot/KxkYhYmw+dZZNeGr33Y68ghNKRiIKx
kHUQE6O4y1WhsqTmunAvxVQ142CHBmMW+PqrbDdcp2ZtNCgpELDZTU+W1hIJEC5l
0chrFI+oxbXQbu1wMTaMXe1yq7kF9bTucR+oGl7sdT8s5GGYcfePp6WMZEp1wjQl
D6gH9cV7THmSoj7fQrPQBANrcn9ikQj0QcV5yfK0mh0EFR8Ln5wvshZtAouc8n7i
GBT3TONoFubYIpbJEKmmRs/PtkK62sYXu+0rCKcEgAqXSiWQbLsYgrwVo3ZjwGN5
GyW/JOF5QHQhVPgS7U7zRY8KdyI5FrrJV8UqzhQdxDjGStPAk+VETo7+rZM0DZoe
0xesKX8LEJ06NNquF9JA/wlMvfJ/RxCDSvjCAOw+foz8ed/TnJWgatsq9X1m1s09
zxVdBZMp3XtW2JVeIZhAI8QKg1BdmINNyUsdT0hEnpZjk/R/iPb8Cual56gdoUL0
9wGrMT/gM1H9yfzFbZJpSb8cqDGmw8MPjDDpBd2AB1AR4esCHSdQbxMCwcmsAy+L
gauczQtbXu0ovBh5TE0jea4KkRhhe+b5cTnxyPRroluV54HChEMzVqO0XejKPa9I
Ihd1j3s4mGsgOLCTeDrAzDNFE6gB7u35vICe+lW/ixK9y75fzmUcjGVuWhfaNnA1
gtAgrZkoWCj+cUk3nzO9W0dZy/MhuYxvfcSp/Cc86ws0fN2KAsFsPKGqN8az4vTy
ixBKs2S+AhDjLHFD9ifZ5vbnkYiI1zBFArExhgqhplGDHVevyattyxrXXHOGXXqE
zFEjRjWlzJakTL5R5iUy49CJal/t9715EyBCcGd7Hg/7lm7SjS0NtP9nhv45Gl8I
vCNFxkwpEaaF/H1Qgy7W8hhbaOM+dyvL93O0JR1Mt8m/SAgED0V3OwfnnVm7rZr8
uD+c6SQAD3deri7o6jAe036xCIWDnddsTMsq46LU1R6XxVtCxELjl4r4KezMHuTE
OaSMYmRntg4HyZkxt7MlhQoY47QvXtwdO7Qs4Bv8uUAMcnJLvKWgRD1E57tONSN3
JvsDHfDr/R95e4q5cy+35OhR92CM1MHjpULkkAP2Sb7gAOpk5yVC2R4vMpHd7CxQ
z3DEzr4LcvEj/egVpcxndbHhTpv0oG1zNheSP0KgmyNcWTc3z2CUmsfTxWrwGlT/
jNCxFueWE00pOuyXMuoshuC/dADe6HAL12EyI6xF2dMu6HFg58o4Et5ySpMtEPUI
2TE0BeuNoJva65kEMpkTciDR1S0F371QCcg67w1nNyAIJToCfB1nMGjDjrIZS+wl
AtEikRFDEZuPWo0VYSjwro8zA8powPiS0pIHVPar5RfHPVXeCN4J1pxA+MhEE1NU
4d6quhLa4tqlsYNn3qmKt39s0RBmEXwcH0AwIsd5zWbDFT8h4qIdfnhIYS+4IHRo
N2Xx8r++NGuNT5EFWs1NBS+8wlF71uuBg23lqc8dkH2NB2OeKY0MOzLhIHwAbFpk
RBaqEFhWbWISsUyldhpbygnu0n0grOFKbsuil+boC9Suz7C9J80ezK22GkO7tVWt
FnA6zId2EJMeG5iblsEV7ZXArcRRefY2MKQD8mnwn/Arjpf24IAMmhPVhvubgNUl
xfeUi5+SZvpkwd3BoIo00+dGkQx5gsKSTdSA+WmdpBH7f8tUlZuMKImsio5J+Bqj
Ts4j06XdJX0M2gDeJWBEIsY9ckZOMkh/4oy6UjDUK53Bdj/SYWMEr//eZpeA3+L1
g4J6pE4eRgJhJvdVg3O5wXhooo78U+k7hoJezGaLwuODSrHQFmBk12q9JdKVShsM
nEHENT7pXR2fKmjOg22Ip5RR7SLSl7ggdAb6m4cf7Qrg0r1JXoIn28r92fhVeuuu
j3oua14F6m7uZvWg5D0JXK/Z3ZGFvaOwbqiH3I5hQOMso31AdGxSgVaZtZHC8qfL
NVgOkJgDE7cUdmZ3ezAO98Vl+nx5JX2oezVzQuedRzxs3SLopipctdU313LaHFgq
M1jJrrX+LRyJqvHGwmvgivCEy42fLsxmiV3JrNIxO6cYVraDDEqhjTrTqb3NaXeA
A62onNUL7FWY/AFaWb8gO+Pz0+Mo+35oQiiHxECWhCxvZGwFGnwcT9R7u9oXvCrS
2n5VnyfUMpwXTyNGlgM4M776yLEnqZvlZEAVYeV+df1zfBaDdZkV6yedC+Uq3BBN
4pENK2l5NApuYMoBwqtEnKKJJ/Vh5suYPKyx4nLfTxHja91ZLIL8T1bhz66yTgiU
Pa+YxVnM1xEyCEPBqJLUvVcycgm0MuARR1kkxgEMkV8W8duaOx0VlhgcCU35kAMo
Ewxj+Zloap41+Hy+f5mHgLtZJAvrtCKSHvAg8MgpKj1ExGKT+rHpZ81pWq9Y5FC5
xL1EjpwqKbeqHstwFabOukX2GTdMtwP9u1C5YnxOwgKW2vq0PIcmtPZanWILm7VQ
f7wrw4ZUUqB3xZMmiN5RnLEY4Fk8lkDSHrpjz3FgIy6GUJW2TWv+4xfMXMQt942J
cLpNGOJW++lcFKagdKdeUT0N0iDRY/B+4d1uFtyfXvEhi0A2JL5QIdtFpAsI0dHQ
EiSmOypEK/BPMIL4AIyOznBwME/pstd2voAAq2d/xTSoZDOjMVFTaEMaDROfjoKD
lqXEYYm592sWkkhroEE6sbzZGNNTaNfC3+B7AY+K0g+oL9jNvc3vl7pPfBoI86Nw
NsljrDjlRoKDOENtKxfyuwKi87F8njUKbawtnxURFFjVP/79Di9rCYPGg5AxyehK
OnlJIFwRu2U/41o0cXr52w9dRyRIrTzBcUbcuz2ls7AD2z1EQbbje+pw5l/jwMAY
7OFpv3la7FaIK002HzAxsxelORdf8VUFkmBxV+o0Jw8uacWKSujyZJsFsXAZ8xrk
AqaPLSUX87v9vnAvchyrYv4nZs0QJ+gRfKBF/bJO653NyzQJ2ep7TaK976jvdKpK
sgBDdP8xCiR1JWbmVKCrD//6MC3NXQR8LZcfSyxXve+vOcFDPtJHIx8DffHZmj3Y
rzXGmbNS6IqlNN8BCFCDRcaALsRd72U7dhGgKA1vms46kDAcTj03SUfptaiR3NKG
5giJ0DYQKPVzbh6uiYuZe9rO/1VUSll0O0ou3gcAxY7DYy82xSwllFkaozptKkAV
NOJsXtsdaarrb5TViZoI0c3grqt2nsiwnTI/wbMuT+HhI7Wp4yLXHIztmOeJkdy6
2YmXvZ33pf+LiHR3r7/vbCGm+2+SULxn3FLBXbA9GqJ2TVnbvtHXIdVESblOcByC
0gzzUM7Vly7034SLJBcOpjz7NRgJ9PouV0c78RToDcyIoDLi8ZUVH4PBXGS+2cwG
8CwwKky8UZCV0JZN4nCC70I5Cm38hMQ8eymMHTSvkWf7tgdoYgYgwgQSjHydcUGQ
HYWZR8XmBJ7ssG9+9pK8FjXsu2TZu2gUlEYLQuQbq29Q9aFGHm3K+qdwjNvH28lV
6DIC+49RZIvAcSVkHlvXy+AQ37Bfyli9Rme1fFtmgcZiaRk/OBIiZn1tKOU+TjPU
Bn6Hg8/bHbMHAI+B04tdoO2JokonZy+TKQPklVNfLcxJ3ks9SPJE7IPuWLbrKIki
YAdiVDTZBdsR6Mx4iDp973vOQsAB/5LslIVvdFSWGFvLHo+9JuBPvz5cW4okz5ua
Rng5ZcTlwQIxoNtk4OXqwARlC+fjNdsGfWAIZZ8O5BCbyvDGfmnLARJPgUTFNDYY
17iAQcZX2Utz7AVlkTZ8MdAim9on62e8Kuzj3npKyOXuRY481BVGByNtsx3nytxz
aoGMPChf1yXQaZNQTJiZKQK6Cgv7dJN2MLNvmSdZ9MRDYuKr0hy4aev/lKWRiVW5
Vf0yV/4KbM2NOXddAdzyqUl2woT+iJrrxqNaiQcjV0j277w/pYruihPWg0cFbjX4
rPdoPdYDNH/uSaiaMfqRAt8F9KcMTHBX0psXDH8GDVzQwOny4xdewPBZZajX73jZ
yANIT93XxH635lHJRPM4FB2y5OklJrKfGLhAujUUEd8Xgir+QDskTDP2iJy0ksfg
V9XawdzrogPXtvpZtso7A4G0WHhQpmTd6D1riIQpZQ/wjCaZP3+QkWw/P9CW3T2t
qt9FoqQGc7EYvUjlkhwe4FEibqUeEoeE2JsG1aDJN818TdJOT506HDxJg0Giodo+
6fZzmIRxSp7sxygZ1Cl3mXa8r2+M0RWGdgKHbdgJhNbpBbjlUsEgudhoZZU73Xlr
5pm6prPSki8gASwBL6D54f+4mWKcPFbezjGCCyOzrQbCtxsRfzZa2HVWlxpz4aUK
xXFEQucTr5WjK9bEdrNOTFzp/Cie2Qs/v+mVzZnmXezS3gY2pUaXqfr27pboKMuj
XDmfxw6mkP2PxoiMoN7qNDsK/nmaU3yxRptMZZqgiGjtToSRf7uMZQ6KEJ4j4FUR
qgAuVYNkifENg5cWRjrEkiTc+ujAEl2sf1YWtRuxxwN/kKW3v3xBTIgcWAgCroK7
n3XC6GwRAB4nczS7cbU+RwOt/EkG9pcQdyJb2x9nLLU6Orl5GvreR//sY/wiwLfK
ccXpuwSzR4q8vAPOq6j8v+Y6X+V+HCLVfcWHmUTIuuQxF1jOazrm7jc2ki3aXw5l
QRdOxXCS2MdCXSOhMLVzw4ycKotUIYQJKPXUtP6mr5K4vpu+WdWyj3dnfQN7Ukzz
cm7agZTtnS3lFgJtj3GoXM4WTxztEdBvHTis3xRK5RC2UQUAM5s7yI8u8E/m36D5
xJUBTXjZSwNwqiiX+3cMhXSYwnecQH1u7g/QtoupJ5nY2cQgLeohmrP+ZnXUcqQQ
8ce9GK0aVK2MM0J2CDHH4fMRfSeR4bb+Vz5/G5TLHa+n7uvzusfZx9b/3OL6bsLN
wqZK4E4yAylyeIUWQ3sAwhoO5GWU45Uq/CgjK1VR6YDOcTWD3SegI1rwVQqSdL7m
I9hiHKCzMHV40IIiTF7KquVOT+WElGQ4W7jXBpq69KFQjvpDSK+8pv4u4gl00fGh
nowTYXhMPgGZNLHhjPOjLu2mZLu5xdgrtwJK/h5Mc6QYQ/aM5fER0vCeE488JFGv
FKBxmSmkjllssKJvJuw+NUATWqBY4zPTwS7UgntiG4zIFXr49ydU87xe3ngIxqIE
MyXbNYLjdfJX299PxSeJQ7QVuJXeDagwGe7BvfnKTqvV6zL+Bstw2kFlo5Oi2nwm
rFjQAzrdZeM5J5xfZTZQ4wwgpiUpzqJ/qBdu38GT6+VbadqB0M75oYmQulDon21b
HAKK3TcF0yenGMZhNczCTN+h/50DSoGaFhAldKEtQnA605/C7HiyT3mvyLHybjm0
SbIXmhlSr3Qc3+GctermdOIZeyvCS4am+mB+kVvJtAgu7OPlGHeuyQZpH/zaaE2f
dx4pcAs/Omgs9pFuMQWvyHkM8jCRw6hV/pxJfSm2HJdpNBSHVlX0CjlbWtee2h6z
yUIQCeTf+o+hFvP6kmnQhQjTdyn2gM6BwPeGxU6ZHSQ01qlQfVrBK3nOXR6WQTox
IS4ct4SRHFjPibBsSniT1S3A3q/bB6ycSO/tc8/p2YuLdi3DN6lgZboftiIjAzsc
57rPbYX4DGv3J8mpXuegrFM0coGUnzcrVM4AdOscPa/9goCGmWwj01R42NloVH5f
ZotId/CSUUROy4Ut/e7jFYb/bgTzk65oVFAYSn7682SXNCrPGqErZES8MVBtXvEf
EGHzax98H2j4RCJYH7yFa1qErHKZHTpm3wCuasEVwAWUH1r/6oZXW/NwfdqPZHkY
7fb7+TOkt1hcPVVorrUMPZZi0NhvjrjMXrhyCDcEYw3+cDvJLr1nxYEwRIrIn1uz
WWRjSUidDK87r6ppreXy5x+F6I+Dyg7/Zh2aXQtZrD7FEeqU+76TnWnvLzUMSvzA
xvwO6lfk/EuyRjr3O0Pg8gdBoNcd0Qz1tFzLwH6cmW3GIIBvTcjRLqka50cU37FS
McrzbQXzSkxz3XXs0FmOQUxsL0syBkGA4CYLj8ISpFmavRFw/8iqFNj7Em8mHIIO
7wlJ4AH/cZWCnnprFg0mD+X974VmeS+ONqlVotq60L+TL6QYqpqg+aPDl3OIdw1A
UTN5AvLCeJCi5xOpAmIfjCROUNVjKIW3lhSJmJX9gVoLUBk0ZPzxv6ysp0cVmmUm
q2xpCmR711F7P6DTFN0Setv4r3tiLPNQ5aCt6XikV7YGf5+DACynz0BLVKwxtbMH
yzPEXyHglmPmKCof6+yDorsWn62KgbcEJ1g98c1iLGtAAQQvjYovvccpmHT/ABtI
x099Mf/ZPU8rGb8YQZPVpr3SitfQ9dAWNQ3wKCSTAa9x2CQfPdPdSrtMoWtqOf1Q
kuOJKBS167j7xRT1xbMTOzqefd+DliI/rW90HmmoTluxPFvhzrqRZK93L+pfBOxY
dO++0Y0UbiLfd16KGv+yQjX4HteuLS1VzGCsLoNQqB2Kw5j+RsibNb+PIaEkigST
kiPumNQYSNFQsx+HbQ8hLqWd+WQVLCw4wMFDQg3ZkAPjNCiI+kFad2tlbnSEJuoI
Ynis4ewkshlBrVXwG51nDk63QSvG4bBSgzj8n2dSX+1sULtAJ39+Y0flIUBRM32z
YIfZUvri5JqShWQAErboFjyEjC2KeCW6f6x4yDR+LDBdLYfFZ24z3nWX8F3OsP5Z
pCMOnRcgnlWNnYaEy9/Y+RvWkx7aVS23SEIeHHICtJl9Gvf65QL3aTdWHNTTGugG
RvOkqkXjqpKLWo7nGWQJiDNngqjcKzPlNotVVGVyKBooTJCByHxrQhvDTwhdagtt
cWK0FWKVG0P4yt9LWgM2bvPN5W64cu8TeqrdteXC8a0fN/9llTaPctvfY6DqNplE
J/Gbzd6cJLYD/vpq2la6f4T1x+5jcZRSy1mEK31+m3hmxuN92B3Xpb+BOYABvrqz
36sNY98WfImJaSaod1JxkObbRW0k2/fxiOfiPkQbwoMsxtzxtH1zZjekX8eFMJx0
somKz6Zs9iNWNp4HTYEQWpl8Ql/ozYM9CeHq9CPBNsTvMZPcG8NqtNClN+CWmDav
+mUbeNw7YXfdZu5bjD3GblcHkfeybZcBnGkDw8Ww7YHpdlCg58BMZoizzyFTMWHn
HXnK6WGCANIqXlQ3bgct1MHkMH0k6Qc76ArJUrraYABsma4laBjt9HURdx8E//Xj
wNHcidlQhvQPm1KxRxU8ql2MrEpbwYzlEukocV1z+cZACNeIOwkEuUo+4qzmSxk6
qKJhvq9IMEVcM4Gcrq8T2PaR8PeD1RPti/Vid4duukFVNhy4AjJLT81M6R6vuvYT
uymmQqf+++wNeIsWIPijTQ4Pt7KA6nSIkuZp+Ao9HTiXk7JH25G7XMD3SyLry2ql
f6ggoyX+5miHh57RZ52x06OC/n8QW9T5sFaGyKcNt90Vjhc25Z8yKQG9OwXi9JQf
3CMWcf8iKQbIRg40BJqblphGbLDnmk9fX2fLUlJHplLmNvu/R0DVVG8vELW7vW/T
4KgXmy4jpvIHwkWRp5jSwT6BBu7TdgaVT8VHSCHF39bSYRiNfHvc9umrwKvz8N5Z
H2iPPY5WROld/3sTLCXajOlbbVNM3vvHHQ4WWjsCSjJksjy6L2rMVEKezL2zA7sc
+Sw0HDZRA8i6MlKqAAwruJ4ubuj3cyumh/q6xf6vjl82WGg3YlD537ZsYF6QjtNs
ZHwx0gk1BoWm2UWZ6XwdTyHwdx+/Fb2sBsHBGG7iTNHZrWcDuWqtM9QRDUtEcftF
uiG+lJpwCzWOhnFk1dHLy2Bn7eD7+LzR735CPfV4VdoXzRRKGgMnW1qx8ZI9ke5D
lnflnKsw3pXKOTiXFQ/HkB5FhN0IchVEtj7KL2pQet8U9C0xovB+H4NWhcPF3deD
6oiv48TqBoZqmb8gd/Se5HT3YUuourGTXTUePH/5v+iqhpj830g7wSGgzFwPhk73
8ie1hL8N44dQ1CHXunzb6Xxx/70qjiLu8xR4a3aMqzco+KEp7lzqQXOx9qzDXlKt
nZRrP9vuwTjDcebSVkF+peidSW4wd0+oYXcxNugMriwyy+dYUG6mibahf6mBDHFh
mXdlH7fI/gxp7xn79SFarKdw4CWkog55zmqQUyz34XxyVGvEEBWGlQTNdomgdt9q
Z3aZ6rxTWkJePiiuvNC/LBAXk4V2tfHpdgHIabFH+Z/Qlwc1uqiJMbfhyXAT48k6
F3melin2OYnKWjqUFe8TuVpcZ+k73xZqTrsNCAZLKSS3v1OHKOgH1++yOAlQtUe4
NdfsHjdR/3tGgQ7eFCckLXC5M2huQOnwHEF2wlbPXyLsKNx6/UvGyIfba9DIy17k
LNAvM7RDxUI0P5lwzuXTecHkQN5kOgseqLQGZ6aSXZMNlQpA1XFB4eEjX87dpi/E
XgVSUWnTx3zRydcyjA0rzJ5rTtSnwaRDhBBcb4xdVMuEGbL6dFUjNo8JkBem6wce
2sSABGwDtTBEZ66rT+qXISDEsRc5n7MgorGSsGXhdyrocjHWhfcU/1BUNf5Gq5Ny
GR8QpVm78NQOf4NDwjgWDDyxE6lDbIo0GYI+bFL2SDiJao9miw/tJV64FT47/ItM
zXlrGUI7kCUYqlBG2sKfVm7yDcDtbliH8bk6a1mts+q9Daecors8sm020/5hDTqy
4Hep0Ks05YFg3nBv4EJ+Wdo9wnmkl8+ddrTgE4BFDnJg8o3Opzz4p9/XXIPpfuex
SRrUx5tzs6b6viXmqI201djuQf3UAYcs2BEhgcd5Z+nFGPuBRqiPrHraCjByj8Am
wCoKynmQ8wCV2xb/L59l3VVG2uKVRUfum4gp0fyw30X15gZ3vqujhGGBXZ3DYGMP
VYDnYPypV59khnsQ0TgkEp4DyLLyYHpob9jeMmKA1I/Ngv7UuyAkHNrcghzxSLli
okLVrBkXCac6u2tusWPG8AmJ6YjKGd2eakgwi/gyipJ1h7SE1Bj+QbbUAjElukl/
yqqJLe6aq++gCbmp4QXn8JVnwJuISawuPVKycnlcsLcpxgwoAwlwvjiWTaWZNn52
ca8rVXDAfOLoyAR/6F/ighUs15VaoKCmc+MZ7Of1GAZuwNqj7t85P/sKnf+JBTNz
K1DGJL4IQilIhndT56PX4/pXrqveIwk2gIPFgnCIXSEYA5M9YyWwLWeU8e2Re5Km
AWTGnKSEdNwAp5Q0lYrnGEWutKAbO8nHf6hNOfhdLEskalq9Wsny+LzwyiaVfpo9
nWJ9uFnmJl6RUANaaWskuYdU+yqEXlwP07HxjoOgTcBCACoMHGMwxQ1/i1sFA55+
pou/qhK2UZcYTf/1KEAUrPr5MxJNbFMspHV0IjI90ene3QR67KbzNWX5IPMHd/fT
NuAO9FjVYWXkFyeCTUYDwPfxSmj88xI/5v58jH2izoAk7+msw88tADb+AUlFU2UK
4jkA3dFhnVZOny7r8K5QDgLMxh2xEOBhW/Hr7Emi5gZFHu1gy9tyC0+OtmLZmezl
kMqDKjIKPMj0+qk5ugMMf38l6BnHcNJH9vYP8FajbOzruPLefLf0/WQLQMA6KuL1
+V77yAiw/1FyaVugx6IEG9mmxztv9P5e15BWhjg+gXoIewyF2JiVcQdYbH2WhuGC
FP1mfBQ4pvET5TOgXtk/QbCPglbJGgb24fD9Uw30FTNPMyyfY8IWoN056rgnWM/t
uocE495ueoMIMVWoEi5TUjmXICMNI8u0nO3a+npFjiMxtzAXe0mzW0nHcQPlZxEG
YyBE/T5T7k+fjOp5u6RMvtsKcLLOkDN/xdRI9RS4RzXRo2IdhqmRoky7EQ4tzLz0
yVN4+4TBWw+BETkxTHgEFPMmUqt8TMy3eS5uVO5GMQfGQRZ/gL+13+aJsz7Vl68T
fFtgQGOz3ejgU6biBNGPt22BJOQO59lZD1g7omSvKkbt2sIFOrLICpo4pimCx/RY
JBph5LuuQho9GJlNzuWv7ZL0ffnX5V+mZa2ssMuClGuJaVhw710m4rju78cQBlzO
+FP3cWcJj+iaDKOfKuSGIWoX7s7KsYXsf4kS0Nvcr4I8kOkrGjmRCmklZMPX2KAG
weqt+p3yO2rzAs+j/RH5OXjON+i38zUzchomjQbWKk2dpX2ZSIL2wyDIDsMgVYDj
UFxed1wZ1IPlepGcLthPaup7KyiwL93Xunsx7gYzmERGNZINxgC64Xy+FppL/39P
91K5ulhAGy4pV6/EEyuCovgV1s3CQQq0o8wU69blL3nulG+JSrzqMI0v27E2ke0f
/kuIM1gVHvwoSK4L6/ICg08OSnGXcjerr7aFg9rDiNAWlKg4cBU8kp8xaRTuOPUD
xxdeknOHPPbiPS+uAXtNQlg7Ec44Pap/GZiq8cbMLHAsgXDYP5AVEfLEJd/Y0A3M
07f74NxGhwyn058xwdAUcCdClqBW8PkcKGDu/LBzglCR8FjLkIbjBrB5CzEekp/B
FMgftZUs8c91agXW2sHk5/skkmI9I1IXeSBJsu1GQWRNdPE0i9R3cv4cXqhKqWqo
X4zg3Yy5HiMP0vdpKoaOwD/96j1c230JTF+sTrdm42zOsUpHK22bAH8z/5x5AhuF
H2jrsRwX450YKzoNw2Xdf180aIShaw63F3jkHV6J06tNzrPdoHDqmKVwc8Ja+/cb
k2mSMNv1ApTTCBL+GIbsJOtXPMDJctJcQZSbs2qKa+66RLDyK0+TFEN284ncX+6y
cMaLUlbR/y8/wV+Ilni8+IOmEsX3ExOOssQ7wwl7YBPIQMKmu1Mx3UXaWBQOWRUg
4uZYhhGT0xPRdd4cnDwcDU9X9Nys8GNPDnqslMoqBYCsrAxmf2NCRn14RuMVImHb
I2wt1tItTTNsRfuBQFIZV16is7NuucfoUFsw9nrAPpvgTHb2nJdnaw1G4Dex1NiW
hOrVnPjRgckPAfj9Hce2SyZrEPYC6F9XHJ6SZb8SGH4/MiqTdtRr/rZuXz2kZQ7K
GvinQO4yCXhbiCV76UUnI7g9WV1eE5EBvqjzPYg8FMwbUkSb4iFL0O5Qlx7bQBLD
IUExFaxLUvgpjbR2auSg2uZfej9CaEL6HN55nJMeKLAniFtwnxcl/7tPHUWxaaur
+dqIrb/8x0X8ClQm0GqLybZvsSu35VOcZ6jhyizJb7eUpTPyJhzC1KJEbWOr2V+I
ie6whrG8lZP97a21QzqcZ6//bWotmfK3WnI9IecsbUbhV9+k8g8d44dX3pkDiTAV
nGY8dKGj50gN74bZ1mDyRVm3OBp1q6m/Pt5ArX4AdZENt/xVlj7Ur6KxSNGcCzNh
XY6T2h6kXzygUQvQBb72DL6mOEMHJGNBwrGIxaMt5u0+/J6hfhRrJgoazvGLxT8l
QBgEtyERjuWdKUoF5GbQ0YPiln10eWfEm0ELwsT3QvNrmAxPasLtxJbb5ClxnHdd
QUZoKPiVyRZdcGEQUt0gobBd272dr/+DqSRTYEZI8GMWyTn4QfB46++mvFCp90AU
w3A7Gm+i6n1x0ZfLwelRSuELNRdNHflPgHys5IeuJjWO6sBEgyU3Y2ri32v82Nxg
oz0gullHTY0q4wcEqSeJU7raeG3a3UrP0hWTgy19eqSGiO7ySE8kMISJkxk1PVe5
1L4gIyPsO0FZAV53Rqbw0ZbDZrfPJZ0cfqpZ/m2s2aqzgjEqck6g9F1evEimVmFs
Txeo6BX4lRa1KmWJ+PWs3+9se1DKKBG0e/bfsjx93tRKozs0RpLB0Ktc6LrTPJ5R
OzNPStA+CEhqlLmR35s6X3jceFRBH30Nauez8Fj+JPoz9uj/hzyAaAj2IgfUrYWV
nmX2jnCSqAgChG7D6lz3XVFqDYlPRzfeZNBdX8GAmNcKb5SptO29isEoX7sOfNHm
D5KwQSfjf8Z06MZs3txo3gQ1r5g7TBLANrEWryC52edFRe3bjQAyg4Eij/1GGuYh
1auf9zQ8Cc3pguzaCSJDroaq4Vtytrk+U3hq0AvtmKkV1ZksVkp/OcUvXdvTfUyF
qZKpn/bprnm83QYTbRiuWrU/N+2nyeCT7peONlj1k22bdOhXukAr4eshJuHKohUJ
iBHsFxrpLDME2uFl5QCwEC56+3mM33HfDbsA2PG3rQ1e8uaS3FlhS8WCT34tnR5I
R7Nig7bOTZKABsHlkW+bO9423Lu19tLCbNqc1pe3ws/Im+P3EszP/zqaCK7h6YqD
jA8UWuYgATX4NrCOxh5KMZZh33EbrEGLr0KPvlGAu7LqedKf8qCNdPmqGiTEzrGo
gTwrEsbimXAJK47JfvfMZNVg4PkZ/crMeCDpokOIHfSfzyEIhQJNmCmsQrrBwZz+
vHgkRERqMJSJ3gUbxaE25C2eKNnPL2WCEp2uww6G8B69TOSIFLz0FWK8K1p3ze7n
AtAwLyXmEtzX/cnUUmIjegVwOYKtzVtwvI5TdrThAAjHEOgVwn+FQL91/MDil2uT
JaFZ1ajXuMmvpUolOtpEz2kF/NO7J799k/r96vX1uuUaWALh/w+ghshDNDo7y57h
1Q750UzXVrc4ZliqXBod/v8lTncQQ4gJ/+JVFBKgtiDSLO490JZ6RPlV8ayykCjZ
PTfnF/efWrFNfqEs5BZkJARdUoXh5i3+moQRtx+eggWLpTq0XjhpqOmIwbMqR+ga
XmrT2uxNdw5PMP6qyApQ0ghWjHiMrW7QUorEon22tekTWTLrgjwCezI+cKIK8fZt
GS8RPr32VApVsYy1aTFSwWJgGOLAuRBHmV/SeqRTNAzZREL4daUsE9AOjvKRNJle
BhDqwWMVBO5zkvWkMhYiEFnjPmYDKf6GDRHJJMuIgP+B1AIghfTDQ6j7EL/7khTw
SgCiQcE5sg4nQTVBG0/DK74T+3z71FwQ/b8MqgaqoRJfVJCBiXGwBGN7usp2o1A3
pUXovSMq3qOPyh9XMuDDD3cOy0mxJjrexJrd/zRTg9LolsLNj51I9vIPtcNt71j7
JulaqRQBUxIx9YFXYKxxOA51n5H2GUT/rlxQlBnF0RFogRbcuxxHbrVCqA8yiGV8
FF9FJdKbmaqtv5B/xcXv7gVPw3jNetbHtdEcJpiPqbHraZEvu8lP8LootMgsUpUj
SKoEUQecB7Vm5/yjO/3bPZwjN22fyJ0d4x/h48REmcwkx1wDL29+xFJXj2/uUbqA
u0KNgMNqHFfRMoU9leL+N06BiMA1rRMadwdhv4qFTJzbjCtxkU1Zn1iTsejxZlmm
9lvXXDkE9fxlVtZV5l+Phq5dE6i7YNjv7/dkE5dFzuVapnV9oGZaOnLGfh1Bu0LW
cbnJoJ30EB71Xr08JlmSMnwNY4bG9yzZsgQ5IT18A5JWCGeMer2e4rwvNP4uFDF7
E76VSODxrk0vrz4vTtFiOQS5Ep5UHcB5MzaBN5zSLhYbWmjhrXFeyLY9XcvfR/kq
55vhrpyxrKomVjBq7Q6aBIo6lwjIF2c9Dn3DroUJE1qVB73zeCjcAenRXas1lQ+Y
8kRODiHKIMzuxDDa1S6TxSWeldel7xFFn7iHiEsZLcXRlIu7HUYm8rOxQW4z2FEO
KBCXSyOEdZlBUp4Qc9CS6twQ2EYDBHTWJ0mksQXfvJfNDfG37dujq7YQ5vrQWXbA
vQPnUROuFYemJ7Bjf+qBjGRZNreaSz6+WGzXRkwZlrKOsx/YzfYjRK1vC2O3rQW9
SC+2yPd/p0z14Mf6sAFG+FtllfWLsBFrQc/sXM4S5KF53gG90B9zcuo5iwgmH42N
QKwbCQJYub1AP9BjAuNrt+tyda0dfcSr2XGwjnmGzSh2ZytTM4hDGePO4d24pvND
Q0tedwwjo/zQcXejNm4KY6NRS7Ug2Tnq0iGsbHDgyx7OP0CBCKKSfxQb5al79pRZ
VWSXscALiayreWceoYJAKJb1xSrHRPKcPA7/5M++nEtWq6jXUapefA4PjAOZxvpS
1O9MDjID8KRvldXWLCR2OklNH/a9mesC/K7qAZJk9HYa1W2PkuRHF1zgjRBiTRiF
xOW0gUDyj9CvTqybFYdF3X1j6cEqdmZmRhxdLlukSpalA/+AcJbRme9fR8KCP6R5
6DDQhUuOm1/zjJFRH1ZdwSuiGbny+CIWohZbguYqINSSQ+aaz795Cc/5WK9FPwJc
fRAOARjhtNgTn28Gkycw4RoMVfn463CZAEzbLpGA7qX/DryA1ju0XDADEITScP/g
Y5P4r+sNwCWMqBe4AyRd6/QjQkimE6Bn9dwBYj6TuoYrRv8oDuxRfF4+6loDmiX/
8OuD1XVwvt6EwY76qV4UZ7uVxlz4z5g5IeJ0oVhkGlhSLCRlk2awPkSOeUrJ1Pce
kHrQxSEc4BBNKsi74sqTaRp9Y+punPmsEKimpYKCx+VriLNiXM3zJCv3KYttw0i7
O7eeWi5rAUYJa2ov9WYUp+vcwlIT3Q6hZAzT6dMa3j9XWCGufzvkDH8Iw4dYH7BT
u6MPoaESJQ+U2UnpfoHCsUhDyxQ/35pd24nitArnITxFEz5inlz0KjapAxLQe802
3vRjwKCFsxLGvYamqEfvZb9x6x458ggR/0OmJ3E21QOUk3ocbsB0YyRAqYsRKyK9
BIJcdHRCkuw7lDUGd+lkzMokFw2nOaTBPCR5fwQ0zVnrtc3pzU0Rdu6TuXR30Jho
qWpvnF2d0YAKGTnA9Om+tND80T7Kiq7BjVIEPvATZfx7IUHNFBSor761+/rqp/6w
4KYo5erCooCNrCBI81fjdRTQmAdtwUsJ1sRSHfJkp0MSV+DT/HFICRgKpPeQW6pU
EBkV09samuZb8dCC+DE64Ega96G9CWdulVg273pfxCzrPQBL1idvb0mJ0ZjdKGXw
n8GtGJrKQjlC3NRBnXXvXtvv6+zF3oQBuu17Z/zwJUN3vZ/3czNobzpx+j4rGcJ9
1pHdVkVBrKG2fVwrUYvBeVTwUt+SGy/CQtbidknwNdaLjfiLd6bvSzvdQQrfCLex
bbfDTiJX8uz1FKJrr7wrGDLfAi7VThxst+GFOwOJYWYZ/AlZGvuFuMIek7t6S9Ds
Jyyqt2kVod2SYGthqCweAkZtSf/zGakuK8W9ngo4ltI4dDrmG6JCjScP5XhDRK1N
7lHjQYbNzasGtXc8HtnhdeuLMEaMl9rPnPRoRDu7weL4dLdhO/Ohh8FDS1Z0+wiH
oQ0uhfVrKa0lmMm3fYW80RgdOeTyDyQravJezEpopa44rH/L1pqh5263gBj5ceDJ
n/dBuCMlioHx4vPEb7yI5s0CWNhjpOsSlNvslEaYIWy2LIFdbbSrp0J1W11dl+U6
nROBzN4UORGQWh+7pnIQTq8D+ZSCVRu4Hu3laZt6I671aal8j+iRXVbI/zS5BVc5
y92mT7CY8/WD3CRNa3RAs7zbkes4hFJ79HkSsHODMaqyQ5JnH4WLgopMXRC9sFAW
JD5r6S3RSsQLPjx5/A9YSCcWpyHb43JC2NuW/yaTMfgpA9Gvk8dvka7LccM/2SAN
qOcOGjudhZe3j4/Qo3aM6+eVCRFjPLxY47flAPpySBVqP96pnGXBBipPA7fBRDtn
3pkcqyYwrfa6hdq8OcUKwJpluyvh+fjHZfW4OeSo1o3iKy4EFwKA4PZa2wNUTRG6
tpnUwkAugmZpbx05BXdxAkFb8nZPDMBN7JbQHCivIcf+tgtlCnBQjl25IH8U4QZv
8lQzs1vZ/VeRh/ALkED6oGm6nwQaBbxtmplE48pdmg39SAUomZD/wTyQ/EQnaRg6
/znNSZA0JJDSbLmqgPL6vWWo9u0avCCBfZPAdM6lfLgMxQuklYyoJIpbd8/gUGzj
YfsSQEVxQTtJuZrTYFqv8hbGlta8Z+j2N6MFAjiwBxrzI9T4AUfxs4MLm8A9y7u0
iLH1e4Qbb4W35lbxl6VOSL9x/qA2zuXOl3cq1LvPdstKXS3j+Z2cDpmKJzfxWVk0
HqmW4NAWV/Bz6IlYO1vZk1ppD5gpV0FeJLz6mcN5GmlFg1gAl8WV8fSVaOehBg5F
uPlqQSfhVvLQHyLVMNfnoBW7z3KKHcUGBPkT+GhffAcvP5LkiAcx0QTM/1QcdcTp
XCzT+XqZOEzL75XDR9sKdOWNBS4baAwwDXCgHKz9od90pjBbjVVLRjhmXfgJ8EWV
YzKU5FA/hpkdQTa+5GVu153q14uCLbBfBzKPKLMOrZenbFlLdmU9x4k6F6/U79jp
6aXqoKvTy47PVwcvGeTBC3PJOb9SuPPdLiVYtTtUkmq9b3OjKHcZTmunLgo/H9e2
limAsIjsD80KINLO5Uq20U3dCNnuFF9rL4DiPfG9fQ0U0QtGhRJcEvNZbrJHkUez
ilStgpqMsW7+4mV6fSBMwY79slJWiTxd1ewDK92SufdxYrbvxnlQnpmbdeigKgev
XNA8joSV7TTjVTP+sx9NFSLwZ3rAN/IJiFOjONJ7dlE3mFFpp2Jp3qCzVfPBSaNC
22Eyq0NzqoQsyuTDc1AKp19TTQkwpU9mwrYgHuDIQPBczL7FyRspnlhPDeHVExsG
fjLrMisRCf5GnwYGnOC+p4rTo8qBaechbugPPxRaMh21/Rw7QNJMIx+Jn9SITNjl
ynxr+9h1zvhdTwFyjIDN5GJ80EDX4lbuoDhdBK9uqLG87qAR+WJvug5xfPv8CKg+
AuAlfzojl8sWMrCqrS+IutfgZ/fJ2zLqUVVdHsPyV1BhhdrmTob9gIQRA4/Y3SxL
QVNuUkZTrvnrnDL7qZ7p29p2/Ul2EW5NyB6Z+CeoGqxl2+KUkWf1LcXkpMntCAjp
RWgPSc7XVaV8BuSQHHCitWS9Iu6PpJvGMe6JW6psePugCx0F3ipZYfJmRVFPwXgZ
4VsKXjwuMYsAbGHsIRKHzMFDIoQePXnh/T4uTnwRQvuqDZtpsEys9mDZtpoPj/4N
SFuenUGX/5/mUBVlnh5oPiDiCYmcfxOpOclEPSeznjC8aOVn4+z4QcSfZYRux3AQ
NOhTCbFmyoOohX3W9TwO72HoaByrqLa0RAa+xbCqa2HmBgjFLpU1VtJ8A0kLv4Cu
3nq6b3OzJw6T6XJ5elw+zXrTSk2XudcjVgYV+lciJbaHaxOYG+SO9BVv1VTH6/FZ
W6Ng2keSiaJLA3wLLYRFj2/r3njEgs/58H2ZN42I12V2Wnu87ucUWxqHWEMg0yPR
bM4bfx2tNYpGBvYykUW047qrhFsW37dhGWflnO0XLwpw6qlIfygouAik8Tccpb/A
EF4voXSreuRTQjBcYNDf6REjL5r9AkQGJn58W8gUATWJIzmGyrVWQLqGhyDT/E+R
IlorlaAIgMQJX0kX/R1lDAQgRdy0U9rN2pOd0jTO6ech4HBL5abqTur82yDCPRqH
faPrd25z80narx4CeG3cJvP9qNVP0PgfE5rSGE4d+MjH/ifBmPoGhPqZMPHPNhcT
t1O+SkbZmkGYm5isKWYpXdmJmhr1dztZtMzm6zNB/Z30e5b2JVAmxSCq4CnW4SOw
lGU8afcuznLLcSvcvMxBfyuxVOxeKuXU+qQRr2ybIm/j6W7v81Srmwf7G3frJtV+
SEUhU2yMwUeKOv130AE3MYRJ3o/VlWE6Z+MNTv1bO8KzR5ISTNC1kAI0NiScnSlC
3POuhSJanO6JZLpc/BTayKpQmMB/uv2/sx96hkTEl0y9thqOv3IZbg8PsTeeMmtd
MxOChuCOTSoKq0WQ1JAalNRejAy2nP7Qlprzqm/4AGVqmXlySS72gzGgXqplqegj
NF6I58I8FkanqHDucY+rJ/EFeEQoMWJyud4wP1/dmEZ5ji9x8Vi0O2ftYSwl9FNP
37bX+H5BIYS+6hcJTIYfxRurJt9akE7yw2TodTwm20034FmTwqPrxbBI7oSqfo4B
4LndVtzsjtDgFuLhlExmYIEnpDHphbH5dS5BgKC9VAjRtALF7nug9EhpiMYC58y2
MhPwOpUFXl/WfaNBMd81kgtN0GV/cvPTHamFsgKvY3sCgBxxWyHrC7nhroEPD24J
2y64d9QHx3unhP6KcB+D4ap67ezaimWjBPuYHDphW+o7u90lax9v7gukRUt6bga1
J/yxm6ij2JwCL5auoonUWrTVeITnzTxGpMHQJ0MsPjYT0Pj3Iv64m2qssHT4xHdJ
lhA+ECqAn0dstn+lsCZQCYGF9sHlIRjQpQogbpvBaUXJ9vszVARQky75fxipfu01
yzh3RdG/o8MVIDInQEDIHhqZ1KXAOa4tr0qGBBRIAdD1LwVRZRTlCZ6uncSW6EGx
5Zolr4F8adVsCKYd6lw8R/IeDzd7lS1qdfWvgPUAj3ss4ZpQKVVOXaPuHwTbzuAC
lNYVJ4N5uLG5ASfmADVxd0ukkpH9ogFEqkOdaXHkxYwuqCwEcAlKzUWICcs3PlLA
N5BtlCPIx18RsqpajpYVbpfxKyc51B7iG7Un1wfS2xdnKWpi1TG+mZxQr/XZBDl4
O45YaA9+b0VKKrvjg4ntD01Wq9yDhO3Ef2Z5T7kLeM88WLVqatZR/i0TOOat89A8
wEJs3cpxfK69uhMUQPpvnebGRlwy+ibPyE/ztJYTHRYz+vHSfykTa+9rfm8Yy7lm
CC76Xlk/P07j++AJhuXqqT5Ub2lhBSptIbIw2h0ZaeSCCgm8Pjx9qXiwv6X+ioMu
An3GW5LdNnfh3XlMKglHddCa6ow6RxXynjQ7/5gSwpSYMHrQqGl47s2QAdAV5aIf
bKE+k4P3sF0Cm2jIbA7hTYZLy42xG0WmNW7kEn3GGu/IfqTbT58SECdcWiLbvyOy
FNAXC0bUXwTLWmr31VOM2RqUtx8HrPRi6l6nYEPQqaURY859e2P2gUKwXOOg6b7e
THc1PlssmFvBFEmwkm5cXOsFS6EpD3yoSRXnH7soHMa2AeR0jj58Wogz4NSyuE7T
++fK1e0iWT5vEPv7y3lZT7Y6I6hxg18PfNH5k8p8UzsUtXa0TaBRcZ3zdvN4D6FK
zg8Qq60JoHe45Ho549iDRN7iYYHZFnRT/QpGJJgZmkekhlzfvR5jonElxw8wIqIf
HCd58UjAUHWpGbtLV+S1f99PEuR8EhRBL3P6VpuQBU3bUoDV/IwmYP179XTC7oa/
unCUOtfcxX0r/+7lu+WabHoCqKSOT3FsEzR2HHtNV4n+2rjJlcv2sKOUQxA8nSX+
WZqavFdIuq6wcz0kejIxVKjVM88tDUvlUaNgR2m6/6EG1WKVyN73G/0fY2STKFWi
GHQXyJDiVWixnnGj7/UQtt+JFC0KFNdJ9Rm/N60zhibE8JFauReVHQJ7Qhru9ZqL
HvGnJYdIkDewFTrGEhVLFiJBaQTngZtvqqgOc4x2x9k+WwAOGWxFhKlNYtDjbrJZ
ejTU7TegFHgXew6EzjGsWnGy5oF2qm3baGYNbbjA516ueE9QHHydl0TMrDvRNpwK
KkdjekUYXiV6VNF2/yhGK5MBJNJQ56w+gyLDOmAIr5TCb1e3OP1884BjxrDpQBKz
gyXVqWc4X9aX93cVD9fPDGGF9qzQ/Hbocv2WKW+7C5VFY6qYfwIt2LIzqFgT1tGD
j78Wmm6cHi06/39SLueVoseuxOkAaZlOHxxs8H126FdAhujpP+oGnwWHwfozwOpq
PgwGb0uUwNFlvmqo9XrLvdI75iNwrPBmdE8nq33htWwVRyK7ftbIAD8TibUOZo8p
c1rXeYbhscG2w/q2sL6ItUWP7bu92OvsUW43wQyZ2jy8Ja6OzLauA7y/HG4NIrFD
5iluA1llfdnmHRenklXFFmhmNhQg8/YaV0omiQNO6A9aESvU5zIUXldkBgwr5AgA
TJbBgsPObpZhAgtu13TGvt9CBgg+THkuGj6SIxW71AVuY/ypXLT5meLOgNm0tItr
JobJJUyx0M/rPbR10Bkboh10wIozWBHEGl76MsrrEG81FGO3VfwBFK1+FMaEJ1ka
AeHBdOC1SPiiA9FElDFRth89hNtNywTdsb+Fm3aowdEKV96WIv1cZhvcFf3bfp9W
j533NeAoxdxLnn2WPb86ew/HNS5dFMTjYCRmCkPOUI3bHj/Ryc6Jt+kHit1N+BcV
ltyXtK33zYkzTVU+QqESWlS8dOX0KWiB3e/+aJplB/Lwzl7hPzKdgSodywfwoDQD
gUB5P2l2a/oP+46ZVaB2pZ4s/YOUG8QA5NpaiTkNByZ+rHM4r+j4L2ZT9Mkdpdc/
XCWtZSwSBxQYOftUrrERV9qG4Snv6iNlNBWXE8QobSqzSwM/WEKuEKZPrnJbGjke
iB9L1ozeaoV/uFAruaQctAAYLfUsjHNGXzi79c2G6iKABYp90hzOwetL0G7IXALA
VlejWdRwxtqVLIeQNpjbr/trLCZBJcmaefEQcY1N+98fnpL4TeEu2zTvGj9Gv98A
hk+zLxxjRiQOd/bEMs+SAvM0idkc1fj2cDU0fVLKShrE72raJEE8cg4SNIuujZ4K
gmvExESL7kyk0nJFqyDUPfeGV9ZmkcD3vkEredD9sseGZmMwSAqY//uqRNxPov/8
TYeotW3Lubk8nYr4JQwe0Mas6Oi/vjpv8wt1Gd3xdADMhzl5TtrvEoyCF2/vKKbZ
TQhRw5KmedKf4XzkRow6wTkD6zQh6X33XpFlUkf1FMgYtDLerxglcE5VQ3dvTC5L
Srus+TuM6Hu1Np/gaIQkVSrKB2qA0k2ICMlpFusC+GLnrfQdTJi+K7yAwb3BvQ8E
yU/ep3DxNqErlUkrdZPxmDSHhIs/OsT4OPZE1RXPi0tAQede+jIqS0tsAw8XnVLj
mx+c2s/UcH4CWcafZxoFu2xhCHHJcb44b/qxOUXY2NT/Rlf1EUIOO8GvLs6FND+E
lwAHindjSBiUKWdvou52QafUYkDI4A5oUUTtrL5yqZ3SJlYiStr4HruMHqIXRBz2
d3CON/P9FM0BPUEO5GYocv93AAphZ5lwKz382otVYB9RvuiIMex8EYFk+lk85Xgy
o83HZ+FdNfraCWf7BJcwreVa6uQHD0LM3v2HgAMrzFzE+/Pp1VLvgDfwvPz3aBR4
0tpX+TPlS4odIjN+ZzVfy5sAj1uTqwa5gl5XaOQlbvykzhlwwdjiV8Aej1oba49N
DaUogbsPqCEYuAZ/05fksuNtZh1FTPtFDjIhdLYu+1w3CqB7O5KNgyTD6oyea4TG
Pwz/sgdiEUFrBfumlBcCm3XoHrR6UzEmLHAYK6gR90kuPmuvhQbHulswEDkLcwma
N2R6Vplxl4KtBDSzXtcyvtfowJuC9NfsYyWWNZMua84580jfN1+fxxXF3kAVs8xH
RbH0TfAbkUeDnFlR18eNSHkdFmfdU0sEBjItMCRxqganQZ0ASzImhpS24SNQVyLf
JD89cc82eTutBdetDeghz1P1tpyu8NFrqOmg+IiawVBFJ+NtiUtuCKz6UyVz4fID
QUk1+i9CYgMqY9u+LWnTDm2/X4TRjvOd9J5bCcnMHABpNCKROSBiOoWR23gXC8wq
V+6al5c23gAB/otdKYLVQGd5Rqj9N/fGMQsCFGKME9BQkw0PGnabkbQw0xfMV4Q4
HxWcNBKXeK953qbjar9Ik+R9+GhrP976CmYTtsAyZvXwMBNxv+yAuar5hye0LD6r
YSfVEYG38KBTwAglSBQUN22TcNhUyMChQWTkZILqm8SLOAgAZTTj6IBz6ptgQM5f
GjH0RuCenhDbLFPgQLKy308GxG/W66650ZefBWbe8sKM9YN9/hnHlq4i5oIoDagn
LpMkELVm/FGQs+DJfY/czSp34Jyoxz18ily9/OQELhrFe7x/i2xKe7QkmWInk8PO
mQrVpu0bjC/x8EZH/5NOqOAUvjjSNO1YDb5d2t6+LojSclRtUKYyfXu0N2hoyjcX
aelu3mtgkLJP2ACJPWNk6J1dlHADSMcOR1UIG9JL1n1HRAW/xbPrRixYxWIpNyWk
4Ej5kazvdkAGyzsbZVbDi6VpoAmP4Qr57519w/fffvxdrDSUQsXOvLxpGwIPJ5cQ
UN9Ollh0DWD5FZTGZvpISBqpqaR5HwrFEn88WjwSEq9Q55l1+EiF2w01WXpxRzEU
C3A7W1R36pEh7xgQKBpnI+H7R1DiKN+2YxqAofB7e6YYhX7A0YmnYKXxybMr6adj
v/krXuXrWqQlK4lCVJiWqIQZinHDmZksccqmbZ3AC5nZsVlq0j1xh8I7mhceat9I
zFu+FQ/CwouSPWiGYsm1K8lkNMwXdVdvsYXq15CjicQOyRNCPsrh35ENrEqO5uON
syDRp+UmubMY4hZ9yxAWJKvchQEQmjDKMMS9Bhr9hsiFXCnQqp2mUngOHOQYshuj
yIwV+GDa9QkK4OFiCbq8bIfESBFpmg8M9zksJwN4DlQHq7cAltXCnG69TxGIaYhg
VPtjxpXZHLlSN/Ujv2IhZ1UOVM0H1Fli4XQXczo8uxdG2oCpx8ZwW4UHFrVuZmp/
Ajf4UJwXIKkR49z7Yc45gfY5OKIh40AoWPCSuTWzZaPfuj9is/cwqQ1qdCEkIwBo
SS5PyIMP+Mcm+naF8QdoEUfKI6VVXIbtle7NG/dFuaIjLecDxoLlZdl4wiDoKeV+
W+qYDgHczTh8cQmCqLfdymROiuizWmnQ9kUyRAmRzXlSTOPEXdpUV+3UT/8OMToU
jBMjJJSWphqMNbTraO3GJLUwDVStMLC7XYSpk0qpPLj1fR/JLbRfMZvY4K615BZH
4LH+aUZLo9WEqvVFVYtHYIfG2J5VkpLVyk2/uK9+JIjHIIPpwnq+t067Eu/X2g6S
eISQft27ibOuVZt/gZrtSCsSUW2zhJ2jjbSCmcNWrtw/35Wxm6+Be9IbXGVOyJRH
Yo2b8DRMIC85DhBkp/Ec2VJSTYu3pM4YMyG51LClAB2FnzMaJq5M9gQ3kAU0NOLr
SpepaE5caOxs3kUmcqYm6TgbgUwZZPTRgBCPpkNCcPBen0Lmhu5lbij201R95MsR
jRokjntsX5KHbUu6iYiKeduYESxSWemWk3q2UurB59uxh6lRbveHYlCpDbIWi3Mi
JQAxJF1GN/zqZEx5M9qqWW2lHArUjbuhAyA9Wh24yGKlMl0UVIPMfdCsalWuo1R4
FGjvohZL7h0B4cuS6/37Nqdt9z6PgBb/eGXzAvH1FKyg7byNUCiZPkv8T69i1NcL
4vsTdD3B9fEJarY2vaI2+9XRkDgMP5laa04u/VNAN5kAGIn06ufqwc8erPUw/Qtk
AnjnGtQZEq4i7OPVw3glRuvHPzvh2fyfkSQGksCDePL5FZp4eKWVxJeKF9dIED8Q
bzxFAkUG6kNjN7wZYfeMw4VwAbTyOJ5v/LlBbM1zPk2lUxBaW7Nl6lCKfpy1z0Ot
H2O5obOqF/A7u+rZH8IUR++usWXl5p/7Ye9hBFerb4/lt0Lvvi57bNSWQQt+M21h
fhEuSPegsxrfPwWVkvDrZJRLHpT9NiMAHgIHgNtDrDUynv/x0OhpyroN5mkO9AFy
O/Dtt+NqyAbksqtscwrFWswCuztPECj/l9V9QyD0qxSdKGEkAWTJMuxo94SStlzM
zrmg0Vq4NuiKDSuWoBbYAUbsZoCOLsQtE5T5/Q3jNZmuY/lMug4hF6WvZCtKw6B8
8vUvdnXI9YgHSVdje4FXU+ktdCYjljPkhiQwAoWEDg0Z7EKyab8+/W/AWlhIIar4
HYCi5y688pPn1MHPwvygxUEyerNOtZouKygONMxJZNQFQq3DoG4P0Vplv1FiK6IV
9/ONSUiov0AS5qn/d/HtDW1J/Q9XcEddFl+r0qBmcrDl1p2gO/M5qASeMu0QgByG
/9U/21NV6fUkOZnctE/YcLJfPlxSI38j9X2m6Quv5ExcfOj0LX9PYJknA5sJca7g
+XCpANC7azbXu7VWoGPxWmBGmKL6EBTWFMIcOdoJ7ypVavWBHan6rRJROGEhYf8M
v8I8Bi4fy2kukeNdxOwGF+B5L/fWWPF27lBhiqQ2daIva56ly9CWf1VhKfFc+gh4
HlrBe5L4WroJ2ymjVd3wLcp3+d2KTN30dPhmVffT8lGJqlvZU37okRdF/vLpvbpr
F/pCG36PAZYyyT+c9rTsP72XMYqiQiOYPKi6Pbg2yHmKqpldbGxkRromZaXS+f8L
QbkyS+x0GUN7iACOckJT/mzJIx82/a2V8tpP4BT4/qmbDDk/U+DlWmh2rThkt3Km
GhJe95p3tSypeHM5b5E/DSP0SGiD+i4x+ZaHClOJ5SUGEaebz0DfvyRQQoPAtri3
JpwaBvJXyOO25CcgRGTNS2BB9AfhGMhMjNQbe4Z0YwanqMifimwiDQudMEShpFL1
+mcxO+/BcG3YuFbBaw6ovwlW7eo/zJCR9I7ZDuCUQ0DwVhRUgsn9TcHJWKKK18qX
Lzwak1HfJPAWVsSfqB0V5AIkW4VnE0NuS/D9/KQhZIkhPoJthC+tjf+iUwB4FXNu
F6o5WZq2pTlcmNCvchfNs8FSeZGC2GqSYmyz8Dd0SDXnkGuI1oibUzLcgys8q61s
FGeaEflbz8qW9KXwDd7XszpaaLL1SyfvI+IVS9/5VR4MYJ6ZINfMzvG5lNxEBlhM
mtildYaHpbv59DN+EeS2D9hQlKbsAYp0Opcc+VOy5Jhw1qahy2b8etrNrxShRwgC
spQQm5tvgsHya913q5n9HVg3ieT88+dIvMTlHBTsVRPvJ9pGkXClAxNnN5xZaoMs
yhBEHX1zv/DCfZHyAAZ/+ORYS4x98zZWnNlFcUCE1r9O7mMv43fzXpgrY3T/r70Q
2c8qfg+iSNWF5Rhn9AYxH3Y6eRYJeIT7sqApSl+ru0dTRgiqZqI6WQXGrTfgYeww
pDe0iy8eWhrzSOXh9pe7qMUfk7dDHHzEhcje6eTwp0P75rQ8brkIQP3byVI5X2it
CGu2rwXzspy1n75H1uML4c8ucUR9PqbRI4eT0qRIQSaQDSGpL+ABsgAzosO+f9Dm
oAP4NhERoh6G/ZIZED7e0BPTQde1DS8XYSLjvlmKKn/xdD294GW9pZKjQdv3tc9S
q2NPaqv4HbcBt1BwuGXL4cXgjSsst2QacZKYoOJyFdE3pIKP1SvDdXQkn761cNHU
8P9vtMohw2cxvBYYs3whnlJeHabbs2OyEQqGKbZy1Wn34RKdobaqR98BceYsAPxM
QmgEtZzGjtBySFJPouVna6X31ZOa3WXouh8arFhY8E5Db6nSoi6leHzyjLmqfwcD
F4fVdPrxIWjTRJG+x01mpZQuJLuU/e1LfMbc6quTfShR29JoHFOltUsm07Ucs1pB
q/tpurT4AAhXi9/fDZFz9FX6P8J2WquoDPAO6Ya/80+rNBi5HeNafJu9m7XkqyRQ
0vL5Nh8siU4kxV75XMqQZmyhvXyTh7ztgqXoZQRMUc9SMT0uCCJipcmEZSb0YoZJ
i4FXHw92AWAXynaYyhGf7+QJyEQYfgo4pqwHnMpbF1byKZgWncRRFhr+3+n4YKwY
fWdek55PKZCN1DWZcC411uKqNPW3m7gvqvex6iWhvPntNaZsCZa2529exdjMGz52
6RP9Cb5sqR0CQzzi2ITS40dN+shHo/N10SVynyxWQPPoE3TTf84Hp7VQk1BlqQH7
ttIIth2msKbHBHh5Ic5v6H8ClyaDMeg4IRf7CwJaLexFyKMdjCbI+Zhrloxjk1yW
xZ6KVNC+rsaUW3RD/Xq+6Nt4XAZhaUmGfvyEqiqib0A84c5ZcwROGy+p/a3lwSRs
dKAaz6I0BXnfOUVDfPjLydo5R6xiMlhBJq/yuGrDEP2V7cJyeTT/LGEFktQqMxUN
YpxC5tx3wq+LHsF+K/RmzAc8fYyG83HP5n+EuT0ZjpfPhSCNfqvcAmmHEpOxNDu2
96AxEPKSqKbb4fUKKzMPDJTfruIQuBhIPCwrwNuFzUsqrxadZSw0qmwBmetlCiAz
ysKGZdWhSfPg0pfFLbCJj0gDoaAD0j4KqhC0L2Kl0W/BKewWHChPduQqMpn+C+s7
KXb0NJYBqKiuYnl/r1/NEVjJWtmxl9sbe9r4emNGoyw5djFWswWxraUfJRnPKeOW
pzGJGkGrCRxS2VqeDiR25eL+xAnq3SfEqC91k4P9X62MX3p261UiqzZlJFxhwLXJ
/CkBk+iOdsSI196Ijk4WQ6CW68VS0e8AYlBq8LZmXaX5Tz1vx+hM5npdHj7qq9O1
F3Lr1kaqIfvak+4AbzOAF1dtCPpnkOAj63lG89vnBVrpVBqRjvwX4QvFQWArtTuI
1uSbros7K0KyIvxvElIFsdSRpPj/QlN4mw/85wtZn6TsQBmmMOhAScrAdMQRjbg0
fFRdq6iM8kT54iAm25Js5SvM6/bZltheiE4wLUOefbiidpluc49FFHYOMcuRyqP5
gpld98+LTL/oYP2jo6zq7qtSFfjZHtKbyewRgJsbFGJu0UXBb1DzTpD0wTWT5fco
3eZHvFNQ7tReye9+Tppa8rSYcXZQ7OBWEfQz1StllrJB9HRm9cWr8Oa5pz8lU13b
PBfbMqK/gTxzZsUKO3s+rG9wDpk1BXvQtpUqFyqOP839aIz5rrM4Zq7Hj+L/xBse
ZkQh1naa7sWgxuPTzrDXjBw97aMzvrf41HiwrB9M9ovytK1OlgH4MitGTDzxeXMz
WGq2evhphL7uhfptJqiOnTJRXDsncHlUkzHUoabywwQ+RuYTqPMSXld0Jm59VSfk
q8KetNo5MVW91HYSVHP+BncbFSM3dEzcFHk/atFzRA/8zUsyy00n6DSL/VtQHgoJ
wnv2uKaunyNlA5D+phv5y1sSpXOm5fb8+ZyjLDPxwrGOd5IIVNcI8/ptcS18LfhS
mqy2ebGsmCeHFKRxiwjoaT0Q2s33Nz+Y7/ZkEYkRepKKEdQQOdmVHUCSeSi28AGU
LjOcDpnvy3DX51Af2mRN4nXJjaHClYothhI8Xn6/TXMxjPW2XiO48tzvPl2XGF0P
QD9tf+d82zu+8xnox5+ZvMUG5HlkuDZ5OAxbxHXMK5ESvB+CJqVn7ckG3VKHYkGU
k9lmUprurGkvTpdkXJWa2dHhQjuqob0DONe4CHxy+dtL0+2IxP69IUYaqY4t53Lr
+f/Lyih/C0BhtdwYRDttYPnJWUUnczalOFkYmZKRNNsZAD+o875w0mTygm3pqApa
5EBiYb7M8O6WZYcn/Ae+uHZR47q4vol2DF2yAfhnF4lcGXbeoqyei1nxcDVt4szO
0Q9jjQK26im+Z4vJA6zstQdtuGrPn3rICHWaHoFmC7/UebELeKqk8MPbQ1wsw+H4
nhc/PCfnndhEldDZ1VdVdyjxrRRtXNCMiPOnx4BmUdRx5SrPUdKzi4O64pHLQ/BA
uLe9fdCDkjvG1/AMZMZmhey5OgXK+a0m6CIOYCgidkPR2m8fzPxDdXelI3lF2wRI
1y4MZbm6JJN38IpfOazkYGZm5UZVTAy7U5bvI77b6ASfK+nJUs1znnYrFnSG+G4x
XIcAoEFOLgunkwf1SZ5BwqHhUTIT1gImQ4ccYI8lGOTSpN6AEEKvko5FP7gSGgcO
5bTovtJuGGYqALJ21iyXHBH5MHlvAh8JJMChFplBEN1t9KmarANGIAEJQy88CrOI
ChMFJKVGio7ehX6hkJBb9U8by3pSRWX9OT4VZQRrydfpz1yaXgWHcP9s8nLeLVP0
UEicUyhdVFR10diF012fSAURc5bhkSgU7Jds4IYbGsFG6JasGHhruRFjJvpK3CYz
UPvMcqCbmTc5o3pKKlxTHbjK2DQzqPjG5t+B4ArDucmYY9Zeo5dI24M7aN3udi/D
4YmM3vX1pY7PQQVl2uf5raqZTfC/unPmSVb0RB7dCLkGmKPTnWCVGYsEMQCpkH9f
P+aBLgHPKyRzjjYvZecN2VydiSInD2GyvrYAPDik8Wr3lsXdPzyW7NEO3HjcmU3I
BRk1Z/DHD5WLffubh9bHIMbeJUAEHCWfGIC2tOmSLtlQ2Vvto6RZRSxaZLzpLMXg
rfH6MLjfqiRzOvg4TWkDTNx7cQhHevuqdV+wZ3GhocEdhnpA47jHpldTRKzBPKoA
IvfsVJIgwMXmTSR3D5hnlU4xZTU+S0RCb6qt0WVvrVxr3XaLeYSacWvpoffqI7nE
ramkPWaRZ3/rTAtw3B+cNrbYJCg+s6fhHidAkQn/1iWll+WEUenkfZfVyv/Imct2
uDdKj7lgz7fYmy1RN72zHqsMkR/xEhkMj3HCvqjRKYpwRprNN+cajAl4TMsrcO+7
eVQboMVEuedV52p5GCjkdJ4qqvx0K7hqvNS+fONxi+RMqtkQZLhdGdNbBwuQMuI+
jXfsPSWiF6Dm3XOrCNsy2d21JugqyjtNcil6FTikYhq23xMW7ENhIF21zJeNoHel
+XwpsSmP4IryugLmQEvnk2HGlLzByF+MaIFQGdY7EXoVJcsHoc4p7GrvWgmQy7E3
gp1vhpezPISpibNoZR3ISQGM4Mf6MvnohzKjOevJF8rCU5AgQdRTcV2r+cZgxSQ/
woi4b+J+f9EvjKpKq9ZUO0cu6SnFD6fvVyMUsa9PJroJcFmPci83Kf24WQf+UVBT
GFEVWxr4vuMYvWO8/fIxpOC7oRzCK0OmdZhF65w0b4ys6mkI1beCZNMxCOg53aXn
/upEydT8OIZLWRbdzDyREUPgVAwV4OYvdYS1hSSefpguoowVqriGbLdlF6yp2lQq
xe4DqAWGYMNn8M63AkuMGrysX/2FmEE+phJJG14z/j8i/EkiJZ6CzfTuJ+uPhXDH
rh8kCAgFrtFY+D734xjCIqkT08ViLlBJLCKFLg8Om9rOWOWkF8xviowBj03Maetv
9rQTklg3vsVmKp+BdzHJC55LLGXZQJK7NNvZXdKIc5VF1tgOobIDeYxrTYlTNUgz
NOTMtQvKfuwK0QEVQ8VOMraPjAJPa6K351/yRpybyBwk4P7rbXgIeWrkDFHuRGhB
qCiYVh0OFE9YX5pPn9fd0Q2aDnao71W54h5pOnV66gHfHy051tVU6uDFcV74H3Rf
5HA7PQEP54ef0g3ruVmI9apHwDW/creUe2FjNB5g6npQhnDIXqEbYnTih9rnTbNS
0c8lAM0ZzgpPs2AbWUnm1FVx+GSDT9grvDv1wWwqVmVPhuXVghRHBLSuSDKrV1IQ
6C9RlVIgYerl1PlqXUksG7QphZWqOMoKr+ga8wa6NW8uh2to5tXW150a3jUq5asA
7IgW9CmbQtBz2xS2AyYT3UszybHmotr/hYlc8TLEzqsFm2McG/A3zRetSgVbxH+Z
gs5wowssZkIclt+NaAs+cqLIwAXqFnJxlz6TsOnVhG8vrwTnXcMIiqVknH1G9BtY
KskLUJdHMM8JsMF85whUKZXrJxQnRDHKp4eKe5EvFm+NonAX7c8E/XvWwQYtL0yj
W38yuszOLAeVMLRwVbU4pOckfCQU3WhxrzufpuMOahg/iHChrFK2Y2c6H2q/NAK0
ZsBuY2uH/bpgPTFDc7qArmmmim7vgk2V5qbSmWs5WOaXiClbLyb8WzpZfSVkxWaN
5hMBWqxE27CtAwyoCEQILDWXtbAIB6kl9Dkc/hwBeuoZJ7clvnn5+FqcqmA8xZJ7
gW6cQ7smUyC2Iz8SlxrCwDbjxBM89sa7kxSzh6SrCHlpj/tzI2B4ONLxUskg1Sas
xqTzuWT0KFLQlx7VT/QfvLizpJyYucvGlfHtAUWhdalZ3M2ofBjfX+Ii7cLOFISX
oVxpIxXruwa35uMCSAsYbIAQIN67jVVP55vEvnknSCc9ynNyA9uvsqH0G38FBjdU
3swtr9TINlUgTI/4/5LtEF+KGQspvC6qztUy8ZvxM/NjodXB3jHlL+hFkq/86kLE
RcIeR3JjP84JgFGtXKYbTpztnzECzL52W3blZY9q9kR+eFasQIFdxIPZ2dVVvlMb
Pv5iTVvSLxOPuaZZa1gfI13V9RDbyAkOkZ1oGM7w5RU+j6EFJRP0KLULI8Zwopsr
jx2BB2fVHxYqa8g8cXZmOgVpGrZ+AOrMV0SKjiMbk8PtnmA1c6/b+vht1JhkxRRE
gAQzfGeb8jNAsVanxe8dNrWcyW+zmrsh1qwAESzh07Q/JtfBfGCozx21SsTyji7L
XfuV1jIzFrSBDXz/p2S5NWliEpXiIHm0utsnMCEDK6XiQyt8xi/2XTP5aUyGYypE
ND8GBfTr5W9i9tzsoSiSVUGL6WquVMjdKu8lVdExhG55yBi0eCQOBXIsAl7tlJUf
pMrpxsXHdMjvoDoo4QTLZ7z8oxJyCDnJi9Il+eVvmFBLWgYwCKclp96rFujS0zni
2fsB/HM6ipjzO/Q/emLJx1JD/o9TpQm0V/E5WPzHrR1gqXohBGfLSQFZULryoX1T
WTFlUQJGnuAhgQB6DFa7aMZcpzW2Uff+qNjbqhh3E/X0WznR715eQzzWqqc+mcrI
CU6UTLI6EazH96fh1TU/hto+GUy/v2xlJAfhLLLUllFh3BQ0sYV1WLYd3ppwoxzu
YUiqtA6gShczkNJFsMKq9Hs5gp2DgjmJ5XAxd6Ti7xrckAioGi47AREHQPEJQniZ
BTzazeikXjkfiyu2E61RCbx+lAl8s+fSLFQ0nz236QRI0RRjIoyOh5Mt2lCewsRI
P4tgztN+xgM89b8n39ifjmA9tzm6D7FS5QUNAjCWDsRG3CSA5A1SWC8MauiZ0y7W
GMNbkQIZkZVNDkrJlPuhZOanxHWWgy8nH5VX3xst/7AgpAQqqBX1BBizYBH1QVhO
Uz3uhpcQXlauOa00rxqpSn2dP+7tz0447Q5IC+M78HALSwbyUmgrJrNIlopgq2Nz
hrYMxaqOYScfVyKkBccKRy5rWBokmte32fh0gNWKWZzdC/k4wEUgXr+vkNhID1J9
Nkf4v9DG5e/Pksq+HsGrG05KCFSY2ALnbFyAOoNEAQjzdPXTtbA9YPXN6Ag2pPLr
QevSzzxnaXgr2Sul+hAGM+T8t4jHjUxEMI0MmhVqUkoqGsJb6CuGxrZK3rnN0IME
DvSQpmf6sfX23RZcW2PkgLr0Cy7o1haXCfp9z+vFetKnxOclNr+acTC8v6wX+Z/H
6w6l+4ioCxo23unm5ItwTXwt6q1kQqaYGJY4SzCXKyV8oPJbUY4mgn3HbQjXbDBV
bydjTZ9tT4iZ3tOLq4y1dH1l4V+NG8jfn1krUY64Z7IfyQBrh291n+Oz7dxXia11
yhvAjZWraIEatYpv4WG/sPKoDvIdnWX5KYOStAa0JmaDQ0TSNb4nIpfczasbNlQ9
wWBSvevHwEntiVRvaCz3PZLhyCSgpB6yl0XewZ9zTZnEFcIn5I38U0jCl1W9GzlQ
RaOV4YMCmDtUA+oFF6/Xk2GKiOtYIx5EtQr5HrhCUrzDmsqAUtTSWW4Hjb4Zx9Yd
a5pstjudE5h9vP8LnDmiNjHWzuJS2evssZvVz6NmEBwOQ4dOhhDhr5sPUUr29Ywn
idx4O4k17OHLI2S9T0jcTiBedPqaEFVzQ/bxOBRP0Xgi2Xn/D+d6cv2YWk6OXDxQ
WR0yMBbroulc2nBf078LRD4mpH26o2r7tMKDwV2GAvf7At0PTp6lWtj0UgPDhdmP
XfwSj8f5NxEVXxtiM85iiwPm6EKlNtLQQ9vIZfydy4NsnA/tBzZ53rZ3H8aBHxSQ
kW1Y8NY89kWWyXF55ZZ8Gjo/r3kHq+JmqL4poThIQ1xmGBCuxZ2riJNfMr+ZuNim
GDuRrmshWMyNW9EMmBcTwYNFtPYZXfEDjKd15FuIljokmbUXOg3wUhHNrJSkliVp
VDyP2iswsf40Egjn5q5qPyPc8dZg3kN+Km35SgfQaLJffaHyefRq4kKXHYjFo0Yf
AzS2f4ppaROQL3sCE9+A2RH8RSjwT6YOQmjSWM/ig3x3ugetWu4aH5T7Wj+YRleZ
vIrsmIGtSmC1xYtvd6wMzPR7P5Yo0KBW/s3dSFB+yiP967cEql2S7quLRBMth8lF
xL08sgMY552UEu6t7vpDOW7RAF7IPdNm0hvKzVT0aCqmpEmBadFzWcJb87O6LkWv
PX1k0i98t37vyoQn0Hbn8Q7lwX02E7UY/OoltVBXvxde6m00VkjQ/HzeATDDGPmr
GmzK+OQXRYNNRdjzIKjPYpWBGVGLXnkUxC/xn8zcr5gv9Jfj9/GeACLA1TEwJZ40
IwZRA9L7w5bTSt3hDVYwAyEbYFNunX4Tnw+hpjz5D5DM1oLex+4PXiBPTizAVZ3H
DmN5nr5cqrBUq90KwAMffRwT07hZunkMt9NVfvdkDIZDKcI9Abv7ir9TzVfKMhvz
no27Yw+UG9dj2U+YsFFvXe+FbAHc1Uoy57QhfFgDl6ZpfxVNx/M68m++XkgqmCEL
Xrk2cHqgXVWYKRgrpf4t1z4o1KXZzhOEyw+mhAUvzgr2hmUQpyL2nqdKwBW/Xsqf
LhNzfdJSjc71ByBbJproJttEoP2hUJ/VLswU8JYnfphHGjUk6TcAMHfergEr0f7J
salf1qXhGocOcGjxRwmh3yirDR+VJY4Zsl/8vU0ogwdT9S/bQgS+FCXUlFd/yoHd
bE0Dwyduq/UyuOlKU/2rQ6tc4mEG+a2ngHn0U5rErU1Tv+boIZS+EhoKb0CCg57C
Erdjjk8/toIVjXNAsQduNnT1OkGsb2gq/wDo799DJQio6xU7CF8y89C7qjxDO7uk
AlFfxpCuGgRAvK4xJM4BAUwCipTntYKJOVKq4fWlyfIws/y/Y6yvZ/9WXj57+I6s
1YlqE7kYgH68oICrkfFTicfJ4mma0S+vps/5GUglgTUd0NWj+AeQ1rhLi1F7985Y
LDQcDNeNap3Ag5oXij69GguUL/MYHtLPFvcRUfwZuPyNI1fNMjccVU2d03FRN/hg
Wv1vjOCZ1D/x6rI+N8EytWgpul7wSbg/2kj7JXlhsWDct8JRXjD3cTNY1XJfYfzH
69R0T7CrTp0RD1QENceadm8mxh/X2R7l0oYs8kCPCxaWiWqYWGw0tjcGIcnlLEzM
UqvkDMTj/QXfaFqMkKYh9ZJ6toegc8GHUzH30Hz/GdQ61S5nk+T0v2QfcK634fPF
jHv2hSNjfDejbOYlaB335MW7JFGm2+qcxZYd7vn2NegJB/rXIVeul//CnLrGdfrV
kapXeXMI/ksdONBXgF9DqzdrbJ8cTNgkwIsYYvJSCZSpErpPmkKbMdD7HFkPUVSU
azqipC27nMRD1g6Bl/5SlqPIsLH5cl5n+4jKGrLEjLXxkG7XKa9MjZvyxvsnMPLj
xOlIJwKCau9e60nZ+GerVEQbj54rgsgqsFVKOHg/rclGmdsSf7KBKh0MEwaTjmSh
ni4h8O27ReTjz+34gIg05GPty4B0x7mxKSv5wdb/x1m8rVPoR4ww4xea66RKnuYe
lUETzB3nwGzkX0+ORCo+7lJtPNCeM7+M0D1Lci77As+CtjWkdiak3FJBbTJO7imH
g/Wqcpsw4WeTy5Yr2rU0f3zCHwz69fP63DpNtAl20VZ8Px55tomaMg0op/LrrYBn
MZsAGGsaf8OXPQMb+U3K5/uH2IKcZriqSm5sNBAq8FGpCc+btRupxl/+xY2QneuT
9//htiIThPqkgVKVKlEUSLLVBgUy+ZppR1gsGXRcAt8hnW27pmzZrtW6g5SH7a22
K1MEUbUnlwjmRJhMdczlh7YqqVgTM3iWGxm3hQU44Bk29Xj9xArXtUBlvMYyXCI8
Ujtde/0rYTrMFKW09lJjSuXKQtQ4ZHf/r9eKf2SOJ97Y9neOQbZm8XkmUEtCksFJ
mb3Ly9WhZ5IqC0/JY1T3KAJ30J+aBszgcIUmRUgAmvl+macdPHpATlS1kQDmSUqM
zF2vpE3z8kvuQ5u1JvdP3t6ioxQ72gndYf7M4WNqqmyqN+joyLJfWwZK+Sm/GBPE
ZcH/4uxWdt8jNLm+KZHEtfO76XJsNbBSdrT5Jy2GLO2O+6ih9NuxRg5jTFcJPxwm
MHHf+G9qtzehtgwPz6bXYHaaVXZHOWseUdV+f/5+AK/+rl6ON2+9FIUcjCpsuhq+
rlTui6P0E9VRuWXZZg+I6ulVZdPpfrPtCwEozivrlcqCDyIGTYD3qlK/LgByQTZr
42cwJ0G/vjBLz6FKIkOwwLh63oqJfc8Vb3XXtBD+nwib69CAKrVzH9UVjxbAG+Kg
n3ejdiUb0fDQOBC4ZAau+307iZ+EBE1THGO80lr7WTRXjwjL/t6i+dRNNF5RffKo
kmv0if3+1QrMrXAGi2V2rFB82npoHSOg+bq4+M1mC5k3HQxxfuppipE9hml7GINk
7uZSmqMK+9Wa1ak/D7AHecjdidMju/kgPj3fnwWJEUWRnCFgW19CMaMiLbpHus9h
2Blo+ekWHNEZq1Nb+lrmnFEjsNSm+atkx/SZgIPaImai09CnqAIpO3/az74DlaWP
wNjMlrUF6HU0PiUvba/eVaIBrxspjZNiX6KGO9mygG3+vZSqeySyLnGoKIzLcMxt
tGzAUiGarCXNuSg1xZwC/0FZTmlmXMttcVrEgB+JPeQADPWHCVzlsYeudF3NvfOs
X0oOc6YOkhhtgCtuoAGRXbm/ZIrzKsX6CYn/xbNuviiotemtyc2fHC5urvQRxhV7
qEpyfXoEwzTgv8BxqKpHwFu0eMs3wz8dbW9Y1PFtoUP2PCqybtXyWn8qpqwXKBdK
VNDjLpOB0jASuh5Jchy+HggedbYRUJnAD4NLadrsfx6ZPAzduxmr5J43irZEG4Pi
x+mwkAQ1AQXhgW/cO/ZKQ2eCJ+K12iRLB7DYN/W/Bf8k9fVGcGAaLeEXHA5xmJ6Z
WmbWgaPvZX56eOJKIoRHIs4wgHVt06hnzhXjl2g/mvLYmG/ZWvL5oUJ+KmM/q1Ox
EB3gby25IFQT183N4qh0bIm72zGzY99GeNHaqiSFZmQuKRKurMfLhXwv6xOrFicm
9EfmwrzihOh+q42YMULou0inyBTd3g1m/sHgKsdp0n/Dr4oZ1nwtnxny5aI0S+tG
St1htf156jv12ZZIchwwI2mWaUD/vfk2hbz+MQsvLuMcyMXKnT0LZMOiitFiEdPZ
vfpYbBS/GPl706lq+4db87DyC/JDpngStYueoqypkiA5vWrbdCRvo9p96PmnP3i9
Oqfzb+GA04Qo6sFSeOWNnCP1t8a8v+vKrCVXZxdJcTRQfflf/hoblBuLXJPWiUOI
lgoAXTfVOAtYnh7YthwVNjtIqT3zmKBjwEjgXDq/KMT63AAMxjKVmohfagig4Qpx
jiy51gedNdDXk4LL71FrUOfSvqYcMfdFuPr9uTtcJRJM0IiIQ7vZtsPLait+PSem
xEII+1OicN9RY1y1PgVrfMOaodluaTuNvyF2356mlDIrgaZTEhKBmX5dB3ECr4Zd
o8ueaQtLP/trbnB4VlAAfmX6UGfpdMrohXohuNAG0ZtVUJFIYSEq0Jb809vH5S71
H6uED8JDLqTzpeNCqfZZ9mDR/j7HYZ5h1rmrnN/9y8AbasobUqTDc0dvcYZddD5F
oMqJdFj1OoKZIgFIhjlB/oITYpFmkpE2+Fg+2FYD3EdHSY0f8sbHz07CYywDBViy
zcSm880+BhggrBmQg9oIcBf8CtuwljLAuCBpbFKfcXhOdfhdi5cHfndCJGgc9fNu
kfSCJCVkcOetLlBGZMFJLaui2TzlsxadzzgiY6qfqvwFEJvUC0pTdVqw6/8OFGNd
aE9SHSpIiDfBb9+KBM+TmliTHzlGk1rnYCdFZwHf/5hlfy3qIkjSbVRRoiE0g2IP
nAv/5dvohxcrwhpOrfBtaT6pGZn2k3EL9zVbGCJ23sROhU0awn9pETNOxiaWdNky
LCu1kIA4cVqgKCi96v1Vf75g2AMFHFP5X5xX9Ym9UCHVXWoNbl0KVC1ipNKqBkbs
8DkIK9V49faOJ8wjzysPy4o8j9HfsQ1NNL01EfvOZ5ZFeEPQAdmrSPNBXb+kaV6s
MwRpSd3Hl+12+W+szCOed4dns3D28TPNyEYelZWF5zM+w8dgqonDjNy9gALo2UGJ
qoxrpl/FmjUNPdP02QWk0PsYnC713x24Lwy3mLrBIlzg/+HSu94Jje0b+zSE6IlH
ENnV+O7rBSFuFzSbTkDaLJd9Odar2/e438q5msFCaYs+b95Qx9yLPkvb70tEVBFd
nf7BDWwE8DkeMXLqgvkLRpfdDXg7rOGhw+A0I6/n9Bza2GLFaF7w8p4hBYXZopN1
Fu0d7vfUBNVGirsQ2GKAOcErxI0sRcImw42SKYWI+POrsM1LpyLS1dYmXmbuSVdH
ndUDOh886/o2YmzjV7+GouN8ipfcjW2lJbdYhE16T0AYYYvTKY+d+T/iwTM2Wsi0
2dhDCn+Klsjjg2APiqFxRlVGtRgE1lH2tiYsK2V36bU4sAzEQnWehlCXLWX7VIGB
z3sZr9VnQSZcMqekj8Y2k3Nsm914BaJ8w5a0RHleWN5//+qv80QfvXjhAnlEZk/B
F3Y0a6bmcm641yqEDjH5aCiTdEpWBpC3ed8fhj/sC5eUmWjoq0tT3jakhWA9QKwA
LkJOwg7kp/PvKr/g4+VrATnDpR1tU42ZXUAXxQA3ZBlVYeBY5Y/+LN+xCXwNjALS
n5AWgQ+be5EGtgtq+fnHgLCcW0IdVxbh6gz1gZNLZQ8S96GWXcKuIH7c+6XLwdxC
ThCfd8C0E+YIF5kkAiMo6RGL68pT3xdNvNsPmQSwgGWZj9ZkEm3nw6nks05ypuVY
LtVwVD/lBQ8ASVZaFKj6Mh36vQzdx+Ck/aZ+pjLUHeF7o+mMLXQkVuUDRyyc/xR9
cWS9GhIdHC2MCTZZ6Ls3q/XSlhJNmGXL66XDUznrpW0jP8ULt3fq5S+G5LV85Wzl
mlv9WlNkqErb2EjRXLnOy0s4XS0SnmU+zHiW2ewAp/jUvEtyWB6yrH4bxCw4NVxe
BegpMqR/xlur3Cf0cSjthCAyLgaD7CXI088rSbCmI77VGAxy0Kg4z1/iWa1v0X5U
/r2i8tcf/9MlDC0NQShB0wc9L7q4csDhB5s5clKKPaK5a0/Gbu8xNKnh0rn6wGhB
b+mRBF+npgT2v368Q727KRUVZvmiwXxcgEf1rOwtPY1AYK3kuQtB/xbm07VSLiZ2
ItGg8WIrlwDq60M2+CRpfrlEakxcfQlKKtgUPxUSaO9F1rV5pj38tDBfxCFp7jYB
Yq4ytiqb3zNCPo0yOVsa+1igJhHot8H99eMnwkineN9Lh/abMPyKaGmNwOJLzaDd
/LBPMQPDfltVQsNS5n5HAxbzCeNSTGp92xs4C+UAjz2N2M+XwP6q8+rbwR6HDJcI
MrPpPBuS8KufD67A4cAQFYfm9H6CRsbiVZRuj+hkxsz2LxvZCLBBiW28PgPrlIlv
80gHCrKqL/N9FjT4AVS+i8MXO1WbzPnOI0nJJmB0DXA1gjgMK8kH+5HlONW2Mowz
cdA0YJiLX2i6C5hoQVda0TOLs+XwUtG6N80RdwjTxUqvztH4f+o2xkyeoCN4GBkW
85M0E3CzXqL9AACqTmWVuHO5RvKOXaLRYxwxPYp1u3Cv+dVRSSAIBzP4swhxwDFH
sE2mLZ/7wFeNMPa79JCapdvJMt2fhhHovFtJgguqwnOub7DzbK/b2O4uFATfe4qO
pPSVLeBMopjeersIk4Ny3gSKEpCgvaTomIT5ThEft6af7drPS45MKvmFeGrgshoc
WNkgqmBiNbzng2IE63YhR2PB5FZ4oDbNkB1k6Pmd/Cej1HXdUe4uGNkLeSXG0Fgq
j+cJSrg+wMbve+n80Lvnzr4QOfoIIILts6Gq3ugVM9CxQ+Bw4wBYYdGbDVww/XI+
AuZq8gl4js8hXE3d+Lf4yE+m/cEOw5OKkgF4p0m/w0ld0ofXN04U/nPqf/vLCe3W
0x7tiYE/XsY+r63hD0L8MfDEy5vgm4NKPdCR/q3Y+fXze4VnG1vD3LLoGUQLFkTC
KKqvL874OVDu8biJI4hrMGeLjQ309Gfe5iNN5gVxAADKuIndMghamHhoXLDBA/I8
6+yHfOtft3jpl0Eg1yR5fpvtHlpMbyk4BiTHdkCYIG6eM+H/eWAm8kISme4Vpw8k
rVHa5HilOWbv7T+otKvmVH7Eel4x0mNpZ1qLHoWcD+HxS3QaRqPbqL/C5hYFmPA0
6KYnPI4fewxZRh6CzYH2Bq2DHKk1HIlr4vL1RUi35loojhQUm6lFfBeY4vvXGeWi
BZVsBMwFECGmgH/DLHrL9b4ZsFqWv8z+Rhi1o3nhfJ5LznBE6ijYNXTn6nkbd+jz
Qd+BmT+jauFyzKmIls9o/975wB8xuFqzm/+vw5t1wdziAsCKCCONMQQcQBdwMlAO
EQBJ6c2a+iP2Rdm5Ww9uWRGClE5QOm8vkZVP/xJ4H8/OqAJbQclVvBNOaDqWDMtQ
OKjLH7zrEVQRRd0hqqPQYJ6uuqt6m4I0LjP9WTrGLDqLDHwgzEQ8dOOBeEl6P0ra
Leac3ugSDQBytr8g9gqrBHfbKv905QRNQbqbAidNIIy1aGSGTkoBlkfKFeyweTpo
KvIQLmqU0eucu9JfhSCdTXEhA/1iXcK+cTF6PxxeqmsyN4kGfwub/PpqwWO/p557
pcsPrQoNDY3UbI0zxkG0wA6NDXBDeraQ/qeuE97eFbU10uea3pz82RY26a5HE50f
4hAH3ynOREjj3rCZGKfLwRLJhBuEu/tODHCYl+Np0yoO7ALra2uiVGKa/TmoavU9
fD/4PUzMq4UvMJtUNB5yikt94izqvXix6+M6n354iZQYX0SCecW+1wqVOO8MvXGd
n7cV3K0hAl724g78TCcmyOJmINCU6rMFjviLT0Cfa8udk9sUd6qM5XU2ZfQnQx6w
ttNTTWrYxAFc+DYoqNegbg/OnybWuhbb5vTW+LLhixDjAoX/B4G5CeI7P4CmsGno
U8yoVBoGNAakoSFeLTPM05rXQV3B8YinGIiNRsKQ30cOYw2xDhtnG2VSmZEfynvi
bpIUq/oBD5VKtfwZ6sh1vcBP9ZccqNaRqmSzNmH6YfUfoXhPasUAt1KTkqGleD5Q
OmeD8fRpglrclz3wVNf1GPBAR54vVTkrOV3F7DhSlh0CJ+72SI4EKPEic9Ffm28M
AB3oLuj7WiQL4nz5wXptVseLWTAfOtvKZ7PD+U86ggk1SoBz2XxiRCtTRrlyQdhW
6U3rIzM3eUEVeipqZfaL0JXbkKoAVpow3v3AYJsVN1dUSP+HcnJAxf6KDEjcxmC1
l3pLsz87hD/4jWFu3Jb9PWDGK/JbbOLrqz5aaSUqhqDfusgfIQ7kx+Z9+5F28rar
bmQ/vW/h0eS+q+LG7Eof8OieXeHsBT1j8v+R9AeTlVw2xZc+EUYI2E4+seA2kBEq
lVjpSO38GGY4TmrQN8SIsq5zcKxbf5jqtYdUYm167EWimGVHkGYlg03tECEzXECH
ifc+S/VBbykSccHc/bhUt6qMawS+murmozD4gKFEk1zqxvu94VEFUnWaLaXI1XHt
BYopmge/ltP8PI88KrSFyMfBRPJ6Q//z1N1XcP449n93CgGnnHRKuZ0VdLlMVl7a
lTqp9Oc623xOcaEcI1QqZeoJtH0VNyYWI/7QDl56/jNM4UJDoRv2EfqfdD9dFxaH
LYYzbTHon/SMH52TXz7VgiTge8kE09GZCXWQsJkMrzgcXnlb5Rqn241B0pjXElP+
xmW2PcQ39eD4v6QZVGx6QCNJXoN0CiqSnfl4gJjmQ4r2NA7uvLgt6M06kPipxU5t
y8OVWczJVXxarD0i1BJLYyG2S3/4MpY/Sr43A4cMbbCIH94lyhGSO0dDfsQ6132r
MD+XLHKpjKuX5EDHF7HlUkzW71q2bAmAfRcv/TAbThAVCNf2SfxXEbvdhlp8lK76
i1SekEK43HuJd+vOIizQ+bC+EMxXSewVkNhHYrU8e8KI6yaSeCDM/DgPafBb4zBM
46RLVo9XJf4YKRUJYIEBXR/6eOI9Bn4F/nL8sdiElkTPohzerDS20zglJf5GiXhw
hVMw07YEFwUM/ZtMNkN2On/ANTPufuAIzyJhqFskTUqge2e+1DtL4C20g1vyGzBm
q6Uztv1sQXirJ2nZsYp86XbGy+aUEBSr9dnNqY2lTMrVJrjI/IiuI2Ux1Dkou84P
dY0uapxK2mkkdWdGkfxga2x00a78HOazvdKoMaPeGfrEApxNuadggWEnPIWI57n1
J8O35QqMKDt2u6PU8PEDR4r/d4fJc/9kocJJrE1UydFWKD0YOOo6BFgZbK7Zml6o
vdg+sQEyxLY+oVDXZFO9gemExou+/5B7ynz/BSJZGlbgKf3KIcwhbyAAPBNqOgpu
Xza/zXUtfry9vnLpV45Xu3VHJpBoqfxsgS0mzjLnx2b6DKScCXgdztbhU496+I9S
/ysFPpNfjubeFHXWeCjrFYEKA6ufXAYBl8UybCkW8D9dvPKPrsNYVZ3VFkzyu+Yn
iJkjNEzNKEuKYbrkMrvwRYXI68x/ycwwzKbEcW5WvLS4LP9FgNRyWbbvEytbuzuc
XjxWexU6EPYzLodKz8TS7xnx+ANTBZnhsNsS60HPXBdSw/uqeQN7FZPwkyuiivml
C9rEe/+OFO4Y3pJBkk6CMPErgFqBH3a480H9Iouu4yTsKQXiPC3SvYd5/XZIuoyk
LJqwzatp+pup9U8bZTc5OUwq1XrReCkz6RUFWmyKexPjQIQG+2j+OQzDZrnzBzvv
1LpR+W/uUvBbam5azd3NKtxL41KKprcQ3N/SisV4rx5v2c2zpzXgmv7fHlTk2EH3
MxFmx0+yRSYZUc8SxqhHcuFHIerHUWwgbhhG8v2zFvB94jNcoLmI2gebaYW1l4ua
tV+feKBYnYkGs5Fvg8kJWBwwH5xS7GmsO/7EaAvuZP8WYQoQLs5+4f3DrMDsx5T0
lQ3+OL1EktQBaJIj1G392mv/IuH7GNtw4dfVGUF/qHejELsT/W2By7GFkgkr4nUW
PxyT435olOoaHK7sS6CbZjeMJL/pmbkr4MQRE8q2hcTtFYC636qXXb2AUIanKq1s
ZPhOl5hfFvnGEAbDDET5T/PLf+QYULJXI+4FbqErIqXq/HiqGb5EKG4V/oShAjvZ
ZhzMHxWRuRVJ6CVOgbKWafkR6CFS8JOkSBPnjJqgWt6nOoqIt44NTJXnRcg7rFsI
o54Lp7ZXdJ24zsUIXSKAUzNXheowCiCcFQPxwtlqJ/iac6wJAGKyy3PtRG/5gdSs
3H8r5Gn3CVi+5ilu/fkcTlRk8ENNNfAgFky4Y0GUT7irtKwoexctYGkw3Oux8sNx
RRtN2ms+x+V/8PwTm0YWReA8zcvQ3ATHJNLbNh9MHypbpasdWwEOBNaIhffsepWi
bN/x7K8y0QRy8/Qke0Dooawd8ixcjdbpVcROMBCDLsa8CuumMgVwYAN9GZpwYLkd
V/Io1NKrIe6PGe6i+pjiTgStKysJDREAoyyxY0p6RtUqKEPrxFZIrdpHj/7iXCwp
RYNO2VCSoGjjS9JdLsN2VWrGZMnhK53LteogQhRvDjrudH518S9+YoHCqIGKM+dN
nnqMzyuAczZ1cGKcI+8RojvN1p27rFVRBuv+7zbl1dtqSdqMv2KBtDjN2Celmcj3
QcLtz7aqjvvGDUwt41uYym7GQxV2CSkKIFr4nAfdYKtiCBB/avoMKaBZB8yjhD0W
Qv2KmFo4cVNQ4v5dA8Lm4jksOwhtlnQKi6uiguF4BHsu2TnIiaaw413BiTEBOfCA
kRCM7hGhXu+AI0VBjGMjx/v5Ewc3XnEPQOZILJlWI7fJxEyEs2p8SVjrSSJQOBw8
Unuhgo92w0BZ3H2ssWAbicoakmc8L4G9lb36D5axtD3/IlJJwIRHpWUcYCbViSL0
RKGwsWp7iv7o95Vvck56urZz+xl4WYvoxr/0N3z7KxenDYgYwdXfcRyj0+Gw73N3
3Z7byPGIKWqEGW60096GgEJKQHFr8iCCCQtcDgLphY1IrcLMilbmP5/PckGr83oc
1pUZpmHBVnCaeVPMLNLWfVHsdygNpu2DTlZuRaQojNBNSjWDPTGE9QAjtfAbOelM
5IIvjDeQFVPrnHivaMy1rTbKAjeK6Vm1+lkVn1sZT39+mP8zZh8sy8sumq9AlKaQ
tr9/INVGlso1a6mwYd5O/QgAmJoAsoQW+Gb6QmPxDhG6HCYfDhgP7dkCiKczepec
TpjjKkd3SmYF+ekw19JpAD0u3ORffDnymBA9/qohVNb3cjTnFBrWvh3vhk1DIYuq
cQLivvHixKJf2VTcJ4tZ9SAqutmI12Ks1X7jgOCowV/U+inxgPSLkrOVogvhSEwZ
IlYcyLVSmy4YHT66B/B0mXZluvrgdMWpHropC3hsPhJBZ9lFWvucKsWPaObtYU7A
D1QAannXySulXxyWYP/IITza+guUxCVFHrFNQ4EPsf6TLOVfMzEG8iXq55hkQ+w/
5MWN5HW1QnWkPHTwFaXAdL8y1csQ9xp/71NC9byatTBIsfmwbad5Oi8yB5EDzixb
tEzdTWfLw+yWSuhWaW04gCLpwwlRPVXyZvOGH7ktN4OmSdSpPoTtKbYT8Xf8qjo9
CiAIiZru4J61pHEzWJSD8Vika1li2AYuH1K1J47EGdsqYuiwaGmipljglduz9tkq
a1DSBD5USTYvD5JxGa5tLPKhqVcVfBF7X3vfv/vr5GqAgUB3x1yurPwhXVk8jb0x
d4VZWUlAJ+WbTAHz1ox+u5O3V2g8/RkQcd/hgYGGrr1qrv4e1144Z9pulPZjld2I
Fu6ixDMCsG/2rFV2DKsa2j7R5K/ZnvNLdsjwfrBzYPsjrFBvw32swNDLeCVjgu/T
2nU7Tg6uxm0eQqvsYwMKwZ0aKzpxbO9HOwInVsSm8Nrr1qhchxGne/PxXiXMH0BS
dpE1P45FiOc8kLYhhDBrFQcp8Fq5xjbkiFd7ksa28sYdd5u7Zm4Xh8Ax8bdoo8cI
vrubKIXGnJpKzvW0xCCJL6wPkpQnNyg24wmwPNRTBxmrgLYuHdbJdQOMVIbNJM7v
eOHtNb7H0L1a0ZUmFRJMdiUuXuG9UIK++w4W7KOx3DMrK/Ahu21lFi1tV36Y5F1q
U1U1gF4fIewt0Zykegj2y/YW5d/YpRRLIaA2Ffdd4DLKaE+bRfwMmtwjCM5UNH+Y
Oqduu6yQC+gLbYM21SUi1DfZBjuJ3df0vajpZj2fdhgzDF+PuYBxWiJ/67zUs9iv
+BFDAtfQElkH2XFVh08RseNFGo5hbsyuE7d6yDNWzjArKuHbeKyyrYcOZP/DNC0S
QCoQGpv/L1KtwZbDEtfRNXsp+n+wUqu9TtuX2zVeuRTR+OtJNI7MMHeBz+1NoDPH
goEQyuVW4h4hx1RNZWSqInGvvbcUJ0M6MWjII3L2NGIGlqjZZVlYE3b8TOLsGoCN
K8/Ej3BdrJrKF2M9Htf49ROab7YV6L8ibStb4GcL1HP4RgUB2RAJ3X51Bmz8gVSo
JfW0NUeOud4CeLMV3Is7y+x7Qx9Am5Fmqu/B14Zrt24K0HVODp2Xebz+W6vsxF0P
M15izYkiIRxH6AjjSqGCrBWTfkrNUjqQ3qjZNHYrILgHHPkT9w3/ynvCDFLphWJ/
8B5Bkggt5ehYPCNBNA4bpVg6NiJEUoR3I9k1WtR5fRUrJjimgHO/5BSfYrWRsTr5
6fk8tSHZss5Lvct9D30idMvQriK90huJdFKHetJyNftCOkEweOhcrfbcLX+vLCgR
JKxjXwXkuXO32PY09ZxP29nncunc8dO9UaMs8LNk91kKJLetZrAK5AKqVsvt3RIW
+RYWnMG+Eh7uU5E7Lge5CgVkdtDcxh/2IbjX29EYwk5fcwYYT1PyaYr9xz43jTec
w0ZUYA0avKMszmbJggkV1/g9TOXJXfXcv9n+GuH5gxj85kCvzwoibpnTI8wHjGaK
YNzo45zCGigMJlytqmchZu+aGYpQBzeJkLi4JmIVo0pVq72CXIDkVlPAyZRy2RRh
UA/bXSgcLcFNSUzvGQbDR2QDO2NN9lbC4330U74p2HhUzRHuRXNqqAQh0Pyc0KYI
RMRX0NRLuqaCQbaVHNcf5zM9CZgNcaGhI0b1ZAod9CL30R5puPlGmJIwk7SMT87I
j5PWx1yusP5KC5AnzpfwfX2ep81u2krsPnBoj5QE8Sfias0Mo0ax6VN8DXy4To8o
ArAUW/Ue+0c5VO8XvCjyN6UK0Wi12VwLK4715WLq1a2H7eDp0m+on5ru2eIZ8Z1V
ZOGoJAbp5NulhteOMNO/twQRlak2G0CiW+/SgxYmsP8hsKKGfk6fsGYiziDAdwWq
TG8MQjmXhNMtFiTclCnK80YaRCLNT8IEQsa8h5jNmxaunuPPgtINSOLX6S5x6OdS
iRPhUgpv14gASvuW2VLl4gB+qdHIISUCTJNxjitHpzOs4kx0vqUXaGj9yMc1Vt53
tqguOTpmcItVJp9VU01T43C7dtgyXclV00lcQWDxVp5vCSUmEFvlCUBcZdHYtVts
4mCuVO3a2sM0K58Akry1YehvKw9cvvB4BRNHP6gJsI8bkhLKPYApS+obu3v1p3in
5qjNwjnI8C7hwERfept/Oua/XDho4akwoDcZt25/tYIIcMSUzU1EnojxO3+Y1lvi
75bl+KaF6rUy7HYePN6tGdn3SPVL8hoQA0IpYOlUVNs5Kfad0n1w2HI78oE/LZh7
in9L1GPkd7wtLyVkpsexqqQYXLFUeiaLcyyqv3HXNaYKe54YaW5Ks4NQkNZQRFNL
xSPIiDQ8nKy/YIZO45gaKgtMTJyIOvAoIRX++44Q7CLdWbAgbEYGkowZdK4rEOw2
XmFTJ3FwEp418/G996dgo+UJk0/M9egIoTaud1khonn/oWEHFa6/AfE1YTyX9rcB
EgB4lMXe/ptjwNgbqRHSQK7Lv8kRvDkIz5oA3DLWUMnXs8pd49Qb5J7LG3OWAWWz
EDUB9/18Hom1Q6IW8IN1szJQux84SA7390ukmrHnBVJ8iRDowXG3jy6jzMYBlemq
TZabNpSe6HF6VBTJHNdJ+iCbd6xjXlkO26AccJCsKymv2Z9K3zqxCt9RG4LXsTkG
tbTCCGzKL6rlcKC5OYZxlb2IHzS9NEfifCLW9i77fWjeUsRkQ71IPRYN8FIwQog6
38Io0zxVZs6ZawTdR1M19SJYu8U/GYnEWebsc59tE8ffjU5xnufarZGUxP/Q43ra
PIC88J7UmayyDfkTwyggASw+Jy7ejJ4Dba3TTKNpmZKuw3wpxvvpyYsGTKgvtmFY
JSHLTEpPPQRU2dktIOdn/588L1shcDod05tcmk7q+z18RPuJd95oblvuJ3UNo0kE
lJXpQPHByhxn1mjgAMVIdHJ1OHrBW7MZiX31XcqDiEY8hltysJn9HkvIa8mpG6+m
TutDh9vI6Q8SNV1FZpjNEwIa7geoJzgKOxhtVBU/R9uehPUd9mT4uVcpdHReHdpB
yQLgEjdnd+Mi2ToOXa4z/ZjUjeorl1E9bXtGpdKb1S+WpyKigUQzaXAPCI3ynCou
7HE+dQ0S8EVI7NlmYiSDlywZjLJHROsGPXSSwRFlXB9C+WrlpTNGXHp3KbJ+nZW+
T+fyp68u0ou1udHfHFkybxnwlO4H0o76isSrUtg3Wi7LO6KMM+yM2JB4Ebz1Lpq3
O/k67HJv4UTi+Kh7fOZZXgHEfYhnvTMffX+M4R9jlAEX686i4I/1ystfGo2F4PB+
jYKPxzLP7WdaO/WhZZEFcdLIuIcr/dkeetrhK2lb2W4/4OO1Ka2QQT1kOyFTH+75
R1CNC8TXz2HOwD/qtqB1wSe3JFMeXa3mQjcp0XbuzxgSMef9rSplfktd1UQ9oW0o
nU2sPFnIeCEXvrR9inRleltAdVchgMUVh5alNdl6kNjl0+BpWL+xTEpL00p4m5mN
jFPCTgjmTDFhw98E4vE7x1q9FLAECfsP/+Ep03oMTHG7Ay1Bys5C48Sb4CSv0zf6
MdE5eID32u3DCZztklZbBdxidnEhFg2mvRApxvI7LazTuXELPOpuZUuWmLg35crb
84RLlb2+kXr9URIq9YjdWtOSiGVAaHtB4dymNLkUaUC9TS/OloAu4wuvyJdImsAc
0x+pccQveKQqSI+9zliMQ6tJbxhQBku9IRXgQumBD3x8COEC77mbwSaEudCKSi74
ZMMhCYBJaD7MqSnE+qXI5G3kbOWrIt8XjVWjUX5g5DkP+FYMRdKSQ8Voi95dpMn6
n3N7aqiY5ewvhipVa+MUj1gvx4VPRtlAnILjryKDjMT05pE58w5yZEcjfnSpGxsU
Xl9x3iLTSyLMNbTB27S2fWAGAOiKs7V4il+m+TdAvxODSTQye6S374K/IXx/PWeg
vbU0OeWzDAd2GygQHi1qssx1gLbQs/t4NLAzTmz4j/FxrRvaEpf2qmZGLlo9qq00
d0NwTdfOUubyWjiK2Ac637KYs/4cYdnf+uwkeZHxAvdtQ8nfv9wUOQoczJ1kRWh2
bTap6QMA4Gm/pU+iEgDueTn7iUBh1hO87T5fgGptGcD187SluWEjXrGPvTobtLYM
jm1YUJ9ysKwZ8ot47ul9ENlaTX5h91C+vEZpMKly4PcTp6MCQHcaLLdFPXac98sj
6x7d56i/OtmYdmBkoGwiDuXsuAn5ySU097sr5MGEEuNYwuRXiTNhPk/Yyhplp11S
DR4P2nih4ScCsiPTX1bKMp0Htx9EWDO81PysH3GImTxJLV5ftbSNGis4Z9nbppqy
B2VP7d2Ytr6rbrDVYVPcNnckI6DEiqXSvumKq0dtN4wQ39JtaXZtEyKNSWPgjFya
pXa8uxZ7+eUf1ddp79kRzk7xnCOs+U4USSvJ9nRvZJS+9E9Pxv9ehu5qti87RFQ8
AonuTxSeiYL4QiikJQpD5EdfBqojPMVd8oMVg4VVA710s+4GU9a1k+8XS2M1kmwK
Mcr5G9uQ/jrvYc7+ZO7Fl38Qc3bQvdhrwb5Viqc26gyM4DsT+rh8Vkt5t4IdSgHF
Q1nXFEbZsb1qmhif+JMNMx1URyOIRZawVEugSWU+z+mZWykYNcmJc9ESDzu8Mtdx
nfIyKsdTjYS6Pyf2ykd1MLMiHuGtdaR8Cf1+ME3Td+I0X2HOG3GMnsDJa5UXUeqy
0oboG2hAGN6RXiw9EW9xqDy8o+RnsmQLpzVmTdoluHXy7N7sPWIlTppESU1BNM++
xRZAXgpY/oBSfL2dYarEJLfASihqMoU506R+XjudK1QkIrnG8HurNPKJUeusmwks
JU0y5A4ioyT8BvRJJ6MvBa5kwaYfdwqy9taV4kbglHfNyyLzoJdTpBU6j2+UVBQc
MBzL24/aV44fjlJATc1VaaL6k17dUZPcFbwXtgR03nELt3ZN9QRLNIz79PUXKDLh
DIRZKqF/XfnhOaynjGQjPkbgZ1E5HWhRDRR92H2F+Sl7e7HW01Lc95RO7nGEsLsl
jXEoE4/FYse3gf9DOKs7+vq7EWRdKNTD4AfACvynehtGXLBBZcfXgtRyFQP5XmaN
O7UWlKCkZuPVllRteNXHWBE9dG+sO6j9PsmkGj9pRSz6Mq/dQp4ZwRguGIF4A6vf
HklPVd+vXOXANAbVfnMz+IChusbqPIe0mUwA+Hbkp0ue89fbtkxtfhbQpww/cv6y
PRfEPUysZJhJMivYPtZaU8hJnwsOuFURAC2miqp1468dLsk8gixUOuyAirjCk4O+
tS1F8QnQpITGRPWUQ5KrmW71MjlHgCq+sQ16Y2q6bOEDHpo+i6OLJr6a+yNFiMjR
ZpMWEtTsL/FYf1Lf/4veTXCvkXW0GxFzjCIh9C4VFhpHUyvQSJs6t9OxR1ijiQ0q
fP4Ilq9c1+K0S4p8EHo+oozMjnr2lNMr0QIViIVWJhR/BWW3qcQ4ksrRgLuqUuam
9hCvivqGFQYjuAtQnO9fiPhZ/w30N0M/gUoJfi8xMeVd98Q0KYRd5UgJuNCWcQYy
L06ubArZuxGerIyLGrORuR5heduERk6fBkBz/a7sI2jr7use9mhu122OvkwM2z4D
Z1equeI9hkN52x0To+Kd4xJOqx05zSBm/sil7gUKUVSD0KlBqnFrgUT1TsZSnVRw
kfkPiTpUojv6ZyC1pvipPKjLV6bGmMEA2f/9G0EWJX94kW0BO6Bceeiu1jXZbfK4
EGRsxBWGmcQlaHFCGvgzXX1aYzVFjx0F3xc7Hx/7Y+MH7sAtzpRprHMM67qB0es+
by62/BcNuxHAyi6tMYH8QtkBZuh/qDNegyy2TguVmlXf+D6iTcIV5qI8uF1gIaSc
m8LUv0CdqmOplmgQnEutRULV0zzxzuvpsNz56kgs2NXn07viTu3SufhgbGU/34+p
sBdjiQsjUXKgOwoTcelZF55TTvJXwQgxDlxI5fqKW6PX/bVur7KMAKnLSPrHo0Z0
IFlHmfsAdiQ6iq28bXHY4g01Xpk/NOVXN3T3iT7rQ+RjGbOp7p6Qf8Ah+rN0QAxj
KhyT0j4CHCp2zYULSnbXe4w0nxOlwSk2iE3TVorK2jmC219L3xhC7E2Er+bvnFgr
1L92w42DJCM57LDa12mcW6M2CigJl1DZrmP+nYSRd0NdCm6vn78RMXdFOyhn2EfR
kuQCExxwNTFmA09pacSE1K+XmzbnZeKgE25zl6ry34udN6D+mXeoZCBMZU/AWE6d
zUOUPWPe1gdWjcUXxnPBKkDvVBsF3jBEh+Y66rzs3XN856EQd2mIbDQ9KSYIe53T
akQkOBdKcUsCka0AihhCJwaCS3O/Y6CCkL2+YS+PH7owbwGUXpfPjnc898VgeRMg
ZEDRPbIoeLWnSokk+uf542DEv6M1V8EdHEziTOhnHw1HoTh+cJbPUjib5Xb2M5aW
bPQTG4Sn3D0zPUg2hw46Qh5BDgmAzT6YghWkzYQxqk0MvQiCqlzM6cWkqHc/8uEZ
xI2w3CK7c3BWVAC41BOuaGfdh79+Wvy0b15Vc8xIBocoWKECRgqWSS3flGNdrBtE
/I70Vg94aRN/qJTwvvXHDXdPtrKutf+pe8i+gO17zCgrEyLUTr+Kjygl/4g1dg/C
iwy7081S/mgM84wVKJjPuIoW6cjN26bjM7SVMgg8ErYs4+cYME/A3uLt0k+LJsNo
sT/ynAxfjZO6j42QkVWdc44YLf3kVOfReBB3R0pR0BY621jCQMCUVtIeGkgdEeKQ
/3Rsl9Oc+nHVh2YyEQlsxO4ZVD+k0wpk/5LOhbupscDCJEdKs1H/Bum6WEfp7eMj
teJRa6bUNIyRSykr3iLga4dmarAOH1+kNW0jcZLW1u8Vyybvgny7dffJkds4Dl+l
w3+1ZhLP2E+QvMwjSDxmL0R0/Nf+uYyZJc0dHgartGPbP45A/2QhVgFJuh9ucsg5
sh4SPfDSq7G9iEiOiCvuTwjaR1P6pfYp+QxQZJuS8ui8glAHpPINUaZeiz8FHUxG
yeB2z51m9B13Bbh3RWtLequBJ+nFUlfCODyX0r8BSP7mMElpkSlpBBAUozVEqMUl
WqjYlBMTEjEMArB+3jpRGNWiAkRNfeZ/NrQ1ifK44DYTpv2mEeHa9QXp6drKZTPB
ZdQa4vrRcSQ5J6AfeiXky3Kyd7G1OXI0d9DZcNojRttjQwo2H0f5StObwzIGjzVI
K0YTNvz/07aAQS8P6/ja+NzOmsAaFIwvD5qvVjUqTGxyEJoU9t+wgYEULPhM+SPD
QDRvSzZUa/DF4Uq9hZHuZUzKWPiaimfmsbVr/RXnmGxFxEPDbpiK305Ax2lYvhbb
4On7Ex0OJA3Cn6HFx8+gj+mGBRpg1E9uKupPXKobbrNSksvFnA8xMM4a4C7kRUZE
Ghgyw+X3IEw1KGsg00kZX38hqzOOYQnNSt58dhcFMJltr6U/ydL3PMYe0M88OcOB
sc/L2Tm38uwYO28TVP9YzrtnXphxd0YCmemA/Bk14nJKjLUS8Qx3RtxRemQGQLlZ
/VFcYQ3QmTUBDxFWWkD4OIOBzIlQwHXA/8/OvidZazRxFrHe0jF62iJAJKaPBj0i
CLei1NTswmdbT0jAYZNi9OanUlt4DqK9JuGRGhvkK4RjVTW4F9n2YYYr0x9MF6bq
cGcTS3rNOhNfGysYa+ckMIRFBAjvWuhBzeRENO4H0e6W8JNl/I0dqg9n9RFcgWPm
KzbNHqNOPYFfLRsngeChTh/pJbuetxNcDcTTnYxJUFvZYX/djBEx+v+fxjoM7C7T
3mZ0V9chcmknpKeiVzDhgFR6pjdg2yvnvToeT270sw+cnfgliFMTGm87sD4mCfGc
3bKv1sfRNzn6K2pyBQktAkLzKnlqSppHuETj3cY9UWBzQ0C30rw1lWRiZsUYw26U
nkU18+qX4EG9KqpjbN6HwBsMwiJojgVvbO5sgKLCQ2NJ90eb3zPsGObIKU9xhk1o
iLME+daa8dpTeozYrBYaAFh2GrzoV9E47+wHdPRzC2Ha9p340KlXup53P3wfKWMy
e0LaIz5kbLLwvqEXV1isMh3vawj1fV9QZM30orox/lpIdPduFwRhqMZk9wMj80jL
ucJUbCYpxe/8e87S5yVmdL7xLWf30YiYmpT9wzBpwk6GvcsetheRpGUetziqAnqH
uzslmWKZjymBjB0gxBvO4m6eWjH20ez6ZuZ/f8WyidojMzq1SoKrtrSDu69iOQp7
ip3mksupagWJinHFnhoj/aKrNjqitSzP2PnR5GH5oj2ELRwvFMSiGU4BIyXiN3HP
0l5PKwxO+QKYsFUZvzBlRrN3eaBW7ZKv4J6SMJohMwFrUBBGNFetnVG21eNPfIHi
LXB5GFBLUK8TQvjXAen0/4cpMZB17b7erYb5gDHnu5AbAHXL9xeZy6W1jcFK1zfH
eLfoY1/u/8eLif8if61PAGMArkxumdkZg4oVntKhDN/K/CslH/Qt4GcfM+m5ulir
tU5mcuhL/gpcOXYlbN78g1kURRvt2gw6/CaozsZHTikIN1oU0q57WWVzTXg7B/53
QptpYh+ldt0oc5tFW5Rv99/irE5jfZqV42jWIx/Q2xxx9GMBnQUOu9W+vHqHG7W/
7AY7Mu7oME845y82XJuCBCX8gZxZRTcDJmiAOIu+VT1cfMOUuM2Rkz+Mwz2qp8YB
kTlcvhpuHx2eX9X5g+BSJQBqjkRhD6uVWDYdmDDHkB1iT9b0qdPzCp8cxqHBFn1q
kl2+FO880V9t2S6oc+74w3XRPv3BPeJLUrtggMF5mGpGf49stOOMo6A04p/Zzbq9
NMKe8Azk4CU45oGZ9uhj5E6Tkpf42u+bqaM/JTR/8DrKSyuQMdHFVhbbEp6sCvvn
r3D0+Xfs82HQqCzSFdfGt1kn107EZg/hk1lLEyHeHHpTZvd8+l/EkT8F3pWIgmVd
GSRgYtlGRnfO7nIWF5Bho27DqyC9YyZ3LlbBgfxlKXYF6NBh+ma+0RADrvRSIG1Z
Q6VaXhzO/EBmAJus6UN8wECxZOaOS+ZctH0sOd07J+xSskkF1QK0//zm2dO1EQpD
MNC4e19yNeIydJiBx1IPtE0H5jKRcfl2LJpjdNwqZorMSfMiEAfEPhwUTKTbuX6d
zZ9QK05oaO3AReOibcKnBhPfiZsBClsbgOE1QpHPGFVA7h5jE2sg5MkxTwMa7I+z
XhWFjKk/KW9S9wgaCS/u09h07ijDV+xRReqF6MNGtkrC5aoEwFH/LrNAuSrK2m43
V8791x+H93uGh2a+Fb1Vrxk1vhbckwjRgWvkH/xdFghHKQERbo46eBZGqJtMLThX
UHX0UikabEF/DOBSNCvNZM4OJg0ik/bfIhPYjP5MevgpjiveYHQlhiDybvvq3kae
8+UnFdxuu6n5aAKFZl+sud7NdhRMSiAOi/RUNqpREcmwoN7Pv3iWMt2t9GT66zdZ
tG8WmKR08HXczDsGNlkzFh5BE6uXYmWnHAuaSRP/l8J3fDrisoJpNWXr5VRA9d6U
4vt8G/jKiB7IONYRpdBWU/oR9TcXJ9B1e3rba/h6gSNQXpuFcArLJcoAVYOWc5oi
/pOOmU8gw6Ig52m6j6PWs42K7WQbwX2v7btsd15fhpyhlUQfV1i5S8A0F2mK+H6u
dWCrLLTf/IgwrF4jfiUWCjbmGWk0au3H+MlcRq8J6IqH2k/PEcBiZBleB3g1U9ly
L5fEli0jj+Ll3aO0trbinc64Vd9UVOtcEi71QLtoT2CzaNRZEG02ri/i7O6mxe3F
LV59a0ipMonw+PDHd6S0+Dhag9FQW7zU7HGmthtyf2htlvHUxCDUxhDapxW+U3/+
ZmgaKL8zUVmHy0nS+OD83XZhpUik8yNpksVknM6yFs7n4HSFL7qqWoIWLNgRDg6P
h8eoj3KLmSku9mYMJ9zajJTwaz9VkT/EqsgziOuyuh+LSdr3aBIXsEQo2TG1L2tj
Q6moTOnydA+2QVgRMzSLFfNWnkEFcX0cEJ+sBJ5HChSIrUd6wCL3/Tq8Y7GUkDza
GFjUOFErw9gOOc/m5Mq3MWF/mTvbf50cP7VCzNWdvxek/1X7Rrq8qCPFuMfsLIiK
9JBZMe4ZsF/Q1KEAhCUGj/Prv7mJlmb2A8paiExMbSyIVKnbI1KIvBodHyTpqDB5
m/o2LkIMWYkbF3hM2cvIO4oLbnP9lP6HHTvDK9xmwhWayGrsHbZsrCry70jAT/iX
s2OAoFuSNdvEHkDX4GOExkF3fJUmT/vOSnXM9O+AIoovve40B6yuzsC3rQ/S+ry7
qpLMmSKpljRad/Aa2gr7nSfZfvn/xAThfoLuLXkNEiqcLZ5DIKWjX4SYKipKXauI
d2Pgv2oaAw1DVaAIkbnZyDKbf4uPohDM6Mgngrt4KyJdyQpospM5HjFSLUVLKwfW
gsT/DtXUF2a6uRtQUpHQLQQBANmMV9wvIYZe1L4j2cQY/Nk9GNzNOxMN/wxqnOdn
tcEF7+KixmwI4NyucflipVrq+aQFEvHqiGoaUqs37g/ZwLhHGZEDtcWA1/mrVy7O
8nMqz6O15jzFrD1Wh6c8KSWPFVKi6cLMlYA2u4bX1FUFgaozyVtvBynKgR/Ue0DD
D3TDg8MMP9l5gUsYMOG8K1i0BytLhaR9ksK/kWCL/HdDEpne+9s8OKfaLh1DszSz
ekzpn8GkLeR7LtpKI7iUhAou7Fb+S2HXG+HoO+bcIuwfuLPJgLMu0bgN0LjR1z/v
Cm6Ei98hwqF9c29mIl6b/lLxALw75aa41Vkt3npAi7JwtLqix30Bq/1avqPx5OQS
TNrx/Jq41aXEfa9sohRiWmrV3JF1ptGH3BhWLSiiwb25MDzaeERO1da3SnCPG+d3
wtg3aWOGG3djC0gzAPKKQE4H4Da+hSXfQjb5JjsMZ7V8DTt/BAy6KqfFtlWVNvbG
yG8+rTc9b4WxSuee7htSrSrgdqSkArv2g8SbJG0p16Jcay3q0rIzDBiQJBJHAT6s
hzNUkZGfun29VzgxNPv1hBCmeQY5jPUUDHbV9z73oD9Arnm1Ga0BpmVYnF4XFQzi
kRfUxTGhB5D0HbMVXNyV9siWXnJMBiagTtKxTxGI2AeASNLlkqYn11yBsAFTUomj
U3/WCCL6ZEsGoKkcQm/9mXFOKn3yWijSILMU8JzJ9CCxw/esTegnxWNTpqXclLzI
LEykPm0AE379zUO2ykip1WIRD0WBY2h1eEPvnoaXsjEPpSTQ2dAV3rZ3YRZZd1KX
0gJxdrL9HbQpbzFhopITJpYyZG6dwthl6eYnT5DUIVqtAftV7G3WrQU+aisImzOo
7YpBXU5o8JMqLlq0eTU7TwIfiaf6SDUbDZj3BUvImDMEs8UP8OOn59yB9w7NpiB2
UGmr5gQsSwTjas4jWX7xD5wUx0r26dltOe5tzr5p0X369dPaNAMmGSFD2jtilnGz
bye9V/02diZAWpMS7mNrEsdkDLaOgs6taMb7ipOG8pMa5og/5Eu87B/fjzd4kDuH
Xq7BF5PGcCFblWP4DS1YxgcC0SVtqxTKR1sYAz/nr68cMBZUnJ+OCrsYUGFT54O7
ybz4HqNlynDKfr6YY5COU0GpP2DFjCRGYQRNvTl6eMNYOkoDbJ0+b+p77cFyo1X5
s5QFJMpG4VbkBETGEOQBGmCSXJPmrzfe0I8riXKkxYVD/at2cymGn+z7ihzYNcls
m5tt/Ix3MpvvAv+0nNF3r01nW1oTO+6LqclFsjx9ucAK5zB8/ElimzmL6oChSSHW
2QcjC5zykFNhFp19K/47pHOYvdrsKCnMQ8i3cWhYGqEmaUBb5plwGdFhklf8/MMC
oqojsUlGGR0FdFeL6O9y5+U8MNxn3tMjdBsIJFVQck0CaxJay+QT+0UMCB0S+gcD
G0/qL0SUfiatcMQCHE8AluyN1IerwM7rGGd4r8vOnOzfAGqXe4x8ct5ve5iuNmie
WxjDZdOxLdNWc83EJilWdWVZ48bXobqFTbZDEsV/n5omQuxL6cVDbHwfja2fwC4b
zLnVuzI6KRLjlrtMIBERMFuC8ghwwGqeD8GKUaAGMK2mBVMyOkQwdKKHesVkFhyz
IseqlY/W5vF1f5tN0v50eDzEInwjEm83Nb0z5DJYcmmYs9JloaRMSPcH+WuVOdTa
D85Y12RE3sYB82SEpo7aXxQ8vgIdsbOQEdHmAdQTOG2FBywQTKgzYxuLlafHEhj/
PwkMKaQMeXXGZTUw4NM6+S0ubpH4IWDaQ3zstzbPwC0LF7Dgwrr2h5x6wrIHwKN+
qk+ssiW4G6yg0my7oxL8+SGGRhXxCV2hApn0GIVD/IjZaw9sD2N4rYD1r4XU71gT
HetDLgvd3KxLwbKlDkQdwSt7ge5n0PGdXXnwDl17uVboA+DdLFEalSdx+Hj9T8Jy
xpYMwOi8tc1KxGPVnv/b/Kpqc5yYNgMMhIWgmnyEnPNfPTs7Iwgy6zMLb1a54UN7
0XrikeIpD/X3whqs/j318i4cQlJI4LU4ChrueNDaUx+HCHDRLM1WTZL/aF4sqS87
P/GA67FdAFkUMis9mPS/lSN++q470jRDBApiPHHb2mT+6jZBg0OKTF6Dm0a2J1rp
vglrV8Pb61m/KC9hNnk3I07MRKIykehlWOwiSDJlWE6mnYyQ02Ky4kdI9M97DL5+
ENuMubtyInazNUbfjwY7D8kK0Frdwpp23FMppDYpqVI4jeLV3lo6oq8bH67IoSNQ
D31kdR2ofc0NdpYwt+G6nbQvYmz1bkj6ss+lcJ3OAOMlFk/miJrcnSGDz2g/plqu
UZpNRNMLdpVClSnwULxiOIZDeFk3taa1m6l8c7ZGMn0NC34TSzQWNoSmu++ZRXCP
uPRrdz58INLPTWnL5hIAGCHLzQt2RRmsknEy/CMsmm5oXgexfxOBqlT6SndzH4mu
qZtBmevESs0S6aK2vWJrPCvoW2P1SQUA5i5/wln9ujpghHIu5g0Ia16wzoKtHnWe
s/BEp8gYSQaWFCrsZoUfK3TS21rV6vNPlTudiq5Uu7v33M3S3q0U+ox6IBpbML8J
5mYJMOlULlSTOGTsnoMCKasOn+7m/6GTJVxyWakr6nI77aF/EHT4MLqAEuhylCRC
y8GcJ7V6LQvJm4avG0ibAq1E4bD5KV+rCdsda0b5vtoHKFP3bLSPa6vRCpr0j5fL
bR/bxNjx6ZCGsKXkVmeUPSqsiMabRZPDgqz7aQul1CSw6pUM95oGrCzgnmjTAVo5
xGDYSiz6oyqs5J7v0M/WPfgQFe8vP9qNpUz+TBAurupaRpor3vT2JYk/lK2/kwD6
PrDaxY4Wfihj970+dB2lE++AoYclJPBN/S9794/V3vIbadE3rI/TAvJx3SboC3UQ
Xo1nbykUOj+hZLeMrd74maPd83GVfwhwcDRMNgY6B8M5DKoD1VEtya3BBi4K88UT
Y6RBxW8m6zrrpxhqVpCwtirjd6U0lYbPrLau4v+EYH6QhvMbuvu55D4Dn8DSvL4M
AEZvtR6UShGYqWXA9gUnSO1t6+VISjqps1vpoTzXMp1nGmioToLrWpen+vEomikE
mTn7d1ur4ygbjqg5bXSRQ5QygaX14QBAcr2gA/PNz76SFx0IDQOCMlxWPwic9ags
FCDj/J+SmxA6l/67glpp2cK0mBoqIxglKqsZXibraibZv0Vaurw6oK0tOVAS6WAx
gVakQiTtfw+/zDUPwI3OJT8e7O53pzt3knoAm3TR9GyQeQRj74XRsPq9K2c0S6q0
kxXtjjaKFnG2rJGz5bpGGq5mEefgd2uB0LzkEHUQfUcbKzZSO165P7nbMGvenZi0
0+vMAoANR2FNQtHOwcHRB/JoyKK8bI4YGX5gaewSTtsc8rZ3I4Kso3U8SOaHbRRF
84UOFt8Ka6zf1KQwtXfiiFDkhvKNkEeTHL1vd9/BeKW+XxXEgprn6M2kwnpcWN06
90l00TmifYhTUaakPqLNULC9gltzNN6833mjPfjV1wD7rM4V3HIuNpWwsUCAeaZI
kPIhJvNyA/ebXS5qE++RWyp/jrYnzbhHBKCVkSlrPGHcPCjGbblSwx/ri02gJnSH
FS4Cj1FTzx850gNPD9A+J+97pOQ2k0OWDezRP58u4utNnJIBI8Io85CoJmxDSsjn
lYc/r1lMxIo2XMB0nFaz2lGJfnaxg9pPRopWck6Lm9whtxZvy9mSq3ysH9nHdB2O
Bx/9snVGckevaHLHoZVjee9uZvCV5IIZx6deIkI2eY7G5qm7Cl7fZoeE1vMzEkC5
39fhgYG6ReSDk8pEk1UXUk5df2kEwbX5DDUO1EBY6RfzcD3sEEJ0tAT5IrM7oONR
BIfqDUxGRSnC+tOQJwjDLwCSNRuceRyjNnwon1HgQRkP/89N95M8+bY2jw72UDky
4lYnGS6Bh73E7cIf1uds6FYHe3dIRrhe4tGmFKPjl+1srLUa59kD8XER0A64hWUD
ifFEVEnbLgj0n1lIfQiZYVmk29PCCIU7Jutn5y3iMxz4iT/Kau1VF4pWBdRqviSt
ROZpDZdmXleWJ2kqQ5m2ut6xDxNSsl3eZ26GJcA/BXA5l9Nga4xGfuKOSK5+0WoU
Eoymqmg8Vd/jN4wl+x8jxWwKtZcHep3wBtejarL0zFBHPVlvDAzAEpLXGM8Aju96
+dMMJyBjg2EdS7k/DOYvC3A48G1jhFP1DAACCPmX/2CQENswS2Ceruemwbc0YU3K
0jrYzE13sYaDtQbmPnEtP/aap6PcfpSFiLpLHka/xuEb/UHpqRbGuNh3Ddn+S1jE
xGTzVb7qXWzL3SNSzlrAyRgMSRUOv8dnkYUNznsVJKY/2gWsYUNdlYTUX3Z83R7c
clvpKJXTggT2iblJfOxvGl2wMDxtEMgF5+cefRuW62nGLuYA4cz6adJPmoapC5XL
O2biVsFi1ZkfHpAvTPXjskqK8g+hFnd4HYx3o0lPTh4q3AfNSEecmcbkXvX/wwbx
CkCOnTJHD6hgS+l5CxSVoXDh2q4/a7SNsX3ZGnT0118O1SQ/oWGEIW6HXHh99Jg4
pj6PKV/z2jVkNqRO4IoWpbKDPY+coVpyWKzS9XcVp38tH0iNgxHeMGlA+okr1inU
yaLtQqJKv8q1F5/Q1a5bWepceeAL0BV6IcQgD4sR+wbmyaKNfzxS8A7sR/WTPFHK
h19EBJCzq6TZ4Jkm/pfwZPaWAqbsNQDLu4jQqqrQ6JsmrsmpOrN8ERqOw2ZEcKEe
d0ro5Cl3fj3iEWe9QVqAUnifgSxGRRLRbZezA41ZUUKNNp0347SYmk8dqL8WTsH2
U6kgkB41cg6N68t4LjjQrkgeDavxIHZn2hsb6N3TKM9aZSv99ZawOxLYHgAoZMmd
1ccX9/f83UAq8hCYuXapEVQfTK6TTbwv9AdyF2NAEw2unyj6ip4t4UPF5bhW/1Fx
Q4K36E0MtiITUgr818t+CHkOQApx5b2V3vYCGIUNhgroZ24T/kM7WH/QePss8v4j
Yg7C7hn3lpa3TgCSL1ExQvsYHjk5Hixl1yGTrwKFkeSoR2W83UUGkfTpCPbNu8BN
UEXPXg8JxWlL+TplUrsM9V4CS/kVKpvs67sXLplhOLILRtiz6DykiICERynAKc9q
fM0jAK52MNVpJ3qGdMuGJw7B4OqM9A5a9MXmTSZU6I3EkSJ0UUUH98raB/PsptVs
OS4bEZ4Ib5M3YeyK8T46dqoua3Q+aDZbOLPzfVgMG+TosgEcTjshdnuG37YDQd8y
Y1j2VGoZGfH3xtTkdHGJW0VaqHCoJLJivJRUMSIiKOfEN4/RnlKIVbLyHALuCMii
bYdRC7qccpiu3nzJPEiwZzsVB9ZxV63H0T7n9qUuYjHa5c91SBwMpIu1BRl3UKe8
zm66+ThRmJIKCLg6k3N6+G+SJqOIjfen6z2t84R265fBcHGmXWedjNmVT18s4m/T
50CC22Rwp5zTO4PAVCyy+lJIXJzH6XiDgjFy4dEKEVNdn1d+qO43bnm3msXYxI1i
DMNOoldNTbriWfLIYgr4SSVAVLrlymRwFvSm/LgNwvJpfiOK2/Tcw8r+MPAPTZMS
3IzCdCHIsqqBaHoUefkt3lpfi5qz8sxiatq+ZO8LoMROosb95F2Sj9FAjFd7kpnz
/LBMpWFkD+Op4fZ1YxUcK98E18iZWfGwtDv4cP6/J6JvR+T6CRddaEoLkAb4EGzx
efMl8g80lK02o9CXl38S5ks3DYawltJ25gtCZpo8DJCfq64EcWOTkG1jT6BsBsRH
gMsM7UbHeRVtfPY+VbVCv2ScJzXTqkUfyvKYetUpDomWEiEMRDdbFFvvste8hBaV
p706dwS5WY2FsL48V2o9uxxDmnzPTZmtb1oMl1WnccLU6ceFg0EF7qsFy+fLFLZB
JflWIIqUc6ldnfpQhv0BAJEQXgG4XrHB912F866agDoliNGHg+zk2iY1iHDZbo1Q
p7eUU8a7G8jcn9WAdNi516hhWyzt2RsGCY4JIF42sLQ5WJfBRl6ZdxqUZ95YUKwn
5dbl4xRkO1EgSoM4GV5NFH622x68EdMFCmQIGIDQMrEOLRU3oOeWoLH50G4i/4ep
yrVWH8cQuP8kZ94T+l0S2MojgNGCx0xDYkeaxiNVQprQ5p76iowOvKgns8SDo0ie
2mQCLAGjgppKGnDn/wjuvnYD7Z1ceX8CegHIMRYDTxznH/9Xn5+ueBkGXa6i1KTk
ijM1vFlMQQUGxOsCpsmx+GZtT4hlq2kdtsr9TaOXnbMzixDWn8LUxjefoq0vdH4a
IIjwv5+/QBUsb8WHNYO7WwNAYSzY14l1lLpMN5MqN/J+HXtHqIfGvHOZLWq9YM3n
CT30MRn4RuwbE6K/eLmtZv6VULMtWkiPsJBDrFZmCcUA8CSJ3dgoEpk8QBfYiNYG
EUluQVnfI/RhnLw1HfXvbNKAvSQwNWueLmPEx4ENWgUVZtHR3NUPy5R/rc3vdNwE
Os6BsJOau6mfSMdjnw8H3bLOXa27/3LyIDA+yfldgja6F+dLSZCGyNm1JU8nij97
Oj+IAvsqY8IIjZdUYqWbKS9ukNGJ+ZeeX6oxR8urxHeCk0VLgjvigWwLvLz/bS1j
7f4kS2xbsGflSnK615bdJxBsZUGHcnKG6dYGNE0NGA7XWcwEfs9iY4pn+Jn6Qffr
IekSacLoIUZwIbvuuDFyLWlhnHtxJKiAWUPUDWsIIpEyXPoBLCBqdA08oBlef5yt
XsYCj9rbonCSrlQtq2i17Ve1cuqUhvnvXBnEQsBVs9c2KVgaqNoNxB8m/Zyyr6ui
CvSo66eRr7lobpUiIMgF2GNiJVOwUmtyr1omYy4NOAf/F+gT+xA3sSs1Lf6sNeR8
Nif30AaXoP4lpo0W61wBRJZyjnXMUiJiSx6+uympN5LwQ4z3Ey+wG9IImIOksQdk
5A3KRdu1IGY+L4qgHXIWwjaTYCkuKFHpWcnoskjTTKCU7Ys3Ztx12Hcw9ARlXj9p
VxaPKBW8OA/SRT9a7JTnceRyJi+6vNqAefa6ea/7ErGF+AHRaprI6nT6GmSxy+Aq
xl3uO6Qrkn0+gGtDMZPZInLtDMlOq31VFNOdz6gDsWeHfa+ixGjI3/3kCm91+mci
PpTXHckgtjirYJIUqPsXOeTtZag+oAbXwMy67LHElD0tdmy3AJVE8UVZhhEkB1OU
V8uiOwSCMcDjSw+a4Dznxm3CF+Re+cKPwRMCPxg9x5nbmHcyiGEpZ5M/YetZ3K95
qNhZC/rZ0zmS8iKbeixlT3hfgefZZCDUZaiY67JZ7juwfCS2ShMJmsh8lrdy/e7k
ej2XYXxaOeZ4L3763sNyYlNyjyHpUcDmUwuS2SFY7w+QDrTN6yH8hlIcFUXomH0P
gh0l2sHeD6zOPEUIWe/EJBM5/4rzQDEnKrnUxX75ogE0ru3JEW2oaDaGYitjf5Lq
0dEC9DV/+/pdh3y7AwobutrClSrM05yk1NjMY0LLmriHBK635fRLoPS1MvY8Eana
HxFlB7bEf0xA86B5Urp8fPCEwX4rrbkyYOpZ+52fl+TEXAMEGo9cNxRLsfLA/+LL
jE3X6iQDo7KmUfpL5x2buTWWooOoQK5Tx00PI44OSveqKaqfCx/AA5fEMeaZH1Q3
EKaNsviXXF3wI4/FCiHpHDLz+sPVIE96lTSoeSFoQc3De8Am/+yUDXn01TwisUNy
Xfpp/G1vUoeeJoXn4+Z8PIEFCQ8V9eZ4BJzOl/3jWXi7Fj7qm9lDuw3CnfcsX76X
7+cGcPwup+ERMud2cQ3MO5puI+39TbILqf2RBoAH6esLYB2DyNYqqI6s+OYtRy0B
tCuQUW4lDSllqcP3tR7//9xoW3v693gs8esVI0z050eFbJQE65SE38f6jwg+nucw
WbqW0NOa2tzG4esUoFKsbw5Pb7QOqjSmEtwXRNMI/RK4doJvivkQcLvINO7YjGE6
jnZH6GAH7U1H0TDLEYaxgqGrSQlRsEMS71bNfXpAMB6JGAfOeaFIty7lk2V9/kvN
OVBbdFxd4cCM6SHbAp8VSWFtjIHhn70pzIL6YiXyHHu6l+k80T07Q+rGIfFRvZWz
RBSkGHop7v4ZunSBDzrQZ1+1+peIZaFIlbTxgKrbn3b2xBDGUqG1ZY6JzcPdMcaS
0qoef+rVUo5ebu0dPsIqTs9JeaTGSAwME4JeDcZbIePADX0gAQWP309iXAlq83TW
qLegUD0S5N5sKpgPBPzRPinxVNquSVAAkjD/f5W3SGYeGq/Sv7aV4hqQ0k7VaADb
daH/kcds3zpPu+ZhFz5WqDWu5SMEU2LqyEZLcL3exm/V5aEicRahlFVbY97O45BE
3jP40ZgPL4TXHhD4EyheO39ZuflZSLnGRxiA3Ymi6d0eafim3SddrqQutHNaJD+h
xhj3qRmjoNKZWivIEXOoTq43iaSZOBSbTyfvQKQ3QV4layIf3bQKqQBPpItpaX3O
BhuAP843QqvPLVwK4NkJCB7FtM2m6ppRmpYMPF9Q1L9IAKLSUQ4FdvRFgJkFQGyA
0prusrPGRL+lvld88NhTQFyVZFQavJIi1b/X46l+rs6bDXb61eIWwGMaYpcwEjPB
hbEYcWU78fJ6fO9CTpfNotgoV5geacIx7TXk76fufQG5RXf5TC1Do7S9w/RWNNBs
OOdncB0zsOdLKwC4nUt8GSyforKq8gZvxArgqAeMRTwzU7yE41OF1exITtCFh1zq
v5KkfPbBi8P+15EM8jsMbNsWCjCcK4RvQlwUtqdk0Iu57U1YDFEHSZ344eQNT690
RuG2wYYXsZrtObA1v1r864KT35AKp9d7pGCGzF0FWcKHAkRNb+1LbSgSC1T7pqKi
cEV3QGvARBFvjm8w3L/UcOmDhEfFvVJr0JECTJKyLMuoaaXwZc+obFDWSCjjfHDA
RyEBgjddZffSOpgCtmZ22jXIU+cyEnnfbA1P1ZbzoqwbbDJ36CtFbg1lbG/gJi7D
jMTTO+NcUA0erw+h1rcDnaavbnIUk+ePw1mAbfrOvuELaPCYjh1wpmJaiuXVqhmw
0ijAI9i1UtbDWuTjgtLgAgjuGrAjXgMAwmiqOkT4fXi6Y3XwCj0rMGw03PJxQ4C0
bkaStqBNro/FR3aYCty3tSQmoyQ25gKoG7no6YT0KpzgPMdIhAYmB8uj6bvA+0Jv
PCx5U9MKshidUdN87Z7U1yB4pne0dTbvm4cuGueSqzLRVaVXd5e41caQ9uQojhu4
SfuIXW9HbcakwbdRLWUodO3AFKjD6NrkYrqVeYXcRuKMv/jiaWbtrbo99HhRtYtq
rjzbdwLXRG29fo+9k8nTCrbn4eC7ygIwPNK2yh3TzobD5q1a/HOUUGAtSxsQ+XHa
y0q5Xerv/N+5cdqdYkoaTWr6uAHBHS1VqGsx79b5U49/REa5Z41tYJ1CG4B1fa6a
d/u+5HD1eScht4WWDrRaFKRFJZacT4cTzKG8v86nywVWi+9QvsWtOXqtFby+sold
87gPaqif2K4uNPHCllafhqF7JwDAidjxbzUQzDri1Vo3myNfwWZeL0v62HM9bLlg
Mcwbj8paNRhwYk9wv8Wk9MsYJet4A52xx2AXs9JGqoH/HYoY25K0uHFadqxlx/Fz
3A0Z9UtNIBk5T4yiquNhivdNqAwoIcN5sWgGrXHBqNYujUDK+F7mP09aucf2GAgv
L71I1MEHLATT5UgZgfcyT871WeZK/KbjP11XsGqmXGp44s+3PYXf5WPHg5ibzLbs
vHFsPo1kaB3DIIZJaUn/GnFaNvygddPAJ+iGfedKQJKlVriJzrJhpJNVa8NCi/UR
cRjhdmsIDiSkLwz1XX8r6OctsBZSuJJi/u4e6u737mg27QjRd9b35+sUvthHflBp
au6mIP5pQOIq4nq0Hm3yUVO05eDlG4ipR9BiRlsFCDKBMXbwvuBUsqWDL0NSZA+Y
9azC3HQ+/DlU594wMYaSRbvYanNmbu1MfBIAptq7x9Pv2BJnaVeL2MQ9SqrgIY9/
hqZ32W5mKsUpAku8IEQkFHrrqIP8TzWXDk+pjOVEV0CG4ZnbXvTfN9hA2kDvarrj
EGQuJIorQApPN3LFAvQALZ53p5qtgAkzK6ffCP6fv26IkqU0DGU4leekweJzSTtQ
q2Ang4rMjL+jSCMxVrp8lmx4nHoVG6duNgGrc6w74nQvadUwMuOZ/YTZ6EQyaGix
X1Cq11sSw2eziAFtTJ4XY1Fldx5ZfAfhaV3YJkvM3/ZDizUg3LBoEgNSiseqPHiY
RIC0jhE59ppkjJncgPT9rcbguWtfl2hoI7Xar8o8Ve895PI5JXJ3RYsYrJqVN5Xy
fcLwsg+4+P+WyJs4GCSW9qMxH9jJOE4KFRaeDntAV3dO6T6OX5QFL3Dgog/DkaTt
6qzeijgKKFFRQ7dno7YepHsbKmVj4uiqXNUHgxIcAmASgbiGfw2mAHX0lQTf/ryr
RY3HGfNc3+8SQr5xyJNvrf2sp7bYd43bbWtaFhBBKtixjIfzYLztVoOa4+L8HD7a
oghzarewwoYuJwi00LvzRRKfeHBL7c7nDdIaV+hDOgK8uCtDJCb5kCjxYcoWT2jh
D94jSNnuiQnLjmct/5Jw/QksX/sdHkKmNtxtcwSWGKW8Ooo8ZFsVOcPqQrZ6kbuz
+v7fYBz3Xr5iRBuZqszO4qPju03habs1p1UK2MOsbJ8EdCsSvdIoNrB0PLYennG6
9GwOukbjLNGnBkgBBdgiu2YvlZSSBKxhbbDTgtTppGWl8P+3aKCa9XAxEpp8wlgy
MvYbrlx4WWb7cIXb6kpfwQgDIj2USH6BgIFIrpYKPfiG0a3ny36p1sn6aMNbFUtF
obmQw0i7laMmw+0SfDVimNR7ash3NdJUb6F+StTMOCEIspdCyT60CCkUheqR75Sc
SzHgcIAjAVNWrpiUH+VBE/U54eERkd1ne/yfViaLm3haBj2jte4Jw8NYsP3SCYB4
XifG+blOD7RDqjajtasz/dDggifeWtOADUAmEwEoZxK0yTnjhkez2aV9z8rwOl2P
IF+MTCudD7Wv3LjtDgcjy2fl+7KnXnbJpwSrO9hdzzhg3l5d3OIt8GDxZPIh5OFL
cb0RAgPIaupl64XZDUmuOPW3sbw8Xh6wq3sJN0gP1Dm6maymssknvfhexL9OCI6Y
jmboblPSlS9Tqc5YoO0Qjm2SXLnYpv66kh2GuiGHnrK5wCCl9ZE5/ggFlHUzcR5Q
eCTBzbyqO4F/fGpHh/vxYeMdLFmLG70FFDHnl2Tb4LRV4VMez8m+jP6WfFKum9Cl
x3ZFLcVeO4w9HS6jQyrGHfY3OGwfoMP4/koz+Eauwf8Hsn1T/oBajGFG7R0JnE/j
e8fsvCVBUMLfhXjsXwpIu97qoSxo5XqsGzFsY41oSYRwgSKiTXval4zfEpbdn1Jo
eUv7lSac4KSC5OaGkxmame+ioqLgOnH6+I7XiqyPg53lOm3HLK8jbQoXHFrW0Z3W
u1kMTdfrjEiKACsPWmDmDI1UHobXoTDL+r0YpF4/zuyaqjmiI35holTwq3p568qe
psPo1DtO0b+S0n9gy/Kbmc5+qLPjEPqM/ZaZWjPYjGFyBUmwlFXCwv+YJ8Dx6eOC
WkmKQgjNr1s4b+p2mSjDz/xunoqpDckS05fzPI1CYOaKC9rSWol0AgbMDnL+r2I1
34y/cr0gJNu3+p98IQLMff3gL3o7Fo5A4n/nLMTNgd+IOocdNW1E46OrqQBaElfj
C42258CQxUDRKECIHVgFgyIOFR0QUqjgr0yYRQ3Nlqo43gwl6oxb1Iw19GSntAJz
sQvubuCIFoLO3PwIwggFLqMAQsjBjD/msfEmvUC5DFay1Yq+4U+9ni9jWHJB8W6i
++e/B/kXtKfiqbULd2Khub4e1tmP57IqVngHthxHoTu8lzjqDRCwqP3Ni6H7EK+D
DbHElNzrOjPmmmo7+VfmLLzLRsJD2jCA1jxSlwmAYCEoi6P+czcUkqgGKklDgg+0
PFHzisgVTKpeBddm4DXsRnUxn1brLOmrd5dMNLGzjCLw7etGZb+4jtCikhQ2377H
nkp1roJBcmXpW6XmHSmwgfz2G04GnkzFZqo6qBQq9wrhYCWF96Ble5zYtFy0CY/i
cc3xGHs8K1zAVUYG9LkOv7gnK9QWl1/njjlrW0UcVGhBteL2Eguar4yzDSPZ6Zfk
7iMelCHGHfTsWDSOvjUnYp10Sxiz8iDH/zVhTmmt3phPpqJ/XAiZjgKkcydbK2nT
WwG+xf/mgRzcYyAERren+d4kr9RyLDCQluGIuHw6k2NQNzAwaOLXEQP8P0PENGmy
qxLbb7MGmVuEGEeSzEbFEkJBRlCrZ5zGLEJuJK0P1dXVJfqaO2PTs3agYs6Y9xBw
7eWQHL6e6hOsjiMIFSTbGqaNMTKJBcZ9Y/5mFRiN+PKdGWpK4vIvoYV00bRN8rh6
zk+j91Np8XTbKRyu77CS0IFGuOOEeWKVs9XbPS7UqZHB5gZOw2TjhToXiTipYV1q
x650jcrmzAHa38HWvuBzZ8BoW/17lZ3XimPMHWaerR8DfqTarf3al2327KC4dttW
J+iL0s4noGQSur6j5GMxBmzCzlhdSvYgE6v13eVrVp2VUKmpEOpRGmRd0RPtLQZF
i7XN+xyWWYWiZ6Xv9BL6zqyXB053qA/n+KJ5QGtaLnHKFEPfIQkCLRrLgqdyv/Z/
nlNN6Yke4ZH7wJTrwqjXJXF2RxmLoRNE9+JEpd1qtQNEU5VGt9ffmLWw6s0ir1xi
EWaeAxDmCAxmF5uxBzLiR6fPF8DI8qrclGElYfAalNqlgB0iiBtIBKbgjCLleLCz
0ux2cld0dAhx+NvCo+iI+W0Dk0+Vg3eUgzpS3Sdiyr/7ZRCTIffKegRtDhrRkafp
c/r1rfbHLhxSJOGqTxZmWBqOkJiuG12S+olYyxjbiidpB1r7nOhOR3+zzhF5Fyu4
mPtv5SOBg0a+vgGN3+kwE2cXjV97FheGFjxF+2UKe+pzHfYAVeVwzVbydxwOZ+rq
szMT+wvBggBCpWiqFS3GrDGmxLXXmX0v0Zj1npSG5BbwD1CbQMbm7TmlYV48uCGA
bzghR8k2c4ICOuZVEaFmQ0DBTg7h8Z4eYPW3Gye76Xb0ABlPmVwHmh6I9yYOLiLx
tI3d2TPqeYttgdMinJIGK60ixXj6fSAz4wQPnx4GlJ78Hf/qxtl3wlSMs3+prab1
lmh+FzQ5nWVbiuX5JYlAAXJ46026AlJe+FbBEjAFs4VWvWpggsjF2hm78u14aPcK
G8QlLTZSo0ukRhwQoiLGNBpxKHx1/9P8UBTDla7DQ6b2saNeJkv0Xou8MFC5gDnJ
ftoOgpC+DjcBF9N3VgsrGjXOSlXge016B/p/OFh8eXI3OWD43uOk7Kyl/TRU5cFr
AP+9R4ngxaUuHTjCRcAFb94dU1rysLLb3nAlfGehV4qHU4RLv8GXqxhKXE7v/Hgg
o4X2+qyQga8slEz1hYX78CVieY+WOVtFhAh6jgDUXBJlMUuji6pj3U9xp9FdZ6iP
GztI6l3E/lVlPNXBB/VKrCRUXNzAPUdsWhMieGkE+7CvHDsLj7qSrc2cQxubxT/0
jBNj1e2iIeoT0rGKOVua3Yip5/Bi0CsYP0pniEI2/czRICFjqya1mzGkBWyByizq
Tj/of3nmpHnHdVCHlPiTesAjhUwXQskz/VGBTebxmdz4wTP63TSAWRF0mnI6lLWm
dTD8dMSq3xadtxKyIy8v8ziqoJoSBlHC7e3A7mI40YgPy9RZrb6Ef7jdU+mp9cE2
fmr0sQaKxOPg38gV/4RQTITb7WD+sWemCL+ae0LdGI8N7vAWTtJMbg2h1u80NTIv
wjCL5qgD0G6D7cQ152oRHkvbnC1cOjT/qzgZGKjRafhpMjdquYc7QaDNNgO9odCl
XSqdkhK7X692BTSmmWpQakunFzL2+lSi4eoJOC1g3oMKp205Vd6oRIBpksa0ZjMr
qTFJMgzLE1aW1r6iwropXh4XxY4SR01SDtt/feo/wUZwLQ1hM4D6B07OgHVAd6k8
pcqdPbx1Fw7H2M6G9OSPvKrX82sD0Zv6lT5sQjJfRucWScCtWwvDFjcGpn5BppB1
bxfN1Q/s1VMtv5DmtcgLoDnajCESvvESfm3psRiHYRT/GmyVQPtKAONZ0gaMDJPV
Tdccx8aUjDW2+cTLVczIg4dyLcL1qaaCj0VzD0wd+wRromAoDRfVgpbfn+QZx9vq
8lrqYv1IvCjS0QQxhMS3pSGbByMVnhKYIsCkIW1pcWEZF6rLSWwyPFpzK0UagIMT
DIejvm0xVENH3r2BwrWf7LHj6X21k1cYk1n3TORzM/piM6/+7j5jifcKReFWdbhx
OEGps/Kv9UcSL9eiJCmfngNSEg0iYFiFl7kOHzoWwsMeMV+zWBym8WnEI8a60v94
5C+OcNdPLTIQW3nFgBF3DLdfKz8Jg+UX9g3yaRUBcOIGsAN48KcUuPXG4R21qz/p
iC5l/DfoEFA1KOfRpMUpv6xZOmxSCus5ZpIXhx25LVjA9aV1CiAUQLSM49zWOuoH
QGfZDd6YUt7ZWu9vkQ6z+zOrwYjVZ988jQHyEmVUEIhX3hZHzvmdMUtgwr88jKAW
+N5R95BFr+rjC61AVIg1dzA+xiqsaXRm15gHXNkwbNIBjjBUx1FZPheIpbKv7bhH
E4/wc9kKI/gcUgfj7KJJjs2/mq9NKzVairMouth77sjTCcYniok8UtomldKIiuf1
xHbHB6jUBRnlfMv/QAxT8z/hAvoHUQ2ERMfnORkhr+rAuo2Pd9UgNMpmjvXS4zSj
sZHtRjDKKLHqCvZ/xw/crRyjLPBk76vJwE4tgxVTCaYf97Fr69wlF5yVr2KzxNLH
VI3KAPZHBaZoWEqLm8ESUiMfkcNfWsqj12CO8dYmo4KIokeAamdp+rc9jjT8uFOi
9hLPK3AcTnsx0xzxib8ZmftDBmrR5CclWo0ylmoqP8vt5q9Bo8NRFEbBYSG0LTzn
kt5cA/G7P+lQebglUhrZzvEAK2DqReLHUmR1d88NcY+P4dFyBIHjpxI8I5S3I35P
pGTS4AMaNlVeAA4ZWrv783S+vYkKXe5e9eW73hWuoK7a89kdxht6YJ0CVwfv2lLS
uyoSdvgEdqh9VM44AMuvK87aEX6FaaPUL69Di3qwRGE4ZwiO66BL2DAxsP1BLjzG
rai5oQ7Mv7kUUHOGcc9f0WjAPduOsjM8VG2qJz5kJeYYDTaR3di8MZkTLLLMCNrc
5XFuNPoGEEVRhTi0Ha5TknzB/ZdkIJJheTI4pX8MUiqSqMHZ0+AjJzCYzn6NCCp5
LpXry7qZJvWnDvfL2lE590SF9gjtpidWgXapb9tKjaPEscAdnOnKwvKWFb1b53DA
VrPLidM5J3kzNi7LQprg12qfeBzyS8Y076IDnEzXv/5Dxyym2NEBZOJ3a3egkR40
NUOFte6/xUcNtylrWkx4ghdo0Ym8RfFgFLJpTm79gQETha+X4LbsvMLp7wcHfTAH
3MnB+V8QmU6zjE4epbOqTG3UNQjViv3yVZHRndKUylP1CIe3Atqhj7rwogjdNKev
xrify7OKWb88kIs0G/OGyf8ZBVBCPtVlRpTtWedP3Y1bUXbdY3oWUKgOru/qCB76
FHtGFmEWSJExD1qTyH+CveNjS4ZJYJdZMPM4rk/0Arxir3zGkPHonVAdpgRwF7kq
/aTJZ9Q0S5qt4VSJN7hXZQriG9cjuVsv2yzN/AJSF/mdiJkANdJ2S3oLHkuTWsge
oAo+/xRIlnQoI/ySOUk14Lh2DvLl6c1M8WEwTfHlR79bxBh0JjbXtk4LoyPezXkA
9xVmFXaJhIJNg0x3R1pdcacJvgsmuZPSQWv5c6fYojrNbNTd7H/vyH04ffzLWihn
bdZ4h5rfV/PMPqKFbMQkoB3BEkJTZ3ZiQz2dv3KXF4iGydApbyx2bomliq7MG5cF
lx80gyEurdexIY71xly2AmSW1H67LIBkJ+MQKRiVYTeFQJrtuVX/u8UV4yUZL0bl
1MI7VrbIA2qB8CX+FXNnWnby4rDCS3d77MjpV753Zf1+rrX7FN9xO96/wV+j79xk
Pl/l38l1rRsY1q3jWgTSm2/0zNF563XXxUQ3o0+PzqShzBLgdFFwsIMiley/Omg/
hdT15boGH6asoRvPPncUmCKMg5CfFcNR+nq11KiuhP/nNQs5a8Jn1VF+uH8i5cYQ
lgV7Ci6w2a15CbmjYQww/ycYhk3cFlfwsfVjdqy+O0WnrFzu3ff32jhnGnO7a+Dh
QgnGV+WEQB6hdFBKDkYpgpCk+iXvHT7l0wIzSL8HapXXZ07ERQpnMylpDcaxCJz5
pKUku2qwocPR4XJu2quXXIs09SYWqCurLOdLbvhlfmT9vYBmIf63dZ07tzehtTqN
vGxvNrY+CzLykzUiI/byS9TZmsLuXyH5kh1vmp/6DyFRDwoQeyu+yCfSxGWAbjC9
Ak9mqWCgju3wWbkmeE9R4N04AgeTJ7ODJHGXnQ381IIptEYV0zO72Ut9tU9fnedc
LoJ5M06wIZU3LEUMjByyEd/TN1+iiPeXKcsmYYOLL9KcY6wa+txMUkdmFqQo86O/
mAEPJVDgPQXpYBYKiNQbkohtvPtrPRdFJAfWWrusKWSlt5XFEMksITV7ifspPoy3
xtOxSl+lXEi5DXh7H3AIuJRoCCvOwOPOADZ2Yq6AwJSITE1AwTftHQS3K4jNiIIY
aav3QiAkw7UXARL5GLIIydZ3n+qq2V7h349gHwqV9nyUTY1Hpny95AulHhPJ/X+4
iZaHuefBdswZ/YjqPdKSbh3lOGj1P8zVWCtZl1ZeXPRci9mTh3kZQc5ODWtKFa6A
fpd37CwI5pLNL39ESbILw27ERR6HYHEdF6bqVi0ftdvGTZnXiCF4MFf3Sepfs4rw
7R5yOP9UEcmkFqHWm9KpRuMrrDiSM3n7/3S6OAK4lQ/4E+rjNRIgyTfAuAcvceka
15cnYke/oeDWs4HEzzBKxOzIs5/uP7vc0JQP5KwWGGvMeZT48NIjPZBd2ynJ1IrO
jSW39rH0Lt6/DmbdT+VGFnkVWpOgQtK4O68V7jwwiZX5WIOovpzIgJThNRSTF7EM
Zl66JTyEq7Q3Aayj41RV5Y65GtRj0YHMwDHANsbJ3yFuu0C+pNMyHry1PMYA4jGR
6hONVDyFtoPkBCWx7KwG3lFGpeNGuoM7ln09VycATSQZZ7kjvVOtDLf5ReJTFvqp
01vgJ05/GBD47RA0MZ+nMMtKaXeoX6uHkAuFyiJA5NruoATHi4HSvktqoH+3n+eW
8dqHz21m1/9YfmoFZCXygr0xpJu3vodqahBYh3tu5KJ2pMEH4PJIjEG/KUKzVa0s
lGwDFqc3dvRz5jQQkpL65IAN58m4c+tHuI5w7160VNyNgBN9U4w95smYTgbQXJoW
Ca4TII1KBMAcDP2CxUrywco0svZzZEcZYG/BTfQBBNA9rYDuQLMeEJ3WnjRDDgDm
bpEqhRyMfupjD1h6MF9J4cHarC3XYrn4c3E9gIYZhBJZAAFiDOBaIofRyEg3tepZ
WnjY0SN2PhXfdsA2+MxtGCkHexz7pUVS39GlPXBd9IzGOnkP5j4/tx10aoQ30E9V
l5gQVuluhqMpAd3Xk+U7S01fqZ4R98LLUR9zpQ0e1CCSrFeMlMoeLzBn5OPUh8Vl
yOtZnOmstrHao/39OaZwybqEw+jWBpT0R+PRcn3jlmcQQauMjdwpkUfnXjl/BTXd
3EAv2lMFnqY9Cn9wXvwnOKD3yvdvPY457dGJSCkAg/nUb3Nx0IA4QEGAeAg29cSt
QdmhiV82uOMuMZBTUnbkh4TKtJG94gduyY8tHX2MXBhZ490Iy74Qr+2zCCHzzSc1
oluQGy+hh5PXSsAYYympYZQ9e5lRE6GR8+3i7r9P9MwdZm9XmNFCV+Gra+0MMxWm
lNB3cC1uZS0Ysr1r6rq0LO600rUVGb7kkF45bSobnQfDnueDIgg1ll9JpAujfA/E
pMDXDidu6B41zAU961xkapJVMR5Sn+4q1xeid8ZQVgspOpYsI9wiGVQK/rnNveWS
GjIo2YgVgOsvVJy67sCZAxwBg2B9A+LW2Rtk0Zkk7eFqGECTSCa8ssMJlhfJEjxz
AlZs0VqO487n3IXCIEbT2yv3wNZ2iIc8DalhPOEPwNeLPznP2vgmnAwy8yQtRXSG
OKfsGhLtqPYCXJa0qqJDgenyLgwuvksTjjNwfoVPIPAjspB6Pn8bq2LFHzrTQAdQ
SKVnk5aqOP0TfBfXHhL3A1v9blB+rDG09VIA1GFmLt6nQqvfYM3qi3Omkv7vKb1C
3U+6XrxF7h+VNUn717Fu6YlVTlppSxxdz/1eYZ5MQ31uvFsaU9LRVcpFBQUPyB+x
lVX8H33G6EXxgj2u+wNRGB70Vl36UgQ8CaUdzpF91L1+jwzevIl3DWzV2E3MU7GM
AQJhE5Gp0RQPa+T03flvbCuP1rkfelUZI5862oLheSqCfwHnGuv90sQb4fzry5+9
3q6iydw+lKkjm30YXZnI8lSsVsPVQSiGdxlmTUpMXM7HG5k130XIl/HQjwswEr+P
bp+ju0vZtENW7T82iVR5hm5cPDoHRfcHfRHKbwF8T7SwvBiR+D7/McJrpDM3PNpK
wrVCGSiSbw6izTIVODFsOmtosHVTxXCovtwKkmUxYFA1lQcVnbYz3rZnLzNr5Zs7
a8rfAclkFBMRoU1ifAoApwl+MN4A9vURIXKweFES07Brso9xdwVOrGpEOjFQo3gM
25IDu4U9j0tr30HO63Ky0pIHriYJsXdOc01YJlJpaA3Acpiqya6i/llXz8uK0Ey/
/riTvz5KcxPiQ4MeJpnSqJgVqhoe1QkQ8GZptO8E2SY3O0i57Nt2ecKzMR5yWYWa
J2Qa5lcnkD1fiYwhgw/+daE4MZdH6IEFFo2JVn9pAVoUtMKqC8f120/L3+raWawc
dFY/AvzESLcW+RFqqPolrAI4nxdk2ntvm8OBP1y7rN5WYLIASLXzwuiDCxkRlfvd
x1zTeZ9BOdCpY9LTg0Gff6bbBUiV1+u61YfHyIuMV+aPDYXqj4lz8H+G5gfFtPqx
wBObGu/pAe1IGvt32R69ccCLaM0tR1m9NfM0HfV9J2mgLUFmt9aiJNsvg9QARV5v
mZtDvUCVSMCF9J0Hb26lzH6rQy/U8cl6HwPouiXwVSH4a4twuI6K6yGEk6d5L07L
pT1olrFj9RXb6vYyzBpT8yQLaw/g7qB+zy0sNMrDhtZPhiOtXbbEDFzWRlQ62V5v
UiwrSdSwgICRqxOoxuAG1b8Lg8tjKQ9TamqVpcrTFqclKqYs25S7m0ZYED6dyA28
ihbJCDCx+bf+vKQA8nuRXNBgfWc2EuDd2M+vrtimdB2VkDWIRGg+L8VymSa/MwB0
p5ozr0lhRNy2RWoCt2sAX3jC2yr5lgCrx7UaXb58I06JspxO9vnl9VTCYkYsE7qU
1p0KA7EuqUcXPNwPPRJubtSBmX91TajPRNLOv1S0YvN2FyZeYGjMzJZEIXI21qNy
1DXsYtqBE5uAngI/eIZw2mufhzXlJA0Mih1Z9pG4yp5/fV/C/JbMFJacNOyQWotG
F/X8WXXf/DtJqF/9Ub2T06ho5Hp6WtKcMQDMftZCmuzLFI5UcVl3MPCk9UqGwKQy
lWEmXmyje1neaISIqfzzM/7sGSlcqg+w5Ks60m4DpSR26QbMZNYuWWjjEjr50hti
XUKXPHrgBuuL5ARYLx8+y86oqFUWmfnr74/b553Q3N6UAioSc9kp4ShyKPgOCh1V
DTWoNRcXi1ShfJLoqFmxn60wOx/JNI0HmsSD+JHpn1mqbxo1fTVlmTijGa846OAr
zdUwfxlwx9kAlNsG4T9BeMO+NjwL+IPT0ECnLU5+ggVgJ8j47LA810w5CVEiTJ6L
0LdeKO/iT38Eftqw4io26fLXovnAHcZ6XNPrPEpY9lEMD9bRXxkE2hkAgM4q71JF
XF9K2+uVNyLtx2x4TvxPW8sqKRljkKKk7vttglzqp5RnaoIrrdKV+QI1IU2TeZ26
YCpOVZ99/J+/8QPu9GWHLvLmg3ilqEgFDd+uePTjZ0bLT4ksUV8Oi8Z4kVEZ04fB
zQkexRvaBROHcAVC7oIT13qrJlTZrDUVrauxV9x9pchMp8IYzhqNmVv/KA3NXYy7
+rLtNmO+p5LmRP10RheYhNTjw3jlpZGfQOR1igrfrWwICcOv98+SOwRmEvIPNyWh
HveHog/Lx8qNNBvTNmiHplMAEH4i2sHPlZeHnY12KyZKyn37tbYkeas1ee3wmvb2
3Y580sZifSWvMpv+a1LrkpFwbTGOo1WsL18YvyQ3nyz18ypm+EJaTrbTKPynF8fb
++i/KZdz9Hc9tEi6ghK91BqKoYGgrhnL0OWPWit5LVJtwZn+gUnTHiQdYli12aGh
WENDhDUX56f4boUyankjx8dLE1+ebDsuwaWLtmCWp/JK6/XAvGIkt0fIFdTX5+f2
3l3+ng6oyowMYsYPEuSM9u0HGC7wmIqB4WOmOoBLxC1pQ4D3a+2elbtNqNq5gskf
qqAAZUE93M6FAom8+2sdXnlzUHSm7w6cFZj+BWv7B7nS5PRxqLrbCFAcBGcVmTV2
2tGh/B31oASAkDCAJly8cZ/2tSsm44Lnwwfl0zZuCwKoKoUSLKw7kHdurLC9KKt5
2HutbcbrmVasQFeyP4Q/i7bnxX/2LUOlB9veSiwQl4nO0v4gbdNsSyldSQfM+gmk
jk0Iypc6hUbQ7G1ShsCQX9lxsM5qQrLBfZr9HK+XMNkSy5mxP7ll8jfNrFKsv2aY
RwS9Zm9lcSEuC+VVD6bmUTSYuO0C7wspGOFe86k4mTjum79O3Dv24kIKww2O+v/g
flCWxN8FWDQ8UUsE9IB0SzOi8/0txETop3qiJSA83Qmiktuo81P+znHdhcaiovLS
5X9wJCtBX6d4yON/RyUvI0lIWM+o1VTLkBd3cfk65B8GtNO3w5bZPZkyLjIHZuKT
HvnzonNvpeHS4ERHdXQWxEkTTbbL4SF6l6ZhHZKPOqvV9KmQX+NMgIfNkmIfNI/K
jm5vxY41c4qJjUqcOAdRxA070D4JmVclLu35ZgmXTyc4hJlQQwyBwfF+E7Dbac6k
KCkt2jIJBl01xwlvNOD1D43lYhS3F/c2uNG702Z27fxVYY1S3OnTu3+rOzUQ3FMd
07vYBZmTILG7RA6Nz3tVZ5tmumpiP7EnbOaXG5CET66ssk0O/D0ke/lqVAfcB+3d
4vUmtweZXdedzYdtxMrs3hEtClJzrGX7OjnuWRUmkHf6bQXhthx7Qu302ziizSXW
yg27QUhYQEZhwmaQyDJtNZZdBzUSOnYchM+LtQYRzZUahMqjVhzU5X+VJ9r8Lg+z
oAcmLsPQ5K8d3R+hpl8j2Lj8Dh6IrODfZsRnlj3GsW036lA6cjkbezm6bEpL9qdS
6yTVE+dLmxOs1q7zXl3+e+BV2sUykYmvEBRYUWuAs3A29fr6h9Vv5f/fMERNXLsS
rLcDsU5ATThUmrnEEibKCiE50efIOfzbZHUNPxvBPPygpvTDlxgXa+lBFm9WQjqc
ESXNGmK5qPdKIXDqTDiWm2ROO7qMhsvzTaMDbyzDxn/rooZixeBmc9WQk0UVINRF
PKqky5D274jXO2OxAd1e6gIgHIMl8Rl4OGornGnPJPttCw5JlOLXBAA5AnZ057Op
b5WuU3MUCuJ1i6YsQoWmjHFGZHd4XLbrA2L0OA6eIFrUPbV3KX1If06fIKADihfx
BGXdhj6gZCUTZJ/9SllrSC4JGBOhDWxzomnUefaknsE/DLwxIPVcYaNtgh9swVBu
5RXAbvo+7Psm6frH2MFsBIJdV46QlQWHbeV93H3UDxi+8LE/cJu2TxcYqqggyFfP
zyxJY4V5lKcY+5Vi9UvRtVSzcMEDzJWdmzAD8g9pwWEAmsK90A8QNI7zG1Thfdx7
K2idWOsKJVgEw0pZakuUFur1hJll8rFsYr4yUqD8W40trx2ONCXYKbGWUB/Os6c9
SYkyEEk2pHAFBZru3eLnP0BLSuk2KAIbX2gGfbmMoS12R7IH4aj8Me9o1JLuP/I7
Ufg14L6GBnmxu8Ah73N898hf/l/2ydz3BAjfjt4IIWtdeRnVe1BNQPiSKkeQ2xrd
09bbuxMwxgHohQ9TnLefMwHTSoXHd9LwCiFPBOmbCjTq+2YdhufmNkzCZbOT+YoS
FRBtRcSS+TwN8RCiUCr4mqRnUMtuEbQuclbF7YxYHmm08SAVW5m65zsn29gPWC5R
VXGwu33yOwXz4EUbcFSXZBf8ZWPbX21mLcglgXQZtYRff1cilmuclwrncTLfyaeV
qeeGbyDGkwV9TEJVCACaIwCaJ7n8g+jnMK80qWk9JcGnNnDsabYZOGeWkZ6sOziQ
Z4G8h7OiYPoAArtzIBOOD6pUUIr2bd2JTUca0t4mbd6Aqhg4nc4cq/vXvW85cWq4
NRigeJCyY0d9dHICaqfgTBt8BqOmhT+GYoSxccAMWO93CbDgkT0JgK9k4ohEMa3e
UhVeZtPv1bwTCMzPPhhOr+H/Z4zJTBLbDGw1DhyTXHIebm7t19Uh/GH2lTn1YRVf
zwa2V5Uxz8gdwRF2dzg4kiPHiDWIdnUohm3+A0rkGnjTfvPc+IEUpXR3wIql7OKy
9Qh5bMxfo3XAE5CF9OieFjwuuJUBp9wb8u/Ur1NGUQPHvvZTn7GEKzESN0dbrqOk
JtxnJxT4Fs4j308LlYiGaMNdR9S3JfWnGAz5+A0ytMYjFR88Qx+Nr1oo4tHUOaHc
wTTecNu2s0/ovj92ObiZJmDY/MsTaZrnQHC4YGXjQR8+j67+khQ+T6vXOzqRUWk0
9uQf/nfsTBl506k0N5J8Ae8/NcCkdVmyv1rF7lygxXIP/IdPTkYfemR1nmNyem0z
juWWAzoqc+clo1Pjg+Ws6qJuLN4gJqy9E7MohhBl0bv3pl4Rym8s/uYoVo6NzUaB
6leg+ZDw/SUbk3aT5/2YY9TAa6n7a6jSVDvLw3F3awE9rXwMVfgkJ4GadywLR+LP
ksEdxmOHNBLONFqxx+cmxkVn/vutIZOK9ZjyHbJhJZLU4x0rS9/3WQrq8tVZBReF
EG9Q61Hp5iZxghdW06nkQdH6m6kJ/iirN1DcRxjVvUjAi4uomFj6FO18fFkpzMca
kRNAuZInqsAhJ6HdXm8EaFQi3mg5NYfh9oLYLDLqJNNu9+YBGkHTF/bpUss4P2zJ
q/P53OCVYA0uchP5FRuvm+WMn9mPj03EAEM+KqBKjiibsDQvcLve2x/OEAk3ivb6
qmlZp68Eo3zv55Knrzx5XiKJdfloEAhyFpFpsSOR0+f7kaL8pM6WzPyKsPs5EH2h
nZzhKjdTxc8Hs9NAouv9Ez5el67HF9aUsaWANpogyOUNhHHghgCR5XQ/VTMjyHbz
KSPSHF8bKZkCm77VxNSL+/bWaj9560U4d6L86NhMZwkWLrPhVQ2RKXqRGZHlyx4q
lzRMcuMvv432+ngJ7eaTHQA+LRQrelnj2aomsVuHRfiLkRJJ+IHTcEp2CsUDp1j+
3RSPAoqQiznxWbeWGN9jf00+S1lAIagBVWpPAiQjOk158ZOzjwbi7AH3UTLHwNDq
XgbS9nPtWOzVp+rkKckGrsVGytmKY93rI74Cu4ULosO138EFJcz9OYg3dPeOQxwE
q+RhS23iAbvsNtHU8sRiCtGzEm3YWq6xuq8hoYt3/Dr/wNSj8smrvks1LnNSqMcN
C4sPaDUK2ABh5A25jxhH/7BWkD0sLxU60TIBXU+JxnCLhYuJdnanN/A6Isr3x6LZ
gSODuuoqd4vKNCI3x21LrkMZ6lDRSCCXfbwKmoTGgYX1qW4hYSR8bAQbEzcz30Jf
Rxp2OcpaG3pIKZbOymSPtblNygA9I/ZPCbX9E+79TZtJTRQGlM7PsONK8nfT0JjO
VMkOoB7bDcSNvTe2VK4JUYwcBztUcdWZAuMrv5QdndirEEjRebt+Js6lRVls05EP
pf1P326HQUVkhfFNlTpWp0jowDdcCmJ7rUcRDh+MjJw1J3G3ufSk02tcDhDjj9vw
EX2QNhaeWdzySEjbblU0ycUGmXFOlhcqfBmoHx1JQPlfydYXGLbrFcF8Wt1wic4T
/OW4HeeitwLk78AUykfs1jygOxNvYgCnnARJ86Wg/omyI/ftQ2kFApRF6PmIZxjF
FqqzW0cQRwe783O6SKjWkpabV/ppwz/KHrQa0SuTPV8/0NZYbAR+z/UGN0MG4dDn
O/iR+DuEBbvDwHqEgrQ9Pp28M4KSG5kfPcLVqmC41/wSjADrVWHgUHhI1RbblsPf
bwc4q9ZnsElaXnvdvO14lbU4WVyF6pjWKdY9QK3bLeg7OEpJnilVJL0iHlkL69ed
cKNCozg0R9dd50HUBmskps99S7/ZZGYOEL4k8koP6c++hUJskiiXtyr1MTKZb/SK
uP+EqQ4y9sbe3Tb06YfEDNIvq9QaTf2H+jUfL5gKMZ5b+Mie5s6ZSK4U8bAyK5Qm
t2QTWt6VVvqusNmw9StlvUWko4zB+7tRDMy6+rZBgpbKrqw8SLPI1wwowXr9cZx8
UrVtXJnnaLgDwOomECidZRWQtYcqtcAXbwGXa9uY5UrTfcWp757DwQ9py9Xyfm+6
GTpOFEZI8t/VRIs9z++K3FhRImqvHul37Xm6XNJvUhkg37brHgKydg6/bRey5b5h
GLcsInSOSIgcRzK3b6C+gKvcQ0NYXC+Rr7ArkBCS5wbKc4/7T8CrEfF0wfW1eEvS
NI4uzlzI8a2C7vpI7XdUgESaHZflM7nJ22K6lZfqbAvKiDYQ03I8ChMjfEsUJ5+Z
mQejF3rCHCmMdWwd/rvS7KbfkwNDSnob1yxSr5Yr00i6cVJ3FGu5lsx/pcj6Np4C
t0Vi9dVljbSDrX4x4lsM7kvg+FHznBh2NaUueZSR0fcHEghM8YjBqhisM5jNA/ts
Q/SVe3pJYNbrsYOPKSvcACclEKqVC+zaH1jrWpEjn/rUHTYFsTzQhwGWascEtF6R
+dyW3dLvs3jBRQ0uhRI4vw2XuoErL/P+QoawWW5F88BomGQbSh4dzmy5fIL0rjbU
mwn6ZlMXP3WSyiuBHcXi+Pi3Y+dnCG3TiUEMaf22KWnlxH8kLFpaT+tSjnoP42dW
CTmiy22qX7zEWDyaCnUt7urbvIlAp30Z75TyFkDzxC3fvyazZEyddXqCH5wFBDqq
ksBDfl/7rDR+AFLMNLO4tgWbtFGiq3tUzqg00/yY5gghbirXiu0XzG4Ki9eI8QTM
ujHE60d2kmmNbfjNBLf35s7yNKaiRBCcCN74zhuubPvugeP4bC2IJFsl5dP4qPxA
BG7nIa4/+4oYoUe4ydk+kuVcKmCs2Rz3NFnV1n1fDYkM6tU7pQs3Yge8km/ZdIYg
aFAVjKUHznN55iin9vjX0xYJSrHDPLj2Boqt2zcno0F9IXDo+hphrn3yjl24h9m+
f6TA4KfLGppE3FN4g0H6yTuC7Loi5lbP1pCYuQVQxdl2XEgD6t121WKWixOIXrDq
YIYjwQJ0HMIL+W5j1+yQjCvJ3eB/pDtmBlJWsdWr1bK3h/1HPDekdTxbM7EJQIDx
H2xPDvxqG48wNWZvWFJiunK+ci3RNhU5LtazxoQQCDQezlT99HW43o/h7ib8XdGc
aI7gyzrFX9Un5O397Z3J5S8cQfs6OEYvsdUXL4tlb2MwMSUEk4BMlqTyQSs+19IR
CukfAVQVzkZvld2F5dyF0ya+Riimx5+xNeSpfqrE9RnEq6fdODDWeAQvhWnexz++
V13IELYKrNg/CePIKe7ENQ4muyhThtrmj6myNPYwXlsvcjFA6bXW/MB+bppK7+OZ
TBxL/obBmjbqVjA7fWIQprrz9aCBzg+J5mwve2FxZkmX47sazYEupgAS4OgMORxU
6yCEaFrmeWR9+6w9K49p73auOaEMqo8vuDzPKDVcHArVuj3NlbbHgU6l3OMxfPXX
ZJYTUCN/AXR28byk7tjJ7yi0QwJYcL/eOrHRdCBb0tXqp7QxfhMGbSmR1sWEZFFc
DM9H1AGaDYu6MyGRASBAajB7F9jEYHRqGcX2xJsWOTDZ16bBtaJukWzQvyNc+Umf
MAoArr6ZtuEHte0bJQ3gB2+i6MpxkE6zm4jPjo8Wbuq/JNuAR1A0MnixqCUvsGyf
3Wk/I77MuaR+W7InC4ATbj4dQpko5oPBq4S/yZBCo6O7tr4P2sdltg3FYsoWuq3z
02pM01qdBdnZSWgsMthiy6OaHu//1+UqIKb9ObmL1dW3f/1dKEcfTPRC+g9/LMSA
GkVs0c5gyVkDZ6tjWZmTX0MA9Vb1Cs39Tztyd6J8URK15zGOIK5SrPmNzLTcb38G
rYB12D5ndFNveVrJ75zdiOeC2WlGjxrX2qCz5uOjvrAllRA+vD15jedjGzNFNm9V
lQHARt4zQjSWMX7ts7SJGshuRtMKLHqWNMl77FWK5PIzYpYWFcs2q0vrlyviMo9D
PSbTg/cL9DSc+ESDpc/36k7sYPCeq8xkxFyTuJgHpIEd+El7VeKIRQ1I/wA7aBZh
+BKgFq1Pue3hAsaAh35VulcO/B5ngS/A8uH0hOuISOABvpq/QWc86dkDYvrtJysP
DCO1OQDLuNnmxwSXcRyUAAcXEOSMj0m1j+64DD8I5gpRfFMuYaHb8LpCtFC5pztE
UEjJXocKVZMpUDTTMe39VgbcuFEMwfMuNzSaYOMWAe1Lwlpa4u0iBGCxLrdt3Lg9
A9QnsKTMK8WrPyFPWken2h1SxGP+0eu6o3yAy2NncMZNTFVnOxW7BQq4IEh+V6/0
bf8RtxFMzKWTV3q7D9a/+YO0mar0mU/K17tgui1ZrxQmm6+qS18xTPm5BGnfBkma
reZVHiz0vdoy54upQJfhHwbHy8CWdsbek1OkPFSe3VB+tWYGxhBbjCdLVDS7/R6F
OLIz5FC4NSizbLTdZZF4TTt7BTADMPUx9S97t4NIrXTsOiilh8bLmldqsKRBZCv/
oLjxjauVqJU0AdZu2aCXg1F+Xq+VWwuRvndCv2FTXoTN+5CSPzIBpGVHsE2KOMyW
YhZcq2YWBAAsUcUAgERp/tnZTNboy5i8l45cOuNJ6kvBavXda7fwUqP8G3hhOcbb
XnN3aXFLneJRiM0KKey5Ohk356ZKcvUxCy9XOpsf3lMoNq/PC1XflusYT50ErWhv
sgFdN5BFxlwqOLjaJZgu+65zmAVmGXy82JJ+hWovVWbXzsQFGa73EXh4J8iTBVVt
ewMbhPjH9ajVsIVM6bZK42xOwcwBlkmlvm6r50DEoIckMySDZvH9ZfOmunvs0gsh
ia+8cbFKBPmYcjmxBZOBHHoqaefqvM8hvSXoEHyHWEr76zKkcjd6J265qX13Ovtn
dVykeW2BOHKJ28o5ZoLBv3fPWTuEpYDUTLJr9mn2XvlLVE7ovrhXUHejKfMr0q+V
Wg+jEMoD911YElAUNQnclZQaH4VhCj5lWdox3Q6V5oHdwTDHU7b9gQkhCxYZm7jy
Byr9sJ6xIZ9PZwP48sHnnY64kIwwxgf3zRQ9FFlkv0heYmUNMtutdlaTogfvycRG
r3BklP6Pmt0L933VYoZoeDzdc2pMxahtudFHBeadRUXZv78iqzAzwyyo+zLTMSzq
4LcnjOunwyxxhs0wpqfjLboq+OhvMUnOAZ/R4Hms9kjxxuNu1xJkbw+j72qejoby
NUURhFh4giGm7WnQ8IjxBIZyPiUZgSpIrgaz2zu9A8UMWCaKaEOtjJmOoLprW1HQ
P//soB9ndLG9nUDi/RKdOsRJSOI4n9uwx9HGJfeeKFxcmuojXcdAFohJxP/W3Jku
k1mPRYL1oEZXSH8s71kJwmspzdQdLcz27mP6KmfqVfv7NitV9KTa8CIupipv4s+k
4Lu48LXh8kKjhIOB5mJIPgQP49A7VZ2OCDnPSfapPhREvGvx5ZNvRdOFBgBLAT6F
Jaxw9lv5p/EhI1eMndTCGHlHeTVmvm1SifNOxQzfUlRxErKpXAqqqKJqx/jFlEpm
KsAjSB+GzZvoQgGXKMDjgGKuOIVZsR3J+EbGU7IyL6FH+SRHNfb6NBubuk0wAqkQ
P/2JoIq1KuKCgxJptdKtLWHJp03AfsQhM9/lXbmhOrvrwHXGsV1y/+eG/7njyBB/
3z8SfzQvtEj36xEgYytdHeXV3ygnvnYl7j9JSDf12N0qvtxPNhys926+ShWts+pm
zticeyAThDQIL9oQd+SS8KSiUl6seF8NZVa5CoiGlLtROkZN8LdWfcK7vA8Mb875
36aT52GojG9jagnQeiPSqRWaqeaOVk5XNi3DqY+kdrTotBq7ya2mhEBidFaqR39o
U2cBLGikv2/UnPtfDt0oBPiHMNL1vVaGZ58UWHfQTKFZfCy0czx/VJ3UdOMjOZcF
MXqhEFQqadaPTccxjZiGgD5hEBhwGT/MPfKSBcgEvyWayuV7tF6eQ8PAnELJCnbR
dboXCDEBgS3hq+PPlT5a/c4V3oObS4/q2/qYFkJRjea/1K4kn/CekijL6UI9YwaN
jky0aUujGZ8YcoSjVjyftsx6vpXHwm6TIGFWqt4THCVpYXXxfdu6VZE/1fKJ++gO
KqWWLpUEtfRR1EI3PqaUS6idr/O87VYr5SRbyqTbnN7MNE9fTRPunGP1VMpSClV9
hikG7kIXK7YVpAIFvt+dI2j37dtko6mjcmi7k1mX0tRGUqV/bSjgTVWreNSjtmeg
O3a+Ns0yNw7CaKuTCIMtd0cse6NO0Ke5P5PWE83E7EIz37ym5qVPcRVfCJtt9lwC
uINsTLAXLFp+1sOLg3bs9cSFPuntRVuByve1+VL1uEhwrGfjP0D6y01uZz/i7k91
eX0PpFP0Ktq9V7RP6woyaM0MD+kAAGt4lZ6Jd29o3EmFB0I1fJoI/RQb68q3rRbN
x1GJZN2666sOHLnbhm4LjGa/UMVAasP8ZCca50SU0G8XsfM5OIdHmTIMB09FPs1B
Bwh1/ZuEhBYlw3EKlsPpl51J6nWTQ1I/OhomyXUG9ubycFIqzxd6HiVRsORA0PoD
WqD5XwK+G7f8Uot2IJRRw/+BCSE6xh8tnqqRjklIVTog1CKspJYFKZ4vyjpdSs4n
Uf00Ua9PAOdl8g0KTyg9jnXF5WOGBv9l9gfsj1cGsRp7fabDLrQX2KKopPE0CXgG
UdpAOVAaqSVnDRWlNdzLMoum4i8Xk5O2+if9LRa/sgRgOE5Sb9ffBO4mH80l2lvI
4HUpd7iogTX/gLca08R+6WBdWmZdDv6dsZmw/XbhhWBzs5FgdRUJRs8ZwtpCegLz
hh+RDXaVtryWP0q054NVLMe6gg0chPlixMyMyQdkz7KNlsPVdbaP5fFunIyXPpdQ
PCeV9b/TVBsK0AO5fNHZuaRu1yqBgnOTU70vc4RYgPRK17y2N4p2P3ANNpJzGJC0
ctefyynmYARHtaIaEIQJMF+9+QHuNdw4QeAD9nIokBbH2nhW9Jj6YlCIn10SYR1B
AsjyVqlyKjLiXasIrueDIlIJje9PGSq2fhsDhUY2irznUJXkVTScpruenB4Q7U6t
NrTXBKjrYNNkKXEaJfy85wAmC842Vpfnm76VlAyGnwGwNbTyk3fiqQGc39q2osv2
NMaP8lrUH0K3ryMzQJisVX7qH5Plz2rm8bcrNNW7QiQlnubtMGx9Ma5jma3Ljy0N
GvHaPpZD/y9okY0b4E/qkOsA3j+63Si/1MWjvbbhxdnFKW3WzZj5mleU/sKOImQt
IARNxnwX5b8YSHdgPb/z1jaXdrZFvm2EM0iyva7oEFU8D4sPejG4Pc9eLL2AcCY/
e9KKFJzUJJoEhEdxaLdZY2N2USF0eANv+abZpsBTUdgmrteIUw+0WsRYfA+v7AEm
MTJMfWY/EqmyOJJq/H7QAuhI2NhnUY1nK4DLTZy89EK81W8/gZafZjlsLKgmdHQs
bqKKn/lnD16fgkMvbhrLT+CQgsOEG9ysxKpEqHBqm6slNwgVAs/ArAwewXPw7cu2
NBQ1WfbisxtMiG3Wu9IBMLMynrjS9zyVB5X8h3+f32VHHY5awz6MwBKlD5QgV9E3
oMHPtZHwGt2TXRJTo2lsc5dxX8iK/2JPFDBYK2ERgXbxMKGQ+7IA70S4XAPG4gCp
RI1dOfo7ttAHipjwCgFl+YrqVK8zZuGec2P2G0Mi3qcAeapcUYKHdJruxy9z5FTY
dsRS7au/VRgThKiTK0u+in112goFGIl/xT3Ayl9MeVwVO3qPFPFHJvS4f4EpIfj8
6aNbePD2aFBmKe29uENmGaMI7YuryW6ReNKKawOUP1KRqBYwfh5GtHN7miUEHBUw
78jMu5Mgp/AFhdse1vWTn8htEaVNYsW10oai2fD2siPuE0hlRLI/kb0FGVIVt2Xi
eHUNlKmTsibKEvpoyskFr4oU6gQ1fy5ilcfSqh8YK3r+qFIP+AM8UDiW0r7qPmUl
BBE4SxcIjl904pgY6a2wqh6bgU9EDg3FRx4AVrNhP4uPjtf2U3lg5LZki8cC8xra
mAS+j4uy9p20CpRQyTnwFA31+M+fYxOpIG/8T+wJ4hrBeKwCT5cA3FSco3LWxYuZ
bjVW5hscHSXUUpMS0srOnRVznUNunqpmNSUQAcUfbQVajqpar/ZJgag38LdQR52u
aO1Rz/eAtwp3oF8VWt0IQMRZfOeacpZcXgne4PWesAi5t9doihcf2GW8ZbYH/zcz
phQk2/LpRcm2hg7c3pEsWNVPcgeUlV+KAzx2sKcJ1UabSCc+I2A3E15kSClcu75O
gN8ZX7/PcIBETZcSYBTW2KnWUAPcARQKWtJnHuyyLS+CnGeN6pH7qcNComV+RTTr
6LegaiWWbj0IFHvRBHCku6t8HlXft6Mga6o/1wcpio3nE765YcjZcnBb2tRRrR8A
TBUWme45F9dVzHFFlKgws9fzQnhSEEDa8ioOx7ub/oCiOcllmkoHJPHf4fBMZQDn
dMLgH871OS2DCVVAOz+zk0sC3lD6wRrEXHVMO3VrgRzDLW3A8TcNPpZp2pKo5v9p
oUF4fu6Z/nC3JlfCQpfqzIGmvUne3XhvDNp91bdEvhn737R8luQCnkifKWboz8pv
P9Ndq7qdLDbJZECHx59B/nFaar0b6Fz/AZmCLDNla+nNz2xftOx4/s6XTmO/UuX2
aB+9g13V/UsB09yOETKEtz4lHaur7IHanHORVVy+IIqqZfiRJKuw8tZ+hEhbwRph
Amm13IoRKGkezPm38QNWQb+lGfZCtMd5V2WiYqaLuIFDkU5Z+r1+loUypRlUnrvW
yfsD4SfQedDX9hHElhz10qcrYYJ4bCZR6vz95twxJgf/r3vGZ2RN5BBO8mCjLE0c
uWSScUR20hekwoPWdr6ts2AqG0/byKCyuinGy+nFvsoeOXB/xmwde7ej1Bg4xbNI
XiLA+/MHTJzdud8G2wzv7j9aDwuDO5nCoH/SGbgWRTgUFbrRi1a7jUT9sS1RX64A
1RXrBCj9B8Y/Skgg9tKVH2ltHo64P7MwfczkNDdScQKSLEgCdrsCsEJPg/oaEQFh
gFkz21XxHPhUA3odav5oL+an7XmG4Aiz4SMDDfCX4RNNOTpeJQsGCLFImPVVx2Du
s6113cvFzapEZfQY4eda68qR/Lo9dViAhPksY7ztxDbBahDeobI+wv5S3PWgPjCR
XHyS3t5JMfTzZ5PGvkdQBIeQv6pZGL6J+1dP1hjgYzoHuGDewfRhJARZrl7b9aVU
jLY3/OH78ikFtDAY3rNYEjVyqav1RsKUpEXSvFsK6+NDYDAwqGA494FNIXuDxJRh
SiEReOKcxQZhUYTaVYDIDi8SvuiL8lQmSRHLBDj2/eSxUwQGS5nvemJCiMLs62sv
cio0dpbWEbqY34JWfiV2JQ70tAD4bgEi21P5h6gQVd83bR5B5tqoyHLShN6f6zZn
wVJm6Zkq8FCE+deH0QfcXa3jpg6cMnNTXW1ul+4q9q0IPOVndGlqRxX/xRsrXcTl
2yOTZCO4O3NTtEDOIUvZ2kKbA4TosMUTDJe/ld8iCK4iCHj6zATveXD2pixdD/Wl
hf1FKqZpnFvfgZaPBYwyYOJpp7A3xrtAuuPKRdA/jyanCX+5w9t0q2J5sYayINBb
/EZJfQt4TVy8Yo5RWYtAv5mm2O/qGnDRdRvF4id/xR3qvSUOtMUGiCaiNh0QfYqa
yZJepZcOpp22xTtMYGktpqL6N5Ci11HFgpQSxsVyEGDmg6pqJtMtlD+uS+qhO+rE
Sr2PWtQ+m7IJCWKftHbL5H46djN1oGNqfxzvY4EKLYtVSlSW2u9LXMjLc28HSsWN
OgHtLzBaAgw56KZPg6LbYo+3R9x7m9aeYQ6pn7JTVunJzcJ2pBnvNPduF3HgMvnW
5SwEowySAXRcpoWmSHR46b6KG2/I+87Jzm9rrCKkx1yDZC/BPHSKYPvq1kuxmG3r
PbdMZ9fPD6aTFOG5qQwzgrROyxm1AupH798qxf0CJ6t4M6hUCPtOT4l0Ozkdj04a
QkRFcqkCWjbKk2n7Jvgc1wSaKm8Kc5EpmkeZA65t8tLkOaII7tc9R7piJ4OqSIN3
Fg73NG9ul16hiojcqbLBgAAZDulRxmzjsmnnCJuwqxPBDWWzxRn+bgUqe9GtAl3s
YXujE7W5NdZbjs0FdRr/nBnf40pkTJsJqmrhQx6WqlUKJJrj6OWZqRvSHPC6BqTC
WPtt9wa42nPLmRPxAoXJBumVHx229J4LQwVubXNKmtMLNdfzougVrji3VwMn2Zg9
6078PnghkQAR2N4M87jqM68KCoEsjIlGu2dsX6u5pzTuJ94ujAMV4UBQvTZ71WO4
MANkGrzbzatH6VW0ErwlBc5hyzqIp4Hyt8msQdhfHBC/adcbnlKBSRfLmRX1C3Mu
uOTVsbT+bK/ZsPbOXfESbrtwRcc4oGEpUOoU7yFhUEWepZP26rFMT1Y19rJgZsv9
wWNQ01iebuiCWvAfyqxzMQ7DzU61/KKBAAsRx9icyFj1lnxI6g/K8vTTJ0r+jWyz
siHt6DJRvXX6AkYF5y1FDrK/9y/P1Fi+v+LBTHbsFExvLD7IABtqxMeG/DGdCuaB
y4JKEnR2Pfu48HBcqi5NtAtnQobKNlJyqItywUjS6I+RVJCmySWBZnMFHXP+AfIh
uCtApzJQKbLkgUv8y9arHr6qSp/IrSClDK3jaxaqCIwheLdnfOVXJ24mapxrH4jn
+wtKvAtFSa2EuR1lb3+XqugedwPbFsvKMscAmLbiBAeQc3dUnH+FefiletGQb5B4
uH6ejGt8Ngnc2oy1HFCOYPz8h6Dzq/w/AkB7tdCZqhoZOD3O5EzDPd90xFQG9icQ
uTEBA6wQrRSgkDXH8uMY7zqoJ0eNI2BXDvwF3VSGu2wol6EyaRvSF5QPYoxd+K0L
T/4v2tSubqtjLus6Vs+U/nnk/2Wbvy5UezjvdBvut2GpW6fOQ21lxgnjaJDYZDwp
YdzftzHlWhBS7rDk176yi0HVw1CFmXaXJ4WoeRJNfbjmD8uaQVa/eJ0VzcpJttMu
JAPfAXLiGVFQHQNNiyPJte1PaTgRmkQJU1ROQBbDGSPryxKEn4AQRn0zkPjlHHMo
eTcPuxbvk2ToSozd3xXbNpLr7CjCzBPu6+Kp/FWfRzKDAGSAvROXftSNhZnjrg4Z
u9Khwn9hqDsSyPzgCCdVDtwTJquIaoEFGoR3UUNxFOKiBClRNrtBSnCvVNgjFRGr
kvVZmYY1nuKxI4MJMjMzuVs6R0zIN0tTcFZOiDPcQeeqFwf8bDNzVUOsYkF4QKfd
DnM+TXFBd8QOSUWYACMZnKuNCGJO1xQ5oIy5TpCGbbWMoEFDLz1aL/bgjBEFUHFm
Yx0rk/O3+TdmjRS8eDHH0GxZUtX5lGf1djofoARY5sN9uhNgHHsEu20KHdrBDYas
fjmRL54pxcaWcWHUMj4Bb8Zds7dXYezMDH9I7D1yP+MJ2esckbfOU5S4l+j3Auoq
FC9mrM5yqnxapAnEDT7eCYLD6Tg+AJUQkrPZF/5IOJ4EMlVMHdkflCXgIT1F62NY
lxkXtK9m/HMoXU6CBciCp8ZJ9g0mVc2bdMI59etPsEWP91zk5wM3MuDr+yN1QZro
uyhVbIdzRjhjdoQpLymqScrN5F+xa2jvGt1h/8xVA7Lz0fR5tTW4OFfrCpC/Y/Mr
KnrQnZb0NUJS6VO5On6Zzfytm9v9d34DSyfhyrY4ezv5Kkpu69lIvnOKzGZvjY7+
TrPko8IgjXWYkwDGTSog1AOrfuAhAVZY5cMOCdEO08qappr4LKYXM2RM00tF4q84
n01+GjprcoMYQCi4JKrUpM+uTiVxIDkQBfzpnW/6tunXjPVwScnMR0xXvpJJ40xo
ynuQOzEB+Ufqp71S0SBP2gp+Ppbu9ry2YWy4hFEBcFZGMK7rd+HdiyHFU5AqEmKy
wO33BFB5TRiQXT0YTw1VMFkTz9gddFztp+GbpiISNeB93hlWD38B1sEdDfrTFMhE
iPgFmVlWsAdIkNSons8r/0x217eIxZzev0FEN8Clp3JFAUakVUw6VYiO69Mufc/l
p8gSougXsAncy3Byqy72oO24gNeXIH6z7lu5/50bDDdN606m7Ty4XG10cOtZRgdS
TphhUsEBV55XF6j8kukOJNBVQAPvNKlaugPE3gzsK1o55Aj7qT3fhyxgTdt/UyAB
Dszb0ehImTGPAnEWhWidsPoxTMJNhYxw7I1AooVmcLeTTyO90YxYfcILua9HwDhe
hs001iHUgsfNao1dDbK5yvmrJorO3mS6SL5iT+djyOYeRZnhJcWrnK6IdQXV/hgA
N6H3DB9gTL823aPX2X74F3nwCEmJCEivcYBtMxCjy67QoOtnEX+/7R4jGAmyPV4r
ROzDEdyIs9dt31TjlUEaOYhRHTvORERwP1GGt7/cNLvXLC9SeDf/f43phPVrHF7u
0HYBvLyjf7eF8oLPKUNzS/fkoa9p9Z5R042GkEBQuhptwlbae1d0GVn3Yf7xAdu3
SpYIUXaWrklNIU18d7XzDdU2aWmtM83n1gvM5KLAqhrrK83XljKoJl4VmHofY4K5
HsANCyEEseyDqzHZGhgYMjXFAhqFqW0lnmWhf7/d3cww6KRMVd8Yw8mUsHzIRZ1w
Ed9BX42GCR+hjolXSFqsPMzDI3twYJwJ7JBD2Z6+2PhOmYdxHFRT45a5eR6Xx/ut
0Ee24gfwAm0sPWyu6+fp76zw/jEqWfN1SraaPN8EJ4+LjOv/PjCqHSbGtmd858Qw
SciMg6lyCMxZfYfgCeaMi3nljAEATYoL61tYhCZ3I5/CbNMUvFtbFJ3KPQ4+ZuKI
qPKA4ZsCRFPiJ+7pL5ZQgyi+noyJ6P+EMgP5RhSpsGUXVcpmSHMFMIaBWkvXa0Ns
HBCrbirPTPDBEeSur4Cg4pAf59kLqaBODB3d2oIS/jYowXhOZ37xcirkumSB9h0z
H6urdEtHpvFvnDdQRzZClaXPJ06VOay+VzItm+0al4G+rqy4e1WTE/Wo+CunN0Gq
61r7SeSZRv5pCHW+5fRYsQVBASEGhC9cCkFY/dds9otVoYVM98/Bymwni2R7Fyl+
AA+pv7j1em9K/puSJ+Uu339cPMralivphcsIfK+s1mcVUu6nuD2eZxZJWv/BE0+t
xvp2wHICwWB9uROIWVs6UsWTRpkzrsBurfkGf8s86I64JzunQqi5B3a0qP/8JVQv
Yh0v4se3+hb7Aiz44C+7wofeULn/4l/YA9pHyGfd4Lg+piUDKzD4u8Z25q3JIwPf
pjKsRv5F5Q2GW4xbn1VWw6ORfIrkAux+Znm2AyfFqtxNSxdzyPlfnP3kipcOFrqr
S8XVLiLXuURM5h/rWnoEAvKxDPhkjBnnzx+7l7ci4qVxKHT2blL3T1trJsRNZSyE
PKapf+smuy0OzO1KHYsPLfzOLrB4w5xqqITWjBjoKrh64EO+sHDTX6avGKYOOU7O
OhlTpOMEGon4NRWujtQ7bZf1r71TaEV1h+kYCHR3D1CyJBqEM+9/xUAigxgEZDPC
eY0+wQB1J0TKWDZr06Hp49dPhPIhizELaBeWymZL8saswkiM3dD2wjnGVzusCins
Ue35/y7pqJx0zc44brjd13XfPPsEENlbCwSHbKaU/LPXrWDfWXLhmZugrx0LqbaL
x/Yk06f6mxzqNm7ERt9doMK6nY/K0AYBjH7bIMqPje/MNqAEfGQM67J+2Pt2xHZL
6KaGyRz0sVOWeDlgzZb5sfzuptKXXJA64Le1S85xX/dvT81PceiLpTyP0E8m6rfv
NMIN6lB8KrCjFBr3R3Bs/zY+fXIvBz9BMoJ4UEFit77jzFaTC8ZJlcmJ/Wn4H0RC
UVkQ2jOcUOxpxKeUR7FZDn0Kg8lz2Z7STtfvivUj/yutJslB1aZpyVJglj9ETkXO
JYzZGh00vlVre/fPCvd69REV1zidkS675TL2EhFG5+A29lUj1c5MvSkCfC2poR5o
/6bwoEnYTUs5M1jZj8Fxlkm8pEFBqUhqvVllJGITeYGBiStfpi46f8Kz0/pNbDy0
lfQk23YWEbQUwoi1uwujP8Etn6QJmaEJUo26jb0rXoo1y69HCGI1rnmVmP7BYaeR
nF8VJYNAG3jU/Z3VolmK3m2M17nTAr4Jc+JRO/l/PhXzfdf/f72eP3gtpfi/kIEF
YGJQVDXdU/OfFlFbjoikuDnm+xrDF1LNreoPxw37yHXUWdM041Ll8Er9/f/P8EjK
FIS9mI47nX4MffVZAyLMXFOaSSdspNbulE4M7kxX6ExW06sKDTinyR64viNAAEpu
LYhhO24BM0EWADNCO+gSoZWtSM4rVNYDbqz6DS/mYcRRsa4NsnBBoj+OuwsThetg
sD7bx1l8IO1QpNlvcBZ+nApgOH9koe8RhXTw0lPH+9vtKdzxsTobY63xiT9V8v9q
JZSCiXVyMZp7+iU1N1dhGTk7fN8WhjI1s4QqCrc7GdFRCwfpBLV/f/QDPnZIFiQ+
Ry18kjCprxU6VZbcQAwi3EqXL1ND8qlOsqZBZ7uz5/yGjBU7nu+xqv+wHCLQKKkV
xaZo8IscXaM8uydgR9OastSkquk67qiJ+3fZExBsOvL49YaC65XVxsgv9OM2A8H9
gaMn7/jvBBAN4xWTtoe64WE5GaWO8KPYXJHbR/hfO8I5Q9us+fENnGZW+03GeL8M
+wfZm2jH9IQZcW5z1UOq3IR/UMNJrBfqU2ASKPLCjrLPz5lb2aUbaQNTPX/d+33g
T5RTo1m2+ZeLkX9XVj1tjAfdYN3fYBkjvSYYIaI0dwvK0o6D+gAo5zICT2izyS+J
T3luUhUj3IdVlF15QlV5Y++p2H5oS9exqiJ2zZEuc19gxsXTRUO5RC5SbGmRndeS
unLnJKlcof28QZRFVAfuBRCOWDahj8m7msNr1KyHcFq9b+WoqgSqnA6zYIlSafyl
GvxhCqBkq/0VVnU/P/rGosWmoNDWO1VHOzsOUWRI93IiCWhwA1dGYsjJnypS9GMQ
9NGhmn4wU6BQUp9iXf8ye3yiDvSNh7pSI3UpYR5jkBxRIkIuO/A1s0cQZfYstAbY
JNdmxSY39Yb6VxgZD6hGJvd9dr/B+0nco+uC+nHDtrxtIlvRJzjp5IbGmClFAKN1
lGAHJh5dgD7/uLTkUVNlIS4Dg+wo6wz/hGRXf4UyDvVK4u1ugL70U14714mGkPXd
6SS0CR77TzBV4RzMcioHDvyyc8w7hNoRcAxjw0CIits1uw+KFSAW+pKEpsiQpbWd
cyY0G+OwjhgF3KDNU/Eop/f0nQfXG7dq1x0dqusSzCbPmPDXK1dfU8vOLDqVTO/n
zk9/4SZnBWVgHdOw4Ea7zw26nQOXptTH15Ai4IH/EpijHW8UPVJH+gzRGGm2uuHy
Ifl8VuLkHCzzoYEaVMFqvGD5liJeVRLQG7RzZrtMwR4qkLfFeAYUFQgUPFmU5jqJ
Ui+CtsGABnMUM2/bq+i+A7JE6gqJGPnSq9tAmsoWo0IvcUSkG6hRvUez7fB1yu8I
YxPqiV7AVEr4jq7u4up3FRDy3vgSEzBpxqtnYxnS3fIPv/ll6yXl5Lqrc/UWofbO
nAi9efOZ6HsAqliTaoEKacxJoe++2+eq3vgTpTLW2jhEFna6dGZ92QpJd4B5AOiS
8dmWeaieP23dah322UApthjnqMc2w3BPAPLFcC3mCoN0ygnFFQbKFLNIIp9v2zV0
eV/VOG1/5lV2iS6rvLhGOiVXeVD1IwGOBjZJl9nUHIuApRwyQY94FELu8s+dpJ9C
7r4Tzohk57Dhg/D1uPAKc/CxfTyTKVQRvv9bgDn3Jnh0yWqw4eiiwFrOl0hxwAQm
bLlN3aYlpgrGolKh8NFwSGF3O5bTqixTcJnF+Wu8jYInXVyUZ74hqk55GnWUgKjR
A5+qQ6lWUFvDXGuCY7ZB943FChleyXoPDG88oXpCEKuTwL39SlEGlyuoMXgjpcQ2
MqVGCQz+kyNootj49z/JnxeqB6N9obSzpr/UbnoeMqJ737DOXPVMOrodppe4Tjpn
5bgmLpGh66yt8ntV9kbaAFrv1IOfVNYRatG8omjciyruJhCQPLV9rSuTb2+Z9Jrr
DSYoZGCNMNcDm7f8B6SitbZYHGisZdMot+graJy3hupw8eK7eQ10ooi5WiynkuRj
WGXfqPSSXeWIz5PvT6c2fC5S+hHA7MvtKoTHq4mEQjYXbPhHduXaww6u5Lruwn0U
Pnituqocs/TE7pCnHOZEEpfBd7obJJ3x9XZwAWz0yBjqMas8pqqg9x0hazpRGxOx
QfBlJbu1z4QpznFBgAVRhVr2icQoQaA7tX4Uf8TzzO31Iey/HvxkmvXYStBi4bNH
MguToTNK9a5iW/KfrPO4carQ6C6VRI2oVvcmaiRZS+y5WsyifNqblSmHz4A4qLEv
75TQIXfEaqOd5KG7wZwNTKe/6UST/mEsCgxSaXlplmOXSaDR1AXZESueIRQm+VDs
JM0Fm/XUxD3wuFDg4jlrEFqpQREK0vN1CVb5iSL43imKpHjT1YEftymuLuQ4COkL
5SYehRENtuO/Rte978n+GetNMQOw+1bfPrx5J+tqmf0YqJnwHVPgDimarjq55YXo
oJfEh3WGNGwQsudtR0Hh8FnFnssQD8HBi9+BfzixlFd7IjS09X3zJEiyMmkhvvKj
Q3CODNBaXcxi52JBCSLM4bLjKozCYqvNUZojNZRTA6IxljNNG/jGlu7uBxbE5p9h
NyOPjoYPNsV7IdE1kiUE+zDLC3sJ53NBEw+yEqeNgtOXiYKfOx52y44LNowXdRzW
mPir0quLO8eR/5vv8jEYCHGy0nmVop9VJXUuwJQgtjEymZxh3zNWvr1WxpwXQrag
4GfOoPKkh1K9T+pmcXC4HdWVkEckUFVQaf74wnktoRHS1peZJMrutcM2HeGRnBcG
FObhETAJAdKW5ruxnYbEvWp1VzHby39Qy/vX9NKcgdWsEwNcYt3wf+yE0XCllmf1
j5rho0BK0Xtk5m/uNy0cKvGJ4n2Dvf4ycwHPLWCDj00KNmnKbmh/Wi86TCSBQaQQ
KT3C1rb9m7+k0hc8kZOR0W7vYGWBv6XzVtsNvs1yjsMkQd6ty86cBoCHOeMJ4ak2
W9lI/+SjJp+amBfDuqdK86JcrhBduUO/NNve9nVPa29jy+jePcB553pdLQeUliIa
yU9QDYisH/mPULX4KMN4N64T4gpVe0H+Ncr/Ghxfdz84oYOdvB8sI6s/+KXf6ze0
Xz//Jx5aNyCuKCAlu2f9zi3k6myWx7bT1e2tGCqt6JqXOO0ZXnP2Iw1Hk9/VAA4y
1M5M195Pn91aQnfp4TZuoKI8SPJZqwq7aKB/P5eBapcc0pdFypLK2hZ6strzqzh2
bqCJD7c2Id+o8jb+fhD0G5EwFpF1EPSqJKjDlddKhjbeYR+p9SmsShZGvdldqmVF
NxSBhSPeLSjk6n6w3GoFuCJxRqqSok9G+98znzByTSb42AnfIHSOGtnehpngH7pk
jwlxImfRmGPBZafAwa90z+sJSCp1W6JyBhj13Aht6VohrTUzEF94g3dmrCsLaHOJ
dFy9Omq8upSCe3koyCqVu12fc3agUtQq/nbgtHu30zlcfDvGo+1wqc94Z8INdC4x
0nVvsUpEAi42XZRxTNHkn9qEZ5J0uDbb6F/Lo5g/T8coznETL8LSwodZT9faLanY
gYRzDMGzlhlzkZOguK6YXpIR/rCB1b6xFYWaK8vq83f6ZRkoKu9HznuNQI/JCKNa
ZZEedP3Hxl0tdYDFu5qzjtxgVmrSFKAPSji8VYf0r3LKVysio2yEEQpvVezNsGFm
Y3yXdT6v8GbKj0Mi0NXMm6NPacfGjbbD3JHbZFjif0Ur/MwG7Mj109ujx5oACoSe
A/nq+YxjG4bRPMeu94m4bjERqnUq5LpESgJllQEOlecEVca/zONhBXvcT1RkRdUu
VeH4cg1cjuK90M9Xc4gQdxFFaIsDY/72E5JcSWHLJTfLUzn40sZ/bUVj1QIslGXf
0yC4uU/tDSEHepJicnNhLK40whrQ6uZEecfKBmFislUi3omSoHYDwpjzncXnwRPP
eCgjtiOvGEa16IipUi3G7GM4sRdyf+1Th6DciM4x5JhXn2AZnASDeXA/kqZP/M2p
PgRC23akOLqpTo20iSQ+PWNjd02+akQSMpaMGdrlrxU5O43wn73SkhrEU2MoGaIZ
JwaBRBikBQde4OYDOSN89kevHMkNTyWTkbJpNcPDqwevzJ2z4jk4Cga5norAcZtX
81MmzvhnprqmB8zI3djqXmnsalURIdBY/g8A0KCUZ9UkdW+n0b3Y6gCwH7pfVPF8
4ObSLw6H3lYs+p/vKOlTi5rQ+GrRBuCuBtRPTaqDhQigBSmsYg7h5+lOgX+FhTgw
aHuf3n+jzYQhO6JEQkWwQ0hyeUCyvk9MgqKyZkvifnpojKrfVrB9JMVYYpxdE6xr
tLiY07J5hCYvGgQ5bkZy/xNRncmOKmZ/TpUYs3EnPE8cTFw0pN0P3dKGsLA71WRV
tGabL8LfnmozEz//QK+IHtpFWSGHF6jSUqPvWEFrWISqWzW4NZi4oywdzLyndhwa
E+g55iNhOIVkuy1gjc8TLhkAAKmAWH7b81FsDL41vRp5pfMzpx12DnvD+53+w9c8
ITpXmKGkz+1R9icQgSeiZEqOdyCKPtIjuYhz9E7c1fmXOy4+22SnM4KVq6HlIpeH
hT2AwjkTNKlfTlPhepAjPMcRNDVu8qIAvyOF+t5lrhLi5LP9XZcbQlThSTICU3tz
Qfpm9quInH71RGEKMMy/1ZeiW5OzaNXQ7cgQ3ioX2ENlevGdaqz3yuL895+1YdF9
YMx+LdAhV0jrj/YZTmqjYkv0mzTPVDh6ssLIHdIdXVLQ0uh38jashSUTjEGNaQJp
t2Ub/g6ApCsX/k/vgjkfUSTm7p7qJ1OKBxrIuiLRWZnCX0cuI4PNAwujHP1dsERL
hdn870Tn447eLRH08Unz6Qtb0QERB8mfmG51CXamlY/OowiDFqZUCtqaO/RDi6Ke
q85wJiVMlIz6XusFgsvcxl6rmt5ylJI3RIebs52QfrGDZLKNn8uIMpUn8J6ZERZr
/XVJseUVBLs7PxVUyUqrxA7t0qbKYDRsmNu1OdzeT/5mVz1EjngQVYxnHMe0HGaF
/5ZzK1LnMK/aL46kSX0epqaeGq3mI6uVNHUC2LCCl+bA8d6WnG1675SSSWyGDGhj
cHI3hgZz0qXEcjzklY1ClMEZalJ8MmL4Sm49KX7btR4Sgt5lwge0S10rQu8jZko2
ob+wNM2YYjml5+UUq4cQrey0/dCXL9QDbKSvryJFdTedcRu/BLMIchM3oSBWch7n
rrBg4rPss5uKNGxhQxg3ZkUoCWuJESfw0pf9htERQ37ds4rkAxdOSRpR9ar4pCKK
PNPJEsjEDpyyaJa7JC+ypu0PxBvlggdOyhFmfyJgmWI2HcNmg28Oi/hXMDyXXcKT
3LTfUd302wv/aH74fcVzBkBc12pEhn54qrtlSl3y5DrZPUsFqFFbmIn9LHsGTXJM
qs52B7tKQNloPXfeIGXhalMVeGkIyCe2fBmB/X97LCkNI+p5Iv4n54Uedz5waK/c
an7H6Mz/nYWVbP7kNy5s9lxw7EujUKpB0WDd9QFFcdM26lBsNQe9ZgSrFs3vlnHN
CfJkWpK1zEmZpi2qiM92miU6PEkz4GP9YXWHSiOWYw4h1zFrDoo7BKeAbI15DZrD
FwB0OmGxpJfWAZsADK7x8qIRdYmHXXEG2CQXPgzIBX/MEo98dAS341lcuTfYxZkl
JcYzOyZxe1WGXUoq09fthiVVpC40dQBT1zibaZSKs224etarA+alcvcAaRSjvMHa
+HECOL0fZakd/LSkSX1HWJlmR79DWe4Oeyx8TvdalRXZE4zXlK3Onj2adpflqb0o
4hXGQKV6Du5g5tJvJ2puIiWNkjLXaY81xA1vEyrHfrr3ypX6bKjY2G7Hg3hHSAcU
RjAoByXX+abcSYigcD/LLN5+ZIKm12lv6tbnQdBqtyBxj5lUxBO0TFFpASHKj/U9
5CWLMYatCzYVpJKH2NsXYMfr8cQinbjmf5zM3j8bZP/i1kzuHrV0ZYgwY0Ebe6af
eEJ0O5Dak6dSTqGuYXHLpubu0/OodGZis68mHnuEszDVqS4XLQAbM/Ux1wyw0/YO
gqJ2546k6KeVe5MkXEid+jgBUgS7SzMOtjlaNp7Go31PnRCwDPc+EqJ8TYARkgWw
Keiw5dv/5Wr+1/iBeR7H/qWqtOKC+WJ2ouxYERoAhnt/V2i8gx4vU2saxCaiYiZj
IwvnYSpHzioaxwORC1ViVIYOpSgy+p0T07DQdXwm5bBTCnKT0yTbwQqXf4l4Nrni
R/x1MtwPJf3fizQk15kVPrwe1HItiICk1wqRYpBISXfN3+jvIiTR9Z8+a71kri3d
9NcVIYRb3h9md3h44uUsak4uLGrcviUjLyUplz+k48eZp9diTFdckOg+xdblfiLx
T55xW8K7vlK4jKDTZTdTXvMB9AiFRaVs9xAL4jWSs4gymopjNdZ5qny/hSVT5YLZ
XDnVTE3Ti7Kq052G+XOMH7+VT8xuzNKnJJZUxoqoY6AtTWP8qF+Ifkcetqx9pBLf
mMvh25O7SSsVrOed2H8rIAWtUePtj49oBpVogZIEqJejPBDMyiKbOx8A3m/4DSZP
WBOdMOuA7Q8ENQAIAhFCcFsJ4ITb/cjDGak04L5gbxU/bd9DpKncwg6lgG/C59BT
NkVJrdxkJPkCLnbMrdA7nqiowJ+6ZsSllsaPTGkCfPXMjeyZ6kK2AEFBf7lVNXut
1GiYHw2Ab2We922Caxjl2iRFCx0mJebdrZaScpp0o6uoglPBjKCyr/H3QXe2Shvi
J1pf4SF8nuVPM5XcWL/+RxxS25YQ/IV4VsGv5v7iYznNK3QLKUASGhGTiOwBnbgA
C2y5BNbSAOAJ4BS5vXqyyACYGb9lQau+5yI0LJC/kILqj41jAQ9z7EoVXfop2Zqo
9NlIrypx2hxiLapkunHkls4Mga5uO1zmawaL+7VXyKVajCkv9qulaxP+5YX3iR3W
XScd6YLv3j97dvdEZ9+rzn62PYNXA2BgsNJxHahzMp6rSZ5TPkPpIchAB3EAEwRW
OUI7mMLILS5Q4+cbi/GzTdL/47t8O3m0HNQnEjJHcJux9jI11LxwxvGg9F0T6vg4
7+YrZH2oMv4rZfuqrSbCotpShj8EqDAh8ybulIqX4ao88b2tF9SjbANMua5yGzy0
vWCemdYc2+5tiwQd4XpsQgVfGN7DeHic7GjXQgbC07MNQ7/p6XiPQ8ewVofhPriq
D7WHNwdTj2zOa5Ciiz0w0Ttf7UsnufKui4dgRx8/tDPbVgKI41jZjJNhpDFzltzR
yEmSEpo36M0gHq2U/eWGBo/k25GYO+l+qioOwAiPzjlwo/inR+vRqcDdHcceKFU1
15JgtzlWrRGET7WsNAS9vju4H/h713LlIsvMJl4bncpHRsEBI7Wp/SX3ZpTpHCdt
7ZFPgyYQhcMchbCoH1yY1SyidXGxmnokYFph22kSWBnC2Gfx0e+FkP2NNFhzKmEa
IpZlrsQACHmrtljsrXhKSezGIJnBQbAfuYaEn+fe96UMX8vTLV1nU3Ys8NsG12qJ
jeNdIph3qEB4QBenP44O6D+Lm8NCLpgdY9Xu0YbdP7ER+Ozz7NMILOes4LGvA1LC
5EwrTFwZbkl2Gp/zD73mby7t0Ig5em5E7nFz6KbwGcoCDHgt5n7i3WBDhn9E+xe2
uh64M5RnCF1jyuazdQJBee3KtEpOFgMgjt3qehbuux+DO1b34RcNQKWxv0s386K5
502z+Epfaq47LdQ33ThRy/PWElzBF09w7tH1Ozp3xep6goltAKO5etmQi3tf143Z
0+UysdTcih0rWTgxjUzHqss9n3kksFADdq6OoVuJU7QC07XHd9AJU0zA+3eAMYv6
e+X9pVdSfOcUo9bd6DJOvHlAy3lPY2+yspU8LMs1meNyZNplmGI017Ds9FZ/3Eh2
o6C9J84fD/l0tBUYy7AZvXxRzC5nyA4lgEcz4sNTw4LiFkKcGNqySzM7pVZaxdcr
/BgRdkBvKFgQ1l+E1JgXB2u/KhCwdCztfrbrmvwKU60OWWaTFXSZSdRmqvm12e5z
9p9nXzzXk/jjmEcuJXxnYFHncaG4Kmd7TJy+6T4HUXJGkoGjO8KApBOtHT4Q5htO
3WukS9ofiEKgTe7O4Gfaz4bFidI0HXoNTJRMLgV+oW2+Y+EiaRwFs1Dz0qf0gvuw
+uQYPzkoxq0PxXmrEBsn4Vvf69of/3vbEKZiCYFrTM87Ar8AvifTQycosG2klS93
lxfNZ9uBqJAc+Eh+osBLg7iLlivBcIJffZzEY3dJvnT7NjN9g0ZD4ad5QhZn3vmF
aLt5HrJIzQPuDN0MywwnV4/ioGhIFeG+GYi1OTc2AGsaLIfmGPdJJFQb2Z+I6gHl
klBg9vsAl1uCo+Z/VeR4HNvmO1V8i3eFfv+Ks3rFNTnzxCHbVS9t0L9zBDFRWW67
r7GKE9ZysMY3xavRFNKoZpdg95A1Zg8SbTloAKS4xsgMgzrZOMhGaN3yHKm5kO1k
nrUjzrawpehBTO7Qe2p4Z6JB6zPCQQofB8CiJpfsepSfOvQvau01cbjOkBBEUspM
gS0lY+y0cSDrHvEni+oos2qOOyCZv857KtXPA1v4F3PufSi9mg6DccTyoqizuKZc
eJehrv+x20KNQguMeFVZCrSUlXQ77Y1pBpRhvagKO299Pipklb/NDxGcSxvChkYd
30IXAq8Bu5UdK+e6zAzZaGRHwUmMJCmJK+WtiZmUXw0T2DqC3k83H/Oynaad9+j4
RdRahP3bevBHCIJeOb6TTnJyhWUVASbFSSh+LqY7Hmc/zoFo7lI6EhrbKdY3aC+q
CnqDqW+A+tmgL8GnXtsI2DOnYAstdxRrSxb12PG6Hn6vA0os4bTgdsXzNE3vZqlh
sYSbU/BCsj4jRwqcpCzbqfdGPgvw+6S55MVwVisYU8MvqcrKnbNeJAyxjTo1kznh
meiyDoblwuaZQSD5T5tLFx5TbXcHnoJPDl8uRToLsCLXuO69sh+r2MSXf69n+do6
Bk52f4UFCH8vK/dsh+A4euVu6yY4Xm59KPTmAC40bcTKyU9+rd6E2tMtyqfwm5Sh
x6NS2lEHxqgQdyuQ68A9ImTWQnkgi3DTvL7yDiUxTypqsf7G1O+i3nP6jPx7EYp4
OWwsz2QsOcti7bDKZPA10fZ+SOMhwLrmUSLki7jB42xVdD9uLElQP4XGwXYiHCvI
w18MRtuCtOLzcNlNHRl5gRAaIAtc92867YuNRHP+qAr2tqAu8WCHibrJGW0Kozvx
uZb7Vv+j4o1MCuPrtnsCx1C6BFW1JsoFbWuKdMBJskP1mTU1/Y2cOFEkntnUtz5g
B9OWD+kJGdAxAkfuCq2q/2Y+S82cufR5UcCNwuzNUz34TnBj2ZTWwS9slSm9wlwF
tOBtyTM3TeXqNzzvtEMmQJZDtnMxaNw+0PtRmqefYukN4oPbfE9up2U+GoD5kRT6
z2biMZLRgNd81m5XP6KoFaR6MhUayHsEhAEtk3KTOxx2VGXxOKvR2aRI+vp9sSRz
ESCqjTovEbUicBhd5cjFKUJvUBY2EJAludEjENHbsSehl/GHsEmr0Juq5wntBBAS
uFHynVGKofAjE64qHz0jUJAkPV3JbG+OuA4KxbHjH6oZyOmrTfiYle1BjFLHnPsp
FIEoyQfGmP1O1lMpIIxytNtNQpH/LgM8cZz1dL3MHoMK95hMZAKa5/gw6aW79KhN
wpXPfVx8Ct5hiM9uuKpbHNLzq/vKRZzXs4KN6NwEm1i0wz9BetJznBwEZVZ+Jgk+
vIitDfz64pxPZpdTQ7fQcXjtV9nYlFrNZbQqTUbdLs2nvuzjYWv+0NsZEEPnajZE
IrATULrQ+g/8WlHP8IPHmOIXZzK45qPdFgjsQmU4rNQfgNZR4lbWRZYBAbOSGtg1
48aXxnpDB8uwWWWn141D2ezT/bzQlqJ1sbEemV4aHwZ3p9sWcr6+aS6LvBDo+h2o
E4ndwgSf2PqzP3ntLdGUyV/ufVDLdrQR447ZKAWjdvdwvBfIj+7zR2Pf7bn4HFvr
TXyRFDlpfFBWuYY2+AGbJiLXY63SbTWkxAVAWImeB4By9x5tYR89V1zwPA2Kqx6r
rLdDpIASaIPn+fX06gLbqI1WcpNyhLDqqrg1RZp/kZiF5Yci/sLpHuL1DL/1lB+5
4thBmcD6CwWUEjvtG6eWyZNRxC6FGEabrccgRheP08cl3BSNm0nCUNIMh8bRuoms
ZydKrRCnUMOQcvWizXx98DVIaJ4g+NGnpHlfxDyGklmpYoBzpz2vwGEAXeu5tHCr
gTCeWm0Mo3O+ieiPgKH7s907Lfpikrllb2OKIwTGOjQJccvIeJiO6s4lKIzpu00F
RNixL5VJv8LIvtKGay6jGsTsNtPPCyF+od23rI0cgwFh7xqlAQEhRFcvMbxoPxUA
k5QRQMjWnpVvciV8254p4oIFSAU5dpkqSEHdaKcZ6zeSOe7HlO0yWAFRbTKuCwvE
SFGMZ1nF+4MTsd0t14wzXURrpiuZMETOdwSiCHMr5cLkGk8614pBV3q1r6KSnwJm
3BNwHVULUEfrWHGzphoKnkmJEF2Sk1MrTziNhCbX7aqnodVJ5rk+1PGyowd7Le5M
CbPIIEt7PiFSbe1MCc9NTBd2lLn+rxuRUAAaV45OtW1x4H0L0SORg1ClR2fjMRnO
lYyBQGk4hU2YMaQEl9Di7eCa5hVKUSYYhY7/RS8IPMzGemlMPxznQhaKEd3unt2q
VC+Ychgt3HBp1QAbLX5982JHX9L3RqVCFA0pwGwVGKKZTR65l687FfAsftwqQ3Pf
UW60GA8vhTrf+ZlKL1+MybLPSCL1PJNFfLKfiMzplKw52EPWrPIBUuCu8mlKIzUx
tyllTt+3veZlh2/VC3lGRbMLa1MZTiUBtmOFdbmoxKjN73D5bRCtsGz2F3OfvvA7
9wswjcLmhGOh/nX1WefzHU5wQRlOSySwz0b4P7IbHK3sOn9725B4xPL5NZOSqOCY
/JpD1bfPUA2zeDmdD09g06Sman2QmEg3Ao0N/hPEcAcqWIDz7/7UmVHnua0jNKzp
WGx83uhK+7MuXCbBd8CsN9IdSqX5/QCc5K/D/4KHiG7htVNGkmBEblDCJGVd8q8y
14rBP1P5yWSeCMJAv+KbPP0xyqKSlG3RREEuVx5ALGCFWTnVhr0lJ5EJRKvTXPj7
VsJmPNYvUcL5VQHqnp1ekpFa9X1i0uFQ/kCltinQoPmQUQcN5l5VF4MdlLSeTg3B
cVGTgztLXR90VMwLk43EitWU8tmtL3BnTHftlOqdIeV2LbM5JcQMt8CDdy+/70UO
6EeJWx1Yk4YLYq1DBX//J3nEa8XN3vPQY2ozQlQgxlTWwTC5W+IsWHsNDnHJv00v
G35Thp7spjAKmzHuMkrknnVwoLXjagY+ucsasoGKN+20iLzwLIA/W0nvJZLkOQl+
br2pB7MNPbJcyr0TVPtqxZTYCyu93UcC0Di5ly8rjfXtwQ4ABx0U03MlamFJXPCG
iMPto+elxBoziPnI0TvMyj9HgApVXiUYNSQM0K2/5qe6J2ePB8j4FLO2o4c8gWO7
PF4ZEYTRD/RWPxruUA0pa8psS2SeKSpev1zx37H9dO3Cg1NEMCPAnPQx8Eb47z5S
YzDO4Q3AL2Wh35OwthJeOT5nc6+AH4RxHUR+MgBsWn2lFrahW6ntlakDOuUodVHk
SLtuVcXt3lt5O3WpgzN2ss9EZtPs1j7vhAyjqVB0hVo1PWSJybOF5slc1KOjCzdV
uZDPoesdQjXnCQ1sMMrUBLKoEvRl18wqv8zNu2YoxFnMShJVDGEbFY6F5444NG+8
UtHdsl+lfciCHdsnklBnz7NBfsyLjmwnPp/C2XR+2cF+OvvEUhrsjudi72ol1c+M
lJUv800Bt2TvkbQEKYTVblbzRqaYYVkXatSp+V6ILFo1D6VcytYRLx/lhukhFAYS
G/Rt/tTgRjDyneHGaVxRArewEp4nozOw5NVc6f1H/79YSgOMTxx/15NgkWzn3UjP
rUDwRI4IdEhaf+0SAuQv4yaxTphHTS7I6izSatPqeOpeLydt8QMrAdScl4hUd70L
xVQ+AB1e8BI2xcPOIdQUii7MTGe/djf1jSn9uiVtXnpYEHkZql/ylx5hfiQWzE/h
3ox/WNHafw5Xk+erbNGqzlnivU3YKT+K9EIc+v5JzWSL3JvLmtevpw0Gd6l1wgSb
X9qe6aBljK6xyMw2gRJU8rk20VVQJoynN1YMyeGnTJyc3v/DXh7+kACccnziS2tO
F65wDAEHU8IKN+zNgdrhVwzNccD3roSKcX21bfGnwqrC8/OUbI6+7CtfYt6Wje9B
WC1aqBA34PE1oPPAO2eSSrT5UTEio99uszyGw68n/AGEREqwZc6QhFIO8lg9ZKFZ
MbVCfkmMKFhm26VsgemNTjPxkQRjcq8P4DSTCUQAjk0fzZ+HAWm8P+Iy68gYJJyr
NZrc7H5fJsTJ0BTRqwOknZ550RnRDtNEh7KTzM0h/f6i6eNQuT2+aTOm1AUyerXX
eU/Ec1d+VIa0qoFvwMd0na6LUyUjSIy/T+1y1ZGW8rGT0Tz8IxOq7/a2bRJdzpah
4k0GjW/suf/5rvdkWS9QCm05nDgvGyKA2K6Z5XChgY1/BznfgI0Hty6D7QfvNYvN
1y7RGqP5NnhlPli3viq8yu+xMUvBuSZLK1ZQsdDuwT82oFZopQgtwq2F1grCrUB6
qf9UKn8oBWoiSuxyLL4EuIYYm2tCV2ift14lBL2JYkmOU2Gc4p1QsIyzlUARpELX
6y82PZ0bfzdTFzZjCch8rEAFZaTMzt0dp5EbFJL2YCrA47mq8yIDOXP0kgqspAdP
vMYxXwegr0ik6UVPHHEzA+9uaXn7XONKraTPaJH6xPx7kgfSHLH06KC0TqkXV8Wv
bKKB8CdhqrCaAM4x4tLZ8TX18vEzwvLiAfvANYLMKJCVxq4PubeWw3k4kYgXCyA8
hmbniKZQukLtmBDgOY9Klrl8pcwQTNnmTf+6fDgQCaQydkU4O9EyG+u85ZHu4FA/
4BpNl8QY+KpfoM8OmfwPQFruiCq/kfS5oVc+xl4unoGdt3wqhIgH7ld4q3bV/O5s
5ZHaVbWo8lE/36xFsDvGFFdZqLFsulbxBMU7jFvY38dp0GXLxUNKIFAsotnfM4ce
OLl7fGBCogcbGuUzEgK2yThrxO8kGLQh15ZHSy/AOnuiFvEm9IRYKUJGbzBAvhWV
Mtrycg21IoQUyWzxe4KvJrXJZzmeI/ssaRBZS1oDU9VpyRnUM+LrVCxDpvhegiSU
5xPNSkO1HxeUAPuMSctWk41IMLKKLMCwVu+WCzi8dBpyoewOaTYeBi9uC4SdZ4Cc
lyojbfK3YGTG8WGkfz3d8y30BgsOqm7FmCXefsCutkc5a2tDOXS1KS8R54sYEFuq
6EM63suUklzv2r3mBQHSqqEfzN0hMCF7nNKA7SM41f0OehMHYZ0pczy5vUzm9qPc
0E8D3b/HAexH2xthanyY6k9iyVW4uqUGPDi8rxZtFSD5ScD9bAKWQUbwNfE4BDdH
2xx2X3RjWGC6kf7N7rzstg/PDlXMd+367sNiwhN8KojhnWet8FocxGNK6Sbd1OM/
RoSUT6FEzrfZ8O98sPBnQhk8otrHmzIciMBM0I3J2squwqmnMtSfbcly6J0V26He
a+GWRgdrvojdWN9zIKUP7VxQxcvBUkyNhEOQKhIwAMptxxBhSAFSLFY9wsIAnSAK
Z3gypfy1tqpj2tjzUysjgTJ49/wEUbTzW1bDzNjebi8+CXoyzy9Y2DU407iLVF1x
vOEPUdF6WH6bnVg4EP0fysRknOaGX/R6UIQQl18yyuv9bBsD+PnN8KY+eo8+Fu7e
Aos/81zF+nPI00GEcCRsZw9XEMrohfT1Yk6zPiaiGEFJtRpSp+98ClAy1Kr+AxRy
vItUvfrAYeGWpSbE2irCtVhT1II9OgcBrC/elzDe8W+POUmaRwf7MP912DMvAdXZ
uOWrClrJGYHqeIqHuB7sTvjF4S1GUznMwcZQ5UwSl58iYptT3Sd1hnfDcfiyuNds
zSXGxNfbgOTwQtTtA+8O29pvE3Q9sNlpAKnMqY2hbg3jeDOp3goJiksnwDmgmzP1
NHUusS7cDVNsVWDK6UVkWWqG64gpDG9yWuJDC4o1RAXoDDAbbVx9/8eQP/Z79GJr
Mste+b4WDnF/8AUllQKnMIlSed+4K72Z2lin8WAmMQAKJVrOt/B5aRJbWRQH4hkF
lK7Sbvu0h1vZZYUIyqojHuywka3I7fUFLcUdI3cLK4Q4wr0NSlRicuxPo66CiIy/
FZixyWCfM/PXm3wjY9TiO4xnMAV+eUPSQjLVKHJukDP3k7N0sRhk0w6J1zVj6WNo
Z/7SkXN/Q5Y/7R0ZzlbgFU3Jz3caZgmf1bOy6v9t1Z1ZTwWWwN5/ldYOKMaAqins
JdqBYQNvXKy9D5qHnnYsgBjJPox858PTesZc02VsDmn0yNho+RPl9H1KBMfd6dZa
wQEvj/KGdLmfwk00+oTVqNQ5YbudMJ6jIekwQhbk4cPoGUlrERtVvwt73dOuu2yj
j4r9E1PaUFYOy7Rrkml7z1wbHVa5OtYImnjkRkDesUBWe5dJNn8fJCAKS615hf98
S+kjmdMQ0jNUen9dRg2cvwQQ0ELzBQNcY8RIbY8WKZhkjP47c1rcsMRLeHHqNbcI
ugzdHlmTF0kCDNC+ZgheUKkDJLWlLU89Wr69vT0M4Jb+nbdiVoirGG2m/s9T/6Z1
fod8u9h7uCsLT9jFye3Vt26aYhsbtolo+ynX51zQX9G29zGRik1f5SBI45vQ0/on
HomhnXCoJq5ZU0DPVLo/2/44DELUG7MC9Habdr99YiQ6PDHFT9zVoQFjGGHVJHbT
0h1Y5qM8DNdsuJkXZpUXbh1WJ70EA6csKm2GKFZg0NA4f3wS0DYap7DZPSEKHsiu
ColxdFEyGikGjg/Z5TtssSwDF1vXrYZNNMxtDecrdAibvYRQNVMC9BWZD0ceNUtp
kMvEHMUU+w3P3ImZ79Inaw6e64UUE4r5krk1D7PpUFJMQHYLxMt4RZ/o1E43cga4
9Aha8R6gelji/KVysP5lHsWVQu0zp7HSW1CGMB0neJgeDx7KVYu6GDFVed2mJ2OW
qwThcHlE8WRa2u8HyhOTeAxhkfyJlGGHoyOe9WPNeOshnm+5a//BzAAbQusH6BEX
NQYFgpfI0bhPDyDrAFXPVKQAp2eXn9z0uyNF0p57DanpX4XAwGu9wk+cGGU/td5q
CGNboe6z2bYxG3frsh/hdn/S+qztPCMRL+shf4t2dc0tr1pVtkunc33/vYNS1D2D
PSrv76A2duGkEWlc6ZWoHXP7WL6FV1cXxjYRdw86lEVUERBMV9QI/slSTk5J2fTb
yVZwR6HNu6bbdk6D6URQv3ty/03+Q2Vloe3kQd7WZnFLIRX+aThFxf/hW9KcH8n9
d/De/aWmnWpfa17Da2bonQL0ksUrloXKoMiP7yaIdY4mBWtTwvHXFa+GBHU5TAWt
S7HVo99hu98EqJMf+rr92jh3PUV4pVSZOSjqMNfnyHA510ue1TRjaT8dFpb06fE9
uwmkC/Cd53biSxwGirswn1gizwsqSTwvc3Y59deRgkOyg8D1zfq+SbJYjxGhZjGx
x4We0pTNh4LlTBM0XHrMDbYV2nlGBVPnJdTOeS3bairVMvy7quDXyQ3kzUKI1oPg
u1IFEBEV1bIR9JwIFh5d42IrEf9fwdnCA8VifL3FOiAMs7Zs5GfXeWpcwCjy6cA4
JC9hBWaMaYBdxzGbeLPrQ4H4KyEdJ2VpMBFTR1UpUSRz7uMRwZXJDlPxFtNteBT3
DwNxI346otNz2cwnMEoY2XUWuRSHkQe9xocORD1ACC/Wq28ESHrdGkzMu5BPEGC5
z/H232aKMCi/We6YPk7rV3IKtDqRG6sej2Jtb2l4xTHCZdTcXPwvI6aSYy4I4aYk
vdmGYE7FgOLv55OVlqWfsZVvTduq1XBkOiOXZlDucQUj6a1/meIzpxH3id9KX2i0
dgs7JCjXwH/0hWDrXuh/Pw1PyS4avLwBo+Yc/L6nlgsS8EPEmNKd1JWvu8duvZ/Z
G5MQOAZcFlkh9pYqCrzTqKsRzbuPqHa0b3pDN/arVDy+zdj5uZn4c6Q8dkiRcO2O
G10Iod3Hr6FT/3JUEVknKjRRMWrhsGHkv0Ijbhzu7K1AfEF8WRW4ZC1K/3oDQTK8
Qns6mAmprm5uxJrK/ShT/eHGBLE5ecabFcI51tYj4HsmhlmTdGxBtcpxQLw3RgIu
MtTRicG/9sbf73faqg3bQRtU3s1LtJC9POMHvLuJOmv1LMIYfJlQp6/uToBQNH2m
uCzqLnEzqiGizk4TusHXVCL1MZi27fmBSp/e2vgHowqHzqMHclI0q4+Dms7vNPcY
3PLg4HOHd/HWsXxDc7qBiM/ZpbPIwF9Gaxb2OFQdkGdKVsVPPkTFLcVvevaqhALu
7yCrilHUqpDblOTAxeYGZpFYOPnttcAL+YxNjXLOKEHqtTL+NnQScG94PG94Woke
pUom41pALjc/9QEsw9m2v8ctxU1/yBJuIDPs3jyYPZAxEOXjNuRe5Oeu7719HBVH
VfDJEFMmBFlAa4xjNqm7PDA5KndOoFf845rxJx7pjTlnpbViUwRz+1q4xHWI5COm
rwUpaBOfFEF4nIcufDSGQTzzyBvK6pCJAcBQRAfqgxCBrpEKjCqZ0LjS6I9ruskR
e7y4jPjuZQU9SikVKTYaEAIILza/q2EJ0vV0CJQOMWGPD9JFbFsWHGDfE5zBPKee
KfmVLqvQwzL5ImwZ885JKwsjAJOu9hHqU6g/hbV4q09Rli3VKBUTCeICaw4k66zI
SBRYNZhDQ/UQcsQXusFzh4lH/OUWkY1S6m2q7Bn14YF67c63eACdbfcyIgj2ZG88
GDWWWYrhiYmqNA8CczzdSJYoEzd+mQAqumf8Rc+x5LJoxmoqtAWqxuuzwyoENe9z
w6iYP0xIgJnRXSGDEGzTnMA/eKkVSVe3OadHgN/Z3aAbqQbvma2AlB0pA+2/0/ND
q3y60FgiuaI5v0V0xs9l1aFnE0oMfLZ8d5gc70JM8Bku2rW6ICkUzvSWldlxrnIA
Gvb2N+grVI38yHnGGVKxjkjuOBry0utrgF4XBeICkmXC/6sAshjgja0n+WKa8TLp
8iZJPC/BSEabTvtYl5gY17IUXThDhQo4bMFO1hkoeuRFB0N0tgzlWTGajealtWBE
KGHb89J1+ljgajVhhQf86yOhIf6HFzEtRUau5stUfLdkSczd4emDHgI9FgqaYTZi
6IpzC3XVYgBn+5xHkMFVhVg1jQO8k46VOSX5wXwN35UQbfbHoK9Sxzpwe3eNK9VG
56YoJE8IMUxCZOihRWCX02fTQ3Uv9kC402S0m7DQL+9jrp4JSEe4cNPvz92Y5RIw
UFRPfrBHps0jsudhX0su2Nryx5EQdGr8+eua/gYikwSVkj0UFvPAXzJAlxss/7Sa
ZXe2mDNVlQiK1jirGa/Iu8tEHjfYw7BY8CV1PByd8Ib+7Hh/yQhd6BrwUbJSJirM
cttctwyuug4rtoI6S7je5xBwfcn+z24IBwLqaHNAsg5Uz4pPMANeU07UDTjQdnyt
8IqxYP3y768Y/JOhklRNoYo9upwH0GoG3Uvs1gM4atRb8aophpoGbKDjkggQl/2S
vDaWpwmbUyniefSOFz0bRdYNPGdY8y92PpfRg6P0YOeq2zM3vI/HExBHbBxFpWMX
Om1sdkmLU0IG9r1Aj6SUS36ncjejcCJMia7wJnpSrgo+H3AWPU+03aBqo9SeC8Dr
ByzEcfGJFLP5gKaN+uevdXQs6d9t5D/kyXXTJgW9VJG1ejC9uCzJbQmfLRKaqL7T
I+nDkin7/d7yPvovM5WDwfm86UM4f1fYgGfrseAVV5GcBF9GL3/XGoGWvDBxJPw0
Aw5tX425HqyjKHEa0PAA/FAQb91DeNMmDiZS9opNd9k8XaZ8xjlaCWPT+QQOpdfS
psxEYAK02Lif0BWrx8ez9xmn6CO6s0x6SrXoxUx+r3T+JTJQ6AS5jefsSbvFu86Z
fxFXa/iS3ESmQM4JgLLSf7IzQnPwEPqsno4j9mpm3AtI5cDc0i3OqcoyH6yDzjGg
hETZ2vi1DRnaskdyth3mL45tP9uCsFIhBdZgkcs7edbDVtEHoZ2JmEqUZmHawahT
4Dxg0b0lHtNqVTv6WcAuZUYT4rR6LXJZuhn4Nost2g4MlrFb/drzCRNEeuk8IwFm
/owgvgsbde7wuI5JFYpeWVHKSfx+fuxDqAgdH4fSDmM1r9MCq5CSmNM/xRMeNVZQ
Rztr6X8nsrzpmTuq3ctKcM9owbY0ZQtKbhMCW7qSoHQOvUujNwcA1rmvOabWk9oe
rnohYiusLz8dX+cBMo0QyKclDkpcuHFYDaFDCuBSDdY0FiXOORc7GSRF40WvN0K1
FUfF8MmxqrzOGbVFhjkX0jorauRrXX859CGIIdeUDW4Lk743DvZNwXh7UCTbepQJ
FP9NhZ2qbaCuTfppGsaUueLltg0rT1BA6lk1+0txxv7GkwXf0AxF2LhdtQDBNhvn
27j6EhMCjP1X1cZLIV4APsmZqsffiOiemHjarFZ2rYp5rzgFR9cAD1C6AJpZ6g+f
kPvcOS778F0JnPejdF0xP/K3s26m3L7PNI+PS83+QgisIXTac7sbheeQwZ0YNND0
VMwOuOlaenLBPg6kZouqUtdjGswJgqnUBB60AihDAZkMExw7b6IH9xKP3Va3IV9x
KIAKeiSpcNqPN3g5p0fK8D9jHVSw/R5nZEOfpDK8deqRwPmAjXDMnK9Kz1lIzlxB
TvwLxMUpiEp3PXBlLHhFyRewaGdT7V+nSm6ilf1wxKxfPN+b1mtASCjEcj5TiUWL
wmSn+xA845gbkOczppbzyGZ3xKdEe8kTEqvNS7P52qLcLOVfJXV3rxW9VhDq7MTm
ONs6q3Zy294f1uyA8syVAJP2iVI3ZqujAJMKKnUcAnXrUDpaTwqEo6Orkds+YJ3o
JT1uljskisfWpzYkpk5zGm7zlCDmBxUr7dOf3OtRTwiKkK2bHZWFmnxHKkmUwSLc
M+jq3WWtmRJK3SSii7Vj7ljYBJ9PHDaJywNI/AzKRkeDuuVsH/BgLXppyoZsMd/J
XpMd5wMdPyszNLs8IRWj6jZ8DCfHWjj1hXG75COsq/UfWbdawof3skpWFfjXOy4h
+bl4ISr/mXLd7hK72RXnuCtrzp7ZcpVa+ijlO2M9SQIiPoaGIDqMPQx3fdPbHl1q
WdA56fW7rHOVj+TKb73QMuo+QNYu6vBErhavugtcfj2SXAmZJp9ap/KSBTgtHM/z
IdXfXbVttwdilQ5dflkRCrnBFLyeuqJTu6MzzNV90b3bx/2JspoXmr2dxnno6sEM
yAclUUHcZGmoHa1jfSPWpG6gZhuxkgyW92r5R0evmwrSdIUTCy9pDqf7u3ZpGY6u
GsRevLAQY6aHNDSXc7Y/JPtPTdBTL4p2WhSh0DCAq6HnsSQnjv0i5e81HqHWJ3jz
rO7V/GkaeNHo3Q7/5eSZTh6qDfTuXeUQSoW8HDDxGG8w3Dyn+Z72R0tMwXev4HeO
gTNsASP8RBPHzpaPr0WiK6ByKNljjgbQ+BbXii7rkcRonn11ykhwracerTJ7E3xZ
AGHsBA58KUiqQeXLRr9kM4CXJ+ryyJUwoYegTfnKC7Fgz9bYiWLcM+a1Qs8WQXPE
KC6C4sCag/h0+OObTVsnbQZjPBuMJSVHn8iPmfkPS8eGxepX8De5STVXWbu+Xt+j
NsMRyn6IgDioL1rrm6FwmZxrQytvAhLv5CiB7i8Abp9HbkiAXNzA4R6J7Qi4bJ6g
5owDv6MCMVD5bqBT/oAUUrCbW31ZyL3baB4UDb2YlLAHapsMntECXWWGZwPHjN1y
NFZcEYeZfyRu66as4ciKVyqFZS0OQIRqnkJdPBsXZBoy+R3QzZFNOZW73mnMUpdW
9+qbdLdp4j9x9j5Dzew6diLd9crQc0gYoQobuCzZ2pYjBROYDQu5lybEvQ2nZU3z
a7lKFfcx7lKzagX2LOlxY38uV97VY36fCUC7xyimXJ4tLJuauQdvKhsOvvI/efM+
m4nyx0gDfW6jtWXIgdc/RXSXFFHhAQtluc/eXbywG+Wb12hsN5/sEztA6fNevNyC
hLP0JjIwawMZxOdVBo3EYbrYCB8A2s69QEV/VKFl4UanRCdrf3VipEZ4CQt9LqKF
JCaJn4Yg5jFi2dJKzYH0RVURxGvVekVvUsqZVZKi8XMA5cj5NlmQUClKZAoUy4EH
S/CkV1lZZksQeI9PHa5LHhCijZmvWHA3gExIHRlSAaKtF5IZZHf+V6g7hwxtAFYp
IY4nMbcTusGTkvyfQ8t8UKOgIgZwsj8ZEksnWV7yRPbWywCrg84OOruwq/TWYmG9
BG9p6MsxWlkkPFUoLOoJaKJ85c7BmqR0C3cdYVduWJoTS+EQiZHiguzaVVw1+rgH
lFtTbO1a0keUvjhs/irA4xOeA2NrT5CHv3Ib9sD+jsJCxlX05GfL5iyqHLPzZWO1
QoyJskupDqjV8la5yen7sXvaHBJrIosbihDI6Ngl/Fv92vdk8cjs/tzjoc6fpVJE
8qXjjv9j3IQ3NSWG4Bzn+I/t6OkG/a3KQgd2KtJ9BW5r/3hZq0lLI+djh8V/bOMY
nupfqZBE1aXH1PZt3+bflaoxcxu2ZyGNnHcy76x/qqI6vY1ZLArWYlFCWFavkVvP
t6CLSTU8braq20ChtdYUpsRKHcSFyhYoCvm4+JQvhCZLBEIjl6PRlDt9Nl7jLs/6
bKLIRusp+5CWYISKsdO0AWo5niOGUn0vOPDJGqrelWyZlSsfVReOhzghW3233O4b
9OhDclifUYwTyaIydN7aWxruepMkIJPTRDI95BjAySSXpFb7CCZFRHvEAnTKfXLb
c2CnbNbHbz9aYj0zcY30gzHz2UZhn/UyjnND4sv7EZ05XAOFfbRGOGziEe8Hlsut
Gqb5jrX/HMaWsCj9zWWLFG3WA8Xz9oDjqzkKZbVm4ng1vgLhsUhathOI6bELqev9
XCmsnBMzb6CwuxbQDpLtlA58YogVYNolPBtblyKHFsue6/w8XhT4gHAb/G4zH3k2
1Ln/3uBXB3Zq4fkVyPVabmI5ZLa2o2ejk9KC0IwnUVQ9J2JSSgh5T+VOh1k8oNgw
JaPJ1VxVoxqbt357qcHNXFqrGxC3PdHUxUqVqpvmnW9/BDzvAV335U3Tp7AOIqep
ui/BI4ELeeO5U82AmbvPA2M8FSIGxnFzh6i4hOyBnCjhbJybPom3Gq77H4sVNaK2
YX7ofeijyoAb0yzIKrHdo7mbQLuoZJ6yF1+rAf5gDgANXDahEf0Oslcvgrz1Z+ij
VBJVJ/48/zCySjqA6R41cel1BvTx9pGajoBP7MksbOIao2hJe7U4RG3ZLtEjxo2y
1b47krbcmjYFNWv/PD1xu+RLkWUsNt81pqgTI1nbwoCUi4XYkWiJZDqqoEq5SnxQ
XNvLJooEMBEcIUi7S+r93B3jXaJqknTdBWPIx6LGpr+pHw0Pls8hxonrgA7ZwTsv
n23PjY44++Cj4s2oZcDYoRol9pqDmFojU8R5QCI1kd+lkSHa7FZxv+ngm5D0VXcV
TO3SCqq/pFoe5wIan7cmWf3bc9zhwTZxMt/ZWW/5/s+MYKGNVU3CJ4HWSA7sL6Sy
oTTvoLwqrC21KcA78Ifv4v6A5APjQ6XXPAaHUtZdpAA4g7dllWJpxEpuxhfaVbIM
eg7ZZVssMBHGb83VMDfI75pRZ3Pmgbz4/8XntqwPIwOFU6W+9C0or6pOUXL0MyWq
hiiL1PdZqjjiYSrg0WwBTEiYBj0ZcXQUtxEgUFI5P/irWak9x++4b9NK+xb0Goay
I9hQYeJJOHvC25sC2ctKgDlzRi1ZCcOooQxlmthA/M+uNKmGR3QihD4LucE0Xn7t
M+ZxJ/AwiLsPnBYGkaCw+Cb+drOt42wY6XvbZZ9WqzXXDIQfEKsyG7a9sNLKrRI+
/jvmxK7nUmZOAO0/HaHcy++fCFgmboWryP10XW5Ws2LuUyGBQbphkt5pKNA0QTiK
s0W3aoLGYpbOk4J3rg/7RwE8J6yCo9usWo77oc+GG/a7r15Ae13D0rLi4UitJ3N+
CfBxM4Da0RReXNx/XI/vLuC0sDsUTMjYjzlHm9nQt5qjozWJbyBvIPYtDnrG/d9b
44YhvvUGvaAHS2EGSPzAhdNtMAquU9YDR4M0kw6UeDU2i6BuSfWbcgL9k2bLRi5+
J0/mMapNrVRxj/waFljMfB9wbeQjrAZOHxV8iG4eJsDjyPmMsyF6yEgGXjZGlsgg
BkIGsJWQKKRqckTZXUw3kwtvjFxiVXfTFxS1uN84L0uDU8a25pIUpxQRAL1e9uKA
fBRE5uHkBnQeO6D45Y0HhNwhIwuYnQ7Duex8bCNuMjH/0LYzNPpWFG9z0Hbm+jYD
EvBwZv674wmr2gLIOOno1XMWK4NOHgxygqRd/mavIqSA9T+bvSvk6XSSitZFqeYk
iSC83D0uOlTfMavNsWRhSuJxbz/6uJTWGcCokHRS7GD3szXJ234HGwYCl4IUYgyM
UT4vgYKQGBpI9Nga9lU7linzkMbM8BryursBOZ6jWgy6WHg/1mFJ4d74n7QMJZmv
M2fnIyJ7KmBO2UkOd6rklbkV0np4n64mYN4Kc1QgO08QzMIb1+LbpBEwR9aGuRNi
2Tn/+NenKAhEz4t6M2VP8EcW25Tghhb0Uemy5FPuIHTz5jrDlR6IOkexa5rh3dK7
Qj5B99WVGZy0uAGNnU9NdPhss0wYGjgcGZfvZcwcus+6GxwJgCYAhx5UVjeLjHi/
3cOyFndsmaGZsA4JJXQkfiiFXDEGt8b9TPpFEJZxGuii97KXeyP9FANKONYGI9pp
8UdtkFrB3eINmvIKnQ/QTUwlPUOSybhdGd54yumOlVOrjONM8/renJ6et0xSefLy
ErdCee3TALu+ipQJ1SXkgI1eaikU4QEQ6kOIc6oFRjBuDGaEdkPsEhZJrAcjB6my
JOdD9XIw1wCG+vWJvzzZLHLglq9bBNt/gXj8AwGC5Q0DK1HVVUiQpAaFbAgPx8Mn
vWTo3ahzBrKLl+9RaerlnrRYTc1wyq6x35mbqkUWw13ZbcChIOlYLIjSOco/53Mm
IC4Lpm+OLSr3dhD6MF4RVeanWqN56AFytqaony91K3l6UWv/imVYG2qMtkPE7WbW
9A9E0nAQRgIYOHjkfqx2Nzh0sZxfSNdy8EEfs1Al86gF3+YggnEHAwPMZpSFy0g3
KBp4f6YjCFHTWO6GU9KVZG6F1E65D4ytFS0aJwoFc9WL0tknbCMwBZ/3snjcVbfw
naf9MvdCtzTZtJ2WkmbTPXJBgNSgTQ3BmoxoZv63ILv1eS3BAIPHUZvAiNHs3uy7
qEpj1YDHadW/D0qlhBF6ZLU6lE2p9ZC+K2yHkArUvQh2APUfjUTDPyD/XQcGKd5f
E2JCk4P9AeAzvD1URR2gGY0cZFb40pCGrL/wIKq8fG6f7FfGw/64YEK3aJ37pH3L
12x7msXwZ7mp4tYSGsyIVl0dFfD6nDKy1JH9MSZ8gn1ebAr8BSVo9tPfYACYsZ91
aoiDfPKcos2T76LNWnMa/UfrrPBLXxcpCgvteiuyWd/miMDkxOm63Cj6GWRPSVKP
UCu2c2oYyaJLp1R0MDlhq4MTBxnvIKmZP7BYdOb+KlFaRarvuou4Mq5J/bltj05K
iBuligPabGgWJYHVyzbPglRjorjfLbnp/vzqF6GdfeBAlOMX0g5wxiCaYDGdfg4v
/ZKyTEcreZGHfaii06Za5Hf/7nV/O0skdAB/dyNCzNlA/lbggbcjjAbndL0/fwmB
wifyYWsUmDJ3EpWnO/nN9kvHudxYROKkrWaw4w02A1Ek5frTGKnRjEfbfQf1RHs9
bzHLvMGh6+WjPkOSSZpIVfNtOc/VMkkb/lL4v6yxDR/T3Lp1NKHk5k3mP8/cpU5X
ddY+W+ZBa2r8uOIG48FuspGKWrlhArjmDHKCQLjgRWI03L7MX/e9FkU5sn9MPM7V
i+OvoK9WiDuQeMXsnwfM0H0smpky4p8i2yUAvDa9Ekv9UecQKOz1QT8aLr8FK40q
hZpjr/DJecciXvxkVxSkGs8HdWUJljFwYb5IJd4MiWxh8IdbBjDcSTDopKZoBZqn
zEvxiehAXlwLnXt96eOmX5XJkChrtX1TFmbMgKs5CPh1zpY5zNHKyghaaB5gmUTB
0SnxPtHgR1Z73ZtXI0hJOcEE+SLYOADnkl3j+2A9LtOQXy6+gQXxFdotNwpdC/tp
w9Q4LcdyMcd6TQS0rXYCy9hDhGQddNZmcW4KO7Nm2qBAMgSzudUX5XG5htQZfCM4
uSQrnYPl3hZuGAKDJqKlZI0LZ5KrjlGomA9M/nkxBHRD/u6pTmHLHWRe0F4hALsY
zUt9v7ann1NEybCwbdu0hH+ozIbuEj9qa6OIGQtsV6a9BuAamcunteTvM5YH9xTG
EsYZ4J3GeMA9ecKq0vF/vVtKQshE5pjhfIr2CjL68JErCjgx++uUdhIhmPsYnzRS
oySVlp+yaLmQvy0BNRHHER1FW3311yhyThRh3xautKtBRkkaqJRI7nWyXWcau27x
ylzzAU3HY0DbeG4Ehtl9JjRtGIgfg5DwOFprklrKZ5OucPEIA8VpeBljvjCm191b
cnR27pzARMYE3bxC0a6xS7i12CCQRywbx/c1wRjgzK98DxvTEUiYLsaMNn1c21Y/
hZbWU+i2J0LS7dxO7b2kz9t5P1D9OO79Fipv6EtD2uAUD0/orGz8/f5eAYX7jJjy
2uyABNyfghHVg9k0rw0bM1cwV/CGSar+IGToBJSCMdvZjuMz7+9yt7Sf5kzzvYMt
Dvwpp3GIHNQ1pErIbBu75InGBtnjten4nJ4aMoFHDBzY5w/9MgPgGrOa1N3S3cf1
WONm41uLoAMgvRmk4XNe1BBE4RQgS2BU7qnrPhqkLofYdbyRET5pWbRrMJAhV6rf
+iHCz/EhAklbKyqdIP2Avd/wuI2RTVG2p5N8I/5iSRQf7BjRduMSdhp6DPLXiYv9
AlTMXkUvEKgMCSuyLMaTN2kWbIeCPrbuTOAowEvZSCpkxtBthl1zwdko9XsrQRrs
kj0AwaZAjEKtR/zy542U33+RqMvsVh5h2Fo7IEsqMewFBZTQsLLDshU78ydG+sCq
sRPTcK/e7FN2NYwMHDuF0ToEz/EhOZdLYhycLQkt0zKYHQlfBlI3/Ucl54q1IBeq
NhMi9NOm1WaSAltTABDZINZMAnQIocH+pZ8IB9W5SIvqULddDksPT5QlnIzxzALw
4nrVUJOEpGOYGHOARtDa/laVUfMm/Stm3kD9KTH34ykLZYkGd9YMi22hfk3/LvLq
iapzwvDoqfqvutGdz5EjC0aKBpwinkGv0tTn0fdrKUtWZBBqWzXfgCCPvp9SYFwk
vY4sOXbPuxxYAkBG17I7R6NCSPhjEPj+Y+i1otYbP9YMJY2rS4p5kmy+DQxzEFRW
O6oCHPRgFqPsoInnk72IPLItCmo40ObjXXqNIj5W81sUd7p5SsMU0w1W4c9FJKHd
cjoHP2MG5zOvR98N38UyOCR+Kr3VERV+PzNSUbpqY6AN6kOE8YrnoLvZ8FvX0pwU
JcDm2RyZnSD+4K6e3/Omft/2DCNcfelrSVRWv6L1cS4PsC7vV3xk3BF1iQo8DVls
lI3j+9uwyhvZAgj9M5BvxWgYFdRgXlHFGWo+Oglv7T874fwb4BzoK9JgF1gvpDke
SNPNPv4sOkk1l8c0cGrYvkB/BA8Xsj2GPQnsZ1NoTrJ0awjd1IIKjgPudRdslmTj
YZJe3enYdUOBsMH+XGdoLDhlRqMkCLD5DtXBxvBrEJOWXCgNMHrlB0oKxhbs/4ck
gSyW5q3oR9Zlq9s9gUfZSRvoPb1dT4LmGLDEEZk04UydWOeNtEt6MeM4TMavqAc8
NyvAqU0O0L9Rt1B13IkszKzhF0DqlGmrPvuBhdD8TMQWIbv9C0yYEOX0mFYnTtHX
u6Z8v9Oh4MBt3xJPJZK4XxwyOkltv10Qi742YQRdpcvKyO4yVSC1dOYETGCZ/czh
6iPV23BhPXlrkguNPS/MjPepVVnQ7MKA54a027NVmCRi013zn50zqOBIEOLeKk10
91ChG2ryvGRemzT+ZMJmKEbfea6IbmgIfpOeljLdGynsPUReUiByl//egngFAJyy
AVdlA/TS45x0m6sNd56m1K7YNxCFqZnQ0WNN/BdhALkyY+3ohMiipKE2/GdMmvaX
arUhsd/pA1H0cR4CMsbNMmnMmbxVt6p0Tvh+lMKHZmc8lAVhblp9s0o8YHTkA1Vf
rNk3YVoc+EJsGrtzRQ2fVtswsvegAthYvzr5QL7YeDjMfM6Ydl7ykrNcP+IgmoTD
jg/mmaOiyFigGSG+AIOhy5F6/gWJV4Siv39it0XPeTqMmtut7KS0265DOM++FQBB
nhr2MrdmxhOvZuDP73vlscJN+DhTzFSXB+I59ysG2x0ReOO/dyStuCz3iefCJM1I
iZOWTp39PQn0c674GQWYqsGcLFwxh9npNK+1ax9jeGGW1LRMCyhpBeslhPq78YqY
Qn46I1uc1h2E4WRhmESWQqsJb0+D0nSPsjXDU5mRS9lM3ZezU/4SYLqAQi40Uid8
+fSrMWBdfwKWrnfl6rEJceoqjjzc1x45ljMZ3atRXlwoBhtLRPTVwEvxXgKeafIo
mhynD5Jp9lmkXCU35V2RN88mq0z9YS2JALIi0DJ1XTbV/OoZlJ/VtU7kDb1zeXaG
aTVWiR1wDBnH5lypj/i9NjxfkuodTXef7oBlKBX5kKfRNOcbZtZ6KwOUbAYRqTQn
mTYg5rPsh4C0LOKGKnioqcFjRh5yWYkhOY69ZYC7+mgUVWYCfeGCZk5nzciMBex3
O7hY1twxUPQozJC4de6s30Em4odGGH5rViEpbmGYYTAhvx4s/hPKHaEhMtccOcs1
bStwPAcRFxNF85RisRlKgEG3vTvDlP0UZvdiiNh3Q6Kccq4ympTULm9fJ056E1bW
2NDCTk6IwEpfh0Repz4b/5LBmDAR52ilajWnLF0cQO1QX8FCv/XfiGix236p91rz
Omt7mGOD+pQO49JmZZc5nmPRbX45UAJM/JpS+UVLkOUFCSkry9MubJdJkFM2iQ8U
4a21zBrnJ1E7APZe+2DWBjJZGTYxOU/9aDB7QTAC7fQNbzhmuR0bqYdxgleyTaMV
u6hFyBOH2CrJpMTCqbYAyH9ioe6Kt7cnA+mbsN8WvLZjj4AHxpXaiEqak+P45bEg
ZmCJCdciNd6hbKN4jNFSFZbN/eEMlK6AC6pgZhWJAed3nYmt0mFqYUEJyUkQ7qlj
yglfbYv1heerfG1sS0mMrQIabB7Ijw+fHeatb3PFkz6+FYDBmupeGaQyyw/NDrSR
BEVpeIszWKXL7UKr1qjgbqkwQIuTCHm+w2tHViut7cDKMYS/k8Cvp/kki4pj41kp
hUeBeLK4A48695OWcLOPe9HP1IvuLckNck7o1xHkseEB4aLVYJlexMzy14rfV7qA
QbNcLuY29eYlPtrT1h/16GXoyAzIwLeHPxjXv4vCaeeD/40pTJgLc9Iw7Hqm17YZ
M/waDHLpZmJV+JEt/Z9brmi/T3MqlfN/ueB9CL9g9hGQcfhgufwyPXm+bciIQUj1
zwakABrfZ9Lk0QPDQTM5jy0VIxkk/VOIIrkwCkAPr/rDtpFYoRdUFdOoX74ZraJc
VOB6NAGK+QSZr987/BJ/SOqJwd6oH5hcxp5GHrQJAJSO8P3JGSBCPh0ybMBBdwyj
OaSvQ/0QdNekDK0H3gvDvKJb2qeAWa4dg0nIromZiwcy9At2LAWBmK5iDWZbpLvs
wdxdF00n/YcS3oRWATiE3mJV2kTeUnOYOQwq1ZPQLVrUhxu6haDUlHys5dl85nut
5Tik3Dj1zojBVaHutM+CfQo8DQgbzNWMwZ79xp1Bnv6+4N/qwMGKzQqkVhev1YA+
2gWDn5sPr/236wEW7mduwmPOt8Ft+nJf9MwSC5QdmBkX+rN+zIMO85BicAHBcSBg
JsdJF0M4Q37QsnbnjS5UMlDOb+G9wrs3yrW1+dSUW8rvvhKS20d+a97B6LtSzxok
ECbdNLCUqpf3iHKFZ9SZSPXqPnlBtCqXmTQ+EmsJdOlrfLD6J8kL0o2ALnIlewv9
49ajYwaeXOiVWa9U2laJjEO9kDTufJpcIwv2cH3sV2j/vvl65wxTG2LD81yoilDY
pKF27WXv6X7iAZIV4fiGmD28MeCbX9AQlkhSb4nL4XqfIRueHYzi1WQXfqrr/5Bw
ofOD0ISXlGA0x+L62PW2VfEqgTXKtz71rjk9A6JZzHl4AzSbRGG7RwAyf66ZiLO8
t4ClHyfnxuKRHh719MX1jKfVxYApKdkWXo3Rg7chF8GLU5KW67LfKq9sR9lrM1t3
vVOmPS50MVCsi3UicH6FD9wXz+UU8zfs3x5TCekhkbiMGxT7HgzUAM8MT8aKkbLw
GXVXg8Bm3vN+qt3HFKSi/c9gpPEI+3dtYHInUPp7tC2M68NJ/wusKWkyV4Y+0nRz
GHy8cw6VUCgvGVGGLcc4JZlk1vIjedMl5i9wt82xnERiwZ8QZoZXJP6yUDH79ove
wGKyMEgjyRsyoq57oJOVCaBSOXNbgYzswSZki7IeL8jmdG5tLR2Zlbvm2neWQIzG
+oiny/Rg1PoW7PsJrxrbMTsnZFnEUXlnMd8hZAMcnyAm0eTgqus2aXgKmPH2g8JY
uD/9k6RWJn+slVx9eAwbvEjiwwUBiU08zy4BE1NyhxlLb6HmFToN0guBR/KJ7mhF
I9+zY8r1oWNi5V/1R3IS1RMTBiKxM+yZOecfADYoTWC+o2UBhXAMOPvDhVuYo06/
dDNG8IYMtZw3yHNl0fy2IWVC2cE+eg7ihZiEApS1L5hqFf8kyQalWl06sZ58Wkr2
3GSboS71Mzt48o7ZOlhUNfFTows6dgi05W6Hys63NBtS2kJIKAPFUdBnS1q8TFH3
x+g7jZQ4T+9qnd8QDMSCg+yK0XwQmhkH3Z5RJrviXt+4aRtOOsh2ejiivm99ItKf
KJ70VHBK5twirOJOchyjkPjvplN4Rtw56KhIvCl3Wujvvx2McfbOUSmvnX8A6xLd
DV6BzyD2lryZN+by3G5XgvxLf+2WKlTPQWorpcCTJgE8jNbfDHe8DH/jgbGbyDNq
cfagfWGdeSmruIwvjLFcPNuRuNvIXz0TGHUuf3LmpmD2fgRiiXRCPIo03hQ+aTnt
3TEfgn/+kfDn8X2sT/iBidm/kn8ubBOezBppwk4qf1s5NsmQVDG+pg6OxgvtkRjS
pUAr/icOMZWz/SqOJv9EG9e0SiuKUBqhn5KcUkNYJMeGPRqKYQIPEA8tkw/SkNla
D8kryu+In6FXPMJvDX2cVD9Qc4bOmuX2cC+GZm8YOuuOdryM/WhMqYFDKe61DazI
loQy2dQ5tS+a3nZDZ0WmY8cY4XyaMFMafEwNg6PiC7Kggk08FQODSzIngXoGs7Xr
oSxu9EhAAqvy8lDl17jBIU+emBmMTtytpBFoVM6Ay+SKW3aBFm4sG76ghyDnTEXu
ICzlYiqQsCQWn+5YxiylNAKli9hLHjFgL2MXjr55cLfAXjs9Sn6p7qRRusJq0/HU
Kpa2ilGBarKFPw1v/440C+88QJwSKubjFV6sCNyutVTtQ+foSHFg0mYEKxwMQNxa
R0BYsN7W8dv5Paz0kdh/ajb45GkTywo6epqKJS+Ld2YrUYstd+UKJPae07zCcC+j
ULd2RAhYfZYwq7UWSddG2pMswv0eMdxmDQqm5GHWntZtJvZB9ops9HJi//+X6jvJ
6tMZkHbz13b2e2+ViwkZwyebASIH4CtLW5yXM32btXBE2lPb+xEDDchZptHJ1q6V
HpPlTNPLREYLHdfjrxqGTuGx1cZAcYVwKJ6oj+8IvSGkWK2bqRhgkuHfbF+sfQRL
v6Heq1QBPsBBXgyO0bx6WgGUvzzdK25qtYBSfAKC6c1nabRyUJiax9JM4PspQDKc
lE5uZO1HgZxqMxjpXmIvl7mRM2Mi5QbUwIu2sUwzQQsBIMcw01+lXB/81l01nn3k
wlb5O2MZEXqGJFkP+RFlnFKvMLmoFNYX66K+HAxpCpd+8OHbF3LGQNWA/xfie62W
prKqnD781OKPcxyn8m+vmDb20Vwfd3IyBRRfRx/TfNaKd2Egm5P9LppuQUtzICfn
99ed0mXKunqasfoArDKxO5SWPoI1+gRxdjOPi1B5Gxr/LoWhOFWwykMxhsG5VplI
JCtcFpVJY3TGZo2pRwFH0eALssS638GNc99iR31S6eIfn/59LzDWUmpDDYqlsqup
WjP2DysEliHcEOH39Af9tVwLfwO2KsnajiQETPS07hM7fmM55KEB62VR1ojzQjT9
FdMpdwKuh9lz8p8qC01pQRpXtVLIjMbnh3ixlKOdX0DUtCfeyqBRyyan9Aed/An3
AdyFSwNc3l00xf1t5Qpf0Q2W0r5LT9qA549fs8MwdBjBPKfrV4GaVfX4aB00JUv9
2Af3YnxnaqyivbZ/y750ZLdtDFUAbZ0HmUpEDAlqui+YUWuth49u/QBF8P8OoGwL
l8B9DEkf2kWd+ZYWn9yUrXl6qOdRGRWzwnYzMjADLMhQgBCEpA9vDOEQsSxFPStL
yeWI+gSxIsBbcqnUhTgL5E4zvVDHpYsO5a7rmtuw914DvpTHPI0Us4lOlL2eboSi
W4nB5tB5TGlDeu+AhjF0KdgDodEJi7c2M4Ka6TcMqc/zQKxzmJFmDKkcS+dMShZp
NI9rR7XmK+wAem0mR/hIodOp8n/tgPFnOSnJx2MSZ+RXokIIpjQxHsDxJ7FgbgFb
gXJ9Ry8C62LYIzDszfW1DYDoZrC47DKNNfUIrXsVd0CGk2ijSg5CWpNTV/6lEIM7
yV1CRql+hOqQjR5pUziQJGwqTfV39bgYgVqAskz70H5RvsWe3CzvwZaBpVe0zewN
2c18qoy2sTwedB0uxKCto1AiAGoigEQB7+p/DH0OBko7y1zHyD54GVMm6c6m/Uae
yR6q+ISyf28BVNQ85Tdn1ANvVhmt5FUZ5EWbtL5dDIvpZsrMNZVYL4R95UQX3Ts5
z3/7Qw0On6nRQiFJcHZjOm48eSGZl9iz9a6gedXZkmGlf6tgokAr6rPP5fcNj7MB
VjxtOtv4rYMXNzTHcUOkGnoTpgxnSo7Zjdxv5tQfErrFgmhiJwGCUG/qvfdq/9yT
lUjryfkbVP72hZtOZ4LeKimnPdW1LLV9HNuagF1/sHiHwPlJNQVgjzTFTkYO0rc0
3UYUoQ3ceIdV/d5t24lnmqNT7q3hcr1pJCcx1djqQsQox/88NQDh1voVmRZNOfmD
Eb79MSm2Ou+tUyI/Ipu2tQFHhX1lSn3h+7XjT75EuTRzToKP4oSxYfrirbrKH0RM
MU+d7wofsU+4+Bu6oXkH+wYwpHB30oD17gkfAaQaaqVW4EqoCOYpErWwxNJyTo6O
2nzEZwhQmWWD4VPkzm+LcMPaYB7Y5YT8p8kP8DbwZvkayxGwkRWWAcAIY07xAeYB
3gWHU9WuSYANsLKAHF42r7e27A4ktEhqix55AxRji0sIccRtZBKr1mhTeaUti3uI
obDq2vDQpzDBVo3GA37ZHGb17ocOrAzhx+8fYYCCHOxRGbxQJOMqCCpzcm3aCbef
MC36GqzFXyn/UiEzer771eGAeBBGgtiFXZIs4D71Y6KZ5GfbCPKkGGIuGblPxIqt
oLGE73MWETIQP1KHT0Wa+rX/KK6szoeXf1KeRueeMOufBC08pqoEahIpHhlbcz01
w+8t/gGWMwkwhOEsLGnfcdw4XeLIuyYwbW78uRH1w2qYG4ClJLRXwJIY/MkeKyhw
w7B21eGn5dgFc2I94OqMfgFkp9HWikIMKu5XLoHAwdC5ujgrtyeRSPZotlCmJ4i2
pwJmatkfncFw2vsqq4iicbzRGYTwg5M6ehxrjAt5kBKkrvwba00vfwuXrV8JQvPd
0TvkrsDN+X6QwO2qmpbZSt1RXvdmqw7LUlqfjXCNvov33zhXeoLIGaMnxEKD1Xfx
8ycxOrslJX+iLidg5hUFed7JI5rVgc5FxsGS98pfEj37HSCiWBoUFgpM7/fhiA3p
uB4XF9jwXoYkkLN+Rb85d3Ct9Je7aFVrrwXO8UK0L/z/9N99fD6fimXhaFjLu1qE
nThIpG9v26/F07VQpsN1nEaMftdiqJnt3yiUe653LUC/cMRNFzCYDTMKYW/9+AH6
TGLHR+wHX1pbLGE9zpVaAIrwNnKIG9rCjMA0jfl62p97reP2WI/sgZHkAIz/DGuV
EOwKq+GiphAxewOTZ9nYJVHLoLiS4GYc6ishxo4M+uHbojH8WEWho5AiGo2R6+AY
sQ1WIPJf8eWv0M8JtNlNYC4pCAGfNFypH2DH806MVMyOr+Ni7NB4ecP2Nf1Wz2Oz
gyhNVFmesyDW3gopGLPSyarldXB5G6N05st2G4byyYYoJ2hANjSVgKfzqwSk6BRv
Xnki6ryNXGP2SkJPmOJzEgnUHxzPQn7tppfMVcM6J3oER0Fj5BVf+byvsHdXN1hG
qjdohCOGrD6mcnQKEndSwu7SQnEEt8BN86IV4Jsw03SNPxKbw2reRc84nF73Tu55
BQ07Odqjgz1gOGDtPWh0XpFt8C+oHoL/AmuqftiG9PUEJ5DPpU3gR8KoASmhwyy7
g8qnREzNV67ZL2W/1mZN/X7DbPuRoh1dEdGbdyDfOTUPaHc9Go+pihtZeFtBtpU8
NqyqpcvIuxNzLwVTp+lpoS4mdcDP2iAXwwb9TK9cUlBbHOq+ujFUsOmRsD00eq9S
FM+xUkx5HE9t32CMtwQeKNflXogEPeOpEyIhVbuNDzCYrT0CfM7/hNGaOMvjA+QU
rnA+BaD+L6TtutOswJQpiWCS5Kr15uHaCsjjXSqkDLZviCPGXum1fV2qaLdi4e6w
YTlqyGqBZR6E8h7uZYxPx5Jn1VK1WrjMP4pYywd8mk8B6N992sAfRyjNQdRg76QD
V4GbfUv76aDfN67rIxMHQqSsZvI8QKoQlxd/B1QRAAqhZ9hb3axRxRwVRlpzo369
I7J3FJUM5Tjs4w+h2gUf8QZE4/LvZOoCZckL6XX9ofK4zS8cUACBb1qlMzb3tVhR
kpeWw0hpiBeZQgXPUYIeICJR6rfLBddk/MiNFhhzxsXXI5Xr9hnFrTfLUWAHKnGt
0Sr7FuvPe/Fvb+2zbVWossrd/k9xjf7VIcmM+4x5IJYqboqIrWZjobs4SwPQA2un
pWZ7ESQcBzb5cc0rSReLSjKw31BKpvlpfD4qyCieVPwmNbYAVRa0L6IU/Jf/Wxqt
ZeZ2FWwh+t9DkbkvPAZE6G5X/uqrBHVhEacpGR7y4g14G1UKEpVp4DN7ulCpHlck
OKzFA82uqJIAUQoKOEGed5gHNFGHomvP4Qwban9i5TvH746MNyWUdASO13+tS9T0
6qkpZrOl1e8wicyRz9kZ9zJ7YmNaU/9alHjdkdEwXSbzdWp+gJFGs+vxqQfNLlkZ
NmJLWnF+Tq5dR8lBFiLc2OqNLBQ7VUPPYl8tLR7RbYc0kaX4YPwDIzJJ0W0NXe34
01MkulDXpSztb+bhSfw1QkwVUMbeEDJbqADXx8lxVY+n2phNV7NPcy+eXSZg/aIG
B5/YQrvHxchlJHQ8MmDIuPAQUKVpIqTdt3vSn1JPIWeF5QqzVphTIp4ndkOYvuPy
E37ssP3yZVzSSv6EIBQoxecMpQS+uIQ4nlA3xdMYkdNSlGW+rDID9J2oZChrNA01
a0z++07zqe1RIckF4AtlDMPPTjlxKhFxIXNFJ6qutFi+ccPrFz8OyEq5KgMc1Dhz
azTVGXmSVeny7uNRRPh9gnCQdSLu3Ib8nuQ8tavSY5jKnbXt9aTMvadfF8OoRvxd
mNlm1SWROS7rWWSfaA72xLhs3PDbZqr1NKqOjgl38dsUBWFW1fGZeUvPhcf4uKZp
bG+oeQEI6EkIZQecslyDi4gg2RGVDgwPvmGZis7x5XqAPKqZOoMjvBhVzBjGe5uk
/ojzIsFSiUu8YJp8nconmlqbuC+YJ8xOr0BgEBXL7xu5iY97egbW+pycuCJh+gHn
MtT0paMiWpfV6S9XwCwEu/nLxaZpya0jXwXFPKk5AKFeVqq7l1Xbij+fZwIsb+LE
Pnp55Qy9mtxL6j4axljzagPPOg2P9SMnq1qxJheDywAtBNSQYDfBM853X+oTx1jB
mPUWiXBYWpAUar1P+Q/0P19VArvPwkDX5t0jqg9SgjWEtmhwMVlG6qcMVX/5MA9k
LbAwy+kyzpoddnP46oBqWy7vnPmSUzuLDACszazEgeydxYcuUu4Pgn6xYlxXIk6p
R4tHs71wnvRJqDbUkuHCkHbpEfNmT5M5BbWYjLMRlnOyV5sRfUOM4H8OqREJA3HZ
7W8+Xdspw1HWmup8gRwuIFKb4tdsKx7a2tKnSrxXIv2TWnbrjN9X9PcK1D/vsFov
arZWXdnyw6D62akEFrd/tQTsEG9ZggwBkioBdM75JfN1LnRMUgCHi2j3E4itOf+9
fh3Sf2dAj1rtJENK9c1A5slLEGtqz0kIzfQFIs40RSUJQNTZAYI3fLWHzTJISFmI
WiYy6K/nIob/L7Ez/uJOuUZ+BiOfPEe2YMxK6eBMCt84mtOjacyuK3Z9/pzegZHg
JlWTQ9ieozvsjrlz4kEPQNW7bmiuIklyRAifA8d445k87HRtqCWm+Lss2J3otcGh
s2MkFYYJ1zoMrw+rKIkfoJ6m06Uh4cAkjEx9ZEubg7wwB8lN/UMoAQtMqeyHxDj9
JXdrFbPXxhFjqXGXiip+wZ3KtoD/D7uEyVjpVRN9TPp3sO4h4FR2kaXW5u83CFS7
0aQ3Up7X/MxvTAsl933TZp60rvCUvCGJriMv59za2Sjybtk5gAnrq8U4gi6EQG60
AZs3EHtdnw4A0BMUq8Kx+TIeLD9IW4hrIN4b+e4IPjuU3tDwvLf5LPPV9EGicFb8
uOXjtBZoMaMIFLJ9D39vplEXmwE4ar+Lwnla+reH3RMiKl1u0fRkvuPSN4TXX4No
kFL5BP5JlADljqne34gzcP1w/e9no6NZvar/rkRbkZnqGAPx8v+/I+WoRqcCVV9C
glkvEztIPig0hlYOMJjyvLEZe9aUtCOH/FdW8iCLoBNQjQ0V4OVJF3GtMZVDdAO9
DnwL3zzZcCyL1YLYu2bZd6qV5QK6/+RU+lsgZ9L8v34+IqQP3cqZbOgj2xrwc0f+
h1pZb7iocG6gi9RsCc1dVmM+uGKLlfy/KXc9AMOxcu5S88vEPqpOy/AWRfXCCMIl
s6JEM1WZXP+XzLLKQWWN66YfUtUz9KGMw1zcUvpQOnatF2SJ4aSaxNf/bSVne4EG
VFbTfThtLshdCvev06S+Kmw+EOMehuP5y+/yjjaxK0BTDE+fSnktknyOv3ERDNMI
/kliwKznO481vclDx/s1fn976dQjyMamPza4eXgEo0fc9YOT3sxRCOhdjG5233/f
cLmhfwePti/PwuhSd8DY6JnsFr/3y55KewFP3t2AUIh8HXfZ7SvyTSD+Mkj6twQN
6pm2/uB0L+bl78VRRJAq37iTWqrMMIFhaYhG6RRWsRq7nzjyCq14aq4nsGUqjqsy
Wzl8wFEgKr73KeeMMqJ/RsPbcuXQs1kPPYI1NBGc0WWS6pq0/efDR+D1VF1KzItO
vFChHJi6U8nODdpjy+zki0Y+E2b0Izr2d0hNU7oZATgly/FqHUNU1b+SajmF/Qe1
YPjIGkBQ37rgWOsb+Abn1PwMDfr3Bu0IgCnbcoI+Nmpf2TpHSFsJ+bY/9PnwI9Yo
w2RXh/Mx9OsAr4eglMb6qtP553TVJgL1E1VtvDI5dgfY24Pjn6Vu4YSqfNBJ2lX0
SrOoKcdBgFcPe3+FiSbQh+BIHWnghn0re/6rSsTT4/VkPa9sx50XLO049mNlUIsi
ANlNaiC2+oXCga76JApTvd06HRVqXaokTK24QLo7BGdbJkyg1do2KONrIKWsY8Ui
1t1dr2oSD1xh61xrDLlQVbxAOQ7acm/geZ9/9O/UAC99Kh+X+1JzVTkEb5gHhW2D
Yl9S2jtGnd+0k0pxFYB79qnJ1WsYdiBsl7XJ17LUXz20OnoM3N+DNKpIISi+9GRp
JJme8zjO4bES2gaMrMGG+uzVSMouHx+5lRLQYHjNDvLH3+MCd21rLVrK75ybUGf9
xuDhTyeAZeQeuDUbv/Ugwk1MiM8unXx9GJy+U7BCKL87lsTiRtjcYzghlrEIBK4W
C/xPHEduwpze9kAjroJCqzF0qE+yQ/4y1Iaz4u2jYxCGCHoDmJ4UvInC8/Oage4J
CXjDRqnEyxmMs09PgOC2FQ2TgoZtWAJDaBNB1s+YsCHdhoV3pZBEKdZB3N4/zUxT
maMS+wADmqHpw6Gmmxc2RCJfGHzjbWyS6NdAo0i5r0aOSrsBJdE4V/PjjBSQt85b
Z0PYjmQ3HOqVMSKi2inmLnWsa/dOInhb2yGoYtzHFlmixi0X/6/hSwspmg6jo7Ju
iWjDsISeDzGV7Fe+99VCk40gVYmDJy4s16rYG7KE0j2IrDWrj9cj5fti4AtitYkq
5a0dlLkJjgyUndPyPEl+JoR7PPyy1Z4rlk6f6pcnBkEKh6U8tsue2d/Eh8H9oDpY
I0Uq4lv1Uu+PP6gQ8VBsVqYH+SWE8MlkgbRf7OonGKt0EYo75KNu7XpK+rBNu2Jd
BRGCNZ5br++oapoLHH0M6PXRbscBv9MTi0U28jH4bJMjkDA/KLynE5rMnoXuEekP
7CHdZiXInqKzkBeznMMlPaaddEAoqJtgjLUUSotEwndAl/1gL82zjBnct0GTYIuK
uzbUv/Fxxwwb41GfhXtHb00qkHj4wlpnhQ1Amr2PZXuAAbMKFfRR47FM9DmBRBLc
xIYw+vLYSuvxviV1cUYoHPE7E51BulQvt2Q8Ii3RZI/tNuqZzgQQ4SWB/E0C+bfF
YdoSK70IFS6BCz85Qj/FA1/XXq8XYzcp4LMgweVnWJm37JoMYm1RLkEf1k9vHC0U
0+4tTNbG8Mztpt+LHJBzxLuGToEDk+joHnH/cMVmdlyD/2/oBm121ntcoRZlVJDP
AgSUIyHlFNio1OEGxz6/XTj5D8ZXPEudvEPK/cA3+F0hRShZfoYp8VvlAmmRUsQo
pmPIDbjNhRNbSjwBj7U3k6u3W9zNgV6KEUea9rumLkxp/BaMYlPs/jmAHoxacHeY
H+10I+IemqhwBmJ9txPM/jzNnOLWaR2owcWk9tFTkyddUrg3V611gprLbjP+M93u
c0nbbwn0YZwynOkhquDyFhtjDQHtjzW6Ln6Sr7Rkp92ZKPHSTaj2GN8e3sgiO3Jy
FAN66HA21VzwQUZCd0OIRnnloDYdtLxg7Yml5z52YEqVklXJOlFGZeqmset+BQeR
Zgwl29ZD5O1qGfbOE9hiZwopVpG5Lph5L8q3yGtom9ipBikFTHQSXaog1JgsbCs4
U7RXEtRP8BiwBMbkIwgD23TAktK0m93IrPs8jdUvfYFpqX9o9Uzmxx6lYpa4HLgS
rccDqz3sq1XRDcpXW9NqXVIwBhb4+KVSbXLYDimPsAZ0oK4GeFxmvDXNbKCRSAyK
wgJTJ5N32sy+gPh5voNEqE3WvAQuXxG6GfCmVHc0yNDCgWZu+sUYRXjCdoidE3qp
DPPavfuA+4hqjMzy9V1pfqKkrKXgfrKoktzyy3XRrnrIhDzQpJC0Tj6UOxWXIc5l
Q1iQ1UAbhhaUE9ueW7cy1p/HwRFs9aS0MNPwWyfPqmSiXGsTsZtv6SvQFQUWUCfX
7/iEr214WPGhMNuhRgBXfqpesqNJH+UzX277q9jJIkv8HF05CEQbfvWR7ObM1c9L
e7bneiKNoA6G4ZQVUy19oD20eMDjQqqfDDhGz1oTZ6UJZ451GaBwHGLBVYrLA5Gi
pyHhsn1NWHas/ejRjelaVF+yNbK8r04YrwQhIUPPX7pTPuQJAIW3dCjvYAprodhm
qXOAkF84taMFWe4JOP+ipvOBiw6mxOXOiE6P8IQTQ6ifY5VGkQLyrr5yUmJkPoBp
IHzxXKm0qXuRnKCgr4dbR3qO2zQ93ie3HLGUiyrY2yFjoFue1qgNdtHOlwiO+Cqp
KNvGuZfHZ0oQf9UKJEkj9mMg1r0XNeb561Jx0BwfBcSx7IYhYu/v8HYmpXX3B3S7
5yl8BviIB6GifK+55yYMBB5gEYQlNy4YPxePPmGxTlrkzRdX9cRCsYW9wmUjuYz/
juhIWbhqNG/EJ8HhvvOKVySfetYHLGzHzOATm3n65TPDBI5y552yiDhOg/IsVte3
RlJHPgOxoYbndpkUUnoCkjXBFFV8MboLzKcoJnmRkrMq0QXYtMcxi3bZ3Pxo1ygW
YqiOT6dv5gGxq5EIwaNq4f92BfGm8r430RmWwDzOawxb0GmsRLZZLo65SkWrho6/
lRabwGEN9ZUG297EPwzZvPDRx0jzsa0JYN68LouHLhNh4OWRD7ya/EAYpTKad+lq
ewvwoZjVQOwp/SP2271F61y0mWRA31PD7jQntLPOsGpgx7RufbaIR7VdXxYwyBlw
YFDY/TzbnljqjqrbgCzDqyo/sJ2oNXmbi3oNeeHCATb5e3LkyX2jiqyfrqFhVUxL
2lXuXSTllRY9S+mFsakh5jKyQWzMJyRPjAn383AcIhcUiLB/M3IQJiucYpVGagk0
ZIxIhG+garqV9T0S0ARLPo/XoO0pLJ5rHX6smkJbzylWCogHk2aorzd99i1qnWZc
VJGvUiFdAJWfXwkALRgEarmUeSiDXUe9/u85hsVuDiP5GjsgbXbaefv9/0y3OZG1
45teHbTOsEUMcAsvyM7V3LFKVWqQVpYo8jdkw2qp8IBV4S+EhO4aFhqPUvwKxxzm
ib4Jgv3XxMuGIsmGKKUDCkLqbN7wN3748D4DcOBsjNP7AYL9T88FXCOrW8LcYZ5Y
S1G5LanCbxKi61X8Yu/g8MQArbSDKKKByiDWVbGPEEAejeX0dEw2vacQOCN0lYjd
Ev5L3JjDLf8HxY/E87h7FzL5/KgDxPF2A9DBsCwt9ZGefuSf69yISdvfsrdnuI4a
N0OsFVYzqBq16DOXQXbVKS1ngeOTKIhmPeCwEwdgp0KSwMTC1dexvkCKJwAvsxa3
YUY0lv6tCXXXqVqG549hvQhPS+kyV/5M9M9BQAgGC0QyttUUhcwJldxOL7uiVtkn
y8aujOqS/4cpxV+Is0OH+bSSI96jmNmKhwCp/xLunQBlLgTrVRn5pUGhSLQqK3rk
sRwf5bO0hYg0OmHN/w0vUXWCQwFEylo86McXfiKmN0OUWrAWfYXCw8e6b9660o09
ZOJbqpL4kUUiHddVjQh7Kb9aeoeG8EmoWKjeNfLHXCn6fmq+1yUg1HB7z1KUQWOG
hXp7HoeXQRKlqyGbmiSkhIOYjDOhHNc6u9FaxLZezkPiT9G1Htu5qIrn8HLqUgnY
hzaDSHwXYTOsj9eDYQGlpr8peaB/e1Xdsl4mtmU+EHzyzon1o3pQ6SL/Aqwy0V8n
005SvnwpmGQ3XdQ32r4lzgWRo9w7/00C4eDBgm2zXGAHiEgf36Fah5eoUzMYRTP7
hy3e7flfW7eEw7s40/5KxvhuXRqN5VQxDo8+o++ZE2zZfLUHpuA9xgO3P7iM2qkx
mOjnjhhJQh2CeeCIsGZXtlD6AiMW4HxuEuDC9mMssBzckUgFAYYNYdFZIKBpoROy
WcWKaZImdmPFEDAD7LFbo2JKPacS6cx7IoLeMd7f5mp3A/wCljYoGEl4IrHcDouM
crSx+43/17kHnsYIAxv0DoSqW1iqzyGuF97Auq9P/Mqn2E+9/EPkjlGD0EDKfvft
JBmbPseAT49VAuetnhlh0UDbPTzZvkVAgXRKWE1No1pld5lGNKUYs3MXs5hMaLS6
b2c8DXelQT6YsCZgxiD35M6irLQqFWeJGRBc9JPCvCPEVadc38XTsfHASCjt13Z2
tYlt4ZxvhrsOoDA1hx49bXYBzRg4QuY3zOV86GvJS+mB8I94WjCBHcnCxpN2Iskj
MEuk9Vd3Km0hWrCtv1kBxeVms/Vn66xG7myPMaihzJxw9WtsWVjQJf/V9ueJdWzS
D66KCAvBftkStKeVwcN87vLEwolUBK40FtB33aYsOS7cKQ57VTCtFFQL39myyFm2
qF/BR0dRc9H8zbH6k/uQzSF0HSgAAz4eXIC1RUZhIDOF9zLnx0D40WvfzxEKPhP8
CZsBiJrft24BkmGXacgcFVicWA8j0Hktb/XvXZZS1irHuEd8MPwqDoFV09+gGRlu
3dMKQgktyjcEwSynccWI+5waRbCg/L/OvISiQoRZXzcieJBnq7s7Bs48jY+GNkVA
FLRJzOOsvlWHuhxKRY528EqhU7TNN3Ibqaxjl0DaFpbnNbF0TQD+/XRMgB4b0H6Y
aVUN109a5WbKXdBmFV+iC+65E2BWSmdsHO2b4kOxHPI6CrcAqj8yrkLd4wQXxIIT
w3xHJRnAzta3EFLochOzj37C4lq/0oHcNNhthD/cx1mdY1Z4fr4+S6bRV393IDgH
onWyjYP+G0FZn72ZlPNV6xTyiDzjtgo6AHsJB563VeE5rpUdP2wBSSiL74YJ3rbj
wxQlofVSt8mFflAFScYA5DRDueOE8IHWJoLEmcQYh4FguDveMCtRF36Aoy7qgQHy
/VNs8/7n4ng2A8YPRcqYRCwj/qz1K0lHS8Mtm4X7OMyvSSYDuIhdenCw/IqaYWnW
b7cCLXMG2ObEtvNwG/VXWt6KjRDAQIAa2CiwXf2rEttlI/6uqBMv271iM+S9E9OG
c75wzfGFwTXmFhipgNERqUxBJoe9Dd6pB0tc0/SEWZeq4sLspbg7jy9/9cxziH5K
n75np19+7NMavw8FW6l7XblXBp6pf5UXgru6DJlp9Gnqp1BKZJP80JhIQv02s058
PBOWwmgeiT72LsPitygbnt7KZKLqynu4N0s7BTCTunORsUR+zSeb9OdcbSbkxU1O
11PcB62agBowHZitiyMYKDZRxnvao+BMVlloFgCmLk4i3IYCfScdwjUVl9FoXKFK
bofOpnh1gNWaFN0E5QddARlhHw68HrCgotJ7lORE+WQbr410BF/EUgg5o6dS073e
0t7hXatinDU+qiMeNE1mrs5gaRD6zTgHkpPuMcj+xRFFwRl8VgF27u6yIjMRtbG3
lOuLYLicQrAn0k823/Mas4kn4lhAlr5yQZ8Q8y+9mbdPYGOGAXvIoZasc6CNvd/q
RL0AAw5gWG9mPtwEyT697KTiXwlXKc+/u2/E33u57kHb9zfG2juflvjuJIWTWke2
AX+LRnYye2hKSKm8ZNmu/TosSmIeH87FjAf3w8W+AT4qJksI6FzBnDqeC2QLT9h8
ivTPGTy4jJ+wGrE9ozN5QT8E666W07SRsAS/R1dIcwrlybOvbiP687hglCvDWOzK
+8AH38Uxm4zjWpUPUeo0SZA5p/fMTwdv3vsHkN6gGLNntcqo2AetaAnEebbVzLQX
OFl3/4Zel3sTAQm5neBPNu00TrbQhp6Kidr6gVG+rdEZRoo5dJFaYPIOSRwi65J6
MWBRLxq1yj0fuKhoY3JFFfBbqMoErcVEXyqoIzkIy1cEa17Ozn72nblcL8iE5mqy
9MVyD+PJFiudwn9EgZAvLQUsRYB2V2+UsXiwlyT2xyLqi9DZvMkq1T9vCaz2+2L7
zP7VAYMXQqhJca6K6CMrtdBCJBDwlVwbKHfY9xK7L5au9JeKA5LKdTl4fxCAm1Gu
agroKBRVTLtAtVup8cMpw9aJYTuCizPVnVB7pwuyhkt9OQq9y4Pi9ldGQEjeGeM6
tOMdWOoK4vlxot89waz6pt9O0sbpdwtq2jYpmAxV6wfh97tfuLZzcZehIqPRscD+
jXSxoTIos5KJFiGrxWxfbPT4RHkAQHsypHNzqO/zMehPc0d3bltSEZ+OmymyojMZ
6MAomHgW7LDgDY02SzoxUhl5qwzNMmXnAxFaW7koi+T9sVhFzDktrMEupLZTY6YK
3Bu3djaBObbT8gT8r3PWcxV/W6+JGbrREmyV18KVJsqB7fhBzRgMO14huOOdxzqq
/kXrt5Q1cmZOqqKJKtIfaVvUmgYCh61vwfHQMi0NpH925RATtixIghh9+Vk4ghpY
JKWaXft1SZHl0NZPCP4zbuDmYmYWE9b1/28vblCgd0dCDO2XBWo7FPr5XGHjpvVr
gjtW0lKDD9ek2ZNql2rNOuv+FWpfTlRu9XHafKCzqLWlxAg4B93fyciinmfYq7Hu
709amaOQB4pRW8NyWJJQkYr3WFAGAGkzEAsC3mFlsOl7ntMAr75tc22tBPPdwDax
eF5SBPQGf+FdkGqX7JYB3ow1d/OXX9/+H1woCbJP1e9Q6tQeeQ6squh8u6JLdM6e
ODQOMfl4Sa3ubFnTejilIiU28aGMyYbuHV4ulxg0c6NXbQBl8KuX5Sv9wqY4hJwa
51ztBK6oNhsmQZBGLMySUEABOzN/0Iz7jHfYjtjNzBlEtFevKX2jmU0iMzx2zUcy
ANVenPGclF+2bLkI/XfjRa+bSqa3qPIxeyrPRMwnPG0q+Gryn6O3GibbYMZUKph3
CAL9xFqByZiRcVWqVzTtAFUzpKMVbqgsHt3ZIYMju0FQhq+0UyX05sOgKd2LFe81
2WTH9ENa2ezbp2+ERhm5qhuPbU5/rSx0ZeQEk8AVGc9JSjY1alGqB/jzDhYKLeLk
NFUGjCmP6LXq6evM7vCtZC9gAzx0/5cnC2c7kFzrdxdKSipG8BObJIOCEDx8AIxr
t8heghpbQZ/1hXWNQPSu0+jq5se2FVodi8wBnEnjX8Kr3hnbH+trzZOAu5uYAfG9
eREaEPAh9BJI0neQDpO3Mntz/7fnCSUt9sdR0u8XMKN2PVYcAQsLzXwheMbo7o0K
OJcHMEgnJlM/uZ6WcUBP66q2uNX+qNWWOnt+mJYOqLAR9MGSY2tQyE7hE0pChUnd
ykroaFCeh0adyslM2Yxrz2IZoMBYrhGjXuF6XLnaHok1+ezdaTn3CNUIG37GFmr6
R/1olZPXB03yZGeZnVT/2WhqCZNw4OuCmw2GQocW2JGwMzBZa/KOHWvmFyTl53HI
eM4D/NOJPOhORQDHGk45iq34IjDuPtHKdeLVKjVZQW0IWn1dYwLx7cfKuBZPHkT5
eztz65+bXSFRJvuEuYHQxZjEo6ahQ9jgUKq3VC5brzUPUN+ZlmiqdikZW0EXmP93
Qe6zO+5k+EM+WoxvagifvNnYGEjUCr3S9fVFDRrEj0Dxj2Dfs8EFbF6+CwATE1JX
80BbCkVYfXS1+xjrNj234RuhnFmd8NxyS/1SrRphO/xK9cNc0poNWPihRCl0YFsD
AZow88HN7XLddVyEsvTDn9W0khekNDrCMoB8ll2ssJHK1bkl0+zz9ebKwarHeBUN
+YAR0VOafz8QXGBKjEPADPPGBVxHJXD1ovf0LDh96C/nAUD4Ub9sJN3cxUTpUiij
hxoLJasP01FC+FsKh6BieirediQ9M+OIABhCRT8rRuKVfF2pSg3zaTFRA2LciOG2
WAzSq/VRjY9fGJkKjTAKvRWVc+IqV/cHqloHmfk9CvrMFadLB6jliMQTL3g9VWuv
2IC5unc/TRlFlYw/wUmFIYP+i8jb8Cv1PcVb8IoTzgEEKFRGepkH9nDz9AmpXGh4
ySI0KK/95iMR9a+9K5fW32UTA36ZckPq/FLRZrxjEjQ5LdOK2k2Hp4g+zM1yy2J5
jwRZbODP9/HrF4LBgSN3NYzKNHji2zMS1tN6IhwtHTDTdISXRdds3csztPcpp7tD
Kwdqqd3bKxlLyIlNcjJKf03ABY40REje/M8cKZjOCrOhqwVgSFdI+P7uXYeVdmDE
T+KWsSqI3gttFvhAiJvChVhOH9NnEuyFkA+WZrOWYwQM+0XzIZXRpckXQcWvHa2I
rQonsOwjX3ZGQ/3MCVPlb7OB8o3ALWU+hZFXoBV8dQLFwoCSRLFPgEev9NsL2OeR
b2Z53HB090EntnpOZApJvoRtoE4brgrVAFoBjJADKNdWZWDpJ1Zugl0VAE0WVFFX
1xeH+tD7yELXDzUWaxZhezLIsZbO0t2S7A+Rc8oqV5k4AvMLmkNReyiTWGK4abIh
e1Pm41YQAoW1I9Gp5Bd0IULzNptJtNeeAjvTePqPJeNAhbhQqv/lTegFsr3ROl+/
mCQjUqlcy4lnqjNIyEdGLoARXzutuixw96Qyrcdy43YevrJrvWJpaTXcVMODlyyT
V7SKBM70salm1NCUgqTg9uJTOqmGIiMxBAe0/975aWPfXlaQWWIh+7Xvo4EIBtcX
1kNaR1zfrn+NhC3iUJwwRUaGCKVjZro160chB9raja6nb2j2LfLD0g8a30mQHotu
9DS2gxVwUt6V0YMwZ9W9vYnNWgVEFIIRnxYV72HroTQWeblwcBmPNCXa6PVQpc+p
Qxy0bUiGWDBcXQzQWi3WMQTWNH+CN+2JEYSNa5trBFTJD5BwGlTyLrRAFmL2wdOf
hl6/cgRTPR4UIlLnqgq0oFTFilcYV7QPnezTeAPPTnwFgVBamH8D8cErxpXCCVxx
10exgKrptJoDt+RmI7LU6qTWVLjTVBzv+E3eZE/75ZoZJn83OGeEzURFHKDWp47O
tIgdK+PuoEfcIieKkrvPxm+aCcp8ZvcWHNwtWg+2pBTs00WZ/Ycmj2X1r7Pc91Gs
fWu2LNrOA2Nkzow0UpIcCuRvfr7oVykxur4uTqecxTzi7m9G9mre/Wgw0u2fpbcu
NXBMPqu459jFg/AQ9Ki9IiWQ/iTHuMx75YUXFQdkFRNfua4ofRtYYQpXz20/4IG6
vvWDqoPXFXzrim1OqZRm0I5xE+xLmLe6fSb72YD2FJ1Cn815mPqzb8YTHmAA6reV
Al4IeHXrkX9yjwjyZcX5Y1ebDhqqbhVVFK5UOB5w6tFDFw0G/kbOKFRO/jkt4kwK
VwVQ3VNTdQRLL99p64zM4DEd0CPVx+z/ohTY7IPdwSvLeAaxXya8xDH4tIWFDWEU
x6FPTYhO9eCeSy6lObzAnxpYyufczCKqLykXl6e0wHpKGFYhvtATpmSKZpldl6xC
yo9kclyfJ2F9ek7z3JP0v0Ry2sBWdc5zhRHzzsFySEndABmXrH2y+CZf86gYB7Jy
7KkgHj4lCQQweeMbHGUrFskDrkA3jcfGBLMZFmoF2Npm+Lt9WM8QD9IBa0OmXvjD
/EnQP4wKe42kuPIQFpWElZYzLUTT0zTA8xTGLgfTMADTxGyFx+qXfEQsH8aJDl8m
H8pGORjrpb2b4QzlPadMmP75DfIUEbb6WtWrfr1oJ9gVTCWhBLNsqewSn+JTayfg
No8aBoJBDA1pWV8OwS5ia8ULc/Px/yAmFeuySgVkTRpUAqp78axwC7epz/31FRs8
laKqUbHrsV7iB02F4insbK4IK5ZQ6lxCOCN1lTq4c81sH68lAjZJbNNvX4Ayy6Wr
EqNXnNNAcojp0Ri74F6iX7TZNFIvfgfhOJa15BaUVDUymBPvt7GI21N0zTW0dpMX
+KWZ51T2r4ZZv/5sDOLgKH3gLMbn0zdLI1oL1/O/Aw7RFSzvN1cgJx++gpjH+LWC
8f6EZXtzRRZ45EtCGBfLyl2CbNdVwWuRR+Z+5ryDAz8jsnegqsppoIGlZRHEMwHD
arcfxBDuKixTtxBqpVH+QXJqPUnh7DTjpQp84r8tuU4mAuddChZVV9Z6RrRF3S7q
H6twmMMJgzQGkjuAGK5AoEkcydOqqDD6M6t27Si7ozuC6BAPRMnZLXTepy0GFRDU
UhY8+swixqfB654ZExDgvGO/IXkCO+dvKVKBHz8jSPIG9ky1CdzRYsLXQ4MbqBQQ
JgdJazzCVD/WjoUjQ8tJRPpjg/ZESbEe2myJIg4nknGGBKsPlNse4fAelDAKwO21
vqu/DfloHt70PiemnnDLsNlZw/yfd1kce1vhco/psFtgL/ikWjeAeCIt3YRkMuJT
lPsAKMz+7yKjTcVXst83fBHxP+lhD5CgVM3DSof3hJDkHkoI3YrdsSHiu8iB414l
GCbh7mKBknXx5EJdGC6o4XrZVSYB7gEo18St9Hhmk9K7xcoLjTE4AW01bZyBgfEV
CZ6NeiuAi91zTJWw+8iuEb+BsLkP7PSVZLb6TUwn8jNpLdXjpDVd9tL+qxbOB86Q
+gMvY1UbB8wdVpxq/J/sTc6g3+FXYuEi4KACfI7MlS0aR6jUgzHmcvVoZlY2J0Jt
AioMbxpwhR8EdLOu+18YhIvC1ED7Dd+6hrjgfMIEOQl/ChVnoSoQ9sRbFpo56XsC
sx5AdA/EvzENL6cSKbSCbgNgOH6rrltfoD4mVnKyn8ly65MspmHpLhhCJvPg3MF4
SQVuDZwknZWA2MmS4MsQRrTZEb1sfDd/27VSC+ndm5g4escoxo3QjrngMBBJH7bx
jhw6ur+3GtUGEm0w+SKf5rIs7RNgyKuCPa6s0bzIpCoaAfIT+bSVF1QbAL0oWycL
gIoAPSvEtLl/MWaw8vDciVRo2zPjOWD8AoZRYCL4aGBBJfrmRxV8mNEqz372oXUY
cbxzd53xDt89c5N5D51gPLFpJXHZvn0bCWK+6m+1bnGUSMjZL4SXEFRhLdTb7tOi
HheMET4uAqgUqHV6xDEeH8MaK8yNRTqnaynEOzhfZOGr9R3UwgtFB43AZo5vNTtY
r9LBEoUrP6R+gJBSDMWkwxxD9gmyt3bqN7f8XgkaxCgP9IsnxkY7ipyMIn74AK3t
Yv3g2eBHjBRXqIDkdrJN9j1yq8VSkRYpi1NuM9CqRuTIProDyYCMpS/7qjf9jvTb
Q3lvWszf6SuEiETf/6ikoefZSLMVhJMtqH8InUf7UOoBWQZFusdzitC3m5QtRVm5
ULJcGuVjBpsAnt/k/Q7x6pafB2ja46towEHnrzvhdDwdEwkfdHhHRooakru0Imvl
XcaH0O+Eaw01YQiLuVcFh4bSDAvHpPxg76d7LD+IurcJcjU5X00Z8BfQwNF7EoZF
SicSwq5cgIQtKkKnpb2j0w0SFnDGK2xqL4zE0L9NDvP3gBIW9a7dk8LgOeu8dSui
v8tioqo2ONsgVV0CPawO3t+5ohieAzH19dAPGbLzJi2+OXlXvn2zC0lQsRzWxbCA
XLEwqaiFHo/KLs0N7LLzLvVeOThsltCfD7EIJhYRmOuTv6/tEgAjb0YLMVplxrZa
uyeL2f+SmpCngocSl+GSHKCiyjEeKXVSGzN+Ux8fK6t3+A9TommpX4fF1urgw7VJ
uB12MSPeoSRuU/v9j2YMTiyg9ZS48NQoIs/aWuUR5RvT0/8a0ZDMyWm2LOre73SZ
l3EzQ3+NeJUBfF6EVdRz7DSzYNgJJZ1eMg7M570Q5t+VYsS4ARsczi6f16d9XB+Q
ZDnknR0SPjluCfXVw87p3xkwxJVMfHQrID28AusvQxJVud+1Qk5RhyC4Jf3OvUrK
+lCpPfeezC9Mz01VTUK4u7dRCOa1lE+fO8rQ60dMVYYjhP5KVbu7ZwfqGZTlQenY
kJG+ZrzBh/q6IxHdnXQ86BXB3dtR8Sqk7iYZCiErYiMXMhfEzopteRuLEB2AS4OQ
xQKfI/+2kpt1sjOOI0yavwpq5gkO+r/p+mRonYhZXIvKl+/a/+bB4ZRYkePRcawA
nCStEj5dzQJ0kmqSK8YTyacr/VF+yPGJiv5pKDSyBXvo0lLrT9ayc09rHulELDVk
fQPvP2EMkOvhnaAkV04ShFetHsAJ13Jo6vBB4jw8Kgg5812dc4xdnYctW5ZOlzc+
UZSLusDN4LBGedlLDZQYjd6xTIDHVY6vEjDNjAOd2NsJUtsjyVDYG6PjTK1NOM+G
wH/8psWV7rj+hDalagNXhmOGS++C25P3GDXkVatBfyBsTbENxR100k/toQ3076d8
5Uk1IJJ5HTVjKfWPuaFqg8zWS5/7NVpos1tncNgm8HT2a5h31nDP9/IsVoyAUBv0
ZlesXo+aMbJjiW/YffNPE6DECKW/TyBlwTGIZSlgOR8pCvBzLUKmdISfzJMG8P7s
RngkjyY9ofntwlF6JazS3rBSo2Sah6jsNWfTxjReav7SApQY0NkgA4eqLyBzQFfM
LZShfEqPKuTupt/Tj7OLLHrndz3wz6PSNzGheJFD74SqPoi5+DGl0Ty9WpvguWEw
j5l0Vfyl4wO3D+xnda2vp+DNRNTHfDc3b2sNGtgLErod5I8i9RPQJjp459/wXHrn
kh3DxFQnHORKE9sSWu7U0PHJNotrBeB1MOUwR0z65KqMm2yV20PByCtlv9RpELoh
DZ3GM89stbS34AA8RbR4MQFVU3UwFO4A/TIVcOe1oIpaBqe5AK5ZQTFH9f40mNTW
JjbnSmp2nVxVmLaSLI8Y5K8rV8s23DK9a3EAOJDxfXStTZpz2dP2PX+EOsYKKM1e
y9N/WYXIrv7F0UAweHOQ1+1P2fEaObv5hFejgAljd3cp3DPE1ysr1fwjtlD7xoQa
68EszGPHgBi/m6p4KX47ZjdnuAP1iNZgiXqvdKviiOZGD3/7PrbNKRPLAB3Cj7C+
RPdM5wcaKY9I1JqVUmOhw8f+Vsx9NWJWuKy/QCWBuwbQ05pgfN/WgltuZ64TIovC
8tWpj1dT0d6XnTYqLaBhGQcVZO+EIxjzTKQTO4ZTqxhWVAU/dnrNcH+kRvfRrIs8
hGroMc8jEY/YbUsS7jaINWZuOtTrQD61pxhIW5OAdBm7XVmIYQqpOs7JtSahJq9z
d4QYi8XN37+mIkOy5lWR/zhk77CMZW7KOd54rhtx/CKaOoe6C/2DVsljTHzk6Ufa
KT8w0RnbX7Yywb7J9H1bWcQSumcj5PhhnrPFjplRCtyfYlQ9vWDd2eEdzVd97CCS
MMQj9pcpjOUlU2Hcr3VYvcsA6XkCppbSuhY4SfTwSP5HI+6SBAwHkn3C3o+JzJ2D
M0lKDMtcRmkwQDYbwhAkIFJj6n7Aya4RmAr+f4+Rgot7PCFnbxLRmmsnXJPBbz5K
7fBlLNP7mQD4M7r5XmWgxn/+I5VolRUfeaISh+bYAYnWFlYyNaBPv1mfVOEGd1/j
Mlp9CaM/GdOT75yLrpS1NcpeLbXRUiJWoAGXnCdYYeGZnMjzh7EF5baDPpWn2iIh
+WjNRbxVXgRqd5wuKXDy8vuYTKVL+x4asOItzkpWkI8KFtrhpIoo9UqZ1aelleo3
75YWQaIHnt9654JWkC91aiIfu69bzDh3ze1Wu0IqC/k3jUZymVAMHj1r7iiXv+fo
GVI88UwQ3IO4jKvhnXbQfpA1FMOsIiD+ec7i7sTcJSDUDkU6H/mQJAFCrbAjblds
VeJqrgv3xRJQtdLfgjj6XGWlgengEwYWxurTDJF7moZYSYVOhNkPPiYiAm2FWD6T
2xQl4FARpTiCm66Qr7BGMFpWmgJp453jBaRNz4CGf4FzIFUH/AgjOtONwu4B44vg
PzF82spiTsgFiAGc8EoJuUn76F6E759aGJOHndVFB3OUyd/xXgKxuS4aFBCTCyK+
GqW3j4fAQVrow3hdie2lf7OzQh0D3RswRaAYw3BJG10/V1es5y8zok0sKQ0gJ6JW
fr2UJ8I24M8/sT1Kb0ac0cPEpCN+MAEZLtCANkRUWikY0CafIR3e7oNEOifIgk5s
xnUx3Cz3zGg51bL9FJFYBQi/0U7xxMu7vVGK9z3IN46GAQtR0BRVCSmpOSIRyGSm
H5xYWl2x8kgY7yiR3hGhFJEEEZeEPnCSJ3/E6NXMSqHSewmCQeNByKe8LgAOhEMA
9JYekRmmXyL3MrfK/pU9HSIKFL7dQYLkosjqtTQOOiKTdU/jQCHg6MIY990TRCVQ
ezMbMY6QpeVXAWjYKUAm9JtHrnTJYo93pLq93BEaEQz6DC6af3tw8Cl+YIhnkEZI
2fCUVjSGd83eSbKE3w4UMUBxx5JfX2fwdwCEaRsRr20JCYJtdpxxNMp2jGaffwns
3I93tjK31b4yi58AUZkmKtKyXbWDCoWCu3Rl4WsAFhNrVH79txYvEc9Nyb8WHKmd
pbYCXEQLi7I7L6RVhqbwQk6gtkTVp90/9BT8ewYskX1mxbI1IT2v4puUsDYz8gSN
itqyhf1j3oGsuHR5qwkXdgTTiFuhexxc9RzaqdoCEvg1K9QDf7mBILT1JuLqhixv
4gylhf1Kk53+HNsIuPLXysGgw+lu2kkE7C0hQ89f013F5lkQNa5EwVXH9LXh8n0w
2ECyIiRUCqwaT78Lqf8XYVSR+zTGrsIRqw/IbkUEfdyJApY6ha71iJfHxkPXZ/8z
R+EQyDeGjtyKVUylC1yx8APoLZjiPusXrfXbA8jHhdZLXBdtoARYkknjZGyV+NlH
NssCZbs7p0ElZ4gVQXdEsl9EuhqT0VOT/z3nfa4NJst5lK1jRWiKCg7Ewvhjoz1b
UZw5hR4IFomcitsu0de6FESCihUszEmO01wYFWk1d3kEUtiESCW86jHdFvrUMc0e
wNGWIhcGR9/moiTvchoyfYeSRzOfI0i6gj3rfDsiz+yx6SxakaibiR9yXRcIqljN
KRhvgyJUGVnNi9RzUA8n7gWNs+xRaRF7XOnS3IEEvORR9gABellmH02xgUPerrEN
btPnuwMCGeMmQdZqQB4rt7DIT3qW67y/2c5ZLVLSi4uygk42oaX5j4f4v4Ho1GHG
fhPrPmhBP/hY7qMuH8iICc28Sn4dDLHkEBRAlpccS7dMAbI5qBmXVf2CroRnKr+0
i8kHU0zVzbu1CSmhof9TKykdZ6Gaski32MMR/jw708TRRevfSG640XqS2bUgpkKQ
U5ASe+vZGnnCev0ySdsBeGFPiM8QValIhKtXJpAJx31gbtU46demvYzsD0LUmX03
SJMMWUP/P5sQVK9OAJSyJo9969/6rTxAiT7O+KtMDmXA5xiz1m6odd3OASBQrBDo
tydZnhiRSw7hyumvQc/MRjT9Gg4NWe/AZpqEbBvm92/SAt2YLshT8UzcsSHNAuwp
XORC55oo3D3mufemqg6uaoGy8T5sUHshzRcImTtzuu2+MDYvLXnrghEKxgQyF428
ZcehMtQQzCiPIEJOcGEoCaSCa/QVO4BnVDj/cKfKSkpRRo0b4Me5qfSRkxPKxU11
CMV3LnCmdJTwKHYKSvzxB3akClKWsEHfh2Yl2diImJ3XVdH3POsoC0GSvT1fi18m
F+xOZHVzRWsUdsFyIkdi7Hk6/pG3tICEzX6OrhICPXEwhnkrWpTR/qw7P7og3/mg
o1wuy9yBHmCqamInX6br42eQPUUYm6DNMQJC5BvXj4t6m1BlqOSpl+n7cIth8Qj0
ieCFqBtX1/DvsANb5cxWZ50w+D5zEUa3QI0moEha8gWuFJ4V7s+gfZqRiJwa7Dg/
BzIhQZVB9Q7x9Xk4Sson4d6eyvCb2G/ouK9ikIIa6eqaVwJigQpfnmtD6lPGq+eU
7CnMECcpDjbUO6hn5seiEWC4axpVBUmZF66iEt8OUONH2uBPRdIVZBg+XMOLjqpv
1goKuG9clQyEVfC2xcOs/sYIFLuXUPEZZY3XQgn/d5KXacbwUAi/TFMZiqO/b6P2
BT2wfI1b7kgyynxFHn8Zn96z+PzNBAjcY3QQW7vTaabP0ghaQLMUTLHodNHbEO1l
qzRAeuQJ/cwOlb//Waq0mOVtuc0ZX8uSLDpzBVDRqQkwLFBdnkghlo2QEjKWaB5A
jMqiq3xdrI+hHF5UB/iGWnpU1IxOkqdvpaFpAtXry7jI0m0fNGru9Y+FTnnOib7p
5uXxTzatIauQhbNPy+VfWmexIAI0j0reVRs4Fg4Z/lQ4FUbQdUpTLRlVhc2pVDyR
PYsfSbB1eAjFP/cLcLdHKzuOpNkMddW64+lM+gShT/ryV9rKI7GacU3wySL2LU0w
foYi7HKLGXoBV4lCek0zKozUuHBu40ChTIjPBAvC3xonBS2nn16ZrybKGZ/KXxXF
Hn1cgNySKkZBOMUtG1BrWeW8Qe8ZuUF3r37P2CmX/GxFPJAyDyagyHgDm7L2LFfC
bkTc2b35HwslRmUSwZPxU0D+vtE11KubJXBoXQuuiMq6dkq0NEiarEfDo+lWS1LE
+zAmaTMAenXojv1AJC0c/PWviOzGs2BIXIRG6c+TsRjuDQpqQWX5rq6S05kBmsJR
Hmbon8eS5WzFRppGFOdcg3AOzCXX7XkTxTyMUgq4KldBnWdFGdDz6ndWPGm4L8j5
kulItaJ3vdD3dxewN985KIYfqFoFNEe4TdWVY5PvUQGyaweJ2WfOkSGiZJumqU6r
EBksZq0B930aqo7J736lM2jfmuQd8bPmTYqMP03ppw8AODgulHuI+h9L1FTjAVLX
NyKf0zoPA7WrrWM8uRXaT2JOVT7Y/86w7ZA3Nk6xEmLCznu5cFNlZECjjDqsjZZP
8jEm7yLi/U4KDx0jmFECu3Up2G3Mn71vIOF51ZgyaC0d9NLGS7lUX3kMYp/o7Phf
EeA13eaExeldHuEMEhx3tz8CcN6Y9nNcgq+a6PSwMwd91rCJe3BsvA4F9J1a3TYf
ol4v7G62qbJY2rG4/1JWq2cmMjqQ9driBnMU4LkL3VypfpT66Eh3z/pThqVtNU/n
PyxevOgy12h4bv94T7rnrWrLIgbL/KtBFWatQ7qsiaR7h0eDWS7qr9hhnp1hZyX+
8R04b/Ps0JbmuujdVJaB/XEfXp+awh+wvyl7GrqGHlvd6jEajx363F91wnT29xs8
cD/5E3kK8PqQAPTdhiwtew451aJYZQWpHwyjsevDM4KL288hQnVDmr7WdbFOKDPY
KRhG24d++X0+gBJqftiSWgBmO7Y1cUgrXgb4Gk2v+XtoqBZJXkrLRMW9s4DxoAh8
noxOcNOB1GvVsU2lBXgdlvFPncNwkhaNxfToiHrqvVcHwbh8jRe5PIezW5955i2i
/sUrcxxypug0OT/mjnB6rRM89njFTcg2IHBMUuiLNuVti7mcvpgVqErQGh79SCSp
022eM03nrm1TBcnycfUSe/n26AllOe1+fG89guuB1zqAfqx7+S8xI7UY6RGvVr5d
+pe4bLPQUTvAJaT7STzSU/p94Z6p5upg/c22UzTWm7QF4+KgSChwGGnjKns8JvUB
1MXY+FjbUwz+34kOROvHNDsr3I3cEtXkvzpbFJdFDU5giq4ZwjRXgEzGoaAaah72
oVG+aku8nw7d4ENNxYPGqdw3QqyTxDBVsl1hfGmwrzD95H37c1yAOij8Nx+63sfG
hWnxnS3He+GJ5EMuX1f9WvD5jZhrYO4LgtVCw3TUufW/e6GU6AZfnb6C6arKy8GY
t/j5/9zKdhWwQ8zbZ4TTwyuBDHFExVoiJZKrLifVnmFIk7TPuWnO4eI3L4aSQ2Lo
x/GXD2q+RCJ04B2AvOpuFGqqYimAqExlFXrFl6GhyHZXluMCpKPJ4wBvlOaH/P2B
jf2i6yUPYZDGvLmbF/ecjxxyAFvuDDzujMu3OhR6MQ4cJKTuKTRDuVljoyk6ss6y
QIDrn9PvJD2+WRuvJ7r+tPyFR66ssLokWsZVMYZ1sSG/GK+8ns22/ducwceGtGJI
B+3zsjh3W9Vc8ZYE7huEWJwtG+LToZThKubmNIg4wdeNsLZCTQEpyEOSJg4jnsyS
rad8fNAlh56gDnzbDV8c28cZIKFZQrd1pYNJDsWEITVPw1z9ZbVXsdRK9/E89AaX
DaOGvtCQWAxR0Fj9NgLZ3U3oUEnVdG+ayR9P4+mNhGfbF0JJ+wA+ehzXqD4xwIEZ
N4dvMqGoE/WYOfjAP/56/YG7FYv2Mz4B9rvr+chSpKqy5uNp6y60MyArKtaKIQfy
i5yGfcBkctjcYc9Sno0E1G8Cw+J5Fja1iuprOKYs47mOrq528jVoA1Q0wpz4P/RP
7nPBMQk/moJzQ28VfmlysP12g3XyHmtZ6dNVjvJXLLoT/J97r1K7n1Ae5QYivz+A
iU8QAVZZpX2tSVLjidgGKMocXQUbQ39m96mu+ENwdann9l67MQpZJqT/Uptg8NoH
/8yMOvAWckr2zbK6A+CrPN1ykzJiOsUK+sg+UhdmgXYi2+hLBUi8Vfrqa/TSVT8t
oX3KuNcSperEXlmE40BDlIaUDzMHR0YEh8tijagleqC4oSO5Evzk1qEBMRMsi6j8
wSs9V3cBvu9emrWrySqtFfeEQg2ogIhvRdbulDdNv1zPJLn2XVe5Ypbhk5tXpatN
mkaNlGJAZJDXD6/miaOgrI1vEJebvfgK3aNC3nTlkRKwiaeQOTr4xObFdjvdQ9rR
68x+e/8XQ98ckJ9zyixdqQVNVJQwvHh+TFa8u04F+/dOCyHl6KvTXjrguxSetPmx
QXQuFggkCCWcgW4GdeBCdUeKFO589jqpTenIreD0BtSF673ZIRBDxdyVdWoPneKh
gtuxkkusQnz6bdXs9jiG5ijtWYex+C4Ivr67MNL7ZuNKh+qY6LaJ4FHeEcE7gOLh
Oyi8f9r0ei3r0TfHF6pRDPjMFG3cGO9Vk5atDju6UXcqvzSCkLKmrA6FizgBKo7k
BbVM/nWHEOUBxm0FHExWJsgEwtv1DMkljrYk5IAyW+zHeUXY3pJJPKtt0Txp+yVa
LHL4+ZjYMo3wM0O+kRY5vE8CMyp6tD47KZTxCynPRZXsHoG+2FZX60h9uJ/oU4qK
fBbdLK9MDPGQh8j+d39DgPlRScMXGI5qGvdrp0nkC9oHCT+Nraa8Z2APS/wDBpmP
LSzJX6OAb2WxrrW5PxqSdPjcQltrKC5dk3NBZcFRtsw8VXjQFR/1HPMa2DxKubAt
JAGe5RMfJXSodX75lHSBkoZjALdtdeUkjtzfDcuBlRHPPt8NM3kvo5uXnGhzM+s4
QCR5NUQUvAgsgOpW8xD0X8vna4RmyHfcl7u/8PwPUpMXTCj87YJey5WDhYzldVm2
LlEd8TsvNED4t3nO+pA9SEtPyKzJMhcvLmh7Ug0O8GutHP0z1a45cyza3ueVJxgY
m7XLwVtixtW8sayOnx6YRb6sCTmI/LTvPSGcN/tn3HYhCpfMae1RfvgkhYQ52UO4
VpJrU095tsTFxagLNKTmqu+d5U9IIZo9pNHvGpt7KCdL0d0zC+/Txt8fZAv55Xov
mBBTbHTOYStO2kRgnOqRjYN0HrckckaRJpf6FQzbQAs+vKPmV+s1iGr0GrzL9n/4
ajrSPLebFCNPcktpqxxihJEW4wvkPXuBK9OlsUKhT2LW5GpTEBPDLO8x/Z4kZL/l
wlmvmxqNb8tAcialE8YY62EIqbrgD+jIY9MwNeDMquNGoekjEpOpcJ1a3dgJbVPt
ho4sD6O8Pm7syqrFVLyGO0YUZ1mTFQFTMQLTKvZfwJm0yRt7OXG4UgphxlDbtxGR
`pragma protect end_protected
