// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gLOP72amY6hwNh3sNc/MvE/osRJkDybsNpRBLIpP1/eZDZRg1NJLxTG+zGS4yram
vhH9ZNfAndUL8lx0dGsRHp/KJP3NXqiFnNY1MkYOEKsWNjUaj6AmwuvLZGpEXwOr
EMHxIkLAcLGzAi/afBfsu6S0Qgqchh/DsrwuttbEyaw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14544)
Bhq4IrDXWj00XBv/EmaCYm0SImYxQ3Sf+Uy0hWfxVOx40pOHmcUaHSaCSZ+Bl+gg
PmWpv0yFOnqa6wPGZRSQpMYMG85Uw95SvwAVNL3q9q8MJmjkIIB2yCAQDrxvl85a
h31c7eghkxO8c0eXkw3yb95QQAw+lz33thdf7oKGK84u+j/KkQIyH+59lZTUvqAP
YWuGR8+OU/Ymy27J4+yMrk+JC2VN6r7qUhimWuvB0dNAMj7g4lEPgyqbYgzqVk35
BNDco/9jwAhNzjFL8wAnwr9q+0lum+KT55enc9y+xIB1g3gYata97RJYFV3XVpbB
IuwAS9qbRt6ppPPFlLWfRVhxBH2Kjqj7Gl8x9TvaXwAZgae1MMWj4CLzHj1RELbA
OJVL/HulLy2L4BYU/bEdW4V/0fbVG3sOGg4lLjhXW2saz5R3ZO3UHQ6ognEX+YIr
yGVkb7nlMUcPRVyKqG9C4WqwZRmDadzT+1PW1M1aWndcmY/P2DvNMDgJE6NO331P
2M/TiG6HG/+oompoB6BGUeQXnFnO2shZIjTiIR0YVyepRVH1g/ahWQ2crunn2Pfs
y9Wy4i0FgY7h9ZIsBCcSQro724t5wF06sAJlejMiwsKuvknO5vQLqUeaAjTc7FQm
XixXcKcD5P+RpEDX5aT9vF5J8N1+zFxNthOHo6H5y9liixgKHdeiZJg/TYIz6Mqn
VsjQKHUSXz87xaOJQqAeGJmjyUvCnh9LAaYT87qT0Ee0VCumXymf0YAxPhvbEYG9
oxq+r51SVcaK/3cQf43BVCLmt+9fo0Sx7+ml2fWbQDW+yqe9HaJa4VbfFVZuWuoS
sDzYkVpN4da94SAWraXtQe9dsHu3rV7/D7Hm25dQQSEzFIB/C/CrTwm33M1JzJXT
ykSQMaqG6LSu45zWW8+2jgvQkwvSn5OxnW5pfjgzcGqrsdHKaMqV58bgWWF2oQ2Q
MEaMi5VURgc/jys8zDkznWzfR7rAmoJtZ2WztN8fndXicT841m5n7c28/aNIdwzC
W1EMoPVJt0i1iu5ITNdT0D0XzZ2hOI1UEvbFNnigl4R8bNUFxBgCAwQtX1HwL1WN
VrBtzuJM4FM2gxD4BQx/9/5uj1xtoLZIf9LUyM66JoyECbektmEmLOIU8CopRHZk
XknRutL2Ai+v37Nx97cn8P8Lhn0of/kfMObX2KzVTHKYADQDetXcWjFIGsjTyGdN
cjbhHfLlrBRxkxeMoS0KdMtxto8HVYEh6hJ+Gk5QG3TnbeeK9H6N+O6uaQvZP6il
k3q0vaijpkjqrY6eSeDaimdjlEnp9RLWc4saTITKBe0RRrdXlYYI1gCKSXF50Aey
nDo+c/BcQ/Y43qjJrVJMET+aC2JDuMqnzm3E5/raNlZglgmGIY0dARr7smcb0XQF
SkAD1aPrSwWVJkB3gphNKnnA+ERC1Run5dtjrifOXVYcf7wNL12gccfsZiXHlNR1
tbDjqfUNrtswbWjlW54bfS0JFwzYL6V+czrRrAznaPqzwGDFFAhK7HUTc4YvYXMY
b4Q2wDiHCcrpFgeEdKhounXLqdbSNzZzey0peprFix9SvvLE/HLb3lBBvtEPuE3C
EAT5G5B25IOtemBHbtvjSY6W+D++h2CP56x1+8+lvuUJitunVQBI0hrDTkJzYgvy
VVbnl5HZOluiCiz+1cRSmC0/exxnODkqb5ekBkDDM44TJofVUMRjjcb0gk+iQ1iI
XiEXX9UIUnphXd5rhu20nobugu2Hsh1cjkTGOuZeXeuw8qoZwXcOBuxTGxrp62cr
UX5fYsYwrmKh2JRuwYc6W4hYYQsoIsD6ilQwjD3T4/h3cQynAjKjBY+IubmQ58gA
yaZhTaXOi7ZEHB9n6ZbSHB5OVpnqXZ4KnQggPBEkGCH1EczW4SMifeLohnI7SGJ5
Mc+fMtqA9ypSdAkDRA880h2pNR7VU0uAS7+NJqSrHRg3OnXavgvzkI/4oZzUceFC
B7DkNEc1rRNAEfeLDcX2Xry5NAS1Djsq32dsc+ie5r7dqMIy8TJWA3P9UeK+Mfg0
AuMtHbJUDNwFRJcppvyh3xeEp+iBbGOzifR7/dPEKd1c9SZDB0l2CsfXLUIvcSu0
rauzdd9eDW806Ufu7s2gsywv4H8NGI9eMGx3vCuOSTV3WinZD6rqkswenT12OgCY
bSahQ7fZi+Eh4Y02nsthMSiQiQGtIo0baXxo9PlADseAVNTmVsgqlverkHLDDKlm
XTBuNWqwSlDnCr/2/dHzh3cPsJj9CZWdfLnfHafgdlPG+VASJ+7rHWi8GT6EGM5F
dr3nrpEykCWabKPgbiRQU/ywDC29Y+DVHgzyNZCxiX/FzVI1GblaZf1+PT+Dw7s9
+s0J71Gugw4N8pe/pUF3q6ka6VcmROsiyX0PcG7ODagUUC9WkP7Nx6pR47nO6gB2
2a4NtMMPcgcZSW5zh26RUbw69H/gsvZ6P76IlTXnzHl/WBihWPY4+TtkawI7fPXt
Z7s+9QvZKuw0Gr8Jc7KIEgPbZ7xj5cfwYguNhowLutdNi6xkMbDtheMSy0pRdjyq
vq83Q7A5dldHHUvOfiA69/+fGE+3yElN2+XuNyGO9ua9KfWCuhE8R9n5B3HnK3A3
uRNzRdn4r8h//Kt5uNxie5kL3kKFBmWNnSsSwZ1GNW7w9UrSliVNQTV3Vzprw1dO
TbVKFxIKC/g5f/hOnYhE0A2lu5t56iVAShY1+DD+d12K6Aqp2e1e4x77RtvwP15w
uQpbM8CZxSY0MJgkYlHbUcAZioa7MpVA1LN9TDg6ODEn1fb8yO4/tewLKk+Vg3Ke
n8uj7KLfdR1MIOnOl0CbQLBp8tl3YyUWtWv/VsxwvPsj51gCTK7HZG9xjUA6YuNl
8UDFgRF9mctLIOELfiZd1tj5+S1j+vLndAV4s/u/nnLuNb5FmN9EgrJCXGTirtkM
I94AJKPyvbwFWbSleIlIC04pnt0FzVyhJ4voTE78efDk+EpeG8t6PeNUcbVtobF2
N3ANeV5JjrJXBnXTVhdhvy+wjOPDZsI8UP3A9nue5uBYdNsDcW3VrnOIBSdUNfNa
OZU9PcvdKlwfa0wyhbMa/PDdA09wRoPJBOG2sRPY9LnkYFaavhC+grUtfz7jZwU6
FN4mzRrwnnd9sXuehQXsT+XRXQyTFOKdQnqE9lfY+7IXAiEqIz5yTdOzsQtpkH7y
PRKSSMA6aBd1SHj9RY83jp2zKT0ZNdetPtfm6fjpWeTMJ2On51/r0PTURu3Vs8Of
xy2GGgFQX7zZeihjYyoPoGYcXX/+N4HP3jC5PBQWIke1/wTbbv7UEiydSL++lQ4l
+co6ky0S0ul4U+miOGfjwrXbZUA9jXGNiifwq1mj/sdCvXKzRBvpN+fZVHqWtlv6
nuyGmQbey91yod7owE3tJXneg2rhbiSlGQ22dMS2Qj8t+O3cRcqMPqlZlk4RQrE7
fp28GKkn4jFuo6pHHCMk2f9B0V1daatfgJ5o8RsP7ENJNXuTwBn6lpuoO1x3iEde
KBLm9Sb3E3xKK4aP9txwGmnL32XeBvFPYxo3e1cI1kaEWTgTc10IougiLFocjxwZ
APlrQHkZL5CBrw4W7nXnNyc4GQqP+2omPZwI8LK1oKO1K9a8Z3WvKnPT8SVnwuu2
mV0ssROCVOgBMBjbK8OttbTYvThGpogKuiAOd+opSGcpsRFvDVx9LZKz12FYagtT
hOf0s1lEfr/vwGaktCNBTxs7MtfeO+8GbQczSrJ1T7q0LJ9mGCzRWkDjfjfV3YZj
qR78V2mk0aakYOwk5AzvtXuUruZn+5HEooTU4CtM96QJhK3RAIgqxq0OoNb20Hr5
1Pbno00Fe4urznaK+WokXlhslmSe5TYuJ6419CtoAegDKsd4JGLMr5lqRp1EhETE
Uk24ib5DmV0HNPvxwc3jl8A4IURoZHi6RId1LbcJiEoat02qQ7arpqKPeKTS+sqn
BNFWeByQdFmocgdiNqovGxmyTn6w28P7ln8lZrF19gxlrDkW2oJ8VTD5vrriQaMT
CfFjBR9+88rJKkrRfO3VTBKawamO+LWoxV/nVHyicheHTcglU7nPtGjVs7aDQ6Cs
MnK9vZyl/M1mEFwJrouWbLtbSDlH8Sguz7D94T3FKnJI4oq5eIlao5NTLRR1gk5+
dokgvrBh3uRHpmbPqQnUqenFg7wL+YhYERFZV4/htQRIvygVfMg16pAivDnu1GN3
gKkCI1VvGlTWoqS3NWyx49f8K8oNFeOLBWhNAkCkBKl33Sk80PsQe8wJAk43/Lxl
wRaNdVUPyPlcWgAmRwkkoSIXnCWKLqmkR3GKvtU0+M4NeyfdbLV8yehVwowMrMHJ
gQC1radFlTSr7M/gwnFW1igZvB48c8In6NDYefHEMIfAeu9aW4RA8aVGbRfHOFI5
zeAyo7u8+WbshUpFqmihQG8NQyol5P7rXpiSu6V5b5fNe8aoJ+wP8ZfbItBI14nO
L72GQKesuXBbN2hQR/BCP4tSUNaEbc+biVIkxYVy/4x9lhypUtwJsigE9Uh34lOD
wGso5bU0Pj5WiQraJZXMZfLbKMWvKF2ISy1QkshTX5WWp12N0UehkKNi/TXhtVAt
K1PtsCs78ljhLyJh2G0BL01ULIzVvO+xT5wrsWGLwXp2om9Z8U+uODq8e2OtSXYx
50QlJyKRWYwiWaixdQcsMcKBXyAyJqaNMDg95aMi0Bzovz07JmOOyYL/XvXta/Un
NZ1eMjJg4lvl/NHZ9dxpVH0g+82hYRJjWYpvHXr5AWgm4oC90wcMIU5d+na7q06U
8IF5GIUcLLapFFsF5dR2gfGTyqRJT/zR9ofpAPZ6fZc1TVVlphqRrZu8CDlNcuPN
cF4oMIsaarNrNgwDg0dxjSpJhQizMO8+Fmp6rw7WhLaQSy9CzZ1sODAWdkneLjcw
G4nEYoxVoNa2SPthRq54wTFelz88IgqAI/cGmScwBAuPmUIHDulvUKd0dcpSivyz
K2/X4+L3c6rrymNESbzsJpdFcoYWuBbtXyxTRFhkt1uxFFOjGCmcjCvwt1QMkzbE
RtcUgScZLjovFaK0nOPZZ77eUkmxjScTotovE+by3SWcmJkcZq8eXvVpS1XhkCyT
0LntNUvkvQjr3UPfa+scPcE/fVNiwBCWmcctfO2hElMbUKHuYCybqSKQd1YbwHNp
W3hFzdYmC2H9ARlopbMp+NmivX/IPsGBEKRR4sRaFPZYKqtqUhXRt4hkUvZpQWTz
WeyUn/aeMB3PqgJMz/CXowZViwGBKcxOl1Dvb3rKoGpxVQfV4Kh8oLdbxY5xNVnP
wS/kAsjbI8CO98OKaaWIcqhbkPk/+XW8I7rQS4Ieghjf1Go0qEdMsFhvoyza8woc
8LXE/WdYydFI3A7nOHU09fkVYfH2flq+g/V5NDGy2UHpibRE6K70cOotQJwt6T7p
X09jABi9gprD5/p0A+6zgu7+gblYW/Q2GQp8DXobcLtOc0PHbIw0vE93+kpXEFDR
XeaER+8HoU1bYfFTvNa//6O7vWRDC1I1jSZiWP78YbZN/99rx5rNDCYF8b41jJc8
T9iDytjwe+5WrIba2wMmxxEY8xDwes35v8wMW6uQuqGq7avhm+4bHUieefX7lxgC
evwjsu8JIWd76Ib9TIRi1Ui6oFDgO1roqq2s/dsvJIAb358K4bgY6T0oQ2E68ukH
zwcUVjS21hYF31+A98UIss8Rj7b4jLFwTEhlYM8CWIdSFSx74cPpa41TGBQJjxFy
hj/MoiN4rNNC/aZGbXvUvQNnLJ3Jhl1sfs6/7ZEuJ5FN8w6ihm8IcajFW0ON17Uz
WTUMpvmTvqfBTlFNO5EUWcX/j/86vBK9up6NShQRF3SJwKJi/2c3Ye5MY5c2MtUT
EX4QBt9TWp1wrAxM+5LfQaOMq9fQXRVC2KG9fDMSYgX1I473J/FxkeI5DUUYb8gD
emD8SOxWU90bMjwgMgMkK73H38yaKVoDQq0qhbTtoDbxJ1sMoGQyXAEt9Xxy2VCR
SKie23JUo53mZVkQcP8yq10B1qGhWIlfAcBMS9raQoCPutmHOycre3bnZqczO9A7
VINaq9RZ/90S7d31t8jeYUqrR39pBDdPUNpJnZxFZjTrkJ4omMD9p3h/uUdWNjJN
6z/OiewAidu5L1aV4JpXANhXhyRC4M5f5FIOUXLGDTM8zfxoRYabXmANJDlfxJ7q
3fQuW9096h79Ew45GCF8W3609Jkp0SwkHD2eWssTeKXYdRfQnOLm6NvCLxVqkdFs
aISMGRpLJgbnoBuoxzyUZAqOg4J1uwddPKYAon9l+J5P4VynBLBejjZ4WcxBx4JS
9kz5pAk3co7mNGtTVFJBsjQwcuK8L3qz9pocQc0RTkxyATqG5cvfp3fG/PyuLkfd
7foqfsPQkOavISPAocT+vgdUItyhpGdurh9J2NxOSq1aM0OzC0Hv3lQWOscz26mH
2zbCz1H/Y0PX5IAIQ3qmlAoI3dKnaC8/DyEXCt78EtMKuzKeFQs9JvUK64dfo0ky
192qk0AIKSsWGVKuaH9z+V7ZxF38IfR8BEddTb+qQa7il4nL55vVYqhAevsqI8Wd
G/tTmWQlDA6H8sI5/RmeGF82MIBv1hcHcfaothFoDnsDZB5KkIrxDqzIJ+1dx9sR
b44R7syBY7Y1yfW3vH/UwH3AEaY4e99Vpf3n7lvkJfTi7wWWoapsY3XkCsffA4po
RQiWQN9KDQAULeUfK5V6opaFQoRICB9EQYDO8uCCXStzPhPPeBVUu5JXCUB6d7pF
NOGV+jnq29Mimqdy950Du2ESTVIVBdovBTHnjPGzeR5Fii9Zt04Z3k9wFgtQnVe5
ZkmudPYdCinGrqfaGX6ymNOvZcHfnb1irQva2a5fETOn3W9KA7hN2RAyoF50t3nj
CQ/86ZBWhG9LOJTu1eVVD/fBP4pciZR6ALDRqanFNCTitSAnQBpv6B0HQ1Vdzz2e
MmOOlUUq/DY81esllRUtSm5UbmVCoRLsXCnYvOTUY0qbiVTmgJpKK+BEHbjic66A
Zy6JtYh1Lz5i/uwFSYC4LBUhX1NgauioSmC8Vmf5ZE8h+CuFnwJuZEAt5+MyPBmj
6pGFKLFtQ8K58x5nBufvHYbCF/fPNZQMdtShV7ln9s3CTvFIl591F95GXszdTZBG
puf4hdj66jzYzZRHxfH/zn4IsLfoy9umdTbBPGTkL8CGRKBNzflKG/rezCrkj8GE
VhX72lh6nUfGIfGwE1MwlWWpLRYt+znUMaZs7t7Y4K/VRulhnNS/IbtmnqTaWAZM
IK4U/lu3Sy6qygAzqGbOvBkp9zlHnWSITPtWLA4F6cRc1XzSqsxNjRMhNu9kQ/Yk
MSQzmXzoU2iAXvnjIWRSfJ8oe4EwS881OHlLWBESXcRTsXJNiWsD64B4ukcoq8sD
Rjgl5eRn7WV0mD+m3o+hqmSAuGNWXpJNf89UEMK4VZoetqcFFeIzaj7n4fw4Fxrx
L9mzffvGhvDutH99/Shggm6V3PX8WHHU8JW917NN3zontSz8RCU44UOsCgYiTXqV
mMUxsaHfAQG0buhNDjHq1Whc3St2ApwSvPJ+/ieRxD7XLIS97br1nCrQpXNsBO6G
56xFO0wTlQdyPPvzrHoWKJqOTfT0aZYFXKOXm+xa6PhHae72K+3JPMjJoU2oLLAw
asWQ6Ok/IRBdgBQLpltV+c1SttlnYYjoVtxzSXs1I99o6ae7ejC/yIoB8sLCaERu
IrDokObcp5R9aEKn1TR8dfrXP89EJ4+DlI31ZzmCzOqZ9uJnvmh+JKa90s5QaWNO
MbBSkvquU8PFsMsb17t0obGjDdwXvb5mFIO203LLIfoEzRQ2fBJYmon9ETFRIqY9
znUk27ufmF6TqImElVNg59pTsmVyXcwn51x90sSCYXMh2i50mLjUpcthnkTj55RY
Cr8xi6rMF66mknY2X6950M8vsIq9UIDb5u1QdtOJyWAYlm4y4E+BNzvh6E1oGDxy
3anVxoQj1rg8eufSUClv9uNW1dtTtCG0maafEhaYtKaw9SIp87FoRjWGfsS6fquu
x00uUlePHHeGJHKD0cFCpofM6behJsnznCkMG5AKWtcotpKjo75Rf62cUuVjy2rk
3hoqpt+gxqqzk5y+fXcylWZMXEVk/Y++e7C1TplJNPjyoguT4vij63gbQ/OzSnGk
Xosk1NmeDTnJh4pPHniM6zSqu5LPO1PCjAjEY+J0d0d3gGngqZ7JIIAQ0o6kc6G0
wQ7ukruRupDXBxEli2DHQIKfEflgxgTt40ZdBViPugDYShbVW8Hf+78Sx5vWvUDt
wmkSnA2fIlpNoXjEdU1CVQ1aiIn/uzAM3Gp1SOlKgxeFe+V2ixb9fEwzve5+DmMd
hk7elU3N+Z51HvwZsDfOtt7NN4Jcauku/55xIeJbk+46W7IRKFSBM/EmlBib+6Vk
cRFeZtK8p/C2Td/Kfs9IolzcbRPNIfE5kGpPDVUm6MAzHDXy4UQCrQPNbunLU8Cu
0fR9xekLRXoBYjXrB3XZpW9jCGw1ro0v3o8N14WlTJksGDgah5fPWGoEwXUb58eR
AS05HX6hMsm5gOW6m20wf6uBeZYqy+aypXnX5m8XmmN+8B8WDnCV3lCjRenevHHw
C+VWRxFCR5iagKGdwEWZm9WyCn/PvZwK5i+u9UbsG2oOMfLvvcDnoU7WSjwjlGAl
yLAFtMuPRhkgsSx5JAW1eKcNRyIQOJYU6KZIRAMCs7ckgE7Y5gfZAh6ogvcomAmV
iPY3/S6iI/sFj2ci01JMcxlbqTokJ0Xxa748N+Y/WvEP3cwBWT2vpsdOWdF7yUAR
bbkdHvz29b5uXwWmi06citvgPnuRF8KoZhjsV9pQgzv6KjXH1gbFO0KhHBqOapSo
xF9CS73dWHse8FLRCq8ptc4vNuN0ZApMw1gSXTPuGzgLOTCjR7xfGqEzZZQPi1l0
lRwuTXcpu+bjf1CdH80af3nai4OZZHOMYUZApw9rHhqwCpqdz+QJK8bdVTvkYxbz
YGn6E+XqjtfGUogsnrsMXMKdSW/uYKF3+BMfGH9NYg4BcwcqT7yyGRmRka6ou6SL
uTxsQMt8nikWqodxj42l0bYLPWxdTPZoO3pfpEtveKENdIZyFag0zBcCLQg66XtJ
5EynpCWeA2fnH8oDYDVZOXv9LLF3BKbK0g44Adt/QLC4BVgSHOLFoYT4+DC1uYsm
mg+53CV0biku1d3Z2cGuBC74c66EGSqLuz8JPomJMHNZE8hQPRV9xOWAJE/g00lb
I2OcqLDZ/uaCP62DcwsFHxqOcb9XRYUpOwwGShOx5Mv811uQVytPt7XGAyChiSat
9fzBpyiY9tUzRwjxMbGL2XzWsEIGCFhqXMmokpQ4mB1P54zJyzdhVjjTRxG8eAFU
jdPJH/4j44zAUE2ool1xo1ybtw7fg+FPebm4Z0JDx6LOfHHzD3Ae55pDr87ZQKXp
e1f6b0aO0L3zLOIa3GlWGecHOz28h/NPhYtI6B6vuoDoixodSK71KpZY+i2VRUA7
/4jp2z2km0C+QjIwBV8dXqeQznjcpn9y87IjgZE7dRsDujSFCvzC8t3JSlTcagu6
6kOt7CxCBf41uNGKEqTequZLOaGWWdDubWsG34PBcFhnRpbBsKFw2tG9KN6hgnFh
V3AvOm6UAfcHVdbGfH5IXyjBJAfdf2IFE0GI+Z1m+ILYDG1gF2083WTbV0SBRq5y
5JhnB9FR3HwiumpjdK0yZQjjziS4NhMmNuyzDYTX6fzK37bv3qam1ad04UlpGQNu
W78aoUfw66M48UA89+km2XIWHiAVEap68/osB2n3F965DMWQ39vonjxrH5m3DN2P
wouUqOAVlpRfUVIJ5rWR0LeGyeBgmFEA/aF1Z4F9srd1s/j94Nl45zWuA3m027ld
st0a8dQZnIOx6UYPwcEILlFPUf+IIJ7L+Y9PUZpSxQaTHrR4W4Ikg9BMTsAkDi58
dAf0YJr7HFAwp5w3CO3DlMHp/yYCKkr9fFTHZ8jH6Dy5Cs9CXRN2daq3F9piTH0s
xaSE5uTOuxhctMci1yHKMrnqpSc7kwrBNVg4Zb+OsZH2JD/MbRTuIAn7vNj3v6E4
hEuUNNuotq5oOUSWXJtkjir9zV12QfGtxaf5fE/zXDS4jagscBzu8zuHZFWrbJOQ
ctj6fly4qq7ICe5sAR9svmgNTOi/oBRkpQ5s7pb3tIXN4LVK6VdZpMZaRIc4WcHO
6y77KxanFCf3zFMMEuqgxradJCv3KOhAAzNneGUonZvFy3J6kCYOXImboHQa8g/x
jUdqsjyZNjAFS1hbs2qEcplGjMvfTn6wyA6EAzecMisEyfdjCVroBXOV7Q47YIJC
IIPMNcAj1sr+FJPbQMv2SvNB2A9pUeHw2+s5G69HQuRM4u8Acth3As+i8WkoIPu6
gvzvmipRjXqJ1eKWsZbSiet3YTz0ApYuPRm4KUB+eH/c3a/kO2I+4YOsQ3OyK/vS
fHqzKzCLU0uGRJsZdSHo8iGUliAtpAgtUjovh6FoIaHNYMF52rj2h+schHubNxwh
8QWe9oSk25Wv179S8kI1mdA3IMnf/slrmCjFLoWXFtDXuonTpVZxzDN0hHDfKuWr
TcjSlOGJlaCP6gTg6tj1x7Jqbwe9VHsL5m964F6oTtIulutSXg3GGBGmA5XlLdDj
bD9W4nd/8AFlmJGA/MVscjUwM5Jp67kuZdhAU7DmI0tFzj6lrW9Z/egit9ajF7L7
n7WArPauiKUVaPhyp0TO3ZbTwcGI0n8Fm4joAeRWUsco82/HEAVlr5FDTLx8U2jj
EiGIMIR0tsF0TL8rsGnnB0lZ8vT3TEJlZwSCx5poA3pp3W77riXfpsKJFgcJ5eRd
rg/g5d3XOYTK2du8F+MZ85TpceIibRYG4xVuz8PnxegG8w0VXrAyBIPsyzJqCJb8
jQWlA0yeiXk+VFNJqn5Q1Y97p2xnXTLz5jOUgqvybwVI+zIxlJ1pFkAJtDQ9abSA
JbdoM1Gk1MOA2gWb12WtJwKRQYI/AdQiwJkxonc7muKduM+JI+JMZ5BTwKEUk8lf
OFxEwu0ZDCyspiGNqs836VQjWhgMsHWq2GU4SPT02Q7SCy1rcR8lvz/RhT4pdK32
v09ugb7fFmNqr1JffrA766lA99Vyw3OuP0CG8spcPi56bb1usmG74wJP7xxkP+74
CnB6b9gah0L5/au73fPwMFeJQ6soXejOiMVE1SoSf1ViY0/7ylknbgQslgjpcOBN
OT/ueh0M6LP5V4b0QqhCLJDjUz0BonHesPh2/1zpBKfwFOTy90UoLYtjAEyGHxEe
KKZ66fqflS0VsdyQ2wHkNPrBT4pbFu7j80blHUa9ZQZEaifQnvloOBdpJVXL8tTa
chTO+PF2K/hyKoVsGNjKNmZt5kNlWW2gtANY9dIWeSP2d91EF/PWlMl70ZlTtofR
grJl/HINjELK17fgs2i8PhlcJCcTAlHEclHM8ldsX2bAd0Nku+iPzzE1PUU0ubxI
B+XtE83RoPWw6imEueZaqFY7Fr6HaxwsOxGaA+t0tNEAVRhQPGDzkFfD7cC5k96t
ng7INoaork85zYNrmT6wGwZkWTT2C8b3Z45uWsKJug88eHS8wuVEjRcv1JwSLDkh
XPesYj8REDYPl8vOKsxOEppICxXSZJLb6Mpsw7jJcezO6is1le4WDaADB5zrqXNI
Z9NeetwQCrwDcqRuUWo0x0s476J7o633zwbCgnk/+VaiAfwNVY/EwvC+lgCjSYpw
CJINvQCUTjKaKnRb901pXG5sZcXnhTR03uSo8QAz/1b4fCIctehfz0k+/0z7wxJv
KdRaLQ9o7qNkM7UjLZOVn3QpBukL3EGuahIrhkThqQ0TwfSqQjfpz7qVWpoqJQNP
2DkEzr8Bu50sdUOnATflpuToVOYXqKKRTytc/lxN3De5k1iuaAVeh1Ip3mwoRlwu
7AsgSpAhI9g4woyzLmRqEocJdO6mkR1mWfFvuoXctOfkA5OCJWmseZ2snS2mg1np
k/8lYU6OGhoiNrG4z05HIzIVylF49q9MYcKqEWocB3oo6bF7jhA+cwB5CY9n5cUv
V6DLYQbcEVBVK0Iv84NuLLNOpoxpgnXTM3ioaiMy+AeeVY1gi91M6eTRTyJCvvl+
HzFwAha+6N8sKg8+ont9yTY8QRSUoprTfgjIj2/3SvosSaqUq2q2O5X3FSghwRcA
eUlspW5mvVdFdX5pRaCkkrLuOa5hSsIWICpXIbGY0EP6cN0s3KMfhScTvdHfZXS8
xMF8KkAzT5lbM1Qvg4qPg7UGEdLrCEyU+HBbJIg/xDDusJR+MDTFGGDyNz1OD/Ak
l7D5VHOeWoKtN23Nq+OPZeE5DQMMXN6D379ndf/dqn+oBaCIL3MWKoUsVAXyM9Qv
VchAqdgJ8dqx/m0Iz+yEDxyB0UiubJIyWMnFjBo1rxN8+yUp7KvUc/hDxwawCz7y
FN/WbEV+UIhCsUPNTOX9oKZYx2/bpUL3EiWFouIt21rMt2m6DjtblpLFf3iE1N2u
KOmTtOGymEFYW0aj9N4Gg7VGb6IfilqT3tQSn4ena8Ozoef8wZxTXgBGN7QONeP3
o4J2hNjoyr8iBvyEc3N6iU0+9vjfgWrYyz0+SqSbSaZaAG4X+KeCvIhyy4S4kDza
Avuk0ubo7rOK2qnGGhiLeyGbFvolwl2lLvFZ/7pVX6PNXOHOkAz9wBKRk7LjvIW7
kcOAQ4CBri0vSxLPpWWyyAhkO+/+2+QCj93Wg0DcS/K5clMqpqCW+9fRo+hO/y8a
WITY+IxyZjBKQVLHm6TN0CvRZCVW61ddw7ziEuQ8IHmZcy5S3AQnP7DP/PGfabjL
FzglWP+1X7RBbGBXfqkotTTibTsotKC4EOr4oapGO/AQXvAzARfvuq7Mbb8mX8i1
370der/NtwlEHkwx2tizujsGrpgNV3ScFPba84lmgiyNrlTm7TbtdMl1J3ji4AmH
WRK5ANvyAJ5IQaT9+yrGzlr57b+0u3FxIh6Py1D7uqX+/xsm0L9SsIx2QzrcNZZg
rLjBJ354DM6tC+jLG+FLO2oPhwoi7U3zvMgTPminidiCIj75561Cz8zXD2y66NwG
RxQ+14G+uVeqT73DtKaoC3nY1OZRogh4HM1ohuE1UWcRhEq69zHOc8fHd3mczBme
Zrs3jXUrjZTkSL/VjdlVRZ8Ko1+KmUAibFR8G3fYtDz8Ywl9SAM8uJbo5vq9Hm/j
1klDwHyikVv08S45j0PGJrDuUygbPvQPs6Gs+vcTdO+slI8Nr4DFhCSQH7B+PT+C
9fvdP1ME+8RQ/HDB4essrzNc2V+hIhn9NfwbJIY9EjFzJDqjdp+bsqsTVvTZo3ds
ZnHVCh5BZGfQg2ggIQ+NZmNU11g8CQQ0smrWzqhi/kS6QUjhybdo/6bEsfECl/AC
W+AnNwmyYiUZB1Tex0AjdVPLMdcjaRV3pC2N6a+ZWynxmjFOGMk0lg3aM6zYWsZp
k7s4/tRCwHzOmDfCXp9Fso2b0bozHfHzkPdgv2bQwisiWuB1qRxR1HWOna+1ngvx
j7MZsnPCL70hHJ/Tei9p7VccALLG28CwztSy0XG1bz1dnrphzVcktaPO93LJkLRG
cs7xcoYY09JaPGRA8k29ic1aserCopQJW8oa+c3n/lCtueQMJRSbN/L6g6dRB1jq
P538D6fz5gXSdhba05WImIuMjMdJ5BDDk7/NMrH8amfuKBluOlLscjdgAt5Covsx
tWBYfw+EJNpAywox20z1P+V3nvqexDSGnQuJVntCf+tSRbMqFnSIysf7NPoIDOOZ
YQecz/E8pFSy2oiCGpbXK+ZLeOW/zlrsBMvKAND/291H84PTDvayfsmPVp1MM1/A
Efh0R90neqvZ5zIIt8jpAKKPsNpxEfQOpnjwYIh8cvp3PhZvukOTdbvdfBJSFTra
IzE8jIDJ/OnpJod2pn+SBZ4tQZFMc5dnZnhfpDFdRUjc5JQ5cvCRr2398p69Pjra
1jHUxi1avlWAuDpXYtBgbVIMAUC5xWYyert372LmCtgJ89SwidP4IUx/hkyIZvI0
hfm20fOEN4+xq/bhF54AxA4WlGcQWlMsN+rKI5x1GzTTTcVDlmpU/YSHQe7ci3N7
seMC3itklQ8Gj+9d0pMzuG8ivULV+wMYUv59dJLCzEVDjeA3VTvvaoQ2kqNcgoP+
QanaciWkLWhzVe18S1LenyaXsvcXLxFTLGJIbQ1Uk5CwjcJYmoIgsa/QN3C59lHF
/9GMks5yMBfimv/KyB/jKy10qmMDoXZmKecll/gF70d5oNLmdmQF/YoiEO4viq46
IXXG2xOj3QeSFO72V2SFAKoWdHgL6nI9gqev/XWidTLuhEyUnE+rjnZv3rLO5y8Q
NnybipuLi6wvwKUy/o3wbioPLClMC3scOpAhDxOuoOpL6X8lRiEqtkmHowQOpoXv
JWdMrTCltMu0s/S1EyS9hM2Ccl4a7IwahEn9EsF9V3CZbLOsvjn4m5DBoscNKRWQ
Uun3kDCTdQcxzOgkWJe28bSfJAyRPK4iVEglySXxyVynfj7o3KXV6SIcyFu2Q1Fu
GYfZNIeCQw368DxAsn7jLAC4RMan9lbR/+SaRzbS7gKvOb0qaNE7IbfBYt2wzEZB
hnaLesbb0Mrh2YrNBy15MHjScrGh+hieOQ/q0/pOk9mizDwJvjmSCajlkBT+0ESz
8Ao16nU4e8T9NnEvWjDyR2h8Qwt9OeNh26I5Nq41cOtkVI2ziR2Y/Sc6pyBHxRCD
51KhYRKLBPRZkEjUpis6YshH+Wu/UGmMLLLBnw3EW++bFX69rR+3sOA9fJUY8BC9
eEdJWB/P2r2dgh+82IwAoSWFzwhcPLrSbBVkMznezq3JrvQ5Ft2+J2rb+L3VkNfm
zbLaVZNEw0XboFOB7pfGm2p4T2mouvFPyUDjhDjdTBfRycJ/ctxjmvjtuXdyU2K/
eLHjXJuf+/vIhztGzQO2MZcKiTy+chDGyv8MEpGJMg4AMJe+S/rDDp6lQr3vPcTf
EW0OAkqILeDWXq7jh/gzxujERBmQoPHv5v3l8FcLLF+bJFj8v5FPE8uRxYvuPYnp
awmqc1rsrAykZDQtDMb5rwfxp8DKHRCs6shcvQZVh63VV1AtGNrO0NSORWacz0B8
z35YAX2S5y1b6ymKbxJHZDrEuzLs4W6G/oUL5BbOnpSzqkhAoxJJza0c6/WifXkc
HCP8FSWxEG/1UiYy5f6gkSSNDhP+CMMKStczUR73sRZOJSqNfv+pq705f3haC4IK
0ymzJzcVBWcpGXsS7bJQ0IdLcRBu7hk6vlG1DYZN+4TvSAtyaHIqYdDTCuTnY9lY
NuZ+icZLqR2GrVfmBahyL5QxWrN+nvp3HVLd/Jme919FegDp/sKwabi7Yq2uNRPy
Fe0/rYpEjPcEAcKoNQeY6E8QqxmfV9y6iQXKbeLd19KNOmxrj6etoijN0qbhzuOd
YQWIW/50nttDgTU0tgnALjwB3OdXg8TEIT2kwYRFJ2pARZ0TEilnPhlzXSixUb1n
4QKlZuiR8QvUpLZL9xe7QyboQR+QArUo8RfG5AUJBQIaT5kvFRdO/EhvoRVesiyC
mJgQQ0D5qG2IcJGmSBi7OuIgstahiNCI4eAXtwVhyIe6t3gQ7OGc8w/zrrXDxhWO
msnWUXg0NELQWjyPZsT2kilDiAkIZq961pKsLU80zvhv/VrZMKvba4LR11gYtmUL
dCf88I/R8zttAXB8vGscoJA6vJSmSAPAERz8/t//ztqO7D9JAISMDB8j0/oZ2sbB
o+fEIKEZL6zObeLXJp72Mak9Ppl8ZFOHw1kt/bgYqEeFQZk1XoK6SKGFXsNs7345
R9VwmWPQQmA7thyO9HFgRWMMq8sy0cFD3U4OMZnGY/CvDnyAjfwTFK4OWCT1Nm8F
U9h/0AkB5UT9v135akUOnzbCnPE1gIUR6EjVt4f2AM+Soq6YJrgnSAkb9T+KymDR
8oniHkiRAmdqGhfCBbcbHT/b2I3wzwn9DY5zJixUlVHIgNa6jMbUZ5yJueMbz/Da
jjo0punnZ2hYc6XWTrp7GEYdLWaFEz2gnbN9aHHRIuIoQgLNnvHmjv6DDC6stXfx
lq5uplcSOVBEr5uT/VSgN0FuFWhJVVjtSxiN2cvb4Uz8Yucw9Rus/JFW4PdEIDGe
t46sx+5/KaVTB4i4Otic9do8jPLGvHNKxmmT8BcsGuBMIvrStmtscojOF5Wy8O8E
3DCTYgXsENy5/XvQyFghbQZIyClpm9iMr/Jrli+zAm8916jNJkRtvEyaCJh1whF/
Obn0jTVbbvkCYIiybSNwfMv5gUxGabq53F+mpYXJw1kvV3rbgwlxESHHfXcuvjqQ
tkjrYzQqgRJa6lGZ0VWGSbH6lU2Y2XD0IJ02mm40hbuKQ8dbbIy2JefE2k1/vhc6
l8iJV7bztdgnUkoyoI49sld/Q9357CR/SCu/uxvobW/M8d1HDbT2zaII0xx+avap
wpvGKMXE1CV8XWzF6KjBIiHQsVvlBIkA3B3Cnly+Ok60c+mXfus69+YgujzgCcMb
1MXctu05y6IDIIF2Kmb0rCS8hUtYfwglh/x0FZM8vMEdBg2XVsLkG76bXYxPMF3I
r0PqDj9RTF4AAXEs43I5E7VfUIH02jln3UGauo37VD9zJ3FHfTMpyrWeMj69B4PF
/7UPj+9ynASRuKOvuEXj53aixN5ZhhKMvjFkCghxecIv2WIfYzvN09iq8tfCZsEv
wCLI2K6BqHACr/NEquYuDr1t3oDREdFO30f880BpungYnw/wDV2/Th6XSYUdI8SF
8cgLYKCwUlds1lW8ef6k2Gv7Tj0eFN7hjwtE5/vaWokliBsXi3hqQCgAC5glZJzn
HNYxtsTtKmEFxzLHBMHzFqkEW0NnvUx2FBLmP70kbdTvXQ1q288g5tXXgnPHQYKw
zKT62ILonVeKSwYKD2tfAbEaXxWhaNS6QWG9Fv96RBqo4MoXD3LVOPiPaAWXyrVX
6s8oN1EaSEgUVqQWJmr+wNkVz5imqj/e8e1YzZjTdGgfz+zZNxzdi6n1GNXBVcIR
mUjTC7NoAX0kHBgYsdG5od8m4DYDIBFsMMd5UZA/KI+6Q3yb4fbCIe7jqGoIJrhB
b396RujKENx7VgHghGavrXs3ZwopNxvxHRdTh70GabCNFDRqB72aqwNmo54ZGV67
qWcb7eedEJcfVAYNLC2aNj3r4ZJNLESnoTZzoR2Il8RiwVXY5MEynd/PWPUD/mgB
R1C3/bk5yYcZH0k/7mCbZjHsAy2uitOP7Mpjkwcc7oc4yFQKITXDTH2atV3+4S+y
F/9FOIrrOJtV6heStgtTeAr1NyF4imONFn+EsT4e0kwU5o59geg7UJkoEmR4z8kg
ZhheqENornwV9PnMZZh+VWxLaNJuNLvfWYXEA+wf81E2AKU6WSIlujT21E4KBlng
qY+qTT2xgLRpTMQKjNFbgfzU5w0sainoXp+rc3yTxd76xaHqfvMmrZr4EaE4s5s5
JE4sxiVYw6LLHsMFdi0y6UHE03AmTCfBDEARcgQkd54uRjv7xh1b9+oqAWNECG/8
/QTu+lZoii9Ss9JB4rXkT3odcIg2t6Bn6LneYWG/BL+JjGsn+A7MbO+xZxpmDXZ4
ns3FGoSQfhE70jDsW4zsRvn6CtDomcUoGhWKUK+gpHpqzmwsaqiCiUGhZsT/cgqv
4vyFZgJ7jfv1jtx/dgPTGyDsyQ//xs/w6xOc/WA5h0EN6VRXiEmqdbFfovRZ4Tmi
/ZTBDucA5RE9+5xVl8JjV1uQpMXZSe2MbtKfI6GX2Qrg3X7ODIyPGK95PrJGKLX/
+Q9xpPwophPDoIkHo37OwNkKBV4FvFr2fuQcgPzX1R8NyUtO/4H9v0JYclWwt4oJ
mf76+MBwQCD8SANIpx6PPevKn6xp/HLeFGGv39sXCj4+NRLgoth67efEiusnTgbT
ZWEF2qNsR6OgZdHhQlAwBDko/C1/x2GJnF7TvVKiVPAhr7vkPlSnWWC3XnA8wHo6
qWbepi/UWQOEqN9vQVTq7C3zvKhw8LwWkgwv8Bp5A/T2TdzdNppnafusyNR4yYbo
bmfTjxwsTpCPkTr7jt+80xV7kkiFmaRok+vb7U5SNg7DvF9KfUAqMJbm5oxn/i41
ImPDrRYw9I6W7r3shyNtLxYB4SdIqvQITAXUs0Wk+ApmsuppP2LC4PlpYpJYZYil
AuAvSqkxAUcQZGnKJ9Wg8cJ0W1pVSKgWjcjPOp3X1JnYguqtE5T+pTTjJXyeVNs0
ErxqMBw7ybt94vTfASxJDQu2jd8Wl8Gw8p53rZy9ZpXypItDcd6ZMg54adLP/QGW
TlGbbTYL25+jz9bwVPsHULwFCKlgHRyewCeol3eZkJy1eiFrJYFa0srKNVevGQ5G
+C7JNMoqOy5tNsKSwbJh9QnGXRVKe6h239IuS7CNBVy09bUF/kLIqp/bQBIqS071
AxOQcQTPiPAH+uWZz2LNT8PwcafcRNFKIBGodxl+tJefW9zDJha1MAigGyu6f/+/
8/B8cb2TvclLryncT5w4qq9UOqDxQidZY4COnVPZoBCGIPnggtT/nKIkoi3SoUfm
nL3PaHllKMNqxFZqH+UH11Ymt7LY7ujJ2Iq/ByJVLNJEWj7MhzDRVHlnP55oArrS
AmIPfSlquqDhe/nVeAc0YesBnkj6GUfFX0yGLMdNKRKnaEBoG3ShVWr+kw78QJWq
ca4vcmfQr6Bas6h8kDztHXJ/bKcIMi6c8+fQD0k1zo88KJ7MEf2uQTEGYCECe1dh
TsAsSeU39QBa4t0MhEYNCIWXoRdohsoDupzutjgEMn7S3yixCCa3SA6GuSStL7bD
Xa6yD/Q3BS+eIqMoUSYHSiCHttxnDHgSlCce47/Y9akfLHbrZDm+N88fGZtJ5QWg
jrXKcvtKwrbTW2Y8AtgJJ6NdfwFyia3maua5w4GcKGtPo0okYvCYfSXw9gPfO3h/
YSN8FYUk83XGQRUv3xi2u9V98O/5+YGxEQkmhNldbYBW8TMx777FkNgVub0kgv+N
WJqUGev3d8rCcmnuUhIzw18xlYhbhWqpetrcfAYxEjIwphzQYW52Adk6KiRr3T1n
9qbZBymhR/8Ubvb2NBTB4ubNVV3Y7JRhNk5zVdxk6jRvfaXptRCIIT5T9zHDpaai
hSoR5iborNvthqkonybjAtDevC5GKe+fjJmzvPEGMNeoFEJHHMZumxGp2CXTvr1p
/1iMBwWCDzD/5j3flyoB4AhQAHq8mbeB5BZ9IPN1W+1vehEwagJwCnHiCgz4H0BT
E0GNr2wIYTWxiGZM4uixrGIF+fef3AH1eABA+gfMzBorPC1iclZVWHB0i+BAGgcU
`pragma protect end_protected
