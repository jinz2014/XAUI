// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:45 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rQ7q6kdOojuob9lgdK/0YguXxkNNx7wVey0xL/R91oPT4DCGTVvJIEUeN4MeWGYC
GfH/0vhGcLLHgS5YjAwUwzA5FfeWqV5sL8hfJHd/OPHMFYoIEzzCzSSjBXkbuyhv
iZz/45raOsHfPQZ9O4K243+WpAYgXl1+oNoOB306Jq4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 54176)
XrcPa7DVftXqjDhFPYWXOjk/YwrWosuIudaFZ1MKvFCKWoDx/VdMok8laPg/8Qb/
7bu4wKcqQFvkWDWsDgq/ObWH2jdzwengz6RsJrmrymNk8NTbzP2WVIuqi2Q7Jxu8
JOEbKXrYXfSIMXq5OSAPID6gDusIsjeNkoXWhH51dl9hYqR0XGjdTe2OzBfvNlYL
GS1PZlW7FqUrhrKjHeYHGFLt77pWDTQZDaRz8r8KNTxRjKXZIrtrBcP8edjm2QKd
bi5dwKig6yr8zUN/vTvtWrIcrmhDg0QZH9Sd54C6ETCw1p9TBgMlC2PyP8WUODlZ
UwTynrrWjZDgLCnWBWGGukHriP/eTPM0h+gsE3PBjIGtA/INgF+H4JGzMB1y+0II
fhWB3WaqNlCZ4kBTW/XQdyj13dxmgz3ksHp0uWASHy57r8buhFcHpIrEx9yDkDJT
FzOC0geQJR/AEtjY6tAXWSjkYI4d9lTLYPIxJtC94Zeh8ptr118TYUA9kOkDDw6G
LQgTEcebe9Ku+7xyTfY/6d/RjaeiWeT1rsFy+dj3zbWmIinWZyS7pbGJS7OcD/WT
tpqWsO/L1g20J02FSzLk9a6wYDhzbK8hsxYe5q3X3gJqAspFK7BLnIzgi8sS/y4w
SPFzzMj0Ed/537j4gf96NJ+NNOomE7SyqEp0E9e1bm0WC1itla7G+WXvrmoeyUW4
hAP6ss9nwRz4Cm9cIg3Rv/BeG2kBq9+rniLuAnu9zPsT/5jTnmH2giiJapZDX8fM
mBFqHi6UHbh3lTjwLJmrllzNhneD0Y2eLYftxeuzbgLhKd//1mgmUOAYKLJNz2OP
pWGaJ16yMzMv8Sl/RTfz4rKwYyTHx7iPzKvImQ97mUIbPouUahNIqj6viICnzoaN
1jJ+KdC9pe3hSdu19Dhme1CuWL35bux6ktclEy6B6GBch7fZdi2yYMe2eubNqgT7
bGGxsNrkSYS3ybUvpAoJvd/R8Vcu5ZL2f8dcgHsvzBnzeO8den89ZojAvuMZe1eQ
2FjxVrZrwgs2ORvV6F+UDgKiko5Hm1iEOQUbw3V4AZWFEahow0A8ZTJNjkyMdBrF
12olaizQYtBimsY3s56lxTxlXDbedbxAmrUXmN1cHqYtszov/75mc3i1o6DwcYmq
Fr3YFuHwb/XExhkfNMDMmq/jhqfRAyWVh+krjUHGHPJMl/96/X3M3NkqBUg9LeAZ
zmPCr/73y2GdKV4PdggZ4pIUc2wyqBXoacIGW0uliitXCX0oIDAYgFXdqkmNFlLf
qesDcADl7QU5oqHir4glFNIsiP9AzK/snL1RYFDLW+anExb6p9yCv2hHGysDVl9U
3a9BrVczf+JxJQ5GryNaECAPGcHzWpSems2M5DMckPBQpzkL4Ho6n0aO3Ti6ZSs1
D/dTS2nOD6ruyMxTjD8YvSmET7FBvwM2JLvdo1vJxLm471f8oTqqumcumaQn0O7d
IX28ddA08GUWdfkTQ1wun618KpXxESUwfqJKiqJsobbWHllMDxZQFQKF40uEkZQS
grH88+sWcLs5wNjqz+RbYNNzbyhWiFDWg263AcEMNO+B3q7F/YCDNnT3NL2idPje
aQSzsE2VdEeCub4mR3ViBVKXWRzh3VTcz9rP2flVAmfssvWjySARY7JSfyEEtSyu
JS86hrmmromVLPvRia7u3+vfRlypKsnMZX/1cbflus0D6qEQXTcp3J38rQEq31tF
9nuh+UCPEAkg+pWCmG3pTsTBtbkL5H92SDv8OoLZlYQdUB9S3TT5sn/jkDQRCRt+
+KBQADQ/jB0jID7rCqDkm2Y3h5oMkh9yLdU4xPc36ZG0JT4nZJV5o4NfxZK6THuE
eYRVhyjM9pg/e0W9bp4Srm3bZm68l6xLDTeIFPFm9iVu4YnCcqyedT4bFW5Nt7zK
OMW5PCEJoAaAMhDxLLefbZErpzGtno4/1vD/SlFvyo7C9LZvNDZhCuMC5+Ys1+ne
DQIrPBlM3EABv2NK56RUh5qG5ovj/UhVd+lV23hckopWVKHbRiv34Hx3EDwlIYh2
FIJ3bfH7wumyS+eT1b7dot7/JyE03xACj13KGNmMFXE0OxoffWCzMrMGKRSuMjoS
uVPI6HrxtWuhbZIsrRFXhDU6f/37D4r7GKkmAd/TGFVH3Gu+ALetbfk0PU84XelQ
9p343cDfTmpgDXm3Qua5otsGvthc0/Kyb5xHt0REXiNOjU0b4jRndIVbpnfUXsA+
033d/YEM/ysZ+q+0d8jOoIrkdpSD4YEiHSYFcUzfMMQo0bLFaZf0vuACercw5lvB
6OGa04/BBGUdr7fOPG9WkqIxIfkxLde1r4OmvPEERDnKFksMLxCRmAVN4b39j+gB
k3kpK/f/KO/gYTEsmtuTRs3JAy8Pd67Aw31ShJKwUu+rDwp1Qkuo1kcUh7J3zHab
FoJUsMO/AKXy3In4iLV1cdvnAVoBU/b23PqUFEsff7DzxPXe9/ps/PieDWmwXt2W
rkcnvMufx0/SC1FEO2i7F5k2Y2KpVLjqPBO6nf0620LQDS+jom/dWqrMNrd3MsHO
PfIFW51YFBdboDeOr1rhJ2/ZsiNDXto208MtIvDXehZjc6cSLWgH6lfDaNcajnQJ
zx13GM+aVSAw+Y3pikjZl0jedo/R7TkQGRpq1oBXF1tetqJ84tn8sWTB/+gXRbk3
3kBzJTTHOH8fA8Y+tLg+XKB2SrpVNWzqTOORQ6O3T1T44ZVQncNAn6C6WDXL4TOD
N3fqIMq6JxlknU8VDw3nNCA4IP1rNkvoqwu9FMK9urPiDI48h0WtnuOLTG1jEjdx
8ZQmId8dBlfJx9gKxBNmHYPgEXleL2S9YKpZ0LmIk9KMrmRqa3tnNEEpLdvY9utG
1s0dGMJT1t6x1kzgdQ7W/p1kRi0i9u2UzUWYe5U9oZ1fImO+KLpZ39bQfnCIZePM
/qikza8B0kfffsnEcSe4+Xg83+TE2aRgtvkyzievqK8cAcGI5739CJsOd1R8tkPg
rjG5uws5tyfTglEe2t0NjqtKr76ArCKU7yAPVu701OgG88S8CFknVgA91DjpwQVs
bqkzx61ft3TLZavZV+9tZojHPn68qkSCel7fywV1k6U5P0tqjiXw423RC294OljI
Uw/1j4oARbCSdi8mFYXmcgcE0e70DDywkcwlhdOnR37Xudh5CZWEkKhOggtkSCjE
dvjoFJNON7zGFJfoqS1BX8m+xyD2ezKNtFQCAlYo8OFbxW90O2tShgdrlc5G7JbS
tgh0KJEtByS+Z4Ef5Firge/M9JJ+sPEzS06e5u5mWuLCT3AIH5dIeNaa/Ch3HGGV
FA/FwC/jpb8m/guTvytD4qnapBYvcx9JqDei0PUJgpuezdac0mgBtCKD355UziNv
Cm0/q2Nm/xY2b+AiHkx66Cc+5E9qzY/XaMndQxpgcQEzSyTvY1Nh5USHISmzt19M
jtbm0m4ulq0199nOeyIAUYvKtZw4Ofv65ka2ZZOtnXJ4r28+ZDmcfTrXHr0A9eW3
i/fmYFQxiTam0Tnq6AmmGNOwiA1AkWGmxRCX2dpZ/oeh7kJmmBrTzXOus4qV6fJU
9On7DDn+qKuRCEDFsJUcSPgNi9fTs7HPAbTyI7zEjj6R2lg8EtQBpKhH3cM/Kk/p
A7BMFwojVVKrNuxVUMX+dko/XiJQPdO/URdww/fbQegO89iJLSnIIQhtN+wSJ4Jb
aiRkvzNEMq4hbJ/3Zfk8207mGKLljIcbaDmCqyCtSehSyrL5iKX3FVcJAvrEkjY+
ly83VPDK4dB88isyXOEQmUhYObX2TDXLUg4GnXwaSzBq7jvTiQ++dyFsD0/hsVkI
GAXXSLOidHqkMb4pkNex4rkzJUBB4BZuhO2NazgXYrAWaqxdQnmG7VpYBnAxMsQ0
bYkPAQTs9CchPUhk7ciu86A58tawxxHmT62hvl+rYhi3B6t8SaDM2lMyP65jza6Z
5njNaTGrSfgnBzlksAzurz2rzOCHdU0pHmiwY8ojsYtuEjaIUq/xa4KRwZXexihi
pRndc4mrjkPGnQpt3GKLL3p2gkYbXVtBy8fpBnWt4+NvglMi9wFIa4uGhHqKnzRM
rhZCMsS4cwgxy2OyEIN+lvVsTJk4QFHe909Bq/1RmIOJDttcFROHCPeqMGvvFNrc
JyV2BVoXskFACEx4E8eVfqivAfX1ry9d8kV4L0xoReGxvxV0punA4yThWmv7klj/
f+kv2UXxq5dcaSMole+cwOx0/6Sw+fjqKrCbw0/Weve3gmLKqvRUKPEfZREhx4MM
01mRuj28boFFIMIYOJkSYveSWsXqhXkNOfdeICdbiDXCNE7JChvxJmfJe22YIzqE
9W2jx6LAOadgDPrbftZ808nTCImC8p3a1H80kcYFR1xYAiGMHYqZu/OoCGpTYOwJ
go+jpJfTBdMzlnJGQ0CWyh0bpp8IwT44s4032kYkrxRkpH2spb/ERuq1gllaVOdO
eAfhd3nBg+b/DvBQR8o8wRN2oPk2TkznPXI8G225TeX2byQD6gynT5Z7rlLV1Ies
vsQ9Q+OW0IcHH3PTVYv4Qc06iPt2AkACkL+Fo1jUbt/lTdtgZrcfSWrYnES9AULd
BlYGl3lXEFCiDl6PFfw8T191Y36xWrzjgX98I5oTn9sZ35r4vU1EUmauJ2+H6G1E
ykLalylG3cyRyZbjQT+VTf2s2eoDNQcRC5H/p5yBvxZOHMFgXwp/9gaaxtoavevr
OBw8PkRpTrrOMtBNQ49zo67cyMMuE7NgfmIg95cyjGgvK1ec1pesdGYv0ZkEIZwn
eM8W4+7D20GAdcbx92G90iNRYXjrIYFavbSORjVsytaTlVMNOwF9Jnc8avBEE8MP
kph9psaYsSLQ889DAwugOJtFW5gBF/MCW+0N8RcCE6PFcnMeQ75Yyi7zH28E8wzq
GgLgC5RPYnEwMfuOTTsQRgUyUGcuq7IXXo3GET1BGWn3OFLAQ4u0mglHQpSqZV7V
HHBw7iRzJem6BuZZqxDAFNyFA64X1ZtddX7LbkqJHbZuYd4C/RtfZ8yfn4f4MsSr
8ytq+slZdRi6P+VW5JRIsj/vQo6Bay2v7U9p4LQwrpbP/p7AWFoQgKICWVwUKN1A
d8XkAlSH3tcwfV7Qx8IZvQfSbichFiu7pluZqoJoVezjaAjmSkMI6Q8Ve2Yc3Qvr
Q+TVbvJXqfGN4Bgg4tluN6bdvHSQd+zu3Cp3cOAZniSqPDTp7DUU1uh7PgotqBXm
ROXPKbVqPfLtRhZOfGCAWY01k57dYjqAaMuPUzZb/PxWa+CpxlMQKlw3caSAcShb
crgnU4pGOx02gGob7e4KHqXEio0SDt0gWmQlDZMZhrAdgxetbIViUioihmLcTqtw
a04Iw8Z5d7seg+zfcdHYb/RZ1e9+MY2RZ807ypddrgkzpJDW3orMkbvJSDxQPRZi
1TaZugVeDrnCRsDTmnqk3FpGIU5Aul2aVocQ+wQLnID7nE93bEq1tP3Ww0PV6soL
VNpXjZodGJpjTELHuXkhXW3aHpNzusW08ecU9ZsUw3nh0ICglO4aKt0zUr6dkgSY
tKJQMCnOR3s2RVdsTJegM2OXbZKw0aaQth3VRYILz8VSmnu72Oy7bxoyrsb1u41c
EJ1aqNU6C41LHkU8x1ZGXyXfu3hHf2uvp6c78bs1HPGtsZce19/ufPG0M3XW/6ba
6O/shWfKyFHGKk49HKxNbzWwERFe7ISeYYJib3nHjyMjQsuJnZqxqKFmXk5fhEPl
8wzAbmxZ/1fDgt/wdgZThPunGbVABqD7uHv3HRvT+OmvhT7PPFLWdrehIfxvvie4
n11B0vfVFXs/wCrfI7TOxM1fGBqJQE1Ea4Z0th1up9HxRAeqcAOiSpl3HnckNEG5
6KJ9V6Bifd8AvFU2KNk23TAF1ILG5mNIkvRtznct96OUC6k/yOiDK5FztyOqEAQC
VJD6BOPVYCdXssLlkwNKJ+LegjiAqsta23vAxKtP86tfkAqGfFn2zVtq0k1N+wRp
xq+IJEp3Z+2fuTXaWIoWnFTsu64lYGmDUBNs1FvZVP6gX46iopgRqwnYhpxGrpcz
DSG7TFmP1FVYXIKciQ7SP1JbRggOA0wNMNp/Y3noypholTQlUsFp1v7RARcDwqPG
tn3AF6lrFZr1FugRn1qI7VUjBwpn7zJrxpySWVJ5ck3aVJroM+PpGiPoa+W5zmtI
3ojDcp7WOelrkJl8U9LsfCJOletFHI/BcaXFIRo2TWz/JhuwOCzC8uS5iI7x8eBS
DyXBkMmQ+bqedDzuyQozJ5nuRnEDI+F3UjsSwkyLXPeKMkCaeVN8jWD2TihTQHt0
MFvK1AZkl00w/+9OaiIsBWAxobDp6dJ+OFmPz5odjXOq+v5PdQpiC7mUnd6LwlE5
a9Lzn9f4TGALzeFVwyhWgygtzocziA86KchZRHrHqTau920vlx4pQYj8NZ0GwsfF
egKlfZbnmRNlcJd4dDhB9Jx/A/bnlJKxjIfNnybCMvt4UccvZR7d499lODgQUK2z
UYBcmFU3u5tm1kfeP1s3H1OJuXeiPaw033GU34vsal6T32HApzCmerKruLZWhJh2
CVX5CRFlRvRF4KKp7DYqTIJVf6Vn1dqY76HIPwMWiXT/xEBiCEqxWclG8npkHo7m
d2PObTE5J1FTnMin7s8av0nlrOZmIDe4NJxWoFXVU1vGt0D+Oeee+pNm9NqsbLii
u1/u6+mJfS8IouzDzwsmKw+7Lzc1D0UFtpgBuS4RexuYEkn3KdFTr7jweiZvRJxt
bwvxqT1K0rFQnNSLbAkmEZJ3+P60lW8XMoozZAGhZyi8jGy4VVj6cI9CySQlUpz7
xlcqkDQehapKHBfCG5+ml60N4F/3LH9PEwRpQs9jdKhqHllZ0vvRGvRgpn+0JEwf
LDvPCiiTJz1axzKxN56FLhrHLUwIuqY5+Ko6oO9PDg5kS8NqmrC5vmsCwG88ivFP
aSDQ2B1vIIVQG+ne0lttYWSZQ5W6CnYqu6MZfB2iuk+ANMKifzW3qAnIFcaV6yZI
Y1sgVlbKLWFOgxQJXPWXeU2i7a+UAUHRbmk6ch4Vbhy2czbD4L8r3nc35jhCXLh/
JLf1L94FNOcPefb4j1mz75/RyBAH5cemkWyt4epxKKp2QD6z5seh24U6yo6d0Y1g
LY1v7fZtEDqSnJfwh0lKekemugmVnZ2uUcCretqpAA16zvzj+ekRIecTCoBawZgJ
xc8RVEilhZoGmeTwtifHAx7vw37+xIQnm+eBi67zP6bnT86fUNpPeG6CQJmuWfHo
hWqOPSYh2SHgK/y3MOadT8JRxuHa7OHXs6zgin4DkM3qdJseqxdBIrljUKp0WZjI
i6AJCqVr9qztkqy7feIlRXypAP/3RVuizQjSCTStyftsOH7/XVg4lLT+xgMtXD34
70rdRJ8u0Z0I0YKYaP8rDOPPVGK9ud7Y/G4a94ZjTnCEbIx5qrGHJVXh/aBnmMsL
3ibWrhdcwT42rcA/8VHpJX2mvTblrkfXKhSPmn4Codr7Nd0oleIXxMKV0pP/pRCm
Rrpq1TaS85X7IddNbw2ZlcubSMiHcuC0tRljHyNgjHL2y0Qk0AQ3Q8XwDPM9XYCA
JYVR9DAa34nwW30MFCt+kuIcRiXncRt5aXFcQvOzdM/CwkP/3uwLyMLoRYodSIvb
X3WkA06sIqs0sUjSasv2ja8wJYxYsCVwqSyffPCxSl3IQLof30WO8skAtoxi82WY
xsATstT2iRlDtDUtUHe/6+AlN/o+AmMsIOwX3RHqLB+1b5EBxB4sAfQjwoAEPK8M
pwSsRqS9iuWTNhaaALts9gBO4BL0Y1idevdY26AdUjd57GMNg+qurpKN1F6xzaXY
YCOJGaU8Z/+IrW6XezQjVrNdypIrMqKT+pZHJFsqzDznaUk2EWo3maar469Byd6L
zUOM2hKl43i+CmeFHo0gyRx7N3x//XkiykrPXTy5XC8WKoh3F9R1Q6oTRZ3Y5CyL
X5Ef5CVDUirpK5nw3ld553PY6Y6R189UIc5BaY42nYJp2/qLjEowBg0/zD/XMTmX
s02QqdUNuxkR1tTVyKfbl9vqgjBp9gBvxxWR+4zfYuRBTWCZOZtlPUO7mMgkGWrr
Od0oPOdJFDle8rHqQV5sujs62UpngaLQmX1hqEeQ3RW5Bgn2tm4dYmUCRi9LCAMP
j2eGRPZ5ieADzj2iyrSv7ZDdnivxWVB7ZTC81O30Vzt/HxQoyjyv75Ioz2C9+fsN
ze4U8vi1WJMVtRIcs38BbWSmd2OL90jOug7cF5O0fXawDAUiuiyv8tNjmfBYoG4A
rC+1yjUgRu+Pnvg5NB9PlRfTKr9AjfSYeYYaBkxdHb02uukFuKvccBuGxyHyBw8I
QbcdHlngOrkOT/YorqVotb07wYw8cWRxR87EO3KdmLiY9YRphoJF0m/O5ZbqFmse
aVnmrFnp5fOzKvuiM49/8iubzkFtqbyKT1Pgq9N+drtRt0Sdv0OT7rgRZ/i6GJHW
bINHOz6wJZn8/Xq8c7YtHLve50j1k2wA+7gBH3UbhkQ7ld1If8VGgzTwEhXEKwhW
943Xl77jiyNWCDhJSqtbPpRlhxV4lGKchAsPHAIGkTkHTNQHILy6SV0cZ05gkRVk
FzcW3GJOawrXV4Y81QY7NmsK+hDo2Lbhm3ZqIbht1e+CUxPXF2QUY+cu/cgA9I2P
QZYM3Onj3AXvbxvMYOQpMoxYNa0Pe+c13GnGgm/lfnbmx5nG+yKdrefWv4AviRBU
pjg2Ca8XSyDa1csT3kzEGUQDaJ8N5f0lCiD3vu8DWkyY+g2aPINKPjN+wXFFQKsH
MHWf5u5TG+689hO5quZ9QW+SzvAvRWjybMpsM2r8rJC+RJ5urHRWI09xz6ZXnYkU
AhZR/+kuqYcCnnwsYL/6//514e2e+v8xtvmGqh4urSZziJ99zGr5awMeJTPx1U4D
hcl8zdqa8pzRtFyQl83hwxPfjIf8XoNONwg5vJmBIXsoLN8qwBNBAjgsFjZma8zS
IawoyE/D6/4h3oTlNHzjOnu2pDG4VR7+tm6sv9ZqONURPolrZgNDguBnu/7oneKw
15PCoONVWL/ilDOD3ocaZ0Bkx7SNBS5vwCkHIdAbt0o5wRut5E0rzgveyHJZdZS3
UxQUehV4zWyh3vYCwbznvQUOzf1Nq5MaRgVGY4iNBSeTdJCojF+8IOYmzgZCtRjj
cpS/YEvAhwrEm6bxQ+AzFJP9LLDjfROYq8qHavFH34s0m5Ypt14klMe5PvHvgD98
Srzv+oktKBfI1VLtiNVaN6qlvRFA7v2JbkN7X7MTFfKZ/RmKnzfsySq92jHj7B/l
7X98QzKbAZKXqxymRyr/PEd8nh9ogpb/as9L8ypYQYdoHW0m9EbAMzvBI1rRFfWx
lRiSi9n6v4i7wzj34ZWjGDtnzCRXbXQD58nxqMsnnofdyLDY1UypQd6M4zJNeCnm
QcJHeEIsuGfzcshuZHVy6BhIskzb6JkuqtLKx0qbeokJiLcl48klTve++/HSrKb8
InUXJK27AatfKuShp+PZTUkFK13tKnmLligMomoenzitoGAxlE8YYDOdFC43D+SR
+vdOZgTzg1q4HQfLI2+blftCQpdKdmFXK6EYXS48ONBsRuAiscjnso/bnFYy8lHW
3987++K1iCV902jHxOWwZVMz3lWk5jKwbloBG65JBOkk5XmLZHj5RXm0YPOJjbxw
ZdbSsKOLQ1mCPDmckBfruhnbvXRE7FQNCLfS0epZqOymc3kZxL2BSfZnzyb/S1ZG
j40Sz0WIuK90e2jipKIZH94/lqAgtPTqCDQRrCSFEvoOTAvIpey3gmxQZ/EsBJDT
Vu88pHh2F5+W04kGDvNqa4zfmc55qnf8XHjek498+a1pii3Hl4UGpbYmPdDvImvJ
cabmtCi5s8/wKft2vpq7XEyZiLkHRIuiKfKFGoAuHNIOSk6dpmRiCtkTNWXF/wN0
PmFnZMwO80eaz+/SBFGflhELMCYYoQrFzIHITW0DfL/OoypiAAMHj0w6Xw2p8kOa
lASYRRqMscfSH7A+idbO/EBJx8jqeCs03mTrFPAFiJpxje8/RI/bMAUPhoU3EbyP
0YFF84ikqs+zhy1enJXYy4NHoWHI37SYsIylpbBaAaJj1fXuuFUBkxvRRHCMNNyZ
gWnblhaQBxJHDfRGspiImn87zX56eQVHlPYP+Jf4XG1aajVyDWPXaaG51OhXXV3A
9S0MXZKYKa4sO51PuSJrGmPX18R6YqbCoEyimgJGPMzi9Vwyj18lgK+cMhA5ZFkJ
9euGL2Aytq7Zcf57j2EUudV+v2CZACiRnLCs38JByXIbkIrv2TugKr+i4KiPCmlz
JMxoqlmF+zmWV1pRPpn3mgKZByJ+xodKT8FXdl+HVEQ/ueaYc6ReG+HoUKUloQWm
88BsuB+lfOyT8jjBxSxD9ZQPiECnSb7BwitU3jP11XB6qx1Jh5GzSFkVRaazfoqx
6LCNxIW4L1Db1og5sM8FBYunu0vuS7PshoL29UPblHG5yg/ugkhnbP9dA7ZEESqk
e1Zqt2H6RhH7wpoq3uB19mGh53pnTXj7/hGEdaLzxJpfYDa5uP5/5UmlXiotoiKt
TVTqg79M1UvV4Nhc/faUB0kzjuXpQc1owrETNE3QiTUjm2zwvkGoAF/PV1t4jOyP
i0esNvuTLe0gyaLsLeNx1v4HNHKXcSnqftAti+Fum6XPfUBm2FGfxwTNosc3dcOA
EqfrMKtmYFIt+nLp5HQbkGXvNvAuxXNea1AvEBPX6MOe4zziKu0QfAsyxAS+Pzkc
sQ/icRlNW5BjBZr2Kp1PGfiA8/7jtwn9SeVk4AiW8vDepOt0eIS6LW0RbjLLWE4C
BN2QEGqcmdAWpU69CQ7NhuV98P3Kwgwrv1Xzqa0IukDq+MWkVH9pOsyCOxxKKQuq
JdNh4UMDC3k1LI82jQiegs3Lo5qUGMq5jNxShaABwW9l18bXRelOiW7XBpYLi/kP
LHu8fRdi6PXFUsA5MUil7D3Ogz5GsQcIY7S6aMvrMUghaATflqaAhcx6d04VpXU6
fjzZt5+64dk5SIWit5j1FuXTk23R3tFmIpP3JW/ofopYpxGFFTE/o6AOn5TTQ5IL
NvjiOxL5xHaKsvYUdPwc3oMUZs08luiu5S4PskAFhSQ6lVykLSpITbJ6xpJUSrSk
6d2aLAUa3ckRhFJPwpg3BrWd9hvtpJ4DjCUNGNxxSc9uUMKUBteB7bfB/iSYaHbV
s6rLm8tqxTogYt279lTqWqYojUhuDTE1FJo8ual2wS1so3e9FzjUjAGUwILaW59s
WUAHx8xqY3UcndJhXzjFj5xZ7e9WBHLWisIqRUB78TObgn3qfrFAtHZeAwFpdKGH
6uumZiHntv+1Q3ZqDEm+JGI8rTlZIGqAT+AYKxWGYFi2nwIzasq+yclQJnu9Fokd
mtL+JaBWK7A85fg8PKjWV5uVOyq032+Ezt0rRsXWFyFVlJvobCR5UAL8N6iSHTyx
IiFF0kFMjfwT2HOsJevENMEeaFyQ0snhQrIfuf2SqqwdXpKu82D8YiAz2CtqNfO9
JIMJGoWru8i5lb2ur6g7bLvHWDaH+odwjV1fYBX5z17lThodjfcoJpm2HJpUW6Ix
8pJ/pSQwrj6gm7iRWqojuX4zR5pOjOiICAX2YR+g3Pf76OegvX7LRWVMKOTzi1Im
TOFm+NxX0nHA8GKQFFQdx6st9O8t63xbqP+CUS0/CMiNvOrO6eKdMnGjfGJcEqoa
7JW3dodPMOUO0dWbknGb3TjjqoZkOHp1bDlC0PEfeNDAYhh8uMbS4hZWxgUHthFs
uvpf/V3Xl7tN6iqn6ReiIEzPLXJJXeA3BegrUcSm1l8f+rHadif7oL/CDMvGUxqD
zi4wWyKysalxcQX/PG0UT75KlrpSEbJ5KiQxcAXZt3amWPDUQ0yosfqSk/BojMdX
Yw9OqkpQfM11KBSz8M+CInDPuZANu4bevtm1N8wnUlsBIHWuC4189nTdH5cc5ycr
WUCQHpE/bJNp2vC/U/4c4a7QppghrNyzwkny9Ns9urcVTbDyoBYFmRiIvOhN05S3
1yI3MvNxg003gfUCO/RvuxDfuHG2lcn3FC60vvZvDP45RMGM1XmVB2Mz/2NJaTva
6+2mL54+h7Uyk5LjGe8pFdAMON92+89xFrDDkPNJtkvKBX4QyH6wrRD+WvblsiaQ
vp3iN+8tU5m3daAk0q+Py5oBn5YdjkeQHv0pfiPbGKs6TKp7nAomVfP6U+hztaXx
yTlPOU+rfIL9WVHAaZnm4rtHt2D9jbp//qnIqES2nfZS91RrL0FLwLQyooPbsYZU
QprQL52hR8b09mBdpNbRWF1rTbLd+AnzvbHj4irCpFCNTXIOH4d2U+dDjJeq3gDa
6QeWuabHiXnB5f37EvwhmqlUlKDTK7ueNyc1PcmZ1L8s1Vu3a9+60awcyaPZVJJt
EdDKKXAPdZkk8rs3nwyKm2IqpZZmTvsYIhTMX+BJKVHE7hXklwPhbN1ToPpVrVlz
JbbbuzSTxFAgN+q5R/iqjgLxxTkmyzA76AsFNemNBGTED1CVkJD5iDTaGX7WgL/8
GMHuELY9LhYe1iu2zb7RK94BSPQa0j92U3kd3s3HSRemAw7He0ew1Ncz1lPUtbi6
Ys3HRY31l2MUL9BJdDJ/o3qEb4flzrEiLpHOQPDzQCkkf1/z8j4XQ9Wiy2/GtvYV
+KZZpMk4wblaUVaQ9xP0xTcf5+DpGtnKpZqSfS6sFEOk7liNEAyTd0d6QmOIu/N4
uqZIWa7RwNfwqziHcnVMKGEhEhlH+fjfGlI+faIu3mPFzwqutaYLD+JAT4noamK9
Au6wx6+NPgn6JdxGd7DTAYuhyiI338aCSv8PU7F5vplAzUrgmQbAcMQIClaV5G3d
fJLGdFhnylbuxqhLkzhwhQNcbdAhN6ufQr1IIoN4s0/dxaBuT5kmbEmtokux+E45
9nN5zQf0Gwel6QlAux1AbfcDrpGh7md1Xz/2afFoji61Y8q0LtkqlMkKrf9Qx29Y
021C2NEmQl8PeTXErS6Fk8565/wtC+8Wx7Z4xmSHos3TwwuBXWi/vHhlxs7PxYOc
7T4uiJUT8b8Qcp/4nS1dTkjMcQYdYTyKEkAOmZBfxlNLxvpCaB+Ceg2h3ZDWfYwj
B4yZ+mj/mLVylbVhzcnLQ0vyLYcgittqr5eYMB1hd7bRcdzygzGXO94abxvejbEB
rIOsm12tjsICHUxRKv1dVi5V/FX2MGTFpzgK5Fh1d2hJV49BjoFxKsP0Le2NzaIu
I6ZalKlPLkRr5SqmElWjeiwa6pRagQ9kC36i2rOK9eJMk7u9Ar5vbgVeU110qMwq
KtAa6v89TnMBpKuHnEcbe2pkrNK+3194b7MHJJVq/NOGwpv2AvsrJSfjLp3Xp6+P
1421YkEtHLvA/zth6xDivfDwPSm1+gniYQZZZ3CtwbjnnO3XBPnG5bOvAoMDtUVQ
54omGgFau8JzpT4sYfxaRr1ZgWeTRuc57HuxaVM8A70b2Ad96yVJc4X4WOa7ISfr
fCYKzbstal5vcJqZMsi9cgWbWLMBSNgO6Ucmb4eSX+kRYVn6KrnVarcjeahkfaD6
DbXNnNCDn8Lfe8Vewdlb9AdHMqPpFhKq7FEhblB4Y/2F9ngxR5MRksxGiAWHhH0O
A9jGJAfme2ccjA2LNlhIUZ4z58VkIdfPn/vdqohA1jbAD/USwF1LO/g/Ink1qtAn
BvrUmNB9rzoDZijSYssBaDWlDwczdZg5dRhiBBnGOTvFnmJ6Lug0bvxNGMOjinRH
PlRNg90NKyEJ5eXo3FajXoLO0KD76eRvnLOoJjlPH5RXGTyEufc6PkCgDywHeGix
3e92y/hlyC5gLKyTCXVm8d4Heoz113BJvzMKyImSDo3CljeaMS956wDd7bhozu5l
AUQm38QmxHSZ8vfwPVpyH0WJ9Owjh2vyhWDfcnErxcYLJ15MmSaYEd+dn61AZFmU
QH+Xr3PrONeiatguKRWKHFTRldCQm9QZnZpqJMGF2uQy91Zr0gJ+oxjtCxoVA5Uv
pVIICthYtaGX9cpG6sM7b7qDy6nVOoBIFGuaSa4KMundmwnTvRmEbCt289OmJQXS
J05TjtNrJw86WWXvsbAdtdtoM7e2zHt+a6arv+PdSAqysqLKxxgTas7AgRQfRwoG
3PZyUD+3nyshMeBky/jVGLcW9e+YaNAwrKNZhny4jL8EmdYQEqD8mzaOUN6Qn8hM
W/KsQCGbI/vPqoF4ECqLVTktHnfVN0kDF3Xd6vSPCm2Kg0wWOTrlYqqAAUqtvNRj
zKxJs9PnpDelZSf/p2Ho+EnIiZPYVNiectnZe8h0lgYZjyKZXju1iXH4kwzJ08ew
/t13AZ2RPOFYF5RHpP6mbQEmg/cNY3y4XKVFxOGSUF6UCuXoHk3PhldBLgbU3r6/
rKi7XSgGmTEqnWguUNRUJmxFGUMYjBvmM0Y6FeNgm9cJv1H2PGvKxcZdthAUm649
O36yFzKpgwWf95z5cDz/3TbtxRijnu3cdS4nYueNmyFH9xbpI/vJeYjHYwObkf7u
wfusEx+k7tHVvFe+eItY2nzg29JNTo34uX97esC8CRuiz+WY9z9Fzmh3f6rBICKn
J/TMyKaZISuhtiwrY+1fXmi2mf38Dw+qvfGimGJeZmIovfGtLuel1Yade/sriw7C
uzHIw9U+/oJi6MlOD9b6xkz0jRAN93cfwsTBG4r0Opvyn0x5vJqJ5X/mUXlTyqed
yES0zkuywqCoukM7Me9RWm2B31ZhFf59eI+YhfmgaixS33Ewhphc6E22rBKwyzra
SX57QH6ejqY7WKim4r5nhYwFV3fkaQQrWDJ4aohSN/3VmMMcFfAUL72XOc6/7V8H
BPsGzUcHTPkgjekt4apZDjx32SjPMR9jvJJgs7QtvFzyb541SI+CbGC5v2Ok3Htb
b/AxnE5mNGgZl3nfbOBzUjvwvxGoZGyRLnors0+yxO9eupbUKa41pRHCN4qhfpJM
y7cIpm6o+6SQ1tx+uYkO0Ddj3OF8nCyIC0Iz4asdFuISHTo5YiueSjVWFKkm9ccO
Z5SiBhLtcS+9WbUu46gc/I+5l4ojtD49sJPnrXDrRfhVvGfTJFP4Pfi5FyG4TiYo
1CT/C16T53xHKeSkV6P6P2pX2YDQbOxOhgyG0TWXWtMYrm1SD6GF7Fzk6ryaJ/4+
iAyDTjFgU4rhw7i6mUx/ibbqo3ivl+srna72leVx4YVoIjGOu4i8TtgtAYJf9PcR
RCT0HEHr/it0mlURiWJ7u4E11ZwNwpD5xzSUSo47JXBBzV9UkDK7Ixfgdn8tMCtK
7L3o+twyi1DyBkWe7SuFcMcNRh/uTiNhqF1xmSA4t3UtZCUbFIOrYVJ+HNUGQPdF
Oah0GvepzKL7y7ZGygLrhqaKPGtsud/VV0xhHr1k8lmXRQiuS6opwjBpQL5ZbKa7
uNnX974Rea/KRgB0es7grhVOPJJW6M2Dxe7fiDaTmF14+y9C+o27HRDB+5a4mgAg
MxuCSnfdApNGltEwbKxjwlBRwFEiV/GVKuvHJqRH1UlECvVJvTxK3oVuYtSqoulp
erqXDI8Vy0oiU2leTnKQc9uqDhfB20IaHRzVuX9jr+a3dd51+A0TtXEGoGMndoT0
Zm4v4H2I/i6uXLc/KNO2PvEDXYzQvhNeC8N3ABbrrolaPDwtbDHa1KEbSNfWhU60
WJj1+A4wRXpnIac12z4zVnvBPfp9bXz1yei10a/Qx3OVOQp7bXYM4R5wciW1/Y/j
oWeKqg+1JtI+B/+Bji+HtnE8or+9PoTchkXSwUyPxx1oPzmmmoD9IACAQzEd17Ok
rEgZKvj672GWK6F27sdNsE76plDW+NHcii08YCd1lWbBhm79Il+YZAFlXegSK0q2
LUnagBOKNpgZHvU/QqxdoFx8ySaBrSGTUMKo0DFsElb4xM65vR2FfbslcUmt8van
bu6rXqeG6dpZHTukfqLYBst3Gja9YvrzsYW147mA02YtfLCx5R9Dqjw6BWEMHD1z
uT2P7yC3/HsvfI3MF5/0GcoM8M/gUPIeliKhZCSpIiR6bVscIjeyzi2aycuozRoK
/bADVduRvsOgpB5VEEp9Aop2XNKE3o63zYHUlnfTrwMeaGuaQE4bxXTrkjfycE22
3rUZIF3e0e3qNz3HRHSGEEE3s5wg74l+rhi6NxcwdMNq05lhxdX+fpOAztMNOtXq
OHxWhVIw2o6PSvahxRpO+Hdp3+EnArjqZvM8a3HbrK4+PYUF2Dl6bGZ7lAUT5vJK
xlfN+Ob6EihlVBAvhT/rFUuc+7R0x/OEFZ3pnqXxW0eO7naimcwHN23c8smwri5X
DIgx8yhRwoDtQ+DJbQIlOR8j6tzG42sf7c4uR++3D6EyoxSQ10r+pykwLvuuFqC7
2jofLCDHJ1txhKqB68DwKl8Sbit3OB6X8GW5FK83SovjNYRsIzLJrBfghT9m0r0U
nmkQqb6vc8ita9gvj+7GDiReIRyKLsslDKrDob0gHxmn/+qAer6TIJyBKTN/ugAc
JEX72v96Vk8FiG22l4QsDwyTcodEebYDka1aqVa4dCtcYaUYNK9Cavu9WZdwB7n+
lRt/lZX+0tDJ4Zt9vQCXNcaNx99T+62BiMvXuRMWfQZa5Ou5QlaJKNzYmiOgyyqf
7eFqXk755+y1vtlWB/YDfZE4TUdbONkE6LeyjgPq8rkTeeIHEyjDWc3T18GHzYEa
r0huifcFJwiXd10Ef84gYkoGZcOYkbRtJhWCTKcKNvb1p/qa0GWdc/D38H7MqLx3
a2RQNs8RYzlCn2EkTOMmxrOZeZds8oq/1kKhJXj/YxbWKsjtakR0gB6QCPppryeP
c48dsyT44G+06GlsmvF5eYgTteqc2XVLcNd4LttnOSek1DHc1sCVNGOR5TejDJ74
dgHcriJ4j4gfljIJE2GSUc0adcd71SlJM0T+6HGNkTV5lWThA2TYvG1rL6Azx7Cp
I4tdBd3QMb+R7KCiU4P5KxNPO8xmLclS/+WvULGbhkXser3/hlqP2GE+O7AZ5MAF
IBRZEUEae0F9uviD639EyfarUqr8O1nQirBMpiXPHtPQryEI07X1HrvyprzUcruQ
N08efphqB+tXmOqlsiRAQEphH5uJ9AWYR/k7cGfkv3TWsCCsWakQjC4Go1FmgZ7e
Q15OC0oeC9KC3YgmNQWbfR7mJXw9rS/3hozU5n/m2xjZ1CzrTikhOMCqdqz79gZ8
7Ufy644qNHf6VeZLHttzdj0F4n9GxHWBHAi1q0YC8A2GBOKTVtfOZ7hpObisZA8D
bIVC8FtBEzy5Wi6UVtRLJkUj/+GI7HOKFHI5DIGEAbN/eYZpeB+LSQEyK+TvX5W8
NWc9iA/5MviONR5TIeg6yd2cj/IwiP2PL8Fp5mZJi5frbSkU41Ip4Ak3THNPTMKv
z031U1Uxxd5fD4SGcamVSHKDgq+jWLiLNq0/9f+JVKQejB60vdjenNgJqIswOEv9
Bf5PDANT6OnQo7oKPUFeSEXAyCY3Tr0eGkxIKc2q6pbpO89QpMNPbxBAo1R10wot
AqZV3d4B9uQ/3dNFaunzcdUr4s/7Zwx4FBp5EdJ7ORAcSl3cdfSE77fGgk981K4j
C62lS5fYAvd3CeVPkpiFl3H90tu/j1LkACEE9dps3GNhBsklvaDSBmGjMIEuZDgv
AujzOwrVtc+m5C2m2WaoeYhMAFU5I97ek9LFBWBeJUmzIkAs72s7beBhw/NJpKxE
M6Md1/ro5Tb2fvTqgNw7tosTCpTiZFBkKeeQt6yZaoW/XfZcwCZXRSnHZ//yEfqF
fgk/9UC9nbt+m4mvOzFeyM6sF/crWCsvilJ2nlB24xvQGGelj7TPxH6wG4XRFTai
7wv7ZAb7DEzw4xKlpz8w980wPlJ3TXIFApImiyumcpbCqfJBcLxGbusj7sR80RE8
gmpDwy4838v8H4YlM+OsMw0qWbGOvq5p0CSELSEPxkAXsW8BZFf6xwBi5Dl4C9Wr
lPs6pxKR1iUbgZQ6w7OEQWsxEKgSTNyIOyODrJZ7B5R0wmooERXRrz3CmwncTOZf
45I0l6tY59NK9sW3L+ODZiFrrR6bAP/JmOMZttxuQ0p0hskGEK+E38ILPn0oRXwD
JWipDN2HHm6ZOCnmqfFvwUaIOjGxJxpPr2ia6PNEOuKmYsgsJ8t3+VKjm/aIYsAk
M1NnhR+1iMOv4+s1aFFMolHac1qFSdrRUw/EzqHiVWoHBz8iAuLwA69N2S1NctN4
s8VbA7wDqTj6wNgQDzt4DBzWJaqvx9AnkcbYgOKim3k1aRdNoSWc7ssf1VPXDGr2
nisJSjE3G+WFgOaywW01fGovzSV5/A3ORqhM17AH95hmJBk6kMMz5Hf4mrWJ8TKf
pOwZE1Jz4QZcNP5R4km1sDvXyQqsBuqhxwuHt/6SbFE0DSpHwPYT8X/ZjiRh1834
Wq/HXvCPVrZXtaizcgfydRir2nARzDJZji7LV1eTsDUd/QGld/JJWhNvl9SFMsvm
D03USPglgRj3A7kbH5AYuDK8u0cVuqlIbadxO8QAfuvL8I/Ra4JyPzl3w4SGxzvw
8tlb9nsm1/t3fts5tw5UllSTPdKVCI4our7I3HIQsB07M1dE9/I7l2icJIGpLK9e
sZK0J9BVL1/xK7qrvg5gU09srQog6j8WBYF/g6DwOsDbqUT9eAYczUoSJeCVA9tD
TX2w6wuu8taNmGrCOIKcMYmsgSBU8pTzIgm5wNUoEJHpabvBhnbgUn9KiD9aHdH7
W9bQ78aDW3vWhzzVii6UJbYdrTPYPBtdmNEVa+ULUAqNMDAMWK54rOb+HeykOoBq
oLVmSFBb43MxuMdP2rzqqpU8+pTMNOc7XHcCfYsIua3W/sRycQL97OQ+Zwgy+lVr
FEaEY7B0d3QcLS9YYyhfeoo4D/TezwG/FUcJVMpoNBIi+1LAJztABhIuWqxQ8N6f
iSB/+WYoijvc0duarTRAKkegVLqn5PkZvcjpivoi0o26HhtRs6Lya6Fd5Mrvd/Qn
Y7rd4oawByvSOYru2o/66RrsqyLj2gB6AxcdKKR8qvpO3QLj4J5UwuV+3r+Wf7bz
shWaWVGJKEZQIp+f0k6Hl2OGXdlHxPVtDLbseQ/J/56Sq6PGaxNQyaxg18MP+Xqn
U33Arm4xbspZPg1f3k/IZNyxEb0sewKV8q0VDGNwNyeMZEnv/ad7hYaDbP8VNwiC
8SwWFz+pTS0QHcPkdmZuxMUMPKOweS0eGEcvkF36xq9KIZxSnRwEEDJ/KVDIdYCm
v1ugv/G0xmNYQx4ZrG8jq0Jv2kKEhQfEwHMKZRCH3u6hUvYzd+JYw/gSCj44vnTG
TNKqD2YL+MJYDNdUJFSSngyX3khS8/3wE1NOX0oD3b5gdwz9hu/jY5JMxNR1JZcA
C7GVlGyG2zKhGnuWsvKuZ5qnEfVcbVVLcYFpin1RwyDFcDpp42SzYbRfNngRcEBf
T72/fjEbAGo5ECZURT5ep4uz6TfPafdRQORg6tgdjfUg/KtwtCwEY8RMKG/qp1yf
L9LJYTz9cKw7sYrf5dHvinkwqCiUcv8Y+B+G7Ox6ojvwtWPXXr/NVwZmzucuKuRt
CeO+0xqGO81ceuJIsA7Mi+Pgguvi+rZxgF5GyDkT9QuiR3aV6MiKkF2QPmQu4ZsM
2s+NgJN2xTDREIj2zewrTDj+V8gFf0FF57BUS2oBalEs6S3174YNfruodZnvEwr0
wu0sMln19/ewKFhuG7ZjWeNO3uwT9/8j1U6F7RgVD/UhKEtrKUIhwY45auF6XxuV
R3HeUm/8cT+2tcqswmYSnMYnS2KjgMxN/1ZsLZxu7c8SDUi6Up+v4HACNCDt876F
bhrrTGOtlUJo9edumFRaXT/2xaLDa/aNkAy+SuLpH21q6MKtKYCiJNz5B3Ytw44a
5Vs6/qCY8uZmqMigRsAHUM8AMci1R5cb3cZIfpK5isw5tzJoOAFGFr3D4BeA2nMV
DQgjN1yw/ZTJeFb1SXCnwe2Gh7xrMNR0+yp7SOW8n8pcqL/ymtd1KIremZDPQiIP
tFE3D9lEJ2gJaOEBg4nyTqqvEQdQhUSSPcD8l8iQ2ySagJz2xOvoJKaAFIPbjG3f
lPdrAtTLtFQubIvQMmxqQyDQKn7kBfoku3lVQaC1+e7s1pmzGpePMnsYYEOkaPOT
fCcVyUyuv7lFVJ/N+Y0S5GD0vcbp3sg/u68wzW0CHQcOldmc+4j3jSrClGgJ2F1B
X70vO597YLycV3iNaz+JA8IXyWnEWLWS2TLPE9A3UcKNSAxK9HNjSB0kEg3YIkoD
k9TZXUXFZM8fepYE7vZPcSHExE5C0gMjrr1zAWlgnc3TJvCzykOIH6ScVhrJe2Bn
pgpYY5g7S5+eLTAW6Pw4FtTXfgPYs1Ewe38YMv55shgJLV+2PTeEurMe66Xz1ztJ
EbB03IutCGCWxR0uBbj+44wa9eiYj09Y+USKuHrlWY+nUTmmV1f29wxx2JL5x4vc
TI7jTte5ccXR8o9kb7gkDFOG/7omNjotQ8UJ5kUWfMYSKs09ZBPJ6AN60ZrEbY/k
cdha3WOk75+KbmOqC+lpfx0fBIzE4stn1hrQ2ypVdfArGPk0/ophrWc3jtlnn0n1
314JH0FgulKabiVisDWvdGRjAfZUq+D3swbm/7UBOZAeX4HCHCZz8UUWi2Ru4Kk6
eCZ1Mc62WJIjm+3SIpIHTM3ht5+t9zI+4YGQVqe/eqKphbMNDlMneYqvFe+iYnAo
4SmhoGERq0yIwTIs/dHEmH4fT5xTwKUW/KwID4UOzCGlN3q8x2lG74l+yLhuQL5X
4BL3JQJyZ4R1H5kvfBdEc8xkBKIdqnjdNoxd9KBkbXe9aFHvCNWXorXiUBxZy7xb
l6lmwH1fZO+wOT8G4E6kL7WTzf+50jcuefMqxLPpgsRUF5bgF55AHhODclypcpA1
v/Y9OFmyyjVlCzmhghaURTc4plclHDcs/caTAVeU/+ubwekvTV9WcYyZUCXdEh4C
kCogIDFOio/mFoFXP7gaTDEw/cki4F/7bTSLaKlyr8dCr9fkJYS1oCbPL7eTHoDY
1TmxYzZJPnB8QGFTNQvPDY3N/3wokIec/f0aT3gvQQiJYAgzCmmrUkKZZ+wSJrlx
jq+2hp8Iv2ad9fKa++FVSxORTzDH1bEjgn42iLc+2Wc0hWpCZe7uXJeHpoT9pkb8
E81MRsGeNCn4Poxftb2kkArG+kFz3+l5oXJdshcH9jAIWEH3ph/v5fNjyRUsysRG
4bG/vd+/fgeNix9VQ+5ykCA/Wkod2M0MUg96QS9jJ7dehBc867vxfDuAkE9qN5zi
wp/eFER9iPxbAZctJd1FFyO8pzqJngm91QAYnE15cLqIzjTZ21/vqFRoKSZG1dlT
YcKKiGM/gpdd5YagIExf2ZJEjDhgnmKsT5nJ9H3HGXk23l6vmEBr2jHop2gYSo9Z
gKA70/V4rpYMbrDvC3QLcsSvgZ2LtgJ3KM0zEke7FHOJ51hdlDuBatz62cto+IRh
ruOhlf2D3xLhSfODsFIyjoSG/W+Rq/8SJlKFE0lt1yRs/WUKCmQQq2UxsO/waCCQ
1QLRUDXxROhryXB+rtzrvYJvQPIUadq/rIRO3jDG4UImhbs9+CiUnUF9FLjrw7zE
565My1WdBKnKlQHssp0JTL2PUOX3fatAUaUIiKynm0NrUKTUGZr/Q/KptgPq1ipG
3FKyx3kobZbgOM+kSOyjXM7Sgh85W6vrBKI5xKMnp9OGIq7XWKqCgmmY0gpoMD6Q
7ohvMOgfNqZDHXc7hjVxzzx43ZyXKjno2e6JJHlk3x1vpeSy/Um5xCwJvyB87H9a
5zzfqbrTJpQkpwE9MBiU8oRGT0UzaOJpqm/O48ckpbxHSdf+22cCR+wzsw1mqToS
Sne4Ba+ZbCvas4oYg7L4IV0HujdYg4KrG7ggNHGQSAoQWnvOIGFG9+YPv9l8DYA+
/cBOf2FWS351pmTFAMBelRxg3HI+PMLJDZHsz685UNsCDrW75JdNQnvNjUURbqSg
XPEgl/XqxfBY6LaHdha1KRjW1wtKw6rUDjJYmD3tNFRSNUYu9lvjkNoGPPwScnOk
Uc9O3CbcscfehL+ouZ8RbQUyc4StUTYOMXmk09usfXL4zl3JH3OAq1U5dxjxfujH
tTJd+FtElSNFU8voou/+gqq82We/epRRLGD7g8/NISf9vW2upJqYSs4ijDLHpa8U
0RlHLKfRrLG0m+OXyVPy2wcQUOoCSa1Ujxb1bqvvDj631hz2IWe/eTfusO8eLoBA
e9kON6yw7ZRr4btMlA+Itt4sCPVRg+6I17blWVZEyC1sMpgKlA3GkpbYe63/rdeN
uTmLfRgTZG5sygWQsVS565Ie3+komN/ntoa3Vw7sGhTrndyXCkygWnzVxBgHFq28
nqNekcVa/IIR8IOBQYT8ko6Revtg1k8sjmLQVAcKlYb/+4os/G8uO0IGhjk/NJJF
bSpV4q77TARgJT2nBwiTB9aO5DTYqeLAchTA7jiUt9oo0OZxPtNs/PoKzSTWYEJx
cfmDYxezGQpAKj9DTOvwuBK8R2sBHebEvENNW66J8VaHYAcqfxNJ9gFAoOBFRckQ
Wi5Wbs0Gx3WJHzXT0RxqxCNCx8BCLRPKf9qkZgg+rhJHuFoOuwWxSnv0g25nQltb
2mWXbarX1//1HgUFxZB6CVF6iB4tiEVOlM+9aIGtLX4e3aDySR81++YuHRhepCwK
RgELRwfd0nzD59U6mri4NeSlSA0NLvtN59dX6nAEzh5c70NDdWx+7cgtDin5e39z
MnmgTuaB+wUTRNwAl0O/6zXxE543v9XLPftCW4US5gdvDd4QQVWGHbCD6ynb7MFV
7gnMqJ3HCWr+B/v1g0FH0ttkZrUaaI1x0fWl7E//WHlVY89QYpfCqd4W1xXU7OX1
0RtoT1wAtSZB4Hxr81M3OtfB/3IXjKfMsOJMmgcL5nyxvbBd1oxNRsizDa/GCbnG
bEaFK5HVNbre72EccgormVcWisFNFyxg+OQNxzpf0WUfpsc66r5CBr1P82/W5DIf
/DceOl/cAgxnmoByAq6XXdBbCawBgD7Vkp+Xwo2tFrCW7FDd0VjKZfRisb9qUpWL
fSx+LA3Zr1hNGkZLATgL9Ks75ZNW9aZTyRKWp7FBEN0NbY5z72HXDkoqsYMMwaEh
oH4Dj2L+BYxz5AfXP+LZ7/Egph1n4SyAci57SSpTuknjQ+iKdvk8vo9DV94TGFjl
88hcuSoSljxP+swCExHEwMk4eUnszi3vdCEP/BFFxD5VQcm+W7V4jGaRNEqdbMhi
NRLt2dibcBzrBOHDVGo5n6ECFidRQOtd7HO53J1lTpt2G1ICzQO6hxyKrFDx49Av
G4/plaE5dJnQk3NJDJ6GuZvyAPkTIRFyFNIwRQ3/nNlCv/2vqbOWuD5vc77IDwbc
YR8lkjRDYMAXzaPjVK5g1j/4BKVjTtGtHZs8GbZbzflgROiGvYwJQoBFSYBod3Sq
jaPZcweHbphUVidpO9Ugc08Bfz6jKmsGgCLretYj1y8w802HgSU5A8AldmKLQ9Dk
y2OsB+pQ0zwg2Sk/tSH+2a8y+3kXwECPA7Gz86tVLizlI4sGLWuCFuvJnMXNCKid
mekNS+H+hU3pwFvXYs3oA8Jz4lFPvSE/8ZbmQAjSkLCTqip53GlxWJ8gYSdf68NK
awcffXpWVzcLTffUbi1CLg7o53aMUkFxVUU5P6jj8hWhNEbl5idOvyi/iPBmQKBN
NmNvPnWIFJWjX++p4/v44vIHOKLLYHrx3mefeM6RlVMG0a4rxaij5uA5XizupxfI
vHaJi6kgtdAFeqxuW6yS/rUm+97kD1GAd/guJ7REr6Rh/WSLXSvBSPJPIdTWkqMz
jMmgpVt3Phmt5/2R4aMtrS7byEarqppxmfXWSZJEbLOifgU5vtaVreyX4fgPMTho
tWeQ7VV9S6VcKTN5OzVAEiIwnULwNdwobH+i6JwkxRH0rVr26ZbZLwUQ0ewRQa4f
rVWy1lSw2SYbNX1XPS9BNumJzCykPIYYh542F0yoChD/7V9MJk4nemYMhkirjC+D
MehVT6+UFDfEZ+1xT+MuWHLEjFe2tBOiOpgrUsoja1xONVoOvXxpCafOCM9IN52q
k9h7udb8UXZdnumoEczVMcwNY4igyUe2HkkAtKE8g1mZ48yuIeCbHYAMb1LbAl96
mvCoEiyrgjFTNsgZ8QmHm6YPWHXPwAQ4/z6xn+gqqP24QBA8pi6qv/5i4VDygxX6
anoRoWO7IuLDiO4+dfdnsGmo5DywrNu/vhzSkvHrsVW/jvPsRbUZrRPO9Vvojb98
al5voewVetd8MKlSnrqMQOFWRqWZCvFIlRUPxPf8zC/KmNp1sD+FB3Eanh2h5xUz
rHvY8e2og0QvehiD+byn6oLVKLKK7xeWxVLCMsLjhJzK+pLMgI+1HFnPywHGIMvP
KziJiO6+gRxtwPGt2KOIVf6L5ykvkHNmzjk98aSQOqva5KNgd06vhN7ExxbKWhEQ
dbzX0rNtOeELx+eDfhx7h8S+1jrMKzaf0ZjoHJm4Og491bEh++G80RSinUkmNgqF
c5VrnKH2aKXiwOkbLCtJ6X0N+bPzpjIU1bMVVqeEZA3wn+bX3MLTEHojNamrMSxY
3sTfUO068U8TvD2z+ez3F6NJdxmeF8kxs88zOxxt7pIQ9hSF1vW7K4vC37djvIqq
6Rig3rg4i5DYr5y0jlswP0OZtS3x2PNGD5dCEVOh8UlJ2UNNG5Ob9EJg7tPTMlyw
N+qa/uVe8hIabQONfvr0QKwkn8KWZsp6ORdPC1TaQakY4/lS1PVw/G9C5N2cqAzc
PgY9FsW8rCw/Th5GVy6T5H7xHvDjePaKyZWUA/O08Ut8aOm1whU1g34x+RcOqsxl
M+QcICMx4ElIlbNYxCaGWjI7L6OsBwDHvJ5wOz+cF1NZsh/iXYWzPiASH0hLf03S
YtQkyUEMaLklXg19NOi2+TksKlGzHx7AKl+xxOEI0Hl3yyLo9Hc33Tb/Iovi9oDQ
igAKnL29WYpZFoGWQKMabx+x9p00yBr6YIfR2JisYgqay1jV9zmlZc5CT4SPEouE
BAvxogsJ3t4ufJE2UTPcshYnwGLQ3tKU7O7ndriOAbUDqH0EeUpDEbua4mLZlwGO
kbp9QbKRLYWVr0shWQA3OGi+Dm9eo8k2W3X7kw9j1P8foWqpjHMgdTp8DzQopI/d
tzQUyxzOYF+GmQp3LLUyTTHEKrLXNbjqDdTvnV5KNxlfeiYOnxe81i8IrKmqYgve
x9VgDlYwZyRtoXK75+ZwpDF4OuA+HCSYo1SYx7a1FdX6yMmxUOGpTCtalRf7JTEE
zGd+/h1DE5ftXJM32Ir51SYMHo33fPBoNERvG+eQngt0GQrmsWt/sQH3tn49LwTx
d5nyTrMx2C/JPM34LDGQt2dxd0M6zMyGTQmUinf6pjlrg1ec+DGd8uHp0iG9RR4v
fK+8vQ0/TxMmQfqZDGm2YmFiYy7q9sd9mcBBZEj0U2YSTuZ0Uo9F4L4NNAgx9sNy
Z3Li/ji7kil0ndPpfNS6cce99QX2exkn09+hTFKdEvEr5j1Pklgzs+e33VZatykw
DaeGs/3DMaYWdoSXxyISl5jZGRchung0EpAhaMGZgzjOhxUchkV9s67IiVfkxXYI
bVn6hEslzxGaL1Cll/DJoG0+Vk9lIrmN/3ISsxf1jnszPp1wsc/kzd2UPSFcpzyX
knTwY29VdvP6/M0bEujiH+Xe6souE/mErXQ7+2L/SiCQ2CYhS0jZhYnoT+uwb5MU
7Pc8lV4qVeYLqQbzrbP9nXsuII+oiXTb9euoJNyNd+BQPDBEaNNBstilsjYrbn/8
3U4dlVQaK09AKBi+OhmHJg63d+vt2swfqfN5NgxOtMGRrlBkJTjFhkMfys0/PiCn
1Gb7BQB3iNNZ5nnchpOwjQHoPeJqL4vkYytfHb92dZr6xqOVk7jR3NHJLTNq+OUb
nRBcFvM98zRwgIDDvPxW1rD5E1T3+nDpb68g2eVD5GFn6czeARS6ieD8EhtWTEb4
ZhWqXldhf0cT0QkYsieIGqvys1Iwi+ruFZZz8qnoZ/X1josuh1w9uDVJi4zsdqEl
DiYcU3pVClfxtsOLvXffweulvX855ZAjrq1DI8ZJGapqfmKyhrvNWxPbJGrInk+h
sULTqHQXDppSRkUmw2g5NRfwB0pOHsJq+KyJ+YcgqVcz7b7EcDyI6yR4JeRPADuf
Sa6yNt1FVOpjKYg3mvKUwZQ+WzIjiKOsD2zKJguMNJVe6BgcS34h7ktgotlCciBF
DriqxLjYpKCv8EWbyE7DbL4wc8qzlnp6ridKbZpuaEihhbimgK/p3q4hFSP2s4wO
AB3Tt/XdGHDq0FU0yiPGZEBmDgrffzWkelxrrB0fPK6gPqJ9Fz8oWflcw/LC/qMw
H656cBHm12NQ2ftRMrTFNrWIODGR7ROsuwEAydcqoo4PRz00ub/kD9Wnibt7CJtT
xwrjDQIUkiOsZJrRBz9Wwl+/K2V7bC6BrwqAQ3Xi/Qbj+xM08bzW42bzi/ZJzxe5
6PragFlzzjCzQKjQIhOMOX6AiwYjL9RnXVMJ0tZQHtwt4TNgpyp9cHNZ4bqFLtBE
KBXp3GmkMuIds867VnCvUt8lg9gLs12V6+ao/vGbH0XLnyJS3RhuyS56G/UN6FCY
P0MKorKiOjenWicFiFy+dSougFVUlHJ3jgB/qKuyd5UMSncAFHLfj14nHrOPsPjn
kJvTdSCe7srabooiIIi1sWX/NV0aTVAErDdsFWtXCdVrzge5FGf7lv26Ns1K+2Em
uF2xXXh1W2wKIvmsY5OuJC6QFPLCnahjdvYxfBIVmSz2N9EzDxLFvWf/Gb0/ZyxM
Nhbalr5Jx5TaFw0IJvixlbfQeTPVFSjVtKimhLlnqDB2N0Ngfnc6DfmmPA43M1+c
4bLizyrZfPFYu8QqRk5mSo3rEoZgx5DhGMp2ZF7SPJMobZ4jQGAbCQsZnpzDccFh
0Gq7MlxPWXeWrJfeVwTq2H2/0zPN7IP3bpuCPsazZ607VfDOhRj4RgYS/gTyUMCv
KRKMeYVel3gbQ6oq8hHXUaeCA8gBKCik1uFL9/agplomBMUNwudDZk8TTCzZiuaW
P5WKk+XgVbjd8xZTsR9B2gCj3ULwPlIDFh5Tl/lm5E0ujZY0lDgwdIRWbVEhQvdp
Kye+U8kYr2XPoQgrlBW6/8BILhsg5uWuzTefgHdYskGGBHnLrTk7TiwQBsWsOBjZ
1om3XO1ib3Qn/+URVNdlJSJXgt0jTwKERDjmcKHlmWbRdzJY7kiP3CtqTtXFc9Qj
/0KUaZJtOJGF+r+zueVvXAbD6hJJwpMjjPjTqrBf+H9Vu/0zNaUrGHVhD4d3szv7
+LTYd+T1y2jfUftjv4/n9zrTQ9Zvw3WGc+UzwPOAgze9mewWZ2YkXOOxX+bPEq3P
YBycKTykOIN72YzCfWeXlDvC+audbO0Tu4IKRfNVkxTiemFUOt4cpYHcZuQWlwa4
jPhrAWBiGl3i8OEHJuPQ/dhYbFT3eVWH14g2X9MYcnxVnpEmq0/O8bbPnv+er7U9
lXKJkXwfOo4EjgQuRaVhNoSzCBN6jNbiHbX6Mw9AntkWXdgPuJDRsDD/ZMLtYSx9
41+CiiMi58X7Oy+fpLQVcgRILgwq5NmfqS77rCHZ47mQvCExsDP9D+y+g115xJTp
si/8WObwlsnOcmD5rpFFAuhOb0Pp/+ZyKv/m1JoKxE2+jaktVX2ueV2lEXaew3jy
Fqwh30WiPUCQihwM0SUZBrxr+68OTmn6D7Nrlg8ZKjDMstjHLZlNdXapV/QwWnAC
OvkvFXDupNPJuHNIOhF2rsNJlGNNJFgGiEg+CBpS5X3Qft6mFWze5W8oStWyYxtM
nxysFbxCmgvQGO71q3f+kRRbKFuRGY/iUxbhaHBpdqDSFdpYf3N8PQRSoI25pXWt
Bc1M7y06PEN5NhUQBQ/vQ9Vfa61VWF/qbSn4u4YoQg/LR+ojb9IXM1KWe82pr8FW
eMLfUOPWMxj2ZaqFWiYScP9RyGEl4knMtVNHzr0CJUpztdNiHpOTjnyu2RDSZjFr
OoRwN4o7t6IfWk2bxwD1EIkuyKUgLGSxRT4gzpq4hLQv5Nfb4vtK/xz1mNR+PDvd
mwPz/DC9+2bttnA03geencBS4gqtIYhzcedC2DqtDlAoKMYDZ0axwU0F/7HMh3St
maYhkf7jbG5uPXBx6Opb617tdFk4QDFl9RFg8MBxSTHCm2LFhBzfUxFxOurdxd2O
TR2Tb8VMZCGo6gMQ7iOFC/q2CGIKDTP7Fx5XonS7afl4ojcU8iTnuLKx7bpHvDWf
5PFzDAfwgjHzTOrp4rbgAAFokS+mCk5z/9i0D8I+AI10BIcmbKrbvPLHUmPUNEym
S3QT64YqgRXhzC4/yCvg2whrdHka4KaZC7a7Bt6cm4J5wTsaqk3rEOo3ln0688tA
XuPxNHTBfs7eb92KNN2FOfQQASj7Y+yCVZM7wSKGKJc4oCLpj4SOtyNw/WzrymYg
vu7dnnB/qKgHuV+st1P8s/T7uKaHf2helrEDGdjkM8CWYpjizBgSyqqmNonOpKCp
b6F2iZsLGGORKjNQ7mFMin3fv8PwBGwdsGgsc7XKFjW9udpfH8JOal7HCuRmiL8r
+jKbtLwbVN4RVvDuAU9rha+3NqEPFgTWBwhrsKVZZOkrxjZwX6nGr/HYJV8kEfiu
01QU/b/qwXJTfIH5Qa30ryyqqRX6/vl9Ost/+LBOHLUWEO8Or85BEpnZRnAQUauN
cl+VZXbUsL2RExUc5w7/I+mPWB+lxKSNdLsV8O1yMHToD7phdF7QP3OFYChEsmHc
eK0nD3SJdoRgnk71JHKMOo5qKX21v2L7DKYZ/oxv6qO63y2V9CeFZqiiiopj1QBW
cWlTqvuZmlYOCSlaOae8Jd3AcIaL/SB1v3/gUxDUvPk1JETh5bxaOWn+qaMRXik1
5GFVAg9IY8xwGk3NMWScvB6/usUZObSvTm4k6za4m5kkWDTgC7un3cZt2x4+I1z3
0nZ6uJ5KlgGdEz7FhhmuCvjj+WRhqWoXEWOBmvDJfbyrftSLtU2Tv3inHexYIwqL
P1BwKVbgpfSKz8Ms060srHr5PAfUdI9OsXLlF7FLsrdPc9EfBSn44NJOnDQgrHJ0
n3nDvXdLxY35xTynetkRTuxb2OJy46pLBWbY10T+UKXRHiDggszPeic26p6uK2+/
bkuhFsEKXVVmRO6uFQg6yXlIuyReNyKpFOUa2jiXq6HXrMTj7xJoJj0B3lUKES1Z
N9BYyfyMc/1SSSW2Twc7fycXRDkcc/FspI+mQphVlOZc5EEQ+7b2YAUvY2DF1c15
C5Wmmwh1VtZxXSrsye8JP3R6KpcwT6ebDc1UNQ4Ixtwhl/dL6LBsXt3NHUpGVQJo
ILOQJ2tqDyXxmr9z5sZCEyBA6Btsechu9iF9p6+x2BNWzeMhxEqkhaD5clBEo/AU
1UFCE+jmR//HQyXH9oHSEQDs9YsHWW3Yshd6+e8NWmeygccrfBTQhHY4MUgNSGtP
IKMTyTeurgltGzTKE78i1u3PRD7W6piDLLVUky0LpUsh6/3fK/ME7lNwmDGjXbK7
Btnex7UajWOcqued8aM6J6IugKu6olNO7+eGZZgdelaf+66U32rwrPudZ8rJV2AF
t/T6N3jwwx0JatdiD9Lm2tLxb/Lr3zMgy8C5IcM8p8RPxdZq7Ta5eZ0xisSKcz5F
vtAWQyk/GivTI46WTN5yR2SUACSflQGT6YitbJNQTx2f4eJ0uVnw4UF+DnPzO82j
tsVNr7IKr149XXCX0OWeMGbMGhv2T7d5M1ObBif/Z39jRydbeo2jj97O0Ar7ih7m
ny5ARpMTdLFJzhClpN6AgEy1kdW5PzdQBR1wNbykrUqNsAOGlZ/MKi+vr9Nu6rLd
SvLSelTa3CaPillcMHrtvBU/jTCD/SElclsuajlGdzcVgj63ahKVc00GaC1FvuXY
qTUGuXtCBAsHUR+AQHvvowCHp2BaiEOUOZWgm9SWB9i/5rrO+LfAhLz91go1HymB
gYUfHDTLv8GEMvxBRQLFO1ov0T2DiLq17fgb5pZfWkcNdl33+ixHz67j2ASgnACH
/zRAKaUMFuwhT3w/C1u3XBZQl0TBBikVKDtYPCAYTFEpDCNqXqIlWSl5SWuop1TT
wSD31mot9UEqUSea/EbGY93Q6uHfeaG3kq16LaHpdtW51/U1B50isEaaJIQQuTNg
kYhBnEIJ3pqt7yahzWK4UeEwTRNpwkIsBSGjVi3d04IbSJNBzB0RJ72JmbrVVOQN
SDolSwphHBcZEA2vqzWMX47EMomGTKkVMsluVde3y7DIPKnSkSQFCXNGrtswVPWN
S6UY6IAkOSOHH/Ey8A7a9yWnAZn2H2Vb+9Jpw+eYAbm3E5uweIG9WVdTPqpqa6TU
2T1/CCIdY+lF0Qu8L0hUh/aNjgbjqEKjkl88Ie9/OmUfOHGhAO12iAjO9juoin4E
9VJVikAcPm4wajMnx0ZP5TslZNpHczqvaVlADV/ULKw7HIudsCE0/Bg93aJr7LKJ
txjIBLWx3fvogzbgqQU4/4Q4tJuvE7OZJi6dbFN4ZRoGJnK1axIa5ismCjT/C+Kk
ARoxuOHUW80OoXRso4jhF4PwuGVVHbBnrybIqx/JF1f9ip5mTgGKZBOTqcDavorh
xzjUQ1tLFZ1YVi7piFjnmjf6L/oVHIyMAV95w1FUGJ2/gVtmfHQMLYreOhtbWcLq
znY7RZgsXUU6rMh1bPwnjxmBCF2mSOsZCPDLnOl/MfR3KliR8yOtvsVrGqqixnWS
40JQojiQxBOLZkZZMrg4+NAXH23rbi67KHPfZLyPAxr9E+iGzes43SuByRxNaRnJ
U1XB+IPSH4cSYCcC2TcxtYC7WMCUbk4fv9gtBxNhteH2luATMxVj5h8clEmUt5HB
nW/CTCSKKbjKzVJvKG7TCspXsdPxGPCDobkS52hwbPfNPjIuaZ266CpYfLMW9zXb
xZe1/+sx7At7D5FdCJFFNb8ggNCDAyVe+TvsvqYpPldnVYcAcgojn8irSZKGuAsJ
UMqX//nfFW0q/d7xiW/nSeYd55/qYfyOL0xdFDMafpiVMa1mY6q7h61VicoDrFCr
8nCQJyn+I5LQfGc6D8YNOw4WslJts39nrcHs3/Gxu5UH2WIfUlKJdVAlqKzQs5IS
YZEibejV9EvF3282FTIkSG/VKC6pFzxOmY7MQKZ9/6IZOpsVxHo7V1HhPZOnGg06
u96kG00oALewyd1rREtuIE2QAw3FTXoMEfJU+QnFmAAmEUpxG3uoL1gFCSQyULRo
Yl5wldDZ/5riy2kNeTJ5/TQkAhCPAkIqPKy2vWmowJEzUivdNYQC0Bu9t5QRYMjE
vW0LCszHhwP2+v70UZRdc6LmT2Wy/qjmNB6CYnQNf2B2j8Mf5idDJdz/8Bdq6bOn
dm7/sbj3NbMcKWpFZGW7fDl0Hjrp0SI+WsiyEk84IV9XfduS9IEGPVs/JKQk3e0B
Ciw9lLx1EVFqNYTTBwc9vwN0xmZSh2nVp1q0ToUbMsFQrzekUCDgNdjnT/tLRJsO
1uEuhuCzXbp3onwMyqafke5cCfklvW+CKLL+n5SQ2TTgllSaXw4IxalbICK0Arsn
z/tdl1PxOPWZKTLK1ORSHoQoTZe0tYk6yokGbOkMQxKTne2sCp0+D/H3Eh2SMtkU
d+z1oC/0tCdlI20CdnrbrBdFWY0ImySvUNtM0cD2chgUpHVoNsS+5comgrM7zZbO
aI9G86W7LfGHE8mgf6ZjIzOa0LT0kmG+fT4uvlh3JiD4d4I/LEfRj7ifJ17jmSfC
nr1HPsvdNvi24tXVQfyZ76Kk2PIcDTRJosC0ZWQ9voY6SrGfl0oY3BJgQVpmWqJc
KnGrn+CM6OB1RE4++XrbCx26XWoDuVCpVj8tWmUmYYYIdFboeJE9C9mlSbI3Kp0i
T2ds0iAhFmRdScVz3ZYntoQtZ8MAvvNDfrhsJdPMGhrvQt8HmsZvy1/repe+R2MT
9e9v//bF+b8i5iPhDvNhfF+p7aM4c/sMq7BtpOLpTP88/DHhMzTDNcDSmEcTJ9q7
HuhSAEtBuIccn3j/BXF8k5owZpBuWINPQmt8Zk7uHvo5ga0YGPjMJGOiRQJhGCHo
eiNQAOrHTiYeuhKY/AeAxXImciMx9djHYLO8ZhTlHYStr9FKZ1asMXjoLdso9esK
Dn+Y5y8G3ZrhxRqYGInL6IB4SXtrbXK2ZOn8DxwslbGa030TovnZWVIvCC35/tUH
VDjn2RkERJtBFzBl4Q4266Scuq893JKRM28yQPt+LDFobUjxRzTI5QwpD6IFPy5C
eVLnKolMUtphDySDIP5na1hvaEEgWew+yl6kuTlpG/MZiH2AkThM6OytjxAnZPjT
phgPeD3bhrjURa92SnztmHLLVdc/i4EFBPyT1lgzI0uXPBv3TjuvGzpDwu+2wuJc
3w67M9kXMYH+GNhZZrK0dLRd4QQrwZEUcpUDj4LiWUCrBNPmrZf3aDkQRHqy/UI8
6ATKXNt4Ep2yhG4wBoBTFDR2r6MEZA6eIm5CMNe358P/Uo5GGxhDgg6aLdLE2si6
CaWVHSvWmZb8taYuTCFRWMn6mKOm362Yt1ynfrqNYYujVscQG1EF7EfCHmhYaPug
BemHw516oPGximM9l+e6gCXnwmwS9wAC5Fr81CN6MhQ0tIfSY6H+OeQWQN4zkkXE
tXwf1kSxUv84rudjUxpjARZFJNcGBKlM/bp2mK9JCO50LsiuZhPGEBY6FQ0g8gvU
DwZwHBozh1X2q8GnRiCvvFQV3qIZKmqb6lHeWXa62hXNZKCIe1FOiDSw+Oi41kto
P3/L8kpwMjClARRTClXCEmzeBPTx/oJ4BNWUD1uFizBA4MIqJEJQS0F55itiPFMt
vprQX8DX4npOTi44blrvw7nUHS5RC10O69xfu9CiwV0a/DBosVQyd++KXIBBl3Hs
FMHuaGiUCk1SoMzPR8DGgtJyGROkWEbUMLUkyW29D70swItj7sJ7glPCpNbsfZCS
SlJjlpJmSRnjWdM2pl8+uk3K5Rxya0xFaNtx61xjZwBH0rxzH73VNFw4I0sKk02K
gNQDqBbiWvmjPC6sk360jivGX7jCCoPPT5tdKggbPm3EiNgfl4w7+U1XjWxisZEf
KxDoB1es2sgGlMt12RRh25kIWJZp4z+dwEol1bsZGFtu/IEpYtFlNrwsmz4706hn
4CBfmcQdqxnp40j8wgV3ypcx+CC+7Y/2IiXJyxrerOqGjn15Nhn3s3rjBo/Witn3
aDhgUz2+kEpRXkUvwMX858z7bXLXf4YAjKQ6UNyLi6UJDGMd7vam4B/FoN/0gGrk
tLHOSaMJxOK6cvtr9GtBO6dq0bEwLsN3HAOij11TjC0EuzKXWO1ueAVciVRLOvAJ
i1SbjGhDU6cm2pexob5AkjfPffuZpe96IQyl/v6X1hVqTdHuQtAkoV6PM0n/TqjW
mWNZDg7uQdFP9h/p02hasvE/0MQ4CRS3QpNOq12AJVWh3QnDsPXoVwLz8HYXWgZX
m4jrOgUAKqVMsRqnE5JzaWavAAH/JfYUxJS6iEkU50F7zV1n+JkoEc+W63/bF3HI
Yo3mWVDJ06JGBWeoiMsq0HFFq5ft/fip0lNtBY0M+IixdVJ0eDGsSOhSf5bfokop
8659K5mV1rVG5rmSR1viL7McOosQJO5QFFyFkDccDo9QmqouW1JsKJ3IqFuprcHe
ovqGm5ESh4zfrxVBL+a/k6Zlm4z4myHADGJA2369i8gJskkFq3FEzSBGCLWB4YX+
xCPNOtI/7pZMb3uDl/rQmDWwPaTFH7aQY9wph+RPu1NOmMMXlhWmmU/lcImVE7Tk
2MsqU66grH1UqNI+nbevEUpw7CTOLJlylHl6TZWHshjVHC/fEQp91i+3OBuQp5+D
YyAMifkhErK4a6Jw6r/uxpCdD6Rh5EhmORQ6527tEXivFmh85mbA/zxYygmQbnPu
bscagq9zt88L1eEJsLK4BYYjURBhu9jxgvN9G8oxqyaqX4Ms13QJS1a0eZeAgxII
mkC0BVCHol8glTpWPW01vDo6Ro5EHEyTKSnay7v0hEE1psJ79/q/ikZjEKVv+Tl0
B2CdX8argJvMhrHSE0dRv42rLw/42UjlEicwl26FPGFcI5oBo5qrAz63ZPR+ecWh
1A3IE8bwJe9tytztQEXKLjrU4aCFDd+UxQLkA6EnOSOOkbdIZkT/8B7ghiRNQcAW
a1IVr5jkbpUOIcGW7hyzGm1OUV3yRmzGODpKQzWs5F98L7YdOfG/LkYjv36r8YC4
s/qMMZyD9gyAl3GuaC74zetWj7MZaQ9PF/+GsipkSTcLJ+reNwvi2yH3x2qUyYhN
FjkpW3zXvxr7GmCC8wjcMpC64e2T3bghAFa+9AkNPBcCBZfT5PYT1ZvfgoxgbtIW
cqBlRtoGZLKGCCIDPnzRTaycDhBlwBgsZrvwqmAuRx+v6FZN7lOf1LthbyZU6/06
MTuIsgFerqd5XOe214UBlnO13X0h/0hOOBDAgNh/3gs9db5aohwkqADdSCrsjpe2
nfhrs38zyj8BYQvtCPQqogpu9ifub98yc7AXqZyeOwcGOFPW3xbTb5bfXyiNvcHG
wm0sP9/nXxB0SPkkEP728N/n1rhfQn8AYBg++uUAYKCocgYXJittr6HGzQDtpQOa
/kiT9c//OjPp6cdwo/zukY2DfZtNNAJpW4q2MMqX1VwabGwFF3xIkWtjwaJkyxkt
nV7sGv+B3GWFtxYwyGBIwh2R9ahBQ29pHw+1Sjkq4kbbE9pYznO06fWP+ylhp3Hi
8d2M26CUf2i1BsC1mkiK2eLRc8x0LAvovs8t5lCnqFEjTtyjuOQS6UgeoTkBbHjp
UwfHSbkGNdCH6iMwMwmfG5pyEcaN67C94clWy0VhpcmaJCSEsDHUhCdgxA9BL3Bp
SWMI8Nz4LC7OqADC0aa+1Ms5juJ8qFyzv6emJ4DzM8sfiFqoy+c4iieBUHD3bjE6
sllfhy4xJ9Xn9VZpVj4V25TwrqnO4QyBTvDRGi4849ExvQXgpUbxtKRMONfBcPQX
9nf8CTnzRIrXTXpULgCWlcqlsA1kCby94XwAoDKrxj0CPoBdp4o6NXUZ6iyMaGAJ
MDWuqmhPS7VxbtoUior75lxheZzBB5CJ58o4EsyiCQie3yN6O0c+9RU44bZU0A6/
/CL0gBrd/f0N2Q0QyFP0A9RrFlYqRqPOcXIw1rO7oJsF6P+cqa+UKv18ayhys9Xt
AHSzxNUP+eBBVWy4v8xgeaGSU+S5FWKln7SSYxcKXMljsl9TAuGMp+YXXsWk93eQ
uGYStePSxQOlKpNmL03vV5UlMWuvCEeS/uRm8KMMANZvHVqoab60/0EnnuQiavmD
8elnCcdCSm4ZSCmgzfuRlE9tswpkPKk3Os4XIntB01zz+0EgAUstl+MR6iyKSYiG
lOI227BZ4jgMBlQXaF+v3Q41J7+jwKFOGuzcntPFSCmtuz0hBARlBrnhkOB9AidC
wrja7jlgP/KFm6l1Yh5sVsM1LargMVBc3Y0x0V/z+7s0mBTfq0jJWM1uOjcdxxmc
KJ6GSd7u6Tn7hRCtsFzSBFcLToINOJ758LwgGOhMDwFXgELyuRlECXNh9HbpydP3
uGd0Y2FvlxQCyeOevBSVESWRpBQsglz9yiW0byIQI3cXrhhpf7hsujr/tDx4TgvF
ZyPphpiT4sHyVLRDv1+WraYOOWUioOAuCMUQ5pJG6fKA/JbsGqChsrtzwbBcMyAf
vohVpQnzsyNm6nUhvNq975ziCwqC+6kjsT9EvAi3D5+VVU07HB0ATvJZg1+n+dLa
837N0Zao1D4XKYoK8JBsSJsCh88dTidVW5cVrmxEpT7Vq336E7DuMqoe4GHFonhh
5Awnnsdrz4zWdChXcs8Afm/PEcbx342EwKa8K7u+oDxPDCumZyWypx44+z0ADZYd
LIhy7BUZUzejavIlP6zY0xyU0TGrG8y1RYGFQqGJj8giB2XfXKQManX8/b2wtye1
T+zrsPGqNdyzmAFWeSW3rOxK1gyN+6s5RE8hDg6Zl4bZduNQdd+wanH5sgNCnfP1
omMjUkbKQ7ekqL0NoFltTzsLk7La/8K1An3c4vV651JWQaxMNOcfDe3sVPOEj3YL
FqRTpU+UMIqVAYV1UJRRkwebS6bg1t3yhxh9yUJ4/6Hng4L7cRnf1IIZxtT9Pc0+
LZA2N3XPyVLwYNAlDJMBbwgtSKIHHgOHz8vp+Pdb+3yNZ0tJ7rzuXbDkWDpyLFSi
ZTgy2NPmc5U+74WuZY4y/Gbn5oA+WKPZ+5xXGD69mICumvYUijATy9Leaa7hSycI
pHMkENX18TPJzt+CQnnRBtbeE0RFgPKwMC+7KumwZ4rYpfh5mtU+wfs4g/oEJnYL
rHmE83wMotHYRXjmgKB2VCaM9JMym8gPOWvERlOAOEG6Q+wARr104s3cQCkAtsRS
x6ZX+6li2Lt3uOZMFHwnSad02zMgePHtRNvqvycP0Z5aivpPz2lUyY59nk8qGYpZ
+CfU/hR9sO0tjxa41NLu2GQBkMUDRMKJkz/3vaXA8abgvC0y4IylqSZ0l8QK25mS
zKYP40YJsCJzpu/YsImAx792wpDJ2uFtt4UgzBxxkphO0nW7lf93HgwSQ9AV6Rst
+5C331Yo6JQMVx+joUFMtt7U5i+wprHacVBh8ZWCP8BP1wAFDPl3ynE6YorLUex3
pa90tBvndEHYebXwEiWa3r+Edwkt8jhy9hH01NsMlHB91L1N1fxHXLvDEhiezBoO
iJEBSBIoU9fBoOz5QP4EGb/7SoNaOBpjg4+5iGK8l6VXdcAJ31m847P2Inj4BAbI
1WivXmf8oS7iMqEh7IPNN/DKrJQu6u50dP/K5c5ajmiG1Cy98VCW/zP8HgHUGuvn
j31lvlqEIKBq4WjRMYumOUzoTmmL4j8ZJO+bE4hJdOv467+xH+tqsw9KeiSAaByr
GRMVfa0IgWkinE+x6aiTG3RKrdz4xs/6lyMd3D93pSYEdw4PwbG97SoneKi8IVVr
+Ld3jRt73vG5uLlY8/OkGnnL5b+IWn9nylxxfqkRBEHqCwSFc3gDMerlSnogATX9
/qLW25+Cb5H/LXylofplE65zWR7khf6ZCk54f4XZ6pYVOmbrh+bN0lt3M6Fyt624
lTnZTrXvO8TPeVyFdJPWBGIsSfzggGdiql+jsByx7HOWYcD27v8vqdPikaWFduus
Uvwq2NODe5uFYG6TJ7KnAs1jvGH8Kp9d/nZT/yCTv1YyztYXgqBF6D/e3GGSvlxV
DK6nlnpyx4hfNeoQMC6iWNnTboak3frzjMiCQwCksjqS8PEQU8FgYo5MrQbsieQo
Kca/dx4lObovnYf25IOmW+XVZICjEhAdrrqodfTwLxZdTwH1Q2aL+O9pYKjEBroa
LZ1LfV+0LZs6poZdawAI+uuMwZ/MSoI9E5JaVxRxL6iAFQGgwNuTGsj2pwGHAaOU
M6FJnVfFM+NwbuxuSPPewpS5PpUhfY0k8we+soUxL74e1SeWi8wkXj/5v8Lw5FIX
DmKSkBt+Iq7nFiw5u92eLcyRG5hEysxliDfFkhaW/5hduCIu9JoLpZrgXos7HfVc
zWQXPK5A1B1A0adxeRvzbkIRW4TFWAm2CP1DCVM++p50DzJC0yS9AgfntId0+/Sw
Ndh9rCtC56vUDqIZkiUEbeVi7n3H/Hz+rUTVeoxJgfNikUbl1gyPPkUwsfGDi3pR
gZErFyQMUwWMApk0OkVrUwYw3LmpYIBum7VASkdWshbpTVTpOy9UjQfPsorQXikm
rWrpi3QCeDaseJ1vgaNpXyMyy0XSseEfT8/0Kq9EFnFKNPyiUGKLqq6VfAj9//4A
IAgQh2xvcXyR2BkBFZEgRO5rIH3elbygUpUlFWW1wrZxhqYIZY5rsvsl4XzOlMfS
49cQBqNBLm7z18thbPrI0/T5r+JZ5bIwVFs8edYgZB9FWyoQKUObpLr9v5mB4i3g
JWKjjwr1Ej56VhwqdKcmTmVqRrPIOkHgb0nIYOaq08HUcPe5F95w5vtdRJzhJSVy
iYsMsSqkB0Uff5hFW6IZPtbgs1s95qc8md0fQAThU+7Ba8mIXabroX60xVX2vPte
PzJVpms28+ZpHvUKA/xUyBzpO0UeuH6dVkzcKXnDbB2a+1vwjVfESZMOTefCOjY6
iTJg+Lo9mVI57ugFlWyyJxvGZ2r1JZWPVIJzHYuVq+YTOIUBQ+SLSWdYexP+i+Pf
Fo7J93x8ssf4zev80LSMhOu4KVCfcz00dfW8MR/ddiJYG0dAK62bd5ASl3cADqt2
ZlRwRrYuSyATQ3CaSgupER8ip5UCxrQuPeZ09TC+UMruuc2ZjJyeHnCmjHbgksyD
8pOxtENdInSszaGiksidb01stexX8Mvlp0s0QA5SMdC9zk2HhdUlgWHjJb1X3hRH
KBy2FBBn/SfbGgX3pvSblNhAMpnZGNKytC0nIq8jwdEj7YUp98tQQPkD5lPGf29F
Zgvs+t9DkbkZAIPICLijMt63NIPpFeZ2jP1SqlxR4D7zukbbgdP0sW8AFXa0wRPu
iQk0qGAmDbALAMqTCdY3ViySkvNU/tW3/yl23wOzV83KrRmo5cocN8siHdbwZ5Oj
YeVMM7lTI19UbHZGjdd+GDLMWXm77d0u8Cxrx+J4HmxP2Whv2GNwiIfA7+bcK2LB
C9sfcjMzAXXdPL2hlVzUQqzfu3x2Bt4Q8RXmhyQXGJNLwWisF4AdfxYkRY52sRtl
bXPc20KT+zxwnLOtkDfWe9BUD8oUSTEkDk+E12dngUK28KkPg4f2IUr8KC5V77GS
S5SYTZkrPclHpRv0lsMBPBzTcNpthF/V/2yB40TxWdnqNCH7H6HNy25DrCoPDGrM
B7ke/V0ybPCBGlqDO/rwa8riDCSw2UC/Wbov863EbkTAQxSN85SEYlF7l8z6frpc
AXvDO09NigCrNnTIO79gKb/e4ex8GNVZYXOQSQ7fKuk6EBp/qbrd7V0ZK/5f9/3g
ys77rhglHfWFIsKMveacPTOI7lOOiLSxuRA5xWP8yFMndqdS19ulhD77VP+Iywcj
X0WYOQz7IXmm3kDQAEaC4naruE7G30+9pBG9enEqaBy161RxTEr84siCagNYjlfb
3JwbxSSCbKeZIqkcu5Y1AOVHoog3+JD29qYmakvAuiR0DncxX8r27tzTMrKb+fzh
uvwbu9PY8cftIMdNa+HEamQ7wGrFcguuY5W4L9RJYBWfkxrXTSQ4AMe1Ku1s+Z4N
QYSkRLodRYiFKnq3Yal+scCOcyRUtt+Q6lyF8z+unHbfaZtWBO3mrH9ZbsQCtA+R
BpK3WGwd4pDKv8Cno57IIKheM6hMpHmePf0a9ffNXFcka4aiwIJTIFK+IrR0EdeT
7Kros96Jqfy6GN+PiKay4q8i6bmwUdKNHRY/2J9lqqz5+eU/8z++PrDxc4AGubCr
07BaPSfvQKe7U+P0jf0r4y6zVz233BCiVBfmc6FwMrBew6z3gblAcllr/FpWXtB5
lhdDziDecoQ9vi2l7ivsjklQ+JDF69ej4a3lSM/PmXJe0RRYLMDzwc3m42YWTu5f
Ri3TWYQnkFkod5XWrGGrzhSpNwgF6ObrQrfOV8BW4PkyxGhEFLpGGrA3P0vJdnNy
DR1Yd0m9ZEfuNTT1ABa4IPUA0dRL7YiftAtGABBBmFem2m51v7JiQCKCoSWE+8Z2
N1NjOkhTF6tLAtwQ/E/e+KHEYp5Ka9U+ooi0dw8FmVvE/8mVe1xaG9ridC9VdGX3
0fYEESseR4kizfR/611IZebR/YLolRPUH49j6I+flZEAZmwduZwpt49IVI+ij0Cr
+oe7TQZS2BnIqRpBJSQuoD1O8BT79QYwyAmm9243N+hAN6o+UW0wUQzMGbFTcyt4
tIfBPXbcX6mUZIr4ecsS6yuo+DkZnjbwtm/Ku/7LIm29gcNyI3x7mtHvABR9IOE6
FDZ6PGnaIcYIzyh7EReVQbBpB0BnQphsaVOTUAD2FA1Q6OwhDY7LZfIDn1fRNQ7k
SjLxSdsnah6J463IlMpadrKMcWk3+thky1/MFGWUz5pj6rZ6cgifRsv53DF9A+a5
jsLTevo0nc5/1J0TBUWk2UnoYHrxJ6JIJZ40lXne8iTClAsiLvg3TvIi+XMDFzmI
bXmRKu9ONyEzLH4U++25rvIfcak4GYtK2obKVkgCrWsa27747HPNo2Rg8z8Bebc+
r9FyovnOO1abslrv6DM+BjD4jlYKHuhq/3YFk/PRoJbWdk3itHUN5iSiwsSaJZkK
TdKvgWqH0IiU3t3FQ712ZGUMO2XtXWNwmz4eppCUrXW+adMbqsYIEIHXtAjtDYVX
z/eb/Uwdkw7zxeizDWcAPEfyQ+q7JcIdE25BpWz/g331cmcPMzsdQFPEF6GXvZeC
oPyh7QUupuTCHPbpW3yG7sVF/JNvxgmmqCPHDYKkpvOgLqjrH7cLsuseGTvokwR/
kTQbuc5Yr6e6iWEo9bIx3WFgUwbPEhe9OdSXKCoJ+Aewrc/yX6yeQBdsuaz+0OHl
nzM457AHXQmu0dQgHxCSnp4QftsluV74jK1T+j4SjAYKzo5wafpdKRbyVdEx9ROG
4R3mVp3PjTZDZ7tx7lHMbjlUssNaDAw+Dl+L4EGMlME0ENAW7AposBpwDCeIT/CF
L+ft0V1zHaYOW+6+ilVHTtlpzxIqbY3Rc8piyyu2ys0O37ahWfjvuLc7RxxkOShG
KwTnh22fmMLDcX8aSI2aYFhq3B+UOc6bZkp372aXlnRWJlYn9rFlC57Wfze3H0pB
7M63KP4goZs1r7dNMMoRYGfUOQ0qBn5wRqBcI6MmjNzfYN+EokeenMXIhxQxlB4g
LyT3Q3HplVwLgs3cTzh3xRu8wZIe01WZNvxzSSmCKrA2sECp9oLVGL4JdmmJN8mZ
oXVpn4Jqled8Ld/zyjEKS7ZfY4akpOUEtysZoTLg3W8rTd7efgZIGO465zLj6Prv
XYV1AFlFw0gYCFJxgE5H+t0Nq043c0eqdAhuRj7hp5M/mS3+hmJwewQz1h+IYjiQ
C5lDMN6p423wg93nvzwRzYilhgDF251NGrzNbGk9QoL3kGe7AMU6rjDjZ/f9XFxk
GBqF1lByIk7U5zINR/WEp1KK0A1s6/tQG18qOppNoTd+wZo6yQILoP2sNr+0RetJ
AuPcQH7KwMKpYafNqlfxn+iDgdzAfN4Z0I9WnMza74p+P4UNaclUSS4mKvvc660S
R8jb1pM/97K70odjf5o661YJVcqECXOVDKJNurmlXCGvli561kxKUKIKIyYmoYWK
ZiksXPQUVdsBhp04fpLDoxZRCiIgpNZtB/J67lWymGBD71Q9GVigvY/phGFHkKfP
keD07QrUGgeJ0+D3B9yUnewSxot6GdPhg2yWHq9+AjYvjbPzUHktlQcvxkeXjAMq
px/+U2R6LpvcWSwRqpCqMM0kZq6OFyFebwHGIreWc1LQmeIpqAQ9kRrCkDS+zXJ3
H8mNkEK0dRoxaNG/lPKpSNg2yNVPym/r6akG+VTZcl4OzHPXSozF7sR0cmSkRJvV
H3dJgW4kym3esep9wmtHd1oPbd/tdz291yZpROFUL4vFAsX+4VzanILZ4e9fyPle
EDDw8Lg7qL2eUx8GslxFHjk4reIH7pQYh9ZaOnlZ8tR98xN+/exVdCTquZYaXm8F
tEz/wVUgP6IXjhdIWTWRZYRlsV259D/SC+7tEbFM7k1OHb+IC3H053fPMcyQ7ChX
YHeLeA2eoewnzWuWDYQTl4+hO7oCe87YiX3FQm1BF5f32VvFnw1CaS1X7gGAmLeD
r6qfkb8evl/CTqSFAR+94/ahaxxXfxrff8mmLno0J44xSGOBzVNhdGGALOI7tlr9
gKI/TBRYy5M7jd2r6YZK7xcyz/UnZ6Yt9Wdj5Yeu1kMDsmAYpAwLvmf+zyVd+/Vn
OzSZtA3eNT2VouGSnR0onMTAGmH0crF7VXrfM5z1/kLEXugxoZqruxo5iM7v0gYZ
VHCNXFDvHdZhv7RhIf+3jnMP0092p6gY31L8IfbGC+xf/I9xbXaF0S+PSsHnW74u
RqrJzJm3/LqRo7ACqheZK+8B9YJacf0ARssTPomYaaeC5j9blE05n8bowFzbS36q
YS5q//NeS265a7lLmPYd8fsBen7VSmCE1PCv1FQy6SfurbxU0MZXk0mbh4UgbPiq
7VJBtAv3p5TxcrzRQm1MmBS3KsaQ8Hb43JZL2TZrGDLp7jqM23RHdfhaXe7RW199
OJLME7TrCS02/AefUjNH28m+IGUZeDwcgC3ed/K1vgh0Z4IWWssnxd7tRxd8hz+a
ygSo7z/r069UoXgr2AokmqVcF6BGadNxmd7JTc86+M7AV946ApJT/eCQjpAhYEgx
P3PWfJzg2wHgGN5/VTiu3v0qLPsXvgWskuYrVYfzXoQfyaaDd+mwUZ8waIv/sLSe
z8nwlpptYXEoI2ee6s6nXXbM8LijJXvIEld5qGWCedz9lrx9SrKJHi8cTeC6m1vU
WjP2Cuiic9S8OoFmvdsMYpCLupT7DnVg6p2BqC1XXrEpmTlSv5i+Tk6DgEK7opWY
/wZtGsjdKG21QEY3i/ROIcXq8nRY2jqzwm2AlqWoSrFKDIvPqytu93vYLu+WBEp5
NH9/z52KlUCrlC57BR24wXc/MHhkYJiWonNKUpZ+5dBgGNf6G+b5IVvQmTtFZL3n
Tqps82f3ecRDMsqO3KYpMUNLMIu6JY66i7aKGUiJaMF2ZR5HxM1PcKF0Kzhg107j
8VsHOKG1RSSPdLHLmRsegI44Lm4mrsbVafTcNw2Uau/Pn1uIavXWgZ+M1aQQUtOK
M4+2Gf1KqvYj2UIk57AcJalAD0Q3vNDtDmwFv9Fqf4KxwLOjlNYNvSv+/9ueOrYv
JsFRTsj8Hkqo03wFr8wDlkYowqi1TUMh7+1CzfoUw+FMCcHc0hujjBRvk75mE3DR
To4fCSa6wwjjk4M/RTknSNrm+wsek77qWfKNXcuy8uwmXQrD/CWpqbOKYVWGRyIR
R4ay+1xRPQBtcRhSN0JFV20/g9iiCuA5m+Io4vZooK1IRqkKyNwKYAciOSiH9/6G
ETbVGyA0k2tGtmIxh0OZeK4z3u2S0wl4Eiyp/t8VaeiJbCgIbeL3H8IBqgGrgdbV
j8D2jNOWeJzSpFnlRisClNvHmsV/6n5C1fUiH+FhQFil8ck5s0bThYLIDPVTdpSD
vsKHOV6Wh8B0QJTuyfEOFf5xulWRWh64G+YV3RrNR0dcOk7BQXkhvfdfn6g7tfQC
kOTvGbVFVxiW2iZEgFH6TdgjkAcCUfEDwca02pSc+yYyxVLGS6bY4d1/copnlSeL
KeFjsK9hBGF5coGmgHwCBGdpAlBEBmfvOHOUQ0YFGUyuYKxjbVvIM9WqMmSvsG5x
FRqsLzRuPMsdFYZyAD79Ys+YSwUmkXTfjPPWyb4eDPuKzOCP1ZoyH0B2eRQiHbyd
mcv0gLcgw+QS+Gr4c2JhIDjosGam4q5r7DA2Wvisli/13y2MBAcPywWVQFTohci1
l0ZIcIEYBQeR++2ud80a7HUHzMbc3bopfs8+kgj7vU8ubkF9C7EuyQbmshuYjQor
i2H4cM20AzOuxzY/WR+wqdebSyBNk58iZR5YJzwuSo7OhcU4C1UJGTOYjs9dKSwo
l3ErviAMiWAhyyiFLAG4QPvMXZM1hHpJkn8DxuK/qpETQI16PW2liqro40evCuZs
YPnoGJ1RZFQ2c/12TPcE5cZayDdRRGFRA2VBQ8Jwtp/odnNMuVVtrxN+bzstyDf4
VFZbSg7fwoJj98D4XRsviDqsQMrT3iEr7ESWo4kUup2UMd5L3isKKEyB2uk/QelI
/y7TMtAf1uUkEGttcykEhxH81Un0JZaDvctKqmbLNOKwNNev+CzgotMmeAsaEnbd
4sSPQ005PnqR6PH/Z73Pp4V+2qyC7xYaytxMmPtzK388+mYCP3ROA9VGWGmVGaFk
gk8+uIXWWDUrRHOJW2AB8drBfrIBxInHmiJX1DXffyvHqM7/lSvGHNELgJIHIRgj
PAnTz+oPrJ9r5lqEvEwZuvsgLyUQWl+lz4kEmRfPst6rHdYDoNcQARtEPHF2s0tv
X2CPWUUB2HAKeYbaMOYqPnAZL256lSS9z/XyPagRrEK4Ji1VkY2Y48Mug+4ZFMqk
hhigGbLD5aqImWx7dhaqQidclFWS1S/YAJjruBTHsotH32Q1HttyHz6jn5C+rh5U
cH8vh/onbtdpnBt+uNLMioN8EkXEgZLtKcBu3+F2fPYjpnAgSRl32JKDIVZhZXHh
u5JQBLmhlxnQ9W1UZrem8XYpvuXUKIXK3lrav26s35RQjC6fUyKSrneErDusMTp1
dFdTOS6EaYE3wezY4nVXYIw3Pte3QPrIPcQgIXh5qJ5vBMspu8eG9kcyj+jHTSu1
DgLfFgaHV9tyzwfIGRNw96tmTa9vO+gV+wC/ltehK52OErgPUAqQqKX3M9Os2AIE
X4ujXBoxDfhoUjoAF0T0pJCwwccauyP6A06ZfnOx1D9IrNJhqwZk0J3jZ5RT03Lp
SypDyJnLFWzCZK41Mgq9qlDRUlSS2Iw4dXQ0JAN07sUbxlywMNpZPLAOlSf4wHno
uTDj04Njv8MjytsQKg9k9s1dqsFXo6s1VTDP2nuTfVqxeJX1WRNQI/O532zZzcRj
vc3ZhIV031xoxtM7gTOOkkKSZX52MT/Cdc0PgSKviSh3Du7EaTy4jFs7TeRXy77B
QHG3q2IH9+bBcqzki595ZYSg8HS8hOL5JMdRjdCzsZvAHNu6Gxru0PW8n2wJH4jA
7flB7pW5CDgrkQ4/ytvlHxg8X1mNu2GT2Yx7sUwz5pcZoKEySsYujV6l8oP1vXwt
NCwDcfzpSD6rovsQNkZWFXsmIZsWI8AXYPQ2+BoGyNmnmEB4xeSrX2lhPL8GNb2p
ijlzeg/iqaXomqGL9gZZxA5LlwaU/pbWgZupiJK69SZJN3tTLJJ0QSun3aJi3YE1
h2nJMgFfbOZdxIg00ayexu8ew2Z58ti58JnN7PExHu7PG7BBsY/CHjQaTLg5/3/7
j/FJkuCh77zq5my+VzBzOhVc4XZEiyirVzYUDqPBIDpUJDswlVgRkuCgX2jrtCBk
hSuQ2m8jtjJOS3xqPS7JMOkr7c1cmJP354nYnH6JEjzu11Qs5Lb3DtyWfC7tXTAa
Uvti1OSIXA1+3cewFxp2bCrABDLqIso+Fr2VNWZKH+UcHDob8SChhwo47pnDY+dv
BUSkRdb36t8743x74U2EqkWNPEUB8zV7h0ngnhUqEyQIgEEmvtp02fLMBAHt0Ds8
8/CLMvPi4RIRlBwtQTaWM+caTnGg/VeeRmRrcdgiBCA4QUBkBcz0dP1FknvxxglV
u6EbQARW8pr0BUumyg9yeZfwA33NkQTlw58B4oUs8LblPSzfijE+VArtkOdvT+RA
mzVTCHe6GVl3ZiVWmHkSHXPt0Hw78VnfQhH8k/D/UJ3gpaO5tazvvSjFNYDGmpYB
6oUvcbx85HXavIps0ikjjDjfsIuuSwwRo3Mm/7IsT/NsZO/jARInBZRN1VjN6TA7
iDnuVXA1RY6tV/UHodsiZj/z7ek+nTqFXklLjJ+ENGYuJnyak4QQO77u6Jvl94lA
7qP7Wfuk5ng7dFcNzEk7NKyIEAazl8C5p9SNHWNH6O2IcqV6Ls6XRtHfS8T2xErs
0EOliZjCUSi+uiy7aTro/2fH3ZG9YdXOACFuRBR7cjnqTUIc9kBV605+zLuCl12J
36aIQBN48PEIcscKNF7gSR3OIx+viTPZPYB6tVm+PkDs3jVH4LCFxS1RB4j7GhW9
Qzkwa9sCrL1vQp/WDk9k732bY1yz7Fxpgf66JeRNbLyldBjP/yzBp++O6vDD3kof
V2HUHwVyEROYbgRHqtvxFs10yqn/hqI1Iry7PYJzSbW7zErLq6699yUpk4L9oLNU
GUT374uKcbapnP4sP0xBxGjEE7rxXxc8LHpoHxYeQadhFxpi51u/faKNSQXZbqKO
z08JSwFF2MIoWaEZ1Rv5PCgpB2D/eQHnbIiFk8FnUifG+ffawrwrujEHzcsWPkxH
ehwAdShQx4T4yw0MKx9k1s5x+dAEXQgWMiY5EyZsT0fGFDFdsKVtMVU979FEFB8Q
gzMA7wNrFW3uodWVVPX3+le4j+zL9GuJ7i9bGuI2gCQnBxdzacPQVSK65Zs+ghhu
ug7U+E9voIQr9pwHDJBja7EUcvm6x0QOHqtrCTOVwbHc5X3Sn7bv59+r71YcK84b
axSxYUE7mAEAAOIQsELeCp0NSEpI6bZHH5mhxL9EbYdyKV5SAx0OLoAlMn0uEdNZ
09ImoDtX98sw5tcYb0DgkZeGG96d5LvwkMwjOfIBRxXkSg+zCxXJIMpZMIMjl2sm
Fi5eRDapEC/rGc+lSJO7BsGNjunkJZXufqnXKdXWPYB3CrnNF7kC0ABnGmNy98pJ
4U/ou47rZuqkAUPu5nWpN/W1/lNvmm0Vy3DCIgUzN60FRV9EX3L/cxBJCPIpgDOO
wqVBVECVDy0eFALvvXNeaUc44J7GvwtNJjkLhLrD6A1/kadQyAtrfs9aRiTPMvmi
OeV4QkH+EPT2PRZkTrl8H981lwTY7l036nD5NmKaPOdm976RMN8gnlfDq0ZfLqD6
gyIBQ3BSiwavXVXNAGkk1WJSyE5VWJS/+DHgfy3SGDWHPibUzUJ1d0jnCeXwozw+
aE078Vnd6LPs/dBaey5sEA3DSzbsoid9r7wKW8Lvp7bGuOad+E9LYCBat7RauaRG
JtubapWmBOpuR1UYotvvfOeYaVIytym678lO6XQq4XrRiS+c3M46goZx0BsPF4Ed
SQ9G/eAeb3fpGxcNBvV3sF/z5fkfAd9mpCCvIbWhvRmZQDXMciTD1reD5aWjLfWm
LjY1jAkub2+v+KkTA+3rlSG0e+v1omAlYAWl4bLfE6BCnb8olUtkBtnwbik7jaWL
XkV96GPKlbCbWz/0gQmQHJdGCLpikpePSflbyZLITk1kx0kWR7gjxEX8f2QwLBHt
ukYmWl2JiDPp2T7PihxVdpd0yMBobw76LcQEFCgdw7CoiGpBQzJ2VR5bUszpzXrn
xS7S04dG8BxLiyI//cSk7l1xidqdAXVn/9RH1orID7MINwD1dj+wAeus5LJbxJX4
B7PAzQYavUxzs5SMmIBF2Tq2kTlKbxjeAcclIE8QZKtIcxCDV1qYEcqjxVJATll8
g2/HdcxxD37scbvLxJy5IFs6wst4P3VqsWPATcdmWofMpkKiTrTWEj3ltmjn/DVO
iowFCuXYdTyGjqxpR/SB4RObMA6IzxKIOyUcPmpCXldgcXGbnXPE7ns1ZuoFVUEF
Kr/f4euYAvCOTFZVz+dInuU/+HQN4731/M5flJwlL+kH5DtxzFovhh4kLCNmi1vA
j63WNoBcuJkpLItIQ3MYpKjERr4iNGp77BEEFJf9SfDJRbk5HKlHInqeJ43bVhaH
EDQqxYAobttk/VMzcC87euyiQQbmZnsLnSI6C0NhdFDT54SrAg37w2LmZxsV5Xwh
G1PKqUS6zTwhwamzN8TGWA27AP9vEo64Lq1i72AJUbmqopeXrybQNp6p/LHlvGZQ
EvdIHGYVNIUKGBeC+Otd2mzxCCORvS7DpypBrNsNl8wOsP617I0YzFqsxORJkHfs
rOOVhXr38iH/s800WYXIC1RqGuTM7zKaooKGoW+OfxCurNq4yOY4bzQeraneKVZt
AFqgcgOwtD8ouNNilc+JXF0JHqHdFe1eCn2uswfm+eOuoMhIQLgCo9+i0yqqA3vI
z+jbhubEunvilMk1kXqiQtw5wKn0t09h1B47LxH+wV+qmeIEpJqD2i4qPAehev2V
Bj2phydf9RCWPFS7D65JOgdJ5ofx/c2xG/moRD5VDdvqOqDPgY8brbzBP4iyVzM8
dtV4dwZsN0IJ8IQ+bo56SO5BZerAUB8FmMgvOVJeZz0LCt2addEq0k2ny3T2Al9l
NUszDZHy6fZQ9hLAXMDFzUT3hAxZSj9ubxTmRclqMi4ux/B3mhwoRJaLEpzqSwqc
sqEw5jrkqvrvkiWjoFAQaZ+X9PTYmkZu7U7Sy4KLqgw7QbJovo+/HAssbAjfghzQ
zjCMRxm28uxlOTvOsLKtJR1jrDCcg5GBZaHLvecMlj8tXY9aRTPdJDl9DGeur0jb
/znVswKcYFWIxCSDyDX3K/guOwbghg66Qp0dvF0vfALyAsEqZ6wyFtz3P7xtnAkU
degu10fJXPHOv5s9KWUXNQQMS4J4prmVVaI/YY8m+nY/tFs1pG5gUkmy/swdC/uT
PBjJ0DoB69t0iQaG/BqqclapFkExxQjXhF+3ra3BgKk0RAxswRRO1rP4eJvGSUmo
OJAis0ujBu+k2RdBx/h0fNbxRPJS4waKmXoQnocdIutmCiU9qSyu1RLToH3o5SXj
Rsc98Pp45etgTJWwjqcxX+2PGugALLvjIp+zLDrWORzJtALy5hLbjZiz17C3ssKp
pOWgZC67Gd/gX3P5aGvUADZck2PUW39wiflcC1N+X1gQfeSshvqVLgcp+oJ8OAsB
hRhNi10VhDxW8vRM5Y1srG0D61or++l6bcXw5PB5lpzIhX57uphxaNRWLCl3p/xe
Wtt39UqDmTrT2jc0dNLSBxgD2gqx0xXZiHLXflseXsKx529Cdj3s9Izwo1pARDdq
KXY0s6IFFE9i+pALShgaiKSK8IKCZbE7tDtfLRkpJq6T2tnEXfFO2FwQHueaOc7W
q+F0oUNwKaeWvkRObosG+zNncrtjaXu2/+Kb9n9Fjn1rYIEB7ur92IfQgWPNt9A4
t2x2VWHksz7LQCYvmFgQJmAk8JIC8bqCIqk4Ak3zM9F6utoJVKBEs5pSopC4PQO3
zLKyD1ypJYpAxFgOhwN1ukoaGWKaTDSr206f0TuhypC06nCWYJ5gpsgcAroNWti3
3HppQPjVP8SMKKpGlP8xddxpfvAQs2UFq28DdUXICbz7/fP96wH0qNJqcEuk56zP
WuF4+ciDXnXGFhDKte5TxXNH2bosyYaLxRAL4C345B0gNhw8Du0SiyWYJZPWALlr
+OfCWUt3km5KkxHYFPu2oH152lrTMWRj45WEVG0FbFsjJLd03MgE8jV8Cjf6vkRT
9zZ0wKjRlwiPoR/jITyuaTX3IYiPFW6o+oh4nuiH6iqrouwxLPo8Ursw8DpL/y4Q
9dm9pAns/g2P0LDwyTnP9g5LgrsCFe4D73OQlj18u1pTPhA2YEGW9p1ndQMRVzHe
0d03HrhXHyqdQ6Ehc6AkTJT4Mw3bE5/ejagSVPUXTWfSCWmGVdtwWq4HnJkoeuSv
Xt7/+NUHgsbNqBcfDj78cHM8YdnV1tkB+FKSWW3Ve7iRg4Rl8dqhNzgP7a8X2USE
j7qoRWZitBnGEn5o5NjQfkj/dpTRx8uywZHtDfjUQJs/00TsvEWQRdgBQisSORwZ
LfSWnH36GhEgaXoZnx/efr8W42iyn2LdbXNYwaJyZnoNdA/B4nU/xFnLoUrs00gC
lB92pd5EUmcpwC8/luWTDBiq7z0FDpnNIKyrkdzRRC0uQ+49Rv8QEYiHZhDJuY6R
xPbJhpVI6xPz75E+d1viTHaHW7IE8+1ulJIrOXx5ra9tr3nsl5Ru7dVU8RWqwWVm
q0esWvOOkNaG/5gzKb81mz+vs4tqMwk/SssVXl4xhukaetM/fmOOtlCdFBUneICo
wyH5Wn3ud8ZHs65tkssTTU62Xd0cBMoYSptjtSLIZSWB9KQxUKUqi/xJ2jpZWcho
aGwh6ee7nnnLrHWncU0LbXeL7HMvKSdzw41sYQ5iWh5RboJLSXWdmQRQa+xpEC3A
Fgh722xMpyHvFrM6EjQDhyS+sl6+K662gBk4EaRYW3klNcqT0qjIbqVwFRXbHqLK
w0cp7qPTsYJsK5+5+W/1V9cNNhkUBQITJdvEMMnmhyzwjOjVEET2pLAnEhsfZ288
zLyH6/w7nNQNmck8I/m6xjUaRXOt3v74qOX9lO0BZsvP5u/CDJ01XkGYDsYqQuQT
x+IvCZQA8mND+TtSwyRR9QxA6osSPy8Y99VdVanUCollxJIHkh38Ir4F9s3KyHvc
uHTf1lDw8tSVgPgy9Tpn3bEhukV5G3eq68tXfaVmiX4rLFeIqX1yivrHtRQsNEqM
H1clbyNjGtp398IP31VntjpVV2GYlePmMzCvaDUPkvNAXaqGOEYJ4qbq3re9SapX
N4i6RohCZOlTw/INxKchGonoumhZw38O1OAruNNziA7hKl2o7+JALeIuChrO7kSa
TgpSMyJxGrM0+X5gz78BBPquqq/tobPwp7oZ2YinQZ6fK+Hi7ms9M9eP0tCDfpp5
LGDQzQPKJ8srkpexqXSWvGqIVRH01ZZGIslQF/5ICT4xx9U61cIrkMH+Mhw72CaB
IyDUnE1ts5VKnfaNHwhfn3NNORwbcU5arziFe7kq/bhNtTHE4ompF4fJ9o+AUjSS
tlKYZwrJ25w4KUiAfxSKhCr47kjAfT2Ax9bB8iTGPd4CcCr6YMHzEkYjI72aycYy
lxhmnrFqUjNeiXdxpfUhEY5BfVdJ+1B+319k0fWgW9SxaDmWSDazlsbI8FdWoihE
Mw2klB8xRHpQZQKxJpHWFBVPQnKGu8ul3DOtZ8QTtj/T5K+hg6D7cnMX65E6nuPU
Jg2cU6518/jjVQL6MSc32XaTcxeNHIkqFAkWwAYSTtSJDafD3o7B+3/U96iNzmI4
G0B4RXeCtkaBxuKks7UMYdl3fRpqe+Vwtpq/UbM2XyT1n0lmqGS4XRHW2tCvalNu
dZkBpmwAwP+SQXz3O96TLuU+OpAlq4smWTPZJImcykR+K59eR7vby2kIeocZyEC/
ksLsDohU3cRCzrakWOHMbxWXx2xuz0ShMUWPtqGC4yhVW97zs0Zhkg31O0U6lXOT
YOfVgZ0zoWwJvBTxo+rX1vo0wO2fzSrIFaghH+b4bTwMOgwnhCojsNL3L2WQyonc
KyVqxeR0P4KaPYjrXU++F/eXiXTcDkO3fKfFVrLPZVlWHKHdykoa+kysuKmpp/S9
aDqZSuGfwhc5wBc5OhcCYaaGT00AgJRWoXBLWhEkbTiT31zVbWXDuzQyn+9Pe/ET
mYsLXj/jF3C5Kms85P2fYA0mM0oPW6b+L/4ObLtnwiVmwL8ewTZAi9WZWi+sIV/c
/t0+yULKwOlcM7qkw8zCiH0JM8KqTe2rofsHQjlfbwl8cgXnKffNmD7FDUh/ceyS
+bsMT4Z1OB/i5vjvPQhVr2lLWYrqO0kv9gZHELYdFDfzOFEUfURt0wPNBgoffFkE
WUFHl8B24W/+UG9apYwBNrXS6Adkrj01isrTIwqGo0quLdYsEtsSXouBvUTvh2I/
NR9x4P1IRpQLebnMpnZ2/LtMJAnq6ra5/Gs49sBeWn5NAoS5SmZvME5kPV1U2Ean
qy84lFnbLsGlvzdZXZKHvASKVjIUYYiQG4uK1nrbA/1ughBHC/JTlpYkrbr/K4LU
pM0VqQDSZcdLBr5xfuQSYbdFceK2cjZJ5Go/oYJmmgjH5e2gvotwqTPvG6ggl8s9
xCA7qqtjGfEdxXlTF2UxuUNjXs4a9pDTogR+ueN2AAqRLHSP0AouXA81Qu4BWPsT
rn48hVZZ+L7wwRCNQWTieSaf4RTaGXJmccAVyANekruA9DSlg+tmnYA5FlsxNFN3
nyhiWRJe+vsu4YB7ZjqHrQ29iS3PzkSPPuYt7/VCCUQfR+T1XGODRX6sHSVTiQti
UygKHYAFkVOZK+0yHxyZRmXdW4VnNxkBZNN7UClPMeI6EOWA+0reDjOVVX8rB0Qu
j7WuS79P9+tNzFxasSpkS9XjBHgL/SP3uBPVMS1jCQQOkE3ekH69eQQT5BvnE09f
BqsvZ6a0cKrSsxhKqyWlNFudM8s8DBoGnNsPODwNCCz+KwcC6fJt0p0h88Qic/jF
3bKYBGdO68MQKc7a0d2xWiZ1RdOK6UWJhaCMsGW5HLnD3ErIYJHz9H9DLkIXXHHo
7aRwm2VofHU/jrw/dkPwkG+av5soF4KguGj3vlX+vvW7qIkSJehAoyrPH5KQGfvz
pESYCRJPn1uvgjUkeiXRT8L7CTI3fdUIZmHztt0MYzbSkk4i2Apv1qW0pUhg7mNM
Dscwdr9qk193ghzs/Zs2V9EkjIJ0g/OyN8SJHuQ6dmwX/gvY4HjzI25VDtymrpfz
peQBBrT33v0G84nEuHbIX5eD3v/hXs9T1nEliTBNh9cfbUoGt8qBLeFwBLppd4Qr
cniOvKF+/raLFZxbEVCCGVGLWIAT85SLNHccIhoMkNnuHzdOl1nOsoxe9hHZ3KgK
00UeCn5dsxW046gmEU8GjIsRck0H8ycRuiqs1xm6gr9OyXKRMdwO4DRi0csW10CX
65vMxQT/IyoA0ynhbgQm0u5QTmaCdRsomsPrF1BwxtiKPuF0JBuyBmiLxJ/a/1xD
9FjQLGKoO85idaBN2+J7cmQVnv77B0nL5aqvGnCZLqOfhrkpL5+UoCzGCgz0ywcd
3gLXppUhmlhUfmzfBokN3uqdvJlG2jw/EQ79fYS16dlsbOqEbiUf1prIN4HtOStf
HcH5+Yjnr+EVfDLw6ja6716L8L4rNIRF02qWzsUjcNcgAHhIawJaHe9L5jK9N4pe
orPBboJNsffw9WPRLQWTLCFmhu1u6e5vi3fgA2qEfEzwCyZlJQtRoS8XLIJwyPzT
HvaNE3gR7fUZKkPtdguKdn0gUnw3K4DLtxOxXXJW7dS+do3sfXLqfKyTlPOGQQlu
RlL9WmGxwkrqujMRYvdqd9c4wECX0+ORQsQyfgN3vEZv6oa9lr5ayxF8qmAUb6oM
JBG0RaOO8/FaccCN3al5IinBoSL5mQxsp09MWM3f0xM+qwutZVh6+VjCWR8SRhwU
hb3JHpLZ+d62KLzMjHMNC343X9+/D/2yjBQ9/9FVFR9RbGlDR+CNNf335p7hnzUQ
SFsMbVfhy0rDvPc0NLmkKam1VXb0kpBfkmNASdtBLPUThs95U+pya1RAyAdTQl5V
FfR3rGIqJg4OkwmRIoRZ7WHiTt9CZXvNHRuit40/nWWinkBoyLtcZny/UCmhtrE8
j0FRcN6ekg0l5mnFDWFLqF/Ucmj1bbA3gZbWJySBJkpnKQTNjugTXQZqXwnVJSWb
Mfx/9v9MZQ9G1O7MIm6JBamtJRkayfhycTy6ARzYxmLJbJpDTmXHCmxsWNMNKGu7
dW7q78eLFQPPG1rUL84N8hx0+oqH+lEsNjmDu+jVs8jqyoRVsK1Ax70T3LjxLO5k
5zmPJRqZEAmE1Zh8NezVXRXQljcyloRcGlssL5VKfqOrxq0svTGVnzGZ1TL4p3C8
u2ElqM9taHq01S9WIhK+yWV3S3lqheMzAXcjwYP0FhUamtu2dhoTveOCepFTLu3v
4EvWW0bJaH38378kmS1Xsb/4cynQ5ztXmTyBdPzcDP9GVNnrutfjiFWlxA5PweII
jVCSYg4nbf5bBRAeNTegal4NG2MJEvfYkumbN2ikz0s7agUaWX37WGneZDt/+BQf
FkHspHiIg2/V0l6ytaiInZO8xb/jwktuN3EvG5g+a8MFTOqNxUKc0fHPa+8e9p2+
NrrE4pxU7iNM9uZsMf/02hmr7AJOJbwrmBD7E0NGshINVp4UbPPTEzwiEZusxqAm
NTqdVUKV4167KX3jtr5Re0aQ+kLYeRc3zoTCi0wsSM33iw8IrozqmCJMEoY9OiSS
0MZwhFD9MkglIhvM9MSyaJtThyGd3O0ne5Mt4O60eLRgmoo8mmIkSFAZyXd/q9he
q1TmtdZx1iMs/lt/GFZ5+uNUm5/T+PpBHHV5RFUpQYjJh0al8wr8lT3bXkiBm7oh
/soX4BN0df8o76MpfEhPahl+zobhM4V7iNZHE9SSkvZFfpavws07fzqlq634SVX8
kvrf0LBYvouVAOrUGRsaLiT4e1uWkk4zbPiVUVN3hRzDnu+kOlr6ehyR30c7B9pU
WJUv8y1SdfJ5V/xisZs967sEX0kmI27rb6Z9VQoDelknPmMGeh1znVb5ETn29DIq
NvGRRHrvAwhRtryBYgnFg7rQQgSHEj0SmQgrT4sdYIdjXcpTdyPCFowW96bkFCA6
rGGk4rAlAXeF8jgSP27XJE/6nxHa5CJXjPeMMYoiE50qJEugI5smnFHxNjnX5+6b
kZExXT3bVEU3ANdBGwvtD5YwF6altcHeZILjL3t/opxPNWG41PznEXNzrlqsKJ8F
AIzy4EPpsfVw/VM75vSsNQikzcNOd3V3H5h7aLRkBpcFe8IRfjfkOnTh3C+2GBZw
iH1fJXpeM2YhU1AtCvdonNbp/XAPJ5XIkRavScS6Lp1ItDiuy43E67ADkfXxqtJT
qvsDt5UQBpa8WuA0bJmtiVxf+9k9Aw/9Kg6YmDSdHBnGRJe3JluNkrSJomJ+0K+k
AfKd0NwrKU3bbA8JLtDAtoWw8f75krVu4o4H69YdLpjZtMrYvTyaHvh7zsssPmdv
8dJjveSKgukqhxHDGyFFNWNvXjeH06D1CjVdBBDsATFBzkWhp5CE2RsQ+xYWW53z
qeXAD+6oE+XYipM2UWBa0Y1/HPYlY66ELetPExO2Z+kZety2YexD+XgynOsyO7gC
Fb+0ipCO+HLOOksV4MMysYLdGuBx1rq5h+B2ZT0SDmKURgb96R3nljkBBcKRBIzg
Z8gGBWB5ps/CWcXX1WKgWncOIvQ/MUS1mx4i+rFsKlpl/GroLzmaxUtVCLpcQb8S
t8MvQBRhYuLlwOmtMHjD0ma33Tg61Vyc3FtRY/U19hvirjKxN9SvaLgRsxiBa6wL
oWI3lwuLP6L7MxuWl0YogmGtjlGPAzTX/5qiD/Y/E2X90jmfOMF8iZORgdv1yNaP
t9IRV2LTK/DJjQzj6ctxW7FNLLN4DhQCMbebSe8gfy/5S0EnlRXmgyznUqfIKyV2
ZLc6Vyc5thQlQcxSxIrGJC9DvAAuR2fc2dX9bLxcWL0zm+cHlJb/i1r366X7MRJp
whl9E8WKwBYeWAN+FlqDDAdueEIhnFvM4GM4Ebsi+Uaj4mTUVqtEGsnDJzlj7YXM
C4mVH3uawqvC6OAqnV8NQMm4v+VDVnK9xOi6KKIllfEovoNQCse/FNFUyRrN/eer
K91YePVXjXccr+8GfpcHIhdVEaR2fkv95SHRVHQDMUha0U+X6aKtgqsEp16tOy2H
Hxi4AFEmhTYxDPBQUOZK26TiGITFX7Mak2/6HJYEAWepZ4DpakVOVWjOl4IBDvS6
GJ8rpcKNYFl4qN3nv4vy5fHXZ9PKHy5iwK2Do0CGpGX3k6sy2a8gpYqFFA4BfW6p
48bKBYLjzRtqwAv9UJPJ1IXH9QYlrGQydRA4cPQdD0knuJpKcIrsngPKZCs7xCBz
x8sU9oK1aEUcnyglUc2W62NDEOuG85p3q/gUl49euFFJLBlKlmjJleeITkaF6oKL
4y2BEPiHdzMCJ2WM6Ulue+tK7sGBRA+P5NGoYmoxj8jYBE5+UvjdmVI6NpVWuFLe
gfp00z5H1heEbgVLPjtYd3B65EQVLL809fEvoXXSJU3HB2xXPd25guTkMtQKCzSi
4G8/MJy0eUWeiKNbmFxAfm3jvoi/V6uD4mXx+aRszS6Fu2/qzCw5CEzSeR2Sa929
nHkslKD1CIaU67uFtzabujEdRxP8Z+AGhMIq016gRbc9FpfZiFQ8m5Qs9EpifTQr
1pjOjoCrkwuDeS+IbMRVl5va69COc12QhomyS7FeVYDduoenW1QxKrsVMKNFtw2j
N3HZ/Da5Ygva+B4lFCL1xJ8k1Qgbshox8cmZ325EkEP0p67nnej7/7kNP8SgnJe8
UZBLUSgkf97oMxkvC533AV+Ac4rVFLSf0C3Ztyq/SkCVBvejLbJjdXxBkEftScFz
wmnqEn1+3AljY7SX5n15io98/FjOM469KqRYr8Q7P6Aflr8m7xXKWtdndDf5DleB
4uuvLYcEgc7mHdfknakil/cuexhZl+GMlG/5cLUjPSI1IEDl79VN2ITSYIVPtPNl
x/6+rPqcM0v42Y6SGx7g9cviov9IDsHft4sK8DMsf0Z43jzRqe0+TrYZHxS0ZzKp
RcO6mrTZy41h19mKEzxWdneDedZDd6OhRDKGMH7P14Xrm8AdHhNh5zxQkMuH0yoH
AoJWpchplALOrY/S+92MD/uRmQzx0azmFQakrsbfsBel5bePzXEmYQHVHqjKcDbv
cjKb8TDNCWHk9vMVB1bp8shNYcU09/ML3+P7nH1NefuEYGkd793oLxTnjwZDQOoc
WxA5ameS5cidZyeS64+I0FYtw/eXUlpP46o0A9u8aSh5yY+pxfk2Lsh2cWJYGCjL
vy1RsI+S4FOhodUYKDzOcbj3YeyXMjOR9C1GsPadzoKK2lD4r/HT1MmsXFH2oTaB
dG0hyae/Zr03YYzuU+oOClXCSTZ0V8e8uDYji97NMsoCo2AEZd+o1VZbJaS6Xuy+
n7csVyCK5USjWRNL/NuoUWHX1zsFezrgNGAKVGc9sjsONqN7CzZ6lXiC49ABG2fn
rdgaU07coTkOdyZOxOBQF1LcYSAsHy353MrFqzv8KOQFwWrAX1TWsYWTnGpr2MMZ
4cqBo4I/e4vZCkhOm3RD8RFWsYDt8v/5haIZLnQIMmfrFdreajdKMu5Qv7+nhGZ8
JpdjvibYCwngQ9e4fWekVDlfcpB2qDGPtswyh5mj5R2gz6tRPhBqmV1CCuWMmpMS
5jF+Ygm5Hm5Nqyn1E8De0RA84gSnpl+aeSi6xzVguL0o2HtUn+B9uRE9/rFSxw3t
RKR/35Y0b/ZLtaEACDdodI9GlXb+7m72H2I1koMUHwgwCoSaknx4e/0ywRxa721p
FJ53wGekX7wZXnyI+4FoXsfibwOv06SqXQBGdwUMbR2XSrVbVbXatM44RiEVYXtE
vXTRKdJdk3rU9pCwNTX1Cq4KOZ559DifasOaG0sw0rgxkM+vz0bqYPYWrnZS7D1f
P5hzdrKY8WnhCZyl6e9nX0+nFjUjgIksoOZG5QJnPk07xAcfADinl/yaAfEjGIEa
wmDgCwGTaLxOI6+SHbLm9UM+KAllWMo/UKMe0Eco5OSgiLrTq+OmeVDX51PKcLMv
q47FljCxOAb0vL3ZvrnnRCfzwOCTUeUbwlpMl9JpyY2Sdn9MZ1HjMou/CGWJudW4
kFXspOyiOhty6GpiMzZEtrp8riMQFKDUzrXvWGKEDYp0cEF64opa2GBcoAzsLNpZ
lDhOf63MZ7fM9kUA0wSK3R7TMpOSp2DVRKar+zsj6HZAZeqQ0Iuw1R/joh3JgIPQ
WI0G1SsJI6nQMSxS4DXIOmPlj5eMnfW0CBgJI2WhM5Tiwn2a44iWmA4UIAd8c4Jh
aSwNzjoYhKCf00lopIuVkB5kiiTsTTVPGaeCbBiCZWCGn9JHA7nAF0C4tZYbEjLB
8yDXaw5XrAu8eyRPI5DUnGy9VQqx9SpcuVN7vmviIuJ2cty0YBNrj0TUFkQW9XkL
iylwVcp+RA08KBAPbrM9iczI2E8SMGRXnXG68uBEExh2epIakmXYXEQ/XzIm1fBp
+cZ5VBT/dTOSCU4PFrzk7B0PiloTzvjeZEXSKXKOysf+mAnSnarnJnIKtK4qF8ZE
U6J7C0PeyafG8PF76PzLIF5XPAfaVH15GwdpFIuC+L6zA8lyTWVYjqZk1TyCBqiw
3Fs4fj1O34AAgEvuiKrvbmzTEtCrsqWbLUZ7X1rEUCL76TmQU4cOaPMBmbDpLm1q
8WN7c/CCe6G37d9jAOzZQr2lL1dSbvwnes5oKVrLbtidgtU7Jt6bwzwGJnJK2LAl
EM/KUddZUiJ+zAt9O1ORZmBQUOc+DrGutUqO9+fR8xHE0pUkqxXaZDhm3qGwgu5E
rnfuyerD5mRhX3pIKTTCcsJSwqkTL0/ndZm0S4dhGudYmb1y0mprhHQ7y93ySc0I
ZJnjsyCTsVLiAYSNLIuqsChpTHZx4DIeYTtY3FHukF4i8LfhpmDTbd3QVcPZVLEC
eQ/uJSq74NA/yViVD4bzGEN23ooqHe0CepxHH05+MzqTFZgikpfbE9DIJNanPajv
1hACGBSH4CVs5x9q69x7JZqAuv6ExCaRrYSMJd55vXflk+U+RAaFs4G9au2B4pa2
J/biJDR2RPn9ZkYfBb67xrgfiIjfXMbyyhHeTY2OpqGgnfZHhIiD1cF6HWXQ43gW
1CxMibs0wz3LqxhU9mqkyPcku2rkc1csf6W8nTuZCPkIDiSTUBDTuhTm26GWauRc
Q6T6ym3IcQk6iEpasIolYyf/ym0XhVhRqUZKJT9K9C3Kei/iuB1nHxzqgB1R5oTF
IeWuWLwyfEd8dX6XxWTLyCcKLAqK101MXa5k9utJeWfnL/k21tWH5go8xPJVK6aB
OHLuFrb/MkCqFOsB1TJ8na9Mo9vaLgt3xB7BCzHJsnGseuWE1VWUf5qUkl1JqEZ9
hhZNS6ip0APirJ6A2slhyWxrMyGdnx4lUJ7tbbHzR0BKhWmXhWYI2Cbm4onw2Lak
HvzlUGbZ4HNuE+JJfavekBpc34wVEGN/xAhaOiz+i4WaT8VnAU7TE5CV5U8yf/24
uDZ469tRz5gALAKOe8rMhDnG9gdTlPJoXnbIWeDEO8vSPVf0UaxmO/D0LmQzJ1PX
7G0ezlF8ynIsQhcIHsCzVked4evsmnqgMj31P5Ueta+suXEZxihTLovWOR++IMfS
mg1hHWs+95gdj8SvaGPeuQyOuMYlJ+LtutIDVsKyGYKv8MmxsXPcQoetkPoYq1MT
uk7B6/EaPD+67b2iCA7/D2UTWqdwpPxuSGaTHOiujCN/ytiaC42hK0n/KXoYxq/E
AYG980g8vuhW31bS4veO+aCGRxyG346TJQJVwZ8XVSghJz8cBjoeGKy2frtCcHZ9
AZfVlnNYZc+Vpm5+e2C8VqQ8CDIN8w9FtMTCymMKqxOEyqOZbt612+2y1Kx+JUrs
dNl+5m7wFGG0gKkxvYsDiX9253PK8fUk8tqyfGxuFlpOgx9OzyZSuZf/oQtgnl+i
PFumq/mlqrR2d6US/o3FEVzUjNxuaRy/cv4KAbGkNiUdjid6abEh79DDjdVQaBQ0
SzqlS/9T8jLl587LK3/GaUle8Gfsh2IOBVLjTAUaQFxn/+kFA1c43om5pvZamJ88
a6OlUAlEzXELToGZTwqhdTtKHaNWG2cL8jH3UiEznw+k9YBToEKuve8JwZK/V2Y1
XNTvfRab8otvzzh+CN8jxpCgz1IwXRHnTcQ+U0e1C7TZ7ZoSy1eQtZFvNaD8zk4z
YdvrUwiwSgQKL93UjxUJDV3C2gb+UmsVP58wyROJewwCuBm6ngQh0iMmv+O4cUT2
91j8q0y9EnVOQT82u2GdGWZQfAYJ4S1qMW3aDKmaoE9X/qYWLZwDkAMBTwnUdVVK
5CS0NkiEo563BpgGKz7EtjpASM1gaJY8CGKa3lM+LGq0lHgpdJxS6Bb8Da/CGCtu
EZY1yw7Nq474DgvP9RqhFDzX1nz0V3h6dB7CPlmhUopg20OF8RLRbsDOErUeITQj
8yrUxabzbD7dvWnYuaes3b7I6+PBDxNJV89MNRxVHd9VbHXqxY4li27dq9JYjiIz
BBCaGWWl32+c22xwRkNSdzb7t/LTzFtCB2IdeS0OJ8D2nsU3JUj9DTpzlH9OEf0y
JDNdEVj8mzKr8bjkG3pR7iYhsb8cQW0xo+/Ts7cAYQiubVkzfrcDgmC47u67IXbb
wQxdHpzwWI3BSR4w30+cGUa4HfKVb1Cxc4MtIfCA4XeydOozzp1Y6+ezQOwkyhoc
0YaT/IvxMODu3xh+3Iv4yxvm5iXNJRHqzFHNUqJAmOg6X44vBA9DxMxkmv46Y2bW
GJ0Yzd3Y4bwCZRBeqDy55cXw4wazlaUZqWE9pVBqayFrpzQ7ns0wM0aPGA8WP7RB
kigjqXimbk9+cLGMaHdtkzbQBv5RPi2mQlJaVCLHUJk5fbJfZBfVuNx+F5Wh6ODO
tb7sygtV+K3pS5HX9KGVIVMxEPAoHuvwf16GMEfVIAc/kHfWabA07W1rL7GvLR/i
ZH7Zcibrle1X0jBFYHsZP35knaD3gDLIGCE11duh5nOlRst8WIYcdmgdAla1YzBz
rsB8FB6U5mEseo9veuznIvOazUPo3lEXO7nzqbjs5ksmg0KR0o6lvg8DTukWvnJJ
69I1ac0neWjbJaICtt/FkdtYMCgZO+hYK5a989jR9EvjoTzPVJlkUp+Zr+KG5mTv
D53tzf5ID6+ogecgrusrY+FPUHn+rCmajqbZ3aZ0CECGrD+SS8aRgb30nUAjw2jz
kl4jZ3X04xtuTG2dJ05rp1xZ3OZnZrF+C2HXOivH+j20p6FA48EOfW7qieuv8Npn
/dxLPpW8HE0RVLzuyJBQhg3B4Ez6eyY1ghb3ePp3IWqkN5JSLIT0Z0yBkBLLa/7h
dI73UbpOZoD7vLaDNe/h+cxuYPaYge+zfolbGyhNU07/Hqup5V6JmCvIagluXz/F
5SXnN7sTMLYqz+wOwrOgPpVDl6LaQKBu2JX4OVW2MWvYa4UEFGlyVYFCObQF+W/P
7VPRHVVMb9gjyR2ut7EfWROX50KucE3hBQ5ArbkDcE9vVdLBd7xMePlj4jMOjh1h
XMEUZ2vWm3BRURw501fGuMgCBpw1S+Ho03pyIij6WaLUg6Tb+pjCmehuhIdU2/li
ZQ4BTlqX7kk10xG90431tl0bk5f6yevg8HAwhqX3Sst2WN9AGUNOeb5fvATo79Wh
ULo5Ii3AHEUQ/G90EbDwewOLcFnxUBnQwXyq/5yltjRw/syqnq7kVxnN9ttPr8vF
XNjM3mIC7yLoYcFQPMHOJN7T9NbsSU9rJ2UrwCza6wfyLEnZUsrDT75q8+VGAsR9
G5PRrweyR80KRFH1Wm3In+0UTnhg68zLgrNwnO7GJb+HaSkmpHRydPmUoA6M7fHR
J+AwVp3eW1HajCy1LxxJNJWkjwhDKzDOQOZiknbZr4o/zwjuqW1KNs7+9Tm2MK/2
3+K281i31f+wkcXMrGdqlUquuUDCOuTmHzLH81HcZAH+ss+lzwAB6TaX2Nb6MSKz
b8YKrDWvYE/6GnjHUkNSBTyYDc9vfrRP3af8QAetSqnXKimydd+pHS1l0oAONaIS
pvstJ9VsCY0Uku6xBd/bBNOZh7pbVzWpNZyJzcVFnX8QctYCMKK+HOjGwYu8Zxue
vG2IPKexVZ1pe+9DLcKaeYutaF3KPzkbjwxe7LihsQoluFdLu2CLOtPapYumSgw8
c/vYahCYSY4Uy11p/id91PyU7uC6UFI/CXhsXQEIvR96cC5QtEWIED9dOnOLIcbM
mB2YLtsLDKdM+ovKUJLCCOJa3YVSxhGPDjgl+Dj8MqKjyM0HspGrbiJirYrEJw4F
NRp9c2tyVar+CW5+WRuzssGWoKQBseWDsiY2fmu/7Dr1Y16BAntPIXRLs9/mO3+A
ga0VIxoTXH3d8iE+yVKiUs7wHvn3uHLGIY4/bMUADND1cmncRBG+1lGr7LVcCG6e
8ZCwZGi4e+5tZzGnacKu05vsBdy3RUOAKeOXlO7lngqSjfQfz1oO6PwI+HeCB8Ud
XHijuvdjMEKEMpRTdLC4iSDukG4ZftoNO1Q/m8F7QVCkU/T4kxk/vZl409bpStL+
aQjOKIByIxEck4n2jk6CL4S1pX9/nk6P7+wHI54R7F91QhJjc7d3QTu0CAJ2A1rJ
Q0IeSpXcHUSnEa+3NWKvrLpd+oNKWIYZtNYhNXTruRmdA7n7WnDwScpgQzL+uyo+
BiQsiMPWmkvudnoJR6dgwj5U+6VDDdACXVxfBm4s+VyUDzCoV952ENSlrU0ZER8y
TSOYdK57nwMPkGQW237qWL6fIhSHGN/NRfUlce4RKgdqezXs5LIIVo1Pm6pxdr6w
YHK3UySkxyPULQGskI2bvOieSh2Jg/2M4szpE3dlDZ4LjY53KQSEOntxF9qRgr4P
4LtHQtEuqkfIZkyQ2e64FfbzcJeE0ZL1eiePArStvi/dUhaiGz0DSwV1UhgvImEL
g6JhN08hBDMUhl28noCgbGeVvQUraxqMm6q0jnACjtnkHGa8r3YeeyoN6B6Xxsuo
2aHI/gWM6ZJNI+we2nu82PUsmQgbmFggT3sc1+QtJKHgRjgGcZJTlnH9XITCRZWb
lvlfAWXh0qRdH1bNCGvDD6cjnxOpHjUVzQ5r/YVTkIhZpFQ7wT9hoB25qXlZGcOz
gCdVjr/U4ly14vi/pZPJ1zVzpGqz59VwxWk2Xh7kyN5nKnKFf90iPHKQyKfCzNGQ
vwv3AEEinXr9/p5rFPespBh15cfqeJXcv01lOJIKdczI/+ALYDi5uURWrDhCUzSn
+l7IZz/L5cEVBW9U1Zq0qB5S787v92OCTwOLXaevErz3rIAD9vhfj4Tbzi1h9nWo
Sb2m5IenM8ylJwZH0h+9fV5dWimG3CFNuXb/5Z0bMAv3wpzxHI56xiwxnJt74/A/
znl6Y5TW+LU/8B99ShLirb/H3T22KdcAQjvTPWmIaagSWzdgaDlh/e+ghMgkf/fP
IFKd6ifB+SL3FQjLzqHA3pv71jn6ZmMon2aqwLh9j21Q6T7db4KFkBiV2haNR0bL
prqZJds7P2gat/KF2oMIdGueDdfcDRWL6AQTTHe5bjWBP9hNoO7gtpZb/S1BMuob
Rj0i6NolWmHqTCLkMt3rHCUrHlUE9V1tZh9hQoZahTR3dFPdhifsXSs/qBVY3H9Y
47UjzwiYf9QvQog6/05/LRjQjUGHukWbjNZPU4jRe/o6kypGKVh2UfevjqSSKg1h
UjPvPb7IioPpbjAN/WpMC+AZVFFvybDUD8+GxZLyeYtzlK1THQ8TdIYTlPN26pHb
bU8dxiQYHbHu8NGI0A/zop4h1Jp6SRWv6IWGsjF0LURjrFIqQyxch9AfAcZ/amtB
xefg/fsv+oVRMjeJHvjI27/ucudglrDaleTZsFjPiBMpip04BPvnx4hA0bSH4kfp
SFxUQoiBLw74ekWNJg8BgsWe15x4wClcqzbzIOmxDs9RdCLDxNJGOGytW7E4MumE
nTmbdo8C9uXTD83JGYEy2bNrT2cbuh4ydgim0qJaJ74Pp0n1F5f6JN+bw88XGOh4
nM/letzkCosU7SuqXCRmRZx+3kv5ihSYVl3HxMD5Z7+WOCp/Dnbh1CG6ARkpTD/t
ClCmwO7zpxJ9//CUnCjwmEH2FIZsqAVttAbZapP0MRSZ0BaUqvraysp4N3FaKGon
0vjTRH0wIVb/zu2o6Ov8sS0Hmgiyns+1NTAIIA/sodsDaNwCwcYZutyWRqKtaRKg
yw6d63L0aFOsOlloraUUgNXVvBy7RZsVhKaJTZTJjsIQfaO7xTJyeRKIGYi4MSOc
/sFMUArL2SE0sFiUy6j5k329lCTSoP5NquSo+ws2qRNQUYTaQJAE+jh/KKDVF//0
s5kI/X5KZw//V/oGhiX7hZQQ4Rnr78lkHzr5FY/DTX6CsLvcq4RaLrs0yUHTnZez
dLV5kaY0gP4v4x8Gf1vmuTtkFbr4wFAlkhW59fUZ3IQTlzlFryPPBrB88bmBgSdS
ThGVhONqZJyL165c/XKU0YLYilP4DXWPB2YJ/5FrqnMhXOYL1XP0R5sOJEGMTjrK
16e0z5MZA2RJ8wIZV51bRvrtM5UCyrOYByt+oOzPgfBRQ4O3oKZtYfCNeI4J71LK
QUA0HrvQGLuSDZU7ADVBRD3CwS6fTA4wWAKn5XvkNsbpDE7jJsRBWTC5jeeL3cx+
d1i7noHMKQCNh3y69Ujr3QqtFDcKv9x2YdiWIW5dFvQSNXvud67glsTA0EL9ZyMr
kUs4k4NmWUBJgKpUnRdvU9zYHvt7le20yeS/bWu/jCUXio6xiAvvWmNsh9Rd1OKw
TmdZbpZyj1TKigdddhP5vFeso5JN5w/wJWijMX3QcikXW3/yZ2bTukuXgMFFieX9
Soe7SO/n1wIuux9evKxD6xQF48uy5wCgIjHfH5lPoSoDFoX7qWcYmpcVxc3w55hQ
AtK0xOrADdSiJQ9MGNyIdHU338CCeUcKV7DG3whJn2slSFhqflE8IkK2ckRmUtR0
TOoCjaPzociNjkXz/FOCKOcPoHgCLBHCv8HgQyldA8XVvHi6eu4yHv6jjwbfjLsH
lpNhA7IdLYiev6vMfDnvkHab5sc+KtXRElSIYrJzNmsxTxG32erWlR3pW7H1mXpC
AbdV2CquPIWeHzb/6KxKDZI/XrLsktGSHHqUwH7HVwfLWG5k1rMsuYaadD2eFsmq
a1Ew77giaTXJReJG09n4b+n9UvmW/oBip+Fy614aSDcCvKAeLePFDUpeKKgmwyLI
w2gaceQANSJ0Ia5txy0Kj1FGpFd/5opT+WBi8xO9j7taegMSrU0Q0T612vQrDrBb
SgjwEpbVevGcBSeZvxmoHamL/gauKZVfUcTAe790+MbcwXlmbFxnBG36q2Wgljqa
Txl7BH3HiZmE/UGGBiLpMVYL7zBULVG0qYsV05ptw0B7zyQeMkiv7ZMGCrDWCLI3
GeMXLeBfmSF9S4rKjJGaincSv2UDp6fF4zYvgSCl+Hfk3p4QolyTc+G1DLJxbcoX
7coe8zZxlUglyxWIQu68dBnKlb+sWRvA7OssWyAOvhA5XNtFHQWglS2PuUEo4n8M
DfprZ4CqIc/rOqrZ+SOdONeiwPw2Yk3X1C9gWQDwGyDj22cCDcs1YfIRThZT2p8O
YVRJTYoh+X3NHQAg7Z76vts5wD0DRhRBV0wEoZWR+AgzXPJA2x1wvDMJNQiyz+NY
h6Kf5YWyaNZsGUbNGzNOLm53nqYIfujCY/bDISS8KNjos+UY9mK4f0h+yerljDwy
krB/eNs42IEfBVuGrr4LH0VQKM/jKoDKmEiVJaCFiQ/g5RdbMvRk6VAJnn0rEVKN
Tp1h8GpnsDXaBfZQjmffyM0HwAOdUKCYWRV4/BO61yANn8zSb1XVk3O3mEr3iu+Q
jBVIM8yQaSfnsIZc+FHbpvaJ5yWA3tDaA2QFxB2r9c/Ad5IF7JYJaU/KH1GLLFx2
jn0Nyn96ZZHf5uYTAO81FdfXziSnXPdjDlNLs74lhnOVwvKAei4KrHGLNT+l1lXj
dPU440ee/V7dkJIZdL4D3tdYH5aU68gewfczEBO65PxEo/KIpfV5mx51TECZnqVa
O6QxfcPp9z4Iw1Ouiboc8/OnRo/MoJjzR9q9gzM2XUzmLsiZYKDEJ4kJnyeVkl2S
6SpyzISGaAV+WQFre7xa4iEeN+w4Nd5f8bWT/RxoE/3sx5piLEk9PZhkw6t7b2Lq
wx4MuLwfzMw8zyvNg1Ba5+HHqJgIwXo+/pqwaNhMG32xjm7R4kBrL/GlIxJEaSRK
v73wqubWNi/Xq4SRPhCd/ZXpwI6cZhqzxUNnUyWiuI1PEqSyfgqEl53q2WRYXEir
a1BZ1PAi3T3aMQ9m4o++f/zUNWJ37fzE9vT9bjRNDK65ypEh8HmZEJgcfExfkxRV
jJttvYMf9D/jrdlEtYfcyv/MH+Uxgg5eBtMXiHK/2boCsDLWmZJ5PwLP7+aKzA4q
BK47/7cPXeZ8UFJllVLexXU5SUO74Jrmov6uc7QdyJKHzpTR83JgwpTM9SUvyPhD
3ZfX5gv3yrJTv1IkfwhX690TAT6IFF6MCdh052qLpvU+kh3igW7wBRhfOWBTPHJF
9wk+rf03BDuCWcPqLQNlQXoGmjI2pZwhfh8tSegFm9knrfoPXui1PRgtM04bYBG5
UeQpyFC7/GDXj91oRY+yUx02sp1Gl276s/e44W7X4iuPrhhttVMy7iA52mUudSe8
iWF2Ri1JBu4rAUEiPDOGjKx8t6kF6xP6jwqA4IxIn4wiwezlROc5KOvZdt/bAsmB
nyBOZ7XXUv8x3jUmLFI7hnmmZkCq+x0hRGWkqO4HYXRlD7oSYV10iJKxgagJ3l/7
hPTerbcusbkXKQNbNs4rBidX/myyi7JWG4fNwQjx6QK1NgjAIrRBJNWjpMwuDoT9
2SnUvNcO9SGd1said13CmEmLg18JQwjInGrsWENvbPJfhDfnVA9KtkEhI9KE9ulD
+lbX0j258w28XCbgwYWv89w6Hn+wNkQVGBSzsd2xT3rWUx6pbYHXBtNllzlkwj4c
PO2dtejMMw+PGUK4e2ofFnIP26gJZkSeNpM4PfYv5OoW7eoWX+/VfmAnkmN+9Wln
B9kLF0IehE7nXrD6CYPKt6VbRvCw6avZOjcxeLDfjtOpj/6LPRZsWjdh4EpGtswE
PVi1qboFuXnQGJ/v7Ax989p+WmtBGUkHwfBBs2bgKjmdrFj78hkYmVN75A4Dg0dm
T8LTmwvTQLffvUaqNMuSmceSrtanBA33GDK80nd6EksOdPVF1TBONC+FFSXWvaaI
WK8BvN5uDvbXRedIBVskZxEHjTc9Q/jzojCXenTb9HNkaSusTIz9hsraa/pDR8On
+iwlkV5KfDreo5uHOtpE8bVFhHHsrDQY2CLj9aIUqadEWQJM48QoOx4KhGrcvfXw
7Wo00x07VMIlCKvxSdurzxmJ7tnhddLOFY9ypT60ZZZllWBT4KYxAozR8sL+xxlk
b0y07WRc9yJpJQb+4E557ZAK4rZaT6PzYQ9FbOZSK/KEwg6EL3Vu4bn4tyC89Ev7
ofS2KHYccI+5bcRZCOcV9r3pJgFY1A4oBettHLPy7dFucp5igjZjOPttIGp26RbP
jtF/U+ozoclp2bdjH4xnJlnoYpWhoXY7jbNPsxjIyNsAI9m/rFivN77iuWG9UE6d
H5sQEkZpHMbNivF+LiVL+O3ag1qwP51ELY2KYOI/ecuBUUdBDzGksFzWQL/otfQM
Mp2JTIOYWKDHJEFoBCIU67zwFdWLE3W/5c0PFXPhnQ4c1aNVXRW30O+UOSsfNo6T
dVx5ctnVSu/AcMFHYz5Lf2Rl+r9KlpapQRGKn/ymE8oO9fYUArJEMZN7u+XOKiPm
RVeVgBbGr6IJZVy9BmgTPPdsIHviKaw0qX9Ia/aE/TfYOXmSJKUB7CTEzKvHee2W
G4UU3bVd4AACbsTqFKK37f0YmdcDnSwX/RnNwtoWO8Wl7QxpeiaGRwlQ+Lrnepvs
xOU8Ob9Cs+4e+hiROwFbd4st2c4+CxTF/9j1XAUehIRqH6AnUm3v72s3z4iI1AYU
JfyIYT49Ijv3w030SiQLjWQfwSoAv3AO3VNerx84advphJlpyIt3JvWWq15RQbOJ
hbA2Z6zMUXSauYC7650W4/c4fmgQKu1PVhnVLIV9cyUw90M1cXBpz7+xfbTFGpjN
Jhvna8vJhDIatH8t195ZJ4ED4xfy3sn4x/RNtOJUXpU+jaYlcJVjD1zkdiL0q0Xl
OL2affxqb1cLw3sMf9stYYvGq7tlqmniiyUWU1PmoR0/MQxqalJ6wshimk5c6mrM
XaUNQw/A/wYWVR/hgOhY0kRcyta/BltgnpNDVNnf6rNoqKMTOh1vPVYOKPWHGxnF
94tUyko1JtDQH3jj6SuKAjY/r5do/i9j21h8F03GXxjcljIOsyrOokS6FiNJoK6/
p+9FbLJyVxTpYWrniaKflafHMTWSDJlG50yHnIBbmYBs+AO2MkbjytN7gCP3QmCw
WaN0uTIKS92RmbYhXkvRvgVBzvREAvWyMrYvcV/kZj/zNQgltMN1E3nvqsoB51q9
73eIEL3SOOKB2CLeeoxQc0s283MUB2kXWXGgecRgMZNKH/ZsY18ehscqylCsINSh
k1Yn1TKa5fqMpHaJlGj2gF+mhb9ezD1SYoPfOfOvjKkJncCfPfhe0J5yfBMO5x6r
W5qZJ1LT/GOfhzaGiU0NLaXjFbsPX0BP7IvMEq7prELPeIcN4sC6imDllXLbcNis
31sBStZJimT/fXWYAUYgTqIj0ll05XTw9AetpREkNj2o2zIp4drTIFX5XoIQx3ul
6EqcvYFKxqM7/4DIKiphtUY3RdzNc6DixkCXmWzk/pG4ZvutfnENJfYpTOynkgRh
2KkTvq9U8aGwZxOqkBdgvnHPvpT0CZPeKvKQ37YAaZCpqXiWMULcAP//caJAZnWQ
M0PFfJQPenbN0dekey6PbFEJ+A984bBUrbt6OXd2a+nBzKKXVpCp3iKkhyqDFqXK
uxKs8NG1nBO+vz/9H7mRih7bfh2yf7EJ/lEGRF+slcWJ1WhJMKbcVSNyDiejmr/i
5PE3rphg+NorUfdRtYB28llrQKtmMAWoIO7FTnBaW+5OQhJkW7Wb9NSLNy3gBzll
/RmsOEPRr3ywscEiq1fZCl9sDcvvdnAD63WbatW0hZ4WVRsD1rw+vsHga+wb+ikn
J/ldfOcj+6dyRpf/fYw/Qt6RloOhSGm/nE9rJU26Pxgq3ha4snBPe+Po7KsCd4Y2
41V0Qaf7riwQDdqNdd165uICVs8IO3Sst92AlKoIa2un6IlKmVSOkfKgLJJMv+Hh
s9tNU2BpNza1kK2dOfRV1gMotFyfgWN2nX739s+VyrsEHEvQ/AnH7VrFfkJhHl6h
gGJPWyKvtZItq53tfJCYLHbgxs10wg3EwRmDp0JYIkd1IkfYEBo7RjGgCbMVnXmz
2H6AIF8SHJdFYGI12GvaxoSVs2fmJ7O/yCcO3tc4YafAHNU9qoz360Z47UfTGO2O
BSDYo/EAt0fp4gU2yYzcpIrj5PkPOtQ7IeXnPE4zqIbWfwz9hGCYqul3KSqIHz8r
vhES8VV/xk1NsFjwA0WT/kKOBC5WbXf4tIXOzvGI4kXMJFeB0rF/CkJbx9uEM8bT
GjYyBmYgfuwoG2jwyocbRdFI7LQtxW4/xevn43/tGhcXPmzL7IPijDkksM8XENdV
IwPX62I48ipGsiU+5IZeljg508pIn2sbCF2T4/XM7mGwXFrF6Q+7ddTMLtLDeiq3
42DLN1425WLgVO3igTvorAGWuWsqIDzdw6AVfQ3Or4nmhlyZrT6U7yknTXjabEmA
o/zo4E6aVPTuVCYWkBSME7V5Tafgsm/Ft/SR+BzLaUXPljFyX4/bE2aH2CcJGS0G
gk6OSijD2QfF/yJqNC3LMQhIOOXkNc4XG+BgyJC8AM7bVi5Uawgac745vELfXaPP
TXDogiDINO+LnAzPcmLx05qxiBwsfg4cjHd0BNjT84Uu9rlxo5ArGfXeehLdELFm
CxYJVyAJIFcdWOmQSC8HrDtIUF2C7KL+1DkasYItWAR1KAzpIfGPm/agM5eYebCR
EuZzYNf/Itt1EZI3VWSaBgXHEk3ATXLzEKnCL4ZizoIWkhPKlRvKK7/HCwPZ8qMF
jcsPak/3BSHmKb9lycPeM2irQTeN0Pi/PaopLzf4c+gJSnhWwBEEx7lr43dFMkBR
61DNicFZnrq31rczVlfT+UVu1FOCCoVn0YjQNol1bL/rsWcMYpVdGr55poR758IX
Fn8Sburtn7tfbuumRGvRcuWOM04EvbDG76YD8Fyws2jtnOgsMLuCeAsZ5BeYUqNP
uCy6YhGlhotdxHGR5uNS23JYh6dF0c3hcjZv5dNuMbHUvWkVDpo5VVt7MPtNw992
ZEx109+Ed3ox1KLmNsgFyaLDxs52TX8Vtu+qRiXD+yQ0PwxZMIazcqYLz1ZVSJHb
22auTvxpRdjB1MiEtfq0xXTMU0G0mlJwsIzsQShkLJBGV8EWbQY7I0oVNVWmdTrR
FzZFqHAeSgdITh7B2kmjWfFzJzIEyngMzUzlgxwoys66fHm9Yynvas4deUBrZCcb
tYryLuL9nXTANwHPZhJh5OoVLrP2wKP8ZlVbSUQRL3KYYxccwcykftF8zkB+d7Az
SVaLREPZG19Ams6VCXtGgVwH5p+jxnPZp3nhbAyYsKYvgPRkiwV/21HfpKeT9Lsl
l+FpYzSfqGVmJxP/Pd3TBzfEsAMCHi91eAeEQYEEIefD0R1Q8BOMUXzT3IprJn1C
tHsLKBOT2itypbD4EfJ74nw9AOAbDx7MYA/Ld5zqIIT32/0H4zgSyVonFSqllQB6
lo0gFiTHV6kOwzA9+wMOId3KR4oDCQ0v1Joar7c1rQ1s9MIabma58SGxIilSph7Z
T69cRFDS5baFNzaPsFhrqrvHiNIzapGJDXieIH6r02If9pBZZt6XN1yKrJIKQ22s
/aqskQP9tk8rr8xonm789HdVo90sqKIVGCKeEfypRfYbT7bv5d6lZNRJSTqWLvOd
htUMHNSfJJHARU2+70pPavs3FmAKsYk9qOZEFVoHTSbcca2Gkx5N5NTcEnFGbrNp
8h7naNhcu66+jeX5pGYLWH90t2Lgw/57CLVhMPGvTOLHCdo7VA/NhYk4UM0j+C3K
DusodexWW0xfpjMNfBYuLX2uWaBGnhoLq3OPsYP0qwcPnlsCIPAlCaMJtIOXZ8MH
GhGLlbEWrC1klhLmJlMp2TPF+AjNzINxsIcml2/cPiFW61l6hWnkSqzHZphdbfcN
EUCuV86Oyoo9/9IHKG8FjA70D8J5qHy/SsV3/N5ElnYJeWmYzw/eNuiNhN3rGoey
F5z7iG7Ag81wPIW7gGDL1vjhEtF0RUG2QrjalvR78DQ7T5gTL6gA86tRGzDtGu4L
TKHrt0kBWgTYeLwzVBloaMFeRFCB9/vpTqk2g4F+o2Q6WGBI/j1xwx90xx6SmtdG
TsFizqaFvAv9vjTqy6ItmGu23+DFeQyXJwXP/kqn+UN8g74gBcNoHYBcwmOLQmjz
4EN7kh4Lz8ffJFcM63o77I9AFiuQuFKxNcXSdaoUBAgWuGbVvtDEBveq4I34+lA3
QiX3giUdXxT340Y0e95U24JLA2crNiyT/3DuoVON2dFOb8P5wcaYFEWAA36bJCf7
u3Lpqa67oghpbYMehAbj967ibl9vXP4UruuhFJPMbXPQRgH/Z97eSWefUNOKJt6c
ElYu4vi34oKFwJBtk2dEY0BhgC4F1QyhZuLIwFtow4bJQWXWkDc4HLu009MOpsuj
2fvCmba/OIp9UbTfAnmxWoFXzeQXJ4ZixHlcurjVE2o+4pFHL6a2YZGNxbMIBd4f
xFjxwJFgWA1WfDuoYdVYRzzpEYO1q5RYl0BfVMt+sJMnnzvXf2DSH2N9F0H7pJ9V
mMOf2/mcH6CO3iLIpPzzM9tWIRqd3oFyrkTcWTO3yi6xlXWcVRgxSD7umZCcwJE/
mpK8fdbFVJ/kjR1OTkg0F4NVFwa06NOUW8yDJg4pC+BDHaoOYjBs3pPeHsKpNqRP
D0nmxHGmA8ddmccpRsVN7qfrfYY4kv4+6t5RAILCQQEDHeGiw7wDUasBjdPbzS/O
qV361mmvJrYLojWzawiYBkQ6D4c3FkjCP+VlCBLR9GI11bAwdbEsdHr2YqOw44+p
HCarAjqiUHPFDtl6V0Y/NYg/Tw3Vl5GnYXFTSPZ7qRpj0p2wAK4DBW/taVcg8co4
p0LCXEoVaRk5jt8azt16lAFmdsx1YgAPsoHM3YF0yIQ/vTxRmWsPSk2Qh5gNycWi
B931yrSN/r7dticffoVN6WWQ8/p/00f1YOCTKkvPO5IY+nG827mwAXU+Ab40gRpj
q2jn7mVgcRv9vLITz0UVPegG56yH17uvBQJ/akOzEKVewHbzOjtoHFeEE1q+JHQs
Rsoz9QYrDyAEHhXHKQWiZm0D8mScOKjp/YPTp2BtyE0FF7jOw9VMqJ9bseWcedg6
zLesapWClsae/oFkf0Gl75HwncPNXBP0W1I0hel0wEhZT4nRuhfKdUAyeGKlpsCg
hBsSsU52oboOsGSfFsJivKh3vvrSKZ6xBeTzZewYbHuRKSmng9K2kXZZgMpTCj4X
eHOoSSgJPlATTS+A0zwPEqRPYJEoNXxBa/XRnt2K7Qxgik5CakfnWXB9QQePpxUB
mROuszrzQShJF7n4qL6In6H3vayzsbJ+c2YdogDw79B+JhsO+HbmV+G1x/v+8v3N
nXHhr68jWX86AbaieF9Nb/yQMtcesLTsQad+ld4H7txUHk1GL02mFdXiceGiCdUI
IMKaiG6xybSZEo5Jx3mZPUduN1IPN02tGDmHxaKOIF0=
`pragma protect end_protected
