// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:32 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Fx9LVy3NdMHc52uLMD9apHRv2AQWLPNTlhX3feJ/PjDcHValXR6kvKJ/XOFqTJ9r
lrNhRCEMEJBg0DeH11i87eSqrkTsRfMF4zelwmvyp7RHD71ZlqKdJ0XUEvXnIwT8
/AyVWmZCWuGkI47Mr8AxscNPr5pYxK5QJ+qIdgMUJhw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28224)
+zU++y6j1FZtegYOXllvYFkJQWuUrtKc6J1fbn28e+qbXwuYEGjKtMZtrw/Fe0DB
IoXyxqudYzEOL2voSx8W7/c9Gz9qeokPxqX3U3ppB4neu/V+6HN8GK689h3y+AUD
J/aSxXLKoshoJQu69DEFz1GN0CjMJAUez6JEopvOe87xiPoDhX5oABR5D2zasGjx
Rc+ltDaA65Spw/5J76crU0vx/7CjOKGgwLlqA4e7w1IqlIBIrvP8jERBAIhGSqjR
ZAwM4cKNIiKtlH+OnuMVaN6I4bCwjQRg4w46501RAfMucJ/x/V+yQ/FARSsQsdJU
Wlumu1lh1bh6+Hg/u+vT0G2Ec+XkRbNI6ahEa8e+kUd7YhImiHx0UzOPXk1gHXAY
XmNSnaGHht2oHFytZdQ1vvt2T6HLAq6Lds2fVWFONUQV6/iBLlshHLWGfL/6POOc
WTQZN+Uui2fVbNO9kzQpMUnEuvCQ7x7FKd43o3TDK0KMsNpgoidWO2YCftlC9MOT
5dTSvszOttigDuxmtj6dUCZySwpyZmGrAgHa0B6/KFhIZfVZs3J3JMlJP9TCsHLf
y7aNez+pLMXO7VqRFhg5ZmKb2Nmn9ofRCsikcDD178FsU3iCBzqJ+GZPZ9KvZ6Yv
aflOihaMn6QXkqo3kxBH4X51tLOy20dXX4U4o0BQGWSOaB/TuJnLyRbe3UebkzMr
3dgB7dC+iXzLFO2mWcUvbzPwpIb+rbamQ9W9Em6fWcQ+gCnA8uODWLZNrWO8jzO2
zEWYl3A4Obsg1wRo5ix/8GQKqKgaEY3Y6tyz54BNL1cthrM5IQhnyv9tNtARyhEc
FYUqM8EeU5vNir6WUgbIX9LkbWdkuaMND4ga94YcDzzMjiMuWWh3QHLm3z+pw+1k
s0xw7dR8wDEKDcoGNLMSx51Xb05Hve3xmz3xONeHskV9Nepk45IJ9zQunrgnQ8Vq
QsH4t1WDoglVXSsUjWUaICwQpmKiF6/sC8cV6kVdhGToTgcxXDI65eXrCaYPXDxu
JNM7tnd2pDOiVR5LGcMY2Vcgv3kdRiSfQU4qlc2oeVMO8ik6IFTqu83AFumUvh0o
olPOSXPH1kq0rkWK474MOMFUgXCAhJesDOjHZdOqeB5VQh5F7s8Hm3dFTVx5F5ja
mdEIcq+iPbZRw5hfT/8VCTQjW6EeGF9TJIt+wCCHl8f9+2LRzWTQZnYKRF8fyLSK
dsMTP9jZ7ZhMQv/j/vhuhNobaSz8f2DHOVWzd+2CLvCE2gGuGW3s/KBI9M3hgHmg
DdLOZI1EqAmL7jLMlxArnx/aXgLL/KOc0c4I4dSZS0apYkE7hbLKZWe8f64MW0ds
ARtCraoZfX2Mu7UTvRhvQhdWKxAZmA0GBmEQe6JXd3mfiqXc6Zev514YPjMWuuXI
zx+Ejp+pzPleKKOLZOvEij4DeMxByIBE9fqj+2Rls6li6Cv9KtIJKXpeHcxjkWoj
bJjcxbISZOisabMagjPsgoA4zdPndm/rV4/ZSC2VWo+eTn28Qrs1w68qZPhz6GGe
Rvwt6Pcwsj+K+2h7xY0UUbJdvXd4gNMgdhezgqN6uXgGs4H65uyz/BkB9MgkoUAb
qQq1uM7JKruyCJjow/+shEdKNKVKFEA0aO9PFd1DFnw34I1B/PBZ53UsWQF7TVkn
a2Bj1BTBJiFz2ft1gORaNNRFLGBeYUPpIh+tr1AciZC8+pXsiPFwJx1SWGiRTEUe
EH3zV3oSWAXUg3F6bz8kKkUY0ePlOLuJr0Wr9AknbdzP+TpJwlBzVB23tWhbpNoG
t7LITzJqDuKdBZxHwDvqwOrgg8Z0o5aDNiPVtJByBMamOyd5UIjm5V1fW/rq20Mi
qjRkmoabH/I9vHGojtTiR6BSjaMf9E6J8p/NxeN4fS56GbOfEgGCmghLQnDruet8
DzJyz7xnuA1YTKZjTxlfeCjxpa4WRHoqqUR5jCXf43Shv/f/5PbZ1X27vQOxes3M
oMuOpOcGhb6ShQx5vgtr24wgCrKbwT+h4A9oZpn3Y8wXoMi0JLZcsw2t75kpQG8t
L6XCAVA0MRFMq955AiBYZkQSWzcu5IxahifqoxHOlAAma0RhHmv0Npld9l0ws3Hg
wwkIufW6RRwaig7ZmDBJ7mk/l2u+YjkGXCxxE1HCeYXe5zIUfyQoCMnlkmlEmJCP
yqaZWBzoH3/M3JUow+1ZTWHeebR3aTu1VCR2VaLfT4ylCx+B4h/bs/+Ckk44Z/aj
0+Jjv4HhdmQoopxxIq24Dk8r3tndOXshi1cpFOqEvarQYcN+OyL/WOq6VLMYI2Cu
3Q4ExiUZDiZXltrUB9fINScnOWn87SgkMrodhdjT+ZOoRBLjy2CzK85J/eWTQTAN
avxBdkeqhWxdvru4iJspz1CN4++3HDRE67Rx42V1SOdEZwkT7DOTvqhN4NLILNHg
jYvDNiOspTG40RE+QkEcIXSl/0KJfwssG9Ts5DlVI0E5sL1709tjA2wNfEXOublN
jsaNVE0M2ui+hfI0snsHRRT3bmJS/FLvn8XfZ9W6HIa5TRWJlqt6aj6gbmG6Ux0h
S5AuaNGnKbNziPVS56ofY60kDiL9TNegmb2xrjXb8J7q9pNMxzHgO6e1c0WuUhBR
PtAvpmEBQ1QJFpH3h5n8IeNwiBuDug0F+XJVgNuiSt0qyYZXYt4c/pnenCB40uwG
z8j/wT+VaQky1OUDtLZ6rGSofFVzUdwSkwJgTxdz6T3PZ5pE9CPStetOlwdHUC+A
jgTrsNcykPAmG5VoZMhXiYm3UKLEV6gZnqgC/rerrQ+nMrsu7Sf7+iC4AeGoDEaA
fSCsUp+pGIyASDjeEvoEHuhMKPbXTEjgACAFXQOdXZmVpdtn4NSWPVWcdUR1f1rZ
zkiuvbLqQakg4p8f/RDjHaL8txglKOql5hL/QgeKSf1uBx9GarU9mxVX62vCE8Z/
oE6UUKWxhmN/0HK2lIS3UwOwivhRatBD4D41CrFVyAMUSQUdw6cATA6o6ER18/5Z
h7MS8tMJmuQMNCVVVqUzBFNEB4QJjYFosxjGBZ3/7e3UUFukmKP3gLjt/9Ez/h2W
zv8utHiGeISNfQ22sGmbeGkP8pEPu821td+rvbpQbbiUm90Z1ZXvgKuSa7HDeaVq
krc2WGvFm8JJElde3XXCuTu1hhxTO3c6LsWBfIrS4Ry2kejDv+0zFy8A3TDWesRe
YUvFrY+1EOYFrM1gj90zFDYDBk25ae5La9QP/K/eopw25TAqBdjQfx0+K2XQFZZ/
zUuGoUYDcLuFs1AuIylBuRMTYXtbCyQm++fsrRhtNRQLA3W0/kkOnoIUIm35Srz6
Wb3+qpguxSdCqNtahm+vNiYvVRdSy8O2yckxQpRuF0cNjf5M87C3GtfM7YbEzDEa
9UZuj5DBRz1PGbwMK3d/bKYXBrcHluAxmKUAizBLQmegapvduupEkYdqhGkmFdwg
EiuSfQjnh8wJrAeu3E/2NcAvIzuLssVAXXLBOpmO406Oru1FO+yCFYVhbZ9bMoWa
A/iH3mPe66Tq1kH/JYQ9Ydqu/27pffSSpw7voHV287Zyv2YoeCNwhWWof5iO2qgs
+kwXbhrv3nW438/QP5Dli4h50ZiL9XQ5jadmxcsoPR5suPWZHYD29vRSQhx4640U
wPYBZda1VPB+xNSreILHhG5UI8b6t6d9QsGKPLV3i2+sx4LkHBtuz5NpbU/dOtWV
LwRoYSUonZhTk32vP36PJCVzTpO1DgJamTxAEz6OpHf4EZ6kBKg9hkcLZ7LdQJa2
1vNzPGxglwtWDj1hEiQG3DI6ICj7NFl4xJey50vJggcVU3bkM5Yf8s8U1uxoHlOP
2ttRCcgRxMeY9gktqcANWSqueT1Pw9F672woGRzl8hXmC9RQ/vkGtOsnU47NdVfU
Kpib02m4fQv1l+UKQSg6mYnhmO9CGvqxe61QT/YZzJoM4eC3n4ihbaxLc6nHgx+X
id943BN6yg0y4HNWcchCkBesTrKpi4BOup6nXL8zCxKUce5mhHMfYyoSm2W+U8Rv
E8C0rdpva1CcE5vXGEtnt6Tj9HIMZ/FnRh1ag0jcg9UkhiiQIshZx6DXkww6gga7
W9BIZKsNV/su+fFvbTkhE3Y7WHe+s4atETnq1iR66+IV7fQe1ofz8iBicCMh5yZv
L7o7xnPgdNBtdWogi6YunpPWf/DnYN/PfPD0wARITozkkmIKgg6i6oXGBkHk1bkE
quzvlAEnJe9MNpfhQG2vZav4lQdvF0Zl1d56rj3OG8JDM5uhqJqbnZv7bIS0luOi
fEpuEmniXfsAVgf3//IcqcNTUHWHsH7MzhQdM/WfUCY5OnZq68NLYU1KYnOnp2bj
YxwNx7sP+vSQuCLMN9XXsLlEx6EaM4nOD8vtabtvJflutUh4ABq5zdyFts9N/FXS
fCyEP7apo62Y0wPWtyFJ0aSpf1DddtPgdsHJ5L88sZuYxzwEMfTVCEi1E2qQR5Vt
Am+jAkJNIulXWz1MeXNtwWpcCKu2EjSJd0ruxkc3IbqDafOPXiu93adQCiJXbf7O
bb1/sEnZyQhoRSs6N+FuZIH0HuaQ/jezuFxNHzpzUeKlJJeghu8SGgZ2ZQgPYoz9
zmtDleuv9PZbHkMe8NCgPSnFFqjx5czB5J5b77Qx+OG3VYHpQNvqwaMRnO9Glcxo
Cs/ffthMMpQOT0Rx9D4i5nW5rHZfqyxlfiNQH1SvNGdVYhwEMCzW81ROZBi7cbOw
uyKUMo2fzkooJLPTbs45t/1wQtich4MLA3b5o3w4+NJ5zd5aBQxPN/j3DKRhb2Ep
ZXGHkL+24NnOxQOmfH6IKJMj2LmdTR0bRxM8MVXRGxhAOsL8RI0j8lC4M4w0Q4Gn
xhF4s9Ny5Pn7LwaE2ZUHm+dXWdTn8+l7vLSBcfo4cA+Oib8KTuBesThEaLBj5vj7
8rvmZlYMbfdjXvGdo2/yodU6U6Lde1knIa9I+GNYXJ/90X24B63M7hfi2zpmRIX/
Pz4q9/whWlCzlKl5jMR7GelAJaX6KuCmvisENgkIfpLd1EU7rC8IigVfNLhuBZvx
2bxNi4q29vI7JsdEAN/TTP1QO4MGCFuWNdL68lv1Vx7ZZsKZuFnlt0iulEKS7z8V
18rEO67pqOWqom+B1aY8coq20bExrqGsjVxwgXv2ORdEyfPhAovYt09ms0LdCpYf
jkjESbcZ0ILQsbIsKhA0z30A958lgguhrSTX+wa2YQpnaooXXrKNRblZY057N8CE
Qne2DCSIAThevHOE8lfF9k04Zcay8I053kN8ivu8vLdR43QMHZvsOqJUlWOD2t4Y
sP9g0cCw5lCvuHZ0Kg3S13CtRQIWJsM1rEs32sjRYBqXR+hhBB413LEWjrCq/Ew+
mF6viJPrd70YeFhS2TqXr+I07gUKZyGTaOvJx/P9bYKPXmMJ5e66LNFY9AVae6NZ
0Zf0RNPxze+M/XAZBhfCaZmvBfqc0BXMg7IttWtCuwGfFXEgaSWAw/IT6haTTiys
WV8J0jKprbhvGco6lTUFRKk6AZHMmJWwTPfw7rnb5ZaHZrbYovwr6bL32WKxUnRq
sWFSv10G6FwGoZQQqoa02aXCACxbtVtr5JMaboyJz1lmkTatM8/zU8v93HYpIZ/D
TDPmQ7lnlUYtehmAIdclQvZ/IleON5MXS47Vh1qffRkZn/OqQSYNu/uIQ1UYAFLF
MZroYHzY61Bo623gM1n8QGvGZVb+xS2iXLTCizkfxTkGOFGZeG9XHJHcYTKkjn0Y
eUnEqKP8TimhOSi2fRP4RsjVzzLDQXCcFIQgA53r7lJJHpPiK5iC7lXRxu7AeTuK
eMS+XQLUWwU3H0rbWwVKjUrf4Bjb1Fbx2nU/jnhqawIzAlga5w9YLpGmIYZIbwxY
vP8oR9Ut2Gh9dy+MqsWti7KI79Nk2NKG4oME/zF3KZJ6i1VXZQ712yK+MZ1xtegM
HVy85jBvpOWOcZLiQ23kOQS5cMdrawt3iNdEbqfK5hKLmp7pCUXx8aVNaLx4jqHG
MCRxAAJykoKma1eyb1UagLEzOBDG4eAhEGaC2u1oIkGPU+yFlIRTmNQKraq8ZSQ4
nZ7j0xaJnc6gYG+32/HSLNOlk4eVrAfLvi0CGHLdJ6cP9X34+vuleLqzF11/2XaH
5aF2OPw9JdLRCEq3QRFPxksgh5+RZXOb8VCx7tc6OmBRcxixD0V2c+oIzAe5IYSY
WuydyF8LDWoLhhK27RInoD0yAL+eLfn9FQoX6PLKUaKrbX6w3j5rB8IBLTCgc7ee
W19VGhhOSmF+t9LvxAQ2huubhQAH/zrytaH8l6fuY/LTzXtibeH2Cj9Ibs2H+Pyn
xvh8cd3pAEJ8qqxdS4UVg4Mc2rm//uhERJbHEvJeBaFNNz38goxaF4yZ0Y6lviIy
SShcOwna+TT52bP+xVpfDmUcQHWceF/cVGWlFLZ79MykZ7zeXA9dWeRQPK8TffGG
YqZNM6Ih2r91Tk9NjDhiJFg7x4qPfIr4A6eZZn+etSfyNH2a2EV7ZuZHOKKYZCHv
fTCy33TJsvIYTlVlSSh+B2ajfqnBI/Al0P4CHihy7G3F23N28k+f9N8OmU4sfU1s
U6xukTK55cjxDoUHgRBKG23d5HtssBzMcbu25lFkn0OHZiogVIwV48bL/hZwXjCk
S1K9g/lWyUCzm0Qg7i0JtwYevH/ZM8TdTaf3Gp8j2pfxm2A3rdVRe8R0A65FdvRP
tmy6u7qVkUViMDZxTwh1s3p64+/gtN5ASqnK+ulofDxxY6hXd8LbBw51uM4TXPP9
v6R3JMgQeJltbUsJ0bCHN6eyLcb+hihTJKOQNcLPj/CjICXL0UZgVBe45uWY6rql
Lq6B1966DmF1Xr1U28SbDU3OrVnr4caZ3HJVMIDqi6b9CIFYuC8JalokEeUDVRSz
rMYDRNLDhR/XCBDXh5q1474s/pa62UyygOFqLiwDWU9394o4dYEZLHYy0JAxW1H9
Vvqo1+ReQIFN88jV0GWvfGmwk4UytQe9pf7pjGbQLEdpCUKp507EzMJKYQOHc/IS
VLh/34DxMuql9jNr/TdmCcueT2iHLfbC2qSWeE3wsAIokXcxK96lQshjOskQgQNn
tUAJNTtG/6PFANb5XCsMmvNxBM6YuNi15zGkBXWyeeyE8ZRi/84iGPnE2GVrit0B
E1pFWsiFO/49RR6RXJKMCQuy0hdnQDzvdbsZ7nflm7qhCxni8C0Q8366px3P67BU
uiWt8rFlxbCCrJrzhVUFmhqrhAIW/XC/F+5ChgF7zQJnebOabCK4TOrCgFEucmd5
yY3WaKIKy9Jp2VEkKN7z4c9u6Isfq+98ym9Vb4a3XJch+jNSDH9xrlGvIj8zkerG
bg2I8hAomGSSMG0rVqWnCFg6AUM8QaG6ik5B01ZTksIJulJxZKcvT9Rl6VXKiB/B
x6N7GNoFfhFb3SqA3f3NkCuRx4wQ1XgP4XTUjCxVNZC0BSNHldhCdpViEe+AESL/
hw4O87UgyXX3ZuQI1mJJJt4nCtvkEBgPHhTQxtn8ltUr5e7Lp3Jv0XVb4JUAmsi8
omEaZUDmEZy9EWdz8OPUZq7XpCPfm6xnrV0PiWDXazEezJ63/Nuby9maBdYhMZJh
8R/YdfuY4nem1lbwGZsAPOvvSd8Og1f3aH3rcuyQzHRU9eq7zFNlPDKEyKmrl1Kl
minEPLdTcQU/JdMbXPP6iV2MWHsxHSzJZWAtUraH5AVOcwkNHGqX1oe14mrSi32z
nxn/5qJ4OChERs6o7V+DFs3RUeqErpM17KWlY61EwR0fC678iwp6yAcIRJ8cWQYe
vNQkwapiVhsVVzqLxawfh3Jn4MXkCjhNoKZWQp0uA3FxfYF1GhUWpInMc1J7Bd8q
1dn3S9qlDbv9fhxvdkALzUIDURWZCtAuTmP7k/oV8MT1njdIa0OhChEYFB0UnofD
ECyu0J5bn81DC66EvT8XbQgBqHMXkNihzA7bu1ONGBAcJZ4zqj0rXRRQoRbvJ2IA
Bz5tGh80ewfKfHvjTVtc+5jBFGRRN8EqtOSbHyXCSEWUicSlOBTpzXj7AOtENxZv
8nNp1ZJfwiQxTAlc1XfZ1xCUWBBbCjpP5WEhlWu1SBHjny9LznFVLgew1h0q4zEK
7vUXlxXJbqkYHXwiNUoP2OdCpNtBk2Igkpny5FKZJ916Q2L97IwqifBgVmV07fDX
NBJlsvo7Y3bbIfOWHVrMT/3363UU2HhLTba3lUV2UOJ0b/qjAEchZLvr371L4gNW
vKzHkvV2xK1OdSzKCd4My1T0PP7jU5MteF6MqKygBHAR/EGhAWwMDGG8M0LRd1Rf
G1bsKQtA2MpzYKfMWkMNrYl7vNAiugQsxjLQ8qMZ2BEpzeXUzvB1eTPWp+NMNcve
wdvtSLIYHk+YWnM+b+NbFRJYyYn0gunEg/RD9ywQpAnLinNUWOPa5FqUcd837tpJ
1Ptr0uo69riM9PDLpaPkpcPbHjn7udrMYy+1r53xDGKgHyy3Vbh599Qq6+oq+woc
ZalN2hGcX2Pn6WxyvvTkEC6qSoRrHzHwab0P9ehUJqyOLKvXxnT58XJye3n1WdC8
OaG2jWDjBUal7LkBr+WlHxCKsIq8TyOGVRjL7Q1ZEFkpneXd5K0QUk8gSgFfaFCU
2LS5+HZELpqgmo/Bw3EpewkkOtUxTKrhc46AEMgEx5QluYPS633KD0NwpH8m1fuy
4dFYsD4a9POqgACUNVxHoMwOItB9QOXe4db+4FEXGGpaKv1noVSMm8bDZxDHUPi6
cwvDHhkY2PNiTz1wVNZqvb0usOK+tozfL1DzsTkMz1KMuYjk/+w1JG+gg7QQZYfs
zm6FnXIDZrM0VCqyybIn/QygfibcYaL8Ukg/H9XWNrCt7LggB5UYklx79wc9+2iO
tGXF7P7N0ctfaQ1+kmfsn4z5leaPXG5pgtCQ+kjK71QwChQTYQVZh0uQQTdlAja+
DFFFQsmOeeIx/4AH5ccKbQvO8dYsrQDoHcVfbbDk/n1anCNHlkn286VN4RSXup22
f5UuLbcZbH/t0d62xAy4c+xtNExMyKuLKZVwxZIukLMgOIpfZOm8wDfABL8WFdxM
9koC4u4raORXABw0UAqZt0Xz72RcVBIjOtk2y3KNaWrxM50q1n9X4YsF1/M4SbrX
9exYV0IeO1Lj0RvsgWdBn4vPP7kV5FyP8c8jq+juNDWZM9ESofPF5UUArWcv31Xh
DNyyFwwZxOUh9IdOQf6UcGg6GJgpIgeNIOSak01xUwzTf+lWCsZrKluhiXakRC95
jUkiXKPrzjiWjqMSbTVMSXrF2c6rIpU7Bip3gAX1WoWKp3qslpVX0SJvSRc9kmAF
rig7bV5G0rCOnEt8lOIMGvwnlgCjB7mnzEm7dKDP6/ZeZtopeYscjYvW3KSNmrCG
cz6VQgWot4CjXdyZtJoqiFVuGlGh9PMzcD6HSAUCQmyOYdmP4VC98yqDkBytxNqo
2Zge884EIe/x04PoSJzdAE0nBYij//VOVWkIEJXm76/0xfQORa0bXhzPifV1QP06
Qn5dsMCsIPo6PcXjDTqf1yUd2dJeyAQOJJS3udjyYHi0aFc6h3cdrutPUwgZO8ZG
wPIh9f65TTtkcYv14hfCT2Z9I8E/NdZB4QIEA9z7YB1KdQ6IBborAh04cZWE8Agm
3wHzqTZFN0GIjN8agw6ri8YR+Fi4fARR0Lp6stXFgZFYBs4MKMldCfveO9iedUeH
OPBYGtxyOByXF9I4qfZKIvChXdUvLmtcLrzkjUrJyDJlVrntEYJ0es2G3arJSwTp
4TT5jRwGNPgC0Ih8jLjof1h7O4DmHk1f+c6ylZuIVbnyNlePbLMnJt6tJpmO01iV
VVGq3yURzo6oBmRSpKBu8i9MK7ahX3peHM+CfN2ciZ/WquNsyjfWPOmZ7AO48wfk
LT8Gp0rqCIODHxEyx+FlqqIyf2sYknzjUYcY7EMF4ju/K4+3aejIHL1wd4XHynjz
OfRqZYZrNby4o7CWc/BnCe8W5s6VVa9l17iiRdB6d0U4MxNUR+e6UR1AM1DbZuDY
I+YhQnB4iysZZxkqBbk3SZJVumB3sZPGmGSyZHj1xOgiIH+whckbDmL3PKwH6cft
PvL6B6O7hnC+IMURUb7ls3OPchlN9ZcxS7WLiuDGxWTTKTBPTtqlOAXsMD6YGhvc
GbJR2mdWpVU07szVItqrxKBu2MFgrN9VNcWieUV1txYS8tV3MWywK3g+UEz2LN3V
sVoFoeu7wQvcPU+8Qlm8v08u+twSBuPSGXSuzQpXzyRBrmb9oeJOrOzYcRumVe92
URoZYR062JeV1vpb0xlQUCu198qXq/+oBSiFdTC5y5PfeHUU6KW5rS6ufP2DZ063
Si1yeO0YHORXiNNagdadwx4CYACu/WHMYS1mSWlzePl5phKX3eTcWR+nlMfDg6YS
eFzC/Ar6k2R4Xg3qCN+UR6SPiXB/KvywaYDSAuGFyaWKI1PgJkQp9X/U9bPULukg
bi+fQmbclE7yaUmaRT4+nyePHd2TyWJeEs8CSAy98AJ6Fou/cQPU2Ihc3DacbciV
TQqBbAsWBhY6LjFTRumsrocCXSNixrn0DOTXEFY/eW8cGatby5BciV1u3PooEnhn
OymFpGqanCxNWLD+fTft03nsh4RLfmrJNdpMKQSMgcXE3F3PYHZo8OkcKKXDXBri
nLzmjOmRtlSAScnOrRlIPk3fhtcJ+rl4kaTcH00o75dNxm+rj3Z4zhamNizk61DD
+uY3NeubEE7bov8/ADmkfDuRApSBW2PqW6FHYmqeOhYdT8f2hWHHqLudEJmuFx9t
HmzGriSmRUICS2UuIJ5QPQWbRXCAoxQBHGdb7V0gfLc7fcW8vxNrvR5ZURced8X/
VxWJzKA8Ye4VputO6vmgp+FFT7kAuJn8b/Ux8kdLZqxL/iJ5jEd73jOngD/fFQzy
BiqqAOUiMCsxDeTfcMz8o88QqlygSxmP3NZMY2neM/jCfrC+P2AWyn0goKJRzpW2
RyZyx3eKzIWBX0eB71/fQedJFHdvvrdomrqe84+uDNaHbYPd0lsO8QLX/MBRKd/d
QSLjtpy0hi+3k/4wXp7FVugxSjVY1x8dPFI0JB/IV+pDtkll2/LwrbLOr3KStvut
Langdw/JapNV7TGlxICUyMbEkZSyP/S/FrxJLwm/a+8igow6U6n4NzzcpOs2uztL
PurtYRO/g96bhVGt7R9L3aAVmEuLo0zZnC05cilUCiquQd8EPtQIncADu5uBlVau
nvxPXPVlWwe9CYyEuWrBPR975b7Q8ULnR72BbdJcL+HTilzAArqqSn2yVkC1LDPn
gQC+kxfmPugGiMWMdvgOsV64Rq3mTqmxPXoYbcmUrYcn+RRFlnoIDp2PrZ2ERNt3
Oizzqn70KU/s72RKZasPwxgHS35SdBUNMdSQ2Q+kF+UQ9J97cSHeMchtBJTrRcyH
KD/YWpxkG7zxwtCRNMC4wH3oZV0eWzBWAq1O6SVHj0nddTeaIxtXLqHqjYtA8fuu
j83dC/DeoiVkW0DKtKyrfQ8asEjVqg0Lxp/LTmcZTwYrd1JlrKzpu5RRBPUWO7nM
t0v5bhZB6wU+RnUwpRnYa+PuqxKR03Ed1OSJeWALEYjIunaW7G0NoT1Age9n5fWP
ubePL7A6qVUtjD+88Hwpx9//NFrMtTA60AxKapav9tWrAz07SlpnOSgCEtCLxwUe
8IiD8yAncYk6+yqIpRZvNFOm8WCxGh77r0It6kGiNVbu/61NJn7TaBgvz8162LaR
rO274Kh3lxYsEttoinLUA7wqcpEe6jP43N8KyNvT9Fi/SKU8gmNY7ojQBFicDB6C
OXtB0OeWWdNWRz2762UhMD8ZBjNnKvlnbOtV5nqOW0TOySITbMz94+vZscnMU2Gq
KLmbIQBQj+0i2PInE2P/Spu9Rnu6FtiqX1+nKSsWX4TZi1HkJ2C1vemnv4BOBF6D
KmzPmi86gXnPJdrIbBALCs78FnXR0hVdxUm+cr/DKdzePvKfPmnlhn14pO0NSn7D
/hsy6VqP5gn8RbnrirR9S7I4VwV3wgTFLCDxUJgHRtCBGnlEVtQZhD9XBk5Vu+CR
acRz5XPEBq/Z0aZHnp/LTWosxDDbrA4CDT+kkDQMEKCFp4WO2rdJpRHl/f2LJIwK
cgykuRGLGtXvxr77cPHM/AZg7diLwVudOYoEqSIwz/VrJKurReKG9qJ9Cl78XwSC
bXgx44gtNKv4hs++M8kub/ygQw8xXn5WH7NmhwsQ02/xMe7KzLrhjVfnIQYUAsTW
oDnFqsns/+f0FsspTZK6Y3WsK+2xbtOC0AjwX4bdJvRBXXrnvpg6/RufXF0nTBBi
vlnk+c3A7Sh52Jti4/2YSgxdO3HuQVe8lDumTz1p2Ygj5D8HXkWCbpZ8huvL71Z8
VcB+FKKjmv9Kw84CZwMJ3na+Xc3Y4xJ/9Yv28YA6JDpDG6Yt0c87EkYJrkwbbMiC
PcQLsbduvA/uH360FLZF7NyWEY4IqwwzvwY32shABuvef5Jwi7P6unaiHENzxeG/
lsKK60cFlVpd/pXolSLOf/ZIhbVNKPQdngtIq12jOIzCaCpSeFV0JMkXgAlzEeBM
kP8uqBPVGKIMCxHcViIhqWnHdBnzuFBoN8B7+bFtso+4UWjunEl8R4UeiQD+Jbh4
YUbRE0JbBueHXxlGPjueNCXW7b45gIgEILDc0SHuGv8ciJX4dKcxad4b08ikvQvG
Wp5H/KgMOto0/PE2w76Jv2L9JjPdtbQqkymGrbavcIuU03JiL6oMQKL6Q6ooKamB
/YcDg4okEZ0WOoz+t1UnHk4fj5J2+wtyMdYCEgSHxf1TeNEIWImbMRYv7v3v/YnU
AW3KK7pPD/ARqadJy40zBaxqiCxAggsxvfTYqKEnIfUwaMVNNqOuyaBTzxFahZop
bU+ue+0Apo26bJjaiC/oYHcs12UyYDakjlZVquz5hDjuu8Jmv6M6yYsx5uIPCypf
M5GmoHYC8uwYyOF3YpH7KijYe/hg9HXfK1zGuS1o3qewnZnMBL+JhSIRvwNvzUO0
txNMc6Q7erz2c3Bdg8u+pIK2vuv6oUhM7TQ/4c9rF7EA6REc5VctFeRzsLCZJdL4
ssc07gp7IeLze6Ixyay+v/KVyN20ytIi9hjU8J0uybo9QJnw4JAGrJYmbFopeQJQ
Yc6HN/UagcI4Ye4zE/pklUlcV4k/DPz/quKDpMuYeIsY0mWFpdDbCS2UGYcSqGH2
Pc+N5NHqMOKu4UUI2GzIuVPe40P6HZBfenVM1j6YlFX16adMoNUausG48KTx/viv
1tQCNoSMiYNpxKTZfJECtLp9FI8JwF7WDGjomGrKWVF+dKTxJqsujCwdjTbJfSYY
kDWzh9IKDxwAgKOoGeYO8bVjitsK7dSpiG8sMmhw1WJ8csR8pYt7kUe+KeqZmteu
HFVyBzqmazJM4OQunyIeYjbn61suLsJ1eIETFyU6S8EzI6RTq+jy9IEFF1qf0mR1
7AcpH4BFMU4cF4ecSx88FjYjp8CSj1TzmxPq1QyOXYqQFJsQB0U2REG/jdfrW1w3
Nl6NKKnvjEtq7svUu+SyxQtuthSmSegNFi8lQKFTI0jW8igp/lex47G8UqfTSVPW
P7OsyevNYJSrIx3N0jAi2hs19rTD1uQXlFCTMxQmcwB+XZZL5IQ0iufMT6B3CgPM
H5+DlPzTKWmZrpJHN0oMhVPA3zhu24iEmGKjbbAv3K0f8ZmpkaJVhHvsF9UAWsfC
dgftzOcHjqJMK5kwaDYV8atFnK1V8JonSt/DkJgNFRaJA9XhX0QeOxt8krvAHwaw
xVtd2Xp9ZbNL42gefniuTgfSuwapWD7Ob6Tk5MTsgskVwQZJ8FGhFdyMKbjFVqKq
KKB4U7txdu3fRZxkltd0z3y4wQ1701o1flxwauAD8D2E1ev3ooE5IhqyLaHkejxD
2PxYJYNgkTiiRM5yYYQ+o0TwxSgn3ivFjb1+ftR6HQtk7P8QThM1JA10XCHlPNfj
p9JNGbHK9fozZH9AKyT9jCNO9B3nfffoXvMHpLaSreSh2qKU0+KAsovOqui8yPVr
A0Y+DK2mRecT4H35eWk+CKueVN4XqbFtDY0EkcBD3lt4wgh1PVtApTo4dIyV0gvP
sN12jvalOxJBhDSLZRqm4nK4zCW1KK8YRpNU6bfaV8DLWKA8J5/T1wGUzRAIx9ZF
K85loMYXxV6X98iOsw62NTYtaZtdem2ZBzlqzPXRA0tNeMq5GRv1eJP1XASDXY8k
L+KHothTDu78T924vAli562rCEApF2dtpotJOJZaZtIJ1SlDcx+igPwR9JY7JNTL
apjUdmCS8b14zZGTxh2/nmZoo9xHZ3LXGPGrCBgp+umGSiF+H4ftwiRP+eNSHx4j
hh7eiyYB3kyfJQX2funj5+PqBgPrz5skT1r+dPs0uKNNqO+aYgqywPxxqnJ5pYKf
vef+Bjmoofs4FvJR4vb+D4w0UdDy16y8cHWhcJYsu8BXMArTdqis4DygoTDsItc8
xbj7sb4h7e5LhexoIP658/eOiuQ0OLhEfcBUNBEY4YuWXk2Dx+D5noAhXpsJLKTx
7H4MwG92BQvw7gjyyLL8QvUux8DtfTBgU89SAP3J6vZ2x006BB3+HDg4xUQdyQmd
lhB+QC/QW2oZaqb2K6xc770lDRZvAbawF9B9PIQIUwoEIQPLZOr5nm30A18gHWeN
weY4DZ+EAz+TCHvhIPLeeL2wppk6Cil6HC5l7ZrhZjazPqI1ltUovH4I49h6tmGT
yFYoRGk2MAnK+Y+GddJwBYFooHl/CHiJHZORYiedd4OWFWC4Eer2LIdPsJIT9f3d
NVi515c4fJB+lPtgsbRtY9KiKYae/BpLdnTybfLx0VmNohvVqOQRNFWOXOs+DJ7S
UO8n8mCZX8Bf+cMDUE7LEHN9qUjUletevnfL+w/Y4AdKvLkaIQ7lGNn6cRRoFr6J
w083Re+nP43U6UlE0xZRuhcds8Q1LeAp8iZhfZ7D57ZKmPtu/hi7h19RhtTH1cSv
45kHtAb+12QoY91YkZkMQ1FcBiYihaLjoebyh6vsMLaEUcVKZTJtnAaCwhwIchoT
wV1LSpETe2gq4Gb2ZsdgkqUJvyljcQ6x5msCFDjILgrmh+kzYehNY1jhdr3eGN6x
LqlxkLPECDxqrW7JvqnWYExGlF8eXJAgzR4YHcMR+EpbaARmxcQMsMQ4lc3g2iKq
firCZtt0SpabLeYFfy1Bez3u/kBVX6vi7Z2ZUFUR3BfA7lhaA1XiNuawWwedoPIl
Kw/k+iMpELt2oPStB1e95XgLVcncinvno3d4sGNPPwMuuEWzeyuvRTeYD18MXPgc
NZDOa7mD5Obko1MvnGPaQaQEaNYDTRBZJywAXR5bH7zTEL5J+fslWFe6Y3nU1/Om
STnHnwXHoaEJgCCubAU0JqAgdpdSp5i74s/9xK0EzuX01JCRII2aqgWWL43Z6zjC
LiiEl1wV/tzuDF8l7eCB55kxi14fVx6HRuDN9+O6N/7leI+ibLKPKVnrnnZbVfHa
NQ46NtEysukZEUtYgTM5Gj0LyHYgzH42um230XYfe/E7qIav/YmBhO2AoepRarap
JuEw5L3NW9P4R2SDjkwbpD5xVyMRtvyQVLSTt4xwUlU3OK+KmSIkcvGMkNtComcY
o1nhdMb5tqrQtvizeDboNO6nrj+kXsZbXDuBdXiEtEuNG4LtoUxqRZQPSt+QL+mP
V/nDyeAh2RWKmDUHWekW8vDna1smDjefVHN/tLD1KsQ90sayeiPEscaCWM58drWT
HxU9hOYbd0hAzIuMlXbhH1PrTOtnantI25rH2+w4ss39B5Rcev2L4n1+3V+9+pl8
CEUoLwM43eJFUOPnKilj1tGZNlZlig6M3zro7qlYsE8AA68njxCaAH+wYGK+8IBd
ytGLFKSgB/ofalFy84D19GhjNW5nUHnSQAcg+gpFJMm3Il3gZXFXR7ABiKVv69jB
1NEi3KGfffwdpapLj3X0o4FMjl5rki7cvQa2EiP/nd1FPTnv6XFyMIDXQHtb0xOa
hIk2CjmmIgYnZB6KaAB91CwM4VEh9xLBd4dmyQyVYOIUri3XHdQ3peL8YRFbHuLS
0g1+v8TiITIF8UxoJuYmB44/iSnFif3MVxkDHfA28cct0cZYAwQaFKG6nDC1djXu
88aSWPJhEV1Elvvz0Z7F2YKVID+ynf57WmMRxRiEd9Vi/0fUMtHMyxoYKh7uOk+8
Hef1B3T9F76HtAQojazLWdEF2Wz+RMf7irxQWIqvFjs9uFJgnt1a3cbz4bhAAfza
sU6vf44zHntgkEpxSXxHKoggJ/TSjbqJxYvMYoqC8RI1kA056laUlLSJS+8FobCb
GKVe3KVCM17HzUeGCogFKVaI9Qt9unDmfTsEvPi/WUmVap/FtpLU2itm6tqP1x5f
cTJityV86PMMmxWBSwj77hMdrLsm6UgjkjoSDs0yAwIUd61v3RZq9aOZsEl9nABC
kZL89QX47pui3Zi+usuQMFH0E1pAb8Si6p+Tl9ScuhMpc03qPU0/9FeFS1CDlMaK
HFeuOrjuRHd52hsNwl2+ZCUaeX23C+GwdtuNuTV+6SlZaGWhRrp3C5xlVTeGHUrE
3QBPSb4QbNUFdmAlDUilrog/A22rdq9DEfvPShJ9PL2XBG66JBojl0c6ha9JsdL6
jHqN9/kdyxUkTqlRTNDW3FkiIEUr0nq1zXiiqJqx0AStqUysz2UiL/tTOODgNakP
NYNTL5Y9BpQwZtN+3z9XvkUst+RoIpjEp98aH+K8YjGMtJAda+8pYGeK3GSd/iZl
a1zuVYmpUi0HcYSpvV2WLpArCMNOv6WI9wLs7DIjgkKS9ydVYOfguwAMwFDN9Bls
CXels+3Tsh3P9skVF/GzoxrsAqhizsBHSLbqjXiF9M5GCN7oWAzDw6CCqYJp7tz6
9ZAy3Qs6jIYCpmTZj+/sWMyHd+y/p9I8HGMp8UJPV7fj4Hgw2PxQLN13XW+7GoyU
DCWNYA4oQ4FCr7ZZmLUYoejwjrtEB8S5fRo2xwxMstdayR8jvhQy5bo1jR2EoL6X
H7ICSVtdh/WGeLkBkqFq/x0jYdWtk80w7Hl7EGk+VdndsRD2qb7WP9cL7CwLSLV/
X6P4TJC0F4H+nUqFUbi9QlFH1tgO/3R1tOFQuOU192FUYuf7AAjwuZ2LLHLruYVJ
Ud0oCljj0NQI96P4bo53Cl+APcBYJpmFGPDHF5h4IUi7a9zkVyLFqJTnWVszOUGC
0/Aa3fPt+8LOMNfyqhYutCqSgFCiF/3EdZMtDWKykUhQzw1MR+FqwKfz9jcmAwTt
2+YAhUgNSpT0Kd84C9zxgLorpdegr9j2TQU6bPeq54afNBa6LgIfqttM7g425UQI
iWwKThAMc55Guar06AoNIVWiBuYenPtZ1sRyFDUSbiiQOaVFTV5xZyx/fOmjQlO9
gS/e8rewccCCBl8MME5qoGpCq6np8JjifGZizWOLtPZXCe1DPVQFf34c/T9CoDT0
esRm6TFY5iNWE8YIxSxINIq0PJwmgyj7jPXNf8XdUoYYPOZJ3KkpvG0JlPzf1iTh
BEdNjUlpgu4EsZQhBb2bvpPQcgSmETMO8XCcu4l1/3cu7o0A80O21I3xy7pSroOG
GDgeG9N0eiNJI9c6xQPF7Qx5CBo+z+Hcw8BfxyxlMsRUI27uEajonrJpMjKKYeg4
bJoLuf0xnaODueo5fuXDHQm43nxjVLiMgmQieMti3MXQkhLJkQKO7fUcb5MCIDPv
WiGG4TsloiEiHQ0wf839LdYbIDndMYnm0mt8wBWMsTO02plAp7pDRg4TRqUX4gr9
02XlIv+FrufAe/oRnYaRyk+WlfjPtc9WUGLPUrPbCzl0LeXimbZu1yVGMNHVdxw8
S6ds1KvW3b/vxoJ59Sraipl1fsDq/25BQb418AYjDax0cv1jtpgkz4a+/j2nVp9+
uGaU9CkeDzk992kqbHXDvpGzjqhLCdIoikpAI1RQPSadp3p14CYhls5FiYZfANWJ
fWPAzZwpLKLSQDksOM3YaWpdbcyw36StR3hZeT4YOyoZqJzs31XQXCN7Y+pqMTYD
KB01RtlbvcEEQGE0W12ZA+Aw6h5cgOr+zifMzoZZ8kZYX1vF/n0TryfEv6AD02e6
nyKpaJIJxdxWoHoQNTQ8z97zxzLztetHWrqdKZ9tFsjGctpMm8DgJscPtOa0/O0L
qqkik4nmbTu/AsfDQ76jduZhNR6J3c9rvl1LuXMpEEpQgN9/CL4A0liOIIYdRDg/
4fIqBMFXK7LNv3PiydXrhaO5dJcBjZ6WBr4HGWRLl7H4MWFZTp6VUBmG8+kDnvGf
3lEkdvvhJ+iZ/nepahdrirKC5wqbFCNgdHgx8Z3Yug56ki+JXgjGLr1g9LIAcDsg
iIspkTw+uIGPd+JwrxrcggDWEI+jGLcmdIoUIdKVYS4avjxLI31yp04oGFnjg9HD
yvCuEW2pJyHZTKVYW8Fv4+hMyH8bGZ0HyW0iXCmoutwfcKrmGlLXBmytbNjIBBLi
PCN7h7ZH7GyHBaC0LP5nDnAwKCgCGF/J5EBfENoUc/QdS3qOZaLobzXi0AMbV8cs
Z5X/pXRZTnC5J0+scYQZf5wRCOXONTkkj7QBScMXRkMqEDrI7vrtd6xmN7K/lqN+
rEJo+aXY1snzBYUYmubiUX7tyK5f0EixSDUspIIjFoPNxNbNzpTLOHPwlrC7wWzy
aC5dxXxbJXQ1ihGiqGrnv1PTnTgPfc6TpyVMpZ+x3F4s/egv8gIp2jXSPaD/3R4Z
lQeMzKBGzxsOrDL75gaELTP7qEW6buUkzatBZqVnzCyMq0pfPBKqx9S85oQ7+UPe
Vx06DprMw2Tz3IpZIwPOPmL2NffmeIy1h0sqELQ6zKftKBfXSspZDqrwu3Z5eCrn
vQsxKvo1kfGKg+6ezZiQBKFCNU1ZheY/dCjXbGvpxDvJuMbXWPi7sLC1LScCgFSW
NI9+iWASTgdjAPbbtPEwFQ898nIV79Sx9vuZVpqtqn93iAzmPMfWaeIvSJDaHvdE
sXHNkWpCXuoxXDo6yVgyr9yXIiHdpE6koP1FWnsgCXgX39mHktfiMq6PlopFdNWM
ID3j3vOQgQitMEKs/IgqXQ1wR1opjvgPi6FQTDh2J2jNQzZm9284aqHz6TPBe9yV
kabCoocZMeyfRjstCZkq9ckAM1R0XX89Zlw4SI0FKuc92ASf2BiP05dR8NWkD1AZ
5jusfTdQQTJqa+2h07p1HirDyVP0uL1FKOQKuZXp1ZFtdoM6XSL65yp0rkOpLcz2
Ipwa70R8BlgXcaCMrja5BILxw1TZl3dok4VlB2x9uWH9Hw4SZfdMib7CDRMWPBi+
Uvo4EioD24Nz4txFVoRN9jOkZwMAibtCw7/430AgW5gSOOXG5tR9m2MaY9Q20gDv
W/7BjXykRyuOgRccDNzHR4rcoKEH9Yi29rH2Zv8WJ26WIn9tXQgT70dnJDjTzsaO
WbXGfn4Z4WbIKcWJzcPe+6EzjWv/UN1PnXvCmTZOyywqMd5G6y3QZs7WmTuh44qZ
2f3s6mZR3+4IwtdhmWW8UuBcy5gceUGZLrs5il3zIc5N3NbpHOHdz0y28Li8WyoY
+k02G7lVjivFZU+JyynOzd9jsC/DbIWXRO/N+09BaeDVEOamVKypBd2hjHIe6PXT
w0UtGs2IwsliWXpM5F6lREFYpN7zGAAbKXaoXH0qDtQHtCxnpK01Ts0MnrhTsuSQ
IdkQVobzjg9MlLoYI0yycnHgBl0bh6Pwhxl3Up2uBFh+oLeYl4bSeOvFw5xd6d10
VGPRq/KrTgeLQfRbtaVhzy7DPim3lQaU6anJu6nyVjvYj7H16gbpJEFlXel5Oqwm
dnln6EdWyIfqjTSVpBhmFooE90b3Cn9Wh5AjdFgYhxWDAxK9CqmHYuL5t7695W1r
3SKP3Oatn/1JPHKwSxtrZnv/zGV5F8ZLJQkBy0dq2fpkq3LsbavCLtH8di09YsxC
Q/0gCqZU0ThZP/4OmWq0mx/gNHQIU7Vrfanrtxb81J1QpG5UufNs1oCMEutgGm9i
XDgYlIQvxCYsXYObnKsNqtLyeK3P6rwh9MZt3K5HoV9qH8jyGHDAVGHtLpRMfmPt
h2UQuwwiUyndvu4KZSFs3Wtr0ptbMY6kGfAMPUDwZm93v5TefOgOe4vRZpkim+Bo
ZtqTmslEa428kxUtu/dAUK33y2zm8ho1Vu/HGya3No/qyC467kjXJbmwh2wtYjoN
xxwoxDRp8IODsQpF0cGEmseNPz8cFLi1KzJqpWuGnNvxda28pv3lmPVzMVhO0w59
t/P8WDrHJHF8V58MHHKPoNtGOEzu9e+ZmFLPQXSZlN7fBUkjpbGaDhHRLvVIYKc9
4cN1Jwg9s7GpgoJfJQRNZOwdFO+ucsHORpcU8p4tGrz1JxDvJGtl7cNGRheAbM55
d4me9gz5EHQETWQDRjr1k0WXniI+8Kk2eFXqqblapej6S+BNDPG4SWJUMsPQsE+A
V4jA3JcRzj8+Enf+12VY0C8YFRTscZaxqyFu7kAEO8CwX6n5SzQMKXwZVuls2H/g
WN9+sC32IYcSCE8GP/LCpQIfB2k9YPTbdFvQ4JcpkmIz8mbpmUOVUqyyxB3QLZiP
ABgbXdO8KeFSm0YpkF89lbei9vDS/PSHqo7hFng/zjVc9IjnYHS5Mcnh6tmGtRH9
5fRpLePa7Ix61jAfW0meUGkqIDwHoifYqCISA00cCgvpo16htZEuR/V7NSUe1Vm2
kmWbVJc2VAlYlaC7M7pwDkBGVpcTeHvxz5U9E48JGm/wnL3JWESjePMc15iLzWgt
t3D1ecHWAFY4bM24I3ZUT3Wj1+7ZtjouVhwV6RiwAvgDI6SeZA+691AIHqBwB60f
aIk4OJ+8MU5c0xIp6jqVoJp24QDSzHjCG/9twdpBgy4uLTfg6exAvI2FXaeA9ORe
zEm0KWyV3kHQFibyFraCXH8k7Tla+vSTHJBfue3FhTiWjoxYhV5BxohWgtmNIu4Y
+VnWtKFEDkmSUZbtH1gnNIC8T7zp92IIgcPZmBOEux7jO6K5wiWfLONkFOlieCcW
U/qP6+U6PxVOxIuPmBenEgW41KOFfyyOz69RcBBJrTzJLOG2YZ7ZCrcQAtLjoQfB
zCvaQmKCKmMUrbtUXjKRali4le390d8NbUM/VW29w7MBRbXgm/bkvmnT5fQ3lTqH
IEbbYNk+AkNpYD2a+LN3EPnNmW9NyZ1YXaB39SEnk6pxkjtgZPKb9iKPCYsrooE4
fxuLNbfFppDoVsqUIneH7CpCKYw2/1hH6PaLq9qihU+VBGwYtk0ZwxEcs+ldjzHk
nk6iM4cwLfDxYl5XI50HC7JAcqmdiZg9S2XuHvoMEYVAro9VJi2DIcFPQ5/iI+WJ
YCANOU8J23ai0xjQucSO4qWe/zZ7jllhzj1SwMn1AeypkYlSEfv2eIRW53e7dMu3
1AoiMoghWN8+cXX0Ieu9lrGhbAfdWr94y8L39X3ljSHlHuvvfADeOzaRnwg/kx6F
eUn3lQ6VHCSfAxHmEOVYBEvJg4M3kTkXQ2Vu5Tzpw5CBvM7uqknuArW7Gv/qn5tR
e7xW+KVyQf/ex8GAXu6SPTvturbc6u0UvoNoJNlccGyRh9+VFHqqft2pIvFMIu2X
Dfd5K4peKN8BPa9g4piY20BZ+GFhijCvH2nAjMCC9MUYDEQJhjPbav+4JxsfUCoS
tdqtFFLS/AtC8E+glIpmL44nQEiCSuSfenjVCa8hnp09jEysUJGTHg2h+7xUwqws
HIFWnQFmxqfMqV+hhM1MnXL+eTw1ayMWFDezO22BWTxi+frveg33pz5RMVrmHQ7v
aV5AlAmSuoU7OLjG1rULuID3DZrtALX5ErZIuMXGecCE/bHr4QEoqgHS/qDIk3tn
LQxbr2XTT/ZOpqlMYR5PWff5XzO65hoJUsMKom/4mCxVOnAsc0+Zs+LvKMRIqJXu
8xqOxMf7ClKFiK6kUlrjgl1R3YNfYWAESZZuwf3HT7WBQgcIE7fPN3fwKfcoNi3H
1hJwO5hrN78zBPqfpCwZ/l0Gmb2aY1a60u+8wG77D4NtyK9WDnoAwJntvARXxCV3
FIWrOPJhvIyxGd36ft3HEsO2Z1OW2qfzFzTnuuGxtFJLftSSQwOb0179Y0yeG5Qo
YyK4dOTt8r0+vF58LVInkBLf3tICLgqOnT3CjyJSnKTP2PGrGYc1cJMbBicaMC5Q
bnqU9Q2STgubJln75lZwxzIAvGLB5EMcwpG+DGqm+/obtitlLLEyUDNivk3chbww
NgOSzdjpZiTo6jQioc70rScu6HFsrH5Pp8braPLLj9dqZtpemBk0OKRjjJccmGWF
xI0NqqN8vJv8bU37IqcyOoj+lc2PpcDu+K1iJUQLYl4WToaGLAp14I30WH6VYYqO
WLCJmkLEUybkUiN6fldxL3JkwxQKa6ftJTfuOrnzv2UqWLfkzvnl3TPig3Ea4SFk
Toc/KV5EdIOSY8TqgT3J83+2fl1A2byiEnqn+u6dOaaJLCpo+WizEMMHrc3rcrQg
SWxTh/iwcA7wfZLMpcOQ8pVXL2SZ3LJ4j6UCBfM1vylFG/kcvklN+fl/11lTD1rz
onVbV2+FBjVqVYv6hrTdNk+Rmiwg4S5Yw/ZOFzInEpUebwFYMkte//YFM+GsaTKa
pNy0P6EdiNRtudwh6ShiPjG8vCspbifsfnubT1wYg2iTwNjMYcSKWYk4n7GGwQLw
AK+r9PIu6oQ+1wZkMlCnZ7i1rLBkxbYxTv8xeeWiNaixp26tRsg921Ub8XpUhj3g
i4wdvodGsLrwwM8vmOG+Dz4zuvml9XYIEN/2KzVGIxIo6r4n5BOKs914sgqL9R4z
LLJ6h3Cl6CG/IXuRREIs8uz+1TiHyZf+oEtz8cLC7mRsAislylUQLpaGFSDjwrOm
e9/6yB0uYUoM1kWwCLjxggmvHfUAenpJoKEXmCTNm+waMxnH8y8pnTfVo6x3kRVJ
IErAsQ5Lzwc9jL4sL+YxjCy4RS2nFsZ56XjdlxFFFcBX2lcwXtKnQKDdud4zNfMo
k8jbKRqfCdYlW52zZjw844s6wtSTD508AL+ENrBtt/8vFAsD/GfKFBkdJmkeinX6
0fvPux3Pr/DcnwOTnuDta5HvXXBReSM14BMqeTSe4DiM8ahsl11uyPGGPGiTlcrv
bxXx7T8XB0pF+6Fx+vTo8vd4qtP+gOLXG+5to8yg52fhYvXkVntFFOVznEQLvdm7
wTMS3jfylBM5nwIM+MgJ7vTUrXc6oFnQJpYhRvpAlzyv/TYUUSmpbnAGSt6p8yPm
1h5lJU9lAqa31jt4TdgYas2XHLOP3JtZ3C6d6NDVSz7caPdWYA9T1lMPUd4/Y+fW
ymUxOzv0eScDrfksx2TDE3ubk8yqz9pDyb/q0GegqAHpBXFBYsu64ub+BqhyU8Mz
jB1YOtKty3hMJSl/rEFDCApjJKT26owzPINd/MN5zQxICvHLhnve8G7CfluolQZx
UD/LqMa7YQx4xRpWj0y+Rn87FkNsXr1eZ8xnQVd1TomVJ6frYoh6fbjcIh7bzDW2
uUFJjkHwoQNtZ62s+rAT3d5+XxKjiaHMv/vTOl9DCODGVlo5DpIcq9+lmdOgiRJf
3XuGGDrAcJpRSBvj87SaUNTsuerB/G1GAFUIF5yW7qYM9p+eZH8riFoJ8bisU6Bw
L3w7Sq6peRoSN2Vj0NfrRJHSlq+8SkB8xSjuHuj3aE3LH9p3eypgt2DLkeQV9M02
ynkXAoJZt9N9/Z/bJlfJZAlavKVnyKB46pcA1//zYsEuyMVzd2+LtI8FPnCh8YVw
zVNbD37flg1GQhdDRjkX7GVS71S7f4xhqhxhsfzJa2Z3S8c7W6Q6tUVCfT2n0SeN
uSPkoz2zytnCIQS4JYxK5Rs0FhD8dAxUjvtZ+35Ph32y0PZctSn+Rk30lOlwlEB4
MXXlm1oUDG4hQaEFgpTDljpqpTQPRkEoLu1T1aZAtoLpTY/+D0RiHeCZDbVRsjGp
Q+i/DNzTr0Lap3lxwJGmYmcCVFuItLgM6nxmQixYqP9GNXlrekWQU5nJfwtMknR/
2AGpN4PVQby+1NvghpQ+ZMIkEUxFXsn3UFj2UZRjDkg4vd4mIphbUXFB5K9e3Lj8
CTIIjddVTchtF89b6rxbece+eAdkS7WEN4tJEpNwcicUUbxpzpdP73uG2bm7VvOa
LKaJ6FEmRwcOtoLKwAqvgoFmixWc2WSYWutNCkjxGNXT54JnOvTw5UgMbVM6fdl0
7z6N11uQUk0fgq6h6PSr4xWmhNJC3OGIihj3GSBc4vxF+cwlRFZ0pMExKpcGR1ZL
1hHSoeUM2WM1roZiBDWEml7Yh9TbpgfR5xXeCG567SANP1GwNdU9zgFSSoBqBZP5
t4PzxHcbTobe/r8oYfpt+qtC6vXHBuB7vfFfBS/CdwVPrKF3v/j26Ik6dgNuyOaj
XNgUzFKEeFXxf4FxPXFvUll0Swfbi7WA789CoWzyEBIVXTpopMuhfGLWDl1xXIPr
CcDV2eRWAM/WWUByNz6rOGrmGRhMInwe88cMeWFhUraWLszvmHSlwX3+nIMBnM1k
YBfK4VNw2CtyBOCBqvpObpDiWI+Gc55ESmTUdiMDYJhieXfUKNP+C4lEZ0PTZNW3
DJfXm/DLhEEDfYK0bahx+FBwiBtpw49utLTfu6MhSfS8/kHLahAoMk+CTeAeBcqX
UZDhITLT/fRIoPDX6x/Lkn3hNaw5rB7QBbqjZCRimKpuWNJVkPxVa3NJIw2/xt4b
MRZR7/C8yWvivkskLO8RGps4WS4TW425IwsqxV45krjywW3oroEV9gPGFzV3TCC5
FDoVCkHL7tHo4d1FuPmDXzCm86nIMklMBqZRmIwgb7AbBMoKS4jLG7X6VdOY7+ne
OWDxMU+6ZYktRTThz4wGoO/36bz3AkNOj88iyl04Myf0ryZFCDey1dhUGg3bMNcZ
scSvY+jiaV9ftasucp57EtbFMmtY9J6HE2bSHCWC07i9XVeSi3Q1rk9VA4FpTqJ2
tSA4VFVlvyiphpjICc4QsG2iO8IEiS8qG0JqkD8iHY9XfmMQ7C2uAQmC2LgZ6RRy
qpqW6GbJXH1UA9uwQiNEF7059Na9SNjSTy2c1209WpW2tBah8eJVgrfz71okDrb/
HVQUMn5FxAUTM9a1LeKNUwEvLika2iimZeiDK1GAo6jgZJK3vN3OyKAHflH31Wjt
v7XslsU3Sgp/Ftc3/+CBiELJTWpRE7l1ZMzB90UNcKnnvdGlgZXeZj61gBF8bAQ3
cLXrKTgvD2Lr9huMYK2M61TTMci079Qox3CuK9zB1SWXYpM8pQ+yUhkqLDD37sgD
SM2Uh22lSQroEKYEvoXetNQGT6uY9hQCjYzw4sqUpJV8hvKcWlPRrB8sUCaU/mOF
W1IHS5tLpi/q7HJ5rAuyEykyc9+3Ey3NUJTkzwYVvEaEPfX0RQAva7A/Edp+BHYj
zzZGCb1to7smecwvCSipg/DZRGVMwuNPC3XuZA9y5SR7oJaUYGevMVPmrX2NEoji
r0OIMEP7sVcd8JfVBbp/cPq1rXvAcH3RPmf1ZLFBxlZzETWYz4ZOvEyupeQymuUb
J++9uI2XtVy7L2/kuxfgbEFd4i4xbvyqOQh0VkHvzuqIGnhazq3kqqeSwe3XTeCX
crVc5WwPWw3pG1hHhCTZvY0yJLoMKwHNSuNwefPOe40/Bc0kRW2rDQ/RyT/Q1pso
KozGXoXABnxTC2WeRQ44c8yQc4WvKacvSoNLkNtbr97TqXFjq6bQCAdZIUlEiXbI
26+DFJmhz5H+iK+gJDQGxRJYjgnEnyrF4/Cin55h8WNhR78FLYeeR7QVegxRidS0
Yevg886g07lkSQsjANUj/p8eIoNuGK7/+GH5HCA5geRcLawSlLMRyxWa2aYV8NYw
ONpODdMYBZXCOyUeal2rO6EhS26P/NF92+MtrSQ/E+PwB7Mt5sR0iOYfcQoggjrW
ezUpgK+QNjowDJKc9GJhbEZXY3bSJkS7kJuIMR1KRlX1JPkqPTNp6djpqaB8RinW
J1s4IjhIE1pQNTVqReVFooQq5W6YRJntVsXdm9hY+wd509jdra04T9+PPa6ZTpU8
q3jmVrcGtNz7HuGq0ZnpoRO+Aq7JZD+sLI7SkvLM3krHlAUzRLrm9vBlbCZJg5T1
GQGiRTISongK6Uz3XBXkSfMABhlP/Kd7DB/WO4vyvSNg24x0Zf87TOdsr16WbXHr
m6MDvkTWjZC4xiNatDl4EeZl5SADCF/bvLsymQ8TqWoXvY6QqpKF61ilRHeGiaTu
qgGS/u2c62oou7fGahYjLtYUxWa8yxxE4tniMZ37DFcpQggz3MBfev9jCZlNCQKN
MmpYx/fHq69++z5pSofcFeU37qgu4Jr+g2P6Cls6grGdQNvc7dsBzaSD5FjYenYZ
OyBv6TOVo2fNUmwecNSuTrX+tUu/PLcXYnF9Bv8vZ+CPdt0qMxC7Vgp44EuWHNfD
MdOOyOzADSFl8oWUa/MYkf01Gj+tBZUPu/9hS6FKyVCo9O2Yv387TGLexQKbpHeE
lAm/aeUaGcPU0Nm+CGzb9/pi5BbHUKublBPTyMNkHQDZCQMviPp46lwgapLjNQC7
jVnztAC6Fpn3pl2XGM6mCkPvftc6dpI0x9lxaBzC0Y3aTckyPdVXXwqv+3L5PlqW
HZ5eobL2O1TQr0Ze5LtsL69Si/1rmeINDcKsYEPiwX+rxw7HEBA/Ft3BjB2dFecp
eeQfTveOx25DoBvBWxkmkQ7N0w/qcCMPbfmYVwGCTuFuF1gHtpv+S6R4+GzWpyOL
A6stEIFLehayTEnzmckip8GOWGw8n0SN+yCVFg6Nbidqq2lam+RdLa84CmSWseXx
JRBUXOCmQCXvEGXMuMPwGCzji5q3t/jVrirg2hwsqETDPqWKTQfSwluz1Skals9w
oC7U4R009eJ9nflmGqj8dYaGAA/mI8B+803keeYQhMfxOhkHYMQm4LIbPxr4mev0
5tiPFE4VOuplV7GFgjKcYdFR6gDGiscZKTeJ02qfCu4bZyKJyker1JqH8G8UkzVt
M6oaMQDxx3pA5vKt9XhJ+QjcNOYH+I1rwSxuQXteCLhXJVpaqF72E7CCkjOliVzW
lKQe4s3aLprant6KkFshksVpQ1nBNciPedpOYBS3qhgH9eitbzYhIVktfsSwZLW+
2SkgtDOZYgzd+FnCfBl/VIsbwfNe9lDVohVe911hE09PiCfBb1NQEK+sWe9BzCMs
NasgR1hJOJCfmJBg7kc61XCWkofzFnlQE05NokbsTOfS/84m9ORxElIURRSfFIl5
or6bUdG1JhkSrDD7rM7E9njWOPQhVPP1HbB4kVBUev8H8zxGTipmQigUs1tYTTGE
74X1E1k79TH3t6RijC0+tYR/Wt9n76DQ281OIG9asNUKGlQ0za/B7V/U7gynxoes
ykiktyQeKzsLlHx8APDcVxDku5SWnVSYKqd/+lQP4Rzzco2wy4efx9Ovgb8O44ky
y7Uk3VRcsmyIu7N5z0TxA1jhyZRysJT1PFt0sAIZBL1C2KwGOOofGVfuW5zA5CVq
TyZQMN43L37925f5Hhlr4+jNpG6gzTEvAbB4mKyTu9dnDbAqgSbmryoCNWobXepa
RVrOckvzP9KpuLPYkeoNHffkswKetQOv6uGA1/3feU5HjseCwO483Igpf4REv69o
bLnG4TeLQe5M5yg4QWXXJjg+3H7AY49n9bmjVBLrq4MKCMEZGo4vkFshEbyjiwzJ
cgW5f+kEOyBu75ooOjXJyveeQgOhEnt7LkWQbA4NxyoexEZmaHLGOhb+f6NDFpaY
poTpYyNeG1kDP1UPVM6dsGiVTYjFN9TSsYfQO4yxYXavT8Z4ZXYdL57G629EUKQM
IAvq5NfVdKodhpHBBg+Q/HHxXxVlX58u2WiUzXf+UpsR/LLmUxqcM9GCrLo/V1E3
qGlfg1IUdFPbXju9B5BKNh5PEeiT+TJmJDDJLo92/otZwm45jrioGZQJrOw2MsHx
K+UbsU7c1gOMcfqQPpKtjjPCri4rkVp0FVrpYvCIDvezIQNOc9p3Edz3NEPvpyaj
XgEgYgPgB3282oSSUGmp62YD25dTYnYxAD1f29b51SuogdBOZUifigBibWBH70mQ
gV9pHUqJHln+AW8REj9f7VV7ksg7NM/mGqwKtOteGCXlgFDonM4lqLmCXsdsPL2w
n5vIhKrY9FIFmTj59Srr+vaALlyF16H0zBg3vJftG1fVw8aaG/2Flxdq4xGMPKj8
wopUqpu4frw09exjxRJmqncFj7suI2GlfddT/NycGwEKXbTJda0iig1J20+F8z2h
wXVITce9bQRV3WNS8lcSAK02Ztrk9GWHizWKqqN6iUvGw8JzX9HQ54Sx3YIRexv6
L5aBzJat5fL0ci0oWFKgpLpTvbIkfYXGjUlJ5fZ3VaJbnH6/ir+Nz6pZBbTap53g
eMf0W/1gl3HXbt5RqvO2/UAt86mgJqkFNpfjxlgk81WaK43Gfy+zxsla3s55oqoT
c4exTESX/BXW9P5ViSCiCSNDjNCmXZd4BXYatMe9fSSsh26QUf2LuQisZmqEBUhg
m0OxLPSXYRBjcX1H6l2TvTj7vRXPmG45UzarjPF8MJiH3B08vy6GaFQAPSlUeIHZ
w1uPbow60LD+m87okZnAzjABv5J2ESc7bIWyLds9+4RoIHc55X3iGjlqqGD1JPVg
mMPM2coKWuTvySPyZSfdxlQ8GNMUTuli13vPVCIioPNiobVrU8Qv9DMWYUvkzL6n
ANfnuFJno+ngZucmatIqd9LpKNgmqLXB81QK6QKrkSFoTQxhwCcdqPx1VbcjK3TI
U6cr0UEBQkh2oVWc8N9O/9ygTsz9JlbkAKnTgU6EFwZasz6abddqmWLRtomex+W/
l2heNS9jVHKhIq22ksCkBi4zANZt98kbBXNVpTHqXUQ1mivTn0lC88S6XUjgWdzD
J8TC6ofWVJmCiOU2BqeROmpRzAb5NNTj80Ju1wqBWfII+MynfWlrX82RS4v5iApm
tiGW+5IJZLJG0zz97qezgD3Ib7F8kJ7f03/MLTqObCeyxIO4BD+sE/ALZU88YRD7
ujB8sm9VVWi2ldlcoEX31pb8117qYKVSGyrbzwtOXttmZwF5nUhSUggoGTKV3VRG
XFXzLJmXREYivJBTHRioxYg4cltPfyiCmgJTumBsQ7HQK4yhVvJV7FrfSF0bwMN3
23Nzu9Dy48eC0HuDb6lXpIHneLR8Kr8TDt/nWudZfvxkJJxzLdWIf6zXeppq1aBl
4Pqd/Chgyt3B0sOTbbbC7i2lCvHja1VovB7DTAu10geZqOwPmbvJoBP3ooISDejt
wbBVgvvVFU/yaZ+caNqdNThG39Snr4LjJP+6zDd5MJ3fuv9ECouJpwLnp9dL18ik
ifyO1BWYLzTlTmb0+KeTFug8mt4RfzpekA2xOm4Kd7mBJ40s+Ossn7oNye2qh2f8
aJsnRZ+5EGJznxQOajmUHUCZ9p+ospl268UiP9IP5v4ExAplLKc5izr5HohAzyv4
AQSPY60SN0mo8IGdwAwDY4aUJ0qHW+Q8qAkN+23QWiFwMps+KRtPLc5a/tfXzxnv
2ftMdvcetIoQJkFqawul+7aVJItMctaYAUPvouDYpWX+6o+vBMH5rbpV9XoZNCFF
J5xZVMZMZCYwiKg+VCWkL9nV8fjUPUZU9j4FdUk6YsUmdqUvBDj5o2Lbs1APTgxp
A8DWCgiUYK8wSTvfPAi5JRnByCfQNgHSO5JlH1QYEof8yRpDrxjSVBa2aBeqa+b0
O/5t8JBHSbnutjNTRXBp+OobZvmoS/D/OE5w1HKjNQjd5pgEkfTFrV7Gjx3uhpjE
ENe2LShjR4vb8/2MVwTEaahqiHsLHVr96PYP2puVx+2ZuvdiHLjTpryHnyponO/b
Mj+8BXZPvIFpqpqa5hUM0Fws3ZhCSOGpTGr4+M3cUDXf0krjhavvO2iWFlpjpG/l
HEyFYhnD3nDi3SaCt/E8bCd3ov6f2On2iRj6gBoPaQrXjLHaMd4R0gQJyqw6dMTo
RDSSpUhDO7hfhGXTSawerjtNudc3tGZZwfXlE+CT7G6BJL68y/1wE1FMORcvB6HD
TAuGGmwOFkH16QyYY/nG/6NHIddoriYfkTo5JOpuGWesmf0YSiJGe/0mbAzNKKu1
fPKe0VZOu5+LEuQw/TgA6U29Pu3hgqp26kwXWidVRgub6EiG3ZmUSEL6e6GES1p1
Vjudb8zArE40k4tgWUGkr6NjYfuuVFjSw3RI5K4lMguagIu0FlouOsTlkutf5a2h
Ro1Uq5BQtsEvY2/qyVGWl6f293xU4C42QfAXwHkKc6ES9iMo7UV76xFeuOzgfXh4
4Lm7UFb/ReAtsW65FJHr3S3zvzwxJ4kaHPf3/3JealNCbbeK7nki2x71iKX1rAt5
1Kmyb+EkDujzBnf60UH9f5kWnvu6VK/ClYcwqeSd2lD2e3veFYBC8g7dPcUX4x7S
ljEg9uE9IgzYFv8Yj+u/qosgh5HWBAP1U08DpKGlG1xx49k/0Uq9iMwAXs9IUEDB
hxf4kv5LpIPAHvv0DI6lmORrJOTw8VuDeQtuG5q6F7TLjnDEg32YKFk2RHBYS7KU
7vJskI+lOOumXYWgAjPR02BFG7Pf1YjcVKs6z7xsdADekZaHJ2ruAlPQeSGbgf5P
Eh0aIpjGYXtncx/Dx1oZaS5HEUw+QMWKKf2XPFgK8lAh0tD1NjMz6Y4ft0lYzO50
AxZB4kKaZD+so9h5Caiu7wgq5XqdM+by+trc1R6UcU5LxPq/TAJbfoxbtLle2HAV
QqYgss7XZselv5kkpOYJPYzh0dZ+fdiF9jZkhNHRu6GACkA8Wv4FzihuM7TcwlMM
DDwmwN9yHZkbJXzoovEjgJt8zpGgpSJaqWqXH1A/17RCPGXImhB7/QM3hgLbp7Zk
EBbymkt/DMUEwryPZjrUegECEPbr2g4b+wPqQYa80J3CBAv/KoF1X/BR4rbwtPn+
KiHmi9vQW1yKtNXfx4n2rjmP1k7FjdtVi5ueyPWyEA3NeV2s/vRIast6GMANd02F
oW/OpUHQD0FYNFIGHBkPBo010kZxIlfRE8ItxTWMsJgolf/Hn89x9CLL0mOu6Kev
61ag7DjWldufkqbzgZu1fqessfUOU6tjqrUPg+zT5LcLkN8oIloLaxObwDzRPz4W
ezCUPYp0+IOY6YdhZAU5EuTvn6A14tWVnYD+mKIcjHD1HMTjxw6pcdJZmD7N17lR
cZnu3Dp8BogLhgvC6pXA0DEXmfrYqh3WnuX7gXgKIhko1ascQSv4GAvQJ48/KE+H
PPof3TaaV7RcTcK7vMH2enqKA01XGc4Mq+nt5rKeQVS0zHcrNNyLIyHE1d61qj+N
5N9fL5W6KGMEdIBEJ5OiU5F7H+G0/J5/SjMcWnwpC3iBkFDlY/0awnwQLsesBDir
++4oY/pFKtfo4fA06+SF/omSudZaZ4xO8q1lBBpUjMNLfIZVFcYInfV85tW8/vsM
f10hbydxeehDPv8RhszT28UKs57qNySNtKxk7+L4cWV4Mv74ak2A/9y3+LrGFmby
Dw1w3s5+5I6xKf1r1JXk7IuYTxgaQvv13GyjINg/bZ5NjhITCquAoMIo4vZ3xuzc
qNa+Cvb6gBaHcLhsKLjP4ShjiormFB41TVHvsXFioZkRg8qCy7sv08aqLcT/7vnQ
q97hWyiKX9igNs/IMv8GvJ0tcuUBPoj6t7G2OErW/wPXIV+HCflkXoDXI1IQdMcC
FFfbVN6+x+yQ6UrsctDWYtwNCOmN7H+cnqYvowduOZ4s74GCGTiPkMZPirPJYCsB
7xx9foyCk51qecU0Gux2QHpM5q1U3xqS2DGCbRmqX3qJymuUpASfpCWYSx6PDtIJ
SggNo9ZGTzIzHfcy40IwXuX8wIF0iOGVzK1ZcslLMk5kh+2+8KDC2zoZHD4ESdwm
/7vDBDhCVtBb6sOf71GJqk5W2X3JywCJwIa9Jq2x9uA6dkrBUebu77YMjvhSC9YJ
puwILq7eN5CU4uwUi0nWRjeI3BKUijkmMukJYNPbQoV8kc7QHDfL7xiHhktdCA28
gunjOhuEPoLEPocP7QurmwYLufRzIAJNfYHALJ7a9SdzSpRpKq4/YsJOMLJ7GbK9
NXO0o4nIfTyfwMBj8HF3t4IcQNKywsyetg77we9K3XQhFzZRyYSYkRS7s6Dc4r3t
Hw6EWkskJGgkeWenPUQH16NFlsoaoCpDvT6PvElP8NfaZi8g2u3IRg24J5coeh0U
+L+L9QUsRReWgCYqPR7luXWj420f9SjzjNV/UdW7XCVsuCqwDGT3rXcjGZlKGxv7
v7ppM8k72Sp5Rdv8sVRcXBLIkd8AQDITl665OQWkONEieKREQjBVUKzYMdU7WpeZ
+QhyguYTbeuAxaahKhBMPNIzSAZm91BGrUt9PQ1u//1k4pItQzFvXwP+2fuBrQdx
CUjmpF+/KaUdVWSBZwHEPK9lUUEcHEOvO1+MN7XOEk8/C8plJZewPqe+ah9ohqKR
47ZndeaxCGFU9JcIgEVpNnwE/RS/iq6ijNnDed0K2k9VJ7Bbiny2BUkw+1eeQQCQ
ki0XMu+sLmn8Wnqa7B2qiKgwQoqpl7TXfRgvt++nhoCXn2VHr94anDM1OjayQUQd
H/lDHkNTYF5DO9bMS6kPfSuz1AYTYdA13PwmVmP6qdc18Zzluh2xNwjyXoTlcDTP
/W/TDpym4AXxqFJois+dNwGeAud6k9vDe7SABFTIgXtS8lNVMGGRgAF26zjISxmY
el5iYTz2A+rnM5RKyrAHMf8L/gUGVr9OwDRTWWU2yu8ft8PsU/5UDUP9ZB7NyNDZ
LZcy4WgwRk6gP9xPHthRMGFn44zd5JaUHqKIlPxd0Zq3yK5rngpqRBLjWcvmQZEp
NzuIfYhDFAhDT3ddds+mf6WIp8iU2KlVqJAJzQfra+SuRu9aA+XkB/90WX4nVbuk
eRNQBUyzS1VwX0heZIyaXIZJ6ZX+s/QYX3LT6EccU8FAeGVa3K4d0Wd8svqir9wu
t4I51AZnPeqt2oFr7AhIjItkigUEJqVbP2aROigteH3o/dGswtDZ2oJ1S1LCZcaD
+UzDdDPnZ891J2Dnft9oRGYNPztAQfeq7K4YNV1UdUoGq3/tcAzDmnVnn58aOkwe
6+59wJpzAydtm19LRqBMcFpssucWRVrUcZUq8GeiORc4V+Ov7MBiXMrzqH8Mcvdh
csY9NCEi3A9VStTMsgLiEU+Z4q0DqWE9Sl0eit6j5WAABHrd+M1EGBK4rm+3nv4o
Pg58Lt6/uynplVHHvihdjVtLnZmTIxorxPQRnWAY/NdLpHL7uSlCL+QIVHMGMRmv
d8A2uBR259Da1GvoZWpDVq1jvgetzfcZS8o7k7Ir7aIe+kl08NEgQ6++hm46xXOy
hSxbKgScIJ1a+tsLrDOXVZSlk3GR/O6kF9qA2VIAo7TFhFmeAfKkMOEp0+voSYVK
M4YG3CzJQNLX1ptya3Kru09qwAb8+BVEzpU88y3mTMjys55vOumjb3WSLN78c/T6
zGLo6KkY87yERG9jrD4HFv4pJu4zlg4jIcu2jmZ/Nh/hVRP3d3jFUegBAehvpOpj
bfUFIJmJ4E9YOy6xqe6PVBu3+XJsNU3wJIaFuYvVMSGzpxPHr2c+e7VjmjJYouUF
PKnP/oc9Po8H3OEY4WWFPZJAXDoVAyKZy/jUhsTyjfUcixSxhzwmXNbZOXeZb7C/
Ve0mucvANMjtFuwL5ny/SJ9yh2FmU3XqxkQdMk7b9Xn/p0IvEtkc5masGMqVEddp
mRYv3kDjBnUm1UB7X8XDWGuGOR9tCr89gmuYhikY0TV4bW3rPLzAdjHNiiTBa6PG
rP59jwbh+Op0CugdFYrrm9Skz0EQtAPTCiAA/TOq/xBWAoqvb5/kFoBEl0AuU4Hk
U6YwSp8cxu2bWMd6IMvI07/W1VPZX4/6lIplKwYSDD0ujKSMvlWFO/XL7p9xbtGU
jHm7EJyAV+Kt+4dyHpH7c+QJcyYDw6jpf1INrnsmQYsy0lbODQ2NFv8nYAQA8N14
8rEafxeaoirphAN+4w1F8Ri37FLERbTe6Cp/ymN5DorkKFdlxcz8mzfNfIlFdt8m
iz2FRauYCVoIcAD8j5epaZYymQtbtETHh3ohPQC5UzNQZ4ol9nitH5YdSbvgz0g0
CG63UI9QqefJ9Dk5FppG54dZ1d5urxcQqc9f3v7462/wwsomm/bHppj7AIo/WQ9n
LgE+gUFZPVES8TJJh04TRyL+Obuf8DH3pimBXhb202X3Qhyxj6tTwu0e3wKtg1Fp
xgyhrpSdgrZ4Hc3JqP3MDhPHcgQa8XtPgJ918ojlCFM4+aCJGJCNfY8W1iLox/7i
qZJIFguanAsRi8c5lkEFNkhQb9wURODkBSVyqEnkvtpZkOFSvuqGPbX7+bk/DLGG
W2GUd+7eqWhdozhPpkwbqZPRHN0nvvcogBW/PbH96e31pxiKjZPJ5dzfewdssoFn
H8J4XnNu75I7PjJvX7e6CWapMuxKjehvIW+fvVuKnuyB3AuoBXZ2YG1omZ0EymHk
tDKWpzmEvBg1+yJQmP2jfNDc7uHD6NneZ3Rmy3lBajNVTxr+THmI+r3EkX8bdNdu
EClpVUZ224xry/4MkYRjf6Lnk6TQed0F45DXAKcORs7xKVTPJ5qtT788Mbogo1Oe
o1jd1OgCGNstjrSe/Zw/dWI7b0h9WW+Sq5tbQ8I+RIEbXmd/Lj/SPiKHl476ls3g
2Gt1cHYbn6kr8odRcsDHQ7+zEZeXSmrjzZcSe63DM/8hVohrDAzmrfMgFVl3ajWV
UXYc61GOt1+Zy7nclxVdxW+8+/vi6I2ec6eyqXehufaiT4AUzOYCGVnw9oW9mQr7
JGyf49Z7qdeT9HheDa+oYXUwvus4pjA4zUphCkJsdYouMMY6wtciHxuUeUK5f7h/
Zf5QnOjtZ6x2h3OYnCTmx4L+Lz50N13r0gINIiICe4jSloxi7id7bHDg6P10yshn
zjAjhDeYN0bxFu+C0fD/kCfEowwY7Vvr5o97CiiSjEHOuKrPFt36jG3eNokxND53
TOqfFWgw9bipP6u0kdn/+1lmUjDAXr/mpczPdaDd2x/9g6hMPll23rYL8pW1FvSZ
y74gInQV3elq0WP9wh80xori/IqLJH9KGxEnA6WuiKjX6WdsIUGu1mR5DxmCuuMp
08uOFRXsMThf787I7dMSr60mbIAwpLWbuoZpcSuWuq61P9ku0+htvrmkAIfg2mZt
kcx6qdBlJ9NLDOCd8iyAfyR2YBsUP/+0gWDeAaj1YbHW3qkDx8OXEXng9eniedtE
Wvnq/XPWCMu6lXvucplIIn/vKGR7b8N4xcAQSAlSkdlPALtmszRF6fBH0Fcn0K0W
97YBm/i0hkL4CeIRMgfoZVfVhv2yZ7qcDw8JIRPQgaPtVIcJnJOPXeDZCOEh1U+w
nforJaBRYTvlHNoY6lQcMP9nJNcrSdLii3eLpkVSd/ipyfs/9ybmwPpDsxeGtDzJ
iKLtgvBSmR1/1BcqTsyahZ+eTWYRZpsQ1vneundHWrQ6lubf4cFFF/Wgv93D0wCP
nlhUIfNFPEhsHTchWTIHfTYNm/0P0Hd/qmaY2VMvzL6hgVVDt2F19dT9tNMn2yuT
byDMcnL8B/ABslydteGAqXZo1Ch/tyJNbch3ENQ2yIXFbf3bAW974Qg7xnlyxuYn
SyftNOt0VNoxxfjsUAYIY1bMbS0qOl5SZgZzpUioFYWmVo3pzXERGaoJj/i8Xc3j
LxsIyibsOyHVxHx0jDXziHfBlbR/S5/DRSWqxztjL1XQE41krI8ZNTcutDkz+HeS
K96cB7OQYYO1Cksrcz9YM2GYdV1OYC2dYPHEI1QGPL2HVPZfGAk0SGn1OJvDun+p
z7ifiuZNkjn8LhT+TeQOzdloSoB1LMISUZSGEANxJt410do2S4dt4bNnCQhkWSGa
OhTe+6+YXXTjfASgaMLq9DB1kw8bDBHNVrWPiQ+s29jeBBphJK2UWtCdGzreN7hf
lG0iVHrBzO5JDZLub4MWqjfL+I0H1khkhfnNIWceJ99jJBnYcHL0+AFU0hYUPPJf
zf4JL8C0d4MQ1b8IsiGn33Od/OIJjHh9UxAQy+rpvjd56mLcGccxE0KE4KXvfw59
h4KJM4Mu0QqCyKwd5uasr7cfTLIb39xmaobXgXrhPqn10ZsC9dpjhlvCIZnDctuU
8ldoBdHrIi1ynniAHyM3xRqMWqSORcKXAPl93yF77UZiRq0QF1T6NJjc7CKBLc1Z
2HRvxJW2PFXeweOPYPYAlHMrePNP+RQX0rZuJHY+7DLll7sT+/Gp4yY9jn18wqOw
Xj5SfodUmMPoLvaEojtFrnHgNTTIW5L90QxbILjd20mvO/+BmDf4AcmrgOC85DyO
6N5MJtxeb0ohByLnT/16WO+UODR5Fc9GliLewEfUv+3kHo2okzorzYJNLnpiwGe/
3BQE4R5MgrJp2BvbM8FB1COoFQmsHMEtOWuk8boJ5fOG7s4NogcpbE+tvCg9d7oq
uvt8giKMHFj9LreWmP5o0w0xfw/F5wRVLuzPuGEsAXVTnySCVfffgX+X3VaLEpjl
HRd5F+zXPvmjZiPGubD9dzQJ6OS7/7mKwXafYAJX6iI+K1QxBdlP5vV6pK8uEgXP
qPZoCBr+JzNOCDrSBv7VzrzREw7USWCPhfiY5iySBsz28eZl0HXvJ7WogEcSFSIm
l/qXHVbdzMzMk4utFnGwWk6Z1LNCXnFmJ6d3OLuFzAFzR7qR7wklBF3E+c/3tqLg
S5+TMPoEG8d24K1UBmVZVgHzMj5Nr7SE4zV4e5BkFXvTnSGH/pTxsZ98sKWcM5B3
AjwkhdUobWZhTX9oglOyzVQCdfrrE8a4p9SBM9tTJp8PzZ+YtLKESFi9fZoQwOXA
PnpIRN1dOgEONYephXW+AOgbd0/rYiUjhM0bDn2fajano3s02bSpU2PUfv1BLlUe
Htn15whtEX2qCw8KhLb+Y0yL49ZVJ1QyDcJCosZ4zukXCA6hVE5GP9489NIWqXNZ
N6yu5KiuHSMfIYmfTdLcfaYYtBt9RRMMdcROYuVKAGryy5h3TjRRja8IHlhYIJN3
tFyQwUnSsBIixjQjPU/QrMD2aU3SfjPizK/mnv0/1i8uoJWZ2PfVQkxOrguRwRfm
dYMZnTJ7/IeMq4mwZQ62JGaUTYgr5sOeBQquj6mWogw00ExvB5pzKD2mPRABdKlu
B40dg9kOT7s35tSHtE5H4+r4/DOkYCJBmdD3PeF/mlHy+Q+W2Bc30vhmTSmIXpiv
s0at04YwNGGxfOepP6JRpagkhxWut7jaGLHOA5uEL0LMVQ0HxI4KddFtLVZitSvo
2V+No4A0wzz/QF8b3V7AUGGlY4vfh1tUghqNi0hXDwAgbi3KXAhd5jmOjYXpp/sB
qDuz6TSaoRE9oINAIfB0dzaE+BbYbpKyboGaDik0aj7n0Itc8mwqLc3VojW0Hc+e
`pragma protect end_protected
