// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pEABeI5aogvOH6UIQzIRMw/chzc19H3yYR66r8WNsfSjQetOkqO3SsBG047dB+Mm
+NX6KWq4xogBAeJbVMfg4r78uG7MumHirn1/VAO11EUaBJnCKxYwgzix9mmschKU
Oc9ccWhXiHovFNCu+U+jZU43OS/itdNJZZct5Wf0DtU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20160)
3Ti0c3JdsJIUI8ZQjFtMpKW2ZuxlRK6x9oyb9krZX3fxneXIZJF4jEmizfjtOcHL
tUjwN/o31hrY5zXk4G73xy49qbSKf/gpyzFHY8ZS0sFaPJgpo0xhiQmYzvfuFXzY
oKy0PZF7dfU+/jPgf0OyShOG4WOEtri8sUgsxiJHlXiIrucBKAxepjlRczmCZqIE
Vju4f4ry5j+p92zT+30WbZWG5rQt+IJYoaAEITMmp1auC4R7b34qhuBFI6Ga3hIt
g9ThTHQPUBmGdaSAevpVtZlspbcQbmzKJ1NrS8u1uCgds0LS1p48E1Vs2oXiClxD
VAUqPMP5jdsU9BrX4gu53wSlmOdWi+VSl7R9jwFEoCzi6mzH9pNh/5X8fBDpjS9p
mly1WlExhhbnNLSWdFTKMiqcEvzmt2zv3ermLY4HfEsh/z3alznSgQ+i7jCAaIOx
4QXVdSmQjf85fCM++g/7VvlDMa+FDpSt8Kh0Y2XPI0BehNYjEOk5CN5dQ5DqBlpA
RM/EPs9r186OyJ/DAB6pesUYGEHFW4KyIBM0A/pfjWxZkp1XA8u6pKiVuh++57HF
p9xC7gJxnkjVfHWsSjSR83uYe9nM4Cys4lzMzWk1IOSge2XwFx76QgI5+X8/OKu5
UrIO9Lx1bINFSqZ7i+8xOoVg1mhuONoXhOHM2Fh0aI5Q/D5f51lVcIp4TTrgKrhn
Qkw7sPEpZvhoE2JiJu+ti4Vc5vtAQwsFkARdoc4fQtuX+AJmcXyGYyxUv5m98YTI
dlo/RFRj3RavdsMBSc1cONknIN9qCoIOnaWCK8bMWtfQ+fVZI+PSwOYfYMd6p6nH
2D9/j1O+Rr11ziKM9Jq7VT3gzuYhZnSUa1id0i64JT0c4b2RzqXNBKkPYDoBvRki
IZC04h4L3xThEsUlLYjYIeVnOioDm4cYMDbcn77oDCq+ivE9HByZ3HxmcWQ2MqHv
5ak0uWbltqaQvWqWiBeDm61acTOJeHuWwK5JKuBammDMuYQaaLr7oKLsdSt7htPp
ftWUqCmnzBxuSa1qtAFxw34oyx1ntyxNa3xsOLIJvwZm1Mtulep6SbRCyK1oRBrh
7YqeATI2Xm+4Z+bnGo0VEuh6eLDseRT5fSWIr9y3ivj/LeATf869Gi+VrmPqnLRj
0sUR8y/4itoNJOyUpKcvg6t7euKhii3iCJPjUOT0JiHq1If5vU8FdtbI0ml1Msyv
Lq0U3XtlzkTmTTNOTl8jvGt90cY4iQQ+lUPbtEIBh1NxaydwtCzMoQYH6+5CCz0v
Ww0xJCUTugB1OGARqhGiqFXLFsq/3nXcKgrV4bB4nzSO83DG1rPNBo+2aJoaGhuB
p9SV10MbFnNsN5p8jOEjK5a1SyK1UanvKKuBFAJ2KvDmcJbdC7vdT7bh5VeH9D/5
VwNpVmI19LfH5hIfTIZPW3de6m0aD4CWPoV/MOm0E+oOaZj/IH39r1o7EwZSsGLE
eHBWI1M9bb4BP8DVViD6r2nz2bYKEPBdIg6CI3rMVB3OJA3tY7rLmTeH/CEq5kk5
OQkTcGzu8nR7MDR2moRvKeidsHhOzpvK71JD8rwCCg2zcZLm+44ujBoB0hCFDbz7
Zizu4nQP29vpsNfXQx+clResppTquBu8S5xfGcK2zErhvzEXIXZmFYgKjE3Qr3XH
+C0xIqCQou8rXaBE3n7sp4XTl4cHMnyTfP3FzlJIrK6A5clA9Ur8kGrkmIzf5t8+
FMxAe3SJXRx7XxK5FwtuEmqmJ09lBjtDQ1pE3nJNDa8rgyfoyliLeicdlPp4BBCf
CoEtrxe5EmoZ1+ox8nDh8x93psqV+WOFsfZ775jXSn6uHMOs7WUEVzdIgDtGaPkU
gd1GS1jlg0l6iISPRekwFiqkoN3kmCfjbABk5Kb/ZK71A90k8RBiqwSX1zakDUM0
OmY2ndeeB5Tk06Lm/3tZGaKfeRssXZ3LtOrwARPF3yZ3hhvWp2bpeEPXtek90e97
nhHC5AEolYo01nh3YLMpGApjZw2icxMRO4B4YwuqWgQaKof1++PKk2mjUSww4P6Q
trJzaSR/oDbvQrOalJoCHzRzFiZvyFyIqHBnr2giVVMHkvJwyHPZaEdDBmY8cG4q
VjqFoka0N+x293kLGlVDC6v2XiSHHyHUk+pqUo9mCBF/u3fO/dAcQa0CPPHTcrCv
6iKtqb3iTFpVp4VNFDTU1G9WqfQt0CjsEVGYS8MDyIBWU804CcfjL73fjc/iUg8w
91/klM9Nt1t5WSXyCifFciYvXUTGEPxiDEugSG8fMoabwxVJeiXVQ9rIYKZkHZq3
vlyPMbyblGN9RK6SKT+3t/w2PcnI+5eYTShAEvQkZuPMkLPfDtgdJb762i6xKwZS
wjNbRYQlzcbgyxMmAVwRFIfofY7JD0Hv8Mh37Vsuj59eVEMvJQ7xk0YdXT3nE4/j
Zycr0VuliMzbspRWxGWyFTP4bDmuQDtwQ/f3DI+e2hgxNhvwUXR7+VrtS+/PN916
wtPg09yDEyk9tdEEsmjYkFxH2zR7AgFsnCO2qe0FbEGgQKaP0aWwdc1ZmHrLx8pH
DCAo9S+OLPZfU0Qv+2iX5dVtPOQL9GJ/ioeN6eT3L2tBjQiwfenmVv563/OZJSiC
aEfmB0Q7cill2wckiF06jeZTQvBP+x6epA03q6kBGmC96VhBMDvz5CruidJF72dZ
xyfRwwnYjODg2bR0Ih3cAtFsl5tr4WLTLXjl33o3968fbZDKdn1TSdf0FqjbZNad
I7RB3MlsPmkJ1eKp+MHKsUyhxao1Zr1xeQ0lrV2LPuwHvw1UPpxvufQsPKUuMZ1W
t2Z/bgJ/FndO5I2UjedTRhm4tHNBAdES5mLo0MbL76nZN+htyWtttKjeyFKfhVyn
hrXd7zfjAP2JeKC55Nr1mHAYu51UtNGlq/fweouOjlV+xCXJhJrE9ktQT+JvUvov
eh/a/6/L/b1eTnSYc6/91wIl2eej6UoqsSLY8wQ0oB+klIq+YkLI+J2XLH2YCQIz
Tqo7Cjk9vdRT7VYv+hEcwOpDbSkH79FuzGW01dFU67C8IpFhbwH/2lyxJINNybxZ
XYC8hv7X1ZPmq+ISGVr3cySrzT6Ddwn/7ILqptpyzxJlm2ujHI8DoQxPy5FMxwhb
xORoNeZ4ATY3NNdU9y565sZDESwnH2qWkw44MmAu5wPYrN1OPIqKoluAp9dBOJ6M
9PO2jApbsiYuQZVtr8nCr0Y1ECpezWPGMmUl1+GoQScFTF1f1pUZYf4g7SvxLjBS
OZ8tjzWvZtYYmWejOfSKQ1qzKdVcxXE9gmCBhnWYNH4+/f0ZV3vmFvoRm7TTFSen
xoZQ7bhMXEtD300v7PQTg2XhbUut5sl8Msi4ejAfC/XFe3sROLTs70/Bckym3Wmi
A5PawXGFNDkU787ADM8ZWwqiCw4yTj3Vu29mWF1RlzpZO5x6BDloAXuXbWJZSaAI
dJg0GsBSOa3UJT8QBA7e9autIdpFYQA7VXhYOgdPf6FvAdqOEojGM0a4txRK3fTU
U/ygsRYpe3w3/rYyb0NFv6Ldbb3zBNfyKxPYR9fOvNN3P8a+H7tVuDGVHzbz9uhS
QoFENblJJZnHIaBCWvuRtLHryUAVHFI3FE8+g++cg1b8BP5gLclVQ+TQ2i0aqf8q
jwr9w93EjOc90IzxXKgUh+MFjHwQ9RPlHIZG7zrzLt1ak3bXxYVO1Osd5rXRy+3z
6iokQBqQzGP+TmIG7hfy7cdY/4U6Xe00KfM/nOjk76e9M1re+34SwirGRmdLL4q1
AwEPOTHhNFCHrgaS8FOhg4bI+0+BDSA2HDKSaLhRoEdLLKli0Ff8PHN5Y9MBapKA
5G0Wdb86kcrVkud+lZsXT4UgaystCyjGz+7xfhU+iOd9A7gfhOtAUAcuXtUbRFed
0QlGgEBVW7D2KkKtEjCwmHkvZi2VZhuFshBeKAQqwLwe8ZjKXvYr9c6vq/lUaoIY
XJU14UtDBeNiQ+7TzRW4L1B61eeDXrS3ol62pvy5fz5AGy0Laa//rNcGcM7Cgnwy
QlGEldUwNGs/EUnFmJnFii6/z9SfVOSqqPyB/7QuAHZzxSQxHZOgqhbUf1bhOaVO
D/4rhYf4aswJd+yxheJL/u0TgQsiAbCdJC9cmAnx0vNitI9e5Q8DU8rMQUsKFp2u
0nqaCQ/wVBMlvitkosRP6NOTvL2z+s+MZ6jxBm0frrstCVyVEYZNZVToSt6Ml/vF
7DPKJNn0AcAP+ZcYs17x4gfQsNZhMPhL4BmUXIZTcAk8tAwh6CbXSwjURcYH+7HS
domG2XsJn9ajVGkcOJSYWZAZTqthoJfmmBubQBuRffc1ttzLVqGs/uA05Y7aMsFT
1Dvelh5aS1EBMkl14DvmjdLgN743NPe/I8+56n0gKU+Plh1b7FoouPN972VOoYhq
F3ikTTJUBKG7cUVPhfpSUyYEptftCEJY04dtwBcObW2oZXRIPCcbJSpDw49Ke7HR
vUj/PRX9Ul0kgtWc8ughUrv9gztWGa6OzY+j/nHTkds79EyvAfDTXyIHbaecgmjp
iydxhOaJBkRrtHBFGPv45kYYqxYkyYaFJNk0SqQ0ssNGeZbQgRj4ObxdFYDQc/yg
7nuSSsUAVK+DkgAUlLmYjy4nV0dcII1nKxnkFARD8EmPFX5ULZK9OMxib0Zazsgk
UkhSzALmzyuDO3aO2kNedNUUP304jt235WR00Qr2U5V+uNWmiK4cIFFGE6kW1PMn
wmUR+C34IRfZf1sJWB/yofO2WqJLNwQg9q6ovkf7ljd5c5NSwyZi+3EwZO3JC5Bg
SdvUdFjIS1eafsxvTn5s1SNtJRUNvxuoDPX0RL5j9unKakSUmhhgSA4WPrURfBiT
zZDJQXGIhark6OswsMdXszPrDnnrpZ6xkGa5H3yKO95gs1DQPmtN2WvTAnx1T3+y
rfh1IzJ6XVXe5E9ZHaF6x4KQeqswBqon3b1hDON2Ax9EMRtkGSO/zdAfE3Z/ta2q
cCGAUZMw2xdR7Yg+HrVfQXIcCuc5/S4FjT3abhwIJB3tmn4/3m3usxcWhvcgkr+V
oK4+AiDDQUPfBN75kGziHxaThOvJDr7ByzyECz9sFog0qMDvg1FqaT2Zu3HytpEy
hALtGSaMjAXszNWKw0ZhKQdTVTiUnKyqD+hsyaBgu4a9PBiEAw4/KDFrw8F5DiYW
XtCYZDOnEOVMzSPSheeFwVzHbQSBR6ZecFb81vsiLx2U3NCAAryRfjHXiY53wN82
L2FXm/1gyweK5qzhiwKXiCbyHVc4tmLfb7mQK/5WyKiuvl17GdCR67B5UG4lNU7b
ne6e7NXloUZjaq1K7N6KBdP6hJDqpqAX3jwB5XzUb+IHh9MkeZ3WxJwZYQ75+tKH
aTJfPAot/TFu/kAlxIviDhxAqbzuLL1kMcCZjA8eOyKf+RxHsuAL+cIayAin9y5A
cwLFBXDjGj/absA5tmXxL28ODP57h5eF/rjfUOZHStkmoWFTFG/OnS3NPbZ/cNfu
rt0d8oDcbKAXZR2ZzaZOTu2MyffbFv0PtnWaDoTeD8PDtoVYCPNPtjDp0d4ER9X6
VfrNrE8viy61YK/U32xlhbEYrsBzd907kXQQ9xvzjzv/XKMZj61w8fv9Em0dBODh
3rrV6Qdk1Nk9Y/ZsrZopmrpMHOTokOky3MRZorkequP/USAiexcH+SAcO2oaEDCf
mvC9EMY3dEuCBAhEnex4gOF21v6/ea+FmJMqOt1MguA89My6mzSMss1WggGOOldc
bh6yRtfDnrKnnTSQkm1pK8oM756c873g7v9PVYku3+pT4vGs1H1EaqqPGwGZ0Lzz
QoG2wzazpq0X/pyXcIC4OzguHqNISivi4Ijj1N/njQKKQyqgu6Vnfvm89dZPhQOu
CUojWmekFS2ltgt0hmBHGyjrkAltGVmqDD7QWynyiDPu1VZJjyiPpAiyyF2wpEUZ
AkdMVaxdNS7uLv51yV5JrrDubZKqen8+IzP+f+DiXVGN40TXvvzaVLwBbW5fAQDX
Fw0pNeV5mLMVB8essujI4SVrHMc/rWCGL9gtvEEwu1Quw3NgtBTA1On8owW7bF+P
LE6aKiwR79gUcokA41BZcGFaZIZ478+64H8Im8sde8wjb/icWyXy6TFpWMmc+QgN
jE+ClTtjaLwQiyZliNFjQ/GRnM288gSPNIpdQrYYwjekoUPu0kkDtN0k84tibDA5
F+3pfEGiANZSHihStTV7Hxw2Fg/905gEQdF14g59VTW5UFg+f6vkLOvQVXmGnRgN
zTCyc7IpvW1uY6rijqhTw/BfNjmepUk9/MJ1zqJBcb4eptXSqPZ/AYlaRCs32HTl
RENGgKXA/BAlUmyu7TbwVLrSYoVpNpOTOZHpVUSkdwBVqBmF7dthCr80cDtNMK6L
5wecbZcMZXWGw1vjApni9ElaLKsONuLuKfMOyPE4xH6VBKoY22dyyc9ZjgR9Ke5S
1riJDQ9vPozW8zOMp+fnsKzAcdZoQ1DjgHdTNpp6zmC9QXm/al2z/N/oWSsicXRl
xEOcMg/7F5JAwayz0QrLlMlPNM7UQohQZi9PJ5gVK+g+LS2s3NGK1TTtUNcGk9us
W4uC5qtexd+wwCCXR/rqgqLZ6ssgonEVRZLt92E24YrklurHd2PHCgEp1qId2e0b
W1PKqDVoLVWpoL4QJh4+ZAtoLtAFrBZKaiqESpA1E3K/IE8XyrUBlo59Qzh7Y3qx
/2g/zMfa725UrsS/c+qOghaq/xI/8aEp6XM7s7cti/QupkZQ0RC82a+8nSx2J1YY
q7kGc4Aw3O8oKGY+XBaCsmn8chyrIYud58jsKxnG7xo1j15h6yHzDo1CJODsHICH
Rx9QGkjo0Y8kWEBVahsZryetochx2vggu/L2Do5mBswc3Nb1sm4W3zCiuIeGsYoW
6piHPvThZjydDVEZg16hhAA51Fw7wYVR3EJtOmzvailR1NiQMO67PrfZvGIQ/R+r
lqyDa3Q4AmrnJEVUKVsLkLIwRwP7A5/DKjGLBGQBXXEwQ1n2Xl0ksmSyEb7GuTo5
prLIsUXESKfKRNXIaz68Y+PFhAzFr//0WWndxLD+6YFHD1ECrNZSQNvmu+cdzFiw
WyOLFdeEkxP7TRaJD83pYqP1aPZxNCLUFTVCYmgluyXPor5JGnZAJIf/YR6+Ih4R
2PExKgRCKWKig5fDeHAd3reyDNad5BbmQAXL224CtxT3RGhiEhCzCrap9xvHdyry
NoiSfYcTVilTwTKVfqkT/lsEjINTZO3fGpMbubqK6z7FW5e3w1iCsft7ltf4GHqK
GW+zCNX3D0Y8mHzafSQ0Qdo9cnoX+7j7b0FGDyc9YDraPYnI5CU8P17HBRaS3ia/
a6p4RFJomaAtf1wu1mB7ETAc+SH8nWI1xEliUyY+kHHc9QSD4S5n6FVUMXf9lgXP
zESRfhNkHz0eX+YAP43ZsqFokiEc0k/q2cKQ8QdRQli+zyxIp5dNmxxiC0AgL+99
0h17vPoTKCSivim22IEwFwTBQ4Gjur0zWpYAmNxeAiSo/3/srNYGmzxjs9yyvBmI
oC4xgWHU8cwW0XXeGVnLTzYq+bOpiUDDNWyFHFTAwHRPBWAEFCv/hrLBvR5mqgoM
2vgKNrJ9Wjt6gQU2iDKrcpg9mL98iKsLzNBQXwysV3+7akXDrVuoGhmyA3SP2tyt
C2eq/VMIHPKkGEIJ03ms8/JnZTeavPEcGAUC1L+0k9fF6v5HIl2PtkKatfOo7hB/
98IACN0Vfi7t7Oq0Tpg1q8Q1eWvQOhLBM1Ug6qaKZg4k1QZcniIwOraJueUn7qDT
/XqIdMVLQ15fGBpZbS4LVNWnEigRa66uWUAfujxyfchYD1eMLqRNOEiXcS7RTwtO
NmbIFrT79Vczurbg+lkv6G81iVoKOyLclFpXiOyC4Y3oZezM39ALP/PgnJNvoGDE
BbRPfpDetdt+4c5RZH0cx/evHIH0t5MWTqhJjIQl3dXUk7p2y+BWIn1F+R5eLB4g
Zy7pByhyeSZwTyr5YujNuCUg3ke2SA4XnlfckofihfMyskd3hdnj/CdVdlORB+2n
mf+TjjWucfwdnKb8Ve0SRuwrnPUxG70VgQdv751XFWohxTOrkKBuurNwDdk1KVdd
OxXOfwD1HwWbXDtasnIb/akWRZhwSTtpx+Idb0xJ+zJqL8ZQ+qkIwewTTtvLL26S
76zNleAMxo70PdpjlIN97ExJJRMxjODR5zfK7O9rK0qr/rhpBrGnYQXEj8VdOd7I
Pm5+u/Qm/b4axLrzjYmKD/T2kO1+5ukD+0ze5/yHUtBwqRHWxsb0T8nHSWINPnqN
nNnFtSwvAQKkEgyHMCj8N2ZJQzf77nujjESIku42k33Qjd768QJEMCwiKwUrXjbo
IEUIPL7N0ANhJCXTcuB0HP3hZNQdCtQeBwv8172+dY3pjvwX4yKYVI74/7SqF77r
rFVt7Z6hmfwRW5trKzhP86A+lKaEepIQBE2/HGf0FBa4nD0gwPLSJJXdBTzlfbQO
ZpZylQYNyJib9/FEBzs2x0W6dhwACknyEznMoL0DE0doGdWOVcSfL1qITj+uLnuG
96YAWBN7K6ikSmSGBZ7OCiaJwswRHbnn1y90AnJNM1iXd2L+d8wdOGLnwajSKAdW
ehENFuOY31DaaPGA1wUxakoysGmaWBWFOGu7PqmRdkBXecGE0rdBXUFsOyZFpMTv
3UDSwt7Qa4SpgqNwIbvnuNUVxcgwkQ1SGE9riXdSfcg1qazbzW3Q7ShALzjdLrsR
wDiW2sQuucqbbvwHzGUc2D70Dx6A45pMWL9wSzDW28sU6IBTLLqUWNBv8NQOmnoG
R+RaqILS6BxwfW3fZoQ2ljawwpm/CDkN127GvikVd5xgsbnj1ymOcB/pZKKsQ0nv
brL7V4CgEV3VPzuyMy0KP98b3kt/U405dLoHR59VVD8qTY0Ctf3BVSzvPTejsRUL
U6f46l+L/3janlT976WoPW+JR8nY7lEalAp2paUAY6w8AF7+gRRqsOjwFRBsKpPQ
rHrbFen3fdziM6ZfIiDvjEI5VZhIIC1MF31ptVF4geKvmEq5fB5V6x0/AZfTw4jC
qxrmNfFWxrFzIwcQde4P5DzWdfL+JZtYiwm7LBP1Y0u/LltiCEDQlzcM172rJE3n
AyNi9+HrhF4k0ylyVGPuBUlt9eCaRmN9WwBlqOIV+gsTyKR7ZZQPmbfIveVF5FVz
hpMa9vL2lfNwpL6fg+h+zYwuQ3l7velmq6Hs4qkdxXbdgllucxvktXAH3enQCCmx
szENvrA79oCI6At/4rhzIaxTpwoo7rkOcwm9wLa6qxIDrVTo4O91WiIyrW0OZ8tR
daAbeitUwQX+OyTHv6KEYAKxWOeeXiwwDCiLSHwgx8Na12VqzRWWPrWVNwNUbYOr
OIqoL0lqEHsTHz0RWkVPKXJIxIb6vnRp5M95bIb5yJh1+w1R1mT47ppGep26IOej
PbZuI45iUhkIbwL2ZrYV/xKRUqfNQKIypcmBaX5ddmVGuw7MYtUwWGng5S1JBrwj
iDtcsYA1kJIn13taLRA1V7n47rf4pNyZRkCpQZA86dmeOio75WfjoPV7l9qC7zFG
wOS3WPgQKWBFvx7MmmJsfEAhr/fbC0blx18xmZLWbmet+661voS/dCB0RqpUPFiF
kaf2718bWCgO44TTrJb0x2Ehd86FzRYF9ZHRXcbtTh7JgG4pIWASaw5ZOuODPAgU
oXXKYc+Pg4St9wxRrBgoDEgTUe2RpdhQd9CocFq3uSv72x+uYjOptaHawrpEhTyr
MdC4w5b+GOfS1n4l6bqVjQFRunW5L03xtp7Ml2hoY9mRbjMkOIp1Cp7E0AhxNJgX
DWGuVlCI118joHYSydXjUJv0MTM3OcAHL/iTzWiDm1FVGftY9SQLvq8B3z2qVo05
Wk9zl3KF4DtYsWDXTSohL1vPLOv4WqabJbp6vts2ccXG3lvkWQRCqm8oSmaHupJC
P/zwKj0Kl97HiRkPzViU8E30SggR8kkC4Db9XWSkQuxa3xQjZnEaztoJkuxa6NNR
cTRLT8rfl+Dcv9kcQfLeK7Z9lylY5RfYkIhKOOvndpEVD0HzAt38lySqIvX59C8n
jnv/ru9FfbCMdfUd/K9g9ByvdAraaRUOyUg18x3nehOljpPjLy75sN1ppg2G8BUA
awd0zmX5MrahLLU7ACGlkTKDV0nwK/g561JO8qYdB51aHBT81iNYzYFADunLt/BZ
glbDsCsYDOmk1nxmLS0xT2w9oaogzO1ZT6wY0Gd3fPQyxeZX65CbvmuYN7eBU/Wc
an0yDcQBO6VqZTWnCy4Ocu7N+ftnfYFDZBRXseqJFJlmfDPYf61MvJgKQhHcqf46
aB99Ol3cZ/H1aKij9MI2VbIcu98ScjZLGQgP2hhrX1SBdoIFL9B9NVeEK56zGArI
SJF5qtwnMbw9RW4coPe9KtRoaNgOa2czQDJHWZ3Xvk/oei+YXnsgmlfFwi5o/7BA
f3Za94UZHqbYejw7w0IF9lJ0S36bOjpz1lJWmdWYSkMUef/wKiAXWSLR3AU3hXq9
23TsmSSU3RvbttqZ/YuOjryf5CaNJQnFWiulFVFIQdawIG5Qh1A+257m3epoo1zJ
jgbKVsQ9NoM68MnNTTaC7CIlg0mFau3/LSq+9yNqY36uLw5+PqN2WXPrvuQdmw9S
fegfWd4gYfF8+UCETorXGs8c9bv2TjkjoUKA8NunjEjzHwRQY9CJzhqtaALHSCL5
ixb6vyYoMLzIoEufsSRQaioULVuUECoGVRxjdOlXkQXgAFWSuBvZug8vu8+DXMww
qrgGxX/JZNMCs2+42OwWrrEdGaX3TVu5J5/lrERvug+XXfiGzFIuhv2hlwSFdYyF
YKPcu/1O0tRZA1ol6Svur0sS49eb4Fcuw0d+ICFbCRjxDVMpFGHocguHHQXz/gOT
/jPjXBbjZmLG9aQn1Ypd2xVfIeELA4SOdv586dbykKZaZTNTNEO5a4qwYs5SaO9o
0QeXiqCmj8BbVj8Ptka55P2n8i07eenrPS/EqqeEbcg+zY5Vyq57AYOGZRNAK98p
801/eB26UewjDyUfV4vtn7ZGAtKH2hjdnST0xe/9aouBEgwqOfA1EGEtzyXpfwKt
rKZB/Nq9Ar3/2N8buV9agx8/2BTObwxDls5S9Xw9GyIo7qXlNGQeUZrfaSAPP4y5
XuGAsqSUhkY7g1j//rUlE1Fkya2nE5l7MOKu6vkCwkcdK5sN8biOuYhF3tgWQ9rB
WVxRiyGv1jV/rsHdI04Q0pW7UfI7S5fmWViS9vWzqMpKrl6bVoSeaPtAf3McTM73
tvjYmeb/eyMDv/O+oe4SV9uNzjWdrbYxBAKDatSTS4mHYnxRqoUMHEKtv3+9V/PL
dFY+/7/lSFOc2vx6aZYj9M2OEHoxVaDHHmD0SS3R9TyHFm2jrjWUMPo7ovRzuRTC
vLbzsPUpBuBWkAUjWdt9DRkMLLXDs+9px8jHjWQR67gfwiSdiSiZlyQbCq/PADvW
SidgcIn2zEbGCkZ+62BCy2GSadjGEPUmFj70HD3Sthpqwygx9esfkLydK7NhbFo9
mEc6aFuoDjjb2hRGSU3HiLbV9AjieAeehruFQY6KBdv1BFFcKB5n2inlMXzkB+8U
FHZOa7xQLnL75o0gQFthRv88RmttzvU8USYHlXqhM3H6mfZV3vM1x9mKGYH2hgvR
AFUfsjdtGXNiY8ta9z2w0Si4UQZMl/rgA4O8XIkazc3Wakze1p2wmkpvzjT3XTid
GX4vEMqxA72Q2RuIbbkFQX7zRGmkQ7K9dEvz7fNz8xAD3HCKgd9zHGLioXV5Pj7T
qxwWh5rcctaQ9npPesVPE2UHiiTD4ixAduJ3N3dgPfUq0+oTm40UbLOkwXoDfaer
J6uRTNCodiLnM6VXzbVwwjix0Yjpows4sNNYJaq/0oaaKeybjtKWEkqfpRR/qAgu
byFDJSbLjXhZjuLnkM88nxPkY2BC/6Q6SZUQxp1Kf8Kv2aO4scuLT+LTNjkpBWpw
F1+yf8CVQg2/MaNUnFJ/6CLyNA35UmuRi6JA+mK4oBsN/4qjdiTIjUgmCE6U2BL9
rPXSx2kxyrDHvZE5vDsK1pX+Mn5vqpG44MjqUs9c7NubLPZP/3szQZfTkVqd16Qw
qB0L2QhlkCtMBOIKeDauUIOOCivvOjKHFm18yk44XKfqzYJs7eDiTrt9hqNEOam1
c6wGmsagoqcLxVyFxcSjHtUizoDvU+/dj0P0qMZyM0ZIOc3tbSAtYr246kWSsqR2
oB2NOlLlkxXWFIQoIAwVNBK6fT2GOkqeNGsIyjnV5EuvspUl/ePauz8YNgG4nLVC
kbyUXiBwvzz9cbcEDn8kFpGIVe12aKeqSl/RkHEr9bgymWA3OZh7Owm0bdtuutvK
bei/9EWjFKrvwZbf9S/sCyXItaPtWTcTg6WxEKJHCw0z8GTS/9lu1vMx4GxNnxNU
hPeJGMiZwKexhxeE4nYlE9g+C6xUi2Ty3tfW8s7DilNy5E25cJG9qvrcqF0BUURh
qDKVJyYlCYrQNQ48UZe07h5CiI+RL3uU0w+kuGqFhYXY44aO5HpLmDC/0AM9xDVr
gdFYYPJo5MNB4rh5u0yDlpQ3MBNmMzqBsvLu1iTFQIa6NQBmlPPxlqN9Ve63v2qw
+inadjzCDCT6lvCOftf8FgQIh+BJZuOiCz6uS/VeqJpHoLizAS0lJ/3zJ50V3sdf
eYOTYfYZIcZTqx45tkuJm2PvkijohbyORtPGCz1+WYi+KmiqHA6qeyUT1Rb2hTrR
CFw+FVo11BmGNGDh6GXwib0EcxIIQFFphP1A0avTl1kEa6tS5osTCSGoAomQCNfx
YiqZ4rBRoERibDL59rD1ovZqUHrrAO52WiauiibAJiZNCtExuaKK2zgy4YTlPneK
V/JMXq4qnY/b6VpM6ZoxsM9LDv4plNz3mTQKyHw+DM3uohzC+KV2tLMECJRP10y4
xuh4O3K45dX4wMUboiNtlHIRtvjQaoKrKYMTxi5uyX/q+YsBV0f7jSgXv0HMECFA
kj8laTG3N9RvFKzj9U7AtQhyQOPo1ryzcHrttJb/TrQ5r7eSdJjx4lyDhW0pBC6n
up4SHjkSQPg89mZa+NtZYnTBz9U8DZXh+/cPY3T3a8tyjAULRZ6PKpk/ytQSVXIP
Fd3kqXKvVmc2QIIK5LFiVFwoSYFyxAdd6GpQCxm8XZVkCRlWyBCFI3ENxmnMYhuN
pD8gcCc48v0iRqKQcw/xJJNI2xfkhV0SxJui2UKY3alksOBtCbF6z7U2b7DYVwnm
DmBlWymJ1dGbnl1AuNdVBUfVjPEz8JHH3n0mhki+lVO/459u2A0MEWKbkSdGUzza
nyDd7I+e+XoRxhjU5skPz27Q4WSFvybrjfVjZOBwwPP8PnfWu1QZ6ISpa44kKo71
Z3drQVJY70DeeSV2lTgNKRPLUy94n1TiXiHq3AoDwVBTX7BDlkdITi+MTSkhSxZW
K6mI/2FU3EbCp+rOmj/CGYYGqxm7RN4SKMfHO2l7MI3wGrIwUZmSxIooHAnPSp9d
jWrrWrxTwYjetmm/eFig5WFMeUsU7XLZZIPB4T+oRvs2SkUpKgg2zhuIkZBnmTPF
WTYXSOLgmjO7Ay3J69ycLe5Nc1UH/+P5+tGUVhRowOBaA4ZDgKp0ptSwGdT03qWd
q2Webuu3lajW5oHV6Pb0RHlIoVPSG6gViwiNcQbp6G+qZWg5SCYa2rnHVmRyciLe
cD2D9qjMtREa6CQ0agFlm79yYXWiLdBBx/OHPILGRPt9qBIfR6aDpTYPF5F97NNr
n+G2fgpfP6Wiy/sJtTY/0WPj2fiFJPw3jpT0/iqf3N/iEETVq81VTIcPpBmmK4La
h4LJgldtbwK4THJ+nd5jAkykxLdG8rbkig13OpeUmGy/VLD+nIJ3jvdoq6fVznlU
IkBJ0jbTFHnwY7iYUzaOce3V2FfJ4EaRTMCFraV32FuFY9uxrNXpOlBbUWSZrcn+
2CKm6pLnXxTMwJ+EjLOm6OsrivVzXomJwJcMzoVg68/IlD8NC8feb3O/9rTe7aAa
OKYG9/HEiy4CaTqpWGxAbu+jMIj+ScJlkIpokeLULNEuwyfloFXLqav4ffftkZd1
VHV2iMsVQ/wxazPwzTRlVyVPPF1P7i+uZnE9BaIbSBOtfsZzSpdxvRKCoINADjFu
ErRLPzoz8LMOO3XbwUTKOPqKDTZkDY/QgDbs76z6sKLRrpD+Vp62WZCcCCUBU3/Z
3sqKPiRz86OF20VASHISVx7EMG7Xwnj/37r9v86c0NVNOXlguehCPLyOh/vTEsMr
1jcgYlbGK9rIIGPJiTZ1/hGjB0ixepOz+/r+v23kvESGOEr/hjOw5Mduby/o3xXS
ifrzhdrG95UdpXmq6CgpmtAZ3mLS77c+Tq+3GEuASZSTpmqmH6+rtUPVQy95zSOY
1x/8KoRbY7Oob/AsY1t8rlc9d/cPPrgQ4c6IFVhIwMer+//HlWpZ6SUIYBF/O/hk
+JOjKREs645nS5pfHQRfV3mjKMkun/uWY9BBjBL5bj/6k54ODDQ3WNDmih+0k8Em
MufCg6D8sMcm8wUP6qpQPkqWtCKGjEdRBLYBbyypWnT9jgxQymgNsn9HKSaRd0A3
mQJESUKQIP2UOn1CsxcLGmwTN/U2ZVNlA1gj/VaF66j5r7BKRmtMJb5OCDfE4Lmi
mK9cZXUNnElmytawks3TLbIMEESnquB/Bex3TCTnafi9FicZIiqaFFJXvnpR2Mpt
1gZSj/caYEw3gzTtfiVEDhkfNqj1gDPlIvqw04S0074DENrrntHbW1lO9wjBSaWn
rhpteG5b3xK3e82vxYJV/kJFsSRel8u/NdfBh+y4zSgoS+joWgzYFpu51aCc4N9m
mzFQvd7VKFL4cGf9d1Gd7ChOdEDCkEO3jrcyhz0/90h00eBCtQu6FtMp5ZWHnNqE
z77+pyzpr5koGDU5GxD9zLppSkNTaY6b9HqOTJXGBt93x83O92Rx6+mdZmhdKVuM
w0aBIiyDkiBPUKkOERJety7Jxtcaplo3C6TQITlEIpyxrW+ZK+Wjfnp89hU0hvF7
jaCqJPuBYS64tYlczXzj5H0x2lGm9kmX5dhobX5wptbSV6aOadWEMrglYoNBRhx6
JvMo/Ov9M8aG0E959yVCuClrrmhEkjOcKIN3DTHxy12GyaM/j022Grhh8gmquUHh
1Y8mzuQUlRO54jXVEukJ1r2dSy5HG2RVP/TrYQsFu2Ilmach8hNiXZ1eBdBc9IVs
PmOchR6kUkFJTfhcR7EPYaKkJNFUml6oDZ5jQex9RWkOxPCs3lSFDNedOU1YqwOk
+g9FXYVt5n0Ms6fliNgag1MhX3B7q6/7MOWfRI3PNN4/G4zmwh9Jw6etUBXE3yrO
9zEUgZx5zv3iarjHRp7zK6PFWEWcrlkS25Lzl2sl9kIOkbSC7fBENbIb562RAGL+
rfzykC3rRVpSLSxjbGQElVbtwnytM52AeaY4zefqdBobM+HoBiGcH3hPvBAQKaxP
rZ+cVaSx09V3m5WMpJzAIVOlH97he0K/B/L/uLBNhtPlU+77udJm7nhiQkDOVYrG
Ru9LUh+2wbHZHPyJx55oOXEvALbG5RQhcUSXlLnhGcJmk2Fl0b4ehcnAzuHBZii/
V/bPTHL4iQB6ipEi0lSv0FEi6tgHVKKe+GsEy0wcsMA0aoki7aYKWlHJzfuUTUEp
FPbm55iVEVreRxC1VvsbssFCQnlBD7mX+TrBVw82WtDFUdRdJDMRmcD4/IAET4Kj
o+zUAKFjt/O19NrwM9FY1vQph/FTxKyD5bBbsef1WXPUvloHMqO7VAQyQs9jS3eB
1xr+VcL6qNfif5Xbq7IXeOVBnQBODkXVHGOgMsaIpAb7FZ/MO25BUaYjJNTS/0UK
KWdJxYBnfZjcultxehrR33By3KeQkkHSfNQQ+n3FuzakxbfQ1cGF5SBq56rXZU3D
In7V6nS4TdNEU3mt7ylpDeLEx/LyVT717g+KS1Pca4oIMsOOFT/L/l8NdkAhciQo
hXZj0MW4iMhjp/zmfM42CGwhviMJ2xc/N3+EnsfUjjU/t7SlL/PTmCnYxS3jQFPV
0O5fsjSchETJV6RQChYwoTF8LMcsNEOodHQ66F9K8Ucqg8rEBb6pFSgfKB4/rg0X
KH2dKFuVbSxMtA97JdFMCI/Aa/JJ3Ft1edWMCtQkbfr1eCnkEha4nuQczDcBJ8De
Nh8GNwljkijdcRUWKRdpD2g3tDJ2siTia6ywNEAlJsF5/EyHjotylyAR166NLY2G
vs9Q0Edhs97vZObdsHU1XQZYqFflOM+pwXPuhjxJ9gKDEqpthtdrGAKwkpBK743v
U70p3ef2I30Lz/mXG7PZk0Ye7TrKYf5Ypqfwo9T3pLp2zfTxaC1WArS4fxpRm0ka
TtdTaClRA79aieIWSxCMvYZssmVSlz/VhPyxwXiZ2tJutXygT7rDoqSRDZNI/8cu
mmsp1cev+WY5Ch4Lu6i41liKabd/ztqlFxqXeEnYizNoFou5tasd/9eq0nL6G6tB
relvq5xKPOVFxGj2IUZ4yacm4ScyWljwOmkRGH8enViM7OnN05VVzuCSV+LKIvAH
+tm1YWEpWl+ogQf2mkMF91rlt7W56J65qk/vZ7w9e3W9+z/4Rh0DvjYUOaFqRoLc
AxTkAVWvPNuybP5qx5XOYELR2gglXp5Y6J4FQqs0SDcql0uy4/35mLNZTt2LWGxj
sefsgFmkoBw+2o6OpsFIGcraKZ1VGx7tInNpoHHuUP9b9NCIYvAGCeMIeHJw5ymb
agS4F+1Ca56KNLr6ErilhnzBdEpWabCMI6wGGnykzjl7vUtqx+rPOldHSAKf6Vrz
f3PS9Z8rEJWC1GHcPB3ePqi2Ubwxo310MxC1eU7Dnhrk97N6KA7zmH0j0olvw5Mg
Kqg6mXEpPkk4zUI5hese43jh2ikAecZyY5941akb+HYoM/y8r5/QIAXnONMJ7tAs
4I7IzfSEwidNoovlhmptfK+tGMIo1T5p285EFG28kDHBb1seKR8/QreQIBXLAAUF
z0E9B4A+FtaE0kt8ZZRO0qhEwspCSLmlW1nBzMGPZfkkfPP7Ni5/x45LxjAdbG6S
b3j7zY5kH9+nIEkNWbinhgnkwnulS+WXqD7KYVAQcM8u2LHCAGoB0DMPUU4cEeqe
+HXrLllrnnb+tO/YApQmfK1i/AITUHilUZo6obKqNb69VutRNBs04Cv2ocU7umoz
W07SbaWQn0+kCLmxXIfDEGLCHVvQ8VTxdvUbR3IEVfLZ58lBZnIrNtOGiGA5RWnw
8eGs9m7vYPXheH5KCOUazaOnF2vh3c/WsWykEjImRF4tTsICkwZMZ8GKMMfN9Bfc
bL7959hA3kmDUqBCfSoF9ih45I7/YQOa6vjplM/YJcoMmtAZMsLrarHZuXhI0Zjh
cD4L3uMrgOuOUTKpjlKVbUrBMQXyeVXjS8WF3/+FqAKS5vX/oNRQUAleaUwmIYDO
T9M61q2aczXyhh/EzJRXuOlFyNvVr2slHbUtBi9xt7ZjQjUxWWYACqiWfFrPAyrk
o1kwFn//r0uAjPfqHpLeVPom1utdLCMdatmTkNv340IunbCozAQRCg0DSigV3r6+
PM0twhS8y96xT3jBnyvohK/c/eGx3KGvVCIw1/ICY1SO5DXFpCeBszn70SC6xudt
aGpOBRuDjZVqGNEy8Izf146T1QRrm6hLG1ISo/RxUEI3XTjgio3JAd1/HFaL5AZV
OrSPOCcJFm97BPw7gmB93deKjFLolsIi8dupHiRv+S0ZL3HKvSEMdw2x6vWlsN7O
DWzj1B2rMKbHkG1HLo4q4JwTVoLE6VWhqWEmEbGVAUB5+Ug9EVhY9/H3jSoUTFg0
XfWHPnoQcvKD7QtLwbrQkyDwiBiWyNj6O8FAYDJlQ1Z/i8fy4mqMco7HB2Pg8mf3
QdeElPsgl74iievryJQFcldV/cqingWuENHHGF05TgSuB3og5YsnDEPxH8goxvgW
zo6LaaARIZ+vuYClftogWI+f3tF9F/Z76o2Azm7CCDj9zQI4SMkMTfssdlH+rUxO
E2t+N7kVC26xlGIX5FcSi2bwAJMi8YL3MV34qb04qH8KfgT77nmxyG1/7Rw+dtKe
03BEMbjljbRCpZ/Q7NeFCod2C7Z5S1RjCC+EgZ6VzYDEh1xzqCzUb1QqlPdYUPwI
NdwTyRrelcmRRoSL8zPulLgRFZMHg2aGixe0uCObpqqq2lSHHBc83T+RNRmGPUZ6
KZuTGE9z15nhbEvBvpxsDmQ42AW2lVvxdPDyfyyUkhoSobvYk+DJgIO+YSpBemjL
xbAlTa07KOVOO/7llH/Zcr7k9Nspm0YBwEgIl8oVMbpJ7HvX8M1ylihb9znqT45Y
07rv+LN4TmAwOxjiguF5Iv5qDZM4T1k6ARxr9su9vYGQd2cGYBi0e9HYG6+6tjS0
rgEOlt6vQQsKV2GcXfiJmrJAsobfLrkEZYTUpgHEXm2gNaQw0tjsO/dmuxz40i0B
eT2IKsWxFgkcVbj0ef978ury10LJpKVIo+KuplJx1yoEoenXzwOdZtFhN3rC3p5a
BO55pV3MHGeEN1Yw1pcyHVekONA/UZJunTrOo3N7VqtNnat/3luX0Z/DHN5ZZLT/
eAGzAWnvyoEHVB1A1w7dsRH71Gtjk8XNA9nbblByigyDCMMg6ntUvVBjWLNxGfUA
N5VY2yOyMrVZ9CkwryWDtOUBZZoCRxlxD8HdPKYVxuHIN+cm3KOHqb0yHqmCxLM5
rDUsudfD2jaExHWk5D1bQW1EUDbtYCDdN27KwfKABZbecKUV2Yz71nyCV3d4xsxE
70HYj/vi+QOiYZJWBC6tvTKu+yMPL8TDIsb9rpC49CuXNE/B7IlHikPXHXh28rMJ
AtmXRGrzRtJTdRA2zw0JbanJwAAKtB805u/yYt12fN6QKcEcjS6Glup/WFfJaNql
pEGswWEVC40VgDHEwS6ikmfnunNxgpH5p0RUlIyTxeoqKWikUvfjq6Iw0FUQN6Rw
m41tonDlEapWbriHEAH7AXR9+mUdPx/ymy9mJ2TlsFw1Indzbq1jDh2CUYxJgt2U
YuHwCPtwMviqQvOHZrGLU0t28t3tn6Q9gKiHHA+nSjmuPNtDlT43o/5VybLLimki
XoG7bYDwgkamWAFQQ7uHH5aVE+5iGU2OqgyxrO4DnxIllZENC0qpQGY1WTETzwH6
qBAKi0VnIIbu+SpRSTb9pD+U0YjzhAopBqJgzQFRtUzo6ygBACe2p5+XV4hXh3Wk
St/2fKRSrh+bFkuA4b+j4MPRIuX6bGuhLta00yKRpXgZowzU2chEIcqJZ6vuUI/t
lVh4Sx6KDU8LPvETXOiLL30+eIGX3NFYuUz2xnnQro5fUmR4lzHtgtcMIKV30eXK
kCZK/QtdoYuqRCW4ZD9LE6d/P8AtDyf5yEL6qcit2R3EOMW1aC2AbD7unIBmpD2p
8RIv2Ypamf2ojDFOk7b304dk7YplJ7q0UGnAxln5288drWqANSlESkGw7DJ4cne8
SZ/gc0fLXxkn1a0rPWA0884/FmZFmtTpZXvM1mskjyuQh6OGIYGJ7l1dbo8WD2zT
0VyerxH3Xfdl2BIgvD1ss9LuKnn0T1wkhPicTHY1iPAy0IM2lrUzbVkAvd4p80Xn
5Z9JJo38dqnz2Qz6FUHZui9hTH3zGwABRzLq6/+saSr/z6lp2uqizrpwpIZZE+Zq
toNA0r16kGQjfharC15ou3Suu81etBFzIXRHkYGIjGFM3AtD8uPWXOInQhVOA7xt
2PCzV1Fo9/DDJ7uBr8N35w7GH3copiKklIfE0xR5Se479QM7zwMgbiExA8oaF7bX
tMd1/UBtq16xLNE9M/+ZjOuT80HVQ/1u+wye8gqzELBAKjS+TJTl4Ci/17EdkJ5k
NN56YhBwlgWw1FRjQfA51LMPO1Cf4UHGDATkwG27yGZlhDrh3ztNFltPzchfsnUt
jBmWHTFOpVSpSULKiCGM6Nh73EnKb25Hk/DPjRxt+XHTbgxYzyc4CIY7ZI/6KnFr
5vg+RknGkBslcdcxPmhR9YwwGWWeShlCzPa0sRizEpkG/vvQtKFrjasCJk+rGqRt
awXqHqdpZfmOP0FLRL2wbUMjdB+WC+bg0EbxC4JlGmDV0NJMPbwRr9mvN6CNIPb1
leoUWwa6xpgnToFsCDIdW0O3DPsmFjc+NYkZY89UO9cIjEZxUXRVy3QYhzm6FUGI
vN+wmYBeYm2QsLmZZI6PSZpEecwJowj+YwhcHD/MrgCtbPX7OtSX7iVULQlISt34
icqV4Lr/7JlL5QcsTGs8KtT8F2vQCO5TKVmJlJ9TrLAgfF5x8MhXy3LlFsM8+ni/
Vi5aiJ57OPuTqBTgaW0mEgv2cIK0oPd8tIM+sUIsbZFRMWi/2IEyziRXYPnpKYQD
4PNMLu6DBcJ60UAaAmbNcWstDoqOwlROfIApQdqM4dMXM6e1uhf7ZK+CjtOmJk0v
ItiE1ncvMlSmb6x6UxyjEoOV+Sj2oZrxIyBjWT1kg8XS11zkska6+PA6oqmku2Sp
RsuJ0M6v+oocKFi2auxpfa7nCxBpxYNVSPrEuElLKGeQyUr6gSNQOTXF5ifvq/Xs
nt/V9m2OmCS3HSRXlGyvKCE7OTp/MshlSy3BvwuhYaKrkkDz7UIAqrndwDB42fGb
yUamOaTXBylIReZqN8OhgwW84Zv9ZlUTJx0evZpi/Y6NRoC8LzD1nBlirPSf+x0r
LRhenjmqz+pfxDn/JQZJXTf+udpKNf34IEsNtjNrBe4gjbNvxrXHcnpHkPdKwz3F
01NKsBIy3jD664nllnrtWFXIrz/P3dkMgpT1asJW9dpw48U4Jbtvy9YvlNUUDcRe
X2+eS3jzN/xxv25KWmnxCaurnItpPxb3TAw5K3t/V01uyD9ezGGG4IXPfXdT3oHo
5T8Ir6fwWFmBL/fboyUqBCiNQpTHX45TttmLG7HwZvv1opUHr61fyKt5MXMLGuje
/FWvVfdO5LIjBklJnemDFAJBDlpVMFd+7wGVzwGXP1hQQYAkyTC4VQiTAt+2mA2A
mQrFvD1m5HjPGfelEIvqceYrA8GOYGT+S1cjQwPccQgA+cWGlD4jEjhro5qYTLrk
0vUW4yZIEvKGbWl8iN7sjk5aoCczw1ovRPRNtW3FFeI2LKjnOlKZx3S8451vtsHv
aNZ2JGqhJ0Q99rK+I9xnvJlZSm5QdSP0fYfWHBQac0FlhzoOviwESdlBFOPJpL4c
W4dvJmVkPOiZBhL2Jwxdx5H+f6K7+Mkr8JTZXAZrFSmQyX84dp3OpQHFwk8NboY4
utSlOb4VpgL16uDL+3gLfzHlL2DSZhGUVARR8HCHHsD/MZU7Hn9Zbj7oRaF+BbyX
5RNPv7snlsmwz9CDGl4y9sUhV3pIXe6mCbrqlbXBfiTFN9vkAggdP13kQHwek0Ae
P0rGvcyx9vsKRxHzLljJtnpHy9j7JyC/Pwv4uz4MpoMfwgRnGcsJiy65hrRPr8aK
vhq+aeha+1iofKs5s0+PkzLbX7leil2RpL+nEFFVn6z7O7Mr2k6eof05Qca8r3UQ
zRAbOvXch1GVEnEZG8ZRS2PA0iGPD34cfQIZTL7/yehGq42kr5n3cXYj7um/4yu/
kdFzYFoYEQfGRZSo2kuiVfktEZ2eW98K0g1kc8zu58KgDhmD5spq+PGDuA3eum09
z6vQR0luonJMV5fVKglFWqA6MVnQGDA8UopMIGSDDkytQGxHwPKJLWj4QxIEOokO
R27WT1QnUVfykCmOIY6g6FDJeqWcxeX2znElZAHwK+YxPv08nLT3UY04VL6mw7/V
eSHzPy1xg9Au8fVxhkcOXDQeFRr9SXva94AuPyXMZaozpCxZxKBuJuLt2Jdj0vIW
FMzvCVAcPY38pjWkfdxZJLC/tU9slGR9oXIUnUfxj149JBZvpTRecxRXfiJY+spo
uRFNequEXYpmCk05Tw7nT0209DR3xoBdNSifqo506WPMj0AjypOLaSZ0WRzjdcO7
8AKmxkzo8IGFLc4LyIw9FKGORBZ3WHreholaSMUtyYGhLKHsXHJLg0SrX8z8rdlg
/HjP/upZCCdjp9qRvO+Y/Tl7IHJFq8HXVeevSQHrn2jUgDrQzdFgqgES/LK7aC5J
YF1xSSRKVg9lyfGTuEuZyDOQE5fReBoW9l+6BSOwdVWfFb8/smBNXh9bRfr03uUi
zJ26sNGhUVs8Un+Sixn8iKVtTqELThrC2m0PuST6aw8BtftK/ASfog/TrkpUBpnN
hxOaWvNicTWZVDYyqXI0ubY9mc2CAs/A7xWkZjWfpfl+08w2s1DL2LPas7yl103F
OGWrmTHEZptYooDdaIsvmuWyi/8YF9yVPwlEYgX//YcqVYZKTde9rvoRdGLSVVYM
HmLea7Q4i9Rk526dyPbwYNFpi6MAM/sb4j9n+qkTpPNfVvttfDct+7/OF83XbF6I
ZA4GODUWqH7MbAOVOb8ppUNBptvw+wiYT3UtJTAWexCEBUKjTQLyjx4nO4K/fiAJ
XfOaj3y3boqbePuohlzC96yJtila50DzdOPwn2ijt8+A01RZuWYqZj+i1QW4Jg+3
bf9XrRN8J8CBBeL/Q8dye67QkXnISWnZLfNnSUbr1uPeuhVTyeYeeUX8b+NwJOoV
vI/QUMmcbROmRYQ8V7u9osJpLzlI+2QSRBXqp/acAd5LgEvKRLDPL7ku/dJnhu15
pfopge/NJ6NWwYSGqlUy5YBN/czpMovxkeAmqneIjs9uh5/aG7pdd4xZaThxcfSW
Ph6GJzohFEM/VHo0pbbsVN38rGWRwzdRVOqurL+3oy2k5bepcVZOMXjVRi6Rbvhc
yyx7pZyABKH7zlyo3NzWygUWBQOyvqgeYb+737PWmwitbKRLr1PyYKn3yDauU3fs
80v7RMwe4tj5+SM5IcKxS/S4y503VmN58xBahsVyeWqCmUCH0YtByCl1KKCXZ4NR
aDVxprw/7/cY3Vki/nIhGTNYbr8Jkc5WVYlDStbiDu13AafL626a3kbNoggs5JUJ
15zdsUl3o1OvHk+wHXeUPW8BSawWMnN81SWqWjFDSGgMMw2gTLOHu1WXP10CR1tX
JSETARcTiy93upr+XmZGVAntOtbjodTnwes0t1vMx+RE1QscYVPkXKq9rmBbtwqr
plIHlF78YuG6GYK/moZCay1uJiUoVa8TwwYXkzguZqGtFtVCHfIWO1cz+c+HOaEB
g3J+hzPfdsEYdGkDXqk2J1xICG8eSOdOAIHC9ebMU6UrBnt4P43/ka2c2eiqYPyL
jwAYeCN4lWmm9jwR8H1qgk586VMjlahEv9RDmSD/8hJJNmDc4068a6Lc6BGdKhs+
kCa4uchT99bUAXZ1LAahrCMWpyF9vNk0kijvnU3GvDem+12hzsmJB0Jxsi7IwbLX
1qYU+pLfalmnm8gz3hvEDcYbeAgbGUJqJ7Cn1gwtQzb5vuv98U0e16U3KJMJztQB
Q8bD37YQAxEzM3BZBss0k9VcejzAND1YQON7mt1f8As6uA6t8wQ0+Mp4Sityt6ou
wY+NgrfQxk6pcZO8QCkgEAMnSnlBNrwnjzbxgO/jIeu2+EwrjthOYgWeZbsoSBBX
eu/1U5GMxuQJtv7R3tGk5MkJPnJTpzdWwLpn5b09OItk3Q9PWoyda3NpcxhFZKJj
DFR7DBocIb7tu+19sFYUi9Yo78YSMQx4FhHTnja7LYllYxIwpbM3lbzTpxuTu44u
l3v+SFr0t5Q+kGRwWDdExjSGXB4kW9e3VSMzcX1lIXFbroN/kf9IbWsmyDlpWiz3
BPovo7CrP+6vQQjSiLAWSobu9SreJvdV8cyao0JzujsHoOMtI/oXG+023Mp4Y+mT
EQQTysks0rhgZ92mhSBWS8VZBif7Xh3HuvTO8iaGeQc1QyJUq1MPUN6ODJaOR1hp
Wz8CmtOrjlSYofmDUcYbBA8SL7xcq5l4a8nZyK7J2Bkx3VCBY8XCfzMHUYz5aqWj
v816sOuCgmhTyYmY07RgZUC7YJWWt4MgEiZQYlOHUguA+WUW96FZDKnmtDXWE6wJ
bEkV0/DqB3gVR+aX+l1ubzoL2bAgTmvq5/omXE0FyAWcMKb9Yz1hJvQIbu72VzMP
cowY6D07NhOoSGLGBOq9mrjnZRTovEFyIvSDsuCOa6npNvk5LGcl1wp7+KBGdaBC
Qam4qe13E9i3Hn0728uxNJ9+VwuBQNcSfIMx2m35goQnli63od38u/tIk5gVKljt
KpaJWvbmPYrzdHd+9RDS1WFUGZA5TRi9SRDLWu2h4YE3EDAGT+2gEPVi96/bfefN
6T2ysvN1R+8FByKgXzi00gtXUovJVwMN9o9lVOkzMwT56wMFpPIPAX0oFBTjJdso
enNeW+1iQW49KKlNl5wChLjbaKp1MjzadV9VjRi8pIv42pVSncvncjj0y3MJpyBm
QWviRmc1YeZouzirn1R4LeG0GMu7wW7fOlVpQb/dLQ5UcYnPQkShLjcsUTwbwJOK
g/novLTMxnEYXXx/h0hOsrhHNel1SuBpHLF+Z8eSkmXTvQGPoI7BCrxHPrqZoIAZ
L2yY8IqiYJj/PGv391HSuMTxhYzd1a4BGyzSFgyFcJfBvzPWG3/l2nAWDTzIzc1d
UajMhOL+l3VQyAsYm8pfvomrfQTfifLv+Vhbu97afWnSMKjbomSOSigxgp1Aojsd
if6rYu8UtfUXO1+6YSoEoXT0RTyQNf76yvIJOTE5Bt6610wCzQD98Bkj0Kck7Mhy
XES8B2uR72cyB0kWQmz/o9pnkB8h7I5ZWmXdGhY6ftcVUMg6IFCZzJB4V+1BYLSk
2L3jFqQ5xuiI6go+TjfvnbMpFZ+6PkLnDxFlfNb5mgdSwaYXyk8LnE5vhdyP//mQ
c9N5pd28PF0I8cPL+PWFODx64b6INFIBASBjeIQj4A/PdiF1XZ7iqkUlBlL/yHw3
B59xGmzU1gxlwMpJwMNaN+pKBqXhNnOepr7zKPzzByjQCDY09QY864Fc5NVcPe61
cxOkf5YgBUStD5Q7swjToVg9vEc6dSonrM4sag8nXJgDOmU/ODdTVtxH1DvnRGE7
QsOmxdWzGQilxZBSbHO6HF58Bxh8BpNy8/DGuvbQi30OyPZCKN8RUhB+p9kbpb5q
+vN2BO0wau60WGBnKX/eEQDlPY0jYaW6861oFsi1HCUA3OhgIrd0FuRESbb0EpMr
tlX11apY5iRmkFw1m7d1GbgjaNYEwr9dtP13ZTMMiBgPw9ybvMfA4W4V9i8xHgKy
IwrdIeeHusMowzyDkQGMvfgZbCIBoTmQqEXl5xiW3ssNuOK+QUqb1p2w16r084W8
oZAXEKJmM4G/X0UcAkg22ERinsuZzMTktOPyHmkiabC3KoIMgseYC22Ns96R619l
byEhoE9VH9c93qFsQaXwjISuYZP9jVhOJ9LZuwtGhrT8T9sn0atjlSTZSRA0ihR5
KmYJgOTesaN5xK7rvbAa9X8p3Cbrp4vJXf3LMN/nPlNY7HXudFJQeZE6IqFMUDh1
vnZ9CP8paINDG+jr9z3S1yOSTqDnCk4s5PlYWSUgY7WXx3/RTTjcz7tjtjmr4xdw
XkZnr7gFOR5kBt2u2OiA+uuHb8VhgFvb+95ATsvf6S0zPy5FDqihnaGr6WvZfHkt
SWURcpCyy1gggZ6JwEtEPqjCNgbYVO+l1SWOl3Ielw7YQRsLtjSR3CVR64ZywrtR
z2H5X9GLbqrnYp56GAfU18j4SxNz2AM4eJfRIvwSwScw6PEZ/pfIg5yNTL4rKbNj
W4vZBqRS4D5hb60a7KhfmM/2nR13mCZwrKCq9QRm44trFBY/gyt72kHI2+OpUXFj
PZUdkPPUTnnOYvEivauUc9JsBtKFu8K80bG0cny3fimHsEsIxMqvozUXEtSFmnIR
Ca42qlMcMNz4QPwQWpWjDvuhrA4jvvCIA0Nqiz5DNbGSd3ZyrYIXj7ZR7Yi6KlAE
1LtRnrVyyJ8Dpg2Yy1fmvq+j7A0BclX1sNGmy8qhSpmq8bKktNYML0DnUe6QFiQ1
D/7S3prrIXO/lbr9YJFQWLb4CTE2takRofNdyIH4Qa3oyjW1pwomUe93GEJZicrA
J0YYKwaVAbiyl9F+l+gCK8XoubOLhaoG+bpm20QtHWOLQoy1W7WeIvDknuxY/ygm
dZoJThkyQDDNeuv3SR5a6aiPZLD1HcV9uoiZQ7YFAdsLjO3UuqnllRqxXDZFlC7f
gy8H7u3TDysh+GTpWmv7hbyYzY4qOL3kGYNTh0HLKuN67Vns8NFP6Pab0UuoHFeW
TuI/eIFNYA6n+7TX9Qf7JarVAaa72pYnZQjKQfhpT6rjucBcEUmlsTrH3kUkS3Mp
Z/odtteGFGuwOfBiGcGBkqDO6OYe1kH8u6FTB5hJ4Gn1gu76sX9K1n++zdyz9v9e
hBajBqfNs3++yUOs6GdZsYagvUNMz7SN0wJ7kHaFGioDb6HxF26wgie/2wLxt6Ji
Ax10dwsDLzJTbOHt9ddEJd1D8bBbW29F/JOvvTjxwsfC8xYWi3jLTkBqwohVNpw0
MarQKM+Lh8yNKUUJXodjYLuqo+N6hsOIcR3YAVsHli7XcrfgrCy7AWAmECyG7SB+
EXs1FVugrSAL3mi1KTdx2WHuL5XQijNZAs9Fl+Dv2ZWoRSiP/M1XRoZUMEJpyTMu
uGj72noLjBygH6F73rMgDiz1rfhFGtC8mBMPpfnJ729xbCsrN3qwcvkrIpJG5cxD
uFi+86g6+EGHXCd+2bcVefWFgg/FZywTDqLQYRr7IDxkcPHgoLYQqV8rTLJne47h
`pragma protect end_protected
