// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CrEigXf+FjWbSIvHZbog9tdGX+pPZNWD25aH7WBVLSojQQocSLEG/YQIXuWzAiSe
RNgaCyM5u0QJUyw52bVRrLIZzeOMeHpJ4g0hnEUYx0ijOTYoyFe9ahX4VJnwQ3Cz
6wk+MtzVIIa30Ar/Arro21b+HkP/6CyJp2P/16nqlUs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5456)
cnf+j+12k1i6M2Wy1HhuAOYBr+64blkNMwXpfD6SVhwBBlb7ioczOZAJZC75OlkS
doidcDDju6swb47/wHZlOykZgVNnrmCBCHfupYz62NMGcvgUNrBhrgy4ZFWKlknL
YFUm9PeH3G1QltKGQP0FIcMF9JchrK/fiHyOnNr4Kl5zwuDpG6txpa3sXLbmBOa+
IbWYzUBNKUDaT4Z8jdpW64naJySJGMIwMlBwYNSst6Zg1pO3h3l9ZD+T7krLVtJS
Jg1CiAJ2dXVp+HmTUdk3NR5G9gY27GdB08WLmFLobIZEOZbrIaYmuVTmuCbLuKMb
KL7+RO4gKH0B1tExL7nrGiej8r+/0UOY04ouS811zguKBDyNq94CDtaZ17ifulXA
00wtKLoNefqiNkZQ6IZIWbI3ZJoc9KcXi+nfVCePTb0Qght1RdRrH++bQ4sjkp+Q
Lkx8avMxtnzpvGX+JuMBGogBzyAcawpG3wSAzvJ/Ws34blyZHF9KhvZ4IhL1MBHO
GSAtXz3B9NKnC8rGn3S1H16AxyYCMA4AQrGZrkVYpykgRJWvC4vDfCm5p8Y107vV
th8CeQovTW4RBLSFBy3+PX3hxvspUNHi6kIFQrRWLgkUgIwz3VhG5PycfhtrGE6y
uVGh6QvyZJWIDvnD1qI0yiZJ4VwZo1GF35zxhMZE3SUzwKROS8xxprD+dfIfOz6p
jxrNGbDY78o1wTY2krMRPkilu0rptY0U91our2TgewGOt7GuBig2AsMvA4rBX6C2
WipmzrxDbMxtKG/Czu7OmRHmDEIl4Ui8d2AKmkPGKTgewt0SZZdGo2fWDW7qmqAQ
+uAGGF3pIedA7WFjfCeVnBI4fO/8zQpKJljKFMsmXfR9GWuVpZ2nFLT5UTeVAPOT
QQ1gcY9UPiE7F4/FPCudP+/3Q0QU+rqHFf4Ubhqz6WM1oWj/dZKxPCktIX+KF98E
TDD9/M6mKEcO68y0mpkh7SiAbWFiabBswDjobi42ywVs2H5N5RYFfjALxTQDyubG
q3lLoevjiDDMA7kl0PvPl3JQlnrANVeqQZLYe2LLzeRkQUALSdRgVgpvgacoUx8G
8tNshaRP2ZYWyYgdJ7bnLgbTkd2Z4o+dB2FVqbCse+fRtm4VTMvUKXeeETNVwsvo
g+XI+F1bNioeI+szQNw+gCdAkW+56OwMH2Lx96KSmgLg1FvDNksO4qvKY/CyoxP2
475iI+Fzztuzb645dS+rBoX+A1kNd91B2psqSY1LuO2DyWS/fKla9kBK7Jtbxelj
rGlnZK0uaAX9bX6z0yfZjkrsnZ0nDf/dbq+OaQk51pyfCOe5vbQOcloV5/y1jT61
s91WmAZ6hYiTs/jzGlUYm6BwyJQLkl4eN9c68h26sFuTeVesSSYMRz2goyt0qmXA
hG0A9rdb9D0ajB/xzl6tYOB2iD4VOPhnwNGUd4GgFjU+pznb/ru8AP1cHc0163Ll
evYJCnGulom2i7ttcMrawlSnzx8FdXVZ4bdmhkpoKVAjPsuGX6s3nYAorxUhWQfL
Z9WnxvvekT9k2VEQkvIHX0+nfCKVzx9PqfNdywNlLmzcr+S/G9vl5I9pUbUpQTBp
Gzv0CQdkHdhrcgkfd2osfX1vR2zVOnUtHsih8yPTqBQBvhHFYoCswecq9V7Gvg+3
m1rVOb4vhCEAMrcElP77YoaDrcjC+42CYrYSR3Bn86aLSUDx2zyb2gZIskgXWj5U
spXx3NBK4s6EtrxtW5HzmtE6jVHAWk6DX1DDkmex9DMJEJ9Da82yJUeKTUH31wZ5
SljTTI88+mo3RDi8oRd5gXvx7Z9H/Ke7VJJBNi7Fg+Dka1qksOsD9V4G1ISpGn46
ETtAZf9u5qKH2NxNCV6hXbWNjxhOSOywVAVLVezS12+uH3J0YZ5aIDkrRz2pHNGn
LE0Tv9TX7dwBxEbaaYHPsulWd5ZtI8SIg292wTmwE20NgMLFGFQljJwmrzxpiHqa
ZnZFUuijJPsgU6+iD1CPsZFWNaTdx564YF3YNjh8HiI5PmsqghQYXcFSEcSYe0cJ
i+y+jBFgzQIca9DDkSjQSJwE6PQVOkcWP6UlfxrwUCBoj+7UQdrrcet7n+Vcgcp6
tanTY/70yk9VzgaAB1sap8QSfR1vjXkPx+RILDW9TbtNAZsR1zPuy6IftakMCTir
w5HJ/VVRXWNNbyeSKohPfe/QmRN/l9f0XG1sSJSfnGxP41qCXG2HG2sploan3HLy
MbdYDqi6iw4PhgfGGEUg1eMpviGXoWUDbFoM4G0YCtZmKuglgEiCtzK6uxz/0mWS
BfAam3oSihsFxYfQ75CbGzUIJCF/YiqX2UFfdW4uL150Tt/hN3jy+6WQDlfuHIOn
E3S/gJ4unxqLC0jGY6xnDfZ+n0EPxSlDcRja+nkWx7mUqXW3Ac2KCXpCvkY/ATl6
k+5gob0Ca/5GPvnXUE/oH2T7Ye5pBcI3d7KBv0Zx4SuM6dIxDSwXNrHCWE+qMovH
2OcPXqPd7eC1fqYTa07ryi0vzH26O5vwJ8vk6/SRyM9yTP23WTxMRqEyizjsqe+o
vTDejE8TegaxhRj54uK54lQsO4Ump/qfhBpPgCaVHvlj1jBySq0xiJKjHlzWu1kR
32AI1Ud3M0p1DAmirHl672wlD8Q58iL/puRTP+9MvtFAfDniETyziCelwQtjm8hl
ySNwxnIVcvX4hMxoFi69PqOyzC3D0dTVhFsKobC0iueNrbvTbTBvX/lxhnjEnp6p
cFd1T+5PCGFrJyBMJEt5F5XlNpX3k3OvB2dGPAz170KTOmNPyMsY5eCF539LRQcw
MC4IAJfJqdXV+Lii8k39Er+lySK2VXbf6OFDb9EnM357FhXr+LyewKOuoki1LOab
cnhXVAcAKSPQWvzjuB5AEWRwQgtlx0+Z5xT7Zd1uhB9lR0eVsd2LP251IBt7anLr
cPFLPTZtGXjBAU+SiILeEFOgVmUbE82HufdWZtB5MVNJjXl0CszW+YyYc0PPqOli
tgHUtal9VbaZJVI5Ck0giL2RV5/ciT4dEnsiiHPWvUojB9SKnmWWBdB3MAn0Nl5l
ljr0a/KdF9iFH5pdhSgMROxPlYXlvlz2NbXJE0nZWgqe3I3QhHtUjhMDi8Ywfjl/
BzRmcu3EwwLpJ4O4FEAsloWGIUeUp1Dse9IUQ4/hevxKN7STyeXZKS/KEhU9OSbl
8P+UzsASU9Fk5yPisogi9sW3u6MsdtLZ0QBKr2kDwdeg1pdx3O8CY5dFimt1BesO
6uTGrNB7Z6+Z51Bhs1stsdlB0dvzG6ByddFXpKOez/AnRed30IFNnSsaKVboSR7/
eOXrtEgGAI2sCavNGOgWIaJ5Kgt4YUaeluD00b+1EmCZi6YIfaZYRbH5TyY6c+6o
GpEeOKOgcEFe73FSgwHpNnmtdR9dca0B5gclsqC/DAFp0iYP+njnGkAYpV5ZduQN
mh8YSnesdkzzIQVJgpqZNO8+RksPjamTSF6im2hPd3MbxLtwkz2BwaiLMrMgagD7
3RboIsq4miUaq745U81OvLy/X1BjXFNDPQN72TDzlEMfdaZUnpncvcmfb2A8wfEl
yIYpKfyGZ/kdP/sxlRbHS4Hzaotn3ws4zMPOL1fAAF9F71zjTzuEr0cqLxVW/PV2
7BZmJ4qaYMrZqmFXtpDeeepWMR7pdSDPyShmAZ8m3X/CkznnjbmGqCfX6rqU9QNx
aaIsnbds/BBprizQGacuQyk+hnboUM5QuqkaimaMCpvb8iEW/vB0WOIySZ3PfezT
cEM/ZbFT3y9ikWkqR3X5Obmeamy9GpVeE/jOB3+9XvkoL6eqWB0D/VwRTag1KxI+
O2s7dczSC0WYO33+x0eOyGkBAi2J1YAANxceZriq5r0rps5xnaH93ixaokkV3Khs
YsO6ad3mxW1AYmK9LlA/FkA1DLhlIn4MXi5g/WxgXocJw7w4ruTHHTb75TLMhFFP
4CbzFCwJAGmISdUclzV2NX3uTNyfAVucJ7ErCTU2mi7+FnQ4ZH0sjRhSYhZs0/y8
NMDM5dcQCiE3+qMdwGjVHj9SPsinnxkOUp0eqpCwbFWG+idmFlAiQzl2fxiP/iaq
vf/ABeKmTQTKGE6tTG6MkqaqGs9pblhl7X/fRRnEiR9YyB8EtuizpWd2pYSqvum5
O5WkKaXE0ZORE+B+s6ftLeUS5pqbdfqz6M8YDxNIPM9H+2HSmfP9it1DjRE+mgjg
28QK0y3zODx4xVMiJF+Zymhf6XjCzsTpkv4yRcTuwJfLLM9E/m9GT4ui/V2A5NLN
81aQClwTAWev1ge3yXsHLbg0/V67DMR9opg5FubgJ4PDaun8y2HWDF/aSgW5JUIE
+b008KBpAWYSdZoq7Tk8LE5UHpNDwpYPAdpkvP9NAjPmwI+vdTrJgVarDeN34+eP
7O+5lLA0iYRSNiCohjBybcbnO7jxOGWUSTRN5Yvle1v7M0kXRoKxuGnKZwr6I4cf
RdtGATBJ7o/zADwa7SOlV3kwj4b0roTytUIt9F/aXXZx5ziH4V8c+cawgHad2p3m
cTTpzub4nXOBNi3eV2mUApm8zmISK1DI2MYWIuw0dXrOJSFEuIaQmn6okxmyeHEv
dJYrG0vFQ3ToROPagu1pU3c8CjkAMOWQ5DhNuvpB3Rrvjw76co6RR2UhLx43rsva
DhNbIESL/i0nnyjgo6RhP8e8lWSdolVzz5sOomSYysYaOU8re/NE2CLEbYoggw71
SvCEL5SzqieXyiBkmdwRv9bH4kuPPkj7sx2vdxHvciJNIH4EWVHs511lkGwH5cQO
2urcwU/i+AmVbQa2F1XzG/qmyUS5Mr7c6KGIO8u4zEiXitULeZa32XIkf3dlqa8/
2hV1oRAgKrThl2VL44ysccc7FTSHu64JiY41RTyhxm2VwmG9NMLmIPJUFZSQdceD
t9Lr+42ROpoLxU6iOFd2MBf7L7aXyJkzeVeWpsGD/aBXvgYyX7lePj/31ldLSihi
ASHCXB7blwL/8VnJfrnyTa0EaYITEFp/HrvgIJ2joRqv5eh4sr1jHP14/FPyIHP9
gTQlXG5hCU+Epg89lAFMjbqDq39q1lmKly19Hmoy7qp6zJk2B5wdKQpb5unIa/Sl
5LBx/JL+XSPHLoIbKuIckxRKOaxHMb5ITVjwhZ5hVV4cMokR769ME1ESWyLVwFbY
zps9z6cXasI69+vMBRfSHrIsSMj9z1SPxT0wzsG0PAPt+U3ao6sHTF8aH888pElo
IinRA87rpq5RG7MGa6egY39vc/3O3rvf2aDDmS3ZZFPZ+eLgMU91m8rUQCaZeEP2
ndHwbxTwptZ1r/UKNqK6aQ/iEUm/h7C1nuKnX/lra1UHbjGi47XocBw+ayMpM78u
lTZ4aCsfqAJngOuUmY2NfF4dxSHGsei84lwhUyQP/QsmQL6HPGe7yLysFCUCJwto
Fvv3mrjjl5lwA9meraL95o5eMxQ5zdmPhY1Mo1E9XOw8aEJdnDnZNU7B6qOgHqUx
+s5FDmNpy/2CQ7hTvTKNT19p90EEgGVyOGY8Fnj8ihHucmORwL2dpF0X6VjY7geF
12JEu2jVD3Unt4XVPtfYEizWvSd6i3sB3SXSUB4lLSf+F0Ozjs/+PRX4iCTLYvEF
3842n1LePc5nKP5/vD5woJakR2VOeT62WJfsReq4p9oam9ncwYoj4bQ/tPkhWZ88
b9DdfK0OqrtG4wi0m9jSfNQxGurqBZSuAs1SWpyZ/O0nk3QUIgk145z2nAfSJ445
fQFGlJB+mYT1ZT/D7zDnRV8MPOt1k8DOmlyfhqQY9ItYMofMwDxcMOYbIeQ/yy/M
6vJeVQ43gSBORq6MH3jqLY+5EnOoldDbdDNszJZsB5MuSpfEiGlrs/xi9yLF1uab
7J7zFzB7NHZfqCucV1RyR0AqY+Uysa5B6hbkSg8lTB/iMEjXJvsY/vM4qE9wTtql
02IarxOquiV8mr35M1iehgMDKC23UaqY7d1T9Gm5U2z5Hi9QgzPHRJqJshNFVzdG
P4XDXmQJdtnufiNYvmAlV036JulTalYM0+pktUSir0MlRFlipExy2Q0tEtTxkQNS
tdhrJWmZDWspI6nFdq2D6XMju7frPRM5op3yIzMOj2RuTUt+pOqMnxkRSSGqn7WO
IjEGD5yOkq1/h6EENZtlZMnVq8ECsFm/HVez20lQTAdTFYkF+iGqocn56+UublxS
MSY/Ts+ZrFibDqF4TI8EjQAN9u6PEEe86sIyFx/f/P8vLSt6LJEDpuryNMPLZRLK
g9SJgW/aJXJwZdHNvKkZLxMrWFDy+JQ6VyW/gpnliNalNaUp0Eda7wrim67fm+hl
FoSkj5gnnUWazYKvB8MyCtQNE8B6GJg5slewHhksnIS42Jr3v4on5SmchlIsBpFS
X8Pd6RDpPJo2Tf9NdT/MCxv/78VlbGyhUm4RLt2SHlnHtUt5rY3QiswB4Ojg8kMv
gXK3edu5ZJI15ZO+bAi9GOzLdbr99J0SUda1U+pj8yg/YRHO9dfucKUMjIwjDRUk
uKlilarhtKg/J9aVUbZuWtao0CC9A0ROqAQVpGCS9l89Rr3UpiAzgxnQrk8Tvt3F
B/TV5gcSk+h2iPR3+R1xCuSH3PhuPyX8vza4Nq8occnkKLSey0cFTJ82VUjh8b01
tXS72Bd5/KD1vut6qtS+KwvnxbsGxMaLkSULldfjxvENbixkd8vDV47bz5fH7E4Y
Nekytv5ujpnERhuZBe5GCMWGzEPHaSVe/OWGeGfbB+hR99IYgVQGTza8TeKvI7gG
wL0ORDtAIF2b4sf0jOq363eCcP+5VjNHDZPMcoL3uXGoxlASvA4zB4N26kEpsrOj
Wpg9/hWNO1UFY7a09KhtI5IoRvKWFlsdFv8zW5DjbdzxB6snlxER5Cd34Mb8vr3c
9LSHRxGVz+C1/z8WPytLrJphiybt15rCxAJ0u4fDokbelr8qoLTMOUqoDXad8h9W
VsTYxzXRolkuK0u+aR6VAiyEtv6C9s4voVwwWpGBDrAsS+0SX3oyQ3p0rX4hN7il
8yfQSNacb8iMrWDMGBv3HXFA8oMjwHx8dLKQGNzyNL/9Fd7O7X+4uj1ZZfDl9AqY
O1DKXjqA63toMKAnEZx6DQFaxLld7Gwagoy0A6K0Ng+eq2bpGrSd5yFSSTn/BLEQ
5LFqdSNUWmNq9Bdj0sPckNsulVA2mBasvsXBeEB4VR5uWLwWoZAZ6K3LtZxKNoyN
fSg9j6gzr9hFTPtsMPDkK2Oc/ytqcqVa3wLIZGTjB8o=
`pragma protect end_protected
