// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lS6NrYXeoR60C1bBaHtWhtQBYMHnE2gR9fI662k6jfbPJzO++UQW9yz0OfVRGqxL
CK7+XTPD15ZMdU40zBrsFsy3DiuB8GUT4Sa0uGqUJlcQ0NCuTBOcnV1K7LMI3uaT
L3lyexbmpDP0yO2kj0GhI2j28f4WEHTx8uKbCU975f4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19472)
M1m0WV88860qsW7SyNfBPRGliYq+3AYXiW/fNP88OWQOllwmcnh9FDJWqf1SJvUl
CQf4yZkteSnzu3102/xq4ShONf42kGRqL8gXa9wv6kRC/+ulX8qN4F1gzzbY4f7H
eQBMCr3ZwRgM3o46K5nGBRv/RDmOFqPOqFvzyAjeoKS2eiEr/Lz0oNwNSXkmys22
nmy5SIwZ2v5NDCWRZGXstj8sg817b5lsZbNT+D0nuvLede9bi0AqP2ZZNi2AdXH6
FpbZlvFwUDHphUuOVV0Y6ysUd0o+Acb+wn124f8rbY0Hdz/637EFbGxsrQxDoCPA
uPa5mII8TdRKg00QpdlIzMuljdu4ARw00bz8ItXN1JF9JzAs+jhYxtrPN/QEctJc
ltWJHdCRk3xUXLL3owZQpLZR/muwn67gVHHwZMw3DR4xQC/qAHUlt9jaGZRxuXve
VdyxVINp75GJsXt0hQIzDJrVdxDAiZyKurnEXbg5ALkc0ZgiKWkeyuQ7SM+F18fc
lxVJ41uZPD4X1+ZEss/7h2kNYcZ/qahgv+MsTunJPwdF7lgvB45qvw3AlrXSU1wc
zDpqCmjVatmYvD8pl64W6Wmq4vjC9fGIrX+lN8684HKHSUb0rbj0Rb1H//jOFOvz
1couV0p5822wBbEQ7EAoPr92HZBmdRk8bhUZtm9QMFmxF30vZBUpFVsr8GcoQTPv
jPC4uBTArW/dGjSLPs763djYtwqVL7ebW7Tn5HpMr3VX08U81YVD+f+gO3iKopaR
TuDirXsYcg1xXYesWHKDdFaubDizcgfW7g2UwYydABWaZpWCRYp8YWKdzaS9IG7I
SwY9mbG0U2caJbetgZj2+4RInbSwGYpyYEqyy9z84UZbZnGkB3kbeA7pFTiMCfIE
Sf3cA3qyAByyRZG8ucOguug3UnSvNJBv0sSMmHlMH5C0QJfNtb7gO4GsMOCee3kE
GUHKCXJHsTovtBsDXTwbyrhB6FKmvsaK63S7EhlJq2cbrSMgn8LwzBwhVTL1UtPT
iCw0BSlFqwEQdA5UJU2lkIPZAerntgychkcOdDTfYiCrRLtcpe6B7MtzVYAmYhvw
U8WPcpb5XbV9VyMuYr2BCZ+Ow6kHEJ74NZgvYAZ/NNXu+MoREFtXRGeqb4D0n8oi
SAuzpGnFHxw1SKqz8E671nFscCRvFGQtrQt0T4U/m9+kC+HJ/dRc9f6pNoxaKNuk
ABjPoFXFieJmn+OVanPZIPHiEANyKcLZO2RSGjRo5gecrbVxeuxqQogkexI6HCYz
BgcySEZusC6XsTY/uk5jA7+V284SUU2V8gQmGPFfUku2n16bBw6hRLPf6ZdzHtZU
Iq5U+wz40LNFzA33iCTGvZrHO4GCROLF6Ha9nlx4S57Y7uqCUIHnmYGc1ZTjJO8n
wnXnEvipfpHKPSDNYceb4gNk1mKPvfxCVCGOI880WvmjOLEVoWialV7T84/VGbIA
dGghmeD3W4YitAkRqz64YbQFXFV3lTcuOI6xk6CDNfI478meMT7OG4gpskG5Jbgg
5akZdu8ThD6zR6D7FejLVGaFMtjGrWp3iWzvGrA2LFpE6e6qvOcS5sdCMs3G+8yj
BiaYRmRQlnIBZUhChWOTbZPL3WIkg3bWVURMPtITNAfMPcJbgHZpIfZAijKRtN8Z
B0SUuo7MmAnXwh7nthJXE7j6gg4rupnBfZHsZc0bg3OZTycjnHFtntUFXSJU+ag+
OKqZRXqVezOeevMEKJSM1xmiIV7RjldYEgSEJgAdkDCOXmOwDtIijMmT67JuFjF0
zvalUJTblYGf+L6fz0QcvsoGgiKG9YF3S+IUmpHzUuZePNy3B9+g2VvwhD4GvoBB
gBKkBfH+eJhpVGku72f8yu0OpYcslLk4vlLSSQX0w2PvlC5lFf5UGIiJW7Lfe6sc
6Tp4gARATECiHI2CUuWW5V37ha6SxURDli8DK+l+ucEHOJxDorn2IkR/wVRL0PSR
jSDf6YdSgX7DmvYo73uAqBdSdptEitjQghnesQKxZNb0b46YGIvlVv9ryliGduS0
O+v3JunUmnanb2PxbZPkLP9vwMrMO78WdkrgNjcgK04VBci4bgSJUXq/llJi+Wa2
7ldx5tJ43It+5DfMrwAn25HxPRy+Vzo8grGGMpsPephkloHU8uFG4txISSmk8rC+
lJrYvYJgsA/tRTwueYHkCp03GrSTdf+ZXPUwuPafoCKRIXxaPLhHmlWX5CFLrYNG
lNdsifXmXwP/Y4vSBkOekk//4/zfA20NhnwEJ0r5L5EvApVDliaM5Imc1YPYEzp4
9Q7wkE0FBd1JE372rE/IqzGEMXqvjApXO+brD4Fr5xgn0B1Jlg4US93TnMlO8c21
9FrNoxd/ZtxLuEzjJZhjjVodKvE/GkRlXaBBAKdTn1VnKGtMmOP8P+/Vu/KZu+eX
jgLmrHzOZJVpmioHscnsXSEjickvvtAWDfHa0LqmQzjpYxoE0LtqjtUfgubb9s9j
P5ff2/L4EYvnPYtB0Ud8s6PE4xh5Tp7IrZmOK+W2ddjocFZMu92XZ+pE9x1WI1d3
qBb3o5zsbrvUZKFEW8XmwkXZdfsHpJij97elnrC2wr7sb9iH7Pvd80xssZOMD6U2
bkuvS04qdWG9zNx/HgVF2KJ9XNKEYVZDjuL+9kZp0lSlRnZOjOryXmevJFOfmnr+
egb+cQ3WIrLbXkkVBLmB8ZgKCpRfsnwahswnYewxdwaIcx0T2n6GgPqeS8AMSQxO
gTJY/UMkGMO5FKj344/ymgN5VhwjgFEAe8p3dsHr2xqfP+/gi8+TqtStt4vrMUC+
5VXAJMF2sL92ciczA+rnUqKe8mhXV8fI1NdKeagrU08wWu5+lIiNSnqBZ18WcpxJ
8Ce/+RkCOfAl94Yxe23KTNq4n0UTOj0c64bYh5BqbKrhMluh5rzBYfTMJ8OfIE0Z
Ugs+05a3YhwLRUwzcjHQWxS5bGyvzskOYiBgo1+tIp0E2c9hpzMltgRABlG7MCpI
c9TY1h5pkHK9PETV5d47dCND9tdixIOsWKmMu+cG7CtjZGdK206EndW6ntXpleNp
lVoazUtpQn+ZT+5gd/Ik5TX/lL2KQH8GE6H64z7XlTA7gbnSYXevEPth1YVh15o8
P6yV2utnlcknaLRlAUfuKpJbVnDjD0fYjXgvERAepW5U0nNcK+mcm0IOv+5l9Mxd
W8GGCgwr6AcA/HU+5ig7YPyNcxI6jmPiJr9s2V0wamBUeVgGCVK3kffWPP/J5DRI
9fNCBFp3NFJlhGtvpB+e3ZEAkHZKEjQNcSrlD5GLmzpq9o4ee6ahd8ym+2y/oEwX
fLEb5kaWCvopU0SRV6zMNuqcNlnIyqFue3foZdMI9MihUCu/QIvgwgsyTJRJ2vv/
FbpWTd4tGFa/3mcc4gkKjMNQHCnHMQ21TKsSXb6Z53SLlY25ADXWDzP0Rc/RZbsL
7xIimNTTnysw6U6KocJ8FoG0t3kwvuoK4XI7v5DLKQDbb+72ia9yUQDm8LcPmiYD
yAE9LErRvsfJ9sMpxLN9X3LJ34TcpVe+ZhsjSNxU7PWGF1E52lYMvtnNdiALnejT
f0f5xAMpXK14IIS3djxGSuXU6cYGZ0qvBjSCqAv8ms1x17+CxFDlFVOm7pgnVpRX
5xlXVfA8TMvi8QQ5Eb1aXlMCnts+6gDbiIYciWFX1gAEhTLJ8aeEdE41VYUwo5JO
n9zIng5UthKJzTIDslu6V7n4asBMiB+FnJ4vxZjn9DmipHn7bRekkW4ac1TFIxbT
LRgRy+8mYnFkgKJ7wz2G2kJ2zI9hxxkgKbkY/zOK/IjH99OIhpJTwmZbFkKrysVQ
vHeY7opS8XzmedX9evp77UFUZqBQJke5qTvQOfHw6huWx4xmvGKLfZoGfsYF/TfT
vXGIsqNDMA3Uo2eQfmCwM/DWqAv9dU/Ha+lVKr57+v76WeQt1BBcakGwlyRRjmo2
alt6fwQyrqIB7cvGNEwGqpmOVNCHHNBo8b6ScTxpxPBc4Y0ulSSjWD88SpNOENqf
eThDaKiRDDmt5Lvdvl+Ie6lEXJh8Qgdsafaega9I6I/C9elORdHXhy6d7koRthoa
KN3cNHhKhNii/RB+mXyi+4T+TE8pnZ9WJ3iRK5cE9de85KeHSt/lzozv50tVAV2N
Yb300Qf8+0cJBTBp0lX1ftzIl/P6IPD8S+QdbhvG27+/NUu7f/yWIQwcElgPmZ10
92aFwibWkYkdzW8khy/4QJEwfH2Qhm9jrRobwcHbAniof+qWNnTTqZrNXEiai5hn
uoTbaELlzPCpidgo79BsJAgfDm/JBkuUDy32aXkfDxbhK08SiB0sBqMcndhVxZNV
so1naXQM4uoOc+rI/Tj9SLLo4MqmKfbZs0Yh85TVj25eYuwTbnKiaDTbHI3tt500
+aIcpdCb3LWk/CvIrd3z98egxMtQuaMfHf97wNB6ypCk8tHOtvnsZqNKdPRSECs8
FfQ+J6b/0Rv6887bG47gpv0754zRr/NBn7SCZQ+ekR7Gd+dU+/VCsABQIgVrkfOF
dOum1tQBlhG0t8hxf09wFx9bgJoIZjo8mNPq+HGFDpJjQC1onF8fKKzXuhadn0Bc
90E8Q/58jQfRK2d+/fIN+un1DyE99FGf8arZYkisUUUa2NNri31RNeKobbIxFxcH
h6gqBBFRcN8RJMX6ZDu6pkiIzT6E+7Qpk8PWc6IatuVk5Ux/yguA82PsEk/oWrzr
nTzGYdRmEDeaVR2J3SVvs4zwxjM4LkcLCpib62PZTu2KKmQXDaTj3t4uBjpbuKIQ
6yAOxrcBBfMqTYFMXLVdQwwVpJMhp/3zTGEX26Jzw8HBpxy9tdTNiWEjgOnZ6XNJ
N5aGsKX9kfu36srTjHR12Qo8kcIXLxadqHQWCeXx0Vmp+Jl4oYoYQHv5BraNlURm
dWvN1sQnWtw/KRRcMHxv/ne12D2MbSJxHDB8Kar1Q9mJ1ho4JSRSr1csj6LStKyy
T0bx09/LwbnFZH/gU91ApbtVca8hGTkxIMVlG75b2o7bXTMX9d/XjLX9TRzea2Cl
TXlLZZh7ZcmfoDFJkYhUZhE/K6dwGdfPf0IpPVsLh1D8yW6FHt93MpYdo9IchUOi
Iyc0+JiiqV8HS6RnpUoSqX7BcnhNe2cisP8YI1GuUeIRcmWtfq+njsWRq0MK3g6E
6dIv6Aeb8sQBYeGY1Jj9Wia1mh461qvzO6abODvii7AOYptnyMFoFlD/0z8XE9Py
b4HwP0USv2KX/kzf4YotwJyI8JL/cOaEy/8PWQW6breKN9nGIPtfWlb3YCczEa/d
ngLvzuf2aWae7RwPTQPm0V5yAOsgJcjUCLvcU0VvdknfwCkfzgJNeB9SF+yVOOhK
zuUWSCm7iWo2fUtoI799HnekltYcbmS6T+7OYvTFBhtItjDKxjYGeOFw5BLlamSg
12HPYCYWFOz1Gs/moackjWjAi3qOtLMgAJyHI4OYrNEPjolkyc1jzkIZtabh66Vc
gR75LfFMfCIt7AubE8+VQ6D8lF6RxzJFh1tIFwxWjjdVVUxu55DmgGhbrWZ8bTSD
Jzy4F599e8U+GFIreKMWwpCpeqCQn6nY32sgMyTEUDzYRtXg2g4HLATx+1ehJbBx
7SPrF7o7l5mu51+VII0HF4TCD+0uE/eqwDMAm15URCZ4mXhnPbW8kAsDGxzU09v6
IIudemH2j3plofhkLZ6lkhvLfAAVfif7nZV+gsTP49Nr36FkfCp5OHXak3iBVHiO
A3aYBpF4rQtBXdkvvOsk+rmR8IHU2+B4NF0XjPLXYj4QLKOxNDvh07v8o4VhjYq+
LR1DR5a4UaNIsxoyFqv0AD9q4hlRtaS4jlA/wxqwFwscNo4xIcE1i26wpyydU0FJ
aDLUc6ODGnj/z8bPlYmw0efuI/t0w3830ju+qWCSYvGwLOAsS31tqmw2XDBhjE/p
6APqyi5s7/3CL0upIYCaDe3cyCphPddUnX8Xaoy6Qe66ktIGRK9WlMKowYAyH1kH
fn6ZseB8BeQW9D83toXCa2dLwXBhT0ztkvM4hCsEkvNKPR70aBqyB/5QtnQLPOuS
JZ2Tsp4t6ahzy5GJQhVzSxzOO/3RFQAb6YuVo02RL/JjAquZnN7N7Fm2WcGKQLNQ
p7OPLN4n3ivfl/45MaVtzP3z/7694Xi+ahb5C+pl1GVsgtewP8OvTNXm+jnhVTew
nHiw802xaKegCx1copLdrKbtIF043xKC1aazgDhM+uwR107SeOVwSCE4QPG3kflh
IWD6O7jcFdKz0yOTjvFJuE8fYqz15NUve4QIpnhaS3gqoRQDCcEFi+na0RtQOj+R
t1DFIPq9Wm30R0Oqpzqu7JwLVqA4PQrHpmPHWl+YYNFtS9L7d/zC17YfxcPfT0sr
MnQ0HrmuECKjqqgk2RgXUQt0ONxbbButW0ZdKAzNJiKrvvKNqTDRfKx3c33Koldz
oDLSj4+izCSoInYFRybA1ad31pn8uOJjOMPY02icnVAeaPWPuW3WJkPad7YxdZ6u
F+nJ7ZbNyViqlr9fsC4eJXTmGyPiNr5wsCpWnvCYkEAudSMTkwIhV/nZVTRTQLDN
fQMq4gQqC5940nIHhDcyltDQN/E9BYDm1KlZjdqH4m5ZtGcBEfRvrPTzcmI+Lld8
yQlZ5w1FRLIguQu/ki/cJdDMWfIpQe2JA0Z5Y572Bcnmh84lGVDBGvMVBA++kfcI
Ue7W59fI+KkoVOS/wg5GiicqHiLWBtoFdu6y5FkDVU8dMpXWT3TGvo1TiHUibFWx
Id+dNpTw9brySrYv+11qaZm9IUJ5q22G/SCSOhcg9r93F2hkmwvmANVMP6uOXpbP
ntsOYEqGJNmxP/YtrYVWajQYIpiWHjyOnzPhi2IE/rDF6AB6UnpNWs09fYvQzKV8
wC7NY5oDoF51q9BqVG/YXZIkZ33mb3dPu6C+ySnVLAIrOYrhbuJu0X35Hg1Scnmr
5aaFzwVTv4dbGaBKksmTSiGkK7zMLObIRiVJ9924FJ/TdB10/uW+e5UE2e3bXYXz
5cs9hlwkSuYsJIaiMoaLBN/3393+Atg4Nsm0f3cZuwQGFnfKZ1FZG9ZNMgfELii/
Wg0dXYkYDHGeF7vN2kW8i627EPOm7krGcuNu2ONqCseXPK/aR7rs7Mqeu5Mc5QFZ
XNVVCV6Ncfd3WTwgtCyOiGZmpg1JuaFKX8AHbsXA//ZuLzOUH7CRpWi/spSZ/Uor
wBiNgkLpRegkX33kHU7i8inEXrf3E/AXV2wARRKkwAMKNgn5cAAqpcfM5O/92B9s
2tagNvPikwFStFezCJX7kU7LjcGiARleKyE/huVsYlbkWHoCkLGEfGx7s82JZDzt
kVlu9z453PmuJjxmpFFe2QCErrfnpeSwxC5MacnWyJ4xh6VvtxuK7YpjKELNpwXi
S2zJEqpbUY4PncPdbsnP8dZNEAHpPpbXtvuYZSo17Ki8BZGxQN2VrgAcfX0upodV
kR3D8vPiA7lyh/H6LbfjedO4W9BzZMX5XYRM9TK0kmd0399BX0/bKnrc2SXo9/tW
bJjGIcTa7PFhLbZ184pP2t59+Bou4aZeILtpUy3LQL0OV2EACYBUbQT4Z3MvgHgc
oxyprZgYwbWrLP4yw76rN8+FCj1Ti1YVFYtCLHyfVrlUYDfg9we5Oh0WKo3eIfhh
0RNFx8txwWRO/UD4hS9P3M+0ynCk9rODgMbtwILiWzRw+QD0m6phK4rQpAQjtHQV
Y04vcXI+G/J6yVsjQMYXnW5PWVZtFxDv8doWDLhqOKS/XrlgJS5qNo4GtWeX8M6k
qW8O+1WgvpP2F+foOEm3MtGuoFn2GTQGR3J8S2cWqKs9iqYhl4JlvQ6oe72RqoH1
s8v4BJ7UKrX7emihM5WJq9eIIqw0N9Ne28CK0ZUzcSHov8thcg+bJJYxFpH2nEw9
LXaOq+pHxyafr5p+CIFzSi47eNhaCQCO8ld+jTLQsTTmwYy4u2sC52W77kgq6RJB
4HBxgIAuAcgMhYWspdJCYHDYS5IC2c6tItqLf0WmN9nHjZyPtJJ48VmNQ+LozdlF
y0j1vSJAVKjXxaexQ/1j3mLyYSsRCNPCBfSHNiTJgSh5zC7EuTgi/SxBt+6tD9Mj
u565X6wOffh/Pdd5ZvsaLy0bdKkEsdZjn556yR3BYh8CYGpMgmz03Qhw+enk4lLI
OcCfQ0v/irzqOivKMni2UIzItWODrLyXG7un6FbsS+jxwVUXr+txGB6aNV3/B2BH
XDL45HZWAOhpzIcjdtaXygr6fMtMHcO6vgmUXAYOJDspJgvEjVsPggngYnsuboAk
TvEbN3XESU2hyjRVYlThd/g2Z8vYN4CqTGIM79Crx8i+KZE1S/jhKRy+nIiv01Ke
panYtlpwS4hdib9XwEB2S2p1gMYCx84HP96r4/XsUm/S14OZMTBZvBfgMF+aTiCj
sIkIGfoR23JrH9kaUFntp8Jy6Ndz82T8fvf6FWz4AQ2wnHhdP6MPKpDJzprDDMpP
5rTqUhNq6pg8ncdhOgx+X28OItVpdhVyXdiLg3BliLEybEWVkBvkmlpoEEgN4mag
h3EKLbNeoBVkTw9txmf/0344U+keyFpjsNzQh2e6TcftagxAWOyUSoDQt2YntvTQ
t9F7Oh9w4PFZSOjKCnPburI6BwFG0bYSgVGM6SUESlatX+yQThspnMFWNbpUJ9Pi
TwXbLwYo+DDq31HJDQmDAYRfHihdDor42cxnj9wBMToqQUpz+kJKaYg27d63gGQA
fNA92MQISv9FmQoaaZ/VrQ4YgU1T+USsPzYc0ApPGg/Qc/BLh3R+HRzp0+WjfvyD
0Uu7np4Y6f9C/vJ27zDFIKRoGMAX+Knq5290I95L+i41h5aRaB9yharXsm3ylEmF
vuQf5e+sLXi8KahGQr73LEwma+wW3i6QfW04z/hg1/RIQIbiW7OGRNkjv3qtSEAb
p3KTcck7qwasR8xpu/4p81KaIcm0gNTChFhK0l5QtDrlzHN86Kq0WtTeOK4LsWWe
IlyjZResicv+vn0Y0XSB8YjNgZBSfsuis13wqLzBz5Aj4UOf0qJQIDOYbX85w4WB
ffRYEH4xdHRZpPeYhe7fWQg9lPdeJKxmN8e/2sPbMe8kpLpQ6qWYF0IePd22ydrS
IkgOsVmve3pH6KC59T7xCElUdQNxVgTJnlzNb970QQ/hCC8bFkJdEqp1gxJm45Bz
1jXM1R5fAqRCdZjqLrLe9W6iqbVIdtBFDJey+DYP6SwpZgxbmwnS6LpAeHtU9Shj
Hc0bT+I8A9xQ5Hh0dplc25M+iwN5g010bR3WHvqe2uzVQ848WF1hrAu2eMtsuKlz
NCvK5KSZQCK0Qyi7I78uBkWskhQtT/keSHBSJ1P2CaBpm6U8losCTluknCXa6ZRG
8zru29v3pYVQC6+czUe0YRTumOJHBHld6aDpQzD5CwZI184U94PKEGpHM9sK3m/X
JAK5N/EjstN+ItEQZCh33y5UHvbQZnkr8dn8SEqRZWyzlQ2/HaMdNhg8Z9QtTC9p
fQUBYH/Bfk8+KhBaxTsTksbm00taY2forpSZ5Hno7w6vXryHmfqjRQKwu3zzU8F6
483NhTfatbNjeZKHkNRqt1BKisUQ4Vjyjw3HdvA6edBzn97Eb4sIU7sYb6kXLbcC
k91zCcyZPNlJmLG0qDqFJ+7O48G4APZn6zlidzD8BFNioT4s62BDh8LTj57WjEAV
K5whWJqpXWchQHogHNjZYzAqjdWA2MPb8wfuijPc9KodPidE+7g/eQU3mP0NET79
me28gr1UoT0DkAL3XpkPfofqfECCXILsFKwX2NG4uOc1bUUWOg4FQ0uqyglWkagV
vMo3uJhgqPZ2IXwC7P0tBBQ+miIBqP4OOloXRNUuW3T6sq1T9tgIvTZR0xBQbKic
jrrZOzKOJq9/PivWW4i+DoNJ2W/I27CZMFQ4bpp7u/KY2ikHrqf8jkDwB0HKyarv
tOp/6wwlO/UK9VEVYvT/lix7/hhHy3zL2c+y+tc8bHr8ikYYgf5BO9UsKcRuXnhb
Qc8epHXxD6Lzd4DcxgT0CAzyGmpiPmPuYniYIg+mUmJ63rQSj/VMeVtpS3RolHQz
TwSyRD/zbXoF3vFonve2b5RT9KAi0B55CYgWXWQipZvx0B3lhZxqnMrtvgDoI4Cj
HlrCWTo1M0We74bcT5e8ilSstlIM40k9EukRNpQzbhcExkyxcGAPmkQwy9YjSJ5b
2hvK1jl+l4a2lDddCpnNn/NdmzgIJq4DSSoFyaJSboOHSgSypdY3r/o13OyuC5QH
bffJo/CNcl9feregKZwB2Ie9OubhBFnTf6gr7kn/KKP/bx2SxZ6h6sDxXSsAqRcm
qFuIWhdr3YwbfjzgWFLQZUUzt3yzPwc1M8fHWc93F5SDv/IdGIRFhcBp4fJyn2k8
dWGeVs9ApCnImj/FyEsWYMkcnqwTcHY/6i2rdi9+2Zp0HWMM0yj0eLMFMTxiT64y
ZHA9rf2R6vpecv+gRb60ioGnsgkNDAzzGjZ7zgPSz2UdanxoF1DpdOFj5W/Mgupr
6Uq7Tv78pVON6QSnt1xmTf8rrqNPE/YZs3N56BETcug5okMTsVz9/m2IaUmATyWJ
acLnaEXWJmFFBAAAtZuSuD6OcNILnlx/UWvG4NzcEmGu1QDQSegSHrzBb3DSXXlN
6BM2hifLO7Gi+D2+NBUqV2xRTZSzHNVNRQJqkTUGJDoY7Mo4+7yPBWLwjmiufH8G
8sBB1kGd98RAJtPh/UZQ/Ef+q8nneeX7bR6e4cvEBoLeucTdu+wTBLJ6kZIsASzk
CaPFTGe7YCE3WxKRDaf1gFTxTU5riRobp+WAfXSJRGFDl1FSrwIJMmqvNqEy8gc5
RPGkNeiCYSTy4UuTVGRJZtu3u7rLYF9h5WZeoSXKtKD3tuQ40/lCFimAkFsxr/Oh
c9MG2Uao8OAGSRnsy2CfY6me8ZG7QTqXNs+oJ4bNWxuWDliGxUtSkw8H4kHDTi9l
985ocThOKv+kqCShyOJZjHtzOYliTdZKYuUQN1dO+m9H/KCkI/dnErK3r/+cB3fO
VkEBeG72X+nQ5CzsZyTqdt4omDsvNoxaHK4d8Ydb4MmHEC54B/YgczzbHox4GMok
HbPASnUzkwsf+FVVBHhqtV35ll0KIRHdLguu6BfMtShKwVHR+MN+TztMXyZlCIsN
+r1HQSuSvdxa8nmNHWJmN6ihSZVJ6vyJbqwjghTRUsJuoFTey0cs9FQKuj8Hxqj+
1plrUJK+dCc2PAC9R4eJqQtM2Kz+iOzwFjeStcFJCsVg6HMUTMkUytEgAFMZI7e2
oX5V8mxZT8DeP3aZoXERhMSH6BMuprh26gAArYaa+WblIBh6tfDXYI0I9wMHe3yx
AxoI+tZX3OvRNT0UAZFcRCehY0q67PkG1Ho073pJ5LbyHBBf0i+tZi4Ed7i0VQOb
DGeu6MkeUeNO6jBEddsDjAhu7fRlNT/G/T1P2I+VJaZGDutedUrumFeYJDLRu1DW
6HzEPZ+ktuwRy7idhuFKqg/Gm5t9RVfjTj8Q3VqfWPIEexGlaIntBZyCMFNNZyqQ
Ng/pDy7TeHdqRSBFfkpNshz8cjxa4JQSFwT+9TfME5JW7OmasbhUSVHw7/swocio
JBFJY6aNMi++di2SiwAQgz74FPNxrbTW6r5M3y4AXjX7s3OMdtjncWQDJSZFfNoX
fzBPxLVR+bkOVEglXhcHTiuHCKSuQTAFwYd3YLTDJW1o6JAqFuJ5Zddxp19o+bo3
mN9YEeZrVC8deEnug5bxDmw935veXwKj7fj0tIN9COb+wVmK77CIumGUefm7zmCA
Jal81wFGDWigHb6/DYmEFw406eRW9LYwRI4FU9J3EU+o3sv7X3+B/faaEm/uPqRv
CS3w5PgWTWh04y8VShEEJ+g343KQGRISyG08udTsWpU8pZylQCoRklv1l4+lxsaq
1rqT3P7ZLN4He0hO8nrO4zMc5MUUVPLciZl2y9lFHncMBRKKRekyWiF4L51wLKJz
19QJXIAAWkutqhUXrBlM41oSVJNtwqz+oGCxJT9MhRlRL7UmbYy6MBrDzXjJV+um
nJXDOaVmDPTOTA7fq+0b40JUD7uGqO3AusHDr0jmzRXkgG/KOe2DHQiMQ1IpByf2
hRaRmD0uUcHLSWPqYZzdo+Z+5O3m2oYRzjgZhgI1z/GYXzElRfRFsqqME80O4LUY
5YwJktmA6TqF521f902sRMxrhgflGelOwOJhwdugs2mRFq0z4REikyTIuBEwQOO4
W/QPXNaw6De/nQ04FgjZa8irWnCi6ut3MZlMLORXH9+a8Bn6dvpb1ZHC3A4DB0mB
wM0N94aHZbwMDdmPuOrInfD16Py8ZwvhkaclC8WdT4qD/gf5TSDj+sozRCqWAziR
FI7NiM2RAfRSyg68fFVc7h95EjZm3QUC7oDVdgUE0AfKhLDvFWiyMiV/cVVDUA7c
3eDBIhZbq7g9nbyxvYxlZo62o+FAIFWEcDlqWelnpzy36ZdQzBZxSGI4UfT3lp6H
9cUXS0fT8nwVeDtCH0y0CdXY8KNf6IvZ0kOXvKHuA1NCHnBJWUvCNkgP2KCqdZF1
uIS63zVdanFMuqh8PA8zYKNwcr8SrNY3ATla6XhrWxrrRyDLu8eIG+9Lmr9rSVdZ
X5vhUkvLTh0dXqoxItiOeuDwJa9bByUNqYTB1ZLg9B3mFLOyyiREOMg+zF3TIyR+
XoEaJ5cPbrbfcJtMiinqMyxCBoYLGeo11gGKbXge/X7LbZ102qI3TrwFMvgqZA7f
kxm23wh4rpZfsYP0eDT7R67KAhk8sOBt+mAkfSo1QHvvwCDT0ymU5sEY7VwclaOA
j5i60RwymYj9s1LGrkobWkfwbK3XnQanF70jMMSHJpb4uOAkqzjPcRPyWc5J8MPC
SfrL8jw1sP5WcR2KRl9kuWwCyMysa5tSsy5gBXfLcNB3JmwdT4pDO66m5tszF3iw
B1r4dXNYhNmJ8+68pE9g4wubTuFlVSoYqM8OPDvE6TsN2xGW8UCKTelUnpSCIPCu
4PUeTS+ghm9J+U8i5j74bK2YUFbFbYMLm6jxPXldV2IHceh5vpy4tqUG79quB0IB
MacDjf38sZ/1+2J2sZTKhbbnAYRzRxnQJDzMubTvpJryFAjtnH5c+sFP6tFR8hLW
UwCbpkxNG4vsjGt+BcC37ymhcvd+jMSmzeY2RvJ8r6BaN1uHyNWHYwZHROnWY+ol
Zop6SbtZdRKPg4xXudbQ4Yiwk+ahCTzzwKPxridILGCPiPBtYmTYppbLL5Jh3hpy
g1HLTTHyLu7jc6FebYMFCNR8/ayj3ffkLNw/nWaHAeb2RqvUXnnGggjrl2mjKaKr
1Wqf4Ot6Dtz5t0JiCr1UaRvIlvIFYWAfnY73qxZfFJXWKusMZIgSnhIWFawoIHam
B8a17kBzq7VX8M0Jz/OVcEE8ORu6LYIge/8K6kEK57zrJfC/3sQVBgGFpOKougTe
y5nv0G7ZGmwflCoifNPtI/CMdwgFTuEd8yC7oeNDakwNM3ZmKJmRhtNwE3+w06Ni
uA4Vuk0u+K6eq9gjVJO9x3gXE1ewKvsIARrbsE6q02fTUClUdYQbj8FP1TZaLRDS
N0ZdhITVenruHhYCG9ApDeBsx3NA7tix5WZUCVv2uBrxOUeElU+SMh23w7MH8GzL
p5z1MWh1K02N91vckRKCkxinhgpzH8NbozJeV5GoTKRCN8cH6BBiwyfxxjCZYtJ5
b0OKc300c0/AZfqSEw5J0z2Cx+daqpaprtda/CsPGLvCbp8dbaHPeZvPcX7Tb8Ks
/fQkLyPiVyQtXJivOazLsBGReWaL1Bl31TnBIYVdqSxD7HwdiVgYGPDEcbgyd6Ho
08Jl9CM80thg0YYkjknwezN4Sw2jyEAzKqiQABC2CwYyaracHy9QY5T1qrC5Ffnc
mgcnTAmGPcSSmc4jN3wUTI4r6GJdEz1dvkal2YWjtiwl3n424caeQa+rdt23CrtV
6m6+ZZgnO/91xT/DQMUnildU+1zfhu0XNBRocV7tgq/CSEnuWcp/BFj4ZOakjN4a
O13d9incFAb/vp7ff6bZ0vZWulDN/+8ezpGrAsdAo1ASjxL9u5GTbdWsyfwEKK1A
Zps1iMaRZmEHadD4/KFGvC4qsi16WBmw+v0EbD42/UW6Qj+xkKGE4IAUXevaDGyx
0D6QCwk6oFX5hbUUKbsjYaxdulFfye+N4594uiz6tWrcYW5Uqpkjy+vpRdoPqlWu
zD51sG70ItDOvr1bsP9tGoX2iekljTGuZrTg3yRdYRzZinsvXdNwWg1DQ4zJOebF
CMEG3Vl4IfysIaqLtylaHOv8CDSoZ4yDwrblsDGMZ/v/GeqoSA4N1AQ8aUwGvSRy
9cODcCj+EqEES5DRvT21UUkmfIDstcxcGbWlabGwDP6i2FgKvVC1rR9q50JiSure
LnPcLxsUniAiUluI80K0QbOvOBSS6mAMaxXaZbrS+6/dabkoZAncEbclzrG4kMu8
ubndM6m8nEENrRsBkBDBYTKPuflrAdf1BS1xatRtH/SPr4PWXwvg/eGKkyLwi+l7
Jl6+OFIM0xxi06wLwj2UE5nh/112/xyQ4D7ydv1Hf8i42THTrh9GiTMLkOgmA7WZ
jdPc5/z+nyHaK9AhtT4lFapJ2F/8/xMWKh44pqucIDk0gGKkgm2xy9ssyfDkHR3n
xdscZuIlFMxekXoNx/VbfR6UFcDapZeXNv/0DxwscaHkMNmdbpTsOPbLadocEFs6
rAB0mQTljiCsiALMpcaOZvOcIFATup9GiHeGhWzyuEumrJ4qJHN1kFFrdPTaLeJK
EWwqKjhK6xDGeOlTNyHjD89tHKBloFmzHAIOD/8LdE31niAbJMBQYA3u4CnZKm91
9MrvN7vkcUzh6pMTDIDSl/UXI8mWOpfiF01hfT2QdF7xzeiUehL8REa75S6dPGB7
rFD9q24r6NfcsTOveAHQq2epW4rNszPqXky/gtIdvtGdccc4X3VMbKN2cQVBBxc0
+me0Ja0hTJlnCrN96VlvyhBxFEfVSVpdBnmGeVQe6EEzAJ7sAgUgJt1zZtZyR6NJ
xKpaVPePK4bg5rxZ4v9x+ZNsqTE0CYAoUZ3LkTdcPBwx512rEWj3FVli9Xodpjes
BX5vqUjjwuzccbvyfzrfReudBe73NtJKHxCsGCxio6c+CLnwCxTLr/VMDyvpTVQv
uFU4uDwgZFROTOxDtepORhQ/vuMfTv1Rp8QLOhqR75boFh9npylbZOUT+j+GGRPG
CGU6jlXvylbIquaC3Kn715R58+MX3/7Fxb2XK1+bfW3XSkqLheYRNELnl5Pm02cA
MSuMJQn+4lkRAT4Oq0n008rCv6n4imCXZNVvvEn/GGRShI7rnZFTIdeL+x0UeXNg
LX4xSOBGZQ66IR2s/f44CL/e7TG4FBxrPOuJau0RNCKK9JW+JU7Hz6Bm5jCLnJNB
TZEBt8acf9v3CT/eUYT6EUo+J4yCVMm3zj3f+k7GAfA5rW7rZRT0gwFp6NXeypOK
pLLtrnD7CRVZ95O9G8hPXlTLBbolqadS+dLxAR+GYrGmo6lH8J/EYZS2wMKTDG5W
DhHoGMnN4DHtJOTwmZbqjxBh9WwrQ0tTE95HiJpk8cH6NYtMSp8JtLAseTz6Md9d
qoKvcjhlPNPVguHET7K4TJR27rpXdBdD5kn+/FxwZw3e9GOwJmYtbBTt9EFQ1ogo
8QxtR3NJ1GkgPEXHKD8aklfIf0mO90x0GQoFQ0Ol9DAe9tn116YnmzpIHjwqFHAE
/jV+CXC4TYcMc0N1Z1QnpPvI/J2SusfLViFlm1tIx8xZ+8hFbuQT5Dr6I7MDcmtx
iX0jIlaoBm8Cc1j89mXCrmFy4EcJm3n0iSdBVooEYamnASDca48A74yv1JK9SLJ0
p3yO8PxgvPQMgPJbnMn+bnt/1KIVrRRMWp2qMTimQkXeE0cTkZGAsrqKLQPc/KZa
nxFZPqhXGJR24vqt2CDcJDHo9OEtkj5daXkAV4gBkXXDMxbTbCWiK/GStrHrAwyG
sHnj3+idEA80ManSFyf/d1wSWDp5+fimY2PI9BNmPLY9YetCrsOtv8E22Bcb/ZT+
w+qvhsJmNYYKw/Gh9YS6KXrEtWhXyxW2JCDtTNxMrSMaf1p05Yf6Ih0saQwmJGZF
NDeg0qWdS6hvftOtjUDrGzh9NXtLEzDlX8zTzYgevg3ALx9QQouz/z9QL//tSfOg
4Y1VemsdfcLkdC5Ebzgh7P6PT0c3piDfExA7C9/p+BveVBeNcIq+Nc3dEFQnY4SY
JK6Feua/RoWcw1AZfRJh4d9hhPO1qaGxflowyaGNx1OLFEQVtsRXLWM3+KfMSsmA
lBKmPTi8zxTDG0c9iEFcZHlVhVYgsSgMPlyURaMEjG0j1lFLhdKYgQhRW2+ujnuL
H7agG1pLQrtD8p71ViI6gMG/KO/CayYr+rf7HO8wdH0gMR+v38nA4q87WKB4oGII
fNwOv+bvvKQhYDKcbkxjj+erRl8+0GbT/vZj0VgteybWhwE65aF2FILlPRTsy6uN
Gj6ZDf60wV/MTl20+nNZ1M/omEqr2vf5lmhi5Zx1Jo8772o6kK5yYmwFD8sJmAnq
LC4oRWF59DAXU6EgMnAjJrMJA+vNfzE8wvJe3MIrWipQVJeRY5VGxBp/uJa5b2yX
qP2JLEayBLwoQaPzEo/WP6zN2iizxFAqi0BSuDkrXlZlcf8CMrqMNCpV/rH1DbxV
0cboqjnelQgPD0os8WdSskKeNUXvtofMpQUW9N7fXcYFkkwhWRN94n5Opl0rVCNL
IeHWyP68KTnqfr68npDh4WYHg6jR4eZUwaq/+nYiyIjq1V58naIb2yxrEXY23nQv
KajgtbcX3t9cgcoEhZ1ZcSG8p2Tz1Zhxjni9qRKWvK9YjiKNe3a6NsKIYod8Eqt1
DUOp159pxT6uGYwosnuJu3QZ8DwW9ew3kgc5RSjtpPOy3jBdOA3j+dTaDSdm5zJ4
gKyyCjPJoi7D8SdDHdbYqxBVFAvq31oDH3Unjzcdbsys5OZqEFdnTF1GslhghYkW
M/QlTG5xMjJxcOxp8tvyVGmzHWUdVtHd0m8NIZT7ZOdInwSxH/HyNWhT1RcpWaar
zQNc4iD1v6UZRvNRZbcZ7Trcy2M/rbbbacE4pk+koXZhVem9SK6XhnwF94Op8kUg
RG3NA4B2qehwwgNqsJu/7FzpvyVh9GCAKnWj9e64R8+kA/uneGcbns4z+TjkWs0y
ca0iFd/oFxUNdaja4e2wLOamhu0rFqqy+5CsotsgYt5U6ffhytnoOThI7w1orJ7H
azwce+dPGJXGg+UtsmwJ3vxNw7Tmhgozx7ll1aPOqPo4ytF4WKmYIkgWAXmw4z8a
9iqkweTaCsmd2KHnPt0W7t04mB35+3F2u/KHeNX/6pzQ+mUxypTyDtHk1FLK3wC2
YKKjFdfZQIY2Q3cwPwTIxFtzaDzcJpxxG3nMGSABc4cv2w1FCxkmbe4G+VYInFAt
MFkDsV0xjnuZE2eTdW0l0R+74AF4fR5pgWE4q3N7REkV9PtBgr0326sIlwHL3zP7
K7N/6p7JDCh02IERqdhLDviQdCcqB096Ufzqc9yerbJWQMlvfxsumTEZnFmwjeeY
jqm95kUhLey5htYhjIkQQDOt58zrrCbekFsdzqGpNJiK7WrmD9AFYtpSZk9WtMTT
pCwj17OIAyYAaC/OHK/JhPHOY2bMMBHRugowGMQ+KHwgznMkgJ2MST1CsKF+4zuH
9uy5QkSnBmBS34eGI1GtaFKWYszxoGyBoRI3TSPPfbptw7uXViTCYBuU1vTSVTc0
zQXO5DjDWPVk3/YhkZS18yj5L+fbJdRQHVdpi58/8ZIRbzjWFXp7I+A2dDb68+Tm
0tMbl0sd5blkHnD5ulM3nnMsy5qTN/QQ9eEb98RypQ1QckgVYRYApBvC78ftaOiX
90xL3n/+uVZqodlsQW2xYHXa08fi0cQll4UaVdpj8WxHo+zLrtG9w2ZGjmGI2fhq
9yJGimi/4uZt+zIoWUY2rgu2kQZ2Xt9sD49t5eICE2J67w+BCyTpNW07/E7YJsa4
mAg+JsCitlv4rfx8rq0ycX/5qUOnXfpul+UyUh/gGp15iMfgZD3rCw/xuoUUSD9V
H+fwAfbBTriKtbKZongoTvOR2gIgEuzNdWutcSWRQfshdwRXKLx0aGFRsTxLMm6E
t2j6Qvneozr0iC0gppE6FaG879MDUbCs40AUWtXBB5ItH4EEqxOeAT9tCVcfxhmp
n8+o+vHaBeFo3sorWJ9ekfDBSMAz/4SF95wzAXBHoIiFDU/HJU6ZLElxgQIK0pM/
iBGOoNlp2SrjNGWQz8vRddXcLp/0Wz3/+4omEHllTuhk6tiAk2CmUiATAd9AreKr
G7q6+h86s+2ERdmSmzTd2CVpKlEXynp9ha1g6L0ehbViXYGKXf+ZovP7R5sd9f4c
k7vlGTZHbBxFRDT6YUB5M/ABbnzkV8QYf4YKhg++CLPKAq0hB0vIyqiJpYfMZ7fj
rF63Al0LfY3P821OtP/LL9YwVGoeORvPneeiFXil4hPG3GBR1U/I0yHb3KFh7zFy
p061gNRVyEkB3Y+Ur5/nglMEmnutyHRO/jfkG1oTvy4d1RRQlrF2FN8jnhtXs4ZK
BeRxN/1IPxskb76oVEVBTorx0g+DFSjNym1vpGVIoHhUd9FADmrgYAkqapvkJ4wl
ZtoXHBOIHcvhxDPTIzDPxhePyPPiuLPHS6c1oeM+7Ce9Lw084bh1R49KFRxeMsEF
OJAZjXHvFE6MNFs/V6+N4kWdIeNdQWn/ze0NFyOzP6y+5pDNL8f9K8kMdrqSh/K4
Ev3bhL/zgg+dVb6heZaEXEACeJ1ZcBvKCJlynl+ZPEj94md6g5xMDOu2Db/yf7Px
xgBwaCg1xrCmZDMcSpRVvSHQgO0sPmhz7xQtpUH6c1PUBaPzwzSxHlEOCurkTWiq
Pac+eTieMP3kjVRzQ+lJkjA/8el6H/tBAQDbGVRFKEFYH4ATfWUL3szzRV5Cwjvl
SmZt0+IuA7sTUSm8J3+cJJUfjBvUAJlU4oRxOK9n3mNT4FRLDFPQ+w93fahzQiYD
Ael9Npde3UHcBhp3gvK7/oZZPWJIZl//Dp0WOOWaDVma8RrIid7mnwVyQfz2/88o
aoDFlOpC12Lx7vqUswCyszec8aIyh20fSNm0SuEttvTznfzApAs+F2LDXv+b2fiv
rv+CLplIUBBPRhD8ed24kH2q044djxCc9+FBbPBWILnEo5XXL6TUqEjkmD4IiDOc
FBmWm/Sh6qb+spR4UH5q9e9NpnjmIjy5ow7guns3DNnWExPmY+98TdSoT+CKYNy9
YlsBeSb1arqIAnLFTJXj1nNCCkLHxuqFd8zlHoU7/f6IqCgqiBxGik8Ld4ol13sq
wf1il56wAT90n8iqWzc0RVNDO0yD5+bSY5Z+EbuQUZA9WSo1J7DiCmORbf/qwRKu
1OullCDMLMVizue84B3VCNeGSRq5b4EQPAWV2/RuuGFO6pxo4RwQ2EYBTx/rYLIu
Msgm38LH90Q3jNELfF/M0REoNmrhY1P3DUezkuGacFLKh5cXfyPyupXiafmNjoGl
R3BaP+AQB8DBuZfByq8F8y99qGHckzJEQ/tvEGjar4fVI10gt/KSJUQPQ6cX/Jfp
iE/Ivh+wiaPgQ7eDvBWbr8V2yZ/WCBtBlhGcpqNbwfWgvzFkj5RNLOByEed7ElCb
t9unPLH9otI/5FlFkOmt1H38qKCxEp085GYNGlzFgJs7oTqDXrve2B361qdhhVnN
yRfsO9CG8i3DAtzSDw5ehtGJpANFMSf4JpIknkxtsHMzgvByMRTgnabMzcBjInik
RI3ILQT7Fa0c6jC9ocPHvvhVnOW4b8M5d6sCZL/IYG45+VlQIVAFfwBjT+oy/LLz
6zurVZm5ooWWfiQ4bVO1qKtkhU7jniFlIlLHJzlLD/i7YIeOjr6IOCpTWhqaluAY
eyo2MqwA7l8bWQCF1Vpgy2gTW3fHsN43L+qMuIp4B157eXw4fv5Ez881apJK0fAe
g6y5W6xB2NI3xRZS78dJHqXwPclK7S2yuLckTHAT7IlwJne/0tmwh7EskiN1MLw7
hoPhV8tQd5oiOmMd74l74XFRJ5wyer8djS+emTDHi8sIWQw7eGyUMNgSQGidEmfs
KWH4eiihOgKlSGrkIYtsjA4Mq/AWsO/Q1GfwyU383Tx0o+ehozLE2LQh+6WG+T0H
HRRZjiMyQ0LUS160n6REj+9fdJ5Sd94kJgP03yS9r3uFJDAyU/561ulO+Cfr9Dzt
AHsypRGG7cOWwZ4KPZ5VGZ66QOpZXGzZy6Eaw1VqE/Jp92PKSbBmsmsMINChQLWl
GHFUWVDiMcZ9Br92TlH9FQa89gMKnPmfNkalHdz2LBFiBJx9XHDoXrkeHrHelTpr
xBOdzNlA6n2Qb9TgaI4yVBsXPaqyIR3CjubkIfIJH4ImxPeOiifZmNaIU5p0Hubx
RPspayoGTG9YKS4TsCMgA6bJPt5qvDmPtX+w9a84rMQv2KixXYKQtHlj8MU2N62c
wKwFrxindVpOyEeN6gJ1PaF2mGObnfgi3gV7KbUXqfMKII0x7EatPQC1A43nl+q7
y0abAhzB4r7Xlko9/FicsUWqIcarpu75wKuwcIsIHCzqATAbZE9Pu4fz1wj6r/Po
epRaNMRB13sQwDiQWzQVtOLFtjCESuz6aPFDRIMevw19O5m3TYFejGHzRdu/s7/l
sx7wRHRZST2iv/8N8QnZpo7dvW+92DkDzaw6SD+WDZtJ5E5QuyEoiAIdofHSt/VG
Mh9Mr/fX49KA7OgLaQ8yihvNwY8CJtcufJGbF51fm/SCa3qGfb2oobUSy39ZenBT
Ns0OjhzxKJq6EZEEiv9MTHGglCjAvUN+H+/uK7sX6iRnweuRfLshj+qV74lNQBfM
x/+DveTyPM7m4qfI5ANtz8FDseAgVCWrb3xijGZY2IjoSOE7id/etJucYyPi/gZS
5HCmitxpLqJIbXkXOg9wN1OvUdpXgZY3MB98l3nD1ATwRi+hSglhTdeaTRzM4dah
2ZwEWg24oBDO5BTZXnwGZLIfIOl4t+t5WCLlJ0sEyXPpbkdTbC/X3M5OrapqTOS6
d29mJwGgwoxdpuhyQpCGzAvukfgGpuqJ66DbwI/S33sUqGA0IaexpXJXcB22GPi5
6hvdCiw5rtJXAig3oHH9AGqgu3qXLF5dAaJw4iMjqT7uNJDOLFiHUOYLIRQAAQ5U
jvmPbRA2rqSGDi/WxvYcymJQMT8tXnOHnVcaboSwulOZaFci2ZmSLrPubrHymhxL
PTMTq3lN4NznFOUf8kKbgOw+qizELYftwoFVF1IOzkHi0KPHuMjz0fpkA8qY6DDD
aaT1q7IDFyklZZJ6IaOOPWtBxQrV/5HHvEH0f31vwG7ARaqJipvkqvhdG+JVZIcx
UtuynrXBv5mhwrlYsCYKllJyWbaLhyEPDsAarmUkf0/6VmDQC256xVJ+altMsmIx
n8QaWNouaEd+6A4aN0tw1XK1IqJ8sC3gFGN0I3c5PURHVwJ9x6unYy77OvlbWyxK
2J7Dk7FORv8O2OPAppL4Rh9enqYx/MLWwj+v5Ouc5HhMoDcDrZI6eEX/A4d4XUJN
rub+Sb2U2mSrEVjV1j4Md6dgAcL+IrZbzq1/ac+AtN1mp8dgKfFPV+5i9yNYwuPp
FUTEBCKFQlffQJEKY3Em/VlTk7TMES83Ly4T6+TSlq46PKw3jL4D9PIBg5jsWMNZ
sOdf3PgIhA1pxvr78U4cHo7++bjaJV+OQuBDEkPx2lnMdSUqwbJ/7Ozj5bEa/71d
yBC7hqzOitIWlyiZY2VAb27Qd+JfIiowQGcDMSHBzhGlxu8nX5lRJzH5a7lrOEs2
PUtqospMhS4Kan67s1nxAZ3y0rlVikQeyWBAC4KvrHOe0vP6gJ/RcoPcZ9SDiFAW
w7v7k8jMIDfCdVRbZPKWv0AQY2XxUTBMT2mwpvVZoNqZ7u67S9Wdlih/z+kzeZQv
VBdE9rNLjS/RFZOLUvTl1fkOroMx9P9zu/ReZa1sPVHdb/ARV5keeqULVUHoMIKg
g/QvYlzdJsr7elTZErq5uYgapY1JhgjQ8F9zrUmIfYewYsqvWLFf7c3zwbAVZcw/
IHOrc790rhPurCXb8VNuz9L1pFnQfgJYcT6d5PhxPxlM2aiJTNLK2uCdQ4JlO0Bb
T+Shdm0nPwmhRKpNKIuNpw6LxOAuIWRdTOfIikij8BiZzxb88o0HOY/7DfL/LwAl
DED8RluriTRun7N0QswPJSS4Esxu/EGqK1BpoqljQWx+vdRCExTYb1SWXSUMHC1T
dL4XRFGCR6qTUXiJRhnUTEBRsm9/J2yJcoTiV9OXHjkwy/Ry06B/sM/BaDlx5jvB
ui3JZdXZfgrT6t6ABRzIjDiuXzc8HlpvyKXSBNSfftlYemsuN7nruVQQGUvkHX9k
fXSCOdWBc75mYErbU6qB7pgaLbu6BnegC7F5KIQ5lFoDLJbh7AUkiLbyVo9RwXi3
+UAY61ReNAIhYCyfJx0qJJncxi6X8Ra5H7oUu6Enbipwz9PMoQoA27FTJrMju1tM
Lo7zc/4ZBnpzAEgxs7K78i1OWtxYExEkeSsicw+rKmZ3PRV2XTd65EJQijSax1Mv
i5bILb948ETyYReGhyLydKeim9KaXPX/lMK0KiLu5k46WxVPcP4zSotqJP6Fk/aR
4FzCuF2x98PHtVR74f/ISo3rWsVxm0sGlwQ5Pt99wBcwMWAo1peAN6+WT2KsgnFj
3YEdz7x/dBNgcfekF4NgxBlJs/eUaCYa5Fgb1ZHLTyTvKtE9YDxK/EiH++cBCpA1
zlnlp9PMcmjTPtNCRwkXymodp902i7T5XQ17Hzes5oZGHlf3P1AT/ALnlGFN9r8r
vYrPkK0FbOJLS1vf8ytr01c7iaqbx5Bj05+3/QINgWZHW98wITiPl53sXVII3VSx
vYxy5dV6c5tI0TGhQa1YNEES8Zg3q2cwGhf1w53MGmj4fU8YZQS2fK8oQE/1TVUF
3yg0AtgM/7Ihm1+vDcX9CJ1e4ZxeBHnUmGa5BE37VSCaJepHtBTmox5LubkrePER
xPtfsRNf9bPDQ+qikTeFKdnL/b3wKSs7nDafxyM3N9cmXzIGHyj+4y25h3HTmBSA
qM/orG5U3HKT+sKdXPj+DJvU6v2fk8sD2ef9v/i9YHAIeHZQmzwZhZ8bsfH6gox+
T/AAb7OOCyWd8cD3y4W6GjdKiBBaj3dCbWjG1WfPZ/ErqhObjFBgBneI5zbbaYpf
8n8v8YxjJIrKRlWWuBMhFiKe/evfVQsgoj7Y1qT2SPePPqnwj7WeBzZHhkG+cFyi
A2aD6BkO945Sglv/8Ag8Wdz2rMn5UjFXPBcyJk/PsAfLVyT+F9ETwq5T0OyOcJiv
s83/KyZGH2+0v5dYPbI3yeocQty21oiyekeTc1bXqqHS66+H/2CLIcqyqj1wjYhT
f8XmKdF04B6AGgv1O+7Qy0MAK7P3iSaPYyqW7LPqKLHL4Bg2AAAVcbnZSzpiTCHq
O1cOCWjZmRUUTyRjqRrMs6u3Y3OvFGdUfj62NXg9eM6KI4dKwfQr/sJUX/MrbUJL
iofLn8ZDh1cFZzAhj5PpLKtRCKGlQsVB4Wc+nlT3wbSIg/Q4dS+9+tMTMgV5KS3N
f+qAn57yXDfykh5uoqAaUIaq357mtibrSU9P+S6eGh0NnmgOk4CzWDrX4igjjyPO
fYpeamQa+3pmkpK95qKaBOtM7kH1ER+RE7Y7fJglKIskzFexZgbb4uN2Izm7k9Tr
3R40i3SMloV6YFNU29DbVUroIj64n21V5B6p9uI0roTdpwYZKuwhhaxdA6gYqdHS
/9ETYaTiI76bOybOI0nuRBsRlMQ8sTJl1XC46ljnyGq9T3xnfJ+Kn7+z711ir8Li
BpVzfDcHKvKSjIBbouCXvDVQmvlwhTJkhT+xLufQE04vF0r4wC6LytC5tbrkZ6qC
D9kw4e+/e3/6UZOB3XywWkvDL1308ZlxKZRTgGTMA3Wl+jlqNSidQKCbPAatGM/N
OuDwibbdImEia+b7Silhv/lA8A9Y2Q1ZfSq2mltj2RVLovH55rmx05Tbbb45lAQh
Ho4qgn2aTLsmlDGynPMJCOy2tHjE8t7XYZ4F69Yo+mmts04y9ZilkhYZgGIR3A8w
B8LMp0fvbhtRLb6tOu3xLqmZW5XO4bSWLv/lZnjQTFb/YZ1g1xmCKyDh+uX8aL/7
ZNSN62TdY342BD/uR4q4m4NR/WIogscIqrhdXyap5adKm7M7zHprb9UBEy8YWykZ
VQhbq4GaONzZstqqvzx1pd2WJ3hG5jIdt89b5wFFTz5iTEs2HzbiDp7h+UqjF6j1
0g33OOpIeWXBUIBYheFbd1UB7s5qKOUrtvjDNNkYO1hwTn/8kpSr7WCAEFu69Hfe
0naRntvSltICE0VxmwaFb5DXV7pCDHPRWfJaQX8FQBS8Y9d4IF3ANvdEInNHtUjR
6m2xDKoyZkGzLs3MnqurgsIvfL7wZj2s3cxS0xj466D44aZiWmEkly6KvlcB8loj
pUuVhKEg74243QJBSmp2XLD0G+h2rUf8J5imcJuLoWLJyAU5ROLv75qBqTTPVJkn
1xlrdWcGMT09wIXp21bd2SJ7Y6osQk0/8ml1wqFE023tI+bc2Hap/nwzcC8W4Hbq
gnrQkK+j+g9mp2xRBuIcVY1tR/sx09pBt8/ZydEOOr6JzyOWkULRwSnxLTolnMpS
D7JhvxMzzsEfSUCfXfcvgACT9QWnciE9GUxSCBsE5tAmtG2V2qS78L5lvZ3CUVSZ
qxnKBHQRd3RSVK1AJ9by+Bi/ovCEBbcKUkPMIt0dkSmogOFW4EoSYDCdkm38eRM4
2SKXT511aC+4vi/vab+ElOfwhzOP2R0u54NpSVrHR4PHJeV1zK7fS1Fs4eTIay1K
TH+o0VOx2Yg2bR7pHlYk6uEnYNKBLgIpSI33LXi/BZvuEUTHb6+Tn4FzWsz9Z0Lc
YrZuWPlub87D8BYwUl87483Cds58t///RrQcF9hkf2wMfsFu/jNYb0KXvd0Ph4qf
7DWV/9njai3IZ8xUY80zfa+3tFdPjkmX+xBBd3ANHyGoTGVOua2yq5X7KDMw73w/
mP3cP33Z4aXelgfaRe6d5wF2oMnvIk7Vl0AgoXcmGjkRLXzEgztSTmJH34lhYF5G
80qfsEl0v+uKJmF6riUYUs7i4gliPyEOZXB20m1a9cJaETYy6DaAq/5TwtYpaTk+
REAXcny0dUrdcBijkJqkPdum4PDRYePnIGDCXKgjC1GraXJB3ew8qJBxgLFP/VhK
jmx1G0oIdp94Pxfrcb1yANjdHZTPQt7D6wj3A/6FQmtrXU7aSemw5uNEP+tsRvNT
KVgNwBKy1VMiop/6ptou+M6/JeGadt6RYrxKUyS6VlieFrcTu4x/8ZS50V+BeXsY
RmsicSJuyYLO166dIzFs2T3ZVEuTZhpBStMKQpHuUkJOf/dau/ivVk5qcegJAq6s
AjkbMWkLkhOZpFpocnL+s88qDQbAFxMbaZv/JxwEvCf6r9uaGbySsVaPboUkWVAH
ANr96Rq65Rch9PVS/a5czGUNwRv06mEtzaHoZK1wadIiqmanceL71fwP8/lgqx9Z
pzhX3onwf5H5hYfX12SKS3OqsCrcnsMILkb7ssuAjVZp395U1gt83ADXuJ01J+cL
bZhM/9gxU1Sa95HIfs2CnEbd1f41XO5Kwp4IZ1Xe6xeqX8HVwy3NZ//KpY7wOu7R
GZRZjnB9q/BdFgRpEdGMSRjUXN/+8EKi1nRy8v9AU/VeRwIsEh33aGsCAHgEWrut
7x4mIIxd7mKQdf3+kwu8AYQRNU0pm2aDYtMKt64UxXc=
`pragma protect end_protected
