// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ogupK2RUFJ3n3QVhF8OSBM8YqeuXeTDQFipFT0oMM8tPJWzPtWF3rdhm10LEQ+8L
txgW5GgXtN71clwVg01GQzvC5EKt+DsaQJHpCvprSI2jig0sBNF1ERi377YQMk3n
DOLjjUDTunsR+/JO0jN7b6fVHX3pTkflR6/hmQfzI1Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9328)
QqlDiW0QPoBdwI3r//Fbh4ddbFZaoMdT371bca0E/7mcx8V9gsZCBE0nqFigEOS7
1W53sw0ZYq4nCduJ8RFSdMitf8yRUMiuh+9fRjmg4YQ18ly0IEEBkFPHCIdkVgDe
7QYmlDLOqwxmzZRCBFCJHKuKv9P+zT0yuI2xQvMhIGf3wN4lvt/oudh9azWubvjs
LL4DDJHWq0sBuvKK60vC7qEXj0k8GImJaTijCCp4ZuHVdvs9ga8OLVi6ORq/j//S
UAc7ffsIcuWmfPmXalh+fNMB9/wGqrU/4mVTdLkAEX3c+1IT0vFO1g0QY+T2+v5q
sZy2mDtGMYcteCWKPEgKbzokgYYEQm0CHWZ3AX6xVuvFH/uQhdeOaODW4Za9wckq
W9QmDKRv9PKVG+LVp9vFS9R4vtz4jm4TX4oQAH5wJu19tIRA77CKBn4s8fAlGJcH
ClL3jNtpvWlBZldADsvrHP81tlyolgEJW13eXkLn3LHP1Jd9bI7/Bepf9LASDPsO
MGOcO3lp8uXYKyrLH6enbjdGfZQBTMPQG4gRsE9yGGUqQZWODqZ76eoFASfzURPg
ruZp5EMbDSnCzml9Adus4I/2c56wILzuQ7BIW+Z6hC1no17pFh/8vHeTInSftli8
XEX8vw2zO6wiJmBlF0R6NwPQMq5hfWN6Jjo+C3jtOJ7vcNniX/ygqvoEVw/kBpKc
1Xaimv6ZEFxFt2t00n22+tCOqmoN9Ysp1Ur9ojaRiBc8ArdF2y5No3rTzdFWas7E
NGrvrvF1QJdc4c5c5WaaYppoaRuHMw6J1adWeQaMu2mhwe2UxQihI21lFyV3p0So
k9GjHCkx5UaLK0xK0WldKRWj6saHSxhQH96xLJ7C1fPEYCXBO+OvU0srdOqgpTkB
kqtoUmkcW4pmiT+xifUuKkYsuf4uvRjDu91pEnP8JylcI57sAPzEsl0gUnBcwOTa
4z66chnP2JTZM4mrej5NaD0MGeXy7lMzoHMaGnXD/WbiPrHM9YhdMn2bOnasiv/z
nyQ7J9brH/W8bZbcWUiQILAznLZJGRghaxI+r6bRzc4/s8z8HnEbu9/TWns8d72L
Ukh2pTDdduzrJEb5CMnGU8VI3S0Mqe+bzrRetCCw1l9Nib0KPlcGKDN6PXOFWs7Q
BF59+wxbZOMvJfKO87cRzyB77C3cRqp68IJxfQIJbw1LJgo3OpBykdA6A/KC1IKo
mL/p9kEhNHVNhSRs/G87YcB8XakMnYCxf+BZZOoLqoLO50p3yAPnC/QSH9xec9vq
BugjkyFkmDHSPDIh3qCYTvWJtj3NnBI3vluB5vGuKfOzXG9SpWyyN2r3AQjNlCAA
or4UQQg/bc5pefdYRIc0XY2l71jAl8ZxYbJN46d39qPLwWsBqPLl2nb1a2Ei64aF
UczPlpzKTf+j075VUF7hdTWQzbyBbH0h7s/4wW6IvPnwFJ8c0hXjsb6VVRLy05LJ
LQvKBWzxx1EF1pYA1fbR0YnSk5Vzu/zKJjY2prtBY1HXSZJbbHHv5HBaO07v2BAt
xNBI8busw9DMrT8tyj+DwD37gDUS2oDWsBlyYfBOLjWAsbUM4GAVJ6RPqNXZMmqi
pf1tmE6PUu7P8WxafJAOdnZyPEj6FIQ67fJ8/BDY3BahwAxQZYVz6m4NlXfF3n1e
CISi3aD014B4nq7OOQNcRyy0tPw+oGcC4GNlLR6xeLWu2za4yX+T+gavWTixoBq6
flB9RZNZzeKcPtp1baAOo5nhIiEe75Y5L7iLlRoIX2/4F4Vf20ScShGAm5QMC8Qn
UjneRlRCH88m+WzqGkK0OpdvGVGVJuM7VEB8J9TWY6zGF0TO+4fqP8Q9dM5hsFkd
ST2HtyGJ3M0DMYUZ/oQHVORyBDajCLkd/yUpZ/EMs1akhmMZSzh0SWY/ABeuRpRa
ik1veSj1XS1HcnsWVVFnGyW18uqcT3wJVXS8ZFSXlI4FAI6vWM73yyoIfbRLZNtX
bzCuReH3AO4tzgfwsZ5ugn13JV0xp2Ub5ecPVwf+hsp6E+JLTxAKkIyS+IF7qhlV
ivqCJHxH6qbZE1s2BgVV09FRbmkMtOWcs3MmI3fJbAFv+x4B24xTk+fRfqB0VVNR
LM2xM9YKsl6oDmN2C9ql4jtP6BjxQqyJ82HmkaiopcOgTcnseMCZnURyEgnU/s6Y
F5krzQKHUT8XiVK4JIqcVKV0XCVzqn4/z+P6iKEfK1JUObeJf/ltNv995Ttz16Sn
mrzBtkTUF7g+hmg2f8dQBZejscav8umGMezXFLTqyW9xnWEr7kGFk6BPwQVzaPil
kVr9CdUxdAajqJDyZ4xViJ39NqTc7VM5oeCK+hnFV2asQBQqGtdIA7DLoBRja5Mq
rbxD74PxgdnfSLBO2hdkOmeTAt4MzlqL9iVbza+zfG3wml8w2gVqsRSapGF598y+
EiuN7pQJ49yL312+ICtQda0P+Hhz4bkmldMbUnfG6ohz8mhLhoBFnWYk3nFbTbgT
mm/3RVRlFTgtKuOjATwBmAtT5vWv2xMoGV/3Vm8/GvdnEN8/SuiXUILyuJ4/4Hyx
rkC4iXmG+ITRZHjOykAgGtyd+P0J5gUdO1QcTuomGCju/lrdhlES6e5OOq9CJY8l
2btvb7b4olYM+m0WfLSEjFVuwZpACrdkYxBwhIJIZm7Gdpr+6sV03jgaB+JK7ouT
AuxtKsZIpdjwZ1dewvXyCTb3h4XjUIU3sRP4+TMzwICi45u61eAYqaj6Im6Hj7jw
j+HbV5mEawBpmmP+q8QrAETtq3GoWHL599EuyXf3kG9ZqxTYuxJ2CznflpJJLYRn
mL1OiCoPYop5D4VtrKkwS/GjJNxIDHCKVv2l9taMFGhPA5KhJ5mMiUrW7rxDDhK9
dt7A4xyJwAkDoERWQmTVHrEzknSxa/uW+AvYft5kGoYJ3b4zDJ+shsUwdyJ/X1L8
vUpFs0IhmgfXz2PU2w/sGzheD8z7EvQNVyWPvs6iK31jyMGj7rQfuqGqinKtUeZ/
DuIc9KUMEM3CRq3nB60tyt+VVMDBIaqla2bxERFWB9HBfPD3vRSo8Gvvtu+X7xJ8
IFwOj17FRFtu0lxBtygnTTOm46B1U7A/rcodC0HBsMw+XgNyObc0cAloKQ+FuPSD
R7fO3qupgRP6K9LB9uX4t66JeYTNXQIrgyv2UfIdmUCjYfM7LkFzCLds8NhQ3CrF
VjMNJ8A8r/TYXJx7T5tdbo47YWMBbQkv9uspik+/5ey9wco+dwb2xvej2Fq6QqWg
F2VsKrofPBAkJsoj+XUvzwwp9VGNsIVUFO/AE4EQpVHTEmWNqS1x8HvIBNWwyeEV
QoikkfZtUrLIHa55wo2p0stLjAnSY5sLxeozcrEXVCbKrRCUFNXqfM1dtUJvQ/IJ
qzIYdfdGISD6EV2TdhPxbbPeNUHiSUzQ6RDmOB29bwxIqy3cGxlZRLi/t9Gd7Cg2
KP5R3OCKz3ekAJbwD/nupAF+BGOfoWQTG2QP9nXnwgYLotk+6eumPjP7pFRyhxWu
a9oDlQ5l0oB+U4DLujncRwr0Fdksg7A68BWfyo1Sxz1NdRUawrCw2HjaR/NgYSjA
1+mtdIueD9h37MEneoTtyX2lJ/RJ+O6CkjYFC1a7C2RhpKmKddr4lAUO2YltzPnE
dKC/8HoLSd8vd2nBMBe5yTkDQrPjtJz4WCiQsWZ2dwAFBpqPR5WyPGrRDB9jCzcr
rdvDk1bfa8iJwTsFk6VEt+HDtrqmiqEx+FOvfvR4MvY8sDhenlrFIKC0A+8+GUPn
UcUCigKDtK0jIPwQ7MuKZvb+KlZscgoCYKY1XboCJSCpXZKDVp4X7co9vp6OiML4
aqmRCJOLTgGggkIxeHzziDB3NGCbp3S0jwvH7ft1suiqBXs8iQ/eDizT0Ovd2f75
uUnxV6l5idOVHxvFI+CKnrktkbLMVb31rtGrREFjx8Td+l7bkmX/LCeRfLtglUh5
UwKlbrWhdKmuJYzSE2/rYI6/daUGFd/BrnQ1Ua4UoiAVDflNn3MHqvYY3GvfY9qi
DkF97F7MRo9QX/2B24Cu4IMxsE1Qa5uRGlR5MKroA2Vg9mzO5+mm7AEsatejhyxC
tR+PTvS2x/HSoLuAcUNYWFuV+wgrzXmtddaaH1yjbWgHGJXOmphLtaphj0KO7Cvp
d4NxXxYbLX0zUxF8iPC2nAt1W9uh8Y74QCvW3O/icS8p0uqT2+mpSry+YTbMCEQX
1Hf5cAtJPlU7QL3KF7fMks1meyWm4XC6NuFBDdvMxNBmWD4r+kvbOkE8j5NCMdGc
CJ/L9JWVgaSurv35RLoTOQvrF+6L/RqLQopicSsYmdvXauFykCdFMf3Uz8CcggZZ
CKuBvUYLlixGsIpcC106f64O9XdW2BlpGxavVP6UgODguXf1IMWBDotRROkIG8SF
BKqWEc/UmEF1GGY2xWCrTJMc5R5I2a4MrbKraVO5cWa5qXaFzLVxnW9BAf3xLGoG
uhSskG2s796JxKNT5LGHtBBlSZcc/ISX365sHPrXw3qeUnj5cgNQ23sMMzH9/xZM
qY2w97EIpPoyk8TTN5+4ZMWedbBKTLyIryZV0/z2+yN2jn4LDKB/ZL6YbqdWTCXX
P4CW0MKKaXg1kgQNCg01SAHjMKaYs5kMCMsOjcraCxdWlnnDI3L734aPm6WHIfmx
xWGEHdSv6DcBukxe6eoncdW+NP6e5+FjlXz2Fm6HeSDXR656tT/pBIYD9vChXZ0T
wqARff7jH3f2i5HpvTYtF6U51f20pQjzxVoR9vUiQtY9ZAYs1mIcOpkqzDuzkNS5
HCl4XN2sJp1bSvZ7PYQye7wx99Q5CDaN0umpO5uz9iyKHGoN8Q3lt0cAFyP7Waoj
tn79tpr3xg5fhpEWmFHrxsyeBiJw3w8fOrtkrv0Q5XQnUJnikAYD0voHc20GYya8
WTjlnM4YDJxhPGV7VXfUvl2xCFY7CMKN9BNEYe5ceCazOMRC/6e5u5lU+BTwc0eh
jey0NjlyZNnda8m0WDqBDJKDNJi1kZLjgAxOm+9IBrg52v9V6hxS1Orin1G4p06j
+WGM94QwzOCTmlEkFWyOJ2XXPtyMz6TDZrurnY/K65ipz4CqvUkqjtBoaeIUMx0a
gsXSMK6U85KpqDbx/8xolJOKukSd/IkIDBYpPY7LjoNglfKigKl2jp27y0amZG0k
2xqX7c0Xf9Qdn9Mz5xc8vEzbyq8f5yfhRtAObDu3lVJgyjjiWYW+lRpM5yCdII2Z
bCsJmvaE7lQo+RHcHDpTWJX1FKHWhVVE0KrBmmpFoioD/+Ws2QOWrymfBEo3p0D1
tOPHx9K41PnkuCUb5LHqAzFtA19s06QLhLq2S7elZ5h4UbG0xqcIbcNi5tifvKaf
xAmg5+Kf9/J1HnGZ/l4kAAj425YZ6xyZywuE4xb+2Pt+XekRkzaTZLeihr3VY8vp
1ePmg5kWMKRkDj/vuLbbASa6JXdeGj5tdOV3hlGWbcsmYeyTcynkCXfNItJXRYqS
AN6w0Hw0eX1Td54aUF6PjgpklajCW9bAhj0AzVuzR58uHBjlyqJPP+hFQxlOEmYb
Wgvv6c4IOX4fLz6MaDmNCngtc1fgmp+k4oFv9l8Pc3psLl6b0ib1DPp6lqooHc32
U6qDjvDIfX8UUBUMHlYpKmeLZHpdpT2xgfMeYCzrHG5DNoHXDtLChPLVbiX77Onn
HGTqcE4o/O5exRtmTk5cgANJPPOifOIweN9iNq5PjVt83GNfV0P/NOQGdSfGMxaL
IENlcv89JjRzYW61ctOyxmEfWwNfXHewonmYEvLzfR3kvbgwNjiOFc0eZwnRVlVd
uKO/oEhhIPNWzSXSjEeqAbmMxnTJOHiKh+pXICNjoDAQ5qi08MYf/1WHlzlgJgxV
UvKrkyPzj0MnplU6keJIC/MnQtMEa4b3h/0vHmmoxYgBlPyo7Z6CPjaNCjD3UpvV
7NG4lE4P3Es1hjI8tjoSv5FJJrtv2CWEUwNpc91aNigkJ0qBgpAakpjUG8gI+CEj
hK8RhUc/8HVTKcsbo9/AxNW8vyCvd0uXMXcX8Ed0ZV80z5BDP9iOED3ttkf9MaMn
xfkQTskeraVNenTCeXULJbRFAr6bEVkfm/OGFP7XGFX9/RZVHpqc2PZljHaAni1g
5hNf5/2mWgShSyGy9ZYZLqDHQyVH5DBBKjVQrSOM586qiTFObu2ikircxwd7/qVV
gMyj/Aps8r+mXH6WtW48+XjIFhncSkb3PxvdEX9s1Lvx/XzYsQhe0iYomnxrh7/0
hVFBnPfWRxScPVdyNz8yLGha9CMXzYIWOUtoYBnyF703M/P3jrGsqpCMsEwHIGYG
bTtQJZWLZkNrYuGqPJ7KfecZXTMuPb4FQbrVP7KxGAgSZrcfSoxfIVX8aaPAEgIJ
ehLz8xRml5cfYLZDOKO1fsdMF29fWNT75qVRsjcnXqOJ/OUTx1wkxiAdNPVyw3va
4QUhfqSnPtubK/yGc1tCe5hle7DQGoduwrqO81ptLaKBlCsIcgVLj12y7aR/v3Hv
z2SK4Tudk97advimEeyxPwYxcRy5nMIzmUpidSzCRZkMGGrZIo0IebgdPQxbO8Ym
RI4tydyq5hV24eK45bllrhJh+fBRUwuxIS1GEQQdm/zBB1L4zQKOsnb9yXTHH7VP
yDiA/RYlFm1NIJ/JU1hJYT+16JS9z++lqud/lmCRh+Dh+WHXlPfhHzp2UbLCc5ru
Ce5HKxclQFtR0tCAujOXW1a+ZF5sj4pPRr0wqJJGMUs/x5yWXay6cNh5NT/9KDgd
1Qnun3EXs+w4hZfTCorqYbXBTrOiS4nVdSJ9HqD1lar7wiE3AKWl9pZUVRwutbYo
kesahTwKTrKiApK23UOlBfzDBE0uBHh2JNzq9KdB+s8AwUR+qwCRnly8RVq1WPS0
Eko4Xu7krjC3/i6IT/gEN/OCCpkKKfdnm4taEmiCxpS8VxSGkir22DivDfiVIzd2
axent8wRiSpyeeRDeCjSZ7Iz5PTT1ZVVX7gVgY6Tv5vG73eoivIrL6a+LDEH1f7f
ipnznl5TC0BtkL9yGU1yqm0YVgO+U2vgcwXD8e9C0j37FI+cazTfW7xYvd3aMHSG
wVBrq5Y+CdGB8CTcA5c94iVyt8SCTj8GD+0K6DDF1g0czUlrnaLimjcf2ROJNYOi
gkvj/ru2KM5KSdmB80Bz03Y5xiP9amJv+1SLAz6ZPuuRQ1CeAE7xDWS/bFQofkq5
Jc0ysBPp6Zr9u7VT5MziJ5ClBbX/SH+Swy48hre/qcaZfryhBsReYJWX/riGjv1z
dcjAYtkwa0QDDNyoAIxBq7SK8foFH+pDdQLokgPB+AGPEgl/LvBooQ/o3JIPkarf
HSEbq2wRfIPqOzmTQI6knWxRtGgJw9ltQ7FKTIh96uLLTXOs7BbltM/6NiOB2P+m
4MJ4kPxy7pdfVvhqMo2BJvOlUc3BEtIDX4ec0IH6sFms8t4IwdLHkAP19b/PlAZh
MQFRPJXf0ZdQucK7NcwFS1wM1HVRoDyZi3Cih6AlAGa8fvCfkq5pda6MOmN+8tt0
jpKTWmS0YTqnX1saybemrGqyT7No5FFDqEVTYH/QFLhYBpywps9JvpfLGbLeNuoO
rsZLfYc+zXA/XkAuSUHtByuF5HwZtjx93VfHXMnNi3yBWobVCbudjUttLUN7LAm4
6l7WuOIbXHFK7fGDyrOCHzKB3d2IOH60VXEt5vEk1iZTYS6uQEFdH4efrOlEvtkQ
fDUiyK9h79ZA3PDNTodsL8UVKAT+ZsXXin/Ya6o0gl1sN7SuUFNGPmn7GlDF86TZ
I1Skpe9yBG/BBQ6fHd/oMuNTivy7frixwwZnSm0JxoCfxHzIoxIeHEzq1LQc+nVL
yfmGp5f3JjXdYnYcYBvGj79+JFSpt88kHKGUNu+c5ghSR33jCsWJq3+XensCg8/z
recvXCC1Q+PCmbantEp8DwMtsBUWc82IPZDiT9wjPy5EiN4KIxDkpO3NzUQAtBt2
uWq/MpEKUAZZAKmbI/iul4et5k8A3vEMKugcs+OfNCilpkqN/9nO/qEXlVFt/U8d
efD2t1+Ly5+UBiLiN3dmRfVd1vVTJxlFaP6eF075DUoi/YAolA39YqMrm+PI0h+h
MhHOmD19smFwBTqJwCYFbRcnktIOks//p0VMleZdAI57lHQ2ousgg1+YQDe5JQQu
UXCP+W2+N/VomSU/sJAHYcr2gLyEBMUT2MVbUwhSRtocCm31BinQU9f/xmojpv5U
atoTDcuJkMvG7uCR0m4IcFq4V0pFQDucJTpsQ6bSVsJnVYTxNqJcYOrSX0LCVlI4
cwxB14gXRQTkCWNOepmXE6Nqt9bdEzTEq60Qd5kOQBfTPLqaGZ7JpMykPIFyBh65
2aM7e8I16HgiSojjAafeCcGDK0Q9QNDdlnlslBmxyVU4ewSSLGQu0ts6IDKvm26+
pjYrt5yn0IXkCAWh9Ws+Pubj7cBRf8TzATgrIezvjLXd1F2o4S7yjaJ3dmwM98sG
Jh7GH0o9xxmlbljlCDLoNgybZJYo6G4PoNRQLNzn0NJS6V3ny6UKDe9wxNujRCMm
paEGOrw9leeG/i2jXRYAj3gI1GUNbsORyGI354bIbnvoR8iigLcYCiam2f7rftBT
0Sm/Ps0MbEF+OnrgF3FtOdOSbcfzmwO+AFq573WBDeggn1GH19x950zVW3QDUTmx
uRpvZUiOWKkfN0pA9Zoh0mYKSpmrs+o6JwNVt93rlXNxpLDDm/56J7yTTfkxtd5q
QClHctjVWHE5YDXcHhBRHT9rRV9lW++eOEEgbztpxIxcCuPEP39WQJsqgGZeKs2z
3quwp66nWzepRAIETEdvrayR0XMbSHR5JR/4oEGDXYnVOTA/RRMy8318I4A6KZZS
C/5TigHVdm65eo+vqeqFp3bn+J052Up2yKOM0glxXV+FRDAwsIUhKPMoDnKnktge
+QtP47R7vsymPV/onqEXHuA8kWJRPmUyn44Uy4inJ5ZVSEK06j4o/Hbk7njBZvjA
yTm2l82rOvIC9VOd6I4P1StB2wxRMSO9g43ij0huBDZwUu9SsspCAUmgY5yAPXcL
N/EXSciw0KcU+W6DEEWxXiBvA0vHhd7lNGa2dhOG7wMiRRT5TeV93luRC73gdVf/
LlxBqwZz1rpapwCvQTPcBHwwoJG6DpvPJkuZ2AkvX35D42I/ebsU0QlpNAEYQUSp
vWZyHMfzkjkP/6OYaip2Kqmn9763aS1Lfedg3YBvOHMSHZ97hsY/iOFLCfpt9Wgc
iFPNA7kNtrXU037dMzpfwbbyUmjTFVwXCinlYjRfQBPmKUIlVpvdpv8qvUHDu5za
OS4hINU3/tnC3Rvi3t6GycLZoMIgO2fr1o58dVoV//ieg3RCwJQTujZ0tg2hs/K7
S3GY2FqZJab6Hbo6sS6qbrJCiCkjujWtOupnRG8J5Vesi5rdOIQzlzEBhsraR1/x
UkAId6ryaivjq7wWf+jofiStcCCbmQLmjWgB9WzAzNSfY4nb5bVCPeqIh/0/G1rk
eGyP92ReYa1B4TTXK6k1QagjDOtopkhnRWjm2fxmv9vOmK0GdU3iqlUisYcAohkg
ZmLl/7TQSvgczTaBvVc0zsyYCuCHji+CkCUHKPdcMjM/DePZZsUyPsPvUPGpW6CU
dw20TXbeGDQBH9ex0xRRReL52BKQYC7NGpF6EFTCL0nUcJ0eyk0V7vgMdnz6GBNB
OxeHShb/A3fdFPmMbCR0tLg8Me/Xvz06i9o3f7+Gfpct/NBxHi7Ad1rnB6MR0jUt
FfCpxwiBjzVYZwPpURCWJ+pPd+xnSOi/TZUFHOHqUsIbBPoU29Hx6OWZ28kSO+uW
f7voksRZvNn3m9M+68vqVw2sLPNaxw+kI0n3RGTpkQ6MrCuplIeiBH/CsUR854Fl
mTsImv5LLeGvI4zfNHS9bgpCXRbmDoHUcXSrwOqYMyAA9NV34fLkGipCAQpn7zhd
KcdNm1zPsYEnB9e1FVBQmlVfzy6IstNCowZoO4NN8XcPMROj2rGBSGtzV5XsLFpu
u7Hyk96ok+M0MxnPT/CKFUmE7j4LFniTMB2NWGmvJODPoiqIaLr+X+W3Vx2QQfxv
gxGQzhGX5eR85Ug7A6xSVXdkPrk+XsPOH0w/xT7B5LLvvmbTo38/9iXdgVy5JdW8
NbMulCDf6580UC8y7jPosjCvHCzITWq84/S4LU7jiSSajmLaFx+eKPa8CBGvINBK
Bio88i+pXrNXglkm6eQFHmQto8EfyZ3mi2Vc3oQNH6V+wP0G22h6hSReDLqwoHth
0hLSq1p1eDYmBJK+SvoeF+vk29EqsInFO9kIXPVncKq87DCk/EGIbMoeFEfR60Lb
fR8eqkrEHUo1t206xk0aRRNjxoOe1/5R5ALciXGouLCA0+/YeX7AiFcTZfyP+va+
hQrYk4ORlYnboEJAJMN6Px4Lo5oeM6Pn4uZa28dKWdQGvPu5oK9Z5sRj/Hi5imlv
xqwyL7fNCvo2Plw4cwL4gX8eLItZ+VzYo90ghNSo/Q2NNlGpxJ0172V37QJWE518
sHbLvubHb/R99WEo8CSidnzyrSEWDTkFO5QpHDs1ICCXhDmjD8ybQBf9vzQFGB4g
Rh/KF8/JHFH74/7rjYpciiL6B22RfJulL3FLvZvnZsQZcBNkHWNImB09wZEyOvVQ
brb/2kK6LveqZG1j52zptZVYRKwJxHnR38JLybtn0RPrGx7tk/UghHr9VJbjmpqE
DjZfJiQ6/xMJweRQTOeMZVQBFEsGBnxWu53StAVuY3cPDh77aiLhUaaz5Vli5V74
3yCcBypQnA77+2bPOoERszC+RGemVdKltvo/pmpG6gmiP7Dw5MH5zUShClQ1lqU+
jlPTu/3IpffNeHopuD4Uj9uWlxSC1BXADmffXGFrEiUhMh5/twkZ68x80EP4IKMe
iOyoB2DRLWtdk/ab35KHeH/6Lwo2I2eu3ovhy8ClhcMEAUh4+/phgbyG5BxebW/7
Kq0Xz/n8rFxe/2AqGSQd7cvIxzFb4IUHDD8MA1FQ5Z5j4WssHbBTHMvIpGCOKKkg
5iBEYb3ZyDZYztOL3RKi0282kugJq80GX9lf+gzqiXQ9hNvJGblH0AgmaGWiECK+
c34P9XjyD/+E77864IIKfNbjd6Q4h9SJCbQ29yR2dk9JFJNonOFPtCnIrFDWh12c
rW6NWpBiE6hHbvnE5B74iiIQsKC2qyAb1Wn2cGJvQ8W9q1wziczZeD2kH6a0avDW
hDdUMft2LR7eBcEuLfjQ0Nk9SJMjrAoUqwpG4ojKSKLO2jY6IDk5sXQVtb2+QNBM
nlnQh2VLxBsTzNu66Xaz/Af7IyKjXk4nIPtpnMGU6QKvqtSjQXoEmPq9Ow6AjzMX
M6/gXxKQrQ337zqksn3u85i4fk9RfBvpU2axe+5ztxm28FgbOVUQiayalA6tv4DM
HoeE4AY+oN75zMhwCOUIbE/IHXFhTZaaHbuTJdSft+gxumQ8ZE/9bebMCsVMfa8y
lSSlhfMx29jiIg0GZ0m5+hs9Y7pKOzKa6O3DBAgm3+7hTcFdwlh1IXbCfVruKRfE
bzElM97ZnAK2tcnM1CU4FVgnpOOPzCZvqEMBBTDKKkA7Rl0j45NVFFR0UDb6/gdV
BRxhm6mih8ut52591omizaCjAjrM8WQxf2atY/kQPsQMRJgYNUdCHe4AfauCsXdW
orjPhHHZ2I2YVcUUj4Z5IOgD3gIDM1v3Gy2LWwZ+m5X4mJYIufVePDMd73NPwUDy
1hnej/+OipMreiv2/pj8wwbvIYm31WmrF4ppmLHfR5iNBYgOXAGeTynjE8SDw5sF
y3Zyj5+RZOZMzImpLHmVuA3cDe+s42cy0sToGoiypP3kfXW9Whx7cV+58ok1pwrS
ypUDbLaXaiJSDVr1iDw4rlAyYCH8mUFiLoCZ05Ze/wSPApqldR7t1cufA15Huv7T
9wIZo16ASq10OQpMqw9pBhlQn8MJw3MdXpftqKIPf98CNEHmxW6z06vf3in42h8v
SpEu5SuRNsm82V58qLJZ8VQTxKXcxrCtXnKRoEoRo2zq4LN4uq+yUIHj4qC4W6LH
7OE2b5e8gowm9Ms8V5G2yH6W5c34wx75vsyY0j0L9Jt44jiLfKZ4AHOrHMIlWfZY
nl3iEe56jK9mwD72enSFSfMlDr0ts0OkEL0U5y4VSicYpwwXCKqcXw3T0tX586n2
PvvnFlJBlGIwNQmjtZzzhfHeTTspKfLiPn5XkSIfEC2xvDz9H46xnPmNCrwEh+f4
79vXAviIr7aax24fGu+m/U1LrEXfCzhEcPpC4wwBIYFO9WOYy+NpLyzjkjR1LgoO
og836gzQYAAbfkyhWULGfHLm5lteYomfgL3M3EDjZt2CxEo0w2bHuJYINF13CdHH
vmO5lYpq2pbN0Y53ekO3bg==
`pragma protect end_protected
