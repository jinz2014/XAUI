// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:31 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dkdiVTFODJkTKMhCGAXRA/0pikGmKkstSG9qOVWbWEZmcEFDKZJSS71R/7QY7297
s9Lat03aH16i2agOaG4I48rGLq3X/DaxHi291+4RkDc8RXm4ZUfNoHISKJJQVZDt
6qP+JJ91Jv6/AXvTNOOASJXNsbgAoCNaapQjsAk39yQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9632)
K9KlnM+ACIkfKDZnxtwodCycRDCtC4ZhCroKGMitNNM5v11qaG2Ix1FVmUyNYYOq
Lr9H/UmbM9sSvwL2k9c6x/KFshlGa97Xdwqj7aZuoU2fhuwYb0pNuGgfyMEnEvn9
XRRS1q7SDoJzCWu5ydXW+0JquYybi1xvouQLazDIAoCXirZ9vPywMJBcHi3lUuUZ
FZLwZxNdhbgQ3XVnIzEfgFBamtGaRuevCdrSd3oPFGMIG7sH4O9Wb6mcbc/1kD6S
On89WmLpfGtBGM2tFUTqJ3rMo1r1jzOlFtJvXDvDanfyj4aKGYvzenFMJBFm3fAm
gC3HjJEuJuwgOA2JjUIgkCPgDqJseni+V99rlNMSFjuNC+LxKXWY5iJ4tq9H/fn7
tj5JuHgiIhqccK02Zt60eCZsD64qUSMmLzX633bjBhNEq5jAYBk/Ujqeym9wCHg6
sb20koyvhqla5Qb18S6MoQ2/Uwzan9vJIbL++C+VytKy6FL5mCLoYWiuGzOVaxuy
G2hUvOlnlq3neHnPq5NGfZ0ew294Hnfcjw/Ah9dIAaL8oBpvleXdkQ3SuIW88SuG
02f/0eilWXNTJokV9BwNIQi0mRhD97iPLqWVNNE/H18bFuncyU4bgcKAwaRBbh+k
/H6BiiITYd/ieP7NUNe533Gzo5Vvytyz0cJ3Hb4dZ/skgVMWMxRy5482/uH6XarE
7gvq2VWAryOwaz4L2BrTkXuwAbkBBupToEH+XL8im1+WZ2cJ0w9wYyZJ9mmzNWce
N/iz+y67Wg2Uwfhb1jnmgHOeSC4up37Ho//eFjE7YUvif9HUJ08bveY8CWaI8xwy
ByW2Cjz7RrUEAGo2eeUkVuVGAFpY76mYtVRjfiUEyTDg7IrbQFk2zQD4NqfIwGyV
ehHF7AJ7slrt8laR/1oc6VMO4giiPZUGFGZ7H1gFbsvAGgK5d1920v5nLRp+rY34
Qviwgtv0JCOrMzKkvGWzAuN/WCfFH5/Zqj0PwXO5gjLMkDKTYuZoaKq2TbseFmmC
FkBo6xwx9CUt8zXZecXqKVJRQxjUhFWRAkGg4zaQQhEoJjRLKw35tOINIDHEWHe0
vWscGnRKze1a0lIRGdDZ6VuLRRFQq0fbgkv3phSP490xPaIWlifzaeT8h2BdPJfc
1WIugyb3zYA4zpZys/yDaFo07AlvQEMmpA7g9gQ0zMUeSo9nfmKqFG3EXcNZr6bX
iOVDoXWkQNOAcYAiYs5icUlCHrW5KjbLcYKYDC2t2J870nbY5A4bPpTp9ZufPI+o
BVFHYlERRoKu3wP3FAAzgeLjIJy5SedZV8Luf5gPrYTqxzf+wdFwUE+GOdReZA8H
uK4UjlYUxIZ1cKI4FWdIAT4f7l9oHOimeeor1CR+Etm4nSCY9FXYmy8InJmfdnvk
jQiK11KjdEOXQwrJ+mp76hxSH+YR2GGVNASGnPDr/00A+C9LhlpIqZ0w1KcmdprA
9OWFxHYkrIeETZGxbcdQymI/X3pd15bOzx1VZLpfzbvc2KZNHJG43T/lqlFejO42
vgRimdDg29cbW7ro951K1s8betfg3ST/7BCEQ5qlx1Jhz1qXVfZz/v5v9UgZ7e3U
WydKNAKym1LR048+1PrEugzPOPhAtSTUuENqOV8dYmeJNIwdFgJ6hEDLGCiUrDRd
bv+Z7vRTbov+EBx75lLfd+DaBGHIeQ3qVsdEkwFevYD5dcodoXyQkPsB5Ug+igKP
4longNQk6Y1ldeko/x0LcyNEDRrIvYzAgzMIEn9ZSd4XnNRLTYXqmbvwONwJBH2y
cTGG9fzEGJNUqLGHuaIK4LrWPYerl0hT0ZI37MxATeZi1FgstlrbdPXuI56EvE3A
HRn/xhun9m8c6Ym42YNLGvWraJg1T1tNib/kXKzICdh1Qdt53Kehyrb94Wd8cBtS
HeV6mgyjBL8500DnfEGZMb3ioSXFu8LbOpXmZuH9w4dbnbfNlIwesubVXloKFKBt
6l5hKfGGZbc2qdTFQaOsgJkL03REFqP2M5foDuywP1Ez1J9wDakpREe962YVRBXT
jKr20lFcpekVi5emEmsnsvAzZiMvK9QbVMpPZcfEdZbYtvjMGyyA8/MpKddsIkCE
mry842lEnP1jOcCskS4b5oOsGyqIJuR+gRJ9O70Cllgn36fbjBFdC8QyXax34zbM
dexfBBB3Dnnu47Sy+ajeCSgxzA0d0si03oTHsgXPZCEzSwAXypD2IMR3JiXzLa77
6jqFMkTQhW1kVtdmxnWkj6GfnuxeXLUtzmaxX5kjmx7MSHWS/teS9OxdYV0+bzRk
cypZdayEGB0eTA3+GcrG09WekSFqZGlhVz9EpLQ3ame8BBMccswuGt822XamMYPR
KI2kKKyK3yYsPTCkZYRC/tgm8mbY2Ruh1CLLZ7hmXBvwKOnUr5CPb9Wr1UtCipmu
V90kUxjq2n7tWlPtrK4H3X2EVu9L4148Ti0Wyy+xabYQL8Cpg3VnZlwSNEQC37KX
wLzCOEjt0sMkTV7nfe6OpugIHG1lGJLraRGaWq/B/LpG9f/Lpf0NGR6mAASdZu1H
JY8UZU4mO4RRYXOdBk8ToZvRAGR6CEb2eo5yJeIAIdCEehOROS0L0IgZlu4h+jHs
kq5jBLOTxMbDaAUE/bw6BRs/1+jsago0ROmucpVijOO5YeKElCVymkFg8vH4PhHf
CTBDp+vL0P5hfsLHc9jMDFpwy488cFxD86aEyU9reZxSPgLiVH2VIuPtTSx9rm1J
aP3WtoAU1wLtoWpL9DBhn1yANfqTbwwxEX0MfgAqJXkXHfJDovuTcez6HfdP/jq7
dKgFZBWakiHC3l2fnxAQexFVg4vAvEb/F0n/8jGwZi4Oi9JZAQieHLEcS200wE3p
5TaE6RZ3M4WUHFPhNrt0vldhU9y0Nb5OGDmNEU6ZgIvjXVdFaQnuoz+kZy9O7CGH
zJ5OavyBgxBpZ3gg5Q4JfLaaZO6/d38IzBlWilqXkbGUGEKaMi6ZPBhqi6/GSLaj
Yz/pqjnQIIDRz8ZK3Sq1iNkQvFISRe0D9W9H8GhyccSsXlWYYKG/oBTJhTiGzfqu
qukwEViKef17aNG/ANB4mNnGN7VvrJUQYk/CgjUe+RUjQhMpVBbeOF6fLaZzLRAm
w8KbZMBss6XUBy26dRs2QS6OkaDU7y/v2P1PJO0N+pHkfU8RvNiH1SopcYvhGZo6
eqPfnSsYDHvNfBtdSXcqlBDN+OaWIMKLG3iw/67TZPdQBX59g8E67NhoPoq0T7/G
owF6L9BZ9/2jl3a0M44GcFbGhZ6IHBfno6WdbzFI3/y/RmaTeNECbjnh5sh+TcFo
8aFqkaaKocf9xB8hTF47IxfJwqenF6IzDzO9xJVf4tsLUhVixRkXVKxTH776Ud8n
sxcbF5L6NxBlc68wCl9GtdlxyIShovoZCShFzcE36mmd/vDLMtMFY0m75I0UDSc1
w/lYSCvXiXJftzUyCCzsQIWGZiIda9cscgOsIwZlGj26943N4Roc3Z87gchwjzu+
8+UhFIuDa/xFmFQZeopmLLw5hfavcXfmH+7qnHkfp2lvk+tYhpRdBRWwaLDN/vea
bTS1Gm+7DBeZCLddK3veSDBXjJ6RVv+/u1Yq7HPc7hw3raf+2WkkQKqSD5kfbHSG
XBNBoagit4igF05mbpth7ZQEdb/sdBnp+zibVx7oBnmntPp2urv6a+HyxnLhA4Rn
CyBCTrl5za1ylGBhnyDj3Z+Pnt++xHmfAFXsSNadtjtYbSztV10E27kgsUDjyY1K
+XnOx+AfHKvnqtUreWoC9TC8Zc4DP3fpM0/0TGd6oQfTvbMJGmbpsN1GmpXAFvxG
Y8wpB+mvjffH5vMJTnbwC00bNdKX7bhPQzHUYgOmpffhTAXG20c71f0GE96oCpIL
XVLM5RajtKKD2KfMssXFziBiLjAFRABu3HbMD66VAnOM/zn/exqzHKX01xPeos9y
dTbVtbS1N0abFWROx3y0S7qHAJ+ggwzgsBcNfiqBFklMQh9+mnvilGKhd4PUOpdm
yhEUnlxpwy0qu/9+zPTCDfhbNum3DiKAkS9i96u14uJDFoRRmA8Tj00ZgBPlnBNq
UxgmOxm3G2txA3xk7pbV2KSN/7xWsNETK3jcrY8H6+IOu1nD7x77OcfAnvn+1f03
QuPDdvEK98mTHQDMfuOyPx/lorcy3FIinnzZ8OsTnuDac/J0uJEZ7sQifzvY7UDw
H3L6JpgT26PO7MSKGwNs1uWd8wXCr1Qzk1Iy3ysS0/6BHJhqUy9nsUfbx3TejRn0
0eT6zYpiX2Hbjhv1n2DtKyN6XUI3J+e2gIqI3DY1hjnRd/KDKZEJXmxp4jYDNWEm
2kO6oG+lBhBh7G9ivGVMzWAmYsoBYqoywC7JesEQAYKRbZatNYS2NsEJ4PCAgQ5n
LwXmYMLueCppnGlyT9RboXAmMeSocAjvGQoo+IbuapSU4JJdTX7OKpWU6d1l5wLi
/mgm4TByuWYF7r176Jhe+4uYhzacKgDJ93eS7UgptELo4BzSAx4vDAqiBMOR6hT7
qJrdwFn6c4fznJCkybUGPUCK8ce60L684gJvGMx94eZtJiZQiE1tsPhHkV9bz5Gl
ZFZ+GJfpHMUHYhW8sVMAM0uxeDaZvKq6krzJJ6HXdd/d+9kdZ9RWlv7+jhltQMgS
8WYCTXENFhBVo+fdM7SZ/lbO2/vuBy8xPTutq7GJyVzUpDt2EkKPeQzaFk5pA1qd
DpMcRLCNC2shYLDKxj7WiTZbQj32owcc8xd69cGdWHB+qzvhPuYmVbHzRqTpo6lb
sm3VImUmtputMyPS3um+p1w4La3/6BHs1ZJOiv6fpwCZsI8lE/+Oxt670KZfLk0f
ZfPQAGu5/2IWy69iky+/xsKvKBWgVobjvXJQ45Muow1RoCOfpq5U7BcQSVPW6DXh
zzUgsNn2kV+o6X4N7nyOwb3Cir7dC9QA7uyRvtCb5TEbSU4cNmBmdPCnUziu87Ha
ffUqoyLLWFoyogWCISt539U5XCML0QXfCei8A5yyfp3+kcNeLQKnDwW5qEZyd3iK
0fH0YFdo+PTBJBVDWjBZkUrgIq/GsQzzDa4OemYHmfjlQATkX3lhqHT/U4kNFqqt
YDRdBZorif/QfP5XigSHFIpJOyXrYeIkdmVlkMoJBrz2N/D/IxJ4/klDeBef5kUQ
BIGDnHnwKyaMmEFaAWVdhK1sTpJnXICAB8OJxnNhZR4KtA67Rtv3m0oRsJTIv/wH
D50NudSDRE72iFKIk2nwKbrhbba/z9YoFUWENZqbNRjmljVcFBciRAi4On+4f5kV
MuYSKmk9Q2WL1YUwiZp51EtZHjO8ojzbh9eyC2Bu+vgQNrFZDLk4qUoVCL9I8C09
oueZsdTOQN1PeAw4jfevUKiti5EH7JNnjEDeyBKJlbcwLjqE85vyEXeGnpTKw2jK
P+GjV1DiU2/27h9d6/WYJstLiBAAdGgOz6BUr76cY0ejUuXLnr0W+RhW8xorGo81
Lr4UpJhvKCunN07O5mYlWEcykkNI6g9JPOgqjw7/bUfosiER218FI2r0f7xutEJ4
3olukBrn86vDgebZQWnizKhL51TzT+iRU22qjhgXd02hAuKZ/sAd0Qiu5Y3mHohN
hkvzd8I4Mjy16N27Dcun1AJOA6G4oW7enR1aaSi7rJc9rDfpyhmY72lY7Q7fgac3
LEZ87iVgfwVmi2o49QMW1jUX8r5ClDYZNqgBccHRd1WKHdXazqN2VLX+Po1Pf9Ss
N4b/k54eWojKWEit07BpojOg+YxSNq3Sj0KUxdsKrXBdh7IeL+imZTWMrVsG1iaL
CnckMpCW62fnw8ax6i7ny17R/2Y2k/vvM4fEHIgGa0ZAW2zN0hyY9ym/Stk5v/y7
4ZFbcQx4xWv2DyIzM4eRCEVuJOlNjW7aN+S3JvfEVYo56DmL5sHpRAxngpJZVNR6
bvcF3gnLriAFiWweXuueBoEAGGIW9EWr3vY3RSbE3nhI6k5CAnpuqBImGEUlcDrN
BSrNmcU1DO/6zlCtldUVkE48AfWsVOH49E6kOVxL8tAYydrfIIos26XbPFkZPV66
4LaKl2uJtjZ6Gulq3SBUSTMW705+WsgWlMMSdn8zO7kuHunrckkcmwUL9Bo2inin
pQPtEH1/e4g7ggZ4J1i9zxYTm9c9h4oCC6VVK7oMvEwUMP7XJORbsibaWdwY3Rh4
y1Ra0WVOy5tZ0g2RVgMNCQEKZST4TvNpvIGhpBO4DAqSy2eF90GU+ucmKzNOWMbA
SOvIW4QTtMyY0jHmz7Tjyn7ACWH9PBLFfqLRN0cFygGxrORhYf91xXnzijjd0vjw
sfvfHSPnkYtQGu0P+5H8cWTlmHKHuc4f27j4KQUbZYYWGauofs1ciE64mZyZ3Agp
ftuT8BxwK1h+dYojZUelusRdEMQ786xEt1Usza2VsWdSVj3o/P/k2MOGcjdtWAKt
ATTqfyxkRwyo6XF9v/fSl/Yypv5Sej/K+9NPvOy4uSUaVEmi2cKdRx4M/DWYpZnX
ZgASew3LbSNCvIxMrw8n+TYJPyRN7ZHLwhXwZLG5VkzF+YgDnZKYt1Dp+PHKaFkf
RsuaSLVZ/MVVuwTgcY6nQ4eKqWll4nugVPlohXK0jZTiAWG3rN7zhCG4kxayfZUu
DjVM+6yywPXSx6trdO2YXYwkV53ZPsTHWZZsRI70kHOoIXjoubH390xWGra/88VZ
TrgKDkQ8mFT1/XgJIyQPeBjZPsdnpWcz3yo0QeX7h3QVb9bYB54+bMujbh6el67B
uP0no579cIy+A1HiC1CXsmGvRvOJupT+uphrHUZPQiB5WlWG3Dlv3x6BTzCA2YYI
YjtpBeNZcuWupiHu9tGrbQqaCb12Adw7JAs2RgwA+HKLei34FlLMg1XZUlgey5rR
5gQjdPAEqC5ccaRqLNKe+8mUoJj/hSHbnSB9GJmlWU7OK7fI1+RgIViGu9Hj1AkD
1jWH7tSS7YaddCQKgN0Ecc7dRfxJKgbqWbGNFRo17170Y5ucMS5/w7Y/wSEh6kcU
Vbpj1wMuce6/azZs88jIwC6R62Aj0QaUvFG/fkMVGa7bhEt0YnhXOd9jQZxo/hs0
N7Nfql28Dbcc5ecbyS7+225culzPSQhCZL/gh4U88dk8nhtA3c8DIUQiO18gyQeN
YC/tpbu8ym/QJxUI5WUkcPqy/9kb+G18QOPRZtuPo7+4766wg1rFmU8ZpSQyISap
X8DFPzCCplnI6VJ611UyXunsmLKsfy2IgwKKP+DhLLEewlJ58wmJnzSTzJtUhdDO
pU/dcn5Y/wV73OHCv08Ua5sBlL0J5H1l/4dcYosxUpexsWNE2/my8jqVl5Pihkln
qWTYel5WcNyLZiEekLvFBT9kvlpranvRTe/DXZR0NctwNS+vy6lia50upcwPFR8s
n084GVRTV4+/d+xssBY8ByhFwwzaBoxnBRJi8lSGEUPRHQauQd1E4wmNFji+bXj9
q/nHPEHveDYOcTwA+BH4WCdI3/fEeFbbtyL0tVXPmlkkDhEMthMQBZI5oM/HJMgK
DEEgi8h2KaU1ndyRfEbnnhEqUZM6Mg78mYTUmC0xTrEW2loqOdCFFjj58J6lCXvK
wLgAu1SJgtuzSdEhU5m/4Qvk7tn23S5leyw0LE0UdDHpISUas0rQOWLSrNRScgap
xkIHrNk2OoR5cltwTMMPdx+JNYEhYfRoD0ADa5m3p7/bbNY+iE4ShEZyMyNqDeBK
nKi3tm/ZvAZf2P8kwAbD8fn22LKDtS1Da+deUFVgu3/PLRV0WNycNYnGLLC+TqYq
0xLKbweZ/feYuiRoizytXJx41rUOoqW5f1oM9UV49RS7ONZRlTHcgnHYG1QotbO6
NjlPD4wELGS/eozhAfG51b2WfgTFrw9w+hE7xo3eqAmTdCXfP/rpGCoD3xYfm96t
bL2h5mpV+T/M20ty9g476g8geGA8dVYvFihn56PATy4GK0oPZ9U6GFZU37A51qRq
szF+1vIbrrJwrhKpm9gcfPB9cGunj6ghwWFcrUom6JT4zhyo55QfadpKMI45h28r
xNDbkEszIqynPiZLMKEEMZG2uj+B1RR73aKlLUBDDNGvSfgvJUSrc6qOhcWuH3ev
oj0SOtUK0UQRvttjfod98/paXRdaGInJ784M/kbUoW3Z2WKW8xVlMVmnq7vVRNd1
I3P5LqVX3n3a4EsZAG9nokk4sbMQJkDZq6cxn+HG/IkK9YR1QAaCOztB+0lTe84M
ECnd7NpWN63cEeWaqCK1CrJb/2X3yNdq0qSYh/DGzjTEZ51++Bhj9qS8YcYhJ/J2
8fKPxrz0O2jFB1g1mNWb/IlbBEYyPvMDOrY2R44TE8pAZno85JMdC6JNakQbCETq
DSMEciDC6yg9GjswMR87BOvsB3ugksZG+DNOtI8U9LdNWd5k1J6OPu72uCFVGicd
D+WSL+lPT5A8ibZDzszYJMFErFBwgEAZyuPEmh5IZZOTmEyz4duWjpnCDtB2lzPD
YQEGv7yIrPu/87oTwjDyYq5OxS3H461zqUSDnFO5qhXtKpRwK9jUEVTxv8y7Qt47
1nIy5qXzQdlwSd6gQfMicOplYsdaeHiVtJDO+BXMa7S0zJAuUfxmQI9To3VztqTF
PSLVv5aGmYrnFksOy+WnK5gGMf438c/l9x17zSJfrLLm4VaADb47dzZjo0WMF2OE
HGMILogUbKByF/mkV/uwaTp6MDgC3SP2OxZsmgO4sq4HzXKaDUTJ3spJSuRwRKsR
aZgyq6U+EOv9qfSWEWdsO0iBvFkRT1O2n9+gHjUWsD0OaWC7kJwY4KDmiDxvCVls
fy4xQxppOhsY/tLgIYrEk2W63D9BKN1nO2DCbHU0yy5CanRxtdeqg6S6MKB6F7Kj
sSqdcmZlbI70G335w6ZsPCANpOuxBUzlLtb99iBqW9jvZfQfFg434kb9RFWEtTHB
hDWqOZQrdDnnqj86RiNm1BGTZmNKi1ufbXEicjhZ1OPkdTmbQzTixqAyQ+5+SDdW
zhx4JL8bKz0v0AR6XzCRU+NliAw5S995PB/dmNlOaE6zKCpcSxgfBX8n7ypRPIzY
Oa+Gn1MoA+Ozun02X9l9ayoi6tkEc912P15A39NP+Wwd125tTdmaYhYvLA23RHHe
UE/DM4nxC8uc9pYmf1V4Qiy90MuGfzAlJf6iLThTbQ+arqbc0cJbt06pLmLssUoG
X6DP0tf/ilGuQZsQ7Q45Ep4kOUTZvBoR2OD8fcXo/agDA1tNOX3AsZGdQ1JBPk1U
NrpbGvSCLoysTQ2Fpv351torH7uP7SSYpIoCngrGXgW/cuBrRAJBTMF/bkIhSp5q
IKEc1FNo2k1+2l6zGm7gYzpcu2cjPZ350V3wOipqFWAkiMoRUHZ6T+dRhKTTPLf0
N3vCCe3qKZBBclYieLgQxCzoXj/nOij9o47K1tGStFXaMsUqfO7avE1WG5frCNSx
dAvhRe4Tn0o2qYsSfoyZKMH0nbvnVd6dUuVo7C9DIhqRrHldp5nY7rd/LsQhA3K1
/rP71IvXojWZbSywYHV/1q3kGTHByNvcPx7EDQtv9gIKrhCiPV7r5RYR0c3Xdn8N
nwyhx7fZF+sHxUkbY5odRhy/xHLCLSknbKvy5aVqdZXABCatNXZfrLjUc9+x8GTP
VbWNxggAsvlxIyMNpm/I+H6ClJKyWCT8KAw1KKFT9dM0Fv2eHCB7BI5uNetNH7nH
I3Ig9emCWoDl3BJXoyLLayiWSPDxDphDVUyq23RaADXmRrN350A9otHqBzUITzaE
QerUkRnSk4Ealw85PKskzNxbIjjSSwGJO1k4PcWyP/GfDvx/Uz8O786ysjU2dZ32
bshjeWStN82Zym3P8s0RLRx8LD23Hcfgv4XL3O1iO/ZwyZUchLHwvUqf5WJ87AtS
/W4bv1IET80NeJyjY4ZFp7KKXSDMNJDDuPkCnLx0ymh6XXUmxxwBLSybUGcajyeL
/tl3wYTA6gO5HIAK1XadIN3fQxp5GgvxtSolsK0IVPdDDISHD5MMlVUfheCDvBEE
h3qA1vckBhZCsXLO4+JhykvysGIMhB9XsjtiMRNXSqi3d9o9yRpLCWPpRuA8Gy1+
64Gp9v3jdy0TcBjqcbHq2e9zQghNzVOgktMPwUrMqmQ/XF4pKN3Fnw4R3ystfV0/
ogqMa0i4gedIX6+yjZ+RDnJlxR2kSEmJr6OZ4zHFn5pBz9L4yMpuRu8U0yZakUwD
lExO8+G2HVZuDBqyYFoLHJFZeJYFj7fbhf/El59KJ2fHOTYRlRi/MI3k3pKSSmTs
gdt+Fq+iOIhH+6opLpix6CpCHrTxKPXuR3FK5BKBu55bjqWPRmjggqnhx795F1bx
Bl9z2XlGJFijfUCwYQ0Dwse1ZPw8hpgVSc576edLE2wj98dOGIicAkv0F1Vcw8or
eVew+Q5WLDK63VUohTSQ+WO8CcqiHsuDPpGy4TH98pFaIstDBcoG+bI6yR0GaNFZ
qdlPR7faP2xPrqsSghvEIRe7j6lRlBP8ghyuBpiT2ujgKHti1scfGhv6CkrZHjwW
JMQ/Fe+7tNj7P+npkHsd2RNFI2nz/pIKX4q2qfmRXHj7jeArrOhInXK2P3sinHM0
rr2vz7kCJPmVlieHDs3oRN6341j5JbUBRC1bdeumAg3aHUP8e4gAjk7ykXSn/Fap
fEFQ2ktitP6QnCv9JC8gtWzo28pUlhx9ramnfYoCvHHmEMrhaeBWA/eJE6Ak/wXt
xMFAgB6MuDwNn8kt2btIQpJwMs5xlLoyFfcJoXigRyrq3BFaRTMLB7ijLTRlvSsh
ILnw/1r6+r/2LKmVhgl2iDa55NqQ1qwAt6lXl+ToTIQ6MUfW++aEgkZiLQ2FSfvg
fWPl5IWNFLXQ2Gqyf5Md2O4X/D7Ij7LejDhK4yInkNrq2cD3FP91zkUJuV/pWmU2
qaZGEJ3CyGr+NsbwR/t5ocRuiNzPugezLIB7ejrUGpSomiww7E3MMX/Y4sWiR+nL
uiKDQ/Bg8kTuY5S/Zgs1NxWXtsytnBSyWXqLsOCY2GcUrCEr7WuqUNcIBd3LHjRS
ODAlGO+4CrdcMzcDZvxmuaQIxRviO6lZ8aXQFowk1J/RnbWvYSezYOEabAgf0u+T
N69AFOE7Qn4b2+kekOyk9K5ljFJhkQtePOB5jOtchBtc1vBqV2lULW181lC/653u
wFvWwrjjryEcL7lfcYEJIE+JDIG0RAPhLE6r1YhHInAP4vWcQ8F3qpfrVEYP9RoF
d6p0jdYdYQQigbDSSkkcAxoOWbKxDjrHkU+5I5ADMIPTHkkhDgrQieEsx6+HHLUF
lX9wzyS7EL6TWh3fMxt2HhgfEEbltF/gYOaOXeWG/jqUSKrkEKTvKMepcj0qD5Qt
wQjhuvuJ9+EOJ3+U1COCXNcrdQ10WVevjjEiz6AzVBwrXAicXoZBRBWcmu+JOCCv
SxFCaknuSvSX47mgqKbpi6QjyhlO8rQIu4mleH9s4CgXH7MSWNT9xkvk9D2sjtIa
fOR5E4Nmx9Mx6LGZlk7TohcECXv8LbTFRDBtgPfg2fq6xGvTe9LqRcaHPT9/9VTU
RGl2l/7Eu4H1aGZX2xy4KIpQ17PfLtKiHlsdjX2fAJS7rSN5F+sP1do2C9fdXfn+
El3f0NN3m2yOe8nUuzpz6QmoavD7pRZUV2ZS9fQxXxbsG1zzkdcHQeDi9wDh4Ekl
T8hOFRG9bGl1NIvih8MKXBY9YjvBQWMjX6tyNlDeybGy6gYsYbdEgi46wwhRPxZ6
KF5Kb/6605NJCQGPMCiiOm9Ah5VHVaDWZKocMKfHbzw7/e21xo3ezSZzlfObY8ex
DzqR0+p16tMoWmNDmbvdKpeO006ES8EjdQ+idNLdxklxgeE66Q7XOpFM7PLQS741
XJIuA+a4b/bh3WEb7EOMJ9/2cuLsq0JyTZyIn9yaVhKtv/gnRYXN4PbdVliey22b
a4g+W1lBiToDJAsOMR2tUWMcO9aCm8RF1DTFgLqYo+rpwnY5BccjXDVyYpuMd5hP
GPs8iO1pDjq3IHK4oH2FQPN6DG6VEF5rjD2zRU8gKHWlh2QHiIdMpqL6ar6O65fq
vs3kQOUKyrobHij35L0NE5t+3fJECJKFiGHGcit8RpMqL4dGrIqKhjT1xaTtHch0
HoZYbc/jpDFvfiin/CqkXSkwfCennoluBTfvkYUo+zz9f3rmFxYGPfaRk2DUpCrM
8CkOaW/hbIe9YEDQt3fjnGp9Z317+V7CsVyxXftOn0rRVnQrJoTQ/CVYMkedX+D+
Eoy0Kint/vWCVNXVEub5wszPMyWEkyY8Oa0k8dZHp9IkFhC4lSpaF254N2XhuRJp
DKsDfB3hlQMI7vALzIX6Qa1ZlEloJGfhav5gy6CtCI8D2BfVZHtpp83vCgeqmGUe
9n29gLhId0vNyECMf2O8/i+s2zHU36sbl0S7ZdNftPUCpXUJeZRlAoDmRmk6u3Nk
GE86cs0DjQvwMwHHFaX29a6K/JyPDM48XFIPmVTJc8sbX8YJzqnnPVg0Xsaw86mX
8bSdgevOmVWEyZeFR5Pte+XaHDct0FIsk5HRq+k4l6+x7HULC4mxKTXEIhPaundX
XzX2OEcEeTBc4+Ccw+C3WoYcewJhUYVfb6V90ZZANvMhsDsVnRcBRVM2OY6ZZCGq
EIKfBaG51FBfWZshR6ZjoxLL3eY2wLRCAVGdHsLlYFYN78IWmoKVQPaZCgFe3/jh
s72mxulhKQJTWfQOkQHymjifHhZ8tOghBt95xKmQPZsUlkd2xSUnWH+U5DEp9gIt
uG4wgl541g3Wpkm789oyJYmG/7I/5E1GGjO3uD96MUs=
`pragma protect end_protected
