// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GiuXa9H3LexRCWQCH+aROwA3Gkaj3WIzlKngNmMW09ajMgVssr7zP7ZqSl8kp4Lm
ka8nK0NPPAVp/mnShqF5wXWEoVfoB0IKq3sGCDJHb2AZbBOS211w1o0xxvWIbJSS
7Adu5q4DiFR2q68SNOMsI0BlrzGtZUuEGtW184Xe+Fg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5424)
NuR1+K2iVsVAuD9ExqsgUGAZVaeY+1pt5kEvRezLyuRt+oyUYJ0SkzOf/MnBWF8z
Esh3sUFfz/k15RbNPSKGm+q60mR2R8nYrDSYFyd4bGHrdW9G4sisHw/wtFelAYRz
/S35qU6VfIv6R0Ndh194Eevh5LRHhs2eEY9Fc54V8Mu4FvWVyKK+G8ENwd17sBeS
9xY6HWwkdtTmgXgocVDentW1UAKU8bhRHpldUgei9XmfvDM4kISZhlAW4+MMr+Id
SowF0z83oUa0qI3Axs0HgqlKXtAVF+N483DEM0MNWpRCUxdg03mHYKxbAWBiBMTc
OkBMcqCFRpH16/zF6QivWe5lc2ubcFCocqmRN7uhHsoLID29tada9tmNsASdCg3D
d6yVo2wJQeIjyAxxZa7AHJxnw+WMX6hB6fSW5WpZOyHwRVJQFEWPIGoNfWVn/0Vs
HE4dA5i2GgBV0JNmjUnpZeq55uLRN3b7ZnAwdL+GdyUiritALNS2IHcGCf2/+gHN
w+cCBRuMAXII68yUGg6T9WtibtoPKDz8cwOb7touvt+sJyur5+kRAXZA5EghTA1N
rWSeHVeBBSRXU/RNdmD9D+wdh/eNpnizUMU15hg0yLi61+S4b8BbdVXzdamQKGan
GrLyrmESCo4774yfi2sjTIOy8rOpkREmmDtDyyQJdh6Lz4NKv6Dj0UdShhvCX6tU
o8gfWt4ekyMGGudmwdRviJyFXOwS8EtbwwXdILH8HDcgz7PJJahLA05A0hLyaAQk
Jdv8Cv+HzIPS0+4ITWkb7VAeHYbIhADzDwcZ2Osf70DSrYxLMxDJv55pP2neHGj4
R/M+ZWBxQyos2LZsp4cUm3NPkJLHJocu1PPDPOCf7dCMqSyMLQOouBEj3ug+pBG6
x+S3nUO5tXTmrlE6MAtx1j0nofw6Qwrs1vjqEpx6UnZ+JeaGmXW4w7WAOIzLDzuF
gCI3wrsqlhSYCDiD2gbcyJSgT6Zm3SDz7F6W5my4RJQ0tQ/6la1qYgv9p1X/gR1Y
QTcou4wEeW6C2FpApfGXz4XLBiFPVfWdwoAJ3rxUQ0XlLclR3hTX4uk0tElYbTsU
n+FQBlGWPaPaG8ZF7FTOcxnGwD5KjRdg02JfTpDKehKnOqvWg7G7bPHVlEyG9zq9
RVIScSQE43K9c/bg9YrKqMEwM+1PEZ9xPVQ9wc7wAuEhr4S8yueHvqupmjaRZGzm
gySIm7HVFwBvb2COPRLmR0ONy4jVXtOze6UGauG+07MiZjomyaEQDfrX94BkeUNE
5ear7wVla4yYXG1mJlGQk4/3+NmC6LuQJGWKvFtzPjTduJ05QeZ41nj3RgXQ+569
rAc6PzR7xc6JHX3KOuEcbVT4d3SvlvPhJj533wXr4SQfputQlZ6brHF4ueXmG6tn
FcSseEeY/lgCpJRmz/b4aCO5WL5KnJlBWiBYIz/AEdfHlr39LMTAZF4OYD7mXglP
pVv0EE8NstI0nSu4ffsI+dtru3hKBFR90k4FOQKHwcNXcjzUzgn8z78qARRnIXBu
xedwj9ZOciC0qmDoTQ3IE3VtxGSwMOg+XCCgLA5ZqvG412BfBbqnoLTPaJIVeGRn
fwOfvvoWgn+y/BhCJo3+JCV4HUv691PEDpL9llUf0uy/bCwm/v8BY/iHyCYRk6ax
Vs+CVpKATpB3DrOH/ULPFcBv311Z1aWUaKEk+BLk+deRHdn0wUO8ctbhzfEzagLm
IFNhkghR/QeUvL39kCrWZsaThkE6/WPcrvpNzloTS7P3MuoYpS1P4bULmLXMX5xl
wiyw0xS7uvNIXusjb2G+9GyKAiBhCTCKEjl9w1Lw4lFmnxwnb8awA8Sj4ZPZA5kq
pplj9/QiFSnfsh7utw/x6QkkYMdENBi3IQ2av+EEr4+bySXrbPsn76lF4oKuikMZ
DwVhpobvhiyNSGuedBPQ/nYBumFmoN70ednOcmxzicbC3uYo6x2I2vFniQ81xFEC
33+7FUmhW6Bucvz0Rs7NgnUiu0ToeOewkjEvI32KNE4GY8tOtNwoz/DGRls2Sqp3
1lq1njfd8efy9Y/mo6gN3z420MUPgeBSo/pRECxRFHxbYuZpDYy62TuMhVY8ZNSr
x2jau9C6WhvwgzNkC8Zcr1yDH94hAwXoiWqMe/+FTprevHlqwHiPchu21paeJQiY
bAi1USS2tqiAqsHdCSEuu18LDxs7zrKlnwleFkJfWV8lySMijvdC7PTorQQ5Dzk6
/aJ9vC+Rrup+cJJPt9KXpEtByOEEyjIbPnN61IaTJlZuisHqqtYqiC20sEUwbzxF
rYjQ+McTe9mNVohR55OQEXHRIVq3duSZIg8Ievc6H7UWYAO5OScFisxW4zcfbDiH
p0zUtlhAb1LhIPc+fOWN+p/0lmudWdm5v64OmsKv23cDcUs/0gz8piPJ5swbhyqO
VD3OOGNE/crjDTHcYQvfzt6BXK3nCaaYOAPOV/Tg75qXH7PATYWbwJfQ3GahDACO
Dukn0HOFzQgbLFPgCNT/KRRqTFusVwchbrk+UWbW1E/vvkowi5KeZ1h5Abs48YYO
V1fqqWTugRdHfZNhE5NHWeh9kEsU3K2RsT9lbBs4SJEm0EVjrQzD6BQCxYyF5C/O
Z7askD0Pxhdz9Qd34blO6GbIMFdDfs9s/c33mqbzswdbJ1GBfh6HHtC/Y+RKAjFl
HxBdpLe3cZuMCsO2/ccDoB3aKnDg2Du4RG13xDU8oX2uFPLfxuuy4KoWPxMu7ryS
gQVeXSkEnXMhEneJvMu/Y07fKGLaRGp6jmIgeMC9UInXz6BpjCNWT1btVLmef/sX
0kZL/oPBaVtYQi2N3PMmfx4bFvmeZLD35L7Z44MVAZ/wcMCX9SG2jjSH3Rm2oIHp
Yoi9fhmUz0GorPtxosotafFmT2n0hkl2Bh01vSwokKvATeSChlOQRcClnVB7lztp
SS68ddyPExHPAFqrXQSCh4ChBfNVOfYUtx0XW+B+JpWYNqk4C7sufC8MVGl+5uzD
HH9pZXaQWySHAtnGNaDoJ5DUVHgH0JczCtJIhGF9BVx8+uZC/UlHgSfMa8JNxOTq
R5KLvj+fEnNixHTRtuXADRUKZ47qIDXUq2HvXLun3ysxjCt2+iwMZHmLzEkoJFpO
VNW2JQgGUvgotz++2a7x2yvVMKWtfGys2Y/VQPot2dZxAp4FQzm7w8rRGXl3yhlq
l29ApVWPap1TsCMJ+tj7hO0A2pGhBbd2OLDbVrGaYHrfBEJ2BKTxtIolF+qvEkZJ
KecAsACE0MpV4V5dn4J9RJchgGqyty41AxLtjVG4t5dee2pPmcTu5TDSOXpxZ0d0
D+UfxrCYMHCmkLzBxaSqBZJ6EAURAbVq1tf1gFXB6WwTsHXpHZs6JnAculStRiWr
sC4FWQTlCdAO8mlm8hUvNv0+u0R3SZxRY8ULVYp/aoXTQvTy70yGeaH0Muri83+I
oXyatUZJCbbHGyXazLSRnJxGEb86+eWGnTL4loksPpcvi/syh/o0mJKO8Vw89or2
E493ytxkyhJuDLrmjazbBgO+6Ze8C86yramLmpc421/kZK6bt0HUELBqR71Dejws
ftZXGWZLE6T0HpLJUcvZCerWBhK5fmWzGwE4ydgTLqpuKa8kj9Kla7fSa4C2HkJn
vJKunuSrvQnrXUOsFhVL8vet78/A3F+dT4rMqoL40reGyiAQhOmJATSTY2xTak3R
7nvy+2uDosoUe02+UaVsbYu9yKOzCbH/6+ChyY2uMuIOGtIVpS1iROAFAxGgEHwj
tbJaXA9LEHJiSqPmX5plhn3w3ZkCyStZSps5mAl2uy6zBAHvVVign+aHHyDxAnpe
pZCQSIlaZSj6tKBMQLesNouSjMpDhlpmltRILxB/D8s9SHtW/CRkOdmylGLrAuoN
JzGmSUDWQXN32Jlk+RxO2bUESwmYUVv/f0rcCrHUxNkp/yQqPXwC1nA64ErocqYc
s6ciCh35yQ8OTia2FUTxt5sQBSZ08E2obveCaGYfO0SZ4xjM7PKSNgzyfubNKmXK
RFMUFkjPuvu3UrgDXVzDvHprR7dsWBenCLMQLLRbKjKBXSh1B2HlLFj2gFjMppwg
tWG/lwUSHxx5dUihHDUygjtS+5wf329yLEm5KVBcpxztRyy5bSwoqgBo2+39gPK0
tApGp8XLC0r5liDVGmUqvXTENcwkr7c92+IPB6mbUZsnr1d13JjYZWFqtAxrdF4U
K+LSOaopN8o92te90BkJPJiPzQIw5gY2/UOu0d1ipRzRDNCi9ssOceKgtppxWJfn
QLZzu3SDgMjehV79pjmVWf23vJZ/eKkZXxNnPuJwpo6S5sTh2SpWTlR4/lO6KEZM
o7NrkflP3BfBkMTTtl6cwqVO5NdNzx8BITD3i4gy7aH5OElANA8RM9kkOZXSl+/d
hK4+9fR4iJTUT0RhXzLhNK70TZZXJ20rXChcjVwcwrfWtDPrJE5jHAXJM2+54xVI
jhXozCotXDcQKMuNDY6NZerbv5LMLHBeZP/x3VL5f4IKfZVOgcdiJcxP4JJjF7fU
EGWp2SxzHMTLyv+zFjUBtW4YD3CwmT5SrhMMbUlaSl79AryIqF0AGYN4l2HgeSQu
hqkSpWIz5tJA8CzIhovz2ab3wwTQ0L+7AgF4x1hRdC3lRvXjsvRd+zlJkgYq4MVD
sRYQ5BmBuuoqBiW3yYLR8WFxDtorJxOhiF2X6c3eBUC7zlhJ4j5SRDGwTfqEZpuK
F4GwUwhVNmXCmW2a/cpyPld22WtW5griJKS0cAroxR1GK7vPRNTO0AMg1qD+AMTB
ZwYc63t2C5ooRndJOT0nF7XMbDZrjY14f8PUgsxLZMcM5TMNU22wnrROhBUzGm5O
dSeFaLCZCZbhnZvdTawaXmT3vFPwmlekCZcDvJAIjAt2kfe914HMIg4gg6swmqIv
rOaXS2vW9SeqafW8neXYZVWsTsbsaACA6yuuNk7n7H+zyDGhLSkYmJsztKJAqyoZ
1kLPvp8hPF+ALMtNqGSWmqnNtbP2vOcht94fc92vS8ctrQoIgpxjn4O0eKs6fX9p
gmTN7ecJIMPG35fBuxrJPu5uUakVzlvif3cUGp4FEhghZgU5qa61XSVkIkhZozde
jm+f+B36mcMVzWFDYUcLKfoF3DaHtAr5VqZaO64DBIMvbfbkm5L55qiKTQXMd4z+
UARcHkjcof//vsICp7ECP1m3wKHhLV5tx0hlAC7p3R6OpTcncwMH+S3cbfeczJ8y
yb7Er8RpJVEhDq2Pn+7C/JzFg/YzHKiH3GL6evsg/1FCJlMQQFLpytLKav8Q4hcf
R84lN+uuJl+irlojuYxowrrtbugCiw3PApcNnFDu4wRyKutzOxOF6O+cJxfOGM5f
/J2MkgA2rg+bSZHTqy6260LmIGILRo8syG9ulz4W0iA8sVRwxRGPpSVYebGM1KF3
lJ8MOZAIbk6tZUhzHLsXCDltjFnWn/jKWv0kZAnYfv6NAwkeiyEnJV8er5dlWNrw
T9907pj7eCuOAmJAQpCXtcfiyHuQIJIfgpmor42HoWz7zbyA6y4JzR1DrNdBS7bJ
jWtOgdh6mBblVdLbpLHZtAhG+PfWsi1R28V7+BB/rTFl5LfIse3BczYyKlZQKYRT
HqgKQbj7lX3GjxzQue5qA8vO6nTmwAMpVbBrOCwEBalOA2TAukm7vBZz8/Ky73gI
BaSGVOZHhAW3Yo7eH9NTBTT3uaLBVenNCkfa5Q5tm1I8n3vemowUqbPTUR8nHaK3
yWHdTIah9MmhgcTA/TQ5DCybsfFTAmWQGGL1/LCeJu/vgkH4RWx+uCIR6pb9XFkU
cWwCXeCBB5ut0ino5aD5b4l8LbBs7j/HR1N9fjcYoK8ibAipeG0wLy3h5zLHJbhq
Fp27eARDNg9Fs8IxPmHaUf0Y5g4q9cMq9bYgpdMvJDDNaqCvuzbX1hD2Fv4sXsDP
6NKg1MG/NhjU0yy2ThCX0KjAv+WiUmAoRxoiUItLIpkSt8G0+SCzCxSuR2yAvqli
dR2mXT0SYVusD5ejKoBIf4+8Xdrf6HHJ44mIuApJOF+HqBqXTQcSEPMsxKi7PC6m
6e0B07Py1sJAEdSnZBWO3bs3Epolcdog0rZ6qVSVhykCtNNootG4vFPqWVC/Yb5Y
e0LBTISBVcqFc1ro/G41zHTwaqAR59HZAkZxRUYBxpUjFCLhmP9iZYnXLmfWMFTP
nVlC8CYQBR7mcOoCeKXXg9SZTdILkN9N0rTY0pWxexR4/v/7GqYNvTUMO+fidJNX
1CO7AK/xsGzOO51wkgVFkPB2z25I+HL134vI3PFBDwCmI8iQV0m0vQb1mkIysFMb
83f0YZNZSQyStkrv2mkf1XEkCiBJo3xHQf8jLSsuGT59gDGxFp8M/GpND1JkjIsr
PRxwrcQJV5OQ6OdXBUNbR+J6D4rjx7jWk08eQwJh1yx5K8ds9CVlG53zXaB/CLDv
TcUzv0WhQmuwhPCD583xOxiFIBGfkjnmLALoYb6u47G6PZUb0OotVMb9c1iVkWEz
p1N8H3UnEmnRAwjxZne1lgGKVUZ3kBCXvJ8Zu1aWwA2gA4Z2ZPwqmN+8wQ0pKxpc
jrDhR8H+FcCTdHEkjoUym+bI+SXI0wjhywKEsGQMSsnGaT7zZ1BQ1ZpvFBt09yps
ZqcKJgC+KEZ5UKqGI9toH46O+yA43zL+ghcmidLUu80K1LhKaemay3qijVJNxNLA
ULRFLa8PYh5QNH8jKldZTwhMLiu6gKk0aE/wtWVn54xeOsxIRPIcPY/IMMC+jQ8x
uAptvQWT8oDPMjFyDA4VctZ3NbJVFDTwbwSa9dDXGskt0fgWgpnufbR7tYvxjLCL
VIhP2hsQ5TjQ0OTspSj91MFoU48oiXTmDdNRvYT0sO62Xi+f8sMGYxPjs+lBQt/g
woiRW3uKrfLZzEcyhfnkI25zU3bSw8JfrlxgmuXitfWI4GLauKe9gOCr8ZSc66ki
1IwBjT+k1PX0xksr+ByGZpWBq3wdghi+GHkqr2qSLbiQ1ieMWkPSabqSb/57gi2n
WcKSMYuu/CqQWtoS1c35q0PnIaFzLPT1OL9iXeK1TudHYvLMuvMM/gUkfobd3xJl
OVNNY9cymP+bCztPWigfPcahN/bAwWJ8aVMWYnYdSCx1LWhOAi7Izkik/PJsJN2b
Mp5qJs5MlfhVlxwrws8AAScp90utc+S7X8zFHJB4LyeLIBM/tSR9bdzNfiNF0lBa
`pragma protect end_protected
