// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gYGs+f1xbjvagOUlaztKvc0woaD28dXC0TyZC9yoAcvqnK9VMtNQnaT4WSxcjSQi
cJjDwpkee4SdiGpkGKjIlBB9M6tswD9XaruejfIRS+CM6ojAEmM3qyyU8BAryfIS
zNl/6Gb9J5mL5XOcJrALjTp5E/v7IyawhwLHTiUqOLo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31104)
JMPPWghCZxGDpaFwIOpWYTOaKiYJ5gnJqmnGdp3iW8eRTOfaliv/nFQrovYk+9s9
//3ATT1MpsI05vHQ3SHS0WcwgdvLW3+RDQP5XEr66M57tyoTXdhdM/IzpvKS7t4P
1Uiv+ZcEe4AfRJjB5d7tFPOQxvSQekfDh0ljy/X1qfndshUrQKS67cJQyfhfv+QL
hn1q/zJvm5Dfcb9nixnzFEPtej2qjhrStRMED83t6CuRcQjMVG9sH/QMsgWLeFUt
m8kyuvh5vXQNx4Xeimv5vqEOXgUk4XNn7LX+yjAM4oN37Xz5o681+REA4KiCyehD
MAJHPtIbrsz0U04X0h1stxSDCWK5VQCPsWLJPj2kpSivDFLkjXZJMh+jtKH6hKZD
Vn80zMaMeOVyfk7gRdPq9JgZic/bVI5et/fuS7yWSP4WiZ5yChfmBmh8wSMcq7Hq
R412/Ft8K+1l5SJ8QZf70RC686SclwXlF6Y4QRNeJVtZdJjQ6frx8SlULV/H98hg
/QLXjA3xpm87+LwuH1r/Z2pheb9ajyB9iSK4xFSDdEbs+Y5wgvAls9CQZC9ftR/O
BMEruZwmzJC58xbUDoZC+5nTEA+u1iHZb8BjDkpZlivHMR3HWT0TT2Mxmr7FlCEz
5s9cUZ5fkxDpA00lTphxjgUHd/LP5kNQnltNJpul5UzSkejdZ+Hfom7W+ChEMrvP
6VmFf6U1izcv5cNaWAjo2khrT9CNTdEQwLmsqx7+QxsNs3DqPp3EX29i/IOcCAQi
/lfn8Qn2QYN042yTLAg4mscxvsMfqpA1CqtfQWwPQER1o3dEK9afVQl4io/ehJkt
jR2wlHmBM0zJkCOGScvmlaOZO8iqKARDcLh+YDAhC74lmVyg8ubzVznUo/gh7LGX
DBL/ny11qM4d1XOCfYae3zbKIcXCGoRecbRW8/yM72ozScPJjdCBF76i/uar+4fB
Jn++6WBQ+C2GRtHPeXWVXfafFNIdoopStE1TUrsemfUx+LQ2VikS6t4zhlqqJxWV
HCY7LyIfGLycDFXtOicol2Eql399uII1I0yjfDD4JA4XPxmJeJHv3+3tYODIawxk
i3vbnjfRDC/Ukg9zINjW4MTXKrx9On9tAVLV580b9S6hULOEuIGjM1lZ+keBIDsf
ogudDc0SaxPE8E3aLdesEZ0ZKCN2Qislb6ZZ+61/SD0zNSwUiLIUPHbzVO671vpf
CEoj1qGP6C48s29dUr8sNZVOTB1NoqvZ5maVgg2OW0ya/+iGZtjGoSBi3aNifuvI
A8IzfdB6KZURvpujWoQk1sLOnPWdbS/q9lz6zF/hrldFn+kp/7orvau1+/UcA2R6
1d/+amMk9RyPzcSYSpE0IcN5hS+ob1a/aySjB0IKIBDOCvGK+G9N7Btgu4tHqHVX
j3TFryqFl4L5ofsrzr6BHkZH80q4EVCAbVAoW1aghrGBDQd9widdjGwuAIz7HTgI
Ln7gqzXJOuGlXhF7szrFGdRcbjE24vGAgLADZWUTlziWe07guXndTI9IRxPaDGnD
6vKfnkIp1CM2S+09HWUSY4+JGufhjm5quLwX3BXOf1aXMyt77EPWQUUpn6Td6UZP
X74Cx0qZMUCkcmDxD8fKhePc658ucUGnqX56/dXxMj713tEOiGHfHj+bN3LK8Nvz
nsE7AOBCZikg1fvC1KBtlM6UltJs3tHAFVRP5d51WjH9h/7QW5lKy3zW/DtYixis
E/mGlo88v3t4k+5UH2LeQU4gZ5/If12RvSEggqWhtF9IhS/O3U/D2ihUnagb9J3y
0IlVPcKHfnybrbyOkkFOFDjiIddTfyQqwMmu6BEUDcDCwoF/2CnqX3Mcu3Bs1f0F
4YiP9xUrehJ4te+IqWFTh4Y6mDkyHLx8kkQLH1JnRSuvj0WmZ18pchD9qnsc7hcv
qabHjsLUp0Bjp2rKnOfMXd2v2VjCQZiOOMf1QO5vE1luG/z9figw0KcFboRwyau9
xql1RhUOG3sKL7SZ1vqm6I3Y2j8tJUIm2UuML3jt3W6HlKwJZCfMp7SslB8S+cqY
neItQsGemdxlO9OPqAcjuoGmbFYW9u8NRewX9T9CGJ7vrW1LAFG6Dd2NZ/Egz6mh
203lE56qnUY3CKadawELroVQTN8LGUvlR6O2yH0dWuy/ccodaxE/EFAUnMbFezcS
oSBQ/9hieC04ywC8M7lnqACtOBb1u6+X9sW2DSckrMCKoH1vJDlbdkiHMEg6CYGq
z1SloubKKnJu/eo6Pt9/pL90sderVwtEccVy9dSrcEL5vm7FvjTE5FhuS6pz1nKg
FXY2hDGq3AB2P7q5gh/XOwSKMcSnEowXBhRJA6RJcXg2wmhrCyTr3BqsmL+Lw58/
M8jMqw27SJCa2AZOxMrlYg7gYA6grEYlOWHW+3RjIxpFiU4g/QTtXmPPaBAheLgn
6eTtgsHRHk2GH6+je3xp+sm2+LxHGt8Ab6nQhBH2lvZGS588H1a7dm55zYAmcs6o
3WdueaY2SdvEm6Z860Fp7lHo/+omcYNz7wCnx0f+DMEEn0DDvn3dpD5toZNHSJ1U
vqKSVx7JAJm5c6cdEEfDmhGJcmAUDoqQ+nXiMeITa3+llNs+6QepT0ifOCpkfH40
NiyzQYI/x/DGQ3JXLxv7eCd8fTGWK9ayhcXz4nN4aOceDt1g53KFhTD8yfXZOnUU
1p6Xfj6lmD5KGYMZHbIexly4OrAm+rkz/QZsFJg2YNmp4VuuPJO9rYnhiHO4ZpjW
DZ7owePnmZMKr9p55fuMAynOaCq7E9yaFhD8CnVUhx0lhAjaCe/LfRyT0PN8N7ED
BzDfi8iZ1u48pe0rUmERkEvsWnda3Vz1pjLdMLi/da9Uu2DDeuyHiY+Be9sbydKA
kLn/ukNYIRplBFke/ySztxDkhfcVp/E8WJhQPpcvNqQ8aiT1/L5hYLvY+k/xwUtu
O1qEsHVT3BePtcrgc8hOXFqIweflIrVL/SH8oqMGPcdvB7o79ogOdNCb1LFhsjLD
4KFl0y1Fn0EWFnVU557+VGUk6K/rxCB0uCzwm4AuEadRoANHecqMNSozCINonk5d
Ur4bDaQO37v6hObVyltOGWopbGJ0+cyCN7aoVRG/S6ARHvNA8LV6zaAdACxX4LTe
5LDOy15s5iO0mezazBIyqaW2tngVI+JleW/GCYMwnSOVlaO21C9GUcLY/AgdfQwB
eOZqDOyDGaMNZGsBfVylJBoGKlCP0macjkeVw1FicK8ETXK8ym9xa88w5ZH1y2Xr
VgmeoFlCz1DZ2ADEyDh1bJ8qkgejBXE796n0Vf0ENAarcuvGCXqWs+93mPwgBbyV
z/UQ/QE6Tj8m9AtxOMTkIt6bpWB/OGWv4Ve4CcS8gJ9o6x4FJ/17CRaDjiKwpUqq
hDRoWeSZnK9dFbtcGCPLDP4pjDvXsOSgUlSMmNxATp0IAyMc7CTwqgox6VgqWajL
e/pf6EBD2Vv5aSv6tjD0Lckn1olegHYhhTk1i/l6xSJHTYfImImeUKTvTNn/vcDF
5en5BV/7JBvjVgFUni5srTwt7KhcX80Zc85nEz6kcGxy1SwpVhDSRxFfKniCD183
nmiEujb3G4+eSEE/1A0AyXcI8rFlQuNFHUW2zOAYJNpe9sY3GrOMzviAQFpAL9nz
TvAhQs7h9sB1MDvwimVwbg9JOXolGfLfatpF7rDizD9JJauLpyPiNi+LTrextJH7
j8DwhuOwsYnqOcyKmtRpcPlb1lDjd2N6GZci6HekQZR1PniNjqx3DyrGri5hwjH1
TOtQyJDNE+XAPln5XM4ZOOU/OfYO5MB6QREkRC2dFqH5WC5pzjBDK0ixIXqFFb+L
RUXycuivkrpGWq9ytvPkgPzDoey2OM3EB1K0Xgn0RCEWlXPDTr0PlJxW4C1yQGPk
X6xKZTtCL+yXABLvKYsZPLlepcaFmlbd9nbXCvUcoRs3gHmVnpsAbG30E2V3ASoE
z1GXSavB+WNsEe8nhCqTfiyrvOkpNdsTEAXWgcyUlhCgloceb0gczi2dkZGVvvFI
ZRlsHTQwzLih2Hycupz2TICYP8sqzaSvNtfLQ6h/6kNvD1wk//5hAWzve0+Zr0gY
e4MpGo4x5y7xqgyID6MIVFj0fzZd5/Oni7bY/6akD01NLfMQkGHUZh7VC7s/F91I
N6UYH72buOJZ1X4vZp0ZdYGGZl8CaCSEP4AHRKis7FT7rD1NZJk9ReRy8YICBMxr
M8gteFaGLZVWcaYJp5fvBF9triZMwfogFMGVkAogbeXHph5VFOb2Agr64+75umsO
HnvboX6qbezvj8721cebfrNFJloLFyxOEHwlsGRS9jhp93DsfpkZ9hQHcxmrX5YM
LO+u8guEBKCLUkrJaHmKvFkAx4z9Xv6dU/3f4vAByNBT/b0ucSp9E9Jy1paAZCWL
unsAIdVgYrVsIxluzT3frkNv6zIFKXmwlpvxM0F6lHf5fCd4WX7c8QxQ79KzcIvU
v5FMvb6eX4iImOeV2IXaldreMlaId5GJxlW8j2k+rpIqAe6kMKvVCQ/8REud41qF
0bF1ljfz45HJcfuJzzOOr6Ky2iqEn0BQBv49EfsE29d43fL0VfWqpVRh1U8zwTbA
CBxA0xs+nSh2R7VU88fi87GOd7IOnxg7p5pHExzvuFPUoc3fTNiDYrpohmMse7pi
tDWLDl4N3uUbd8kaItKDqHT60tFbIPIGDFZRhp4DduQYgsZxE52wtNaB6eoJhxry
AIlYuNr+KfbcXn0vIfkPDhv6OWLPV9Y+Qv8obmG0pl7oO/ASZAN7SVzGcPbByftu
mK0DVSb6Mg/rbr8Ve/OshSiMvqZDS1bgxt1MDN9u8nJKron3EV83yuX+nZ1jZRR0
juI9toARFO+GHI2SsD2Ag0YBqGc8x0JsVgehgiIQsVywhAYbvToZDgcuJIUgHd/C
IDxGPxMSg+0zTkKLrVOStrbxH0UgT/vwHGj4l0dGkASvqRAqXf4C3dJBH6IaUxrh
rl2FBBruuFWX4GBVOgA1enoFQovBnSZZnlvByU97KBwNqI+VGs1UlHe3/FYRCCV+
/ewWYs0N/VvB0M2kOd9GzJylwgK8cczjfxzG4wH7lY/kngIGKurud7GBLSGU1ycJ
L0enpOwcyqLwnYEzWp39TZR4vIoV9T6PSsDYIHe4of1ArQUoxPYpUbREFMj0Z9F0
WbtTRyGQknWwReKNoEb+nzMXHhW4WEN7gNH710LnrBd0VSYgrJqJUGfNue4OkYuW
BbNY5f5unkZhD2KsOPkqppeAQiM8EeoOK35+/H8cLU1pQV0vCTYmllS66MO/8lKn
qoxJWSKo0DKzIA5vGhZHED5BeTNJD1xEokJmqiZSSHxrXfyKNhUBJdCIDcRBpiuZ
qP1bx6UCuhHyylgNVpBvmSCBorevjXtRU5pBPNgVb/LCxr1/JhGwkHhq8ZSxF9c0
Yp8NSMJ6AG5TlXQVQxFywuvzM5zCX9PCw6BpYpoWuSu6UU3a/DQwvX5AODMSJdA3
+G0hZZvYrE3YkM0oDzgbB+JAp/jWhOklAxJfCw57anYSFdygiMhiVoslm/flldwV
VM1JSPKOiigG6pq1YAlSsNdijw8895zCYcDoLX6UHfHX25dOJsEnCCYvXhG75nuO
FOnbKWoHBxGbHAax5vcjX32kaH66fgENgiVlhpAEjVHJP5jxuIxh+JhieaoPzzgH
5KzlWjdfkp3gofnpA9Z1JbTJzn7YyPRLO0C7nEuUZs8cfoV9yhkdZ8gcHY1GYZpX
TrL3/Tjg7ohtNAovyfPZNqsUYtGbHTA1+XlLMmzbkHcFblkoD+HuOAdYGMhHROYH
2ljhAtMgNWyo+tQXIIehZIJJn9wvLNuYSk9bcOwAQjuKG36I6W3b6hV2gribjMR8
De+BwQrmAuXbZTQrbx5mz9wgrDd7pKRoHEm/RPP4vGwlpDCxE8u5bB1p5HP7mxSV
cgpGG4cqy7kGlrMChev5cgWQF7gEi2hWVi6fFts9yM3+fmvt/k/vzEfHJs84Z2qR
MoySrLKqCc0Te96idXy+exLNEMe3wZuH3pCyyd+22qV9dB1aqWTpeOuPapigAGYB
6K1bODi833YrhV26Eb/rQyamHXVlturB175lkDyXvs7koMTUUFk4jz6PFsx4oD51
LI05V9tpYAmZ98lpqVf3559xb5Cg3nDqdZrKjViDqy5N6I79SBU0wZTW+OOtVJf2
O6bSfK4/riG91GEwMPvR30x9YycopU8wOsAJPSDbuW2rit5L6LMLM/u+uAY/3DfZ
jzX2iSIWIQU/XS1A3F9e2lN1xz34W19/N57MN+EViw/y9ER+5c2Q/4Up/aIC2f7g
4g6Bo4660vxukwFpuVVp8LNIItHatDGRj11PcIgfEs5Kt4GeUzk41aJpi5EO6rQ1
c/S0E6vY32SWD23OhSG/NTLNbirTrAUJB4faHAzdgEyBIN7w9dkLUnaFV2zCGU6O
UmhnhzaBhRZZmUPKcYQiBiZUI8O/tHlpLLzEk2Q4SpPZwjYL/peV7GIKvk8YR8ZQ
Fix/9G/CN91XfQ1GEvYMQPXYwOtTW2F02zEuZjfk7q//zX+gfja1RaU6qQtr9TqI
9GTqVKapGe0cwe6i1p5Af3+pxg54jIe9w4ULoJOokb98d+uwvHDF0v7xAiJO94OX
CSZUk1Ncd8Bj4A5urRF2gQSArFTo+JW2D1kpJXXiltCtBN5IC/LdmUkbmjWAvtHV
iGYBqsURwIALroZzQmYXRLzAOKHIY2lu4U9/FgRdny3Esm64zqTnUJ7WDB1Fz5QV
faU7XtCRX8WzLJoCyAmUpFbv3UFvdzcSASL/415CjFRoJRc55tKdIOqJbtx02ZJa
n52XKjIOYrAThG6X18z4tTOvraKmTXI9r0aW64rIcTjEeliQh4KpkpYGCqVK96UH
JVu5x5Oyzz8rn/2WZ+KttHyjUC5EnLx9QjMTvAxwmxn5l6UDmPLen5Aayx+AKTis
z4v+l/wNIlS67kEhTRWNlbqWQIM4F4OSIsHoyFoHyfzUHDBRwoJbw9oY7ILzf7rv
F65w27r6IMgfnCmZm52XhT+Hr1WLXEYDlb4Tt/llaF6wv9LG8lXXAaAQCXIIYRZQ
bYmtN+G6iXCQ2DvIdotwNxv+I9OUnzgTULCowV533Rjo/brfmCEXDL31UGlJC0Yn
3Ud/Wko0sIGY1Z6++PkJMyNXmN0lhOUBPKIjrbxR2NKh8dBaosAtcZSSCrOKvfo1
48yEjlCOhvlDe1F5KUkoJ1k6QdWq73V7S4ExvXxhbWjlGHKm8oI/nj0bFzpiMKsS
zPRFIvNMD3wIOo7Ca4I47hqLNOGpGSXawiWjKFHKXiEepJRpBRCcudj9+Cyb8Coz
R5lEDh40ovd11hRwVob9Qn1wX2G17cwJwZt78odVwU/dUf8X5nZxWGyqChYc7aL6
q5FaiN1aZSQR7NxUN8/boKSQIAENlfxixurzjRQksG+6tjWK2grMFZVJvrG3KEub
FVguIV88plClsBr0pZh7hRWc22wnOhAdhjfcSKfi5gAcT960an+d17ix00/r0wMb
htnspI7mGJnvZgYlpBdGsdTfbNdMQ27OoxR2212Snym/l3rFH6egDx2evgf29xw3
gO3tc2sr15RrsTGoVYx6+Mf9HRq3AsGyEh+EhHrgBUJgb2ncjT1vKgx5vx2dUrGH
4rCntC/aMViSyj+ZDTm9IU99ngWEsVL8xTUKu2Rl+R1xqMDri2a+OuGHzEO9Wudb
c6oBkQak1oR58TyCRQwxPS2rXQ27C6GW6JasFsfbAZbqmm7pf6YdiiAKvSj++Bzx
Hl+8q6hIDItpfPaVNDgR6cjKRaXAEPqgYul4BOsjSH9Vjo3lJCpLMJK7b2LqHU8F
o8Pny7RlEtKDeQ1WNzRnHvDXvEna5s0+uTcHN1m+iNX7P3lw8QNg9yVZbY5DRLKl
yRvi0Lh4+9UmyrsDPKPscibQTEmFCLOoxYh3MqzaprqeIcwfNuaNLenZqCRN9lk4
Ulw4l3d13PlMmwwWlK6yoW5gpBpJw4v2LQ4gBqoG8Ns5xvn8MOVCh14HzdkYGWUH
b9MdJB5jhdG2ULcUxWOBQ5coP8LDQRv1rKR/JGEPD/wtPHPoPkCyPfK36kkYmgTz
I0FUD//vcvzdpQJHwagLx3Nj65qcKHBLIS0D8nU4WFH83WDE0/L0M6WZXqcmIRTO
tePR5vUv67TRy2vahWg2zyrV0QktFx5tkItQtKDpJo5iaz8Xp19Km5rh4hoURFiB
uEcUXt9GdlcvgPTMMFdPLd2uFgurgwVv8phF68TTQ9SHthfHe+Jf3TecJv9ekJHA
36zSBsTTNtGVY6PtPX8f/kYt2C+r0eqTaKRIksQR0MHFLROKmEgrR9ulUA8PVEyR
IXAVNl+nekHRCpnPWU43U6d1WC2DoDK/MSFUpwVV/dWDG1+JtsYO0ylSA7LU8En4
DRq0jrvAs3ndovRIN/2RrqSZ978axLVQ1jnilOT3LD9txNuvRgE3EgmxvmqBX8a3
ExCiCJ+UHZkHzVSA2ea63vfnMXDQaNY4Dgfxa+N1d5KWl4IOK3iWn/moWLmc1MSN
dAVRFftWNCk+2VWaAQftGXGI8I8YubmLWgdjGNSeOpefGqWoMlZYxjbO/Uypaan9
42K2s5edBTrl02IFnUqUf0U4P4RZFplvbZDbLpFb6knoyTE3MDx93D60HDMUpSdM
h2WHaz/jktK7Fb2O8MW9VANJZln3jOIvNKb9MAgSJV+vMouw5oRXft7y/Y5guTKl
kE0rk+t+VyiiBPfmwWQ8ct5QYtlt/d6DBRh2ovsckXR4b1+UiadN/WwcWTyynvVM
yM5dhMjyVFjhvO5LHg0p0LCBdSWSeMxiiQSBUsKX4lPEx9aGSkjj14DfUuSZmK7P
Bxo3E/Z1RTLxcvbP8uUydjPfzja+2vRvOXD1xq6qr3zI3B5zCh41zKLxssbRWpWK
zPEJMTeXAJfBYyUKmsh3KmdXUKZlfIdDV/Me9bptdBUm5gSXTlV3XxXi7h7U45m6
T6nz5B4BfLbXwBPKq/rnCuPUySevowlgTfIS6hIoMG3NFSHIoRJ78LP0zvXW8WYU
W3qwjWN/fbX1G57fMEb0lPZljAzPa4e0pFgyM4q5cHSxkHQQCHUXyQ+ZhIAFBb9c
aVcSoeMwccqz6+FFBcfoTJXCBZYbTlvCbun143PAd2Up5abEiGGXmB3mMKkIUkKL
PueXev7RRi1Px0JkLFZL+h117ODp55gMzbXv2XVzkSbabzgrt5R3ocj+cttGgIDA
PKJmOMqhlCc7hgEKWR0vw84RVuMk8KGOHDXF6JNYwL7/QAdllcGgtOdm0kaCKkui
4fJf0jcMxwhmDQ2QhXQXQenDLhCwGoHukaTIv86arVVbFPZI2XATtxyF4T4N7Z6H
/M66+5hqACouxB/wasRFp+HnjLX3dxp4E4CfZOu6ZtgRnGUk0YabokGBTz+2yfKj
LS4aGVNSkVf5BzEafRr6ENhmqCqNIgXTlspuFA+579stlEm6veaLZvqF3OptOGE2
vBq7kNmLNKTfsS9TvAEbNCsT9OuhqZY6Gc8dGOoU2TwKLIyYG75ItfvN1/GfHW74
MynnN6X7M4YG0x/vuf1VxX1W1SmDWlfKbeyYJ6hRL0XsWUvnOElWMn7YbZBK53nc
WuiFCUAVWkP+RbAg6CRNn7YRdXrTjVeqHEEGZG0uTQ+HTTicAyrGcHPmSgx2ifDZ
vuZiO/Ic50VnCCiTq8jtQFQ+B+7zvH3U1QIYpNHlMN7+W/Ff683tHyGAqLxK/+kR
2f0dgEVgGrr9DKB7s93TwYOvuSYLmLSl/n/GUPoelda+rUnv6JchokyGKDh2CepI
1hZKDfARyKvrLJ8nAypUWqeqaT6pbwi1lSSMPwsodNBOrMFT0U/Zs6+rmmsGPhqh
t/Bve6NX8fcvU3O3WvIFHqKvVbx3YYYOvD3n6R/JPnX/hMAmrDDjhcGkTmlH7aOW
5Gm9HwFdMSMlvblb9a2a6kMONMzz9KJwyhOvaS3AzGXfwCqq4LVcu8lP8fj1kcbM
5V1Zfpsy+A1OhDSjjhwcS/K5g3ltLLo22JJ/6LlMw0BZWy4MRWav29a2Ejfmtbkk
J+2rcElR05nN1gBc5cQREN5ZUhsq268Q8kAkqjQIyBJGhK+r/u066LwSrfD7RGxS
BjKq3WZBzh0zuNyG21eCmCKAB03QfT+HQAauquWa68eZ0d5Hog5CJc2PDXpCZEH5
neywsKuZf+7rx/YWSumZsPBSNktM+p0xXIRq+Ao5jlDR8zIObldZJQeLLD28Xndi
lTKcoin0J5lEpcMrwu+xZq7h+c4mJdOcEq5uCi3iwmWqK2gr8/I77GXHBmlTrrI1
GM2UAizZ7dF0ZBZ0aiHIeOp1muttoYSgPoYvO4Hfi69MsJwOh3c8E+ZnX/y5omX2
pI/xnASr4CaVawMlzxvolYmqKxg2O498P8ytxZOr+qJW/UxW0epezXt4Um8cIDUO
yH6xnNlvgc+iCO9JVANfHN15rdSkv7yFm8wdyt/6xcQehBU2GBqyiu02E1hlxbO+
P+p/aTjLcqWcCZfwTq71Y86xGFwn5i3F55+XZUcvmkxqv9Ost1J6YmnqUz0PV2i8
YEAWB9YE3HszgNV59w0U1kce4wTyp2B+szUeRZBecFnOXo5nD/WjPw+mRxI1jGYg
SG+HsvsDNTDPczfxCXZgOlZ9pH05zRUPAMcm6P30v4YgIdnobI3FxnzEcw/YBHX3
nPpwpkjbeNOWbcXCvEIUNlWCSrGMNwJ2KUz/HiFEb/9NLkE4iWmLxorxWcrCom6z
Jpkpu382OOrPaL7M0kx2nY/yqIpUoI31JPfY+LECTOWyusMlnSbFQ1e2nHYOKQQl
qJzmG+ixqqOxQov7M69MbLJTvp5GM8ALtQpNPOXxOB1EYvQ2+1HQkGlXWAKnPIYC
FNN4GHfZdafRGQJSx7Z+xAZUsz/nRE1qj7FaeA1aV+Xfb6OJLqVRzzEzTRVhuiYm
eQW/puUpWgNZqNjpOA39o48M7LK85TLrhRMbQP1++ZbowZgBIx+byQB0qXpwkf1a
oiHm7wAgHLTw2BQFmJNlQ80t14ItpOV6T3o3fy3IVpStFmeNW2Q9wmP9gk55v9Qb
Nm7B1OFEc1No+uKvxz9+rDc+pTFQynB56l/3BEU9KrfOYjDGJfWe0dX9acdOIacJ
67H5NFyEShOVw8GSEiMKJmaCxmgv5CHgEUNvfcie/ouSKVtxs92QusZM1kLI40FY
FlLsBv+JzPi1OUnpY0a0DwUgT+D0cz8lH8uFsFroUftT5MvKn63zndJkxzBWmdYC
jwbF47r0KpU59tJDDXPpf/rWUhgLfavchA59lSbDN0LiHTWrEMs5zWLURCCpie2x
kw2hzJA4z4OF41StYYYYBXShCbY4r2Njd0mZXIHMHhRC0WsCObFpm5+wqU+RfF6n
MpyyGTQd8hLOQ9ef2BMc4bi7Svjh0SFXYbpEhcl8bMzePgk0rEEjXjouKKWfLEM4
YDdXtLlICWd4VNzvUKFvr6MnQpNMninSEimkI0kbB6Qq5Ew68cPOJC0g36/mW+bo
bCXXBoYbMsBVCc2qaZCDFXIzD964jkpuND7+FqhHI2LVNmiuI98EJRF3XI8bOqqC
Rq2VmYCsVm4ZA3+zVNru+VXfNjlfjn9K39Ri5LkTEMQQUbzhrTMRonO9mqjY7VCK
5zizow3Ly+NtBLK8YZPQvxlRIbskyhtBUJZV6BcMGxRfQD77nghamKm2ZWDVoPXx
AWzE5WRshxbd/Qo4bRUvfvALCFGU/l/ZXuWHfkONn6UaUlXZ+vq4r6/cWhUKNYlB
U6mpzl4RRHIkMxUDDLLg5ciobRVfbjSmhLQaEod5TOL9+QZivGdBS+pPl/g5WVxS
o9hYizDIU5LpV0gkHp2ot0QQtokFf8JGTMZ31z2ATcORRivBDPTtL1YM5W8Y41TT
+nMOq0kCGmIbXg2IWIKUPOSKGSxnfA2q00UcOEfdtT7LHjAW7MvKdl7PRNj22ijF
rEggNC2u8Pr3cPcOk+0QrFuzBXBoVjZ4umoBHqYtr8ixvmwaDU7sWtPToyEulHWV
vLrRwYyylG7c+DU/TG9vLIf0+2BbfUws6OwPdFukikiMGxe7BLXwExi80mCYlYUx
+BI2V4ua4gEYKrkCOMBMYd08A4NLh+vvExZhBR9XvnWbDXb5b+KmT3nr2GuzfHBS
nMFsk7sPzJXZ1SQ4WkBZLydMh9GxTZbRK1P094UH6Dj4hgvaOuYDbU5SKKlopYBI
nPRHv6Raijp64JRXuYnJ0uSk95StY7+AGBTnNFNZ4yX2khPERbj1RcgyNeZ2G7CD
MZqBCTsUGnKQxxmo5Bu+1PZfIgEeYHdZJqR2gaT/eEY1oYPV1AtXSbFYALiWHqFd
plqxXRUzq7k10y1mO/eYPmnfQMEM3L3uSK4b8B0PLK3tasYjLSyut1+72iL67Dtb
56ViKnCcjU+QibA73WmqDuJpjSUzTUbvYaIwbXZICsgr4E5Vs/bT9F+C5dCB/Nd6
hrE7/7vpIhbBAMuIip7QRNBRSNbnufdSrqHpc2CZgbKLlQjDf/7tLjaqqHSHb/yP
3690ERUC4EbRcTJ7AIDsPqDtKrcncIhdVjUulvZIKySY8wAF3GW/NFmk/htl/js6
TVWntR3JIH48SJ4oaJLVMyQOYrm7YasYfCV+LiYthBHtqXdHKuA05Lq2oTK3/gQA
nH8d2v0ea26kuD62009Qw6PVamFz5lPVCyH5TQO6HKjp7TW0xfA9UuaHQt6UBqnl
Ce4jWtindTKYuHwTCZLDXd2JclSrW7PneKfRGCRAegNHnbxcr5H8NaZ32fif34+p
xkNr/7OVpjxduKLpbIJBY6o4iDrS2hPuzZhV6Z7LNzdwc+ZXrIasqCpoLVvNojie
rlfKkFoqbTgiwp6uJi+t4EWCmAoNXxjfl2CF6JIyqnW+xfOUfKtnKGKX450/bJmk
VJ5W885XrdlSYQ7x0udprD5yaS8I1KKxxnXMi2fj97X0UlADjMXvMSpN+munsPvP
9/EaqMZt427emxEI5Go3zlneZkc+Igp4CB/0kQlNvoIW+QTAZoGBYZVbDzkKwgSN
IqTZVqWTuwTz3tB/H1um+TKJkzs7YLrh8yUoVryfAPuCySfHP93mgTvVbaRuUuwU
JiEdzIvg8+ELHfgDQzQlMzRJBz5d6l1+QSencbn//bMJcsAdxVTngLsNS1L5/i+o
dxv8ymTtZXEE8ZIrAMKVRAlmMB3QSkRM7tB5saqihoin3zkj0G3CZA0/bkIQxJJV
2v9VIfBu6beXvcEAMjD54xZjDh5Ds0ULO0ETOayGjCI9PzbxSpLWCARA9Uo0A7Ex
reQ1A+UiA5xEY5tCmrZG3zuJqL9K/LLS+LjRUplDJG8MgBAWtzeVSBmrL7G/E0mF
0VfIhjlWK4bd1MaKl95HHzB2tXHCyA6Vm43NsmS+mqYdd9lVVHVhcB9+xWYwVT6x
ko7JVoY/rUNsIXyBQt74pBMgW7vxUm65/A1nXXJR10PYw/yihGPiFwWNP4Xdpa4x
+QLDEMOoTE1g5L57IgrFuDE7Qjk7/H1yyF07HfB32+my4Sm3Fdd+BTPGnDN6TW63
zGUO+1OVn5TJ9bL/cyFabQIuFuOlxZ0jXIsyxoBvatB97WcVNvc8wbUrWT2hDXbG
OPGTB3itXlp+oI4GTJNtTfZ1O+bJ4MPL8OuF0eHbDOq8pbu3aOnCPOvbTkgJE1aE
x4f/PPBe2WEQT+f52gKmWX3VxJNSpvxL+9vBDv4Lcfucg0+CRQjp84C4PLMiEXAg
zYXUMNCmx5LIZym3JoThD6XmIphF5SdXY6P5Jn6lCJ1ECXyEJcKz65Nlwam0Cu9O
5N36eSEMLUhfPdRpCNRvSdL3UhF3CmBrS9BsxSjp3sOVJFdtibgk8iw097UrXFeK
oDRewYnpeSU6n1gQ2NCTIzc93Zzt148vR8b6ymr2Y4iTO6LbWVXvhaquPDQzKodh
5pnYdxJV17NDd71G0+ULDr/Qjl3qzifyGFkjZtrVw3DcL+gdOZq7oP6jYT5PeA0V
ygyAHxomvdXB7RTBdZfwLZ9jGpvo0uyeSDQfBcVFynRGPvfSGdaB2ttycNIEKIlE
XzyybZ3IhB9fwQjBEKs7IegAN2nv37YrrnRqB/uZC4KQv4QIbL5n38EMZszArmsh
pcfo3EGgWOpMSCOx7vgHWXZKkyYqBuCpwZhadkilXC4DtfzFcDmm9TNIIyt3+NYg
+PU0dtZgRgEKvXUAaBcc/lRk1+PgOhp9PyC1G4SXlzfZUx6JcYeb8V7MUqVAiMg+
WC4HrOs3BrFRd7/5QVRuiipHE8oKFRhz3uVwHmEbanF+E8VrFHqz6yTb+qEFJ6kf
QEbuQjQMSKw1uZ4c0EOUmSmuafg6wIpZFA5YUm58HWWvL2QvB5oCvrB30XyQKNRH
VEMGalMFckTBhsWkGCP7fcc80veQ+hJvfrvlysTCbsa40zTLVjwZp3bX/ieHq5Ro
TG/vfQzzsI83Vm9CoDsLHFc2JHgyTzQlJpzp4Sd3eojVBPV9fW0Xgll/N+qFols4
QRfXJsyhTuEiCIf/Xaeing8kc0o32c/fXmKaG3v6DrA7t3RswUevWVEKiM92mfox
A8mdD4iQR1sHkbtScLXJduuvpqkCjFOBa5/B9khLPohltATCirGG7qxoaeIho4Iz
yyGfNDbSg3eMrIFCoP38Ao/1zsBdVOPVPdinQdy4ADtotQ52iCgYMm/G+kanAroW
cjrsMges8NPkfVZz1p84tz5MloGzUmZAiOPGQ9gd/ZeEQ9U+jdb2NyLN083K1Ql1
NbX/Drl9Um9UyKFZ/n5/9iH61gTDez8idtAD9a4Zeqzl3RlI0pydqhVjs04L0Z4F
z/1W3yPyY2C6ciYSxE+F3Ttu1TT09tVnkUPhB8B8pRvOORldN0iAc91PmpEVBvFc
7pu6HfGulkbZOyOoofvbhkbTX8U5sCSVHTLBPl9jOdCV9dWSZR8aZRcEGAprriuv
U3t5bf27C7cTIl4hAaKfwl525NL6jj3RuFkpdtcucsGlJYaOfcWVCp1a2t7wgTSk
KPh8omHbxM8Do5qAvyjEDvn4N9uKQBqYyj7UT8wUz6Y9T8qawAnli6kbs2HceRHz
AJ50FzbJlVheqtZ10c/ysFAqTfPES6s1P/mrks4RTjFYBwnWUrBgkRUr1sLyVNPr
uthH17NX0tcEAfzvavWTF6MO6uFlusnHDB36j4AojJceoRIWjZiusoUxQE8rftfb
Aak25kOZcOUpoojQWxZpDHLVwYrumRYw7Mb4QgpG+vZ6SVni3LNgej9eHBqddI4H
RL4jE8YOiaGKotxvEDCuf2apI38ByE6dGpWTmR3WtpuLhblIqMLeSmx1tzt5P1H+
bRaA/sgQ5fz4YUF4Dt4wSxAM4gMdiz+sC6TNX3uVxKA/C3kt38SFvZ8NJZY6B1Q8
ChTOEidExNJ2Yzhtabu4dKaB0ZnyBnTmWBIvi2hq8vwwN9Ma4gg0yIjzbzxELUVs
r9S5k81yOUYQknFdAV1/MLicJVe676ALZht1zm8jYvOUeJCt4hohY63eBF0RsXYC
fX3KqCFUEmhjO19boCzcyUmvKmDEhUXCE7hlhrypuzr6NYDEfJCmq2TXN3jSZPNv
+rx5jtXbc+9xruxmkxQqqNL/MwXh2t3flxJaDnKuoaFrgzXQ21hEOjnFyeb2wjVO
VqeasptQsWyTDlVnc5ImKat1JN9AuJafH2aKb/yoSo2RJV5FlD436/FYjC3beQ+3
k2zDCgDNie4v3dGxh1jk862z2N54x2KQx7ZvLEqDvHik2RykQafYnYBYCX7tLUAA
cuJZUH515PfTg/c2dp9rWXjPQ4WUcgrdWY1yiADBm/PbnDIe9U385gfj/OJpSiGs
9Bn4WBMureMwLuMFkCMmv9ez2nIJkj+1UIb60MwmwMUJrLwyPa7oQaGMP0KgnIm6
IG3A/lVBb50/iNOoE5LZv1SfIsMlmVadw/asrVBQX3i2sWeKRRPr/MJRhJ3BLSO/
gYasptSrW9uJVzJkBbnevatRGz1SrTVV4PgwSMjJSDu+xvoksDYBQwtNXJPvTlwA
KmiRWYZmqzGQdgPw3DyzdcK/9BdXVFol/f3qi538PIBweWSPnoRqN6RKR7BjtQlv
vE3ogWCz83WNvo7moV/ML7GSCCTPPyis6Ih060agthvffOOV8S3Pxl66RAIMKRgA
lD7zB/Sl0+Bic4RSsV+ZzmT6JfOXDHi2lIO1e+8R24XFoqyFYfF2nkoQ8bayyN1t
7mqTrs+xpa07Mjkt9EsvxCEiNqJ+wMAYOGGylB9R6YOEO8PPduO7GU8L8yqHHbJz
G5EOnE4NsvWt+48tVEfN2587ZGZC9jb0sIS8GyG4sHt1Z8kFQ9bJzSeR4cXh8XCl
5QKpM3UJr2JuSlONpfM8A7cSwQF5tCNCPTksVO9vbuHnV9++D3H6I8SK/HTfjUsY
Pt0QtSNQJnWpD7nOPPJOVld0n4+NOHQZ+3h/8sKUx4zgfUUi589Uc6pIz93+bSBb
Qe7gZjGKuCQlmjrTTrdaXsF6LYAS+uwkp8PLSkWE2643STUJPAtg3tApKvm+68n3
pHoAL0Y3YWFrn7ZsDPeV6jn77xXl9cw/iFPeI1O6vZTh7nACG/59PPZp4+44irBp
LwMrCECmW2ytp20Pqw8pGCpVAk308voFHK8Sn1uuSkhUyTbPWbLk2+QfimWPonez
svfm6wRpZijqmXacdvvS2oR5qN2sqlOblVs2nk2LJsLhLb5EPujmqPbYLkSmT8LC
BRZ3ORmASWq52GM0fYNiJpV5pXCmNbdWyj6K/4c6k5YZIkd7ZjwQ8gVgi8S75RKa
JnsrzoAj+FjLgdQBuJ5rS7VP6ZU0XOESDR0/1r3A9cFv9/c9s5qNmKXyrnw6r1Na
Iu01NGhbYhk+hEE8ChAYoxQYDm0Cudb344QT7mQks+FlR7Bm7OsdqHEbG9Vb9epz
YfTTZJm4gMORQwZaSRolPQtMi8ezEi66ASkSM2z3pouhWHl63UzW/jue+UNi7ZIm
jN/bfJ5mSird9AqynkZMnLTBPyzvFyb5fkFOn6z1JE9E8n4jr2ta7Oerk8GX7wOX
iI8i1lK4xymjxmS1IcKRRXUA6hRD1pILWHujn/1piZ9ThpciISAxDG4vGSgMmVa8
H8qk4RfKEXau7c8Vgo9z4mPs6Ho889qNuclW0gk3xRxehG/DQjeMyQSvjMwRcgIt
oipbSYvkMtij4timpQOK03ScRwwYybZ/Dr4BRpf0N6UEx9jIrqfRB1MptEidw4FC
ipLKFl97KaBkAFx9e+KLsuUUqGzDlgu46g4Rt4c1pDt2X8345crGDw5a/YLmLN4G
PvBWWnldY6yt54FfC3o6sM1dPLiydzpnuh7xjZ64X8mmTQCCX8a32Gih27VsYode
VpJghduQE67GJOKBLnQzG0x71GZMn4/JW+R4RLkQlIZMi6n4iNlIXIBytYS98jq3
CJWwqXitIoeOfeQM7djodFTUROf3bGkSKxuX5BbamFzT147uih0n7GbQzUmP2MTA
P8jKFHQj33Yfhn8sN9AP/J2DWxpKVg0oCe4H4PepF2cyoUAEqqkPqBUAjZ/kd5KU
Cr2vvzoX15AZNSws7pg8FGBHrKdR0jdFH2WZIpvTwxpxiFP9qjJv1TcS8HHMDwcJ
JccuwObZ1oZI0iaiKRJRIFYGgDnH3rMO7f0ZtlOaoLkLnU3ApXQIBte2iz4PSQLC
aEfxw8gETzciF84V+kB0XZjMjkcn4N+7WuVNPT4PbNLk1ixeLZyAV4q8Xibl2P9e
hlZt617x3juNfT4XwXcQbivFwdWHnm57rySl6O6Q2C38VT/dQpWP9OXzw6pnnHe4
9GHypClcuUrujYcFl702XC94vhaGTlf9UDf8Oax6UoFrKA4i9rxOnOGxGiApneKc
JKejQSrJ/2C/LNRxp8JyeKYckXIP+mXBSOB4BsyJcC+ATkwCV31TJujegUuk8yxJ
7HPIHI1zfhJDdt5HfviPG35L1tY3zm+AcxWF6yDOjwOQedfzz4XVqqANrZ+DldeD
vMxhGLam0EZfwszGd/Ht11Fk/Vd+O9SxJ+OJHXWlIiHm11NaDzfYnuYeTQaiH14s
UzR8OPteX7uc3EgkdNLrkshLSI7kMTR6uQvb+U3pe1u8njCM9TNqpD7ce4Ez1yRq
mEvOLaaSo/JV5AzStLyqbs88it5hDSgii2oF/7K0wAr3J8SUiwYCTj+m8a5DtnpK
IJlJUZj35YQb8jC1jdWBIEL3hT3GP36qcM2eIMIiM+ouchDlQr4vXrxQU/Tn08z4
WAgA0H47r5heuOQgHmBZ/XTDo8dwm0Uw4GMeRePuxA8T0WphUXhXbqTLkMmg4LTw
Pgnl3xmqTDHxBnGikcIdvAD8EfGsRraNu+5pUsk97IXhBnRFgyikf++t2lkI2Pxu
j33HWHvooH54MvTg25W1agX29ddSDT2KWjP3YJ8ZMEEnzT9dsmMi9uK5KitS2JdK
M9Ddkbs8UjaZX+OG1iUW0zvYNiqxdWGNbOsJmmnev4IB3nXcpjHmg30JM9id2yaq
UxKTGgiW3h3XsAQD6oByhs6fcPc1/xJY5ERgL4eUe0/yFrNjdQnfGimOVHxEpJFn
MrWBQd8hXV3N+juBKZd4HWsfrKC9fBaqf8CIoDluBqC3TIGEFXF7myc0IppSXMzF
ft3QQh2jchMvf9SfkXNpm+mRT9IjU4oYPIpmdpcKhSERnq5xF9BXOyGQNb4oxZ5H
OqCXijO2MbN8iObLaNkZ+QC5O1K6yQqUXdKbOgcmswSmCRXRPoH0CwHAqSL9+zzn
zXPJS48PQHlPZj3EgtyU12bND2jx0/6upk5tFo0NfbQqZLt+3W53i5vY48ELcbDv
A1hhzdPhjtIVpXXvTlokVFs+zk6X6MARNuM5CkTX6Tk7i+hAAe1r6XpJaFNVOvnH
NbaD/QoTa8ITK/Oe79DENu1o2s8VkkkwOxS7NqIDD+1dfLVKpdvoRZiD4q7DfxwG
O4A7Od/TMj1kQBPfuI1IEd/2sF6Ot8scgUO53BzEZiJMHsKee+TOUqX15Wil63hx
ga4matZ3voImHshcy2faKNM77ZaqnsCXXYDlGDGLMsaBiB5/Yia94Zj0dsfWDpV3
UhklQKJjlYigwCuCxhVdes6wKRN6nhfgM2qEc6sl/TT5GrOYI2SH9fFjDcrir1TU
i4DBMJnqMHuNYGzrt11w0Icg1aTP7eXI6Istx5DhEIrs92qfypIMsH3xrnfyZVLJ
a4Hl57/pCTPjnDffAXVsQ6+rzPEM4J8E8I6P05qZjT+r6ee5yOBJTWqyZXW6FPoa
OK7cTUp1PmbSFFWuG+fVMvmvKRptBeNd9iWnvyLxDYzRh+6wY4JAbT7XdH2I2uY0
+FRyQYw6JkLsYMoxrasxrvF+S+vXNSvRik587/WjV+AR6HwTV6kdY2NhIaPvB50T
KK1FhRbHgv/P9ogsLI3LXbiBDs6984uqIsQWaFLpg0N2Ko7vI5lV+vbWNJrtHfvR
+goy+OfCjgM9cS614PfGBp7KpGeei+h/Mr4GFG6ESLh+leyeQ3uZcZiguMOEOgWJ
aiudq3us0vpr/jd3ICbk9bPsbzWR6pLRyl9wlS0boSXOLKN03Zf8bvUinENFQ/bc
2xvptsXJerv5oz8GLR4fSo4HaStSAqNwSIsG2hf0qkcgooVKjFf0gNxJTaYeB6PY
FrV05xftw8F9m2tbeoBMABVwPodft53Fu/LL/fAMSD6i8X9FW2R11y01GYkWp//f
IHPF4kElDOhY1hmAZC02TR79ZmBIc/MwVjeAuQieVe9rzOpA5EzcKCN39Mno3r3P
Q29iWCa/VeALRxvYRXF8iCVnmv5Ot7UhPbhJ7JQ5yh64cqHogu1JbPGySJzcnnwi
Tihl+Y9vW+wh1UtXmG7m3PCGGw1pq0Nht3ubMeS5zMrcozS0IuHk3EifO+33/l2p
JOrN7yY08H3MLar+BBei5m2OspuP4Uof7IJxhwt9jFN37pZfCOH1+qrVhsqEbAh4
NaZJfg19lnDSGoJZ3/FQZnAIpqqe1WkpSuRIslGUT9cJY03SkTb3cZHp792+kDPO
09hW6lB8HLcsuElA1qvq3cyvjAwaJIiWmRH23ed+m1imj1qS3Y6rDoHlPFTdOzGW
lxAgyzRyBtIKHDijKlwUwQzPF7N+uP9OFvy2ftZrZSZPhzFLDOaIEgxGVRLBGyB/
KLIrVVYTq8OVHwVkOmVvDlIEo5ttzstLZ/EnixCpNWGR+0lMnBwLHSCNmZgHFW4+
9x/Dh9coxXyaWdlIxJXQ+wtok5K83pox8gEfWdk/YOq4U0WQFVRmnOc2ztsymowJ
NC/DygoLbLUY60Lgn5XeWJ1LthG6LzMA8wZb5otk3swxFQv9mUhuYu7tnj68vRWw
CYEuxS8tbYbBRf8olSigUytPo0asnt/GH04vbCF+TTw+6kZ7w36qXS7Dt1ZOojQ3
3VhqQ8k1b4Qm2nKTE2wezkB4zsI7vtLM62NqpVODndvbk6ltIk4/Tk8iz4KBP6NQ
1Pz66kC7wOcSaS64DIyqzqwaIze3y7a1sg78p/e4NUfNHfbTbEiQWn2p878Cmywa
2b8SoRvrFt9bSfFxAletqMTL245Wru7f+ze54mlBZyykCfhe+sUeC+MEunjTQ7SB
XDzLD86Vh3KcpxxkgsyGIH8aEm8bfw+p4LGDgrxqoZxfJkPA8Pc015fSY4LsaQcT
gOZ+Jac73EynhuXjCQKlkHJi030tzYYTiHNxtym9upanY7xiGk9PB2NnhF6CQOs3
BIHraUfescM5QrjXXD7NnwUJ6tykE7Vuu2+LFSA5QtzBRJ5zMNHVsSmgNk5E/NS1
EpNemCwO6dasnOmceG4aTjE9fl9khV9sUbAsSuqZt+DEYSGcyerVs+2xPP0htQgU
Jbs4wbOcCXuF0LS7tWRT7t3L47G0NDquvtAKHW9MGkEFhrmse1aQ0sg97bsw1cOK
2LiziEKsbQ30SYz/7P4XD+7B3UghK8ReROKgPvey9l7flEunM13Lnm7Fi4lD1Gnb
Mz3BNRO/w8vnUTlN8XMYi+cclHjo3ocNq7kGrq/cLWNl4wxuuY5yli1G6U3ZHN5R
/m90wLhWSBQTdpIsQpoquTNht/TBZmNHSDZNZIwLfbc3nY4iHCUItPiZZRZGflMR
W9AoJpffuLZP+wxZp+Ri2zSbOH0j2m8TAo5VOCkm5tvGNsdtirFceYyyxvW8LT3R
06/HebZWwld2uWhcbvfOu6L7zB4+YLljvTsdzUXa+bA2wxFQKoHhY76yBqfoc5Bu
xzFYMCXkRpblWeGZwGRQ1zfEoU3HGyEF2iGAWuVjW4eBYM/A71YK4r9ybK6gywvK
IID0zVfEL9R+7cftsPJ6rR5fFolVnTyAGRQfL+iE4xltuZYyXg1m+Ceqeo4zr2HQ
Bf18yhbwA02jsVrrhKL1kSo8YaxKuoCFI7L+fIh2CFO52xhRkrp3RDYanxqOy0uZ
DNGGEwrp9twTI8mJr/IGO1IpWHzaE57FVffyTbmQlxgL3Q6MyF7EhJYgQvKsvpcx
6n/i2ePBxVV6vdvfGxaVvcT/ti/yhl73MfeaLlQpmr/aBWpfGyhnmxbLZRki+GuZ
8vKBJR/8c7wREs0hmfFRHnMJMrvtk5Te5OHYoPQFT+BHpgngClOxBgLy/w13rQnk
jt5kES+bvShvlHO+xxBAq3K7Cv6B2UOaP7luQDx4yaOdZt2vipuPNZbVotQamcEF
f0Ntej54+FlU7mxG/yP3Q/cEOwuzlAZCdwAb+mZwpN257voCFcw37ZrazS1f3OTi
gVAy/it9VzJ5jK8Hy51CUqTSFSDwQGOfK7JoCbhhtrsHlQ0cx0jqSN830920+vZS
MOxuQi28bGFLKOQCQgZMweFMR5jAjNiXsCXD/aaXId7uStkINIrr72KLNXZXUNFW
Im7XHgY/i2Az83Nl9olJiC9oBzelRaovAn5kxBOk1LHUbc+F1D19QtZDWVf5bkcc
Q0/EoDlLZtzjf41zZjH/IYXbBprEWS0oNIeZxKQ+CTJeXRrNQXCjJEbWPQDG+P4I
S6SAA5DT5LBB/TcSUqaLQ0rMFFkFIiXU6opeK+LOyRr8SZBdDSnBscELzdEhdBNh
taLx4fi7D8TntaCAkERYOboS207rsLIqQAjbA5kRuUJzuYT1yoysdUpkFM5kCi6b
bzOyrSu3tcuXrET4P7ufEVuO+a615PIt7il2IHzmjDMT+sE0RyiSFHFtKyHk5xJZ
UyGA6bSEWwiR6atriHmGJJyV93x5eLQ806eLhLJBP+CIWGuq6jf5SJVG7XWhoCro
fqsZvDzhB6PoYpuqmw4GbrXkt9w8MR6DAVle0DeEkClTiv5CE54SfY9vAkIfNg7F
um281RoPMwdOOmVixEjKc7+Rr4R5PfDAgM8UctyD/lmOMyI4yC/ccPZ9ALFSxeTn
oqI/3N/MlEyZqRLw3RtJOhLkF6Qx0m0c6SmBqHj3mmH0E40CFQuFWI1mfshkt+te
pL9PmSRYxMmCPp/oHZAJToYbjtjH3QhGeSpLqo59CaO01lShOMuXF7mF3fSKgMs6
MngFrf9J9F/AjF6xaHVpT3/CCSjitwhGxm/UzY/xysXQ9HALRv7OWpio7DDhGoCa
DzBKgOm94jU0cxFubWnbkO079vQbSTclDAzE/qmqUOo4d9y3p12Y32dn4MHofLcH
ONvnR1SUgaERA0UO9skDPXZjmlZoh5/kpR7KBdy28tgEoOh8nhzJ2ln5Dj/NnpFM
BwYwVUX8cy79tDNLZMm96iNG5U5XbvSMruhiVHlhw944JwHqZ8u40Dxb29e08hwd
WOPNYlR8LK28o5ODvIT7lmpqSEh7c+qARGqYS99kwu0vZamcZZPvC0cuO+VpnUCi
G+GghRVEcxjmrXC3s9ryIIw55j98eByUosdpSjtE7O8jr+BZijbVcY0D++MT1x/F
RAI7S3UTo8PKISO231HBiZyPHQN4VthQ0LHEmmFo83WfLbbsr55D+GFvtmrHs0GP
sJvoN3AtDOW4XYCyE7/lDrK7CGEYyJYf7QwuKfSuMSS4u+3AJvjpGJqiMJWhMISh
8j8pGzHIxLUnxISRRzqkvmG1jNXIib8ecENzSbY+fUca8665KcDH2n9ci+Baod+L
lrGYdKmCNhRV5RvXYEq/eg+k2W0ttg7N8RahyF40f6WaD0q0Rck3R8dekvOiII1+
GajF7WleRfweyi5hJz0I5ROJYyF5+I+rDe2VXMdf7sPhSEqZk3avII3FQHVYfuLk
UQViE/m1CqU9MdYIo9XO+IoDTqqlTjaWTtXyuDs9RzxT1lRaVIzUHIFktwKtktM0
xtb4486My2RhvPEpYjEw7NG9jKiaTHNuIq6gRY5JeKeep7Gk3YTHvW+ZrXljrMXC
OKPQmKx2NJ20TVhYBhvm2vv1XvXUDxHwZfQi4vLWkO+4GNx4Q9y/LDd5YXcs4Wja
ndtBXUxvxfZam4HA5JtydW6wDjpyKAzHzaMNTBdjuIkH/nzbEB3QZVY6Gzszc6O4
N701CuV893JGW777QMeyrgyOpSaWBLfDumIYl/VqAYvPnF3bq0pDGbR7bbLv5loy
0y53k81rAzbi7QobYCSqF6C2/XvmAAf5FIqEh9NwIm6pBkrfatiL5D12V8deK1sz
UgyM/d8NN+paX31sVRYy+btaOqKn7pzmZYEynM1rDG0T6vUxCa2FHx5hDaViux7n
OJhGEtXalgBBEHCkre4YpickXirOIpi3KxaetUwgSfcBQjO0pG6Z3zNasIMIkoHD
wt4KtnNCNFWiG5Gk9iJ9v7OZ79iGZRhKqtLAVHA6NT/1JthFuMtUR8dkqZ8Dy+P1
s263vLyGmmwDMmN1w3PZ3e5QfRdBZXKq8C0Qt0QDcn0ma4PIwCuP4705SNEiUZQt
mopoKoJ8j1pj10FKMBhuk7IRmDo9AG9RFu6QffxXhW1rJ4mkr2dFw8S1eC5eQg3s
EV3dk5Vr/CYW1Nk2Am/guo3pBKvIGniSwebIk+h50qiQ0JL1ByeZEWdSDsvrmdPG
We0JvDa7+vHRpGvu4gt2KpHwk3LUjge4dYu2oyvqB6g2FZSCNrH/7J5Djrcztapm
7d65dxqoAfy+k6hIjIlGW4JU+7T6y3ycybRKPEBzTrPenbphr5NX2qgOU+mkS9cJ
ZdXJnt6Q6ZNZR+hkwKBoNfkCvvo8KidG+181h7d8jpFnU6l+KyZvvbsAUEcluZNZ
iq8GIGGU4cDCoYfwwQ4SBi/5U2nyAYjSDLHZi5TKIHvkmpkrZY0EA/qGf8sq8J7n
agtbFvWZuByQb7ArMEO9fGRIa20RqIv83nmsppj5r4yWpqcmP+azcJuYV1aWTlvz
1i+JT5M8AWfQd9by0zpRODhLbOc5j9PxzNP7qufOXMdSy7m7vHi5+YSyfS0oQy6p
MFXEyCdsr2rA4Q/0SjzanRc/YOKF/Ug/2baVSDfq1Efm3rdh/elyv0j+Bp3AJRwu
cjdvGWPpY+clhmMCU8zYARGFc/GD2quOjqDc7Uaawn1ULFTp3ecSD4sL3rJijuVC
nuM5kX/Vse8yvCRLdZxUeZlyij4UYJYRqanGg0wTmV77d701gV6Pk5D0yxe7cAqR
CleoTf/qcDcgAa7kw+wd/feuCCJ4WPY8LgPezI3Qv91t+i/q0mr8kBugVUjnKQo/
Lvc4seeU98dm6VC9uJ2902zv/zHRNATrdZYHAXsbXhryHPNd+srziKkBOnugyGoA
cvQUGUzfgCIpb9L6TGrXXb0sjkTRZ1FAy6yfzStbVejXEtrEPWvGYV1ukbsstejl
EzYFOyzvogugJ35vDJLrHXy6Epq7aVltZwV9D88WNbXmZAf0G7ru8Qo9bp3WMXLc
2rLd4l55YSHjNSE/Wqyi7PJN13hqV/PvifugC5H80S8pbse47IPDGUO/1MKaTZrU
gO8C71EO99b1pvsvG+XUaks8ZaSkuVqrgNAI95itAmtcg2LkUsSegMz0I6j68VEW
B5PwqeFtbEzhsFZkFwGiPUPOhit9d6iYW2nA5rzDXt4aVYl5X71XOROTJr8oYCsH
kzSX4m+s0rlwNjN6pe3bRoOA2oeL/R+VxKabP8CPjc28cbwJCtcK8zIDmGsQlCax
ONXYzYh/tK51na20hgEu7ID0BXQuc92gGQ6TaHLIoN8XUEnmO/VGdBnQzwZnuRpT
kso8IkAY0aUF4rxsYDv98EYN78/4FRBjfY6bKk8PLtp4phBwLtCsWDN1UKx0LgWC
/ACTxMHxjqOCV/al0kE9sUCUv1FAiZGMG2J7GzooseoTvyEyw3z9bdkco6qEhjmL
UwX9Arvp/LKxrFyCmhqCmLtsra9Pik7YbX+XvM3JHRG4MErftnvthct63Tt+/M6g
dcLuNGIeXFGn8cva/DeLgR9tTGodbIGIkmCwqHt7Fi/OoJKTtdovpS/bd4y5/4h6
AAkVLaDtalmvrrjKABKJW+VVX4+y3hNMALnRuGJoHlsTkh7utH6nMahw4Pfo9AfN
4MJzBweBKm7gvT3C9q7YQKhMF9XgcNxAoUG2M6rCZ0jHdMgxKE/fB97M7smUUCMp
+twNNWlQvOO1IG3QpEVxkTsNYOMArGX8Co7FW6fFItJkrZ0RI9KaEBcDr3HfyIcC
tVk9+7h3fD79Iechs7BZGAGRosIsHWi5VLq/LRtkC4R2BLq1V6qG/IDsWI9XA4V6
D3f/YiO8SekWT5vu5iPIf20AtXr/1cwiD8VpKizAOpq7HpO4EKkS0rAJsETRpynI
lpUE5XOEaBMllT8KwT5C2w9+LQ4p53SA56jJzXqroYfgD8kii20QAbEDlcFG+EOz
7OyGP9r5rtzuys1VtKSaXqSj7MojNg3KZAhOneLJFkOm7LOWhropSt4UN4GYpZ2f
9yEFMz3UBziIbTOh9T+FnA7zuvJZJbHw+5RhBzCkhzGt40WpjK1tSAY/Bvx6RJNS
I6wKsq1pzTPa8gye4s/m5Mr5XxzehK/MWwt0yEcQDHOmWjDQp1YeSWLXzygoilNz
sUKyNZ38byj/B+FccLAmC6bdxMROfVoTdffALVfYA4kUaknWsHJwJrvBJjBkPrew
BnWIdB42C3BjVqYKmYEiP16b6ivBa38nDBrS1vBkmrVSwG3rIK88o1q3x21afb9c
DnoU5RIxkVyCZ/AjUFdXI7IMU+PTMsVF9sQPlRro9tqhukf2bzOq6BEXoMkA5D2N
YpbUvfxWS+zgSmfaXr6DzX99+uYYcVou5SddLjgrJMHB34keBsyInd1otxKa9O2p
8uPk8QQqflUn7EYNOMkzZ7IOF5LjR4U/dnM2Tf9K2xWhocxIIEky7/t7HVR+RR6E
hdbcP5xP3+z/jaCIl2x9CwLQhPmQe0PR5KBNUxznUqXfXvnt2shE3xQ8mZ7XUvDv
H6urS/Mq01uHaKPM+OzAbkTJcxEv6l2QCSyAwbEIn8239y/i1BFenc08c/4mDZGQ
/g6QbZsoVhMdxcY9nNY2FBb8DO+xtHZk58cM+LEj2MhvNGtH71TvA0ghnYXBkrrL
7Mr8RKFFbhln7vA17wRyD4JEAKOfRaBUwluZ9IxtbxAZKzp6CxSE00qD1ai9agvK
t32YXjIx/GHc/2XNkMw5Fi2anSnu5Kq502T1Oim/f/sIuMOw42lvt/4RoT7NQC8v
sIH/VoTAhtE0cQ/S8ESpIji7Lb/fR6+ECInttb6qgL/c1AKWil3CS60zGSD1i9Pm
SKtJ1BTY3JSs6h/s5JV9202294QmpyQKLDJUBxJLUFRJN0bS1pxs0btBdpMRriPQ
IBU7jJ5qK39GybUfyzmwTKpj7gCHVUWFh7mI2upxYyTk3Gr0YDnWOjSEtTAcTUXM
x2wYbdy5zLjvz0dsQYmJAVSfyZPg+p7KyFCeJ8MrVeLKc+y5JmeoSlR/vjriSCXe
T1cpU4zMLzUeeQfDYlAALRYc+SwbKkgeP8cLLj754R1vI4LfEHan5AeMuKN5ENL0
JrzQA5tdvWq1hWg+nNvAiK6GpSBVr2a6Bd/qsyKReSG6+Ouu0jg4CFS/75bK97FK
m2KRgaGBPqAt1cM8KaLo7bL5VrOULYThMKay8vZyYAnf4PVkr+MaJm1VgzezT4VO
XmeO/ZXGbY39H6LwpvMh4D56noPD8JNkxS8eRdGG0d+nJBL+K4AslKrS832hU4xA
hvqObTs0uWxDbtyr9Bb0W2cp0VyxTieFIr86C5Xw8rsQH0+V7qttOY7wxe5ue1aL
mjPIX0UNQA423ps8rb7no8/6NThIhbRsoJ/g8oFFeWkN85T3ED13FCx2Ty9Dp3KG
34/ADgKTHTZIl0o5cw6uAFdRWloWdYb1wh8ayasPNUfRAJIDTqVXUxEzxvuqeYnJ
ND0n++IXz3+Jx1XIaJwd+K0f7OD2KoyFsBioPWgWvx8CXFIsy+qYTTcT5FHyD7h8
VJ63MItgF8XHBt5gbjFRNi1+99j9NBV5oT1jXfAxJUS/bgaY0XwlocLEfG/Zftnq
kJs6CzavDQckARPFtroQ6MUBHYbnR9zfqs3usBTR8zKpbFK07E/ucZvQm5HuDbuJ
9Shk5KvjkkejwnVtYVegXpCc7ydZBm9nuBINHZtHGWZXoirv0BtHPjPF03a7hK53
77H/SDNbl2YosnmAn/wsLXhMd2QELftsVOXtpC7OLykm3I/KY7vWxP99LgKFwFZz
aFk2rZBwLhlJtqsNPcfRkO3Ayi33KTlgymgf9tjZZxZvurV+ZkfLBYmpJUEIxP8t
mtEUi+M4jKSD/kYkGeMZbXwtUiTLqNkSQRrLrqzlh57jE8BSEIlt2nB/d5aHdJAA
LBC2Ediz9ysr4rCRAUlHbFSU9Qxp3GzwJi0aea4C1jFmTwUcG5yOBXgWHjCeEVaJ
LT5Ons7JDGPhPoX/ep/aVhKbg3h1K+r8yLixen2hiMZL77oEVc/HVRRnh8MgegFs
g9EsiuFzNJXgWIQaSG4V6mpGeOyxZuWmR8oIYa1HPQ/KFQhD2e9CxPa912v0KYE8
yEFOdtJTqpqb/2QmtjsBeyjj9xMaiUCChb/xx6lz8uIFsV2Htqeb6GJREAuIEQkT
yWg2xnNJnPKMD73JYcWtuYG4G3Hu9YjxkkCd8Sss1HOXoqIzINdE3q+wVdt6YQ5P
bvhAyOAGyPYj1ef/cHaBST4gJBeuVPuw4wv5ienjv8sLc4gEvVynbT6BjevONrvX
5aXUaESVYFdb0oUCntnEt35XI3wPvoyu8IxAO881Vtj/bzR53lMTMAMGpUDpeZVz
9yTJvjadqHVx4IL+KWekUXfyP4ybzFjNcLu+dhgsXoW2OI2fEzgvxmD+85IK9BYf
gogzam1wG4SZ92YXsp5mlSAbV4opZoLJjbi1smx/M9eyS5IWiRFLWxfHflIjphBv
1PAFB4mSc5B5s8SFmtulVzwt3faSW+syGR2fD8VzWvn1zvuUWj3oPkLR38IdKmQe
lG0KHteNQY1NCvxMV9vKNcSUjw3RtRSXwcdldBom2IbP7A07iqNH1EH6UmydhOWC
Nsrn7NC2p95sjwCOUHc1p6n+L2nmMfmdLPaRpZMmkKV7gwdCPNimOyzq1E1UEKHG
XtFRa577tn2hTOkb4XgXSTHOTiTizPxyfjJeDdAvVG5EVISw2ocEH92HFEbXbqLI
9z/LNOmbsPn5RuAFSP7SCd3k2W64hFbHfOke+yoVMYKM+sZOGAXaGgu1Ca4OcV4X
BZIJ7U3722xoaGcLc8ZnDMRjlDDIsJ+maZWB7CAQl0FL32BGT3yCcdVyto/Z44J3
4TdKLBCZJwzGD4uZD4h0lvV9zRCHAr4FE4UmH3EL4QJjT2FWJIwsBKAdZlpoFnaa
rKjIqKSLFQytziFViJKwvrdv1G80fAy0gxgm8FtTxp0JbLCe4bfYdMEb9wh1/qfo
HoEZTzlPtUzT/XCewwYnQvlO0FuHPXSNHt9bR88aozHLIVjzPBi9+h2TfutFRGuh
1zIMHaeVBJFYTHWokoydxEMij6oFAKxo7rDtiHrC+H+aeopB6Ze2Y0gud+sxMTPs
JHtzsJWAxCvYfxt5pnGWr1KTylRDrncRR5j3eflgVt46Inqx16R2VVIy1s/nT7pZ
wAlKpdzQq50GY2tN2aA5AWm0bcZfBcCH6zWnUaLQK2kgn3ZLQe5m5JRJeNixTBm2
eDQdgcDgA9zK8DytUvmUrrYmPfnEWP1XTUDgUcqsXJQEQiF54nSUgf6trQGWwbC5
QJPNrpJ8iXKy+lA2CKWvQqkeaeW8RwLkzlN0smRQTDqzDswJiJ9XsQ0E7cOFjgu7
iVP6bRwgGLWhYK/hwhWHcCX77/U+cY7EGCikdX9T86P3HbNo62xgpNbP5dgCD9bo
xb7RJmOyzMWGdBo60RTTQ8mXGBPQgUrt8p6GzU0CeOr57XLwTXeP0a2wd+ue38a2
X7B6QKIZxpLwfmK8o8nCas++2k5hP4d4BQFG/Qye0dS5G6V9aq3hTkq+7JeXDNv9
ryf8EDRHBp9kp+ezDcO8brPRltzN7FrWmd0CYaGOgjf/Cb+VxGmPZJe44ovMOeQS
3zj3EDngPFnDybetp7kz97K7aThp4e5CAv5Rc0JRh2SvkWeYAy/Vs2+RmdKAstXX
lv9vaIflBKVElBO4vFv2TcWLveXf4c6DtzeZryeCs/JN68bfQ1FeCh1IMs6itRHu
heieWeIU26Svt1Moa51MHxAX7xEKrRyU08vsjCqJDHuQp3MxRkfEtFs5Rg5rZIYZ
+FguaUvF8qmH2OZBVv4f3ht72M03BBVQqAwxX9lvaOpiYlL8Axx3vYnWVLlN7t9/
XSZhdM+in3K+Css34rFCc0ROz9J3C6QfTF5E5lOZs6iND3kDQ6ZPY4HwiwBbRfy0
aKe+TQcRcYgbPupjsF5Xr+IUOrw+9MCmDlAcE6jlXwY6zu4BEuZtQ8MoDdGdT3q4
fdZtRvDKgCy94VR+ZFNrmhZbHBbdJ3d7sY6hYh7nEOA9PxiRHzrE4+495sBxypBY
IhXuIhpyRaZyXC95XKkyK+7VCm7yYlJkj2rbNfR1j+NZIDkaAdIjAA0zi7h+vKhE
079Ko2K7/eGVa9H7JiZFScAV35aaU5+tz7FZDqRFHkGH+qP1Jkelt1VNkSSoUqvF
O7jFPBJJGZXq+gLDlMODKdyohpgoy7QV486PmB8FbAcnU0BZHPAChRDVHeKOKgKm
ww6kwjx+womk3B3uDagpg3E6Vjo2nluOA0pKezniatSfGDcAfjEElrXthMNIHtmf
i91DxtEdlgE6KSdO92SLEQt2SpSsXerJIdBC9b2W9HV2yXKc/wp5uV5cjs5RHdeS
bxtjxGIRlcFMfXkImtZWP71pQ4klOD8OAMwq5lbCUObauUtiiozFB8iaSaHmyp/o
+mHrChtoZF9Fc9XxHdlM3sk/IMUldjn8KmlZY7qHDYy4sR1biI1ozWfTvSI+qYE5
xrOTvi6tfz8R4p3cZk9mLGIy2QKSAuQ4a/O5rg7FaYACdHU0Mldf/T0BgAJHBNy5
YwFChoqwFg98I6aUINjQ9b06z/2xcIGyEwqP/goZF7K2rJ4ThR14yBM2LWcJP/9R
dfcfAhQCdnUk4AAcipmSHd1oslLJStUlj78qMu9jM+a9zM/yNjVtYbWyDp3FEE5v
IciiAlyuVTPpxVX3pPM4CplEq43Ex0L0QczwQp6FFEbznBOz2O5ZZd36GY//lSS6
nS4Y02ysTqAj//2+kfZM+bdcYWWqkN6cUscSX4qaqElNE6f5nv+MjIfMgVWNXSKP
ZOe/hBoZ07Wm1/WJsQAEc+S/3iJqQ4+mC1fnlUwBoQWv9ir/M35snW921Sh+f73Y
KKRftcmqRnniliLwNWwjLdU/8pdfvTs7fZ6OnfESHQ2IT0yXosSVdmsq/6LsRpw6
H95fRz7bF3az3n1Rwo4ob+mb3yqywx1jO2AEGlZLos4u2ptXCA1c7yb2UtB1pFFP
RXcoLQlTPqa3PmFDNq58VXptCxIjokPoB1ldXhlsm4OoSMs8utc1HOvZtg7vHxQm
sWbculcF18mU3iVE0yBibqMTHEdMqk/yQY6RqfWr4231QlHvuKSHyOMgR8p+8+wi
MvriFiqlAt/5cRHK3LaaTwyJKK6NGLYAN884XD2Q0oh+8G5GkQyx1J98qdMqZjKl
/XDEd96FT7WeopXnSaDf0UYvBNgKc1Rx4DOqPhEpIMbgbGfULSH+82+fAgg7vLMj
67OGgH+BB4okuOZ4GoVlmbzVKHJPtxin0OHP967UXH5WaLkOiX3TrDtvdwyhN0cx
Eq/CE2deoaZ+nknFUWgoICrOIcr+BqOLCO+CSf+KXVW1eAlv7ywpX9VHdiyi/yua
Rs4/HlJi9lEhIhP3Ghn2g7nE128qimZy+sWVk8p/Uf7G+8WyFhGBz3yeYjLpuWNO
LwtBOioZfFxoI3UHgjGfZ0mm75aT7sGCvKWmoZCPW2xKwnmkaVK5hXYF06agodVk
yHA7M3wGinNP6AqQDhzoxOOMSWGGtxbtP4hl72v9NzCjYz6b0eam6qNesZ9N7FU5
Iz7i6cuHySV80sil2MSU6rfBa4nns9p3t3sNdKQNBijn9yBlcdgrbW4EYaN4EBBT
eksk5ruaZSWuhLnQpmIan1d3mpMbUrI3QRq4l5RADaXq7zFhDUIykuOXes5yJE3R
tkCTbWF3/dnfWBg0H88RPXAD/BDWE06W8ejVDe/RW80NjTOer5QEFiDovDthy+dT
hT4g/13Gs4SbheUP0MnKUCiuv9EJlPe2Eyg7g4zR09JVtInB4dY6w2mAgQK2Pt8Z
FFZKDyd1ZJbGIaqxphlbCujboLdHSf50hMtKkXNPUhOwdNhM7BAhxbkHicxHuFlQ
N+f9NWB95budHmZy3rHQ/lziis/Jr/vayCLwYXtiD7hQx90Vmh0YaJ1UWKqYJL0n
Ca3dHFOTHotZX2pt1R3lCMdT0mawBrDfyXAloyKFwHYsCMWU+BaW88l6G5ZOrhZf
UZDALfg4fwMbuGJmlIhJ248+XD1Xy/M1IGAOQZOpVDoRF/rYz7tlk5xenwYS9HmT
sy0lqt+6yo02C2n2Ml2wtjUGLx4d2opQsiVDXWIKgJS+8+c341V+TGBsCzZcbmai
uiUl+D3n/tX/qBNe5T5zdy8reVXJsMR0IRJSxXz0WiCPvTmhVdki6B8fPt6E9vOL
iE9zy/mjaXaxGqoEAg5jYWZHAZfJD6+AEVpWIh5y+5k2hsSlQLOthc1q0fbVZPGw
svbnHTuTNhvn8ZzhkmGhmt2Ye73RXQCX06n+5sDXSoCAc5cWJTafMaoa6sIKthtU
e4EPDlrfVedRftkl3SnWpNiVEarQvTY8rCeMrfY5tnA1G12yfitegPnuY3YD0AWM
CwbEvnRZPJm/AB4koDM0sloXNyf8nxViIANiXKlNZgNhhMfCkVDak2Ppqb7kq00A
BcGPmu1JAi3yJWO7nrhx9/1LOhDc7oz8X7HOeNASTvaw04I25k0rAcpSVkgYu/3s
ZS4Gss4bFdSonwHzMrPidmajTbOY1NHZNxR1LAR/+Q178gPXDTKI8nVsO0fqD5iO
S3xWSwUGRZwvWXgEzr8n3ZuBJzLgtu6jp5RETo0Vu9/mxSOSJSaOq736GlnVzQ5S
biqN2PxeKdp3l5tPPeOsLQCvQZqh9swsgaze6QPa4XFAuq/3C6K64YHCl5vHkMZx
BrqpD7VxuDDyFau585XS93NvjyvY3+rigkRoTd6z1U7EOEv5nTSMUhz53r+aFpte
wh4cfi7op3U1d+T9YbTTLhmsl4N9gg1an6HMTga1fG+25Cu7WnHF257gogZ019zl
SPROMNSSZPVtWhXackUFMfpMJE37GzsxXSvvPocrBbb2L1+q/squFGTv0gjypIai
NJSpZF/Y6dDlYGCIFNYRFIliXODLbnPr1ZpEjI9ctt6V7as7r1EVDYDCjz4cDs8Q
ElTAbHkxWZ0C6QoWzjehffw7GIOIMcVt0RAUghJnj09weXlfSzq1xl9xnDQtwDMl
ZMJsQhTjB/h45Dx+NfU5htmP8mdMfW13qft+uH/VfMqpr100lw2TwqJ0YQFzHrdz
TtrUaop+m6QEcd8HCAuQYz7wEmVf58sgZp8eyGsmy1XuOsdF5cFdFEdSFY3cHwhb
cxJqlqSsHQOqXY/hV4RFCJ+ld/KXINylh0gqOjYZTHpyCOiJsrGUSiB0vfE+khjO
DF1UOcE7S2HI1Uuh89c6GXv+Dx03WA+oxGxoqEg8fms5SDrb7oXw9N+CWrPDedWT
cPy1keYHbOdDGK1TZx2Z8lQRo1FxeE+/k1DTbCFPPkqkRPmqyz5U3zXw72dahiol
T48EWl520lBkieCBS00s77HtpQdT+p9+Cf0CNJ2NAeyePQIHnNo7WJpZ82wmc6g1
WKSyao411e/0cxHrMtFdF09+g83ipmnvLO/u5ZbqaZYKeJFRdvOtsKcp5dgMTISA
o9TW31oxAGZz9aSV2hg5Q6mbepS9JSeXW4TL8hgoZDPX3U1CguWQDWrKKhy5hTKA
whRa+XUkZA4H9UG835eNzfZHKlWEOehJITfZibFCpfpzhS08NTIk6YuO8O5FZ4Y1
T3SHxuY+HcFcpxhzeQWIIFvz/4I2RxFLowMcf44SEz/5gGbtIjlFz3DGIW+VKbHl
LOURF49tlJmxyc/4daIhN4MjN5EvWqPQj+2ylbdZjdji6IhZL4MfVnRtdnDBrnGr
TDPINww44ae2aH+0gJr36ukoR5AKl1Pox4xUePgqZI7Yz4XOPY2AbBoJNUVQstLO
PXruPmIz5qE1ZSCZlEstwROmpa75hcowQt9WRUqsnxS1RPk+1DtiOsylyq0th21x
zOkrm1QcT7rsrWr/c0TU4rPVRO3K9NOIQl/Y0eroX+0SwbE4avGGi5aiLtu2lOfN
3DTdyMff1w1NKUqpxFAcKaBcJizYYUtPI323mniu+pWny4mlWaxrzH1gZS7SqGqq
tvpaVwL03eDW1pY8iM9RJeUNQiswfC5FYaXeiqUrRiTVlcCr14Clham2KGVaB9hy
awj+/KKjwIBIu4ZdLAZ8e44ZD33B2i9jCxI4OP/x09Kpg7s84wdiTlWspwHMOlUy
CX8xaT0F8IpKDbVCfdbZy8M53pyxttP5XRWd2Q0wMH9zmbQwvsfe3bmHbCgZwa5M
xLdt2yaDY0EhohbV2BOAQ9GNvArCxfl758Eu1w/6ChWhR+nkBQuX7yQF1iijzKe4
OcBksAw5XLSPv1oWwFUcJSeYSMnXBTS2e7VEgOwH3ciWCVK5no0o5fgIWrjLiXVh
PXfScUi7kLzHZETi33DID2ON+hHvLmdpbXQSdRvPZ8i8642P+m7geBUYpolaXW5K
LSs+uRZshfU6LKkVGToM338sWmTPJQ3aK+g+uAoFSW4cf4YfiHroC5ClwvPsbMPV
e0sQRkACOAyqwARw2u4PZNCfX8lC3EbhHDg2XbFSlt0EKh+kwtXeMhYYJQkPaJvZ
S07Ekum5nVs+pSt0Y9ZvyP8Sr+6ZI2aKWw4xTBqpbt5Tg1NuLKC0ezCl0CvCVta4
M6DHoTtPjVl5TMq3nO/pYBK7/UbivI48Fc1LWl5Wa1Nq4+i4HSUSx5swJnK4SoRL
iJ4R4wpZw2qg8cDjXNcqM0cS/Yq101XhxGDKpW1YFcDZp3b+JpI2dACQopUPVZ/m
uP0nadwqB47mdIWPag7fcMaAc9iEF13SiysMgGIZjeJrKPbK9XdCmGDnh1r95KB2
ltmWG53mH6RIKqB/m91xFEMNTj3dkGgRh3KaVO8xnB30Rbs/F/dyfPH0IM50UfYm
EcL+ObkJSUclAGcWpcWj5l6EmKvKPAnD0FFMdusu+mDRHYAhulI8w6+F0V89vIhw
2ewbbBNnMdBOJrwCdX02nyn13+CbpoyGcAxQAkR789Nrs5RywasC2efWNcxSuVTC
prOSe9nxgFCzhuUobU65OL4YmCnO0matpyt/EFbDNIursl+ZBYVyh7JGFjgx9efk
DazSMqoz9j5Lo1XPTCfp5WM4BAaMxydlOscNq1WkrQJ22KHF8Rb57nes+ciWQIT4
x9b0Xlp/iXydwQco4DXBbzpmK1wXFep90pf+ap0oO1vPC6qwuG7+0H4L0V0iNrSy
1rwO4LCDNIAOL8JRDp9jgWgXmNh4uX6Xru2cM0G71qwdVQfgBHcwCUzSBrNMbfjT
XH42nQwOD9bjmLW4sA9qFwxD9ht04Aq6DzAdMRbJ9Cb5GmMGMTCjdP80vcYq9vbb
LH2V+OPxQTgAYEHyZ2rbyAmYWyzcGpSkVAGypYm3cogiUd/DyfsZ5+Vk8bRg/3nM
r9ywSgtgDftBuEJDBnU0NpSkvUQ55lEDGw/AAchFnj6vmVe7JXy+yjAxyhvsuZxd
Dz9mt2HkfMGTB9mg2lDvC9GOc2nkHt3ZXm9Pqe1BpUQka7RBaUueWGcxd8PkqSPK
vZZQPfUvWUSA2VvDPTDH3SVLPzNPxmzgX/GdLOnJHdZpOn/3g78wAxQ0s6ZMQ0Es
DMLwilJZ+1APiM4vJmhG0y+m5r1wBuhY9HrQjggO5gh8c5oWOzB7lQVnlQWuJcKy
hFoiPl4KV9GvhT2fOmcGyg2yTKmg3O3cqt+9+Hh/zzifDo/7yv7NjO5VxmJdKR2L
OO+3JhseKmw8eGvt79v5EsMnWqGpDq04avo07W9JhQAzKxqklP2EI0vrlo87rwZ7
tKzUgBpVxlSLaf5/lE+M9FyHqINl+U9bkSfoZMA830p9t7hyGP8jq2sRTIhQKdw2
u7GEuz7ezZnpEOac6IvBd9JnFM3Fk9rHYz9im7sJK4PeeJfsJKrEHzsePaOE1k+5
ywk6LmtyBhZVtTbOuiZaeifzsGJITugDZfcU8Cv+VTefkS/L54NLcRdkahdIW29Z
HRTqm5LRNet2r5oMGjEsI+VJc7/4EcsZ0DtPdRUIrqsS/7qGI/MKAyqleAW6qCyR
HdKWYxK5t7g8dYGP/Sd3+4XWqxhH8c1GusosMv8mYXBYnHuWacqgf8+Xns2ExFBf
2XF4nAfRCq8UN8LIh//iHv/j4npg4COx5Mc9k86sqgJLSFsHh6kLfvOAgvANfj8d
pRQ1QB91varSV7eUoANOiJngF828Gv9RUrSAsAji/9KSdCGz9A9WvxC48q3MzsEU
X28AaKopR1Wal5NJv8vANlLUavlrzsrpqAr1Dlfzy/IBsy7GATunpHTAhMs2Rea8
PeHZC0aqHKzOZ/BpLabHo6ACoWkbo4VkWee/bpFSIeorNBKCgHdTHhU40cu4CaE8
/Dv+euQR/gaav4yLpEd4kmBgNoYLEUXZ2NEWhqcQVBHNxHho3InV/KAHJmzpDVl5
MkIdelNme0HLBZf7t3ZVKpQmkw8uuTx9+iI6jhn2LBCTlsOFKrma2M43lE05Z1uW
irjni2pESqgkTUAPv0I3aODSiv1NLFjiTo/WSMhT7dYVRKI11gMt0C3OCRCKGFqI
RttguWtTwRQiA/6xEGfsn08LYdmGcZGYGDn/VmY0zqlINwc9iNqArtjP0j8cybts
OyHts6Nl0V+6xwehEnAAXJTnOGzagyEKexVRrjcxSZ9LSkAlOV+ZT5/79iDYRSUR
x5FlxtMSniVACdarDkVsJ63MYRL4Mol11I2KcxXSxZSx+DukvYGj2pKxXpasn5Vp
Zdg7/RKDXzETMKaeWO+g6aCjVsZFk0h0fAAfuhJyakCbbORS4GwB8wNDlR4nazJC
np7a/sq0SDy1XspiyhQKzgbXEQEJ5dAQuiz/+krIFKc5MabYEexlBqcEomjC44Qg
58pqFIAa5enDGLp3Ci8QRT7VhPNcbhHWu7MiNAfVyrK8GZ15pKjmtmcMQ211sdeE
2U/Cw/1WPtE4LyVbJ2sCHVl9AHdC56XgLhVrMllqBR/MyL4hvuo96Dl3tiwB3fjN
OaueqfKRfCDv1Zeivi+CVTa/j4Bdxajvou54F0KHbQLTqAdvXTDtZHX73OMPZDeL
IKKkaRgxIsovNbmxwjxjCee/hnEeVppEF8gwE3fd352msx4S2Sy7XQKO6gq0TPNz
FLIdaPmKJEr+gCl3G5rgl6e15YWZRNwMXiQRKjnhUsHnUSgIWgzYhPeBTnYaayrZ
e6cmK6doeYHohY/L+XlF1BsIoIFK7hD8isPfML64WkUrXl2z4RQ3qGspE/wN8IGz
zrAO9ed+D4+2NZ96r3y10zpLIjhdLrMETyojMHk9+2aMspb/keaYMLnomt2+6/9G
OjorbZG3eAdUztVaNG7YcYcU99UhMi0nem4VLLc8mKurGcAvuVuMuaCuKRprOMGr
iwuRf3QPgZeAH0A1GgHG3PfOwzgigCPn2rMMDrNjDm3eBvAHRAAAt3sUhoZFVnl1
5/GTsZDv0KlmaLzqCZEU4Qa370n91+qacDEkmxCA0JXU3Cxxp9XrAhePDFhqiTi5
cCaIlGRuxoF85pOO5ow1gDtOY4vJb3qumb6Np5JwqVNsMKU2ur/6bw+c5DMEtFUx
QxWmJOz0OzKMxNYPpyp+d/YZ0fuKwVh3rpSOpSZgRHhG3XbORUjsBpm3XRRmDvpB
Dc5Fkrkxfyxmrp6VTyM5rj9x5FxjDMIETQSczSIpttjoPua9wDTR+D5g4uVv0yQs
IdsVUCu5ANxS9qJwF5e6axZbeymMIdyH2qJKnpYQYXagK+7zk+o8FRsPc5jSmHPb
2JrhUU4QsKVeyltliU4H4ZGvwlKjXA5iw9jfZHu8imSmzJVaH4TvX2arxO8/3/aD
wI4YGxaQal4c4tqPWqh31+NW+dUo89ZecT2rYhvBmH8ztZA3TOgwxON/+ysWaNfG
vtnmysM8y4eEwxNl+KDmUxQpGAANDISvm43/SwQMyEutGCZJ/oxn6A/UFSbjsCb1
Zl26zSa6S8yiCReAIhlr3OSTnfDcXfPyARLD+quqe5BeXPdAgKsDBkgVZmRdb+jw
ItHH6vwW8FHbLpIHfy+9f58aPV7Xhp8k5zBPu3yilH9cA+cWe+lXEShAsow+3NWr
6YTBpB9L+wn5HgMssgo/0IKic+SSMa4v95BSks01taKKYfuP5oM1LUmaECvmveqw
zZ9xF9HTcKXhQoBifmcm6KmrweLVu/I36ujnuNc29vxaCWzRM1vHEJwHJ8sj8ftL
358xOFstG2qyJZMvBJtUPm1Td0pp+u0y/EeOEaU9hvCKPNTjNbEWubFRQ4FHGj/7
4h5ZXKeizJNCDm9MuMLR9Hh7pmd2T68LzDTobiAHf1m8bc3c50m9iZrD1hIiHDZn
ye0ydBxpqhq3GupklUH6VFuGq+UT0nRVThLiKEqActlM36FMdWY2fTHpCucm4mBB
sO8AKRg7WztDEPKyGkggVc0HA3WxyB+WS1lHUDcDb1Q7ofy3PZEf2qFlemeoR3lM
8X+h4gzWcdsIBLOMLRxwpV4gKRIwdPhQx7Y/wgluPXuYPvihnnUUjLTuSTp0PBWM
/WS5DLyaA7R9yfF6DSpGas+yry/+Uqs6K1xTwkLaMC42IVQOVZo1O8LdnaFW1bsd
ewajH1U5xu0iiEgSfSF2Yk16IvYymany7LqZ3W3cKTitY0HEVL9rU6QSn2UULxMx
OeVs3T069YH0w2L0XKAZFgiBaze//M4v+Ed2yI7wHMgzS6IY8zP9ROrPUyxe8kEK
10g0Cx0J8CX+qCKjt4odVHnKQjXhduP39G9Dz+QXLKv8GKr4a+1RCwzGlZoCEOoT
Bdw69+EcWoj7oWvhdUCMjhcz063shiVc6Xj/BsNSpR4rESHwCC3uR5CEiUChqI8S
MDqNTv94RTftuQG4PmmvHPZfIsqilvunmTGMFLvuXH33MA/h7aw4xgq1v3bYdyTJ
F0Ht/PqUlZHCxnysXOikJlXwtxss9UNFfNxXZOc6QWSCX5L+KlEzMmOmn1Y57yxF
DmyUtEH5bigsd3kjyxMs2qpJJ0a9ydo+Fudqlve1TTlnkxESwyMkQK26zfZEQ/gZ
99iM932pw0NwtI4Ad6qJ/uZ9XGMpI8nN0qAkBfQrLvy+ZmyIGitHQxoTcxVWnw6E
+N+iYMi15wE2NDNWXrhCu9JrRkvvd1yYwBvIXv2eM0Qegojt3hnK7hbJto1FYI31
lm1qO9NLudq2KeLlLPYNXn+fIAiCbKVp9w31Fi6RaRnUfNHQkOSlmECHL2sglAA3
wpRmSCeczNWyWo2MQDWI93XzOBDLZez4kaWIYRs1VrYZjZ+v1nFNvZRbjxka4htY
uTsl73FjRBVre9p+EnKXIgfcSd69Q/wYkMi4mrisF+fAMm2DNj0O+zWYwmRjbt/D
dqmpsNbGhLNDAfK4duYR06Zri8phZOYdwMA2Z6RumHarGXhoy1zJNuQH+HuFrFGH
8FH6Q/MQYx/ZZ710sROUKvOCa2w6L1cuKuAvDBjgdJeJ8xuFAMHGicO2UZP3K132
7AFWkdrFrUbPgcROgsDMdR6+pGv17EsJYOZ8YpHxCCGyWiYLnXL2PjxA6RlGNNn0
oA/tigLV2pzcnkMBN7qBP0/HD0DW/VQTJxc+q91dCi4kyKPNUz63N9XS9787GBJM
Rsmot/ap0fA6ZI1A28aKXWNtG+mdcJO3gnbKRbdWfvR3pyvuK2YgcI9VssOgbvp1
IearrRnCLvgX2wOx0drwhWgLWnQZjc9Wbc/M/lm4elT/ofpZP2UiupEIMwgJdRvY
rzxM/4gezQIH76bEWGCYzkxWEvKFINLki0byJsEtacuxQaRbHChLFnOSYth7IeFW
/g92rLhEgAhp5igsdatfG0rdkj3zxU2aD8IzEcWvaVnRI7Cr7sB7iY7HGjyOEOS1
oZuZDJ55Olk+7RviKacHBwaDWXLbStVCc0sNvjB+4XsY5r5QsJ/c6EXq/Qqfskrn
gWYRWZyfNwI1OdnDPqjyj/TgX4BCs29g4+v2kKaaE5Qp9aCwxQubxDCVn4lwOBmH
/aWJrtaJoZLeN5d7bA+xLrBiQsEv/yOOG1OpMFkPMN6lkjb+Br5z+1gOH6ZnajR+
WWYGg3RXL67HBxMYkzPMcicKaiRhu+1mHb5nAVghzd64VuEDJnVmcf7D1YWs62c/
blP6M9mwyjyXrfCaFrbREw9OXTKkXAXQZHjQJ02DD6H0Ei40J8jyytwRLSN7uEig
sMcuS9FUPRo12oma2zt2JaJfA00El3qpMzmMNYg71RjKPUOU9Qd6HR0gj6LN3GEn
6NXhU2hvy1wLYjDhfhpEdLQgJY34m2Bnchl59qVRZVAHYPAvbbQnmEJCF19gRyFZ
U9beoJ9SA/v+dYrWuDwu08HMgdkyDRDohFcXwrrtphtJ0sz3mRFDpIlF4Ulw686H
xP4DYE/TAQcghSSCUcBO47n8MQhvIuotkAIL2MhHI1/cHTQVmOVzb6hQ/xaAyeng
qlSp7qImtsbumbviVl532qHpMegCljPR8fGiZ/IaYfqPh+LsIrhjQsmbI3PdleLn
aFXjkO+aUa0p3+Abc+1A1a2gUkfOhZhZv8xqnmlXQbRBb9UnOaKcFl3T1dxiLwkl
Mb0Aq8/96yfCeBnY+kvJGOGj6bcBlKD9/wbZX0n4JFWtWi0DBDvvQGRK7GHlnnin
dCy9i4Jsj6TliJzsTfKNU1bpLy7RSY9CIpF99o3Szp/IlkXV2CrcMeDFLt0GYvBS
eW8lmXP4RCb25emN4HfBxV2N0LEdowuprEAk0AdI0h3gI90DdoB0SKgx8JjuASAi
BACtKeZensVIeyBgyg8wjBhvRgW7o/wY81Y/jne2qEzKpXKp1k7PnGo661mHdBmO
UWDc9EpqA6fSJETvNSR9rDR0o483PGMqjiKLRB7Kqyoo9sqCNMmqXzVQ0yOT0bV1
gTQeIuc7Aw/ULrArB54n3cENHzzT265TlesRb/aOJks0EYflpzjQbpWZMKfAp5e8
Xc9V+opZMGzZWKTiDlqZWrosi9ZZGxACLtxmz8Ldw+kxYHYuqqX7pBgOobF8GIwH
OeYJUfpqmvKRcuxbPvOv+uVki3AJf1/cUC8eZrsGWVXlZ5ZeJ0qfLeBJ0/4N8NP+
yW+PTp0B8SWuJph/3X8hWf1wSH8btNEV9yXXa02WnKWxbR/ulej5340ltNbQZwKi
lS+cqxxRj8uGBC38U7bgy51TDkJ23DfnMGUJIFRkraN4HrIO1nQ1zj5ZnUYnHh3S
y8mDglBrfbowUY+JcFceyMbvNIqSBzg925x3tmP7hCOcV9UYmSuaAxj+2GjdgGtv
kqFCipzxh8EU41yyn8AC/NEkTrmf2rnSuYivnvFvG5AZ0pqRa4OEhZXHrGvRymsc
I8UMX8pp/WrbCZJErZW685FuWALEH5Mzoxm6pHI3SYeyDbIOCzjP823cBEH+3HXg
/tTANrsvhPNAZRG7jpRw2lgyeI/7SJLjcjLIRRaEAbwN47U9w+y0M9OtNFSxqcpT
`pragma protect end_protected
