// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
f4TEC0ObNcBZ6SlJgWGkomvD9IJq4oxSBi4UmTZTiarFhSS1M4wWbJFvvH5MU+00
cIPIJRacFCFDCj2Zil1/6jpq8OZJWffDir+dcuxTtyotVGrqHFo4+VthIUPwJ93y
bws6sXD2jCCWqSAYau3+cd4KA9ONjs3tYMD5CJNFfUg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 527968)
WPKFsivqKivMYwO2khLmt9klA5DJm0q76vDwoqC+uFloW4IzCJ8tBt9NiiGLhBDs
t9504cAyuwnhp/Vqpif7E+c2DFtHihygVFWhTxgtnAN1tOPeXOBrCpqd74/2WQLe
fijmH8X3S2wdoDIW/7+TF8mrtBZY7qE7PLZpfFhBK3jOyby0Fuw21YEwSjrnXQOi
nTWsNHxP7dLcw1zob0K/8MN99z8e/vP8KZ/ENQBj534u1DziQD6CCum1hpCuJm3M
UQfrhUMzOdxHy6xO8Ga15EmQtUwKJ1KWhAXHAotrcgVcO79f4fdnWX7ANv9z05vn
5LVsYgCiziXblKS8RvC+A27raoPua/MJLS/iyz1CL9S/LSxJ/O5sZp/jGX1zshKL
0SzjLPU1Ea5bK/lb2SUIdWmW/9nq12RLCSdLQBC1vcQU2K+7rUsIbqyJhulP4SW5
aWljng+fuWVP4nwuKd8YhIypx0H13Jlw3ysSGLm6gnJaXKYNZdV6q8ONbVWgoTju
MAnRT7teWOw+vHi+FX4vkufPVVwkgHeMQCFvu3JwjYZQrQdFHJbviViywwSsJmJJ
5IAyCbsYZJjluoNM8Mb82hsErRmvb3ozV0/JADJhQUMOoDkUXT8YG/RIfHtMJHLM
QhKOzqaETLsCvl6Uapja6iMYulOadELe7m16gObHsTHkutSsjPgIdvFcSJ2HQhSX
OztrNi6WPoeXGKaLkGFK9KtMgQ7ChOStVz5uhfYQ/pgMEwCbAh8U+u7k1ZpIFOdg
5NUMJJnu/OVRyjIuL371GrZ4u3t1GUsT3VWLyrdCUoCMKlH0Hp1yeUfPTql6sIpl
l7KExo+ODJefgayTl0UPdgpjxXKaT3KUcmklRfI2JZhZap/GjX2x6vO6SrRZCY4k
ylvQvp4ncgblc9Noi4SbqHKRvtY+aShlae911PEvCbyf88aJG/r34u5Qcsrred1h
swJX/fj2tac8mo2ADnFJKsVMHV4aRJ5jB54IbxOUQtcYJ07Q6ah6Gf6bqVJhkou3
4OAR6JCKscK3w73ztnR+p5fwAgfQQPFnZsBRIQRo/mhZkd2TQ97XAoYwqzSI3HdY
TXf8zkPLhbjK4zvCxrYytg2BZUeRccNUF10jjB0ZXBQ74FsKRIfhx8bMvdIunrfD
Xdtl3tbmG6XoM5gQeOrE1LW/MCBN2a3NKA9kvmwdZtLayNRe7n3vWghCPvR4kBIV
k7PR3SeXDbZFVNDm34ctDpVI9nWbqACk8yVL/BWUo7kvv4762b/S4Xwm6naBFjrc
TXvJQP36272WXvehF+lJycuXvv9nPGtp9pgx3CSXccv5V5ugyR3hq1uy4l9of8te
OtpWXspDp/W75V5WYOaoCVURdoVvFg6GhyWROf8DuxQtkleG/tA9jdp+YIu+LK1w
0RGa44nfRV5GdbqF2zqypG2791RpKJj+FBNFiqQiHCc+C26ZuIHCdI9Ww7uNh6UV
ZK4ZJdX+yYdDHcgGrHPVzwMLGO6gE18xaEgIukXzqbSGVcV4OtYRq1/UifDl7q/i
I3t8pvmRhE0Q1COPlUR5hPTlzAaNXhpWKhD8F69gnukxu5MCOs9Oa7vsH9AZ4Nnp
eLsNuQeJ+QjAXBon5gCmb5a5w2JnjCcZNRj+UsyPru/gYW0G7EYBW3+j/XVdpZHM
pPLbdk2IInzyemYPNH1TLHYc2KK5HF3Xl4a0AfDn3A3k560CTG4OwpLfI2SVdHtl
nRdBYx8a0slf0BzPKRwdF5AoFdcKhiiUEd3PbCXYXuJ5OYCmBQO0qvXV13Mrv8JQ
3pwsWmwLZFKSZztwAqiaerTCEE4nukdwMR9jvlCEKM2Fb2A5SQ0pAndKLnjUIE2G
kCxILY08wyaj/8khnNhLIb2h3zsWoqsgZralG7GgQ0ET+1NK/dBe6ZmeiF25qtOh
6of4nA/DUogSJMbTGu2hcT0X09GjDwvHxUaeH1lDg9jVxdbpapwSJc6lKbXIp47a
1SmxWVed4kXPRSyVHd02yCVPitRfkHxNN7pA87OFkEBj4+pfQuIwrBNd87ICanqu
klKY9wDHEtjJTYb5kOIApGOtv4+Q27D83hM4mCoqg5ePhKuIjqSUexZ1imjh76SR
JRir3dAX5IBIzHXv+Xi1p81ydeSvF5YfczAETE7McPvmwcu3QGT/cST6XN9QmCMA
eJ5yTqdNWuH2V9RPWZ4wxD/x+KmUKRKXHUVoEwpa/3AkQkH2Oo99dnBh639bec5B
UlWGaA3ediTyjJ3lHNAVQxhagQQJqWBt/x5PBAxNiorGBp0jhE72Wn9UCDH7K8se
9iloidMOqDsIoU7e2nYEmR8kdyhNkwPgitcpEoymFQ86IDI5Au5LulLpuu8J7yHH
viB5ZAj5p3ZRVmzXFrDQKsUWNZnn45KpA/IMfdSMi90Bzls21gDbZcIufLN+oEhx
DBZ7lhYrRgpwECOtCdeYS++ICXwRJQX04lZed0eosVPr39mcRcCJvXS3RRtAELQr
/Fa8YjmJpGRbYUORMzQEQe9lnwjYZAQ4bXzlbglONlZE72i8ziLes66yYsDvgbju
b2/IzH+16TkcliPw5s3NgYs7vuaCscD7HDG1REhY41lkDr5k91mD7zVeUt1N7P4B
3Lj5BwDEUKEDRVNsv2sfqsGGW1xat44pIywOmmr4/ZgeuVK8ebuj8YB4zd9tRxy6
1usTf+jK9lrVSShM5xuTXskns8GW/RrG75Th/QfuNERYfr8jbkNzEQ/BaQlwCFgJ
mypb4fq4gRul0VS+oi+0LYnyDW1AQfqN+Xjrduq+hEl1e8wnvxt4FHAgBNjcnK/P
zqYTnSMuuVE5Xs7duFonGtp6eXhu6s2RQ4mtwVIARwxBPeFLACeCL00FVp8TKFMO
aKr1C/Ye8hWfGc52W6uZSBcyunVoSejIODhES+HobHvwrXMoDQwbN78Ne9+xndKo
A22dOz7aVJpS0OpufLVxmsyVbT6kcS7gX3bxy2p120nFfeO0O0HZ8+7Qz16W+V8k
gjtOq7gwCpgCH1NRXK3GeenIXo9OnmG1cVmvf3zD5xgIwmzTtw6sH6bgNQxREtE0
RKTwcnjECvK4rNRxOpicPj6/p+TZOTC53nQvF9QsNF8hA5oWkZnqFVKkRBDFi2UB
DB7mwdz8B9hNXUHO47D2ziyE0UVuey4qwKb1QmrFaizzG1F9wXUjRd4fbHSsS7sr
y5wJsdFdGsa3BqPs0P++Fn4btT8QIU8MU45Hr8geKnJYEvjqQMAgPt8fnv88mmMI
Pfdi9fB2VGf3qFJlPsb/tD0YDDijW+BFS15Wl+X8ffORIDOpnixVw1vZXeXFhqJr
k7HIYw5zkR8WngT1mSXA9yf6CTHMVEX8BqJHrFYHrN6JVe/CJsxAC5NVxSrmDQUn
J+3LIEuAb/cflbsEfqMUoz7ZdizYJ4Y5jkzucGwd9KgFfJTZDZiulDSDYXi/AYTB
v7ZX3HFuzAVc94Tre+CFPO6XMQ56W5jdUTH7HiYKPHMWpcLmGjAj7ILgCMhLeNEL
0ao7Lil8DReAUcoZuP5sCg3q5ipEYoEMwFAu2oDTw9VIPG1ZaHOdJNXEXHrCZkW2
kNKNMaPgqSXzjGwPv5Gm1GuVWhKc1bsSdqeiA6M3AYuwpN2bH26PamvJPf2X2ax9
3wZ94JgEQ9QuAj5ue6hN8JADacvTKUwhBRiXLAMrFG/EdMFZH1qc28m1swvQ9qQM
e5/ToYvIBLY2QWV+4VY+ZgMBe/g0wLTjJQ4gw5vb5ph/z5sbqNCWr6ORnevia6eY
nprwk1ChDSoSDozonbgr6+OdpGyCUKRj10e56a7GKDSItRfc+B4uBgPSMHtBFMiP
Q26axkc7jZgv80vbvOICudfqggIOf98+UXycaxYnDmi2GXyPGogicKXM8QoOcO39
b6gNLpqnVLeo1OkCHDMuHSwYzLp5Lno0c3NF2ZoidGNLb/xbIYahRo2k5KJ3i2aO
u8m375C5tg+fhSGZjohZ0/lYJCYA2DN2d13lkop533hxZmVehr1Xo/dcUxEz97sm
++H5rFBM4F2Q88MAbp2umCZWd/+ZZ40JuQyt10RFl2EJ1tUV+O5e/ZeR8jQTHMaI
GrENxSsOHpMkljLBftAhYQ3dxKx8SNRjacyb7l8JSVDcBpuqr0Dd9k/KR24jhDHO
MRTxF/J3cSGv0G8oe44jmPEMHt/GBH6hlCNlwZ9NvA/trC4q6PkOjhThkDmrTJSp
tq7+XDtG/2vsGmwnV/SMrUrZzj6AqLFmDWzWBX5Rvd0QgAY9J6p+afC7RfmprVNM
daMHbz9fMmoese+T6g+OCQhoM29PFAYsHP4fhxeTVOAot6Xu26/WB0K0GffX9zJn
OsKIqi5rgGbvbhQblwHf+rDjA8Vtcyh55eoyCBuWHRTXVjp5XyV7SGhHT2PdmUMK
jY8RjN/5JYWlvZukRrZjPc9quPyxYLVc2ATlvWzduhU0lE2YY+9sUFaZSNqU+IkC
IleAdWUWsNIEqRl3dPw8Im68yn9FZe2GYZUcJ+rErnu8rWjMN7QjY/fhmY/llnzU
+qChjcAzc83NLtLPHpjLa4uX1ybWRpcGr7Dv263x8UwFQVkBZx+w8z5sMg/PqUut
gC6V5bVTeHBC074BUgIfEeSJNguL8bbbMW5LZYB55GzbRdZWofq892reljokqaf2
AVD7IM0ICt2hvGtLsls3agvTinj+PmswIAstt7hU0RnZDEH3mRRa9JYZke7rL8jd
aDy0XgIjAaqKuHZuyqfr0HJVaCb4oA8Ib0g2Z5TR9bMkipS1Gt7eHWCTnfyxxBRn
f8OKSxFKdY5NxME2/Yp4rrL72VidWPKzkxUPTz3sr7ak2/EoH2GQbotsa6B7t12x
K5Cvi9AECkPVr2Xpx7G4YCwnwbCaSramrb+AnG+nYv6yo9k7o3orXa/zBGjnuwg7
ozogsHHrq/0M7VsuzCsVH/sP9y1bGib7BK5ltlPScu+maneeeEnh/4dRu3v3IcL9
TlYVWFvAbK2JUe3R1fbwcx8+dGu8AlMrNMTUGqC0Pe5cL98hiCxtBYmA/XGiQ0pa
G3CYWRrsse2jDet4GRSaQevh5LZ1DPtPfgINajE5Ce7KvZ+gNwP8x314kOOyX3Ij
KoMkC/GgAH87CrD5C28YvL6+TPRseWhJCI6DS0jUL9jdeB7BWVEH/4DEbucJfg8D
r0ZsvLzghn2RzfCHYnWGhPW5803MXILUN6tto0up4v2Mty07YbTx89DQm/LVXKsc
tz9ozOkJE09GnTkF2OQmyJiNfGSQYuKYyN8XxWxx2/4v60aZgYpxFaEHqkJq3US7
Bh63tsTUYlrshF3Cw0vK8R2aNUR2GKuehHO3SPkJZ8YQS78xvI1vtdoG28VjQH7E
agoBobFQsjmfH8uCVW1ztZtcR0C34y5VcXyq4BdzV9UUWT85dAIAlQWsQ18knGur
8D0LPnyVwTZ1uqvjES9poaemKMV7QF/o4a/owKMC+i5cpPIUkdkZBFpZcpXfhAyO
/3y7XK1nBu8sIzuU+jVC+BCBnQzRkgyqS03ddExVS82X+o/X0KrM86sYNPcX0lj2
tqBm5n5zQDh/4MGKcEfBD8YL4kMXpIcGR91KUFfOSQDVPUxNoOhdhVT2xQQCk6K0
ykmL8tGX8nkj5UtsH46HW17sgjptL3sXcOjp0t2co1Zug4qHSr+FEchPfEOGUkkC
bKMiJEcvp1MM5+cEOe34STbhoY0/ZbikV2rzfp0N6RDm/8WUgYF0PWwifK1eKVL/
vBUBXbOhBb5hRS/lr0ovJYhHOW07vjMruyvLpzaAo7RZZ36xEuB/gEVOd4FzJIKR
fehyB2QUFEyngLMW5jECGeYzTJskX3caw9drKL0YkXtmLfWbdIxQ35e++2p/7O9L
yezbL6zsDZYQb32roxavKG+F1sbLRlADZr/YpZAC+MtHO034BQRXtP4XyydbQfKb
m/hbe1+7A92iknSQ3Ns/0KHEieDDGrZfIfk2FdBZIFR6OWv6CIekMshjRKtbepeV
WLvJJqBJCEoVHll7/fZR8PfjTj0YemOY7aQBt98sho6cfsYN8RvwepcJ9jYq+c/h
9Y+VZsUGKUHBw1w0E/m9mTl2RHi09SkJqWiLeSsehTY2HdDpd0w2S+FkA7O+qTdL
VRcqqG6LBZfTKtAeMINICjD6oIBpS8FXej0YmecZ731/WFeO9M1W58xuAcT1Mn28
eAYaUdeDxM1B4WwsnTI2Y2hwApcVJn+lUIoxmg4AlB52NP9FnocUJBSSaKASTeyi
mCdevzCVMrz9EuVnxy3RjWjq+O/zh0yqtz2bumgOZ2N3o7As2C7IMiZs3X40z9gD
lOyIQzI/1sObGZVNalRg9H4hwsEJwOHALRqK+jp/ZDZx+7zuOxo1vqMSKXZ/crBK
Cg+0Vbp7PRUww4Z5KNMpLdphiVgtkvYw81SqlJPdGDCX3kbLWkOd0QGoCbCNtnpE
31JINbtIZzBzIYhY18eRrHWtniAQ+B2YP2CpxWs/+XZfKKoFso6Xc4Ndl6O6J5ED
RMpXgYpi3yE6MjoV4IcVXO3AXrCG8o+HGmNK1nTUj3ERr7jDOoW08vGQzBvxM8+P
JEXhty3vsbvOCE279Bf+febtF3tjHnjR1+WIjW3AeoUOReLPi+461OoPpY6t4T81
SUDVEduCA4qr9sH1u9zJPXFHoQ2jpIkexPcbqGahq3S3YIWnOqBCONyLCnpCgdW7
FzbZrV0dkiGvTRnCphMu6md1+hKW4i3HMKAPZT8b6/y1N2VS503l0e1SqFm6Dmwn
P4+m7dkbq8BRQcDlxPgUUOvaCz1m3q46yUX5nQ/8G6lq8219jRwjeQdXyTIPYQTU
lrbVY4Ea6Mqi2yxLjdrAGspBWiLWMsAFltGOiSPbU0wMP9o8wL1peqNIUClqtZZ3
x4leeYcfPqGwVxedQx5fW5c9IhU1DsFojGvQB6LMgL2gM4bNwXtvm2bmc+qHhVxA
b+qd7D6oaw3inoowI4ZutPe03tcj+HFC2hg7oeOFT5eSq2PzMcJAbRPzIuqlwoiv
uwb7FYctQP9Ua9par+nGFz/7VQg4UFbN5fKb3BMby+PQEU/VOofosFXSYBMLu4qc
UqmqTUH/amO8ldTBlVXeAcjwPIXnbvudUyfvLqTO8t28MUeDr0dYKFE4DSemXfbw
jN7CS4xVFgoLcCkPxkFXpAuaIaJeKY8Ss9Vk6hHdQG/YazokQz8lr/CbHrAkzNQO
B8Ixtprbi8v5NicNBUvjqlRW/uK/Nvn8MQn85HglaQ+y+V6KccdiFVH/JJBC19/C
WbT0PnNED4pi+M8DXImKQ6Lm/Fs/48D8A0hdR5qfEKHYm7DkONl6BcCsa5yr3G8X
jub1IW3pY1VNQDckQ39KRHdDUYYxUvon6RAvbkX/aWQ+1E2qGECGG3aKv88tVbz8
QFQqDgY9R1tqOrPF1q7F2Vbzsd5ksx6FXCUTEjnF4pqCuAqlAGWTS/qYrnxt6/Hy
vmewUlrdru775kSrSGQ2RqMpQWiUIEtWnCRw6L4S9+e2ZvkArZlnbiv55gi1Cp4P
yags8ASQ/ReaKxKhNz/3nb0kc8ALPdPw0EAMTFokXMFs9CZjKsw2OUDOw+HTITjy
oRbGDbMnnKImR0CalbRQSntEn4l/7RIZH/GAwcdwxMzU0RbNlw4xp3SkcHMECtDL
eBPSGLjWyH0t0DRu4Y+d2fvbehNduAajNJCG7Qjs3om4aLh85kyXT7hlK9vFbPQr
p+MflDaEADKeAiej2f5vX6A9oTfAproJV/PRqNsyU6T9lP5rHAm8Ze7V2+m0ECp0
EJHAz7yBOQIgCzp8lUwxXx6MEPsM0LLAp6cUpl20mcsG8mBG8wIvLdNGWupEVzBi
YFgPhXXaeIhsDjlmg1PuRYsN6Lhn3Q54sdV3uzpS8YdnNDDEOyX4HNucn82w/7Ij
q9iT0lTUjTsKTrkRVzeAozwumtMKg/w9KaE2UcljxVXfoxFRKxe6rThPQhJTa9Z2
sN0GB1SfmlwlSnnFk1zcUKbkZgKP48+C1nE9+EOC3Bnoj6eCbswosV3ZT4Jb5XPC
5zEM9P+NNI2dISG3Mywla72OMBg2qMllTEDD3oRxh4KRY6wb4qufta8GGcaRdZkz
AUyaw+vIE1uxFvtBwtsTdSxux8TxdCsfXUIJsuPLebpVLCHfODgOPdsa4UGIw1Go
F2bUfihts6Fa7HG2lYMLtDlZnXKP8NYE0UdLL14FMd5KqzAPzjSjcXN2vxnZSFti
2dTLAPtXTaVRtIGJsvt1b/VjJumfNwE9aliQHcdyDZ7ubvdU7og/c8+2P45sbOFx
9WvR4reE4Z0jhxxUK8QlDVOMS2zmpL9uRj6GpPCffZNdxoyJ+F8I8IEFeR5loRvy
fjd2BzenGqNQVXG6MK+1TLfZRy3Az6he+kV2jyVjzM36RV2GWvLXyPA9EWYuc2LC
XdTjcxpnkHeuToCDZjl0qggvMi3ED8ggOseLrJRA28XOLZkoGpqmep/OyLQrjmcN
LWg+n3orj+SvWCIfU5uOnDV+CbcZMplDoKB57hkS/8HtUrLy31QqBx96IV9ZRRMQ
h7On8Dwdy8lLKtmbwmiPvYB8Gw6HRH/6/54CYF0LIDhzodaxj55DJ++D0WSzzpTl
odHzuzf9SN8MZrKAVgGVYKgy0qAZqBqURPPrw0UU2sRqbzscZeJWHN2lCrdI6kFk
TTmhYB42pRa+mDaOd7bKZAQwX4X1Z8yUTMXm/ALZz6xH5YR1Gl00SluDK/j/xx7u
Y8c5MuvKKUs9Rr6n6cOsV30DSnS0agwv8iiTWcS1wlr34F78LAm2jPd9+6dkjJnA
gZpETFB+J7yD4wfgBRNjxWVV0vSYZlvt6M5aF3CAWNAet+kJJmq++SOUEXhdLIB/
OswW/NzrOBfQvuUUhorgT8M+af5GfNskpa+r3ASU+RQDi3UqCCv35SUOWxt+s3hs
Jq/MJcdtVOrptNRZMYMhtS/1Y4KF0A6SIZFqsPwTJaAWSK+6nH1JAfsTwD7uG4nK
jQIA+h92e8J9UHq5p7LOCKGvf5Z8kaEvDKY9B4NQLcePe6hWwT2glSjlktnr+M+s
Iy1watinSmDNyDkH2uzewaA5GYiuAmw4En4MBrSku4kcApGyK3UB4vNtOQgodoSd
epQN93pyCDzVdj9gvq32UnHhmAaqsu4stDv7ri6rce4F7V5fNIv45MXZngL/95Wr
Hwvn6U+Grz0+n9XPlZ6RsF1A8hdA7EdlyzyDAHj68ct3AM6COxe9hvhIIBi3MrJX
EAJft394MjPxvLK5t296B9GKYh1thUV9XqXFWeGhMmSgdBdMrh8I6WSWY0KzF2tY
10hfL3pOf4TxL5bGHkJXp+ESIUWynaxZN+nFvydnPtbzXP73hyywBKKX1/yIrakH
5/c0y89XoPqrdQWKXhsjHiTmWcgCv1W6MIruXVfnQv+Jr6tGRQYPt7i4lhY0p+9l
Q//k6s3q0K9MWF5zAB5WNoHts5CjvXluhSWqU6lvXCqmqNH3p0700KLNGyD/NdRQ
tV3I4RXTOTHzMnx9qLci0Wb6Y5O3NLytvto0L9zgipFiUvoGi4CCJMY5HM1AvmX7
WJ6eLrCIjxmSYcxiHX6rUwzzK4b36AHIJGsxQ5ODJh+r2Lzid5sElmNPg3otXhZH
YJOHxVKiCSjgb2NshpXK1HR7vWHNTGDz8S6zs6estnd7V5uGuPtJiHTwt37+Icsb
JH9gS5GkvTJsqgac9RfrHgq8WJf97R2Ggcx0lLj7keynLYD2zkBqk/n40gcsN/Ub
6X5ZBqfQrXfnFV5AHOZSWfic+/GO1hPO8J/kqxZLjwmnzum6jzitJyt64/osXrdi
vX0mlWwZYuEpNTuBtSD9jfBra5ARKEBOLhggFOt1TvNp2J+zT0O+z7YQ9JVsZoAK
NBN31f+txhCfWDz4ZwejWoVeDHT8ly6wRK5RAWArzxL29pZnDWeCK/OZDed1ayAX
bud2dxiETrIpksGKGeCgLsewAvCKVHeqDqoEK5Eu1jaI4XHMZbXUbr4Shl5FxZG+
05DKR4VUTBpp1mvGik1uhNacr6iFupqlIdkiF2uiYggt/sIM2WFQVhoOkaAYjVHM
CsJvYQ44usXT9nfIz0GIQIX5Lq8B9JnSgtnz9tgnTv18xBWZ78c7aC/DmqqA25au
1so4eNOq/BqR9Si0r0Jw2aP9+6/zkd+NR2CXwEZsPHrFqg4qmcbCDMN/me2KKiAI
gwTjV6jhHhTkH3U8FE4tcKypma1oWp8ZskRq8zFW0InEPdPbia/6OeARNIT1V0su
a5onSlV00i1k0YexvasXLXZgDa7FgGAEuDc7aX2DEWPCZj34Y0urvZ5BWT9XzQDD
ufqW0XloD3LzdsxH4XksfhPDcWGd1iFuyMBHDCNcS9K2kYcmbMEAh0yN6/mZrtz1
r27npL/YRm0Wn03mNews130A438OrNJiRPibOn688wy+Gp7QYZFgO3Zt6m/EneYy
Qhfr4F01OCwFOvQkaex1s6OR6OwIqdi/xDNkT72qWiga3K5F9BODdhsK9+LZp8aC
3ZaELLY1CYVdICB/Pl1Zqhy89kdqFT8sArTjYzy5tYuJFzPojls9BIPWnxSBgWqx
V8sN9aC/R3xu/uJemJTGAqXDVsFRDvCUZh4g+P+Zs+WoVaaN78yGJVeN6JSTBgq7
V+OXzg0Xuqd5+lNfUUOrQ+70j6SazfqOqoSGgGzL8pmT75gQ8Imy27MdSjiDDS+N
f1bjSx72P4S76o8drZuDz1SWIrUa9e/0dbxGZOGNvFOAhpXaYOAGNGNDnYF+pgG7
gSVFvyFu0GzyCYcPQCQ+HniV+NcwgwGzzgIgXwyuN7meXnA/COuIkWxCHEEQHQDG
2HVffLHcZdf5NEOujdlCG+w+G+3RSy3NR7eTqZYYtXlq7iA3EzDXrsppXlUEWySZ
u/Bbx0USCKe6nsbYhz3ZdZi2EYYep80AXGc3eq8+ey6TDMdX0EfAtP0xAiNmlI7N
EoxiElCBCvBLTk/D+lTgY+44aCvyysKcxomnJI7sxqQUuKsfk3yAngFDmts9w21I
nXI6cl62DRuGneJuhRc1Qt7l0CNNtOMNFWyLruxIKLcF06ROOY2v94zdHLLY9QfD
t6xHYg4liim/EFaKtOjnsUvdZRnS0PwY7wz2ZithwXgvNrv49FsGkVqiLltrH3iz
/gt6Zi2QHeSw30D2UZZCLa9Z3ZUTxbXyd4nOUSL9RlZO7symZPq1dfRRYuKbDjby
LC9tlSMMm4oPoWv262OdrOQ0IaI43JMmKQQQoqz9PpAslXBLbQEOQah0QDwfL84E
Yn5X0Evdq8HPm/1zh4JzUAAzC6dz/dV/qPVpBpxwMsIqlLjZ4FeWS2wnVYZHTekW
SCwwU8O7TDaqxhTZXHEZi4/u0u4UbqsFRlvjHwZYuVn22+S0wsgVwv4/8S0/tt6L
d1JKDYo/ztEGpHP0Vo72lyR3NZi+4JJc9Fkjte3MYlusSo4SkX2X5DL7EP1Li5jn
HAas0Z+z2892IdzDxOPChlZD1MRkL5/zzFpv0nVZOLi9bMYMziH+ZfbNxYgudRT7
aEViiZRK45TvE1bvSfdKLbVkK8EKjoP4a9OkKfNU4/Z1fOu242t6EJ+csG53fBHo
GpIVoHnRY77bzavjVNmA5vCXZ1Y2qZK99Hs4ilpPbMjjtu3zBohjY8dYhTJb9xVq
u1Z1GYsi8P6VXfnoNiHneNpaxiYgiA0t0TZOHD3zimO1BTppPFB31l1frjm7ZYCy
ckTVKaki2aQCfB4inlBEI3KWtlPpXdlAx5TWv2VRWj3Je7STFA87FhKw5z91NVnY
bFrjuCdanHBL8QFP5S6S8Lw2PGC4buMmYR4EeBRY3XiPO4oRjLZIclEoFnv6kXAk
7aVG+FbrGOoWMVdZXTVIXR9uVBNHJIIdbltOZFMij6/I+FWURvUzx+ooLuyJWrMS
l/0Qg+v9+Ru8fzceCJ3mBlmne01j3KXpu7in5dLhHoGVPHmRmUQU+zjRw5/UnoA7
7kUk1+diBU/XDkS3JIUwgnzgy6j6KSHhlNEK25E5SfBJOVhzGtLQY9nXf0s3qbgG
lH03NimbsIPbWxwxqQLwqFz7esqfKvJf7vzlzPtSJd5yMzlyIRtRarzSf4HPtVUn
wAD9hQE/ebcClO6z1dnd282wwbZ8/nLqbAjO+wJ57poeVZzGdFNew9iKB7vtnNci
FxBxSQ4MWNT4uYOypblcf3ad7RhRBrqumY1vD8rIOkYeV6eBn1hu1K5WpAFwxroV
IozP8YBtZJCpyQr2TTHhETKGTFw2rLmQjPgABiFiuvlpTkojVZxvpG6cfnEn61Ao
HjTjeCHdaAxOr9S3JsdWmHXhKu+IKKdd+ufQVGHqGo3ZVFyKTjLY95ytE9lIQm4F
pXgHs29UGk9d9a8fT3d5rssrnKfUPYa+3kCF+X65l0fLlqHgLAPpAHb6QrmtGYTW
6uS3YkTozaqtOdfzAJTRjdPHvwHSFsL8FFKaxCz8eqpA7CWP3q32CMbK4paYdjZx
W2eXyOecJp37998KnqKAMDh8VlXgFwKyLeK0vHaW77DIgZvWxt4shQbRZCNXNvv8
vUz9VtIRQVZyfBZpfgb2s5YqlcqwLL3lneYuDUm0p0qYwLTyjC2zQkD4a7apjquD
nZxJ8z7fF7g1D4eOo7MibtQn2d/eBpUJfP/X+yXEa37INnNMlgZPSKzimpIETLcl
qa6yJIApy+chggQacSuMexgjPlkqZrS9mlOMrqFztj4LRrDZNotpqtotR8HxH458
1/myucsMv3IGmTPnB/hmxp+N2qBb9nXQTbSgJqNHee3VW2sxP2uMPbajGl8oMPbF
/tw3cKMFMpWa8x2bO4TNkfjwnzM1RNbvMoOW+0NOxeHWrce5u9TsgaukXk+FjiwD
7wNRmsTNSofo709x6uwYtWaXlSSXe+HDFqGbsLSQxypqj8lSHhb5dYQAJtpPNRxE
lVRwYukHTHlr/hFYPyI42P5WoG1LoLcu/4DCuluDnX+pux1xsyLTqU0NXfXNooSp
VQieGlQDs4Ex7fqCHbKiHHqQW2HLxXb9aRNIjr6KEDaSKUzAC4hG2g88WY4hSjy4
B/AKsH1qfImvgsZYwgcFJEOTfGDTULOCZx5qEOEwXa4L68YdYPxFYB4zWIHKb3Wq
vitK1Fs1akoOCK5S/EimNckwyzZMNcflAOLViAVcCn8rHKOXhbYQzjKwppXRO6z9
grEVvuGYsunAxHDiha4kBxC7w+Cc4At+OZZ57aKeQjV8X5t+2RDWDR4XPu4JxGvm
zflQEjbl5N74AF9bGhm1yY8CvCinh0yAh7KbHQ00zlgE0KB48RJoKMwJVeyM1fZS
uaH4tzDJDURnbBOXItYOkmb2dsMcXsqi/1jMo08Eq52Il7jbBTbFwsBn4oYI+9Py
SO+hT5T0x+0flqzOP8G8gnHgBxuPEG1RB6/sKHZwyGQBFYABAgvfbIH6+XTZ6iyu
vDAhkU4d2KEvJCuGT07uJWK9ANzsU4m3+leJRrq3wDPjEoBC9ExisH4Y2E1kTOhQ
2DQj9CWlGgxW6rmkANtaJCTVZ9hm3KTDHz604FO1WWyqt6uZNPR/f0o2DvS4esXO
29T6+WzwQWuMd6iP8LBIua+QwTjiRIsR9/9hiOSfTwWm1MXCHDI4JpvGihHj7uLx
lwnupUjyOVoZLZpqf/krQauBxwVjOB6SugY6rAtFhRjfRXpKUKGjLZJcreZf5sQi
oxUeyDGMYB5tjzgapE5abeCCflYAPLnFrU5kqit1nHQQEtpyUE1z28vKrRHt9r1r
R8uZKje1BSK9zb+l06JNZB4M56LLlSLZWg+MIAVDxS6K3fipb2rSHDwN1itL+db2
0NyVOFon+pqB8ZlTz0u/4bUpBJBXI07Jr++YieJPzlsNLH0l85Z3WMLM8CMhjRTB
P6iaPANitpBkJWLNxdOVN4WCsYQufu3S7elwj9iL3GRJksVTIZy0QzMvKXkGeMmu
zLZcHuaafAMTHx/7/Cbd0wcZVDusraWMvYn/ERwHekFqBQbOgW+wP9cOBVV2BCME
/4xCAahD/EyceyYOxFADxpUKf7SN1d6R+SFSL7InziyiVEh3kEBUrkakL6sOKvKc
o+2q5rnn5JWemOFDrP04qYEb5Xt5NE53IgbXsUkCRlzNRy7dHqbzu8c1cYG6FKbp
AYf8cRHm8t0kAT4SqkCV9FLuaQv5l5cLd7cO+GIcXb440zsGv2OQR/GCyJC+LZzf
uL+ehgyTaPyuRSfj17mFrH6cAWj2BufM61ZH5GLd+zuqDwtGRiXn7cn4j39WUhve
THjwsFzz4jm+bWWBYa8BLuHYBBUFcgux6qCxCWGeqqcZVKG7XXf2sqMdpVE9pRWn
OxyF2V7vF3RZS4vlu6KnRSe2Q8b1V6/jGgTD1mcfIvYd7GV4REnO1OrCeJ5fabZM
oOxJ/Tu23f32xuAWVZ9r6xoPbZO31emq5/0fj0zPM5FQZO+vrl4FTJf9r71/ywZs
Yr4sCH1dlmNbdoh5cd0fJyzxzASy8xmj0JBmmoykOpcgaI542JUY848PHi7EycB8
ViAgKtfU2D8RJ+1wgjnkGfKWrs8A/cAAzsYAV4lKsAk+drq5oSgCsV6FijYzHu+N
7Kfm1SfzRq3Udby5mfpnw/qXsxCgDUqJh654sry+eN7HB/Xbla530hs1etiBzAPX
z73yucX2Woq+RD37+6n/uqzXJoz5MHhvR3Wmi0MvihwI9rU4z9tASgKWPJcSjkRd
M2BbarYndsLZwHbW1Jgr1e+zDt3PGpqlAezIeb+VcYb2RDnAWXc0tBi7g7G31Fj/
35vaXaMdkOxcFJiuVv5v+PT1ySr5MijKjoelkv1Q/n1hHS9Avxk6qU1iGSFv8z/s
FXw0uiObG7cLwfXSL7A2C0iedeGxFv2iQEAzfhZhCK4FEicwu4xjUZxMDgP9lnQJ
CvEv+ZG5RtwaMtR34HW/m/5xr7XQy2jkoXqIZZJ/aa5TihLWjzXxHKpQWm+s2ak+
YlBnYLNkTjkusitTmKvn/Z3MpgiaWMJ4S4IBgUwRlYV8rZjl4N1zrxZJ8dxYbk8C
MMsEylxdcJRk+sL4gXXvrEyYxDiNzzWdnceisfGy4IGOtmGANd8/x3Aw2xEImRMm
xTFf/LG1+cNVMQ94YzltbSqEgKHBG8bcMLI906iHjHwqWRvKfrh0TAkt7ElXDXBD
DmMcUY3ptpei9p+9DS56UOCEM2uVYtCVGutmKuj9jTmA0p6aX2tcNwUOmyqd5GHK
eX5EUVwT6suxAP0f8h9B+onaxLkgwFxo1ZdeL9Wnexx/yrNd4+o8hREf2djkI94C
XrDiVO1M3ZbmgjQ/pcF9NLAmct6aZsK1NlRCmtPTHjMgQvDHTDo3T6snjIPPd2EM
rHjzjMSfSntghH+/PynuqcJXQvCG2xQaLt6sTx56B23vPMUtFAvZ7pPqEpgnnCdT
4C8u9cjOZ8p6QuOdkJzb5R+LiHnIo2Q0vQk4tOC3k2IO9w4bliCMb5Lg1Jm/4N4z
noWfXPfgVGD+VvHrf3WW46DtYVNuTd/UTmrZk1N8jz0bXbYpWAesFcepyj3WOp57
XOJIZcfw/+Ru2QXWesy79WgL2U/rmI9tgfu4QWPc/b7tmOIPpLxIrsqZOyBgzxlV
mcMsNCX62a6eHCTWiHqpktEw5z9cH+42IOKQL/TW3KMwq/fItU0WiLJXe8/KmYEC
JyLjm7qGiyfoA00DNCF4abTeIbPLyfn4+e3+RYieuM1k9f+jqDlMX2l+KEv+UDo3
FTfJM6Zl/WaQWvq48RMC8BKMKu+BY9hNR2M3znEsZG/H18hvzwv7huL5oWFbKmOF
LR5dkCJQ8708iv4s0U564f1V/Mm+Ndsf723BSIMQuLF1LQx69YqO/RumaocCvDK8
HcWCzmMmA54hTBv/prpEzHsj0L7FlA2rbsKC4ATYE0MlDseqazCtEQFzKQXT4szI
Av9aAnukFDMzeJOkxsD7CdgkM8dG52/yX6w30wrLarVJaXoOdHEjwG1lTlTu3TvY
RW07DlJ1p1S0Yui3sRLZDzxRLUcMvQ6mYXlVqNEL6xSgesDMCpGtaxEpGHWGPLfL
GdgPJtWd+QbwW2/g8/QNzplu6nldci04yqwmnBnUbzSDXdKRGJs33llTO3gxIgQV
gU1d1hIxfSXCCm2ou8LcKdtixOeFWA9llf7ZL8MamUJjPjWtRlJBhENDDw4ybwPx
oMOfSONjf1fRzNGozeBTEG69ovxPvF8X/c8g4ePSol0imqd+PXfE6fWlbExkwHto
g7YZU9VU+W4w1tXWmY5+YBAS4XmOPndRd8JIUKkluWoARHaDgvyEQnYUDmeY11pb
34QXUGdm4kuI8+rt4RHq5DMjzLGtlON+88TP3cIRtlqLFB+thwmbtZ6to62kHnqZ
XM3mHKLphu/dc/jUG2znLP2AqxVG2ZPE/BG2Tv8Vybkk832Fgrx7W/cUG0seiTxE
1U+FA9JOc5ajTwkqaZDhllFLDtQD6nCHZ9+Uojfe5v4Ej3lObTEMjnnT/fNKFswC
Nt/t3Tay7pHdPOB76NUX33lVzJVoY/JgRgA1G5KflhEjs35bYYwoGnXbFsPRqoQS
yKIydPb/tgzelHkZkhcX8WnGwqxiG7hRMOF5M1QRR+F0tfG8hiAjvoepeyaUJFps
wIwNah/+Z4FfJrtKVAsNmlcJxzTtCBnWahvDMfYPbM9D8iLq7AkgQIozCgrLPu2h
NwO7jvbnjkS8M0yjKERXC7CZEPAE8hH+9JOBiKufapoy+Tf+bSWAh4ZEkWUh4UxD
w6aUrklNoKe3/q/kY2FtcpwBK6FjFPZJQONO4x3dftIoY8o71Anwc6L2RB66IrB8
angEfv/hvW6mKjW2VAwDQX/w12CMS0bGS+JGIBdsLP7i2HJzr8LybjBFXUpWGK2e
l4hXPRh1sg4LYZRXqOJdznDjO22rkJCJiWn6UKZ+JpIW5RdWfLCQ+Ea6LZlGFSAy
B1xCmYdRh0sPat+aJqZ6O/V4qcJWB3R1W4phUqpW+2sql56PcPpI/NFvtug94rQe
4nQeay9WGRRiCINKLYkf+cLaC9g/q7SkwUWBBeFavyaZM1ckuxhC8IvQ4H8KXGBN
AtOofqvuR53XkCG/rt0mP4La37tb05vhWf3VEPSBcN0bNJyocrqrm+5VLxIfOWoa
rFB+61TPw0iurMvWgd4Gqr/0wbTXntMX3N3Q4wwuhmX0Q586//LEp93o5fy6PZWu
1aqR1KoeNUN3GilUJDwKhY/u0U7NcpWRl2oZ5ltOyraWr05SXr6M41nbHKm2j3LO
guXhI1XsKhaBSKbNYAfmZW1Tocqc3frHFu8RlStQy5xBrb38v4dDB1FqUAlswfJn
HUpneMRZF7QQTkjQFfNCocIzkGQycZymbjLHniQ4E2I5hOyJBP1DOSV/lukSPodc
It+COlMvJddaNOD7ohKJ6CwSOcpnC7IWDCaf46qm8ZQfIH6sHHjJxK5lqROqnlKU
UuEWU+9WdFQ3XRfSCqsHMOOQOe461wdmfzsbAxskzAGQyFd8ZASk6YH3XbS2xOSH
Jx42qcm2T9VZ1pnhjgAv4kFuk2cWKoBbBj9JKAR41x83KnyO9VffmU700ahdNkjH
PLfP5ShjK/seb/n0kjB0vQB3w0DB36imbW7mlyvnZSSF+DCKQc5ts981t+0x0MZH
JI940jiZmNEE+nvew9fjV4MUTO3WAgISf76DcuJC+ZOpRQ3lZGwXYuTrNgoFTbH5
cvEh+qs990hSbXgbU5olpNM7P3FPhSiTQB0xaufQRygVvJrGi2EPvOrsa/hQeKPX
b0H5awNKuUbOd2Ou8TO+2nDyd7Af3/PSBpCRx05GQRDjppO+WDMC+k0C8OocCGQQ
qJejoBR3ktAqoVZ1Gu5mBuz2zG9YYiBTQDXymwr0iR04TANatVrZsiYHJCs+rQIB
FrwOHQ4U7WonXFWe05nwTslXhyUbOesBpnVSqWHBa2sGIXlec1G8/NOuKWl3JVLh
YC1ipbMPk6CDifyBaxvMjuc0HlDuuMr+ekDrYJAqx/JA/SZYUSrCKGM4DiEEFF1B
zrD3GV3+aeT/Et9hmC0Uq80ehtGavBpyGIMbiLQyyO5Tf3UIw5InprueDgcgZl/H
fiGS3Ne5EmaEqnWT+EGAKOjeHeiGHU97yVbwle4ie3FiIdd0xFSeOM4P6FpqEtpA
wsip/f4i/fUgkTtoo9XvabKH0VYQKQh5I1jN8Go2dUAkcCpKG79vASf0ZLf6i48r
xTB1LMEawuLXG4PRpZJ9MpCATDwNpnum55hITDnR4+cKxfiQAuSQSrV0V8XFiorI
6Z0rEznd1qtaEmTbJWP9Jbd4LG06ZpIIqwjpKdfHTXCn06e2QvlTkJulJQFqMN/p
jMT4QHS2sbUqXmUc2wVXA4iwkES9RCRG6m1eVJqa++5S5E5lcPlnBqMybChCX8oj
hUwTScMAmcmNVoevxE+eTy31PiuP9SfwanL1yIUFso52gPYCBPxoO1HmFIQ9aNnB
7pPmexPql4RuKqY8fESG4jKCr6/rKqtwjKBhvzCXE5faqj8NRV7mUIL86dW/1fnn
hTbYxgR1BKa45awKvURbo5l88Qmu21Eer1MKN0+shquPYH70Nw210zYiXZ9Kf7DF
j2DX5wW/rjLAuXG1JD3R9vr9wZbc4cV+vO7OrmmxHxfNbEMHqkw/CML/eAcVX//L
5wwL8U3CYhgWs1zeWxr+fwmxfU4esskYtPL85EtfisSqZwjo3j+Xhh+5GUjI4OoV
X9C9rY/vIEYZ/n+MZzposVFvQllR83egV6cmh0l8eNckQv8WVCrj3ksrf7TiDVIy
XYuiwEtIUxkm/7aGhupZVE781PythzbbZ0SxXbBtgPYByjhlzrnAoCquIArEdAqi
t2ec/LuXwr60NmAIwlyZQL6h0+orasHcNU1HNqX3azDmY1NfqXU43KszBC/xhR/9
nkMvUs5AKP8XipPwGAcpRCRVnJ/D/wEI5HgBQGSPpAqDbAzZuCmzXkouLmDgrrec
0OMbu0Aoc/RqXpuvlo94hWYk7+dGbVbv59QRB/JEcz9jr1v0EuCsUpLd/iIGB2Ku
kwwU3fYujm0uF3Knrp9cPiPl0ITnXLtchiLVaza54lOHhWGFaas9X8NihQc6Fhou
peW8E3I2zL3HxIIEISoBZZ2tCxtxeExPbiy1Y2ty4+ocGoqUFsIHfIuE4E2w9DHq
mzFSmLEUYkCoHlD6lREtyG6pFTkbGTh3NGVis21QpvpgqcROktr28vLeOYhZhk/P
OMg/nkqiHj9QIv2A67ooIOtCfNi3Pab7C3hAD5WKQX3hDBpfotJIgCJwlTglqjS6
wGLFvyEfljue9i3j9xlQT89u2qH5DNhSC9rH7xuY0SsjMP6kj0sxjV9+orgVPpSJ
f4ZCmmW2CSyRCqVohG2D/SDx9WJhRVHMR3tF0MsTwVXHdnEjO4xnSTGFseX3b7NA
ljyOWoH6qGpFdPFEmUADSsSp9uk1kMKDu5OddWklYJ9G0YC4CbAf8hEEFdSovCT9
nzM+44/zNHbb+oXqB0C307adLC7RsoI3UxGpl3zCvM91mm4/w2JSROx06E4/6aSb
xYGjNUV9NI8bisNYL1D6VptGqW0CWw5gS714vPbko1SQW+xaCtG1pwnRsPup+Gu1
Ka2GQG4G3WX11PtmOTgTQUKMC0gcvWEHTBrHYfxcHGoYHJ0BmXQg95yFP065Gta+
JsKyTCX6X4oPiCEk07y8Gszwnz4e9aeYY/vgtMXPfYbg4pKwrw/Nodv9GaVNhF5H
czzvb1Ao+sVARxyRfS7K41ZykJhVtuTTiV683KqeVaYU7uTeED2xWAr5FtuUN85/
ppicrrUgSNn5oO3zMuN2zUMD2TWS0273Z9EWgqauJHXjTrNCRYtWSQzOd4+4Trh4
lWr66DRUgyLdW3WJYs+6R1vpSAjfPVBr4082Fq2vW3McFggmyvBIDx8R+OHtbL4h
P8ybsn/03eKW5d4MdFT4OiSmNIUFg06FvGwiotLH0AcAOBDHVaV+E7LN3w7hp3tV
HvBhUEvvvtgUH5HdjZ4BEaFpLp+iadhX2IJ6Y3BpkHNQPgfotTRVvIsbwsGxpV8G
IgSQwD+rat6zW7uzZUO//Bo65GqvEsF6jT80OSTbWsyjt5ZoLvp2GDz7hYDEW8yM
JAc7VwltyiHh9sbbg7/s+KSQz0qI7LUqiKHI7oKWVyFDP9hVVidN6cRbItvD/Hs2
eRczY+O4p2GoXvLZbJNunSSKf65MpqhZBidOUCc/RNB8D8noyoXxFh9mzAr+keeZ
4vk/wl49yrJlFsDHjzrQcQtCpLeLMci1ENjO+nh6dOd0gs8JeVdAzC3VIp0XnRh6
WlL66TLXP5XEUnEK66Xb5V0L7IO0T5Lk7liZdWeIpklquXBhdKVaRNL1+kF0VplP
9YkvhXHnXiSFbOj7nE2vNisXM6Qjh2AhPnBFy0lqohDuHSSPvJGt3cNflqVEuFvq
LIEkARxsg6j5AJrHwDxKFGIbHcMMcwwFqT5trDfF/1If/9cMfb8wNYFZOT+qm+7M
nsZME9ggqgutQaNDs6Y2BSRWRii4iWHFchyJI2pbILG65lecuiQBT7Lgtc20Iy1y
N6AzlQRvvz9g+TarNratLDsQl7RAPSWcw+f+nJ08XWqVdnVhzQu6c0+NHHw0j4Uc
psNRvp+j8JQQt+DYdpGbe3qO6ODwvj5QhNrF7YvDqVeaPAweGrwFDrQe8Cr6JY2q
rDWGA6KTAbYwWVN10+fPioePsEs7dmYYughwRpIT6WGOYJWW+c/huN0qUhobDJR2
3cV2Gw3UHO5VHZIBRS5rdav2lIN6MS66oxHaPuyuZBqEc71mjYRJ57bzcXi2ZIDS
fF0GXJbSXNXDgrC3j/N+SnfdX+4fnlkO5/E0Q1/KO2ec1HdIGqMPotZygnU/L1jt
hPx25efOp5BAluGSM26qA35beAjikXRGl2I20yaIr06toAKC20IXpRwSRHWBilny
Zk9eQWLoWBX0sKFrpUkmtoRcNgo6QHWvgxnMld+buFzGTxZRbfFwfXDvdCaCMsUK
vRBuB3hFEYsuf/Fv60zzXhCOBapl5CVQ10XXjHIVGt/EW11zUcQlCA+otrqyr7Hd
0j5AMWU+oJcT3HH6/hF0LOpzfWU+kZTSWqVQ6CGMZsriVYyff0MXgd3s88JsXnJj
PCcb1oX3ijq5NN0G0P/XWCo2560FJ9nnANdZH37uDSdiFxv5W2TTF2w+bXrD46Xi
YJaaG6TQVomymnXCTm8sSCrUw+bAt0IHdbLSf+3FP8OlDhuvMsMzT/T/yRVWjJol
C3TGnZ9B/cZcYOGF6wBvcSgah39XbJJBfMLlGEQ1AS1nMchqWIv5/72anoDgt7uC
OuxNdBvlTnQuK5JBoaBLJOCQDQAWeksMrXxoIy4J9UkuR9BjSmiy/mIDtbwQf3ZQ
oEYZb7k/QLhwoWC/A/154elC6M+9+M5IEjOoOkffLTim8mmZkHiqyh94f+PiAr26
z/HxqDoN9LIvk0Mj7xUxLxPBF+lw3FmjFJppgcrqDPprcnNAKaTD15Yy8mPbZRpc
i7xZE2OZ8FTa/IYpbdLIOQW4vS8vBWeIZpWEHpRdXai+gxzxpk1Em5V6MEwvUz0C
c0X6dlJ45YiuRqpOKBCYDHYijBstR39AJNS4Y1iaVWxCaDn721qBCB2SIGxsdfmW
OuJDnqE0brNZBcIBWx0cyRx40H7z5a9c1fQwLTFQU0jaOXHDGcmDoO5PmmA2yv0o
ZoBPblzGtfiAZXD345kN//UGUjlMGL9R0hRKdA9A5JeMiUoqEJ4+Ko1BOkp3ZLWL
KhG1o4nDi+ABYmsr5wA2iRMchr7kHQqCXQWcf/TtWOoyxXdEV9DXpNvy/8QkZPiz
xxhNF7+pUWe/EIHvviiKtmy7Nkf8WaPgIfPCSikmjmKhs0StwPcj5e4XguqQ9p5m
9CsVlB2X6vjOcfnrYzD7jxYffsnzUXijYIlb009KxzpRyvw2cIuGlv2JvzXU++rE
3tTQACX8T2zeRTK97tyqUIofEK+U7xa9R/0iatOtEwaGUgkua3fqF0AyRdBql2ao
26wygr1ghIN8iNfZduwWxdY5JhEil4vUfbUplniqmUaSPv3yIJKiEWj8F68x9ZPb
xvBZTUN/gw22ESUJh2nAbZwEQw7ULT8EqKxsvyIns9EgRdKaARhGNwJ88SpAO487
H45N6JlK0uZwQWnHBP8TVemugZqT9MNyszyk6Ce3qio1fkT2Aaj4x8p2wWrqyx9F
Onp/2KzZ5mf1cukOdFq56qb4mqFOHjDLOLMbjhOchIK+qDvmN2L0XpXhHQFL8XvR
6CFH/L09VAMesQIL0he9YWNN9T1kPztpPJBswH4Gz2N80iIdtjWtkPe4KhXznnpK
dWA4KrrBX2i0LYBZOrvg2jV2+IvV/G2vyhy+h9YmGBwn9xI+KsjLoBxKHT04ayjD
44T7aXoAo1Eda9hueFWWSZhEN6tmDgAfnnRCs3eFA+/lvnNJkv/qwuWqcmvyEtlG
ONXRIfzcLU/fHKc7cgYwHTB08CjFQWGypkqtWJzKna+fwsloCgTFP7i8tGPyg1MN
ltbRgaXwlmT7hg0XXE2Xqh1u+Oq+b1vmlj5bihja3DzvsUXgfBBHga9ZWef2QlNt
c71TnkRMsnZAJ880Mq+bk8FB9B7pE2cb9cFt9GPEBlxZoeB3Ff4i6X+hDBRYhDG3
0aEYIgbrw97APOXhHgGEj6ltIe2NRQGSD0gBE1q4idscxnvCWHCiSodCEr7Pdhbv
VGfHXJvRIfnn1kG4E7PxXGg3PSRrUYDwXrY1VQoEJX3eDiQdwAst6ZatC/QFF+GQ
VPxGWYWnsK9e5p2xQVA6MSgp1vutfFsJEqBVMkyBqkzng0pPOUrx/XMr2UW5BAqO
GffFgemTD+0o3BnYT612isBFRxRRc7HqNRMsLOhi1sTVigwawYgciO6q9LwKVUJh
dgJN/Ke+4AE9YPgt8NkCLRuS+cgtm8tF3maLzF434BSNvANxoXxq2zPAaMq49VN1
9Zqc9XYPPyBTjqYaNiSKvSVBcyFyG0hrWoyxNiMmZajkRrXyVlgfaV0yQM/evsQI
YvV9e19SS7DPlk0IOKD7nSYJVuq2ZWJ8HfHt4hLAfPOZgZZuyBzgYhFNbmHbzjsc
5PFtUVT91AboV0VlwafB8g+hDuj9s+Hgx9QLSXNluQo7ZoJnH0PmmnoYyqPUS5L0
lpTCC3XWz6o6RAceDKXxhDbpS08/zMI0B+LVIWB+h5l660+pXWnI2FoI3TRODSqy
iDx4LOlTIuTe+bMznNUy9Dp2h+zJ/xn5WseEq2NL119EJU6QeePEMeYTKE3o2fwI
YRmYqA30LFDivleYuiuImOEPrtSiZBxaBkl72gaWtvop5tYMIZuhYN0u8B/rAxhZ
kFtYBMIyKrwv4hSYgXv/FOWBM9lUU2qvSZXJw9PwLqhai+epBErKsOohZ1Eo1QwD
Rx89lqyADDouTGqf9mylvSwBYjepTWhijTYAzLfbHvCDekvVN/oeeheivCJPj7lc
Y74oLi4UVtGWLPik8sW7CWdJIpNAE2lg3vlP5DjAvBLmnRNdQJAtDykLMe0aUvsB
rTHFpCOcNmqy+FUGPFxxS7DLqyE9FNvIT24EpNEvgznNC4/DvLDmTnvn9TgvCPZ+
8/becEtXM9g17fCIZt8nT75BMveWVstVAaMPJHrNJeJkfgUmZ25xc9utUvm2mVLq
kav8y2/3e9K+vft8nLB5Z6vxG2tctHQNQQWJ80TMhdx7dAH61miasIIjbWLvBmHa
dnHPJmx1TlRVseMHfz231lQBwR3e9dXQcxfF2hrj3WCnRTnydMff3ewEOOBB6YnJ
C85UVKxTZbOUC37rIRewlvE42/6r0oD1XrDWoYJiNBfxOy7xSneajlksuVscfsIl
j4DhsV4SpuXDnl16vQGjuSABnqq7pSaCO15l9xm4skGeUROZ6RqPtnsw3D9NYXaP
2E3UgQcXt3P94fq6zLhkFzkNi9Vb33bipzARtNa/Xdzd8GUejoDihtIBVhNSPRZf
3ij96nYC1PjGGOg19q0uvWeDartiWERApfjZqJROR/75uW58Wrgsv97uqO9qSz5u
UgtaP6azPZdpKWoOsOhYwimtpZx3Nk7RbM71PDkVPmq3iQPeUw+xkSV2dfye+vuA
9XQYmduZjF91gCEQHhpzH+N00O86HkelkazM4eCDapEHMSulgTB/ybKwP6Dvzk8N
tjusJW+EYxw56CFR4k6LTYJVoYzNnN0DQ1EPdFPaNDtjt+WVk1ifnHAenX9tqukm
4WofBYEgvMFpeaY7nK/PH3SAVE/2msqJU8p1/vZf9lrPercus5PT+qhJuc62+FKf
fzdSthSP3L0zrsLtICzR2UyN/GMVtkioF1TKtlCQHZt3Yk4jutaHf9Vc3ZtQYHeF
VBmBv1WCI9NBloN22PG0e8NpgaNM1hxigKYciVc/jmaQVxuCKiU8tQ4NP5hA6Wjk
BkNkyymRmPsO5ToTIoFhsU1B1NNJq6whsCPph63EgR/s513f7gWpGg39+PaH8PXW
LJvdJnESFolb8fAPsBrrmCmIYTm3DI9urknoEws+H+BhVQfqWP27kMBnPrQz5wZx
btsOSWOjsWAdkImywnPyAWUgDpNfpcbiX3gejYofcE0POQpzZ3Y40M2n+8EVQ107
xblky37x4Y0S66GrZ0KxfMwOoOLkkChEnTd+5/dW+TYlWrzXoZtJGZ18C9PTxXMR
ukiMT4E4nlSjlFRZxToJrgO0pjDbB/FvcNBLNrQe7lbZmcFb/W6BPOsFfFAPubWY
tRQtF5MN2QUHDQR3/L50TX+mRkgsVYklHR7oYgCKBBEAsjmTv4zkEwfebGs/a71i
kNIMUkjVbVZ/rSSG0W1MYWVNRrPKw8DNq9w7dtGAdsO0WA/wBDnehcTl7bP7E6LT
Wb2zuOcJg/C9UV7CEgRskd28Kd3XSDBrq2q3PcJeO13Q9sbRGewfwlCUTcndSyPZ
wb/kG0NIp0+91iqQ6eMD2IO/ZuS8g2dHsYVDIwL+N3GdPOc/9b43OomwEs35duix
yljA4ODi/dg/woT6gVXxx0Gl9YX6MeD0P1oyG55S5sdQfqTYChHjXhqyrSNSSpPO
5+x5pHw/lXs8dO79UY+vKTQ5osh7UJZba84NpzbM0vZPdo/zX1MgajHqmHAYeuj0
tI5xmDmFXDcK9fACoxUqTRjZgTtYar8AcGMfEzT2WHWBVBoIv2T+IMzsIUqfgu3J
Go3RvhHrdNi4P7NsAfiVyPwBkpfEqA84DIi4bB54DuTFOh/vS94DElixFiCiJICF
/plp0rjWzFdiH7ZqzDqsOMquEu0tQeoCNIupX881VIkHj3SPszY7GnU2oB5uIImU
57CofW1SLp5ukssTKgpcU9dUspPfjN0P+9zAVyxJlKTlNWD7/aeELPVrcK9tAxG3
LcPkDo01134DUkOowP7MFuRg9Op7AETr3byjf95v4OO0eFwCbeyNKj7EjbO9A1w0
6BfdeoRRdUl6Hpi4m21XwZQfKZziFOp/HA4UI1/16apzwM62jDFeCTNPDwT5zPUg
IcS+3VwDiKYDrfcfTkXvOIuP2WBljEbaWhiY8Iu0OZByUf2hG79Zk1y05Sw77l+V
ECxi0aeq5NvOQMMy86EqHniPRaVqYtNbZ+mhrJV2u3FMdpfVnhGPDASi6Uc07u0Q
cshgtutThx6OjBP61z8RRokIqKlTzB03JhNagPwLoUuvmrTrgmVu3xch8agDMTQ4
xnkwNHt4qMawEkc2bXvCTP0+BS2w7bbv0qGVZJmS89XIyPi7zU8asUHIovALYigb
A+767P/sugJemFE6S/RO0DGeL4+MWxurtYmpEW0p2zdUj6vbZ6d67Tjej2NptpAi
Lwpxnb3iva9sb/quOYyoWtm43xwhBYdb8ExjfRUWKBlWiMk2EyYc5mW7yvDMItcc
Kg7M5NZgf6rcdkC7QN05HRfF/A6wjX/luZoYoR7L/hmDsLuiGrnOVFntSbtTzoL4
Jl3KavWXJr8kZIyvmkBZMNkpTDC34gm7KlQqIB0AoKAaBoCVhOZg/NQLJmOgSBFn
4uzPUfhs5AFoxLTP3BeDZDL25njU6krW/sL/heTKrPZUR5yFmdvkfxlowoau25ch
g1bSqztUTi7S5s78CtfoVlhaxj/9TmEdGCFotH6RkOdKFN64zblvhAml9G+1qvtZ
H/p0jeHPFDbOddRGpkPPWBpUCwkOGReS3LcDikzJdzPc2vKatw12/PIz0DDiokBf
kaSmPDKX4WLTICpq7vUzusB0GAORtVsg2Mrp/zNTUaxv5VdRJ5zK9Xet6mEL1KVd
iltd07Pu8LK57rxV+4sPVX+rsPHTNY2d8mZzhUVOgdgZVIslHBuNtUxAXXlDs+aA
Ur39i0RfTZqV79fO0ceaS+r3S7mhtziHUF6Nc/dalkCB8rNha9yUGzVfvF0eFSHG
9aPh1CO68KLlmA9HKApGox5Ntp/SksZDkllm9Kt8UpJAMh1zLu5jpEMRIW6fBC8j
c34x7adQXYhESqLLKsXvA/q2EriX6KhEGHR2FKgpsTMcyOHQXCSlzzex9vlXc1mx
sHTOlkmV5cUk259hZZtSYSCtt5STNgjN9IgGyiH3XzoazOrbRVTEnl39wGFDOfLH
VoIXvqHsV9LEDRlmiTLUV5seUE2Rz0i7rb/KIjNfkGXMKX7/ZtZl5hifV9hIEtmd
1iI78g3LgHD+m1vlf8BaMYjWqZqikkTvalPkDeUuRNPI72rgm5W1Zqds/bsmd+Pa
/VYjRMLsWciiNLUxprEsoIvDi7Ce1b46Pex2MSros6WmC0khGxtuVlGSzQ1bJcqP
K5cVFnFzg349ggw/Mbxd7MUgYboiHpwMsbI96fOIgnSZbhPF+bP6aNS5C8u0314l
/vh49kAN7U/uQrAnT9L1uxsyt8c/uvXcWRAXuETjw/cvJOsBebB0aR1Jtb4PiRrb
Vz31D+ZxYLQlO9WkNfMY9Pn2jw2OSBchIjSueRi9rDBCny11aYWQUxAx6lckqQ8J
OW0xu+j76BO6kD76uB0d6X+Mn8bJsIpJ7/Ayx5n0ycXSsDcffKy/pbiku2sppHIi
sIeCOXWqlcbmoEIr9ljbraJic/tulpZK9Jidm/OfnrmkUnAzyG1/shWnFpWhwDWr
E7KIAeXkdD5B+i+Mgy/tR42B7FHdR/ikAl6EWQywwvdg/Xi5KNdeeLiTlpnYuAiI
O4VXrvnrnAOzkwiWRcWjKC60EQvZOoQpUhUtTNygmSEPjVKjMJBFun1WekR51fKn
HOCjQV/i0Ok33tJEic2vKHM65It2m6TEV3M9IJbVzBucNuydJCq+x7Rx5fjn7I+/
6VKTf62dAGdaSpF2chQR+KuIPIgA8ajV0sT9Aex4v6g07BhoUsXoxSXA8MShXg94
YsN88MJ3OrUkL+M6VMX0xj3STOJRyA9+nmyqY1cs9C5Y4bC7XHA3YFsaNi0tgz07
/32flcjXmjNjCeqGKp99xxYCaNWpw9FbnvBEaF6iySVLg3j4Y7/teKBObWo4YREO
PRTMdPrneA87RxXb98rAnsM9272G+biDzNURS/fI1eZ7YhWyICwGN8CRft0oG8SE
74lF0gYRKKPXSr90/q/jV7VgbASXk+dei6TgM68zkcEIOightTgjyo+W3MlGW+jy
QCu15gGwnj9eohGXknaktLbIECukngyrQDV+lQrLysuGvDcMWFDN6Y3biBN7uTre
ByW6ObZ5vIsBxLhpXnrk5Rtw64N1rNI/LIc+PRL04DTksherFXghP8lZFNQUFwe+
6kaT3gE6bRgVLfR3fUkUZnDm9vk9qVDY5nvdqBaiWhnczxBk0ANEuPHS+V+oBMT0
J35x4mJX8F/Ggb7NYk7mb6eihGpBd4mxUCOv/9ILuGA2hGUls+9VxYfzQyLeVSQQ
F22BPDcvQ/rTfMltTUh2EQsxRVwiDEKGjx9sAHYJs0U06g92t+LE8E+/DsV7ExAH
0UBJx36AWKJc4SN2TH5gujTaGDKVdBLEvH8CHAUiZJPD6m+4lCv9wgCfPa5jwAVA
5p970PbiqTKVX1Y2FjWv1kJ2USSEiMy0oFD0wMpe2dTuZquHhXfGdhKXxqz6B56g
Yj0uUqZGXscI17YSAKCFTvp/tG0v1QGQighlNv0opTwG7lHD1SVxclvLP9vuheul
mK4jhAsLenHPCPq8XtrcEvXwh3PU7P1uDRPoOqjKqSlc1VuF0R5WAA2fzP57xRw4
ISkmWDkUEhXhvqJpQZB+DaRRN0WXl0d30HqL0+/QbZ+AEAOj9LHgWEoZD8mfS0vF
T0EoYS93QPmy009N/SDT6NgTot7vJK8vAPCtDEWaKOgMhw4Sn5j7rhvAsmdP5HdF
8Gm5npXyykonahOCheulPXbNqRCi3gIdjjPVyNGTDZ5K2iOfr6DqL3PUqeEwjkVu
vjBFUvQHeJVBt44H5iSa0L6x6KT7JZlWrgttIJr9OhlaxRkKm+K8Pz/nNP6MvzR1
4GyQrIm8XfSKiJNJ8U81wTXvAIbEK/4ojQqKxCze+4ZRlg3vieGYUrC/CfN+s55N
uTXPC2gsE8mcjyHebm6t5xGM93XWpL1alRBd/Fqgg4KL3yI16Sj/6fXDfL5+i5jo
xYCjdCJjcyVnfJ17KSRD2beiJevhTF3k22khwJ9lwsQvSWiIutotoHWU0ZKIWpxv
KqY3BYXe2aP9w8ba6zsB+qSj/23RkqnP1tr/5mxd0VSTIr2kU3DugF6XFf0bv69y
BlE+wH+OtGCLScC/8QHODE6a8GD7FySzakcJ/lbIj8d3eChNQ89jhdFF3zg5Ussf
HlsBSp7SzJVYtHBAsGZ12GbPzwZT1/VmXIv44q10GB2imgBRues/TvHgX1d8e0EN
DaxWRjEAOG8cNS/y/jHov20aVw2fXXt7Ea874TltlkXnwL0zZvLKPwmyRlb0Psuj
ro+3QWhmGWTuBUfmQYWBtPX1yNZHU5dMqS7XDAHsE4ORiRTsbtj0xN9JbQBh72mB
pO31Tc06tB8AKTH09aBhM0yEWR1IRwWa5N1yzEKntIr9nPzQ9xqrdFrJb1UlBnRW
xaYx/kvRKFJLGSvC2m2Rdt9dITNJHf/NACtASzf613HnJ8ItqHHVQ7em+42bacRd
Mp5be2TOTJ6yZhHknGsMb2gaWj0EltzFoBrqeuHdj6sC8Og6qTiYSnPod0bGXnOU
4Y2m2y5MEoRF5ww37nY8A7pUhVujbaorszJBxU+xv1W2YXl+SpQSupu5zg7nHoPU
zjjUi2r9HY/WaWjptiNgMKMqbPcdYqEzcZEJ+oRi/yQdhWXjNoxF580ye4xsz8Q5
6kKbs72IeJCP7jvDnlke0Yvr+RtaRWLWdR0oTtZ9SSynoYS6fMKqVplEnUCSaShX
v4FbS9O7JpAjzCuY8PKoNwtTMbbWqrXJQi+k+TbkesLyCztPTIXTaZUBQ7HGc8GA
MUOMf7V14jNvlTIp7cYJUEKxdbn8A8YZ5YsHIpca3RiSuClobhvjX2NWXioVy2sC
PHwMcR8BNiOz2dYT3BVemkqBqwNgaEkU1M2GzTwgusRQt5r+yaphv2DBaQoW+NqD
VoJzkpx92J7caLWyob2144YfpKWm1qwQsfmbWEdAUSx7o09JS5NKcTYOU0OEsWAQ
MNJ9gF06n6jcNLc2rkXzO1C6Fso/k2RivDi4cA7H63yNniFkr4I34h7nOTCkb6pW
gYoCSUlN3M63BRchLbLb4CGFUzS5/9MUDUzZfqXrhEif8MvFBHYiWGM2w/SsXO3s
8j2lHoOZgD1hHXVU04OfwFtYERLLgkd27zfSNhGfwrvUHx6WwMAn2fF0OuNQWaQN
vFTvNH4TFzMAPnPeRikD8SzuhXaPXRCGv9W4JJIESJ/KbaBssbjs8RKA1sH3/Sqx
x94tCAD5mcrkeljANQsGuWTeh687GlOAqHtZoapJxyF6yRViNbX6BXKSuf/ZQIdn
U3LISRhHB8yYT2GrWF2rEL916NVJVfcbDs2i4qTYUXluONzB2hp4sMKi5rc8Oclb
gL4GnwyHbt8i5o201oshuNze8eGe6XA5z9s6zmFRwXbnSwadTfsdDK15sH4fp37T
VHoBlMA3+dxUBZVkZ9jCJ8rkKzLN8QeJ384D+oMsNWotXRSfFYwAIjePPBGrP1OU
AzIje5YTsLBWLQae9pZ0gl0uTCDMKlEd97sAH/plFPli8GvURvMHuYd/92Cugw3C
+NniTD2yC4Ns6FR1NkhPRtozDXy5UFAd4oMip3xk1otLk6y182uwni9JbNqxoEai
sNWDQrrgHScDvGvwLb0Zo9kRwk/vuqS+1JeKazAyKiRndzNkcXF6CvyYjW1F4lQk
wEyOmOIn+9PUVwNDFJQRb3p/yKYvFEwU152e/sxs8x95z+viH42bzHH2Pdt1t2yr
n+dvhuJ0BdBuAC8FA4TA4CCeeOjPxgQ8x3eqi3FhkYjY6gAilXciHBhTFlp7oDIS
r9mTpfRn5aU5NTe+QLJbX17iBV5wSeelo/lB9XWuxZzFkeWCHcEzO0eIqd/Ir13k
K2KMnStLE/60hbeSKXVG/7kiZzmgzhbetG1IFESFqey6jorJ3W3q/wZo/KipQUdO
04o/rDBj0+LFRgNZbvSW95oERWE8vP/KTfsidtKxzESqlOzW23uQcpwnBTGxsBcj
BDR7UOjeeR2kXbD/+tqnyXRzp5qSSjxeAr46vk3tufa9uBYl1YFclDLIbJU1hm1z
aQgjSQdkJ81fCo8+FV4bpj119QYPefI/NHdUush1GfVx/xJ6xqA+PPzQTeI5peFY
rrrBPpVTDIoWf57EbYaauBDN9xUTuI38TKF2LPTPHIxSF2zDqXU5wfnkfPpe58sq
+xZh6KxZG4HICINSMhI8i+trBS2WxpDdJ9a8KpAttTEFiJiWCtKlqn+P8euVsx2Z
si0oII8m3aqi4qeAgJvy9i/6hHLUqDbj8Yoom0XfO9MhngfsWu0Tv0zVdx1UBN/w
+R6M9Qfw3uh31yO/JNGI6lb+XitVbayKBSNYMABkIKhoTmXLXkrgzKx/y5kBlEIL
he8d6tndG/GYqn8Yqx1VQ5INe9TOBq33yFMnSITaGYpdMB7BaESytqh4MrIoZQDm
QE6KC+8GT/k9kNf6pTFed24RkK9EKj3Me7CNLBhXYfzMOuQaI5XpJFQxy+VH+rrG
5iDzNLaEHXUZuooYwGqN2lqN1xvrilroMahDQcUpOuQ+PktDok8iQ5PQ7YjbdRwA
NiEtVGTMu5C9soWPu3RaZ6td4IvEH2rAHEtE0LNPxcYWyXo37QsuNd/DT6uVDScn
lwT7dxTRpaYY5IrBW7X128VhEEC5uxzrBxNqzPCKug5hpFkd1QwzUcba7Ma6qMyZ
A7ClrlF1pJv58WvfoxG2bibmjNXL/0kbqjzBrB/H61faIhHnO9fBZRm8UBmLwLEy
MIPPwaepkBgcvwsOucyctS9dUVQHf4b0yK0Y+GmHGb2i3/z7m5LfqkZUcRenErC0
9pSkxlJDEDJiPppsVkP2ZeBcjOtvvoAFaMSyClYG6abdDBHMsx35F1EJt5LnZwzv
LzMW1BLDpY57/L9xz+F08YrbBtFDALzP+1hoc2YX30+ZzPmXgKdsYqWR8/W+4p13
V2ynQfK4CBID2kJNHuCpkSPz8aAgAuQKqW0LThBUEKBG2P4wLD1J/QH4WHosgN2C
oHICKqut1WmU5Bh8zNj2XE1khsfNvp0WnX5+CvWRscW4jStON7Jm1aMr5jqzgiZM
FnYmVEi0V/t4R+iRMQe39P1tpbOb52v+rWOMXxMTI3wBYHq4wGcndoyrIoCoKu+3
JqBS1GN2RWAULk6dt80dxXRDn0WRtww9kOyaAFhT6l99jIo8vkvU+1FvEf7VyyZo
Zm3AvxFpu1LBTaxkD6v2VCP1RgpNmWfNjrw7UQ/1TUMLRad4dUAwLe0q7gg0wGWQ
zzLKMhpWhZI8eaAMtJzo/UMrgsu0lOf5FXNRnmf07ZM5JUAGOJ3Uif39kJKgyxMl
DIGZb47M+IFOUlcHwuEGYOCfleKHLRpvHXQgSBBP13R0l+E7j3YUTaKCszqTl58r
Ybbpo8xZ4MmQMwYnk1WidKqYZ7t27bQ74K1NT1xErKJx+sBiI7uapAgbJ/Wl73rl
5BE9t25/wSt3NL0MYR1+WLWwGR4UuUBVOCyvtRoVCl5mSsK4vwN+n8wZW2W4J5AW
TMklBLZYZyqzuVrFE/D9mSZGR1ktIdnABkqrr4gAevy3tnWl44FE3QflfVltf9ZJ
lR6JRIEkCh/ZVMXODu/5ufZHyafvBIjS0iOou12HmlrjyfZ8r3AcnxPXeSH6rnGm
HVfkmhZnAXwlwiQSafGCihry9wk8zLaa4uULnIO6ZtfoBqq6yHdaRbsZ5X3/pUfr
G8XEkGEZEcrTFghjDBfcT9uZq5nq0XeFMKXY3TXZaj6LCaN27KXYeRgXfNpAyENN
f3B5iPUtgMObUImWFhd6QjQIyrLz+lyr4JfR8jRHmmcNCD/+2/G+yre80QhS5L6J
o0vdRApcUWbV+k8RSn78el3rsYAwUkg951bxElgV9FifA5UbEMBZjfxwygYMtsqG
UhIK7U2LkzZkRpdVlwYk2K2tQqj0Mhvr/iUV5meTDWXxMJlYGgnLZYX4snJAWJuP
ThK2BslIgew0TR1Z842VyTTPxgHUuobE6+wgwRHTdUVIRSk+GrJkHVTPq4txWAnr
XIIcmGbFsOJhbc9WUbsuUz6p2TEU9pH3bmAgv+6gNVLpoFqGYY5C7iSkZas9JkKf
WOhqKlFh41Ipag9+b+AdNFrId1RPMMU7papokNKFL+EPxG3MoM+6aC5z70r1hLFx
WviMk7Yd6gNVGzFZAbg2jtnO3uwZXq6PuU5toyltusHjFwcvsxkxWOB0FsViZrzp
37H4P4i9vBZ/wZNm657UneLuBZVLbDFoxmq01tZnT/fZQoXf3I6tX3FE27vds96s
LcjoZye0iEwC7V/6mwa960axruzWAfYM2uIpUx7kJWbc5S+g12y4RAQUpQgCKIgt
sUE2LPk20q5YS3oljy8oSH6nCOZwM6whkarEWorxjx0D4S09tWgyPzGEGel0dL7Q
rPMjQefa/93ZQoeNr8PEICUSWIgiMxGwRxvggKk1UL7NpPeKzzP/fNjx+ZjYIez2
fjIYsHLNvaAeeephueTYvqitkvbHB4tLER538MzYYTvkbNfGHLocSC3OtJj022ni
uf/6v3+/p+KZQEWUrg+Dz42uuQk97nQ5FUbesvHgn8VMpTFtfZjYoB8qDqFC9ftQ
EpmgT86sI9Cbm3+ppswemTKFToZwX1G9AeYFBtTx2PyN006hOJMSuBpdHXBIPJOQ
B8Dh8+xAC8XgO6Ig13qIZF1bcyIBmCZiz100jlECTezAa4Z2eySRb+nIovE3BwMX
uxGhRFl5Ya0qo7s/b/7bFX3iLv3taHC8pXEChh5QYOayyobVmaNFmZKZd1rvWO7Y
VijSkaka4ud2OKERVKfoztmZjO50moIoskJYrGdb6hXLVkokHBdHHqjaATUpaCyf
W3ZX57E9LAO24HXVRTggWIfsMLd4Mgc+Z4Gap5p4bvsaMD0H56011OdIFo6nlHwV
B9F5Ko4d0HmAd38MaqWkPS7KZY1YoilsE22pQuSHsrob6fq40x91h8LrTD+ERjHy
kpfYRyk8fq6HxSPKY09X8gKUiAeLPNOhaWyPCiAyBbaSoZ8+M44WWQ73QdhxH1ci
RW1kTHigV4orTdBIK9IY5UiGgOmtANRU19SoPJ4KQZbuowiQFCe/U2cwW2wH0tpx
XJmoLB9A6mkj9LKCS6n6+0ysaSXWDtaWG0jdASwAKZ132G15uTB0yyh8gKieFOKK
cpYp/VQLxSDW3+a+69fZFbFN3JntHUcUywKGqu+eX1qpGi06G+jmlvDH4D49aezR
B06QokYsYQXxccAlG2ocCwvLf5TSlE9BVyl9RFRwEcbkI5Zy1PFWdJaea/5l1b15
DWA2FjozEqK3lJQ901gPxuQgFOLiz+UTtewMuuYxeSPFGpMfzSQguY9GFFoqC9do
xsDHUSOY6gPbh2VIjgixKfXRcIGP7m5j0OnwEccXidiDhoav2CUgobRFjHCFoDfE
XzNI0hZgvlQUhlg/yJ1ffKq/5LPkb2ZVQiLZWmDgb3L43wNLO9i0PTdHGVq3iMxf
pLXU+ed1j9WhFPxDBvYiqPc78j55r4s6hVkImfwRdeYN0SKelGFNS/t84ddyKF1N
YqcA38zI9biRaNK80hRiztLr2xdarPLPqrNCqCAYh1mzTju/zZssD+2Gk1GOOfBz
FCdQZcbWnJ7lIxWMRxlRFZOuDyPmqF6wtc8PCAAJkVNuXK6QxJsbmqRAVrcclR2c
1ml1rpcbWO7bEJdVLEssggeE7usg5q/p3M6fBcMtpMavwcx/9VOLdQZQqSjk8Q6x
ChxNgC0muGAw2zYpDRX3cKL7OrSdxoDn5qgKQamL3djXbpwGTu6nIepILzTzD/Jn
j9roM9wtitGnOEFDkw/TsEE/y9jtEoRzpK2E4cpYSWQMI7+n7mq9VK/VDzssYI3e
YLH8wkII3eJzUWaKk559kLWQtRwKRVKUw7c2W7SC7jeKCC13J6bMuvl6Y+wxg1ad
l/tvagTdNoe3X17TlsfD3vw2st18CDD00cksH1boYy04yg8Phe+Wo7YRoc0Moh5g
RJLn1M/pUivhM2RUrpj27UL2Vo6+G79HXy7Wp7q1f+e8lZpJjIdqoIT0Y/JgcIXP
p8EFn32qdAqbleapVo9jg5zmwRdd/7rQB5f6z88TPoWuUzNz7lJMlXsTLF9I2kna
bKoBiL7Ua0l7PeVLgzRlZdFvt2pjLEmssnQFyPQ2Kpu42+TW8+EYabErDN57rE4y
XKq9fUgSRrgDac/gHnqKcx1WTNl6Xz2HVevpq7q4BlOa2kStnP+aH4yv2bAM5KLp
wph+f4E7IpMj+4+5Wj5YYKgXXWtJxLdCqaG+NQqjKmds1ya3WPADtQRb8Ceatedv
kYZ+K5xouXKXXLNVoOGVlCuTbchleORi3c6jsLXh4+Z3TXr+KC5+1u9fPxZV2nig
VQWPQ3ASPHcID1sznwAjaE42IQilRWC1/rZ3OVwZvdLb4rtL9jCRnha0jQeBjVEv
DWj997M7Oa/mvYG005wmCKseVop6UWWZiJ4Ehh3caj3Ky2RZJQ6OHgPK9KFKgvlN
yXtAKYG3PMbR4jq/0+cJAmC3HT4Jy0EQLl/h0h+goG1KxWtJguI67pUau59y5EEe
QwD4P2GIJq5sevaAKigGtkQlpq3bfPcSLWAN4G/POzhf7Co+Hghbc9Y9Hn0of2oN
MMi1QhusW0lSuw7Bw9eq7sJ6wJvjflqp5IQxLInj31RGD5XR7r10KP8KbNK/0PBm
go2sbcicM18I793+OoQMAEbk2t0qZQW63RXm2SKYxEgoPP2SsTkWWSbmpRbyYPEB
VzdLFmS6ICiOE1O/frv5r0fvuLyMHUZMaSpl9gBeEImXxem4VVKke7mEJ0FrUm3W
HBmMQNkjWlVDxFvBlZGuEYsaGnrke8HP4zhFuE3gyRiGKAtZ/HEfvh4xu3g3tcCI
Mot0u8/+0P2ImHIrF6QwQNbhnj3T4YWzjZ8kUtLuTaoG6gEvQzOY2I9r+lGXxgro
oQIc/L2UZ+HaaxSlR0BUoWtWA8qDCiuh6HHzzWt/98bgM4gqBe1PXh6KILIUfdVt
3lYDzr1PIHOgSXkilmRBa0HXCHX54XS3PdT+DWdlO01y2bBS0y019jAphtf3hRqX
Rj116w2GaGYnkSc92EU9/qFcqcgj/AP7RuYOhDutFoVBuM2OwtigDL+HOOfnaTS0
74h6EH/D7wIvzqbb5Ervrw3HxkUWPwpwFrt/05pYY6T5feNaZ6XWgX2goKFcgxqs
cdgnhgDC28XrBHhX1Zz2qvDSR6GKflID4lIi14WI+gbxnKsJi87CMd6Hud2AgKzW
GKZuQxLxibuXHoaOYRFmOSc4AZWgyRjhO35E5up/f3UNYE3iNGRVbBVtrYXCStGi
KQOp1tDMXJq1PNXLpmN902zp8l4VXyBrg9Fi4STaBk7il38L7TI7V4dDF1dzq4r+
+Cy65CjyyV+OG6ciED+EfiKxuUmE0jk5CP7qk8np6kSscPUCT0hUx5y2Bw62Hm+A
r5TWqMjq6svvGI1c8cL8yQP8/Uimn5AUaldCb/FWBrjqb3ZFKvfTYX582Dq5Tosk
8jxvuecvlIj9jnecVS5XDqA0h8AOKg4RxXkAiNEz4Os8SFWVyOpStYhK9ConFezd
7tPAi2v8/tMRVQBJcsdlss5ulL18vsU4rdx1ZxEsfakNrQj3mNk2B16lly3JRqRI
Zqq8MY3FyOSLmxoKlphA2Q04i9MMkcr/UgZZ4oZqCxRmTpLJiz8Mvo0sqPFfFmBI
FCMXwW+wGcQmFnaejxKJ7rRhZqBraYC/Gi9obyLVD0HtDj/652gMHijLN5dCrThp
NsyHBCwZVycB5aSUGGl5m0643oe8V2Paz6J32F5skLunWhAupJqnArUBZPX5ehfn
3wsejJIo7yoQYQUJDhq8lXvei6MfG0S0KWHy4Yn6Yyj51Pbg6t086P0PhKITgUEe
ylRoPQnYC4oGNnjgmQlvpmpFdEhUXKrvmLJ6QZdBnOyFOq5UBGNt4dOdcTrJI+SF
SIi3BJ3dDQN+affMgE7OUt/63GkaW5NFbAnGe2TE16sX9SUlw2YFx4fCzdH7Fsm4
Wr32503Qfbg2ql1c4jgMZ1FmEQ0GXNGo8doGRE0d0q7f8av2YI8z2T+ENClZX4NS
46ORaoDuqWMX5NFHVtcE4d2H49ZMmok1z0RLMv+6k53/L4L3VHUlL3BwcqNSvNRj
MkG/AAFgpt0l/NCRwftL6drEU09OcWEnCBTO/c2rDGXbrQVTdLofWuUE1HsGH1rG
ajEXA0j+fqa+xSfSN7TifTr/HjACB0kwid70VTuTLgNJ6M0Z1Y++C/cREGEJqKsV
Vi0Q3i+WlphcXN3AIJiOl/+eXyxBVmy/svjItT1PNQxO9p0C28MS1QsDc3xF3euo
WGs3xuH6sswwy77bL8NW7Amjwb40wC/3xlFvs0EpgMXF+0RyrRHL4x0MGapPLHFA
4ceftDzx8ozM8gPEC1aPBO+vmYXfyG2xyIo3Yt9+dLKJdyOJpt7oASa5j7fHGmls
nEJ+2ftcbHP8iGae4+8QB/A3rAY+motrAeKLuycrtxzjGQnay+0QAOU/CL7UBPWO
DcKToD84f5rsFhvw8CZ+rbeGU8GreiZUl8Hm8vLZBulp75E9FZ74Dka4NR0Bf4Kg
DYglPae9dg+pqv4rmLZODzckH5F2tQtZPXvD/5cQoHak+PXG5HyHxYPEJeNmhYl1
n+GOO1Deij/sSyuRTGB+HwG6IYQXo1Pgrv1cByLYj2L/o/Iwh8HCQWGmx22OssOa
QX1uqEj+hK+PYM9ACRRZgyNbz0ClzFK9cJqeMGxRgiK+AJFZ2Qhit2zxv9M7kfwS
Fx310JSqK0Em7xepKv2GrV0HFRCwwAlsLH8nUCX3eJPUzRw0wSB/kRHXWiss2o9l
hWiPBinWnSbjMCrcyIjGzfO+2JQplYBXnM1LeuvIC9Nunrd6vugwyqpKukShvw9/
p/hMdVEdhSHf4zEoz4FCHddDVWdBIE6k5aS5A4Am47qvheV4aaNlg4cjmDUz13ER
lJ25r2CJVMuldYSDyNTn8FyfcYBGAaFCGc/EEWan6u4H08RBJ18ByueYLXlvepQw
2o2HqDAAAmxdFzxLct/oX6HB54Mm77LRsB62IvRpaeHHo/Ep8kVcmh1Dn0cjKmMB
fj7wETJ84THfc9s4uWgh72CJtQzB2FK/Qj57a1BYhkpHBuc+Yz7mEP2pigTaaQAU
3S0+qrNOHYmR3oJX7JMKBRtnrylRmxyR3W4Q+JuhewbeS2iVCbTRhdqZcxrRvS42
rbtc+QHxzO5/fhTAIX+2P8scyAa3yNU3y4zgwpHu1lf1pPZEG3QUQ3CCx7a+CJSA
PSeXEJ1Rwyp+CJ/oRaC3DovhY7Ux+YJf425jMAZ8Ytq0XImeY+uVPYIeLhSU9GAk
PnwvGyBuUt7q/Bonoo1emj6UFk5/kqhbOgcNMc94k+wPIT/UnXmEYQHTPPTemoiU
cHvCJP20Xyq9XsI6G9qss5pKlDvNyjXVkPvFI1folpeltgNfFu4riMwkklKM3ufy
EqmuYcK2Rojx4Pq087Mu5+sGjoR+Cvf1/VsGt6keuUxWLO1dqvxEyCjD/i9MAMMN
dbhpAHY/Llw9fNECoi6VFhzjlcfKl6XOmvDE0XzHDzFBJtN3t72v92WLTcyEhmpx
gkaCBgMkvRRtXdKnPKUtjkBgvS+vYsuqMXleMnuZiqFNvmq3mg3fPEuAAOmMNsDJ
dVcDgQ6aT4t0proCYPqtMHLeB9nzHZzcwt575AUm8gJdFgidHHZb/ocu4Tv+6lJb
aTirIxAuz2mqscpvZkSktEP8O5woCGEn2I0gBBF2x7cEe/ngzVs0tb9GYPLKouXP
snMZjLVpV/t1Nz9mQln1i7At6KV2WpL7HB/SWsmVBF3vHgqR0SxueuV5dmzZvq/Q
O43c2lM+ILT8bR9t5yuYNoXaaYlEaCsna2Pmv8YS5cCWCSoS7E++scR4n2OMjcUR
wa2XUwoqDQcDIpax0HTr7FgN8w8zBunrtpQnWT/yQsGxAaIGsgVyqhO2TI07pdjR
LmT1o+mhfg4lGcqpZL0Uhhh7ei6/1nzlymX8bWa8H24yO7fKZG/FJTYr7jCpKqzG
ynTQbPKCfBQsG+iw2Qtwm/V+CqvWaPNCUuH9D72uu1X5OvUYQriQahc+pcWAyDKp
fgfme8PqSLt4k/bQ24KbzX0Nqq8zKRoO8tzpQTtE06Mc5L3fEisyuL0SD3WDTV2y
9cO6zFIXmcRkes8h7VMyCTBw5a3Kbh2LEeF0igX07VuYyfGt4T2dYRQIGm3tVPqh
XFy1TqmcuiFB1nNSVNwbPWozHqhm0kmbwgH+mWvIB4J1MtEDGJw79Ht+McQa5Ndr
0xZLdh/PfM4D84rX0tuS7vibDWBbq4COmpfnxTUF1ijgruTdIkj1fMghq/dpHEY3
ZGSnONwco4GT264Ef/gNEIt6q+uJRPb7sidroh7Ua8XVQ5vn7earMA6wILuec0QF
INzPot/1+scZ2T5hT0kHYKsyezYoMkxzxY2UK7kzt/DG9Sfs/7Cg2HHMQpueeh8u
jxKYxGNFDvLSHljrmu256BXGBeNXpjDNie6rtfdi1Q6NpyaA63TKmxbi0Bdyx6Yn
n0ZK1lqmstTbWaRHFRIN0QBKWFOm3q1ddorIsE77W0B6a7X41rKbELJ2uF0W0sUn
tSxuGx79UTorGBvoDVlRF/Mgw0piCIf7F6RaW9QTxW50cYWr3t245Ej/a6+t5MYq
qhlQNowBMqkDhMsae+fH31f5MlOHjrkxCsrtaypCYfAkZP4UTMhsdCI+GMma/RWX
7/8G/0zFJR/QwlNFLq5gxLgzEmLnxzAK0AI4ZFHeg5Dpemt/d8GTiGjGHKQ62D9s
RSRb2OTcpgpF0440BpMhHa7+zqtqJH6OQhMKLJDLwtl8XNsbSthp8QO8NugY2hPt
Y53LV+g42ZDgqnr6HzFobJceOZb793QaKBaQ/ICl98fl6T5Fk6FvkzUn+0297XtN
rQfXqpsSy6o7gH61AKCrT79kuGbUk3sbPjSeN3tx4Wz5vCK9bN3kE11BtIkTCC/6
OdVT9hIZg7a+4GzMOYrd3QSw66mtnBMI/rjbq6EmfQsNJu41Zo5lFjbHF1EleisF
q9MJhVHnPFET/b4bikLWdao11keRefmEkXMhZgs6zKS12/Ah3rp+sxLpF+qZtpfv
Z1ILe9qFctua3uHXl2MDdFH/z8HysqPD0J0Arl1dYIcabUdMjkU6jKMoDQzyKH3O
4VpNziG7/dLj8v1yAhOEFDtoR458FT+oqG50flyG6IaGc0vjG9bPeqFzd2WQHWPJ
AW4vgzR1uUu0TwiL8noXYjx2uYwyE3yh7CnNLAS+0D17Peluo+vnU18ql9XP2CRv
6gxaibSUefujKPF4V5XX8D2uqa+sOfNlkqmu+YVta2vhwfMOFcF7hDDOVr31DnXe
1KEdBY9cvH+zmGtna+epzkQUYFIRgwUvDG7x22rH5nf9jjFb+pitNBS7t8FrezwI
zztOSsCP0eLbvYrkpmfq4uJMzi88r+tpYJDtp2UiYKsexVDxxeI+SvpJG7NH4lup
Dv3awOb+PdrxKjahqPqZkGpa4AcIX3TH5iPy1zjWDY2EU1My3aOx8pweQRcyZt3r
Ydf9mKb4g6kdjl+QA//lU2iivF5pY9WCRSUhgowxQEZTZZ+ueBf6nxcgnFsxCqln
+7nCkC/uYuhdP2chD63FWO3gfy+/wGFXtS3g9Ct8Au7IBxaASlrW1CGfBAcLJR7Y
ueJ+zpqYgw4jbTCBR/MuOWgIrwf/hp7LSSKsznvDa7gm7Q07yWAQ3Uui/lcPGyb/
ILhaH+sTbFtl+oJyufd4ljNjxooZzzoc0BHD6VPJ0uhFW575xQoGhGs5ZUASG4k6
yeZ1Fh2wvXDIzJ3rqkOLCH3yT3I2djnoJ435oGMmILJBC2B3hmHemJvDMprXDIax
YnkJIeZZHW2Naz3VKqbKjRh5YNnfJFEXr7dM+DHrQpgdlxx9PsbiAUkxXCJF2jeW
pzs0eA/OnD+EQglfOt496Yv9jrnDyR2TGX3SbJED9rCRnHwwTJYajMY1TeQw27KW
aiIGxO2guGkEbEXxOVRZ8Ok4Ozn+H6bZ+MV0PyAotahUo394smIAuKPY1ix0tENf
CIoUZme7wtRupjrBpKyqxirVEGcBDSH0oG7Ff6buCilY/HlXlUGU4JJAdM0ZG4iW
nW/2iLnGeEHaRqjZlyDukMxf9Wri/nYDmVB1b2Sv2PH/aFlgCEBZCP4Gugt6pOTu
vFsyHe0ahKBMzkNROWS0QrVYhqTuOqe85g53fDikxZfqVZ9gn5vvcH/m4rEsG7Za
lwpsdNKkEhAQ6nEhWhaqOEqXq7IWJSD43M7L3Jo51H1juuepuroKhOU+/ANLi4yf
+noONZFME1QWCrF6jhtl2dKT5ZKb/4DXHoeqcx7EkV2O3Z4Cgyi+KpR2bOnqaHdN
guoOj85eYZ+d8TSC+CmfX9jjHAOIl2om6H/LB+LIahuxZxtR0En0u+npf5P+8czd
6CGQ8dAiG1CYkr/PJsklOKiAsK8sNlE0bTlFNH3lNs05aFlGHh8Z3sg9c7pWKqrn
uBOT2eA4E+qTY6PvdbUEqHWceCBWtibjiVNzWy3C6ZXzB08x0TCdp1ChV4n2A4Qk
RLQC8K8iHHLh7RLy7JncAnJQ12aKbm8VhZmq/W/odTb/PsgA2TbyfiMBZhoZuDyj
A/JaLSiJHW9ipR9f5/DTC/77aVbKlLl0ivYKMqWXfUk/AGQxj0HJuvlIsN704++a
U3wyBfp9qIOs9Es2ADYHr0R9qH0SN4lYZmWF2IkWxBocaz+5AN485Iwxro+fCAVS
65PtMpfOG4DdVAGChUMZ5HVvdtd1yehgdzMu8rmCycdgPWDe7AHLNvMtvwB9iiJp
l1fz9+/wnS3g+UOs5feffl3LttplJJyiW3Xk5nposit7u8Cf9JVz0BplfFm8w+Dj
+E6/mw2mQMsWbc60tRw8lJZAef45khTXwDfkr7dhS+PEM4AftBiVp3lGRF91X88W
OIPJjrNwVBXIqGTsF3ZTKzitV2nReQikd4XJYwkxFQFUcMVM2kv8HtXV3akh0NG8
Rp0sufPuXEp2Q20Kv/N4CQqfXRy0obeNWNYxuy+meO+Fxt5XhTIG7xvhhnR9BhJY
NFLSjRQZu1DYlr1SCDrixatpfXwdKR8/E3kSC90dxfBsp4Ch+JW1j3kEf3qB7x4R
AI4A2yraci48a89h8tqE/tNReNK62e03G9a9SCg/kaKOu5qAfEB/z5iWINtuD6B+
NX6JhaqOWqIxpxYTefMSaFCLOc5Eo0YOGjitXQ4lHfRuItYDHKp3flgk/Ynuedxr
+E84mX8umllAwEdi9yLXG7PCXMBs5/cHxj6rrfqSsdbmmlmOuTFMZ12Yu9Kz+ebV
XRJdIdxJEtYomjHZhC1Zod4hyjBXV1O/+wLCQszY7RkYyIgszqQKPruXVGwY8egC
LH01t0di4LMmnDnHSgJxB67VyOP9q+0TYOYDRDYndSipfntOdLzG+W+RZbTFCB5B
hq7W4iPHw+L5VEH8qouYwRNqWqq13fsx9tZFa/2r1YKtBihS0Rw+QsvxisEBRKqE
ZnQcet08wqEYTybEjbhRZ+w4umjZvQzPmidqHi+aQhk7R3wlebsbjASnsZc/Okb1
o3Lhxf9O7fm/vtDosio7WvR3nM6L7cANSqmEDDCoDA9e9fZeK5WtuTxH3zFPNsAo
tExkSCs9cNOw/M//5UoZPhV7z5M8ixg9UaJydBqdj93LGKTCKBbz6zrLT0ioAae1
NWTXJWKE6tIa+Am9yuEY0bkMpZip7IfWgFdJrvQT+QcFq+65RY+Lyi7xn5U9IBCT
TVudsNxQWvGCX249O8K9FBb9k0i5d/QuR/J4SsUu1QQ3doGfrsydyQW/iMOPGe4K
Oo6FjUD1uVTRByk7MTjzg3erUbB3eHXGCoDZeASLasG+uSSsud2KZjWvJjxDdDCR
xdSmKhCuf0w0Twlr445T+cQ7qfTrizG1OW9Gcnugj5e3aq6zrXYtZXD9TIhWpgXP
wkMRMinX/d9cOWvm/bBdCpTZCY41DzRn2BjDpvAvz/NbCEUtSC+Mmc25CVNXEbz+
d4OQKDyRihZWyMIPgbyd0lBKFK09Vfc4rdl5++TPqkQylUF6tXOtamK7JOm6a0lC
qtqQC4V/kmdTeZrp7PgoWcsculRGm0oIxoinSr7AMusZjpHfApQCGflitrRwfK45
pFswcjuzJ2rYWXsDIFTMcgQd2JzQ6Ngsi3jjoCJv0mby33wHsC1EaWTr7dFGk58j
Je75NwjeIlmVITr8oEYtdVdleG6CZBuvkbrlphpc0/BN94+BTNWpl6G/gzsVTKo+
S9LfdjtWqpna4IxJE0Tar0C4wHkL5HdC2XeZRMgDZ0YHwOKbzlaleQVgttrO7bA3
iMdbd3mXVzhgb4jBbMsVrD89Ap0h1jdUR/BSewx+37SmGjdS+chxtFRY/h+ZfRN1
xJpXezlfQHIZF1WQjjGRMQJ/hWi9ftukzrX6REfZK5CzuCwpKmYGc4COQgvJKSe8
Amz7l5f6leM4mLmoVMIS+qu7hqoljSX4s9W4lg6s1dqsp89/PjNQWCKmjoRXeCxq
vu38tPMJUugJYUudc44XqUSE78i51ZHYZ0vhk+IWmhrPtCWq3Yyxt0DsqdFeyTKp
3fFK6042KX8UZIce+Uv7tb6pzkEfPnsVjmJ2Dez9paDElFZo8r/0FdwHKE5pa5Ic
B0fXgb9b4IZ0e/YR1asdilVla5UdxdFZqo6pDwDwDUVrBG15c9U9abGEnzoNiAwi
rhdIZbTgnCzWR3JUtmA+QXd0toHdgD2IoNchZnvIRvBpg5rMstcrL7YHPSyZFkwK
S+LjdEiQhqKk5C3V6MvRK3bHrqPQNiNXVU3mDi9bMJEXWhQY9Er4qldqb/nYxzNd
J8GYmpCZ6vVHL4k5ZThkWnDcpgsBaO8XgOV6c8xcrfXge3QvQ2rfD5Swe6RKZgyC
t9ad412dAEUmeqBdkcTWRi2T/eXHc82zWmdwtDxa7345VN83jf8t+RlC84t3Uhmt
KLvLTsvEIDK1OX7cNIcqplQ/DVHSU24KgyJiGx83yshBhZZvM0ZzOG/XDKyCFgJf
11rtQUvNVKJKmUOkc/0+bSNND4QpkkDaKewWCIFuyWAgZ9xq6fUJDvXhFqHmABtb
IcTqXr0kHAbQhjHGY2jRVtqiyWmUPbOs/3O4lZ8ptjhtyTAMRuIR/wERI+NStQlK
Ol+GhaP70BBV6HZY/7eSuj7ab8EQYcYAEWlDbtaddQ4w3d+fqZBpgKiQY0Yzjtea
z/QivJ4Oxgj5OVASrZ1sNoLnp82IMXnShuxGqIzitj44i+nxdsDVxS975z9RX/Vf
KFwoYWCZ1BIofOpxgcbdPP8shDdfOcIm7Kqn3w2GrH487kLnpMoRKVFxkSiDklP/
5uFAf4XlyAO63464sUCmCu+TfBYg+GjdedW0RVupYyWr4xJmpmFu9he3MK2mPQ46
3UyRfJneYQio3cw2qoAQLHIRpQiC0gI7q9q/Ky2wlQoQPAw82I54Jl1PHfO8PXoG
H/aPKFhsvLNuDC0PeCrrBrJmnuux8l3Arbtd55PJ9avA8zSwuDvoyjTNEgzp8s77
XIy4gpK/Q8GwrTveMfwdUsd8+Xren5vL4DO5bfpxbNNfTlCoZ8HERzTDj1CSGHhK
LkHVDLRf+ol/2fgfOLkd5sP5oDaQEVjOnI1YjVxdlMv3yv7VY5WpzfHqKplInIX1
0KRTXlyG7tnTj7YFCuIQ3TdVf6p0mSfBKka1EniaQywKkS2jTdRwIiCJTNrnqzt6
aC/srfKaEB9/J7UqGFVl9C3NstHpUGwguQn6v+avbZGvGtBeWB5FSES4SFSFaudy
jkguAk9gdlIM+/hRzSzBMtZzB0R0TAil744awQMO1TEOsZIa+IUpLyBtOvjzQ6KX
qMGM0343HlMo2uWYPGZ4aaB5eiuuS6eqEXBywXHfUl4dPqh29RX3ohx/eC6mC+o/
tSJS1eHIWaQvRsNpoC/Gk0+Tq+seNcIMZhCWLZHSkOszvsSlr51wxXoy4hZc9BlX
VlRH293PzFpdsPKbTiS+NqW7nz8F1He3hUrV70xlJXcua26cziNE809VIojwazpf
FNRW10sk4BwyzSPsQlt0sAaj2SceNwOcmzwvn/sX/5CAsDprCw28vu+pG+ccGdls
QfqQjikHhv1zm/+eEO0kiEmEQCeSg/5SzWSeivdSwkcYkbsIPSxOt+/9mS6XLD1T
mdzKamKLAvL4bPC60E9WYuoAK9lARpjd2wX2oQwG3VElmsJVIQaNxDor4KyQXG1V
zPSQ2GDiZRVFBOp3jaz2kLDwKGL1JtmBN7+W3N9zODWvjWRhHDznAI2Yrq/PqT9H
OASMcsSizbbVW4BxosWWiXQAhGo8nur8eiUpke2y4dyma2GN7Oo0FQn04TTcJOqG
treMsSvDORHKQ6MDV6WKHmySJMy8SC6MeeUI5ecLCJNRM0cBZpSIqusD3NYw2Foa
gaCt1t9soIo1mj88pCCl+cP3C74Gdvqm+mYLP6WMP24vyaSvuSG/DzLkpM3vsm0K
p28rsAsrOdb0bGiBnqyckVRdRxG/SIqEedckdUnr70vWiQ+0ktYLKOy5OfibGK9y
Yg6H3Xk92jab90xMQ7KppipuTw9xu/5FVA2vE9XnxzQsQjvwsFm02cAH+YKEETFa
v2WCoN9eP+2uyHS/DsWbRrpiO2qhunUdg68YwLCa5vgmRb7pwvoJge9LFA3Czf4W
MMKxL7qT9ejTbVLuk6MMdTtlzkqVIsC7/hSInMkSuCFUjZfHaVRHJVSdQGbHiwwK
WsCmaQTcWiPDGiQPCgzstpgGyi2ZsBjBuEuYnEBLMyfV04Yc3pnrA/gOMUhqZHNb
3FNaakA27AitD0RQIBzKjER1LDtCWhuq16LQXo7hGqBnAp9rmrg3Wb3gwEv5FsLA
2bPc/kLNITNZ1u7hEJUAXArg8wctuMsFawXkykbgVP7CRWvvK2Zj8V3R56i9kbTA
VLTBpFAIxf/+JMuDRRhcLHIq5astQsgmPMlZtzfIbLIAnDt1I28GSzzEdrH/hMPS
jQOljGrzgPd2NQkvCPfq4+dy/bGDVUMNOLs2VditzPM7TaQJoZxhhgd0uDDzzusn
aYuE4atYTw8YWPyu059c+ytiYTnEgVzZu0qkiHuPHnZ95xKjz2sf7QFse7hufRcM
z8cNOmAKP/tE4AkP521ka+pF17/2+IV2MpxqZdLDqyWb142wvOLAC6YKJ1EMDF8I
zxpFB3W6Kj6NIjp1gHIWW45tXYUWeA5WS7lXLVFpBIXldgqBh5nGo8GJqfo5VKRp
kxdPppQoPdmm+mevH3YUyeGoqEgDb1EDEH4qDBL8iMjtdi6I5NrrvzfytDxsURS0
Eg/WYuQlJt5AhIN81x6P9+tRQ409o+wWaG6SH9O78cGoSyeOcPihS5iSjHEMxf2M
/9OTBe5V9Ofuw1CcEHF/RcZ6dqyvSA40Fyk6tW8N5UBLIV+L9GSZUeoFzcQdd1EY
jXzFyQIw0mlUbPHwCRtsL2grRGIulWk0xG/+yO3Cw/4BaWz7kXzP0b0Ob0zLS25L
zd8aX1wGWMv7HA1AF0nhm2LRqwunkaCS35LrP5JXimuYg22Jv6dgu/3M2AYn1+VB
k9PbqCjyrhF6hobo0K1Y6JlHFko6+SbBcC3Re5V6w98/EtY7bAKh6wIYminIQAaX
GcUNp3iTF8mShpqUhg/7CkiJ2ZrWjIWFdt42pFndW6IiGQnj1onNvR8EK4ZA4MwI
Usd4uIa7VBjo/iJKV+GznDx5Zf+iGNAk0sBxoJf2DuwcYL8pnEF5f6x+JsaHWsqK
V0u72Mgya/JVBntYpodZ+TWZ9U8KwcXbQZh/HoDnrhdimvLtKQCLU5+suUnPIjgr
pvWoQq77Q+Uaz/SBco9ab6/RftryhL9Cdf1kfSelse55yxJItuEvjMO/9kFJN0c1
nILSRrNoY4dcfRiIBVBUdIoR3D0X7M7xDm5uJ6qT02LIViI786mqf39wgbNcGJIX
UNtrvmSExn6sHwUuj4ir9+jWQsvLqzgvUYfQ4HhiZGQas4BOgOjIHtRLtzzw6ElQ
PFHZ82QDa4dPEb8VB4GtOSIrbUBzBKFACRO8zSO5PJzAb3/KZ9J6ZIl2CLwD9l53
ELRurSTJAY2gg8EOCE6lzvNDyUUKaJt0PWSVgZMnTM9YN6i0J+DBrkqwLlcDX31p
b+xs9OCTLQZW2t8o2nAmF65HrxTXJe7nzdx2Gu5l1QYf3zYXMg7WYiHlYn7EVN1h
R1dmmP4XTI5PseuMqIT9R/p3B/1vY8Nw7ukrgY90FhxTGG7+B53EKFA8UsZCo2gT
eiD859RYruHusgnJnKS0AhvEAEdZPtww63a/7yAABj8w4hZemGK12fwirRA74qLz
WvfHd08bTh2L7puc9fS6VQ+wWfFuA3FzjVLAkYUBf7evp+jd4UxPtBvOZu1i5wYS
3yN1SEU5DdBxFhbsBhLncpvCRMn5zu1T3g/DBaSV5q7sHRY9R2rNWRrgzEad6jBp
v+tyXYStGxpBNJGmEeLTIWHoABSKZRjDIuEBLRlmDSPQq5DrwjtJ4cd6n9eYfOOm
zHOuvF07RlJY9+6CpCNpq/7h9kuKywTb5lh1tjnuheVIhsq1D23pTYIMUdoOfXTm
K1h4EQRgs4QkTjpMWOAEkNFxgp9oez7ouhPUlP/9mseIUmHRNMccW3JEnVkClaky
WpQ/ny3iWOa9B25Ps+S9swhAjKg+VUU8xpEslvgSRpT24niJ7pz4bir0n4BZtgpv
vuvyIfkSFyP9P2UHHvG/nGSTuK3xWJ/qHwNSmhVxjsFcbM/5FE3AcHpHY5OLMJeQ
B5eCqjk+GdWe9lmlZpYpHS8RKog2R7KbAGtYQP01z5bZcY7HFoXSxF7xpiXeaVBs
8aDPzXjgHlORj/3cHVVtXB0160rh557LNc1/6G3dkLbYDbJHHKL6ELcNA2DEDpY1
JMezVs3KLae2PXqzT8vM4sdckQFqrnBThkIBDWHK3PIBE7kMlFfiWvRUx1I95esq
K7EWsg80iWRSo9QlTSOSjzqp00WNQciAykfrGMfHtVZmcHLco4Nk9n7v96M/tRzQ
VXW4owvf9YFAc9G7aJmX+k4N49z2YxHukzhpX92yk+DFmL8aZiJXrxRnyA09UTK+
kDaLB6PbzxQ60T0j/qXSV4Qu/qRyibYk2GW8dFn0FtgxH0OIyC38K5LxW8CcmZ9F
+/Mm2wD72cWUF+CQruTSWV1sv/qOmFC/EIOhvb+H23EBcs0nAbPtRJWhTll+lLjS
Aaf+Ci734jcyMXpvIvBxeoFgmfJFbJgL9i+avKwOh7h+sxJ1lx/TQ4PWZich4+/2
PutbdUpE08qKvHwIcg5fZCXOsUn4RGMJIaQzjZCc9Mui+jwlA9gOedggd29k6DN2
+C+F4jCCmF56xwwRCfElYtY1gBfW2ZZj2T/6T3X/C0wK0jHZQvw+R23Np0nqb/Li
HnPFeGGMG+I7SRfpqtYQhb4yVtCxG3D0VH5yRHnkDjdtItuWKVp7aAmK/pcVSOF7
aCeucrxwHPKYdnHUX+Nuqjx9drgx4ujonD/i1fKTcKQGDoIpVDdB5wywt1Hunf20
B0n29W/7KCT+84CEebdVI5MsIKxKZFjtGYkRll8rwesFAeNL9NB3ZTOQePyby3kS
J17nZC8nPifVFNvND/tQmrYTkPLvB48tASZTU3IJxbBwXQXnxOIgAGKl5/HVsnzy
6MF31obC0mFjCa9BA+APPW03s54fFY53WmF7ikzQO9DQX1mLu9wq6iJVA77Ov7L3
zAkCLqTCLrBKpG1P5rkIN1evUcJqgI0aqrtWCkqrfF/tkp/K8kJfl+cKOsL+2roi
BhhiYx5E7sWeIWV6rFYCc8uZW6Y4albJHXFMlXie1oa27PTYgGf06pdymDHIMIiP
wErpUitve07sDlwzgvfG3HZgriPODScKdrOXaLvDrPDJabMR3s2jRY904DUxU1Ys
AVWdkIOwx1bANeclOrFPAH5zP4nZyuzYa/19yfxXwjrZDIHzFo6bVPb8OPDPU9e3
wA5TXexKA3yKaxpE/wGsE+R/FMK8Xl2SNg84G09vKJQP5BwlVgwlwhVvz9IfjaUj
uYR10OwWhv1cmcNebJL7Ah7YDVn51vLaUR0K4nJteL6w6MUBkI9yyjygrsmi729N
6wNpQA7SYeBSpZ6waaSfRznpCMIO8G/UDWvqEdbEqwGzpVsXzg8V/BPpNoEoKwFJ
we1GL6hcHXiZCIwQAjgDWeRazCgLJKPQ4ZS/bwD0nybgsZPxBrUGObAYCeyOQ2Ol
SqX1ct0exYlV287bdBcwAm3R+x2a7fDw5S/DFe1ijTrBM3uvpT5G+I3LmTlPe6VF
x/T5st+Na49X9NFfPNOI+e9MimfVIRWJzOgkQN0Ut2tNTsryIcW1U1LlZzwIeAKM
l/azp8Uf7+Zp5pbM1A1swdiPhd+A5WDSL0u5OjjshwX4BKuS022UVANCYNVmWRZl
PcF4XMgeyA0LOaDsk0y5NkbiqWUUmFp8plOqxmqi1RfLwmuZD5Tq5LOTOg430k0T
pO8cC6WYBf1SLdxR151Bb6IVMyNesicYpgw53qjczjm79X4RDu/Iz+vD3yww9G3c
Svf6cyX9oDpYB8EIIqR0jjzTKDz+nl9hXOgQQfcrCLxocZQuVa0VkkocvG68pl7W
TAt4L6gNZkX/pw1BR7StBbuU8GwSK3nmJFHiiUhuMOqH8ReT83uxyOfDvBSdbZE7
Uz/IWzqG7zeEM4rXXQhdZ8reaV+6DwF5qO9jhfnIY5X8/abj7tGceFPdxnQLps0X
8mFrINZUzG8fchSzxIMtIwXOeSXnbit6/rRd/v5nMWTaFweQKiPGDS7q8pxHGId6
d3BKlNOdtH3EYY149oSSFizXIKBch7phg2VCOb9HIxmUaPS4SluWkR/EdjVb1tmj
aS6KhEdhaY78Vf9bHbTRZX64tqpeabcCYIKw2ObnzgZ/eS2CWuKaFcaCWogglLcR
rAgflJbpepCzxDGkMgaq6bpc0vHWxAaJ2tJOOum4eBuyM1M+xxPSNsMjnpliNppQ
AeQSBxWiFzsZK8/WnW/5mGCGyTFAfpliHd7j1VnLYz5e7OekAgn3czaaZhklZ9h+
nt2ulf1/m3NiZdhV3v8m/+R3ULi16rKOawb4Kpc0PoZcN/w8XkzMIQ3gqHFuIYFc
jl7t0Qy2a+lBpD5b64JHpa9toE8mnI4xj0QKJvbVsFw5yFj8T4LRxv78x8JisLna
gdAV/PudM48xBWHQcYXmclNhF6AChTU2y2jZdNxcJ4XinSrzGKuU4EAY0/B+rQ+o
z6LWIzoD5rgDnsv8tEXfWVLdteWxWmmA3JKkkfaNpRhW4OsnUWonLmExSEUkucIO
4YoNS9tINP8Kv/qF1P2xEcIjeMLOgBxqqkMr0mwgJBkNti4cOZ/+wxBZ9M+54fFw
MKsMsAUCfyrpZ69h0bi16RY32ScXG5sJ49ww3kdhbYEsupaubQElobWdGQ+U62/w
98lAaZVQy3+g+Fx1SoqL5gII7o1hQRdocfbAXD4SRt7bK+AsBwH4Iht1g+6kziUF
XPn+vEKAVzusb6MF2U6T6Wwp8y4+EQR8sJxqYzAeEbQ2ZZCQZjsHZqfaR5ARx26v
MlJnRZHB1VvVnzr6RKqiF4yU0jX4VOkWPG0ZGGM9PRaRHPEmdk29HkVfivK5viOG
K3lJttebbZ0DTymk8uuy5eZIAqqshg37Q8+TayBWQ/ls37nex7qPpOK36bxjIcrS
x6G0R8YDSdKwWOBDCBsLGWme9ez7YrQMJIPa7JvHZ6S/1lXsLmGrlXWZNUjXJdQj
URYesxkB//v3aXS2reBpHzcdzmglUWmWOa70ea2jyDWeXaoTUhiEB5a+wSZOViw0
szgDWq5xSOmuZClTl32N86HpBRvHQuikzxnKcchTzYhCKPWQ7A3I/o2PeO+RQmTk
UYTuNge6CuZ5R8j55gKRH1o6R42brqKtyXdlQ3O//Pqdq/2jTo2GS05sqY81iNGC
VkwvpNliFVLaxumOHHfVz59LhuBprfsMRDHw+ECEGBLzthkbTIXH+qF9/Sm/Hgxh
sYNIm/VYPDITaIQeWl0kv5ARjaNlr5K1udhAFCdc7k4sCFPwi6lTe9coOMWiJY7B
Y7fF4+bYPoNuqtu93NaVc/fLxAK2B5EdbYwzqBcbsptSefzUoIxZJcj7RZAHe9w4
2mBiiFZ2CQevp8IOch+FKxOobildx1k34fM/OzmPmdV2Sse63+J9J+EPfBhYJgTU
xeFYahxx6VDDUq0JL6mrBU3WyNYpZ7XGLTZSRHBPmDCciNX1yS8MDML53/KkNsfF
dd2Vsi/x0iqxgTH5kZQL+yIJQbzMIa/0PHko6H54zb2dKOBu3gK29BLciwcpUa8V
vFq4y5367RBARZmWOdQtdC7P7hY7brVFlknekZLuZ5AwrYPB+iP/tTazt+th4qqL
t5hctJ+eTdES7K39AMHuUILFAB3HLovcanApSf1VnwMNCpjLJie+XirFQh0HCZLa
69vTy7LhpWA5+RM9AWbQaaiWkMFBrVkLCMNRQw/pBTr3AJQrq2n+cdX1pd0LAsTS
PCc/UpXpQWd/sh3ZDXYoXpM5Y87VcMxOIq7h+48vHiyOflhJPst5LqG9WsOgCNTF
WdxTIukMrywRpFsnsIfgKAYclzBT991E+pKQgyZ4s04auIBPHNVGaPG1mX9QmGDf
jwP4xtUzGcRTsofcvyQgz/ia7vdrARDvnz7zXBWjzrS2PxrBv2SvZx4Y6O3rjYWA
4Ds10oj6hU5KhLTiBaLxTMn7jS1r5xl5h/MmMiWku2x4Vi8nAB8pBKVVomsEykTM
djb0Nx8N35jn/kMEWh5AqL8hoT1Gi81G3L9it8bk8m1C02T10pZHkFJDSU3FjJRQ
RkGSrqmPtaZZ+PGqvlO45Jvjd6mbMG+ElLfxJOzdcuikh3Drzpv1n1dImASJgZBS
kbSjNafo2fqPUaVRQRZl8TNcaGTQ5YXS0JmKG2vSSCWC4jpV3e8r02kmPV5l7c23
SeNM87OxgG11VJd1oz4jtUHKmzEW6p8i0+avV6SG3x5scmDOW3i/KJ+fFW66eWk9
BkmvP5EMOh8tA/Pa6LCO9GF8V3wPcoaz63ldLQOKxxy2k6opo3injf8alvHBbx7L
k+hzYMPOMXpnzvZ+j2HQkx9WqzZK79ANJR2lDlxdVf9fDCmKeD4ZcdLJ01nbI7cF
HWOpcRlE62EbvyimwoQIeT/yhFn5bbRadgIVvqmKegzrEnVtL+HcMESd/mwS0D0z
gVBzdgMkaf/+qXR/SbKVLrOuxxvaZSBdkpGZrArsJXnONc5sEvw0OCVb6B9Ue/mh
rnZOdOSFBwmUC18I11CFtoQE0D+VLEs6zRmEsiVvwmGro4nRq/kcb26TacJhpzly
T29l7+V0fz69MTIcLmKrU2vMUbEejV1ksslBMKICGGjv7rGYJwRitjQ5tAtLb/OQ
AUNNIxKd4/wVukKa4PyPqAAyzSUuLNrXgaw+UOz5t/ZLt+TfrEQGD3YcpwrZn5Zu
UTgdPRopdATc8akRaFqAo+m5ZUrm6EVarztWejt0UZLc1wqAeatclXF8oNRHdrR6
SWsTwmZ/L5YMTAwY8puoF4nsFZ0MnWLoFhP4+mRl2f1pCSLgS/c7WiX2nppN7DaR
gbi+ftWbP4qN4AF+YPoTGM0rXxuIyXqULokgHBBeSnhwoDNaQdDSOiBrSZnFiWhD
N5v5rSsDkSqKm2jeUIlM6wGvt15wErfS+ADFkSnxRTHlfLRimU6889uDQ2/XCs4u
83CcfMGm6JNeIkfdbc/SnmX7NpcLi9Og/HoHYcERDeOwmL2YOU1Pnd5QDiYqEmew
AoVL84G9msje2y+SSOdL5+PrKWAbhc+9XoMPLvBcQuZntL2Bi7ipvJOvjKGv3tDE
67x2YM1kF5MDM/FmsRnQ97qNj7a6NIyD+90/r9HoRm4n4c4JIux3Jg71ltMuSlO1
/5pmGw98QQGft7MJ6lkdhqKCnAHEkCWsQ1S1E5xBULvcfku7RPalD5HJ0PTy7tG+
w1yUvry61C03zZRaEGyrmVaqFMCx7Vy8mW1WP0WWwTYJ+CK1cVmZlsy9YweNsB8c
xtdf88Ap704DZ2r6Ee+jhJUTnS8XvFgu6SMEgHPa8Jt1RJCEllf1NDUnLCtt1iJp
u/oARx/9azuL07luqUsaNKY7pM9VEBE3kwQVn7+Xg6q90Vt8VZ9mPkgengRPXaWD
xTmUSduPULXSRv/Hmcu+ljE9pyoBW8VArqS4JdJpkUnrBklyJfsFZZ+bwLp0pY6q
G4FkCFr47ROLtjQA5QE15zLhQhIxDuHM0iSkDu9V5aasbiUU/k7hPVGC/uF8ugn7
j22XIBmHfDHL5Df8BcG6FkpIzSpvV0zzeIbGqldS+xgZmQ6SHaGiawaQv5V8Bk0V
6xcBLmNf+4sqaJnMxNQN4pPZ6vmiaxDzVEMYOBytvLn/N65zludRNXJoDQbKod8Y
+pz+NUOkvLLKlBMPQuaUfuT7m+CjeMeGr3u2eOtU2VZeYmi7MnadWAyyTosVUSqj
+bSSFaYRPIScIyRp5KOOWZhTK67GPvGBS/cYLUdGdFyxyZsje9O/4qkvCvaJ1I7E
h7jgiPOadWt+o3eTOWQyoC8Tdh6i3C/X79PJHs5V9boxfrvx9Un/6YMK7ESWuqNU
zbgZ7FGZ07kI4yKahYQh8RzjIFb0BSakIAvCYHPRjpOzX4PLH2J/bRzLdlzKzikJ
M02uk9hemgI0LO1SzM8m3Fbt6qy8VwOEcznPhqXYttTjIe9m2NfP2GhI/6ubHO80
WgJMfNRthQ9u3RNfVr9CZcmr0SXBsJArXGg9kj5lCrRlkDO5RjDxtTKeas3xudRG
kMDjjLJY34Jz/BZBoxtg9GCxYqRsVZm5D4ZNRHvbvYz0PqeZnwPhANc/dI6C3pMU
SFNNp16JSBdvpQxup++yOxJ8PajpDu5QuamhK2l7ByF5O4e506ESatPTKzJUBfQQ
h4wyw/AOG1PmZD1GXD6poL4kggywYB/OvQwDO+TgfYNCq98b3+CBUyuDjHE63jwc
xeP7ZddkYJQMPGsIVXhXEiYc5PZvACHPYq7/lpm4dPZ+OQBBSz75mMPZzIts8i9b
5Bdm+l0SpuIAAxbPAi3pw8DclN4AXlWfBupG5zF54gp5vOf4q8UUU2HepXtLI0fY
EWsK6Iozu4vSXkbfYBdb3fd8jeto7cjukBJAZ+1VuXqbJ3G6fLV6LjKuIOy0hRAE
tZo7hWqD6/Ty0TOIiAmwS0Ivuj6CLsC6ejmfYXTU13Kc2tEByOURObBav1zv0I9J
VvWCIJl75LMEr3csL7+L6EWoHSXPaZiioPtrJ1S9zbEu+FhhFpUjja3mM/KypZa7
hMqiC3MRm+TXaWhzntRkWCDnoES/yznplrbiSxo3blM0PH9oYjibM8Jgt3n5tEfw
vR/3RRRZfordX+xJov87R6A7Jq0HaJYH0ZG0VolZILn7KFkZvR7NlRmVabLRNN+2
SGdnuwGx82PU5XaZbTrCvo4TbmwGHVai9bvEJW0FG5qaVS34BnLoJdvcu+HRge2f
UBcBgNTe9B99eWt4FsNB1Kzz8aEu/AMkrdgR4l8KWjzv0oTLpJsM7iOHD9kozwpl
3KRUnjSqrvU6CPJqOXL/FoSRHymMyqEQs74BMCCUmljmS7B2UN3WTtXu5S7/Frfz
lVK18U4E47QxB1vmaFvo8QnJiTbi+rH+0c1CxmbxTL9O5kus950KGeoKHGl+fP9H
/Rk/d29cTw4aXF6FmY9jRy24N2y6h11aChLX20C3iNQtgWtDi1toUAfKB1TYEPpl
U0MPUjJRBpZ8JTVNRDCfZbojpURZbYKJtu1+hno3wy27B952gygNqmN/eZVTGqQI
N08g1U7gE/c99SH5DLVjsae1B7fWw1KlaAHCYqRKP5GrSwAaDPCbYgqcrYN3lmrz
8S9UZ+0+0GzzsAdxFovh/JIenhHwwG64WEaS/e8w3i7RUNsLEU9JOMHcvHyfcE29
NZOoC7rDSDdv+xbbwGgs5+NsefGNY20LZn9Em3EET9cE1gYG/KLvxkxAl/ugtClS
arsFEje1CP9bHV1+8N52l4xuJ4xcblxUZQEt1dnW1oYAf8xbg82IKMp/uJwJw0vM
0enJnyEj1eJLVtXNWKS8LDuhHEHJghVqWBowjBfxix6R81I+vJrKe4DnU8ddAPDT
UEuJFLCQ5hRLOAYrKGK+k+WYuA9qwKMGpAxIqiG7YeKZm3PpugiIE/Y+3koNCCAS
eCRiLT5wrwxco6YhX2lHfTn6jaZsi74BK8ZQ+Rid4HEV1MMM0M30l8vwvWM7FtEq
F4E8zajZMjY2NsVi4eNLHw7ZStCF/zc0rA+TLwUs73kceRvURa5k0dZqsXp90aik
NhO3hu9JIe+BAj2WVjHP+pNgOUDxUAeW8Zfi7AD/0wRqHMyoDKS0zoa0XGPWvttu
X5kEwrXx6hhkWFLSRJVMFagWoo11Lb+7RmlC/CXsMxVibG0HayUEQNlSngw3FMOg
xJ3t4f/noe6ohrh0OWlLqDodq+qchiIm7ebZxRxOJzf8eQdIzErnbOAOXrTVc1YX
trJ/EkOTOm5Lq7adCyklqVs0CewQbYSFr+6iwcPcdRzKHkMbGgXIKuZu0nMl8Ftj
fMaMMbTgAxFOm4LH0zQEcIcxNY8kZ/etNXaJFBS+H6sz++lvnHggwPbxuhEj3TYR
8VcxLMJWtxFSAsxXjQ+kRx0B8ZPRd3auhcWAFOfjL3iVaHEA5NqRp4vpCPn7so2M
D3aYdN2tvlNYIvVkl8+1fJqQD1+8U1RrFLhoeCGoAFhKqab4/auFF280e2RBUZNi
zAFYtQZ0/0QOtEFz+8WSAVwMB1apv1fMKq3f5549ZbpV2i/yN2V6HZp6EHgOC8Wp
lYU+RRuxER4oyUGNgwLBY1onRa6/NFn5dft3A21k+nczfupPH3o09qtTE4IdKPSh
KvB8Vjp4T1Y7taoc1o3eE+owxAC9OuTTcDi6LN21TTahMDS6lEHmpJTtmNoZjY/j
YpvdrwjVYbKdft08c5l5ru2eO+VOiSpQUA/HSfV8deM00kzi66bchDs7IsTWLiPF
iOdROJ4T0+Bfez5tlGriqyTyWkZLlyDK4KnQc/hTtfyqxk0APgYYHhItoUjt5Z63
O+OLNW7DmJfm91R1LslOIVMFdd+OIZjMOQnAWuNeBlvHYcoqJ2IP1wiVPJDPfHxW
5F3M2UY+C1Tj0umK1amtssi01cXM0MU4Ac0pQQvlmFzCfcJ6dBzNRAviCZANsyeC
85IAGW1uopAc1HiUiQ4rBegFAoUKDoXzJ9yW5Qus+iTQaoUu6/jUayIUQ5rpfu/j
HGmp7SbVH6dG9GZhe7HUTZIskKgCDVNhGasqoAwe6s9MTfWkIEgMUIrTC0DYepf6
gEz3mgyzkjyTAs5H0By2EmZqSeKaZFd26tVm3GSYkt0f0BldmGSt+mp3HxEd4/rD
2CInhswIcufM0F4w7oU9QyoVm6p4p4Eq9CtX0f0xikQ76ynn4DVB6B77gW34/iu6
Jel1GTsVEYLymiBPkZzxClwWE0ENZRxqzVMo5B26LjcafX0mxPymA3iK1QubsxmR
mUM7K7DeGqKbDiWUPz76jt33WstEHfyPsxTffJoYgJ0Cm8W7z1dZMOonnsnWD8hB
Wg1u0Uxs73qEcQDQnDev/7hTcJwK9fXaiRVQwEO3Zf6k/6pITjKMsaLThGkTzCEN
3Lg6NmgJ5uPUXqp5EoOw0J/7KI3ZeoxaFkvka+s3DXVKh7XufhinngTCyynMg1fx
LTL2SuNT++Bb/I7rTj0ivsZZd/+pmsO2V3uZwyp9pyewKVSKoatSx60HK9KHoX3w
GhfdUsxTHeUgmkP+xJpmuJLEgYkxxxm3pNVQN28Z5JHvHwGWLvSQ9zVwCT+gLZNc
WERlXMzDvr5XuEdgu1Y3NBFPHoNldTZ1gnZAGzOpvUwkfPbrgXsTO8LzUZbpnHxP
PSM9HpThSJG4OWmrJfCoWGzatECskgdLqkBuhYECqW3vfp+LGxY2l7Nc0mG3qTXb
beA5aDhiUlz6DxEIb7oHwMwxRurB7A45vjhFXAUar/pnq9g9LvYoCNomSd7UePTG
3M3fBW5Ka0rwoLj0u+iDOLAEPDbToUnxDFfFsF+oAifvZtDNR76KrSqHMYJ4q/lq
GKFNAKJ9sYFQ/TDXCoAa92dPYYrq+W0dJ5fK5PnE0QRlCWv4lf4MG6Pr+04hjDiv
AlUEUyq6K058AbpPFt0DjEtL9sZZPebUUmuhZ03S+61Cm6dFoW/SgHSZUz1zfJTU
FkyUsxFY7dy55rDE13mCuDV8/EVJkbMzgys7IGJCh0OOCs3dgusI3J4lRj2aQFYU
0ih3huq5LR9BGKKhMi+tEpkgKgBqwf2/WVPaHEEgcE0oVvkMj9vGxz4MlBU65eKb
YxLoBV2Sp2o2qCkuQfFG/FGXQMZqBZppYY56NvwprfGP6T6K7Tf+ffOIKNFCjfr3
W98jPskoOA2zQw2Zwc7axoAaccoiAKiO8UPhJD8qTz90R+Cmb8knwSvOOknQhmR2
x2yx7ZTLKAYV3ufDvahTmWeezF80+Wu8G+meeBREiKBPhit6CRkzHPiYPSEIVMH8
6xNveg8cgRg3fmZR8bGnOPnaP2bUtLU7yjZ7LNOLwCQ9ZKY/BoWX+DiwxDEE4loX
xvQq9iktAv7hWHnYLCvPyPy16+OXB8bmODHJOLlAngiu1Zz7IBHd3idrnSC2mKip
P0QE3qalsyiOb8/si1t/sb5PbXkyLZbTD86Bmo8bioAzfWc+o0oYP273yQ9+JQId
kmzHVSQIJBZY8/4Rt63MaTr9b07eg9EQZHFgY4WBvZUWFMqvhnruVW52oDh7qLMT
/WhnCl3fGyO2IPdjCP8B6IXYd7Ro8sBGfdJQLE8Et0yywyyn9u4gAOYKrdeVcGBz
r9L42jnqGhdxYRTZWk1lmQ6Z+rIXLDejJnZUSz1xq+eQre3bwLzxkYucNdqLhezR
y2JkyIk82zuqkraD8s0nfenf7GjXyAgRsnqmTf4NTSfkXdBxG9nVNNvrsIxKf3X+
JyQHFxHHtwEdipD2LASl2GYi0ttvnPizgKwjpcMUyclfjNra29UQbDzFgvsiKFhW
w7zvLW9E7YJuLOlPJIlbHzXDw0bcc4VYPqQAiLZmGmvcv3wd9V2VbGcJ2Tf1j8ED
+ZKAdshZdevD9Ay4A/nPsVWGnxxrBjNPSEuXE87P0+LIcmLIl4Tt3a/j7cC7Yz9z
F6RxuMInruWJj85TsAkvSfgQW1UdhgvG8jk4AyOujGgne8bqitfvIQgTqvBP0Kw6
1xdUwNuBstAwqmLois2PtmCojQcrXLTdlCDtn1rYxyQ1XWbQtebRBAVzj9iKPfaO
akoRaG/crC9iHzY1Oug0dpJZcaUbkldEy1bp1g4RCW+nS8LWZGernpByNVIb3K4A
QfPCnAYkkk2sLVzZKVAQOukZEm5OywbouFf4IUbOaR4QXIpFLaZM7i7xfGJAEchW
20jalDsSaV75wuX+uKLP3iujCpHe/iUF3SFrktvVOczvXYUi4YfVMbhmMJbVVMtO
9QaSxpErSINNB+GmzLRiG7acNcF39Np+0LRRfx030Nu1lJlrUv+bWNw9O9EZJGJA
dw46kFXU2bGPoJgcJqkQqTz8euut3uDDK1rqsAAU93MyFSfKF2c0FqWbGWSXnPjp
FAiydFk488c3P9Hz38H81Dc+nFdkA0HmkNNkd6qDjzZcaxGzMDSRd0wP0v10Hsn1
Io4CT2mojrMTU5GmvjGCthP1HvN8QUpmIkQikw19qMUAVzW/qaASDWW6qF35ySx3
XVsDcZ7bgrbU5wUkkihpYT0r1wHXq7DqkMrIl8VBELhLDBuBw+BiTXQCN1G3g7Xx
+fn6gxvhb/nA5BHdH7Rec8BgXgyeIPosXWQcCobPHHfjMHJBlDeR+vtyoCFQoKW+
44rOfFkABYRmx5XG4excfVkALyvnKCkfJ3Y8pHQTh8wNcCuOcQdM/tHwZzQhbTpD
OrcElzNWCjrK5pTy6fV0/BxvMnoiteehgrp1QBedVeSw4rHSehPUoIX+JBMjCZKi
tPTMZmDPRjcsRNv7HZodTpBsoPGoND+NXBX7v8ZvQKYWwAsChvRH8UHOEf1kJHoN
zyXS3w6xJZfgX6jaC6bZzCxdaFuN3QXMnHgecjpHwVxpYARzIlXg5O5fmtJwU2VE
PflV6FSfYoRObcj4MOu7cjWWQcQetU6oPW1wWIwLchvQ0cOuWhlRiGsEmp/l7Bfa
GSho37P6a5PfjrylukEvJ8x/yKs7xBbilIJ+mYdfNAi6x7TJGwf85YB4HGSBGk2y
N8CfJUr27OjqQhLVbma9inO1ooQuLqQm/jiCRF0Fi/ALiPstw8mjyb1AktY2ZcNn
5WiYE1bBd7ERdKUxvIM7XFGvuJr3ehgLH6Gq/TBbNb0eKDRmp5PnRbGiOM/TXBlI
eZANlNzrhxicap7iXl56uZpwmq5i9G63AwRK07Izwc8XscX0kqMqkQ8q6sfP8cdd
c1kq0Fm1rEJxvEijYnSrEEOVU4IcEGXaO2MpoY14fAF8VOhQ9IwKAvkDAdyt1fWY
Yz1XmNB/PRni6Buk2vS1syJQE2SbDtzoBN7XdllAd7w+gIsRDr1HHknJ0eljIfOb
FcE6J5HhlpNTj3n2DkH2u4fZ4hYE16rYzQAT9OESYsJHkPclgcNusr7hI+0MAuRy
gCpAHY0Dkp22L13KnV1y4l1XXfyATv6P07zlnGsv56jKa2f6H7+bwZ1VYrqs4iwE
o284lXlMnly1GpRt4rgPi5b78MEzYeog3tUZcIS+b07rS+b5ayOWQoR7gtImWVV/
XsGC68TBkwTs7lcXkjf6yfbWXwVMdDui9Z++JQWNOP7/kUWuCaB2FlAID2kzG7D6
5oa6ifg/eQ/jZwvm3O/Uw0H8Ne2cgyChk9Ilzq3i61F3BdzkWqpXtKLBl0aK1BBA
3boG1av5/12UW+oGfKv606XAeNAnkx1cUkEAPvWFTVaIBU4OdeTVal73PIRqJG7a
Pwb3wGYJrUrVIiMyAGH5U6FV48e3JlM1YbBRJwbFnkTFrAl0z6rj0YfEHCNv+WL9
HHSDVo/e4xbN55JpeLC95rZDYdGZ5rLrWOVfPMHbrOJbmLnvU2MLQ8JDF6LxupP+
XFUiBDJPr7Ue9i+pLptZLNJsVyzjIFGb4Sp50qfUtGxghShtJnMN5OuAHokijQXo
7uavd0JZZP6R83XVXpCRd5ZfaW9f97s8gBUczvFxj1b3Ny35Fk+x2uG2qM1OCPwD
9+F+iuQHfe4rwQdhicAAsumSgXB/2Wi3VFdAUvID654ogXPy/S5uhycbxmP0dih5
eh85E2K4I27POFhtcCeAvSuAwdD/Jc9/4Z1iY/ZHuNwOQSIyvdCfsmLjc+CqVP68
SgYeqxRM6F4vxFeLaBOp6TY+1FiuA5dmk0TehZiCa+c8ZO7w+Jo6kp2TeYYvRcVx
1w1XKf6XPxiB43xbJwK4NbVpDtEQg3N/N8kwYKt/iqwiZhlQBHkbzn+DMzVUKHx3
x8W1oBA/ekLf+lMwTAEa8NrYcmx3CutlgKveNNcCe9EW1GvP21YjdZp/G1P1/cv+
elHG10JCq11fRQkKKP99KpjXd1x847+rOUEQPKKVoITTCHDQwwYv1wXXjlYc0lUJ
HV6kKhXiprYuG2CbW+DXrS13IYBPwThC3h2B8tGoWseiN9e4TdiOHKSHLEloSFdc
ZxAZJfUODYSEaiOyBsRiF37WQtHY0yZwFErgwT1PKa/2ZfKxMn36OGiBH0fpI7Nt
KLaLEea8U0h/nn8P7ZeHuTDSFIg8fXagpHaMfc1LjjH3PyaeIZ4TXuDSXbXAz3pP
CfDTrAFZX6+haNIuBGvG/OlW+2SwxR8120JO9CBZV21eNcnf3yi+GYse8rY5jh0S
ABuTU9AJvgMCHNKge1rEzqCxsRXIpr/j746V6IJoS+yRm4gdrw7tTfb993pKc6gG
a1wrH9FbrUjbUmBdjTTyjyVh+3lJmFsz/woIQgNWRE6R9RitSTys62cqgSD21GEA
991AqtdJqq/X1eIN5O5tv5GW2vrvc3IUwwjUkOL9Vvu8CqROi9kg7lpJUwMohwWZ
dz2/PcYQrlvjFmRMbae9J/5YOO7bT+nEteeD4KRrDy1GyXc/r0//tt5TEexeKAdQ
begjwzVCpvWAVl02Xr8QSH3xHtCElTqea/Hxo0UnXZP25LDdkHiMTiuBJaOSUwKZ
wt/U6/zVLyWhDYcTg/VOl6xa0BGMk9H28OlH4SP+tcIkEFHpMh9eP/AxX1rxtudE
HCxSNJpEjH3HYjVmBLVjweETYCG+fQ3jTkYMVPr30Ym7AoRL1yh4ZtM8W4yhFhC/
VWwXcy2Us8EZY2HjICeiAvCEswvJHK7384ulIR19DCdsRB3r3NIm3+hYgDmyf9eZ
etDRd2YovWyLJdXHSbZOURkQNO8V450075bnVwY82tCa3y9895RShl4XOSCkhqA/
qJ343ol8ABzMtK2E2rC8L09mtv7G7r8tIuysDtLJrfGXFaNxcQyBmOv34ONz1lh3
NhyEqFWKnUT1yZaRymskB67Y+3GvFsUEZqYyUChGc7srV5PBFaV51fUP1Zv/cvML
36U3LqSNel3biYufLNK8v6+oy1QK/q7PHEeUXW21E6JcMmgyMbLt4YK1ibZdAjRj
DttFry+fp1y1uOo5vzeGQCYDm0KQ/Zx8QlhjYdLdEhGK1UiSV6J8G9EH8nFcS1Oo
K6CY1MZtJhAa41lM58SHGOLFR7hi+kpk6FHR+JR30epdyZi5W7vBGedHmvF2AMed
I6huD1cyPlDWtuBRys9zisVmjd3KzrGK/hPfP6KT1gl5E8rc9mfVlPU4hlHnWfkH
dip/WgY62oSCDUMKGNvN1vy3H+F6W6ccXE4WbirKC3Bavihag7YCqPAa0jAipN3w
z8SBOJNTqYTblqfMG4RMNMOCiHDYrbbrTOn0oVqfMr4jv/MDjrwwy4rguKrkAHrm
Ek1FOX3omwX8ulibN7CqUFgPPFc7nY/wAdI6jadAD9gDqtdqD6h3IKfafxiWnm7f
+1Ul3KcvI6Hp5brucOc7vDH9VURy/bluO/3uG+rX1dPhRmiZQqofS7IxUasvBdjq
Ja9t25JtiHMl2cXb8NlXVVm7GZu1A4ZClcoj5bn8AdqdLbNYGt84EIor/4k4dEEg
P6UnfV8YuWzBoXfNrN0LhEULG1SKItGDgaajiIC7MT2rJqqZyUqBJVovS1fPQoWL
PYfS4CIV/oaKxFlAdjRUiZqhmCFxMhHd3FmpLB/B2JH3/Wm8CNTJ2fYzDq/7YRsH
yS63lVuJsLob+2zWkw2IUYWc+yG5dx0iJLuoE7LEOkzwpNMezGEbZAHRtFt+jXlW
o1OOhocEqvuVu2ImYSmP3l/oH0BiBZpXtT/gfwVG3oM52rAfFHtWW72DDJyWPBHG
wRuN2wmB3gKeZ2JUIgUchi7yF+ZEqWDfxf32Sb+Fe85bUiS04xX1xQrP5GsuHmsI
0yS7taEeROrQjaM+wyCvP8iaYoqmbKjenT+1X4RxILSguq7ra/jATXWMwwtSOp6n
qY9Ps6E7jadDvh2+ft6lqs5a6macNZz3up+Ncyifs3gH4iqG18vQex40z62QV3AI
bryUd5VpyvnGk6d3jRgure9fX08CU2rjN7AvSVHEwbuO3jzalehTGDAnw5DOoeao
I9QEXyeUYtoTZgxLcnnzvIXxhAiThMf9jxXK4lb2x+K5eL3RGVtLNAXpVykz1u1D
ewwjURWgOiBk0dlkmWbo68EpLCacloEda1KPOLqJ9eINRTTiowAL9P326P1/hJdM
+eMuCuvRUGi7V5jYzhxzXX4FOzxnQfafNy640h4v4oDN8jU/CBkwJdyl1unKnpUH
Ks6IS+Pcp+ZTPuwqL5XzqeOSVKqQofGf9W4spa0PpVcIOWAK0GmhahAjRhnRgqqt
yi+VygB2SsP8bczyY41/51yafh0HQMCfq2tckxmTeLs02UVQ9MuJGpGWILGC/DIg
KWCfwrx3b0O/4xTM6ou2GgnrLVYbeozWvBo6gufFc8mN+Pw3piDK/teMKyKfpfPA
1geUEPYZRGxZsuQUKsyzAzoVXQyCZ1V7C0DWUbCN48fQZP03YFHlMcHxzIJW4f/S
7A4qsXfDBsD0eLICAYBiyzn66w4UmwZA7fzsfqXVztIZ9schvBYM5+7r0gqsbZH6
aAfkbdiM3bch7MT8HgFuEMQ27oSdXWlxqpZGZCcxOykJPSmWmkobM2X3IOU8nJBq
sVwgzzSIAFdUINhanPXBI2g1JQ8BQ4ZFY4iTRFagD31ntNZ20Ep9YdrCmrbZjZ2L
U/6A1dghEX0eJZfcnI6LSHrC7lTMN3DxSvB4ApRZiViXmsipGiBD7+nja+mHN1CI
ED3LCnZZYhqKUHFO8oxARAdZXDUMMeV1ohyx0cMVzFHLjIhcVV/Djna0o9PuT5oa
Ytrh5lKeGkNFCMKHk9ulNX6hEdGXLphI8q7DGYX5PrvH3eSrHGKoaQLWIEFAyLqQ
1V5gb5f02XvHoBDgsgbwRcfF+2I37VUz2P6OYs8jt0AvSH65CE+qWTSvjd/2pG6Z
khycK/HGqyHMOcHCFWd+78sV/tOKdrQo9jdd1GFUBISdDCsDmFlwGcGR/tQV6RfM
eiM0p007xQZpEhE/TeV6ZL0RKeDH5Mmw5QOOsDBHvZdFMhd6NboBAuw3MgjO+/GG
odXVD5BuEkAy8SJObS/Ar/95/Hajz2uE0aJxvcfsQ1rXMx6di1m7jCQPrw4YPvQ5
xtGayTOqSAGVUFNKMYXjs32CqyjZqBp7mCS9bawQhfUG3BgXlfDXkQ9fBssIclNA
j4jcnz+uod4FpjB9MWplEVAlPEtVIColwLlzdUEIl14KnINmTYmqPLx5KfR+mE01
ZVgDKb+5LLnwXRk8e8iaSWT49nobf/YPM3N9LkAE/d4qP2ZcVIKPktjse2Wpo1s7
U0ThLoBNL8YfrjMkY9+KoLoYW2675IhyifJkeUNiMpCY7BqNqi61ULRdLZo9NWqc
2VeLjxwGC/s7vDjOKZWOdICEB7suhXkVKgwaZJ0mwNNiSaQKMu/WOglUufWQxnpf
xTHjfS18DtKd7eYY3BnGiU/3sEZcU9be9Z9iAluP/alFIDxTjwwIevzX2SOBnFqq
2R34GrSmqsT1rcJGsaV7tw6davhjUZJrTr/FBSqMe/GXqFybvvpgDX6qZTCvCyIj
GA2+zvReI0Z167fyOgGJXKcbBHgiMtd1vEFH5PeW+cdc+6r82I4cC2XUal+jBGPd
Drru2/ve4/My3HJZ+qKA7DiFwPdnYFUFh0qkr1U6jI+5AwJ8IB9VZnEcgsA0+Zip
iKIzz2E6fJxqyyokHj7aBROPHr0piraAWpswo/rccWBtZKjhi++cPrIJ6VbwRZs7
fTsBZpgRc13gW8jiQsJz3u8teFmmtNhrobWIGoewKiXTipImaXIn64FkXunCen9o
a7GsqWQJWU3PK0kW22PJA3ExFVrkB+GV0JVYT7V6ulTLk2mippW5LXGjEpBUtBCm
UUhf4Sgu6F0+RcHrNVtLZBpdA3AAL+lHA9sDSgSNfssugNiA2FwdCtz06jjsb4r3
mF7/lfj4yqpfmVKQrHcWhUmKiFswZbcygOaPN61VBKvSxiZ+WWs1gUFpFtKH7kE7
YmcDSfHdRrmFAWBF4Ze4GJF9Rbzen/QwNT3TfdIfZmHQzK+F0MO/eA7bvFALuIHT
A7sEY93JYuQl3hGw5Q62te9mx1hsLrxWrOfqK21/FaCK4N+hZLLofoVYl7ke1mc7
RlhZkpuKneGAwSApwalOgdFEClMN9UiiBisMUNejNfg6jhowWmd1IbKii9Ohu2Ef
bVMLHtQGCTsjzyvRchHTBJ/h9GwBK5ypwjxUgdMtEbz/NJBO/Dv3CJty/Y+RxSkG
6G0dC08ireLPOLwuFPZR8gQ3SXOXC7qwwh0PW/wmcL2VJcRlVaIlQcXcGdHD8sEd
zzlg7MVvEoBjHcdxDbSeUkeBpf3EIlKXFoDrXZ6cofLQ2RINV9UKapHSRGtUzB79
P+Ro/P7DF2gtgzrao21el0utNA3rcA6oVTZ31gcMITirKMlbUALs+RgAs8mwLpsO
EZawY7nIHaJymmrsXbxmbnEOnKQofE3kVl67NubEEnGxoEszcsAYsW1KFjgtgPfm
lTWIGB2+GdrP3Ay/bFJ3NaGLKAYzPHnNqVcvpeXwUrWxqfFIefYY8VoAxoEX04b2
lPM/R7fj/wqEP3skz/AcAQZUOEQNKZCUHAVJgjdAQzadihGrz1tw8BKWnnJ3EqRR
3VqZgS/957GTjg3jKmnUtosPyXJHsOiC/5THHQURCPsAxWTx96kifXN0tMyI41Hh
Fy2EDBdgGBTvHbMGEK/9jpnRwk/J4BA/htZfvxjxR35Oczl7lD23g9z4fGsAYx58
XjQTMbGOsy6iZzwCUGAyI9l/UeVfiR4aQ/jHgYeXBCbmtlX2o//1GUWxVFC9yUsQ
nzN4lOz4/RiCafoHWHYi4plMaCMjHJQZVYqK22Nh/2HycBFy/F6eiuSnzFdzZ5C4
bW2rM2K5fGWZAaknXQlCW7rfc5xBueBKmeso08Wrn9+aWbG5ql0BjrBlCcue1OvQ
iHKWOeMBgXSaboFWjlTPocdfiWdNgVgbzzovh4xbys1tNveFJ/hI8UqN9q37kAmq
/UCmsuP74AyTfuUYrd4EHxCl4ybT9/gggtpcoaSQKYH2d7XHV4xfWSTwN6FRuhF4
o2lMjLvCpTKF2GgUVtawqR5820Ef3j2fLo6M8klwy259X8BMFo2/+CXVb3zw8FhQ
hQxZLGwH8viqV3nOASL/8aq9VXJZFf946QY4qCyw14khjiLruufJl1GAXbLb7P7k
X9gSUjVGHtFaGUx8+0htcQonAk0Vg8dVkdZBISgD7gZeDzqqZ6fFOrTG//CBneb2
3wid1W45xl+yKTJ1TFUz04nYV8Ws/74mde10aORze2h2U3aAHo8MfHXUopWfOdqL
WEuJ9JXK28xeBjlGSOblTceBI88GrAii5Zo1toq9aVr3EvjtYKYIg6q5+MxT+p/P
K/YfPiPRbf1JDY/AhdvEBPiV3iPIKy9qd9yGwhSg+AGQPOhBX3WuSScu3gWD1kfO
L7XkRVlfJfSDwOPKQ4R+ysQ90i8zHzDZVYCVpTh3hzG+FtNlw/Cm1ZOGUK7yHTS1
IkGwUaMHH5EdaHzYPhqTklK7Basw5+G4KvAeaBVq3jL6MSycJr/Nfqi1FYJZc+O9
BLqMr5hS51gTiCKjlSXn5w1XOb3lNjOx1t8x2ksqsoiIti01J6SwWcbl180xamwG
OuBT/ECQ76fWcqJpkvtZYVqEfcCE8cuDJ11k/4HqZHd5YksXi+C6CuM+opHOI7Zq
yJlA/k3q8+RE4MpIif1vo4cPBnyY+KgaGv61KxZB8UZdaMtOdgUG0BAW+pQLodCJ
KaC9QHBwCcAWVYoBZvH+QRls9AZ6GKphR9Oe/034reZT5txtDjF18pGT4VjFzqmy
Cz0TjKimgFTlkM4HRDE/vRr+B50Lll+zbOn1FBN4j6Rul/t2UXEt2i1jggPvoc9Y
tB3kPFHngmnIhdZjvkTsarIw8pHr8cIWkqULAdff7ak3cXCbsUM33A8UB5JhX8SI
GQNZ5OEvnLA2hE9r9zjoGogcbWgGRh3zc7It1q4MbyZ/jMuBfDG/A3kSM11ZNYvj
OSA/fiqO+Wc35bqKY4KL4sAIQgw9CGtKuiTElOeGQERXksM8EjyL450jDp5dtH7f
zLArCYEta7LUccbGDTc/2GSiR3l0jHTbnDwgnn3anvpU8g8itgR8rtPXpwt5i7GH
e3J3jgaryegyVfqfiAX9hwE6NdAmSqrIgcOu8b48mj3De0sTqJutkYwHce137Iao
8VNRTur0YtvHLaUGuRRJP6NZ5b/4DML0jaeWaTzx9JdHDwsqenill/Q6NjPnt6TL
CoCdsOdsi/HiifnEGpTaG3EwMHiwZQ2QOPxCb5SaO/tAdIUXCylXUQgyjS/dkjb9
oQuMY46ZCAfJecMpEs+NrQJDaIMhi6/NhI3Z/pgZLwkAlB4BXC4178GUfHk3DPw7
Zq5/ZIcoud7J8JbTD/lHMNwC4rBhsD2DXs91LtYqjmaeEwAPa6G1ufVeoDJNmbuy
UVxc6Ozw/XcJBA9ueg6WrpQVkvRIkqlNVqNnVbImGu4ia+BRmRMbjih7d60zhVER
ZXkxTs41bLO//SA3A/9v9BzNWZ5BW08VQ+Vk+27TJ4ndU3X0M0jeQLYP/29xE0Ah
seh4SJqfIB/t31bZoFDcRKltXb7IJ7WHbhB4zc5EmUYYm/4+7fv4F/W+THpN9bGF
Vh7cs77UHNsNFS/9XSsVT/qtf8YQ1Bh8HwUgjHCzxMdbjOj+BtDom83s1KAV1gxs
uDZPJtMabps863TGS9mdYPdWUt5vy/2xACT3x4+k0Z4FH4L7tGsAtm64AvmZZNNt
+daUEEaLfjwD6u+h8V6FTiIPEUSaTjeTDKSkXDxV/tg2+rzlsxMyj8k9udFl59fX
CYsgw8vGDUz6V7bwTXbIo6iM4MzCJXk5JSG/JyxQLur2UNnrzrfMUPmmlaXvR881
2BM90AZEyYONHTOMew2OEQoUccUQ2HhNILtoihI7LOHwI5SupQVOvzesDnKlTzuc
fXxzKGPXcea22fiG0C77Lu4ecVu66XhOzUkcnT80R+lNI3mcRnLwSP1kytVgoGbf
mywGlsX6HbKUhR8uxl9CLImeIFn2t/xBLCf3zvmjswAK6hT0VDniv8l/VOl1pmWm
r896Wb1/CzgI9yxGjT5qcz7yLO0w6PxcabSKGYrvLfgwX4czDTpWdYm4qQUnUQSl
Wa20lkZpQxskePISXaKt9nErHCC7u5cjtQV/eZOwRs8gGkOPjvCipWDV2nyceD9d
4hYuYIvdY5SfrgO46cDz2UHlR41H2w48cpUWA3ryDyJ6uhWyoNk5HiPk+5p0c5iM
CXvArEnDJN4y3Z9DwF6RkLTQ2f4M7mP5JY6WOFYT2eY5Y8jxK+X8UoE9QWnmyRbG
vEsU1vM4vnBbjK52HdxommFRJyq/0MsaBqq2Q3Cj6saHNcceUDEHC4XdvvbtWdja
zIKh+8uWDWUfLdNN4M723mhoFiSaN7191B9cm/BDpTmKGdKEFIKFi4hJEJb2QRk4
/NAjyIi0InoBjyIsldNgU1Hg7Ohy3Juc1Z60h4p6BPLpl/HPg5+j8yGyS2I5k8W+
uIAoAHM6LWOSmze5z4nir+9LHt23QRpeyONeI7qwryULXXHfiJtYMEK8j6O7QdBe
7rmmBDO7S9rkxhCyc1vnAoBetPxnZSSdJTv1e9Bdde8u0wUIrsJveEFyDu/mHBrY
wwIkICIzl4sHwbzDQwej6+q4hdm0VHabfaHcJWvOpLzLfcZIKy3Gc6weuUVvnU5A
0ozRJ4ATuqFqgSFNQZr2dtC01H7e7PmPU/bKYBaNvaDlsGm3s8JTVjaZ4KiFkXIK
c+4yZ3jWe5kmSbRuHu/dKVVQ8a0/hxdRdHq8243lgP1bT8MH3hdNkAadQ6JQU3d0
vrIiIVGRQAoyhc3StSy1CnemBQlkvkinMt2B+aaTK+EwUVQPWXw0CVc2wNGronPU
8b8HLT3CDbQfnUFLtnNuMS0HlqflgTzV6eu0QO1L7D2sPIBd2cJqV2IpjLPpYDdt
/ssyFv38mOzRSq/lCrNfIoGzdHGQhb65W+xKQ68/+h9TKzpr9MvZFYNoKYCASb+f
WWKFEywhBSlEKnbbxJdkZyvzki/oDWG9DKzsceLCx5M6Ewd02k2SorzgSOE9cBG4
DLHVHMPw0NoZxH7OktAma00+v1PqKXLi8LYryEXEIiU3XxMEUm0RuVtKTOSE9Ul5
D7HHPO6oOVJhnm+zHAskHvI9Tq1oenl1db6tAocrrGYRXcm5iomjk1i0men31Ena
uAfouW4WCHppeyhUSgNNVE5ACL0LpQ+J00bDHsu8XJgz6/Yv6L8Lbr/Wzg0mDMYa
xGUScNdmeZrANV2+J3wyFxiJVA7eDW6XnK1Jggbjs17TCf3DH9g4hMc+wWjuFUhi
aLN07NbABMifsoSH7/0pagX+aTSIYO9aV9cvAQw5icy4d5xOhkJxeJ9PkpLyoXZs
vfLbAEPvO5dFa3Jv8DPSHaCTA1W1/aeVn1XqJWX0xemo0qKZjsmXOb3H92bv40vY
heIJjdskgDPKkAzH7PiyKKbiSQviTg3SGBPrpPNIhj3empvCTYn5/idWORU1cpaP
bftNZvPv+WWbHHrktH1aLHOu9CGbuCoJWrNGFFGzmwOh6y/EvtG6EIleosgELXTc
pYP7eCPq7Eo//KMhoA5IxyfsFoe89G6ndfBQK74st0B3nP2QZlxTWNy0ae4bOlU8
ZLFkQg3EtXQVlZn1MF2bT+tSsL/ixXobr/xjpP69Mlis9YSrlBcx34E94qV1/pHE
qVV20mu4qkjEqoWWHxgaKHIabSI4qng/01B/0hcxdp6I0dCX1e4+l7Tsso8HRAvp
9OOuj63rgjdHb5Trzeih86sjREStR02BSiSBYYJhEJKlZQRzfZmteVno8GZkh14A
Aq7O4gzwUePrs3oL+hGDW4Mh9aWaAk0PlsvFzkONhcqWQ15RrTX/C1YMGPJQNMPm
ZSCgdYDsSMN7TPCE1vM80PoSnMgidsND3QWmuI7mQB9sQPflorwJzt4nRTjjIzCv
mjyEVwn9YzYIKXCGpLvFbu2l+cqU+JIOfKb8DIuKZ4hkiCRbFnOEPpJmXN6B0Fze
6PCnN8pOxzHTkKCMkCnegDSr5sA1+rYicfWysxSJ0mwlr9mzQB7jtz7OHIyeQ4W5
w1We+8SE85XRPYRSLldscbxuOr3EY9QrhgAcSlXYdfKQn0Hy8UzykeFmAIALrhIJ
DWz/RCkuj6xDKdcZ8+4q2yJ88X4YxvT+TbsdO16ym+yNsFuf/ZwIs4qzMChiKUB7
OImD5BDUX4Byhdx+a8vuyk5Wmm6dcTrb5JwkVrHtKUwKFiD4LcvI6sSjJ8vZZw9t
WCxuTFZQL6179JGRThbD0itH0bLtr3eWiApkK7Uw4yuJahReo+28IRnq/FQF9Gc5
Cc2bPvus1JP4vwMNwiQeOYZgzTQIamVgRuxvsUgWoRzkaPQv6JPfi83EIgms9Cjf
RdKVVTMf/6IUJbalzquwiHsr7Yw2rHLaoFHbj3rAZ6eq3xwd0ydFEGdgnWpzrjcR
eK0gDnJI5gJ5esNOfbtqXaTK68EmmUV7zsHbUBYD9R9j0VDp7XBo47Z4F/EPcJaO
Y4MiSjvgcxf2sGpVg5Iz2euRDgTqNazyEZG3qKiQAOMI2Rj35aGKUbH6hAU420jU
7xxvIMyWU/tK/0W59BkI6q1olXZ9sc8T/77ESM7Tnh4jvV6MJGKNUNhx004qF8XU
7acrEqXgj3mFEfeLBGDlKAVmVuCJGV5bTyDy3KcLRIaDhJZuEBdXlQ+FquDUb2fF
qbCoiY0tnhMue4GGSmqg1W6vQG3099LtInBAQvB7qpvOA1VHW5FSQXnAEnx6hyXL
yfJli3+6F7FGEIyC+urWcPK4vLbbe5+ArdAOWAZqbFFEsU/k67mOJu/M6r5Deg/p
KGfPw8A/PBbLJeuHLzIapmMXSICVykHQ52mAS7iL8BOt/VH8wmJhAqqFH4UI6yaY
WLziqGv3rEwalbIumLcUbzhFu1otNdhinnl2HPZvH2QXGvGX3bRb1wRoaXPBwHKx
i2N55ZPSoeOtANedjR0PbpqQ7CGLZqNvA9stRGRxTodaBzbPdW/Z71Lyi3mHEIo6
k8kKoYMNJHKN8VTtMJCg5v3kEKMnrpFJi8xzF78WWbK+JywbgIf6xpUXnPWZHllu
Cv4HG63AH6ZEftD65hxeE2BPJR+flT9d2oKSubkhyqfvl5FFBf8231jkhxiH9aZp
yYKc6hDMfiS9Jd8mItcQVdrS25uUYDdKZpAnqxPh0qzavJxLocF3ZRknX34yCD4h
PZ7oO7d0bEsBqsuTQU7Gfs+4AH6savK1vJ/IyIW3hsvxbIcYSFGtce3dRpm8hfYE
JDQRR5WVyrkZrwAdxvA0UHNuRZkCX8nVtx6uhJQJ6EiT390/aksyDT/NsQsc864Z
yWCTI4xbGcjyr7dVENnTWgH9y0m4hbllwwiC1bOg5OmM9yE7BJD1CrSPyEpPKMbu
USOJQFLWDBwFeK/cKlv6k9wKkJ7jX+TpPBc7hVImg/WAmt3+qGQvYOcxXa+Nufel
TRZc9Fq0uakC1a1FVCQEfbP6tcwy4cmb/ckfW2KUrexntwC0Xah7AyTzSKW7BeZ6
VhalRWk5tkFCyEq/JA1yIOpoE+txtuWrCeci502Q8Xkc3ehxdoyqy3AhycrCOKqB
fBQVlAHJqBRlBgeUKaTfNoHjMQ9pgDQRAgtxcUuo6JrSrqMcgoIH1caYH7pZ1IH/
i6TyXPka46OlFcZJS8uPkyedPg+JfFFvxbBJHA4efRCMxmSeXB2Z98jNv+D7ft1H
8t/jryuoF1GPt/I4hWTQggCfVebuFhtNRNBCMkoGVwgUvfPI4vVil5GBzEbyUeBG
vmpANDb0VXGXOPRLSYokJ7/kZuZP/Y6i7hq8UJsM9SbIgvEep5TM8JGh06P7lyR5
R/6yJSgZiUMVyOH6KlmIWux5OmT7mWuAC5rJDnVmYmLend/8/QxmHx0YI4omHQgN
968/gzLL+ng1+rkzjRic7PYHJtNuKUAGnrdIp15h16wmwokJsU+OUq3p/p+xPbBd
o03XlScFWohfqcb2Ed7/LMR1ZFvpBi+zBnUDib91FaaaTDLMOqQtyRT9JRStx8FF
bkDkUsp1/GQ0u/G27/s2X0iToRib7L2e4KvpgHHJUoJXYorwxyg7Rh/C/9XaWmif
4oEZ/cY6wpVPzDH2NdNcg8SjI2to6zJxFz41XkPwZ/3wMpC6iEZnVIZMH8b4DaEr
/JXgjFOpO8I36UUu4PyU3rAo5oyHPZsACm1WJGvYY7vsJOiu3eOUUI57MPVxqgiE
fPLskw/9/ASnFiRU+JEYTg76vT8Hto0ArMTzVIdTM4W7GX4TZvyyQ8lDa/vtGj1Y
+92Z0MWJI4Nfv9xorOnHJhAkQgEGau6qYGdE5wUE/BZfOHAU7+/NV7ynn6eigMAP
gsY9zoDv1hpzWZkotQlpmR2F48tp9rMOlvBBKBJfnoNt3qVZLh0x7NTSO/T0uosz
Yk1PKaZOuSeuXdClOkjQwK+ZGdmfp/P3TV5rl2CcxMMv5McB88vIer0xHrd1Pg5F
SfjmZS+qMPyfN0YuWjTZLCxoyYpRYz3lgUFKnlLt7zoXAG3B/Aznf4/0FyrJAmZl
VmEEEp+qoea1+/3VKdeZnz4J48ACFCRDl1jycZJdLCaMYQ+v9HQvV8PFVcMH2DIr
QmvPI1Zwupv4Nwqs3h6Oxhru+C+gELgojqiEdPgX6hYS2xFaYtnYWf3nDDcRtZ+K
5EsK3q4/x++MkvQ/bITChbpKn1LLSw8K/9U+P87JlXdDEseJGF4lXmOx8AjCj6F8
qbJuzAwPomqzwTzNWxbwDEg96tIPd6xmVpZZAWccVM9FU/ixtVItfOsT3AoRmLc5
VrZrjEHNcdDiVwg1fXUBAEE8Yer075cgHoASgyIcB6Jpa7piagbLU1MQYu4lr69J
oCIzO1JJlyQUrZeUDNFbFs8KPyfN3vWPb+8oy71qzdjlPuNOW0LDPhAzDrYi6fwX
EzUU6svCOZVHI0JK+VThSKoc4P26wk6HQLuJa3811VJUTyLE7BvFH8RWQO/+q3h1
0JOPEREKgsD1JPzUbiQFLnHntsezyH/fLFnr9v7BJ9xq7FVWtKzI9DObSWxWLIdg
e65sxcNIyCloX0bLZsIQDjqqfoxa31F0ObfKIcp5uxSuzMmFLVruH8oCAtQmot6C
2KDHkhV2TokBHpCqBY/xb3+UqH6N3mj4un8y6pjlqlBCBmT1cB3Q3WsPuzFFVEeU
dKyF0+2XLmDtvYAOfn/jzNumhcSO8koKGg/yzfPa1Cfc5BhB5FAN+MgSVNdIhnLM
Nur67H6OjNWYj4R6R90Z0tZVIUhH8ZUd9fCp6wMQbhFthJtsout1m7RauRZHYd8e
8O6y7G1/tYGFbXojY60zi9IBVUH8UIu+sukY+/6mJDEchC7YuczbGuft3KmdiZmS
pEYr/Se35HpQ+5/29Q8svlVhU4ZTULYD147l8L27cin7n0pW2fBtGMXxOXFjW4d/
MIXZgyqmllRsAx+vwAW8BVe4w4EkeDvYRggbOzALFSAP5cEHNIoEnmlK5v5gQfrB
1/o+job+tQPjUXsJe62CLyRQtYaGFhsTqg+u2T4soVmOdu0bXhRGiRhLFHUTQYSF
xHLy3RramvryJW5erz6zUleJx2amGhSFNPeot1IUhSRf55RIjkhdY+Hm5DzpCQvi
sw3tDCVdsrzae5XlkHvRFFvAkl8JPih1r5BVTQ748+MlHZdYtaMbpr4Ky1+6Xet1
655fzsk30upX2x+5J9vAkQQCqof3AJpsWN+XoBvAkIhiOFfoqpYcK8OcKyU2zUB+
0M7bBnKg5Myh336f7gS5BE/yjXg7pBYmM4Quj8wWdZ4YnuHNb9MatQcP9ubqd8Uq
OVHmdu7+6rJvdvDBn91ZNEKNGxB/nWrLaCuk4YnimEgoszdCYJv6kdCKGCgznZgi
7KEv65Q/MOsBg7vSC7QMVTsBxM8n9X1uNf6ggTv5fuiYure9UjUAS6Hwui4YEOZo
YJW2DkUoShOmhQfFq5eO6CZx1cGIzcNmkj3rFd+GQaEKxxbl/qam4jj57TZjlw/o
tktd++lIhuEgdPr2BAaivemERGcJlhwsch3utuusgJR2vL9jD8bZsR7+jNc1AoE3
Px6wrCh36lB6NfUERw5sifKhNq+QlAVQNcbz1amnXSruXhC/8brffRwk+37FGLi8
1oASqaxboWKfXIiJh2fFBUn+2/bJjbYbzp2qVh0A2WVBfnvcTPPRRTBxz3V7qtpB
qUmq3hDMUwdeKoKMT2oFVyYXVV+7KfY90kW0vI4xXQS0RUybkTTFQPZ2w5ELu1em
1niFhPar/HWFjMJHWsZS8oXqtv4XCe7JoC4BKEfnhauaIEh8T2xDyRHG3UzxDW6j
kTH6K9RSuu/jSYJ3C6oF8QEWIqiTYEVvqPTJtZY37kaQBgdqqEbSpEH2YR4Jc2gi
6kBscAe3jPUiFQZXE+KZHPlfJgmsrV507YiS8mzyqFEsQqluq1e5EtBtJyXgdufw
vtYmo3n/k7k3ugLJ7TGPI7EW6idvJ3uMpvqVULze6gdrYXe6Qn7OTd0tbrw5nGQR
eRZ3s5ONiI2I61BgEkPMoXvIJArIIwcRiqNAoIND5OprNll7j8kgT2E3QLLUa68y
NJZjh+ADdgc09qj3PiP1GYQe8vDXgsjqQC8ZqXgJtJZeU5Ka/KDFxX+VTNxMg1WM
X6tkUFq58Bl6hCzbZZ5ydcmIGg4q/21zxIljHhB/NHv2YoNgm4z722n1vHJ/tMB0
hBSRaACtafFAGdtnywpQ1flgZBMtTyVzlXbHGNrQK3KyL+vVfYrqMpJQ2v67ExFl
zkVWRkSJcUcitZvDpCXVzt4C6Eu/AwJ9yWiXoEAKLrkaQRMlQSJSi8MPQG4R/lK9
uIxVhkchF5wQ2A0oK06w+ZtFHl02+FSa3SPkcMEm2hAasFb73EPfOIMxZnutX5fZ
sc2TnbWV2YhwGlbfM9LBdUUmcKQTmVrDfaUPFmfqpZBwJIf1UxxAqDUCIkoDDDh3
tiCUfcUNOmNVi0X4IIR5629XFd5hjycdLD06oLc7Varkd+W6yZjIbUyJ6KHLgDnH
PRmhJNDrKmBBRjywcybjJV+/bHX2Q9mGE6g4ctldx9bbW36l5s2vNaBmjRs0f8u+
En0VxPigtJfrFmAuYSmUEG2YxFJZx3BwcbdPOBIA796H7Xzvy8xlvZO4+QKh8sAl
BTerP80UH+uWEDSzKmoXhXoTpwnwp/BSJQXRIc3U1+A9ZI+Mzv0B52prQBDwrkbW
1v9RxAGiDXQknLG6DBU9aNTmxKIG8ZN5Fl73akFCaQEpmml4G8kyRS0U/Shqd7Us
a1+cl4LUl/EesBT2LcuBymcUmK/To9WWxQxWpcqmfESPnfvWdkK82v4dtM+WwPGL
/4R3i+EbTvTLl4yjXt6/GCpmSuO3tliQSVSOuRBk7+h/KPcsPRcwWpcTQy9bW+DE
sBiBVMORzfzKZokCIR5qV7RSOKuqIfQ98eOmhVpr3rFGizsZIMKgle5sX5yn6r4/
HubPinyaVhONjRoOD47l8WjmYv5oUZUS088DHWC8e026OVQlk1BEGs0+HJMxew6V
P57z7/WQq19Kd1RQWHxxj5u+OJhWGmg0/W3eDviP1vPYf5v4ehaFoRsZHTAzFZEF
+znYUar7d+INFBiclj4dEokwr69vqZ+gE5niKfqd25fCVlGFgp51nd9A6SyzhqlH
0ym38LEEaxgloCy5Ux1qahV6CqitHkf9zIsOevidQay9wKGThCpNVF5wkODt25p1
5XjxVp7Ofmbocitvta6R7hFvUMy+c497HM0v6OzRsb3xbMEdiAKvITncH/TTsk2L
NaZ8R854bayWasIjP4fezk7F0snCaQW7pFeC9IwQQ/LAD6JKU/TzFgCxaQqLDKi4
t212uBgkrWsRxuJwqnXjVVZbFlKlGRUGbICcyxZuMTHZzjxb3zfY/iV9DIAT0jCF
VqjWSsNjRynxmr9is9C7jFw1wVurbeBH+s+pspLXYKalgROOyOwcfE7MAPG/wDiJ
63dVHadKCVo16fhsnfDibMefU5UjpFcSmDLg9vB+WMzxVc3H2kwqsyjRXAJy3ZdA
hS08jTDeA5JjDQkrhMcBhu3ToUcheRMWCE5FbU5HYyW8dCL0m35nZQIBooEse+Kk
9v+Sma4wBN899bGQimLi4NXHzNi0Cd0NWHI0p6I0qThb/3Ec+fqGOapooKKAZN0V
y85/GzLx5RmqLjbvZ1NEV8ZHxOGA8zFacS350eQU1YdpbyGbV9kxCOL9MnO8bHxG
jkGJSkfNTI75QEIH5U2OYklYOpQdJjy20GR83qGIlMBtZWe4LchxbtRRFJNTVDNL
E1KLdQ3EVi5e+35BGxuZFq9hRq90RrryFdV+CW2/dZ1N4rrRSg4pmvCpppWlkR10
jthHvXIAg9QvRF+4VIH89g4h7hawTN3hrkiEM4c0HpSSWhtzmveWi4uBncHAaWNR
fvY7Rt955Dt0UfCTyH+hx14VHztdwxStdcxAzH/hq7lCZ9d5MphcVhCt0hnqVhcH
Mrn5mTyJ3DgXVajGIkiDSTCjA7W34rnFBQVLhAIB8rLn2hpUyBBoX/9YWi/zEIFo
CtRLnl9Rel/sgyG9U8Mn78RTAbqrFdDNQX7PendHee+wy13NJkFKS03898FpEVk7
45un/IifjRJ1z9Cm12UDCEN+D1Q/c8DNuMjDKgcO+3j5KGoL3PdJ0yPbp4jTyyRN
+6QZTeo6HX6bNtlciIls1RvMDFguMwNLEu7csUq37IKhlA+kGY2SQw9gu9RS64u2
Fje7/Yi5kWkviW9tqmxvTrudLdVaRZXyQswtguSNi2leR5ngt6M2QibOdG2mF+iO
bxuK1AE39Hd3lD+XaevKvir/21cOQoLg3AONOYdiOZhln3LJh2+flOiQRg4ZRPkz
bf5xCL8RWjJvTDTG7p5zHWVmek/IBERlPIxCuy1rN5iyhPPpzgxuHHD6CRej9Crk
llp1IgMm3uG295Pi5zOJpJCNiJRMJZHy8bAaLTX/w7rNuxpib0YlNOTtnbQGLbje
tKkNaAV62Uh79AdJlvhLmwI6oxz0348YrD28I1cBfPhYWWM6A8HRNuHg8NJTZij+
gGZ7b0j9WT6SYj3gs91BFMihXg24eFpff19GuqYFnE50XwhoDiJEkWaVyfhxSQkQ
lmZ1+0O7e3WCKB3ynyy7iwpo/AIjn2Cp2aIhOwrI7e6dYfqV9wwUx+yHlIwvguR+
fxZwthf23vkvPeK1J/3zFX4fam8hYuVmQHkYkV7dFBmcaFcDppxLLYWtrSFWTjaD
uaRIrbLjYL24OiQ8Z8MZDf9Ry0uAB5y9tY4LbfwaOH8tL4b1C0jDYYU3decKhG17
BRjBdUG90GI19GMNqE1C4qZ54KYOldPneVMn+4cXFR/GguWo8Tk/TaXx1Ts1Wgn1
DXaskhTQnRYTf2w1F1OjAfMEnZAI2fVk//91mxBECPdwNYnO0S3P/Oq6YG7aDuvh
ze2QAAUlxEr7TNLAG/+7ScpEvOZxJIaCnMDsaLjdVcPGkA7qM/sjNZKp3x2XtcuY
s1fgHUV7CauIMceYWuSzkJx1qrAiJPbK4LMT0Q54f9s6FvanZA4iHVRPWLEQ1XNx
Cn5U/71/c3KbmthQTGOtWn8HnJmTry1Sw4YfAPLqhnHG5cG01eLkQANT3HpDLgY7
5JLWXg+bWIpkiWCyPV8GyLrdbBlNvNBgTwD/+p5qWOZ/EMFcFJiESC/sVX4g3qbb
S+MiMWDrrXVB74mGtSeyHVtA4rXicT3xlccFNJ4/dxLFK0sSUx54w9H9OKHuK6zf
nDrd0Fhd5wW2I1VdJqPWwfEXPT8RDaOAGnOVY+Hxl/Kyiy+U7pqtvQXvqcsl+rni
MtxlaE5RqEJQACw5bgVagWFXGr5PiT34OsHsX3NgNS0rM10rJCNBqgSCFFz7m0hu
Dks3/W12yQBlMoufNHBdcVL91cMJ2v9npj8EDPvAgCMoFIS7to4AAmWBJsF6VdG1
LR+JQ6nay/JqI9BZHUrbVeNLBoOs7xePpUFxrrhZ5ys4e/3virxTDnz0T34aQRTS
CnSAyM/FuklVgB6z63QBkHjP/7eIDApd/YUju44ZH6MHmXgyK3yjZWhrx8gi0MsV
9CrGXQ41SIE40v0LAF6FpYH+wmcWjTKuTgAR4Jq2ZLOHSSGHMS2d9DowXjz4wbjw
dm2J73mdM0PXZvo+r9K3urzcIAbC9mvgWLVTQdX32+9esG2hS3SKS/KPl53vvgUY
GdMmS06UKkYLdV0vBRKRmWMRZ4K5NMiq16Tf1VAwet8BjJvAvmAFdbojhPNLv7Ft
vnrG4MAObmmuO4wZQaIPSStNydd7T7J+0ezEBVjODfIGtRkEfpjX/LCRoxJ2a7X/
hk0s+7Mjc9oa8PPkaVqXm4E2hmzC+8maImc5Jjv7jWNSAW5G0VHdbJcHvVU8XXsq
0EiJgjrcDVcuUqHQaShr/P/Z4KXL4Cq6Yu8oWCN0bwXLjelDErmVrs0RxDDZ1zEr
HTeXH+HLNB83oYOXDU2zhIVOg17GbhUTxHjMbzkMKdymdBdpxz2xmNNPMcJ0MQUq
ZmRlhQJtoCiuR5ta0hp9K/+C49Uf/eBS3DYnLaapovNMU6sIOyFAtCjgzIX+hfyZ
D1ntUuxgCvVCL8LfjwyYOaadRHdGoqYR8D6W1zqR8sAjjLqpAQ0BwQbIdPAwLyLH
Fln0FfEu1pSrwmo974vBKJ0ykxBXUBP8AYxBvbod0RZCjLijxkslFLmwuV24PpS+
4923CnC/aNScy4T6UIsSPkUL0HYxgIrOjqIfO8ISsqGRvVmwMzGuY+5UUWgXEcXU
PqPR8GClMHJ6Z6SE9DSio4uOokWioEF7fDE39IW6xB+kfEM4oZha7/Q6VJg3zaGM
m5MCLtvu+8D5vZdCKCkGDTJfKs/gzE83dEXc/zj9eKYMIMaFqHtBQxzVNbyCSjpg
0lpyu44/CTL1sz9Hn3i9DcSVtfzXLzpKICZYUbfWvJhIAmWnMv6oSA54TShLidCn
/ewD9dwRMcyCXPpOwZ/iPqO48JgE+/j9/gdzuW1X3tWaqssK86vrVZrvred13bcK
1+bxv+/ol08C8+J82CJPYkUzfC7iwY2ub+eZyvERRwmeX+AqzAK+sPNavifBr6z7
oEL/4aEZuOZogUoKxV8P40UgNIkh1V7S9BF9bwFWWV7WOBe36RE8EAPU6ueUnHgx
v1sWl/956j07dlpmHwa1u3Ew1ma+p+EYslnMPuoNYin3n60jjq1Fo9NyUiCN5gSm
GX/Bzbe4WepxYHE4QXQvcYxuAYccSCjt7i5M4ND2Oimq99I5guaVIa9DcaCOGxhk
0KLK/nYGbO3XUO70f4oZ8UXPzz5PAH0/L3VGsyxcoXnQaTW9PHDP+RcXeJ8uwFBz
hXOhls4r/3a/6IK0usStIHtIDXN9xdBsI6pvFqZsYRFFr1HwOfkwoIiEgnUPtLRa
mTjF1JvSVIRtQn/uWw7Hfli/gbSsQ2B4prjZN/u0NTrsLdGft+39d6EBfCBxm8Xo
/Vkn7aMy4A+Q9SrTF63e8CwEZVYXSuji8cukiKj1la6MGPk7Hp3UnaYNnhH3va3X
pkVkw0BhJ4kPM7xfCZIySIAMAF0aG2omlNlwAk4BpXBsXBR4OW0E1FUdXQQDScN3
c1qEpaMqMIA+bkwdaJKj45bSa3ld+ZhnGDhcD1hplo8UcwTbdplEBfBQCZYqMFIF
T4y+0Hl0ceWdd8ikxKuKdj9K21jKMGZ3D7XS97o3o0JV1JhGWRjqUPqMgNzvnXKF
HcXa5H0w1ObO5zVIQC5ovQg/Q23vMaFEb7MDDs3+KO3UcK3WOvQK2sj8TfJd8mEQ
St5mDDFdB/91a5fH7kIGrXnFjozL6Ub6Pa0Yp8ynEIP7V6++3PQOZLOtdJLN4kk4
1R9OTBs0r7ratr5UENtk28l/xUj8BvWMs9oAPDjXCvjPDAhQ/H+Xs5QZ0+Uksj4F
ncezL/re/1/y3EqO9CQ0XuOeEA/mnVga8VyrDboMPWh9KTSy+/Z9J8fKiJqvrOq/
yguZUdZv7XZkbRBVt/zTmTIOjOLoyHqo11UuhFP55B0DNkWdf2k45A6/UxGR6LwI
DQlQg6kZ5fH5X7/9UVL8JjC1KxMM8OEMZcFnIwZhS0+x/tFvszgP9ZqoWZhpcXnh
0ua1KTqLiZmvUQcEm/Ob4Wjxe+iG3qx2apZ6QYBq10+DGSVvFGtOEPTU97hr4f9f
u9a06W5TTgrkwg+o7Fih459Y1GpNLgHUkHtG+vNDrTx96m1f4ExLSphh2uowPfYL
0nHj5oyS+U8ZQSbW2mMjytAIaqBCOOt4fASyqL1SDx3JGegg8yqK/uQTemWFG8qc
102yEIqZPHF0+3dd2sfcK9BmYaPYl/98Lj6SUlh9q0fuFLh5O5bRz7ZyK3XW7Iif
sF5uwE8Pk1wkyqK4By96+ipL8QYdn25JS8wSeRT6rAN8daWQ0t3TxhJmL6fwWJyD
MDmMCrQiXK2p0eCTu05TELvgEYAWl/a47Ruu7YvofVB6y0F5eUmyLWs07lnmahx3
PvtxRw/1EIYleLzoRmLVZVVSIEPuL/7TxqPc3Bf+GMpp2iwpumUU0mkGK6SkNNJy
xojTwgemtrhbBRiozqUjE/Mj0AdZQ9w/x4hYHGmSgXNsv9VnQ/cqKraOR3TgZVnK
f1Fafjto9teD7gOP9hR4i6t4NF1x8BQFNVG11FhEgM8DaO/LriRaNr8EGBRQeHen
rdQmcJKhDBHNA+rQQC+v6nsw828FTFhxzodloTRRQJTXnQrnDac0ADtLAWXZNPm2
Zros87D6EVFk3f260CJ9fezVKw8gMqnVM1jl6poa8GsJGEBpLIjFoFi38r/URFBD
MEp0oBO8i2BxpsfQTyRL3jbBrbWi/O6ZUQckfotUqLSjS7Z22tC3tU50w2zKqhSZ
2fMTG6Ik/nATVP0BTowdl6JrZArAEJIFBcvoysSicd8mUX+xSXtYnqGiQHCGo5Gd
GLU2h3dNhaUSBc2FAA+NlCQ2sME79LUUIUco1yP/CcMh3GdmyUaKaWox7pqRB7SP
TRr4Fyf5+pQvq4t5Knm0Vi5X3tE8rj4xduDSFvq/D6fkRc/GSMLbWPsh/xZ0yc8Z
eEIgKSxFexsVFxVIb0vR+vcwq0W1/byMhxKuoY2mEg/gm4eC4zqnxMnt3gGsucD5
rDLLjn6mfrEwY0jEekOsnMLXVd4apSEjFTMOv7f/of5qzE8AwTs9JE/9fChHMth0
nC+J+3aNfwaP4KeZDYeEy4YuMGr30oEwrgEKYjVYajsI+HCDe1lj+ZW0PsDNNbxd
5x6rna/WMS8AUeSqen9jvIG6KJsA78JQtcaLLiHboTxRCyYaOBOAeaLr0LH5AMhx
6eP6qlWDleNCguKa2NMhI4EcskXYyh9L5z9AFJZYDxDgRJ546xb+ZaUQI/pz332w
I0SQicME5zDzBHiUmxQzs7IjW4/A7ta3rK4bPhYfssrWmJQchP5w2Gs289qDqvtf
ZmNBzOYh2ov0S3L20kkuFyAjK3ghBmoR5I/rtnuDpfv3ANy8ekFmKjRCYuLRe1GX
BtYdPKyW7eJsiIlVubdYfevYvKgZiZJhwx+G56ziNrXxjPLdsWFZm/Zaat/MNHKR
UvqCcchTbp0qpl7Id205mLfvIpcjcCRIj3PFbd5jTKo+37g5Wy691+lGwRfpWD7r
VVORbtXPydqz/lRsz5jcNkij6xR9GY3cL3mCIiMTSVk9GKwMNoMRj+hawCGRV7w6
e9m7szwAaIXSI2aAkQIO57zOqJ38gwzmLFE9IPqtRT5L5VaWtKs0RHS+zbFRSOU0
FzTQ6YMBrT7JIaICi2/cjfSWibD1P2S2/yE5n3m94sFPMIQ/yZl04fxyQMBKi3gM
djjVjaMxjye7EAKdAE9lgnQGNrw9dfoN5DZDk4Jc1y1PsOYi8zZ87+begZvvw0D1
+ShwgOIqntTEeO9Yi7F2NemYbcv1j1+loE4Iua6yqWpKv1gfheC5RQvpMlOLsg92
ShZJX+PyXOIBcJjP7tCad9GmLqPATQqoFWvvjG1XI5ZD1d0D1zK2F8YINKJdV314
9cFZJA9T/bTTluJVqkkEgF7jph8Z0k8Q7+y0bPUccerNl1NBayPNqkVb73Rc5ke5
1SQ6fAx1cf9FN5MzifCevy+apS7qLDav38/j6o5i+M9v7MmXy9ty1ztI5knAyB77
cwbXsw1NgTkH0/DtJTi7i9KbNRGIWo/drOnlzS8t3EmrQluRyUMJ63K0lnxQlxSe
3LpwrdMWB5UO3hxZNXeDx4mDmObgWb6ZgAeI9rXpMI7s5LuDNEKKBDVb4wZzy+xz
SR3zrevoQXH49+vXk3A8D2rULix3qgJZrHrzHAFGDXFSUL2eQHMFzYuLHlJBquh8
eaS3F8xh1ryccL621DZgJ5R4rS3D1kBLLAjKknQQeJTR1Pv3eGLSIb8ejHKXfT1+
6ML1oHNPYGNlheCGbNdWsPXgv500bu4PQquFJhrpCJGJRvrB/y65N0cvT7pUR1Y6
qO0G6nJ5B3UPXInYXQCEnk4uw1afbjuZ8zY2f4/LXHZbeZGCoOwvuC4W4RRXtrmD
1s/ADRML0hzStXFoBk4TKrg4BE7/QrW/Hw4++VyPTPobyGhYOx4PZccKAdGaUgVj
BjytPeH5IXysaEW4GLbBOWs0tGb5VnQF+hge6dQigbZ/6HsL4o/2nKpdj5xBBAJ6
Q63Smq/iGSsaVtN3qrTJlQQ2usDHU5ruda7LHIvhuLlpBqxu1bxWwDL753s97PhX
g8I0hDoS5S1HdqekIzm0SNkyhNSahSruuCn2VJUkqEtIP08OMU4vNhS7tB6G0EeG
Lh7r+8l+P7vhhg5pqzMDrYuTvim2psPOhRXReKT6LSIYBbFZ7HL5I2Yzi5+nTT9H
McVTFlEUqiO2MF0hKkxYYRMK4wsiBQ44O067wRFVJRF7SeOpN/GZXC/zQmQxwBig
8n06vvxgHh952j4RNBC41kDgztAAX4+CE2eR4BpTuqgNCavczb2p+/asuMCxlLBN
T35qd6yxREdTBQ0E/h5vihBTOdksk5y5zX41PJFHWnqiak08wTig0B2W3iq2NekX
MtAGF57OJuzyP0qCu5Tk+uZ6XrB7LmvCRPG8HLkD2x/FI1cEI7c43XgyuFvHHTRV
mh8TPcfVYMxiEqguLtxYhYMFRXm84hMbGg8n+7u6w/v4rMQ4FCwG4yL6MvqrCHXf
TZz7N5sD0A+h/jgaCNjdRWHzfHUvMvROKksU9ZG/bafaLOwd/SqysnCaDtyk9JYT
UxTlI9CzbdkcdKIsKROXrvqeSAWvGOWKCZv9uvmJLY2xr3Z4pTT0g3Q5BUu3OvpP
ZpKZ9s7ETTZbM1y3H7rtzkEflHBe0AsAauB75/bMHw83dBuWMAlMY8678aVj/mZA
HeF4ud2zGQ/ghFp3z767fikbiWBWIYIAe2Fvxa+/1gnIqYge+6GgaGIFZYzjTkUm
XUo3Gz5+eQHdKD3i3LVrQ0O7G+X/dnDTAqPVPzemSYvUk5M/55H6oxHkkPDw3qgj
2LK6KtdBLXjihPoGYJxdGGwwgrxBO3CFr/cGPSvUMjXMGzm1bS6bwljnXQIfkHDg
fmn8nnI9on/L9qTGhpCgmb/o2D9wIE/DDyoCvIepP6Y5OzJGtdp1Arlx0N77tUKf
oo6ERLeekrEMlmN4IY75CON7rtWUFj+Gf/iFxvX8x7AlXvytOa+Vv5oooB9GMXlm
YQpTrjKBOkPYYhy9zorjMBD8wzV34fCG1HxDowAx4RY6BmC+T6r3y1XgmLGL0ISp
u1j52yQcAK5Q2eDpRGWh4LbMOmndU1SQQnccOeVE7wifNht2fHc+BA2PSm1zRHpW
2dUcQHwHbixuC8uycdFMPRlS7453K7Gfbu6WrXYY5utJAIeSc4+S6uGfJqpdb1Ls
3pZKYhi66Mn7NNCCkyBEvHVThVDD8SAPKkBfgMwDZbtFo8sEgERAKwPnY2JAxpU7
MHt0cE9FSKz+/9lFM0jn6gtkB+5gfl/lg8GAz3eWeFYz99Sgi8XR5Evs5tUoC+hs
v8WscDsh28BglWmO2C9niqcz/NN0WxU4Awy3aD63nQKMpFgWRXJD0r00uGfL/KZY
0W/3nfwsG/SXjmZLfb29vB8bvbj8UL+ZA/klPNVMdFyQLbefMh8+qnNoKMheS3nG
xhOeHwHe/Gw1MYrSWDB5VB/CmPUk/ZRb2Tq++1LxUJ6ur+SmuzfwHCXQ/vw6CfoB
pXOo3INoB2ug884tlUDHf8oc5BAdCXXQB7LwcMQI1oRSJF9P4+PyI8fHq2tpgvPi
VnBKKgA+qmCnrGrsOEvlgEgI3KnCwJ3+2Q5Qo12UJQ1VweFYdeBd31oIq9/J9eB0
cJGWrIV99RVVfJiEkcWlooYHwP/vOtJDh2eo0IkzhbyN75AZazhU95ylYgq3cF97
ei/sitZzo7FalhHAo6FAaQDXNFgUuCue1i3dCr2ZJ34oIvH/f0HmsSfYDmAzhyCQ
yP2e1I58Yy6WWpvxT+q6QTYk29RlnjTzDLjIKw/tpZShxVZtZL5tAYy/kSBMoReX
8alcgUxKYPa7lkWOBnZFGCp+V/RXj1OZKj46GyQ46YbGe5XwJns8alpCeN75yoAM
ntjibJxNyMwaBiW7jbofKENia+B6ddl6D+nwpiwjueBE6PTgt6YzPjwUJQc6iMh3
1SXthRuIdfaAcQl6H4SZ3ZIlcrdWWBvCCVqLTpEN8hPnyp+Hbg9fTTeLzdqDnaH7
A5WKg0M0w6KWmAYb8isBdmXRwGlHGpu/D64Hidfc5f3EBvPfess81eJeqFuRry49
hxasHNnTLg/GDKIcHpjgwtMD3B2kVx0j6r1JcjQ1VKer+HpVbJ1tUsxvA93lhbHh
6RXeWKjqFaciD7AMSy3Sw5kEe6VpLuSnj1FlacttMkvsEBnMjBvWRcsh2skPjNg8
IftbKKdKoKHWcWa/wvEQdeEIX8Qek04focqGAkuhclmEaZ1w3MHY1b49WaxhiAvp
pB4NvLK/XhpdozlhtMtlsbvGE9A3cGJkGHGIp5QNOf6mbBoIQjXM6dTH30jlTsEz
s9Kp13zyPlQivMdmOrkrbCaB11kmgbDPGzHEsrlTTgXDPiszImz1na7Jy4GHcnDW
cLIkPZN/aGPR7EPku5Zh0T5x7cdCEtp2gBvuECECzDhYmGjFop3CC75q5jrAnWPR
QhrSymItwA6+bJPpK/L14SZgMNT5KA5AS90w1vO0bvwh/2EOvlDZSl5OgjfaRc81
4cLhV6AZu9aaIL7NggxnveYH9yybxsEwS0kCtpaMb6rQ9ZmzVC/Kv5I7KJ+BywJY
QSHRMH95q+FoPd1RovzkyGRTSP4A0M3c2rpqrU5V6Srw6SSm4DmDNBx2iBf4kizt
8BTjVpF9YkxRTN0OQKuATDLPtlmM8F2bX9Eh+IAdjf0gwxHWQ9Rr+8ZV5dJUnIgG
uRgi2+bES+3hQgMkaNu9nfcPfnbZEIak6kTxyBNDWJ6fn6kbxbadaNGcUEl4yWLV
fKdPHY3/SfjJNneVyBiL4Dri32y4J1Hdp0Xoj8ITHWWXhNFDy73aYT/bHLAw7bty
n/7rUpcGaGPRTYjO7MMP1J521QLv4dgN8s3mW8QLumyFqoadM0aI7WbY1sIJTBN7
oRbSJ8eXNJ+PAit7dc3Fk7Vg5vxjgJQojqTF/oOx/N4LjFAlV8Xm12aJgwKq82rB
i9EwLE1VbzgWhf1ZsJFgExCb3yG4A3N2kSZ3P8sYtDW+Sc+BRHLr1khqagKVasbG
BxJg3eZcVsI7VFo4beWQNtoFMoPv4Bs1c43bDqVRwTrCouO8JW7Y7tJ/kOHdbglY
h89I7BlhMtFKjUC42t9uCO00IW29219o2MYQyGiDHUc2jpSgRb4K6NDKgc7K6RFz
UbwJWnDJGycUT9loxnJ0DcXSlZIdXbE6x00ycAm4J3NBLDxGLxLZCQ9nny+z29o4
QchbN+GxZHakpkYyH/xhPFZEaWj/N8FStJ7n/hA+/Fl0o4dqcIJUIcVyNqle4lhh
ip7IRRRjYlR+O51Nfbb5EDZBaV7vRXX7Cf4YVp51/dhQMH4ma48W8MgIi7jpQj6E
ErDlEU3Cjxz9YnoZq7upNHObIPN1SR5ALsqZXkUMHUn7hOQQ5hFVd3pNWQCZ2xZk
UbvxJ/zgd3YJc6xSKJgMBFfP62z7N6IyjXmei1ph5xb9ily8i3ddXKYSiVYiwPZo
8DJVevN4hEFJ1H8SspVblZslZMENevaoOA4r99WBCstcWX7TaPAJ7A2+dTLnbNf0
MjWGJ5rCLY1NsaZCoUYxHcUTTm1OtBhmbrJgQQwKJrkcI3TR4DK0L1LgZE5ldKOH
yAaj/TJ54U4b4sqJMGcrgpfdnf8/jnjP6a1AxNsW/BVXNLH6Fw+cMB0V+vD+BsLX
LloahkfXv/jID0Q4UGrX+Pil/FUBRtKm45vb0mPlhEQb0sZy5iqFZyejeZxhJorz
m7KdNS3IHuUJMkaOlIc06ZyzBcptTQhEea4vqFLMDsyH0q8JJZrjZlVXc1sw8FGi
moycP3NE2hfHEp36H9kmgHz8boTw0+H2dNJZVUzZ7c9DcdAaYh1LEdG60yLQDhJn
Vw336iqGbv+XCdhI8sbkGndpj1cN3kYffsJxW+0b/ajRbM4FLkwoofQXo4GTvHh7
d9DBtXK9GF4V9kV+qmginp/OSj2U1eInS0JavtWa6Dk0WvMNJdSOOqASc08PvW0O
w7tfWZzurS3x9SwsZB3dtOjkRmoth5xB4urFy54fF21v7ldBoIe1GczTzvnpSaNO
2vywHF7IKtiI6cLfPUuth1HmFlZJNyJN6BbL2XhhQwOFFPbAec1aMoQcSEv9+pqz
Nc6zbjQdnbfEYdpKBP/PeDoY0DhqVLsmRs7B2V4tHLTD8xeitmUoRHVBRep2Wl0J
0dxJaYBA3xfq4TZWi2SHem/fBRF/YJjiyTYCPLOhUcXw4/AYPiflS37PzWdRYi/B
N/3zvWLZzlQK+XyxXM78+89PrbZIIHVmTQMAJUkpPJcvE2ly8X+qLJpvdB1rKu55
1QR/QkJ1NSD/idid7ftkBdoa5C0+cU+d8UCsMEaRZh0n4GylY9MDzXiPy8hfMheA
EWFuznyFWjOz+tws9k+rzfs4VXnuc1Pn/W1cfiPGvtb9Nexf3r1KdM4M42R9C/d0
xb5MDU6KFRgWd1IhGr56uNCJZgz+FnaBi/dbOBoccb6QpBUnGGJIrH+vs6oLWAsK
7HoFvlO0psUNuPqn047Rg5bFQM7XSbJbzxI/fTvyh774xS7qvcBkuTuTWxVl8P98
f+jhcv4hcdpMqgkZVtes9HtxW3bhZ+9H/M923EFbs4Um6Fz6mGmRFMUGO/Xt/Ben
ouG0JjAnbGsoQdneDMojz/aa7Q7/MGjXsQMLnllIuzX4D2ieWDmKuhw62OyVEfkn
UaOGCDjhyqxzIz0CEzUUJhoQAQxzFL845l6GFKS9OFKgYNElagRJxvn0zhhJpDj9
6vJC4yOlsGrvD3KqV9j86jCmT4GLBIL3aN4vV6zoNHJ97apYhurC1w080NJiaZ3M
uxywZUiuftxOWfqwVF6ErLy1soXTPKAGYBpoTZJqsdOmLvCx0SB/wrIpIqrsF/KN
l243Z9Vz4MRXMdJM/yybvhIsf/d1fo0IOK/5vM/bL2QhK/zemeHWk4ivhY33m731
Q8vCxdmDsyz9lExznLnH1iBT712rGm2OivHVy4OhjB+al5NACfXcHdoeHw9OkzWa
1t2aT5WzCl8P9EX+3vLrai6twoDYO5ODafpBR/+VcRJReHmRchRudIU76zxps/G4
fMIeREtqazke62SOibIiaoyk9+LA2i/R3nyKNCFX3gz0yW9wLIUBBMFYmNVejR20
kvKv9AqY82AaoiYKP/yGmuR5Hvw2eeKiy8J0AcFdYJecNUNeBIwPXrhGdRwCkxjZ
vifTxEzvFg3g2u5vmAON2smFkxnsjHAkrW5CgZ1qJ1WgVqczU4kCYPcA0pIwuY+V
r5YNVTlGXcxMGt51px4eqiLaTN8ECsBJU/0xoK7zF9qNftuvCb2D2SGly9qHHpUN
2pH0lQ38RMABeVIgU3CJsyX0iQ44HOY8QeLdoaJvnd6cejyoSrx2ycULT6hqoYT9
kATIsl1algO+enPxLaqguPZN43+f9gPyZgDJqTV1tAOK2S6HNheRa/psHpSkSIZ2
1gfhKlpqGTwebQz7h6DtBPmSRxevv7GFxtCkWOYpiax4205YdDYFHhBcIfCTigKv
cohsNei3zIN65VxCSA7n3GPawnqYIEmHuxnEwkXm5l4mc8FEaKvCpWu4H1h+qi3n
3StNAq5h/JjUb3y7NfVE+1Ef5mHB/ROxMBV+T+cdXG5aR13/R+vFZv/o1AYhuv51
AHBeEkMVrNG7384rbnTKc1fsz0wzi0kgc0q2p8DKKtILcMIyqtIkm/xi66W6nx/c
ItQdmyGUliYSyiTfJr78fVl6DomaVn385ZZGK7YvJJ57axNNRxL3k9cJN5Cvj/gm
RUqhnBdDFFjOoATCsO2QPaAqddpt4WTwHa1Iu9YpWFbA8hJ8+QFFpjnuchJ+jIO0
r2iRzYNXD1cPN2uf1Yme9T27ywZUxA+PWVe3Lp3PI4FwD+lcFAgVaBN8BgjqcO7J
E7FqZFkGHf32jqThLC73USBOGZ2jOiUgZeAAufiuc2ZJf44pggS0+Gk48psXcPXs
2DAD0wajLncw+2xTIr0Co5xQmQk9foTSnGhR/Xndggf60LXejbWEBS/2zFZ5VAKp
T4DLesiqWqiNAjWNwMCOAELR8DgKzLc54ui7dugHmhaHVsF6ALFHgQmu9hqhWvcG
RIFi2AtVBqDeo+S8TzPAm9qwOURnxboQC2rOc2kcuVK2YYklpSHpJrHL05mPgbVN
OMdUnZ82nTKfX4KQSLDduI9Yt3osGnGQMfWadvzPHLE/Ns8jgNKxh93aid+EJ0/D
amvIbpHtatM52dIQl7ddheh46/hA9SobZJznvvFvaBW3L+gJZkWQaKThd+Ai/SxI
FZ200nu9phdU8aeEnZM0wDhqlY6D7ojB2ksMW0ZNJd4+GEDa9iZrgMP8eL7X5ckh
vF2XIuetahnorUBW2R6Gl52LJKY2sTTA/vDbzNuZ7lq+VVBpLQrsLuP9NRCBIzkE
xSTiOLdEJJGfKqvBnNUXTX7/wrsdItEEwkhIwpMxS93wHOxLkU9+NxXE+VmdAysc
/pouSF/Lr7TemKld2nz5ff6ZFNJ5zbhOMwUTHSWWRNOAMjFDaNqtuder0iA86eb4
xLElLzjUpC2CZaF/rW8Bny4UUhBQjknavvP06M8WtKPX8pdnKSmlMwsB8rn9xqJ2
OwkCPMwvUmLZvaf9qg31c/pdjmmqx7YUOoAjG00DZb3rCvzPh+uitH7xDbAaa+zC
uIcYoZQsPTVvzf2IRsV93S/YxaEqrh6m7P92wiIdW/6MEjv0iFWqhijGHrFMvp1r
ta9ApJFXCFHOiRO9Am2zu2+p+n5FanJh9FBvgAtwPBBRNMkFeQ2O3whU/ig7/LVO
igP64BQt2x3PY9/EaUk6uh8crA1cZ6OUFj1qR//HgiIi+TROgzvIaIh8vF3JGQg1
Nf7N8AMB/kf8twF4G3w5H4dIkJ3yF1vyRbzQe66/Yuq+CREz2/asbLQDpjE7pn/p
hAZCPUEXnl+11+t0i1E51I/1OHs4lXFh0x4nUyMZsQARrcPbfyQxP5gnQEaEWll4
W3zV7h+Zp3DG/1VctsMCxwS0E71u9sEOPMBf4zIxnvyDei5V2AfaU0Bu5KDilxTw
u2i0PZJ0WrrmzFo8ujfGuLHNynQ2Al0YQiQgR1gYbrn6UJonQmQYoej7EHNb/EB+
g/GCb1gyj//ZqlbI4U0bjCAixq9RMtFiHub7EIlLC0JId0NIfa8knK64gKdkVY2d
tfOMeW6hyVFl6qJmqgCQ/XsGL/bEL4gp38LsLiX26ybGqFZqOUNbuZuAZNGPWqQl
91psJTCGtnw3YSCAw+hb4bTiWY8VxnZ3Vk10gL+9kKbQUUL3tPHNAM6r3RJybsXG
9hBE6fMYVFE8TxzZpki3zgfHPrl/hPZJRQX3P6WJNpxJQ22yiGjz31L7Msl+T80S
1wJf4FvCqz5i2tVc702sNpHdmI42hrTV7Xx+k+7GgN+46GoX5hkmfk3MJZvqWIFV
TS69FYOf8VTWrA3hqKSKH7OykWexJZqGurbCJ9Te2KqWKAmMTuV2ifUbFIfoa7hZ
tixit2hdNP4+eIj+z9OAsMhiYY/zv1XI3pX9/xL0xFGT885eqa/hGAp8+1BYVad7
S51LZJqcQLwDcOTNB9YS7VNmOcUkWYkJS+Cm8mf9aF4kiyLAtgAnAoBUvGv73Sbu
+W3lUUo8z4SLVoGg0eWxxDT1qqbltTvoZZNxNIhJdfFXq7U6KNdoPhw3ht3pQER3
vpGCfXBq2mVYF5/x7KX1MQot7i2+eiz6Q6XKPcNBpfWPU3B8e17pnk8tLlpBTUi0
cElUs7MBJG1K9+OUCuq1faV1s8y/AV5KT3Abi9L1ptrUSdWzfM+nZZLsnwZfJwjz
3wVTlK9RWUmkPCXGi1Xy4A8HcWbavxWPRFlQvHPOHIQIKWew+01MWJR46qjrpMJs
t9z+Nks57qPU64YIA7JPPzYn0svaT+be4VNuSfCLIdULXoAxXR6b/vuUrSD92ycn
pHzUPMCvi4YfuqN1N/xXJbaCZToeJz7GVAsCZ9QzSGDjV4zganjARjvd8WVni2X7
r36xGKwpXeMs/1Alp+LyZdFgCc2boUB/lAYAbW5OTy12WBmLrAHEdzGOtN33C/sO
VinCr/EodOrdSR5fuLqN0DoeW4Qd0thD1d+xLpitjl2vCxKJnbj7qMiuZKuhbJ5F
PSlkE+LTqmLuhNFdbAgYqfgk078fuN8BgXbC5jDfd1+f9OkGDUTroPl6p+QtCYAD
dDpPFjlvhXBwJm7DV+S5+m5/HILS3/9o2QInVJ6EPwfNujTKof8tqQDWr0bZBh41
CPZr+xEYG8yE2zKbj6DwxKcFlItyHLJRelUX0YjShfAzAftrQ+vSCvvDFeDaHbjs
YpChh5p3VYDfSxJEsNbIjKOhp/n1XVvSFk9RponpDLiNaFjnjkRDkPdOfxmoAYDS
jljmcCFSQtyZny7Duv4dg0OwWZr8vfuyPsLySkxWtCyzkNcpFrmtHiMwdD2O493d
mbPdw85Ww/kLgz1IKy8sVvK/vdaHPnoC74Ce3rHWNl1HNajH0/1SVwvurcHSLKvX
Un4yVFAWKTzfFGjMqRq5YH4gM3BNt9Zmg80EVhgSchCwqMeFFRLCChn1NE7sjeCV
FuUlJAqwgmW2NIP3wcMIfkAvmE8DpBNrPeBdys5chElhW9kkBFJFBHeoAMdtHE4p
KYMFHZUs2FL8GhIo5taNy1I1VBcYFBzKmIx4q+LybQxmrbKvFZ2iblO8md73tgYg
EKIRBCFpU5VuJ6U7HVWd9U6VXKcbQAPKSr8H1AWEPs5P2gVuwuVvY3BK/PuVYNbW
Ry5HtRFu2ZwOPuW7MQkL3YB/begbzrVZkbFF4NniMIZfl/7cAxiwpVNy7jPPnE2c
q/Fm19B76CcbxIZGmEq5MroYaqAeYmqrp+HPgvDr8fKIaQlGYZ9lHrCvF4szW9iL
WimDkdcNwGuEM+/5s7ZcTJ7Gn83AvQgxfiO7KBLBuSAp9X4xRCx4NJeXH8zN5Z+I
/kWXMZXD96QTlGacNGclx3LrPIeChituQA8hxIy9aVISS8jRhm4z1tMSRKBmVI7X
fDicEv6k9NCYE/kKF4yfyvtsq56649f+0Fb2cKw1ck11XMUGDtGWw5Ty6ImpZvH1
gvFTd6navnUPG0eOALdibyGvifRpc34y19RqkXqFs37DJvMlrfBgCQSqAVB3rN1T
x/JUBfEMIgCMv9nxRziNnH/yOw8GAxjKLHVLPYBkZutrIDE7SlLyQrS4rG8GVt5m
bxBUlMjXe0Id2tgRVc70urrv1zpGbTcngVPLj6dWaa/QxqiA3NCU1xDdZiCDVfzL
tRBRBsE0Q7++uBbt4v/ZUHl3yImMY69LyW4hMrlmRoHCreKYKmw0WKtpaCKHwrCh
IjivPKLPDR5zCDwMRTxNU8K9VgXufq33sh7FH8quSWMjgsaPvd+yx2XSHPcb5WKD
ynb2pvLFjqQxC/7V1+DzR6wiwhUNz/W8U8VoSk4aRm/nsbdPEpk5gnisNILEjkCn
ssXJ/aOqCV+Z3x3OEm4Hyo1uykMuC5/1MOBOeqRtY7fpF0hUfWGK/yin8r6WoWGf
B2f1jxai4ukTkqcNCZz7ZrooPXsWspX6xYPCp3a0WgAh0QXMVxXm7gCr/o2S7GWi
zER09zpvGSjs0swYie7/P/UzgLCrGBmFYoFBf+sm0c7wF2kAv1nTheF/jxXuF2lP
BWENnEV56QQMiTiaKSUaolJrfNtntbN9HLEzR6SUFS0XAATLIHz118ZZWt/qBN5c
/AecBXJhNw+sKCjZ5fzZzmWTCptAcBV44D1cZyMu/CjYa5OvDKvP8+ai8dJP8AWh
DXPyZrSpW1lwt4Wsh+pVA90SexWbF5t3Ijg2kKfTL4/2Nx6NCXNpGUT2Kh1SJTcz
1votjdfXQl2cS447a4TznSmBTUwoF33uFSjYtddiqhDuvzyELc6V1HaK2DnXbDuc
xB4v3enEF/+z294hhfJ+iwEfEDBxW8Qu0hT1aJM8dKT3RtksA4GP80VeMlkSaGfl
ln0EHGYxbvAPBu9xvpjWu0DJjRnXVMwlv5bDmKDcRjM5+hYqmBQaQddIBAnz4ojM
VojToU6N6/XmHXRWJ1ZLQcO8jXosDlJxIK5ENRwzH4a2/pceShXHVNngLSrSP7Ht
rihM6rv4G3RprwaKmQrCDwdkdE056hX7bnHBcAoKmwoSR12sQwXe4kG28mf6mP/r
OEuIODi/m5ClL7fl7qLoQM6oOekHmgjZ7VULigBBqDCKfgCR1R9LnLWT8w3fEel/
2ZQjQ9+gMZNLBjGaCv4rK3XWpuiiXUL/kAt/L8cY+ePo5uKs8eyHBq3uB7gYE/rO
rcP0cvdxeIPvCsWE8jKoYcpsxECkib5hidEiDDbyYU3Cd2so1rgvC7AMiC/7sMV0
gl8VPjgIJIg1PCokhrh+4A8Go57AzrrFnflo0kzmPCqh+wpMxyo08eM5T89dNnf2
Mp7lcRuIvcxMI2J2QpaqU2I7gT16T3o9sfsnhOMjHm7vfibMXgQUDO9lwT2uToFx
+CrfQ6LKuTibxCnUBbb/4y+jMeXdJ9qrOHIf4hRbuDGJYdULUMXNug4vol63cL6u
2FqI+sGEWZBGsBFEYaWQlYzQ3iaDoLfKGgvAA59iTm6RWqD1Nz+Rq+UbV/pq78hr
o/gD2L4m2Jnwu7lRE7NbcbueObyURQiwmInERnw85x84IXZyEzzEhx87f5Jt2Skk
ElDVxyfcSYlIghDMZqBOsnj+kVzkrd4Pw6s9CNcWO6AS4CXN54dFL4vxXl+6cGKQ
jU5fqpnaGWNCYpveHxxIXqFSNLzRcfSWUN/jo3IUosZBOZR7bR0XkTZ1qKmOhgdC
b2FEzC9bBzKSMalb5uuCpt9IHe62j+iOstWaH0n6LnkNZ/up9tRbWmsNXP6FKo+n
yIe+XDcUfHPSnx3iItvkJZABv7EHVMPMROw3AdPgK9xoVO3srbCiUlIbVgEVhMSG
yoJRJWanySsyNa/VGoVyeVvLvZ+bgnGGyIcSkkWCK19lz8PlSUUDAxT4LFMeRKkQ
B+2l3dCB8EJO3/1jWQuy19xFCabAm6Htfw2hhfhf77TvWI15kVeig6UZArxYVZAr
QD4mYRJvEGMFZ9h6rDdsEZZUHtzn49kZcoUDpRQcbOFHp0NkwFw/rVoodf2A5VBl
5eFi3rIdKfSZfLsFL7+Yo2VcuM6REDnuec6YyvcoDJVU4/7zYLsMl91Mky1NYkSz
MsfG0TGJeHvUGkA/kik3Ds8xpIezdsjjionE90fYP/1IwOn4GwEnefVuHHzaj9Ke
q3Q4T7/hmTdtQJnHi3ZQAobaEZA+k7uCHRyIC08r9/OJRBFP3rhkl/D+OTmDEsnO
PpKeSkKVd84qJp7Wd+fA+pmkNb/th6TgSyMV1AXaq4SDzPfAlgJbhJK43ZS2f/e9
aiKVj7OwsP2h9aV16q5PS0UOWUdA1lj/8zHKfiA0aYrf1HElr4YEIOts1Ovm/llZ
ZtZuAvYuxh4WBqwFSGmWYKgDdAAOT8dTDny6xIjuDSzamktVXFs+uPxj/93T049+
+dW03D3EbTR5Zs7TlskEr1uiCZG1TjtlR8ZrMu0trUnSpVQaQURWWddo7iSOn/2c
UUJRTIKx7MS8R1pnH7aDZOMg06siocZbaPSsYx6JF+Ii09BSi26/v/GytuxjMrXZ
s4lMHLRQ62WIcuzlosa7iSf1Dl/fCevRUGIvytLY/Syn58Pw7UZdShVqOP1+86Wi
CaLUO/2usIlNkgAug3q7XYqROZsM8Xi8puCLOJJoAvpxOBxNkqtLEerIoC2scsg9
dT8dC22UFCHIAGcaq2btTQwOLx/jzSzlRljtBnicTRtzxT8VKuqcJR76TZfFOX2m
vKOPaoPtrL+anp6G0Fm1Qj1YW6DddTzyLFWtxJ8++gxwAiwELr4CGjJzH9hKoX2H
u2iZS3apRoA8juhvf1ZTZCxh37UxaP9+jdahHGdbbZqucOy2F3c+58SdZnEpFtsa
uNFphwgkpj/VYLIk8P6VjZt/UYuTm2B8tnCZskcP1drZ4EV64AeU+y11oKSYDfeK
6Ms2u8+5swLSnnkn5kShrWKzllZWLRxBOkUgrPXFdNDwsG6tjRELojis7bp3JzMq
eXfxkErD5UYMT2A2GdOZLelHgV4+X236GlpmHYT3wqUD88eVEWJ6NYdnbVg0b851
fZsqpc/1YwaqZSSQb4Bzunux9vww0+KLE7WdLobLLye3HIN4cA46h92HDyPzlXQs
Uofv90SutTgocHd8o9UFdd3sNQnOpSnq8j3U6x6W7A17YkfaVrAEuFHBB5c88Grg
0pfhL9GSVpDScu/Ox4hwCrkvOYlwJhpsAN2V19jKCRKskNe5ivulV5SvQ676TRYY
PjZv5ODITU0g+GNYqDlybobgnoISBRpGVeFDgQJH4rD1EkH+RcZqU7SM0sgKmAqV
lqipB5XBp4x7MWohRbQqQlw2irxW3sgYIqZFy4v9RJhHpklg9dYfOUutkXBlzcCp
rWhIuqpodLCYeUk2Q1HiXHTILI3SzmjjHP9D7UvorzBu1sgyKxV1XQTLcL7Tyem9
zGpZ2HffOZZNwp352/tHVtHujNbfF8ndreeuRR6T2VnaM5NdTLNFTexOidXJWmKC
54uRpiw/OoPjEoXfaB/YKVKOpdt1mg746xWFcsFi51p/I+2zLVJdLeuL4jh0HkdZ
MhPgAnUN1T9ElBDizKbM01xzn+giuiBRdmo2mFBzN3duG78EwIotcU/rfMIJlK30
9gd1MxCDDhpDZfi21NDhiI1rgg7X57qCkTMZ0SmGnTKyrEpmuoJRgsiDj71B2pxX
iWZGbIPs5cOnnQ5jxHfvjWRuy7u9Ovs2R+VRtnzahLDQ9sE4d7GFHBBwRfMwQwVv
lcFmnfMCNvtCoSqKOc9p5gSgwumuBZ0mNIyiK54HguCF5ngg6CzX5TjDPzDz6afE
W/yw8nDyjexjH5RvuGdGmppULb0PCsKaAt24o4ri4E5K0pXkzugj07IWHWV5lKJ+
akYu0jZrh192+KEjKz0Ez90RJs8BkyqB9Wvpwa7YMQVN7JPoTybUV2Ueq4BNyR8A
PPjkuSOVD+db3daQu8yfaC3jraO7JQnx5Nt4uZm2Hf3q4PIcOXV8qipavDnGCzUn
xrOb+MfNpD+nGSo4ZgnfYJ+RnVFXOFTKSVW5wiM+7eVDE5owYMb4e13Ke1E0llCH
ZrlszP1wZ9vwFdL39txPH5nXsDMyH2rBLs+uYsJa6lS/HQX5P+q+ZFPdh5xcL2K7
XYoJjHk5PbK8WjfLHIuLT/3V7K5dEv2FQpdeeN/a035YcrqlXe43kifjURmFCvIp
ovR+lg7DBTz5SDdECAp+NT34/EEYLpR5x6ZSo3EVY4gLULf3L5uD7Ytoc4HJaKNf
qnROWl4bbS/JT+h53Ki92+bTPTz5txK925bmziehqHQ0txVYM3qzDpRD+Y1R36lx
o0stQkrCioTa5N5ipJ3az+wKoCcO0uTiaCRYsV0ykIn3uPtbkNd+tGr90d0dwA87
1mnMeqsCUUa/0vdm6S2P7fs3ExAix5jpItPsJHZNREVT86ych9YqJQs3Z7fhreX9
fzuH/kDDlRmae49SwM+TAOkslXRcQZ7Dwtq+astVss9KtcdzndcMPjsPDUZnUo3J
DQYC113v8RgpY7j57po9ZGhrsijVCSgr2fmgWzPhPDPEm+yV4Szx1pCy689vI0Sd
5dJTCEFqlKo7htrcAUGzaIKh/a5LTshg0QmE7RhamP6nbhmT0CUTAfdWwIcdsREC
YHz+DgRWvH8gRh9PzrvlovDD23afe5aqVAiL9k7nbQRGqORLd81317pQm66Z50k/
OpDAm31or4P7niAX4mVpbrh6VvujsDtObB2aALacrQuKCIHUt8mO+fEyi/Hemsr0
HV5gBb/URg1TnU5Vojrqob0AQ48nJ/ruig6KTyGUtj2cNYaQAoRpO8Jy+WUH4rsx
0+Vt6JM+SLHNiVPGeE6StmmXJAahEdWUh5lCyrD++/CkEzvO/VJXWz2wyFzFnfPr
K3x7EHC4Y67RAR1EEf/POXZXOGdgJOXCOcvg7AGUWeI1+wx7Hv302TvRhM3O6Lx6
JRRyGdaAT0pCuWswPwaJcOl3hwhvNYqv77trMrfGez4quUgt36ZhvmX+dLhVVcp1
9JBE3Y9NParV8StxaXZftXOgmQUlldCK0Y/Ef3VZ1+PI9UJwkkf07XWVOlKmRKFZ
j9qeMMbOs+9QoIu4b0j6PrPAAHM2ZTN9knYwI/NJKdWtmqkAOPdJmlTZZvlHo7QX
BFZZgP9WB5HClAU3+zVLTTn9/ePTg57eys4DASOQRSUa/Ojft1pHN+jK5LSL4pcI
gxQlDQ3wpN/hrYMDXIR5EDX1Zz3lEq937nIdloIOTwOd5OvFkg7/d7lEM0mjtJr+
MvwKKsXr8gdl7pLHXWnbrclfz9t5pcWGZoU28JaJf+RUA7gTEkOUvlP8eZtIfBmw
t83NQpVI0LfkQjNuxMYAmJaBBZvEg0kKSXgklps6mo31Kxi6Q1hkgb6iSgcr2i4I
XDsE/uzqVfKeE01Yp9hg15qeXIK67NoK7IW++CRGTo0fxKRvN/dhIkL/cA6vyAVE
EHaNrcCDMSndt1OGiYEfvuVBpLlVyGXA3SFDXf5PRfLQ4Scw8E1aZMPU1l0t/Y3q
RxaNhBt4tRPwFN0pkmFHze9eAg/yDV9pQQb5/6iF0+U6PKdTmn1Xl1ypUPB0Wva7
Po6bwjiwqjGb8/rIwdnXBUk2MiEP118djd2wkcqlPe+ScNIKg5xWDv39L+yxJj9q
irzF/YOdmqTqxUpuvDyeDEd3PRjpqdgdEd0B8G2AmAVfx/UY2og2LWACzRoX3di0
b9XjaIkZDMiEkEGL4HPGpGxXaHlYBQMWr27ZsVFnv+SkpaDwSNJIZZNxauYlHl7F
cALzK+KvAob229moINvXu0/IVTCODaf9f711/veqGWuG8B1hlRpesr/szWTUfZwE
WrM5knBdj3hyjSiCXKzq4isRdfBD0RxC9Znx96fbzKlyQ0ywn+f1TPOq0NEO5Of8
tgAuYtKO0N9Ze5kRc1p7lbvb2o7PMEqt1egtgrVbQFFT08r50T1n4LS84zQUHbhR
0rcbA8tk+GcCZJYOLK5Fhu7Ye4K0c3Dyg9CuYSulCsPlx6RNzW2+7Xr+WWaPy6ZH
fhh0whh4Hnifm1Eybs2D9ZAgp+r9k+FI2hfIBpMF9vEiOrAhzygdPs2w43IN5mEV
wONMH+9erV16BYRWUCkkT7bzvTJEahKAEnZytWnWBNg+3DJw3m69YNPwXfpp5+As
E0ap8Qo4KQ6COLmpKtCT36eaxrsivXiUmC75IKMsAAlTiBwHqSi/gplGyI/YMIfC
IWYPfWySv6jQicKFQO/k+uP5gwdEvMmpioyxcvVVv+CjPFgInuUmTRbgX9VyOLXc
mlzvb2fsnCURMb+bPkZi9Cgyj9Yft2uS3zY03jfuOZxpFmYrRQB9iT/cXhifdaCm
iIWFILpGkaRwVpMiALXXSXz6DNj4dNG4P322/NrHtEuoO0ec4Mc89TnF0Ex2/JxU
2V7shbGaiyhEg3iqPYQ9bnp+EArc4cyxP6yARab9sGg5j35rSBRS53rYkwnh++99
814lM/T1/xwy54DbmY2Vb8U4OSmWQwRzIgGugwOXILcZ+Ff+gh7KG08IhkAAGW+f
s3qSNn/NfXeA8Bw0/kn7Hl2hzHGSHi5/9wCFf3STT1FJE60FbBfPyF7egbbg4/Tg
tN9DNKJFAyiKwFNoOqUodzq7g4g8dTkiFjdz1nAC+wqRptLnbKzG0CgIgVNvCTXj
kco37jIXUKb6qWuFacyn5pKTI3MPb/cHttXx+DT163znOPln/TFH7Yp9TdTQytPz
h/BlhxKqBI//AAsPJEz432cVOydYcZjb55MjcCo3JOejD8TnGLecY/K25oW9YQrH
m7BWrK5mM3D+rNHQrr/VW4+zl7mmvXxL0hssIg8oPKwV3BdBUvfUI30SpRq2lkNt
P9s30qytISneUY8wF/Sfa4sxB1N9K9alA4F8SUcFARqk++7QacWVw+uG1oalXUqH
q2LowrQ85jOpy/8E/m/9NqGy5lbUbX95DTzitwvgucB7cqyAEHnjvSmp29qSIWjy
t0jHcqMvBQObyA589h0rwNvBqLduym6hJke5TBjL4JFB4PAGz9CBar6lO41CAgN2
ZiJj1NoWsVv8ulGaUulsS89oYphbDlJrHWed9yd0A2h/61fz1MpnQ0SjdvzrHqAE
YWWsijfdjl5GwBNngC6oFc6b05OSLiN/Bj9ShsHfOOS/twk2Rh4zLas+8upJyr/F
nxWo1qw+xGCjuz+udfNJnXU1dOGdmr6wYptNAwDbgnoflBVGXlbicClY0Wid50tx
K0W7pQGc7HXYrgQ15r6/1cTHMnlyxeBFKXOop7riYVr2iVKR+IBcc93M5kNaXkOr
mlGaFK9banXbHFo0aDDRrzJfLT2tlKbst6ip/QxkV8nloeLhbtHAy+LcJwNNfcvL
29gRBvLzf8wHUpOJhOnkzyIhOCky6t0c0itIlscCiudpTdHhCrbXVjlScEjLyn7O
oH2nq9WeY438dsTvSPjY0ZkNGXhGuWf52g3WjnuO4T68MBFnaPsDYClo2SDh/Y9M
lav8FOozih6sXRE+RSLFd6gELawY+9TiVdP86G+RNNc/N47n2uDhHCR4oZnjKbe3
aoBN6z2CxI453wKG91ZfO8I314ekjpo6GZ7mgTRExsPCGMLtJzYQ7iTuWK5CMptD
7TUZs3YUu3BG8JCn8XnY///TMplkawlxxgRQ2uZV4q0Y/BUmjNwRkVoDeEZwyK0k
AzdFwKgV6mlPqpg7lFYJPywQjhn6PgmGW8GGmh95vVrjXTR/Wb6KiDD//xSJPzuk
mqCVz/H/i9ufYKgS+CPTLjJ0+W48jXxyHommbzHZFaiD1DvgcuZXJwaBL2uL/N7l
OViMx3P/oDXfWH5HJbrbCbHXhLQBUQi7PoTo2PDdK3RLbdCOkTNO1a7HwK7cBNNg
25+OX2G/wy83KE0wG2IfWuJUXRIlciF4+6iDoN8r8BI2y+ENPE0cesng9BE9KTa1
M1h+DG5JObqk0sRCG/hGfXLGHuz9YtGwVErs0bYCXh3aS07yBHMcZyZ+T9OpDYPr
Bml+xArr0vGzmyr1/6pZm5SOZRYTcFuvSZf96yY1ziAZqIyXpezDnXbamfzlgKnf
ZAvFs5nqvneBrQeqMjYhRzptwu3TF3IrKEn1gpwf82GqdiZY4sEBvi4pS3gzhJWQ
j30cmQYCbsqrTPMGujOXOzhdnoTFZdAzu/MXJURMmQ12ykE6P9/v/2tWTrLUcLtc
eG2x0wisryH1PKRlisWilGmszuimL2tk25yvkkCrEpDxqbsAA9pqydlhDis4QoN2
ewFhuMPJEkI1nAlGvv44qFTVmPLsu7JtLO735qYjIcjaAwtLQwsEt/RlERjKfhXt
jo0dAfDTqIVqZgpk37x4uAPX+SWKdCS5fIw+7zEsulQuaY+LTYBWeMs4X76cplWE
j0l2ntaZgOtATNtR+iiLwKP5+/uRE5DqsDj2XsXbXHrgCqQCbWZpYKTvHyOJncq7
/6BIx5QaU4tXpIKAg9mt70Yj0jUDiJW2ebu+UCyaezZoJOsjmulEhTAADinrFuVh
AZYftLjZwcXqTrTf9yLpgtQemAMHF/5YYI2/dfV1RSqn8+HniVPxpPLL3IWG1bJ2
IAB2egeMLun6/OKLCbiuqsAQCc+SLKYu6rTPtLKSJQulRaB1vArKcvmHVeM0LsMt
txRirWhnj4W3tyV+M/B8VeqWicQuWyc0yjO8/PLHnUXcIL0L3pliGTfh9N2GxAvR
8rvOhCHAZCYOrIUS5tleFgYAujYZLdLjq2gznOKelLYLruouHojQdQyBEG72LXhj
jiFAYsxLfvqLPOIDuAUhJyhpNvAYhBWYdAcsUhU8phPsWy67WWunoMslIV+PnK/m
lIuwowLyQUf9gNoVUUEY8DcddGjqwQmgAV1oKtr+rR7ZGdtVeZK1B2pH6fhKL0B4
etIOKmlwJ09hhGa5O8LOIQSbb75PcK5xOWubQ8iZTdbIdfvJkRPA3g3cXlmos+zG
jLjWs7aGku6IGvAQUvA8/BJfk8lwz9iOBVKd+OuviM4z6ofW14yZIFZBibFCrk+E
6px0ZyuQ13c6RyOfoTqYPeSu9JckTFTBZedLXK43yUmyU3687vBOQ5AOs7FOOtRL
hjLwDuGqhjCZaz1i9DrAxahI7Iw1UdiijCdWPVf0YjV8azDG0+XfZsh8FFdRQ5ot
Unh3uaB850GaryrrVzvE6QXGKhI79LHuPqfl2QBA0E0VkFSMi28UN2zAYQp0R7Au
KT3yltaQ311C6FeiLv+eowp38ZEEJj50OVrz4NsGDnQnM0GEZm8NxZpIHghrF8Sw
j2I8XttnhzVVz54I+cFvVbA+aLQcH5u0GAOJWzngv51WT83a/05ltncs8Bme6bDR
EsQbWjtmi36iNX8DUz5dDRZwJXaOBZ0rRkY2y95wygtBma3xV+N/XfnO50o1bkNU
3fehhUbVmO6hdbm7krILL/iPw4ajFqqjT2aAxTPLNDurxryXlvqbnld2XR9qi3ng
xiXUOD6cMDVxQGQc36RkUxZAEUEVZMzFF4Cp4JAibW+GXmXOiLPFWXGTXEixiHVN
KVi0mBqwMn+s/TtBDTNJ+adU3scuq7S/8HpWLNDlFoNV9eFZnnhIfnmJKp4uNIdK
9QH5Sc1jcvdx6D6MUF6AYNsZJNrzq7RZRNkXRbP3EyDNwRVB0T2bP8sf1aLKG09y
m1DB/DZ4UTVVpAeM9ZptXnOVjZ4hNF8ff4F7AZbsgQADdGiaRzADOBS/qJNkmODy
TZwtxknBH6yuFJZFpjEn2Er/gnC9oAT0UD6u8IvBGd4bCh5ojM7jW4s4U/LJX6Ys
uRgZ8gRNHXC1Q75FnGNsR1/fu9+vfUt0roKJkQfrIpGUVZaoGcj/gcSkvlZUGQjh
QgekbNMIeqRByThItOKv99h/oRg46zcznAptBHWHe8zXi5GLizA2HmTWpw5pV1Dt
jCJNHlr1MGo1lXr0ZtepU+vEtt42ynAMxuqB5RmbKX0foE+jb25AX6IjOx57ZPHu
EaA+iz9N8veI6j87Wn5HMEuTIGD3P3SSGyWSluERkQbdgtlvl/tfk1pRPR5PIcKd
fyXd1ByqsJOTmO3NUMzfK0B9fPQF5tv/oNw20JMcT1reJqrrjVtyYviV7uc9Kivr
tPNxNB0Af3KveEEEtQh0OjoPJi4fjI2BS/2kbEolm9ZF9fCX/TXkeWokB4KhFaaV
YCoMG2PR7zAB8mKkhRGBR9SrEEoZ1V25ekb0cjfx6d+ZovkZnwEZQff9LmCaRGDT
2eue+8TdPRcYlQFTqJZgLlnGL+2+/ue8oUkTH6F+itir0pgi176XCoPc3H21raSU
ojAmOXFyBnpHYFgTlG+JDDg+z0b0Fpe+deReaFl4lsqmt9ZbXRkeserSGVKg93Ej
tjJH5B4MpgL1/ZrWuf/16e2+xOoWo/jkNZsRmZ/yuS99gANmx9550l6GTZpMMxe7
TEnSVfr2zpYG9MDetaNrFtzRlV1wdlkcHmd8QSRmblfeeOt+oUbXjds4U2xew9Fp
jIeKWAdVZDK6sjaQ+6EF3Z6yGSlIsa26RDzTh+052B1oh63jxmrzpOcmhDut5p+o
P8Vhp2dR2gJ3D+BuyWgRdEA6/NGcxgp4f3ER/hATJSM0+J637+7Xvpep0WM99jgE
6WJ8SYPB98og2UusVs9yMEBgfOPcYkAERFsWmRWYgA3IPy/qSu3fvqOc5gaL9rNH
eQuYyJ8EMUHzJ6rDQ6fwH61tfI+L0Z7OmQj6+uAFsC0GV01jHareoCiWH1cfFoXb
9Spt6h5IsP/lb/8COvbD3wiYAH7sMQT0RpyS+pr+ZaPbEUHqdfZEgyoNYvA/SlkQ
60AjlNiNVaBNIUBChcWupP3JWd3obTq9mptMcAM5QjimTlwDiqlJUv3GKrtA/ljv
sjK+0iC+/OJWXRWp3qwv5rTylxXlY7mKe3Y0SsI1jn7RN1lpmtcZoJdc40s00BQO
0c/Veg+Bm7aY1d04mQGQI4jXV0tCTLgOcLUD4OfpxL0e6Rr9hNetoitBv8zeUBIf
gKDCOf2v1N7UGicgs/6ufRFQul+jjS1T1a9od+8s+cOgJvPaTcwiUBPkgkLozspb
MMsPJuY4Pzbm0+r+Hgx4FdrsHHidw/PIbKVaQrUfQ9MLcEqI458sTRE0GozJZExa
yKEzXwVACCyyUU71ZZ/fOsv0OLo9bDJPCw4JToCV2lRM+o+4keUocjqdsHKb9XE4
zrv/Ua/FDEjvrq8Jk+XUdyOMV+VrBPLtAke1Na2zTQBEmrSY2oqEDNJ3WHDZ4EF1
zyf6mmoEIGQZF7OXv2MPuKxc4gwdnoiQLwsr8rq6XRMtYdlynh5ZxoMbmy0Vki0T
jhuWNGOOazS5Q3J21FZ4K1c8yPpB6JiglI6lzb9ziqb8741WPpBW1fDqO+oTDUYJ
FW1XBBehR74XhmsfQINViS6bl2CNwVOW5VWYm9TaGhtx9+bMgpCWufuejnnwFd7T
qcV75XDonYYbl+XCn51LDe2AN/6LfvlXa15aBA9ZOnLX+i8ahDCbowVUWV4hfcpl
7672vJBC8F7uBNbIWYCSm2N5OBpCMh4vx5OGvgZJEcEekQcHoIOOrA0LhN3vuSus
lVvmugv3CFRywxgCLE5R5bwnnqas7kS23SoHe9lwXxZV+0VQ17ah7FkMdsJyO3+N
MsyXT8j/tUgWKVzWa7y77Fn5MNnXukjez34uRHVOX15RJaZ+MAjbTiNgUybiWkHJ
3uE4/ogP33FpvwEh23ocb1o+5xB+iYl743Bd5xO3EhfRdfUx3CwOEmZjZHiHl0ia
0AD6cqKsabfPwSCvTwodm0eqPhH/fgddREW8nWR+8s/npT+vPayChbgHVIuKbI3Y
YuL51U5L57uVdbMk5q0ibIqRHFcd/TV5KeM///aYwob05OEsd1lqbwgkzivNzjyb
+/fYBqR+99l6WxJfCWF47k4Iur8JJvEhDb7JbmwosGvdPBAWk598S1H0ZYft58Bw
DZV4+rVfQ1L+3Byfjib16syhJU2cVdM+IvPfxiKGKm5xxyQAVK9b04U0bOhqgmot
KqbCtfBiVcnhwbdgMac6hXmbYCPw6aAj7/6enlOXFQpUBkQ6k5QJ/iICN+FAbuhI
vArY7vuqYIWRKxkbAg0l4t4fOGF8wdP7pSFHpBmCI+C2S9HZqMsbUuWvyRnSf3he
ExbCzrVuzp68hY7qpOF/aAzEdpiTCCxM9TXiXZfmg6p8Q6QaUSaqaqKHPmzL3S0F
qelz3cTzp/rjz/8rPasXQNDkvPXqCgHg0mrzSO1KLoTZhNpC3HSd9XrEnOvywkbr
DovasqJLBlY4CZmAS/lOV0M7A49Zem79MzIfyNxIcjs/MbGMxx+JgLJ1kMLu6Zsn
Yqa9szpLzrtJ/kIdopxtQ0ndQmwk7DPzWSKV9DVcXAbZapA9EBdRB8oL7wtgJ7Ts
VXVubjzANvljGDNPxsYJudYrmcMCLNaxShP8FcCWSmRi6M8kEU8PSDJGvkfYWOqm
gnFhnIq6+uqOzZrQ8yb++fjOSEJYVXR/IwmhCPAIEREoNCmb/iQ1xblJK/ybszf1
8HmvqCQdTR0vtvMXGco1CE+d0CCCzY+qynky7qzZl8hNrWWp1cqi20i9S+b+PT60
j3+j+eQj16h0fr/kPdc/GX1FNppTOCib1dDMATLOwRd5cPwsWdL8Iewri2KODayV
UrfB24HYuD8yWN4iO4IOazK29Z4kbNr4U0/0ZLuis9TnAo6MqU/KLNCeLreQbCf5
ltBwb1zO3mLTIz/aXs7WR3lgIC0cpBdaWTzDfKoiw6VtKfGcR0cEkwWFGpDbAYva
N4UZvrp1TStilCRns9+wfDzye7nEyl6v2Xb/+IPr3T+8yPOs3tx/olr63wB9Oj+Z
V+/YCbxm17tWyQtsjpl6SJ0AfyB0oSf7xPxWpI1oJ1xQQrViJadb6fuky0gYGiqh
XxHehCVNb9hGgUMnG7wTfjXYP1jphcHt9FTdoT0q7ytUTTI0v6MPY+VdjA3PDuhe
ZRDJswZElNHsfRDNP8BLyvZn2i14+nIUbGDyIvxsMCA7gJ3iKk6tD3L6XIlo0ArZ
L3w0RFKJTapItxqwKZHaC1/rj5OQO6z2nPmJBfrGJVk0jJ0BkyyMNaK7Omj58TTC
nEP9vCIyq0g2HC3TlsGnR/mZdgbYxXh8ZaA8XTYbMZTj6gAHxqS87EZ7arLV5wV5
/PcUCsMb/a4kWrjsLcp5QS5SQEubaapkV3atRLhpCJdU/ryC9eXUU3T/agOgYzMp
IVMFIIaDOrprD5u3qP5ezKBcd5nFvBp/zQ2m3EwmEnLLKZRm4GeR3Q6ig5Ua7pDB
tlSyT2Q2Bvxd8RrlQV3Cl6ROTORCdUJZwkLS007MEKE/B5O1MEaRzQM6YUr4pS8e
S72EEx3DnWl2Mv6cgrBOK6bHvVt9yu5wHwvPvwc9fJd0XMDB7F1mTqPJk2kH1UMg
mTvuOERa7ze6azIEz97y/7P+EwZajVGMSqCbGVvLBPsXRDkf5nA1zmWWxp77jtOx
BczPWVGSnw4GG/G2qtxfqX/31gxLhUJbM3W/IW0vUKquBnFKsINwdjPiN1P1fEpj
nNbjRMmhCWvy54sBpmMDGX2OgcBAtRDVXjZjudujGNbN3mPmlZI4DUu8/AAsp/Tg
IgvUdXeEv25deNQdRIx7iOJA4DSjb059NE43aonEQOEF4bxrs9pFSQTi/gX3plLG
Oc7tBvb/42v7iRkGjjGtQqD1VCvd5XPXR3GdMBKLylsib4WM+xhi47dRjv1anT9N
U1W+rC2GTHoyVK6tA8IeDgj5I1MT5Z3oDUIoSaTYPVz6TjYCruy62yBgrWwS1T4N
e0ZOBwOGcbTy2FzqqNswFxQiQ0XUFVF7xnpweWWFKtog24DI0NJ/4w5dKhEVptQd
X4nJdE4mBe2O9OS5JPfbPyCoVnIKaXXwS9ktcVxDeu7XC/lgx+zzVmllj8xiSPsn
bH+4hz4ifUwMWw0xA6rjFWSRiGbgxhyZWPlnlvJ8p1ibzNVspAb6z+Kmf1BzFdV7
iTVikfypcg5O+JZWhecnjFkuAPbxuK0lu82tvtGYTxRS4EgeTlGIvw27wCj+bH+k
F2p7rh8UFNli+gaKU/0ZKmJHn7BmoAJzKa5rY2ClXUuTuXJQJzfu82DWl13Uk2pl
eNmnp0t4cZem3jPfRn0Xty1Y+MvPn3Q9/KCv6FVRhQXm3RSznfWt9mrBpLQgioly
RVwiDCrR4IR5r+aNvEuPilcm11lA83K7GGCmzbwAgMYbWfkP12BeS1Ff2ZafGnDn
tPDnyuNnfLUHxr94V4Mc4lIcZoVDaTIapK8VtEBTh+VxSPsIdtqroBlnreCFwpJ6
8xFl+VXOMWjWj2a3FUHk3ABGwyW2VPcknWimagt/jO7GRmElQhjOAuevjTsUUN4z
EO00PmHCvxPCIzVN86a9ng1SRTA4Vuf28gSDS1Ozcg3pxnuG2DYLgNkGIKvrU03+
fXdvFoA94ZWjt2uU0OIZqpELzQ4OuEmyex4g6jMw1NFXUU0GCdX+7UxTbqBZ5cmP
fI06jEPviT95Qemf/Bn1X+CDioi2bhc7Y2GqxJ9xYT6exWvA24WFxmcPpxY5hdFu
uSEmrjaRv0ZZ/AYCGbKCHRus/Ue98xFS5/YJR9nLI2qUAI8eslYvPLVnGN7zf5OI
idHU1oouV4RvdDGwhPABE36rO+oGariZax5nvDxEnlAr0HubRweoPU5HZ+dMsWRp
h4Oma9QATAfl95fX2WawRMuEv8KTYsbXPdlRLnTdtvFJbruqwQISQvLCanG6elfH
fYybcoNNduOdHq8bHi9fGILD93mJgmPlhlFfeSfV+9MLsZK1ia1z/HEycsIwTB1i
nO7tMnsNAYtR6syffk4llQ0ioPcrMjP9OAsXi72wOFk4L7AvmXY4JRTaQDOxNOrX
Ez3j4kJzdpVwovwP88YVAgcXH1OxqmKhn69E+HEZb6IMMc/Eilg/5Ocibhr6xay3
aW3tJ2qrT/eVYTFKB6L7Wjwqabslc5d8D67BhodnAotTYFOrMSqBM3UadMhPUBVw
2ZQrbL5fyUNBoqLC6h+HFWWdt0ldOlnZiR/1KZBFmesvT5xnPCwxjH8L8KWV5ZN0
IuatGA/yx8IIweKm7gzuqVTKwkrLJaBYXyDTWPjzr16dUc6+zUNemptJsm1t9ILM
5yvjK+ID/zu2bmOL7R/PklzDPaASS8qaHV80U58kgm9ZKw9J/jDPiFUSXdHMWrF2
GvnT8brsNYClVx/KjXYAYXUNd0fhNZJZUixTqvsnbvV98rq67hq99s+/J47MAI7e
MnCQjyua5tYV6brkxFr2IQ3JWq3AjZlWxqXD8eJlGZe1Wr6B1msDC0yunjmg/RyD
iGwXwD7LjDAmCtYTWIWN6s3zRmalmaE/S62Sp8kxhwx8M+XNx4LQe4njENrD0QC4
Ithsuh9btSHPGXpSeziH8TpyCPA54PVvo+B/MR19mnUaAcPMIRWjYBk75+QumgAB
bWwJ6iRKyr/Q1h9IL1NAXcjtaE9RuGiM9DWcrXkyRi3I1cB9Rd++FmPDx1v/g1ep
ibpgxqUOk2no2JSkZwjw4wmQ0RaPbaLMiUoOVL9AABHOHGsfAit1KeXv/3YkiNq6
DE3mb8HwTNcy9M/W0PthMRbOY7J3WJLc320srCthdiy29320upkHZem0kKRAiN4v
X1piCwfGflmzBW02u5H6U5XkCoAVFor/JniaQ+Fyt8ro8zdjsDmSD/qnWPswOVOe
Af44ZGfcbk7TKxgAPQuE5xyaXKTTk2C/d8EJtrAKnT2CU657ARdvhrUbprJU65Wr
BecQWGO4YEI6/fQCEWH38XfDqDyEVP3kV9LDKPNSQ4V6D/hb+kENIsicehY7zVP5
RZukUWJxN55+SUfGc4FpJEMPAN0Pdacpq6gaqHmDvBViqUXBX/a2t0dlDjJc/xku
1p7yFso/KMpwr1wCNnarOZfcFyzdDEmKZTANI9JokRd8t5DifoLfxc5oS4EjJpXv
7hHkMVQTBJwgb24H7PhlBmf56FbRFEDw4ag5cd3mi0h1xnNn/v8Sgel45bcsHI08
GhN4LC+i+5gbnJyl4snWwiF9LotrdA2ZQclFuZoC5Q7HQviySF371cP3fB2pg/15
clR9VhUYOWymloWpYx0sZOh8EvK4YnIBXjjwEGewXhj/uo0jOOaPkyItOvnKr+mz
smPkwZV8hqPQk5j+YwPE1CcuBinVhVsp9t7fsSPc5rDZbIMNlwcfnKtSpIhsHTsm
DegnRl8vz5DOdAXwGPg9+TkKkuJNqYSl0FG8Lg5q0c8ragOVzz2mYOo0GgFC0DEH
bsls8IlYHDuRuynZH2S9IO6qzltzVo9xXWKYen7G3J0qV1Mq+1m6sei1h4u7oNVI
C47VPxzgLajhsc9D3sRTV1XcXB58MpNtY8lEJZ/BM1wHIVWCLI2iOI++0AT6YPNY
HvkB4N/tSyAK7jrcpfkH8gWdjDkAdzHGE8i7KTOkw5v86wGolG/9TVhAriRg9wkc
5A8G5C2WT0dl/N2xMpeimZ/vzgkFTKaMKPDLCqeDtX/VvYNTI/EL+x8h8LbTgO06
GOrbfQNSnFelQn0msVn8bfROU1Cwaotn4hygSbT6TfIhl6+GlqlUH24Kq5HANI8Z
7XbZ7qXa/Oju3RuwPk+lnVgdqoMMG0AwgkPAZV2QWab7qC7htH/ftVIrpEr0cGV2
yp6M8F8rOF2x+74guNcY249biFJ/23D4YZ3G5l3nuRh/cJ6U7isDtFtWUO6Y68tU
EefOn2bh1V+CvRIOPEIel+AMJCK05xU54ilqkCOonv9pqxMAYYaaXLbA5bjUJfgN
ET5OVeZpfoTH2Zc15I1h0FTks7VLzcCnVY9cL+thaEEpNFFFlE9DgJVhtH079vue
DTj14NvZnltspQhyb/+nIeviRl5JbNyKY/jAKZgZMzorwymeVO0JzsMK3LF6tDzk
GxpNakNtPlC9PB5yVPDq0UNT17xTSPYf2FUV+hIfYaD+OdcelyK+lsno5ej7bQCf
ZRR6W3DD+Y4eUoW7CDJWOJVT8rYT6161IkEfrvI3itWP5wsGlqhgSTyeoGHtZ5nN
YN6lWCdiMuNBLM0OwFG2QLl6jtEmfr00Xt6u9NoFi/r5FVogRRmjpK+GqGmlSKxK
uOf2bpkfkw9/t0nVZUvdl6TgpCUgO6z+ZDsN+COZE9yQzj4AHs9Oil34auBLTDBS
WkxUUobDzRelQZGgiQti8CM9CDOISpd9Id7S09wuxjCTbZ6G72s1mWnM03OwOEEz
G9U2ySKbXBsUmu7ek3334M85iZWrLkf+4g+y9iNeNaf3wPPqLeXfVQJaF09QTe6v
JI3VOt3tVwK6SnP+KJ/QHygSkLx8OF40nR0lI8XUf1lpcaIK6aGXDqBjfwPdmLP8
QBS0OqufTHRHUWYMnj5qMe5fWOrX4FBTNxgP7Xiup5WWCR0jUfg9VIwcnr1jxXyo
ydqIiA+zp83RCf3FndTuhL/sxKEX316AS2dtxkYlL3nTa4apVQ8dlc14nedHfCjc
dhhN5gYKoyqcUhCOOCMplm8XUJmtsHtED92JuQLvuN7kpXCr0bt4gjMLP+1IesO5
SLUPfoa1USHZCckZC/yzRLB4cqj8BAhpglcOsrC41kAD+a6xq8d26sADXHPXTulJ
V5ZDeTFrqJ9+CC/gSwjXFxu1X8k7rq0pksqW5R+bvmcEQ+FwomqXYbTCR040TDKv
5AlaUWh43s23L//zSsW/081C3mi7Gm/b+HwdkVRZtLXZ8m4CPHJ1KKCeWm8mo19J
kXc7k57jxWnratXjkeB41H+VQUP43U0aTQaYp8yBAxJ++cjK/+eCikd77foq/c0d
XNgrrmjcJGPCaG5kC+eURHOUP4USh/VGfULVmYBBOpsmNdYjE+cIjZWtNVOuixcN
GWgXylZ7VU0a1eDV4lrQwEbCNJYeUmBBooc1BgM+jGZ0wur18lyn60c/AoajYG67
V4l+Mhlt+41cKwS+3t2yJUUiAbV5QxtdVBSpscALy7TezqV6lAXowgiFM6rZiSy2
gO5HbbqnHwXCbDhdH0K8ekQPLUBI6hj3qBBYimydzYYkG+JAXRXmHru4BWoaRq4f
TPovFPBHJML9PxcZBcKI/fVJ3JP3ua/906/FgheWjnqxL/lRzATo+jJQCO2RoOmj
lFYdH1aHWAIUQp9ioxqj8r2DbuBDi5MJYGtC/RcjADIuHGJ5mkZrt4+sAfwclgIs
QfCyMnWl3/UDB6dukb00syiw8rpEvWnmbXxnPcJopeDstc8COro/H+MZ20UahqbW
VkGpAfTItKvF+qEC8bQQScZNKF2hUhe4ISbPhqmJqY0YNYEQFrzfM+YY7KBi+j0J
2rQUjbhw1H3Oac9f2Yy5LeyQLtXIjX62z7fKLK74WnPmohVduQwlEw1AX6eSQiVw
ujuPOgrEJze4NngcLYit3VDjJEeYpuPp3pkuZEPCNWRS9E3Rffug2BrUWyH2+sqe
0VjcZbf02qbNV8EUkld/DaDtQGwuU0iQx0tWIIC+LOQ0ZPEMxZc8utXbzXrh/z0h
BNWIE/q0K+DwT+KWfRbEcUc4I0fm9nLH+/kcHIj7uuCtwVVV+ub/vguuK1g78Heh
Xl45ruMq0N7kH/31x+zHstxbqiog2j9zZpS2W9hZa1sqzmKVuzmCvp741Kj81OQ1
LAgT+k/ynWixb2MZtdNVeovVxC/Q5AvCyYacXz+4Z0P+Hei5/zOy0fP31c9aNEJ6
2ij179E8hD2/ZciLl1hRZzvQ/hd7GGT665JoFtXXLTSsV2CDO8ou6fztzMS6a4EK
AzNIvWK92htaGiCkYKWOGlMdXVvml9uNNQNYd3ZW0R4S0yIFE2Q+PeK8ovDXdrX6
0aH4+EEnESJm6GfmR15BT7mcUJsDtSSKAPc0y21Tb889XzbYQiVo3h1jqx7UXOm2
BpMPVoVBlZf5GLlopkU+PbF93Nu3Gcr5pPfaypIpmMJ1EgZQ+L1uZyWgZ9FBIx9i
RbFDiR6ToiOSdQHKMlwbUFuY8n+T1MMoltFpmljZtWvOMErHyW3twwPxzCrwPP7+
7VrtcR16//5VO7YTohgcyncsM1hST/8Xz0fDefN7MPIZCl2hkypRM6eI0MFaIj9x
ixllAUMFZlv3L4jD3T6ZgjifYZCQNrV0u7/eutd3YR8+Fokc8kUFMkTh0VdTdiYK
cJsXyT8XkVprYSdTsDrY2gmw54oLF+FUSNd7GuEvm+n7O+Zs3s5OqoY3uLB1rKGp
dP0H+nciv/s9GDRSp83HE+NgneYcWfUb4uV2ydx0k0HSsBYLZ5bPJRVHT8HzEgrc
/b00DIEWfTulCaYQno9GjpQBMAPh8qwolGmESrsuqG52jBOqzsCgI/C+Irv+eEx2
pC9WYRGSZ5A4TD6/JxdUAmhJzHvncVS66bsBAL4Z+MJsRlx3EUCz7FOOtXGDwVlP
1mtpwrSQeNnyYyJgHIMeVFencJ6fAoujxzqN4PduseFdl+fzTmaWHHQy9jMUQIGk
V4e1PoV+uGsLespj9lCPeH5u14YotusMP5gVM7b0vTYOj8LVl9DJ3zEfXzPhmoQM
iDsP2gqoXM3PH3QV8bC6eJQf7gNTeIjRj1LLoII8vZy8ggZucE/gLFxLaPtVq1Sv
QzD6rfR0TMBGFpUeqwY0uGogilTeP8vTUfnU+nCMJZKYsRT8lx9immhyZ7W2SoUa
buVWXarK19K3eseQKw/FTbE8XEaZq6ldzxjWsm4MxcgxIYGET5FBVecGuTNeEwOy
Z9P8Acg6wR4vtfHywsXRMNBaHzwksuodltihQcnEzGH38YMi6tpIxCK0nHZSNNtc
DTKDAKt6UjTQYrify18b4fHMwelZZR0iKnWRvOdMC+pVYvrhybOPxOluZ575/91t
Xhhc3ikaOZ6IGC58F9V3NsJA59GW/qyLDAhmfp3jLkN0kWyepvY0NHDLmqYOlZh9
Wk06d5rD0cEnUSux7LA6cmWTMDzPGrkV1skcnne1E/5QVlgvS+3mwmQWn6fhCEds
+VsRKcvSvMEgJZkkCG2ii6sseGh2J8YmBP8yL0+nw6cpaOsKPJbUBo4bNIo4+7Jh
lC7qZWcBm6Eljfx0D76gWG5hZGAvB2cCkhBk6semjH5sdZRPpC2zqyapag3GHZUN
bdzfedgUMwdCSiCaA89D5xtYLv8WlMQqdqdopphkkUO25PdlFCKDS477sFmGbqRw
KLQf4tqrCulzODv3sNyMMBxWRtr13HDmYLqGw94O//bkwZLxUfLOHbwS2WJSNxfW
m4+16J+V9SROMgBaDxmAez6J2G/D1la0biEexSPyzG1sn4qHB4H9wkfaU+N3wWSN
7UagHHk2Zp03OrcsKq6gCfnOzls1HHVal/YKq6CXDNtya0NzK11nKfvUoORioLHY
eZptxNmQwxdUcif7mtTo9PG/eKsjS/gsturPV4ncCldbf/K/egZdr74htKqhxJ4r
bLLVfyvmRJEwn1mKsqQY1Lqfa8sJ5oet4l9aNcJtIGn6fLekupXxm/z29fIlDh+5
b7Uff2wuJ464OkVHBIsTnED2lFqXabtHsyA7cGvR+eh2pr4pVatqeLAWgJVWW3l6
EMEMaFyGYM5KL0mWxx6fu1Q8PrHVBV0OrYq8g7qXSv7aA5v1I5b+bD40tlvbxuP1
7GW18dGuZiYKkrjVXVCo7Ff6ZlzxcjgQUKbVe6rbXM6IXULiX0rX6KJxwH+yr6qp
yMrAv/aETsJk3FWWseBsPQRi8X6EpslDUEcfHTxYYHD7v2TN3/AINmZRyZxvPKxw
DqtmM1VEXe1hvzrm7fbJQ5bTMkZL/V0JTKEk8reVWL6jV/HouJBUkiIPwbGe/7Ro
VIq+kevT6EwHcDTGgKP62wGELmWwS9DflfhXizht5RjYHXuvqbtUzLghDb+pNRM4
gzUOChE09aEIS/S5XG4QWx7JDrpuRnMF6zWfHaHetUnlvbKSzc0rX9Wq7HM9j76v
lDB0L0SjVjMn8ngEmJiz6bx4hjnZoorID2MTW4AXtKqOemCygK2tCUnTniOjLgd3
Nn+fBWGmfdClzWetiXPozh9n0mGe/9NB0CtTWXAQDHXkVtkWTyhUdM+mM1q8qdhe
EmSHUOZUu+aQpT3mfsGaweelA/IQzBEReTdihZPZ5isFX96Wom60HmRL+4E1OWme
pakUaHlgmFQhxdr7VXcPa42JkbURvc5l77whiwa+FKIHjloTYNvEHJbbAXSqpZ+j
kwXHMEbfrk4GwdSeUQFUodcojM/BeD2xtsSb2ft90OtTu8u9onNJKnrRSfJEvg+h
ueJmE4StOrx2vMS5RtkIPmSmQDVg05Zlk4VpoEWCwz7mmV1r7JHi9FcxgAhv/0zW
tdU1EpLwPTTToUmxpWyfu/BUCJQbZknZblfPiq9kl/o6Lo1eFaqthZF6VP9ZqWXh
zhKwvE8p2syTd+UYopR7S9yRCWI8xtVePBcOZqMyVIMTEAGVk8VE5AvRTtjKfAJ8
DCTBUTRMzJHQTIpiupRvjG2ytJzkXRyqtuYhbbd26DyUStlJUW0NX4IO/fNMIZzP
Kqhfcd50DpnhBq4XOZ1ssMrTzrfJqJLVgqNTZl2zLHIFxEIFOpR4bnSVg3IDT74H
TmuwNqlyGTIcFeKlTsb9HnBF/2omnmOE3QbJqODO+uGC2IYcQk99LuYKgZ/0ZyIx
93Dcrde6jhZt9N67i2fXO7nueFl15HhNGmP1JqygaUT6YKp7id6rRumeNu39RQwE
rMNLx+unvAg06L5t6hHfkIcpPX9QAnfCJWF6K/ruM1Voxe+ThIYtv0xWnDrVc4P+
yva3QcEdR82uhrAT/iW4TCc2cTKMsPWRSKtjnqVcvtMo+Vry85/2kGX7vo4Ti7rY
ixgMFzTciWQhagylop+ye/vS3+1buTOS/T7HKe9lid7FCkXB57tHsRgAzaWodYaf
l7w9sDs6hJa1i/QgxSMDKAUFLRQHy18sR5USvheNBkGQcgXAUo/xwO0tMB4b+KlQ
LmjVT4XYciOXb4VewM1QWxZG7TZIQBjXJHMcIWUAMFIhOubR8uKCm1+q3gJIE4N6
hPlhSHTirHrI/4gzZ62qt0IBqlVpwJ3BNX3AhfVjFghFaulXvJCsyKqMSALRlW3j
llHhHy4Z4Jo2NYlEznedjD4lIht6t73ptLA8ZjL6mYLRd8OYwDpcCmZikrEKH8es
hhcsWJHLfg+zNLGqE/Zf3YaFcARDeT8jcwON8A07Fw8lMcDtsyB1RQvas48E4jmp
YpzzOhikwluM+67hJVeBG6pZ4Csu2T86EiLN+1DNd8FeMq6AdR2wKyTCT+aA7CJW
V4mVh2T9TOM1LbhsiXOnn78G1zj/B5fPIJAoP7TuB6RF3jzR3adnCF5hawRhlPSs
GdKKulM3iiOa0GbH6rkczuPJVZykCss0nWzseJhx43RhThCb6UfRp1/tic2NAvz/
nSIzeTcS0RP0GGvK3OXocUpVePDeIcFZ3uosToWf/2OaJs5/eriC7temla/stJE4
mdR+y4+0nHmenVZLb1GnvwRS///FvJJ2p9pR7Xn/waaWgN951r31OpBu6njYhcp0
D6qar89NzQijOjf+AFwkGVhAfOW4xRXd4bBzy9WxKfGdN5mdkQiOG96Feca9b7BK
S6zyhEo/mMHVZXhlS3/GDM4WMzi6t6nRYZAvKsnnc/cwh1CqkdDaDSq44b/mvph2
UYdJ+BO7lAPefFQ2UxKcX9rUKvj+ZHjN0VyHOZzsGw9QhituvdQGO4/J1uhva5ms
/XZYyrKuxgBUJNe1+ifNrJ9bwH0BwL/dZqYLQWUV+fi9VJNrf3o6vYG0OIwhG0Bp
0rz9jx9p8U5LjQKyV5z0pSuRx45UHxT6jjJ5ejcq3o2Vs7LIbFX2UGQQeAsjPJKF
5UuqQq5u2ygXCTDkXZ6LLyI4HLPz4FhthvZHwRORsL4YrAjT4A3nbCpTnLMVRanI
pLVSndARGfcT2XLVmMUGG0adE6GXpNN8Dq+Jie80a1Knvu2l6jtS0iUkK0bJWo7W
hhGTR3VSegwhGUsbsjD/JhfjMUIyZfFaCAVcnMJSyyHv49DRYdc3ge1kzRhMx6mf
dx9lB1RJT6+WaKI1D8ub2V1uHt89dhUDj1tSjrl1uZHNNWUHjQKsFJ6HGzEWs5sD
kyMNNciucGTRqFY9I8mLSPkNiyzqNUCmRJJ2IqEPUk5WbPBX/yWiBHnXLji04EsK
m5VjNor05jr5I5Afs4p9JQCAlll7gz/Pfu1+bQ/ZVufSqP+OZ3bf1eG+ONVycucR
jHB4issTjSfguVZb5Tio8ZRqThcsefcivw0NCZFFsUFMXSv0cvUY1rE187kD0JKK
4eCitwfPNJlXFX+4HpC486Z/IFpXQM/PRAkkDn010SZ5BBBD63jyArREGyxG/rkp
a5aa9KiJla6XYL+qHY9VZd25OHRr5hivn2g4HMZXOQeDyDpK84EZtetdF5ga2kc0
IddlL/k3HO4pYieXMUaT3Njb2R3wZDzYAIkyeP79X+atjhKh04ljlR3h9GNoarba
wGz4oelHPcQVwHo1qn2TYh9/AMFWn7pEvt06tSdzxs0X0kqvkFCbcGsbAPPoyM9f
pfTP014aswjb1wQLb4J/v+ysA7ZUMYas1Zb1o2W+hXmJUhc99TvbXn9ZAzENAi9i
FvNZY3bY9K9dUUc4vQDFilyAqyv3vWbHNla3IC0C5sEUq0gDM/pXoNWWI/UhTCJv
d0eA1uSFMpI1GVcIBmB7GiE5hDEIVu0881o3oDpylj5qxUUeAv/KrZSRVyUAmWg+
d/B4ZYem3QLEekFhRur69IzADCu8Mxwom5BvDf5vuM8dYzBTC8PrxrMj4YuZCn5Z
71Xu82pW+zu/rmlWMygY2A07dPsJmoNRI2c3hfXdKGa3BqrzkVYCaClzuYLL6F4h
1q4RCVBgCf4eOPWlBmemjOHIj02VtOaMGYGqKNE8PuGZ6A2eKufa8MRkbnFlowEP
CzCvZ5JCleiT6rYClynMllifgGmkr9eisUgyZNsPOXDUh4gahl6C0k/teezKZ6m6
bDRYc3Aj1g+auyIwEdTHTIoKPCFW8hZaszPPqwDIQeJo4myh2RkwGf5Z3mcGf4mg
DMPnUincMvkFQuZDo99sEzldTosYxfLUBgZZ/PoP9bni0BheWNJVk2B5ZQOeLmzo
TNLr1KIK6a2X0Pmq5KWin3hGLd7CI4ATLXxwXb2keZt1E4Jw+XbobjC11LHA6WM0
vK1NNCaj6fUkZHEtJGIYhNoOyHa2JgM1NIbfe9ItXfHN0ei/BSyLRYAinB+nPeNn
rSsCjgMb5opWJOtXLw1Hit3V78any9TKBdkfyAXkM0oRqLC+KVY/2oEH0FJuJc64
cvenGfqV05rstudNnOAkbO3dJHXOH7kQpmSUdaMPoPrpBp/z7y8g7gHO7CI6h9sw
/6ZMOsjC0bK+532YrLCZrKjfg3MXW3VIUngIRERaRFZ82HIrsgF47dCf7Nu8HLej
hVqo24Yt/N5vUxRjjvzyL2dnN9iOg1EWoRP+wmCxOVF5c27qQzJzzdf2IKKZWUbJ
kjNoIuGYDlyG8e/u/la6DzQ2Zdh3Zf0i7RogEHbEUhhBBOCwuFKWg4pGA9PYHiZf
tHCRoqaV1/IrqkzvDar5FuB/wxbk4nsy7h1MbJ35kcXS6SMpbFSTzMokaKf/N456
hPUTjc5ol7KdN+PRd1mxD991vpOStlnluRIBLGJXALrFEFWm0KgbGrGlPXu4hmD7
Eh7KRHtOIUeGtJMex+Or3g1ZNIKqMHqZowsqsGC2DmuHgjPSiCXiwzXTfyITLeVI
rXBLHKgTYZXZajhYmv2Etkw3mvU7yNsKcNW6yUnAgVbl3WoW3uC03eYGPxs0EFJg
BJbI2FzBHse1D9XApdmPPIIkx1KcARHuvwElA7tYOyG57MrWBPi6VRMeZYPvMcIO
fBWI0MV8UL5bhrKlbM9RPBeAY5x+X3SBm6Qe+N9q2Hf+U3iIu7ve+YROZnTKkf1U
qqD6GUG6nEI0c3qlhxTYif8hExY0xc0wmslk+pXAuOQxDg5jccX3Tgx2S8rPpIb4
zRbGoCrx/Q8bXveyG86pSx3TnoIi5scMLc3sUo16flbeNTovoQbUWCgtHVjq7w7f
LHa3/c1umafNbwnLHtxH0AoqAL9EaGxKC8uL23WZsFFSUB/ubhnFKTnRJPdpE3wN
hclwMrH/sivkbEYDcMS3HBPC7OFN+VHpkqN85V6HIhNFkCkq98Z0md37ZPaB7Sfe
jZu5k8XgQ9Z9KTL/OpkQmukpwm6ny6xlXed5jX2o/wcNbsxUjVQ5apI7PbMfnWPj
InGIE+/dYGN0QjEB4HlEerYf4cNhAqkRAyjqRjNx501SuEwRkoMmWIES1a/qhPH5
AqN9wmuXeT6Vf0fLFQTzYGes/MewMfOYjzr5jnFxqJTL4CftB7UomzNxMyNDoL2z
6LinHAyEljh6g5MARrOWEy7DAihVAtJyFxGIPolx7/S3+LO+gvCoN2jlcrJy3fHW
KtS6GN6dBNeRUxFmsXq7niEz3H9kp/sbxtFXiQXpctGpP9oYYgd45V6YTyInZPQJ
nf2cNJqm1OVhfOxKLHEhLv1sFhZFdN/ihprQ2x6cUTP70guX+jY2yX9E4FdarrTH
16XZF97CTuMpzEUnnMous+WfiOZF39zesmRY4JhCbOqvFLFxyH4XzI9HkEOw6OYH
VUg/93yUskkb4AE8hmI6k8GAFMFHr7dTD0Rdz7/SClf3pUAsxtGxrNXLv7W0bYm7
fO/gPJWpGdgISIAJLS4U3HYYtatQUS3sN36jcXJoNL0+6y6vQ1TYDGeryHRrkpf9
TKX8xptKd5sI5c/ws85jRkxLKjIWqjoqZ5bzIYkxYQygLLO8ogTJ6EYmCT1eCvE8
s6rG06OkxSwvMae+o5Hk3WOIzZNepV41PbAe0lD0YTMaKZIVnE4MUdBG6Lj5LtII
1iI5EoGvzDg5lBxdrSkab43Jl0DJJUkIha11YM2HHx37b97g/qVLGIUsMU3uYDNF
BwQQku7sx99moVTNNEki1BrY98ZmKg8ZFQXDXEDIpLOeh8oiPbRoSbMF8Cs1wSmB
C72+J08ajZzUPoNkzu+27UQ8rMSLgODkl1/bh4tMzbiJ1EVh8RwjjxznDoChyN5J
qkmtA60wqe2zT925fYAjd06ulIvj3MflxCaTGRXH9jLPhJwTM0KwcgNa5ChzyxJq
Iml3FhxgkBq2dk4kDT//1hBSAATiiSLtAHqDQQZWgiLqDyAR46lE3wSYET/16Bg9
es83PkVqNq2EO1jqGAB+I8L2KGNIRCnEqR2tGcsEuugRrD/3iVjrJMN2BRJUmo0d
LS4VhA+F7BO0GpN0WDworZ5oxeSiuCOjYje/J0PrWU+UjHTvXxbEy6tOH5pL6JAh
2nuH9MO/gpt6pVTCDmuCcqHB6a5Rfjcw3L14rhLCzJLZ46Bcgt+33x1rHu56gJWd
BHn+PRK3TShYwyNUtg6PFLcQRnOS8cRgVj3O26oExBG7CpflprgUO2CDsFc7k4ys
yBvJNItct2sOkbVWqwApg0oc7DlbuEbQDibmCMl07DKNZmqZo3nI8t+s6rKzjIJk
znkrkXsndhdBH8I56Ah2yKeKSSZtLDofLPy26F7GuTj/iMG0UcFxWFZTEulnfDbs
ySZ2yrtZfKbuRMGxQO7r0rgSISfSg3lgcCgVIldFiB7AgE2tkBCIYRj8QklA6XdL
msoyLsn5VBaq8v1FuRnyLZAqQ17YHUnF4WUtQAEZyM5XPMecG0VFbWXFJaqQCqA5
rsuHzSOYzOhVTKtyj5WqD9E3V73FODU9Uw5YMOBKwF11YKC9t0zLOC2E96K7H8bU
k+2fheoclngN0LJPSPvKzKNXHmpXT/WFn0izujPi57/VJj/C7FHYIGUzffHMEldT
MyAwCGBdMrdJy9Z6Sc9coVpITqHAuTpYVshua7Dml/Pm839Sxh8iQCQKegieF+SY
xM4oyMq+tiDYaynVGFri2QOVH4aYYg8e26cNBffE54XomLwWiELk/kk2CRbB9B43
MkX39MiWO8wRpc2Ui/t5i5soIviKaB0SzIcjewmAyrCKxPA8aI8snQbNPuNxR01j
MSm/BJZ29LZ6UTUtRCZsQasNwFbI0Dj+6Iq0yTRCwXDHDF97TSxLyQ2BkA73MeAe
9V5h7sJqzQJBSyb5NFTnrKucpk+4sI4/N+Me4OXcG67h8QoYDtqEflK8lZvYohr2
tYYV5LiFoPD3z5Quxjdxgwg4sFq8zj2vWnLxWP9mut/7HzC1/SHkMVv02ZeWHNe/
oo2immyuk//1YFnHSkK2e0p5UxJTUxiiOF0U6QMjD0mxJ0XZoyiSws9Aha5sfbIv
b+GlyksAs2DT9RCHDzwufbiC3SYUTkutGXYVzxpbsCqVFY95ljmUrWd+HIOiFUmu
aeorhlqwdZCkvUg9N3kt2l6ASw0VVLbwtvinMMbT2XfuhS4M9/+p1QrcN5l3I9kR
lUoG2ruRYHelvDG/V+R9FlJRE/aRDdKO0uSxxU16CKrXm5xh9vW1rGGgusbKbnrz
bYf5JqNICTQmjEVRiqLcz7f6duSDHzDLx3jJTpkmhYKHO0f5IqCS5XHG+kO/lGkf
3pcFnOl7IqO4iRz5YWKe/c+6p2UtGQymMWwMtdd+uJBmJcjTOPVz1xMDuR/9vhit
gl4kD2iStwhkoQk/fOvO++xNLTSvYioFAdJgc9ezHDguPDgZz/r5IhWD88QLlrlF
/TgLSaNCcJD1TSsseeHW7/YCiRzb8zuxI6zoPe2ekF8f9mf6Vp+1AuTCtdpaa/i9
I+Oo1IrWC5Rdz8Knrb3/zCg18mM/5H0ek1qnB/twGcq0vqwyy+meigtx/JlOG1xK
6WJgyHrHa3mLMGqdZokRgvE8wpub9+UYkSxNPJyYEgTav6219u7I8YeCmLqv+DLs
3Zg1lhrBMog6Km/gUXZp386q+0vvULE+5htdqlrjLyYl/DWimahnm8YoNYihf3fK
DiQOqJLwxI1XdhPzC1KXIQFntvtMrsKRi20VYin2K56nSsLX4JaNp+DWE/brIWVX
cM41d0Rk8F3Y52uFn2aw8/Vmovfc40D0srTRBfinyjSUDIQgCM6p6hpVEeiCG3Nq
5PJ7Na+rPB0LsnBEdpwl1dLZphocZI5a0A9jz1gW2n0ak18oSniupa6zqw1B03wq
j+i9pAKdaNrjWo9d6S7LyyU2fJ4zhSJgb8ANUMfU4Y4xgTTJpcHS6yhJmk26rih6
oEajbjfTDp/W1IAf7/YDZE6SCloYE32tJ+G7Z41XJxPpTcpuRdB0pVo+IY4d5Z4j
F2va4s79tMaSyfTIZnwGCeTeWRpKda8ciiB5Aa3Xnvny4107zhgN0vxvotMucGxk
IQkmwDx9LMhn9Fs8NtQSzthkbal00lQUBmI2qBXNFmqWnm0bOZw1p8noK+QDJnVm
HsRtps/wrETq0FBGO0PzS6wWGAT/DxqeulJvYG4q+jn1rMKJlc44IMUu8NoJgcl/
f7dbQFGCoBVtPfWUB9jPNQ2NqGfePClmpbR90tBzE9WY4DmvW9pBG38P5WS0XyBA
zCwljYrXS2dgxY2WkJpsERLFSnj7ov40eY1a03PdDPQufAsIHEBRYEI/oFUC9X8h
06vLl7QxFwWTH4RqP0VLbC8FL60N8K25r2c8n3R+o2vJ33CkBiymrOOrPYeOcsiN
CUkm5qjYu5eT1Fv6tBAZY3IrKzz8bbpWI23No8XVAHYEWhwyhLtlFgwJmFyDi7D3
VcL6UWEzqZv1oIbnGlK1dMYnTv8jgvEcxyDQGX75B906MOJFJb3L9MAJt2u+Ac58
tYC7k7DibeKItjmaGh9dHfdUAO/TNdConfezccQSzar5Ew5uNcwtgl0kxe22jxzX
KzSogUrGYxZr+dRnEkNuoLigcEg+RW02Dz6LlwbuSZ8P/mwalw9TsL0rHB1hYWWL
FWGcCOGiNAtVjXAb5Z0hOWQ9VVUJi3kMth8U4lJWb+gRnILLkZEMup8uzBvnFkoe
CTe2+N7MIPUqzuJMiBgRVxYw+gWb+9arrPIr75bbY6pxIZYIuxtATbYn3idDjc6F
s8KrpgGmDkhn0g2MhuxsuiuuHIBv2H0JyJniE8UASRkJv8JnxwtRA/lJR5aVKKfV
+5Y09C9OMMY9lbo5H0CV0hIfgAu621Rq5riXaC5rLDxGY50XcXd7FTR1RorCwjlt
cKjgo5Ztt/qdZTniVAjokOMrcl7wt0LRjmoRL4SkDOjc3ZXOdYJdwTRoI7UWVy1/
Pr/iGUEqoTYfX7MVRa/ueI2PG2NgEjGn1CsJIMACpbHOewJjNlhe++cvH8Pzeq3v
HBdfI+SAZuqh03lf4hd91V6eq6UsWbf9i901Buaq95xgjQrprgwupqgeoiXgHhEL
tIXUnsSsVmD0I9iqSANzciJvzZUGhn8v3LsJ3YHWQ831BAFNCDvsdHH4cUYAFO26
wx8NxpLmkj5g6huwKuG6p2ZoD6EdBI2lz5di2WKtvtupxmFEO/SNEqhfZ8XUJulu
4nI5KPDPJ4PI8m1VIS+4TxDfrAklkp+XFsrdxVYE4fC57ti3c7STLzFsByCDoH/G
6pZQCggeFWWTFu59iOlVUlPr+6JDj7Kamxq60VlhPAUY3LbwdU/raqxJJH82qvGf
OODeZ1iG4WIH4NaCz+4WiT1oWjGtTOzZ4MeMwV1YkZ5OgNffdY3TcGHm2STmVx7Q
G4G463dWNd7qVNM6yYueDHVINy7OazZkYRztPb1yg2w6gQGRUPs1PbF7jB/nc3Xp
v0qru0FtIoaLz8LMjm73fGv8NShQzWLtUNHLhbgZBJzZ7r2Wlgf/8BzcC8GI7Bie
omjiF1P16cI67r8QUHHdIt349n6C9Er4R3d1StK5P/vq/UW+BIwHAXYSKgXWMM+S
xZi3Bpy5dWikMB4/102a4GFXmBgPiOJKYr1AN87ZEukHXWvehwfKmNoBO0hHtvIS
4o9bLH1AyqqQXeLYbmXch/vgf2XAkbYj/UIVqm4I+fCvk0jXidy6L6M8dLMfH5fL
lKFs5ICxqQOBAfEeVfspwLr488tkhqW1plp/BmhO9n9yrN+yXy9qst0Ani746dsw
qmTdWqZzE33LEgrF19rgd6qi1+rn7fuNDRzapG3Ajfix9/bWYB8pdRBSXW/ydytR
7s2dXjAZB8ifdIcZZkHvDufKgXCJMFLa1DC8H/xHvK9pLz+mYZEcI1rzti6QmFjD
an+HTiCQ80BKawxSgf+SwZqCxhL1hbojdfUyzMHE8imhWRIWEEg+gOs9Qn2oYv7s
TKnOp79o/mq+MaeINOlEVfHJJ3jf1fkY09Kwnc5DvUWJ6o6n8EV5Z5KntMikRdgp
LqO5Df9md8IIx5Vhwvd4B+oUcDPP+RH5wyfweQp4aGAvicRIoMrU3eQ6dpqCOkPH
c6zAJRyvePD8U82dyI6XoxyI6ldC3XNWZEWywd65yVT1/tBtMuFH4C6oat7mWqLA
gXubFrJGggrFqmfFs9VzjLNFTckOeLzzJDgTm9jqUQ6t27sGnFvf5ZEq0622nV0C
JQMBvKZXykTbrryfmnKTRjiO5vqQy2ntq8Jrw83tZJLDlUryi7SIJrzg6obuL3Qt
pViMj7X4klqt4An1lrx5xcRFH52KqXpPBig6IHHnNz2mpARBAwYq/OwILKsFPQ8c
VHYRSXqBzDxT3Ku0+R3+DA/UGIU5LsHlGDRrq+HImQOOpQeDdopcrTKClMULy+r3
7nP/2IlR3ViQv/Kurt5htPA0S58xslKFjycP3YzuQ6oEZOEJvsvgomSiOEr45Xhr
QCIgh+SHN7xyeqSAuGDcNTm+1BkfCGaqHlL5YwujRHLmp9NcAf2Rx3cFKzw/TRRR
MtjRe7v1Y8nYjk5pKL0IOwcJoUj27Vkm5zO8ClpaGNeX5G3qwmxrDUoC/zex8jJy
HAFH1XMP7QToQFXUwSmnLqubNwzrs9bje/eY0HO8k55qDPqC1XgX1vc1EUjlk3TP
VBXYxO55TJ/8qi5/zyBZYW9WGMjF8qYF6eVmCEbNWpSIesOolNcKK06hDDG9FlR6
K5S9StpjMKun31AKHhBqbchGg7QJv0SSANtsqKnjhsvrYFn2vV1T9hvZHg7vNyml
Zb8sPmYpjUZLCXIU6MFf8Z7wqKxjkUUnhbCM+i1d54FPuEHQ3fMhICdtNXcW1Qsa
hv/5A+KlyXR070i7lT9wxFDwJsRXQjyBXspKV9Nwn5LkUwTjY2K6sPKfh34AQiO4
o8D5dQUcDXlH7MFKPM1IDdQX6z6zVrFIVPkunuBkp/lXPzxa9ONasbOwX8kvGA3/
nQyzxVnygaLf7BwIWjsMmMoTPKWS4oj2CugQfL+PxxxJe28K7FMu10IvdSdFNHts
+LNWkcnlj2TOez40O7mxy5/ThiN/FgIHwDi+SglZjOkel2LFrwzifBixKDA/zdxC
BPWKDBi75bfXgAu08GQj4sMN9qIq5ycVLT6wyTdcSWR7ZT5eUJg6VtG2bLXWA86B
sVSJbim/WTxViLYegMyv9fS5qh6m9ezoOxTw7vnzixd/yEGKMEaS2SCp4wIS3TvJ
n8FUQQ6ADqhnlRdZbAM1NJY4Dw1s/ga9Ds3gH/SqkqBrGPC9umqWsdPAXL14EzbM
wr/vKZPY6fWPtqRh/5bdj7OofQrcitH/gUe+2bhNToatV/kYlRb2Cm1KPKpN2nnY
sv7TXBktfE1zplVnUec/dQxeejK+V9M4mUs6o1lI5gd2QomDnv/H3O0wZwVKyEgk
eKzneqQNKhFIf7cCStH8m3T04tflRDfMh9pGIHeVwvMc1Ps9yMXAWugyONSkf4vb
4xZDo5/x3J2HIR/5XeMyhaWMC76BPJ6RyP09s/NhVDaWLf3lGRnbV9de5j3fg3Rr
EIuWWziE0EDPij8CwEQs9uwScLIJJNNDhs8AnU5JM8/CaetWI4E2pkuI+kv8ewOS
l9M4ovhxsdFOKu+S3GRCMyLbysjlKIBkcwtV3iGKT/sYwPABu4NShK/p/avHBQCC
zilolkpmgsRzSN+/lnC5YlKowAF4/QXx9byGecac8Ycgbbyuu4OQl4R3y8TVYIaR
t4CyxRZRBylHxZA2y1Upju7wOMhpkFgbZX+aWR3Wb+XbFONZ9foqkF4guJAJiCV8
/ScHKE97WRmq695s/kAUAmAEeHIeQegxacQyZlaCSj/GxSX2SyoIdwUuchSWbESW
vkXiWlery+GcilDTx/S5/CidKxS06Cf4AUXgHB44lGD49DjSC8ugNR9P+ZW5+Cz+
VfDsr1MMp4kEy7X/FalhzpuEnShZBgrW8/DpVWOjq3p2g3gRSbd2+nnz5Jk1P2pW
AOl4XK51nximQ1h71NhdJyw9FD3kfFQYOA/cMFb3dYAvBT1zTO+/8LTDAWBtlwAZ
uIh7GGvtnC2eXASc81SCj1Fna7LZt1sDp5tH5MNbiLchaXghxWhNA6J9NDFoz3zB
0fegiYVmFrmRJ8cn7JEucA++jXrrz7cX/mJnN8J20BvVxZ4D+9ZEOOmYZ8cAzTfo
y24f03oa35CYS+84/Kh9uXZnmDU7djXoZMVmYTBewIvFNevyHCPAiZk5Tv7FUdUp
evNxHXZ8I92o63CuzHX3BRfbcsfZv5B0xMwjcYeENHo1p2VHWReKncAbXigdJhGg
miuMWbsa++h0qW8NtMcZsrjUshiUEbrAPFqYrL8A7ACdMTA/OW1PFXP1OegKg2Xv
Q9T3JlZmwWJ3W24/t8NULto8c5OqPM/w/7g+70ET3m3lsPgi0C8iyaf1ACp43XBu
9pzroF0s7atHxIfmF3XWlNQ3XcRSovHSi3tfVJ2zC/rvaY96uWsz82/1IUHW2Tiq
EN20C+8txJBC6q3kqpG3VhStE6QJ5avvITlu/UcPl+sDQK7xMML/WgkPcehbwAHs
Z3ckozSL7baK3L2LohtkfcOMuqjwgIV84BbYL5+nS5hvLuAgHKefIIVZNYzjCZEu
QDi4m28oNLoikpoOSFpWmQF6juffNC+4sTN3fv/9xAvHYWKlB4RN2cssd+8Ln1Ck
E3GnTGU5pFL0oNhCHzh8WsWoUBVGu99f3+r3WRJ4ewsVcqNAmWsZ5j6QRGX3UhcO
I+VeZ+b5Ia1TcSSkNrRWgza+jssNY3My+Nh9gtUPd8n636hc68zJVkKlQQirgiZn
U9UUcZuvlRaOpFlaXqrUAbxbpa0DF0tt5MW+NsRdYkj857upeTisecdq6iBGt61Y
g6Z0qI+/5W81R151Odmxsw+LdtHJE4TRdcCV+DTjuaeugLrQSlMBBbunFVItzt+m
8owr23Ys26AIzzAtxD1ZcLS0TRE2BuFb5nxAetE8ZUFeYhY3uZ+Q4ZIuY9AKg/vu
WrYhHmTYqfkPVfo3nRxvKOZ/V2WOU9H4NsgEJB5+JEhSBqsXxOhKILpifVIu1FVa
HK17FN8lWVvB5fLn7qdw1j3BBHLKJyKAbtBh1GI+zikqtvekwybKSCGOy7ZCgbKk
ASy217/G02fNf0JhvX50M7SCxq7/wQn6oBpIVdj0724109cy8n5Bt8RY8XSJ3Sdt
QSLDzbth7ybUl2jWy0tPfqEzwqeQole+4KFjigbmEIfururZMsIRF0Bb9PGsqzaR
YBRuM1oW0GaiuboPtAlgUi7XVRH7iZdJ8T13VKAGKTLNPsouCx5xhhhXfQCFgY+t
c0/891oaTOqfJK7P0FsPFkc/leLX1UVDARI3KJEHVb4d4tk6DepSFrjttfBSZYGB
DsDrE4sI92f1gm/xQeqX8iez0N2IFmKBZuArPi9AycLmAsGMMDWLMtj4gosvyrly
DYX12FOUOOO2HrsfjDjpvo9yMmrJMdzI4M2nIaHMqDbbFeR5hzp2nhzMlWp01cdr
trBUfZGyphMyhOWHZps2fVCXRHD09RVA+cgUvRc/8xD89Gx7S82aCVDEUD2A5coO
1SGChhqGYSLh5GcvxTRfgk/8o4iT6JaoDGlCikx8VvSNZMoL+Fwzr4j2wlH8xtf5
y36h3+PgENQKbj/nKPNhUJwpFVnXblcnYPNZQqZXD3YPURyvwmjNVdWrUsn6qsUW
U3zFrDaIYfbnM7v/m8X663CPgLgu1npH+v/l6ceqOqpaWP85Iyj9AvRJ5dJTknqF
5APQ7Si9GaxOEAPSAB+mkDjiS7ePJYtl9IcdX58epv2iFGuEhm/SVwP/E9Ah+miZ
S12MuQVdjoGBdD9JfAMCdJWvIC6ShZX76N5CHKimQihGbgbsibvjfXjxUUnlL9nd
tLQtS0ThUOmq5X9UCAINDCA/5kL/iXq5heVzyssvlJIOaIy6v5TsHys8fHWjbT2b
a2dHpyxCxh4AoBjAfp8sHS3wp8gTAAeOOPsum9IVq8nTc1UioGM6Q5XOgpVnJV/y
TDku1xXg0XHd7v0KcvVkjFgZhiQ1t+Fg+JEs4C7GoQeh95/OEnUHhfbi6EWsbN3X
qnks6VScvqlKLsB3ZTVsHU48PEpb9P4qsLGU9kP+Mk3SkLyEqDB4hKf788BXvyZa
yRBBJNI0QFJYoihKGYOZbmcUnFTfW9NyMwNPe49rKGR3U/m8IR2GSrE6xH3DgB6e
Db93EiMy2qXFs0kn5iFp33FNIOEgedkpHhqyV9/wxN/X30FiRYJ7+duJ0iVMWtPf
bsbHL/Qvcdr7BqGRKInSc93NWGdhOlYjfc3/IC3X4OdDr2pDLvzYPo5cxrBYg4PP
pZYUSGhSR4mOKczOI8qNPLJkk1Za/eEJpkEPvuE4qmSlEmcZKXf0VJ6cZBZ0RfM8
ZP0Ijaibpr47pnmvUQZrudH01KayZjCBhh0kfXPOOZqfN0ZkEjXEMRMhg2nD1NYM
WONkuH74IHSB3s+NRELabb6nu865rzeMD4kZ9W440kgzbyrZW6L05W3W92dAKavP
hmH6SSJjuisTDMLd4g8YSzJlt4vXuyv0XXGE9xGBfmB8SrX7PkyE+KgrEN7DC4DK
48TlWXF0pFbWbIMZcZm8cqW8Z68dg21jt+/ZtOOEXYFDjvneW9oIO76MdA0+zdq+
Cfei+Z7Jy5ioTd7f6/4B5Mvc+kMo3k5uq0wrMVIZf+78nKb+GGLFyGEwztoZqn69
eK2sEyLmdyjS8XECQy56CJwGaoS0WHLxvEgeUH8Y5R4p4ejFx/EYiZX8mjhkiQEV
av1napV87jVXfmRSDWxAH/2c4P18bOR+mR4R2oGrXAARML2km6jw7xzJJUKy+pSF
tAQ9QmE9B9B5HWpEjjXf6tbksKZjmyF+nrgxzMgom65YGBU1tXkk0XZvMS4wFIdK
307MxiOgySMZsbBB2+cRt2J2ydhSEG798oR9B12Fv/uCuCxOP1rB0gxVhMe/KPfG
lxG/TbRt2ssywYnqrtLKr6hAHTUeXYVIKawSL6XVvh+reD5FgMhhz0P/BTZeoT/M
rQHbytoN00Ah5XDpfrCSUkCnDfHx6AQo1vGSt5mYBHxOTHjfE83ooUAzwelu10As
Fy7nRBccOJqp90pYq5OOXj5HSoDrQ3vMn5ppaBOYImcXRmQUu1yhT+SuT6PsUIHQ
aRTvucasXxXiKVIbWf7hgt8sUrfxXDFKQm4jkE8JPXHhB/peinqbNC26qUtx/S8d
YFaWhNA1/jRVogfOKHMWssCnqsc+NjjyBBapjYlyOlvEZxMs5L0KWFblInkozKQ2
GJx81EMKFfOn4PzA0wa0aw0AREuLamOpLrF4ZZBcPm7e6/dqaZdI04UZ3vKTqD9T
RkldBgK038DPVSyrQr9erVvDjv+eNbzWWIbSfrC3VHBi2J/5PuU9ShHR0ns6SnP0
z3WXoCrn3pmNU8Q3PIO6JB0AGjs3YBN37a9lAFG/nvpUeeecKUfw1oViP1Qbfxpx
RVhM7UwLrk2kntJYvTekFni+mZf5xa4L18I7dlIBOSlPI0AH0hdjK99mJqRQxY5C
WSpECHfP12He+a9EA780uToZlLcMH4t6UOsOjFERpOYqM4T7UnQHya28BPraYFcx
wNKnZFoS+4P7D4BdIc9GTugwXzEYMLy1NT+0wMFeZJYeJodO9fufi0ByKhE1yWO6
0X8tnyvUVoYsnCEHw4ol2bAszuzEoTPG9sG3GIBqYIT2x3+w66ZPXFVktnbuaN5m
EzaiUomWqqHiqThPg1SfyPVZhWfocWS0KgQBiqybDYFeusrOG4x1NObsLcYJkLy4
YVo0sKiY8gsJZ/ytUmjVbyuLpGugbpX8ZhuM4GvD/hGaU1D4fzy3uOabiBkuhlOX
nUe5jvEyrku9aMkCM2o8ZFPNx9H8AXBE4QLgw3QGBOhImAlhWmOEUQLLloMRwDf9
+BBa8dvRgP3GApnGiS1EobKV6Nt97PlDieoB2g1o77KEtnZorcqIGLwq6pIliNoQ
g/cabO8/jjG0kp3RNz8O/cPwolnzz2nCnudoho5m4XdcpnX4zA4LtHhIljFDjxbd
zanvH32tO7T43aeCQSSbX101x8wLH5iq9/afivc1kcgonjoZUt/Hv1S4c9jFi6Iu
wuGAzADTkXXY8JTf+j2HDS9IBLOPX9LiItR6VWaieQcwhbg1IrjbwVevuE3G9yb1
H7Te+Y260L43cW1ltsp1Mk308APo5DDLzRm98h3VfTJ0pxVgIrpuz9iT/zodzBNK
hIhfyqR3eTpfO2GhpU27x3qvubZbrFq9yoAdRdQZb2Q4JzkPKeTN+ZaelYiALwwD
AxeuwIj36Fz4TCG7kK3eG+UfEQNOcJHflLMpqe/Gnxn3R+qlKG/xgEfKwNkIDXSO
QWmQCkdGxMjkRSrkD10lNhBMeq8bOzKnVd7ij8bbnp/o9oRFw4MP1t2190Pzh0hN
YyTovCzIhkdzxh6CIFwEvQaOXgwYwZtKpVjKDHdhb3t6kHHU7d+WJbqy/croRgy7
RL0UZKTUmsNIqYTMc9rmfBOIX9JQnpuG4Zou7B4oNCiVzdIfKSfScbenU9GfnGZq
4wVNb68O6h6NhSacLIYdEdK+aM4Hsasd/41F6zxjgAiQe1xs2qCvWe3ZrkatiwLr
gD4cwm0voZ1+cWNPOz+LNNAMSbb0566xIYWsto0dPYO3E39DTSNlM9HM8i7PZprM
akLh0yiMnd12XTyGRHgPtysWtxDTFXcAgMIOARMPqfFsHpRWAiQYP2Dc1zqrqQwQ
qpsVY7+kmBP0RWxOwziwgdkpwgIFHn9kkILJUSfO7ctjgkGRNzZsJIZCiUmhyXfY
AXU8poTlvw1bdoTgc4OHjRK+CSb41SxksHU7dpRt7D8jNafOiPhzS7AblwBvps6b
NBTn0V5a7TT5zGKbTZcXmlFXm3Dq3hvboerrjBKZvnVTwa+Sz71G+l98F7oms0p8
ReduAJ3d3fdZtyBcOxrxzskIhK83vfQ81lIxSiJPOPZkrVvlRGfLVhFqaKNM8hI6
oDgcx+j322rFHycdjHuFGXKQdcpvTCNRwKfO7Qj3W9c0eEvOmnJ/yCXCHrl35JLM
fO3GivgF0z9Kv+xnpEWzAdh5d5hUmlMjSGwACMq8NfQy2lzVkks5aqCXFFhBdj0U
zVWwsPdx+LBFFJy2fNsUnf14p58L1NNaeI4zuW1lnnfSn3DxvMAqe3nHstGHriKV
/osILqHYm+ieI3fagIV+8/RCxORo/c1yhq5XMdApqwdZdTqtIe3cXO+gyJls2vXP
naBpu850rTA7uu558UMgQqUaSeAkkfZXXgWpSOoEqfNYUhfm4cmW/nwiqXIdBA8g
7br2CHQIztAkDecR8I5QEynrbqKMFIEOsdN/50IZKn14lX3oFwHJMQhSIdwzyPNu
Yzo+9FrOMPVsSEMgFcafG7gIXjSO6JtZnFPoNESPIIZnCC4D+T0tOGMDxtjSJzuf
h9LV5WloSUiI7z0Jc8Tx1h+PKUMNceOgn6ed0QQUmj0pdtAKCqOK5okT7Tacv6k9
zE5c5nvdldcL6P4M60vtrIFhaBS3MBxoswOjbSBY0IQKGx088/lph/R04gCtKutV
dKQ6rJlB/mN/UTzCubFSRhj0aX+rBjon3r+RE6Uxm8jH/PeJXsDdTC3cYeVRVYy4
PSOtJiMczJBpUbYz4BPSzOedzGYwdYNgFyAYMLJDmLDKTDRrFOs5LLsJOfFosS/7
Uy2o0BXSWt4VgT0bqT1AiiUnTQ9zqpdDSkYL0JPJ8Qg2p23mrGM3447apusebx9y
NmeCoozDAxaF5VZpozdZ+srgKCML6kYLtHNIMkKz8hBGmDbdkxVn4/oQOg5A36Si
0qnF1O7ylQfsZvUzlta1Xzq6XeeKFHbsXzEADvgFjQMdHGFihv8fS0FjfzgdJOnj
M7UQ+8sxDAHMDhCXUiSirD7gXguhBTVQeEWYC0sCmZ3cfNXfgstgfDTAS/sMlIco
34BaIK/1ujvgmNNyJhgy4s4btASmqJkWXEJzx6lAz22qyjeBK3AvE+iXx7IQVpIt
9j2XWAUgEtoyi/ZnBg2WkOief6TI23OK4OwLHtMvWsiEGLx+rClyw1YAhKlj9a5t
wAfVgw/M/n5udd7VPbXkO5nJBFFOHciPMvLT8oaXtKsY3ro/YS2KClwOJTB1+Y5c
apZSpghk4JehkYC+AIjRgcz10QNSuFa5a98bf02/Q6VR5LIk8u1WjUoFA4SFIa3b
Hg/qDlYGWPguUjcUEm7l53fUp0B89lUbR7s+eeeel8N48FfB61EZ4Hv1zS67bZFy
nEqoOjUzoE8WIt/IG8DTZFcprag+1iY0fnHXQqNexvlLV4G9Wa9cxpgKGMDrGXrD
P286ULm4AQyxdjj3AWGt1PH8c1FdjraZCsyldU7JcIpj/uZhWE88sl7MX+vJ8vTM
WOXuLhOtov2uU+Tr3SAtjwDoB4FGyRBtBAvkkogvmqj5XQxKJicj+fxYZ2dLSiAU
q4fzqH22yRFjbVUlCbvLabv8lLuoyrlVJ/b3j9lJ+6v6KF7a02Zc+3ueaa8jM3MM
X+glMin5/Sti95R9bqQFepep3pXIXZyr7tmmHWJM0aq+eemjKqvAvas1UDRdYkD+
HKIjIhji091vc/8n1RB4eMZ22B9/Rs3TrlbhLQd7nYpiUsNMsUodSrFoZ3PjnE0y
9USg/f1EJ1mPQwUYUR71YlJi2pbg4klL2RI9DLB76BkqJY+3IZXSX8Xw100RBT3H
xHzuxEj0UuDjIjNTWPssWtYObHJ2c5KxjZG8LDCjcJBhmU7u3zu5eRTxwUB5OmYU
OoAfzd4VDDZtg2CECCb65AuYhvaS/cP1b1X2gyP8dRpsUYpCmNwdGj1BBjJdnE4g
R8me/9mUMEboB1+pxCsfqO09myPtqsTk3Ie6gNXZ70uedOE+3tLJnswWolDJeG6A
KzG9hazMbrlSfdlBkamELFbLKZ2PASG9IV+/53LqBeYy9XkLYx00IhF4qZjg3eRV
QEiYi87gOcaPRjBb3vvopnziSm/qfjKSWYszeIkU4ua3IcTUcXtWxQRF3RqjfJoo
jOFyr+w5YCqor+RLN9l2qwNQ3OuyK/ImeOKaEj+JCms551CNvHgjAPUcn2E9vd2i
Hs536Fx26KolmsaAOssGw76JZqX38Yuksn7+yUEojhVkKuK6eeOU/0H+2Ru074EP
OnPMPew1smocrta8FoT466P4KJG0TUosgVkFdIIIfdT09FWNaZ2STE+DzDMO8OZr
b8kjcaeUtLB8VcXEHo7nIjxzZebWN/uPd4pWLLn9HrDZTPamLgntaFoExvVcphV4
Y7JfosROs53GPUB/Ds6l37T9TzVWyjbgJkAM3xoOrHZMwbaSR6pvpoAZPgJV6Wr5
x4Dok9ihnivahCRLj9hEL4PhlcUXsFmmmzuLoRAat8D+ooILPe9Ios7QB3R4Bavz
ddDkyCcf5DU2Ltk1cLaJV60k8RTBoPOHRGRGCDHBixCaP+LssZjopyQ1DJes6bFX
OQUXBAkskmJn109/jQAzE3LmNugNTPAiK9DsetHnf/BoPJR6A7TSld38eEX3rxit
TeVW3owPbTygl0CPH3nhPhEYzNZNC2n9F90eaPDTSdieY1TQs9N7Zss8OpWG6QRi
I2/n8Kpx3gjiE7Wcta0r3B+CDIfmsMKgjbopjDNhQEl7he3C9RMwEjZekHpd7+nk
IEFnNQ/uN7Ut6MukHkRo7ErISP+aJYhyM+rSHs54SiUOCm0NLEdOf+GozsMOnsUp
sSUTpvkqLQdYP5hbvi8O2yWllydvFRHL6Lfox9apAg2IoxBaxxAeiOxws9EGMZwy
lT0yy24aminhuW9tpwSx4aJiodRRVVY8sl+jJndxskPUNgCjE9jsgnYjDYoGScaj
XKMM4snz67z3OtRgQ5F+hN4dNLVTdwWmSC3+HitB/O7wjLsWrkS3ovSg8tYJtYPv
dXy1lJj06IuzBqz6oAnSrKvYGb4bapQ7dKLawPIo3sI+sDXbrtvoBRxt+53GOYe1
jiBBeQqndt2Cq3vHDh5THxqCf3pTTjUuEYRt1jy69mwe0hevqsq1L4x3KQPDySWh
lm639Do2WoWZA1TOLCWkXZbE3p5SRSqC3yEFJUcDABc0UrJPmbnQQctWCON+ZzPe
U7ieGCG+JIsMwFBeB4s4R8UX7yJ/VMS4CZIGVmkOjKZnrcl74L/Zct5X9tib3876
/3+KyQfnz4WTGoE+3T97Y13qR5YFCjov+TaK7s3SSVW8XrXMC1vATKj0WjvQtO3F
ks2YDo5dFt0pk7TUNaq9w9PUMTcbGluK3VW9/BIhM9nB1Z1Nv8Hyth0Cw6i4wHGv
kCgTrnWiGZ3t0qwjUQiNJvkah5d/JbPTR3UWJnICZykBn0iwqjeQHIoLnC634uyS
aFizC97PVhV9xbDqRfbEN8eVq2k/dPceeyVZ/3+3WHXmef6CMO0iylX389joVhet
PX05DUIij4pRZGHEpl6CwWdeEYoT5a6ZXPcWafFseeF7n/XkR/AyWRewOG/LQpdd
UnyNuI5KAFv+l/CDzT7rNtf/OTGcCyZ38NPRq7yd6R4c8RQ0q1/JLYdH4JRMQGs1
EDZCEycILhBNK3PCba/JzbZ9+o98ylyA3205BBdo7kFjQBtczhRMNM7jpUcpeTMk
kIw0XU3iTK/f7S4ce6GRICA0BRk7r6GERz5k4jq9L49KqyJ7bVWKVnImaH91u2GD
mSFrkO73jnK1AlEPCCpxgyYhUKs0K5t50i8eQP9Fr4IlSUwy26pu1iD9+MZxfJIR
cTt17jOllUzrYsCzgvxWb5dnc3Qh3pvCliyKzpl030n9yXAdqfHIL5j3P8InseT+
I4Bmwp6XbVato4GDGU+zBKWE835290/Svqx0BsR2gGYCqTP/dx+t2S7gCQfSZUba
ByMtOQeqkKcCRw167SUAzLTawfrGCe9QHdMIQ9wP7VFQq/wRq5lPtnjV2pnuWAjL
CMU4j9ZXxyCjnhBxcY4Dn+P+ouEX8gKV6R/i34mdMneU6t+FNletJ3G3+xK7CCZv
Dp1/rC1wjTsDtrSAkMk/6V38+QGraZVSpmUb9YKhjNSYd0kXhcWkRP75QovKeUWj
MIHTz4OUoi+2Cx6qM4Cnfj2IetI4h81N5j92HvGHAoaFAUyA68r7O/OnQjrv68su
SksEhBMeXAKBo6iDvlyQU2a1K++RdKsMvzLLfVD/a5OGgUNPzvRBglW1lvZsOlB6
AUVuZV4IQD/dENTvN9A34F7+zPh3zmL9JIYKiU27FvAeVTTXD1QbLKxRp71kErB3
0Hw/7cY/lyRuUWNMHpm2zr/zralNTgSfLGgaJmxaCMKVFzWKHL2bBwyM/3EH2d1r
Yn/NFoDQlAGhxzIHI/iZfKw8toZ+3kT7olYi8gkHz3CtntLhItC3qIopqAS8ELJH
0ocl3U+Jik/ZkiWATd+BCHMoF/UVl+qA2lRCHGpY1C8NCS5opzipDHHhS08nEJSd
wpU0+7vzuYWNd7v5TsF5k7+bVTEr+ufVOXEVleSaM627EpHPdTjduu4Ho9y5vms1
AFnN+1u8JSjQLaSN4fez1i/lBHJPFNkJybT5CTO+RalTsWR8C92F1OntYTeEMDqe
iClIudxOqP94b2R2/cOvqPDqL4Dcw/euXMBUuofaoJBK6QdtMv33TYNLvW3vRth1
xrF8xEV5RdK5BZ+O9688H29H3NPqnjca+SlahPk1G9bWDCxVGA36ALarLcWDPPRp
C7mm44t4QNTxSYK+Y/lsaBexmUfvF+6cFLDZnVacqzs0FjaEo508zv5lFiT7BbyD
HCLMDggmmu92Z0YOZSiJrJ5kTF6qwvplfBhY7b8geb3TEUJxmGJVkCzAQRlrDEGY
KQA5qKR8+ZxFiwhe9mTrKQ6aXgNLJOzjpnWz7CTLGpX27b0VG0uhbcWpcAAt566P
eSwiBs/UggdGcUPMs8x/o447BqP4MpLhSuKuXLAJutidVbb7vrlnp74eJzteq8GT
8xVJ6Ubqh0dAXUOgBhtuAE5B6MHMFXPx6GBe+0THCbN+D/izND94q3uc0Wi127j9
OTecsFM4ei0Pq92+LneMxZh9TZ4AFpnncMTaHv2oday2cq7NGvfN1UrVOArbXwZ0
KkrRuLHxpCp4vTCJo3M3NbYOykxb8c+W47lQlEO8f3E+3e/ltq5eLqAK1NgkA/g1
nqKXzePrVmj2OCV64hhd6QjVuEkwjnXXpuw5xYJbn2iDHV5fk4fS/EAaQeLuRHov
ptVNmKthQkAHacZVELZWEziitUBWp6xeCu7WWWjUuKpksyAq01CfC28RZUn0qL5f
Nb21v6R1H6R6XQdzqi2jnaaTfFMdB/HBH979Jcay5eON17D4FJ0rKZ3JiZp22heT
+in4WvnW2im9U3yImvDKuAFT3Q3VcLMTM+OwJsRqHqisuluex09+Z443Rl3OITuw
WaddEBpKkU6y1HTK7Txr+ELqQtlSJrOGmjua70RPzVhlIZd/j0Zz0AuM4ET86Uyj
Xm/z7hb+uumuvCnzkRDf0CDTJFhXQt51VdoSkGxcbm8J6iGJXweTwcdkforslUjo
NXRVWsQpblhMWIrVVrm8jJnrVUGepJChCyuPkrx06P6G7x844EKcUVEEW/JGUEZB
o3TCIsiNvaMejZSJ/Q87vsHM/dUqc2vAmtLcBfhrNOsaEm8BOxIztYpGv5FxDVMq
6vMhTWS/pf6aaZu+RYCHiW2Ux+wgVobxB+Dv/t4Hf29OzUcQNvzWVJ58JpXGt9Dm
/ZGW25kizjjU/vFrsb4Qqkoq3M8wHXMThAICa9LYNWLxw7hv0640fQZUeby07v6p
Vd4z4Aq2b2UJybE9SiaObIKorEWCeeTWMV2mokPpXIznH7OwLO2t5XrN+cPU1evG
nuZv5KF6JtgH+Zb1RrWPIJsJGJbBwxemCRUdqGpclQTBGAD4yemnJ3HkMdZaoGFP
OIWt8znvuzPs5bKZpV7HK6HzTC3IY+60e038IDYSfiTrY6jwKA7OebMlxZ1VjCG8
gXSHHZ0ll/wItvL1b9Vfe7tGhL9/7W++fz3UQyRH4bt7AgsALwem8WMSIs1kGvkn
Aw7EX6dBXZlhLtzD8TG9BkiIaDGzUth5qpiaN2FYn5HbqS4lQ/qlZXbgADf38hbn
wIgkMOvX4yIsYrUeQBb6zowJ2w2JIQ7VmE11cbeCrWFLjSytP/IelX+k/XLWNss3
Ft7vgHPkT0t0Y+sVQGebI+3hD4DJ2nxZkxHDcAHRAKqo73IoJrtQt1NjVLZOrXG0
fYSaGi/ZrszcFAXHJ6uVyO0rggwOpv725IA/DEQZs3UkVmt5+7tnq+tzs2EwNS+i
XDJXZNapLg0joOyoecaMANqgIM3JwBMgvlonXdhmqtuRcfWiap1OOksUCpUQb8AJ
EB9R8R5T5b+T6WiStb4pwSSJIESj8dBqbHFjEaIigayIYDBUfzYf+QF11v4tk8i/
6THLfMn8UPJRty+u1sWyrCViG+eAvJJavAoNHKDOGfLsv3qBQ6XZVumr7gNVdxKp
JzdrGSJdYf/PbVwY59HKRYYtU72iOrCZIcOPzGPKnGSVN6ZB1b1aZDuS7jWuaGlw
xSvhVcFCA2dGcjyjeSpS3BLjSb5NUsz9lako7CYJcup1X2JVgZYnz3RMZr0tw8x5
rwjmO1kZnvPqwuB6bKzJgaEKJyYvKubcVHwWNsfyLYRkY804uWD088URQSlc9p9s
Nz2X9lxMm67/GvSXRwKo0CMDAl5kbJRqBbLMlDZSXSmMFUG+rSsk6NyXclloLT7F
0DyDUVVoECu2khryzTw/7fniU49ze5pLlNob/et115qlYDUR8Gz+rI4aljhk0XAj
jfSWn0xChU/hbSMZfGlqqkNhnWj+80RGZc1h5OIi0ynmyX5Zog8pHL6b5PvmY3kP
H3wiVLMI2HxQxM4/bj3ZPKQcdkSwKEtiTswUeOWeJdFX2WZpefRgeBfLfWu8hdMH
EFvaVjgRLBkEBydhHZpVdBCNU3jacbIEnEVjgEM63MUht+7QVnUHS65kavnDsoqa
4dESMyN0tX2kZkMsd7IumCCPZbrR6KuOf3SYlFpx+M4I00cYGNKkZDSyFzC702sO
rLVcJ4Y7qgPSlsHDJFrZu+6lgFsMt3LoXS0i29pbwvTQgUrA7QB2KzmFHmuckSJK
oprxbZni/F2oCIJGQ9/8nnQ9T28STPJqQI65HQuX+tmq0/JqLhOfrM9DhFpF66Dj
+rqo6W2zABqfz5ErYfH6GDh3aGJx+oxpQi3qo/tC9KK/QJZICwla7z8LMDbvVU6J
PbjizyG+OI6VnCx39AwBjZDQn39Tsbweg0Nk5FxwzG1nwi447mHx93TN54rci37N
fK1CeGgjP7XXxWItnrpNoQTH8geRIfIXxs+B5QQHIqZyvV8vqzIIw+xyVsH3lxiz
ni6B35j7fDMqBQ1zjabiAt2pL354DmKuZ/JxKnr0HC21TLItNQgVz8zgOAGjTDzJ
tkqgT0DMTpYiF5yBSKnimDWwbz+jLW/6wv4iEDmX2bppTgpLQ2CJ1sbbSHzzoKT3
Ww7W1RxNPfneo3AXuaNt1FK5rpQep202J+i+2YNJcH3YX35eOeWN1Ym2+hb5ZRtr
mXkZd5m0kq7qR/Wyx3DkhXKZS/YWHNw6W9uzQJWJD90jMpttcXA9foDCzPu3E17m
vaaVXQWOpi+b22SZjO/ljRzECrQnsPS2lkfUSMDjDei741Z3QuFq5EJCGFjMEx82
N3GHL0J/1riTx0qGttMPDrVdhdBKAbXsXvNbdoEpijvKR+WRQIi3xesURi0n64WO
Dn5VuIDn5KhyY9g2GGVxjle6K34dP7Dsln/iQw8kxkmYnWCNVTIpYQe1LaM1Ib3j
lVARZPsbXbBCD8FhDqz5EDcacwTZSVXP3laOr2Vr9eN7MLv0KlPNPQ6jt32DOkd3
Hr3TI9tIb+4U1K67FvVgix4Wiu29dhaimkdOhEiZOyuEjZyhWENe/6zadUDX3Jwm
oPBnbgWnDcx2U/1rp1grFwyvsZH4iqocKcSEmzegSgjVEHBtTp1LbiWqyJSC1G2u
5PoLRE3k2e1xwIaWTZaxbhSdw+NaOqZ0+zMzWWGQ21eKVJezD0rsO5HtQdZ552eG
/aEMOsnpsILuPkwsL0UmX9mj7BrVHOo8pgAaCEBnRW7q4U43jxsuaBu4Rn4gOT/t
GJrruZga6u7mZtPY/co/v2GODwuWD72g3E98M7pSk5Y1U+Rkp2yXhTmS+xgCNKxx
uBnqBbk/tMVUX6+soAaMGTZxwTmpmdLIiiR5Tr8H3ejgHjXlVljj5X9zTX2AJb64
+3uqYO7QYQ07NUdn4lal6qFLfvcf4gj/TvigIr0TfEiKuzUCQ9fa6Nb/gHlyUPQR
fJq9gEJE91yGWKjHjTPn34ls4awc9PiowbQLJrnYjDaXpI7QL6Qd3bgqMJtL+CLG
16sFzo2Vel24roDJsjqRT4m4VfJZvEm/flF+/QmAb6K89ZJxk6NPyXpaZP1x3OgN
tuS1WTZWqfHDI8p8hwXds3rMqmtyhcEB0/M4tfuzh9ADxNBwksrCSzPRNmmq8DCX
0bUsu/GYeOHggYdgpoKAINhzIn4hf5/kQya3dKHbOjdP+Sc37ZzP3oGQ6ZyiIFGB
z2UOOQI2NtqAEfKSTuI9a+Zrq9sS6lQF7LmGPjEK9JEfgguvNJwQ7f3OSIbY88RY
jGjFbUxBie4lacPxUVTmKqDCh1GOfv5c3475FN8d2UOxuld2DQC7ZI3ZK4reMhcJ
BO8Z9MywWQB4FQgKdMKaR1aDqcK+qUD6rbzUQASrdqBIM9BLk/ImIqYfkrfjkNak
dkRx7uJAf8MAjmhaIMm3IcYoILEWnGwUZLs2IEKAdzG4dmm4pTFyQStwrQxwXosT
iZAlp/sB6C+cPk/LnGJaxlceOVJ2IAIBmqslI2Vve52vhNwjewwFPb+bXw6I+MC9
PoAisglTaq2E+fpVltony2Lic/cS14aoWH9gfqdREumLVtQyyBf/V98fym68cj5m
uv5pzYVryzj4yT2gO7MX+b+6gTn+hC+BZcRNAXeLkdUf2MounkNZqVoXedO43Xjv
ObFEgIGdIfBJGy4leuEeEafvmL/ASana5xqhDAVBlTaEOH/C+frnl8+V+j3heTvS
o5PRBgzM0uQmBvlzJcLqQYSvUhz1yEuTSYWtUjEKn0uvEHbVIJOntEf3j8aShCby
VBoFGWjEeNMXygoDR+egGjvjIkyZIro0mJoAmGzP1Jn+m4frRV6rospXU1hd/6+i
WoAeROhmnmRLr20rMWQ3mSRHhJHMo3nbfRsWWUId5I8515FkViekimmksp3UoN+w
v386UsP6ZV6Drns95XNSVvZcBUqfLmGZj2TFE1Se9YKwjFp8NnYypIO6ADOTe/zj
zT3eXP/6MnHOgXihDaUU8yHp4/ON7DNC8VxDPqv5KYxOvh1tXXXW8y5iTEwJi9tO
VDBqcvPBmh41oWAoX9L62u66wJu4XKlgHq24ZVHMavplWn9sz4NLRUW9CXJDtPIl
41krFt27ECq/AOBxOU6mGZdYEc5VBrxqYP33SPQlnmDBrxb+19F3AmZIE+Or4VOP
xYr2aVWAOai0Ed+QUasPWAypPFWSXp6DbUVwa1pTSb4sFiGO1GWBLRb6WHm7NxWB
zIKBgL9uwWJ3AtH1TkoadcpuN6SLmUWoKAy0PxgYgi3Kt76Ga3P9nhlIIQ0Wc0Vp
vABQCo0wsijvuNM7o03uXsv6TPV7Ny15DNlIwTVO34aUY2DJoylc5m2A1/ERAFpg
LE11S+pbmoFjM0GCyrYhMnJiafFwX3OgVGZymhLyXkD3Wo9ZVAVeEZWe9tvck9gI
RaZPLS4xLHY5PZ52AxfTCbb7ZZqVt5uBJCcu5iCZMAhHKcweBmPana/Y53PdE6Q9
brvVdk6slKIJKN0fudWYXMwHhQkUB0Dz6ZpER3Pg4bC1HfyfrrLi25v7T1W8odqh
gl0wEZpIaw2r56zd0Q23IurPJt6GJJfrD4qc5Xfj5bpWMEnSZa9LiuISFVdjGBAo
T7cb/NICkcY+qtL4/L/Jf/2rAL7IRacrZnoPkeVE6g+78TtsXoDiTFhxXcoZiuAl
8Xp85/hcdFd0CM/zuEtL/AGf601/x6/rCchc/zmOgrwNIoLDZgQmunfRZvAju+Cz
5u8phyJ5qXqKnlvddDpDS12bSrXPSmNVLJKilQHy66RdRmO9BoViim/BQ45oYJbP
AV5wv6CVISdUX8tZcELM9CKFo73U36l1rXF2mnWlkmf3z56lOjeQ4T+AAmtIr4Gw
+cBi3nUSceNOWVyxRmWKgq0vNuhs6JqL4Utr0B/Kl6d6QX8iAcaiYjb5EFkgLGMS
LC5RtIFsoX702GnX2UF05YJSRPOeI3I+gAZ8CE1x43e2BylrGTejfuOJ+myPlqs/
lESQ9nAeWrIzVYzUvo5ldXMiK4OVhkl6yXCHXApjRZHeA/DiIZQ3XhWLwwpPOXDp
1VeIPh6Xb+AukeieDzyAf5hVCA/u6/G39uqt/nJuetel4lNaV9Fr47DDUr6jrP+e
E6uN1UCqgBnSZqkwMxkBRu9uOlT7fDSsPUfKug1rPQ267uvGf1RnGssuyYmTSQY8
aER+df6O+3qw+zqQdPGJe4YnmM30ChpcBSanfj3ijRNzMHqQNhuAa5JZ8Vw0EPeK
uU37c0eeedIUNButB6ZO+35zocFK01nKU0ZggwHoSchKoPHdwIiOoBLNLR3M7PmC
1/fRUDZSosRXHagL/qoW6PKxLRdYH6J3xVFCuy+Q1biGXVCg/HaDWzv66KKt8XOK
xT32QBrFqz/eLTPnTtcj9rtafxcyXOoeA5BaCgl9Whzte478m+aHOjuTqrDi9fGA
ROUSUStBwqkhVUcwNUuNFX0AYg5vB4DqjJ36a3IO+57LKtFUmIWJVxfFQcP2to/t
gA5kBSub7V+wnmekodBBtpG4Y6RgdIl2OmutRvx6U2pd9estAKnU2wxIsxTI0+e3
jF3jxu2DMcTMwlb+dq+c4RWWbNN/w8VxPMXY5ZdbN9ZHQRQ10gAepzwOzk3Hck25
VAF0KU4T1L4OD3AjTW6pJ+EmcAQBkP6h2J9GJn2ks2VGi6zfu9BhjFtsdXSprbus
mzJcDg1Bi6rT3kJpD4QM9qewDlfza2SVoo1E2XKrHsFkG04FLEttbj7Y37K6AKZR
CRFKmVpgmI/Fr5ik9NzN//PjioKNUQwTxbS0lrPxvxAJzVdlJfNwPSic6qWmM3H1
5Ad4f8fFEk1ZfuSlsRv7oTbnYtKJdKjmtiEZcP0BePip6ol5rpBS6C78uj1jvrMH
H2vjpnXzBSl1AjI8y34E8lENDq/xKCDlkHzrF7GoKQpzqv8IJJNuM10PxNBUKgUA
240m90B7FqrHmkdUJURWK/XmFlntCRMXZRANlQEzTWTwEbL7SoXFGwZDeSDI+r0w
kXRfzf5wYHIt8lJir0mW7HIljjpajUVE0juVtMBINHGhg0ggf9h0KvybY8224I9L
fBDAWrU7WckIEfnbzs8+s3BmoyDCApUqnKO7gMnjPp/4NCA7SX4DXSK7otMHc/TZ
Ts/Auh7Y7nXCXxyUgaSeHJVRAaQ7eI91yB3ZTs93E5L3184+6MUpAyUwm9Q/bhQV
N5aLjV0A/oHUPIkXyRqvS9Z5m1Pbj1ZJD9KFigHL4yaNItzBr78Zl/NZTWkQFHrf
OAbfPer3qX8W5/6BLI1ERPcMDbJqvH4WIpJhSUco/Oe++n8Q2J16RS6Gwp7fBlYH
baehkfDNQelFIOtKWeRhJBVrrBD/VhtXBUdFd0jlTJ0kTV7qQKUCt0Pzzjfmut6P
dTTWxpn34b+MAyVS6fk1G0PlHr3wJYdMXEuN5yUwZg/OW87YkNdB3P84vz/Gy1tl
WcXpKaEvWqUxVpg2UX6fAG63jf6IstHAeFNImFJcpEzLbP9c7DzkbgCy6aSWqQ+3
PTpx2cP1FroP1WXW17q0f8eHoteCSvb9e9UjMY8uY9lcEJXqywgi0qBdUxhSbSB/
VUY9M9vnJSNFaKHoaSyRI3emdJ5fK6SVJRgbWRpQQmL+mCK9jJ6NRHx/e2BBXJ20
9EQsevPKRi80o1NN1w3Inu106hTKW++9HSAT5q5Uvmq+M3U0SepTW9h0zxH7cv2T
/jTMrXG/KuZf8RWEHYSPxYBwNw7aXtQnZCSmFgPpU/3iJNRqy3AcAtnaCZAuDQXm
pAsUUGrcfTW2yPUpbSHXpL9PaaqpXf8cX53MFx30fZij8OChLoJFbO6itcCyN/jj
7Fwl56rhhXqyP5URB623H5bmLJ2tk2cp6RZ7bZtXuqN6aL5S9M9MUClEaNY6z+nj
28UKsaMXrQ/ydsewnEYkxPtKdqCNogGDUdsB8c60B5wDHc5XPHe0fdZ00xw+zbRy
pmWSddVWZYjVpT/nDrRV9N6cPuSXekZYsFap8CA6Sd7Lx0UbECC/JR50Nv5TdQmb
wjS1+mFxVhPPbFvMIVTdKm7Dom3nBpxgL8uWGr59IXvTT4QJGPqrI3fB0R8ksESB
E3Hp35PaOMW14hjr8mlzunfiu6z6EniqRRay3PWLmtYNRNOU5e62/TZKgDkQhqt7
JzxzhmdgoDrF988e8n7ZH9pfe1zN31YKxCb9xQQiv0GERLABxlxKdwpJHylz72S1
cxyO9Jt3j3iIQMoySM8NqIiMDUa+QP3Z+ic596x0wInURP3CcCndsikD6Rvb7SkZ
TbEC9cU6VE/nrmEuCi4rLPcq0RaIdHk5EtY7pt0nYwRvM9ZGkvVKkpAFdCI3pYqQ
qeuLA9AsdR63faoQKgSLgwgqF2QCZKP9T9+XPZz81Y3l1hJiDX6lvDFo8cWJgj/6
VJeyvOQ2MGTQ7fgkgXgb//XHU7bies0mHw0uM/ZCWC6GS1Jc/zB6eJkuNqdNHPdu
3XPA9cTUiweGr7e5vNm5Hk10iU1pIlN9ZdeXZ0iEcqco0NQXv07hMLrjKwP3cCHG
06LMPTkK9ihEFTN4fIlELPgOygfn0khNT0qP5ZE/S5tJxuO4WmZz4olPvTWQZtaw
fXSWUrZoBEcC8qbgX42AYMd1RTagAAdtVj57p7dlAeaAkgduYaG7Xy76qgE0SBW1
FPcBEJwBUvnHTyUEA0hv9eRYKzazLtSkA7YxQBM+CsL5uWkxmV1GOOddwXSrIhkL
HMAvwTZy9xCOujRbkbGbWcTfsqNWcgcVigR+0FRijPQymBSfoDh55Z/SPXV8A9xS
F/SpeP1lgl4GQPkwFN7fM8mPDxrxupprvVPdlqVA8CzIsfFUM+gT3wOh+ax80seL
MTqlP0TrtY0ZgKhKzLqDXFBLI2V5b7RHs5bDBQLyPAuz85PhAUgSyTuANmAJkIlp
ZkdtieaqM/8lB4vxHwTvsj6PDakCmmJ1W/3cyfWjjQXA4nM+7kv559cVmp1lpA/y
EuvbduI7jSo0DxPyIuIdi09MBoWOYxlqLpvtyOycAAuK52HdFTOH5DLLs6JGqFvv
MDjZvVZ64FAm3DW4JqyHWRPwRh8vFCWrNR3QpzxsFawGEdcyuFEi2drlxPBix/MN
Y8e0NLCyjOkttM9Iz2ghHAu5L48i3X61dqB0/sf1G/FzhFtfQ6bzp6hynBJGV57/
QcIWH8Bd6Focs2k/GSwTmIF6yIFCluPEbL4pAV7StUoJ4CDSlPWF9/uBoC0K8l+M
gOgHK2zr4lIksZ79mjeB3fFgBoPtcowm/yZQgvJu459leDaKyvzRWM8f3YZXMOwC
r8s18Jf4K7awe2oAYQPCkhVU9DVrHmDSzWPT5RIiMVzO6N9p0tgYO7CUKW27r0Xl
TodqI/mOCLW77gWp3clGl2hREqdz2h+GETEIA2x90h3092pt3n/No3+B6e2J1+w2
YM4fzommKU9h3Sz8S4N5B234OuHK/NPEEE3pQHBqMK865ynj/JYsG/g1LikcEzPD
LMcN0lIIvAPBXctD5Yx73AEWSaMdnxTr8iLpDtlv3l2PRuNZuxs4uFF6u5SJ+dND
XTnYfViVN2GljKL46FeeCwILKQHMJr6s9fEKjm83QgbQ7UviS/BFqXAQW1kQFo+h
Gld/WlcwewGCcZYxorsUHsz9nQKbgEEn2Bx2bZSQ79kAzTO7gCgoqkMhJFIWzTU/
SBZbfR1fq3jhXr+VZnWJGSRfnMpvBVCnISiXSO5kiAjQgPlMkK5VFHrbczdglm1h
KG/Dd86YH2zYyC0HksduJNRlfaOPD+yKLbDt+m98iibZpnhxpub9Xb+Q7M0W0Vrd
PCIvosdfhxuLJl0q1VQB/syzWbgEDv35FZY1NkgS3fyUsVSOlZFHx9CIUhQQ0YZI
Pd25R3DwS7J4sJFhjiMOSwPcFP60Ghs5SrICNTyfACbsXyv078dUbtplM8GXzb61
OSyY/2MITYW9Filk9WEbLItgLe9CiKolB4qwQBQF6TLYaVtThYF0M3W2OC3JIQVg
QDamI/JjCwbIEiij+ak6yeUMCwPYa2DHiZl6bQuuJVvUFFJmi8wF8gS0XZCaCuq8
mAaZKgiFQyAAWKJ94Ce3Cus+4ax6c50qIOpgE/m7edZqSu44T6HcKoOjsII8t3h1
zMPAXu4JdIvzZTUJ7vyzDiim6tSMOJxH/tzjVjjk7+jStonQNG8PPqkiqmvByXkT
n9XZy7ulxjp8+EOAGaY2eIty3diG60dCUzpclHaRdRlMNVQ0LthksOLsR9V1W9FU
xEZXzbDLhuNdyTFiPQS83AthNNuaKWw9UHDQKa/lQNRzBF4YMSPQpZHbpSNEej8j
q6h5sdyCM7Ak+8COyGmfNodp3gjj10mcywWZ+vHVgoQOMLGfap88lQwHKCSnZfm9
wJD4Jx+jXi90Doz2Rwd24gMKJwBOcO1nY4ohYrB88F5j987vhUySYtt/83v7DrrP
g8dLYFu6ozXXl4dZdCUBJ4Nw2HOjb/hZUoukTYeeqBj5Od/nAK+1eTOTisNiit+k
OWusEjeq1ZGOuJPtn7Quq9L4cF04S81BF46ayyWZQp0QBdOCvm2NwqNzPqtXZ3MG
N3us9DRcXSDCcCsoq++71gH+yq4lvSUUJB8gc4cFvFWrlrqLqzyZobNcHhWfS6JM
ORoNO+HBiDx3wGByXKY54qc0iYlNdl7dk9uOlt1FnFnWz+qWLRQs808O9jjpHJpP
Tpj6amS9Hp3emJlBl7Fm7TJCS2DoP2AE0jHWiHwVFockGXlJ0rzoWP2sBLzCexxr
rtsZ+9ffM4iRc0ukSOCIbh/wXxM8edV6uc0h9nCRDic1l9WA5ddp9KcG0A+QzNfa
rtUICYnFNOH9jlrPzWl2kk8vIy5cDNZskVomjbc/ObH8v/pDXrdw84w7DlsKsXX4
gFXvPvK7enQ36KAx1iJjLtyb4HDYiv7wT8TsvPhf8Mgg5qMBkQ10dg9rY84nmq+t
hqBvbGA2LAAA0104wuviLMxIGtaXornBoTaVlkOlCU6fmOnaXnmv7x0rRqzgUxYD
VcikdQzSyNPz5AhwHK5DHJZ5DEDgV04tmw7pZ3/QkUSMAZhGtt5c0HIX/XaHkI2F
uh4C8sv6lnbh930mM6qiPCxUp2cQNsh1pP7Vmmv71w0CljGfBXmefj0D1R4mu2dX
eNeNjYJcwMPsGfzvOci+onh1dcT+tP3mbqUdDZa+V1Hjq+jfGNhIq6rzBDg8WD1A
Pvmalni3MuNmG9cetM9HcO0x4fF00M25pq3MYSzUBV0ctkJuJZ+Bg1/KwaDrT99h
un8GhRkHck7cbcCnf18RtVgPOV/4NEFT/a9AZK+Jk2RRVWcEv7lahHWYjqOmgFIV
c0mxucwjqI6jf/xlhFbS4WF97DBRNnYip2HHevG/m3NtHVQvtwSbVwQtRRHIX9R7
/yq/UaNm85n02Mfur3ruQ3gvcdQrxGJgYfR+qpBcKUGzxBtqTlwS9ZjB0dZRp96q
7uhS3DLGxGDZxFDQNkfVZercjLUg83KOBoUI/y72pjWIYPhn+a7mZzVby+9YuOZ8
GuLfOxR3RBK+WrRmkkSNv4xV58UodXQApHCpOadn/n5ej9lKAbi7w1MToFvZRvZj
HYrcPAXSq2cP8Sa91hnxaopWiKsIkypS7PuTh3y9cDM/2uvrhTMAygpsfijz4/Xz
ATaG935jOfaqxI4dD+0gJ/Hv2m4+SweHjujqqfzKDf8j38GQfWXKaZjGW/6IEpVu
jXkUGBiMEykr2BZJ08JUEAHwGzcCR0G9YqUKhifzK1UmbDPmgpjnT8YLnWTfsmoZ
A0V0R3YvfAROv7/HDsI7XIupl3LWn8PIG1z9F3imWNpa3cpump13pVwCcFZlRnEl
ORLEG6Ps0QI2pdoVh3+5TXi+1DOmoOHKqRULYPvqne0P9yp1v5R1LlPPr0R3btLr
TTffCuLUSpCEZkp52/K83KcBVH8YsCr9eNvYm43QjE2C8WcLxUQt1iJfJ+PmdgaB
KfOs4IIxiYVk5gH0eMg2FvyiN6lxc7cbC1qpePfuG75iJCHAAKUWwdgVnjQMzDxK
58CcTuL0DMQW2oMWuDzRAuynX1rB/aIglvRCSSnGphsSam2h7YHrHZL+aRCQczmX
Pn3/zh6mDZ6cRAwt84NGHSzScEZ2IbZGJpHLdXzEwoDSOT6kSwg5rc1OwbDjmWun
uBHjHoCPonJWVSV1Tva4gnKLcXSV1ggY+VsY0MWvMQmGa+P7vOv/yF9v8Jw9UPr7
k+B7YfliwNIFD8iXowCgWxKANfw7+Ex0L2D2q1RJvReN0f7VL31TDdxbTkWV/tcw
sGR8KJwbO3geITO2/eDCmXodmKEjz9M7JaBy1W33nukp8m1TTyjfNEmM5MvhmH5H
5ISLgfxM5lb+GqWElmbUUE7TGPy6mQbzDbU06M1btuSkqE0r+XwZQpVpZ0vUJHGC
OrYj8ZMc9C2A0EICL/ZVnjk2lPlNHsKqQZ3v4RuI7HaxCeAmHLrCH9UmFE8t/PjZ
hrzP9h34djlnrwP28YkBw56GCTPvqVFl+2G+lMJbFxY9n46dN2IPxPvWFfKeM1Ps
NgGvJrZhI6KFTxLFdDqnnz74PiVbmfUm459v5K2uuDi9Jz0LsRw0yeYEP/6Pn6lH
rUExaQVej58jDKlMN2DZ9vV38dITtq8HQx5MdabOyTg5bBnW3rYdMjRgraJmj/vX
dSX0L/tPhWa3Sj3DShh6ir1OpboFulo9BuMtNtMJevTkAD2Uvjf0xRZpdDHiHV73
c9zmmLZpno69V6Aln+znWnw7jEIQJn1r3iR6DalrUpMsqxOGZ6iuTk5ksfs7Spl2
Hezl1vCLSKBPkUAAW8Vq4ngNEeW6pIoWZ2SF9OdMaN35kTbwc8Ifqdnv9qGUjobu
rV19yPogzAknKY0BEBO8o5kLEtJ5pVOZNWAHKxge9NpY1vKbsxRjbOLVcqVY96UL
fAw5xt+PGZmYUxiondXiz1V4FeneQpI5y8eYHzSgT8O732rwkbioR4JSwLVlh5pA
2rs5w0Ra8GqgM4gCKvDW8NoYTPi724Cc5fVLQI8POQNR+llYcEycPLoDmTXbwnKQ
a1uFC1+zyANc90xIZ62vzr/qXIaKcmaeLN37LBDrpHwLsBe0NpoJ+rCd8b9Yc0nP
FV2ndqbdiRHSOH6N9AFoBrMyuEuWpOywTky2S4aJb5rfQgnKJRTtR8voVdbeCdXK
EPUxCjixXf+vSLQZdlysOQd0+mDeS0dlytVHDslF2O2a460sgw/JwOE03VlJClw0
cIdNkaHelVcWCN+17H/gMnuPTr73ml+cyAtRkU2EHZPYAi45NUY8MO5HNNGSIlcK
IPTmDufbsLPZLqhj+CEo+Wo+OlY1ZasbaGe1WWDSptlDMApkI4SuIpFakdOgaNCT
42o7BPBkdhtLA51G0MB7Cr1Y1nuo4/wzOHajr/xnwdBP/7sPPCAWjSO7OyAcoPzs
XVNdC0Rru+HftbiZVhovWTDObbhN9pAYSKmQgZe/HMR+KIImsuoxiPz2SeX1g9gQ
J2SeLiXNUKidVWH2pbieCy3JpcoESK7g5tkqgEBqExgZEbdZp+atP35WKMb62+0U
dOZIwfffSNrpJ5IfPhSsYbqxjKS8yqOZuB251uQOQlPf401HB09JhNAN5fRLWnpT
32ZNip9Rq+G5jDwVgZOgLohkEZv+hL38ZzoOlXS6PZHqbkCoY7b6T8Rg53oENQTz
7QV7y+ZInM8gvev3Jk/+eN8V1NFgsc0u60kwkPYQQ9AlqZWyNZRbxA0ZUhO1/ua9
KORdhweZ76s07cpk1yZ4gj+jdC4jkWI2FSYbD7fxxTJbuVPMoHjRF+EZIE+fxCcq
aYKviv+yYCwA0E90BcjwH8xSxRIw9exGGWulTXFOVw974mTpCFXljDnWmDADyJeD
Tdjcvgq3i1+dXUahGU9N0rq64cgEBaPay7b94C9rp+BHw4LAC8f5hoMCrQGd8Zp4
NJQ5eV5rLKCJV1GTJngixYmg0PQN65jKEeGSqAaXXM+ghnd4mAzTskfwrdeeCKE+
yGyOnjAV3A7baR9pkp7O/63Qv5kbqOXm9Oe1aLsG7X3N6Y/ppZMySeKbRb0mG4Up
5+q+pZscf0gL30mB34hSEJNCEcKtA/JA21AAz8Vph8t5QEAKuW87DXmE/NGCQ1WD
PrYpy2slm7FecoMYFyly9kj9mUPDudBnlLvIaP8zbYtbpsLwM8/pTxd3SjFGl7Kp
k4PVOi/HTZsXAG6Sbs6eKsXsXfiGjeT8oQq29rOcXx7gIdOfP6SIuraqKpvRB0hj
PeYABjV5OJLtroyVI61sMPikYs7umu2e2cn+R4JFoax4tbWnZfuKYqhxD3+oVScl
JakObg7AlhGWcebzRMzmQehpyCHwUvOpt6HM1t9i8GWmKa0M6/AzFUKBEW5ycSba
O13+sTobRJty81kvHWRG2jlUziXKaifkuhp/I4cF8SjGCKisZvpqpY3gXyYPfQFt
5d421g0E8Vjo6jYNe2juSq4GOtQyh2ZBhkWbMo/A34BeD/a0OqraPRvN8PKKK8XP
OzjzLzMp5SL8hkM1y19rimPkxjZHRBB+6zo0+ma9GuIqfh0C58ekuVDhMXraOsri
HP5c3U5sQFmfxZqdpjuXdpXAMIvlo7LzdvgwH2UM7Ya/b2VUQVqvpW/4EkmUhHxD
AZirf5RAC6Sch6vMLFKkMFSXun0KvYjUqSAqnoCTVTqqNqJYijXx5gBR56cxQhk/
KSDVG6ov3VznuD7Q4P5Js9v3K1UYgeSYYk/4Zo4s9bi+CHERWx8TTpCSp8mv3ilC
Lhk1AaCxhS8tr2x/Vzu4iPVQOpHRNo9kqQQM085PUWwKW/NZLYXcq18c7NIcu/Pe
fG3FTP4lUS8iItptBGeiX6jSnWsgwxrEmUESwprKeE3PYjy3Ksj/0EcHb35mapUp
SkNeVu4KHnFD0A/hzuYw5ZjgFB6vADM7RtC55k5qlrPgf4pCtf51k225f+Rs03GG
Nb7aPu/mW5PYUarcCVk4QIhr2PfIZKzWQQ7YLFpUgYX7hPMxy1BWeAszI43cA6ar
/qPqf3xjfrh8KT4IsQIEx2FOf3VrJsTs6/5+BiZyUvsPI2An2s2EmNBwBCvHZEh+
ChFvf00Y6nPY+TdTZm0QkpJfDogH6XKJRaj6DXKmfA06z4TqmWTafPLDWUcVhqiB
ECtpKOGN5o3JCe5CwRw3QxfeoB8VEu5eM98UnWNP8vrQ3FQQ7vJ3OXP64zKGyund
qQj2+/cd+bMqdNoplbKBvxggVWAbkgx6GJnqmpwAxOagt9A8iNqXoz/gB3YGr5v/
LZjm+04FcJkNkWmWaFH+iPl/C849AACOl2djI4S/AgWjCJ0HPkjx0y/JrCoC64xg
AyOR3EtAVEn5QKQN40JpfoFTWQ0h7oTOj3vvzgfCCuub/R43HTMygs8Kblp5TU/9
g0IzMVkDgFbC1nDMSNfslaXpb2AuQWtbh6uJow6XLn/XS8t5tEVnIvGe5N+xMzb8
YRuT33C9UN5BxbqWCeJZxdlzQj3GOTfzLloenVd8T10f24xWcaKsDwunCnD3JGyl
6EKm26pb5JNq+Z9YHtH/QnWRmra13XfJbYLiQniYI2JOvhgefZY5ckhKz4ip+MVv
wqyHsapFu9fPz+k2J/fmy7TmND31fsHcJzLi0wUmDpGG+6rEIhrI2g5YC5SNbkPe
t9hcgLwWx/4tKfKzs6z1tGM/aVM7nJA/Asf3qq8myejmJk8SyOsjVpA+28f+MSbH
kNTAYb4/2PNPS4LedjIAcAbBAHcRAzDod9w9S8mW11nAFeXx5JfVExcV9skTOi0k
HW+9TOKQIhnWiSBV0NV4PcPXT6/nuO6FdZpbh8Ef4r3ugq+hXHtlAA9atrwNdHew
ZaQ2KvNu6Q1ABSXRnleTT2lc1iVpkD1Fer1JBuuTWicJi55iUljerMDnDg/RoTvz
keX96J0kNCjy7m/Rk8jtd8F/fkxRRLyfM5nw9okCxG+F12mVvv0NfJfWXVIiPQQ5
2UsP09vOnXfRqH+zjVl7mdejaePNW1AR14u32kmT97XT2nCLWESJJsCrwNIQgakS
gHd4FxdG0pL9TDVc6lT4tihI0J/z6y68PcW5jksyXxy1ThHzKHyyNkkDYqXfY/Aa
kBT33GUDXTmLxQo5INITifRN7ALSqyJVKZzSXnY/2yA6R7RpdeEv3BoQGUjyxeJc
dq1Dp6jKMvAnvWvOtjqHKuusgj9Z6/lmBUnKDfg2aGtc+c8KBqyGlJgJ5fDuN33R
7363m9nP4oKzlE5U1TZQOA6P47KH+fqprFV7WRVjKf6623ghgsDqNNY+Z/uvVoat
MpwxNu5R9gqnir159wLf1t6Q7NEe1bSXIx3KHNCLSBGWHH/BnJ/a7O+caZAYjx8K
teZb94ZULNnM/nV1ns+qLCd98HeLAfKLk4paDe5j/Dr8QjlJsD6utmNE4BpcjxCv
LnbsZWMUQz8IEXvtP1fhgDcm/KLVjt5t3vcGZNGnctwSGLyxQ2MQLVxwP5W0jyEl
jAFQw6FjKvGWvGm/UPYkRQ4Z4bMkLQorLMLac7ruOv6Qs/rjtG+MaHEcDc5uo5mZ
rXWvuoWDnn09GCZUmK2qCdLwcaYHj+3oWYIGU9XJ2GvP0g3SkUsZIaP6LASALO5E
9U9IsdJY4W5evyZHHk9rUWH0QBbvgmj8jUy4IxR/qC9TyPV3PJ1riZMUxZzBxrjQ
IlgqXJ2M1S5ociEJCn49tJxwWvXwWn3/fx7u5eU/TANlYNRJwPBmGxwg4ohPmVPE
BiGog8svAWvvlxrWIBKs+1OHyBaR4aY/PKXL7MbOd5WgHoSpsc7ENxc9mZaCTVat
H7lHxcMtwgMLbuuR+Ub+1yuDAQ2IS3zmNzone/LsE+8Ul1AwGbW7QcpgeIjRkD3S
XO/0eJyU+buEwESnx2V/eKj+EUmLpvZD7yhiUl/1H9Xof8kZ9FphjESOr8+oSziv
q2mHjk0Epc2sjMnrPfsPcIouP2ws//M+aRN+YVDc22oSGXhaj8e2EFK9xIjjsqR0
JLlI9NZmtH8MTg7Zpxl+MaYZzY9kLGRDTnl3xPJx9UtVUulQ0hlw0tvn16qY+UvL
aCV0ewaGXuGsCWv2ZYEridapcg2Pq8avvAN/Elk/e1H18rLoXjGceLPhn4Pbk4t6
7iVsLQ5NVZt/PyoDfhnByMooeGn1uvjtuoVag6az3b1y45vBSFqlfYEvST7H4mCZ
gai/EuX1p+lFZBBWGlPwyD2pSvmX/Vb2HOzDciZSoUbfJYK7b8blSMOfFNGsVK7z
ujWcmVsdSAahgS4Y5+UoXFW5PkYO4PaWwYuk2mjDPEt8hz1NLmlje1lHK/U9OUCH
lj3r1EDB/Wjdyc0NGjvqdPaR9WSeAw7yJzR1SBkl1uLLbyAhQSOynW6QN5MvjnYW
4SHo4LSd0iX1AydboaVhauCD2wYXxaSHmRIpH3tghmY2dbWBCL8vePKcc+/m/Xn8
mIX5OT8B8m7AGUZ/dZfgN+AOWJxRECJAnToZXADM6lY0mNl7/WNNy/r6Z8khRx+3
ZPECj6Gjpi8sdb6r8wi+P1q5qg2kLDefVoy8LFsSXjeTFAVodHjKMDl2tnoM2Uzu
eCK8SGn3Qm69oGp5kjL9gXp7sk95hN1yAf4aPX76ZyEAUcxPFcZCB08RLYRLiy12
eT8Zo934ujAysAoiBZdH1YaSUOWbMpzp+/1GuyM7V0rLoppq+93OsvN9RndvNF6l
Gnwz79oH7cl6F8u+/yE0Fakptgl8QCxtTB0sADZ3Uf2VdpI0G9RMTsteMLZ1ck/Z
e+lr+vXHegQusEzQ8S4upseOxCx9HTOJdwj8jB4MrDKmJoJ0kznghJOOK6hC2gNY
2op3M/cApUS2QEoO/V7d1BmLoAu7Hb/c2S+yRTHgSMo3kwCc6bUwJBDV2S9FeMSI
ZaoKeNbsemBBrvcUyVd22Rn9704+6u90W5VJuTadCDmMiubPILG5OAfEy91sN6U0
sqfKGh13HnRQYisvXplbeCzkhxp2uAInpe+1GDzEtVxPkdIqknuNMS9tvu5U4KuO
+ubuH0VWBmWwU1b2YYFN4OpIC3LE49kT3qhuIhN87FIt4gvOMyO5eyWz+2Ixrk3s
jWYOrYBgIArPasmv3grcGOxTsYeuUtlercV2Z4uXpM2galvy83//TDfRD6ZLy0TH
Wv5w+8yj/rLwVJhED/HW7XK1N3X0YBPHXFhdMPbzkrkkfAl0tF5+VzWoG5DpeuEb
miyk7ptXx+KYOOqFBSPimSLZ42oW7zofGN1p/4xduifAIaTM53VhQPHhIXIAALPg
d4IL0HEK+4G+5Yfr/u7iiSW8qWwSHRMy3dK43AOHHhAhEePXafIftf6x7koJpJ6j
TPAav2hfKoDL/uLAeiRMGLfCO+NIft51+Wi7xDMorncasleTQWMsm9Vm18Q9mZTa
IX19nRySOt7dlo8tmiujkyW0Z3GXY7wVpn766ovnJJoMnkuufqC2aZR3vb6fSGZy
kzpDSwWU1R2lRVQlAB44chpKz5nxgHR2I+1RPZXxIYJo9k23AGCWO8vzXo4GSUbx
IC60AdUh3gW4tij5Tyk6oXaYv4iyPwBUks8aHLiCeuB+7zQcM/Nj6+23ZF59HFNa
FCgsanWsRYQlnpb8iMip5Vx6A+aay62U6yHxBxNwufdbIGEDl8vE7KztycGj7OeQ
9LtvDfN4ecUXdqDjriWOaVZ9YUWWNnr/cY/LmlAd2Z3Dan2Ppz5BgSnQe7y7BQ/D
aogYjVB0EVU6rvS0UxDe3pGzjAmsKXESkIo0HXcOjvIlLEyFnPLvDwn80lcdI8IW
V16GtHH2TYSdvDgI9IwEXGv/a8wepaEQQ+QLsQGYc+Pn/tLh5NEmDCNq1EaWe+aQ
o/nLhU/Wf8oPDsUdrp9dVRQvJjKBtxfr64f26AYwDErH65jLyCLGqMH2tnBUaGM3
WauTb2rGdXJb/JrjRfdc3NdJZmHMUVKUkwpB0z1kSUoCv2AQRdPhRjN7U9sf6Ssh
vzgKF5oY4X8GG0eBgz0Yfjk/tFLJBPUFsCKnNzuU0dwjF9Smx0FV4SA0Nj84G7cx
jWIN6aJv6YWnjY7DYkbW7W/PtmYhzKX0vVMh7rkiYtMX2/jgfBofpLYb1rNRcCQ9
KuUjKF3chO4WleJQgLscrAwS1YoccCKcg7gGcaEuGRehDEyEOtM001JdpndK3F28
ptoQZZxA/xcR5mDUSAsXCXrMYS0jQhJp+WObyDThjwhR+UakdWNNq3r/lCNDShZW
RketkrDHgNgFyLXCjs6Djmx2y+E869tAXDRFvwxyP7OfH9zIqAwv5aXytP3MbqZw
iwD6Dwo6qTKL6ucxHuwPRFxyVnVOYYFu29fp8gaqLPIRXs6hAMHBl3IvEvad79Sw
dYRlccmiHRw3pvAf62cASH0wiN1RK/+6N17P2JlCv5/JCyssA4YNey9BjDuULeE8
5wzxg4LzhLOBL6FQwysU0gxz/sCd5Qqbl/7mt5BHNJ6IYJt5dVR2TbphDStV2GGu
2eBHGDbhCDOb72TSHJF44pQczlaeviJFNEtoHVkIFQ5jS4qgm6a3bnSP6ExO0Ml2
rt0F7H548y3dtkSWUGXiiXAyURB8Z5LFqzDyEM3bVVgQpM+JYyrrW6xTRVwNa5+B
EuyDZtfQuwHvNXLAXzUMdP1uK34F1Kam3rvbLYGu0vnww3QdjpwDcDEo2rU5GNKz
bK9m/PXZyv3H6MvYfTWPLqxoazST1FdLBX4dzRXKNLi0hbGvcQvLWvXT9deiif8p
FfWeIsUjxo1p2SJ7zIqCsz/cIqdBY20SPIJ0l90Qp0FvfuUwg8K2jEFxgeVwMYvK
78N374SdPSKOMNxANMIk3w5j1V39+G707oBfNcJZY/uC8fh1vT+yMyIFBgoaMSDi
eE/DO8Yc0oMAc77OKqw99EnZ9uQgWKkj9LcXcLFLeyIABNHbDcFguv02iyE8T9tJ
FbhYdcYEBCcx5I4y/WI1z/EF5aJytg3XvT8u3PjD4dDFPKKKoiYexRGKE44dHXgA
UcdmtDmhyOF3RhcWVjqEwOnzB3G6M8zbynM7PAAk+Lh/txteAscAa0qeIQ8rSh4G
oRFMgLJb2SB5rjrh+JyvNmNh5RLcCpiI+RTl5uehlmI+6cuCvLWnVBwz9MoC1OQT
APZ65hGlMlM2jsoO+D6JuT4kvyM9ES4qSciCJ2DE07yIbJmaRdvb/WHr5u7+ETKr
yBVkquiNwyQS2QiEAzKqSNNKfbYoeaAPG07Ff9J6c1kkCrAIIMNzqaPa+ZNwBeG5
w0fbGpri58H/sHbsGohICWSuksVNOF/6BB6DRW5IKF7BweMl8KyHFcVsXdBuh7D7
MaPGZSjzBDsEiTq+KEUrfekv6eVxzBNOuBeVf64T0miMtP0lBB2buPz/w+55rk48
Z9utiv/DVAb8th8lJGOhX053dECgEzCwhIktVE3pkUoiuS/sZY5YeWOeEmgFuv2D
837iVMJy5Eepv8QFmWsGaLqw17FKHOcR7UTI/tha/fHVknP26jFEOQ1TmlMD27t9
l9X5f3dHIBSlIGUUyEicPRbLxANwdmXNCTv0jr0spbcRiQtZun6ahfnHFZYLqYp7
MLXllWFqokuOHmU60NWjtB/S5qvC2JmBjRcDdnGWyBtk6ABXXykU4694avdHDquH
HKDFNfYl68jhkSmLNDsWpMrS2RCoC/WOHzRb14j5imN8u5t31fE8S6uENQBTW+ul
c0LCgtAp/jcCjPPtyENSDZ/kbaX57D80yI3nejd3NtM6HIKoQ4QT+4jzJpjjZAXs
SgGJxJiIXbQgsvDE6r07+qGQ1LzGf8hxnYisqJzhQFCPOr6IB3J6BtmujqGWJb08
X24F5l4oW7oVwbsFY7iqr+CiaQpPlZespvjrybYma0fQHVyRv1iu67ae8Vbh4DT+
GpZmQB11obbTlOoTS3N0UaiFQT2yd9kdB2LtaupHBE/qxeDVlWEbvg6GnZDFihH2
eBVewrr8tcKhYkgNRCdVET6uC2ImYOYnCxob7OYfszlIBWm7qix0gtTEv6EnAa4V
g/lDkABni9TQbFqB+OH0t1UaF/4nV0G1cdw2pUArxEtam9oD6TfYSMOu5aWbr9vm
V9UHbMnIQq5WpjybT2LKJYUv4ueRZRv+8Gimbh/l/aDUQQC87VI9Llu9r4Ngs3w+
lF0GO6ETz77gaa8rdrjtyhM9h0vhybE6RJSoYSXwv9yNxZCf+6bBUTantiMperL9
3wcFEnimSlp//IR9sH4itzB79BZKL9VrBv0izcGPbJ8JjACaqlyqydm1zKttLDjd
1fWIkDQe79k3X5KS4H3c64mSeiJxlo3fOjH79nz8Me0bSNvImnL2Da6WB6MEDWmW
kMroZi/ZSExtDp33RdWTyhsJo67HSUCfhROdPZ5foQy50qjpP/SzYOPxNEO941hI
MqgFDjg4ya+DSHQ1qYRl9uNFDnJhWxZ46ROVkJAE96Vb6syUtEIIeyf41+NTiUhR
BVApMkTGTgo8j61yQuqd3jz1pLifRe4g81Jmfq70KV0Qu55Cm+uYPT/NE1D671Hi
BQRjkWo1uNYkcyhhrGcTZaRVNuxwt5NEJb/OPibsz151uS5w8HYrZqTlxAwuQP+S
L3GyUAD+c6QJ8AyJCCNwEQ1WTuwZC022HdxhxwkSy2GT2Hfiik+/aewYmvwlyUv+
4lkwnPnrGbdF7gBZ9EtUlnv8YwxzkYShGaSWJhZrxKY1zvKTKsxpcjM2v8q4010Q
u/8ejR90fzUWk6SgcUiU/T58S0nqO/SnIZRjo/104LnLhDu8CsyJKGfAIeAKxc3F
mZ3/T+eaAfDexUZBr0XB7qmM8X8JpbuLeRwPdyRxvjAPWUs9hxC8O62o763AvoHb
oh3Njt6cjZtB1yPmPLZvBS3ZrVLYnnZsXuwkGKQhko7+XS8LBFe2E3fnlp9C8RDv
Nd0HrImeKePE4vftcQnOVW/JGEKwdPNDcarqx8o4OR9Cg0leg3kO5IGqrI4b5Fhr
dr++DHtvwHv0cH0KXRn0zGklzSFIxAIfLfzzDAO3JZkHse7yhKu2dStZLEUHP9/a
at6awceiRONYdZRPiV7B85XM8uOiDpT5SuRgbP/QWc7+SydcAlQNdKyeevzxwK47
fCqHVnbAszI3y4KIC3lu/nUIdOCUDaiJZjk6i6bXY0E/P4tB+rhaPAKUUukxzuGB
Wzx/LOgBeGanMa6485udh0raH1heEhME/u9huKjzKpNxBMQQlzsHPzse4TlVGFNT
inKcWb/M7VQ7gYwAI8WXRaWswZ9JIZkrvcDtOA3ZxZl8ZFPpp2Gmi0bcmYXfBzuA
L1FtY0Z4P0QpxSm2rc1HK1lHqzI53TIOXcC15t+j2gFYa7FQSonHNcc90RMNRAU4
LzqfoKdXe+pxJMtJriFV82ZIFhwBCkRuTUs3qEVBrOAPlCx0JfJHHDVq4QI7GMeU
4aW8otqOTm0o7UmukUFFR7fFR8aK/SFUl+tg4FNvWWUZ2zlu9kdf/qS1lNBSM0+J
XnSqTwdXPH42QMiQE8zdsZOuY5s3dSAFDp+6ybZnxfPcOqflNuZ5MYRDV7m4K+Xu
LIFPtzPHn+cSx0PC9vp00a7qtbi1fRoRMoB6FGNLkOREqyzJzNk7cauHbrGahtU8
VMvzo1jctxyHEgLtmoMonX4nuTWRwmqI0M6MzNflUF4iPSqmKVzeV9u+LVGCid8O
2TV/8SiZ5C2HTL9ckVUrLe405zuIJnjhyjEr57nNL6z/toSPf4a7gAYzukuOdK8r
sJDzNLK+tyLe3s8Qv++gpn3IRUTF7iqmHerlU4jQEdjnB45WHYlH4l/HXTUU4cXm
CpedQYSMOdoLHmv640Syny6hfl7I8r20P4AZgWky43JlUTgrzLD1f1c3Z2J7wtjm
PFLlq/rSTeN2O1ibUuTJgJNFrw9PMDoCMUZQuDYbjyM74hJ6Xg5g0EyQXozRzE3Z
JUj2DNWO9/vUFjSlKMiwfEfgW1WLQoGO8j6y9FhHCPYu9PV79PzprUWX2tnjkHNB
b7kqkR2stjfJhjw2UZXprRnoFrbyCQpp5oUPS0hOMDN2CeWJimOth66zCVFj9Kk9
uncfkdL0D4s3kb2hdpGm5Z/lOwLNoGF1WMmeH1mJwJypcqME4IR65iwEQLa7rb6z
ZRX0voo9lX0NwubSLlZaY8bGRMjpx/u6e6SHbJt2mIplzwPCGFXpN8vDEXMb9S+e
/Zw6muNC3xNqmRqOtyziHRpq5pa9q5ZQDbR8PKyNfczxU1eM7qAYEEIbkRhrk9N/
qRrcfDEDTX/Yi87zAoKidG9w6lGZQRCB0CY/107YIboZ49fRVMZokumLiyihHOhh
lu8OLXOeR9EbJ+omtPH62+wFNxj3b/6Zg+Ianma2kRMU5swaEaZBXuJgSPuAPfE3
KClODvX9TGJmZhjdOeXHqzas7T9RxsTCYe9efokp24UJZM4+CZe4akyf/4M7aAGD
bh9uPMu5qh+bFFXgIK0xxrHfidnTxefIWDR9guRPfwEjWinjlM93HfUL+8wwJIEh
HkB7Me73MIojVY+zhKbLTPtp+ErfS2Pbzb9qboHoYTZwXxpjcnNA0hErmADZVfUx
FGnJzFEZ2t096jIPm85WDoWSjEZp6BETCy0kUHfLtiRhQe028PcOhi6TT4+FZV5M
TwozjO/q07EJnpNSKE2NomJAlPL3R++iJUqjI/v5ns+NQE97fbl+5LYSqjGCyk0Q
SBhD37HieR5m6Vhh1myvqFH9rsG3NEDaOYmeZakGL9KdqHX8X8LWNej+tPKBuxNN
PGxl/hbteR7Bfe1WuFek6X+hufL3e9VzWF0Ige9/91W2Tm9U3a9TwngXWw26WdD9
EOXx7VgV8wsnRuJEASXiwr282k5LpoQtpLJ0fAr5Nw3k/AiMvNQr/2ukTDTknia5
vlYf0ExvOa8DKCkRSjN3QLkYQQnDgC/IU5gJx5jQBUcLttfoxUYpij2FEN1NrsP5
6a0dShGsQNXgbiv3MKMcOKBY/Qljxom3F6t6sXjowronmpY5Vm0ak5VqehQIBnb6
XnYvuaVxzeHh6z/os7gvvqDUHnNVagOlHMQfu5cXfRV3Bcv2of6ifwMoTs/pJeEv
+COjDFPXHDIaux1C2XA6MfzyIoiurNwz5NalQCZ4cxuyCUqbrXYufATACJZ9pyb0
MPJUGZpiFmHHJswS2tUd4qpIBakY8URlLpfG61Eff9lQ30mHVxeDQN3C1Aq4pei7
4cciqd/JQFvYL2oAlDhwLJT26Lh80GykvX1O3BVNBJt1TIaF4o2s4h4Uz67ok8gg
2Rdk7Ujghy2kM0oCe0uZOLFsMXAbHh6ePnQdcY2v8SfTjrkBUJ8wkiqt4oS/TRjx
MtksQsowJzjFCyQxWmeDyg+QczcQFCfoZ5uTkpvKqYAni8mZmt24tEf/uWYdacR/
7z0ucbxM2EuUpjKXHfSxD+V/Gbwa7rQ+DwiCDo7A3Tn90YaYLFbHoqJBBaoTwKFZ
pVVJG9ACiCF9qFFkLop3hc9tUwJFcEFzmQeLujp/N2RSQC5ziZXsAzakLXfwQgNL
sujM1J1licdNFMQXke+iu91Z+wN6yM/MPlYMOBBk3e+UPhHbq1bzw5TVxxkApNSf
dH7QOQIpsToqvWyQKjgacl+rV/glSu3VZDLvXSPPchRz2qfMF/qH6qC89Ftz5Dh5
DvitYQulgyNRXBNsdH+LvO3SD+GWavSpD8o28s9j1NqmZIBWvpTSwOiKfzJ+yNwi
gLdDtPU3hoiFYttk9zza0/yDt0RNClrhTosxxCq0dMq9Fr63cMr3D7IIpdUhibxq
oNZKpYRYaq7yaEDE4zAL+4UyPWOceQUcZqkuF19zdXrRG9k+8crubpIt63Q5WkeZ
hg18pGGYKPUsSJIFLJtK8R1BVxuNgWMR+OmWnZ42XxqlJbVm4Ay/nXJL3o7ToXFc
r1nzGQJl5WJwAWM93J4WOE1Lwk6BHkjRH9rLipUyRaPuA817rddjzwnUV3hbgHZG
n3jj/Ancz/HJoqv2d0PG6LVzMv7uE6sONIOf8yc/4Y30cfpDzQvcj2zRx1kEbbfW
diYNGDKociAWn3VsM7lX2qrkEjKig+FVKn+/fPCeGOU9F1TrK0wnYQs6jhkTyKil
cD0+Kb1QM9w9puHELSy7nw9OXTxVoQz+fyAUmgXJwEviC8+eEyDJS6UrvNjneO56
FxQQq8A+mrCGjsfKSsAfZh3Aor8eXKQ5cj5FrL7AuwUBx8ZP2A2IeUD3tS0fSOmH
oqHwd3R5YE/bEA76Robdo3bbXhsCE39fqw7cBN+nq9/bTh4WT5cmQz3PjjpyevB8
R1H/bBcqBKGUf/gDXsxbKAT2NOux/u5Yhf06kxLGi63i3on/aYUeS2X9odq/fZAm
7dfKxrzXezPHv7NzSIU6PzAClRZx0FoCFgV5voQUyAhq8o28jmLlsP0olgAk5eLM
/+JqvqVuvmEx4O2bnx8E9fe5U3ZLWaxvT/WR2+D7OlxhbBhndG+cmjZ7FbA/5Siv
mWkKUmqw0LEwXrc76AQcZ+0Z1a/pqOL8vXYrm4acNcbpcI87wqd3UJ00JZEM62as
lycZ5tOq8Kgkx0yCXnGxSfdgqG67O19jpc3ojmKxe1RJ0KASQPtzxQfquQtXySY0
mEoOxbAJRtQX3CPiN6jeDzvaIXcSr8LZAR0orldoAsTyZvt4UJquDh5zH/9+/X71
5jZhKbv/jhrLmz1NX+XoZs62AuvlmCUTLtydDEEYCsPYy2YSswHwOKKfVJJ/pgla
Xp8jJrDLR0aCvC0CkS8PE5iM0Z8sEngI/ba0snMJRq2AA4zgYIUvDHpWVjb/2VzU
BZMVBlOQTRwHrpUTMRos456+qeewxYyOUIM3g11CQDSfdAnSj6v/nu4JHm920yDh
Xiyy3+xd7BgzlTrOno5erj11P1l4DL5zrb+wbSbfmJFWiPSv2T0JlC1WIlj5tzFe
L+fX+zRH5xDQrCebosHM3LrvzS8lSBkJXXVGzJGyKG+zNZenZ3Icflf7DdpvjWss
h8+5w19hSVU97s9+HZlpI7gQsgZjl828xyAZlelvrvcuR56pw2Ir/oEgKYMVfWUp
qY/dlCfaTprzYBUTzsGptKV2HsDHzce5sfhPAgL8vgmodMS90nkblejNh7213m7t
lm+afima25kORtiMxjqxMHAT8Hi1mguniZXeBA3vJamseTSYMmoz0qoCT3oUAwbl
b6PYo7goUIXHrbU8E9sSDnDDNKDBAUGwU2BCrc7LBDSlN13WV6AGpER+AQWi92vm
ADLXhjDZXrbFcEDL7gV1MfcvXjW8tNmV4AK31yYKfIugpEilCHwBCY0VbIpCjJdl
SvonL4pBnfdBFpNXrRCaGKMMSLGXL92ca2sHPvLMjxluAY4Zq2mege2UCHOuDAzD
GxV9lCIXc596sYtszZ1221BAo5zbpOAcEsohEP1z2iY3KTYLXqqY0lVGbAK43+bB
zLoQaRmFRSlV1YtkPAQw/JG8ee4G6AOs09PaTskSBQBM9CV+PfgQaQVEMrWK9dok
023n2EzTMkDoEubRWz5lvnfQuRCrfenTdNtk/2tcAz4rpnnSBl+VnPzKxiwELkYi
vjJ9BR7EGVAOdPy1ocnPJkWGP6JrI+l4K/rm4tcJGoYmNPaFbTe6f2hLUv3DkE3Y
4+5MZ3pbaCKFM3fDiLgWKbd+cwa78a0LmbPCOA2FZ8ejmTfSMwG/3g3q6VIlDBZm
fL5o29VUcPAIDgG31CW1jgDf1PrNb5B58fBuD+WoLKsF+4Fgb97tz1aGI3NNvGTl
DP3+j4o9aXQGhxY3QrLB8mBIxwQUvGWpqI5IwONspuvSySVVJuRUxhBuov7fUSKr
70ktLLw0NLGS2aDq757kmQV2eEH4ukXbBZ6NvKC/Rnj8J9qn3DBmOB6pwQaQkrNq
LSZ21GinH3p1f7dztAczav1G5Yf2RVYBwCEkump+LAzhalazOrrHXmWWBA7lM0yG
7iIX2R2pEd1jcsuM62X6AXLNqLBuq0+aYMJ58btOA7BwcQKPB2QfDXn8QRQk1bac
5xjesmbVVVKQalQw0NJYbiQVfY1opLejv45Kd6caBcYXMUXLAGMv+Mc7G2BsZdSz
icySZwoYd1ceMPav5rd47O73pHnv7DihKWmkP1UKut3wmoPoxEyAhky7ppYBI10C
vpWlmhVWuXLIdJW6MsPY7mX564O9EQpibM9CCoaXXF3UsfPsPwLTTvULa2ceulkJ
5OAQsLco2ZkO2+oG3YslT+RD928rO/Bcx8Kq6rogzREbYq9CdXdS56yL8efmq3RX
DNKbqJeJl1RcgFFlim4bCQwX7ULrM7W3AVJWkp7G402UJUO6lIXQHl74wL4Q/SsS
FV1H0tcrBMiMDVtjPOPd4SRenb7Ph4krIYAcqY3lO350JZxv+r/qrmIyS5HFUsLl
hN3ecRTMnoioqtDX9LSjmgpVNPN+1c5+LkHkCXHvF9Qo1E2ALhFhdgXQxNYlMnXc
rW7C6RXIrhLt2r79/8X227kLij2LSrOQttcbtgC1BvlvDWQH+Ycu0zpFHObTpIz+
a4Cn5R1c2H5zq36iDS1S66NUIxVTPLDZn8HlNtWxLhuKOs2PKPkMraNpkO+IHgh0
iWAmI1PfwYC37Q6hh3+c5XIEeW/vvKS07aYPpKGFkGzbbeLLS2+p7qsxAoFhB7j5
gahavKUxrq8iVQIT9Ob47uNNMG8lf7D+GI3DnJRYjXntGWCXpjbKuK6mtKjen9dR
qHcr6GXDxbbZ2hdJh0GxORqks13qsg3kg95+DNy7oBWj4fO113MJDWXv9m8kOQod
kjyaALzQx3BQSVb/m8NQEJ+1Vye4s61g1GwQcrzzwsbXe7DLl0BSUY/ROF3/BCxF
g5xyUvU2Yw2fTA72lFE5XBA1jJrCdEBClyAWU1fbAUrkpK7sGb/6Po9FAtoHKRWl
RCvtRfxXCjNIvcrpJ2AfsRjN47yUErz7gGRJBb19bxYBYf84TWZ2ZN+orQ5YIRNS
YgUqtNiGXASQ4U4l/2xszSQcxfRhyXt6Go6BNQlrMN65uX1h6dPMzFaynJMQfclH
RyXjJwqPhObl1mtlw6ptnF3XZsBffO5zQZ6hzSPFVcBLzkwYzES25loKpkyhFbpM
iJShopLZZq0MDXYKjfCsLPV4kqhC1krjikm3nqG2hx5dj8bMOAeQVo+bZjq5qHI6
6VOe+BglweoD9qNvQh6loIFx8CejzPwYJeFKq5gGHoS7+9iBySGU5j6yAQEGYwn1
/ydi60uxaPSZbRDZ0g35lJdqHUjjx/z8g11r/biKXQPD8RU7XFj10rKibKIZAAYV
FWcvKHw0nAYDclp5N8bCSxwfLjM+dbvOZZp3/1lUBlXQ/zRlv+bN0AJQgrQ4xt1J
yr5gMJGA2f1dbYpLm850UoKUy9SB+gfBFmV6E8SXyti9xFpqpOsPa5qQXW223mAg
TV2He0mY3FBChXAQtnRQ+gFCqOrkimMJZjZ8f5cqWI87rbUDj0+AzsdoKPJnVdd0
pk6n1pQ0dO6CXBD55GQVDIT0g24+1Rp7/s6Mk+Vv4+wMleA6L5cPvSHMt/BhvNKP
PHaVomI2Dsx7pE8DwYhbDPMc8qpu14loTwP7Svm8gchhr6FFxa+sZSL4JDrJL7Yn
0QLOVBw6Q5Q63q5g62SGqhoo9WAWLqPOg5FYFyuONOnmWdp/NikKHQQD1s/ETM9h
gRf5q+X/GjD0bK/nwj3I3+IZJ0i5LnelvzXHFs+EkypsUlpf78dRldYI7Kek7h7r
TS8hVPpcLS4q/r9aVQzfZcD5tC2lMU/J2erzXeFPMRv67YSYpyL0uSBFELK2+uJw
Hhmr47qi3ZEwjQbQ5LKaNCZaKDB/Z4WRlSys9ZcGoN6tkiULSyKcQfDHtyoOtS9e
FA8CvT7Mm1dNeXJu7OE0Kn584IENa5SP2FRfom97vBFDuY6If7XvBrtjxwTqrng0
T7Do4q801qy6n032FBnLf7qAlIpghl6vLbMeHFac9zar4+XQVU7USbfDPTyDSCsr
aHfFbHc7e0/8ur8DC8cqda7aS3JQFhXBW4xScfgicZHgl+Wete0vnRfNCKTsm1NP
DbrTgI0wmoUDcOI3DQHNCgYoLMQLBE7zKwcjnoP38cxZJtAhr80Uk0uPh/6ynSls
oKPbJjTfNzzVMfWRnNkB+m3IvfqCA/vHuBJZ5BQBBHCtBZaVVAX7PJxTz+7k2CYY
W6gACNZToQUdzaizHv5BlzYuVssRyuJEX99OFexnZfPlvC0mI6TswlbIISLSdHzw
yOGA3DU0hfx9bFtnNke5PuGsQkk0mIeMQDA2ZSe3H0FJB/fjBDLRtSjZAdwiEBbl
UA4g4sB6pK8/n0mpMERz944TvVi9p9Ccx9X2m+RRmcgrl3IdP5EKoOvstLwWkcQp
25r7SELoVZSxmOWGEYyo/etz60sJT9llPjaXDOgLACP7a4RXb2lJNM204MB8TxrF
ix0AKDCKmLG+dfzHbDziEa5Qs6c6+aGH+UsQIaV1yVTk38Gyg7UTL+Nl8hn73x5L
3q9g03s3tFLmsk012f4wXXyBwDpQIljHoL9sXrugxvtluYWxG3mudyrn1XFmj2Hd
Ak+hQyQpgi71RZmBRklhiK0kddXEMVlWJ7fflyU7xYzHe6aEY0RRDjyFW6uCuaM9
ltYfLGo+DVwhLBRmvacgZyKILcCHsjhFSiRScCV34h2nvF61z4+kHk3vGwSbG9Ix
ZKXMjlbmICAM5mjhS79l3wwzU9hZw1U1f+r1eRVkfAy7tvzpVti69ryEeYr8ehEo
qgiqQq5PR7HYXiWDWOIzyNoy0pLSX8g5pRHKbM0PjEq7LtRNpXnlLGLBkIZdi6QV
ZdV71ISQMdrNzJvtUhJShkq873iwnHPJ+8J/Ze9JAvqB64G4cM+ULl2Y6I+3Pfke
TkfiXIdMhgN7/pF6fcKLB10bwdDTK8yQm92KGvOzUZmTmXt2StRsurk+nrq65oHP
YNt9XPtU0PDAgIBgl5F9yAfrlsO1AtFLtKUDRA5q96oVrQisACdAv4Xznu4yLqQU
em0v2B+mSjV0yU1QQjERmctOIzzGhq/KZlI0Tc2IAJQ0cRUmSRGvaD+Yz+HmLHJ1
t+arIVAobKEJI8cLpaHae5QEdEkyEBv2bNVdFNptm3B/3dXzDt6hp7Szq3BZOMOe
YNXotWn13ZNRemoxyTUmKL3lNUaB+2eoy60dKPXhk8XuPfmQlC5tc9aFYYDefCSG
gsFmeG9fHTE/PwW8Wg5RuEv8eTzwcT/sK/clrhoRZwcp9IcxiGwah7n273nzLARl
5ccy/hkDV6DyU037SNRk+NfvxtKk3JqENUmzgK03qL+N4R/e11v1Ob/xOElDiUC6
Wb7d48iEgM8USP6rYoGcWxTaimmN9D2GpX/pY/AgWqHspo1UdcUlykWvoSeUU7eY
gXPTfJqanVxsyx+dEF9kcG25ZJREDpuL5hAAuCSJtLHluzyuTQloCGwq4Ju5dc59
CX6lWXONAPflK7qT8Y2Kfc5k7G/dAzKlox/TrdktezM2rNg9iDFPfk5LGHPihjaP
ggq22fS4/92XMZ7CanzPCy35A4nAnlFkR78QgcAwxt3Znhm6ahDg0xPvNCfihPbI
e2p7rbasprYk+iLesQPXI9a2C86FIImfWHj3ShAKRErDuxcB1KRHtnO6VlyCDt2a
ysqzOtLq3Ps2f374OeDuhU/lzcPiu/YnGyr16tjn5/4MC7p51Qr1U7uBM2UKSilG
hBXlp1jnbmW2AHm4/x0KOxTes7VCzRD3ZD3zzNBt+4BXxHz1Q1BRZl8s+xKLoxmN
Ykst+rj2YxaC2zMaye0eYnqXY1AYKiKUIpLa+O9shkGrvXuLQK4MbVQJW6McI65k
OYSXuGmB/hewUmi1U4GcYswNeTBiJqT3Nz2V2RokT2c15dhoxwIMGcBYqRJ5iy++
7RvMe+DnhvopUySauJgpzdVpffiOQjAJMwljTjDVLaiCVeBapxrO4lvh1j+7GDp0
u1YF2hC7cTcNrIoqFfslj3mHDRRFJg7G6T6vWKkNc6/azW32Yekzvj/pNjYgpzyt
gVK9wBta9EkcMy2EWZc+PFDcJ85iZtrgN5WfyoCkPSvKqHpyLw4iPwM1c9ON59uS
zUmwYzIx617mu2hWbexe+q1jIfmZGHpqqijrsYCXl/QcRKJrq+iX2cW/PgA4DYqT
0MBW+kbz1T3HSY3Wnp36j9kIEIzZYZKaZoHKOLS9Xr2L5/eAdPISpxy436X6ZyID
ml4J8zb7g0MQmuVi48qydLHT0QvYbbNR6qccLYB2HKI1TQYNXE+4WGhTlM9AV7FF
ENX5JBxrpXoYH0MivNZNKZTObamxpQ9devJVKZ2639luiXjMWAir3eKWWfXyG2v1
8K4mSzWuQyupBH5E8jgLxZvgTrsH1WU6pZJZ2wo1KLKGCTrPNYf7E/MNCBIixrLt
ChbdfoR0gATMrTu2omDM9xoX+2r+JnceDmmKUb003M6GU4ZMEFzmuzb0hjER0bQp
cRzMK1LwNcJVyg4OBJ3MHdXJeEFLMA9UHFnU97UkzensjScIYEhFDB1Je4N7GEj4
oBdCBRAoDcDPwtSdgImY51ajt5ePE0geBwTcitlXXSbmA6oQUHu/XgTn4EVkXo+9
1ByjiSvHUEi9tZUQ/h3tCoqw6OqJFhxeGerdVPbndZuZppg83PZpb6HGnfav7j4c
wEtKmihBy4uI/hB/ynI5FoSbUkjywqko0wJHVAHnY8u7xTlarpWuIIJnX2bEPZJO
W7sRM1BtLJPzm8eGQSm6JMLyQmmonJNnxBwiBZ3GamkrHBDddtL78s6vIgQeKVHN
l3vL2NXOYfGBi3Bu7sgCiWMyj+1vMA/Cvwcfxmkc57ihIz0XVe78mxoZKLRquqgx
T2WstSRYLGiYIAvqqNX7zai0SdauqPXFt67RdgI477LRLuaboXBmot1EUTa3Z1jS
jiHgoEupwM5aNqFBMK+G+RM7ODoW+Id95qDfFaQKpU+D469r8ba7VpxTh3Yeilc4
QOgNxf1HhhmHNAPdXHv6+UR+upCQr0KrglGMIkJ4YzPAQwdezNtTRUlFVPp1OwHY
zLeOAboLqBOlQW3JG4XWkss11ZSKWLIsqXwdF9P+wsTfJSWUdXUtz9igQ+slLhFE
8cS7Hl+N3856LfY4EwLwGy0Yf04HItwWH6sLRed+1HklisVU7wP6YfbWGEiafT/C
sO9Rf7b7iD4+2r2iKe3sgCnJhBRJ2PTKcrbbANYJl83EikwriJ5yCMULGss1W5LP
YdJlfebQLu5W0ePO7g2Jtu/wrKhCJdjkVDZoIDta55gqPbWnwKOiPnVzz1tl3Cyd
GNWmh38guRUOLnHRRGjVTCF52qjVEh3uszawuzCFoG7PFMHG9UjP1k70wOr38f7+
fpxlwIC3GWtV+GT89cD34xA+/HpxPcSHDNOgLOcgwlaO0vnATNCzc2tW3ibyO6e9
9NjVqY6Bkej1ky2Ri4r1uEnhiOx5uCZ6l7y/FkeGBd/QxUFcFm489NtKJN0hNumz
ITxOrciOFKxxlHoIOHly11sUxkX9ITsK4G+PJyej51zK6oD3OwmAQ0Xva20vbw/P
HXtW42Em7L9wG4kywC2/Nj8NnYXfbTnhOvcJ4BggXF7IWRk5mkpdmKoduqgQ8DD1
5tDhwLgjoy0ivf4BO/xf9Iv7mxG/JsQW8q9IZ3iDOBVz1svSneWdbYnaYykmIvvo
5Qg6A5bK32XDah46oLuoXiFVBnd9uDv72//R6GyIr2JwAXyOtumrr90twUvly1mY
7dMJWeiYMgH2b9Ka8KMArr6nU2VEaF0lKKroq8BV33mm55y0Ghdy4MvgJU2AidRp
EGNNDupcGUYK1OZm31HZ0NgBOR+u7DrGmPaACZsSGKaY77IAMLSjU6lnnKkaV/2g
6N8Mvb2BKuhgSE64uKjfief4NDlhC1901FCFNxUVfpgFG0AzIuT/UuuX9GLNWXuJ
jvxQkklM5bvEwwHil4QIzmDxw9D6VD3eIY2uXaA5EdVrhcS6yuDWZAo/5cXcmL3C
VLIJMc3L748LXzGqPk6R2RckQ53aD2vokVDzCItAf1DTMT8tktLeHZHZWzFrscUN
k7joXJYjvBCOxerc5w9j6Ic6PCEMbkS+b3LX13PUQDexIG/xnmPHhZVIO1eiO6G5
501s6snVxIo5rmtWYNqhVYJR1Hh6lCLN263XPC+MU+BhuhSMcUAFHi9Jpl+8W+tj
TwytodkBXiqKIj1D3hYi8wPn3yu2qZF4VyuGilsO58Rib89LvyunxxNnmv5iBr2Q
ghP1u5Bd0HCuxPc+deg1az3UWd7Ty/TxAG59dqc4fLFpksXp5qhxZgjI2S5hcyy+
io/LOd4wkceEodWyj1d7KgTnOemw7+dvXLWnSdl8wsenJB/fem+ir+cJH4Rpi2jx
3K8w5b4H38Gl+qrOCPQ2Qs8be9GuAfji4VtYY5h8X9NBeVuMLs9Gk1hZRSPwprq/
zEr8JyIxid9tMnJn8s9s66Gd2oaxp9opmA9fIMZLeSSvZ+8BnY49UE0SZlNmEnmi
B9bEboD3v8I8mghqAW/q0cYPJGGgfq8541hZDyJphwWWSlRiVYJCXqPFSaI7LIXl
RVYfI+79HPeTuCOlg8hcQtSJcHISDN6R8EKUh306GYJ5YVRlNDDD/GEz5CcU0q14
QYHJES4tWKhBFmUPQp8KfjMEsHSh7dFmhXXJama+v8xPvP5yI9KyRCxEiO9ygFQg
Mv/Ea8mlMrDlTprQ71YOmj6/wg4lmVqpIc5+TNmGTFo8InckXo/4spxvvz4dHNwq
IA74rnWKLXZTD4J8y9C0Wn6NaMeGc4njamq+wfk8H4BlUIz/s6+NjgxXA1GHulJp
EiXhIyRMbja6XixeTyMxi5LzP/HkGDJu9ekztklkRzfvneQOl4htMGOluQvDHtmO
JeNUenY2Cup7Qp5ZojN4G/gKpSZSDH2crfnk/3XIvrtW1mVgs16xyfSjjX1hx+SH
I4UUew4JoHiGfGOawh1PG5lp8dUxXUF6G3vwDHmtN2ZqKvA/3ThsKmBEQ1VolknB
4kt29KX00L81tYeAhjCv603KLlh7FyQr44lIeQQ4ju/cF/O+ayLBXDYG5Wpvz5w2
bSzYI5LlP0lq6g/0yXWdFaLqdbtZ700xse5nfNpVvEAbVJi91tR5t+a9vgjn282N
mtqgMqk8l2WM+D7oR85EAYbPFPwhYlvM0KIcpMdp87dKgZmvrrlj+AbqalrwpPkU
1fzvqFbW5/Aj0UHRdTT9sAORvOIIY/UchKinqY1Ix27+Ky3AEFP2Yxt28HitbBlp
lLHCcB2jOEZRtY4niVmn/vvkWB9vkAjZmVwS5VDlnhZKwakqyWFXhnGZxCtrabjI
ogEk6cfeTrvhnUHkc5DEQvjmjPKveDuOHFqm3kZPxOinziFoUUayp+g3USM5Blyp
JrTh/+2BpV8QolkFrdolgpSiOc3ojTd599Lt5SjnRXRDBPhYcjDatyNGhlZ9ZrCY
//GK/txoTN0bSdLwTCvJYe4IT+qhzANm9ld6syjchhbotBCmfBqoQLeUIa2aDd0a
yStj2pyX5MkfFYLeqJy18ejou+fEex9I+lJDjhPmDAADNpdTGwm1ROzX889JHpF7
HGsJoP9skWw49Xmt4tUK0dHxrEOOinEEpF0k+Z87bXmGpmQDl0PBZPtfFww3Beuh
N3qsK22yomonyOhwHBbdozmDinDk5W4Ghd/V4u9K8hSorVu34o2csgT2+O3WjFw5
6/n7DX9fSSjtht46wXRk2ZkHhsIBrmKQJ35XXWhUEsO7DxHEGydRakqnlZUnO5DL
6iHg0XlNccJruEuH5DuRlRgGkgx5wUTty2/sW7WHJfNZ21dTw+GZ59mCYVjq6BmS
iVdvP4bCPkFmMUIZCN9g8Cft41q7Gjc5AN+qGnnUFbM4viW0LZ9lNZVXq7Vg7nzb
+YvYfMppF9XzUxmOooisqSoi1CMgy1f83LOKpyrvjLvIEgqSU2UG7v+KI72ZBqox
7Ahk9te1lY4R95rDT/qQ/FX+QMHNWD1BL4WNFdkQZzvwKUiBx1xgcMr11Yv6NPxW
TosOHBximQlaVVSjDPRqGi5bCSNwhaB2hULMoPGFafkFasR0GwYUdni64lMdqKxi
ed7XbYjZpL4osFdyh62MZAO1KFed8622xOzvPgtApzsPo4ZfCGRyMyIqH/v8sBKo
uYFYHA7FZizWyOXMRtf2y15b7YilUCsPzaskk7hrLGoQrj3x/xOPD1R5X0ecSVc6
TdfJxk2QTFBlqeiXuClsb6Qd+pWB91yTgbzTHPDxmrAIB1NAPNfNmZqo/6WLCXXW
5k3O8RrWeeTGebISEFLHXEEQsJqkM/xFZz7RRhizTwAPQtc3ehAT1PTh6Ega0q5N
2Ay2n784Pj6jR6OFUB4czw/Q3d/ch8W7+Do4kVoKDc12simVAJ7yDdhMtGZt02jh
6s7cbLBtEUk4P/SI4W5iTNTyMuTuios11vRe/5XdaAJqUplMznLQWhVAxTzQmPGD
Gto7KBbLYRm+dy2OpxCPIRX8tcQKURnteqMUqU1lr8kWqsF+5Eml7PuIdi2gbuAF
EFUk5UFfLgiHx+ZUK4f8YdUEHWJ15e3oLrpuUgTD7QlBEtWSmbmmuhwNU8ARslDe
yLYoaU6QK8X17fiKGj1bfJeyFnoa+ZKtBqNdSMq0V3UOENt2TEDJD8iCPyvJy/nU
ORxTRRYU2tTe4EUy5AtRtX6196PhspuYCBHtet0I34jungC5ndWaet8HE3qEjtHV
3Z64iVFPSd9Q2PXGE6aLEiQu5yCDRUqfQBWICq9WKhuqh1DhZPww48MM1imE5FSZ
TigbWkF6RU6MLqG6dp/FTpLnHWb9L7NVQJeB2Er4jB0JCCVQJN+XS8jpt+x24tCf
qsMb3e2J84URiM9ZwmKLf16iHtJGyPe7TjmRBFlQXURdNkC4fE7sqGJM2pJCvXbp
1m4fHXfXIKv1V2JS5syZl9X7qHOSsSHX/B+nPb6XnFNTAFliPq7vzIAqwAc9Qvlq
Zwei5i4BPwpmU3xMuF9kmdamXcCSx2JgHwIA4X3Yv6WiGz+kv01SaZzuD3DTxpip
eFzbR+usqgFNa/rN2tH14yLqbkSlHoknur+XD1UOWWSF31w/ulOP7LHNXEn5rJE6
dGHiat08+f6NKOgfh+Qf1137I7zZEFGQsK5/mdMy+EKWeq5r62XEFoaHBL0u7Yag
RzkLvdTivoN814e/G8PvTPjWyJUSp23U4HOcB3MTaAiOmr7sa2BJDzPldidImGS+
CWRXoKoM4Ked/mQwHHTz+mmfHXCvRUeOBZVHdDCPzvaODGJ5wEJwjyp5y2g1DUNW
+gZIYuRprT5dwuNUId5gtMzfPcT9Y+6OBAQBuBp68njUYA1ukV1Wnbe69zNEwoSG
461/RJ1jDYOXNRRjcDvUxd6cqaVcy5jXFBIZI1+mtmF93D9OHD7RKWiznX/igjL0
R176dcEi9J6eE1rBQHd5YCX2ihOsjBe5CznWlrETQMj/fKqK4JKHH+/uL57uHO8D
qwhuIcFZgb3NrWWYMPLI7R8pTmpLd1Y7ZLfeGPHrY0v5BsxDYUIXp0Bnr3RnJvp9
flAESR+fr3eTzVmu9QMK1QAXQCY87sFu8eh6h9YqYFnZtwAD4NNLITnmGePYOzVL
xlqxLTZTsh+diflPQvKDzEHNjDqDNgad5gsTUxG7qDQfvpXd/PHKs0BaBZpvNxMN
dB6h/DEx5V2ZUBokSroNltsaNnpS2DqJWYgzBROZFSjvZ8GMdJ+Qm5RTDHqzaaJQ
owQRVmHjaF4/kc5cUXRRHHOCync+lFUaYc+279WX6QNpUpdpmvPKLFbMnW5ALOUz
k5iqEsG6mdjJEHeo1SkbxUKKbSgHhjdlo478DKVV/95X3gwlj1Rc4M/Ao+YesVS2
xYJfodSs5koii+IWKbLcQ5dWMDjACdR3xurmAfZ0lJcOPGltbUF6DaTis9ICwwJM
xWA1KIQWuB+In4XKBO7ukbqN63uUjWjXufsHNYOO3gXzCjBMKDVlpCcXd5WfW0D7
ORGF4lfk9g7d9skF+kSHq5fvkikxMCd9St/UDiP0gZ7EcAWa9jmmf7GSAPEBOnAJ
AX14ujzRMRLa99PS3csz7pCcI8oKl/MOcnS6mr9IN4HBGs6jSSTVTx7Yf++3js1O
JnJxDUVGY5TVNY9YObT0sL8x4UVTqjN1w3uAiImn+qKMcISClD9+1FHGXOKZCyNF
gVZXFh9PyvFTB7aL4GYHX7VYXV8FWYggidSy+pHKuTz659mhZzmkyEyfjNyQJuZG
yQplr9MmVZe5fAGqRXJaPC8uGTe8maJFTFb1Nj+h5wGJvObXHNx77rNzHrU5/LgZ
M9LSuYcVTYxKhvIm7b4iKlz39XW6wBb4dE052kEyZXJUZ2coD21whZ7mW3Ct/CGU
VxfJGGNpQwusbq0dxWwMEWwIHMR+opXhBUBa4ErZozcF4NsSt0iUzz0POhDAW2Wf
i4PLoi0pRxr5D0wwoPelbqlSSCRGchh4DX3poziX7SqNwC3qa3a96aJ7iY8sAYIx
IndoWXLj78bg07FaXtN8/G2J8ktJNBrqK4HmU8I2UO5wtyYDTfxqkxwd6OiRJOxA
wFrfa4XDkwG2YSGqtAXdvcUVz9d3L1+ui4IariuHO1PChBoUPbC+aJDbtocJaFWh
EbyTZ9mhc+WJYvLBcx4HUePL3K3zTL3fHY+nsAKUcoIEgs73ogQKjZIPJdH9w6CC
N4d66pTnWzlqcACUADfU8no7WHy9PVPekvWVaE1paFsG22qravZxTruFsQ/HRjDZ
Fw5DiTlT38lqDRkZcp3nX2Tgx8Pbclc17MJB3D3Nv4MJ4WfeDLyvCRmQo0YqroLB
ECxy3L9oVNi+ckmsJb1OTlwfoIeYgOrvKuMriN1chN8nlCUsCn0G/AHXXgsDc5p8
vRt4XXgl7ML8jgoQi8CKugHI1PDL4eqzxneQMyx4R+rwoTK6niW+iMAvntILjYdN
AlMYh7nkt/7DOk9codDu54mGexAp1ibcDe0BO8GCnjdoSprw7UiKMAX0Go0/eaqU
ENNd48f3fVol6r2FHGOn5UP120IngJnMlvnBcuTZCm9y1ptU/cmjCPKZdQ573oA0
Y76Az0jBdD+nDEOAggzjJjIHByPZr7+jR6LN319u3k4XAk3/O+v76Bkhkf6jXZ/4
jE5xLHYED/23UUpOlOBRWpsvmt2+3fdo3G/q+NYg++jtUuPg7YyDk1cqq9ixwkwB
R2z/w+/hfxQtzH6Sd7g+6fJZnNKlAtAMEs1HGOfJEYYBznWtpqc2QshOrvNEtR0Q
KdJ3j9ssRRARRdm3YZ5dzQSPzySY90PfE9U7w/Y8MHIGyHa7xpmNKvs1TAFjq/yE
QCgdfhXZaH5GmkMAW9gXfma8dnW7xyuYZ/Mkm2rie5nJ3nu73epcqzth/TzgxmTd
yPQ2jMbKGRSCYakwkA537qtptpGkJXUjclpdkn1Mzc2fiaV5ew5s6VwGySAiyRzw
9tpdZ1wNLtsHhGy3coertYMZ2O1pvaPkMibE7ERRwVyUGsPRSBECucDeWSmmoFgH
bNJp2mf1jNaIb3SVLOtcYg+17Shjo78RCUFdGLE6lqPPJJ/PRT25p3bMuLDEsn4L
eUwbKO+Z7u7wq3sV6l2p4nrc1zKlXT4O/KVL3eZExhKPZe+m2JPIIF4Hu56KYF7e
LEFTQv4flXqbAjsYpfTFCPu334EmW+sglOhYJaULQK9tF2dtorA3vRHCLI3vnsnj
24m1GoykjQvYt+VUhCPF37+xou5Te9++s95U6phTmlQ1I6jogKP8Zam7H4TFUWXa
5uWbVBNBu8/2UvOzNslC3WclgMMVycaf1SkY8IIqan2rB07omigs4UK83/p2mUtZ
8tB+qlChbOcsTlRvaukyWjeaOLnNonk9EDF0umlib/iygbQ3c/uigMFvyHEmQMK7
iMiGtO0t9TujF1BzlGyjI1tUKM7OPBxvEiSU1tIrF+VOc3BMVsk6ViUJU8G4qqBx
lkcwi/w05otyLfEmXf3rDqs/Ly5fs+jHImq7+L3QFT8Otj7bCcj53i30LO7NFRkW
aICFwdaY4mw6jl8lHEpQi5f30zSSl1i9yOY4Q+enEUt6+51tfF7pY1q6mNR5bA0o
cXRKqzFVjSLDnqX4ShHpxrKTjG1GhEgOlx2Y7SDdCDbddtgCWd2PFXXdd619O0Mi
ZjUMAyx1uhqzJn2zj87GAvz9HuWDfJZbv9KOUnYjqLMHe567qHZxhohoGC9hP4uj
o+MQ8x3x+XpCKRGOGI8TBSgY3jCHKE15bqEFrrFk/da7Acxq29RiIT9FqSqOLIEY
RlpQKW4zSy/AW3g63AqfOeWBw4wmZsCb96CaALWDhncZarnPp2U8Z9pEhLR2g8UH
/M3rY9Xe1ZeXK/3jByYg1AdXuqIZx4xp+ffNAbKybAuIOsAxKknd7vbh+UymKZ0P
C9Q3xt344UiGD8jnTm3gTdPR5TvfoNsx6V+4fYf5N1OBqXlkITbou1RWdUKBDsCs
mbifescHbwqlwmiPkiMDBJXK7Qo+l34lOkBJWGDQNAHAPorD3TPbyO2vBp4Afq3C
HmLeM3MKB7gEnsR6Mgl+i2mP4H88Y0IvFzOshUMDcaL0/jwuTBDH2o78C4Kr2b18
oYuXWYcY/FwQs4VBtxgMfrA5V3zRFCgFsSNeZIhj0nylfXfzcSM0a2F0UfaIb+i8
r6KhJnL81Qro2NoLjDfIq11jsFUMoW5DQifpejRfK8VFsof5hCFXdb0kyiEJVl59
CEoX4WuoOSGjAJtSulfZVWLRKNa2DB1A5CjMXMdlh4uphjWKq2wQDFEMI6gSxtBR
icsEBM+Ie/mCDlN+F2YjfJ+jzia0peFq/DqD3zYEdBlm/e8ZsjfstexXBaBPBqUn
6PG5pNUBVqoB5iGTsm4Tt3iELIz0e1+SNKxevZ7W8DVQtWsdmtA3+2kq7w8hPif6
XtJq9/FsRuT74zGHGqzcngBZX26f+enSQ/gBuMjtBDzmNS5M0ZIjY232ORyBvQA8
KGHhUA9GzP11+X2Ptz3U44CDwSWOZ/9szzxb2UARFwsb8WjzLNlUf0EltlLnuHj1
+wIaBDg8mpXcFzASQNXxCew33Q2jtYoelD5c9kA4qCNLaDQkBwRRswc2IWGruppK
xisrno9OCp2ETkZ/wCC6+c2iP/nhOQxyolS8NYJZtDpG3uScK6tjVcmHYt3QbPsE
ZnimLO8E+pqsSXfZvofIFKlR8Y5y9DWCvuwKItzQKHvzO3lgY62KQtM3Xr2HQJA7
KR479qX/m1hNgx6gShwyXElMebv4Sg2+lO1qPjeDQR1w/LKMJL/z/gj4jkeFp5yT
RbXwU5/CB8p9xTRLE3MVcq/qlmCtxgS/YwRtupE9nkc57kp3t49/Q9k8XGc2m/bt
gzw35YeOB7hopEksTFlYRLtvvYTC6RCqrjX0bHkU6LFUJ2V9tUiU5+i3Bl5IA626
MhsNEUaugaZiXSOqw79pnShOFx4pYRzxptzJrsFBLnNrlCd9T+ruM4HBqmRN9EJG
/yeoQOUjRvS8qM7Y2LmmuUp9qgVOl9Lel+AzPYFrdrfH+M4mUNKLJVp66jUxCOke
nD/AjtTRWlxvGzhMJ2oHfaBBaSt8x8D/sqgcvXEHkxLhQ6EPKw4iXoYNMiiSwXdg
81M8KL1gIvx74lqwaCibRAYrTf2McZEj8QtXI5tigeIA8v+eHU2rZL3hq0uUYwJs
oi/T5rKEo7xgNqJBFhwAAyFEVEo1R39s6/T7z8dck8FBpMd4yJ7RY/wEJwOTKoWo
d3IPcjsl9qmWW40xGcXOy8n2FEWoGGlOD0uwOdbAmcrgNGYULdlhRfI1HaYzoccZ
k1CvG+soPXuPrNDHl9C0YL1Ra69Dix8BebMdlXND0utkPDPUksJM0zrKsevlNi4t
ogFOIY8mmEfil8iZwJB8D3MjX4+HIrQ5N2/uL4UeFw1NQ9LfwNAd9m/ZAz6vh8Id
4QMfgmFo76IhUo+RWSclFK6yLJTG1r8WwByLaWrwQ3uQ6yZr+MebxvcsKiYZ3ehu
5hkBaHgximsGNFn2o1PjxFikR9uu0xU5+yz2GLwGSp4W3aZXCazpvcqbFYzfJZp6
amrrwMF/DSIOQx6lww+2cylsNMh2mIhHxl+Dw/1dChy6yd7dVwfXU8yNH3me1LrX
CJeTXb5QiB/FeX87xW+KIToFYSH/nIY70h1+hwQPGBZUDxGV6cqUYqHO9dzfDXaN
3vjX0lVinCVz6UgyWt3MoIYJK9ayKMY9r2C9Y+ECJ8UHSeuvZKeQJnuNg6bUhL60
U5b+Plp6qCLDhPW9y+IbghOnrpXEj6/qMf19WcyQaZ/wRmMjKdGTF1ggiD1BkTid
47HHlS9CiJGLTFF0/qb9wTc0BJO14+DvAfAKV8l7T4oRto2mICTzw0yPbwHxe/3i
XP5yKJmvlrAwrUo/LHgprlE5jYMKp/iXVV353UL7OxxHLZrh63m8eDvhl9pZOBO+
/12BLj5JrdEFYSfpFY+ugaGzIDm6Nijy6JU6AFLeZr/j4a0fyCoNoqWt85vawmkj
THZWAeZKQ/o2oPQUJk+ZGuzr58dKy8/lxGe3SzD0EtAIi9sjAJAxldEJsw++7fAb
vHKmZkSBW60dt4IBXmzZspwxlwR8JhL2RWvmvGFN3Kym880zjDK2F8wUeIJyPlEa
MoSReIRnPXJ08+30DpSoKgF0a8+xm/Q0m66OKKbF5BY+hoePjxViZP4KjtfLyX90
V2madjUatM//cGyOvyxJapZ7QYFu3ZOOdgu1xHcK1TwdYA07Lv/DMFqiqC7qAXD3
elGFVltivT0vMgW/fwCxq/zWlqOVzfvRKjBVmK9XmbTYuzdHWKjy66Jo5hra1P3B
6Qr5xxyAJnba/yF3cJzQOpEci02i1lvRCOOF05Ax7PiSr/EddZ68I3xqAFlHAvSl
DryZQsOPJXUBSwxH2pSuapJxGsYp9jGOL20zJH9qNcm9x7O0BXqkzkx1UD985Tyf
S8s0aaHOcoIgJfe/kCugjoXJnRscOcHmRO2Arj83+XFuF+UT4aeY6yK+cZXhU4MX
6MUUq9cIVmMzmxmnVhxEIBfeKwQGMKtLrwFythsmcPdo5C8/ApJypEAFbGRDcsyo
ohsV3NhthAlsezR9XNG2fE0EEnFqGzAVsWMVZssxf+6hZ/VUt3pzRyr/x2s0rwgF
VkLVz/QbZwKoSe1QTDFseDvS8lm8oKzkUhr7wz8oUlhJvlawHlGZmCN/9o6sphNJ
ZB82tO7b95fVLpPrNl0inTXq9u0U2AYJnEB1M7S69cjcq3kOkt/JztEsVZAWvOc7
YeuP9PGTpMEoer2XTMR1w3IVIJAM3iDBoxdI1q1MEio/uFkT1qzbNvSsErNhf2GB
i3koWR9E+NiAAACJssyymD7gRvG79TZ4g2pIHT6ltEt3sLbvn1EVLG5WlFaSizbV
gUO7C8ffNIr/ScDkjt6IzkewSpW1ROla1JCQwxHL7cqrd4sobzlc6Sxt7olwl1pi
kyIHcMDjwATWeQn+CC+lbZGgckay6DjuGKKB1dzoLgCmNylL8qXaWQf2CkKmCqd/
/xyQy6ZwCynuLZoRCR++/88GNaWIceDkZ+jQ0sMxCLEN7+pAOq8P3TCnO4StaJ9E
TbiYwzzdAuiK6ABC2RNSzubtex7eCv4Al6in/km96J09ewusjGVuOrM1By7rKVJR
/cQt7utHkuaqp0pxTG68D7ljVkcUgi8wWn9xpLrgoLVfkB5A1L5GmvDPFcLMiVq2
XbENQbM9f18girivCbvFfxVf6OMcR+A7hG2K20CWeRQtjAc1aTI+73rIRzciDNol
ghxN0CEPuagDPI2Woadze2QSpbG8/Hgp8nkzgOFuGK7OZGJNuh138ufxLkLZcJ6n
F0UpaCn4cYtoYakB2spooGsafWcob/zqjengwph/3mllC7IATro1c4YO9cIdVXU/
obVG9A6w3AIGej9sqllbdR/ZTy3euVRNqdy4v1HlGmGSl/uzAxSoK/U/aR39UeTI
omIHdM8TUOrZOQZe3GN1aTNxRUTSUPyLwK2sSshm8cBmZAQjjnaadExuBUEixrrC
nQjbAKZX0sYaLf7iu3lrbO2CiwhTHpB1D3T1473mYyyx65vI6gohJky+BKlzYfHB
bAc/Ght4JMMnpB8pCYRAVJ9VQZUDy1JWUlub7Mo1VQjssynK9n2MFQZoinW3XbmG
/3CPE7G6JTA/fM2bv96BJYEzYf2Bb317llRI4blzNFYwgF+OYdq3Lp2c0g4njf+s
4jRGhAKEgjy79g1NuNV8UG7P1b2cKMry8BhsIFd+H4MCe10caah3nMwYFsih/PTx
Imc+oTVmLyCjsqce5G3kQhuzw8ZHVTBKwWCBois59riqzarSYrlF8htTz271fC5b
AUeTFCwz6YlpegIgKpnrUYPjdDb61AKEGTLRHvpbyf5bON4j8cVoCf41ck4lzzus
Nft37mzwff1HMaJmdnT7IJjD4r2CMz0qJXGLa3HCxxwbbuBWhrKbHAT8uZjzaexq
TqkcSCKvAHNL4tZUn/r9PbOKXxnwZ2UhMkI+5p6hb8Wb7eA/Cbi9D3WgP9vqb84x
vTTdsSuJgwcrtrNVFdCqQ7XVTQtN9AfHHspG679o0uqHi2ZPYD1eRxLqdfWCfb4Q
ksDdoJafl0J8lG28x8f8CbB/SfbmPC6IF9C+KnEyA0dDaakrfoNaALs4YV1mkPJh
1LZGPNjI7zMp8coDdPXy1bGi5pTRZ3MskY0GDlas76QGbJJujd/c7swOj2euLh3F
ItnSKWc/mrCFr6e3/wvBHbeJaeM0kGSuR8pjH4yzYUOPkfqAOF2m/X440GcZ6601
NY391GdjZulAcm6nigsvJ8H4AJJchV3d9nj6YAHWHskPE/WFbCPSk2rxL2C/E/vy
o90AdYL+Hj74i5SprCk6joXeKAzdxFbQKhHvJ+/NgjgE4Qbc6BHTq68VBd0vpV0a
BHU0O8Qrg/Dwcxw8U4yCvn/LSP3RQymOxSQMDmaUGweXd1kqLxtr2d8YOLDXz93P
78Q3M6c94xMPmcigmyudgZNN887LlCvv2ULi+RLtGyJiM5p59+t676SqCDCFhOpl
F2L7sV8+b9VoK1A6Xp+0m3RPX6PToA2aru0YxnOg+O5xFHjrr0yEQE6+8yXvtxW+
P1nNwU0Xd8d5yf8uvmb57U5W3CoNxFDTxDi8h56n2VQgqXPDlF48tuksS8Gm4yss
gA3gt79ecFfLs1tTIHJxFUHwYiP8CZPv/BogzU8zJcgCOJWqfmhGRT0WDjviyEB4
OTiSCRjKzKJqhyDehmDOisQ0OR1e6HhnKyc1gQOZq251OdkO/2K+D8h1sKo0VDw6
fy4n7jpooV+wi7WVXGTL0dZcUw368DxUof6gL0VhZatoqt06oUUputqtgD4/fZW8
YLR6fY0yKNeIebttgsnsV4qBlviZWHPS5vvePnMnAlS/m3NW2NzFeKTqidpgiCzr
WQnR5r61EUyOLwjrPcN3nNQlLCqjv5aWfaXqMDvtK0K2XbnLZkNCq0JrwZfjzKb7
ZhAFbNw3t1MdIae3aAV4oKRladfJ2CobJbz3r1E3IuXk62jJcciAVVJ7OSXlAdLZ
mGPtiuHE3Mz0WxremlYATnB4JBFvZ5UonSAFIbFbXTlkVAN5pd6CZjE3kZNVABnY
rMszc9UboB93Ga0MUm3PaRlocIWv8CaBH2gOPxKBtgi/tubQV/eT4qhdU3MA2ngT
WlKSO+u0n3aeqEGHC3UGze+5HxtYCW7FQGJp/h7UKFP4ziKrKwMjwuVGUXJIM1qJ
nQjKgz8xfTYClYjtzk+d7OmYZHzx6Ek6PIQek+ad1V+GIOE9WjG3Q6ypqedoXDvL
VVoTqpwKvyLHQmgTARUto/+LA/dBtQMQwjHUznDDr+NWp4+b7x39z04QyXas9NwJ
5mngqqKrgGxlxoB/rP+/qdyak6BUJWaaPBE4FYtGMFR8tAl4UUh1HkmNchl85WBw
lFxLpdHKIw1vsiLc27yIzdZBZg51Ur82BVH9HWN+GJ/F+7ZJpgYtT/zIi9Z3bcmX
ubcw1X/Ds35PsTkjMm8kiZIOZZLZRvuct07nOY1j1wrI+ZcALsiFWiZkbG+/D+v1
peJSWNh5wgztnUPUvMjwPnT9ONkVbL6dOEZr6Mx926fTqUljPt4SaffSvTkMDuCQ
3K1UADFB9hGluYDBUuONcs8KeOG++atcHcDKBHA82rmPPr0kFnXpU+Xmo/K5SsmF
nydnKJNrRPT/YytdLBpb+iGPpzP9JsnJ9hlOD1kmJH6+uM1SJS4l1saYQ1rRZ2i6
d0sUIMTksGYR5qQ3crq3zKjtpFdBQwd4cVpUYLUiU4k4hFyzXYgmGCWezMYdcpxV
ctJLWhIMmYY1LvLsLBP9zFFm4g7uxVQb2htm/x7BHfok6WHJuBRYPjM3znHUlurj
GbwsN3dedUGECJDMPulFFeHfqoaNO9ytkUoHjWSy01G9GY8W8mDKappEjqglguHG
XwA8GXjLSvVAdnU1r8JhHj0jdqrztKE4jLx1l7TfZPterQx1DgzR0XBHIO6gsHsT
LAXJcGdT/s35F41h+5nAQHr30Z/qaCvO8G2oJ0gOiUg+hSua1oXK6YTYBpgVWYAK
n7oeQGNdqQPlU2TMnBgvWM+vp1quhPAFQSyj2kZmcMNs1lHg0xRUKAeqrDlXeo3W
Hk18YliBMf95MQWn6OwsxF8x/gGCqCqQ+2fhoKZ2J+b6FhcRxunGh0ygN/vg4YgR
sIupjt2ZcFeyPlNSqv6xfHeU3TbnF8u9wS2vgQikZBnWIdZApEl6/pHO6dOy8oce
wF6V5y3PUzOj2nOeXN4CTMwHqms0OaJ6CufAYASUUclYniDtlN7W8YBLcy0oDHO9
b2tYAkG2lgsF7qkTN3LJJI6e9vKMxYqveSqlJd/ttv+FxzdGalxOuVl5E6O3eQ6X
MNlVC7vyoyguLlhmBIqcoHp4ACx9AWnDFCDenahF9cn0MCj1dM387XInmKveOYzr
Fopa9TdtvfkI5BOTmFMCnCGTbPovkBam4WLo+nIGisSdzIooIfwa6trVqDQ0hpxm
l+UCyoEzQ814MFih6Ayxsp6ADwsz6//Lhv7mKUDpjS3YWlZn6FtHs7eprzbmHeDn
6e7A2Nslp+V7bURKZejfSYc8meM/oly5Mg0lX4B/pJ2vhiqo3NgZkhiZECNf8Ujm
dawOQ10N5XXUfcpBGFMT9fpZeXrTK8G8dIf/HlLQkVbU2JjuQH0OFzowOQN+IuIh
RvP7HsRFQb/0GtIqYEegWGzjTYwogQNNlS70Gj0ou6ldE9M/XKdLkCBGeQ/sgkZE
JFwqxJWSh1HwVyiYQTIxREjM7IfPWxG1qDzR3iIuySAVrNqTssseLds6rC84WNdh
3xdYbIPPDYEvJZIFvfzeEswLFQMy9g7ETEQ+uT3zn1qsfmpQNK3n86f/btFxim82
mXCjdxc8bb2yclINi/0jVoAQA6783PuJvjZoEtKtypgFXSnmFzXpOtn3gfUg3hpq
hWD9TIL9cqHRDRaHqPRSQMDX/xqll0O5t8rkGCERiSKJl2092fDOcIT42shEFxi7
8g7yAAMBwuVzgoRAsIyae2yuoRpQRGsCNV4iOfJnGg3d9yiQLZz0oCgXxwffDG9D
5craWpzWIrYlu0ky6zQcnlaH0bVw/DYvNu/TlL1gskUujmIxpAXungfrOaNdQq45
zfvSC629r+xwi4oVRpI6eKfDe8/0zkUJLRQoZXyhLZdk/Lq12v+KIQVV2HrEJvQZ
w+60ofUlgry8jh86wNxTA1NrpqyfXqhYixJbW+W9zO5RUmXQRloocq/yAOrYrLdw
R4two5zUUPrQg6u5daqtL5BbMOqUipw7manajPrPT2Br98P9+4OEALD1PTL1ufPe
9GY9IFma9HktAQgTroUxsq3WIDinPGghu8mayn6jngVopTbph1Tl1YDQ+YKk+RqI
H1ywLjCgtPkjUqhhSZrsZ4t7Fdq9YGXhg3ZCFpY94Na0UFG2UVDuuzXV+SiqH0Y/
unHXBRcRVXx9ySUo2Nso5tPQ6/DP5M9YEyhfSVXjyCnrbjYKO+xxQYO3FV20i20y
hKnsePMnDZyjUXSGOfIm98Q0eWFHwuVOHbN175/OWcBz6izNGYpoSabdrZlyN/WW
PrC2HLIFWbYbnNzr/gNMwsPLZicBTLUd8oo+2SXsme5rVrfCm0ADiHjcU+AehtJF
kdhuWrYDKIj9aA4RwvdSDGZkkqCft2f0sKLBZ0t4uVMi21DihIVlsGPYdrOtu2Gl
JpMBvRhC7AX/1i+DqpIPg9U2Zs7r11ViD91cV/y4rIxID4Mq2C+ShvQZs/9h7Sjm
kBBk7nWxCs9uBBeR1wMRB0Ge3p983uKgPF8HGdwZzeiZ1AZJKFIzsVrfSgGsCLfm
LgIR6Y8s+0X+xTW8nY/542Kr9XKYVth6QrNZ3qzsL5hxz4+8bb+rgJST7oJA/TXB
NSHGktiTkrQwy+3rZQUb2ug4wHqdxOTuROj7pMFaH5nvO9ZzBMYajnyOIuLEnpBT
0mvglAZLypvGWRUhkPKtJGVDMnRHULYJXO+Wf6Z2110QNp31w83I1Hu4x5ge1D5A
0MMu2gu/4J0/YM0E2ErcyTRcrDd3Wd0DlxUpxufWDbMFyf21I5rtsGRDMVoA5mzQ
ANYydk2LyO/rL3I7gxvM7JgP3yf2aV5pslgNpw5eT31j1uw2fQNBVAgmC+WlIJos
QTins2YnEiKx3I0TfIwb+BCh+EM22iVokKNkuIhwu8GHtaS3OK1HfjGPO+TOaZSd
Qz1RM1uJWvzkDVkWvpiBbM3F6BhRunFc/HkyI2AcIacgdbddAXuSer3OFGNHV2k3
DMIEyADRbcQRDFDMFGqELn4sKKtfvvx2pt6pDXk8XSnQpUpy1GoTKiU4lg/7Y9Dr
GPxU/B8B5NwQ0c9HOkygiHDJ+MZiWwQIjzHCO4CjnTQdpj+AAPGpe0ACED9qldAJ
V1YHyO8yGVdOQTyIXFwwFLKFqt9Jx8A2QRT8fjzQspKUmQwdd7ZznE15URhXOKWA
TvqutfICiXbB8j+bR7lyc+k1P5XIiihi8x9tQl86AKpIil4gzMtDBuwa2Z0WSD+D
4TF1Jn+w0iNAiCmf47PEHlnUc7ew4HPAgwzvYZLt5pP9LZlu5vDETLkHYjKOnS4X
OgStgnhqQ1LesioFElmEmalESj5RQY5wNi5vV0j51Mor0TeudbgF4GDhjQ4iLtRZ
CRrsuJXvwTHtz9hqToHrrHTqv2bPRoaFTPuOAEC18MgWk08p53wZDBjOuOXwsPuN
f/qG4iUPy/pLArymJMF5GYzzpzPU77CZ6H00+IB2A6lcEwjRh5TEa22C8M27Fu7R
NUg6HVVZelJ8bBAIjq+Iifh1FOCR5UfY/VTd2KAMGqwa8txjBwbyuFkGJb3AfIsA
+5oCEZcxI89iPpmJqShfA4jg12fUory6Fpe/hW+rX1FqKxTGS63O3hz/KKQmhinw
toefI8O/ITFi/+/ekX6XPEhFXAXzM6AWCHRF0Jiu3sb4DqVWuUWzwh2iwopoixId
+nZ3b2zTVsQEM8heyMamLm9swAVPGoOs9MKKlBx5o7atDMsdow+Ds9Stjgn0r2kS
4Vr4l3WtWxy4WMx3+w416wPzXhueETlpHOowOFh/X+pNFCFMHnZfSIbSrepCD9Lz
6dJv9Iw82bwx7wCD8y9hFC4wUYqbz3ldGr6Lk5qfItHj1vY8zN3xDMxRvXGzYopJ
+qHlOsPz5WeKDJdi8GIKdC4N4gYSNInYl836jN+LYTk8ckwCI5J228gy6YGCqWFm
ZedYhpzwgGm95hVWcOCkKrNPd6CdOh2ekn3zB/R857cryvLMXwEt2S2pl1aEafXF
XMliTCEnH0VJ0n3HXHMzkuF4/6Nm9AdW3MUQCmPVEijd2eNF0rEdDzIx5qyQB/k5
4DDRJkC8sZ3Fyu0dS4ULrUNJFLrk1mJFIPVT8C41p/Z653xDUopEiHc2XKXTpxzN
ZHShy5fXQTxOjfWIZv2oi8DkPrxrjVeAsgLjjjqCsZsgXEfZy2uoiJy11r1+EeAr
yzWtrnX21l8yMiyWrc86XGd+LJ/ctevW4TaiyGWfZqFSJRoI82q+yHJGwudqHPuc
Sk03Xbh50krw79SvYxYdm2hHSlcs4JhMNAFZ7E47FewoIsOgIi4UqpUDyW2oFGK4
5uiLcGnIqbCEWpvVVyBXM2VLbI9psUbk30FQImJ032KtJBIOjFupSQGz9vUBaLu1
mR/T+uR9XKoAvmEfmNyaIuoJKE8jZ8gxp0T6/DGx2fK+lpHsWp32yw3h1/IyBkIL
vDTzE+UjZUvd1WQbHDVdgxVJmt9zcnj8dP3so/RaEcMMTiNdxgKix/uY3PA1XqPe
x1gyL7wPoXdfOt5TcATa/RwXoDi0XlC6b1GQifXlpNzAQmMWQBNdW8Ja3XDuyTVn
D1DmPCC6NtFcI92YN7ZCat+G3V0336N1e1SOs/oOH1TvTclHtZm9zPjsvY8PQIFU
7XanTr5tfFGhkWuUgPmFUXuMdvDyYLAmR3eU62Iry5SMV+d9luxOO8OKH5QeClie
ptQX8hftPYt3OQ+tvDfDomkRIx+o1Yl7wQJ/A0nvcVnrC28lfNjXWm/ShMVKwvrc
scFmLg7hcFzdwTVZmL9HEUE1IiKE/c8VCA5FgxUuEoiirpp7Mb1z57wRV6Huk3Kv
Ze184nG4wH+CkrOSaCZNaeWvOiMJ1Jid2JI46fyg0MwmSP90ao0B4CwuOrn5uGXA
Pbsp0fIwPdL+/rA3mEb+Y41riG7Xr2vB/mIA2Yterym0chnQ+dPxWIHxPC/W8yow
CXTNVR8XzYjAxBzxqr0zTyF3z+ulO9J/8IJFX8a7fpHv9wz5Xtwmfjh48TNfwMPn
jzWal6eWFAZiPWB5GuYBFGKk66K9q8YEkeaHKXJ+tMgtcCCdbf0IxN4iv+yFPw3y
Y04XK/pKbDY+kEr1c0ADANHZkb3uWiLeYOOI7gI1PSOWh5KOtWuFkp8Ot5D8S+sx
0+dIxmwNt5HwUatU/ZH1IRexFemso94DsbeKsZj0QMvnf0u7pyW4EWgsbB12SXvY
h8cDQxTHcO9B9AgmcKWgwO7k0BQJYlVM5M3FaWl0Ye/VF7epgqthfhTre+oyldwW
DaCfrfOPBkpSCGY+qtrHDl9lhdDe8Vp2A3xnHfTQw3xJFCDvtClmpDSH0ERx7xgx
NXqbFzipGdRdkHK01SgLK8yW6vMOiNmP5doEZpKJ9GuT1fk8L2CoeDhyd42/9Mb2
bK1qY9j9+UIbIcKVG0w2XI2hM2gQPkiRvihcPoQzB2YpGTnn/4lTR0vUDylSiRnV
3CzMU4R9WW8nxKND5el14qH+9vNkbNXTBnswnNOp2fp6XEgvTHtTn9dl+dAymfJ3
lkn6k13UISTg+RbNfvDuLlyPbZ9iQ9EUX5uS273KUbF7iCzDXNoQ6b8nreygamWb
0heIb5hFCY5FmKdbS/CJ9GaUXAjdiQfiWjF0taTRvbC8NlIIovNiwHUW3PX+vFpl
9I2r0klsRMcNmi5pZM76Y5JwFhjMfCnojg9jDG1MkkrDHdmtgs1VmaMO4Axl+aep
18Lfp1mB1lNzRzm1DkNeHOs2wibVWrIZh5aG/Pzaq1RZIwfw7ryzCXAuF+Uzt4Bs
+b7sAXOWyF+WGGaQi3h5RZ6dXvzV2xB8G595cTiiKDq2FWd8kP4IhrejrQ/oOnOM
dH8SUeIdUY6DUHusxr9qahex3B6p3nju1SdZooUKVe0jVuX6LxlRqx5mkkCdhIu2
jnPb/2YL11RnPWMii69UkMo5VRxuc6+zEebzgpywzg8FXBHpVmDYEu96gVqbKsAi
1wC8df9S3U7EkY1+59yHTMmGea6EiRP9v2bKv5f+cMiMghgw0SYLhOniCPnMTwKE
Y+g8Oan97HlJ+zhA2qWgasbY3w6yttgt46KFu55msQkTrxYDAHhIMfDUj/mxXo4h
BCxHpHLxKHmkKFzEtfwCxPgLPHQNLNfPl7CU1OI29WTU9/crNqMILSChcz/Zbd90
Dm4KzvGs41N5JvxSmnadcK4+XM1I0a1cMTdQmhAdY8ZeyJ/tE39mXp2bf6LLt6KO
BPFsuo35qMevNrAlpbptnyYOfQ4tYf2ZAj69Tyors0I5rgrhW1P1edaXDBjNkS1Z
NpByxrdDQe5OQSqiQcdUKrE7uf9plIpdLfxJhizyL2yaXsjAqde0ZclVJyT6gavk
niMnXa1tqw4Yvnz1hZY15nwX+jxtcnDE/AcejDY2+DSyGs92HTzWxp7UzYOlu0h7
fhlF0IJXTNuGShCOgSLyBGYkZmKu417p4lqMH+nq64VxZXaasQQb7tMQCTxUUcuZ
FhZs4JLOqWXAfzl6UJqOhWlTM5P6N21tUXxSRBDBd312lOwVOokNM07m0OOLuLTq
Vk+OGFFIC/Uybq6c8RjzHYvGkzyDavctEgSoAZs2GqIhuTO7efBdrSdc7dBRv9rG
+/0puvKOz/d1pQRiuIbfKfymCPIRuJP7XC1/J0FP7ABPX1baqbDQJ7sS7XT+2ioc
EvaK1bDvIJDhgFkmO8vmzmqpWLs1AelAvRxpqDg/uy9fyjKVtvnm1C6WSy3GZz5h
P5KvPqO2GeMNNG68opQlhk2sIcmdPtttPybMknqUJUJZ/Jc1mAGSvpZsbvQUY3or
jxrFupvD8DAxve9gFGAs536vHckTsyRfJfQfVRgpc+qsl/IlG7YJqMNiOW/g30Go
Lp9hGELbKNpUW5OgoR2fID/3hNiCPZ1erFyoSV/0myHjHM8a4nvh3QDqzWJVk2Lk
NNjAxJekvDCy3kqXLE6aVxwSWQg+qzSd+Yutv6Fi2R/xkEcc7Qr5Xgvd5gOZuqZ9
JskDfTnw22Y2t2bGZUyN/zNi1nvm3+irxotdISbBfYTmL0KpdO0dg4K0IylKRpIV
HNxNzW/2oD3XOgpEKFtDd7eTOcVi7o2pGG3AoprnuCmVEY04PDbMqaUuTd/GQHhP
ivaIcqlvx90B0I2yxr6REA293sblP5L0txsF9a0UR8YAk9QIHtcCsYwKcSIHUyrG
VkMV1jyUAxUAwy+AMtjN2ZqPve2q/CPUKqUKwlCIkkIlHGL6xcSvqhuyN+FNrKki
QUq6q1bVrA4xtJ8jhrCxkobg2XBNG7P6XOStjb85/bSxYep/1XxjipE5nmqzLHgc
KXCaDcEFO4dh03bmZRa3ozTPwUanEHukWcipRImdejVEn5quULwYI8lIMc2KvORL
5pf1EMWMaAblYXOL0WWK/JRWiTVa3U4s9CsmR9y36OMrpwtuuq4ef8qBdiHY5BWf
lw2+8C7jNh5DZNowljenJxr4MvJleoOa1PRr/4sf4/hIuMs1K7eggq4S3kZevZSp
JOwjvb2/BYkypyHghAT43qCBDEY6SOJaBZZrQ7kBgPCcsDNB1aCIWDEBpP0wyUEW
WQQv4TdyAEMrHRbxNmAQ5lGSvGNu2/2yCeJCmQkT2apj57kUsv3Ldpofzqhu8zU6
sn1JDu3YtcatXPa7A3beKNaKdkudkz4eVNO12F7JMP4yZ22BGsk8U5LhC+YEVW06
EsWYWdkVga+r5AYiu3OsBDG+OOk/pDUHzr1oxhqXSmwCTVhVjCdJzSUeRlPLHOgS
JpNeR0BCJKAmBpy1hJL0DL3eF3jecJx1xoEVYPnywcyMpIgJYwYNFgHVCCMHmA7z
sx9QFhYihN5dsHFDIBhZT8M7skyogUvYXkOsBM73edioqK/KO7pbXn4FryAHFZwN
lSgsuJly/9L4vASo1g7EyepbZa5Q62lG77RTm4tcZkvQAesXDpnViege2OycTCO9
7URC6MDi+JM9fSRlXWpIJ2RY1jQqbcCrL/1TEq2LOmXuNgE9JDCf61fZdqbtsMon
1/aPuDaSA/OAiNpdnOLOLM1O06yeIC0LJ7o/auLMBWhUDa8tpYm3uvN+8EczM8tr
5KrfASAzRj4ZphJiXBtJcuYHKm+QoyZkryM1oZqa6IW0JMXc5Ip91hf6QnvOUaxg
ViAzLhQV+MI2+e4ngEog6P6ZzBVjOg02iFuWbpAeWZUJTaKo2IilHaZrAJNCPNYx
klfgNlzZKSZ7fEP28PwfF6xbcx/KepEyX8cme0gyhtglKIIX613P2uS49+bAPl0e
vu9PcEvU7sZR5WBd1vlVXS+njYp36S1EeWpp43zfM9jrkNl34b9hEFUJrCLuW5J+
FHwhK82c9EQzeJKGmYVgdQmCX9dcFEgRzxamkb80rlGhRVFWxfVtki1pjpJFOURv
T40T3nH/QX6jSjZyprEdfmJq1OUx0pGF+RDM4fNiJoqxr5Yj4uLq6fKs/6wC9ZjG
vNWnV9GMrCkFOOgYN5DgQpq0qi9BP6v4DXgQzjZYCpM8ptvql7/yolAfgjoxr5Ox
RSTW9Bkyfp+5r/1onyEeJ9dFgHSnqOTWS/BeKSpgruIZN1kEj70Svq/uIBTSySYC
nOF5MzD4Gf/5Aur9aF6KT8a37YmQEtmuP8c6jFkEnP9BcDHrzhU4007uSF2TjxB5
aPxYawLhx9DJBYtPbHbXxnm71mCUDo1ZXnql5pSWeTXnnzD9Qr8RmankL3kkzKd4
gibpcz2Ew1+zLD9Em4R1vyR3Kq9lcAqR2JA76u9mUSGRaq9AvS141/qw3uPV8dRi
8cOrMBtVzOhwxbFRYVtSjnq6r2g7yA+jJ2NBW91iieNtstv+loNmYidWsWZywld2
aUlvKVaZskO4ghR3qU+UtSU8tnWltQZ7t4Z0F8DQ74FHwBWoJkHyC0pmqxJ8YNs0
dEg9d6oEMQ0UEvGsiStqgX0CzK3MsJG/ahsQibDHU2K7tacmHyqnsMD7VOMawfNs
Jntkw0zitVLplE6dEtIbdntCnFtve5WbhqzLiWx6LW2pO8MV0npEYRd+JJ4/5rCE
Fe1OuuwWj4+PO/E+is41rxsr7XVTB2/cyxbyv7SQK88HeFqiayA3gRvqwI89DyjQ
ROpBdloCNAGRJiVoHzXFdxqaK4l4xoPGiedNIpk88X8rC4wqQhE0i+ruHt/Gkd4h
KcLJKEpV6W5JA/5MrvsWS1Bryl8R5XEB3r2tqJpr1qhGId1K2tDowjDkESbIBovE
zd4cs8/Q25IVgM1VCuhwAOGPOYG/D66vlN2SDjtPm6hO8ILgoUccYhIBSgH/KNoZ
au2PnkQAjLdWWS1JoEvyEnKJUmSF7eXeWBmmO31jcHjqj3gkxzpu0Wjr7eZwlUNc
nTjDRtqx2cvAFVAjJ9mtwXNUYkrk5DCax4KXaTzw8Lo8ATw3hhoOBQ9Fb2oZsTOv
RR1w4Q1c/Cl4LEKIuKGzX8aypczrslh1U1Uz0MF99HJnqPCpXFmZANPMYnCpev0r
lp5A7/ku55CFjcJckx5u+OMDRA/vBN7eiiumkGZuiFqK+/gEPX7oGqloIw2bjW1v
GhIoY8buaa/p936tMHIbxD9/DJ7jlwGRiSHqznUziWqDXIxfGCGcdWF1gvlCSmeg
JlttYMTB7BTAyC4L3ftbq8BUM6MbxcyPlmBxTjWf4SNXrYm2ruuyej49hogKojy9
LbSV/PleCen4QhIrg4tXUAXfdo2Eiw+P4BF174UhJjdytdIhmgA9IYqMfsTyIAp4
wdf61csZDagt+uKEc6NauGsAaSM0kWdYZtYOPdWKxNXv/EQrxXwz/YvnOIVzKzsd
Skq/gpsa+44GSKZvyP3rTDSr94EJODQhpkqc15PCMPHI860JwatHzXQ+OfZe3odl
T0o7BRju8HiGXTv+OABr5tRkYEuMYM+bUKN1TPTupZjoaMXGZ2ZvZZE+wDh0IjL6
7tt/XNA5miagfhISAGkTsNd9Cf7yk+nt0v+aoujQspE1t+GqGI7GbH4JYqQeUfFi
H4s1y7gInFlD3CtsGX2Q9bFH15AWrmWKsTvahry+FzAAuqyh5EU9HdKi6Ur0yVQa
fD2M0pqgmN4+r91vJSvzBdfqEt1geOk5kKNw7LwdLguruc+mD0uHjRzJVal5koZE
nR/YaopIj67ajB8jo9lter7HaVvuMfrV2zYvEJqvsCRA3uFWelYozgt2RvJXnPM8
8+dviHqP+CYfD8cbxF5NtKmngeaTWWnmS1NMN68zSWgalBBQ9Zzd7OXGyHHqRheV
eT9vD3x2QE3F+cXNn8V1aIc3wSlpgPjEZFG7cjxAwvjd+UkKNHiYBNJPLKis0/8f
qG+oayO5zPrxuZVz3InY2woYsSmUsyjUbashg7WWi8FKSkZF5Kw/MWlW7vJfb4Tp
y4WmTl+7lklJXm/Sx3T1QrVJsy+JSPdsZepLBQlMZUkovMZr3DsybRTPBK3fYiQq
CzAE87hcC3XE21zDIL4mxe/f9Z/snm/evLlY3mG2hP8K4Cl2pRGf2hz5TlKd5S9U
uTd0qD1Swvp5SGxL3yMCMljq3gN0rloVgOZVrpQAmKY+3fnNfl3OdV3JVwxAnjXj
6fhalzDSyNQlSYrCMT97pzeh5EVh3DTSWzxWyAa1LIU46IPHUUdDbXXQlwYPPQ0M
nvmlmVWpRllbQpPmAUTG/2VMSaSboO9tOh8TungdL/EXVYQ3dHfzMwH6PmnJc0us
4KBcyQVmQObWMWQL10fqvcpyPWwkXHrTCu2F1Iae8cBFcxl3heWr5poXNNDcSLD6
6EkxrlT+t0wUGqF/N7n3OSR11ACpzfz/hinvqnIol/J0ezyURDuAsWAQOSt0PF+A
ihgFWQPLKWbOuG1jS/d0tcahTuADFfQLGG8t+mBLZL6gAPRyN6ouD9kYjn9Z9e4d
DBUEtf9CPUxLZ8YIPerMve9fZyR2SmJxwdMLHgqo4apXFJ2sJA0hlczKPYqLfrYX
5iRViQgE9/cZUtfMZQ7JMdHnPv+eGryMmqnEsBF+tWyKRVJFPaFj5WBCkCPbRAwg
wcdtyCB1YAKeS8Dv2VIP3hov18/EMrQcSU0jKgCQcdJhBZzJ4rP1HyuPdei95A/S
+JXZI7MQt16gjt0u39pZayGKTXmhITN0AX9eGWs+PM38dD/eKLpWWMcpBzuDC6Ij
1vZ1U3Up1d3jGkWgJo/FMHXRDteMOVeMz1VRxlMV2ZsdWCCwql2Ig0iTb88qGAHV
tkVgF0YUdBcyRc6qcXl8TUBPU5dLJ426JhHEbV6M9YD0WoNN9V4f0YEAm3uCmiKk
K7GtbsngaP8K/ETnCZoL9FewxNsJTH80vM1DMlnkq3dmIyQCBY99PZQ7R/m+u5IT
VsM74GuBJEdHDcQaYBN3IXBpceX9waZ+as0VlENjdzgBjOurTFTjrOIp93Zh5EMh
f+r8pw+yxynBtySXhqsuJmur15gj995b/21l64Y3ZUHgLll3JJb8I9yI2UCCSlMc
hVg2+OrBFmk0RPZhwNHy20pbIkH8lB2HMxpESHmyNfXn2b+Wf0QGGJMOpUl5gXH+
uXhLlcDLJUdXTNDvua1atyLv99dNUB0j5Gka/bv5ZmugqLj8Wzhc9yeZlC+NihYm
9zRzzYCDfQf8gwb+EtDLD1UPBSCjGciIp5K1B95bUJ7LnpPDzdChqCWAOIjwsjTP
599+6Cvu04kgMPCn79GJwqWKWE4QjSDkLFMUgMlbjMXBp2+1QkcGH4kmQI13yPjx
a7Xqe8EJGTwrxVZpIoRlEZrTFDa69JlVwvl2xLhDgPwvOHwpaJhtA/RUyS3w4Bbc
Un54u6g2l1qaQ7qTdLxVmdTMucfMiME4gk21uQwlHdvYyUCq5VlxHvNyUbwZeBc3
LgeY3fVsaRvWpYr/6xpiYUYJSOOZYT1eIEFpAV9JLK9TqUVNKT9FYblnYcLioj5E
TQgC9wfPiFxfp3i3rIDCWZU7L9/InUhrXXaTka7A4u8nsziNh2bz6YLDx47gwtGj
GSgwJ3ERs0oJy577u7bwOwcxtZSJ+rmuSPlfTd7RYUUb9C/aROgIRQgp7mzt25YG
bymcTB1JCIyy6ZcOOHExSocMSw3OtKNl1RfnurRnPstEyxy0cy1uceJvAU0SnYIs
0/qOGb4GIoiqc6TTBTCnNKS+mxFc+TaCtoRwiUKMzWsDUVaacD64T8YpsspvIDZA
B89qS4ltUwmds6ALFUDy0mQxTu7MhKVKvwNkgbQ9733RMEdudAFvGcG0VR8t+f8c
MqcELvXhEPwJgaRJ8rJJu7+Eqd0PSESYOLoGS0PFVmebU6wLSb61M83CuezS2rbk
yfjjVLVgKplAXn3t2QSn+yyjld0mOqDkEQDLEpEHUA9vmRJ2tqV3+eAaOQRn5SGp
YfaqTJ1BhtSSjeMwcujxKvzFbtjSbcGRnek8Ja8uxYfjbSzthpk98REo94rkwMuC
fx2DXjd3RoBDcRnV4D9wo2Rj/vX1RQOpL+M1FElVleR1yPN84jzNTruG48aLb6+t
gCHw/ZqQ7HGBIx2lxH9GBQ/J6NMVNOzWnVkA1vSt30OQEJshBsBiNis4NUPNSDn7
jv+2Qk8nTsxEn4qcj/hZYb0odcc8wiVkMb9zpkntjeRx8ddPz1ciiaoQQDdML+3A
+ydDy45214E+JCXI7DQSF3ISNs9iOh4BiDpIa6XWfG3avdolZ7gSCSdXRZ7WVgqV
01euF6+o5VoP3Ry7jzZXxp5RRnx0ZvOrkLEDGNlBqgoNS7L6BuapUg5+lAGVYlBk
BSYQxItTH54Qswu0Xu6RY0wUxlbkRVhcwR/h7jqSVfPvD5Pl6quC9Tx6MXPQ1C8q
1djuVoeyRLQEzCWuRYM2EfsHoVoDRFDhy1DvM7vAMIRPN4lHNZ9Idrldc+OzxXJV
5YQahCKL96zUQyMgkWOGhcpkXk7nUcZf/qinUQtyDRs7Ycv0kT0B+Vw1l38alJfk
gSd9ttpEgyQlba+fMyoMiX/ul0gNhW24UkkId37hxBOh38mg4mcqwLgztFsckbNZ
NG94cV6IEM5IvWdgw7uPLJP/ahERuvPDhOCT/7nCpoi3fgte53yTrxco32MLV/sQ
nyqhJEH3uNZ1YfP9JJclUyOGMI+dLDyZDIzdBFkcWT0l5r31zmbI5cB1hZ4MuzVL
XfvSJWXyKr+Csz0By4+guf4CWnSQEAGC12gaAdwUKi3WAE7DDgX7oGCCezBMvH3b
aoCl84vXopJFeHxnvs/2n4MJMMxJKthO9VPoEv0MOhWtF4x/9Jax1FAK1AUMf0uI
s+/p2fy6RCsU112aqJPekLl6KYtpuNdRVQ5jRVJ1jfAAmBz+hgpALxh5YgdPmmU4
rVt96fXXEDH3786mtjf2sRIbD9LyKfwTzYJNoW93YCTKIEIzTHBSWPPDJBNgDgt6
/+ZLOC0sQS2ztUxSQ9G8cfYTUY8HXKBY2yEInNK5aza3/FPNEytwK/r9CPr0Ii2p
2qVNimK5eZGaygeGTeuzSJGn+tGS+Hd/49CIInox2E3KiAvw7sTOm9wGpAaoKbX+
sDUMbuWkAyy8nawTG8nW7zhRqWJkZu2UQm5Dtfa2XEXI8AY2Un9wv2xnnvD96qlj
QC6+TcJvKY0ZErMx1RA6/kdRisnrMeU4MDpLrat79PlAw27NbYWdTZrVV2fRQSBV
e3z1fa9pokQ6i4Q+NgP7fJn/cjMenFOCHotgQtPzdMs9IHfTbqhcygjxZ1r9UUfX
OXzMaJ4sEnDCWQKJ7D8YEfhdzHkmBniP6aM11FL3GodTRChYi3uVSewBTO9Ud+GO
iTccH3B9uQrqAWAWZX+/lx3ak9Z9PAP1DX0shltMZFyA7I75k6AMdyu2Qakuc+O9
r1ueGz7PP/J3coNIHhIBzEoadZF8msHvIOoTGURqCSukE3RO2XFvIJmR9rfqzUs0
YDk3OcD80LzyORlsfNrsGSJTnJ7q07b/E4dwI+Qd6luCLOBTy2ydGE5sltQqFfjS
Jw4H2VHqeMoieFZRVW/Piu11B5Az7CgDXKqXLlElqlEsh9ffCNtEN03nsoPAcgCV
Yy6XTKQnrHBWn6qoN4SFbjg552QPp/qyMdqnLhPi9S/DzdmEGC9ZwVqQJRnjKZtG
1gm/b3e9BAeLAL6AllmmQ7Q+k9xZDx8CZ9LXM72NVtj6VYm9LwlQm8Cg8lveJjse
F362KmAoE3GlUr1uYFXciN9uvJ6SqDC8aN97WQhziIQglpPH/ZQCX6fz8h+N04Fr
Db08vvmX9bhsitHc2AsIXHZ3TBpR6HJROuCM0+6mLYPuTA4UkMzbNTtALW2FXvPD
iEHK3+wmn5GtrMNfm5VD2gUbsRVXB9O2WmEkhPypKmjH+0bmVMC19HAXLPpufKf8
J8OyxXMxGfgV57jjI85ZQleyMEEmEBIzKymxvYM6ebYpFjk43nj9jBR6km97jmck
pXmDlCvUWzKfd4P43wszqq4AVmCiex2kV70sgiZ1noBgXPTbCAF3jqIo8qh51vEu
7vlYn2DgVm6hp6msP/uwSzHhz40bLYgGYx4amkI73hSIkP0uLgB5yVuC4tpYErLC
8CgYXTZAj88qPjNLyY1I6HDIzvbmn8Jr1L45znIAxLcJZIZt+ysnz16xs6PCAZIk
MBjyUxfPe2e3zk+AP0RXUotgl9iIxmZIOFeoQ6exwwao2vnPR8WlHQ6jMG2/W6uN
wJ5mZ9rKPtH+Un3GNSuVsVBHk7HeLrIZxL1eBZR9w4xqPuaafLY3fNLZvr4fkxtI
WqRp7vIn8Hz2ds6tk4NZNlroxvt1izxSl6D8hRXPAByyQa6PwNEUnoDvDuU7ig7n
26GZiG4ouo9itTLQ+t5alhYDgtvsjyeN9j0iJJKbRQeshGpVsAzcPBUufk04/Mau
WybzZYPtpOMBhoTTKC+m2XL1tgRB9U2sW3s349wVyAqfAnoUiHHcu5etBUrv8nnk
zvO1bHHTKvziGUWGmkxuscyJTwSDR3nciS1dlUAsbYPHanWKmA2XlDQS4SeuJf82
M2U1049sdiKDXtjfhWB5+TKRYfySgy7C84O7jHn9ME7ImUpMS8mMH09+IJ8KDC2y
WScdUXSCh35/2V+ru8exfQUKEQ0jIotgwq04f3d0690WIzLSdQ94qma59NPvBtFQ
+bIIgtlV1Uqyftz38GrLSAnZxMO2bO9MFfWeMwjtv/AqUNmyxUmVStOkWcFAoshD
LIGyC5nfKTEcaY1YYB2RmtzaFhQ4kvrzADvDn6CHGSgp/p89Fcxo5gm3iYv1Itjy
5GGn3B9qz3ko2t1Cbmbeh6HWUtxPLr0msOfvcqHj9pQb5CNk3aTvsGZXt0WTO9J1
tFo57QMnFEg+XLt7Svjg9Pv13he6DwOhz3A26fpay8qsIm2tVFTkGKnE0hW932Fl
nwzYDvKq7TFYWpXys58EtJjGdCjDRcDdicBHZmZBb3lx3v02Ww8aWRLUDtPExZpg
qVIxA/2R5rCjZaYfR4gSPDHIyqgaoOr1GG2+o+e+zMgNCPL3+a4CV3McPWkoctHJ
DVT/P/EoSGkmSaST6dHNVAzYhs9TgEM6kZ7jYk8+wS08RH96vrmLbKUkSw9DPCR8
njOR8FR+QbKwm4m+DlOrdfgVJuhaIMkVHNTFjh2ZKUD5Zxus7DP/IGKR8doH6GNV
R8IUQD45ACYa8bYtlFj+7WdGzZ/rhzj0K1es7lKANU6OgJ0b/fR/BTFQUnJ1Sknw
zb4A7nzV2xZ7B/M2/jLTJ/UwhMfwgQxLDkfAhWT507p7Qe38yK/vOGlmB/DzKrZV
Ipj9NPPRTEv5uX3OiEXdY4NyQohiOxyo7e5JqWlmQMEwuW+jW233+jIsibXyUbIy
iVjIG3RzwzvAIOjwyt5I1FWtiUsQ0dLw9D1yz+8Xq5250/QnVcuCSL/axvowjKNt
9eQUblZMAvVGp7+aem54xvcA4/ywv95dWe3WKAbbq1LgufZ1h3BcNLk4KtCMHut+
JG5J2mImy6ATpKkeCHTGX5WI/VUQ/WT1TtHQ60fcwS1EeNWz6eHd6XccJAKPKIhy
x5GYLPJ9TqtUvJWVAHNbu+L2wFU2ps9wgMZawdB4LESDoJC4P3BAXYZXaciDzg6i
mMbxaaiCMt6eDxpspcY1001eOdRdH/O/CVN6IsKa/fNPiygqRIB8VPUjpeG0qgXt
l75ne9RFC+IG21XJ43mYRJ0GCxHmve9HDB3Pe0EDk3E1befRVu0Mmr4l8192YXdv
nH9LPYMbNGVhXg5C62iS7ZTh96hFklXLBgZIzXVM8RviUitAbkUMw3ND9PzExX8w
dX+uzZtErLrjs2+jzMi/spv5f6fzwLEYh86/QELQ52XL14QoxxL4aokI6ood5f16
4qNJOtiZVkOwnb/G45Wu93LZ6hd2imLsboS8ETXDdTnkGKDV7VoDsjV5BAV7yGSm
sF3RxbS7qoy10k7BofdlycgoqldGT7rBdUQa9smim2HjqHvQ+Z8f1u94E7XqNNNo
ydS94KFGk+NJiZ2IBmhvfY3IkfJCmeV4uMRWZdRa27EQXK0Lv/r9EGPaOBMUpEhi
/C6tp760yavu28K+rTdPNAHhTcr3oqb1VGALzt8OFK4dIhCvPnGHR+Y7Dvf7JgPI
1V6I52mc/H7PyCNRiZN5Lda5RwI9Rytbtc2es8J2FJLlmKWc5xrGOZ1Xc0KA9Cus
xbA28aYwU3UFVgYUjFTj5sUDxvlGeQeFHbvSeuzFOEVConrkICwdLT/X+Mun9CjQ
eAFHBxG+rN+DVC3F0tsjjN1rcnS0nQ1qgb9c01/lxpau2ge5nIQrMR1Y3jstN7TE
QKCyYJO8/Y33ASIhz+8AcLmattqqnDcRQkA9stFFSP0/NlHN/ALXOt/IEGsB9QxP
LnK3hpB/dV6DkT//k/YJZyreSysSKpZMr6PDOKoS0e9O6mMTvurJaTlBAZxMJl2L
uyJfKx2/ZnjJlyn3criWFz97TNGWWCDdWOsUilM/I0fWsWH3JoOQrSjWvRzKjL4h
hVuW/x14+5LELlRdRlFr0Peu4SoOwW+jO8wG5LvEsxsWM5QOLi2JI+b3FldRzEs3
v5U/zGjPozWyjG6u6NwKYvZ7cg9uHBNDjmmwY8O8u7SelFUiPag66d5m2wihrqF5
A4IbFtgvj4VQCCBzXSlM/3AToVMWzaeJNBv5HfQduVluuOXHs7K86D0jT2f8neRi
DCcOfTaUi0YCHLhuaoErola6XAwAS+gfHVmhHQ0xCHcPdGEfFYTIxLUwLxaPlrDD
QIssuMC4OXN4KLTHQNK/j/FBsoEGWPVOuNdHbz0GZUSoQrZzvMg6TFceqtbMobpx
mmSJY27BAitZ6HsJLmYTV5k3Za+d2dMN0ouPW+8ID4V1Wy1pHRguOyt0T4ED0yMX
iV5wLgWMCnGyENmx2BpfA8E2KwG9+WgsAWLzXfIJup9nxBgl8PCMRo9QUSJ5gliT
oKyLSIEQvyXgO1SMHl1H0srpRHP7gUz9sdl9EOBr+qjNVOf+rTaC0HwIzXH+5AO0
iegGm0xur0Kp3T7bddzvKmROIOu0ANfbwxRJ9ghDC7S1F8U8ZMiezc7r/BLbeGS4
5c/X+x96RzKvCGlGHY85dkkHFxesQhClO0rhUNgeqtqeGgFBubYOAZeMKICXycJj
21KIHZtxFx/+TMI9bSD82F8RHJac2Ox+2P4YwBu4whRKZ3RaO234Hb+gJt2lT1am
IYTXQXtLryFMZexFVWFB4S64rfgL6LeDRa699lOpo06H6H0Xr8eNvXvm0jTw+26D
6+FXpC6Hv1vrSJtB2OItmLBDr1ttfAB4GTEvB8QpxpDR0h4tgyihBON0sKooTodq
iuuD+YbV4xZors3a2ABSHblwO35kfzq3z/hUQQb+fQ6MzbP5Eu7UXsP8QMdWI75U
W3Y9349cTIEkTLSFqH7VKa7F2raxQezW5KoxKHMukPa+4HhlEComTvN1ih7qfsZw
XlQUghXtLHGt6TbTmzfW6PXDaPqsr/J9wfu8NWwrP6uFxOH5qzSkVLMnlyuEw56J
F5gFkWJ12/lH4zBXU6mYVQzAqDK+c5ux1ZKBxa+ZE3T0QNfaq6rz55kxk5DnKH/M
zR65oX5E6HipXtUlXcpz3KPD6f3kXwM5NJQ+NAb5FqVbBUN8jFim0RNlJ6K67g1h
Yi8Goqi6VlV0Syb67JPdoMaH5UIbZeqvEadQfKwhxTAOc/4/rTsQVcagwZw2+2L8
9BpO08Yuy3qVf2QJnLyB+IVaps8+rxX1mT4oD9MHJgKy6RMDz2kvB0kzePtolW6J
oUOw41ccgFPcIFlGNtWS52WrS+EEtRKuskwNGu/xOsMz2ynvu6DxGtROMJXPTmr7
4npYsAS64TV7LooUQ2CcdZ57W/cxOj0xhL8o4sMUwd/wcjBN6CBextVmRLC3BT20
zz8c1slPgiteBsVX3gmp4O3KCWoEvqS5AFqh/Pbps2muSsHBzR5gsDKLRvBoqyq9
islzMRCV5MIyWvhcZb92vTW3A/KHG3h3LE+2TeqTS54DJeyDjKxRKjQSstqpInFJ
QY6tN2rmWt80AOJu7c7Zki7qqY1P236N94SGBobflFvuNCPe/fs7htJrvMLD24UM
gaiIFGSvx4GgrVBtGJdFlY9Tuf09ibETrM1MEqEy/Tnbj2JIyTxlMECfjDN4Y5d9
a6Q9PSf/bjFnwyDpcRfFKHYX8NRuZxaJ0pksPxob3ZBRCClerdHI9omEYdMK3wep
Y3onNSDD1pDV5b5Qb6Dz7s8/od41BaCuHoBr1D2Lp1unXwMGLLVVpfVe+9A6yAzT
WBJ3G4ShwRXpdhqYb1N1Ao6Ej903ZmO5Yw7fQkcnLk6t7YwatnUgoeBJEOmY6eFx
hixaPqV5/otm7/3HFjTPOQuYvYDhqKDYSm0SCc7b9q0RjiBCVKx1NO6EMkSLJuLK
CjEeWQ3/z9a/sq2tCWaeYPeIiU2P6UtIAt01T5tveh7uTmMtmrFE5PQyrPNefoce
XsaBDuwTQguWaQqd2zS7sqsornafqy8Bb/KSJhPvbKy0j+ZEyLHJVONa9kIhuSpM
JuTyHgYgsPVolm9shxcz5oN1M49w5q58yScZbVzqL1yYf8/Hz27/YXOvq7LsY5He
Y9eXwwKVAt0eot4staTFgRY4myhUkgxo7D+LTP30RBxBeN8tF8E+i2q37kz4LdHa
vXvLhzKOl1Uvq+bEgLxim/hkA1du3jhHBZ/0K/IebS5SYOZ658+Ns0hCnlFvitgn
z56wogafgqOx+HGihLeTLHZ6kuMIWbr3EUWyhhX9w2pSlvmbW9nMMkU0w3LzExt4
dSXc6XPDlED2P0jxY8brdpXdIMOZp8YSd7ppMDYq+eXQBQraFXayE8luLDFgF4+g
PonJrcL4gvPG6w5itfIdK/8At4TY8sEC3UgL/QLTbmqkdx+qWdT+ZvdbVdFAktI/
dg+kn4CEVkrCc5ahlMYkHVK/g/RtrRIzturUhMRpEDlyBng0fezoMP/Vp6u+q9tq
N5ugrlQwOFXRjMSsYjRPTJYg+yhmzkij5pXVSrdR8nqEB3HTj/grA/jWHj7xS/ay
5bQ2VRYqDl58z6lvpA9uiJMf/X95EYvLPuRhEZyVlBLIcveX7lyABPKuSNfQ2DN4
aYYcit0TcEtsH6u71G81M4WWQyyIpma458iMuCnzf79bveMg1I3/BkgWAFNOvHrT
gDen+c33hQaBQVrasdatE3WUch0U0/eao7GCeLGIT5/ih9krISvHLgJnCSmTsyaU
POBtUchbh0zDjuHj8sKcGWNcngxT7gs7HLLWDMwm95A9BC3+ZD1lG5pVSAWNTgxE
90kWYklCWGdVw7CrWGSZjcyiUoEx3g2tUFkrdgQV7EXxuf3ew9SXNmml5xkdc+Xd
m29BX34Qm6S+teuaOCoV4gRU0WuEwTMBJ8GtfHMJGhpRU8al0TYoTirvipB3N+pT
eKJOq9o/hRuvv+zwKShVygLfV9xvMMiGFLx9+5e7mUe8521lfUdu0kqCB8UEsCg4
w/USYL22USWMADzH+xUdOPsBqtlzANHoyy1lBkfqCyuslFNrwb3GWr0hglpFDkM6
QflM5CTm6vMvnX2nmvHOUSvGfq0tBOR+ah9VU+4eIFK+qSB2uNs+y95+GvEEc6ws
csFELWtF+IC9inxpd7zU4kdz6zc/9Bvv/wrWhj4LJ9LarAjm2FymXRsgba26iHe6
TL1D6Kd+yAoEwDFXKuXqzdW+u5f7l99wOF/Bqa8XT54DUVWjcuRjPahAhOoPRI2O
E5ppfL7uJMZTKQANjy5ZT5aiQbB3ROn0mldcOIzxtuer9dBCpOynsS6N2Ge/SJyY
eHAMEapY722XKLNHnRFBxyk+Nh8wpMQP2yiZQxtZ5+EyxTlvyXYGnbstczemBNV/
qqJTXLzPdfS41Q+JrdmD3jdlgoagv04NEXvvs8wTK5Zs77a6R9krY319F6fd1+5N
DpFNgdKvoy1UUcvz9hgVB6FCqJ87jsSLhhd8/qPSzI2fQhkZ0FVRrMXHRTsDDGnB
Aw4CkKbS8UjtGybmZhsRNcc10B+dKSnF4yliOImtDZZkLnHfgSjZWy9kDFOEd6Ak
N9Ri9fjLI6Wp5qWr5SABDicbpYzyqAxDFgPqLMt7dbIo45FUm2yehoM6uE+P8K7m
Bfgm9KIvaG4Q3WP2DBzQwi2vh7CDaz5+oNhaY8qZhpTZHCAsVyRxBvi4FGzHomxx
mR/LIJpCIKvXkVYoKWhTtqn9T/vQHdWPmp+NNGVSqfsNOEgsvF4qXzVf3jnltbtB
HneGhPUx1PLg0eB8Ed3D6BGBLT4GLaCnZlBKzAOYW/a3M91qpYFI85tjcM9X3jO+
5aTcucBWHqYqcjuLq70OWvx6Udr6IXsbBOXVUzJcSkD/4GHr6mZZKgmQjH9b73le
PiKzBvGl90IHnJI5dIPbBqzIrMumrnzKNwG2zHH6rAhCNvmoKaGhdRa7r+nu6Zvu
8zXDb5tN6E1Lhd6TwDB2M77StqEE7VrkNQEBX4/Kx1YteG1DtAXHQ9fOZqESt6C4
G4NNaST3jsjSiu1Sq+BFE935vqnCshUgfMpOHCKZXVyR+5jiH6eWON2lcIOg4+RH
bn0yBEE5OUHKt/Mp66QhnovCKpOGV0qBQmA5g+0Nrn46Oivy9tytuwt1ZnxP5bGE
qM+DaPq1M1F6rU5DtRlqYPzexsvjgbh7uN/PMlmY88xf+VPFfRT4KX0qLf4IT1eE
kFIYgHin/ynpyK3Cuwnlv0Pv4vkMdEpaRLvJ+dQVY1BehIwsRKqUpNVawATFquOn
/NKQu+CehBY/2JoWwqjZ8gGvoCX5jAYPbxTflmMaUHatZMCLXZSfNolgewPLc/YK
7Dfufq7muUVVvDIl5JePwC9G5rZ1QJjts/A30pgHDTQcrpMavyY9jf7d7kUMVNoL
QNCep5HhDlXz32Bf1bchzJCozv8lsm8d7ft/LbK7buaqlxmPHNAn39dE5wQRX9eS
DCHRYCNxwMboZJctW9LK3eVnUpSUV8a4lOm7kCea1aSlikUblq7nNz0gjVBs2/CL
i88pb3bcJLGZQV3CGcyhhPyk531ZQJF6P11OHOqnPY3rLh0vtcj/qwl2w0gZfUTy
H0YZT29o7c0W8aYJO9DpdhSDiR1StH14P/9Vkyf6mSouaMhaquDDQs1741VcgKc6
7ECbYAj4x94OrKsCtXSmHWC3XngPFhKvQYbiCyjtTKoRYaBv6UXBI8WupRw6NxBY
YJqO8Cb0WM5f1CYT5mf+C0rboYuMXJm4ZQaofnhIdLcD2Cxz25ZG7tzDAJ03NXPe
cF0m+GNvZ4Y78+XFwJMP0OsN2ULGvvkaNUvazHeBNw8aF6Nc+LHPWRcwxpVCD+Ar
d5ozqnCq7THVvzWAzTOVurdI6dQ+V2eMNAYy2Bmtteh4BDpHUr3EvNWzQvSxtRZh
0OL8B4qtg1VitTUdcsEiSyUCV2uBRe9fj0aBDrrTj4mSVe3DjByIfh90UcI1xHte
jI1JHcTeVBlSX8FEuGISQ/0A2XMsIy8xgAqXlh1evhRbono73Mi5tlIfhkElXtlH
DG8KHz8vJHXoUPuWXWOeplnu603nxIqvi1BRrKae5enrP9VcBNk5dbM67bRBZSOI
BzvXkDYkZxQkFMsoJ06nTmzX1pjhYB0wM79wfLgzhL9poJHfrqEXXztP2LUw8ZqF
QXzle1fgyUf6qvBDUSTCFMAbWrZJMJn8s5ZiTP4o6EOWy8vMBloSboZw8cLMPceI
XomeuIGN2LKQZGX4yh4wQ1rw2qEFu+k9U32vfzxQ6qTsXXkuicJiA/pckP2dxnKX
Avrazpsj0VMBDalH5lSFatBwaZrLYF/FuetENt3zgh7YJIXvIrWGSPzu8ryMK7bu
k1lGzw/os+qGQDBkTvo5u+3Uv8AgPoLHYoxNzH/AF2rnFsGQc3xsGdqvVK85kJc9
cDf6oT7oyspuOZ14UJBjGacUBhjypVfTh9GdchbsuaphgZocFmJX3j+jOgZKsJSU
VZUWD4c6Wn51lRvDwCZcTIO7oeqk1RXivqC3n1Wz+IMnQy1O65hjCrw49BCYTvRm
gh4SiGmUZApRKEynGWyyWya47TPZElWaiO9qIClTp8iT5PBdjWOOAKQOIZ0Rt4tD
mUaor9Wr+UMKW6D/RvV0t6QOlhFcc0oS91Plx5+RkY7o/wrbZu1T7bckQrBt1gAe
nsi8g5Yr7FcjSQzf+kNBjzGECrCaIPrCsotSxdtJ6wRC14MqGvwDZBOY8j5zvd+q
ljgRv6oCRr0FCUnAmu95T11WUr28ao1Vf+QVt0DVTjPVQ20qfb4kX+eFnHqEY57y
9D3u8Z6InHrfnh0HT9ln+ChYvUwXraq/DCTJY/T7H+97EoR3CCANqwdFdlm7zBq5
S6D/FiNj+nsxZ+LzhOp35hjNT5wDs+POgu04N66OqvksdwDafUr/3BUlqNVCv7gE
/PVZoLwYHEU0T9mwhYcEOkDLwhCnGygClWoyK3z8y18DjALOJV/zCq6P7MSE7TK2
ROnQLlzutLFJs5khKrEE7Lpu4wpFNrzQKU+9cTEBGMI5u+oUwvyM8MF3P6KqbjJe
P15FwmMZrP1JepYdTfCkfx3ZSjfSIXw2JbOvATAbBfW8o0x11/OounO5SowCu6Kw
eF3v3TvFsWrXUISBoVNSASU0O03D/73zG79eLThtGmfk4flFGXbRYjw7T32Yabxp
a/1lSBu9G0sMLgtfSg33rE3CTDcL24M+CluoYxKgBpQZOyZRoKMQzfEnpgXhE5YR
i0RWIOwER3BE8bgiMQ0J3K65nVi94yNn41eM4k8nRfAh4WHdLUM8jvmiINODXswX
fhOIaDbFPsezcLhqg0vz18gHQE/kzfOI8BpBJKAlwA6f2KV0U7EztkBYEPhWSSgD
xAKB7BfrFO2yCPR88lwPkrTydJSRncBJjXvo7H8rV1I8HNC5f0x2C3H/JcvLe2nG
BEVr3uzS5z2TEuo7RdDXMd6pHymM+VQRm+dzUngSmsuqoxFsNms0uGZiHvi25EW0
NcqU9VWLj2tNFH7N7u0XEYiUUv7/A34J24hgbUB03WPNtyl/WvBk9rsN7rVAquhl
08sMh7hDvKD+G9/GhYohtfACTkeLGkEItOQLKJlcBe7Nx6MOS0nYT1LVP5fcLp45
7Ob6cl7fAObRwpt5yiz3NKMmwZG8NpgrPBfeXzllHh5Y53AOuI7xrR0rGD3t5v4t
7wNwWX0LKJZ/sMiV5vZXeamgrGT1FaOb0cX5ZjmkOVv3ZvDfW2IH69YMquYPruVi
ac52LCISZguoDk7YXUbr6URlNkjfmCXwMK8+RlAaNLiG4krl5j8ukzYWdhxPz/Ez
cwS1AcyaCdeq2VAO3OAlTwZgZijAY68l6fzCmKYdiaGxu/s/PKO+KOEr6gHx8l4I
VaagLBSDyDpzrRYOIUwPKpTUHGqBbsj+LVhxRpUhWXNCY+gYkbWLEeraZHhgg9cr
p0ribFPQl1htHqvzHo/6Kj5SCfNaNTaOtt99SZLlh3YJa+uoMLuqEqe1IAcIuYBz
mp0NvH2WAxDS2F6sXH+tyDkiQEq41j7+f+WPONoJttofYNPnSuv7HDnHKdN0/v6j
McOkCx0y2T6znZE0ZO1jFdOOsbcuryC5jNuDTwKO73BW3+gYxdL5ZNiYnLAySiJY
gS7VRdzqjEC0TNf48hJ7b0WUxe3k8n+UYT6D4tNuDSxTve/5COrvgT0v9tbl025o
pYC+Kfa0RtG2CW9+MbZF2pYT45RNzhGZ5bQ1X5uAwWdsw4+SwSeGbXStGCdxxULs
miE4e1+sVmWRW8Gg38m6DxkygWjC6T++S5TchLryebE7mhucr5xuWu8XJ0wFDKoM
lwosWx6V72NLQJDkNz9AL6uGLqZdcdcWUEgeleapMiNKkUswGNvUWxs2P9Nw/jg3
ocPNX3LOHDz8ILMEdqjAUJ23Qq+s5uCqOOmFW6uCIccYaluojKbck4Jm9tz+Pgr5
kgoGq8AZKLbImhtXvH8IYl41fZIUmrUB4umRF3v0Y7fQ7TyOmizM1SgPwUt/Du5D
W48g5GaEWnuRqToFnuVCzB2Ps1HO06CzytZI0a5vJcUR4LEeJVs/lbd7R/fDrL2K
ajmEyt/Yppnw6K5ycjcuGgJ7IdY4gJb9eb5ETji5HzSf7YCDNNP8wyOOEwu2aMdN
euOfqsa/sLLU2cYIyc4kCFIWwpp0v6HVEfdRZeb44NA9XQo2k+YU4hW3xNPHR2l8
0ErR9sEV+8GBkfP83+vxpCP4zOtJaCGv3D5/+oAZ9cpZuawU18jlAKfvXX3BO9Yc
OAq3cWeRCreyX88nnNOAYkw9U9vRyH3RaEAdyOfeiI0HIKJHl9ugNOqqdI7lE5c4
/BWAFOCkSrWJPE27HPU9XJjQYs4+ni+LAq+mt/SkIcxB/aDVDTk8kvLjdtMAoxFi
yzknMV0scI+IBN3JhJQaULNNFYyeeahYdpH6FF4t66I01m5KxKUAbqlrpOeoYCnw
nDI017dMysgQCmwZoka6e41n3wH5QGL2H/d/w4zSNsDt4mtw2A+/dAlgdYvO1rUE
iXU64b0rTl8DMIlMsfN5YKmjRadS7aKNRGEW5buMeRw7615WsPMPrs+kRtLq+J78
LutDKGekhzMLZ/5w1owo3TYzaRZsGoD/hdmlfloDT+Np1KDYjY4FGIAH8WbfArle
tVvomOjBMsuD1IxxLrYdfJ8b4R74gMZQv4xClZeNi3vfCyUfmeMivnPv1HgkjqpL
3QagPe/nQLZiUCz7ZWc4tH3d4lFrE3bjqFtJX4oe4sa0CfkgUuN1uq3DbmWOiUmP
cz7ll5OQ4PSOanJrAe+72cawBpVlyoMjtYLuBzRy7cft+g8bGMS3roKsyolwfK6G
qyjmsAlEPgO1ap89FK5+JLvyd+2f5YnVJVctbjMnt6ISLg9ozO0++EspIkUR16qL
ofj1I3pG2CMH/qdmfzYDCYV/kSNeHzamukPGq9aAWT/ftcM0O5IXwenJA5NQ+xJx
1W1CHkhMITKA9XfyF2vkSQv4KkFXwmmWy5WLSGMOswKJ4lLYHZoB+RQcpaFkTa42
J0FR0kO5ePaJ9R+tvE/5PCuU4/6dkQEHofqWrcLTnZhsnHaanTe53yGckCRYDUlv
oTRrwIWW/6DV80Ksg7Aw/xXhCd+bRHl+T1YKUyZvCMY6GfvR4JyY2ATLlwtZpGBH
0kfW6C56iL4tMVr+M0O+lhqQTiCUw4koDO5rD23ZFQswgVCZmiAGWWb5x5NuWfuV
f81mJkUJsZsnRH3/Dj4D0u6OLlRW6Xp7BZ/VR+RoTFHfhFRq86ta2iWM9duL0gIE
1aTRVFp3Ib8R+tLHgkyX7HTgPwI76AQS3UbJfzB2j/qfqEyaW+fCLk/UWYaG6Oly
1Rmn01ZLpRBirbL9dpYoWaCFK93gQVvJeE82nXus2xrlUv2tQ7FoQFQi41iIfwOp
s1GVCfjclFG1klnJNOdQoQuQ2XekA7UCIMZ97FKNj2HyegLyhaBurszankiLXWKI
/nXx+JxDRoGCSV9Hu9hGq4w38Wb3oaoAtLt6i6z72KyKGsV0mssWFDBmlrRzLN/M
E5HdGxZR2Dpm4QzKZQnAR4mHKB+c8BAQE9OyHH8qDMCUy6fhdnYoGnkEyswWTr2P
ejd2TbsMU0xvd1K4ytLOQVNL9g8TvSdyzYvsiqKmhKrA/cC67InysdqkI+mRdjCr
ZEtB78aaajc4RGGsCdOSLrq2kgGYEXd8HG3XVthkgi2CUygTJYUkrp6AW+WqRt/Y
7qYhXwqYu4EAQYkg9AR0XFcXrR6143wAnJVRza7VeAw0TcIngQiHwozdFt9SKlIa
MdTwMZYhOm9d3pSQaLWWN1UECtkzRVGRrvHB2uqS0FQUaZE7zEqGTYMPggRyhpKU
Q2ef8n26idCCsSKNNOt8sHxu6DxM7RjhH5lXUi+pj8bNIVJmYoxZVTtQ/pkCQnKa
Ckec/jJG++CS49nnnAsi81EYhBIlExAmgUn7JR5U+2pKhmUWR61WxoGHHR8ejEkj
rTx0ujE1wim6Je7FJqFj94UBXO23gM6Ql3FwzCClmvNSdAfbm4LqPlFsD3Jk4A5d
Juez+beJDppaNWV/z2HWrI7cq0CFlkkhm29n2Vg47gFDkVCKTyo9kHPsmZ2rWPxI
Lptd4wnoGKvAwPIh3Hs/Z4p5cNkWiEfvtfEB2dcyRfT4vyou6LllNEz9OXtoq207
69ywmyQju0DIBFwaBZybU89zQKFIVep4hflzZ/jx6JWhhwC9B8SSIjL8SCxtHCF6
lObBI+B+/sxFnJUmsOsh50PA62xLLgjsZqm9nfZMt8GLqzDlW2Co1LXFMiTgOyNY
xFEo8Fzd69P36XRsmsCOcGE3d0Evo5lqBcXAHn7LkFN7YryRCgdX1aPGp5+kWrOk
oiwClL9mWVhiRVQbnwu/EwTGwJuMe8osy9WfdNPzv59NM2eqHz8hp2LiNshdFGMQ
2ZDRDwjsMSPqJmwODR5RYrMO2H1+6lF5C6Lj4U/ZuTx8/cVtsh53qWj8kENeFJH9
XdAggTqf78fZYCYbuI2OZ2cLr72Fs0jHlt+D/tK3UBi3jvMS+A8Q8pPnXV/27UPM
cSc3QaXwOll06wmeNviIqt9AJ4InEdDH2e7jpLtnZ94KGXdIBCnqXhzGt2k/gPta
/mbgXfN9LzFEWDYVaK5bTfoWuvBagk6eOn++kc5eSpduVpiklPyCmG9JFK4ERIax
EKjgDyG293OmZ2Q/ksKLAu/udBkBA8h/ZnBqVrLgR6UqIVf8oho71GF5gA7ZPvy3
xcYA6VwzsEXjKAw67xAhGpVGJipPHhLtm+QwTFoct4wRTfOweR0DNFV3Ci+5771B
tQTgfcvoCr/8AZfv3PP0JxNo044cFmESup9ugAc+KKjdQq9U1p88mEC0g8IDqjlX
2/WAjiMbuNO3/PYFQ0FnuDr1QjHdGd68v5PE1mvijJwg8vrWsus+t0dZREDOb4IC
QVWOTFylI5WB+1njQ46TzxyyGSZmb8MkIbL2rD8Wjls1pC/oBQBVfDhOUQIxlgLC
bgel0nxR0jRU97U9BAF+QS+h7tmL4nSvKQEZoeV/+lYM0n9/SJLFKj5FMGiBBxCc
CzzmILGQpwax+gaW0oS1D4BUvdZll5RURpz3WD2FkHZXC6CU17tqFz4RdZRX8+qS
RrRk1WCrPpGHATOPQFYUva/HqfjQu5+hS3vi3/SbLHbLwVVZaksOh3h7JgztQjwQ
9rB8NVISj5jHu7asyYsQjG7vxKdVb0JSf+o1FpDvI9INmTyTiPKe0VQPU8sWCJX9
QZ2ZSHujVa2FIRS4+q6a8dPympIoykhuLRW2oWqaFvzsff+iZgHWfP8hCR1d79YA
qrpVa52hiPjxL4I6H+stJlKF0iZ1Z+hhDBwwGLayFbEfxhwXHTusvcT7s076j5IX
YkWLtlJ3v87Jp2nYplHuEp4VCYQhOICsWLjW99S6tHpV8w035ROcfq3DqOVdtdYJ
2JGVJRCX/ttI4VprF99LvsMNYrHEnBy2899NArcHPKsGZvJKxOxEUgOqXdxF6VpQ
HyuTWsy26k5FlG1TQXWClm/gRfATq5fSrsI4PX6I/XWIoq+hP5nknNBUVsSkZwjh
hFrqNYP6oLEQHJDoDyNzIfgUdLZjypNTEQ40VcoqXoWgl+3waAcf+XE/CbrFCDGC
cjsw04CtCFeC4vnPHwVClata3nvGJRUft0v0ZWGjh7S5L64IBOSdn4831TL+RVlQ
pfgTLUE6lJRZzIZ4XMq9N1qqxq0GyCLS/82gFbSICli41tLITED8Biio+fufQp0v
XdqXMJ8Cr//0AK2orSorcDiUkOvJL3EjFMnCT+3SOHXrQ6H4PVPha4qiITVwx7zk
pUIcI2uiFTEFenQdK+UEIhfaEqGx5NejKk2grQAXZS0Q8oo9lnfsTryN9hcy7k3j
R7YMvPSTEom+LwyJXQkb2OasHzXSu7tnt4/5Kjb2j7jCqPUKVjNi2H5FgxRYVJfp
ensYrqjPGxAntfuFY2aiG9lKXbdD3l7qtP49ZLT/cszBRLsv9eeBjwhm1B6l8lGf
/+Kktg41gEDriMx514kJRAFfj44J6oU+b4v1jh8ZTdU98/VTmK2YXkBABxjBbeFH
lUhZvTFwAjooRlxoX0+Tt4ZbDPxcK5cpmINQdMomeMrM7aa4q5aXzMeEeW5l5C7g
u9zUSxcHFz7H9qhkJGhwuw3WT55Yz9dJKYyHO1E8AolcqAPPj0vq7G50nf6Zwgvb
iCm6G82AM1KsVxrYASMabahB4nna0hI4r1oA2Iraq0u6bMk2L50PIbc7nnpCuaJp
r4ychuYlSWXuabYpbkoh9KZiXOblHTzT9etLugl++DVRiEVt15zLoUt7mjlJ5Npp
VWKVBiqd9meybOIkbPsAmvZxPtuEXVNdcTTZ4+W/I+WmZ5IjHzm8pRqTuyY5dr/f
coVmylDXDypJjnSFkjPiLFwKgayRdJ/G0K2eWYXuYRcDL7gfwa35fbEokEDES2ya
R4cbeoC7ci60/2bFqHhhpmolg8ZdEdpdQWuxz34x+F/N9GD5lT5tVfVw4RUGXVqo
UqFgbKukymlxaA4moGcyfGFBb8ob4YmUqFJbEXujZBjUv92e8fpHFYUZKkOvo+OJ
O85f9V6WykPUC3P9Supo/0htkUMRfC4nm2Bv0CtSM2nOWi1GWNE5U0T1NsEglP1B
YeJPyxnqMkq9BMGgLjNj3pxFzG3XFjIMN/V7eTNhavt6hZqS+7UOtwycYDD04rEM
7IFjov3NsMh8S5b/SANSdLbQgLZOYAyJTGXomE7VntQKIFiIW/Nrj0XP/pWXTcgc
e8n0eXiLIJSYFaVKIoLyrvca7W2QwpByp1SiHXnupt/f9FvoGm8ncJROWeGsKIEU
LBLA17cnqqOHmu61sV9XIUDuu6HxX0Nv3/7OMD6Ky/r3UeF9kH4Ex762PnYCl8Lo
JUF181oxgdZwSvEyUUJrHj7edNvqZ2fQUb6UsVil5MPhkvS/Jz4g2u6LRdh3Xa26
64YCXS3VpnWvB22hPTWe/8rh5aC1IxjfPaUo/tAmfvnboCf7LxOYS1mHyNuOT4OF
+60Q5suI0VXW6W79vIXq7z5lXrNlFeqeS4Cxj25+/e1eXzDiyWufJGiIn5mITMp7
DiQ68dJgIqHzwpbniDWC0rABVNHFYHtr2CxTfpIpc+5Q5TDapvXhznqnlWXdvFHE
eTY8/KqTQ3tu5pOnXJBPAln+sIpgp9A1N+19hWV5SbXiQgwQ5O3isGEgFuuei2Ws
HwA2GHf8g5jA97BDJp9FOPqlSbeUP6HvUnVTf5aORin+nLptFebZ2kx6SYdxncGL
my30XUyDnFy0UAetlh/Dch8a8HoyGkeWmIasbaWKBFU58zPLPlBQ89v4zIcv3c3S
BFC3JFlKxBv/1FIOIoifC8IRHjioJJF7LyZAbKpHrP9iVNwuo/M5UoV20wXE0a3G
1ZLHR5FXnCyYk21z3GCRxYGkFSsTYx0WUWXEQJDBDqaG1GG3y+5zrxGzicO8Mfko
qi1o4RYxeGeUbFyYShAQKaY4Y8XdZ/MIQjKGcTBARrGwAeFU2gGI12AlMW7foapp
LHnOIo5GbFGtYJxQglLjkdqFxFyW/fwnVtESVhop4cdH7FfMKZaU+o0yjCNRDHfc
fBYKdBNQ54Us//armheGUmulEpoyFPuy0WgxsZjRYhcQ9abRk4cYYxkPi40B2+n0
0aMuPDrq0hqtZJpiZ6gw03zx8c5qXpP1uAjePlwRUAzsL0NzKgiKcUtv3vOW+kLT
9wlrcm30ePLETqDCbzgSDYeP4uBcX910B+QPNzhExcnD0aCfPHwNlv2ErXtfPy2X
Qs1SHMJOZUDb8H83+ZHSOaT5jzyaHqIhTvVOHh/DHJN4H2wVzS6KwyLBK8TQo1ae
9MtC6HXoNwzoZWhruaYUyBYkX2QOgt6ZRepiMWvxkSpQzuNLepS8U14fVe5nwuGE
JyUrLBl4PLFZX9oHsSOcPHYBhxdA+ChATsgW9m9VZjMIY9zB8ahlXbNFS6CPGB+Q
NrtXPLSffEIZOGY7sd49iwipxEnSBTAisAQkRndtREbJVH2+rkh1VtzKGsdp+rMW
dZ0agbaU2+gKguoQH5rXBUcO0hGfIPavq22M5PJFWnU2n0iukzRM3VVRyBTPaTuR
qpOurM9TVxcf3DNI42UVHwfiYh97wXDEfnvhm9ozRICupbQGww5B1hKxIr6OJBAy
9s3Fwbv6Pc0r3At6Pzh/OdHkqgkTn84YqRnT9qVElqKbSze1QvzrtyW0H/AJHUZi
hBqEStcjZ8EAifbmCSw2qNnqtrTXb+bUNJ4QUucHTQFHaNWofccX6t0znp4KirWH
aj991qUO47Ar7c2V55fnRjPwOeuE1ex9GsqWchgfyRUolMRJ0v1TiUAt6qE+BEVl
hbOwRahyQV+YqbDAfCPI0wQc8vCZhT/jtxH3M46I72S21LFY6XWnjINoxv6fVUZd
rMVTCX7lrRG/xg/NF9E4pITwlKgDnW4A7OR0sAewm0TJPt6XU24egwqrOWOEtd3c
x5RsX1R0X7m7+B1zEZrZoLQYt9wqTDddfNkfuRAbxZzvc/0kh4TEFqWEcLnGPNWq
Ld9XRdT1q74SP0hn87wAk1X5DdNA2hhI2LGXmZ+x8GyXgeK2wZI4Ovopvkm1UWTr
K0XSersherzM58mKu1mviFTV0czdoX7DfOigp11Kmnb+B8wI19sF+eD44sG8OdjE
sUs61dyTxIPPhZvHu2oI5Lmi7Uir/5eXL3p1sqH//4mo6j0VCi8ZWUegAgwuIDrH
d1QDa6wW87lt8eZY8WTfTPWd2r/8wSJGdguQU1b2J5d+sbd/dhicpoFKvbrR/WNY
aFfWUYydXwFzRPbpXTZzZ7C1+lP/KjexNopo52Qpk3Bg04jliSvabtJNPKMzYWB1
hSFXZmXs6e3xxC3PlqNJLpzS7rBZQyouW9cLokY13VZH0de6RIrzoOVqFmIyuHdJ
O8v5jKBsi9WXrjz1T+uXHJpkR0zdrLr3qRXZ8Vj0DdVdSySBXfIu5l/mt6X3LQVi
tw8jEoft6TZjribAGX7bWw5LaMek0KHkf09k2lRjYeeER4fu5nNy5v/0KJePxaBg
/b+Cv7AgjQS9AvTOvgQKnyvGOErqDQjgklkBk8t6TwFqoVkm8FHmVGs3qwY0rB2d
8+nQZDxAhK0O6EMiyGFiFt80ICXVsVvtkqRgywWFhGrsNnicvtJDgjEL3zsQM1ur
AEv0T0vKzmhDPmpdTKKyKj62wNbukH5jbamYRL39IYh0sbHYoFMIjX112mfWLxdQ
gLAeAGn5u2NZ+ToCtOhBIPcXhoUuOnUhAa9utGDusHLednjxHr/AUrlGDdu6wg9F
oAGiK2/1AamiT0dDNSaj3ihC9nj2bdtfRHdP8CAN4Lp1iJ1DF7SKc30rj8kTlwhT
u1k6K0b7UNMbcfZZB85S6DIhQ255XJhYM1D7/SIM8IBNwCNveMXlH7PBgo7WZMqU
wLaTvSyRuvdWQMvef4Av8Efc5S48FGANMIYEq9Qn/sd0l6xwkvivJJfaqMCPbvBB
Z2h1wi/UM/C9dRRHDKnNXbyZJsHvS0mgzRbdx4LO7xxpYfATjy2aEIPMi+UEfFTX
zB98CdVxCKWTSF4/5WFQFYTZsNy0GuVflGsuGxSPX49ViwjnbOscI6+9g96BYZEk
9tjpHEryg5ybHbLHrKtzGhQx/+Jc6ncg9FSmCAJ4uQwgOTk/fL1TLreUS2q62/n+
7hPOG+KGrtDM/B7FfvIOy0U+LbgZULOcMmFUO7mXtZk26FNMwgBH9LM5IKkKzuRf
0SPyRXrAXI5++SlXJx4L4PW0BRPnDLoBIUmh2pPBL3DYZdbwxRPN7bGM/zCOM0iR
X2LWnrXtf470lG9SlQsWZqpz2MGq2fJ+r6aaxzVbmPwA98D0Ksa01ue5de5XInKM
9/8VqyUwW4H1YbvO630FYAiwjPq4oY5AAk/qC1DVfxx1N0bj8C2IcHEpWXStCz6w
g3YObRQnxdDAOH1h1QFcOwg9TLpwbmmcSkqKVXnRYLdr/7Cy2oTsFfYzjxKATbdH
ByQUocbrnvNC4QSGuukkVKXW8ZBksFQmYrkkgyXmptja2uLOkYGBaU00HQ26aFyU
NmYeMTFqbQgTku03aoHJrQUFpLpvOuNRbNd2LpuFb9j8r1u2aRNNRI95yYEVfTFA
AOHV6F0AeZAYcHoVZy2tXdiKEyJ/BQzWgbfGGZha3/QxNw8uV14STvoRXavRq/d1
JN/OMbc+My9GIQqt1UOR/YD2E+L3CIyh2R7FhXXqT6LHXOS2M5QAkVlFLxgSqSUE
+PmI26VUkmHYqdVMPdX3yfxXFyZmnkLeLBHhmoEIbm/TPlBN0w+CaFrEdkDYVtoB
PeZwn5+j1uSiQgFygEgCh1TyVkQisynSoncyBqwxDjdSeCTzavLFmQ31UNJ8i9AZ
3eF9K42UwGx5Wpubgk0PZDGxDGNnSFuxN+HLieN+jhub3EOkMr8RRv/ypZyq3JYF
GSbtc4+1YdjDwYdoF+WKDuCFQYfbtIMZCIWPqRk7Wlp9M9kfTZnkLyJGR9kD0wjB
Q9Pymx/2Yyfm/c00ut7wBBijw3J8UEy9LZ6EfkNcMM/C2Mwde0jHrg1J9fhUqw9K
H2Yod5Fw0hkD84oTfsIeqamiabg1tnwByhZXS0qgLnGNMvmmceENTksk6aa1uW2L
ElbkjW+07CUlagSaO1Ban5kNvOJ2oFLSA11pP/s5/VNlTLrcZYmHPY/b9Eudg7zG
EOQ+xL1zgZT5Vw7NhMWpA1t/HRV0hHxIkjhzzO9cXEpcu7tUBx9c2ySpb6AQnkDa
ibmsB14n3Bcljgtm/ctksj3otwP4SS/iKNaxBfLfDzev+fzEMtTMoz377HLyW6Hk
tMNqnGYpJd9BX7U1/8cw0NH//YdMbBWm0MkmLS+JBs2YGmMZmGsdReHFSk7SoHHJ
Usrw6lBmjRUkvYuJjAIG3HLb03dnsE3e3kfcDqbkKbpGtxvTZYcPYH90Hbjlg25J
GJuRnwr4CEKPoFC5TZY3p95OAqT5Kx9ISyAONRqTaizgEZN9q80Pa43WdgX2f5ci
7ozbzykB5wZsMpUsQ64sXO0RCE8hfSMwrAA018fdjmJ/6cc8RDTSpcNdR/kIs5dI
ioKuseoun6YcnDSz2SNqjADSMlxgugO8BfkIKCJDD5mQIgswNDwmfW6ZyZGAWtop
PH/5tOvL40Uou98I16jz6Co+HJi2oWW1j7gPB6fm+IWs1m6d6a0fh0GhKhgF2oyb
PrfLEamvE0IfJUYbXYYXBQcbTmdN6wzGnjFiN0K5q6bkWs7UFSVZVwc5KixrEMt2
rlvmhmfveMDGgzHS+nY7NGoRO/VewQHuwY5oUEHAMCH623hylrlAH2hF4443FskP
xz6jJGHWlTknl/9cKN+fmgATY1hquN6B0BHbvUEJRVEACvs+pu0Y46Wxb+cV7Lww
2F3vDIn0oidvpyMeg0rHXJSVrrv9q0KDrQr/puLdJOg666dma4AQPT5vfbXCu79c
+r+2FokQEU+hMsFOA02w+bpNv6WQzb8f0UasKQVKo0vH/D9KfflOwGWe54/WgVIJ
PSzrEQYXg5k6yTX5vz49pYxMPFvjylWLSXpzUp5dY/OxhawuIf60Ld6nzaiz4I2i
QREDWe/2mg5HfcBQCVp2dT9CfeW/S9/arFRjR/SU1CRdnODv/wEsT2zmD0rV0SFG
C4Gk8C4e4bDCMd/Nrhff4hLDUR+iyWl/CrKUGYpUL7sTbh5qe4i+t8mM7CUiErNn
6GP5CGmYmMzzjQVuWv4JKcpHHUS7skqDNDzhdXGyUz645qvah9GQ3CvMzYsudZMd
MN5gFujm+R9FWBrf15aT8T3aYBLFw0Et2cV6DzmD3zKr0UtkXyUua1kxDs7RDcRd
82yI90WERRXM4hS0PoeGZ8xc5KlVvC7dpOIJiMvOi/egDp5He7ZRjgC3z6SQxT0P
W96hxaWVVGG5+f0qynpNSY1VEX7Wtre2BGFcJYCspOYjCyZt11vgRyhNHlSsv1+2
LZ+JJcDZdN4HoBJ6PjZXGm7alzc0NsD6GTkTPJ5OZO6OuM19wzb95Dp9XcUAi0uH
qoX1IgMpl6LsxDuqoat+oVaAaQwvgqZulA3axqWxycjIIGredq9GX3fadlkdbqjB
tEAU9i47vgAVl2JskHQS2y7u7UpjnCCyFwR96ReN74FISgwIgW+cg1gV1RIOvBXx
jsHjrrkJHKevdy6o2pjbfYJX6ZmsdPo8XZCiFv6bfiULMqEUpWU6NF9/rbU8arIB
4izWW1Qcwoz9tlQBangCHf97lHhw4SCaDdzCOiEcqgrg1He0sYISHFup5ouDVJzr
DCdhxoEpLUJK3TRGbRIzxG63u//atMcetU1rfUQkNpTkx3yjpAFCRG2AxsHia0lU
UUHoqM+usaR58aAOX7RqM88d22VAf1TkSMrrpbiebhVOCfbgnjueijKQbX3CMlA6
Zw0JWH0+Rh6PmdyI8SyB3VFYsnv/ozbFfnudcK0KWn6NiwZvCFl3sQj5g9FTvdTD
tAjzgFWViVlNoQuTGkG/aH12VtaMlU8jqRzmXR9wkLH1cvh84BntFqIupvyUQrKs
fWbjf+LLXrZdgaQM1g7ARuB5DGPYdBRM+ylVa6bd1jqt7x/NopI3by2KikxmQkf7
RVC6dyvTcgDrVsk2xJSeb+RAc2UkikcV24OvCHZiM23m7p2nNtvQ1MD0H1Qp31Zc
2R3zCy2nDdVWH/TdXJ3/DnOrZrdc7aP+INb8usxaIbPigm8aVMcUnw1dJXwwHN5e
Y/OQRU9/1grQzbgeTBxpghbXHuiJK0PNMvaQ2XjxEW8FzQnP8NNB565nppfTBx1Q
S4HGd3q++Qsi55pNbiJUWqrxyuwH2QNgEeGXawjEEBq86QOMMS1fWImVN6ydT/v0
CL1jQMv0oJtN1X6T4JL4jlxTsBW6Hr6zWDvDjxLjlTnKGXJGyKTvOPrPBQIJolnF
hglGvg6Z4Lr3XvegF+2Pt/qkD+9SVEjAE4CcqZhZ4u2rfcK+wO1NTFiiBo/ZPmvG
HSNvBFpbNUAcjPhtc06YvmWAr7SleSyFPpcm+8j5j7aiwJ76mrXol37W+z1jTY13
q9cU3owGa5k8NXIttiT+6djIKmYE5QraOLOaEjtGhHyUYTU9LGEgdjRNqZtanEoQ
c6CxqpNKOKpGFgXdtRtR516WWcgX84Edgmuos5UwFwzSnrts1hL/n9waG4Ax2bHd
wlCauYE+4GOxFHZ3vD6rMVHTuwdBG46CYKwMCgqyQ1MYTM9iGY7fdgPxtXUprBhe
sIUoIkodqG6sazqDHtnXIvOYJVRdK/G8cOfEE3zCQtE1HcrmjUxLoyH+sG99Xcys
vmY4+xbK+TU5ta2u0hINNG+uLwtkme9adbBPGkcnBRzBErjXTvtq5HIv12xOUJqQ
uk38G42jt7puBKvdbhvWiX/nkhiotgJmAdc865F6dhPEo/6yX0zH6YrcCXfACStQ
sZquqXeQ5h5B8FcoKhDcHnX5OEsGN0nydXAsnukrCZzt+sSH81LknWKpHJO89OJU
hvwaabE450ih9EO70IE9uzDedhsuwfGKVK+JNSjbX5gBHMXXIAvke5rlS8Pv8uGZ
Dvu3TOCoK26QkqeEjXM1sQ9zItXCk8OVxBR6sCWWruB4QXS4oqfoMJg82wQeLXZG
3wcgCz2fLvrKC0V/YjZAk4rekkA43siYebpn/5Aj0BKw0GzQbw4wGgskMYT496tU
vLXJYksR9K2R+0G14Bk7QRjPmiXfsI13+YeaLyzEaYlEukMYOMPEL9cKavMrpX5/
thIkMgkj7WlQfYEHGU1KD/aPj9G8xBg/hOknNVt7Lr0Tl/QWbQ8cFznPv4uGH0Qm
+4nnjXRWKmkHp7U4OxputYiUpF85MGvEKx7cfXf7biU/Qa4R1teWXQSf2alt3f82
gI6OOGVTY0ugHEuLCbrhruFQ0FoJRR3ZTuL1n1eq3fe92qPLUwGAVUZFqS/Tg0lZ
h+jkPVXH1dlHYKtJINbrrEPxrITjzS+f0ULN4JZa2no1bbgZ4LX2duFs4fbBbJgX
Q8Mtblh8WE7/Cjlj2iqbcBBYP7jgU6Ja7HG9iIItBysNrEdWRMtiTty9SXPlyjmf
g6qL+/YHwItqcFxf93pcoqIeNsF192zv4zm1485gGOg6Hje+e6jIm1juis3zw7wT
bWmaimK+r7AUtH78BgWVS01WKh+bk1B9ifn3ey1B/1wFhENEsXIDDIwFbIFZ6f64
gEEJObosfQfgBiA10tgCuZ0WATshXWdDkH/5et59bmUlnUQWgWE3JdsWnz1aYZAD
zze4/6ykduIGuJOJT7tWkSn0GXEEwRID3oQlNURvSu+gkLRk6pMAaRHnG3uyyl23
7k6i7Xrwy+K/IGR0RwoXh93H14hE1xqu+KF94pwTVKFjJGFHzHL0VloQNfJjiO1U
UZ07lAJ09ralIvEf30ktvp3IbuR1yF8YfZoDs3fxdPcPFNaBxyna1S55wD69Gxpt
v5iFzkfy6LCN9yUn3atR5/y7CWRgSoqdrsIdD56biPVoBuM1mEWMn7l/nrRagTPF
nkFbCMHfF8Nqiq96a8lkQc+48rOPTPfApM5XscqWECLXeTh4SbwavgHNuxA6rwMt
tOeyRtvNSJMvd2L5LAamgIrTCDL2PKhMdbs2OgMgLo+sgJOcp0d258Pp7r7Sst5/
srPzvAUErYG4Ieor71Ejq/qddw2SkqlaCyd/Mws3r93VEl/HD9GumVt7E6YDs8yQ
39XJJbJb9IAxuzBULlI+GghcNlHNF6ryTZl9xwMMt7rkg/pU3wi20ghMzcKJ3cia
zaQydYdpJedKoVJiwW9Axyw+65bFDLT2WW21tixVJa+HWbdSG2g+lccFyEnue6T2
X/HLx8PAfsh8G7rVKhAn47cQnVlsI+QcrZzvArib7CDeFGy39sowy5gZh1z03Aw3
w0J7iVrBhCmfFWxUq6Tp63Nl+gTjF2XSM1Zl756lO8dADH959QY7VH5p6PrE/Vrg
7N7yx3K7US22zq23Qfy5i/gU2VmtFFOf7/JpD80alQy/aXhge0FDs7ZT8o0RdwGv
XHpB8oMYXCRNjzWNXcpnu0HB1J5wDKUVM4qhnANOSGsT+4jNcodAOMIj8mM0VHjH
ZZHpL3793WOiiyCwUSFPaPzFptoVyCsBN8Bm7Qgb7mkgGLhfmCDIRfwplX7Kd811
qZGcFzJ7qePHUBsymn6zOM/ZBBvJ2V+k2xqWPZfZvTaPnuBdCHZ8Lvpp76ixoy2K
0mzRVtHTgt0ThamLTeIszCkI0vMOZ/2rbmoGr2K/bw+H03MzzIQSPh0eEi2uVeFG
Yiuh656DBwUcecfpw/5KBnBHn6yYGsS9MUyhd+JpJo380gAdYy6JA8lGlgFtTtVF
G7zro714MA1fpBkxrkgMlqReW+ffuegd0P4dM6alWYEhI3tr6jH137TaHtsMDp+7
RaQbo5TP6X4TbMUHTK/MC/b1SZc22KibVrVJ99MhcDB9d60qTpyzt9DVDtajEeMu
3BHA36UhaS1Haq46HhmufJSZuuCuE8WxVVJZDTi+FKKn4boyc2+KHHOi7dS0eevM
olDqbIxv3reQ9L385ACa0h6/dP7rpWyITfg8y+hgjg1ipkf4HC6DsyegdMBKL6sD
+DC0djqZ3XRB5SUqIB9+v0kjQOYCn1w+PHStLCibboPSMLjdxxAhe+JMiZ3/RlSN
28TwNRU3bR2T4urt3oclyz5byfsKXuSNiNIF01O6Jjd+kkGh+YL1XwhGpAAI0E9q
GLNqHrF3Vy0vF8fGTpY7OQpfNvxuvPeJhtwJIVJB66dOOtbXEusz+GSf9z3uGnAy
J0YhwigVPZ6lyPOFOeQx/Ilwc32EIVb3bOcnOWzuF2AJvxpkH2lIWvjyns+n/3wl
WETGmhYxphTGSAH2eW8xvqYz4ZB7eVQMwiSYvoMDxoral0BjVx19Tx6P/0/o/iz/
C0BDbR11VXNGmBB4pqw4z/lpCxjJpUgBqJYC+RILtSSeLd63gWHXjA/R/M+Wo1th
yItrobExygcuvp86/YlKq9ig44yCIdjEA0v1wQ7T57HtS2GWj2mAdWeh6uXFrafY
LxRRBpCpJC3JQEgmHtYsxt6Dp5PgG1cg4wpGCszKFnVdwtLj4//E4nPMWNdIOrBu
jbHWheG6KFEbhoIiRUAvqEflzXdP3pMxSRSjpOPtw3rJvIm7DjgCe3+ZI8bEPwNw
XFgI5oloXKF0JF/LHi1rsNVeyYF0rSRGLkQdL408De96PdtZazNPk2zxLQDJo0/Q
YrF2dfZpRbBHns8g2H8ylk/Fdwtr9L8894Fge/luq5xJ2Uv9f9W+7m4AOVoMkQ81
tmKuWw691UKDEXzkIk7BAQXI7elkq5qXHl5TH2W2dQoBWR0MAGMfGStFbqBrMmDT
VFLU6DHSquTgCvfEDC93iipGHejFedJ6nLB7KSi0w4mEy5OCf57P933gYYn460q1
ytqUgM31suy/8Y/42zrbhGC8HIFuoGlLtSZqdG6yggen7lpo9tPsWvqxewdGG/b6
YyoBS/9VCST7ncuTjPgXKig4eFCmIdizG2ZjDaBVAeWgvCxlNX/gAJgKa57T+MGC
zm6l45AeiFzDCEsxsqKMUlux4dqigvePjLAphgx3nPrBWbLUg0Xo8OCq/ZTJF3hg
TBeq7U+ehPEoi4MYov3bXawhe6cNspuywZ2aw8pVQBEik6x1WVk6KvMKjqueWjIk
nKX41SS6+YXdiZikbijrmRzZrdV4D9WWuHf1/u53u+ND1bgTQUYhFdeiD+NmIWAW
JS3AypUAonYvjI0R0WHixlbGGTPoAFnLH5t9vUMFVq31jJ38UdNIwapYy8u7j9Lm
Q22L+me3op77yMKYb3+Ljue9AvB1SS+bKQWfEZqTKdftpU+lDRzukK14qqHMHNZc
Pk8jYgKUAzBicEl4A/re7AxeWTQbVsjZilJiSuAWDoIOGkDquIPSf+Bap9YRq03g
PDHzhlwuj6DeOCyLZbzUuWfaUOmNJEFfsyAmSwlr7xLY2473M+2HPIgOiamVZxDB
YVgNczKCuWL+y6kcD13RjMcbUGagKyjmGCAvZMEDo89oPiRi5hEzx2v9akbcquDE
2jAjT5UGfHB0Yhe+bY1DAiOPQnEp/klvpNV0SgYW7ZPT0e5gpRZ5+KuqLl36REZb
FFDlCZXnTKh/JIEn7745Ezh3T8jygS8x6K90ZnhzvQbvUgf50DDQ2DQvxPZL/iuh
/WoRri/0Nt1UyiBg/cZju1gab7RG+ZZwEGGWIL+CvnjdfjpXLZQ4C1xw8ZSeVFPZ
iwLPO0sVs4yV9348VIe6HdZDqc0Bii9uwScMSDJ+G4tn2j59gi4vKUZ6zSL/V6vz
mpjX5pMCeublt7pD6Gv3yNuye0ZHtJTckN0Cd0SP9y6s0goHKEVxr8RsNalWLEUA
cSpeK4hLxNPG8oHZyN3OdIUegpBBMPWv1uj4EBK0XsTFkIWTrryGZJ29Qk0oWiAy
k5/tOa+r+OCpwYbLti5NpffP6YhK0ORUVYxRpTtE9esAJYCE3yJ39adCwQCjYccL
ErB0PtSV0LEFhE/oQ7/ZpOYbJckRNtY4E/Kk7qQ3WdJnuhW9eU+e2NRxD3ZhK+2e
lNz6+TYYNu3MFR/y0skRDh/1IguV0JiDrx8fWr9kz7VLDDBsmmK5hpGQkPDkJsAW
pmNOxgh2tNe3LmvylmpZYqjEVJqde6FRDfLmdekZ6gTa9VGAC6miwvkfTyt0N0k7
glE5u6Sa3tqAWt/odmu+QNi3J6z7vZ/NaWIL5nij8H4QQEtrIoh8w1g0d+/RGAdA
GePey9fXsGAVQT7Y7Xc/LQg2Tc6vgzZ3OT4hk+5mAuOqKhlfWyOHU8Nhr25v9fMz
TaYDsF5a8h/t0O3MEhT8FhbXpBWQCNbWlw1dc6HfcBybta3VgMSAfrbo+YDuCfU6
uEzEpNrprh4uW6SZtDbuUATLRzMs1lK3jLBfPyMFmkaMIVI7F8mLTQYr9i9QgmuR
vFoCBgp9npVMrMcvszIGiVRzFXIvryJkEIBpgqA9096drko41fE7V6yc8Zjq0u3l
brPXcAJ3dzLHXVF8vwii5ZjCUF12D8hKIajrIFquABo4EJalk2y5YyG7XteMugWw
N0AqzGdP4Q+RTQER3ped93obavXZMk4hwOnPMQjbuGBgDzKFJK8W6MzXeQQ+/EuK
rAQLbAUSF2jc4Zp7j5VWpginTfKAOurIv23VMjjas+tiX9rCf5mMMfyZxoNMXzZO
/gdV+JvKqUhD+WDYRcUL4iPNDToXu31uPikjCZQ6gcux4h8tosX3cVJMWxdXU/jI
pWNY76L6FM6pwIIlUy2mepyUw1VrjxHXb4IoOFkd9SFiw17JOXctWFZEEAvOV0FR
CKkg+JzBsESJ11WIqQUCU0jmpgKNLSMb7XqSDhy32bf/+2ZcmPJXP8ovryAMYchx
4GZYioZ/bKDfM6Yb0PPu+ZCE3woH/EvB08G3LNPKZVwT5QiYV7oxqlneeRWiOxaR
HVtC0NjHOzSHklruzyZe5H609Yz2zYoYqCJ9cdYIcpC8/BXCGDDPVuVODJJsY0cV
qfFMdetCHebbvlTkr+8+BJdUO9tIaR2mDcoUKVOK42wwpVZB9v7p2cmh2yOa2YZh
IeRH3ME/crNaD3aDj40GhVnQFw/3KolOsaYa6X6drYBAnP52X6RHB/C7l0d0ro2S
Hybkev3a/I41OyJ91paDCGiRE+jgTHK/MYO0plYp76RzT0W1x3JeUDyA0FdOM43E
nZjSYTLxZR+wK4UGlXoOSt4T239lpSqbPVnMO25VHPcqn/KHzO0B9MJt35Gnh5ES
AWakkQQG+S1B/T8ZOrDsvmRzR2G1Tx8nTfzXIBBeJpdjGJTe/xqydaYl/dPE6FLx
Ugy0Gw8LubqYcPlT7CZNrYHzwZCEN1dPPcBl1tFde10uKEk9Ze+sFCqCGmVayo/6
vccJZFe/O6z6j7VOk5423IkNxtzBYl4AxRRKqGnipZmQNShTffxhp+dgsAow22Al
5/a8NfxrqKA4txPUtdZDz8DOkA8CdarlfmjFcijsvugecbA4sN4wCQpiiO08EaUz
7G5lpHNVqgrDnpBnKlliM/bCCkW/T5pLt2OPv7z/LO+61zHf0hnC5md3gPhc3jhJ
AlC38oE04Qg7hPu4bmhN2VcmzsBLdXa27RdN9W6gSyMn0K2yLlwxiTIaZuSujfUQ
KAA2bgp1osa+Ia/cnXdmFsKV9gLjAi7pQe3qAabdb8Gz4XOpCTwT2t5CbuAluXan
961WAhyZyTgb+fUZvtMHo53DsDriqounudas2VGnMwKCVOEIKWDjBmGZvmHlQ07C
oZs+3pDH43EBgkPPmVKIJXxQMjdf+/Vt2ZRxjzky7NbTDre0u90J3oZy/h8FAXgN
DAEjXGIpTTCLGTQ8RsZN+umOwnhlNUJek74inw+wuRucMOOBceJIkgYx/BNKd5/X
ld8lKMhDKDQLom9m69lej/ZySodZAuvt2wr2FwOpEfinkqgqY1XuMnHaA9KCADcn
u0gdJYc8RVqgvUqL/d4p1uMpKlTZvD7uBDReS1/vv42SseQqDnULMiAgaoISHEyF
t3Pz5IiWueWCcXDe0hVE8ab9AVsGXzD4bgzBqN+Ra6SHCJ1Sb5hJ2EosCj2tMhOC
DuXYOGnWBl8xFsTcB0+/AHf3+ImEhxerifkH4VFqmqzlsrFf0466Ut0yv3U79URo
4XICQYuy4/UE7E/HIWwiYU5FNVmNpWpQAevN2KgIl2cggyv6qLL+LoztZA1Tctyw
L4kWtjaIi4tYziOGCnHA+DJXwJyiQ/DCVCWARbCJ9jxHtv7pXa9pK5nQWujwFmL5
qbNZAKvuhyQMWYdcTOcc9YVBx+uRWLO63eS0DRL8HlbZKb3QmKaFIztBJFGaEx4N
M6xiZaXtMR55t9P7J4rGahcx3Kqb8IUgg+DQRY/NES7ojSSwaae3JqthS/J+ZwXw
hDtPfF/W9vaE7ZStPk6Z1yBl16ETcEQtcS+kPV2W+ukGEXsGbVIUAO9+8Ipa3t2W
vyB4Qq/c421K1DWXykr3oZm7JzBVGl49O8EVJihm2/BDC6bekxrAkazeJ1tVe48R
lNQAMYTwYp4NwYEeJvVA4WZ9Z5q5Uw2ULqFWk7hGTs67GiwIDapbjkspP69U1rHA
6aN8oew3ZvdrJfMw+CCQ2THb+xnIfzV1VlUL0fO3eHUqkA/FMfX65ss9LwkK9QT/
K6GVDi4q6iu5sPbdDA4v/RDdaJ47nTUyVMmQPHPCFj4p6MCPcUQTB2RzlGQWyZf2
Bc51wu9Gk9WD6ej8cVj500acO08FIRS/Ho+aNCDDXIxE5kXTGMp+TlWFsMXd/GXs
vidxEQDdbHo2666kODM/e4AxvY67t5rs287qJ4uRaUzTaAoSMaRvMBLjhOlTBM76
yGT8GiCEQGnAxjgbaHpE+h2tB/8WOg1WcD1XMf2ZSoSAaPXMoCGqI7/riSoAsW07
ylNgz9cT0h4fcIb1IR54cosHzBuIOORRhgusLfMM4nQF5HVwuIx5sm7E2/zI7ow3
hGOtM+P7rxkJZl8E2hDGzBNygMgc4lna0Tqss43evqGOXTSLsLwlIgiFHbUjw52J
UJwzQuKANvuvCjUlyCvDIgcEfwhaHFqWLEX0q/ToPlv4YNg2HYcPMo/oiTJgp6ZU
ShL77NYCkRiFKAIyLkbQs75nAmtXq3SgMITrqkpD6fPmVJfie68aHzUVGf6n5KtF
NtPFB2z6nY3i3yuocbqaf0UEHYLpR0q8n4Qevxon1q5LOHMXbjXQpQwg6pi/23oS
krNMd16hsPUuUFkm9uqNd5dYi7izx0qCi1TmU5FrIAmC+Cs+ErNIDTQ57hFhKn2E
FqfXPpO/JLkar3SfguVmBqgVYG+86WFxyHVUIuziUB8j9MX6SGqVPu8KHZ/iL1k7
weu7B996NOVgAOUiiZs2F6Xg7WEW+cUYCiD/r1iOV2yCRRpJWPCVPJ2Mqsk5JyA3
CjPOEmbPfp3iof5WUCc6Ai36cGtwA6yfso1LZCz2/A2GQNqu9OjRun4dxKG7cr4A
iXO/IfOWLMBiIlFFMU82wveoid73sjIVtA5G5YXQ1WNly3mBVKg4vLi2G/dDUeJn
943GGQNpWrS/inQZTOXSmlJgft2OvF05VBezawVFuYBTDqOEpUXfviPI2zeEcCN/
jEi7iEumKxrJ9LLZi8YqOD3jiJ3WwxsOxx9PBf1SH9EkIN4LdKvSKOFZtxf/pGEt
Wb9mgJ+pYIaUuexiamr39Bl1EnjJ1/KbNnf4Cyp5QSCfRDretsiNSM3WNBd/+4Xb
VwCoHUzMAMKJlAGWXPCo4yl7hub+bVq/EcOJZVYFkN2IvozEzigP8GUxDPNVY2u5
24EwJBMUTobYXSqLdepiiMpK1S9ZSVQWK0srpq06uDJaleJ+SFRR2OzJjFaynGm7
T5jPy3AM+Xb5gP55O2A8Lj6aVAw76i2yQaH32PwMjGgQYhYxy2eaYvBqEeZDvP6r
JD5ozNIGGhIzsJGyABpG1lXKtVxX6wVv+XgLZDf+xyx57g4VFW2EoiJTOuC7O/4T
JfORGZSO0zqLhgOjklyo+dRsE6vF8fZl3Ln2/2bhwN+AfF3bqUilIzS9pPUm7qmg
LsvUfKnhxJDMcpXX6AcdHnOX/o4l69xA1xkoYBgVAMf0Tu69bxAKZ0gK3YTZzseZ
A5cbjekcYsDFzbYt5LijJ1wXNyGtgsQMhUiKchekIwUJ/EUSb2HVI+5iMD2pf+Iq
2VpWGpgjCUa38Pq9ZysJ87MUTleNZ+GZUUTdwW7hJZAYRxUPI8kHp8T/G36oD+/v
CTOByRXE46aSlZ95DUM7khvW2ovRWNH1oQBTNlgZe/QzK53Oh71ZIWgVOPanZhMZ
0TL7NC/M4fB4M4iOIcHkk53roEvMZxAFewEGOgR4rFle4oiXhKTdzZCCZGSTbXgI
dzLo3EBreqpwVmkOA8exi5sKxSUvAEBsP6zqo/DZvcvuUjk94uSArmtGn0s7tNuM
UyqZsDn5Y9OaVUJmY03q0bOqUB04/IdyuzgPDqHmnEWSZtQrk2TrBm64uOfWHss2
cVKTeToeR12PTKsIFiSiVCWuiMETW0jsbbB/kfHTMqHhrZBXbuM0VQXT4/Jk44qi
hP2pVoRBhQ1W4x7Ig8Ss/C8kbuH0Y9h2ouObmRvkDEeavYFuHrZI7REHQTa3VkIc
eMgRRiC3BZIbEwY2fD2slr0Ys7JjY+4OT/RXrV3MZQWoCLWTm1SWc6c5BdeH9Ywu
fwKNImipj4pwy6xRIqkARh1AaC0fIgrh7G2tDaHMlD9EAQ8oMXlwwLN8rDerqMCh
pt4dDjptga634zLj8p9bpYRzlWonI6o5mv7hPOo7MmLbi8spQjQa+iF4fgxx5bgZ
J4v42Fn9Spqj2gv9Y5VgxtMpGzbLESCVHuixbWGXWM4oG7r7BV6atnxCo93qDJed
CLRwUKOYgXkZybzkhi0YQtFS3I/0XccQ1yJwE1Qw2gYYhLng8lWbuRPOxCINx2Z0
fpLuF9YrafslvRnvPgSrque/fXX116dtJ2MjxVSl9Vg60HcjBC1EWg1Ew50nl2Ls
Acm+yuVUtqAXy9I69ELbH/suAa+9bvJkivoxDNpe95oUiPs1TIk6AyhUQw4c1ygh
2/WoSpwZ0W6kcUu8OltapduWkH2yBUVJ+I9v6RPD9lMeMyTWV052XolYKkcMuxTA
kNcIlxM/8NI7KPplxenDuzBPpzM3AE+GJPuFF99aJF1ZheKy7QUpI/q8uHDnYK+A
UVGgaw4mbceM7Oje2jEyd403b7pP5pkAkyifjTLfYx/1wQurIH/+Kdu/IZ0ks1/e
9VsJYT4M214zhB4qzZiRoRbe+M6977sHgXuAIw2xHhNnInytmNk+BcL9j7Zs5OrU
Y+TU1woIbVswSQf0wvHnij+NVysEV3gXT9gQyOTYs/wLTzoEbubv7UGIHieyY+y+
EiWkyu7N+rsmtOtkm5Bna2LXg5sv7o1I+Dra3hA7oLG6iUPAeCwIhZchSL+D8H9i
YneWEqDB9n+Mln+77qX0X4vmtjVJfYAvP/JEECiSNk1VhFqK/RhCIE4+6OkKXamo
C9CljERxC7M/Z82horl/Ur2IEaiORUXxAk7etUgur0c+B5fjeNQyEOOh23s/efF/
dZBwyrdWFVod1Pgd0C/6nYE5AJWCqiz4zTGNiR+aWkbHf30/K1c2kmMl7MNfrw2d
SWevB+vLQZXAgxTLrfabJVduUhqU8gGZUV0Xck2kzlMW0nG8SF3p641NJ6ibBTD8
8kwyRxjcOqmVc0dPgTSzEVaeY0JT+c5cOWmc40U73jWFd0REq5yXTQiz+kWoKSUf
5DBIwKiMl49gY2QujNreRSi89SyES3o7LWKwlG4m4AjFpL/Z3KMcByF7rjPVb7LO
K999+SxrBLZS8a/GFfeix8OX3UVWXbji6NGdWWHh0X6SBXIAjeJzdOf5MJV5xtDf
TgG9/3IPdq77dgFD/vheJu2s8+4AH8yzD/1hIGc5WlULp2xXfmD+NxIGqrWUulyg
pj6hnXdzyOe5fQ+/U0C1UqBBku0myKvo9bKRMlCZilGI/53oPHk4oCw4cLDor5nw
hKfbRl4a3xRZM3HR1W5NI8qGR3ZLvCJRvb1N3zMYtlOd0wYyg6i8a8llu/3bXHws
KBKiEX19ry6jf1EJgsLJJ7nj4SIGgGQdv+PQm0wUzgyics8grXqDiuZdfLSPiHIz
ycx7ZobfqsANnY4UHuK/yVLGQ1zb0/+XYbQ/OTcTNbWJmNHoDKnbKYRlAxXTBOqp
Wmytf4j6fsjeMX7ChErP1idn8JmwSKVhEfS+eSd9iWO6piR8JoMO5WU4jnnSrFmI
M4FowTsGf5o+O9NQwkkXW0d5iKruEXDpdSJCf2teLFNxh8c7TyDHYy1OT0d9+3MH
0J5PTUmCtuHgF3bBL14mDM4Vy9JFuYa5iOs3MeiWst0+NowiX7iBGiqFecr0OPFE
sI8zpx+w5WjvYnHHqTkum9ykoMi7f/S+IMxA5xMUtCPUUzWx6gU2Vxc39EYt3/4/
KEaz3g3isog1fDhCHhihA8AcnXrhEGET7FtBNsiT2pT/0L6wf62oLb7tvk7oJrtL
UMtEDgFKVGiqbReZN4IFHaRkg/eBBRvEzM+/9mgpZijCLxDY8ixYHj68fLLYtg5a
0L0r72Txj/kue07vZJqnep4i9qVD5qcwWBhxtULS4zdh11Pz+1IklSW7afuBJnbk
b70MsSCsJPPkKxWl8OtdSTuqLJi4jjc22fxD8FTADi0xl1/sbvfBfiVxSasOAk+H
qJo250YF07DUt4B2I87nCziRgHsHE2VUGli0ARQ3hzgPBBGePrAvYQ6uZb07uOMG
fvU2mJ6eGIIuDNV3e1bdgMLo4WxSMFUvCEvcVy1LU/ZZPVjf0k8bNvfXX935QTWO
1xRuY/Uzf2Qgr+X4yL4YCp5XH4gwmWeKoTPv0ifNw4iJJ9I//VVTb8UB/g/fx2zQ
aKpLvHjPZ56ib8Tou//NSi+HJTrD2JnSbwtKK9yt2jaaGyKPJUOQ5FDbcEm/A7f1
1tRtu4ezYN7PEWrM0jo7+HUjeV8J1NHeE4Xnk1gmmLnfd06/p55DCEMNA6iH5+L1
hNnbv+MO2vaXq5wPl2xYuQ9o1ED5CooGt50U6n62x6nykV1JqqTD63V5Azyf1u8O
VGNmltqgbEmChYXKk6+7FuG5aAl8fH1xYbGdKpLJr+CNEku4oJ0XSmEO356BR4f+
8urnR4icZeHEHYiMNliim4/5YpQ1FUSU4pUQ4K23+0cXX5ZR0kWhSVcUMfVcjaRD
5EraIT1fVMTUk1fhRTEa1BfJDDQN53axdtVooo0YkM2pUrP7C/Ikap1kJpeVqotB
Z1xfPc0Z0x+DcbXmoANh5c9XKOj/KBemneZK24FIWZChWcaR+NhHpTCV3QicXQvF
ZH1Hy+rJRu9DASb/sUEwCXK5pvFiBTR4PdMwsuqQ0TAsaZmbMlxrTl1fZZrPAo3o
HNbEpo+4lBMahO9CRoiiXBu5uJ5+IKvpiRIS4kwzH4elW6f413ao68Lc7p9MyyBr
ReF/zgpopfbVxgwV2IM1uIQJETE6EXlnL4vNvxM0HE0bOvd0NoCB3GE+3bzyD2Eh
mINAWzyY0JWWog3z+p+5lytunprYA5BRHVZWNIRAOucIIbm/SnpZzabmo77iQUGy
zdFsLk/PX44eZdHB49zBSKI/1gVIPjjfDTP+XDccAz/BvB+OCzqB+yHU7iaW3QY1
VH4l/8AWiiTFrqcnT/scYzZWYrgPpKGajOqfU6bVl42UXfjWLnrIAfj9h8pyHwN/
TeiKtT+qtRhuMoQjauvzl8k4DGy9JrAsR7EAI0S5JhzZt8b06lKcBsREKP2LNvjc
bJ8zSOPlab17uJj0sUK61eW+ZoHe42rMvdnGzKYwPXVWRZtuFHiGsVMcV1Ts5WVc
LGGAcHfN7MNhvJPW0I5bSseATWszzywoRlwssquWrqDVgZKwMiioqzplRJjUuyvW
BXMjws1vUDOAZQiTEWKaeykAjzXmfMsN6Syu9ZYZJRW4UIR00JyUZ1LiMo2Or+ab
8OvUJGkgeVgDWtJuf4qTsAqsNoEaq6DQPuMoLmiabkYtBJFzf+sfBsA8REqAxZ0t
uR6Hc18TM3qZJ8x9yoK+ch0Cbqs7X3Ir1XINo3meSdjDFs0SDx3t4XPsRlimRRGu
/0dbgAbuucPyFjxIPJ7s9pdtxLjmJ5kuRTcz6OlwS6FSHPJwSHhtB2TKN/Ce0KwC
DXHVueeHMRvvvzTdhWSGuedIc5Y/qWxoOzVJTOlUmvxU95jfveqGnryAXDKZidm8
3X+PlxUgPjJL9Z5KUIz+ZuegYjv581qQZWM+xB+mc+mxfXMBGrGPLyKaAiVOVMQr
Q5RlKC1yflO0s4rUtV9fpSxMuB87JV6qrFMeNKR0rqTiO8+d+ncVADw1rAn9lLJW
7H07cE5IqR0D8GPwdQ4fXD7gpeSvR2k73WVOfdS1XW0URLsPfjed6j4XJ7QoG1Wq
EARYRx90J62ZOtM+q1laS/rI/XVbFGK/DUrQg7GVVoQuDr2rS4cpB1n9tQPmc0t8
WPAGVlkmcnrChUKZMaBnQZniSg+r/oe1qyza7lKDeqy3aDH51OUCHaMDQ8GHZ9gy
W2whiaHF03cemmfKYLXujRimCkZh/aphMLF9uQba3+wxpS+BfZfQaRVMuljSy6e0
TswNXyQ+GwXCSE88fUeUPJYws3gZ0WqEs0AZER1+R6ewqKvNoFPwW/JCQXy8ubxj
Qu7dxSl9zUUFbBuxXvZrLfFpFGC0wJYMXfYhPT8QPJcAr9LeyA6HPuOD44LPMMtB
JNbv55jp/9Nj1H69FLThxaf6kbArtYZddS1jgliv41B97IWF0otb07ZMY/L92qSY
tkOUrIcFIyExZk30yV8APkGAiqZJdo5Il1hWCrJGQtWMYeBT4QtD847pD+oUU2TW
o82tTsSaweASYpDDAM+gqaDOHUumFNU6GZdTvTCLzqJjgcMk26RhEu6VZYm/K6Cy
qnQ/tyGOYOoeGe0IxfEjMGe4qBqBd9m//wRnGDGa2hBt0QbaKkIFr7M50GuA9hPH
J4Q/yzomA9HDHKqyDGEZYjJlm/qg15er4u0F/kDWvZiTbB+HghC4VT/Obj2uhOd7
hXXwD0bMkCzNUu5W77E8a2D+9Q9+NWb/3sv+oYA06EPeqDBoF0PhLodtuhZTBo2Y
nZkjeDbLc/Hdcdbzc+ShnEvaS9o8aXQN7E/hZj0ip9ycWPQoCGzJqAwDQkEuV6TD
XL5qaVSnhxh9Ad2+CtziY6dxa2CCxCwxqv0udvOCwAi15wHWDTCfgxB1ML4CL6xY
Vz6T3vfh+l+kRtTHDLMKqw+EjuCANHaESE8RmXbzaYoZiSf/4HV3HHDmJEihvg7k
ORjAeIGksNNBkYD33u3G9dRuPt3h+U6wB9pqMkhn2QaiionTw9Uonv2EP3BraXMv
L6yZkaZMvPWn/ZdfyvuX+lBsK4pi1g1h6sVeOAYmA3aeUosx/cfL71tWCKoi08qR
JZxrQqtrSrh1/Kv8pRaZJ8Zz0d/yiT3lCBAagEIe40hTWZu2OvK1QrMzsx57x4BC
F9vaoPWH1e8dkE8Jrh2XSVSp0lk4WF1q6g+MvFdmbK1EimoqBwxH9kalT2SlFtjR
4eeMB7n/XqMSMd15kYcJjVXK+z/GwtrPeRC7qxqcqk3EcLkszqyRoQtcYM3lRt/9
NhA+et/Es1tJl+d4yowmrjmSz6KO8bv/Onf22zKOzS5Jj5GkfO1aA8LSpjXixwP9
IZUGTKCh8qykEX8x8D5y3QG4YtVF7owf0JZye+hEHU69Yi2Iuhmo2OdgM9WW1oos
QhdtrgTezcjxqqgf/nvvNtgxJpzWObH87NzjUezkM8RxjS3pE4Q5Q1P2iTbcxt5b
pJdDBhmn2gHJgBhkYmF+qXiK5x+4jaZgob7lXeidtGIhFQqctZxY1hZ1ZUQGi2+w
j5OBpSZnPtndm+XQzwaI+PKMH/SOHiWB9G2B5OdfN4k20o/hy0lOpmE7s9TOy9AU
Jl1MBkueNHfDrE6jxvd2YK4VBlnjv8yKsMgtxkwr+On1jdpk80JCp5GymgsaJs9x
qgscealXdyABE8I9F3purA15j31MaNLfyoZYRgwEYp9J/A7AKTeXpLv2HmiEdv+U
3jDeo82mq8GExpUIGjwemjKvzm/SRN346FDlr/z919pcmnoMLNr5GegX9uvq13aj
ZO9GUt2GMcffZGPyzrJPSLCHnCafAG6DrilH/QrRqoZPtYQ5AU3ZewL1EvfDb6tZ
6Efi3sTzz3N/6sZATpD0NQmbAEeqJmSAJ2agVN10XJ5lQs/zb82Ocpsd+uxOaM0e
fK08Z2xZB8tTyg7a6o09rtEUT1icT0tfzfNqGyJSiQN1ORWhMht1T9kOn3w8n/yv
KZVvrGialk7YCD+k2XbACclCdAltNuo/fEb5gOh0y8N2zU29O+zTUYMYcRF5s7Pq
dyeBfRrnqRLzeGTTAIjVcAWlgGICkyrDbElIyddFcHJWUXCa+XLD3aEUNEwNZp/a
LPCYHeuCujh06kVkf3A1RI3dpR+jmiTsdLg+hKg7JVpyWWkA6G2DB8OcaW1v2eyC
zuluHCl+XZ1/yFnJqyxz3Z1bEFL2PY5I6alVApqwvNnOh1qsDv8I3omeA2wAcmVc
THGmhRyxo949y9K98A5wLyYWGarRQTU6aJOxAY2+gqFi0u6Y1hqr/IL09m03g79s
DSzuDLW8LZuASM/kIUtu5XrSSkLDPk3qB+6RnCmaTJBcMwVhc1yPnvKpQxi8LPG/
qmFrQUDcTG8hs2wSSSN1H2iM1e1ts+euoJdewD7lgWo23OvNuH9adC8AnnZqsHGA
57pFrqMRLr0I0bNhyg9rQIBcMtCRruwGktj6PX7w0Rwts6gKCi0CZTXymINu0C3s
tdepnjJvzBp7X347epc5KSlFcPMSKTXe3lsT/P1d/NBbhYETywEUU+upx1lK7LcY
/CdMweHgTsjwHVUo3GSXzLHFmQG/WPg3uCNjk9bzoaOpg+9sonzHPsPuAcYUeTH6
4dMnVAZKQEwF+d3oVvqHc+57czDPl8BvndjQgxn5QSBdeFzT8tCvPtrCd/QhEF8v
mw6ocIJXCzF0vOxJfRrZO0O/pP3wZ0hIHLdVI9RGJhsqVEQU1rEjWzsvsaJdrOQ7
CgdWa78hge7GerXnE5eKglAjCup16CuBu/YIXGg+GucEdIZWEEPMuLpzDmm1zT3r
xhE/u/1LCp425PVFgC3R0sijKlNIZv3UlLZrmqnK9gCksXlLC/Bh+UovmzEL1+Dv
NFKplY85Zqcj7fsv+CgC5RS+gRvXdedmDfzGxh5/rbeIp7oqBoAENd8dY41vUKWz
psbVVQpMnPd+3OGmYbLEPon/K1Ua3i6ToHc9bmaib14TfwaSUtJ2DY291ygQ8+Ip
s5k4JX5L8hCDr7zWot8V71GmVArbffCZ0FEWUMDS7XecUmlS62Ytsu5iJ75R8Prb
F7MsYnCTdlavTlVc+hM7v3TQy1VGdQA+Xf/bUYdv3wzM45nVJ7ZQ0JpeUUgdwlaZ
jdM8u+QU+Th7SCwjz9BrvevM6CCI9/BdbE9zIihjqqdQ47rg40/bVVnqytxm6YR3
f9SlTIMeVZgqQjXpcBme0gzz3XuC0cf6OkM2XXhYHk/DNeC0teE3t84w5FiFW+lb
52V3zWNvF/s205M/ua1LdX4SxtD0W9l3bPlDZqJnWwZlo5+XXBdzKJ528G/5zMmn
JykRp08nc97c4ZUmgQkp8zETqc//8VkcFtBuQdjru1a1oJ0vENIcZZyhQ6nycC3T
6RMh9wWxAobXVMQWwqqcKcUjRWugq7Tx3+T1D1aFx15AS6GoHWY3bPl2prG8mjJq
NOosahvdEAS0lFFZowVCemR43x0Uneg2UQVZpc8A/vK8wFuG5z4CJjMAOHJl4bEo
+yqYHTs7t0a+840KaZ+/ffnf+n5uv004LAeCPKWNqtaR//2uSeuejfdxKakC1U6v
RzTV5Z6A8j5wAFI0kAmKJybLY3wraVX7+hvmQunmybpj/aIwvdEqSqnTG62cOP6H
ser5lXGkL5jiYtBqXuMegt6gh7OYyS8esk0GHtVwH2Wq7JtgwDM4bSlxL321jT9U
xT4QRxAj3jOyg2rDoYQ2Yu4YFSpY4eld13ea6B8hBVOYMZUacMq1e9bdoz2RX+Mm
e7r9bOEEDx34wEYv52bPQnz+rYQw1qz++Sa//1YBwhDcCxzayhsznpU9j9xlw1n1
LrmYC/4C2liXUXb44K3aaZvNvrdsfNY//YoJXq6nKLwHlecWDpp9D7JJOflA5ulW
g+bDrDFDOP087gFpWAt4boF8UdtuEer+RTa/6jXKDOHP46L9SmaeINQg+8H5qQQL
i+6ioqOOduzJkQYCbu8HprOF8019BPBpc+dIWukuOfLForsPwcCXZniRyhXKMsRL
d/Kihkhu8r5L2k0rgwD5IirIxwHf3lsnrMCujA763nEreI04smPjsM5zwEDGsgzq
S9G+fIqdUm1+UQZ3BhCQXby2RQ3XAysHNGWFH7OFrJU+ErIDXKveC1eS5slIqAWu
x6nzv+ovrB6BghwHGAd7iHOqWwLvtqh/GOe1qPUzxSzi+dlfI42Z4HtRc8jLDTwa
Hf7BGkXLsMrKXeu1NK2jTFN/+mPNYrQELGeS6hFfs8GR7Qrf+pFKbQC4jurkK2Ug
1Bx+vqk5V5H5k2KOI2bs7VJyvOpvR3MNlvmsvePkd4HRgyICahH3GRpc3myhLrtZ
UjSBWqlkWG5gca8KSRCVd+CAABlzZ/GgU7w3OCHZlGmRGtgbp67d12RGBXlGlbPd
6jGbNW4ams1+gUoDYuuCgQtsbc7djFsI4TcbItaWuT0e1rv3hYvQ1wwoOCoxlgxS
yYbFWRSbiQoNqSS6y5O852ll3GhBb9ShjJ/3dHkpegcEJn5Bt0/e4NgBIKeeM3zM
oqRKHkeCrInUR4rnE8qNWjpTE2j/Jd2Snx+cRfEyg9HbtucHQxvYaaSirSuTvGSR
dDeCf7lNgeofYUdi85yLfrhy5mOqTPxjzoaRcxEoDEBIvzbwdglGVqf2crbCvDLG
QdddpSMoilGaL4I2nGGiWi96B2NeRT2cBcAwReClNLxfuiy8beMlm56luZnzBVB2
Vuc/A8S9WILgfZNWPsaLsT8DVQUfVY+Blhioo9aJu9hCOERj39ckuZ4O6f9GoOKH
V87Gyu6FlwhkxxdnsHi+UDE33wM4KtLl7UBIkb/rjkspinoKXhoHm9/+T7y3oknl
9hb35saPVNTs6gzeFc775vmq9Wl8I41G9i1SLf/ou4g5tnw7fYWkAH/mtZvGCwu1
1auQvLyVr4kYKFA0jUB09EMuTlkjBPgMEbkbmpPTtO1Dqht15ivfNyh+h+Uqs79Q
DWF9DD5DOVKayLDs11gzcxajNe8VdfrTfOQotZ3rQedugBuUZM27vLxVUTsdZeRj
AMSQ6mOYwBXynxveviDREeCaswlwsMwctrclDEbUVC5K/P5UnVY8dJ8ITCHNVmxf
7nJxLddqmsDOjwsw6ZfNwS5NRHUn9zEh0T9pzwgk54XXOm25KWRBUh23E6C2yB1R
OZySHxbd76/7HFq3yrMZ5sllGSgPQbrs08gm5jiYe+6taCZxAGt1HaYe/lQ0s8Pe
iCaayxF3v71aelUXplinB3pwuzYcjglkIzYYUfe7Odm/rMLf9zd458EKYJakC01I
wRJN5/nT4Xu9hdnpK/8oVbOAnb3yEcDuYiOBD04biyIjxxAsPb8geQKxoAG5MaSi
b+H4RhWZORoFxjRB6xSTvXrQl5jnni2guv438RleuPkadcjpucXD+5zz19F5BMvd
KtUOyFdh/2JGAQHYBko/uunLVFHEUwIL7QFOOlS1bdVsosxgt7pUu8IiWUrVU73H
bd0wNzuGs1pM84spRECf3rLSSXGDBxfmz/W43MRXvG1IKnFL9eSa7yQiqerWoieI
3apDSvUfO19LXRJ53pUsEmd9aZ1tL0vcmu0jul5WfWtWV/9r5P898MNoCfIrjubl
QlNSDM1fE9/IbAlGos9/fRLWeWwSjTPLgaSzo/jzDtCMhe9koplmV4f+4mZXdMLa
tOrjfXwyE856Oi5Pl5uNMTQ3dBUeHsT66wecIugW6eKK/9mgdJE6adBUmXlR6BAb
K18vuDjRi/7pLKK4SAz8BQ9nP/+A7sVlV7HXFg9K3Lng2hLMXM8d9SmvuF6s8qSM
SHgNIvZ+lBWJXPNBBqTghluj575egXud20oGiDUXm+Zd7KF3wLWuadYyc2r5G3zS
UxyqfCqnO5cF2BEChtUwCTfrD+5gstDTgVWGdJAcitVPX5rsivgwEF4LuBO2lxFa
myc/tamNN3LGPw8Nvc0txRZMId4Om9lmzrcDeBrfynFtbobA5xr8KLj4lOynMhZd
5I8amEv+LZXvT5oRrCzNeRv0HFmoFzEPh7R4E41iaY/rmM8ab10yodKrMW0aOCIv
QZcdYYE+WpNZbqkw1PEqcIyBS/NWRiH/OJ8wTmuwDu/WRJu2BT2iGlUykVsIwtkC
pTcPzg7KUZfb2hvWer0yLvqggxx5M8xq+wgh4fe1GPcFHvLDpxUUW4jtgDRmDJj5
3cRSOQxCWrph2Ckpqo2StmgZoqP7GtdPfbeab/H1VgKOdwHz90qKTd/pKNdAIekC
NQA6m0b18mI4g4dp3wE6m4GNGM0dCx0IlPDjDtiU1+aud3c4L/iJ0Mlp1W38WNzE
pMzaYblF0bUzovgdpz5kB2BzUiFbcwIzphpLWmHDgqZskhzxaeIaM1LP9aSSOI4T
6f8Q+wm76h9/dh9bg2ZoK5azpVSQMF7nxrT3fdkgWY4Fy4h9hoJAYfczRMnQjjlG
++olLui0dbo8gHtuFJi3ThYUgzAlzgj1fm0vrDHWpEsmXTPGguKnlwVEI6ADzdKK
maQIf5osJ+YTCjxDvG8fdfu6tkvAMfiKXMRfT1Vp8cU7IGHmZpf89ohWVvWBAqDf
ThTVvUbslMQ3KlGF24cacT2MxOH3Hci8+T+1rKRVyrmzDLsVrgId109mRTXi4mr/
cAU0yBWWTkgRxw4cPKHBqq+I+5/VLQG2YJxA/7bRgwQcU0yrrspZgN1oH9AX0Nly
+eaQn0PzoKn84vEpppeLnwuxVWjh5NkzCAEjE+nSnvor+zEuoqktkww+yHZjp0qp
oOPhKlrQwd2VnivJaqw9ubt0e5lbXy2SMK4/HlBvv+L7d9m/jQ4PcztuUHexF5OW
pzH82qSlf/cLkZ/MPljhKXRzUu91QC0Tf81oBztwBFJPwlOhelMcaHGfjg4CbSYO
p0VU081KCyOqSCq93SdIBIeTdqAF7Iqf/c7EBVf20LFgdf63oYA6xvG6donEBWpx
yI8P7+V8+lLFmFT+7y5Uq+7f38LVIQecWk/JRecBAZdQCXtcU6vF9WKabbl2IRAp
N/bCGr62sU2GvbewURsutsw8vz+R8k6vACxH0sSJTfTgQf0qZaE4zho2h8CyRVcN
2nZatobZ3EtpEakfHXXTa3/e2dggKDknV9WrBt1lb74pSN/rfaUvr0up5AMi235f
hU+v2CQsuaBsCuiKERa3v3gSBiSIiDmIOEv7pq515SEsUX9LQpOh9hCsAvXziNs5
Dzdrxt9VbsjIOFujEh75sUUEHT1RWW1vzGxeB3fssWnpHmlwvyv0IZ1rp/Ogyvl0
K4fIIyGUEXVSlsLbUMS2lVxnkSgZlVU3EplRMsc3+qV8nye0I1N8km6vqgLOuUDF
qzZneZXnA4khCRLVQ44AUjUmGNhsMf/+2/6DbWxrr3Ki3MEyVe0qppxuO+JRPHa3
PTx8SHcxW/teXA43JMREvHXoXPu+A2bHFgaJoq7a/j0g2W5rfOM00REQMxepzR8Y
gsuoSvGJQEMJUBknxYuG/xbJUrXCEFOlrexbwxc7NkQVshhb0eiD9GUaoqYX1H15
nZZJlHoMd5fh+egAcy4rkKuEFNjBRQUXrWv4EoWZpVTNnXn7FkZJzGmGuJpNrrP6
AB8H9fSKT78eFJzsJGmlIZxkE87/9SBTS8GYS8Gv6U6muqRvnsoqS5+G1OAdnvyN
c9kKzLTZxKtwZP/ewWRtkVdsa5NVx/wG7CQ9ai+DAZLT8SVlr2gFcvJO9ov7ZYZ/
BTqyD7mtw/Db6trgOFEZ6tB1xfTyJ8UCnRQlShAjG3GcGA0OKsOQXm+T1mhJBkD9
FN4pnhkZO6OxVw1zlmJAeGl9KFUpiuIcy+Z0JFCEwAi4SR9pXz4/IK1ZK+lvFXjV
ioje5dbYE+++NOY02Y1ju+SC04IDvRJl39ugDnCRH+mBnEAKnYMRldXS0cd2uOqX
YWNgTXbJjFVcmySW5FZoTg0t9VJnFGlGiluVn5nFe5Hh29SXzWK7xKRrrNneoDow
lLHjwSkyEC7wwsLXFGqrYLRiPIhiSXiyCqCleWnsBBMTN0sXfDIva5mDD24AzFwk
jXk5eeb4ZTPw1JTZXCvYO1dGMr+xwcQ04obzZ5r6bcgjXxWUnOaowiFvtV3MS0sD
sKn/5nGhy3P+quPwkl1JlvGaDI01px92AN5giYa/lMF7VFFtxVlD4/WlQtRX4gl9
6YLns131e7P//CELai4+VQ7S3fetsOBUtXA+rJLqJegAlZAEwBptN196UxWGacyE
0MSzfgrwus+YoBSVNF6k8I/LFNKmhXVlKs3/eAB4JtCIHeJ1kdbeR0wDchTtUmag
tEV3GvEwhGDbIQrAPZJqZiJmTcaBz9O61NuOiYF96vljtD8Kr6EURPoVxtz8xhPO
teIp0YOVPqcJ2YywPeMRv/mQww2VgIpCciBZguOK0sR8SLpofmfLSTta7Bqb8aLU
yOuMWtdTaJYTS2pHyVWRP0uUxn9tverqwKEdSNitdQZSbhC5cAaXHBUrwan/MG/U
bOrnNglG/VYfm1QECmKk2jQBA4g1oCDI2a+hDKvv8S54qpCISURHl/L8xEQObsLg
Xa88E9RtzvXqofSx8LxwL4R7vzaROkGL4nK+RttUm7jv1bV+cg6coQcvxsVBvtae
CrAV5i2Ojaj4kXjWPTHgkwIZ3AAr1+bbHgF9CaZFBOM6FHOBSCKM6iwJsTVOq6/U
Pxx59dvgMBB27myeJWM/SC6EnqYActLnYVBuADnrkpjtp1GhQN2bOTZgFu7S22KW
7PHi+71NekTjhi2VM5Vkj5YmroiPPgkOD/NaNQSh9ucGEwlLBf/pa9p2nPx4uIHF
QmrwuXNsMA61y6X8SADi+nYI6UA6o7ASiXoKKrKfzm4ebN2pkkQ6pP92Jej6KgjC
nkdtSYicoqEXScUgdwHbwfNpbOm5CmIVzYpLNufKIsxsdz6IO6EetjjP5oyvBbJi
s5bJdeo9KLF60OQONaaSXpCr6jjxmJhMLWgG11LTCpL0L/zNOE1vGndxgM2jd3Uv
Jr59aZlws0Yl/QZxXTnVwjFhufnuIPUuCMyL/xUhFiqrSLO3jEEYeK4D1NHskbGT
a88g1eXwVIKEg56oBmD3fVpDchwfYpWOcWYsuJtD8R6ZN0xFzikh1KBMu+NbUqTf
CKcggFuXDkyl2QZ9WUUYaH6R3WJef7rG5HlgOxIyiTH24sGpeQtdiyoiVexL7WXH
UB5wVCUqVS8WHyjwcC1/KfbKdBVMlwI4cGFfM2LFXUXO4QeS2APCDUaHLt9fxiEU
gZTYcpijaz3MCmHApbGSWeQLyLAEFQGSLHB1oiAGgkKulBU+IQpM2kqLbOfCmf7z
HT+QjxLvpT9M5egrCFUBSVDLFr6+uD2C6OsQWKgAka2OnE8vFdqvr+cRsiRl+sp6
uHFj0IfbHU9K4n42YPV70uq/oB8dehKkos0XNUkfc1MY4uovqGZ5Z9HexrW2fByO
XTpJGE3kfmQDD1sPrrgtGNKcgBZYwYXFiFoLAdy0nCEd4V3sfdFIwbj/MM52PVr0
NK0R0Fr4oqPHSE6FHHq4CkheX+RysjDe813R10/Rzs84aUJcWypFYHxpddWA5cro
hrCxx5tPLZakoVd8/OmCG3e25MM/iVr7L2T5bC/Lys0FrEkhCfLWxk7IgjLd7fGJ
KbInnnqukVZ074sTq8nSKLsNGFjmthu92AouFwgjt9nvKjEZmOC02m/9JL9ac18P
pGvQuQ6ZRmHx+M8t6gk7PxJ4nDN+oen6jFG4acy9/iUrH/IioFRbMFIkrQhQp2+O
PxfBu6YAiNB0Jb7LANXBGki/Utj+NgyTDLfcag/a034R/gDhp0alXP2mgdU+NF/g
Y4zZ1JatWIFQMiXc5BVo45tP/lWKW0I/5WVRMcOU+whmVubf/VPnUfH4tQALWFhl
Vpu2zthBo6JpaVbQ7IIOLkNf29Y3cd2XdPD42CLEOWM7Vx8jvVdzltHmc6iFy5Lx
jVURp9zysJeh5HpKMW0TsWWOlJ7AhuG8ivaTth6qtZSADVCSkKg7eay7xvC5bxco
f5sqPIvkp7hqvLbwTmdhIjsVBKdGxNTA3xt7KGcMWb088cXAcVbOocsdRXaEuz12
xOon9wCq79nUHLuZitLQlgmON3eayubUKCVqytH5Gr1kyU3DxXfTdQwk9qTQXDSz
5Mg9mOd3+kT6kxroWUAwswvOCXFzDtEWHAO2gsrtUw2vNNnFyiBFSkrCovNu0tgW
AdHSotA6lfZhWaNaaVysG1VVKAYuaXkom2UR9Y/3vXhstUr+dds0yt3PWbCn15eZ
AO4p7bm6eb2dHtQZ7c6EsMePLwCM2Ee6R730bCoi7utsDfC77xDVHjqReyrX/Xwg
gArq5nchj+T5dkzpRzuCY6OtB8ncAbQ/p3y6nk8kXkzNNjN2RNOkcEmQkC/BMGgH
7/ltsCyxcO2Ii+nPCak1Ax3XIqAhw+m07+w7xtaQ+uWyEAhHGyfHh6zsAKCkEuhj
AY4k8N5GKyDj6YzYpJY+HPWumHq5LzA0VIfYgUbgo9nf48O+9QKSmL4sK13WX+/E
9sWj2WU801rL4WVlbN5YnCb23yZOD9Pw4BsxgrQEk/8cZQmKEpizcOebNDF4wXmx
N2bXp4bpjGHq4EuJ50UvxI5sXF1KGsnt51lqsuQ5xwHzSrEfaoayCcBx9y0eJQT6
zk4SBkm882hpu6Ypvjkgmw+szjKx6g/qaY5h2nbqwKBamJ0n1SlnsuWtI5kmO8/g
nB0AoQEpxaAMbyuylWFQJAk4YE34ZhlTYX0IHuV4fLIA3A2aLtaqsYaGZ8PbWpKW
wf3AaIiLy3Zhj6dBYnbOLxES0ZEJnj08pG4CvKGw1k3vE4yMLdWoKzdLtzb5JQ5t
2dMOyubCZYv+G74WRdbYLlnAUEj5EYwL82OxT6mVY6raBiuLHQ0XoHqFJ9e8wJ7k
2m2oV5is8DrsGkg/VrNv+x9sSuHJxNRaPO8hy2pSo6cy1Fbh6WZ6ygLMFsNKieM6
0iY4dx8bfa7QeqTj7vzWLNv2S9ArLxhi77CO720ymV6sMwojC3tkrQGn0E7TZwYU
LDIrBzViLriIj6hitESgKGw/RmVgfhJuVEfkQIhYa/27Cfl3IikPSqGGizJcZbk5
0okuV5YbhRp07Eqi/IjXAYYCSDsjERvgzY0j59wvA1wTt71M56ept5rZbudMeeWI
g4iuwjYhBqbnhno0N7mB2UKDd50bJeAYVzsRF5iHHMqukZWgohsiPQ6xKwc3N4BT
RqzlCyED9CAfb8Gpc+B6RTx6irOic9XAWH6PelPTdyYH/j4clT6C2lY720wMRoC/
RhuSOezhpwKPCzbKJiOeZ+lAinjRuz+f6SSUbpKALiy4gpB/lNXp5ozu3K2zLjMp
Dk7GWNV+BrLlTuE0a2QG2RDcdkb4r5qNBDGEvDJAeThvfM9yNQpKsNWAyPhuj0A0
EBgm+eX8jCpt12S8imDtz4iTGZgtPLK4IWR4bOXB4WIzsC7RhbwZJERjznpub1hf
3za8tN5FZ/cY4iV3mQzjv/VA/lSDl/voiOH5Zov9Suliw/GJpkpcGghseqZM6lBx
Cq8j7tSiwDCj5+52gAfCJ46xNwdqyiG8qmN8zoFF0e668QD4t7ufafWszIKYac5k
m0JfBLChp9aKuWYckmt88CUEcIP0QvP9gpi6Ief25Vd9sYHjrhoL3kguX6yPPqJL
pYBhigLIejuEbGefEOl+T+0y+SocWdFiILkRktb5BldmOnL36EAcAhTanYvQUPki
il2O52vOTSsQnfx/N1CxAXxiE5i10dE2mO/4cCNya0Pl4nYON/UaABumgjo5b+oH
GyBJkHxYzYOV1i2I7Y+YF64FF5ytDSzvWaK1CbFeoz8z9TRpw/XvhFZ8JReHimOf
R4zTfJGwLGBbGzgDw+8hq4c+CVsS/qj/sIlqvTPtEBHnmc5qMoaqMlC20xd61/Uu
BhZfIB0JUEjRJpdxNRq529oenpHoaz0vStF4tIr4aMarWpZ+oLOfdNkq0ea4Hizh
xsd3g609M0nk+fiLy86X1w08gOqY/3TT5ioNIU5GPeRLJhRaUUPhGK/ajsVP9NQ5
hCb5lq4P7Y+cCjujQk6y+bW4PtpZbMJYYy3nq09B6I3H/OykC+S5aIDRADnkzFP0
5Yc/mYPG1pv1j7dtECSlCgNP+cemTTTL7EWlUzdO6b02dKGTV9d54GHtu7LffNn8
wwHPvoWLg9wNQITSydkzkxxnr86p2tPXN32Gtb7+ieLtTprsTYG6PGJk+JVQQ+vl
AiI3UAC7aOcH3WVuJJMBKpJYv+ewDfbUhkNsNctD5lOow7Yr//Vs6dRFGO4TSn8f
U494xPZJicPXozrHfZOintSjkzukZvBK7dqbO4T/Q70CvdSbDN89l0LlPqeVxita
kgwBdSuuYCMioYPeti3mIjfH+mB9Y7YvocxOrRlrEQ86ilnJ355qqsmOHeOWDirn
/LpbZ9i8EiGSD8JBZkp9PbdPo//SmX6DZxSl83N9jFHqll0gnETniyM3CyHjCPvP
rzTK/oe3i5hM18UwvyDclbNfIzMIjt8SHqVm/+WgaUILD/RW06S07kIGWYpmwWem
P7e2pAxyESPS64yrpXoW8CYvmHqCUeNwwCdRoYVBtNn2Txzhycb3DBMBfFoaN62L
LlsGi8NwUdQppi/4qf6lNy4k2ghsbCrq/sIf57VSFSDUwYfqrrMFDgKfPUGXyWYP
w7oHCYXdd1FUhrKQEnvAtYLgtziq8SuR/fG3khYP0cc5lhTZfiP0yC76mGmQSXg6
DPLRkzNiVDlcq0JXT+fWK0Jb6OoQTZ/mKdKtWMkjbI2sp8VwfmpZsOVuNxHNRXrA
FFELIZ/K97ubKvKXhEMbFyaB9BRIzdy7XG9iFWz1YwMgDVzgVzW86ZJf2Lwo/G0X
iud/2qUZd0gcFiPNyr/apyWNVXa1AbsxvUJq1IdatNRvkWRdAizpH/ItpqyMy7ui
RgrveifYcYytXycCKCvTG6hbo0Z+o+SZMkW4aJtXnKPyAr4mBewJHOerqQLgbJM6
uEc0HBshzjhEDrmh1Y/bSG7bF6EJugHDtmSAWRaRbrtTltYixJtj7LLC25VZFyG2
qHv36F5sYmAcX7xYi3D9nwycQFDpuctPJDTOggW8wcV4MFKp8uoe7kPTGWYiFxAF
t778i6k0ravlxtLPgk1K/AaYBtPd+l3B2YbCqoaR3lpGK4wkzdRhVSCYjW7nzAIE
Fw+82rO1foIUezH+46jEU6LerNnyyaO4DHxunAnUT0RukSrEO4VgHXkSVsVqiTgG
8h08u3aAW6WZnEThV+TeP2TqWO119NgrLMlSvK7ffH2DvIPjk/+ha+py+bkM0jyi
zdKRLzEhNrNduv/jpt0DaeLIjpv4Q+g6BZAjMt8iXLPN7A5B2SGaOr6wd6NUVn7R
3yzh3xEBqFJkrdw9n70/3qyvMZXyq/yOAxP9U9sXbcrDe2Wk/XTA0wcDuoOgqwqF
X+oDx0mwupSV2bCbnCUtHh0DTJb9qXse+qTBHt8PUk3XR+d3TeAxD0UMefzjYfJK
1I5lL2B5RpxZR7QVnAZaaYWUYB9CwCIbJVTzf1pVGMgjj7TSxOYC2IEwuZ4eWFI1
Cq48VurR8Rxx5NLvHjxBQGFllWvakwaPQv0COMk/QimyNmMwFkwMIh2p6KTjTEwC
3fOFB7kgs7j54J9OBaChnOyR5COvA0huKo0+3v1mHWk5IEKEaqUwn5ZOXatTfhtW
eVQk3JN705FTAlPu6/mcvPzGhyl0m81ekULL/HnoL8CFJJ/9cyKWwf+RQF1YFkXC
L8e3XyguevoRbdVE5eQs4aictJ/OactwduHy/t9ItZ7Vx+ZjcH8wvnCDVBXkRrh6
VMcw9NrUDkuiEAiHAtUtz2RimQtxNwNYCsye/cZc6zuKCWIM5rkpSMtFPrKnveuX
bOXS7lfKghiVtaKdGpQm5F5JQNEdkkefWgrNoxbPgNrdhkH+Ml/mBHzCTnIk2pDn
isBR975na8sh+1oIK+j/O20+Ul6AcJ4qEaPEnopqu0aVcSdeemMdtLdcy0ouLgvF
3GEC5/kcrsiMv+7239k04PgyABxKNv8INTXWKljL1qtN8dGgh5/aiXF/alhrn1uM
SQxQ8rAC2p3i987W7Ba/px6HManUu2b2av4uCVC1mp+EVsKzoFTN4emI3kxMHv5s
28NX12+Oz4hhnsgERLoEhD91D8/V2UBl/BOahrhnbKwu8v2Y+XTRsJ0ezh3c1gNh
w+SX+TRzABZFdH8wESux4IN8iFb3fEOIy9FmZQvg9v0zFxtlQFpqdxZzX5M9I3LC
6n1GNhsESjAVqQVYMPTeQVFoIMON58z41Q3jSuZHbqbD4l6vUBsie8Ba/qPKYx1A
ykh38rEkvnnXdAs8toEpYLiIxQVshO4Mhu4OVSx5/EbwBWZxuo6lPxHm83kL1ubu
4P8DLdSSkatYqsFGupcLiRYZdmzDi+RPwkpk1OJBFuBkSxUDfwBF5QtlJrrZ4awA
R5ROaqKby948HjfVpqqnQMArB3Zj3Zv4D/ojTu/9Qu0Sp5/BksJknEkTFFdj9ETH
ASbst5wcZQUmGyJoyGrZHFr+sx36CCGTelzKTUoH6J1qK8yC0jDedftT8n01sSJN
5UTz1S4LlfS4JVLWNWrwhhQIFj2xg5/nd+f0b0qBcR215yS8W5ubkdoJ7yeBsILJ
nuoENutPnaQdPf2bN500eMgDIPaVTQNtsh8UOAg9/dVE1z9zWD0syq2tLaveSpmQ
UZapFTnFecJ4FEp1Se+LCSFpiHuH6lLA1c7wrnI1KYOQAxdUDi6K3DrdHlSIcj8N
iwW6EBBd25JH+v2ACzKPvpfbvCD1a5eFUIovutBdTcKOFqT7+a0QIzoBJBwjfJXm
Bl9ihLlPOdirznW8+uJ/c9l3EX+1U2iQKzf4PXDe7u1AlpI5FDG8UMfpEP43pbRF
0CxxTzstzVKJ+wcAMRJL2c3BCl4VoMMgW3zxJy68MxV1qZBFXGx7bghXZbNIMOzc
nZs57NSWY5jJ4gblPNvbViRZLg/j1SC60m8/uk3pohsLQq7fqJ3IukD1rIyLsGu3
dMUD4eH+/N/QKD6/g5xxnzkilTHxeJ8hrlSPmvQcf8jGgXLmaztZX0VbzQ3tX/zN
ksygXvIowzRhjX9RpE2bKgDWmTXDhHbPH4D/Q7vOARC0kqbHolE8ck3uJhsrc2aH
muLkoAi0hTYfYxVggwzQ5gvdSHCod8Fctf/yxJ3RnPmUPvp20RMRPt6erO5AhJ0H
FgLxcToAdAx7PDxQWIMxMJifOpfgrbKke8br/pc1MlU/McN7QWhcwhLYFDPSgCdn
AdK+RCrfSrnbKEjropln4npP/8uY4cYmELqnKbZfyW2DOLxuRQbtSj+kAKHHTe+M
VPQ6TWBirJN3NxUD9cHGnv2RuHeTX7qFOsbvfs3j8TMP5b6hmoA6oWLo9PgkbBAd
5vPB9Mcn4RkggxJCve7izB/QTq+KQnREbWOQR4oTw4mzUjEyqceu4kMYlAU8lWrM
Nd+oNes6/mgSP9LKUcdHp1rT0BYkGwQ4fgtAOW/rgIFT1kYdVdqK56K2Y3FtycQk
UWGRTZBeeiHWdVzLCDvUikmPTaiJyZpRqxAzw+xwVYtU8ZDw524T1SJ7uZxWMU7E
7ZiOah00yMp6RbLfm/4ej+fAti78RPkjxVwClr1qxpbFigZe08/GG0DevjB8Cgpw
np5zq2bk1RQEhrF5RFNzJ1K3JU+7EIjxHN4ptCyNHRMizzWY2/JdPixE7E1kTFje
l9qBdvpFF4FrnYbtzisyx/k2EzN0kIKAgRFVXC0R5sFqXHuQ8Rc0y0S5nmWdLKun
RLwlizf6QZq0gfTVXR4P3YuHgv+efLBw0vhOEOKvyOa8nAXiPmBXOJGOjKZWqoRO
cjsNRCGqIngZ/MgTxqhj7YiH3OEUiIsjo3moOkKDl/8kYQm8tmZClkxuLjCPQz0r
VYvoepv1m9x1vM01SIdc2/nNFH0X/9QC8PbcAMbPrlJmjsX6zP4e/oh7bOJbsKfG
XTgdzjESewZdjASdpVOImp1yh9SjAj10VmKVKzeOG5Rf2Yp5r7ZWVMs5i0fhuVLe
4oB16iRZkVu0nL1cQX9t5BS2mnAeZ10TPcfbHvOLhZFCNo0lModxP2WoTaUlGt5Y
31VDbDemhUFja53Esh6ZoUsJAUtpyXLg/zwKAhPyEnzlP9HfAUD105rN7Xrpf1QW
B3tR3KHbTl47puAlpVOG47JmwyBIjnQ7n/gQyGRxdevIeXwlOCKBoRh5jSZCod5M
A7guuT/bSZ6oyL0+ReLbPO8oNV9akhsyZknXLmKvKkdXkOfTNaRpUMAUaZ7mEKbs
OEHcVqVG6BFe53E1sAvN5VBmRtOXbcQ8yWmshVlIhqh4JQnntu+LLQKhMYchCTV7
6Civox9rGz2P3utNCzWaMxyltMNt1KS4uDq+tEDrlhIAXo3kqaRMgaWQbQZeJNQy
dOrZFFHVA0IGeYTYSaETpDTiwS23AC0vCfjqmr8q1V+onktDxhJYLumIrY9E0pmD
YfYsBt45aGKn5I2Xw677rTNKkopyhcgmaZPPDo5+aP18mALHnpVJcm2hZTsus4v9
J0c1Od0gR8j5hsQJiqvyUMmQ/BZ3tOrfq8GjVhkToUhngkt5aStM8s6ebLRd9O1+
/aeDN41mlUx4vh5tAGcoJR/e2gZa3rfDVRleJEW5PjP4sD2zAU0mVtC3Iqkv886i
6824b0o6i4YCylqXgxv7I8uj3oPymqHa3Ejkqg+alVdv2eTEAmCV3MitygS3okoc
9KWfb9UjSknNURNn/6thFCT+rp3qYbiWA5kqnGhhctlKm+q5Oa2nloujfvCTDf7f
RZ+VL8HZw0Ob47UPLGiwWb36n9X3R4ENeOPXkmSuqjCiWbVRatlMgRq77vXD6zuE
nHj8e3wAXBtOPZhA/nxMuE/tap8a6tnh77W9OXh/ZKTM3ZTVUqP7x/GkbcPya4ZK
X7TdBIv+ZcHV20FKzOp7Nzr0/ESj90RmsGzmGB+l4TmpR4B50t50piNd2atEKPgj
oLUlVnTF9DaSnyrgrNDioql3zU5QX/tUJoS0QhEN/l9Q8chPiONdmgMxb/mOWGr0
aXa9v+l3FpdSBRyt0FfnKhPRJH4wkw/JnOHV02YinEB+kPPTsgvVWUo88+aPoba+
C53eYcUWC9K9X0jwd0NrQccWepntBgbs3nC72d+jkuYZLsTRAKAZ4i21HH3p+NET
PAEu0w5DOgUeRpm8LYQ/VkifCWvz2dgVXl8BXVoayi49nTKYjPIZbecwW5FSNY7Z
86YuOPDufjcMz3DyEGhaGrdqfdO7VcT8+IGSix42JP+4cyCpPeA0NCmddGnceKE3
t766VSNctu1lp32yfzy5EBvegBtLAKRB8KlBR0TFHJKmNiSpcsjlPo9vkXYEiLVs
DFTfxWE03a39JpZlVPXi6Prfhf/B8F1mbCAi2DET6hOo5KVlVWoY7M+c5Z6nN6mq
WlgrU8k+WXeVlFlAXOqqpAw1VnoyietlvLoec55ALiZ5E+TNsjr7mcegm6XrsHvA
uITt4FnymhwlGl7m8N6p33a8EvssBcyIvCJ7L+CyDQzAi5NRNYgAIHmzc1gM1Gu9
fkyBV4BZv7FrMuMwRhFh7asgiL5GCiDHa4gzxgEMnS5eCuG9LuFv75036oV+UL/Y
qNLMAkv4sZpHs2Zuuojd/oxW7mz5kwDUjTj6o+Ex6xiNTxAZ6WQ31YUyALbPNH8Y
FBX6dgefZwIstvtVpTjv/fub+bFq/qD4UW/wbJ2PYZECqX6KaGvuYTvOHJaCQla7
8tlJ+EorXgJYyU9rTGDIe0msHaTxs6W/dAY9zcGwPQ/TmLj1INwKXTvSyJrkEsyo
FQX45iSdTw5lgt8NiwywK+lrTQjPJ/VXsC9uvTAHFMrT4riX6JdoSgQS/mZVK0Cw
39tqole2MIXGObiZMRw7I3x6YHQVgW0tGVwEJZS7soYnIYNVj7tb/tqRDNV8t1GX
nCB2us9wGILQcuZPp2cDw3Ku/QmHnFZhiFF/eZUOFYx6G0wKGTxbi1t+0qQ6pV43
juPiS2uwFLj7BiSpRVUQ/wLjW78A6PAILLpzdAbgwP9LRuEflQLOejNziJ8qlqOk
N8nx/rtrm7QMZtAF5oSJkfyBoOXKkplGObb9Ozw0Ao+/8eJreWMwmEyM17If7/fb
P4Wg7NTtz7XYS0dIQ6UJx13Y4u7QctXmaHLXYDSZ3OS/5+Kb3tbJmf4UtvwGLs0f
nJSs9bjtNixmzC6e5f2GDLnL5Kcw6zWMGVrCCtIoeIExVjXbVbNhdBoYBv2Fr7wz
6qaoGD/YC1/eT8yej43PLgSASnrjLtysEQSi9x03zZwLHp6nahf6jjTYy0b4ahG0
tdF2x/WL6PR7QwTsMH+IF6numF0JyF9BKpqIIeS5TV/lfnMm2jszZJUvW5Q8Hcch
TCh7CUA9uSykO1Gl2mlY3KI47oy6U39Pj+taJrUotpHZX/s4Gg0QqgXaguimNpD4
mU445sHq4CgIYcomXYN9c+n86rEra+8kxH/osyqukc324S0kEcXgSeNjWF2Cz8+N
uCN20EY76rvJnFtTjh+2KGW7JrapLXggiVh6IVPElsWbiFKl3K0uHXUphYHY7wCk
YcjhLZ3RypHRVJisFiZ6MY9t65oES1nu1Fj6S9bvNV3qcCGhCnhw1eCsDYCeHO6Q
U/VgxgV7WD4GPdVktZMMi5MnnzhndZfSkuKi8nxMR7rCwNeq3tMzn2yPvrQdcJQV
7P1p2IK75vMO9gn0n6r+yC/L19HolHEBf3fK5h36nDAXmz3gdLM22Xh+zDh+GB45
tE+lSSiFkUFj9X+7OzD0SQ9A1gcc7Q+RZD1u0NuV1hJs055c1XTHgFMLqg250+Hd
vucmHDpVeyhqZ16/UEwgf+9D6d+sDFGycLRKBR48YgEXMlLR73erNVhFmfs/Q9vZ
A6bHiIEEqUCHMQMOizSv1GvbVnH3wTjzQuRhLVDbz8PdnSTDcPvqSMkhSG/2j6QV
DTbgVFVQFRxHgI3i2pCfqphnc5M0X8zHIVYHTnLvoIGPsKkmCdzVhl9CYsI4nZoX
0em/scrtImY2QRyuTh9hu4qI9neW2BsrJkMNJCu6Hw2qbCHayaruDNWqX/bGwz1A
FaDPbJqzFfUGb9mX4Umbvx0/Jz9xEA04s4dMsugwNeWsFPoa9ZJjoY8nWuTZrAz8
2fLzT3AicpUQ17BIvjTvcdew2m2fRMJCDiGI97eSxEZYPW2k2QmMbFCpm872t/cU
FTqOk/XYqxeIEt2cMwldUzWknM6cR7PzUo8EdQQwTB2uJWwlqetXskDrWkIWUloS
+UKrMw1alOVJ5YFwCew8YQRJbem/1OjdxVDN72xHZzIHOlsSXejWFsB9/8JCqf1P
f6rV1EMQt/JpjVOLpWGklq9lQB03Sgs984SD83RaoQTdDZCFXVCgTa6vTn7VQLF5
kLbGYMxsWQ/VDhN+Z+OmnNBIw46XWY9nV1cbQCmmVw8FjhEDf7N5i93rjcAh5M+D
Wx/dnyBgArZYlumykMUBWhpgsqyZoVMiJ8F9HP9OlIZZMwcmEUZOEtZxMr5Ek8Bc
sKF8VSWEMtvlzUfRnZZScNxr2IQjYUk+RpVWH/6r+RquNOtM0/AAUCI6pkg32kD/
PyKWRS1X/50tmo9fcjg013jymGyhavhZEL8DjVmdzqYy+zDVmS0nxeNCiV8Q3wTE
yKOF8reG5QKxvRJMTaVGiVzINAo6D0CDSANDYpj7Kv61WavEf0P5Npl7J0CgGmTV
idWFEbHO2PYFD3xCUbvNeYD69gV8M7YXm9OcWe2yJkgO1TVS5uc1nCBzVZqra2Y0
JPRwfI7WQ5aHhLfBVMWq+0j8jcGm+qB3E7nlY8AzpuUpXl2Gd7UfMRTMJQ11Tyus
4c3vSCxU44qRbjvRrKVaGK8MN3w6HgkST97gsGRYqtA9SaeLYOcO2zojkGx3y5Qz
yETewf8f1gzCJ2mJoco/kO5YzA44ZkagtjjBSI6XdsgVc7viS3+WEm5/y8KlUddL
rzcnLLIbNJyuSD/FLBPIj248jW5KYoUOS2H2JM4XtbqCoM1NzgwchcHeVQjUMKT4
pHzHxhxZYpjZKznq80I1LH7jio2NBAG5lz2mYZKi19i7sUnqwCc1yTMvlPLeqqLN
2a7ArzKh29X4F0nVGSPcCPgbTU69oybUiN0qsB09cUjRVNlZmAm7tgMi1awgx6qa
W9SOS/N75QX1ILa47pdDDsn0LSDxEdThT0h8us7OLB9HxCpu9sXVG+Zaos4dhwX/
o2gnFHw80ExEZfR/QbyNcZm5qTncQOhD34mjIoVZYI/cEIc0uksoL8AKOoL6sGix
2M4pAWAycDety7BRnqTjWcjg1h+EX2DDP46NAUYQlXyV1EtI2kMGADAv2XrEc9MZ
GpXQ73+NGiKrWwtqLGkcDMLl6WRsyTSzTM2U+wYWRxDPmKkKol8S9QfdZECDAm7y
1ZrzDsx6qJl0vOVx9l4QDJ5rtfn1G+Jyoc4vLL2j4KppkpwLgls1lh0zw69QdezG
nKnEYl9CrTIQ56DW4tQq0iA7wJqcpBgu+SngTeN52L9RVkL0gVyGp9Yc3Zce5meD
sEkeeiTnsm2Ny3HSDioOFJ3098lWfd3uBXO+c4qeMD2IkHrnNi7Bs6+/DVjxE37M
YXYDGmNUkiO8425U1tv/tlPyHW8aiUbkzOIiICmt+7rVsOkZGRvuF30FnXAcZ5lY
ar6DtDCEfeF90T8h9v9QJQFllP10AGEQGfeV4L6UNch1RSpWx26W6ftGFLody2ww
hGnNin7aO9k9Vz20tKVzLxA2cVex7lZI/qql889yMm6iFtQSYCQx3ONZyp4A9YnS
8cTfOeGEgnlUR987xTyxMUrazd9nABkBuHE5J/WRoOh9LMCAqHsuwANmZXBOF1Yh
TIe3iEqJsx17AAVQEH0ow5M/QQCHi2SGMQA1qjacQkoO3AjLWKMjYfb8jcXu2yQe
J6DvwMZssV5HF5Nq7azc4dj5+ov0OIsE4yUB3QOnyLBsmt8o5qJstj2FezdUIt2O
wZiZBua52xF/YbKTmFnWVoSk9mozoUPz7JkTqERceN+Ub7U4V9Z5lHnjO3kpdPeZ
Kw0PRs64FpSVPaMgo2earv8NHoe8qyTDkQgTuV71iEgU0sxRSDosGMPgQRKZ/nXo
zeOBepdnUWeXG9iW3YZRShghNPWJ2GGUfP6OXCm3XPE2G6YjFwwurCS3Dw3pcbOQ
nSsb69aOXRM25yfZEhBOMoN/WYR65SwjCN88Pbq8N8tFyCTgjXJRokzQpNQtlODT
qSnbm2Cjm+nhmPIgROFkRqQIlkBppVz9P4y9EYNrHAzlraTeTncuYe6GlX+RzbRx
/MNsnqRWdIVDejfRYHHm8X93QUTcA5guUIWRs/AlMVDtctQfpWWe48FPeIBkVpcj
WFNb68tQ4kR352giAz72itieitv0uuT0xNoI6LPCqsNf9Pe5yWRtl74DLq/iR31a
8Vy+az7mX/leZSurMRnjvK4h7aExkk59kpClIDuz210qlVnHJBN8kMAMvzx4bM7h
0n3hGnjbEsXfVYXXtQBBVd1zlpwiOLdKZ8m9bD4sD93sR8jnZlOSdOrNLZNjnwaX
8FQnXBYnLwUwu6Pqeg1wtWS7MR0qMwWtEcbbs/SzatemnPRzPwXQzeQtvREE0jN+
eHQP9+vaREOzAM7CLPB48BE2XI/gq2aKDYdeNoNR7T50LHyjP9BgsWJi/9vAAci2
lfyOruxvlIgfyl3Mk8o25AqLreW+pq1zkTm2dEH+9IxkPWqKeAhhMHnIYs4QFx6O
lKp7uInX6uPhaHCsPTaC56vWUKKwejv0WccL2N4KKjlXQxWqO1l6s6SWF30cm//M
CsNRHNTH4O77Q8WfTe+I1IcfReMH5S9NQjQqdf9GT3yPhvebsV9stBCI//Tq79jg
4+mDf7ChjrhWAt6LkO9ZGS/aKn03cFbA4u003gnHoA4Wim64f/kYhNUj41vTcLot
MUYJR9zKlWGGOlp8bOiheoZQL3ZaoBP513+zgztsSzxx1eMk3OnYsSQZQSCinhNh
PjXGOEHm+LRdHDBPL7rmnHsWGHg7Gb7A5lXTjyfhXwr+S9HQ3gU12o6fx1HoWNLK
ula/O6RBxeghzVp9C8V//G1HR2mXo/x+q7YtlVMGy06kfj7t+yEMR3rlXGWdchk7
8HsiqMZVUcbOteyJyhg++7rs+2Lg25OoYutCJgklkOz0GnEIcc9ovBrKemnFFoah
A80PEqpq0vzaZYmHyYusEiYRGArmDQ+Pa0PK+tbmBeqssCT1AJ9g5WkSqHlcM2LA
9G9EyKANBZnr/p5w+NpUYF2Z9Ve+5mRzdT6nzjuGk3ZqiQauydWSfmKPpQdHV7Yn
MFXVGiocZw+altTBfnnsRPOaH8iDmjN4xAb5PWIJD5rKgRd8RvH6vUnj7uUNWse5
xNL9DR5J5qMLH0S9X+CC7rvcnfssEdogzFW5HPhUUjMeoN7C5FGOJVxObzTbI6cA
bhVMyeyCS3yWvPaCCqFNN04WdzE3AEZVs00FEohOA9DkOuSPeXje2tF1T3boQbkJ
q7BjStmkiI3OG1uq0qUYQvjuW+gRQLPNplkQvbRhJ9suVE1JBdwjyztL4+IVohPR
xOzvFRiZDMzv37di3tUR4gTFpooodVqbeN+zMPeGcf+NDMLBUX1/nSmACm72dLWs
d2jH7/2KdWdqjPDNc9NtdxtNDT4Pw9D16605VAb7KM8sdKgYcwJ2DVsgxXBc/AVu
4For3lKNfLIaSxM4c6hVdam50NY5y1hVGWBWRmbu311/UY9GYfj66lnoouTpO1Nx
U3fqmkZx/5jYYtC5cqfZwEk1wHzs5XjeMbmrK70MmC2gjWB99vr5Z77QgYODAUE7
D9p6azhuCCjE6yEyPEqlxj7/V+9S5Mg4p2OYo0I3xfemuyR1WhuSvJeHa6+gmkae
jcyHg//4deiAkCVSkVjyqabWulwsu5ebJvZjTVbairQSU4UVp/xzTqZONGgDffsJ
WrRpT7duPn4NGCQgmvrYR4GyFMpIyisxSymEO33eNxjmxi39lUASIu0WsNP9VkWS
C66WdpdJfzy9+WJFb7sLmRVyFArsXZRipH9lQTbhjYuwPkwMmsx8qqO9byo3ndki
Zo4hic+Kn6hRU9cV2hJfCvaMam8G1Ve9AclMe/lTllup7bLbPcLDvbTZtcuZZE0W
kGuQE2na91JgQc4voR8uzAemlDaw23f++9bWIYozQkKtLzAvnG+orJ93oA3g4Rkq
e9lWpKbqma7VOOGabKGIiZPObghe/d9tPD2/4hYK51XhNk9wSa4sk8c4W/tKGyPi
/PNuOsFmDTm3pU+Hl4++S8YuGzRAKuel0wNdG7968aqgwkM/yLsmkxHUmAf8RhY3
ctvbL9LVefhxFLEMfdl8v+2qgOhp+pJ2xphaqQSjjZbzq+TWaMkg2r2UAihZxYnx
jorb9cLUdpMBbT20i9Y8Kb+3Z77kR4y5NoQF+N5X6amugnxm9QnjYaqGRPu9asUp
pAo61S5xXFbRXd26daZHPTiB0mR05H++8Yw/FBODogZfmcGhSxO6xH6joe18OnD5
Y9PpfA7tmPosL4z82EfFFnXbvT4dFGkXyhUqFuBGrO6sZHpeNUJjGBgz1MRZZOLK
x/tTpNvdU8/sA+ksu06ajLtWs3A2KKuOrcomx7Cekm0DDbfxdnO9R+sZoYSMtTTm
DX/JJ+ZUvnuIPB5Re9z19d7zi7RGY4ytQq142r8a40zAj0lyzafoyJGSh3hBLEr5
2QQNJeVEtr9gMG8NhtHGG6+WCfvqzOEZY32Y0N1RI7ouR1d+JsD5brjaqtHB30fI
T0ar28PeHidUJV3ceAOHCMikoGPilR83L7qa/wcbmV8kGRQB/tMRKhvuipyHWkIz
kGoC6T1eTJGDHbxnuFQFPgrfvxtmosLovX1SmZfZVYoqYgTZpdLjjbhM+x+xD2OK
oezttgH0yplcQhncoRVsMm5MkQKCyrw6+UkfkWvwbhsDtijqozYREvffpnuU1rik
+ukWuz3FvY2NjlqVlCs2+1aCY9YIXmd0IwM3JkTXDim8+sU+RCIDU3pI8kdc/PNJ
xSyUKnGyXIH8j+SDOUReaz3nfSnkWIGOtsS/fF3AifNHvURer09lIh0KGpL4N1r7
aWKeALnKcEJJotdKhGT7kAw4ZkIqQnSIYoKIMbDOlnBMv6lxnIcRrcFTczWa8G5h
k1ITyfhSm/9KZXgi1XaSwnvH1lRpzlq+2+soh5VMlJ0xRsWpUvg6OIMnVB8JFz3y
9uit5wehO+LR1RQMy7KWcuu1PT336oeEiOhX1N7lzyAz89NXKSHbAeBDhYPxL252
L8NDItKX8iCC/8jvw3GTZvw2DZVqSYjAIijZglG1jl1LpOYCUlJrD4Tl6+4sUU0V
UdEIsnT6kutR6ZULHBWgfqcbZ61uRtJHxCLpLw59qgFYJ6VuMLpS+yh5AXoS2jF5
wdQ8RKZB7WBMHn5+c4BGVqkpRcSSghKoiOFd0TEc7iBsY29IEMQ200VQWApX8fVn
5QvpgAdydpRgIYiDRPzJgUQ3/ReP66wPESES9HtrXeAccmA3Z5RxgZHbJQE7vGet
OjV6koMJZ49EWiGCV3iQs78++BicddT+jNfkDdeMPB92UyKVFBrQEMgc8cbjGaSj
djy7hOAJmwBq6D94H+GhQgH2zgeLnHkkmQfVrzX2l+SbaCnfaswLPVdrx1W8M/IJ
RAecgZBFWxsB9Y9484icDsMey8OmA35xK4DIrNmsEyxEh1Q3ak8LWnICB7+wZRUk
opVa9gUzpnfRoAYFYTXsC7Kx3/wzoOlQ36oXV9+chEXU1aw4hjMhy145sIuRZE0X
8AHGoPyfe4+Lxnui0LPjxPpo1tWSVGYQSKCoqfal76Qo2ZzNVUEJJtECJb6SatS8
Xg0YZxyDxjI5dofEo2pGT2lBNj9Y2XAhQeS7+sphiiN6wGinALXM5TGfrlXvaqUX
9mFLF0O0Odi0lwC9gAjWkPQHnMDTA2FUHisTyIL5gxlTSZ6jqvNgyJGdFQhlWyQb
I6lbkSrob/t+A/MT5KEQ8TCelJeRFULpTUOc5lLsFn2BstDpG4Xts03Z7rU+BuZj
aC2wivTAw/eivswQgHT2G15/mc7U3Dg/Cvf4GY28tQwEIjqlhECdl+4LR6Fdc3MC
6tbXOi0S/Y0liuZBR/S/lte6oK/KZPCmnUYCEnILtfBJWF/C98i7BFTWeYdru/7A
0AWbIU/1MlhLTOfUJmCarCMmFuhTfyzmOQ0PJ95SjdLSbfq+sNms0AB/leICig5n
fVPJF9qq6aUIaTyi4uYMXnzKI3NGs9ep7H0qQTIQ/6X+OXU5A042O1wKStEb1s8M
9zyoLBNCo3ANwB2i45cCAKGhcIYtPEa18EoXEDqTmg63hFPNMSYYbhMgtrfRrYnJ
YyHRO1Y3lNPUG4V6m6LuegvG0vcbfv7QjOIz7HkytZIZvquIIKmN+h9c5S8oqZo/
z0/mgNVVQF2Bmz6bjMSftue0rbWZew1OJSHBUaHt3rT0Tg7orDOfo+JU2g8K1aaS
GW9RXL9b247If904bCCulAP6SKjI4w5fe+n+N40dVxQZqyGIf+SbFOLlW9RRnInq
Bwfng/8ED9zrZ5/e/bZw7rpmf0Zea0vYSpMQen9JyPxSPUa/CyX88wSMg8BqWpqr
42i1eZMrlrIDCvjvxEAoGTTKm0524DIL2yfMILNs2tEPWWYwiDPXp4UjE6o9D91K
/nvCaI13tmKsnYOadsO9gXZBcVDYNssG/nQb3Wpk4B/SWICQAg7d0tZZSape/yxC
66RPXGCyvuPd1cWEzTn2AZSyuPl59Lst5owuKHzlo3UoJFklQLYlFnu9bTpzofAW
I31sN6V30N3RcqbK42xjNrGtNeSTjJPtK9POuD0MsBjBsXFdZ9kVK8kUzpmy8KDS
csexkqh/9uHR38BCU0WIslYn/K/wQWpjEEDS2touHDRnleGFi2yRA6Ink6sS/Hu6
fbjGlxcRKQTzTJkCCmyG8sQBgJC9z6X3vTMXw+gP2StE9ph2hU0cemV+2bOLha/a
5H36Q73mjZuFvdXO7HursV6QPNr6YaHAd6jixKerxZzOGCP2hsqqiB5FRRbOaf2h
KvhdzAybK3XTUw0AtXNMo7ENjS16aBOsdEGdK0wlrM9EdsLWpBVvcchuDwzY2VRW
euGPufFA2zVvZStQVyxI4g2mu7gr5BUybiZ/zUj778UzljSLJREC2Pr6AaysgDxK
WyHW2gnbH//a9HiM9YsHkJ1JYemm4mHLDB1hlI4ht7NFEAkcAflP+W/uNf1/nmE8
eAvJCgj+PBXjtPaYNKEtMtVqLH8L3VzH4wN/GtLCog5qEltWQ5CutUYhGcL2y2UH
TKGcQXNGaG1eaUU17F8b7R6N82x77wRGU1/hSRbtd269E576wcF4GM/7hpswjjvo
GvplcWZhJrrQ/WOPu69uwkKKOeeNF1WsyomYXU16Ar+ey2T8BIaNiBmVm+qk5TTT
4DJG0IGmY3zx4cW1J8R2zFuf58/3iHoV1eHZT/qr0pVLtZlfXLS3szhoYjC0H/6j
eJh6oyeVHDld8mxXuNzjadhn0OQdK5FJCPb2Tu90PoPJctLyMLkaMVE8uV5AlY95
E5G1KlfUD29EC+OBnGtS2skMcZuc7hnA8z6WjIxQTsNsIZdfQmWKcqi8hxtEu8zF
c6iF/oBzKngx8timP4C4QoScz99vuKfJoopCyOMqMSGURUpunuG5r49j+ZQJnuzU
u0otUa+IV8W0TQ7Q5V0kulcvD4wMVQPhAglr+rr0T+qscLsCzmEYuJKLc2xM5QWW
i0quiinvxieB4gJYMFBJGDVWj3r6TOvxi8UTWdOQQkRTfCVKpW1kmwzJxRWA7PqV
xbDQwVGSsKjlxbBO0PX3S53km9iker5ISE4Jn+OCZN04omhmJkPYFQ7UC4MBRocf
b6Lm2l4ya05j5GNd+rTiO9IeIQDJOtQZl4c4ARlLfLfGxKVx+gqgrHqvajd8FzQw
eaaLfJi7tF2B4nfRz+ejOLMEr4HaVyFKIpQjcq9MVsqjkpsGm50DbMWBpQ5LKbMA
lwMo2yWQ/bBD2xkso1U1K20zLg3kNhXJ1mQv9lp4jdGQdFnSlqx7p8OwKxlu23R7
MdpbPka+2VvuQBX+ieWsmUqqDsDdfgrsgZgX3NCV/6JbyCDhBx1qWMITDzp7WUX3
7qKfr1nPvq8cIvkwuOIirEeOP0nKuuv57zs4gKVCWvnGpJGkbeVSeaAZjC/yVMnB
rTrgiXEzkYuzBML5436XBEVBe52Oi3yggsQrjpWhp/wFTB5axDt5Unp25Gir3qhg
3+3ceGjeGuqstZNGadiIpdCLGfHNb3UC0XBnqL19c6KT6n2Ces7ecQrAhP9VXS56
dMyokyu4hCpbsIZRaejN22ayGFMTRteu7prHXknCDp5/Aw3da/o8WxFqc4vGYWa4
/KHEN7+KWynn4rPhDhOQSfCUv/+Uwp2Y/JQlawLec6/ABHHU4nBk8jIEa1lKIRp3
ly7X1NyeqTjheAxBSOe7smKKlqX7NZW7qg/E/gEOdt/O+phz4PUTqiNh2b+xJ3qv
tZ0SEvtQfMb5otIAljWSHtMaa/nnGPsUF66NXd4AauCCKoYYGjWYBhIui6RWm6yx
j4jpLIYwhCRwdQIwqJ3F+MPJDQv9/whkUiIGvS/xedkDjB8IgEKCIFxJjTzXrcI3
AMy/X0wtvhjJENVz0IRQzwSuMvi9zYTiiA5Tv0XxqvNTkJTfAptnXxIVG1ckHvxZ
q3OQlBosCQYenrXt6pT/7dU/TXXzLwmhTnyzU9Q7DSugrwsqiETo29Z9qeeM50BI
gS4nlFyBg11HuBtDYDrtyKdctKWB35svmDYqSOn63TK1JW8aGuaOYTS/6oiG1Yrw
SPClxsSKr22ASvZL5YYf5eDu9PADEy2Pz+1aehEL+GGgjTEa3pKR27VP5k0mAhwS
XftzaMjCVkQQ7Bi/O1tg/7j9vdoxJCh6TYrLLKoJgcmaJ19OzP8w2cuc86PAhrF5
8KOZPwYvsmawdDTRzMvXfcLc53KQ+SdgB0KyYEXjnd+PnOyyj0nw0R/TSHNoynZn
HIR3df7OlyVFfHT6L5+xRUn2bEQKDsRjq8irPG7pJWyJDomVc9hA8PA3t3PIqb2C
8VLoSN9oRc+GGQi6ho3gVSREKxO3GdURQ2NChdl3ITWpkQ8Lf2pCluMn9e2nSNAn
yGOBQBlPHnZ3a1EVvz0dPRP7DDymb7IOhPchgmXiPSOlc+use6/ecaOjrF1VOGIS
mgmfeqURhqlNBY+BlXzDS4SjWhi2dmpvyFUCU9wXG2kdw09ZMfEHgBo45VemCJ/T
ROvrFSQCkkD/pnqT0OU63wbT3vnUf2gdGQZwSQY9YiFqItnjq+gH7SIJqrm2F4Z0
b6ixVvYiNj8c9TBpFkB4CxFX7i4aov9vkgCp8mfRu3nSYED3px0juMaMPml/6Okf
axGtejUA0TGjntd0bCq0dvJUoXG7GZOrg6XRIRb/sCija/TFck290CWuPPQq8u5F
KB8t9Gbp6jnvGxvK8m2cRSHlivmsp20pKQjRAuabtda3xq989pvkgttZ64BZELiG
KxIKbppGEbBz6f3/n9J84OJxYL7/MwEvOs0RfHBFJTgTWeeg95PWrY2OwEMVqeYl
uwHaSW1/an/wVHiQ+D0m6+GrBhYQRDK1Rr0L4l3UTHQ5LnuXHuVjZsqCG1a3r5bi
pVxzHU1GasiVGuw8RKNxxcVi3Myfx249kq9oM4K904FvAYHPkS0MfB5pc7lIgfLW
zwwPGPt+vjqVGb5dtJMiIqCHSps3f4sJMDIahCNi83rcrvCsfgg/6FjsD3bDAJEx
gbNPR6w1t4v60vGV3EgY4UmLJTpfR7fPvt7hA9FnTc1B+1zNFpBxXSyGDqaYvb9v
D4hCnA2UF3pN4+fc2iTrRY+fG0wjZfZLgD1Oswwx3Ta7hiGccTUM9d9XnH8Zx+1K
PiNBJ4ZAuQB+d8lqif75JX7k51AK2CTsq6pAkesmSSMriVR5vG1iwcikKw1ArHRF
Ufrqhb9v+IuWhL4lmPwNH/8tbjoSndBVDRpg/JW1lZUYf3aqbMR3OxRtMhcNXDUT
5F5UeqwFViDoBvpVwRdlt7za1n5LuUSVAh88NOWV0fQPKgKGnsjfJZDcPHtuPRro
k/biabXdjZtEnkiVxs/dCYV5hTxYqzNKHcZC3cqvDeFsyCNXSwwhj2LThSmE8PGl
eE+NVt3F58SDN5wT1/3xerQo0MYgUTqGe9Ac+rjCpP1LbnGGQPgJVtOydugCIsy2
O06as3wAyYDG/B061EoN5B/z7E+EpVlcfoDStx7xe1FMYngAN0QvpGVlMPJUGkv4
je2mAagdDkOim7RyTU1iJsYXXtcrpnIdojoXIS8+7k1NMugSGkzMRs0Ox9GDMajC
w2SP+9YmS1A2CLQ9rImBFKrpHWP0r9jOtWb3H0pjHeJWMK10Rl7yXhUyXsb4Ntsm
DyhSDud8n9itU2NAvU35RegEaI6ok2PL/wG3Kz39EZPLxtwmCEKF1AzO6KQxI4Sg
0DXWPa5r0yrtZduA22pfkTqj074Lr909MRIHvwAtaPXJk1+1K9PKRXouON+tR3kt
dhdQ2lNCN8xq2Yb1wIuJbTsk1vo9J6xlsF2njAKIUzaxMwNjVwDWtGtlvd5A5GT4
eh2Sd3OMkJnqT6KytutEG7pjmcgrfbGZBYHgYo5/RElcwqlby5CCfFWjuvIh0iAS
zuDf8yS1x/0ip6M3GhqpORfHqCqmepW+l51Bb9nY9rElpDVrmvdJ5mSLuG2Ht+GZ
QIoVJvAxn5koA4E891jPkdefvt5M+58zO8k8oPZx683BjzK4Zidi+e0XS7QIfkrs
yr65UdmQnpPhqOrhWuKu1PEhraMVOoAb/eotOa89XSQYgHY8XA1z4JuuPkSmZjXA
4HxaCqulW04z4yaOHUa5owLjvXg5jE0QJ6ky4lzdaADU6/FJFqn/5/esuiFfFzwh
wcbJcFiV0Xj7DQe/xhnpWA40Mafde9MvMJ6igmlzLUTKRuKYMXqbQHlncV66EK/3
u8e/xAge5hIavzjil7rErPU+dBJoTUYhVUARMZV7J3a2AiEd7gTeXEvzyQK2j7T6
pf0TKhZ532T4hwnjLTo1p7jCAaO4j1L5yOIfheOyx9zlxFmQdKfkjbl+jkuydn04
zOgCEYm8IvKACG15nJb2OxFQ3fEqBHY5CWosQ6KmiR6aL7pM8hWfbDrL5vmcJHkA
as0c4nJ1f8Yw8qBzNtWo0pszI3y+Z5GEVPaDBXWyJYnvV2S8gIHiDZ5oZxzleDyy
VaTU8rNemyJbsL3W1gnLqIJ+BWmGM+fH3S0vS4p34S+yK2Izc/XuuBOV4ur8C+7z
qQcO/AEozdyGkWdCoKzhYsKqFpH2gs3Mf8ZRxHG4B7yTWWIfuowPPPpQfmhl69Me
26EvHHhU+qtTyDyEJW2AAD7lXVPbtXRj0lt12Juk4va/Xbj0f0TqtM5jycgbpdJo
DnS60+T5J5pYLK0C/tzJfyHQ0mpZJ2z5O0MAdsQW4z7muzwcnNqjGKOoSAKZbSJv
Zmn7lLtW2XxB/bxcwtcv9dAIYULxgP7LKJqV+s++3HX6oJYWiHLABgLkrMa+UgyC
YfN3SiQ8vdjuG3Wt13itm+InSFVPhzfAPqQxwqoMe17cxmDbI9fH2mP9d32z5oEk
RtZj7ssimEK379wLuFTqZP5Jr0KJ0lsZkPn1VpxslvRfFiSDGmLsQ0GWkysR2a19
I5UcF9ETMeJaKsj6fcmhKVEnZpRcGKQvD1XF/WNnF0f6WfBFBn5RrEwu5pbQZHkg
I2BNTNDpOB7+duY+JBz0mnWKLB90euba4izQ5Ug5NpQLLYdtFoq5612rUmIMxoD2
nejYg3AIkBlwUPRoAqkmR5DqSG87IhObDq9YXajjLoFbOhUvN8w/sblGTxg4/pDH
Q7BGERrj5dd4K82oYuc4MpyGrUBP/XsRpGCe5PS4qgnR+4H3yMH4zEMGIR16GZ3/
Z9SNkLQ9DjhYOdKvERNcJV/C/DPOnjT0EX2ognZymYyhcgOs54kdTyNwCT5ml2nE
aWAdc65f5GeWy12rm4HGLvEKfGTWdH+s9W7RxbP5K6EBvuav0zg3/NgRkcyl7Kzg
U8H+XuvmEu9G1sq7fPGPy8dg8wMZHZkZ0f3eTjiGjlW8C3B3U5zCePFASToGnmTw
ZKTL/umPKC7jnlAyo4lSUcaob5embIsMLWUXfeVLYiL8oEGDVAqxI+5rOWf1dvoE
eNi13lQeHR3O0kG3pHhbd43129JjTS5Px0vXw6CiwZH21lZaAJpG7mUElQAyLVRA
oGgmyalleITEggG+U1hhhoGlV0OodHt6nQwr9ZCzeLCA5I3/w3XIrVUK5FfO0ZM2
eUK878Y932ryMizjdyNYQiI9O2oyn0lOFhbcO7pg2vhZLRV4PKYaQhgJyDhxGGL0
tk4XrktqJZkVIeNUS6HINFRkryEhibHcMj1afH7JTjgiXIRtI/CkzYqFKbZ5vBwu
81pYhNVxPjLVro8aHa6/9+HTtIt09d78sgFsE0qiuQvUlcnpmoZy9kMZMXAqgdVX
NUEjKmrR8xJhoed9Ipz/mBj2aODuP68gfWMlRMsGGsLnXJWRBSIBqoelMcBrjT6O
ZVItEtJHzusjYZXIiT64uBFnQU/n95AfdBd49mk3yinPhZsKBqaqEdL/NZhmWCUo
FAZbeOrI0vYoG9pV2O5o+Z94A6H4cmlcl8IacvbMfu110SR8g9SjGaFlD3aai+42
OcUgP7q+6kjuQBmIcqXh+pPRHYMouPFrIBwnSy0nVkXbP1ckjRJ9dToo12uTnVtY
oPGZ9+OIKRFm8HUzVAebS76h9LvcI9lqUxuwZWv6U1ozVVSkXYhkA3xLMEeqCp8W
V9SsV7HuRbuGS1cQ45TB5rRNYiMRtMysK4e4C3McxSfaqOu+cWsnS8SbKKi6sdUu
dwK+zH85MMPb4EQnf8nuDKPDCwKXuiP+C7QILXIjiKoSgR7XPBH1sBlXRz/APYh5
uVB5CFEAQZI2UnOrsRwrge8l9tHfGo/rBvjO1JenooLFgxjEh6S7Tqda8gmJ1wZo
4FsyRBFUEI6SwVQh5vwf9TDICIwmggq9R+PJIRw1IPOdlMra3bmXjkKbhsQH0xvy
82afNQtUivT+0MAicgSWWL+V3r0MLv3ahBxhZBtN7c5A7FxHg7mKWh2qDQnRcPSN
LkjY8I8xm0gTLEhqJs7JmiEs+e1yYRR6YrPaxHb4RnE+XP/42+JATYaPxtsd99w3
6Go4qBsdV6rZimU5PQ1NfzNleau2Uqt+m5nA6Ydqiy5ZNQ4GeqHmEMaab5hpkY1B
B799r9ZhZH9J/bC/rl0wu0AGMH+3ba0knqBBHblNFWSmko+/YrQTKlsMSB+QQ/xp
Qz4NjkxZHJTdgYlihGPXR/SKCDBKcHTKVvPtDEcV8cVSbxCXeNrDE3yoavG8iRQd
FXCvYE58EhrIMEoX/T7jFHxpxSOfrwHASanwMZrHoNCsf08qGVIi4w4pw1A4UhP2
5RGTlojoQJAoi4pPPqLIxwwEbGd6wKal127GWRuJwcg/ePgeIy7+tRSEdqd8LhZB
ulFnr7NH/D2wBQ95QYu9vCKtK1LwlYKDs8dMZk3g8KFR/vhHKtuxaJtCoK/D9vI1
5/RXZ6yb247HAGDwLtWvY+r1Fznzg1+i/J6ykOZ0m+IGofFMLbExhtagugho2Md6
MvF95U9Ro8+kStUGjIX8yvpSGRYnb/OVsEVS9POHvrXRRV7ly3uL3VO/8izgoSHz
ievarHhmhvKIOvINR5fQKUh0edlON/RI0K2u712DcWRJA94crlcd1LIfXZDdmAC2
HaLVLmiC5M4YpvJOVtfcMCaRR5c75XlPmYOmKVmKkbh9kyBB/0n/zSFabWStcwWh
6UObrJEnVfBJytXh6nvZAF/AviIT5pDLdMAmMbPMlna7jYH9zMcLIHS15QbxS/I2
hQ6B9qpeFalXdBuEQKk0Pd6jBJygeTn8oSJqQLVumER3ILIb2ugjmkvg2Gpvyzvd
c7reOKKQvXTZq56+Aa//Xpmp6Xw/2hcGksu3k7oNItQRGjooVex835MPX0q4RPuv
u3cigisre/TY7lECf1gf2XJ7XMRWRbfm2Wpb98YbnE8juG9cHJzMg4242qHeo1D/
HOuwl2MTCgpJPdKgLBvDt8Ml0dU2IlZIwU5stohhu6DfaWStq31M5DmEh8UU6/33
O1yiWbhMG+y1NhwRG9Fo/LV0XJZZ257uOPL8AtlJeLnIJab9Ace9xwuapqUvRG20
+0qIt3G6po3iPVBWZqD/GyaZ6vJ8JEWhL4S+EdShsfn2C3RTR4ri4qBijE0o0ZEs
A77xjPrW/kp4UMknv7a+qu4wnaZY6aNwysKsTF+J6SuanHRAfc7/RyhVN0rn5XQn
RVzj6FvbIbQ+K25lYNRaDS2JaDKeA4aX7i7fN0me9YFuuP1xe+TMUwNgRNBEUtIx
t/E+edvQNoXZR42WWrLPi5XX2Xbyl2O4drUCe+7wKPvwqNbH5+z2szafscZ+6xAL
Yd89PNDJ0ift8ZvWy91S5+wDYR1j5cHqX7M8i/ECp5Ro5o6MKOow6wcfXR7SC7T1
HmXDOY0MS/J61Lh80BswFfPrDYmrZZLNPzVuRMcl/E9Q9QIzyocxMc74ZDSuVPhX
4A8bcas7IdjZnsn5jW9zG7lu3XtW1h2eCjqG+NvsQ/OZY/eMarlCdgy4N/pS6QgH
+oyREvmi0U3UySe908LFxA42hJkpOypJjYLNZhP6PzDh8QF0wz9m0xPrZDQXGiW+
iaaQnYizqsliMYlhIuGEQIY5tq5ep5atd+m4KvkpX1h53XY4sr2c28cU5g5en6lc
BiFjY58UXXcrGq1j5WtKmtWAD7T7TiZmkFCdQd+CMKm5zaiI8WzfesqL6JeWVd2N
MRP0aB4vVV00enU752J3vMyvEi9CWo0EQNprb1os1GdyW4yWMQ5lX940x0QpoVto
8riQy39nurZWb6vwbdeSCd4iNs5zaSSFob5LMzbxLKXRIKn3P/ga3kK2T2wq1qL/
/d4QXjh3CgEeAoVYxX8IIMpukikLh/RmJcc08+r/mQExMFJuDopyId/L8jAFdcW5
9TVq58Pj4AYRDjdp/x8GhE57ZwwUMmPeXTkISy7t4sjpSVIP7dorOYONBLIufhA7
V/bmouyUNfJwDP3HMjCJ68biNOOllRwjE55K4z646gtTeA/pj0ywRDKnaZs9P/lF
QcMnyOLdCB5m62SX+QGxs69JKa5Dv4rlvYs+YAB04D94gkxSwat1dXSv6b4BA5cP
w/y2/c4AzuU0qdxkSx/zyVp/g5DP4FrNvYeRr/10RYgSnTSEK1Tti5CSYE86REoi
o5NRQrqeYNYM+w89l1wdCCI28mu8nUrpvLhRoy2/2u5s6qw6Ixu/irK4GSA2bVc4
apAxA388cysepyBKyEkXKBDd0HSwo1W1DKOPm0bXgAT7uQo9FCi+KwKJuiIV/dfp
7ZHT7qe+3flzhxXZvyCOeon3FrTZ4FLVZ6FoA5PsmxGDEUksoU+ScgQnNN0AwW1l
21Hu/uUQoxMxrME/t0/drN/29hUrlkPb3rPCeYxvLtU/KXtlGP9EOMeP5Uesv7FH
7EGe/4y6/TsItquAD0ooKRMQ+9qmxHiQ03uhIzZdnmpo1MHeso54r4EJhVYEQvKm
8a1iah6DRruZqJFjPMWnKqixZfUir4Cwgc8fcitnUrSAJx/4prme0DqNwtk99K3/
vrF0ZmmNhnigzHcpoQZGlaXHLTzucF8oO1XAQ0Ekhp6qM7mj5YoNgv7Ei0bRKzAm
w0gQbjyg9EI5saS1OSwc5bKDLWDr/92cWLFZQWsCbVIa1KpHxbG0EihshKnZmBny
+fs6zSsKFxm2bZbcxCzXHv4b88kpOHAIpWNXn11dL+3H0UowgFi16ZBgy9kOKMhw
evgaBXNtjZ/B6zulI8tj2c0tcs6ioYVilQl7gSWH1RxlGB3I5m/lDA49pSo8ys4w
OFQBypXnI1DYseWft17ma6RvWahy5q1s4pqt31iGSXIdjvszqDEsdBhD7S/iQS4G
cmc+g9SM6Qj3i4YPgPLlHUZ2cRlh8MwUJB0oHGG3jTJFCCTApsPHhWV7f1+GNun3
Sv8AkLCHMpHob28oPKtYioK+hx3tvBgBHwDQxs/TLTjNCbpl29i+uAWn6UwYpcD6
RqBTH3hQgHGBkP7lnaedUgp++BgazVImXTfeY+/sUppnr5to3lpsojwv+f+xBsfd
3OT1byk+7/JL78KA4FqCckG10dCfZcA0ac0Nx6td3YQAutbUuYXmEKL8pYj/ylPF
jx38D1qUimFqbetwBVRHzYthWvu4o3b8bd+jtbCC8veFdCRGix5M0soYXvwg2OZm
SfIuGiDFNgXm20JRu8SVXH/sURERcqX9LDv6nUtcq1ajDs0Yb+ANYDvJ/To4vK5F
faSO4jXTnNNaFdnhKyNjB8U31bS+6UhhqlYougiw9Extj8g0C4PHO1bKJWKSBREf
Je+ea5R9JBfgy26mHtySMEKZiveFCymj/gAuZHO9XeNFhcL2iv0KJpsxI0akWl6/
qhxLnjkan4YP/8vJ7ptzxmdvv+6C35JhwvvpgVi2OKdvjeeCAlovmQQH6NSQ6Wxh
s5t33QJmEGAPT88eQW3lcRXGzDOwlVXqejHv7R02Ut/owB0vZ83KZgHYrRd10tCR
b2N7HUtJhiwdfVZ1Q+Owu/Hw62hURHIdXWWJtOFH8oHiWWkydavCb+o+WlLyck19
nknsRz/AKVwvn74m4Gw2T62WA1BuouxgMwzD4C15QwdtXgtQFJAAe0sTvqYiOtrM
hy/v4ekbuU8T6dXdt/JQ/pMO+1tETQrk/QkJsvMWZ8wr57/at6dyAkWqMehVxif7
r3ll4L1+ScpJlH8e97EnDdlxT8HWwDlGqH0JlRyJTUpCsw97+xqTNr8hXQgOaw9F
H5wad2nP3i+L6z4WRwBqWnCiPWMSfFVRs/5Hzwuj8//oKbpw9QPjCiRuDJJTh6F8
dv1YW7PWv+31neDagUtUkvDMOsd4dxcFwykEwZdrbuhItuJIaKGX5xkQ7o2RGVPg
SkHEEN4THkp5Jl1zzmHKtu3LfTOrSLjgoXn9L4GuUjz+Sgy8ALumhZtyzw4AhhOC
piWtrezxyoBc7j3IYKzD/RuLAJAy3mLCxGAMQy/sHWXqyPloocTuTU3k4xEyBOaw
+Zs1pZh0+DAhZ3gC0OicNEtvj1JaAKHK8DfOdlI0pEk1b87lVWgY9x7zWS70En35
qPLlM/ih5/zxmqZX7+vUze8k3orWj/HSGWEyj2PQDwBENIoRXcO6W6Ldw4aXc8ia
DyDlyEFqHOmD2k0ZQeUPrmi3Vvyzf0/u5+K6lqdcJii3M04fqz9Hgn1SZY+LgSQq
WsXebQ6F0ZHeQoltwZlC3SpO9RTxitmSEFhIjLXOhyH59DTIsg2Gs4uB3xEyA3R9
JG+qFcGUC2ppEH502eNsyVwN2h4P3QRFfRfne3pwbGfXb46+QgbukSsOj5sVeJlm
NCmkrLhhbQlIzUwTIQfG9twbOEJ4LwTGZV+zoOxXprwB1mZByo6xpTcF/Kr7OJtW
lLGlfOZspmAoAUpPvH9vfthC4umas6qMxxZ9f683uJOTKD63r8ekV8DMSfLM1Weo
LFmnmRYcKGhkqyHVW+oD5icV2xYSykhrrullfVjLkGJmCrJl8cdoYvADnQRWy9Cy
hhLyjhnPYRiX4AFhnPM/mto3WIf5F7exd/ukhTuv2638G/DLlR1sicnO2n0cVFxP
BjumLLu6WUHPPndeDrafx8c7vEJl1a3cTH8O/sX0gpFpOWjXIkSDq5wM3Mm2usdz
BJ9hJpjRmDsGfXGDavFMrBS3y5/32ObQ5YiAM3JTvMs9AJnu8Yw95s9sFJ/RCIOH
A5MDHiuFzW/PTm/QBUYd7CGbyf/54/2VIkX6HxPi7EeekT8sIBd5kIfLVd0ygB3o
biaGI5ci8FaLx50fNi96+OeT0su9k8Y6D/YXWW4gljNX+2oTfBCMmKTLEftFkUyp
yEN18vSthMuk4f6lm217TKnhIpzEOQAm2F9d0D7qhLDfdS8uvsNkYdEtNLkrlrS3
rwodTNqorBr9EZrms8NwBKInT+++Em+2TXY5U+5I1Nlg9G5PBe4V2M19CertlhKO
JckUAw9L2HVMaqCgmXgJilR91qM9F1hX659slWRmBAj8kHWdEb94TxoQ1ZyckrMw
tg5hSsrNQrtuVC8PZimkymrNonBDPZiPw1jPgsNdlWTFHnBWAsPjQQnMMkBzvZLq
g1iWnvu7weW1eOSvg1XeJZJnd3PqrsC5hAaC2WUunuS5/4XrRTt8TYVyXEH/Hagb
4lHcBqsFtKNBP8ubWtrDR/lrfNLJxrZ5Jl4O5UOSvegpcXII+Vyc4yicd7ovXz94
eLqAsCIN3Kk8ODAPzqPUQ9ZaP6/h/mYAcvevhxlyi6AANPbhwbJqxi+pLcyQMHPv
gVEHQTgcMRiTuDDGNEOf0NBXfGPiVzHS9Rq6r4MF1e6PE3f1k+UIoa9Tcwnj6AnD
IzuymkeXKsgA2J4WlY+NuVvPPXF77tFmLxPqwu90omo/4vadXfLviUAVCZ0kbVUl
NiTlwTaSAdpFgoI/0tNh0Qw1HNG+7LvnXlVF+JtqUbnpjBBCVQ2FuLUeM9wQi0J8
zMElq8gI8HtStyb2XwP5oXLjVMuPGKp/wN0ebjGcM0Euwt8YHTJKJMchxtTriBbq
JEw+V6J6b2dyXKRuiBCYvFT93Tj29Qcms0+GR8QNP/yWOvcY/mxh+wK+AXJxMtpi
SpKJz1te+dZ6RjyVBKkQdTc7BBrhm6iOUqy7fhI8E/DJ+SbrFZkz4M8pqqwzU2pP
frJ4sMaR8HWzi7K81Pb3UDfikH1FER4EL7V4sfHhOKIj7xqB0BvahMHZyqNVlw/n
JlXX8OxT7K2o99ULzDFRRcoouI6F9C7TZ7lqGpUKt+I8kBxr9QUYXU5G1WczR4/k
pWOz4e7bF9sDsaWqVT6wXYv5b2ivD1wFDePD4rLe8sJgjwiEVHnUiOjO94k5lzlX
v92KOpnTgnnRpvbTw2yMoQYVCgqHMuSo56I6OYcvAi9k2A5orlWKN84ovQM9GKR1
YnE7vvyjD0kH6Whv9yXVhQHGFk9JFml4FNHqbYktewgtBqgQPvrfNesp77OabPnN
PAlvvrpMaTIK/GxPl/Lcj4Xghf+M7WSYO16nw9Gi4laUqesZndzfta8YlkIMf0QM
/h41UqUek+Bn5Ea9SfIgEFfqTOVpzHuIJRkLf2ElQyVyRGGFTjUhJ9epC3Fp/Zo3
nwmuCOxcfVZ/F4EDhR8JGyL6SHH3RWYIHykVcPeV4Kw8MC06YI5G3rsUItRZ1syR
z0odmFP6jzF/HHnp54urSKWY7AYoK6bMMMVcSAJDhw+xmU2/e78SaJtYGH6RrJCF
r/gxIJpT1wUSSglqJHxEYHPgN46dng1kge5hxyvaQV6LuKDFa5AfjJitrNpHCTQO
nvuSVY6RL5+lasXVARx8mga1ILZT8E9Wb7SFbaWcJfQRGnwZqoOhV9+VuAdELn4V
jvdFPRtv5uoQ+IPr91vkdeJ5SKVZLfA9s03xrywuiFjl/nbtyDjqFhKXBB+pFzDz
CARETaWcARdQRyXQ/feyBWdBnVCGEAl36yryjQd7CdRXCX+ZlVIchZkvKnhNicxP
1CoseM3Yt3qc90gQ706ez4/pSu+vdPDemP7146BeMsDM5vS+f4DcBJOn5D4rFRQi
bkpk7EcLo3vYfAW5ImijG8aQ0z/Llh2UILn5blOqzD3EfiChkOSj4LDVH8MbX7ip
3rOC51Zhfg6QTH45YGicHmc9TyN6ithTTlE3G5t3RNYimQsFKELwoKOqWQA4hC3Q
5BaGEuk2KKqXk+QITA8uf+KKcyUxUG2QM0K3OZcD71OGqZXHiJPtFiZtASwE8J3Z
U7F/grm9sAE5YPMOl5e0PmabctrngbyUtgBJf5mqDqcVGBoggO8tnCJRSnbhtV4g
PQ/BJBDXLfGnowchOubiMFFOFzQMXwYTik7oaYyux3qYsPUDZSLfpbfwIg6/sNUJ
qd4YaOsLVlLyJfdZY+nrlW1Tc4/RWET7CiVFNoYPA2I4qunsoldAZ3qJYIM92r5N
vFCAbsIJVwTqB+whhbWg6c35QczAC91VVeO02erFmYXLB153EFzAssWg8fL3WTrZ
8oMyYon+NeDHiSp7OyGXH+3KBhJIrr9hWR2d0jW9v4Qn90ltM1w3nJhdNSgS2xoO
RwbkE2w5Wf5UT88V3+mj8Llrt6PuJrNQbmyYX6Z02YYDDOtR11uy54xkz3/TXCT7
8GZSGr2uT2GYExh32cEgayQG98a7JPbd89bZfEWxGm1tCOM/kQ5oIsjaS6+lfe6A
cteecES4wNZ+0aInLDGVE7QLrMBigxnmzS7BpDyiGdPrJOx11eXXtjF5Po1fkhj7
bK1hItZ0SAYDUPBcXBZqTgEG7hOW8wARr6Tya+w8r6iBGlltW7L2F9/nzgSS3mzX
yo3cIlCTT8Ni0CzBOdG8xP5OM3cxZ7zCaGhs5oHEZSUVUL0t/aO1z0PQ7mDkX/dE
q2EUY048x1TZJul8l8U2tGThprIGSTBKHm1zompLMPmBkplg5sivN7L2WIuTTIaq
dWfFywfux5Wc+0oRr/OW5hVOmdOD4xbvWtR3hstvUcRkiV1iKlm3/2nz7WSvkW92
6R7ASS2iv8DNqR01KZd5/SvOYMtQaSFpca++GQGn0Uf9ZQRE5jLW18xu7WGtR6mb
Y2gSo6vC+NpStRG/iVVHtmgJPRxwSLw7lsDmCiZvraQXl52azbD18+qsLiuqfxZK
lxpuIdtyJfbfq32CvW0ymqc3jWohAHtimf35Nf2+L3PBuf69VLnDwyXrL/gxPp60
+8aYraOQkac40nU5UarkpnCOkqsmRHpneE8/V8ysTUdwuesV5yh9LV4ZNgB+qSrR
lVvwgPXOYV3Sgk5GEgK7I4lN7fbaN3ggUa3mHu5bhZda5QA7ajULwk2yUxLgK2ve
afwnbejcJ4pUDanuPMS0kqQjC7UF2U+gdIflfkyO+7ZXP/BahUGojdcYcFxbs67D
CMYuzigTFnsdk8AvrZQT+sQvcXQ6jKd9A7GqukhTbWo8zJ0/9M/s5aTXajuhRtLs
XALw7efsFw6GqU4rl1Z5X6d4hIBDYtZ7ThK5ZvgBg+NeqVzldy0cSP9v4lAnMhCb
JQdxheXEu6pXtvpp+l+WJaxQ6e/q8IbfSeCYfSSAxDfDOX6QxbEtehFAF7cuPQXe
TAigcsQ7EzmWJG1vudwSKWUtfHZ/pXNavfH+wzfhapclT/YGjYCIfjCQvrOZ3c0P
9z0hImm7EceQwXGXsezL3raohX0qmXz0RSRbXe0FHMFPEz0f9LpXyPmbZ7qUkmJP
xyrt1zF/MnHnmaf3pFr9xFnY6bqox5iTlzesLOgb+oWbXCgWucSVi07pNrMQuYme
Sq7GMruCiGTd97Y8aqNvDMQ6KV+hdUkPPfJn6u6yn//3YFFnA3fxXUmYeIQKqMNB
OxXPpqoeObTaNFD0tlCbSXqz+p1yu2pcnYeMrIzH7E5yQaZaSUVR8KxPGPePlb5a
sLgAopb7NWUrBLp8snfvPOx3sNJbCUZ6o7BI6I9iVlbFIUcmpEZK7WUBsCC/hJg6
4D03aLRhCKsyy/SsxI+rkMQH5s04vwcXg53KbpmJM1HapHXnEXoZ5PwJRCB6Rj3B
HWTM5CiLC99otAms6WB5TOrZwJGWMkN8BMq7nCFtxLY3etM8jkmjzBvZ0Z4h/CXr
H0SJq9wRfgK/H7BYonHhDjMZo+SO0XP+NfsJzVaTYARf4njXSmmW2iZeyQrYs853
56VdHdkk4W7FpTM+bgVJ3qxZz2zXOMW8uQeqihe/8NQGLtJxrIOgIGzjNAIHaJ5A
ebFvEHor6SAtjUlzUq8kk4o9Rcu159Z+MOKpXkiqM73CLFaSgRjVPDJ9O1IHC2kX
DsgjB1P3K7zdjZ14j/3STp/rdAkKS/tpfTWJ+YUNzh7eBTi9uKhaz0mmkPL49DIR
RVMQD6kpJhdqyd3qDZ+anTAn7j4FOdZ9zBgeqzwzfJBAJDlegd5dommYy/UAjiWA
jVaWqSrZ+3e7P7z25d8yhUcZt/wJ86lArmwxKzkS/MN5qRpXPOpyxZOQ9JdMgp4I
8vFRfxB2rUs2fTIRLLlSQyGM5mUNsBI13xcpDN0Dt+EDZD2F79Pq8wTp6NpLO5El
pOAq427auy9sT4lOHQCdeln7S70zfn25cES5YZ429asMOgbWo5qny82UKFCcamHg
7ZqZcjzv4EXzzOJlczM6CijbsSyO6xSmNXoZ5rVS81uUFPZKDuMhjhGFA0NL4Vtb
6ft2OjLIPajcA+p8O+hKQ8HHxfwD9mmco0lh6VxyHL81Sy+uKvLounPRxv2Kk+8Z
t/sxDFfopQbaRmL5aGYyoJStFpq8AYIGZ9Bu6ENTRCbpnGQr5h4vaf+JnV6l1ROJ
zG725e1EggZoYmDQCjTxYXiCkmBdnMKT5BkI6qak+VvxKIPqmSIl0Z/63DKmEdyN
HXWsrwyhMBIPdN87ZKvXlCvcrgwDFGfqMFM6uJsB4w/4YvnxHHeCEzgUEAxQLdNY
KFWQ3wL8AMgCtxUekyRNVPXKM1Qr5mqvupR3PUu2J32w2we+SMizDY4k+UG7wUx9
eRxNV/R7uhrqLB0DdT8nzSzpC6DLISRctNznKbYTZE6GPGGWY8K4iGhGrTyIc2If
woeVGL6tjv08DzP5q3RGf/LXy5AtD7fKzZGWX9LNEzhTD4y/hEmTU+cK5y0BM9fu
geIPcXzMLLAI0EcuKbTdx+ShF05k/GP1NGT56UnGAZyRXX09QEzlceqnOR1S1jPd
4gvkhEKVKx8IT/+hnkHK23u4WWl5U2sxUQBuO0DG7XiluFxp9cIIU8sU8WG0pTbU
Uo4qTcN4KbiouCw07y4YyZpxyvfv2dLETyXgbT0EPKFFsvWzRW6asDiCAikdrF9w
5lRz5BpyjaBvDXD4xzytknp7RQu5EXYu65Bu+k2Neh+6CJkATTPTHHhq0wFLNtq6
7OvfW9Yoc+nVCyXeRxzELpUEvZS+qEx1yMngCN2B1y523LFOYPIoXzPcymZA2GiN
JFEvIZSLIy4W77hRrQnulU8Xgj35Jh8QOttUHeG6IqdFGcx85QuAk5c7NTJBVIkt
gXqQpOVOYH1g+XND2tMQJ47KZ9bQCeENtd0Jt5S4N2Byyoig88KOyrGBD6qf01zs
075eY+Hox+IWRhdt3tpP8D4R8R9gcTQH3Nyxvh0vjch4oJEWMx9NvFiEPQZUztPn
Sb1OUauv90URSzz3nS8zSyb3MuLECj3O7JnPVAktofn+PJymkZPRZK2xhOVev4WF
oMOA0rUxlV2pzHnRJ44vtdFADjxaTPrFJe0tfwIHi893SyzxWm/n8cjV4ks3eJup
zhP5fRLmG1CfOmzgJ0E2qrRnUBcIdXM/MG6v0Jpf+7Hddxg8W4OXpBmhKd3MArA5
Qnk6dGjMU5pu0tGENwCzZa3PEVx+os8eshqRBQrUnI2MZC4qhGT8dtPoyegUS/XK
R0o6bC2gjG1jMV4+8hF2fKn0sUfoNP2TSGum02vhJiydXo8pZkvzXs8jkAFBrqO/
W/HAK20Mlsc8IUnzEf8pipWjrZePv1lycRkLdbvkRu61f53TkRepmNnzhh51r4U8
kZHdjfMObeTyZ18S/JItpVS0dRQxBdmaOI/Rpv6huVBlbw8P/QhDAkG5O6ULHu1G
axC1p9L5GlSomlDI+f1mQ0NxEmvPh62gadvFxFZLa9iNuL3fmIvpp+6LMY2aW08j
05AJoX6NqKoTp4zzkJAYHuLHEH8fyKPk7YPBVi3M4T7aU8bH1BDYoC40i5HRNa7s
Flge7RyP019cSlygIHApFAatfGAG9+p/q5Oxi4+0EwyfWbr7sQo9ATGoKds5eD+t
Yjjo9JTihsjWZTJViAxvkRiTY+9E/uHjtVudE8aMU53lOJUUH1BDSxp4fffcKH83
J1MWmFN2DeJLRD/aLTkIZVfbGOTCGoPFNVNsQ1Q82kKMmdULmb4OT+BRR3M8g9+F
t7AEy4CZUwIj1dm0Yudi3p8LaPiIlFdTi/43qEcQj8aPWW0WLOMDlZuzySp7j0pS
xaHSZ2u2nCZzucRHv1vpqZG11ch7Nphdmw3WgC4vqW0SA92qHMum0o3C1c8isBss
pQqMIuz1kvN3DEEtAeDOaompoojPvNJ3lE6PRce2uJhR2IGW4WLcjKhJucxbxXS/
4ITOlLWMXUWLe9Sra+76HHchAu1ypHT7RBjC/qCTAHkUy1WOC3VE2g/miyS55zuA
0HryhnUYpMZ0JJOPothLm822Wl2T0EPuFg88Qhv58ieMRMzJSBXiEsCBbKDm51Vp
FsBNsn20IrZ4MGydWpP0qI19uRmKnAfl/gNxa4t1BM48mUXgh80aBCn4GKJtl0AZ
RcynYiG5D+lmTudF9lMnYOjXI4WWgvgs5ndL/CRpvm8Ly/wbKa+tm3TG18g/Srv7
3vu/csrEeglQPdqPZXMppMzQiGMCV7NZ0C1ZrkDA2m0//AjSMXA7yONxgCtOXlsa
9L6eVGKP0cf1dYCs9HUQqnwB+DncTFl3Fz+mHMVfuUPEj13vu6ppcsm/Pp4cWAJX
kQBK5r67XY7ngQNbJ/CZ+FPqwprvRjT/1vSLv87KvRa5wwy80MDI3akYrQvO/aJf
E6crB2u6h3980FHhq91TuW5/dm8lMVxnT0GoObDcFELwfNTviK30FdGd7r2bMqy2
o47LfSMpYYJDbRxG/9Mfdi0MMhtLAT7lyBOUpmVyiX0bPcM1SRb7BNigEGhrXBBn
6/OaUAbpwln6aWGtTRL9cr7cLKl9xX4lKcoris03DQQXhep5cdEXjnbU/zMhUM+m
OUxhIg/RLYODKv0YJhwH+nAic9NzC4x6nk2dCQdrU08Fio9Yi+KOWHvNDDtsz83G
LD5yHyYjfDNXaWHm+Qlgx8MKQioOQzULZfFQyhjAgyGNwXVTeGhNnhIXxgUyW6P+
dP+STuUBU7lctUGSaWQpKvLyBxOr2HkeEBc7CO/sP7VuJzKA+mzFeCLOgqbNs/fm
TAS61BoSoE6lbSbb3tbl2EJUv+G1pjqPVG2DMd4Z5PK8XcP40nxUOtEr9AKyFon2
ttaILwVTAri7FqLoHKvW1O9+NdraGFU1gjAkdlDrVqZszpRPOYwyFJ0Gn1Z6M82c
wOdKu7Iq6iaTNXU8dgtvtooSw28G1FOEGphnmtXJ2+0UOLrJD5Ioiw/i6J8K9m4u
c+Rd88KIZVpN4BxTKJP/Ph3OlaZNBJWFxUrYZkVAirL7no0kaVa4K3zbfJ1xiSmV
aq4stHaRuzPKdDn/bW7/LTXlbk844rJeVwQ3ksf7BvADBAGCmMle8fxZ4nwlSjAp
TwujoWZG5I8B1jnuYy8Fql4TY4wXFPtl6upzZT9PHB5sCibzrviq5vt2JQo4aC3j
5eMN3sGTYjFmrHr7kINCy11jyzqtu9GeG8lNPrDrvaKzQ9/0U1SNnYsGdlIOfYSQ
A1chVdjNpCn9GtDf3LbEIwglaIwonOqQdfNif06UEA8HkI0+54Us6X4p5YHfLhJ/
Ltaj7Q4NOYsiW6uPd36X+wm/jXZr5rknDWTAguYRRxjwkkEtOjYDF18F6tLtOQYd
Mvfevsn8FuMeorn4s72hFCacSb8xRIQs+Esh4NbBU26H2iJTny/Bev7JwVH8IU2p
KA7XwI4mXJV2rRgP7yCGwRvceSScBGSxeKexcu3T/wOVVsyNR+CRUz2qnkIuYaxf
ZPvHSR1wCCL0M1WTKm2TcYo4mzofHceDDm3hHaxeT602naJSDejR7OqD+RMoPkxD
BZF4JrGjasyyXvR6WY3Xd/1ewHXuKNZvh47yHyDwLkQJILCsRm5r5dAqUulDXt8E
NO0uFJooR9H3OBkcsc8OIjG8AXDf9GxOckEef6iDbK63SOtLfY/uTcncb6lm2pIb
0pDGXhCsT8LCvF2D/W0Kay/inKJXFbvI0LvlKYRbVsBor5MgEGFp44I3NJk9f3eI
OOGbVIn1EyEehRdcdcSqqzjuv75/6XEKEnfl/mAgLmvHms+RfDz282SVZ9cV1uff
5zvXChmY8G8Yz6DsBXcc4OT2Zd8X1UoZVYOcb0f51/KHVtInG5sdpp+PJKD0qsOt
lgQVltupZAT8e2rLF2U5wP8I7cZM7Q8XSJYSZMam+N8UWO+dv6MAKCSVfO1sUorP
+uCvYAxsNGJGVGj2ZrWfaALRed9DPt0EkPdV7ZmXeGAsdTlWtr28TJiJgbUwtqXK
XEjYHoLRmAviUcB2EmzqDo3/UMUxc/6ZxBxdunMOH+u+lxJgG6xeOwjvEKfUzSeX
NGKwvbiddE3PHlj30mI8nkKdwOaBQ+hu0Jf8kNmnReRblgQVgAsqa7AdCMYJ1kBN
DI7tH8hBXdIGUkkF2+w5eGor/5WcQilOIW9kzqGiFg2aVFqNipfHCxd44b4JRBU0
9IFbqelELJKysvG47MPDtxRdpJrDVGKrOxBLe6QBawHzzhq9Wt0dp5FSV3dgLIfY
k2ZQbyMWDwoLWXdHizNOsWUnHlNyqozQPRb7b7v634SN7OrlPpQPPw82jAZXybmk
A5Izu3rCz/UuoFi0VIJ+Hc5azHMZ6R5JqFcAXjSYMStPFkZOj+7X8nRo8QjfpX1d
Sc3bR1hZdleeaqdbdfRLHHI/7H806kG7WVHKNmmnRrSh7C6MfV4Z+uqdLLPRYXXS
aiQ8yPPuz4Ge/+6/hlB1BVg5s1XCcsVyiWJrI6QVQfjCu7f6RDnthlNgg6W2eeIw
0KsqR59rk2oMwsf8QFT9ut/bt6JEoliCl3B7R2YUGM9Gy34cf57cMTj6eJObx2Xg
9ny0UiysnNGhXiBmll3evvFUBU9QnK9j4DAaM0Cm2jueo4nggPEdxfbVNjGm8N9z
+re9MbnBIpYkaTg+tnXwUjwXE7YRL/uxmbLV7Vn6qVpGOjYcIGyq33OJQwegDUEW
Ce1s53+ceBlnkkTAYE/B0bRVArahrhkbUCgFFNlrOtbyw2Eh6Au2Ks2QhlN0w07Y
diqIip+B9NNCehhzskTkM0Q/RR1NL7ty89/EM8WbcImv6xW1Ds2Y+wYa8aCHm9bz
m9zvb3zM6YTONTk7b35Wgq5s0bGQ1mUz3RIkrymujECkCi63xHI1O/YPGPTzhNOZ
MBdKUdu45BKF2ABNxMwnLGIokJLUHU8AhX42PQluwdPtJzRleom375Lh5P+ZgWqN
bOsrQq8MgkS1q4O8vavQ4YehPDyazDNE34SXGLNkeelSYQvEBkZ3yAsF/TmEQEVK
3r+hNFSB3XcsVm0FFU+fYBBvLspVN5uvN7ilaMfusRcndUtnNeV7mx5Zp5wJuYkb
a/p6f7cJP+/vT8XdBb2wnsGiOn1XuZtgpGAHdCXBSdzStrqaE/nIlOPa71jQcQqn
FGWkOxnGrjh6hTiZdfshZZNJFaHHxY6z5Jtj5Q5EFJRqVeGkXl2er1Bz7NZJsGXR
aqIbg/K44MZz/ZHzdBA5X/CufA+cYxAy+Aal8NmI8/gdRObe8Mw6SjQ0TFie38kA
cCei+xl0VmoYLvZ0SKaUO/txDDWFwqMIuwWAQaj7LT2d9KEL6hBcN02Ir4QyUgzR
CR86S/I8E3dCJXzxe4B02D0yHJ3Re1vBhNi1iwl4Z30qwH8OJhkxEdWyrMYkOJ+D
1zAvXl6+A1kZAbgCaDWclc2Tzhn6PyH06Q9UJomNbVYigVO946O/sKLDfR0JREvs
83mfQ3I9FK2Q5KnpowrnVnFRHmLg43lJTrNm2SlJ2d4iVKokgfryWdcPsQ7tH4+8
1iCkL6sIEw2oRBsk0gsRQ9rfYcTjIgJOoyfm0cWbdDUhHlXKjzjRLWoRCFcQnX0b
O8wwPmkJ7LZsSzXlkDt+2FFydxWfQzRFSzs9oCqWZqd+mjb2HzY7Z9q9se9gGji4
c1+KxuPwdVY9eNA0T1sBz/OufBY58yRp1A6BAkqXBQtAj+h4QICt7z3szLjaX/kT
L5ITQUG8Ap6tjVb9leFK9Ve4yiIkPYywAbgR9IfhE1zpcDpLLkKc7d4uW8NVSXfF
aPRQNPj5+1SRX8TXUZR7m2lmHYn1MAcE+XoaOYGI/4CIurI0iAQ9PxYWLPCqIOAF
t88EYzVMQCDJdZG+dCRPy8+8OIydfDzv/qqnhuaQKaOD3lw85+IanMavE/Q4yWdK
zEMBnHf0EtcxrOf7z51XpyO8ureUqCSp2gW6K6FEgr8tPvgCM5pjWsfOOjZXVfNg
LbKwbhH1K4XaZJ+k2zZSEuPalbhkI8Bo7HwxUq7P1X3lInHJyeU0jkUg1sgNMkFp
OXqZlwv8hkVjg04ecG4KCZMeLVAqozEUZeyEXsdltcLGs8rU2GERyNiBhipujBY/
mFbynjGJWiQbT0J1hFUno6g31XdIg9i6ObKgS+TyvTh0CI1WvAF2ZNHwpFaiCrRN
QRw61p42yQc27oawbtMMupcjlk3Vl+7RwwHAGFXrA9KX8MIpINY1/VtatJp6WWPx
j44w7tYhoxEiOKWnWTdZpBrQh/6OWhTqimUcsrkr/1OFAEak3TvlHpGmLKCGEotN
q7YIqFUVhUqBh5CLcrdSvb+aX+Bqe736GxoavuTnjkS8s1e+rtHlbrLjH4WcZY+i
VQt4XNbnIMrGJFpdQW+Pttan1TG+bmizfkQKxWYQ1QuN7u9oqyahmFE6d5YNcHpu
rMATknAsZ89h1jVfuCYAG6h4XAYvTqB97HyAZ+0DFKoqO9O7t8gL4KimeTbwuRog
0497fHT4DtLDgBLnBpABGGf1MlhsBa4Jsu7HMR8I1GtOGVg08E+7EyUGymXURx36
aUPR2+LihgHfbM3pPtOFd69oYbGX5Zh+YnfEJ0EQbgmRW8skfurRUIbqfS3igYlA
2dv6xxed4ddza6nznEb0TQ6VkY4uBqEE/dx34MCZ+MYZe+MWuA6s1gChX3ePVcgu
L74UadyUG8l21G6jTOKv+Sur37vmFPc/SECL8T4NPxaN99lbIWd+5o6NaOFlLtDf
aOZ022PTiFcGIZQwFjdNQD6sIne8gJ5BQ6qYd8tiJnu/+2+NqY8WngiUmFczoi8j
dz0Fs+M0iky3fw9/ta7fsiutTrRvm2w4HlmPbNqPr2JS64AwlvpPdO3ckNkJmsMW
/Vqry81I2ARiLiA+gW/Vj5jbp7fYbds0QmC6QLWhJmf3CXJnNfna07JRDF8vpgx5
VLZUR3rQKCVd568ZuhoSjJLd2zoAeO/Z600kay/tqiEYV5Cs1vf+qKt8EuiCQtww
XLQV+aqLC/nQWzxfRVXHHKTvhelij8jo9FdI5cBHv2cBM0TSrZb7DwQaGe3ysNDl
UwEhDPLMqrWmEyrcDFaePYc6zCmk0wt8Ubdkvgt4CScJuawGWKRrewy+ZMA/J1AN
LTdasR2G1aJEIs0mf/mKTNuL8KfxaGVvoyWl79jq8wSkKXgl2ZPPeseyK4XIT1kf
+FQ+y3y9FQrTNKJcqo4k9AZxaNVV6h8I+jb2S8WlXGyqLZbBIAUG8tX8pIx5ACnL
hbFAf0toADYMXdbLPWok4b0TejeW0MC26JYuBj/DcL2fd/KNnXy5kCx89Scd/r1o
E/QuFxJ7Tmsr+Zzxs2LRzjwHoJlEr2gKbTpJ+Vh0CXDF6EeegmuG+5sRCrL0tlkD
2pnOCA5jXCscwGukZtPLUAizEU1Cj+fTEyMTcg62ElFbCNxZTV7nSXjLV5/hkwgF
cG0Ca+00zgLkN0YheU2KPLL1HbAcG/i6ktCSWnb797uNPwWKva8NJPG1Sm5PalBx
LBvFUSEuVJJC2dCTMMlWLbvYUn3Pnc+IA3GjoEsyljNhTWDIT1rJTcXdF+v7J1f1
ujqkcvvcAbOYj1b/JnzrMNo7n/innzeh2SjQQIQB+v+LFhzwLYjBT9RXY40RYawX
Pn9GEtg9BEHQDXxX0SRs5uXEqzG0kZVP76GWvzJ8km2wsggiA2rJBdOho3nElJeI
Vq/02Y7ryQNAhFQHF0sVRNVdcuAdIs8WW9W12CwIYpx/Njm6fB5CrR8K1WkBBYL1
u1c436YNxg9cAscXLG+BmOaun90ZtCEqvKWriClblhQd7N+ppYOW8U0pnZc3TEqu
h80FWIa5DUwcsl+zOVOZpHEbmfJk8D6aAXPMrWo4slFfbBJQ/qC8rvFk4PX3hQgq
iX66m+aRQHtpxnaFvop88s2UF8GG8rlaQDXPDMfn+k4UX6iSkGbuYpy5JX0RZK11
pkR/FwzOJD7D6YTK07dXgCMoHa1/n5MFN+1MRPyoLwBN1K8KNqugnj2as1j9SHLF
sd/KgaVG6UiEr7e9Mmbnrtk8ETKTzH+mnumz3bud7M0bnC/+7d/Lhotlh6I/ZXW9
zGs295wJw5kFGkUVgwCp72a2vcjTt5Vw/ault1wVu3sAnclQEGOXbmMcRvydYUH/
qTQG5FIGdiPZcnHEX8lnHWmGdD9mkBM93Tq1RGFoXkRipKdBZPTDIq9d/KK3ZaZW
du35TdF1JXX94QMMzqgLAZLO8R9utJr918sXN+Xd1rzDUk9rgr6EPGdluQrh5DCT
0ec6ASt4O9dhw/d79Z68X9EQImjM78cBNHVQaMHuygGzTc/yIIpVE/D1JEw5DkxP
7VlJlAR6DC1S5iuGoOhXHzKAfxDSIx/0KRbZYAJObfKSlqOZDrBfmq4sQifqrgGd
GYiaEWvlLsuigABXVtBZOZvcLmSA6lI4JRhqTPn5P+b4Pynqe1+pJ8mUYri5JrJJ
//Y/mHZ4+IbF+G1AhcIRsicF8WmBgF4AzBHj3mva3e2/Zq2n7L7gi4Nn3Sa94Gmb
q0ni6ezW1RSrRQ2lpYawvBrGeVv2r/SSvJMPlnKE7HWn/ICoNcweVkqkg/xYfH8M
bCz3nwzuWxlBMB9WJ0rokJ9rf/+hP91MQKIpFrbcW8jxo6mYYYrFfGYG/pWLUuBm
MC/CDJ32q9Z2WGe0gNvLWmpSASCkIJrkR1oaO5ghZ8qXVceCkv/vOSvLkxww2nx0
Dg7O+SWstayVUl4M9ouiAp37HJ7qd9IIL41mt/pQfE40yDnVjDEpUM+ccqkRdbMw
ITwmXLuI3EBQySTYOKmkdea58ijZVmgYD78GzQbi1PWsTcogXkZJWtLD6BeBkGbn
BEMY8zmKw2XnUV9O1Ya4vScobRFZhrXczN2+DBP4Pj3ehesMQ+coqGdGWn8pEMc4
S3woPmBMrQz4P8P2CTp2jndeMqGres9Z0Lo0uUHkKist9iD/LwgvWZpgBB9yWKYj
aua8ezdLAUK+ffNMGnzcgkq+SoY/917g96ic/W6Rj7kuK+kqsKT6ejmX7w2XX30T
cIyXk5+pSjLbBY+jc8XRxaceYIFHCuvZUMyj5+ve2QZi83w2rQRZTSutYcAZ7ItB
fVsgz2Foz+OQhaHxlGBbZ/UVVs7HBmrWPFTKhC/B5BBS7N+vN8z4XQF7aMyrPSAe
y1m0oODxE6p9xuJcgdr7DDUNQtVPfRzX0Mg7z/wxYSuxQOsG10ftMYy/LGx8bl2l
2BYHMD2qaORVomIM/ZTT2zYLnsEw4BKluoJyWF8ndIulE9f3pncTsGrgUCx9kG5o
eGpy9Ug3O8PwjAaCvZwYczqKX/A6vRuukgSVcVPk59wAVdeXalsQfndydJOBMGMM
iTWT4Tuvhc/Y4Xk3UtRjj+JRqlYDdT0Znfdo4TWzzmcONz2GCJKrgkImrRmUwUe1
xyLxYv3PCPen+W8O57imQa6mMD6s5ju8Dy7Fc1/zkp/E+fc1OzDbq4+vWC2RArE5
sTz8NzHtBD6rB9Cs6fmbFF7pKHnnd0lB9vwgE/082HZ4HSujFlI9a8lJZTjGaoaH
yo535Jlv0j9ZsvtBCXZ73Lmwx5Dt14Mg6/pLaRDTAIs/Pxx2PWI7Nc3j+FTePa93
IGFkteFe+Za6xibg1OpBWfDM6v3LWaokU3RrEtEVzgdiSqNHUO0bX0gaIe4hZX0x
vzy9Lg5wuIWQQgJcm8fFmYHj99I5mDEDuWC6arHIWovjqVWBKNjmu7hbOlnizh5Q
a7JlMWrx/Tp7R84VK/76Jy70d0OXfvr2rfxv5LreXGmrqtO4Pu04XyCdaU7/oBm6
w+mVAJVeolA+Y3xYvNvJXi4NwVlEWjN73qTz5HhX6/I+Z/WQzbZMU2JyR6djNayC
l2CLALkLoJ0fdmrt50YrX6/a1Mm4vWuz65zHsd5kFMQSAamwJluriCyOTt1hQU5G
WkSm5c9gbuB57feA5X4vJeLvo3Iiyg6jN96TxmzNhxq2dkfA7dCVpd59ZuhJWSOB
v0Wl+Zp9+SYwGi+djZIRCnYivJ/b/hOh0t5NtsH+Z7FvEy4/quXI+7mveDFLulXz
E/PBKDh+/e5Ycu5Md9UVv9mhYQeDf8VtUtwE2/40YsB9H35I47lgHG4+Pu6yO6bm
3D4dmHdQyHwEkt/kCykLTzfiTazUizEL6d3PvzJHVA5Q3xeYIDIe/YrcyXjGKYYr
wrx9yjS3AgNqEswtbU0wHv9vQuACZRxUwKYGbc0g5971srcA7RexbP2yWgHW18MW
ARlYZmLosoo4EtGp5TRFMm7YQ6kEdI97Rig7jgNm4CiqGOvE9ujdQvScWSRN88ge
scaN8wOdjOP+L9snB8A/rtG33W51zzVfy7eFHGLXhd5XxgBWAuWpxT0kjOjJswP9
t8mLtA8KWpvLFwgbQXy+dG4mhXjXjFOgdjYUZH+d85tbz8WqdbS6B2EUpVlUM2N8
n7LNXDlOIJowqEPeMgN+/wkrl3IEORPET2xJ/TO2o6H56C/3ITPCIOU0AEjWy76j
5S+Ro4zs3il+zd4WsZxHYc8h1BtLfjThcvIzlHeVxtmzAJoIA2b5BiHKfX3DGgxQ
peRzFuf/9nFdDGPSzN/3A8nuf3KgGJDVZHkbQB6nv93KJWZhH85yv8yUYZzh/mAQ
emrf06+W0WZcTHXYLvD4nJWyul/V1ejObejvtPqexLL3TzUbTsDKOpdTMxLjrB+o
ZQRLU1bzTrE/lKjXRCam/Qozq7B6S8tVXfueamF5BA2/LR/KGlLhAuOObQOaUnss
LVHkV49lLuBaZqQf9sQYiXi9KdJ2veYXikj9+ti5K0xjKmocMeN7qlCmo43pchuh
XWi8DVx6BxmmlQ3QUlKtQ46bm7gCCH6biqmM4fj15U02qcmbMg4iR3IR7cVbBhVt
a3H/HupFx6S6+dFl/hiUh2+jMVsBVGEAyptiD5iKorkN2u4zyIdcTjdTfR3n4U5t
LzRyCuKFKfUjvFikdTsSUuMU6gp2qAwv4mFCXI3ccJBmutr8MWd9ZL0l+SUOcidF
CtxQMrYBpD3weLUWt/9rDSiRoxML9pJ31p2ZBJ4URMN2O06X7X3Te4be4NhfbEoP
M91mB2aT1sbvFEqMltzlFlmmqngbDx9B0rGVuG8hznk18masK5E+aieHtkMblHXu
PQc3AKpSiiZe8MZe0WY5wOj/iBcfxWNlMxKAp5+ecjYKOb4UsGQnj4s1rMIiDRwL
aK/VoTR2k6IqzmqzNeiCY9m6+iaEnH8OJejpivRdLiH3QTUYi8wgjMeyBwBS7m2D
Air6FpJ9U8ziHuaZnDxvuOV8yLI4JjsdV6REhJ9PaZJwqt7sp1N98bhYxLBs2dEl
gg3pivQ3DF2b9etXlX2v44TcmEREGGhsatkh9Hz8d+irkE+GS7XcLj6kP9JFafrJ
qvTO1e/sfymStRfZ7L8JiTvugs0dKjaXvWxdLBuLZssrZBeMQzFb9JUgU9H0YwQF
qQS8xR9pG+0PLrtlzKhP19S4pFaCzrHs73m7hOrZmRr+cpo0eBDvFP41q23Vb4wS
Ggmgg0Mzcjw6ETlEaEtxsMlaxyCPxWNlweFxV1j9jpeb5jnO72EXFW5HCaqqE6EX
GHJdj2KO4DRzgbsuCyw+W1YyFmvhd93DIkaZoHWr4B4BjO/qPsJhdeEnuf7MrLiy
0NA+nGAhWWhq833TZqmg05nDgV5d+Sl0ej7VcfEgJGExtX5nhasXHBYo3fye241t
XUZsQJ4TusofBFWkxtaltjgmJxvbiOBzBSF5o+pVcSF6spSGScOEdLD1I6djfGqS
VFGFYL5sTswMppxla0qzDMY20NjNyqTeJ//3QOc36gKCXbj88Jx8dVxVXi/Td0Ak
TXMJtTUz30VqpzhXLF9RYYWoESuhfnI4nrTsDt+FS/vvlzyh+9M+5C9E/7DIgUj1
SADdjxkLUOOtr35+bbHCDXfdu77vjQSk2hEAJwMGwlNM4/daoHDQjeJ4+L7B8Re6
tzQYCgyi5VRA1+1zxtv2MgHA1s5+MFFW9ABRakAk2wHIBCpvHn/pbutjJAsFMLq9
uCd3vsqGo5hd7tNCmo4r+dZ25e6ZDrax/p22T9whZuI6/wGFuUDIVbSrCpQNIyav
5uzDLe/Wg8cFlIlyzdn0bGcz9XN1Sn5HSCOVATkRMq6fncbajtGHJZbLkcFyFnMi
WkNYf/qRHqhHaMnwFLO+7sc9c/vGX0jVsniXNfxUy1yOqe2AOIar5mZO8Os9xMIw
6sAx/7r8sZ3QrpBXt4zOPSmEk6fSCVQ8h9uRrQ6tXt7MFHxBe4v3zQpYOuWgoV+p
dU6a+NGqDn+ms04cgukdQlCXbx4+VZkUwzA+2hA1oa9SEsZK5/YnL3tGtehqJbJx
a4UMEhU1+O36uycROEGm3rIEpkWsTYx6PO50iuW1P+3Zqks7IPsimMAVU8i7+GnW
+/Zd9tKiQ4BqYzkKbCnVi45n3rPeq4fqPpXdrSxjpvFJ9ApwrVKfUDGED4TpTloD
YFARZCXqv/sGb1sTv++chbgKR5qaaS8W2qVh6FH5Y5POHq38XQ7iVbHWX6l/3ID6
nb8t++s/lGnYfcfECEKLAH/rW6zBIQ1ISNO+JaGGEV7+8GWmFczKuKs5KWaMHbbP
RAPzFiTLmBl322mjhXfYaQtU9qCK/OblGJ6B7MOgLE6dy6kV48mZ5lgIJPZyhjSd
702iMaeVbxgvO4v93XX3hHJO89h2XYI7NnPxvVBrzfLWxCqKX292GKjyZwxExlfr
rEAT5yqXDGVB+tQae4Q77MP+z5MlyM2Yz2wk6Nmas0FRZsziLA92L+wmYBtjt67C
akgXIMWiinwwnFJEpjlzL/sPxeUWfpc469o+/ZRTkJfVFt6noQpf0RsTAXvaIL3H
CTHiJP8luHqr+xZQcCv5Vn5nzOKsgwwOCjEFKUXOUHjx9dbgxLME35uRDxqR4CKw
vkrBGQgPJ6FylKPgO5E1fMHeRnOvpJDvMQMwXNg1zSnD8aeJf0JvsT2YYNM6ABUS
l0jLrPC5TlDWkYM3Cb4sRIhn7g7fYbVmqfjWKnmTBT036wbhuAIeN2YZC6lNew3j
CfrBAKLnLpE+zut5iR9gUcKvx7pMLzpn8zHhwDLFU+0cPz0Uas4LbteKbI2vQd6x
sFLx82Cw9A0wGaKzfkhw7BUMnWo9HIkvtcWpSwg7a8y4nDwt/HawUhNafPTdFceD
QmFqd+CMzsJRE1epGcEKEyr+DcVA2FSUF9c9M2qSn3CYb+FaOMPORDi/piZq/EOr
SPBQ9ZgWSN45kblJZLdwz/NrfY5WgZ4oT4+KvZisca9SaTv/l0TxsvzZ6pl76K7i
GDKJKb1BRX/2vwnje71tuq5FrWMNujLMq6anIg82CFHWC2iXrb43ljhjKf/4ftrH
S2uF4ntyZiONe5gS+VbymccIvOeSqGL1nDp6W8txQvi9q5QfiXQf3Wiawl2SF2pI
V25zhXJHAl0JJA492DEHtRxpdXMNhzgABA3cwAI/4Io1F69So7fI5Aljd8/z2f1v
bSpgFCjgKVvLreD8CNfgOEqRpAKAc5NsaSUvBRo9v+MShH0SCmde6pBjEkolOo6M
v9kuv/3EB454iuMOgy+FI6zqFNmWhLnTFmtLi4+ubPR8SfcqXNN+wauBMBVe5Gp1
g2hSfJq2az3mRGCihCW2xfFkEKNP7pA+9vz7ZFivPfs+/6fT+VtYnKo2PZ4UKcUi
FVceBOqep0QveDioV7n+wjndlU5A/H28H8I8JWKozQMhlXxgahwl18mOOTRzcmJR
1n8fkQ5ne6EP5cqbtclUslmSzZ5mJ1cI3zlgvXwcLSnU65jvtbu2hYi1V7nf+qoZ
9k1BgBR6iO3bf9cJMrHYW/K/Uk4DRdUHthIByYa5uj0fDFY958mSHcUV+RHliHHy
NUUVmkL0PAhJyX+PhttIXcKdm6Y0WkDokk2lx5/lIliRScOI8MGgGJmjFh6wbUyn
imTiW6R4Pkbzij0CQke5VirNghzYAGfh4uuIleWSx88PWONNFscTz2xP6nYIq+YB
lQ+4pUTVLt7BqqIob7V9dsIye4blzW8lKa1rJCKtDwpnSpjBI0Geb7tuUrEsgHD7
6xwLlk/drrfE04aBKCWhQ+HzLypqaAN/h78A1FWfP8T+kbi7fRR0UoTCgtfB1Ai2
mZGtp7daDinrtF7uBtAArXvSOpK5/pB4xq1N1SSeHdxzet+g0prXUs04DEJc/tox
zYuQFccH2fZtA4vijRLnjCmfDjFDrB1dYs07rf4Wad59GVKf7pnx4nWwZHEhnFCr
5uodg+djEc9eUxKV7AgDro1Sg2Y0Il1N8oW/MGqHCyJJ0pmC4YvmxMheNuYBM14b
wZjX1qEM0to3nAAqsU+/gwJ/YGw1AeIOp8Q7YWlbT+nOifzi9utOn4mtBDWa3ARd
fAv50mn7tKgLzWkKdP7w/xAXUFVlP0PKPox/rSlIuFY0EtcA0mxpOy3i75fvT7JD
/PDP/iavxaoRP1zpdilk/GZp8sFkCFOOGpvL4aDwlEvqOrnAmIot1KDi5RlsjK/W
D3YAF+RIkbatowN+BVVVXPs/HuNDuCMzKzFTlvFmf94cCfBp99L1vCFOE5+OOEmm
my0oxbqDG2XpXCnMwFjgUozyHoL2zLCPxPOXzSGYEwY7gN2+rt9R7aKUv+KHS8I6
cPmfLwMybRm5uWDndH+iKIx88WBh0HYOf3sp9CL0WYj2YVhRo6jmB5eex3tBGAa2
kEJ8f+usp0UaZtBxbcJN7xS1d/uvuKzXHDBbIGo1KCktBhJiKxlLsDQJEYH4LhzV
N0J+j/uOORqycHyUobJEosfw16Vjvavsgu+JgfGD2/VNvOET6c94SnnIiAgj+6g7
knuaFJZGD4QECii+piXN9YYGcoSIc6w7P4B7wUGZ6sGP2em6iowNXkFbox1OxylL
AI3bfmiaYqdBmFmTVcmlSwyt1Y65PWrECf+Q1LmwSLHur8q2aWSqp9kFyzEEfoDQ
Oc2HedOsqY5dj4fNcvSAk5mEy3fjd06Z/R1fPqJ0oRHRVjd2Gz6davEyTGUqnlBe
pmr83wbO1Po4sSP3T8bZuZ5wZ3B/MsECMv8vxzvC0y8Mvc1NlH8RaKKex1blTC1Q
ubGxrnO7dVgAthU9puEm3aUT1KOLl8kwFxe+hzXN2kSVYIGkd9RAYG/ZXkE4dCvV
b/H92Pj9kjtzi/8nigqDHIJ9m+sRfo+GJWs81TbjyJbqimeZ0F7diQvWiwyXlIVL
eapWPyiAhKoMxc21vsjt/c3hDpjoq252jV7M5xL23r1HVZtAOWltLgIX7f2+prci
6FzM3etjxWNf5qC0bfZBc9lzOfnAyKHSLnhyN9nfehuRAFdJPgkVbVEl28X2ucVO
Ytf7GycaM/ixGK25MwoCmkzhdExmRBjGffm0qeM/ymxJiVtrSp3ubROg+3v0ZT4K
b/BbPzVyBvONE93Z/11Wog9r3tT/BmjQyw+IuGJr4pvjpjYeQ8GzFgn+12aOlu74
9YvVCkVKBVenM7cau6ZrognvK0qgXFRTyxjsnLKmeQRZAxfXxyZo/G4+exP5aiAF
B93U3V61JRRxUUn8k4YdBFH9p33uSXJA2hLExeg7ofRj1BJt51bLc7z0vm+1gc8a
+JaD4Mi5X8HDoPYkeMuV+uhTb7yL5fCWimUMH2+pFpS8Z/cptlEMydn6C/qn7B43
lP0bglP8jFSEd576FnsEjPloEwqfXBV9ZD/orOeu3Ig/skGcS6UlPuFOML4a+baQ
hdy1Ni4/49f/9KAN1/hePQkiSdFmJTOoPByOrJdRJVXX/XMW+yH9b3fstD26pnla
kuY8GEBrB3fTEHV8M0ld+Yqh4JoLZJlFVFSn9MVRCXnDApxKIpLEAWIoPp5PMX4v
BEwe7Ir2uy1tObp8hUrtYzlWrkvlAt/sR/xDF5gIh2VArqWLZXtx4M6AZ/w64VVe
1+MN3Vl4zpq/zII6ic1iPGtJMtzUOvzJ3ykerUi5bVMTU+cvZXDXlBjdy0fmXX6l
/Yp5h9470VAR9lmd9R/k9I46ICk7R5qfSwy0OLqH5BeDTnWsYuSlWWZOC19F+7zY
nPiaBmULWYWs6uV+gAHEB+FEC+iMlK1G0kgzUFep44Xd5z5e4tnrzDFa9ub4EBnl
luuEoSk1UrRgmLoFnBLWhpgCxUzdZNMUPiuZ0UCSGRoTzIAXqFPVuWEVVbVbOwhR
VtPBsvGAZho32sPlCCLgzJG2hzgbifjRHFe4G+P2B0iKxK/KQrAB73mgJinNWaES
ENLYCItPzdoHsdnHEu1MQB3R/O/Hl83WMoiSKMXqt214dazI7IPyjUMdR10ONxGo
XU530eBgeHLhp3BwvPDw1IQpmxIh4Kvkz1IYinFNffzsxsQntTbRGj/mU4HpjJ8R
0Y+dEiWsGS5ujgkeZ9S8Av2zmlIEMA2j4uaR8TzMEtMP6HARZug/GiD9FtZOxd8d
ob/lExI218j0NWxVnJzL4XNLC5w7yy7vJCRdUEpYRON7XnOQYhPrgajrfr66UJuS
LQtsXZR22vD9FeJwvrpMK9SDkfQUqCABDQSB+vhFqTfwWP6pq7fx0PzSPKxG6Oac
NBI9TnSO8bGt2/E6NDCn6CFn8uMrheabeMU+27ZTgThXbGYCslot41g1gzqlAvyk
BQz9V9OvsTzftED7terV7JtJeWnkmpT5ItnwW7mf4mQdVqQ+wLyR7LG2tAmvX/Bj
6s17PgYNNvseV6uHK6pOEY/BnBVJFrLcu1kuqInKEskqoCgjYIhZfJpD2xKXgGE9
XOU/AjTD7f+4r26qXSV2W1ABTJ+r691V4cdL4XAHQMNOkKSgAdKfF/3lWoFVm3RJ
4+PZ2sTs7exYEmldt3di74UJnctEHeP8CrZdS1003aeGFhjgH+ZNIWaDeNWUqYh7
RfhtjTkQL7doUNfcIscwvIquT+8tnGYnsBcmJQTuF7AAhsigvbWHxN0Di3uCHH9l
WaYhtrS6S5vvb7utI7+wltmRVNBcTtQLLne3XdeaPxrMLXgdwheLS5i4V4J7eCs5
0YqMyrdLE8dV1rM0GozGcMwcWKTTPTr80pqFdw3lG6iHBN8cLWMuxh4dtNBf9+O+
/cNHg8uCZWvjUuu9JrULoTrKh47/U4d75TWuK+NF3v8sQ2gXzBNlP2kBQkOjSwLV
n5O2x4tA2XSusGOqGZXE9uUsfrLY++p6R314JHZKmqeXVJ5yHJhBpUiVW8Ilab+8
QtZrvC7hqYgKlIUBxWdpdN3qDlcxDgvduyoJRGra3ZPFUsR9VkIhtRn2O7GgPTUb
HTuQfCXRdBkuITZJ2lFJ05+nNG62QHS1wpbaEAb/lAryDFdMjZieEhHTKFgh04PP
UWGomTq+bUTX73s+kujjRET2+Nm3td30N5jgMyOpeCCY7LYGxG80OVq5+CDHQO8Z
bBf13bN1IWl5b3pkghmukJTmvGMxVIa9b+288n16x8sz00Z904Q/AhxJ2KGnWvzB
GdRxFuKp9OknwlBospo7YPZMxjwtC77BkrbULgjT9XCDgJ72cDK8jN7hyPxTpUm7
ulnbH3Lqqy3dh70LLhJR8f1vNIwSbj5slvpm313FRh7MTJR5FqyHRRPo3Bt9LgSw
j1OBZ5CM6NGVJcAwFG/ydOdej91pVNbMPFQvYw3tsKn+FeKA3qf7vAxN3peuUky7
R/MhWK+KixlUUd1P1bIQkjlC4PCMp9DZQnVvUwX0m0dJ8BD3GG5nTobx2H5Nc0Xu
tm0yA7Slij/8idDCcEd2jn+bsC4xlbGqx4Wysn9+yEQhDXfO7yG18ClesxmAweI1
yibjvpwHG2n6zCJKyxSyZnnio/xJSr7/OKxdHwoSd1yvHd9aRTbAPviKzyVj9AYD
q6NFpAY9n1JNF5KMtGsIWh7HR9oEKDH9QdZ8lNI7t73Ga+1dwcOuX42L6Dt30sW1
wLORG2noAPy2W9+fKMBzkVzo8s1bUZAUj+Z1HEUkItGxW3rnN2VHE9JubnRUpDLL
/eeNTBZVLhOYLNzZaAvChe+BptTNZw5ILVSCkGNYBKu/14xOHHLlM00NzT7hyqQW
n6dOqynK9pxq9nbTgCMynjUEwWoIpfmwlrhNhR90TS+0+xrvvkHD/WbH2iJp+r9i
7WLXaVcFZHUI6ebtXNDW/HkqVy+kC0YElfoTUGBC4r4euQ6sJaFBfLcHANZk7SAp
PUN3DUS3Z5Jav+f5Hp/JCHQiYhizHG1zJM0rX6Uwa+yw56gAmNhLLVyxLPKicFgV
xzM7Bd+XnLIB3RdOHlD2qAlwlSzvpZwI5S7Etln+IeIEgJyNWwHiVJLAwBJdJzZr
+5ZpaAdLCP6veX5ogX0AFr3Dj6WEGPn9pPYbahP1Wdu2164u4Woz2/3ssRDCy/Eu
pOG3F4DMoexEeaS7xWN8TQFGVnuuBqSsVyEJlaZuUMJug55BcDZw6IazkXSsNAvO
bN8vpjYn+LOo3FtCKl5xcvXJACKaaB0VyhshQ3tpvtJfEPV1Js/NElfR0lNn6/5S
TtizlJZM6sIIRvHdd1SJXho1mGrInL2JGpONaNyyhV4rniFeMA5K/rDXilTPyQ26
bUl2ayKB5O2DXb+9PAnLmR5zTNUD9SiF8eL3JX7reFhegqfi+ArXfIATzu1KtUGj
AnZt946uLt95zWqxBxEr8X4Nqft54qt2bzvMCcJvD09AyzVG/lr15t3xyu2Mgcv8
bWVMxG02Fo/J3czdl/nxQqeTMd3wjaK5t2G52sbOOr8X1XJjZ+rux88tTE+jWjEh
raKZpFEJL1wIZK4og1+GCwQb8aNSfK54Zbjyv3OBGnENcTyTqzzjJgRxyIpBwvjz
FkFTNKTUs4Cwlt4VQKA/OKI/qBCNZ9CdUtl/yY6IBtuH1CFGV23uze8xa+7QiHS2
4SVDC6atObmtWBgYYiyThyEnJ7iTxR5Tq+I9tRh+TZ9saa8ZSG9ZWzKlE5IDuVo/
hG1qVgnhywAax5xa2gkvUxgJcBe2NSTNeNXVzrjOf29Nb0U0mbTjNJXNCuyuF7hw
HUDHqWBSx6F+bZNmJExGNVlY7+62WH+LRWMbvCFQSBdeB7NvBhYGIvgYI1LvWhU6
z0IX7558JTy2uwrB52TZic1koe7h/3Q+bzaG2TwGwEGUXc1IvcrcsNN6H9EjDy//
nZHFwH8rjd9S9i9SFjIL/LMBsodTt2PgYCQb3xXnNc42HipHa1J9zGToVMfY698w
SHwROXyr9coVkCjgNBJClLkLJDtZXmIuJePD8MGn9c/lySaw8fPvx0QCTaSWmnis
MkpsAxlD19iaowcGyMS0wywpovXY580kL6Z1PBBXz9e2LveEcyvDhVQTxGltaPjc
kbkPMKnZqPWhYc2m7xFQ+rYt7KmzLiUAksQ/wM4MNBag/snzScap5IaEM8ZzyBGT
gpBEAJzAFLlqFcSAAACMJD1XA55eN2ZE8/HydD5Lo2YLwXw27XKOE4gLTKbjQ1hq
Twuv7eg+NGrpq2kCzB0nRVeAtqS+hOyuVqCcHxoGrGSvtL3S8DtE+LeQzitOEH9F
rjNRLd1i+oSeEc0Lpp2NR0OLyzTVF8JqXT1knf8tkx1jCYsp7j+OJJ/s2od9jLIH
pi5m/XRj8u1z0scpJSdwdr3/ZxGzfs5H+A3VJmlcD8KCSCpyKoTYX7RuA+S1K1VV
IJ7ldTMxIIuV06QiQAtFm/8cb14EmSt/mTZyWhSpdCLqbUKqreeVjkq+FYy8ympo
A+80YYHMENfEY1IR2FeuD8m270fIxzTbkPcI6dfkbFfwryRZLdJEqkO6GUjkSFYJ
7WhYbtMB8FRbEdyL3YlFhnfgC0Hpvi+eu8SoaQwvo83HqK022UVgELYlE9C6rCYG
QvY7ySJ2at1cOZl37m1/I+47G481mZ7yo52k7uORrfYWaITSxM2kjM8E1ny97BPa
42Q/jCddi5iyvkUN6HVtCDDREemw4Nlvk6gCw7/B314GeV0pQVHB1VyVUiswdUpH
jKZOmfhWDB1x66yYraNTBYSB3yb1hady29sP0kBqNWxsLOsIcFraYCGQULIRJpxW
IuwZ1sGwxT3lWJrCpy903gFlcmuPTGDs/FhaC3igG7+HKJ/IbZoYCVAkypmeiqCL
2ONgBVpgIGPy7QVmRmvhSRLi7wj9WoyhuhiJNb/ZSzHC134ncanOIUrKJI1no5TE
Pa6z9n6GIdIZRMACRBfgAunSJgCxMw5FZbAQW0vQSiiLrvw+jWo3+sUAqh1h4zcl
Vx1WfXRiUc9JXQGXYm04pOvkSYcY7jea9CUO7OZyv9B0RbF2S9nV6n4kp1j5myEe
7P+N6yDKrK1D5ElrTJdFHAnowDKdKnTfQqZObqv+BscfPb8m7UoerrdljddtIfNU
8QYLP51qPT0DTli01b9q+PD4OdngNG0w8Kutnoqj2uUbwuOc/KIscjw8vT/xQbxT
6BVLDwgFbHcjDi7km4411XtqcPz4dCMA3HZwWEq12PnI+2UB7kjdUU8RTUSujk31
/Jbz/EoZVBGTg/fXEsngV1bGSr1J/IFb4J4XXbj95GlsEeCjUNqkl7xdKYvNJ1AT
XmMGxTxnsvyazby+6Vo7h7JJN4cMOoOgbxLIVyFCbXj+LgtFqS1RlqRi4Wkai12W
IkDj1gwGQ5fJ3hrDjsOpTrBrJL36Ko8a2KHAH7WNr2W90lB/FNhPdaDFfSp9nzZc
INpzMY8gZl1sTFYH/BrhpJrdAikJc4KnwyAAbDCPFvYdJusbkhX+wFNeeP1vjhuH
tOMijKTjssBDFyyHdj11A7Cx+JKUBm3sl8u//TvNYy/Iu/EiYVGqzxXFp6GjATzV
0r3MpM09KpHWm4f8eQgFa95X2WZUMcyl1JCdiagc8Iml+OcuyRk/Ghc5FpC7OTUI
kjLOrTFHOum2o8gHyPFQ0IEptaMy8V/QCMf2aFIgB/HZX4jeKAEBLtmZBszIJoJ7
UFVhWbwqiyKxEr12yYmgrSZhR/Ybw9S6ZOZzF12VLwKUnd0lW4hyHB40WvFwTUJr
0JhCPx0S47033C1t0rc+Q4VxOniKJWfVa84koqgOMzutNSdGXr8/bKsUioFtKJLD
nob7rAOLWp2W5bgG1bNEJC0LkVxhuczbnli/yhbCodq8cqpv2fBt3rFVhCBHGzUx
BKJqARAstql0n10Xm+pbB+rWQBxoKRruFAPGCRZjo4y+ft/hnCQDPmWAjk+7EAI3
Pau7UWLTJ8lMy8y69b91JgPGjILNuWG3HduQR9kPDkkRh8zy9y+jyVq5VFI9waJr
tUNniBeErl6X9BK54gqO2tbM8IkJh16DoKgj8r9JKSMeWeY/3iHoKQ/SN4RK+jPV
G/F2b/TJjBWoYEujMIqzKI2jhK78b3LGBKKrJvH2BVJ22cG2MhjFeZU7s87Qb3RQ
DMSz+W4Jyz3WafERss7d2vuecP+CASNKVuMfd3KVraGNoKctMSoX1CQS8jnoZFsZ
NGsOX/ZlTXpCwhPmdwH1pFXfFRxN351uzPFglm6a0r3gGrOAl6nv6j6BvAaykr7j
8oQMZhyvzha/BAz3yUO6mQDvMfV2KCzC5zDg5yZtk3oljQRHmhVU3MIv1OmEBk/S
Ab3BdLRzZ+J0AjTSlxE5H8t4zN2sirU1tvhR1tFmUu+Hae7p0oKTXYAB8nj569J+
j3rvK68S5r59CVF5pI5Z/+xCZnPDi2D55PHWI9tDpCdfDQIWGGAd1FGsrGUIq5bk
apXDuXr9mJZvECQwcU64BoqGCaI6Ir2THB25dMl58pOAyhexbDF5E/zV9pSZ4Fs/
m0XQWiXPRH1cVdK94/nGHA/gAo0HCPQzYzjR8fZ03/t0vuwlwbwjpF70+dwsKV7p
cArcTIXeKXeOOTT7rpxlzH9wtiInWRtmHqxvUzkptycX+FXljPxq02cnwPOFE/VS
FMbLvF096hghEveo0yTozcyy8d1aJGSlO2ns9RDINt0mxx92vXFWVshSpDQoLHEZ
UIFWjMg3SilKN9lrcBWusACOrIDd0Xs9i+bpe/L81l2DIFX5sRPGVTM64ogAjUqC
Yf5/GlAmquwl1rOeSARG75B2T6mq7e/8Xl/Qxxdr9H0gQj0f4ScgEV2nLQg59VAx
e4XT290iG/sr82sMY9A43lM+IqVKVlPAlwpPTaA9OeNpPD2LKNqEEsoLRVi3hvvJ
l6x3g2WFs2x9QsgqIpw93EJcu35BSnVax0OBynGBx2NmJifvA+tju9ZO8DjgeDJJ
u4nuFoD63obGsqhrKRLp6k/iW6//Vu3RsTr+x0WnWI0ygvHgTXA4DS59+SNsI4Nx
rbSEpAsJI9OYrxdKjSXvqdfChBKh2oeCkdiQZUmZ+LI1VQ22LiD040JAdakz6DIM
hU+MosD92CAk1TjFEcSxs6CyxF9b8aSA7Tp79d8RXJK2OnBnUsiLaAT1moutn3Hk
pVY5qO4pbyAsvC4yHnl4q3xeENtvCsaQHi+pnRKZBNzqa8uGVYTZ7bRFcT0+CZ57
kEG71z8/Z+zp9OQVnZ8HZxasDs7DwN11TLjDZHp2xp/clnE8G+vASb4/wXiRDxzp
KO9FyQGIGA2cc9lZIndG2kuJmZQHxlfeT3vlFRouJMINzfrLOtkMjoS0uyY2EJvN
Oh1ouqNyJfh1SnBAd1T+DtixA9Kp8fFDioOQLJIrXWV7luVTyFneIuygvYhP4MC/
8QUQbSebQGcljFjzZLpfrKpWszcR5eszNYVxJowF6kPfG8M2Dgwmoky0lZzVX9cl
g+9L5iJNzTdkJTCW/FcTIwvufYsQ7eYyCPDOLy1m+dSOdtV2pEDKwydaH1pGkzIM
pY+Ogxi1ZISFOG7VhVPve+KkXSWYhJOfl83ObGzQ+2U9xq8pMUcS94vz+k2s85pJ
HJ2kkKq/79VgAlkzNQbUNx7zb4OKo09APP15IG7c3NfSKaYfxyN/dxdaU3hIBv0/
p2WpikkU+xJl56OGQweDF/pMTMUxLJEU3+Ja/jC+uQZeg1xwgQJmEw59lMAznJAP
SVQLH9ZXFY9I9P+3v8vdzrcD20tujOArKgm9nrPzpvmydB65JpGtcb1CPSmYbZJk
t1lkP6PSyTjgcuL+qLzVyRzVMqgOpNV4kzEcnI/aB5MVVX6GmaPztrUNvyg52UyW
DsLX5xcOc/Uy33wpba6eYlA/AxGv8fOm4hmMJMwVy8E65ae2owPrpkCPCMSBP/Cu
r/lNnTVl2u41SVVr117qEJZ9f0yHzgiUxKZNO7HENwOlVRb4FIgjhZdh0BVub/Rg
VKmk+HIr8AkTcg+zTgPwCniwcL4XnK6lKEqV21/wFNOtHxAeWY/cqHMfI43ugxbs
VfEfi+O2hZou9xJd/nlRnPpv3R+Izmn4jOr9tBJL8PyOV8snkHELFtDRERM7c8pe
dBzNtkITNVnjgjhH9r0fBBr40Qly8gPJ6wgKhfxy2LjmJdUyAlj4b7ZE4PzUcfqw
rsRLvd2OcoZIJForwsoDGjq8yEdcmyKYQURzrvNEaICq+niyAsDmo15dfHMVRETV
gNuUTLvHwTBKP6294gPQUHkIgpjhDV1Q5XqNqeT2jw3MuE/YTQpeTSP3/HIhGkMH
S8HlLxk65zt6KkYZlXVQqaQWNraYcOiyYStT6xr+ffWmBDuW5AcjX6Yv6HM/10uu
koqCdmTTXJbx6ZKXZwvSbKrbeQPwKkV3vgNaGGgv+QDSKlgzWGE4GlXP1uaSjH5O
GYV3nKH9JLc6uU8Kavjg0+iOtEk/Qs5bhpytNSPEgZfiqhf6y3fvWata1bRiRnby
e66YWhllwjsMku64fJyKGTfYzjev6hsrqoXRRwhW+7usosMy676mZh0Sjfvdi9CM
N/lLwZC70bnr6A4ALo+46arZdLFJ30vdySyNA0CSzPJwLOAzZavpE+/NruX8KZuM
oLmNNOnTmHG+bZx6FxpSwx2VbDvLfi2AG5fHNOhTuBHoV1LuF99LSJoCzXaZAxYx
NvXmf4g1+UYbS71R9mrLa+oxsmLLQRLB4Uax7PTmrIMgzEe+ohqKfrfkXX5NFYCp
bbvJ7dzBGgB+kGI82UV9sirHUwNx5LVjXtwA1gYY8iZjKi+775cvB75A7Y5qeEeQ
PxWMEu9oa3GEGjWf8sU4dlRx6owK/IvMtKJMu/xtVd2vjyhFqdSIVKATGW87t8Wh
m2ilB+GT1P988K4kO/zGJf4Cg7+QMO37yKku8FVMqzdp9EMa/luvH+6iL0yMONPi
pgTcQR/FmzSfm/iRaYPPTmYdnhWqKA74VmnFcob9PYCLGKQwSZ0K5MRYgSUtW8YP
t3HidnGUVXZpi0jqceDMYF/5IfY+oF8Chwn5BfQuptkRgMe27GgZjb5jDerrse6h
KG+eLwgmZKADQqlsRVYnHVa1SKx4FSftaYtRTSTCl2vScF2Y0Sgccv1qHW75K+fv
XCWPX3V6TGBLYT1Y+9Iud7vVGIBz1JMq6Gci5pfvS7wEuAR26bcFW0YFioaz1NiY
eYwk4FE1M0DI/z8jF4jBd5hOedN43glSrNCIDH8e5/QfM+1PL+/6bXH4IkVMN8sa
EGSBNCIa8G6S+Yw2Vu9AQNi1EVKEZx0ZPeWLXQZIgnOgz+U4/weLD/I48JhjpW9d
d+yJ4soF06hQeLpE+QSRQCKowG7BVSmgXd6xsi6IzJ2lVghZkIrinDRgbYDJ8AxS
g4qY5l2roXmE9wFHnx0qlrTc3X5e86MMLWzNliQchfOIZl01UhYw8MMgS7ai3YVM
LOukYr6do6hqB/XV2JraGzKF30zS3NsO84DKxQKgT3v9NC+HX6DOUMQ+LQ9U9wmB
EpEhN8G92obriNhZqS6DGGxyTZ8QLabjCw8ll86MZrcOdfd+uT7NNqHrwrcGhz0b
G+S3nKhXnxRjE9Ne7rT3TfeefZQH5ha7QHzB40UlmZESzGMeo8h0WOpXzpOuQzI2
j1UdgG61nVDNNRSAsGe47rZPh1JiMcrNDfKBdwDUajyIDZ1QwSl7cRp7vuklY/6T
7qsvNKVZuYz56pnzMYXgjzQ9ZEbfO09qUgQtXfu1rdHVGt+ln1FyR0acRbvdGc40
u+3aFk4L3xu3keLBgRUSX3WYFEBxetkrwoHqFqveK0fZfCmZ4VMUVKEkFm75Hl8k
05FMbY1lLliLP9eTk8H+KFenRWp+ZOx4FzLuL/4abcD1MvfxarKZ7Ybhk43hnU0O
SWrwmIGD9antUpb4ZjJ1gCzm2Qck1zQ7Vl09U1D8Bku+FifsY5k329P+ZXla1JoT
dNKQfrTWiBSQyyjfTiVjdYgJQNggorTy3PMCtXNvZ7UVb6fE/vSj9hCZ6MtRSP3g
oDWoW7vDhyM/ZcfkjGqQZ+3fngGwnYjyyQoh124hDXnqtDQMUEk7QdmWfSXjhEDV
JFgjj4Y4NgwpcPRavzcZVo9b0w9w0yBl7aLN6yOjcKElO67tdeBFfhDOPBSpmm8v
VH1SM/zwMq6KxSslxl76vnmD4G5pvlK8HZ9zSJgSpuvwkzrMv9B3g54qoT6wFQhn
dlmRFnY6DszLxApZ6aymIg+2KPkO+p3LvIx6pLEG8KImxiRpwOgR7AUsulzEXQPu
95/r5wg3jiW+5njHVAkidfiXutvoIeXxcvUCmmjNAgv4mvwq/G3W4PdF1HBU9Fjw
hPO8nuy9u5v8cFFIbOQzOF4NTB0GeM3psbYsfLmz0LNgjmsP3DL81Dk2vsxw6sFV
48wwzLKnWAJFyR/0UlqAo22xSgvxIbHq7l7qWhxwPS2ygy9PJ5Kf2qXYPL1xOIEv
g/YEdAFP06BURTM/S7/zIjTffhjV6Fo/9BrdmBSuxfzqP4X2vm7DceapVJEtKNDk
SVV3Bl8R8D4ESuKqR/kwESs/xRI+7gjScl42UHyJqJD0Z0GnSfVhbFyYf9Wq1Kuz
NWu4WFWjfVetcDzKpBNL1AP8ko5NkkJpF3KBihGiUHa9CKendVWCi49EcU093JUS
LvA0x4lNp4ZbFe1igpXzqte5w1Aw+37nq+OW9QGDPvEFxRjdcSyONE3+8mC094cK
gMiXcbhXdaI5zV51HrjthC8jJf6YEU8fKbzj1sNBgC+xZmxXLKT/teARZTrop7UB
YZumptOtSXTnNr4Y7u150BOLfUii2SV2rUMSRI9YWgh/3D9j8yPaY5GELv0h2X5Q
USrd7DKK4pTlzajF5TOfG41E/JeXmt3m+9Fpqs4jGIZawkjp+yTSjjXLBO61YSUF
xhqiXifIG47KglPJLkVJ5LKUEf95XHdP1e8EnfqArZXY6nKe4OiTYZzD6rSpIc9O
qyhcPUKcqKPj2EXIdHBNQTTyoxajOLiDZX5b76jpX4RTFotUy7VyydjnB2+GG6sz
smeX1GKTH5XuyJDaWUndzCsvh7b0FNbeARIjfahH7VElPT9PsCAiRjbPeQ3nrw4R
yXNSuSISXH9HyEVocynBoDwfErtqyZxWEWxKaaHbsufX6mg4sY+9FqbqHuW7h0sH
O+x1LC6b82KmO/N9EPk3ZryyVGcOKxyZdTLnnwor77dRINpTzxd4VUDXSAGdIve0
nGa1Id8ztx9CHW+9wYoRK37yDqIgCK/3A5DWkAC+97p3avx/WuLaywNJzekRGDAF
rs0KAqr4SGyDdh0fKEUVaes2UTaXfdpo9egnHvxSSMjDzu3N8bD83EMZ+PAIMtdn
N7Dwetq+8uhz9NwGvIEZOG4Xxjfr5xt/GtEx1DEBNUx5WLwnt6NyiwofSunpvI/K
iTz+BkUrrRo7L4LWKP7QGVJqWTQMyx/kMWnM0+kmwDcdlTamh2bzDUmMvpLR6Ddw
TICALk4NJJO9dNFIMcOhn9HRfvzKhd4Lt0MBtqQWqZR18+/TGF623+K+Hs20yGJn
IE4yIMqvTeRaAokXwTfE4XPOwUOY6NyqX5TC5IOUP3S0BR3HaR3apNqFTgmf79g2
LfS+etloBR2vtHnD8caWPcL38e542gygOYiQZE81KJ2gK1WzMKOGNZQxdDcJZ0pt
fZcNQia/jv4so1TZmsCG6mYIiycCJFgBXuhnQOKBn5L+0rCRkmwOSkF1NOWWT9I8
v38FggeztU9ETd3BSC15ZttBJd6pG5RMCt/i8VR3C8xq0my1BD0tXYU6CxkzgDDK
+qBkogxkzp9TVhU/3qhe1j6lkH+HGElGIAGdqbNyczoODiMIRGiZ8UEjcZ+ezLZM
pVabWniO0U4CcL9nC3jZzIg/62qwsUxmXEwcv+2Mnuax8QSXZFifMTcaj1EaV3Yz
c4w7GDcWUoNbuWXSO/txvRa9b3opmYk5oG0iWmN0x+NTi9p8uEx11/HmUdEFOOXp
NfN8tlwhxnPleFDyqTthDeWwTM4tM7+leXiIpHKQt6c8VslM3C8oNtgxUdSqlgNz
AJxkOajr71xqGLLjKVq/5HWTcVYtvE6xMu6a80aZNnKv+p58ZvFkcXfjvUKecfEh
aULEIjkaG2O0oexZVIsLjeR8+slpB4mNY850Vtj9eI+CxVO0FtfLXzNx6wqreM77
KJ6agQwrVk3I4eELc/j2CnXOl8jOURE0p98mTpCcYuek4L6azbSMaYOcJd80S48c
wXfspOtENrKz6xtCXgLpAoI1KEvZNNb+QBJoaVFV+4aSJqnP4AsNYprGGXekM+64
JnKZTQBLDo6oiE58f62iHnMsjvkQJ/CFipnxbGIm3j3oxEuGakroqFkfauJTn93Y
i7zEXT7E26YzLg2BTbFvd8QTEYS4QJDJLo7ye/M/xOvLNX801kwBuaVoyfmWlzdo
YPgKaMQzm72a2Ed2WyImUj0hJCh8u0dnXbQnzNUWSa/H/43r5lU1KvTIBd94zbsL
4CuTI3nBUWB3R8recxX8e4YJaJpCwZ2JJLbfCYZP1S+oiI+8AnN4hR6eOTERjzkS
UAgaGnE6YVOAEw83GjSCqr2PXp6SdDPA6zhJRwmeIwVqEvGqa7yaIFz+tmIrOcPE
MUeLCkynWaJh0c/rvSjiRYemUtHBj2/Q9SjxjV2aMbIHsywjAKGD6oO35xYYpzTu
gky+UNcTUPMckP6tgJVeo+8u1b6Hkl7Z6rbrjQ8fCD2OWPjKeUROsh71LgDM53FE
5FDVO4nEOoJDn3OJrVZxHieibMwTMwPF9SteT6GYIJPkqJJ0mJInYGbFP1BMWm1P
cYKVS0TwLhWOQngJkrEz9sEt+Hwl+YrIDaPkD51zdSVZdmr3LZKmq156zV5dpcMg
jeBD/2S+SRrOk7LeFTGlWbCwlc9ueie7EaM9C6kFBM7SpW89tueqRAjS1PnTecGr
v/8LeNqs0nfyRHo9e7Xvkatxbl1ebu+a6vSXkpM84rvOQPSpeIv/yF8anOmk+NOn
YgEOmRWQ5v8vbdNBEqIzmBXCXZllueQ9S5q43LdLA+K7fL5uriFBiKd4oJrKOd07
trtKapQmnKw0Avwi0qp2I8H2oOkV5ylAS1EsHSuwsmZZWmMiKNx2NyUiQUWaFUha
2IdpOxshVNrzZ8cz5S+/j9RQqyO1ITi7Zfjli4xOhCEGK3E0umMcBIJoPqks9M+y
tUTTfMlkK8+NDH6bunqX+Ygqt/jXB1cmiWGVUr4LDiVFg45jEvnT4yqgrDhLRCNY
CVe02WM6V7iau1C07+ybdImzizWOm3E+04flgy0HedsSN7WXBCopBXtcZm2Mw3Hz
GRTx7dEcQtdfHsq5h5i6phD0bMhQQXsZzloPsefz/v6cMn3e5K2JNH5LdZTt0P/k
v4rWDyX/lmAAHPJVu2bg8vRgh7T81dgdbc+wZqK0Q5zn3dwYgAyB161tqB+19cVL
Q5fGDihvDbAF+zjZkoajn/6tJ5H1zVCqrT6/8yt1tmS/9lHktOKkvBTZCTQXaLSg
GU1h3faajCLLikokOOVShTskv+EgrwDduYiuZGQegu+Dg4v1oyYanjdVZYpsY+Un
/Dpk7KivLFw1mz6gAdYd9f+nQKUmhIEYingky9JBYww23m70kJDFJd3ikZCvkxyD
lgFqfgtRM2DsiWLz3snqXqS/JalUDsyW5AbkdAVycGvYMRNtZVjAeEi477OA62Jc
0Y/2xD0HefDxwEVIcR6ag/4KnMqGZR6fHXp8phxdeOv7voCp6Oe2aMcSEXtL5dN3
FUp8fsXHf/scSrpVdTIkBXz5GQU49bR40mjvLnh+1vA1CSkabmv2I6StVniwdmjX
3/8jbapWIu9K+oLz7qgEceKynMgdbBkiHBg1RrQTzyKkwDdAAEPA3UgFXRoNxYIU
O1kJ6APxg/PmqC/HW0X9tx7iG8R6HgQ8E4Q05zB5yQK9/bUymW4oYp2ZLjJjXJkY
PITvb9i2Yso4BsqzHMt3s4avURa+SAUT3MAYALF6Sp6J2xoXzq4is8sbJ9bM3PBl
YmD+3Vhi1atOYw34XMG+PjVjFHBODTWXF7ejTOGqK0CYIlq8/hCa1QoaRgUFarCh
ymS+ZHZkEVgQ8/y9cM/WGJ/ku2jtgJZ6xlguhGHAUMZGOxj57fbOfb+UZVktxuBQ
xBjuZGeizNaTBxE+BCfmKTgu6ui2IFwGT9zctL/508L+hxDld4kgpaGDBEpHNv0V
7UahGHQUv2QH+ko8yXbC6eNCdzJguDe8d1R7/DHTp0PhVhM7UksgS8yOm3Blqix0
fZKRNm9pDEtu1qHEl5dTu+IaRpURXQkllDMD4lR5CSP72sfunoZR/PoP7+lE64e/
IufmWa8X/VSi9I4wY3s3ZvRViWck+G3+pznXDLICughKTwBqNOeIKL03hvlnVd4x
lnJ92gs9Dadiheg5MU017cZF0ZtLlVo4rbsjFFBhqDE1IFyty7unCR9CcBwSJ/uO
E1VInXWPc175JATlX6YVoZ+1ZfQlPzvntQPQ3TkY5CK+ZBhE4d8MR9plZGyWtcn5
M9kkgvojcw9W+pEz3ujr2Phwn2Crd9XtQmaa4f9cFBcXLqh1YFYz+MMNvYYlUFZv
y7wnZAp7UqxcvpMQjwfPuoqqmj57GR++4e5vN999LZx5W1WdqnN6i5preZ1Sg7Q4
4AFSsX4Yh1TnAtehXCAIqK6Wx9VJlFBJp+GgaWzRyyQpm7wDk1kMqWEzAeT2waf+
CuHYG+LHDlWkY2GxXoPAcEFOIn+wyxn88BRQeFWjtYXle7fUNu7SYa+NDNjRE9dC
HUz0Q4H+etQZArEcHZaUVr2BWow/uUYDWdRbOcjx9zDI5vCI1z3DvPQW4xEN9OPc
wKN/ABBYC8uygHEHJ7CncCd8U7jtt8TjgCj2niDBvYeTvPTQCdqXHAbV7oi6toC+
mK2siCf8DSz2cyAMdCZZTCm88ZOCplyQrU5ccpANFgAXfV1/WYD+c4itgH08+u7a
+a72PJUy0G7Wfe5bXtMTcdP+3LoiFxXqNF4MQ/k4UQY7BSn98aK4KnV0OLuwxvQ1
I+XccfukT4UBM1lpKvhWfTpjIwsyqx6ovZZgMjfYT9dEX+ScnYnUkAfPlJH5Tf15
PmzxZhOTr1QwcjiwYpyTTvONqCuVeP2H172bB0FgMxshfR1kGhmSil3UdqhSHFI0
0xa1mBfJiW3pBsCQ7r589d16qb+zdIgsxAMxGHBcpcGPC18GTn+dxUpuZjnt1ckc
9dGJfxDGnatq3/p+FE2rFfLt7NnC0tDWlxqStulTVAaSXPgmfb8u9h9QUPA+46J2
h708FbUeOuGuqPWFdHSrq5MefcWDhx0xvhFLA4U5+bwIvwOEJYdSdKZOO538Sj7i
414OsDZKF8jfbMkM9ZUOHf/GBZRrTCqBfeD6slS6qI1vrg54pH1KA/bsc8F12GgL
29YkDrS65dw95OO8GVMDa5KR9B6cS4RC7UWvp9ZWO67cRW+La3JDLo3IVXwEhUca
gU3E/L/6IlXqQCICs9zL5eQ7yvQLBhPGQcprQL83GKv//jfr1wUYrPRZ1SjmhNWM
ASzPFbv4Z+nMEZX3Lclj2m3NsrFB6j+wpY/Rx6zHKpG8cRClJCvUIcyZvnlChouy
di07V6sS3jB5L3N87JpTflPNKxYcexQhtD+1tikYCyrVVGuzpAgPi8BFtOF7eZc4
vWG9ggcCN+XvxO4nTBMcDQi6N0ed2ZJ1rSpdbe4UQEcgedUwQNwC/6PPJ8XyOLJj
J6m0nekyOzjsTRldNH6Nuj+llTeSBvYY89GnV9JAI50/qVMLWKnAL/9YKJ1lx2r8
E5RPLDMI/i3nphvzF2CypfDQbfXhKcKXrc1uh8xflf06MDcvvnEL2SpgDSk0QYAV
BT6yQyKl9lmSqBgPGB6D5nDPtlUSWpMxuo3oPizn5tbofl77dWFMQ41QMR4T0l6W
2344jrPQTC3yn8h1FIuTOqK1sjzhtBK44UO6fIIc+Xuj/K21MqowE6Abrq9u/gwg
Za5panxLmlAsYP87DJk4cVa7UTJDM1e3UqSg890Ry78LsbQOzVk4E7WiSQ0smaaG
wCbuye5WuKQd+uDBeEgU50iMFUdRhRpe7wSmiHt04JxWWgoVmR5XTkladYadyCEf
e5Hcy2jto1aADypuAqhSRanzo5M4OyCVuUaY7/xEm4U6N1IPe4CVbFM6d9tFJGIB
uKh/QxtqenO8FSEdiveockZN9vnmHAyW+CVj/s0yrRiyXfpRo0lBCu5XPc2X+upz
9yIsyMvMYK4W3EEpw8824jvysYnOkvwGfEbF+U5iwEEkgy/N0y1iX3eJLvYC6XrY
ym4h+EkElLRhAclNb4YMcIaIyUaQKwDk24uXabuYunRKpVdjH1WRUFRqu0Py0nVN
DqfXPVFn5TrvSUhnQrUK9zjwqeQZc4NdO93tJYMczttdmmruA5N4qjbjIrV2G+fR
GMg7EUeV5P4rGKn+CePIjWizAI0fWsMi9v9H9zeM+UfXixtj4Fz2wFfq4acZzORj
Z3EvcHNZw0NTGVwvwaLn0pvQnEWcDTq/SwGUxsgo5yhrZKGMGWHh2+b3yff5T7xG
Q9tjuPTqdssU4zGQKdRB6qAWP5CJxkTiJ3LxigyWwa0SDUO1qaaykUMMoPaa2065
BMUL1OndDeTWboYP8HLTgxzXj8tiPWBd6aSzUiCACQcdcgn3kxvhsFvWYYm91xP8
huxCQ6JrEa6L5JH6+8OYmoAWLq0snqegyvGzb893QwA4bIKamT9Phy4uPGYsR6c3
tRy4NWyL4MaPfdNsthDhKg5gAPU/U+jxoKcwe0kKZ+0QUuriJLRmgZoHgL2EEvPo
Lc+xA0e8G4eH2ezJhtPKAjlW+A+eavbJQMvqfsnXCmDG5QAeDQh+FSLGM2sUzzGg
UmTBSGxcuNfD22uBwaNjxVjnNeYOg/tqLUqxXXgBwqXHsIbs9FNg5vtu7uOIuYfc
i/vj9X+PeEw4n2QVnFiMrw7fSkQDYcpLaM3UKCbgaDIFsuQrd5heW1dQSv85VgpU
h+xk7lNGNE01Sj9AbncSiGnJK9pUTvYfD54kXpJQChhmkr3VfYfmQCFNbdcehtz+
bbooA2LPQdymLzV6Gd+jjy2it7K+AUDE0XlOXjoxOlfGG6zJa7xWc0nJX6VPv7b1
SBaSelv+cPcnrUSzkvh5AnzCbuQjx5nrA9RbXdihHb4A76ZbyDKi9UhfTgB2k5Td
sWjuENMck57wNl2//EJBSFGmZG0Fm7BWIZaA8uVtdC5jWaWTtG/UP/CPEnv6bFTc
KrA8ffuiAxKzWiZTrnAYNL8muBikjv6YBRTDuwc0WxblwiON9oCCQAdTCPM4b2Ly
yvHm9bgNXiD2AlROyYowC1308CYGOk0CBYsyNuEYlKHYObdbP/FHLGnmbCpYNwPF
FxrGf7zXurqd2xDll4hoIrZt5ERkzRC8fm0AWltEW92E7yTnM5lo4LDRpXu6j7TE
FCWqinpg8ARIIwzzWMpU1bePnXQYtfX0qTBbmAqHUuq9pG/E9wgR4897vbQGI2Ei
Q4jlW9GIAQL00IF3NPXTLvn52nTKOtRRNqYysi+BL7+cMj3xgNqF7lNd3q5kEIg4
z/7TZ+QIpFwLlQMjjWd+7o3Oi4ZX2PzPNbPHZq5RA5MK2a8PVdIvniL8wHtdqb0w
yHu5YKcuQpTudtNEZfYRPB0gBWolQzmzsNQlIbfVRLwi2Ou5ZUpdmLnAmq2OdKoK
BMooiyZrk1ggLgzU+7lgexQlCVxXPTaxkZbII4fvig0iiWhDSUE5x+1qFj5urVsr
VtiRxe0kHIlYtvZmVNnZ4coJJiDFhv4xA2vHlrDd3YS+nDkZd8isUxGZ688lxOAP
VG5fxJPZupmqvCM23JOFmIvjHKsQz6xWzZt/T9+PdV15arSai0uzUHnrAONw27Uw
nCaX3XanjvdecNICGCx0nHTXlJgWzOGmWF4QHYdvTSsSwfaS1KKUb1lZ4kw69ErM
sEH5hOueqcujYwv66zoPODQkMRw8yg7tnNKqWMSaWz9IXfzRWCZQJlUsVu3aIUGv
A711aomvJVGMJyxDtjoROhYt3YS6FZGvuYMDjPlvh37QOfKu6TxKR/323TtL38IU
ce9xt+W7aqtwfVXKxYGj3ZLissQNe/Uyv4eVKrITL0EKjTbwBnTpZ7vetiKg36iH
L0RSjX21kf5Ww1B423DlC+ad0OACsLHoM0RgST3xz2VGWv/NeoiNx0bODA5mgoyp
/rMj1QTSdCLQJoaJ6VccRQqibxagL6IvlRqiElVaZ062wJ/nfs5NPC1k8KCDTGpR
Pr4v/CDdoGdca/vf7jI7+z2+YJn+Pp3IyYgYnuUd9ySJQytnTRVT2IrUsqkVBTut
lKenq4EZNFlGxWxZ93mIcogtbnMM2YGsaPpWCfCpZDqgM5fX71bNp3ISq2k4EK3G
4tQocfjLtM725EEdKqtBO9d9yS7YHEIRPg+mjW0NWsNUjA7BB0KyFs8PwkxKQcAt
Adti93g009I7xp5N96h+fBoKj67jSbkzc4HBEPNIN1tyk/ekcRHoxj2zJfAXWGvB
nIE4NX+Rgmlc9tr8V+OgaFJKRo0opTV3elwsaqFGm2U9wDGM1iCmpMXds0eRK0z1
u3h2EwIsCZ031HzJjSxDwM0qG5JvUZgC6z3EIra9FDxvJiHdD8DzrkMHxwh8m02j
VZl5VxMruTPMdhLW+w9pr3rqhe8+9vQUKeGcUX6cNVYkEoLlv6cmTCfhHr7L0sX3
8GNVW7ubEKTJWu6zpwIb2gXk9fjAUb6ryFbYKfBkvI7gwOdpzGuntunzCG2wRVUL
sw4YFxAS4WKp2hr69UX9cH9VU6xH7npKRInti27vs+mU1IejkI/0AQXse7KoZUfe
BcPqu6jLPZqzIH+RPUJLpJAIx6LRC3eXMryeetN1DDo0AQjBwdR1aHTgZe5VfMCm
SaZ+6U/vkZyry/V3dMGQEpSpTuRzVqdUfQtR6g3TPiOTnTp8bfbaXag0zeGw/S7q
xU8KL1X9T/3PnSgrmyQJFfG3CdEPGiVcv4PIwxF2PeZohp4wRY/kakl9Ke+JEfzx
CeoktkTzxLDCrVb+ZQPT8OTmr/Q9JzjfvFwCcjKDmpJK/+EFgOHkdwWtFr48DUDD
fYI8Sh32oUsqs+sZX6sTv7CvT+YOQfz4EnnRAyLmHn/HKsU6r6Wx36XIbUsONzfK
Mymz3orIL9r5mt8ACvEVPuUG7S21t+SKxDycR1wniEMoDsYvI/fTCVitrBxV5BLa
4wm4B96ygEkT6GmEIgTkpBvptAkAzgsfKmIkSbqFF4vjIkx/C/HJ8UBJNXyVSEfy
IH4jLfoDU1KbkGb4ZoeybJYOhePnEGEb5we5shZ6gXV+2TD8s8ZcIfOEZ7CPcQ3B
GbP/TTSNJp9eek5ltdJLGFFLbsElOOfONEDu8dC/+i23+MGGBis5oE/7AsC/WHs4
6jfBufa8p3J0cOmJUuH0qbKUkrWa+1sGT0Avz0qTSXz7bclm0kjeCNbGWF6TBp3O
FbLl2KM9RAXYIfL+7WOmETdUdVyv+h9sBKRaw40WnCLHhP5sycZHp3yGlevQO/Ao
pBuPnH+8PtNFc+qB1brUUzu7qj4C+qMbhg4SDSWFSqIkZcWhiGmlj31G8YEcM9mY
diPIT9rhji9Ojj3Y6pZusGmBFI97plT7Q0p7HjL9Uxz44a9hM/sNQCfe7G/RTYMF
lgKQo/uDzcaNUJh07hPtX9YUrGzBJsd2yY/5MajFBz16kMOJVKBajaCzVbYy3ms1
F9+u+rwEigLfAayZZznHRbavbhzawKKcOoWOmZa3kXPe0wESsL6rg6MHkd1kwCf7
qG6GukWs8KctEw0gg6FBno7EEyYQgEDke5lH9aACUzUWkAl7ggNnB9daB5N+dNlq
E3wQNmVSk6vprgZySFUSz4YD8V1+6MAJFptSYiSe+RgzmJDdKlqq6tysbEoBvJl9
NxKhFjewAD3CkiFLMgpwvBsK4bgET9P79BxTKI79tYErx+5/ukEffvHdAEw00dfW
0qvIUndKuRYyVQxFWlzVhOo2ruv6XKsqQtRSOK0Nb4ePuT90+p/9WETyXyDXm7bH
6Oy/nCV/PcJQdxQCLt29LK6ADOrp0S0xIaYamkOgvcmALV7qQlIWAbf5iE8ZgcJ1
rUMWSADNbnCbDyhE1cSf7s26JZJzSmmrcVqCulbCt3pQstmoqWyptA1cUl3Mcs6b
Y4y0Yj3takhvzE3fFhKc5m5AaQa1xprlDClEqm4vq2OPpK8qD5WxKyS1r8fT/m51
DrDAvq8R4Hz0Z417AGn8tpFGJDahD7keUkEbPFOrB0dnSDMOMPmJUcXqME8hI5kb
st5VpjTPlB+W6a2tcbEu1AiyXPvWZXc4sSlCGO3KL3uD34keYC2PTyptuavqXN9m
0bgA1XAUfiAkx9EXrE1u9jvlbaCXDCG1MDDjGEqBEB7fE1+aUVSb2nvVRoWHf4li
htmIHs3cBLxdlPC4I6r9uyU7vk9Gb/fXWG1KE9UMCFAhuCJYqZFYH2vJG8l8+3Ic
AcZL+SnKoIQeEHFnLHc06q3LfE5eBwiQ289ICYap+O5LQvO2Ww7C7OJ4K3UF6t79
z359Q3/fyrdqkPU55i4mPiSM5Sm/830iafiY3Nj8CA6BJI/X2sTBTR/V6P351570
fVsuBFECj8cKzxZ5vcDLyxwYzlYVFJm1BHHkOfin1m7ELG+FvtPiK19ma+svGHak
qt3IesmSjSxfKpkoFIKDNfVVe3p5KixzvPp8473zULjwGwErodooPGIfSO1lFIN0
RJXAdtCAZTOn2Pl3y2aVPsYYZ9CVzNCtu5qHVYdgjgwwS/6wMry1OjO8525TnAOD
IIXHxak4b6duoEEhsCc2kWIaFdxEb97q/Sg4UwYZUUdiudmwe8vhgFJt0Mqinf4Q
1bIL4DJGW67JP6uiMQ/+aT1n2oEYOP1xWjbqpDka2c32oNYwR/ib76/gnP6SYdGl
JWJiPTNPa9P4mcX1m9CpyH2GRxLLujXc8d4BGpL/GYEAt2Z9vVeB/yhq0Lm9vYaZ
Jh22oom9snJjbPxJUiMlpaPPLgmhtHSC05YKGJ7zLcSZ5p3NVRcEqz4KSSv6e8J9
D0wcdf5C8jHZfCNg4/X4tHf0A+FsBokiB5JVi4+CrnFB+wVtee2UGrVgBllZvuFg
J37sdoOq+ubim2VIDlUmU6C09DpLLUuz8tPFDzgvKTMeFaizBVQQ0i/hmMCjceGf
N1LnZQ7jjgQ1CZkkDGN67FivAaBujoPyk73ZZ19Bc5fJcleRLbBnSSeocbkO7gK5
MmraNDjsEo7aBlsgzvPd97RcoDsxqoe1ZYmkWK+Z5PFcRKtZeX5aU+oNxyu7G0U8
fR73aaumDvI2lFVMOKdsvl5BDFLEwa17EFUT4aNwfgF0byyuL2KNO7znDAHAaoUC
+D0zeKyepfvsra36jjg39lqQWTxP5Gbtzv6Z1qjKWNfaWOweOHxfMABrOvLxIBQX
HYuzLtU0oJcpPD6IMcgKKICFEkgKNoQSW40TKrAbqfpJ0sD7kVha7b9okC3mHle8
Okbk+6C1oSFb6tCy2ipSOZ5qK3cE9GQGS3iLq488Tz/6B9jQpQ8TQRr626AhHjeE
5r8sxxlYVrWkAazGboUFi/tqUAIAI15mRQl/vsxBU7yRgo6OJ8sPDBkde+OQ5bIw
HmOH9Yu5cFAOo4sOoCta9PZY9QOeO4j5zLvxircAbZRKUvQKm9cDu/mlhoI1ahOe
PQvAonz4b40YDAWyijNMP0g36S5ZlcFGaE3jlMZidknNjwF1xKaVWdh+L3zSEW32
G8kGtbGEzPDRiQBZJSMHNSTKV2fa6R3umH6eysOMhcRFxr6dr64kdGhRSfngEY5f
9h2JGzFTp2FopiCep03yc8ZS+xcZLoNMPDWhsPJvM7nUXegR++tFHssXFse7XqE6
YHbY/MpDFwlTprkx5PrKSRquwFXoLlVnpbCTG5dsNpdH+ps+585TG6tcYKeVGQx1
PDeiluLBpUGbD0KcFcn8KgZImm6dMyuyRiRK4Xlps3FGJTf26Fa9jq0+TGXq+EMV
oJsL7UrjZOxXiSAadyKwnn5BW+9KmYtw23A25FvAsibI75JEmeXpdFIuZALcu5Wq
ZfxN/tw7qHo07ltxzNw4HQ+RS5KINQUFdcWQo/6v40aIcVT/jN7SApSJfWnFoTL3
JPTfJWLiQgd0Dk/vNEsDgiKPKRQFAnFFOILM/IclOmCRB3oqSSPauFaC1UckEGm1
cpJxWccLzAV7JrWv4HwJIow8ay9gWwUyEHGzW50+qOoTC+9juPw/qfk+ueF30xzf
nVbkaNCJCOoDKBVs9b3lkxahKkxvnCtSVVMGIWD+d9ZW+IVHZyEsOZA6Nga4oPcD
OlfZkJ9BIXXLM7HY4LWgoEw+Dlsi4ATJKGxlAoFeb/RF2CsCOBjffR/HDCLOWSyf
23Gxv8hnMTRZRT2Fhge1+FL6xTKP6pHypWqdazS9XBDRlNZ2+5nQTO5qT+YI4qw3
wFmUfQ0wwTwZoRCDbHOD1HFoVLQX4cvNwO7/b5JyIvab4G/4lq1UCTSXLgHNO83p
Z1SSrspu7DhsD26Wx/sgIQnz1WqhnCub0OcSIo9+cHZg0TIWLsE5Uw6SFDCVKiHm
BxAEdtEipZMPR0XpWUtwXgjzKAL3/bgXi297CkH2K64NIsAy7hwdf2y4HKjnNm/b
BHPX8jvMm2RkoogmaN5Ci4XJEc/glfbCin41EGIdXn999lnA1wH29gjezYUsPB0L
KtUA84lWPGfVS1QZBOjiBeEUa6HrReNhLCDaTqHAlEQlqaQ0M41PZReRNgukPfg+
3DhNBtXfQWaJlNXvvEkBE+gnPHbwpAyhH0pbG8kul767mvkWhwWTBgYFK0sADHFN
WiugCEXt6GL/Qvby3qEXQL1LCtw1pfdr8dEt0hr326fqLOFUO0VmhD8Idp5TqDKq
uNrg6cLeV49DD5LE2bVFgtZ1WIu40JhQpnc3l8wEDzgpvI2X7ybWgYJ8jAHSgrc7
VYA5mTi+bhAOrYlQrHG9YOU04S6q6TLC6EHIc+X8/sRE0VYBSPb+vJzZ3mf12Rsv
hdCUG7GzAsaGasTgp2MDKcIvd444SdbCOySpJcrQMyAklEo/mfWNW4lFbViT5qbG
u0hUX26VKx6ePE526TFkivaAA3BOpbLWYlO5dVPliLLUPVsk/e1iBuEl5qWVWMSL
kr655P3lrae0Rc4FZiRBjiSxOrrgL+7HX+g4qCr/xtwVQ1iAyaBHwI+1K2ur+OF7
IG/wzVKlhs+lWKQkIeW5J2ffCDNi63YFIvDWNy+56ex+B9JAbpcie5+2FYB8WPhP
Di5iAC8yS373O2et5e8HU9T+kX8IKDQIzI/E8I3c6uZH4HPSkcdNc4SUFgbARPkU
+IkBuSX5YZEsAEHzYAsgr+pE5ua0zacCMpBCKIMKZVTXHA8HZJMTTDOlOtdoUOfI
4TyDnD7plCjoEpwYAORf78wAlloYJpdRvVmYtGurj639hph9i1P5SIVhcTSNSm47
R2xO1V0xHF0+SgKJCKyVToyD49OAAo/rNp0CnDftEN0i5/YpJWRdyV6tFgbT23dE
Fg/i61HB3aqex4TxOT4VjyOkjYmsVIj2uP6HA0gOVAoWUCf2iFdOYMBpHb9NVVrl
vf9KjXKYwQIYm75tEg6SyaRf6VWpL7fBgoQaxebt37PZPcgp9OdC7kaL5nUhjd06
xDmzZz7TdSCoW6uB9kWN6GNRIyxLSO4m6TgBLuyzmqZgwi9lUGvrCq2xkf53QiXJ
jf6vjHQLLXhgM0k3X03++oCQ9EkknANLr8LYyqk6lMpjncjdi7rkaynXAbCuOKF1
yliT/kbYko+BT+iOotIDqMX0ZSZRAsItlGNPoCqcshg4djnRZ6o0jOD0cd08uSME
FhMovebfOOLFlZ/KBkxcIBnO2CfF/m5BZB3jTSote3B9iTAjp0yMM5LnGnHWpsC4
n1IhrGXpxPDKqqlF+a8mXCo6qIOg+B0kuGj4QEZ8dY4lTi8HFW/TRugJaRCBYqUL
BRzpWUOTIN4tABQHiDFOGfuGIvs1ULiq7VE4trI5UDxJyrnc+VxXo0sU0feqlt0+
vNxjUeyklHMzILmbTEs98kWrPW5yWUd8Teefwh6nnPFX9P4qpYizMh/WbEgHpXgr
DqSSqP2hfF9RGXBh/cesATYqBx7BLtCZ8ZfMkHgc3n+V+uESQXpcRFNavI90i1Si
L/TKxYE87rjfHUP2Zj/O6q7w0Cc6bMF/9PePNxkMnm0BPftA4eUE4k1YGZRW+KfA
O7lFhLww+dRlDmFuxOObJPuMsmDqesj4AklRNZJIjNogaxGSUy7jMzRlds8W2LsN
nQs4dSoiXHYs8piolFdW7FXAw2UXskYL1yK8VOsxxBC5fm1+yUxfIM0fUS1pR6TG
KCV7/uX6rRozwA24jxYU8wm2OWd01lvBQHysK4HQOKSYkIM80iNoZ7YS9B1ne+gP
bY6DvG0aJigYexA0FPToWLcUEKCda6wcNz+J55ioVnpr6AcLgcCwgvHh0Sbzncvu
eZFzYmB3Hj0q7zdS+/AL43RIjOLkLsEjO7alQcfM97gHEIOiOzXfuudPMZTQxosu
YU5+TwGgvAMJxZk6Rx5tap3M6Y7GE9WV0l/QRwqgc5QOgyrKIZaqFVO9q9ygOWpX
zCeHHgnBA0R5nDBog6AMx1eEO3px87EjKlHV8lAiiK7sw01DCYpFOe67Mrqi6bji
qwGlmVEPQOv10nUH7+GQcdGoRDbJL+fiO03uY0I1MJLv0pVPnGzj+0L2lCHC8+ed
wfk+qKX+qeDqVlfQe6jmrfALvzVkkFEXAnWk1DJXQK4je4PypZV1ZktpB+3thJQ6
aeCJ0pZw9PU2oSBRHqUdDtHteVfKJVSrRqKd19RSEpt7D00JxYOCQR1cW3thxZQ0
yPZxOd1/aN7KTBfdMMiIf1m/sIpI5wq/KP0KPuT0VLLyJz6Qogo0oCxC6weqwK7Z
IhV2LmEqivtzcI7mfi9EynYDn5hY/NEXn5Jxl5DeYsfZtV8kAq57SZlrcFFlRMt6
q0/jyRyuIliQl/lciJCy/IzEr6L9VJmorIVnDl5/4rLBpuM8ZLyDmyROqm+J5H6O
5UpReWK1oWVZjnip5WQLQmCxbPJ+crd5XKN83aH8BMmeFdP8PJPMxdggnuBe6hen
ivARC4mhmYmqa2X/tLFhfvatMTF+TaTZGztsZ6TnzvJY2Y2k100UfpwZBIG28jdc
URXGjSdo5NYMb+lacWz+jK/onGkA4wNqk/rso0mLdYGWv51CZAgFFW0+aFeu+T61
jtDbLi9J03PgyKGV6Nm1XqpRQuG3CARGWMHC6tDhdhJl7r7Oncz9jqhuUn2mYJ0T
p0dY605pS1buAkC1lB1vX/R0f0aReECKWtnwt3lAEt9QN8yl9DZ4IeHHYU2sHmZs
7jsAShKWXGX8kwIow+J8OH156kBLb7dGqAE9uRd9P+ib8cHvUvJazVEFo1qv/BDd
2ufqvjblN8O//4+PPGC41/OwuFm4mkEFI3txiiudiyHuIZbv+OtwXyZRQ7/ZxqKS
jhWle9Jxbnx4NzSRak0+BeXDrhHNdNg21NEIPjCVCre5wbvRYIXrBK1LpeMyZJvT
DFaotD5RAKF+sD1WBZyfaYB50bvBH0S/lNt2JkQh+SERlC3FxpReqoVlfBrp+g2o
1zPmPUjHCFax1IbpnVPbtVKZ876aM7cIlo2DKiic4pOpq+P/+3d5rDejBAzwQxoP
ZmJAS2607ixSHHflsTLKhwe8BHhvU62W7uTVb0mXLH1NceZRzkXznOcjp3NBr8dd
lVrggsHK2veDXEX8rry8U2wdjdpezT1gK49FgYF+pnFpDJbOjJ7ey4KDZdiiuZaC
oZWPzaOgEoVTFmV50FlXsMaYOewJv4Ocq7clKBWWfKk0e/5D6jXulu83vXRiMrh/
iBdF9K1CQQt6g8e5I5FMcl9mIsyWBieFAxsecWQGoKYYva1ZDGFYZmZ61Py8hz0b
Gv4NXDO70ZarpUikqdH8Ykl64xf+6qhfZSnu/fswe/FMHLTXWsrSRXQinoSwVkDA
1d/wEN3CLhVjdzFkvxZiJnLEjYnPob26lRAwD5/8X+B8FrIbJEfTI51q0yUET6o1
bpCEm5iikhm3ph9MFMLzDYJiA8G7WhanBfCZNov27JDrYVuipF0P1zLhbuEB+mi3
W2nSpqixLBvN1E6uXdoGI8wl+gNXqI5zPg7UE5WabnwufC/VqhsF7rgTEM6RMXt2
dnLxWoOc2iIDdjv9sG1EDu5EcV76AXnp81X4lmLCJhxX71ugW8mLJdV6ueHbDjAC
UXOqG62NB7Qh1nsbeX6AFTKGvdIYAW0c1IMeXIE5C60j45Qlne0pyiEYINnGVgRj
87w5tkH4ZHnQ8OV0xqXBdJuoenANW3NYOthpESnuYY5TojUFVz5NLbNleIrrQSMD
ThADGVcKwLWpz/efsn0TPjNEyl7RjKwulEQLsmFLcrYEyUZaaiz2lVv/wUiqh/RE
2CnNtDSW6/26ImNxpxEbD2Z4ui03V5M1Vizb3xuWDr65ZyAwaNugBoue2Ct8eQDw
in3zbalz5M6E10dWYR9BTSu5uq4Q+s8MWSuvdvQTmcqPIwVZxoWdoQhOlevXEU+9
b9OVZfrdEkYSBfyIuK5z7YgjXjpTWT/uiUv+BVJkemyFAv/gm10+YD8xh/u3f298
SoNG858DgAk4rgFpJVt7fHslnuVIAjPVyN3z7EWQHZTlaspZlG4SbPRgv3DnXKTs
64cJFIHzlcFilGdhBSmPvNkkrXM0n0XKiS886X292PFLvg78/xI+/HVRYrBo3oIU
fBwEH77HJV0PodxzdThTK6xRnuH8CaLeNsNblAcPRLTTrFAnVWl6FX3HLY0uGCFb
yQhKLmuPex8dWcwrf4ZUPTOSvnLsdg+wv3W64/6jxxv7PCW5oDekiJztGCS67mTQ
83tuAFIUiYFzMpKh4QXW9fVrYrvWwyUBZ5Ij/JWfKxvsc02ux1RFrRHHBny8XiNY
cSudwS8kCoOvu7DS2M01hm2+9xvJaRqxYAagqQJKCyJnPoPOChsQqznZmk//UAcj
JRCd8lGKuIfUPLFKZoCOd6LfrAbluUqNAoHydGoAoBRphLo58U4GuvdPPXXKvxEw
+JCAQennQ7zEto+cWNN9EvccrNe3a3RdvToImbCxZi68RmCwfqlwrC6sXRaCRr53
Qi7yOuVsL0Y0i3y//vaAx3TpeWTPHfydjydg0ugniacaQ+oyOLUWjYD7wvEM7pxT
BWpPKJ5vDpbYhVT/RJjjEzlV/tfA6e6Z53Mr8GODdu9YeDqJfUXUBVmfhfepj1XK
EWgp0n1UlTF/FtKoQm6twVNeRbHbSI120QN4pSOrsmdrik7aM+26eyfyLBJBnQym
mR54yrQ4yib4jI1MYk5XgUg9uxWbcQGcSPrUUheP2A9eSLoWxsU8WxTjbso2du6O
FKUuYZKP6zwEt2vAifOFJ64DYtV7zeZZS6O7uUTkvrqcewtdoCfhklroj863dc29
wrdlLdEAZf3p24hQ5C2CadN84mKpXmBvFqnejoj0sOD0LB1IJ2K3g0+1sNjSrDNl
7RC+A3Kue0rlbqQvl2NB0cT3IsuJ1K8iZjKyBrmcylyQtIBwp1ttQ7UBzN3y6TeF
juKE9SDPj4BUV2RGHCuMJ8ItjyHTNLc7YoV7mY4mfP8H3THGFWlIO1hqML0gNYcG
EUxknGxtSXQ5VLL6LibOuwcioE3kMFALu0/cKNkS6ZQYpl+/+FauOkiWsu7cNBX9
l1YNIhDofakD8p5VWyTrotuFi5ArDIvI1T5H1QmhjmvHf6kJhZzL1bfsXtizWjml
HM9GXfgZeS+LBebMgIwEGTcpsi9Vvms1jbM1oGObwi5R82/tTbV8NUsyvfevRuY/
cdSDa5V3YpHjV65TJRtcYpa+Ia1DDaKUMzftdd9Zmx5SOu8BAdFohcT7pYn38iZB
u65u42ipw9ttNZRHpZdbL5HDXEZlQ//hh5XK72U7AgGNCkY5YNeG0xBpjCWz9ZOL
k5jV1fhJYFs/BMHeqXyVfDKp2fjANHfj2nkBojyCkhqcJQM2ETgUEK2DtcMS422m
/xlXmGvbaq/88AoIDETJfgtvOm4XCLEogvquEeXC4lmsa9mU0NFk1cxYenosm0x7
j1VdF3wqAngpn7L6YZofeXqLnw6Mz+evZaLHm0taCDaB0zqjjfqj2MBUMl5DiQuQ
9Yxf7ouz5pgluqsqWNsdG8BMU56xV43l44YmnHYkjGDAVdgTxkfAbtzmghfxGymH
kPLl8Wh3If4AbeyeHRIkAFLKA4mPqr9yoGqDQxFsiHUcvS3yaHeYBg5hjr1SPbWv
jDlS4FCPGHV3WHwwpy22ZBsWBRx7IMDtfeWDiczPdHrBnOn39JBrizj1f7MAmiv3
QtH75K2NZj8dX55nRAGPw24KmGar/Omj4LthZg9IfaT9vftM7SHlUao+W8E+UFJP
2Y9d4rwqSadX9cTT/e/7HjlmggETOdXCmrgAspNBNZjAmLuQJWkDV6LR5cP/ob16
79tK+rm920GedJJSPXtJwpsR+LwylLPqs4En0gAxVR5sW/V+RJRm6pIpiwEt5g5i
DN+fw0VMt/9OImuLGeqp8Xa7x0qUTvZOkG0jg9/P3Ftwn/UARUHTWcjS5SleUqth
X/HhMXuqoocpr/kWHQUl4s4FrymMKE6eXql1FFQbz4eBMjqBa3tlsVy+AuaK0B/M
mbEYAUQaaE8RlWy3q0dgfjEmDHPBhed6t246Vte85Saqs6/K4kQWB/ANExd9s2m0
L4Pcip1PGWn/iVp6GkWh2J9ZAorG2orK3qGYcQK9GAWtlxfhirM0Y4LISI0gXyv8
dWpNwC5WwZ+a2t6bebfy83d9XAFYd57LoS2JqpGtrpkJ1XUyfSt1AEyJrHYHGo1u
XTl0zIGIR2L7M+wIVWs23MUUuz6RFzqrdcaVs8aBjVUoaSeonhGwPHHInRa1uucq
++SoCB2Ka9OC5njlIf3FzwzS4JSSAYhdngwU70kPXfkk+GSJNC01EanD6eiOoSOV
hj3oH8Hesy2klX3KK0H94DppwAMawzGr+iNykq5+BnDvm2XulZ6Lih3HSY4NZ7m4
3rRG13Ru8g2WA51ZPhvKecTnMCXgHWMKqrUFLUh1hEHTq0IhJlhFHxSAXJToBHA6
BWtAd/SL7Ijqet+BT71JrmE/SgKTNXV7p/a+9C9anFKuhl87uSCVtga4nzzCpcwQ
WPM1CyOHUpq2bNe66g9yhReu9juhtYD2SjYtinC5hbGntWhqpAqDn8hXblLC+uv4
E9I+YNWHozmKqgvRLqZOlBq+tleiGG0KkxMG42fVC++AcEZJq9nX6yv/DrZTQJn3
n5plD4oCzE2m3Ir3SbtHvBmVXJIkjXiyJIRpGvgTKS6hLiZNuFKkNxf/ClZVmIPd
Wy0SF8PW6pso5A8mTfOi4BH8xrk7r9bXnm1X8i2qY+g05yJs3XnXWjXVLqOsIJU5
X2hZezFPEuhMkmHzVf43eIflJp0Lrj9CKQq13QlsbgFovS5nnoDLxDWVDuX+tpON
5QowGillpCxeLPmoNf5uMrq10QGujXC5D40xPeGamSkkg0hYaAp1iiZKlvkp/KSS
zD9nEEk+k296J5/3aMAZu+MElgSv/Hzh4P+NWvbPNYunnnBFbxYQfXsX01uqyAvs
y5uMAC0uh9Oi7CiwGBHUTT8+95vbCPvinjjFutSQ27vRjvgeztdmwL3UvLpSPGAZ
lEXClHzwlkd24G09B002N0Nrm+IzNc/9Zri0Vpa6x9HFbGECm9mng3ns73xRPw1y
KrgxBTg+B55mcVvwC00FUqmzy4lwHxmLX4EoGbeBxoMENIFFe7hRYWlaNjGQTisz
I+mAjO/RX0caU/eFd3RxQvw/emFgIYVfGPOrC1WlqofpZ1ZOED9nror4vfxkQaJC
dAaydnoU+lfen9QvHBG36lvt5Rt3xnsnYwRKs5CoHANamQrYXrLiU/LzWyQig858
Q9TAFiOgXuSGt4Hb2PCKAp8zPBYzpWQx/MnNs8n97Rb/MxB/+tfcu9OPxnQ/qpJa
QLgjybo6d4yenzmvMRXsDQXZEUHkzuimpErHxD52V+vBT7bDdFeqqT6kis9nlXY/
/1g0HYsb5mhUmI29mRF04YvyJrvVxy9Wy2pomiolSFNv9a7n4vKNhcEpAMOE45Su
KESAI3IYD3zLbAkK+lqsAk1dINFaYKu7cTHJvczi5Fwt8kc2uJZPO3mDRGCueTAZ
S6iBaBZtRGrEcq4CrKgZXMVt3SHfKjBnCP1NvfPrU71hVl4P7RUsndlftp3KG7X4
ibiCSL+FzhVwyqBwsuHkYGxrYJJdzuCNy+7vVprW67xGKLTWMV7eh/sPfAHSAfSN
/9jOi0q3RFqb7jIpgZu5vUGnP+q3b23nY3CSq/ZaIdEuSbIjxaq6gfj88ShnEQRH
sEi5H3SB5JJQrKKfaphn/c0q5F3H4cGRMH4mD5Xwt+IonzW9uvffp52c83yJyEag
hKicY850DoD1R7XXAzNa/2akq0fzH833E2EZt3pkFbeokpLwy8u4yleCD/gkwEUe
sAzTZEGul6TIBMwM2xNaXyH6YOIl3TYNAGZSNYZs9PbLq0kCFi06Vv7t2Z3LpbDl
KVODRgyJlJJiBJDvs46ToMWJF1Ir4naMoCHRzuXkEJEvyVDfR07ZxRkqMeN3C52U
q6uvDko2//H13q206pxEMazb5ReS3uTgBpT0g53TullZneZ2NkJqgON13lRFN8CJ
FkwFubPOKv4MZN7utX+Z4MbRg3iBvJpioiZBfqjmDedmOiU3XM6h5WZ6LRz7DAIp
29wFAC+Y+Kw7Eb3hXmVX8m04thAnbIJyHyMfUZhYWO882qRdKmE1eMyLPnsF72WD
XdZMilRv/SQspHIF+bPbjr6lpJV9kdQA+XZtaHmIGRVu7QHk6XjNZWVjjfToDdbb
s0Oas83u89oi0p8YtfZ7WwNyaHsEVdQWq5n7cdonRAZ+AbGD82q8UPbGPf4HUjm6
ythQ8q10bb4QLAALMjbv64boCmcehiK/eD76MA6RAMllTOhXigxtAFXF4t9JQ4ju
N6EOKP/a3/M560wzrofPE1KcVYrTrfve6C1TZ3Uvhx/ZjdTIiJyP18SXibWio3Ar
HddYrgrRktZmjCXnG15Dj3dIMkhoNtiZjCqjGZxj8n0wJPTUsc07E3mNqiV+Fz4D
wY1pItijmdWixKWIl2iTIKf7wOpqrILd+VhKiHeTD2pFEGLOFVnKO634xpR6EUhD
h+RA8Tgm2+4A2AuZH+bUcIZwHPBKx0AFc3Edpp+aj9mvSNdHs3C7w6Ovm3UgTdgk
d80xH4NTaABfp8o/Qw76u0rpLCMZk/I8Ttrvcr7Qa7V4i0O6Ly15wNJL6t+fVvGz
LoIFmro5MHwX/nPM9OdNjDCQSF08paz4MqgxKj4QPIThPXBdwyyMJ9RiB+Z9KjEa
LRZpx9ImroESjQSlWTgOpw7M8DXjCtDKrFOLNicZthmz3p/vSOr9EJT/lsxkKMxb
IRvO30aHEPU4INmkuyOJMENJwJ5lUyMuwdvBv4BFsf9YpbMkyl0OgiQVVfW8cyox
WjdYP5al6YCtDYTBGUt7CTZbBM0FYfU095b8JOG4vsCeFXvIgZNnglrRPQeJOxAY
s4Quly5xUc7z6jQrDU7awhLMu65F7MAeR+dStKElcYM6dnENbJ8AOBKDEVOXJdgs
AzXCh4rhCue8mqO9waNKCGr6/rZVbPcZK40B/OEePzfild0YmRF1eA0xUM+wMt1V
mcj1UO3mClkSZOufrPRoihWHvZG/AHOENPdkuMdbkkl5Rm6tH8C5yzTlJlQGSnJq
r1/YiiXGsfvOZdKF3OJPsjjwJupwKuYWHVa5hX8TpQjcCOX7A865s55G0iYG+oFM
nklZw9lOsTyGKv+TZmEOQ/EI51o0FRsDndTAmy0umjxqHbfiB/ysHb5cDRF2WHW5
CrkSdLNv8o/Xtr1bGCl5GJYYD/Alr/6H3NZj4ght/GI06kFMQ1nDpZMeESuljnB/
YtxYxASOGxMK3xamS+VAUiqr55VTnZ2OC/1xKxzns3Ull3MFyceUXQVID2NDogV5
3rHmxy98ZWS6rhTi1T9/2llIKnrffMDkAn0qQeQ5mQH1u77AMdeHrjE02Ln5yEtC
A0jFjyko19vnGDK4swGGXbdrLq+8K1EWu3Nf1MUecYLeQGv2RgL6y2Z2ogRn89uB
oaZDvttATWdyJtag/CT/C5NNysO4yWvd5fNM01Zb9Rv4wEwH33BneM9Be4NCzrR7
R+x3/gQ/JVr58847j7UjG0EQaamHlJ6OyChOhj2Toq70dXVayzzmoPi1X6hx+aD2
2m7p5/Cal1hK7V1uymjZBoFp7Jv0ALF+hpJOf/62sja6HGWvRQ6t1vlHbYaOaqz/
gpbFFCUjbsbFAsr5VZTz6FdeZN6+IiexEhM8+Q0PXLRLlqGK/EkI5wWS0EsfufP8
VZtpYZoWg1IMuvvFVaSCf7cNRH2hhpK/uZZzNstHhXYnJmOw4jCWATEBPR/As4Kc
NzzJnMf3fuJZBzzljTYqiwKUSTjPQQI60uCrvPMqTDwYCnyWpFNIPOp4mSbeVm01
S+KTSN2bvB5Rz8OTRRAh2k1vACIWoo4KOeh57///V4ItCMYSTAkCk461z6dze3/c
2eSP9kYeAQYPpFHbH6fi8BMCO5u8l0djD6sC8R3di60CWT9IEIScK9sLERp+gq48
07maPdDghr72++6epb2CAAKaic+iZghzJC4fQcfVbFRHY0Q197qXiieIp4K1WV1V
cyYeO5Izb7qydXMBl+VoY+BiB7LL58rzxkTplIeSQEaN9uQRF70ztLGc31k4q6cC
1VJOm9UxFvD+IkWH8CTnq+uo7FxHCYKN9x2qIEnOR5reUzquyXjDgwBuAEU1rVq6
tmEbNGbcYLLTD61gWWY5MfOEn4Kf/SvByep9mvevVUU8lsnHbcenmpG0FuyMXgfZ
P9fad/Jjb5zud3abS1lbtjektHoKK1MRIgfEyZ+bqLEJlP4+UNZRQDRmp1ZooNpN
jr1/BQsdgwkl5M2NtyWXqiUlDvKRWJTQL/EBJHX9u0HkhGVM8PoYPRRqZJQJHgjJ
4RQ6jZro/bIJk9OcHnmI8YrrwgW9qwtEDfgCGyxXldR6KCc81x1o+5AFfrKtvWrv
DyBgpTUObZRO7SoSqfIY9SvPiSvoofrBC/4hfNP8T5vsVZQMEdzw/Onu3NxRtRiQ
1DiA6be58d+Ij5kNFluLUS3db9DomvdfUg/Hu3cqkS5EadFsXyZxLxMKqRFIxnG0
Pl4q50APpCSE1bHv5pyJrNuJ44IiqWsXP3MsUBKxmEArQugSkoIK7ZAV9H4Dc/lV
GhhAGxH8aVP3396uvNVxRRXTbpECGLBud37eHS/bhUabOhkp9927ElOPpfXzndQR
gCeF+MsTl+bSP7WjOoXK6XxQ3BLY9MATZPTj/7dCNtW88my0TT+eyeqUbmTB+JNp
161qsORAc+/nXh5XNHduGWFkYUM49yafwI7ztOCGi62/gxlGdu3v+uUB9LXoVl3o
ouHZ7ojUGLU6Dt9phY9Yfzff2R/0KfR/o3zTT47ElxM6d6YugkTTPnb6oJEYAfC6
hX93Y09ChkBHRUHEKTrxonowYRve1esoaTXKFbYuJd6xsJfiTVsmswnbGUWXgq87
md53WZHAvyCuzxvSBquPhv+Naa1k0K3CHSueklr6Eeug6LGjKRNA87nIVYYYIfEp
3NS/EoG30TP2bChbiuy0lSMtQCuwgnvI2zfl/ssAf3/UhO5mqOY9B4EFLmsW6cUh
gqjWiaMwMWAU4dCN7Dg5NhqYCHmcDfCXDQEFEHyfPeRHbujKcGtTD3hwoYwzioa3
9rDRtB+bnfs1hlpM+TnH1nNssoHjPm44RKp0bZS/7MCwEE6ifVmv14dH08dHFHj0
WeB2i+H01xKOYOhq8O36XA4hayTCP3BZJWIHGKp3yB7ae06DUpHV5qH5qwxaYkhN
qqgjSRLYgE9/0eydoCsNMbWNALKgQ5XLtfpOR2yGvTAwVNmBnyeCvlFYxwONEseX
ufvfwFw5216NPH5hnwIZSpxO75XYjIUd/Y623bfPhMM7fAsURA4Qg/Gy+xEvfOXi
yI+KOXo20qn/WxrnkeizTfhV8W6EPci/MzvRdUGtspFUs4J2/7u8h6uztHdxutN8
i5geEFKbVBYSjM71UT5g6bLQ1btPgnIowwGRDNlbwV1UFJZBx5T5PPoP+J0wRT3n
alWiOnyjJpPOFkvd4AhsgkajIpM5K2OINWzVDU4sxp02KXCv4Cc5rhkMRes2YGo7
7SvXzN9XcMPvuAFpTwFwjCCq4bUUY9kad0YcqrtCyqPUvQIMPTDGm1J2MeJhKbe2
LqhB2AzHteEBlSfGMYZxiIupB3cDk20AiqUOB3WjaSBX1jbe79TxwoxZb9ZXW/vt
+cVS7a6ry456YdYdCy5w2oe98U8JC3xRZsGDgkECf25OMIZpNwJo0Zzv0Mj5F8l4
dcb71Mwu76ikepKvxi6PdP4SQFFsiwxsnKvlpKyBCDFg/Pz6kXGza4WD5JARaKt0
WVwn+EY0JCWFxzqjRJT41PqtQtjj9YirO4quci68dkQMpZBTweEjWIWcHuQC3a48
BHIEvzWDaHoyfMyUy0lGDM480zjYrWXKZTU0vTv0eRjAHiXpu3HKmx62skajHyPT
dB08Jzp+RQdeXO5KiOgU59DPCosgKp9czQvxwtDRw5z0ZJSU3cpLUM4aNcZ9Kd+z
HSfsNjgAQSOyDohk/Rk3A/+qgAjWitWHae2ASwxkF5Bo30BDLJrBVEOo7AvyMDhE
y54Rm4T0vbEiqCO9268ga0Gub+F6JrzuMsiwsuHmZ5sUIlV/JGKscOvzJz8OJwsR
WN2CQ4kujD7l46YR9O59OdTdfS/ufYPf3cIyn2NfMndufLlHBVQ86pZb9sbU3ZNH
RXA8BLW4sTG//dvjxVLFsZE82Zj3jJBr4DirBHkt2yFDWKvl0kQrSTR5W/4yRDt7
7JcNqY0Vy1Xe5wEi6s8k1emohAgSuH6vbWAbm/VOG6pFBDv8Gn8djVOwj+WzQvgk
mk04eS5BlAH4zaS/mLvO/kvT6VTvp/pBi3Q66FHEBkRQ3sPTVU3qkoQ5AP2AQyL6
PaYVUnIcBB+z0xDy5oA0oKhr1sL9q7LXxTtvDegz0sMkc71ouNDsRrt7t8DVsvwb
/iPk+y5mevgDKQeXQLYp+1dKykby/qgD9uG234F55c5yv/ZjIt3XOq/DLrKcgffU
A723ogv5xPw0dJC27rwB73zqncFQvw17HAU9wqAfvUK7kfMMIGUdGWg71kEiB+G5
lHtIwVyEdXhI1hvVk4rsRrY5AhxTbF56Et7cau3pIb+U3GCYOrXOnDszUw42V+7Z
0fexTHg/rmBrxSuy9i2Wg4xQwdElcoE3vXOH0SghB0u9DVmJnIIME/Rz6FMFCsG2
lzqPrD/o6UXAwkoCU511DC+281LVuXiP3zJvvxwIjbtctyUKgcPrRJ4YxqGlpvf5
SNrbFKOPQQWRsGp7suSJkO7RXskeVg39SX8IXVKamfylTTBW9AmtBgm1O8l6D3/j
lKFq8KQBeAkv2r5tpFWn55tx6Omm4nxHDfmMuMrBBrzF7rsclP5ECAvyQl+EeSV8
xqijZC0WIWkyjItmhyTNL0PSkOhOU7ffGTBCQ94LgzEQN457NG+d4rc/JL/7DABS
OXgIUfmC5WZONbNtMVYwUK8pWhu3NiDzwHJQKkzvZb6gvUw5SNc7DwWQ1f/knGA3
MnQpTFOlR3tiN/yFmQz0L5faf+OszXcJWa4YsUJ7eiAE2qL1FgStFECKCWqnoU90
7usCv+9hAGpFC9J0mNAfxipkvNnrsR8cbRZCmxayudvHHHnrKM+UK7Lubfavy0u6
do3RXGBxtB3xRvtAlZcg1JabZOeFLm6a3xHciI4PFEM1vHkxuceA/XrUrGOTrdvH
qAALP8F2mbN49aMmdzzxQ3A5xKYzQQ9h3wi2vl93/5gf5n+kFBYQvUNJAU+QzYZZ
j5uEE+oOUeMDCyj3FBsYaNtDJd4Z+nDa8MhJCmYCijvW76/3Q0suVvN09ZaDjHkt
VOSMv6e3s2vkcR2y0VzM1D+4dKXV47jjkCNpmz29RvNE9vLpYnKcLQYaH310VAK/
jnDzmjF5jz6CVMd8gH+r3A5EoXnAopzmnePzSVPcRe1+bX7gc2X+eh9DZnD6uzLh
eu3Eh7FHob9TDUZF5+3sJdhMPiKNy3wu25zV319hoiAnoYN9eSpmwBa9MqKKgC/7
cJ26EItWeAzvZ9Za1xmOy0/Kq5ZnwQ15VXbO3kq4gwzWAQfy8p08bw9vQX3swLJG
BfjFH8J5pNQTqHBQ6Y7AeniwZS/D6cVzjg9tALC02xw9ClHGpJC52Hux0pO+mXqZ
wcPn8n/JUEmdNs89Cxv6BKct+AoY0D9+USS9zEOCQDAjHvrE3CEBCRWX0gWO3h7T
L4h1Pl9gkHSTBiFk1Ay9uEtWYrPr1R/aLxqK6zNoGyisATwLv7EjjYUatjBB0OfC
BAX0OEAW3AnSb4ZynyoOUF/ngCOhnXz4ohKCCH8Ez6hh8c+kE/GhJNjVxo9jKPqc
xjmj9Fap6QMeDHcMJAd+wnpKVTsErmAavLMtc4s/LTOUI7Rc+VqCF3R3bqvh/gX7
u+piQqn9lJeFNhGtO3QEWkTbg2sScPAZOQfo/PtBdCWoLxC07e4dJCTJx+WTVm0E
qYvr990isFtlNoQNR0ohLZ/zlC3FIiCaOWxao9mY6V0Vq0ygbGmtumJgon65THKL
PWVRnLMtIa2Bl4B1R3p8YPDwPtE5Vc150YyZnCMZ4J6ds6EP+uTxp0vXvEePp433
eF9YVBaa9HgeN6gICwWRLxrWeL0IV9Xth5IvTqjnnNl/h1OCBrVt+643YbEAXMzV
bDtcY6HUplNqRBdPu7wZ9UT3FG8fUhf9RC2mLHSzzYM72h4sUjHjC76FKRE9l4uT
rpeL2naBAnjqbFNybRO+NhhNgsP3B6vAqwnswUwNgwNxDKcy6t9O+hdd6X2kLeDe
+bDM+lss+DwKZmVaPAbTvuI8+lP9RpaF8E7/M3cN4paoufSDsHZSeaG8GvCQ0tXV
WwZwNpkzmzAdTfsjPUDfWH2DZXWaiRuO4t+DQPK6UzzCWgnZbqWqiZpeL/uNHm5z
hWzQXMlET7vwyGdS65HlIqaMzmvAhOtrq1d+eBS6/E3rYaSTQwKydj5MrNQK0Zxx
nIcnYK6nrbBYTHktmi+7BoeWs+HBrAi/K1I4FtbvCmSNcAcealhYZMJ6p72f35RO
SGiWV2/AoSf/+r9+1ncQq9LeHHpbNYt1mcOIxaVQob1AorNbsG43ZG99V8KT+qnK
LEr4y2o1xnyg/YitFm6it4onQGwsoomgZD+wQzwAZaqyCufYKMomd6pJdcx1u1rQ
A29sARGpLX73Wp3bXhOSHr1rBVusVBctPkNW7AMYjKqfuxnZoh85csbinZpQX5YT
QNs0divQYlKkf/jhcjtn3hOsIi9FsygzaLlHL32mTgD5Oia3ExV7BlfZ0Mu/+gNS
0XXcGTAmPUgwCKTqkrl+qWfOwEfCZ3M20e7lqVAM3a5faLfgpo8HGV90Al2Dqx02
u8ysEjJjMjCyu6DRagblcrQtdQF7LGcjPjOdZ0AVYj3fYdeufTha2nPOnZXz8Im2
HHRgqNwsus8qR4rH6x9QM6ylm9NL/R73pIcRSAgEzxAPfXFm889LkLq8fCQYL1i7
NNrfegKieNM3j75MZ4Fr4tisrOQZ7buKgeKQHzdzCqUVxvPZ3XnwYBDK1oKL0a7E
rEg+dAnuOgXUz4B/iZ8GsA9Rreyj+WgjisC73dJt/U52XY95WPW33J5AykGinmhX
yfB36yewzyaJ3ZWdf3iIUUxeKIt5TH+PVuq1qfIxoFaYJ5mgtZAPmJzwf2V+pYjj
5IDHbeUO9X+EeLouZnCdCuHsjqCyS6LP7DQFcx6ZcHmH8i8zQmBuE/mKXP7+b/90
C0Xb3sjE69FEagrxzwohy0ieYqMPe+PfhCRI6rWa723D1lhGjWmxq+Sn1xEUT7Pe
dNOxAShNsdSUQHZPDyDYeno9oYfl534CQtr6vDZ6+G6iR3KumGyTIfXPJmkI7Ns4
4pyH68iM3bkssLq8rmzKFkzHff6De/PqfxNjKSx0tynKmjofynoVnz/UII+xZVC3
p0a6P/MeGZP5++bo2lZgLqjjO2nDCBMgr/Y26R8iwPp+Ax42mu0lNmHPxVgpYm3+
yLba5qdGf97hSMXJAONDATiE7ShIODxexcbs7RAPUiSpQNFHlFV5EGi5IgdHomTn
YHnxFigL7vpNmFC3JSIcT/Ku58CHyYqHPswVC2rmDUh2Ry2duZm3CxzRRmlKJ/Ih
w6EnbT6UYxaGUx7aSIdrhFFSsQLua2HE4Pfes70JTQWbRX5LJZoKy3VZNOAcazun
Q8Mbq+MdMYVZe5ElX60CkvMje/iVn0y0S9L+ykQCHDzig5Urq4cJlCp3wvATLoCp
RnSfpz7O6MvIMxBeJj5UiRryWBZMf3WwfAWOyzPgloD1TfjBipzolyG29ZUOfLRp
SRcieB0CpRZEqefkVtc68YsZUGbS6I84uEFIBj2XvaYkLp2mBP6xvyILW0PKnVob
xgPB2q3ONRijdQqjDxhr44MR4ehpwWKT5ZTx05NXc9gj6j4CVTkS2naqoIDM+doI
IseP/Kocf7aTLYivPmymVbIdpNQXdwXjOGCQTLAaO1IhnTdIqB0p/TQF8hlp/CKb
qrpbDwDDX0Xy4W4w1UrHxIz90JP6VRNd4E1uvr59N4KP3hfWvz9aBXNzX+c5PVjL
biNV40z9JOuaq1f4CANCkCUWHOVhof3U3rMN7yHDMJ6SrKKQlzkfkQVHEO7E/B6s
baZT+GSaLKGrWMutuiPSA313FYqGoWwq9Pc4mw7QbbJiRxcMcTA1LB71XdGLysmN
n7/xCEynt4lhvziBm3QxfSmayV3+34niLC2FV8xN+ci5QQIxm71l/XX6Pq+jKOqx
dhJstyKHte9uO3WYn47tg4Sxb92eXYJtZ5QxsVgBgOt+Gb9aVK5G3rqdQuQaJw9A
8m/LQ56t02jAHLhHQ2GNjLb6EYTuMLIvt/wPkLJMiK8rdxDJNrV3Xe0cYvJhl/0z
r2SzY6G7BphV3l0NkQ1KMeHPBeb+2t3I5y5+kPIMRV3l9y2FYO6H7UhMNUEZOraB
gQFXEFncBgSlfcggJ7T1c3LyNaSMh7yJF+oqW/K8QDBYoZCtc2d2/bZcnYn2sde+
iSvcgsBBCsculWQsVWzdWlhscJTA5+w2L+WMIusRmipkN4CryKEACcPnGNrtYpxO
9zOpzIzd+9O17osjkxQcFK9vPmiF8QWyuiZs3a/qKweRClS/CrK3L0UFRZRECPJG
M7PPJSipsr6HMsSt6nxM5aOWpEKt8dME++9pnHEkGAFnMvoBbMjT+Pi4oJHAccL2
5YyWP0y9h9n7RfEN39AFdOIiiZdcs76mg9ACEueRz4ofLCVDe0OP2SrFMrhggYU4
BhlC44KhYswCZpdS8quiE8/74UVEkFROrx6g4z2WG98tiIhAZzySt/9J5qfUB6Pl
QJbW//iVpsM0xj5Ef/Sw5S41SjKj1hRKLPA4wDQTHEbBrxor2c3uuKMz6hh1tDxk
QSdU5FoNlVmXeuJ4XZ/YIk96FOLL9WJuWd6aNOqa3dnHurJKcJGG80meD3XowMv+
2q/o5Qeu0mffcbVXXU7Xry2iqnKaH+edK2s3mfaBzN7jUWVI579x5/Xlp+0ShA3+
3r6rl/QtzoemHhzesUrZ2iUe3y9XUiq4zGpFVylSBMgPSQzw7dfhdCvTcr6+z37I
pNyOvBlavKPo/gL+Qgr9taOhpk88zCykQLymCQ0TlstZgqPl5z/nYLVCnEgv4O6a
dyweNuVTYuK24v1+ESH33URBYLgynCUaXhOlIVxY1TTsSY2BCirh5iR+GOXqDhEX
idWsCshWF9qA5Ws4L0zEs1ZyiO/nJS8wVUoCDNysEICEDWnccPWvatn2eD6w4kXu
wlx0U2Bt5MauefLd77lv4pG+fdVzKipQjrE/DBe9Hz3OvZdVjzv73bNwlAkOydjr
dczFg1Neszxnbjs2+3KVpuWQ/fz7Pb/9Qh84OQ1Ph4WGrs773KnIUfBD3A5O//U9
E9rog9RgVWlr+qVXTr2CFVEFchM7+8gfh6U4FxoCKeI0J2kQwPv9wmD2VXAiBkF5
zu15mz0aFBEVRSywLoIG8KfbP/OGtpuKhwdahKJ8k2NV0m3ESXu8YL9Rw0GhXRuF
UxakXJKnQyt/bJnjJfhkyFh0RF++XCjZrelAgzZ4g9NaUcyZJ8snGWOAZLGJTSru
UrBF7kcSdTct4MFJnaq62jFOv/+BNtpXlnI1xyKilAuG4YJ9aTD6NAVNfe00J+0u
QQ+u5HA92/iCNFt1oY+sCHkZ5u+zb5gc+/WmUAOnsStzAQbrzAyJ6mlOdGok9BBB
EjyHcqe9WSW9DnzUKBX7hguu2E2+gajlAw3+wgb+hEnxLv1CahXIsXlQ6Fu6N5ou
NsgBBBeWyiEoYxNGQPLQLhbPkufR6AIT6Ihv5cuX5L9Alw1xVtrcefLegnpn53r1
yxHLjM8QhuW8pgVg9h4FW7IZVf4vnthSEXkdpdKgCXrOfRRyhFqchm/kG2eQNBGs
hOg/C/Z29P0N3YLpsMinPN5GE+rsxFXVh/bghB/cxzs9elEBTrrZ0caGU6NmSjcp
hDBe4Mr539zScJ0Vh54Orkg0d8nUbA44f76KvJ5XtSMo4PUuERgcgTvQs8oMm2JA
PMMgvjUJwJIh6nUu0sYOzYeHb7SRx5jIeSzMbm0aEmTHiXLehBlap8ATzC0cr/RR
GODba+nRcaEWwt3muLo83grOg7vP361jkBjgDD+4PZSPtX7p7SNYXsi3c0UMR32t
6PQghDLJG0CmIegJ+DoV8uNcX5A+2A4/utO7Qzjv3WHSiQ6+m1L6ajWsNxXPvxTb
KtZzSy6IXp64YQaq8Ozy6PeFlFP3ksrGX03QIM6cDfjQXhQlrsL8RXS2wPEdJWHs
hIfCzFVgnqbuGauafwfrcKlO0+38QgR8c5EQ4WuX/s5WfjZ2M2r+4PUNhH2Su0Jm
XP+KtACD6HHJs9NNpuiaXmacrHb9+m/ieu5E5u3B68kyi1RJdg2PKIPL1NhaBNQ4
a8n7yAQ9OnrJJp6m7p3RmfYpPMSKj11JevQQ9JSuGkbfioH5pa/p9Dz1pFZG/wgp
GmEsQYKykoHeA2Lrpnpu6gvaMVp1BKoH8kE3HDByNo4/RxB42bQOIIAziWLyXQiN
n0E54VIMNgioTNaet/r/c4O7O/2ng4Ku69kiexMPw6fwVKQsnfyTJeR3MTNMWfoX
KnETGCGDfccISw1g3B00VLOi3EGRSchSZY8qy2IxmPtb0VL8dNrVpuD2k1z0BECm
u32pm9jsImUOsgxRsvv49n8P8zj7qnxpw8MxJnyIXzYk+x4Ky1pi5/Zq43W72u3V
E0o1Yhr4KLexK+QTszk9MOlJZoVydmvQFrqgKlzXcJVopOhLxi+Wo0cm3WnHr/6I
xvF48Kzg2NZE+mGtTYiFkBqctS9eritGPynPnsq44XeB1alt94hxwMBOBXRiUW0h
bUsDmBD56mQ1K3M4l5RxNQlloilOcN9H3E95W7vMOM1+s5d7eu1hcZI/qRxpR6i1
5u15qQSOxIGTyfPyr8kCk9yFpNg5tm5t2smHrNXbDdblcKR2raVYHB9hXQju9Wuh
as5sYbQ5cC+P1LE29kprWgcIXI9JBEY6FWMjXBXQZQly7rH6VGAIoe/f115qY8Fd
uNrNdNYTczPasLExjNAQTQEOXniKZd0lnrlWzSPSGo5LjXkhE/KhDd1g02bpkS4u
JZLO7o7DJaD46E2bPKIRd06L/5ZTNnVlf5oIbHtZlSipi2U7jGHcQK3wK8FdTV90
a7ZhvpUDI1RfxvLzN++A9SRTP7PflMsSKO4ubmNN4AEaN7O2fCNjwA/Z7etMle0f
1VD8zAvmCjdcv7Dqeb8+I0N860DHZMHYviXjkE5KjaxxVMWrWclDQmzjsks5Xj2T
ra0NchHdoZH//VfuyfC9K1Yo7ZSQjH2oO58Upg/Lwlrj/5bBrj6u93AF/ODAyfzo
hmhZTNkACXb1I6zvvdkOYGZLMUS5k91aMnEqTY3R4lisAp9m+/O2oPokE3hW1rYq
8klH34uXs/9su437dPlgsf/DjgkNg/Jg35LGVTaOnaKw0n51UWG+nf4ME84/piRf
Zt5dpCAHzdIP7CyAoltmZ+CAC7w6Ck0AMhHeYR/uPrx8IvjxBGHtf4zm9nJ/xviW
RE2Af6JwNGax2UjLLSmq8gJ7QhqdJoQRw/fLFEf8z5W3y1IKfauw0fx2l8npIYT9
PlRW0gn1syjfaS1xH7dSkmmMZkAOpkAbZEsaK2Nhtt4+O+SIfMIqw72f09Dg3LVC
dbEwOXdRivYxYNXD9Werlkt+M4CUzT82DEaNoYkEJwkDPTEC3pPr+aDnSeqnk1Pb
FLY5uf/nb5wSEfeelWaDgUG3uUTSlp7aD/FpF0iOPan9nIXCy+9h4QaOQqOIAGS8
tG1K6mRrOAMdCLYj5+qXE4ZOFgoRpvccJWUh8rDRWY1TWl10CYPxXFixXcmLabyS
OI79HMKfBIJxYFuNUBvAwUIWwwx0qMT2bX5zID7g7wiVCP7TcuL3BkF4gw7XVdJ/
hDxyhKnM5ROl01n6jFmRaOSSVs4ys7X1Ej6ubAr9VguVUxpPUuIF2NgH7N1hB8GE
Q8/kPg1dOtcLkvtKoQns+50mompxtaI161f6ELEoHATtULlpLXrzFGe4rtfutgtc
vWaA6mYt1bqgfYrj/ouYjzwPARG2A3wsYt2oHolTbJayHZqf3e5VohgSNLDb8rno
WQ6N6gVCyMQ84KYNd9Ma2tOHGtM4Twg6ZpzdpipEQD6ZBSuu0I9cm/OOgQosOJr4
hZBooc9gEC7ZzE8Q9uJSGLlZfY+DVFKsQcow7Ne35MBLTOLiwfjI8WG8jbN3t9y4
T2MiOm0ffQGO2gOX4hTJNF6C3dRP7aP0klz1jgXkujvkxnKwrzmiGhKLBkc3UnhC
kUlx+iGKJVlHRd+ztoCIM6XQYhPVH0W+0lcV/bSOEPhsuib0GnEWaFvULqB5ntw5
MAyIGoAD7hkwH02LyFCsqmXQDJFBlHU6MSSC+SmZVDQwsXZeqtwZ68B6kX4XBzX2
zak4xuvs1t9aO8ew66wnEvF7Xh8CvzIGSn6GudLYQBdcARRO+KJIAbgc2z/wgtKQ
Jhn4ZN07YL/zSfuctTNax5q/0AoJO1IU7+iinkLuNC5VGpoDu/N6DnB06pP3WhvF
Y2wDN3kZttH7S3Q9DLLxzaiz2ZnKT8QKfmvFBPHBpwPfe2/RegBY+XxkLEhBUPoB
ELTB7KU8VrmjFCFzM4oKaDE68RUGOSjRc6e/MylQ26IknWhteo9MVZ00sk38Fuop
ab4twC6vNgmcdrcEgZ9ErGZVM7MuwoodRGX2Vnz0xg0OhpKZQRTsAHPaFDLNME/w
yocLWu3LQK/1a8PLElFjRwHSBuxiA0RPcuRsnr58VtX2hlERCAjbLhyU0u/VhvuP
WPBF7QVAgO4686oHu2yhIRF7biUJjwIxbZO0cM2jRlsxnClZyFKvfQ51uqDs62m4
6P44yqs+OezU3/VB5HcfCF4DLkQgTqMfsVLh5QxoOaB7PuWskJ79KBLDBC85II4m
57lGMKRE97BGuBKmyYWH/1o33jc3GnyNyqpu9VpC888w2PJCkEQ9AdMA27XoEnp8
bhUFHnTqg7be9KRyNwBI6/KkH4LGEhJjAc8UCF9j5Yo1oN78BGD0c90v8nN4NhpE
XK7oddyZzk0qJd9zW7kT9TgvXxYCK+F1FOKbCmr48aJGYKhIw0ISa/IRi6Ky3LtI
8n0dCuAsX0QgBrthBK8osFE1U43dCcEfKRf8xQPLHiYD8Y63yngZ8+Em5y/cr1zp
XEVfL31y6NUWWcRb0eukWCu93hunOo1XizKRI7Fkhm837zKd7cTDoSweO0w6LC97
Bu2KkDemLoLUs6uIu4AXPQLoMEI8j+umRNkQMOLvcZrHL6YWabtijN5yNFTIOk5i
HgiY+MXg0/1pRjhvqod+t5k8JLKKayxLe7GHzYis5CxixIKExB4qeCf/LTRN9uIE
AL/nMDrnqnFTii4EMOqeoy6dhTQ0XagZuE8W/qnPfY0zO16IKMEfRZ3IwjFYwZhu
+iCHD8qdyL9tBSkDGElklMG6eapzzLVSonKsGGzf5Yoid+DGZJ2uaca6Vv3X/YkT
cm9nQYWznvKCLcKSaFB2FO2EYVAaF8ZCjDosjd3N/Gg9xLXCDv6YJBLqoNxbbo+b
97AH212f5P9AhR8qt8gPVPsbF2viRnf25KVZBBApkqamaVziKuhx6x3TeC0V4xTM
oiNqE95YtJHDMO9PFGbLVcXkU2WqUnt33cTUHgv716ORozI1ukx2UZXmvJTFIXsz
whtA3ldBQV7JdT97W8LcqJscIgSKaqkAN1YuFpz+hd8rfyt4IcsW5RLkvgepmuPy
Ol+iWMQ1XYJ5lh3zvQ+gT4EVRAa5WHjANapSvHU4uJoiaaOsyv4pKfU+/D9uobLY
Hx4vD18z7ejBNJNjc31GUYrHENDVhtmOJ5VLUxoPGDn/KkS4JI1e1+ODcfsc5ETF
qZKjElkvI04W0bFV+0RrTKCkAE099+sDCWGlT59qhS4Fam9Y1XFgSIbM4H6c9/VP
wmmR74vFNN2CL/z/rWo0/NvN7YWzBn/Jsf07kIwe8onSzvAjCT+woZMt5kNAgMnG
qQj0d+4xNdONBJfZ5Z+/I2yUPXczckn+JZ/tu9gCUO/3iBFA9fUFjGsf2Ee4536J
o1mDPsZ1MOCOcWsFopyNE2vMYELdvGgHSrJ4kqQgEPSdSB03eAjqg1mv2T0k7ny4
RPCNCKXkslH05Uh501AXcNse9Y8h781LIwY2Q1MMUdsb0Bj5SttxqHTwuWmvWmy5
vU6EDKiSTjC6dBIoUPwhaAjXlk6CoXixkB0SHpcsYrIxjzZkGOkLv7lSjoFyzbrD
uMt+ETUXqO7XdMJNiaFbnXzNeY0wDerBNAeP0FdgB2dtBhRbESLSd1GENeYxdvlv
QZY6AoEH7nndzMo6o5xsGe+UlYmaG80ohFnfD7jyPiXP9zOQL45/DETiSZumwacw
dOvgXcaNJmD6XJwKqzNuwKGFrP+IoXg57tKh7rxJ/eBT6+AIxjq2Hnyt3bP884G2
Ak2HnkdAN3kqrvK0ap9p9Z4bHeboYHkUY5EjgGtTseaulRpUfZnt1Vs0i82O//Yu
faRJvBOiIjGgNwdEj1xWq9v5QF0XWcm/DvvDndH4YINu1OYIJSyMUcphyEI4XCbs
DUXYJxWwFODQpFyMVz8pRfkMQGhDCQosIOTCN4SOUcby2oq6HbbN8ieZyrEKVa/C
BssktM0y08f8Zc5CrFhl3q+5nGB/gk3/fseAbGpYXued6L66DM+dU8BonpcyAeYx
7foK2WS54n3OrpkXu1/WzMuDbQ1fK2x1kHIIyRdcV40LlWCJASr4g0lwFNKX6Ko5
BgZc35tybSbcSG9vBLjvOguO5vMjWqxZOdzDD/zs6I6hRYe/myVfbRIq9lYAF4wR
OZAMBC1FPJbZgZLE9BOYFraquXqrDwab43yXjM/M0GgL2kp1ez9ZwoY8n19rGTno
OWaRr/sLkpRtVFhyTEYwRQdycKl841yXBR/0XvgpEEZV2w6bUIfAHprmNG+wg3I/
Y9EgFQo6R24JQTRv36fnG7m6K0Bxyl2XbZNU0eY/d7iYP2p1yTJRP+wonYQspuWr
bMHQ1ajUZo0T2Zuh9aHrA/iORf96z7FzUhWGTATvxSFHq8FucXyQHg0/jmEh8itd
BHfTyf0uvT67vEkaBa1+cCi6oZ707DWiiAeesyLA/eT0z4M6xXmqQzZuQ4zuB3/o
fFFGZhG6m9shoNUJctkTpMRi+Jyr1ep8M/dnN7JFD07CJCLjvOXMuGId6GtUr/uZ
FfAaNt410zn5JRTf1drqU5hBXtIEE0davV1jhJkPq3IJX6a/ouUd2anAapkiPkE4
Pa40xKyxLgiOugwdCOOuXoxK35Y26G01Ldm8pRiKzdSl9K62kDUTowQp8oeTiFqC
usATqC73N/jIAM0hLKOdWHud0mCN8AG67+/C52xZDHbFu1CForqheScXCAUke5j4
tMODHmXKieZ9Jv+glPa7AR6KO2TZjpOYmsTGasCQnh2+Lqk3RNKamCuOeKLIV9fO
27fc6K3sCiqrYWQbIyqHHyJ2sxEPzykomuwN1Dv0L3zCoNsvDTV/BG/1iPfbxQVF
98Lh5qslNIHBTSCVw7pkaJJZpG3o0fpwkwrQTM/MmbuPbiu9QUx4EnZ74zxEY3A0
E7YJ0/lSr545T2DvDgIUamgO8Jt7PYk6oF+DoP/c634x3YFi6FfV1YBBguGkvftO
KmleDynK6u8iprMYQZzsWHFQUH+LmQ3UxigHwAURmPQdhEIKzh1Gu16qti2TBpPS
Ql3I1qBHNX8Mzjz1eZ//7ye73tooMcMl6OhvOahioyawGH5BK0gtAWUMr75J/K/h
TFZtjfnv7+Mun7hSzJvBdXRjp8ziaNdFwczMJZIFVaUIVrEtTexHKrVQrOycwu/b
7h0GUjRxkmexpSOa9LTbzpifsN4+y4E1wc8s9GVjTtBO8mE+7i1Pqzl30FKzS570
kHYBAJCEZnqPEDrLsyp8Wytrbl3bMuYR86UAR4kfq3y782el491brDKQ5ZzMItmp
OXy5sd9OMSnM3ixmE+xRxwJKW7084X3ImSUfqXTY6IqOTYtYf+9Q+9TJiR87EP3C
1QeOjjQSLhsA+m8sgxZx5OT8jORK3wasOpiMX/zknI7SG/Ms1V5Jh5sQoMRFiNfO
2spYDVjVD/INSkDqWhJ7aGpZewhjnKz5cE2vc3gvWm+JmdNZf7AuL/ke3psUY9yg
Wl0xa/MraQdoBJb/KkdSDeYfgSUhTbQek43tbFLYXlXfxRTr5Yh58Jffi+dhzXps
kDCfHy4L4HRZ3w5uWV1/TvSZ6qw00PNgQTth6ZIxXepSWKcTLVPThqn1vzbDqYiQ
SfNRDyBgJqpyT6+Tp4r34gD4p+c7WSXdyqFkhEt1WKb3EIWzQgkPIVT6Jr42D2CC
O7MHnHA2fesAcRr8VFxNNuYz2dKVgNfQPT9WHUJ2c23C462yStRU2feZb4sopWHH
FQGCzIPpOj+1OX+yPSw88LnEsQwIy3NUgmMTeuTRAsdg9+kZAeT/SnKKM9CmA5ui
k2jlC0qqZDbsJ0SZht4M8HlUL35V1CXG6f7rdR/lp8tWAfexReuDkWRP4WXJWrT0
2lkXq1pwv5+DKRRBkLyk95kPkX7aDjqkkMkvovu1tVodxrH+LhSyLM5Le2aiDJnx
bT6IFLita1exvS9EKBU6kS3h5mlZa1fdrG2EnI2skSxZTNDC8jylFwsEvDore+XC
KY+9IBGzpuyTz8+4sA1xPQkDMrfyfO96s4vT6KvY82NAUyI7D97yEEko0FONA+jM
CLaBn2UJHTgwsWvwIexfootnkXEcrb6ArpcxCxs8OzxN8o6jFDHGKwol3OWi9o3/
R0eFpkjD192vzgbNSnWVOrgVFHzw25ikZQxeknRKvTyLaIkXkfvVMjUaVJIWS7w0
i43rfGA5ir29BOAqhXYAWmC6PSN4HQ/LqecjZrXvAPodMCvomQlI9Dj+Emzu7WRv
yADpJEZSr3eCCOrmCjR0i+vpySjIbWispbBygM1KErR/edHGw56l5rVtWIjS/cZm
n8K9/6m4PsJMEZ3o0C1TGgF6EXBtEeZhh2iDjTnb83K/mzTtorHpVzM/drkjIl0x
Rbex74Q8Tnb/02WLchbEtXWvhW2NkqxhbnAkaVHZh1cT7Wzivuk3D2MCl+XhGxi/
qgdJedu72WX+LvfLzMILq+oG2v49gE11vWUx9/eEbu0zZuuWdTc6S86JE8G89EDl
PpWxQS3t+hN6Elvq2toVKBaLCy9mENX2HmJgOuwVKc/bifR6jWZrXof0m3dAT0sn
xiRTFEXPfValWSsgDJM/NoEZnKt3qzoOmNZ/Rpsh4QE2zg6IPqKXCrJLEM/skSuT
VUmojLtXmp0atd1KiRsC18Kwyuc1nwytGGlMU22QdUlbepVFkJwBTY8EYP/eZSSV
SYXeUAIwaf+FVhGQ9jpUpLEXm8bZApuSgo9GYbLeUkOkX5iyDgoBqqh3ThL5FQ07
LH3VOO8CC5QeRNgV43YcGTEMsyDh9lV2kHZZWXynxDDO7oQNPlVDKlcYGyYvYotB
73wRCiTMzIgjijNDQE7sXZE/52XVCe077m41AQ9sg+riDZt5/55dnddAN5Yz9pgq
8N4U40ppGGbAE2EkUcyAzzQ3bymLnEQJWqxvx9MBHB+0HPCNmfyDVem/HcwkgGmk
BbjtYFQWsjxy2PdfHOKqRBjVLIligjybVLNtK2d7mSW058sOp/OYpRcP3ntkvcoF
y7bt31zgqJP6LUn+qDHtfGBy0PiwFIyKHe6NxQyNgV38BCJA3TdYYA2hmJv5KBOc
tnxeQWMHQV6sTou7qhtMeELU2dMnjUbncdiidDXf8yT3Ooha4OmKTXsIkEPgH6yh
33Y70wkrBxc+DuQuuc9Pc4LBc0umjpf5wiy0V7JxemWcnMfzTPCFvykGQKlk1zSA
YGiJvGbcdlcoOfuMZofYyNGCAA0ByBzukplvSaauvYhbj2wfMZEO9aWBRpAvS/4U
Y6TiufnX7h/sewRCBSCb1WFu4uiK3NY4vbrhhXI9WxgglC+gnaVfvGtP1vF2sT2b
tuYkk4GQrrS3+Ejh6XTBxAqtwAIuRZzeFPp05ZlJik0EAK+M/O/PBxpqopgKLEkC
v9shkUPz7eZCNghiSj+bOhuvVz8vJ9pWd0u3uoZQr4m3pO92yghQ9pusLUj3Tjah
jrxXps0Xoijn0ZCqEgZmED/NW4wkfpy8xPUdUpTujIdVjcPOAWE8AOUxX0bFyYpL
7+14EYOtA0860fKgvhzcA6o8hvKHZfEq+2iHD6292yFEBXKtBlKPQnz8NE+1J+bI
0yPGnXpzkzfD2TZeJu4N+IW8J0kuElwkBOzjMugp1MRm+YBLTyAfQlrw55tseAK4
NdLRNuvWNF7P9AVS64gIhpr/nh4IU0wJwCSWkrY8BV9HZvQ21fShE+aTtruP9NMt
I2ASCnLFD/5lj/KzYjLgLkSlavir1iNrJVqn7wr+uQA1qTql+MtM+Zts2PCL4wYM
Z25AuFmbFDHrtPG1jbm/EmzLBi0frRrvLqodGmi2oPG8zgdE1sk1ejcERNcDw5oP
3JYKRg1q2wwOSXTaRTjt5OBWZab9lH6II/Turq0sFyA9LsCprKwbrNFUNGpKKH6c
y/7K3AF7ASQeFHuFeAal+xAXlHC9/JCUPpG+5xibatZqV3UAZVsSDaVxz3xb/2Pq
iI1au68QAm94506ONkUu7Shcf+J2ArcvaQ+VjC0Tty3TwYv/D3goL+JN16ehmoC6
zaebqDFbIrz60QdB1nQUF2WwLqxmUq9hlwQqtiryJDdyIqK5B2/A5m5roXXSw8m2
MfDvPBRz5u8QgHzcqrFC45ixwvltLnSMAJZFZ88CrSTo3bBTsHk93qbEK6+At44L
uux8SxHVxK6wpQEX4TX4sCqh9oO5CxK7fp6G4JwICtel9CN7RHQCv2iPAF+5/NPr
03pp8RYzRBoTQKroQfp2J8exTpN16cU9aiFY8W6pHbrk+zCJoGAqtLxV2jz3rbkh
bldCqpXtL8CWIkOnAxuUc9ZPjMAKwdYkGuJvcW97nrUtZELDjZW/oKRw7RfS3xzz
E0POuAQT5ba/fC7t9ZnZWsS9VhlcOBpPuxfZXOWKnGtq2ur/MpAaaJ3t4A3JpEuE
aAqAlfdTA8aE8hyxgvFyuSSkRfiBlYN0YezZkJX8AtqrLf//R6BWXlxMs2Fx+ydB
idk/tRZMdS97u2J15TYSoS/skKhP105GrAryB+nDu2ezL06PA7owhBqV7Y2wZRVf
8LOZApLLoc1MzvVQD8YQyEWU+Ic6JeAldIYuGw9XixvX3GsJqaaWSD/t3BrDLyiV
FyadmDcZ1jUqiTMySp1QJXqAJw8RrjMlTIjTaSpa8Z277otjq0B1JYzrX2HhOPZF
Y4vezAYxkhxkMCiWK4M/pfmR9ChVvxKD6JQgJuyKd7SPkZGHix393Y+ZQa+rX/EH
JjDq1XaiEbg5/vqNlVVyxa+NWQIAriImmUMrEJJN0hIFkTWMM/HqY+RqrMn5CjUC
TI1xBLzInnGd6HD/DkMgGu9vzeRv5lPDhjI4LolOS8Iy8ACzFg0zrQ8AG7eRnvWb
ZYE19uDc/yNOtgmDyCKFMJZWPUi6F9MrtWOGAzQKo0wRlSoAD9U+PEY6MnkdIjxS
ceiVKR5AokpMfN/i5xx+NYbqClP0pVp5329qzLv1qZYFWc867O7g+soQHt0D0Xrh
Rwe0rCuVhtK25TyZcOhmQmHHK9rz6TlbRSLhiCkX02EQWs/bc5hDNux9YXE8qQZh
ANLWtKgCgP+1VBPYTFwQsJVgbYzDhu8AnxkoTCZjIeQLPh8hhFNPs5JFnSvlTPYo
7+Yhkp4QEgUxS6iDJ1xtSO7GtmdiyryHlO6j+f3PxDhU9WIBITEIF2z+9dzGUzQe
rd9JxsfwLQeth01ktSuPGUC+iARvE0i5dEMxdXvDdaIqwMpMZP+BXnMzug8rs3XS
WM9BwsqjMYoqE1rLhdwWD4ol6MiK/M0wwHAp0kKjpynMPB9+49UV5y1FruCjByeC
KCBdbrvPsfCtuoVMtpoN0Iq2fPvH8zYqTqcjyJhbVZG5gniWa1r+fTc6jgevm+ws
oymSn8wbI69TJQItnmMLttnp3y4LLuIVFWYyB/7Ww/2ZPIIeGur/6Ay2tzCL1f2o
jHqXXgx3+sk7zywAIGz6u7XX53H824Gz1MqfI6BC9wKFB/QV4yGTsWhvgGW5ydGJ
fkkpnld8GyEMdo8bGhc0RWgnY5hZxuB54oE2uJUOMpnak/Cv+2ayKYClEnM+Es+F
SYeZg01mN0WgLmifjEBJqUmr/Yvz2DZvt5J3Bx1p5IbIWKQS8wWkNBcgBkGhqAup
16E/635XIpFnIUaMwu8zRKr55vhwyJfenNWGAhTc2dntGDVuFp74FVJkChwzr5R6
FrxlqUGidemZQ8ZtIatbP0zaMYEhfu5j9Gx2x7fceLXjfA39mcnGa/k1ayPhfsdt
Doyq/XZKCtOaAbO86rWjYIUN23WYsM+0qHC55FBE+DQNNKLSL/0tIREt/nN/+Xir
+yS/MW43lHaq4So/MBBtGEa1BtbrgLc+Lu8uWzbuqxjSK0eYo/068LeeB5Wj8VBd
rov8HAcidiE3QM7gUCsnf/YA9DxosqeMan/qCmlktQ09AyKAw/fnIkkIMiyz7vTe
Y6q9iikspdqKoYZBLgjneYyoiKC7ojlCscUG9ycUvoL9LwAmrq6a6GGfJJ2EN4t6
+qqn5iO5Emc2bBuYWxrc07hC/WbGQEGTKA0ra1Bzl5XUyDdJSb0h8lhLELZ0vZM5
RsIabErYaZU60agYGV9U1+rx3yo/Qh0cspkhw8ppcaRaKEMMk+XDSXodOj1JvrjS
3Ivpb+8LRnJUQlg6xO682xarJs0/LXYHlGpvWYuKYy8A0qGcDvFl7lfbnUNJm5dm
nkOuzRYI/NjKSyPlyKIjXFQixDu22Ih9dtFKn8WCUE0fGV4RzlI2TH7Vqe4Omok2
8piSTd78/rdSBlnaI5ZDlt/scDZI7o7lNjVju5WT9dpD/cH/PpHJB/wbDXbweQuY
nACge1eLsPMoPkph2Oh4gtNJ23oYVG/TV4to341ht+9bhmj4CWtE58XrgSmXMG1g
M9P+iDAuMBOy0rhkFU2UYYK//z0OMqQjd5mulX7H/XUtyZDsNBDNle497HOein9A
R9lID3vtn9gEcCYIp0cVZydF/n4Gqmn+iTqYONzf71Eu9ZHrWPlB4j+becaeVp24
1LHU/jDOTZxacJ9eQ1efcylbEcgAEsPRY30JcYD0zW66j+4MkUPXoNdxyaSdtnnZ
6nXmA0ngjr/y0BXJqIqQbVWNeMh0j56DT78LwJbrB4HSJIRkfurKwXMEbUspTkY1
ut6xyuc9CMTiAy8B/v0BwsE1MkkPT40Vc9qHIcHI9K9ZrpieYDF6ZPoJbiODDPtm
fQtPn/dvCh8XJpKIor/RnIb1vEtZNcbzO2+abCU1X4kTEmeNQ1dqmZu+Hrl+WJaZ
y52RG6vTeOzkSk0sHZD7SejQDxjz2CCjIQz6G42F0obpXVJ71XeW2qa/AEJbzNqP
ZL7RHfUd3EHfTCUKtiGmXD42GQNIpNll1BPovqHt58Pnn7QNohx2kkOIh7kpfG+6
Ty6wJjjNxmUiXEv0+wbuMVyRTZSdRbuzLqBQR6s81uND48b9rVwOJyUddLfVANL1
a00OH8YUGl/jYAM5XN/siZQW/c5TkVgJBPw/12VdeV1XDQ8d+lAgofRbfeZqMpH5
FDl3bxuV174ZmEIJt6oRf9dOLwBX1dww2LUAgpmO3AyAoQ/LFBjVa6F2uRZyhZef
oahhU0bt9x76A3dexf2HGORtYRNUPSL0qO6mlE+NMsKvt9SAVvObjgGs1LEXhxM2
QgBnw/toVEmzBsvM29fuD3Kl0S1bCOma0GCSuFBaWQq9y9muPbi+n/95RUNXUAY6
faeH7x7NI2RxwMqg9Jg0EB5TDJE2yAiCTjd+PGfriL6NOv3mBdnSUN8h3S0sanEZ
rWzNxG7qLYtUwFGXq2px2p63ijd3ySaz5mQqMar8RY1Y7SoG8qkszSi2u9vMRgSY
PQXxTNhxQ6Hl6VdJouaRFYN9haQT+pcQWvW+gOI2mA0QyNv18Gm0GuAq7vxdhvfZ
K4LRgf2BXIry81LUl6g5mv/xOV7JRZSSIdkcdOWPFkSqJqwtVeX5cgcrghr3T7ci
mjbkwJ+NZegPaRQSMnYAQMpYHF63hwIkydIhNtgadlCYIDMpRPJHXvdi7Nh4fBXZ
RCPsS5pMdp5EAZuxmoLxVtea0/NNg1fG8xMGL/PlpuEnF5Rn6wjxDtzWnE5hgRNx
ZHcvel/zH5Rc/hqYdxHLy3nsBtjPf9NKYRg6JOgnKqg9lS3o+vBzVqN5ZHte+RUX
gesGBjQBVWW+plOyAqNahcAwy2izcv6yokja3/3GlDnRWcpVTk7fzBL8J8k3tbOY
EFLBRqSfuzPU48aiWM/Vt3XG9NIDUJPJ9hbvXTw2/SLPC3bsB1e+Qhx8n2LCy7QP
e6HaMGMvzmvVliakBU9/89RWUGwqZuY9nZJ3bUdFzew/6rtkiPCGtX/6WnfXXMse
u0s3jtLgSLt4YEoWTUbaX4elt7O5wZWYwu43n+4IRXRDzDUm5XXbvbAiWChHHLQh
OucET0VwrIyxOLXVx08oJROpJrqfm05MTrqQh2Ll2+tmR1WLsnDRvLySdxdyTfUc
GC8+cA14DCwXjzMjbZXAwZXcow2wvD11QEXRe1y1+1tF2Ey0gvgGdiPY5VY+VObC
ChdwcDWWW9IqT1h5+IXcnfvuZXfMUDtR8yfO0LGWks7cTf9mRK7gNXpvXr9Q7+iw
AgLNi+0a6K3Kk8jsXluFHBsQlNOWNW60Rr8iKx5yQB/dzG2uyuabTFX47N21YVkW
euF4PyhsPZz5PAD0RWbAMOjcU3fDZQbqCuNM5R5Nac4ZdrasjUlMJDqMvwkebilx
44T0GXLtWIsfr+7M4S0YB1UGgjOYOwLidUtFMFIHsSMsic8A90ZOwZGPz1LGGvyu
Y2dxp/b699oHF8wDo4+cr5qSDmtBmbVl1szMrxC5H9c8RcsBFGk/gkugNHo0hKzq
FvSaAu/ecUcgUhtq8kc/bUQ8Ww8z+Je3VYnPZ6r9OeGq/j7zX0l0g0DRsIW9+/sj
jgFAPcbf9vVpPLe18TRIUkpf3CMpZMLCpnTZrAszDBWGG0lPty5MPhbCkNcz1Yxo
aD1ga0FrNob0+rwp8w6Jzz6+rksL/Z39ekUrOMnqSVjmia6gnY61ObLcybBaQVhL
8EO+0FEWel3Aj2yRx2HIIupERqZeQAxcKGiHaf6ccYN/RQh38vev0/5c6ALBjsyN
mfyeJfS4I/xuTGWMur9AKQn6Y6taMRMJCqxkjeIqaORI8wjn7h5qLWuZshbAg5jb
9GlSQho3xzLU8/e9keM1h8uS0iP6aFHEB/wqkypxuClY9X+pvR7wvTwdMVEiGA7X
p86RCOqXq10e24+v24clogb3dz6kLRI1Evau/87/M+WxeKZzm+8942Uf+lwGTXks
BrIJJCvTg+cyioxnYDY3VQjZ/VV4DOHZMRaMWGnVZFMYZks8CKrXVxiKwGvnyI6E
cwEFx46XnEMOSuQSjTGwAFBtGQdMbJiN+WPZIC1j9yVY0MMRPoEcbdMOrJd7hpDw
zWX8oqKzeoyKM2d8mpS3rnDDIpANRsHHUnF2f56N5X70jiCYWfHI5X/rKXdxaN5h
nbzUDe9nWtxHPJzQNaexaIq3QFeXvYSqnpDm/Npro9yqIVDwPBiRyuqM0leUbL7R
IRoQeUNBMiwc+g0tmIEGmlh3A36ponom+tbZxk48xN2jpklom6YHO42BqtDwKRSh
kRivjicv+Gze48enOJ9x85pM2iITbCKooCqg1u9BcpKYf/dJ8IoF0F9XSzhvVi52
6ilL/fsIjtxHgUyZ2+pJw5CrBMzZi1WV7XtlpjfB6jZ4VOofGqQr+7cEOFDyi2fg
hTJ+94e6PgNTp3OAPBhff6Uw5Tr0ZLYQ1mCR6rXlUvH6xre6wbJxLjsbz4ACXuhY
8yg1rI4yaNRQ3DNPuChfrgueOvYw//Uz1b1NCw6r60ng4qlcY8dha/+VqMwvSKax
g/LmHvWAFi4CU74SMVaA4P4gK2pu2VmdKBBPqPUEbNavWBYabsScYf1PFltyd5x9
a7g0kODx/AJUHKK1oqZGgE0Ci9s5QP+uiln55SOVDQfLQDRh0FXeRE2gb01MJW7+
zic38y9jMV9/mHR5GNM7h9yMMF2iHBCgk2IZVplqnvMQVFvDn9ozsOFjRivFtmgq
JXgZYJCmcwNIXf/hh3TbM9UuOap0JW1UJRv4xqllz5oc3SG2LhPvJRqLmufbEyLe
y3B4XWZ6YUndgyngr7IIfYAyIuOJrdqvmQUIT/ClATDedC3E7CuiO6tvqaH/Eicl
Rxwt0WSjhBOpCP/gnDatI4PU15neKA2EdVOBJeyHWZPsSCNKb9z26ZNxDA2i1FtO
VKjxPNUHg7O4H3GhFnevSg4Wo6YUlkyrn0j55k3LRI8qeMIWHQF4hVVQacUCoDTq
tjbs/ORf81b4VqJf4sEG4mtpPnVq14kFARLiWxS1/oAGUa6RzBNJ19fH72LpY8X4
kvu73wgOkFDJ+jtVxZQb7Lh7tQJcyNpwbjut5bD6fz5WtQ0vZdVdxE1XKQsrwhY5
0v+Nd/8bwvA+O8EcuGk045GA4KVaYPgh24meAhXndvYxkHFQC+EiCGe/WKaPYGiA
Yrit2n6lWmvOyB7diL27i7vd0hDNlxROjcQ7fEd/rnXB3jl5hoz7cCl2GMCbiLWW
W4og09I+aJHQzvAC6FXLlWmlCrPAvbmbCXgFnFflLnufNA8XM3sqWk2YIMlwnuO9
7HfNnEPSp9VQZu4yjkSUkzYJUA74DYPukrb9AgKmpvbZNjW1MG0orax1ZoSQT51W
n7YT76BDVQBsjJTs4ytYOK1oMS8LA5PR/BEIASL/nhYkg76vuKC+evJFsm+PeNS6
qJFGCWAcfk+tdwRgw9403b2ecMbriH3VG+tqurrDs/C1a0gGzl9UonRpebKZjkqY
7SIJ2Oz7rih0L5CIMcIdaSwAJ+SxDYJn7a3DWFmD5aPFbhHJW6ygu2tD4TPNm1t/
QJNnOvF85SXNxOcLe1knu+QnAL6pqKVULYOYUTFp4sBoTaebzSNQxJdDd19UnzPr
Ny+85Ryib0Sl7yYU9YNy02NDqq5ufLiLxdhpZ/LpWAi6iQIV+SBoI/KI2veJu7ED
ZJrfGLW7vGSM/D944RRZM52hYqlvFMD/Xm/vqw7a+lqWV5eS1l8fIEObsyvVlncM
Op7u6TKWosGVyMVNVCx/WknodhZPG5/VlVo0BI6CRgnhw5cdH7KH0MrM6t3r3jBG
a71bs0SJxE1CjAwy9gGFOVspi2TPFplfr61Vyv5PZi23p9fAFj/ksHgiMuqw1Eva
AKg5el5i2PcfdRk2PocLhJjAvvouOA9x4cDb1xTsdsvPol2Zb5PSST0pmOsxkmCi
sJqbtX9KRRwOsxPMxoNEfTSNQmV82EIAvm5lv5/v2hP9S+6mU8o+ee9WhM/Wvkb7
SB0OevfdJQkrZvat9v6FUOTzGa+D0OAPvBqgNJXn6ga23fJIigpBaybln0lMpyTf
bTw2ID3lzPiyEKKeHzom6lqRpii21MoWuy1RGLfv3QyZ+B/T72s6NsLXlMqPipIR
YQtmLb1KTROYSbdjEwPxzWmdhob7tQf5j4t/ZJebWdbJkWOavtSBK/r5Xq6MdGl0
XaKF+I/XZl2c1MdZ0I4vY6Hw1zTPE3a20KvHsSaXmGh+aAhkJtpVXNaBqIxKNOUV
6gHZgD64XknCaMdTr84tezL4bYyRUgYcfjGGY1Q9zOtM8N+VoMcJ23OwIXE4gfdy
2dk4xsAOduIXykzyZ7HjLgItjgRggu0XC5P11tLZvl6kuEUuyYMkKFPON+TXP9l+
kuAWTI0yxu3ipY7fMbJmU2VwOSkPXv1dRpUcx4XNS5l3lmFoOr7KE/SaVBTzoMIV
jgiGwJ87j7+K2+mDSes0Os/0Z20CR8Q/e4KlDN4rqUFQ1qDiwi/Oi1O9Vke1zcdi
ncOUmw5ziiQyoBHk4QfX08XZqrzHqrDzWR/L5JrBCiuwQpc0OysZ1quy0qGFC0SV
6gIk2NE0AwL9eqNzH4R8vznwV95y44UbFhNoVtExoyFIWy7YkA0+mvawUhF5Z682
9i+AferO2zGLCqzxeLMrWvR/XmyS8xDSnjkP94xmKdKvt3TlNP0AC09Is0sDo9WN
w6sDPjEjyDhCZAJlIz+LqDfoTWscaUI2Nt7/G67Ul5+5dwSwzAECD/4rh+mElYdD
ZO75zz6N8Mp4jdvmACH4EpN4LJB6gwezOPZKnEnQAdzdI1zq0y+csCByNO7CDuUf
CYScrMbJH/+eGbKI9XQWFPi2CRrgX2vhbnNKxupbbdlpAWL9h9blpyUUyTlBDffm
tFFJlIYabBe9HhDnJntQB66fxLcW5YpkgkL78OGCgLAJ0WfflUVyacCU6zukqI+c
HEKpnDLw600FFkXkL9TGf4mvcBQ67+I4g9XAz81lcec/bzYFEMBKXekSib6SGpZY
NHcDK2SY4DVmzsuivm07yHA7xUhe+zpwdEkpju2itekTLkQYeiSTR6Tr3qBb6mYw
IORrn3zq9OXsR5ihVv8G/mGPZxm0gLdfdNPQ6pNWm7XSv8ZN8L2cd5iSpiVjheEh
HgBMRdqdE74SQjWHDm30RnZuHw9/kUafdYC+hXXXxuatZYEAaZwaoijpgi/F5L9M
jOkH826Ksc1WibNui/vDrKW2YrzEXivPnG0Qj15KG7bz98Vl6qOqFwWTUq1fMeI4
Sk9l44RrJJ50fbf/OM4ETk3PWMB9+ZwJLIjqRNuN/VtzIIqpTr0xBj6c9Of3PQms
ga6A8/0cvMXojrDZuU07d09dpUXcC8qG6Xds68ta2ghqck9Rz+9RT2fSGDcDpKEm
5QItKnLpPR91wIR98ZTq+xeHU6TWDbs0gb4Q/+WaaqyZjXLBrynDE+T6vBSxtOYP
dcDoDJxMBYUCaZnEYomYZNmI+/vTcZG4IF5S1tX5WzM5Zj/aiajPN8ZMjNXlcXZN
x7T/MCHwTXeyiI5EWHU40hZQG7PdHv9awRXe7VC9Kln7cP5eETd+ASz2XhYCQRCF
l1oX/y+vEPrxQtfcVD7iZDEmSEeDQ+pn+0E698+8TTd7PgogCyCdLc8TDnN3P7Pj
+Wa8TtK4IGi6oGUsampifCS+rLWYbKBOLlxoXKzGmyemj1iC7P4UEOYb8tUPo8zm
5uhlT4mnMJXmNxBTrmDVqMvR3Ov1CHlaO9dLarGW/MEQwy1346NSkHnBuwmSoLKN
Dyfke1aTttTOudAcIda4aii86jigJD7vsxoM+zVIBwjw95sl02fvIUUZgjGk/Y5N
xuUDAtdw/pVjOz5YpRM9OpSZiOLPzvkdQadj4TbtRT5gzqUhvR7Bh1JasVeXKgYc
RJ4wF8DttkbtYRMJjc+HJWPORLzBgdNrlfmw228G7xcvLDKNYpM1Vk6QSRZmtD+z
bRxNWXvqtvLphQpyezKOQdffw062jJ6bu9So3ghCM6GmR5zzX8T5xdNosQ99Wo6B
01L4oob3IoGXm9DCZVtE08vDq9hZhx8Cv7RBsImONgOLCnUmqKYsrEdV7uLYLke3
tgko81hfm9/DSiKs1xNuhrqh6Be7RJaUTQMrcizZpTdcIcrVvSTBzMGygm7purLy
H3kPbWr0iKAh7fIDYbstidQK6WMdNiRI4sxLFkOIUhNyGF98Rjm+cZsXly0/Oao+
X7z59Ac2P30a3P47xoQdfjeJgdoqwgbI/pPZ/vthagQUCDAeo/Sc3TlVV67PE1lt
kqjqqXVioaeQ/1a7bJUnSGvCwkqmmSegyNRYcgJgYNYTzkcpZ0CupyDvupwuGlz0
c5Iyme5lrC9XlbEN4+yqZet2KXX/DpsdmEw1YHUPRyecGI2ofe3gtJy4ZRiKQMEa
MsPLRoz2/1Bponm1DpqKGqUF00Zv6hY+IeXPzxQU2doNTVULJ25wDkvkDnAkZumm
L5XXHaeQnDTQsN4tOU7Cbo3+1d5X42EI5hOv7zZSQ0ZaQkXdljoi/awr5YKAVkBY
BV5PW2C2O2hS6rNgDmoJ90eYNlnKJKrJ9YfhuEB8W17DKbwFCshsXua6AThoutC7
gkLbQddfZlEACu+djF1owrE2lhZ8Y/t1BedPPp6Vnv+PssypytmOoQazp+aqqKWC
dkSa6cPxSMmttYGhron3fRJ58xSRSlNfRXRr7o7yme1IM6KAueSsjkE/f0qtAjl2
iRqp8O8hO3qNuP/93HFQ+RSywuc9/nOcnqtC/nQMucad8qCDwxxy0dZhXBYhevdW
XCSRxt4WBsMzWb3nVHL3NrOmUyUUCPpmdkytf455AZtBW5vAYrNs9HMVxCxUE0BL
yJhA27jdGnHGCt3uJUP/GUm5BOwDDWS6jNqVLhU1iSaN6HuB1+PCI8trAMnXxxtp
+hAKfQ7Creb1sIC+vT5Cs9NAFXYaV0xtykrf6K1LUfe3epDAPkLdvsEXE7OuaYUd
k3n/DG9iHI+X5K1Nkh2j3RZZBLuTBOg9GtRQi+0VwxrjPvMNZZiLCaz9vO54EZT7
BYJHEMj8iXGVEooZqxQGmUvXRn3HQQ/Bx5rhcEDBKValPXC301p4Tasv7ezyM8nZ
lQ5HU0W+D8nycvrOuWudC+6mqNoZSqieXl073igbcjmKGp9RtJCbi/Mc1TKU26gn
xouFiI+584TnZhZOE+KzB82GrtelHDHn45JjjGJASROtZLqHbtyMLNGesa+KqNst
AtVpWRRWF/cv2D60OQBFKHPEw5xEe4jge5bYMYEUcgcj/NG1j+ZV1s3zYkIpfZje
P7ezsDlEKYCjLzK49pl7dK5T0IITmPsM5IVSvyj1M7tN4bxIWxFnWxk9Wbrzoc02
g0mz7eml17Kl8UBKbX9uEORGxg7mmFe8OX39q4+aZ5FJOxAxVrFto5GmgUcrvu0I
n8S9zTEGEfmNjILYWHYQayalTTGNjLd2yxApNgAN4v/zzQkJoCMH4j0acnmLvcA1
bHEB/jrpdlYgKaO5jBC4pJ2ptRlrjAOh4dWHo/e16XjumYPk2GOCGsoFKaBZXAfJ
SN28dLrkeqzBjRwvvbNgkXEXFL3ONTDVKE2XF2Dx0cpKnTgmptCDYnmS5/5w3qyW
EDsJ7dq25dcouQCeTYFG6wO18uK1yBNhAORu6IQnBvaIoDGwic2XDg3e84KD0C5D
/5FqLcLIsdDLtnOAkhmakv91D6ogvLf+vqtjTTnmRqbf3ovK8bJNikCIXh9luCau
AeXDISQi446pDK5uVBIou5YaTkLmpOQskTuJfciJwTCweblzGOm8JCEdBKM3I36G
LySEAAzbeno9JHTTu+RW/j1Dml5j7SBGHuL6QGV+6Kn1/8jvfokCqqw3RgiOpfjD
DN6WBYwG8eY2hTxtSnSjT8T222rAqIrzhqXRM1TteSGiHg1TmLjnTDZWXhL1wcE5
u1/l7Z7upYodyC2oE9jJSop6AHaPJ3w1bSTBAsgVWKMC5yzd1F2Xtmh2DTDHmFIh
mtMgpUw2phYFlUDirn4NrwlHmiTI7G5C3HsLluVooUBbtDL9Dny2hB5zoEWi+QCN
l10ppd9qSFkU0Epy9w7VLKPty/zR/rSFxQ6Q6YwNbvzNZEsSzZUt7WdEIAEIpfn+
fDOERKHBECLwYs4iQnYvqEoTKS6owh3sKVSvxBku42R/Uvg+vqxSswYO7A6hGCZg
BBu5GpoFlk58Nj9J9v9L0C+u8tw3sxmBy+2RN448A5VX26SHc3BimoCPiY1qeCNk
KPF76BswCnddqE4HalCWKztxrfwUK4nPECdeYPPxsuyqlDMn0Nwm1QIH8aa/scR7
3k1XCIm+YBJMZcKspvDQqyPow55BIZ9qiOAH0+XHmg5/u3TqaT/8Pec/50loalwO
00PK8wP5dLE9iJ2/TFQsCvlAVV1FZujbt2L8+fkZHAfrjgaueelKj9bPHZzYAFlW
1oAxhbvbUV2WP9dzHvbE1EAJtR/eaNZ6/w/rnDLXoiNr0+wSTcDf4L2HGHt7eoI9
qR7XX5PrO52Tyf+YKwCPbukayoPkprvkdOOyGqf9QAZtrhOUkk8/F4jvZ3/qd47j
N6ZYiyVhxdlq0SxtPruCkL42uPCx0zQffeiXyHN88cUgQYA0cB2E6Y9ujjNMARn5
pWabgy+3kP+c3x1Z6BnGluFMC8kCP55CNhe2d9fpVabhZqAuDjCQTv3HutTYIfJz
WW52cP2i04rFwvpMTYD65TxBD2ZKrIOiunHmGv+SzvSIaR9HTdiUpBCeVbthd7PU
0n4kqH2JXZnHRwlKj/CikkYltmbgtI1RjTqTclr1P5Ny8YjwBIgOgPsoAhpmgh30
RBjpbbfmzjB44vkfIM53o6rU2oe5ka/eZWqnbJZcmDywoAbaWuZLtg17PscbUfUI
f3Gqz/8UKc1w0TtmGr3d3mtVBHdW5aNuW58KNs9v0P1IECexbWrP0OGok7xJD1uX
3gWujwibv7YUTcRMSE4308JiaoD+K1r73RE2Pu0KQBPrLPglz3vveO7ShomJ6VdS
gnX890TQvv0oZLr3HW7s8h/gXMEWsQm8epxqQco4tLv+WpNWJ5WWpP6kg2hQvuGH
os1nQX0GoswZHSuEeiIVJ4oj2z3R3Ydk9N82mTH7zZdiVl2mO3eyFwdECLGmtvQn
ckd886Sv9y7njRQLjcwbnMOw1Mq0VbfVwL4yRsKcJD0ho3LCyydBX5VyBnzagJh/
KbhPF6HRLJ0xwxrtnM2XvO57DV3lwMHEBZS+8J5LPqID2eO+ezyPUpHqJZhVzZr9
eiV/lqq+7tobOIywjIuQV1Tvjpx+m66QGESOpbzv17n0y4lfQFgiy9Pl7UrnnK3l
aemQofQLdlhM0FnZDXLI3g5rAaphnfSV9vBEv6D+e8pv5rwFMtVI0wbpln3AmOrS
eGidenHrGecKY9Ue0FW5CJB5FjId3LXAUtGQ9Oc4VxDckqNXGIq/qNcJARx3b6vL
3weoUri9xG2XIYXfV2CPZZkBuhFm0JbOUB04spIB9Ho58/XibOZ0c6XkSgIBqrmI
dAD2kcIubTyRdzeM9JSvrou4z0oKGl7qLYT4GsBACfR45OeVksBO0vjw2JMJ+87h
1BwCJrd2GWj0Ops+lyEkwM9U8BnH6+fXbn1FFqK3PcfRtrSSzxpEPG7M6PrPpM3q
jyooRLNBCi8UBt8xgIcKIK20MIXt9ajUGJUZc8bfqMezfJLLXkUbodrhfWN4oC2X
P8eojI71A2ITlW8FJjDFmaJyaHCLVVu3YnAGvnGsDJHBiWyaDCwU+wBzJQtU0g0T
t8DQNI0/lr5gYf9rI0t8eWaS3lIyMzy/Nt9GlGB2KqSxQJ6NvXn7qNgMBU1DhZKT
lXZv9gTjKvq6LlYwSnzsq+a8fYEXe5Hm1i/VpDM1XkZcTRq44zhmQAvScA7nuQLE
2jR5u4WKzGDyPCxVmWQypgVajJcdZnAV5PRdtUy5W97I7gyNyUQ4d+XUVA0ebJwR
u29cI7x9M+E4kutK5StV0O38mWqUMsy4VU/bdHh+lR4h6q2PGnZjaq241CnZHDhN
TREwHzhOROo3OycXA60wwzBtBlm8xM6QzUrXfcmxPOETLN45/jIV9QxBgGHyxmKm
0A6HqoYE45utcvBSfU2bb/0JBz7Tv21WnvFhpKHLIFCmdlAboLGn4pHEpQQc6puO
aPIjUGgT9PSbm1qxxfgUc/gWcQ11t6uDbC4Ules3tduHSoUfYPWldS+DsizAvWVh
V1OBkU7fguYhtlTftI4XqLncOAxw+ohTcWaRFIF845hoHoep9dUyjT567Wx1pxry
OXEFh+irp3PNS8iZTfAO9iccISoCIuGoW796FBsZ8snjSIKtPEDK1QggJ3oCIKkD
VsdmPWNrqMDjHHr9Kizw9ElOv0DDcQbqMo5N+h6DZDqVf2/G+vE3xwA30Z39u4kA
BeOTXoO4rgxJNnZry1EKPNhUlyYzywwprpfso6z6ld5y1RDmYs+nTR8XYhKztVFd
pI2r554n0iK8Mu5T5iUxLQPHxoUxGSfHdX86EFR2BvM+L1ak212OJqzsuI2QZTaT
1W4KeSDmXpA5+NEGU5f11uODpLb3atxOL7qnP/oT2NWYil/wN/QjqNhrEsUwBDtP
Rm3WE4rYsy6XQETKvZVD/urR+fOSiBTsalOVeihiTFRJ3zkse5wwi05tgG3GShPw
1vYcqwMsGxuZIrItZ+4YLYf006ne3E2aBdbsUQJvawa2pku4I5kiSOgaEKNuEWYN
0nokhO5cJalTzKzdKp1HJPTx/MEtDS6RE02Tv/oXzZ6S8I9tCfvVkOr1htKKFjab
ZNmbta15ttVwbvK5h6aU+Gla7ZEBHD7R466LvuxmjK6OGcQiX9rzsf4+b2o73+QM
qsyqVh2sGQ7PQQ7o+8e+qb7lyMfJogFjIRbigS//7hP3596PhgDfd4ortagQz2vX
XKHrWq8e5wn9UChU/f6NQfnNV/5X4c7W5qR98tOwkCaaNQ6HEn0YOcm1RbR2i2aq
WZ4Z+G2nW/RiWmYhjJfJ5ykx4WSCyCLaaEiVgz7ZeuiI1y2APyQZYY0hnyHu81GX
+C4LcrIUFdo0IdKgDMeThmG3Ie3nYxqF0FGulPm5NkvBW1Ea6vq3bEB/EEzMCzTr
1EJ6nViZVRJ0iNa3uxm3WpNlLzf6MIBuMHawG1kpswopuiJnidrBP424aAGy/6np
LW0nj9zX+tbiD178xhyhYaPTAJ1OtmGyXFbCAKJEsXbgPWIehaJviiGlhfygs/p1
u8u/qXnOh8ZyMGtOx3mL2SB89pwGaexxstKBZqV4XPIl9B8Or3ODSBWIDDOXaTQo
E7nJyVZdd7hMua40DM2veMyt9vLv+5rkOxNHddG8iFX3d+f+/cTyYiuv7jZJDIiM
Csg4y8aFIVGz26NC5AnCvI1zAB8hC4roLeOZuaHcPMgJA0N4VUqRQXmvlAhPalqP
t1ldwVcAlSt1s7/IT8cnvqYXX44E1nkIr4xEbPRZxY/vrVkTSi+F4r1T+Kj53SdB
iDF3y8z89G1wT8+S3uVFp/2XbHJmJvmN+th+0pQrvIVOKLniQyJkRTslq2ABJcml
jcFM0xhsBqeLr7UbKCsh2yJbfsZG6qTvHoZOJ/Lao6xiDP7OSelBfHr2l0jJdyjO
KRi7Qcol/6eIjKdXskQ8kcuax6+f5oiChgCFim9QkK9pljdJ7dSdbof9pHF/nvJU
a7e6gcI8ppvhXM+CoO9s/QKpGUtCCsNWLnk2BnS0fUhzm5A9nxD2c4hQji4fqj/M
NbguD/5ZwDixyRUn+dnmVKxBZxdX5052rRUQWxfx0ypcR+HFchuF+7pMsPjPemjp
m4a8qjXBX0VcSuX2A1vBM7F/wTjXhsx3TKzEzh9ghcryY1VB8zxu8yLnu4JMvqLg
qexV73p+tOAXjK94ka3UDe1vQj3VdWQhXPzIojU0tPRzZlWc/dU8j2ngd/Oswtf0
OSXSL82RyNW7tIb6ca2OukWKs3CYr5KmScCpMjHRr24FgL2yKP2lJsOI65ycj86f
7nu1uiSFVQz00NswdGoT7HAdr1PubJ3wUAoPATeI4LCQE6uEu0GRAvrOstE4ipca
E/JVMvvXngQyF2yVmyMPVWLUN1lALJy49PEZCrXOpsC51y7HrkKUo2u1AIT+vJhx
AWLe2K3Xv7dZMortutvug5rOkB5hNdmhow7v/0oxgZj/2Hd7YhZ41fYTkVtjxzEY
Bso7cZ3tsYbjSwIzpFk4LP1MHRpb2hjXXPxatCaqnyNf2XamV4aAVEoUCjpcyhdM
sXZTE8sOWma05RFJodfZSAP7s25P9dEeUKQ8e44Kz0lhWBRr5nxJG40MUAiLUu42
H5kXbtqvsyeGFG9jvv3Lb//0TcrT086ODUGqzkZdTDNGh9pIxuE91usKTo5Q5vbU
AUbyy0W7Mg9o5M1ZL2MqGIDM0mVUQtXL9hKpbiRieARqJWGIl4NQKW1aadKDEOMs
dYZ9xlOaw3j2Fppc1maOFazOf+cq4QUdQxobirdYGcL78wi9zFOExo63j9yQol2O
eu3zcWTzCylCdM/hNJrzeV11KJQG/v6erhIdf6Ki2u7i8V9+x4XkneQINMa7b3JW
/Hr+159ROtRCTxcwXaQXk1Dz85yQfDuZZdfcG8kIKNT+1FaHxxsMRO0AUsX9PUUh
uYkNHsoYSzk3pTXD7oyHRo0dI2RcXI3BeJ4g/ZRwaywxkkxXkm/o2vuK+eNfWutl
tfVTWHEblQJCwb0EiAkEewzvBKuY3nro5VqlnJ2Zop4BXxUqAtgZDggqadGkIUzC
zAP5lCfWyL44Ne8JGy9D2QHoQcYL2nYXaCPtdo3YMNhGhafBKDp7mbA4nR1FVlT+
qh2yDzS2ctT/TXhbQOs909QEN/BlGvVffv9yhhQcYT8OpFJeNG8ZNZCMI4S8GThL
kM1k7bJm5C9l7/SOAoh1b6qx4SNj0/nxdA/l9zoBC/HTUhk/T31/0unJhjYkvNwE
B0XpkQCRuPvDfFCpZX/K51TQ/buSIEGthPtjwC75oZivHq6klyV0wJAgRQ0VtWsa
ExKXmtotWsEvM8ESY/S/Dwo6Ov9y0/n8SrDMTAYmqkC+mGOaz6n2Mnsw4LlEiRMf
KXBWqFBYYKhOeFk/KmHE3VCRLWcWrNO8XLKkkWRT8IvDdqr82/02sEPE/G0Un1uJ
FqHaWMG4skUeDcgorBO+bPkSMJ+QPpS0htp8W1EeCrDL4hwZnZ1FwaELZ986NGxw
x4wwaZUDGxQrjRVElcGwG4EasYIAvOb8AZ9ull5IrQSL/AWy3Jd0mHqihN6SJMY9
f+Qkgb7L7rEAzf/PhkwrY/ACngW3CSCwj6xY3qdnA3I9i610qfLf35IalXV7gvQ4
C06m7GcPLRAwIFI4ZKy1VB6k+JOwP3Qpo7E1k+ZyCMySyzQGljRmi82CMBVwIUj3
c5/YyLnOLCyKC7SHK19miiKcsXxFeCLnGN3La3zirltdwx6eH3AKA8m3aJ7SJ0JJ
HKd/frqnEr3DQrXwxiVCFdI/gInwmlL6q+TdWvKmXkbNG+cY2Mdn9dIu0AJx4rZh
dI2TbV3VD8kZsp9E8zHbEgFSe0x50T/w0CrEgPCtMaULWa+FjPDaByn3WdCzTkva
0K8YFo5mKTO9UhnI1q1Qc7ZBstZfMa1IMGYW0aq0p6SOKeri3aDcPb5YXkESEcdj
ZsPTGdvS+TgGeTqrdraf3i+X4Eotx2lTrnmxNnFNjKWWrUXVnI38NZMehsnxBaaZ
ez4hTsJv/puPrJqWF/ZvAd/hI1iFBdCb5l7oN3eDAB9+UmLlMVNy0ituXzvDCCr+
k3cHlQtcwKC6au7KNzpJRFPvuexzOC/bJdmiJWBdGrC15MobQBpYGVoLh60bHlQx
cttUf8ivVVS9FFPIxvg5zbVLJ3g/FswnO9FC+LSEGTk5PFrgrhqvmLpJXyTcDgPm
+kXl7R4OQTEgnbA6wHcy14auMocO0UfpY6wFh6EbygDLnXv3xGViZhnuMEU1T94y
/tz4q08RHZzONy0SxXU3CrUie4yrQ9SD/nmCoFVDqrAEZAW2p+wLdE2wGW4WNvY0
6cROpB3go63rEczmsGgWvNTOSUmaYRbuM5/sDRCA2OSkDbCWfjQ3VChEnPZU2fpN
yW/DftKm/+MlGQWenLMTJ6VMGZj3lRAPzy6/K13udSeSXjGUjEms+8u5PIGiAZHZ
MKUXOcOiogVi+EG1gTqSeuBfGJ8lyAyGGpKmbOgvZ2emujV32IpfVid67xkJzDD5
dZW8+xnlIbxqrMEO9seQ7jqQuSgpdkLFT1iM/tgQxxIcAaJODR6GohmGurcMTAYN
x+yEe+IgfKZOzLO5hmEmbck6Is3sjAipLDjI+PEMtMoYsdTVKpu//BhyMigcnyHU
JkSIdJ+0a0JWOTuiTJvXdIEv7r9Va7xaAFbov//YYwbuSSBQ1IvcXz+EgzaNwamH
PPyn80+DgIIek/mmB63ltRk3CH4nC5+s00j+IMmTPiAwL2FeCLA5+ZiszsDyFDx5
p2Lwe4H/01NT8dIyv/EnR/Ob9ZWIjGTBqk6jjiyRlZEp+paIzAahSYg5FhpXgxkh
qHziwFuaYh+rmjZl6hHHkO0tzFoau3Y4FYc+yNT9Q77qPiKDLBNnLM+dYYYVYtJh
PuleYe1UaxduYC3v1S5CuU2enbxmfv13sdwcE0gBGgYen5OcgfiZaU7ANB9q8auE
lGIZN+rNj6Wti8HtcF7Ns5RXk3fTzeb4vBStTzirw3hczqX9pZyo4mCrkL7A0HR9
0Rrzaje3vkqo0cRowDZAvd0vkgUouLVbK0OczHzVecCFEOIJKKn6XF4O0qBY7hHO
GTb4MAgBZVrI4V/6nCa8+xyZvicFIsom9XCskTCj5MN5sZDu/A5JIFxji1m08JQr
kklc38HnGgJ/wvyMD5LRfIQN7vKpmUZcz+bBQcCnoWLE5PT+yOs/T9R5Z7fy4jNj
kClEXEXAIG/73ZTL8xKJLib/8JuF5VCNtNpQginBDN6FrL0ltjPkBXSXDMGg2hhc
ELS/JttrOawXg17DV2guyIgBXVETlxw7FOPFN8HfmcGq95ll+WwhZjX4ZUTu1zpr
WhhnIapVW+cNZ+bWCPROu4OWnk2eK7Ba5ojHho6Sea7JUOd2oQiU9cro412bO6Dl
PeQcNEQizexhIieyYi6PUQDeUKSb4XZhRmMsoHdr0mndh7NPcs5K7H9ywkUiQnoD
SEsWC0U7/wQ+2iFR5zj9t8qqcyU0y7EEC+8imxSpMEtNjIkq5tsPhrc1iWi+AAFe
Xfnx7+83nVOKWC+jzLlOvAex6S9MlfYtN4Oqp96d1PMqbrN8nS39Mf5lIysVd9w9
3BCEfeFKCcbYc1W9sdR+oq7IUV5zyzMAQtCCBQb0QaV5yFTS2WiPr3Bu5uwmqFvm
b9f+3wbav8v4F1c00Jf1o5wr2wyW+QCUz67Lz2dHNRGTu5PfatGNvCgoXuv2CRbJ
SRZjKsyQjLS/QOfdvgmdif+fPRuNis3+/b56R4EYJZWQr47EtKO4PF7ETP1Rt/an
YfZXU7QB/GxH/le1USk1PVnFTs37TNhn+o813SdaXqgqjdAPzdii60rqH188xaQ0
bsJ1pgLkfbzm+hIK/2QPOotDI8Mrm9IftdvOEKdKzXtzSTyJgsfZYWzi2XEUPFvV
W333iXVxlq8zox61f07YWPy1+BYZwzlp9/2ODLzwB2DWjyV8S0bPmUtnrrRN9H+N
4MjMcs2XmVxrMM1wFyP6eO1pt8HlqHN2vuRE5NUlLiMEuBjjPmmxG3vBQytJ0Rj+
OnZHBUcGoviCU8EeKdNa9ef+tDcINWvDs/pWhM3BSO9O3jQS1tcFTKB7crprECwC
1OQiHKTSsnVxNA6NQ3gnScdNdnIWsoAg6fqGDHPnU7sI1mEND/GYJj3eG2cyVy7d
NcizHyBBgNyoTELStKgtCRqiWE6Ikw5y8kJd9uyFB38ouKZY8w3jsB0MLUUN0Otm
eZ7BVFv08xnoRlwmud+6DVN0DY3HrHKqOwWEl+OjUvPosKRKQGQtQCsln+qXwT1j
OXY+ko/cB7pwGSwmEQ3KlAx08Xb2uEM9244klj6ig5E3t2fVVppoHq7wUQgCtXAa
rYLrgUR9LSgjoSW5bpm6KQdzrytO5qWFDpy6C8PT+fH8go6UOyJFMsnP8tExFHYu
QbJBQHIMyE3zgmR3aO8BFh69sh9Y7Up/6BSTjuYk31hwVAj0VN6Jx83E/J2RdE39
V+kgV3oV85sKXnB+cCxzefY3jqPn4WPicHcHQViil5ataRzXgmtorkvB2qhw63UM
I8HVxw/thHXd4ric5BpKzCw34h/gsmFK/z+XOuyZ4O7hWFXrkkPkJYF7pOoezQRH
gBcBtq5DUxp4Id9kjWnBD+VC9fnPXN/gtA380pdWugt1uu9hqcud25bJg6uYL6s1
m4EbsEs6GcY05f79qsCu8AGo+r7I3yM4XEcQmqCySlLWL6lk9cRiz+/bBR9Mb34p
mmWxROxxs3pAhjfZLXj3kAE/tIw5x7rrhJMdTAizh9wG4OU9HKfhEzHdNBQwrN6l
rsR8zVfaQzROJnh/+0g3lUNyHVWQffP0Jd4pOxoA20xtdbbzex477ZcfM3l1FCqM
yRJr9CmoV7ETtnoUZnHbz3KR083P9R1mSo8z5VRDRZn/h4H0xf1zFdO7SDvHk/Oh
2UlGB0dR3Bq6i0tyxWi/uNwy6UNZXbmbeQtYwgCY9Y2cTfA1RhNJrtZlqFHKUPZZ
sGV4G2+6ig/rYGzRk/GW3liHSXBoZlx83rJQJ9X3fnnofih0cHGY4D1zd4TPKczT
pPKCfnPUgjgAfSjaJa6Kt0P5UmcmRUMFFKVL742y5l4EjFQveG4IQpWg1XYLE1uO
4OfPdBIMc7/E6hjKDAguy4V7a5NxVO2k6qChjhkdDpxbXMV1IKYtwqWjBzpIDEZX
MAb6haYb5M8y+gCl3fZ2OfISJYaSDmYOqwo3uTk91hhPv14bx33VROCeZMq0aPKx
g+Vwc+uuQzpawvnRFXzh/S9ux3sWo/OONCyYOP+cdp/GCnUgcvPM4o0MUTecm6xY
DG8FrUvtoTu0I+Vt6MlEmsoh07YBbBtgupJJSGpQe5ufTjYOGmUSb4CIHXgLfIz/
D0iJIvro4m20r2xBw2OOK6bvlVku3BJyoRhMiRo1jWDgojr5rnG+bnqBwoLDbpzb
lVRXVqmClqbNXKT5XN2ewuarW938FxmetrqTsWx/DL+D0k3UjLZB5tbDeeUGTELq
/eHnLGmkoUfY5Bg7gyzMVK5cRWerxAwD0LnLb9MTOH9mnuMNCIj3np6YtarSpgx/
VjKkOLXWi1+agUFNGHcL106xvfwMVyisQGVCXyDbZXSKzh5SPY3zNWqrxuPpCQDy
mab+wQUPmSBZkw88ca8GfeEdkv31o6p5wtgULoSMfBnWPnYa49+448NQ2/XpsR9+
QX1GfUOnbJ2y8njJqEwRKtWWPHe/oGhI6RxuQZo5MA5fxEh2o28DCsNWYhpsYc2y
Llkbz19zsjQ4hEkPGwl9ToN5gOt3O6OsAFP/ix7oru0zRZj3yW8QgA6kqzNZrXNR
1qfUa36CsTFr+XnbD1a6TgUtK/T7w5+VyrWGnsGlbPh27y+7RM5O4v2nITuTC745
wXjIvNKVc6mqF2tdJZmNLyvuno+AvnY/ztTk6Izzv2jL62gQFjYd5WZuCPqVvQWJ
LHJo/rYj65mg+nhwjgbBDTjlvXDzCLsKPQFP2YoZIvtJoi/SahZpmgXUlP75VuGf
o6KHHTSZaHNVUFc9yXUPhKXa0U8QiFXqzfV8qiXOMbTKbStJ43yYXEw4p3Z8ySiM
Ii5YzjRXZfpL0e7j8fejg1qHUHeKVv07G4G+XQvKAEmR8DVCo0sFRxmWIRpedSL2
6gM7NpVdVEorNhivHANzlmrSXYsPxIbcSIJixFgq0C2L945LwQpnzF+LCsZDA9Iy
99TTc0IS3vXfHhE8yKzRDmJGuZxAoceQ621CBodnxZ6ZdhnPVK2A+DpOM266syC4
HwrV+Mv/+vopV248wHubLVlzyS+dAeXzBBfqk/ABIieJzT9PMMjFwMmNV6Sfwa+5
UyRzxiYosuTybyiQ0I7mlnSYt7wTdfRfmKHx3Mlg0IU7DVE+o7Twav56NGDNCpb0
Jm6RUGXd8uxTxgT755yDrMQTIDKuKVsYfPRMk+kRxh9/qpWLJqNaNWas4O1Wshs1
dizW1MD+vyHh1GPj2eRpc/4LsOEj8JGY4NvgWmNkoTENkN5ljKZbtv1CPP+0mFuq
AO7woK3e3QZlzAF0GWsAmwA/FZwzF4Pk2xdJts/r3DJ64y1qPX0WnhBMqjrOBh4W
VYSb+onIDVbpwX02s7kIZYvPaxLS8TgBwn4PmQdBduv+jXwSRZZqMcjburVTmIGm
4c5YmNg17bXnOzhH59Ea7+mKEBcUW5g1a3P7Ytj9oWASkom/5h2FBSH5l5bwDaPR
doT4wWdjDNpUiRTcEzM46mlenT+ivc3H9EowYafxa+wQBarz36sXbHB1wFPdYAfC
m0mgh0ZAivNzlrnbDEvL7UsdjwDCnTa+eZ8KvDkbgRXmLJNAnu9UoFv5wEcLern1
JLkx5TqQTn+oOUgUS5xQIYWJX8b7DAMuMEJR3D7DKGWqGXqi4W/fh2cYyk/tc/5g
WexFvutEmf6o3Ps2ucArh8KIkoI1FelVIFoAZy/AaZvLVGXQJbwgxqS41lNA0t0K
b79cRrAB261RROVFJQPGl3MOTvjnLALo7nwC38S674gfJKXr+R/FMCJ+viG5fGmh
8QAFkkZI9DCOKyznOiufPNuF8oJoCc40Vgawf/FjerkV+xgw4Nn68/wCsEFctlTX
ya8kOqtvquyIv2xzO2lz8PeyTb4+5mbHSdLViLk1SGm7NIGlt3STPDTtkMYZJl+x
4GIormPJJTTvP/L5X9OqWBIg1TL+G4CvIiIQDJ7nyhufXHJZO4qH3pPV2hoWI7lj
nSfTAAYr14O4N7PGj4qR5BMYJG+YlTtupXCyHHrFUgVXwfHR0G7AnsDMLlOqDZbF
6p1uSha7gbnUBZqWa0Hh9tbHxyfESbOGVomPKhaLomYan445iXWx5gpAzUBpP/gT
A0eTcjpLUEwDXegwnFPwa8bOSLBGQ7CwZHe49aRXuS+Vgs7AeNSgj8ZxrVisW4g4
ndGRnEmPBCGY6Ngt1pWMUzN9T5ynaNN9oa/EEFvSkBtxuAnaoKCOcJD3qlHa40tG
KbA1ABFoTX2J3yEdROFYgb+tE5ruU5mzpTV2KnIWAW7RH5DUx0ymdhCiNRbhXuYj
0xN3daSJjopO3pyKuc+MvxMNg5aZ7JvU9I3Mlj6cINngZCo00hercNPLTEJy5e0S
unZTlzVZw66GOgOcE+TVHcZL5/lo7pQEnUtBJMiVsT7XyEtW86CNGbywzjCvtNhU
bFNoGT6MS91Tlbfgs+Qkt/+PasOmRUsNsrPXU3DdB5wi8czlDEzO2tR+alsobBzq
R4Gat+Ch/3DdWrM8gbmzIQ6Eh6skf7haQVq10mb81BsbyQBwKv9EMrIBANbcSOFB
aLZ4gw6FcX952ICkcIKKodimACGh8O+cGy+dRdFW2XBlxLmGi92V3nWMRt/X8DX2
4zuf25x4DPY/57iFN+3OxTcOLoz+WXl3MF3htw7St1KeKfP87Ied2JYLA0vlJmyY
eQRA7qI5Xo0DOC38R5mTuWTm5W9qfnP8oOJJD6RV/sDCQwHenbeelXQI4nibqPgp
pesbhMo9uLfhjV+mHgBJHWTY22JimOVLX+Gym+DvbsSsnSU5DFOzu0suQWynmpT2
oUAOLmKyuBYU3LbvkXmcPU2KLANIcvrwz3Vvy53fNzVimVPzNM3knV4LVG9WF47H
9+Lfuxogyml6qVFMOP5PXcimKKG8DXQE+/qbrR16RK4vpzwKy7nNODnmvudcEEeR
TM901+CYAxDS0F5rJ0kFxxYei4VR6HelKuR07XPXM6E0gVOIHVUZLIJbzNTwSfTL
o6DZLp+p76ZhNccMMcX62oMuWDRI2EcXirCs166ZevTJgco9kon+Qj5K9UzrOpBk
hrJ8ocvdIKFTxDN2MWt4mVszwtPXOjPrB5Y4JY+H9qSSnsxWqjtX7l2cFpYs9MKa
uLI1svfL/wTIzn8cB8iGVqJUabUaGDUIqRlnTrTt0dc6+atu+LFOr93n1t9bLECn
VxHxqBoipxvQbHnKLP2P534KSlEEKPG0Ygks6pdpG+SYfSuxFqJsy04hefCMoUvw
XIogdlelyt32io/TRysSlyQL5xplxyff6wb3LndhmcnDR+Hdm3Kdm4zzuygz8ZcX
niVb1hTzqPoc3AmIPOwQjPFVBnOEGuiOz1Ic0biGRwt6hR95oer1g92ez71JN2Md
RV9aemHdRBKn5l9OCm+u/fmPPNol/lH/yfsWyVEsrcZOPysmPqPlEJOFs3p+WTOi
MhowHKZI5mUM6vSw0YLcqkBqtS6O5EmKk/75bA82U9yPLhCQaFZx6EV0cImaUBvO
xCiRMRFzGbSFNK8ZzYcatHO1tK+Iy+oesfbp2UIetlFbrXnoae6x7NrLCXbG8Zrz
ZCpjawYDVF6G2pe/Yu/ORTxSl2UCZ/hynWt7+6T/NCapjta5EuQgm66faGVMZkqj
5K9lAYO5hDMnsCJi7GPN/rSLnVlDewxOSVq/nKtYHk6C+/l6a+0X2QSNk3WOIuKu
kwVS0iETv2c17sFaNyQtDoeJxr7giqmadKqE64DtjB57HdDQOIjd8FCfLvgErTl7
FWO9sMg+JU09GD4UCbMt4hXDj56ZCohdB4i/7XATNm1o+/3XtZPxNOfjv7DrjWRl
mO1fZI1T59hcVx4qh7JLjPhb/SUj5wMqErs/hhfc9p7fAaig0Ia1xtJSSqvqZ1rG
UKn/3X8tjqN9sW0v4Gueb5psEORcCROt9mugEWKKU5XF6GVFN6wkCZm9QSTp/JjV
cRoTP4mBrJTLyg8eYiPDYFt5dDg/9vd9PHeaWqxWtAEnd8hvYWRkXR9PZup0HslM
pgOv1xHGdmehhps7zTxdDvaegDBoofh7IId3lp/I+NXCQKMMuhu0o3BDTNmiKnNO
p7I0WyOz8RMyks6Bw820Z3UcYm4D1VGrteUMHRkhCxaiyNvQaDANMCGNfP8lSrBI
XY1fGP4u6/HcnUpe+5nfjeKjdHwBocKTYnkOIAoenMoXGpVXFiRxJE8CYWpNNZHc
vB51Wx3Y4a0uiWCz2km4ZzlM2egD4AM+nOILOivt5h39483oyAMv/cFEE1IhDHkb
MhaoiLS1zv1AFffYYxv6J5KD/2NV5WC1zCE3vojRbttbiop3r6EVEucF6vepeL9Y
y2foAe3CfEISimgW9c/rEcyb5RmAfQPG8TueR4/TRY6LR9h+VJM3MIn1TZgxvU5N
tjNKFebzmB41fo2JJb2Yz6geerffmqtfYOLsexAB+WslEdadX1yuqG0CA129R7zT
u36q/QvFGHtwjPrPHDRyjX6KhGmmwy6ciA+EO9PyFB5hRsta/eG8mbWLaOsQ+2uG
Eqxn8bfBM6qX+Wt+80ECZgGyCkq0ZdUg79DEb9nbTsVvIaXOGtgkFu20Fw+J6E+x
8Dy26kUiHUPD55CsvdTAWpffZIoELyYODJrVKqQOl7qMuGblmhTrZVm7p0MAxFA3
zqPEAKVI29GJhE4aYrG+pfkc32vfHpoG6wR7Yxmh2eVDBYFGenPdAQmkjU6HQtdS
6gHcivK80cx/hBrkonTIQVrbH5pvKCUseMNFt+zOG05PMpzVm0K5J15KT3Sdq506
MRIZNkA6CvJHMRlFS9eApSO5v+1KX1URgaJjn38E1ajIJpiF9wSvwOC79fYgwbUN
0DxJZwrgInHm3XXn2MbzddHOe1P2f975wUmFoo78JGGX97ULYuD3ZLo1Zwh1q/6V
igxMTUdRbq8UJ5Cmy4+RR1y2N37FUpaDP4CRkgBaay8045rgPG0Fp2sh2ubHxKuf
HVC1O6Z5Hy+VQtvteAN/PkXiEUeU/OuDack4hD/ZgnbMW2aqt0Pq1cZ9d1qPfEpa
3LwhANUfuqLrfQxy7t6/6dXyHoiqlSnsmLQAWkRvaBkS5o5iK+QJ1EauBDMGLBh/
oo853iFfBHRe5R5EbPJnrG/Jas3GaCKp/KZLlcglUzUAZXRXmvjxEmnYiAT7yxD9
aKcgiLUsc86jhHvGny7wdAcq35gVLY/8CRJ845N5iG5EiiOp+k7+Imm3RFCS6G0F
eIG4K2BPsYWGDNvPtsxE3MRzFC7D+GmqQ4IgImKRYB/FWB62T6aRwIUVzZt++AQU
sJ5IKKQkne+63/VqZYkuoDr3dnHWUcSOI0cCGluKhr2tuRzuusYOOd7ZwpICDl/D
c8fKLdGPfbEeeGBxo3IbJYrP+Wjf9gyM0w4ODDemG0y/+swfoiw5rD7G7kxl/SYY
EKyZPnEY+rHYdhXlya+qEOOHZCSJopG0YMEQpa3DgdLmxEj7s/8XfwacJ0MxAg/G
6F2NQCOhj68XveslV+cfN5j7LhrQevhOzju+TFNuo7ikkgQZ2TkxdQAPkJU52VsX
GoZ1AEAoU3+H20z2buKpVzHnlDdJayyBiVv8L5wI/AM/r+11WQFDi/A4pO8OgpBc
bcvWCzjHq9oJILy6gWiGFZGEyoJd5onMDSmrQwG4CZ89Y31XxFLLjqxx5j8fIsY/
DN1brUht+RqLjTlSSeTfC5d3p6a2D1nA7U1fc4QD+NGuPp3IxdWdHkbKFJg78t8b
wapzDk7HVtmrjPBPrEMEnDIUaYJLPTnulZxl92HPNx4fCn4WmgyRSN+33ono3LCU
pI+4VsHxvTqH8AnXnEGmssBVkXr4G3HzxeAHpVwtQhTFw3yCgd+RZrU2R8nVo/e0
UOmyxFqt16O9PdhY4IuYHofq73cX/DHzDPDWPuHJ2DUsQxirGHyg+ONH45qskivy
gju1uF1L/+LGlSpn3gBbAxHRzVwf86rTET6UgIXgZYmoTxoAbGJBxr0tiaSWIQj0
EsEfpCOpeE4Neww5//i3z0b09CclUPsfec0K6xuR21J2qDXiuORrCnIWhojUeFYk
tlvYHGyyZzBNz18eOTiBtrM0nQ9n0O33cnS8MSmMDzd6gXpg+0N1E2h/sJ3zJsbO
wZjITRCOVCVpCtre7N82JCJgQP5PrNiqATZgU2epGWJQNea6gu9iPE8Gyz7C1+66
+jzqZCAVXuJw4ZWdGA6UJt7HHfjvnlleZuWvkNVHoPqdhrdiMs3Xjgj9HKMWB9WI
tI4Q2DOB/KHqiiC0bFmlRGmiHKA5Xycf1goappFFh3R4vWXCt6PSW4xeIiYUSL5t
alINIY/TyKQYHpGARdpGWhRomJU/476ZQdvcVqO64N/l2QyXjYW4UuB6IYUbAfBp
ZlZxls5i0brpXIi0ViUVpsg/5x9+XGBLS25PxAhF/vri8PxCzchSToyUH6UVZmXE
wNhr6RQiZXQqHNkHZ3WZizIWWCNYIoxfAHMd6vRgWmKnRDxZTxjoKZqDVB4ANaVd
MIrGYcM/AYZE5FPJz8r5oaXbT7eChuKXJs1bDC2190ILsNg36ux74a4Wsceotf8l
t3xWd2pB8Xv0P4Fq6JgK1yoTdmngZxXI712Im/biIJ2aJ7ZmiJ3ueRAt29Yz8xOf
pYgfhzXviPZUgmnqwFedjXvB/qGPd0PE3/s7VkjNOlN2HoDdHkKsyNRd8AYKA0Kq
qj590DezjcMCDWEdqIuClHdrkL1WcbqdKUaswmIXmbu/Us72aodTzdt+pxT+SCj1
D+Ra+Vtn/JUrXGe79lqdEK/pN+1q1LovwMP26CMw94ki5IRARAVWPGz9sFkiiao7
yGWV1wMc8oFgEtqkt8zOBTQP+NSzx5KmtwTGjpE9Ycj9vMFxAvNF3OfQJPbYngcV
I2eainXZLg9y/WcmRxFK1HaBRZ3PC6+lJRYmHsywzpg7jpQCOJMY9uUXxQCDYabq
+YK7/YGXSinfWijUfSMTz3oufYJXt+QMOG5GRk64py1lQZDWDDVNDNdYb9wjTNAI
AwdlO15CFo3ZM0QYWkXqf8Z/7qyzN9vwTs9mA+LsllAtaoTqVeO9Q67VD98scIYB
4ySbynJ9A/YCvgFkqPuqVYHvanEBxxUCbNwqIqsIepxStu4J+C8D5z+EgXGPMHSX
Q+g55aOwCFJOkgOzu12R1tQ9+DRcBDI2DeYA66rX8/YUV39tHeXjaiCKbBG74nIq
IXFYViFiCQPACNjTSiiFo4xpDU6gyNDbeb1lMZc5Z5FY3k4pAs7A9fZlaMz8OhjM
vrm42Mso/uhvbj7rNS+xve1pDrX4LaLS51uetUS/D6kpB85kdtqpC96x2NSrCiEJ
KYWnKIwHbQNvjvs3ubgUTcXtLavV9Hnz3/NUGWSL/LR++zfHWpcFgdB+zoFzw/Wo
nKvndia5i+Hf7A15kYVNUBYtlXvGLmYLrP88waIKmkFZlS+Nhxfi7wHEIJyBr2jF
kem4VgvHKcJQXCzX+gKmiu9kiGZ5aJHhdbBLoOH2PNEjA5j2vlPIZDWt+riyJoqh
gWJyghXO5RM3BMKH3VS7o0NAdQIVDdsEg9JQrV7eelpkpOFEY2HBElfuxr6t1w8J
Sht9ZI7kr1q/AaRrY/HOWkV0hYh2ZlxZ/HwVo/MkTbeGmBwcfkDMSlOlDUxkIU2r
JpYwK///7AmXbXt2NHXxndv7uN1Ch+S5bUEl029ML4C5xB7Vv/zkAe3jH8HXtQIw
mif2ZyIaB0YygVZFE2a2LKLax5o3Tzp43hUYkWti0Ty4LVWn4nRsrI1d70c46rzU
THvELIFVhX9tqvIvXCCGH4huaxsYJMhxowulyGA5II4svyTloMHeBsc45FGl5oy4
KqJWNA0BnW188LuauJpYzqoB2obwHMJO6Jce8nlfeVOBEbeRGYqxjL9yZOabh/Jf
i64AEvdFBbxoqoH6k3xiNWZaII6VdBqmf+gi/LJkV3tt/HHWUof4Qj7SJk6V0/u8
wOtkjOlnBR+oHxyVbayiBoYMG+XcAIFs4/wD56hTVTMtGhnShLJE9mbbAVxFUgjX
/5ewlL7preGY5MZ7nuLzDiTwFOZPpUOanfrP5Ke/+hIkkk8mfOIjE9z+KMUD5m6b
TgMNgqzbHgGozLo/C0ELdh/zRLXXmEORZAPG7uUys27OUJZDo/AL8hloEGqW2Zx6
++TtR/AXoJoitXJrgf4/IhsEuvg/d+TWWNeQfpNfiOZPOfkNIUyIMvo35d3v0MpJ
jrtF7ZZj15Kep0MT8E6PeSq/JkmHbY/k4BS3oTaYDxjEe60siVrnwDweJ32ZWCk+
3dACLAgBW/8nxK9IxpAPp9/8rJ2ACCRgEIZyLrJuwVJNmx0b3l0haUnPb0QEixqf
7AsU3jbUDhzMelw0zxiGBBD24sFVK1c9N/L6DWEQ7dCJiJulbJDKN0Gyim7HTuts
AUtdtTn4ZbNZzwi/mVZsWOzGCjTvQOx4oHg1+DY/X17O0l5OZgOc2qvDYdnQHDhR
9m5pNprDz2vr0/dqNNQfFxAj/MLwV00VjOWwAFQ8IJIcVhF1jf7udrf3aassNB1V
byPZ0wUfI83GtP1egaUfwmrgUtKwv174GAnprRQ43i61uioWUIsBLUhGBzQiqLbw
m+RmNqk7zz6/YJK6byVP6KWdYrJRZ0nmXLf0UwPQcX6I9VY8raAUFs6mJfmPxts2
jVoqpim7JU6pSXkYmaE0NBDNZGdHWGR9VBGonFRMjr9F4+QQ/rhWK09IeNAoulJq
YKgUUhKG96415g9vJ4236bVdSUT65UxftAcih7EKhun0eWApvExkRA+YjeiEl/yQ
IRJiWhQO4w0b0R6oU9WvpNC4aKOhHbs3TtkrYmcgiqurOqIKO/buJq8+pxfF57uB
MH2yAS73e9JMMFmrZcmqaKKc2DTHjOWfPIIBpM04k58+JvGHSkx3DwDpa0Cav2y5
I6wsVbbPH5qyh6qf4TTDI8IHKoHUyYzXosUZ3kqM3+S4Bv0BnvhFqW4CnaPsMy0h
i2HYmMzRwdBPP9EAVgxSucxktYsjNRHSdQqYUdO8J256JjvifgLSgOdKzxQYWhgk
GbvHlVRd1scO+FR1QqptkZjMPzWJp+edU8/J1TGwJKYj6V4tSIrltPwrRotmdvji
8JAZkqASMeMMiaMsCeCXmM/y4P9d8cUMpwLEP5OnX56hEe0/EhRxQz6qvkgZY6Nz
frW0G/7Z1ObJN9Vda5xkywxINdq51lyKTP4jhj3ansW4NutJEFS2nY12k7c4HQDf
b5naqxLFMup2bUqHYJ4Kew/Reh6T50hyq7sh7bpo3BVJVJ9elc/wCKexPR51NZef
etUx/n9pqwuKg6TNEi2ShrIkLoF8nwYhnnruzotbiad4azrkEFxA3Vc1SJ6Pq+49
EZKGP8kRdUkg9bsKC220psfbiS4jVonRapmNQRWMF161AJgoLQ93NV2I32xhYJ8F
w1xVmVT5Ku+co5vaghUfW8UknJwdHLwlW/SenWvI70G5Hy487QyBZ1koe6FzF7ch
HCjiyQIXP3ulDq00jOGXsbOJjrMsDlwAEtk8c9X85AcgBfBDO6nubVTFsuxcAV5w
ALT3Zu0/BmedO4uX4BzZ1AmK3j0o2vUuswzT2m0ILV4TCFWTVAQyKT2iclxy6Jzd
YBttzl24VBnngbbpxzOZjkqwgLVGjhin5AWOt0M0yYdr1JYfe4R6IdiY+5aiHmn5
+CFOOJf/t4D4ID/o0F+oWa1pntuealKElsa8gLDFSr1m8Pgamvm/E0bjrHw2Vp7P
zKl5DR81wOJwTx0iFrXAdpfo4T5qG8bpDXEDg17SxUGcDoovjW2crDDcXTK+jitR
ed/+C3TX5xn/ZcUS2DeDc0MiExIVd1buGOB2EP843yUv7A0VXwe4t3rHD9BFUIpk
H0a3/eEyPPWcNoWWKt3LZJOZYE6cnoMSY55EssT+9BCnN/V7Av23Fuwv0TbPB5ex
9VZ9BeogvlYD4TVzdZxlpFEIhhW8cww+WkHf5vM1Wa5YcszF6JRKavDxdHq2UNry
w9/cuNPBKZ8Ik5pMhZcxpWo7ecEkpDsUyTaCM7Hy+h+/icloqW1mZgAJidPuU629
/sZRcYDLtFRrygasycUltBvAGdRysXKRRP47mzCStM6lSAN0EPKuRNTi1XrHWscW
gXX4ut1TkURPLyMgpvJkpiWD8kcTeYMi3/BZlR5v6e02E9DhRuhgXdHlBAExb9lR
H9Vn3MPhRE3Wf9sNSEh/4h5FiHepoELC/zLDN9uLiEHm2yBwZIBBSivk7FFdYwzU
2oMx1Z6wNXPJ+h44EdBFwItx4pip5OHsQB3o+1XesyASvk8LbZspGJbWKPfH3s0X
mZzmWbepVmBxWrU+Urer0u4b42g6ny9nXWc89e0FM7knOv4VRM/QQb8DEAiUYtVF
A0kBdVf9X1uQ7xLjOpcdkJvwsgv83zCd/FbRsVBjoZQ2GE0TYi4LCTIRcLUuzwxH
AAuMt4jq4xA17B465KbRud/+unImKhF1enGGuqb6Qj3DiGym2Y8baE87FwJm/RAj
kPg6HfoSvxfMVRPVoAM9DKaVTkSonOsGRjPGoyHAvPyx6witvFJRlg7gprz8JRmC
iZkxQVUAdNgx6FiNEo/i88HG1Xu6ZKFQqYFgse1YxO3oJ3ZBslO26aoqXVkELa63
UqmK094zK5NPEwqPX9KzIxanKljhrlfy08rNcBpdgo8KnCh3L2inorBgf6YBTuvR
WVB6QECJ9ULBvnLfeRijhIH8oNVwAgfDdkFB7pYwVsQbPAuJ26D0/e5vU0VwZnAX
Sdayfu0dUbDXU2fYso+3w2HuCmeNidduK/IYM+q6J2BSEhGJyhQW8jp4lZ9bHLXm
9/FEsplQYZHK7Zjo5+Z0btns2elaI9u+XHzpgIWW2YjAk4oBGDKLIAF+cz8t6KkZ
k/ddfeCTBBCi+xyVl/Fq4wdMspd3gonsBmIcs0z9OhlpDgJ5liaA6yyz5WaBkRJX
WZStxzgHfe4cPqDr3reuOJGGodB6JvHELrWdUWHMn0K3jJBEqSz2TRVxypzdqy+E
+bZbeqT4ODBU47tAyg8cEEzSWvFDNn/kaR1iNiqwF3VbrRRp7bELQEuvTTSBp+g0
5984gejea5VTW6wxj12Oqjas0zAGDti9TzX9VAZYzLFlYl8WB0s094vwapQiFLKA
kF7A9S+uztOIUSvh2xXgegy8c239KfX+Mce/FSego3mJUkJhGxATu/NGl2bOo5to
thR2Uw7jtV0lmSHQRVK5lfY+KlodfeQUUTq3fMrJU9AIG89KdhZmf4HXsouH+yZu
jjJ4LHEzzD7TTfrruhh+wEAYsgsLGNuwONr9ldYLI/QMQ0N0uZEzTYM1gZxRVPTF
xMIOWJzyjLWwLgmlWpCIT+tQNriHMC06MYK9jKaaAsHeGF8llcw0alkiCsDum9qn
SwJWqC77SlMiniUtGWK+jvonPoU+aaNJBCTWnitRioZKEQL0ktx5pAvliZu4a2Rp
wITy6JdbICZQnSMDja9KRyGn8G635mFd2WaJ+Rbgqfj19cIZjdT0t05R1A47/Gui
iT6OHEJF9rjRh5QnYBVQZho7Z87zaM5XAaCkFDKUinltQdAQTwFKHTSJfSUUm1Nj
R+sRtuTg/+iigJDKHt20APs1fyu+sc3/s3elSEcUzhAlK7DXwXnMWATdEB3hxap8
Luuj6/FTe/X6/8DW7+JmyvXOG6aACpQj4PhouJKVI+YVqdTPqUJbvhDX9Wn9Oml3
QvAX52XTXWH9BxX9VMETfC1QDssf0AME2eoJg8yFvlL/B783uNTJXx7k+tvukjKk
lYvN/4G0O2YzMj6oFOCtriQIMJ/WV8kgGCZRYSgAwCZPu7kzudGXRYXiJuptO5QE
dClkiRmZY4CohSf7CJhH0QZkaVegAqIuVWWWIQ5bHB6Z8MeXgfa15deLIn7XFTiL
J1b3+jEW7IeEeiOeba0DZfNBHDfw29r0S8ERWZ/l1BzfutUg2KzhoXhDxlkhvmxZ
y+5qMu/MR11pAtdzHZS/L8txIhYGZSc028owdW/74yUGlRrWuluJP2cTSPIlYm/f
pwJdDTKHuXkxZYGYw3z3mUBSokNWI/x67UqLSPtnGBAXRY6Tse1csaGUAbsrN7Gc
2Zw3fBIAvKUIUqUkBmUaWmNDpkimVohCWAirDzbYGSnGo9JQfII+pBa3/ekd8aeJ
RnNezt0SQPu1rqvOwNS1F9V1Sel7Sap5JXB2/UOqSM2aLGfHvTMqll8ROqxDYMxa
g+YDy7n0R+qwxjXCYlYWsGqFl0lfp8HO//N95aSltBmwbXfjoZpx0IJ2LdpTkDYG
INFItBcvf0192YvlOrLut/nxABCEYxZvqFZaR3goKIj+um8qtLzbZF3E3a8Jp0xx
fBWplksZ+ukhWpdozXdAjOc3tlOh+/LdHwgC/PIWwM/AmnLDJzmW0PnvFa6dBiro
weJNYDMvAuyO8fD8mLXNLfaCiQXbWY6RuNbIaM5CsO0If+gVMTA0K2RqW87VyPhk
90mvakjb+z7AeN+fznoKAtX6Z6ar4qNP/gM/fX9qc3wuwKSqTmHDQooG/xHA05+g
dmZSm30bwAiz7nRxTtQD7eQzd07qKsJhKXS/gENpZPHYrnLfQgsuvUeiajEu32m7
QDg/ujwB6AGBMnbQYDw1IqqgLvJvAj/ZZGMF0tgsluM631y3IbtMsjmRREDjwVZ+
KiY7OsjVdKuLzKgd+ckmJGOAhvP78OkfBmdVnN4KX1fomZRXD9SP6yZYNuvvo3kD
Rm5hRT6Y7M2XANTX5xFVMMtumdKl5oSA04DBc+h4Ixag/B72kaUwFrrpETBj8BAg
lYNgBDSg2t4GQiw0WMpefmvr2ycrt8h39XVTcQ/OBv7wKxYd+pNrsvp3hjOqtETY
RFY5nUXZIBhQ6bHiNt+noMxoaPdqKX9uTk/ZwEzWnEb45f1pd/mRcvNZ69GZB1rK
1+KOQyXeNU3qPVwQiiEp9J0L3QIIyMhF+FeFI18vxt6/7bE3tm+yhuIODfBktPTf
mCXVvJQ+76x/0uSvnFPbYLKI+lcizqJupK+2CkREcVyJ+thhL7RVRPIKpt6UdWUN
Mtd1MqnPFDt5bDoOU0LURUiCcye3otpbrBSAvCeL++W6bU5dDsOJ/KGbWt8n5j6x
L7AuG8ihDoonep1tKL/sDTxNlh7F7khxRKr9jb1u3qYoXV2evGvNOo/ZYdsm31R6
VFy5WtrXippOgWiX6PKEgjriSp4OoLTIlgxe54bwpE4yAabj9DshOJewIFmxSRO1
OdcTl8ZD+SK3/GvIU3gC6uluVx7PeRuuIPyLMtJeaUErbpzisMTze+sjLM7SSGAb
fQT9oWDedWjkoaTMZ5ITE9eMa2+4tEZS+gpr5odGQHYq60HT1XfJsNKGyDWMsSKX
ekKJp7fovfU8aX1C/fDw/xooUntTsjekjnb/hMi1ubJLl3WN1Zzku8dW18C1y6ek
G7MHeiL+G6kThdF56wdIVqO62+upjI0RbiO1CZYgKIVDjbgzx+xmFG0WJUBrUlWv
KM7pxvAa44Ea5hDEWLDBdXQkqU54rg48vcrhqNRxiDyCNRP3LgyJmA217DqyWo4B
9xelWBcNKdIYL0R5N4E1ZdBsDo9Tr04Zc01XCC3xbju2KHt6fWhxQuEjOD7SLhJB
elwewPCM5kXR6Ipo51gd6JavPqYL7Lw3G1QpwRQS50Q5L9O7xdjfgcguz/a1uzdI
g3/w7QYUUZEW+XVnXDY8GBfaE6UPDkEihf/iUqenqmT9i5jMHssqD5+VNOi1yK82
khU/BFcZ36lz9NH8NRdqIl/EhwcipXLG2vNhYQ8u6I8ufQrhxtoTD408I1Qb9TCm
Pq8gXLaoeHtxHUmtcWSoZwgzM57+SobcPiJ4lDbfXOqw0RmwYWYj/JctcwJXsbbR
BkICtPNyQvPNS0CzsadbYj2w2+GCj02zlHot5q4FRNXsdGj/8Xc2XmH46DSMU0Ey
ZNO1qps7J3qnlFR5TnRaDaxDt+6lcfL6QEopM8GqpBsE8U/7XSticQQKWTXR/nqd
QTm9Z0AVXoVJL2iles3JodqQY1aMkOCZjY5t8CCYE7loKHCfhYlQSXcOd0Jv49vA
tFVUPtL9VNxS1U2FXE65VR4YKrcisVBY6kq2vVff5BipRM71QeHmYmokkxwFzXgS
L6T2tFc5NORARdymyqev2obMByOcmDEJvSgJPrNFDHuw7T1buM1SNdKP8KmidaQ2
8qUM3LQKNSsmFH3nYphzNDN+8VkhOZLfOOh5QfWhnNVy6nF7lT2TTiD8kcLAxv+p
+bPKnBnHR+3GeQRoKSrLILJdgTsTJx4pUPuhk0jtFXwCd/6HAQrsZHUBqVO5wmsD
uCd7PJQ36RKnv4O1XwEdz5WLF8um2SUV3l0Oajs19ymTNP/BuzxGMS49zXtCss6C
e3vzXs3YMDjPv1tJFqvimFz+AfqTLMk2o5Gl3BGbDQjVA4jRW9JczVvCtFZmDWQT
3SageJpadZt5BNvu9YYcCseuyi3q5KbgSXmr6wbcz4FBE66DaDdRUnTcIagJ8kVv
jLLGkv3ZRRpSPZFZqHiFseg6QF6rDvHuaIbRRzkCMGIMZ+Ut3JHzZj7CGpS4l8Bl
4iC6BJeSvGugt+dBa4wAReWYCZUBv6Y6oM7pIcry9vt3kaCG2nbpR+nusSSqXMT9
/+GgskVYRfN94JPqFGCgt8ATXIk2pw454BvEqrqwhcQRuyY0CnERip9fe8fDKadR
tEmr/gDd3+1kanTd/UaLIXLAmnmApb8lRQUkdbPq6YPyC5HTPN+MptB+QK32tCS5
tWGvWwzFrsP/2hNNf/742Or3XfuiSP5SeSWzp0fQ+Qcljb84ZcA0tUADUrSR2xa0
3tNohNI7nFYJfk+52aMTl+hZrTp9IfeSdoeLiBOH7pNRY25elhsKcKB5ItvQtoC/
hpEoi4Ck2FwNMTfl77KNQ2+S/nctM8/qxjg4tNwlBkR2VkVXobeEreCq0A+GFbj3
sPAYyWIrNiAgr0pPtnWvMztLJJyrh28PU/MS/vSQR125H9NFVuBidJ8UfvvozN9L
4XmgELS2SdETm2XLg2qbUuVVYNXOx8i0o3EiLY7LGJyg0Rrq0/94WvxLMJL43RyX
qAUN2COvSjm4jqLEYGmejs2dcujhvvuS73LYQf/Rnl5dCxzOQUcv5VNNznJRnADI
oM8CQmcCivc3cEgya0s6XPBTjilQ+I3FmHoT1D3lZLmyXTeYXFvNiPWmNlj7Lfyz
lPHc/rC5dIPeu3WuukAdG8nWva7ASF/khd645C7W6D8Hb5212eJawyixr7hhZO9/
bUdAQSIXmark5bGkrpIj1FjpqF8DvfZjHwFL72Ln1LrvQr8l2KSczNF2wIcNRDsR
eO8pp/i8T21pDmksfBXTbTpVbzndUmjAOS4g7kvmInyAeBcf/eYI+gP/bc1noytR
PQ+SEBzS5hIFJFbvH6CI30nFM56P0xhtfzibVxWXDHt2WN7z9gVmM9+GOZ37h8wM
vyEdC0tKX0hrHNfVZbZcEpS9nxE6B4kZaTdr5F4qG4xg2TC0YII26OiYVEOeMKse
nyZPCgE+MHLJEtp1t0ANxjGiL5QRkBSSisWA37VmUmZtjNHzJegra+31XBB9Qz5T
6NvoV36IAzB7SoL0JKd8BVMsrP51Gzq2UdETEbFGb1LPqXvLRvLGmdWxMl8+gM9e
a2W5PZrVtMCwaylvH3WBrJLR31MlrHLD/PPFp2dYB5bS4tmJhtk4pFGRhmg+mqlx
fT6qmx0j/72hqKawlGm8zK73sS4telDgJuZFm/dxS3VbUHIMbY+EMEBZfmz1QZeL
lskQeI10m1n8DmIip0Ih0aSiY8lOAiN64u5IjmFAuRvbqe3KpJoVI+ZptrWxavC5
3JS3vmmDktUtwF2w1cNspOTD6jQQU2BLyeBghjK/GoJSGFstXYm18b0NEokCb9xD
bPl5xeLicK1THzj73EIyEzlEGWT3wF3xRriU+CNdN8VVHaEbE8F2LJALLgd8JfD8
ZA7YRZ29H77N/mZftQCq8aA3g3tprKW7f+ChQS4tgmYE2j0NX3vqCTcLxyNZh2ly
3FiYMzPSfjcIRgcv9ru2IdmNQ1s0sL5x28W9GcXBlaufgpsGPzT3oJ5YGeB0QIsh
3wsebb/WnAWJ10MBTvE6vQDzgH5qDHXjWlmEwSMQGv126KdyeZDTLVI8RZ2WsrSe
m5+LUoigMKFjkM5/LH/zS5timnVzO/6Qf19tnADWVEMrvJGxIgwBiUZgNrn0yJp+
ZETH4TZpI33lJ7phmO7fDbJfD3cagh+AvwfH9bB1Wyc9st75DgPtSCat8R4lpmi0
sdNDBiVX+4yxFT/Pl3gd7BWiYjVLlZzYT96BW6ovsZwfRx3Ip9i/wD8P3Twt+C1V
cDsitsKT/eKJSYmtWbodcbf7nbOFlbNxyPiJ5SB691hwIWktMbCjjkFXQld3cXqr
nHHXc2PoX4bMcxh6VN/2WAEBrLaP8sPhhl+LcBNgsa2cTOCdCrIhxSpqbb7l8Vbb
Qpvk30KGmRtt3m7Ems+IMPchNJWcl45WkwT5mF/Ew8T7YUhA+ycksFMc86ULcFP0
Z/LjWZM0MYvc2XayB2jpUF+nk1UoBvkrFHHZaxlP1u8V5Dd7d6NbeYa5fRrKws+a
G1kdZQ+qrk9motSd7Jky/P75rtA7la9OsxjzgAy61brZYeItmonzyjLxRq5V4SH1
v47segvnHud6YHZWxPCMuTG9R2V8hWnRKW8wdFZsk3o9wfv9GT56MAGSiW/YVPNo
XRYoKGdsHS1EbiC5YS4Boof9+nRrN8hRNWB+TfJ8xaotdQQjmJH3X8lECKb117P+
45MZzIm6i86E2MBklhrk1OZ2p5qSYH9oMBrkrYesw0U70PxPJgw5rUoHw29RzadM
wT/PXrCksbMxO30CrWx7Huv68pdxMCd6fXKx9JtL3A6KI9sysfn2xFufA+IeOD4j
EUOu7Bo8S7nZnrwZkMeq2Mm5PLpOWtk+d24dvofUjY2vcomWhRXiYvjV9Zhbj7WF
4Zo/S4qZC7ZiG5A8eftQWvGOuQtCsA1omAHDkAJRu8dXQSE6UmIXNt6DWnwtf6Ut
EPraiMPcXud69ipvScjP6OHJ5DzM8HucqmQiJWbYmmuTVH6neP4rTO6YIs7WZ0KT
nrkwKp5XWmIJ0I0SaW3rYYak6ZDISeUpS3XFpGRwUv2K9k+g/fTviRPNCB5biosJ
+XCNcan7SL68QdGPB5UL82Eq9uCTmFdckm3h4jz8DugGudqOzz6IcDSzlekYStET
lAfwLHnA5tw9HCBKvO458HrGDp3FylQB3+uZRpyYwse0JsWlDx6MhzyRR3+8gk61
kptydWE4eSmAoe9inJizbl3X7APHbbPOCDGf4adns3LAPyIWlv8JCQ2u4TW5nCGD
F87qfa3lBB29pPwP6GpUdgBGMow4GSXHCmjQXAx/sgQp5tHYQPoVdHUK4FJhQXVp
RCyAev6MfK/cLsW3vztnm9+0skvKlVBw5siaMGi/kLoulr8x+EqMDaVhETKsrd1C
+Y1qFNNeHfO2n4sW2c6xxLAx1omkmWd8QerDMtWsI+94UroYpL1TLubGMyq1OPcR
ApmWE3m9vutuWbzyrATRZrGYiuVC0CIUefai/o2cMSvrW5eiRCkY6WQ0xmmKr4QX
QJccJdIEf+ZfsX44NNW8f2lq8JAf1nfaxfDlw5vX3L1KcyVucN1POUw4Bn1I963r
LwfcoIWkJrB8W9A1CY3ziv3X67Xeu/XRIreoY8ZdOw+qkq/PVqQTr/odRfndYsty
p7vnO2a34ybVomEAIQI8Oq97oC4jDnpGp2RpuMYq1tS95Ay4fkTtnX1Yu+QWrWIJ
pAf2srs7v2Bx6i1P/9bGbohus57wkiL5GPfed1bpCm+RD1NeFn1t/6wtIbVUFZ/c
ANuH6zqtKdhZOFl7Gnm9yyUOs0xgSZc0mzB09znDolv7x5wiyaOh5PE8YprGGdrM
+BJXeq4zwWLiaxkMJYPt/xbqdxOEWhalckQPicw2NNEdorKVHZap3vTXyIedLkIR
BRzQzAmUINUkJ5z5vFC5/ftnFCnTwCosxRhjp/uZEITZX1iZsMzDl2Qg/hlPctJn
YJ2zzK+szpbxgs5S4z+YSJ4Dd4wrpus/rRjilMRLZaMQ4ML2USC1EpQPUWTPAVmY
uWdLSxicoW0UqoTtgTZzXzkt+fkLmztAeCPUeYdaXEB+Vsy6sgvhwPdQMuvwfGmw
XJeF0gf8vy1FcBbsnrOJcMyoE+5FNeK11UJpH49fE2wRmouYcqGaDR3qS9AByV57
6/Bf0GHRJh5ZWjPQjLdUrV9FN3RrK7F892GOujLfYPJW0Mf2plfYOOMV6ijLVr6X
oTZG/ZvyuKLbO8aP3CGXmmwQaMHZTWEvE90UeKKEpraipTDZc2v2Vd0oDgQ8Ftkj
tzkVfuwPdc7muUdXuOeeOuOrj2ZPolnxIXA+5bK2a81jDMPUeT84aMSM0QmFhZu7
LcpChsHM1uRUvmSRxvegE4xFRgZAnzd7SCC7qiSday1WEDrdOLqdx/MxWl/WB4Zw
cQf2pTSvbKMyzt8tcK6XhHJ5V32pLFAqEISMchc5rM5U4fT793QrroHNq2u/fhn7
5ws9zbPwIOpAnvYu9Q+X1vV97vSAFsiHsdrlbQf2nHXOG8bFug+3TnUvuviSUPk1
jyaIyPkPxUdkEIKEDjnNPlAEreHR7eVtsrfM+/ZBEoysvxvJ62Xn49xYqc7isrWG
rvz/5BtMNKd8y2e6m79AXV7iA+JD4xezSHoAdxp/7hxumPpBHpvKDtddFHYhJTyo
ptCfPowvhLfy3tqRXuKYVUs+5Of2GWH7by6vJZGlSYXbVFDwntX3NYGLmIjVfnrG
DjgFAa4jS9+Me3WvMlmD8kCXL2fBOS3RmmwcffkSzDXX9CTlsU/D0THjnVxL9eqQ
Ze1d6ZKrxdjqmEIW7USfBF6YwJU3W0l8xpW7gMuggXmygirzzmHyk+6MlziDeuFB
LMniU/XouuO7qkGtgTyi3UnoZ+f6tHgPvJ5tj0fE0+ZHhUOSO+v2xQs+Wai+3BS6
Uh7xbsU/04O/9qj39+sNdTfSpAJrSlF0RuD7ACNtAYzoZY4LRT1FOLpy3lCRzO7O
jzzlcpVOEy+LcQuy1SfCl6yv2tnfzBufXkhUorqyhDB5cmQ8v8WpRlez8oX0JjdS
vbTIhx5wIud3K3y0SuFGudhsV9NWtS1ySUbq9R77QoT1kecraVo8sUH19hqDZnxM
1JzpR70jlilbKmhRVUrcKJ5TOmrih/8PbX3flvJdhPA9hEg6QYFuSAZNeaR9b/CK
Xb74q81+XM7tKWueU4IXXkGDLXd078sNL7gg1y3hMsDooXKPSFxQM6NMoCSXjSmT
RfnFQ2R5un7jOq/y9N03keD1xYc0EkMM0MJwIlscgoiDwGVsfhcLAxY2uEjUk98F
SPit+sVY1HWRhBgJ5L8FTPQ8P2d4aEMZ7NDbqu/GtW60V9GarkhJfdAvfC30g/M0
3xcykZjufxGvKl4wpH/SGuPjnubiOj1uVsKcUoIkTNoRurEhC6FiWR8+Y/D4vbP+
QoFldOI2tNhvKPwlO+pauXALmoPSnuDa+5D2sMrZ5pyQwraHqbNBbEr6eXoc6XSn
zpIENmat37wNtCViwbueXyBEPBXdMwN9X5r3xOw4tRTXYuRzmdYo0LVVe511oqDK
V7Z2rWOkVfmKwkFDz6J7I+aoEygWw2uXB3Z7RpF+nTkdcWIhUKPU7VGIRz2au2Ap
PSIE1JauVOzmNjGM/mJj7b0wQXW2Nrak5fdEhPg1YBq2ySLgapDBEYAkjJatk/H4
TWm/sK7bX3SJGdOzwxOKpkPt6lfMAvdRLVLchPpzAkMhBTaWHEG6fYvPq+eoceBl
r1D2bfFmehm0Tn5rNdg1gpisKxQb/jDyDZusA0TFjsoD07dA02mRzCnSwqo2Ra5T
l7aEkqeHzvhDF/fzXC/5eykSH2dsxYhlqzDaGmmyFHy9qS0aDp5QqPkA3Gl/y52a
VaBgQzqmFD+hzY9e/7Q6iI0r3ytl0yVHP8diFCHjgKaH+hxe6EhDVJ/+lo+cjeM5
ZnlqebF4nU9+/SUTTxDgQQ2KrdbgFAqgc3xE5jCZpCbI1GPsJEgB+rD2HqqCLjME
ljMYddzL0bQsDWNspeOMVS2ooRLMtnv3Y87V11pKoD1JyKENqPXjwm9hRl6LE7h/
nauwJx+0DSBfVxQtd9ns35ppRpk2Ey4SFjyNAUizQelWO1kEIN0qkvL9XJpM3gSt
aJWoBIKea9EH1WR552XjueMMW2Y7+ZG98TQ5KtpXDrsATPzVebXaJGwxGeO/0IqM
/KGlSAHgtXhoJT5gh1Nq0WZgyOrE3L6wS6Qs1RE4Rr65+HKPPDA2kUYO2oExZb6E
CmzFLC0rKIUj7PybAIb1pU8HewUwkkctZNWgK74gXcQGhv7TZ9+y+cGmKi8IdG6W
RORMFnXTgeG5sumGL6ejrBHYzCSmHKW1pLYB3ykDIdg46hucGbxb1zNJScpzqdfY
A9ba/GS9bBd1mA1AlHzC9ByPPxj/2yITRHAEAIe0afYxRV691pCNOGz2QaRHHWMz
TN9eKd/QS96LP69+rKU/8O23wkwDjfwXhVb8jO8Q5LMp5HaqsMWFZFBoFAK2b9mR
UMjhqvKHl9hY5hGfWwv9A7zKolSJuC9BLYgodkA+MdKeKTmz2fSfLGvKPpz5vQpO
45l8S5WuIof9SMHfGksOnerROqOR+rSXC/TwDG0Hr/tPxyg73O6p7UlHRmR8CEEl
KjkRa5l46PWOQxQybQ+ikqI1iTAFKXK4sLX3gImwrLutsRgOezq0LynUo6Bkz2Qn
HGQkZdx4DGKpnCwDVZv1d9NlGIwgweou/BLioObhxYH2mRLdPBYPCyjqoAtP2iuY
7hqlkDVFQpI/CbCsKYQJDGBbJDVo6lX0/hZKFrF+2Hqpuknw8qhKpM+ZAQV+ylBg
8BemBlu7SgwsUslxiz+4MWXtymqQz6FD7nIGjD1tGBCvjNhSrXZrwdpOqMe7zmiK
3ORLRbeXKduHlP2oBaCh7xCJ3qZ4WjSDkh/FNoudUFOFWNBtPUbLDMyE4rkyTcds
Cz1dTXrFHbT2B+GKMu1znvu2bz12XPeXWMj5tEc8OzT2grkxRppuW+8YBHoO8Ukc
PypT/lR1GHa+HQPHc3rZv3urpHQuhS/hh0Jb7oz+MCVa0jDRqf2VNtYnxB9YNNw6
GG25/b9FnDzYvLKJnX7Ak9N3aH4GbS6eBCO2ecAIDBhDtrLNr/7M6V5/NhPlrose
9v/yHUfTSr3oFE+VvV4drA7cXr8fEnx/iPK2roDG9Um7+sAbXo/T5s1VbfxtoVSy
F4sgo+yjgzeTKrvR78SYIZ4QY5CfvnDimihlZogpQY2A/SXRiHaCbD1X6Qk4yjwB
Thbwz/4dArYd18rELCrp48f1/NosyEr8WrIm/9VoXhC/O9bVpycjFNj9dB8Xo+ni
o3tI3zMatM0DgWkWpcrMsAkh8LvN9njcC7eepDso3eVuOcMwUimeLyq6/cDx+ONX
Oih3gbo3DyWmVe0j8hZ933qmmcCGt/rRVuqaGf7nAEcu1nAFJldkekt5dUF7gt+P
TbhgX6UpKLofaQ/A3DVm48VQXahsS405sIPaPQ/hdOfxD8Nh/+10AcrEikynTi0m
tmTNKxVLyIeYTL3vqUKekgEvnQX/ZLkzhDnkX7KgCGU0d/3H7fIrH4ix38ueHl6W
tk27YV9NDOCkzIIF51jYWKmMTwU0pAm2svH+ZsHwUTFMppJsrRf2GCy7KLYAtrqb
6wehtlwJfM72oH7+yltlcWGUwrHVYWJTR+L33vp7rP3XKmwpCtDdXrl+hbOiyKfH
y5K+/IfvbCVOjIHMiioslp//hX9oDciq5ohZlpRIcrnLEHFSkZQfkLuVSzAKbpZS
mtJgm4a0KFEi7z8cB0zVzrlKgY7aHsFl5xvp8KbJcj7xZccp3Ff43w1pWnpiKsoN
0mFJyWcoUurZtX8B4kfRHCWbWvpMGIfqwisgjLncvG+Ai3pQdiwQ81leoOBDi4x9
oUPAzSQuAbctepAuq81dJsw5VuHwbOEn+0tNz77iEIPA5eUl0xUxXEzPLL1TraAO
UCpi/rj51igRiOTDBg9HnPIBFoWsyb6St774Coo5VAE5uaWg/AEn9yrVBXyKpfW5
liNPHv5JzLDXrJ2L85gsfcotdL3OuFXEaacnObciswLQW8gaHqDXGCUpbPYfOmrQ
/xWI8LiTunM+jRCGikZLXmjjEf5ktTQtxknCB2WuZ/hAE0aaBqVe685i1/ry8z0m
0mWiHckRH8bt+lFYQ35j/spdx2E+nyMW+IHWFcGR8gi0jkDbEdxvDrGVW7mLrI2i
Rr/KINCKmYgcYYSormO7ftxwrC7WaNxd8bKD0enVqLaQcYrcnPDHs+NuafNoHZtt
lUwQK8WAHtE0Xhv4AkI1phK+zJ9TQEVE8YpazUPXYpOw3WDuvpYtOhXld0GII9E0
T9znLBWRkhKneh3KDAMY+FvvsO5B5AvLrg2tz6C8cJH8UFXzKxq7EH7QCETUoFQL
tbY6cYuOYfYypgt3YtKZeQprglzI9CCOwyxi1YUibSptzKHplYCSClEjD3674ldA
LpDtfqzkPJ7+LTr8vAPsVb+CO5AMabDbhPccPk58MV/kz3ZGW32TSujP2X3bSJ3J
lKo+SNzyCLD7EcRPNZHHxQBqi5/0cc3SYswkDXLQ7Q3fEGn7EtWomVCEeQRmxfT3
tGNtnvVUzgsrB7BahDcgnUOPJvgxBz3AdDoVeO23RRc1GqDiJ6s3A1j/KJzUNJvk
bzmZoYCXNxekI8xl8U29J/KX9jYzEwX85DZ6MWCR/5SY2pSSGha3BzH8qWv8iAj7
ycpxQJPFWkK2m0wvTD9CIDR/BUE8lIBYGU7ln5aUEAACAxWDqEo/5xoNt4dwVDge
6AXSuYPDXvYVH8S3kU1HA9BWWr/rldYyN58ayuHByNAVhDSeM3e6iq4uYpwAkiBu
j/ocsTBaEt/XdYN6UAF8Y3rJUtcpfxvp00Omifo56Em2gHRKzkW5B1oJpb3jW4M/
0gn3dAALQqWE3jR6h3ODBECtlS9s9hmc4TVHkNGwnbwWImTBvuW1mDjSIloDgxpi
58Nw+gXN8Xq6NAWZsx1tFnIE1k+bdCweF0iOwM3E2AZNdvEGqQkjd7WvKgzlso5f
D/9g8lQrf35TSCXQkOf02pEFFQ26UcZvCTF0xWjt60mwgnp/dXiQdkvCpfqTezY5
+aSD1lHm+3EbEe6K3LfoZRAIUfNRTKOsOYliGxxPSkE9eWsBk+Mxgkxz0QUphhfN
FHQkVMXwaHU/XiOuTMi1G6A2yvgY8YZndj3TbdQOcY1Ofuc/avzbxEhMrxL0hzCs
3Pn4ensGn0zfZ9Jc2pJsG06lwHT4DciEXJhjB4c7XcUU9gsijKu6CtlIUxIy9YGm
O9NfghxF02E7Y3D5I/sVu9EgWFFrI3460XEET+Z7Ws171TGOOGf0Gk5UM+bDNHz0
P1ftiMu7o9Xj7wUIRfXRwpbQQ73wSuHpZr4spEySRM0nrw0PLaiqQ/DSWeV8HWsF
nEOdNvoIghm2qooDD4iX/39BbdkuZ6mcTRNMuyXwK9QlMyF23WmMksWfX6QDCQmX
5eizo/d9rQo4Bh0GJ8/1+c+Ma8+NAYI+m/Aw46P0u5HbKvWr9nJtmARGt2ai0yRT
NomXPCbEJdEyEoeNFhw4anX61CetO29armObPSDnq8c3cntQXcmleCMosiA6/4m4
UgX7bT5Q2tDuCVXpqrpXreXjXGXZNF8DH0CK3Ez71FNLktoVyxaFyDMiOypwnYCV
KtqzuNOFjOPcf66PJP2DkrV3kV178IccCgSPpdAsWHKPY0+T6+mHT8e6Ry3sd1rk
MltwqOJjG2Guy39FlDeuioNzgDmzTP+2jP5Rka8dtsfrZ7SNCLYrMrWbNI6CfeRr
HQrpIKLvGnAnyhTfBVs/ijBUUvp68O7xh3v0elGGWB4Xt1fa+1Fo4f0Qu0fPdNkp
rSO1KvWethjqVOBu6rxNTyOotl67+/Zm0OsMXNqt4Go6wcOz9RfT0unPKoSpgzKb
loHYbdKbJH2X23HCiflOv0doxXpG9JUHc4Ih1igxI1KUSbE9W8f15kkFMYaPAo0S
Ckb8i3fveJlWIIYQQ5+i5bc6fdkcP5mqpU65UfrCFP9+VJsMsjlafbHfLoovQDKL
4wWLIjzRWZG5o5cm/pTl1rOUpTHhJhah/Gcn6SYQXEHgVvA/EvSyBUqeuRTzT7Et
IoaQM+AuVCaBepidRvgVX+LPIPbjqbhq2pyYoT4cECLc4W/w3RcBOTmCIzFSOwu1
SEhZPFiC/mmj0f0UjAlY5bW0yoil4VueAPkHkHoq58Pap+8jNmxWhj0Jr3DRaLZL
/RXeoEp2hwYoDB7AvINa03kHMPsv38RO7E6ywyJS6cLSHPXOPPAOJ/MOpm4nldct
m9LtTAnDrSEP9AgBS0Az0Ynx2zTMeIu8cGwNIr6EAEz4KG8gbFEtaK79RJdOXBv3
1Jq3qktpR0DlvzyORNZC47jZFlE7Fu55IfrJLIGZnYMAE1z+k58l09NELAay65Bc
bZmXokAYVxeaSTUwmIRxsAScW/1vN1z7jDtOlw0tLtHgg1DTyQny5gGjl1Njhjx2
xzMHucXIgJ3Gx/9JEWHrqkMr75Cpbh9Cx+eFPlr1UUMrzbuISdGtuVvi7fKFM959
W/gvPFcTq2xeMDk3L249fuVhLfomoD48s3G+VAsaLS4zKgT0PeQTWxfKsa4CNgkU
8Fsp+G6mS517WQcaEvluH4M5Ym7dZk5u+zM5mt/y1SeOXM/imlG/++klpfbZzyjF
3yv3ZJuV16I7UNz/XtEA2DyQeoeWv4i16mZbdYs4otBX2euV/2fVaAbuaeVBZKBt
/IFswmcLgifmFwRrqUXD33YYSa6Odbb3noWRN9uQL5CeOuc7NYTX/jPepJKwYs+c
cw7/zOXAAqsWIceC7kLWyIpC9On2I24CAVPKnf0LNGKqCj7DT8KQ/Lkb4Q5Rejxl
yO7eyeehDwgmV8zu/LFiNsRSAbFWRj/xeuPf/re3NgF1Een0F8Y1fRacC8CX8Qso
SRNl8B2Up+vQFA2w44ANgKKwyt5/tJusMtx3RWiwIaWk75QyRF7lPCJ0+3vESDhd
/KuvABMwgm85aL5XAktLdzkS1X31167gnTeyTdoHhqr27EfzBTufKSj0FFYalXSh
It0dGBOf3mFUJuoO6lX1SDBd0qLCDvmnP8aGrRJBBbv3mUgof/EaIpBV0UG2biLe
pTX/lyUYAsL5jn0K6BsFyNiCjnNY0urbEHCfVHFGAPATmFriAjD/Sxst9yfVga2x
NO/U7PsWBk7VuvmjcYEG7jxzstIBFjAMJvqoD9/yhEOAzpkXLhxWb1P+1ml1BpEd
ko75kZ8KNlhYpl6GF/mG+u3ifdSnWrY9JjQ3MFZOWxKxpKoBPePmAmpnUi8kSKaE
822spsO+szl8JAamWM2GfLJ0ux5Fc+Z4E6Z5xFSE6G7Lw1Kn2nlRHQRPR5Z5vF+O
s7g2PmUVc8vCep9+KBHSNyCFB3Q97leL4EzK50vDk7QnGH5CMNUkFOwLOApef8Ab
iC7wxnbO3nbDJ3nqA5a6hm+Ewx8auUKg6BcGKv8tx/AYo/nW8WsOD5Pr4980ncFo
QlpfOBupDbv1AMNfXgbuRu3Bp2OmhVKQRxA0iT3dt1WXp5gG4pnzHI1A0u6l71US
L7OgAqCkGPyY1llOmDf8LQVyc7ePBlNq2/ukLAFzPXvzt+720JFfO0S3cAA1T1p4
1gptd3a4ZT5E857XaljUz85s9wLoZwQStNpF1Vigg2WwBz0018iX8DfDDSjzSb0J
3gbSiltKphXwnAyZJcNfrn+Bz83w6wtYQxxiVtzDGtk6Nr5pO14qmaoaA0ClZbYu
65My03zUEPvCh684j/qfwNmA2H1ejZGQ5OP0uWIdA3f8MUyC1PKtzN7hAiJqgdPX
XPDX1F/E36x7wLYj+Ah3OVmtODZ1+IE0XbG9krwZXzsslNr2sVmlEXR6xsHw/Gc8
OFwmA51VPq45d/CopFgmT63lxhOVqdfoxm9ax32mPDUWNcVvqp0yKqjH25Z+IgxO
wDMxNKqsFTeEx2NXEhUt5qdhKoa+hRJngz0cRB+nL2z6esAQERsIQHxa40ggPU+/
D64Ey4f/ZS28FFzwtdwgOPJ+v2cHiRF1e4P3N8lUpkRhVHqntpa3JoBvQHNOQBrX
QeXdpKZFUs+2X2adUyZ7dB1lIcuARocWZFy/sJKObSKw60i4uv0Zic37RX+Tsrvj
JRSVPSiLS1NHBuQgAb+5i333xfbqsJDQAE3/sRLf9Fg5tDraSm8tDoSQ+N+OQV8g
Wftx3K0RWjvj1byA8n73WWuf3pJ9CinB/iv3jmIW1fQeFxuXRNMNpGRka/60fyRW
AyMCEWHi0snE5NVLIxSCSLr3ZJtCBJd/76hVCZH/BKhZY6usxQNpN4zEZOPKkv2D
sEKiGqjFsfWhexjlrVyNyu27j/u9THOka+fRL4nMffp/pDxTnno/vCNQC8/syISe
dP3fQOyTwMqiF1WDR+gBKRpSBnNr0lhtnAl42b7iApMRtI/yjgJ7chytwebEDWIJ
w0RrH2vnj06Tc7rmGhIJoGM7aevH/pvzUDCLyCLL9azTPridMwb5mJiOhZqTyUo6
v6Vx8LF3+AGZLY3zWBhl8CYlnhpjWPzcSWGg4uRecsATEuCkoCReEQ0UgEHCqhe3
musWSJsRsIo1bZCBG1IkhezoBZh3PNUGoVL+M2yeXC1/Ci+ycL7TLDan8ApKqtH0
jvnpoyaMhNW1z/9zWwfwdD0+omzsaj/Y3ntw8wUE+b1ZQ4sObMieS/PstiPeBlLh
qdXEwAjyGOzO0jWzPOm3U805H/99jFdoueOZPBdXD9IwNBLuLUtzvmOeXEP9dAom
QPsmMTjW0nRQibwsMaYktbFwLD5ENYL0xSyx8pk25GyGpCKky8EGznpHNmUH8m8e
8uWTTf7GFVe1X5PR8iCE8vA7nplRWZojbuURr/ZdSa9O/VaU8TzXTpqnUl+okbnV
NpmYGueBWFROT9+DHD4TFJPNupWYx6uLxvL8bri4mqmnxXPO/bqYevJEenKZFluM
BhBhAcOFTSaNPB1m2Cge8Si62LyxyRNjYL57x97qbyr1TZZF46WsRewGS5Xf2Slu
k999mecs1q875iQeVbT5+ZAO/aui9k0k3UQZLfhckWA2S5AQBFHKpyM+ENaLwkmm
KO90UxFLjaVbu0M3Q9u2pIdfp0MAWicmibcZccVjNoqzTnIZggGKo6lT0hMbXk1D
3MQTu3XHtiyyXfk6UTR9cDcSIQMvpmE1f8cV41ejxQntB6z1xMPXfJhQzm+SxjtQ
KaCmhvy0P2mJv4rVtp0givnTG4p86AIF46ep1DdUvu2jgaGP3XceG3/JsfTQpwW9
4s9yQZcuBGXfovhxz7GRFm8SXUbdnENPI8bdqTqivVsw8ekvI4l/pCqAkfPCaQfS
P0Eq7sIyrSOam9n8+8mrNxb8A6oVngw9K1izx7aDVpgusi30xCqwtZr1HjlC4h5m
3SukGwhXrZLUdnFovyRYJDTDQ4WZBs1+Jip1Fn+dyzmy43IetqJy5P58pHJuJMO7
z0vkjHIc+vK9/lZ/xEhuu0dFlG80jUEMO1G6X2OkxtXjN8LwN/v3+BWlTT0Lfc9p
cv/tXCYOF0khwzI2THb3HS0eDK9+QN29gOUy0ak6rhFRDbS9xW4lwUPNwI2r9VKx
hjGeQKSk2F6FwiG041Sd5Cbmg+kXJDuQniNbKUR1Azq7Yl19PU+aI9RN5bdqlytt
3gpOjqWCmwpemWjF6k7Xc0xCl6nlhi0MYMPURxuyas1+SOzFXO6DRMc/Cy4hyjCR
qK4jS5NCQX5gpHGt9IhEyEWgZrN8N3BF30Ax2EzYZdtvR5gqaI5Qj70dxTP9+H6B
BEt0K2p38/GleBhg8hCRM0+71UrnX4DqJbW6q4R9L+x0NwB/t7or6rc8JfAz88vj
q00ObitaUpyTxCghgkI7d82rLHV+OaVaQOMoPkYc7ikvboXtdesFlKHEPR+CDkjh
HDUOHslwp4hMBjy/dmRBqOE3tALbjAwMiZSINdNGjj3pYCQrB6cdLKbllw/facH0
S34MNIZZkfmDfH5ULinpWzUHGx0axPN5/7kjKL4FRcP38L5hY58Q0nU0jKKT9OCP
mqotle/NvcF9FKfjxp9G21XWuHk1SU4Ptw+L4TE58kIEmEyM9Mu3r1PuJHAsMdvL
zQbEOL9z1IRGKU65VFMhK1bB2j0hwpxyk4UOrf/H3QQ/F6mEnnqP++z8/ziUTF/D
dHOM+OwAtRBGkxxpeg1VFYKx2yklCa0hF1uYHveVBto9twUAa3sS+ult9Woqmq77
fDKbM3smzm5hIOItY0GJ8AZ6Q4NxvDNPMYOMw/xb9cB31hwAruwLG9vkrYllbuRn
OgPccIDM1Lnuucyndjaezl+p9d7V5taxci+XJ9Bm6Sep3RLoaP+woDtLbWY+EXak
LSsuu+Q3ZD18/iYMqzHjrWyccPy5WbvbyvlLjwpmPzUvSYn9PPL+KfHQGDO03Rc9
6qc0HTRs8g9fcEQjzxDiMVKDeLPq33kh9PF/XOJswbNzk5vvBiYWu41PO3IQSgrr
W10UXuG/N1lBaO4C3XAlw8kNJnkMszkzowfNkmGqWyh3mmkRCXpC8GrKQ/CiP878
OlzkXDOEpTMX6Fbk0kO7F2RJADveAYtlr5TsF1GyrXZnsmgqFqebBXZAIndItfCZ
ajn1Npt6FBDB3q8ctN48+BG4TjKQMc24uedSOIAo54w+aDgg5Zk3UAkK5w+hYw47
nxFAEBl/+f+J+UqT60Vw6qKbezie7DmElfGvwJpr82h9EHK6eNt/oGvYvj/WxGlT
QPspEdnGLm8xm0XqToiXvtGyFOe3vAY+f9G9OzRcfP/a/zW2ql2r6sRTVH592UV5
Z0ftdXu1j4IGP9tel3hivbnfH6m4Iv+XDgvvTcyNRB508nTP7/jkXDQiIqQ9odXS
mMns64iToZnQHw8M7BC7TOikwCQ2y4GShf/khD2e6N7kAmyKuSTTrU0S3MFj6uKh
kUO1Y6SYf8I+5URlua/cXV7SVV6M3WQzwz4zzMNovdnmMg18YKmoXDQX5Nq+R5ES
iAo0VwmMtmP6H/Ztqelpi67JrXx1NrFNHTyeJ7H6BO0gWCRxg4DpfvRCWs3bOSO+
dbbOsfgUe5FaVGe2mIoKecXciIsb4YYvrWTWVYOQ89/dqBfPtk48gq8DcHQe7NoM
jM5YXqi1+PMOUwBCUTl8MmU9xOkfVSaz1ycUxkQT/7R57eDt6yJuI68oS2C03Oz/
PGYZQez7bjmUdQ8RObNGj+xDYt4JMzlKth5ZCCdnJAGwULhDoDNsQxCNsJdbKdJe
zEx2a0Bl9LKniq2sIHblV3PF/fypTdy62SHH023NAZ2kQlAX7zDHlULSum/smjDk
JHsgUJC8Kks4FMADhhgJhwzAhp5vluK/3ltGbn/EatO/PVX8ac+jCTXoh3YraDCb
srD/oAoMi/kipYG4ukm8ccn7D4p1fAVfoYADJQ64Vn+Gv+vuFOQVnn26uBFzWoSq
bU/G2FuQvpYYHfMjmEyToz8DLmdHW1jLq77dl16vZzBgOx3X54M5GqIe/geLD3Q/
0GW1osTL33b9i/szvaPf2QEZR1GxOSaWM7SBLFP3kp9MEslN9J5VubrkCKws3csM
OE/xIRnu4MAExkaJQAEjkM4UoN2DaQPqIroxWsiepARbbbqKYl/H+lUpHpCdRFcD
EU0ccfo/xJbULlL4DDIwfZA2rKaZ9BojcSXDiqrLhuuTUalA083oWnCj+HTIlYut
OdONJdyfjy0BNxhwQzW9vS27BMKn77DKIFB5SgCSZsfykikbWfMYXGqdDjNgXyAA
+5XSE0tZheke3YukQwhcaOjbcViGFGD5cHRCfmbFasBwSu9Ve7NQc3ov6zmeTv4g
LR4EOfWwdz368n91KWpqLhvJ06iBA1Dwia8eRtZM7g5mJkG/VUBnFXDSqyj7opbH
8glclZT5CEq1j6tmg6AMolMPCohv5mNoWX/fVNA2+6CKy8iGK9k76D5Qg4ijlX58
iOf+CEmy2oDruXvlE0psvtG8daUELW8I+K8Nr8WjV438yX2t934leOZA3VfnTQA9
bChGALqANLszldZMG0HbuVgM1h00y+Qk+9peWn+tdhRmcj9fT9rmDiwc/yVzNPkl
3ynZ8ygKxCY2RCYnPRIJ0qoIATXgZ9Z0e5TfoMmG9PLrOSihXMvBVHmRgA+TaTSb
5ZEVoocjd+NGJzNLiHdt31yv6QuORPcokT1D6cgLjyXaCWbQcRGH3gikC9Z7v60k
OpVmjaW7klHZc/VPg+NwtPo2KFc53hp01yIBkbvweHjjhsrtkBL/LG3shwNrH3u9
ah+GfX/Y+7ZlDhqBfxzUT53OvDARW6A2Alkf3PxDgTcqzhg1Pj1XFgi7RfhL+i3T
tyRrd2vdfq7bbesQA7SnENYrFEMbEdCViv4EVEoqD08I7H17DDiv01YMe4xNW1ZU
4TQZNfJ0cypdTxi1G7ercNWuFIzxbmpUoX5GywtVLpDFzoNaOor2zD9M8P7TSQff
BnzKzxC7hi7GE/nKV+ZM8e1+NpDiztci0IQ9Z837POkVyhh1ClWOsZ9evZxelp3l
CZbMW4fPYZFAH+jk4MlmUPDyJq9f9FHfwezdf1VuVxiMEtYazOb/sQL7x1jSkZJm
XZ1Xt2C/hAWvjFKzcIoaA4PHdblmLkoHdOOrwNyvcrr0vLV3nyG5EOZHg76gHNhJ
pb5ecACBEKk9/30/HADHVCed6tBT+rEOqs4qzignhANioJdG+Nqp1vqU4MJ2n+kc
Kb5vZAo8xMRzIB3805gAtnnaJ5B3k9CejPtUvrSYPnBb5izZYQXbDFakQa0LZA+1
MpVbKm7YHNMNiQFUrkDwwDij3hm8KfswgxAgmv96ryl4Z6ouNXiZXn4dDlls6IZk
cFc/OnlRdqPuRkJFHs/Z7x0TR86LBhihM7L2i95Hc6onN8y8HxR2+jETaR06dKbs
fw+3Pfaj8PB28LoQOgwGnwmtShOkq+aTrW4N/fx3G/nJ7+Pdlzuf3Csek/bKMgm9
1FZZABuAXUhQ57MNl8w1DqREzWnRKk6lMM9h1BqXf1ZFvysr68Ld9xiCDD+eVFEz
RjXUYxsZl5108ar1Ohmv97Au0xAPc57j9iovQFExGn922wPf97V2bcRNKo6nAgZd
LVN5UYGj5W0AUsl5g59ed2bAJha63yyR/PA9r1m3LT/Jr7XDmOlNnUoKFP+FLtUG
U4mykuo4f9wMQjMy29sue1qI7SOQM07yNUFC2lDsonhPGIAa67mId9KsQnvtQJGs
pHxSoZzUdVADVUDSQPAQEjJEbunMFV5QI7JROMOCsP4kn8VNCZu0Mb083d7m+SWU
E8JSBQkQLdwlwaDnl9vO7MoNa+a91PoN0fWb/txZNt1UE8Ol41wB6P0luE39BjuD
UVM53+lY7XHQZqqdgwnTHehnxFqdDDZgAjn8bjJolCDdzWr6x8BMqoDV7Xt97ND5
73MZhKxJWS/tI1Z5bSjMclx74j9IQ1G7YLKzFyLuR1UxMpuDqHtiPtku6W79enxu
1U50GwwWNdu2p49Tu54Ikhla7LyVqcd1btT+PytKRMHUnuVwHf4Y0hmtmOmldQFr
kVMgCdPtrtjuTZLaCKRO2Qi/Z1dVmZN20BKQo+UHLHVBy8EfMGgx+cTGDEdlGvzv
1ZTfac8cGfgpdNdQx74e2gVBKLA6qp0qlSbL+g2oZ5AnL4xXThmT6F+tIaVvx8F/
lBsjU7Doly83m5Jzj6Zy7HyyYM694uS8Kp4sCnNNHCEeB3h4pWb9Gir2UM7KX0aA
08XpCN5I3TffGiTINrpIFSHRbv8zmU/wHnh/yGne3R7qyy45VjzbWBirXwoyTgCE
Q+2/EsnZiWb5SSp8VNRIK7EJe9MTOHRo4eNxP8E6hS2keiB5mZ09wN1rhUEWJk6V
N8/IFQ+NdcDpp5j/8VQqyKrJ+CmjG5cWRQey5kQgdssjgrGFIxOH3SIg85I0YTTP
A+z3DNNSkH8cHZMIGBw3D+nLo+RXo9FDWefz28snQ/pXWFcbvzqohv0P6ZgX+di/
ySNW6E//EPpD4gWqkAIzcqi7W+O5LvjEKsgeA3VyO0GTdumNTKJpNyTu2+Iba+vX
2lsBGBhD4mVlwJy2qxVC6TFOH4pWAVB30hu+WLE/BBAV+8m7mCo6GXSnxXT47pMY
JmBDS5nkUbs5pNW4iJzqH8yEhFyz5H6kHFhntSTXyfZXt241NfcgtdkrNfZshrCS
zAk7Nh+xVs9vVmlWrHKYfxU086o3Nei53THG9OgNvG3N/HeMY31ThuRGD2N8KJVd
Xca2TBtR1BYsCcm1WvTJkNG4Fm18c9PwFEVwFvqWGw+4lctqVEwUqOx18Wf2Ka4N
1A2IBiqU1+FMw3zq6duXqOWk5ickX8CwAUSUaskoMJR1/TejtfXS8J9BzZQHDNdL
Plut3YShUgWgwLH67CWkKv4BJszZsl6p7zZYvIbo/TCwrnalcJO37GmNmyJSamR6
mgZL1hBHWPK5pGDqhN9RH7zUdJ3j2CK8KrDDB4lD3WBjq7OifhiFru5VCATOBGyV
6DHXzAUJQkIgjEl7HCcQ1PtYlt9irVAbH2NMb7RsVtGu2SmYZA8X44aoYB2S/8nW
8QUJGtZHZuUeKj74m1vJcLEiguqSRjHjN0hcfpRIF3gjVvEhldPywHEuOczvwInd
2SDdXSA4sOV5e47p/zy7Idax0sCksr4s8os1IqQAx2sVgCYlepzWxcsfpwK9ToSg
7IVLNw3BOTeBS64WsXZx/gCXDZQyCJaJX6pJIpwDUVk0CsuE3xZVTKLvkZjxM0al
opzZTRhhFVUEIht23SNGeGGIu2eEfLUIQncdjiGHYc6VJHw+mRWqLtyiEWEMI8EM
eY5+cRcl8s4tvHo8TyFopZsI6YZVbZbppzsl29oqLzKIOKj1bMwz5vmBh/cxtGqL
swAHo0mmyV+uP2NtPe0FHUe4206jzQHO8sCrFVWMzKs1GzlqrQpRD0gUDKCTPJv+
iMegwB4MMst70s3PAzuWeaO1oPJGNF0E2W5mItLI6Ccf/Xxx51bRKIivXnTpMpvW
rTGdZhijFHM/5vhO8jQhwN6Bq38RE5rGAFI5kx0xsMTvSeOpaQGNhlmRMjI18rpt
YWE5AfkhVMt11u6qFM6iV9F++ibV8aO8LhQ3DHX7TaHgIMm6bTnoXz1gTF/i/xtR
ntxFTwtJtiSIDhXpkA7mA7BYmsAb9PfN9brqvSaqGkfaZCGB4ElzJs0i8JNCCS5o
Xw4MnUk4dQC74bpo6eVN4AC/9i2QYQik3e9pIHHtOLsSdTplK50mbA9DLP3Cb3UO
SxlLUdWm0rNOIgh2yU2L3NErYqcYOO/6ic4t+qzIFRjI6/Qii3reIpFG3GhVfNXK
Pfxq1MCVC7Ou0TTv/vniQm9bDa6ai0LW4mki2ctppYGq9MZCNtDCkULmcehhrdpc
ZifbaNg27sMf35b/8QHhQh51V8GcSHj1/vBn5XlgavR+1X2Ba9s22QWsxClCHgi3
IH6/QFVsAMJTwtB0jFArIMiK8AUb+DcSaTYUK0QeU5+BUTmV3wRJF0UdgyhggDkE
fAzgQJD7DvZ9FcV+qwCXwDjEG0aQ/fL5UwYwfqYeJnqk1X4H1T3zuNuguc3WX/gv
RqvKsAqrKfXeD/8Uzy6M2Fz/jtUlLVr1xCj4Gz2W1U4wmq7NL3CEzXoZl2TbTS4J
h1jMegq4tT1kn91pAC3yF2igEWPx43TT9EDaN99L0JG/oI5POSjNBqheOAqU6QNy
G4gJkvLSiVU/r/KLo/x6mMLVcT0ka9twDkcVxoo02E/L0RcYxhC9PfovvwWqDNAS
qCa5sE/uHd4jbGKyorJDEfYWw0pWYm6Mv13laVDwfvH0AHJewx4Gx+mVdPoUHes1
3yPxw/WXoprAJ7ReXpwTw2Efox9EREi1zjq3d7cIPrKVSDC8G2PrO7Ntar9D0tEy
E1JjL0BvBqLjVo6w17v9eyw9V0B6Uz08wUFlbJEPfMOBLbT4DWrNrfAsb8FHLR0b
U0LtborjO78PEa0BZ82nm+Ee0x/GoEc2xwcjZ/OkzOnMne0RfdArMDtlAigh1wPy
IpnCyk4rUgL4iDtVsraLD6GsfIAWM7QVVgdj4MP95Nbu+RNzFHXzx6/MLNhudXKw
BWUYM/0+ftaSPtnbTVZe0ewhi+BVGR6zXF3y5/jSM4pK/K5zfDOnk4RGefAiG9Ev
pMAzSuTx720+iyvxuYLpyicBV77EIp8gBPdi+juveKxQsgEtKme7PD7R9wnDnCcX
WSaEeYU22bX1GS7CXxruVo6n9ZZNnMHQTlJPEuQX6qoJBU8UdIsbi0EaQeNhgroV
XF7a+ucOgEUwNiYmhY8zFyp0ab32BnvDEdm0MhoDGgW3mdoWwHq2FM9l15svKX7h
ZvWMoLJI19w9DmVr7RUERmiAt0DYasDoI6BSGNQF4kaWteCxBNCHyCsKFM83esZD
7/+AsNBh8SuLTh8Cz0tdt4F8p78P14B2TyXX9S/4BHRtE3KRCKvHDSddD3f4FmAC
oFard193q7WhP/jkazjBnBPEv4d2Pmc4MMP9PhjQBdbDKCOXSpMVERFk3PcvXNMT
g0Ca5QqOb1Mp23DJFXu+dOzbKwP40YH8p8Nh7tLq18Ps1XUn+D9Ob2qHpGWeES50
qkQlmGa2RO6/EYfchPHyvb4wTWgtBLEsgv7CkDyxhkKDi/mZr1AaShrqe3xZLOUA
2+3hRfuSKA/AWOfSnL+ilHYZSJGJGfuxfbgx2DCpS9V9dS7Qve3S/Fg+9KTkCfZ6
gAhNM7deO5XId0lBrVMafJdcRQPgM3mo8Pd30TksnwyESfn2BG1QRFH3kC8vgctF
QlDgB04QTvTpXweZ0FKM6M7314plLOXYzeLh5G4GPI8/NNOmMHRaDNt//DLTfBo3
pci0ldMFmcpqgsm1nUKmpzSCna5k/5ZYp7gpvc4SN/Yw2IIa5U1dS4WRh4Cw14Lb
yEITqvTyf5sg2Cc+uyPC7RVRegDSoue1x7p2eimSGY85p7q11XYPsrRW2LVy2Buz
jG1KsWs+actefu5Q0u6T9LAtIiKk7bx7EAJHcjeJZskRC7cLLjFggJTzlRKuEPPf
zfXUG9L3V3r+k65dJOkOCgBvOOCG3xuGEyuC3MT0jZ2ubPgs0F983Trg221nOgwO
BGWlK+whD20yLkFtmguxqCHmY2dBOjdD/fwp3SnLPvHkRPz1bUEhzNQrYZYuAg5s
n7+qcrD/JJXPQZS8PYpVYfOl0gvNiV9D1FdxqSzdVNShx3xUyDZrZjh6xugXqDFV
J5X0MhhkhcH8CMcet5vYTpjq8K3p1kqQiLeqD4NbuRWAEiWmTk3ia4N9Ol9T8KkC
YLuWR+1loBe2yRrsyOSfPJGNDC/Apg7BSgfjwCwVf8NQ0zbUx1X2IOUblDmFpiaW
jO1zSE5CdzDks6T5azak/39diTBP3/KHonD02OC/wTn6RzCZRMpB1lq5aaWE4tBp
PTk31+5viJcSquFlCq28cvp85M8DsMDzkBv8MYUvjwIQQYmUK1HflaYL4TNuwAvm
InTrahHyuKoyRv2+c3KJo0HOlJOwz+gZIH0OjzWa3SfJdRgT1mIWMe9w+nc4O6TO
McaKAwlo8019q4MnJDkQB4fYxgyBoUlvepAimJXe0mLZbMhqkr3jBBKxGL1eelQj
uJIhXwqAoHomiKZE7ejfzf4TKsdseV2LUGYNQndefIPrFjpFRKtRogrUNb5GYy8Y
h2fScyM1atFFwOJO51ZVzLMiOT+VwY62y2NdxyeIuXX3WjLOV/q46L6Ppmv/Idd7
X4x46AwDEdwoP4aMpaqTB765KhA6lTxAfSzDZtBVX+fI49Ylt6beNucAkBatVXTu
0BQEsvfKJe/X3+06zkhrtT8zBF7COU09bhMGtvaa0Fg9Vz1PYlMqWmGl+bGTWYeY
slv+D8B8aeVBHgRHdOXcUehpWD1DO1LyG9XDnHkcrkRMCsKOTKpdCMjFAvt/87NX
dh1eKN+hTmwxw8QRdA8FDf1QQdozcvsBcrn34wViN+RJ8xTeg6nr7D5laWpG5k7d
ZowcJsByEzOquL4UOS5UiENyGR17aVFUP1j3Sh8Q3+uQ4THufZLoTmgGCyLB9a2K
awVVMwywJ7lt5hndW19FS5y6CHRqQlN7bNpG8ScC0xWw8RF4HkBxPn0PpJN/GHTk
JThXtWUANqdKlDlM5jlX+wqUwfN4iqctmk/mbWg2am5EKWLZIgJ6R/lttVByK1Ic
0DzUUyAuKKjrgjnPLOG+gcjmaHeq13vTiwTecOqE6rsa3JsMOcEk4ESh+uAZN1nv
EEMtLr6Gg4jLh26w2QjcsMdF9G31twWONU+ctC+dJbkjcER2rEaEINabRRQZ9kCV
Ehl46AV1Td0qgdf81q+7UXKfk60ky1tu+e0D/XhWbzfDcwWuKfjdeS8+1ZosddnE
S9kt4JzN1z1at3NUSKELDLQQwyAMyO1qQlTVwfMDPoFMxVSKEECeKIPn4QW8gDYG
DBzGd14mfw6DCh+eDXWOd0G/mSrZ77HA2pRF23s9+6WE/7iAlZHUACEg8Hodr/Vq
lWgJHnCPSiPszK/YHTQygYSVcfAgJjaTQ5JhwftgwYqOnvZHqNeqqkjrEsQMNvHp
glPLaGln05LHHswU18ftuFELhH0Xcq8xub2hQR7aLmjaTUPzKk1+X31d8ydRp2dM
t6a2nCx50dkuvdQAdUXTC1mVfcVsMM7jPftObRTPDwSLXsUiof1ex5Ug2oTADYOA
fJ73rHJzsQD0RZSUish9/zbZV4V5cOfJtJ36D8nWkIJo++XdiopHwPyd7L7Pfc+k
pnZLlwYG5YrtVjbiz4ZkR7xUIq0JPzykDeGTrfGx1E915bHAmcB8SjvGlUd1OrFT
EeXUQf3luO7+aFc8FT3Sn5Y5nrtzgkf1+iiSCUzty+8+Dw5d/51MsHoEj7ff4sMU
NBC78k8BAyF1G0Y4EZEOiE4eOLbf8xKZ/Mw9AMDjS+B8mt4/uN3fhY/445Ep5RMS
UI/NO6BBRa0LlpqP4/5EY0srU6aJeqiX7ePtMr/KhPtzvtxWZmkjzm9+kuvUfRwT
aUE88dqYuYiGDwTv7BokMatxaOLVffo11s+8rY8woXR+NjznIobfjazkittzvCJT
EDZ9lZA1CFzCPRRe7wp8keGmoSW13dxiIdA0yqvZASIdSA2G6IlFSskASGjft7Bi
smjs9KozdzCf8jHSVLe43ZQ+pQT6C6pgS/qEqdi+xs9tLDxjGM99Ow7JvnUfEunZ
EfSYY7C06MA6AIdyw+A8W8p0noMnUtdb/RLU7SSjjbDdwzaoai6+/3eyfo9VO5mP
pI6kHsnNWUrjcN21nLcVcZKI16oadMcLj3XDGb/dhs4MS0qaj5eJ/xTo2b4/zlOS
fpLOCRsrGRBNxK4yRTQ8ttVsWgXUVbB3Dzh4xVtIBQv1waIgCpFNVrnN7Vtt8cs5
ZRwA8MuGoef4xwU7ZLJQhus7o+RI0vGvsZoQEYZWtVaAUquU20J41KJnWZBO9ajR
FCJriRaSLy9fRH7vHJ2MX/iO0CY+m3r6R/CQQf+twkZ6S7Wo7ZIUDQBo4HRGog+X
YSuhjZHUSkrkVdOAdqMa/4mm0Q4ZQIChT9CFl/J3bW+xl6CCMr4WTgF0Y86YC3hk
t8VtSTamMGGuNvP8gYJwJjNevhQy18yGosheGiqyHts+Vqk+tQOEvQhGwP8fW3vQ
/BIpK+0DvDZpyfp7WCzHrTHXp8C7l/n3h2OLvcWs7BVeOznmmXIqRv5bUHZzonBI
SvOWGigoFtjdcmu//C+g6mfRi0mQR+VtmIadeVVQq+ZEj3MhUtkRviDiuDhLVWB8
AOw9NuusOjmYY43MXi2t5TZDdRuBhxDRXR0kXRi7jFn/ssHnovCL8g5yqmGMc/kI
CUQuKSCeeA/w9pZ3j9uBPmrqapzNiRJYW3tAHQAbk2tq6y/km6JTx1pxkb9rO1CK
qLPx41+kBMCr3zv959WhOpgVkc1zQzs/AZg5HlR4RNFIID8nzcnQZU9Fu6RxbjBv
mA09e+XbMOFcsb1DCv6UEmNf8fb8YbbhIV4Z2cs2AuZR8s8aqyeblWF8TleXoc8c
mZ/VVpMld83ENeyQfDUsa8Yv/wZHQPsENCb+7hylH2EPKn/wJDiGs4nQXjSyWmmn
Mz13V05I+68StiYNPoofBp3w3gdvuzZBViqNlA1Ga5gMADge25c5lXAjhIxCPSNj
ALMSTm5TklsvCGvug51acsg4kXAdZlwWnl72SwxXfXp5iPX1fpH04Sm245BI0Sjk
xk707rsQV196PxBpO0mthZzEUssEjQKFCMfg0uVCvWMHE56+RIRe8NOpcBKlX7Po
BGLpLFm4cvEBa+6I8B7xNhGD21g5SJlMUFMX0DpIuLgzUhU/QUflK4plTrnimc1n
FXqbFDda0zP75QAen68GXi0UmRaAi42B+pwv4kLh4cGslEZiPf9pMC8qvmZRPO+3
HSKQGe2U51ZDM+ncs1u5MddQxPhbDqUxnwac+Bc6tNoX7/9Para8xC3BBJK0+eYk
UbK17MQAPjpMAhjtEmfMcYgw1KblKSnGBiX8kIBDHWs5/do6xndWqD5KW6OL4WYu
wjW3puVr8CSPdhhXw2WsL302sD2plhJcC9VMOn7PvRGmkyvbZ1/IKXrSq1LbMbBe
8ugJDp9x7w8hyj0dfO/IxV/2IyLBDGw8xDoAu+ciHPhJV89JhmZKqm+61JoRb4A+
UsLkHqWSByjJOKJ2PcEfPKxaVMIPLAl/wFFkvVIdHDPENKzi/4CAdBaNWCVtUV/Z
ChlgoPt6JIqlWPFh1kx1rScYV72h9zrNeQ6/DGprf3o06tgo0vJArHJSb+Ga6ThL
9e1KqapJVAW88+vN7f3zW7FEFrzt0XyytBxIrSNcjbQ36tzpVpq5Zc2SJlZ9RN9p
qJEH0hLHb/3gHYTLBuSnMsRHYiJsCegGxbPTWFus227RwPXPsGYNElq3gx9REyws
TpJxyhwm2q0eKHkHgXSEPPNIO9s9uCYU2FmNQ8zTqMYKqvjK/0+nR9CDUIWzvpQ4
xeSd3s5CZnLao9aue1khLDpwnlkZ9inJCoR0eo/lrIAuJJwzmYh00xApnKvB1Anj
j7qAw3wEhIkxjunoelcQZHn5Pz6+gVYMgS9CziLOtlvXDcIWyXVHWQgqX9G2MCGo
0P6BvlxF0lzanHnzAyLLYbrp6zD8ekMAHVYNhUmQELWSG2tqFRM1qpAEmW6pWy9o
BhgY80oCM6M6Ka6zTdkzjHQf66zt+1YIce2rlWRA3GQGQ3uzBIpSamjmaTU73agR
55u80SLh4GSRNQ+saWPUD87t+/T/TtwpfOa0T4g+o0V43/8n0VRyPSAsbcKhMKgs
brvqn/yGRCUStMee57LCqJadr0NCOmbmuhvVIQpVkAmhIhSNYNcCn6rhMZXAEpka
hG7YdOeXL1YjQPqk9qi3gDqUNgAq93lgz55Z1XHWT5vbX7zkGQO3Xn7VC/SY/nyx
uODB1IpnwTqYteXG3UqHHDVySGZpzjvkVvhETrGllB19fvQ62WdEcCCdrCv0RNsz
mcldV1MGibl0RLyMI5Kow+ld/9aOg3c3961KeCy0IhxQEb7S3WzrJo3zWB/lusPA
zxWKaFtP48y1owsaK0PhHMo5HDT9hgWO52reMGeRM1EwxbMlVm1MzV9CTYBDDzb5
0b2fcUKocXpkpxKIGcu6GoNpHOQ6B2lzOx9dnsrdyEC32B7/gfraHDHtCIhbIXRc
2mQqseGcKY6QPHCB7FoozeJvMVMjB6Xvn4gb0HBjoJDqc6ZRuZjFnp7UzB1vdfRp
mFmvCFdpvxk0FZ0MQI0V1d0tbKkl0sNlhckoxsNXsR5vmuP6rQgGjXkjYz7/oGYM
H+8aJucATqAfMwIzZMKU/StWh2N1sOjGyY+h1/N1zFoIdtJf6NveIt2JvJO4OeoN
lpFhfxfLNx+C+E4fZ8+kagjLvO6254dzgI2/76b8W+1NAub14vTvMVUCGQfcl0Cy
9Zz4/BsBqTgHyPcQU5PIjj6lGTtz03uAuk0oBP5jGIHbgtFH2/VGOJOOwcYL6c7E
oEZxZsCAIwHftoerxFOPKq7l7AXP4XB395zWuEf0iXnzsur+ZbE9Q9auRNG5ND0K
fAyS+iLuisFMIDxx2JweoHpDWkAT39j6DOO3S7zuE6A+IlTV0sHVBDDF1LMlen/l
JFWW6AofuBgWBJjv69dMGtuDKw+vYvHjK0uIgKUeEElfQKbaXLLlInANL43XQi+0
k62fwRQFWi/+g2uU9TOoUifVTOMqqr6nj46K/24N7mRVd+/la9h1gRGne9e1F4yf
rFJX8OYG4RypU8c7H6F4Bg+UPly52n84m280GeN4DFRyUJoTMUAGWQg8e2l8pE7f
UGcJph3DzjwIgd4TBl3Kf9paFv5A+Srle625Oju+3YHc9ZccUrSU3WbKlpPcHsWY
cJFg6ycqqFn3najuFV6vFNhBMtVgKPVwyuLvOuDrRD3gQEMtDNCFJdiAAHDsf5DU
Jk0NQCJR47o0LYLSiEX2BOYIRDNjZ9NB1cWEGpNNcoEHgRMu6TJ9fE0nKChguTkk
sBXg2VO3iOZL3edUxeE/eZW5k7SeL53+6evJPebzrdPoeIvrbj+dbZlJmI+pq9+A
LH+tmdH0IDGX5tRyv2T5EuXDeH6DlHZYnMNLpC0KrbpEKPlo6saqd4WdwGBi07Om
NSyoYCoJNaqb2ckbsds2HUyhMRHJd/Iok8f8JtOun5FtVtomQFnV8fJyNRK55Fbt
dwA/1SonEMpLw9pYw/34TW++ivFCqrtFc1lCG9SUS0Wg0Xv2j/DWrpiQl52mw/o8
oYkvTF6Vh67+qbrnoOJ0NT8KNEswy5o9nbbmHDdNVQpwpw85Tsf/ARp09Dpq5Veh
FMT8QoyAoLkZ6Q2o5J7WSw5OcqRMNFymtan9Bt6Ce6Thz5zUPQqrQ3SQ1T5mObJZ
peL1yzBszK6ChEeYuMyPoDqWAnyDyi1g0OrmBwZQfBSE0kxJd5MVIYjb7aJgmdKL
ExZuGkg75ENo1Xi9fpF7VULr7t+fZtyStvGjN13xm/acRlzMiEFTSi3V3187fmcA
h+IkfSFvs7Z+2RwL+4fKl8phetLXcglAJuhulxX/YWgTfyxfkrpYAS5U8Iv6mW6r
1y15dxPlV/gyoSZLFuV9ds3PXtlMTAWZVR63N2qyi3HtOFEgzM+rfqnrgKvWhPnj
gXmayBx5h7QNqLDyBSsyzcAXbFe8LQO2pOgG/6cg4GDnhjtNhG1TvEFBo/ZMwAs+
D1LHsyo0ufEJNSyLkNdlJW+KWlIi33WGeHIOC0kkp3KbRNNcL2zTdlU6VY37EVzb
Ccak/5jJfQ3AWSn0St1uFFucAiMKjTFXnQM2240WsRiduGvzDZPVOa5b7ItAswab
JzsIVtrMuKKxJ8RiUWbyKkgUvGCHGzskuo0gJhnDMGqfZIjKX1JormVFtzJZCL0C
EZf0j+4lYUHZjcLywXRlG9WknAQ+vmEvhbQStJOtw31WkBMmVRTDxlW8cmKIY022
s5HoVV6zFsQpoCfJu0/fFG8UO0KAed1cf1iEC3Y2hbGI/PeJvKbUH3BxCWz//7Wi
mXK412rD/XorTnHtE2LQAJf5UfNu0SNcjXVkph6wFlwpHn2ESewZENoQ4XHZmLrW
xjJNvSS12R7aEGDh7Ab5jTncF4A3mwjx2FD+4jQxLnloJgkHcPnxsfVnJ6pM2iRF
84qrKXVmuDexcTuheLoSZBJUY5DWeueP2JOrWsWqJZRudNEe8ySYoiYEvODwsB2U
Mifa16fnQKvQ0SRzNweXWw0mwQ+Tokl7DZB4VOLOHQnBRF1bdqKcS5HxIqFpMCK9
SJYU8WJHmsL6bJirQg57gtDOjUf1aM5PAXxqEMbijbV7uGwrkLWOFGBQOi4OMtqC
DFPFpURmsfVATB593bGHS+OqigAxjr2MQy1+y1EWogHzB9UBfn9G6WL3XcdQxfUG
TDDF4gBu+7f+dtONIdptvg3vd8aGaNoxd8zC1I5gnx1QDc1tweMHza3ZDAx6mINj
Ak3yXzIX838W/v9RKzvdOEhWHSrdPdmfEhQSAV7vQjRTZ7rLMisY/p80zIEve11V
1gF0B9qySltPoHETgiaNdCe0m89mL/4CTyF9fdsKdtIxnIsQmg6EheVTZOSJ+XZp
Tyrvwu9EKkRKm4tOngkq4FQicvDc88HDykRNEyTn+2R6wY4cpZG8TJm/JEsgkbNI
JEZKKAfz/Z8ZtT7ylUtGEUAcfdWXt9aawf89TmN9FN89SrRdLfnGnl4rZh1+WDRS
0WCcZCxSHG4+44bspsN2IdXk+zRjSrNJEQpwID0i4mT0YU+szuarSWK/U8ICKTnQ
liIwn/wyrKk9NxHwRRgfe4gI6XNmrKwfqvH/CeIe6o9PhCGR/J44uHBZFGz96Zow
N3WVNM7rpYfl+8QATIkIGZuOpRREsBRlO6ImVbXvxdFQ1NfHAzVftiHVde973aEc
j473xr14qBuDm6qWljLw7vaHpC2+qnnFtSjo+EIEHhLCRvKvgfrCsaTl8jaPKLZ6
CUb7jHxw2Du1s/YvdxNT17SGAlfwNtJmfFpAtcTGcTPIqfBltuUbfhOzhf9dsRD/
1kT/SpRKGHteqsA4BA7ER+GfoXMltLKLPdVf9OjIbIE6aj9r8wXApypki3GxyrV1
7BhlOAAD1sK/WSjNenjfDnnvP3oGnbV+aEw1ZYx1h5IgEdlB/Hvfddt9YIebK7GK
z15JEH2K1u2EQHP0p59yvCmVf515EpYqggTytjhlX7TlDvQlM20/xVPVVh9s/8Qz
UF56r+f7ySylwQxnhOexVcM/fU6WnAfOgHzzR9LPtrYBeqEb8fYIEzn5S2oWJMqb
5MV+iEv2mH85brvBHbcxFgYbmPyEBtS0eFXvLXWZf3+ap+klAe5zRSJze890WCTK
1OiyRxciND84323z1lnM8FcEjUnrW8xmWXeu3J6wYw4xKVPEoA/WKyUEc3QCknPH
JqG0lZlj7sa1NtBXKjVOWg2jjVus4QcIoTBhaPMSSQkmabtYcGtXFJpKRWLLz4wI
sybHAkLlBe6H9cJJizjXorbuqbO05r2z7uUphJvybvOrLtW6rLWWXveqCv9pB/nf
Zdq4fCr72d5P1h5EF9FwW3Dh06X2seV5/6iDrZ3arT3dPC9XASfv60YuRBtDBSrt
Frci1VcYZhAL/rD1z3ysx5TauxEcauYEbC3h8/t+Fwk/nlpZUsc34figqKFonJLC
ZoZM1GnY7TIK/IzVDsvS7+q2sOHjFJT6ZPM+0ceHH90kRVYS3YEKkH+dnUDEEs+q
NYMGWXl1v8Qq6Znw7Q5gymYyrFxFmHKHRk+pEKEo/9FDUraYCXAYp+xwFoLTahin
1rbclms9HiuInX1zwyGb/mZKJPFaG4qYzOc+atD2dl0JvQMp//hLQXnhg//wjYiG
Z5dxiEbQEKHfACSb8MS9lq/4WHCU/XZrG7PqHFUppWTTib0KAspwOeW0PO5V5ctj
/Zps8Ja3hg3ScSWOcc6zyX4daUvPTX1ti3qpi0VdNZlFOgL5APWmUMEFulzSJgsU
+l63CZw+XBDOtQZ2A4G+4CDysxmxfgZpKOUgeh+Ad7YEP4IAM4FiJZUXL3jHAtMs
G7kNZfp/sakZ9b0vdUbD6b3ZuMOXO7esefgjTujCtnwzPRuCFAnm/j52+p33OLv8
CCMxlq//JuvHwU3n/giwy4yL2fRWWV4eBpwZZ3nRxLjvb3/AWBXTSKxmgAN9DTCp
z+bmCM28nGnPyqMZi8WABtQ7OzdhC5bXB3UX3AY+8TI/DeyTAAC7SdqeHnCfioXY
0K0xEXiETLF7nOEnP5Pb07X70C8kp1REPtoAxl5ceANib2cXq16T1UvRNUEUvjiR
J6qQ6zDFeeeBngERCvO801vLfr75fBil4sbmuwFox0RQ2EyqgAisgfGGfRbroKrj
8bcoxN5tplkwLfZnCsF5BAMQg6bXQmkSskH2FId26pOBosSZXK8MDQH5AGqrulOA
oqCYOfU2C3E7P7BdUXAeFmDahwdSreiJX34SyDGvSdcs8Duad9hl347f7DEHeizQ
tvxxWFFLgoPLkGYZT3vcqL3KSB9uRuVPU8ZGB8u15/BR400HQkBJvsTtvT49WSeU
yoALgu8pJwOMKUxaowqdErMsjs9bJ57zMhkOGtmI8wvOBtrMzLHiXDtW9q5rLQZ5
HjH5HyL1DhNVf04nq/sQbG61WMoolysnDCZRE/edKVNrjg5zOs/FVJdDpb8i1eT6
LPqprirPa6WOKof0cmvkFKC6eCQiP/XdhMscuE4j32xxW7eJw7zqgRMw8JlTwTsZ
rXWRJrCR0aEOVnRHZ/kQ/grQSWVDWkjdUZiEui+Y+LNiRTDGS0lF+ADpsgqFGJsk
Vn+pqo/rLQ0gIRrN7+lQEqk2AB3byBQbQ3YKEidR5+dJr3XoLfvlwntygAuqhHwo
RG5oRw1yNECHCzTnWBpg3axNhMWLwxFISVGYzQ4/X3No36FAeekpPFHXmkbeBX1/
OtQrj6+Of4t1TkB94ALOviLPAx7fY77SuJNj0xB6v6hBf+LtC8geWfH5Z0fUP6gI
q2oe9YOpRQuy+E1DFrysFdUJIk0p2RwGOKTXgtWmKtnq32V7dIoaavxoC83kyVjz
SeAm33KlfUX59/fuEjT2yHJY5f4FrRhpGNBQzrBXKfWPVMmVxuOTXpuDsKYdVl6G
FD/1hxawg8lAZ2EXNYUpaMUxoblGhAbiBOwGrHNaTnfUgVOLyK8GIR91yXJdg2Kb
SsessgMDsMDyvVOVz4i2AngzKVWuiaGGtPUdJot2FUaDcnd7cGfk0IIHknst0o1o
y4n1HoUOSJUkMd7l5BCoH9hG7qcIsqnOcSl/yyVqfUPJ8djFw1R35/638n9MBxNC
suNGupvyzDq10czeMjT/arhsbeRrnB+9B6jZDyePz6Edt0ib5zckxLppRMpGMbn2
lj/ow7xuJ/JBEXOecfjCL5sLugNWOmAPW7b1igvOwCc/Wc22t0cR9iyHtUPQJv9D
MbDBMgtB6pjwWlFv3Mxp1jnEWXep8mBtt5u/VbcSQiOxJlN2/49rPFsvFH9OljPP
P+1lXbzKkygtLpheWzjV1F2t5gJEoBOB8DVc8MxaQjPsRIYiWHsy22DpbKH4s6UH
wontIoHHyy4j3Ihislv37FpRxhb3pi8vcGFwNYywQEpX/HLYfqLQ61qnAAkysNxo
nGQCX3HGl6NZbOtfwXM+ZZa/D91zB3TQAf9Wul2dISO0acf/+0bqUHBskYmG312b
Zt2v7N1m+q+PF0pEKo6t21AkxKaaw7vJf+cbqTqH+yW0e+t0sJson5brb8LfUb+V
I+HJ3KyKuKCc4AbykCBzV/jlFSKlwkF3t+dkjHrlxzXyUvT8eiBpKCLeewUFGbiL
Zr2N9TjRXbdM4NFiWile4w5JRYLG1JgkpGZkReUV03rd6292plF2DkGQRX0MSejC
Ml0Gg7hb+wzpATIzt5CRqO1VZpXlKvCul21G8VTRk9sjt0AOekElV6ItRC243Wn/
NHFL/762Z4WZjowAkWmrHlR58E/s5uZUdFa1qtAtpLtTxxe6Q9Lv80gbRjot7WhH
fkh1i+MWabs6lVZWrDyfiu2fhqWHlLeIuqrK1idPdhgVLMCdRFkQj+M9jesw9Jwp
+CxAqyuOh1ulUu3SASEjQMhDVv0e72LwEaUtsG0o4uBTIqtEQVNyGnXpWLu3puT8
JCJrIFuaUXZENrtdW5ls8o97y8M/dxYPf0vOSoZTt+RBfgeZSAhns/mKtgBRlXwn
XTa2eyA2HKGzdxlYfI7ndY6CrUoy45ELoprSFm3d+nIzOBN/VZ8RAdJbDBJ64Ubj
6KOx/pHIcovjTs8QlmbpYifv7Cc/oUAg0dLZIF+lTzh2NdibvVlGcbVsVZr/Mmek
gCmt54Rvzd0ThjCtCZPDte5GJZkS0JUREtLLxlpGK+4gPAp4eZOOi04dK6sFkGUP
MwF8N2yCAN8r+3rpaVi28JX0yycvR/KIup0M17FiuP3XjT/VQlAW0QpSskDRV5Ww
+LYlAo/ANMP5uZwOzQal7ujrUEuSzaG1zWuBY2c4+INtA6Bwj4c8yqsoYT2osmpa
brhJXjMw+SXGF4EtgECvIXeWu7B7I3sMrcokJGMg+KicKZbvG6O7SsPb2JOS7F0v
rxJx/7w2X2M8C9QsHgtdez4hXrH/TUtpyc4Mm6e+sPQR+BaOa29bEAluU5zkMndW
8BMCXr/yCftROvffjlpQGNOO/R/k9xHVPaaRLdES9cXlbq0q6Oy/wrfiImLyG9t5
X5qCiOZv5LDYQkEWHIoGC7F/wQliB/PuGWseSTA8Wtb0lFEI+gemGPt01k0tP2gC
1hECZo8tmE8/GWnl5f10gUbJIG16KZiYyr7Sek+maDQOIoyEJ+8nCS6lLbdp5Zpi
QnzulWwLnByU03zZ4DB1xA1SwTge5WAjJcea5lGfnot0xWgQBPWCsHtOdzV0tpAo
R69j5vxFvItzPhjButUzI0I+yLnjx/d0hrwiEk/QQrVneiRTbl9donIYnLQ9kvuD
1JnMk8klJyoCJADCmG1GltS0tHuwdO6lpc+520H42vXGhe6qRMOyDBgCyosNfvje
G/qBvSs3vaEGTi1ZaKVo4UCS4//1aM30PwMwXs8UX7buAe0P0t46SkNmCdGd97LH
bJDwt39GGSiqPCcFWLYi2F+XaKFbvMCiBhghP4YdMjcnht35IHlYM2cg3SHwffBi
HTXyIsFGusNRhc/ZU5WWGwGhDKRz7x5iiT1+fXb+Bwn6k2WV4GysqnGSD8RaRPDR
6IvG42lTi4xPqVGSRSOyFG3zCIBtUeHIuORaf5XY5n6zLMTYwuigN8vinWawqsO1
5mn7mqztxq9NtHhWgZ3F0807a3Jv/oeeNcjnkO6SkJmZu1+fQzYb9zwIomyaG9PR
AsspnjvjpiEFt7h6mIDbFMMVHy1UBQi5iY4sAv4p0q/hP4tdNlmxvPv+pn2V5oy9
Mx6UhqXfLEWJaNiZZYM69y/Xjq7dRTRq+zflxpRz2brA78zGv1EhXBtaroCMhsc/
ZvalWp1Wg53uzBWtaJLeWfho2eDd8EFPbh/Z12006VewpTSo5hRHd/MGPDOL9SDo
v3DIcdu1dyF1fB9e44/i4jmVheKJtpd6djGRPis41/B0TXCkrX4wW1VbGq4mTaz8
ip5KP7BQ/QQ3l/C5x2IudwS8A9aQulizjxYfRjFcWhnBveQqYHpcBoNDbyIqNlQR
AFGYgihQwBSiXG4IQzPPBGEUPRcDzvfrQzydjzgtn7DFOo4iggHd3Rvnrux7b+zb
3laevr40MEGfaTKv4WJb/oB9DlLj1ZmVRZlYfrJhyB+EnEazpz7WQ4OqzXBcwyOP
JCr1IN1qA/j+VNsW6HNcc+0AyqwwWBG7RgOrTi5a+d2R4ZHBtGlYlw+9Rpfj+ID7
7KCpgG197FKlpdXl9saOab96GPcnmv8LjTx5CuFtyA+BSE0RHH0Z6qST/U4Kpm7T
WxCfnfOcc4Cetl+6WxuRXpUrY1oEz0D7hINlBQSJ6LHSSN7m3EgLtv92OuJURB1k
QFjx38eZwJQrAB9ky1fYSW4J5RldEZKUgNvPwhkPpZLaCgWG30vSFmO92hL46DPS
crtMps/uaTnAM4uc+6Sl7u/Ol02Qg3/4C77nuMKDyiZ+lsX1/b9F1/JlIKr+VU9k
Q0bVT5aRarzRpn2geBi56GRFkaZ6Ke3JYBib+HcR6CVC9zCIsPkGf0FfqTyZXJIG
SlNg95dkpb6KHb0bK45mNW737pDVanuPJdjqROuFgDTTsIP0PObOmU51cHBEgvrK
DjNTEDaPEsynsfkHg4eBFKktJVymJ7PVBn0bGL/WB6knfCGCqRpgBNibxtKZ22tO
QiLLYUzk7qNVoyoHb8dNtNT3D6F+tAdxUB9yejU9r7jLMpCAECsbheslT9div60T
0Zn0LkLSY5Cznh4AWhYEDDBBaJEhc3sBfV7aqO0pb4USOOQdaGnI/dWy7Gl1loA0
5MZ/0jIs3Kbmj2tCfkzrnRnE2/KyDdQ26M394khSOD5hKcvYwJ4TN/PjtfGnSHLF
Bnth81L2Fcus48ATtHVsNHYJIubk3YO+kJjIq9G7psiHA7u4cJM3WHtBBCFADh3R
vx1JrNyyC3TuWxan+P+1+ysJhTAmtvH+izUWG5F5JfL9g9pXk7FQ1tw2b054rsaW
3ggl8y9fgD3ulrmA/zSrf4STJG/ojrdL5eq/PLIYvGjkfMw3XvDz6JvIDvGCl6RU
tBSxpgv/N004EN3DB860zzHMR767QdtiPZzI25IXx7rorm/nTnXG/SO+AgDkME1Q
eOsBpTBslvmD24VCACGb1/WApeN9JS5gXKMYAQiJcf7TcZZ8Opw9yyL4umzP+vTV
4pXBjPjbYyfVq3FPF3GH+T7Rb/x8OzTBUn4ZJ0SaHXukbGQxOido09WjScufUelP
00cBav5NhFhbGN4D74pALN7qszowUDTOr441mnjficjbQK6U+KPHyV0UREK4O67y
To4mS2eZyFFWkn+TdL3fEolYduT+SyT4S0x/qLXX7UxY5+Tpi9sCoUyJi5y2zGG1
G0ZQoKPXeZ7ekfl0A7K9OCpApRLpviIKUxAOXOrZnhuxUwscd9E9Me6aJNBEw/KY
GKYCcBAbdYtha61k9Y5jHCzemtVpG7BZtoSHgb0ZftwOvn5EQntJYr46kVLas6z+
QuUoQGFE22+X5mrS4a99W5xvCTXoWwNP8P5QdLxCHvrflzhPIX3SkOG+zC/VKBa1
f8qpjlwUDjmCdl+98SVxTDlafbqMR1giJdPxwhhTK98jX6P/7qC3AClJ4mIeNfRs
INuyEO1qCEhfXyrhu+W8EqrV0DSVUGUA5EdUC73eqMVrP+xF91l7KdpvcRLp+zgJ
c6HuLW7MK1lQg98gps0f/bzQBLsI7dQ+ZIEgQ+ClMUaRv5XLihev9B3khsm36OJL
lowhOGSWXHTjrDDof1+QO8FNYXajBhE/IiRfyLLAFIeGtX+B3tqmO/wzS7jhXCQY
mg+Dg6dJ5n3nDstsNTP4pS3Akw2KZQQ10HieJwlDc7WAfEP4zviFwE0ZbL2vcdAn
XYEHKE8qdosKWUMFYljxr+BXMHuFitfQS9webfU/kJ3NzJ+DJW+6rWb6ctHeFAwS
nrfAppCEvU/gWtuyfgFlAy4pQXd9O23+klI+ZCA3+LXFjwDsWKsw43MrboMCVRqt
gsm7UldPw/42yb9JTjVbY3HNc0wmz69x2LbXeLuEg7mPskIS9w9A5rRH3lVSrKa1
EEDfsvg1AB8pNfrBjerMQK/GK4HS+sgPkQlDRqkDIP+xr3FPshPlqlXQqz8GqeJo
gzzx1H4DtLYUiqZpTp2NjKu9rorsnrh5rBZSNdXoey/XJWkgemZMCQbPnZFhA+Fg
MNz6a3bzER4a1/OGnqJZGxWm9CeCMHSc0qNVIq1QUfCiOnTFmVFvDwJU+q45qEoV
3CNtjKfMulkx3ZHpSWvOanl2Cq84zZ+aGD4SUs5n4Enc9YOGpM2MhMLANgG1NUie
8brSAPm/NncheiP+w7ZQVfpif8242fBSK0B9OrM0Jz7kYegX1WEzmuTo8uASsYSR
bqRPHVIGzTVG9AgmynxnpQUMRfpVj5xeeWc7Lm3+lUi1p9qUsi9k72OCGu48U9mn
Qm7a0jR3krnezfBz74kxzsrYIXy1NnKUoVJo9ufDasRR3gw6ltL14cXH9csAAlca
n3z1Xc0YC5HwR8JQCgvi1vEV+THwVFzJXXFBtDf8ZZMdA/HgHxW21YCyZdUxhILG
bWrkaZX00B3db64Hq9MF9oN2QanxPTU8+AgyZALOR9+WpI4aG/S7WL0tEL97eKGM
vfl7SwQcczBT2i9qG9GA5pHpadfx1n9bDd2rGLShZYHLmSyAHJLyETK44prUS9KX
9PNG/ZARBrfNuCfUgXN91VXApT8ErAOkSpPxdrUgmy/Sgw/28Z4QE8FUJHK4OSaC
npKGPqfX46xy0oxPSWndkO0M8pluCE1gyfOnhKChOjDmoA8ocbsXKp2noxPjEfhK
ADObzqycidmFCoDbAcgBy37fllXLgRMQCVXEc/1FBVMgKDnZp6/nT77goXHcLXhE
2Biq3+BqYR8EywRhF/r65ZERQ6kN6MxrCrfK4Jq9y9LmKjdjmwtBG3nkf7E93GHl
ibIMYG801kUX09kqrCEdtNgHlnGfogWgLF+QnT3+n/TH9TJFAKenHmH3kjYudbHe
a1ZNQx1od4S1RtrmPU2bsblydIDh/lvJ7wSmB/d6kRR1LO581enbeBiVLUCZALub
KzZqeq+3xn5i5lamdaAXCDq4dDzMp0zpWlgW4OnVLGVZYRmR2oNwX0cxYBBlC/vb
wNNEfntxYHGRtVsisvVfDLfOM61FsgPkcnwNl/OGvTzaqVlxE1g03tsgzDo/SMYR
ADXUjpRMD1d867XB8rRu9ZAb4lJGugPP6gbMAngl1zudU/3TgSiiX5eR0aAIbpcA
Js5xLvkMLhaLg7xj4jET+sqnOC4a3uEd4rmUjb7BD11quv7Wd+UVdQgFqq1IEJgt
HLqfErmL63Ln49imv0QknDtMrQV7DPeFOnsZtXKvZgVRWjbrcs7dLuAUApa881+e
GzcP6+OMXIbr3xYZlSlw0qz6TQQiPGTaSSjcJ0OPketMVMlGRSR4MOMtftLpKE0c
KEXDRSFLq6ap4U6nshl9hyq7cIEAlndTTtuODWVMsVnor5hmGQXi6jZlFXoZn3dJ
W8OWZKUSED79rYkbYGisqC2rSsJjPxRhWBWcaU1kKeVB4YkzEPyp2CSxhswJbvwl
RSBgiXc81+cM9goPbgGB0tQwjUJ0BOERXLVX6RxLmQHRHDumRFY1ELg8LLXMR87L
tDa4JfXBHDKmTIbmpPmBJA6ymdr43D5XYPLpWdPdJkJC0fg+BDhyho3oxgDDf6QK
1mkraKDavDVYUHr2dOWk5urAbXZhiRgBb/OF4Ww4qyoPpERFiwmSYdafm821IJ5c
MHBaksV9oMrBtAGWLYWiKQP/SdSUAxs5Ozlc3r88LNEKWgVzwsgDQk41/ugkQfMF
R0MiwqXjFg8BJ2yTXOXmPRyLPTEcCwbNd9OvAeLDzkUVGTgELjhcohSAWPEwLeSo
HNuNp+h5qcemgEeWSjTveSX4ySyhH0dclXf0jauYkTYH6nsO+LWp4hd0KvphKjxW
MJRSBe4y22YPsLRNODbzV1JxFFNLJQnHtzPzO8twIp/K/gVat8++BxnqTt3biRZ1
DbGYa/yPyD8jGZBFdG+IoR85h/pP0WDMNFKua0Z2HKHw8LAiKT+oEFF4G3c7pDB+
2FfuTRaqZfvx+zR9rsdK55Frh8Qtm9+ugbQFBe3l8Rky+fqc+jhrPUc5rwkBjW25
o7ipQFIz6gFzi34QYwJDJc1Sul59VP8TKowLoZClu8+tbgX+MDvlDtcAHo95Ukpi
DrHuqvKnXgIU9iTjH7jw06a8feNO4vKMHjCcQmCrhg7eG2sayqnMo5VFFW92yWFN
JLO73sDK68cuNMdi5LmUZdzF6m+Gj+/eIp5fMmkldX1VuaExuICgpPQy+F2FnKWn
mz3ym1N3YO4paej8huubiX/RAHqw2ygfX/R27nvnrAkXrZdoELr/Y7aFz0omddW9
qH1DGkm36cR0grvJqLd30mbXK//etQ8/dePOmaNiTlbEUVtuY8KMTmnuiheSEyvH
VGMUdkkMnMe0RchTb8xV2MQrtdfeIRQGLoZd91uckxkKKJ+jXJkQaZB62HUn/XfG
M0NNevthhwlGmjBZgNw6m3jh5nEakgePKPApsv6qqwxVgwEGK3xgUq+wIpqxTKVW
LMzLOlHr2IlyEX41aJcnxk7r7Nhq7+d66FbkcBysfX8i7NNc/09KEJvochk5QPnL
WWtlsAtstqaN+OBaopB32g0dmesq+/KdfJc8Y8ILlC1Ljxd1kOCKKwq7o0bLvdnu
JZvK7NJBpLzdvTOLGhCdS7aL0I+BLXz5WC59lL4cFgNPdHhZS9SxyBMoHMujOziQ
7Z+cn+IIJNWzK8PMValQc7sdrncpmGviZSks08RVOFebN7QV8zOZxwoNW0sg96PT
/gOOFPGFI1R57pv9MdofbyvO793p9+NXgucJ313IJOXQicDIehtCWEnpvzMlZkE9
dloNdWCVzhJM5R6WpEiDwZKMedBuRSSAmi9vu/Iifvx/PfRps8cjQysHlggngMa1
G9a0shA2SPUM7dsnAnJx5joSKjgWSWT6uAEFGlcnFHIaj8TuyFJpa8cQv49S45GZ
gRbt9XUT5hYdvZrgCVySj4BhGFLgL+oKpe1YI9mE2HNV8HLgxO1gYFqO9PHTarzb
plv+xukfb/pjVG8YcBWYw9uzzUepU1r1B2p1tbUK0kCS/E8amblrXK+GfNXNe5Vg
O3Y+K082AprEeM8QgelN85s5SdZetUNXhMDfYiKS26N18vWVUJvxeDr7pzgsfmXu
78LhAjTrOEmKkTgnm9n6xFXJZ+VplwxjaSBcJIF5JBviFkx92laoYh3SjEGFP4gJ
LtngLe9GiGAX/A7SSL6A6CcwVfiO8mlvC3eqoIblTjdV3AqEMFvbrzKtFBRu/sLP
51DTSro/uy82413TglxZtoqxfnGF3Ht5dA9LqRfjNvsbQnUgqaG1n4eqCQlSx85A
lvwzkojJN2G+MCVICIH1S1s+kbfCOuceXkhhieou8H8uIuAcBQphNo8/nvp2VFQM
kVtYx/TichIDommqXE4JyQc7rJZxc4zOa2U/NB/v1pbJ8ypFo/RjDhtok3MCb7+3
iDq7uinLjCYDpoTWKgqMW/BZ+meJP5x4XUo5PhSyHW/n8eTgD3a+hOw3pJsGDhz/
SfZVrgAi9xapXkF50EjFc93ZaIdqP+K8RNUXbnYKyZHginK/6XRc0/UvgrYAD45t
CXTDCkJNIWTzL3XOVO8B86MnPriaVvoKqVagYEnIdG4RDnsirGLqFdiFQtNREPrZ
jH4VNSbc/LR2etBjw8fn/O6mekUnuNpxt6kHC0QBTWwdhNqyHL5mLny/cwjoQDKU
fJhCgNx4DBXdKveKX/Go8dpi/pOCIbcpH52JppoF9Agr+s4y+XrFS5CvJvw6BK/V
tDwGiWBQ2lUYHmTCY7IA0aHVm4yGu9wgXauI8twZJ0akH7Fj35Y8GmNLNOXRA+LE
ZepPXvoc097jVBTQte+3nUqrLSydc6lFqILsEBcS5uWN/rdwhQ0MerwsGMgvLFFu
sa1mpmIToIAdfFTWdvdokNV7ooIkI5qyWm14MmeS8KAjYaF5bNp6jWRlNohZWjOt
r0WDdZA16gn5v+zHedypBhqqAj89TWdyhhfLyoTIqPBQ0PZvcnCp5DaDfTKUBwY1
OTGusMTyDe/tyIvRQeoTPFCc4RVQeVuiFFuwAAmoiilijYpXEeEc6eHNxe9ZUu9r
bdW0WACsMWwJUq81guHWIKGrDtX9pqZ2IdhfxAoE7zM1ZrfxGUuzfyQG5KrzQ4hg
qYvouu00mJ/Z27bMLKGuH+7ZORFH9ljQPhlVGLNC4CJyhP2wichjsogleSRg+Yrc
EqDPEMW2j0WRvpKi2l91s0BymTM7Lcc9lYU0TBT2kubo4kfRSjqDilHVP7wFD1Ua
Bu3LQt4cvBr6K+ph5vcGC3MJDqoiq8LRg4QfLU48XOa0y7Q5GO00sPaMQOe9GUyP
nXyIs5MIpe7jX5FHZ0ZxufCmZ+sXgHSR3vRXSPeiOdyO2grPYI2bf3RVFpxulDdI
LASzvE/yjE10edkOfYf8U9ZYDWMWVWyBjzMbNWlywOSB62NcVizHXgL+FqO+LXI5
5qVUqSn10rj211mP+FXz/4tOMgQvd+4lbqzgsdzyqbWgCmDlN7ANaxp0lkGl20jP
r4fI/T6yIpIQnt4UZ1sTUGopf+l2Xs93QKOJNGMxQMf+Lv4FALoN/yBwJyXUAOBU
2pTVfDlHm6TleiyNa8FIqsLVA3cDcNZ6kppPlwGIGeFekN+HKKqhb7iXNIFMbbfS
v69WQh/DyaK7811V7sA5s108sWXnHfFjHil5g+eIaFxIxRL4+mHsa6fhTCndEIPD
VEXaekKq619P2iCx6108/OoefIoAVUkRXzuLl+6klwlzVMupEM6RE21Q41unh4vg
m92gvH0oMnNztLMFyMlcyGRV/sdzudrG/LagJP4Z6h7KG25hr6lTJ7a8uQAs5aQk
72Q7ov7XUfMgbOZ32sV8X1kxyu/5QoTsyDSgRAd85fwpIFU+DC+k4JPp3ndOsxXX
9X3xqYVmCwqEqGNfHG9pU/WTeFeOlmtAQjRXs/VGKiID/KlMAKbm2693A+DdmDK5
ymn9rAc6XFyMpWzoPNqjpv+txbJVEQGTdm69U/V5wd65cDEiWfKBq4mncJkhqcmT
tpcraK1i41qMqBij5ABroWZ96aeqPt/9YqeW/51HImixoVlfL2tl5f4SA5PIZqpa
DMgYOdfTLLY7ylvlldAIPx8dyze/+UcPy8BdgehoRuLppb7NPO92myScXLMC7Ngh
eC+d7dTZEuXpTdQpuzwTQUTCVxlErqPBtMBqvNqExyDuQycXCcRw71WIyPp0x6pr
TCWVUWZdyl7rFif8+36WyHKLozMFq90lYCLmOIt56lBGVP0HgUivAM2cWA0unx6l
OewnASJtCyZLWxEtCxY9iSrnkL+Ru6GDGQdpQkFqB3Xp/CU2bvo4Yn+U0C6krGYb
Qs6PXgeH6xmj9AN7l5en/VfpyFsbRH6beqTw/ZkBIU1cSpJbcj6FmuNMWI9gjYJm
sN9tjARXjnX5EDOchiCzxZMnn08fNCbkGIQ7rZcEfdzcCZSQyw1wzp5+uxMDviT9
Jt7uzndi+tGYlemXqJ08z9jClc0vjluDSsqezpxiriUCTpB4kTy6OTfyMvNFHgvB
Tl9ubYVfdtQqahD5Z5L8oVtXcpG/d84n/hMBfW6E+zLDm/YMrvQwiE2Sdre8Cw35
K25GcJwQptMBGRJgrfVZ2FXeIAlHrrOmyMdSflf4wyUj2Y2f31i1nND+zquNl6AY
5/IaWN7Tllo+Vuj2TOwsSVWnXu/+uXeYFJBaORYec7WQFqAbJAdVbz2D+BiFAQoP
2l+Os4+zNQXMrgX5kdjcNtvSjs9VckXzTlyP+KqhsDvfXkIl4UdKBOxQtI3cgSXC
Me2sWLy2dRJaZCtU4qtq7pTyEzE3fasu4whcnQ04OM69ohy5WYtuZKrKlY0vsw1/
X7haYDJWexXaeFctImOs1h/62tRyMmeRYszF2WGK4UorLIvPPEFM7lTgsJUAHJYY
JMya+NMB5d/xdRxwxyQkZXAlWvHPxrlMAQrB0qJZsC/D0XvPGmbL4auuJLnmgt/P
75aSAbUNSqBhXP30Khquo7lg/S272xPlvFvxdJRwzLqG6o9wes1kF2Wa1Gd7hhRo
WjuWCteuA7s10MAtS7Ta7Y9KmxD+DsXwSAnWDMwKeRptuo4pPGgsRBu+AS503ekJ
hP+BrHqGDseqREYdbNh53ZmPjJhhJzZpqIuW50tLEikW1Ynidxz4mkw9pLyrG2SU
3ntlOwQL3mtFM9XkZpTSRaNFz8L5VMmdGs7WM/OjT1lzcedcyBtEWguE5bL1o0yi
0ZngX+43MO4ANTTOoNWgeH9DgroWV1HM5K1EKlf3H93xJoa9yaK9IfR2tCX2W739
krUvDMUA+0PuOl+W7yKxTb/ljXB1iGIy8RAlVYjP+E7yynmobykQ7+caj4ns9csI
GorgwGF2TIRYMy9cxO64Rj41+o8AUyENKlPcz+JY6lfETkvSr7EzzxGMZDSxufEG
H1X1njp4HTWG5MFTyHUb5Rf9Nn/TTBRlCfidv4td1gCveTR33dVZOCPZGmMumOYO
/rvHRCphDW+/oOECdEl/cPtXfk641LCLgH8AjODPw72nznIqrRDsvkYLABTHQs4c
MqMSyO5jyxjsQ7IXPg9+pNETynMeH0evaEI+ATldBLpmyK4gwGlLh3HlZKYv2R3n
DLudWoJM4uYKW8oihSWW5CXq/4VtbquNQadspTYcpuOYietKmQwmD6AYgPKSgcN1
ZEj2/jRiuFQxGBTMc43xrU0jXJq/e4RR363lPYcvtrmiydiYN4Ukg7npHl9BlehN
lOsPKadSvpn5wthPMoMh4EKqckba0veDs/OdgyGMZgV1sS+bVEvoAeGJjCZ9ar7S
MpfPjeqnzic2gqkhKNGG+9VmUykOOy8nzfOfcn68fHdhlUf7/ed9x9baoX95m3ch
nLApbb/sqTZGTziFLj5MCEQkuaL5qm4SLtqt4pdqchq/g9MZX9/r4Fc8+OK12c1O
mDYaetOxonxyOF4+DipVJgqzr6i0AAwp8hd54Ofya6wnTkv+5jHFawgknbQSQHn2
NX6L6uJhbyfAKnEcpCwsRdiqWaGsQ5Q+Qx8IgZos1DXzYJ10vap+q+J3QpLJQAc+
A+APS5rqVRUdhPAkoZDpE4Buq1rUy3/okiPol9Lkb1ysPhbyBaY00VU4q7SORY1F
iDaiU7cDyMy128nvXKTZ4Uwgu2YB/p3X2KzgG1NQyUTBCn70PLi5lQgIKRUDZs+Z
DfS3/AzlREaswLuyAT4PuMwv6UN01Tf8ymnK5G+Ms8f5GrI/S7cS4db7vcdDLCi7
+sIgFlQ9DL+KWbyGGLkr2yMjRC1596qc39+e1l6WHR6K1Be/FAeWCt86jIj467J/
rUmv3Z4IOUTN+l9EmXowfZUFlmZq0uP9E6GLv2RloxQpMXrBHFR0DiN86fMI4eQQ
39cQf2+wJqiB9xopiE1acwBDWeCPYgLwYrPY/6FdAWpj7ZrbBxmt5kEOsAkpHzBX
npDQj080Dr0niUCsbmJRyEuLQ+MUudS3nsh9KPPBlS8qVi4ga344mN4WZqkr+7kZ
yuCbtooWcoVjGpqO5erPR5MAQq0OxlgOM28kqHX5UcxpLvo3lXlHyMHKx/mVM2sP
IV+84k8ad9lD39fjohEuXBel+xxaeLDUhJWYlDhk1eqm/NgzQN6xVRraCmJMP2rP
HMYO0BQuD5XgB4MRk90VgOzBDYoohk+EsNjx6JZGFA1I2HA2qii2IjX07mlreUay
vn9xd+6IUrMMb1Q1gAaabo6y+wxl61WvCB3Buhe1dIk7EbbVYJCiajdEfXDp1btm
xK5OyoLeBOARb7YxYFIQPmeM6bfWiDmINO4yYdVRPd5OSYaoQ4DUoZk4dpL7T8tX
6TBznPsrp89QdJd+4811JCjXrpeTXJZA4TtfaLq/3VmW4zkG3jaMyJcfVAZDyWKm
Wmx0U1NYFrxrvsONTNqnLHjFX+sQreJD8Sw+RFz1+DAMjsONHodRhQA7xCW469sG
CEZvtBsM82m5rkEPC4dtLuC9W8vP/S7oDSUaHzFmxgJUCt4ezHjGpYOet6OYQSiK
Cb0vMj2z+OIyxSrS2ZNWXe0ieFgZHFuKv+F6J2Qf/kV3qlpdDKQ8QF0q1oiu4bSN
HoXfubbWUbFG7nuuE178GNjBocLh39GLp+QJLcHem6KlOJLpSTwkCemXZZbUOIB3
U9b2WlwVLE/knHWcQjo7SXia8SyPgbltSMu28DiYKZaiu2ejSgH68d3EmTY7pCsy
ARm1nzZsLKB6fs7QmLWEy0ayn73D+NU5jS8YvsAacVn9snS9Mx1kCCHBIhSOQ6P2
p6IjkqTc+JFVmop3rGLNlacmIg44EcpprOZ2w+TXth9AUAyy0QSLL6xINXaneObB
9p7zA9tlf8M8gR2DR4KnqQC2tlFsclwPFoX9K700YY24+mQVjJzaE1EbdWGn9KJC
CocUZ6KRyDRDsosrnlJLR29SCjS12YSEL3R9d4hqPhF3jP28HVfHilK+/8/vFWiC
Y7+l127MXkYihJhsu4PQ4OOrDt2It2wCejoz7rG+UtzVNLqFvRhoJg9EmOBz7Mci
pyN3WiERDIdvUiPYUipvfhU+Ldg3tuUbCyFavv3pE1Pj6952su4oCuJqBX0UTXFc
fxAOuIblEesm9WCRGPUmQyUZmmR0+XM0Wlpo02Yi6+sA4qQJZasERqh16CEL5+7C
oeMq0NU4Q47sUJzh6j8Gj3eFmXKDmaXBYmE4rtA+XZRKfDQ95p75FxdvboycUVtZ
2fkqwX2gETeAKNBeK4XC47ztSyOzUif1R7QZW6WO1VYDXUwTopH+wt1GJimSBcHh
Ufn9NUXMuGiWk6HsAOdrBqT0nhmNYf+dvIi36ffTU+KY8XcaJftbLGALoLaUsnsD
WyG4LbVclB5UPYXkR4/3UGF1I8Uq4lbwYxVp0ybn+PJaE5UBZh6ui3NZQpHCRfCC
hwDlEGq5FEPfqrwFZwCXshOVNF1rIQokWF098Spb4q1x1X2dwEYE1RC07Hp/Fh4q
1xSjgreZD0/J6AR3dGBhvvmOqJ16Ix0bEld1oG4X5dhdnjgKqLRTCkKmb9Q96hKU
zEqz8i1V8ayoD+FBOQxQ1Tf/0hEEdc5eQkz7tHGDORGV2ThFWrzg54baTCiUI7Ss
CTXazFj1+0QaR2gj7QKBDLnIYA9HLW+Tafmif9elbYTeupDj6HlkV0i6c1g03r7X
Rs6q3lGzVlSHITecAblf1qVThqMmRw4Dsvxnhr7KdOpH7lit59imBmPdFT1zZZ0r
hyOnqo1wESQrKkgW7izsuVDHwhW9OK4mzN4cOotYsg+QwJd4Zd4Yn8BGP63v1Ypf
a6Zil2l9s5hC3lu5RaSosU20bKnLRgDijwqdNCheN0TjYvRipuWUcHREk3/BtIka
IwhfbGDlQ9pZYyBaKAxTGNHK6AVmAanXKUdC0Akj6uPmYSMxomcPJBFgXKnZ2Fgw
8Tjnfxe8fUurasKAYPOVLEp1NwtfDn487Ilzd95uDsTh2Ua4RaYaf1uJP6ciW33Z
KbTmrOhsdUN7248SsSAzBj250XkdiI5pI8XncV8qkBtdiNOTPWfMGTHITe9bjSj6
g/bpf6GKKznUimGahNoLUeFisDHGdj/mByZf/G/esrkmNwge2ViHPFomQsDaBHPl
3Iapmf2BJWdHl1VQ/I+vyecHxWc2Cuc66R3YzkCl4aVdoPUD5yORVxxXfO02tsd4
QVbzoRVItU1G2c3cWHEbYu+vRpOP/K/by6UOjeD2qXD4n/4vb0cEKDRq2+KBxBK/
Rud011VQNsTqaCzBwpWuHO9ZTNEedb7Xp78B/gt+H6SfI5RsRHsQNq7nW83CjgZQ
0mFdrCR1mT0H9abIvvVSqHqnuKFUz97iwzctyPgc7gKfka9NCRhoVVxdEql4p+6a
dbmsamWLLWMOJnq3LQ7f0BjGPG00dymzbbufWvFclZTTLrUb0mmHVOCRW+QcLVVm
3WRjPKEXg6kuPW1VFq+nW/LC0M3mtucGzmpRpnRwVCYPu7ouOLE6LuQNTY44x6ah
YHcQ885ZV6qho6QtHsXyJXawLa96Y+J0PdmOngGCcTsGAHV4k/cuiIgHVFV5ccOP
mrELy+zrLif8UVnVWsD3+F7xFZ0E3pZ8OHbYcvRKA2y+3CkMLE5DUaEM+fvL+04Z
+KZvliknJgexlRacgkK13pMh4yEZcfnWdUv2ZySo1wRNTHq9HF2JGHtEtHLjfAOg
oazdWkv6P8UfJ6+5xyxsh18J4xZANBH6KQYYiVa/9z0pfBhekDpOjibPCOC/KpoV
/nPPsNqKQVKSh3ij78OIYfogxGhOmTaDmD69o+z1xzcEUlHDS5kgHFgLVVccY94Q
UyVWE00oWONf7QfJ8EbszyWeRv5hdTiNaAb4fJj0AZwrdMq6Ivi/t0V6Kzb86Fx0
tkcBXAjdMfBJaKetVCZhgbmLXu2iqLdWcDPGbrfxQ4BQdmC7aBAYSPlILyV0+C/x
ZNTICUBKOacuVp/mg5mMs3BJ/QBTt9hEfC3p9cAia1/+YdgOomR2w10nq7/g2qDo
mqbD6PfrNqR2Hudmcftm2nwXEjYQ7DKA+zludIg9YtxfoPPcXCBcfxgatRTvK0vm
h0mToN+ZpFv6eGyNGWyv096SxfCUOt1lZ+DoCeY8RAiNV5i6o5MTBVGsFLa4pD/s
D1KyTTwzJ6biwBwdsG8lDVKFVYHZtx4P04geRICuKfQeSFr0LVbab+35F0bVLGXB
/iVzrNDJJvJ7FRsdwH4jVwpBKF4mdz8uD5mPAzZgPL7ApXL4h1QW45slsenFh+5H
2lOoHviDmo043xXLBJZTimBBxb/GtRjycpJjOYP/bqI0ti0Byp5oQDAU8HvzfgxV
0tyvMTlHOEmdlEIeEG7nxW2PV5WyuOEtDBDeeYmQ7hZvc8OduNbnof8MxG78QRRg
YyetyJSp9G3pUo3k+ObAg7X+VFXJ/NHeZbZlw5rXiCRaIFps2sgqvP9zbIdk0R6R
D/Nz+gv4goeBBkuAHnpDT0ck42i/nEfl3LGei/HxLY0bM2dP4uZH6H6Srj/xQAao
uzpp+c50m9iyT+SPSn2io5SZEzZyAeHbjXdjDKbMFnQ7DLNLmV/SOv7jXeeYBZXU
28QFqg7wbq4YbOIMmdb5s5pHYeRKMINzaNItaegbFY3mvsQMWBeEm5Fy9GCmXUXy
/P5H3Tdxi1C7ypV/PkxSimITcKfA5T3YMDvB/9dOAGIHUhuzb6wXxJ9w0uaWbNAD
qMJGOPGN84qqaUk+EOSSx1ijemGZtMtJLGLkOU8l/X+tlotElpiE5AMYS8ib1OyB
dNqERkZcioJe4y/Ze6UOZO8yZ1QqQ+Ro59WRzhqAqhhqHOiWfV5sjyPQbweBf8G/
hkzhTo1tArKyWTVPIXK+A36K5041ZyDSAa2AHCGmR+3vyGZ54JR16UnkF6WtdJ7f
WLL1yPZF5XexPM7MXQmN0kUEP8cIl7gme4zN54w6fuGVYxFJ7DK76zS6taVvk9ko
AQfaZxo+NxhHDc1nPFIS+QrBnxO9nTJAvgB7/SuWIxu9ycshGkCPDHhN8LOm/8jt
VSWe+idauMUVf6GVr/PraMfoODjnAiWHuDQWXlZSBeFDLFrd3QuHCSqlTzD67t9N
IrqRQsC2iboz5i0Na4LaK6c2d8tXv3Lih5MlklBDAV0GV2b5qE71ufYaWFEj4BU+
n7tayLtUYOHmIQONQcgI81Ibxf926/y+zkcK9Gsi0fzNA0fHii1cfD4pEgNXphob
pnl1PHfxU3wxVk8a9QnrfZdrnbDts3PFltHfNzQApJjBy7dhG8JtU5AFMhuTUBPV
WWaTSxRFExBuHuRu8+FB0rW3aQ69q7I49wkUzgBo+PvkJPXwh0t+JMXGDaAW6vM6
giF3caztCHbDHNPxXdDyhcC52be3joH8tY1MjAtTKgfxNgYpR4cS9gQ6X1gMyTXl
ZUE9Hws//7dsUFC880VB37fjJhuFlPTxmLP+qdsLMo1K3hM1eCiOUvku5+alQQg/
kE1kdapoUuB7OO9yTSAcuG3DfIqxEbfFr1Be6Sv0JmDkpSJZhzTAuDLzZheZWMFN
ZH2algzVpnv+TrkiAZdyq36DRQIaN+sico76BzqAOo+TLJG5HcqwQ9BFG3shEeKh
SvPEPTFgxHdLyXfDgneIio9kFLNZldEuMuFBOq8/ezmnEbAoBv145KCypxUgDD/5
OVSBnJv2JLodV8j+y7pAt7k/d4m7zVdCyBKta4uvfzDKrqgL+j0BGgL+cRQrQGq8
O01cugjMbatuKnigye8jwPpc/LaX/041LZmfX9m4w0/7H6m95tk6wdDwhExmKbDm
5sjqy0lgoebPJcahEl3m3LYBaMrtaAuPf9kioSmeHAA8B6ybI3tZgFRYpmthXE03
a9JlDZjfT+u0J1rhb/tdSBenQVpoQHqr2CUGDM3nb7GqCLaesW61gQbG2c9s9NXd
IJmOL9eiXrlZ795vP2BJAaTRwbIJuPZ+9I5VBsO1oJueI95CsLSA4lvzscAnqTod
+9a9u4ZJqcDwFPYFiCTi6kKAFnwk20vVxff+IGZj+rwPNA3Y0Og6YnmbZjYVQivq
kdYQJiTiDpEstJQKB27iWPDHJDNlvscCwsqdbhgJzK5TKUQWxc2MsIHSVVKrjNeR
ViMUbPrsyQ6wPQYSVezS1aSi2TYSzycszcet6ZSH4RQh3QbuNKdJ1Rif4Fh9oYk8
z/++xtEiorjpah8OIPpFqAYWNwUYFrIwR2l+4MKunPgqBpwAs5QyoH6NOLJ439MO
0SOrM5GXt2blb/Z54PUxLz/hRJVr3WokonpydQrpRZ3A5ViKg1TeKMJb/JdLM8eE
lFeB27R01Nhw3WedlDcmWxM72mRKWsIGRh+mHjSufcUh6bTwHKOiZseGencpVkdi
OXL1pzIM3xkIzGQ1iV/xSK6dn/4rDkAzEaGa+iBjy7Gf+E84+vhepHCUwv5wQgzv
fbQenGe9gjtHOT1xCtoesig1P6hMdr6LFbaXeedMFR33UlpmfoM4ll/ZeepOb3eR
fZ6ewEcK3rjfc2BedYqZT1cTWd7ErXGw8twammh1bW225ggvALKl6Z6a95kEg87X
B9nsdC1L+EaDHj77Ey20qwbJ0PXxcOXmnLIhiPQqlvGl75u430o8DBEIpWk10R8j
JmVyY27LTcuwTecfVIX0WUIBSgu17CMtPuhPiw76ct8wrZIWAKhfz5lPOUNgiesq
+9noGSM+/yw4AJ1xcmxJsyc6Bo+xnujGfBtnlRjjf3vAfeAfefuIeMahX1WiIamb
Qm23GffdUKiAZB8HDiW3cYFVKOtQZWipPf9hikaIgezqBQeKICvcsayAsDyTjE0N
pSXSDsjN55w3BA5b12SN4K0PWUEtwOOrA1drpa4ONSkWIs60QVCccVvnL+dpdz7q
jrZ8udjXKEHioGL4FxJ6i3I4rYZz01YTNSlOt0nI1ZWetMXrnNFDuCpMnVFdR/ks
kmH/gizvH/piBTU9L/zwBbubDHfYSu5nQO/duxjGOkdNGMES3gkE5sM0CAIi1ITb
/3v50jjU/OMru+ITIuhQ63UStNqZE+eIYMeuohR9sgWBZJ5f/Awb/L+4g++E3vYO
5Ullq151RnEPxpp22DSQU3fiIpRoeEItSgI4ptkCARN+jZaxnGrPTru25HLcfj3Q
qK1KijKePwvGqwXEpzNZMO3tK+NUDLSq3GdOXkr41K2HAXG6I2ZBeP8IeObsEQCs
iKe/AoSINnbjtuMCyBziAcGtKBrGUeJXuug4nX4XCs2jnHlgv0gQG8uriTjSuttP
cS8g2ebHGJqyO1IoSkmRB4Zawz7oWBsNGM0VxXuPmwyBejTJWiODl1A1B8lzrF1v
nsYzrEox2ThjM3MzL7doAPWCtpk34eZIsrVXRMAaRM1vo1TJ0MIQ1kEnk4pDgQSC
bNzc+4DiC6LDwAuhwVfx6AhAMWZ7sZe1OhDHCWdZN2u4RJypq5m0MBKYFAtSxi33
LedKeI2QF6B//sQQ0s95qSd1lRXzECF3Ns+9AdYunl+o3Hn/Ndk6EolSaFB+nVk9
yp4o3eNGMekV3Ygl2CYUPKu0PX/LD9cas0cMXi2XN8Shq8XCetywUgW1QBSl8PBZ
m+ylQ2MpBoXu9HeaTZoiMIoCTuLw/vGLQrW5c20E7rVMlmSeskCIIeHz86Bp0YFS
5Ov0FHHZ/5a5ok46tF749dv7bT96yjzlbDLpUrNYMZGMwy1LOTFPVEuFD3K1Sv1d
0+faMQwDqdtTDL7tF392IkqUmSjH/2saH7PTb3Gh+c/nBmnXfQGzQ4fVhsyZ6DTg
F0+Ep0r4mqnCK9M0uoo0fIX4BDPtcGNJWahtlS1jBduDgTJq0azDvQLLFCJWKw27
vDN/OYuJmQEWIRSfpMtwzSZke1nG2hkehryklS8Qr7WVAQzv2jN3SKgb8e1zdwZE
aFFAt/ExuCDEHV65/sfqcCz6uhLAAyLv1UDfesv2NHoDuLIFVQuQggjdR+x9nxqq
kAEga+E9pR9nNb8N7BoxaVIeXRlE6eoliTT5m5DiSc9SLvf2/FaAWUd2mzWw4tIP
+OFe2U3Aw2CZpbPbWgRXVqnechR4QnZrIXdTHBpxNrgorHHIV9O5lNrMC5Qq+cTd
5d46RY1q1SxQAdarn73KOc7whbP2MJ92PSAJ0Iu+k4kIgs6p3lrhhOls3L9+X2bF
8I2KkTv4ZdVOZ5uAjdKWVNpy0XMZW0qkpONZbSPq7mVaVTAGRM/TBZDAyHyuT/D3
TLDcRbgSNGN8D3/oMYT/iOszd7Iho7kn4z+A3LBQVeQLsLYjd0iDG6hjoOPbs9t9
BoZAcgPxUYuY2wB4Vz82Qj4gw61b8QEGJLkhqS+VdWb/qJJ3BYcPWdeTFyE1wm62
tQlFnsmxrItsVP6a0q2/QGUP2a9B4QLXD5MdFTFh2C9WOJa5SRcDkMK3EFTuYX60
UwNEbU3QbyH1LIYpUwH9fFXTPym8vPiVQW9JSMhXtFXZS17O89LGU7SpvMCKYk7D
vrqjMA3J6TA9BpYjDdcJERgAHQxrUtS33nXAvi2RDMXQ9B56grP98gwuBTKaww09
SYBJNwEAUMHHFwzCOSXQwteCULurj0JXIrQ3asmgCDgBJUvjkP3X1zujg9qQfd4m
uIugQfR/RVqORKYA5aDlerWtEdlpbl1SYz5YzBoM7tB84VNDhyxKr25EL1XuBzF/
v8iYDbbVMb2CaD4T2lqv3sFh5RbAVhfwX5ws65Wmcdj6nSCIsPBEf4DAee11UFEA
iOpJKI56JNeMxShdjytpADDzmYair2+qkgAA4z/ALWcL/x2rpob0vW4uH/XKGZkN
2f4sNeGSlzbGk3YMfgCU0V7cJfXPSbBsfd1FdbTqGXfl1PSLVxL5tAcnYVq0yP49
WuJaH/zut7jHuvIvy8+DmD5V8d6waxmqp9M5anXb8sra2eCsawg32jgP9Jomyowp
k63fXwe18Ad3vWA3lV1xCDqWDVtUhPcUETeuaPZ7zLbJDnj3WGOg43ZP3fzYbfqi
XGJ9bGO+0lDciSzPM+O3G4M5zSswbHv5c2OFuAIC7Lhbs186zp7uYIHyZCBTwWt8
gZpH7R+HaMt7GY2pHywwA+MkMGdjsn3UpiSnjZMtA7psRvbg5nPDZ0hr3kJgBMwh
xLVSK29dk1EMrO8uD5M64TVYqQv/lc6Y1VRbuHX5NXkHzOfTAPgZOBAK2mUryyoS
ujaI7VIryqnMz+tvhuwYZAg5z/vLCdA9aqcHx7cpTdA3sUwqdwn+7w19rhx9cQeL
H4bngd7UBHDQT0zzoYdeBODS7UDrTnb5cSZLGptE7D9Xv1U/RyHdx+WiZKwT45RM
SJiZ+dxLzeqxHS8SmEMXrr8fgT1Sx3WqjOIE8XeQzMDqy2oaIL6TsOJ5Ybu2gLbU
JaLP2L+nD8f/yDIy5y1+UaDXwWxL49Yebd7ZgTAtSfX58x+V+psDR2QNP6JmSS1N
q0Hj5PsFNxAo1K5Y1VqXdlUbTR7qjZIiKaWohTHBibUzjiW7kpK3eQR0V4d6TGf8
puSrditJtVmVVT642grsr9jJ9yfNIKCVRnjcLGmmmPBVXRIIAZ0rOL5CGi1QVwSI
H4VweCXNpVK+4DLK6BVLz6c6pjWBRxVMK0ieZBjpANmxK+SZ8YmfPW7rGNxRKWtG
2hw9r0v0qOVjF01TBQjjK3iWbH+LxN1Axfkn4fLuRy+2YFJk/BapytgYJJJ6vRHP
afhdbDT4zWxzbI/FBSJYh2UOTEizvlNkdoLG8/iTiJYoUnNrIOtL3FQ3IShTeOMu
J7UuD3laN9L748ZXiprOJ6fSe4t7hHFEHpxwOAhuaA/iafhgJ8hWKAesrNVlrztl
ljBRgho+OmwMHirMBamAycBCz9wb8+HDkYcA3GXuH3wGTF65UC7q82A2mYmtGyG6
OmVA9FzCd9LVCQNQuZWuH4xzENaF9Lx8lC0pVtWXhunawudLwhvwqytaCo+4SAQB
b2mZN/A5WBuW5TN4DkTRl0xx8keK1ShLauJ6Knoz88or9qDDNHURaw+KFCDecT89
WHFYENQ8rJfcXwnG0YYEnccJDU8X19bbPnvi6da5rwN/wCtNBoQrG0zHwhPwh9W1
2F5zSHhIu7vUNp14jN48UUXeq29/u4MihF1Bt/mxFuH0FjGrqluMWKAl8CNb5m1y
I+P8haBdT4ZywdHn2XxagmmYHzvtZuGanHYo5FC+GbxuTKFTfBfuB/NX10KnNMVv
yHkn2fa/a3xt+hx+XoL1bE1af6NtrElnkcSOM1j6gqpv4jDNyHDwOo4SIZTZtlUb
6Coz7y01lwxCLQPZzX1xU7fma/DZDhYlwDv94aalaolTfMcRsF/GWqAOdXMeZLLU
3nszfXAy5moXLXWzmojLkRehOVOfPJlTL0CUYtIBHlpE5O9MgM2eNVojv32Q2FVw
SkziXcgk31WyIZinBNXPLLqTEPGewMMdN7zez/VBVL+ViA4wHWQX/tenFtlrmgwW
JjGQvyC/mwfB++f4Jf4hUZeEo+/9K6ZlDXkjJGHI9/d3hrQdGiiN47C1NiVHSMqT
hLFnUpfQrawSP1XZVh63W8vfH4Ow6XydkUvCcz1X0evsLKIoV/f4d9c9EDLmcKxk
3IEHmaPVuykPUEB0KlkdSzkE64ASv8R3BGIWSD5oeccaIcTQ77uNXKUyww5sdMS7
tBFZRRWerKvnBN49JDADfLN+6rPJhTKOoV+WP3Hc2wbsjH/B3uhjFy5o5t/B9Urr
ppq/2utwOfbRpUPyTUoG3dSERdUFy3u+4zPbii+YtGJSFe0lH9YK39RwriKp5yQG
pqiSpLwibncV33b7X9RBouB2TNJdUZpDD9sJTSw7J7dfetWSocLeU1CoqAT6a5mC
Dob66Qji41QSrDiKMWEkgOFKlcCXf0dBvjKe3ojPEypr+CMmFNpnmc+QiVm19vK7
PsHG0jr50UJO51U2pq8e/RUTle1DT4070jL0grXIXClLYz1Ji83OX0GmSD/3LSVm
xuWxuipcI+CgQ5+gT2rTH3z/MqNN9WZZO+cWYSStp0ztOqiWhSsyg7BnfFt5C0Cl
8fVlvN/v9Eia7Ez8R4+o1XGuZdRBTJAO0PytWU3LGogQarJEkM4OpM3bqkY467nj
zjmZsC1dbZWwNGz1RIiuvjaj3brQthTSXiVgPjQZK8kMxxYq10k2Zu9lvZRQDmKi
EdYZlkxZlGMRgc0nwxbqiPlyj4Hnun604arHxvZXDxrFz7dFHcVPt/51XZGAS9Aq
+XuxLFcOeXBCHoGVS1yyjsi7Z9X7KNdkB55k0e41zg8pEJxQfKSe6Gn2Z/lz8UUT
mnRazXIWp+fAGRvnbF/P/h6K5MRo3PblxeAd5fNOoDBzwbXF0IDvKcb3/wOmOJs/
euWQHbdHXT0qAK8NRd/HYvk1v33grQWCgxbgYaDzB7ZTw+4+4LPVgtcsxpvw8B0N
xXU6Mh9p4C7NWKosMW5PR+lXkiahLhrcAtoYtl6sZNjfqRd6MWdq9+06fEURIqzQ
AibrWdEDvLbuihGvfFNU0QMlzblY4zklDhuCFxZ//yWnWh2ZGLScwNjYDZsIKLxm
GIgYsmw+izrRrSiI/L7v4xi/OAmmtZrz9uJFL7NNVH1qk/GPhgeAolFAiVjqQFkJ
EDkeJJfjL1tHC8UW9RPY0YwuABWRslQs/afJ2rHRzUdUtXIxbRtr1glliwjmg4mB
+8aAu2dQZoSoUg2Ntc23zS/7KKmFhIgzq/gJj19k1/kdSjOymeps8a9UxObcEv6x
sZ7Z4ZH3JWAsxjVR6129YbcTPzmmmPt6GBFeHkWxFldQmPon3f/grH753UTuoqDe
xV5024ffOsX0maFO4NMmf6PCvNm54hyllBzTyFfAyTKiw6Km3BriEUnT0Qxk3m0y
eOjEeQIyxwdA0brhG5WbDR/pE6zeWMvNGAmGmwUZYVKkybSuYCCADOJBErFifSoH
sv1ze1tLaMWtvXGL8JpaG0BDkuT/k2D6l2qoL5MtWGKbaTNW/hl0mi4rwrMHKJqJ
1U0WWm3eje75KhksUMadQJa+J28k0GW1OeMvMVL9BvSe0aaSdQBm1CU6ISPW+Z6q
0LpgGuzPimq7oDYjcfnAAJP80oepQ9iIKn73/dS/1RDd1c96sRfYqy38u+n5nDfJ
xiXm6TptTyTKQyU/siBWRz4a+vHsH2cf1xOngYCe6iIT1lEsGL/BltI2jkGHK1JC
tl8viKvVx4IKsoEH0JAou+pwX95stxI14xQfgwxP9r1KP2LTWYyj8KgyBQvkkMci
ctt3YDB2jnxrSkR/QwMNz+swZacXX9A6o2/dZn0nvZjADSUtRmx1VTlYMyaOlVrS
3zn3CxwJH34bpyz2VAjlZnWhKNJFvN+HIn5pPOWr7+zkwfG6gaMUHWiSj6dfJTLq
oItxKvbPN/U3A+GY+wW7mjsWL42PFdVWiJynqDchKlEP1+KZd6PujKVncdWRVnxv
a7nU2976qIEOmfOdVjdKHKyJM24HV829fXK+gHsrLipD5w472+eTRdDl0onOd0y+
x4XoOeFhnbjk9Uv7JBEFdrHqDOpJczdQUWgbbZxlunAYAwf+yN0HyqrF5Gof1VJO
gSoplkvLAMztgZtkAYyAWU5Tm8iX4JYEYHxZ8W93Dklz7hPJddyxdyOhjnn9Lw3j
PSX/rKMuYjyYnp0cYywNRab6L9LLtGzkyB8MLA34IoUVtnifrw8D7T2G6Tmtdo/5
Ql6N8oe69c7QD1mcjnOSWg8VHR4bqZewODrgw5qc7cikHhMb/Wap4Bxqt7L5P3dY
O2jLyDRVc10jIbP7c93hMZnFEQiZpVKrRloLgFTblHzQDsNt/Cmed0ate5OnvDnr
nZTHmoXmcC6S9TfMyNOC/cnUtW4rCRKQNcE2rNSDbrP8d7wLWgfkSf1/GEzrK9zm
APvvnddD6ylvkNLR9V+ZlqSllIVZVKTVS85eUf2NJgTEZhaCsSqSn6WWwwevUwcI
Tol7lXrBovE4DzeVkdlUZtbd7YHTQ0mgK6k+yjFAJnWAemv6tCfi70hfOjxzdYnN
55A7Y6I9e2vW5Us3TSVjIMr1NG48ZkASRX1dLusECAI61q/Uk5OcnKhpijfcyPX4
5MkILRF4UkszhvUAv2Mq707mpBZ9GCAkHFjCzC1yxogHrf3WEHpzCnD+Vg6xIDjq
GUJ7EvBS/F22MxCGmRoe1hLqWhHqHPKcg+2P43DsjLvEytQbF+9TqnTId8hQxcZ7
uH0idAnIbZoez6VWIvV49Ll2rfb/+mbB0jqyPkKT7CfzSM477qaj+U++gnEH5kyf
jEqKqCu3Y+HVsAr2u0cvay8liqxAuBChZ3AH01mvqf7M1MKlnqVcGr3ancjLZcch
oCDsd/V+wi/qwBGDIAATivXGTkO11MAbGM453BEsohGet8hvGnzFjUHTKKk+/tkJ
4Si0m7qCSgHcpNqt+nBcqTyeXcfbzssGYv6uaJGQCKdMY1WLGzKBrgxnb8M/lmos
D46irujU4PoDCbpcxnmHohMPXcAfsuRVyaKL9sSQPqHeDoMRNTnKMryD3DXi8U0s
8maON2gTCgFTfmHYP91zOnEyDSXUlSQzcFIXiGMPounmAeYNBKDPNHN0MxEjs4jp
hj3uaoaPb3S/cwc/XqTgf3LGxju7vsizmJSmG+KpcWlvZZphDDkb7uKeen9/xcBl
1VI/aNCLmyIbiOZxuozchgHM4D3lMHhfmTQCoVM3i2maRez97cPg0M3BnLymKYF8
wYP6QvW3Is5FnQkFE8fyhYEJl0pq9zkFkesF8/5rGC6TIjWf2NfKNR6NS9u2potK
WQ0EQ2AaipsGRN0bugJYoTZr1N/muz+/hpsFBEFgRYH0OPzcMN3gB91IJ9HKInf1
JaIeMFj+kwDSVxzgskFU5YrHkVvNRbwndXIVsY8uUg+670DwGK6L+I/R6Yh36DdB
QkjtSQJofKsrbHgtub/l6y8O5Wm3bFBqs1tSRxP+mmSr+m7RiELTi0BK1gIjLZi+
bQoN04R7qwJ7gsUFDxXxrszbTfTjFPkt4wdgZTy90fKQIIQjWMVWwxXeBlsTHU5m
tlj++TZoNz6+1PpIoFtpe4kMZHY2acVHZyOWC7O/sdDQc1o7g6+LS7bhmG2UOvuN
XvYsiCUJSq/EOwxAp4QZhV1Nq136cuEgY8wfQORdyL0PgkIDsrxZGaHBcSbCOMpS
av0W3lvMDcYzSD2FuQjo58NbKxZQAovzI8HKoETCvMoNcl4/6NjoTR5eouwNssgv
KRQMCDQbEFD2IdQXVMpo5ZJEhsJJc9YBYJb7mfYC4SDw4Rzl0H0N8egA3vEMuyEA
IXrzx1xXVdumBRAUTxVM80LswGRIhlcq7VY3mQ7Fgy0ON+CAFzUGZ+c81u3BERhW
HYLgeknMNmIfcF2jSLrRsJDDixV/Ez+mQG1aG+3HJMhOnOAdxJhjSpw21UO1IweY
N4eWjzHqabdPpZ4EQpJLjpxhw583yX65ztDUOdVP4KeYltXUccP16zTgqwFHNevZ
W1mD+6UHy0aFQ5XNWgsFllWueiqbhm3Uy30O2eHnBKrUKEzCAxo6btOFl9iJiE9a
+xcrlngHeW/4A1NnOqsNKSHgMAIPOEZlnKO/Oezjte9F6GE1dYKH8wwJ7YsxYeWn
j4IuFjdeNpA++SM2jWZ9AgSQqjtrctKg4xW8H1UWRAxtyMZe5+EREViB+XHHAhMw
LMuGbTtyTMGPELE8AJcZtSh+qq7A2G912AALwQTND48UgoAwwflGK5CVayKkNB+v
YWbeBrbwG8rDvs0l638lz7vyrG71pJqKpesx7ApYVsqd9CHdPa4yRqrsbAX09JAM
gbPw/cUrbcqeFwqBy40Qb0qRuwg0FfD2HKpGI5my94gaxNk68SQrlZPXtP8g0UJa
nl0mjOeahAAmE+vxiyjKG22orMLVpmzPAum6TdCGXZYWsNICcPDDZNUx5sDmwIci
vMV08mvXiEBS5whduUurns4YKOt9W9duqG7vvqoFwpGAxZwq21GSvbB6rQSXG1XN
4yf+Tj2vqvSSRyrQASHLumgvLfmKXcHlcdoqe4/7MuLSuu3FNM/thcLBuwjvODZf
Xqx0aNXTYXoefWkznMxRdJmvXxzQ+fjHvW3DlVZ8y9qbyO29R0n5zMj+fIkgmbjX
jnxC7k1SlaIGcvAgqlxWfyNdY3ghnIHdzoxZstKeIrqcAfCFb1bBKAffxfVerz1m
wTXRn+9qWXTYvPAn6NQ2s9i5POmTHoQq3yQCPiIEJ7y7h83MGjLUfbPWe3rY+FVA
mC/rzqUSR/O6QichNKP4PSlNM85+HOTnL8BEgI80yn7gii5f/sWErZjd72SNUFcn
w6BEdsQz400KsGCNqc/JnXcZBb0oXRh8RsrvKA7leAZY9sYK6WXgxTSyRtKeEXM8
Rz8+iOP7V1WCbSMVsGnSK1zpUW+5ujLde2IrhOQhT4jELB7bfs0VubxiueGu2V0s
/kBJ8aKvcoGmFDX7A/remDvUv+rNb53+HzDdZsNjZ/9pVwPwESKHc18kqj+tpLyA
vOk02/u5xpwg1l3eySM7xfaxQZouxwuMWVeMYbR4HhPJZAO4AXg0BM/j5FYS/KOz
2J+K6zqAT95X+LEjcmvpzslg+/GnZJHAYX9PDuBYSXuurrQQ4NyzQW8JlXHjfdKo
++JfE/8yyMFH0qdXTCJgxqAebMqojobzOIb5sOxIx9mzFzqhNvNFYRmbnPITbROM
CsTjq0FBlNwCpVW4lAoOIKolRQXoa0DjM843QmFwQ8UMAcRihL1tAXN9trY2uRob
Y1yWw1XlIfH64jcgpW+vehW6H8CvVWbx662oRYvSYOHpa2vZgsued1UlT3ezy2Ck
UT4rhwztAiMahq5bKggJ+wGTvNJ3W3xvXEFX6P8405J4AuwOh1J5EIjkm9wRXU2P
ZKtnm0+t2NgfJMI44CNyxLayzkoBQxb5Zep1iMfrgGyPb9i4Uv9kJrRJHMEvCcJZ
6h2+e4UpqZfq/DipxD7TYXz4wiX+ir3TRahDc2DaY4+JrtTNjbvlcdrvR0j2kN/P
HQDICa6VYOGItJ887ZiiKnIFpohQASBp4lXhCeuIocO/zc6/fF0RQQgHjIVhzWSJ
9WpxrgojKvFou6h3M1bwA7qUv59EWEeeAmGj/PzaM0iMKQWzqk7cT/N5dOgFuEE8
5gZXrsbDFoju4V0/h13i7XvUiOwF+uis5j42PSgiNfuJzYTyxIizHclriUvcwF3l
/yBLSuNculhTMzkR5M8/vXAgiuLhJq+VgPsmkAxUQWjB41/DGifQvumeZp9OT/LW
YGSemIb+3vgyE2rI9kHgvfXbJRhKa4i6RtGCM5u4jHPRGElQ96vt1RjhERiP2Rn5
5/e+UTe3bC7vgAzKFtEQDdsueHG9kVsJezvA6FL8I0nETOoR1wSBV67J54qC3Rke
wUXAKVTTehClsB2GQWWEQFf7sMROEyXiINgZpJKncnX+L+Wpb69AsJlflfHn/eiX
JH4CJIkz+UnETuZ6Ml3TmUHZancQjj9jYf8rx9d1h7BFu6GQkHd3lhudQtM5RhrM
A9ySd2A5/OhbBI1fc6PUNbtszA6D02d22Vl1qBtJz4RFem5sp7/MsSimqPf8gxD2
XDggqUB+7rMOhjmx8awhF4G6BDqQld6JEZCTgLZHcHwaPzZPiSS3Z2y7YobGZUcX
xOh+3vbcLMLjvR1zRXU6PoCqr4ozHJYxCI/yvAWTR5bav9D54sSRbdyq4Y/I5OdL
q/cuUUzPH6P417Qk6MN1CS3TqN8zxnLnGJXtCy1mDGru/Vow4EZy37zbpZT/kP6Q
dERsn7fHySbJgctNu2H4iCcd4yJ5ShRm4VavI8GSmlH8yCMSvyFVTaDJDt6dhEC4
Vv2d3YTjBXP3gTXeJvX7qmG2LTE0GaxKlQjZwenQMq2TUoOZ+BNTyCFeErvM60GV
XNgcAURze6qkT63hxbljsRaaDHWpQ9bz2YgkmmDU4zFkqPkDi54otaHhBzQ1pQSD
7FzSPwzP8PdDh/BA9/nnErOVQiVrhSKWe4IhJa2zkm5VI+w1l1UUvNU7DjM2QvTu
RHR27b5iOYC8JspYVkhm+iC9IFAP86tCx2iIlXAhMVKsFGrxRbxcGoWblsahGuc6
DWsuGRhm/wiREP/vHeimp3qqinfirWMohjuv6qemZBXeEAqCBvSk57fyI2DP0sup
rf6e+Pf67F5m+0YRoU0aE0xbp/mnTt0F+ZEQ5Nj1FAkIYkSWtpQjqunp4cyY8WtK
hny99YKzhSwcdItUwyB6BtHVJws4AfHj451d/2mvqvD0fzTVVqUpjKbT0RB6jQXU
3ktynvidUVQlao4HtbBHo5zyZEVhiaVgixoAx+U65F1QKYMgphX2lO8nDzzn9P5S
6CnPLucU9V8C2fEczkNRTNOTzJ0l4L0zK3BQ0vQr7wokYUD7bgYsXCIw1NgzUmkx
cinhDqA2aDH+UwvSZ8iS+LHiagZlY8JZOx5Nmo6L+enLh+Du2yAjYKKcHpDrJfat
YZGAlKN/damyYvl8cuTROI0eTezu6CPybNBgVFkmz4uAP6GY1f/tZBTsWdpyE03U
J3XRRAQuZvwrkJKbTDbljtWorVn/C6WVYShKSm/NPQGp5owrinoeX4soMkhfWEwI
Wk7WaVdyV+wMZZT0Y+CUTk0ircMp5af2yoFq7UsIA5mG6taxSZjM+VBUbXT16rsM
PayeCCi8JC6o8L27i8j3GWlXLgdUGljbyiZVin2TapfXAdF8vm2uBfuPSth6Z9Kd
d0K1/E+2yyNCQnVfxBTcjJ1flntEKcoMpR6PgfqaSkFT4AZqyumcLE7R4ACW3hKl
gxn+9MRePfKL+3JwlT1iCEBYj5qbtIRmi4Ted8sKFziQIeRaM3xWqFdTtAL9PiGR
4zkvyFx9gVOGr7BdAEHhO/4KNbTlih3Iy/8TP97JLlaP5A91KWD2sG4n8swDNOVA
YzJuhxb8H/2mMLsNGsYs4hD201GfIH9i9UL/qgOJLHZnvLwaHv41gUYnqD3io5Kp
Gt1CdljkoR02zI7K8NUe7VwSjhOemHvhMeBSFNb9yjCJTXo/ER9oVq62gKr021zA
VVxH/e3aggv1tkv8TL1EX/NH/rEjGKwSWSkcpokDCct5x4/XYsI3aCTZU1FLJSBj
ivrfoTuCTql/5nTMygg0dQfs5qkS1iO/QfdqDdWbnJ4rtlnJ17E7RbzkWkEHwXD5
nT6LCCBcj2rJKxvahQtzmU506MzJoerO3x7pe6lPdAtu5A89LaSOAsIx6QAejf4f
RjHgrs0x87OYdUYtK4IjV145G/82a6+U18fg06GXpy4muE4LHejykXmV8nk1JeBk
98M6/MOL0colifVotFOGmP664yoXEomHM+hEAwqA14nmh264ePClL8c2NuCOhy2e
7v+/xEe3w2B53a7Egts81+SbjvH3kEhC4MyOk2jd8FGsF4xBu18NTByZ9r8cCKON
PG5Ti69ZAuB/5fzdy0Nus9w2H7IvATzRRTDJfQnACEIbee5TtVOVwAi3ucK2kesc
/rdcqBxAgjGUw7P7s9iUPRev+tOC+PnVdTJotXGX1duVgD6cq5jHsyCIvWXs9ucl
bc20ig6xGjhkr5inOErFjwkMj2x3elX8+3AoRnggm5JfOIzK5ei3hRhv/xeTcm45
ugpFPb68sZyupWWvDg4zcW9+ndh3sOUV6PPyOieCZYuQMTOPpNoHJFL4K6hUXiY4
GPK8B6I9lubcZd3+jaOIkht5C578+arE+xWtJZHoGP4EotKo6vPXVwJXLgzclMPJ
yvYPGSVXGXV/W4IS545FGUs7N8G2dLDPoT00hbdz3vvhsDCQU33lQVbrQjWHLQmW
W6J6mfPZOOW82vSeMa/gn5V1mTCz33/mzCW5ynH25oRkuGwPUnLCHuO49yPPRpgu
QKxn8kGQjW6dhmwEmY57DcyVR7b0/dUrZtHXfZHgw/dvzo5PjnKO2w66ZXPVrAWZ
ab3RUU3di28V00FUyutOav/+Sk2SqGX/58IcH0rDH5gP1Lwvco63oxkpJJnqmW41
V2XOIySEDono0l8igs6SH00ie8IHGeH54ijf/qXkXBO5J2RO6mz41r/nymYFttXr
83ZUTxmGhrQanIKCw9YTBwnN32cl7pDtv93htxB4L1M36hcGWzOW2UwQGnwZPd1g
+kYGrHm6x0GAZjhS8NP/Opn42lzD1L6FxQJGNMBp4afLerh4kdcHPQVA61mpc2k4
/cwHCkOziD+lmPaelxSAX8G3eyjxOlFDbNQvINsNv9E2t9GIjaZCMXkGaEYr2Xje
w5+YqVxXumf8yaSD8BGV5CQKORSxYPdKusxxQCbRbrWLaXmNBYLaIAgan9NUbooO
JDzl97+UtTjXSUuvgkpXNyvCBPbolaYM/tz9tNCrm5O2VvXuUpKA2zyZLkgddiKo
d9QshpvkpKtL/WJbZx4LPIS0QmgVuk+imy39RsQLdKX5WSc8Lxukczyjgf9ZZi3k
WRof3RrK+fexQe0vnFH/4XejCnkLiI4Gs6sG/lfy9MP59RucCbCeybKZmdAnEKMF
i5khx3/jgpWD8VtloHmaE8WyRIwmiMUOGvGj0IK1b8XJxRvVWmW7cUnYU8DohTiZ
z7M7wH5RtEK57+QVj7XwfMla2q5qyWlBTHzWERgkbBsBXJJmtIJL43RnC+ut13ZV
uLsXkO36i/4TcXtoP8sa9Omfe5PaPupT8ftLB7zQELaHOEVx2pZMxVYfSlnEiTd6
t3uJbuJDE4ER7lUcaJZY5lC2VQPYhleuUR52JVKKeuicZYmredWeFqHOieyVgke7
ArTf1Tgj5xVS8oySk0UK1EW45jnj8zlCfe1vYTSPcj4ksR+/rv0sGJg9ZrhHmOGt
/rde1NQO6ywjXRXSYRqn1WETiAZDDRnUkTCQ7jo8Q5iLRp0Gc6EjX09HIF+TYIwg
fU/9KUEmmbFMCtTchRYwbqojcEsMETXL9OZB2vfvodNPT8bXVSbECfMwmhNWLV2j
CXg3SY2cXQs6C7Q7ayHZeb2lGlDpDZJvVd1iJCc7MQt6OJWIuSMJRX4qo2OygdfB
H5R8N5QDvuiWqgOjRwm6mrKm8ZStTbNYyj40hXNqsde3hQUWH1wcA62w0pG0wRuE
TFHsDojFvjnF2PlJZtHHJlkJs0sxgWH3vM9kMjRwrk/qR4NtdE/Qf0Qteo/9zFdo
BqEfPS3UOIKQ3EzR0YOZtBHY8hK1QEl1oSX8blB/tabeafvxnPKPqUGFrFLINsqv
78X2jCyRJx3auS59YuMd836pbrT+USsEgz4Qz+HCN1eYhIH2Ari1OcptF22XegeT
RYU7YJFcFVcLGiTxKdLg4aWdjkPlLCOfoZWbPiO7sIhs47kQ+woNoKrcLnCNwXrO
CMiZl4+Iyf4uNm/uufJR9/Z/RfTA+H5Uh/QH7GkFZIMCX7XmBfIhtj0LocUd0TZd
gZXpl0n0XXJEUdMQx4sela38Oe1v/GhwgW9WucFK67g1qGHzzw4qsLE7od8Iw6Kh
kXXVS7ThYZ1it5xSM6VIxkykv8AMqvY/cGI6M4FfJmD+BuAa8hbMoZnTchF4qEE1
lRFPjtcu6tGPIypm8vveBbswcaaA8a/uUQiRiwE2yI/0/SJsrc5WtRc2nkkf5IPm
Zp22dsbHpwYmSD/UazliIUz1aKynFgMKBV0p2UoPR0IC9miBPp7gcV54ipZZxl3Z
9bp2pajmV4C09exzFlXwCEHzJqvn2LCGKLCXahGqRFjPVA57z8XqyABwzDN9cpt0
f72wdfEcxjbKFm3+T2fGCIhjV1IuH956CBBhGH9Kdgmq4q1lxOLZozbhfZILjqK1
Hgk8N9fb5aOwwPOQYYw81ZOiSR2Q0tbGGWZrDJBBbVX3BM5+RfhUryLfERbs0ObC
pknAFR6YUjlxPkc/Bk2GJ8dlWa8fIrOw35Lv7N6smpL/kkDJ6K6Mok9PwiTNUxj1
AY6yLgKeAkJ2K+eRu8KnCKZ+Wr3TtM4L9kcbcpUDjWmaWXZSEEYn1d+n6JeTY3j7
UsznNljP7E9EOBKKkPl8pGXvBNz43IVYA6vQ0eoDj5xW8l9ETha0iPgVFHiaulxj
t8vd8ucsUiSv2VGjwToyCibSBtHM+6IvIUuBxp2D/hrQwP5CH6YZmP/FtbFOugAc
EFdbe1UZKm+dDAqG12SciowWmcquFHyBKbulmv9Fu6LxYh6L/F9MIahonv+xWOOv
KfyINfwdnWsvGSnEOP/WUtBKi7t/qqtOiPVkKzK3fo+RdaAysNvXhs1T9vf33ack
QZUjLqs+o7U7pKbAJKdyEGKzaMJAYn/jXM7g9t7PK7Z31u1MacrD5Iy7Pvl1m8pN
hx5ByfEGlKWdHNccntm2lhYokDXC6vTgcwX9jToe1cx33vw6A/6j4c4W4k9cQTE1
/E/KLcm0qHrw0eYaog6NisKG+B15EjOFLGMed07N70OgrcKDE2JZ78WtHkTS6aMW
rxt90QcUXUirvaTGQx/1AmYjMtIm3uu6X7io350zQ17y3c+Sa2maFvs73rSniKL3
ohVmrwaYetfYzW38S3ofOPohSKbqalFedw1YEIPVsdKRoLCuZitq3whxszqsQJ0v
pZUqtiNrKQTGq0NuxBcbkDrmSQL+02iWv/oxDUV2aujuW4UloshIzsOHLf1gSQY0
rx4tQCJX7lvvhkNVYtlJJ3WjKWNUdlo81z5527or7jQWyNOXnfLs0Y+nfAx7KB7X
EC8r996REifh1kBdDFjSVci4aRvQjn9ICGl4fLusJILhjkTIeE844OhneFtvEVqP
+WGMjnQAagToqc4QrBJeZ4SJQRzEsZ3Mx69iGHZ+MNPjZxxU4fUqJiIH2xCAhaDX
IsQZzchJYbTqpwc+AkTtxn1+xb5dqA7cJLsbKnZ3nnj+aOHIHB2B5fjwpUGNjGVN
+b6V0uFMLRl3snOdGozm/yJ+8fE8DKHSqpHSvbL1TVeg1YMo2sLLMdy9SnC8/pz+
6OwDHlxXq5k6l0OkpupDmDS6ZkYMc7mYYwbrizQWwEli1mpZSXm4WUa1bRIn6Kpc
DNHprIZxe2x/vuwkewH4fgl2UTcPuN8xjV+IvDvtAHmk+XRm42ogsVpSba/aq+FA
0kGAmVRhZtmSSARapWBRHCFCPCxA9WihMWGjUsSnjnm0T4KPSCdR/Mg0eJDhYSYw
nkMR6T8h57IJaE4QQ2V3nurIUp3Kv0EpxkqqGDkAE465r/V0ec02HCFZmY0OZ1lB
c8m8v9bX7aScxCmTYZTlpsfj0VD00wJ46zgUyDjcBlsvR7iwe8wB2jcwhf2r1dKF
KuIHrn8Itk0dnMe/8vXymG4c8h6vG9wp0cxvnpDpzBucJs8eGLsZW52illpS+1O0
d2ifeNZANq5HR+acYd8tb19KXSoh7prJc3LOaylr+mCoabm1soIDCEs5VZc8y0bH
LvfOG4IE4iAugvIw7kALdVLOO2GeEDVuDf0UtnOePRHvVkxCTbIhiJxxzTw+UH32
0mWTlMrwp4IOTocq74hKGJRtmB8s3zJ+gBb65+GBisWYxF66YnWvRce8Y73woNW0
Nm7bgy3W1GLJYIEQxnccgGu496sVn/5Yl4LKXehv7KZgGKpLtogx/mHOY4bXbw4p
7fo+eczZl0VRlicxDLXmrM9OU5IF16WqqWsJUncWps2bDpaG91LkcquhgZxhGubR
0hXOX7egVoTAUeCtEEJTT2nHR7EFXS3ZNTJbxedtOG0Oa9VxqaMKrx7qk12Gd0yg
Z/ji1YeYH4yHbU4E0ly/zvIefRJbz3JsqvugO7JlbF1dkifEJbvuduyOSINbA8Cb
9LlfG12TbaZGS6TGoFA+gOQKGCmKHIAI5wcyUXBywoa0YRM3voQmF5YpblbBli2S
BFvj1oS3xPY0Mfe+PdfM1ux1opYWTmLRKlM61zIW2CQ9U18ScECQO7liv9vIOWeP
nBbzL8Ye+6Nm2378f8kMfvz3IOGnG9MExJp3g37ISFKESEDvQ/G7QNEYlV26mP7S
dU62MstAtNih1ydHW0u4BqByEujOzZhAOy4gQDV40PBlCAexAoguF13VLt8qqgBK
604sO//TSPtPoan/IAZvUVmw1B6dF4BVlmIWPvwi+CwY7tHeyAdMGjb2/HSm3J0U
MhPrVwZkitB25jXeE94jCZVHJDLabBQXcsntUFAIe3bm6JowmH8ipGuqrG+Vsuxs
muX18/1bDTj4XvkuzvfiP9g+09tesGiXhF9m768q4jvjl2xlq8uTu0aKu1csgskj
75usz7wO7V32BLHVwyF13lTXT2tiqNRdEzGmYe4Ok87JDJBOHQejP+kJlk1gL9n0
rLKQOuSk1E4clR/8BKHQvHD+tCEkIYyxwOpI6tQpRn+NKp+6M+EjyKgtwER7qzob
ufA+WOjKUNHCHQuJboWHEOdETJKbiHehrRMNbrRH3r5Q9pB2plwyFDVIu8sxWy6B
By8tPOlN+WCD2IS2hKKz9CSHlH2MFhU5dyslUajRsODRKeuHTBzaEcM2TX2y55C5
B/iY6A29A6Ob8prz+l95DPzcnOV9EO4JeCrltENw74RGgObXh5nMN1DcTMobK//+
kTdnR4SID+G62nAB/FBSlpp4T8ko5K23RsjWPDvjd+luYIYTcjRpxR7R/FTHJa8e
K+yBIA6RN3t7liDFH5zsDuqWXcta1lCBrVyXL49BFJQHHY3xwy2nJKNWmmHIJXJC
6wgaMJ6o6WhT+evEh/gfUPT3RWv7xHEsWQRpyvF84EqywIsB/lYzwn2kkUW49PR/
QwcNUvBsyXSYuCMttlbrWX5NSW2ItD/oXF1xtVJTIXH4wBr+eN3ZEMmpPu/7raVN
uYMB4pg66rlGTiBZJOK5YotrINqzOuZuqoq5ayFAxcQFYf5j0n2X/t5XHxaExT8k
FFihcaaS2G1TVruCE9DnPgSP5ogvSNDbf+BQNdLuAZmaGzxT323oV7huPu3F3Jzv
ZT31VyHLARs6espsLftlFgHQlzYM+GmweTKa3FQqrYWnSyo2aqgfRnwpKcaS6ANw
xpc9mVG9sGuXSP+cubMkLKHnMUTOPdf3mE7wYixyCOM0NIQi0nDm+U2HD8ZblSKP
nVMTuu5WfuXiZhCmWAehgxdj81yq+7+vCiCbXnabPwd+A0zsSzg3fsXq8MAJtS+K
Q9tlt7bqwfF5C+zhzzStK9+1rOafXv/DcjjE7+vhklXpXrkAd9EbU6upRNuKbh8S
M9qDc6WmwxAV68OcYzXx2sGVE7tX0EdR4UTVp2RbFhssATXqGdPSI1fKtEAncKfs
hDPp6AaMkKEQZ9CgxE/zek/pNuwEGb5YlgwUa3/ZHL0w5uXaa3gnd7NvcJXXcCJD
hbNgq86VBDO4wqujZHIPzF7rwpNK1MHt39lXLDIKmAIoVmhjh2tzSh0wZ3bdReIc
GDDFbRmG+LrThNzs2c8kB/sbTxaVEOkNYSQb2C0bcFVniBqTMi61FY+psyRgUMRG
0/dHY8mQSGvh2Qe7wTv/wVYL1QVDeKT0L/JBtRK+XoQ2i7+sh2QVijbaSB9ssWRs
rgPqb48DVuR+z8Tw3mIoF1akDrSrqPiBJnFlf7dmeUR5122DxPHl0hT8tRb3DZku
hNSNfhESQjl45/brMc37rK9IO/m6lE6z7bA97CrPS+8QFh1lpAR1mJYtA0DIn0XL
UBUTnxOlDaW6FWzC8byF0o1tnm1zChCUeEyFiclBND/ZaXE5i8vXa7wJxRL7oAuc
43GIp3qVOSbPYuEyaXizyJusJ4hyJFbRHixgqBWcd9M5RS+Ri0pJnkumlWz3QWFu
+EOH/4AEx/iLPGjT9zJXUEBjva9WWUhRGqE9Wx/ukdjLdvxCBevgTp7JaWLJAryL
ZUX6xNSjMjd/lovhzoaNK9HBwvCn+2S7Tme+ZnivGkZ8Ia/Ij1nfe0j96F1r1ddI
g9kQ1uLN/ofM9L3vDf+Ocx1bgKSbhg+1i1vh0MY5ykZaJlgnZ/ZP9qSVuJHPVgp3
82VQ4zO5qK6BaemB36zrH/EQN/p7AbBw3/XxydXX4iAjnopKusULhWMzMHBZ41QO
kLkav3aRF8GsRUHkLeRIB8vu+hEP3QDMQoY/02e46KWhJ3qod7ryYaCz6sFewMEz
huxW93t7oet4cz1kkqHHXGNdP4Gk5SbDnFSGHKpospTqowagg9dNX7ATIOVIAqSV
64GkxwFPbHpR+/ZrWATjXvGYzTMh7r3rE+lVqzDI/kxJegbrIokOpkYUZD0tooAQ
FuhsVs7UWQnSYXDZJnfHJ5KEIJStPpalp3SMV/XwLBIapggGRIb4ZnzqlqJci25N
ZRfYUy2DXqg3jK8ED6nm8E1waiHahledMVw6RwE7b1b8wc3s5mgyYhVpL0G9GORZ
jq+uXaMz87b7QenR0z8GDb4+BNxjoLLluP+KZv78jCvFkJEoP8CVCyUy95Ra9V0d
zIJOmS47Q+UvOIUvPTvfimQO8F1hvFPAv3Y1MFp5BpXtp4i34oM9uK5M5mwTgw9b
bKkXYmw/QLAmhktlKWuF4MkT0PefMcgAnLZVbAQM0gsL6GLoAxXJy8nYwkLDxm6F
P+ogE9cFKujyFUmnU11VNcKGHCC+zdV+AX7x6pRxFavKZ+DYL3QRrDk/HWIxozJ9
eXE++9T1Rj+UHEEbfiAMU0raW2yBFGSGs4nkCboJhh0LXBVppavzl2u/Dla2oVMP
WAFF8mmeOGSvH+ryRsfu+nxeZ/nWV+wzhbPMUzqus5lASM3Qx78hynbEeSGjczRx
OB56p77V6HJN5QB/TTMrM6t6MMlbDOgesgrNW1lF05wQm4EoMsppEwWUJoSZ+L5B
nlaTR1VZvWFy4yYtT4OfSNoYfacJOU14wCdmhYsP3QWVdvVrIR8amXVhwmN8nTWh
esgHnTH5MOleBtLmgE+7tws90dcc88Vt9ZDOwjax+HEM2JXHyaO5Z0fm2WjQpqiv
kNSgwZVNNfeWW80r4sLoaVLh3pPf9uJOCYAVYIK9suHyoNs01shIMoh/9gzR9dSg
e8l7uDdAMOjcL+77o2uwd8MUVAqgoCne7xmm1Ls+X9MOaUIhB6XMvfLRzMmCWXCY
RUKHCNnNBAKChtYURZ9SDSOsmY8369edLSIH4Lz+AcX5nHZfLcM9B2SIxqIrFTlJ
Jk4Jwug7kvr5RwhI7Myt4gT1la9zbUhyyCQcnUBy4kcWz2oq5Q7D3rsKSVGK0lkX
9aCWcXHcM1vsepdE/JA92PHqWIEu4zz/zwIA3EJLZbHGwlpmD1Nh9rNPe8aED8v7
ZjJGJXkzOzg4hXpuZX3PR/BDiRxqVDZHeNQs6SjWHMT7ESe4Gk7W0nhqis339McQ
X9aNvGW96T/AKLwiWMUwdGHbr4W5DMwTuDA0FjZKthabTOR+v8Ue2clHg4bHxngv
TZYAVsgLqNubuRP/7bX89uTpQIvPoAM6H6ZNeM7o3O+uM7DoUIHuOBXQpQ3XlTiP
EAn5UApR8cusQT5axzfTxicEFITWdkYkb8wSaBn9DNuzQwlEB5ROLW7SL206dkvO
N31TkQpluVIOlhB1WIHLijaFtLcExjpNVHUl8JSkAXJGZy+pXH6IG8lC/MwoXtXn
l57KpvztJ0KHKaRb2Y/2Hw/XtHsRzW5vdXBHLZ4M3fqxV5s0hzdEhn5+qxhxqVaE
pNzU1/Jimz+YpeKAodNfGqOst/uiwsfZaajlSyj7Inf5neQER3A63G2XN7anyVTv
wR9crrnOek5k5RGLsyK6nZ8XjNJIPSGxCkw2F+AR8GtCKN2MTtg+D9M7hWA01Hx4
yONqSen8YQ6lkL5sW8ZTdKwbXyoMHrZUeNGOV5O0C4eZLcitv435e04Hl07yJoDL
juweeRINsZaa1M6mSd69zB1i1+xM8iiNxHvkIqh1vhvNAcefn5XgQq5FWY5G7tMH
r4U176KT4gsH8qhwg2DIFRZcd98OK19VvWOqYXVLzOJfvB2JSNWcLPT7W8ykxfQi
8RnKQ1xQ/RHqzyznowhmEvVIb+276FBNyeD4IZbUDV+2/gaxDUHrq6KYY+66G8i2
aLXkLUWariAb1AdbJX1cnhTVIxuw6jfzFkmOIiTPjyGiFCT4HgKOP7iaztJgto29
3XLU3HIJVNx1L9gHXiPJex0dMMQLnGDPyFeUfOEpMfPYxferoxGpHqmCto60LfyR
RWYd+/adn77NIchzPxNsaEsclZJGApDNfjPxK1lCkg5ybYVPf3PWDNIc1zSjW5Sd
DAFtX8z7F8CyrdcJ8ZOU0ZYYkxx+iGffxCtiWQYeKQ1f0ptmaYv3iA3ik5/nNnk2
W5tWaRfPTOguEUpSmUe8YWJYzFGmofoy381fGEVwoSUs3HsmxoS9NhQA/krHzuBF
7lErFWCku8CcsgCwJgsimjxvlH+504MoyjjHBtkH7LmtCYr1T/lTpYxXaqYlN8Wf
jKndrX1ngYv5PbwR22lrNJqVf2xS3yySCEZCm+F+bsTi6LO/riVTVmYxjA7x1lU6
SRNAnjNqGLZuWu9iAjXLw8alPhxgSXt5wGR/pJyMZRTdRc4vSQYUtd75tB1qU3xq
PF8x78jff55M+Q7RbWN3LW33otb1A+fK/CN2UV3RINdWivtn1HlXz96KCcs/mnKo
RWKVAfo2AsCrAMbYexR2FnctKw/bKAdCGyZxOotHf4FPpk7GydEhVM02HQUy3p+E
DcxKzPl5VzQLyHgytZWYwtT7pe6wD2qvqv5AParGFt/gkSgZSMXmETtnHT+5QC0L
I4O4MjuubKH0Ty0dv1Q8Eyn+jJ1BCspxt3Ugm6OOEXW1N5Y4EzzvSO677p1C/D+2
qXR728WmoVihyv/mOGDx+1wlxmprpEwYBXn/2rzU2X71puQdwjqfVh2z14tcM/wl
MdyAkOGCgmvOC9qghcBJS05JI00EQB6k7iCLntes9Oc6taPVXeaeRnYeNILxek71
qlMUrGJsB1aoaIlrXzb5wYKEAi5/gkcOPgW32/gnBmbeFc0Az9KA46zOg4XcElcu
59UkVFSN0LuUFVSyjlz/AVTI4a0vxn50BNJ0zK9LOpUPqhhgvbBk5dOrh+xJxkDN
8aO6T3g2DZ+2HhW4NwyUhipVtE5DgdWk6AYbD5lnew/b4NE6+kcpHIMfthHO4RD9
nMrib/VxkTA/dBMCMxpFStyhbiHgxW5xU3Cpry7YKr8IEQgheoN1HerH+Hl4tisJ
z5qhU1/HC5jeWJpgk3etGIHG8kGvzuCguX1uo1Ziq/7UtGGtYvx4wOW7JZbh3BRd
jUvCYKlFtHHxp81rwKHjaQtcCgSmfxnOhqbf1WHNbfc61qiIyC+ROFn5hMh01Vsq
ZSzsCpPO3nwcBXcgTxUG9jpSM0y3DFltUDNlhDcnKUYgwTigXy8se2dQtBQtGpAn
c9HAolh5YC2+QxOK1jvwWUCHWZYSDFRfMa9gJuURZ6iXWUlLoJkt2IFdOmjptJIs
XDCHWSveh/ecy27Excy6raZK0AAmem2qu30QO+YDdtV4OlguyVnQtaAWQbdPlkJH
vh03D/Gvl06HnE66cqg+MHU0XU/vXwAXiDI0veI7xprBjRs6Y5UT4J+hanow8sLP
9/mmdhlENhJ3gp0FTD3vP6ecpj77wg82lia8JXgS/sq5LtHzTGfe9z8jXgV3RIZI
nL4TPZ6Yc4uwNLZYX0mW+KXM0rEAiu1wuyhx1fFchenpRc1zPSDbk89n+a4Miekf
l+L3/WgKWzyHCigDCq4D5qoxPT/lo0nPtd2k3P+r1jtu662DprqEwNvyB6Pf0IcC
Az1XtTUp+OoHw5LWh8hzKM4giKV4S6hgWPjDF862y8Z9ofVKerK1LexVmTov7b+J
8I7su943XIPcofxuG31Zsh2uN9LWobQ3BLN2OzHtVCo+/uNhyQp0BbsUDVUsk2zi
AEOneBJdORQ/2Dq0gv44xkXhwbSEFSCcxGxmwEzaqrWLbUlK2BTmrmgBZHQ0ToQq
L0BQHCUgpqDeKCq7W+MWi3ZMHPGCCPDlePelFBETFul5tTPMr9HHIS2NQdXT42W0
z0hI+lrfJHiRg70hZ/7awY1zaMqYdiMzw5fNPkQbgVJCl0oKb005OyBmpSj6xvmZ
nc0W4fkhn79A3RCdz6Qst3YuMf5qH94JJzApG2KzOeilBBlSUZgfWW0xwJ1Rni8P
4cDlAF3dkjcFYhdGmKE3oZRWFOmEDksT/pJ4Qb9kPWr6XwyR2uJiY/LZ0UptdtJs
NszxA3/DXvATktOMwkNHWZItVgU+9qH5KeBSEazNIigtgSP6wM+30LoCYFKiQMSS
u+Vl/vCxdUcFIQ9EnA8NA/VH3uQEOsYMN+0IHXPCn/5gZzcz5uHGlsOl3TFqQtAs
j8fFxiymRvQFCm1DtG/s8xCH6jWdIax2pfAP70u1XXtSzMJVcPSrKhdTwjxXu5BL
dGM7S3+IwVZQ49qDq/r7Honu+3c8hp3mZqwLtuQl7aDyOGompDSQ9yRwzihz5YGt
hDw0aY5IozTqUX8XaMxx/A6LA6nMqZx29/wXiW/fFXNxwaC60VAcpL9LmnHLLJfj
ZwOeUfhbCIdktvVfNdU19gUZoac9P2q+AhCY+1Q8SU/e5hbwUi23kPq2r4OIFRaH
hSAk1WASk6/GpbiQnJyBdkz2Xl7mdmqZrP9wghhRy+JjUuwO4jsFDcG3r0PdnSnY
EAxBUoor6imCV3SDBolTZ9jJQ62nDGogXhPuLDhYzyUagoLPqi9xiVDoQVhuxH78
BbCvG7rAEON9rZF+nM8I+4DIYZHWIzElkO4LnEdDLGHzUqGPOnlUSjs++LlF/NOK
KE7rqdVC4XW7lGNNm0MEVvrlnt3iPfJaCKi1L5xHB6esNcYgKGzN3f2YYWg2aBIF
JCS/V7v0oUJokXjKLBa3/sT4EjSKCpWKtjKKaFAAGcKFwN8R8E/HUU0VdMOSKZd/
NuFohVzRlGJ+tJKNIEg0cLAw8wC0H4rkEVAtzm5F8RdsaoDZUeATetLehqLD9xlS
gDebeoaaLq9CSPX6INFs3BuVMG5b2SGtDLbbrM3tLljTam6gFbsUPGMaS27B09Ab
NLzH4wlduBptkG+EzOK7TY/r+1f8tu16bOm+YpV+Mgv/cHC0+2gt5xnW/c3PGq9l
vTZplV8gpJsS9gHJeTjSbQMkUduA6ddeks+sn/i/opbO6Q8gWSU1JIFSs6lS4FaV
Ra7iBXkSdVOuPg/7vxdGTxvwU3ZlRN3JMrbjpBAdesNtQ++U4xlNhZIWOJM2blpN
mQAVJErwP5i0As0HHvwnyYtjDaESjv9L9W1qXW6xVJ995ti7TjWQ86h6Tr9ezzDm
vhr4K/Dok/9NZexf5xwQdbw6J4/bl41ycSctEmO3NHAt8Ol1yMEGZ1afS69t28fT
ElwN6MU+kX2M1suThATF6bwATVtv10qf52Ccnpo2oZpEyax/b4OkK+hwMOds/GqE
BZbBHjp3BVy7tnqcifekE1aUAK//SdfPlPeOlvnylRdLr+7UWHADRdq8gWtzCmGm
bctSZgiDbT6bOzrXOppPugYPQ4HT8IlIK7sT7f7ugt3BW+oz3Ye4AEI/nd5036Zl
rLfyR82zjNynyw7yioCr9WhDVPZRKvKAVcf0gce6yQ92qj5bWow0fJOo6euCqCYE
qiNAwarUphok/Qu37Z8NOjroC6tXVKEM8oos/80FbA+sim2s4NPhE4Z/1WLDx29e
2arE4PZ5TmNa/rg8OD1tBlNTs6wtjac8E9Xcwlj7wSAxYkdwxBeJDpfQEzyKkG1i
7NAilqkYpdydhX5QGVnCGhImjFya48x7ItMbVp0ERrlMtSQ7Tj8S79ffKhDxG5/S
LrTq2+F3Vf1xOkcZnAX3sSkJTbwqCfuNjMmKZ2bqE61gf23LQVntJvzRdC1Kj93x
qvl/g5unrkMlCmK7N2V2w6ZHYdX/zbjDJYV6v5oTKzzEFQLN0w15GjXwBJtZ39Uh
2JgMFGSvII1FO1Lkz3bGKgHTwInG1RO5BFmd3dJKWw/ZBv7pB+O+0HihM7P/VAkU
AUXwlILYH7kZnFxhl+6+/JtUvdRSX6N0b27L5gWideOWg1hj6UptZMxQR+3Xwsnj
bB+X0WXYYjJjwn5FdeoO9hSpHLMqrrBMbZfvRiS8aqVHvgHUtdWcbDROjaFjulkE
G6m0HoMGswoz6aJPkQK3XrtCAvtoSVlxqQPOwPT2ITS8FkCCBRL+ze8ZElQTrd9m
K0la5250JClKsaGWlkhPPePAkv7GIffi29hlOOE2sseleWNA1TOxhbEXSAJTcg0/
okHb4jUgFgmcwrYt35Uykf+DyAlwuCW0YICs0RHmPSECOzMZ5zhK+BiP+qKO6rhA
dHr5hL7bvgSzOaECovfU4tvR1cK6A9cYvuj00jm4GDO+fxXDx+Mhsi6CbrkcrPP/
LvTyddiFP/96tmFAmzPalW3i8yHiNTEI+kkZCq2HxG0v5Vk1duBo9Cp4SY/z3Bx4
K1HQj3n0ewMSZvDEsjzfxSFDYlLnKu/pa5ijMRMARGPBuLDs/yZ+uiwNJ1lS0+kZ
9yuIsKvDo3rTKp2ULnRRgI7pKfT7s5YHYE2o/euT+b6Ruez6XQdW9L9eSvaeEdVM
C9v88QORGs66wd7MG7eqOtg3xspwf8o53zb4IgEumfFaBGwfEbYXFK6zf9ZBxsZ0
2oj38lBw3wq1gc3whTQWQyAiIYKaekljwWpVX+1ulZzguOJWNB5hF4Gw/lg2SAhn
lZGNZbkdIFU7SsTZ7prmY4fOucLtGmKpMq7/+p8oBBk0b4DlxHXzU83Cx1G4ouvW
uSX4sM1uNaOQo+MqjtFbOBEODG9GP9r/aXb88cBcAlMcuer5Y5MBIQtriLCt5Xej
yNFvQ2QY274Q5jZIdA5Uj0a50JKofHIs39mOHYTd01VzV5uwIxvl71UDP7lRFIkr
Xl+VzAE8LRycQd+uVY/ur0XNFQYUgt/l6ZdlRWOgirA0cGmSX8PYfM7wOzstQSo9
W6iThvRgf1kaqwqrzZLF5Y2nxqK7MtDX1vket2nG/OkjhT3WlWXGSoBhLPswXmZH
E3xTM6HEUMm3TaRCcDZ+a4uvgHzIl4sdBIzB5ugXGZPOfAq42n1LuoMJ6xeI9X4C
PXUThXIgXEbKpj6LFBKWihDg6n7YeeEqaKe1qX0dEBf0mPX4nhvgUV19Rkv9ZWii
vi0I9ndAwuL0gqzvfHFNeDQhZfPkk7D63eU6tsc0K8tIVMKz35pRghuNH3xlWTVl
DR8kN0bCQW/glC7D3PFhRyWIZhyxOO5TtZS/J3THgNNk4/V8R/ZWVcOTwEzFri76
zPfzLxecIMDErYZFGSYoT3rcChyYgYp/wm4jlhka8u8C3MdtHPul8J/+tDYD2C1n
hAV/xNfogDGC2ui2tWX4VOufIR28pLKLEqrfNukelbgw6NB++KhgCGbpP7hSJX9k
wKsX6sN8icsBh6Pclv95Ia2kqOkwFDsvN8Gb6J2gwHc1XNdawgBrC66gKa2tvH/L
nQdNCJ0El+7YrzDmK6g1gdJpB7QbsOaqy7KAq5Nd0oXlnYrLqQ4LYdeOR/ng4quI
NQG5Bvs0DJmzp6vWH8LSfVYRTAH5EoHWPkUADtHjWdqs0sJGa2rwlJpkVIPLKqh8
Sv0iptoIUUoc41PD92uM9pKLdb9qIGwRlxLI1qsoM4AcjX4B1B1kmK/4Wb4257jL
iQlhz+1yLzJNfPaKZa8TAVWQ7rVDJ/dp2Q1xPhpUWSSSmfKiXdUstjO7HmFVb8DV
voJz75o+/KSSGjy5zUfLK1WRgKbD1Et1of/8x67MJDYmUM9/E3BTh40SObfc7ohW
k8DHwk8GwJR2/wkXiqqopdLTDOzi3HlGhkdqKD8YoC94L6HEppVU2YWRImhCh3FQ
jvZqCywqK1v3hQUma9XaoYtq0ip6AZJ5xPH67mE9HotHKX0Ebznm8bfYrnmUe16S
hi8YqUVnR39N5MsWn7reVA9/hQCWG4TsCf09gDv5kvsYugQHOB27jKqJxYQ1x/ll
97fBZnJDAfx4r9nX9euM6QE5WDOf51G71HfAqSJySoMqAe5P4Ff6TQAB/qXjq8j0
SXxdkDI4uwDL9vr77V3AMNsstIHBRTt9QriPZmfSj28N96kW8Moi5DB5hS+I0X5d
9Kv29LUFzb1oPN8TLdPliZuYueaJ5YQuYmnBXbHZ/hx1vbXy3lqRVrjT7mNtAMae
papp+hTd2+/kx5bQ4NodXJBHZZLhdxy8g4ROM0xWUJfiQjZ4TI0LKJmzZ2N3ahic
NyfNnBdplD2F/MqiRwH+bY1dN7IfmieQYLydtt/+BLGfO2xk3vVUWVYyoafDXpp1
+z1CBqo71Zq3BJnWAYIPQ3Q3l1xR61mIwlTyF+ISnCAmdf7A1eWT8FJMKa9yQgr5
usHXPqMVwCawj+xRJZlQPxJf6jsnfJTy5cDvsJ/r3nn4PxnyWsgbSglqqyAAXqtM
7ydxdXT0TlLUjS8cemVqfucin9F7kOPourMdNrxS3Z1AL+t3xjm76yYNK+XdInDD
ynau7B2GvpQnWSc9SCjA53gMJMGwaXxCufraVwD/+J/X6nqWy5bSwaEFYIbv6l0Z
LqyTBHhoP2yObnR2kh3OaZMM8kYZuUSd6V9AYXIGI7dCL0Ko/U45S6cqkR2CdQon
yA9i+xDniupjeXguxIgPWn3KgFw5i2qG4ol2cmi+ZRHH4CZpLI12qy9xrphBZ1lr
3N6iubxAvK4zlQam0QN2GhYcyTQmakGf077OjDhvXG+YHoLqU0NOnCgfPmHL8QGu
fwuTefyK4Tg3dHFIzmSqsWZVvIl11TQXeGKCi3P01/IHdQOzSu4ZsrZ5C+2413cG
5FdbdxBXXTDKYoTif82MJME5wcS7DXFGMZmfcFddoPUrvj5WKnB1M0gG1WBkz8SB
0locKPDjNcJgSwILVb1mpHK9qkIV83yVcPW/e+y1J/yviCDE708F7wCGelEO/8iv
wA4itHgjWoGck950vW2sE9CPT2M0Nqdj5DEQz64/txVU3iErgR1ZeR3FYPjD4Mdz
n2BhiOuV7TwRv2OM8Uah1rcjTeCZCjeZlq90PKRbg6VKlNc+p+MIEsRk1Aalyktk
/9u+NHSn6Jxm8zqOu+YiuSxKkT7SyxzWfgaDE2NwFUyzJFlgocZwpwdidUDpvIQV
EFB0qIhSDIpzNwZ0AR7uECn1/aS8cmN8kvuE+Dee5iwO59wmpx0vF/q5bdAAy/RN
NDk69p+Za7tO87g6OIBWtVIFnyVGmdCT9PFXw0VoCDuB0W/d5Z8aJ6QZCVQEz8Ra
XsDYrSuIRtnbPAzfFIwcEKXlKfgcPXIRkGLSul7TwY8Up4LuUbxJhcROQTcfbgNE
cgVibNNjMy4cbH3jafoyXx4VDjTFh8A577c0eQi0evkiIP3mq4MyvgcXC3xqNR/7
hwcl646WsTUzRThqdkSpI9vvKLMSA2aQhlezGCpIWt0WaYz/ZBY9zqgpbriAk3tg
GnLF+1JjZBLoMoHjS0HweYPzKi6SqirL/6SjsdpHcsr5YCGZVXSzpo1rrwISV9HC
JiiwAT6RSxcnqYjFieHrbpB/v1dUGooAbK+GmiL3tKvkOBQLTpsfg1o5BpUn1RXq
IO/wih4mpxPxLD/9QptAYnOJMGREjrMFZl7wmLxm3N6bYqpUAolbN7AEWdNb22X8
mjWdRubNRtdDpeA3ydrdbad7fGT1/+SJQfKiEYR6DQKNbe+N+xZ6R80sbpUBKx3S
h7twacwflsa4DfZaRPonBQqiKgJB6WOuHlfbMksrVSA4QLhk2bk5h3H0GcxKBPIa
TGhBTXPlKrDvAjAUB8sdkrd1rl8czlT0aDk+2M5KbHoCVreYongyQMAQKLfWJXYO
sWY+Q3ajK7sSTZp1S/wrFfOR1GrWVRvGQSrYhSlqr8YtSiayga2S9uWSEzBnVsnL
p4+NOdVEa6mkyEeNJQPIkVO9aCDEhF5klKHiDWLGMVJb9Q6Wpo9NLsspZewMuIP2
aNDfSsX3QIv2K8ji7VQwgSvfuJdpry9zbDA7ie0Z5AizhKKzj0Gb/U5jRlSU5VfJ
C2CexLpm0mpRhkPOdHl+Pnd4cA1Umo9Oqhn6bm2stq0fVd+fanj7JA1sk5ZLHJxt
kyKgdZDysGHdhNGuVvdu7TahMe3I/nC2VYrFw5rA2xfaLWxq1+uarXDYQWR/hDdq
VTzkipeF+9lISsTw2pVnFK7qB0iz3U3GRcC6eNb5P1oWlN9wqAKFZgcUadp3BE9g
HRyso9u1hSiJtXNYikC/osQFY+1SOua+N02Gehchqyv4JjPPvAjX8MduWvY6VcSj
9xQkgJQvGOJwzJMmbEbRMHhymOZW0fiOul31xv36q9OmyL2kLMWIyWAELgrsNDfa
oZmvc6nvl6V4wZgq1tkhkzKJIC+fZUa7DS0LsiyfiMeuBgVl1myBLGs7+Dbyktb1
p/abvNvSu5XygxGhnEPhfhZOVMOp/LAaSDTKr1XD5qz+m5yqN3hWxJ1y8qGzlsGF
ZAFPxy4NIC+FiQicCbonjQkSPWeP8yKy/CPHGQ5v48dRCIfIjOEfkEQcbzoHxMPH
ZwcM5jHOguuzWZWLHUrVHAwVOc1MJxVw/llj1GcJLXlHUYKFubEMvcf26ZZj/AaC
rfCXiO8dK9gBQzN3SLeCgpaB7gUCvtJNo0yQ25kjdjYFafb0E199K9OpunFA2nMz
3rKE6+KcGLEL4famr6W/5C5qslPYf8uDOSpNibvE7fBHupysW8sjKlOhg8FV803L
U55YMbtFj24Yl1SIgTAdlyoYtUVSEuzc6PlYSqrFbipehEtMcPNCwee2XgrG6qOC
zYESZvVSqwJO5kF0iXjPGooKqQe8NVNNbAkqKSrTeTv1uMAEE/JiTO4tq2gXNucM
U98vMn2Fn7I8vO5b/nQNDgUt6ObtQAK8hfj10kdJAOTwbo51K5u3fSGu6cwYxD4c
Jkg7JpErf6+3XWjImOSLohJyxwLounDeeWT0rTkkRSVYbep5PrfRQvSTJalRzkcY
Dg2q9vZw4XVAL7+xBM3eIV9kj6EImvnlMiolGfKbaYMEQf0Zw4BCvh0Z/PCuuNpY
6A2cHdGQQrKRlN0UJQPR6bk73MZCu8qbZLU8XUFE6YKdkc0osRg2Pb4qoRJr/4Ka
/E/E7tNS8pxzp1okZUw4p0p1l1X3U3bHcAdOAERGPq8AFZu8ehhSUNIxpos5O/qu
1zR29n+DkGeXPYanzPX+3kwaprJEgzdXLfY171Az4tw8e95NQnHiuISLfgEfOYqd
ILjLFYkLZny+7UxJCL5nfaoQKTQpOy+Psa9aHx2a92HQCFgSEHHOeTdPLnlWG+Qo
Ag9gDdXDZ02H43GuM9drDvY6Yy59zpXhbT6ehF942ZS7tjXmnYa+kv+Ptojsu5N9
8fiBSHV2rkErDyudgQYVhAkn6N78biIc0aON1f3fSUk4leq14MsiwnK/tRdnc0cC
ektAqANkJJZwY3LZqIobT7R6I/3xLDPvUQovwVRIYH1SeUY8UgFwWmJIe5/8taMG
PB33JVIutZ7xdwbJ7NaFRume4PpiiGfcrFRTdFsfRn3843EAI/wAYmecEfV5ojUd
ollXmQ6l+SD+JZBJFvX1swVDkYGE1fa69G0nCNQv3oFlB60A4kJ5rP5dMl0myLx2
Fqc2r+SLLB8XUrO0FR1FnEGEDTrwb4RGE0YcZfKeVjCV3CL1ZguDyCeozL6r29ee
BoKdF+t4tZnrNpuVAiyNPSbdUxcWSkiyT4KRsTSvkwftcJYzpDPLcmx5nbClTXFq
SviHRUqWV3Ydn0NSC8Yof7hzAMopmYqKC90tkUVOErq9nauPSEb/AFot9dJfPsFS
/RgflAff/Pv7Rl4DVFSEp0WqeNlPZyGEbZgzk/qyfOS2W1f1vigzZhyojRvCJliV
zPBN7KF+sucAGZ5lUcF4EIf1iKcvQoc0kTyottJjTZ7dBNE8rSi4Y0o54H88wv0N
zaY27FaMWfExLGMO/YH5aV6wvLtYGdcZiUtwmwS456Z7BKQAYtvW80/De2wA6goT
IzP/ztfPeB56vyW73v+HH9ahASuIzpovraytUCW8qs6+TQvYZs9fdWs6dPw11vT0
d1UJen1IdME2ECbYBYbu51HzgXs1s8Jd0xvgKxXiiRf23iYqs526Ul+gFN/xgkuD
I15wHDjW/H6l6Dro4QU2tXzn7CKjNBZ0kTBimbtZSwqpX6ZWmq45gGc7lkmjj9sz
2nADxFC2D547sO9Zbk9SaK+mx6OXT3unWyDRYxpFR2G1zWWyxC973M8jrHiJZlNW
O2L7BY1vasibhUHmQzmoJMFHKFHQwsuCORI136zwFkpirvbsctosWHeinsHUjQ6W
6zqG5wxFdxrHvRmI6quWx9D/mUlpAVfF/wRS+QI9tIfB5veLK0T02zEX8K7sZ+Vo
KwqOUZK+ZlfbyYJc3Fv8QtfJleLTrj4m7BjvR1lZjDl/aOAWPLnTr5fU9W6nM0G9
VVU2qz8ljNwiB/J7paspDq1IRPgzt0t43rRtLKvnkMs76lu6+DGdlIQToBQ8Yk25
73F4iCgD9MhlK66pQt8svhQ7BD4N9vkCyN6ew3zn8+vHjcTaEU26SknOdAR17S3O
hw5VRhB106ExqtenYHSm6xoD+jWuPqPzHfUNxgLNPQEKq/dstRMvFhdtWGvLb9CZ
Ybx4qSM2TpNjpjZZCOcTCtrDKg7ewoV55WvYPWB6AgxQJh7WB9E3vLZ9Mv/3M6b8
+tuHflpTyWuVEbSNKuU33fjAQJJitqu0soesPfS8iPFPeMTZq7OxKUzikmFRNulX
iSUYqTcbp7E0+xwGMLHwrsJuqUUG+4PCpo+l9Yqkd4K095x+SzELiR/S4kIEUzwt
4oDSnDpG47avvLCpuopisEvcjaWupezvaJFo2R4vfuLhcKow0MAVsMz9K843QM9d
Xny9SDTBufsz7hWrqBGOgzZ0qplSytwf03kAYQsqCacF2hZGYe+gedNHn4zaNW8A
KbCqMgCffg2zeeetjRyht8L5jcI8cbwB/FQ2DpYeRGNizE0Iwso07MYuhorqI/nW
F0SgZAlS//k/DCy0gzliGO0N5wNFUzLBFHeRANW+utETyDEJXGLwrCiNH+BJXvac
A9GBxd9KFVH6Jz165lClKWn2NQGlPfwXnDCINcXaGJy4wTI1UpRpZAr9LvneJdsD
eLhskUWjFU/8VlsjNPCoyjL/yAdNqoN9JVasA8/BtHSCGGnf0ZxuD1jWNEM8f2b4
jmxaNenfHG2mafTAcPW8rMBG86kD3Yb9uU2xzhPs7dYobq4KHSQcctjR7CmnRL7I
6ZCLDHrmTS6i0OWklRaXLduZi7du94es/wvXn+8Qn2uqWWKAqX+p8mm6sTMKT98y
fRK7zl7AgI2SMg62++Cej+EYhLw8jdFPDpuJ3wsLn9Jh3MXa26/yOG6C9RqQE0ez
1Jo2C7v0DAG+A8OfhPqND+BOcyXmBN3sKG2W50jCBM6PIwrGP/2IFFRQF7ht4YiE
H7b1rrrWPpc9woeq1ojA3gX1jktgVCZvxWFd4vVObFCgDEX3kJnSys0Robki9va7
kpJlFQoQTo0GHqFMcWaPy3mdNXi6gELuGSnEjHrBxAnLwgXTFBY6oWE0ryMSjswZ
KvskTjainpr2IuzLwJ2LLYSKvFUs+6RIiaGOLVQICQfg4aNiDi+5KwicMmM6ud2r
VRYGf2mNv/Y503OnfU1iJp1EgK0fjh0cCMhIa9g5Aqv5dn9MA3Ayyb3p62JcKMSE
8asXo7iCqZOJgcDh3tn3VJEyorToq4D9MrOMaFFaOhy9BJMXfpTJ2XiXEFIQCx7u
LS4KrAoR8OMYHZPjr+MJHp0ve6qKE09D+wpip4DC3wqJ8X9oPseNefcg8knchC6z
aOYsKd/JBGFFfX9Jd2hQu1sw43DPdllSxU6izTiogsrJD0tEy5kT2dQJTuA+ErQQ
jxCMVKRfoHInw3iICtM6XCId+wJsXWnRh6wWsCbwGFCKJ6XiB869JuBNOwA2qaQa
YCT+Zxb1HEEA6Th7GJ7yE9ixbrVwlgdkDCooVmsjPEhiOaLglA8zSgh+923VlPg+
wcqmXmKCMB75ueTJPG5jvvdnQr53O8HC7OaQf96Dty2XcPkrlghCRZ6GgC3U5Rpe
VsqvBuI2e+z0jZThwAFsom9CN9VrmXODcwRVx2y0MQjUhEwlfx7nCETwdBb9qs5w
nYTeQDtLAVVlXlb+AgGHgQPSu9jUZ4c5SEeq4BL6xO/kr9eYxGF502HkmM4hY3lD
CA5sUM3FiIFPUCXwnLZk3zDqik1xOgWnCBy2fuAVTs0XFXSWg/k0Q5Nl63LrXSRF
2BCcxZIQy462HtYHgdxdTDLrNKSiNZb1DCRYY9NaR2I8U8T8iE+Il0QDvD86Sb5X
HCNG1OLiKeMV8XNRO6Ibskxgz1SGnmlQhV+PlLmRJVBYw7e3Rn0zM86OPPKgy5ep
n+vL7ZzwiqOnWG0cpsi6S9wF6QWzuH/wf1WFd8DczTsLKw28H3aHHSMYcp4fYhWh
NkJXMLkEPM5fA3MDX+JpuLjkN5TBUPC7D3KUATjHvfYoUjW1A7XPIzvDvo11dtrS
hP4pnQftU+eWdtqrfy5q0kInKXK5t+D1RyEmtQVLgw1H7uYU580cIwUucrl4jO6v
unyuGryOhPNsppmnDaKtQg0o8GY4iF+GOV7kAeA6wVYLDws5x8EJzaOWDIz7P5RW
IGe3myTF2YiAmgJw9ilO2Pg5fzvwGdsn6WQ2D4ljm8qoxHyQgf99Cf3viXFg5nqS
0sS36fnNcyYnrS9GDA3mPt90fTF4eWRvd6wh0Yq+zqLXki5ESmqM3D/Iwcitc8Og
j6av47bj+ZnZc3W44be88cJ7aaDgVXzDLqILJztyxNEAqPwcCPrsAWkpEBpGdY44
6C6DUyOeksK8pVOs7OD/MyZEifglklIX5T4xZdrm0dM3HMvKLy25FT6LR9/CAS9N
pcOuOu3SFTudhjXrA5IzMmeDVPKkIEJntqC1eVpKguR4WVj+cKWHQkLQROJnnGmP
0W7mDg2ZvP7d2vGe+hiltH/z/KudzGSyjOdOb2WACEFQjn4wkUpU4cUxG17EFGWC
FvSbNOa3Tj7zW2uNjZGwPXOulJOfBzzSbXOnbqqZea5D2eHjPOKz3lQZs3Vd6W9z
RoKJ6DNCVGVjAKaWD0PUE+0X0GBNcwuJ9OIKw1Rl3UX2riHIljRyYflsEcQiS96j
l78qcEZdWikMLAiofqK1bfuGiJ+dIBBTLY4CvAwuyyC955LHkOpcIXXiGE6qrXSm
B2V0xKxVUh9sxsU2d+6BAXLcK2kgp2jdf67U2GIQgJr7XKodxGoDmloKI9TB4G7M
2BE1192spYbVuzKQptgnmWgh9hpWud4dJdLbdr4rL25rpZB0G53J0HUqG8FsxTCr
/1gzIvXRPNDGqXu6neqRBVd0HI6cBgx92b8FZrfDM/q09LuCiC5dbPEs/0uKVrfk
mWkkA8dr8IDqYShNxIF5P49GeImwTA6lwLmWF09eT66P2KUJNG7QLk5NYZOBccrt
TxBTmrbHVwvx9Ka5ubRIBkxRgeaLFnffg83DpMEID9wA5xR9z2hfwWRrWac6auBe
WikK1chHOxyjRp9kUn6WoRVS/nqNtrAItsyWkG9Izin2T83Rt3ySoyFePNI7oPbf
C1YDFZvLIqWAZXuMiM3Tw2LzAWrif5+hmyYlruLiyP6I5YSU+8p+HDZY6kJtN79w
ZJQdGUa2htR5jjdtGVbadHjyyvokyIRPlW15czDZGE+uvUQljKE5cdQyFYcQxT6J
6LW9YiUuYSZcDUnA4b4XsgbTYZazpd20aCP9UVzRVw71Ook2bbQTJgc4uDa32oDc
AY0eA/3swb1B3IKuknDBj0v2PyCApLfFSDFNADZUcRFFyb2smZiBwpgP6PyZGgXV
fmTGKmDSEh5z7iBdNppv2xkUFQTEDUp58KzfeJWbN86VX1w11rh4zPV6iVNA2H9F
ssB2uIAiUmGwvYW2vqX0MrlReVP1VSeE3MI1Qu5BHpva00R801bzduUnH5D8T2SL
mD/o9w0Gbxa9zitRG0kRAuDWdVq/BjHtdrwa7XR6sTvb8K49g9Bduv2WihuBnk4v
XLcVxkEJ4xbF5FIov1N946WxEYXyIKYoRiCVqebEAhCNR5f7YCc9P4JCrRWyqeIm
hJ1ShhRITdTFsENwUtiF2MgRJTpz/hnjlTLLxH6nZ2TUSjpEcQyedH711ZePVRvK
NxfwoHcBubsy0QWJvfhwZhNA1nZUuxWEB8dDKCaQK1J+pI+rJVnjAmGxedt3zm5Y
+NhlOYVThGPhVeN8URqH/Fpg8mcnW0NoqAorfa2nZqOwH9tSRquV/nZ3S4+NOV/5
Ldccr23wO15a1UUvAxz3ugdHAeSfILHALggOZn1ZmN5drYrEaFX8IkMwGpaRXS67
AEIZWXp1MtjYcbdixJnuHCyC3GGFA1OiRE0gSaaowc72df+8uKm1Lg8MFx67AYBL
wNKs4pa/piK07bxwgaQGEwBAqfaxJOWCOni7BNrIZWs7VMVQGDWg0Bzgzg2/NQJN
KtlCPzgjZsFrfRihNCT9Bsdv+fVav2j6P1nFey1tg8ueCUlGuyhGp6jktLJsDDjp
onsk4ltGcjJCLxN9tUJNOzGgsV4NMPyQx/yhc8N7oxJg8PJJbLq3oHxf5F64NB5L
neeKQTANUVreb/CQcRJnYCPsel22Tbg7ZQIPAXRqkMS8K6kVPbXN3s+Hk0TpT4p/
C67Er8NFx8xh4ltpdt4/AynzHwft0fjV4FnFPSuDf7uRbIAeMjDQiIguw1b4ACYr
UEg4/G9uhoj4TWw/dLbohBKj+GJOveZajBx5EWxUNwN01jxLgABBrIEeFyo2PTRW
s6jL6V85hureNvmo2vh9T9YeHJVVAVgAMAZBxoDTtRM+e6LZrDxg+20nR9pXtnhN
j3IpEsJ2oQNcJy77E78NXaUHo/pzInEZznEJFUOPylWdChcZT6DC4N0fRYL9+RnU
W68ATG7hMvFrbI1wjWi4PqFEcC3gw9UKrHsY7xwKcSgkrVcWGI+tX8uTR3eDUbKj
3hoRrgyL3cjjGX8w+y/rHHzVu0460XmzaspWLP0tQb8IlXtsPDhk8HX3yNkfQ65z
a6S3t+zVNUnK2YDF6W0CEHCRmXogILn1Mpfq0w3bLeJhMOAcKO6kZHl68VCTaiee
dLC5D1KzuHOUa0LlHc9PW/s6MWQhD7aXw5/T2ZvXnE3mLv0gm3bVl6L9PyF11kLm
mCOnA7ZkqpaRd9KNsgz1yOEOjqZHJebkqHV1U/90T+4M/TxzJX4uzhISxrt31bih
Mqpxh3O6slvKCtOKU/FvpiZ6oxMMN4aG1y/rXuFtVwJeez4aNma6dOQEFMU1/kkk
fipValA6Y6LMxTwbQLDaxytHbY4wcwRQ6kLc3Kj/0aZkYH0lgxHUThn3c+U+irLQ
3hp5C1b068HTwUu0tyGCF4nETIQS+NvpTfjmLH5GFsXLdreI19mtfuSHmQEAxjuI
tlNB5KTdF1cecnRnhx9Rfn9IG4X57WHByWBjODkaYJ/rMC4PrCJX6GVKFZEG8A12
pGnEPTAOl9ML6o/bG6ffJeTv1KPCxXkKEc5DCAg+a9Thm+Seuj8XpyY0RcjM6G+K
2PL+ajr5G8SPMwEXJS9Am0J8LaeGbo0fxWlKPB6CXtpzSrdslEQiF5PLBe+r7vYb
MxlGZ9BpwroYvQXvI3F+CoJ4hKVxAvqj2aqtTUb9BQtS4bdRF4ncqdDLYVTzctxc
kZw8EzcCBOsjGcMRmoIlnae1Rh0i+By8BWkEvZExfuDvfMHYHjQOCdbiM8dZczck
sZ747smC8FJ3Ef8Lfb8KLY7WoTl/DfxfNXlHeRgQr1A+IeWggpX1ozMfSyYZcOvi
xANeI+GPfD/zAi9+1VV+V6Qrt4cCqZQiU6Ji47OevFTc09jAmAMTRdzPX+CcmjYR
6w1CgQsUh/0RtNP7kRcZ2bQhGw9fKXb2hL9lB2BNtLvuoCAIyteG78U+kc23Ynzl
cNjyn/49XTwL4ruB6Upi3CZMnMtMt0u1eUb9nlhVR6KTdWNAzK5aPXJr7aDFaIq1
bDCRYrsM1SR52gwisJa1hIMEZbDZjlWz3taHIP9TRMbg3KRquOkelCbOS4OZl59z
yhaF3g/F/JhGYlpwC3h77bSi97VnJzQYBpFzDtS0+O4t6UmY2XAzj8POW4lkU7Ap
YTrejcE6SDjtOEoUXYPmBAAN9bjTU+HDc+WCZKIZ+dEO7/ibSc/Ca1EyhrGATKI9
mNzTPaQ9V8Ly+U3RqZs4eB98k8msHPiJgDK5a6engmnkIGw6sGnVkro+V1dos5m7
ye889s1xvv0MgISnwFk4b13669AJohep3W3kkcuKuYMdGESFbVDQ1V0LMlsoHd2E
yJyUbQVt/li8FSWBcvsnu4By+mc1oqXed2lgv9SV+PtWZwQKdKNxKZI0q2IPbefE
7e4mxhMFlsqDDPKsW6yku/c89kk947NL0viKj/IWF9EFIirJdr4+FBdoe6ePLa6s
5qR7KdMoiVPAX7Rs9S667VEnVC8GRUH+zn7gHY1HAeKWxzHBsLbgzpP2Igxnz/mD
JBstGGzXgNi0Eu5kS2qZauOSoIZnMv5iYaRzWx4nIlw4N4DRAJym9yPhyh10gEsx
nfh47jauixpQrhE02E9zvbsMQOEGpmdYYuywfgRuXIQODgap2WJDVADWOt+BcsPF
8yZ0twuFkTqx89CejHOX0KR8gkAE0tJIerqHtK9f6BIfALSF3XyWs5CjXORydiUl
5p92IUfqYjfakcU7uITAifhNFLHxz1rsPhXswi89C8KSRtNgNHpk0aeP8zNG/u3T
7eX/OGWJHynCp+zCP+rr+EtuOgU8TwL0l7ml1P3jFko5AxCOL5N82sCLs3K/OeLz
hBPWeMz8v+CztiIK3lGeQYl1GQEYp5zaz9b8jjvkjmeEHe4vUwhaV8u7yBMwSMGr
st83ynWLv0YWi984FRAGaFT3EEXiHrP3D/AtiwSfiv7idvSIuO+0HZRiBH71UlEQ
6CaF+5XzbY5K+YqB//OWIq9e9v+H10NIMskY/iVSYQsuv+7MXIhRwjcMyY5x5i1e
ssh5g/hsSYFfobUVDFJdwPOm7uTJ4GSc90pt7Jz8Jkk4n569Hf6+Md+mnDXFUm7Q
KlansnDE/8sAjjMTU2c7+X4qp2+n1oFdDFH68bhzEXaN7ijeB1CsYJ8qOyd7HftR
vt9g0jKBmW5C+mv3ku5bzKbP5TEl/hqxfA3GgxmClvC7DEkL7Hd7BAwVepHAb5f9
jpAQR7juxUTCMD4FpZyes6pDiD8+8sws/4d1UFyLaUym/U64mlH3qlXtwniqmDpw
E4CiSsHYA5HqVgtJiN3GQHARa0nPiT5nKIcZFg39Vmgs7kyucpryT8hhCekg/Z39
QBlGZ+0SE1Lus/XK4/X/V2IwC/rmgWsteii3JUHEzjzKWdudyYVWfIQ8MZjazOQ+
2YZm2wHOnl+TKeuUAieNnrBP1BhdxiL+izWzR7wyi2Jo2tX7sLLs2nDxgGW20v2r
xUdXwpWWVKaWqADVsQLB8y28Ln7PMNznVuWE5LELzJjFuzyjbRbGpW4FBBD6LKoS
4rziLQyMncjzOdpTKUXJOCVKU0PHUJOAkCpByBSI/u7E26BuCRFF6DPzK6y8PHig
+PfLjZHFjxNJEHRn/FCibO45jojwtAqXE1Nu6VBIxtjG5iiu8Kso25sa7T3iZBTC
JkXLsC1Mkj4vipyqr9j6RfmafsHT1JCqAvvimPRfzXJE3exw1BmjjLt9Vf+7AWqL
vshvJ00vAZs1cSWa53yprNGM8JrRgT6emgxCUX43Sd34Wl31Zu2IzR2y/xhQryyo
NJKLI4J4fGEu+U64lf75pxmNXalz0kaDhlrii7guzqjXHxNP8UKycWon2VN8AYfG
ozPmzZGN5uqjWmsmwavVlUEZth4gcpRMv52keG1TY+dMkIPlBmJtISBQb5Tok3PQ
iURC3TQdrS5vMtjwKKlJGP4/f+Ty9TbfTSq1u+kEn3ZSjVyfqy3eaOqiMnOpQ/LS
0FBA+fPM9PCTcVThVryLGAt02sJb8+tWHx+1BC1Tvqf40MGw8419JPaqC9deyr21
cbpiG4d/Qxq9LcgG7sTxQjnX6eg275S2RtTCDS2iz29NSTNSiCB6fS2t5kRNhv3F
8Q0mpAQuZ2+6DnW2iecet7H0z+G9X4cJi5n2xTC3Txudnag7G1/a0dzQhkkqTk9m
9J9QiW7/21SdS9PrXYCrnqfiF1MXnUcitgBT9FOwrgAh+pyKTt8vYPGIV71b/d34
Mb+XRDU9c56AmiuakS4HtFCI20SRZ/wsh3mTbJUqTRjTAaG8qDbR7DRGSexyd70D
MbCF6XZu94MoS8jWhkIV2YtS9nahtioA/J2YmkpIDT3AATHICt3G/mdUsfPC17AP
qxSokQ4TIQtFslL5SrbmaD8D8BNTLX5D7cihO2tlMi0lfZo49soafc8BOZi9TzyQ
kevCuWZParp5esu/8QBKpB06rsFZ5CLWFx4zpqTBH7MsczHiCldkPM140CLlp0Bn
UTUDm5FsJvapvLI786Omd2dj570QeiHKWEKv2zYh/VK6K3dQs81qoWCGQHDUTYDD
GdredOatvzDFrwZAUvAUcLN5lQVx3fsIREgg8hMnH0U/lzf2bFVUfAzIkaIiej49
koF/N5jZJxRWcSH8i9XZ7I8YsC54FeOHoC6lKNpEUmM/aaApGiMtpi2rxRAERZ6X
nSbT92Rb34xOC76VH2X6pp78woSrYQpoQpt2yojlAxLmsGvtFWppYV2N8SGwIye+
yqjV/UxV3sXK/0FvVRk6TG08zbNeE7wn71I5QNiXogBaXUp5EjajhyBNqNoKeprq
0Y4p4K5voEPLsHd42QRcYzd8iOrIjGq8ElHLEUu7a8hTo5d1+V8d1bhp7JXBDDwV
zTl7kO6GS55lwOiaI9XE3wJwRcUVe+jhCXn+F164TlxIrbzmAGMERc9HH0IHhKYc
d5xAaRTR8UtA/Rux78GOhLdjC53mUPWMaP14E4JlBRJwR/VB7WrNSMwdE9M5wk1g
fg3dPi7Uj52tDLZa6/VNLVZIWwwTBKA8BQLamJr0tlGGo/mzuAmZ+1fh09e/JEa3
NfQK/GhX036/Ak1BAsGVHPpxtXNuEViFWFUL4k76GgZ1IzzvZnvyNjZzB+L9d4lF
ayvuQmcSb8dQs7/21bBLux1oPStIS1430nnujWtSu1aiQ0t3sCdKivZdndMCsPxs
M8HL1Zws0AReYXvkSY9uKFLVkR41xc4GqA1Q5csyim4HXvarLYeHYQLuyNx9taP1
yxMj+d3CdhowkLyoaZlMHvH74K7YpZxyauUadINiHb98bymGiqPoO5kfjRsZazEA
9ZjzOabofjfphJT0b1VDTKc6iUZm7Reo6y717OBITxW9VeyvWgc7TApD0hzf//r4
2awpEfiYM5Z+WZzn6QkSzzPVw1rmwNlZX/5RAHUrjP3pzUVMe5zFnMaVWQ8IJyXS
OH0sG2Du03uMNyPkFPmZi63HCNwVpiZOfZlsrRIQJuwkl7/MIN2OoLAXcdp0yxT6
84l9NyFwyceEl46KyXHN5g8h+SM1lPbQ1nNWWsMIcA7gRIyUhHPFT2Uqkt0JJ+vP
P9r32B82HjdrE3BneQlPPvGwPjyhQ95kB2pPmXU06Vt7MizjUvST8AEV3cuybeoE
XX8dZQuD3NEXtxxXptDlD+m1b6LBcN8dn8FIf3i85kkmlMpdCsHQ1eLP7vkCS71B
Vgtf081/9IhygqRQLKB9zU8ZSqlvIGYFWVUggC6Bt3zn3ruDFtcOGaBTH5FVvjp2
RQqFbTJR3/kSr0sdBdeauW/GJARMFR1fgX7etB4OFhk9nW7ofGSVqca/O4t0cKz+
4pTWJCvNa2EmkG345mA4JR5gJ9TWRHVBoe4nUBea/U/1k7BLLiuVFIXS2mcfCNiX
FFVImcwO5KE8hj0PFUYeQODl1gkDI+hkz2dHarvOxx7KbVJMALq8x3W9WW5iJ8Fc
QRnJ81z3iQ2e7x7vYq9N7S+g2y3G2RU4a05PhNX7AvmUAWt0QAq+oxeyL2RyL1S4
FbCVaEIVOSffqiFjMIo60eKbtrg5tNc2vr6VhAmXSoZgaVue9jk+TTLEr2bDaos8
FQ0cl5icMMDjQiGpshBlxCMC0G1nrHg6p6xO+ArgKaIaedwNlSBtaJBRiLCJ4KVG
Imi9+MciNQASt6K0B/CA3/yeGFctV34YvA+gYbPw3HTDLlIJriKAm2+Zp7AH520V
NKLOsRU2xnLkHaPNlxFt8vhpeggeCrm/tJiMdaRjdfCIXFAgpkWh1Rsdc0NdZdwv
aoZOnrb/VHjBk4Gsd5rabfIjUZ5i2aOQnEaA2Hk9/Qyk47DAflhW+x6anaCecfea
Oi1r4ho8Tm8IaXElgWMETMLI5dW1McjHZ3+E9hE9wkiMdTkmp9hV+cX3frWzSkIu
qvRZGntuYrn+oNbSQ4D5DSYSr9GKmFMx/8ndsbwXLxFngpdtkYKt1H+tnuXY5ye9
RAdMxqe+eJadG2SahtixOY31aiJE0zVSmO2BBdfKh+dWtkftjdmELnhK+CmXYO89
UNziRwQ0AvxBnFJKzulE8hg3GBoSlZynflW48yjX4C5N7dv8SRkHHGBhtv4e8+aU
OKssjm/sZ9CujatQITNdarJcGQ/ZbOUJOjGcmHQN1J2lk+26AwOa8BjJmiDVL2FO
dFvBat/eYLiwuN9MSRcJDOtn4CXew+iD53zdXAKNfSr9pBWjZtWYCwYgA6tlPxEJ
dBoO3EFhuYpAvvoYfAiKZWu3czDpfFd9iBjAk2YPIx/ssRfaAMRK4Tvp0kicLwU/
X8x5gJb51zR4eOtl0SL8gBafqeRBA21KN2AE7fyLTPZq40Gr4h0J7tuW8eHtNuX+
VJQgDH+mkaJJuxXT2jS4g6nDU1DzeJlWRTm9i/6AUBboFJ7Pvk+mMIsStwUQtp70
xA6y0Pz3udstI/vumLot17q8G1j4cDw2bt/e1PC/HhnXuuEQnHhwpz3eQ1eElTDU
4QF4b5jbk0ReDvVjfNh7KSJrRapr0rOKurzUKQJH7ogMd6bnPO98dqal/3PIjrEq
HIElem394xndsXtw5ywt6Th0ByRMU0ib1pe4zSx//1f9OR0fRD5uwKA6cLFlrH9S
yXiVsVrjDjIL3BOZYiEZYjieKQwZEzGxZmCc057CMYu63fQaIr09J3Np4M1O1IKx
2+H7RvvBzJu7HIS74qRVqCve+sJKGjfKSqK0eBtNHa7IZTT/xl9mdz8TCb6VdAS3
hgGa3yxaYt5yu2Q61gIwytjA6wh3jPNEh73M7Nzd3XZavKq3zfUqDkP+TDKSLrta
8meaoFvIRDolz/h2OXeBq5oEmirqKTEQ//+C8i83BaF6JW0ERPVwsJaJomiHNUaW
wHhd5SNPZeABPSTZ2ekz6paEMa8kaNaQ90KuDxTaBzo0B+0f7SBHRKTsCkqcjspc
J7qj276YenPvLqn+rA1f+8MKm/N+7glHTkEAk7ZD/KxWCGX8vgoBBIR1e88B5oWk
mQXwJ8Zd1rlQhisEvkG0czNCYkUaJbYLn3eW4ufQOyMka1V/gfiHy7FbjHNCmiTr
iWpbqPIXG6JXn6Vs9y8OsO+HTUqXdQbnEwVZZM93YzrU1ejZ6atBzsGLvQSeADs4
myRhBAIsayCyv4m0rLrXfTYHrzIiMV4Cx9s4FrYLdYfWKOnUQhjJklI/DbHTtb77
/tnrbOxDzWc186yhATosJXV9mTAtktz9Z9Xf92byaJymU4GAJRahvmTkpk7yimYW
dsRfHEBUU47p727Y5HBpZnmyrsWCouGl47qWnOhm3a8GVGQ/DSyRzyzRWgrEQ+z3
I1ynKQZUiTFyikXXa2/tDdul3NiV5wnKgTCcPPbJsU00EPxEe/ZhSsxmf51ocolq
agf8r+hViahcy44gq+W/uRRREgUNjdT3g5650t1IrUU5y1QHjqSCLyqIIqXF6814
LafhhjUOLwBXNlEko652l/JN/O1vwGCGoAfOTQl78Xk9H9pEbBEs1AbCQHYZ5BPE
AffwXkZlmB7anyR8cT1NWsU0Z/luIX+FTQpkrqzfogjqpNb/OwtD6pC9wLp9BjG5
Zkv1F6MZBjeSPJjRcH5UUcTaG08qNbwu+zji3dJ42COBgkYhQlsibhlb+n8gz77L
TWLI4zwyKwhkyWU04amHGLGvPzlt5INqR1x9O1qAdaxFMaNoHRZET9QPVJlehjwD
SktA3qhLdwjTrotec/tKb14JzDlfz2ic4SfnzQj7oOsQrP6F82bs4gCfUv2zO2fq
Y0vAO+al5oprh/ZNs/BQt9YCjESryOj8rGkwbcYPc+aH6fK17iYUXYR26CgponLF
CYF6umPfFs0Xiy404UMzMh9GAJHmYnqXs2OWwwN6igzPM/2sAdunbbT+xj3yuNPf
+bJMudhBUD/9AdlaMI+qkSH0bWDXT2sLmB3d6/l9OJYISn5tiNdpSnb1J617E/AC
CkrS3Y9cx8BVHY77Uw4W6w86g7ELciRplJicRD3w1FZgQKV72KNjGUhL8nD9BxZf
uW5ffSn36JR1G8RBPuPwVUNXNRaRHMkIYvalEHM3K+0qaUPYFSIIHLKB+4zWdIqw
aFTiVgnuDD8KC25Ws34IPtgkJFE+S3eYUbGpVZ6FtHaGb1vEwbP7jNrtxmMpbNWB
xOjkczGTXGaQODmkejUVQcZ3rwFbUcrZ7ABX1lkCvOCPc/CcUrzs4Vs+S+8UA1uS
ODyyUJHknmGffddFpCHPFzLaHKkRbxXW1Qf2sS8Bs6lto7otvO/T+2QhzhWeg3jg
VKH0SaBEDGCam0QmAM2yUCNPNS1HlfPkZ1j6W8B/db2HFLEt0OjQYOVwzPWufedn
CJn/W/cBIofLvzxsMoCjL3quCrCPSTrTHEcFb4tHUpE2rDlSxs8IZac0eG61eDU9
CQj9XVmRv0rvWTn46Mki9MIlVbfEl1/++8o/aUIcDxRYz+eXVv+VKHE8yQld1Z/o
e2D7U2iWG86/s2v2uPZKgI/snRjK6j03w0aGLIwGXpCOdclMlldA7IEH/26PzUaO
VjQ3vCOZL+GPkoq2wsC8CbtL/XE8+EhEyF3IPiIi33B1PTHd47fLOyssJ4/Oi1Wg
7htjnwqbjooD1i4UCxT8403wpDlmZXY/Is4cK+bl7wMANBFU210iix6FClv34vJW
K2q4VAzSnIsQwCT2l/XnpXM+Yt51RZO3TlCRQrj9YbWV1SjfiIY8tU67p0KBxeFQ
ORcr46AgZpmI5ZkwiIT3wYIakHWoK/tAr7L3OArGu3B/E93yVmw/QhwB7dI+MhWM
wuAbl9IJBM8LsV6P1A3iLkAYmtgQ/3cSikmA+7/AmSxqel51CXbvTLQQU4JBuSsc
L9yMyj//QKSHEjSNWL28qoSabZrhB2VDyXYCHzx3fpLwxA1KrW/FTJUyDKux1Hal
DKOmLwRz1TWot4oHv4FzBV5S+2+3zlTiwVGKZ777WSej1EsDZUDSIvGDCH9t7Jil
pXDIgFK8TIwib0Ysps/1MJj9TD6l98/aVqx1sMaOWpA60PE6cy1fUstUkepjJkvS
HOsVL2rJ7k/urHT7CuOpbnYFuHVoIcPRM+RuWK7pqifNuaMnnT9N/HtAHHISJvke
SpvNezYPdSYoqdzuDOdZbYvd4CXl3RLDl4dIapcA3Tl5aGw7F4DGTYwAMzwYrva0
qV5XNpMHVFGPASA7qHyO0FlxAwCpf4hjmGZFjnfj4rHBCr5nQrnBx8XzONzX1EH7
nJL58qCPkgt9h3Npv72dEXdrWZl3AkORxdG3J1ZnnqDtORoEwQjpenpbgh0meCQU
QIoSKyhtVr7vp1Lu3IRozTfc341IceQ73YHLZmXOsBGNAlYuZSiDc5RBmsWJdnRy
yepSShOwrog8XalRv4t0f+nmsmq7aLpLkG8OcUWg57yYOVQ4eABuVByCB8aAJpza
FfF3OT21kG0lq/ZBghEUY3izuWwcGFeo9WaApQqUxypyvYEwWGNcZCt9dsaHizQ6
0HJf/6TvhpMaeWjVm63SIUIajIl3TawUAzJoq8uPaG69znz7i66YKTeMkV2ldM9c
2M3ZD6qEpNJRQCfoNBj+4wZfmyfQhe5FedD9JohJ813NG6knb8RfsI0+gQXvBeRA
TItcmo1FOci0IOCe2rCEaLcQGyFwGE6jpmVyMjSwbEXPCeTFSAsOkscN4enZm9QZ
SZV4FfMH6vwYPaSIstctpoGO/bMEmnPVbcg4PjsirYPLuuZ5mLXR6HJYG9cub7/Q
g2EqzScztt8/yJcruQGKf12ejuRIBlHV5Ow6FRuyYultzNg3N8Om9Tp1tiLZzcDR
hKYtFlzkYF6Gv6IclLFiySQmP+Hy1QX6X4SqDkXu/9CHo0qU75ISkBVh6IVvjwdL
VN/IAXtkqpBIiGZFKFKcBDNujKQoUafijtrCXmWtSAS69kod5DT7yPxSBJZdIrEY
9sCoNA1FPjw0gqZKPLFPt/3dNhq+No21A/3JE14qEBip0xOEaDLsvcbffVxrVkYv
u9gDv+nlxLXwGCAoJCNLqnNbSBC34aXOVeM1uHIcKl4VvuuUa8WiYZ4seCFIX//X
Y0lrQHHI6gMz8KXZ2cUrXJqOQpzvtsq2XoVkuQyn1OXxK3NUc4X8pycN/EahpgEZ
WATWEuf7m6xKZvmKet57yhRdksWjDx1EyDhvsDAGye5OsBondbfChCVK6e+AVIik
FIUPUxQmgc37iH3tBXQg/cKhfH+0IlIBJimrlFbsF1QVISxRQFiKi7zthAlzv1P/
XA0t7U1fhKTBIAHv8X16hj6Ymln4pb5ao+XjsUef3qdRqheh7GhZ5x38ttW7PlHQ
PZGqg+IrAE5cWliIVwtOIWCkiJlfJQOvJE2sOeBf+RS3ge2lZ3CvfGu8uKz7l2Op
Q8MnOir50uwsq/1O/okgiPEDcwYcStkto0QCkgP2zxq2eECsp0Bt6jAAuDrAE6zJ
WriZocbzYR5Y4FRvjsIyRNc9/big6CK1BIRpXg+tDcLaQJYK8eSsYGy5pQrJtAf+
W8cC2fDOyIG8nGpfwW1e61uGFd4ugk7797k4Eft2loawr3+o4J3YMLRwaoQje353
uhidfeb010UFh0C5v2gpu6xC9kmmsQsGafrB0an3fbDm3yF0lM+yldof50P3sTtY
Fo9noHB6/42P2NisMPFt2akRHQcLwTSx8mqOthXit6NEi+xlssSFx3yOcqEzUuYQ
89oihQyYQVmRV8UNmyGvC2aUA42AqR143WdTihXJDsRIAHlkRDYkmmVRioR/zMsB
Fk+3dqNA3yJ4Z96x+jWCJHrusyC/oFYUWz60jKWmyt3R8i4Qu3B9XHm3Mwrmpch9
xcZ1qfDhRqLzubPLFIH9f1Yiu7e6cFIBtnocKdKK5lTcdqCspH9L/C4vfmSlFBcT
g4lHuJl2LD8OXzg7tm8LkE6f5Or8IRx4ipRIGjXaSQu9DVLyHxJN9iM/6Vp2Echj
DrdYJfJFZ9BJwGBu+vYcFCx7wqEsfmXMrKp8ZtMJSNBNn1CsUdx9Fo4qZYMT/FTt
Q2zZCAt+deNLSAZJEGySr7tW62r8KA6erNxFxE2E7Mb6Ue07EO9sGhPVjnZHfHzF
nUZqInOuI20m9dyHV3cP4YKNBWOOWRaI2IXrSpNwYUXfxOVRUvsBdxjfBehDsf+Y
R9/lzTZ5cfWk2OnXjZmZEv45RR9CQ7xY95Gi8ainNgyCTyAwEHloOBxu3AvJSMqK
AJA25qk+5QDFK1WN6OfiuGNRT8G7VIjsvI4hBh5pjUADstx3RwwRk5i9IBe2x5q6
w0slOJ33oRlFR8tnSJW16/ZaLESwzZClnP28QbsZCHpu5IiH1OC+9WUEssXzj3Q5
LoVbrYiG1BaCI4Oy2UBwvcVQhIF3t31AXqYibo8zFYRLKD+A0jGbNsLPNzyX38qC
xEInGKd6dF5qzvY5ZFtB1ULgH89l3VxoG8SaA3d44vuMkJyc3Q3SdpbKM7Vc6uLj
fVr94yhHk/QhYsdUOtBHKeGjr4HSAa0G9cY0zJgs/FODLrg2uDakIyrBygbTzgP2
3x3Qc+wYFvkH7hoUMHhcs/ODA/SjCxQzvJ4lt/Uu/FlNGw6z2Yb7C1+GkR79pD1C
k3AkumPIw6qL8aeGIFQ2EeTXf3Olxx+bH2endCIQG0qEB/6zFiVKmtH7N36ted6/
AFkk2CgB59z52T1OyZQ2S4LEvrsq1Yt5QtH7YN4tCDcamR3k7maZe/9uKJ8TVBDm
XZzl+6WLN8UEtfFGbXRHYpITPSN4aUrcGSyNTv2cJefCtFdgedDUazYqvh54WmKl
5OjnyQ87grwOHC5o4FpsJ3PZm8owH/nA6QWUQULPDfDIHJmIsiFrRODMavxftxKf
MDforvO/H4tJYe3eLQ7mBUVxAHChoEB5lH2EuzGfFbcZpEnEAH3XpZ0nlnVMalgY
55CJTmGabADFdeIGD/otQke+/TEEB4bvQhRK2ynoFvw0KgcXTAYBFumsRJw++dnj
FqFhqjFDd7YNx3/m7FZeU5Hew8L+aOOWTDz2RjQWSEsikEeLeNrSXrZBnIFfqkA1
APPlWWENx2Pq/rfxfZEcFRNcduhWPEO+yPZ92RNOkEQUdnwKTsgP3WqILnEodAlu
UY8BPyZXGbGGVVJ1eu1owhO8yFXklBTWEEYnjj0J6n9/8NMg6t8LCmMyzrA7GYNi
s5Exv4tUwKlAM66k5h2dF4NiXVd841KdIOgcUcsHrrZyq0qTKJ52pS7lGBb0nyNP
xIYI54JKjtAfC3eObdPjIuFfgErTJviCe+EZiosrBPEcFjF/5VGz9czEFJu8f8nt
tLZIR1EXBjnY0MSvwrp+d0b7uxbkwVh1N8EWLqhrq3bcegtnzSKSZ/3Mm6AzMtPl
Bbjc4GsrWgnc8wIK7JBq/c1kK5O2NOo29bV7mXqmOMJa/TSMdjXh56OpXi70RfMW
r+NCohZ0nV5pJ4AWx5HPciUDwC2s9qC5QXcJ/+pfOdVP5pJmxpI8OqiDri3+1BqV
NuxPSnEl7TdUJ97ksXYxNaI4AQmYASNa+txImznp91xO9kD9yOP2RDpLRMs7Gt9V
QEhtEMSye1ckk2YguS0XJfwjpZPUm6zkAtSt14j/InLbpG188+TQtTj4pppV03B5
RcIxEFuGOppvOMyMx5Oq3fVGb8+vs95jbJGRzBul03eehS91kNf+qoD0Qw1NGaea
GdhmNeK81Q3hHXMKgo+EPNKeR4XwzHG/H8bQ/ZYsfgX9yHt/+kUHD8QKcN6e0uiC
g/3zqDBGlGZy3kt9yw0jdXbgkq7HCf5XwEVRpmcZOu11YofS+ouEQQXwbhu0eYJQ
XffLOCJA1cECn1EdewBwoQxJGvLaCTBT3X6kt+PG/1HH1Vf6fmEV2imN8oh6T+cf
WNBFlBZsF/51//g5VYpxAf6yyI3uH+6QFwHRDDuqQAZov+hT107yBsXabuV4Mla6
rbYzTyVXmETigwcvDxzzXJlbbtVkJdae6lz5PqL0AV/N/WuEHK8HgDZSrfVyphuQ
eCq5UFgkMrMiljtjVtB24JnRCs3+sCp5ozyyXcAX4UkbXw6v/zfA+lcZ1b3FgdVj
xofPrtIEw1AfU2NdBlmIotx+lnVz/DiSxzKu8UgEsMuC4l3MMKCd0KdRpRhGaGkw
kOzoyyAb0N4J1pMYnDFfS29r5UumzeSUK+GGQQlEHKC7qsjU/OsLkqZsUKOFpVbl
r4Bwg3SDaHXbaYTd+v/oy7nqbYlY10F48UorIPSAq4K+7RD6I3D+jukTRcKYAMs1
Q2VDyU7IiSvtzNRrlkqJSVVyH8/xUAAf9mkTlyJ9j2vKEJouBaa3+mJxZiMsfqSV
4rIkGJn3Nz5mRvXa6NtCyWbX/LeSZDVEBFh76WnuloVMa6iL0gdN9dN+X8Yb9/5b
eyjQN8DQNopKZGCF7XAIfbif4Azo/ryZGxSRuG+q83HSpqDNBOC9UeJiggvRojv/
xl74ZjevD8WTmI/7Nd2PUykIgguPicGUbGXPu2fvczSxiTRr20EsELPXmdk7zP3T
Ko+TFGNhZHYRCknEg5euO10vbJSjjHvJo9dn9RpUOdhh+gvr7uU5fQ5PGlTOQmJ/
G6eUdPviq53Lq4QN4n/5Mv1RxPgCq/cgG/iM8bH+Ju1P7sQycO4Y32tj/cffj/ax
vCVq+Ue9RcMIorHc4+/l71x9l00RGjXZyk4ysFPsajqcPIswliIjE8J3UesyWvfH
wgvdVZmtTilIgA3ISfueeV6w5LaDOxbingOlbPuoJcGcQFBBxvfVQ/pOYfDGxk6d
pGNzSRUBlCWg5ICMpx7h25Qyv4KKTXsNJ2MGcQtP6IObbzqd5oMkAmR/HzelTxnl
9k1iqSLZw4t2ZceyhP4dkeM+ASM5XKoPMd8Laop3+a1tywA2lcrkuh/vJdjNcBOl
v8jhnx0HhZOJglYMLA/NhpLfyC7RJ2qJFtbse7YGYRl4tNxsHT/8Vm7xseUFz+q+
O9V9rQvlV+7clLmz/8KAoZnrh4NUoZlWnPvHZlh1xV5SaiRlEe+x0cO1UtLH6k2D
Fi7cnBuQr7mUpG4MKFajWLyg1NwXk3alsxRiJ6tnMZauKi/VcdJgU5B6Ie84XZN6
t1XxltS4eV7UDw+BvVfTjUIM9th/p+U0xVQdXdQ0K5l/5zScknS8odQF5S5K+FPX
jn+RCnPrYTRKhEVuVc8Pv3MsNasWLIdwkVtbNCGft23HL1uCas09kYeFFCNz3CTd
xcp8OnSrvzxv/APyk3hw2JkXP0DxefoqRlQX+EmITQo/R8GJ/e7Rj/3C52AyrJfL
72b7TI7LdOmvfraXhWSSkFcsRJlJIisbdqow+JPe0r7tZg1Cr5soQQI8ISSLx/xk
95V5pjHe5XQXnO8qdKNKbjI+OwH2KVChxrCTJaGoVSgLPnpvmN3ZbLKhHfZlxXMp
7LJ34PouVLwactqVtW4tJy057K7wZhHGbp4a4a5tX3+zBdFp09ESvDBGAfV1uAHX
7bcN9mLeEXHGxMuEAhBkANTblyWkQ8U6fjU95LQ9OOElR2exTaBld3bADMVfEMvQ
2IyZDG89DSPDaRa7ixz2Y98XD22RK59iXOM1btmk+6cb0ZPXwZrIfNHTjLvW9KxV
f4XtUVbbxkfTNskfFEjN66mAn8Gw5eDnWWCqaSDhk4obFvKZZLAUd1II4HVssrrP
ESsgZlPTm75uA+xmjuqOyylj9DxpdR3DHx3En/NgyHpH6Ni9bvmcQqkp45y3KaS6
ZhvRYbcfYEpurUc7iRLVyNrxfN3WeGX/sp7bBnclQZIrY7PKIztE6kIxpHo+Ik7S
MhkSza36+xOqPc1YtQmxxYGEDg+83s/rOUU90rFZ32zu68jk1zFtMnNqjqiSK049
wVB+YKNjD3jO/AK6La6d0db0GkOaQLEOydvN2Cf1ULAczrlQLANy5OKskq4vkFn1
wVhFn0OrR5calMci0zPmyGgMiFmzrVbN/pledZxZbZI4Ll/+C8DE45zGRa2V54L/
7GpTBI33c59i6ORpSuXfwGvaPzYtkeaSu+kKyB0pD1PiT0MlFmpytDKRkqzyIME4
2xZ7HovYML1IMOhQeiIyCC00N/CUW3pbBShgbdn+0ciFTDKUoRxAEgy2GeIZlGTR
oceFeamj0uFQhdpNqk7QFBi74ddbh5y8gnIVVCS9zVJC7VLsculksjY+rLP/EKCn
4rGCjYFtYracs3uUz9R2gM8TxEj/V4hkvXyDI1yBSvtSFgpqrD6DFWFXISLdxvzh
xEx7cnCWSmMvW0/94Zw8ASA4O4AnUVpMxKvAPtrlwS+3+GI9um/A7Ah9ZNT4bFmw
l26UCyUqkDtGbY2QTKe7m02fgV5X6VHkdBE20VrUO1BKItDHlm7QO3xS/6wNGqRa
QrUMw+LpCi/VXs9yYRmeOzSLIj+8xRqdkmmYbte18NhU540k1NFy4gUoJBJEajx6
rv38QU0usolYDT3zcOjrf5+o8N4eeTtSAbdrVCFH+crQkmlKj7GDfUn6ZvCC31Z7
Sq4GliV7WjgFi8fQ1Pc4bBs/tqOuOrZTWA9eY9/Vh6QRpTDfMwiaOuAZHwhsXsp8
dxEChCX1MdWvx1PN5zxhtOPzDIEoNkpvN4KF2d8RcgLnplzK/mTRwardrM9Pm02e
Bdhg3GN+nFrj5JXQ+ClbjLnBJObqM2Tgjc+ueJF4pCVY0LY1PTtGi0XAKiGj8n4b
fWwBIAISNBPjp/9m/yciKLcfaqsLboODzwNY7DtYd1BEYdwBBBqqZybGa7PgUw3p
j0o8rNTZPxsQzn28vmZdlCqHXUCmOSnjpEmYj/+a1z7iwsbdHCDhrNlywnVdjJdG
8ojtb8sdMBFghAJZ9w1mMpLbJTA2MhEcBe19jDiiaZVdzYTZbEW92VxMV83NHqCe
N1wER1UyRr09LnWxFEt/8mT3cgyPupz0l3/SviE+nSGRL9YziipiGELrHGSG8cFa
+gdTIQQifEYKAySZe1Js8gQ4VxMz0OFa091/mkOUOMa+LWEMm3kX0bgKwCFAEA/Z
NRmFAmtA0FY1HsjuVO3OHFe83CI3p6+OXHZze3PA1IBYSZRVayF1o0Lzjvgii0SH
85tWyGT0d8kRLCh8FlAD36iqZ5bQYFe95TWw3DBj+goOTfGXeRIYQ8zlN3BIZ8t+
rnEx9sFNZErSdWhksq25mk4bz8lj3zcgNDAbUsbbGmqGa94sf+vPJZNHPzFTClG1
UHtY79JeczikDMksp/n8jb2DXc7V8F2MRBZCSSSZB/VDg82r5c2c/+f0vfcDOqIP
kSBEOMkp6OFakPVtp8KEoutN9YU/FbiGzpyMhDJVffZgV8eJdgqUodznF5m8MEfp
xQefOmrm5rFt5Wa2Dq6xlrZHTXHa2/7rBKhwKda96cbA5NXRZ2SDF9eaRXoAECcZ
RDf1JKEYj/u5VGBa5m5LJaC9gETTxexX8yLUY2O9xHj++5r7BOnmqY7kPeNRvAPk
OUYbV5ENVZbtiFK+7fWxnBPL8+HNR7S5dWB3x8d3UWI9XOLTkLbf27qRFS7Y0zqx
RslCt+TidBCN9Tjl1WXjxXCqyM+dXINrZ4I+rbl5W+ry7iLx++mnD9KPwF/O5NSW
1XSLGuEexJzngo1xBbvMz5fIfZvO8ujZk/gtRe4J1ZzWK/Slo4XadgoU88uIfi+p
uj8PHfdivgagfGqa2NSK4jyA3cUML7Ah742qzPccfkatI6smDU848PuDbULQqamY
YHUTnS05939vBO1fumGTGOC/ihPwehcaZPDQD3nYvNaD4Fb4/MEb5uy/I/8Y3nBQ
yF8TfwC4T8AYycvk2yTO3iRlC5Gew/evqKQgEkLr3YaIltWrH4wusg7MVOVRWVZP
0t+0oTiigD7w9GaNOSBbWz9f61wslR+g4fSq1kYv1Q9Bnomfin7PCVg2a7Hrl8ib
5jus9Ki4Rvw9YD1oCR5e93dxamK+cvTuDqjZszN9KozoD3XSEX9MyzQWJ9Lnj304
2DK+2FBSA4uqu10s6BgWdHZX5c8VZQEXzPgiA62intzoAl/yCvZzoCoO1/j2PBRj
iKXYLTFXtqItXyq4E+qSHmusSZ6KojH3av3vbQaWC0nWCFP67GApU2aSF4yhTnai
KJad98RVWFXyy+awVxRk8w0NyK/oLVVI1vj12TS3NspfdA2+9lpdK4Qa/toAWl13
874a8brK7zb/u/eD7KcwEJUtR7Ooe6/4shos8/Qg36akW89JtKGWqdpZ3fG/0u+h
2F7PE7AFI7IHiXCfYGaXvQqALAemRltXGcvVh2xQKld8yUcFcW4WJ2AMJZZGgMl7
xMLCj7kJ8bynP1S9/OqDknD9Po5pA/A28gCpQktWrxbTFknNdWRGlmCaUZ6DtpwV
roTccuiFNeJvUt93ORrHsw2FNSm5C3UJD7i0Jq8SVEXL1CMSRCyO3s0aT8vvV930
MdJoQeiFVa8MO7PhGXWJExLeab9TWvGEu8tLBQsZ3sV7EdYbUwZ/KFrcvK1Ge2uk
W9P+wrjHJqm1Xl9kDOvF/1K8L2wGTnIv+bGDAh/WbhLd9cg78mx+oKJmNTQlKHlD
i87DhdC79OEg/p9IXFLYp0UH1Iz8Xo0+KVImAbNAgPlIUidS802rtqduWNjTiaDR
jk79/253c2XhqtLHGjp1/cxW8N7JD+WsKj5ic+W8NjCDU7WdjDzt3uBzE7l8q2T6
t5OWRiSdKwVeX7occM/QXZNAul+fcJFtHR0dy/S9P3cR4plZyKBeG0GR1lMtd0fe
MRMqtkbyapDXUGZBGDrqF7f7OHmQpqOCxnACR3zm+7YFqp/1qG8hyfUnUdiPKW3C
4YPjiNt+vsVuQsybF9Uxmkq0MdvI78FPsUtYLVhBZBelXYGfahmB3LhCjtnMWxiJ
cTOWLmJxpaXxqXtTqgV/VNvY7YZ8mIjWS4O96Uarq7igL3XoDuYN3K1fiNZLTLqU
U//oeBkCMbj/eB+QFYSmkDZZ/PAx+y4+ZJCSrYWZWorHMT3SJo8SUTXXK+gClkWW
32+QzrxaQxatrZr2kzIiUWr91BlXT9d31YxA2/sh+FRR9Dzbh97NyI1vN3sN7wdB
n3QrNKhR0KIwGPWCiyYxWmAKMDbDowfQCO3uUKqDfUfdyoWIoihzdGqa5heqRNif
2MnO2QRzFxW97k9OhcENpXKUTeRkhFSAXNUZOVmt2ykHewHuF03GvCUGORRBB5c5
G3HfxsolKxOB+9ZbYjfseCELj45Ni/ODbMVjQOEZnil1oZ9/nRI2txgOGM2kawOn
vgjpv2FINRUzkrqE7bbQhExJ8D19mNenoHFNcnWtMYLaICDziyMz7+sSEvLyUAHz
AR0wxWgP0b4h3G9yi5ZL3G96s5KK2yf3cUug6F41wSOsogFTwm9/JqHl+M2LinQm
gisCEI/ysAc0OrWI7MABubivibYNlf8ebLYHBy9C5DCG3tSmiqs9zIJ4jEznOtYQ
JGd0eswJ7dr2DcVv1vZvVb4qtYLnlQB4vN9Ncofe8+2EiLvXS/LLFHk3e0OTitWY
036AkB4vf0qawBKKoGJ5/6xheI1A0WDQZKgGd5P96Zeo5emYQV5u/xAIf7y5kQS+
LSHONQLFQT1ZUeaUrSoOjfR0zfdzY4Im6GPSlnX0f7WKapuiD4fYpuvlhqhwgGam
r1N7m+Y8G3ALaHZ7CtiyxiW39kWjjKKw2W0PcmZyOkI0R06PjhG+IH//3S9b7CFm
5rYFeWbJVWFJdr/iTGrxPx0gVH0LuXzsi2g4R6ne+DaVcxrc03rRWpNcGJjDA0ZT
d9V/DWyv4er3RV89+E+3nA+g/vnLj2rnXjceSS9Yw8YhEx2hIlsACn+CDHslKK+2
JAHBztAXvIIxqVlemEOdxWCqztO6b4bkePhiihKt68iK0NYcruXaTWki4StiWW8k
y6655ShY1TNfzzmKzTOA9BbtJsiAydbcdqgQSiz2IuJuz82gU0KEyaUpnh9Lh3O6
cN4myyMxCeF0Bdvn7OtXPdzlGARA014hu5fUs3y1oeuvsj/f2h0lUtk1TCoN97rV
EPWg2tLBWY1aUkFf6FB2GMSsSYX8wo7bTWkQ8alnuLMuXW5XHT3u5rKZdiYPF/CF
jzqpm1wncrB/haj3SWTbKSaufYuiF6CRTUtwim4rP35MSrVflwRJ9Q1u0LSv/3zl
Fjfe/raxY+UnKIOvFTp5aSHn0ny4z7FdszBXK/ffh9Mi2RhTrlcn7ZW/XrokMCe+
ZLHtvh/UQP5RmA0WJY8Bvsvy2NoPLDZAU4vlZU3KB3M7tEDfCrScU8OQopZje7w2
NRlxrS3Xph81abIE2pbpWpdjUEHD/PE/Y8Top8x73mAEq542Z9Y5h/ak0sojEIab
3NTXrBtS5sW4FChUpx4bMzjEZGG64Uex3dkUE5FyIi5chXuRkoI2kbO8q+FTs0r0
0x9ga6Qjl0s5VtYMo1nTKkZ/8xm1DO53gsuBqchuqLMofllP+74VYYAw0MoAyDro
DTmkaBqMvo94emvENC3NSpMlXiFxU83dq/tsPXGS0b4TcCZ6d99RFHmDXi5GrKqm
yr73+cHxrLI+YEqDSYvLXD6IVs5LaKwbkUNQIB4/DVpLWcdBj2pDL74MWKfXmfAU
gc3plTv64jVxm2Vin2ESFCdI5ZKSlA5Lov3Vs7LxXWFHVVyNUGwo+NB67n6mGnsF
0BV+7LdxKcFbe5D+NSaJCQQLmD4SUZpwBFxT9YSOEh7UrxKyQXHWuB5zRew5EM3s
UNgJstJNYGrGnJJlalVpPHNe5YsmteRo1362jdD5Qey0oM1oLtL7Fd7KGuvvYPQ4
Giv1xECIV4ZlBqic6nClHsbYihmogui9DBYNgVQA/XH2wH6opaiRtFbZLYtTUoYh
CB4giZx2U+ey9agx8g7WuG4451JBHQqmRDWXaHLpaeWDCAbVoZWlDMmJ2F3VqaAj
bC5vsHbnpBegri6mBy/tUMHpXuSv6IdaItBwR4NvY2zKWt2m+HoWmv8qCUGrq9fi
SM7MZTTKMrHgfQb2336DXnl5xLZZBfkhrGh6tR/pn04ExD+gE0sZBMHXZgDweZjJ
ktnxKZqTnIyCe6iW9it+Vz6GbK9n6LSvK0wxqim3taiqMpEeQuJ43cHPAOs2BG7w
4hWQ5Eg5U/L/8n+TYSFczoSdJUwQy/o5fnLNbPiXjBG1RqPKqYEUbTiIXvHF1/nE
RDxry0u8sPryvgKyHHdW/sCoirnRpxxMEfUppdFKVNvg6sNV/a/XFJKCrF0mO0cc
/7iaOk+7NP+6GisvMeck/Luucz5TA//OK/9afF2JShry7l5yuqitSyNUfphd1LMw
zhAAdsIRdtcGXQu1erJwNs0JeRfITz0qbzRjYU1lU5nlZkVcSicks2xSyFA3r/ih
BmHKTRePBEnx6cr4II0loeO5loLM0YW2Qp+3ODFQrE5lv8dvh+ZwmQX/sD5cAYGc
42vJvewB7B/6E7GSYC2U9LDciJCE1WtW3G6Mgx7bgLV1ldmy4erRK17Z57we81d7
zknUBaShAhmETDptJAOIDdkak1pQsNJQujrePb1TnBQs6uN/3PFM44/KH9e6uYsX
+WAgOTZb3GZnOkGRoJWxJa+nr7GNZBGoVGTfMsKW02Op5s4VSXqmImvGnbQYNgJm
nYxQ331tH1rwtpRNEowVR0VzTLp3VA9LulDv95qaB8A9XB7zhlpsDgzzuISyx8vv
Odr1olBD88Nh/A3x2UEojAuihT98Ce4As2q4ma2sjTFkT3BNdFK0pEXEnYAnHt//
EK9+upCMoJIz93d9AsWPGLAfpkIG1Tb2TuKSpZz8AZc5Cp3WIjG6Nz1nNcTrJElB
LQpHDlH0tXS6ylkyshrTyIfD+Wun72i0FipWRIuDtY7lWpkeDZNIvUErRTq+YrhY
z7O2RUMN+RPXwoCGn7juDIbEJGUlvpZWfN9z1Bgz0tMja9wyo2ajaRiMjf8bb8qo
zho0O82BjvwyvwGLfbIaWxJqzODGTQrM3X9n7dJIn290ncOodiq++k/1DDPIlt7D
jOGwfeRs7Rq4tzDaQYs9QmWHVJdbv3gr5XICYWxSH0kD0/OaMC08HF7FnrzVXbGO
fzoPs6F+Z7PB8+EOgo3673gAdktA5Ki+o8oTqiYAMWXUQp4expwLwQI8Mbc1Pd57
5bKwj/CWY+1E5oSFdWIVSgXXkR9/tpVVnsLiKAnEAOZPqLtCu53SB8TbMa35J/od
D57tskVasAHgLKInidBQkGvtZUzCFiQvzdJOG+0su04LlIDgIf2RmAH7hlOpERN8
NMAFo69ckziWshkquiFEs5FiGRiwl08K/q6JGh66C9YTv9XR14PRg2651LX13gAI
KwGmMzGUoI+axypnxRg5Io6q3GGjHUKuwDVga5Dx8Zh8d+lBB9/Kr5XEOF9+paDx
ZttHVUqt0OfGWb7fIc3bMFOsA2DmUrrUzXxLrREuWMBM0Vv6LERgRh67NIiIp9Y0
cQDJcvhpQY9sCLQVZFFC6T9br0/0QJ9hlx7KnMSBXzd3VwiehZcwGzfycRumdzNP
5n92VHuOEhTdPYEjakRYGl3kpvsgdjSyqEes6H9uA+gQ003d37bscwYWo4uJe2Za
v9iIA52LPsunUW6ZZ80B2DCksoC8KMYRAcUCWXRKRt2obXBg5vQ6U0wm0fxfjTHx
YnalN54cEn9noyZ7mSmea+NC3L0qOUZ+r4qHiX6YUhYvgczY7nJH6qqJXF3NENFJ
HyDylhXxOOmBIZqnc8DKlHzau+zb7FJUyh7Vaxf6t5Q6UKYLiJYvD+nRLO+kp3rm
UWU6gTdVVjS4LEoR3nNTTIVkYPrksh35MLYiK2+tgsLv9LFlxNLwkSRcH5Pqj0OQ
kPxvoUHVIr0kyRXkdA3hYtH7z9MlD4QhCzuA90eDtG4v9mBP2mJxRrrLKtoOi2XE
AQf5ADhuAoxaC8QeIVp/Yj82u/EEXtZSy0jcyclkTMN7OuerYyVmcJcPDJu1AOya
7TJdJ+ZNDis75eXoVv/Ol+hEjnh2p8+z1f+XNGcIXrtET/5Zv0wBPobo9T58Kkce
9JIK/KYS7Vxh94dE4K6wgJJ7mrdx1HBAHltH3mvxB3FGobYQAx82CIvVi2/kHGyA
F4D4jz5yJnQJMcQXfJYtbzrR7AGL+4Fiv8/SrtpwfWPF+8sUMRXKK7mOih9Fwk19
BChJGZrQGBcBczm3+MHDkf6R33mCM1tmbjgzK+6S5SoQdQzIBEqBG9ssaLwawM+l
6l/npdFg06AygSgV0KoC8wsUJXdKCgMG2F9LMJMPuW0VrzCvaRsYXW47hX+JP6W0
o6XW1bemxPRDSy/EAOc9QiQGp3hsxRFGiJ+ylOcsrN3dDUWEAAo6i6qtW6rU7Npe
KwCIAkxKKupYxfoks4nP1ZJA5mhrIlqNsarn5IyX6bbsxkGEWlIc7CNULdM/tEHr
bwP1AxaQLio3NtjRB4+7R5/I+ciM4r0qVodSMI/7G2VbHmQTGFUBQXYfxg+YvWVu
BBg+iJAu2Y77JIGLxCLUxcDhANJE05VZz8HV7tx/VONtcL+0UxAbOHArHi7RyrUp
blDUDv7s9TM74SE4wwJImIBOFfuemLZcy6RjO2+Hi0Qi32jJLUyGMs0vwJANWmKQ
yDF+Ar5gOHhhh1oeXr31j0sxMrsi1F2ducx6aHmPAJFnNKyYllO/jlZ0V9+885zg
QVo7Km6PRyfezGjQ5m37220ZyuLTE8UZRbspM4QmNaDTdjWFIm7yQ/duVD16t21P
302fbfBZQRGmreZJALtZwMC0y1o9HK4oMgvQU621DUHCFnQIYdf01cQ7LE6Fq17f
IQYKlavlhw2OrJW6azaK6XCNBRo/RMOltPBEeQFn+c/8XpLY9fysXvhhlHkFZQpd
sITipCnBm/pGmsDGHnTec9Xu7t8sdmt/7tz8F0i8Zeb+PZqqnHNOJKsMs3jfg+/m
Q1ZwvduUJFNPkvYZt74v9vvs0oEDe9IwOFrRnVynFctRp9JlsL/CaiQ+jpapVTVz
2kXRyEP6sY10At3GcPhwohJ41LjQE0fJFBOCvRN5IJvItST2eM8pairprFpjof5J
6KV/2oXgoDL1TuE550nCnf41y4THRCRDRhH4/fhAGHGcGuXQnN20K4UoA7vm8RmT
B9HqySyinCYtFjZjNgjkkiRj6O2FP2ueIaKUL33z86RvWZhb0hwxMzbZ2miNgpvN
YYVM+uWaLW9IQMLT3RbPrqFuOuhq3ueY8pgAQU+F+0hwhRlxEBUVVcNGQOOEaElQ
9zeHYhi1WbkBGcJDGPcWymElTd1Roj50xqeWRc2068C0jVG/OkIQf/+bmf21VwAT
J9zagxpc9dhRvpg4ajK7rk1IgvwI2wOc4xhFP2qwv6ewa9if1aY4s2muNmxi8v8F
5sLiYyt+b3mUkgUMz3tFsgMe9N7ZiWY+CjvhIN/F8lYZsJBY4yqEP5FJgV6dJurv
jFpW5ZllEndiZbySu2rjQFwBV50+Jt1WyNgbTLTnVSRKBae9ePb3OCOimnx0Hu0D
fT9jRwppU9zizNrRIuikEv3HItaqhzCi39+UQdhaiemwhyDHvh4G8QWz+N9YtqM0
LUOiTNF7QkW57E699D0xa6ngyITHPTwRWpAG/qndEUv62PR9Rxu9GYvm8Je4eWJu
ANL6tfxux7K7BTEfZw9a/hs9b9heICiwpPA3Tl4Gq2ZDI7OYu1PPSPvygLDx9hXo
4fTIlH/rn3pblzI+91ECiZ1NMxRysHgk/St+eitEcECOEQHlpFs+8LM2JECtW6jB
yN5ADu0gBqnzO0mwT08ipPrh5udJV2g+CAUq3bpeVkMF3vDHbV9KGqirp/23vHLJ
XjpeAix/RSUoGjRoTC7BdrAbAMvy2n37P05ckfOWjOxxzkeZqfrrBu35UsH9mmNo
CUy/3WwnbT/vGVzPa93p6f8RHen18Fuvslv7/RueEbrTq2OkKxtxWDHz18Frv7zB
RQWhweH8WBfZNGqkC787ZCerXZ7jES0kiAoRWHOuysiW0vNtsH+TrMWp2V5k+Nzt
KZ3J7N9wv2vMPANe5mpkcYyWyToIjLSVdspeulVgVC++/ILV4yp4HIJWIbXCLCBX
09RBrjctE0uNJBjzcFxJjZ9ZJWaUDweSrpq3w5Gc1BbTPrSXUjtZgpUuHs+8PFja
xMn+JRirWnsIKdqpYbTSJjVj3VlO3VqJKAnVAb34SgW+AF2fT9a6suRWlFD1fNtP
GOtLowF5vtau71NfQ+3asFyD5jd2eBx4fkoR93ba5RdoQosj9PBgHefxPZGrv0AA
FcnJV38s4YxMTbmaK24MjWFsMUTuzeBLh94ArQLGsLqM5cjmJVYA5USewfLiNXYD
XfoccyGht54gl2nh3IGYenV0sTpe1K/qhn0GCWZCLIVai1OPuvq1Q6g1WSMuTKXK
hOVG8orzbIRePw5SoUQzThNfYrl9eIBTVfR3/Q8QyFew6ktIl4WOxQ8mH0/0441c
Hk54Dunx+QccYjPuhNPSHnxZrcXPuPMBDJb+CYNX7sR7SrP6qKPTUu5S1zZkGgfc
EYM9MO6SpY7qaTr0zavZTbBQiQrb2gWtjxyb88K9NOEunYy5KhM5MPDkhlXlS2Lh
95RCvC1PcRLyzZZnmfryHPigX1bTafEBOByGlXusUlYVxSiYLPB0rJAPCHHwiUAi
cknLoLQsUGyYO2vNxtI7WSycC0iMreX/IfoYH1GDW+4uCLTbwSE5a8D1KcysuQRT
mhBL6oCe11NGmJmxk2DXBeb76b8Ev50MHB52Z3n4poluPk+LHr0knDcwiKIocyjR
RmBRq3yPWhbt04kqfqoKDMfxPsDisUMCOvsq5Dso6LmaYFEYsOUGN7e5chZFr4fU
CAHt3pKXvT6z1b8Mnpx9sYmjJlP302obLBbp1Oe3iRmasMppDhvfAQoDdIW4yLGj
p9eTt0D+aHffYHo3XqYIYnrtGkzT4Q5z05SP2uvQC0CYWQB0arDOzBv+Dbu7yK1e
Y9tNQXnNX2TrYN5kIfuqfE43DpdNim5vzeygJKjwmkY1iexVUqwCq+prjGX1mrww
s3k5bsFhwyNmk0nYaVHnPK3IiU+G2lSCGJl25pqHySVnpi85t7vUe2rEgIuXnkZl
/OGyiia3W08wY9qgUMZvHLIk3jSaf1K/LazMfG8vHOVqfj26ZQ7EhxVDZQvy5y9h
fVPLajMgJSGqjhzTBA35sW6I4xZC2KdqFuVp4VKuUK3M1HxqTadY01FLvPYaspsP
LdzlFpc1I3LUbihbWUSUB2Bo1bQB6mZfUfRRxFhRkIILEDqel5Z4pVE0Ohti7gL9
SIek/ldWJ58tKP3U3lIeX+HHFNZtXfU/OTNIIoAt52c82BIeFr653uNlK/sg0Nhx
wBoBvgyU56asAVqdC6fmaqAh5T8wzNO9HHEi6YdZ8kj77b9mYewzxGBVSJMaM25J
70C4oy4NowU5uwtIc/UYJVCSpilF1VpkVmNQ/p6VYA/VCWQNzWOHCNDDelSccEaB
teGWyV6xrpe818YylhVXVSvyQ9gNsI3JPtdKUR0J0exy0j89seCQ6H/W+c9vHL9n
VzJzEepbd74SPJiEDFbfUygVuy1s3UC0IVKb/qP5QEAlIF39LcRd1i0HNZvq86Z1
K068MloHZgptvjWLns+QDBzV4h+9ot1Yo3cMb8FrcKsKaykeufYFtzr8mVuGZwKS
oM2rJrbvfYH91/fnTWU/SiGOxzCgHSOAJfe+cIoHNH+Bw/4EGEOU14t3stY2TPXz
o5REv0tmqGSYioacaJgjXWdzGrmk9LYFq4Y5bmPDHjGU2ypuvgjKc48R4xW+Ur10
pc2p1zBZX+dkDXvjBjt8hZBxtkAPOxqIqkmpVNe3BROFGXoNPspBfJUCE50oOwsJ
z8iyTy/YjPNzKXeLexsC/sXWjNTZdTjIfb7+OHYM08u5eerL+W+5/MHxo3T9xH77
WBbrAo1GhdJcG0ZwAOaR+suiuZRxLLw69svy+PZ8fiItlHFW5baanw+1oqsoYSHC
ToXDMaj+CGKhWtWUSkeHg0+qDWVoxrRCiKo0Ps6zHw7GNj2ugXsZh81yM6hf5JzR
xpPwma4PzT4CrbuqpgrswX6W4dduV3ugKjd9HrfUWxQfZI22l7dNe8GpteQPqfMZ
ZE08m2Yy4fr3bzrqFsiZVJ9m28yNwJ71r+UFJ7NHVxZBHDvBEeUljBxcnSzJuSDr
XZoe7/B8ytW3pgznGqqmjmZHaT9YWfuNqsGb7XQx5xo/iZ7sDIFivO0n7CLX9x/U
OMvIy5jVIgdtirds7R++zCL6QPRLtkV3vUIlZ6xiT6bpL3qaSDb3NoJg06FSGT64
TjVv4qdegbJ6MO3fBwqxT3/gMQ56X9JheeVCA88tKh1Pn0jPLUAszdxh6p8MIpfP
QZIvRN05nZPOyCxyCTUnOGrR5/P5eYollYjv96deCgwQVzghskbore60qX7tU3Hn
qCiLfN+c/Ct9ibL3LATaijWvEJUTYciIfp0+gNcGqUAvnFb793QPH9tsI1f/CJlP
Xwq2Cv1PkaHDNCgXir4SdlHpWHf9DUbeVw6DtkATvIcW7oF3/bZafNE/Zlq3W8BU
2iGTUxSp6n+F2cGnQ1TkqzwXjC7x5isf4d/MlKwuZaTQ7oqG0N+Ye5wvEmLASNCZ
+oj4QrQVmI6gu/DFX3UZ9Cf8aq0JGIvk2YlIi4px+rH6GITal5VzW5TqmY3RoICr
ZteEZBEY+YOrYTNFVA5VPp+PgGw/dxOPejz1TwxBDdO/w91VjGr7n2InEGy/AqSj
YI242Y/h9tBNyqgU97Y91POh1Tu76wg/8NYWAtBjzqkKy1SDhH/LuhxwOjefKYtQ
poYCoyvwjF1AaM+h/5DDT0QbYd8L518oBrXfvhPm39CZSLaRd6inMGBnwV84pFdY
tiyKyzQ+GidR1woJROXZf1gZzkPSzfvyY2VpQmsti+uBgIhUKcUF+fdRosfD+l7+
dlXoY8h0YYzs7CMUseE7F9W2dPjIBe87gSxUnrApEMsZZy4DxgMeJTZUwbvdBKZb
/XfxcHSFjsQBXasjSfmMUUCu+XcvEzExajuMPumaQIWaT8PNE3t6mEoXVgQqisSd
NebF6Mgn5e9+f/CulNdKGNUvge4eeClwGSvxEqEvMwPNfCgPsDhyFqTZ39wMR12b
3Oe7ldblIqsg8Mivwz00KLyO2bvmsxx4CifWcRCEOBLWTh4twJZdL8V+edK+2zum
SaVjyseJe3wlfFeIRnnFq8PKCEI0CV8dq+UGoCKGTI7TWM8QpsvB++JglSOMR0Ot
NocczUuFRq9An0ZmqGqDispn1iKEeR0AGqv6DjLSkyq5ldvZc0quHxpAwtL9Gecd
qK/peiuHQcGso5D4+78Xz8hJuMTqbVJw0pmK8dTT1WMTjga+yoxSSkLoXCPuj5tO
ymr1KTQ5syyMQqSy2PuMcMBmByGGJO2b/0ViKA8CVbMtBIg7kFlD9PdJw4pj7PKi
j8+eJXgWmvG7MZYoXa/m2ksNfUjUeXNKY0zjIzmx1+v3V8Hyr7SiZlwOF6LAIzfW
57ycbE++hDaoahz5YuHZN/kufZERh8V0rjiymu3zXYAPpT48BrQbbveGN9WRF1J+
CSmq9VJ4TtAsct/b/qErCFuOx2VO2wsSImP0NPH86hqaAniuCPJjTzOTnO7x8uFZ
lMXR9eIpTVX5hvcAHkmu7O7pslfqCUceztCUkureKovDDewljdHhov2u5DFVKK3O
MJOxgVYU8HgVC2CnI0xAXihWED2eqUCm6WYLyrQWg3oumpeCNY9Z933jZuQQqO/d
Pqzv/qEEsfhteyGVALiZ2Zw7s8u5cl+9NSk+CAiDR84ymySkuevYWS6U2qEJrTMo
1p8BFVmfMIJcmTBaxdct7rwq7E7EfqE5mqekXWq4uprDdqPYJEJFElO7aOcbVL85
XuMlOckeh+JDE5nzMBuCGTjI7Xc9xUTRVfEFKRpz58S3VKVTtjriathIT+hgVd7W
nMc45T23JPB/8K7SXwRXwgVvET9KTB2rSV5vsbateTf83KTPUZXxrtw++yDSixTi
7HQq+6rrUXKcnm0MX01El8Cksejf0HuziOYy8utMnSv89112L9e9e+5G6opwE+2s
cLpYTrhWfpmyER/VIc4W6OvXOPRvQTl0x/EKw1+xuOAj4vGnFp9xP/1B8/6XoBza
eftdict9uQCVFcSbyNLfr/2uiVZBDyUL5iIUeGt0vWaXHIgVou+iOWskMKGwI5+C
e6JFbDHX7nTAs2yk/KD0gzOkk+gDKWGfU3YepNtP+YWMW44v/n0OKx5MBdn7l5iF
/xpXmdTf1KXiEurzxYP9CC5WNtWQPHbo4DFZzn0ZiwNGqdnXVXXZyKMgU5w9ICFw
EdWY86aC+G0C5uiwsKrKYJ0ea+fofHmUWaYXTdK5Q/qDTEy/wleATQsXV1Wcpsuh
B/PPM+VBecTpiTRDTCpicyMa2+Iw7xedNGRftm3iFTvusfl9anovC50AcukxmYG7
HMpV0vLKKgjQ5+zpnM3qEaEZ0FTmLNBph1AMGGtH9TQbN6i5NlehSZKAzn9S8C+P
lE3UAG+l+HyEaGVXA18aoDH32GTBaaxMItK/P1rK7LuHZb5HxjISFfn2UhX3QBSD
bjPGpcihs9dC8QKDhHl2gwVSpzSqx2UAH3dfqO4iK915Ji333uMQoCXEtbSAoVyo
e1Un3FiGvgfz24cZWsYwlbLX0XADuAwpn8wSwzrql5CmT+LKz7BveK7N9djLn6k8
HE1j58ZZFHCNQBs6k7y8+QOhqehY9HgZaLTJSZTh4oktg8BmizDoNiCRXkyOXlzp
pKbM5poSaqJI0q8zBWgwqbIwZwO2qaLq5vt7B+0w3abHJzNW8qkOusIlaqqze9b0
JHgJ5jyX7d3IlH0ewb+FSG9QQiflroAqi+6hd+E0O1xV9ExFE/q5YEVluhhB0SYp
axSUbCYnSk7mOuDNppdlro5L08hdZMF9ZCEhW8bpfpS/tnkPyYE0fBxCMXRyi4q0
KWq4ZcQUq4CsWpc5jmN6xppMD2iO/JtmyvwqeeYA1fnbXbuPJWiyCH4ZBZARVI1f
MYNhHgISzJys6+Wc749QwYLYpsa1LFUD7BnwJNoUXHKQgHa/85UrqxsuDBwoFsqk
t2KSREvguhXSmEEKp37YqifhuhGAzvIZ1TaMXfuycIt1XDQMgSPT0kO+SG2FG7U2
+/goQwGXdPDWc5dWNQ+vFWrWrgwnLej7+ou/uABXohTfbhT60w9mpmY1Bo94wzWx
zVLnbW4nGddvg3DQ+4kp83hphGPH4riY2MLrtcbid7dzYgvBoFriauVCGg6mICKh
ar3PfH81sNg2hb5u+a6nLTm8TXqF6V8zfMUkYCwM5x9j5xooOVfI2UXQ6nyDlnnp
veHNHrOM4AqE7toQcsjrxAT8jyhiR+Y6NcXbCjKRelJC56Jc1A/tW46gZBcESBHK
id9BhcREJQOcKCpYkTLmXOHU8abf5itgkStUoIpxgk609JTJuHbLfM/1syZcxFEl
OUQLv0/pnaY0Jhb898OeO3qlO09AxV6LlCX/OWNxK3Zi/Hl3FjZay1S+QQr+RkO2
/69AXqZWdkGgN0cBesrk6InAYSwok78PcZPBE+GFKI2sOFYceNfMGqIDEt6YBKEb
ldv8bx0c4auN4HFw+wcInSdTkuEH4dXQHQxXcJceUWeNNvkcHj9W3kShx758U3BD
JFxrFLMySWxxPusLaPa6Jc8HyHAWv+CP4XIhOk9Z65f7o4si/q9ZVBMUwRhIte6o
c1uL61dVUrXIJlcJOZomRByK/ohd73Q/5rFqQCWuL+shCk0nqMZeMGpJZz+l4cHx
+Y8XbUKBMImX4ErEFzA9A3kiD8oOHq/yhb6b2PRTRbFAaN3nG/F0+7/YJOw5pHD8
GWyrLnipz8YpoMMu3ls82b3qYM45tboEL6vWYLxB5U9L63Nn3iM375QcQ8T6RsBP
Koez2RznEtPSDe81c7zaTFIubB5aKRKjBnKFn4tupPwTTiLw/d7Bk38AHCya3TeJ
hrx9jLMEseeDlorJ4henk1xz3BLoj44Qb1UJKY98AvSw2m0shfHkPDQUoICCeWLk
2r6WKleTngEYLHtcuuz/ZuFXzR3bGga+neKEBrKEo3ZP5ub43L9n5E6kyyFmGMxr
VwnovhK5AM9gl70YcA9f3KG/Wic/4s39+u/vJRdD/CMs2JAQkEa1nwLMK13gss3E
9Eh0Zs/cyhnvNaBDhoTRw3/x2s4JdhulKSznxbLS1fWt+aDdCrr4HeBqIs8IpqxC
ThYxC/Y+/cPzRiFOPjJaLVLIlT78+r4d3idQiNCjbBBIQNM7JiqaD+fCH/8nSnhE
AwAm5v7IuTzSosQkHOh5N++nbYOSQHhxIEqySva2JNFWOQVFb6nnWp04aA/bRmAl
mVgRsSLY3DWoOTwskgrG7m4jxGGlsngX1b5Lyrbr+ocvEdx6FITFS2nskUmghvFT
cZ+v6ADfHP4TaCcEnpKWbpXbYl78esKiovl0QrxIOrgdx6QEe/VPYebBmFlwQbFu
AlY7FNcXWOEqCUIV6hYge1Zx5O6K8cKTxPKpYFuK657ikoufbLLKNhRNi2X9OnmK
1IszeRM76V4P1krLQKOJNIRoG09v3L5zFqQp8iOaMvNQb+quULYKeC/1q/N1rl9D
yl4noHAysfkRRFH8nuF2AMyZvjfRjukVH24JI/8syju5kW+zN+RWlwrqva11ORiZ
A1wdOzeQXCfdp8f92exmp69Cd3/V98dpW6LKgNWAzZETO7u2LBBckAk5lJfWJHk9
H0evGbJ7Dbg6r7Fom76R1FKRFNHuWdvJoaNoEt5ILEdkyKe/YsMEjPHrL/IUbnpY
AMV4KQ8sA8K8A2zzkHqIx/pVrNBrJ5U7/GxOyqR5g/Ie4LUEHzrHlasw0GBtYXJW
W8Ems51LO/J5btpYVhpIb93iFPMPuL6c9BhivsHk44pi5xK36GGrxP72SEZbvWPX
NOYkmDPeMhsWcnGbrhVwT0OJwcCEZ8w8m4FbYNeVkRh0LYtRx21Lm5uIXQgqy26I
7sApfGX4/GPb3ZsAvs/PPX6QAF04ZJxboIf/Q3MGW4Fulwy1DqvdVKsI/uhPc77G
7XHDaW5XnVFcU8St7+pQiZkzfMmxNkujGy14uF3crzvXpB28IDTzuK2eMSq0tlmT
Uf44bOr2pvEVZf59UccgHv31IHq64Oe68PpeZJOUahE783gAWj4Olrym74DO2R/k
Ox20KPgox8LfKMZ7nQQiC1onF7/k7b8PFRhvHxK9hQJTQP7FqU6bZFhta+SOuu3G
jOM2DrmKDubf5sznYPHHatUGIW0MzUSD+xfHUX/44NRhx3Up/KCYWAFzhSaTxr6A
5O94NrWFJd30XEXMxd1jPebYUVXFA/SArYB/F76c/GMR5Dnf5WorTcTxn9+S/b8y
G2V4CSPtAVTWTC6qJJbOA6TTLobusE0LUyuAXiHnbqH0OW7wDhvM3U9qhojOlql8
vnP+8zUR+SoXtQCbRa+iuzCkdkF1WZJ7KF92Y1qqu2CN8ueuI1zCWRfLfP1WPYUO
jwLTtyvQ2QE8vI76fBLFfEDHK4LeeZJn+aCL+kiny20nhXAvoMvHqk7TP7X8qhFH
+3gUHfMJ6DZ38+Nvv0MB5HO3RBxz0dsxmcgJGnf+nk+jb6hP34TLivOW9Lz2lvNo
/VyU5duLgLPC4MCqRFPUTvkmJZHMWo5Z6bAPv8lWpPQR6rsUuahBv9zet4h1FhkG
xFvcGqF1zYufZHdfYoaAcDArSQxpooJ9LuLN/y4qA/DsSiChSQwWuaxTV5bNfUKq
0tcpLBNLUS+Hk22pbTTEyygOaOvSKamKxkRYDA5OToHdTu0n41uX1hf2YH0/D4ex
HG1zsWMJqgzm2SZ/QpOHaZxsf6ilClPMEgbxhrV3tpBTz76v74NUaLb/76oCqgn3
BU+Qg6+X+vnfQk53x/CxtAzPIks5JKG+k1P5yLOCEq1FI8+AJxZ6UmnKoYm4ETMJ
yN4HxpjVUBNJDQ9sGiNCgrfownWJUF42rugKc5QwDxmpui/wZRgewXaaeZXgd86H
8/k6c8xAGbQttwagjU1+stZLq0pomIlnxyD8bDfuLQlGN6vQV3OsleR5UPnI8SOI
YzlIMo4WqnRC+8n9v81QBSglcZ3xsJ2QpxjYxxRhxYSJyx8dKywzWzNCA+GPlSLr
2fpm6ReZgBdt7oyNfVjIeG1RJ1tKq703ikxKW8QlFEQyt2YlBkfdiICoY74N7AGd
WAjk5MQa4B++CKeU1sFDvwd00VrPjPvLDbH5DtjoAfEopnNo3UdvsUSqfel4Zw9f
eOUUsVaYbm5GCzb15lz6gmwwi4MrCgtcnAj3S5/l/FD8qtDduXOISdjNwMAPGTIN
PAUEwSuaoEv6K4bKQQcZSGafPU560PJ/1iI2BU8g29mk3SNXQo88zKHxSEtOQ50v
+SlOxf5MGFRfpAtSV916L0xbYe8rc6NsC1qUBl8+v9TSCACtTLABO8Y6VZBMU9N7
ixZvFS8dS0JJ7aU1aQ1e4bXa6rEVUFEHwhBzZjnQniH6yzH+HiefLEsSfmBqZtb6
zjDAvcAfvxTQqnhZdZEXKP758vWxtAvq6lXYjDM8tU0kVLkj6iET06G/Eog82TJ5
galeVmORGMcFuNCq7PS/kvZEFgdq0xcMoOMHVMfyhU+2MV3a/0CQjHz89n1t83JW
eTkI+d6Ohm+EH68LFxz4GQvm0WJgJgN0T/5ttS9mMtcvo+fHwCeaV4Cp73l28Dx2
pqQ6iBGKLtB62UBQ5ItA6nin71UcJDhBQT+IdiV3gzks/sEtiTrrY3DvPW7aSA4X
vYtR4vfrqw0jCHF8NWQ85ussuM/jES1XIrQbHmEGlrpW6YlGB2DdUa4qXrVq6tAF
7+06p+Msi/WnCV2LVfkMXxEpp91F5jSgzAHnpuXOuhyRHuxr6qWSHawDfUZ/uQeo
Q7P4pdDZ0Mu9SLNml1EAfFEVYLH5MjC5GkR1oMEZN8shTB8sQ9qjFKx7DHOuRXIc
tDc6YfDQmzM+CozuAnezNgVIuHrsmZo3aqhxE7z12wLi74asZG0K2F2ZI908m0wn
3BQGkOQg6b+3cj0pKl1lR+wTSlegL+2ClW2VLlpJlnLegB5/ZQmeQAxjTAqSMqCG
P9uKh1B0kXo8VClxQQGI0Ez00IpB1w3Fsx6fUcoulRwjJygrLiNhB6+nn2OYdWn8
yElNKM+e/y8Yvqu7xSIUTpAqwcGxWB2FGNZOhnv4My/EqVFQN4xHdL93aWzvh0k8
7FcJwUy3a/JYb3RmZ0/8fO59JPlIEtEfuYHua0DY2jSezd7nM4ap1P3vWnCi/n34
xSe28mMpYUSyPS1JMqZv6Yb5mruDytDYdmJ2FSWkQW09mBKvquTrlGy1uTuF8u3S
CFa8fQLnLsi8W9L5e75icQULbc16RrdzI0NdvGlZwELNebMZGFbitofHv2rhxkXo
88zb99n8NBVGk7IE74iinUqr1qukJSUMlxQ/HEqfwP1giryA0FJVUoXMlmN3Z5M4
HKYegb1WigTLnb7S/6+dyHzs7TJEGyxII6ThTRPskYM4THxr1zeS79d7kRnuDNAe
Sb9XtCmkeU1a1xOgv5QTwx//IJ71iP2PS4NwHtyAgO2f3soZHbIRYtsjwnNi6JrH
Etr7HwvXBhneoYqUF/RcNiaa0xDFZqCHupCQ2ktl4uPikJ2Te0Oag8JMDzM/d5Mr
pGbvAvKh6j9vZoHNn6LcNdRJmUUXcIYGQwKBM1UICxTB9dQvGs/CCzrxjX4xs3QH
lnHp5/ePBqDtlfuViqh+mBV8EN44y4R7x8BTFpzMxqs5MRPcpZmJyxDQu/5G+M9D
iE+sh0UspajUrO2F0WGB7wDEqdTDVZ70zWJjBW06KT6h7rqV8YXxixL6SjEjxMqc
q0/j5XbMYQhYtBZQBgkNJNAXyxkXqrlo7nexJweoOj9yhs11YbYloVBUNDF7d1uH
/o1GKpr/JKdEGdiSE5+FFIS7AetNyZ8Kmtvag4WhsUEydUlqdzqyI4Tv5MIv/O4r
AKtH+QagXQiq2F5qxl0VrT7gz44Jftb5VDLyF5AHsUb+3Rav8zYS1plM/QkCakvi
E4sJRaxg5JkauV1nqXe/5GGCH0jd3cnyrNywj02GGpPyu63pMWGO1rPzgwHxyvX9
JkUmnTLBpNBKcJ5zw9MhI8AxtCi58S2xpvYdzL64ZeIPAYfLyvDo1IbVt/6ySFro
vpBaihPxHbEWxsBvNeATCBVn2kv4eXgZ5StKQFTxGspDGQRl5KPyUK53h8JYwkAL
/vpkn8FFHhSFG2Jyoo8cm3mCqGNq8CbXa/EVR1T4DzY0zWokBHl7Qz2pADi/hPBq
rC7gtJQ8mghSwiX3YCTuj0He0d2rcrtOqElxhzxdUjQ1f0iK6bQ+t3Ob+nk9ssES
05k8EXFcRZVLxY/FC4m3J1tFh66vZukYpZ1JnyWpPFoI+1gv857XPwjMiJwVnkeO
PM+kUv/YB877IyjpTDpDqFLU5aBimzcaoLsweCOfh76xhGKvxkjLdT4YV4MnOkVJ
jWqrTE84j70fI0ROpNEMsBX9bLH8FbQJCQ2adoTvJuFyTkjuVbfxcorPmcv0nDyW
E8kvEwO00UmnkNhpAiSqc9avhMZcEGH1OJPnS4d/l48veDo33zKd4BM9dUk7ySa3
sWwDca7DYFdeVr5mts81g/K5ReMz/IjyGcPbvwVAYLUzmPAAuADmw+oEkef4HLJd
iroQnoA0HGsMifvBABHm9f4vr7muYiMrWJAZ1Q648bv0E75zlDBU6HdummSyyFKf
eA6Ab54rZPy1VdU8v5E1at9+XjYx00mDMClwFxjgcHcyZ8LoZdIirYWEFVP6iy1Y
x3mafQ5F6CjDez7DJDgVDYkfjI4+y7EjG5tD0YvdmMnrihTbR3+2PzpS98iI6Hrd
TBteEEYXj1/dI+elmDqsLhkBkfIXlv4yt0UTUVsxAljADLvJr5Tr9y1cn6rxnYJR
8RmFry51S5byKRuZ0iO+EKb4AmBT658rL5kiyRTBnnI3iqzuftSgd3MOGknVcogy
Yzm7LZRbl6QEdn6VJ4G2zr67cxH16lpgheSDz5Irbcf/NtIPUsm1/RPBbLZQIvH7
0UTkGciK5jLrGXO4UnPYxCUVLw5Ztmp+TWyyIt4Ehn6jeFmn0A3qjF7O3qVIxbaj
X6TOJkPmXkHVXrbvtbleazN5mnIhgS9q6Ig7xGc0rATxDUZwDmoDv1S72kSw4dkB
szRBeS6MF2Xy8EM3/OiJVXXjHC6g0MBRk1VpHQ0XugvYuZ6ENhimE2wv+vaD34aH
8PiDeqD3tnqQsINLy0YGSr70bGP8iTx54YfrnsRVxzg430RLkL/1RKNmCxBj+dBg
JJLWFycMhgKzDoLYGpIziWvWdeMLRBcfTjUpfCI5nPlxRX1yLb9BcVmbpDc5uRdB
cFoKYU0PeZ3Oopzu8/F2U0dHW26U9r/YetrQK9HkCluKHJ3zkb8zaN7tcrAqeTa/
jGZeXnZtCtsgYd9lp9Zpp+ZoKiPxbkwrtRXsZUEmMDyt0ygF63mmYQLvxVPfUOkH
JJDAeguAgUYV0jaNzNStUerzLryoh+2RTGu5agM8sN1dmKyMoyYpVSughY7j4b6C
tCKfjU90Ac59z8+MySXeBUE/18SjPSWjTpU2cmseWDU8XxZ+F9x0T9TM4Ns0ALZu
UiYNtu4tjEnkBBV+a8lDyIoOpMnOFstrgezId7eXpEscBW6tIE6sLN8PeXisxfDg
GgWDlFZTZFjmqNM5rfdch+7mKz7mHLIbeU0Bf2tGaxV4c81iso5wdPd8ndeEv7w0
INeDrv6ZPrWNGuzPLw+UJMhR/XUT0Yo7OZKyGOW6p8J6dFyJmaucesA+RQx4W0Ep
hD5JolLZSH5MDpIzMkyOO6xcUWnLqadMkHCwY7IsZVYb4XQpAI99AoGsXkNuHp0+
D24X+YzH2dkji+Gc59YDzsfo+Km3YgSzeUn+sUB9ZtuhjtKciuKjLsiEh/JrkYql
+etjTiuYwYjKODQFDFng66J5nzo5VIWrhODY0EX3WXWumad1zIWL7XSvY3035mSJ
6pfxBB6zJIlYAgB1+w8pZQ/9gvCw2KOwkVZu4Th9zAZWB2+OVL9jCIVH7Zc1w4NC
vIQ6a533vv6gu7iyxGoaJdcLR4mBsbP1fJ+1sEsSvrnz5gf32ninwzyTZ4hCccZP
Te6rVGyK0EaDYX4uhzfDV9zKhqCLBcVHX6ZsrPFXhzxNPzFKwEXg9ioCdelGgB79
KfGXgAl8+SsOCvvPGOaHM+6wfPsmJiBLiOyJ5iSh4UK9jMlXDzjDv9QMxgcrpiyZ
cyADazhxpj6V7KAobwT3lzeO3flR+HYV0yIOoij8b4nakve4z0zNIfqRyMX3i+6A
3/3yaa0LtOfftLW6vHSW/K5SsZW3zTfFwEi2pY3FaDVxAbzQ07orqpKt16QLhV2a
J6cDdMRo+v4RKWI+gmoQBZoOoxWTo6HyHh69Rv67EBCGnXlF8kMU5jDiZhgah+8B
tcnFdHbcTxR9GiAiUgidZizjxeWD+xcREwThXo9mVEMuyzsBp20bxreEgQffz/ja
r2yI0IWQ3nt285/eSmy8WasYTkrPwSRvwzRnjBwQswhSQtakYyOOI2ZYlBnvDRWa
jre2Jc4gsWp847sDTUhDEyP1MExsUzOsCPG+NCY6sjcyAR8d26y1UF8mCnGgnks3
FGTYG3CH3kh3QnaeapPRfUEkrP2xdu7sDqiDawrQ3qCC7Fn/RfFIImOPMZZcbe2T
h6JYS+O8jHWWPYxMt0zHV4u9ihd4e+4Ok/UVhx7L1bzKxDI281FPvUV28w0m8+cc
MXLSdppPmIkkiJg46SkFHKzz3Co/ilWlbE6RtsypdZJAAuGjTaIhEfMJbWe4WYIE
aN1XRdZwZxmhY8S+4j3vcbBigLuisbLAg+ZchbE3MNvUcRcsZhEU0wMUjXuUx5gb
WZ9zFVa8OjDWoO2GOHcCWwiALsYhrpsV8RWsfIhkfmZ9FRBZ+aRsjcyMfurl8O+2
1cs/PY+rD+M1yNtnEZudOU9iueHTuWLA2EBC2nuYZuqPlaApmiy+xa4406vgd8/i
YZT9iEbqrs2HzlFqzlxPeRNm9wRh4ypcU2T7yhbskBqvzbZQD22eb0Oi3/UmbzT9
J1jKQfnIZmnfuCqqiGuWaKhOWGYLaH5eQN4cQ/88It8Uh+XJk+JGWq8VdJj6P6ym
KXUJ4Fx+uiQlTVm2AwjpgTz6u9FR4mNAqfM4qPNCirSOmLGKrOGwIN9nk/9L4jUt
dMC7PkexkrWu1JAUUcGZs06dqNe/m/PwUP/+wZwVuSH31tYuhToJl5UCJCV8T3Q5
al5L7Ig58U07uQdXFKQG/kJkhXHyv5gV3/AoQbhdDst+vYTmX6UMkV1thhXBJ6Gn
eIQkTxNi5vjfZ+r082N0jmKBjukzYD8lw9+yHuA8hez2xiI2VvEGbMLUsjTWJ5BQ
6ZiD1cqO4ZJRIlEAS6eMg7KeM0mP0ZJb49cun2BJKs6runlgiOLNVGpd4UNjegT5
tNxEPHEmQUjGBq3fLdDKi0b+CpD9rgu0VhP3Bhr11WaN6Em+EQL2zrzFFIASuNwF
0aFeDUkjoz1/cviQIwnFVTB8U0l3tcmbS6ArCpPDJRt8EYXQkCgH9aPO6Tq18bmd
fRq306zimWc5bWq4IfOvIMhFj6fOUD0FuuccO8nQx3ousrtjt6Esmget8skfxzgq
JV4iq+1v7rGi6xlgS3eZIgmK+jDqbY3MSpkO1eUxDA1+qUTXvcwzdkNRTNZr9oFN
KutfmsDqDRJduj6fAMTrV6fle0+IpMsjeisj0SSCfrH2kxhUWkHmaJXu7QDdwVvv
9QweTAVIYXUGkAsS8c5w2oaTlIwp8ZUqjRz0fSenjtApE6MNDt4PRZn4MxWij/D7
2uPJE+Ng1qrjNn/iGjwzjRTOhYuDzH/dnH60EwBGOtzHLyxkJtxb2PA6+5caHjB9
DnTfxO/oBi2PcHj9ciHubxsmQLgKbizT7Bl+E6oKiHb3ncd5lxqT06WjjBAX9ltU
TE0i+ggvCY1ULyms4KiLr6bligCDmOLYv45AcX54IY3RiicWEty8TDr2VQB962H6
Gv9BeEQ7ZsnmlAi0JAkIabvgNJfPdOTsfuIFfzFviARzDJ1F7VrWefQ+mram7sdD
wj9MWeupcnL/2y6ZkIAxBjFvJHzhNep4M6PjfmwymhE7+tOqjUXrUUi1y5ARvp5q
8bc6gc+ludiKiOx65ekxPW+C9lCWvPb+KnCVtsvWy5CNOYACwrKzQzWOV/9tNsfq
Apeb5drud09rEDupTcRjq8Dj6mCqD9PHFPVK9TemAr+TU158VTorWF8fKnS68fvb
4iENfpPIZkMYe1o05Ii1couRsjeVzg3+opjyLuy5V3S1qx9vm+IXqAOq9mnmCtvs
i858N+O3kcngi8tehtunMPZNIZpcKzCWgY1nSA/AVzcZq1ADeWCm9F/GiKgKuluM
Qog3LkfK58J25EDqfy1f9n9X3TK8HlBkRNgiMgUwAihR4IrrFUtGrFYBm43f8iYy
Zb9TPWI9QNJ32cgXUUr72wZwS+ulz9PQIm/dZ2rhSG/B+BoPrIAP+0pwl1TI0Bld
MTFTasXaRdgmE9l+89DhwLSAcg8tbUt/6miy/RGhnkEzsOFyi/d+iOZKfogALPcq
aG3NDN7kaYHNJIIfjdInJZbf+MTpnKlsB4oYhflBp0eoikl0Go8zKtuztlVM+cjo
jJ2OJPTnKnSZawBSGd7P8Q8EwZF3t3BY/xE0HEs8+XdLGIvL9AxQH6OCY3pzVEws
c8dNR1ZB8dHHval4m6/pDOGJFTS9x0TM3QXaJwPKD1V01ND7YFQCeQIs226hmFyA
sT59dJ5TurT9c4dAJRhsIQAn6sdS9+6Xifm+qQf3O+RvpGDVVGmbhKKq0xxYcsoo
0jO5BiB6aRe1KPOl5AsnPZhN6CNqBSnn6Ho7cL4NmYYaIT6wouYWhXE+HEh2k5Jx
S7w0aECihaDBweYzuKqBJyYpHkA96p8EWIvOrQtB2xR6HRlYnc//qDtjS3/y8ILs
fLPzU9ZjDIGdZhO9L6ZuMlDl1xRWiPF5A+5wh61p9Ryqfm7Wpt6smJw2aQTTEti7
zhc06QvBRUGQEvi3ALxuBe3OYUsCzoKa0ZJuKxD755hTd1d8XQOruU6kS00XvVAe
QQBnigp14e5UvQTgY1yqWlQuVydPsSjMhG4MLduyJrAVxMxV/p8+fnNKu9A0QZY5
8RBpravBe9h3o5V3n3LT83ME/+sln4W1eTHXDT2R2fUr8JVDt17lXfD0JEh7zbcx
kyY9Z0/svOrrAtkLFMpU0jLkNzS7hnSDzZIeJc9YoiJwWp7fffuwKdhnpH+mC0aT
MXG3Pmmd1+Da+y+CijK2RuPO8SlSQ1nMVeFi+UgawZEJ7zjt7HdFBUCXm0eEfzVc
XY5HW4hLqbkPgW4/4gmkwP4vtUqvdeCZ3AODN3I4NcFQAn9vpIkay5EUHYbq3zfz
oLsxNkTh8Si26d7xuo/xn9zp17UcdBvxgg1DxpfE9FTiFQSJKUWKXe+Do5Q1wvau
tmvE+36sf/3doR064d5nolRu+cSiwZQgDFbWzjZgd79GGHYBgH361Gyl5npwCxQe
0PJF7ePYqJuTuzswsM+oUJA/Q3er6D62RX5E8/aqJiLniSVYaOGJyNpdDdkcoNEK
02NpG3493H/5XdnrAOafPoBOEWj1WpUXz15WKNuaYvA6Q0/WPPNsgpXuVD7IGO6V
L7Jhg60q6dqW5I5q5HhuWk5KpY1Llos2w2t6Dzw9Mn1phX4YOxGoNdC8qzP993c2
uRzz/+MBVqdEcD9ebh0BoVLT00o52T121P52od76yf1cCsK/yfw2wm4BiohVBiPx
b1IBdFg/gTXBKtdQ5TVkt5T7MY3iSM12d8eIl6mi85P+Di2x4/fVIHsswr6GIWkY
fn/FfV/PPTldPtJnkRPxctf9VsgJyDeQBer2oErYUJwrRrpva7fux8ktuWcCGIut
clwgMXumvt1kUkZYxANuOj0M/yci6Q3sHoVzxDVoYyCJrNTQARrKKqNVpSkVip+h
xaN5jwx7vvTsGcRNV8vMeOTgQY00BjeTjaaqaUkesaSarZi9IOejeKmH+BUSvMlk
vvdOHrK27WNOru1YgPrBfEECkv0A8dAyigcGRAyOj6A1hiXkI5hg4BS2ETr3yoq6
RpK9iQxplPg/Dgre55s8LSvpLAACiCbdCsQiCFMNz9gcATxxwKtaXx/hpUotHyWu
rs0EJJMbme1RnHS1xe76giJDaP7pwYJrdKjXER5awmcRR6f6nFwz6pAYIxcaIIVa
KjF3S9CT19Q8Hmv3G188jrgV9Axf3cAou4cuDvgjMDd5pEQkip6t97qUePPsZz7a
vqf0caehHIZ1g54HHIBi5zZyv+eqveUadvu3p2fXfor83JWdHNVG269D1WxfMzNK
BO0tYk5LlgebsMZmq0r192P2/3h5JR3wap3naA1PO6qnnmezzEWw+x06szvIJ7z2
7he9jWCDf6mCOUtRGdaYI2IL8NHYPEl4hk0LNCUTMuEerxSyo0qpFV8ikjAGwVFk
dlaNq7cFaDXJ8PSCdxyu5XlXhN1zrhVsHa2PId+SyPCPUjGwuQ/QQ/RIHXS4yH5R
Q/G+X1Ma6W+43fFL8tUwkqGfLIKeSGQE0VmilkYiIminabCxDQeA2zdwgZnCMeEV
1gG6YR0CtIlaulz77ZUAdVoDpzQPWtaw3k5d8Fp6N479YwChguhWqy/dLRN8Herk
xA/n8i3LCHlNNSrNX/+BifSSjug+dWgVe8jRACVd5DtDWfWrf6Yi7JiOqLEL0fLZ
Tara2Q0AhCV0BS4O6+raBYCMuRrv9OlZKVKCGVOfdlitfdYby11VwtEHVbNIH2DU
S+mt1ZkqQ/bvNJGa+3yJO6BusDg8iImzrwUMpUfhTmwqs/fGXVM/OXxvcpVwudZi
Cam/H2Egpl6x+waL/GmAuVN/ISndg17RXZfpX9jtBgAk4AN4iJlwuKmjXVKzBa7P
i9nCR6uE8YvrqvORqnaG7/rHnA7/bFbsqahv00y8XdM2x2zUmoBfYoQmMGDUKk7l
ENs+KrRseKZGMyXazTuMZWr34bmbUGG2aTdSJYiz/nKsy3aUGMwgAcONgpx/mLhD
2nnlhJitQw/1PHYUlFSTwzpXXjkstXN0LOVZIGLrE19OXCm7TaH4REYkxb6zlyjG
n3dXi/t4rN/D9jfocXm9UUgOGi/7x3PFvVXURNtyu0tdecrKHXRt+e6qRbS5xcmq
udr0blfNESpzstJdAOCmT3mDXqMWks8IyLK0mtVw8/BDC9zq2YTW0w+sroRMdHpf
kibyW1eC+SAlVseLgcGnJWNmDdzQzWhrpjW95txshWyzdnnsjJ5Ubh8PeaV+AxC+
M32rNkhvHPbrd6rnwGyRVO5KxPmAowV+zh7EDXElw1cxavXvtm9XmLYG5kd+bZ1l
kzh/09Ebiz2KHw7exDMT/mE0ErOboJqgl3tdQ+cl5qNNGYVOwkkKi9Bg6obSJte+
DXshAAcm+cNtIO07dUJALS81ytTNFVPdUAeMRBFH16ah8MeCEeybbv0DYe7HO7Os
kL9NPYOh5dFPmsLIxFpNsxZcwnJvGIeRnnZSJTP2p8IskuianQvXVVwBgRwe/jry
MqBatszQzJAmx7ZrKaWgF91edCuRCJ0d7//dQ1y8g113K6HE5/HkdvmCnktcyVC+
IsyQqsIWZoMCeALRFVctJPb0OpArJuanVTyy/vVQv8GSFi4FFAnKVrT/V02Ekjn8
/lon8CAiWf97CmYZC6XojZZMzk4JLgOdDNGCVGn2lJkgHdaOlzHkB/sWtzvsXNhw
ft+4eh6fnwCEeJMy2uhXQXKxVDE2Kb6iR3ZajvxlMrtY4LvzaW2WPLr5DieKgvk2
+0PZj4lIVOMhqfFN2lsWszI5xN2rWStC4YnonKgz4gZr23qWgG1Xxg4ny3cga7gX
EnjESPcaIyOivDFO9tWKOjTaWBcnFDbV2byNgt/2pbvmi/2wWfDBGJGu136l4NT9
MbaPSjbdtVYQnKcuWAIHjZ/VaAZ4Aeoq3nKxuR28YHH1JSZHojEfIGunVfPnttvM
lsiKb4kuUvO4xxVHRxBtXSYbCHL5JPj1ZdAeE+UuPKYQ9uSf9fvWNhpQC3sDZSbD
OYyJKULSXUWKP1jKNrDD4wtn4DIJpJCiSXEBoaihu3YPDaW7PuSNkD8U7G0LbiL6
XHYIEGcI4Vpnxmrq+SqU1czyuQEObNpmqorFB1z98/XtsLPvO2SJmfIYAcL7c3jz
3J12I0pLDUHpP4MeVCQHJDk5iJnDIcvB45VsZCWqQY08d9cMR+Zu1wYXgpjSm+EW
PyO5fKIcA79JeuvAjXUL/n+gruzRid96Ok4FiP14mjoevAfruV6vpQW4uTaGtEhe
uUmsOH1r1r1N557ZS7EMMuvYGxWat9TlM6q8GmqzDv9+DUEu4jFKuKVaV58+DP4p
ZCGwAWvQayqf6R+qOZ4qF4SFJ6ovmeieAhKCDyFNzzCIW5veBRRcnMjOJ92IySly
nPR+m/sYHOHaDbFaC4E4I2NMjwslsDCkWkuVAdZQ3gOfFflOqZ7qPgizEgvc1RPZ
sS74CTNdfRYkNPv7UtrZKtq60alXVL+e1ZxpwcptrXKhGti5fLCBZO0mXbcBYg0w
M2N0PX5X6DWEMLkiHFCp0kizlZHFQMoOeySCKp7R6y2T00sGoSGXwTMMRA4d+HpG
QgdRl3CgLxihL6siFG9yfaumNeqG5ju6Q8Qh06t2WwFIKyOrcAP4AUoDbvky8Ksv
FZcvV/wJ50PXpxPBO6wdJPKle47jlYloo61DXbPd2F5GKUaZcCRn2wf3CgwpRLB3
symn5ZnX8IaZS4p1jFwBJgeexythAwGocD2lVRINnW/mRDUU4l1xHOi/xbkTgVZ6
j1Xli/U1YSWHtLLbZa31ai0HO47s1D6ICAN1bfo2rv5aDZsch0l8Pf6fHlNjNXIJ
ZjYAfkHaZlaQsPU0GvaciuTlwi5f86NhUfm+2BMgOsFUh5y1Pnprk1QI7YfDMI6B
/gLoaz3E0ZbKFqWfJ6JocW9NOxuT2l2YJILrBXHxqMW/maL1FBMk546z6a8/Ej0v
xjqZfv4Eek5WMxG5WRMIr2qaSAxazpCVeOVgWyj/ANPrqDzfhcqHJSDb2cwP8BxW
cL1fC7St3z9atc7evdA5JAtzymqLw3zicC4kZ/u5wEL4MwB3bmPI1t/LhGVheEK5
pOulmJCNRuGzXdCCeMUXtz8AbScbsQFMGnkY4mSTYtHY/gu45NkPMMOX2r/B5Vg8
iu0JgbMmpg0V1yq1Gr15nkmd5ek/MPoNpUBA91zBlUHqUeZ/rDhg7apCehTBM+k/
HqjnLdeJMsf4D0toB5qowZJc4YPVFl/eO74ud3vEmVXYpdpA1AI59Kqf6mSsVU/u
ffc4VQ/Slbg/8TvJb9VO2jRB5/sYjn55HwNZpvLu4M8JqGbQz8HrOt5SgT+re871
hNWfVJ5rrB+VZek0czpO3v0/56GH9lEHmxx7OyBbiCuvf0PiSZfQdpfoLotnibLN
UejY219tJFCAIIWhuCn3glUxMF53FKAnkpMSmPVcwMCisoGZ0AnsFLeMQ2zVZwp2
myWct/f5Q1dqLdW6KAB3PccTyUb7htBESWEImCIJHreSq7XxlbDVERRAHuAEdh/g
KOTI5d5QXZBfyyluQh+lIgWIr4ZtiuF5Hj2Nk4bblnqX7SlIPm3SfHheUaKSaVii
/9DV9F8tXOCcUam92DjKUoakcvx1iEJbWXmRJh22jaDlABzm4vbtVGR0iapveH9d
sh+WnMe5GWsfGqeH/52hEcaqjpaoRzEZqOiIJtrgy+6OM1TR88Jv//DTBAL1CE+h
rawYaGD1DVRrNB9Gg6dA9KmtBQUXZgRDpXyazYYC5AISJZCZC04FyxSIPuWpmEsE
87RzdAtGgoLR4rNbRfjUoi/4mbOwwi3Glq+sh4QpiPXTqJ3TNnF0WDzYPXaFX82O
YBcGhY5lyF4QjdEp/lLmHTx7WQMapP0NqLMUtPui2PBQZ1H1wC+cu9sWisaXGKMc
gzhIY8cPWU9NNU5VO42O+WJ/OoIKWL1E21ZrQinsI7bkccLd/c1GLYsWlUpgPb2b
vM5K6toXKGCCaYhCRhpOngf+Pwm0/fBRC/uIROFVbTFf3CVta0gaMRPd7/ugjfgS
J6K9eYqNl+h+bs2wdF60sHPqoIYJByJoO6cATY3yQ0x5tLWic0kPPISNme6xwsNx
J/i1M2VWTnu+ol7NQe04isCZ55eMSg20EIJ/KGIq9LqQy4iaGufAe54DlHBS2gLu
/4YDY6dv1SiWXuuC8UZXmehQEEL0h89gE2vbxA3W77uKqXgylhzKUf8ooQR88g3O
ryX7NCmLEG5xpOyaSFrnvzpTKUNcYMYl3ywLvNfdsP6MoqY3mSvWthCrqx4U273K
weVNrQ/XB3b9qAueQyql4cB1Vity5rblJXS3Tyq02C302u5PxFgDUjImMhMIA/vx
ds3DT9P8BoGJ0eJzx8YJJAgegSigIGn73dy027QHPU39Lms60JQNK/3rfg7kcAI4
TIacGCwzZ+b2sNGj5edrfNV+QUn5RTeiH4gz+E3R1Hyk+eae6z8fc25gY/cTNUv4
wmOh66zGiPIVAvsArXYY1xHc2aoayq0DIRcyEyCu7mWvcEozMQ3L5fmLs7viYiSg
niVy91LHgO1nxBZMPBK5ATRDXVJGflTwGZj0AHnZR/PzAXq12mq/4koDsqPshVBc
JV3ZXhdi9ZMwTWLx5Q/GphwYhxw8USeXHyQ78eFUoR36NxFY9Gdc+dJKv91NAndD
zxIUewsIzYeVD+YfdfcSl9SpRe3N6P2AUXNSr4IdH0V1I8nBz3uDncT4r0AwG6z+
BmYRD0JxfOzdsS7p91BtCY5tDKO6FAE5Efi8TSeK10qk+J9rigg+eDL4P2ZS1NnH
+iRekv1J3dCV+Ke1UhH6KH3B5OG/aFgpGF5FEIS3fgartywMo26KFU6MLwRV/mHA
BEKaW5FsFWD8gaSSBfKJ4i5pgYRsibmTrarGpQKck2BNvv7oR69UL2cWxtmDk4Qg
1bFgCARQmStIpYTI+KJKfgemxr0QLtK+c1C8mJAwG3fM0RAewcl7HhYb+4xWH6z1
UIde29MyMH2myL27TqUHXG7Bc7P73chb58sZvBUp3Ua8kTtq5Iy1F8DOHGiWSkCU
cHUqxMOuKc9dvXhUncqcgS877ns3nN4lNYrr6KKubrvP0q6EugIuS0xJBj2gCvf+
os60XDSQH8HTGklnSekEsIz4N8p4rVXCiw6b22zrUiAiOYQD0vg10KuFcjHe3qR8
K8QUpkQrr6fckLdOmDCnaGve2vxCPuCsQM06/Fa2k6Hb7RPdPgLzC8IdfKqLK5xB
cpR40xL6Gxbm7ALoRgQdHU31mj8dricvhzWS6GnuBqQzYUhQplgo1b5hCH5N2OO2
Z3BmUlJDfghQlkSNeH36HxsGyPbsbMPL1cezNB3ygF1qxodv3ckeOyEiUObDeZju
QXyBqUauTH5U72/hkkGdFZb87ZKfmTh9LtjZoEUlpclGiUJiCHpEU2jS2u5k6hgC
QAPANPNRYiJrhXeoYV13HIiJzycwYXqUoKAxACBcG5xqYS3ju9ANuNbhEcPtNRr+
70K6T9WuMdE5Kv35B2GsC12KkO8vpkDHKWGyQ8UKNG/LGTDHiJUO+XpVEb0dmPYA
rsmBPVYRN+wjUSo+Qy2AAHLgdUTQqRSPdn9mye3cnVy1UpAUsXHW8R4+qV6f6g1B
9Xl/3oGpeaevKgtzHMY21wPpnVexYBc+nZHcjTHfMxza8lMcMDhP51b1B08R6NTF
HXc6XmONHQAjnoZImMhX9zmsC7vzZPwyfXP16J7t1ENYzhm12DI7dlElP7UkSmm5
8bKJRXXBBqs1bnTfHInoC13PET+IkCAykuzlU3NYwi+aR/1Di7lx/BXZZWQcpl2P
iweI2PNeCtluKMab81zac4GBaZnj6Z/1cAnwqy6ckjRxr81PL4zTKt54Oj8uBXzn
q2GNOPJcKvxX2kEUKawKeAhAVdYOX0OT1bKewnaZT08EDthfA18fWcqvW1LEodyG
XT2DDWO8YvAt5tSHlAq1xi58N1GGXowSrQurgESHU6vS1fV8y6rfswmwglzd+goB
pS+eDjSNCk1CiNIXQqNqAVxHxaRILzfO6lUt84LuOzbVYDTGOaYsona/rvpasaq9
qTkBvrq+egBN6WPxGDAzsecGIBr5Dkia1zJqFaveoj14AWOOZa6LmVYlQA4DgPyK
M7mHKFDkb9X40Mm1J0bn0ryrz0l2WrBi5QVrsReAGhbmEY3kRh5nMJyx7oVx4D1L
CqTFifrVj3mnzfA+zKMEemJlkcgEMjfM5ebCPxc/YylbtT+clynrG6/Ed0zhDrvk
rsDOXXO0BmBGWzGyx551B8W4WS9cI8LjVx/KqZl2tmHAYrPktGU8DB9u5766xPrm
G4LAzIoFjUZiD8cs06FwRRnusiQwPdWvOP+aqhO5Bs2SZKti1RZh41tgpWbE59n9
rzd6gUd+q9CoVU0c+0rzZSyzM6VR05VMWE2naM57KncN7c4cYQGiuF2ouYHQsvGG
bdKfHy1SvX+pKLrsLQievR/VDW/Gbf+Q93GMz2KOmwhAitygUVLbY+mo+1nQ8t/v
HSp9JTDANBlBzaAtyomzv4C152Rn9u4WQ3pNWKh13RuSGRxp3cOhNAF+lFoJiPnA
sZQBiI8+RY7DpBEivsUd/4Y3WK3paEWcNQdWZd+WmVzutQUxc76AkvUnSlXfRf53
xcdH9AChXCL7c071IVQSwCC05L1BSlNuJAWytgrqjNMCi+l+DybtyyZelOV1/IHa
YfFqE7c5oorCDRrInBKK0K/Ikbo5MKnORUTnE9jWzYn0WvN6GBMVOD8NACdGU4CR
ppgByzy4uc9wVNTYrztgq0qrbP8zqcWu7LeQ8XiFS50pQPbfaWNbjkw+M9MoBWGa
J3JsKYonDZgp4pe7rNfK+kL+fx7ww3LLS+ZEMUxT6jK0SdJ6K/0Ef8yIdIIF5iDP
p9g1PdZz+hqYI5K+llHmnoZyJEiDyKlD8IIKYSQag0p4cug9ZaB2FQ2sXQ+dM1DE
XqwsWneQxrwz90nT8VVgXFmyKayjKteV9R3Kx9/0F0llypXl0x+0diiR2Gr7jXi7
iWDAFQOlx/qA5kSoDuI5CVXVv72CPkjOtKwaKnWyOk5/IwNT9P/jFXxhs2V//wtH
d6oEo3IgXh9CuxtIWCNSRvRjXwPmQ5dNZ/nSYZEJJxGnOKF6/gy61bSBCkpAbuyN
iGd0WyWhufKgyRvIJTCz55jsFeXd+6CLh9qlPReh5YM1v0CrqIwtn7l1FzpN0dqQ
hsK+58cA7itvo5EaZbeOq6t7q2CMeXuPo09IJtBXwD7+oV52l7uvL2YA9lN0TJJb
mPHKXcM8fk0m50F+yXEGDlkplQNj1FQI7/vwCUyXWEHd5cCisK1/Z/KcQqoRj8gx
RPJo0byrl2ryAvKs/XTLF+icUKTqQPbWIX28P4UoTDkbEG12j8qwEkppMZvLH0N7
HvOdX/0oTeZ33T6JWwXICCmwGm4RxlkmZFUiil7QSRk7j9szsbiwEoxSElVCawTK
k6HN6jX9z30PaT8fUQqGo3Wk/llR3f5K3GCI26We0VNXBjZMYRwb3O7gxTBKRxkT
MPTGNK8OASJbQdWGMPMqbdwBYyP0LsPf1iI50TynjnVLEtcCvTMeHCY1oPj3/wpM
GKbtuUoQQ8vWztc05n8hLPZHW/md6V+r1Yr+kIAAySmtCmxpPM/RoalnBIKG93hl
22attVf3FCbBrZF1CV72kfr7MklhDpxDDf5ll6mluJTACCf/h46hIjta4kb38G4m
4vrBhmUisUdeaVSMwXDp1HTLmpi433gcwsATH3a6xxUk1ZzcQ8vW3sZrK+zIUTpK
4iTCANWNuuhGDgYzsw505A1zEYv2/qmqJYR3sQkGuW+FRU5z216Z9+eat5WzuC45
2vcHg6lPPnDoy7ml1lpVbX2sBjIrc0giz7ooiAaVBz/fYqO5Qo/U78kuHlcyIam+
gz3xk8nxiBWt6kmL0KU+JjBipzx4AQebPH3ysGd+tAQNYbc/hYYsFesvONP3m3vP
FER2AcgVess/CctZv/FaqWOUiWmG3GJG1/KWeqXEfhJcej0OxPpFaRo/jFHQ5uGQ
PuassYCjFxY/sqaHZFjW0NRUPABnkT3tm+ui3EHJVIRI/OvADAGr3nWiZl7q0Oj2
qSV+HW1gn2AvXdAKKTzyTvb4rgp+YYWJhz8H3rwsVoS5yx7Yq5ATLWbKtA0mRI+c
EYj1tB6aVIuPOR58/GKLOhJYJmmZn9LctsTxBmO9CQ+l1kM4zyUr2ORwWDtDwXad
sn2KuZLQ0nXnA3oLf/Vh2gHpaLgV28o/eu2biruUMHJ+F3t4Flnoz0F840uYwX5d
6vwdt9TZSozO3DFIPQ1Sh6dpJK7/neR54MnmNMOWsikipLYwC6mhsysBMPr+odLZ
jD3qxgkRVdBzlvK0HwQJhHeUSpicA1MagDklt6JGXm09CMqJOtasYDyEnmXwmktz
iQDSeCDwgl891jphqf0meGXTCQMsG4RaD5gjbz3wVFmXCt5sV4PNcrBf3l/L+OYq
WM8kuFsxRocEE9baFCY6r2B68Fo99c/zY3TXV3wAnwosqENiqhkBCX+CzLNuoYyw
CgyIeVDBez4b2h7AWSsuBDNOZ9Vw/wkTtHeAHCXxY8oeNxKmUuXTDogjAygY5u5c
znf43mV6nxSCIND9hw7cqKvh3eNOc/IC0RINQGvfhgTKDHp1XAiKzbnqsSmtIDcd
WeC6T56H/NS9Zq7tGk/ecjePBHgJaX6XuQhnt4mB9fz3dXdUTeBL0NZ28tCA9iey
ktgucsW1GN3fln8biQYO5av5YJLW0yEWolXgRCuFL9VEVXE9frMEyyxEQeuq9CBV
RGFSGYf/wHOwk5442axudWWFjNrDBgHNkMQsyZMvwo8U0Ptk/CdFoFsitAqdmulb
bDf/yCL6JNAYBSi4ZCRP4PQVGOIalWwtMgJK6m/7FYqQuTDbDXd3TyEJcMYbQrX9
Yz/WHDOg1VFEDvgbrTRiMJRgfmHhhCjTnk2G0hkpH5KIkNe9jnQD73X+z0bDWw1T
ZUh17uMTOjmIe0UjWrtTBiCpcRBLbRCNaiZj/ktsVxyGuADcurdkkwnk2h/3dtye
vzS7ypsZs+frL37qe2SkTHSA+GdxdMwz71v8b+Tbr80IOujxIyG1EOvKxjkkhw0j
F3p8b62NZPm/wmxsddDVZAywW/LO1nEO8PdtUal6AU7XxKej3NUlhwcVxmekgxWT
HnoyuTr3L2vMUFYlKQyIfeUWT864cndAlGcz4oFhdl/ne56vfxeO/ia6Y3qlqIW+
xRpjlv97+DUQXZilY8oT9TvNTI3UExKO9cKZz0ySa4F7Mi+t5a1MVXUjJKgILsKB
4MTfQX9aOPv1hZrbFNW4B+hKmpB0J7+SK0oVjzDgRLaaapy8eLTFrKuG61w5PZCW
d4xEfcGAkorm/AgmYM9Y+IwSPESXT4h2hHElrdk5CqSBQpXaI05ne8AgFRp5O8gg
WVFd7p4UV4yA5nhlRvghAjA0oFQv9c5BsPx9epCPP7UeQIr+AzQmrLGJuvwcBwD0
5HtD6UjFHrl47eia6ClELVsgot6JVVlZHVkYOx1G1LNttzoaejvZniP5XH68tvGI
rWTz3dnFx2BMjCKj9z5FE03s3bIH6cbH7v/zpMRlFaKtIrDzTMSLQJ6S+bSwJAXM
UVDkoVJvJmdNtrWqwgA35ZJeFi2vJg8J4AjqPgDWXV0krIfZ4oei4guJB8lHZcw3
p/aPgY041ssHpsB7I1Jt5KILysu4H2IDiQLu2WU4E9MjJyhnxA0s7v3GGv3PqUcC
2iIP1o6tkqQg8wYGs9T3OJrA57E4vwYPLgg6gPRePdo0uK8vu8UxhaoTQnZnoMGu
oqDKGpqGFq+ESLZnVofUY8qjLm2YKr/IWUciDOW8E0jlZFT59zJ5hHevzGFPQPio
k+BnwRIFvbYcTCFsN/SBQG0btpYMkUR8FABQlltNfQqjZYCiEVfVuNAhPz8qJ2QS
ON5nYh/RMvBrGdpF38SyqAFnn2XqSy9ESuyxhpxPqsap+EMd8iJiAx5Hfbr2hpTa
Dm/tv0mcxZbVxMbSBbobtgmm0kU6UwLNUrr16/uJEcAK00whFfRfRpuU9+xc8kAo
cAHPB1gtxLmFb9xmnizEo3g08Q8aS+iDMmFJOdXqqyb4y0UXAqbXhPbZmCKCt70k
udWLq6RKMS7lwQbbiFW1Blpr7ITw+zqDW+0fX+0PDiQR8lC3Jn9UrA2vBSlozGlO
Km6dX/eQTQOibH+FDDG4xDjxFS+OS4NHEqYk2sdmbPZgu+wqVcvtMLubbN2sSscG
OiqfmSB4fbnsMj+ZbztwL+IGwOUaGJA8u2x8QOkirVZdkJTkXZvq0FbDI9jSbRVm
4DD0HDavBKyR6yFr+5mQS34dCDhHJkkGoN5RpLp2jllASZDaf4cpDDmiGPIf0UUU
1MgsulhtA6m72yB3po9PHRLy/BaRGbVga8YUAdC8z3YKAxncVjNivRqz4UAXcLSq
J5lg28QgWA3u1rhXKNsDFOJP+dGAJvix+xfEtupkuxOAELGCKgD47de0Z3JFS8bX
qs4K/bMifVZebu81gAsT26mTBrX2lSxKDWyNA6iMUJwmuhDIWhpa56L4SWl2TdPM
Zx29EhyRIOIjSLav6W5E1hRo521nZ6WOkTQuiR1TftbnLfpE5lf8o+gMkk8jzXOW
eeGJGG508nNUbsQ73qe4PPhsK5L0D7FjiJ0Jq1cmxWDo3Dxv7YPiBwDg0PPnR7WG
gw1kLeR7fh84IWJ2AdRdWIUzd+VCL/SqTJR7FtT6reJ0l3On/hLvOM1IW0zujmlN
WMFdkQmwnTxZ8zu2ihW4ESe7DFNKGeKFDF6yo9LxFezoAt7/8zMJAmujVOtoO2fc
H1QmGM+vJPO4kycDOoMmKt2AENUs/3a08wYbYeqY/8rbSHRhWhfBU4LZPUg3e0uI
Fo/F4Ei7l/uSFwzXqdLG8A9b/lD8fRjPtMAfJZkl3n/rI4l1S5FMnxEg8YWRaeFL
j2X6+EJuJJTsZiyTKhsLFLb5d1GnbSaw2DfdeTWB/jYU5wAVskdVaZkYEIlcwEvq
0F10S4IhQDYh5UbLziN9RbUkQ3LHIFwxhvMWLmhxcKrUlnFnWzx3Ku/b3QU8OfzT
r73uFOjAz9n9NtlfzR1fvbeUv0evIgf9uaalUnmGbAF98ZYwqmBENur9Bo7AHY5J
F+lzQmxGDgu/SRZuKrtijL34MwYiOLovzqcZdcCNQAcoVAgV5UDRRCEvOZYoqElP
mSN7Ny9RPD7npBC/UqrWSawc9naaKLL7LsHVaQ4WTvhhGOQjDy0fCLJShzSawltQ
2zUT2J5AEJ0cvFRhwpBjtHKDF0Hx18SPfYZMZHVGbVaEltZ3n5ePtOTKgLdJUawA
kVnBtYOLKPB9UIkXzRoq9JQEjGYjoufT2/guEKCt5pFYOwi67P3qeKpPl/MIrDrj
XszFoNlR/MwJ1meF9NswFWP8QpJFKxlPy21IJBhZgJCAhLZdG/iDnHS13NxqufZd
iHDAZTIdDOlIe94VSudFjjwE8cusPmv680B1+r2tjMoftGRRhM3zQtbAMobQKfn0
h8VvQjrl9tN0ugW1PcJCuNbT6XH0KH+PlcxbLr9O6ICqtCqnkgxeeJcYyhsorKyW
6FIngnc9+R86jiqh4tHGjKy5w3vmDvPeyweWrWBnokYERprtHn0wuda1Is7MXzO0
vMSKpHoBkCs03piug2/U3z4NtbZaaWOiObDWVANamtABPK99N/xfcXqauW+EftwB
Sqkbnx8VD9d/VKeapLirzBI7FYxUgtlGAhGhQ9mSZhJJqyekJw0atfHwKwyOsLz6
cNVErG330jITofLdZW1FOaWoppr37J1J11tIsU45lDnrOl87Zpw4p1s1naTol9D6
7mn2WNWgqEFuzehH//mHnaIpIIfZiGLmxbOVqjrJXHahAntbcg8I81XVBGNqFh/7
AE3Fhf/rQrY2VNAwtX24DM++dtghxaX5lq2KBx5R7OIiFLDyXnP8+Dg6LkNB+rvo
L73pTy6rL6g/x1TCGPw9iilgTG62tX/VA1uLjf1JWvmjLnKjwzy4uu0cuuJLP7dM
8xCf2NSVLegsQ5suqGSv4IbsTQ7NQ6hAY0lBen5xD6C6R1F4Ftf84V7MR2/855U2
whQoiimEEJXNYYtzumt1jpnqr+eB6m4GrkniydaG/I+VBzFKKhG+7DcCC0vv95Pj
c7wJDmW1o257Q3UvMOoTu56EtHnNvBUvoCXqsof6V+rs9++7n0kQEy5KsM7LOkk6
soB/d/H3PYGFBQfaCDAs1FzCaWGx6iq6/sCngMAXc3/QvgFfgElhVWzTVyt/LZj9
jTcPsVWOzGbU4iU3XaoEI0u77NOqkIsWmJlgPrtCzdrpgmWRbpqYV1dhfHpI223T
yBXJ0bsQ6GG3quzG9M7v92ptIIL8AjfhZEC6IHxBEWvtRNXJYYr4TGDJoRerNi1C
9eeJudSNXePg0mb4j60nKFrlW0tV46MadWf4I3v9DlNpXa26QIxay5RXbjvSqDg/
Zfl33XO8/1fueeGXnR5Zzv6EXW0kr5OIgycYoiZGRM60KAP8CJlJ2FeWTgki7it6
Uewh1G+5Z6YASzTQPKT5iW7fB6Yd1WyrK33l6sTUQNqmtCbB/NwjzCNj3ru1EQGB
x5UeLZYIsLMFChyUspFqZj61cZ1/Tl9Xog5UEyqlNpiVWiDwKhGT8cG+IFYa4nTt
Oh0PONsI5K7zuxm57/i2AfS8QSH4iAQoOtykLbL1CPDBD3qn7/oaPKqkufo6/w+b
cc8j8lljuoF4t74sskROeJpShwTzgmfAz2F8dPhI/6sGwXFMOdEKuRfVlRsIkUB0
33GlncNJq+YJo47osCMm/okuRIaIrg9IMoKIWkyutPTrKWvg1GZIyfAPaUq08W/9
EVupef3rotyAKgZThz+uxkFvYndhO3DnddDgcUjojm1WgBuYRHF5RTkxoA3VLmBE
Jk1Te1UG3QjcdnOI1Wnb8+vYXQqyY0S+WgoDJNOZ0mrDH/MU6kU4Lei9w6Zgy0TI
SU0TryvRLs/H6X9XfnyMHlkpm7uespY4CmX78ADf6fjqdXMRZNSlXnDVhRbB+Qz0
DQqg0j5YV6Mw4JkjP9jxqVHVdZGWlS06P/nhvbsP2eBuJBLJ98B5XKMHHZnZO630
cvNdo9Fjr7SnBeglTpeP6P9PLPZJZH4NuVNu26a3EKveKOa8Nq47HiFk3+RwUnY2
i85mME3hz9ZkV5Fyym/sH/eRSpSWpL7E99wCRs+X+dXRwFdSr/9k06artGKrRXI2
ODE9giKP874jVBBTCrTJcuDUTXGU0AO2xLuY+Ir9A5DJy3IwpTMxYgkAatqU7Mvf
VyiAYbwtvgYBUOAXsTcARyGgZpoTpLKozTqUWd/HKo21otI58lA6vMK9N61VokXy
nfq65pbMJdVKvjq7JGQnJ2v8GQ1BVa/LPmEcPoVS5Cp6hhNQ8VPSwtsUzNkHUrMy
qhZMdgveLvcI4QwKWSMEL5HtSwWv1/dWM9rJMl5oIIH8keK3rfEnW9pd94D6p2qd
i+aONf2eEfNa3llGoQyp4MT6P1Dnf+q36OuEbW/WM2AZa7BRrWnRvrHNIDiVLjxe
E6tSiP5iyxRTpdHI+PR0kt/Y3cNbPVjzNMhOEy3PBxKU7cPyqcP8EibZsJoukzVV
rnIiFWWwhGTpx388ENRzNADONHwng5yWN6fVt1ZhTKLldCNhNW4i2LWH58Mw8nGD
23fz0K5Fjo6Y3/6yxq3lXzBEIW/ANQsMa5utzOiJ7zyE/NeFsdFkLvhkd6EGep8t
3D93wDKOZXzD/PWMza5kTF4AnNDjuLw0JiTLf56hh+YiU7vbCe2D+NnMWY0suBZ4
H7afIkpVseR4tEX9DNPNuM98nVokyUyZ+fXLWEXgr0AUa3GxLu7t1aKwnKsOXsLA
cq1QcxpSgFhSNkQflDUrLcaWFAkTgvoOeqYNuzhZOgj93Uq/VHkCGPLxtkznZ7Zi
SEVfipWAont4yPUGyqOmTkbqtf1QK+YW609uDLjiu8HFrEmtpxMQCfsN0BarKHEm
xmHpMaORzO/NuVbrTrhXKMStoyEdNsc0ED98aYceBafnvXVy3tbsLhv8uADbBjYy
1uKxhVROPuUAvYxy+Ro/19/QOXfMuxDlYt2YuYCqXf6FzAw7DLxIqw5dKYt/cxe+
mQicFi57gtHWymXBa76I7CMQbniduJG9af7yKFDHns/EMndOSuBpAiZ/OQrj39So
xRPD65EFr0rpPEYSodZg0Mb5ki4KDMDfotjPWDHfl7eQ2Y1DzJG4KvLowmW5dh/R
7DHAc2fqzEjuW/oItefhDitPGcl7rttE6+3WdykXgLBYZVJo0XXsdXvKZDqEvZXW
F6G4h4YmeBAyGfD7GSnRILGV2QDEvjriKNlsvkkCVPRWU4mUk3rTGZUf4A16iIpQ
J6Nyauv7Cm15t0fw7GSxVfCFHqsir6uBQeqxMXEfUS/oEK86gp3I3+lpDOWLdODN
Sd7Z0Pn7YpLtALd4yuXnFVuIMmHccM4UdpKWNwXFsphIn2SdNN7ApQdb1p/V82uQ
niT9dcx7kGcYrwGFPapK5GAOg3E5dEYVLr2q2gA3f55nGiylwm22Vr0d0E9Ho+yt
KQUPb7g/JN+8uYYOvRRljuIPtf7feapitvRep53eMSr9MxO0Pp5CTSWjE4Cch7Aq
7cbxbYyGEVXrTrxDSKhOdyqXHmM3CKsi/bXjSDDdjafd9pWzsWwDdUktfJeSPNK2
mQvp3vtS3oGjtCYxBwJmQ0PynLnduo6uhqVS2LjFkRilVegQOkmrNNW0tq9e0SEV
8Luuv9lG6ylJLjizNgJuPyeFyqaeymR2whPguw8FTtVdYx7wyKqg4Zw9IrMMt6eV
E/WxFKYPAT/jCIm7sngNIdFbFbDXyAWxFyKD6cWkQlwuKzG+JsdoFjYE+FdjzGu6
88amWgiBSHVGCxxN2wSM1FDt+flaa+XB7ymmQzoGe0kbUkG4zsaPprzePjonLfn5
76+PoZYwHmnkZgeBCqa5TfjCSh31hoUSE5pDTDF83bupOk9gEBFNTD9bPzpsuItw
v/bEhQ9uTjfV9cGXy1KKskyBYOWo/X8/d/6DJIdohBpGUmlynWAbO9r05EJFjyXU
oMWMde5qGtLKYwSmzDoCEcJ/CaiviyB1BB1XNb28DcGZMi4z0gVL3auVhE+TLXjk
z7V2YIBPxQ+hNZbrqIrMhUDgEjnWIkAWbqxIcb2fD2vIV7T5WPSlEESj5ZH451MG
oiMlYmOnma23cbKJjW8yXCAZFB4bVu9KScUzhnlVWiasnzhiFnNlZhw9QJ1MDJur
RxreLPYHHJqc7B+52wmybyOE3k3ykCyds9+MK+x3w1v7eqrvmg+IEHk691sT5fwa
j3Cobfwu8YUz+AbVIxNb6iMS1IpkHPnpEZWykneipK/g3Ava1SLzYde98gbzkUZE
3WnvnxXUxfHH2MYZt4bVB5vDSJtId5ry66bR7qE+pg0MYkTH4pv2Kgh06O7pDxTn
pdxDYBx5hlPJ/fmJ14ni7FmkFr1ezW2hLWUptkjbQRxN3PY9bMhGq5INCypnuYyI
eOOkuHLxp/pF2L1aTVBmx/SdDOgCTYVKvwfWxsFvL9gPeE5FExdq+ImFN4zAzYAI
BwAydQ8yXC+v97JVXg/dqPlO6/LQV176EWOUkst7A6qVdasQ7rORfbB6XuPt7X0G
bn4+XVT5ViizNHq2KieRwDmViQMCc05Ri1/g4FMBexHnOeXiNYNttLtuBE/BqA5M
JP8cxjknd6gtl8HKLgDUL8qqVWNqFU88kWXrINYaFohPEcV5ruMvZh9kAOUuCPqF
Kn0aXSPC/vvKLJJ2lDZYm+z3iy3af/Z9uLBBIVGFpbdUOQtHeue5BYOfatQmeRI7
0xMSu+6iYu1vli2LUW5g4H7NCsfHJXW/piPBkm7tr3LjhCOCRG4Cunj7m4RSnamb
giOvTDCKJUBhYrzp4TVn4eE+0CBq7K7xOGR+8+aAIyA2yhdxFmoQ12XjEvrATANN
GRanZrF2+UENJJ+AlbivznRqz8MwksNSYOewzcJHxe217nOEy7B86U/nn1zmJd35
ExurDdNfLkNi3QZ2eTmgsBGAqPixNIAObj5XsHn7aCcIagyrRtdnPr6i1h0xxqo2
yP9bRvczpYK2hec7saDpE+Ww469YdLIYWYB3vkdiktcsmGIyrR4+QB1uWlUBRk9s
DDCzZh7qhyU83PdrX9xTsa9FS+3xGgiVvrYOkxHg3lFadkWs1H2cKwM3jjAZ1i1x
1aOKWlIvlEIFgxUr2aBlqxNxkHK6liRojltx6T8yvpWS0znpRM2KkPFz2gSJfzcN
glw3ILOl4oqwy4BsUmawpSCxxoTywUrKfF/rphyyK6+5nwzmLTz6pOgkjWuRDXvd
L3TZg18nMInjD+v4X9SR6aT4FHsiaR6gpOiChg/KZ13HdYho2dqflM5b8sQMy0j/
3k/ffe4UBDLaILn6Hm9d/qwXXGLBPamDbrxWYC0PaXtybTuFwM2CGXh1Vu6UQAZV
hsqMwOPVPBr3nfINetkKBoAV0bmzz+lQtwE4/iXfCsNdO1O1vAADlGocySESHIdt
M8NBnrd7OwOKRDzLNe8vFtRFnyptYqUDxGlhddLLs7OSWRu7++EP2VmhFrTzcOgS
wkbdl4ADflyGoH6s5OQNHUz8T0/7YgyCJyBRGS22uo0LIoI5m/gWOWBeRO7rCESI
ot5ZQVQB6+DU1Ww2cb4gDEKPlvH6aHLVMr5Z7PfTqkPILKD8qOocOkK914IQFm+N
vEzaCZDTCttfrzxSr9VjD15fPRacEcwnZRaTBW0T3cZO6wv4tMqGrD7JK5HwUFKk
eD6XDd6RfcGq4FE04PiCveg77NeIMKSBGcbe99KT8HgSbkxlFPOkCZb+obe0NYba
xrjPRKWUnry/a181O3JJEmN5+K7ecFyrsG7HwVI8K5BZEJunv0WuPAy0TYgNddVA
nlbXvK9J+noFcOXdKUVjE3cqiv3QFRhdNyWCHVSGbPc4FT+ty6pxyCSCeroZvTRZ
Eiho4I3X4O9LkeR3wKYHZlb2jKcxaiCEkltgQ+Jf/bXOYwA015RDy797tOrzd3IT
W2hnVrV57cVVGGTZHXj0BV6p3Q0GmVoMplrfjdR2pJ2gjHkCfPCJJBmwRzqwEW2U
kPHc562T2/dDteXkKt/It2PqSXMzKFzAelZXky1yQxfaVdmvFClPJgwX0SC/urLx
WIq3KPQZtUNsTB3xCJmIfZLHeA0/vUYwdbWxOAae6x+Ld2ueb1IteFH3yZIpMuey
BekscyZ3B1H69SplEfn/5rUwvAhf6MOmU+0OH99DOoL8UvgjpiMP70hiqmPKt+u/
8XOT9kqwJr5jXGuVwPjhNstPZTJO+zcOIAV9uwViAEnQV/J18++GhRx4zBHtpjF3
PDS5CtXEeC5ACMZujDtVrn+AAx0JKJ7CdyOX/G+uNlddkE6026DxOU7R/Xj7rqfB
iwc6BEUtToRA6r4aCLUsv1PaAuxvIbSKCfVz1c9FrOcvLrhGX9JwV3uDVrws0XrG
Kg00hcePsImA0bGui5H9DiVjs3CIZxCkbhSuxG+Lv6T6PXd5L/4I8P9KSkb9rllH
uDbsx9pfUrMRuTli5czdTdnX4OKRKBHc/hQPGW2fXMe6kVZPau9xbu3Lubq213aK
2xmKHN7Q2qM73SRiQldsKVrV+KMToBsi3EqTY4XdwBPSTFMeOEoa384FxbUNZMVf
5P6xLU08aaXuIA4zJq+oLKFDx9jJwfzY63qDv0l4YoH+O4Cs0kHeD6dbreKxptX6
JQ4A9dkx4QOjFp1XLiZhnIc2Js5VRml5Eb7+D8dz9Pex2Tr8OVZbFbkG4JUolAyv
w4WwU4YES6ULZ1Lq6swJNXRjNdvdTJBunTZ+Cs0fn039jGyyZWd3fWnoGrQKkTMz
5aSSIqMpQIfyBSpwuaIfVEpHA/Iz5FjsQ6LGyyVitklcrTmjSaWhBFUMc/YcATte
5hrJWaYf/4+/cjZtUGHwaZc7L1oeDsjOCstzlWbIxvxvRk+VTwFhYRjkjzeRlEdz
AtuKUfaCmiSnKT+0Dqj3ZGNpd3wlqDZ2BMRdIBwu+L6xkxaBk5NRcN5Och0p89/u
Si1FCY61QczVKPed6PSbQfXWs2cFxnjyD3bI/+qDGXQePQstZ2hi06cvHc4gnkNe
1YZTXINIwKnDxiWPO0NckvqNxsUT1MNbinbaeis3z0EFtY6z65ZVjfDMjV3KlfbD
aLgg4qopXlBjDkU8KxbV0Jr3Ua+dlMCW0Tzj89zEGj5tlfE+W0vxvBUMKtN/1Bxw
GvQbDtZt8oSOnJBFBc6mq04iDTG6SOS+A3nPCeo1c+/UFH05UXvBO+A4VKXCt+jM
0ILrctP00e43WmI4f0pgcQr/DU7NeZabllw+galjNWkIfSlnNb1fUidknau3V+Oh
hoasFzQmOKOLYrN5D6yG7zlrfDOBVdovHrS5y4BhWj2mnQm4hoNbUUF8tVbIZFn5
gjuiLShWj+8hJ9Rgm2WQUM+NnMbWRlpUFpoCh+YyT9ehSQMDgLKFw7kZ7kbfsPFl
YaWOLTHL8pMT+9o/s+YIAvIOMB3zZ54hQHRnHkOAfp632R6A04zVgBMkSP9G9n09
LWaw0to459fvjHvY1HhwwtkoiP0zUkUnY6pfsYPCEX7dyIwHI14T7PaMVs8LrLRL
eaBzONmbRL6iQbjDw2WhE/9z4Vg1kV0aEcpDowoE00rdAb+nHZl/xQpjVHuqvFDB
UC5ABUvMv4cdYpANshMInahVtZo8c/QnwncihjW/lCQ7mhPFTkSyw9+PxkuYWtuN
go3mxolzJjRy1bkqQE4ZiisWf/m1o5jsUY4QOctqxOYzm/VCaZ9HF9z9wRiTEjjl
+RbNsxCBmQNFr6NRcEZs2dWBYSyOQuxLvyLic4o4s+/uuXol0bapj7cIm+tcZ2Kd
8bISy3d/fMNA/eiJNDcglFp3x4wGTDEO7crWc0946DVEw/uhuvkAA6eySznY7E9w
Y/Cg7d5IOJ27mL56nRGMaoSwpFJlEAwhcJVzjYNa/P9plA5/aI4Uh5O8tPOL1nBV
7GFncKxTv0es7gcjsEeOz+XZ1pTAX283zDrmxkzgu3qaqtnT++Wuak10wcL1V+5O
rxP+NEAw0/8KbrogCbrbihNY2I5uV2ZG+Q3odDs8FSRBrUShN7DSVqmCQ/OY/Zks
8oPgCzl0MZt03vY6jCDzWk7hPHBtUWhDcRY3z7jR0Yd71cgxbqXCFZhBHOHvCPv8
eIAUjpSbc/2z2FEsYF4Ner6uCs/TYbHrxtxWq3TIHzDJGh6hy023JJdJqAC4iQti
Cn+Optxv8e3cFMKLGGrg+1ybb/RMTxxVS8JT9gsIVLgnNgp3jIYkunYh0LLenjQ0
I0hZjkF9H9ob/ZlnejUHZ8XJxUQxkMoCIiR0Y+sUJV/CNBzwJRcmmMIxXh7oHVUc
UbysehLOL18QyzCQ8G30BIye5gPFwJzOZPdf7+53LP4oPmmGSV4ElpMJ5dl4tCt4
S/4J6NIr11gSmyqCCqRbAt6UeiQXZ0AhNEyE3fnbhHkXdfyoGzWN4F78G9Wkva0s
YZr+/lLZ8MOHWItsphWeqVypGrNaMIjDJLr/Yl/wJbxlfBVysKqGvB6cMA10JM7y
+bsobX9Mh4LHleUNIRfmUMxrQtORIPaJ2lFJ6Fk1PywpHtVj4wRQc0Jyiiyfg+C2
ZEl6FXFVZTYSFwgPmCTSzWvwqabmX9PZ3SLdLhEsAoIRAztvTL7XYZMxWMMago0p
xi/0NQKNXiTGbgaIafv5syKwcxEOyN7CxagxwcS5hUs+fGCJByVTAB+6e11GzGxY
Rfd6xzcQ0mfUTdtwhbnF9jotgmbZnHrllLGCOP+WKVLjn4kpb2f0nXSVtVBH/65w
rkSx98i17VMr7saXs5B+WWkPAEYJY2z52Yy+Z4kR31I88BedSjbJjYFcCdebUrKg
q1oKJ93IJAte54l9Wj+qhua5Tpd7Rw0nntKnamqMP/aYVTeoxjJYACCCkmAetpVO
rYST2wSd7z3qymGPTj+ers+81rBdoC6c59HahvsBebrzrxS1pc+UU/yjQAvZMl+9
8gTvdxDFPuzmLL/aKVLF0jXIzuBWo7/Qh6Ed/PTF38RffOPXZiVAgO58eyFKZcvp
lfMkPUAPAc5zx4X3Y9n5nXZpxrlncCIFZciLYfmvM9pNHX1dC8tblroGKrRPSYiK
8ZQ1l9+vaotJH5fOPD6RN9M952RaKQpsVVblKBpDT+xuQ0Pc1X/Gt4JoDJIyd+9K
NfJNnXq72sAIXya4bYuFKY3vo+6uw5YNentiQ9IkbN8l9AZDT4fLYWi/hyTqDS83
WNXH08VIHa6nuf7zBGQDDQwo/pgwh9VfZ+LWw7KW5Hz8Ku9c5F9RZvDJcRUT8AMV
9vVoDQsskBMh6DT0mOVpFn0uT2XPi5Hn+dXoW4XlBWdjV7e1TC4mFRd8xEjxSCtG
4L/FJaNdMsVldcmZ/VhotUKV2EVSi5jElIQpXIrKMDJw+ere8AmR8FapuR3TKWIW
fUIznD2d57yZxLuyoo+S22sV/WslIUXfFTuahVDI/DTAJo0Cd48HHuD0zDqqH5ke
psmhoCdv7HOQSH8RNGWeTh9vsqUM2x9wvSnL9kHGXH00PY+rHIgfp5RLC8d7XJDh
CcJZdkb3YkwNNh3lzsbeYpeALGDe7GHlieHQ5BXgqMnxEIowOHl2aQyV6YB9xri8
Isq20YY1aHbWy9Rs7zVomnoh4k1/6cUE2VRwmIV46hI7u+2mIKlo7j+zk7fsoQNA
8CHhKu38IjEe6X0unmllHVR5nknhG3XjU64I26qe5kqDe63DpbjDsoW8DsGJ9kjJ
8IF+7iYiooWFE7mQbXhYrQTZBR0py33ausXW+ont+o0Ww/jqsmNce8lRMyIc7y6B
NupZZF++9u+dTcq34VPSTGQ73fMYNryD9zKsBoRaEDRjr8F5hzWcff0Ria2I89+e
Ma/aqPf6f2JBwra/l9eCpj+CLmuGaO2TvPZTfBBTboWNrjPTB5cPlNdh3UwUAjV3
TWdHN6NswseIJMxSrEs3b6WcF2lq9cB7pvVpPpX7kJorSLiBRKuPl7tVIq1oGDJp
ftuQhwgIQ7YBXJzjylTnFzsbeY25vCtxyAK0A+JSuqYcs9qvoLJtQDzvAjJoKafM
IbBBmmJQXdeBArOjh5Fg8t2JRiVExmWd/WhzE4WfqOY7HmAoS3PCplyBd2uxNYy/
RLuvvz/Qw4XvrlJ2AMv3XfURDy3vSIVg0Ckx4nuKWRhzQqiUzg3qrF5i0hSpOtfu
PFa4NQgyAyzf5O1ihf6mtZWiMhuLLQl2yIyOHHn+XaGk2dEvRlsAuC8i0GBuSiom
Q7QLr/LHI3hbq0Bjh8u69rpeeLaPWMDcGGxBP+aR3IPzZE4W0wF0WtQJ4XJsOAoL
2efIP6l2BHINuoUK2lMd6qhUs/WzrT+QsoZNP82xQ8pffLcL0vFctuylivrghAK4
vKRSOH8/S9sCK1DXWdfNdizxneRDF3GjKdh4DgQKmWfi/CmN4LpBoEsc75Ib//L1
N0Fj7jxpg1bfYy1mm5GrHMF7+4yF0MEzjrORrLv9l/tBGKIwh01ug5VheLlivpFq
2yCAZl3KoLX7o/EnQNQcbFHqHioCj0HfmszM4npuO8YvIxOcThKCpO/70ZnGkCUD
+6PrEyqapj/2n21MOl9WNnAEDjNET2f0j0cx2UvEfSUUwtDu4sGpt82oq/lSuTuO
AyR3jTkqDDbUxbns1rBdD5Xv35qwcp7Dn/Jp7aMmVJz20haoUPSgMO2hkcorYSaJ
8YRxoFoUc5sdnj/9qilYEP0O6PbW70eXgDVBohXmIM3aPlR4V+3DtrXTFh9XVBvD
ak84kYHZKHfH2AFf+Md9Z6uwYg/7c9/6ea+LdP78a20+rj5AQXnjrE0BlHAy6uO3
8eaRgzaUsOQDnL00o/gp3nboqZO20fym0MOIDxvxmpY0QE8PUvAJU6nipfROOlCh
22TSKQZng1GJTha3z9yq+L0JkKmVRzyx/EXiVl2eQTSk7fAKCrjiNL0MF9vQLNDp
jDVLXyqoRXctmKxo9HRwPyNvSx3L8vitD+na5eYrdGzCnShFa9qwi3Hi4lxrvzvS
SQDKKG8wEw6svefoemKeJcUvRNj3lUsH6HUUDNS5GP3oI3EBvNYvQEC2HwcjQKIB
yVeKqNX+WtaR7/82bOs0SCuGS1obx5V+5T60x5WUprRo1DP6tGkSurNhKdJWFZTM
X0VQF5gmOhl8N9Kiuy1xeHxHo9T1LEbr4NFWbYeYpyIXCfkAWGfV14RX1U23yH6t
NenNORPMHHx8JNYoFfPiDRd2mg03ezUL/rFbtXftSTQAmM+pQgNaT8Aj2taPgIn7
BjCoXsdXDzUJJ/ce8it1PtOPBBPQV47z22tUsWYlTSa3lB39IBtC0RPx1ro0vu8u
FVkUrRLTA5YQbB0IRrz+37PPdz3NxVSxfYdoPoSOe4jI1BZsW19zW0gtdAu/TBKQ
MEX/G6+2DEo8DRoixiuB4/e8YTkijhK9EV7+PXUrw9e4woWgmxCG5Ap1fq7W5wSD
h7a2dP5JxIr43dsohUdAiKA6XQix+S0n9zYsZ2lo6LLHqlGFPHaFw1WjGtC9h3hF
2PjmKfst/H2E7ORARb2NqoH0h4RgP1uIhPcOqWN09ZMtubRZJGdUOcNKhPNNooYN
X2DU6H2lT9X+PjYm24gKWnvs64zg57lCDQeklKgtEu1vUiV/TMaRxAuZa0ZezDig
Eox6Lferfi9x+IVRHoAIQy+yzmSaoemXxWlbDwdk9pclZ3NB3xYrbK8htAEA2Uux
7AK0/VwEkk5JoNwK0FBWkRXKVjzA0NYAu3cWbvq4fP8JtuwaabtqtCxUpxzs6UkW
tAJeRDJsSK58pS+YfRUcsDh4pVx+R7SDMtj/FAzPt66FGFwfU4rjkOuomFdShgu5
IG7EH1NHKkyecQDBkhDdRDYGpZwN/H8N2daF2fIT9QDCKQ3Xdb4o/XLIYYDFyxVT
o+SDlFJr56ERlXkDdbQcbpWlZVLrW9P+yxpirgG49U4iA95hsJxkW0UVI4sj4S2f
Kalv9LPln7p7SmuGJrCq0Xc9lSem/BC1mhjOlv+NPiZeO3tdfGR+w4SbUbiq7oKN
XG5ylWmND8EBrGHi6iEQKbAtiA7sjme2n13WnctJktWcMCUfDi11+VNjXiER5c2f
SgWicTxD0+hY7cnaNuHzbDp66lH1RYncoD/fZRZMp+46LqUI5LHcr6+CuQWCryWv
qKRVRoKi5kpDkWOx8J1zT7XtERT2pCOpcoRQx9qZcVdxSZwwospsDpNQBKiJ8xWr
nPlxb7i3Btvuv6jIqLGXiLMQeRJaD2NkgxVv/v/NDjY2ZUMCvQ3OCAVIxz2O58uF
RHgYdxAw7sxw53ttC2WpYVjSTOXyWROdTaNQoh5D1s3JB0SN5roxRi8J4sNbKQNS
0urYqWXIc1cDVVkzrp3jIKYqmDzFiAg3ffgUOz4/emKyIY+X4C55RZLiuBX2nlP+
CMHdtQX69Ut8pXRvOJrINtTKGKV7CmRMMBlfeB0PTlU/LptN1FimdwN0yqLuEBbA
B0oRpiG5TrZM3iLpPYRfXg3Z4v9sGDzOrlL1CHV3pnw5rvJL4sYLGaSToQsjnOAN
QBMil6gSikGJnL6sEAx0Nlp4lgvKL5PicfuoS33t4BVlUvyDSmFDNSdH6yz6Le/R
pi4yWIKOIBSBLGglR4q/6V4ZDbuOhUnsIwJUlH+8fSGB433IuvvyAqQ7PG9tLSdJ
19SFeE7ZjlQ+VyvQLOoGzNgq/8SyuNCIPYb+NFFHK8jELGDdwFPxKYUVum/k/uhJ
RLv7hY5A2Kwn80O8p9sgLmATTOipX/Xpv6btUSsMiFSPUQLPbqGOysAz/ovzBoTx
qJixCxdI5KCSs1MRC6Oe/ySQW+MAjEXVp5BdD6g2h8b1CfCkgW2a4INYOGpW+aaf
Hz8YFE5KIxSElVaWQXVaUiCCrnV77PjLcdICAINaktrD87pKPTu4mTo0bdqn6lHm
t3z5pdhan9uPVTedV1xNIoFIR0ykevXMp3PKADDmiw/G5KEAGBwLy8DFvmJokr7B
vdVxBcnNwlnDdOCt8wcZO8ofXIt4DbnEvRlTOKeLp/ku9X8RmuPIs1eETuGgJF+v
WPww5W35Et+/WY6ZVXvnZPiRYoGH/ozp6e/OY8g9E0kiJXRoi51bfztXuxLsV+s+
evd4AtT2bWcSSU4x2Hjs3245c5ydUkXR4oLenW/k9/klY+c2mCZOoLCRwt9yuCXi
bJz13UnrcdAss0QDvdbHDF3zacyugz3MYnceRXgjeG4ZcQFx0J+W0yL5FnkzGiZ2
WYtunQbucG0tP8ATVDUNpeobUf2rr7yfDpRR6uX2HlooZQIdTrfa4/rdhOJjSse3
sWZAcGD7R+8y4yLfVg8DDV6LAJI29NWvyQbD9ga54V1dQ7heECrrfYKgSznBUl2H
N7+TIKprHOrGjOlHnIK9v/wo1rrjzqse77svB9sIFc6wIK+wvh7gE9q65Qil9YQP
FPiYXBZib8uct/6I/SWd8qkGXn1TJT32ltT6MWdblBOx3m8IPfFF0/dpN67Mb9hO
Ojsu/hqawRgRxVN/YC3NE8ZManZsSG/magPcP8V1XTsMbtWN4iioyAbmT9XTZns6
zZkHlU1l6V2jtqQ6RZhWYw/GuFFu6SMWWVBUKmPnt0vagf6fz7RAl3jxVbdlWxzD
v5iVKfXvmQmtEqrzNo9X/a13eiicBJCUq8oU3kFW+aXnHfXAeWzxqNiXqyLBocFq
TNHur/XrVbMfvLJsf3koDzuKwMD9F63chwn519ALHsHBCt8n1O674f+ESvxzsXt8
qvOM8d+sGxRwVh9GjnlOC/buAy53UiWOcxyfK+sag3gEbdUIMwYURqtn72UdtY6l
Y3IkFOYKKE6zPYbg+MS9Wd56vwdwBy3SJEZkYsO4xCfWsQrMQcqSb4v2dXEsuygy
9HwsY3S5JmmoXeSCnlObWxZ9l+zACIqAlKfsaAAB89bVV3hsBzrkU5qdj99VJdlT
swaGI/ztRShd7P35LgF9tPruByVmf+/DGbwB0OTvpgW1pQRKV7bDI+Fr7G02KpxX
F+CiwHiJf/LPjaQGKAa3/JC1QD77udLljcy/rPM1VnHQyOiq2hh2RAH3YgXeGxiL
2f/rrEnWytHPYFO6e5DkBA4aVOSN5VcjkDnlOzG0fZ2q/KEioa+BwWOHJwSs4Ovp
ZP80cEGPAE7W6BLlR2l8SAUicrLIq8koXukrf/PAFSuBqCzE/X5STvn82VMRyyPz
3sUfcZH/tx5nYfUcGEmm0+u5Jbh4vmqCZkcXPnM05N0BYbMKEaCk49OigEe1keoL
zPN7p2QKRxi0ceZIEADYmftMxdQTO+NE/BVk5pTd5gDZUM3tAlty7YaDd6bMpIai
LIgh0hz8+JdCIzofL+lhNKlJaNrblFYTEIR9dAclri6ZX8Ro9051ad4iFBPnk8vc
DTolRjHaK0V7ma1Q0ADUrEPJaChGT2Dyoxy6EYPS1mRfwiFMNI4/ZGnk4F3n6q6u
UnSA8iBlMQYmBvz741zD02SUCUK4h7lYCWrwOvBP4/8z8ZvKedoUxwS1uxZgZlQU
hJGEn4/AFwonTf+CsnzRz522Q1fL0zhANN/s06jW2HTlCPJIMMCnBPPBOv2Smdju
8bRDlTyqPWYcSh3pipkIsVAWntbg2VFmMJbHlJjjxQThO8UCQectAWP9NnG4B7U0
HCkBLufnlFbVKntqdW3gTSqNi+ln43tCLbgQ++p+bCisDnpmMDICKxDbiPdL1+2Z
sjRI8xE1nlFHfZAPzQAPTgx8qPklPp4CgMzYUF1AyYTMs1K0hGPBkUkBr6pnniII
+K9AJIMASSc4fcVFwi9Bkzwn5YvSpbf93fGMCkGiXNXL4P45M1CGjYV46BDyxjuN
23ral+R8NPvMD22mDPrWooArWEWhtMkqGMKceuK3XbgECzKONQlHVaTsq6HSPtUd
Qa5saqqWHKmG2gJtTJgO72mWDYjG9GSijfhOwXWF1uvx7S/NjC6h5cBtk/ptL13X
tKkXr+sgaxI88EUNLzbZScUydyiM8lFId63eGej6IKBJbsZ8OIoILXKAO9GA0xRn
PW64RwMi9U1qGP4IiY+67apHJEBZDM8xza+E+Hii/PF/8Z9uC62rXfdulsHgm/Oa
HRK5Hps/EyNgEMCwjFamZaHjgxP8pHKpd3Dp96iZ7A33tRMJyUfYcsmWA0FoER92
l4TEBL5JdB2O7DcCyx9QlFBq/h43Ynh8Tg6esj/tccqq4m1YT7YEhNrqAJIL/p7m
ibu5f+wiaVcIYq4xIYsf7vVtaNxpJkt3SxRwW9SNIqVmJnaVAiVpqeyoHPY8PYbP
fKew+Gm7ms5cr9aCRNL/leZLnpYIKIhJVBAJiQpvZhg+VcX+73Pgx+wTgIusGAeP
gwwnKYC+26WGOSWjoqlUnp1k8vc2LUFJ6oU7VigzPNw1XsXDrViS6Hc1MMDVeRn4
lTyOe7iAP+hv8vUNYu541hgbeOlXAayuei2oyLCXZZ669Ada/IkAM88kIPnsMFi1
nktrIa2P/dnKcxXgNQUH+sGlksMh8Zd5M3i6IvpJKyHJfvhGy33XBeVjraNJmB2S
VWt05lOBGXyfMkOF1mX02iqMAl/UZby5TxBRPSmcV8ta0hZw13nON7rXPaDATDEV
11XlQzxhJHhlg5KE2XmnOSG7zJGUWdEBCgCs/OyQWeF2Wih2ZQrPbUMmxK6mqY4A
quxj7Xpg9kFoRxW6J8Eb2Dtfz8E04HwP032HucXWP+k2R9Yvx5k3HUoE5dCTJGux
pN8aM6vM7opcIU1DB4Arlb9923mxaQlmX+l9V5hj/ZgP/mW6ttc4oG6J5+3XXp0S
X8nv/HF+F944loFc4GyCYpuTyZho9sYHTiHbFPqgKk45baISGMdNL6BS8RGTpgxo
1VZBX6y3MuSL4oIgmHyBOAL/MpLExYEO5MwuepSbo8jjYNiwD52MaZiYNpdcO5mL
fasgD+RMz0lfchJfGkeC6oHObgYOKi500hrCrfdloA+Fwd5vojjcDS/BwvddUncs
zZF0qNMa88w08TvwAzhc9NRbCdk2HB6EJT61AyRdCZ50Hw4dwX3fYFkilcJKsNKB
+I04UTK8iEKWkns7kE47c4Qhj+W07VbU0Dvv13lrQ6CuItG495Re0CMeyJXeGrTq
WuTlk9T+msVJ1345wxj2omjivB3N+Oof/CFqSnmpD+v9j5t+8PFg1Y12IeIbQR+v
/53BvdiWJLcqwVLTLmCLRRHj039tJE3f3azvnB8XwGl23AXT47P0zp/yIGEpMWjk
6zleBDp8L2REuU1TiSVmvBTjKS+lZEerLD3bNJL/WlortPRiR5pp+JjWCkLrTy9g
Xkdf1PO8QApDKebMftBEyq+raHZ+pKjX4rD+xX1l6lWC9Wl3GgPZDWUR19s4mbBH
OdMkLnO4NqnKs8TLX0IO38X1fApcN9cR/MUSQAv14a0TnOsmbhRKeFzp7146ZX+D
qiy6GYj0FpCXgOCLnheNIAbjIZP7bDAT7pmZvMcZ1iAkRvlgHvLMLOv2+EvH5ATw
liYwyOjJfu43sqUD1CwdfS6YYXABygQ6Fv+An23MYknpjXHY7TceXkvwl0+v2c7K
jqIfy69DxNqzl72QLnQceFkFu94Ow7iyfcVME08ytkOfxIsBWQOnIrM5H0B3hA+7
CBXNDEKevw6TkA/oAy2zGelkiFiYFOd82MvZwTtUEZRrcb04P50pfGR0eFz9Dtkw
+OAWTm36T0PmDytNymt3/C9qRs2wuk6cSkgdlFV/kfqf3UqTGe6kQDNrM16XnTq9
dKhr0MRo7i4qjS/2LWzAiQaa1t3H0NxhFRNiGTCpAhVppFTb+E9HZr4HFIQNZTwL
obDwzKIQ6xjOSBy9MnqJF0Z1iqf4U8CK5OWRR+jiPFLYu0RvkoNB3TA7qIM9+Kjk
h5l/I+O/aYb3gv/8bfrCcFO2H8o7xhTyEnlSb5ddCHX/gk1zCk5a0/2H+G2eVaES
xhfXA+doQ/eYuLf+GyzijTtYB4S0EBDDOxZRC7ks/kJH9iwzyF2bg6NYRNcAZHIr
9QJohzrC/KAMiWcWe3ZanNF5drQ5t8EhVfv3eQ2a14CPxuwywFhCuMR8E85sWqsF
fZpL2SfO/gFfLPS4iHeC8THZSuTyBr7Nz1h6DHEg4d1FNsIW7Iq31u11yA2A/3tR
NNNVYwbw9aHa7tXrFV6w76WVW2mVcZ5dSY/xjmWg5mpNtClqhNMVvQXUEI7f0x2y
LQ1ZaZ5vjsp1Bgl4JIUDEkRqcRc6MVXAy+RCUeDPsHTgEuWBnNOK9KdahFjXU8Aq
lPoOI0Dbp8i0R8PwDNFNanRnZNeJDMRVPIKPzSw/cMUx8kMVHky8PdnNjQQTrDxh
qR21foe6wSOx2lYt5Azix0bQe6z3mO+2lXX9TxWqkSkDPY1lEfTfycOwgk3Ne7c2
zHbWYb9YYKlI5jjIIahJMWHH4Nn06t09NJsBEZmrQt2jlqVM7qdCgJnJc3gH/cId
Fq/6MCl9AJMmHCYyhUeAVbbsV4HBPlTi4V9iwxq8asafie5+qmoyu0Ez8e0x3NIB
BSIwVHJ+7ixRWXd2FMBhsoIXcDDfeKvbT3S/0ItTNSmHjDBakLWN5mfC+8zf1M/J
Tlu3D5ViQCkAyLQu5Rn9/H4hkyX03LFLSs/KwwLk74Ruurk/DpyFYwOjR+lD6VmR
298GXcaflPtKT/KzJs1wsH2wz9GsCHkh5jeiewH5LZhhefyOlh9SYQtZzzGzgjE4
1mXLLYBFuLgh8170GhlypqlhbJmV3I8jOFhrtWVztMoG90SUpGtFKgxLG7sjQ5C1
lhHweraK7Yh5Hq8P7zfwu+CajIicamUVIm8PZ41tR3clU3hSBSStOea7lKV/Zylg
UIBMzWIE8IIT6xG8zdAzWnBxSiIYRGefNT0jVdNuWAwilX39gUqaPXNLN60BnVEp
1J2EH3s8HQjE1IQlbXvGEN9S0YI8lG4gQ8/V+uECfwyFnNiouFWNj5owRxY/fS8e
jZA5oi7myyp2RJKGJMUdsZ21vAbb5qGRrZCmYMXILq83ay6mOKQUCzZDTKacUum9
g5/lmRS4QTD2RPA4PEb3FphtPHGq9aWcAi/nohCqhlh5M6oO17dfRG8tTYa9jwYA
7cG7ewGg9ADe4HrIzbCkMkvjqvLiKS8dbk2LeiQIEzkPO+DC1x4JC2K5D4JwhyhM
UiqmnoqQLjOsYaOpjatKD8A7QQWgtyKh2/zR2xXGA+Wul3w4Kigt9zEm1tWSH+XD
GqdtlnlXKaEXPOnDh0XbnjIbiV3WsxthTOV9AijXx0zSgs3Aav28QxIjUKYmic+L
a+n0Yw5RPmsoFYtw3vkCTOuqm/G38NMPDzBvAmEhFXYzzj++g6yZWMFsPykFlpRf
X8P1G6yut3eiGx6jkjgL4CUaRcCe5F6FR/UKyIALYGgYcVJAEvWa5Iz80NDic86M
a1LX0N0W/VWVDChwZT+jKmlIE2t/qgvRK9OM1KYW4dgHryshJHHzuDbDxpDKyArR
8iI9iHDBX2L3N13xOnIHPa+460LNeGPdVYtEz4IGvyqaxR11ODSmyOJ6evr2u+UK
b8ynPD5kZFg3EFY+4TorOAxhQPsMRp8qJENpvfwgai9iZa5/bk7MrBX0GUu69Pgx
ZC+syxA7/DXbkzHxNy9fd4Gf1FQbBOPjJRKwf82ZYwHyjcd3RYx219P0Qt47SGcG
dAV132lHS9F67kMFBM3PUeGPKlcHCJf8bDp6qJoQRQRJOY3nkgkc4SbpPy9uJQ1O
f2MFA9ttneKdmtPi5SI0CmNGTAyHJ/vtP1hmlFwaIc1NFib8owsikNlkW1rYz5Ni
ZuR30tncJMmLCf7/bRCSN3kjAVR4RaKz+ZpFftpA2g1gyrx5InvLqWpikP8zVOCr
MACLzbfEAp8ez3hwEFrC9fRWVbUhkOxakSAgzrSYkfY0RkR9MXag0VVpVIP+pdBp
vVgfAveOfDHAakNTna0VqcwKJYNrBxQfCpXxVx5gaey0ENcCEJv1Mgwe1EAL1a8o
MH0rGhrX+M+hHWr5sDlbX+4lizodwCY4igZ/C1NAzakx/wOvAhA0y7vDS6Na/EsZ
5g4cUDjLo/jbeADk8DId0OVJ+omFjvWEAxZHgSwVD4JO6qMRSSfLjaX7DyORP4sa
lMyDChwAdhym/aPN94ihroeRkjP60UU7lBsqMGknc81ASKjMqapnSuieE0d3CA82
FTWWtb7Sqbto/S+pdqmjUB6OUP067U4JcuGAPh5wj8ocFp/5B/cUG9AtQDu8z8GN
FiXmQ890gTa3F22xeGjvLv35IQ9ZBmMoaAXe70TpYS+LtUZd8kKcPSQj5rCIC8Is
VYwdQwOiXNg+w7QtcZVFC+TyzCEY7fVKl5oFzlhbnl7PrYQ3ex+aETUQuhBA5lDP
OBSp/WNYMKsKQOzxT7kXo2s00TNiJeyDIksKnVCD7OUDGvsId+WEmCd0CC+CFLJ2
BMrv/Oej6i2IQ87oX9EPSCg4z9sZGpWLljiu+n10zw4QrXItkC3Nl2VFm5uTjxzs
fgYOHOLDDxuxjf+7ImHhbe2V3nKbqtQgUj9Hb0s++SumpH/fI3igk3VHm3qQASjq
EgQw+WeeZ+amgVNVBl8HjJkZojmAmg9Z+19Cjt4LjaJP3F7t1VlK9MNAg5NoJRTy
OyAsSchkN8vN1OM3MY6ju4KAZoPtfqd81zSOHd+h0+u+3ZlcboEsRRax008/kNvh
LBmnvNXRl5pNaT/yBHfsw1pLJmuGsuu6oe3dujhDzRLky5Eu0P9QllOIEc7sqctf
9jX2IZI1TbPzGxEq+XVZBtfLHtmaVIdCE36lyACE9UxLU/vHiLqfU40FTnmpeiLf
ZxmGQRmBmPEuChxz3UBT7Scy74WXGcFEr2nX+umlfFl9C2XlXld5yHTEh8IHDf9P
0nL5VuYb0WSwuE2d4ZPqeIB8HXaP/QiDiSxd9RJZQBS9L1TJVqHiC14Mca6OBCWI
GB8gVAkNRp9ALwAvI8D0/vn0bkYpt7LJSm8hihS9H1cubL8Lb4dPIQnhUBqICRoS
zuEd4svTI0h2FstpgRO/5vlGRndFQ4s2jfFZeqWvlyL9jVpsDYmVoesQ23gJ4KV6
S6sqwtE37qhjR5S9DjRcrIDsGj1Ww6XOauHeveHYrhdNhLcQSZBtmO902V5kTglo
DfoW8+j3QC1zu64N7JwYg61iqAQZlcEsKOos35qCCt6+5013OgFq92FfFzqOkiEE
AZmHsSONbik7p/lx7fef+P0Dzzy4SF4UjnPmguTXBdZoP57m+HLiSpZ8uTb9bWil
RSakiOFna1pa29RHMGMQeUWZ3tD2HsCtx9p7E1WfGI7dZLLd96/KrlH5exzB1Paz
gXQLMFZsvS1ZJdTd8YsP+SjUfaJfXrIFFiUzs9T9qewHwMomAYp+wcJxPgPACx7I
70GGdHEGahBfehXUeTybLQim8jRdhEp5UuUDBHd3DQxy4VJ4WrDCiZ+hVBwBNpRo
YLqtLkOCuU0DI7LdPwTWUyrgc3bkJXKW27+aCK1JawBp+qkQm69cMOdOkxANfH7h
16VSvB/rGJOZhWrEyUpUknvKD8aRf8631qdiFgr1YVgPd+xHDB5gKxfmXongtQBG
0Grqxi5+vysM6N02ptoYytBTl5Xtah9W8kL8mfCtU8pyoIpfDvhdTKGXjMXcJo3U
HM2dg2KD2R+0ELa47LGo8sLjVdhuWrc/eFAJh+Xmzu2WmBJVWXg8r8pL6AbShCdo
9lGqhmOT3emJcmDFEKttiDO5ZpqKmKZ5En94ybkXDajQCjPgM5SOty0KDl8wHxAw
cRTClP7j5FSb5L3nhtsxpiroA28j+00W/LcQHS3g1I8LOgYN0FV2qVBwbKT8P9lv
YVD8sXKMpR4BSIPvN39pLmB5a9YJcfEQumKc22bCZLx2YWYWnlOy84769MI+M9Mo
YVasGF1joaOTGf+HG+QPtSjkTGsZFAIlkL/Zny201l6sU7pzjJIZ4Ru3OnW7MdVG
DUOSoM46o7lAcrRvyW/t0NPS/nLHm2efB0gkYozr3Cf5BuoyaKF3GMN6KLZT3KtD
UmBfcpqzn43f27Nt6lsc209Jlmnc0f5/O4lRuaRXcPdrEpbzaOPkZJxWoBEPdtka
CtScY8kpMFnSIw0WNPtpg2T8ZN6Soax0/0zsWmy1h659OtEDa2Icumy80PGAJgOH
lP+vHoV5Fo3F9Z/Ql4UbJqwU7pbRBzo/QgckGvW+GAOTWdJZHTJS/j6egNZ/iw9u
fhDIax3hqIDUuX1XlExp2vo74DXHk2QU2MvYwNJOWjSBrK1VIn4QZLHRcCRGLPjW
XbuL5ITv3xMktnRShIi7/8d/KihZHp+kp8Usk7Jl/KjHSKWlyDYyZ4Qa8ZTjQ09t
Ii/s1uwCclTuRM5LbQXXYXxi6BTbLt13oEen//oSUuObWWfGLcVSKTVrwjPdznYm
OoeaapLgF65u5eHnSEDYisbfwgyiFo9u+V/WtcrHONlc8UgJQp9n+k7emIUkPxGF
PiDttB1u8Veal8bXKDe0vIhyvtAyJg4Abco3DozLVoq+7+N7KQpCp7Jf/eCRAD+c
LZ4kt77FEaxeR5nTZKMhGg8mm6+Ga3qRIBGslZOw1uECl1QUu5aEiCH5n5EBdRfE
YD07ATjJQ+17mt1emyzlx3eig84dj/6KHH/PhSdC+DRRt/CmYP7y8J4vdj7N/CBM
8YQJhrLuUnRpizHiCOWLDjlPguXk28Ti+7YthGYCtAaTcRs6Zq/8U+4pJxnIZJJT
wF55k96wMrP67EglJlHd0w5embB6o0vyZEMlLj6lMMLP5rL/1YIed+1KTRbNwfwL
P5hWdYfAFk5V1iQR6LnVZTLtkldvksTW8m5H6Jo2YzwaoYnx/7on3E+RiiLUDEw7
9BPQsMAmvKwtRlfVeUKvaFRIwpDuw7wwc4ng2Qt6UvFcUSuefYDLkDj3U42ypH7e
bnOkGUXI2ajTNswC7607JEwUB+S9Og0y+NN6f/v2pzaiiznvVyRy0DEh30XJR9cv
vrfxR7JCn2IH5Xm2jdxTiyIHK6vqXgRDtAX07g3Q3aivFgztPdvJgE9oeHl49Umi
DYJjb7jqpZXpEsnG/iuIKHOhq2dfBNujbPm/khnrtfGg4zelU4H7X+mHWcDs/Qk2
O2DyWIGuzK4pWBcRTQqmEMdxeNcbpDGS4YFYXKuDyV8dty5RteSbQgDCQvbsgQX4
srHk/tIwIxTdIUOTw4GKSk6iB9efHBcbjLnCeH0bdfIZe29XRZbJJQY7+ZYEZgoW
XF3R0cg5CQ7Z+8ORir+wRT2/MgeZJO8GJDZh2oEBiP6NFdfmln8paPeU/xXPKe1E
fMKvfkh0lHO/l3Dzz9waxFuzBn7/Q7Sye8uYtV2gdL9VKJ0PWjvltL+z3pqS++OQ
DxiyiM8vb/+Gk4ZUlZu0V5LDyR6vXxwVzGVSmPYNtTGCEfaiVIbeDD6z40Yd4rqc
d1x9cB3NOLuftKM/uSiGbJlspIWy8pifFlnLdgikov0D+qSxTC47qcDI2KbuHe+8
GoQNZCgnRJ1s6IHKbUb2NUqGpDUWsrMOwPi8qpyq8Q4FboVmazbeFHzhPDsHQsxu
adPqzjOMaRuoeBu+vmGLlnmIoBLX9u4lear8rqPdB8utLD8co0ksULg8s2WZO0oR
/80z0SXyxWlzkWndKabQrSERz4sx5p8AfBEr9w/TIYWemNRzEAb36qKMdSuW0dzm
YREcsRba3PQXGgLeWuzMQMCZOjWksJJIYfJdMx0QrtfskVmA2aHHuCG+XWplaqzI
ZxxYG45QA5jA1qOeNtskjfNEfWW+QP6ebfHg7jHZa8NCyQyPjdhCgS6ptweyhF7V
GSOGOj1NodkST7fdbGSeTisgmrL7JWhfE486e9fJeEeTNcGCbA9sSZQxphXoKLZ7
u+Z5zi1WkDmfgjePxS8RrStVRMZ/hKUmilMOv0ZUCK8l+YueM9TeENrO+yhU5Imp
wAZ3vN8h1UZbO1xtY+NIgPfn5fb8oamkT+yojrHTY7gh6S5IGWZEO7XApfUASCVx
C9gvryGOxFWaVyMfiBpYV9iInafVBEgHykbK7DoUxwJtLbUvYB/YkLZWnhmRB9xH
MZTnLcJQzZy24Z9QaEKFiuLseJpNxymraDwIm/KTHoFBoHPdIJghy1eUe5nG5UY8
uQmwF+8/QkEGGR4cxVcFZDL9zJlDy/p4lDbI/gwFIrXrNl3ZGvbYjKnhwSWglZ+O
HQVGGO078BWB0UCAOz/wYDhlDuY/dYxf6eWlj122awrE6ocjY7tUJOxSl3L2yN5y
woUbcfxETDH01drT6qOmKhrs9e12GOE01y8kZeyG7/arVvfxdO2wEAjRAyMlpEDp
15lW/DUBO7ZNi7+2UDTSHVcnbFP1mdgRI7KOyvJrJUUQMDujxsXkRTKHecs0e7So
2AujotzGwtIXr8yfsL0ydVHMyfZIbJtjdIAqoDc6demTywMwf9Nm0pfY8msOal3b
mk5rLlTyAGjwVRYEIa4g8jsesxe0NmfMAIm0q7tm2ugqRsbihL5JfWDxIpqUUl8T
UhGulz28eT8S5idKhwEEiYnGBHWU2dfNx13xcVdgaoHAmm/lxNHvZgq8OpxX+xs8
3xQ8Sy+chIgyErw7dNCDX7twckKLL0OZCuWigKX3bogVU1Q/LCC49Z2gQJ6bk6fs
5Z1X7WA4xjp2B0IwtuIYWzg+Ewl4Um91k/p0GCRNSz+KLVM9eiEI/Rr3t0YRDRbA
JxsJAiFfz/tTXHlwqqAxiD9Aa+mxPsbPZK0VC8zu9FSKh/Kfx0pBCgckghMaQGvl
tc1KolnRmAhk0U52dImBpHgVEKh4QcDURppx747hl1u/25TnKeyYLs62OSTNjfYV
hPKOU5t+YDC2YGC4BHCAZK+gMrymxtQhUW+bDIcW2p13NiqvP6kwUJfG4EmL7qCd
h8d+gTLO5MRZLoC/flamh9/s0lEaqftZaAspjR6yN+niyj9S1Le774Uq6kBcFWih
VXm70p8xeXUE+X3bWi1PQ83wUzgitihGT0cuXJOEeFe/IaNhjxCqCbZMEYLFyCP8
9dFs7NdwUPoytrb8d3uTUq6aIHyW+dRwSNBONKMdHWPpBRgZHq9p9ltWOSIfsIRJ
HY5f8hZt44L/vrZd58GeAJrCR1/NKOfW2UGXB72/6O/7KLFTly+xw4R5exzzq8PV
GqTJHB0GakF82hzDKtgm0rkZh+UsOdFgmHUnOSpjeatk2gVGPoHdzvmccPIS/msz
jK34ttCgtWEBjCD5q/lb2w4SM2fL8hrOw3ee1CeyQWLxbCh6I+jm1sBF3E/t4nWD
8WwiV4g2wi3Ol67fJjRpuSnAytmTTNXhZNX/X/DUcLThbiqixXs6rqPDbUvkUZBN
8kq2+7BBE1I/0fpBPY06vv7uEzec7tzn0K0qmzCWg1fFR7BhRlN0gxIIHVkF0JDE
FATtVVDJ0cUFR6SO1Onw/Z3kZbWPswQZsL83/JfDU69mzPb+73a6kKfxKIOwVHJC
sqzdkHkc1mTRYiAnc6UWjfqn6nGhSYBEYuIn8UUrDzMObfuLh8+TqvUfPiChDhl4
sRBQX42qO7TnT+xT8460SgAFkXyUVfXollVH2r33S/j4sCupVyysnA7ddsSN4+rq
XVWKbAWnjxQt8C6byDY9yiMZPmGZsKHWKep9ziJvdKvDNF/FH0heVlpbeFgcei/q
JhJ4YSXSTRIJrUhIOOexGw4RtMvL3ZuuM/v7eMKhh53rdDt0T0HZjuuJCDezjKe+
QQXhhmZOup/V56pDZ4140Pb4HsIzF9l/kvNx020GUNhWlfq6xaIn62U7XktXdYPa
HtGRC4ZIMXfMZB2OrZXKTSB/H8Q5cQqRVf1nalu7ZxC+QJelRnKeJyp4Qqc2BvZR
ZDcaKVGdo8qhLgaX1gBZU9NHtgKBWV3mx9DFpecXyHRCCvfffxwWBLuAzBQW5tio
qD8Vz8PQ6TCRdcnXB5z6TiloyeAL9iabj8T0M7ZCLmvY8Z2MOh6RvmZnL5pdQNGT
9fLobibrkBcjEOtO0+y2DF5NFUan9kQZTKo+U9RJXNu0eaAk+ARhWf6U4SQC6ulo
cblOi9T7MRXQ90lHbYJU73Tc6VuesNVJxITGnDzVejOnjnpRrgw8wyo5wlzRcBwl
hdxeX9/Vwzm5MROxyyrhNjCKDBU1NNeSm/7C2YgYiNrd1w3Xp8EKPzHjf9Ksg1gC
6YMBy183SF2YdlXoL9pgp/8mx1u/Jf404vq2IisgtEn43M7nJBMxa23yQbUwlAAW
oKTWNuW4sezntZLAKzCtkOPBIWhRDakl9+4xrCanyQftE/lLA2keFMmiM77e6EQk
FSoi4Uvk2Jo7ZRErRknUvEsO/6Kag3zJwOHOCVilFiXBtKlDeSiYxgYTYv8yFzJU
Ym/LUTee9G2MQPVfB20Y3rdF31CXCdSCgOVf3YVxcqA5AvJ+cxvWUV0aDYuziSGM
pqd7cEf24zYitbeG8mz/WZyr2liIhMUR9MeVLf4zazbaIz3OLBDkRBBz8oKRta/U
yEqHT7Fl/r44hTLSIw7tIBd8ICXqpWEaKTVW6jV2byedDfbu9SVqRWaXjiLXKH4s
UZj80b2/k4E5kBoXGljZVtq4HuOPnhzeurgPJC4KP9TY2v1W5YDpL7m4xPiPfXId
SPfApJHZwlTagHmL5O6YMk5gcgfeF4mIUZhbejaug0CkZsFA+yf8zn2mFSIphAkn
RdnB27tSPsY3fEUp33zszkAcckI8bpwQpg7+4zPvae4vyeJVO3xopNTEygxmk3+S
0ShZsGv3Rb1atbmKlIAw01YzDg/6utfxJwQ/REzIUevWWb1Ufzj0zJhqvVFN+iEX
fYqSnjLXSx0mBuk8Aywn6on027E0ajlOyTI48HyS1cxv+BAY0NvEGOAggEPmgTdL
lKFT/0Jh7GVcZLSKtZBOODGRr0TQoFQ2/DXuSpcg+IHFHbA45L/dkUhGoZI7ATqA
W+l40tkjqjzmK2DnCBj4t+7EiIFrAv5uCC8Fbb9UM0YVn6o0LL9WfUZsc0rQmCjc
62U5mORZr0X9s7INeHo4ixFnjWBKtAGUYvwmcIzl82t1pYCZ3J9KWPe6bFeUoPFm
+NiBzhO9HZlcq+zwIbV0X3Lk6N1gWy+8uJx7BIKeYShwGl/Q4S8/I4GS26EUWXpy
priYcNFFLDLqVNUXmbuZSYT0dGpr9g2Lk/OYoIUJxhpghQCj7+X/oamEnBbyjhkP
FDwTOUlc3dwMGTbIZpeWTH76za0Dlg2xFcWHQ/M3AfEwkLm/E4mxXay0kNMoaKUM
aR3lpkveDHrgX60I9nawRw32wlYXOHDjAffJuZ46W2tjond6sw2zJOOKMl8Hd5Dm
crVZ9cgQP+qwzh7sc1H1Kb68AaZAdXRoNeolLFQ8e0GgUvbNsEJy0pjAss9yQ2fJ
BbMz5gjbuxZwL+/jYuMWAIoaULkGtQkJspLp4WNtGUmCotnmAYuxK81EYtwLZHhW
9GyyvTYmPTOp/ZJDYHWWcGNj26e5mYYK5K9xAYfjaULc7xrM5YiikM+xe5nFbfBd
MdotKDw8q3Ab3oz7q3OTbFi3Iby88YtqtJ+v0PTSmNxV2JtLSegQnIZ1CjDM5EhB
wNG1wwPdP4PkeXcNNRYIiXEkNFZz6PjyPJkvQtZqWMiOnqr3YOxtYBG44tjpmwea
fLT64Y0OcJnBj/VNyMwYXvawRCsS0ciSk7z9eRNrO6XSYqqwm31pLPSEjgyTuLXc
hXdX6Tjxr+XxWPPA9PcLAV33Dg1UEWwhsr4xDt5A9ptux2k2cSKv9c0cV4xRceVN
HpZtdGR2ndWcjNiTH/0ypTakEH5n/SxjTdD63SIK8y2lcb6qdvJM1REvL3xJv6oV
l7W5ASOi5E2KzmqvnidzRn56kG1L6T1/0FbPy0eoSukwfO3V0IKG9MD5V/c21oOk
/7vpY2Dql7gX2AXLeHtaDo+HT2hg808Z3vb5a5s2Fh2xNPao87efPI1H0gAkIeFt
TAwA8stsmOZQd6LOwhzRTVJPf8dtwKKx6w2gtzMHpUUDg0kAGdWt1jNAJml/CqJP
Q7Ly31aaqjnF7VH/+9VY8gMAO9Vi5Rq/KIhSuXIZP0NQBca/XFD6OydqBenCwGiH
Csv0zDoMGoOEcx0VCxyeVQV3J1MTNSJruMeygQYMgHwHrLgTT0FfSsoTNLp1MDPm
Ep58D1IZFYhEZjmueNE3O7dO901ZmMP/mIJdE5n+2J+d7n6AOlcLC0jIReKZnpN4
hXgKA1Pp/TyApw6NddTzsvJYWExbrcXao97pJNUcc1LPtK5WtQcK7ZVi+93NC2dI
YZ4eNavRdJtVPrnWf/bo46EMuPP+lvoIaMs1QMYj2U8wyaGyMTuFQJ9qSdtgsFqa
4/WOn3I4GYH5CkPlhl8z5las6L0xAddgPmN6I3Dolk7w7m8MXKwwZDE0pqB41lzk
lNlog88ItejidvVgNec3E4w8ZEnpDZFsC7LKzyJJfjBQko0Yx9Vz9L9RWIK99ZIL
k0t1raFOTZgRCROW8m/egQz8KYNTgXQlAQhPip/Jyv86LzVEDZlJtB4GV+bIUjEd
GHfvEJy2174du9kvnlufkfukidVFn6/JB0No7e4b9YoU7JtrKEuAquti1MmA7x7w
QXbliGH6wyqO3XiVXLBTB6lQwBi7CIbceQVN1JfFOjJP4AkVQct26ZnCueg3XfGH
xu2GZM2gLycKRTJlEvLEnVsFCnfd825KFbAFPtCQvKQm/eAKLMdx4Q0Z2cSiYW24
17rxMb7phWggsZdfWb7AikvLx9l7dixOxvkZQxRo6B0kKCTHsGaPR8J+UWhT2b/F
a1U6jYKQ89Qv1bR4x3QKvVNx0gIzkh3zJW6ZsNaoK3pP+mrPFhqGYsSclYvE7ia3
k1sZYDfmiaqMCTvo/KOKFQcBfMz2s7EwpT03AQSNzu+mm1N2fRBoelpqm1vtWdkr
shl/Z0ZXExFWfADvkERYlS/tp1P7E5le/z05mhLx84nKT3OM/s1eDNxC1g/TOdwI
q/JTF7Jc26brsIweQasunFLVxSptPneCGW/jJ7fbVT2fnYeqHDQF+norwO8euC9v
Q25p5Up6Dn2pmWtrlZseDvAA5N+QnHrRJM3gu1RYU9AddJnPvJlhW/uxE1FQs02O
UBb8cgYE59GWh4t+ZgaSRbyQTKHAvFJmdUd1TPlcl6qjHSyGGN+UksW2ndvoxLxG
NMuFsidF8pDe6eP8rB1o2J91tv0gUBfXCngFapyLooqvdo5UboQPrXuQFNp/jogd
mBjtQcV/9hNAv94gxjKDueFsmPETCgZbORjz5wQRlskautPXQ5ZEHuEwYhlE0ItB
FwmpodtFNR6QIgcpTyL8aAV3Kg98sGhRSB8XrYAj/TD9vDNO1UvltWUNpYxr69fF
xfYNybc7h9Mni1997r2gXGdPw4Fz4151zwiQZrTGtGoRCLl9HnLp+6VXJeCMA0Fb
lkHPR/6bBvfDSYmYYbr1moOZjSnGNK/Aqii68YOvUPvb6M9ysI65hZ6357cQQh5J
BW+aSJEAFQCPz435dSgOrG82ytE+XjPQfdlwbkH84OLpvQHIa59R/nqGBAoIzXqp
c3Od+IOw65xuUQKg+HBX/8C/rm6+tRJdF7g13TjdpzeeriCA3wR+O0knMyOEo92/
eom/j2j9P3azskcRiT6BUV0oRtp4PJ3UgZtsxgDuHLfyWJJPAtJ6ZYatGeP/j/7h
RbyfObDhPetN8+w+uJkYuNXmp92QcgAMFDhU0f3gPPAIFbnRq/tJed30HqvTkx/k
Ny1owAlZX0M8UgXeAoYftcVBQxhYy7hmOxfwj4dBo2j46JtOPfea49HxPlZCblcc
v/cKeelYh+9Ho/6Hox+Q9xA4UH8zJ+f/cyJzN0BPey+/OEciRaOwkvRg5H5/osAa
FiPRa34eqHBINQgW1Oqm8pENStWG3frMRELy8wD2XEleHDpuzxKfOwdBkSAPHLMZ
xAsV45x1lbMvHYHP9rqCRyLAQy8WH1m5EpImqHU+rmknAtDaXtgy8gXWBfV2ve2h
e33HI/3R3dH1P569tTkUmhnv5ON3/F7w8IO8i4yoNCb8QrA1jZRKFpWYH9mlxd/H
iuTuQvHQl0Xko7E9NeRAxcf7nE1/kIBlql1SYbhqg8mjoQzK7XXXaxL2sUG/rHwi
EGOreSxz0h/9uAipZYIr9CKQUZwnLCLBcLWIr2LtivrOdk74gJmnOpvABCmalVnY
Ev/vYW9r65MBfFXp1dThY4z1BB71UotCe9/KaH7aA5ATk8uEb4zqhPvKSI0LV+M4
CdIiT7AmaINoClwkt6ueZEAavKhykLE5TUtAm+CAtHcjq26VvCe5389GTKNvQXMH
OmuAiAXhX30mhU43M6Sf9N8fOPeyPDM5opRugUXZBpLu7aPNySWVxgDaVx0CMy1v
KwWORF1Fnd3G2vjqkJ/Gly3huPu/YAQHMhaG/avTzDNQIM4cHhvHKeKzPmKPWm0U
cTKsat1vm9wLyPXFifSwe8vHyHzkBvkuDWvkNOkMZIB9zmz0pIkwFT5EPu1Ooo0+
GNBcKrqe314AHV/C1lI0zI/bRn+bmiClg941ii1EWllmPVclU9zwozkCQXrqcLBk
f6nIHQ+3dSuqEp5cru06kgp7v5NktoH8po/1HnmT5+xSdgLqC2ZKwU7UAQZA/MZk
eR4pInDRSijXPBoeqRa3xCBAMipS1o1QaN3mqK6knvGnztAAfi+N6UgfwvwU2USa
dpk+raFAFomBm6czRp8oOKNZUhBP/axubA+19Q5hoTpM1Szy+cU00gFvllPTXCLo
G7enBg8A6fN7QoEEERntPcspQwB3iXWr93/K1L2zNuX+8zXugnoopq+vyfPTsI2S
7/rAzF7jn9G50aIyPs6khVdBPJTrup8gMWf8K8oOKlOY0YW0nEfWTanJsPmwzlYZ
SB/cKJhOKs0TpMwR8LX7cP9nfRO3gxhdvCcI7ekJo/pAtfkh1HEg8j7Q2fFh+fd1
G+Z/6kKuvjfbdKbJwqHY95UIUiUXljwh2vvv8+Fco0OxjjzNGf63t+ru3BJwGTvS
druZYwLr4ZVmh7Ylx4RTy8QamSnuUa1wXZ1geoCY7h6UbKCYY5yl6/8l/KJb6g/X
RHRY4UJhZBNU4mh5HlDv1L/A3M1LOuEynSD0qkH8zwLcKx+Up4JByUW652dmtoKi
NWpn6QMxVZjS2sL89Sz9Q5l8PvUfgxf51xx0bsDnf2pFytA5mTkQTqTNqG81mHv4
9ZwUS1R/1rZkwCypcr0Kavd3r0Y3d6+d4NKkSYbADXIaz6MTqWv4nIEfLsSg0ck1
IB4Gs8DbMLBdfhOnVldDzKsZu2xXXNkM8BB2EncOM8NKaovWOXBLq9VpB+V9yprF
7MyN/pbFT5HhGil1Lqdo8EHV3/2E2K6PzFq/vbct6GMtg1H/FlPD6VitBVtjjbgC
6OMZfG2FCR5u5DA3mqFDSVgCbbTXBoBgL+QqdCSvo4bCTOnKot06KuPZFf4KTsnu
M6AeC50z7mdZrwm/zGTWftJCsWgJ7QM4QnmdjoyVv7XjH9IjVF64uVA/rrpnH8z6
Apch7A6WNbVZym0A49C3qfo0ZO7nRuqdFdhhWDFs/7rpWa+mdf9CMZd53IzPeY82
rZbe3rrKuvt/7SNvWp+ZqJtn3EybImPjc2zW1P9rHz5TmRbmwZsxFb6p3PXh6Oc1
DivLhkn6qOBW15GWETRbUMxYjsNM6CA8WjWBJM1DKrGnPp+HebtlW9FJOECh0ndp
mGty3/OpJZ7q2gwl47x+ru0BKtRKjdGr+EnTuhQjoqbMkNKv2tiZ09mTEmWF4LKY
d5t+74mryp4YBKJ0nFANLhIzNR5LX/X3PwY5CWv0GEEsz46rQQ4ThUVO4Xgvxmkr
HjArCMOtG2YFMXkwg9PIrWGWM2tCYlx/58ci6OnkOpt88lH5IpHlW8x0FA+BouAj
29LhqtDOy7xoKPy+s9Frwa+1S4j22DWU95wJt0JOW2rut/LHoDCKjZ1AOWmYj4i3
Yyf5h8ZwHewINFgnsmL2m65ZkWRVL4snNyHlNkrcGyDX67fhJ+e5C01yRbQk69i3
P7vPBWOQTUOu97nhagnKhEE1TgVHgGYwISlybR1E7GZvlJ8mAFKNN6jZat1Wz2X4
h5NS20a5uj2ZmKy9OEvo2e5WxXjmmHTX76Xfj4nISQ1pUVH2MD2AuxkmPJ+m+TyO
69Wg0dYcYC/G7MMbfwV7wlTDAez2N7dDw2pSGjbRsb7IMiqkjep51ZZMk9CspVf/
wzxiNn5+5Yxad1qhMm1J2EC8OerwBwX2cAT8dWpmJ+C4XFdx9tDJ66as0SdGfX2M
fg0K/vCETUXljipzekOfki4BXfsHymGXO8axsNUKbEc/5g46LucjTdVZW4mM1iDY
g6c4cmK2Uibt5DGU8XIrI/o6e6f7iCKnhudTOzbqcr3XcA20UaIY6CyKsswzbjJ2
0Cbu3RULdPdW+dGahd1MV/Ulkp+DKCWiwfjbbOYsmUm+luP0O9X3qUtnp7T4zAlr
9xgnb/yVZihdq1ZTAtZd+D4cnGP3zye+RaVJ1rPQlxr2kJxYF8scfsXNNo3X58Eq
YqTQurYJjWsm4FVXkq6rzdVmeff7/5UuHxT04YuzKu9T06loCFGQkUQ4606ANRwJ
pUh3dJcXSEbAgXt/jA8ba/wZCkK65Y/Z8c+6BkurGVNXpi/K6kBsgPGTusm+f5Sf
IrtnUzvsUfes+57MDKQkZpD6s6+0I/bfXQoLqdpNAVYMCUdFkaeImbIKSIwoGdW5
Esve4v0Fndhz01/0Zguw+9m5GsPq/LGVOrJvMhXP32WDiEFTmpVNkltQWShSmoeK
MqHlIjqfoNV3qFO8g9j0SZsImVNF32H5trjSQwy7RSWgfwl2mOsBc3uiD6yAniFb
r57Fhwp7nMGMNeG9Y71QaRd8EKBgMTzHXiuEhDCmxrJNMbXpBldtNwzEVqVVbHDY
BPT/DYrNVErPbFAys2cnTwfDQNteDDTnGhCfh0clHD3sBuiamaiShOWQC+bdhe3a
Y1OtMaLnec1U5okIGWb3xCKmj5edkWu0aSqm171NB/Agul5mylgbtdWWokcazW3y
tfIqOg9pGK1KA/0sLxqr42NcdK8fcEMLQAc3NguqUNg0lZQMXYycv/65c0PpuZ1X
0fjiKyukE+8Wbf6le0kWL27fAh1hMkm9lWdyeonkO5sybpiR2f+j8TmT/CAXFLVt
5sEYTOKyhTV2z1CJgRaVA5fyKzeebcT/m/+1wzIlqY15LrD5MmKgx6Cd7/PF8Z2C
D9IIJi+VGjjQLKKigdZsx1N6Ikd3Vw7AZ00ZJv5LrS3dGoDOn+JEPl3C6B3AXI6Z
pgMkoOAIRUKON5G/RQcwIyg65RbsZJyFigl6w6rLpouqsE4jTlg3+NQucogXdCvc
Snem4RgcWaNdbkLIDjoskzfuwFwShcrqjXv80E3Gk+1rC6xuBGo3Z/D9Fq6kcn0j
Yh+HCPHZUCsE11ZsV7GH4j+2e/VXVgKru3ibcOZhkXcaIros67aq48un7snT5csu
YOhY5T0AOqd0o/1Oyeq/fNN+avLwg9ekXuUw8L/hk3Crfn0qpmd5i4p/CeeO1lWw
6B+A4wR8ivSQKuW4+f0cdICZSG7g7U05W1KaC79L6kPq1L/AlU3BewJtH4SfSntv
BFrPiUzCBTZHvTs/Jy1FQ29+aWL5Y6gfOo6eq+CKEmXN3d/pE+HKdUIMe5/etcEF
IdioEMTWuCe9bVjxUqXcZnZzAMmT0b+io0gehbZV5lTH72ZHxNpj+ukh8F35y15H
cAwG6/5uyTKeVvz7uFdMP3ZoYywXnnAG8Oz4XoNiIG+nEJN40/VduA/zqql638Lv
t5pCzK1OHGEK9WKPl459WHIEctjjSQ1/nqEG+X9CaeXqvNL4R1DkD9LzwHAQ4046
4A1XvpqrDgcXursivm+cMp18sU+s3wNTHOaJg8pIvmbQ0KuOKXoMFNsWt76nmUv5
F1iZSOWcU/SUtm0lpapqkD/8kMJp5eG/p5ey4WkMhCcZRSyWJWUgj3rm7jnLa88J
bLBFMS51hrWvZfNCQDXt/2pZIFqiyEITeWBGyWsosGGJNIaE6GE3r3r7kk8KZNTm
UKeaMdAVisBuTpIwbrJNqtezSR9s7HJ8pZ6BiQCGYSsVGmCEfbz1IFXAMJN10fcH
4G/wa7uEUxcYayCErvWCOc3NQY1rzzkaeULj8I2e7iFRqne6EGyeAwVr3fxAlGIC
R1kcgidwTMLrQu5PRf9Vxb6Cla//17D4/VEh+/Y3nqDqZDcfbX7IkRm+0FWBUpI3
t7vWtvGc9SQE+kTcC9E3kuzyIhHf0Aa4egLbryT4UT3DIj+hbnV4WauO+DXsIBHq
/sht7J+EetIZI6zU5kAaUOAc0K7Mt/8P2J4KCX7kmUANojQbdEB3Ra1AFOEuN+ck
8rXtD+cOz3ArratpdahUf8pCxHP9FwQjYQXacj9nt7eDSlggxx0xUpLC2dz0WWSd
R0Ys4/Ek2MH7Hpgbn6UkItS2vYRyrK+IEZqo6gu/U98536c5l/yRoUH320ES2Q9F
8q3/DjPDvObVKwWqwpU55Zjkhq1sEhWCChxRyLgJZjoLWCBL4WbyRmx5yWjptgBP
cNuNwJPOz7Tf38q9jSxVDLGBrSHnGz5/1MFBNbRTh1uwDMRo83AzhLdg2SfKZjhT
p02H0gzI8yHYWCjMeDv/frB3ADWVKaIAgHOBxbMIedy2FIyIzSmJvJzpafakepBO
6pq5LNdR8OS40kPpgTZrnzCyU7dv6fD7Z2CpPEOjgVSIf7aRk2tLyeya3UsteB+l
9lymcWo3pSrnAbcYBAs5hZvxA2UOx8y7zz/8m4AOhsZDzPNQeQbZ0Cnf8eqI+1R6
DHTeaGZNFhNuD7z+GslbB+uoz5pnplObCS2e/ZKMN2st2H9Ut9HCn3Q/UUZbh87n
OtEBLqZRBvgHT/V6FlYMK72SshW8mDHycpaOugi14ltyfv7K7dhtbIudVdS0Cs/O
Q1BnG3nsfKK+0PZTNpp+kwvTbuSqYlayiB2Udk+V+X0J2nuJym4rrumAZf22cUEV
fA+MHr4QkR68lX1xprrOLvdb7JHX7MXhbIFqZopB4l99+UXrAoNSZEFGVjvhXP4h
q2jhEY18iIJ60j2cjbnZCtavX0dqSt/BEzNxUGdp4cfH0ZC9YIui45sJMYZQDS3j
UIz/QHTQZDz/osqi2nsUY35CNBi1oqB0sA6RbLOXMzZXUt06q/2CsjP3nQbSBflE
Z3QOggORrMPs4NCqu1TxXHvaeBgpdsG/9eBsnQx1nyZKpy4o/auDOp8q5Hjw/HE5
MyZ8fkKiGiYs331IsfPVbQqVkrvLrAkl75D6JhKyc+ilXr9+cwkKlKk7yBZXfJH/
rtXAAmPddQT5a9UeKl78/YjHWOJ+DPJckPFYOuwhLQsgydifaPxd8rvmCqr4NxjY
ZoxIN69I/Dlo8FibdRbFuApCZnHa7ywAj6Phl0C+Yba/oxpYRYJoZJaKvqlh7I70
KuTo5LUAywzUaluEtLvGoKnKeGcrRQvtQAM0F5ASfAp58TQ7o/g4cGPOEHQ8lNS+
DR5qLlnYrPGBAayU5nnYHgCNnz5oShtbl5aFc1WQU/bnAMb6iLFS6BhY7cf6aHvP
+aXWNIMt+nIpKEipkrJpWonrNaLDhbjXFs4EMpgJqHvlCfMG8isIJzJdwnL2NY77
IqhxfWY3k4F1FVegQ0SKzp5rBJmeO1EhG4Y6EdO2L+3aOksvMnAMnPJYE+tmzA1j
/lAsWLjs9p0eCTX+sdjqSTqMIe3VmoXOWPTdoYZ19Bw8H5TD0NNlsk4YO4TbEyuy
pPvdf2iaA+eUpZF9GaQfGHOUydAkuflRuFPonvSQ7CccigHiPM0xBBZL/t0rGQeV
sq5GsBfAcAwmUOxxwcxCnNpE8ueYlgB3gDhf9uXOtks/ahkNN4qscfvtD80tNiXo
PPBlA1BddMuRFT2RyT3J5lwNMzslCqnDcgExmhQGrf515vCI70L118RWLAJNSt9s
wMbbGqhO5wUVlfbDzey6oMlEwkNi7rE2ZRUhktBIhpEkRlKvkpqN/OFBuXHbV7Wx
VxuiiwwDZ4Rbt/xQ6ddiZ29pxOjme55bMWQwbXRO6cIqV8QBY7heHp91wDFNKeq2
SnIdO1zNbhw/pQV1VX8xKDqpkXwo5XxOWR5+h0sCdAk5HYkbruix833X2rahBJq6
a9x0oFR3iSw+tNBwIbxHAxImUM+MnbZsSI/Em/TUv9ZrXnD1lAcQ7TIi4dmT3rg/
y10LtmDvbg1TN89xxESihq9Xb5GNYEUWQyVtBBi3j2O1icr5MUJxTfPtosImV0uB
Qy20esgvsawuMFU/HDvB/U8xSh7H8+pesQ8mMaXpxnu796FXdpUHECePKh6I8nG5
lWwq6f5oZWXsxAzUmHHkEt/57QxSJj2+mgWDobpV8FUi5kDIxBMbrFtovcD3Zzij
I01gZlR7YlqWkstNGhxKPCYKVrEesLbQWcT1a/E1aHt4rmi8i9yDwGiwYBTG5Yku
hhnk1BxzK33R5TEEZgzz3KqxMQGAAFOop3j9wiEA/bKXNuAm1r78pAOkCTpYox4/
+UpFPFLUwHw6N9yhpBso7W2NslgikIUH5zodsCk3QF+YeQzOi67cwZnAxWg7rlla
x0Xal0tcZ9sT2LY46RgGCoqdpl/5w3hCxq6WyOQiuHGyWp93NKqFKURo3Map25xx
jw5hkriKIp8jv/sA/4vv9rKQG4IfXiOB7riiryYg8j71Wk1PdrCPPyLr2Np4/G6w
cGSUc3trPpyhvBS5O2gFMQ5JmrGqiHxiAbJGs2glr6G0hUo/3enHZ09FSGpzpe2d
MWmBVDQEzOOxpnRAwo0II35SuBsgFwC7SwueDfZ3U+5mh8AalTk6SWHKpLtuD6UR
ux0NDiJ8IhXkCBv5xpcFoY4QQKMzvBBQQ7SfQaf38fMMXMnNOwXvPNeAGXG3gPfC
2ZrO7lN584r3hynwQUOLXXzlHXGlN60Fak0KOtrB5HLZxL+I1TxYtavfcpJamMJ8
M2WxHwXKSMO9mfRDjnPEO3f59Qk6Ox2m9F/Ph7SFRfAfTRUFlNjc6vNg5z504Gif
iUluZs9FohJmRfLm8pVIB2YVZjoCL3Ei12s0DuGnV2LSh75RBW/jP/TkuQ4oYy6u
JcdJlXENFyscPLzHc1JpynZGLh7ZsuXAyWZi1g5/g6hpSoKgmNyWLUSjgJl7D8pR
QJK9qR3o18gi63lQ9NAViiLvRVwhS2LYqGrWxVuMWAuOaw6TKjLXZhXiZY6dgg3s
CXYKLBt3DG9BcuYf6W79Me3U9/Y4+yMxSdtShMtcDEVrfBYjErh/TfH+PjqfIAR+
kdRMYteEBoGwP9cj+a3jQXkxZuQlZF8tg2uYNm5HxTFcFMmyN2WuHmmybmbVQGRt
kQcQT6CDu9cyk6hGLZKU0R4AecwuFBwx7bP9ELu6vbvDO82wTC3w0jokIUmOFARA
vVVVXpE9+B4hMwzTNLPF3WRT7aph7ZqWke1SR0z2YU+MSCc0LW8N+jw1dlaHQwT7
lk1iCdN4tyNxR1B4WnxZlXTTmm5yDLXJ5zhggw3zox6IwxT2qaUaKE7w57uZ3I7G
iiD4zLVQW2KdJaGhMOaZ0b3nhnMBEJ4QpIqEZSlJeGvyA5rbtU6dcwo2smXBHhtb
CmMOWNDhqwZe4FdpysfPl9rOVgxgpKOV4LoEhqViDlvRD/veT9bOyTG5L+Pa+pqW
kKKlrvWupR72IWUPu0TN/volNtgapYVRE9OT8+/hHXx5RjUyAGEWxybVSRmL+TpI
Ebjd7KZdyMXOSyHKxo1a+udgzm9gWhlfMmwcJayIprflUGscNlGoeZFVnIWbRwPu
HFCYkOhtixGf4lu3/Q0KPTrM6SKeyA0nMWlrKDhvoss/z0iFpxExEOIShTIvOKIE
a8/zOBPv3UcLx6tI7pYS1yyTqTwe/nbUZLftZ03ka5OCELF/fu49Q1oZsjqfVItN
wjidUibqabcIXo1ec7eoZaspeZES3ODlpMGc6NBXbOQvZNcCT6UxPiGTdDhCMj++
RinicKZzqbbIjgyQcYc26yod5eBZEkPF54/SUKhNqNhior8K0Jb4Lm3SuJv8VQfP
AOVnIbI41kMAydWUWWyHpr2Zj5LfoO5MSoz7MFvquTMVDo3zUj9qYjQNlH2Qy1ea
MiOFCAej5eZo374QIL2FljVRFsEPQXguqRXYttrlcdC9pDnCPbsJQ3VhuPXC5sdh
TaS7MtOdmdxiAhJAnweS62z5kMumvXXXy8XkbP82M904A0cN5IfwXbfcvaaOZPKd
Pn1d54b2NI+yWcYOPJxW/eBFnwi3zyWYxBhWnldPbHQ24fQzO9A7DmxcdRAHiDF4
S2m7AT7gVDHRkMv2IX1YV+unTmc9cf+7Zutiz7RvWspRc9R9PhLGlvG7PZQKNW8V
SqRiQUzcP6LxUbvdcWKLwHCZfbdepZJcxSbChdZEkTCzF+5SLuNsoYZogdFyFHVa
bBanIibD6/weyq2li3hu/w1ElAqbv6xqYQf7b+7n5MehxjsBMho5P49lW1CXIsNy
Tngv8M8XBnEFSG7HjoCV1vBxGxfjlDw5qJRgYdjsKPyltGFriZJ7MwOwii2pOkt0
E3Gmmn1BQJ/V4B5j1tmqDHQ2cr/Sdd+XJAMR3sIjAQL+lIViGDhzlX1frbKFjHeH
8DvAIcP9mtPgd7tJyoq7o7l56wW1cFX/vXHQcyqbfuu8QwedTO/3Sql4MmOCWC+x
BE5MXYx42bIOqt/p6bkGVAQ/QU8Iu3xzoxulDLPwzCbhmRkntm1/eiQ/Fj2d3oLH
86mOpPX/EBB1dT60VOX6W+ZXrL/6M94CCQM75KiK89AEvOnoPGM6QR1QNcvAMJFx
hpYKhV4Asousa6bxzaBaJc1i//Fi+p9nks0uRLqdUwwQ+Mxft6XZZeKJys+kUN4I
v7QRheWOsLpQrs/045e+fU/Bw8LQfpkP+79GB4Y8t+2Uz9qcxwHH4Q40JGlGCoZJ
PXPCvIdCgdl5xVAUUecvCwISXhRY7FVuloXNdvtUMLFFLYiwE0O20Z6sZwmocZsA
q/5kFO5xxIXCwmzfUsf8oWkV9x7Jy7oK+8lEkRsRZaBVY4wzpKK/1EtgHHBzIm//
fRmu+v8aeI4D4JTo9+4h0PpgIpnISvJ1JgdiUoJLh/P9QDMEP2hPNtGpEUlwvAXF
erX8QUWpOSVPUAC/pLr4O7BC02LOx0/bF9Uf9tVvoKSQZqFOVP0uQuIp98ci7eVG
MixweB3fueQoY1JACThZndS5QP3d3A7zCU1QrVl0Tk6Iru8xelI9AQxfOy9r4hL6
bJZlvaepTlJKsyaPyb6Zq/TqB8cdZKLs8h4J7etc9MzswvfVmIug+MFkLcxETVQM
xPf7YZQ0DdIp/mC3FlzXhFdkkKvdDo74fNqr0tFcfHor26d60lEuBLzMJpxC1vS2
ZMBQy9I3KUzb0vguqqWlEN9f0R5C6rMx7P/9MllYMqzC9jX5KQIUeVJgsZ/ORO+E
PMNodbF0m9cFSslhkXHy7D2rt0LZvVMfJQylW5r/Jr0fquJei3W5ZrgKtIxR5fdi
45TI+/HD1GGKeJLtGsOrQip4gOo6L0bHImB7FQShh7RJQHWT/qsjK/wDErAbX+kj
sirmx7hTLj3fOSYb+ZPRS7HwyYBTbSCEvo4zCQ338DINPcwSc+twbPIn4mT71H02
4kniblf0kHJwANVpTsDzSnGLQFMht6bkV2I0FuNXHHiJ4oFRN6YcUvHYZitAhfxj
Cr0puOUUpwTcNGIJb1dUycER8Rzc3mrRJ4hH1i2u++I69vyt+yRHR5BBfAYakYUm
3Gv6InWvbR6hH+KMqOnsQCboJMUGm5ifQIxEVI+3ZLFkdx/rbTz5mdndW6R41Fdj
P/toVCTLBdqCrWSnRCj1sa3zDE2i+SrdcyiaMV0SawxaHvQcK35dRylGzRj0sGm3
bKQJ7ALcF2/FMmP2QU+OgXwO1WA1W7DUH0RJ0EZdNFldBuSnR5LfhVX6v/SDmQoG
Cq2E8Ynq+sUk5iyQZzWdOxv+YKou49CRzQ0U/j9dRQGZajq8XOhpTYDhh4U3Gz03
08x0RiCBl2IXmm6bSdamV/7e1voZCzn0TkcG3dbhRh6ueEXnsPq3w0ClcKcNCCnn
7LklPVM9nZ4dHtEMhdzHSBUpVhBjHoMI25dYduEwkoq+Cu3l/qXPNYkBvVFrU5D7
fT01PHZkxeRY/qU+wkBD8cq2a0B4fqYjbkqR1yb3tg9AhUqTfSoDCQry4+3DuWxu
9YqAnoR6IDrfxyj+wwrC9E1SYKCyBUv6Hj64S8IKRPWJrLYocmrWOrESyvRX9iqS
BbVBQL0mPt4xo2aauW50P1ro5MnYAw+qkCxE9DJ2L0PS7u94u7p/sZciUFQ4tKV6
zd2Mwhq4XoDJmH9pPU6jdy73i0g6PM73slTHzYCb89rNAeusa27xV/ZKtWvt3iUh
xQZ4AwcBfIB3cf3GAlnUUAI2Jkueqqxk+ugVHCzFSq+mEC9X0GMEezwWE4gEnm7P
VcUfNHm+EabGCeAHoj0Ui2PJe6DGBxdQgNBuQVa3e/wb1FtO5K6wjQHtJB3/gsQb
m+NynmEYclmQJkDyH0dReLS8tbmkjqGc3DxbflrJHxt9C2OlKHicz6zEf/JbTZym
2Xklc/WniT9p+07aWydG9amTpu+3CtN+kW6VHevyTyxN2Fz83pCwqmFDuEa/DB/1
LFnAaPpZV2Om2JnS48t7VnDdRa0bCyq/gSpwkPU5modYqxH0AzcwshI6DGaYL1uW
ak/iBXaMXs5LdTUKnI3oknSQ1WQgHSwTEBZ4OVZObEQDNd4fLtW0QNuCdeNGJQ7l
Pcx36qEPKhWN6ZW5FvBdMFxD0cMUIi2lYHR6T3xIMGJWMgmJVHkwe/OH2QiJ59uR
/yJUJVIY5fXcxBruB1v/jjOnTXt1igiAQ5J2MBnrj+caSAG0fMpDCjsBU8ytFDG7
1aML9ir6GNhHUCuSzWXd5/WTg9CiQU53TskFF7Yu/TwmkY5btQb6dMPuU8UtuIyt
mdqUkgGPW2y1MB0YYrI17dHgpYZ51ETjQ2YqXUXB5IajVvI3r8Sg2qvYoG4OTxod
t4+nUIMzmiQrw3x1AU0ElXIL93rRcWK1ZoFzlfzzQ7XjBt01JR6Yx1hhsv38P4I3
zCrjay6oyTkj8xQ/+XKPTGLwvn3FIKiSB/UE/KJmVoNvgkFYwgHjz8pHZNCBMb7e
5fixrBCtAkEQKpdt86I9pIHlMnZ7+mTk7RJEa+GgZ4n+betWnco7oTcC09KL90Mf
ApjDJ/c+8EcsD3S+GDZTbzPGy0fmwqmPGss5soVbxQvB1s7Jv16EHbWyfZXjPMor
thnict+xWIkTlu+26fTPvSxkaAQxfGremH+BzNn8MUmteAPBCq+fXVILPgyzTCwr
jDOwfrZJXq1Ov6+lsQXC4N8yJLsSEolFaGIHy/sSrvumUiw8xDCJT/t2K6MTggMX
XHkD0MNV65wfNGf7mMKbKPX1xom6K5Bk5gMHMxJYl8nrL0RRAcwy0nku1ByUM1rQ
U/uhv7wK6Pz710fpy4eZVo3Tdsq5R3aEP3/6pdm406nckmz2UU+v7C404ix2Ggk2
SQDYf5coa50tfg6+/MHRa61eX+7YgL09vBmy4fdtMfvsL+Y4mSIJpjTrW/XBskKM
NGx1aV8MNryhv8GvBNGSs9GTTADLp9pazA7oG9oCMqJuj790TmrvSHrL4D80Ty3J
8fs8PhguzPkmG8XpC+1hBlaaWnY1adEcflkco7hzvb+4dzpYNJgjLxGIYHU16oh6
Co3qChhq6qqQ/ipxDYgMktOj7pG8w3EFOYxfm/xt/5eNIV87nvNzaf5gwb1diTbp
rb5JsncIWezp/vgYePGUDRk7AK/m1XHKfxjapTvGbpUimPnVCqUEY0OtrQdgBNn3
/qu6qSr8b+euxmeIxqY6Zp+h9by+cV8FZEVNGVdQZzUiZPT/1CG6qnXHm3HV0azA
9lDMlFGF0KQ6sJ4PzyiVTBceRx48uhq4nD4DQdNmSYN6fpAdTMhskdRncNbKrQyI
1Dyq6G8S2ZoAZn7trfiigInSo8RsB2KyGBMCv4jaA14TYM+EZg3FJMF6shvYUXJ3
6Bi6a59CYhRgOQpJZrKF8nM1yP8XoJsc8Vqi32AEjT4ZmWOEB5mpBwxTBi0ii1Fl
FFz+XNZEKjrsSWsZMv+hfXzyXPpIqihGLZ+hB5EeJvSBynBV8pvQNKsWRk1TtQMu
kngXGggek6hm01NHq99T8wfjjKTcYL0JvkwKEH9oLrz5Ib1pq/4WCyFdpOeyxEBT
mvl58RetmiAbCCl57uZRBPS874SnhX7rA0tsMxqRwrRCjlsoY+jIQ1g1boycVsEu
IoDnlq2lLlAsWrQ3qieeFgPhOuUTv/ArQq/yDVDFOo4XrmfbM8UJV6NeH/IdIdYF
0zvbEdEVjftxCLMfy/RSa+blHkyhF9ZHJpb7vBisKqRK9EUoiUtSMdrvYmPJp7La
H5T6WoJ5ueow8MYiS7CqktlFK9NWYscg0bXXTCebQAuORDRuFFNXp1t7z5a0FhwZ
ukcLHbLHC1PEaN1nV/+SDOKLmqFAx2K5nE8tSbGiaqURvqQEcu4ZLp7DEdonz+Ul
pIfLsAwG7O0c6qlSY1szGW9Z0XfwTSA3zZmVSkO2wgyHhoR1ZJQfcJUMZIKvvqkG
f72I4WA1/h0BKyOYfNhQ1vP1yOOzWQhQUN4cUOWWjy3h9CxFfQoHlFvP2pBx+cUm
QPdcZXU3syDHriO2yCTytLtnqH7oNuM2WUIM1cBHxaIM85xJ3G46JgxBALsoFahd
bjW0IpmYV/+o2LczOTh8fax6kSGHJPBIIDoiQFkH0ML8aQgg9yq+JhZRuvAEdKj0
x+tmWCbw5N0OpW7GHF7J711HUMvY6wbS3nM0LzBxlOfYvbyaY0BNqjBGy4pioWFY
ZTvF6BBXFyMkjRWf3FD4HlphRLHGoeQ+cRpVPdkr9XsMfN8NmBbN+BbUaHMqeK2B
zeZrL2FjAHu/RETrGA/tPLeN8G1S+vRST6SIEdJGQbhJYc4OQIlAnY3VdohPGMnl
3ZyEB3y6sv7xQNMiGXkxzFnZERLIpFtEXV80Ofj89qlN+zlh5sgD/uy6uWHeucZl
zHT203Cw/owgWl5da5t7EitXKPwthm2zdqUyOcN8twlu/6s32hexueBNo40HkK41
rbIsbdCQv/9EwcnU4wTCLEGLI9mVv9x9u2tzvlBK+I8IBlUFME/4WIl6twOurd8V
vdfYueNDjH7IFGn/dWpI952fRkPhI439jQE4n0UhqNuSkt0lQID3ymxb9GC+fbHn
lY86ZBAyFjtFoOsjDa/3xDu5N+gxYdpZ8RJGvtgDEjs2LPMhCs48hpijP+3qnU8L
QJs/m6c6I/X/30TQJovzBg1eleDaUkM1dFlvV19b8o8V1He/DWck1vd0Ih8ZG3/S
UEOmI9V8eERE8+oqSaqGMBjhALbGeh0nF7haIO++nQ0Xs7ihMumTh4k/4AqgJhOs
WKZbZoeGJTuMUiws/OHlnYM37S6unLB4wwxGnzez2+cUjvjcPhyW4ujL/8BLhOtN
OZIzfvtUfLvEH5xHcel0O6NGRD9wHpZpfiTWSfK7xYBGnR8O7fPTG8etL87JeOiS
hrt8Q07Xv0LfiijoJhqDiJnlHFKKJ8TV5iDnuQKJGcy9MNxS0y5UzI0R18B3a4jS
eIhRYRF/jVQeOygGE9gsPe8X+NHvxrQiP3oQzjF5+y4+EnhGCmZlHbxBcznS3miR
rHoQxYyJqBGfDji4jDHA7MV1isuBwuVAZMo2qnk6zomPt1Q0YFcp5d1tS1ApGc6Z
SlCKP20TgetT6msIuZzUVQ/1wuA7fLQAUnGdTlsCtR+7fYZLQwMUmtojsc7kvUPx
deCIc/LvbKnjqmUgJVD2/XRMp38DOH93IMH9jjwpchStuJdmTDbv6plXMHnAvZwK
Vnc7jCS84thDZBZTNDJv3SqOtss9KN7YOlWZAWFoE6ZfBCFQC4C70coifPXiPOfr
xbX+1sBGJR+IaeO80L6XhSQs2apyz+xPaIG8Xq2HnEQTCxqrT/bGYAlUnqPjhnna
SDf3aLM/9qCXAWVMRc3zKgmogtLOUPknBsbZ9oMfGc8B2isNzAriauLZg+fYZlh/
Sm1TC87YOKGYEB8KGv5Fp+jUhnyDZEhdxB3Ac6aNhBozgMTUk9Pz3IVtX+R9mOc8
OETM7+KFEx17+53MPWW7nHC0xk1dpYFcMuKxjFtzbyT/rkNGthZurgwCuFYOJ3ts
i73NU+aMvQa5BW5LFA2oTNgMHUFWXXd6KYA3v9SCToaAh5HmtKl+9pcfaohWoHy8
ydWDJmrfXJada9XUimEeQQisfU5WHxlGGih83MmIQa8KfvoaGuJ9Ze0lMBNI8e8W
+/LjYbkdUhRNG6GO7UDuczVofZcQQt4SGbZh78mp3Pwluz8knR8jivGSIuKrIN+f
UHhP/0Ri4duKPjlIZ41p+mBY2BUBnAqKMTyciYeCRbwiPxchWWnjuaIstI+1QBvt
OPoKzemW1vFese34v9KRWI6bjAA2TrJ6K3kegmaeyMyf4haXxSTT7rSF9Nl+ywMY
cd52S7C2hv9wcv1uEoZDOMymYixB6kap5aG3thRDfmCnctvuQi0B6Ga13iuqYeCk
Qo8912DhH7uET/ZragEC6rIUkFaRlb6olkHJArCfpp3GmgNeC31e0Hjl2HDesppw
HAG2/58avRlCxJDKWN+Gjp4LcybLIZ8sPmppMsHgC+xW2DOcYtJYUQQB0BQ4UoFO
uSEkNPEf1Usord0Q6hqgDHxkktUq0AWoVJxE3UmoBo3O2PnZ00gEy2Qcvh0M82o0
lTBkUOsR+KOjOAtCZagO7h2wSLrbSMMj337fg6mj7DhnceYKCVbNVnVlZA/p7epc
Fw7uX0229pZGHCocYjles2cJMXAyJTyq+DsA4pD+3dt2d9Xh1JC/a4/IxCtJ9ETi
iIcIpUOlNWpScCMuUSx56vL6rEPqru19sRkeuDw6Tki/7DtoWXX/bBlPnM8h0Gr2
C/U6vukGn87ZyeYxNX180e+iHPFwGxWebPdRqamhmJM9nO32i6Y0TVpCiEJydLEJ
RfG0VW6gzkW3/3YgYYPLYVqw2JURtBRrB6mAM3GUFHRfmcRiMbgCDqVOCLVpLN8z
gSXlX1YPImRqQwxDFMgdLNt/J96njcaBTmp/qLtoyb5TQsdhXsjxczK+THTYy3L9
lLVZ7sVKxNvc36grU0CB6ZpIVefBltxXUNu2ftWN4ELAsl8M5EvsnIjfgB9WDauM
FTvw9eQQHS4QvfGg3F8wpXrQaWoLPVxp7A3pIZWdTYhrbTuJimu49ctx1mKfYndt
pLr4d2bqQ/WSlsttaARToetKeX9fZDLEX9mmBm+yqZDmRV+mg1ION6kFT+GHVIDl
kB5a+SF6TDcgf3lcKiot89dAjr0jLYb+K+waArabv17QSokTtyFSdQvPYi2pqmZG
ajxh0ZJUG0ABLPO3q0PVRlV3idFrADFKH7kPydW7g/rOtIQocQpxc3cA0JlOaQxN
SkhaXVN09X7jKu9mQkrXrRJNgNwNNm6KUnCLgZJgpoduo5B1qNfMTxfZYNUkSBXB
pNFH5w4oEL4Czr1a9QIy0SPvZede4bQ9SONQWYsk4BXQKlpNJMGefagpr85Le/Me
n3ut2URNPMc5emPcil04P9Jfalh93mJ+Fo8aRBllU4wZfgKDQtPsCgsKM9tUbxxC
UFDpkyX5v2E1pfgXNgZellV640xE2vL9guY1SAeiYSb9lpYuN6X16VoDnN1MDM1+
XTFQiqR7vRXSjiLeunNeiKv62vfnsrbNjmqTJVyPkDMkVrfxUe5GLgPBa8u3y9j/
Wdyoi5LQ49dIRGbe4JZc1BIA4SkaySrG/wQ/ylfrqKBMUAj70ZwzUBq1Mb4a620H
597t4aulKzPtOVoBa9W78HlFbdFhBMEssEqN6iAUGdXc/6BWzgc/o91CWqsqKiJZ
aiyQh8Ykmd2W7L3BJpl8yl5AWcbSjfsVuqM2KXrtPLRPFTmmfH3FheVfg9UuQOTR
X2Xf6MI3GVAEPbcjAKrhg3GnBbp64CDXf4n/Bv9nZffWMosO57KD3+Elqz3l4JzX
v+xa+RqAOb9LKtMvAJaDqjnVEIa9juKEcllgtMcwzoG8ucSmgxyAayDMRgYCRvrc
JKNAeMRsnSGgEvRDZdDzrXSnjsPuhn58kLtaO3fX/QIHm1DMIkdfOb4o5ui+xvFN
/BdAHj96Yz0eBhYvPPvaTIhcrAqMLXoplvnQ87ZpzcnVv5ehM7qLTBA1BUbW2ccw
/Cqp5DRzsfce3ytLa4pkoeJQhBcD86LIFEN48MzNoUELABms0fd7TSWvga0ABmpd
Ckv+jlqxGpvuNpEyBi/b4/Mkii8fe7ofi3aqAOIcXqIFOsI/ilfurI9Nvn4lzPRs
aKLAEC5WzauZJhwKNhmgWgMyFojrAmxGfWj7427p1uRSEURpbJGH23kQo15E9Zqu
u8iWF+wFaRy5R1RuxdIyqS2qN22Ci307RWMwbCBS/SV/OZN++R486cP6o+qC1sRj
Q0l3Q29IOvauAjOQtxLSAisf7dA54kEwkPl+JTalE0C7i3r0CYHOWYQXPL+Kq0Dp
MrB0+sS/3sb7dAZ2ICP0PG5dxPIelDNOWnQ1c2DBLl59LWBfytxPSkIcISy9Kvxt
ziMcncWUuBYPafLREiAgM8bgVImihyV3uqfWa/e4vv7F/aqQUoVUIl0GCaPGVDi3
dJp1V1zYpSWfM5kac41CQKoA8NGAd/F/KcGrCeHcJq3xY9YXAk0LqSIlS8SpFud0
4k0pOgKSzjz+G9V6ST9kNWwrlhB4BXST5v2VjWoOOeISBaysmc0KIIh7FIbfP2bk
AcpV/PE0RZvgjhd2I7gHCN9Yx+EKxiVWXho/zi36ELHpirwD2L4pr6JYhzj8ETZM
7BhMTalgKwtqsjwFm68tDcM/aIfbLdYXFmMcu9NUeE4XrBcS/nblGS0lb2l3Q7in
3z36iRylNuFa2YvABBipK22NJLhkCD2r6NMrOiTgwblCprGIMbxxd483IRce8LBg
vnwitcssOO5S/z52XFjtg6piJa5MydaST/bQPoLLB2fRy4r28K1nmIMAUSHCUkNo
1h2X0J0oqgUbJx0rvflLV2j5mIxbOfXokrlNYnufk7SLDLilKkI5TsHJbPocvwPL
tHPs3zD8QviHIiKGDQ3hLHV65LfwfaJEKLO/iz9YNAXFb2GSa9Z1kWtJDAE3JThA
nnhTFeWselUZDOEYok0O/GhLCaYk95W93ghxrA2AiYifMvf6mpmOBDgd7k1D4qpO
Osjx0b8ro7sP1HwWbBFTYxvRTyFa6nLWnPLHg8n865ETsb8qyGPuQKRoWXWASZt3
MgSF2mrqa0EgR4A6MGMOm1z33xObgVzH4iL6jHHKQ72VB6YmIQqHajLYkmE2uZzN
/CRGoO0CZGYcizu0QJRgfwWz+R3tG3ahzrRoYwIlmY9nOhdwG8n38eiekcd87ZQa
wGe+E7a3sLUZG8nhhBTF8KsAdVRM0LBur0uxc92vQLCwZ5Fk05USk2DFOeqxWG2N
GE+6rnFQJZ18JdSyuCG0xFilX7OKtNDARBMxoFjoWkJ/CUjk0SntTxIOZV4EUPC0
f11HxTXZ7H4oyecUq+pj7nwp3KaZe7e26MbS6vmkbgyq5naG2EFaZntLaliGjOjo
carnkKnpup86w24mxppK50lsM9XewsUllAqeR7gD2Cga7+4Gubj2nEodDEbGOPNO
PIlyQ8wPaVCniQjkurvoeAXsHwBKZEJEwTwUR9vEMkM1SB0XjrR4Wk0ufdLH32JJ
WJrk3WZV1S500A14azx1vF58wpsGm5K0OjaxbuokFJ6qyJTlp18Btp8MWQjshNfC
RRCHjfKq9hlphkd2YiVXrTSdx5neyvqD+NTSJQs/yMMTgcwsfGjg2x4qoxIvbAPP
k5JWGusxQcZO9jjYSkr/xRfFgybJOrvVWZB5yUHoYbBazHKrBthnUcN+6LV3zVSa
BOb2Wkl3G8d4D3iRAbqv8Ns9tJN57DaD/vrErFyuoC8GYgmSoYPyji5o2R1ASlap
Wd45YE9vFH8GQRA0mhuyRZiXnGoFu4SUX3iiNkJabQvK264CHw2wsrLvnUJI5RMt
24+mjqTjDPg3H8e/4K7QtXe0VV6+KOJkW4ehskooNIPorfoZcp8gfwG64tGfsKMv
TduoTP1bPQYyLFCjKGGdc/aqoz1K4oiOAIErezTm2c2hW2o2zY+dgKoPTSZIWTmZ
7wAE5BA6RytLANzZC9Tp3yLHAnQQLuR4zWZEMHGgufJc/4RRLMdTUdS4m08ICf3k
WX3DvgU8GFuBTPFghCvwWCxabQRve04tPrPQMRiBJo4Z2vtr5bB/v5UKlg8U2pnf
y/NDNNQLJ51kOyrLPNCbx4lkYBkFU3+fhO16km93lWI49aRXHUeMWDE/oVKYNCHp
gL8hnH7ex5FVAETegm6GPo8G3mSUdshFzDHx301KrLcKCqYnFwCH/EEAfhhxQ+xQ
gI14gitgEGbp9dfC2lTwN/MZa05wfjSnkl3acGIg5wIAKHHjRCbM2JzoeWJ6sexz
kvbc6CxnxaExTVcctbYRSWO0y9Nd+3N5V+wllcbI24rAskVM49mlghcQCAmBF8Um
DuR1/gJUxck323gqhA3jm8Nf9Cx4yTkojVlj/yxqVSulYuPtDD7eEuadeV/h8Sda
4Iei0wbMI6HX1Bc718mIcMimxuPZNFMQfhoKguLM4oS/FJrxlwGj8VY31L9Ff93T
xEmHMj2J4wGECgDYA++oTWSTktHCccog4b/rkTDDu5mYjNDQbNv3EuDRGKuJkeWN
JT7Izzy0bJCeJOtqCoXlb8TNE4EE3NNa+7v9PKj30GvaHvsYpTgHbghCDVqcCzLC
K/PoYFN6hcwLYHUzQPwXhpKd/v6lOS8SaKK+7ggIPNKDI/v5cl85GuRNkN4rxFb4
ttyEaOB04dWv+3tbsIhUAAQVeKjJl81zbUQWYcqrXjOeaRIRIOE8g7g8R0mxDPM2
BidpJlC7GMAh5Z73sSwxkJkMnbXnsblXv4XFONDLjdsUgCwPlYiehpzLAMhKSLFM
FaGgkQz2uT1SFAesLounf8gU0ihvbymUghYskYL+t4HLOAb4KQnIUyYkY8jbwgCy
FOyCUOxOZFV2zCfmFMVX6E3TWDa7ldwtaO3sPcaf+BUSuGUh8HVjrlR+YW8Dqooo
2mer7wBTowJDiZENqTO2ex78/pkwuoQMxIwrJIpEEB1ukgM03/kZmpRmGB4ohhB+
y0OpBkkNvzqB6QeRjvvHS1pvTbYtAHSkPOXwDy80HQ4bBqdVnPX2ol+TCFRDK8Se
GPQH8l9IghJv5p8I3J3o7UIgvH5t5ladJY8kdCqizJ7qUMvQ3+xR6AK0nRWS80PJ
BgUcJcSafsVzPplgvsVbzI1ycT8Aukkwd6uiMsPzICcANZDOHzf0A4b7nAbZt2Jd
iNNOTWkB7QZLBMblJ10gO/loZkSoxKgSdFvpXB/dyNjf+BC/aRobtKtG+zEc9WuW
awHTU1wWUYQ4piqvE9HtZE06TqQNH6xvgVhyW3AC75gv/hFXJyr65ilLpvRMs956
E5+WtAa0GtEGTcnAi6Ll8MER5mDNFt1TNhccLBTrJ2gET2q85dTE/Ld+XM1nSHK/
YP606T9yPIFxcak2HWSroi1zcq1mfmCZ3jLNVIH9yMkc6wnBnDWIh+8ZRecG/FlY
9jr8WN5wfgTnobZIufEhI0I9f42pxO3lqScrIWElncl39iTq5Tyq47VKgXhC3ZEv
/xQDWaPQxQqyFT8R7/5ktxcEocX2RycKuqWwjdg81hGusFbMf7QrkqesqlIlInyW
3C6SWIA9wlvloQXGxkfRBQTWFR/+vPVBSC8WmWw0HVBvAamnR4vdbiHjkSsP5Hsk
hxerNkg3A6jKg9XgFSfqqOoSV3YgBRTh5kaTz07kIiGzrpvYKloJatMjqJJP1xSx
j0r6ZxZysd/sKEpedA+6vW1uG9j7XgdIng9wmsFAnhUKI+udskMEMc1m1QCuaEbs
NtriXVijXq8VqRsADY2LFH4P1ivijouuexx2jl7t6secwZ2tnUfi6LeEjBCNPAgO
dfsbYOiKcIQKDGCmFmFnOVDuHyCpe0m15egJaTyPIkWPt1fyGmhdTsCkV7ivxy+/
Z0QeSnd5K3uFllhmVsK6XfPrih4zPEjaOJfZ93T5UCbzx9b3Gh/G9fos2LKDvJeH
gYx2ScVNmUuqEG8+n8YkqcwxxMcl8eGdee4ADsyzaU6gadnxxIHHZFnbAtbtCf0A
C6Kfe83JJHv/D3GfPyzB1cMR3b3RyyDsyaKidGJp2YrCwEhT+ajmrCKnbCyr4cDd
WnRy+KR60Z7DxKifgVBtgaeZp6nC+G67suADqKQUjHyqDADYpuTYLYrzwC0PNKkF
mLV3lERIZ0paRaymsR9VVPRczesjVAp8hzRAq7Pflyogb69naP7acEK59HGI6CWT
5/V7qlXlD/1vTjdMi2BCI8gXN7elch2BF5UVP3SW+I2sokebgDa5Omrsk1wnBjlo
ex1XvRMA/YIaa77Mu190ctrDKCpR/Jt8yYu+dGyYU511LUezo8Zx9Tcec8r9UBMT
tjOngzadMI42bgWeNHzA4/AAJjz18OxFsV8fqBHmR0f6MxZpUE1iyvpgVj8NXqDf
tIKwojWSUOPI4MxGA75EhazqnSNgKvvlTFECUPffgFKEbq6fGDduep3U07ClWAOn
HVuvHCcFm87v24PpcFFff4aA1KZnrmiZElegkfCfgHGquiHq+M+RI395t2tWSy9q
C9Xmb/pjR7gPsgvlagpKqLbmMdidNuxDCFkQEco0Z3Rf45DjBHZfiBww4MkLYa1r
KNVofkCKyzhrVCOAgqwTpLcRpbL/NcvqP5FG2awosLnPJiUjJYUGEhfyxwwHFLg8
Jk1837zQjHG7FwebEk9RxHa3CmxnIREI+RP/CpXP7sktVNGYH1KKPA+s/AVoGjvq
V1lRI+NnNuJe+kiGxmTLFteRxLA91WmsRTPf8vr1R+Oq+dVJhLfq3lihIMningd7
UWiNh8rC1kgZaKhjzlxlsYgfQaxaJXUJELiinmicPPBmJuxSbmc4sL0QeKMbeL/O
EueXNFkonw7YEAaXiiK21cIjhoc8hTKlA6wn68g2TE1F8Wiq28fztEwAU8d7SrkC
oPQZ/3YogyfJEDDbHWVNRcClWsWvaBQGzo2GqjliZo9wCx94PV76jfSpxWQA8fRb
j5KyUaKuZOhM0yFPA9v0wztNdfBOb2oxGBvq/+tjfgW8WTTbngT5sgP09M8MmYDj
SPZJQj1k74WXaRR2abJqYYfFdRCKepPlaZtraqI9LmE3rM1qfvKqrm0ydZbgbJSd
KMWVYn9VfQm9vrKWHvNANfz5dgqQQzbz0CF4uex7y3Hw7lMbjEi7I65dG8FPjGum
YBaUh72hgCDD2NoYE4nRgYlE/ssEAkzxnS2kyzx0ocrov4VDbkuF0C7BehBeQYx7
AiV9HYsBxyqlhOp+ihN7Oge83zr5NZVkb8d9KMzZvUem7TPZgiuvXHRDaMdJ6cTR
nuzYo3QBJCQmREJpBePshIJ+3ihSlyGh+0wpB9Y8K48JBDwIzypKJzOCAk0iW9k0
ghW9sVOfKRuLyAxILXN7477W4tLHzuex9eOpXFDPHXYEnysmBYUEV4mGOt/6nZZ4
/9AwN0zdjaqD7Vvg2+tjv/SsW+4wJV5ISzzGUn3TxFzrpzAnqEuio0m+bpNew9Or
2zvxeTtSKWYtqnpCQUyS18xN7bGob1FsWnaZlS0us9x4RI2bioegbThXc1AuOWNF
i6vaTKbcNG5djnYEV5PBng/lOucu4W1SNYOOVXAIT7mbrDht//FOZkPGapQGzKh6
5+hRAulGvbY6gu85b8umovd8x9Z/9iv713A9amKaN/lOGSlViX5FSaojXhUE3j+Y
L5M7tOBTB9lCDQsFPkBKfCCObDrJWVMqct24Jtg9530tmd0iZQojjvOguJEdr2RM
/naMCGtTc+jjeCUjiH1P0BivP5TIgGa8mNKpx76MgT2VyQBqntTmENyi9J33q3ij
OXV+UescZTkW+OtIZeW5bYNGi/uZUwuB2f2RJn6CsSIUfe7EdSpn0pBqog9dP2LG
XObcVwb1QoTGWfnWAuU8VIc6m6LJRr32X7Or7i30A5pcWCSSkGC4+OFvBDxf9O2M
NNS+aiIYcZ4ZydJyEYRFE64l0Kn1Mk+w3Ya/30SPB/sAxDQq3Go/8/XDZZdP70Ti
VeROL4yX1XLVA6D42szS4zUXnaDdHzEWEiC0CAwBX9oXoIjhMpt0SpdntSJ/VvFf
x3UxzsLAub/OJzW9W7+NmagzxSchkE3etOOkOpQyTheLAtbO/DPZIb5AFNKtthF+
RcNJj7pH1iu6sxfTbNY3Z99XecGw+aOCTV+ZgXHgD0l/c7fEeMP+IS9VzY6Dxgg/
jb9zgnD14SGtwU39ioeaQ1hKtfgX2mPbcBi7KNQVVyU7lg4U688qqxPgMQXq6WAn
xtF9kWY+YGCfZJ85Itfe/wVoU19L/weKESRSsIPc7/ox3a3BiNNr0eUEaesFpEKH
mznHySlocRy0JZAw28d03o4wPkLNzLHy++qxbOmXJbSN2/+zd87yoLCQBHUFqX88
XO7CXZKiA9eO772/jWfgJf7FKlIzjXCwoVp+qooM7506UoHgfg39OlkbuWIb/B9H
pWKZJZO9f3i9yGry9tRA4K9uQ2kdIFsh8yN6Uat+iV1jQgPRhmYkFrHjoeDnqB/G
tZIwaLfIRW2sB117oD0Pa6OYenF9DA2K6g2v45kEXJBFKzu5pPL6PYwgOpUasDM2
XqkfjPjpivdQBV2fF+hcOv9Pl17tKJdskrPl33XPRd7YuUAZV9voswXyFV+GRvYR
Jcat9KtjKeyHzR8XrgHfnh95+46D5qUR+VXh4mNFzwWfNvjWcnFkP2exNO4hdaKB
VAwoyABP9jF2wxieC1mwuEO5f84JwxKAsKZxR1ftl/Sex3xjaF8x7GdkN/F1UVB9
T+3sdyqPfkeENz+4rbF7nltukLytGA5rqXfdjrOqiaUXXFbpam6NCRRF62hQhmog
SbpzELzuBaPnIcH0YQwMRcagbokojcPrSSuRVHsjp2ct0sBqRUN12m1yLSy0dQNC
Co9o2NIeS1Plcpg4vtzo1Ucw+JYIKssft/nZKNAewc9ZsSd8vkqvSubncitJY2Uw
wvz9xMBRdoPd7ay+6He7ovdysXDxRIHO2a22mNeC1wztRODA7hnKpnZD1fAlNG8Q
ZmeSEWHaa5yUKVuMPC7Du/8O//jYckImFBhCDPBOQISciirlFouaqK4RzsCYjeTm
Db6/cvwHDPXCQgsiwMfgDvC8e6XTSfOTgjSWVyqzpkBkRWurka5HRDio3QZbEIx8
1Hd8aCIwrFZyfvJyvlGICdTxvKEUCXu0biy+izNm02+3w8k0qMzgVXyYe/sYEhZZ
DQLXSuZnsijKlVdia0TS7dUaM/9dV9CW7CHQQQQIfISSJgCJUZqSVnzbcwmxB+BX
dk1gb7FIrbO0a1DX7V7SyxXMb1Y50ovqE8okNiOMdL6W1xmrfRGvq+ImkbQEpz73
gU9n0rQY6DoxhSS7bn8qc5i7lS08VVDUb5LFDPsDi0a9FmGA0Yc+r/3GcWrnx7Iz
j2wwq6K7KNd1dzCxQArbgIkch20pQACprMu3Mk4OHMDPT/zaKdGm1QmxJg74Kqu+
K9pefZUAI3/PxnTTdaCKRzseHcb2R2uiFX6HvXgZ8Y6vbpBs2xgHUCA8NrqFnjbn
Jrp5aQvmsMqBKKb9doe67Ok1+DEMhyZ/f1TM78EO/p3+CwBeSKryQM7c2N3MR9AU
HxuIIPQ3LWWcoSe1DHwDwlajPqUPr4jHXurbC36vXqUHlg0vHX0BAdKC9jWi0eS4
aH1ci9NtbqKKumgJpV5Umgvj0eyEFzsKZ7e5FpSQbccCt3X/52qq+GuTL70KkqZ2
H2YBYymivdGsq8mu1SWrOCbrRBJd6+uBn0LJDHpPPXqwmhRcGXuPeageC/W3N35L
PGXcCoZo/mKVHFnAYbl3o+/+IioAxmMp2wSV9Ip6eStpUunhbuPb+NOxVgSrjLmE
RLF1wjH9IB+YFblLUB//NRZfMQX1QM5OEUE1gB1mjNRBu0jDOeP9IUALWIW6bNAS
cu5UMwv6Wu5HGLvrBa4BKv3vZbzAP5aOS7tVAsKy9agdS87TH9MU8clr7Wf6SLRU
mE0DFN7ZwrXDr4NWnpcNTUHOnBlB88LXDG/co+FuNF0+VURqG+m1zxQJ/8iP67le
Hy96UH1Utm3AYcHnbuK+ki4qQC0+6ojAFowm5lMFbRqbfIGJaE5XO2MZ0dJbYWkn
ee9RP2MY1SLlRilGsTl3YkNsISrSvEScaoBymiz9cKPxpkgscxkILMh06zKJ+VZN
RW2hSHEYpHW7lxWL8/L25KQ1Oap2bBqb1Q8s4yQv5+BHXIw1p+x4UOvUMV8dYOfB
js7LfqCo9j6e/sRuSjF/xs7DvHHipcYjH3oD/Ba/jPjL76BECIi5uVI+R1pCpCRt
k5oG0lz0J/CsUmuY/7ukQs1nOWp0rZiJPwoYeTUp0Ojlnr67mxabnUAHaa6lngu7
aBTYThvJ4SjEZDBsr9c75/XxQZK8Ga06YxGCmkbKclYn4Xbj+6Pzh6DAiV3GP4F4
OqZru8dY7TS0wM4hNB3B/7IrDdReODjaND1UJFmGXuVs4nG2OKigoKsfla4go8Ae
EyB9gONs3avhAx5/R8oM3/l+YTALdg08Jie3DDX4hzMYCZUtR+r8fcCz7cJD//v5
8CjO2+e4PkHZdqxQueEqqf242gTjf3SFNkOY6ivqAJKinSuY5b8PMfQkpGyg2EnG
cy/VaWcyCpaAzi11Oe782RfULbPlu60L1mvm2nunn4frvC7ki2bfUR2pXZje4yjt
4iLhd4W3AIMfZAnANwvSvBSrjF/WJ8UjDztqUVId0HlL+pIRulZiMx1cVAzynsKU
f+J96PBIRsdL4MS1BSEMhNvWk9F2iO/LAxDlmuoFomp9uGFzoLObQs/Z5i+VnM8n
D+a0mvl3Fyl3pbVGUOGmAZzAbecaGQvxnu/Mq27FGASITRswf4qtj2DhOKm92y21
3d4dXaKlyWjGKm7SoAvdj//FSAQojLCGekbBrleIZ+ywJSLIHct4SbVttE+ai0tG
z4WB0cpqBhLFg/DzVZCtAga5iP2Nq7LqO7nl3w79jcnshZ0Yl/CVH1sY4mhlek9e
gLhhFWQfVXt8KHRQW42UTREucas0gJYWllk3i8gfTWJ7afpAff3PLBu6/v6vyWsK
01CBDQ7ehKbORPgG/QMq6Iz2iiyBUXyEvRkH8GjdLNnmWPKDzSFBqYtkRxi2aH2H
Np5AyHo8gbPWvAtbz6EViotQGbK66oS6795oIgPJcQqkd5SG9C9CpMVXDAcm3XgO
CJcvonqu/jHdh60Akx/wcgYBDeFMrPn7vx0O6QQUfQjPd2XhY3VbLtPNvOCZflPF
ERGQzbunZNsBji+16VttGpnsxyVGVAdnpXloua9rs3CWrhXvhGjITewOiiv5rveg
7ZqWtkPqhGJcu4Ru+RWZaAlUOq1U5aAXJSkfMN7pLblyY8H9AuCYKE1oGtic3cn2
rTD++nwrYGeIfjN3VoFXHI/gbI/tv9Zo/VPhGYloZnO3It43wnMtn7OHN4nXWsHw
yjxS41E7JZ5Jek5yxwRkw14XfjWUCE7ATlUDdwww50DbI2Ga2BSb78OZJ1L1eTgg
1EsVlOq7O4bkhgIRZI1qDsl120+TEVZh8xuS7bPDXTRyLJq7XGYXXRk7IsCsA6B+
fN9AV/2zPxnWMHMOxeo8HJuJa1HB/qjJElYd6I3HmQNmKsIiJsavi5LapkrR7If8
ZBMqZMc0gdtQ1Hq8lm8V3KVPxjYj5+riquABODG2gy6YNTnm7uMszbeXDyAG9Aoj
OKKVOkZEJ+74ZcpIWMI5Hc0+Gyegc3n8onldpYM529sQtCPorWdSADY7Fpsr1D2S
n7ATOkO5mtGbOFhvhwSYhGYV0D6JGgKyNIROzKDDF7bYEgmBXfCUzHoWAPhKtK0z
7IyQLX7ir5P9WXJtA9xRtVm5BdlkEtZhBtuBpfMCJ+Iwxe9d8iGwnkS/CDObIM36
IpAQFBLGGf6pThgyAx3WQEL4JXby/yZ2ssxDQw6xHHmRficacHTVwORFyO3wsjdz
Gw4QDcpf3TggjNefndSPWvlGBA8bSr7xDEcZWrX1trRMspvwJNSVQ9mmwdMtrgMC
leOdF8he+XAaH0Y6pWHxyTipH4IClttd6JozJplqm0sEihU+twA3J53B/CBuiNMZ
mKh3Y1j/9CpOk7DVkDmVnU0AJRzfs4X0pNbR5hterMfVxtH2tcwKLLvQBx7n5jmY
20s/yil83i5qVJHh/jCX1AAsU429t5yeQq1ll6YPn2LLQXAmzN1HRFjL8uLJ5TV4
8T4/f0VkGxr39XbY6Cf5SeTye7dTIP9vlynLurBJe4PYq3K3X5GMfWNVVjnDcdhm
Q7IJxQctyLwenbsZ/99w/avEO4PqG97wjrmHLVtom9A63p2KHjOtzEA3RdPe0KUb
eEELbDmRUOWExKUEVI/V3YITVD7pZaFr2WKHQ9wzrQKqt9PpbdR+zmz5uSWZrz3C
HhsucR6nDL7+ZVvyB9tr6/FklydT+elCrPn7tMXPVkh6Unu1A8O6oGQ6rjOT8NoX
QGsWQY0rEH2sxoQ477gBxTZ52yJZeJvGQtrFwV1ueKdvfxIhzFnzqeEO96iZp8Ur
RokulY5thcN5APRnY9HCnPQSfv7JbYTyuoU3NJinkfg9tdfVfRG3L5cHr/WHKcbg
6fAZqWygDwoCy6xazFD340H/LaGYOx0Yl/3cIxugMf/5E04cyxE8y+ZxeKxaYiwT
KjetCXJM+Bui1G0UuWg+MNH5gfV7IDPmAd8RXyyFZgKS14Xih0vyz7fQ6E/rmpdd
HFO/5FDH89dlAJdStmi3tSDH+z3HK68rF/YkGbpGXFOBCqsKVzjq4l3US90TCN3B
TeM1QTjVMklubDKIJnwoCPI1fN45E5tjT6bUokMdC5EmLczoQhSRWSkBFvSRaWIU
7TThdxdJ+2x+yqhUYLjEdo6ouK6EFzWXnkumpqJzBY1WKmIkpKIDNr5Am9A3kOnC
3NvjNbJzHwMbbX6/TPaFhucW3O/xLp7uOWCJn6BtBdQ1NLrJUzVjgpKhsID3BC5w
pT5EjHfRAkNHtLylWjrcdMOsuT18/cULczFSzSG5F+MBKnvO1nEaHdwMODFU4eNe
PlF2YvvLCUyKNYJk5U3uvdjNnQfq1uaWjLyevlaxd94INn7QAbprMagHuyC1dlTV
FDImI3zRpmPG00w0cbFbwmVLFf+F6lo1nR7/6s9MToRrso1ESFWyMm5CrFRFvGYx
TwKcFmmpw5i0wbCW1lOydI9hTYsG+9UKEUOQWdse7DeYe/qQ4aXiprYz85rNdRoa
a9Y9DHtEz2dVLkCSH7LYiVVRaCAf5tlx5d3xcn4JQzUrSQ1unMgxGaaduYCzh67G
qncoXbe9x2bZmJLJh/G3UR0MLybaCOA/ypy7IAFKPf0IIKl9HZ+oBzqU1Bki0iB8
HteDd8A8C8TvETrVIX35uJbGziJPYZLXn90jSIWDzZOuGNHoaCzakWSnVk5A6xrh
La8YZgWdGYGC39xKZL5aJB36cs3lnYpAfSladvu5dcIIBNDhxHS7srZvDp+Tyvdg
J+4Dw2AsjrAtUfxxv+CEbwFSBsmoFDKgapUouxWvXUQvJ3GDR9BYxR8HOEvjCSgi
BdEUi1spxwMkuRYxvlQMK00Y//i3M7gLQK7YsWcmaT0PgA9soZxGYNUP3L8ynCev
OQoOsGaKmO2tuOCvyv07TxNWMxTZY6rvdIOt5NsymZtoBSWYRj1Yit9NvqInalyX
LdMHRhzjSfA7TUYMGs8bQLRKH0TsAUuXAeIxBA3eollvXbirdOaKX6lv+qYJXfGP
krHcNhAi8R1d2Dh9I3FP4Iv8OJA3BDWzaJdJKBpEMXkkPyC8RkFFrFCaQ+sCQIbZ
HbqI3czcZuIkoML/8/ExqKS2TaZj4hapHTNApEvMyermugznqIpvkjl++bdesY3j
F4o230/Zvowe3pYJlsFsV1PDjlezr9b63D/vVh7QmLpqHsHM/5czPXEcPVwrAnU1
UL7gpOUSBGzJCpJOUT7cvytdJ2lUSHsXPt1oSoj2qAnkSpwERxHi/jDjGOZaIWJt
JdgalCNFXGkZk5ARU0BfOBF1WbP/rLXNAmSGeVOHMqPEOS9L++lqYdhBuZR66Moz
SlGVpY90Ih7MJfOxSKNPGroP7ChSlLWQabcyXSM7CZvzjVWTla/+7QhXWJo+jzzW
IhclFNgqMHTm0FM/bNCKSlamBq04AHTNhi75sRHZ86bxEfH3VMHKj+vR9nNgSEJ9
M51t98lQHYADJ/1bwy/6IXYNt3fGdHtran4/ORfeVidJfHq0rxN7dUbQ9rt1KJ7c
CdbAyj2GH8SmORGy2fL4kgvcjntCDoL7qFa8tdVAq9KS2EjsS6B3AjDcKs4o1unw
+yW1jN+YfE9mwLHkhPRWm1wu5U0oD91KCEh4/vGODBV7qb1rhQ7cydZSVBTXR3Ch
ZYdbxbAnhuTONR+Fff7CgNP1MqpFQXjExVgtX0/rl4Ax3TLwbXNxJVQxsGcsKLKW
VFTTiwzU5rislVJyFIxA1suAc7ukDFeAVCJDDftIH8tWOtE6r+3Qky+N7Cg9ohIs
pK1t4UXiHlMzQaCN0Sv+ijN4QqvsOKHXVTAEF9vGNuHU/p1QjDSSV0CNGkhLWG6m
96jT/AezSFEBlF7i8OgIKtN3LTcs9L0hpmBWn+G9WrKL5/UhMJqSR6PpHeisf0cQ
0QDKw/26wQ698xHur4srsGX4031dCNafrbCzOBouKU6CmqXirprvNhZpIuFK+o+k
G4syMANQYJLJNKhHPr8EUTNduxBNii6D9PMLi630w/cYB06/mLaeX5KWfwIfbV6g
xHPW/3idCWf5mOr2BRwEdSEbBVtqJwQxBA5d5VuDYskfEV+gCK151DMVBM/DkS96
ZlcUj7CdxvIPFlEHmASbjDjUPbswGeTiFpcjk8dVsyTUxAGRcaug9NK5K2tqm6cc
SYTz3/giXLTdcYHDPyIJwtp7Z46Y/HD0NuUaWU/eXoa38LqFf9zeeTYeNtCJRsHx
zaBc4Z5E+DZ8NaLhQ0MDjSdkPHYCVkgNxRGpfrNVmZeI/RcsER935VtWgxAT7FtZ
cAzuSUj0z1YgvQ1R5g3wtm1F77nC5ImqsIAgp5NuLeSCgOo90s3i0ELr8DQAENMG
Y0c8hPvIk6acKX+z1v3yxRILYz7iKkDsjfh4f2Z44I+wJr9IZCxtTRxsoMHMAqH9
1NLeIkIob5LBkGECVqeDSGN/pd7Ww7bYW29sKRfPW5An7QFs2LtDcvsy6weSRLyW
HibbvjSrnDx0lkxq9PSpU/4tsz1Cp8IVDV0cAHrAz/Gqvw+MJmKYh8mari3kCgzC
nQQCY2abOge4/8ZbzFWdMIiUgGzFoCGTWrvU2x+e55qWc1OujRa8RrE9fFTOX8oL
PVayzUjPMF6xd4K7cV2lPxKyG315iC919YbaoUkWZwkja6cmjPZz0vb5ELQWhBI3
An0NYvknNpzQnKMJvc3ldhRHzM+Ud75jwmZs4uZFx/xpXAUNcMvy76aPyDPEZghr
QP9LyITBUcYKu8TxbP6Ax4xl5BcHqFEysEU22S/T9gY2wsUDgh4b5G2a5HmVCJ9n
rQ26/K43Y5iDpUSb0NtZwvv7BjQGRmF5s0teY7gftdq8jg4pQt7TmbD+OcqSYFEe
2fbHHhmdMF/KPEQxG/UP5yTX7nIoO23oGZenPivjyobwB10B89q3ZqbzbwWknUkG
M0SH2iLD72z+43bdzsnc333Q/faVxKYxAiAHkQKsNaNAIKP2FlDsxpG27mPH9mCz
gpeZGp6eXZuHWk4HTdhTkevXW/ClUkZmX6RDVdaAs+U95KWRpYdFCxzMwGj5yczT
Bc1Y6+S5QPii8qmf4Hoar2DsJNPts6K79SlS8uIo2GJt9OwjhNWn7T1PUTcskGRY
AMf/x4cTgTIbM359ucAje0Tk9N8u7lR3qeuBNyIk9f9p74dL0juel5fH3amlJklZ
ATxNt2SC2/skG8ol+eEGz68ZYcDHDHBwr2XdkGxqjox/r00eCmEUKOvds7bAcfc7
HVXFUz8BsRfl7KZIeJcN/ZeCPBOrHm+CF1KqUPsoRGVeHmafcCpFE0KIxMB5G3Ll
4TzHrZRfb0W8+eXoat/2UPJOTDyQAf4ki3CAbL7RAs8+fgsxhKC0SGb0g4EIGBt+
tXkpMv81O16eQQ5q9oM3FqLcFIz9v8/Wq5SzmmPWt/e66Q+yCHTPovbUFS7nQDQN
gr+oFHQRXC17E/pLs+owGoiG6puOJa/Z6yxMocanc823RPRnv4XurtAEMOxxQgx1
aIN+BlLaJ5g9wqBpOisD8C/2y3rW0ahZJszSX/Q10wpwZmBi0VmhO6C/XmwlDViP
VHM+LG6bc8vHpC/kSWqif4G6+7qs4OpKuOAHrfeVHGGiHpoJXra5Aal2ZFzp61xW
BDQFSVI4BVTiUx93i1PN2jMpe+6zoCTeHzBFlf3Lk2kfGLd5IBiYRYH+XdOXubpm
2xzYqbq5dWEjkScT8kT65JQhdspxW1PNL2Gazenh2BnOJoEKIZ8bzcTM02n87ftA
z8C3oiJfEKWNt4W9mo3am2/kHen0SKcvG3NKsLETFjIPshZV3rJVAwJfvf2SjPzt
FpuyKcvN2AlP+1nhL0/SVWAu9DyBKGDXkCkkde3GDZH1pst8DvwfpwVISp0N/HgF
hTTCydRUhPkZqmmHpHrRY4k9goSxeYG42RzA1VyyEQgVQHJi7XA8KK3Ks6F+ctFi
IldrWVEG34+RD+70KcM6YxLOZbzXLrCWy/khaM0PVyuEStwybaUNbzJZ0jg1jw8k
WrsY+lh0EDbmkQyeDk7s2VTHkmslbfD4op3L4eozxhKlpZJWgvN8SdbFGVy5QANW
nwLKrSLqdwXFAwE8Eegn2gvrx4Yg89hc/lvIoO24Hc1Is9eebfoaiTP3wpALNVvo
WUhc2ZXamvs4A6yVGblKweB9E/FbVTlBx51SExsJSqNZsypGAhTKLYR4YlxAtX9m
BBxWlgIGYHPFGGRE5BMeuxJLgd9zmorRGBOYdeJyA6H+Ox+kzBdK1H9gwsr7SmEM
RIqYxJl5W8LAvvhhPjb3kwICDJt8+lDH/13hE4t8ZV38LuNX44KVIn/J8QS1x3VX
T3bGad2k62yngS/uXptoxqEf/VwPuyxnql0xbgYUW4FyNmixQD4SbMMcCN9k6suY
2hipvmdVQ4HA8v73OEakIYtSPW6KGVLxQiMFMbT29+XGyw9ZQC2zy1GTaONkpBLz
jIpAg+ZUYoSnMA1GIL4DcCP6HNqQTKDTj8l5SZq/fm52OLPPEPAyS431c8QpkJVI
nl53uBHoG1GSSy92K4wZoOnnGBUepLRm05981ZeqJJ2JCEc/ROK/KtEFoWIv+cwV
3xzsFOmVCwCxta9l/oSUTHGgSMH891KjEbeSn5O2IGvJG9TIphlVmlgsEPMptq9Y
CX4Ee0OvBYxOFeDjq3+iEUaiMQ0Xd29QNRk++Yo/Eyne0wnsKqirv+rEx4zg4mxA
XoTwpjzyUv1nx5JKWp4bYZGQBP4obw9nodFXK5y/L1VZXOXoaGg9r5DcxlZ8qhKU
Azlv+NQRgAKUybDU7bWRes2LaADchaWCx+RAEoC8xKvJs1MxwC1W5694s/doO2If
hY0AmyYKrnnohBGts0+KAqWaObbF0jRDm+DdUDczLQWVaW5wA4gwGNqHsGQKnPdL
O7jg9XJLdVrVCspDkM5pWwOcK4DPvhPZ+X4Xeqj24hc2kOCpQ2DY0y5JH3Ql58q2
cZ7MC8cuBPq3HQpYRLr+J6/2IgUDcLD5vPJMfVuNg99HagyMOTbm273OOnLLG1pE
qLdAx8Zi1R1wPJ4dOl+GvgTTD/j/47Y4MbektsSXsoT/pJwhKGxO+jnoPJIqIUqe
TFgEet6+IMS2qX1iCoTiCEmQz+SEIMABQV7TjkJhgoDztR1XEdO5+k09heIGG8rR
AmzDsFWzqPQ4lFdwx/txb7pc+J1abeJLolMS3DQLMnIdsNNVwQkhD3BdY6tBJ5pv
p36reXrHpw3DQsACDrzno1+1VrkYGMR86hbqaHEWoGkJuAKCywqBvv7IVnR0r0rQ
nnZti9a90ha991HPWRPGQ8GiBy5BRG1Prbq5ADR+342g4DPgVOkgTaxoke3v+bya
J/RBpBzllPE+7uhGXZx6vxyj3ViFrYdf14qZFl01+ekE4KZCcLIGfY4htQikoyR0
S2SJa9ZM+FC8UZ/nIA4tspqaewxTT+6ZcMk76mqUBekce3AYVLfucmbjK7x+gVwb
CNOsBwGhDqgKUCyFrQbDHI9GCNmUyLqVNFqJ1+EXH8zdoQUmb+7ip8TX+5ft9BYV
+Og8KD2V5udwbs5Lm7tQUJISe3zcRTpwUkN+NpjYO4nGOUf0X5F9oT0tlIf53gg2
/LjopbvZjnq7NRx/ITQRn5U8AlecyArEpnhHIuZDWYegNvDC3COFJON2bzEeUr5P
C+iFLck6BLqLEtW0b/cOH4pZU28RxU2d/WLbeCUDrsVhp4RZJPvXpqo3fMc5rrCZ
sx/4XYuwJ2UTIwPXhkRg/MqsZ+dLw5bZwzrQ8WxBVvNDwSdhrCalxFx0WZq5Nj9g
TXaohMDVNCmikGBZ93w5UYpZsGBN7Pcz43xuOwopynNOsWLPKsw+YHfqmZrJDN2O
XDQdsRvESqfPaCKaOSA04osNYywqX5PAInuu+ueCdW8+Ml2oHzuKlC+6VoklOGiy
J7UfLJI5luVOkb0gqAyOO4igjJDHd5t6ZIU4maHNaQG48TePmtzoUn8WPFzpj4C5
LmzN0/mAmBy3VzlaXaxtCOuVofBDp9JYraCUvcamIfv+RHwIjheRDhFbYh1L6fdT
kHXjAoUey6vGJa35YZtcc818afM2kBpHAcQuHJHU0rQTkGGjiK0sh8QbXT+ltuxf
xE8va23GIuRFzA5lllYRIbJARc3EE9z0bgaCVVGjvP6zW5W9egZYKda/XfkOgba8
sqbShbAolQMsERjBmf+sDo8sIvXx/2y0vAkGqbJ5R/euihAXXOAYaYtKM3rNvArx
hhtOvVey1Uzy3pKVGZHThOExLILfOMhLaZlHyPuUS0oUDdjNgL+/vJv5FlyatGRd
LqWvshzzn8K0r+qGKGEoeRzgHLxOE0uFvQ0cA4T+ZyEyoiCl+MUZA4/YwBoUQAk9
Q7PdGYnEZ9H5DyBDOsyp06V1ELU31gbzUgbmbsq8lo8G5Zontu+H5EFJccfNdCDd
ic8/BvkF1PC5b0M/3zbdPvnYnrxuDjUA8VZ5DdaXw77lDAnyK4orQgGl4jILq51a
wvCC6TnVM9e9Vb3zOLuvsVGE2EXUp3k98uK1Mo5P1FDZBPpBescxdPlGjRZkNuOE
xa0PlJQd1nSLdbMF3nZTh6G9X+uxQhWBLKJxlH9OAZQu9oKog3F5YbG75a3zMCEu
iEzxQjT1DiIJpZm8rc+ewK2IkoxMo/qM0k3Xxaz/ibsCT+4r6O+NamXbO2CrFOzX
j1YIwxVttRr/KBTruMjoIorIx4URDMq6BZaZD/kjrwZRlgNVSPJoRTyXLChfgzm4
1nsJcNb9nEqon4ZhGaUUxZweHD0FexTTlP1Oqw883IQLcIoS3UcNuJMsX7thC4uI
37ABGzgkiIMqHcuPkoujwh514Ikk3fJqe1XbFTDzQTjchiyg+x1hanNqNbiS1v27
KXUCBdSzr7LtZxTemaqNyZQrlWCNLfjx0+Sbq8Uj8sFViaZRJg3YYpmZgVUsotaR
h1sYPBxyrj+AEvaAN4UwqfpPqrW6/voCTz3OSfMnLD3KqHmT75EsZAuxiLrG9yfb
e0TaF+zBNsFUhraPN73J/GHOXcM78AOzVWOlXmT4KGKrCbk6gXqQO3nkLn/REJzV
OunTvuR2k21ZK6neO1wU95JgdFElACOCXYgsrU5X2RrDIV7qwC+e/Vld5T6s3Y59
JAT5TlD1Mpr9d02Vss4Lv1+xBnb3gkl6Ni5sXqTtozecSWeqj2NnNxBCbDsNgxve
O3dqjzQBiDLsz1uZfhz5Bju4WXqa5uu2tsdAvQxaq5WZKDe6B92H9lwky2vhxHjD
EKVivWZMBsZNq5+cVdCfLic1pypI7N6E7aKWt/JVUidXxtJOJb7OkeBljxLESWQA
p7gOqRR52jqr8hWRjnppHC+A1gA/L+2V97g/ly5ryw4mc/uzWo6r0bhUdx27XHOa
3Rswqk1mwig39lxBAfc3kaQrqdswYwxgHVxLL1xM9VAVBZEw6UX4+Q5cAF5iBsAM
ouJffYjYdqP2XGyyl4zPdEGZ+nDNGzvK9xKoikxT2bmC1x4RVezuYckxbroJp14w
2RP/U1xCmSA+2w9cH4myk7SjgJBqEqrYxif9iKcKgschk7+f+hjasPXpx8hwXcHx
fPNUx42t9btNdocTFfnjnAHq44//yJidaNeoZStEk9xk6xiSZL0FHHq3nA76DFrW
2IIUq6IYMlZQ/6Nwy/EXpeefHBq0rHFujWWUhR07xYHVEYt7kfCXRCTy1J0jGX/N
QpbPZesXsgtwWZPniS1PnYCnR1LCogOKfY/SfhKUws6ImjMGk2QpsyDugimLixbb
C/MdTcmBEDSjCmLGgYMDATiRg2Caz0ag4W2BwxqhztiJ4XHDZi8WwAhUFsVqn4db
24Ca6tMqvqYNDmfYZuNLYPJM6mDsuJ2/+hSTCZprG9fZLdQz1sMUXCk/2smUWBsW
C8U3Qs5j74Ao7Djl9KCtm4u5myZzNa26YQ5pKY5YtHvSi7b0wwExy7Ku7kqAhymT
cdh6pAbOH5tiCEodl0cWd6hjgrbS7MzBnEjmvHmmHGBibT8kzjv3RxR6XxklgwsA
+00naUXXvWzniRMRUarnyFXbSbQ0GRW0j+cGSbEhIVRpoEdTwMA7V2J2xwuQ1PUW
XqkkWfZdPwOcJ/why21zmk3YZ0NAM6i0wJjyl9oWVU9tTc3N6gDB7fydKACdn1pE
taWoBnyHCnsf5PxkthhElmOLXfaWmFaB7Xv8CQluzxnbbXZL7ho6ek9O1J4jOkpu
npRKZ2r8+wVSIZpZJArSGJQEdcR4nIerSATcNT5Qc0qtWaVKJEz/edgNE3zEySde
3V78p2J5zgirZjzSj0p3fz/yaUcW0UBL7uc7z3YoXFJPYA3TAfd+6RqPzXalA5Nd
Bit3+qgKWYug5tXn3Q7dk8iPk3RI6mj2zumoXaNEMH88h+xRsDsJu0+bZjBHb5MX
PS5Z79+Pm7zutKZCU7kRMFhPX6u8+VJzMeHCRqJ/LD9KCiGfogxS/resUD9fzLw9
9JqHj9/lBVXNd6hwA3Pnfow+7Cnspl0b0YheEo/wKczJmjC8zE8lc6Y1nrPQMQ4C
XWz3JajKpNmeF7yBu+05dbvCR0psl2yFAnI620SaLTeHxGmZ+AuUeqhT4aqeEZxS
ubssHP8kFP8dkzbc9syUpRyechYZxrBzEueDAQ+2TsDdJ3jdmuSuWhg2aCXXF/II
G4cnx/k+rFhnEn2Svz3eNl8acuRfwoi+2xsfRdkFTV//Bqk5i8nDnXp/d+D0rOrP
fzy73d3VnLVp7UCDMtQcICloNQUOjZ2m/aPlJTvJDZJZTEx1Q5LTLbtyx6lFv0ii
iWSf01mCN7dSx6P/M6x6YLXuBpsMHqxM57MlqDS0cIzNd5D40WlmsolxD6G6NF3t
dLYMWm3JPdKhjmT6zqYH4LWnekTK3/0AUbM2QJfFZu4Be+nqBR37wcuVL3lf4NUh
rw0zRv6gBh3HjWdI3agDuXItUsU8nUbRzuUn2oimvmP2ds1eOW3SV/4tmJ2Mksky
AgqfPS17UhBAwzNIv/MK3YLjNiobmz5vTCUslgunxB/qbYszH5R0QC2JCPpmRno5
/4byZW9T9z2aoFgl+P7qgLTRR5b/FEt76JI2wxcR+v5e++iRyFDHUAkQqmooXkFy
SWunVDzY5n4aV6/SuNUt7VJIFBsYvnWprcBIB89GYZgfvhwu4fFmSD8fTjib5hMF
IKYyMFC/ZFyDucVrbxe7wqngJTwFNOVWxgRBjqYpxWZ3ZhXMc2quPqb1oCOY/KGQ
DVQzWBjF6B3qVEKvwMhBEn2I6/PQCTofWCZDC8BknO4vgXM80Mko8VfQ0uQE7bFq
2XCHb5yXt1xwoddZsa2K0w7hplQSO5uJJSlc0XlcbOi6jKx3bHljvsB6tp5AdA+c
jw/bL0ZiYMe04SJ5h2/1Dmdg92FJURr66/8v/ZNKKpEU+TdBS9sgQYHgD2VLa8Tm
5WtVB8uS3aOJNLasPAdZ5DRF1KcdLSrsDGWkaRz8JrDuMYoE+hn3no01EqirC1+d
3uHJahK0YqERVAVnRbKfxb2InwBZicPwhNcgvzbSvTxuTtJUVDkARP+MTJQcWUrY
154YTkfO/hziV8ioFuDbAE/rjwwvi7hVbYu84ZaOBdBZOCGeP/4OiZ4nJkA+AHoi
lY6ApZmCUGchHD/qtkl7sDHm93UCMRZiGA4oyWhllsZJT9PdqAP0hWCVkU11AJdE
HFT7Oy/IN7XrsEcyBpZN181Ah0FZq63xT/I0erqkdYA/4ZYOETQdsOZ5ZdwsMEwE
PJL1dZ2E28xRtNWd2DsHCtOsGGWU+/K1MqW4iaPwxcxaqNu9jF35l455yzBXxEwp
bDtsTfp6XZiANCsboNjxs0udJJeWNL3+fY6O8a3koJCtBb6eNuja+tEk8Z6fXg80
aQTxWrcKeam7FzDoVXBPVvXenkrgBKa5jwo8tPCRHxNIOR6EjtONdZRFsAE35RRS
pS4NyEkN1V6VkXXzrZZ1pl6un8hMAAIJapIDI54W2oTNHoaaTsldzyzZtSM4U1Oo
7Z3YjtaV3wWAPLc2bWhqgl4x3y/vcqh349XeouSirMA2qBwGn6UR+3X2QIESyxqu
lWMxstK9ocgCJk7QUXDuhWx863+PVrusrEPpe6x0vejzfVFcEE6Dl4XLnpmyv0z/
Aje/fA3A0l2MRfUXl4t+MUUKWeofl1d3pND7FuDc2Bt2vSGlxGm5HFq3sYsB4ac4
HJuwL/SHd/IePDaHx8dFpzm66pp4+7WG/yyXyFtRM2zFXxeY+sKvmb3GRuEWajmB
516W6NIIvn9Ys/swZ08KDEVQ5aXJiZTHUAe2dHbPhexooTjGrrV30oPzgK6v6SIB
EKZ6mGv6PKD9PHBaB4M0t4dUPKrQJ1wIoHWAcZTnnPQ506MBwou+MgtksXfjR9ye
q29B63vcjrq8xWk8MMU4+K2eOU1mjvoAfQmTs+qZ+9GrKaxt077tk/etVVk0ljBT
WUCuEEvQ/vM88IgSz6YJ45/3YQV2boVEgWQd6dDXbcyFiTLb4VDQMrizpQXdMh2M
5iYVU3ioTe1TTNiMioRfoAdoljQ7JVT1NSJviyFBtoxFO9HDmplhgJTo6KZBPXcG
weUTH5p9e3tEbLb3SPdPUd6hDSBP0JdxDjsK0UzDtk2+fHoXxxZjAjeKfwt8HpZt
CIErUvxNzfGFaQ7jGl5MXxsWt43em4izQf49QxHIfFWhYzyCmF94hq4HyuDRvR/j
Kce0Xi5oEfFy1VR892vzxCAZ84HI3ytFIkBexsIMmVL0z6Xvia6EWVbDm4mHElLZ
qhcGRF8NHSY9dUKmWcb7mqpdcjLGho0BE/w5a6n9GSD3RH9FqdzuWJEnKd0MwB0B
BS3S5NFmt2wZgoCxbjpMTAhjZjTApNP+q9za8bxwnm0zNPpAO7ima9LyxsgQXfa8
kseliE/6DrHfluF+5Yh+u4PTrt+IemnQGdOAIjEKFNiocX9MHcBkC6TBNxh06rsd
p8hvSbJY6H0Ah0/G0K3zM+AHfRbes8NHtrwKHDHVRllDheFIf8VYwZoj9LT3vFv8
MTQlaMvlclUD7CEEz3kT3TgW2VbCccHxTgOjqRTD8or3PUIjBFzZIdcdTlX6/e2l
T27pMEZMTw+UxYiKoQRRpZpKgTdAQ2fTs985RuoDCBgqrqnjQv8uHobze6yizE/D
ywnGIR+V2Ee1D6uS33kceyojkwA7az5PKFthrCCQWU0ywe4HO6su7G3+tucJyZPL
P5YvozkXlZnH78Xq1buUut6YR88VHSVV5TBAuBTnluu6CAYmwr208VhzrHzlNa0l
QPAt0j84RlAGuiUVKXIpUu1lobKQhDjwRECVoD+SC4gVgcNPtbT/i09W+6iSxAHJ
PELCXqZgU9hDlwkszsg/8K0RGDRla7mGDlQ6EzF5Ghxiznhw9mDI+nY7PxQBd8MS
LeQNhWIeJebL/WeDHOE4Sq2c0S1C+tSazXU99Wz1uay4tGpnt+8nc1zEw5bnFo42
7VayvwopFwYbjZQbzAFHa5fvfx6OkHcP2zPe8MCgDomoYun3ePt5+I0DSHO9qgHA
+c0GvPAm8ZBO4KEvYMI1N886L3GSsoiFC4edyv4U2hu700HUjyyJIz+CyaM8lBnI
7bZuzfPlOUfkjiYeOza73QbA8TZ70ombR7Sb7Vcrug1RdIRkwGZob3SHAIYxU49e
A28n08fHpLJu/j5RP8SgSWqH9/tcHW7IPVEiYIiVJfpDeuRs7HesZv8+Jwqtk9WR
QL5xmCGePH/lFESuwP4CPUF8SD+K6l9Tqy+ApXtwO08SUwGLP/ylrSDvMoezFsme
1Z3C5I0OmHV53wNxo2m9ZeJtWeAGzwKVFw3/3px5Cce1uaDu3HtU7leFkG4k5KW5
FWjRY/RGBjyMCK9FRRyLQNsRgezHQT76OaPhAauDHZOrd7N8E2pK1FvfNxZyRLjn
taFlHbJBths9+l/uwa4hwgZ3eAsPh7QsFliF1899rA23OyVE2e/XPfeJfVPLA6zw
r2ZYqJO6tDzFriBKjwPj2eutMKpoMedGHjS8+6pQQI3px5hd3MX5Cln1E+zbRETI
vcG9CUMS5l0IpKyRd2qCHaw6JwGHDSnxtPJ0+/UY98CFyfqLi3Zk06ZMuy/V19oP
94MtXzivU6IaXiL04jhA9Ko+ymnLSndtxa19Gh+Ymtp+AcvtChzOFy0wHtTvYHMv
pvCQungN8R1WMimthHTeWrBBh9jzzLQol2z0YeGhx1VE2D3cpxeq2TQSi6ibGEmP
NTWX6B4d1v/H//F4wpurYO7Ypv1BTEc+F76v3daiN/6rjdf5l/qsDxk6WGm3alAr
jF5Zj7+2QlUNyExXZviCgjwzqWFe2A52Zey/bGYgdaJt9iADwNHylsOEEk3aajWW
krXp6yFGx4aqRvaRnERGrsbdoDxbG+uyZ+ZNqqdpueX73UmD5eSxc5CEbeYieh+f
gXhpf8+UMtdBvt+nMG4m+EVaBWODnnM2O4fFjKno2Mj+Ey5XtsCVr7soq4KpOHEd
ZP+WEc2OTGYtKqX5Is2g0wW2x+ouJeQl3Ut0HT/ouE6VWXv5QjzpHlB/TwGMKyLt
3Xuf3XtXWnPNZIBhxi37IqDWtYgy5spdqGC6W9bJ4EqxBIXokI2iIrC/ZBVIc6mr
rnpZvFa3AUuy526keh9YV/G0/s+GTFbbHXtP4Cpbn43gYbv+yGpA7gUne6CjjleI
DC8vi6F58OD7Ns4rrO/n9QfFH3NWUlEIBklfH8DfBkxxl7uHV1nOM7WPlhEQiIIG
9OQ8WFp1h1tasRcg2O6VNYr1DqEjnhuCrXwJN+Md18/U+TIxusyF5KQ5Y2Yxt1c/
iJiq5sIpAZKIs40WwqxqOJrlXxmhMwMZKC2FEUkusqfPIGsRfTEQelo+KP361KDd
an08+iGjDdkkcBB4TtGe0mF+WFZ7IXXFaRA0Q3UAOPRFhgj1JQ4dBRcAOlMXQO1Q
Fr5UKVx35sLxO9caHxfAj+SFLqfIYWoEmPlbSnNFexDgbaLuXg2+YpchxRiAQYSM
K3ARzSP8E7Dm4ZFpRsdgZlzl/oiELz4AQ0sk7U3ReKZ+1xG4RToIb5M1rX46ACYW
m3w0nmiWzUBRdZKXZ1O7MvRQDWVzfoetBcMYDeo7HPfTtyse1pFtwhMMUSW+9GwR
jHwa6NPcLVO3R4FChoE1nxUQWEyVXDC3UoSkdsOA7vU9yw+MpnmW0zwjbPYM8x2f
dW5vEvy5t0yhnDNkOLklXe/YuAt8Nno6KEV2TWWcqcpaVtJ4qI85PTYRwfn1vK0U
+Xd5uV8bhafNTCdvArWokujxqFx/ru7Z9y31Cn8i2g9eTRt9HBAdfgg3pd1qLpd5
RJXF7rFLtPH0qn1WSRLM/s1xFIEOtbrS6b/je2mZx0/jlwLaOn8wzhoxi6ddRoB4
DZKH5jkAeNFGo/ZZaPjhmJrWz3yISIY2kmT3EyJBbsoFVZ1LddEmbLaM8tJ20pk1
lwJQPtZi8BPVpYF3jUgHxPyfOdNQ7HNkLloS2Gl1adlYjrvDwgliG5wv51SiYW6h
QO9mwOeGreR/sfqzBYUYGe/wdTRn3p33LEZiQtB1G6Qqx83ZcpGUVadhX9c+x6Xw
cRLlZO/M+GDH44oOw0l3KwSGOWYbQGfCeuI08dIFkhxLcgH0YcKHRKTr1ikS93x0
ypqi4XioDmkJWIoF/kfjHdUgq92vua0i7n25E0gxtB9LQHgeHb1xpQCoNqXKEEkH
VyD4IEtQvHBDHHwiplK2ZCdROSZlEACVBx/AHnt4YPlhd3ibJniIbCMdlNB9boB/
yehlKDri3orgv7NFqWhR+9V1Qv3y3gcLLGAzpatMC0R/rwBsVjUIQTeOqBUQJQK9
Wy5I6PIabGKpwgMJZzG6yxaNhIgKbCGPOw7KMQNPq9lztAv8ulA+g8VGHcQEhM59
DtukNNd8djqrHl6ehcxclHA6rj4KPn4QO4VeUbn/Crmky6INtW8GNikEzgsNSXcG
l91T6EJg/MAHEv2Gy+0yGAFJN4NI4RiTPAX3x+4mebFhBE4GsvTgx5KNtBnh2E8s
tDFyLElv5VBAXPQs6UqEiJclEb1sACeh9SwHIQInfi8kwUCyUw2XIp9MQvjwi1RG
KD5bAI71THiVY3p28kJfSPkL8ASteMSmUKVrHqwM6TL2lWu0lZyE/+7uEozIfLmE
pRR1fltxnNOUm0W9u6gqRAe4YTRNQ6sTZM9FRPHh+6+uogBcv9A9vq+bfAQsUck0
NAdSiYySYbUsO0OJNP+UHdktvdfBJx9WtKTGePWr7Q5gZeCseDzNp2eLQz10dp5W
KPviM/Ecm8GCr0Pg2dA+WejdE1QI5luRsX685IXGaxdmJbDpCWiKJFJotggexWYp
47aqpsnEM2ItLrbzvxWj0QhdFK43wZC9JOXYUSwJKJdH+ZzH9k6q2Dezf9hnvEbb
HVTHNQ2TWV+eQR6jXegSb10/Xvuag6AjrPxdH41h1SAAZ7Jbr7hqoM27/xPc50Ke
6nubYeF0deLDA8ZITfWZz4vKbW53tW178y2TQqPR6lkFoOVTrOKD+0ia87w+CA4+
Ft+KnvoOVnRdDA6eXI8tD5fFsxydzmgsL0CO6Lw+WwDhSDVuOfcoaCVSLzPfmCJL
83F/IFtYV9+gPIYvdchpF//nOnhYYai5yQUZLD0kh90amwTGfiPMW27RPfYd4UT8
zvbZiR0CGsUJbfpQWewGL2BsmjtmI2TkuJ8XaXpLNLfLmp0AQDTZbkO+colFt3BS
ew/l1x+W47/pEEvbQUDG++QHn1SDH5p3fshA1EO/J6l5hC4gmqY0q+z5ISC/TKxo
ORy4vjptXq6UxHjjcztYzw9c1QsUtb/YknhBaIYNKkRVpSgwCRrtgTL5+DFpTDp+
ywNbn/tpEjgY3Xmqs4nJeN17JLYnayeATL3pvbddrzKb2Atq2tn7nBk1czeCGjeK
yVvXQxx4/cM34bZjlzStAYpOd/3miRVLJRIzj1D52C6zYrpaOAgglR97JI0mRxeq
jQguYY8DBOw1/1lBnZpkcSh8hgGlNrvrYaZbJ6lDkOuxIUJR/uwgmi1aT2KW0ElR
LJNJbtXg2eIZjo8pggZdAz9PncGGLmbS/dxZwhnYJHpO7qLHjG+kSXTAffPShIel
ROvUXMjg6KMm7PZLaklCOagieKic/8uPquf1thx4cOuwDzoN+ex3xXCN5+jhC6ic
S6T6ZblDd9g0YgtEUVQI/+cELsmxY2gkq04a6rAolVv5Rh3e5FFeEzvmZHiENVge
KcK3dTzhUmNvhKFAAs2uYAHbbm5XMmoIMD9UhlRvXHkxzRM7DHig1Bopj8XVTpY6
XoBLGqntJl8ec2kUm/R4DhMYR0+rOvk/OgtV31X//K3I4HOGSM0FlVbtPJ5n61kv
dpbio4rtQ5q7rMa4VN+CpyZTJgKCKj0H5YkipkVvF2mDSQIVpTcuFDtrT0ElbfL0
BsCGFMmxq4+K8UIX2haUshkOzdD5G+Ir7TA33JFFMZ313tzN/GT3+vNMT5bnvO10
Ei1PRCW0wtQuLPaT+0q90z5PKQ/r4fS+iQ91i/p0NzhuWOC8ew+B9ItVrKzFAp6a
6N5N8OsVvYOSV9BjTSzsdg2QLETNA8frtkomOeWMUTZ9Io96tfT9ZSKGtmazmbNL
SANCB1YH17Ya9+3RFlZucL28L1P2AN9eibK1Hcn8+RJ43ldvcnbp0m9xhwFQRIDe
TqZVtAPj/2gT5MYnbTUtTO5P4532oexylBY4rGnv63+KWgZUTKRe0PeAbi13xhg7
+ZDqWdvHkJUQ9LnmdAjROum3oRJDCrLQ5hlPGuaN87OUqbEVPzojCXsT0JYpug0s
6kZDdClOyZIsMFyyZXLuNRxurKXi+pgnw52H67ITHfuqHgJX3adfrn2QevEp9grv
tOIHUBJ7hRC8BvUtB9SB3xXrVeqx/6iPDN8kr+BIG6kVa1R5J6aCCsc52BgZRJUD
VOkKTgDXrIVbdp+/qvi9c2oNYl9EJytImqpYGWEv8SVioMt1nAM0KKi36jv5MDkV
yEi/vfRQ/TuhTEqZ8tr5kvlZh+ZK2nSIp8y3irM08b+DXFR14VioaaVDk4xb/L/Q
eSzxANpfqJmVQ2fXOFEq0f2A/tX9gRucJWfnzik0hrUklM+k6V0nMZWmomxHnjID
Bbl8tBd0m5rPsGoNKIpa3mFVY/3l+rubBcephNi6bQK89huey+WKafUWge8Gc45x
mA03OhxM1ccIkNPf9y8JfR4Ei1UHYqLMG1AHgTf40+gRFI6swV5jfwdqkIvPi/A2
zArrkuD3nnbTKa7kmZBR5CsEsgPSJla/n64pfv+3mZWZH+xnt8iwr+rRe4KFAGtI
xWaez7yocHifkPz27zQ44WrOOzh/O9RB+h5WbrNdz/OmgCFrYXJ7xjNxSTH6Bbz6
Lpfnq927Y+rQpLfnDvjc8OPzQ4OTohDds324prc4OO+dKAEii5wIqlrUn31pIbsr
1dqpt+HEDRe1fmHkUhNByz6RS6hICL8y7Q7/usJ+gKdYTX2Rrp7aF9TMUw9Fcp0F
JIoHqkyhQ1APdjWng1BsvRMiMay9mZfn1Gg77U9uix3PLvh+4gXvmXueussMPBcH
znxuR8I/4VNVnjFzSiwCdpPN/FnFCC3H73AqjX3eNCNNJ/DkTpSfYeP94MedacqU
2r2UJkiAHTlzCI9XDGynNOXBZo9VT+XVR5CnWyn8ITP/IVAMesugbCNMnAS+HQks
St0vF2kOe698sIc0GJrka0WGD6q7l9pIw3uPbosk/Vy1zVdX4OVmPfz4swOuSmXt
uGPP1RxNESLuS1POWqRbSd64k3J61QtOLZ0OUOqsWjfyRsdgirMLaWjfojwBptz+
iVwZLzJJENMqbSikUlSNoMYDt1QHXNSQu+XnsYtQwyhLyUao+h2UmGjBbLkruykb
ml4z1f5WRyQY4B1WryQ7NTDDGbnJmBLA2qoITB93464GxO7vsmDLIEFz4gOH4woF
N88F1kzI6wpKR9sMpJ8vu53q6PAXp5qN8XH+FRb4Fjo2PtcRgCPLmWnyvzyxcHIL
X+ZaEm2269flBUZsNW/oNkAqeacdVpnJW5UH5VWeEBnF/49DLOmjIuDxCt/ny7wm
6Le284NeMWvQgdPkOmKh1QaCV2H9Lmlk2bN2hEvpzPExma96x2JxiqN6eyBPpRwJ
12vsyaouFCoZ41aQXsXCnSTkSZqSMO/IleA0iT/+LSWFIlP+SK6L363ZyZeQ6IFI
3OsEefNhEIHNIY2c+QJcx6yDDjZrxVYQXY0an9Aj5NWsAmJZLALhtrVrtLNX8zJK
+6uQ1w6INDHg633bJVa1o0oazxWMK/s86IRl7HKrapDkM9MzMZnnRIjUzFw0Tpzs
MLdJIaR3WUD03SGkC5N8+EQ6fkHWxuC+9ctplMVQC6GmI8kc9Bo5NPkxoOm6ia1V
6O35PdPFw0ZM3kh60MxPCFVvIXrQ7CbdTaDcSTxfTqmmMXCAJc5gyuquwsv+0Hb4
xcQl2Uhun2wAM2/6UGc1et+cMMLal35nQF2xOrXBBrBdfaQTJ4J5eOrE2wlct6se
XxqMJOaSLEbMxNkj+lCosJihQZYDJechWLsNceL9+1PSCC1Jf61QZt9yht2tFnqx
oHXgBLyM8KscnjpsRFKyuy8ToeM09MOpwd/z4yzT7OBwrr7YFNSHhuIWyXjBnl7R
gshy+xP2R6+yfvz6xBowvReHqLGBHvB0pA8yY9zt11MN8N0hFL53LuO9KAhWD83r
sfN2c3O2ZqoAMgQEcCP0gd4GkefjYjxQThYo4tlR2kY9F1wyP7XH+yPomzqie9iF
qBCfyn3wE1pyjm1AwZoB1d6Jzb3jI3Rs5ncmwIAzmAYjX6RRFl0magcxdAmlaFv6
5M6vkC5X3XnZBsfZ0RuaHyiWZnifHmU02nVrJgNXRXA7b39PvWwlyHIXxtnY3kRU
aqTEGCrnakN5gBhElR1ujw/qVnTswTNLO/xdrlXEHwEGKVjByAeEPyfW8uuit/GR
rZ057wJVpyxBia6jhxiTxPrszAjomQGz1wniryiX8xVXKJ1+vl1GKuSifKSuTJq/
7TLWsTS11NSAx1h3sO6s3MrApHm70yIx1fPbPAZ7q3BNCVZ2H8K1frQOmfNqeSC/
4wCizgnsKlhFS8Yqyy8zzK4ZfSJBPFOT0uwbmanzCiuuenKh6WHHkcUB2Oh9fD8k
wyHg4W0RI4IA45U3Na/u7VgFcMdeCZ/iJmxyYQXphJv1P0wbaxblEJTk5wl8hg0x
2VCj353Ca0n5Cx9UhpSI3q7G5SjTk8+DkRfbjK5LFPSNkzuHjA+NHbwdt1JnrnOf
iw94LZa9/7J6jXIZ+lSwdm/32SxUUsWgrT6I587Z5OE0hcDCfUm9WRr+CaX+/UIe
v2zJZKcgpduNWPaEofw7PWHL2kvlZ4qnfhoRZtxC8g7dwHBUoj/7kImAfOSTzwWW
aZpV8sAhTqAz8NhKZ9LjN3K21YGi6lflpfwh0OwWr4y4hyQ2EZ6S6quFRwJzAh7r
Tl7kPw61QNVbacnaa6x7enVA2Lj7WTMup3ZCzdDtIg3lSzkqVB8TQOOpeVRN5pAd
gj3IYObyZ3WP8GeG6W6rWsTzpC+EEAVcIf+fPGy9ReEoQNeavGGeLGRyucrZcJaD
CBAPP2sezG6kCpTew3JLgHhfh50jebgIFwq69XErwzQqAPOsaMuX2CSCXHWIdI/Y
18t6HY4z3oIQohH9Xh5+8wMcqXjE6bcbJuRxDneEAWnU+bqYFGtaX+VdmncN5KoT
C2lksp93n3lc4TF0UokXGVtg0zFQt98sKyxbWqnCKpK6QokRtnGx1gJX4Xx3Kqpk
mUHYKrT6+lyc3Zqj2XjAzI1f6OCoqG+yxpszb0FzbqfWCrDv1C/UNzakrn1zz2lY
xVNAZoeAnTLS+czlpH7BbWh5t8JLRytbctdaaDA/Q6HXgl0zXyjuHXqp425oLDqD
h4G0nk1uPozSLCwJGdFdrcf/ilalqgF+/x0CNXZRjOwexlzkvV/FmocOyhecetUR
i25hdp8/fXAYbS8MRMT4ex6C5C6iMKIN7lAniJQ+4zzjla9wx0/lKSNsaXAZKsVf
4OOljb2l3MZ/AO7OcXlrdC3iB3YHMXDzfNxpC1HHw3n+HQI90Wcqpn6s6nWUmUUy
jZKXhUYieNloFOzGwVJe7lmfNso9mPenr9nDbuYmQ54prxsUSEikZYFfZmXTUuZe
Hw2mvrNQqTS8KahpAdTO5X0IzMnu9DjfDi8ywuy07knjaVBcSLOfFVdmI+47cm3i
JzGBhsfSeAgFjf4XZ7iYao0G4d9U+F46+p5Tmo/awRQrbggrKvaKFAJd/D3f/XvJ
Urxbb4CMVrW0IHo7j/UrdMVLSDvsnWwN0CqVRtmRSntJ6oCfsg4xMnOUMdofYktp
pDI1Lzd2u8LmHee4ELpotki3npCimURXln9qctTRkW8Rt0VaXHyPRSui0ronc87L
K8iYrhfBoeYdvy5AwUUuNlkFpH/RNgbLYuMLeMI1dAOQr831s056qKog8jlm9nhA
q+wTHG/mOk7ZAkq+rXwnz9/D/cWERHvkJEy2xdv7NnTerMlivIxb5YIF9T5HT/w0
oe3jUmY535gvFG4y2K3WLtvWJw/3CG+hpOXIDlw6omC3fudTek7mV4J2cruYf0Sr
kQLMBp9M1KHDB+lTyHAeJIpGJAsrlsOEolYFE/rxwDdBPvSHd2PtXxKNON9BtVpo
IlFFp4DuLsJDf/KGnCLkEZAA6vsomHEuJOczm4XX22POnFopJusWJycg7Rfk3GBQ
hJrRZhpG34f64fsBpC8p+PIHp/AjfdTVIVS4lQ7t7GM1ce8vPtsr0hQVRlujMEZs
vHiqMdkqZGiJrx3jK2Bn+z11kUTqy+Ps/en3tXKuHCRyjeWZdssqqFJp2+1BmzY7
+9xtO3MacWLSb8CmopSpFnOKoo35/ilz8tNBKEyhQ6ts3rnoCX6JWIgGaC3cRzYH
8IDL0C0D21JMArxmkZLFfBC6haOUsfaUxVfTpuo1kweiTKBfeiG+GdiBCm3Es7JU
o5YgWlw9ypH7MehZs92ctvOS4+tzRRVsUiA5u0IKE4TBPPCRNYhtP6dT4Fshx650
gXPIMQILCxKVlTVz0hgMpF3Ty5JuLHtbNqdbabj3yYel+5xzFgVMkamORzA/upEU
/FbUFOKwNoGr5Ks9oxhYQ4q8XppMgaBbhBmOYRlBDptfeIVlSV8f0gxdLAQZ4OeG
nkJXAZ8uuxdaPEb1JPuk/8l3bBOaVbyhwei8DCFC0aMoEmBrhi2Pb8iM+Bb2EJJ5
FUxK+CMzmv9fvgLLqiVbUA2vYgbhegUWCmYtgGzoPv3m5ewxVVbj5KoqIg24BpAt
YsLrq9Y93FgG23PJh3+mDV88yK9DeuHnttPTMzzuBwHzrJ+O6q7ugoY2ZeungK7M
YJpL5x5YBulppLGj6bCO8Oew7TfyU/91S/NDPlAdSuNTscDtK7p3CZUKf2vCxMDL
TOmsddJ5hQxWYO3kX4q0gtPJ3S1WlVxeJ7CwJk6rGtTgaW+oOcYNSTu7nkGEI9pk
DLLOX/2R0sFIM3IB0hBmOWgqgeKblc5c6FbtheDI5DsqS9Yw0tjs2YnQOmG72G48
w083fsIcprKEF6PobaG+fFDs7c04plv6Muws3p1kHH2NLxeD6XNOBnjQrwWN8Tc1
Tomr2KFNV1qXavHYK4vB9JnAcqTIfKjqVKrcGaH2wjSGlF6x2RL7laNCvsN5lYLZ
w60fW+MRg6rlasvUCWjZ4L8n7C4LO1pTcW0Y4hPSNDFNbP8fv3E2K3WMfvmHHIAr
kfclpeYSKKPsI6EHT7mZELLXBYSFiyavQROKcBbTMGEX87caTzoUECv3H044Jm7t
fLosEWD1lnVKBhgKXJbsVgU+oCpy6B3Rha58IXh7hUIUdNFLvnqiPStcYYIXC+LX
jOQtHQBB+GtANRALH4wSudf4P7UXzl3UsKwhhT6+RVfIxfuHJ3yh8Mbmgy7vQLxs
IlI02xhVbFIcQGh2e3R3YtmgmmfJ3UO3OpZWZBqV2YQ2blhmzaZPA8KIyjsC7V+x
lTqPfR3dsiDLKl1Ib6Mr+va1nc1moP7AaM5QQ6luGZyTWukVLYyw999qw+oZTbAA
o8fX/njIMwsyJ2PSP721yThg71iECiPTII6KK0Ze4djg5o70ZBAN3zilgS0LB1d/
wGkvSY8DVA3akdScUCBDaQpeJEOMDTFlld8il7DcvNOk4v1mTkWNG67w6Pk5XJzx
CyXAG0qErWAINLdb83iKmLrPBEpNac5P3X/oIIYVlQc8X9RwJewRw/mT+VfbYF1+
jRGpUVoxFxM7Oy6CWVNKyEcb8rh1hVx9cUMpE4Nwsc+yNHPz5YABVKTb3DTdHGQh
d9CX9R/AYDYOWLEKtSnszq2/0XbOLkv35XnCuREqrTsF7w1LfBAdKUq5x+Dq8gQw
LIiDS8KBLBal2qLbRrONG9w3bftb78eJ7WiOs+UTtRZrLNcEXD8GwVgbGYFTmM0u
wSoKQXvpfo12e4R8k+FXQrKhswsMGpP4sgMso9E07gV0a0PJe3zqMeEnFufkyjMt
l4rIzc6eFtK3TLhSakrZ572hZcDZSsX6FInrH5Um6+FBFDJ2Sh0kP++kndVP+7Hk
UIuMMI0tGzgHMGkI8VpW7Hipvtn3vbQJvTabEPyVKIb6i/faNodm5n/BfdugdyeM
lNxGk2p6r08mbTZ12w3ZGh18BxRYWC+ezGKbt1c0b7Vv8fk3Lw1qPvQQ7rvV2tiq
LJsAboBcuJ8wNopgaqEdY+9NLW7woFGqNUa7JDgCEVgthzD8kgIRK9/ZBdYSJAPZ
CJDGr7JlWIa+DBHr7v+55ZpOuf/RMaree+t+m5U9ZYjJp7AjQn0igX10cCJMie5/
WBYbMngj/3IT1x59uG6ZTcV2m5CoGeTMEmIWZU7OBBpQyGZMzmDJ7+rQGbQLnEwm
FgEMBBtS6O7CPTwoTLTKoQHrNyVpcGBEltCPVyxDK/F/x+jAeLuXJCg2hp/6Img7
HyvRczBk+p9NOA/DCo1ZYLSjyi2i2x0aYg7iV6On0D0JlFagZrrjUcH3Xk2h+QxV
6kXXR+5bBlk3X1IGs8lY25eQEtbdPC8vKvzpXFO6u0MqoXDd4O5Fy9tFrt0ijsOv
mbuxPNIzOK8v7wCSiHVl2Ks1HZhs4NpbJr35jObrimr56PVLxnsKutMWkqM9Asc0
uixfKdXBJrz4rt5VB4oLluysH4T/Q4ELjzEIMhYiD/T7Bcb60fKMC4CJgtfSG/pB
Ak7I+yEfXecxhRcBu4SW3KH36Ly+Sk0SKt/aktd0N/s8MO+6fdbUGaptLi1qxGJ1
kWRv7wBEHab/nJLA7zob9imEu73lvF0OzwG+7f4tBvztVjznznDVV86iwdqATVSd
M+SFyfDeI+53x5wKOyl96fpVzKOdVCM51e4UxgJNeQ17YebuAuEGCjCovWSfVEb2
eor2uNsoL8Cwq2zkGEsGFXG+Za/eA64l3SB6LV2h1LGjcrbFpjbYDfCZjMmup8ir
N+NUaxD2NguJDrOlxy1j7ZYqzx5jtlG1Sy+UKlKl002Su6Cy4dU/cZoypAJHvFPB
KuHKtpsS+93zvYM6xyNAS5bD6pSI8sVKQ7Rc6ZXV1+SUpgpDcYaH6g0YFymnq/ps
JXwGv79Vm9fU545forJsJBsZCi4RZSPVG2JnqBVqNCm8rSoGSv9/IeGN7UtP7Nr8
wV6wvG6hQAxDcJAfYkPFAC+b8wsjcCJyuhy0JL4yeMHC5BvH7YFESY++z/DxBUcf
1FsFIeFF6fJekfbuoaSfvMvRzN2FV2CxgO0rMS0e7awiI6Cgs3JduhjZa1unUtl+
FvmgmzZ+pMPRSdcz+afzHRPDdJTfBanzP9+y//Zofj7o9MnTy/X7jYjKCpS6Jhrx
JVfqvk2Jen29s97OIkIjrDOu/rIdbtQdZbey8Plf05+mL3OLaUrREOjg+lW2A/0Z
hwteRTdy6i75lXzp9pZuxZkSHnyWqbmd/udceyFArb+OKGFtGrSgIdKgYz40r/YA
ywdL3oQpQQZFs8EScjrOWRExyiuO+Tw+mFIfygHneYpfLEabKs6rg10UFGRWaPne
hF58K2EUbsdmCuiQ+DmJcYTkXPkyITjuXI8pR4tU2J37ibsuN0HWlgEmNUsA1gsU
AQhwXtN/nRFHFOcGpmokDxIYPcF4gX+n6DCysjaWHy1twN8akQCUR+hPGFY+83b4
tSGUymSCAHVgUlRj9/gKawpgA6DFrBe6sZwMW6b6Xxsd5l50LNzJzeGOTcsSXdFt
pRRA5Vb78ZjzKP6gNSjuRWh31chdk0qubZU7hJY46ohgyjJ/OSMnT+cWixBv61GZ
s+Yr31h5S7nPPMr7bhaXY9W2zlY0pQZv5Z98Se2rlBvkRvsKuS1zWLBFY/CLkUdv
y2KZNbR6QHgvBRRceVcBj13VQS4f2Qx4x7u23a+ZhOKUeXchhRTqkr0jiBc/pAG7
BuhamoSOpkNHQyC5aPRHJfyv4RUg+3yy7rDllA4T7+LMSTfFcNgaEypvXABNBY1O
AZL0ffDppIjpUDx+4FiD2lHdK4Aozmrq2eJq+Qt2uk4dS26JdLmS27mR5MzXfsnZ
3MOmaLs7hrateu0hdLXGCbTbWpVhO7o1/u8vNJAQWEdppomrRrBJICf9dGFDsBYk
X3aYdePhxBDDfa6Jv79TZHPllstopaz/Hm+q0ZHzySSSp6hTtv7yCPs3x2stHO36
TsHYASartQxhe8UQ5/n5t4v+kvKlo33jO6gWyld/ADaXUFaLj7nDFkAPIOoAK49c
0ovks9SiJRdN/bGiLcJ9Srh3xpZ2w8DQSQm5mhhTU+6zDdWmeX+1QEv317Kcd42X
9bv3qbVph2jaGpOFKS4nxY36cgbsjAKafpAGKJRuczI7ThMBaFjhhxz5GV+7m59c
d1cgYcvA8H3OiRYXUXVITYJuqDIIkkBLmKDTuQmDNFU6goeguc9kLachft/gDtPV
tkDBX7dwgeM7Q+Pj6zLQVMWEaWe3jBitHlminqyyLKx9ZGcJRjG9y22nrzPpWM0C
3/N53EGoPkYNXogKb9XZZ7n8BIK36M4B++wjdIvVXDKJmgMVqYkQRNJsnCE2dGON
SdUvlX/CexPDEiwwxbh4lNilKhsA2PFvdPlVzrJ5s7DBUAaFBM6OzdrgTctkdVmV
vOGpdIl2pBOwhOP3O7z3vVA7HcsjjnEwXia7gox9Pcnf5OIzWjpn9NpzE+SEtJx3
njDgLZttdDx63zaEzElycj9Bh4m1nlJIlYRMq1vsTOm6/njwSYponbBiLKDkXGiA
KCXHSqM60GdjVID9iQMt1zlM7dqVmhfu8t1tmRHIHopBSYO9KS4Y7HIbUj5ZZOqx
5MHfdnmiFJEWMRZxRSR98sG/V1ihL9eN7P7OH3LxMF2P9qhLvO36RHYJJOujZgQM
x8IbXNj1DpUbPaVOdcgRqXPqyCuICQNMrsOyxOcr7vjp2dw5I2HM5fE9fcvz6rII
K4UBpGwNxSscV0KEKdTyfJaP/w3EfTldDOGGFRqwO6aE5dxnt7NtI1uRKJ4hw6cj
eVtm/reDGKYiPKH9xjisx3xhPFDiVFbSyzw7WW6PqHlX2tcJwIljyFtk6NgZWMvb
0JpXjcKFC8RChJIrL1lPCpTeVPGn6i2tS0vnd2nwrB92eS7cX6IHz1CJ/RdxdWUx
UzZCkLuQCeDimq6XFmOXF/4cVJvl9Hg0bM01S8FjHNagU4ZZyqLxjRHTWvwfxU0e
SxlzROVoQsazYeT0RbsNQ0S4MTEQ5mhmncKj3GQI8Lp48SmP/LuVg/ZhFFvTLVdd
dWfVZ/++EY5mFy1t1dgXRWmWChrgfAF1hvTuJPdaL8Q5s1hSgSgwHdjkXwK/MRCc
XbGeofjhblzFjHykExEog15cBPSFLhPASGJDY+xAcvpYSOVTVJ70K5XkEZ8E/oP7
KPiStXB0z8dHvi9hUw6fCVW4U/ydXHejvPugU02wtoskpdqFakzZ20GOsnQ02FcN
RaMLvnU7ThjnZw3ksyxA2enMWTbJy1iLac/By2JWiFbTgjxgAzdm3suTAvuU9AEX
TAy5MBFyC9hkpLE8VLwU5Oc4O2LSrOeCWvT36yUySolcgyPnNK1M0jgi5Z45NCaz
o1P5L+GI9jgbv+dLs5eosEClc3vCoSxizgphbaMKN6yY2zh4TKvMwyi05PDb98EX
BvUwAoiv/n0g83YE0RzLgr9xECr2AF2naV75FPxjj9cnViJwQN2GR0l4uD16bhsh
6lkwAkKT/cc5eWl/4KsIQOefkv/f7drhInBC1WbZZUptzjTeGBEz+YHd9jlflpzF
5PxBQ0iTCXZZJXoheCXtr+gm8yvcYZA27oDGCVp9w588PU60FYjaXmg9ZQVYYP14
yncqguaqbfdZ1nw8JRn+c4iwS9voXD7Pa8Be/rnb3sbHuTCGyaZuj+ObnE5sxlyH
tSiMQulOC59P45jRfImt6v1JUy0csTc+kpTN6kN2u3feuXF2apAgC4CoRmJogspH
hMhB6/9HPf4/SPTcztaIDDgOmUltxjg8fFDS4isvvWnzeerYdT/i0yGlPaW/ySsV
+zsIzlRN55oNEo4LlcVIk3QHAC6sDMDwbknE5SwQPhD/aQqtPDnkSfYxAL4mGZyu
wcI5QF3xnwbrpQeGzGDYFtzP8ZKe3Qup55G/bW8C0Z/bljJeQwffWYr7RUlmLTFk
TRpeNAFWiZfPgVBH4T5O6yJbWvlE6XI7kdNL0r/G+pOCCrhg0QZqaJKdznFJbiKQ
5iHvURkAcKIGC2VpDMW5hOj819L+hNkGkKaLJEjMk1mWI+m4PRDvCasN8+FhPmje
SLJjMVGo+96wz1L3EZj2GjqlwQcm/84CMDKhhgeXGDqAqelLVoiHPM+3Ozwv3czh
MhBXPR8Ql/qziJKXsVf2pGN2PER3nxGER5h3rFiLjO7oHBM4yCC0ej01MblBBh++
jY/orHUlhMT7CnWKw3wjY4paQ2w8NhKMhH62gJDxEH0WTCBks2LIu/evoCGPxRlg
Fqd69f1B8My9ES+XUzDoM9SlJkidvii3rUdMxthZf+CeNLssiKiwLXuBJttQiGYS
BlI41qQSIhemwTMHrlJzFiBBReBoPNyzfnrYXSE4mpuQy22zz9UyMAUrBO2cBAJz
yua/F6mLrTrJMVTswekMJAnf4nWGWmMWE7MDOGm+mAdnqfBgo4DYOuE5me3feabp
6V/SeHl2Fn/D7wMlxHsP/sSH9M95tBmNYDzdX5vF1SKe6JCEsZInoVsiR0f+xagY
2GnxXAy804y1lvc+F9isWaeN0L5sjFtHTdZpf0VtNQGhiP1C+KOjtfb8EJGKJRth
mVe+XMhL8xmxV7aMUFdNjzPRamQg7+MDNoHTdLeacU3yK0bb4D4g4OQGWHRBXtDK
ljxwbuGD2Zrl3n9EksdFdxoL1HIqpJ/NxrE+oeVOJlujNDcbVVyotE71k3khHoK/
cqlvdALYUVhl9byZY3yJ35+5amLBhUiPonuC324rsOJBADR7ZUPlvrsog1o0HrZI
tn9+rYWTmAxWavEzNwSEyon8L+1jLN+By5BmqGsQLjPPGX3bjTuGgJk5nQBwkT9A
DURPelzeYPDyO0E2K6rdsS47UdaXe26X2KUE9Cy99eioOpJ/hrQnLWVaGw0ZvgDc
09tOBxpZDtf7eK2HdHBJ93AFluy/ak6etOsXu5XyWHMGSwMACGigi/KE30+5MnyH
YQsE22dwi83YL2X40wleAx5JuBGhXmLRKeMtwb7KJkFFZ0CH43RFllcw3T+qTrUN
591aCP/tvNvoF3QLpBcgqNJ4J/zyRBA6hvDx/2dNNbjpN+04neV6MnwVAZ3gBk1t
JRHLD3x1qlRgbPQjvjI+uek/t4/L+H62U4NKW3LdsBM45o416GxVJnDRl6zJ26d0
+SXs9a7seqYbsxH1xiRP72NHgMSL4Lywgih7sclxvPWmZNw2TzYE5Vci/SIQvwei
MROWalLiLRedQpvucOv5gb8aEi7KCWOyE71RbfvsE2/DQMF/jpstdiPmI5Fos4uZ
QxVRMWHSgef0+iA4Ae4NZfs3T1cP/STBqeFk0WLBqItK1yy8ckyQb1cMVCGFVKP+
rIihZS/78tGaQO/uJucDX/LsPnWA+neBporbg2H95DFXeAaXFr0DI0k9I/Prygf6
u64+SL0Xcgez0/L2NG8i/AFvCLY4ay/juH/k5U5L04ySzkQSYxBZg1QaAC8I7Tg+
CReP2j8C2Tku/of+TbebFRoj8BZTSa6yt4szwBkjwwcdAcjph/Pp0DMOX9N4EV/y
TdPkl4aWRArSpuSnrkhOOqplHBCzcDYffD9Upb+oCxlNhj9+Nx3AZPWCqt2qKwbH
lX8GO/IoP4kcwEel0T0CE956wViBRbCenR7anHIlPiz29bkiobq5ZQZShEWTQ1hX
+9SJBwT1dqrwMeNKMQ3Ch/eH730ikRnJ1FHER+T/4rlNJjneBetHLhauMm1KYilc
KxDudcRDtYyIS/liegw5ndEpncRJCemlsY6pld3SYHBKct2hHa0PNPhizi4MCnse
v9iHPLsf7dbO8Qcs10bszRcShH1WumRGlkyxAIDVBV9RM7/Il/DxDAvqJZjDYuvy
vgqQ8tWS0E/x2BMSSHUfIul5aqb3dERFIThTkC708WnbXm5LJLokEvR7Owg9Azwu
wfZt0uvk5av6KsebSFxMmBFe+yQgUes1Sg2whypkGQKOuBzrcgXvPTwodUbRdbu2
mYljGVxmYOdbtdepLOW6NIsOGSt4YD2jslLRslplBUnypQO8TpgnvZHX+Zbr4FRu
CEZ0HRkyBziixisshCuVLADKdHYPlabeTC4NwmYb9fZpgZVg705Uj3EFjZhHCk5f
1plzJ31669A3V35xrHZ3PSBNoYD+/NQZpVwOAhysct/S5KEmtrvpB5Fu+AgnTrkT
y3mr4LGM1EXGDJVGRJSsl6JPr2TXc+IgZXgZ4ONYODVrfBcx/Prm+fdRXWWztFtX
q0bkRAWRgakCInUGIlV3Sd2Wnlj+w4Nx1hcb91BtwDcoU6+yy7tQ88nvL+FxJc7l
YEjJyNePkfjVpwjc6td7jKgGTc9MeEDwGGtwQJIxkNwmNbyk9k3Jfej2YAE35QUu
Iqssdk8iLrXz6PtC0ee/HxYWOGG27GlR0evz9i9y5MpgRcI756Yf8mjgOBb4K086
bdsOhIsDX3CKJf30naVUwPHw6xuVGtL143WeZg/Omv+YWH/C0i83ySQwitq1n5Sa
HLA9+Z7Jr1MNYlu9nLtRHWYaHllYRLRrSVe0mpp27zz4p/TkNFEFgwiuwbtVFi2x
CMvjQYVXW6gY7PIkUpjZyZHoyq72dwIby5MegX1BfxkYXG36DmLmOoTRHPFdXl9t
vBb693kr/lnNj/F5eULiLZ3u/Zd4vzSThwbmHjuFD0hvPqN/VO4hGiUVovB7hRxM
k7xoB+cBMuf0wo7l5GiJ72zFAtkSk2S0nPBRI0ztNnKfBzhrTyevc6SfpvAWN23R
Z76BAxca8Yc4UBSz0j8V5Dl1YTZgk3/Rn+na0hqk4iWwidjlHoHx9BjEGgmSZPR3
tgHkTFSGwAnwd2ZqjYuhmxS6uRbSh7d2a/RwvyB1Ro1yQ/OhNHHRiRkk31XfMshQ
6iKhgEqIPejcPDVIXyVbxBU+hXdyRMxM9eVyQ8ZFyQVyM+4voLYYZ0+pbSrsZn6C
GH1xtb9GIleCIJR+zlbVklg6/uYEbreFlfeNnaXnQS7GWLc77+crMI1ezkqYSP3P
TCbp0++OlJMu3Cgt2fXd7NitPPiIHIZpUyGwUsLnAXC/fKNe5q4GfoseyMJz1/a1
+N4Qd7B14MaigaikeV7L13Srzo5Vuhz0tIG2NuGtvL46KXrISRW7AtEgxpbUuT9w
ANk3BeV5xE8CxXvlZtNH0TIcPNIwJSm92ZWgeuAYDn+h3IAuy0V0t7ZRppL+QLvH
knsjt+HIrslVhxZ9M/owcpdwA8BXXB9vgSVk0GTIDEQ2m4J1HGIUzYBhQ38x3J9g
QRr/+a+uq/pU7Y5dCC8m/ww6OGJv/PWJc67Qreyk6CzYTjvKcRvcz9s5WwLGG7bj
3+qQW6mfqNuzmfg31jTqQSvP0RJA6w1+1pwr5wTfY1L54ioUUwnety4AFlV7JXcS
ei/0tGcpq1fVE1TMiMItvcaHjCyvyjGS4qeP0GzhRIgGnNMegGM7UsUAkzNXNtpV
rLgYxfo6jrYCvwwENmQqhMc3GqCdNYGU3F8mO2903NNXujoYNpQVxjl8jdNxw//Q
GbCOqKBgpf5iBhDNPUc2vD+cGmX+oQkfQisQu+gk/EMqfyAy5rhpJJPDmm8R3yBf
BSEWy7A79FIVD1tTqN6Yws9ecZXEbMUpbSqphDQZGB2FzW2J0PI3y6f3TiNBeuh0
SgTiDi78slyQmkQN2/TvQjyioW5cPDsNDLv2ZscUPcZuYZ3IRp1G7pcuCvn41zA2
LDwU3o4THNjlkK1IceO7hzmNYwkyfdzq9eot4jKMF4Jv7iEg6fistoeq07doOIHZ
DANzOFAUEvQqnp4qZ9pQxG3UvLkGiAjJ+3I2q5W/B5tQrBIOa622TwC3/lpi5Tw7
y78eviJ9q1Ck5VBld9xFaXrbFO/7KLMdyo0n2vzxE/8dk5hDEv8PNB11wLSL0YnG
qtMc/IEwPYUpp0USiAhRdLtB+DnWS74kYuEF+BirdkqQX3S0Bkeizm3lGbBKvkHV
UjEM9QjJM8t+nKOGl+9/zSaNfbEe64krpfSFxQXkvJ9zSsTN4u8DhRqfT6215Igt
zvJEeQwWK2oDS0jvNRftD78Rw+I5hV1H1aTpq7VkJX43f/KwGyjmouh17khKLhpL
ueRf6bhgWWi4jKrZZugYoKJZJoHR+lbExueq2hyWnf9PLWzLgA8xV54Z4jW4QyFx
s2sv0yaqYnCdHEAHK26lbqr3bqHOpSpBUk1ge/NwJroDIiO7bPOHFCFujX15qRV4
6eL8O+3UREQaiklTnIWRoaHmep2CG886uan4BkkzYQBRQPNza8oVKqE62cSMUVTh
Pnfafs9vrkhLo6ex5HfjxCJ9ei68NlBINaOfP0R1D6ZKX7+1BqwgNKZDJYS7PBJI
uBicMTTLYH01NCScSrxc7C0YlzXhKCLDK97+36Jqa4t2E1Re9nnuXkI+qu+Y2Lhd
/LRM7hi4iK2vK2IZzBA7kMPH0i6AzFzDd4qLcIT7JC2bg7F1rku3tYglyytntOaR
Lz59WRw+s9uibWKODtFRSfkOtqeh4dZw8okah1kPRNDJ2UlPvrngIZYFYTyZH6cB
KkWb4996IjL9bKrZW4MzI3s1H8x+qb/xzTeYB2FYI87XcLeMqF76P+Jm47fgqXfT
cBsH3zclCrz7dDAqlE6tr0xU+nUnVxy7Kni7VtXhpDanRvroWSs5g8PhiQWi0JQx
P0TODnQVFty2yTU5UhmYreytvluiOzs8QHBHCV64sYpWtuf7P/O8KRKFhLNC3NIp
6kh+4KlvpwaCji+WBB58ZcJddxR0ygy6BYlpwdVtHV9GAxTAiOrP+tIxeJjICzbH
MhQKeN9oUyM4+slLBzAlS3iK8mUiP7NV5qkoneh2KEVlyYtdjDW2TImprdOvik92
NsqMe8Bo5/v3xChmiv0Tdszu89hSkDTfQMYy2l6H7Le77080ATA8K8pzBJjyl1Ll
xSJvTeVQYGTafyrWqv5hafUIxqNU5xfMSTVQI5ew4/5CoKk4ZfAkYUhH5igrVUFe
lmCYA66b0DWW3c2C4iqRqizC2NX46AEigDd4zvawBFNFSJnt1/fC6WEANDSPM/k4
T3QowgW7Cw6HFntKEcfAwLfQCacBH/dUntJ/gE2/bJMtI5fxhSR/qEEP8HSx9Tbx
gMIkr24TE0VSZqY856gD/9o3nXuDiX40tbAJANMoqTg/qDA2+01Rra76n4P+a++R
Vt8FlvGTp2ngDnvu0/7TzsG6e/QApefaLLzvJne+Ew/MpvHzLImJjtaDJgGpaPpE
oRA6/2KYxIMzZSARsfrxdISHRucq4vburFSsFJ+j8gTZY49o9OSEX3BFd13c3VzS
Oy3KNXFnjt6M93xuxfKLFJs0iHaQA9d7Zbtk+Po+MfGeDCcr/QpjZnNtGwMAjOUZ
DnVSrNPa1nsttWBMZAi0Z1qZxY1saYZJYIeu5A/tdfqGhkwvitJGidQ6DeX8Quq4
YA4Wo51zjELPaFN9NMR1/hsB1ua55QyuayyZW3ejzZFFTr1z8EiHbE8lxpz7Y/ly
H8CdhM0dH/Ovs9GFt3Nq2MgGdwBAWbv8ZR/O+Tb5AdzlBJGeYrLNPw+u5EGCEuYw
fbkgxiGBkMiLj2pmTejm4Xz5T6vZ+pbw8tH5PfKDNNdhLakZz3P8ofs34QHswWRg
Td5rABoZLe/SQ7ptHBV/bs+FD1kQQ1UE1h0vlEE3m5SJwAGyE8SFyMeuIGMPeGQk
Lobnxq9zNt4UpYhT81/Lk/kiv+YD1glCi/+7tAvlX2xVP282+q/60J4/6/byoG+n
cu92ruIgBrnrb8EE76XSrMvPl0+7lEuIDdzNZFFvltGlWncCL/IYquWGxAfDjw3J
iwtEWRbvcOw5ZJdQqreqtyik933nqd+KRn5oJ+75B8lfvvnmdjO4N/KnVG8cnNvs
OCgTOTvBhvQ5qw1XAuVvlayEbmpxNBOX0LIbG5xwHlF6erpfNl9uPu+keLXGon4D
7/Gffz6SW3rWQhtL2/JA3cLGWBKnspKUybyJyVRwNe20kb6AFguI9WmimYWvqHGI
RXXUvDbV8W1ylVYFoxD061OBm9N8gF/5/PZ2Gq9NhOx5kiDCHea/vszCG/0V7NZS
6Il5N8BOFyO0Z+b197YWjfVuMUjd5ei+0ZYmtkh6wBhrNW8Lhqvq55J/VU2SAU2O
MrWJh1ujUQFYFO5nUjJSsVx0hqVl++OuZqsg+pKsBGf+MC9FtwVkvC3NAkUUIG49
LJNScdO9Wjbi7xWv9B7kTMSaTA1oi5DMXW/g13emhyNCnVshaU5joavrDPA3lEQw
u9/8o7okPb20oDUrT56v/6QrmLQmGx8k5byvbI2uFeNBdY8rOn0lU+ccil2Vf1S/
2shpTQ2UIixnrBYAf7NFo3dDHjdAtlU09uAneUkXl7WCGM84O3mIpsqcuAazqbu8
vVGhV0TBWl+JiCY+jHX+yi81O+uGMgyL0MuEk/NaenE0wo3bwKuZT3vTB6ZnAVI5
oatJukyk2Az+NIEYELR3WptUa6ZrymM1kMPJ/bIow3at4qhAFypaOU35YOObGp0u
kA9BXzYepxaHTDjYcONNpk8pDT0fP33h9RA4du4ctyKAhQmZVfsqe/TsXM7zXF9g
46unixm7V0wtxDqsojwTXCpdJvCYVOXyz6OxW4D+sapqCaYbuKgZ0OuzkntXt818
AJpYIeDhq0qtC8hq1lvzYNWQvXjpaIK7EO1WXbNt2ibmE9a1pCqxCqWDxr2Qs5ka
e+XquLGp3/kcNI0uaQk1r5gVVT14GHFsisDlwSZaGIvCeKEyvY77Id9+phAW1rDY
SuT9JOvRegx5yBe3bndDlSj9S+u+4s9wFd5mJA2opgBt9KZ/GMD/Mg1BwN07N8Uf
hzf5SkwcYgU39Boyr+s8YGBqBKE4N6udUZmpBNWD7VzfT6QzSXHmVARTwvcc+NwY
KMsOwSmVlCJqBMWcmOdp02Zv/yqc7z/E7qyT4IxgCmOU3eIbaB+7hq4stFNynCka
Pzh3QuA8alGbAi3DwoPs+s1bNPpOxIkGh73cmUhhB9bCG/OMzdAKC45W91DcfBo1
Ss3ZLdUYvatSmz/xClG97hVnEuR0+AFaf9CZMSv7rV9UO1/ZtW5nlhFM+A/NwntN
35Y2xx8O+cEVKewZO1FYDJPjp189kM9DWsOzx4ZTiFjzTthJq5LVTb/h0DVRNgj7
xxctMJ0Ye+6VZXH8ywWgyUYJSFcAeeIE2XN1NMU0Yd9ldPAFTspihnPWlYlJSWgH
IqYDvFRoyhsic7ZTNKjH2LW4jlIy4cRZML5aUbg63R4LYMEnkprpCdTakjegHS6F
3i9Z6aZlIabghTDVZSKwbrlQqLu+hujbGViA6qIyslfLgUMGyLyJdW/LZIHzYT81
IFuWgUh178VwLLE1h5Yx/eRmshxW+0iaRXgXgi8Lh6DnSunlD0GCE0ZpR9S2sieU
ELfMYlShExsHm7cOZI0LndkQQzbPUTAXQd0Mm/tDHh4d/P/ViBbzkwBso3CvMA6o
dseJ2K/v2SLcnpOXtip1Rp84lp/99uOrlbEN/2a34VdqoSQ3hrPkVVHthdS5YUWl
jhrijOMpA8iTibUuaovkMV7F27fGB6U47sm5wmM3vDz2PW3601Ph5YXXVkvafmVw
0TD1mOtF3x5UYTjC4EBCZuPSVE1OfuzMAgBO3hBVIz15mnohmjKQmzz2TDldKQn/
msfboQr75UFeaFkaFI2LBN8bSioJ4RBYxFLd4pCPcKvF9n2z/+6O/NxsA/Sqlsml
XjZnO/erAmQi/L0tla5qoH+0ByQ2HxUbuikJwf9nsmZmo77DuBPapUAPVG3QL+rY
OV2FF7EaBMbse8mnIlrw3U/sEyhp5ZuoWEuI+tWfKPCNShVlK2CwOdP9B9XOVzmN
g+re1cNbyPkyhTWVgn7pvzhYoZ7eiZKiFkUxsXAZfEgjY+4XchTKCaBUyQpb3/e4
nXTSC5A7wRwOFsJDEEk3tGFwT/ZXd+QSUhejoyTkNpF4xhXwfyJYtv36E28Ba1an
2SJHXYbdONEvafyW9bw9yN1E1ofSQhaOgk1XYLUmlaAxU+naF/CD+eYPmY+BFjAM
u8+oklM7HP8PsMVMvWQcYgQLhSNuFXyMr0OPWePPqGcHzMBKhXc7RPuUMKDkWN+W
JSq0wsc1BZFc20KJGh0SYx2Ol0X5GOl5xzDyBPbRJJt4Q5OrL/o1nVNklELVaEx1
KHy7fXlXTXxICvPiFjC6PCCnROxIKkiTerR9Hk66+Wj7TM62SFpCy8C5H5nLjg4K
CUgF1LoV2S18fy7PDLyfk3G6cHPPe6SFZ6EitMMyMs7mi04WNxTFoBMK3LQEfZlE
0+qUn+6LaNmIrYOtIRHh+NMSZNE9VNtNSUm3uqK+Dh+yD2Hexs0IkaYxVQLqpjsI
BTUl+VQ2uBrav7N2hs40DBVOK/VFL6kAn6cStNB0dVOS7z+YxxtDN4THgMmJYcOZ
B+cwDe6tAs2QzkoepCEuD/NzNq9c7LN5hbXju5/0qQguQESgaHHlcGuTzGg2A/0B
Pe+zSoFwjMrO1Rgju+iocDo8KIZ/DugoslYR5p9yiCUOmQ+QgetBkgDUI41DP0gv
epTgig0UWn4WJ+3AWfCyEcQi9xHisobByUQVUKJneNoJ+GLziO2W6RoPM1kDddvZ
O/ctgfiesoKpg08JN62ors5lUTQt8sx285m1fIhoTgye6J2HZhyrdzwfgabOVFuq
mlS/HvS8h5SZ1JLuVSjwp6rkqgCcuq8pgVIvnzhijmM2til+W+9W3hciHHc8POjU
GHGwuKH8Chx8pvGjsZdMdAyh+EqNW4O5Vch77pAQ42Vg1AjnxuYM0w/SukUcyMQj
8O0VZypj++zlbh+RYsTOZT/vS04arhNPTn9fG6hz/nm+JIjRPE9GTUG4MNZpBEtm
T0XGg8xwEGVyljo35Xc6bYopauWf/WKXOdZA2HKsqwDMJDzx5Sh5EWynh3Lkzq75
eegr+fUqBOwVTSQBygcFuFkGzCSltkm0yHzgxfdlep/z50lUtqKfP1K4s1KrsTSX
ixNApa3F+XtKyWiQP7UkNhZWCSOYgHVWz+UlfHHRQVxOC8t5GkuJ3ZCRLqqeeRc8
sopxV3QblvnpSn2crQqGMehk6iMkr/FJLjiI2Xk0vMcAhXznRoRUPDEx5ILFXGk4
HVCYRtJwgAkLqP52Jjr2FpqfoW3g3rKOzG5inO14enZlBmiG8mYlY7wXP6ZDN0h8
WDKbS7kYrPe8GSJS+Vf9OmtTquH3e0IlEcIk4qKbAZ8u4UHGTWKXpe8HqEG6OkHu
EbZoFFi2GEpO4xO5sXUpcBfI3l/32tDanEAmxJw2omtZUsv93uHregK6sz8yDaJE
+LeRzHoBFDLvABbvvVEUn5YKeR8NFEwj5KXzhGIAiw400HCMdQVNAAHpP4+Kf01e
6uo7RF7XUrHFVpZBUd5QfhnbOqkyjOul1zJukgq/g1XhmoUavmzs8W/nScYMCKJz
m9m1TkijrXPBFG4L+u7KuH1IbtMVJcYJp3Up+XaT9aC5J0LwQPuVnSJuGgOSxWzx
ie5idNuj6gy8qFgYQBrNdHFQSZwaQMVpzar6yjawpM+tHrAIa+52oFJgPNzELUZc
iRr5KVqzU5jM85lJDyCGGGQI517P5Tw7Tbnp3A6waeEEele4VlMEbXymURW1OHq1
m+oCRE1HTGXOQfdk/vdoOiDJ6jrZVJe7PBzM4G1lzIcEG1ZG4tNt+vM6n0odS3Iq
OvSbHSdMYNCcArK98CjPsu41tKEwr1yWwVfIXCA6d/EK3mOpwoGizinnBOJlbTHC
wKaMIky8OYEUCaqSmDBd/waa5O2kld2ncHdZAayXywgzFqheFmqapNdgjDPVs3Rz
JbdEzy0vbDLo36hWGmUK3mu3IELefKdikraeuZrPvB1SQJeV57ZNaGSCGR+gk+D9
1imrMGfdYIzo1ZHARbavaZF8d80DDvfEmxvbSlIS7iU799kFZITvDnsUqhNL5G9T
PohCOE4Sk/+5Gx/RSS81QWjQKcQTZP8Peus4ef9X8Lld3z4/VviUs4BIQUuVWkd0
4Ftx26qIvR+CR27WWnDSfihNM2gFWduBztHMU29bqvAsJXQC9gTRNPxWHEBWeaSj
TTp1o6h6SMFQTHv4tidPE9e4KiPDJ03Yzkg+IZnUPzLAuH+oTxA7YobwyYHclbst
oyOS/swNhjkilHOth6Qt/p4iXBL4Fe8NUtzLi1oyzAh5lW4BAh5woNsdC2I52Q5R
cLdQGOcAWJEejDbz/6GZ3UJdyG51HxeFxTTlnIU6VxLkvh///wgw1V1E276lEgdz
x5WsnWmnagPJy9QXEAKK5tUm5QocAJHiMVB1JuyWfbvUud521hBYb27rqCo3XtiX
vIWeLwGYBy0TrYMXnGbWLqsQbrknxVY5pQ/TI83CVV7VIlAydAsQ6NXHv2zTgxMg
55M5dr6wSTNpzNKoHfT4lu6LHSyK3U0b9WAN+pCRa5dgKZg5ECgnr9Zo29JsBdPy
8AMlCHKsHrKdPu9PFlq3lYXJ3+POGd57OXsUw+BoZXZOb2WdmJovm+5p/IFL4Xtp
4osGTTgbBYXRItI1WSD7ILChDpozrpTv5Pj39Cv8PAGSdxvr5CF36vW2Eb9XTJ9v
FZ9b/k8NIwTAwocPmG5yBzfXZdGjJtumVK4G66R96hvd0iaOFPojnubEWPpiz9/v
0ClqBg9YBPhTP0GC1Do6ahW9q0sgcGTm2rdGVHMx6broUzJFmNZAgIDIzigM1Qrc
kneJ//bAIi0OiTQ5GqWWWWx2ynnOwEC9M7D3GojznXJIuBo8ZTNlDpytvHQSIVFJ
39pSTljEYDCe3zRhxXySjdcmx7f36hUrZBNaociqq3AnZhidPzGzXFyenWN3i9YF
oVlJ4RPDEMNkMdnwqCTB1kDuGxfOtN50GBEbnLUHm0FoaLcdPn65UfDLd/HDuLKD
cy9xzAN37q6Aos+lbgIt1sOvPRtB4pUKIQk9AUJ0fARU+clTxElEtiWyueoyJS5K
h6Ewm6ZBRvDGMFEyzvl4isrI0m5YPOzqHmpcYYFT+XdnJD7fVOLXnlwtoQI7rOZt
A6iyKVOtHo2P/lj07vfWRodHjXbxITv1rejjj+rNBqSdfhmcIJoppXHnQHvTwGbC
gyDlKD0KePQhtJ2/LEhBfNRn1KRjEewrScL1XQZV/KKKHuLwe4Z01knzL1laKXa2
oYiijlYl2aWf1WDr+DcTYXGE2gr41qmKl/ej6hwVmaz0WXGDrid2mSL/9wokkgrk
hB20/vo1xNHGAEweOTsNy28HhKpzi5WvZJ3w49vQha2plahyV0+Qphndl1xX1eER
B4kA/UoCAdLKkVuXNR+ttkG8iT4JTKm5XJGUSCn2JvbW0bc1v6FCk1ZA35yBa48z
0liqwtrzymLFnKZIyzuZrmmK7xhQukBpZDiDu/3/G6AmZX9kvyVA1N9C7RY5Bj1K
u6MLtEN4Mbn5OsB9pvV7/eGeYPlzzmP2n6dfT1PpNQYaidtFeSFhX/MAOute8Dlb
YbyNU/U+NleVtv3Fr91Ogab350S+AfW3km9LUTYtz+BXjyN2UR+LR08S8FqxlUIv
Xi/+fc/XOfvU9U9Vl5jir3d6qjfrWdKUnHQrIaSJjNl7bNZON2A/mg3mc4MVqbFB
+wQcboHYH0j5Kt8tClRMYklAQ4B+o+GfD0VLlDi+ayEbGfzOZz22qaTpoDXMAkDN
We/x+ryGqYLy50plkJFjPSH71Bc8IV1XY2h+viFiJ+fOCbufU3FOGoIQwWyE8ypQ
iIRx6uGjKcF9T63EqD4bBUotzxbmrdvH0arCzSTzffrWc4MikvFbTaycgW+BHldb
Z9bwOS5ZvV8ShR2OjSQKlrdeQzoxx2GR0Gyep1yzO4MeExY1QYX0i1/+axdGCQbd
IVlC2AoDjdWS1TMY9wK6oSpWQWx6bQ0VRPipObDK2RqJ58a/qvNBbWm8Ln8P5J2B
91vYmvF28+wAj2yxMPM2hYDCx0TqE+j6JoVnPhnu2zB1zABJc+Z1xDVUSoec7T0Q
VwCyH/DFWtnrikXTcXk7M3+LX93F5245ulDZupIFKDbm//qU/UaQAPSOSznBVySX
ZEU2ziZnRMmDepvXyjPcdvY/pbcThNsKAI1VzfUTL1wsJYM41K1YAn73JJBQKhUh
FdxpmpgQK2u0F1tb9oI9PBCj2/6StwkCUPlCxbgKkemYoDSZUpqk5cGkU+vhd/Tp
E8Lm7cZ+C5lsEYcV6hjwkIt5OcIID9ATiHPrHxtvR/6AALGgClNltbX/no5MyvAF
p6wMSr9FMLLIoOFdaSJ9QdJHefkxF6Ve2AoV6La3mxBP3y4h5kb75e/M/DgtuavQ
QEd4tvksLFKwkmnaU6ceFQnVQp6+HvHKwhN69tdkiOXkuNGg/E7jT5AX7DbVDXoG
Ce2Cle9ggNBCF1tS40JaXamMUSgJLmJtK1u4h3hf/MpCc4C26sPrRs9QgBI+8skV
9mF+EzQHfpxh2wdR+fcUIvlYPtpOYNrs3wsgxruoIuaVFCN5576gyDhjkuUiGCJe
CTjWEIDv+s1vdUiDduAG+vOVZ3c7tFxL1cNXDwuP1Ed1v4/tqD4xRnscE9AzQNJi
UcRVn8ml0LmAaFvf3BMXfRb7gtb0uOWyE5WtMM2ixMR3nhibGhseZC6V446+taqM
xa281sPogq4X+U2t5uQAbTiVYxACxesnVb3WxWAeatX0C7O3AYXIA/gEFmJLytUb
3l0R8u+WsiS6+ga8rARzXkt1zQmFONAnt20jH1LgZiXyN4eJlLxOexhFuu2vlkx+
Z8Mk5ncnRFRsV69LpYgRb9FDrqaoormnycNz8hhKMn1WQo/GyZVuApDcfB2V/FR6
0zXNAzItwuPbT7X+4Ts67QrgOLNb1py/odpmT63cuCTszwqjpyTYRoEh7zRT/mJj
EAPWjCAlspL1qm3S2Vt3qkZdugVnLbCZnX7qf9Kn3KpB/oLTqlj+p1QAlqFN0BYi
X5Pqd9XG3nUbrmN+Jk538U4iVvZ7shr3eSXKHPu6KLJxN1sD3Jvcs0MCDT+0MXUA
ZPXfGB7LSc2Ol5pYNpcW1/eFldfFO++7yBAHsAEg2N07w0neaANa2ioCzhUwmpUv
LwL/mEKbV92n4HESv7W9cvnv+nwoQ4KtdeSLXMuWEryLScG0APKcXTDr0gFtdUvg
FnA1Ak+QvGabdYHHmO+4ryuvnj8FOyc0uNmGNMmCxBbAiXKgCOFMZTWcyEuQ4XQR
FbG5hBXx+FW9vQty67Nuj6QfSC00+kAkrYEfW0DolPR3rxJnq3uHViL2tkGYzenk
t1S7Rnh5uLOjVYSlKddsfYV24p8H2VMYxNsaFP/pVTSE2v+5xcI9/fDgYe4mpF7V
M0FmsnQ29qliGNpQQIeA/0KF9tzLkJG3gDXkJ0Oysn8WS8UQi1RIWOge9JfafNu8
z7D6a4fEfEuPQa4sozF/YJiqr92vWOGVSvvo/lzldh5tcEG7OEJlivfqxsciTThO
C8v54Gwj1SUKTfovdAmP4wGLJ9Lo4O4Q5SKsgg/9opW6lHEYZFrOgY3i51QCysyH
S4XJmCrXy7L2H6EXVTSj39NBHNdLkUGZiZ1syeqSLKIx0U95h3+CNY1Zdz/0M3+y
AnmS+jD8tQDYfB7UKyACtX7pRoR2aj7ld4SjNsf1Cag8iYRXEZCpHkaILmnPAowI
CJsdii3tZUw+dx1vBJ8cx07vC0D0+xcBpoh+PSPh1h7oRYvjTpKYhuRV9fugYfCH
Z3V9V8FXAz5PuMuj4p7/HotdE0nOgryWUaOBo9hyp08MSOxakG8kITtXECzeUGox
Yw6jQ/EbjsP/S2ptcMAIOiVlxrdfI6fcO3wSyvSzwCmZInow2GfghkE46jTqt7oq
DcX82LioSMvOgyhzTZWQXNoB3lmKik8g30deyxJWMNLjQQJC0LgjjFAi8bZrXvw5
y2if3lozsZE1Uv9XloSizj2p6RF66wGYxRArq28h/aOl1Kgdt8Xl1DLOxMDqvPfr
Zh2aOA1vVdodRPgF7OFLshjWdQlg7iaFdhYuNGJPaQBx5IDJZq2ww9dt3fZrBT14
hip8qyDBpfIMl42/GBNAe4Zo/yORKhIirMNdCoD16ooFjaBd/f2uhzSyzCkJwtd0
4Y4Uh8g7ccqYXUSci/E/85GX/CcEFcJRstaU+e5tyIHBv8LpiNJtugllXlDgVc4u
vvPzO/3+xHYt7As7AeRrYvNgeHxikhLAizwSF5hUMcs3m5EVgZZyeTiEfbBRzeVW
8gESlDoktm044Zyi3/HuJBzPE8NTyqFzLO+j5+BxGp/Ob7b2gpwykSsZEV9mKpPh
rjLbEhqUfySj7pLAQkToEEcmAOpw1bvVwPdFSyf9tII84sBqUyjryBTxYv/PUhTz
hDMmyk/bGF2C18QqW+RvPQvBunGnvIPfDgODVy1+y2eDSNvKt06RXNQNoWUlwIeH
WbXG44lQJ9B525WOPX98t1qxH9/sNEokjKDYLlXdL2dqOPexwBX6mz6PZlzoyJPi
W6ek5DpimwGZAsJyFnoQJZgm7ZD01CIg7HAL3CQApiU2nR/SuWpBeLu7vAZjXLg4
vw5lMGSV14MjpwATlFCSZPTWIUwjSyaeumLgdSCB0W77NDUB3k6Sf/T0j7kkaa84
K33onAm30UWstJEs2dtTTX9CZq53TZrZtiNPElejTwPTyX5nGrhMgZTFVD/T5TCF
Sh02KlzjVsSaYrZNW3/tmj6OlLa5CVFVNyElkYr6M14id6rVZySnXjLlCX/zniIo
2YL5EEkAMfB/7bHa4ZNjvSDTM9bIXAHKZjYGoPnvs5yqCJgA/ScYsedarBWZEhbF
9GdxiGzIWr7NZOkN/lM0RKFgL+IqwVbwY59D4WDe1LDvI4Yuy8MF9h8x2/kpFt6l
2w0+vFlSu74n1xZvdaKihGhQWR6Adz1oxhYWzgTNi+pylT8+ysif/7KOKBB+b+u0
pFXWSBmwhfbcfLR+399s686Km2vj8kutOqidgNtJI297WStjiK8TMVoGVfcVVnX6
UPPW5CPP+gASZwGVQ7hlOUEPbg9fDleOHiyR1MKZURU+E/LJ7EfPo4CUEc0esXuT
1Q6aB7zYZNsiW4YJOF4BB7aIyhPcEifeAiQDfE25huWkIYaAX0bF1H5fu9OHIUn7
8Q2kJ+ffT2x1DacPpa12AA807YW8I6d6lwWANS9py6vLuBEXHXhS1fLRdmQWgis/
aQktdzzofWWA/BveSHmOLCl+pRQiRmMQud+5xEceAX4NjZvvhfNknGeekaNojiuX
R9FQjujsL0SW05Y23RKei4zE3t12MawJ9GM0cRKBCg3FMNLUjS95a2X/Z04HT7tw
pebaLgr+8Mb/JEn5NwqPK/w0pXMEHePt5/3sfI37kS2/1Kh1tbQqhn1KgMkh360u
EQny+P7Pv30LcyBcyXd01KWWuO8uGLO2kID/YyQzWF0ZJD0TRo6J6FaRO6WOMDuh
jqmfjnBEJ9JfoeE2uJJFO4591wYrz7A758Dlk+xrj5epFUUv+yAlFNBL+wJWeuf5
lmH3swR1yf9K2JSvW1IJcD2y36Co8xuxRpXIH0Pu1EnLDRtMhc5y/CjDuqKg33Eg
sofBQd+Jh2CFBuKMNWtL2DlQn1AIgSPVEpZ6PNj+/hPszNXulyxTYeAb37cdBWrl
aY5GWgFYp2myIgxeAtwf3Grs6vx6Bd/b+YRiiq/PKNyCWGaNWPvr7HyW3gzEw4Zw
aLpTXsRS3DsHazEhI84zfojwUp99qgLtviYb1BGDpYGKzXYaxWinuMsp+4M+P3pn
4Ro4EQt+HZTtb2Gy/mwxcMOGvYCJMcYdC//gFg5ZdmOy/2F9+cTxQJ80+Oj45+RW
4pVSKNGnrMkbpd4yLkwkRd2Ij6thw1bTpBEwFp/KSilTJWQG48GxZRZk3y4I6IcN
6zpmvqe/0+/6rrIKenoZvvzaEGMiCR0AwjHt3sYX4NywJ1H1uwH1Y7EnU4WevmeC
nYdsNsMiDiMtGwCn6UxGVd2Znktl08OGvbTJqMOfN24ntGvCi/PQZCma040sEIc6
7cbmq4/km7pJNGjPzZhj45X76wNVLwqfLpsgW6PeMHDwluWcpHJMGus5qG4X994d
CyBt0E4wqGnAcnrLVz7jSuT5tYx9NRqAcyWgrotjjYvcZq4ocquAE0EmcfvoddRt
UW82B/HCh54UKGDagA1jR9dO3GnjwrQ9O+41TjeEHEaY+CFm0+Q1UnphGzcb6cmB
Rvzw/Nf9zGHVEncQEyWpoZxwJ/U/w9wtpSUqcoLMx+PRVvv4ni68E1cSmmqJXSHn
jLeglNNjn12QvGo4l23smEI9K6Lh+O+vwyQ/RBhHJ0xL2+Amrj8sIWoLpg8tCoSY
7hMWNdTmJ0SFDTF1nMg4iZQ+rw7B5sn6xVbVu18xvYimPJR60pAuQIrgjk5ICXM3
c1emWEBrLFE9XthQocP4/oE9x+D5NCq/Khp1fY+MVI0WEjfgheFjjpXttNVHWgoI
mR9WbaF03Xh831qVeteYYW6FdbHnyrjeACCU3eRInGXql012tT6zcvTBe6WrisuD
gFPa6G6YWdaTG9PJ8jhpw7MfvImHhKYV3wwWqlJUL1vpMTPAe7JOOdT9f/98f/Uz
1MiJHFdlhPap69ZJH+NNwqob3Vx9Z52O3f1PmHoIHFvzMq4ExYiBNmSdSMMwVl1f
CezbxZ+L3m3z/VmCJuO6jc70O6l/NVC73rfPBUST2zreBpeoaDckwAyrWgi4zeJu
nJHku1MXelHeh0lzlfYJoq6N2VMaAUVySfIwVA5QdVURf8fIM7p1ux5/FzwIZtN9
L0JXDT+OBuQOxzNl2ER42UrV5ZZxHIO2WkErAMLP73X5ktnYTmn1Onxkq19sKgsz
ornyYLiHkzVpt3xQHdJaovahKBlbrJOmjZRu34bnpgPxQfDgdI4kXCY7afTbBnVx
EjGf3pgTp8uCCGPklxGs9omz5M+6xyKzBgwrIcT1RaIKW+fyoU27ISLTqrNXuQ5t
Cr7ayN3zkV2Ng3oPOb528+7Jb1oQ8te9epEcwtgqjmJbkpZO276TkxjOBoYrRXgU
XTQTZgbEN6ru7HZ2/VmuX2OGe6QFsq6lVeOqXVLRv8ps7BAzRfCEcYSuC8gLuAwG
Lh4UZnhmGY0xMmtvLEaF5RgsgDG4fXDFAX1f7sl28LZPXuxrMXDCZfBrGtiFnkUQ
1m/RjDvyB9QKvc85m2Y96uOeZxfJFNhsLtCWBdALzzPKpEkCTodujf0jcGbj3UAm
hjdZxyYBZs+kpzTB9kI3PMmalMBIynhrGml6CxTWZweKUsGuleiIVSdg6k83MxYx
3IwK5y9jfdY3qGLAL46+8OmRGNUGBOqUL+vTF4kKsQ5wud9KjSlYWysog7hE+2nr
GsXhtn4zsOI084Mk11LufJP08XGiyBwqpD2hupwr90StVWUk+lnFm7MMZ1p1zY+l
HcYMDHPfba6bag7j0tb7uZRISGgPl3tYrIpy0QiV0walph0rc40nC/Rw0sbg8DNY
SesMESdTWssZGjI3YO5xCwQqzgWf6pnRo/E6XmDhh9pvemC/pHxtnOnELBDPXt0e
HjA5Fhf+71/ZrZskerUsTVvjFoaFWJbJuJIWlW2be7LVd86mORGxat8SLVi/R79l
t6FR3X3aBM5+Otd7DYvekrbd5HlsOVI+BFqi42bs5Y0BVrVd3lB40SbCwDKfTFoU
rBS2Pegyw5rZPJkXvNpFwX0z3L7wm3ZTvQKyEJk8mBmudp7gyUSCQdknqgBi2m7+
UahpqbcnAf6TaCvOpOhckawssaB0Zsh35RSjS/yJXQYs9wxBpCyNv6YL8eA5FZQt
iGDvQ08wpzBw5zmRk4NY9bcOkYIvoT3UjMMBbFXiu7ghjw7VbQCtYliwCUi/1PZN
TJeWgBPMvzZLmRx2h5+BUsV1IXfx3e4lwUonCG4TWFMSIAlxVsssxa3unq1kTyol
eYvIp5ZXf9d+taY8VltoANx5ZO3DxwrodNmoD0a8O54/HebcubdX6qanSNJBE+CA
mnk79jWsnoKU9TCXLJ8uz+3EfH9nEH8CXAXaX9CCm6ZZnEvmww+37C7KDW7ke4xf
o6/AZJvkXwG3nrqb6Wp+Dit6t/8iyF5o8X6VWimKpgwsQ3g3EJ91MwO3s69YfcRz
uUw7d1unoJ3AnNc+ZcpB7DYaYBckwjhEFIz9QtyUKPPm7Si+iRaNHS1ta6Kw0tVH
8RgYqTeeTfmI4g91jurUAaRGAroDMar69ebmDZvYUU149KSr+2cVDcMSYfOUVkPy
pJCh1jxJ1mpviQAOQj60pnSGikWYfxSEAmQyX0eFEPB98Lnoy8B0dr64dURaz5bH
FJ21tTlv/OipHV4pYJtLQAZ87J5Mym+ZdVCXMZkMxZivvH/CENH1TN3qIxiiTgIP
PxQoi/PKRg0TC0g/tMBohYFa+aH6SZ7cagOugXaJhkQnasLlXjyM8z/CUKICkXut
8KCiQwS0EUV6oGJWPuEL24aZJZJV/IaeLr+0CVO9BfJpzaiJPb99jbNPb+DSJQgE
mKFjHA8nyZ7aAKLc/IXACJgzSzZnbRpjVsRAzBnaWeOJNYg+L4H6GcR4qUnhUKbx
kpjxgSCe/QmeV9XbN0hQK1XQbP6SaDwFwsMQK8cSZ+377q5hhu7/zN/LyIfEReiJ
oiGa9Vqyq8JGvTt99tXsoIrHjDYKW36EK29139YeYJeBaNZRqJXOp3QuHSM2srjR
2sr7auvmtdfChHibQQYi4yYQLEMnpgiVrviUj6LPpqjjGAo0B00tM1UzbHZFCMjk
gbL81FTh6th+GnrBiV2SUkDImeEUigCxHz7ZtqAu1iiAzx22r8pwBni8eOkiiMDj
988jgLyZGhHnU+uu5ItWgFf4l/Ti28j6my/8xIcaMu1J4IyeLbS4c4U+BWmnXrcl
VF4QH9sSHOD5GH1m+3Zrd7HEDBhi5GBtOaMYPe/4jEUQ6zLjUz5y9MHQskBSBXoO
+qgA5XHBj5I9y3d4qX6QXE6H01GsGPGeC0EQn5SuZ9IBDUwCYJ9KA84Mt+/iCJIg
gMOGykLUZDX9QhgVkXIW8sYfs/OBZrjDM1j6JuxccO3c0si8XKNlk4P/luvsDwSM
vDtLU1+6ilQFb2MK4/BFfOwqKk/7yZkc1nUM1+5Oep8cgojwpI4Fg+b65l5L18uW
zK03KC1ZQDImt/3rBzwH7NUgCOvORPea6+LX0KGJaXjnySogx+rKEsBdmO+ds39/
6TSpdHuo+QkCszjGqNUB3Zc9Uz4hEVMnwGqWR+QwmPMUguzBROlxeQbCO2F2CNCT
7b4gq0me5ntbI+xEneGxX+FlQPvGzjsYR8Lj772Dnor1DEoKqReKR5ieZGU6NGMz
6Lry22wKvw+Gzm43RXKJzV9BJIrB2G7SAtw1n6d+/9d3JAVShaUoXTsdGm2Vh/n5
9t1SCSoNRgKLqibEVQJ8Mzwer1rwgbA8iviWCxXKVb3+1H7IXO5hzM6+5epH6QLK
Zz9V55eVtmmIeoiW6T/QFosScjiSR6+1suosy5nG1e7uAznR6oTEM3I5OAsavhLv
QetmSoc22+X6OTfcmDtYEhMFOWpNn5X4dkxIfMMnSnq7PfzT9UK6RgKWAw6Nb9Vi
8nQDtKoqHOgzynsk5TDVKprlOGsK9lABjaAF73xv4CkPOtbtgTMPjPH/fkm97ypS
eltF/84wihimL014IuiJr0FAadv1I+QAyjLAu54Nnfc6HBERXl5XG1jiloIbw6ZQ
kaVzpEBeCtt9g8yuoKHAC5Bf6Qp2wmPuhDE5jBONPhdM582l6H4fjnqUfhgYR2k4
OjlEqvXEh4O9zDm2jJF68pKJLznqhkyxyLT+fkIzF2tMlMDwz00OhrhEf+74G3no
qZaI1DQoKj6S0hbDzAaD9KRnyBh7jYYNbtuAIFZrNzYkpQcwBBYn+ro00FdbUwSr
M1jY0cnKV1sdDVqe/Ip7OKUQxKOrKHQ8BYOBTcVOH2OSx1z99yXYz96ablhOQaRQ
owQ9FvSTxcHsKJ9LrP52/zv2r2lW0Ytx87yTnSqM/uXC++Dj8TNnWYZ3UkOyHXlv
n1pwac253ZzI3oavIB96K7aD4GHcbGePDHNVXXevcFFXkhtxoafKcAcn/gE6+deq
dvdKBgOnvqvBxSEsIvNdTdR17EmbuDEJA+PH40gDDuukx2BxjxqnNvTDzi/1CE+y
JYH1aArzDwn1deZza8X/K4FKqguPHcE9yrRPELlKPu1MJI/ROgtYQBdEMGirGXSL
jML1YF+QQWEy8APWXXLAaKHJl8JgQk7tv+lAIDYFs7Htuh2W5/jecREdQ015owlq
AmMAVGDHu5X378lwiqu4LhWFeO2g9NLjiNthfuOamL9TfmyruKXOUbu+b2eaF7DF
qaWBj43BRr+B16x9avfTJtmX3pfuKSUVXMiSQa8UCk5PjRHagF/vhaJDzLwUDYAT
KaGfNtSHXL2gp5/0n7/8JB61juKo8LvI0/4qp4lp6h9DVIfYfe1jHcxe2CwWOwIx
esCQMxAEc9C9NvTT5Rrgh4HCSvkCnScTM8y8Cw5Ni7kuDrZ+Os5GrqE/eEO9OKqy
8Mr0207uNwseQJoVHUvAsr/J144sTqEjNrdnJFt9H6VPmDaaDprJ46Pc/5YcNc0p
RgYHQkIxCQ26+CbfcEZo0SvdsiJcCs8BJ5fC06h/BnIgDOZBy1shyH/0Uj8rJ3BD
qdvF6dIty31BXEIJr04PTciOcZI8DthbpQpaveKMw708/bkzWqCPSc/dInYugYyk
b6HNTOHV2IQAjM0fKiOab4qqkaw1JQNBx7rOASjyCEVwXs4iVTFDDBa7DNPE6/PF
8+zK3V6wnSrQFU8N89Qv+nsAcNAO7qycsDegGuWTD3W7cRah/0BVHKzcS1bOqHLq
5Ox2fcPx2NeFD1FLDyTEsRbSzZ4DtDMgNljvxqxELRbQtBdFcTJ1Ce3x0dRnLtDm
jrA1aDIbRb5SUilIkCuf0ISu5KwNhsckHjOqYq5eJXBTWVLuZGo5+9WBKUCCwTqP
YFv46nqDFuL7qc12FWasl5ef98qaZl/KwrtL1TUAthti4siN4RuiFhwdB8tk5+tP
YSbPq+JjtUVXSo2tnYZMlV2Jdvf6XRSqgAQe8EMP+/ZH8QukulFzVJYhelEDdbSB
8CsUg/MwxiBfmXH3NaejiepRLEeeu2HbuR8+p2cLXlPCqIA1FGk+iAHY4bFftsrU
LGR/jKYYK0PgnLBnLprjMnisX/oSwGkB7HnbMdZuclr8xPvBB1F5MoCcl+lUugnD
0NEBBHCdyaeVApr7wbGBPszxLTLUpnTHxhZV7Zw9iZ6eTXGLpmKxc9VQg3nKW1qP
kC2dPFU6BQ0yB5uBVHtQeeLYj88X9psl1VhI1CRAm3OITP7EEaKVW03fxQI59RQU
kDyvhmvmGHYBYgyKFUR/u2zlF5RQssu3TiTzQ1Ck2qrUOOtVoIPbR4BrNwPpkT0Z
wOx0Pjd8A+ZUh+9knaTSbDsJo+8GvRgYbD65VS/063DUAUOwufXE9tI1kOHNXQBU
yqkY3gNRlmnR/71NKptdQOVtXHK2Qyf/yFEQLLO3P8Rft//vBDo07qEGwSjlXCz5
6KeMmAvmVD2vC6KtZOcEK9pgGP3oJNc1iZsur+WOk9dhcNnHRglEzzOT+zOm/f+/
lh8DqV6aAPS99WiXJd1XoP/nZ4k/cq7zf02qG04DkXqUufegqweiOt/DH9qMs5UP
0VpoNe+r4B2himLX/W3i+ZnZBI6vMRVUTc2tNjHTHlLFC9kpUq1ZZr6g07OshYw/
Kdfv4glAdj231AjMM18TtppPJQZlGxMrbtVpS4jCs16+qPBgRbrjXlOGDhxU+Qjj
3CmvVNVgvIxwFTwnFofB6fbesn17D/mVlrXvkv7ZEtnhY33pEhJNA5E15WiLC0fH
nBHDg5U0rIhb55Xp9KPItQAsDTpP1OYAbQRR3BBDvef0PD28ntYNIBgYvtyPQPE1
tN99qgVcl+SHcn4g9A3s/pxlHH0XgE/TudWW221rdc+GkMSy90aatrh4JeCEL0Nc
DtyAG86DtqoZATPdG1oHolEblxwrCXLCSFo8Tn82tkIX9918DLY8nz9tKky1lrKg
oRmeNIKC/EJVvDxRMiiqy+fJXXP2RudTvCCt+I2aqKZKJwxKvw3jgdGHlryzNPGW
xg1OnBeAxKKDeKV9jhYMs7m/nUWzgWTQw3z655KeR5do/etTgeVxXS4te95bTwcj
WMo7iVaetKori6ZN90q/jz+PYGMZsRKDBks1Q1KUcw1fLurx00AH2itb24LpzhXN
Mlm6Fxwh2piwgtimDzYSPhvXby6xn5lVfntjVPgbFMdvsX70Vy8OZSUpghSu/TCg
KYFLj497iSOqo/aKHUsV7PAMXZLTIUiKR0o9HYdfY41ibxGHInSZjmI1YvJk6GKX
qaDgdkrgn4+0BDMVCubV/NB0ssnXbO2fdyFxIMLHZvC9Qzza23xgRRqdNkz4PI7B
CBppmFMf1oLFFteCUErwGc6AJYUCcV+duSOLflRfpaBF3CbSaPqqDcgpNNCfXUXt
AR7tSaN9+LHRreK07MQgn2j8Ks+WyR7uVtUAVXmS7+jZpGCmLMaJ9pNqcLf74qfm
HkGpjMWBQODK0whqYYnG0iVAytDj+iD0JmBrEmGIHC+Ds4qltLsIv+ukK7nqbjTK
gjbHHriVirVk+6RsQNLKOljJUcsW1XMTC4iKGXOAlcd7+vyM+nAQybivOMp9svOZ
ipYdAebv2HTSx24AtKPoGXey81TQoo0jWzf0BAvJff+UOPdu4lk4bcabcxaksgjx
WvsLZ7Dyt1Zh5JLRPuwcfPGKSt8gQHGJbYZXk/Dp5hhEu0LZ9O3I3TjqDdMxZdgu
ACKXCfx9tRJ1ZovRiGP/CLaE6XAnjRx4LhEfoJMBW5FWkhqv8vneQHR+dCiDSaSd
Hyjld3aYM2LKOAJFVSjkYehQ2LPynqgNYjdQ2CGO+/w23KfJxoA+uqWtfNjhSlAQ
4Sh11x/yMQ7ogzv2qJfPTM0mk0D4/NJTElxTv11hNO+jzsGkxzby/Magy40cp+uk
IA+xVBfHDTZERBvweAG6gwNfzT08ajhrtUM2g/zpvTcbko4wCFRTD98+eVopgQJN
W61g/1TFWtmwRduFYwIYVj4oM55BrOBIvVjRI+AGoFxMro7w5KZJVktKG7/uW9MM
myIdftw/cUw5R1eGNonbL6RiJQzcuOjswDkTc8p17uQQNSxywYpVXbZpFrpta/id
1MFiAwjxCrgCkiaP8Ef+KliUiabQIEHYelscbRc0VeLSpOSpfqDlUAbhQNWIwF+1
zJb13ltGfPAQR3yRR2QjQXqjykkPVsh9RzIy2MNGjjTHjpQzCLu7u7Dze9laHHbN
d3fA4WXVEpQsBwNfrAVDyEGL1xUc1dtT6b4WUs0tID41XZT4CRkvhFvxYvRjgjhs
GIrewUUZKZaSPDlPPW1uze0T3rFoNOrXSem0uqL88HWobfXqvfhdVyFA5s4RUMqZ
QrP6igJTn6ZZOGO/+MGQzKW0eDAeH4YtXPUcqw10/X7hqGXVyq60YF7zWb/gY/so
nHAezWoUBlx22m/5nLq7bOAsSIww+9pVf2rJua/lkjlKQKXPARApQ1p59CvqNUhR
1KrDIqFlzVBACflXauYpXQCcAl0s1XKow8ThGV+gKID31cLRu/vKgAeoeklZAsuI
rp4DSbbHnLDsSf96nuuenIjE48wKAgniZnXUpA/kY3MwQzWw/hCinjJDs1PBFNrE
KIy3DLTNw1W28BdB/1RDplg27H+CkOk8nMC8a6nFhduWcHpB7vhyhDYTcssOwaZZ
ecwdxFVYmpHIscEJEjiz0Dvg9U14nQnq8pyoQgLkirFu4EpJLKiCWzUpiwKd/K+R
mNghg9buAX6WKbNF5dx2ppE8VNOaPwAe1p5Xw4jGWiPvxFfXgNlQVJ6Ilv5a2ty2
LAIj6jt8RwrlxjiJtvPCQTbmEWCcCkVazGFlcjeJz200/n1loPZ2M4a9iOcSOgXz
dWOPAUszlSq0QEY0yVJ4bmU9VBWyZzM1xm2S7qUxHiqMskqRDVRTHte7Rh6nWTuk
NU9t6jZHjvB4I0+1VUMVKOKC0a4Fh8bqK2dY9ZdG8v6rRXDUMD8k3IWtwJ/tMOAm
atNwmynmRt9A9EDjej/PeIFShuBsPLuu0R5B8GUJLpx8JIT0Wz6FynnZOCkITTpk
O8Pa4ktPqv00GuAMQu+R/5Uf4veD0etfwvIedqW+HKJRznGvAOhgfo57hhihFXNI
40kFSicsiHg595wVJld1yuTgN/tXN8fUxUyEbz1FluYPel2E31OZBBtn3FpTWf/t
gy7RTExWS90DtV6ydZIDxgi8kaJBuJo8EQiwIcI4RZULP/729nOKXGAiiAMq92t6
dHVgLoLmbY/RRvgRbDSwtz5yWyqg1IY3S9nCM/CrscKQ3vtRBiiXenTYh8XB+ivY
mFqhMXcJq+TklqAeJvjjnkLoF2f9LxgRvWwAPUZflTpfsE1zCp6I5eZXqZqr4+Cl
z2UXQarfNPuQ/qLuc9KZYIkTcbAEvRpKSNTYvk+wnBwGUJiLFbWBCOWdYuBe1Gip
B+p2cv6+C8ZIevYanIWDrZpC1nqxhyk6cpbiPcFl1BtI7Hk/GANKoYjp4d/c24Ss
s0FqTztEAtmBc5sRKLaN9wd/w7xqCmPo0DOtOgScpLC/uGR25Ug23jXghkwMTZ2X
kfDOZ7NBWRhRgQ+yR7MAridm5fpL99SNNtvXeP/g79Ltl5FQG3OjR9VFnLFpznRJ
+9DgMSARuBPtg2pAhiHntWPdTmZ5W0uZ82yidATSVloim9kaHdta/PLJwvZbWEkD
NJb2TcE5EhDS3D+wg8ij6bOyb6ps8fIv/0VfyTkY3n3kRG80b/CO/XNRN4iyFwrO
IQQfe/F585NxcqJBn5iU0pIQVzbxIFlaNnoMQNCREVnehTy7ARUdU8/R0iL481cv
bG928DnfA9CdhJq5Odg2RQkRSn4E3+GRp7N9A8dh0zArx4kq5eQBmriHMwRgeCh+
if5y/Nm+DAOvkglJWMgd6BvFDa7ilyqdSdC4mi5Ljivhu8gqtdJnyzzssBWLXvLT
G4NhpFuacaHEI5TnkC6rvwgEDKhNDjflYIPGhoKhwv1F6dFrZEofrz0FocQMU2TL
5N/8k00UM8XAgCyMLr4sqy0Cs92s/3g/GIRgnYVrDbUXvfX6ukx+B/5LG6vGbofX
Pet42O2fwD8c05KP5dKqgHh7gbSurRCSJje5hGEnOSTsw52DMBfJvk2Y2JO1WQAM
0Y8bVBMDkRDt8pH7zolDWbSknmw/ruDfWNFWaN1EPN98Ke7QldU2R0qnY/WBhMXb
SfewSMW5hgWgSx7nfGofwD4kXsR4cv/7+T6EZlYQ17LbLE5VFGUzwzNn0/iPuVMY
aILrU3QaNJF2x+CnXk3zXa5Mg/3ifQJIkgllND9t57RvMEtNn5lzZKwSl82nwbNL
dJri+dYIBaeHEhdZYHEZgt1E7EyJIYolXF/Ge4ADYIeXXBAJft04A85O5td8p6+m
jBfq5ca62jIuckaxXkkMZHgcevAmIbK3GJJtUkZoUDFUpacSx9ZnYPH/qHEuUThe
haPyXGpbweK6lPCQkEhjYL7kziN3SJmd8NsDqyUIrzUXGc5dFjoJ89lTfNzstWN2
LYsL4HvNIjqFTA2s0qNcNcl8VGeECYruEy3IVoAIY4uXmBlG42vEJQjh9IJ5vYBh
785m/AvB52vG4tdUY5prJxsW44muSRyene9qQ/WhhXQHKzflOqpkQxgug5OozIes
kQwhljEEDnFmViPDgyO0/Ov28n056e0tJCHXzp/6efqTz7GwngVenReQKTk9j5mL
8/4YhDmIn8rdLtfa28exYUP2Iogwr3/QZUOY+PJc/CaDotRpFznllqLnGzfxwIYq
OIvbvVx0LbIZeu0cXXArWWjvg1CdcP6Fv3EPTX8biEubeuzBgHgFn+RsZcYOxLW7
rhv4eBpbONl8c+ruO6/jmM+fQ+pWI1pOyLtOxfZWtBS5c8UC5dlIxMzAfVxv7HbJ
6OQCOZUjW77h0CYGlJRHJxFECMGJa5/HUHwpWq5TXHgl0lvEfYBqnL3cBsxEU4TA
w6+REb5xx+k1fa7/CjQhduquBY35Hu9FDaUOzygw3MyGlaCkAj4OpIV35OlNXynT
671wWK0Oz00zKNOAf0hU3P56gScU1Z/YPNIt7+WLBU5lrfjQhWzhdDcMt/Pb4U4C
BA/thnceup4e4Y8v5WmYi5kjmfBW8YaMmWCVpD2PSKTA3bzbdpQO7FxO59EUkfH4
6oBZ2wKXerVfP5Xxuk84TTpEUPhVeE+BS9oFHVViIGtBawAL0Q0XE74Fzs53TSTe
aCnIEMcjSN4E7OnhiBRze81bHy5IOoWMRiCLkXjAyCf70bS8in1QNM9ivS6fXjlJ
UzUK9NoaSX39fuAvlrjPpP118w/9u6qZ8JypeoYN2+iYwVWtSTtLWaEnNSA2adv3
CmuUMrtlVh5U9C+bPkmHUHGX1msfoAOUfDc3xHkq3NNVKVML/0kL12q+iX/jdZg5
7jecXl0AfzI61T0Wwpc8cjAX9a9dKQXwcfgyLJqT6hHyX/8jauVJRP2vOdpoZCA/
+WOhnvJyiUBOCIeAe6MVkbsnzzVbEgE8JZbUhYSFG+Sg6kpSiF1T404c+wb/fREy
Up/OZbEg4AYGXUsG11eu1F1XtFYPIGjdzLPBoSTQItxudecobiQ76AW7I5U6uCoc
iCp41Gymfxt/S0JHMhGJkipE8ENls1gtY32Hyrq+yr1wsuO5x/O6qcT7EzRRQuxG
nd6tUtV+tcH7IYmXKd+h0Gk2UHkHL2vIPdokORRzPgvE9V+SkMiV65SCDYYIRVel
wLeWAoT9iAix4F9b8BKjjoKN0S+oaEAJB6Q8qqEVboOqcIvLJFi4YAVHxWpAE2wg
VdAHZNUrxD44BGjlLwzHO4Q/1ykuR8YX4y2VzpTpmz2yJ34GuWNr/HMnRfHHGjwf
zfqaqdafxOgeJDGYMrpZra6OrZBV+n21qUx/8uYtxa305QaEIW9TUrn6uRISM36N
5r/lpgxiGuvPIf6n0PoMB2go0+Winv2ML0dYZvEAp6bPHaop7Vrt2jy9TI35IDJz
+aTn6+RrljLgg4MklBkoBuN49ERIrbciFuVi90NlOgftn3SVJFWlq0vCG4cyrpIs
0xlnkhUiHZNpqAthei4jlNzFpH06et/iX6sWhiluHR+NHS9MgZleYpILSVG3dHV5
uLJbG6zJcP+5M1ffFpUeeTgwPcoiS/vK4x0mIbcPZGzJr+wtz6oy35Ytf/JP4GEJ
dRfM9ZWrixViW9TN6fDG/zCHAptlEU4bIQc9xQb595l94lcbjR1KHFtP7xe8+h8t
EgJfsNfY48Lygup9lXQlEUUE6HSrmUC7YISHHoM1b/ReNyG6mCqKZZz+74Mcjjk1
q64zb/1mJTUneQnfStqGM+ytwHObSA/K8mK8GxPvpjj/e8NpghSq168ztECID91H
l/6HWyyAj+1FnRMJ+OY0hGpjxST54GE4lKQc1qASbcutKLGY4b7NiD0L9pFcbinb
ABp1Lbp7r3FkXm6nOfDtkKVPzSodBn24X0cZjlAGW5C+AHxV0pzsR+5eR8Eo4zD4
Ytr//0vmnaR4ODKv5AFjGcoq+67zeqkWOxgn0xZ40BGEGDAnv58E6X+d3yDr6P3M
ZNWTjiu7N7pJqvj5fvrBAS6ponlwntI7CpTpAFfAQTly9Srw0lFBApP8rRGr6FBP
HoXCqqueFRjzPBxo3N/bn9v0BbTTPiBUKJPq6U46vG+ZLEG0h6UVplv9FADOpg/6
U4AI0RppUx97OywFy0a+iROQOrxx12idxPrK/Lm2c0xPXfaVf0q3wHlkh0dEaaMa
0lGdReIjiHUdAFZgLNJKH6BHzDGnsCKeYGsufSvPkjO4L8gApR0mWU+u+Ax72F9g
JTcN/y8aH6anBBuTRJgwl2ba4dWCMn0kP5zQeiM5Sh8biAO1PALIpWI8A2BsBc60
7HdCefA/s5LjHXlISArRvaEItB+ZFcrByugpCDr+B83vojEQjaEr7WzbijGUIuPS
KaYt8170jIaZ8LMr47uz6ZJVwDGowknffMA+tkkzQkc6hqjPQBtBWdHXqDOcazmB
TyZrw6FuD8OOlD79+Iu37Ez3NmAUiWBAO1gIlgnG1Ks9JutCxpyt0Vz1bPQ1ctte
ArYpHiqXsb7MNVpw32H0+M6LK/NiBihUD+oARkB1n4tkEu3CXLttHtpX6TwoqMpQ
aUWnhQy2Iq44GJ93jWygaOi1mDMljJ+eB9lOvj/MBwNYwxe+2Mi2Gx3kCKMa8jjO
g04LTs5tRBkgiYJhBDaN7qOA5OpKcwXGUkITwyTZfU7Zji/+vTu3DgjIJDCkApvk
vLY5AlcsUdiIhi0Wg+yGYbHgQ7dmwH6unJIuyAQ6SvJxvIjd+qxrwf5E355xkcft
jjtKRAHHq85OqNaF0jAd+vbQ1GpEQ+3iijFcImOsLgQCiX3DpyCz5C8/gZSkUdVD
PCBUviA7CwgxkLGBhT4OUtHxsdHxoPMMMh9UheqAhjK2RFaDTxqpxERmAGxYz63z
mddCSRVs2cw2ZLcbfIYL1/uu6mYkJDQspGlSpilR2ww8uD6ahvKtexsB6B9fXezB
0R+NHI59n2hSvErnwDauGVzczB2MF0+bTYmfhvf2dZDQ+Mp+0rCklKucne6NmwLI
9oS55R0mYtaLoXaa/AOuZPGQP9iiu65ZvzjR/8InjybGUGLBxyvt5R/9ggU9EhIp
tRiNzA/gsR1KxmUnLps/ztP//cCGv9pFZVuxEowCKfE8sW0yFME5kUfB6bOFtHp9
MyXu2iYNgDmZynfz5zmuR9hNcyLmMxnBEu5uLmH/xxCjsh0/6XhJL7O9NdQ3+jt2
a2nGRcKC9J/3il09WCROTRCKVMoCoIG/m0t/khXlLP4+MpkvHRBavCxrLjoPP0VT
wSbBM/2bh4b0FN5O24bpTptQid0pDXxtPXVqch0Zc1St+8c1o4sG5CvZGFJTFtgX
RRNKEbIWbHq/kZhiupyfRCs9u/Yw5pYnlVhjmEahVVvHNHLKgezWPRgB87G3AOBV
zKXYfVuZO0UNVv4jw/VYeF2a7qDUHFBEX6PsbJAfUKHFn+zf88un716S/HzDrVix
qSEZJTmGXUjcUW0rx+hlatY463dGi2QkRSinvzef0jc5vS8FWDXumLBRsK7zmpxG
ZTJN0p2kwMys+x/1tA1Qql6p/1TU3iCr34S3TycCTdjHQ/bUw9Djn2TRZEP9xyzW
+b52Nq0Iezr0t8zhrNj5U+5q8SXAfhWy7uZ9rpGYJN2s9iGfGCn/9iAz+psCt2cr
mZhUA/EEgx/m/2QPG5tKD/2RX2E88oxxnfY00xPApgfnaIIeVC/pOU9YNL0eDJb0
nMJP42hkE0GrOjH2uCX3oM+POZ6/NJaCPyt/swnfkd4Cm9HxG+TA3Rtyvq410GGA
2028OqfLjdryNsRg1MQ1posyeFN2a5pmzIJfkTWjK6t+DzzUIQB6t4nVhk52NuAL
BQ8iSwtvfVrJFGxGkE5WBNUegS0Mqeb+yfudLyJUvEIWSI/L+jlzw6Hoj5aJwEzE
RKY9EPGq9p+YkcJD7ODyzuf+E6P0CCkZAk7sqnTZiiRvneLVe5FoWxHaNBZ6vznM
s5b2zM/BS5gbFsM7KYwMqK6aDypGeCUuZSR64bSXuLVwQblHEgZech2xbynBcMyR
bZdIYv+eLZEeaJwCK76JBUONciamVTHABRu4d+heMDM8EA2d1Q9WRwZC7sfvz/JF
Rz6ZvQNKqlLlPaTxbhti5xBZmO84PEYK/zxASrO5KBb85XKBJM+Zi3yJc9WE/7L1
8UzsI/Q8Mvge5BoWHX6cEKTZ59mJhOS9F/emnwlARTbdFwaV4nrM1ObfImKWxMRl
M4hiS1UZSfjmpKspbIskKGcMpaGgazoNIC2O4n3uH5UtAzzxqMDJhMwh+uMohaVj
to4qu+eG710Z3ODDYuG4Y4ybFCkW4V6CYXXVPOrhn4mIWTJwtrI1IqCoQ7nFNq/V
rnrGPTNn+BAAPfIhkn1qiJms/dE35farrSzURtDVGAPJQG5o/JE8F3foLNDBOEyU
JNanwpBx/oQku+jX+s06yDrr/O7t09RwDHE4FTcnaKKoy/QLaAkN12AVQ+0Ua0Zj
tHzeG5zUS3FrG1teeF0MlCg96r1jGXeLU4zvSjBtnu+mwLvYWQUoiCUiftCziiNo
3FVPh+l8wLcmxfpZATUsiobBiVOrctbIxMJJleIF8JiUtE21Xaby/ms7FHsdC2s2
vCGyBBMLPgfWaLg1boF55ubM3PMVk5hSyTTazAx/qhYtGhctE57wY6CP3hZvwu3y
J2DCnkn9/Gyk/zhK+Z26+vf+s4teVKul0dLBwDBrwR6q/0DGXm+63qLndJtsmZwz
sErEFpUX54rTx4EFJYq2Yit+juVl+3Tz3vo2w0ZrZb5fDbzePCOBynss1E3BYoQo
tEClN3frhVe3NBn/iiLGAr9MSwqG9RrJlmR5BvVGzEkRRyOgDWr9ozt1VcdN+EhQ
4FwUXzx4T47qA3k1gy2mwdochlzYUDqrLVbkGxy4cbbiJecYmqc/jrqz70fttyVV
KkzGd9GjV/UBUpBKec2OrZaRQAb6uYMtZDEAcO30cS6+vgxR8l5/XdT/ZBJjSThE
qVzwrDH74w6HgocGKp/iR85978ztm+tPPH2WBX7hmXzp5T1o4yboP1X9d+ze6HHn
QS+zlGxLDukk+EMYaH8CtnUmHc8izT+nEbU9X8J1A0IhgquBWH049pvvQYqjh3PZ
VxX6LdhLJHoSVrxw0qXHdg1uPNG1bcgSTXYgxNv+RTgrlQVVxkw5sjJcREeiAxnn
70K8Uhp9ZS5sZLbtOwGjBJ/+0JUCl3MmkJnTxJkzVRWvVOIdGfDsCKGlFwKdkiRp
YHG8JKgyBfQm+sv9iVpXOW0rugzuREA92qhxNGorgIqfZtiN+L6mLfDyDKxpeHTQ
J2F14iaXlmrBWuN7BLpD8fMxT7t/OHmRGUza+bk6C1/FtTtKdUqJ5QeZntOZ1G/V
c0gQj0/Q2fyJnxBvo78ttekIuvhop463ufahSTcD08j7psnnTpWLyfQ0iwHrdQx7
0sciK/0k3Rk3szRCtNtNQc/l7DajN1YjuQieSniYoVWKCIZdDU5C90kNzraEqYTM
sFDMIKXCt+0+tkaxVctkz0cu5i+DV9ImZIJRJGXTgbIBXERNe/+FauPBEjYXk331
Ih0Zuzq1VlWUcGTwiM8BuQ3lWNHvEKqCdwsCDTaUh52Sqj7nspsbV87Vv6G6kBBZ
0GY35dqjaDgxnxlAYN8Mbj4cAuB9GiewFMSQyZLIVodB4ovSlSvPv0EzCvbRLD5P
18XSLl4TQW50ZCyGHSxRw/AYk5O8Lfnt8XR5BuG0rkC/N3lupJYf7DsIYjRVqx7P
QLGjaBOFIMg3qgVNwd465R/g9uzF2WNn8ieC2p/1iv370cyHsgrxXTz6GEE/iUZa
v/LbVgZDj4DsCqwzvcicQMl8HP7NphzaiEJfumQRByu05JVUC3x58zIbKZGgb1Vw
QKUH3Z35l0oCAZdbbC4dwLPlyi2mvdw+5PYHoAiuJ8g2rp4OM2ty/wHn2F7l16f/
FXpcAcHvTe5s6sfawsaf9HcrNLA6pRmv5WjxQiEJnfpqosWzJI+QSTa6e/a6d5TP
wgZ/Fccg0rwd4izTTFzSPVfebv4b9dbW2CBUkg9KHiMGERJTzCxLHt0lUvuaiwWP
lM/LUzqKFrxJAqC6c4GwJYPtmUDDyMcjtqnyglxX0hnE5AcPl9gvip4n5S1lhiHq
7DhD6f6GRtG1PpOklt8fjL11SveGHB85f/84pZskh7AvUJhqQjVmXhdfTfA3XLjl
VZdz0o1hqXavczprz7jEPuR9jF61XBw6wt6zjEDtNZgoWoAhqqHMM/jlvgYlrREp
5TABj+PDaK0XhEuy7ZgTM5tEaFj/fNDUU2TG8bZqK+h004ixSym+vvFxwPNkXSWu
dv1ZbUnEzI78of4tie4xiOjSfGlCQW3Z0V13TBJ4WNB9dnanrE7FUusld/5CiG3W
WWZeHWLcNvNjm/nOYZ3HqntT4x241evDomOh7lnPEViaVwY2gm9M0GAaJoVgqer7
hmaooqVQ4vPF0oQjIhw0W8x+sCjC7I8b8l9V0ZOhHUD8duXb/ZlHlVbPmgyFeoUS
AbhwbpylTZakXTu8+RIKRq1PewKJQ4u+yw2mujhz/Ft7V8FwiU88M4G19c/3dO8U
WEA9//UQ/+JSHgPv9KmcKTeuSD/+rAYO4ax/k6HaYOwH52Hsa7zMn/GbsurfonKh
rQgNT2ke9cD98Vg9vLno0rk90MszEcPm4+uv2vbwlTmtkCfivb7j8M6FxdGarxTF
3YcDwgih/XY+eeq1InFGdcfFfrf4ysSAUvUOj+7mPTqJd2DtTTJLEsxzk9cMYCYI
NPzTTH7GDe1Azm7szqJJNScAerEs3iniQi4xqRkwMQFYECoO+cC1dopzw9AjhiSw
n761saki78tlEcupTZ3eNMRjCYkSm6uVUNW4K5r3SmZm5pGT0eQEGtekc6dx2sZY
S0Pf2PTGuphzGn1spB7M1Q+mJsXUcDPcvUb/VLgW3KHz1VvVIr2Pj8mfyoKub6eb
1mm33SfqhCNtSlgh0IeMaAABFtQpErH8DURqhPsVzW851j1HQYmFv+b+dXnKGf8t
vCLSqW3+T0ohShZjz1JWtTgJqUoi/l6J3u7Hqbgkl7VNj7yinuC9ot3RXnhjROMz
Z+PC3XJntgTyhUE9+sVxAxlqlfgE3lW5t1OaRCxPJxB8si+eDD+LelE4d79rCW0d
vaNSHqrKwr6zyf3YJysGH3p7nK5FLXSnwzDymtExV0MdqCPu/Rs1y9SUeNNpEITy
j9Mr2XX4ydYD5gwYc1MkLOp4l2ySbsZr2QKrJKmuNxemeeWBSn04ha+gpajSwrKI
J9uFt4rkYgDVhrdsNlowsGelp1laP0qar1y5sxSsanbKJ/THpNb1fyURMMyo6vg0
AfaCf7BAkFXP0+oWTY/AoMOPoWvkv2GHl7/odaHAdL0KXfElgJ37MfKbczJDJ9mD
qi3Whs2FPyjLHLa0GUTLH6ojaJfRPTecmWLm0BwBJlrDHxhCLR3dS4vm3K3AX53g
u93fqqOITW8yFo5ULtciRJ6mH4i3r6b2cFCoomIfT2OOosz/9qy3Zcc0nVkVIbwO
g2EYq2qKHJWmwpCT2l5HLgGc7rHn3fQdLgEJL7Baah7PTKZ7slD1RTuxgWJiY3iE
ei38c6L+ZelZnNlm++SzhBhT6pE0iPr/tf5IRImlOdETbCsrxaPDJrXmd6jTEGt2
S+jQJ07ARJRq4rx5zW7trw5O2pLk4UZDCExe6nAnPYCqBzBmhtKtOI5i9R1yLgZ9
BBTJsFSmUtS4QLSS0z4YlrRQN83ZZs17Vq0AOH2S3uT1m2yihEXi9LRmKd11DqS7
ZwxWhHmREhdo9kXz8GPcvRG+AwwS0C+kbXpMNDp5f42+yw9MQLhk1lJqQ2tmTv66
ZmyIw7D5vt2/2saBlxjXKKuo4qAGWi5YzCzlzs+pgYQhSJzekuZFwwW8iXPtai96
xtIDcppfYFDGwnIqzX5v/oxqZVTTH5QNSxm2FFmg5vF1/k57qNGRk+/i1Jgos47e
BE/XeG6sb3UoSbACv6Xoo5f+js8YU9s/RDp4a6UiGIoUWraPz+Cqqt95f+MSNZtm
ZUK5hdokjM2R22dlcnFvheiN00oZRag2/lwfKtT2BgEa9zuqfmVAoW9u/VUSZfZM
5oWR7Emiv8iqszfNi4o67Xuva3M5/QvmdAaXQPooFafHw9TMzAEnsROPJoOn696R
E01trx9Y3Xeq8cRxxdO6S6pt7RejFqXaKUbbZdZQRQju+IFGQLtahUtBaUnDGGUU
LiEvN20sC+Wpqs53EctijzdJ5cDVDZY7bUAeJVHuxFxHF0u3JAVTmvDdYD//zy90
/j1fPT/BSpR9UkCGZv3Zp/92EQBLsv3rnVonzG2n09WQYXAgZPPv1aOARCP1rFDQ
qL8AlMA+e/4qQzhUYp8sazxQzXmBsy4a2UR2HSQgRgfv6UZSTQbqZZ+fUvBt/uG1
h7bA9/s5wMTddtLW+lpA7juospjIJf5wuvnD6FvOuYahDS+5ReQ5nai7b7mBkuzU
WfXUywQyJT+PxWaTsJ1QcWwJSt5kJf8UbB2h1yend6MKaHAKWhDH+dPM9eWXChmv
/eKdELxq3e/W0crQsNcIUfSifpqN/IK9eMCP6S978csT6B5Y4HtNWHSMDz1Gw6jF
CwfQwDIZ+y5bs/b7xGzdc0OuIm3eDI9F+kawEeX+PEKU6fByWm96j7MmNNHRA6B1
Y89A+2jSmFOo4d9E63BP4yXFBZygPoAvV3vrYiL1Yp1QZeDcCicWQuTp/lwQCOog
YhTmUOL3GDPFu3KHRC0uuMKix33Zfvw/twLKDGCW1Hc7re/1us7HoQxg4U6RdYHE
W9BhJvfZ7ExKx22IWpip9cEM4m1pzZOdf/uZupxWdQfVJPhAxRoWqV+KrtE7X0+K
GY/zlSrs/ByQZMos9yHZNIgF+q2ESsCXb1/UbH+zvSi7O28MYq9bDlMJCVO+Mzy8
62Z+oLMBBYH7LuT2XndH20kqbrerzIJYn+/sMh+dI/saE1E3cHpmM6xzYCNFAqkX
g8A1aEllYOGnhB0foZT8aUYZNXtvDRTCyEnOuA5v4D73zVUMUHyUYrxGi5YW2YaY
udyK76Vb3j5EjapzJuhDBLh0nfHDz2J2s4SfyQrqWknfSx0CZBMaByRh1nuDQYmx
hp2NVAwBF0wkDNNYDrf25JwA21Mk603Ioq9Y6RUPga+UP4c8n7cepkx3VY7+QJgy
qDV0Dm6HIb5IARQykyiuuSlm0/vUvZq7u2nAXOzB13UfaBf/f/ZEMNB22PtoDna9
r5wejkXRkL0euxc8499FR/OZ7gTDTCLCWfSg6fu4rl9LfBymtaPMXb+kaegpOt9o
KqCpcPA9m54nAdRPgOiUuC5j4VH9NcWEXBlheN1n4CMO8Mg3EzI8woHk1Ao/FF4l
8FNRkWXDlbvRQriAm8jEMvS8sChYeWI1hCLwijMinTpJmGIVIyerR38fRJ9+C7Zv
5qH1Ew05SgOETRgLwz8th57MfrHe47Vl6PxBq3eFRVQp8YlyGcEcxas/KcCfB/To
bkrrJTsZGi1AoshdnNuIvcX0w3+i5c7ahzxRwvy8gih0YCVFEToZec+03HkRIcHp
4BdNzIdVVd77ewOD5qwssxoM/ThpsB53pz7tMx3xFExI2sc+F1/xRexb9ZYO32sk
buLZJCsKR2LRnbCjiieNGHt8N7vNxbzEGJAcpQgfVlnKl0umu5/a5YUvG38l/YcN
vnTxBvnt0SlTlTPL3jjVyhwp7UE67fbnQ+iZj18vPhSzzSCxtQ0jS4cXLEVQkcGc
HIvLs1vwURDbv7ioGGqwDsXap11L8G23ASOPokt3k9RJFSer1JqlQVLcg2T4DgX4
NhPp2wKV/Teg9fMpgr4jrT4vt235VvWSRCDCCMz4OzVScwUhsgrm4F3HyGPFbN7j
NgXLAVnRSsvZE/IT58qE8/USuisnWtFcoVIQrtdF625DGGFRsswojMpbffMvYc8C
oAALddwFPMBMoFVe2L8fa4zySFfWGW6vtjgQD2dARdSVItvMzn9l4+VAFBVzY9m/
mM1kyM0dP90y96R9pKxN3nwSKknnTYRRny7OMantzJncG54iB+ZuenIVzFP0wK1I
GE9zhye5/HdcoDsVID7g8OPi0YqJvKhiO1R5Ia4YgHh1Cz5m7JD9PGpQnYPLkrGT
NR3bvczk2koOT9tOM0/2lOOEKdp53bN491rjfs7DIMl95rSt2Qwjs4Iyk9qV0u3l
8vwh8R7Et6IeB6+ZKDDgI8yDiFsSkw0vu8eEcuH8yQ3d56WwybAJmrvukOU0G6+q
VILWVjWegj3u3Fs1kkG+TTBOCG/Bn8IP+Vex/0Y9XMXYlg6otmOUzdmsZ4hkw18S
nWquPbOOu3scjTpJv1/u4qj7wMHeYxfxIg4jIQCUxk8LyX47cRl+T+WzJKPnOU/A
9fctWS6OEBnAPJBB6upzMsxvNoNRf19ucVcshxo3UQZSZfbE6lke5uTLEQ3lXe2a
GyjspVs3BVKQK9cSLGzZaaZz5JhydhkyiQW9Kd8Ixghq8KvMg/NPedHtECwdPCav
F+e25gMHcoDGFVZ6Xib+mpKtLgPugYiAAldy18qu9tYDDU4CcBU45QOFF4Yi7XCd
VEtGN3q9t1cJUtfESiLDNO9PD2zjpLGe36OWtj5B5+ALg6DcgFI7+WUJkkeLan88
rSJEYuuZaU7FRU49PeVCLRoWKywCO8kx1eeZ2IRZoQTPYhR4fwlvjzxAYIhxz7/K
eeJ8T4C1xKj1YwAqJ7xIep5i+5toMwBbwp35nvnqhebZhDLN85dHqoTVNPKuVz/S
Kt81RklQAjTCKpBMp216mbm8+uk57jl9wqcyQe6gb9lgYbq7tq2JMzjcrCHXXCUQ
Ks2cUOdeU/FGU5qfAiCjZSn3RBNi96TZMM+Pdp6Sb8EEP0PMh9ouQz7rU2jTWoGq
rW6Sk7O3TeSxhl8ywz41Gz3vax3GtJHoc3/769ynOJSN3trCwBsWgreY9monBROn
gh9YBO9SKj6SYhvHBElL8xmNa/1W/UiemOOyx3UAH65xqSVjUuO8BN7c3F7jgS4q
vyEyidgx/QKNQeIEw50Iz8FN4niq6yFM3ErSaW40PVEXOt2kHus4Yc6SOCCS/uVU
v958kgFXi6v5rfyskGjm9I3rZcUBqhLS6JYpbUSKzEPV3RP1iKKpuVExpRqQQVEo
2jbSbUUPI6QfoQEm/nvmAqytaejv8mc4EIB7dCAqZR/X/lCr3UNGFto7md6qCVHs
WNZ6QBmKMgnR1odLKDZZl13hGSJOw/WScl3lBot12BVPFKCgr60Jv4FR9m/Va33a
+hsdYuyyHuECYfR3/baJmxra1NbppJni+8D0F4yFJE0cjH6LojuV0NsUGfLarP2N
cmArz4lHIzNCLveOieTa4HTUwXd8ZbxIhqUwgHByTwPCYeqA91CdkKPZ7hCueUvI
CnzcGknXJjbDG2U6uMOUUaTFC/VwjnGJjO8CHkmISI6HAvE0ndN+e6lN+pdjHSmm
hRWuVjwF/17eCy1REsNxB6of2kpCvGZaJOzWBSBxqFOkzUkllaVF7zHTzlaSbz5F
aZBEMfJsUrgvgjh93LZZReqHaspN0IIm9dr0lc0JRLuacV7Ho0DugJ9oJX3+86ax
lJWW0fBb25WyT4jl3HOm1p6x4zIyDaRbiR0BamhDyJ7OuPPjKOxgvtLAdap941zb
RoGYVYsguYDrHceDriQVpKg06m9K/euVfcZb8NkH5ZYrUpYnE4hOZ3z9BHlY7dZm
om7YZeV2GPFb9RcKNlfa20j41r5JfjSfsfX+xcRrK9stVWYMcxUuVoXBB78KSKqz
+wKdCHydPWuRVfx+B36v9+h6ff4TGK9Ijv/LOcqmHvyrDxLE52zbaC2M4+6XG87/
gFf1HrznuzNJQjt5J5f4ZOzu7+cvG4WzFnqYRUgOhQuEenH1eH30+PKKc0MFd580
/TyH8Go/mRpWZeZeW1mz0a/T0ZAUzYAzj0MjTXDxFo/E5rf0iHyVrK1yU2vZCgLm
ics2bA4sH1wUY/zInVN53kKA60NS1Ah2LUcQ0KMgPdUiLZJhmLXFtiSgNVsofG5P
kDNj2Odz8SGh1Zn4WmBt0XK/mBJ2prgMVoedj5zi1N64bDfY0YAGUBT9sv5wCVi/
7hBm1ka/NnFzpVTpvbnPYiWCrb6fkpFOWlQ7QrzWVdqYlOn0hMqM5FFaL0FzvgxB
bUvGz97WpJOAD2HpvDLL9B8IgZhFrfvLeiwn8DF/v+q9eZounuwWLCms5ZO6RXjJ
av0cw/XvEknRLV9PVhogNWB5ZHIpK5sIbvR6IEn1ji1lxnpq2AEkB11NtFwHVy3t
Iu37sm0g+qWTTYYRtnhQjg7li6tSq5TBNw9MYxC21QKYnRN5FOf9c0TwrHYvtgOu
nTGCiIvR1HPeNgoVehdiJByLTt8NAF+LH4a/nP1U6PDfWdtSs35ycuOGECVGGvxI
sht9nrv4ACeZpBBFZrif9UsDAa2Mu1mxEG72Q96xhUxjWyUEmqrNrBkfz/MYPE5w
TrKLGQpggwGBp1Pe0ns7hfL1Y7P3bvvAJz3bdcY8AbmjYyzTyEl3Wow3Potj7GAB
ojM7iP9KklHfMgjxxLOxNZaTLuo5tSUMvzYDct0xqNs+dxePj3A0UIozNW6WdPbD
O9oRIF3o83fmUK9Hw2buLZpqUwxEc4uCBjv/sbJmbW+bK9RxQugsRNDEufqxy4sB
YIGqgy3FgT9SPuBfr8JeuwE5ReC2GMYaXXGW+CloO1sL2KksIbQrSCxgZHiht2N5
A1vXNJcFQvKAfLc0RJDajjW1HEHUG4+OomufPI91mXi8harL8Xoei5YBkD/q2DPq
Cofld9+wrfVRBRywOxNuFFEb4zW+XR9/US7sKXgxwdZLYmBbNCmwztLPsmevR7io
tPhPUJzZrWAm3yx/YbrONwzUApSz/LPredHdFtynGoYof3B2QkuPRZksSjeS+aws
OHY3ItpqM/GSMDO97FHprPdjwQRxrg8XsLRcwD/l6voKfUwWFIdXcNPnGVizzvqd
57pkDQZc1b+fis2rC0sEaxppkSNreCLrkHHmtuxZS52Qt8+cd42bWHfBl6CMP/fs
vYcpPFcImbuYFKr/9uS7Zf5PWvUtpydPQkYyQlZgoNO9Ue5xifilJlomNBOLaVcV
dfoxCfe9exOtCrVZ+nHaEimOU+2dl6geg53gAmuh3Q+KcBRHST9NRaccZ10y7NQf
UB8uUcnQR0ZVBalW4l5zUpSUDsXtciahUPJg/uwICoIvwNzJuXajfA9S62z1Sr3k
xkKj+baoyWUysp7o8OaYspcpzB7oTofzduPDVfiyRBc+i4HiLdbrt9Jhi9c26142
U3tKxIXJqHpwgFt3FCWdk7uOwIX3T97lC8KnVyWwrhYGiUj8S11/nvIkoI9biH+H
urO9K1DcvrEe+O4X+xGlMVE2OvO0JkDBQEn2MlSeL2tuy1jsCl4loxlPbFHMMMEE
Jkfd2l1sww7wbpUKYHMSQ2aOsz+xgi9KM3Vb6UBJkrw5nuCt5P78taamhnj4OqL2
nOKGur4wYSa9iZrnTxDJF7wyfp3wYrNK2/PkhXLt5PLSNSvoIJH88DPZ5Bq8+Tj4
g+JWN9zWkIa38ww/Ajsjcur1Ppq/OKcQIr/Jpbzk5YpiLdV5dEhUHcVO5hXVMWKg
IV7CUD/ONPaSyyLs3MoJf6ITg+6CN2Ccjy9WhhxrtScYWTFG0fV2a7oX5BgtVaJH
+fz8WfUz6WD2bsdij+JkwcLHvUx0KmfeX8r4M4xuKkn2oky4xpdcC5FqaUZIZ2aS
5loe5kDip/1Lf4H/PHJ3A+b7Ag8qFKkGWcchZuY6h74WeQf4g9mWcx0nRsH65P8l
iqVy4ychU+FU4WgLYTQQHOAjVMSlMcquooWjq0+p43V9LGohz/3hmom7O6BIhCz7
I4/WYcS0tuCTqPhmfa726BzBPZaagWjvLJQnRAELdwdUHgPvZrK3ftJKU79qEJea
ubQp5xsvkDmjuPim1QR3fHLKiIxsr1pyKaSKuQ9g+V09i8Q5Sdt86qVymgNMVhbV
9X7iLfKSCLl2aHfPmnmIj73MWhDs+CW2TAb6gDCzyNvjqoGPM6QVrMsikFNDJVRf
QYQk3hHK6F3Rx6GybALdiZx3MbrS7J93bgb6joPBNasIK33DhfM70YQUNu5odokW
KFAezz1P7bkD7DDxECg08kIvSy1DS/spiPMnOBLT9qJeSUrHrAZzjkbXS1Jg6fOp
84Oj0UWySPCafNuMzK48XAJI3CSM4nSxSNUB9D/Okfi3msFsFKp30aCnc1np5Rgb
pPySBl9ktIWaj+yW4fmjI+EzI/DsXiVoqmcGH/EFvvjIoMbmqSJljK094zAvib5W
c7gNGXmWFE+/Pgrt3779sJ/Z1Kj3OPWrQ8+ORL8Clr/X5Y+FjinyOEkEtr/tBsMy
OuRH+DMF+xYxiwQqGbUniiCele1B7e7wjyVcnzusjM96dK4Pj+MpA5iAcjLBfu4b
JT5dzkT7+3cJnO5BpbbLeRgMm6VVZFVx/HH+xTjyGH6cW/99Ux3caAVJPKsj7K77
Y1FthG3ewT35gFV9h3Tunc4X1csAfnkpx3gqYTNEsUoXEyHWNoM24PgEd6PB2ZtK
ZiXAMdBwsbK5DOzNfq6Kty2EingERP/lKvxh/ZY43CzHasKzW/ksueA8KfMiJPUq
H7IvoOVM/XEzxWAd8++GWRwuCmo7b4USUALr3Ykjh/3aXyvT7xwul6W5DXtf+Be1
er+gByz0UXUEKnNinmyLgb2ZuydwCnxaPBKUKpyH0m9lupTkfXzgyCyws6zHNk9S
3N37/Pu8fBR0QJVck0lyGGfN40ebl7fip0f5rCQjVSvouH0LXAaBr/7UFxOayFdP
aqcS86eQivpUsr8CcujVEl0qXBE7Ca9nGukDTYbVekriT9dlrbf2Wc7uaA/N4Qgl
C5m1uhZ8RzbBscwGZ294iDFGN0Q3OVh8RP9i+/peMn9LXCURHQr9koYlREUtHkot
iaGsOE9lMgxbgTJR422YDQyonsc91D1duJQU0m730kF4maVe5i5qsAsvgT/UeMIl
ZOAcInW6aEgyy13Ete8daEzJS5S5xo1qTvqPFQ0dAmgiaoGvk3CiD750t9vGsQ6a
rawkf54KeaceqUgva327lctjw5LVT7ssUhhNEdniZsL26IGCClkDvieV8Z7eXoIL
xDg2V1Wu9PbJ+21pz8Bb2TwhxvrpsRdSvi1h6U17/YwIO2YNjFDwF7kBKIiy4XIF
ljSKlJbux4Cd+TpYkubTHgBol1JxO9ZmRDFMohesjuglIPW40SswvqOraSw6Pb6o
V1tzWOInqVUREAKe7+24Y5hRoWyJgOoqw1svbX2Xkf6hzXurwfNECaO/fi8KDgtk
WgmMR5MRfyOyr6JcAYjMWw4UwEW8B2wOb4z2Cl0nQjNBNh754d+gKgVvlISHQbak
HMAlZ7eqR4Q8j7LT5KZHpkExLainv8Tq3G04tLtbPZIGBsU6Fxfcsl8OFBB8f/8L
qBkpHmMeB9ZMqPj1WYVXuwRBfR3nGndOkQwlavckwI8cTdMuAwtGaCVEc22T/Prg
kkT+qBSyUy+P+f8eKl18qfpQll05Xeeyks/khQUv9svkInl0zr2d8/sdThvHI6Ul
OsWmqa+x9VkS5IMn/O9oxTRtGgWXVHBGeUf8v9weYIcW6ljG9KlNUc0vDNdk793S
MSVmnyZUCmo8bpV+ZKuuRKaPajj7N1HJYSQM0Ij34wHiB303BahlsM6YiXqNjC3d
Rj+ucOjqix8A9yWfjiK6vPYrHelY/iJMQx+/EEY5+ebvcPGrYtYJ0BCRwOCNQGrE
ZfuiI7RIjSfGBzuLPMLI2UIRIGHbu7RKdlek2TNsFUp2e6IZr16G4EQ3vxIQeK9p
KgOnKjQnDlMKQ8QFPYN3aeFP3whHO7FK43vTfUEkeBeXLiwvORsrRDdlPPc+qzYG
S1DKTwacGPUvvUZhNKqt6+6dTndMQAgvzzWplIVTBcOIf2eiE8Zat5inTwpJHc2T
VFLPxpeVb7MWu43SNXEOg/MU4+LJ4ovIOgU3ldfG6bnweuASfzZ6srAXpdFKqIHn
OyyXoh8dbFgd0pqJpACjnSIc+mVZUR3jxEvtF4oOVdtkApRYityXQWC+Q4OVUPz1
j8gDRX6YHCaL1ZtipnRXy7u+undwoLxIaMBECgNjrmoKlf1x0d6KWHPMetcwQT6c
D1Bf37c1sZFWpv6FV4x7abt+rfyl89KXGcRsMhklTzIYw7mQeKGtt4EhST9xQj/u
vwdsFOBuZZaQRY9QYZHbFeFbYeFeb7Gkz4SMeHekQkSjNeLXMFON+k/2BQ1ZirvY
WBo+Pt/ij0B87PNIH/U/rkzhaIu3vPJzGLFyiBgiBtd37PODnAVe4/3cyMkr5aa3
dENQ6GYgFuW1s1j7yn9hEegwgjYVPGz3eLvTh3MNqRHz4iYgdy9HFyTABOZR45Md
ZS1LV1+S9ZcKz4j+1a9GyRhdC47i0Q3xy9w4YvSQ0rKLVh1jQCKBg57beUeUk0ud
xAfY02fmZkIYy+deiOnjsnFvA9v/PCWKBOAv7wKlpV1sDoIcWXts9HQQViL0pZ3e
/BZJjQKJqoBBxhoeGPtBB3+KZeeLFpihOqKDSC5v1TUT8cFgTi8nmZfA4uRbVY5m
pCxwzT5BAQXZvR8dv0Yvkhxnm8gdUj9NsCmsFs8lo00K1tE9nfCvOmxq7/8fm4oj
7c8MGLj7v4ZeS7Zr/c6HoMamI3k+GpQQNHBGQfcj79CGiVQU93Wukt8ejydGe2zB
8bZhahN3DAk8VZFKUD7C6HVkmqjZyCMPVQA/tKpV7nHsbgnztU4Wc0pAc57/+w+x
4lU+mKCMIOTfCgBu4zpysthBM+uBFFrDENo7h/lAuG/+HFAXdbtCycRr5a4nRVnN
thK9tVEccpUZsGXq6iKQdaM8eMC1Q4UxvgJ678/XiA0LIjPwEayp96QBvwJ8mGvX
PcF/3cdDLhFMkxHiIdwyq3PVbmsebj67XrlUdgCl/rkEiQsyLaj191EBq0NtQgeu
aFM4nFcuco7obJMn0oRR164tlWoF6bXG2c+HRzJg48PRQCefQPNcRDKwnspr1aJ8
F8prYaviw/0auQznA/DlB88VFyQTEB7UjgQy6FuQMhYPusTP797mjpP8jJnY1Rtk
dPZfmq9M58KLi/7jimW60ybDB+X1HWk5MIlODtIVGDAp5+F1ktxnm09FES7cIyLl
5xIJ5/vbQXIWUoDR9N+yZp2y3kstu23xhvsVJLIBKU/Zh3AD9LTGM4q5OhSkaALF
KUmFh+6Kz+km2jZWSPZ2WJjGEdq+K2Ly7gyEjbdLLnD/2Sl3JyIicTphZ8eHUTws
j4hwHl7lEVjHxSB8jvb4iJ+kDOelQ8GlF+b+tvh3Wet0hmXE6cXCa3rjqGxrPoFq
eNLK7KQ/wqYkzfzXcPaL4WXv+Z47alshEBzvy3TyA1li0KyhWd4ll8HFEsD5r3F/
yaZ1AvLon1uMTD8VRE0R8EN3DxN4CgCkuIXvrgYMMjYkpNr/7dAftnQ5ueN4j8HQ
uo38G+VujsdE3MZpdCVkLNpL2+OEwwjtm7+5lzL9pUDpgJPCPXDE7DYWKdL0x9PD
3I1iZlhTtGG7jWeA84au/zBbQf4wa1NPDNrP+lUA2cQ2SExCZBzMlIiIgDNlW/Mt
cS4/2ilJd5dl4NgVnppAn7Zf6CCa6rgkt7OpWAs2MAbCM7j1+PBj60A7WZ3v3vKT
5VWWVsm7fbRzVOBgXVrNhjP91iliK8j0bRub5L2jAyG9hXK+rW74i025MPDY8qBi
Ok7tbERlDtGQs4jnunopLKTkCCHfPnBmN916czbNHqQHZ/eHDdue17IuhD6oNmW9
aJmM7PSym0GgEX+LQfqM3SmALK0FNOtpbK2+rJp/kgbZFRguHRERaVrQodAwPM1G
UzkZlBM0WQDT211WsrO999SnWMQKah0ivRGGlyMJiUCCBfpLOciMqXKTI/W4+hkV
idRNVTuDOJfwWXY96pBqI7sfTmtEN89hWdyc3lFhZ1CTgRLb2yu/k2NjddCOblMk
jMqoQgmqj50uwQDwoR5S3r0lYHm2QP7vYOgS/ev0ny6aBwM0QszU1dbnrDcwMYFl
dSTZRuU9fkCVCgB4+WHnZrYNU5m2JAz9iUI+/iho+aiYmlYP3zld69LJUQY1sf+J
+G9CRWCxDJ8qAaoTFNoZnztSpbzzF1fxjdRfeKoJOYH71zkJcLK/129U4dq/GgHl
QjQpK85XdtAEoDdWGjU/LpXsEvTNdnPEotV2FfZ4Jq+1n4TARoYXG5qiHOIrhqht
iWyjpwAITXNEjrxHWcxdV0dqUOJ0mdFbGUyPomAGrM1rw3MCfalTMT7Un+BRw/9B
DfdTnJVZT8qEvDZVhaR95s5fO7qdQX2vW/CehfkK/JL/psHGpchnT3jag8A7AIPH
90NAiuEseuiUkYRL33Fb2z1X8LE3J7sOMhoaj96s+BUfGCBfPrKfkskntpYI83Lz
N/SMf9+AuqgKGYwyGtGeJ0HkLcvQeOoxtgFDfcyPjO5L5dMfzthaKOoPUwtzLnTu
1VpHTDojnqdc2BlHxKnwKQijNUwYUMdHq9g2SlTtHh0NmFDxzGYFL5YYcLvNd+CL
2PEWaMk+1VIqLx/dGtV4WOAz3Z3yPeRqYxBSS3z+cZbA5K0wuyKLRTchaohdSlyl
PI2Pdy/ETRJ5PNWh83cgRkGup+KNCSp1AenkLF06maO07OY5yZ+pBWWnev9dMgXO
3wGSdIpgCRvVRcAF6XA1AthHyRPFxnjN9h0AvsavhZ1x/ZPxd6FTmDjH78b2I32r
t3mbx4DyQWUBDvVZmy3yw5VJidQZu8QsEvcqzOKJ06Ks9nOPo340CoTy7lqBVmfr
Ln5INywtCP5gUZQ3eRCDd0imZwiyvgmU5Ebrk7LRDZ2kN+IvPeYN9rCWRCkT/doM
DBWS/N7dNMxT4tNgS72+5xAZcV0TDCl4zbnfvOjs5tzElzGXqM0lQIGxN4S18zwo
h8XonxADgTI1XKBS3vP3XHF4naSaiL50+VESnfmIavrcB6lIFl9p1v6UcPssqVd+
bSUseJIedqVd3btlq2Glvf01kl8ulkVnmXkQazsRtcz46iAZRV6EHl/0s65seGSH
GEe19g1f5xjJ6LhwAG4Xf6DMnk04QA4ck9wlSHN/MHncxEvTFaDtXt2Mp8WGkal9
Xn9LFhv/jl97b6co5S5NE5rm6vMJUbb3BcOi9dwLuGMFdbW4D3J8OdkRtNH9Gk4x
HuMW4EAsbHoZ/5icvnIOhMzo1NY24R257dNhKYeSQFSPW8wxRpIHXApDfI2V+zM7
S9SRWsJ4EBS4v8IH19YBQ40PWjbd9fftQnzQ8nLhQQq1dRf93cYnVUTpAj5dEOqa
N45vgij/fs+WdStBWLskf5jUCJ6R/9Uv2Y1rDS9lWkkdGtoy1bFJeaZnjUGzNbvq
34XYDYw/kPy0PPfBwYwSTxDQcvXwpEskyDCPUiFRl+oj1xEsiaEWKAhAaQ/uv98v
BknzZ5K+6zaq8cqyCi0wuu1YRUljvLe8a0taUiF2SOjHDGQOQgbyQI0iro6ND3Az
hJGrzacNGpeU1aRj/mbiz++k/THgAckaNT3WlWvRl3287YhvTPLWlc86+ChmEnM/
qwkwI3PURQiqLx1PeZWhMKzLEMYzm+BeJ3dMNFDuUXocuM5y+ZhwPFbBJBdL/WCz
nbc5XF1i9+c9vWEoYGKRhDgOhn0EEShTyWC26VtlMDlOPSkFXbj7nirRzFuL8JS0
NxQQ6ArhyA6xpqGrnG1sOvfBzq6vWVM7uFRukdVyH17X1bbVYtGm8WUVF2QAXI48
vY2gowMvurqBgGZfrFT3BeDP0yNMoKBNXVWcQ9fBLvJUIOvWG8TZZ6VbmQNbvtGA
poz5E6B/Q8AC4PF3ffrd1nyz1O1oU9C4d26GZ0xTokhlEFTQLtQUajSTmESys9yY
L8bJ9BK+vTokyBkONNkY9cZHJ5SOqA7AnMUgUKJDruN79mjaj96FYbD7vYB6B8Tj
IrLs1ezRMJBV90/ef3wom7vl8SmBjTuJji2eVNLHH+XL9DXUzT+q9bkNxpDxXYyq
rPl93Mn4pUR14WhU+HOSERxVFqWY23cyCx6gMmQe+XAV1/pfvR8UV/8csQ9e0oR5
oqjQXLrvDkcKV2Ip2QSrzIQkz8h1ZyQhI+fbPi6kySgZXsG7q9q4cIOREnjwYp0B
50oxfg5ffHpcoFk8/32jsoce1mCcyZg3x/6SAsQrx58R+7DHU8fKQDU3t59A+wWW
LE553Kq/2/p8nXCj6KTjRDuPRnMK00D5Yt30xvIoU1FnC6PvikWS7MuZH9LbhF4U
Bp/SPNTxXMEy1sWH934DsaNQ8pcZyk5g5I33IBV7w6kPi/gKYFlizWICdwadeJDO
ES+GTVXMpIgw+lqJUn4HtVDTO/gqtSyu6bjcElbQsFD3SnqbmIYmzgSjpCwNquo6
wFFjqoBpusMEnsU9Einhz7232mgsimTmo2umWcyg5DkXThiCWuYoFsBUM+Sk7zr1
61NlXp8kvUikLAujYj3tK0C8ZvQQkaVCfrdVRa8rtrk49XDyustB0E9k8aD870J8
SwMCZVJg9O1LDQP/3JsNqfYAY3xJHMK7ImK4NABNGaZcoz6ovxwUx+Nxvcy3RBjT
02i441EKMpxMCLSmZwVwP9tOSd5ie0ouGAfnyMoqAsNHPpSTHA62gQjt57E9dnMp
zuFOvqvMTplWtTmkMAsFrUSm/zkmbJkbNGKQ9XiHIZgD0PHsXGRKxGiXzD2lgf2a
9UgUGQJCLWUB6590eB78R+Vm2pZNenmnwuFR0O37F655WUVR+CEfoDT/BXARsDBq
y1/jVUSC3pbZ6gT1C86RTv7FXS1qOWHsBS1G6ODsEe6niPqFalfdExl73hUvzyQR
eduE2KycUSdcI7hjxdrnvHzOTLf6e7MmS88OuUlAg3Yk5f1BYUQ0TJz7q9f6jy/f
d+x7KhWPN61ro85CdGSy0KLrnO1jtV/bydoJv7H3DwtzmdOKb00K9LquKE8bqwnt
qNV78VhSYJ/dORgfDwqjL605qMPOqRh2RCHTSNBZuC06RqAJzGaGqUxu7OP5+fsu
GCwOv/EqcPSYioqsBkMK28Y5QJoUwqni0wtGPDQshE+8BHVrPKF+3YMvVtuFD7ps
a+SOYQ9VStwQCtUSq7xlHq6BSQtNhquYYHRTNEEUl166FjH9qMuicntClnx62oTJ
ubsuheld8R3fKzxJZDyXiIpMaVWAPMb8uHPHNOkIH/SsSpvELd7pWdIHFrMjP4Ih
et/c6kvAWc7OuBjFtwNLOxHdpFwQPd6BVI6K3evnzYuzn/a0bVXg2z4cv0Ba1cDu
UiH3m4PlNMAykhiIivL00PxA986RM82AEEIOGIiRI3Qlf6/wKiKU8XC/afthE/Ar
gHAUCSWvyYBer/79w4GL3EkozIJjZZ5rvuqm2GlIqm10rpYxesGVa6xKkZIrHwgP
Lra1mEqEpq9gFImvPtBHaMAzmpKLvQotpXI82NUofQGS17M+lbl1v2cBduk/ZvxB
gF7GZ/QNhJtlCme6PiCVaEth0PiiBJVm3tmzDpzqQVq0v39236tjC0VqYGMd8hQj
4+CW+Q6+PpeTBWHY3qKlT++YZ9BM9q+8t02m0G8LzrP8iI4s4EupmrBVERpEjXsm
3SRYNzb0l49tZRxY/jSV1pzj8ulYr9qBNRz3wq2nra0YklNkZPr7o1ZPh0fnsvYQ
eBVm1xlPKR6me2P+J/Z2o2frHpW7A6q+oByi80+buvxDk5DDY8MNoSLiG2yj00y3
d4lgWsQwz5moNV8oeYiOrPYs5eakGCJ+KWN9gC266VdhKKgmlH8L6Ljp9VoQx6e6
VNNLulzzSoBEStwOJRQzDTlsVIgY6ZufyRbekUqiunJiwwI9m9pO0jUEa1WgisVt
m5rbme3erfKSig/Vlor+V0tbjwkk3cnb/XHtUyLID/116uQo/+YkNJVdXCz0Tdob
9Cb9ZPS32kyo1s9M1d1allRrbVwV2QIx9c+d7bkaM02WFPWFZXhd9byp4wEuy2vu
G8IrSP8ZnSq9wNo+kGRFd5Dj4TXk1l+jdvOazaBlb0LCWOzRsNcdkPIQuwHPtgny
ywHV+MNW3/DaCKM9GFgkJk0TOT1EgqTek+wyPLGT+2NSG2H4LupMsYlIkD5h0jp7
IGru421/YhzZCAS85PyPX24w6FI1s5izpUNvfnC8Mvppq+xkIbDa7QspV+9asN1h
62avf1p137WOzhZ3OM3qEHciZgoG/wwGPZT2wppeBaTvPcDNy6bH3+FPokF8BM+n
2zUu2Hu8PUrtH5WdGhYnQyrgmnkUZ7px9zr7WgQ3t8bedOfjVbVuQsKzf5X8wZnO
lL3QptBTr8RD8FypWuBrxo4Tig7ITozrIdDAteJuHu1Bvx8CdPqyYOMgO+98rKQy
qWJAxlD3fnOv9pstd/36heJAyOEi1orNRfdgk4MXwBoechOT93F+q0LTbVbsF1/v
24VR6TE6LKo1hN+mUIJcnS2Uf6IcqLeWLCvRQ4cjNlXLmMYuVWfKQeBR//tRysdm
7OD10TjGNM6hguZJUjMCucfGsw9ithZGBRshk/PQKFgyVp751dXvPVYrX8R99RbN
iZeUESm2mkg33jGKY1wqVYOU+dkHgK73tMvAUkKRpsTHlb5iSN3RvpKxvF4tN8Fi
hB0hWC6nSpUYJiHUceQQ+vzCyef0p4CKZ9dD6+/6j3BHGEV4WEVJDCzzIGtgp/Hs
g/D2WaKc8+N5xmmPgIAGmfTMfcwmFau9PMEdNG/woUVdM+r4JJX8/4rcRwCmEZPs
bwqgoMRJ4q3peJTDC+sCU7acfmRXVaWAzrCRkHMkbcSV2259aSeW8sIyTan3xMgG
D1bBHikadxNAPd7aANckYcW2Bty9taFzZjFBndb7ZBmih0px1cCuitUnz/KlxHTv
HR589hw5cbs10Y0xT6+1mERekcumjsInOE2c3uN7WJ80RRFaflNI2cm7drKn3kyS
GTRwyJkny4T/FrYmOJzKRJEDpACI+BRGznu/5IJUPGn4gmh9kPp07bg8cGashLDZ
IhO7VNuGASQTQOH2CXcjiAdhJKE7WBHhK38aTfPmh0vbEXq5pk9YyQDnVis5kP7l
JKS5YxoBMIAjdKPNTS/VcHAjLprvoKdvJVVU3MQZB18tKcv3ozljwF3YgB4W/GXN
sOwD6LF9tE+16kwkgOIYzCgv/b0r1OHkUrmjZ9OG8AQe+m8N0QNnO7/AmnMAkR9d
4+57Mv/pxcs7DUKZA1oRJCjbLjkfYcLP8rjM/9UNjgJrLSqlFYGc7TweZP8BZlzd
UhZ34mQ8cJStqdvNWb13NJcr5moJ1aTaJsstCwMR4FbZuzMsQXUlu9IimNqk3/Oy
ZQadrc+hduka0LUB/AmadCwxFG9AaEQFxAjhWJpg3jBGKYHYUTIkBlpRZzPtburQ
aTsTKttht77nk2Dzkber4ksE0vZpOnapsFvh2cUPwIC4MDMib7qjR8l1/DC+1AuV
wLFhoUSrfV6vkH+4AqaAeWbo3w5HOwHQtbkdWXoxnNuqLVqNly0g708NAa2WeiMm
m47mkjGC5UGykgxTF8UsSBwKEkDgD7uSOsQjmZdmLvlyoUeyuGWEBTQIBxAOawU5
wMgqPJkz9KHTChRHlFWWucY4QtYspKHKSem/7GRvjTHcTEjGFPNG58weHMnqLxZs
tkKpZl5dMuRoNdfX6wYw4Ey30BIZqmqLs3m1dzTuYPAzpFdGb1s+HV+qvZ6Q5bVt
YzQC5Pep7wYoO9Vyl/FR6okLOkbUbeKjxTmZz6ozExSb0HWsmGh8n0zNfI1Zd1Am
EG+kTem/BC7n6KiQR+8lJP1s59ic8ffDCasHg2U3uKfYXVM19SFZr+h0DPaIf7Nf
z1zLqxXDFnhgTP1RnuwQazMjeUuGLyD/zAUp1tOFYJTtLcx3VQCbQhBQVCMFJKgn
9yglvX+P0CHjqUdO8i+ywDGNYDxGgY8aUkoPi4+3nz1eUwXT/1pcldinyjpRzZbx
78zH3OHIDBe3DtVPEDi5LxktkL8f1LHVIrWQiJW20Ot0k5z2ILsemerfbGpNaHsh
R6QEVkKCAkhMJl8tml29Tzvaed//K39gWLVwYJ3k+Z3fVwCCEFlTYXt4iFlYTEPU
0joGpqYIDpcgRulKhTUVy4JFwkGaef9k2EMeYp5OT/U7doRil2XIRhNk0aWIQK2J
gl5Y7yyakbBQTeFFp6UsiId9uIWTZsoc4mnPy0ya88If3Fp5gW6I0/0/nm5oNu58
2qo9p37HkEpkha3ZV8pjIDuGdJxUB68ja5jUuhyjyt5OnhHQpUdolTAKRCQT3wFM
t2EEhNRUdy6KjFoYO6/T6fat22zgXZfGm4kkUV0tZJ6M1SWyX9iVpo4wV1/Vat+C
2wIFitaygLvvKIyTuS2j6DL5m8yIhsk10T62fxrPcumFtMCPpovJXlt83q79Yr90
OnSTDQeYJxPw3EHqItb+nY0rUeKXJ9awUve4kkQkX5ESqH5x3ujOmy9X4gocu7MF
WIllGdRzMn2pfUW0dZpiTTtOWY1EHBsgB7vGY+ET66ulOI7O730iD6aI7WrsczT7
WaqS2B2+8/MA5TLtYlEkiPCOQHhNoorR9sCWxwH1TjjpYA80yAzEJHnbAI/eK63m
TKMBdUqIq1ILCelDR1/Js4ZK57cebrBLX9nN/yK+Fqd9HUgAkRxkJrEvEU48Fwbd
hm9IewVHrNrKTa9ZnBQkBdLVhZ3ks+ZBJlyTz/NDlOySdCKxLxy8Af4AsVkDd5xy
i2wE2r6je+BQAUSB2D7yCGKjkhYyz1MTENBTcb9VZ94md8Ndm8YT4SUKbkdg0ONb
tKPFPx4CVtRLbKfv/lTRd34U5HvlIKHUdTZcAgb95kRZtDfGEypC7ZtfzC9lAjAN
TeDeLERYIxwR9f3mhu72EJ8ywzxKgE2XqTFvdE3BlUNF0n2IwnA0g83qWzoJsf9b
D62k35YadMdSl5RJKDdqYoGqKuj9QuwKAyYMqGYSWHDIJRQT/zYatBOr8WUxQl28
Q4macPf73VSDuorA580IyBIHpv/eGkY9u//yC9rqxNAgDsZ3dbcRyET0sbLnCNav
5YBWJ/Tl2VHks7THLIdpy95yLKfgaTlxygBrmKGjIxoJhOM7eDou9FngL2gaWoMd
obk995ZGDjGh/ctsCCjYHRFk3r1eJ7xjGDJvqlRss1uwJ//eHQnyOOeJdfB774/7
O2w0uyWOWeR1mfFC8i/wSYWzTSPKkNpGjQVTAnCEQlOU42WGpg1IKPaIAvtY9gya
gG2hJc6UQGlUe+Ywrart3gR/QQCaM4wnk+4jJC9k0sw390AQZWSllW1149eSURcM
T1h9vh5f4Zq1kbEzAxH1RnahXbMIDOxsNhJjt/dwChxFZToj7NLziPYuI13vr5in
LuNYr4iJzpLUqNmcUDVh9u7eRzTbw65d22bJWqjoQcPv4BEcZ16aERS319qLowCD
TWPvH9pTj4GR6joccNlD+62u+eK/WRbaLHOlsrYif+8blhd9tX93LXuI3/u1CfRs
rDHZlfONZFS4bRhwZRVehRXP1S+32ru9YhF4DL5k03Cir8P1tials5DDr2EDvAxX
GW3NRof0sUn1UiVeA0bYWkAkEO6zDgDnATFI/xGE1j/oxhmM6uRZFEoB97GgS0pS
hyuaiA7j/TyxL1T1tIAtao9dg23zcdubLsrs47/s5sX4xgURGdHaNfpJiXvbAwpo
09DyDmWUJ9S4XSwm/vxUwzeZBetkOMQ2ntpucu4BOtPdzxvyNF6NB6FRQzJeTg5X
OtvDgy76lvqqJGgsvano+nLVKN/KxRpXoOmevf++msXe9pK0CTnvDbAh4+1gBiIy
4XCQ8WT6njn272zTSYLU1RCPbGtiztagC92VWKIa8SmQiORqJxxOck/KVLyB5VXt
tj0t2V9nyVuOiYn0snZhfTbv8ZZctGWJ1bPRYkUuRZgCMiVUffXz+6OiaKMSIi0t
+ya0qJT9pNmUO8ubKUQondQCJmvOAotT3/tThm3m8jS//IqL9KqZQouwdu9BzTDl
VffuLLlNPOMrRHRc8UAnkRr6SXcRmS5m+Nmz5l6rRzoJwqTbPdud8XcT4TwqN2BK
EkzTYpjgJOK2/4aEXBHp/bp25NeFZPJtwi4Ar25kFYmusPjf3TnX2tdqb8p0isa4
uJcjk7yugxxwFEH49uAE0GQhCaf1jOjRt4pedXa6KVZOmK1ecQQyBm/6cvRgGdF4
gkd3MtW662KKicfoG+QKVdqDLaJscPTvfBay5aCbLFcSvVfsymSfT3iw/ym+U2et
9ZfUR8Ww6VNjjHh9l8akTfttpqE8JnsPX04XqMhyUuBKSx65W3iEYj37OHlebP1d
Uy9DdAP4AdRviFKhpVuFHOEEf/VGOy7Oo/Z7gYrhczYmV7Czy1O8McTIa4Tb6mut
vyojdHeOvIk1Ne4s/TNJKW82jP8q7PI+qwaiGR4Z2fatacD4q/GvZ2u+qivn4086
7RArNujX/A/xeASmXgBteh7zJUdf3nu59mdmNeG/VZum+TrbXYbkabYiV8oLX9BL
6FNvC1MOVME4trdTa053kwpCQGedLOTDjYcyzaup5WwBVTV4KJ+Q57WnrMLZVFi4
6iJtrXr8VT/I56hU5LM6c8YmADZGPDlJaFR+fP5e4d+YHRnEOZ6o3Fa1OzFxSR3M
WZ6JeBqJ1zYOD5FuEimg7DsghJZ4AwgY2b9NaWqcX43wbKRo6N2qN8gtt8hNHrOP
rdFVMd+oSPbRgl8sWT/SoVUhhwofL0DoXPHJ0z0cPGncs9/ME11ENXhHHSnyDUIl
kLTKlH6KFOHjcvUyi2gMXwCli8NwC3rsU84e/bwUwdKS2SsIwdmhAWoHOwiHoJqh
4cYY1Granh6SSOmbQk5mtjGpxp82gxF3wj12f1BDxURgOu3DJRRf8kHjKEewZCjb
lZFAUggaLFwJhOz3WUpI7kwkGJfKGrIBUiR+/5YAbzPJ34eBfNwtwCZbbni6WzIg
cOS3UyHCMJMbsLt7ZAG0CbX3SeYlakULa0drVOeZwBoVw3e4Fu+oDulF+ly561rH
lbhoudTAm9wZ5Z95UoANl6ErAYUpVGI01IBv7NCZKEC29yD33woI2ZVjtkYkvmsx
1mIRYGNJRu2WwYDvsUh/q3BUMdmRyezpkHNghMcEqp63tCHy5GAgFzKQrk0C2Ru/
KPmeLxHEvoSmA/qT6bF6OoNqwfJ0y0nMNwj/MpCSBqMEqIT74qWpgJNGFz3ROF42
TfTKKeF6/6mSEx54+HmZVX2Hxp3rt/xnzScy3D9kBNkqe7VRmMGg5QInlSNGXInH
z8OYMqBWcrHhjiMjouc22dzoMJozNTLNJx9U2ntllzL9DWBDvOTT3JvoK32G7Z2A
xHDI0RYLgA1XPvzVTQ9PODsydRuQfltIHtbTtz3dh6oTU5QXjRK2Ng0vy2dX24jW
Yc70mO0Qx+U6Om0lYtKRJQLyvBqDTd7gOSIo170+jHy3DfkGwcVQsDxnmcx8v6Ra
P7OTZ6Yezjr5+aWh8Jwo39HBId959kxc9t0hrK0WLFtmRNApaVhp8u84FORgT6Mq
oNa5DoMDPYWUzSreNpw22YClUurvkae01/Ct0O6CqL3z3T2WebteXr3XnZrtCijh
8B2VoIqeJm9PVACwFym0T6jkgIxQdnB1a9uj3VOvAkOU9BUGkIdjWfPo1SyUqaXF
SNIgCDeaW3742EuAcKzXMvaf4K8PPCornf50siu+FXz+zZ1osZrMf7gckBhzjSEA
sqxV8SQOvMWfWQXsAsRyG0y48QuN/Ltm+RSVdp5AreRFoIWeZRkqduTR0eEn6Q8Z
SDCfYLLz1BOD5biaJlNM3O9QF1kCBjnS37dB65kwEYAsuLVuTmS6F5hqISy/3QFb
APDL513Clcbwyv7pENlBNe9wTBFfr+crVhq68CPApaapxPYinLlfgy/ts4GTDOPv
GBEXT7WX16yJf+jVHSh7qJ4TJ40o5jrSl+oJT6wlKwOIfk7vPvmkRuPHVAs94NGy
H4MbrFfvXAjaQVhPnMHwdJZXn9UQ0BdLegkaYddBhuHAEHlp9vA0iHoFiH2xab63
TsM+681LYt/w+fjVYOjl2M8pz5FhRv7GFutKpLzLWWPbT6Wq4uE7zg4uCo0G21e7
3GKV4nfJMzHn/e+WIUgzhFPZi+JYtUKCHdR6bkCXPzq4rgmC9Qt2AZRYEbBZOX+9
GHnHAmSOXTilTwW5PowZ3w1VPeJ0X9T7YVo5PxQ00hkHgCpAV8Fbt5FbFyvBrli5
4DQJWFeUxp/6yLGtO/nE8kK6r8qf/4DAtJKY7rQ4d7W8CsRyxIQUkM7qinR4c6cC
u1oByNQrCt+f9peCl631dBHAy5sHFHCj9WZThxRELbIWiqVAcLmT5XfjPgP2PfJI
BeADGIB7wGETdcTtR3qDfq7ZYMcNLTehmxilEqQOZOIT/F5NYF3wyeuK0b8LyGw1
rX/vzF5JEoNR2lJovovHcsU+M3wf7VKN5UXddWDvb4Rs7HAMpvmGe3kPhz6jjprH
NsDzgMpN18N3m8QOzImCibz+Z3xY5sxsnApCeQODNM0w6mcsj1V1bH3ppe1PyaEP
BdrNNJZXNJTmIt8jMn0GVAuqKv7hhgj1rJ7VHHnkVTqymkxSc/JkuFUL92SC66/P
z5ZNZaxEaVNpfhAmT5j/rSJbkorN4XWnGF4PoszwAj0ZNqX1dTMTpD4iEmR+e/EE
k3YLtt1xdf89uMAoMVN849SaQ8+Aw02/0Jmdb0bT2Vaz8r36z6/u6t7aku69K5B4
w3I5skFrycXzvwC061orPXxX/wpdFTKsVH2+sF+zoJWJD6hL42SSD+2g2iiSxe1r
6803KxExrGnGcW8KOUM5pS6zjOGDRevdVIFyveKQ3V2f2gtwJ815GB2OKCZSLwac
WX/0eUd1cUBnBS3n9z7jW7zCpYK8RsTfk18R8YQkMXQzU1SkVW3Ls+CVLOnCMulO
IyJ8wchy+7opZiU01ITBwa141B/5JFPeCiVl9jLhfTSjIrPBbRPkAqRJShYOKyjH
x83piPjdpVDsSOKXRIXer9yhMBM2ZzgXiNR7Ol9Ep3EXZvbQOsFzZOHk8xvwQp3U
9Nhl/9abjCP+uMk7VR/qoyC2CcEI3IyLoYh4+EfgB8Nab3e30Vuj25rWiRyXF6/5
7Av93itlOxBXOoFZ552fV0r3JLWoh/zS2EO0pv09Du6tv7JQ+JPCx1OujJCgqdut
nHyDjfly9OKe/tMbt7JUDajw0srJeZ1Gp+vqQdp31duvTPVbTttB3gwhWBACkaW+
s+LffyqAyVKmpEwg+IkM+IRHc78icMnRHx9OGA8XaVBULbzd3z4R/Z6omH+YQJFZ
04IJjrIKDJmiBMS/jD1htWpaxurFbGGUtM8+fvhtnOX+w9ijoRL0azNzkSp/WAck
AR7i91oefULlkQjcxdRqDvyRpP33wAHlfYPuErYd1txsiWfpgXO4A1kkI/M6gaay
qbO/EkoyYe1521oEMnJwWoDeF1Ww8JYSGLQGgnKkeSyDTUj1CIH1xuhc0nfoN1u4
dkyNzexy/ZrjP/92Xl+Y+pXtbDG5N91WuvWmnRw4dLpDhCuvSMr40gaPbcH56Smb
aqWVD+JgseYee1fWfD9OxcfCOF/zPFUcVdSkr8UXTdBmOlP3I1Ff+/I+tI0xejo7
0k5N9Bh6IYG+QLjtUtFyiIsQEDjslXT4Qgh/1yCaubl5LEoSo/SafVFVF/q22tCj
i2vgoJS5hyz8TQIdEMGVGkuF/x2NBrinyIhjNCxC8fEr08ZPOWwXzqhJVc4mwCdB
3B2iEVMx0BOUBde1vBWSK9xH3Py3QcXhI3Kutf3Xjwt27kj5dqj3xwOVpF4I/YdT
90+95Pb7/FgpvYELgm2Lg4eFXGYmkEsSXCDW6Ce7dx5xVklNqnuvhPl9JeKOiWZ/
rr8l7wAEuaaxhQot+yvc8uGhcGePjWzxP/84fNNnmG68WGM4wkrxOQxCcEMf/qhF
JsbYo0+eOB578ctWJXSXRaZSED9W9qoC9pZjPKj+LazrPiwWnXUPD8yghaJM3rFG
GaiEbKe7b9XNhMXxJjSS7tT5SF7zf81PKUOwRsKhFurbXExDMIBMCJEZQDSLyZzf
mdbylF3ERStHIkr+qOLEGnbgklc8tDCZ4Ogf7a+JJzh5gxdDmckviYUvDV6HXZL8
AWoIce3/WWYM3ranE1BzDMER1puuWwZO37oXRCBkQuRaUnWvOxv84gCsFbC0epPo
tyDWPKPML1WFmfQq8W/3bd21i1tsy+KH6Zeblp4x7I1KVx7JFLC2Cr54CG1PN/UT
Xwo5A1i9HT02SpCgMe4kjdF/hjDWQaGS9U1ykqbkVj1M7Q8F2S/nilLKPFCPRapK
MaO28LEs6PIvWkOl9c4u/tmG3kstBPt7pQzrQdVDlY4XkNQ6sR+3/m0gATe+R8yr
hUDNUNSszykfHTY88fgMCF0lLvw4y7zF0Uouh4y2OASORxN6/P8Nc1CCW//if9Ok
XE7KWEV/3wgfcaT8j+NZI79BagQNN3R5O2exo6BjrHKOQmrSvNMyMfsrZOnBoVTU
uzj4MX/Nm/fmgMUridC2OeFqUvogfiqDpeKDuxQ7rN8zzf93kS01SJ2hN22xfWXz
Q1uBJAzm+9Dv/AtWh/baA5iKbvj/RO1VPy4H3fNPI+k1oESkMd8OjGzsiTsn6lVv
8gyqAJSwIuA5qjDpqeRqDP3MkX1JDm7pioE6YIjepHtXvIaYL+O2icRTksxLxWwo
gC2Mcedf12TnNehZotUMaO/5IV05cKIvMTIvWWyO6u6qTqUukf1/6TNRcriV6D/f
jc9ceo5NwXA+oC6d0Zdsw0Mk11SP/FSYcERjrJCSlwDCbo6wetrIBKeBdlTVF4xN
+y7BzeHcMsGOiyQ98ymd/uFv6jBJv/eGSfP4Jkpe79LXbT30Md5MHYHueeWf02yh
y4tnkUrDbyGUeFOx4Uba94q++2l8nZ9imvl4eqwfT5hfVSV6urpbCVJBGElq8aHB
fYlfcaUSVDYzVmxTlzKvl6w0tAuLKUPDuL3wR3CK2znUWnjBsG9+e85ktSrN3lUw
YVEf9tOUNqYOI0G06dXtgy6yPWMnUe+XkDzQfhB4XWqtRcw21VS5C5Wx1oGeUqj4
1NoWfUEWLfnZZH356nnkhrC3gJDpAJUcycRbNNfDJJBATltueyBuMoYwpvza0wHW
1nlOcxJQfLVox/WdG3jdL5rBHEBPlY9mWvEw9jvhOBFj3Yj+mRAU9WEedfkdikv+
77k/TaNSz6pWrX2+ioqQqSlFqtn0APVv9iA7KfAYznHjoQnYkGIRQltWo4kDVF97
ImtYlqMiA1Jtl8Tkv2bnyZ2/u9+7OaAMf4FhbDWf24fBgrbGwufnE17yAFong2bV
nAh+rugWoxIGOwiHqrRcSYqDGe6mYlE7VQlHYS/EOtPaWsMV6uZa46IXVquW1y9/
Re4Uabyx7msijXjk1zDZLI6IfEaqeOt2OMZKZyjiu+MwF/uX3gpXkEtv39h7ilmv
0LONqqRWMqk8QGcBnaA/Lo25HXDrIb546bcpqCq10bxODm4eX8qzVi8XNKk1XMAn
W4mVubq4fWI7MkVNQeVhKuMGUCXfekcJ55IZwZypZ7pkCly0hM01YwSAYQLR0On4
uvoPdDpd+CpXG5junXj8X7qZuLneTmfCsOxXBaAjXh4w34Q601JrrwnV2tDl4UvY
yn+pDaHCWHJsnprQbmSuU7P2eIijcv8PvImdSUYb/VcfDnuUGnvJYND3S0bz49sK
Fa3GqZi8POpIBHj90D1MTb0A2x+uLrGASICds5dwkEsSbyeJDLDHGyI2BA3epcjU
USO9ugU+VRKplDl9AaBQ3MmEjYe036LPhdYAdajV1XENuGxibn5CpfGziv2Cb8m6
R5hmY6aDlGzWUQdTkC+YzgQKeAM9/NK0Hnr0bIfq6sphm2cUCRRTT21D/f1hhNns
rybxR7Z4d7V6RFB+EoYxFa6pc5dLSZDwUL4yLHodalWZEOg/HvA0vNW4qX633TAl
H7sJYM85g0l0RhlGtNfZznuxoEycpJ+UdNWJyojAg++SdhkSmWW+iz06UntWG6VC
lrS3NuqfRfi+i27FTNgSBk9Kmawznll0RglHs3ALPYHpYaub9lvmsN5fvdn/uMdH
sj5S73wC63ukV01CcB87Kve2igYwHvL3GqbUHO78m6nNAIRqiDP6BRB/LCWJ7MP5
+8f1Qws3Y+SCfaS2J6ocy1R6cAakOc3iXUw1ScnJOcZKqvLuaR1aQotdi5WznXki
/fs2Lg+r6lkxTx4gub6J38geSHyAZ4M9GBbof+DWUv76WcmB6tFmBhZW4LqATWdW
ZEdARZ66WjrKuEc0SagnhPGMHxTow06EUx1jho3+D1n/S2Lm7jH3Rfa6E8X2xsvc
YHk69B8f2d8M04aNjcV5Umxdmr+zAskUP1Pn8zSm2JQCEQte4MQlxMkIuREo6Mcx
ZkDtqxYzxkx/YYqpBJN16o9jWwaUaordhWUudmhm5/RWM21IEiGe8DzbJ8eCVXSG
m0wquGHKSFLYMnJSEk/VpWx482HHSOwbDithi6dVJAYjoSWP+V9UpNU3ynlb2rtc
pppSn00d+qoNp9s+N+R12w5ntyvkb126+kK2LqZ34mE7JkCMWlknQmlQ0J7PfRza
opX5XZ8yF1I1XRfqzt7qBHa45ymUf/D/CkiP2LSpYdHiV1vwnyOqouqPLjXQixdp
OEs0pVa+PZZ/qw4inEW5iqtERM3VEKeHsX7qExtqUyXlIP+OY65S5qKSYwYq0gEo
vLbnh0R0UF+NyCHYSaUK1DsqW+2jaJOm7x8Qqsqu3zjU8i23Bup/lXJfaJH/yNgB
gxHr55OrdCtM+awOLNdPGl9B7E9o9eRltgRwO2Hafmq3+p/2DbtojHM0Kez31iV4
QbFeFoF6T9TM+6OyfTXON8Hkz3NB0c+0NC+BG8OsQw0s8TBx3v3vIULAteFW/a5z
uCyncaR/HSPMPughFm2qZomy7bKqRxY+/mn34UxekDJfEatauKHIhtyfKcQ4haYl
9uJqrixXqbO878XOdj92dDCzjHskECHu31Bg2neKGaEn6tFENzm2h8eLQDe9sL/X
HVzoPx2K1Vo8TQ9y2oLWdN84nOQzWwYOh5Qgii63gwKO9JI2Kh4jDA+5tiRc5xJj
KYeToRJJ/WmoueWI1tnaUFwVF6FvNSHMH2BaR+eaRIBDTJGpKQSChg66XAyMjlbd
2f4LIA5FoE45x5ASWesEvQN5mVL80oYX4bzM6+Iu6hNWIZ5HTGWFTnPvPY2br8Pd
TH5txHfuo9HytxWYg9RUxBminpmRQEEAvfPxlJjouaat5Yn5kHqGXxiA3VrEsafD
7wUXiX22eun7y+JKyCjLnK1OWJJz/2pHutQvWpYPEU13M0hOPCVq55aCkUeTYb8Z
+OUzP/TSuRz4jMRNVZ5MYUGn3z/ZmOjcfNxtmFCqcqGtSdpnemCdSI+ttcMdCnfz
t91APCHlUghP61Uzm51x0KG3di+Ji6IeGZ8JJMTNYwYCvS2F4T8hVfQDdure0QuY
BNvpvTE4riJL9nGTigi8BapacnzyHWP1aLGb6BtIxWuVeMnkenkwhTlYBdFtPM+u
xeNt/lVgr2blXjSNoW1kMw3H2N19ZgLLCGN0+WbtyNErWEDUdhcokbEi3JWWHoJu
ujtauo8Uy5br4rWt7QE4PbYTdQfbkIIP1KcbxBPMUAa0z2LVDE6bk2KEng4GTJtj
oK2dSCF1ZqzoWXN60PTdQOStDC28kdqwURxpkCXUfVgOiW5I8rbP4u+BswB+wdz6
SfL9ka0if/QM8LlckpbacK6J/5Bq11TUNvP7/mjldMgVI8FvKseJOBmxjzhsliaC
JQ6+m8XBofuUDzMndDxsRGAqvH6bH3yYZeBO6SPi3iK0gGbe5qXl4X/oZKIWEhdh
XebxgXo4a7GL+RqsqRnE88BFotQMlM2gIcksbb66YhXgllKkO8hshrLxACENDcqJ
o3lOABtpUXd9feR9a5vaOJQgO+UtbCe+VEeyt5wNNJZMu0yv8Uo/KU0AsEBbq2Ek
YTJCur1ZxRS5cGoAyx5MXW7kDxe0SjBOz6KeHGSdX8GSTVsUP41yO121dKIVDBLw
lCwxNE4In/i9efScWKjIQhvUM+BvjHhRt4UJ8dJhHYJ0vw4q1KTJlRcF+9QygODY
Ng+FaVKhFh6GwykLmMxVUZdcafIZfSrmQeAkwTLks0eluukQNbC9u3CJBC5/qHF9
JFPQKUNW3jUx37UMXJcn/uHZkn1oz86xN3BOoRkAuTXyTsmDS3OGgMndwoaQF2Lj
8FbnUAGArbdg0eg1vXNaFa3aYog+dohgLOFGtBkEFmr5O20SWvrXseTL3uvwWleH
Ioj718mM6DcPetBucy1NxCFjXjY31yeKNpOQmfuA3joDeOV5ZG+PUjPMDHrOTkQe
fGX4nq94UMcpOvowTGTwHwcyqhuOP3FpNdG7J+9AoeBx4kji8HIelrzOKANV2VwE
KnvtPpRFqj56poB4DjsmxNmrPiDZ97bhwDYd5QT0ChWXoNF9d5qEduB0QugBWXHG
ZRd5Jzie+HHI432zmzlZPtzuV7aUq+P3ZBEpY/3i7vxGCo88ZhTqDGlQwE/bJSQV
JaD7+W0zrQWQpR1jtvg0jrbaSJp8izcWdk4iL1BTpca62p3KFm7hk0D9r9ktaDd4
yP8HOteFJ7AAbPf7drrKa69rr4P1E3imDlhLyYvRf5VUL0wrd0cD1y3FAlCSrzSa
YifLvKesR+c+EDKtqZW2m5GOXRlpKIKlZBjtO9H0EtiMiCY0jWdWx8FZzpEyG/nd
Os857UPs8XX+2BP2eHGG4jMRI+Kv8ol5LS+sGCkjhkTIkZTJLqKKhE/Wz3z7F2rc
+lhY3463kf5E9MWm8TcRDW35QaGSzx/8OX5qvleWbkwlzI6LRvAxHd8Xffjs9paU
kAQpo6rqiF+x78JbzQlMpmgbTeyNmuSnrSm5RiGTn54d+3RXJojd2H8l8wM3orPM
R041YAmEsv2t6GRkX+2ihXj7Y8igN8L2ZwEbXDE08gBcPTcKg7IxdNU72Cdtv5us
hxVJsJuJo6IeKHaYJsAZUvNUXje4rENIJ9l12/TaahKuY79Uau0F0hYvFUWSB0LD
iORQnh7u1i9SYVmn5GZbMzNfD3ANSUntWgICHkY1tDB1MA8DdseCxjUD+c/DCuVl
p0TeYFIw7A9NzZdx2Ebf46CzJsB2COBCfqhTOu3QhGfVEO4yKELfDA1fkYzNQD1k
J8pxcx9bSYFTNJRlo0CA4dWroEx2K+Wetv55yEY5cwv8e5vBtaW+nVyflLnnggcX
zKt7kDRUnvSsFrBHaqfXUD29SGHjenyDNRqM/7Q2aq1A1OBNdZxMrOiQl9MZ5vmC
CwvG4qiu6arWP0Rr1CvYTEphj1GonWmVIPNdYwJzbcKys7b6pK0gmuBdxbWA1JEU
UHlDnrhjGFP4fzjpcFvaXh7MoCmpPV57pX9rNvgahaW7VrfzDyaW163pTg0bPY/l
xLE1ctiqRZ13V8Ax+24HL9m1f0ZkGZgPDtWlKiwML15Wn9QtN23DUtSoAFCp6LOU
DLF4HjC2Scc13l5iLkmMwQHbrIqH9zm8pfehGWjQL/Rn9RWtE6ewR3jFAIuhwCYq
yCyfDmbahSndky2dvA4Fbc60X4qfJhtEF8JH2LqAntQXc2gkLqoHQ45c/DCRVvah
H+yCyfZZfb1bCEn4rWURlYqaZgNaiMPukTP3rzs6EUk1GtRXjsv62Nc+3SZ2EqZG
vXx/BoSst1xNDNBnjxjH9XLTOQAZrSPdCEtE/c12cufs5lylz+u++Q7TLf8GYC2r
X3/R1lsfnhOt9qckWXGUe04W9ryxKtITMerEZRbYx30swLNgQ4ue7GWO8GGulRXN
8RumfJYSdAbi5tQ+ZqI+OoYbtLLkqT4DdCOxWn01WDJ7bW3R0paxOE7kLC5OWB/s
OFr/Yows4powm5rnXwWyUgjHk30tNgE6rhKETcTM2mup9YheUPONQwoFkcYM2pop
YgDWcekJJwKfVEerTieUsPA1XP2MNQn76a+/jcD2zn2KLCZGYRTtjw2urbyC+VJI
RWQUyU2RFOCA462iqfQODbG1XcOz8Bxk8yzfQC+d/rBVXgy7psm2sBfHFBXq6pgZ
pzn+Of0bD4Lo/kO/GjLptBnb4UrCLdMKBmM9nI3SdToDykcCj614ZeM5k7Kb4xH2
+UeuA9hYNqss8QDsOhOj45U+qKkREJ5gCXFpMOAKEFoGvZlgHWi5HuZwkppFKnve
lQs3CIYQcSAJphJ4TMATpLHbmb+lRIo600XrinhHyc+2Lj/+lavsDIWw2JP/4Smg
WaaiMe1Q/QMwRMTqOG2VxdGHP20kDY2n92nxnqyXDh4V53r/57qD16UpipfJSwEq
vgYCM2L96j+TBeXKiZj/B/dmn7UMZZ0xwaIdiKAn8iw/TQQCFBUDtuLjmoYabSp8
JR69D5uGOv0bfjqCGkoCQG05QOsoBNmeIHUg0VyLAM9MHn+KXiwAXNPi4mz4nBB2
/BUNfKqSnRgcNEmlvUcDNcUjBYmplg9w2sgxgrC1O7yHg6pvBNl2E6EFM1ibk/lN
Gy3tX98GD/JGqXi0y2VRzBG3O+BfnDVhYPAleycCa+q2SzkpUUJV/i+vZThBhcwm
n55YKBYgYsWPcwzME11IAUeY+N1M9WFokXYGzePBJHxqwF1tK/mU+VJa7btHVzRs
hYEVSPzrkwI7D/TNmdztzhHk7PsaO+mTpo3pwWvaM7gp7GevPAFZGzOQPnb6mOJs
zUDdvba+/eo+zI6kRJFIuj4DJfd9/XRRlsO/LylPA1YbI4jVldxCsJBiGX5tKyPQ
XfFF6dN2smt2eUVFuKgSU9kRzpZcGbzNxPdiZ3jCq4fAKJbsr8C1x2AeJQPsnSfX
PLY4r/aTJ2INRhJNInMzeYb429ZFg+KnePN1YSc4EhWEKe4Kun8RyAsf5GNnYMZR
hA52OpOEE4IYqwtDGXSHkHCR6dzeHHp5YkqWLUYCZdOWqXR1xmxJfxCLBS/VEUKK
TXnVFo6NGaIGi22Y+XjoF+HVtV0NH4KvbAzc5aZ3Xu/iTOzBubtufdxY5xBY/1pW
MPYOOJ+Iia7Y6uMr0mkdILk5r3Ep4XqI6pRBjaPP22tvT+ebB+F/2Ug+luTu1Yj0
FcjcGg9uxZgqhmBjfLk0GmpR7fxyTI6ESVeXDVM9QJue9TGZDKZ7zmYEnPww1T1Y
c3XZ8lH7PQ79CaIHqxD0WwSM8ewqAzgKT7g0jsTxkf79vKo7vEU80v0g15s+B+Xs
2KCvNgJBfR8nLDnxRrcsjiKZJjAK1HrgOc8ljFGMi4USFcNixPvJ3zQiXcwjZPXq
azN6JvWmfLbP6n05arp9W+3yEzI36/1A5MnxEnte5RLS4gFa08ky8jP37+QBeGvj
oBHzX8KhtwP5LzxrWckZy23xuKK4CiYw+8gIpqr6CFkWoaXjy4ylIeI0UHbrO2nL
oPLifLD8K/v5o4acsENj0D/dQvl4CDY/wD5x6wM93IzU0oAsE5LLN8ufgxFPv+jQ
xHjdqxHc/C+Z6QPDgbHMifZcfIiHdTjkHMAie7d6M7nyAlJoe2uFK3/Jx7sfJJRz
Ibr7RyfF71xL3hMEhgw2E+qyUMZsEEBhyPsw37y0z1u0vbkP1J/fwG/qEdN7fv+Q
OLM8JRHulVea2QAz4JOcB1BoLH7ehuaMZ+RmR4qEa8i9tu9yiMe1jimjd/3qBea0
FAaHQfgbCizxNtzv542JkdezpXq9A1J3ctTgUBWUl21AwIv8epTK0CBu2MMSZUML
7KF0J1DD2fO8Dlpf8uTB2Z4X+LqyKOKYsnB1YqkFy91kY8uU/S6N0j4r98D/dD2I
k17EqcMzpQh/2RdQLh3oD4r5o+Wb0Y4WyDNIypdfPY5mN597xvHArmU1ZN8WbV6F
QXoKKUHJrTKfpNTZ6MjsOuXL87DMIVFbPIs8esvmBgbXt7If+v0i3SjDWI5agMtn
TB5ScrYWNi1LMYA4tC9xYhw+dp2PeqrrT61wbnAkNAYkO4FP1TqXenEHkngZG4wy
55/pGpRiuR5TBF4tzHPzzTOTAtE08NlrBTiSMeANKxultNSeULcVTL6KziURZDuj
vR9pSn4w76Iud4izCJiXCYNY0t5jIrFaTlChoFa9W10KRV0RE22xR15dfnpdrKx6
mPr7cbDU4318kiIiLsx8SsiWE9BpZqdZm3+ktZSd9M20MkLqC3T8fHucECZ+Hg/J
L6EOt3nFzqWssujAcnr+OongUHKffyCLaVFHhXl41Z+2qqXGCVPEp+w00QF7T+i0
OnlTJihAcDgUXNcGqZTguZ9M4CnlDLn53atNKt/ViHCGbRcz9Rwoj3HyPeKm1zdv
CEJZORaduiMOfuvGLsPDx2wQiX5saBDjjwEwNQW20yoMpaY7eJmuEJqp5f1lxTtO
EVY6VCIH5Up0KjRA8Cx3M0XpEH4A6ykvAJ+34+6NJmcUqWT5D2AwygBHxl5bplx1
Ah+0kzfgzGvMmfkPBD6JNHER3WW8A5rkGa1Xx5eUVWkGEzup6R/PnjNyEFQNS/r5
o1e6ZqLvdFJ/PImOV3+PvldMCV9iuj3nO8iwD5kMuXTozjr/AuKObKxI+dJa+8OE
dkuPRW8NjonL7dNQCvsTTM9Cg/NYwAjFIE5NzuM4jQDwCI0kOKibGIBQa2TBYD37
hGI/3Xu/Fb7bpi9Ej6BRLTIyAXryzcLzGPXHfgjwfVTvEkK8yHAbJ1QP9TyqqZpl
o0Wu6CbQsYAmDoxtWRlHkyava2iF8r/hueWl6OYfCQVP+m0zkvM//n01kU55VPvL
h2Gt22ax1bfVuiaGsvU2wozJEeAWnRNNo7tQvLCN80DZQcDqz/HhG1Gd60DZV49E
Q2T7Pz88vlgmOmIJX+UCGASRV62V+ndfgRfkwe+iYhF0GhvINBAOEJTer1X4AuOy
XvWoWHqLQ1McLx9nCIz/W23L7Xo6G3a+LeA/KbbaIsC/PxNCqc9i14xS/4O87vSO
CINryfOPPm60nwgpmVn9X6VzA7bDY1yAm4aBvfhYXj0wLgkNFf8dQeJn7RyQouy9
zLYFbhnAcIItpVPPRBQTV2w49dKl/Ab2NtVvAKxBbP2QE7l5PS+N6eeEBxvDNGwM
OfB4HMvC0J9/ub56F7VsV74imvVfchpFFck+038W3NAers2Slk7sidPPUfCJKsaZ
RO+YMe5JYoP5YY6WibQV8dluaUYI4N3kJ0LvWdF/NrB5Goc+H0rHoy1oHGaSG3Ki
g2AyzboBWToYUYuyA3yvJmqTYVpZmG2jrn8tp9GgvM8DZkW/Mb6a7GfET8fAgl5g
kCw4Ay4ZUMIB6ZpIeNCaL7p38G0B8nQba7k6a8Kh3rwkYUwGS5Gqr+XD7vdmZxXD
7ruyTzVBNSHVQgfB8ePldb6VQUi1wjdpjzbZRCxD3rT2rMZOVwK42OKJiVJIDxop
Pu4GfSzDQ0x+lCsJfbF3KmsHHNiEhzOlLnBT7wPlsjF8owLxiP3kNc0kD0ylMLML
JbdxisxnYzXPpbD2Ojrsqs/MPnfd+2noGbQ2RKd65UiJvZXCHIWgwqC1vzhELYiL
P/apg6bx6dp9HJmAYXNAQ6urFHgIWRF8mc/hMKnxM+pPc3VHfQRNZJJg7EiDvz2B
AhqAtHdEh1E/Wg1MwiJA+Wi57cubyoAtdLahuGW5WSPfhbGQFcX9LHyOCdNf88OP
xsEmOhJ/pE9Nz9jx4aBARVVaAc3pVMEgYm3POq7XU7rwx+xC33aWGHcdnn3EFi5e
4zViR7rspPYMDvo/7mJmaF/IzCTKoIWzfYMgBDTHvGJxVIbRs+++EWwRhItkEzu/
vSo775QPU+zSwaZvoduyI5zy5iy1HSCXSN10fn9m7GkWie2zgjtYFpvFdDC9wdgl
6Y5G45fPWyAUnHYUYjwG8f2r+1dGypXRuj2rq2GgueTWHki6e9+5adan5Xu9J7Jb
1J9m8cYUb4oxuToD+k9CthhEZ13W9DdQmUn/zwnUeDdqZqSU4nIpKQjyLZgkChZF
UhLwhVFUy9u0rKuBDX4sbhDhrDqnmo2PaIhzOx/UCQ7o9L5GYWNTS/Gutou9JH7H
WglXdzRZ7FFNj5xz3xhzfdTazv+lHCYi5Cqi6NjtbIgF/RWR9rLIQ/A9Sil9Pyfp
8qtte20arycsxp/PdV7epkFyBfvpDGqfcy5EGTqLFATfsSsJckG9WFqL/d46KCvI
NC5itVvTOK8U3I5Xkee02+d/KeFX1VqZrdA3LeLLL9qvGOLOKj9fjVphScKNjqxh
tTBt8y38CfVWUt9hRlWi+YT/HbsVGxqwMFnXtyarR2f+S66ai7831q85JipEh2Wo
DaWi7SjAlOEnSLK82CLyIlYJY2qch3BM70m27YpRBJKNtCDZZaUF6h2AAzCezxOJ
4p19/g9uTY8a92Uk0W7ALLXvNsxSs1O9x9CSSGOohFVK8vjDrWOZClLM2EAtoGwy
jIUf5c8slPDi/f7X6MAMx6Ll7CrfrkLPbrY6yNFYLUVHhi4vwBxi+a8X6FX7WKcY
nGNBM0vOP39BEhJGQSBRjazadoRIdLwa975TgOw4rCnpJk7+3dm5Na/e/frD1yH2
l1TJsZbb0f6Vvaik/w5+fwQFsrvLYjLT+CRdunX6W0a4Wj4Wv8/zAI8TjhIfbg/A
OqEeRP3kP/djKRcV4jp/zwYPUwVLolZPYVzotVDugX9nvVBldc3lB5WTRIygHtFJ
gKaw3gtQc9N0fT2aEk7Q3YtJ7mCVA+fLfIOwei5L1xTAuRAmF7PRzBBJthSPqTi2
uD9aW/UcgcdnXpxBzd0OpAvg5lcFhvHSkbWXCACQMfRV0EThuSZKhKlfKhozPeau
7C3rjYA/OwG2VvPmF7GWxBzPcz9u4L8486wl98m5g0X9EElz8myQnZVrac9u4fES
Qos9PhPPghM4kdKWN7keZeNLB9I8k1idGg92iQdeWZtU0Q0f9XqNFGBoEyqzK6wo
eOvbei2EmEzvP6g14bRr4iC8I7l5zlXGpS+IfqdHNjJ+n3RZMh9Vtu9ftDPMczKX
nZSH5KU4HMWrj/vmQvAjAf4y0B5RVAEJfBeJ64mNHraJb6n6JjvDHVTOMk/BuEiG
WjfXe95VNDJyG0EgZqBv2KS0ANGyZNFybUndmTTb3t5KTP8FBHieiVwBmLuioUq7
2tCRsQl5tXKaHXyyz5EaLQDpwuDtiqGhp+dVON1N/j0P/TKGSCNl0RoDONjiWxaz
nFewgOJVEGJyAwfc5HMNipMf21ICCZr/SNzxgCbO8kLKA0aEt54JVdEB5MyujgZ/
DAdPzIi2VrsVvuna24cKmpA7Z+72V+lWLhys3E4576JbcZMdwX/Wf8m+DsWiR37m
DBe0OO85jX8YQg/k8uKgJJtAsNmKI+sLOIoEhyOUCNz8Mk+S+PhwUXA/6GT8CEbt
gnsWQD+P4eVCf+J359iemDX7Sag4kuzakHl+GmhbEGTCwUJwFfF0xoiENZplaF9i
P+lNVDVzK+e+0394QINT5miPYqrRnDo3zE4J6AD4qE/f0mDzdP2V4eZ9+XRQOCw2
h3K2YmxwEkpNhNM6OS/O+Tyf4uRjINst460SggWyuhXUgWNFBfLv+a/lwlEsqhKb
MYj03mqUwGS7GMuHJHRtQD+m8aIWo0lORwEajklOsjhm6YsvAXlf2FwJS4n9Wets
3mgFTM44CsE3TPepvrMjU7vksCGcDlNJUzRUbIhQa8tkptRCK4rhyiI5xlniJMTr
gLaWPb8poqs3xj2I+XysFzZDJ9rjytkvVrEBf34zmp/7cg1bvAs9qlzFvWlX5xfT
GoNay4ws1qWiQG/idgXFU99ilIysIEhsEhT4wuGYbbqvDx8M9jSiIS6U/ZCrBuKm
p9Ymqn5ZjBOMzYqqPm/vweKaWJAn271AhFe3xEEe4T8qDbrl7X+HduPD3kr4NK/h
uvKUXbJ5iWyFp3udL67jmKVV8R/MjxDeXTzWErAT3PsB6gDrvzdhgeVLVN+n0EBj
NlbVNn9t0+F85nXDxggC0S9J3FD9HWNuck1XVALvgUwLZCnnxTHjlONWH7Vl/xqh
il1YZHQjCx+UixlDJeAETL7n7Iad+xONEAKvBv0J4e36sbQZmnjzUEZ13IJhbQjP
3h+7nr+FCQNy56dfgT+yBjm1i2h2Pg0MP8Gbg742Zj0zxaKm3bAddnABWf6ubzaz
hr91hc+1iSJijnTD2Djdgu+04K03+pXdRYLo8z844Ab/pWbiG56Lz1Z7ICET6A+Z
2av9nX2u3sAv4r7YilDsuR6/oHGzNynEr/4VI5PysCme9BDVM96eTPib+Gntpfe6
uO9yTYWjOMB2lWb4ghwSMw0/b/jILvQBDv2ek/J1jPIUjoy3/mP+726XqpMlipS2
R4+auhtCLf0H0XlbGawHFcL6i3NLYtYCZh7sCbLxg/GwWKWR3oDVA12ZFKuOpYjT
moHM/f/zbYA2D0P1t4Sz5l6Ysk0PONBp1FqwlZG69pmNGA18J2CHXDoSEuPCpSiw
X1nkooiGN2TMj7UElEa1U75u2+y1oiqhG97czQIIOzcrrjNjYpkp9A4ihnyaDi5U
sJg39MeH6TIWgTNjmjEHwJCxNTErCHF3lDbS2Y8jkeFdJiD+5nrdlv0PUd9zWE9C
IropOJvu5SP2tXfqBksUnPuHIL9pm9JolDZA1LfIXtqG6D3bzoPCsAebPFS4vwNa
nNGlh77NrZJsz9dpZrjPVvegrwON+EergezPbCET0yv3nwFojtR3p1dAXfi/G9kT
xqtHOWvvhvAPKZ6QkhGEglVhPjuSgd8FegcCap24qlUGqtaNJMN5etd/NwPeARmU
tOaWD4eZ3o3SDnu+TemmSQy/d4S8HCvtjkkBP/x/uJDcilVvXGplAgt5RejyR0rJ
W8V3Q8MykLeYmnwFm2vU7E24LhjYNm4Y8bYDVioRVi2P/fH0gjTWH759CxiviEAO
u3Nm/xQ4838D8dndfKtelfBEQoDoeQtjP3y/3CxGGPAy0scLJ4hyLzSfdcLpzF6i
9mGX1khD0xXVZo+5y5hVfMc1N1UhUeMtREGwmMg1rqVlZ8HzmhhJF8JT3OgFWlS2
AcwATqdy2rVyKDWSk8lHQdZFaqDF9GsaOWVkiTe0ns4wlaW9xX5Od8xN9DM5OlWe
JjwluUV2V5IzDguNW+XukAHVpo2KnCYe4NwY63/sFePHILBAEgAnmHMoyTc0GzVi
rNRd9eOxVCOXB/ie7MjK3uZ9dbZSsDXV37LkQ3ebjOyvpkkonRUzcApntz2O6rOL
Yle5Ykf/Qy5ipSbNBd34JFYtGzOWVCE3AO2EC28VTyGxTbucT4RjQoELoDeeSQLA
tIFwEBrd0z/pSbXR2X63PCSR8+7kG4PX+oBpwC/7u3Cxeq0ElRgHu3a4eGUMQymT
tJM7+zBvay/OvCNWFnzyzjfMhvwly7aVjgUKKzeR5ZA0sHbZK65d7YUYLh/DJeyW
g5rBVwRvVKLzQoifGajVJk50AB8/9lX+37Df5PSI9/ZNk4LK9YGleu9/WXLrsdhj
PnR/+Q/K7FMTqmU+fn/LVOFGD6nGzQOVJ976jTF1zkmr+WfDkJxzjzMlvi4ZNNRB
c6dNaVQEpLJwF2MXNa1uIAWxzxmvxjX6eqEKrUePrV0W/vMjnxhkfeq5VNET4KlC
FjCfZK5VbCk0XomToQb0kKbOMsr67hsWCJfTrE9G6h/hGrX6p70SScpJ7fbP3HSO
jdl7jRL7v8aUfHcoGa15NfBUYBPs7Gr90JQlj58dLwuBQ/q9VoBFY/jT+GvuBnmX
AOmihOdv/u2pNAqr1YNOyArTPm7OJACsaaEGlRXoBrANi5OijSGBPdpi2kk15Puc
gGNgvZkFSDRMG49tKCsQ+v/ZkjQXikR1nAaXlpJ3VTl2P68TgYcIsf5E2ribEfNo
GXSFreK5RksrMGFqMcXLJASjCTyPc6rDYTON2heXiYjbmQV85nPMMzk1C6CTWd9y
ySE0Y3Q2KVxE3n32GywM505wkxfr8pZf3fhBp3pgo0mUTgDPdShQw276R0ldyUfD
TGBTr9CzrghxW4SIykAy5JInijNuwvbxWE/mrkZtSre29g6VL1u3+K7RJe/HYS6V
MPVMMibF9SDWx2lj1xuZavr8uNbXmdJ2zYMwZngOyA5qjA4Z/eP6u+772Rn6NKep
imqMlfceQYxxMnxMsJSVoVXuwQhuKvwYgsjh8fsj+1Egho3XJm6blGus7Aj9EDfl
0x7bqnyb7mpgDaSCdy3Zi/cZXVDY0Zjq1/JraZ2onnIIX5OqVcP0Q0Qr/ROKBM84
bGngXIUFMZe9F/9CmxqC3MITe3at0jvuFo0ZoYX9yZIuWrdGNVB00n1zIpuBw13s
NgGDUHgWJRypLTJ32ACBMqjjW3UieIeh0TlDNNcIw9klqa1eTpHRTMDP+0iTfwPO
DYrxftU56/VHw/WX6+6IF5P1G6CyNOP4lkISlc039eooMCSPmOTCbq74dt2hmelq
AJOGTru0/R3KKV8s93Zcs7Kv3AOK/075KoIykrZyPViOT/iT67nxgkRjOW1OPyM8
WhaMvs4wBCf8gUPlnWo1ceyp/UovHqHA182HH8Zy48cWkdXbd/EqB6Z2jybrHZQz
fLLrQCgaKiDM3pYuVosaGYHHpg/mJCY+8GSxUsooeyMGKoldRLuC3hoABZKupG4D
iaRSB/FY9CXkgxPA3Pjzo7iEMeHPNLy/8MBSczExMMvT+gNZLmExk/0ZlwuygmIu
TDtRlIA+rVaJsdtfr/C/6or6FFc1Gicu06B6kkQw4m5HPt9R8aoF2Dkvn1hTGC4o
YKyuSEayBwsYgigMYujR4vqSZt0ZlEkdMETHeBQCcG635r5OwQ87lVTSjImWkjmJ
OTPhfmv6MNxKyynvWlAtHEooQvup4KxJWaaRxGQSxFE4h7KmMn0IQGjs7T6Eenpe
sYteiWCDYCvr+yAYJu4bVPecRieu+JnHt5B1gTMZ8dFBu3ecG+lbZ6aqHCGSHaUF
zAbNSSFAeVWiNdF34D5n/NwQvzDuwT3Yh6xk27i09uNvNhE3hrWQN7RdSamJ93/F
Ke4QQqPUZ/DN515ADaWrl+l8bji/XgwPlN2BhW5IGGFGbwUD5keFQiznXpXnRUzQ
9miQwPkHhSN0L8pS9n7QH6Yf6XBKiKPs1kOjClYPKfO71qfrKLZa5IlsRpENigq6
YEoBzwjamiKqXmnhmLIcsByq24Yqwfsq/64XOO8e/745u8URizPW75Uvq89ed+80
/CSm2lQ5QjZUxM03BvMkRtzsrKB30OREYtrrYzH1Icwy3fBMwt9nRGJ8OFl2/9/i
UlqJsceVJxjiETTxwlUaNv/DO6Qa5x9KsZCNxsvZVo19aOzJfRUnM6F5jttN6jUh
3u09NBEIlJkIA2aYENLn8ZhqFWPUvoTPe8FLnurals2O9d6HIakX0kg++alhPN/y
br8Fh4LqNXK5kPdBx5iGUESo6hPzsYP+I3mK5HRXQWtqcrZsx1T+NxjLYTEPD2nU
T9/DRsEtWSVlIVY/7DzcrbVyvoh/E9Kommktu8mOU2RB1AtVKMYDokBHL7lqu4uN
LLtvcxpaWFB2x8H8QJwXJN0FwQLBrSVjqIwtsebMzkbwWBjHSD6idY7iVbAyNrxt
p2hJiUPd9zSVLRZI8JHaJ4RZg6Tha3ha/Pu9xQ9OXfV7GqmAKJwd+mkA3BiA8fvb
IpyicVA3JLitv3ajfTKtnRwnbEJgrFKR+8XsDBdBmg1qhLWew7BqP1rQJOX4kdmy
XeRP+ZZ5ev8UU2rhQQWNyICJV+CwMUgHe0G42vfThmcSjudbOeDuffj6Ax7kiymD
4pxEGyTTQFcRNhp+0GgusINv+f2LRrZdkgR5jGpUce9fy13QbFIdgwmul2yMQ6xR
dB8zu2eQJ4A4VZ7s00Vahgr6G51g+wDEiZ1KSATtKrirdWElRizSkf8yWh/2e7zW
doHDw7FRBpK0lDlCOJI5jfYBt2Dj06vSLFP37AfO8NU9sPKb9X+6L1WVNEDOzGq8
/J3vOzIzvSV8ZCohbyIuepn1qoa5C4vK4+jaL1hQX847xNbYvkVrU2hZ3sE0BCyh
52Fr7Mr03Y5dL4k/W6P3TZXg7rs8zAUS5BSYv5Z9rgdplb4adFjvt9s3KBsSJSyQ
5nnlJGuSWX6DTXVqVOhqDVdqyFIb9kkQgPjHjOyNqQoUvKTNl+pLIZMzIosWJTuu
YalQov4rscGOBZfprkYwBlN9P4FPT52+6G384fQc7gurI3g4isMBF9NeRlvQHjyZ
Pn09RDQ3+4xRxkGWWME1xxAbi9wjhHeOFAFjwM9BpGTTN3r0HYFCy0+ejE/+5Gu2
L586Jxaoz5wssT7qSKB032lOKv05R0zKvJ7lz69ni7urjvXbBc3q21WvoGw7dLcp
d+LIDw30UwO2tYeIro18qPcpPXrY8qRrTPE8thsbJcitneuDlxLfT/icnAhlw6cg
sFhUA0WhLMJlacTPBAd+NoTXanRfEvCrQ+sXsnMdCJF+jMjKw7L2TZJ2Gf+vL401
n+S2NzyPCsTcpPmq4eAfzbBz55PaFR2PYQIUFu32p32UAb4K6oIIZk0dMdLrNkUv
zQkEmhlgzawJGdbFrzMtNGDYZbPCHCHuXu7oPcEIT1Q++YwgESiVwbXIkv9OL6E5
3/SRQ9Bm0p3aW1V8SscMOXpgrv2uDmVw9qP4SwVWlaU+ceFIeqrJYV4JfkwhQkc1
kdwH8csYDtm6Fx84+7zqSXF8YUcxKiAa/aU1v7AGUz5xlCtqmakhqy1CH6OycbKL
aYFmfbnKlWgHzjb19ZIVQR/6E1PVxyfRJVNx7OL2IS9o4317Por++4o8RSgZ4Wul
DHEkpwhP9iGeuuFrdOhFGsnOSHsszzgyAv4aYDdu4oM/EPB7mLVFAJ/elUfjDz2g
57pfRjmxxXmgLMQJaQGlZaKB5TCP6o9IGvslwMfarbheEwV+tVRnxRHMEzo8iks7
90IXk31GPiG5ahshRJaPGK4jmvRIiDwpI4z+WJOx10HfvQt38NvGptMM0SKwRKF2
jyNkKLNm6eP/lfe7+kTvM6XckvUQC5US7CeHlJV46q1/icrnYDhVDGVL6e/yoAvu
befW/hSzL4/54pqAWxhXuYCttkY+ETeZCE60jBQFbh+HsvDfd7bkqZcEL6Mw9RQp
uPn2hy1VcAgLA5XzBHOAYbINg6ZvwO4jIZgKQrQUnDB5cbAPboeXYYLLlcY9KDdL
cU8VQfS+QSQZuJoKVpg/W1QjGfD2GYPyUFJTh5Z5rwVq/tnV+ROsskMJKhK3xxiC
M0JP+AaWr2vgJ7T9DFYCkFSHHX1hlDNnFqhp5Q2S6twcH5CccxEKW1m9F+V0zDWz
vs9792KCelDvVFGz283kjUpNg5N9NntrFAZ1I7IBmHN6z5/NRKYGQ2kUOgkSmHqU
g5BsoHvQMx5vOe2Y7bJICvMLQ1IAjbq16BdsevO+WN1RcItmcA+WDIcjQuSOY8j5
HRsEdcFRkEDRM+5PflWnKXcD3hJL5gYmSQ4WDewh9grUFHs7ekKTE+dLkPuMHXuz
rPs0ZOXWMNz+p8OdtaF5DWACwdzUr7hIoL0Jr3d4x5cEW6TlQFfgPeudhhoUsZq+
lU7fKl+NYgcWYs0dZtc1t4kxKK+s3v3+iWlXMvKvsj/z4HPphDOjQwkog1dtsNIj
43CZN64Ux7xjLEhgOfQ2DQWpbmwq8aoSb3zn9z10UnEIL9ZxAQenqqMKnyyFVXWa
nrG81F6jMqSYFxDsJE5/sFQI1M07lh7KIyRqTOyWGxcYCgSy5JcK9xKXgr20XtNe
LwEzBv8+U49yBh/+0Z/KLvskgdvdxvx3ChWCYpkSO5y3AWbhKIV5fpTMO/TnwzLk
0dqo4ruBsIC+GCIIOXauNgybXoP0QwF2GxnWirUWrA1yyin+PZncfox9CudGeL9x
7PVAEAed2Jxb8UEEHdlm8bTJsYT0Gsdo2c+pdL1Rib5kuX0LGKucYUCKYRSHAWBO
hNbBXtj+hgcHWW7mp6v8CGSdaPYFkgnE7YBvqbqCHZAOnKkLdI5p6inSdrg9m0aQ
ypSTBwu2mU9lHsYVP21YhMP4wrSsz2WdjZ2GM3ymQVmTuFNhjxzMHcTy4q6anCX7
tsb6viUVeFq7zK4We4p+WKbO4cmTKlwLKYHNTCb84LRwchxRiLBtmSSoG6cvBMSB
g0OAsPq7a1oGBAnuWScSIxVufJnxN8LSQCEigI7b6TH4FeGPf6fn1g3/ylfHAkck
aXCPGfZrV8zykYGnon6ZQ51AohaMJHj67lG9pPnQm0XS90p1Xp4Bev73DrMejHz5
CG6tvaL03k84MyEiTDv3I1HaRLIFGqgOkrqd8YzBlet6w4kK5em5ItmfUMgvx6KL
PqSoKCqU4xICtLWvXkW49B7RavWCVrn/kWqhQZY3HC48y+K+UVbLIhuGdveeT2hX
JIa9S9TtwPpxiRu9ybcYdRQgRvZogFq9Pm82wtYTZSfFULTHiVO8o3U0//73MXtt
SZI4EDIF06/9qglEKW+RpWA3Cnt4i7qPWo+sTWOWyjb/Z7wNTQ7fPmuFA7yUEDro
4K0wboAarDufZKHJmZiLLOnI1x9P/nlq38hBhdWJssAUbExe99xrWYJZqnb7lBJV
Cs174oC5rRuq+IaUQI/tzdAGnHQHwwBIydUcnkQN2Y/Gy0C82sCS9OkYoqZ4gGlU
02TF0zwAvKMLCRd+9mLxuV42xEVyJ+0OR3mbEfCF8xfIvnUtQzeDjuJEWZISdYuW
3dapLmnbDr7KLeCXe1HEFp9F5HWtRADwpwbWOKhxMQETR8P8TV9ti8n4v1/95JlL
5GYlRezNs6G67rSgK32gL0m2PlqaG15CCWG9zH4dO7itbU7oe6w4wTJYY1tC1Ipo
0hRw36/pbUg8T3UN27K+8s285SjCFyP0ci3DtiW1xusGnMwcu9bC38Zza1WqOJW2
5Qg4fAm1mmlpGHo1USChz1+gJNN7JKLbYViHR+Z194GEmMG9v9o5Qi/bK8PtSO7x
Vl7Q0oVN5vZNqFns3HOwkluocKWBc/8PrGZaIYkdltExW9LKrTgawMIKtXdnPfH6
JbAsD/W64Z9LrKssTEqVnEIC4kxzDKH0PqeLHtT3Y7DAkUVIF4IPypGlPCztU4IS
GW0YG4BZzrRGB1pTX90wuNJ8JzEO1zXmErkf77UsoOioAFsmhMe19BFZ4evPsXBH
IskdSjLn6ahEitFUcU/m77m7quHK+Q+Jm0VHc5lwVuSndtT6q8xHx6XjaDp//oEa
bXIKSUUQCPOMLlTGHmtzBNTy3j9+qWyHshGX2uJKjbG+d+LAvo3DrQSBfLeBBYrD
6WCsD+HtsiYRW4ZajitgkBA8p7rD9HCSN4I19wnywvPc07HR3fMT8k49QcEidQKK
gtqv+ogEVcXwKJ4Qkg5Vr5DgKyHE6QC4PkkkAAdxjvYhnQ5QzHKa/Vmdk6sxn2De
0hO7eERlcvoCYC3Ec8IR2EKDLYu/smAIW+HgdnwGBLtp6EpxI90eeFy/rYFk6gp7
eMWjxqk0J78KvLy0tqhdLH/7JRyp/9ADDHHCxtSoKwyANs4r+YcJcO3nGUzYTcAE
ss455c3vDwPn6Tyc165GgzscBtmHdxnw+C1nS207dx28zYA2qBKpK9LGPJYaot71
bNynP5H+3sNc9lilUA3hK7S3Y9idLr8eC4Z/02nb0ZXgo2Gx7irINfkKWCGRSb01
rnXe6HS0hrJXX4JP1QMZzCMfRpkEd/9TcVwWahfioJ/Fo6GpqUX0EKM8rt9zkjCS
csOO9CWX93sbLLOsVLbSKAkCE6bCZRHYKrAny1q+pAzXksUrab5dBVj0GLPEkziY
8SLAz67l2h23FMaj7Q+WCeUKkk/K1wVoj8GvO2clV8oP5//DNmJPZUzGKbOeJYvQ
Fmiwq78N8dQNpB+euBAd9JnA4sLYS8dOhwhid7idlQn5L2odq6D2zPxcQUCefMjt
WzDLzwwMWYpOcJkl81eiCP/yz+52bSYEwR6K52KNcF55GXTFJ6yKyCNgs216/A0F
hSSXND50d6QXfl5eJ5lWzPUXzVT4TzoCOc33iMZOGshrkDyPHqY9flMsvD1dFIZu
VJ83BMD/v8nqEW+F0lLjl4lcmtsEkNBLzUh5wMzEud43YkHYIc9k4bvqwtXEfdZZ
lqpWOXvro5XCN17WAq3mOKOfTyHYVnlw5ng6hkEeyKq0sSBVoxGnFxGlhNVUA8Z9
KKwO3DqiRheAaV+HxjIvMrq0ijD1g2VpIhg6V7t8jnSRJ8rtcQtmaOUBqiIb3paF
VW2r5Njitds/Wh9+kyZgS3UleU39xxGO68SrJgnP4hvGu7bVA3XAEZBACc6NnT8N
ZxojbLKBZGk5V7MP3XTvakLwunsc167Kium8Kz1wyCY2PznoJmD7NvqBQfUnpYwL
Ph4s+/s+3fP68vyjIpyIUILLG6hcM5Q4SbxeFn+I3JYtYnFjbj2cNFOz39LJmrZp
PHCygtweKur34YBG1XFV2nqf299bxt5jy84XLU0RfnOrimw60IhExDskcUu2SMU0
UMYUHFlIWpcMOP9onWtiRU2n6LXIjTvW+kjhvx8SpbL3lMXIm9Pw2rknRvhw+zoi
P0RRCYpbN+1geGSr5suX2QW6o1JVLqMgz4flY5Qd6oDTxncyCfPjY73CQ/hOGdi4
URxAPFkMOTKaLUbAVJSyHlsaHWsw3MY59WrfvAi7JgT5d3Zt6A39HaiPk0D8e1SV
LEwEPmAvwXjR/t8iP+mFpugv56WKDeKKIoJk94nZSGqC9essaDQnsn3k/2xKHLrW
nQgydLkD3VvsZ5krhjggVb0VzxxfampCVtCHgeGMyPjpb6X93ByLxkVy/VG+zYRy
6WwY0os3c/MjG7fMx56MDpKHby9TFfYffqSR/lTUhQxdG1DR2fytj8eQqA7koxfC
GvpFcqQG8C/C7yg2VCC9MzbCY9jRh3t2l/zRXoOwkN2i4J9SnDNPxkezozN0HorL
jVQJt1FiOP3Sf+ODVttKu9uISpOFm0KwgJXegEx2H/0c1ytqYxDMqTaue10HXODv
NRMMvmNq+gn1ZsLKdtoy+mU57xHih4IGriucHOxyEnV6ZmuvGO4XcUnORLoJXOLY
/MKCg/JQXDKC+7ykC2pr32ab5KE8Mh0HdQyjd6rAgqehkYjfHWw2NrEH1JBvXRux
nPqZRLLjtI0yQOmXes5Ne1BcwWzPe7sPm0elaxegtAs0ep+OEzO35yQ6J4CHlXfr
/pOsYin3Mfp4wcZ8vlOrJAieZ8LCHicKL0PumXB1GYjTXj0k9TlOjsDf1fG/h9Yf
1ps/nF0HJEopgsWxLoEArTe8qP7mxkhEUFt1WSb6ApP3BI6Cpn8Jc5cCDXI4/pFr
25QzvIAIwpHyLu5hjYZDq82gZ7Z8d3OoCZV7I/UsdaWnJ8gUIcnQRm4Wl67QYybI
+0sthRTvexmX1rb2twLFvwZn6287E8QLfXx7S4bnpAJEzq0rrTT07qowxcoYls/H
9vs98s3yJ4xy7nUg/cr81QcR58D74Uf+s4z1f0NzTkGllUNgcy57Brq3u6UDGj7O
v3LFhS6nUvI05ngRlOurWuQj5c1lMjOowuAKUxez0u48BxhkuTNc6dgEJKCJ8JIB
aRUFSFEtAAZSzb5DDQ2sZp1sKAUZ2e4LujXEJbXjavvk70WGujlCfjuvIIncp6f9
gqeJSCRIDvnvbJ+lJuxDJcJly7XqdX6CgOdg2KLKXQJgRhgmQ85/eqeXcEecpUYo
QH56r+X63MXQGfZExs6HA4eWnBw5obcLN+TMFR+DEWQnlFtoRomYScf12m3EvOI2
rTn4CjY+/XETI6zs4EZZleJ1X3ylcj7tpHY5A9uaU8w7o8rZ61O7v2Kt3Nx/n3l/
aD4yE2g2MCFuSysfaOozYZ5dMeuGvhvHugo4zBjzmMoirFAIPQRyqlBmqFgjtKzz
cDmg/ytlS9G+PoPR272JIFDQhwEHJsA2E3AfqwTVKfkxj0DRXtTXBO0yE48+NREr
3YXCswaR8hqvktDoxB9NvF7x7zs8o3FHFT7w7PH9b3q9NJVC2I2H8HXnQfaRxmt+
WX1urUzVInpEmn/BlOwDQ77+gQdeLUD7EA0X2oeo6igBqOMKY8hmzPVoXH4j+yZE
SxLx1ALu2lfnvk9qkOibJ2eu5ZEnl1hix1rQ4EAtZ9kPP7/nFpE+6zgO6MRUqHGp
x+WZTGToajtYXRPrMfeAJgxcndyxt3Tp7m2QzWTUNd7N4qjKOdr67vB32B8QF+30
1sBiurmjeUUqIz2x8INDPdISVbYbGa6xWYVSOlXzMEwgi0n/X/8DAG2As60QGO6b
hDZe0nECPjVeGofcRJqh41qNAhtPB3D4xBHLJxDAYgL8kXjwpZlIa2BYMOet/KJY
NIjoeTUQm68nyWc1N+pooPL24H3ajmR5Fdf9cgedeMYHmXSCDLq8k2zZfhu1Zq1Z
v1CsVfWnoVwPO7C5hLI2I9YP0NqBsZXS1SY2Zb9iDYRAHGjgRspYGUpfThd94xi4
xIXmafk8u1e6tVm2/n+7xL26oI4BVXFz5iqt+PyqOT8daj0v09u0T4P9RJJNfN3C
GnRVpiGQRFJb4/FjuMRMmFvJCIzRWnpBLBKUf4w/5md+8Cw+dsXENaXuV2fJ3iPu
VOx3c8LeODRAbkPfQNRBykNRn7WECWBy0wsUg2jNE9PpJ4YNyNcjuRrNaPfGrJq6
7AMQG1lQjKlmXg/MB690vXXXPVs/68WjVfJFG7QaqseYh/NM+6/mATaUi+/2tLJx
hozWOIKmtKSmRZwefwV9laBRI39668Ob7IcZowaNkcCv+Gemebh1eGzAlisMEROe
WipKNs8QXFbqv3561sdqI9gA2HOsSQDiqUUWF8CPPpsEtbfwe7fSdf/VAIlCr6jr
WZPCk97fkmj+vL2JwWfQfy7mECWfBclaVYeqXq85krVP+S1+QghtDrWrANAI24jc
xAqiDk8gLShiYRa+7bhfNlJ99P09tMgSh07fr11K2r9JolEMyx3QLMPpn0StpTv7
yfmBMRqN8BB/K0XNItPlcyryr8qwcJNjIlV72+iGVVmrBGn9lV+lw2z8QPj9jFOk
Xv140NomJyHGRHTl9/cGCsujjxyJwvoORYiMAWjvfq/zhE/vKkBLCOzrfxysgXq3
hEbVLSFZs6IFJWJvFCJATECyV8DTD45tWFvPmxpomHyt/m4KXkozp2gg4SIZY6w2
qspBiHkFn/T/kqzipfwDzZI2zCRQCuTZ/JTO8w4lt95XsF314NA5wopg8hKKXvO8
7oRXTJEn+KJhXCugxqLExv0zSbIkp1JHV1vKeRRczyWo3UqAKny9jCdmq5hiys2U
UFxAztb75ePjP911VAHlLFiyCpC55Xjb1qZBPmXfzR073NqwfCEoPnf0/euVpdnU
shvD0IOg+aoaF5D44pFAWSKmvqDDZQFrXQETN95X98O7rbVXzywZXccaCMDHsZXF
ybXpKFgUu9a/n6wgJG/nCqCTivcSBiqFMRaftw0oylvToKruGCqdzY4B7O9ceYTQ
d/IAKFMFA8CwD7EuEDMsM4Yx3QUXJOloVrd7Ky8AeHSRCAfxXvCIU9kTGdzKN/rL
C2ieXezKEPbRDptai+6c3Iz/mnVVmDtyvhj0WWEZl+w3SyPIOyPxbfuYr0fJiVEf
J0u4UUwv1B+mOVGEY8e9CPBDVpKHXrb4kh95KldIIvS5YuORPeJBHghJMoRgVvhU
G2wPqbnc6mLYfghMUPatFC2PbIijjyiUKgfolIW3TZSw4Sh3pds3IlbzLZDcNlHV
jLd9ulowAj/RPQCWhcDLGHXJfMP7rbkuQhZ2qyVD926vNj6paLdjH5Z4tAdhWiDK
3u+JojqZc3Jw1l1zVl61vx2IEl9Q5OzgwAuKwW0UqQd/Ns9S0FgYTFpXMRlob+qY
mwFus0+1r5q8tHGf03atxW3+qpdLVMNsXcrb+UHw6P5uOg3SdXBOpmRiP516eTzD
jRwMqIInYd7Kwf/1OpB1qbu0e6+8AWfrN0TvKmmzZLwKixrWtOh/5rOUeWeTzOQ0
6cGcEy+BEMsf45du9Hy/FPhMdXZjuDjw70IT9IY7MGI7YDoIMLHSIHClbWu/gghK
k/SP47Yd94UVipmZU37m0/Rjgr2kl7Gnbvq3S2aampysRXqCSxZaCLpeMKkWGwPd
eGLgdqZCc5vvharQ4KACbPRqXkTO/M6qjGyel/9ek+SS/L/++vm2Xr10MasOTnAK
Q0aX4AoIq9bmY6eN5Br/eElsZdC56ehJTXxFWLhahlvfy9GRHg316Y6wettrKqpr
UFFmqRdERxPN6XKoJTQghdCax6cfimRJKD/0ykipbWrIQKVligVBIXgTWiNoT3oA
uG1DXP12ZU8woduoe8CcTF4lhGFtBCbm/t8mHrnlla/5v0OJIj4g5mbQwUep1gWD
T9cptk4ipN2tCQo0TjDJXtbSHcdxnHmH93iBn1isM9EPzIbH/0vB+8bcXXYm9Ymn
phMlWZHus5L/WsnVWPFdOq59/+xQi0ZnwHZUYV7FjKhUrv+uHhTcWhGM4ACEZDK/
SrQszepBGI244qAbpL2dfgT2yl8ZNq5KrstL/dDrE+UVcMmESzlhxqNGnLafCI9j
mPpD9a67fpd/AcXn90wqlz0PImRXJbvoXUKeDWxC1oN6yoqqATv59bgvCYToxA5H
boJgUf47hSeJXIy5zne6LzIb8HJvLgc9i6gzTT+IzBJLnj9TGERYk8Uvbl0gwR3q
BBgvSXDPIgtYBEVTbFIfMEVkNrQRPkMivPrFwYtguxUwe6p+QbR05a+BpGb/TrZn
4SkufCpjVyYtyVzV+CSRkMLCFVsUI1XsRUbKKtamAAoD9jSAYaDe8wtwUj3lt2Lh
PDHDBO5TRua/g5cDlNQ+SIq8b7mwqq8mOkJ6x1npCGq/nYWfZXaoM0koiTvtOm1F
n89bzHEFjCvJ/bXcppqaDxWl+qQ47Gd4ZhIFzg1yyMVQu0oSPZsL3bIZ/rfsQIUn
gaXQeqjxZIY/p1ixE+OdfrMrcFQWhz8d24eCR4OQUmErhSEuNOVPa7Ux7s3eU/Mh
ve4jq6J5J74p5+LEOm5Oe+2bW32JzjmqKyfgVSKTAX1kiaN0dly0SCXS5MknVyE+
pNx0dfogel7KsVpZ00ALhA3UlSiqQlFT4nkXtXTewJJFYvyjoX/ACkjTWaRd9awD
29vORHPAe3gkwbqBf5BXOBMjn7hD1H8JIFPZr78pWZz9mkMRksWm0OwtpxRi3wNJ
ibIql1Q0e8NQgTU5GlH93t06L5tlniwxfpYSrFBBdBidJF1+NMk7lxSRkORHhSlR
JwNEgLcAQvnTLxi3GTQoUhMwbwsm2D/DhWwctNAbqQfdPTkBy/rh6EEsrrFMY8vu
VWIdDHvP290WSBQDxP2j4R16rHmckSHsVxlQ4uuvTg7tbEuZjIdN+4OSztVbd72o
TRZEM0N+Hx4iHwwF9sfsEghxeIugZi8YlBHa/FgsGZnNphSJaJFFsL/5sXJW798u
KVqFGmOlBdLO53O/tFmMi3cLVHe9pR95QPEY9852HVEkqjyhorGxSNScmmVYzfeT
6W/0p3mGHTa2j4N886i+zt7UaLaiOoOQD3lhQt8R2mMZMPLl7Oermd/44W3yILFw
kmVzGm8so0PlFnPlndh1EM0vmpelw6H/lsBhGJL+e/ePx28lmGC1JygAD4cdEtnf
dy26xx3JUpJga8lLruCZKraHzlGodC49MtwuYIzv93ASTbAG0U/UyZyG+GO3lVx6
QLr0imYn+xJhvt83RoaXSCiXfJ0qgumsWLza1cG4XFWLOj6+TDFBHuURDIxUiwe6
Vxan6K+uO86XzCuBSQ4Dmtvlj3m7xIvcgtdUQ5kxKVZaw64p8b3PrIJTT0UgsoTI
9HecNqQWgqWK1+K9izLb0YuxjlVAfp7k79ctm9uok2XgxrdcA0jF425/NeHN7OEN
6OH7y2p6lbKylruzK/UK5hUBYG8ytuUNfHkWCc+M/hf4dc8ZlW7mi/J/y+BNqs5U
E9Hp3o43mlpLfaf+RTNVJ7+WyCOvr0Ms4RzN0ps0xOTemToWwZ8JyPnAQJYQ5B1E
v/brdQB4v42n3zucCO3JR/b/C0zl6GjXJ8Y3g5x8pZlThvhpqYmzlnCwyIWB4zYf
6EdSu+2B/n7YinI4TMTfD1Sg5kt3xWmdWZg+49prsw+N98h5aU/PIucRWoXN/54n
DDK23msZUkTpPh2BXK8wJ0rr3Hh+BFYW9iYk/oiw09fmwbs7HF2q+8cmdGmKQ5xj
FU6quEOUzAC89uEkN0lr5ZnSwVlQSncQIhO7tGlrmc9LdBeEQ8A6l3EiF2Fo1fZh
l0iA9qwZktDquy9VQP7YvUgKWvYqp6kKQVkV73fp5KeI29qRNANe6h+EvQMi81nM
OiSxASr3NFWKw29+wH/0/FFoHNIKi/T9hb7/eoQ9g2HdmlhSseE8tzImbcrx2llt
AFbEyTM0aN/PmymK+7xH0PkTCO0IgncVEFELTzTxMqVcyhktCpT5WyYALCAriHJg
SZKwXEt1XuUA4rNvPca3hsNo0fbdPnpYsAyH6X759SMeJlq2us0zHjq+NfjCmcrJ
jycrWjpmoH6gE/DtHxQ9Vj7mb/zz3h8d/4W6A31vya9d8zHsMRnaWsLx0e97ZTT9
CP/Vh4lWywMUkJSQjZ7ilU6jKI/HEeOSHb4BlH17SxrpL03v5zrfusE+4db3wphk
k47DELcYu3qj6pnZnwd+aGI9Tp6hGrmxK7xB9y0ZdTERAS97P3oB8THJyImMDTRm
n4nsliU1Oxa2xJVgyvpmoQ8qG9gWRiIMWhu+PnWoqHzGJ7yW18BzqH/J2DZlc/R2
o8jHj2vtE9WJX2jUVQViLAcPExTYPvLJN758M55AIAWlpzPjQeldTMOLWdNyQSoW
6hltC9y9pdQYhVfop0BkGwQXa1/AAYH1ykPAaUnMnF+LUZTwKKlKz+J8UMwdik+C
DoAWA6sKUkwZe2VSJg28vL8a1HPX/GDreRSmLga8xg3BrVeMPzv7qTqMOwMTthtH
NRyP6gbUDNo0QLEV4u1XGbtExlKa4c2orMm/r2CBGLuYLHRBbjZxTdAhFy+Fsc1Z
oo9k3ZgY8jkHaH0IK5a4byNMRuq4TWichSVylkWqnZPYBvgur0+N/m293B2BTTcX
tHBpRnpaXz4LkYEeEyJuZJH9eub+ozkSAe6aNkphAlqtdJW8HRbYZz2/8DUgMC/7
U0Y8Tj+ZHUX6wPB1qHSGWbXqf8KmESXLv5OYRDldR26ripdFZA5nvJ0roIsD940Q
1o6irPKdLMgqQQ1xbqxdQvIYodZsSbuKr/f6an+hFfXR2828qnR05R69RHz+IRJ8
djgAfrX3vCRK3Zf1OIr9dxI/Geou9aqTFqW/MS/XPLKtH69XyKOus6iNAIuTbn7m
VNJ1XVZH5batKC4hJHvjdUQu2lCYNwKS5o9HEs3rGYPBRKpCRcOjfH4WifBSYec9
1XYDBNMwSuoUqEdCRXPlHV6VHPV/M/egZGhH59ncBF+pEmKB7TI2na9vJVLCOABP
9o6mt0p1I1SZ9ozMMK+3PjPxwgrvsm7tXF0MdvV49G34295lJTj9zsnsleRzfMxg
9l1ahNT0DMPYka5fbREWa+su1CcnruV9qg5cyIKyg9ktjr+gg+uX2MTOuhPTWElr
UNm6zqsMhY6vmZ1cH54wGd4dMtbAuL/9ygpDo38+EtZD6HZTJkc36eIJhBE4JduA
liFGTunSpLHAiBoADy+yTxCYMxniZjObXbwDk/Kk8Fjh7Q+uFM9oHNgZWRwZ6eDK
gMWzuN379P9rKijuT4yPDYtKd5AH1gl0jdi3pYt08DL6u641PS55eO0iHndTX36J
B2JKoZDA88o8nVW4cDULuoJAJ7PjQY9Ru+q7cx5og3CiXuS8JZFCm1udyyplg4k0
fyVz9fumF0wpxjUpuzd6vkF9bIw8jrGaWhqPmzP+SYg6IuEqvZ5L1oiI1Bv3m9VW
V5iP7ZbWBDrb18Gxb5aK+TSbQ9siGCvoMFOnpFKGoUuK2Rb0Kb4u1MX0osn6scic
e3zQm4YlL+Z4ReU7OlNjZbY8cHEemx+r5ZpuPXcq4FPlRnwXXZVpKgtpK1VG/TGG
8Q9/qkxX6uiurnT+CDwWoUt4RBkVAzELPEBwkBTVFfIK/UvttAvGgWwu4APNRqaL
gS9bzhb767mIBLbk8DEDwpWHpoeK9YBXcTvH/ytd1iFIUeJzcIk1nDo6h9lp5lPC
wCStm/IlCO98+tR7+cw9Kyi8m+//dn3MiyjASQy+rkENn2XosB5ZsSQe0KXDcv0m
KTAhrRrYAthcWzshpFkb++8gnJKBo0l6XZfMXZONNU4P+xdTYRcat3j2X+m/wMKJ
2Z+WKzHS7jqp0fXkrmnZaq0bYjkf9KpMqoePQx/OAGIawygu7yvgsOf4Xug3xtV/
BCtO/V/yzkbiun3eqFix/5mp5P14svipiYlCKebkXoVp3bVeO6OON4a9S4yGQddq
8ovQ8KoiRTyBX5+lBRqiO+3as3QbXhQ8li/9/Q/7Bkomi3+V/AFl7gpyT03ATBeQ
uSKk7I4UjYScSvrbIhmsE2PKNRSVDUAyEW8kunsqVL7hbubS4Na6kb6TWgTjmdrD
WJJNBgxmbEM6KAWHbceTjqRLFTWNFoJdJGNvzdCe9OXrFZS8XuwZVpkbrYbWsH5a
JuKvr/9QHmwbmqx+bmFwgBfQFhEdwfBj1XJLGVITCcHMqxLLL+Y9hmsRGIoL6UDh
VRXCCxiR6l6uMOq21aDTDv9jz02lVuFPAyMdFwqP8zv6JQuwy/EuaGJysXTQllLo
ZypxxPw5THLJWe6LoXm7HtPMaVD9A9u0wD8myPPSVjRYLbNJidZ4pIzRxK11MnY8
G1cFzmf1kNBFbojOVl81a5k13f0AxZqBy9QqOaLZpZDDaisIahsQCYwH6+jV3xKs
kbmpmT8jYZT+XMnbCnIxxsEoGGrWAYYnGBFHDFNruTTlKW8CRA5AAcdNziarSCXu
1JOxXuJVCb32OItVkD8J8CcquXH0HJTn+rvy6tcDULYMvXO2e8AM/dIcwAbtSE/a
5q6Ot5p6ue+Tpwxpz5meNoqwxK5wlXsr+lv4PvN6aPTqjFNjbJlN+L9q/kPJ+cDI
UTAshiltVGBQoRfCrCKYEGfJc3dpPZFDpcS7ZiS/YEjQsXTk/SMxuqVvvEoFEHmh
AgREVk+LSS+QBrAZ3B0Sb7aOL5BTGnrPn1Q3i4rD0fCtp+tFKpCCKikwi/89pDfk
SEITFLEtqldJLWGKniGgLc5kVb2l4pSQLt7Y/mN2ys/1wZw0yG1PAoS9romvZg4Y
YuM/ed5VAEOb44DuIHOhJuhKe+s/jpOiQ224hRcsZjufOHZESJMwsZwxyAwjnFrD
ZTYn+Ym9Urc14NWyjUVDvN39eqTp14ZzYJUnlP6SShHvP1ASujnM9egwnLmU6lv6
VZqr6a17ay1GOAOXy7QUafsdYh+U83ODn6TZxvUri1wCU17JvLgpp3L7v2Srv0Ja
IWsrQk529xP2luNpFRWBmqoYj4PTmaTKa4E5eWwgUp0hT++z5qpn1miThdi8Atar
Xayq5iI419adz296S/sSUctTIE55DKy93g/0AYuJos9P0tTF0tItrgRZcZk6CnCz
mhJpSS60VeNAvfO3U1SzNa64qoFJ5lZfeprRrdKkqQQ75tXKrc1OJZoOTUIbpr1u
oIoNlpxwEr188vQea40DS6XyeK6z0+bt5mxGwji5VlFhsR8s6EAR7PaNbZMBUizQ
Us0a0WQ7gtsx/jIRAFCFmucPTxKv11k3BdZ+teIp+UxlXAJrMpDiC6Txz71wxGg3
chvKTZUA5ftxQIbXb/fGV6fA923HOaqrQhEJ1jFSxGUJFnEpoy3bJNz2uMb6dgm5
KPPM1ybO1HOFnQlTuThmfJqeqilQlTomc6q/aRUfVYqXueE4o9gF8HaiKG9vaXXk
ipItSWDmx2A04Let/DAMkjhUL94WErKohTxgWGQGZeaCO542N+d2dRjT/vqOkdqZ
0NVGtGSYOqzqvLAKKfejHNCrcMWOA4Zy1Tslh9k6r9rw0InK1lb9nlaEp8E3D09a
6UDsLU9gApn0M3L/EmFQJZRKN2MCN7OVFaPu2Ff3E/tU0U65uvFAoXChVLrP2Fl+
igkeBQUv5M2IMk/zLOViagmqWtscjSUO4NIuyBiWorPHwY49uqyaYjR4w/TQjYyR
2VmT0DzJb03zg18rVKoss2K+4SyRNxh9ZNl1nfNUynTL4dzWr95OxYUfWSNGmnqq
tyrMJdkPMU0603eBDQJYScausITuPyrzsKYpHDAEyTpNIrukGXJFsCRUX9ywmCkH
9BuXRPHQ7CwvIY/V8OZFX/ojT1idK8aEUylgWYugC4/LVVyV9lYL03kr4mJ0pdAX
iVWPATrh3e+u3uydYxn/PGIm/fdDcuUrepDztXcFPjwIh/9/YsSRgOoJMUDQ9az2
e0TX3DrzfUROAJ5aCgCSs0TzH/21p8qn0/ARbOIT9FZuxjT+m6XderZ1DwebE18c
LMH1UJeO7oujQNcaDlQL88JFq3/tdiXO3XwViPLRA/GVA5QaWqyPVarxjqhN0KqA
+Zk8s37z27ll32GtQcqxFljLGA+2MCGhrwpjP8xYLwq55lkW+7HnNat7k0tgIB91
hGzJjXg0d9TKYPIRLcyYqCNQ4trE3coXhUDPws4GvwflSnatsv2r3Te4rDmj5z9S
K71O1qHpC17UCOezMjRcP7FfhvNbd5P0TDHO/W/iIGrm6NqaxgU0k1wlS7Z+6ogI
w4fYJN2wS9wn3sWSq4XcgwDKuqy5vvLJGAzrrCN1lP3VYFGw1bz3Zg5+upDOhVOS
WjwlJkEl0FnHuB75VbZsZcDOlWwKpHUD3QeOTaoqOrXaM9xLgtRmSe/il7g5v2qA
SwUefw0I7FR5b2VsbJWLFHR7ykaCzm1DGY4JR8vquQ2dxDV5jUlsdTfUsRQNbVle
W/QfKLA+aYiBLbJCiCfOiGOxf1qq4z1TTp6Yd5V5T/ynV8LJ9RBXKmtKLH5UUIFw
gA5lXFX6vbUlFOXtnnXCQvUNjE6sQNh4zdTmQ/2L5Eh4+2Nvg9Kj52i27lSJRv77
U2OXbNUwRDs5x9gzRvv4TE5Hw4ggbOlrmDKZbKAHsIIMONfDsW8WohqRUMYOckbO
V8tihY/v/1LDHBfr8z5N0jM2IP3aJkjtBi7CalhNE/09XvPlt/9bLkgMyw1aZRIZ
HioSMAsV+CCrtv+gmfNTSjYhg7mkBz6pdveeRwaSX9WMIDUb91DYe2b9Q9tzJXCy
W+8TY65Kmsn6N4CFjoNxoCiviQ7EM2HIW+iOvoxmllOjaXwncAr1p6Hs6c5sR9jM
LaFb8mgVCQEjmL5YhUoFGDw8j8SxreQW6cqIyCVbTkaQhoOJ0M8MutUQde8B2FXC
7lQegj+lujgTXURtBkjNpHROLLMZ2Mw9p3Syt8q4LGl/Rtk0o/ep7MwdcQy2JYvF
KOfhGIHWrzo4VNCsJgZGBMZEn+k1Z7b0LpwrnM4G0kaw1HO/BuzN2CTjtEN0vNcV
WaHJgxo2la2oSDenDCZL2YugrdeTQfTwxTJxwv8/zRJXnmNDgszkIKaRbA+vjfsf
TEXtxQjL5OhIqbpzcOozV2fu2Js1Ibg68ixS057bQbR0ucgY7MUOztuFaOwgZQ2f
UC4xF7J7Easq59W/slAfjdLKelGemMUDHctTwNVAghWW0vP1C1rqTTYIhqPeW7JR
Pbwha1GGK3sdyLJCJyJpZ2vwUhA91i6bq9UoB/vvet58XHOwy71oeYqy+HEf+Bbh
Qnf71uy6OC7jxfPsOzVzoEr11D0pSnyQkE1UgN+r3P4I3sfz9/FSAkjNMLtNWBb1
3eQhLs+rKF6xGHSqOeONZTGwMHbd9auf5Nd+0waI63vJR3s0SFTgIepFXQs7K9fp
+1gO58PjgGh9g0CZ6KASB0izzezrDgVHTvNTUs3f5pNHEIUvC3BNTnxuY+1pEGUU
h5WOsm/LzB471ZrG7aiZbdz5Z8HDQBxOVYuTy4OUTZGooU2M7k67lHhyDx5kPQMI
V1jFRyCOu93tolPTOeR8f5C8onuKdAotS+H8ySA074Lsr6cWU/ywkQGyjE3DFDUs
ucRfHAfR90GosAfkeG7UK3XJTaZ3vEuhmK0XbPRpmrHQuN4JfDV7lYfxdbMyip9D
Y0WYQAdUt84LYv1Am7zAIyhueIuP6+8dTKip2rcAtWeWNV+76QXM50oplaTYyciU
e/VsulgSJ32SFSqeADdyFQ91EcGZRFJaRdMVA3VPp0i8PgvzJUDfm6pHX1kGGbOl
D+AaBNl++8wi5A6wviOu3l2hQ+k2Fut1sHpaY8S6KGYrmiWG70npKfJnq8rokP/p
8l1ZlIZQ55xhVduFlrOHO01JfK780Tjyr6Qv8UYMjq3UoPdzFmkcErqkrkRuc2lF
MxDnVVZFW0d9i2A3u93yMoi+/CbCENiY8WL4XgL/8VQ0vt58jj+IX1R6F8vQ52xX
fnP90bMwQPYHDJe6J1s/mmo+KVZe1VoIKNXc+qI3/RM2pNV2WX+zjGrebf44Ldtd
9i0tMm6Co2m4sJI986tqijqa7BjMjghJ+TRRiNqf3/hM6vxqeyjuKetSQMYRB/D1
msHnuXchCkUwnJXNpJNBrfyklxnqMj1WGJdeU04Tp9QYFVqgnJ1of+/nZKo3wcEq
vU8JC2LTtt2Z+PxvJlaeS89FzSU+28FYg5uOhZ+f/hw8DPwSFVGbCR5vIr6q63bV
pGVVLCCdBjbIVA7sUSJhFZPEtBYcNr2zC7MJCxJvP4h6ZJH1OJIge53bcLzaXton
qQx4aUY84jATu6vVV5MSmcht2u/2CKJqPV2Rj1VLR3usjOdWPe8p4ShBscAXy6j4
HteoWpV7Htm2u731+rIcGqzM+0f9VCp7aYDnTAwNXX8WptDKOp6WlqQPoHRWXwRo
VwJwomLbHd6TwDO0KutmexaQ30wwGBD6IRzs/UO9EkKZLJseC8x6KTuXjuWDkwrN
JRGSmBwH3h7Q2r8pi9dXMvEWMDNaRLGW1866oTQYIobYQEU2mzS2sriFb7pjTaeF
axORwrq+BYmkyimt5p5v8mPt4HEXqEaa2wL/yhAm545B41aPyQbe28MMEu1RKMWp
sBQ0+PKy9NJP79aO9GtoVJ+nlrX56PlsNtIgd8eF7f8wSfWWndydzYPBIZL3qob/
g+eC9/MhiLa6XGST6S9ZY98sNETaCq+5WiimJRgbMlAWHgLe62jO0tPHBg98UNWI
XFH+8GR4O3l1yOZzTAFbaImWTxYv1j/oRRy/6Z1OgFyxHBNuYOpORfHwOvpQYRY0
kx+vyFcd4xoA+NnE/Rm7C6TnHGDRPTdHues5m981Qcm6UhpnTj7qUKhjlsDX45UF
MvO34TMhoilw5JEzXesPqiAHw/+Kmj3PDIqcQuB5ROrqhFyM+TLVQDaVmr0rvuN2
AoQvOCwRXctYXUDVIQna6Cg1L+GD4JRYOV4luVUfKPBMK3XWHljxXwdwRRq0S60Y
UWNT6UOcmSUi6lqKld/awMaYiq9C8c8gXlztgwORsqd8+jIFY2u9RpQbSm8K9UoC
4rj7h+D0gzhTqDMBFXNTTyf6XDwoAE3Nvcmu+s0jjoMiS7nne4pYw9fgfwG3I9jT
d2swQ8ByV1exi2pMXMK0Q/JgYR8aee06VQb1oWlvOcedagpw1hmCyEEfBzcOmTIb
dqyIm8Slo/iJuwmreTyP96QhNWeceCkIBkfyHoGqqnjbowJoMgKD/ugpUAhJ9dNR
S+ocMhHkur2iEjbqxzljTy5mC/WzNqDuH2vj6OEh79ot6gN8zO/GM6KYPj++bAy+
mXeiOi1fh3CnAU7O0aNLoRXd+hFzMZgvX9AchX3y6bdUa/TMSrQ3r/g2KM3UaGH5
kqUo01dzSsnQB7g8wl5rTGumKdCFJh7snHlW7uhTJc6CGXFAnqkAdM6iEkkRMvQD
Fl6Lm3fbDEYAG1UioL90ZRONPuhcyFQe55WIZ9uJ+IT53vuvQRcTlxHvHjlM5L/l
fhdzE8EmpF5EMGbHy92uo/JghoMgQk20XUCSgLf1YbfFic1twqwXbr8vup2v1AeD
JxBcxbeVSxc1lx8LgkPLjdU2jObLZFmjqt5TLcpXX7Hnl286A8yOjx4br+BW8l1j
nnEhQjkCOozWsLi+J5asnBTRTTNe4fbLSPKemHSgFIOTPny8nHJKqlHmwHghPcWk
D6IY1Cd5Mly0khI2tBQQ4z3nzo+c9XEY4Bked0OVVwfpDJ9EoDYUAA3dfOTPmgoU
x2BOFApNW6lRXOn/1N6L/Qa6dBQQFdevkHoDI9xInpFHAXVHEG3AUkdk+rTTIj4e
2u4uJDHyCx/P5IGLg0XVW5e3K/wdO3kjHGgaFPhMoRttSdAeBuZowswsVg1gIAfM
1PiyO287r2psMfN2jtcJFu+m1LqBumlFRP1ide8qhUN+zO81IGEdTNqKqPdIrBXL
nxC00o2lOk33tkdAyxIzYJ97JqTmkyzkmtfkrASSD9FxFnwTh1Jf3li3szMq9h40
Z5AEqFZOzwdJ8tFnUeQYvHxs5KTgBREf3MWRvcmzFncyfCUVJaS2IgF0RQMt7WrV
llN0CsMxudilVyJrQne420u8pwKGb1jr6txDYggAuzJRkgqTpTIrNMAXKS38DadA
RL7qsF/wTtcw0Dz9aDjyeG9ggyyI3Gi3CdiA63CTQ4N6CiBz7vTMZXW1Q1gl60UW
L9jUT5SUYqvS2zL1wOrqZZ9P0KPgGn2BthNcEzsl+SFWlyGqEneH5oK3DhsF12DV
DDyh6lqzuBFP0z72c7EQzhQiwKRBMUJZXFjmuioV8fl0fMQiETs7UwTeXRec90g2
Jdd6mKrykAfqBFmwF81+4v9vA9uLDGYjhViDiEWoexQ3jmtaT65CAlwwcf8UlATr
ZQBAppS27BArw79YZv6LzynOaLO8GMhtsRIZcFineh4qijJhPL14XPSIKDO8v4dr
fLjwWz2AdmRO3m0Jzvq6H00dfkC91L4ixf9qYkRApOCM8jcYIRqxpiNthu270xKs
+o28Skd8aYqM6um76H/RnaPY5yF2OVSzBy37u4DSheQ2IiM50JiWHaMsu7Zs5yNO
t87TbXmUZpj3RcwieUI3G6AiAbSbDjYzwdDjWtQqoSAUDIWaAbE8MCh+7RwcSk7E
LDlXKVXB3AV43GuD1+1M+7fx0K2W9pKUYFh9h5UqKVMar0/ZMUx8MHKooqIOgT5W
m1PTlvbeePHECHSMGh6yc5H3AydC5zOJZVCccNoJ3vO7ocn9XrYNhSWwO9NqAXAR
t/H7+7A+kexqgrfoQ2JhPJ1pluoVxGMWAiyHctLxn22/YLtbfjxvvQwjmIi3cOEu
EdahGcZWlbCqBUU7qRfHeyCb39AWURs7vCn+9JlH2URvADxvxM7/riWaXORVH8ml
RRqGHMnw+WJqCKWJJZ9aIZE6pLd88gJKzCwxqJEMFZEg3ojdj2TanzZ+YUmjlEIw
Xe1+PR+g2d2Lr1N/KkrPzLafwB+cYn6DFvspKNLNzmWyE15KACueNkTWVVUre5ij
MuuJSfEiqN26vMi4YHOklV/R4xT77xMDM1XNuLwRrn15skA2NaIroAosmK86V84n
CsadvggjX+CKieYlUIv0UIaJgCKu8QNJ7nKgnA7tkaOUbDKKCMwIsg4TvjtL8O0F
nQJN6uVkmmagL1A7F3sO4AkvCLDsJlED7nbseEH4cZIvg8fxlBAc0Z7m3ATbJo5W
hLVIsweX0CWLoSu+efjF0dPwHZ3VE9TgpWv0NGFDkOBrlfoC5M4f0btOM5T7SXd0
BqxrRl2vmqCWcWIH3enCC/ysH/6TaV21afKhGJ5sp1HkraGnyRbrivd+0k0XfNUW
y+/Hp+HDsKJchYv41xEtLlgArK8fPWv/rifjrw7eDGWmRAZwJyM+IzhgbCoaODOv
nFiA46xepJh97lSAIbNq8KRyVKJB4NIep0s6IDdfhkANwBoV1XTIFEq3H2fxxEKn
Oc8CzP8JNt7ZiT7oLBZaURngQ87pS2M55K1Z4JlTeC+3ehJ54i2GOIhDfcGeaeFZ
NQUgNZScxbPARjkqL6qY9ffE/pc/EPY4ajA2fJIzN/K+3ErS/y2dYz0EnB0HdCFB
S+VtnT64ublwbEEOEokMV+D8uWPzd3AEuZX7UPrfm6Knlx+aLo1OY8BlRmjIufLE
YsS6qj82P+3cqR6cnPwO0aWsFpbqBvfIVBTR3ye7HSXxj9k1AUxTzu9nuJyizfZU
/UaE310wb4OstgVL5tvgQjPcCZQyetGBbYc8Jkv1Q6rO3CPe88g01QIXIOiHbqwH
aZdZ8fJTsoMbbrdqyv72BBV81tEAlvfH/AwazviVLvGEmePc4pF+5SjAFeT8aEkl
jvJsudrLKWnI/P9pYQDPK6bxjviBMiatiOLRuYBllh6xsvAaSH5xUF9wJE1bRQ6D
GdKAVDtl/zH1hUAZKl+LCQTM/FKzHnkEG90a+r/H9sT8eX8IlesnDoMwqiUfBj2F
1M/oTKDlqoLHfOpcwTUhrT8oSbfBQYOKeF7YFKb2fZu173U5rRhhpAkM7D6hfuu6
9WmGvsoaaSSLwF+5dITXrvN6QgNGrYBRH+2OBAwWKxSarASJ8RaMji/5+13HBkfC
rRrS+ct6vjjEof0L4rClWK+BSt7xvkY0RhS1TdctluvuqTsvV+FFaewNgKPWA5MG
nb42QmdUW2PwV+YMyilMbQCa98EzTvCxNEIZyeXEsNhm4aqrhZkk01Jrqz78S/7t
afE/Q7b24230215Bg77aF4JrnxtOmgjDAa/VrOSahAD5uXmnerdSpuP/KOiq5Veb
EUDPLNa7jwL9WQUPf0EfIS0vgUOu/m9C26ReGXbXf9mQRavqlVLm2kx2czf32te7
cMF7YBmZshIHt9FuLFfsA8sfPocCz6O77JRIwm9Pvf53ZuoBGcu5Vj8BzGSEQ/J/
xBwGmjv2+vZWfuMJqWVfFZikDBFklpTJyT5slEuxHXYVJF3o743iyJSLTThgL8nS
9u37GAXAngHiWUNc1fJVEPpeDIzdD1ahKCi49QIO4VKL5dNVBffbzIs1HeKBFqga
UME2S37h78bRQMT60v/G3mypstga03FnT/wKMVhB3gnojdkp7qERV9OJe5FR4GES
DLYMRivdJIwOsgVbUsubr7nmRwjX4Z2cLQOwlwT95eGfkZqpiUL2QUgQItbzBBav
tNIgnSqIAQukJf+JHdbxo2nmcy5QwqIcecG7m5sBNyPdFwzOBvqadHDb/sYl6A8x
qqpSXyLt+mNAsw9Yg+NIfiTUFOWt6iA7SG5/+JQKS5/QrHqPRydop4p2/HSwnGbY
Pn3FF9P0MD4uTnJf7M14HJ/uLrQkhi0xk16KaNHVjlX9DWPsLL72/kzatvqdlxiC
MQtX8giS2cfA9oaws3XJv8+g/EkLn0DUKHyZTMkDxJdoOUw7NTdWrK3daP4hfz5u
Pu5g3yzXRJ8BQNl2oAOJhjT8jX+k3K8LcKYGbiZH2k5LjzNpDqnOFuCIKgtQ4475
2Q8q3ty012rOZxBDlE6gKwl7yOQ+LbfDr7L9wnks+SZ0CUlU9w3Jp4nlbDzCkUXj
+hU3Ay1qgM81ouUWJ/T2r0dK7xYMHl9B4eNCWuUGImjbdxtsotZJNjpKtFU2Hmvm
SzsuE0DD1ZS0WeABWXLNHvUUzOg5NK1hmQilnSyCbT89WgR/T9kTm9ncKZLmd/UJ
An9lr52RbNrbozwqLWXnIhyOVCSIv+xbOU0/1yYPXsV8vw3eoNjzLa5ywlZtzfM1
hAa7kohYDDIJ9IpLuxn0Y3T6737kbKcRjrnU+1l8H0skUSD+jbc3a4K7B7OEF0Cu
YrhKEmpiFB4g2dBAX6QQQueOMd3bSUmdymHIAhOUeaMQfbnvNMeK4bYEaHBqxF0d
u9J/+lT/w8jxEHAdNAr/Twf56BnsMG0x62KEzvTcF4ZDuRqN3u1PH1ej/oTCv8zr
lIjSW8m1GSgv9v9mP/sf+Rwx87I9TR1lYlR7tRs2JD34Xf11qvTJcuAX3zNteB8Q
+g9PC+87VY1uFOPqkgq1tn01G+1KkE/clImGGZDQhskh2QIUNMCv4HpOutLt40gD
AYeduDKZRG+Y0gyoD9gAi3bvwp8u4SEetmnzYMVsPc9m2qa2Zlj2boxNyUT8KFiG
eq4AerMcqiusysRWMEePGVxB45Ei1ofn14M3R01TolyP8QC1caeCQiX+ws+7YEsS
a4nFtoDiA8qIKeMgqhf6wHaiTvcbzQTjbkUs8OSrv3anuN24b3IZmkRzxCp9zodI
GcA1B2eF31S3fhDrZKz9QO9WfhRwgRH6z7laga1jDbaSIPcVdi2DWN3u0wfAg9I+
eeU4rN9/myGA3sigS/ttrLtL7LW63jAzYrOZ9mOqGbmfoigIljA8msUYwco9QgGS
l7CDGkcRjfq5Az44bIcDDMewp0P++FM2wHjWXbAQsUeMa605dY25ULpm03MKdu/M
OOy0bowNQ+naaNMw93JtPNxftIK0cl6mlmtG7eBFvqepoE1EGqws98mtCN1ooBsv
Hced73GMNJo9xPK0aue9auvSQcOmFc/tM3x/eM9N1ex764MLVP1vSEZ9/bzAjOLC
K8ZD+L404MSgo2GVEIYURWUosQ+LWLR4iLtZiUK5g/oR9+Ur01XHmtgp7o6sCBZn
H158uyMpO3lZPhsasQSplob4kjCWcxAb66YRvnqLBMcXmNVtX3YUGaB06XArsb07
oLsO/9d3Cn9TF507lNdbxobCoXOh3+L52lD1EKzTZTJNsZMX3SSNLWn9uW7iEISV
CYvqEPo/qZSRjD2pPQ2HwAHDFecXfEwGjJdswZu2YqGeBmYgQ0qQxFMsPweyRqqn
RrNkRMle864PDlO3U6lkEqL3KvxVTAgwjpJCUrzlWnE9XpNNwaEIW1ozlw1j1wqr
gMOCmOvYLh3bmy7a4mk0+MSHrlZTW9XcH5bs0AR7oH36lpRmaPWSLuzCEqegxRPO
g5DNm2P7rXzlKkhJ+ohG0NB4sNIYN0vkJ1SHWP5rxX4i+9V8D5SKgt+s9TCCLiC2
c6i7ODNwP+3tRI1til+4AL7AFCtKhGEWjT/0iiT1u+ZOv+TUIpiL1lwYdbTbABwr
Bnb5U5EKIw4Lwrk90TORuVksnHNAKU1BA/5Hleee+M9K8eQsfIbDN2Ps27sVCmue
NxRCIno+prLTzMHlw3Adgh8WKU1Lh5//kYT5xSw4fJ8B33ZrzMEFusZqiIRnhDee
L23mrT9UvnAGRw/AUhnOFOdGTrQ0JcmSKTvxQbJ42t5THyBcFfipYKFuMbzDuuRc
/Sy1MAD+krcIQ4YnH6iC0rwX8SdOMLY9+3/oYdVwnMgtnMhsqoRvMzTORKXZdJeO
u/phjQv8gDKCsuj3YieQits1y+MYrPV6aKCeLA2Dq+1Tf55ONgXLMBsUROf7HmwD
w4I5SHf1eZyBAwgpXx2q9tq1a2OiEwztDpfxqAfeVN2YUWnd8OAdOIw2fiKYnssO
cCFOTKGL0kBh64pQH0o3ZLRtgOCWEbGx3uCaxSTLx4q7xRxTj3m+uBp7fisVD4z/
nMkvU7jUrlHjSq6UOQz0iq+BBYlwMox6SJhqwy+Q7XkVoSub/7mHhh/BbXXoMeBz
sFMpXdTCGb+hBP3SsmTjyRr7gJk8tuRrFuYUgnWEAQ4iDMw3fEaj4CDVN/pPTh74
gN8KVG8ay0PNDcgFaKat+NmPgCmABbSioBWkOoBmsUW+4k3W2kijZWCURjRnJinM
WWXAPrRiMGcPVmd308NNTx3A05ETNgrqBFhJZU4B5GPe8Xj2u44RPEsFFlv4UrnJ
zECb4A4Ipnv6a3YKFlj7+KYouyb6UJ+luhc/GnfDt2bkgbxmtMTHICYmrSVDL1n9
t6BwyBdgcIMha5W1Kk//iNjWguE6G8puD7ah8q9W8SiGEtsLjr/L2k2Utf6iDKLa
sqeQ9mjiHg2H7ympytKfinuc5YkeWhjj65wrtrzStS99mgwFf96JYdIebSgapBWo
kAvbUrhh5GNZEU90TJbSDIWPqDslgUawMGtaEgl36xQFzUzWIZSpiHDFMnYcwwfM
osbc6riHNG0imP6qqcCtMhvC3inTd8H8nwFEJXfqnh3Pb1F90WAPKZy9p/AdK/Lc
DRJyGUgXqhbwqLKmiz03t5Zw9SXYXgTyjw8rmKt3oEZq2poPVjBRpdy2uD5eX8KF
BZJQ1UBBgc1D/8stA1DBFzpYYYqMlTUskv2IWfWhiL+Qxi+KTrnluCrfHmzdO+ms
a50TlnZo0v9l0RVXIpKmgiFfDffrsJR0oecrOEXEWMUBavyy+EI+2BenxGsXiGwA
iQJQ/JHMY5HLz2lUwVthhHUNLY009Rx5Bhg6CSAPHH7sjF+g1Cw00ercPx3F77hY
wxi++CKQvQvOVtkvVPHQdstBvWEensL/JzrlqzFVXfQyqqd7BD1Stt2wJhvWEgx6
FtaJMzzbJ180R3kAdXCac1v0OUQT0IFGuB91oekcpuYkxFkDPbDsJ5d27UwSkN5Z
hwFbCTDSg8WVflrOZwEeOmn2FgECcCDGV1LcsgrWTQTBiMfSh9gTdQ1GQthmjj+W
UETHV2+uNqGO/VdFx3pysqCohDw0/eAs0USUCle3x07BlEAvJ3zw6nI0TGqPGFPX
nrrLRLgcQGRk7ywQ2zKWPrHcFFFc5WSgzWbGc54Ps3NOnDwa0gAz3t+MhBciwdiC
C3glw4mYcmLeOLwZDw6rxciSNw1I/cwD86mWkco4ak9GyYKXgpUA8YJwIycQDPA5
yRKCP3IEXhod5cIkoHTJqIrTGw0Bh97uAVl0lihZqAYo+wBNrZhUr0Y4/j5z0qYy
XNwNy9SAWfmpeiH6cwhpluoGHLqPwfsvFjeDl7Zqace6M7iS0JYVSIwcA5bvWlwI
8Hr06XGxsPKCjTRhK1gZ+IKBh+MToZFDi1pPJME9WSZJUHhr+RcdpAQwrlTbZZ0z
3PskOYO7ttiNPC+/JNn5Th6dRQjy0UL9SA6ZC+fFtFHyd1Y6v56hblT5U0aa8wlH
2kBpBi3gRtXYJNk+XxpHWj1XeLFk45/VsJa5F5P9M0IC1EsfPCX0+tiDKcgqhYdz
0LS5CM4mAfZ0yTk7nvqSPIreMKs4pm3Mc2ReRxp2gqIoNE2o2x/B7CL41yOZPWEB
MCFYZoqUeiDGMbeOFBlOd0TyEh7MrzJeRGDabcTxVN+oIzFdjZF1+xjewQnnejc/
tbqWMjL17MwK88saCBhwYj+7PKOZuQMA25xt72SA1QdWPLULLlSSj3maxkZyTHyr
sdRxojOmbX57APPH89WSIBHL08TyLtR3Yv0ry4v+ek1I9hQNF6Npuoy1ohbqxxi6
O1jCDeo0VgrfrCEzLvFQsz2jJZ5fwo+it9UFcfSYYCDBGUltiTaGk3zxN0bh6gWg
DqyAr2ojcJThTACU5+Cl12PWbgx+NTYKGfpeqXpmBRd/yKrcOjjXgiG9R6AiFMDm
vcIG26rtK3MYxA6t/SIxFG3u+EqGJSUxJvtv6XdvqU6Mk/GXw6Zn/wTvEGpvNueQ
qFsxYw/UTcMi9jvpFPgZ1qqYaynsyCJ7uqax5PX4dr6SKsh577/GNIQnom6j4BpS
KYRH5GZ3pRhGcjWg+b75HmiqVD80IwdFnLFnLT7DaDb8zwWUje7AlNjafW5Y/LuN
qHKS4IN5/v9M2lvuAWaKTUbijpSCaZDAMDlAjRFJFNGEPCFLXETjugyoAoE8ig1R
3PyCBV8q2xwm0JcqHiLhrscAOtIUzP4ojCb9p/kdO7DhtP8O8M6VAmWZMdGB7G6N
SmQUJsPdyFjcOBIV7HY6FMp6n8W2+bzTHAq4DGyhYwVdFG7SNr06ySwMVo8qMfZv
r5VfblqMTOSA5QCnluBT7WgOHewl5gDrQlT1AzFA3RSXXt7zTfHeRyi+7tJHAm19
71n9mNAngXNzldxlF5WKSlGv++bieV5RLUnxiHH0JYoZaFrpsyR1VRuWo2OwdMWo
CO3rAjBwjGMmBMpxcD3lDPzKZQoIc6La7RP8VlR5KCX4wZQ46eDDeGHX5g9jaohN
ih+eLNVdkHW9XMCgJ7GNvawyscyBt3AHKoviCYwuFBSTEFUlZBzhfiemrL+keLWc
5QUA51UjQbRtoCbW644jBQi4zyPMan22iE7aEKbUMVXTF8jaTo5yN5f3+WwzE87Y
UkNQa6mhu0diykdP7GhAxQrbxxqqJQxWvB4FctxtdB2QeWhWECxmezjDZM4jSxGu
dOrjO2S/eJtP3dk7QLOoaK44YPlxFJs5hIctS8Z4+N3zmi7tvZ7OB9SfG6/O/gmd
kw5GJBCUhFqq6TmWe1go1Y3OTDNYpEsr1Lo6HhaF5gdZeL8fentJc+Gd62yqqVcZ
cWFoaRC+LIbJsrIjUgjUh1fK0mI2Fa3WWQi91DzKdy5p9eYvqGbUYhv2AMHA/Z67
ZSL9nCjmJZNEPdWl4FUBXHgZSIZZF4UnRqm5i0ei6W5jpIL2VgVH94eFArIdHFwA
9AFpeFjgy7KKEK4QNyzUHvc6U57UabnIeOO82oH4Ua1bJjOgYBizUfGTslieCH4g
eeLflnMlYOf+u5dPormyoCrK45QDDCBeM8WnEd0SKzoBuDS3rQ7cpX/9RGEvtWQG
xTVWGj8MbBi+alIkWxa6nQ/ptxDNVGlqF9bf/cCjdyPQ7vqQZGXfdUUbz/ngZh9u
EwnKO1VEZbYH8MNbSNdFXYOz4G9EQLeN9oYUkmIpKM9z6+IHEqV4iEh7cSta8Sps
sijSFAgu9EwVZ0H7Qhavusf9a6oyECsp0BuF5S7Ze+oYGp82m1lgmjLupIvUMw75
aquVqZ8roAUEumdVAVVf9uFXBjeImuS2L4Bhps1xLNXpEJ8KTK8oJfZpNY3V/Xdx
ALqHu9GiJ2UQX/Y5Uvoak8qqIMSCzSp9nCcdl53RIbrAHBGmhTiiCftRHg7y5FRE
gl0ngHmbruYLmQK1OnQFboWCQL3tYuBOH5p1CpM7Eore8dZ+7Uei05BjKeQf7vZ2
cykw5GYTWJA6ecuaFbB+gKx6CwdtbOMsd0wLRnbvff+L0GVbWKMDEHTDZoSvuDui
mpMP/wxOEo1ivPhfiIlvSSDk44FkMukgDTvzzGTPe91BtIx2NzVlAv4fK5Va+BIK
8cJWimK3d7l0zooEmdPY4QZArI3fmF6gag57rfMYO5jhoQGx+uTwMzJVg+9uQVaD
gL/CSVzQRDtymtFcUOo5YfLDeQ7PcOgrOYjLbFFtwTdT4jMjQqG25y/XuT2glRtY
66WAU8TjtvwOP9ttmAQ6eF1v8IVRu14Sf0NuDQE/rkszMQ12hyQ2hwEbe1g+Fkkk
PC8fyzziyTE3PUuchUPHXVfWmaWfytkbwjKqxDf7U/4PWi0q7ReRgUr8O1GUwh+u
wmU9tbBKhXliSZ9yeLJuUXveOY8oILO3MsmW+U6adJ8ywmmsnBplWN3HHx52MN8R
nkk8H//wwBmG5TeBRjifd2fWKNATJikn6Aojo2adpgUEBVNw7U1VqixCH+2vYp26
aVuyJSVSRTP6tYpHi++40D4nRMolv4B7NfEjIxKDWtiiBQ/xHaG0JyEy4j0/9Jb/
XiBNwp9r9dAVXkOrWE56HxE5mVaCabforZORUELpMpwgvhaHRou2hceyJbptF0Dp
hMvf6Kfljx9qm7lgpOGSqPkqSxfhVlVs7jFEMHIoh8HV8lFOirNHMwThSsjC3qW+
dl1+nKsQrgGkgEywHUfdhieUfHefh4JzvLoz1G3pFxRrYc/72ld+S+/Aoc1s8cWi
E2Q+mf/r2+NBI+gVFz7pWB0He/fZ1BlWpIGoTrJDgoCTjMG0E/tkrcaIK3oxAS9/
nMkkTnwggiIDc+DbqZMNHzlp0pL4YP5coinL4yDNwx03PusM43QccHCWdW3deZrQ
beLD2fVdFcxfnzwCohebyKkF5XcwDpqfW+m5VORdKU4ZuxPdyK9W05vTYM/3lOJT
wncKDgFSZFccdAFuo7CRqxTtnixKfvN0f84OXc6DrfNQH8q8433snq3EaiVFdT25
hfRZK1w4c4se5QTnsSLgc86B8wd96vyXPtDrXJx6jegTbvF/0f5GKDa6bV2LytRP
r/wmG71AMFuVFRXw1u0PevFRHGkM+GzN8lN+Oa9vThm1h/0SHjoTcI62kiuNFXV9
oQy3BdDaMPFsTUaH4FNrCTL+2JE7AaWqQLm2f9IXaHq3PI1hDjkDqEFC1+im/3gJ
7/a4g+POqTxbT/bawZNArTZ4ETMTeifHMhB5jZp2fwTscH6cZ/ry8DhHvEPmQPZa
xJDfuVQ3mJSfjdfZSb2gbqnItkQbDABbTBM9KrRZau/lvld8hWdOVVgCufHsSpKS
5q/5tybgUoAQMPhbnbj+tXAOh0S+5JtbxBEKhvAM5W3rQgUOOtLdfPdmpMyvzzZ5
Q8vszWf57y4ua/IpVFwKO+vVdDkIm0RuXiQUaSUICpsTf18VxPXGN5lIskMGSdW5
okuy41gztld10bSMP04tBztvN89iTvTIBC5s3JqZqw383UTL4EPvTO3BijBabhx4
dk/0OnyyGx58Fr+fALG63n1eq+BfsCDHCtNjcnVupEgDlWk0Bk2F1o1rDujDYQFx
MBKtetSmfIvw8j/YVuU2gUA1HHj7Rz8sPbuYf1FR9gCkPeOwVUX+4ar5Fq1I3fBm
GwO5FlVEQ36qfe3mMySj8Wue8+8Xe/A5HJZWycX0g/YCpBP/oCKLG+A5LB+PAkfW
NEvVWvlywDAhXEqfy/anAHOGA1fgVGTqTdWIGyVSAzj/4HVoTa3zI2fOx7/q4VTE
1jVP41/B6Z0ui/ax8C3HwIOLZxEYqL31+dGSKhYBYV4WZUFa1OkTQiQcvHFcQV7f
gOkdKfftS9junFFbZYsgP2eWS0aAa2hsupXFsfl4oPOJJOPaol75bMzzcGyWZRRj
WoWQPw2V05pB6KzmyI1cKGWp5kfsxdx1TxrKv17VWz3qvp49od07hrmTbYFsqdSB
+T1eEJjh4KvzUxAC7zAgA/XCKfFRaIOuuI2rlYzO/9Yxi5hjJoyq7c4f6p0r40II
K7DuQfDUjOWq2frmNBQkXw9oAFObWE+e1wT3r/96mP9IK1sLuTPMn68n2cDgodWF
9TT7BjONO06S7WbGVP4EgZUdDPcmevDpaFpV5hnHFJUSfNZ/tRTWcvFOBGtuFFOS
v6fhgPsEMzKu0VuxF3F0ebe+1TWIAv3vnZaDOM4iv+OyYU56dxp8RCJ5cb1ExB/K
oL1+tQmwUT7JNzqS1ENMVNCOm6xs4ujH8wvtA5PuX7xbmqQeVsY5ol3LM5zFcIBC
4TY3mZ3A3EZARN4WmirKwc72iCSxpoleCbc6RHj87GHTF8qgGoMQ8wS3jeUtMaUn
8u3x3KqMb2+ZhYp5Oo6bZ2ghhR0c3MOgsfpKIIrsYAHrcbDpnmafNtdZJmeC2SYm
ayMnnHHT0BleEqCg8JaFN9BQRf9EP62nhI5Szyjb7kedhqm/WRiGHJhleJJ39ZKu
Il1LokCoS9eQwsa+a8eHlwoX5vSHeXJ4w9oK21J23W3udWiNyNZ8FqNgnSl/FrW6
5RWFFt0CJL38cap9zlCjEDTZemcAUFDMT2DpMU9JbhRAdhn6PxFmQ3IJvRYhbBpd
2TDqZnMMNDfeVtV8fIpwrBFuZMK8dpKQ6I+V6ahYwdGz/p6e74x/TFy25Oce2shm
01ofEyAHJ7KpMfj/0J3re4Ko+RG9y0fKZcHeUJYurP2lMH+JqFdiJAxQPYuvEAeX
YLuYwf8uzXzNt/LY23MR0pfr4YfIG9iHhlAJf+jVBLTB0Wo2GUc1A/oEqFfXVpvo
XIpsBlApaAOO7o3BkpEmoU0sJx0nbfzGJLuiR/UuFzmwBR49dnJBRviQrKLJQGtm
eyxpWig+hlSXPfD7rntYT/ZsYCVI76I7dsfXAe+FglOanLImOSaTciTDbvOvKGG5
KTiBonj9pOP90shcWnAMDfDRQCAa9drwzsoRfcpUdkPGg1zPntF5dD92hajNYxnt
4+7OdeyB4YQ7WBk72a8ScNP2jjwTm90k6JPha1k+DvQBXcAy4gtqZdSvfN5G4HJi
YbsG9k5gLzzosnIFPjxE7Zvt51jWzAKInNQmiBp+nVKYLgWabgCeQIK2C59IxiwD
WLm4sK8fDX1aBL3Yw/wRlaUHDTic+6Om8dCbNfIxNy6ARw41yqhMARJZH5m3szzx
uy1OEaS716nKD9Pw+8U1i/c8b29D5biVR2VxpiTiYRnEPg0eINkEF52FJAo/NztS
lL6MJP+L2UsCAGyAJb0q6gHlaG+7a4xj+7dE5DOwQHduRoSd484Z5N4X84e60t8V
B6bRsvdA5xOY3hSBIQqTeZtNSAGNfzYBsPHzeFY/Mgrfb9t2gMyiIAnwTsxOweJQ
WujDUatJPRB+e30si3E1ZUitk3LiZFM8pJT3tYUpoCboQcEfjH92kBZoehmHfvUT
TnjVoasBfLnlk1z4Cc/cgv3oERlWOHHTGqf6hV1hVSNRhhF3+THEtJkO7y3Cssch
suAVixi/YnvCv7JKJXlZebb5/oY8UsHfAvQS5M0qov2K7biKW3o5vRMXdqcjYZnK
42RRcpVqoZuvbWA5teNHP0uwKN+X7+Cx83E7wnQboN6CLbGmPwcfkEI23+tvawyz
tszQwJkPC+PFcGmSnDfMAouQ6DNJhU3AJQcNJR6JoaD/7Vx93LVBPQigqAhauKKK
HbVoqnSpyQZt4qwQqwQfTWRP4Idq+ycUTVZO7faHXaYNUtuD65qf3PwPUZA3P2lG
NqFa7pEfPzq+HBZMP+nlDxgKEnG1a+VFKklZNd0m6F8sop/tuacol6kYK0nMhPaF
yWmJ5v+PCeflpFkHmjwLcuZaGReo6vQTu2yxlr52TZEPRy8H9qnBZQmU2bgpcd7D
p2WFF/iFbyNe/yyqvMNHGWtDpXAYpGa7C5whzZ/CTBKcQ6wb+kx8HOPSSypTT9yp
msmNO4gD7WqKCoW+1IPsBij1k7zi62fvoGho1XXfM3effmx/k1EqucYVmctWxx2Q
cC5vo+wfR7MxCwRbrk7DqWuvv6iVK3Mq/XspGD498Lg+OQsMcp18Te5DOC8+80I4
+o3bJs1ScHOp3iQi9eI6Z/JKBEGs6QkyDFtb7YkvYbWuocXbcCDS6RQexDRZFzyh
qe4unL/yej3IBxkirgEyFRJ71l/aOxgQjq43TxDnTGnmXSZerK45agVZnWZdf+5K
D94r5Wmcba+qHSLLAsFSLp/jGjpv9hns76UG/IqWIcnTQhuBB5Jb1HsMWPMEn6Od
RCPAa0jjiPqiR8Dyl9urEQ92sE1oqszdXhdBZMcxm3X4AS0vgLZ5CvFV91oazTJg
6N4gtr3un3Zw3Vw+Hn4nyxXnzNBKrFZ/JJqvHNH4kNNrnl+QLXiv5Q0Q2ir3Ur8l
ucwgUmOXjoP6LYxSxRfFFo5ulNDp8/PE+Aqb42wmmqwpDABMl5fuP4gujT68cgMB
c/PWbg/QDrGbfphosxIp3gXEuvldSvOkH7yRsJteMdsbxv+ERYf/8m+IpHHKsDqN
s9AFCCXAeYX8eGEwgLtlsEskektNC7yHqjbeMp/cCfjkMRvpqKHdK/yQJ3NToRAn
e69GfAJUh7Z8Bc24uiZ3fOkldOKJFul46tH9Ohd2hZv/gFG6iDxcXMj9JNWnL6SV
QW+Lpz963WBDRqoGQ5WWiKe7DCn/U7F3Z7xbSUmjro3r9I0cAPVKaK1Tfx5kG5yI
BMj1keaubQ0jxsGTzVefa79kjdiqPmVQ8EDerIAKB1L5CcdAfrQYodFIT8T2TPLP
IRNKjPWWNXeHVils4tOf+ETyeZYcbJswvFTQGRLA0rc3w4vfXds6KrfjGXm6p6vp
EM8LDeYwF/jQyTATmqKaRkOHsmdf5Dk6WrLR9Pecu0PUHAKpkuUZNlQT6j25RrE1
PE+CFYw5i9FexZbP5QC8mTHYwc5IRBLNqPW/32NdfSOBh9oDsYETuLd7qmFyvctC
r4IjR7ueRFydP+5s62AwiZouTqMMlWQWFRie0xkqKm7xpO05BMY4Pb5msNnhIE7O
7pxUZwTblj3VbMG5N1ierhXfIINC+6H6MDUfop58ccYGQcWQBsUEl3XS+EpY4IGD
XZGVU2ypeFN7/JTMORXPDz5xCUuoStlFLz5RClEJsK4k/MZ3yU7VWjYGIh0poAKg
gxLnO8wAPzCNqtH3E3t7uiC1om/wNAms8aTGDQ65z87FtfGIAe5/qnf/VPjRBSam
4Nfw77MOy/rUbiwDHdR43pXojWumcq2TktOrA2afTeCvWwAsjhfOLEu5uO4ebCkU
woc+qQuEBbl1vMBu9Pp1iVYqj/NeQUIOMhWe+0ZzS0KLm5sgwTkAlv/LJPtI9ZpT
hlLXVpCa6sgFOVtcR4cc25qCwk1QSi7tR4x93MQjtaJaxEoS2yZs5ap79NkUBmEg
cSTKOMAfm48WhtcVdJzTOBkMwWQLbZycSiFmklktK2I8YFPefFPtr+ewU5JU351Y
mRacLV1dX4ms5GwFbve/K2YiIBVml9zFbcV/iLG3l7h/WZonhARRuO2H/CdVHdoH
E7T6qyHcWRh3J2FRLDdPGALbZV/7aUc56PrHMVzToY3M72ybaCZLSWeINRisHNuI
yQXd0fWK3mj3L95l/8PvsV9IMttDR0UumkjAPb0o6XY1SqfQcbgUzb8KoPIXYv3G
EsFG1WYsR0YxE0s+zzxkPxC8gNOOfR9nehPZdf1g1qoyA4fvPJoaeXo0i3Zxl82j
r6W2GQ32MlAPJz5x8uu5IclW5H0h4RSoaNz5LioahMBNkNXdizp5JL9igpb6j06Z
qyN7pGyzAKPHrXkgtyhGxeozhOKqywPdNTVb02wSb1qcxdTjgmBp/AecJqVS+UxJ
RvSZl0rTVMMHks0AOaICyWX5tII+QlNT+cWgFmi2QoS+4dbkciu7PLC1uQucsneN
QBDIs17ec8QX5AEqqXtsHmkrgdHhniQPcfiqQu2Uc6LhPStyDSRZq0EQJbmnLAgP
kzcFH/PLodBfJ+js49hVCpwgSMxnlSp3oF5elfBGV2r0Idv87DyiP9mGnqWqDFSo
09AlIrqGRu2CyWhw96KnbnywxpZHdGnm9iPk3LDMkigkHQs6eT1k6mWRiBFz0SQ5
vgHChQ0pTOyY0AQRmRG98bYvWXMbT0kiq2DcUPqUCNKFypgLcQzOVzZb6S+/wmpx
JgaFYxMclem7zUbFjENE9q2aTM9emi8cQ2mqDYmpLzC5wa8Q+fskvqcBNYMGghuO
MaU1qZq1tS6lLj/MkE9FE9L3fo4XHGCtf4EwdEdUk2VvmPig4K9D7+3D+rtmMgE/
9zhi/xhbfk13N0aw5E8BAX654bd+1C8KbtyfLyq3ohn3Oin1dEaTHloi8HKkpvR0
q4madoz4FmoTocTG/Hb8qvFjdF5a360w67NlJC9AqO6QKMGGhAcg8Rlbi8hqqG36
smu3oq9kBy3pCx7DsIJrlA3rtaYva9gTMNTSqU5Ub5PC+4U8gvroQg5Je0Uau8r+
iNaf8jnomowvL6CUkxfoa8H9jfHmmvpMe79egnRoqWmJgZbrli2SAiOi0aVN6iSR
YvcH3fdqtmWjhwVsxqAs1nexKUaVUOhnQzniAOU1deS7QfQOE6M4BXsQsAKMOTGz
vdppY2PVkE+4xa3t+EU9oBuUOin0K+JjHU0O306FUhGL+A7+8Obe3+VhRIgHz/m0
IN0r/i9M+Y5Rx46oCc2tCKFaS84R9Wnvu8lCYklUAzLC2uC/ZY8RCmDeU4jazEVv
10f5QjA+7/P7teFeow9d0rd/e4rITrOuMpdc7TbIi22xnHX0JQWW4vQdZBP7NYBr
bwsmm33QY1W859WbPJ9yC92RhNekW4bq1VemeExULQk6T9yWtpU2+IqsOD3eINj/
O9xjaFs8/xvUvN0/fVLekTx+XTjzkbR7G2w4N2GJQIwRR8utt9ITyBZJL6Tdnjky
R6qQDK+VysUsIOF1y43dYAgscg1Cfee6EQ+QpO6ZJL1fPAiO99uujm1tBzSajMSV
CbtVhfQsrhEUDSHQbUTNo9BQKJSnVlnMKtYMATBd0+j6zeFY0MxrA3p6kMHYYjz0
jLbSJuUFBjaDAWIpqkyyv3DsOIPuICXX0SXqjZJbnpqvxpAmxDJupAZcEdQeVh66
WEASefNjZ4XfYNyvc7C/Gt8ugmsXkCsK9j67BPsCsXmocSwXdxkWvo4ajXJcCWC7
ndtqS+AkIduq2d28e6ktpIHaVW6NkbgBaDGkoBJDvhd4BWzeU6LYHgNhLkgFWPBF
mlwZ5yCuIa0RIHu1u3f42ipa0lkdgCBdo8E9hFkyUT1aIZOXoa+lV7jkKx4t/9OD
AQP6mL+kmPvxAJAp4BrCbfCfmuybdQkln4yHDLHxh30Aeab6DfYkM93nFItJOQwZ
hVCbe+Qsk+EIienek3qHdxPqfCTdEoVyIhHwCLI3i1ESSDX1CNdvKpNpia+gQA9x
b75ueamQV/EDkvwztcGsMbmlKMkmEPr9wibx+E3gZROheLgxjkzVUECFaUzqbLGN
LKgYxuAmXzGdPoF4/fE0OO6t5tyjwmUktzkUrctHvzpoN8lSk7fLPKZgRuy0ZKYR
MteD7cGI8q18OUEIm9LuTazx6Kf3pq+x4jbvsEEOdMH/QTiyY0Jq/ljf0M44oYni
7bsVcpzmXnfha5M2NxqZu03SkR8mmP41zq3n2IpgftopCVhcS0pyXJcPMTLIi2yV
ZZ+rdgZBTsp2XAozuCbzY+HS76B4s6n6kQh42TuGW4MPUrj7V289uqv16sU6ppPd
VO4icjUcLlTutewJCrtAmTkluLc9/86aUbEY9QjU/jxuWXWGcqkVgowldavCPWqf
mgeAD+dYX84+AlA8MZxLt9JVFEWZOzFYFUhhqB3nHhAvcUCyy753F5rxPMgd7J3T
vT37kFINXimzUeXs3Y/Q+fIMGK20y3NOZzMtuuP6iU+3aGFJzI3JNzQhmu/CmidY
mYFrscefTskU9QuqODBHwXc6f+p1FdNUno/faeJBfZjjpcdoh9wzFenTTUrsrUDE
XNRYi/6sE0HfzDxpul6vEZW0dbITK54AWG2vjNeP+skpgIQpr1x3fvgdErKubarl
tOV7tDIsMaT4TjGfsjaqrNc1j75EzbqDIY3Tckt+3/PT1pNuwNXwTWXolyjA5Xs4
3LJG7BRgKFDaPt9C8HZhFgEkLQyB0kt9wUzG+SNstSagqC76PLnA+Eh6lIO1vQBe
LSQeo2R/Cc4SOmi4sO6xEqRJefGeVaCg1adzEn0d6UKCnOqAeUrI1FOXRwWWwTbk
FHwKj/7/mbp10eOIk4Q9zFSgNKX+YrIFvhUwvlIap1oeNP9BcYdy50pYfWK+TLu0
0ZGKfaXYa9tpJl2df/yf1rcaB2HyiWMtFdf71KiuOUsw1DBewFHh6E0/DV6sSPG2
wTLDGKDwl9Vn2w7iOVuINenQ7oPXTRPLQck8l3PmB39uEDb3723EvHhK6FBKy82G
y0dIo8qUEj/cZJbcAfOiP1iW08e9abkEFUOkWjPgWLmzBR7+OBEtTafcRpywsdFa
y7Q2fq+vVp8iwfpIPfGRu2iOP0jBgBKluGJQjvA/ymkh0JNeV9CbxKXchuGTgubR
4896F5aCUN1vXhVpAbAMx8SM1fxA8TXk8GkYg4FcPCiopm0T1c+z+M5keXT1JhSG
xRAaJpYuxtN9+cTXNcdV1eHILkpYEzTKJ+Qfab/s/d4Z376AD5l+ynfkKwnvOu0p
zxZtXmFBLXlHPmH4kLelaubVZPgb2hus1woC1BsSvOsbnTfJvM5W1oEf43rAlwrl
0G1AdqJxyfHM6EYApVZ2tjb7vkI+DoCnmipK43vMrOV7eNwrpZnSEOVkzsjcnBfc
Ajt/001C+EtLsfS7cAy6dVOy60K9hdXgH3U+GbhbO2EDF5brW8/OemYxr0SxDayl
kdA6KQvIIQOibO/72uEJqdZu6FDJVnbcbQ2gxBVPqbhQPP7QoqhwU9cFGINsgYdl
oozc9CR2wbQ0xhRLVvOsuyjNX7vhcYNhk3WIMAhSsjE1v61DNeVbfoi2DdU761JS
KPKy3//k9nR3H1CTJ+E4cb7tsCEnXjzfHwidtI48Rr2cW3Uh8fr40yDwvmZKH8uc
1HyDXayxV3iXqNX2pgYHA2ipmOsG3/riPIbUxUxXx4poyncOPnGVLTDkL11HGXBl
vUwJHY/Egz33ZqJx8WwJF+leoBZd/EziD/haPFoP2H5L2n/nJoZ9GEq7yUeJnSzf
3LM4PMkYsNQhIImdoYtGLQA010pYxe/VkVi3HLX/pLYlFManiWal0Ufr6TDVkxhO
YxaH+20BPqJiXnaSXKq8KxHXDv2qGwScJVcyrrrkyr3OxO1ekoFLVusSVUzteusB
1Qz69y+27ck9hwUlNrAM+ea9xrc76fKUKHzhAY+xS0e8SsA++SLdquVj051WxxL1
PAZDob+/Ro9kXwu98xNSiIwPnupJo15MBjM26TMBuSY5DTjL5leUhtnT7Dg7ksad
2zX9Hd/pWJaQDa7ULTtH3q7ArvOf7N43KbYR5nlM8jPJAuUaIniHguMYL6U3Bbfc
XH3mFiI516Q2+4n2ElPLccDZMxJMN/a/eUzqDFhdWBUtpHVwEM3A49O3WkmY/nqN
jpgeMtb1vO2aQ7dsOaGwqOAgMsvbnuMdkbNjC88TEbIykBTndHo3k194xH3bU3Cw
8olkSMB7vD92lo0b7uBO6klWOKWN0/5zrgJGGWhDs1c0z+cDuzdtVcJ0Tcg2frQv
at/8cmx90hrl2zZ1dNan+CfQBErjwQwPjwOleRct4WLqL7UKK8J5wOPw+P15BWLY
g2MkIqDBZfPzn0/f+If6mDhafXVxx+4KKn+8cW9soNxe6Nr7Ngy/3xLnR7sCMT7a
uMqKhASQrU08b0KYsgJfD+5IP4ssKmejd+6MUxMIX9zWdrAFqPy7lskd31Nh4M9p
ED/3gsgpixucSKs87NA91WA2TqAPwN//yji/4m6Yf6tAg1zSHEt69lfbqNsQkNyb
Z1VAHekMSIdRkcZ072soeS14Nu99AM7L4Nlm3/8hOHRVPU1RhVKCQSwIMLLYqR+7
R3rKDI9PsL82KUtqjplbnfg/i0C8wp6+akXvqxHIdUbEob42n1VI9/D3mVnTuIP0
YVhELRCSlNY1N+vFErwKsWemFt6who8efI2bthsSqTTiKlWQJ73KJfG24D+xzqvu
NMNGwGF7XIddohU8447TzS1y3bpfEb2JzHB7bVUxU1dgL2l4c+oan8uzIHvv1JRk
5O9yQ07FGxb6iW3iZ8My6mNJQGtzrypvCt8zZxxutGRkqO4afdR+nheIvSUoE26A
LdoW7mU06dY41uBXXSS4NfY4h4R1DB2tZDo9gs8LSitHdJ18Y66xQEEyC6ye85Vd
HgStkdt3zAlG2fFi4pn3Az3EhYdhhF1Mtt6A9BHIXh3HNZzjsDmki1bK3odT3Qne
BR7H1gfhUmlSJB+etZD+ZGacA0rlnJmUjhVYwWWn0lTnn6vxfAq7joX8j9iQPOaI
p4dD4ynXBz2WEN28/5QNgY8cup2LzHza3tuEcLisYa9+OjVV1zFQKej6Nubvv5cc
ITrIftw0xAlE8Rgm4Gc4wfI8Fvon/xnRpyz+hZMDmvlUA86o2+Sa893ImjswG7b4
62MxQuYPKQGMJvjWpP+CgbtIrykCmYuETBdWUpvZCCVppNCGBiEWQZmOS9e4JhrT
5VTnF8fCGZMnQe4aR1ZVql6m5d/rNCZ0/+GXutHtERA0xec6EOPkel9vKJ1F65vn
69syu40I83YqssAddO0AWqXEbP7YArBZhzMAnXfaMf7vWZAXwbe/FuLbEkZGZA/w
AJriRWBQ9OmocGzYZBAwF29BGJ+ecs71d/KxruszQkcDq7jF8VcvFnXQGzixPqMr
WyXQDs444fs5mgl0xP9x35nYapU3xsOE3BrFd5O6XQYeiZxPAd7SX2Shi31HvGIx
BzBqA1VkV65F0TdR5apjEEq2uO78gI7g9rLB65rdD+HCAleN1a42k1RQRhpw/5Bi
jI7R11xttTqola7MbVW5lXEm7qPJhPNASkqPrC+aoHRgJQ5fYZpLDUhPv685CR7r
tB4LhQWZuxZdWwGi+ArJdbZuG1WrGVfS6QCOFVp235HDPRTvXU7TpExtIeTbEsMN
tiy6/3VPi14X2Piz5M1Tvzh7PJO/K4Exj42h586bACy09iLwTQdx1d5pa1D0xvVE
Qmj0KZd/OgFAM3miGh1Exnx2WKHyehlA8e764noOhNVnggRdGDcq6pH2X4ligMz2
Ef0B1SforEA5fX78P4oiWUOnjma0gpzwbM66gxQQPe0JUuglBvrWPDYHLsEZclsc
IU7UvtCoQxanYEiVR/2AN/vmoC5R6F3AF6lt/M8Bpw2ax93dUlHp1YGQEHMu9yrl
n4A7alFrVgatKORkqPrPEM76vWdna/TIK0g2Y9DfUSfxTvJSqQ/SldeKpmU592Ly
hAIm0i5UsGCkFB/fsT/3KxFAwzNgUEdb0eyw0zgQfY7RcK4F7tdwUyvcOmBt8HaF
omaMS1UQRA2cFzEEKYLz70vywYqgxMqtDJBLni6UH39+kP3SDFFLH7Pz8QyIXYXn
ypVDD2eLAKDMPKqb44CVevvuOZw94+RK7RpvaNjvOzSFCaACgN4nfhj2RiPK6gVG
aYBpOXICBTGLm6UHFNqi865Xm2rUpsAstktBjDoT0Wpddbb6i0VuC6FdTscdBUlB
7mxeA8DxcFYZzunsf1DJu7CV3pQ71IxduX0+KijfQGLRQp8G8Kumq0gMYfzcCkWQ
ROwtJrZAl+p4DkCKQp7EupeytwiBa4fQ/t4ezd+L6D3xY4zjIylxfebM92/KJkRi
Sl9NYaxrM2OQjoV/L8T4l6bjrZjVTjVamtSGVlBug6kIyL8ioZ2xzLBCZggn3ubD
MJKyemjTLqu7vhIxcSKEAjBLvROh6TZJ1ltBkyucnG7Au7MMak99TB5ixwigXuNZ
FFeRJLNC/Gzm6yWr3B9jZW+NX8TylbM23Ic3cL4Fl+hgmC/R0psTSsg87cDObPAD
Ac74091KYOgoV4vd8pIwYZUILokNKLvRrzfy8cQg7RBTPWltPcN5kIhMgPqzmfk4
aN0JdiZZTey0cJPkrcLAKLLtPUcS+h5Fr0on2OVEWgFzA+Q9LLPlkk/6Jaq0OrVh
RDldWVvb6Byjsy4lJP0h0gzUxJa3jwtS0Dn89rZAfASWymjz0nRrl+bJuOOdgQU4
JxpT6GArh6rq0/sdSM5TemgDz1w0rE9qWqAuLx9HjwNxSuStqoZJnKmzlt6jevA1
bfV6vuGdxrvNFDF4+APkN63erPls9K4pO25ZGjKxciPT4b3CFcQuie0w42XIGwKc
WA6cy4fTgZZ3McoUlxwxPOepQAMA6+6BvQgkLhweX12ZnqTEphcHoKxixQXqj7uz
UCnOJiMiNL+M7uzrGC7EUSUNPZR27NXlzR8SIiH/s6168+LhjwhVGn7BzXYwZP96
y2LjyDOHJqAxYQXYUZemjI4hD8EBPA3Yv9ZNIwAHNMw1THeSuyGRYrXacgms2u7Y
F0QSELr+G4fRqH9EXyyRePPjx814/2EQLHlBs5HEvN45paeOJXV8Qe/JkT3RZsPV
oZiwS9EbWoJQk0sqjQnwAxjnTRoe0DgB4QW2a8e9WtMk9FQkqHnEIQBUjn5FazT7
OUo7e5vyOQ9BOIOelyG+YHpSOZOS9TsXe3Huzd5KgDD+yf+/uycGm12PIKiGQTQI
OZU0PnkDd68wM9qwuO0MYCfwSqfc97Ms35bfEf192/WZAOFJC1G2ZczEJBAPhr5o
uWFBoNYv61m1+lXdvM/DD8pm0d/HJFn/bbTF0aWLsBm0nBneOJsT+N8yiOMn/Tmb
Oia77VZad6yEU1S+7OD2u3qZ0MomnQHObpHbohYyBwnq9HRjekUd/lD4mAPiln9k
EyYH+bInar7lpbSRpCuVrDpFIhE0sqVR7TcsGSJDIa/mx2CvBu07oep31ZrMT3GD
kM6QUa+mgIYPT/la3I1cg7cjXPKjof5OtJzcPEtm7Si00+U/FRi8RispwvZ979hM
YheJtPeG0ICUc7lqxHWrk9PNDOVafEVaiK371PGczWlSV35QbwZshhikmo4Q8p/i
nFdYpAszno21CZTgoNWBTkIwsh1/bVNmXN/G/iFkjuxNpT5dSgEBehEtCHnIEKLs
bnvd23aYfafsWbfQ6bD7/8eFi6/Ga3wXzg9xkBnEH9CZwY+kcOmke4PP3m+E1Vlg
FY224p50IHo+uetLsV3Kgs3l1MOkF3SVy38ogmiFxRWAxG0kTpzVLyZSAtgIDr4E
0G881g9YPWwa8qXK65q8xPgxx7IovudyfgLdhMiFru1zK9XcxUGsISUgSAT4c7Pc
don/oHUo7g1rXbVjVnbc54i2ZvMQgIZgTgk2X8BFirGM1Jgj8vD2UrQ6onOGvbKg
7bXoyw+3jGshj8XQ2m08MySg+iSJ/rZAPp3BR4l1mjzShHkzobzt+V2iBi5qduLK
JQeeREs9DXzg3i0ofXVANTbOH5L/gFMBqsWQ27yOm51hhYfwwHaMGFjVNgM7Xo/h
zUXCOOPSABk4363uDWyWsr2IGBynlCibY3VUAYE5IeIa5BlZ4OMk5B+9v9r8OtKq
IFTn2agC3EUW+zYvN4JEt7J/X2nEDSdrzWRFDafMZlRZ6LqbmbByodQr5rcXNOT6
dT87EnrAkkokfWqfxLpezi6HDWHj8yDYAgRTJSMn+Jk545n92z8Bm4S/gUPl0l7l
uj0ffuo1LHrimjt8xN4Uf8uECmASDu2qUZN3Gb8puXBtHJXcU37VpmYtQSJ+q+4N
xObXc80APB9qmgpSqgKI0GOwlZL2SRm0WreZ+/9ZZ19/B1sP+Gd+hv7tYeRlrFRA
zmMh/mMPJrjb8clJQWM99tRbmT04LAptZNK1/DKiqpAV1B8Cma0MXv1TIsH05A2a
QCw+oGnvdlYRtzUHNLik/AkzcCuYOSR5WsYh8CTdPK0gWEs1WzjNi+3moejZ3u3w
FFB0pDAF/H+lQhK8R3Afa77BNdj50DNKCtcXEgFOQS4LH54Ve4Ju4ArNm2ZbSU8T
l/7PZ0KvGlJI4cjLy7U3AR7edP/usf7mTKidHzllZqkccWXdgkAc5HyYo0ChcIiY
fgb7je/83ZuWaXNDVXBqO9QDSwLmjTMdt5kwrsd5fNHXRofk3al6UnVObY3qRFGu
YJAdxJrlfLT5/TW0zvUHVAzvMkeFyvXvbLH08wfOpo5VQHNDt18hlYXIR4NbNcwB
VI2SRgvVvVl38qHY2HuAjoFXNXOovR31z7owXqAL7xoa76IfDS52aWTo/nXKOj0P
NyysR2fdEwDYhfCHUg/JegtQ9aEsnYoOJiZBX6ydOj4ZmcBqJKPtZw0G45eNR3eD
m2sVzWQU0pzbd0R2Tu2sTakvVfy5gj1Ipf1aQHi9CtTeA0EW9JEEsBpi1ApiGgM1
KRena9jyNl+xIH7u2SJDdA2NLk7cQx+xWul9hIDNouTJu6l3RNtgQJRd6TQ29uSr
i8ofsiYqc3Oyj8tMYtj8kcJRjqzrobKZBAZmvBAYO56/KDRXDSa2VulxOrOLOhkb
wQNVhAZNwCTC/jWrBzflYsH1Pf3+j2IaNLW2KitpBTBRKpxqTsAwoZsoLlpnRgLJ
11xjle6uPFuR6GuURGFPCuNnbsV9H6I5bEmqLSWKWqYbycOa9T0S7Ij5AsHclNFZ
tDg7OAswCCrM6kbOgd4qd7eTI02WIllKOjV+cQipkamSf0VLz5xfSfHt7dsnseLq
TphPZJTYDRMWtY0NgeMWfRDQSWZC6GW2Xpuz9DnU6ObMdQBkJ/CscWBmyH8rOYSC
OzGsyvhD8T6I7T+Og/JWwZjPABw1IgIO4ACC9ihTmAIZ8uCvAoHPOvBuVRVJgzd6
3lPpO1z4sXIWAQitVMEZtt1e8Awy/mHH+la43lo0u2CJ/uk7iiSfvby+LiNRbY5F
iSq9Yajn6GCy7JHp7aFgRpApCxY1sZJ/QMoKkiLqtwtuJP0nhnQJAZcKKwGhw2kt
qnClEPit05/i6juIXlTE1kY3qjqGDBm/Ce0S75nTypskjqi6dbFjt92HP8ZVadmN
mDMzbR0gwIQxt7G1+sdrPyqWUG5TZtRMeVSU05gSmE9cZSp/bJoc+yDUGKRmi9F5
P1jQ2RGaxrZlvZKnOkrqbd35s4PlP/ANpvjeuV+5ae5A9cNrXR9EKAC0jX3Awnnm
2oSZZODsNqW0swoPSBleQZ8GbmABc531535NCysOOYVVFGMCvHgnrgTTqkpTKNdh
flFV0iszy5Ha2qZHkVatHul7uhwZf0Uj+0k7Cs0Jxt/fdo3Chervq24aKsc00sQH
qytl2QUIFvnFUw22PDrEHGCz5hrGtZ5z3/XeZAIZ35Kkp3buMbUo+NPCR+fNfaWt
WSla0nMvkVTwSP3vlS1qyXUJLINjqPP2xLRoVry1NBriYXflP6y6qCAriNqh0a8K
uuTKaNNZq2I/ws3Kkn47ssoaVFMEfD1L2UZnfMgAbUbZlWDDGRwplTl3tzVa/FsC
6zM//UTYred8F+xNmN6wtbKy8NpCynOCqmSnN3YX6GlezsgdwGOO4u38VdPT9o1k
3mtiPCINcKfiengWOfUF6Szr9aNltk0d6RxamuVPFqG3RvuvhO3wj1ata8jL7rQF
6mc96h+spHcxGtVzLIQX7bwuADTnZixQGMlA+sXyQEHswULep0nJ+HehwLE7bKD3
TBL5+Eb+usp9T8VcsIprQUL9ODJLF1F7vYUFntluaIHiHjOZKOga+YkO+uLk91d9
8mA6yPXaxvUvViRdo/d/PUYiUDqD+yO85MZbxwXViXJFX6ymGRQWFPttPigOrDcD
WBVkMQzOntarefRQE7Px3Fs02aPd0jXMKsyalGgoyw6beLdQDaaBU6TRxxgkqK2M
L76W9iucTd3aeQtIE41YR60FVuQXIGHu8e+ld/dr11kVxV8d0c+z0GcqTGV62Fy7
As4pm+5CYSmTdiuB63SDWqMWdOryxFqVmsrk9QyGfCVItLp/wNPE4scHpnyBekFI
1nV/VmP63mKRDZFlwME37WLdpFtOb66Z6H35tvOppfOX/oC/6XCiBleZgH4lk1nt
xb9NxD8PaZSbGFPz+n6WH0iggVZ3D5L8dxIQjwaejZwx2D5eSx8l43Bg2ToF7COd
cISE2mlTFKNgZXGO+lai914fIKLa27Y7ud6aJxljL00uG8TRvzOIj1pwPqPgcrwk
jD5lxJRH2eppXLOU1p/2JBlHx5YXnCgvJOxlA5EzsGocQyLL3MsK+/D08fhGg1iW
ncHDM5V1iRmoZy5Xbb2cuGZhfWtUMjqs6oe6Hg3fBYcs1Qk7Zl9b9qQ6dChMu1Oc
6ewYrJSrZNfZJRW8CMXgZQqPbNuh7HcEpW7pjpRZhf5Pc3xPR4KH8fKB2+HVLyqh
cvCwn/z6CuYSo83TFQ3MfcUomB31O2PPfTo5pLpxRW6Zbyz6MAXD32mj9tTv7Bzt
dWY/oR7wBv5JLU3KJHq7/ALRSlgup+nNoMEETEarOaVWgvAILwjrS9WM0EQeRd3K
3ykD7YGjoYKKLO0Vc2kNTd5NXi4g5D2qqioUdyxYx+URYA5QWd/2K3vfxdE6kiTM
VhKq2fI8FI4cf9ihCilKz797F/6jj2/aYYGr20+K2uOFiRIdoSp73d3Jt+Db0/11
p9fgxkRpgE7hCQw5M9qpaEe4Mtws1VG/BJduE8qF3g6FDZ74JlLBeg127JUMmxBW
nUQCfPR+qYrgDBhCpbC3qzWDGDQrbqBCnFXLrHDgTH+DNVEnT0m/BkTvRGcV8aeq
w/PO1svEJZs777vxDqYCgDhsavozzHM+Bw4ztm+5MDMhM7NJy+2I8bHhdIm5LZK6
HDkO4WhaeQy2ARLWGpdMYDZlMjKpcSa1cYDahmdJlxf2thwPliXAnCrjkqKmTlQm
MjeMUGEBV4euOcw+q/VDA7XnfI56PKG8vZ5CQdmf3Xn0aj8luU1kxlGkUc7s4EGh
duNTVEfxDQ4FNawN5A2dXH7y/Nm7ZpVRMKQ7gZFOm7JjOeEjLEFVkkWMdFnpgcFb
Vwm9e0I9n/qLKJCMETOA33GrfJo+hFLvaIeeQKAV18annTCyObKbVDJj/79G7I4S
LdT0Ao8YZvSaL9Rjwc7h7+AJqtafNaS/0+yXgT5guBup347iD5spi0VZYG+302Yu
P7cTOd6DYycxxCGZn2VA+LfTKoowlEyl4xGObwRvJ/uWTEgmIMD/Ze4e9nqVkVpG
cZiG4iZMHoR0gvp0xcaCuPYvtSouDVnDNMlvoi7M/cTh1q6o0t4hLIqSnMr+Wnz4
eMoRldp6b1PgH2Cpy3im31MYfGLjwzmWtwWdSV6H8qOq1jl45zJWSwJiXsupW8eN
PYTdwY+fAE8a+Ter+vD3LfDBHTjPBcHF9JjwHk7+wjdUsYLaiJE78U8iqBkyncay
yS27z0qIlq++RuXg1NhFRzmzM6r886jNcF4lSh8e3Eh209RVYKsi+N+rSMng+2hp
Sr05mwvG88BjYqyiBvocvsqfHit+DBdbb1ngvsOy4JEMy9izzdPy4oAnluRxuxKk
eay2xgnXZ1kuBG19Ai+gAjn/wB+PVyZ4HDSXbPruIkyTqQ5YzZGUQijQOeDD/GLp
NVKuhskO4PfWvooi7jgFOl6ya/2sMAzAzzQ5A9DZR09f/RChvGohSdVNqNasv9T4
aeTUxk+hWrYTGjU290jlz95GV3Nm6/0zxTpIaPdrHqdtLGDae+7UbGR9mpQ5S3Mo
tZ6hxIIWY+VUG02rCf76H5iezAS2MobyauC2wsIZV2AB24W4yPc0TAkCKQPfULeq
WvZN60PI2yarb7rHH1/4/ziOdzOUSNezuiMC/j3lz2WBrP3Dm15tQAQvF36EBRtx
xJLQeAgc5AiNl4F4K0x5SnsyWtgSG4srsm0Viw63xBJwXCkqC3Npf+6s8nZw5Fac
s1aNTQX8WpI6/mhyiDYmlcptQ4gYC4lOzesUhaPkqiE+mmfHz/EWi03o4FHbeM+d
VhdlP22k87hGKWPT7D2rSaUWtvRqePFDVZVdaHK++iJT7d4ADpSjSYjtBjYYK40J
zt0c3n2N4DJcMiak0+U9c/2Xuk/1XbyAAxAan53oV7bjoArqhQUElMVwWR/D0jPq
B9nKwTotfk3Jv7pBF2VXW/vhLi+3FE+IgAQ+TCWRBKlr9/gCgz8gzM1BG+NSmYLr
gyWSapvDv0jF6zTyfyT/uXu4Ezkg0duDEo3tC3dRAyVrKWzlBy86ZJNICRbiUohn
0FPHC6A50dJT03hc5ta56v3Scq4TVXPk6aE6oBfrwr/R9+YpHkeKHLivvZhXWq3O
axqJK4+KoInkWqlByBsScvVpe+dpgZQpVGlbgpcqo0Zwt1nIYanzxmBkjC826cpt
lEX8FP5Xq5Ub5D5kXjdLLvDwu7/lFsKlnuwyDtiMd/ZX1Bj3PmoJP1Y/PMJPz+vV
KLfcKyHyxcVE4udes8X0DWSj+uHeYd8+LZZL6VLalY+FjiLeF7Wd6GSsqu67iXeE
zz35uY9o4yE8fJQA+MAfDZ3wycip2hwS5lqkrsvZ3DAVfr/1GoXdlmvy/3tdmhSn
RwYCEHKEa14bOV3jjKSJLjWnKki9x25wgUGgs6O/CsZVHUHm20vXG3WNmRzr0MEx
sp7JDrbwD2FSPofUmQ/D7FQMv017ZexpfdACMa07wS9YAbFxct7R4tGtgRqCNdUf
D9fxeNHnRRL2voLutB9eBiF9sf5W5u6iIaiSsVZc+ZyPXuJWnUemkkJrVgrOZ1yy
3lnyy9PdBeevns6VVM0fScv4qLuDddqbRo8p4BjmbQeh2gTwReFlXCmk+IvNL0k1
S4KNX8Y6lPFWSGb9rTZx/kleG2sG6LLMGZiHUSSp5eW4i5PsZEEoYmxoq7lLslDc
mQ3imeal2bPWekMCfRLXEXzJaTCYclk2F6ugUvpvjQxAf3vWsJjGHcgWWusz1GPo
eOEQQe+Qu0wnC2HKDyZtNs7uugRd2tcS1QzC0C3w+Znr5FSLjcJ3sMKOOvr6e112
pemyZpvxJ0NcV9eABYo0j7d+thNi8NvQLhZE/NVR3Gbz70IAGx1lUCWdh0BtLKwi
BbfuqnkgLCMX5eAMqWYIGejvt1wcOUzotNYaflHgAIXe/F2KXZGN+r/3hxZEzOs2
RcAZ362NE6lWdYCoOOAq4N/+7yd1LGa+YHcazno+wlwbnAn/QVYSNXyCWcBh6246
vJjH5Xaa5PgpZ+JTi3BnZGmLve6mPW3uz0gxvohKM03WBJCXwuDxgR1iAiDoyMke
Q/e1ZZyIjbx2mcQPUvy3XSKdR5oZpOjJRAdjwpLXw3yeuNJPNujc09VgNlSKnvV2
CL6WpOHKqRtQ2k5fg0jNRQ==
`pragma protect end_protected
