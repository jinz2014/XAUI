// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MtymYyBTnkE5/UOvmHXUiwgaY8+3Ll9YuvLxKyU/wWrYkfjyN+52VrjOiQElcALG
dYt1wx4uywYWjkPIpeTtvFOpk1lQ5ULLfJCkwewm/i3rIoDi4YWDbcE8Qo+Bqf74
fQRMBF8YrKarnE6DAT6IrdzAY8s3ifZgFEH1+rVa/aE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1856)
1wXhlXlsZsKdcmUO2gb3so7K9BMWV4rnSwMIXFOcA6JxW40Cm6uEdv0PqauAnTfE
WDkj/rtsYd7f1nG9Ou3EqUV6Rgw/4CxuuAuCQ8gCvEos1ELh4vKZuialm+MtVUn2
l/AiARc7ph2bS/iKUQ86BX5U8cgE3T48T8VGetNRUVjwkO1kdIuC4OcoZi1joRVv
de3fkt8NE2HQkeHrLxPFuF6QAMu6waWVmdgd7hAp1mAxVYr7Kx9snuG8F77wxTOl
PEQ5GHONU+ikNyaTBAE6dKSOczKXhmBBqmxYMX26IvbS1GqSqLl+PrRaX4uKvFEz
j5jbP2GeYuARPSd7TUsav1PTbhKG32Gh6Q1byOAs8MhJW2Jiaj4yrj6gw/chCTDQ
rx7ou+1VSUKIYmVoH+7gaYjOyQqkQnIv8cS3TkiTWta7gHP/bWtTKHTubo7UF9WJ
siOpSEJu5auuOEQIrjq08i5zBQ1GOaRvZ5waacrPP7GGcZHZ0n0U+qr1Kd0cBl+Y
amJOVqh+NcPZaoBXlaOIltBvg/ezKEaSOKy6d6xHewRX8VeTXeZKjhnpMHvUSpwg
I7FRfVtAd4QhTN1fWCujgktXbbjy1rx92ghlmuQWSltn0qPfxMISQonGPHVcKozO
SIjuoybv7TZQCoymEsOHwbd9HUPp8l2YIgwTsK/garq+lflD/vdJISeycUHXNeBG
gpLBZz0UwXYVmsg9bug/IqgS40ZU0xZqdnkY4i/cVMe32Q4kFquJNtlSadMYnKTe
dklrF0ZIvMGjw9LPp5cvdCk7THPTZPX1E46aAZyJaGHC7S6q8Kv45ccHAhgcSWPh
KwMrSfinpzmV0qEukax7cyr8354lieBzQN+7gszmPLJAIentIB3+mD/RlwjYlzll
jQUeP0BEUPb6A9NNZ4RrC3WCPugliN/TEjCQySrVddAOTHSCYIsxXWw2EKy+2e7f
pWlIn7xlVSI7FMkU4enhYfdM3jsPN/f32GLra1Jf/Nfmg4rAoX74mTkXaGL2VjGk
H5rEf5JJMo4grejC7AfE3+DMg3kgP9oJkAIjvGEOCi7QyiD53mXvPws32fEG/s/+
T5dbj6860eBBFZmrbroK9tcbNGFdV5dF2mvXFraZtQ2eAQqwRTSzv0Tz54YFW6ej
K9+G8ZwR82l/jj3EzbxWqtBZvhgD+zifJSRRX6jo9ZpKzjTnKROnuT3Yk9qHwO1y
fjljiZrBfl3vOQjB/NuNmtVK1f9nnTp1hFGz9p7D+yQOw5FFsArRF+ZtPvIHT5lS
KCLoRlijUKOli6nkYsh8bse8rjV8melJNOBHo01co2+TQVflcPQkTP8RKqdwX7vI
dfBI1xWpmS2+QrCD4JxB+WACIPXUlFTlFS3LptF8xcy5Ws6VYk+8MNOzJ4o0uHqJ
xmIgGZgEwLNcBoHTGruQSHfRimZsPm7jxUmQNMm9JKxSyytSJWwc4TSGJw0KCTPy
7WPOn+WVeIegCafSkuWKOiNGFjxN/WGFBJSKvmbpgGXx92UOblOZ1fp0Rda0vRPB
KAc7QE5Ik7oYyhVztQZYb71+mW60WPJtfMd69DYR5Q1MArA8A6B31J9lH7vGDjAj
Amg4z3SV7H2YI9wJ8NiDeXNyCyLA9Kmpig8MNUlC4bEVg/yaFlr+xDmcoLHZczzN
Z0ZO9cdhKeeBjHCWHF7x0v7EjLXaA67YajXqx4RTpLkb6g3vRNtoudrYV3EJ0abv
sqSH5/L2Sg6xVMTl8hJzTIl2QT0K6+1/fEpVQKnsvZCqztll1CMTvwCgayGtU1Fz
/gQgV414gkQKJ7JJD8dj+hnhchsJZQA8kUFVumQFjqktwPuwtAXsSYd8X/DeOYcm
N02FI/4WCguz4SDOOcHaeikrVAC4QXvMLxRGfQr72x2ugg3FtivQWxGHkGJFb5+C
FEV6UuKFidhPssQppaxyqKIMZuzud/SXwoQ2nXVdg/ESzau1aO1kTvcEeWz31X2j
6v0g9ZRRpJf5uJeB5ermO6e8+sNCC21l5IQUHL4KlvPSi9TYufWessqS5X8DEE+D
bTbXVo2HfPZPtujsGpsafkqpaLGDrYr811F2TNk27eUFXRdp5FFUBfdfRgLyrFri
0FBCa9ge7FqF9TJ6sipGWZYqkDAeo65O5eyXbiyqmNWFKIoxwnJrZOs5EeyzlUgg
zOTQ0Tkr+4W8EmAXII/DLHWfS6+M+wOeTC2FxtvIBasN9/zCHWtD5oYjPerTJCjJ
u06rOzMLnkHcvoNQ2FYMY7LCLYHy+mZxOqJ18D0FzQqMelwplNt7QY8cGmlodXAB
Koit3NArn/ib7Kx4iwsLDFxOl9VxjGsOtI3K24UI5GxSzYJloYit0G4rse636T1C
4Ack5KS/7PPoxQ2V/0iEv6JK2O8QQruA4Igk8hXCBhJbbSZL+4Vt0SqfhJrzI4wQ
6tuRS660yP0KlYM6zkL9lO5GLA0DUjXGfwxMiyThEns=
`pragma protect end_protected
