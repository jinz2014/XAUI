// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BEqUqBCmRB+7+NJzuGEoZtUA0XVvhsljEJqR4c94tjqqHfgrhs4V6hcl/TQliok2
pEaxZ+3OxLEwVkjwtLbRbRTHgNcyqjb4wjDV8qvCqDJoYdyC8VoBPkwaNHASZx5+
QpO/RRnTDXDkTQotVXXt7zXdvu+RKzeTVyK3j5/15EA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 45328)
AR3hGednJMWBSmSph/INrI50mPbrzZC7lqzgH4wcIV0WOvqbzuZRzwVweDbe+KDX
5OlqQ3nHRJieZ5JBBHHHWi0ot++diyvpCqAuO95r+XrKpXP7XKLoZBe+DL+sUPw+
h2aXcmIxc7A/TW0s7KO3j4sfWRMKxAlcrZRXkhjbmaIuViIs59kyQr+dana+44Dy
8MeTZnDZtmwWwmxEBYIjPnesqDTWvhgeNov4FUY09NKoJnvy+2fvftuxxDzfwVb1
4IVyPujmvyKXJB+xy7XxE5IQY+9+vEUaae/KTog3OCrsW+uNUWVyDqoL4/gFvGCg
yGwgQP7tqfdo2KOezk3eyXD1BYAs17SOfNPgddGmNU+iesw18erCYz5Dc2OVxSwm
fXCv6oExHQg816cjPjjp8S/J2A/PJ3T7Pd+HDxqB0tAFqcE+6WxELlWPseyt1LVZ
iAEG8Z/I4mQyBj0ag/gSszdlQSgGEl3srLYbuyPCAN6ikjgoPJOh8fujubp7HV1w
DsY9phwkRqFWJgYxHdkrPjBf/JNec2gITMt8nyEAtddQ8E9VLUEq4grNl/UZs1j3
LiR7uDTmC48+mQkQIILRr1y+rtfxbaOI9ZGQBhQsyA6adJt89nA2IMNeaOg0fHv2
/QwlTZuZ4snxYaEmJ5jnfmG0HBhKIFrf4gT58id16IJDWXjhUHsqIfQ1BElhIBNM
TUkQwPbG2Ie9b0DkOjyvbDzuxbGGNnYQb0/sbIhNfZwCNfbbkCY3dcKT6yrvzo2f
4o0coR8mr0B1Ryg6sV209jLq1PjxNJEsCDaUa/vlk64xUqyY+sFQPbJzAeIF381N
ra82ZWecV1lGmm5EAjWwbVyiu3CU1r/ILV0gkalcRtgssv41VeKunztpX/snZbYS
/7vYIdfaOwtEGzPZ82qjmb81BWGzs2TNQCidlS2br8Cvhxea4J8EBuT/0Ur7EgZL
nAN9KqQfNvbqh6ZQ3NQvGuiPi4mf33S3/R+S/EE10Ojws3ApSurA4gOVBSKKGvU0
dPF2XcH6OrbiJXyKdagwsZxLmUiFAxY1ZZ6o+0Z34/Zl3y7kV4cZ1J4rmqdfsz38
b/RlpyYWhVtKSQYKsDSuWQ9zMzzAzhfiwcKIsw8LgItqPMv9aiiELOv/0T18Lrmf
JoWEgQ02fNahty1w4+cD4iwYxKL6dBkRk5loswCHDhj0OOF0ctahLaX3pcLwNFHQ
C7yzqx6bDvPPmb9DIubgLGkgIlxCqVQy/PbPPF5j39aIvgZ5S7d8FwAKs7rGUvdt
eo/E6sZx3kMvTpBpxwJn70XeX8M/yhaLJ6GWcEH+pD6LmRD8wTgaYmGDDVHd08Km
j1+4+89iPoWU8ocYeofviBupIbI5ILh7aHt5qX9hZveonAyhUrXMO1kZGFVvzhBV
/nfEXbgh0viCiDS67MIJ/fyYY0KxjX6hR+5Eh6cnzY4HD5fLdNSLn3ok30rLHCBQ
HBk60+l6q6neVyhqHEmcL6rY4Dyr0JM5sVqYfsHRlfwATLNjoKHWGzXr/8JUhWpf
R/dhDFbiruQZQzPOZEvHEBCdaovzmKjssf+MEWPzj+eTNnB2j7bIPsbTiv74kE7+
9ytT0bm2xnUgTp7n3dn0jTCHQ3CpLzb5H0cqd11rMTIV7hRBHh2FDovxCHmrxYFh
imXrIrz3KWU3m6ehBf+mnlB2DsYd0uR0X26bAspk6Vl+rK9JREPkQjdC1ossdBwk
SXQUiHpJ9R/oS/WElbhHi+BUNsurM1LRyzCmnyo6vGVb9QyokRm+Wcm2hpn3KWvz
f/97TbVU1pn9VzjX8ncl26NRbmcfvahzWZgqoBmN7KFOftcHnSdUJlEGDOUJE/Qe
Cs0BWgNKL0xPJqIrbkiTHm+00YepQ2zvWXKTaWbzoZI63/29y3dq/Q8gW+pwsyqc
Gwp48h7gwtv44OupfXkzQzvKW6KdO/lUQumGyeJeEF61EehXOShLw4urJxAbn+7S
jMVomQKiSzAcBD7Bs+Ef5V1pO1tMf9TTuqzSB6KNAJfCpUeSfMngA5iMrwqAYtDm
pyoo2WKZTsqgxOUIz23HfQAikJ4uk/LdyKeglWzTPGggUc3ZDURBsdBA0mXC6DxI
+Zn2XhfFWjPTpH8mdQuuZ1drmZBch4vzseOml93oUtmtYNRKoiFJD7x7MJierf5i
UkMFB5U34p028KCvxfK1mEfoRFNYkhSih1zyi55/3gjoXqj6tCA+xk10zL/FG79R
qPYIT00YzbVsS0tOgBPFYNXBfDQLreohWW8tnxdJZ4j9oT7gzVpqGeef3caDYXYY
ijqNgXsVULgJC3KIggrWhzE9simrrSAt325d8olM2cyhj0xquooSlACDPg0llPPY
u6WEmVB0kggHbdrO107vLtVdZQp/iopePlARK9HTtQ7/n14X0tzvLChhlpngFFtd
cquSm3xJMU6wgSjdWpVujN4U5BisgjKsUQ4q+qO0C7Na+BNSv1qvR0ZLIaI1SXON
pGFF5CJo3zZcJr75UHpprfOxGjFqos/ydJ2FGxCVa1wC/6557hhH8GPZ9ApGVmjT
LZqXu2wbOPNkkgotPrzNdjXWH0H1axyWu2dRGw4njC4JuR//ipn9udcfnU4lXu+J
SkVk96MOKeiIGwpXaOCOERWJn8dMBagXKIefpw3DgbSDNKpeEkdMe1xxxwgatQBe
dfmJPveIS4sL1pUe+o86NMcjKpsNy+G2P+HWrpuppvYkD8oqIwWAkGC/XhiQfgOS
VQjbluPmE5Mp3Rb8iA0UA7Qtl3Cl7wyVGwybj9Oebh1EA7+fWiy6sWh2THsVES9P
i0ASCpFnaSg+l/U+lCbOrpLtVH4paem4X+JAQmJlmcDrWinpUfeYvBKMF2hIN2Np
Ia54MVn31LrUGZ2p4zLg0Cn0sA8asiSmQI+VOvif+dgXtVjSZDpuwvb8yxssR3B5
EaF2l9N0Ip5IrkJ85Kd2/cp3rGESCPk4uE4RA6gaCEfbfuNVfOcuQtEwqT/cAXwo
AGruEsVd58OLMTcvc1NMOj1s15oG2Zs2HUIkd2QsbclmZOHokiDzO5MdvGy7pPpc
E8Liwz3Fd76lyaNtgVJ8mRTCHrtXS4pF3EHcr+x/jD1NoGpH2g1WvtQj7lzf4POa
kyyP+0Oe1NL2i4y80Kd2qS71pTbHZsqh9vQFyVI8mh1nyjColl/WZ3WWkgS9zecz
3m3BXC59/P1b1IZw7zXh7bA6xn14oQFHuxrVEWr+w6SUkNhtL61iHzqgjiSDGdfZ
x1Smm/E9YysAU0F7VSukt1BbbyMQd+LymCyFpyYXdGp7gQgCnzX6Bi5+JN3B0DVp
aQSIXai4ggqOCD9kz0S23AfgLVZRNKXNpseh4n+w3begDkNaSFX7I/VUIUbarMH2
SPHYvGlgk8CqvV9QCdQq3rtgIsqqfP8QsQEq3o4YCHRhXi3OBVy5TGt6ql/WS0tr
6UFcAlq7FuDDgrysj2GdqapKVyG3SD4Dka1PQK3rAU55Ml1iCNTOsGuH2Aj61Zkn
Pj9VX1MNYJMF+DaTxnIRU3HK/b//FrXBPHUXoUaq5CEvevwlCcFJ37B5/G+xtm+l
2YFY3hJ/R4wq+PJDbeAxF2n0Dkr7ulJa4SfPMzHNpvYWZ4rDRsCF78vQYx/ae1et
WmqRpHqY5FwxkyezfebEezT8w0Ju3sOPRExnN/eAuqefxiAqLXjBCfpw7Biz6jyD
r5shNZcWzqo0y8Rax1+IUHhXt4+BxV1d7imZabERe/GgBjaz3vLmMCr7QhBXy+b0
7kGRDRVg3AsUXom7MLpHtL3bTRtvwuMWlNuhauJ2ndfo6m8ndzSQDXDVcmFXK2l9
G52epRfTeZ4qrpEHLEMsc4EFh9T2iXObMymGxA2m69DutIZVrZtokBKyZ9rmGhch
P6jVAFmbUUyAsJ2UMdqbHwUBdQdMeQEMJHa/2HZxrQuIgHxSJgRGR6NIsQ1g7nwb
oRjMwB9LBcvWVmev0yNAMss/jEaTZ6KofkC8v+P6S82iCME8ODSJKcIb70etUPqW
87j80drlWsHAuA/C3IiI6sIgWfbqA/Mc+OzuHxogx3ZTeAU96MnD0eSe3fug7v9x
fAyRwWr+cw5nVS2o8RUKM3qNlujqS4VdUE0XQFxpxv3NcG0iCWfjOV5s7BPgS6Rm
EPB8Znu8pRn3hZW0z3LcMYgQYMTAxGWedSHUgZcRuMUj4SsvmIZbo3BTCAgb0RAY
lU50ylgu1/m5pZYxQaMgqlVaoZNmASVzOyzVO2SRUClbl6AKyHYVnenXUTW1UibE
gCUM6A1u//GJbkgt5LQMUNhF6OejejrTq3VMNBAi85RQlrkKs8XswxVziUyW0tT0
GP7PeOgOjigwNrdG6qR2i8RwSP9J0Am3LsDaJcs+xOcqRgQx5u521lpBImpp59d/
z9cDR5DvfsHgilCrtLiNgAcRRZqevBX+bJC01moWXnESZh5ORSii2xbdqF/v2XwA
4kVimAbYB1mppAVEjMZCd5INqFXvaqOBW3wVIFjqP/AQm6/pPGckh3Y+AhkMVOcc
RnhtPXzOU4DlUkgqPPPATv7Ei1rww+dbLegGSB+wdS3GGqNiMcVl4ZGN+MdTn8sp
5HhJM9gI1XR9HOjjwYce0g37bmeexSbvhZb9AC8j56LjB1dxWMcyU1sDdUFAZ/+y
dmT74OcY7EH0pOnTMURtmSY458O+2LUfYrvwdrrLq65mqwu/OkIJj2oUf0Hx8nUL
vRF0e/rg18OwyHUP6gzRkVaxnGDK3N/N3+uztNn5uxS6kioGMDhSvS4+gFoc/vj9
0oioGbhDphB7z/c8xgOuKiwotoM6vId5Fm84zEx00YFZtdoA6HqADPa39yy13Km7
9JcR7iEOCnkxmDifaJWuWyzQ7Q68WqLbrTI9I2VDuyw4ffySw9+Z95hIVU8dANvl
RmqXaELB8Kk1Q449YYv/ytZroK7qm6w4WFtHjWeSvhcjnjT9BonAQSBNVnmeKJMy
P0x6kxNcZuF1qeZ/57cvI8rVCxHlG+zbVbEe5M1htwZMALKlDzGpskhJUj+bVFA8
e9FZYF/xfNX3fKMfl7R7VFf2PofqwsvE02MJS6C3ED5n2NIKBHVmH7GsbEuqCEcb
VEqIcYZcwf2eladlPeTOux88ylC5js1e+H9CuRr9BwfIC04VJYXbLPay21qOIEa7
cmmiIzJxNRCj6q/yTzniVTWaQmsSpWSm5ZIJ6+oARVOcuX3/u7k72v8MZCnDwEVY
QDGLBd9UAJ1M5i6xMPg0An4vUCYqZxfqGhqdROrssUISWeFGYnatHJOO1UhuGWq9
D5qvf3Jy/jxzmiD33+ScCOrmCql54ah8TUZn2qKrhERhhNwSbTmnSWbpvlh3F1Fd
ujynEMUopTL3p3AEjVj3BLteuAzpxJS1vmgjJs5Yt8Rt51gofm9NQQUVO+JSfaK0
oIZzV/Os/q861oWmCXZE9l1xXKScc68t5HC4f9VWVKR19mht/l3kNx0IdDf9nKAO
+F3CCCQiegaQnNQ4Ic95rP5oS2QN1sRivrIAyCwoxMC+b0jPgkGsioWO16Gf5odW
P/aNW2QZg90UpzxZyajXvejPiOhpU1/8ZxQQUuu9qlA/JHPQCaxdoKwx5mA8Jw8t
quRuhPhRC0tyq91op8T0V9ELs8lVGdqW7uL3SbTg+QcAvMy3lzXkCrGVl6CjMflX
KLqhVbUVRk7YxGD9y+prcoUKo9pR2z0TO4NyHtibWzJKYiIhvXKomN+KRh+1aP+T
UBRovnDqcAiz1zAtD4qovAfRUd1tcroxC0r3xonaBuQQ7564jIx8146rN6XznFL4
Rp7VQkZ/91CKMC/pAqpAeXHrbQFHpPyEpB3DDeOu4mIf583cLXFemNEV+dpi3R9G
e0inxV3AU/WdIxsi3NSqbKvlSE1+8R2ZsU8y9Gssp/gSrG4+pXFYNIaFvoTklA2Y
7Y8i4E75hPEX+nl11dWZRXznvM6Yw9/O62muIqRwCgewfP3XZ/qnpyc65j1DGSVv
jIZ8jJxAnC/zj8o/h2yp83AmyEvKnHJ9hPN4qotKyF26vqnesCft/rZvgOZC6USN
8w5v2OfC+NE1D9vdRvl1Mq964lX2HB0I470Ev+Zme6TP0MqY71VW/L35qZmtr9kf
g0nxcX0fmzrUzNe0n5X9Efm13Cwfc02LKgTOHJuftS8DCC5DZ6cok3XrXELjY7WV
1ghMs12ew/A3EKvYL+NyfsIrck+XvodtYympDkIK03D7uwB2wzxdPStx3qRc4gco
ZiD7j3Ljt87ZbnE1z8iA6CBOds/atWG5vCgsJPZFXpztY8Bij96hnBEQ4G0dviL5
t128e3qzrA9Jqi5Q3YPUb/aBerk9XFRqReqBfWs8GBhAllgzf2raWoFaGwF6iIml
AijqIYHmC56nSaxkwZmPVPCIEzUdil2ofmdTDoqaT5r9+FCT+rMZuwyI1xj7iibR
/w3XHWsaEA9KaH0uebIANqTsKMKvn2WaBo3jawf0AHqBjzLusoousPtVPtALPpNM
YYQkVVD96JhOTuqI0bE4EWhCya6g61Jj2AwVE5+RniYuDzvY3dhopl1KbB5Xvozb
S2lZIz3wVW2h1oykBwka+7z6WpXCsEX80nqtvVBGwRZpdWwy6sM7UvpeCBJiIKSn
1aHsossFNxWTSBHrCAL/twFNv8QdzVyjtDzm8GVLZ/qhiXcaQd40rYq0v5TIK399
aKz4X5ZI4sS2AETk45kIjvgIeSlSl0ISkRH/xTaf+vuAwY9RdghILCMPMvpKbbWX
pUaKUGA5cbygH9nlt4B4QTJCDgqyTPBAWAOS15r8w72hd4ZmvuiZJPZOozP1x+PE
QjU+Mo/6PqTjLFdrX4pLRIUSqdKLeDL/rqtSOfDEiiSDNjU9LwZDEVLGKVKcBQux
fo9t8WC272KGSoAVZUmxKOTw/vNcz7+81XToOOAvLwSrVzbA0B2BA55MRPfspgu5
gg4q621M5drF+65I5dEnMjkQQOcXAoDnIFvHk6bLjx9p65uGzCVtZUzC5G13f3rZ
EgFc+kiIX6t8s2duAcTEFnIV6aEwH/ek3xG7d5CKGYFMG4xnuZD++n7plldXiy5j
7kNhsEGFfXdvyRehnld2LccMyyFd75SCLV5G3BV/+CpOesT02GmMQLh5YGZub8do
jvbRCMfRIFe7dytPGIlYvkIkBLUTQfS+NxWk6Y/CUw8hHE05OQvvieAUIZJnfnFZ
OMPrXlRZjPVZovayeuKvJ7qKzNgFoFDVGR9JWx0+j+Df7dxuFh3q79xp88f+F4K2
q8rRNY7sY+IPA+GNqaw0O9Zl63LjBNv2fPeJEiuqGyqsCIbb1JRgGSnTiMKfTzsn
HD/Eklg3bmmyNcRCr5eNy+dYjDBV+83yQif1imqvHgcdk+0Xnq630QklzOcqs750
g/bPNbRcUI1LO8sOiEpHUHKRqGrThuASqzbZ1LMv8JzKdlICqaZzd9yCe2+AqeSe
PiFEAZzCqMDJEz94Vm1POYxQn2a8ozlWLjJBU9GwnFRxuAxxlmAkmDu/o9q9Dx/U
UMH2GoqMWQIYcpAWyqhEZc1GX4+bYO4uwPM8JkrNCOo9Bei9uZ1RlIOVWjkQb/br
glMFFW4HK8L4Mg+Ywjjb++YeNiyz2WFOLHBlfbKDhSvMgX5OXLSX1fPr8pCCvXuG
GXIkFzXzjQCcl6YUshh6MbHAmVAUY5JgXI0X/IdSHfm2rVgxZUbmrds6xLb0A3DJ
MfF/72w1r8+CwflLAhoPv5q20nY8HSUUDliwcKdIKU1PZMu1wabMIGhKQXa9wGgd
lb/dqpYiQO+0lxW8ydkCKntpiSQvYKftr8MloczKA9tMkUPt2rZ19B99MJzeO4gy
OIQJABF4HTeZou+m/ZkN74tNpMc25k3oeqyLCdExKo5aAN29EwgY3YUExoaf0ja/
dH/oHlZrqVo9u/vat6WHakx6oFnaPSRi3ti9qYrYfADfB/aPAzgBe6iya6XTBLR7
0f5EvdAjKsz4AXh3Movnc3tzXAMs9TAWuaU62XB19YhPhKLlO6HchhjmIsiOG3iM
mQy6fAx5+afxAN+yY7iN12v/oPOfxk/odO2HUBxvaNLaicb5DQkLjURtLdqyXTBs
RPlPOwYZsudlgtjhFHt7viFwWa8L5HUlQgJ/KBX4RQ5u9N48cie34AmmyK35/C1i
K6s+0FCsJKT47fo6saRbV1OrlShykrbVmA5/6eox6jLrrI1AEb8BUs+i1tQywJ4X
2zxhM18Dt1p32/Kg68IzckQmfQLiMvk/CnC1/nynbGD7qKqWaMEEStipTUxsjKGO
vWn+kbf4ELcconWV9IGah3zwHUBMRoaCZCY3ixufsthdaDVYyjeJ7uvmlKttjPA1
9WXMNzehmWFmSdfS8Tl4Ydr6itmeKdzqDpGqfLq84u8t+eRP0rpls1mZAyu9xuoC
IKypUgadzd79mVSjPyOMUGjYoTYGnERho8NQoHYOA3vNpUepxNGmsebRd/6EE2DA
gvh0YlofU9jp1ObFvPNyA0fdhqvpzSab07HsHA0Eb6ap0fB7IbvNBlvz3O5WB8+o
m8M9TMAYNeTQdFEDR4qYSj5rNnBiFz0uG+4qP3uKtVbh893MEcNAMohJLi1g8nHq
OP8MHttv/EgA7XSXpnJL+d824k4z4nlCMs+LAJPAhis8yTO0ovTCHRfqszqRNYQt
XzEjSpAWwWks5iXh2W8NsTVIkUslqPZVt194cU+moOrbmEao1LkBDyVe4BPpKDmw
Fn4lOEwuy+qI3rqBsuLhUHNLhEJiKV0XBkirZDXsE6P9gsXrqa3OV7mMutXAq6xu
Fh6IH0nu5TtD2Yus40qKvPBoAH7I2/ULAljbvTTF69KNAqreXGJ4XZpQjbI6iCYQ
3gg1C+ZMP2Ac/wgF5NqXHZ9r+f5c7WmNJ5gC7CL61+Y5RkPqzvlpo0CBCeo/q6TM
eaEsYaUpoRHdyV9a9R3yB0OSUr2Qo4XljhYPwIiwssyAFwS/Ef0kwfDmfQXkPAzp
QJSLawi23F0gi7TYSjWFSLWOFPhi54y90u8M1nMlGsJP7D26N0AoAUL/yvFQBSpt
NSJPNwlOW0iLsQHYSLuYNBQnUFWaHtbKQc6Z7UHkRZAkDiNOaYRNBmKuSG7dQDDV
DYJBVNJAFuYHvQov2nx8/hdxZ27t9jFwq7bMTada72M2GwSQeKRkZ6SkFftAe08/
O4WVq6CaHUZNRclxen+LrQw35yHiVlynAjVQ6D75OFGKbTsdqXL7TJTTG29JwUQC
DpvwMH9beyAahOtcUw8o2UXcKYoT/PD/T+5VdsSeeiRK8U8v0FuN0Ut0trdgdC1P
hrHbES1fSVBqYI6mRmi9IFuqryBLjQjKfMx5hp45AGEYnXvjUMRMf2e5H3qSxezr
QopI8J5H4iySB78FDEhrS4Tb//xzQkrIKtzHfc4hhqtKCkYP1WCW+lCGwRzNr/p8
XACBjS55BwaVOP9DosHUZsCHWjImOOHzPAwulTFdPxllPpRZDVPiH5D3WvLVKdEo
M3S0IMyQMfUTCdn7ipLmlR0aG1Lr0d7xeM6joZ3eJ6pMMvHtE6Ryh7lZu9T4+N0m
2vcc4PmUkESjAQFXiwHq/DX8M6uI/7zCNVGigBtnSPxNwDu1nLQFNx0uLI2ybWPx
839ezGsFleTBNKsjvO2hBpnDHVgyierunCQAX/PhVy6q4iIcAwef2pQxsDC9mNgV
ihiE1YtzNPsZDCJTj5J4umKz1107b/8f/csX4eu3pL5fAdkuRu+/NJ/zdkr1WECs
5wZM2IWQlczvE8WiDax8v/5GCvXTzz8x7hOurscB6LCAVi9cTNaoHyJ8hhj3mkKm
ldYcrrl9GkMh8CcjTu/+3hZFSuv5hsmKYwBuRjmKElTiTPSt/hfIm4cUVOnlV6W0
5OCWSCvGC9T4D9h5ty3SE1UQ032d67HjS97Pt2fF+2hmX22FqxXh6slZXMtI39fX
4qCfHiQTU5E5LUsdlWORJh4FX09vbhldvU57UHVcXyuoduviaoVaIvTGFhol/T7p
dhrUnrW6I4HvRkUDoaUNWIcWacZaPiNPhXTNI/YbEOSiapAC9FQ/PEW2yycZITCc
Qwb90qtechy22V+yAryUKO21NiXIu0WcZaejoqx0LXGwicE+oVNNUJyStmlx2PNs
E0LQ2fSIKCTH7/0bJ+GQjp3notdsH1RdijnNvNLS2UgREbluRLoKEfpFh5X0y0kr
E5ecKinNrSVP9Cd1GuWmFDS6kM8EfAwYH6DH01ML+CtxUly3/ZQvKjsfOlnQLaRB
ML44UZAl+HJCPwwpQxE3C2Jx3FB+QLRCAmwQkPVxKuR0wnznykWlck/BnoVfC9tX
TPdn2j/B15VKKbB4wks8wA0GXqoiY8xFaKm7uAh+grNFFc05iElJ1MGsUtZtbF+P
pJtgDHi0imQ50HvEV+2B4LbstejoOCm/DyqsUp/GEvx+SYW+iKK9YbpNP3fbtlCC
z69grvwUSHJ+qF7J+EFzHvMzjU/gAA1gux4XcoahTWjI4obwYecjBDs5HWphnWTa
2gzgX7iG0w9NYPeDwNiXBAeIivmTGHeQVwgoUHUeL44CnHmB8NVpwQsn8vFFeEcc
krrrT2jPJVBlASFgY98fPhG2r7f3ASUrUXvLVQ6sbg506t7DhKsXZ4+br/YUSbI6
RkJPEoD4FTOvv0GxvEP2Z1OiOfTa1Plvm7rs6ZqMgC1XyTJOfKjPkHyBzJ7mvyX9
ipbcDtIOJbSazLyJvCvF2OU1yX1uVwGiuXrMDbVxmKsFx2uMeL4qMJFOtl9Jz9BJ
bgWMPqBkH+gKiHVnNwlfeFhqtbcbfTrVA0mtcrQfRnQ13pMRu0eoVLH+Wv2Aypmk
7PZYcsfFVcUBK9MoM8HlBpRLC1sCUHK9+sEom1pJISnRebHHHywJNNhnMMFLZQyy
kbqOxDD9YTFd8CS2pRZUImju8HyOk8TzK2baftZFib0Rl7nT2jnMNm9OLQ7egLSY
/UusJCftXyabw35PwO2wFk5FDkBf38UAKxUOJHExHmsWCDIbaBldUnBzSfnrMms8
Cedenps1gLDUl1uu5GqJGMRppcWcW2XbJRqx3W1VaHUfXlP6lkKo5p3zSR25SdqZ
EFgfUxkHP1mEEyUkXYtzgqFUrirkk40YhT8dkgeq26/6oGHkBd6cX6oTRJUsomz7
/YWmAjNcYEkKy8EHQvJom1yswlHTgJjHQSZqLwvQiBDKhoA1CAT8qFGD2CioF7HP
Rl979+hWRaKc9lbKtua1WlVXKR/Fcf3mDVWnjV4Zldo7IqN5R7u7P/Tv2bOLLnwZ
vWXj5ckEb4lLnERRlGHqaVy304m0sTv2Wqh3b3tJXNa0uw83SgFsqZeMwHNJCLvn
ogKr92NiLdWpm/j+rAJiDtPI4RGCleh9X+JRTZ93LYIUZfAWC/kkDvIxQPCPKG+O
kpPfISNe95KpYwDY93Pa7dKwxQx5oyPbVX35jZrCgE9PmFk/YVGqACrqpptWOTV/
EdgPm+PvTyri58US8w0TwxUvW+TcJLE1wD1r+gn/j1T22bHcb9YNGSUwYloy9rBn
K7me6FUZQENdgmZ2Zmc9YdxwG96FLmu27wRU7hL/epd4kLF3LL+Bd+edQMzeq2lx
zmxYeH5/EFxVnxWefB+iS7vtcX034V8bAqiNbeeyI4RQ1wJC6AtrNwLbQ8AF3Fzz
boms8MSudevd1XVda4XymAonxuYzwcUHJDlZ4+L1Cq9ayK88mRLjzywj0YjFdPJG
AwX1aFx0AANA+Vi1v3caV/26CGY1iG5CVjyg/dpvFbNimey5jy5qmJ0AfB83OuBM
IgeGnEHvroZNmkbu4ln+kl+OhlA5+M90pyln3VGpY2ke0v2OdG3VAAvmuP2lLC7r
LjZUVBLejUBWDGX3E0nIVETqNM0qQSinBPKzW2Koy4DQXpyqDQcK7q0onBzCHvDa
AR+40/RsvNlA94tbsEWqZmoO6PQKP44GOe3hD2qH0huFT0swJ2YuZQud3rvkun53
5xoE8kc8doSOAbVoyEsarDjN/MSlON8qWKsu2DgBcmW+zA7w8EOJ+iMl4rWLGPNm
Ax16emJez4Zx+6EPKgv6fcJ7Yz24RJxQY4V/jsnZTL3OZ6N4D/Rfn2Mniouul4JT
OuL0dsWzcPua8nWoCjRQ7nAfpuggIYHRG/rFPkGLiQRFzOu94KV8EqudCaeqQas+
NuW5F2KXfYerqHTeT6eDXbtVYdJbhBuk6WDJxSfP96uSqutjNt9v24ZE2XYCHj1i
bvfAhkEXrT+gSqQd3oY1b+g2Pbw1n4AdUGKFePFLSTWWPCxITNZr1IwgFlsJuoaE
1Q9e0W/c/RS1Vih/Pg0tpWZ03alxwh9CpDzLMvNB0ul4MWTnxnw7vgTHJvO3FdiK
qSefSouk4NJ96owRUO3GIqolTH7PGazBzL/pvE+nt1K+pjyeY9ulZZYpYzA4NfjD
2IptuHXZnQoq7evZLN413Z2qRJv6Y3fvFEyvxvBCN5UHF9pyUpp5KtKXOOAUwjId
J6kS9AuOC69h9Beqwu3VqRdkPZbS1+76zVxTAiVmi7FsZyZolf4t9mc1zi1znlS0
u/AVsH99u+p6jzws4G/IzGgNTv1mor6ZX8oBXjNdvwlI3J+6iiHKyU135x4Ep6E/
b7JyANmPluIQEWCCp4qygSeH7VehBq/Qygdf5ND7kr2AaDt7n+48wpMUqMt07mEV
RkQmqSqR20NCMyBSU7WDkyvW9K9gOeXw17UWRYJBUW9fpqOPgA68zmFdxpSplf3W
Syz6lAo89NJryG0SFIBMGUXxZjJa4C4pz9t9ww4R4DAkdvcYKenT7H6Y9aKdvdcl
5b0C6IUSoCkAW77+2i1aor39Sav3temNXwQKU3I0RA2jexIIfiUsrPJ5sN6hlP0D
mTnBSoDthuNUZtFZe9ZsgvxvEL1WAMp7fIAuCLzp9zhgfPwt6XmrZqH6SMaj/2Q6
hqaWtVYnF4owCFCLFEvcRVemPs962zx0rLAoYf1TkysKpfHtlxr76CvxSk0CkX2f
ntiyc57EWbsKemGo/nh0ZLT5VHuwLP/A31mVjO7A2yeLoPVf8DVTuw03V7Vb7tbn
gvb1LkhNkTMU3DVmVPDk31j6RqKKJiEAkIeEEXeycSco3hGGJvuoQrYR4PZ4iI2N
MtO+XeKtWOfYv0YehY4dMhfdBTnj7y6xQb+kvZ3OnQryu8l3ks9b5QvuwQvJu4xu
BmTJtvm+B5hGQwkIoQTrIprOppEsqcWDnvHYuZyaIpLUJo+ODhJv1QEECJMAPy+W
Fyuk1aa56rpmNXkGJZRN90sQB7Fwes2AXFQYe8n6CqJYQ8wmvGOojZc2Bh93jwWm
q3uHgtAhZAwwMZyBYDZtLekgvNu8XmniSJy77/xTbNaBSwKMzAuHhT9LzmxDZMcO
+jgh1HZX9UeRqvVinmQTIaDa2Bk9JiA020mc+IVKuijq3CL1yGL57yPB2sJKF/GK
oMGPCDiQZNQIvuwnmTEXY9HaIG/G5DazPS/PQUK/di0WHXgCfyd8tOw+l/LM1I8m
araz8bR9FxICpUnvA2d+ef/RP4hyn+QgJm5eZ3nCkOVanX9/zHr+Yf+hg0HI4niu
qEglt4MBTXFVsvejv49BVHQ98M/LVCwEDBi5enwdoHaLpxWjOy993tvxkyTAL/kB
qkK9BLpsVYo/IQhKKXV4RObWgRI/h9iF1k/amlwaFNh33gXbrBx2qMaohRbXaa8M
wQUN0Rx4BTJmx8Cktnt03ZZ3de3oVRe/0U/vvxE7W/SOdTmV4RdZms4rARz2558E
S3Ma9QX+6GRWAl1A7/tMMtGQ8PJwZXyRvCcKUJD+hJISvn762qoubYkTiWqTNuNN
NtPQKCd/n7z05XluWIX3dszBBLdoOMng7gGd5uj5US128AyHgSZZT/cuk6I1PsU8
UPuEZNoh3QKf2OxYmoZvoOVbGuw0ZiRg6MZd69CTz/INXbGU6uj1FkmyN9ZVMRPF
jd6XxNY+O7G5IQRkHPc5jCqO9GrRImH1M+lPcy5rdR1QvdqZ5xsXx/CehLR7rHal
8LBnf2NyiVBWruafjjxTA/iEQ0efJrwJUW/NPiM8nNdHNHrfMAFO63bEjlkceVPm
gZmUb8cN+uWaTF7gnzZteeZuH+4HbvlMsDeKAneKsmG6FC/jNPsU4SvRY2S4amGO
mMEmLY+k9S9WKjct5a2RA75yqrzZmQUbpiIZgXDSfmNYFY6oYUF++0uMsM+JaGQM
zteOQdMPajoT+KgkiRakz6GxU+H8Pu/aJui7UZEu2fH8szv0kfgTZ6d2iTY+2Afl
lF1bmR77x3hh92o5cxY6GUk31ppCb7wExZvII5WsoU++fNVJ8uhcyDO1N+DpTHcc
O5AV1HjEKftN7w/6VMRocr1eyhnk8xTEcjiNS9eYsk5h9lRjmxure51icc2xNI7G
fAuH0LVaGAAuhK86qRzY8vXDcFDKt8L3zvocXyvrvXZnfi5zsZECmb1yBW5PaLjr
/ZoCZrrAua3mKkp1Saf/ZPg9eo0RcjLnPtISZgHZZ71aHGQ21mqrnob/rVKXXlJd
pgEv/D6K4cBUupMTeadpgz37V+yzJi+1Qgfcgd3gaBQeXg8P7IjtQ+bXPCfF4tKN
8Y3FPj5/1fWE6Of+SlwsBIp79sfi+OdpnPPZhuWN8kADZrGJTuiBPApLZJfF9HRO
5KUHgczDk+fLWYKlGF9i6W71qobsVmrlhEO03p3qGlmMwAS5jgTy9thnx/5qq1Pv
X5kcpJ/HkByC6mrvwh5D/0ffcGuB2GHgflBkDg370pOUMzncln9aYCAs4YQoGzvK
3oDxUThSOUfeyLNhusBpItkMrTUXV7EFkj5hoaJTchPKV0LhtIdZn6RVodj98QpE
VdsKHq3oCz/+kY+MbDpkL0//CakSzOpUc6Ns0r7BSwHuzQDSL9hmMD4x7/BRCp5W
Tuj/oD9p9/qn+BSGFV6QK0gIAW4yMv4rS4+QJ/c7cRXTLqEd53peJlRSCVNN5tUT
4JBIYBstc8PTHxMfrzPHuC5gDn1vc8BKtMs1eQxh/ePX2gI80iHaGruD0Huwtivf
IvpPx1hyYsN7Owyu3vBI3MdEBx1BzJAR37ht6idGN31P/IZNLG5ocGBftp4aIIpO
6Tos541/zxcgc7l4aK82ANbI2hYTaPrIpnmHLdCgNvAqSGhIG19utickP3AyT4wf
m+iAocZb0BLIKdKN+W2R2RMUEf14wJc5VlMJa1tdA6j3lu/MRTURbwXRdsvnaN2j
nl8W/98DE41NXqQ9k7Y6hlkywQzkEE2fTZmvrzQcD3Bz3JPcVFr6UQqq+RUzV8oC
7jdcQnOdVh+g7gZRxoeeKzwNDiO0RP2rGaJ0OM3i65PQ6ZnL1TViJF9ajKzSw4sL
06DFDI96FzKFa4XhJVHwOEhF3RCHPNBEu8Eb0F0FtKuHAVTqOSwjFHFNA0mda+kW
ktnVfVsjJAqxj1X4DTVIOfGs5YBDcTZlr+sm/dKvdvk2CHSxAFXbX2OyEYCX3iQv
sp0n324eKWZDF+/gbjDDUSS2IELH+T7ru9EfTMUwHNnamZOMz/38VWohWlWxR+0W
/lsr2IiMaRcmNZHbBtMmcNFCfRKnAt7XKhC9uFaaHSyhT1fjZJi2S9/SkOnEf5EV
wBgTZ1Z010O5BBoPUvp1Sgv8+fSg+Y5yvpVH5JDMt7aaEv6lGnMuoQOUGjNpKo0t
bL9qJBMHJelNs4NvKu3cnPSGr1DLM5my1aBJIxX4gRdgFnh93lbZFljrWfk/6VnC
VXordqYVSKR7wLHTw5RnjXQTTnBCD1mQtIw9VsGvG7tady+93NksLjs/XrVUs8QE
sW9XqTMQYF8mezVLKFY/2lfDM+yvumcZSyKoRSrg6vx6oI2LsdH+7NMkgroUXToM
c3L2wr+qvUE+h9fm99C2/XnCrhccFhyphlvqqi18AQGXg5EygYRX87si0h3G00zz
YZzQp4DxFFoTuQUB8cDaUlfhwc014GLuoxm5ECEwxnEx77D3vc+OHLu16Rxzafma
ziQ4TvsjSXIMzSzx5mcEeb+K1xU5NoeNdVhecMOkkb4aM7lAqCanaEOsCjvAujYY
o8/cQ8mZmoUPRHmX87wdOHe9DhL0MUqWOJtEXIQ98HC4j9T71oXZ8bzs3gY3blmB
aTQrSW2zkObjHRhdjiMuWwTAs44eUbrRjqv2bFjtSNQspkSmThgbOSfo+/vKAybc
nuu3eNkGR/d1pA/UfQeWzEaaxOW/GA9agAHlvI36J4Satx8T6IM60C9KKXhYyL18
ikQuQOSGMx/4j6UixDPRw3CTd/MHv+1TO/o+zpN1tnW0M+zNmtUxLPKgNOdHPtM3
cBYNBFQ82dgyCTMFm0fZYp1mNZzlM5OZettUmWlN8uwq+frZeLgPppMA2xYKzseO
KHsIRUBlaArwR64Wau3hLofBpQxNRXtHfxgiV0wp6wUATI6Gc4WI3fwt7nIrh2lS
FuOu/e74YW3l6ahuFZV2sQ6y3pa52AZ3ONTe/RsE3SW788avRC7Mdi7BwuPLmRk7
Y27yV3jyruDPYa54mlR1CKC1Opyct0E8MswiMpzdPp8+EBIela8MyhCRLJAYLDwF
rGLNRtOPP7Yj6/ak/WoEcAQQ1MjnNR0mXyD56g8SagmIiPfVBeJhk/uIHJfn8zf8
0RvmOo97X+aAXlC5+u5cH3ZCzYjSV5q0CHr4ZuPqJAZ9x7oBu2cIuzhjDXVZtk6N
utIoRWWARHyu1n3yOD9BXrJraJTEo6OaZgYoL1S5hv5W1RixZkdwBpHBKZvO2FzH
yAREbubU2wdBhXwcQIqtrmreZgk3PM0+TkNm/WGvMn1Fbjl77FR54AaTWrGITrU0
NOCMPiEhxCTV+qypl3glGMeH8C3KIPKEJFK7MO+YH19ZicgoNZpAOdROC1TZp5mG
0Vlz6/1fnDsj2Yx5liFghXbJnJRN12iHc6QcKyueRzBpCclGobGf+O+4ibH3yVtU
XRH6lb+jW7y11sh2GvzeILvOG1ekPAiWAjfx7FbTx03fu1S74k6SDIwafA3vMMwI
KgGNv0LwoXKwNHfvVGelO5JSIHU2V3RiSfztB+40S2ItKm6SsNPZHZ0LH3+OsLbL
IjiTr1dujqAqRzxFYXI3SWqnGX30LFQe+S4UrmGzIjE0LPbV63UZncZ5dAS0p0mt
E8reFJ5sC6oDGaOTHhCTmH8ziav4oH+4pWqVTM84Iw788D45SX4/j/sR6sUafc1x
kOZd8x9iBeW2tg9+UBubxIPsW1ZL+qorsiQfpjAVIghfDuEuIdcMu/DV7oqoiaH8
tho4uTLUbsu5EhhxQTxJAWz59QbaTszaMGwe2dciRDoFRVKRGULQUamHdfH9a3fp
qRBcKvS9CF5ELp8W1Tu/RKzTro0gaxsvRy6omsKfX0qYt+k6JsTK2JHjdj/XHo8K
2EPbCMeD4K3rirnDhtMdLZZM6YcSCMzt3Z2u/vMbwcsREl6koC2fUsXLoGSFSapf
pku3mjas8FXeSt/0k7rHaT6szmCMgm5JWeet8kRBg/iPVva2fD6hHzU8nWfjTGiW
Mjg2XOJFiiUG942qpe1AyOqSZ6IxAfM0XTRWA9ByWWI3Ce0RV9evpWcuYg6sZmuN
s0ktGXjhR3h3rTadNk0AaKxZZA/b8b8sLxY0MyvJVHilTMmXzWAKwM47ex2dJcW0
PDE432KXU+yi5DigGQeAH9Sh20591aMgv/ophvcsqFNo3oUxHwCla46+hTmU2v2C
++m93eGtYi7xcc66f4lGVkzvkYjJGCn0uzuLeSIB/H75o9qQ/54Nx51ho1Rkaou3
lW2oqIdWIkCZd7x8G2yNxmguh9v7N50Ivy49CYR8iKLmizxGdfxikiskb1+4464L
sHugnwaF+bie4ayy4V8P+7ZEZU3P7VEOfTYgdmUira3JGiXDS92hHKswS4zcrq72
xBxD+Dqs5TUv4Gcjm1u7ifGbOL5fw2tro9kUzaqjJIf3bFm3+hZ7gOAt+7foKsqt
yrEoCxFX4qMOMiVIxUtbEBWrbsTowvdKz3N44pkrSCNQBPOb6fZQTJspzeS+BGoG
jRGxfYFc55vmBCH0CV/aHYoC6cTMfun54yPLRaUg3yNRNGQcfo8b+w3G6yVug+RP
/k0ljBaQSP/UdZal6LVngF7N0zF5uVwZYZ5k7MXRLTbdZbca6+NUyKwskaxh+122
lY8pPu/egvCj9G7kNDPse7pF0L5B3nRg6fBNuJvWKnHJpsql6x7FirVDhk5XeA6q
sRdTe3sMdZAoJojUFIO1ioOYSyb8jyCciSkJtYOcjKcFdeqGdl3l/IPu7+J4tgPi
PuQZscKBa4e56pbtZG57oZvDlvLvL9lAyvH+SAzUYfPzWZhjDI7DDMa/w2BbBu5m
0UBpvo7Bx7fKhlMi10BRs5hyKl2kVCo7hXcgqeLav4g8nBmuU3bCppCJ9Tdb3Ty2
Y/WX1AnDkRS5CZgaexM/Iqi5YVyuPgB1GskpQJn+xedYXizTDpKBQ6llVdu61Oxn
DnhYdiE7bqz5IfXfXrxzG3BnO8KRSHIdxWlVJz62DvD9WSHNwR2+Dh5bmhVG977Q
YHr8mvm6tvoxBgNihINqjgpQYgSDnUAIPJCrD9/CH7SJjrI23lV7Qgh3lQMWpf84
CFBnwt1yJ3FsXCYVFjSb2Mh0fbaqTO7gD3Cm9vHzSgdXg/RVUwiR6mUsXEIRQYza
+X4bFfEuN/bHpEMLEM8lkDMejAEJBljL3Km1s2+bPbYbMU9+JnLPPJEihnPZsOrJ
B/f3hu4uhV18XTeo0hU9UgYDlEfFGlZD3AePurTMKfAzpDfA0C1aZVkCarh0wlfT
8t/Xx5WvSaJ8kTPCbRCyKsuOboRrRcBKQFdkdZIlq75L9dDkKbjL1ZK8BvB8178Q
JpMHTJ4HhfgT6hEZBa/Dp7My68qLD+je0nvkj3dPd7FlFTs6ksdLGAcDBW6dJ/Av
v7llWEBbHopwYga06pSVifqeRXPPVSXnEvSR5Wvo5Rfb4IMShdU1vE/RyECIB4WB
s9LBixI7I+lLW93735X8StMiuV6qFxwLk2fJcyzvfjvRigSevkpF69CI6pd4uDl4
VDvj+Fq1nRQVWu4R0iQ57otPv7IRgpA8wcc/9pttt5n7BfoJgtY7lVdeSIO33hBS
lfYuRLEq9qXOiXdu9BJ66rgmQ4eXV6kpA0uE2wKnHN2FTSDhY2PWYIpaP3Vs4o+0
pJInpd2abHDUDl02QUM/YZGWf7CdU3fhCMBaQXEBcGhymhbxCy+xDRHccJdvTlrd
MOcdDRmaYluD/C+2iSc2hhBhDCQMqx1tVxakPvdZNjUrSI2tsFNOgnn8Ss1RwVlV
Jyj5waJ2RU2D/inuNEkYT8iLK3MDA0P72YyvaXRlhTMRoa7yQG7g3wAuHPwfqWHX
qcX4BWNLcvw+QCkBoApIeW2MUD0MrCOzTKkiF9PhAYQi30ye/i0uSf3pr6Jseuc4
tcagMwPGXmaGOgzx/0EBC4yQKckSvt6YE813hc/1899VSamsFeTpd5bGlRVvrqYq
W3r9Mqc0xKJ/FtixFuTL3phWTkplnqPFIlUQRPDWjBuu5+aE3errpVGDSmtO51EK
2mgwq/StBBz/XBHNYzARSGtP8101CjDbPMJl2aaVlFoyHn08pQL4cnD7/SI+LgRK
iJOQvP7SUoLZgzLHvRF2jlajDVbkSOoP6FbEbMMH1wYoqApTKWiJzIqfPCt8QZ6g
qeehQlQ+BBnjKb4Blzo62xH78o0kdRqMb+JFbhppP69aftI2KJVGe7l3FdWuOkpt
GBwJj7MOm1a7t0UM3i77p4QUiEulqvsMRnuXgrWGWBWAfAokIVktI/6TOsHADiH8
JZlpkonHSpa7H9f+3Tnrld4Mqimz0LnSEx/1eFQWxnxtZ1VGaxtLx5kU5NUPcyVu
1eDmLx9fu78N21l11bCjeYuPQIioGIxeVaLVRjfs7AiggoDP++tcGWUwybGm9od1
n9xVkccyVcyAQdjFDuB54aIekvarAYBn7hLluGaisIOYbJe1vCDEIpWVfiFNbUhD
/RtFprn1rJbrifa2sdCsFQemZZP2eWjYqBcHBCZreQPRcxNSgX9TT2KfBVaCAQLM
i+scX1tedpTOEO+byInObgqjrFA0djsgTAX+nnI5gR1TueUgx53bmYimqPvH5G8k
VPMqNuo7jArhJp3mjgIMWFiAPPjL/rBGaijrBprcvmaVxxHNF8c9JARFBhjeJ31B
PObv0/mRg8JwSRMXiebJ7B39vPtdZwpiV46v5/V5iNkIG/9dNXh18UWnj4Tan9lt
pVQ+Nhmv/m2gbX8fZzIyDzq1glRYbF5mKFQSrzKZ5J7qstnWNMsEw1kBuugG9x5e
cuyqKK5wTrEm3YbDNjhvqh6SMO28bcpxCNIUo5rSl2wIsKxognCLQdF8o2pPcflf
wqGcSyNSif0DmgQP11Q/p7LDA+ueZ0cilFN1TFtVQ2+N/Vv3464YuTgO0mJnulhX
tReeirLNSGI1KULZ9HTu2Ra8GL4cXAG+DtoNfTudFS0eIXlFXeCdkQuGjerWtgcs
DFtAQ8k9MsCsSxm/3G9e6yZ1ixg4Jd58zNQh6BAiRym3WoumPl3SgQVToWHL6b3N
HF3etz/EHPQG/ZFxzJHBXSrRwxkqN2L78mbZKstuGpaYsclYu7K+5BjSkRIhtygu
YmdIxHjIv1bB12NvVkNCm+w5MdI53zPLLtHcj9mloEp9Pbjm+5K/e5qIYOKEZDbK
SpJyKBbkftPJ6cwfj9C5x2F0y/VA4vSyRls8bt0GarUV8kv6/rYKLTCBjjSMvgAF
p8SCikQDymvq8lSDja3NREsfhndepqmcLsV2V9mzHR+RrhQCV7p9v+Y5jICuXjnv
CxmSfF04PAd5uI+bkPZJDIFLZ1eeui2u6oI5zAwev6+amj/9PInhm0320K2sr/dy
jTDN+6u+EHLsg6VRVuJXZc/VNbpOE4blIkJ3tycQ030Yhj1HHiaDudlnMdMn/9MK
HktJ0U35hQ+39RZwJLqVTLKAPm6FYtaomr5t+NvCgcx9hbInBNR7WsMVcdfXH8xm
7ZI7zZuQinCdDDzqMYhFIPEghWB0RLgxUBQEaRLlc9h7rabaVjaJ0t764d0/13pO
cJHVOi8BgKGCTXVz30k1CJKgJC2duqmQRYow0qaEcJv7WYUVg8jnWeekeH9hjqfT
cnwZpVyiMfrLWKVOrkMpJCxaa7QWluNp7UVF3uiWqlEvDD8YZBRXhNb+Z6ECFVy+
dv0mfKwNz7hwfuQoZ8ZzbMmI1lOs9ZpRFP87cpXV2CFEXtqSAFeUo5eXK+Gnv+2h
FnQswFoleUvZxAl1v+HSPuaRUpzU7RUXyLsPr1sj0wMBrC7aXMiQH9XWiGm/21uK
S+wrZ0wgRj1AJdWJEiRY0VSxNnE8Vq0YuQZCkHPrdOF6G0sGs1JViYuOKqY1P52+
PTlI3JOGNr/TwMiATvncwpM/me5KXtzX3j1fRDskTMuTy/NftfOU6Lo7ytRTpuc6
LrwfxPwCkz61qMfjvfgKoSe4xCAodHG45pgEQ2CAFL5PzltnoD/UhmY/4e/TAuk7
wfIHm7xUjrUaioWcrdngxY4NKzkzRp7a7VL5EmRSVH1vxv4bqt3/Fgrzeau2QJvE
VO0yrEOHsk3F4KQ8BkMefi6jwe9bEfpBmfcrVshOulcWu/yPPgV3t+UlPeb7S391
hIb+o7nPsUVbGmY8j6cv4vhW5EU7BpnAN+ANaHvP0qjBGPVunMihWc1y8Soocgll
docTljU5As0so9SRJ19jmlAqZYuYTOdTzlK1eRYJ/K8VY/i3ifbuPHg2kcg4fwRo
qeouIjv1z7dhICzdTNt5qHwP0dzuLqPTFHnc3x7PW05fbIFqvLs6E5yE2PRZYIxY
oETh2rA/9twE5pY/3VmiAxxFkeeAtjSuw7/jN4neTyycHg5enGXxfrht0/0lPK9j
r2WIC3XhF/4WDpuMEklPflmocbG79jv8uNy3+C5aoEDkw+BcpVS2TD7v2+XynVTE
4Jwnjc9YKYt4A+kA9oDEt1Xf+BarWVBuhLyRTMDP4K2CCLWJF+AeFG9NMSHdNV9H
tOVkPdMoMkHY4vibEmDoT/K54XUFrIfFQnfwpzUTf4KcH2GLPJseFCnjGl38p5ky
3YcTGK2rBHB/r4lVmbyNV5/qMfV3Xe7MtHVgHycPoSNikMgdps9jz7hFNI9ciDa5
8AQ/w7McyuWOJGQNMz109QRqJGPeSq0zYTxpeFvStbtz3DydCWtw0HQb7VXjr4+O
fAvRan35qcYnQzY5hf0xqQEfgKko8q9Rf6NGlhs22RcTuLeNmZ0O/4Ht/q5+16Wx
PsRRY+lN1yiBMKTibSCQ990NvULcXSJcoT/kshzmX5f2v+tUuTRkB4ldsi2De3jy
SIdSmwuxxkNKGkgv5kK7LxMguNmz68vr3p7iEEAwoALKjjJKNW4zw1p54Rj9wSbY
K2OVHER5wqL3aYfC/WzKqtgEm/fxvyDUEHWAlCpjdvv2MoyX0sHDuq+TvrcCkldw
/ZtLLF2gGY0NXlP4VHY/3Pk52NjCJWAdEU1N3X5zUwd37e988N7qQ2f9rwrbrJ82
BmWaBrsgh4tEIoX6ME2gUwhCNpyENE6+FbGa217QEMkHavZUEEUtClY8Ni0J3m7+
LkHPiRTvKtL2JLm3dIdmj9V3ZfCDNbSER0I2UUZuHv7rM9HgLkk3hBLlvoG5dToX
6cnmMO+dOk/ofENGDP4NDzO4U1FbXi+f3qKHaiyF4ORLYhEvgZfXoZU4xMSzinSP
AEotjocuM9zCGVltWRcRnxfCvrRvgRd6KBWuhzpIPiVcG8m2gxJd4ywvJTsO84lk
wPBqaWJ/O/Tx5F9mp8BWVgNW/hD1unk6UpJOcdK68fY5DpRKuiUqIX+6UjAWqsYI
Az6XKRJpkUaPuhtIbUfUiTNRtldUemorzXgxvuEBQzl13rnjNxCZWD0WknG+61Qh
Ewx+YCKYxLhce26hLvCsTAhNcj3ViRC7k0EWTuBV7VeGcgv5Od8O+8+vbuFFJoRT
6/sHA4aiBZeY7HN0n7Y7MAL81pt99m5p18qHOfdXUNCvwLzQJfBwX+kOEN0KVHNl
gtKqgJ1E5YfuOw1te2FDeX9/uCnD5l9pWDXvlTARTZzuy0kt37aC04FKuOZVvMyV
Mb2zc2qgFDsLQFmXIsg7LqYYEOzDeqV3G1nkpy+CNa6+a6NW2Nyc2LXx+QppRjbG
xn697xzC2kDNrWY2pUUI1f0Pwc6w1i6DCw9To7otvR52tCnxMm/QPmbQbcE5qM7t
TSuvjHdd24BpXfcXYqouqqNsa/RTL92KMcPHvW+SoFjtRck4QVxzu/FEzRjZWyE4
kiXGbis03t57VDqe/YY7/Ntn6oYKrtTLlI/pNj6rEIunORDb3ovb0WSDrpa7d1LI
ZN18qL4vRlLl4aiavkTA04LXNIW/jKWgBCjCCKUvkmOfqt4ZGDX5dv++tPbFMLmQ
NI6JbZfgnd3p340xDuglrSoyZcDIPCzg5E2Or81FAgltBehpxhjKUuAL2BlhYei/
/oDkxN1SVoAoqq3APXr78GAXpdwRKbdKnwoeUSu2APzkmKeFZZfHBj/klhmWJCrR
x97oV0psZMqylFaGCAQIAEGoMMHwP+xpNFflr6wkBl69jlOH6cI75+YItBriyGNB
+NYxS+pDBW82BSx353KSQs8q9oUXdi0860UBejdLIyJ+KU0NtasT+/LkQKEwYVh8
LZ09TUu8q5HoXOYONjaxEw9/Zd2cdvxQ3OlR0QCnapH09P/IGhCpjP7kox7bM+0o
TLT1vZgk6rUiRCxoC+ALsIeXyNBMDINozS9LzMFpzhWUaY1if7fi0cwWzud3WPtN
ycl6q/lTG3D3VOm2POZelIdbMxYMfzz2GuI0VbkPJtDgfo279XNG5lAQX60Y1i8c
IHY/k9PmtgYdhc7s4eB3r9tA8WBQOIIeeF/7Eb+bdNDqqRToowX91lZIKH4pSbIT
8bENeO8NflzW45S2P7dUggRjHZ0ebLoOgpvQMlriq3utVUixkz9xDG5OUM5lZggQ
jTQoKYkqZWqYFTYf4/Sg/1yXiHmQyLRLnjZseJNQeC/J08houl0ChZ9MiPdik78P
sUa/RNEs8cUjS6Qkq+juaI5Fzhq0uVh5ffFHWJe7hjmCDrXeq79+HglNchfjg9B1
zrwMMIqId48WMIdIzt79ja4WrE1iQ+/zi65k/iVXH4Bdad7V2B5VRDor54MqA7ak
Cb6RiUz0H9h6OkYLpmL5gEpYOQtGU83X7tHTm2GXALWIr6v68JQgGiaUFST7HoBu
A75Nr9Vg8PTJr5dntDIphdzovmjktslZme9zthVGVmjw3Vkd1CKwQaW49rl/CB3Q
RYGCHATTG5EWObY0OA8HlCxgL5rGClHHB6guH8ONQ2EVlurE6ybnoi4r8Xrr11tX
IY2XMnqkLPzQaoZZufgKo1GHPUp9/bGoY/taDfF2VzS23vYOu5IdioW/aoYV6LH1
ZNfIFWTSeWE9c//57PcYRjOliYwVYT+8u7DS68l9nA4n3NjeABAVnDINLY/cXjuJ
vnyQ162kmgXtHhRdKJEqSDZMVgBS4G7fCq9bT8caKfnfS0zSTehu9clL6e/M9ZV4
LEr0c1mPEOFp3vW1snjlIg7wgWtZKJzrxPAhcMSGC882rDDptdemjFtd3oKYORrS
HoxYf5noTvQDOoUOU3g+zN38uKLWbHN7+FswqDqMSv/df8p5Ge4fCEM0gfOrtTtX
FduMDgEEFC3E8lrPdMfJETOEYbafwUM3UyNZIPZVzby+5IbJrKm67rSgKkp9mQau
8Rdcw2OYM9CqaUnLyqcN1YRGgswCLYgGfQVEQUaFfHDICY6hVwHKXxPfvfvkilIu
uSnxMVqSFG/xpdXMA9zrcrTZg6VZNc+2XBz3h8z6qgPjtn6rBiKAHdCU7AZXWKMe
duXHZcQmBjTXtBAwjlew3f4tT5TD54ahleQC8j+4gldIojNUYyfPxGvyU46VJbi3
JdzSfngU+DZLMUzjhUg+pPjK8vMzy1XpivgjGdnDn7242AZBjGbaJ8EeAb1/jdUT
hagVsDaM01TWv2jP63v8HNZzqpDhQNqFv76naGt1CeQT/aNSjF0qv1Pt/jf2fpwp
Pdqs0Vcwq/QyFoYEKvD17DttPYd68fvRZArci3JJm6m0PWLgElh6wYQev27Ztkn5
+ZJboeNCkhgzHLG0wpszjq0eaHqsg0a7q0cJyDlA/RJln62O5f+Q4QNgLkd23Wu0
9NFtz5ECzFpAXOFarqe/U/j25/pvPF47HS6+GFEEBwZxeG9XBAgiQEVL3Ms22U7A
On/Vl2jo986FDJcyS0EyAzkrtRWD8COHXAnbxYebKR4xNy8rYLPQEITgUYTUrA8d
Eo+l392B1D7C5R/tgyWHoso09NhuHiElF0JUsUzEyEbhFtRvlsCJM/31YlWQekJO
l0yH1SKhFEIZCkSFEeGykF/23n9E5XhOiUbhllKBe1KGIBRZrqw5jKD7cfZwRjWh
jMDr/legNgbQQbAuwFnDPRgj7xvIfB6ImJog28r3N98ruIRKtn5rNKtTWaiDrQMD
YYoWs/cUVOZdwnziLpv/xw0UbzPi+LUQPO7Q/izt/eErTgUAlTZRryNKQuUh9GCQ
cv8oEkxoRmt2zqFdsDS0rAR49aA94kXWn5fEaT3CIapw9okzMvYn3YthDUmheeUO
BExcHJdGU9PBcrW7q6kcgv10DLP8qQEanI8jk55hy+leggkjw+5Cs3AlCd+FGv0V
U3o7vqVZNztjoXTuHwHaw9Kw/pimj3PsqgFRADgOUUJ3UAxqvmiW6xnZJXWdPrdV
Z3uE7I5qrN81NXr9tLt+I3RndCgydYySjccY1XfyaT1CF7soWXqvmbG0o6bacQdU
V5YaCN57dRbnusXO1juYgQH+k/v8wmvE5vTqEiWbbep9gXViFBrSHND+9y8LfqyM
yquHkBTSj8cdZBGk1r1bHEEoGEsi81tPHen8UQCEeKqnCacNO3FzVZt7i8myh6TI
ySw5VzHNxctNfIeZF66g4J8EF3hJppH/oPngf9MnPzyIxaK+cxiNiivNlUWZqWNY
kMkEj8Spq3zxUA6GzNZymbkbLgbgbSmJJNiTqUQ+4kcv0HKX8ktiJN1annbR1ywP
wF0Kmkdkl4mVkm5JIILMAxYAGUDxWEaynFHR8FyJ4a5nKO5npvJwrJooKW9TtgON
k4SJc3f62NAMxjtTz/rQPOaj4aELFb9NnwbHlbNxCvLdQXgOQ8qyncrxG+wigmAq
bNERD3BnOOD0pmvRyqXdtUc/jg2s5g9eH1PODWkLca7bOSGn5X3865gT1euqceiG
Vp9sj3YLyuZbONIoJeg983iTRc1rnuCNsNkybwa89uVwKCVqwnEC8UWoTaaN7Lg0
BFA7P4knrr9RhVDUGEYlIZb49dUbJzDyx+YOXlEqGTD0tfQfD++8DSTxc4JhmisG
/iAGm02ITK3nVumNV86Z3z87+1VtRnWXhe7kwO9UjhJMdYfnu1WJfj4nayRp1M9R
KWDibwcB2y1zLa1QTZqSU3Nvp+9uIYuxwXhSFhlLrONde25p24+A54rl9zIJ1+2Q
u7kAFy2rWJBGns8Vh652S0oXTpypFntPRMCvxX2ObsfIGkbUAPLvZ8xCcEXt6cSB
q7xkG9tsQsFb9LanULDbjHlLDvvGD+vWJ4rQKg4friHH4aeRE+j8Ha44X1X9YJH4
EbzFwFDTKASLESJv45K1wgYAMJ0I2VjYiTzmO7ds/FrGTdMcmEpD1Ie1c5Izklr0
2CM9W5L69wNBMX3PuPijhJd+AguSrOWxk7uPc28Vt+rdhUAFWly4grtE1xXFu1dw
onl9Vi0zPqvfXYVJbAaT7DjBclZSiD+wp5vRvRQyXe31lA7VvayeOKBaMpnqyVxw
F09k6ph8SRJXYj3uAFcxRMe3WZ4ZDXA7NynVIAGKMGzVWkaK7bgW0J+xOugp9KY0
hti+1vb0doLlwCHuaSDpAuBcHtnXA4gF6KztYPCR3CK//4a4ent2TaeUB7McZ8Lp
Ph9t9fNmAtclsRoGCCm/Y79qXmLJHOUVMU+wqgJcDHUw7WoWUMhXAWaIdB5x9I8Q
WokT/dLXblyRXjwOgzyJBomXbdGZrHz+pSJIr8o/2tuvsX7KJqrjk2jTj3Pjgk66
2tDnU6oAA/4UqHF74QoKQ9eDZMOs8JLjI+yLk4dIirJxkx+sseRrCS6uNi0MBQl9
bGPggIS8oenLqxOKOpP6KjLFmxKQge5oDe3zCfh0ObXRnIm5jFANkTPCl77E5lhY
pAKEtu1RmKbhRq6IbDR1HFCHUPsmflDz0U4aKGiD6oxROP7Zwv2Gp5c1hq96shdt
SW56G4yfejXxU7nnxFX2a2badZzg33sRYCodwEktj3VDAj+uxfxI0qj9gmhT4wGp
rqJLeqtf4AemGDcCf3PQX51aaiWWYEH8GDErfEBoYl3MQy7tIAwPpXh38Hu9G/hk
3UJhmYGXbrW0Z9fl63bSFqUXWhLs1iNxEYYes0IaHIh9ePUagNQwXnRAxXiCSDXd
5LzURDr1U1ADZHDKh6+2TBfUMPGRJh33oLyM2L5N98gVSV+RawWscbP84ZXyQwPJ
x/Hheq/zhXzw4jhkGHabJ/zwMHwinYGySzXZUpflsvqjx57JXOMT+Udi3Kn4WOwJ
cB0a3k3VLbRPo8svfDVLF4FT6FHxu0/FpIJieXOeQJcgXH4hDY1jXF6qYHlW51Tr
eTzsjDP2kgai+2pmRd+codKnhEikepucf711v4bpEbYnTyCrn/9k223uEPbLkl/S
1WB53eX7WtpKZ+Mm9bJZmq3+FFLI6OZq4hXoagG5HSSkOoLJQYDWT8LBpA6CMyOl
3kPc+iwnC+NfewA48d+ThJ04Yurt1yGMc97DskuFdzlB3uyCVWjh4xnm2M0BNzOd
UsNhjl08lc8Bd8X5zvP8vJz5XS+Et99+WgrUd0XSvtnmAqyShXCGcwtaDMMIVtle
H3pjAFTUhCG8hYBsinYm/LPuNXPnJZe9p2KpuVwXIsW5IXgWInN6iR4xPX0rGdKH
t80fGw0qkw8vruAmjfERGePsj7/qCCOELpvAHcfwyK0gEva3qCYfmhKrz76nkhTo
XhbIzYxpxqVf44M/8X3BFhkV9xVXZyDJbP1NVMg8nMTabZDI7BJHyk8ore3655r4
UpWSZCigueeG8HJ+zeMapKZW8BB9abVlxXPveiozJCZXOoOTsMfk3SBY5vYr54sw
Sv4RAmi0tD0vtqJr8jJjEVMcM7OTTU/9yYOyXeCtvZo4fNquaNwHWq/CSYVq2Z9c
M0yoCw2D7bzwv8z7gLz7Lix4KHUGEkLgaQhDpD1yEFEeY+FZ8Z2hdgMB6HTFOcmh
vIo/HnSuEmUcpw+1M8OKt4AE8F0xNUTx/Rxq29q7YubnzwjNSvhG933yNCowJ10W
c/NTbrAtnGUK6gjjIlksSuds5E/1qm4OAKqab+Dj17asRpALyKAx6Z9zE/gRVyhb
5cAfsGQwghqd3ks8K646TperY1hnaqlqnl2hEzYXCuqF0QQVipBu+Jjf1yYjrGf0
SkRij1NeKIHadfbd/KgfrpCd1IadYnuo/xLCj72JgWy9h6LX9FUHi/gQvgDNMukG
65L1CJvDkWZ/Gwavk7p1A/XInRB2mjWA6jcRPhd7qCbz8zW7V6CzXQXdMoUj5hLM
8T2HBZDkFE85Qv3+mCFVD9DDh4T4LJF7mqdBLCCF4hnjmSMUBJ9jRZKhDT4q7gd6
znfVxGXLTATVWyH6VPZ0HQQZ27ScioDJjbb1DxnR9PIGaafseq5HsZJz8Wtc+qw+
Qs+GAt0jQ6JTWfxg1xom8VTnJPROzAomw658WB93NhwchnWGawwxwX8fG3m0fVOe
CzddFSMP8yUg0bbgINzBye8itpT5XBGsQqACPILVaJkflAQDwH8h2pJah1gHBlLr
pCwYr2XzVt0vDgotC8xWpPljmo68/Yv5tufwsZEKrLDYtQWxxX3EDFvkLiF+iJHd
nHRTXVVo87d4hArQgDoiIuav8RiLBYX/Ll8WiszV0N5DVW1b9XF7wAV8/zJY+Fp6
nxipg7McTV3XGK2SGlXw3pcSyo4aX/l9M5OwZIYgiuyscqAXDGjFdEWUPMExQXAx
sLD6/YxasF/Cd2QKe//VvuCBPDOoczM5rrpkmPvHciGrw5IQc0rOiLWuO0VFNM3+
n0a6hbWjBTcQlC8UwL4a8I3A2988OH//4/wH01OuTKGGeIOUTHXcE38cO05ILOep
xOiZcDsxn1sRoJkt68HuyegbkM077ls0H4tBpQk8pL4NizYFlQtsiQ1AvzMMUNTx
5N7mW6Gj/AVOIx7YRAnK/4tcG4QGBtnhV91S/ypxn3nqrp3A7umcZLwW4hSZ1i3R
UnTzITQOYYgL386WIcSy6U54HjQJjDr+iVxZmqUMui8Wg56hMb75HZfd6oIZGuqg
JjoCYxh5XmzmMsa4jjT2LJH55ND398gFNcJzR7TMas87t+eahlggvCOBy1Oz2cOY
aixY8l6VJrSOvfoRPRsmwL86N4QOUG9MOddIFMCFByouaLxWcZDhwDn/Sdvg7sh5
ESx5tPR+WANrkoe+OqjAUOqRBcEORbUodSpQRySd0sJzi/8PdrLSpTxTryLMtztc
eADNQnvnkyDDQI1UVL2WC8qPQDOK81Cm21zWWwo90tVLVSnaVIKgbeFeVw41T1x1
+ut4bPzsAAPkEtUtjc3ozWMhXH1LQQyF3qWeSL27RUup6YdCZ8ukcvEsdl1CwxKk
qNvMlSz9NSvKdG0gzTJ6i4ijS4XInRNQh4iWxmpEe4ufGhj3cCJ0dWyyA1tODHKC
Hyns5ijMGZrCLdQ4VY70pmbR6juW51xSuJcOcebcIhO7s817c0y7jPBQKNLgOMy1
JfpyJs1spP9Cm7fkN2vicKiATJ5bZ8OFW3GTGlOAe6vG/eMvH9obuU3jwOpSSWya
8GRf3/z9P+eFooquGyMiDnrle2O+9HRymNWthTS80nm08Kvs2XH/tSpfHZ786SB8
0DKwR9MyiCqHMsuMNPxgg2iQ7XnVFoB8RCInXTu50E2E+h10zqS3/HSdJwpzfKLH
J9SpelFkHEnAB3Jx61Az4kt0S7EZaS4SRdZL000pQoUC8z3qzMQtHmdyZZ+0reQF
Mk9qm2p504wBnde17tXYpBImKGP1jSyVZ0j4PFun8WC7RyGdNzMyPc9rYRm/ZTqR
djLetCawjHpdxXC8uSuF5A1TPl2jNkapNtJCaGuTdY7DAMQ+vMt/ipEWkamP4bLt
hZibqBcavB7x/L/ZEVXRVltRs9L5NMeqWBBNHb+ZM5gfI9l4YscDAQRAaWHcIWkH
dcVzW6P46+ymhMO5rlZCRjRxK468wqnQkfDDFJpysMx1jRWzXqoEOReHL2zSSrWh
raEyJRvDeHPqDuVr81l40hlX/Ixp+bqvAo5UnI/sodC3pMYE/1y0LeVVcBLKsxj5
Nzg2xCbpp+1BkULbqaUjDYsCK0vLPfxFhnk/bVFFp4hhQ8brl2mCvJTn/4owlhxW
CE8bcRcXDscKwXxIZNJWhdQ9+374LU5u1htDQZube2dNu+1MifX2VFVejkTmUl9C
jXEbGLFbBfh1OSOW/w3CsWAoHjNwryqSGfTUlyzjG/S+kRXnxjy3jEjHEoJfabQL
310mACOj85ipMr8Ryrwsnet1Eb4lioM7vSB+cHKhRs1By+7of7VvBE6EBgS8vPoh
BQfkat0kczzfuISfmfJuy3JXzozcz6Xvc7lV2NvVVd5iwc+0JWBM1fD0Mi5NRccS
yCHmb/yRcVlRd0TBTi3FyqPbcdTXYaZ3aJboMxlXuslcV/qyqkn4fQSaWsJxETZs
y57AytaNvNadJWnwV3LfhJDSp57tObbBQb0ym0HMw2xe7OFqudgilUo/ley1X1U0
5ITQWw8IXOpKT3L/SX2uC+G9JEOoFR6kZDuyguhbcUl0sWyH4oQ59uNPOGe/KnJ2
KHKFKjYFMXMWxR+N5/hsCCugpzrOyqINeJZ4xdthhyUL8bwDKn4pklQiXQe7P8lC
7+ASGKe4ipQKXJE3P5ZN1NlJibof4blT2QBLVg2kWxxcw8H4qocP1nve/rhn4QcY
mKwPg5J0KP7FKjzPgbRLbp9PmjEPELzDoAQ8nlybFXmKuE/0qkAHykNO66MoD/i4
u7c6gFRZmcz60BmNre4I6myApsFgMAOswWR0WU6LJhj5gOtTJqG8gzUcA3ayGLFR
TNgEoDO4blHYvTp0+XEmvmR9b44S8VnoWXlTTvk6raTTFOZpoSW3BkYD/ORCIpq3
U6UCPhW/lQ4xekgdo0ixDvLSoNOBGh8NBSDU45ODi8FOgId/OQOs9pjzoy0/o7Ue
kKBIlrQ5uDtaNHVXNPqmdqdkYY75kaNzT6YwOHQS/5GGXv3mFM6wAL273yfKaK/R
3G9Gq5dKYYRmL22csskjXZkScOhYlcIqNFQWdiRGJCBE+xydn7cEkO4O6AL5/RdD
ghU1r6Pw7nnjwr4RJ2N1X1vLzCpJtRLxkK44yBawJi4l5sEHJ4VJxPy4DACpPXsE
8jz7P46kfbE3GW/ZxAZenaOnnvFg/GonJXOWXX0uOaTBfSC4Hzt4LMi+1N3ggRu/
KPOTZyokTaKDOtcO3dPFltAT+qDcVu4wP7+RaBrffohWS1sPWV39OdiLjessCprv
V9fa4xllLCpd1gPGFA7RRRFYZ061O6HW4tSu0CQJ/caopgascZd70V0fKLYraxjc
rCUT3jBbUPaCuwEqtKZmE18SXpuITzV0Gx+XRNEs4da3AOOU9iWG4Ch9k74k9RwA
na0WYCORVtOnzu2nLm089Mcg+ArIWFrjMH09zyq3hU2ZKWpt3+elOGJuXTNq8g7w
l3vt34NJt7JW5awA+ZjLjur0z7befnIhR92VjRboVAYC+G31znApvIHfcOmtLTE9
budutKoYZOHX7BEySH+ozHjV/7yMmr+NBQWAfnfLfvgpAnM3eJ52vJTib9IUsiUJ
r6KTQK7w7EwOreJufxr9WkfK86HfFsiCAaaylZy+ncbRbUxOLwjhMRe9LabMN13A
hgCqxN1P2wYV02PmsEP+3wMblOQQtxyHNM/XQjb0hNFUVhe1wx+19TkIABQN7NuO
tQolPz7g7uRrk5vS4YXQMiud5Qdai5+Bqyf+FlUgBl3+Md75qiLWIesgIONOrJPj
Xa9u4rKW5KsmUFe68ydMUFeP9AmeK3Cn2t/TWxBcjnH6QMM5cCJa0BwaKGEpRBcG
s9NbjxFYqJxaYzSGbcyoOZAdOQehsGm0kvPey7UrDTUBk132pttAauSQbPe3lgMs
Ex9mu1rPn8OHyed53l0fQyEMZkcW/ptSQVQToYbN4SJXnF3dyXtsuWGiJ5L2Kla5
Z3r96NmoUNQ9ev9ifv2U4ObukD7l13SBXM6pF6ElvH57hfySu8SAOkv6zXiWKOis
sTK3d6BKlj+YoHKlH2yQKL+gez+NJcz91BmfWvpdNodvNAeOZlr7ELHQUMnSZSj1
Mo7trbuxV90/14SZRTuImAoE/1XrBbiyBNc+1BBQnE3cJe6Fszg95AezBIjDV8wj
D+h9d3iZSXTe4KHqCsbhDBE/tSVI8RlLWH+b7MI/OgEUfVaN9CRNNm4bEugJ+hwd
jEIb9cIAV6Tpecm8WRa+/3V7V7/ausznlo24e9ZNAWmu49o3hXqlaKGKEUSGiOs1
Ut8S+TTGSNydhffsUT8rR6pObs56Q5XBBw37uDDihluC3nIL/9wYvflwEPo4JDzD
1zYbUuLvpQgQlizqXVk+FbqAGjNKIQfhMpGklEPliAzmbW6wLlMVvaOPP4HzJs8t
7F+AtZsXlNqwatgLT9d/ZAaK1few8Ajk7T2sd39rbIORGbdtsD6OBsaZQMta/wOW
OeWq5GppUdEKahWXaYAQy1ocIXuj+kJwZN3ZVMKpDsqzOUWT0iZb24s9Ko9PUFZv
khmWpChemQMsTcdX6sYTb5uSZolSDUbfWZyTSbhs9Ul5RgtcdoVV/yZIKMi2mMjU
6LZkONJ9F2uhPblYBRYiHTe7BMijyE7oBcbk9nwhuNWCwXcYt/SeOStlAgzR0vVo
JOOnoIhbkEjSpxPxCjwX+DgbT5Hn3auLQeYKESznud2LTToCnQxoEfL2Ac7twTmF
gmDn4vT5bRSTvLWsEMntCOKQqHZgWUu0DLU+OkDthnssw5KVEraEh82YZYtKAQn4
PSpTaonvI3Fl7YWkG7uTe/sV6qQoqXWw6iBwL377JOEgY3z7pApsKMzfOo7pgvjJ
qQ6TVp6phK9oC8ashpLtvFfMLelKj5RvdY9TtbX8iORb3xgpR00ZKw5wjvSeqnUn
oMuMr8RRpej/vCMdVtkOu/r8SWPUf400PsPmXqiieVloFgZ+Uw8wWmoBz2986sim
N1+icnDDldvAIcLLPp7sNUEZc9m32R5UrCRmNjgbnWo4QGcynM5DNXyfAMvp2QgJ
THXNzSnqUZWu5dDkhVUHK2xg+7+PgjlwRqSD8m6ddW1WrBsx5b6g1LZjzJfxuTYS
jvf4afp5g4TKVgFHxc2LhtFc0wF58dM0VTeXpRW4Y1nWlrXsu/J6NH0NIC0+Kzcz
9hGRfh2jlsCmg0LUBf9g2rdG2ZdFXAjpk/677v1qZ8UtEom1Gw5sw+sl40ZZt7Gy
9HhbKwFAjss8saTAHTDwv3ZMUx+Au3PSza3jA3vMFZlBVGGF+b6xjshbCwHaSlX0
4rn6osA7NvkGkvRMb/Ltkn1PQjRXmAB3mcE+DdiTJssELZj+MQkm0dH5qfRkO02Y
5Fl1W9HeS4m4QZAmcpi2ZAGpw5H5AWtY2QkMKrB1xtq9pXRUXdItgRwemgPma0af
X/SfmwGy+CvPR5a3Ux1X9kH4BBJzaP72DSXMX82VtEjhO2POjl4uyr8eLyur0LkI
aMtyHBxa1H+rZMdzTIJXyI+kxZ3k3RLMkJgXQb+Hs2geiAgz03nb44vE8dgppyF9
DA+f4+zWEew9+Bfu6pRhf0DqcKfEDWA+nMVxWZWKnqe42tLf9N/n0U3LAeFH9JX3
Rx7RPZQQIqX8txobuw7bZHzfLj2JMEcNvQwrC+ofzh6oyPdVLixXG5IMUd1H7R6v
wxsEadq5FBTc0qePBkO6mPoMyn/JlwD6ctKXjP5KhKyEqEuXPC/B8doNWvy3lYM+
EOi3+ssamSfyts5Xe8DtVqHoremj/j5YvSYTqpsqcDzpSLu98KN3C7yfbCSbO4wT
coBBIIMeR5xswu2pPxzLrBPtN1YssXQG14p5T7oU22u5eGQMn3/WV/FFk+2AIR5B
JiRVGIRIbsxjDlqCzoHgZTeaGTks6DjTVHSeiM5IhcLEPIFeaJNxatxTpqEobkPA
JOC7h6Mwbl4JaIdwHKvMo5QQSN3g8Cm+MTMBNzGoXT4pl3M7Szjt327Nyo3yB46A
85l8MEPPWHbHedNmD+q3DTYRBpXwd/BwjnWZm/PXB/h6R6novSa0XMYcYHnwY968
jBkT0ec0/M00pxC4B+d5E5euy/b7tL0ZqRTHyfqzOm6Kt0mmVHwRYzMZosieHCkj
woi0U9jfiNeFfCs2gP5tN82yc64ZcvGrg0S+zexgII8xyXrexwdtmOwsIglV6Uv4
cRlolowmS8p/sPIy79/qXfd9yW5193r/XYMqZhUA0wr/9nUx1i0HI4ybOyV8B8MY
cdJS2/jzkxeat+0iQzuUn+QmFqecmFoCxSdO9+Jc6D19x+KrvjlH0OESKB3VuEZe
b7V/nlETcH5HNfCserAKKG4O4LCMzoPYOWBZPbQOBCJHpaKzL2yeQSPJy09Q9Nvw
DY10b/55kpoOBDWCPByc2MqnKVWprbz6HZYiOojP4trFvqLRopHQ3CLVXy4ZnaT9
I0kVyvUcUk48fG00ZPeh7JKqRPz/H5DVb2UVW/Kaq1E2SIXqtLgsSpOH+sTbk5wV
pUGPvjOTTmBEfqANLHi37zQVQuVB2MUSl8rh4b4RSw4EleqkU1C7vXD9jlDKRJZm
cwPy1RHR8N1vAy/ZdgXetq9EYsn6PrYfAqDY6j/FHY1U1Q7DXCb4m7M613rSz26h
rQRwN9PbgIGnKjU/JwW1i/MM0uwRLU0kVBD2Ml7MBEzCv+oLOkKS7T3W3rbA9dm1
A4MnVy2witJnE7IEyCa0OghGZIhio+dSuWPRdCsBXB+oXvj066omYGU7KYY/0Zb4
iIarLf5UNleVG+n7erWgnKCBTkHV2iTtXEkU4avQ/yktu5TVW3e1cSdFUFRQU95J
LnCLifVhESo2tFWcGuHm5WjBLMPVe4VorZIxJK3PpQReSs+pq1jklKtGODbYd0+D
rKM2xFfkJBP/ZOzYz6kCwCIlFvcSjm4Pd1y7KPtYVmNcoSfmAqXPFJ1wsbKXIP1K
gvulJuCNgWayZj4wnBXpvx71a3ed+QDiKHC62L5knkgRk4zwzDFW0WXV9eUMfeYf
EIBEL+CU3++BggH7HL0fwDPKlUsK2JcovXWkdTYyqrGJlUwvTECi5G0nlVHDfIEE
LStxSZLHlFtP2j1f2hPwILKGb51eMsm+6PqT6OFoQv95i4FSB3miEEYbWqpG7dHk
J+v0CWSTXnUI8o3liAQRSidaDSe7/JwRgeKs/INtFPgw+Rvv4uYtJDU8AkTAoFmr
tNC0hFwUfVy1/9aHp2kCAMSrpmhwxo3/ZCffHIE7ujH7T5sRirxp51szeQGhpnuc
VqzJ7vhgJQwk3m248ei1LQlGYsTkpk2PgHoAS60rjMXgFmsBvHL25+7R2mWmVevw
NCPk+F2+83GwAOVUyGlKuckfDZijq0EfFYxeWdf9GLCpBfm6l/Xp4ncYOLji7OO6
Uly9PL3lEk9RaqZcE2rBNQgvZVCzDZtxxLqFaIxGVjVy1CbHvh27fUKrUFzGlvaY
iFAY+TsPlMgnE5hweaJPrfIUwc8oVpgFhDRocrRzEVLAZY5NulmFiAMO7Faa2OaU
JK71I9R7W3daDCL1gFcwz2PLwOoTap9NJPt7Mh/WWwhxKfRC9awTci5sCVPeI+l2
JaGTwkWO95dF7vNcet26vepqDo3BywgujFkEsziA20XC2dBbwK7A47vaZu8671j7
PWKglBWxwtGg2IH7c5IVZ2VjH67y4YksHN4v/csM8olF2UCAQ8EKz6zI9eSbMHdA
/gFjtthzwijunc6CtEORG/YJNjj2OJSlQCSvqOTVSXFQ6MxKfaoodMY3WOvhpGpY
UzL0DVNHaxqXDPJTDDmyOUOIISb1OW4ly8KsNp+7o7C180iSzXgr0lnq99fr5DkO
4qVR2c4PqcB+J/Srnchc6BhHNU0OBQLpNC3zYHVjkk/r/pCmw6zIjPK1BL0R3Mq/
y8EeN/FLQHCkfAj71BYHALBOaDhZ/O8j7NcyqKEmWHzMD26DUrpsKIwpf4lGTcf+
HwKnGNx6D2Xj/T+e0GLG/9Fke8A1u16F/XYoifOF6fe4riJY7p2QVKcVsJ3BjYgl
fD5XohUyQJqLkM17Kyj0erstH4T0xwAiFxYgbRnL+zEA4z85b5ePRZ6AF/vNeEIA
i2/lL0YT4h2Q5CXBz3JrcPrz13bhuXvl8npVlZbSuNDiYQqMva/c+45wJDErXtQ1
6nrxDlFhc+MpppxgCY9nvoSf4bgccZAUdjM57Z6KgDtETQ1RjqMojG9BjZX94XM3
xqCWpS/ddLKNonVzUVBUnrpOG7t6GmcJAXAMdvt/zY7k2yX1KDkEY25A7Ed57SLS
h30u3UXN23hV04Y4xSwfwWfM4uZxX5Yw2NI/2E5tGAl6Er9IhMVcKdS5KYmSfWl5
ylyDz6ZHizf9R3SdD8Zt57AOxIdQlJw1ai+r56LGHqEmQV3jqgFzrSQI3yGpGON6
clN7pDuap+YzH3J4OHvle/ComrdtvyivEgJ6vKPIBFDRGH22MxZmb4S1b+BhVqoZ
WrRaLKU87Gy3vrOMWc2uvVNL0YMItLgEP1CDPFMNQHvIzUMjAdju/k4kzoaMJBJj
N2i2vp5w8plAvIljw73SpAyfrK74S4P5MKzASBy47oSfWAVwgfKl+JxrKPBY/Sku
rgqSysIbIM9BcxahXePZ0qigoruaRIBcBJxfLeFud7TocUOjdSflYtkg8OV0k0AV
n9V0jNnVr0cNqfZZI6vLPFpttiHyIWF1XeySCTf/8jkatBBdkOV5HQA4uxX9swqq
Rrbypf84IoD/86+1oQbfsZFhUEMKuxBs/t9+r3RrtM8hNEC+GOENLzewy3pr+FHz
9cPD9NgiDawaFveqXE+2NwB3oQkkHbpBY4vsYsc/9KwcdPIoTtKum+XwJWifBktU
HL+5ki6S4x9N85sOcU9Y9KJrPUI71mfC0g14VlgzABdnPxYkYMev+8rGhIArffGg
rttavYtOCPFG8I/R3zbHTLxlJyR5RpjiAx6e+TtyTGkhXZbqHkbeUFVX1raAE+rk
brwYmKgIzJFXQIRK2D5qu07hCJaRa4+xS4oWvw7ouQpfVtehVWVH1ExSg2tmB70p
BEcFkqlOSO5vBCLB2/frGJ+VhBUNRQ9+zdP8/A8i2woEZvq1AdinTEZcSKKPHKOK
b5FCL0AQb9llK/wGlNdQy7WmuXWghDG5G93Ckctjfv0Rwqgx44fzWBgzjTcF74hF
Mlj04YFfzQbJiCY5UfKCB3TBdesbMvX/648+IiSR5z9RumrekZ/2+32R9mOP50LO
Y1nGwKytm1L/LYf36eucgpvRM3j0R/yhyaHJigI+vB1km6gQbNtydw5F1MpR0n5R
iwVYI9hXc3785fG6CaoxaHbAGRSSAxGgY7m1r5IcbXVLSHbQgilHsm8g4Qa9AJby
sL1oGglfMx6LGrNi7npcXRcCXwZUBp9VC5JNsMsq0JGjAiep3XNnLJrI4UTQcpbs
DvFPGnk8fOJDP1gt0sqW5ur9PRs+nqzjsikepHYpXDl3LaSVkJt0M/bCaM68KisR
GMjdTIdWf5gJcURejicNNL5ooPLzssoPzH9gFgzheOnwV+dh5yAThxjM6hg6KOmA
izwNwu8VRf64IKUhBUGT+dKT3uoK3k1L3W7i1H6zcV9lFTJq6ywTh1qSb750y5g5
IVkTRdV1ynU/2UC1aIsXPJDgwWsYcpA4Fv0vrb6IN/brqRZ8ZY4V1i4mrzU0n1gU
Al0rhaMJioWH5aIYIjfwmuHj1fZ5j8Rv8bJlZh8P9Sf+AIGiCyKsdNUBxwc8+EaS
BlvGLaTnKV5Hv5Xz5Xg6k9RIMuk2qWeH2vKA6STLttJZsDo7Us6Nlv7J2W/LBqiz
8JrA2MkCicrKc8feGOq7/tbvL76q8jjIvNwls0f9YTbF0epl+Ta7+7ItflOQvcWU
BnFTcwWnRj0sxLRhW/mLPAhGkxArIedO9BtzxUFxOTVUraXFCa/K1afsnVRX7r9l
vlH2x81Tm8j0fjFnUHkGlhjJu8hF8JzQJByhsWD+IJOnZhbKe/Fb3rS11xL/MmY+
VgMpiHmQpR6Tjha4yUya21A8GjWtgoSdRRs7yYouRoXzEKV7lnTrj/HHd3aH6oCf
fbakijnZan1i1ur0Mz8ZNEBvFwK7fq3alizpECJ4X7xaNMHCdDFED1RwlCK//XeC
VSFNVtIRboWjUhSAbdvN+jT0lQtrCSw6aKwTlNS9FqkINpUjKHuCN1Y9MUPh/L7g
YgTOacSy9JTa6JTWpSG8V68siPGAAuWGMwtDuscQRHUevFBChPf7kiR6PShxRtGg
2myNs15YarO2OHs0LD6XRvABTRLlbhA3GeW1cgUfziTp9l9mbQhXdQJmIWkHqTwm
Uw0t5fsnN6MJcp++61LnUNpYF4uFz7o0MzEwXmEX4ho+XtZW1X3Twpa41HPU7SlS
LXJR1qrMzKjXTT5QG6COrrd/dahTpwnWOUM0t+s+BaaDJ6WZYbzd7br2BK8R4AwI
WyVriGfrMBS7GwOITkygg+q3eh6kKq0CZ+oaM3hyoxEl/OkoboIFJUi48a3ofTky
+fS4phlpBXrbUdofLVjhVh4dEBdNJZGrdog+BKuHaJD9Bk/NWl4wHTJR3M51/lnw
wQwgmTKaV4ysbFaCEr1r4xBoBSGjlNeYha5NHGd/BWH03DP/ki/jkVcme3VyKiQR
ZWtsu1m39GOwmbOREj2ly4K2lnsNdVM2SN5LPs1L1gYAGNcZjdS1E2De3pdXaKv7
9luSNq+bqDsNCdCir5A48YW+pakT57IsAJAsGd2jutvFmSAHUeow+IIwMnsl+WHp
yxdjiljbIr8T1N8DcsOC+srw0vEtj10zRUj2sYUF4xpgvbPTFRout03ZA6g6EqDW
O2A8C+aMOFBBq8fmw9YILjEnhjaOhIztLqJIIOZVTnGma3zNO6L9HWxIG+tZndTM
utwWhDyVdZHb/m4GEu4TjIkuCmp9wL6hkL7b9tQr4o3v2BDrK11fI0kIjLglTg7H
pSAi21BLIcDhtcXkHmlLNad+Jx75ZqM1Vs0u2iYoTjE7wIaaeoBvLpovCPoqvk39
aB2VhTgX1A5qDO7lnvUCLcxlVjBVfAi/xwMsw1OfQjwQhaxXZs0QojhxnW8nJzPA
7QBQNcLO9C5mTggqOYcJqslSdbJPG3XpvajfAYntq7oW+2Cyqg3BUVfNDBkI8OdU
fjP7aTa1RFEt5k2H+UhyIEYZzrFzSUqbA7R33YFwu1jZOJS+XnqoqChv/BRE9Seb
xt3cahX8kJEAd9tZHCC9jhnI2gYYYzFN3encHm6IhY/KoVSe+HMS3BCXqfUHpOts
8uLfFx8zPBFaCdTLuxneZ5qidbSDT/YG9YcBedQPcBcy1Z99nQWs3yeZ3nEb862m
15KjLOM3T3zFyXu5A2k09h0cdzRgx4BhYfQSnks6zA3Mwcqqtgo6BxWSJ2Jx8bhM
uLlR5Nj/KtK4IkTf9xqYdK/kKTLEBTkuwQVNj6+T9cP093vzsSs6CAoQ93GdadxI
w97+1/+NIAJR+NpYoFZMFW4mS40RkDOO/G7dXxHrZokDvklF2F6UYL/ZJPl+7WA3
DK6ttGRHv9BdA0YTMsUsU/jgde3OZDMD09SeHwGelrNO19qgaK3ypkep/4e8Z9c4
8Zqpmpi+xFCLeJJEXKBSpHK9mkH1qRJsj5LwBxon6TZ/qLMumDfFoTZaY1hi5oH4
umxCXnmqW5N7kWQ2bS83lE929SigteOFNClTXA2O2QdD46zG/FnAh3PM5oqC+BCX
Pz3fwFrtLk6kQvZOz2/edc+p6B3AumXa5+LEiNEHHeCdjIh4GLqVb0ZS8SIao3fD
+pPSbivlnByULcbMjStUC3FmTvAWlp3MoCzL11wyOM0i4QdGqYbc4GGoO4MI2ECJ
HEH44zGMC5XmaLLWPyoe1s8bpRvaO5ZM66cCXcU35f42tu4ytRTA+Gi8hw9cdUVQ
zL9LMRJc0K1MxGDndg7/jpWKmq1HjK3mW8We3sK2H10DSjRPqhipat7T9alx9tUa
S3rUPGUmAN6ri7tjPc6xhmTeB80fW0QbNa+joqqzha5Ci3JYbTvEltzyLCgTepdq
1IaVJU/Ih0oZuTv4bxAQZSmY5tkErVzZN42AOgJAk6fGwlx5rHmfgTqS4oLdFD7n
q/qyXzUEZEhOiz7CM4sH/53mcwb8wdODV/avbY+hmG1b5q53M5trPkFdrAzvi1np
Pth0L16kXy8mEiTmdI5Bkl+OB1Dh8cjmXv4FXPb0oA3isoSFxltAjq9HzR8oJCh/
39BtuBF2d6QzMSLQMZLTK/b7t+23dtI+7lcSkVL/k8Ya1m2QGVYSaNv5x54qJT1O
mVsoyV5IfxekHMCSqFsqKEukjhTtZpGV8dScbCSlZwBN0Xw16n2dvJx+Z6hJdcrZ
H0LaP/VAxgW6vPR4rOxu4sQzhRmxK8dlQNHs9xgM4wH9tLNYO4/pwnWlVotgnVRE
wopBeeHCnP4YJlYEo2KtdM9ynhBiW4FU6JmPKbheUvZnE7WGh60YCdQ5yfPJ3rnj
tKD1+kcDSjaLdzqW6VGvX6rYx7n73+3YSFSho3oVS1rjq4Wjxq2WRBhyqTxMqAFl
g+FZ/PKZoCgfXgr20lEy+EcXz60c8b+WS27xC3ek6gsB/NIr44pDYRCBfN01yAZf
KHNt5VzaIhgBs/VirEHOiYud9keM7i4q4AZSG9mZivjeP0rwLnY2v1gcSD/SrqTF
nX6JaSk7YOXaZU1piLPqbaNjubHV5g6c5/AHDpcPHXY8PFsfaB5ykHnlkLyxa3zI
BYLPqkYWHCQJQUcN2X2QpyGq3ZyBMpjzsHRlcgwdB63m2ethPom0bSqPDRo8wYzv
PZGu2dmnY4TOzDDiQfVLVcysQxGnTx1PjB032pXRwnSCd6kQ3hNcZI2HdQKopl2w
0+vUcIMCiLZd9BpvrSt4t59b7YXk8Y53U9YZytaE0j5kuboF48xUgWGC+J/1+vdw
vxJwJUoid2FbAkXxKkgmbjEJ3djeRA3Frp5tPRTpQRBeWiaAN6765tm93rpLYUZV
suPZsid+yz9L2/kGixiK1vhYoFaakdpww3LI+66OL2E4nFH/7a/tVqT9B4koldtM
Grv0tDjtl3y49DVbvN14bH46YS5gvHLfG8DBbw5s//PTCZeDQ3LHMbnOlwDQUe7b
7K51k2unuyPmMGw+ide91blV2ZqeALKeHyRitesa2d/XKap2Bsv9Kd0J9Y5kMZBP
1Mkb+1+vrWF0/ZtwuFopDKirx4tXfSOHAo1TvQz7E4T4TxSxSqwMiAeJKF4Yy0TJ
ZQ0JTl+FuVJWo3rBcCwU1w3gFCwzb8Hg0ar8xSc1z+0JP763I4uBATIadCWVfCs3
4D8cUocIW+cb1Z0XuccurtClC2ENWR+G4CHmvWXZrUEGl9iFrme7p2wIu6EK7y5v
0qRf5pOIhanXRJMZ8DLz+qyxJ33+nbxqGt1aubInRn0Pb3fGxeHy+A5cGz+tnQLy
61YDRIDN+vJ4BAwbYqcKUYvgWPPvzLKObzXV3xy3PuxUKzaJQwNxi3sCXEX5fHPH
ObnXjJhUEA87Rn/vtraF3gGiG1w7slXgA9EdzLxOulOLej49Ulyz8Nb2ED2kQO2b
QaaSbCVHr20J2lW4tO14jo5CRtGJ+N2vl/poUs7w93um6SuBmxCvxMLBUJ5EfIvT
ASLXoUKHBNwf8kJQtTcCmIcLP5Whs7rmoQi00ByBBfDmx2lfknpQa0hMDLVAqiRj
J8prDEcgt+oyDj1Xb9+vEsWfMAUvjx5Uidisgm8GKI6c3qlvDTZ1LCQXHdGZeiVi
gDmpIqZFiwAcHdmeYRqKvd+42KX2xtGzFZqW329CvD+svLsLILjNgCR61l/c0BMN
f73KOZCTlWPvItga8jcUrNxLQ8SJzJY6G1xulev5WiSjPM30Evhg2MS3wuMJQDE1
isXKOt6pyC+SVgQMGkPqKdXR5RUFet1szJK4thbflT0tskIDvpOaZrHHDkjHACBc
ayMQ2aQtwGvQxuMElGcx0pxcUzW71fH7Im7yPZp9J2X7Y0ya4TOkZF/v6+ihcHQc
5HHmYZtZtmruiS227YNVTEje/2PxfwVz5MTX2LO6164rGL2CKxk5WWj62opOBJJE
7i5x6AFb7Q00jCnlivk9wkiC2J2lddQjAP9DwJ8LSoKe6lK9KF6nZzQd/srUcXCO
4hHw3FHH3havGIf9U72BN/aSuwev+X1I6z9M+5qihjsvkLZfpIZPf232iS1otg+/
rKHYwwrc65vQewuYEoYw5mf6fEDVMhVZcUQ/b0bfKjgEs5LiPAVv7pgAJPORSmEv
JxvMJU1/LYtBhA9nEH/wtbURXMZaMQRLJstpwV1mTjWbHi6hyhRBM6SRW1i1VRf2
iXJG6q0565S4sYqS4icOaemUPr0DRt9QeCxaHH7W7gyEv7+UT19xHh0qcJ6N0m14
Cc6fRNmAfbpoeELR6ev60blHytAneXwZlIY11mFukpRp8ujUO7esWfIcLQYeBd6+
tldw51S2TKzEivgDPITzAopuTCdsuVkuzxy45Atp4tjkJxkRLKj7LT98MCTiBghb
w8xGGwPFxyX3AL4W8ZuTLuDLiXoUzuUhuAe2cDMa9bLo+9MXPAFbwDhdSDgE3dgR
KCpcaic3ZVgtUGA0PDWyISk4H0+LFJViZ70ZzeF3A6JqIsIlmtkKhMHswvGUJGB2
1MEqDXFA+tLjpgK/wh4y6y2vwCUOnY72tB4iZdXmWn7EWTO30rDEsG7CcSAVW2tE
xwL6YR6rmV2CZxLsu4b7LIJryZQ+2viXLqyxqNZ04kuMbgb1TSUwFDCRTtLKMrp2
/vV/9+4P/wFpmZ854NphnrQSL8/Ckk3YBDF++YQ2j5LBvbK+7jIzuo9NJnc2xhim
UUOQr0unFrUmmvseCV+l2TujYdmHK+kpOFG7Sa6gIK7Ddgq8orzI6fKjGCr8a7+B
MAqxotGJVKcGT+i3cnz72JGSqXqTVzsGNVw+0e1ZzxiomkA0VahTRUzKx1TfmwBg
BQX8GsVo/eBCSIQylyEMCkM6P1sk806iASEVv6VuT7l3Z/uhZ2RNXsg7DSNCNXCH
ANii9YjjiecOKNU6Yqz0qzRgnFr0WpT/4b1GqnLgyVC8VDecUffTZzdarYlwNnL5
UtMqxUGf+RsiHZeQ459/aPZEioQfXQGZWIWpj6TNrBZFT2MSbhDpKJU8O1kVDdED
tLCdJpm2TcUWrOGUBfp9dNM1TGGD0MHfeytORfm0ziiIlnWmaA8dgTbMeCiaYfhI
iyZcZw4epWGV6eI/qDTxqrT5llizHFEuoKkdffo3hOci8Nf4xIrOzPzjl2pg/nvj
2JNYnvxfRR587xYg3qxJbF71cX2r5EHaE6+B4/cOc9z2yHXSWZfE/HoNTF/XDKSG
lWfK9e4D425mmRD3nSIj83xBO11whmcohPd+4FKbmJEZ1dtU0xe+5lyRPWBQrAQN
zkQY/b0XQCnaw3PybAygiGMn2fFFFVzht0YX+4H0qRvm3hl/IpcLlVwIwSLKcz2Y
FLEsMxqcpcd6YaPaJ4csuK6juPaKgMt0rgxkKRm5EyGCQqg+vrQZnkHujf+wlN43
Jax9FHWQlacMn4wCp928JDCCkWAJNGwdjhROY5T3PNfgrCRG+L9xhw1iSo2Wtp1J
X00qhda0DcBDVBhynvPs4OaL+NWGC3vfUYuGBCYKB0cx0/xv9J+Yu5pIuPOdfvnS
pcd65fy/MaJCP5oA//MUnFmHNEc5+718YJsUf/TZv4Rd3WRJFBZJKFKr3Hno0qsI
Su7tMHTSLZlABrvG+B164z5bESlJOgsJV+cWgBLDOCDDx/u8yPpfdd6ab7R4HYd9
FDBLM3DoO1tOaSglWd2OM6v65FAY7QSlkk4yLCscGaTdfOgcq/pKuXGYfp23mGKT
dTd1Br7/F+KTTPP2UYR410oKAo8KQOaxzxy544utuS76/MsumYMOtfDOueNNT5Ht
i72FxH9d688Tvpd4bzz53YzwgqCpG3gI5Gim1V6xNjetsORKcH3ebFuqqDP8brP3
zPyoJQsLmhXxv9Ij4YuIrtwWGIBbqO+J44dE/WTQUv74hnIClLSqLsFX/b07EThQ
FSJjoHLfRYQXvFQCLs4ToSmf4HbuNMs5btoaZCVmoMnscAcsvVn1XzbChvQ406Oe
VQf8Fi3I9stKQAib0LmHpdNkqw62hLLJ1vvcU7W+D0LZuZ48CVkRm8r+LckucS3a
/T17HVG3gxzsW8h9rRQ6uPK4XIOHiIrGxhsPUCEXROKbf4Ne3SUw9c1YuGyEaYvr
eCfKmQ1ilpSAVgRAtIittn15lb79e3UI3jc5QV/gX+OQqCJrqmxZBX/LzsMdMjCW
oNX8uoJpBQq71m0ke59K4/ELssC6XB++Sz0keWIu3EbrBRSUu0rv6rFmwp7plPlH
2D6VSMYqXfuu5YwtaQC37prnF8TA8ovvqCztrDgmle1Nn/KqkjMbo8SqffREbHVJ
p16vJ/ps6+lER+Vi2Yq6lrPRCRZZ0Hfp9j1qO274PTzayeWlBDepJBTR+z1PGH7u
0i2qr/pEnDV/rstYUFi1yl4pC/Q5nqigCWsZ88RklArLOnYgH9X1amr0f3E4Ab+1
vA216vx/QKHC3UMBp7eP98axEhwQAv6Afz5bI1dq/dGgjHaQQCx71fBzuoMpeX1d
BKHd+yJKnEL2A8OMNaVDzDn9F9eroOl3ZSOHXysNRzZHwnpvqBB/RtDhJQ+hq3FU
W4oKlcLtMt3wvxf4c+CKLjqzPwAJD0TBF1vkhy7uvXDzCuwGaVjmPLUm848UFnTa
KQrJ9hyBzqp/CeHaAF7ryP94GPbHBni+01gWpeE+ImV1rJXWwVNpzYXccaDJWrB9
3IlcucbDrisPSviaSRnQF3yaN4inr4iXaFq4e3LVS1xSxXS6CSIjlCAkb8SukgHi
BALa/n+sqwcm7Pclj4wom9Xowmdblg5rU4FF3W2oA88Tj5WBGZxYvln2MMiNyNxv
wQc2thCWPzjU2waT+U/u4i+KIGwpi/feZ/nePRVBuKcUajO+mQvRHcJA0TGQ3cXV
WAcYqkPzU8i2lorTbbHmtpriqGIefHSQgZ0F0LVkZnPfr9AxUWo+PPPv1xjVLBAM
lkW2JMEfKb1tUDOOBKsqKBOS3RGH3uB2vCQEIQxQtvBOGhg5coW/lTM12sXh/QOA
jxpR9OSpHtkxEqU7b1qA8vlKqoU5LvrXtVEBx+ONLlTn38czyRhGeLTQbBIumeu0
jTqwnHX513kaySY+70gCEGuh6TaxjJ5rOG2Mk3LDryTsxrvIADsR0N7jbbhKCft8
W+HZNEa7cDdZQB6B8WV+PniKcCpXCXgG5nK0B3Oy7xogLudqnKPeAOHmeMUB/AjU
OjTDE0LvovHZEVuemw7jezDP6SQfZEQgg1xx3L8zFCWAA+vKePnOU/B6dAxEQZW8
HZ1GAqkKz+jSge0W92hwNkKhI00MpccLNVQImlJsjCRFr2/Erfq2ykpH8k/ZFA6w
HYqBcatbARB1bRaMXkujfSoG3TjTeP2es1BMEyO1FbhK0q/7BePKuHlw8Ket4a9Z
DaB4nHLqS8KWZW72vhBabkwikPRv8ZLaxZeeid/UPUWP6muu/h/en9FJ/OFQbybz
JGqJcXJ2UnK+K/wGABgmbSktHJ4AZssayjL6leqB+lpl+nNOtilOzzX5DEUyyheb
yyPJOOBWWtjfopimOd/wZQyy22NdxBeviCnqga+8r6DAOAmiT3y3NXUm9P9DsTFX
VmuSPUhlREmmIHrsTyYBYvTZ7jjxW5pa/5lb1uoTZIgMobNlAqCykIdDCSYyDraV
VufYT6PatMt/VLGZztJ0lC0pihyge+TEshHAwliUPRb1CEFpqtdbWXd9uXiHv+cA
vgQI5SrkC4U/aeeSJX5/O2mUliU084O0i4qtfTSnmJ4+chze9PFYhKCLqzyO9jrM
Svz/L7IlGslMndnQO52+mGVvmtJVmOSXlJuRfEOWrVdTSkkl0SEtGeL/fFlVkNOh
oy2XvyFfHix0sMJWoPL3zVceJKP5a2FCirxOW5ttenw6AZDeIrLoBWoKpbDDdm6O
soiU9b70MOE+Pgp7dEtqUOaxtBh+8HknfMwPLtBwl1tIuSNPiWWbjdBOVENpWlDA
9zq8NCrc0+qYaTR4YxhUzcOEv6xwvVDzXRIJF43QtfmowkCSQbZnHHNwjEgXxBAk
MuNgZ2kwTeTqrO+hVsBhUelwFlL1QOBfxEkyBI+DJuFshMpuXkOmxRaVzu8Y+UkW
/migT6D5ygaFhCRXYE3sK6qKwr0BTl5XoR/C5T9aUYUMzx+tgEkVC7a5J2P46eBz
JYNI0jDN0ZMushDCh2IsIFW9i/kZb6TrP2bymIMe/TpeNY/ItJQraONmXJw+2MEu
8fbcYUvJSvCkVs0AmgqIrO9F4+ZpKBv/jDiNokwdS8xUiJKxocqoC9k+jNLr/zKf
FD4v7v8hSVErL3xPx4zzan0KDkgB5vn+mZfenOzj9dEM3JE1LWGICI8tZpCWx+BM
Z2TusNUiCJDonNfEYH5T5Z9fxaS0k/mU0YROUCjs8BaANBSmNlmhSRQLdQfbVzzx
nlN6ybVoZBBANL8OOVKd/eGFnc1+oKZFQyzY6m7hWGnH/L5mkUJ8xCx0Ogl4xmMt
6fZJIrSjMk1EChehnptv8H3RyQRU7LqfQbvEDAnD8IScs0iXB1YW83W4nWLT7+Gg
y33oqMQN0YXFRkXfJ1uy6W47NKqKztS4dqxArtgMPyN+AAtdpVNzA7QcmksLmYBR
IzRxK1I9lSB1+DqoAyEDURMzPBF1zbr+g94wd9isDMS1/EmYbD1EjMejzp6UBcMY
O1eL5LPhz/HdDAFwkfz/7mO2YkVrDJnr2QLoeu46Jefj1fRyCzmAPs+qJGLqZ1RK
uZsNnGDHtLQVNIoE+w0FJ2U7GYKXkKWNjkkE2at+aCXI76qvlOzzUKHF9d0btLgW
wKnYt5rk9hSPYZZ0uQJGgY+AoDZazmxE9GgcqzEmbZTNOWQp74lD8a5n5cse1Tan
aBDHdNFlovi8lHOWOBX6srzdhi5otCAY3qalB0j83JbiRDn+tK56U6mql6U526D0
kV/BRPjuhgbyoGM9b+E1fhDbBmjAafzTT+UutKQMLVKuYYfnTLlTFhlUm7yaiIWJ
PzL6+B5iu6rlPMgx+nM+u+1FXHTWcFWTPeDzi91WGrddVoibQ9lAoN8okNeabQiw
pfz3a2u+PgfTNRP7eTx0SWoB0ecwtizgqumo0y60h23fyTgw/ZFdgfbMzepWU7R2
m9tnTWzCvX/s36WHjR0Mr9qXY5skTd5OT4hlEn/8rIKEBsnSENqTnMP0qemDJPkQ
WFKGkBPdnAX4Ede/oSf05d9GxX0xYgPymvJEPXECkYKxlSgI1YVoK6/NCi6WbgX9
90NvhC1WGN+4i7eTfLUmI3F9c2+1qPuy+PxBUjDRoG3FUWdnmUKH+ZWKf1Nxj8gT
1rxpxJu+cf8qxFL9TysYlrTnWwdB9XXT4AsZ1Ie63FFa6+fxXgvFwKHMghjDt02w
JjibMjdYmHFd4KISx7IDGuZaszcAYM1c30JyAsuYkQ5eMNFhNrQbJTIWmhguqsWk
gY1PafUOqV1JwKsAwXKiy8OEj48kFbIGhsj5SN7RTr70PFWyM+zWgXAfTgskz+Lp
d9BR4wUUXb6JX5T8nzxheMVqzpXJK3hnT812EbK+QeURYqHwgyIw3GvitODHJoEX
W1cOSW+OvG+jTZTTld8keKxTV2hfmaulq9CCxvLQRjUXggvO9MDccoQCSl2My2cJ
B5eS9JuYh4ASExRjk8zenDjWosV2kJtpgxCQEzkXRyBcaeBJxZm3Fh4F0uu11cbL
6EwFOiS3aSSPapwecK0VcjpCq6nyXq9c8HPafhph74RZD6clnBVXw/3n9/2V5z8X
P98Bx6zVGbUCmjeKI3uFk0tPM4Tma9jdzKfpbFawgigkMgcwS8ziULbk5CSA41d0
Q2UJFA5F0B/rEWRL9tX8TBQrIw+/GhhPQJbqzTXxi+CflT3cTO0LwmDObmXbDToe
GwOxHrdI4jCd/8P4MGUcXLZd1eb517TF7SlxGNT3Almj10VPrb/uNAFCmUQriohe
vdIFkDu1tfO5YRSQpLZA+v5McaPFuGMOPg7LWa7/dp2lU+ALfmbK+oM1b2PVv/BL
Fglj9GvyA90/h5KpmUDLGh0EmeRy6dFTJH7E0DV1p5r2+jT1TMHVoAp0YbzeKOo7
n3zqdmbXCYjHynemXOGXlIPtPQo99D86xCgDTV2uromgCicfgk+yPFHfmephidRV
+vTVQf4ji4mMhzaZv7g/DsbQHRn3A3LQuv+L9yWXyd5gLfTcjrioCU0hpc5rxRxa
2D5W9NUo/UkyExP9j/dRqDfZSgPCx5gN1vf9FR4kMFHdTm7U42D9iPspywzsWbeQ
eS4iCVGx1O+04SASjOI7pMhCr/GRjzEFud+5M/qHYPfuORyluBitZWQs11H9ZBn6
k2b/vlpxrTPwFrgHgXIXH07cqlBlyAFO9zyt1erM6zjC6yTYhH77WCQnsMQXQ9X4
JedD+Xl9U/C7rCa9pO5z7E2qRD/wlgD9L149MzaleHT3RunAlSjEmGM8e1B0TwyD
dl+pzCNS5xe2nbPVf2xzZpGtEbuE/9Wn7M53oF/WtkegZUx3Pm4hmnZR27LZPk3o
CRK+5EapmLi33zZTU/Iz2RfB86BhnSMbU+DVyILieAtThf4zQ1VLi+GwGG3mPN/z
XgWu6HZHEquqnVSi1CD2ycEqsTJhLWgFV+uLxovpHAq9MdtBp4GM8sXI+rWsGtE0
463SXOn+IwK1x9V9oSLWZM8/NzYI2PYGtdcgauGLvj7NjNC6eoVtqBebquCREZ0Q
Xc2XRd+RL5L2UxohJkUS6hnId1ScWU7IV6ZMAgkLotXg9IUnAiMC6WCduzz0wrG0
75sB2ERHfhPbliNmIZx/BPcOo9Wux7g4qhuHCoAQXxQVCy5CACyfMowtjsLmV/22
OvE3cHbeD7JkycXMSSqHxJxY1osYNlRky8nUIS1qM+Ic3XG+ISCoYxtHsCW2yHpl
016gRW/qsNbikppFLUINMxsF1N0gRjc70yLRr4zG9T8MwAkh0CnfzgU8a1Wsv2SR
8qnyk+V1LLcY1UhuvGKE/VyIFXyZFG+RG/1vnC7qAsI3Dh0KwKhZuGqr15SFKAMl
MnEo7v1lNQgmx2pzp3TPjHU78V24KrppaMGVqSBJNz1ZsJ0UD5xSBsrOUCZ0RFPb
x7MCTjYBCCPuxT+YG3B6Qrh85jMElrKtumeAZ7wYau3snClHm4L27ZKHXQ1Md2TO
Eatv1EP0A8w2pR1xRiC2OM1eVTUFL6ekkuGaiq9WiZWyRe4Ns18pQMjkEJf4J8Bs
Tk6lnZVKIFNBYZdSN4UUZIhc0pMjxX56TxIdL1qVfm+PzRGn0modVYPPTqNH6fWn
SrZvm3TtvT/LMEW+SyBTAbnEBiwFWZqx3EPXZZ387ZuESagpcfa1zg52j+hukau5
rS9+D/9GOxyj9wR50F1sUeiXiEVzhEVoYQYdyI7IRLufddWZUS5/lpeqQsEFm+Bg
lQHV2s0zn/hobmwZJUxni7jDaOsziUAL/yMqGMFIS3+NIR9Cv76ylDKv0y5bVID6
xdBvjkSCPNxHa8aK+bn5+832OIqVzXgssZnd0n2XGf/yS7E8dtE73zx/BWypCfPi
H1n7v5aeUM833UsgJS/Wr9knFbD8WqQUOW/y+2OTAoFxzpQtiXDG0cJObd4k4ae0
Ax72G/fyvJUrGqnC/lWWPLBK1CtHLLsB9/v4q8ATuTokOjU+56o4c1oVjpfD/h+w
Y4fTls5J+W86eGmo9A3GC2QFMYJwlErJMAeZco7YTYP2j6SpIWuZwtifY0zGU/Ve
p7Dcgrf+56fVmbQguIqsl+kXGdJFX9Hf0IeKDwh6IW/tF2iaXZEBRrb8IDqfiFd8
TnidvRvKOVWEWE1fDvFYX4nRvLNXK4FCGGxCvq3BUvrQNXOz+ge2yOwLiVPWehV3
TYxQDTr+4v1FwsFAJQFrJtSbJfDrzG6gFoAX8j74ToO0p7RCGz2TK/6Y3UACZIPL
ngpJ9gBtWiiLPdX8BuOF2l0VKDjGrGa3QiBD1v2/W1JQ1KljyEQm/6wVLnoipORd
WqPsRHje964aqiEyvFHIAMuOqPZizDqpH+di2BXOKEpmScK9a/zOJXs/eUCHX2wQ
L6+i63h3X2N2FEqlT/gQBrR7F2zHJVdJC3Pph8a/L7B8yHrIJ1m7AG5plK9zyQhd
dSylJ6gquNCWKjSJ+fEA0lrfCpCVHeDi/KGus6E8oH1smdvMcAykS+wask5nyJSV
03P9Ddl5eOoPIi1n3OfSn8Lkff/RJmB91FNE6uyHjJsmJsuuowfMH/0fsSW1oltY
t3mUBJ4CzPdJ3KDdzK1H1bmzz0o9wkCcLZJrnmu5l7mM/VW3q1l1WMr209c1XgbW
sQQVQTMjBrybPEJV0mdqJ69HdmIwnkDPMJgu4Jb9HlJ/umsqtPNfBgc1oicKXMeE
Qt+NV8+u1g3hZoIXWFa03rroAx9Ml0Da226/aj/mj6IRnrvX5+suI3SsSdIZGwzL
ihFRVSnXeB47CQ4QbdW3Klbc0Y+b/WexdhsQrzp+Ij6eBKxOCmO7B/VtKlCKH2Db
wOVXI5VhXrtBNUkypmvARVNd410wrohnHZfmTUKFniL25cHBxwla6uGMgc1a0BMi
avWBs8rq4V+1mg1CmAkGm6qBLUuXv74mkUySS7VQKmehivGqGOyovDiLnrbcXb1a
MT26PdlUZiBAzNIVonOpKNjZ8P1to3LvkwGnxyAMknWnYcCM6iaGIXsRxdGnLfv8
MMtdIbdevj4M/iG9KoW7CKf7wbBIojgYucgmRTg0jEpsUMz8Mhiv2iVSWFGEXm+a
CQTg7Zx4+jPLhiEs9kHPSh25IzLYnzuq5KM3UMLKppAP7zpOnOMK2kziwFAnsjye
mGxW0KKAzfA2yTos8pqoQRsuCzEvD+jmjn9tq+jsAylOZHooGWQh+9YCqu/oRiRm
kw/3DilN3oG4WoaeSE47SCuEJvFVU1yzJJSw0Sdkvlf2JhAK2J/ifDP9zWqcJoey
6Jk0gMxxO4TV7YiO/a9QBPgD/izuHOg5pTiEH2kdzf4zWfqFsZeraP5ZCkuwnmu7
jGDEFVXfsZ40g6ZGDXrzmNlyZalTGVK/L8XRU1RYNXR0Cq12p65Opyw4sLbb8Okh
jjZpkgpx8s+y0L9Zip+nQMUqmIcz0dLaBF9RDNd2BC1wZ7Oe4PuhRy1+l0PxRK+a
ySs2atPCTVcBgpjdBDw0B66GZ6mR2c+Gtt2lqyGe8S4SsQJDEW4xhwZKObA0j6E4
PZD20qlWq0sAtL8RFWWReJBIeNpz4fdzdAHR/Ct5Pk6egXzev2CjJBCUyHEMAQ75
sclhZX5bbOa8yY8Q48e4B0zFp90J1fXdw+nLq4fEhKiH57f8/RnTOWcHzdjl/SmG
ry2AmDJGeTYVISKybSBwD4yv2QtibxurvgYMjupkoMUdtYXNcZHfHe5xX1TsvymF
wtXD3IWP+kMpXZSOWikRgPd6157RSpdy9gadjCfXQ0YootwWPXUuTJfj6ei1Kpfj
LOHgMuuEFoEXmyOWBd5P23wKVVPFjBCMi8n6DGCpTUdydxfGRGWI84QlgoNIUT9b
Rak13Xw/tDlzZCom3m74bi7ME6g4v7Tg9lSKBsEfP2rkVZLH6YbTktZd0xCoBCPe
pJmlhAViJ30an+nx20nbGNpxq4XDakJNouXSOk27vFQ5oDHDaKALG8psHHqUC6JB
n40DTdWYdMh5JGgQliucBeaJsuLhaEpo3JqB4cFODLcfjskzOpHwH1m8tzS0qhCU
gpkjXg0TkU3V15YU1wUV+02rXkBm40WH85Cnif4qDVuJSX5Znb5xTtX74pLTixNv
OCLQ/otRis/NXkE8/vGJCxKpHRBISEoDqgMfBil79F88dK76QOuwC5fDVh78yVRe
e6PRNbckOHrq5LXJInFj2pHw+vEP5gBGQOe5COBBL3rnzbTwD/z2vyz5eQizdpEt
nsJcLuKbxzUSqjJE/LNetbJkEXa8KN9FdUKt9UKGfxnrK0G5r9P8Sfdk577SM3wH
vHecZo/MX4EG4QXpo98of0Fa3XGWoWym8C8Jkr4qm/o+Rk2XHLfdkwUGocwVL9YW
1SdEVKqemtXmzeRtJhUjkV6YStVwuYojT2KtOvwoGCLIIr6FjqH47I8LlfmvY0g/
9p5j5Rk8MjqtXLPNBw+TL4BpubVbzaxMQqfA+tMV/i5HC8mjs6l1a5DdzPna07tF
2Yx+4wzYlynIy4hRosteCZ9binUrKJB3yTGmKt70uyxP49ZYaKGiZnCMbLicOhb3
1IgxqaYbSI/3+nCpY7doX6jWZlhMTUO82I/OZiOcTFkNW714aqvA05rTCDqs5mBl
RH++EoGw9242MZgMdk5L/clA4YtYmZtSATIw0QRG1rm5k0Rc8A1tjio3OUxyVsX9
4ONdt12/j0HASCz48mFZx2I9KFAb1xexBxN9Z7Te9OU6bZInSv0Q2Xo+ElcIKYaB
AQjZye8YFCoKN7AKUE7TvFEn02DNG/2ri3n3mYqVnzuRrrbidGqQi9Mf9MkOjL3T
oLBO4xRq0T8LNVCda7QxFWDoOrgvqj6oY0EFWD1x9A/8HcyNlC5hk5zVaO5zJMpY
w3nbuimVLjpPqLsKLkCqKM+yBmj+dqDAqEjz8YwEnrS3nKKRuVdbOmUw5gqCx0aA
xnq1cj8kl2U5ao10nI/Sy61Lk08UWYV3z9A/7MWh20BNzC2PuOYQOpnGJF77CkcQ
1ikA6iy4brJUQ2UnXX5r6UNE8Sqvwiw41CBWuJA9M0TA4Elv9mElaxBku6bRVypr
LF4L3QzmiLCh2ir3VmaPG1zoAuIEoKucLV9Cua1MgRXVkr/LyijpWKzQ8CcUjso7
xJeszUjN1xbB3tVueJmJvsDlYz67UKbrEqgeMBj5YVNlLv6ALiD/gp5jTnAyKood
FOgn9lJK652Fc2TjT56Jh+PzUVQHqXoH3C+cytDIR0rjc0RPEvtIw2yPi37MMoQS
gGNmrflUClnvNN/fv4OzuWAIVM3zh4b2rtRX7zqKgakAn3Ckm2pWiwU4Jx8Y1XFS
HYELd1bGKfhJMkiglbuUurJW5QvjxO7UhG7FK5AvdHzMnupknBSpWNxU7fPq7Knw
vvj6Zr931zuCwnHWisddfokjpjwHyhDBpSiNbRi+Nlx4/y0xR80muafEU+d/LKUi
QmNvb8YkF+wRqRo3fXfBUa1Io1oIiB+U6g3H+keG1aF185aItYOu8+kJCpOM/jxX
fbG70+kzl9BMouD3+e+N7dxPLPYczQeqrhv006qEWwWKypQSdQlGOZS3szvXpIJQ
rV8SRrNvoTudhZ0AhVW5bXbhdbtoydaGRoyiw+k7NGVmSvZTU7fXLgv+0gXbZG2T
k5pigFzCz+8KFfsTL5F2hjJff02860297PZY69qxyyRK6zvalxXRcaiI+SoIvAPN
dBu6agz1CGVWcp/48C/cO5QWjgApf4EzwC9yWedTmcitl3DWgucFyFsxEW+DK9RX
op9BIGoRwWX5i8WNPdqnTZcmVJLyNpp/RNrYTbFhaJEfZw7UUOjB1iOxOBpZ5xIm
feE9o0TLjNdpSzIjGOlZ7E9rfaL9uIeiB2kjd2CrTRBfINoN/x2THBtGrxbU2q3R
CWXQ8UupXpJdg9GrTpNEt+Qe9f67yUvC7edqpMaUcjv5miKoROVdJtq7ViNuW0tU
u5DfqDfFzl3XosE/La9az7VcboWr1TAQYQOIvQnZxFbtCQyUEUOBkq4Vb2U9XdfQ
qVoKWuiwFjC1XAWRR9YyN4DYFf/vBWD8hCl94JTHZ6UNPGgCgQ3YTRKIBjwWq2w8
XLl/TwoZuDzvL0pRKYeMrlBCiWO6K2oEPG7oAg6dxWXIvYQ4ZgNNEj8f2J0JZ5iL
vskXpasyNRB0sd02tsdTIMBqChw05tA9FmchqJFO/UL1k6WrGJEyCB5A4kT1QAjE
wkA370fkI1yk50sV1KKNtAKIYisWFPvexTSQeFxHPRdd7zPOcF0CQ+Lx5O0W8vgR
Lg+QUcvnQigX6IIYVj5Z5vxPmibmq7FXAmWD0IpjbQtWgrNWfPoRpjZNDUomrtjS
bN0KDcvNgkDKtrFGD9MeO8ag/cg2QXgqM711L15Q6HbYRaMIQmeKWk2VUH5Sk2mr
uy7bdMPVMwWPIuDQ44wbKbTkOZ91zZnIqpYhp1hNCd9d60HGpK28aXWANwz/AGwb
XCBJva2d907Vh4Humox/Zx23TFte9HfkFHPAeuk5pTnw6qNNnIt3RWHOiRiuDcG2
a4LOQpUriwEOKin0OnbjkUJ90vajFGdeeh8pKdawo4sYn+Xt9NlpM9aMR2edPDuv
fXfYA6ylME8lIoSiCHH1+9bmzm+4uQU7Y0uKNCld7qLUriU5hozBvoq8VxNlQA2Q
1GWgOGsZDtN84uqS9P9sc+3MzW+txIEe69kzYXOKrXauWfTl4MUEo4PXp1JWufjE
K6zKD3fzo5WTKwfEj4WHhFUbcodMGiwh2Po+MBQYxTe2flFGLG6NlKIzYs5+xQOB
088FwHKFfXFtBwYtc5OMSb6TL56hPFfcwUEIRcmUUlb8k8fGMhq1NfBCExy+xC5x
rtZ0h3UvLz2YpWHFYDrLE65uoRgUR91WD3GT4Pg8tu+JjGcP4iZ4dacqDVlNc2Zj
aSfC3gPtTpw535GTIO56hRQeC3T4+jNp2yGbrd7Pcmvceu/N00CW4uAJ8v/0XUvk
58IlhyF6J3kO9X9uQIRvX5RoHObKGdW5/ywya3LL5uV4zhj81vA9DrvWB1EDFJhh
enpH6vuNycKB5ZTmqFfdtWvOckGIuh3UGSl7xmRyF28TIuw1StjXlovPQDtfz8JR
YJ9kjep5yr6iSwO0utnU6NhaAmB6nC2F4qQrB/23i48TdfUrtPABWGDxDOyvqCqw
NNZxIB0Rm8ICOlatVMK3lw5x6G2k15dLpYuIjNksyyFGLViPFhhBfpzg7DcqFw8e
vlK6v/xV8a6onYwgRMViaFGt8g1qUvcJ5cZofyuqmpmErFuPgL1Eg+xLvRHXSxFU
T0pbozxoImk6gkIroDJbXCC38aa+cMH7lxclSeynOfFq4KVrw5Ozo0m27rlGD3JH
ijFGKzRB7/kNsUF2AzwAFRhYzN+ZH2g+grPQgqTwOINsiqEwLqnKQJjJm3yoirw3
PZIirpo5PPsxYLLhREM/Q9DRI4tCpXJRxQO3DLIdUA+djjJg1NaLuceHjVRqOuwW
pXApVFo0EgqIln2Im6vZsjEZ1MbY1kcCg8jzCKoETsm6jdeEjeCHMKFT4NT8pvVs
zgY2YYIPkPkgWsO30BkDOdqimvtK4qiTnHXSLGnud9Jpj23S8bryq8maCdFFPomk
q7P0z8omed5KGjOSWoF3H8HyILTsfcglEXj/keKH0osEKl9tmfjMJLZBJYkEhgxo
f0MrEm0Fs2sr8aeRwRzXsPnbn2KzB29t5PC8Nxul83gnD6jbLmM1Oux3XkOWpop9
4p/yu42KI47SRrDuldTX03mkq5s/DRNvZgnCarLxlHVQmBDt9A3Nk9nST2bpNuyo
PEvGbGGovD1cIO5t/A1vyoObgXsyNtT4CqD01ahr0jFa7qOtD9blkA+3lXaeoWH/
BldcP1Za/Mfue7/G4jjHuTjd1PqjUgHJ2ZsxRckwihft6437deIbxDRSxIsP1JXS
fR3vtbkepJugGy9IBz7L1EtFNTpnNSSzAxisYEVdmoP2lZxzdR7Y8i42HJsLLuqk
KPa/giN5QvsGyqDdp8/Jf4gFwTFsGWa1mC938pOeATrhL49/2Dr+kz96n/I+DeTi
TvJ9AnVmOcKJqpJZWEpUjmg+yfvF6XMPTV6u8KYsP4s6rYbKyqVRSnmbnwwnS2UN
tl6/RIQnvOgA/nvKaJjRgvqfUvV14/yRjCO8nniAEefwFoyIwTQHqsgMe1zI+FXv
bocNpucJKg43i0UqXmUIZuE9+3Vm/tPfjtJJAzYAsAuEbXvliRIiYFifcSJJ02+9
QcbUmiBjdwvsIFNbPnvZNoh7HyJmq+4aX3NmCpGNrCLVvcVQfI6PdY+skpBktIrx
rzO/hSSJkD6JMXXhrnchJ6HTlIxRYlvvAFZGGubfl/puhz449KzV0VnMBU451w54
53DujzYhTQj5bPJGhcJwOKxJAMOGQcmhbrxVXK9jG4VVciklcZxY4CMzV4RNeeyZ
xinTMHGKubYBVq93g7Kdyujmo+tabBL32GwBILZA8ofX3N8uNZ7bgpdWcA9mdYsF
hQFBtICB/HtkIKc2co0d0RlAZx4EdZNhB8MiIDElJyr58vhR8S+DV6BbJ/s2ORLJ
vsvuUAJSi0znk3AQ1mOcpYNQv94h3EJm67xCB/zC+2opg7pwaLq74cLNzu47OzpB
M36plEFEfq5nOmTe7G6L4THLfQfdrgNjL36hVQXd7/WW29A6wRC0OzGAGHTje8aO
RnNc3V7MFGcHznJ85YBE0xt4d4/0flblSQr3cxp7uc1nROS964DwTX/wyGWRNeeZ
+wtWgGVzGQKQIzF18Ms/3LneaBm14FkRveQhJHr4dOqCIUhvBESv9vQrLT4Atiz5
LMAVp25e+1Whv3Zz+s0BJSmNoH++OqGmklO5owSaQoT9VruH68xTylUWODmTk9Sc
RIPLQoNMe9uhrfZeWmhED31PUSwiwrAXfEU6zxZf1lbbxMl7fh+270DHCo29btsS
ptk8DBxNzCBLr2mbZMXmm990FaKTJfIAhDhvq3+tIEU2Y+525FQ7cCRZ1IoW1X/6
bbr4pVGI0MejGAIlt3QpH5gVp7SolaAKiHMRd0S6RQ/egPjOd7Uf3ld4MMnuDkjF
YQacDz3WYHnFnhPhKUcAelw3FECYkHOMCv2b9Ayk/G5U8tbQ0DdumpH3xuceVszM
4QnDHQh0e6vzTfc4kllXZCICYzMEnGIIDtWwhZnqoYsewfA+Fpz/BPxXIyk4Bglb
SgjL01qd6loKTcc43h1p3PHG+b+MmW37BJImVr8GI7BqsZtgDNMvsKonGtqCOPzf
gSITa5WUoI/UOpK85X9zZ8j3ZzN66bdzEse5MKwmEOxgB8MaZu1YLU2bopGlv1+x
CNNw1zt6ohkV0UJlboInAK7xiq9P8slG2nDUGj+s3k4i4icJ3gU576h1r21pT/Kq
y57eA9Q6kov6fQi+0pJjuQtg5eJhJy+4ZPKDTECLjb7+Qs2pg2g8mu3C+TCKxWdl
AsqnFEOMw68SxIf5Fh8A2TJFP+dYSQQysJ2+USXfBm//xIGd+Oo/srTTXTkCNd8e
FmdA1eWcV1IfraAxy2Uv8OGPJwKXpn05jF6uCYMpv94MOJbrLUJRT+8NKB2mWCuq
3Ylbunb0lQdlYF4Rc680DYPsXSAkodhUMcKExhNmJEyK39DbIvLKLrUgxOXtKfTd
6gasaWaoP+wNzmYTmtz2bXLopYDwg44BsHblRxPEHuaJ4xCiA5MfG4RnBYAiwmDj
rT+qbnZrfFOGuPmS89nNaYYcHoVEkw3YyUY4I9rkhvGq8Pui92CWfA/REEUKCf9F
6+brgdOv9pMsaYcx/nNGt8sB4AjWXsYcLqiZ8gNNTCy0QFSHiWuaN6FHCTnf5cIZ
99ArHjRo5qZItgcYGhBFBHMNkOEr/E3uagzdXxxPKAY6GWoP1dgZXCm/1n6orLoq
gR1EwMBln71uPX/ZaQJq01Lp2N4dz9BnR6eBzqp8TOcDqVx9EkR3K4oVLl8Yauef
20xcYUuQfsu7O3xmxVBqDtwcUZLZ34BMR9IkMLNWF0D36Bec35vxP2kRprRxTflJ
Xyzf7w5MBv004KrgAu9hFtDl7cl/K4rUIDNEVZKwxVYsWdg5Qf5sIKS3UUa7pI6d
4BrVK29EoM8WRSKOzyvmJcWjibJE4dw/upNXlBnl1/zLuw4nAb+Sdgh5XSidUkK9
m4GcQ5RsXYwDZFkPB1Bv+1J6xcs2QBctwxxyM6c6o7LNlLOlFlDWnGcMXQ/rJy4h
oE3PSXEt7zKdNnYjbxwvNiAeXPcHMtp/YjaVg3QbTYWuhNrgoFeiZiFryhkZGN+S
f1s3HoMlqk+R7/Gez21G7SByRJ0Ii1BR2ZepOSL5OQdNzKhv0z016yiiDR0HPEyv
cXbM4Gga5TjuaEsZYVRvEfr3E0Q9+bJ/GDKDgbR8qhjHXgYMrLT/N0Wctu27U1AU
jIaYJWE9udZsp3CVMtvrECp9pbcuS8gFeWjXiQvDFMuY+AFl8DhjBqzshOsM3+3v
pOd+xnybgjWQziYpPGCENbfkON5Ibl6wacO3MDd4lPFa1qtarQSkUuOMGoc2k7EI
QSrMIn3UWuk48MYUtqkUj88khXn/rB7vsIuE0K0S3wyzkZuyBDb1kDLUsvH1arGD
u4HsufInqafysNWM4xlH8F93c6Nqo+E5xAC9CLQmO3hNjwAmmYz55rCfDo2fazPe
bZDK4ZFT5cUuN3XYjNnXGXt5RE+ZuRbPwC23a/++FOLuwYDi9FFKHTLhzcWzh8Mv
P9qXt9/JXk0D2IY1BqFM4EBRT896eoWiuny1KdF1I04hAcZeQJ5pCpeNP+gWwZsg
qijvU233AW/9hKd7or8m2hJtpL/AVHIUO35DDA9eUFBGKnpyf3mjzIkB+lKu2nSX
DkQiyxwvaCLbCYW1QZ0ZcPBMIxj7BxceauY5Xh/F+Vue+yj/nnoSvuDT0p5IhFZ+
SII7tjCE8o6Kl3z2XYb69HjobhzCTBmJBio5D1mZp/+sN2uVi+I4FBXpAfoYNqTQ
ILc40jLz3bzYz9/3Nwn3o88LR87j01x8aC59LrY4WqkhAn1Xhdpkath796pJ0j+a
pDhWz7yvc8tHamdPRuCwnnocBmWD5eGYvYvtJQlOfcpco+n7pW4Pn9yLMJXU5qv7
hc/0NFGr1LOiDkmg2IBPM8TIkvKBJEaAnNAMNW164i+qGG2/jUdpTsJ4uFp5xQ+P
YX2thXDlxXxRbXYL+9fz25X7boEkS6hKRXcDcoAJkt+fzMAFF3ilcZb+bf3HWZmX
lLUhwNvXbZU39XRtiv28IbJmptHzFei7QYdNhdCoXp+JcAn6H4hMno2mu5kz6kBd
SoknYTvwsuH8XfSijvB3VB5xKGV5c4z3Hy7v3p9rmXtzuqRMY5FQSKXyZXlCH4Ro
oN1hZuhCOxMez5V3vGNVB4g0DMKaHUV/m9ud1A+XDCuwqXF1M/oBWJL9lZZ9VDLE
Wcg4QToH6W37gwkIjIgEcgXp++9cBF/cueYQE6zsR6q/x3vKqUXHmOyHWDDcXpx7
z8IRsuS0ETiWL4A9+WQiqjcizXakxNX3iHbrnulKjqM9gKu8zCjxCOh9OLeEUpTC
xZFCHdcyOuFaUHaYLCJ8uOrgA4yO8q1mxrmZwawuxHW/5Wvq9A8v37IUmGUw3/iW
AK4tc8IKDs+1K4mD11Sq/eauAWuhEZaN87s7j+AeYdmZ2utjzkCyE0aA/8FyHHgT
7fM8dLjkA3WfL0kADfLNS0hIWBPeGLCk1hZ+zlKm5nMFyYtlUxnfP6y1MukInRIb
qaN18ZlqaqfuEcGM2JN3bBay1q1B7M4iyyu520yEzU6QDZe/czx7FXeDda9zV0B0
18RgKKZJyNJLosbRyznK9iv9KQ6sQxlxnVwLrR1hiGWwQ1MIqNtN2sIzU9xRqZUL
l1NLip0ft1MEiwW5Q5c2V9SjJTXItYGTB2txFnSSTxz/SHi6K9oFtSJTYpCFOEfV
XMQ1hVzRhARoqII03GHnfg==
`pragma protect end_protected
